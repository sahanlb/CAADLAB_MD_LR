localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTY_CHK = {
  {32'h41b84144, 32'h429c8b2e} /* (31, 31, 31) {real, imag} */,
  {32'h421ef9aa, 32'h43170863} /* (31, 31, 30) {real, imag} */,
  {32'h419d04cc, 32'h43126c82} /* (31, 31, 29) {real, imag} */,
  {32'h415d2832, 32'h4303574d} /* (31, 31, 28) {real, imag} */,
  {32'h3fd8a854, 32'h42fbc35e} /* (31, 31, 27) {real, imag} */,
  {32'h418082ad, 32'h42df4762} /* (31, 31, 26) {real, imag} */,
  {32'h422a5a2e, 32'h42fd44d5} /* (31, 31, 25) {real, imag} */,
  {32'h422ec80e, 32'h431ace5e} /* (31, 31, 24) {real, imag} */,
  {32'h41420e25, 32'h431b9a4c} /* (31, 31, 23) {real, imag} */,
  {32'h410eec99, 32'h42fed6a2} /* (31, 31, 22) {real, imag} */,
  {32'h41061cb8, 32'h42778c03} /* (31, 31, 21) {real, imag} */,
  {32'hc24dcc36, 32'hc229ca6d} /* (31, 31, 20) {real, imag} */,
  {32'hc28b386e, 32'hc266187a} /* (31, 31, 19) {real, imag} */,
  {32'hc2665d5d, 32'hc271c469} /* (31, 31, 18) {real, imag} */,
  {32'hc23e4527, 32'hc28f2594} /* (31, 31, 17) {real, imag} */,
  {32'hc24c0b07, 32'hc2bbaa91} /* (31, 31, 16) {real, imag} */,
  {32'hc190d2f4, 32'hc2e51a46} /* (31, 31, 15) {real, imag} */,
  {32'hc218614d, 32'hc2e61019} /* (31, 31, 14) {real, imag} */,
  {32'hc24b2984, 32'hc2f9e394} /* (31, 31, 13) {real, imag} */,
  {32'hc2061259, 32'hc30826b4} /* (31, 31, 12) {real, imag} */,
  {32'hc187b659, 32'hc303922a} /* (31, 31, 11) {real, imag} */,
  {32'h42287f72, 32'hc1294f4c} /* (31, 31, 10) {real, imag} */,
  {32'h42ca9c10, 32'h426a182e} /* (31, 31, 9) {real, imag} */,
  {32'h42c21df0, 32'h4218fe56} /* (31, 31, 8) {real, imag} */,
  {32'h4287b874, 32'h421da96f} /* (31, 31, 7) {real, imag} */,
  {32'h4218ccd4, 32'h4262d55e} /* (31, 31, 6) {real, imag} */,
  {32'h41f2b67d, 32'h42b7ac64} /* (31, 31, 5) {real, imag} */,
  {32'h4216e63a, 32'h43067489} /* (31, 31, 4) {real, imag} */,
  {32'h42019c2c, 32'h42ef828b} /* (31, 31, 3) {real, imag} */,
  {32'h420633a7, 32'h42ef28d2} /* (31, 31, 2) {real, imag} */,
  {32'h41ccbd27, 32'h43108882} /* (31, 31, 1) {real, imag} */,
  {32'h40e97085, 32'h42b8c586} /* (31, 31, 0) {real, imag} */,
  {32'hc196be52, 32'hc25aab34} /* (31, 30, 31) {real, imag} */,
  {32'hc1a6fa74, 32'hc290eaae} /* (31, 30, 30) {real, imag} */,
  {32'hc10b8762, 32'hc2a83a69} /* (31, 30, 29) {real, imag} */,
  {32'hc1a46e1f, 32'hc2d06674} /* (31, 30, 28) {real, imag} */,
  {32'hc2049e5a, 32'hc2bbfb78} /* (31, 30, 27) {real, imag} */,
  {32'hc15e47d8, 32'hc27dd97d} /* (31, 30, 26) {real, imag} */,
  {32'hc18ccf70, 32'hc28922f7} /* (31, 30, 25) {real, imag} */,
  {32'hc2131943, 32'hc2ce78d2} /* (31, 30, 24) {real, imag} */,
  {32'hc23e8b34, 32'hc2d075bc} /* (31, 30, 23) {real, imag} */,
  {32'hc1a8b0fc, 32'hc27db5cf} /* (31, 30, 22) {real, imag} */,
  {32'hc1b3d17b, 32'hc1455c01} /* (31, 30, 21) {real, imag} */,
  {32'hc2117aca, 32'h42bf3025} /* (31, 30, 20) {real, imag} */,
  {32'hc1da3596, 32'h42e4cccc} /* (31, 30, 19) {real, imag} */,
  {32'hc22f2632, 32'h430489ff} /* (31, 30, 18) {real, imag} */,
  {32'hc205e2b0, 32'h430853db} /* (31, 30, 17) {real, imag} */,
  {32'hc1e3b001, 32'h42e74e52} /* (31, 30, 16) {real, imag} */,
  {32'h41c7121e, 32'h42a98dd8} /* (31, 30, 15) {real, imag} */,
  {32'h423b7a8e, 32'h42b66c97} /* (31, 30, 14) {real, imag} */,
  {32'h422009c4, 32'h42db15e6} /* (31, 30, 13) {real, imag} */,
  {32'h42246dba, 32'h42c476a5} /* (31, 30, 12) {real, imag} */,
  {32'h41e283c3, 32'h4263cafb} /* (31, 30, 11) {real, imag} */,
  {32'h402a72a0, 32'hc21f03eb} /* (31, 30, 10) {real, imag} */,
  {32'h412752e8, 32'hc2f25087} /* (31, 30, 9) {real, imag} */,
  {32'h41e3d9a0, 32'hc313f1fb} /* (31, 30, 8) {real, imag} */,
  {32'h42202803, 32'hc30df5cc} /* (31, 30, 7) {real, imag} */,
  {32'h41f848d0, 32'hc2f0f6b8} /* (31, 30, 6) {real, imag} */,
  {32'hc197c372, 32'hc2a8a05e} /* (31, 30, 5) {real, imag} */,
  {32'hc22649fa, 32'hc2b9f17d} /* (31, 30, 4) {real, imag} */,
  {32'hc1ceea9a, 32'hc2b2913a} /* (31, 30, 3) {real, imag} */,
  {32'hc1e717c2, 32'hc2986ed6} /* (31, 30, 2) {real, imag} */,
  {32'hc1c09834, 32'hc2bc85d9} /* (31, 30, 1) {real, imag} */,
  {32'hc0f50d38, 32'hc283c5a3} /* (31, 30, 0) {real, imag} */,
  {32'hc0ef184e, 32'hc1887645} /* (31, 29, 31) {real, imag} */,
  {32'h40f9ebbf, 32'hc11dcb0a} /* (31, 29, 30) {real, imag} */,
  {32'h4149c529, 32'hc0706db0} /* (31, 29, 29) {real, imag} */,
  {32'h410483e0, 32'h40ff0f34} /* (31, 29, 28) {real, imag} */,
  {32'h4082db24, 32'h411dd578} /* (31, 29, 27) {real, imag} */,
  {32'hbfde363e, 32'hc0413e52} /* (31, 29, 26) {real, imag} */,
  {32'h40381548, 32'hc1d5397c} /* (31, 29, 25) {real, imag} */,
  {32'h40b5bfa1, 32'hc0bf77cd} /* (31, 29, 24) {real, imag} */,
  {32'h4118829f, 32'h4108068b} /* (31, 29, 23) {real, imag} */,
  {32'h40c4a370, 32'hc1377428} /* (31, 29, 22) {real, imag} */,
  {32'hc13f4ccc, 32'hc13c1883} /* (31, 29, 21) {real, imag} */,
  {32'hc24d58c3, 32'hbf3b9010} /* (31, 29, 20) {real, imag} */,
  {32'hc2400e24, 32'hbf6775a8} /* (31, 29, 19) {real, imag} */,
  {32'hc25b540a, 32'h40cf3f95} /* (31, 29, 18) {real, imag} */,
  {32'hc2166738, 32'h41a075d6} /* (31, 29, 17) {real, imag} */,
  {32'hc248a0fc, 32'h4134872d} /* (31, 29, 16) {real, imag} */,
  {32'hc1eb8103, 32'h41a2b421} /* (31, 29, 15) {real, imag} */,
  {32'h40a71ad6, 32'h4138d66a} /* (31, 29, 14) {real, imag} */,
  {32'h41f90dd3, 32'h40b4693c} /* (31, 29, 13) {real, imag} */,
  {32'hbfb64978, 32'hbf85ee40} /* (31, 29, 12) {real, imag} */,
  {32'h40b2a7c2, 32'h41264c02} /* (31, 29, 11) {real, imag} */,
  {32'h41f1a839, 32'hc0b57942} /* (31, 29, 10) {real, imag} */,
  {32'h41db6d67, 32'hc2041e62} /* (31, 29, 9) {real, imag} */,
  {32'h42841cd5, 32'hc1fbb6c3} /* (31, 29, 8) {real, imag} */,
  {32'h429dc03b, 32'hc126d68c} /* (31, 29, 7) {real, imag} */,
  {32'h424d7ceb, 32'hc0a40e34} /* (31, 29, 6) {real, imag} */,
  {32'h408101ec, 32'hc1a24f00} /* (31, 29, 5) {real, imag} */,
  {32'hc10af819, 32'hc1a09f9e} /* (31, 29, 4) {real, imag} */,
  {32'hc16771e1, 32'hc08f6212} /* (31, 29, 3) {real, imag} */,
  {32'hc19cd39c, 32'h412a537e} /* (31, 29, 2) {real, imag} */,
  {32'hbe76fe30, 32'h40802b16} /* (31, 29, 1) {real, imag} */,
  {32'hc0809e1e, 32'hbf3fa12c} /* (31, 29, 0) {real, imag} */,
  {32'h417dff7e, 32'hc0b7f397} /* (31, 28, 31) {real, imag} */,
  {32'h4181af8f, 32'hbfb9dd78} /* (31, 28, 30) {real, imag} */,
  {32'hc175d663, 32'h3fb9fc50} /* (31, 28, 29) {real, imag} */,
  {32'hc1ad4156, 32'h41880d6e} /* (31, 28, 28) {real, imag} */,
  {32'h3f88beb0, 32'h41fa3950} /* (31, 28, 27) {real, imag} */,
  {32'h40f00718, 32'h4209bbdb} /* (31, 28, 26) {real, imag} */,
  {32'hc0a4da7c, 32'hc0466b54} /* (31, 28, 25) {real, imag} */,
  {32'h404ae768, 32'h41808fb3} /* (31, 28, 24) {real, imag} */,
  {32'h41e0838e, 32'h415c3074} /* (31, 28, 23) {real, imag} */,
  {32'h4264b70e, 32'h417575ca} /* (31, 28, 22) {real, imag} */,
  {32'h41830f0f, 32'h3fc19d20} /* (31, 28, 21) {real, imag} */,
  {32'hc223975a, 32'hc20aa884} /* (31, 28, 20) {real, imag} */,
  {32'hc22da810, 32'hc1d7a294} /* (31, 28, 19) {real, imag} */,
  {32'hc215310b, 32'hc06ced88} /* (31, 28, 18) {real, imag} */,
  {32'hc1a8012d, 32'hc1a1d1de} /* (31, 28, 17) {real, imag} */,
  {32'hc1b55dab, 32'hc1dbc16c} /* (31, 28, 16) {real, imag} */,
  {32'hc1adc1aa, 32'hc16bf6c3} /* (31, 28, 15) {real, imag} */,
  {32'hc127c946, 32'hc140849e} /* (31, 28, 14) {real, imag} */,
  {32'hc12af2c3, 32'hc1cbc48f} /* (31, 28, 13) {real, imag} */,
  {32'hc1c8d82f, 32'hc1e0ba84} /* (31, 28, 12) {real, imag} */,
  {32'h41188ee6, 32'hbfcdcb9e} /* (31, 28, 11) {real, imag} */,
  {32'h4207f3a7, 32'h42311cf0} /* (31, 28, 10) {real, imag} */,
  {32'h41ef0d40, 32'h423438c8} /* (31, 28, 9) {real, imag} */,
  {32'h428a181b, 32'h422bfbf7} /* (31, 28, 8) {real, imag} */,
  {32'h42563f2b, 32'h4276ee96} /* (31, 28, 7) {real, imag} */,
  {32'h426d91ae, 32'h426d1409} /* (31, 28, 6) {real, imag} */,
  {32'h41ca48be, 32'h41d28aff} /* (31, 28, 5) {real, imag} */,
  {32'hc1a0e22c, 32'h40ff53d7} /* (31, 28, 4) {real, imag} */,
  {32'hbfd7a58c, 32'hc04a9094} /* (31, 28, 3) {real, imag} */,
  {32'h41854dcc, 32'hc19612d2} /* (31, 28, 2) {real, imag} */,
  {32'h41026dee, 32'hc1b3bfe6} /* (31, 28, 1) {real, imag} */,
  {32'h3fd3a2ee, 32'hc187ab40} /* (31, 28, 0) {real, imag} */,
  {32'h400d33da, 32'hc0bd5acc} /* (31, 27, 31) {real, imag} */,
  {32'h3ea409e0, 32'hc1bdb412} /* (31, 27, 30) {real, imag} */,
  {32'hc1615429, 32'hc1a5fc8c} /* (31, 27, 29) {real, imag} */,
  {32'hc18d6fb5, 32'hc13cb47e} /* (31, 27, 28) {real, imag} */,
  {32'hc19493d1, 32'hc12bee06} /* (31, 27, 27) {real, imag} */,
  {32'hc18cf76c, 32'hc110de75} /* (31, 27, 26) {real, imag} */,
  {32'hc1b64839, 32'hc0ea21a8} /* (31, 27, 25) {real, imag} */,
  {32'hc23e2517, 32'hc1ca3f2a} /* (31, 27, 24) {real, imag} */,
  {32'hc24dba10, 32'hc24556a9} /* (31, 27, 23) {real, imag} */,
  {32'hc1a3d7fc, 32'hc2349a9e} /* (31, 27, 22) {real, imag} */,
  {32'hc0cfa437, 32'hc204fc8f} /* (31, 27, 21) {real, imag} */,
  {32'hbf1ec3b0, 32'h40e18dd0} /* (31, 27, 20) {real, imag} */,
  {32'hbf85a454, 32'h41444050} /* (31, 27, 19) {real, imag} */,
  {32'h40f82ed6, 32'h417fe174} /* (31, 27, 18) {real, imag} */,
  {32'h416dbf78, 32'h416001ce} /* (31, 27, 17) {real, imag} */,
  {32'h4182ef04, 32'h415f786d} /* (31, 27, 16) {real, imag} */,
  {32'h41aa8741, 32'h41df378e} /* (31, 27, 15) {real, imag} */,
  {32'h41fa6eee, 32'h41873b9d} /* (31, 27, 14) {real, imag} */,
  {32'h41f3de83, 32'h41b61ad8} /* (31, 27, 13) {real, imag} */,
  {32'h41a7e69b, 32'h4208a722} /* (31, 27, 12) {real, imag} */,
  {32'h406d21f8, 32'h422053a6} /* (31, 27, 11) {real, imag} */,
  {32'h410a32d2, 32'h4130f867} /* (31, 27, 10) {real, imag} */,
  {32'hc189ebfc, 32'h403f68f0} /* (31, 27, 9) {real, imag} */,
  {32'hc1f83047, 32'hc0da710e} /* (31, 27, 8) {real, imag} */,
  {32'hc17d8588, 32'hc11e5f5a} /* (31, 27, 7) {real, imag} */,
  {32'hc13b96c0, 32'h3fb34134} /* (31, 27, 6) {real, imag} */,
  {32'hc11b634a, 32'hc212d4fe} /* (31, 27, 5) {real, imag} */,
  {32'hc19c34ef, 32'hc2260dd3} /* (31, 27, 4) {real, imag} */,
  {32'hc0d0fa61, 32'hc1d0677a} /* (31, 27, 3) {real, imag} */,
  {32'hc1972495, 32'h3fe32eb0} /* (31, 27, 2) {real, imag} */,
  {32'hc0829490, 32'hc083e708} /* (31, 27, 1) {real, imag} */,
  {32'hc0b16873, 32'hc04c6af8} /* (31, 27, 0) {real, imag} */,
  {32'h40ea4502, 32'hbdd62660} /* (31, 26, 31) {real, imag} */,
  {32'hc0a1ada8, 32'hbfeea514} /* (31, 26, 30) {real, imag} */,
  {32'hc070c338, 32'h3f84d5d4} /* (31, 26, 29) {real, imag} */,
  {32'h3f17ac60, 32'h4044794d} /* (31, 26, 28) {real, imag} */,
  {32'hbf9e7198, 32'hbf65d360} /* (31, 26, 27) {real, imag} */,
  {32'hc03020c1, 32'h40b3844a} /* (31, 26, 26) {real, imag} */,
  {32'h41437266, 32'h408855d9} /* (31, 26, 25) {real, imag} */,
  {32'h41b67ae4, 32'hbf9519d0} /* (31, 26, 24) {real, imag} */,
  {32'hc072741e, 32'h41135c05} /* (31, 26, 23) {real, imag} */,
  {32'hbf78e278, 32'h40ebe304} /* (31, 26, 22) {real, imag} */,
  {32'h408d59d4, 32'h40aa5944} /* (31, 26, 21) {real, imag} */,
  {32'h41bfbdfa, 32'h40c73be6} /* (31, 26, 20) {real, imag} */,
  {32'h40e7dc2e, 32'hc138069f} /* (31, 26, 19) {real, imag} */,
  {32'h4016889c, 32'hc08e2be2} /* (31, 26, 18) {real, imag} */,
  {32'h41051f86, 32'h41390a53} /* (31, 26, 17) {real, imag} */,
  {32'hc11abb0c, 32'hc03b2b3e} /* (31, 26, 16) {real, imag} */,
  {32'hc19b061d, 32'h40a33bd2} /* (31, 26, 15) {real, imag} */,
  {32'h411a3b34, 32'h4174c23e} /* (31, 26, 14) {real, imag} */,
  {32'h40c257e4, 32'h41314dcd} /* (31, 26, 13) {real, imag} */,
  {32'h41178d80, 32'h3d2d9b00} /* (31, 26, 12) {real, imag} */,
  {32'h4164af7e, 32'hc182a3a1} /* (31, 26, 11) {real, imag} */,
  {32'h421f9a50, 32'hc07db4fa} /* (31, 26, 10) {real, imag} */,
  {32'h4200f6e6, 32'h40e1c4b6} /* (31, 26, 9) {real, imag} */,
  {32'h40858d85, 32'hbf3b42dc} /* (31, 26, 8) {real, imag} */,
  {32'h410b5d34, 32'h40edbcc5} /* (31, 26, 7) {real, imag} */,
  {32'h411b4a51, 32'h41ad1783} /* (31, 26, 6) {real, imag} */,
  {32'h413dd7b3, 32'h3ff32974} /* (31, 26, 5) {real, imag} */,
  {32'h40c64f5c, 32'hc11fbb1e} /* (31, 26, 4) {real, imag} */,
  {32'hc1078c80, 32'h4143b7a6} /* (31, 26, 3) {real, imag} */,
  {32'hc1baae5c, 32'hc085bb88} /* (31, 26, 2) {real, imag} */,
  {32'hc12059d2, 32'hc0e4fdfd} /* (31, 26, 1) {real, imag} */,
  {32'h405b8267, 32'h3e36b280} /* (31, 26, 0) {real, imag} */,
  {32'h3f3fe594, 32'h41096c32} /* (31, 25, 31) {real, imag} */,
  {32'h3fb65908, 32'h411002be} /* (31, 25, 30) {real, imag} */,
  {32'h411609c5, 32'h4039f47e} /* (31, 25, 29) {real, imag} */,
  {32'h40fc1e1c, 32'h4143b4e4} /* (31, 25, 28) {real, imag} */,
  {32'h413016d6, 32'h41bbb565} /* (31, 25, 27) {real, imag} */,
  {32'h41e55aa3, 32'h41855a49} /* (31, 25, 26) {real, imag} */,
  {32'h419c9f48, 32'h412a3ab6} /* (31, 25, 25) {real, imag} */,
  {32'h4183b1e4, 32'h41a65042} /* (31, 25, 24) {real, imag} */,
  {32'h41208bd0, 32'h42002c82} /* (31, 25, 23) {real, imag} */,
  {32'h414ee53d, 32'h41149d24} /* (31, 25, 22) {real, imag} */,
  {32'h4082eff7, 32'hc046d4f0} /* (31, 25, 21) {real, imag} */,
  {32'h404eeb92, 32'hc06b9910} /* (31, 25, 20) {real, imag} */,
  {32'h40ad7530, 32'hc09d1ec2} /* (31, 25, 19) {real, imag} */,
  {32'hc0c0a5b8, 32'hc099b670} /* (31, 25, 18) {real, imag} */,
  {32'hc1934b02, 32'hc0ac3365} /* (31, 25, 17) {real, imag} */,
  {32'hc1aac0bb, 32'hc0759cc7} /* (31, 25, 16) {real, imag} */,
  {32'hc1090eac, 32'hc1c5181d} /* (31, 25, 15) {real, imag} */,
  {32'hc11c266e, 32'hc11623c3} /* (31, 25, 14) {real, imag} */,
  {32'hc0f7ebbd, 32'h4128c5a6} /* (31, 25, 13) {real, imag} */,
  {32'h403165d4, 32'hc109ce48} /* (31, 25, 12) {real, imag} */,
  {32'hc01e6f2c, 32'hc1b46122} /* (31, 25, 11) {real, imag} */,
  {32'h411f9d06, 32'hc1582e26} /* (31, 25, 10) {real, imag} */,
  {32'h410faf94, 32'h3f2efc98} /* (31, 25, 9) {real, imag} */,
  {32'h411bf8aa, 32'hc15f90a7} /* (31, 25, 8) {real, imag} */,
  {32'h41c911c5, 32'h40cbebc9} /* (31, 25, 7) {real, imag} */,
  {32'h4178157f, 32'h41d80063} /* (31, 25, 6) {real, imag} */,
  {32'h413461d9, 32'h40c7bffe} /* (31, 25, 5) {real, imag} */,
  {32'h41c7177e, 32'hc0087344} /* (31, 25, 4) {real, imag} */,
  {32'h40952569, 32'h413043f4} /* (31, 25, 3) {real, imag} */,
  {32'h401a2142, 32'hc07a8d4e} /* (31, 25, 2) {real, imag} */,
  {32'h4145e2da, 32'hc18614ba} /* (31, 25, 1) {real, imag} */,
  {32'h4142661f, 32'hc0c68f0c} /* (31, 25, 0) {real, imag} */,
  {32'hc0b22622, 32'hc0fc9f30} /* (31, 24, 31) {real, imag} */,
  {32'hc0ff49de, 32'hc15fa984} /* (31, 24, 30) {real, imag} */,
  {32'hc0a33159, 32'hc17f8343} /* (31, 24, 29) {real, imag} */,
  {32'hc171a93a, 32'hc18396e7} /* (31, 24, 28) {real, imag} */,
  {32'hc2067bfa, 32'hc02bd71e} /* (31, 24, 27) {real, imag} */,
  {32'hc1fa6152, 32'hc0572f27} /* (31, 24, 26) {real, imag} */,
  {32'hc110eaee, 32'hc0f31cbe} /* (31, 24, 25) {real, imag} */,
  {32'hbf5a4cf8, 32'hc10b3837} /* (31, 24, 24) {real, imag} */,
  {32'hc0adf19e, 32'hc1a52f96} /* (31, 24, 23) {real, imag} */,
  {32'hbfcb84b8, 32'hc1a6cbd4} /* (31, 24, 22) {real, imag} */,
  {32'hc0af8572, 32'hc1366f46} /* (31, 24, 21) {real, imag} */,
  {32'h40f1f307, 32'h40bb4244} /* (31, 24, 20) {real, imag} */,
  {32'h406e9c02, 32'h41d9ecc0} /* (31, 24, 19) {real, imag} */,
  {32'h40e4af0e, 32'h4200ba96} /* (31, 24, 18) {real, imag} */,
  {32'h4148f087, 32'h41896ca4} /* (31, 24, 17) {real, imag} */,
  {32'h3f8fd7d4, 32'h41a86484} /* (31, 24, 16) {real, imag} */,
  {32'h3fb39ba4, 32'hc0bfe1a6} /* (31, 24, 15) {real, imag} */,
  {32'h415db8f4, 32'h40fb4024} /* (31, 24, 14) {real, imag} */,
  {32'h41cda8b6, 32'h41a063f0} /* (31, 24, 13) {real, imag} */,
  {32'h40e9a008, 32'h41e0ee97} /* (31, 24, 12) {real, imag} */,
  {32'hc060d1b8, 32'h4126f0ce} /* (31, 24, 11) {real, imag} */,
  {32'hbedac5cc, 32'hc156c0a5} /* (31, 24, 10) {real, imag} */,
  {32'hc0804604, 32'hc20b2ec8} /* (31, 24, 9) {real, imag} */,
  {32'hc16d96f2, 32'hc202dac0} /* (31, 24, 8) {real, imag} */,
  {32'hc1807a0c, 32'hc0ab5b68} /* (31, 24, 7) {real, imag} */,
  {32'h401ecf36, 32'hc0972674} /* (31, 24, 6) {real, imag} */,
  {32'h416c2462, 32'hc1bb3f4b} /* (31, 24, 5) {real, imag} */,
  {32'h411e0c91, 32'hc19f52c1} /* (31, 24, 4) {real, imag} */,
  {32'hc182f87e, 32'hc0cb3a04} /* (31, 24, 3) {real, imag} */,
  {32'hc1c4dc51, 32'hc0c12098} /* (31, 24, 2) {real, imag} */,
  {32'hc1b8ea4b, 32'hc0a9cdac} /* (31, 24, 1) {real, imag} */,
  {32'hbfa5aeda, 32'hbfbb277a} /* (31, 24, 0) {real, imag} */,
  {32'h3fd0a38e, 32'h409b34a7} /* (31, 23, 31) {real, imag} */,
  {32'hc00d3efe, 32'h3fd998e4} /* (31, 23, 30) {real, imag} */,
  {32'hc1767e7d, 32'h407a8ea6} /* (31, 23, 29) {real, imag} */,
  {32'hc121b423, 32'h4092de3b} /* (31, 23, 28) {real, imag} */,
  {32'hc12529ea, 32'hbfe7d6f8} /* (31, 23, 27) {real, imag} */,
  {32'hc0e62e30, 32'hc10a4139} /* (31, 23, 26) {real, imag} */,
  {32'hc0e18df5, 32'hc1b2265d} /* (31, 23, 25) {real, imag} */,
  {32'hbf94989c, 32'hc10388b5} /* (31, 23, 24) {real, imag} */,
  {32'hc0da64ce, 32'hc0697ac0} /* (31, 23, 23) {real, imag} */,
  {32'hc172da21, 32'h41306ae4} /* (31, 23, 22) {real, imag} */,
  {32'hc1063fb6, 32'h4112b70e} /* (31, 23, 21) {real, imag} */,
  {32'hc126ab4a, 32'h4025df88} /* (31, 23, 20) {real, imag} */,
  {32'hc13cb772, 32'hc03c5008} /* (31, 23, 19) {real, imag} */,
  {32'hc18c2780, 32'hc07f3128} /* (31, 23, 18) {real, imag} */,
  {32'hc1a1df48, 32'h40364fc6} /* (31, 23, 17) {real, imag} */,
  {32'hc11335d7, 32'h40d9b07e} /* (31, 23, 16) {real, imag} */,
  {32'hc0836766, 32'h40f6440b} /* (31, 23, 15) {real, imag} */,
  {32'hc052d51a, 32'h3fa657a2} /* (31, 23, 14) {real, imag} */,
  {32'hc16273cc, 32'hc11e0320} /* (31, 23, 13) {real, imag} */,
  {32'hc1d5b3d2, 32'hc1238b68} /* (31, 23, 12) {real, imag} */,
  {32'hc18dd168, 32'hc15bd119} /* (31, 23, 11) {real, imag} */,
  {32'h40a07c16, 32'hc0ca1a94} /* (31, 23, 10) {real, imag} */,
  {32'hbf80ac00, 32'h3fbe046c} /* (31, 23, 9) {real, imag} */,
  {32'h4115dcba, 32'hc04d6694} /* (31, 23, 8) {real, imag} */,
  {32'hc0decd58, 32'hc01db6e2} /* (31, 23, 7) {real, imag} */,
  {32'h40d946b3, 32'hc147582e} /* (31, 23, 6) {real, imag} */,
  {32'h40eeddc0, 32'hc1790867} /* (31, 23, 5) {real, imag} */,
  {32'h4165a0c6, 32'hbfe85528} /* (31, 23, 4) {real, imag} */,
  {32'h4076cd7c, 32'h41113cf8} /* (31, 23, 3) {real, imag} */,
  {32'hbec81870, 32'hc10ec1a8} /* (31, 23, 2) {real, imag} */,
  {32'hc13b5add, 32'hc0e5775b} /* (31, 23, 1) {real, imag} */,
  {32'hc0d1ae2a, 32'hbf5b73c0} /* (31, 23, 0) {real, imag} */,
  {32'h4056c3ea, 32'h3f9ec7ca} /* (31, 22, 31) {real, imag} */,
  {32'hc05c7946, 32'hc1210e09} /* (31, 22, 30) {real, imag} */,
  {32'hc18f5d20, 32'hc091e5d1} /* (31, 22, 29) {real, imag} */,
  {32'hc073f645, 32'h40fd0be2} /* (31, 22, 28) {real, imag} */,
  {32'h403f12a6, 32'h41779b7a} /* (31, 22, 27) {real, imag} */,
  {32'hc09b3310, 32'h412997d8} /* (31, 22, 26) {real, imag} */,
  {32'h41087476, 32'h3fc03f94} /* (31, 22, 25) {real, imag} */,
  {32'h41160532, 32'hc0978b7a} /* (31, 22, 24) {real, imag} */,
  {32'h411550a4, 32'hbf24abe8} /* (31, 22, 23) {real, imag} */,
  {32'h41a146e9, 32'hc1023690} /* (31, 22, 22) {real, imag} */,
  {32'h40d749bb, 32'h4118175c} /* (31, 22, 21) {real, imag} */,
  {32'hc009c76e, 32'h40b87fbd} /* (31, 22, 20) {real, imag} */,
  {32'hc1033bcd, 32'hc1624390} /* (31, 22, 19) {real, imag} */,
  {32'hc19d35bc, 32'hc14d0b7b} /* (31, 22, 18) {real, imag} */,
  {32'hc1395b3f, 32'hbf9af798} /* (31, 22, 17) {real, imag} */,
  {32'hc0c52df8, 32'hc0ec4377} /* (31, 22, 16) {real, imag} */,
  {32'hc0c7bdc5, 32'h3ea2c230} /* (31, 22, 15) {real, imag} */,
  {32'hc08685d5, 32'h400b99d0} /* (31, 22, 14) {real, imag} */,
  {32'hc0763668, 32'hc019e320} /* (31, 22, 13) {real, imag} */,
  {32'hc1101f3e, 32'hc10d26cb} /* (31, 22, 12) {real, imag} */,
  {32'hc1166cce, 32'hc0d1bf54} /* (31, 22, 11) {real, imag} */,
  {32'h40a62f76, 32'hc0dad899} /* (31, 22, 10) {real, imag} */,
  {32'h413caaf6, 32'hbdb7ae80} /* (31, 22, 9) {real, imag} */,
  {32'h412cd2d0, 32'h4169974c} /* (31, 22, 8) {real, imag} */,
  {32'h40ee5378, 32'h4139d0a8} /* (31, 22, 7) {real, imag} */,
  {32'h414972c5, 32'h4144af14} /* (31, 22, 6) {real, imag} */,
  {32'h411de349, 32'h3ecc7b30} /* (31, 22, 5) {real, imag} */,
  {32'h40a43d93, 32'h402cfbca} /* (31, 22, 4) {real, imag} */,
  {32'hbfceef44, 32'h3e29fa80} /* (31, 22, 3) {real, imag} */,
  {32'h3f80b732, 32'h3f11a538} /* (31, 22, 2) {real, imag} */,
  {32'h40f15337, 32'h40f709b9} /* (31, 22, 1) {real, imag} */,
  {32'h412315d6, 32'h413078b8} /* (31, 22, 0) {real, imag} */,
  {32'hc039231f, 32'hc10c3b6e} /* (31, 21, 31) {real, imag} */,
  {32'hbfcc77aa, 32'hc0c4e8fa} /* (31, 21, 30) {real, imag} */,
  {32'hbea3dce0, 32'hc158b014} /* (31, 21, 29) {real, imag} */,
  {32'hc01ec996, 32'hc0fecb96} /* (31, 21, 28) {real, imag} */,
  {32'hc161514c, 32'hbf6886b0} /* (31, 21, 27) {real, imag} */,
  {32'hc12bc0aa, 32'hc0426fe6} /* (31, 21, 26) {real, imag} */,
  {32'hc1001510, 32'hbfdbb500} /* (31, 21, 25) {real, imag} */,
  {32'hc0cc4667, 32'hbf8e4680} /* (31, 21, 24) {real, imag} */,
  {32'hc112ad86, 32'hc11dcd33} /* (31, 21, 23) {real, imag} */,
  {32'hc16cc1c3, 32'hc1167f61} /* (31, 21, 22) {real, imag} */,
  {32'hc1623ea2, 32'hc041f86e} /* (31, 21, 21) {real, imag} */,
  {32'hc0ebdb48, 32'h3e11c450} /* (31, 21, 20) {real, imag} */,
  {32'hbf3581c8, 32'h40751108} /* (31, 21, 19) {real, imag} */,
  {32'h4067f6d3, 32'h41236170} /* (31, 21, 18) {real, imag} */,
  {32'h3fd1f15e, 32'h414c0ce2} /* (31, 21, 17) {real, imag} */,
  {32'h409ae1ea, 32'h4141de3e} /* (31, 21, 16) {real, imag} */,
  {32'h40b11f30, 32'h4105d136} /* (31, 21, 15) {real, imag} */,
  {32'h410a58b6, 32'hbffcd34c} /* (31, 21, 14) {real, imag} */,
  {32'h40cb93d5, 32'h4027d376} /* (31, 21, 13) {real, imag} */,
  {32'h4148469a, 32'h410d1499} /* (31, 21, 12) {real, imag} */,
  {32'h41712180, 32'h4119b483} /* (31, 21, 11) {real, imag} */,
  {32'hbf62e3b8, 32'hc059f82f} /* (31, 21, 10) {real, imag} */,
  {32'hc1105981, 32'hbf0a9de8} /* (31, 21, 9) {real, imag} */,
  {32'hc111c9f6, 32'h40a3c4c0} /* (31, 21, 8) {real, imag} */,
  {32'hc183afe6, 32'h40a13e5f} /* (31, 21, 7) {real, imag} */,
  {32'hc0f9414b, 32'h40801bc1} /* (31, 21, 6) {real, imag} */,
  {32'hbfa97dfe, 32'h3fb9b108} /* (31, 21, 5) {real, imag} */,
  {32'hc15278a7, 32'hc034ec89} /* (31, 21, 4) {real, imag} */,
  {32'hc16b02c8, 32'hc0c2a4e7} /* (31, 21, 3) {real, imag} */,
  {32'hbf6398f8, 32'hbfd878d4} /* (31, 21, 2) {real, imag} */,
  {32'h3e809380, 32'hc03d21a8} /* (31, 21, 1) {real, imag} */,
  {32'hc08fde24, 32'hc0c616c4} /* (31, 21, 0) {real, imag} */,
  {32'h3f32d496, 32'h40722b52} /* (31, 20, 31) {real, imag} */,
  {32'h40f444fc, 32'hbf49be80} /* (31, 20, 30) {real, imag} */,
  {32'h40dfeb9e, 32'h3f2c6748} /* (31, 20, 29) {real, imag} */,
  {32'hc089f33a, 32'hbf22c230} /* (31, 20, 28) {real, imag} */,
  {32'h404f4759, 32'h3fee58cc} /* (31, 20, 27) {real, imag} */,
  {32'h413f9b22, 32'h3fe0b170} /* (31, 20, 26) {real, imag} */,
  {32'h3f372450, 32'hc0a9a3ad} /* (31, 20, 25) {real, imag} */,
  {32'hc1752f74, 32'hc0fb1bc3} /* (31, 20, 24) {real, imag} */,
  {32'hc0968597, 32'hc101e33c} /* (31, 20, 23) {real, imag} */,
  {32'h412d8815, 32'hc1276808} /* (31, 20, 22) {real, imag} */,
  {32'h410f0746, 32'hc0a841ee} /* (31, 20, 21) {real, imag} */,
  {32'h40982d14, 32'hc08e5ce2} /* (31, 20, 20) {real, imag} */,
  {32'h40d4e354, 32'hc0dfedf6} /* (31, 20, 19) {real, imag} */,
  {32'h410e919e, 32'hc09b6be6} /* (31, 20, 18) {real, imag} */,
  {32'h3fa44158, 32'hc0f4fcc8} /* (31, 20, 17) {real, imag} */,
  {32'hbf692f00, 32'hc0832d53} /* (31, 20, 16) {real, imag} */,
  {32'h3f0bd980, 32'hc0b56eba} /* (31, 20, 15) {real, imag} */,
  {32'hbf904c8c, 32'hbcd3c180} /* (31, 20, 14) {real, imag} */,
  {32'hc097f02b, 32'h401b3bd4} /* (31, 20, 13) {real, imag} */,
  {32'hc0013208, 32'h3f233cc0} /* (31, 20, 12) {real, imag} */,
  {32'h3d42de80, 32'hc05b8b59} /* (31, 20, 11) {real, imag} */,
  {32'hc04cb722, 32'h408649ca} /* (31, 20, 10) {real, imag} */,
  {32'hbf4daa20, 32'h40a2010a} /* (31, 20, 9) {real, imag} */,
  {32'h40b69cfd, 32'h3f5d2746} /* (31, 20, 8) {real, imag} */,
  {32'h4138322d, 32'h40b8bc98} /* (31, 20, 7) {real, imag} */,
  {32'hc0238e60, 32'h402b07c0} /* (31, 20, 6) {real, imag} */,
  {32'hc101fe5f, 32'hbea537c0} /* (31, 20, 5) {real, imag} */,
  {32'h3f25d21c, 32'h4120e318} /* (31, 20, 4) {real, imag} */,
  {32'h3e1eb630, 32'h411d9a22} /* (31, 20, 3) {real, imag} */,
  {32'h3f7c35b0, 32'hbf238690} /* (31, 20, 2) {real, imag} */,
  {32'h40a7ecc2, 32'h4097c3e1} /* (31, 20, 1) {real, imag} */,
  {32'hbf98f426, 32'h40aa6b18} /* (31, 20, 0) {real, imag} */,
  {32'h40b9a2a0, 32'h3f9e3d3c} /* (31, 19, 31) {real, imag} */,
  {32'h4102e7ae, 32'h3f8e3b6c} /* (31, 19, 30) {real, imag} */,
  {32'h3ec5c318, 32'h40eb97c1} /* (31, 19, 29) {real, imag} */,
  {32'hbffdffa2, 32'h40b39490} /* (31, 19, 28) {real, imag} */,
  {32'h4002fa44, 32'h4095d2e4} /* (31, 19, 27) {real, imag} */,
  {32'hc00a6d8a, 32'h40b15217} /* (31, 19, 26) {real, imag} */,
  {32'hc049f3da, 32'h3ec64380} /* (31, 19, 25) {real, imag} */,
  {32'hc0f2479a, 32'hbf46a8a4} /* (31, 19, 24) {real, imag} */,
  {32'hbe258640, 32'h40bf3034} /* (31, 19, 23) {real, imag} */,
  {32'h4103e320, 32'h41263b70} /* (31, 19, 22) {real, imag} */,
  {32'h401b1adc, 32'h3ff23648} /* (31, 19, 21) {real, imag} */,
  {32'h3f98b424, 32'hbfe3e3b4} /* (31, 19, 20) {real, imag} */,
  {32'h3f06b330, 32'hbfb4c874} /* (31, 19, 19) {real, imag} */,
  {32'h40780514, 32'h4058fac0} /* (31, 19, 18) {real, imag} */,
  {32'h3f639804, 32'h4179adcb} /* (31, 19, 17) {real, imag} */,
  {32'h40a50ff2, 32'h4089bc5c} /* (31, 19, 16) {real, imag} */,
  {32'h40cb50b8, 32'hc0a5b988} /* (31, 19, 15) {real, imag} */,
  {32'h40119581, 32'hc17fc5b3} /* (31, 19, 14) {real, imag} */,
  {32'hbfd58752, 32'hc115b304} /* (31, 19, 13) {real, imag} */,
  {32'h4044ec3e, 32'hc1016ed2} /* (31, 19, 12) {real, imag} */,
  {32'h40117d5b, 32'hc143f4f0} /* (31, 19, 11) {real, imag} */,
  {32'hc026e674, 32'hc14a0da8} /* (31, 19, 10) {real, imag} */,
  {32'h40324b81, 32'hc1395246} /* (31, 19, 9) {real, imag} */,
  {32'h408e606e, 32'hc1800439} /* (31, 19, 8) {real, imag} */,
  {32'h3ffe06cc, 32'hc11e4864} /* (31, 19, 7) {real, imag} */,
  {32'hc076935c, 32'hc0a66fe9} /* (31, 19, 6) {real, imag} */,
  {32'hc09af39e, 32'h3ed5f520} /* (31, 19, 5) {real, imag} */,
  {32'hc09d44de, 32'hbfe65ad4} /* (31, 19, 4) {real, imag} */,
  {32'h3f622a90, 32'hbfebf586} /* (31, 19, 3) {real, imag} */,
  {32'h40efc147, 32'h41438216} /* (31, 19, 2) {real, imag} */,
  {32'h409f625c, 32'h41095548} /* (31, 19, 1) {real, imag} */,
  {32'h3f8eaa0a, 32'h3f22c2dc} /* (31, 19, 0) {real, imag} */,
  {32'hc01ff260, 32'h40664c46} /* (31, 18, 31) {real, imag} */,
  {32'hc0c0f420, 32'h40e697a6} /* (31, 18, 30) {real, imag} */,
  {32'hc1216a70, 32'h4103c0f1} /* (31, 18, 29) {real, imag} */,
  {32'hc113b7dc, 32'h402b008e} /* (31, 18, 28) {real, imag} */,
  {32'hc0a95068, 32'h40ca56b5} /* (31, 18, 27) {real, imag} */,
  {32'h4089f825, 32'h40759c59} /* (31, 18, 26) {real, imag} */,
  {32'hc0512a5c, 32'h40a8e7f0} /* (31, 18, 25) {real, imag} */,
  {32'hc1103f10, 32'h40b3925c} /* (31, 18, 24) {real, imag} */,
  {32'hc112b7ee, 32'hbf81bf60} /* (31, 18, 23) {real, imag} */,
  {32'hc0e151a4, 32'hc0d29d88} /* (31, 18, 22) {real, imag} */,
  {32'h40ac53b8, 32'hc03e843c} /* (31, 18, 21) {real, imag} */,
  {32'h411a2880, 32'h404e6546} /* (31, 18, 20) {real, imag} */,
  {32'h40db1312, 32'h3f71128a} /* (31, 18, 19) {real, imag} */,
  {32'h402112c0, 32'h3ead14e0} /* (31, 18, 18) {real, imag} */,
  {32'h3fd2308c, 32'h4001aef4} /* (31, 18, 17) {real, imag} */,
  {32'h4099ab63, 32'h3ffb6bf4} /* (31, 18, 16) {real, imag} */,
  {32'h40a1541a, 32'h3ec2ec20} /* (31, 18, 15) {real, imag} */,
  {32'h40a3ffd9, 32'hbe5b59e0} /* (31, 18, 14) {real, imag} */,
  {32'h4008f688, 32'h40033cd4} /* (31, 18, 13) {real, imag} */,
  {32'h407734bd, 32'hbef03470} /* (31, 18, 12) {real, imag} */,
  {32'h408dd264, 32'h4008b902} /* (31, 18, 11) {real, imag} */,
  {32'hbf6681d0, 32'h4072ec96} /* (31, 18, 10) {real, imag} */,
  {32'hbfce3018, 32'hbe5f21a0} /* (31, 18, 9) {real, imag} */,
  {32'hbe4b9680, 32'hc03e9fec} /* (31, 18, 8) {real, imag} */,
  {32'hbf9ffbd0, 32'hc0aca254} /* (31, 18, 7) {real, imag} */,
  {32'hc08239ca, 32'h3efb3420} /* (31, 18, 6) {real, imag} */,
  {32'hc0a1e450, 32'h409fc49d} /* (31, 18, 5) {real, imag} */,
  {32'hc12e212e, 32'h4113898c} /* (31, 18, 4) {real, imag} */,
  {32'hc13dbc4b, 32'h41086493} /* (31, 18, 3) {real, imag} */,
  {32'hc0d12ea4, 32'h40e0a60e} /* (31, 18, 2) {real, imag} */,
  {32'hc12d3439, 32'h401b871e} /* (31, 18, 1) {real, imag} */,
  {32'hc0e69828, 32'h3e8e0f60} /* (31, 18, 0) {real, imag} */,
  {32'h3f4b651c, 32'h3f91e4b6} /* (31, 17, 31) {real, imag} */,
  {32'h40fbafc8, 32'h403cc590} /* (31, 17, 30) {real, imag} */,
  {32'h4031e7df, 32'hbfc1944c} /* (31, 17, 29) {real, imag} */,
  {32'hc05ad182, 32'hbf966104} /* (31, 17, 28) {real, imag} */,
  {32'h4061a8e6, 32'hbf1b8810} /* (31, 17, 27) {real, imag} */,
  {32'h40d02b26, 32'hbf559830} /* (31, 17, 26) {real, imag} */,
  {32'h4025238e, 32'h40cb870e} /* (31, 17, 25) {real, imag} */,
  {32'h40ded49f, 32'h409c19b6} /* (31, 17, 24) {real, imag} */,
  {32'h40b58f9e, 32'h3ee36c10} /* (31, 17, 23) {real, imag} */,
  {32'h3b9c2200, 32'h40dc6332} /* (31, 17, 22) {real, imag} */,
  {32'hbf95727c, 32'h410a0e1e} /* (31, 17, 21) {real, imag} */,
  {32'hc0454326, 32'h40939170} /* (31, 17, 20) {real, imag} */,
  {32'hc0d716e9, 32'hbf187f78} /* (31, 17, 19) {real, imag} */,
  {32'hc04ee9f0, 32'hbfc72814} /* (31, 17, 18) {real, imag} */,
  {32'hc008985c, 32'hc0540c7c} /* (31, 17, 17) {real, imag} */,
  {32'hbfd3e2cc, 32'hbfc0bff0} /* (31, 17, 16) {real, imag} */,
  {32'hc00e8495, 32'hbf0637a0} /* (31, 17, 15) {real, imag} */,
  {32'h3f8f440e, 32'hc058150e} /* (31, 17, 14) {real, imag} */,
  {32'hc03c4c64, 32'hbfa38f00} /* (31, 17, 13) {real, imag} */,
  {32'hc004214c, 32'h407bf25f} /* (31, 17, 12) {real, imag} */,
  {32'h3f32175c, 32'hbfe765f8} /* (31, 17, 11) {real, imag} */,
  {32'hbdd9f340, 32'hbfdab04c} /* (31, 17, 10) {real, imag} */,
  {32'hbef27360, 32'hbeed5298} /* (31, 17, 9) {real, imag} */,
  {32'hbffd65c0, 32'h40715db6} /* (31, 17, 8) {real, imag} */,
  {32'hbeb40d58, 32'h404e8454} /* (31, 17, 7) {real, imag} */,
  {32'h41051e53, 32'hc047086d} /* (31, 17, 6) {real, imag} */,
  {32'h409a48de, 32'hc09074fa} /* (31, 17, 5) {real, imag} */,
  {32'h4040d572, 32'hc0736f57} /* (31, 17, 4) {real, imag} */,
  {32'hc0c590ae, 32'hbfe59e28} /* (31, 17, 3) {real, imag} */,
  {32'hc0c94520, 32'h408bba32} /* (31, 17, 2) {real, imag} */,
  {32'h40476505, 32'h40ea0db5} /* (31, 17, 1) {real, imag} */,
  {32'h3fd6c1f0, 32'h401a7168} /* (31, 17, 0) {real, imag} */,
  {32'hbf9ec0f8, 32'hc0b404b0} /* (31, 16, 31) {real, imag} */,
  {32'hbe7d4c80, 32'hc11c2cd8} /* (31, 16, 30) {real, imag} */,
  {32'h3ea163b0, 32'hc0c0c1f0} /* (31, 16, 29) {real, imag} */,
  {32'hbf10d568, 32'h3fb71860} /* (31, 16, 28) {real, imag} */,
  {32'hc07405bc, 32'h4086eb90} /* (31, 16, 27) {real, imag} */,
  {32'hc0876bea, 32'h3fcca700} /* (31, 16, 26) {real, imag} */,
  {32'hbf5756b8, 32'hbf2db080} /* (31, 16, 25) {real, imag} */,
  {32'h3f2673d4, 32'h40ad1f30} /* (31, 16, 24) {real, imag} */,
  {32'hbffd10c0, 32'h4085cf60} /* (31, 16, 23) {real, imag} */,
  {32'h4076f940, 32'h40b9d578} /* (31, 16, 22) {real, imag} */,
  {32'h40bb324b, 32'hc02ff3d0} /* (31, 16, 21) {real, imag} */,
  {32'h3da4c240, 32'hbce16c00} /* (31, 16, 20) {real, imag} */,
  {32'hc044fdfa, 32'h40172cae} /* (31, 16, 19) {real, imag} */,
  {32'hbf2ae078, 32'hbf71c268} /* (31, 16, 18) {real, imag} */,
  {32'hbf3ab6e8, 32'h404b06dc} /* (31, 16, 17) {real, imag} */,
  {32'hbd83b280, 32'hc0843e8c} /* (31, 16, 16) {real, imag} */,
  {32'hc0b313ba, 32'hc04f3be0} /* (31, 16, 15) {real, imag} */,
  {32'hc0b35530, 32'h402d97e0} /* (31, 16, 14) {real, imag} */,
  {32'hc0742b44, 32'h40a273b0} /* (31, 16, 13) {real, imag} */,
  {32'hbeb6a510, 32'hbf20a240} /* (31, 16, 12) {real, imag} */,
  {32'hc0a5a546, 32'h3f123780} /* (31, 16, 11) {real, imag} */,
  {32'hc08d63c6, 32'hbff5997c} /* (31, 16, 10) {real, imag} */,
  {32'hbe8c3280, 32'hbfadb610} /* (31, 16, 9) {real, imag} */,
  {32'hbf199120, 32'hbf363728} /* (31, 16, 8) {real, imag} */,
  {32'hbf0f55a0, 32'h3ffb4f80} /* (31, 16, 7) {real, imag} */,
  {32'h4031427c, 32'h4080fc25} /* (31, 16, 6) {real, imag} */,
  {32'h408fb1da, 32'h3ea6bb80} /* (31, 16, 5) {real, imag} */,
  {32'h403b5e73, 32'h3f019700} /* (31, 16, 4) {real, imag} */,
  {32'h409767ef, 32'h408658a8} /* (31, 16, 3) {real, imag} */,
  {32'h402e700c, 32'h40ab4ae0} /* (31, 16, 2) {real, imag} */,
  {32'h40b34e31, 32'hc0425690} /* (31, 16, 1) {real, imag} */,
  {32'h4016ed69, 32'hbff46260} /* (31, 16, 0) {real, imag} */,
  {32'hc05da3e3, 32'h408d8ed2} /* (31, 15, 31) {real, imag} */,
  {32'hc0d35c78, 32'h400fb4f0} /* (31, 15, 30) {real, imag} */,
  {32'hbf58f234, 32'hc048ebda} /* (31, 15, 29) {real, imag} */,
  {32'hbfa18c64, 32'hc0a92bbf} /* (31, 15, 28) {real, imag} */,
  {32'h3fbe4940, 32'hbe1913c0} /* (31, 15, 27) {real, imag} */,
  {32'h3c81be00, 32'h3f94f518} /* (31, 15, 26) {real, imag} */,
  {32'hc0295fc2, 32'hbd06f740} /* (31, 15, 25) {real, imag} */,
  {32'hbfb748ec, 32'hc0292c6d} /* (31, 15, 24) {real, imag} */,
  {32'hc050fd88, 32'hc0876ae1} /* (31, 15, 23) {real, imag} */,
  {32'hbf09bdf4, 32'hc06c7764} /* (31, 15, 22) {real, imag} */,
  {32'h3fd0295c, 32'hc0746298} /* (31, 15, 21) {real, imag} */,
  {32'h407b2f0a, 32'hbff2d940} /* (31, 15, 20) {real, imag} */,
  {32'hc0322bc2, 32'h409544e7} /* (31, 15, 19) {real, imag} */,
  {32'hc069d040, 32'h3faef194} /* (31, 15, 18) {real, imag} */,
  {32'h40c93f1a, 32'hbfe3cfc8} /* (31, 15, 17) {real, imag} */,
  {32'h4014557a, 32'h40720cd8} /* (31, 15, 16) {real, imag} */,
  {32'hc04ca58b, 32'h40384428} /* (31, 15, 15) {real, imag} */,
  {32'hc07697a7, 32'hc0952ed9} /* (31, 15, 14) {real, imag} */,
  {32'hbeb8ada0, 32'hc0922460} /* (31, 15, 13) {real, imag} */,
  {32'hbf84e0c8, 32'hbf908cbe} /* (31, 15, 12) {real, imag} */,
  {32'hc018eacf, 32'h41028bdf} /* (31, 15, 11) {real, imag} */,
  {32'h3fdc096c, 32'h4116554a} /* (31, 15, 10) {real, imag} */,
  {32'hbed93360, 32'h3fcfcfa6} /* (31, 15, 9) {real, imag} */,
  {32'hc1176624, 32'hc0458946} /* (31, 15, 8) {real, imag} */,
  {32'hc0f1bd0e, 32'hbe678540} /* (31, 15, 7) {real, imag} */,
  {32'hc008da54, 32'h3e01cad0} /* (31, 15, 6) {real, imag} */,
  {32'hc0a1c3c6, 32'hbf38b830} /* (31, 15, 5) {real, imag} */,
  {32'hc091b973, 32'hbf3cf624} /* (31, 15, 4) {real, imag} */,
  {32'hc0ae4a76, 32'hbdb0dd80} /* (31, 15, 3) {real, imag} */,
  {32'hc0afda70, 32'hbe560240} /* (31, 15, 2) {real, imag} */,
  {32'hc07667d5, 32'hc0ae9c35} /* (31, 15, 1) {real, imag} */,
  {32'hc021ece4, 32'hc03c1e28} /* (31, 15, 0) {real, imag} */,
  {32'h40c508e8, 32'h3f108be8} /* (31, 14, 31) {real, imag} */,
  {32'h414cdd38, 32'hc07f286c} /* (31, 14, 30) {real, imag} */,
  {32'h415b0e56, 32'hc0129644} /* (31, 14, 29) {real, imag} */,
  {32'h411b9a8c, 32'hbf999a1c} /* (31, 14, 28) {real, imag} */,
  {32'h40c5f1d4, 32'hbeaaa150} /* (31, 14, 27) {real, imag} */,
  {32'h3f808fec, 32'hbf9479f2} /* (31, 14, 26) {real, imag} */,
  {32'h403daf28, 32'hc0c13c30} /* (31, 14, 25) {real, imag} */,
  {32'h40b2d35b, 32'hc0aac92c} /* (31, 14, 24) {real, imag} */,
  {32'h3fa909c0, 32'h3eafd480} /* (31, 14, 23) {real, imag} */,
  {32'h408f6e06, 32'h400a8810} /* (31, 14, 22) {real, imag} */,
  {32'h411cb8ca, 32'hc0ae61d2} /* (31, 14, 21) {real, imag} */,
  {32'h40863688, 32'hc0aefcf3} /* (31, 14, 20) {real, imag} */,
  {32'hc09ea9a6, 32'hbf66b60a} /* (31, 14, 19) {real, imag} */,
  {32'hc0423070, 32'hbef1b2e0} /* (31, 14, 18) {real, imag} */,
  {32'hc0899295, 32'hbe8b83a0} /* (31, 14, 17) {real, imag} */,
  {32'hc0d776b5, 32'h3fed058c} /* (31, 14, 16) {real, imag} */,
  {32'hc0b006b6, 32'h40f1447e} /* (31, 14, 15) {real, imag} */,
  {32'hc0adb785, 32'hbfb6b584} /* (31, 14, 14) {real, imag} */,
  {32'hc03b7f18, 32'h3ff49d58} /* (31, 14, 13) {real, imag} */,
  {32'hbf151b4c, 32'h409034a7} /* (31, 14, 12) {real, imag} */,
  {32'hc12ea01c, 32'hbedefb10} /* (31, 14, 11) {real, imag} */,
  {32'h3e96a460, 32'hc10fb21e} /* (31, 14, 10) {real, imag} */,
  {32'h40461c34, 32'hc0aa5013} /* (31, 14, 9) {real, imag} */,
  {32'h40284508, 32'hbfb3c5a8} /* (31, 14, 8) {real, imag} */,
  {32'h3e7ccf80, 32'hc02478f8} /* (31, 14, 7) {real, imag} */,
  {32'hbfd98ba8, 32'hc065ca04} /* (31, 14, 6) {real, imag} */,
  {32'h40805120, 32'h40a9cec3} /* (31, 14, 5) {real, imag} */,
  {32'h40df3fa4, 32'h40c86379} /* (31, 14, 4) {real, imag} */,
  {32'h40a13092, 32'hbe82c560} /* (31, 14, 3) {real, imag} */,
  {32'h40025158, 32'hc04170dc} /* (31, 14, 2) {real, imag} */,
  {32'h40404364, 32'hbfd6ec3c} /* (31, 14, 1) {real, imag} */,
  {32'h3ff98236, 32'hbf50f6b0} /* (31, 14, 0) {real, imag} */,
  {32'hc00dbb69, 32'h40b5f6bb} /* (31, 13, 31) {real, imag} */,
  {32'hc0aeb5bb, 32'h3fd067fc} /* (31, 13, 30) {real, imag} */,
  {32'h408870e6, 32'hc0b4c57f} /* (31, 13, 29) {real, imag} */,
  {32'h40893b34, 32'hc1149622} /* (31, 13, 28) {real, imag} */,
  {32'hbf7c5d8a, 32'hc02d2da4} /* (31, 13, 27) {real, imag} */,
  {32'h4027f5fc, 32'hc0b74f71} /* (31, 13, 26) {real, imag} */,
  {32'h4068c326, 32'hc0da0238} /* (31, 13, 25) {real, imag} */,
  {32'h40b09e7c, 32'hbf35988c} /* (31, 13, 24) {real, imag} */,
  {32'h40ad07ba, 32'hc08bab04} /* (31, 13, 23) {real, imag} */,
  {32'h407f17d8, 32'hc07f7706} /* (31, 13, 22) {real, imag} */,
  {32'h4075c740, 32'hc0ee87ea} /* (31, 13, 21) {real, imag} */,
  {32'h3f018ec8, 32'hc075098e} /* (31, 13, 20) {real, imag} */,
  {32'hbeaf9320, 32'h3fdbdf14} /* (31, 13, 19) {real, imag} */,
  {32'hc02d617c, 32'h3f19cbd0} /* (31, 13, 18) {real, imag} */,
  {32'hc050a33f, 32'hc0865942} /* (31, 13, 17) {real, imag} */,
  {32'hc051164d, 32'hc06e0030} /* (31, 13, 16) {real, imag} */,
  {32'hc039cd10, 32'h40acc34c} /* (31, 13, 15) {real, imag} */,
  {32'hc0a6e0a8, 32'h40e79f42} /* (31, 13, 14) {real, imag} */,
  {32'hc0a641dc, 32'h40895d01} /* (31, 13, 13) {real, imag} */,
  {32'hc0893444, 32'h40f03804} /* (31, 13, 12) {real, imag} */,
  {32'h403caba1, 32'hbf3f8ed0} /* (31, 13, 11) {real, imag} */,
  {32'hbf02f290, 32'hc0ecde01} /* (31, 13, 10) {real, imag} */,
  {32'hc1004f64, 32'h407d6676} /* (31, 13, 9) {real, imag} */,
  {32'hc17b1ef1, 32'h404be2fa} /* (31, 13, 8) {real, imag} */,
  {32'hc181d3f3, 32'hc080ac8d} /* (31, 13, 7) {real, imag} */,
  {32'hbfc13eb8, 32'h3fbdcafc} /* (31, 13, 6) {real, imag} */,
  {32'h409df282, 32'h41385c3b} /* (31, 13, 5) {real, imag} */,
  {32'h4012ad51, 32'h40e9f31f} /* (31, 13, 4) {real, imag} */,
  {32'hc1028c49, 32'h406d8cd5} /* (31, 13, 3) {real, imag} */,
  {32'hc0ab60d5, 32'hbfc7e424} /* (31, 13, 2) {real, imag} */,
  {32'hbebe6408, 32'hbf8f9f3a} /* (31, 13, 1) {real, imag} */,
  {32'hbfb492d2, 32'hbee7cb48} /* (31, 13, 0) {real, imag} */,
  {32'h3fc9a40b, 32'h40358e9a} /* (31, 12, 31) {real, imag} */,
  {32'h3faa41c0, 32'hc0183cb8} /* (31, 12, 30) {real, imag} */,
  {32'hc0a22656, 32'hc10e123e} /* (31, 12, 29) {real, imag} */,
  {32'hc0c947c0, 32'hbfd115e8} /* (31, 12, 28) {real, imag} */,
  {32'h3fe09552, 32'h3f7416e8} /* (31, 12, 27) {real, imag} */,
  {32'h40970c87, 32'h40820d4c} /* (31, 12, 26) {real, imag} */,
  {32'hc0d676d3, 32'h3f94e044} /* (31, 12, 25) {real, imag} */,
  {32'hc08f5e00, 32'h40d6a04d} /* (31, 12, 24) {real, imag} */,
  {32'hc117340c, 32'h400274fa} /* (31, 12, 23) {real, imag} */,
  {32'hc0ee753e, 32'hc0f9e0f0} /* (31, 12, 22) {real, imag} */,
  {32'hbf2bcdf8, 32'hc0e9750a} /* (31, 12, 21) {real, imag} */,
  {32'hbf74fe24, 32'hc113d0f9} /* (31, 12, 20) {real, imag} */,
  {32'hc09568f4, 32'hc0974d7a} /* (31, 12, 19) {real, imag} */,
  {32'hc16dbcc2, 32'hc05f802c} /* (31, 12, 18) {real, imag} */,
  {32'hc18cbc1c, 32'hc10e150a} /* (31, 12, 17) {real, imag} */,
  {32'hc16f2fec, 32'hc06bd79a} /* (31, 12, 16) {real, imag} */,
  {32'hc085037c, 32'hbe250f10} /* (31, 12, 15) {real, imag} */,
  {32'hc0bc2c2b, 32'h3fa00676} /* (31, 12, 14) {real, imag} */,
  {32'hc0ec36ad, 32'hbc73c400} /* (31, 12, 13) {real, imag} */,
  {32'hc0e7018c, 32'hc0581348} /* (31, 12, 12) {real, imag} */,
  {32'hc0d87060, 32'hc0ecfc0a} /* (31, 12, 11) {real, imag} */,
  {32'hc088c4e5, 32'hc14191ef} /* (31, 12, 10) {real, imag} */,
  {32'hc01d2ec8, 32'hc0e33b2a} /* (31, 12, 9) {real, imag} */,
  {32'hbf8afc2c, 32'h40875a9f} /* (31, 12, 8) {real, imag} */,
  {32'hbec664e0, 32'hc0e70908} /* (31, 12, 7) {real, imag} */,
  {32'hbfb430c0, 32'hc0b94e58} /* (31, 12, 6) {real, imag} */,
  {32'hc0aa7a3a, 32'hc0a6304c} /* (31, 12, 5) {real, imag} */,
  {32'h3f437cac, 32'hc12bf204} /* (31, 12, 4) {real, imag} */,
  {32'h407dbe55, 32'hc02793ee} /* (31, 12, 3) {real, imag} */,
  {32'hc0ba131a, 32'h40c42c36} /* (31, 12, 2) {real, imag} */,
  {32'hbfbdf731, 32'hbfe0fb3d} /* (31, 12, 1) {real, imag} */,
  {32'h3fcf44b6, 32'h401831b0} /* (31, 12, 0) {real, imag} */,
  {32'hbfd448e6, 32'hc0eb6105} /* (31, 11, 31) {real, imag} */,
  {32'h4100f45c, 32'hc1705c53} /* (31, 11, 30) {real, imag} */,
  {32'h41804e44, 32'hc187cde4} /* (31, 11, 29) {real, imag} */,
  {32'h416b3882, 32'hc0af9f64} /* (31, 11, 28) {real, imag} */,
  {32'h41338662, 32'h3e8b7c20} /* (31, 11, 27) {real, imag} */,
  {32'h409cc61b, 32'h407be782} /* (31, 11, 26) {real, imag} */,
  {32'h40e012ac, 32'hbf82d340} /* (31, 11, 25) {real, imag} */,
  {32'h416a733c, 32'hc12955b8} /* (31, 11, 24) {real, imag} */,
  {32'h410420ee, 32'hc15785e5} /* (31, 11, 23) {real, imag} */,
  {32'h41025f5f, 32'hbfffd4d8} /* (31, 11, 22) {real, imag} */,
  {32'h406f938a, 32'h3f941b9c} /* (31, 11, 21) {real, imag} */,
  {32'hc0e1b720, 32'hbf71395c} /* (31, 11, 20) {real, imag} */,
  {32'hc11aca78, 32'h3f37eefe} /* (31, 11, 19) {real, imag} */,
  {32'hc1169da1, 32'hc0a2cb6f} /* (31, 11, 18) {real, imag} */,
  {32'hc058da61, 32'h3ded0d00} /* (31, 11, 17) {real, imag} */,
  {32'hc1023b3f, 32'h410fbc32} /* (31, 11, 16) {real, imag} */,
  {32'hc13fe85c, 32'h40b88cf8} /* (31, 11, 15) {real, imag} */,
  {32'hc0e390f4, 32'h3ec9cdf0} /* (31, 11, 14) {real, imag} */,
  {32'hc15fd3de, 32'hc0cf0afb} /* (31, 11, 13) {real, imag} */,
  {32'hc17bd7bc, 32'h41398843} /* (31, 11, 12) {real, imag} */,
  {32'hc0a256b8, 32'h40f2f482} /* (31, 11, 11) {real, imag} */,
  {32'h3fdd82e4, 32'hbfcfbace} /* (31, 11, 10) {real, imag} */,
  {32'h412cfb29, 32'hc103a2da} /* (31, 11, 9) {real, imag} */,
  {32'h418f326f, 32'hc0d50866} /* (31, 11, 8) {real, imag} */,
  {32'h41018209, 32'hc0c87421} /* (31, 11, 7) {real, imag} */,
  {32'h412c0247, 32'hc0b1a11f} /* (31, 11, 6) {real, imag} */,
  {32'h410c5352, 32'hc10291f7} /* (31, 11, 5) {real, imag} */,
  {32'h40fffd4a, 32'hc0bed4d0} /* (31, 11, 4) {real, imag} */,
  {32'h409022f0, 32'hc0fd0ca9} /* (31, 11, 3) {real, imag} */,
  {32'h40e789a1, 32'hc112b60e} /* (31, 11, 2) {real, imag} */,
  {32'h4150ac20, 32'h40a1b6d8} /* (31, 11, 1) {real, imag} */,
  {32'h40d2ede2, 32'h40e8d00c} /* (31, 11, 0) {real, imag} */,
  {32'h3f43f5e8, 32'h3f509dfc} /* (31, 10, 31) {real, imag} */,
  {32'h408c55a3, 32'h40e32c2a} /* (31, 10, 30) {real, imag} */,
  {32'hc07dbba0, 32'h405a7db2} /* (31, 10, 29) {real, imag} */,
  {32'hc069e63b, 32'hc0d78bfa} /* (31, 10, 28) {real, imag} */,
  {32'hbfa3bae4, 32'hc0ebb490} /* (31, 10, 27) {real, imag} */,
  {32'hc0dab460, 32'h3f59dc98} /* (31, 10, 26) {real, imag} */,
  {32'hbfc90380, 32'h4069a852} /* (31, 10, 25) {real, imag} */,
  {32'hc04b0b00, 32'h3f22a8a0} /* (31, 10, 24) {real, imag} */,
  {32'hc0d4167f, 32'hc130222c} /* (31, 10, 23) {real, imag} */,
  {32'hbf9fe410, 32'hc0e1bcfc} /* (31, 10, 22) {real, imag} */,
  {32'hc0059de2, 32'hbfb8b330} /* (31, 10, 21) {real, imag} */,
  {32'hbf9a898c, 32'hc11b8e3a} /* (31, 10, 20) {real, imag} */,
  {32'hbfff5d48, 32'hc1254062} /* (31, 10, 19) {real, imag} */,
  {32'h40a0a176, 32'hc11007c5} /* (31, 10, 18) {real, imag} */,
  {32'h4137a0d1, 32'hc0e8d7de} /* (31, 10, 17) {real, imag} */,
  {32'h4033cd8f, 32'hc0fedfa1} /* (31, 10, 16) {real, imag} */,
  {32'hc09c2b7d, 32'hbf9d25bc} /* (31, 10, 15) {real, imag} */,
  {32'h411fa5c6, 32'h40bc04ec} /* (31, 10, 14) {real, imag} */,
  {32'h4153baa2, 32'h404a2294} /* (31, 10, 13) {real, imag} */,
  {32'h408854c7, 32'hc0ea6b12} /* (31, 10, 12) {real, imag} */,
  {32'h405ccd62, 32'h3ef6c498} /* (31, 10, 11) {real, imag} */,
  {32'hc00bad1c, 32'hbf610fa8} /* (31, 10, 10) {real, imag} */,
  {32'hc133ed72, 32'hc0b1df0a} /* (31, 10, 9) {real, imag} */,
  {32'hc17f81d2, 32'hbff39fa0} /* (31, 10, 8) {real, imag} */,
  {32'hc1220b76, 32'h3f335e58} /* (31, 10, 7) {real, imag} */,
  {32'hc1288081, 32'h3f290d00} /* (31, 10, 6) {real, imag} */,
  {32'hc126fbb1, 32'hc12e3d18} /* (31, 10, 5) {real, imag} */,
  {32'hc11cdd4a, 32'hc15171aa} /* (31, 10, 4) {real, imag} */,
  {32'hc140f842, 32'hc0cc97b0} /* (31, 10, 3) {real, imag} */,
  {32'hc1092922, 32'h3f8a2d64} /* (31, 10, 2) {real, imag} */,
  {32'hc1449d72, 32'h413b8dba} /* (31, 10, 1) {real, imag} */,
  {32'hc044f5b1, 32'h409c8c84} /* (31, 10, 0) {real, imag} */,
  {32'hc0c61236, 32'h4041407c} /* (31, 9, 31) {real, imag} */,
  {32'hc168937a, 32'h412f1af0} /* (31, 9, 30) {real, imag} */,
  {32'hc0fb4a0a, 32'hc0693bea} /* (31, 9, 29) {real, imag} */,
  {32'hc09e3cc2, 32'hc0c7cb03} /* (31, 9, 28) {real, imag} */,
  {32'h4057d746, 32'h412e5c45} /* (31, 9, 27) {real, imag} */,
  {32'h40dc64a8, 32'h40f8227e} /* (31, 9, 26) {real, imag} */,
  {32'hc0fcd53d, 32'h41033d96} /* (31, 9, 25) {real, imag} */,
  {32'hc13f7b36, 32'hc155b361} /* (31, 9, 24) {real, imag} */,
  {32'hc140750d, 32'hc0864c78} /* (31, 9, 23) {real, imag} */,
  {32'hc1b5b352, 32'h41152e62} /* (31, 9, 22) {real, imag} */,
  {32'hc156dd4a, 32'h4116a14e} /* (31, 9, 21) {real, imag} */,
  {32'h41391602, 32'h413a8240} /* (31, 9, 20) {real, imag} */,
  {32'h418bad13, 32'hc154a4c6} /* (31, 9, 19) {real, imag} */,
  {32'h41d3f404, 32'hc146ee8e} /* (31, 9, 18) {real, imag} */,
  {32'h41fc8e18, 32'hc0250986} /* (31, 9, 17) {real, imag} */,
  {32'h4218321a, 32'h40a87550} /* (31, 9, 16) {real, imag} */,
  {32'h414e6a2d, 32'hc0da7d1d} /* (31, 9, 15) {real, imag} */,
  {32'hbd9c7f40, 32'h40808c54} /* (31, 9, 14) {real, imag} */,
  {32'hc1246a2c, 32'h403fc384} /* (31, 9, 13) {real, imag} */,
  {32'hc1352227, 32'hc1095420} /* (31, 9, 12) {real, imag} */,
  {32'hc1ce5b8e, 32'h40043cec} /* (31, 9, 11) {real, imag} */,
  {32'hc1b4663a, 32'h418837ed} /* (31, 9, 10) {real, imag} */,
  {32'hc1893638, 32'h41557236} /* (31, 9, 9) {real, imag} */,
  {32'hc132a036, 32'hc0cf2476} /* (31, 9, 8) {real, imag} */,
  {32'hc06cefc8, 32'hc130553e} /* (31, 9, 7) {real, imag} */,
  {32'h405f35fe, 32'h3fbd4994} /* (31, 9, 6) {real, imag} */,
  {32'hc0d670ec, 32'hc12a0fa1} /* (31, 9, 5) {real, imag} */,
  {32'hc161e730, 32'hc1a08868} /* (31, 9, 4) {real, imag} */,
  {32'hc0e70a98, 32'hc0cf7d55} /* (31, 9, 3) {real, imag} */,
  {32'hc087bfdb, 32'h40122456} /* (31, 9, 2) {real, imag} */,
  {32'h404b5974, 32'h3f7ed488} /* (31, 9, 1) {real, imag} */,
  {32'h3f95f338, 32'hc1231b5a} /* (31, 9, 0) {real, imag} */,
  {32'h403ee065, 32'hbfdd9ad2} /* (31, 8, 31) {real, imag} */,
  {32'h41310caf, 32'hc1af9dba} /* (31, 8, 30) {real, imag} */,
  {32'h41a3e692, 32'hc21a9657} /* (31, 8, 29) {real, imag} */,
  {32'h41e4e46b, 32'hc1b9fbd5} /* (31, 8, 28) {real, imag} */,
  {32'h417acf9b, 32'hc0f2bc69} /* (31, 8, 27) {real, imag} */,
  {32'h41528f8c, 32'hc10a1ae6} /* (31, 8, 26) {real, imag} */,
  {32'h4195df11, 32'hc044a504} /* (31, 8, 25) {real, imag} */,
  {32'h4047e3c2, 32'hc121e09d} /* (31, 8, 24) {real, imag} */,
  {32'hc08d2326, 32'hc1afad52} /* (31, 8, 23) {real, imag} */,
  {32'hc0dcc556, 32'hc209f6d8} /* (31, 8, 22) {real, imag} */,
  {32'hbe03b640, 32'h409c5e7c} /* (31, 8, 21) {real, imag} */,
  {32'hc0974629, 32'h421d2f66} /* (31, 8, 20) {real, imag} */,
  {32'hc08fb7dd, 32'h4206938f} /* (31, 8, 19) {real, imag} */,
  {32'hc13aa859, 32'h41cdc7c4} /* (31, 8, 18) {real, imag} */,
  {32'hc14910f3, 32'h41ffd148} /* (31, 8, 17) {real, imag} */,
  {32'hc144da26, 32'h41febf5e} /* (31, 8, 16) {real, imag} */,
  {32'h401ac7d2, 32'h41a5a92c} /* (31, 8, 15) {real, imag} */,
  {32'hc159b440, 32'h419f686d} /* (31, 8, 14) {real, imag} */,
  {32'hbff475f8, 32'h41e3e422} /* (31, 8, 13) {real, imag} */,
  {32'hc10e802c, 32'h419a0239} /* (31, 8, 12) {real, imag} */,
  {32'hc1248db0, 32'h41423432} /* (31, 8, 11) {real, imag} */,
  {32'hbee182ec, 32'hc13f308b} /* (31, 8, 10) {real, imag} */,
  {32'hbe3e94f0, 32'hc1e4fccc} /* (31, 8, 9) {real, imag} */,
  {32'h3f1b5aa8, 32'hc1b3288c} /* (31, 8, 8) {real, imag} */,
  {32'h4114371e, 32'hc18d1a65} /* (31, 8, 7) {real, imag} */,
  {32'hbf48b138, 32'hc1def9b5} /* (31, 8, 6) {real, imag} */,
  {32'hc107156a, 32'hc1db696b} /* (31, 8, 5) {real, imag} */,
  {32'hc173b4ab, 32'hc193ae95} /* (31, 8, 4) {real, imag} */,
  {32'h4096aa50, 32'hc192539f} /* (31, 8, 3) {real, imag} */,
  {32'h41ba69d5, 32'hc123fa20} /* (31, 8, 2) {real, imag} */,
  {32'h417812da, 32'hc0de3c24} /* (31, 8, 1) {real, imag} */,
  {32'h3fae24e6, 32'hbfa7b3fe} /* (31, 8, 0) {real, imag} */,
  {32'hbfbf93d2, 32'hc0b27d28} /* (31, 7, 31) {real, imag} */,
  {32'hc1aba056, 32'hc111b7ba} /* (31, 7, 30) {real, imag} */,
  {32'hc2002ff5, 32'hc104350e} /* (31, 7, 29) {real, imag} */,
  {32'h401b56f0, 32'hc00cac42} /* (31, 7, 28) {real, imag} */,
  {32'hc10743a6, 32'h4183dcf7} /* (31, 7, 27) {real, imag} */,
  {32'hc1de3adf, 32'h418570eb} /* (31, 7, 26) {real, imag} */,
  {32'hc16c516c, 32'hc15c2a5a} /* (31, 7, 25) {real, imag} */,
  {32'hc1110923, 32'hc19a6440} /* (31, 7, 24) {real, imag} */,
  {32'hc1b5130c, 32'hbff8a5e0} /* (31, 7, 23) {real, imag} */,
  {32'hc1875ea4, 32'hbfda8850} /* (31, 7, 22) {real, imag} */,
  {32'h40837249, 32'hc0609b20} /* (31, 7, 21) {real, imag} */,
  {32'h40ac1421, 32'h4141d7fe} /* (31, 7, 20) {real, imag} */,
  {32'h416b7008, 32'h407373a4} /* (31, 7, 19) {real, imag} */,
  {32'h408af884, 32'hc0bcaf00} /* (31, 7, 18) {real, imag} */,
  {32'h4091d58e, 32'hc0286b16} /* (31, 7, 17) {real, imag} */,
  {32'h4104d268, 32'hc11e8605} /* (31, 7, 16) {real, imag} */,
  {32'h3fc48da0, 32'hc011fff8} /* (31, 7, 15) {real, imag} */,
  {32'h4122238a, 32'h3ec5cea0} /* (31, 7, 14) {real, imag} */,
  {32'h411b20b2, 32'h4104092a} /* (31, 7, 13) {real, imag} */,
  {32'h414f9da7, 32'hbf089de8} /* (31, 7, 12) {real, imag} */,
  {32'h41db2e6c, 32'hc15cdc5c} /* (31, 7, 11) {real, imag} */,
  {32'h414085dc, 32'hc1886a81} /* (31, 7, 10) {real, imag} */,
  {32'h4044e570, 32'hc1063d26} /* (31, 7, 9) {real, imag} */,
  {32'hc0df691d, 32'hc1a6c0fc} /* (31, 7, 8) {real, imag} */,
  {32'h4028a430, 32'hbf9dcfd4} /* (31, 7, 7) {real, imag} */,
  {32'h41613f49, 32'h417dea2e} /* (31, 7, 6) {real, imag} */,
  {32'h41b2c79c, 32'h41c587f4} /* (31, 7, 5) {real, imag} */,
  {32'h4147831b, 32'h4199a53c} /* (31, 7, 4) {real, imag} */,
  {32'h416bb510, 32'h418c4557} /* (31, 7, 3) {real, imag} */,
  {32'hc0cb895b, 32'hc114132a} /* (31, 7, 2) {real, imag} */,
  {32'hc12a8530, 32'h3f3fe170} /* (31, 7, 1) {real, imag} */,
  {32'hc0a48e8a, 32'h404ce9d1} /* (31, 7, 0) {real, imag} */,
  {32'hc0ef901e, 32'h40bb0c70} /* (31, 6, 31) {real, imag} */,
  {32'hc1e28df0, 32'h3f159670} /* (31, 6, 30) {real, imag} */,
  {32'hc1a4b393, 32'h40d93fb3} /* (31, 6, 29) {real, imag} */,
  {32'hc16cec8c, 32'h4103a0d9} /* (31, 6, 28) {real, imag} */,
  {32'hc1e34616, 32'h41efdb06} /* (31, 6, 27) {real, imag} */,
  {32'hc0d802f0, 32'h41a06230} /* (31, 6, 26) {real, imag} */,
  {32'h3e276100, 32'hc0c1b9b7} /* (31, 6, 25) {real, imag} */,
  {32'h411b9b81, 32'hc1f20691} /* (31, 6, 24) {real, imag} */,
  {32'h41919cee, 32'hc108decb} /* (31, 6, 23) {real, imag} */,
  {32'h40213cb6, 32'hc18e999e} /* (31, 6, 22) {real, imag} */,
  {32'hc0c8b210, 32'hbfffb480} /* (31, 6, 21) {real, imag} */,
  {32'h40a24012, 32'h41814ffc} /* (31, 6, 20) {real, imag} */,
  {32'h4175c0d3, 32'h4092cb42} /* (31, 6, 19) {real, imag} */,
  {32'h411c2c13, 32'hc0a4cc1e} /* (31, 6, 18) {real, imag} */,
  {32'h404b0eb8, 32'hc189cdb8} /* (31, 6, 17) {real, imag} */,
  {32'h40e821a8, 32'hc14da604} /* (31, 6, 16) {real, imag} */,
  {32'hc05f5c18, 32'hc15e1be3} /* (31, 6, 15) {real, imag} */,
  {32'h4115921a, 32'hc184f12c} /* (31, 6, 14) {real, imag} */,
  {32'h40ffcafc, 32'hbf6e07a0} /* (31, 6, 13) {real, imag} */,
  {32'h405485da, 32'hc13454c7} /* (31, 6, 12) {real, imag} */,
  {32'hc12bfa88, 32'hc121e88a} /* (31, 6, 11) {real, imag} */,
  {32'hc11cb330, 32'hbfcbb114} /* (31, 6, 10) {real, imag} */,
  {32'h40f5fefc, 32'h4152c37f} /* (31, 6, 9) {real, imag} */,
  {32'h4138cc0c, 32'h400b42b7} /* (31, 6, 8) {real, imag} */,
  {32'h4101a136, 32'h3f20ab78} /* (31, 6, 7) {real, imag} */,
  {32'h410d9dbf, 32'hc0c9fc44} /* (31, 6, 6) {real, imag} */,
  {32'h40c0666a, 32'h41554300} /* (31, 6, 5) {real, imag} */,
  {32'h41bec875, 32'h4136d256} /* (31, 6, 4) {real, imag} */,
  {32'h413c7d3a, 32'hc15d74b8} /* (31, 6, 3) {real, imag} */,
  {32'h410d3217, 32'hc1dc086a} /* (31, 6, 2) {real, imag} */,
  {32'h40b46b68, 32'h40058b02} /* (31, 6, 1) {real, imag} */,
  {32'hc00a5391, 32'h4166bff4} /* (31, 6, 0) {real, imag} */,
  {32'h416ffafc, 32'hc1d6f485} /* (31, 5, 31) {real, imag} */,
  {32'h4196caac, 32'hc22007bb} /* (31, 5, 30) {real, imag} */,
  {32'h421198a8, 32'hc1bb9812} /* (31, 5, 29) {real, imag} */,
  {32'h4205e088, 32'hc1a020f7} /* (31, 5, 28) {real, imag} */,
  {32'h41b57afb, 32'hc1f99c45} /* (31, 5, 27) {real, imag} */,
  {32'h4193f14c, 32'hc1bc5a88} /* (31, 5, 26) {real, imag} */,
  {32'h41f58eb3, 32'hc1edf584} /* (31, 5, 25) {real, imag} */,
  {32'h422c6785, 32'hc1f30c62} /* (31, 5, 24) {real, imag} */,
  {32'h417f1560, 32'hc2375c31} /* (31, 5, 23) {real, imag} */,
  {32'h3f151c50, 32'hc244cfe2} /* (31, 5, 22) {real, imag} */,
  {32'h416c88a8, 32'hc2169267} /* (31, 5, 21) {real, imag} */,
  {32'h4147cd09, 32'hbdeb4820} /* (31, 5, 20) {real, imag} */,
  {32'hc0448176, 32'h40e23c03} /* (31, 5, 19) {real, imag} */,
  {32'hc0a14ca6, 32'h418071ba} /* (31, 5, 18) {real, imag} */,
  {32'h3fbdb540, 32'h4194b069} /* (31, 5, 17) {real, imag} */,
  {32'h414fd9c1, 32'h41dfcf78} /* (31, 5, 16) {real, imag} */,
  {32'h403fbf48, 32'h4246a5dd} /* (31, 5, 15) {real, imag} */,
  {32'hc0baaf58, 32'h42061fac} /* (31, 5, 14) {real, imag} */,
  {32'hc0d49594, 32'h41de3f04} /* (31, 5, 13) {real, imag} */,
  {32'hc1b3eb89, 32'h41f3596b} /* (31, 5, 12) {real, imag} */,
  {32'hc1c27943, 32'h41d21e5b} /* (31, 5, 11) {real, imag} */,
  {32'h414cb812, 32'h3def7980} /* (31, 5, 10) {real, imag} */,
  {32'h40fee3f2, 32'hc16de018} /* (31, 5, 9) {real, imag} */,
  {32'h40b5a96c, 32'hc08d5988} /* (31, 5, 8) {real, imag} */,
  {32'h414ef312, 32'hc022b75a} /* (31, 5, 7) {real, imag} */,
  {32'h40d95d4f, 32'hc0fdbf13} /* (31, 5, 6) {real, imag} */,
  {32'h41a2b97a, 32'hc190b10c} /* (31, 5, 5) {real, imag} */,
  {32'h405f07c8, 32'hc1c75136} /* (31, 5, 4) {real, imag} */,
  {32'hc130bf10, 32'hc1750e58} /* (31, 5, 3) {real, imag} */,
  {32'h4137f6d6, 32'hc1afc943} /* (31, 5, 2) {real, imag} */,
  {32'h40d4a6e8, 32'hc242994b} /* (31, 5, 1) {real, imag} */,
  {32'hc083c717, 32'hc213d4fe} /* (31, 5, 0) {real, imag} */,
  {32'hc0cc0e2f, 32'h40fe323f} /* (31, 4, 31) {real, imag} */,
  {32'hc1aa9fd1, 32'h41988e32} /* (31, 4, 30) {real, imag} */,
  {32'hc18b6b26, 32'h422bbbe6} /* (31, 4, 29) {real, imag} */,
  {32'hc13f6e40, 32'h422ee641} /* (31, 4, 28) {real, imag} */,
  {32'h419bc289, 32'h41c08d2e} /* (31, 4, 27) {real, imag} */,
  {32'h41dbc56e, 32'h41892f84} /* (31, 4, 26) {real, imag} */,
  {32'h4120a4bc, 32'h4197ce8e} /* (31, 4, 25) {real, imag} */,
  {32'hc1a7e313, 32'h4148b60f} /* (31, 4, 24) {real, imag} */,
  {32'hbecdf200, 32'h41d8320e} /* (31, 4, 23) {real, imag} */,
  {32'h403c3578, 32'h41aa8687} /* (31, 4, 22) {real, imag} */,
  {32'h414ec89b, 32'h41bcc99a} /* (31, 4, 21) {real, imag} */,
  {32'h42666fce, 32'hc19a728c} /* (31, 4, 20) {real, imag} */,
  {32'h423200f0, 32'hc22a37cc} /* (31, 4, 19) {real, imag} */,
  {32'h424a53ed, 32'hc207da6c} /* (31, 4, 18) {real, imag} */,
  {32'h422a4b40, 32'hc256c69b} /* (31, 4, 17) {real, imag} */,
  {32'h42019c46, 32'hc246c6b6} /* (31, 4, 16) {real, imag} */,
  {32'h420c87fb, 32'hc19a3233} /* (31, 4, 15) {real, imag} */,
  {32'h41cc84fb, 32'hc16a43de} /* (31, 4, 14) {real, imag} */,
  {32'h416d2a71, 32'hc1d42987} /* (31, 4, 13) {real, imag} */,
  {32'h41bbee7b, 32'hc1310cb1} /* (31, 4, 12) {real, imag} */,
  {32'h40bf2ea0, 32'hc0f5d2ce} /* (31, 4, 11) {real, imag} */,
  {32'hc1c09086, 32'h41922510} /* (31, 4, 10) {real, imag} */,
  {32'hc14e930d, 32'h42265950} /* (31, 4, 9) {real, imag} */,
  {32'hc2087aea, 32'h42450105} /* (31, 4, 8) {real, imag} */,
  {32'hc2259125, 32'h4231abbe} /* (31, 4, 7) {real, imag} */,
  {32'hc1d12ec4, 32'h4238acf7} /* (31, 4, 6) {real, imag} */,
  {32'hc17dbbdd, 32'h41cbdfab} /* (31, 4, 5) {real, imag} */,
  {32'h40f8d6ee, 32'h415402c4} /* (31, 4, 4) {real, imag} */,
  {32'h41156b42, 32'h41995292} /* (31, 4, 3) {real, imag} */,
  {32'hc116dbd8, 32'h41cd425c} /* (31, 4, 2) {real, imag} */,
  {32'hc16ee546, 32'h41cad78a} /* (31, 4, 1) {real, imag} */,
  {32'h4090c686, 32'h41a9a3b0} /* (31, 4, 0) {real, imag} */,
  {32'hc0bf43be, 32'h407d8cfa} /* (31, 3, 31) {real, imag} */,
  {32'h403495d2, 32'h417131c0} /* (31, 3, 30) {real, imag} */,
  {32'h416435e5, 32'h41cad6c2} /* (31, 3, 29) {real, imag} */,
  {32'h40b14360, 32'h41c755db} /* (31, 3, 28) {real, imag} */,
  {32'h4105b56c, 32'h41214b18} /* (31, 3, 27) {real, imag} */,
  {32'hbf1d7464, 32'hc1347230} /* (31, 3, 26) {real, imag} */,
  {32'h41aa2333, 32'h419d4076} /* (31, 3, 25) {real, imag} */,
  {32'h414ce73c, 32'h4081866f} /* (31, 3, 24) {real, imag} */,
  {32'h40c106ca, 32'hc14c546f} /* (31, 3, 23) {real, imag} */,
  {32'h3e36da80, 32'hc1c77194} /* (31, 3, 22) {real, imag} */,
  {32'h40f32101, 32'hc1d62784} /* (31, 3, 21) {real, imag} */,
  {32'h42085917, 32'hc1bf0e20} /* (31, 3, 20) {real, imag} */,
  {32'h4200affc, 32'hc0e5bbcb} /* (31, 3, 19) {real, imag} */,
  {32'h42816137, 32'hc160f246} /* (31, 3, 18) {real, imag} */,
  {32'h42517a2c, 32'hc1197b03} /* (31, 3, 17) {real, imag} */,
  {32'h42023acc, 32'h4106946d} /* (31, 3, 16) {real, imag} */,
  {32'h4111983e, 32'h40a1e3f0} /* (31, 3, 15) {real, imag} */,
  {32'h4116a37f, 32'hc1864337} /* (31, 3, 14) {real, imag} */,
  {32'h419af319, 32'hc1ea4759} /* (31, 3, 13) {real, imag} */,
  {32'hc165bfe5, 32'hc1171d78} /* (31, 3, 12) {real, imag} */,
  {32'h40ad8ee4, 32'h4047107c} /* (31, 3, 11) {real, imag} */,
  {32'hc093eaf4, 32'hc0835668} /* (31, 3, 10) {real, imag} */,
  {32'hc20f94d0, 32'h40521108} /* (31, 3, 9) {real, imag} */,
  {32'hc2911657, 32'hbfa41eb0} /* (31, 3, 8) {real, imag} */,
  {32'hc280653d, 32'h403bf572} /* (31, 3, 7) {real, imag} */,
  {32'hc2679371, 32'hc137049e} /* (31, 3, 6) {real, imag} */,
  {32'hc236eee4, 32'hc0727c6c} /* (31, 3, 5) {real, imag} */,
  {32'h401e0aff, 32'hc0663aec} /* (31, 3, 4) {real, imag} */,
  {32'h4025f814, 32'h40d3aeb2} /* (31, 3, 3) {real, imag} */,
  {32'hbf1ad6d0, 32'hc13e5b40} /* (31, 3, 2) {real, imag} */,
  {32'hbf6227e4, 32'hc1290e4a} /* (31, 3, 1) {real, imag} */,
  {32'hc0635a77, 32'hbfd56966} /* (31, 3, 0) {real, imag} */,
  {32'hc1555b7d, 32'hc1efb520} /* (31, 2, 31) {real, imag} */,
  {32'hc1026304, 32'hc2a5249a} /* (31, 2, 30) {real, imag} */,
  {32'h40106bb0, 32'hc2c32d6b} /* (31, 2, 29) {real, imag} */,
  {32'h421667cc, 32'hc2a9fa5e} /* (31, 2, 28) {real, imag} */,
  {32'h41d9e4a3, 32'hc28c31c6} /* (31, 2, 27) {real, imag} */,
  {32'h40446620, 32'hc290ace2} /* (31, 2, 26) {real, imag} */,
  {32'h402fe302, 32'hc2a7bfc5} /* (31, 2, 25) {real, imag} */,
  {32'h40646630, 32'hc276c3cc} /* (31, 2, 24) {real, imag} */,
  {32'h408ba4f0, 32'hc2b1ba64} /* (31, 2, 23) {real, imag} */,
  {32'h40ff1ede, 32'hc2d44bcc} /* (31, 2, 22) {real, imag} */,
  {32'h40109200, 32'hc22733ca} /* (31, 2, 21) {real, imag} */,
  {32'h42195c26, 32'h428d8a43} /* (31, 2, 20) {real, imag} */,
  {32'h426faa49, 32'h42ec1404} /* (31, 2, 19) {real, imag} */,
  {32'h4285246f, 32'h42cb2923} /* (31, 2, 18) {real, imag} */,
  {32'h42882762, 32'h42d040ee} /* (31, 2, 17) {real, imag} */,
  {32'h4250cdac, 32'h42f11320} /* (31, 2, 16) {real, imag} */,
  {32'h41aaedba, 32'h42bd929c} /* (31, 2, 15) {real, imag} */,
  {32'h4171229a, 32'h42a16479} /* (31, 2, 14) {real, imag} */,
  {32'h3de20300, 32'h42986552} /* (31, 2, 13) {real, imag} */,
  {32'hc1fc7664, 32'h4292c45d} /* (31, 2, 12) {real, imag} */,
  {32'hc20531dd, 32'h42110db5} /* (31, 2, 11) {real, imag} */,
  {32'hc22ec43e, 32'hc2888c4c} /* (31, 2, 10) {real, imag} */,
  {32'hc2819f3b, 32'hc2de442b} /* (31, 2, 9) {real, imag} */,
  {32'hc28a1aaa, 32'hc2d347b0} /* (31, 2, 8) {real, imag} */,
  {32'hc24ba52b, 32'hc2f1901c} /* (31, 2, 7) {real, imag} */,
  {32'hc20933b8, 32'hc2e38978} /* (31, 2, 6) {real, imag} */,
  {32'hc120f5a0, 32'hc2ca3610} /* (31, 2, 5) {real, imag} */,
  {32'hc11f66b2, 32'hc2b29997} /* (31, 2, 4) {real, imag} */,
  {32'hc09065f6, 32'hc2c4c7f6} /* (31, 2, 3) {real, imag} */,
  {32'h407d080c, 32'hc2b7ad94} /* (31, 2, 2) {real, imag} */,
  {32'hc0abc1be, 32'hc29feeb7} /* (31, 2, 1) {real, imag} */,
  {32'hc0218c68, 32'hc21d1689} /* (31, 2, 0) {real, imag} */,
  {32'h40fe3a1e, 32'h4287bfe2} /* (31, 1, 31) {real, imag} */,
  {32'hc102f266, 32'h42ff857e} /* (31, 1, 30) {real, imag} */,
  {32'hc0966826, 32'h42e6925d} /* (31, 1, 29) {real, imag} */,
  {32'hc1bdb205, 32'h43051dff} /* (31, 1, 28) {real, imag} */,
  {32'hbff75238, 32'h431a7bed} /* (31, 1, 27) {real, imag} */,
  {32'hc13d6bb6, 32'h43144a15} /* (31, 1, 26) {real, imag} */,
  {32'hc162884e, 32'h430198fd} /* (31, 1, 25) {real, imag} */,
  {32'h411619c0, 32'h4321730e} /* (31, 1, 24) {real, imag} */,
  {32'hc09617be, 32'h431b6b24} /* (31, 1, 23) {real, imag} */,
  {32'h4030c6c1, 32'h43061403} /* (31, 1, 22) {real, imag} */,
  {32'h4220d41b, 32'h42867dce} /* (31, 1, 21) {real, imag} */,
  {32'h424787ee, 32'hc23fb45f} /* (31, 1, 20) {real, imag} */,
  {32'h4254d24b, 32'hc26628ee} /* (31, 1, 19) {real, imag} */,
  {32'h42467def, 32'hc257f18f} /* (31, 1, 18) {real, imag} */,
  {32'h4275313d, 32'hc21b92d1} /* (31, 1, 17) {real, imag} */,
  {32'h41dcd60e, 32'hc286046b} /* (31, 1, 16) {real, imag} */,
  {32'hc1a223cc, 32'hc30143e6} /* (31, 1, 15) {real, imag} */,
  {32'hc1c9d95a, 32'hc30d372c} /* (31, 1, 14) {real, imag} */,
  {32'hbda77700, 32'hc2f22098} /* (31, 1, 13) {real, imag} */,
  {32'h411a68d4, 32'hc30419c0} /* (31, 1, 12) {real, imag} */,
  {32'hc17be537, 32'hc2b37d18} /* (31, 1, 11) {real, imag} */,
  {32'hc27136b6, 32'h42068a5b} /* (31, 1, 10) {real, imag} */,
  {32'hc239fc61, 32'h425fec9c} /* (31, 1, 9) {real, imag} */,
  {32'hc1b7e968, 32'h428fdc39} /* (31, 1, 8) {real, imag} */,
  {32'hc2720c48, 32'h4292e94e} /* (31, 1, 7) {real, imag} */,
  {32'hc2733e16, 32'h42978d5f} /* (31, 1, 6) {real, imag} */,
  {32'hc1ea5f0b, 32'h42bc78b4} /* (31, 1, 5) {real, imag} */,
  {32'hc0f8406c, 32'h42f10d4a} /* (31, 1, 4) {real, imag} */,
  {32'h41c6d9e8, 32'h430e05ee} /* (31, 1, 3) {real, imag} */,
  {32'h41cd6e86, 32'h430ca99f} /* (31, 1, 2) {real, imag} */,
  {32'h41122bee, 32'h4310d6de} /* (31, 1, 1) {real, imag} */,
  {32'h403e2692, 32'h4287f0f0} /* (31, 1, 0) {real, imag} */,
  {32'h4131d7af, 32'h4221f908} /* (31, 0, 31) {real, imag} */,
  {32'h41ade2fd, 32'h4291ba95} /* (31, 0, 30) {real, imag} */,
  {32'h4106fe6c, 32'h42c4cd4f} /* (31, 0, 29) {real, imag} */,
  {32'hc1358670, 32'h42bf6c40} /* (31, 0, 28) {real, imag} */,
  {32'h3fa5a3a8, 32'h42b1ea37} /* (31, 0, 27) {real, imag} */,
  {32'h406ec97f, 32'h4294b312} /* (31, 0, 26) {real, imag} */,
  {32'h40d7c44d, 32'h42ae4994} /* (31, 0, 25) {real, imag} */,
  {32'hc0111d99, 32'h4296804d} /* (31, 0, 24) {real, imag} */,
  {32'h41b1b26c, 32'h4293a006} /* (31, 0, 23) {real, imag} */,
  {32'h416f4f02, 32'h42bd0aa4} /* (31, 0, 22) {real, imag} */,
  {32'h4158225e, 32'h42ac5ade} /* (31, 0, 21) {real, imag} */,
  {32'h40fcf7fd, 32'h41b5040d} /* (31, 0, 20) {real, imag} */,
  {32'h4117ec6a, 32'h40889871} /* (31, 0, 19) {real, imag} */,
  {32'h40d30719, 32'hc164ad78} /* (31, 0, 18) {real, imag} */,
  {32'hbfaaba1c, 32'h40b09712} /* (31, 0, 17) {real, imag} */,
  {32'hc1031170, 32'hc1cd91ff} /* (31, 0, 16) {real, imag} */,
  {32'hc1a218fc, 32'hc29c0335} /* (31, 0, 15) {real, imag} */,
  {32'hc1c0fcf2, 32'hc2b73143} /* (31, 0, 14) {real, imag} */,
  {32'hc1802526, 32'hc2a4a3c1} /* (31, 0, 13) {real, imag} */,
  {32'hc106f944, 32'hc297793c} /* (31, 0, 12) {real, imag} */,
  {32'hc0c83fa6, 32'hc2830347} /* (31, 0, 11) {real, imag} */,
  {32'hbfa9e2f8, 32'hc186c7e6} /* (31, 0, 10) {real, imag} */,
  {32'hc15a7420, 32'hc14740c4} /* (31, 0, 9) {real, imag} */,
  {32'hc18bf2f1, 32'hc0bd627b} /* (31, 0, 8) {real, imag} */,
  {32'h41b78cc2, 32'hc110edda} /* (31, 0, 7) {real, imag} */,
  {32'h41c1723c, 32'hc1229046} /* (31, 0, 6) {real, imag} */,
  {32'hc004e60d, 32'h427e06d4} /* (31, 0, 5) {real, imag} */,
  {32'h40bf0006, 32'h429f4ae0} /* (31, 0, 4) {real, imag} */,
  {32'h403ccbe8, 32'h42a7323e} /* (31, 0, 3) {real, imag} */,
  {32'h41141feb, 32'h429c6652} /* (31, 0, 2) {real, imag} */,
  {32'h410ee7c4, 32'h42ae22c6} /* (31, 0, 1) {real, imag} */,
  {32'h4103450e, 32'h42122467} /* (31, 0, 0) {real, imag} */,
  {32'hc2147d98, 32'hc2f086b3} /* (30, 31, 31) {real, imag} */,
  {32'hc29ac48c, 32'hc36cda73} /* (30, 31, 30) {real, imag} */,
  {32'hc28b6680, 32'hc36f9c29} /* (30, 31, 29) {real, imag} */,
  {32'hc285b8a6, 32'hc3617a91} /* (30, 31, 28) {real, imag} */,
  {32'hc24a2efb, 32'hc368b315} /* (30, 31, 27) {real, imag} */,
  {32'hc22f865f, 32'hc35ee4f6} /* (30, 31, 26) {real, imag} */,
  {32'hc2894b27, 32'hc372acf0} /* (30, 31, 25) {real, imag} */,
  {32'hc290e5e1, 32'hc37c4021} /* (30, 31, 24) {real, imag} */,
  {32'hc2992670, 32'hc382bd82} /* (30, 31, 23) {real, imag} */,
  {32'hc2a2e42c, 32'hc37d7331} /* (30, 31, 22) {real, imag} */,
  {32'h3fc66cf0, 32'hc30cbe91} /* (30, 31, 21) {real, imag} */,
  {32'h42e974ee, 32'h416c869c} /* (30, 31, 20) {real, imag} */,
  {32'h42ebafd5, 32'h428cf800} /* (30, 31, 19) {real, imag} */,
  {32'h42a5fa56, 32'h42bc8306} /* (30, 31, 18) {real, imag} */,
  {32'h42e083fa, 32'h42c00546} /* (30, 31, 17) {real, imag} */,
  {32'h42e4f01e, 32'h430eea9f} /* (30, 31, 16) {real, imag} */,
  {32'h42a1ee87, 32'h435776e9} /* (30, 31, 15) {real, imag} */,
  {32'h42b77544, 32'h435e4733} /* (30, 31, 14) {real, imag} */,
  {32'h42b42b4a, 32'h436a7259} /* (30, 31, 13) {real, imag} */,
  {32'h42849470, 32'h436f6558} /* (30, 31, 12) {real, imag} */,
  {32'h41f2134b, 32'h4347866f} /* (30, 31, 11) {real, imag} */,
  {32'hc2a6115b, 32'h417580c6} /* (30, 31, 10) {real, imag} */,
  {32'hc30ae754, 32'hc29eb7fe} /* (30, 31, 9) {real, imag} */,
  {32'hc318cb3d, 32'hc2ba2547} /* (30, 31, 8) {real, imag} */,
  {32'hc305d7ea, 32'hc2b4fe3b} /* (30, 31, 7) {real, imag} */,
  {32'hc2b60a20, 32'hc2a267aa} /* (30, 31, 6) {real, imag} */,
  {32'hc2716cce, 32'hc33726b8} /* (30, 31, 5) {real, imag} */,
  {32'hc283a34e, 32'hc3628c53} /* (30, 31, 4) {real, imag} */,
  {32'hc2a93c34, 32'hc35a285e} /* (30, 31, 3) {real, imag} */,
  {32'hc2bd9034, 32'hc351ea00} /* (30, 31, 2) {real, imag} */,
  {32'hc2b6aeb8, 32'hc3526344} /* (30, 31, 1) {real, imag} */,
  {32'hc250013c, 32'hc3020bbe} /* (30, 31, 0) {real, imag} */,
  {32'h41c7c26c, 32'h42ab25eb} /* (30, 30, 31) {real, imag} */,
  {32'h42450fdc, 32'h430b2c4c} /* (30, 30, 30) {real, imag} */,
  {32'h426416a1, 32'h43106abd} /* (30, 30, 29) {real, imag} */,
  {32'h4256483c, 32'h4311260e} /* (30, 30, 28) {real, imag} */,
  {32'h426625fe, 32'h42f2adec} /* (30, 30, 27) {real, imag} */,
  {32'h42816e0e, 32'h42de7070} /* (30, 30, 26) {real, imag} */,
  {32'h41cba4ac, 32'h42e1b261} /* (30, 30, 25) {real, imag} */,
  {32'h41ea2ceb, 32'h43176ae0} /* (30, 30, 24) {real, imag} */,
  {32'h42362e27, 32'h43165076} /* (30, 30, 23) {real, imag} */,
  {32'h4270f4ac, 32'h430b881f} /* (30, 30, 22) {real, imag} */,
  {32'h427fff10, 32'h41ed41e0} /* (30, 30, 21) {real, imag} */,
  {32'h423fcb66, 32'hc33c2582} /* (30, 30, 20) {real, imag} */,
  {32'h41875dfc, 32'hc37107c4} /* (30, 30, 19) {real, imag} */,
  {32'h419abbe6, 32'hc379c95e} /* (30, 30, 18) {real, imag} */,
  {32'h419b0a1a, 32'hc37327b2} /* (30, 30, 17) {real, imag} */,
  {32'h41d530ba, 32'hc352a4ad} /* (30, 30, 16) {real, imag} */,
  {32'hc15aa462, 32'hc3298523} /* (30, 30, 15) {real, imag} */,
  {32'hc25d990e, 32'hc3072567} /* (30, 30, 14) {real, imag} */,
  {32'hc24c838a, 32'hc2d62f81} /* (30, 30, 13) {real, imag} */,
  {32'hc2034b30, 32'hc3092818} /* (30, 30, 12) {real, imag} */,
  {32'hc22ba564, 32'hc2ebe2de} /* (30, 30, 11) {real, imag} */,
  {32'hc1cd99d8, 32'h42be6a2b} /* (30, 30, 10) {real, imag} */,
  {32'hc1867300, 32'h43566cb3} /* (30, 30, 9) {real, imag} */,
  {32'hc18cd8ac, 32'h4375608e} /* (30, 30, 8) {real, imag} */,
  {32'hc1d15670, 32'h436ec957} /* (30, 30, 7) {real, imag} */,
  {32'hc26ea2ad, 32'h43505636} /* (30, 30, 6) {real, imag} */,
  {32'hc1e2b9c7, 32'h432d8b79} /* (30, 30, 5) {real, imag} */,
  {32'h41b986b2, 32'h4320c630} /* (30, 30, 4) {real, imag} */,
  {32'h427a3594, 32'h430af98a} /* (30, 30, 3) {real, imag} */,
  {32'h42984f2a, 32'h43017814} /* (30, 30, 2) {real, imag} */,
  {32'h429a42e4, 32'h42f4d5ca} /* (30, 30, 1) {real, imag} */,
  {32'h41d8d49e, 32'h42a9b5a1} /* (30, 30, 0) {real, imag} */,
  {32'hc0b00f34, 32'h3f248398} /* (30, 29, 31) {real, imag} */,
  {32'hbe97bae0, 32'hc1075c64} /* (30, 29, 30) {real, imag} */,
  {32'h411ba2d2, 32'h41476305} /* (30, 29, 29) {real, imag} */,
  {32'hc1391ec5, 32'h41a647b6} /* (30, 29, 28) {real, imag} */,
  {32'hc1c725c4, 32'h416ab6c8} /* (30, 29, 27) {real, imag} */,
  {32'hc1fa4780, 32'h408dad8f} /* (30, 29, 26) {real, imag} */,
  {32'hc1298258, 32'h41579ab5} /* (30, 29, 25) {real, imag} */,
  {32'h40cca29a, 32'h3feb7868} /* (30, 29, 24) {real, imag} */,
  {32'h41b71980, 32'hc12f886c} /* (30, 29, 23) {real, imag} */,
  {32'hc0db25a4, 32'h416f2c24} /* (30, 29, 22) {real, imag} */,
  {32'h40bd19ac, 32'h419fd47a} /* (30, 29, 21) {real, imag} */,
  {32'h428195ee, 32'h3d2c4640} /* (30, 29, 20) {real, imag} */,
  {32'h42b9dabb, 32'hc1f7a2ca} /* (30, 29, 19) {real, imag} */,
  {32'h4298eff0, 32'hc25e90fc} /* (30, 29, 18) {real, imag} */,
  {32'h42bcf8dc, 32'hc269786d} /* (30, 29, 17) {real, imag} */,
  {32'h4284f476, 32'hc212f5a6} /* (30, 29, 16) {real, imag} */,
  {32'h40d16338, 32'hc191de81} /* (30, 29, 15) {real, imag} */,
  {32'hc11e8df8, 32'hc1ca30b2} /* (30, 29, 14) {real, imag} */,
  {32'hc0c49757, 32'hbf5241a8} /* (30, 29, 13) {real, imag} */,
  {32'hc0e25b50, 32'h41607383} /* (30, 29, 12) {real, imag} */,
  {32'hc1a3ec74, 32'h4178e44a} /* (30, 29, 11) {real, imag} */,
  {32'hc297594d, 32'h41ab4f9b} /* (30, 29, 10) {real, imag} */,
  {32'hc2b6e1eb, 32'h41e2e10c} /* (30, 29, 9) {real, imag} */,
  {32'hc2a2831b, 32'h41cc9b21} /* (30, 29, 8) {real, imag} */,
  {32'hc2a58fa1, 32'h42160f93} /* (30, 29, 7) {real, imag} */,
  {32'hc2a6713d, 32'h422fca81} /* (30, 29, 6) {real, imag} */,
  {32'hc0eb9de4, 32'h4183b707} /* (30, 29, 5) {real, imag} */,
  {32'h415ec089, 32'hbdfbdb00} /* (30, 29, 4) {real, imag} */,
  {32'h40661c2d, 32'h4023c9da} /* (30, 29, 3) {real, imag} */,
  {32'h41bcc45a, 32'h40cc843f} /* (30, 29, 2) {real, imag} */,
  {32'h4136c774, 32'hc1b7f559} /* (30, 29, 1) {real, imag} */,
  {32'hc1017423, 32'hc146fe19} /* (30, 29, 0) {real, imag} */,
  {32'hc02794ad, 32'hc15a4f89} /* (30, 28, 31) {real, imag} */,
  {32'h40b55f90, 32'hc1914773} /* (30, 28, 30) {real, imag} */,
  {32'h40c02283, 32'hc1a0b084} /* (30, 28, 29) {real, imag} */,
  {32'hc055d921, 32'hc2001de0} /* (30, 28, 28) {real, imag} */,
  {32'hc0922e4b, 32'hc1815338} /* (30, 28, 27) {real, imag} */,
  {32'hc18afa2f, 32'hc195e9ea} /* (30, 28, 26) {real, imag} */,
  {32'hc1d55dbb, 32'hc2237dc3} /* (30, 28, 25) {real, imag} */,
  {32'hc182e186, 32'hc1f89dd2} /* (30, 28, 24) {real, imag} */,
  {32'hc1473c00, 32'hc1c824c6} /* (30, 28, 23) {real, imag} */,
  {32'hc0bbf98a, 32'hc240229e} /* (30, 28, 22) {real, imag} */,
  {32'h3f9cc4da, 32'h400dbc5c} /* (30, 28, 21) {real, imag} */,
  {32'h4257b2dc, 32'h423ff75c} /* (30, 28, 20) {real, imag} */,
  {32'h42a7d2fc, 32'h42403a24} /* (30, 28, 19) {real, imag} */,
  {32'h429c86cd, 32'h4240e0ec} /* (30, 28, 18) {real, imag} */,
  {32'h429ba9c2, 32'h42621882} /* (30, 28, 17) {real, imag} */,
  {32'h428b7ad8, 32'h4241ac54} /* (30, 28, 16) {real, imag} */,
  {32'h418074b8, 32'h421d5ca0} /* (30, 28, 15) {real, imag} */,
  {32'h41dfff8a, 32'h42362060} /* (30, 28, 14) {real, imag} */,
  {32'h41db0d11, 32'h42280d18} /* (30, 28, 13) {real, imag} */,
  {32'h4192532d, 32'h4233b258} /* (30, 28, 12) {real, imag} */,
  {32'h41210274, 32'h41f0866e} /* (30, 28, 11) {real, imag} */,
  {32'hc24e6b06, 32'hc17b25e2} /* (30, 28, 10) {real, imag} */,
  {32'hc2a1a9ea, 32'hc2481ae0} /* (30, 28, 9) {real, imag} */,
  {32'hc26e54cc, 32'hc249537c} /* (30, 28, 8) {real, imag} */,
  {32'hc281c138, 32'hc281ccfa} /* (30, 28, 7) {real, imag} */,
  {32'hc2a26870, 32'hc2298116} /* (30, 28, 6) {real, imag} */,
  {32'hc241d8ca, 32'hc20ac9e1} /* (30, 28, 5) {real, imag} */,
  {32'hc20920d9, 32'hc16c4e45} /* (30, 28, 4) {real, imag} */,
  {32'hc1bc31f2, 32'hc13b0158} /* (30, 28, 3) {real, imag} */,
  {32'hc173725c, 32'hc1d7060e} /* (30, 28, 2) {real, imag} */,
  {32'hc1a9c0ae, 32'hc25ad3d6} /* (30, 28, 1) {real, imag} */,
  {32'hc10aea1d, 32'hc1d3b3e7} /* (30, 28, 0) {real, imag} */,
  {32'h41729ebf, 32'h41ed9571} /* (30, 27, 31) {real, imag} */,
  {32'h421ef14c, 32'h4281a0db} /* (30, 27, 30) {real, imag} */,
  {32'h41de48bd, 32'h427365ea} /* (30, 27, 29) {real, imag} */,
  {32'h420aa974, 32'h428f962f} /* (30, 27, 28) {real, imag} */,
  {32'h41cc0ee0, 32'h425bf9ef} /* (30, 27, 27) {real, imag} */,
  {32'h41bc4b10, 32'h41f0b091} /* (30, 27, 26) {real, imag} */,
  {32'h416f2180, 32'h412fe088} /* (30, 27, 25) {real, imag} */,
  {32'h420f83a0, 32'h41b01644} /* (30, 27, 24) {real, imag} */,
  {32'h423db920, 32'h4205f333} /* (30, 27, 23) {real, imag} */,
  {32'h41ebc59e, 32'h4281a7a8} /* (30, 27, 22) {real, imag} */,
  {32'h4187e8e4, 32'h421467b3} /* (30, 27, 21) {real, imag} */,
  {32'hc0eef475, 32'hc1ecec48} /* (30, 27, 20) {real, imag} */,
  {32'hc18ef0a6, 32'hc2590142} /* (30, 27, 19) {real, imag} */,
  {32'hc139c97e, 32'hc240c42c} /* (30, 27, 18) {real, imag} */,
  {32'hc10d6e4a, 32'hc1740c17} /* (30, 27, 17) {real, imag} */,
  {32'hc1829f12, 32'hc102d4f2} /* (30, 27, 16) {real, imag} */,
  {32'hc2055203, 32'hc1688834} /* (30, 27, 15) {real, imag} */,
  {32'hc1f80be1, 32'hc1b43ade} /* (30, 27, 14) {real, imag} */,
  {32'hc195ff86, 32'hc200185e} /* (30, 27, 13) {real, imag} */,
  {32'hc1afa5fe, 32'hc2544fd4} /* (30, 27, 12) {real, imag} */,
  {32'hc1a00e73, 32'hc2461752} /* (30, 27, 11) {real, imag} */,
  {32'h414a3fd7, 32'h415096cc} /* (30, 27, 10) {real, imag} */,
  {32'h3eab2830, 32'h42232f6c} /* (30, 27, 9) {real, imag} */,
  {32'hc11ef188, 32'h41f2476e} /* (30, 27, 8) {real, imag} */,
  {32'h41a44b72, 32'h425250cd} /* (30, 27, 7) {real, imag} */,
  {32'h4125ee6f, 32'h41dcaef8} /* (30, 27, 6) {real, imag} */,
  {32'h41ba8a55, 32'h41f25fa7} /* (30, 27, 5) {real, imag} */,
  {32'h422095be, 32'h420a2c3d} /* (30, 27, 4) {real, imag} */,
  {32'h421e8f9a, 32'h42260d3e} /* (30, 27, 3) {real, imag} */,
  {32'h421c0633, 32'h4271e1de} /* (30, 27, 2) {real, imag} */,
  {32'h422884f3, 32'h426a0bdb} /* (30, 27, 1) {real, imag} */,
  {32'h418cf626, 32'h41a9102f} /* (30, 27, 0) {real, imag} */,
  {32'h407dea02, 32'h3f87dd44} /* (30, 26, 31) {real, imag} */,
  {32'h419254e8, 32'h41023a64} /* (30, 26, 30) {real, imag} */,
  {32'h40c34ed6, 32'hbfdffff4} /* (30, 26, 29) {real, imag} */,
  {32'hc00b33b6, 32'h40f4ccd2} /* (30, 26, 28) {real, imag} */,
  {32'hbf984b58, 32'h410d2ea4} /* (30, 26, 27) {real, imag} */,
  {32'hc0a2be58, 32'h413418d9} /* (30, 26, 26) {real, imag} */,
  {32'hc0cd8538, 32'h4186aeee} /* (30, 26, 25) {real, imag} */,
  {32'hc119bd81, 32'h40b908ee} /* (30, 26, 24) {real, imag} */,
  {32'hc10c5ec8, 32'h41a8aa16} /* (30, 26, 23) {real, imag} */,
  {32'hc186b752, 32'h4126de52} /* (30, 26, 22) {real, imag} */,
  {32'hc1963fe2, 32'hc0e816f0} /* (30, 26, 21) {real, imag} */,
  {32'hc182c73c, 32'hc1390940} /* (30, 26, 20) {real, imag} */,
  {32'h408e2e5d, 32'hc0c4fdb7} /* (30, 26, 19) {real, imag} */,
  {32'hbe7a23c0, 32'hc09f181c} /* (30, 26, 18) {real, imag} */,
  {32'h3ec52fd0, 32'hc18193fc} /* (30, 26, 17) {real, imag} */,
  {32'hc131b39a, 32'hc1503e12} /* (30, 26, 16) {real, imag} */,
  {32'hc15f4775, 32'hc156fbf8} /* (30, 26, 15) {real, imag} */,
  {32'h40d43f27, 32'h409544fe} /* (30, 26, 14) {real, imag} */,
  {32'hc000e556, 32'h41d6b9d4} /* (30, 26, 13) {real, imag} */,
  {32'hc16b9d50, 32'h40c1a208} /* (30, 26, 12) {real, imag} */,
  {32'h3f6c654c, 32'h40f646c4} /* (30, 26, 11) {real, imag} */,
  {32'h4110afd7, 32'h4187b004} /* (30, 26, 10) {real, imag} */,
  {32'h3f21dc80, 32'h40a0f250} /* (30, 26, 9) {real, imag} */,
  {32'hc0410148, 32'h3eac1480} /* (30, 26, 8) {real, imag} */,
  {32'h41058fca, 32'h40d2d540} /* (30, 26, 7) {real, imag} */,
  {32'h3f92b25c, 32'h41182ff3} /* (30, 26, 6) {real, imag} */,
  {32'hc025a611, 32'h40c0674e} /* (30, 26, 5) {real, imag} */,
  {32'h4118ee64, 32'h3f0b27d8} /* (30, 26, 4) {real, imag} */,
  {32'h40b618b8, 32'h40194cd8} /* (30, 26, 3) {real, imag} */,
  {32'hc0acc60f, 32'hc088ad24} /* (30, 26, 2) {real, imag} */,
  {32'hc0d235ee, 32'hc19061d0} /* (30, 26, 1) {real, imag} */,
  {32'hc1147e9a, 32'hc186b8fc} /* (30, 26, 0) {real, imag} */,
  {32'hc0ecd711, 32'hbf675104} /* (30, 25, 31) {real, imag} */,
  {32'hc1665fce, 32'hc15c9164} /* (30, 25, 30) {real, imag} */,
  {32'hc11701b1, 32'hc1789c92} /* (30, 25, 29) {real, imag} */,
  {32'hc18df5ed, 32'hc1c46f0d} /* (30, 25, 28) {real, imag} */,
  {32'hc1611d10, 32'hc1f652cb} /* (30, 25, 27) {real, imag} */,
  {32'h3f374570, 32'hc1b2605c} /* (30, 25, 26) {real, imag} */,
  {32'h3ede6138, 32'hc0f33f6b} /* (30, 25, 25) {real, imag} */,
  {32'hc15093cc, 32'hc1c0c87c} /* (30, 25, 24) {real, imag} */,
  {32'hc159b606, 32'hc1ccc9fe} /* (30, 25, 23) {real, imag} */,
  {32'hc079e385, 32'hc07881b8} /* (30, 25, 22) {real, imag} */,
  {32'h40afd6ef, 32'h40798776} /* (30, 25, 21) {real, imag} */,
  {32'hc0068ffe, 32'h407957de} /* (30, 25, 20) {real, imag} */,
  {32'hc103d933, 32'h41229c8d} /* (30, 25, 19) {real, imag} */,
  {32'h409edc5e, 32'h40b1b14d} /* (30, 25, 18) {real, imag} */,
  {32'h40a5fa92, 32'h3efb9ed8} /* (30, 25, 17) {real, imag} */,
  {32'hbfa91fdf, 32'h41000a1c} /* (30, 25, 16) {real, imag} */,
  {32'h415d52d4, 32'hc04d0d0c} /* (30, 25, 15) {real, imag} */,
  {32'h40ef1345, 32'hc150d609} /* (30, 25, 14) {real, imag} */,
  {32'h41c3dec8, 32'h411c81a4} /* (30, 25, 13) {real, imag} */,
  {32'h41c7bd3c, 32'h4184f01a} /* (30, 25, 12) {real, imag} */,
  {32'h402aed1a, 32'h41792c1a} /* (30, 25, 11) {real, imag} */,
  {32'hc18eaaaa, 32'h3f82f0b3} /* (30, 25, 10) {real, imag} */,
  {32'hc1749c45, 32'hc1248ee2} /* (30, 25, 9) {real, imag} */,
  {32'hc0545190, 32'h4107e613} /* (30, 25, 8) {real, imag} */,
  {32'hc18ce2f0, 32'h4109b439} /* (30, 25, 7) {real, imag} */,
  {32'hc17f24e3, 32'hc14885ab} /* (30, 25, 6) {real, imag} */,
  {32'hc1830be9, 32'hc152d45c} /* (30, 25, 5) {real, imag} */,
  {32'h3f82ab08, 32'hc11c7f5c} /* (30, 25, 4) {real, imag} */,
  {32'h4016d064, 32'hc1cb900a} /* (30, 25, 3) {real, imag} */,
  {32'hc101f54b, 32'hc0ad37b9} /* (30, 25, 2) {real, imag} */,
  {32'hc0dd0d67, 32'h3ffa5f40} /* (30, 25, 1) {real, imag} */,
  {32'hbf85c79b, 32'hc0c5c29a} /* (30, 25, 0) {real, imag} */,
  {32'h41244f96, 32'h410fa862} /* (30, 24, 31) {real, imag} */,
  {32'h41a33780, 32'h41a63ac8} /* (30, 24, 30) {real, imag} */,
  {32'h41e96068, 32'h416ff1f9} /* (30, 24, 29) {real, imag} */,
  {32'h41f09c4e, 32'h41569d6f} /* (30, 24, 28) {real, imag} */,
  {32'h4199ca03, 32'h41738422} /* (30, 24, 27) {real, imag} */,
  {32'h41cdf2a3, 32'h41715c12} /* (30, 24, 26) {real, imag} */,
  {32'h42296144, 32'h41eeda7c} /* (30, 24, 25) {real, imag} */,
  {32'h41f268b5, 32'h42087536} /* (30, 24, 24) {real, imag} */,
  {32'h4181d9f8, 32'h41eda5ae} /* (30, 24, 23) {real, imag} */,
  {32'h41756e74, 32'h4155da1c} /* (30, 24, 22) {real, imag} */,
  {32'h413aea13, 32'hc0ed9956} /* (30, 24, 21) {real, imag} */,
  {32'hc07f1110, 32'hc1c8edc6} /* (30, 24, 20) {real, imag} */,
  {32'hbe0fcaa0, 32'hc1d730d2} /* (30, 24, 19) {real, imag} */,
  {32'h413c9193, 32'hc237f4a2} /* (30, 24, 18) {real, imag} */,
  {32'h3f5e7f5c, 32'hc257cf3c} /* (30, 24, 17) {real, imag} */,
  {32'hc1e4f81e, 32'hc204ee17} /* (30, 24, 16) {real, imag} */,
  {32'hc20f83c9, 32'hbffb3eb8} /* (30, 24, 15) {real, imag} */,
  {32'hc21caf34, 32'hc1a98fa1} /* (30, 24, 14) {real, imag} */,
  {32'hc21f159a, 32'hc2076be2} /* (30, 24, 13) {real, imag} */,
  {32'hc1f95552, 32'hc1bf3e61} /* (30, 24, 12) {real, imag} */,
  {32'hc190a510, 32'h40a506ea} /* (30, 24, 11) {real, imag} */,
  {32'hc129e590, 32'h41f96632} /* (30, 24, 10) {real, imag} */,
  {32'h41683717, 32'h41941188} /* (30, 24, 9) {real, imag} */,
  {32'h4126fd9e, 32'h41462982} /* (30, 24, 8) {real, imag} */,
  {32'h4168f13e, 32'h41e5cef0} /* (30, 24, 7) {real, imag} */,
  {32'h3fe6acb4, 32'h41f425a4} /* (30, 24, 6) {real, imag} */,
  {32'h413e0aaf, 32'h4198c8fb} /* (30, 24, 5) {real, imag} */,
  {32'h41a98e28, 32'h418bf993} /* (30, 24, 4) {real, imag} */,
  {32'h416ee558, 32'h41cbab3c} /* (30, 24, 3) {real, imag} */,
  {32'h416f0884, 32'h41bb998a} /* (30, 24, 2) {real, imag} */,
  {32'h419837b5, 32'h414ed004} /* (30, 24, 1) {real, imag} */,
  {32'h4128965c, 32'hc05f1760} /* (30, 24, 0) {real, imag} */,
  {32'hc033a3a6, 32'hc1571a6a} /* (30, 23, 31) {real, imag} */,
  {32'h3f73456c, 32'hc1563d58} /* (30, 23, 30) {real, imag} */,
  {32'h40c81f6e, 32'hc1086791} /* (30, 23, 29) {real, imag} */,
  {32'h40e6c845, 32'h40886e29} /* (30, 23, 28) {real, imag} */,
  {32'h411e7e38, 32'h40fb2ad4} /* (30, 23, 27) {real, imag} */,
  {32'h40382a9b, 32'h4164a17b} /* (30, 23, 26) {real, imag} */,
  {32'h40f67cc5, 32'h4120d806} /* (30, 23, 25) {real, imag} */,
  {32'h40f3a3e7, 32'h4170d059} /* (30, 23, 24) {real, imag} */,
  {32'h417cb9a2, 32'h409f5bfe} /* (30, 23, 23) {real, imag} */,
  {32'h40966723, 32'hc0d606d4} /* (30, 23, 22) {real, imag} */,
  {32'h40b70beb, 32'h413cda76} /* (30, 23, 21) {real, imag} */,
  {32'h414929f6, 32'h41266756} /* (30, 23, 20) {real, imag} */,
  {32'h418f9bcc, 32'h413bd6d0} /* (30, 23, 19) {real, imag} */,
  {32'h41a6e511, 32'hc11572eb} /* (30, 23, 18) {real, imag} */,
  {32'h41addc3a, 32'hc098e0d0} /* (30, 23, 17) {real, imag} */,
  {32'h419374bb, 32'hc104bda2} /* (30, 23, 16) {real, imag} */,
  {32'h419a462a, 32'hc1a624a0} /* (30, 23, 15) {real, imag} */,
  {32'h400caede, 32'hc02c421c} /* (30, 23, 14) {real, imag} */,
  {32'hc0a7757e, 32'h4063c0a6} /* (30, 23, 13) {real, imag} */,
  {32'hbf9e78a2, 32'hc0c45560} /* (30, 23, 12) {real, imag} */,
  {32'h40d73cab, 32'hc127b974} /* (30, 23, 11) {real, imag} */,
  {32'hc15758fe, 32'hc018d38e} /* (30, 23, 10) {real, imag} */,
  {32'hc20faa6d, 32'h40e39f9a} /* (30, 23, 9) {real, imag} */,
  {32'hc1ddea7f, 32'h40c064aa} /* (30, 23, 8) {real, imag} */,
  {32'hc1d84b78, 32'h419e9d59} /* (30, 23, 7) {real, imag} */,
  {32'hc19eff0e, 32'h41a05432} /* (30, 23, 6) {real, imag} */,
  {32'hbdf55000, 32'h407b15c0} /* (30, 23, 5) {real, imag} */,
  {32'h4082619a, 32'hc0d3e078} /* (30, 23, 4) {real, imag} */,
  {32'hc0d284a1, 32'hc031cd7a} /* (30, 23, 3) {real, imag} */,
  {32'h3ff65380, 32'hc0d83a88} /* (30, 23, 2) {real, imag} */,
  {32'hbeeaa5a0, 32'h409ab4c8} /* (30, 23, 1) {real, imag} */,
  {32'hc057c806, 32'h402d5984} /* (30, 23, 0) {real, imag} */,
  {32'hbf2b885e, 32'hc0fcb211} /* (30, 22, 31) {real, imag} */,
  {32'hc15749b2, 32'hc0a18f0c} /* (30, 22, 30) {real, imag} */,
  {32'hc147291a, 32'hc1162f14} /* (30, 22, 29) {real, imag} */,
  {32'hc10edaea, 32'hc019af0e} /* (30, 22, 28) {real, imag} */,
  {32'hbf6cfa90, 32'h404f6394} /* (30, 22, 27) {real, imag} */,
  {32'h3e904090, 32'h400f20f4} /* (30, 22, 26) {real, imag} */,
  {32'hc0a587d9, 32'h412f4a67} /* (30, 22, 25) {real, imag} */,
  {32'hc1520d57, 32'h3f6a8d70} /* (30, 22, 24) {real, imag} */,
  {32'h40b98960, 32'hc15011ef} /* (30, 22, 23) {real, imag} */,
  {32'h409e6ddb, 32'hc0a68118} /* (30, 22, 22) {real, imag} */,
  {32'hc124f73a, 32'h404b7e79} /* (30, 22, 21) {real, imag} */,
  {32'h40bba09b, 32'h410dad00} /* (30, 22, 20) {real, imag} */,
  {32'h40a676fb, 32'h40bca113} /* (30, 22, 19) {real, imag} */,
  {32'h4181adf2, 32'h408b985c} /* (30, 22, 18) {real, imag} */,
  {32'h41dc9df1, 32'h41807d10} /* (30, 22, 17) {real, imag} */,
  {32'h419fe7e3, 32'h4144125e} /* (30, 22, 16) {real, imag} */,
  {32'h4081a1d6, 32'hbf9674b4} /* (30, 22, 15) {real, imag} */,
  {32'h40e04442, 32'hbd918860} /* (30, 22, 14) {real, imag} */,
  {32'h4182e0c0, 32'h40c4eb98} /* (30, 22, 13) {real, imag} */,
  {32'h416a72d6, 32'h40b9d400} /* (30, 22, 12) {real, imag} */,
  {32'h4063d015, 32'hc0a520a6} /* (30, 22, 11) {real, imag} */,
  {32'hc0b87abe, 32'hc025c8b4} /* (30, 22, 10) {real, imag} */,
  {32'hc1b79bba, 32'h40093ef1} /* (30, 22, 9) {real, imag} */,
  {32'hc1e88c1e, 32'hc0e09990} /* (30, 22, 8) {real, imag} */,
  {32'hc113de9c, 32'hc14f8808} /* (30, 22, 7) {real, imag} */,
  {32'hc1b33560, 32'hc0b1667a} /* (30, 22, 6) {real, imag} */,
  {32'hc10296bc, 32'hc0a275a0} /* (30, 22, 5) {real, imag} */,
  {32'hbfc3d746, 32'hc1be7894} /* (30, 22, 4) {real, imag} */,
  {32'h4035e9ec, 32'hc10a9d4c} /* (30, 22, 3) {real, imag} */,
  {32'hbffe33f0, 32'h40218988} /* (30, 22, 2) {real, imag} */,
  {32'hc0220f1c, 32'hc13c9b59} /* (30, 22, 1) {real, imag} */,
  {32'hbfc7fdbe, 32'hc158743e} /* (30, 22, 0) {real, imag} */,
  {32'h409bd892, 32'h3fe22034} /* (30, 21, 31) {real, imag} */,
  {32'hbf8015d8, 32'h40a3a006} /* (30, 21, 30) {real, imag} */,
  {32'h40c53711, 32'h4132dbc6} /* (30, 21, 29) {real, imag} */,
  {32'h41b519b3, 32'h412dd85a} /* (30, 21, 28) {real, imag} */,
  {32'h41e4ef27, 32'h4156f2f0} /* (30, 21, 27) {real, imag} */,
  {32'h41712d14, 32'h41860b78} /* (30, 21, 26) {real, imag} */,
  {32'h4192bf47, 32'h41614b8e} /* (30, 21, 25) {real, imag} */,
  {32'h41b35199, 32'h415dfecc} /* (30, 21, 24) {real, imag} */,
  {32'h41b37b19, 32'h417de01f} /* (30, 21, 23) {real, imag} */,
  {32'h418ecec0, 32'h41594608} /* (30, 21, 22) {real, imag} */,
  {32'h416c2964, 32'h40143684} /* (30, 21, 21) {real, imag} */,
  {32'h410e4286, 32'h409859f6} /* (30, 21, 20) {real, imag} */,
  {32'h3f9e7498, 32'h411b7f2e} /* (30, 21, 19) {real, imag} */,
  {32'h3f20d3c8, 32'h40aded6e} /* (30, 21, 18) {real, imag} */,
  {32'hc0e19390, 32'h3f52bc90} /* (30, 21, 17) {real, imag} */,
  {32'hc10e7472, 32'h3fa089f0} /* (30, 21, 16) {real, imag} */,
  {32'hc18064b9, 32'h411daf5d} /* (30, 21, 15) {real, imag} */,
  {32'hc1d46534, 32'h40b65659} /* (30, 21, 14) {real, imag} */,
  {32'hc16fa462, 32'hbfc8d7fc} /* (30, 21, 13) {real, imag} */,
  {32'hc1584664, 32'h40ce431c} /* (30, 21, 12) {real, imag} */,
  {32'hc09a582c, 32'hc105e1a4} /* (30, 21, 11) {real, imag} */,
  {32'h4124e645, 32'hc0b14da0} /* (30, 21, 10) {real, imag} */,
  {32'h4128bf20, 32'h3e9e3260} /* (30, 21, 9) {real, imag} */,
  {32'hc001c986, 32'h4078be10} /* (30, 21, 8) {real, imag} */,
  {32'h41b80f54, 32'h410e9f8e} /* (30, 21, 7) {real, imag} */,
  {32'h420274e2, 32'h414c46a6} /* (30, 21, 6) {real, imag} */,
  {32'h41a2f5d6, 32'h4181f654} /* (30, 21, 5) {real, imag} */,
  {32'h41eefaab, 32'h41738e4f} /* (30, 21, 4) {real, imag} */,
  {32'h41b41f37, 32'h4129bd50} /* (30, 21, 3) {real, imag} */,
  {32'h418a33b3, 32'h415489ee} /* (30, 21, 2) {real, imag} */,
  {32'h41379a6b, 32'h414342ef} /* (30, 21, 1) {real, imag} */,
  {32'h4109ad12, 32'h40d77872} /* (30, 21, 0) {real, imag} */,
  {32'hbf50629d, 32'h3f200698} /* (30, 20, 31) {real, imag} */,
  {32'hc08bfcb1, 32'hc11cd82f} /* (30, 20, 30) {real, imag} */,
  {32'h3fef26c4, 32'hc15d922a} /* (30, 20, 29) {real, imag} */,
  {32'h40f871f5, 32'hc0c1ce7f} /* (30, 20, 28) {real, imag} */,
  {32'hbf5af5d6, 32'h403a5bb0} /* (30, 20, 27) {real, imag} */,
  {32'hc0760445, 32'h3f7d12f0} /* (30, 20, 26) {real, imag} */,
  {32'hc0b3c426, 32'h3f98f81e} /* (30, 20, 25) {real, imag} */,
  {32'hc137899b, 32'h40f4ed3e} /* (30, 20, 24) {real, imag} */,
  {32'hc13c3978, 32'h4062f90c} /* (30, 20, 23) {real, imag} */,
  {32'hbf993c30, 32'h40518c38} /* (30, 20, 22) {real, imag} */,
  {32'h415c1bbe, 32'h410069e0} /* (30, 20, 21) {real, imag} */,
  {32'h415352b8, 32'hbfde6a68} /* (30, 20, 20) {real, imag} */,
  {32'h3fe489ea, 32'hbf827808} /* (30, 20, 19) {real, imag} */,
  {32'hc00ab0b8, 32'hc002a628} /* (30, 20, 18) {real, imag} */,
  {32'h40e31897, 32'h40c7d475} /* (30, 20, 17) {real, imag} */,
  {32'h408a7a42, 32'h408ac372} /* (30, 20, 16) {real, imag} */,
  {32'hc027f462, 32'h403203aa} /* (30, 20, 15) {real, imag} */,
  {32'hc106767a, 32'h3fc8f674} /* (30, 20, 14) {real, imag} */,
  {32'hc183b665, 32'hc006460d} /* (30, 20, 13) {real, imag} */,
  {32'hc098bb58, 32'h40061d18} /* (30, 20, 12) {real, imag} */,
  {32'hc0c3486a, 32'h40873a20} /* (30, 20, 11) {real, imag} */,
  {32'hc04b8896, 32'hc0860784} /* (30, 20, 10) {real, imag} */,
  {32'h40c6267c, 32'hc010e47c} /* (30, 20, 9) {real, imag} */,
  {32'h411b5d34, 32'hbf1314f0} /* (30, 20, 8) {real, imag} */,
  {32'h3fd7fca8, 32'hc0409164} /* (30, 20, 7) {real, imag} */,
  {32'hc04a91d6, 32'hc06d06e4} /* (30, 20, 6) {real, imag} */,
  {32'h3f955a6c, 32'h3fb91744} /* (30, 20, 5) {real, imag} */,
  {32'hbef9be98, 32'h3f85a9d0} /* (30, 20, 4) {real, imag} */,
  {32'hc04a2efe, 32'hc0d0d57a} /* (30, 20, 3) {real, imag} */,
  {32'hc0a00f79, 32'hc04fd6a4} /* (30, 20, 2) {real, imag} */,
  {32'h3f9100b4, 32'hbf8634f0} /* (30, 20, 1) {real, imag} */,
  {32'hbdd05220, 32'h40426da6} /* (30, 20, 0) {real, imag} */,
  {32'hc029338b, 32'hbf118758} /* (30, 19, 31) {real, imag} */,
  {32'hc0657c3c, 32'hc09b04e2} /* (30, 19, 30) {real, imag} */,
  {32'hbff36450, 32'hc0969521} /* (30, 19, 29) {real, imag} */,
  {32'hbf980388, 32'hc0afa7f6} /* (30, 19, 28) {real, imag} */,
  {32'h402575f2, 32'hc0873838} /* (30, 19, 27) {real, imag} */,
  {32'h3daf6d80, 32'hc01d6c4a} /* (30, 19, 26) {real, imag} */,
  {32'hbff7b0c8, 32'h3c370c00} /* (30, 19, 25) {real, imag} */,
  {32'hbfacb6ea, 32'hbedf5300} /* (30, 19, 24) {real, imag} */,
  {32'hbf5f53e0, 32'hc0aa0d63} /* (30, 19, 23) {real, imag} */,
  {32'h40fe9c8e, 32'hc06ba356} /* (30, 19, 22) {real, imag} */,
  {32'h3fa45cb4, 32'h3fa1d220} /* (30, 19, 21) {real, imag} */,
  {32'hbfd9319a, 32'h405fa40b} /* (30, 19, 20) {real, imag} */,
  {32'hbf906b0c, 32'h40076774} /* (30, 19, 19) {real, imag} */,
  {32'h40d82b2b, 32'hc09b4006} /* (30, 19, 18) {real, imag} */,
  {32'h4122f9d6, 32'hc058aca0} /* (30, 19, 17) {real, imag} */,
  {32'h408427fc, 32'hbd6af680} /* (30, 19, 16) {real, imag} */,
  {32'hc06f3f60, 32'hc067d1b4} /* (30, 19, 15) {real, imag} */,
  {32'hc01a4842, 32'hc0c2cefd} /* (30, 19, 14) {real, imag} */,
  {32'h3eebe2f0, 32'hc0f23945} /* (30, 19, 13) {real, imag} */,
  {32'hbf0a536c, 32'hc0eb3252} /* (30, 19, 12) {real, imag} */,
  {32'hbf281478, 32'hbf945d8c} /* (30, 19, 11) {real, imag} */,
  {32'hc090aa76, 32'h3fe51424} /* (30, 19, 10) {real, imag} */,
  {32'h409f3c49, 32'hbf940b28} /* (30, 19, 9) {real, imag} */,
  {32'h3d8757c0, 32'h3fe686ac} /* (30, 19, 8) {real, imag} */,
  {32'hc0fa1238, 32'h403f30d0} /* (30, 19, 7) {real, imag} */,
  {32'hc03afe98, 32'h40805794} /* (30, 19, 6) {real, imag} */,
  {32'h3e0619c0, 32'h3f0f1f4c} /* (30, 19, 5) {real, imag} */,
  {32'h40b33c49, 32'hbf087fc0} /* (30, 19, 4) {real, imag} */,
  {32'h4088e576, 32'h407c2970} /* (30, 19, 3) {real, imag} */,
  {32'h404393fa, 32'h40432ce6} /* (30, 19, 2) {real, imag} */,
  {32'hbfdc4724, 32'h3fc682a4} /* (30, 19, 1) {real, imag} */,
  {32'hc031675d, 32'hbed9db30} /* (30, 19, 0) {real, imag} */,
  {32'hbf99f014, 32'h3fadb404} /* (30, 18, 31) {real, imag} */,
  {32'h402fd5f8, 32'hbf29158c} /* (30, 18, 30) {real, imag} */,
  {32'h407c28fe, 32'h40351d83} /* (30, 18, 29) {real, imag} */,
  {32'h41153263, 32'hc0032b10} /* (30, 18, 28) {real, imag} */,
  {32'h4155b180, 32'hc0673f0c} /* (30, 18, 27) {real, imag} */,
  {32'h4173aaeb, 32'hbfc0add8} /* (30, 18, 26) {real, imag} */,
  {32'h414f6554, 32'hbec31540} /* (30, 18, 25) {real, imag} */,
  {32'h416e7c77, 32'hbe374730} /* (30, 18, 24) {real, imag} */,
  {32'h411b04ff, 32'h40beabf6} /* (30, 18, 23) {real, imag} */,
  {32'h40b1cde2, 32'h40a9f263} /* (30, 18, 22) {real, imag} */,
  {32'h3f754d88, 32'hbf97b5a8} /* (30, 18, 21) {real, imag} */,
  {32'hc0861b48, 32'hc1163874} /* (30, 18, 20) {real, imag} */,
  {32'hc0cc1324, 32'hc10e48c4} /* (30, 18, 19) {real, imag} */,
  {32'hbe820a80, 32'hbf37c3c0} /* (30, 18, 18) {real, imag} */,
  {32'hbe98a480, 32'h3fa53df0} /* (30, 18, 17) {real, imag} */,
  {32'hc0279060, 32'hc064339c} /* (30, 18, 16) {real, imag} */,
  {32'hc09e5f84, 32'hc0f24b82} /* (30, 18, 15) {real, imag} */,
  {32'hc1654841, 32'hc0c04d5e} /* (30, 18, 14) {real, imag} */,
  {32'hc188f502, 32'hbfdc0d9c} /* (30, 18, 13) {real, imag} */,
  {32'hc184971c, 32'h403d8480} /* (30, 18, 12) {real, imag} */,
  {32'hc083608a, 32'h405d5e17} /* (30, 18, 11) {real, imag} */,
  {32'h4102cecc, 32'hc0a5401f} /* (30, 18, 10) {real, imag} */,
  {32'h414ad868, 32'h3fab4d82} /* (30, 18, 9) {real, imag} */,
  {32'h411676fe, 32'h40a51732} /* (30, 18, 8) {real, imag} */,
  {32'h40837094, 32'h409d7dba} /* (30, 18, 7) {real, imag} */,
  {32'h40c24f56, 32'h40a3c8e2} /* (30, 18, 6) {real, imag} */,
  {32'h41145dba, 32'hc054353e} /* (30, 18, 5) {real, imag} */,
  {32'h402846e9, 32'hc0aa4e80} /* (30, 18, 4) {real, imag} */,
  {32'h4048ad14, 32'hbfeac2b8} /* (30, 18, 3) {real, imag} */,
  {32'h40779178, 32'h3ddb4960} /* (30, 18, 2) {real, imag} */,
  {32'h40ea3d08, 32'h40823f5e} /* (30, 18, 1) {real, imag} */,
  {32'h41127670, 32'h4090cdd0} /* (30, 18, 0) {real, imag} */,
  {32'hc0e16434, 32'h3fea6c05} /* (30, 17, 31) {real, imag} */,
  {32'hc083b4f8, 32'h409ad8a2} /* (30, 17, 30) {real, imag} */,
  {32'h3fef65c4, 32'h40b3b980} /* (30, 17, 29) {real, imag} */,
  {32'hc0eb8a0e, 32'h406e8d78} /* (30, 17, 28) {real, imag} */,
  {32'hc140d9a6, 32'h40992d33} /* (30, 17, 27) {real, imag} */,
  {32'hc0b1025a, 32'h402e5d72} /* (30, 17, 26) {real, imag} */,
  {32'hc044bb60, 32'hc0443870} /* (30, 17, 25) {real, imag} */,
  {32'h406e8cb4, 32'hc09a5580} /* (30, 17, 24) {real, imag} */,
  {32'h4019cce8, 32'hc038ee08} /* (30, 17, 23) {real, imag} */,
  {32'hc0ab1e7c, 32'hbfb640b8} /* (30, 17, 22) {real, imag} */,
  {32'hc10f2297, 32'hc0b81480} /* (30, 17, 21) {real, imag} */,
  {32'hc02a5fb4, 32'hc105778c} /* (30, 17, 20) {real, imag} */,
  {32'h40e7117f, 32'hc0ec7e06} /* (30, 17, 19) {real, imag} */,
  {32'h40f49268, 32'hc0589e78} /* (30, 17, 18) {real, imag} */,
  {32'h40285e1e, 32'h404d81f6} /* (30, 17, 17) {real, imag} */,
  {32'hc03850d0, 32'h402c93b4} /* (30, 17, 16) {real, imag} */,
  {32'h3ffdac78, 32'h40047590} /* (30, 17, 15) {real, imag} */,
  {32'h40ff3766, 32'h4098185e} /* (30, 17, 14) {real, imag} */,
  {32'h40c8af64, 32'h40cc2c4f} /* (30, 17, 13) {real, imag} */,
  {32'hc0036be4, 32'hbe972d78} /* (30, 17, 12) {real, imag} */,
  {32'hbf4f700a, 32'hc107b344} /* (30, 17, 11) {real, imag} */,
  {32'hc01ae6ae, 32'hc0b324a9} /* (30, 17, 10) {real, imag} */,
  {32'hbfd607a8, 32'hc0940554} /* (30, 17, 9) {real, imag} */,
  {32'h3f79daa0, 32'h3edf8380} /* (30, 17, 8) {real, imag} */,
  {32'hc04ceb10, 32'h40041af8} /* (30, 17, 7) {real, imag} */,
  {32'hc1015a2b, 32'h401fa4d4} /* (30, 17, 6) {real, imag} */,
  {32'hc0e3bfae, 32'h40cff40e} /* (30, 17, 5) {real, imag} */,
  {32'hc03c03f4, 32'h40c92146} /* (30, 17, 4) {real, imag} */,
  {32'h3e437d20, 32'h4014a328} /* (30, 17, 3) {real, imag} */,
  {32'hbf99d5d8, 32'h40b39dde} /* (30, 17, 2) {real, imag} */,
  {32'h3f0c52a0, 32'h408ab556} /* (30, 17, 1) {real, imag} */,
  {32'h3f463080, 32'h3fdf29d5} /* (30, 17, 0) {real, imag} */,
  {32'hc04ae9d0, 32'h403092b0} /* (30, 16, 31) {real, imag} */,
  {32'hc02783b0, 32'h40c3b3c0} /* (30, 16, 30) {real, imag} */,
  {32'hbfe220b8, 32'h402c3b40} /* (30, 16, 29) {real, imag} */,
  {32'hbe3e6c80, 32'hbfa4cc80} /* (30, 16, 28) {real, imag} */,
  {32'hbff2fb30, 32'h3fa73400} /* (30, 16, 27) {real, imag} */,
  {32'hc05e43ac, 32'hbfc9bb00} /* (30, 16, 26) {real, imag} */,
  {32'h3f20ea78, 32'h4066b5c0} /* (30, 16, 25) {real, imag} */,
  {32'h401b90a8, 32'h40a8d770} /* (30, 16, 24) {real, imag} */,
  {32'h40bf2d08, 32'hc008b260} /* (30, 16, 23) {real, imag} */,
  {32'h3e88e440, 32'h402aa180} /* (30, 16, 22) {real, imag} */,
  {32'h3fa340d8, 32'h40ba0228} /* (30, 16, 21) {real, imag} */,
  {32'h4037fcdf, 32'h3fa54340} /* (30, 16, 20) {real, imag} */,
  {32'hbdef0600, 32'hc00ad544} /* (30, 16, 19) {real, imag} */,
  {32'hbf993fc0, 32'h3e3406c0} /* (30, 16, 18) {real, imag} */,
  {32'hbfcbe260, 32'hbf83c818} /* (30, 16, 17) {real, imag} */,
  {32'h3fcd3230, 32'hbe46c500} /* (30, 16, 16) {real, imag} */,
  {32'hbfe2194c, 32'h4013c760} /* (30, 16, 15) {real, imag} */,
  {32'hbd93c580, 32'h3c73e000} /* (30, 16, 14) {real, imag} */,
  {32'hc03965d0, 32'h3cf85000} /* (30, 16, 13) {real, imag} */,
  {32'hc0a4b6d0, 32'h3fcf7100} /* (30, 16, 12) {real, imag} */,
  {32'hc04e3640, 32'hc02a4000} /* (30, 16, 11) {real, imag} */,
  {32'hc05ed310, 32'hbfd67380} /* (30, 16, 10) {real, imag} */,
  {32'hc083b256, 32'hc05a4404} /* (30, 16, 9) {real, imag} */,
  {32'h3ed5ba20, 32'hc0ad9082} /* (30, 16, 8) {real, imag} */,
  {32'h409be370, 32'hc0cc8d80} /* (30, 16, 7) {real, imag} */,
  {32'h3f8da4e2, 32'hc03c9a16} /* (30, 16, 6) {real, imag} */,
  {32'hc10276bc, 32'h4112b8b0} /* (30, 16, 5) {real, imag} */,
  {32'hc0b50fa4, 32'h40b4f6c0} /* (30, 16, 4) {real, imag} */,
  {32'hc01e655f, 32'h4080bb00} /* (30, 16, 3) {real, imag} */,
  {32'hc0ffeca8, 32'hbe457000} /* (30, 16, 2) {real, imag} */,
  {32'hc0134060, 32'hbf968de0} /* (30, 16, 1) {real, imag} */,
  {32'hc01ddb60, 32'hc07b8020} /* (30, 16, 0) {real, imag} */,
  {32'h40c43ab4, 32'h3e54d3d8} /* (30, 15, 31) {real, imag} */,
  {32'h403801e0, 32'h4049ccfc} /* (30, 15, 30) {real, imag} */,
  {32'h40d947ff, 32'h407890ff} /* (30, 15, 29) {real, imag} */,
  {32'h408ea4d6, 32'h3e8fbc40} /* (30, 15, 28) {real, imag} */,
  {32'hbd438980, 32'h406e3b1a} /* (30, 15, 27) {real, imag} */,
  {32'h40912772, 32'h40882ac7} /* (30, 15, 26) {real, imag} */,
  {32'h40aa5fb8, 32'h40a50f78} /* (30, 15, 25) {real, imag} */,
  {32'h4066d0bc, 32'h400a64c0} /* (30, 15, 24) {real, imag} */,
  {32'h405414a8, 32'h4011c688} /* (30, 15, 23) {real, imag} */,
  {32'h40488558, 32'h40aa50ce} /* (30, 15, 22) {real, imag} */,
  {32'h40856a26, 32'hbf65e600} /* (30, 15, 21) {real, imag} */,
  {32'h3ed6b460, 32'h3ec0e680} /* (30, 15, 20) {real, imag} */,
  {32'hc06060a2, 32'h40814496} /* (30, 15, 19) {real, imag} */,
  {32'hc13e3204, 32'h40c838fc} /* (30, 15, 18) {real, imag} */,
  {32'hc147af68, 32'hbeebb5b0} /* (30, 15, 17) {real, imag} */,
  {32'hc06543d0, 32'h40bb2906} /* (30, 15, 16) {real, imag} */,
  {32'h3ff70be8, 32'hbeee1484} /* (30, 15, 15) {real, imag} */,
  {32'hbfd18f58, 32'hc08fb61e} /* (30, 15, 14) {real, imag} */,
  {32'hc0ba6da4, 32'hc042f81e} /* (30, 15, 13) {real, imag} */,
  {32'hc04342bc, 32'hbf6e1644} /* (30, 15, 12) {real, imag} */,
  {32'hc044670e, 32'h406603d0} /* (30, 15, 11) {real, imag} */,
  {32'h410c10cc, 32'h401011c6} /* (30, 15, 10) {real, imag} */,
  {32'h40af5216, 32'hc043d578} /* (30, 15, 9) {real, imag} */,
  {32'h40d8f8a4, 32'hbffbb260} /* (30, 15, 8) {real, imag} */,
  {32'h413b865c, 32'h3f338320} /* (30, 15, 7) {real, imag} */,
  {32'h4180085b, 32'h3f087330} /* (30, 15, 6) {real, imag} */,
  {32'h414ae865, 32'hbf5ebf74} /* (30, 15, 5) {real, imag} */,
  {32'h40cb314a, 32'h40112df4} /* (30, 15, 4) {real, imag} */,
  {32'h3fc3421c, 32'h3fc07e30} /* (30, 15, 3) {real, imag} */,
  {32'hc00387b4, 32'h4005e144} /* (30, 15, 2) {real, imag} */,
  {32'h408b6c24, 32'hbefc8160} /* (30, 15, 1) {real, imag} */,
  {32'h40bb5988, 32'hbf8c6315} /* (30, 15, 0) {real, imag} */,
  {32'hc0ce3c73, 32'h3e836bf0} /* (30, 14, 31) {real, imag} */,
  {32'hc1117042, 32'h3fba28c6} /* (30, 14, 30) {real, imag} */,
  {32'hc1200850, 32'hc02ceec3} /* (30, 14, 29) {real, imag} */,
  {32'hc10b6f01, 32'hc0bca8f8} /* (30, 14, 28) {real, imag} */,
  {32'hc0a29d50, 32'h3fe04118} /* (30, 14, 27) {real, imag} */,
  {32'hc0a723b6, 32'hbf284650} /* (30, 14, 26) {real, imag} */,
  {32'hc0fe18ec, 32'h40161a28} /* (30, 14, 25) {real, imag} */,
  {32'hc140ac6d, 32'h40b1409a} /* (30, 14, 24) {real, imag} */,
  {32'hc0c14a82, 32'hbfd8fdd8} /* (30, 14, 23) {real, imag} */,
  {32'hc147c04f, 32'hc033ad86} /* (30, 14, 22) {real, imag} */,
  {32'hc0ded0ff, 32'hc1016ca3} /* (30, 14, 21) {real, imag} */,
  {32'hc05ca230, 32'hc12d4b8c} /* (30, 14, 20) {real, imag} */,
  {32'h3f9bffb0, 32'hc03e1830} /* (30, 14, 19) {real, imag} */,
  {32'h3f65f1c0, 32'hc0009f90} /* (30, 14, 18) {real, imag} */,
  {32'hbe2b9500, 32'hbfef7770} /* (30, 14, 17) {real, imag} */,
  {32'h40147940, 32'hc0a16672} /* (30, 14, 16) {real, imag} */,
  {32'h4031fb68, 32'hc01fe4bc} /* (30, 14, 15) {real, imag} */,
  {32'h3f876b98, 32'hc0343e05} /* (30, 14, 14) {real, imag} */,
  {32'h40a71f5a, 32'hc125458c} /* (30, 14, 13) {real, imag} */,
  {32'h417aff28, 32'hc0f03d00} /* (30, 14, 12) {real, imag} */,
  {32'h419f4e04, 32'hc0294f57} /* (30, 14, 11) {real, imag} */,
  {32'h410b63bc, 32'h402e9bbe} /* (30, 14, 10) {real, imag} */,
  {32'hbfba1680, 32'h410318a0} /* (30, 14, 9) {real, imag} */,
  {32'hc05f5b68, 32'h40e385ce} /* (30, 14, 8) {real, imag} */,
  {32'hc0e8ccb4, 32'h4075ea0c} /* (30, 14, 7) {real, imag} */,
  {32'hc117eed5, 32'h3f5ebcf0} /* (30, 14, 6) {real, imag} */,
  {32'hc03058ba, 32'hc0c8ad21} /* (30, 14, 5) {real, imag} */,
  {32'hc0064271, 32'hc1311420} /* (30, 14, 4) {real, imag} */,
  {32'hc0ba0f6e, 32'hc06c3aa4} /* (30, 14, 3) {real, imag} */,
  {32'hc10cee0a, 32'h41017d2d} /* (30, 14, 2) {real, imag} */,
  {32'hc09b3c88, 32'h40d229e2} /* (30, 14, 1) {real, imag} */,
  {32'hbfef75e4, 32'h3ed69c00} /* (30, 14, 0) {real, imag} */,
  {32'h40d1ade6, 32'hc0dab16d} /* (30, 13, 31) {real, imag} */,
  {32'h41757eeb, 32'hc0b7f4a6} /* (30, 13, 30) {real, imag} */,
  {32'h40be6ada, 32'h3f9ef274} /* (30, 13, 29) {real, imag} */,
  {32'h3eba0e20, 32'hbea91160} /* (30, 13, 28) {real, imag} */,
  {32'hc12930a4, 32'hc0a64220} /* (30, 13, 27) {real, imag} */,
  {32'hbeab13e0, 32'hc0aae245} /* (30, 13, 26) {real, imag} */,
  {32'h4138a5f3, 32'hc0c104be} /* (30, 13, 25) {real, imag} */,
  {32'h4111c2f3, 32'hc0181f88} /* (30, 13, 24) {real, imag} */,
  {32'hc0b88444, 32'hc06b34bb} /* (30, 13, 23) {real, imag} */,
  {32'hc11905a5, 32'hc073823a} /* (30, 13, 22) {real, imag} */,
  {32'hc0ca6e51, 32'h400d89b0} /* (30, 13, 21) {real, imag} */,
  {32'hc094e706, 32'h40df0822} /* (30, 13, 20) {real, imag} */,
  {32'h3f0590e8, 32'h3fe3b9f8} /* (30, 13, 19) {real, imag} */,
  {32'h3f57e558, 32'h4088faa2} /* (30, 13, 18) {real, imag} */,
  {32'hc038ac6a, 32'h3fa51060} /* (30, 13, 17) {real, imag} */,
  {32'hbe47b080, 32'hbf032128} /* (30, 13, 16) {real, imag} */,
  {32'h4075b390, 32'h40555070} /* (30, 13, 15) {real, imag} */,
  {32'h40c7eb7f, 32'hbf510c78} /* (30, 13, 14) {real, imag} */,
  {32'hc00cda4a, 32'h40cd946b} /* (30, 13, 13) {real, imag} */,
  {32'hc021ac19, 32'h4140ec73} /* (30, 13, 12) {real, imag} */,
  {32'h3f997d84, 32'h41223d2e} /* (30, 13, 11) {real, imag} */,
  {32'h411a1095, 32'hbfc8352c} /* (30, 13, 10) {real, imag} */,
  {32'h40b63119, 32'hc0b0f04e} /* (30, 13, 9) {real, imag} */,
  {32'h402cf81e, 32'hc012604a} /* (30, 13, 8) {real, imag} */,
  {32'h40b8d2a8, 32'hbf668ca0} /* (30, 13, 7) {real, imag} */,
  {32'h40ffc574, 32'hbf202c00} /* (30, 13, 6) {real, imag} */,
  {32'h40be9956, 32'hbfa9e596} /* (30, 13, 5) {real, imag} */,
  {32'h4055961a, 32'hbf4ab540} /* (30, 13, 4) {real, imag} */,
  {32'h40f4f646, 32'h3de4a500} /* (30, 13, 3) {real, imag} */,
  {32'h403e3b6a, 32'h3feadc04} /* (30, 13, 2) {real, imag} */,
  {32'hc046cbce, 32'hc1057ac4} /* (30, 13, 1) {real, imag} */,
  {32'h3f40f35c, 32'hc14424dc} /* (30, 13, 0) {real, imag} */,
  {32'hbfb92906, 32'hc098043d} /* (30, 12, 31) {real, imag} */,
  {32'hbfc6b370, 32'h3d4ec100} /* (30, 12, 30) {real, imag} */,
  {32'hbfeee82c, 32'h40ca8d60} /* (30, 12, 29) {real, imag} */,
  {32'h3f8284ec, 32'h408cc877} /* (30, 12, 28) {real, imag} */,
  {32'h404a9c8a, 32'h3f9d5ee0} /* (30, 12, 27) {real, imag} */,
  {32'hc0044245, 32'h3f9c1b88} /* (30, 12, 26) {real, imag} */,
  {32'hc056eea8, 32'h3f746a84} /* (30, 12, 25) {real, imag} */,
  {32'hbe522000, 32'h409dae62} /* (30, 12, 24) {real, imag} */,
  {32'hc0353f22, 32'hc013ca5c} /* (30, 12, 23) {real, imag} */,
  {32'hc0b02bd2, 32'hc0976b0c} /* (30, 12, 22) {real, imag} */,
  {32'hbf9ca4dc, 32'hc019ee06} /* (30, 12, 21) {real, imag} */,
  {32'h4099dfc0, 32'hc14d079b} /* (30, 12, 20) {real, imag} */,
  {32'hc100bb23, 32'hc0bd19f6} /* (30, 12, 19) {real, imag} */,
  {32'hc12b9496, 32'h400424e8} /* (30, 12, 18) {real, imag} */,
  {32'hc0b54759, 32'hc1191fca} /* (30, 12, 17) {real, imag} */,
  {32'hc0b0882e, 32'hc1101479} /* (30, 12, 16) {real, imag} */,
  {32'hc1208824, 32'hc0926b85} /* (30, 12, 15) {real, imag} */,
  {32'hc0ad9069, 32'h40a7b783} /* (30, 12, 14) {real, imag} */,
  {32'h4049ca48, 32'h3fc8607a} /* (30, 12, 13) {real, imag} */,
  {32'h3f8e7e38, 32'hbfed64f0} /* (30, 12, 12) {real, imag} */,
  {32'hc0bee590, 32'h408f2e3c} /* (30, 12, 11) {real, imag} */,
  {32'hc0cbbafb, 32'hc104bdc6} /* (30, 12, 10) {real, imag} */,
  {32'hbee37cc0, 32'hc12ad5c5} /* (30, 12, 9) {real, imag} */,
  {32'hc04911a0, 32'hc0419104} /* (30, 12, 8) {real, imag} */,
  {32'hc079f01c, 32'h4006d344} /* (30, 12, 7) {real, imag} */,
  {32'hc02c0b76, 32'hc1522c87} /* (30, 12, 6) {real, imag} */,
  {32'hc0abff1d, 32'hc0c5ff69} /* (30, 12, 5) {real, imag} */,
  {32'hbf9a7b66, 32'h3fc9dc70} /* (30, 12, 4) {real, imag} */,
  {32'h40bb7f99, 32'hbff2f748} /* (30, 12, 3) {real, imag} */,
  {32'h40a8b263, 32'hc052bfcc} /* (30, 12, 2) {real, imag} */,
  {32'h4102e1d0, 32'hc0df87c4} /* (30, 12, 1) {real, imag} */,
  {32'hbf29ec2c, 32'hbfb4c8ac} /* (30, 12, 0) {real, imag} */,
  {32'hc120d5cb, 32'h411a1a7e} /* (30, 11, 31) {real, imag} */,
  {32'hc183a51e, 32'h41afee3c} /* (30, 11, 30) {real, imag} */,
  {32'hc180b612, 32'h418a65c5} /* (30, 11, 29) {real, imag} */,
  {32'hc1924c9b, 32'h419a4cdb} /* (30, 11, 28) {real, imag} */,
  {32'hc13d0e7e, 32'h41b7edf2} /* (30, 11, 27) {real, imag} */,
  {32'hc0988347, 32'h41545ee6} /* (30, 11, 26) {real, imag} */,
  {32'hc12fda58, 32'h411e142a} /* (30, 11, 25) {real, imag} */,
  {32'hc18596ef, 32'h4106b2d4} /* (30, 11, 24) {real, imag} */,
  {32'hc0f71afc, 32'h410b4bd1} /* (30, 11, 23) {real, imag} */,
  {32'hc18adea4, 32'h415112a8} /* (30, 11, 22) {real, imag} */,
  {32'hc1404244, 32'h41829d58} /* (30, 11, 21) {real, imag} */,
  {32'h415f7acc, 32'hbea509e8} /* (30, 11, 20) {real, imag} */,
  {32'h416ef3c5, 32'hc15cc96e} /* (30, 11, 19) {real, imag} */,
  {32'h40d8cab5, 32'hc0fbe5ee} /* (30, 11, 18) {real, imag} */,
  {32'h41b18f3a, 32'h3e00f0c0} /* (30, 11, 17) {real, imag} */,
  {32'h41919391, 32'h41069c2e} /* (30, 11, 16) {real, imag} */,
  {32'h418794f3, 32'h3eac02e0} /* (30, 11, 15) {real, imag} */,
  {32'h4121fc70, 32'hc05dea82} /* (30, 11, 14) {real, imag} */,
  {32'h412df4fe, 32'hc0b20561} /* (30, 11, 13) {real, imag} */,
  {32'h41137296, 32'hc1574c2a} /* (30, 11, 12) {real, imag} */,
  {32'h410472b3, 32'hc0f5d728} /* (30, 11, 11) {real, imag} */,
  {32'hc0a1739e, 32'h40780538} /* (30, 11, 10) {real, imag} */,
  {32'hc126070e, 32'hc0670dac} /* (30, 11, 9) {real, imag} */,
  {32'hc1362d78, 32'h407c5358} /* (30, 11, 8) {real, imag} */,
  {32'h40327eec, 32'h412680d6} /* (30, 11, 7) {real, imag} */,
  {32'hc0a5accc, 32'h41b67c9b} /* (30, 11, 6) {real, imag} */,
  {32'hc1820ff0, 32'h41e4a0ca} /* (30, 11, 5) {real, imag} */,
  {32'hc15375aa, 32'h41a37ae2} /* (30, 11, 4) {real, imag} */,
  {32'hc190e4d7, 32'h412b8d2c} /* (30, 11, 3) {real, imag} */,
  {32'hc1a7aad5, 32'h41b68fb1} /* (30, 11, 2) {real, imag} */,
  {32'hc0afb8c2, 32'h41607589} /* (30, 11, 1) {real, imag} */,
  {32'hbfd8cec8, 32'h3f3a4cd0} /* (30, 11, 0) {real, imag} */,
  {32'h3fda0639, 32'hbfe962cc} /* (30, 10, 31) {real, imag} */,
  {32'h406e5132, 32'hc01ffae1} /* (30, 10, 30) {real, imag} */,
  {32'h41460df4, 32'h408dd9f9} /* (30, 10, 29) {real, imag} */,
  {32'h41ab3899, 32'h405f67f6} /* (30, 10, 28) {real, imag} */,
  {32'h40d4ede0, 32'h4163cedf} /* (30, 10, 27) {real, imag} */,
  {32'h3f9fe3c4, 32'h410d8ec1} /* (30, 10, 26) {real, imag} */,
  {32'h3f99c0dc, 32'hc0dc504a} /* (30, 10, 25) {real, imag} */,
  {32'hc12f382b, 32'h408c0632} /* (30, 10, 24) {real, imag} */,
  {32'hbf86e5c0, 32'hc09d2742} /* (30, 10, 23) {real, imag} */,
  {32'h4025a2b6, 32'hc116684a} /* (30, 10, 22) {real, imag} */,
  {32'hc15de468, 32'hc0411c79} /* (30, 10, 21) {real, imag} */,
  {32'hc1935ce5, 32'h40d1cff8} /* (30, 10, 20) {real, imag} */,
  {32'hc17c7ede, 32'h410e1588} /* (30, 10, 19) {real, imag} */,
  {32'hc165083b, 32'h413aa3f2} /* (30, 10, 18) {real, imag} */,
  {32'hc18a062f, 32'h40e2208c} /* (30, 10, 17) {real, imag} */,
  {32'hc17a7d4a, 32'h411113ba} /* (30, 10, 16) {real, imag} */,
  {32'hc0bf2872, 32'hc0088366} /* (30, 10, 15) {real, imag} */,
  {32'hbde08720, 32'hc001c065} /* (30, 10, 14) {real, imag} */,
  {32'h408b8bc2, 32'h40adc44c} /* (30, 10, 13) {real, imag} */,
  {32'h4111f5da, 32'h408cb624} /* (30, 10, 12) {real, imag} */,
  {32'h411f27ff, 32'hc09af236} /* (30, 10, 11) {real, imag} */,
  {32'h418bff60, 32'hc0d9e102} /* (30, 10, 10) {real, imag} */,
  {32'h4175b47c, 32'hc0770681} /* (30, 10, 9) {real, imag} */,
  {32'h41924a6a, 32'hc05fef68} /* (30, 10, 8) {real, imag} */,
  {32'h412fd430, 32'hc104be5c} /* (30, 10, 7) {real, imag} */,
  {32'h411041f0, 32'hc15a4c05} /* (30, 10, 6) {real, imag} */,
  {32'hc0100ce8, 32'hc178d356} /* (30, 10, 5) {real, imag} */,
  {32'hc10431b7, 32'h409d77c0} /* (30, 10, 4) {real, imag} */,
  {32'hc0068e04, 32'hc08f6441} /* (30, 10, 3) {real, imag} */,
  {32'h41b5da63, 32'hc0b2b170} /* (30, 10, 2) {real, imag} */,
  {32'h41964924, 32'hc06361f4} /* (30, 10, 1) {real, imag} */,
  {32'h4102b895, 32'hc01e4948} /* (30, 10, 0) {real, imag} */,
  {32'hbf39d972, 32'h40966f80} /* (30, 9, 31) {real, imag} */,
  {32'hc0eea73e, 32'hbf018568} /* (30, 9, 30) {real, imag} */,
  {32'hc1039d71, 32'h40b2d30e} /* (30, 9, 29) {real, imag} */,
  {32'hc079a076, 32'h40fcb1c3} /* (30, 9, 28) {real, imag} */,
  {32'h40e7d89f, 32'hbfb47b60} /* (30, 9, 27) {real, imag} */,
  {32'h40b754c0, 32'hbfbaaa18} /* (30, 9, 26) {real, imag} */,
  {32'hbf8e3e7c, 32'hc158465e} /* (30, 9, 25) {real, imag} */,
  {32'hbf720f48, 32'hc1dac6e8} /* (30, 9, 24) {real, imag} */,
  {32'hc0823778, 32'hc0fdf5f6} /* (30, 9, 23) {real, imag} */,
  {32'h40821cbd, 32'hc0d34fa8} /* (30, 9, 22) {real, imag} */,
  {32'hc0f75cb5, 32'hc0f02a58} /* (30, 9, 21) {real, imag} */,
  {32'hc1ec2585, 32'h41a7bdf2} /* (30, 9, 20) {real, imag} */,
  {32'hc1e1cfe6, 32'h4182747a} /* (30, 9, 19) {real, imag} */,
  {32'hc129883a, 32'hc0991ab2} /* (30, 9, 18) {real, imag} */,
  {32'hc10764c0, 32'h3ff681fe} /* (30, 9, 17) {real, imag} */,
  {32'hc191a97f, 32'h4067cde8} /* (30, 9, 16) {real, imag} */,
  {32'hc0fb0831, 32'h3dcfd780} /* (30, 9, 15) {real, imag} */,
  {32'hbf42a7a8, 32'hc12b3b73} /* (30, 9, 14) {real, imag} */,
  {32'hc174a62b, 32'hc130812c} /* (30, 9, 13) {real, imag} */,
  {32'hc0ecad84, 32'hc0e4ca4c} /* (30, 9, 12) {real, imag} */,
  {32'hc0417d1e, 32'h3f564da0} /* (30, 9, 11) {real, imag} */,
  {32'h4188742d, 32'h413f76ec} /* (30, 9, 10) {real, imag} */,
  {32'h41a00cd8, 32'h416a55bf} /* (30, 9, 9) {real, imag} */,
  {32'h41bca70b, 32'h4175e497} /* (30, 9, 8) {real, imag} */,
  {32'h422df74c, 32'h3f371be0} /* (30, 9, 7) {real, imag} */,
  {32'h420c6968, 32'h40b42722} /* (30, 9, 6) {real, imag} */,
  {32'h4193dac0, 32'hc15889ac} /* (30, 9, 5) {real, imag} */,
  {32'h412e66d7, 32'hbf2fbf40} /* (30, 9, 4) {real, imag} */,
  {32'hc11a3656, 32'h40fef825} /* (30, 9, 3) {real, imag} */,
  {32'h40f0b67c, 32'hc035fda4} /* (30, 9, 2) {real, imag} */,
  {32'h40cadfe8, 32'hc01d4530} /* (30, 9, 1) {real, imag} */,
  {32'h3ff64deb, 32'h3f8dd7c0} /* (30, 9, 0) {real, imag} */,
  {32'hc1c42fa1, 32'h41a85ce3} /* (30, 8, 31) {real, imag} */,
  {32'hc1b897ec, 32'h41aec438} /* (30, 8, 30) {real, imag} */,
  {32'hc115d058, 32'h41822b14} /* (30, 8, 29) {real, imag} */,
  {32'hc10345d7, 32'h41d9f0a4} /* (30, 8, 28) {real, imag} */,
  {32'hc14f5dc2, 32'h41e09a71} /* (30, 8, 27) {real, imag} */,
  {32'hc15a0bf2, 32'h41816f3b} /* (30, 8, 26) {real, imag} */,
  {32'hc138ef38, 32'h42150e1a} /* (30, 8, 25) {real, imag} */,
  {32'hc1b30799, 32'h42074a56} /* (30, 8, 24) {real, imag} */,
  {32'hc1ce9212, 32'h419e0246} /* (30, 8, 23) {real, imag} */,
  {32'hc17f3b44, 32'h41c75d0e} /* (30, 8, 22) {real, imag} */,
  {32'h4037b2fc, 32'h411654b3} /* (30, 8, 21) {real, imag} */,
  {32'h3ebec8c0, 32'hc1f772c2} /* (30, 8, 20) {real, imag} */,
  {32'h4088fcff, 32'hc220eca3} /* (30, 8, 19) {real, imag} */,
  {32'h40facefa, 32'hc1e3bc00} /* (30, 8, 18) {real, imag} */,
  {32'h40a66608, 32'hc1f0a14c} /* (30, 8, 17) {real, imag} */,
  {32'h415f72b4, 32'hc1fdc80d} /* (30, 8, 16) {real, imag} */,
  {32'h41db8845, 32'hc1bf2100} /* (30, 8, 15) {real, imag} */,
  {32'h419a698f, 32'hc1b8f8af} /* (30, 8, 14) {real, imag} */,
  {32'h41eceb43, 32'hc2032bd4} /* (30, 8, 13) {real, imag} */,
  {32'h422980e7, 32'hc1d5b761} /* (30, 8, 12) {real, imag} */,
  {32'h41c18fe4, 32'hc117df1d} /* (30, 8, 11) {real, imag} */,
  {32'hc0da8790, 32'h416a06d5} /* (30, 8, 10) {real, imag} */,
  {32'hc1066a13, 32'h41d55fca} /* (30, 8, 9) {real, imag} */,
  {32'h413ffd14, 32'h4208ac88} /* (30, 8, 8) {real, imag} */,
  {32'h419ae677, 32'h42072d72} /* (30, 8, 7) {real, imag} */,
  {32'h418e69d3, 32'h421691ce} /* (30, 8, 6) {real, imag} */,
  {32'h40a6e84e, 32'h422697fc} /* (30, 8, 5) {real, imag} */,
  {32'hc1fa1054, 32'h4230f6c0} /* (30, 8, 4) {real, imag} */,
  {32'hc1f0a47c, 32'h421c503e} /* (30, 8, 3) {real, imag} */,
  {32'hc0f7b548, 32'h424e6827} /* (30, 8, 2) {real, imag} */,
  {32'hc1a6c993, 32'h423a9f91} /* (30, 8, 1) {real, imag} */,
  {32'hc1b286ee, 32'h41a2c3f4} /* (30, 8, 0) {real, imag} */,
  {32'h409efb2b, 32'h4070c327} /* (30, 7, 31) {real, imag} */,
  {32'h41b7b845, 32'hc09f3afb} /* (30, 7, 30) {real, imag} */,
  {32'h41a07cb4, 32'hc18d1b9b} /* (30, 7, 29) {real, imag} */,
  {32'h414fea26, 32'hc19babbf} /* (30, 7, 28) {real, imag} */,
  {32'h40266be0, 32'hc1a3c075} /* (30, 7, 27) {real, imag} */,
  {32'h41999cce, 32'h40120544} /* (30, 7, 26) {real, imag} */,
  {32'h40d171b6, 32'h4114586e} /* (30, 7, 25) {real, imag} */,
  {32'h4167ff7c, 32'h40bd01fc} /* (30, 7, 24) {real, imag} */,
  {32'h3f394280, 32'hc1824644} /* (30, 7, 23) {real, imag} */,
  {32'h41110ee2, 32'hc19c871a} /* (30, 7, 22) {real, imag} */,
  {32'hbd394080, 32'hc1380d68} /* (30, 7, 21) {real, imag} */,
  {32'hc13799e0, 32'hc0f020eb} /* (30, 7, 20) {real, imag} */,
  {32'hc097ac0e, 32'h4109f95f} /* (30, 7, 19) {real, imag} */,
  {32'h3fbba2da, 32'h41069165} /* (30, 7, 18) {real, imag} */,
  {32'hc09dc696, 32'h405465a5} /* (30, 7, 17) {real, imag} */,
  {32'hbf529e7e, 32'h41511f4c} /* (30, 7, 16) {real, imag} */,
  {32'hc19386e0, 32'h4099d32a} /* (30, 7, 15) {real, imag} */,
  {32'hc0d259d7, 32'h41414aa3} /* (30, 7, 14) {real, imag} */,
  {32'hc040ec8c, 32'hbf675e28} /* (30, 7, 13) {real, imag} */,
  {32'h410a8ea7, 32'hc0238978} /* (30, 7, 12) {real, imag} */,
  {32'hc142bdbc, 32'h3ffd6800} /* (30, 7, 11) {real, imag} */,
  {32'h408abea9, 32'hc05db6fa} /* (30, 7, 10) {real, imag} */,
  {32'h419e3920, 32'h4099172c} /* (30, 7, 9) {real, imag} */,
  {32'hbe72cc00, 32'hbfa464b8} /* (30, 7, 8) {real, imag} */,
  {32'h40b975f0, 32'h4084f97e} /* (30, 7, 7) {real, imag} */,
  {32'h41568f39, 32'h4022421c} /* (30, 7, 6) {real, imag} */,
  {32'h41b53fe7, 32'hc10ea6c8} /* (30, 7, 5) {real, imag} */,
  {32'h4182de4c, 32'h40a1dc58} /* (30, 7, 4) {real, imag} */,
  {32'h419a4a36, 32'hc140f480} /* (30, 7, 3) {real, imag} */,
  {32'h41e6d7fa, 32'hc159a448} /* (30, 7, 2) {real, imag} */,
  {32'h41377dfc, 32'hc1921d18} /* (30, 7, 1) {real, imag} */,
  {32'h3fa6d82d, 32'hc10c433c} /* (30, 7, 0) {real, imag} */,
  {32'hbef67394, 32'h402faf86} /* (30, 6, 31) {real, imag} */,
  {32'hc0830bfd, 32'h3fbd7852} /* (30, 6, 30) {real, imag} */,
  {32'hc06ac50b, 32'hc1833cc5} /* (30, 6, 29) {real, imag} */,
  {32'h4116b066, 32'hc142fff3} /* (30, 6, 28) {real, imag} */,
  {32'h40e5f4f8, 32'hbd9034c0} /* (30, 6, 27) {real, imag} */,
  {32'hc1473600, 32'h408f0202} /* (30, 6, 26) {real, imag} */,
  {32'hc1d6f262, 32'h418b27be} /* (30, 6, 25) {real, imag} */,
  {32'hc1857446, 32'h41723449} /* (30, 6, 24) {real, imag} */,
  {32'hc17e05d0, 32'h4064924c} /* (30, 6, 23) {real, imag} */,
  {32'h402c8cb2, 32'h3da68200} /* (30, 6, 22) {real, imag} */,
  {32'h41a7502a, 32'hc158012c} /* (30, 6, 21) {real, imag} */,
  {32'h41fd9be0, 32'hc18483e6} /* (30, 6, 20) {real, imag} */,
  {32'h408fd1b5, 32'hc0bcc26d} /* (30, 6, 19) {real, imag} */,
  {32'hc04aaa3c, 32'hc17cc002} /* (30, 6, 18) {real, imag} */,
  {32'h40b0bc99, 32'hc19ab9a8} /* (30, 6, 17) {real, imag} */,
  {32'h4070fe1a, 32'hbedd76c0} /* (30, 6, 16) {real, imag} */,
  {32'hc070edc4, 32'hc08a5e11} /* (30, 6, 15) {real, imag} */,
  {32'h409f6a25, 32'hc0e025aa} /* (30, 6, 14) {real, imag} */,
  {32'h40ed42a1, 32'hc193aa60} /* (30, 6, 13) {real, imag} */,
  {32'h411ae6ec, 32'hc1b8361b} /* (30, 6, 12) {real, imag} */,
  {32'h4062b24d, 32'h400ec9cf} /* (30, 6, 11) {real, imag} */,
  {32'h414f3d81, 32'h41a658d4} /* (30, 6, 10) {real, imag} */,
  {32'h417bfbf8, 32'h4140559c} /* (30, 6, 9) {real, imag} */,
  {32'hbfda1f00, 32'h40d5e4dc} /* (30, 6, 8) {real, imag} */,
  {32'hc1366232, 32'hc11072bc} /* (30, 6, 7) {real, imag} */,
  {32'h41486a9c, 32'h406631fc} /* (30, 6, 6) {real, imag} */,
  {32'h40dcb014, 32'hbe841020} /* (30, 6, 5) {real, imag} */,
  {32'h40a74104, 32'h4180f3fd} /* (30, 6, 4) {real, imag} */,
  {32'h3fdabb40, 32'h41c52243} /* (30, 6, 3) {real, imag} */,
  {32'hbfde581c, 32'h4133f938} /* (30, 6, 2) {real, imag} */,
  {32'hc1359c77, 32'hc1255a99} /* (30, 6, 1) {real, imag} */,
  {32'hc053a27e, 32'hc1c9ac4a} /* (30, 6, 0) {real, imag} */,
  {32'hc1746af5, 32'h423e48f4} /* (30, 5, 31) {real, imag} */,
  {32'hc1e3ee14, 32'h42b46ead} /* (30, 5, 30) {real, imag} */,
  {32'hc1ef82e5, 32'h4297c24f} /* (30, 5, 29) {real, imag} */,
  {32'hc1e2ff91, 32'h4295d945} /* (30, 5, 28) {real, imag} */,
  {32'hc17a6f54, 32'h422c99d5} /* (30, 5, 27) {real, imag} */,
  {32'hc0edc5ce, 32'h418b443b} /* (30, 5, 26) {real, imag} */,
  {32'h40aec7fc, 32'h4201dcc2} /* (30, 5, 25) {real, imag} */,
  {32'hc134f530, 32'h4299e3d5} /* (30, 5, 24) {real, imag} */,
  {32'hc1c4ffad, 32'h429aa840} /* (30, 5, 23) {real, imag} */,
  {32'hc15f89c3, 32'h426f37bd} /* (30, 5, 22) {real, imag} */,
  {32'hc106d877, 32'h4205ff0f} /* (30, 5, 21) {real, imag} */,
  {32'hc100dccc, 32'hc15e8a8b} /* (30, 5, 20) {real, imag} */,
  {32'h41a9a4ba, 32'hc1e27913} /* (30, 5, 19) {real, imag} */,
  {32'h4194b5a4, 32'hc1862d7c} /* (30, 5, 18) {real, imag} */,
  {32'h41baa0a5, 32'hc20b9d15} /* (30, 5, 17) {real, imag} */,
  {32'h419be238, 32'hc2513f9c} /* (30, 5, 16) {real, imag} */,
  {32'h4210cf17, 32'hc265ff03} /* (30, 5, 15) {real, imag} */,
  {32'h41a6a8ab, 32'hc26059cd} /* (30, 5, 14) {real, imag} */,
  {32'h4055cc0e, 32'hc25b638e} /* (30, 5, 13) {real, imag} */,
  {32'h414987b0, 32'hc1fe8c37} /* (30, 5, 12) {real, imag} */,
  {32'h415904c6, 32'hc209429c} /* (30, 5, 11) {real, imag} */,
  {32'hc0b1e33a, 32'hc152a706} /* (30, 5, 10) {real, imag} */,
  {32'hbf4b2248, 32'h41503c0a} /* (30, 5, 9) {real, imag} */,
  {32'hc0315fba, 32'h40fd088a} /* (30, 5, 8) {real, imag} */,
  {32'h411bc4f5, 32'h41a7aece} /* (30, 5, 7) {real, imag} */,
  {32'hc040d18c, 32'h4201c6dd} /* (30, 5, 6) {real, imag} */,
  {32'hc160cb6a, 32'h426d25c0} /* (30, 5, 5) {real, imag} */,
  {32'hc2181e10, 32'h4280e2a0} /* (30, 5, 4) {real, imag} */,
  {32'hc1c44e24, 32'h425aa956} /* (30, 5, 3) {real, imag} */,
  {32'hc1542f14, 32'h42379e9e} /* (30, 5, 2) {real, imag} */,
  {32'hc20727ed, 32'h426ca5a7} /* (30, 5, 1) {real, imag} */,
  {32'hc1b453b4, 32'h4235c4be} /* (30, 5, 0) {real, imag} */,
  {32'h3ff53eee, 32'hc18915d2} /* (30, 4, 31) {real, imag} */,
  {32'h3f86fc14, 32'hc19d06ad} /* (30, 4, 30) {real, imag} */,
  {32'h400f0d6e, 32'hc205c36c} /* (30, 4, 29) {real, imag} */,
  {32'h411e88fb, 32'hc27826d4} /* (30, 4, 28) {real, imag} */,
  {32'h416466fa, 32'hc285a008} /* (30, 4, 27) {real, imag} */,
  {32'h413d86c3, 32'hc2413c0f} /* (30, 4, 26) {real, imag} */,
  {32'hc0d931bc, 32'hc1fc6452} /* (30, 4, 25) {real, imag} */,
  {32'h3efb74f0, 32'hc239e3ad} /* (30, 4, 24) {real, imag} */,
  {32'h4173f118, 32'hc1d5caa8} /* (30, 4, 23) {real, imag} */,
  {32'h40ca7520, 32'hc215fa30} /* (30, 4, 22) {real, imag} */,
  {32'hc0bdb5fc, 32'hc19a11b6} /* (30, 4, 21) {real, imag} */,
  {32'hc2344772, 32'h428a08eb} /* (30, 4, 20) {real, imag} */,
  {32'hc2809db4, 32'h42951a52} /* (30, 4, 19) {real, imag} */,
  {32'hc2a862fb, 32'h42901167} /* (30, 4, 18) {real, imag} */,
  {32'hc291e856, 32'h42a02079} /* (30, 4, 17) {real, imag} */,
  {32'hc2574e6e, 32'h429e7224} /* (30, 4, 16) {real, imag} */,
  {32'hc12d19bc, 32'h428bec75} /* (30, 4, 15) {real, imag} */,
  {32'hc1ba9ea6, 32'h42800b2e} /* (30, 4, 14) {real, imag} */,
  {32'hc1adf271, 32'h422141f8} /* (30, 4, 13) {real, imag} */,
  {32'hc0876a75, 32'h420feb74} /* (30, 4, 12) {real, imag} */,
  {32'hbf09ba38, 32'h41a3e2a2} /* (30, 4, 11) {real, imag} */,
  {32'h4245fd28, 32'hc282e3f9} /* (30, 4, 10) {real, imag} */,
  {32'h425083a4, 32'hc2973760} /* (30, 4, 9) {real, imag} */,
  {32'h42140978, 32'hc2b55b8c} /* (30, 4, 8) {real, imag} */,
  {32'h4255f92c, 32'hc2990962} /* (30, 4, 7) {real, imag} */,
  {32'h428cc774, 32'hc293b469} /* (30, 4, 6) {real, imag} */,
  {32'h41f311b4, 32'hc24561ef} /* (30, 4, 5) {real, imag} */,
  {32'h41ba8afa, 32'hc20fb4b0} /* (30, 4, 4) {real, imag} */,
  {32'h41a27028, 32'hc25609d0} /* (30, 4, 3) {real, imag} */,
  {32'h410e7e62, 32'hc27023a9} /* (30, 4, 2) {real, imag} */,
  {32'hbf440c10, 32'hc1cb2ad4} /* (30, 4, 1) {real, imag} */,
  {32'hc0fdcdc6, 32'hc10f1d5e} /* (30, 4, 0) {real, imag} */,
  {32'h4152e584, 32'hc12c8846} /* (30, 3, 31) {real, imag} */,
  {32'hc08f3612, 32'hc076ba22} /* (30, 3, 30) {real, imag} */,
  {32'hc079c8b6, 32'hc0b8c4a6} /* (30, 3, 29) {real, imag} */,
  {32'hc19e3b4e, 32'hc1001367} /* (30, 3, 28) {real, imag} */,
  {32'hc20715ac, 32'hc0397ef0} /* (30, 3, 27) {real, imag} */,
  {32'hbf804358, 32'h40361e86} /* (30, 3, 26) {real, imag} */,
  {32'hbecf4e40, 32'h421ebf28} /* (30, 3, 25) {real, imag} */,
  {32'hc10d0a5f, 32'h41ffeac2} /* (30, 3, 24) {real, imag} */,
  {32'hc0b751f8, 32'hc117f354} /* (30, 3, 23) {real, imag} */,
  {32'h402e862b, 32'hc10fb328} /* (30, 3, 22) {real, imag} */,
  {32'hc1cff6d9, 32'h405a3a0c} /* (30, 3, 21) {real, imag} */,
  {32'hc296d72c, 32'h3fb8797e} /* (30, 3, 20) {real, imag} */,
  {32'hc2c70049, 32'h40eadec8} /* (30, 3, 19) {real, imag} */,
  {32'hc2cb0f24, 32'h4151bd80} /* (30, 3, 18) {real, imag} */,
  {32'hc2c16c22, 32'hc0360be0} /* (30, 3, 17) {real, imag} */,
  {32'hc29e7aa6, 32'h414096de} /* (30, 3, 16) {real, imag} */,
  {32'hc21680a3, 32'h40b20b3b} /* (30, 3, 15) {real, imag} */,
  {32'hc180134e, 32'h4089c726} /* (30, 3, 14) {real, imag} */,
  {32'h411e4e5a, 32'h415f10c8} /* (30, 3, 13) {real, imag} */,
  {32'hc0de3792, 32'hbe604d40} /* (30, 3, 12) {real, imag} */,
  {32'h416df54c, 32'hc1132662} /* (30, 3, 11) {real, imag} */,
  {32'h4261c97a, 32'hc11803e0} /* (30, 3, 10) {real, imag} */,
  {32'h42b2ec5d, 32'hc150f750} /* (30, 3, 9) {real, imag} */,
  {32'h4293a825, 32'hc0e6d824} /* (30, 3, 8) {real, imag} */,
  {32'h429d0c49, 32'hc16e4b75} /* (30, 3, 7) {real, imag} */,
  {32'h42cbc13f, 32'h405f0150} /* (30, 3, 6) {real, imag} */,
  {32'h4254774a, 32'h40cb7b60} /* (30, 3, 5) {real, imag} */,
  {32'h41ae2e98, 32'hc1a1b901} /* (30, 3, 4) {real, imag} */,
  {32'hc13056a5, 32'hc0b4dde9} /* (30, 3, 3) {real, imag} */,
  {32'hc1c1a732, 32'h3fb46ef4} /* (30, 3, 2) {real, imag} */,
  {32'h4158a7f0, 32'h40950484} /* (30, 3, 1) {real, imag} */,
  {32'h413be48d, 32'hc093f58e} /* (30, 3, 0) {real, imag} */,
  {32'h411482b8, 32'h428977e1} /* (30, 2, 31) {real, imag} */,
  {32'h40eb1dfc, 32'h430cffec} /* (30, 2, 30) {real, imag} */,
  {32'hc1db3976, 32'h43246107} /* (30, 2, 29) {real, imag} */,
  {32'hc0bc5fdc, 32'h4311106a} /* (30, 2, 28) {real, imag} */,
  {32'h41c0b7c0, 32'h431fc4b2} /* (30, 2, 27) {real, imag} */,
  {32'h41e96f10, 32'h4327a7b4} /* (30, 2, 26) {real, imag} */,
  {32'h4216b22a, 32'h431ff714} /* (30, 2, 25) {real, imag} */,
  {32'h41d67b75, 32'h43048cd4} /* (30, 2, 24) {real, imag} */,
  {32'h41859c5e, 32'h42f4da3c} /* (30, 2, 23) {real, imag} */,
  {32'h40418a80, 32'h431692f1} /* (30, 2, 22) {real, imag} */,
  {32'hc2453f1e, 32'h42b665e1} /* (30, 2, 21) {real, imag} */,
  {32'hc2e34cdd, 32'hc30a972a} /* (30, 2, 20) {real, imag} */,
  {32'hc2e23ff5, 32'hc339a2f8} /* (30, 2, 19) {real, imag} */,
  {32'hc2efae82, 32'hc33e660c} /* (30, 2, 18) {real, imag} */,
  {32'hc301d72c, 32'hc32faa66} /* (30, 2, 17) {real, imag} */,
  {32'hc2db0be6, 32'hc33006d9} /* (30, 2, 16) {real, imag} */,
  {32'hc264218a, 32'hc31cc271} /* (30, 2, 15) {real, imag} */,
  {32'hc0465868, 32'hc3042d65} /* (30, 2, 14) {real, imag} */,
  {32'hbf3e9a60, 32'hc2dc97e7} /* (30, 2, 13) {real, imag} */,
  {32'hc181c705, 32'hc30eca68} /* (30, 2, 12) {real, imag} */,
  {32'h41374892, 32'hc2f729c0} /* (30, 2, 11) {real, imag} */,
  {32'h42be94ec, 32'h42af8085} /* (30, 2, 10) {real, imag} */,
  {32'h431529be, 32'h43470e7d} /* (30, 2, 9) {real, imag} */,
  {32'h42fd2959, 32'h43468a9e} /* (30, 2, 8) {real, imag} */,
  {32'h42d0badc, 32'h433b7f8b} /* (30, 2, 7) {real, imag} */,
  {32'h42cc641c, 32'h4344594e} /* (30, 2, 6) {real, imag} */,
  {32'h4257aa1e, 32'h431b5db9} /* (30, 2, 5) {real, imag} */,
  {32'h413f7863, 32'h42e8ab0c} /* (30, 2, 4) {real, imag} */,
  {32'hc17cd3c0, 32'h430aeba2} /* (30, 2, 3) {real, imag} */,
  {32'h4100cf24, 32'h43150710} /* (30, 2, 2) {real, imag} */,
  {32'hc10aee54, 32'h431ef445} /* (30, 2, 1) {real, imag} */,
  {32'hbea11000, 32'h42afa563} /* (30, 2, 0) {real, imag} */,
  {32'hc18dc3a3, 32'hc2fd79ed} /* (30, 1, 31) {real, imag} */,
  {32'hc1afe036, 32'hc368fe95} /* (30, 1, 30) {real, imag} */,
  {32'hc21de24e, 32'hc3758503} /* (30, 1, 29) {real, imag} */,
  {32'hc1cd0438, 32'hc383130a} /* (30, 1, 28) {real, imag} */,
  {32'hc186e05e, 32'hc37cb755} /* (30, 1, 27) {real, imag} */,
  {32'hc178487b, 32'hc3684d5a} /* (30, 1, 26) {real, imag} */,
  {32'hc20bbb62, 32'hc36e8b28} /* (30, 1, 25) {real, imag} */,
  {32'hc2332127, 32'hc37b1337} /* (30, 1, 24) {real, imag} */,
  {32'hc110d5c0, 32'hc3758636} /* (30, 1, 23) {real, imag} */,
  {32'hc1189e34, 32'hc360bbc7} /* (30, 1, 22) {real, imag} */,
  {32'hc22e6fd8, 32'hc2f9075a} /* (30, 1, 21) {real, imag} */,
  {32'hc2a373d8, 32'h42b90b54} /* (30, 1, 20) {real, imag} */,
  {32'hc2db814f, 32'h430436f8} /* (30, 1, 19) {real, imag} */,
  {32'hc2dfbe5a, 32'h42d3b782} /* (30, 1, 18) {real, imag} */,
  {32'hc2b46180, 32'h42e076bc} /* (30, 1, 17) {real, imag} */,
  {32'hc21eb0a3, 32'h4308fdad} /* (30, 1, 16) {real, imag} */,
  {32'h41ea3934, 32'h4356f50f} /* (30, 1, 15) {real, imag} */,
  {32'h41e45cb6, 32'h4365db49} /* (30, 1, 14) {real, imag} */,
  {32'h41a3ae80, 32'h43702677} /* (30, 1, 13) {real, imag} */,
  {32'h41ec25de, 32'h436ea5ac} /* (30, 1, 12) {real, imag} */,
  {32'h420926f2, 32'h4343ed39} /* (30, 1, 11) {real, imag} */,
  {32'h4243e4f2, 32'hc10e892c} /* (30, 1, 10) {real, imag} */,
  {32'h429fb3f5, 32'hc2f32066} /* (30, 1, 9) {real, imag} */,
  {32'h42bf5452, 32'hc3004c2e} /* (30, 1, 8) {real, imag} */,
  {32'h42a1c653, 32'hc2f5f36b} /* (30, 1, 7) {real, imag} */,
  {32'h42942e28, 32'hc3047961} /* (30, 1, 6) {real, imag} */,
  {32'hbf142aa0, 32'hc342a6e0} /* (30, 1, 5) {real, imag} */,
  {32'hc262abb6, 32'hc365e5f9} /* (30, 1, 4) {real, imag} */,
  {32'hc2523be1, 32'hc3703d22} /* (30, 1, 3) {real, imag} */,
  {32'hc239e167, 32'hc37cefe8} /* (30, 1, 2) {real, imag} */,
  {32'hc1c55872, 32'hc3675002} /* (30, 1, 1) {real, imag} */,
  {32'hc008b730, 32'hc2f71240} /* (30, 1, 0) {real, imag} */,
  {32'hc20a9050, 32'hc295c748} /* (30, 0, 31) {real, imag} */,
  {32'hc1c417e4, 32'hc2ff62f4} /* (30, 0, 30) {real, imag} */,
  {32'hc189d400, 32'hc3188fb7} /* (30, 0, 29) {real, imag} */,
  {32'hc1cde45c, 32'hc309c693} /* (30, 0, 28) {real, imag} */,
  {32'hc21da660, 32'hc31c51fa} /* (30, 0, 27) {real, imag} */,
  {32'hc1fd430a, 32'hc32c2c34} /* (30, 0, 26) {real, imag} */,
  {32'hc131bd66, 32'hc3220fc1} /* (30, 0, 25) {real, imag} */,
  {32'hc1a8f3d7, 32'hc325a230} /* (30, 0, 24) {real, imag} */,
  {32'hc250d411, 32'hc3146364} /* (30, 0, 23) {real, imag} */,
  {32'hc208b272, 32'hc30b9da4} /* (30, 0, 22) {real, imag} */,
  {32'hc17eba7f, 32'hc2f5a33a} /* (30, 0, 21) {real, imag} */,
  {32'h40b1c618, 32'hc210da3e} /* (30, 0, 20) {real, imag} */,
  {32'h4171b1e7, 32'hc0e67e0e} /* (30, 0, 19) {real, imag} */,
  {32'hc18e002c, 32'hc0bb60d6} /* (30, 0, 18) {real, imag} */,
  {32'hc1650fd8, 32'hc19e04b2} /* (30, 0, 17) {real, imag} */,
  {32'h40169cfa, 32'h41f5e61e} /* (30, 0, 16) {real, imag} */,
  {32'h416367ec, 32'h430585c0} /* (30, 0, 15) {real, imag} */,
  {32'h41815e08, 32'h4322467c} /* (30, 0, 14) {real, imag} */,
  {32'h41e890ea, 32'h43080118} /* (30, 0, 13) {real, imag} */,
  {32'h422a3708, 32'h4312a848} /* (30, 0, 12) {real, imag} */,
  {32'h425d8a60, 32'h4304be7c} /* (30, 0, 11) {real, imag} */,
  {32'h3b405800, 32'h42728c2e} /* (30, 0, 10) {real, imag} */,
  {32'hc09a0322, 32'hc198e6fe} /* (30, 0, 9) {real, imag} */,
  {32'h406a8df4, 32'hc152b42b} /* (30, 0, 8) {real, imag} */,
  {32'hc17a3018, 32'h417cbf90} /* (30, 0, 7) {real, imag} */,
  {32'hc0c9702a, 32'hc078b77a} /* (30, 0, 6) {real, imag} */,
  {32'hc1ed324a, 32'hc2ba09a9} /* (30, 0, 5) {real, imag} */,
  {32'hc22a992e, 32'hc326c21e} /* (30, 0, 4) {real, imag} */,
  {32'hc1189c0d, 32'hc3240dfb} /* (30, 0, 3) {real, imag} */,
  {32'hc1d5932c, 32'hc321481e} /* (30, 0, 2) {real, imag} */,
  {32'hc2241018, 32'hc2f3d462} /* (30, 0, 1) {real, imag} */,
  {32'hc1f3f8bc, 32'hc289b18f} /* (30, 0, 0) {real, imag} */,
  {32'hc1858fea, 32'hc26d7393} /* (29, 31, 31) {real, imag} */,
  {32'hc1fe9c60, 32'hc2c9b9aa} /* (29, 31, 30) {real, imag} */,
  {32'hc1a7df75, 32'hc2a6d148} /* (29, 31, 29) {real, imag} */,
  {32'hc1fbd204, 32'hc28eb754} /* (29, 31, 28) {real, imag} */,
  {32'hc263e570, 32'hc2a5da49} /* (29, 31, 27) {real, imag} */,
  {32'hc250ffc4, 32'hc2c6660d} /* (29, 31, 26) {real, imag} */,
  {32'hc27803c8, 32'hc2e7d2a4} /* (29, 31, 25) {real, imag} */,
  {32'hc2230b40, 32'hc2d9a8e9} /* (29, 31, 24) {real, imag} */,
  {32'hc1f10685, 32'hc2990b4b} /* (29, 31, 23) {real, imag} */,
  {32'hc22ce712, 32'hc2a8f8ca} /* (29, 31, 22) {real, imag} */,
  {32'hc09917e5, 32'hc227c80d} /* (29, 31, 21) {real, imag} */,
  {32'h427971d8, 32'h42381e80} /* (29, 31, 20) {real, imag} */,
  {32'h429366bc, 32'h4238c4a2} /* (29, 31, 19) {real, imag} */,
  {32'h429c5416, 32'h41ecc052} /* (29, 31, 18) {real, imag} */,
  {32'h4240bf38, 32'h4206dc9f} /* (29, 31, 17) {real, imag} */,
  {32'h41c61e88, 32'h41f356ad} /* (29, 31, 16) {real, imag} */,
  {32'h41b27e12, 32'h4295273e} /* (29, 31, 15) {real, imag} */,
  {32'h423cd3b8, 32'h42a3133b} /* (29, 31, 14) {real, imag} */,
  {32'h41c53241, 32'h42c3af23} /* (29, 31, 13) {real, imag} */,
  {32'h409ce44a, 32'h42a18535} /* (29, 31, 12) {real, imag} */,
  {32'h41a00da9, 32'h428628e0} /* (29, 31, 11) {real, imag} */,
  {32'hc1906d58, 32'h412cea9a} /* (29, 31, 10) {real, imag} */,
  {32'hc2404ab3, 32'hc217e1a6} /* (29, 31, 9) {real, imag} */,
  {32'hc21e3be5, 32'hc211abf4} /* (29, 31, 8) {real, imag} */,
  {32'hc2212910, 32'hc19667ee} /* (29, 31, 7) {real, imag} */,
  {32'hc20bf3fd, 32'hc171406e} /* (29, 31, 6) {real, imag} */,
  {32'hc27394a2, 32'hc262039c} /* (29, 31, 5) {real, imag} */,
  {32'hc207620e, 32'hc2b7d3ae} /* (29, 31, 4) {real, imag} */,
  {32'hc21c5808, 32'hc2eb421c} /* (29, 31, 3) {real, imag} */,
  {32'hc23c1f25, 32'hc2e0d402} /* (29, 31, 2) {real, imag} */,
  {32'hc18923c2, 32'hc2b41fa1} /* (29, 31, 1) {real, imag} */,
  {32'hc100d2b1, 32'hc248c567} /* (29, 31, 0) {real, imag} */,
  {32'h40e5466b, 32'h421f15a9} /* (29, 30, 31) {real, imag} */,
  {32'h41a0dd1e, 32'h4247cc10} /* (29, 30, 30) {real, imag} */,
  {32'h41cd2eed, 32'h425258f3} /* (29, 30, 29) {real, imag} */,
  {32'h42040ac9, 32'h4244a1ef} /* (29, 30, 28) {real, imag} */,
  {32'h42274d58, 32'h421cbd72} /* (29, 30, 27) {real, imag} */,
  {32'h41ed5d87, 32'h4215842e} /* (29, 30, 26) {real, imag} */,
  {32'h41e9126e, 32'h4214a372} /* (29, 30, 25) {real, imag} */,
  {32'h42013942, 32'h42063a46} /* (29, 30, 24) {real, imag} */,
  {32'h41ef9988, 32'h425fb53c} /* (29, 30, 23) {real, imag} */,
  {32'h41fd038b, 32'h4221ba70} /* (29, 30, 22) {real, imag} */,
  {32'h41a4b18e, 32'h40e880b4} /* (29, 30, 21) {real, imag} */,
  {32'h41ea86df, 32'hc28de2d3} /* (29, 30, 20) {real, imag} */,
  {32'h416943d4, 32'hc2bdcf4e} /* (29, 30, 19) {real, imag} */,
  {32'h40291f90, 32'hc2c1b0ca} /* (29, 30, 18) {real, imag} */,
  {32'h411138be, 32'hc2d9b40f} /* (29, 30, 17) {real, imag} */,
  {32'hc109ec03, 32'hc2a806dd} /* (29, 30, 16) {real, imag} */,
  {32'hc1e2921a, 32'hc25c9d64} /* (29, 30, 15) {real, imag} */,
  {32'hc192119c, 32'hc2824f0a} /* (29, 30, 14) {real, imag} */,
  {32'hc1c10ec0, 32'hc211fa36} /* (29, 30, 13) {real, imag} */,
  {32'hc1becdca, 32'hc1c3e797} /* (29, 30, 12) {real, imag} */,
  {32'hc1bda720, 32'hc15b9a66} /* (29, 30, 11) {real, imag} */,
  {32'hc1cfcad4, 32'h42168416} /* (29, 30, 10) {real, imag} */,
  {32'hc0cd4790, 32'h42aa1867} /* (29, 30, 9) {real, imag} */,
  {32'hc027dd00, 32'h4299d16f} /* (29, 30, 8) {real, imag} */,
  {32'hc1637934, 32'h42938c60} /* (29, 30, 7) {real, imag} */,
  {32'h40a935f8, 32'h42a3d57b} /* (29, 30, 6) {real, imag} */,
  {32'h41efadbb, 32'h42801d1f} /* (29, 30, 5) {real, imag} */,
  {32'h40e04056, 32'h42433320} /* (29, 30, 4) {real, imag} */,
  {32'h40b2eb38, 32'h426bef84} /* (29, 30, 3) {real, imag} */,
  {32'h418a5201, 32'h4257c6b1} /* (29, 30, 2) {real, imag} */,
  {32'h41f5ab50, 32'h4204ed19} /* (29, 30, 1) {real, imag} */,
  {32'h419b81c6, 32'h41f475a6} /* (29, 30, 0) {real, imag} */,
  {32'h40c0f65c, 32'hbec0f5a0} /* (29, 29, 31) {real, imag} */,
  {32'hbff2c0a0, 32'hc08ce909} /* (29, 29, 30) {real, imag} */,
  {32'hc1247e5d, 32'h4137d295} /* (29, 29, 29) {real, imag} */,
  {32'h411ed09e, 32'h41cfc2f0} /* (29, 29, 28) {real, imag} */,
  {32'h41208bb1, 32'h40a00c58} /* (29, 29, 27) {real, imag} */,
  {32'h41a8da49, 32'h41bbbad0} /* (29, 29, 26) {real, imag} */,
  {32'hc02211ca, 32'h418c8d72} /* (29, 29, 25) {real, imag} */,
  {32'hc04bb6be, 32'h41b41b44} /* (29, 29, 24) {real, imag} */,
  {32'hc14bc5a0, 32'h40e74c1c} /* (29, 29, 23) {real, imag} */,
  {32'hc169cd1f, 32'h415ec34d} /* (29, 29, 22) {real, imag} */,
  {32'h4147ee0a, 32'hc12a1f14} /* (29, 29, 21) {real, imag} */,
  {32'h41cd4255, 32'hc204c688} /* (29, 29, 20) {real, imag} */,
  {32'h41c34176, 32'hc1b4e839} /* (29, 29, 19) {real, imag} */,
  {32'h41419110, 32'hc0d896da} /* (29, 29, 18) {real, imag} */,
  {32'h4199d683, 32'hc0d424cb} /* (29, 29, 17) {real, imag} */,
  {32'h4240ca16, 32'hc1025c49} /* (29, 29, 16) {real, imag} */,
  {32'hc113848e, 32'hc0ba93f6} /* (29, 29, 15) {real, imag} */,
  {32'hc20f258b, 32'h4171bb11} /* (29, 29, 14) {real, imag} */,
  {32'hc149aed2, 32'h404da368} /* (29, 29, 13) {real, imag} */,
  {32'h41bcc4c4, 32'hc11a3c45} /* (29, 29, 12) {real, imag} */,
  {32'h415b0342, 32'hc1998e3c} /* (29, 29, 11) {real, imag} */,
  {32'hc1828e7b, 32'h4190e180} /* (29, 29, 10) {real, imag} */,
  {32'hc136f8f8, 32'h4257b8fb} /* (29, 29, 9) {real, imag} */,
  {32'hc19a1d82, 32'h41a910b0} /* (29, 29, 8) {real, imag} */,
  {32'hc21af24e, 32'h4191bdf1} /* (29, 29, 7) {real, imag} */,
  {32'hc1d14ac9, 32'h4177cb51} /* (29, 29, 6) {real, imag} */,
  {32'hc0090c00, 32'h41a45ace} /* (29, 29, 5) {real, imag} */,
  {32'hc1101dfe, 32'h409d2119} /* (29, 29, 4) {real, imag} */,
  {32'hc1398869, 32'hc145249c} /* (29, 29, 3) {real, imag} */,
  {32'hc130a42a, 32'h414822a1} /* (29, 29, 2) {real, imag} */,
  {32'hc1af7efc, 32'h41875c3a} /* (29, 29, 1) {real, imag} */,
  {32'h3f5e48c8, 32'h40304c7c} /* (29, 29, 0) {real, imag} */,
  {32'h401321d9, 32'hc107a78d} /* (29, 28, 31) {real, imag} */,
  {32'hbfd41e28, 32'hc1959810} /* (29, 28, 30) {real, imag} */,
  {32'hc184c9de, 32'hc1aa0498} /* (29, 28, 29) {real, imag} */,
  {32'hc0da2360, 32'hc10601a1} /* (29, 28, 28) {real, imag} */,
  {32'hc179ad0c, 32'hc10eefa6} /* (29, 28, 27) {real, imag} */,
  {32'hc19a5ab6, 32'hc1a73204} /* (29, 28, 26) {real, imag} */,
  {32'hc139c6d6, 32'hc1ac8d9e} /* (29, 28, 25) {real, imag} */,
  {32'hc1264026, 32'hc1ea320a} /* (29, 28, 24) {real, imag} */,
  {32'hc1b0c792, 32'hc21426d6} /* (29, 28, 23) {real, imag} */,
  {32'hc18ea860, 32'hc217a1fe} /* (29, 28, 22) {real, imag} */,
  {32'h403e6370, 32'hc12d6f3b} /* (29, 28, 21) {real, imag} */,
  {32'h41d1c521, 32'h418f80f6} /* (29, 28, 20) {real, imag} */,
  {32'h41c0e0e9, 32'h41aaf725} /* (29, 28, 19) {real, imag} */,
  {32'h41eaa807, 32'h41bbbe3c} /* (29, 28, 18) {real, imag} */,
  {32'h41e41264, 32'h41a8fba3} /* (29, 28, 17) {real, imag} */,
  {32'h414da16f, 32'hc035c330} /* (29, 28, 16) {real, imag} */,
  {32'h4197d451, 32'hc1467199} /* (29, 28, 15) {real, imag} */,
  {32'h422759ea, 32'h3f841a60} /* (29, 28, 14) {real, imag} */,
  {32'h4200d4b8, 32'h406f43a8} /* (29, 28, 13) {real, imag} */,
  {32'h4158173b, 32'h40ca6f94} /* (29, 28, 12) {real, imag} */,
  {32'h4109b47a, 32'h4169b6f6} /* (29, 28, 11) {real, imag} */,
  {32'hc1b8356c, 32'hc141136e} /* (29, 28, 10) {real, imag} */,
  {32'hc1b1775d, 32'hc1b2dc60} /* (29, 28, 9) {real, imag} */,
  {32'hc1efe455, 32'hc1e10d93} /* (29, 28, 8) {real, imag} */,
  {32'hc23368f3, 32'hc1ff77c8} /* (29, 28, 7) {real, imag} */,
  {32'hc2232411, 32'hc201d3ba} /* (29, 28, 6) {real, imag} */,
  {32'hbfc1a510, 32'hc1c43c0c} /* (29, 28, 5) {real, imag} */,
  {32'h3f197764, 32'hc1a2c03a} /* (29, 28, 4) {real, imag} */,
  {32'hc127d79e, 32'hc1fbc8e6} /* (29, 28, 3) {real, imag} */,
  {32'hc1ad9433, 32'hc1f06e4f} /* (29, 28, 2) {real, imag} */,
  {32'hc1433e18, 32'hc1e70ab9} /* (29, 28, 1) {real, imag} */,
  {32'h41387747, 32'hc107c674} /* (29, 28, 0) {real, imag} */,
  {32'h41686846, 32'h41a3cf3e} /* (29, 27, 31) {real, imag} */,
  {32'h41075b2c, 32'h41a9f41a} /* (29, 27, 30) {real, imag} */,
  {32'h4194ad1b, 32'h4174f1ea} /* (29, 27, 29) {real, imag} */,
  {32'h41df692c, 32'h41afec96} /* (29, 27, 28) {real, imag} */,
  {32'h421258ca, 32'h4222c786} /* (29, 27, 27) {real, imag} */,
  {32'h4199008a, 32'h422e4390} /* (29, 27, 26) {real, imag} */,
  {32'h412907fa, 32'h4220378e} /* (29, 27, 25) {real, imag} */,
  {32'h41d57090, 32'h41b3b8cb} /* (29, 27, 24) {real, imag} */,
  {32'h40d03199, 32'h4198bc10} /* (29, 27, 23) {real, imag} */,
  {32'h4143c512, 32'h417d5ef2} /* (29, 27, 22) {real, imag} */,
  {32'h41b2ada4, 32'h4177c8b3} /* (29, 27, 21) {real, imag} */,
  {32'hc03e4a3a, 32'hc0d2de54} /* (29, 27, 20) {real, imag} */,
  {32'hc19d1d26, 32'hc1e70520} /* (29, 27, 19) {real, imag} */,
  {32'hc1980f02, 32'hc1970d7d} /* (29, 27, 18) {real, imag} */,
  {32'hc1a6f617, 32'hc10c2790} /* (29, 27, 17) {real, imag} */,
  {32'hc1779e5a, 32'hc1b31cb8} /* (29, 27, 16) {real, imag} */,
  {32'h41446a31, 32'hc1a66eba} /* (29, 27, 15) {real, imag} */,
  {32'hc10cdf1c, 32'hc18bd64a} /* (29, 27, 14) {real, imag} */,
  {32'hc1b9617e, 32'hc0f4070c} /* (29, 27, 13) {real, imag} */,
  {32'hc1cb9bff, 32'hc1915890} /* (29, 27, 12) {real, imag} */,
  {32'hc1cc18d9, 32'hc1c6a34d} /* (29, 27, 11) {real, imag} */,
  {32'hc1265dde, 32'hc0e35b46} /* (29, 27, 10) {real, imag} */,
  {32'hc0f0fa1a, 32'h41aed73c} /* (29, 27, 9) {real, imag} */,
  {32'h41121e42, 32'h41c20e17} /* (29, 27, 8) {real, imag} */,
  {32'h4098bf57, 32'h40f96a80} /* (29, 27, 7) {real, imag} */,
  {32'hc11da98d, 32'hbffadfb8} /* (29, 27, 6) {real, imag} */,
  {32'h3ebe78c0, 32'h4169b676} /* (29, 27, 5) {real, imag} */,
  {32'h418805d2, 32'h41aa0e64} /* (29, 27, 4) {real, imag} */,
  {32'h422ed4ce, 32'h41d5929d} /* (29, 27, 3) {real, imag} */,
  {32'h41bd1296, 32'h410afdf3} /* (29, 27, 2) {real, imag} */,
  {32'h40d51b91, 32'h41752900} /* (29, 27, 1) {real, imag} */,
  {32'h41276e2e, 32'h40e37c8c} /* (29, 27, 0) {real, imag} */,
  {32'h40174fc8, 32'hc032dd62} /* (29, 26, 31) {real, imag} */,
  {32'h4124b6ac, 32'h41893bb6} /* (29, 26, 30) {real, imag} */,
  {32'h40d68a2d, 32'h410121e2} /* (29, 26, 29) {real, imag} */,
  {32'hc17ee366, 32'h4107d362} /* (29, 26, 28) {real, imag} */,
  {32'hc1a0ed03, 32'h3f293308} /* (29, 26, 27) {real, imag} */,
  {32'hbd991560, 32'hc12ad5f7} /* (29, 26, 26) {real, imag} */,
  {32'h3fcd2a96, 32'hc0ff3294} /* (29, 26, 25) {real, imag} */,
  {32'hc11aa1dc, 32'hc0aa4801} /* (29, 26, 24) {real, imag} */,
  {32'hc09e44bd, 32'hc0ffca0a} /* (29, 26, 23) {real, imag} */,
  {32'h410eeb76, 32'hc151f62e} /* (29, 26, 22) {real, imag} */,
  {32'h412c1e96, 32'hc1b7be68} /* (29, 26, 21) {real, imag} */,
  {32'hbf2419b8, 32'h41119d0c} /* (29, 26, 20) {real, imag} */,
  {32'hbf0dc558, 32'h4179ddde} /* (29, 26, 19) {real, imag} */,
  {32'h4081192c, 32'hc0fe0a5f} /* (29, 26, 18) {real, imag} */,
  {32'h414b663e, 32'hc1166b8c} /* (29, 26, 17) {real, imag} */,
  {32'h41400e96, 32'h4053e05e} /* (29, 26, 16) {real, imag} */,
  {32'h40b29b16, 32'hc101c3e1} /* (29, 26, 15) {real, imag} */,
  {32'hc1935a52, 32'hc186306a} /* (29, 26, 14) {real, imag} */,
  {32'h4054468a, 32'h409be11a} /* (29, 26, 13) {real, imag} */,
  {32'h41d8e782, 32'hc0d03c3a} /* (29, 26, 12) {real, imag} */,
  {32'h41330c46, 32'hc14edf35} /* (29, 26, 11) {real, imag} */,
  {32'hc148cb46, 32'hc1b9e18c} /* (29, 26, 10) {real, imag} */,
  {32'hc1384e3a, 32'hc120ba89} /* (29, 26, 9) {real, imag} */,
  {32'h40d2bd90, 32'hc0ba0dc4} /* (29, 26, 8) {real, imag} */,
  {32'h40da2686, 32'hc01fcee0} /* (29, 26, 7) {real, imag} */,
  {32'hc08a27e0, 32'h40ce98d4} /* (29, 26, 6) {real, imag} */,
  {32'h405fe6ce, 32'hc1a848db} /* (29, 26, 5) {real, imag} */,
  {32'h40226e1c, 32'hc14f9d6f} /* (29, 26, 4) {real, imag} */,
  {32'h40e6c070, 32'hbf96914c} /* (29, 26, 3) {real, imag} */,
  {32'h40cd5495, 32'h413d91a3} /* (29, 26, 2) {real, imag} */,
  {32'h40007d34, 32'h41c84fe4} /* (29, 26, 1) {real, imag} */,
  {32'hc110bf59, 32'h41285a2c} /* (29, 26, 0) {real, imag} */,
  {32'h40ce90e0, 32'hc092b3e7} /* (29, 25, 31) {real, imag} */,
  {32'h40f70c04, 32'hc12dc7e9} /* (29, 25, 30) {real, imag} */,
  {32'hc0cb562a, 32'h40ea439c} /* (29, 25, 29) {real, imag} */,
  {32'h4033b466, 32'h41788ce7} /* (29, 25, 28) {real, imag} */,
  {32'hc0c2b7fe, 32'hc0b75928} /* (29, 25, 27) {real, imag} */,
  {32'hbffecc7e, 32'hbfdf01c8} /* (29, 25, 26) {real, imag} */,
  {32'h40a4fc74, 32'hc0a4093a} /* (29, 25, 25) {real, imag} */,
  {32'hc01b8e74, 32'hc0964852} /* (29, 25, 24) {real, imag} */,
  {32'h409fdcef, 32'hc17ef06f} /* (29, 25, 23) {real, imag} */,
  {32'h408f708f, 32'hc197dbd6} /* (29, 25, 22) {real, imag} */,
  {32'h3fc3b0fc, 32'hc160b5c6} /* (29, 25, 21) {real, imag} */,
  {32'h409c0fd7, 32'hc1819aee} /* (29, 25, 20) {real, imag} */,
  {32'h40faa918, 32'h418780b4} /* (29, 25, 19) {real, imag} */,
  {32'h3f8dd37c, 32'h4148c1a0} /* (29, 25, 18) {real, imag} */,
  {32'h40b406f0, 32'hc1189a1d} /* (29, 25, 17) {real, imag} */,
  {32'hc0c57c62, 32'hc1288934} /* (29, 25, 16) {real, imag} */,
  {32'hc1081074, 32'hbe8dba70} /* (29, 25, 15) {real, imag} */,
  {32'hc153606a, 32'hc0ecae34} /* (29, 25, 14) {real, imag} */,
  {32'h4143f782, 32'hc0ba8f87} /* (29, 25, 13) {real, imag} */,
  {32'h40f4991c, 32'h3fb248e4} /* (29, 25, 12) {real, imag} */,
  {32'hc098c8e2, 32'h40a6ac2f} /* (29, 25, 11) {real, imag} */,
  {32'h40619a82, 32'h3f983362} /* (29, 25, 10) {real, imag} */,
  {32'hc14a32e1, 32'hc081d304} /* (29, 25, 9) {real, imag} */,
  {32'hc12aab3a, 32'hc00a2870} /* (29, 25, 8) {real, imag} */,
  {32'hc0dd206c, 32'hc1744a23} /* (29, 25, 7) {real, imag} */,
  {32'h40665527, 32'hc11a6ae1} /* (29, 25, 6) {real, imag} */,
  {32'h408ca149, 32'h404b5c84} /* (29, 25, 5) {real, imag} */,
  {32'hc0c32e7a, 32'h3fb602cc} /* (29, 25, 4) {real, imag} */,
  {32'hc0507dc2, 32'h40a94546} /* (29, 25, 3) {real, imag} */,
  {32'h408a5d90, 32'h4019f0e0} /* (29, 25, 2) {real, imag} */,
  {32'h40c97762, 32'hc12d5c1a} /* (29, 25, 1) {real, imag} */,
  {32'h412e9ff3, 32'hc185807a} /* (29, 25, 0) {real, imag} */,
  {32'h41052712, 32'hc1688b77} /* (29, 24, 31) {real, imag} */,
  {32'h41223358, 32'hbf012d20} /* (29, 24, 30) {real, imag} */,
  {32'h402409fa, 32'h4134fafc} /* (29, 24, 29) {real, imag} */,
  {32'h413239b2, 32'h417989ed} /* (29, 24, 28) {real, imag} */,
  {32'h41906607, 32'h4069542e} /* (29, 24, 27) {real, imag} */,
  {32'h41353b45, 32'hbfce7b78} /* (29, 24, 26) {real, imag} */,
  {32'h418e4200, 32'h4100e819} /* (29, 24, 25) {real, imag} */,
  {32'hbf811960, 32'h41a57444} /* (29, 24, 24) {real, imag} */,
  {32'hc0316730, 32'h414ecc30} /* (29, 24, 23) {real, imag} */,
  {32'h418415e1, 32'hbfb8c524} /* (29, 24, 22) {real, imag} */,
  {32'h411062c3, 32'h4199f8d4} /* (29, 24, 21) {real, imag} */,
  {32'hc1516bd3, 32'h4109f2ca} /* (29, 24, 20) {real, imag} */,
  {32'hbfbdc3fa, 32'hc0f4a864} /* (29, 24, 19) {real, imag} */,
  {32'hc044bbe6, 32'hbf4ec4d0} /* (29, 24, 18) {real, imag} */,
  {32'hc0ff7674, 32'hc18fd2ec} /* (29, 24, 17) {real, imag} */,
  {32'h4045fbfc, 32'hc1f56e1c} /* (29, 24, 16) {real, imag} */,
  {32'h40d296c6, 32'hc1195008} /* (29, 24, 15) {real, imag} */,
  {32'hbf67df40, 32'hbe8f5d80} /* (29, 24, 14) {real, imag} */,
  {32'hc0f34cae, 32'h4069d0e1} /* (29, 24, 13) {real, imag} */,
  {32'hc1906b87, 32'h40f54ec0} /* (29, 24, 12) {real, imag} */,
  {32'hc1569142, 32'h41434084} /* (29, 24, 11) {real, imag} */,
  {32'hc0eaad24, 32'h40112faf} /* (29, 24, 10) {real, imag} */,
  {32'hc0f18018, 32'h406269ae} /* (29, 24, 9) {real, imag} */,
  {32'hc08687ec, 32'h4087f4c1} /* (29, 24, 8) {real, imag} */,
  {32'h403cc018, 32'h3f5eb1e6} /* (29, 24, 7) {real, imag} */,
  {32'h40aad000, 32'h417aef4f} /* (29, 24, 6) {real, imag} */,
  {32'h4157df49, 32'h41a42eab} /* (29, 24, 5) {real, imag} */,
  {32'h415fee8a, 32'h40691aa0} /* (29, 24, 4) {real, imag} */,
  {32'h404d5503, 32'hc089eb4a} /* (29, 24, 3) {real, imag} */,
  {32'h400c99f6, 32'h40b811ee} /* (29, 24, 2) {real, imag} */,
  {32'h40b15642, 32'h418ce311} /* (29, 24, 1) {real, imag} */,
  {32'h3fe07764, 32'h410b63a4} /* (29, 24, 0) {real, imag} */,
  {32'h40719497, 32'h3fda1bec} /* (29, 23, 31) {real, imag} */,
  {32'h40b058d6, 32'hc10d2310} /* (29, 23, 30) {real, imag} */,
  {32'h415442ae, 32'hc1810b00} /* (29, 23, 29) {real, imag} */,
  {32'h40055502, 32'hc0216902} /* (29, 23, 28) {real, imag} */,
  {32'hc048c1aa, 32'h4137caa0} /* (29, 23, 27) {real, imag} */,
  {32'h40e172b7, 32'h40ae8394} /* (29, 23, 26) {real, imag} */,
  {32'h412e9e0e, 32'hbfa233aa} /* (29, 23, 25) {real, imag} */,
  {32'h418c8d38, 32'hc13a8bdb} /* (29, 23, 24) {real, imag} */,
  {32'h41880d37, 32'hc11750bc} /* (29, 23, 23) {real, imag} */,
  {32'h41558d6a, 32'h4130a6dc} /* (29, 23, 22) {real, imag} */,
  {32'h413f34f5, 32'h4180d166} /* (29, 23, 21) {real, imag} */,
  {32'h3f884ed0, 32'h40f1e45c} /* (29, 23, 20) {real, imag} */,
  {32'h40eeca6a, 32'h411f85a3} /* (29, 23, 19) {real, imag} */,
  {32'h4042ab1a, 32'h41246fd6} /* (29, 23, 18) {real, imag} */,
  {32'hbe7e7bc0, 32'h4133066d} /* (29, 23, 17) {real, imag} */,
  {32'h4134300d, 32'hbf2fd254} /* (29, 23, 16) {real, imag} */,
  {32'h4134ca9e, 32'h3f8e5a04} /* (29, 23, 15) {real, imag} */,
  {32'h412dc99d, 32'h400e0503} /* (29, 23, 14) {real, imag} */,
  {32'h4069207e, 32'hc127372e} /* (29, 23, 13) {real, imag} */,
  {32'hc0cfd00a, 32'hc13c12bc} /* (29, 23, 12) {real, imag} */,
  {32'hc1869ad4, 32'hc0b86794} /* (29, 23, 11) {real, imag} */,
  {32'hc189f23e, 32'hbe2df960} /* (29, 23, 10) {real, imag} */,
  {32'hc16e0a2b, 32'hc015667a} /* (29, 23, 9) {real, imag} */,
  {32'hc15065a0, 32'h419088c1} /* (29, 23, 8) {real, imag} */,
  {32'hc01071dc, 32'h415a10cd} /* (29, 23, 7) {real, imag} */,
  {32'hc005a849, 32'hc04b53a4} /* (29, 23, 6) {real, imag} */,
  {32'hc03c05e2, 32'h3ffaae70} /* (29, 23, 5) {real, imag} */,
  {32'h3fb3ee88, 32'hc1583c04} /* (29, 23, 4) {real, imag} */,
  {32'hbf7fd6f8, 32'hc0ce00f6} /* (29, 23, 3) {real, imag} */,
  {32'hc11f8fda, 32'h3fe29bbc} /* (29, 23, 2) {real, imag} */,
  {32'hc13fc227, 32'h40aab7d0} /* (29, 23, 1) {real, imag} */,
  {32'hc0a82066, 32'h411f73fc} /* (29, 23, 0) {real, imag} */,
  {32'hc0cf8e07, 32'h404026ae} /* (29, 22, 31) {real, imag} */,
  {32'hc1390f06, 32'hbff7ed00} /* (29, 22, 30) {real, imag} */,
  {32'hc11e666c, 32'h409b7a54} /* (29, 22, 29) {real, imag} */,
  {32'h4000fe23, 32'h41056402} /* (29, 22, 28) {real, imag} */,
  {32'h3e62fc80, 32'hbfd092fc} /* (29, 22, 27) {real, imag} */,
  {32'hc15b6690, 32'h40f89492} /* (29, 22, 26) {real, imag} */,
  {32'hc12d022e, 32'h4149d2d0} /* (29, 22, 25) {real, imag} */,
  {32'hc00b1360, 32'hc0d58ae9} /* (29, 22, 24) {real, imag} */,
  {32'hc0ebe045, 32'hc0278464} /* (29, 22, 23) {real, imag} */,
  {32'hc0004ec4, 32'h4116baa7} /* (29, 22, 22) {real, imag} */,
  {32'h40567dd0, 32'h41644cdf} /* (29, 22, 21) {real, imag} */,
  {32'h3db99100, 32'h4138eaca} /* (29, 22, 20) {real, imag} */,
  {32'h40a94107, 32'h4044f38a} /* (29, 22, 19) {real, imag} */,
  {32'hc01edd80, 32'hbfc94e04} /* (29, 22, 18) {real, imag} */,
  {32'h4061e806, 32'h4127eae4} /* (29, 22, 17) {real, imag} */,
  {32'h40c95cc8, 32'h4008194a} /* (29, 22, 16) {real, imag} */,
  {32'h3fdd1766, 32'hc11980de} /* (29, 22, 15) {real, imag} */,
  {32'h40d63d3b, 32'h410a5b2e} /* (29, 22, 14) {real, imag} */,
  {32'h40e3fe3f, 32'h4107b940} /* (29, 22, 13) {real, imag} */,
  {32'h40df0218, 32'h4033f724} /* (29, 22, 12) {real, imag} */,
  {32'hc0b38c3c, 32'h40cac6fe} /* (29, 22, 11) {real, imag} */,
  {32'hc0d03b33, 32'h41b30e6c} /* (29, 22, 10) {real, imag} */,
  {32'hc0be28c7, 32'h418aa63e} /* (29, 22, 9) {real, imag} */,
  {32'hc143301b, 32'h41216592} /* (29, 22, 8) {real, imag} */,
  {32'hc0878703, 32'h41483d3a} /* (29, 22, 7) {real, imag} */,
  {32'hc0833f33, 32'h4184b7cf} /* (29, 22, 6) {real, imag} */,
  {32'hc17926f7, 32'h41399390} /* (29, 22, 5) {real, imag} */,
  {32'hc06e6fb4, 32'h413c09d0} /* (29, 22, 4) {real, imag} */,
  {32'hc0a4a4f0, 32'hc0e9ce25} /* (29, 22, 3) {real, imag} */,
  {32'h4064150f, 32'hc1135ab0} /* (29, 22, 2) {real, imag} */,
  {32'h4144bfef, 32'h40cb9238} /* (29, 22, 1) {real, imag} */,
  {32'h4019105b, 32'h410c2f02} /* (29, 22, 0) {real, imag} */,
  {32'h3df687c0, 32'h3f40b2c8} /* (29, 21, 31) {real, imag} */,
  {32'h40aaf11d, 32'h404c91b4} /* (29, 21, 30) {real, imag} */,
  {32'hbfdc7802, 32'hc0b749d4} /* (29, 21, 29) {real, imag} */,
  {32'h4106ea10, 32'hc09ab5d0} /* (29, 21, 28) {real, imag} */,
  {32'h41040f89, 32'h40245a5e} /* (29, 21, 27) {real, imag} */,
  {32'h40bebe7a, 32'h3ff7ae44} /* (29, 21, 26) {real, imag} */,
  {32'h4149081c, 32'hbff2bb54} /* (29, 21, 25) {real, imag} */,
  {32'h414dbebf, 32'h3f5a0558} /* (29, 21, 24) {real, imag} */,
  {32'h412d18b2, 32'hc07a15dc} /* (29, 21, 23) {real, imag} */,
  {32'h3fefe696, 32'h40be6d4c} /* (29, 21, 22) {real, imag} */,
  {32'hbf72d3e8, 32'h412a65af} /* (29, 21, 21) {real, imag} */,
  {32'hc104ce94, 32'hc020dd2f} /* (29, 21, 20) {real, imag} */,
  {32'hc0e89812, 32'hc0c146c2} /* (29, 21, 19) {real, imag} */,
  {32'hc047887a, 32'hbfc82128} /* (29, 21, 18) {real, imag} */,
  {32'hc13cef7f, 32'h410a149d} /* (29, 21, 17) {real, imag} */,
  {32'hc15316f0, 32'h41045e07} /* (29, 21, 16) {real, imag} */,
  {32'hc11054ee, 32'h3fd4568c} /* (29, 21, 15) {real, imag} */,
  {32'hc10f9d02, 32'hc0f87919} /* (29, 21, 14) {real, imag} */,
  {32'hc10644de, 32'hc0b092e3} /* (29, 21, 13) {real, imag} */,
  {32'h40344c36, 32'h3fb79bba} /* (29, 21, 12) {real, imag} */,
  {32'hc05d313d, 32'hc0a0316a} /* (29, 21, 11) {real, imag} */,
  {32'hc0864eaf, 32'hc016e4fe} /* (29, 21, 10) {real, imag} */,
  {32'h3f3392d0, 32'h404bf63a} /* (29, 21, 9) {real, imag} */,
  {32'h400f5a6e, 32'h410885fc} /* (29, 21, 8) {real, imag} */,
  {32'h404bdf72, 32'h41642397} /* (29, 21, 7) {real, imag} */,
  {32'h4076daf6, 32'h3f98e2b0} /* (29, 21, 6) {real, imag} */,
  {32'h40f74596, 32'hbfac7a24} /* (29, 21, 5) {real, imag} */,
  {32'h40062004, 32'h412bb0b5} /* (29, 21, 4) {real, imag} */,
  {32'h41802fe2, 32'h3f7c3114} /* (29, 21, 3) {real, imag} */,
  {32'h413b7fc8, 32'hc1811511} /* (29, 21, 2) {real, imag} */,
  {32'h3fffa576, 32'hc0cdaa30} /* (29, 21, 1) {real, imag} */,
  {32'hbfe1c724, 32'h3faec763} /* (29, 21, 0) {real, imag} */,
  {32'h3f1612f0, 32'h40f1d736} /* (29, 20, 31) {real, imag} */,
  {32'h3fd1b39e, 32'h40d32595} /* (29, 20, 30) {real, imag} */,
  {32'h40c65fab, 32'h3fa1bfcc} /* (29, 20, 29) {real, imag} */,
  {32'hc006bb32, 32'h4067b0ba} /* (29, 20, 28) {real, imag} */,
  {32'hc0cfb836, 32'hc008fb92} /* (29, 20, 27) {real, imag} */,
  {32'hc008612a, 32'hc12e9f1c} /* (29, 20, 26) {real, imag} */,
  {32'hc10023ca, 32'hc0fa2194} /* (29, 20, 25) {real, imag} */,
  {32'h40316316, 32'hbf8e0068} /* (29, 20, 24) {real, imag} */,
  {32'h3ff3e378, 32'h3fae1222} /* (29, 20, 23) {real, imag} */,
  {32'hc01e3ee6, 32'h40de411b} /* (29, 20, 22) {real, imag} */,
  {32'hc1250960, 32'hbf9d995c} /* (29, 20, 21) {real, imag} */,
  {32'hc16dac56, 32'h40cbe714} /* (29, 20, 20) {real, imag} */,
  {32'hc0c2266e, 32'h40425b86} /* (29, 20, 19) {real, imag} */,
  {32'h40c8471c, 32'hc0126ff8} /* (29, 20, 18) {real, imag} */,
  {32'h41008fee, 32'hc109c606} /* (29, 20, 17) {real, imag} */,
  {32'h40e64523, 32'hc0708638} /* (29, 20, 16) {real, imag} */,
  {32'h40445888, 32'hbf2dc958} /* (29, 20, 15) {real, imag} */,
  {32'h3fc3d744, 32'h3fbe0bb0} /* (29, 20, 14) {real, imag} */,
  {32'hbf963e3c, 32'h408729d1} /* (29, 20, 13) {real, imag} */,
  {32'hc012820e, 32'h4058c521} /* (29, 20, 12) {real, imag} */,
  {32'h407dc472, 32'hc1258587} /* (29, 20, 11) {real, imag} */,
  {32'h40f45b57, 32'hc0e25811} /* (29, 20, 10) {real, imag} */,
  {32'h3fa47342, 32'h3fee70b4} /* (29, 20, 9) {real, imag} */,
  {32'hc0d781c6, 32'h3fa66c74} /* (29, 20, 8) {real, imag} */,
  {32'h3ff3e326, 32'h400fe6b8} /* (29, 20, 7) {real, imag} */,
  {32'hbc9f0e80, 32'hc0214803} /* (29, 20, 6) {real, imag} */,
  {32'h405e4122, 32'h3f0052c8} /* (29, 20, 5) {real, imag} */,
  {32'h4014e6e6, 32'h3f1d733b} /* (29, 20, 4) {real, imag} */,
  {32'h3e134810, 32'hc0607f16} /* (29, 20, 3) {real, imag} */,
  {32'h40e12b3c, 32'hc02d4552} /* (29, 20, 2) {real, imag} */,
  {32'h3c2dd800, 32'h3f08e380} /* (29, 20, 1) {real, imag} */,
  {32'h3fbe3bdd, 32'h3ffb1d86} /* (29, 20, 0) {real, imag} */,
  {32'h3f4e9ba6, 32'hbe4fa9b8} /* (29, 19, 31) {real, imag} */,
  {32'hc00bca6c, 32'h40494cbe} /* (29, 19, 30) {real, imag} */,
  {32'hc0a9d9f0, 32'h4105a1c0} /* (29, 19, 29) {real, imag} */,
  {32'hc035cc31, 32'h40759ad2} /* (29, 19, 28) {real, imag} */,
  {32'hbfef34fe, 32'h4050d9da} /* (29, 19, 27) {real, imag} */,
  {32'hbe61c410, 32'hbf7f92bc} /* (29, 19, 26) {real, imag} */,
  {32'h3f3517a8, 32'hc032fe35} /* (29, 19, 25) {real, imag} */,
  {32'hc08cae8d, 32'h3fdd7fb8} /* (29, 19, 24) {real, imag} */,
  {32'h3d001700, 32'hc0e7a626} /* (29, 19, 23) {real, imag} */,
  {32'h3f1cd974, 32'hc1206496} /* (29, 19, 22) {real, imag} */,
  {32'h3f4ef168, 32'hc080e41a} /* (29, 19, 21) {real, imag} */,
  {32'h3cbb4c00, 32'hc0e13b94} /* (29, 19, 20) {real, imag} */,
  {32'hbf4d1fb0, 32'hc0a190b6} /* (29, 19, 19) {real, imag} */,
  {32'hc0111eba, 32'hbfd8df44} /* (29, 19, 18) {real, imag} */,
  {32'hc0b329bc, 32'hc02606df} /* (29, 19, 17) {real, imag} */,
  {32'h3fbc6628, 32'hc03e6c62} /* (29, 19, 16) {real, imag} */,
  {32'h40c99a2a, 32'hc0a20a3e} /* (29, 19, 15) {real, imag} */,
  {32'h3fa43ec0, 32'hc006ad7c} /* (29, 19, 14) {real, imag} */,
  {32'hbe90e108, 32'h40c7e564} /* (29, 19, 13) {real, imag} */,
  {32'hc04746d8, 32'h410de658} /* (29, 19, 12) {real, imag} */,
  {32'hc122558e, 32'h406afbd7} /* (29, 19, 11) {real, imag} */,
  {32'hbfe48530, 32'hc099bbf9} /* (29, 19, 10) {real, imag} */,
  {32'h4005f41c, 32'h3f8a6438} /* (29, 19, 9) {real, imag} */,
  {32'h3f30da00, 32'hc02e1980} /* (29, 19, 8) {real, imag} */,
  {32'h3fc7f0a8, 32'h3e7ced20} /* (29, 19, 7) {real, imag} */,
  {32'h40944950, 32'h400941cf} /* (29, 19, 6) {real, imag} */,
  {32'h3f9f9da4, 32'hc0a70625} /* (29, 19, 5) {real, imag} */,
  {32'h40b5e42a, 32'hc0f78d2f} /* (29, 19, 4) {real, imag} */,
  {32'hc05f8b4b, 32'hc0afa8d8} /* (29, 19, 3) {real, imag} */,
  {32'hc0c72b36, 32'hc01eb571} /* (29, 19, 2) {real, imag} */,
  {32'hbeaa7270, 32'h4005951a} /* (29, 19, 1) {real, imag} */,
  {32'h3ff12f62, 32'hbf731c20} /* (29, 19, 0) {real, imag} */,
  {32'hc08ed8f4, 32'hbff7b40c} /* (29, 18, 31) {real, imag} */,
  {32'hc0498736, 32'hbf5c4d20} /* (29, 18, 30) {real, imag} */,
  {32'h400acbac, 32'hc0b4dea2} /* (29, 18, 29) {real, imag} */,
  {32'h405e58e8, 32'hc090d9eb} /* (29, 18, 28) {real, imag} */,
  {32'h409f7ac9, 32'hbfcafb7c} /* (29, 18, 27) {real, imag} */,
  {32'h40382b3a, 32'hbfc54e80} /* (29, 18, 26) {real, imag} */,
  {32'h3fef1b24, 32'h3f648e60} /* (29, 18, 25) {real, imag} */,
  {32'h403da43c, 32'h40407c54} /* (29, 18, 24) {real, imag} */,
  {32'h40ad0195, 32'h3ebc2b60} /* (29, 18, 23) {real, imag} */,
  {32'h40c56bba, 32'hbf1de388} /* (29, 18, 22) {real, imag} */,
  {32'h40070b6c, 32'h40ec4c2d} /* (29, 18, 21) {real, imag} */,
  {32'hc111816c, 32'h3fa7d3a2} /* (29, 18, 20) {real, imag} */,
  {32'hc0babe08, 32'hc06a90c0} /* (29, 18, 19) {real, imag} */,
  {32'hc0812052, 32'hc05e7c00} /* (29, 18, 18) {real, imag} */,
  {32'hc0a61442, 32'h405cd720} /* (29, 18, 17) {real, imag} */,
  {32'h3f9a3aa8, 32'h408ede8b} /* (29, 18, 16) {real, imag} */,
  {32'hc051c6fb, 32'hc0082f9d} /* (29, 18, 15) {real, imag} */,
  {32'hc0e8263f, 32'h3f1b1058} /* (29, 18, 14) {real, imag} */,
  {32'hc0a0b970, 32'hbf58cc18} /* (29, 18, 13) {real, imag} */,
  {32'hc0422938, 32'hbf853dd0} /* (29, 18, 12) {real, imag} */,
  {32'hc042f123, 32'h40958947} /* (29, 18, 11) {real, imag} */,
  {32'h3fa7e430, 32'h40936ed8} /* (29, 18, 10) {real, imag} */,
  {32'h41056c8f, 32'h3f993d1c} /* (29, 18, 9) {real, imag} */,
  {32'h4104b348, 32'h4022a5ef} /* (29, 18, 8) {real, imag} */,
  {32'h3fb95fe8, 32'h403e9c2f} /* (29, 18, 7) {real, imag} */,
  {32'h3feabec0, 32'h40ecf771} /* (29, 18, 6) {real, imag} */,
  {32'hbfec11b4, 32'h3f681008} /* (29, 18, 5) {real, imag} */,
  {32'h4092e896, 32'hc0867bef} /* (29, 18, 4) {real, imag} */,
  {32'h40ba2772, 32'hc0c4f3c5} /* (29, 18, 3) {real, imag} */,
  {32'h3eeef560, 32'h402f9f0b} /* (29, 18, 2) {real, imag} */,
  {32'h40488a7b, 32'h40ad462a} /* (29, 18, 1) {real, imag} */,
  {32'hc0148504, 32'hbec63a7c} /* (29, 18, 0) {real, imag} */,
  {32'h401325e3, 32'hbfd4261e} /* (29, 17, 31) {real, imag} */,
  {32'h4005cdc6, 32'hc04a0482} /* (29, 17, 30) {real, imag} */,
  {32'h3fddda31, 32'h3eddca80} /* (29, 17, 29) {real, imag} */,
  {32'h3fb4fc37, 32'hbe61fec0} /* (29, 17, 28) {real, imag} */,
  {32'hc05c2240, 32'h3fd2f5a8} /* (29, 17, 27) {real, imag} */,
  {32'hc09280bc, 32'h4022e1c0} /* (29, 17, 26) {real, imag} */,
  {32'hc056f414, 32'h3f91fc10} /* (29, 17, 25) {real, imag} */,
  {32'hc06d9bbb, 32'hbe1410a0} /* (29, 17, 24) {real, imag} */,
  {32'hc0b65c59, 32'hc09dd92d} /* (29, 17, 23) {real, imag} */,
  {32'hc0e2d45e, 32'h40070bbc} /* (29, 17, 22) {real, imag} */,
  {32'h3cc38d00, 32'h3f16bc66} /* (29, 17, 21) {real, imag} */,
  {32'h40010b90, 32'hc023309b} /* (29, 17, 20) {real, imag} */,
  {32'h4017abb0, 32'h3f69e4c0} /* (29, 17, 19) {real, imag} */,
  {32'h410e9f10, 32'hc0619ea0} /* (29, 17, 18) {real, imag} */,
  {32'h41218ab8, 32'hc02d5f04} /* (29, 17, 17) {real, imag} */,
  {32'h408326c6, 32'h40a6f724} /* (29, 17, 16) {real, imag} */,
  {32'h4108c21c, 32'h40d249ec} /* (29, 17, 15) {real, imag} */,
  {32'h40cd2cf0, 32'hbf400494} /* (29, 17, 14) {real, imag} */,
  {32'h3eb055f8, 32'hbe931c08} /* (29, 17, 13) {real, imag} */,
  {32'hc0016d34, 32'hc023f658} /* (29, 17, 12) {real, imag} */,
  {32'h4083745b, 32'hc03f20b8} /* (29, 17, 11) {real, imag} */,
  {32'hbef37a80, 32'h408d1fb3} /* (29, 17, 10) {real, imag} */,
  {32'hc08b8350, 32'h40929610} /* (29, 17, 9) {real, imag} */,
  {32'hc0eb7ef6, 32'h3f9338b0} /* (29, 17, 8) {real, imag} */,
  {32'hc120b96b, 32'h3fa5b478} /* (29, 17, 7) {real, imag} */,
  {32'hc097ecb2, 32'h3ebd5400} /* (29, 17, 6) {real, imag} */,
  {32'h3eab0f40, 32'hbfbec10c} /* (29, 17, 5) {real, imag} */,
  {32'hc07fb7f4, 32'hc04a2bd8} /* (29, 17, 4) {real, imag} */,
  {32'h40022340, 32'hc02f49e8} /* (29, 17, 3) {real, imag} */,
  {32'h40c92651, 32'hc05a7208} /* (29, 17, 2) {real, imag} */,
  {32'hbf4e075c, 32'hc0bb0765} /* (29, 17, 1) {real, imag} */,
  {32'hc023ddde, 32'hc09b2a66} /* (29, 17, 0) {real, imag} */,
  {32'hbe912f00, 32'hbf293848} /* (29, 16, 31) {real, imag} */,
  {32'h3f5ccca0, 32'hbeb70180} /* (29, 16, 30) {real, imag} */,
  {32'hc04b558a, 32'hbfd401e0} /* (29, 16, 29) {real, imag} */,
  {32'h3f1b2ec0, 32'h401ef058} /* (29, 16, 28) {real, imag} */,
  {32'hc010df60, 32'h40694400} /* (29, 16, 27) {real, imag} */,
  {32'hbf0a7f34, 32'h4072e8f0} /* (29, 16, 26) {real, imag} */,
  {32'h4090f5b4, 32'h40def6f8} /* (29, 16, 25) {real, imag} */,
  {32'h3faf674b, 32'h40a3c1f8} /* (29, 16, 24) {real, imag} */,
  {32'hbff7a770, 32'h3f7e1240} /* (29, 16, 23) {real, imag} */,
  {32'hc0a5845c, 32'hc071b8c0} /* (29, 16, 22) {real, imag} */,
  {32'hbf60d220, 32'hbf1aa940} /* (29, 16, 21) {real, imag} */,
  {32'h4074736a, 32'hc025af58} /* (29, 16, 20) {real, imag} */,
  {32'h40787e24, 32'hc05c9340} /* (29, 16, 19) {real, imag} */,
  {32'hbffc29c8, 32'h3e792f80} /* (29, 16, 18) {real, imag} */,
  {32'h3f7af190, 32'h403943b0} /* (29, 16, 17) {real, imag} */,
  {32'h40867fea, 32'h40a0b692} /* (29, 16, 16) {real, imag} */,
  {32'h3f900386, 32'h4085f13c} /* (29, 16, 15) {real, imag} */,
  {32'h3f6a5000, 32'h3f704680} /* (29, 16, 14) {real, imag} */,
  {32'hbe727840, 32'h3f2ac040} /* (29, 16, 13) {real, imag} */,
  {32'h4039d426, 32'h404aabe0} /* (29, 16, 12) {real, imag} */,
  {32'h40abd032, 32'hbf86b720} /* (29, 16, 11) {real, imag} */,
  {32'h3fbd2550, 32'hc00e54d8} /* (29, 16, 10) {real, imag} */,
  {32'hc04f57e2, 32'h3f9f2e98} /* (29, 16, 9) {real, imag} */,
  {32'hbfd20f48, 32'h4004ab79} /* (29, 16, 8) {real, imag} */,
  {32'h3f9370ef, 32'hbef56b00} /* (29, 16, 7) {real, imag} */,
  {32'hc0313708, 32'h3f818248} /* (29, 16, 6) {real, imag} */,
  {32'h401707f0, 32'h3ed25940} /* (29, 16, 5) {real, imag} */,
  {32'h40bd247a, 32'h409eb04c} /* (29, 16, 4) {real, imag} */,
  {32'h3f6a2e40, 32'h406bd990} /* (29, 16, 3) {real, imag} */,
  {32'h3fe4b6b4, 32'h4078c928} /* (29, 16, 2) {real, imag} */,
  {32'h40159386, 32'h40a9d368} /* (29, 16, 1) {real, imag} */,
  {32'h3f034500, 32'h3fe579f8} /* (29, 16, 0) {real, imag} */,
  {32'h4012ee2d, 32'h3feef05e} /* (29, 15, 31) {real, imag} */,
  {32'hc0809743, 32'hc040a5fe} /* (29, 15, 30) {real, imag} */,
  {32'hbea62084, 32'hc080ee48} /* (29, 15, 29) {real, imag} */,
  {32'h3f466cd2, 32'h3fe2e318} /* (29, 15, 28) {real, imag} */,
  {32'h409f22d8, 32'h3fd9cfd8} /* (29, 15, 27) {real, imag} */,
  {32'h3fcb77d0, 32'h40214ba0} /* (29, 15, 26) {real, imag} */,
  {32'hc040366c, 32'h40b263cc} /* (29, 15, 25) {real, imag} */,
  {32'hc06d0525, 32'h408dc565} /* (29, 15, 24) {real, imag} */,
  {32'hc08ea357, 32'h4093d7ad} /* (29, 15, 23) {real, imag} */,
  {32'hc0e0a1ae, 32'hbf64e7f0} /* (29, 15, 22) {real, imag} */,
  {32'hc09aaf81, 32'hbd934d30} /* (29, 15, 21) {real, imag} */,
  {32'hc089c5e8, 32'hc06bed15} /* (29, 15, 20) {real, imag} */,
  {32'hc09361b0, 32'hc079b8e0} /* (29, 15, 19) {real, imag} */,
  {32'hc0879a70, 32'hbeff3c80} /* (29, 15, 18) {real, imag} */,
  {32'hc0bdc2d0, 32'hc00c2edc} /* (29, 15, 17) {real, imag} */,
  {32'hc0e3fe7e, 32'h3f8f00b0} /* (29, 15, 16) {real, imag} */,
  {32'hbffa12ec, 32'h4025ab69} /* (29, 15, 15) {real, imag} */,
  {32'hbfb2b8a0, 32'hbf7cb0ec} /* (29, 15, 14) {real, imag} */,
  {32'hbd5407c0, 32'hc0cfcec0} /* (29, 15, 13) {real, imag} */,
  {32'hc0c2a656, 32'hc04d5f68} /* (29, 15, 12) {real, imag} */,
  {32'hc09fe6c7, 32'hc03f0028} /* (29, 15, 11) {real, imag} */,
  {32'hc04203b0, 32'hc0606de6} /* (29, 15, 10) {real, imag} */,
  {32'hbfd5fb3e, 32'hbfa19d40} /* (29, 15, 9) {real, imag} */,
  {32'h3ebc9fa0, 32'hc0467258} /* (29, 15, 8) {real, imag} */,
  {32'h40f307ca, 32'hc068023c} /* (29, 15, 7) {real, imag} */,
  {32'h40aa712a, 32'hbf6c07c0} /* (29, 15, 6) {real, imag} */,
  {32'h4066ef90, 32'hc02627ba} /* (29, 15, 5) {real, imag} */,
  {32'h40f2687a, 32'h3f181360} /* (29, 15, 4) {real, imag} */,
  {32'hbfb864c0, 32'h403730e8} /* (29, 15, 3) {real, imag} */,
  {32'hc04d1bb2, 32'hc0510d18} /* (29, 15, 2) {real, imag} */,
  {32'hbf5d1f24, 32'hc0184cd6} /* (29, 15, 1) {real, imag} */,
  {32'hbf38d1ba, 32'h3f4712f4} /* (29, 15, 0) {real, imag} */,
  {32'hc0bf158c, 32'hc0ae247d} /* (29, 14, 31) {real, imag} */,
  {32'hc10167e2, 32'hbfe35270} /* (29, 14, 30) {real, imag} */,
  {32'hc12146a8, 32'hbf0d7d30} /* (29, 14, 29) {real, imag} */,
  {32'hc02c6570, 32'hc080e19d} /* (29, 14, 28) {real, imag} */,
  {32'hbea0ee70, 32'hbf3b3e48} /* (29, 14, 27) {real, imag} */,
  {32'hc01035a6, 32'h3fbeac00} /* (29, 14, 26) {real, imag} */,
  {32'hc0a35167, 32'h4042cce8} /* (29, 14, 25) {real, imag} */,
  {32'hc08bd3fa, 32'h3f8fc618} /* (29, 14, 24) {real, imag} */,
  {32'hc067bd42, 32'h3f7850d0} /* (29, 14, 23) {real, imag} */,
  {32'hc04dfc74, 32'h40950919} /* (29, 14, 22) {real, imag} */,
  {32'hc126b36f, 32'h40876543} /* (29, 14, 21) {real, imag} */,
  {32'hbf5935c0, 32'hc06b3571} /* (29, 14, 20) {real, imag} */,
  {32'h40e7ca78, 32'hc11e1ba0} /* (29, 14, 19) {real, imag} */,
  {32'hbe7cdc40, 32'hc0ae4010} /* (29, 14, 18) {real, imag} */,
  {32'hbe20ab40, 32'hbfc79bc0} /* (29, 14, 17) {real, imag} */,
  {32'h3fcecd78, 32'hc0fce143} /* (29, 14, 16) {real, imag} */,
  {32'hbd28df40, 32'hc0aeb122} /* (29, 14, 15) {real, imag} */,
  {32'h4055269e, 32'hbf463b58} /* (29, 14, 14) {real, imag} */,
  {32'h40b93fec, 32'h40191296} /* (29, 14, 13) {real, imag} */,
  {32'h409767e0, 32'hc008ebb8} /* (29, 14, 12) {real, imag} */,
  {32'hbff4e5a6, 32'hc0a0e2ef} /* (29, 14, 11) {real, imag} */,
  {32'h3f87dfa0, 32'h40ac308c} /* (29, 14, 10) {real, imag} */,
  {32'h3ddb6880, 32'h40bd5029} /* (29, 14, 9) {real, imag} */,
  {32'h40347340, 32'hbf8a4b5e} /* (29, 14, 8) {real, imag} */,
  {32'hc02375fc, 32'h408c2ea8} /* (29, 14, 7) {real, imag} */,
  {32'hc06bef70, 32'h40f92d6f} /* (29, 14, 6) {real, imag} */,
  {32'hbec65570, 32'hc0809c91} /* (29, 14, 5) {real, imag} */,
  {32'hc02af514, 32'hc04734e2} /* (29, 14, 4) {real, imag} */,
  {32'hc052c34b, 32'h400f3c0a} /* (29, 14, 3) {real, imag} */,
  {32'hc0fb5c98, 32'hbf6130ac} /* (29, 14, 2) {real, imag} */,
  {32'hc12a895d, 32'hbf609354} /* (29, 14, 1) {real, imag} */,
  {32'hc0e252b2, 32'h3ffbb64f} /* (29, 14, 0) {real, imag} */,
  {32'hbf5914ba, 32'h40013248} /* (29, 13, 31) {real, imag} */,
  {32'hbfd28bd8, 32'h400bdf22} /* (29, 13, 30) {real, imag} */,
  {32'h3fc57990, 32'h409bc5ff} /* (29, 13, 29) {real, imag} */,
  {32'h40876c36, 32'h40b3430d} /* (29, 13, 28) {real, imag} */,
  {32'hbf6cb104, 32'h4085b80b} /* (29, 13, 27) {real, imag} */,
  {32'h3fdf89ee, 32'hbfd54ff2} /* (29, 13, 26) {real, imag} */,
  {32'h41139d4e, 32'hc0225fdb} /* (29, 13, 25) {real, imag} */,
  {32'h4090b9b3, 32'h3fceeb88} /* (29, 13, 24) {real, imag} */,
  {32'hbfa43dd0, 32'h404df1bc} /* (29, 13, 23) {real, imag} */,
  {32'h4006659d, 32'hc02d2f72} /* (29, 13, 22) {real, imag} */,
  {32'h40af1cb9, 32'hc08e77d6} /* (29, 13, 21) {real, imag} */,
  {32'hbfc5a410, 32'hc082f5c0} /* (29, 13, 20) {real, imag} */,
  {32'hc1295453, 32'h407f2fa4} /* (29, 13, 19) {real, imag} */,
  {32'hc046016a, 32'h40cde11b} /* (29, 13, 18) {real, imag} */,
  {32'h3f51e7c0, 32'h3fc92e76} /* (29, 13, 17) {real, imag} */,
  {32'hc130b367, 32'h3f951c1c} /* (29, 13, 16) {real, imag} */,
  {32'hc131c703, 32'h3dc58760} /* (29, 13, 15) {real, imag} */,
  {32'h400f4ef8, 32'h3fc63038} /* (29, 13, 14) {real, imag} */,
  {32'hbf8e2eae, 32'h3edf9860} /* (29, 13, 13) {real, imag} */,
  {32'hc09fde08, 32'hc0cbf454} /* (29, 13, 12) {real, imag} */,
  {32'h3f329c68, 32'hbf80e322} /* (29, 13, 11) {real, imag} */,
  {32'h40447da8, 32'h3f0e9948} /* (29, 13, 10) {real, imag} */,
  {32'hc0564a74, 32'hbff1cbc8} /* (29, 13, 9) {real, imag} */,
  {32'hc0ed4624, 32'hc08b2578} /* (29, 13, 8) {real, imag} */,
  {32'hc04b90ac, 32'hc04a9c0a} /* (29, 13, 7) {real, imag} */,
  {32'hbfbfbb1e, 32'hc0987bf0} /* (29, 13, 6) {real, imag} */,
  {32'h3f5f9c38, 32'hc1291cb0} /* (29, 13, 5) {real, imag} */,
  {32'h406b33fc, 32'hc0e54751} /* (29, 13, 4) {real, imag} */,
  {32'h404aa205, 32'hc0961670} /* (29, 13, 3) {real, imag} */,
  {32'h40375f2d, 32'hc07c830d} /* (29, 13, 2) {real, imag} */,
  {32'h3e69dde0, 32'hc05cb42c} /* (29, 13, 1) {real, imag} */,
  {32'hc085bd72, 32'hc0e2d296} /* (29, 13, 0) {real, imag} */,
  {32'h3f383e88, 32'h3f1f0cf4} /* (29, 12, 31) {real, imag} */,
  {32'hbfeab158, 32'hc079068e} /* (29, 12, 30) {real, imag} */,
  {32'h3f872dd4, 32'hc04df0a6} /* (29, 12, 29) {real, imag} */,
  {32'hbfda926c, 32'hc0a86797} /* (29, 12, 28) {real, imag} */,
  {32'hbf085790, 32'h3f905d64} /* (29, 12, 27) {real, imag} */,
  {32'h40e8ad03, 32'hc00c56f6} /* (29, 12, 26) {real, imag} */,
  {32'h40c4cea4, 32'hc0f0f4d8} /* (29, 12, 25) {real, imag} */,
  {32'h40b656b9, 32'hc15383ad} /* (29, 12, 24) {real, imag} */,
  {32'h40b432f2, 32'hc064dd51} /* (29, 12, 23) {real, imag} */,
  {32'h4086a333, 32'h41122e12} /* (29, 12, 22) {real, imag} */,
  {32'h40854ec0, 32'h40bb5caf} /* (29, 12, 21) {real, imag} */,
  {32'h3ed81e80, 32'h4062af90} /* (29, 12, 20) {real, imag} */,
  {32'hbeaf1360, 32'h3f073c46} /* (29, 12, 19) {real, imag} */,
  {32'hbf84e2d2, 32'h41490664} /* (29, 12, 18) {real, imag} */,
  {32'hc0a9f0b7, 32'h415751fa} /* (29, 12, 17) {real, imag} */,
  {32'h40841385, 32'hbf960510} /* (29, 12, 16) {real, imag} */,
  {32'hbdc32310, 32'hc1094b9a} /* (29, 12, 15) {real, imag} */,
  {32'hc032e666, 32'h40a103d4} /* (29, 12, 14) {real, imag} */,
  {32'h40ea4cb5, 32'h40fd522d} /* (29, 12, 13) {real, imag} */,
  {32'h4123711c, 32'h3fdcd192} /* (29, 12, 12) {real, imag} */,
  {32'h4139ebaa, 32'hc02b37df} /* (29, 12, 11) {real, imag} */,
  {32'h3ff9094c, 32'h3f9d4cf4} /* (29, 12, 10) {real, imag} */,
  {32'h3fa1b562, 32'h40bb7471} /* (29, 12, 9) {real, imag} */,
  {32'h40293734, 32'h415ab9d0} /* (29, 12, 8) {real, imag} */,
  {32'h3eddb418, 32'h40b5affc} /* (29, 12, 7) {real, imag} */,
  {32'hc0bf5ac6, 32'hc013970d} /* (29, 12, 6) {real, imag} */,
  {32'hc108192e, 32'h400dae2e} /* (29, 12, 5) {real, imag} */,
  {32'hc020f6b4, 32'h3fb4ec22} /* (29, 12, 4) {real, imag} */,
  {32'hc081d8d0, 32'h4064f2ca} /* (29, 12, 3) {real, imag} */,
  {32'hc004df3d, 32'hc0d3f415} /* (29, 12, 2) {real, imag} */,
  {32'h406e25b8, 32'hc07ea170} /* (29, 12, 1) {real, imag} */,
  {32'h40aa172f, 32'h40c2f67e} /* (29, 12, 0) {real, imag} */,
  {32'hc00883c2, 32'hc0de2bf9} /* (29, 11, 31) {real, imag} */,
  {32'hc0a05a03, 32'hc11b3a83} /* (29, 11, 30) {real, imag} */,
  {32'h40fced40, 32'hc01a133c} /* (29, 11, 29) {real, imag} */,
  {32'hbf0addc0, 32'h4119b70e} /* (29, 11, 28) {real, imag} */,
  {32'hc1614e2f, 32'h413d80a0} /* (29, 11, 27) {real, imag} */,
  {32'hc0f7dd6a, 32'h40eb702b} /* (29, 11, 26) {real, imag} */,
  {32'hc12bdadc, 32'h4157103e} /* (29, 11, 25) {real, imag} */,
  {32'hc0dfdfa2, 32'h415400d6} /* (29, 11, 24) {real, imag} */,
  {32'hc0d51f31, 32'h4138bd1b} /* (29, 11, 23) {real, imag} */,
  {32'h40866a2c, 32'hc030aad8} /* (29, 11, 22) {real, imag} */,
  {32'hc03b68ba, 32'hc0e4ec76} /* (29, 11, 21) {real, imag} */,
  {32'h3ee37cf0, 32'h3e15ce90} /* (29, 11, 20) {real, imag} */,
  {32'hbfa8a6b8, 32'h40fd68de} /* (29, 11, 19) {real, imag} */,
  {32'hc06c8612, 32'h409b633a} /* (29, 11, 18) {real, imag} */,
  {32'h40332114, 32'hc0b50c1a} /* (29, 11, 17) {real, imag} */,
  {32'h40b452a8, 32'hc0ffc95e} /* (29, 11, 16) {real, imag} */,
  {32'h40398278, 32'hc158c978} /* (29, 11, 15) {real, imag} */,
  {32'hc061817e, 32'hc12be556} /* (29, 11, 14) {real, imag} */,
  {32'h412a2f9a, 32'h3f934a3c} /* (29, 11, 13) {real, imag} */,
  {32'h40fab607, 32'h408456ca} /* (29, 11, 12) {real, imag} */,
  {32'h40a392fe, 32'h4112f6d7} /* (29, 11, 11) {real, imag} */,
  {32'hc0730d7a, 32'h407542d6} /* (29, 11, 10) {real, imag} */,
  {32'hc14cbd84, 32'hc0e74bb3} /* (29, 11, 9) {real, imag} */,
  {32'hc0a7f937, 32'h3d3a6980} /* (29, 11, 8) {real, imag} */,
  {32'hc064c52a, 32'h3fb70be0} /* (29, 11, 7) {real, imag} */,
  {32'hc11897c2, 32'h400107a0} /* (29, 11, 6) {real, imag} */,
  {32'hc122caad, 32'h40def0e5} /* (29, 11, 5) {real, imag} */,
  {32'hc14ec6ad, 32'h41082d85} /* (29, 11, 4) {real, imag} */,
  {32'hc1782ab3, 32'h408ae232} /* (29, 11, 3) {real, imag} */,
  {32'hc09d19bd, 32'h403e74d0} /* (29, 11, 2) {real, imag} */,
  {32'h40835530, 32'h404ee700} /* (29, 11, 1) {real, imag} */,
  {32'h3f1641e8, 32'h40088bae} /* (29, 11, 0) {real, imag} */,
  {32'h41539164, 32'hc070b998} /* (29, 10, 31) {real, imag} */,
  {32'h41a36873, 32'hc0c2c334} /* (29, 10, 30) {real, imag} */,
  {32'h41be8156, 32'hc13ad11a} /* (29, 10, 29) {real, imag} */,
  {32'hc039231d, 32'hc0eb68f7} /* (29, 10, 28) {real, imag} */,
  {32'hc1857b61, 32'hc15598b8} /* (29, 10, 27) {real, imag} */,
  {32'hc19c9326, 32'hc0809dde} /* (29, 10, 26) {real, imag} */,
  {32'hc0975728, 32'h3f519238} /* (29, 10, 25) {real, imag} */,
  {32'h41296022, 32'hc05c4ca6} /* (29, 10, 24) {real, imag} */,
  {32'h410ac9c6, 32'h40db6916} /* (29, 10, 23) {real, imag} */,
  {32'h41837d14, 32'h4126f22f} /* (29, 10, 22) {real, imag} */,
  {32'h41bd41f6, 32'h40ddb022} /* (29, 10, 21) {real, imag} */,
  {32'h412f12ce, 32'h4142f8ca} /* (29, 10, 20) {real, imag} */,
  {32'hc0a3b139, 32'h410d660e} /* (29, 10, 19) {real, imag} */,
  {32'hc105d71d, 32'h3f3269c8} /* (29, 10, 18) {real, imag} */,
  {32'h407cc7ea, 32'h3f770e78} /* (29, 10, 17) {real, imag} */,
  {32'h40062e4d, 32'hc0f73be5} /* (29, 10, 16) {real, imag} */,
  {32'hc07d57a3, 32'h41128560} /* (29, 10, 15) {real, imag} */,
  {32'hc14e64c0, 32'h40c5ccb0} /* (29, 10, 14) {real, imag} */,
  {32'hc10ce7b8, 32'hc0d6d748} /* (29, 10, 13) {real, imag} */,
  {32'h405625b8, 32'hc11eb793} /* (29, 10, 12) {real, imag} */,
  {32'hc0ac4382, 32'hc128d523} /* (29, 10, 11) {real, imag} */,
  {32'hc081d2b3, 32'hc145d4f4} /* (29, 10, 10) {real, imag} */,
  {32'h408d3569, 32'hc1d8b178} /* (29, 10, 9) {real, imag} */,
  {32'h40b2ab7a, 32'hc14420de} /* (29, 10, 8) {real, imag} */,
  {32'h4169d372, 32'hc10dd964} /* (29, 10, 7) {real, imag} */,
  {32'h41207a00, 32'hc1173fe0} /* (29, 10, 6) {real, imag} */,
  {32'hbf6f91d0, 32'h40973ee9} /* (29, 10, 5) {real, imag} */,
  {32'hbf4840d0, 32'h40b6bda0} /* (29, 10, 4) {real, imag} */,
  {32'h405ff8b3, 32'h40f719a7} /* (29, 10, 3) {real, imag} */,
  {32'hc091d09e, 32'h402fd500} /* (29, 10, 2) {real, imag} */,
  {32'hc107b3bf, 32'h40d9e484} /* (29, 10, 1) {real, imag} */,
  {32'hbfe0ff92, 32'h3fec7bb8} /* (29, 10, 0) {real, imag} */,
  {32'hc0d6c3ee, 32'h411fc18a} /* (29, 9, 31) {real, imag} */,
  {32'h40dea8b6, 32'h3f4950b8} /* (29, 9, 30) {real, imag} */,
  {32'h40411ac0, 32'h402fdeb8} /* (29, 9, 29) {real, imag} */,
  {32'h40c92887, 32'h3f4c36e8} /* (29, 9, 28) {real, imag} */,
  {32'hbf99e2f8, 32'h40938e50} /* (29, 9, 27) {real, imag} */,
  {32'hc0c56bcd, 32'h40b51c78} /* (29, 9, 26) {real, imag} */,
  {32'hbf477020, 32'h3ea52ae8} /* (29, 9, 25) {real, imag} */,
  {32'hc0989cea, 32'hbfc955e8} /* (29, 9, 24) {real, imag} */,
  {32'hbf9c1bb4, 32'hc029a3d8} /* (29, 9, 23) {real, imag} */,
  {32'hbf005ab8, 32'h40bc9a83} /* (29, 9, 22) {real, imag} */,
  {32'hbfe8f480, 32'h414d2977} /* (29, 9, 21) {real, imag} */,
  {32'hc15388dc, 32'h41876cab} /* (29, 9, 20) {real, imag} */,
  {32'hc0039783, 32'h3fc23bf8} /* (29, 9, 19) {real, imag} */,
  {32'hbfcc202c, 32'hc122e88a} /* (29, 9, 18) {real, imag} */,
  {32'hc1117571, 32'h402332cc} /* (29, 9, 17) {real, imag} */,
  {32'hc10c7263, 32'h40b01b9a} /* (29, 9, 16) {real, imag} */,
  {32'h40974378, 32'h40b3c94d} /* (29, 9, 15) {real, imag} */,
  {32'hbf53d2b0, 32'h40a2d7c6} /* (29, 9, 14) {real, imag} */,
  {32'hbf9d9a54, 32'hc11a157e} /* (29, 9, 13) {real, imag} */,
  {32'hbf7d74b0, 32'hc140e230} /* (29, 9, 12) {real, imag} */,
  {32'h4092734e, 32'hc1bea00d} /* (29, 9, 11) {real, imag} */,
  {32'h41889bac, 32'hc17a4f46} /* (29, 9, 10) {real, imag} */,
  {32'h408597fa, 32'hc1091e6e} /* (29, 9, 9) {real, imag} */,
  {32'h40e5cd4f, 32'hc14d943c} /* (29, 9, 8) {real, imag} */,
  {32'h414eb605, 32'h40c92c7a} /* (29, 9, 7) {real, imag} */,
  {32'h410b7cef, 32'hc13d21ad} /* (29, 9, 6) {real, imag} */,
  {32'hbff71174, 32'hc178818e} /* (29, 9, 5) {real, imag} */,
  {32'hbe37ce00, 32'hc0e22298} /* (29, 9, 4) {real, imag} */,
  {32'h40faa0e5, 32'hc0e3b23e} /* (29, 9, 3) {real, imag} */,
  {32'h414b2500, 32'hc0e45ab1} /* (29, 9, 2) {real, imag} */,
  {32'h40ef8a12, 32'h4029b101} /* (29, 9, 1) {real, imag} */,
  {32'h3f4fa034, 32'hbdc35b40} /* (29, 9, 0) {real, imag} */,
  {32'hc13fcb04, 32'hbf7cd3e0} /* (29, 8, 31) {real, imag} */,
  {32'hc146460c, 32'hc124e052} /* (29, 8, 30) {real, imag} */,
  {32'hc003293e, 32'h416d16e8} /* (29, 8, 29) {real, imag} */,
  {32'h40d1adec, 32'h41bde3c2} /* (29, 8, 28) {real, imag} */,
  {32'h41823c8f, 32'h418d2504} /* (29, 8, 27) {real, imag} */,
  {32'h412b3269, 32'h40f800ee} /* (29, 8, 26) {real, imag} */,
  {32'hc0d1ce62, 32'h418f317a} /* (29, 8, 25) {real, imag} */,
  {32'hc18d5d3e, 32'h41ca6200} /* (29, 8, 24) {real, imag} */,
  {32'hc116e474, 32'h41935794} /* (29, 8, 23) {real, imag} */,
  {32'hc09d4b1c, 32'h414c560c} /* (29, 8, 22) {real, imag} */,
  {32'hc1606655, 32'h41379efb} /* (29, 8, 21) {real, imag} */,
  {32'hc1980ec0, 32'hc18b8c71} /* (29, 8, 20) {real, imag} */,
  {32'hc0be7418, 32'hc195fe91} /* (29, 8, 19) {real, imag} */,
  {32'hbfd1048c, 32'hc1a1e694} /* (29, 8, 18) {real, imag} */,
  {32'hc0fcb35a, 32'hc1335966} /* (29, 8, 17) {real, imag} */,
  {32'h415a7c3f, 32'hc11e8c60} /* (29, 8, 16) {real, imag} */,
  {32'h4200a23b, 32'hc0cb2f78} /* (29, 8, 15) {real, imag} */,
  {32'h419f74d6, 32'hc05a9e80} /* (29, 8, 14) {real, imag} */,
  {32'h4045f4bb, 32'hc07064e1} /* (29, 8, 13) {real, imag} */,
  {32'h416706a2, 32'hc0fb0c18} /* (29, 8, 12) {real, imag} */,
  {32'h40483478, 32'hc1bfc882} /* (29, 8, 11) {real, imag} */,
  {32'hbe8cae80, 32'hc0e58fb4} /* (29, 8, 10) {real, imag} */,
  {32'h41aae2b8, 32'hc0553bee} /* (29, 8, 9) {real, imag} */,
  {32'h4086dec4, 32'hc146c116} /* (29, 8, 8) {real, imag} */,
  {32'hc11b4159, 32'h3fb02215} /* (29, 8, 7) {real, imag} */,
  {32'hc0c4da00, 32'h41bd7d4c} /* (29, 8, 6) {real, imag} */,
  {32'hc11b8db7, 32'h412a2ada} /* (29, 8, 5) {real, imag} */,
  {32'hc125a118, 32'h41b4b82e} /* (29, 8, 4) {real, imag} */,
  {32'hc091455e, 32'h41621ecd} /* (29, 8, 3) {real, imag} */,
  {32'hc01ffdfa, 32'h41012713} /* (29, 8, 2) {real, imag} */,
  {32'h410cd107, 32'h4195307b} /* (29, 8, 1) {real, imag} */,
  {32'h3fb67714, 32'h418633cd} /* (29, 8, 0) {real, imag} */,
  {32'hc03330fb, 32'hc10e7844} /* (29, 7, 31) {real, imag} */,
  {32'hc047ac98, 32'hc10326f3} /* (29, 7, 30) {real, imag} */,
  {32'h3f097b10, 32'hc132f424} /* (29, 7, 29) {real, imag} */,
  {32'hc04d27e6, 32'hc0e43ffa} /* (29, 7, 28) {real, imag} */,
  {32'h402a7413, 32'hc13b0d4c} /* (29, 7, 27) {real, imag} */,
  {32'hc0c9227a, 32'hc194ece6} /* (29, 7, 26) {real, imag} */,
  {32'h3ffa7cce, 32'hc18fdb3e} /* (29, 7, 25) {real, imag} */,
  {32'h4199b198, 32'hbf6f8670} /* (29, 7, 24) {real, imag} */,
  {32'h4185d4c2, 32'h3e4cc340} /* (29, 7, 23) {real, imag} */,
  {32'h4000ba16, 32'hc03d476c} /* (29, 7, 22) {real, imag} */,
  {32'hc16cb408, 32'hc02db190} /* (29, 7, 21) {real, imag} */,
  {32'hc069dcda, 32'hc0a31e1e} /* (29, 7, 20) {real, imag} */,
  {32'hc06188f9, 32'h3ecbc860} /* (29, 7, 19) {real, imag} */,
  {32'hc114aafc, 32'hc150aca8} /* (29, 7, 18) {real, imag} */,
  {32'h40a7c358, 32'hc0c71ab6} /* (29, 7, 17) {real, imag} */,
  {32'hc1452ecd, 32'hbfca1120} /* (29, 7, 16) {real, imag} */,
  {32'hc0818c44, 32'h40935409} /* (29, 7, 15) {real, imag} */,
  {32'hc1048f9a, 32'hc092fdf4} /* (29, 7, 14) {real, imag} */,
  {32'hc1d03c53, 32'h41276c20} /* (29, 7, 13) {real, imag} */,
  {32'hc10c2bcc, 32'h40e5d0ef} /* (29, 7, 12) {real, imag} */,
  {32'h41b61bd8, 32'h40738cd2} /* (29, 7, 11) {real, imag} */,
  {32'h412b23aa, 32'h40b474a6} /* (29, 7, 10) {real, imag} */,
  {32'h4176b637, 32'h41979e05} /* (29, 7, 9) {real, imag} */,
  {32'h416c5416, 32'h415077be} /* (29, 7, 8) {real, imag} */,
  {32'h410ab180, 32'hc16d698b} /* (29, 7, 7) {real, imag} */,
  {32'hc04e8ac5, 32'hc1d46598} /* (29, 7, 6) {real, imag} */,
  {32'hc0e88ea3, 32'hc07e9ff4} /* (29, 7, 5) {real, imag} */,
  {32'hc072caf0, 32'hc0bd6cc1} /* (29, 7, 4) {real, imag} */,
  {32'h411a00fe, 32'hc1d8a7ac} /* (29, 7, 3) {real, imag} */,
  {32'h418e154b, 32'hc1f9e3c4} /* (29, 7, 2) {real, imag} */,
  {32'h41903968, 32'hc1bddcaf} /* (29, 7, 1) {real, imag} */,
  {32'h4059ac84, 32'hc0dda965} /* (29, 7, 0) {real, imag} */,
  {32'h413c9235, 32'h4053895c} /* (29, 6, 31) {real, imag} */,
  {32'h40bc2338, 32'h41c059f6} /* (29, 6, 30) {real, imag} */,
  {32'hc12115ba, 32'h41a83e65} /* (29, 6, 29) {real, imag} */,
  {32'h404f87d8, 32'h4153acd8} /* (29, 6, 28) {real, imag} */,
  {32'h3f7d7be0, 32'h40a151ff} /* (29, 6, 27) {real, imag} */,
  {32'hc08682b4, 32'hc0c636c6} /* (29, 6, 26) {real, imag} */,
  {32'h40c9740a, 32'h41840a71} /* (29, 6, 25) {real, imag} */,
  {32'h4161a52a, 32'hc008d036} /* (29, 6, 24) {real, imag} */,
  {32'h41436c2e, 32'hc18ed3ce} /* (29, 6, 23) {real, imag} */,
  {32'h4087bd6f, 32'h4023b5e0} /* (29, 6, 22) {real, imag} */,
  {32'h40f22f3c, 32'h4139a9b8} /* (29, 6, 21) {real, imag} */,
  {32'hbfe1191c, 32'h40241402} /* (29, 6, 20) {real, imag} */,
  {32'hc0561aa6, 32'hc117a2f6} /* (29, 6, 19) {real, imag} */,
  {32'hc031d114, 32'h4078a80e} /* (29, 6, 18) {real, imag} */,
  {32'hbf98bf54, 32'h418b5d38} /* (29, 6, 17) {real, imag} */,
  {32'h40e0989c, 32'hc04a6e7e} /* (29, 6, 16) {real, imag} */,
  {32'hc0b825e6, 32'hc199a2c2} /* (29, 6, 15) {real, imag} */,
  {32'hc155801b, 32'hc02ad0bc} /* (29, 6, 14) {real, imag} */,
  {32'h416f7f4a, 32'h4163d4bf} /* (29, 6, 13) {real, imag} */,
  {32'h4137d175, 32'h40ef6806} /* (29, 6, 12) {real, imag} */,
  {32'hc0334efe, 32'h40d8e442} /* (29, 6, 11) {real, imag} */,
  {32'hc119723a, 32'hc038d010} /* (29, 6, 10) {real, imag} */,
  {32'h40d89c5d, 32'hc11dae4d} /* (29, 6, 9) {real, imag} */,
  {32'h400e98a0, 32'h41186c4f} /* (29, 6, 8) {real, imag} */,
  {32'h3d2b26c0, 32'h40e34634} /* (29, 6, 7) {real, imag} */,
  {32'h4144b610, 32'hc10cb380} /* (29, 6, 6) {real, imag} */,
  {32'hc11006c6, 32'hc1139186} /* (29, 6, 5) {real, imag} */,
  {32'hc16c467d, 32'h4066812c} /* (29, 6, 4) {real, imag} */,
  {32'hc1168f64, 32'h412ed178} /* (29, 6, 3) {real, imag} */,
  {32'h4083f15b, 32'h41bb0006} /* (29, 6, 2) {real, imag} */,
  {32'h417f534b, 32'hc0692b18} /* (29, 6, 1) {real, imag} */,
  {32'h41159aab, 32'hc0c92ad9} /* (29, 6, 0) {real, imag} */,
  {32'hc029653e, 32'h416e8495} /* (29, 5, 31) {real, imag} */,
  {32'hc1440e38, 32'h4197e27a} /* (29, 5, 30) {real, imag} */,
  {32'hc14f5ad2, 32'h419417bf} /* (29, 5, 29) {real, imag} */,
  {32'h41517313, 32'h4193293a} /* (29, 5, 28) {real, imag} */,
  {32'h40818cd4, 32'h41964867} /* (29, 5, 27) {real, imag} */,
  {32'hc1550f24, 32'h418b8605} /* (29, 5, 26) {real, imag} */,
  {32'h3fa63870, 32'h4197dd73} /* (29, 5, 25) {real, imag} */,
  {32'h41113e00, 32'h415403ae} /* (29, 5, 24) {real, imag} */,
  {32'h40d41c85, 32'h41eb80a6} /* (29, 5, 23) {real, imag} */,
  {32'hc005597a, 32'h42246000} /* (29, 5, 22) {real, imag} */,
  {32'hc0fa9591, 32'h41fe01c4} /* (29, 5, 21) {real, imag} */,
  {32'h40a1a86b, 32'h410b5f98} /* (29, 5, 20) {real, imag} */,
  {32'h418d5efe, 32'hc13e63a0} /* (29, 5, 19) {real, imag} */,
  {32'h417591a4, 32'hc1a194df} /* (29, 5, 18) {real, imag} */,
  {32'h40801afc, 32'hc1849dbe} /* (29, 5, 17) {real, imag} */,
  {32'hc0e460c4, 32'h40f7f4c2} /* (29, 5, 16) {real, imag} */,
  {32'h41588c13, 32'h4097cc2a} /* (29, 5, 15) {real, imag} */,
  {32'h41034192, 32'h403ab8fc} /* (29, 5, 14) {real, imag} */,
  {32'h40dd1748, 32'hc1c37009} /* (29, 5, 13) {real, imag} */,
  {32'h4127c29a, 32'hc20e9f9b} /* (29, 5, 12) {real, imag} */,
  {32'h41558616, 32'hc1999497} /* (29, 5, 11) {real, imag} */,
  {32'h4170bcca, 32'h411829c9} /* (29, 5, 10) {real, imag} */,
  {32'h40ea1cb0, 32'h415060e8} /* (29, 5, 9) {real, imag} */,
  {32'h411449b6, 32'h41ee3f0d} /* (29, 5, 8) {real, imag} */,
  {32'h415ad828, 32'h42057b65} /* (29, 5, 7) {real, imag} */,
  {32'h4103ebbd, 32'h413baea3} /* (29, 5, 6) {real, imag} */,
  {32'h414810e0, 32'h40cffc77} /* (29, 5, 5) {real, imag} */,
  {32'hc0bf9aa6, 32'h4163b999} /* (29, 5, 4) {real, imag} */,
  {32'hc1428c7a, 32'h4216110a} /* (29, 5, 3) {real, imag} */,
  {32'hc128fc74, 32'h41eb2c2e} /* (29, 5, 2) {real, imag} */,
  {32'hc1032e9e, 32'h419ae5b8} /* (29, 5, 1) {real, imag} */,
  {32'hbf32c438, 32'h416b9e62} /* (29, 5, 0) {real, imag} */,
  {32'h411ae2b2, 32'hc07e10fb} /* (29, 4, 31) {real, imag} */,
  {32'h3eaf5e8a, 32'h403cd2a6} /* (29, 4, 30) {real, imag} */,
  {32'hc0e71aa5, 32'hc15b9198} /* (29, 4, 29) {real, imag} */,
  {32'h41cbf048, 32'hc19b7e34} /* (29, 4, 28) {real, imag} */,
  {32'h411ee156, 32'hc205d80e} /* (29, 4, 27) {real, imag} */,
  {32'hc0abda08, 32'hc1b4f616} /* (29, 4, 26) {real, imag} */,
  {32'h4129dc1e, 32'hc206a81f} /* (29, 4, 25) {real, imag} */,
  {32'h40f2139c, 32'hc1ee0ada} /* (29, 4, 24) {real, imag} */,
  {32'hc10ff599, 32'hc1b4f345} /* (29, 4, 23) {real, imag} */,
  {32'h3f8ceb20, 32'hc1686946} /* (29, 4, 22) {real, imag} */,
  {32'h40a1e0b8, 32'h41941e62} /* (29, 4, 21) {real, imag} */,
  {32'hc1d4904f, 32'h41f454c6} /* (29, 4, 20) {real, imag} */,
  {32'hc1cba013, 32'h41b4ef57} /* (29, 4, 19) {real, imag} */,
  {32'hc130e852, 32'h41af5964} /* (29, 4, 18) {real, imag} */,
  {32'hc18fb6d8, 32'h4208bfc2} /* (29, 4, 17) {real, imag} */,
  {32'hc16f4089, 32'h42363834} /* (29, 4, 16) {real, imag} */,
  {32'hc1146aa6, 32'h41cade76} /* (29, 4, 15) {real, imag} */,
  {32'hc18ae704, 32'h41fa83ee} /* (29, 4, 14) {real, imag} */,
  {32'hc10c9890, 32'h418db66b} /* (29, 4, 13) {real, imag} */,
  {32'hc024ab24, 32'h41308f50} /* (29, 4, 12) {real, imag} */,
  {32'h4080e7ff, 32'hc003ce26} /* (29, 4, 11) {real, imag} */,
  {32'h41fad6f4, 32'hc16b33ac} /* (29, 4, 10) {real, imag} */,
  {32'h42044bd0, 32'hc1245ef1} /* (29, 4, 9) {real, imag} */,
  {32'h41b34eff, 32'hc1a77631} /* (29, 4, 8) {real, imag} */,
  {32'h421125c5, 32'hc1651c9b} /* (29, 4, 7) {real, imag} */,
  {32'h423cfd13, 32'hc2060dba} /* (29, 4, 6) {real, imag} */,
  {32'h42270732, 32'hc22ad2a6} /* (29, 4, 5) {real, imag} */,
  {32'h409e8468, 32'hc1a34caa} /* (29, 4, 4) {real, imag} */,
  {32'hc055cd98, 32'h411f1e0c} /* (29, 4, 3) {real, imag} */,
  {32'h4151f5ce, 32'h41424152} /* (29, 4, 2) {real, imag} */,
  {32'h419f2590, 32'hc10439da} /* (29, 4, 1) {real, imag} */,
  {32'h415c8545, 32'hc1410f38} /* (29, 4, 0) {real, imag} */,
  {32'hc14a5846, 32'hc0ab71fc} /* (29, 3, 31) {real, imag} */,
  {32'hc1ff7696, 32'hc1073668} /* (29, 3, 30) {real, imag} */,
  {32'hc180b228, 32'h40925cfa} /* (29, 3, 29) {real, imag} */,
  {32'h3e540ba0, 32'h40983262} /* (29, 3, 28) {real, imag} */,
  {32'hc068fe14, 32'h420237fb} /* (29, 3, 27) {real, imag} */,
  {32'hc0f87d60, 32'h4200e84a} /* (29, 3, 26) {real, imag} */,
  {32'hc18b0eee, 32'h40bf7066} /* (29, 3, 25) {real, imag} */,
  {32'h409cc251, 32'h419d7fc8} /* (29, 3, 24) {real, imag} */,
  {32'h41461878, 32'h3ff67940} /* (29, 3, 23) {real, imag} */,
  {32'h414d60cd, 32'hc125ca9f} /* (29, 3, 22) {real, imag} */,
  {32'hc05771ae, 32'hc16fc0dc} /* (29, 3, 21) {real, imag} */,
  {32'hc230eb58, 32'h41e7a094} /* (29, 3, 20) {real, imag} */,
  {32'hc2543c1b, 32'h40bead74} /* (29, 3, 19) {real, imag} */,
  {32'hc1f9ff96, 32'hc19cb30e} /* (29, 3, 18) {real, imag} */,
  {32'hc233e51a, 32'h407f1e2a} /* (29, 3, 17) {real, imag} */,
  {32'hc2129be2, 32'h40f280a6} /* (29, 3, 16) {real, imag} */,
  {32'h3ff61b84, 32'hc1847742} /* (29, 3, 15) {real, imag} */,
  {32'h413835d4, 32'hbfc0f048} /* (29, 3, 14) {real, imag} */,
  {32'hc13df4f8, 32'h40e302da} /* (29, 3, 13) {real, imag} */,
  {32'hc1393b08, 32'h40d9a27a} /* (29, 3, 12) {real, imag} */,
  {32'h4105b10a, 32'h407be7e8} /* (29, 3, 11) {real, imag} */,
  {32'h424bc962, 32'hc137bc48} /* (29, 3, 10) {real, imag} */,
  {32'h4277450a, 32'h3f741f40} /* (29, 3, 9) {real, imag} */,
  {32'h42502fdb, 32'h4054aba4} /* (29, 3, 8) {real, imag} */,
  {32'h41d0f253, 32'hc08b4c4c} /* (29, 3, 7) {real, imag} */,
  {32'h41b818c1, 32'hc0350fcc} /* (29, 3, 6) {real, imag} */,
  {32'h41d14ca2, 32'h3fd0ecc8} /* (29, 3, 5) {real, imag} */,
  {32'h4147cea4, 32'h400e751e} /* (29, 3, 4) {real, imag} */,
  {32'h40ed6a9e, 32'hc03e6d40} /* (29, 3, 3) {real, imag} */,
  {32'h3ec18400, 32'hc128d44f} /* (29, 3, 2) {real, imag} */,
  {32'hc19077fa, 32'hbf52cff0} /* (29, 3, 1) {real, imag} */,
  {32'hc1554892, 32'h410e34f6} /* (29, 3, 0) {real, imag} */,
  {32'h40cf94b9, 32'h42598893} /* (29, 2, 31) {real, imag} */,
  {32'h417c571c, 32'h42b8785c} /* (29, 2, 30) {real, imag} */,
  {32'h3ed2d440, 32'h4270c099} /* (29, 2, 29) {real, imag} */,
  {32'hc20893a9, 32'h42083461} /* (29, 2, 28) {real, imag} */,
  {32'hc180b9a0, 32'h4243418e} /* (29, 2, 27) {real, imag} */,
  {32'h3ebd2540, 32'h4289bb29} /* (29, 2, 26) {real, imag} */,
  {32'h4014dff0, 32'h4281431b} /* (29, 2, 25) {real, imag} */,
  {32'h40a72d2c, 32'h4280eaa4} /* (29, 2, 24) {real, imag} */,
  {32'h41a386ac, 32'h428ffd6d} /* (29, 2, 23) {real, imag} */,
  {32'h421f5016, 32'h424b3eec} /* (29, 2, 22) {real, imag} */,
  {32'h4185b532, 32'hc16351e6} /* (29, 2, 21) {real, imag} */,
  {32'hc2311cec, 32'hc26c961b} /* (29, 2, 20) {real, imag} */,
  {32'hc279306f, 32'hc2264a3f} /* (29, 2, 19) {real, imag} */,
  {32'hc23dd895, 32'hc248b30c} /* (29, 2, 18) {real, imag} */,
  {32'hc25236b2, 32'hc284c3ed} /* (29, 2, 17) {real, imag} */,
  {32'hc21bce61, 32'hc23d5dae} /* (29, 2, 16) {real, imag} */,
  {32'hc16fb76d, 32'hc259ea3a} /* (29, 2, 15) {real, imag} */,
  {32'hc1a5b50a, 32'hc25cdc45} /* (29, 2, 14) {real, imag} */,
  {32'hc1b8e254, 32'hc2637b72} /* (29, 2, 13) {real, imag} */,
  {32'hc10a9ddd, 32'hc242eabe} /* (29, 2, 12) {real, imag} */,
  {32'h408e314a, 32'hc1d84077} /* (29, 2, 11) {real, imag} */,
  {32'h419f37a4, 32'h420913b6} /* (29, 2, 10) {real, imag} */,
  {32'h4211f7ba, 32'h428b4265} /* (29, 2, 9) {real, imag} */,
  {32'h4242aaee, 32'h42999cdf} /* (29, 2, 8) {real, imag} */,
  {32'h4247943b, 32'h42a68160} /* (29, 2, 7) {real, imag} */,
  {32'h423d0788, 32'h428f344b} /* (29, 2, 6) {real, imag} */,
  {32'h415a889a, 32'h42890675} /* (29, 2, 5) {real, imag} */,
  {32'h41a376b0, 32'h4272ec84} /* (29, 2, 4) {real, imag} */,
  {32'h4133f512, 32'h429887de} /* (29, 2, 3) {real, imag} */,
  {32'hbe000f80, 32'h4278e085} /* (29, 2, 2) {real, imag} */,
  {32'hc19453d0, 32'h423b7123} /* (29, 2, 1) {real, imag} */,
  {32'hc1d444be, 32'h41e4a59a} /* (29, 2, 0) {real, imag} */,
  {32'hc197be20, 32'hc2440d83} /* (29, 1, 31) {real, imag} */,
  {32'hc17ed0d0, 32'hc2956e72} /* (29, 1, 30) {real, imag} */,
  {32'hc183c77b, 32'hc2b349ca} /* (29, 1, 29) {real, imag} */,
  {32'hc1d78f84, 32'hc2e616f8} /* (29, 1, 28) {real, imag} */,
  {32'hc1b4ae41, 32'hc2d10e61} /* (29, 1, 27) {real, imag} */,
  {32'hc16c0812, 32'hc2af6ce7} /* (29, 1, 26) {real, imag} */,
  {32'hc1f12eb0, 32'hc2af8c94} /* (29, 1, 25) {real, imag} */,
  {32'hc1d142dc, 32'hc2b9acb9} /* (29, 1, 24) {real, imag} */,
  {32'hc20f53ec, 32'hc29ce9a1} /* (29, 1, 23) {real, imag} */,
  {32'hc203ebc4, 32'hc28df5b4} /* (29, 1, 22) {real, imag} */,
  {32'hc12fedc0, 32'hc243d83f} /* (29, 1, 21) {real, imag} */,
  {32'hc1e888ac, 32'h41e7c688} /* (29, 1, 20) {real, imag} */,
  {32'hc1dbb601, 32'h41bc5d6c} /* (29, 1, 19) {real, imag} */,
  {32'hc10e1dd8, 32'h42015a68} /* (29, 1, 18) {real, imag} */,
  {32'h3ef645c0, 32'h41ee1381} /* (29, 1, 17) {real, imag} */,
  {32'hc167631f, 32'h42616478} /* (29, 1, 16) {real, imag} */,
  {32'hc11380aa, 32'h428655b0} /* (29, 1, 15) {real, imag} */,
  {32'h40af4d18, 32'h429938f1} /* (29, 1, 14) {real, imag} */,
  {32'h41e6038b, 32'h42bfaaf7} /* (29, 1, 13) {real, imag} */,
  {32'h4210f1a7, 32'h42eea4d1} /* (29, 1, 12) {real, imag} */,
  {32'h42085c0b, 32'h42b923f0} /* (29, 1, 11) {real, imag} */,
  {32'h4265e188, 32'hc1ded9f5} /* (29, 1, 10) {real, imag} */,
  {32'h424a2b61, 32'hc2894ff9} /* (29, 1, 9) {real, imag} */,
  {32'h41bfd9fa, 32'hc29e65b5} /* (29, 1, 8) {real, imag} */,
  {32'h41db475c, 32'hc29017a0} /* (29, 1, 7) {real, imag} */,
  {32'h41bf19b6, 32'hc2147f58} /* (29, 1, 6) {real, imag} */,
  {32'hc05b9140, 32'hc2794f7c} /* (29, 1, 5) {real, imag} */,
  {32'hc06b3664, 32'hc29efe36} /* (29, 1, 4) {real, imag} */,
  {32'hc154132a, 32'hc29c94ce} /* (29, 1, 3) {real, imag} */,
  {32'hc1dca6de, 32'hc2877dd2} /* (29, 1, 2) {real, imag} */,
  {32'hc1e332c4, 32'hc29b3c63} /* (29, 1, 1) {real, imag} */,
  {32'hc0e11131, 32'hc2261035} /* (29, 1, 0) {real, imag} */,
  {32'hc1d7bcb8, 32'hc140dd72} /* (29, 0, 31) {real, imag} */,
  {32'hc1da627f, 32'hc1fd60d0} /* (29, 0, 30) {real, imag} */,
  {32'h415470fa, 32'hc283f754} /* (29, 0, 29) {real, imag} */,
  {32'hc189cf68, 32'hc25ca8f6} /* (29, 0, 28) {real, imag} */,
  {32'hc1935af2, 32'hc2894d24} /* (29, 0, 27) {real, imag} */,
  {32'h4103887b, 32'hc29f7944} /* (29, 0, 26) {real, imag} */,
  {32'h420beac4, 32'hc2826d1e} /* (29, 0, 25) {real, imag} */,
  {32'hbfdd9c13, 32'hc2179f55} /* (29, 0, 24) {real, imag} */,
  {32'hc1ba9dc7, 32'hc20e52c3} /* (29, 0, 23) {real, imag} */,
  {32'hc21c6dc0, 32'hc21a4c1c} /* (29, 0, 22) {real, imag} */,
  {32'hc23eb860, 32'hc23bc64f} /* (29, 0, 21) {real, imag} */,
  {32'hc06216a6, 32'hc10707da} /* (29, 0, 20) {real, imag} */,
  {32'h4130e6fd, 32'h412da657} /* (29, 0, 19) {real, imag} */,
  {32'hc10f65e1, 32'h4087a9a0} /* (29, 0, 18) {real, imag} */,
  {32'hc1c738b2, 32'hc0dc9774} /* (29, 0, 17) {real, imag} */,
  {32'hc14b2c47, 32'h3f92b94a} /* (29, 0, 16) {real, imag} */,
  {32'h407da895, 32'h422f9456} /* (29, 0, 15) {real, imag} */,
  {32'h41f502d8, 32'h428b422b} /* (29, 0, 14) {real, imag} */,
  {32'h4193c400, 32'h4259683b} /* (29, 0, 13) {real, imag} */,
  {32'h40f7b353, 32'h4282b239} /* (29, 0, 12) {real, imag} */,
  {32'hc0f26932, 32'h427e2a21} /* (29, 0, 11) {real, imag} */,
  {32'hc1cfc3a8, 32'h413db1b8} /* (29, 0, 10) {real, imag} */,
  {32'hc10ca8ac, 32'h4015a57c} /* (29, 0, 9) {real, imag} */,
  {32'hc1513273, 32'h406452cb} /* (29, 0, 8) {real, imag} */,
  {32'h3f934169, 32'h40b37ce2} /* (29, 0, 7) {real, imag} */,
  {32'h413d23d8, 32'h41d65bbe} /* (29, 0, 6) {real, imag} */,
  {32'hc06ff0ce, 32'hc1865533} /* (29, 0, 5) {real, imag} */,
  {32'hbe1250a0, 32'hc2619f80} /* (29, 0, 4) {real, imag} */,
  {32'hc178637a, 32'hc2945984} /* (29, 0, 3) {real, imag} */,
  {32'hc0ff3f07, 32'hc2665c6e} /* (29, 0, 2) {real, imag} */,
  {32'hc1318306, 32'hc20d76db} /* (29, 0, 1) {real, imag} */,
  {32'hc189b514, 32'hc1ca3030} /* (29, 0, 0) {real, imag} */,
  {32'hc120003b, 32'hc203b8f7} /* (28, 31, 31) {real, imag} */,
  {32'hc23704da, 32'hc27e6b74} /* (28, 31, 30) {real, imag} */,
  {32'hc282e3ac, 32'hc284d6a9} /* (28, 31, 29) {real, imag} */,
  {32'hc237e123, 32'hc28d26d8} /* (28, 31, 28) {real, imag} */,
  {32'hc2131964, 32'hc2810d89} /* (28, 31, 27) {real, imag} */,
  {32'hc218de84, 32'hc26a8a88} /* (28, 31, 26) {real, imag} */,
  {32'hc20cfaab, 32'hc2817cd1} /* (28, 31, 25) {real, imag} */,
  {32'hc1dc55c8, 32'hc2885db2} /* (28, 31, 24) {real, imag} */,
  {32'hc25c742b, 32'hc2987b26} /* (28, 31, 23) {real, imag} */,
  {32'hc24a00ce, 32'hc2c1e51c} /* (28, 31, 22) {real, imag} */,
  {32'hc24d0b16, 32'hc2954ce0} /* (28, 31, 21) {real, imag} */,
  {32'h3fc4f588, 32'h41b54f73} /* (28, 31, 20) {real, imag} */,
  {32'h421b62bc, 32'h4209252e} /* (28, 31, 19) {real, imag} */,
  {32'h42222bad, 32'hc0b0fd3c} /* (28, 31, 18) {real, imag} */,
  {32'h421ad2be, 32'h415db410} /* (28, 31, 17) {real, imag} */,
  {32'h422910ff, 32'h41a472cb} /* (28, 31, 16) {real, imag} */,
  {32'h41a6226f, 32'h425d629f} /* (28, 31, 15) {real, imag} */,
  {32'h42461404, 32'h42aea7cc} /* (28, 31, 14) {real, imag} */,
  {32'h42363bcb, 32'h42a48ca8} /* (28, 31, 13) {real, imag} */,
  {32'h419e4b99, 32'h428dc1f1} /* (28, 31, 12) {real, imag} */,
  {32'h41af5bac, 32'h428d9ad9} /* (28, 31, 11) {real, imag} */,
  {32'hc1cc223a, 32'hbed88360} /* (28, 31, 10) {real, imag} */,
  {32'hc29dcfa4, 32'hc11d49d2} /* (28, 31, 9) {real, imag} */,
  {32'hc27487ff, 32'hc0f6d478} /* (28, 31, 8) {real, imag} */,
  {32'hc2851dd1, 32'hc1f7ffc2} /* (28, 31, 7) {real, imag} */,
  {32'hc2667d0c, 32'hc1ddd458} /* (28, 31, 6) {real, imag} */,
  {32'hc23efa63, 32'hc23d8831} /* (28, 31, 5) {real, imag} */,
  {32'hc20a69a4, 32'hc280de3c} /* (28, 31, 4) {real, imag} */,
  {32'hc2061257, 32'hc2715523} /* (28, 31, 3) {real, imag} */,
  {32'hc2153b50, 32'hc289903c} /* (28, 31, 2) {real, imag} */,
  {32'hc179a4e7, 32'hc297ac21} /* (28, 31, 1) {real, imag} */,
  {32'hc111d775, 32'hc21c27d4} /* (28, 31, 0) {real, imag} */,
  {32'h41b992dc, 32'h420393e2} /* (28, 30, 31) {real, imag} */,
  {32'h42107b62, 32'h425122fb} /* (28, 30, 30) {real, imag} */,
  {32'h4206b0cb, 32'h422f984c} /* (28, 30, 29) {real, imag} */,
  {32'h41acfbf3, 32'h41f7af7b} /* (28, 30, 28) {real, imag} */,
  {32'h41fd9432, 32'h423c467a} /* (28, 30, 27) {real, imag} */,
  {32'h4164c19e, 32'h427595d2} /* (28, 30, 26) {real, imag} */,
  {32'h41868a22, 32'h42392a20} /* (28, 30, 25) {real, imag} */,
  {32'h41eeb878, 32'h42265370} /* (28, 30, 24) {real, imag} */,
  {32'h4204d78c, 32'h423314be} /* (28, 30, 23) {real, imag} */,
  {32'h41f77eb5, 32'h426e8c8e} /* (28, 30, 22) {real, imag} */,
  {32'h41cfc7f9, 32'h4120bcaa} /* (28, 30, 21) {real, imag} */,
  {32'h41b71f80, 32'hc29c0db8} /* (28, 30, 20) {real, imag} */,
  {32'h4076e970, 32'hc294b741} /* (28, 30, 19) {real, imag} */,
  {32'h40bfa508, 32'hc2923f16} /* (28, 30, 18) {real, imag} */,
  {32'hc1324be6, 32'hc2a5c168} /* (28, 30, 17) {real, imag} */,
  {32'hc20c88aa, 32'hc28a7578} /* (28, 30, 16) {real, imag} */,
  {32'hc1b5ea7e, 32'hc23bd4d8} /* (28, 30, 15) {real, imag} */,
  {32'hc189dda8, 32'hc2660e3d} /* (28, 30, 14) {real, imag} */,
  {32'hc15dff4d, 32'hc2280ea4} /* (28, 30, 13) {real, imag} */,
  {32'hc1c67ca1, 32'hc207d746} /* (28, 30, 12) {real, imag} */,
  {32'hc1893427, 32'hbfbde688} /* (28, 30, 11) {real, imag} */,
  {32'hc131373a, 32'h428bf1f7} /* (28, 30, 10) {real, imag} */,
  {32'h40b65478, 32'h42c06e81} /* (28, 30, 9) {real, imag} */,
  {32'h408c5da4, 32'h42a44507} /* (28, 30, 8) {real, imag} */,
  {32'h3e9b4e00, 32'h428a2dd6} /* (28, 30, 7) {real, imag} */,
  {32'h40322934, 32'h427910b9} /* (28, 30, 6) {real, imag} */,
  {32'h4190a22e, 32'h425250ef} /* (28, 30, 5) {real, imag} */,
  {32'h41e964e8, 32'h41ecdda8} /* (28, 30, 4) {real, imag} */,
  {32'h41c2fcac, 32'h4225729c} /* (28, 30, 3) {real, imag} */,
  {32'h418d4428, 32'h425f6685} /* (28, 30, 2) {real, imag} */,
  {32'h41cadad7, 32'h426a6761} /* (28, 30, 1) {real, imag} */,
  {32'h410e3698, 32'h42034062} /* (28, 30, 0) {real, imag} */,
  {32'h4141a3a4, 32'hc08d6788} /* (28, 29, 31) {real, imag} */,
  {32'h4126198e, 32'hbe4cae90} /* (28, 29, 30) {real, imag} */,
  {32'hc12091a6, 32'h41147fd3} /* (28, 29, 29) {real, imag} */,
  {32'hc1b59618, 32'h40ceb472} /* (28, 29, 28) {real, imag} */,
  {32'hc04b663c, 32'hc18793d4} /* (28, 29, 27) {real, imag} */,
  {32'h41251231, 32'hc147264a} /* (28, 29, 26) {real, imag} */,
  {32'h411e19ad, 32'h402796e6} /* (28, 29, 25) {real, imag} */,
  {32'hc1896ce4, 32'h41710de0} /* (28, 29, 24) {real, imag} */,
  {32'h3f5f1ec0, 32'h412ed725} /* (28, 29, 23) {real, imag} */,
  {32'h40465672, 32'hc1986db0} /* (28, 29, 22) {real, imag} */,
  {32'h414bb40d, 32'hc0259ac4} /* (28, 29, 21) {real, imag} */,
  {32'h4200b621, 32'hc192d86a} /* (28, 29, 20) {real, imag} */,
  {32'h41621f8a, 32'hc1e3d77c} /* (28, 29, 19) {real, imag} */,
  {32'h40f38e60, 32'hc1d89d1c} /* (28, 29, 18) {real, imag} */,
  {32'h4208c027, 32'hc174c895} /* (28, 29, 17) {real, imag} */,
  {32'h41c89bd4, 32'hc12e843c} /* (28, 29, 16) {real, imag} */,
  {32'h41346621, 32'h41254bab} /* (28, 29, 15) {real, imag} */,
  {32'h41ca4636, 32'hc0a209c5} /* (28, 29, 14) {real, imag} */,
  {32'h3fcd7a38, 32'hbfa4fa88} /* (28, 29, 13) {real, imag} */,
  {32'hbff4cb10, 32'hc1a94694} /* (28, 29, 12) {real, imag} */,
  {32'hc18b8366, 32'hc0c8aabc} /* (28, 29, 11) {real, imag} */,
  {32'hc212bc8c, 32'h4182fb98} /* (28, 29, 10) {real, imag} */,
  {32'hc1d5b09c, 32'h40880d5c} /* (28, 29, 9) {real, imag} */,
  {32'hc137332b, 32'h40cb8fbe} /* (28, 29, 8) {real, imag} */,
  {32'hc1b7f230, 32'h4179fce0} /* (28, 29, 7) {real, imag} */,
  {32'hc1916d00, 32'h41e9740f} /* (28, 29, 6) {real, imag} */,
  {32'hc085a8f4, 32'h4187cd89} /* (28, 29, 5) {real, imag} */,
  {32'h41211723, 32'h414932c9} /* (28, 29, 4) {real, imag} */,
  {32'h3fc27780, 32'h42035cf5} /* (28, 29, 3) {real, imag} */,
  {32'hc04faa20, 32'h4199e17d} /* (28, 29, 2) {real, imag} */,
  {32'h4093bfb6, 32'h40dc714c} /* (28, 29, 1) {real, imag} */,
  {32'hbf94c9f8, 32'hc0df29cc} /* (28, 29, 0) {real, imag} */,
  {32'hc1a859b0, 32'hc11a1be3} /* (28, 28, 31) {real, imag} */,
  {32'hc1656d0c, 32'hc1a9b4b4} /* (28, 28, 30) {real, imag} */,
  {32'hbeadc540, 32'hc17b5438} /* (28, 28, 29) {real, imag} */,
  {32'h4108ca38, 32'hc18cd841} /* (28, 28, 28) {real, imag} */,
  {32'hc08434ee, 32'hc14964c7} /* (28, 28, 27) {real, imag} */,
  {32'hc178035e, 32'hc1129d76} /* (28, 28, 26) {real, imag} */,
  {32'hc1b131bc, 32'hc17c02da} /* (28, 28, 25) {real, imag} */,
  {32'hc2088d42, 32'hc0e43580} /* (28, 28, 24) {real, imag} */,
  {32'hc1e9ecf7, 32'hbfae7420} /* (28, 28, 23) {real, imag} */,
  {32'hc134c712, 32'h40a06aa6} /* (28, 28, 22) {real, imag} */,
  {32'h419d61f6, 32'h417e3242} /* (28, 28, 21) {real, imag} */,
  {32'h42167f26, 32'h418b1594} /* (28, 28, 20) {real, imag} */,
  {32'h41dd7a48, 32'h41c4ab3e} /* (28, 28, 19) {real, imag} */,
  {32'h42373c59, 32'h41183573} /* (28, 28, 18) {real, imag} */,
  {32'h427020ea, 32'h40ce8232} /* (28, 28, 17) {real, imag} */,
  {32'h41dc7882, 32'h41883bbc} /* (28, 28, 16) {real, imag} */,
  {32'h4099e607, 32'h419a5d75} /* (28, 28, 15) {real, imag} */,
  {32'h406cda5b, 32'h41df8cbc} /* (28, 28, 14) {real, imag} */,
  {32'hc05c9a60, 32'h41af9235} /* (28, 28, 13) {real, imag} */,
  {32'h413dbe0c, 32'h41e74101} /* (28, 28, 12) {real, imag} */,
  {32'h417590fd, 32'h415d9635} /* (28, 28, 11) {real, imag} */,
  {32'hc150e68c, 32'hc11c49ed} /* (28, 28, 10) {real, imag} */,
  {32'hc24d6afc, 32'hc0978522} /* (28, 28, 9) {real, imag} */,
  {32'hc22d990e, 32'hc101204b} /* (28, 28, 8) {real, imag} */,
  {32'hc1c6291a, 32'hc0463454} /* (28, 28, 7) {real, imag} */,
  {32'hc19e1408, 32'h404380d8} /* (28, 28, 6) {real, imag} */,
  {32'hc1b6d097, 32'hc170b49b} /* (28, 28, 5) {real, imag} */,
  {32'hc1827992, 32'hc1500a07} /* (28, 28, 4) {real, imag} */,
  {32'h3fd3f624, 32'hc1eb5896} /* (28, 28, 3) {real, imag} */,
  {32'hc18079c9, 32'hc1e08424} /* (28, 28, 2) {real, imag} */,
  {32'hc1b3edce, 32'hc20cc0f6} /* (28, 28, 1) {real, imag} */,
  {32'hc156162b, 32'hc1bdd97d} /* (28, 28, 0) {real, imag} */,
  {32'h4168f843, 32'hbfd065c8} /* (28, 27, 31) {real, imag} */,
  {32'h41eef078, 32'hbf5addb0} /* (28, 27, 30) {real, imag} */,
  {32'h415c993e, 32'h4114d9b0} /* (28, 27, 29) {real, imag} */,
  {32'h4022ea11, 32'h416b82b8} /* (28, 27, 28) {real, imag} */,
  {32'h41795831, 32'h4146f4dc} /* (28, 27, 27) {real, imag} */,
  {32'h418ce592, 32'h417d3acc} /* (28, 27, 26) {real, imag} */,
  {32'h416db7e7, 32'h41c48166} /* (28, 27, 25) {real, imag} */,
  {32'h410b4015, 32'h41b7b686} /* (28, 27, 24) {real, imag} */,
  {32'h3f09eebc, 32'h41cd1282} /* (28, 27, 23) {real, imag} */,
  {32'h40ad4f6b, 32'h418a312b} /* (28, 27, 22) {real, imag} */,
  {32'h40eb16f0, 32'hc125215e} /* (28, 27, 21) {real, imag} */,
  {32'h40a91ca2, 32'hc1478f9e} /* (28, 27, 20) {real, imag} */,
  {32'hc14be6d6, 32'h411f36de} /* (28, 27, 19) {real, imag} */,
  {32'hc193dc79, 32'h40be8e1f} /* (28, 27, 18) {real, imag} */,
  {32'hc121510e, 32'hc0e9242b} /* (28, 27, 17) {real, imag} */,
  {32'hc048add9, 32'hc0c9d86c} /* (28, 27, 16) {real, imag} */,
  {32'hbece8ce0, 32'hc18aacd8} /* (28, 27, 15) {real, imag} */,
  {32'hbf1dc3f8, 32'hc1bc55f0} /* (28, 27, 14) {real, imag} */,
  {32'hc0279683, 32'hc07fe220} /* (28, 27, 13) {real, imag} */,
  {32'hc13b44dc, 32'hc0975b60} /* (28, 27, 12) {real, imag} */,
  {32'hc1a5c3b1, 32'hc1437cdb} /* (28, 27, 11) {real, imag} */,
  {32'h4113694c, 32'hc00400ee} /* (28, 27, 10) {real, imag} */,
  {32'h410c377d, 32'h405da805} /* (28, 27, 9) {real, imag} */,
  {32'h4185b683, 32'h417a87fb} /* (28, 27, 8) {real, imag} */,
  {32'h4196da05, 32'hc0d6f989} /* (28, 27, 7) {real, imag} */,
  {32'hc0c609c2, 32'hc19edf04} /* (28, 27, 6) {real, imag} */,
  {32'h411bee61, 32'hc02a3578} /* (28, 27, 5) {real, imag} */,
  {32'h415f60b0, 32'h41d96fb9} /* (28, 27, 4) {real, imag} */,
  {32'h4135999a, 32'h42029c3f} /* (28, 27, 3) {real, imag} */,
  {32'h4116f89c, 32'h4138dfa7} /* (28, 27, 2) {real, imag} */,
  {32'hbefb5a70, 32'h41021623} /* (28, 27, 1) {real, imag} */,
  {32'h4118f3da, 32'h4136652b} /* (28, 27, 0) {real, imag} */,
  {32'hc1772363, 32'h40b40aca} /* (28, 26, 31) {real, imag} */,
  {32'hc1ffee04, 32'h41a2f687} /* (28, 26, 30) {real, imag} */,
  {32'hc0d9bbf8, 32'h4193ad97} /* (28, 26, 29) {real, imag} */,
  {32'h410ae618, 32'h404e4980} /* (28, 26, 28) {real, imag} */,
  {32'hc17f6f6f, 32'h40735e8f} /* (28, 26, 27) {real, imag} */,
  {32'hc18b79ab, 32'h408c5928} /* (28, 26, 26) {real, imag} */,
  {32'hbe469f40, 32'h40d2bbfc} /* (28, 26, 25) {real, imag} */,
  {32'h412f47d5, 32'h40de4f24} /* (28, 26, 24) {real, imag} */,
  {32'h40b1610f, 32'hc0283d38} /* (28, 26, 23) {real, imag} */,
  {32'hbf587740, 32'h41138a6d} /* (28, 26, 22) {real, imag} */,
  {32'h4091d641, 32'h411c14c4} /* (28, 26, 21) {real, imag} */,
  {32'h4012f9b9, 32'h3e37c5c0} /* (28, 26, 20) {real, imag} */,
  {32'h41161529, 32'hc02d5a00} /* (28, 26, 19) {real, imag} */,
  {32'h419258a9, 32'h4036a79a} /* (28, 26, 18) {real, imag} */,
  {32'hc084b977, 32'h3fcf8d92} /* (28, 26, 17) {real, imag} */,
  {32'hc119bfd7, 32'h3f9d41cc} /* (28, 26, 16) {real, imag} */,
  {32'hbea41ea0, 32'h407ad554} /* (28, 26, 15) {real, imag} */,
  {32'hc1b8b57c, 32'hbfc0fe88} /* (28, 26, 14) {real, imag} */,
  {32'hc18d9952, 32'h404e4dd8} /* (28, 26, 13) {real, imag} */,
  {32'h406cfc5c, 32'h410e0019} /* (28, 26, 12) {real, imag} */,
  {32'h41023948, 32'h3fd54cd0} /* (28, 26, 11) {real, imag} */,
  {32'h4083fef6, 32'h40cb67e7} /* (28, 26, 10) {real, imag} */,
  {32'hbf8420be, 32'hc00e1814} /* (28, 26, 9) {real, imag} */,
  {32'h4161dec2, 32'hc117ea48} /* (28, 26, 8) {real, imag} */,
  {32'h4180d5a9, 32'hc066c2f8} /* (28, 26, 7) {real, imag} */,
  {32'h40b7bd60, 32'h40ec20bc} /* (28, 26, 6) {real, imag} */,
  {32'h407133e8, 32'h411c18e7} /* (28, 26, 5) {real, imag} */,
  {32'h3f784ac8, 32'h40207036} /* (28, 26, 4) {real, imag} */,
  {32'hc06c7c24, 32'h410286a9} /* (28, 26, 3) {real, imag} */,
  {32'h3fd10b68, 32'hc160af7d} /* (28, 26, 2) {real, imag} */,
  {32'hc171a45a, 32'hbe86f200} /* (28, 26, 1) {real, imag} */,
  {32'hc1282a0c, 32'h4142f25f} /* (28, 26, 0) {real, imag} */,
  {32'hc07f4864, 32'hc0d62e5c} /* (28, 25, 31) {real, imag} */,
  {32'h3ffd8628, 32'hc0cc18ab} /* (28, 25, 30) {real, imag} */,
  {32'hc0a8cdbe, 32'hc1599c9f} /* (28, 25, 29) {real, imag} */,
  {32'hc17ae413, 32'hc15580ac} /* (28, 25, 28) {real, imag} */,
  {32'hc1765a4c, 32'h400ec34a} /* (28, 25, 27) {real, imag} */,
  {32'hc151465e, 32'hc008225c} /* (28, 25, 26) {real, imag} */,
  {32'h406b6dca, 32'hc1b38270} /* (28, 25, 25) {real, imag} */,
  {32'h413ca87d, 32'hc19922a9} /* (28, 25, 24) {real, imag} */,
  {32'hc171704e, 32'hc14f2452} /* (28, 25, 23) {real, imag} */,
  {32'hc1a61268, 32'hc070fc3e} /* (28, 25, 22) {real, imag} */,
  {32'hc20127ef, 32'hc1bf650c} /* (28, 25, 21) {real, imag} */,
  {32'hc1cb42b1, 32'hc122491f} /* (28, 25, 20) {real, imag} */,
  {32'h40ba2b2b, 32'hc0ff9701} /* (28, 25, 19) {real, imag} */,
  {32'h41d75aaa, 32'h4082ab0e} /* (28, 25, 18) {real, imag} */,
  {32'h414776e0, 32'h416c1ae3} /* (28, 25, 17) {real, imag} */,
  {32'h402c1d52, 32'hc0fbb772} /* (28, 25, 16) {real, imag} */,
  {32'h416b6bea, 32'hbfb93f50} /* (28, 25, 15) {real, imag} */,
  {32'h419c3e46, 32'h4126c6cb} /* (28, 25, 14) {real, imag} */,
  {32'h3e30be80, 32'h415d6672} /* (28, 25, 13) {real, imag} */,
  {32'h413dc062, 32'h41366898} /* (28, 25, 12) {real, imag} */,
  {32'h4154fec6, 32'h40ccbf92} /* (28, 25, 11) {real, imag} */,
  {32'hbf6cc7e0, 32'hc0ae506c} /* (28, 25, 10) {real, imag} */,
  {32'hbeaa16e0, 32'h41051db2} /* (28, 25, 9) {real, imag} */,
  {32'hc0ca87e2, 32'h4140ed68} /* (28, 25, 8) {real, imag} */,
  {32'hc18ccf87, 32'hc00d1688} /* (28, 25, 7) {real, imag} */,
  {32'hc18060e0, 32'hc111f790} /* (28, 25, 6) {real, imag} */,
  {32'hc0a961ec, 32'hc0299b48} /* (28, 25, 5) {real, imag} */,
  {32'h4165b1c7, 32'h4084c590} /* (28, 25, 4) {real, imag} */,
  {32'h40fde46a, 32'hc051348b} /* (28, 25, 3) {real, imag} */,
  {32'hc0a41f62, 32'hbed2ced0} /* (28, 25, 2) {real, imag} */,
  {32'hc1959f9c, 32'hc085581c} /* (28, 25, 1) {real, imag} */,
  {32'hc0e15131, 32'hbeddb5f8} /* (28, 25, 0) {real, imag} */,
  {32'h40d5b83b, 32'hc114914a} /* (28, 24, 31) {real, imag} */,
  {32'h3ff82ad0, 32'h3fceee04} /* (28, 24, 30) {real, imag} */,
  {32'hbf9b09b0, 32'h412ae894} /* (28, 24, 29) {real, imag} */,
  {32'h41cbff14, 32'h41860410} /* (28, 24, 28) {real, imag} */,
  {32'h41c21a2f, 32'h41bb0eb4} /* (28, 24, 27) {real, imag} */,
  {32'h4180c5e6, 32'h418f926b} /* (28, 24, 26) {real, imag} */,
  {32'h4194bc02, 32'h41640030} /* (28, 24, 25) {real, imag} */,
  {32'h412797a2, 32'h40868f16} /* (28, 24, 24) {real, imag} */,
  {32'h41497a26, 32'h4053323c} /* (28, 24, 23) {real, imag} */,
  {32'h41854dee, 32'h40bbd9b5} /* (28, 24, 22) {real, imag} */,
  {32'hc088b4ba, 32'hc074cd10} /* (28, 24, 21) {real, imag} */,
  {32'hc201c9d2, 32'hc083cec6} /* (28, 24, 20) {real, imag} */,
  {32'hc1b8ebfb, 32'hc0eea661} /* (28, 24, 19) {real, imag} */,
  {32'hc1a14628, 32'hc135025e} /* (28, 24, 18) {real, imag} */,
  {32'hc1a9b266, 32'hc1278384} /* (28, 24, 17) {real, imag} */,
  {32'hc18afdae, 32'hc0b03d2c} /* (28, 24, 16) {real, imag} */,
  {32'hc107cba4, 32'hc1b39b0a} /* (28, 24, 15) {real, imag} */,
  {32'h408c7c28, 32'hc14294fa} /* (28, 24, 14) {real, imag} */,
  {32'hc08b40f4, 32'hc0d144e8} /* (28, 24, 13) {real, imag} */,
  {32'hc1ad904e, 32'hc1966232} /* (28, 24, 12) {real, imag} */,
  {32'hc1f142c8, 32'hc177b9b3} /* (28, 24, 11) {real, imag} */,
  {32'hc1dde6b9, 32'hc122ffa2} /* (28, 24, 10) {real, imag} */,
  {32'h410d8100, 32'h3e65a4a0} /* (28, 24, 9) {real, imag} */,
  {32'h41c37670, 32'h41a39693} /* (28, 24, 8) {real, imag} */,
  {32'h41aa609a, 32'h41957bb0} /* (28, 24, 7) {real, imag} */,
  {32'h4088901b, 32'h418cb965} /* (28, 24, 6) {real, imag} */,
  {32'hc0841ecf, 32'h40bd4bd6} /* (28, 24, 5) {real, imag} */,
  {32'h41648c7e, 32'h40bfac7d} /* (28, 24, 4) {real, imag} */,
  {32'h41223c94, 32'hc0bd2a1c} /* (28, 24, 3) {real, imag} */,
  {32'h41122751, 32'h40c8fd21} /* (28, 24, 2) {real, imag} */,
  {32'h41c64cb2, 32'h4099794c} /* (28, 24, 1) {real, imag} */,
  {32'h4193aaee, 32'hc0a1e334} /* (28, 24, 0) {real, imag} */,
  {32'hc03d4ba1, 32'hbfbe64e2} /* (28, 23, 31) {real, imag} */,
  {32'hc1116785, 32'h40b39a6f} /* (28, 23, 30) {real, imag} */,
  {32'hc08040ce, 32'hbd011540} /* (28, 23, 29) {real, imag} */,
  {32'h3f36d218, 32'hc0512d8c} /* (28, 23, 28) {real, imag} */,
  {32'h40f43b7f, 32'hc072add8} /* (28, 23, 27) {real, imag} */,
  {32'h405a09f0, 32'h40314694} /* (28, 23, 26) {real, imag} */,
  {32'hc1a1024b, 32'h4052d748} /* (28, 23, 25) {real, imag} */,
  {32'hc1980868, 32'hc118b960} /* (28, 23, 24) {real, imag} */,
  {32'hc0ad8cd5, 32'hc1674c7e} /* (28, 23, 23) {real, imag} */,
  {32'h3fc1db0c, 32'h3e6fd8e0} /* (28, 23, 22) {real, imag} */,
  {32'h4093a3ed, 32'h41574ba8} /* (28, 23, 21) {real, imag} */,
  {32'h4094dd88, 32'h3e2de280} /* (28, 23, 20) {real, imag} */,
  {32'h412410c3, 32'hc136b7cc} /* (28, 23, 19) {real, imag} */,
  {32'h41869aa8, 32'hc18965fe} /* (28, 23, 18) {real, imag} */,
  {32'h4189d18e, 32'hc190d198} /* (28, 23, 17) {real, imag} */,
  {32'h40050fae, 32'hc0880b5e} /* (28, 23, 16) {real, imag} */,
  {32'hc05f13fc, 32'h4128c906} /* (28, 23, 15) {real, imag} */,
  {32'hc096b50c, 32'h412503bd} /* (28, 23, 14) {real, imag} */,
  {32'hbf4789ec, 32'h40cc4fb7} /* (28, 23, 13) {real, imag} */,
  {32'h40bf3bd6, 32'h411890e5} /* (28, 23, 12) {real, imag} */,
  {32'h3f22b284, 32'h3f159a2c} /* (28, 23, 11) {real, imag} */,
  {32'hc0c8c537, 32'h409f65b9} /* (28, 23, 10) {real, imag} */,
  {32'hc18c03c6, 32'h410f8d8f} /* (28, 23, 9) {real, imag} */,
  {32'hc15c4e27, 32'hc07e5828} /* (28, 23, 8) {real, imag} */,
  {32'hc09a0a0f, 32'hbf832668} /* (28, 23, 7) {real, imag} */,
  {32'h40b2ea8e, 32'h414e19e0} /* (28, 23, 6) {real, imag} */,
  {32'h3ffcc738, 32'h41c64637} /* (28, 23, 5) {real, imag} */,
  {32'h40851082, 32'h4194317e} /* (28, 23, 4) {real, imag} */,
  {32'h3fe9da4a, 32'hbf49b834} /* (28, 23, 3) {real, imag} */,
  {32'hc0e5dee6, 32'h410701af} /* (28, 23, 2) {real, imag} */,
  {32'hc18696e7, 32'h40df3cd4} /* (28, 23, 1) {real, imag} */,
  {32'hbfc949ae, 32'hc0235aab} /* (28, 23, 0) {real, imag} */,
  {32'h3d8c4160, 32'h406d8754} /* (28, 22, 31) {real, imag} */,
  {32'hc0c01a92, 32'h41077c1a} /* (28, 22, 30) {real, imag} */,
  {32'h3eb13fc8, 32'h40b5f646} /* (28, 22, 29) {real, imag} */,
  {32'hc08b5ee4, 32'h4102c75e} /* (28, 22, 28) {real, imag} */,
  {32'hc1af5d88, 32'hc0e20614} /* (28, 22, 27) {real, imag} */,
  {32'hc18be1fb, 32'hc09afd92} /* (28, 22, 26) {real, imag} */,
  {32'h40160d9b, 32'h4122ccf2} /* (28, 22, 25) {real, imag} */,
  {32'h40a4754b, 32'h41942e2f} /* (28, 22, 24) {real, imag} */,
  {32'hc0f1232e, 32'h40b09726} /* (28, 22, 23) {real, imag} */,
  {32'hc110d37c, 32'h3faf087e} /* (28, 22, 22) {real, imag} */,
  {32'h40ad6a1c, 32'h3f34fac4} /* (28, 22, 21) {real, imag} */,
  {32'h410ed5db, 32'hbfc9917c} /* (28, 22, 20) {real, imag} */,
  {32'h40675f7c, 32'hc1072f85} /* (28, 22, 19) {real, imag} */,
  {32'h4094832e, 32'hc02a96be} /* (28, 22, 18) {real, imag} */,
  {32'h40ff73af, 32'hc0ca0a9c} /* (28, 22, 17) {real, imag} */,
  {32'hc0491b8c, 32'hc10afa9c} /* (28, 22, 16) {real, imag} */,
  {32'hc0b2c210, 32'hc058741c} /* (28, 22, 15) {real, imag} */,
  {32'h3efd5380, 32'h3ef83bb0} /* (28, 22, 14) {real, imag} */,
  {32'hc0a5f040, 32'hc0b541cc} /* (28, 22, 13) {real, imag} */,
  {32'hbfdbb6b0, 32'hbf91d8d4} /* (28, 22, 12) {real, imag} */,
  {32'hc051d859, 32'h40929818} /* (28, 22, 11) {real, imag} */,
  {32'hc0d717f6, 32'h4016c1d3} /* (28, 22, 10) {real, imag} */,
  {32'hc13016d1, 32'h408440b0} /* (28, 22, 9) {real, imag} */,
  {32'hc0e76704, 32'h3ff0436c} /* (28, 22, 8) {real, imag} */,
  {32'hc0f1a9c6, 32'h41180973} /* (28, 22, 7) {real, imag} */,
  {32'hc1743182, 32'hc0805fae} /* (28, 22, 6) {real, imag} */,
  {32'hc15a316d, 32'hc17a7a1a} /* (28, 22, 5) {real, imag} */,
  {32'hc0e87cfa, 32'h4041b518} /* (28, 22, 4) {real, imag} */,
  {32'h40d300d6, 32'h40a9cd3e} /* (28, 22, 3) {real, imag} */,
  {32'h40bbccc8, 32'hc14fb552} /* (28, 22, 2) {real, imag} */,
  {32'h410b0ad8, 32'hc0ddc6c1} /* (28, 22, 1) {real, imag} */,
  {32'h408031c4, 32'h3f17dd70} /* (28, 22, 0) {real, imag} */,
  {32'h41038919, 32'h40bb838a} /* (28, 21, 31) {real, imag} */,
  {32'h40b22d3f, 32'h40b13a26} /* (28, 21, 30) {real, imag} */,
  {32'h404eafc6, 32'h40f6e37b} /* (28, 21, 29) {real, imag} */,
  {32'h40b6a52b, 32'h415c12a4} /* (28, 21, 28) {real, imag} */,
  {32'hbf8168f4, 32'h41715efe} /* (28, 21, 27) {real, imag} */,
  {32'h4021b064, 32'h412bc38a} /* (28, 21, 26) {real, imag} */,
  {32'h4055905f, 32'hc0d9c901} /* (28, 21, 25) {real, imag} */,
  {32'h402c782b, 32'hc157a4eb} /* (28, 21, 24) {real, imag} */,
  {32'h410b258b, 32'hc096585e} /* (28, 21, 23) {real, imag} */,
  {32'h4139011a, 32'hc0dc8f36} /* (28, 21, 22) {real, imag} */,
  {32'h40b1e5be, 32'hc011cb88} /* (28, 21, 21) {real, imag} */,
  {32'hc0dacbfc, 32'h40732a1e} /* (28, 21, 20) {real, imag} */,
  {32'hc0c044c8, 32'h3eb9ca00} /* (28, 21, 19) {real, imag} */,
  {32'hc14034b4, 32'h40b3d16f} /* (28, 21, 18) {real, imag} */,
  {32'hc0c1a044, 32'h4122629d} /* (28, 21, 17) {real, imag} */,
  {32'hbf90dbd8, 32'h3f3a3678} /* (28, 21, 16) {real, imag} */,
  {32'hc12dc5c1, 32'h3f10e072} /* (28, 21, 15) {real, imag} */,
  {32'hc11d3109, 32'h40f6db46} /* (28, 21, 14) {real, imag} */,
  {32'hc13c565e, 32'hbf93dcc4} /* (28, 21, 13) {real, imag} */,
  {32'hbfd187b4, 32'hc00aafa6} /* (28, 21, 12) {real, imag} */,
  {32'hc0bde630, 32'hc0e55507} /* (28, 21, 11) {real, imag} */,
  {32'hbf150b88, 32'h3f58b520} /* (28, 21, 10) {real, imag} */,
  {32'h410df029, 32'hc082cb19} /* (28, 21, 9) {real, imag} */,
  {32'h401c3e0c, 32'hc0438c1e} /* (28, 21, 8) {real, imag} */,
  {32'hbf9b4980, 32'hc03f1f9e} /* (28, 21, 7) {real, imag} */,
  {32'h4126caf7, 32'hc071acc6} /* (28, 21, 6) {real, imag} */,
  {32'h403c1c0d, 32'hc0363b44} /* (28, 21, 5) {real, imag} */,
  {32'h40d3a8a1, 32'hc1406e10} /* (28, 21, 4) {real, imag} */,
  {32'h4117e65e, 32'hc1541050} /* (28, 21, 3) {real, imag} */,
  {32'h41347a18, 32'h4085c0a0} /* (28, 21, 2) {real, imag} */,
  {32'h41200422, 32'h4121e7ac} /* (28, 21, 1) {real, imag} */,
  {32'h3fce45f4, 32'h409ea046} /* (28, 21, 0) {real, imag} */,
  {32'hbe8ade70, 32'hc05db83f} /* (28, 20, 31) {real, imag} */,
  {32'h40c33e32, 32'h407ebf3c} /* (28, 20, 30) {real, imag} */,
  {32'hc102239e, 32'h40a8c9dd} /* (28, 20, 29) {real, imag} */,
  {32'hc194906c, 32'h408050e2} /* (28, 20, 28) {real, imag} */,
  {32'hc0814262, 32'h4083914e} /* (28, 20, 27) {real, imag} */,
  {32'h408def3f, 32'h407b6426} /* (28, 20, 26) {real, imag} */,
  {32'h3f938026, 32'h3f1bd5a8} /* (28, 20, 25) {real, imag} */,
  {32'h3e390d40, 32'h40083db7} /* (28, 20, 24) {real, imag} */,
  {32'h4059fa22, 32'h3da2a280} /* (28, 20, 23) {real, imag} */,
  {32'hbee6cba8, 32'hc0a643d4} /* (28, 20, 22) {real, imag} */,
  {32'h40aa88d2, 32'h40964b64} /* (28, 20, 21) {real, imag} */,
  {32'h3ffe88a4, 32'h3fe503c6} /* (28, 20, 20) {real, imag} */,
  {32'hbfd56b52, 32'hc009ed9d} /* (28, 20, 19) {real, imag} */,
  {32'h3fedae90, 32'hc082a2e4} /* (28, 20, 18) {real, imag} */,
  {32'h4030bd26, 32'hc0b364b0} /* (28, 20, 17) {real, imag} */,
  {32'h412664f4, 32'h3f8a3f5c} /* (28, 20, 16) {real, imag} */,
  {32'h40175a84, 32'hbf964a5b} /* (28, 20, 15) {real, imag} */,
  {32'hc058c9f4, 32'hc0054cd0} /* (28, 20, 14) {real, imag} */,
  {32'hbeb41580, 32'h403106cc} /* (28, 20, 13) {real, imag} */,
  {32'hc0d45be0, 32'h40ad7267} /* (28, 20, 12) {real, imag} */,
  {32'hc0892148, 32'h3fde4ec3} /* (28, 20, 11) {real, imag} */,
  {32'hc01b1e56, 32'hc0ff91ff} /* (28, 20, 10) {real, imag} */,
  {32'hbffe69ac, 32'hc1375371} /* (28, 20, 9) {real, imag} */,
  {32'hc12805bb, 32'h3f9a3aa8} /* (28, 20, 8) {real, imag} */,
  {32'hc0ea8c1e, 32'h400e0044} /* (28, 20, 7) {real, imag} */,
  {32'hbf011d60, 32'h3e860c70} /* (28, 20, 6) {real, imag} */,
  {32'h4049a164, 32'h402411ff} /* (28, 20, 5) {real, imag} */,
  {32'h4076e4c0, 32'hc08a629b} /* (28, 20, 4) {real, imag} */,
  {32'hc0ee972d, 32'hbee2a260} /* (28, 20, 3) {real, imag} */,
  {32'hbfe4e338, 32'h40cdd116} /* (28, 20, 2) {real, imag} */,
  {32'h3fdfcf3e, 32'h4144c919} /* (28, 20, 1) {real, imag} */,
  {32'hc02b22ac, 32'h401fa8ca} /* (28, 20, 0) {real, imag} */,
  {32'hc0728c06, 32'hc0d5e8e0} /* (28, 19, 31) {real, imag} */,
  {32'hc09fb446, 32'hc0082317} /* (28, 19, 30) {real, imag} */,
  {32'hbe9582d8, 32'hbfbe92ae} /* (28, 19, 29) {real, imag} */,
  {32'hbe8dbeb0, 32'h40ec5e46} /* (28, 19, 28) {real, imag} */,
  {32'h3f4566c2, 32'h408b50b3} /* (28, 19, 27) {real, imag} */,
  {32'h4090ffc3, 32'h3fcf1c4c} /* (28, 19, 26) {real, imag} */,
  {32'h40ad37c6, 32'h409217ee} /* (28, 19, 25) {real, imag} */,
  {32'hc0948274, 32'hc015cd78} /* (28, 19, 24) {real, imag} */,
  {32'hc1266ac2, 32'hc0844b96} /* (28, 19, 23) {real, imag} */,
  {32'hc0831be4, 32'hc003a16b} /* (28, 19, 22) {real, imag} */,
  {32'hbf1fd280, 32'hbe4fb900} /* (28, 19, 21) {real, imag} */,
  {32'hbd6b6340, 32'h40eac59a} /* (28, 19, 20) {real, imag} */,
  {32'hc0c00656, 32'h40dd242f} /* (28, 19, 19) {real, imag} */,
  {32'hc0d88fca, 32'h40b2508c} /* (28, 19, 18) {real, imag} */,
  {32'h40327a48, 32'h4032edcd} /* (28, 19, 17) {real, imag} */,
  {32'hbedd7400, 32'h40a5fe17} /* (28, 19, 16) {real, imag} */,
  {32'hbf67a938, 32'h40d98e4a} /* (28, 19, 15) {real, imag} */,
  {32'h40570fec, 32'h3fa8892d} /* (28, 19, 14) {real, imag} */,
  {32'h4071f512, 32'h411cd7a0} /* (28, 19, 13) {real, imag} */,
  {32'hc0938eb4, 32'h41373e95} /* (28, 19, 12) {real, imag} */,
  {32'hbee344e8, 32'h40849f42} /* (28, 19, 11) {real, imag} */,
  {32'h3f00ce38, 32'hc095ee0e} /* (28, 19, 10) {real, imag} */,
  {32'hc060b6ca, 32'hc02adf42} /* (28, 19, 9) {real, imag} */,
  {32'hc0a6905e, 32'h407383a0} /* (28, 19, 8) {real, imag} */,
  {32'hc0d21900, 32'h402fb8e5} /* (28, 19, 7) {real, imag} */,
  {32'hbfcdcdac, 32'hbfbe8758} /* (28, 19, 6) {real, imag} */,
  {32'hc0bcfdaf, 32'hc0c45bae} /* (28, 19, 5) {real, imag} */,
  {32'hc0f18f77, 32'hc02a001b} /* (28, 19, 4) {real, imag} */,
  {32'hc0dfbd3e, 32'h40826640} /* (28, 19, 3) {real, imag} */,
  {32'hc0d3a6ae, 32'hbf9764f8} /* (28, 19, 2) {real, imag} */,
  {32'hbf3cb054, 32'hc06f3ca1} /* (28, 19, 1) {real, imag} */,
  {32'h3dd32ac0, 32'hc0dd33d4} /* (28, 19, 0) {real, imag} */,
  {32'h409d64b5, 32'hc01debe9} /* (28, 18, 31) {real, imag} */,
  {32'hbecb05a0, 32'hc039fd83} /* (28, 18, 30) {real, imag} */,
  {32'h40146278, 32'h40216a47} /* (28, 18, 29) {real, imag} */,
  {32'h40880338, 32'hc066e11e} /* (28, 18, 28) {real, imag} */,
  {32'h3f3b9da0, 32'hc11edaaf} /* (28, 18, 27) {real, imag} */,
  {32'h3f9e2af8, 32'hc0bbdab8} /* (28, 18, 26) {real, imag} */,
  {32'hbf813340, 32'hc0496f52} /* (28, 18, 25) {real, imag} */,
  {32'h408457be, 32'hbdb82d80} /* (28, 18, 24) {real, imag} */,
  {32'h40930054, 32'h3f188798} /* (28, 18, 23) {real, imag} */,
  {32'h401fbee2, 32'hbfa2f7cf} /* (28, 18, 22) {real, imag} */,
  {32'hbf6c3224, 32'hc04085e0} /* (28, 18, 21) {real, imag} */,
  {32'h3cae0c00, 32'h3e16f560} /* (28, 18, 20) {real, imag} */,
  {32'h3e29ec40, 32'h3da31980} /* (28, 18, 19) {real, imag} */,
  {32'hc0b8b61c, 32'h3e2e3140} /* (28, 18, 18) {real, imag} */,
  {32'hc0b447c2, 32'h40210d44} /* (28, 18, 17) {real, imag} */,
  {32'hbf471240, 32'h3d7654c0} /* (28, 18, 16) {real, imag} */,
  {32'h40702750, 32'h40c73bad} /* (28, 18, 15) {real, imag} */,
  {32'hc0f963ec, 32'h3fb41c00} /* (28, 18, 14) {real, imag} */,
  {32'hc163c985, 32'h3f5912b0} /* (28, 18, 13) {real, imag} */,
  {32'hc0d9a56a, 32'hc01083c7} /* (28, 18, 12) {real, imag} */,
  {32'hc0a645b9, 32'hc091cd8e} /* (28, 18, 11) {real, imag} */,
  {32'hc0725f4a, 32'hbf2c3d90} /* (28, 18, 10) {real, imag} */,
  {32'h3fa1c24c, 32'hbf9fd5d0} /* (28, 18, 9) {real, imag} */,
  {32'h3fdd61c8, 32'hbfa74ae4} /* (28, 18, 8) {real, imag} */,
  {32'h409b72f0, 32'hbf2ab184} /* (28, 18, 7) {real, imag} */,
  {32'h404c8222, 32'h3eb1d628} /* (28, 18, 6) {real, imag} */,
  {32'h409795ca, 32'h3ee2107c} /* (28, 18, 5) {real, imag} */,
  {32'h408ba608, 32'hc02db0c8} /* (28, 18, 4) {real, imag} */,
  {32'h4014787c, 32'h4004e69a} /* (28, 18, 3) {real, imag} */,
  {32'h40794520, 32'h3ff3077c} /* (28, 18, 2) {real, imag} */,
  {32'h40a2edff, 32'h400bc051} /* (28, 18, 1) {real, imag} */,
  {32'h40c84028, 32'h3f2e2f34} /* (28, 18, 0) {real, imag} */,
  {32'hbfd04726, 32'hc01bdee3} /* (28, 17, 31) {real, imag} */,
  {32'hc0d4cb02, 32'hbf5b4b20} /* (28, 17, 30) {real, imag} */,
  {32'hc00389b8, 32'h405558f4} /* (28, 17, 29) {real, imag} */,
  {32'h40d618f0, 32'h3f0f0ee4} /* (28, 17, 28) {real, imag} */,
  {32'hbf0aa858, 32'hc09eb210} /* (28, 17, 27) {real, imag} */,
  {32'hc0b49b07, 32'hc0644ca8} /* (28, 17, 26) {real, imag} */,
  {32'hc0291d6c, 32'h40796ec5} /* (28, 17, 25) {real, imag} */,
  {32'hc08006b8, 32'h40947745} /* (28, 17, 24) {real, imag} */,
  {32'hbfe333d8, 32'hbf1f41d0} /* (28, 17, 23) {real, imag} */,
  {32'h3f0224e0, 32'hc01b35da} /* (28, 17, 22) {real, imag} */,
  {32'hbe43e120, 32'hc03e7b48} /* (28, 17, 21) {real, imag} */,
  {32'h3f9038d6, 32'h3fa82b48} /* (28, 17, 20) {real, imag} */,
  {32'h41049afa, 32'h3ff90d84} /* (28, 17, 19) {real, imag} */,
  {32'h4084e1a6, 32'hc00fcb00} /* (28, 17, 18) {real, imag} */,
  {32'hbf4d911c, 32'hc0027f84} /* (28, 17, 17) {real, imag} */,
  {32'h40b59d52, 32'hc01b9cb0} /* (28, 17, 16) {real, imag} */,
  {32'h40aef980, 32'h3edb5a40} /* (28, 17, 15) {real, imag} */,
  {32'h405744e4, 32'h404c2577} /* (28, 17, 14) {real, imag} */,
  {32'h403edc40, 32'h4052acfe} /* (28, 17, 13) {real, imag} */,
  {32'hc00d035d, 32'h3febee78} /* (28, 17, 12) {real, imag} */,
  {32'hc05252aa, 32'h406cb9ca} /* (28, 17, 11) {real, imag} */,
  {32'hc05b9a6f, 32'h3f3c2ce0} /* (28, 17, 10) {real, imag} */,
  {32'hc107d2b4, 32'h4026fdfc} /* (28, 17, 9) {real, imag} */,
  {32'hc00bf83c, 32'h405e3514} /* (28, 17, 8) {real, imag} */,
  {32'h40ba5850, 32'h403fb79a} /* (28, 17, 7) {real, imag} */,
  {32'h40538654, 32'h3edb5980} /* (28, 17, 6) {real, imag} */,
  {32'h3fc5bfa8, 32'h404797fb} /* (28, 17, 5) {real, imag} */,
  {32'h3e880f58, 32'h40a8b76d} /* (28, 17, 4) {real, imag} */,
  {32'hc0ccc4c8, 32'hc09da720} /* (28, 17, 3) {real, imag} */,
  {32'hc107091e, 32'hc11f8140} /* (28, 17, 2) {real, imag} */,
  {32'hc0b41efa, 32'hc01b2ef5} /* (28, 17, 1) {real, imag} */,
  {32'hbf740a42, 32'hbf879462} /* (28, 17, 0) {real, imag} */,
  {32'hc008fd66, 32'h3f8dfea0} /* (28, 16, 31) {real, imag} */,
  {32'h40706600, 32'hbfd7c220} /* (28, 16, 30) {real, imag} */,
  {32'h40b86172, 32'hc0bbaed0} /* (28, 16, 29) {real, imag} */,
  {32'h40a41d1e, 32'hc10a34c4} /* (28, 16, 28) {real, imag} */,
  {32'h40410668, 32'hc0347480} /* (28, 16, 27) {real, imag} */,
  {32'hbf81e4c0, 32'hbf027c00} /* (28, 16, 26) {real, imag} */,
  {32'hbfda7838, 32'hbf0bf7e0} /* (28, 16, 25) {real, imag} */,
  {32'h3fd3c3e2, 32'h4092b914} /* (28, 16, 24) {real, imag} */,
  {32'h4031017a, 32'hbeb62d80} /* (28, 16, 23) {real, imag} */,
  {32'h3fbf94b0, 32'h3f700600} /* (28, 16, 22) {real, imag} */,
  {32'hc0ae1ebc, 32'hc0503770} /* (28, 16, 21) {real, imag} */,
  {32'hc09d93f2, 32'hc10381a6} /* (28, 16, 20) {real, imag} */,
  {32'hc10bdb54, 32'hc0a62d9c} /* (28, 16, 19) {real, imag} */,
  {32'hbfce4260, 32'hc0835344} /* (28, 16, 18) {real, imag} */,
  {32'h40778792, 32'h3fda842c} /* (28, 16, 17) {real, imag} */,
  {32'h4010345a, 32'h406f69f2} /* (28, 16, 16) {real, imag} */,
  {32'h3eb9927c, 32'hbf3593e0} /* (28, 16, 15) {real, imag} */,
  {32'hbfc33190, 32'h3e1d4680} /* (28, 16, 14) {real, imag} */,
  {32'hbfc67dd0, 32'hc01c4f20} /* (28, 16, 13) {real, imag} */,
  {32'h3fe783c8, 32'hc0742cf0} /* (28, 16, 12) {real, imag} */,
  {32'h3f638f30, 32'hc0812390} /* (28, 16, 11) {real, imag} */,
  {32'h40409475, 32'hc03bce10} /* (28, 16, 10) {real, imag} */,
  {32'hbf2bdf20, 32'hbf63dd90} /* (28, 16, 9) {real, imag} */,
  {32'hbfdd7a0c, 32'hc034fae4} /* (28, 16, 8) {real, imag} */,
  {32'hc0b18759, 32'hbf752a20} /* (28, 16, 7) {real, imag} */,
  {32'h3df7ff00, 32'hbf6d1ae0} /* (28, 16, 6) {real, imag} */,
  {32'h40909c9d, 32'hc00d5230} /* (28, 16, 5) {real, imag} */,
  {32'hbe61ed00, 32'hbe505f00} /* (28, 16, 4) {real, imag} */,
  {32'h3cf98100, 32'hc001c580} /* (28, 16, 3) {real, imag} */,
  {32'h40a751ae, 32'hbf884cb0} /* (28, 16, 2) {real, imag} */,
  {32'h409018d0, 32'hbfcaf120} /* (28, 16, 1) {real, imag} */,
  {32'hbf4a57e0, 32'hc05ffc9c} /* (28, 16, 0) {real, imag} */,
  {32'h4005f58f, 32'h407576c3} /* (28, 15, 31) {real, imag} */,
  {32'h40faf4ba, 32'h3ff0fa90} /* (28, 15, 30) {real, imag} */,
  {32'h40474608, 32'hc0a73a9a} /* (28, 15, 29) {real, imag} */,
  {32'h3f058ce0, 32'hc084e21c} /* (28, 15, 28) {real, imag} */,
  {32'h3fae0c2c, 32'h402789bf} /* (28, 15, 27) {real, imag} */,
  {32'hc00f1e7a, 32'h40156328} /* (28, 15, 26) {real, imag} */,
  {32'hc013f794, 32'hbe947d28} /* (28, 15, 25) {real, imag} */,
  {32'hc09d5758, 32'hbf98aad4} /* (28, 15, 24) {real, imag} */,
  {32'hc03f9814, 32'h3fba0fe8} /* (28, 15, 23) {real, imag} */,
  {32'hc099cb3c, 32'h3f7b4768} /* (28, 15, 22) {real, imag} */,
  {32'hc02814be, 32'hbdcefb00} /* (28, 15, 21) {real, imag} */,
  {32'hc0659391, 32'hbf46d190} /* (28, 15, 20) {real, imag} */,
  {32'h3e954350, 32'hbe591a20} /* (28, 15, 19) {real, imag} */,
  {32'h40862b76, 32'h40e7d6f8} /* (28, 15, 18) {real, imag} */,
  {32'h404d5c09, 32'h3fd7eb08} /* (28, 15, 17) {real, imag} */,
  {32'hbf7b20ec, 32'h40004560} /* (28, 15, 16) {real, imag} */,
  {32'hc08c8de6, 32'h40a6aac4} /* (28, 15, 15) {real, imag} */,
  {32'hc0913916, 32'h3fdb0b12} /* (28, 15, 14) {real, imag} */,
  {32'hc081ce84, 32'h40249242} /* (28, 15, 13) {real, imag} */,
  {32'hbfcd0076, 32'h3f84f7c8} /* (28, 15, 12) {real, imag} */,
  {32'hbdf69fb0, 32'hbf9db254} /* (28, 15, 11) {real, imag} */,
  {32'hbfe4a60e, 32'h41118eb7} /* (28, 15, 10) {real, imag} */,
  {32'h3fdfcca0, 32'h4066fb0c} /* (28, 15, 9) {real, imag} */,
  {32'h40618204, 32'hc034db74} /* (28, 15, 8) {real, imag} */,
  {32'h40859ad8, 32'h401efbd6} /* (28, 15, 7) {real, imag} */,
  {32'h40ad7ce6, 32'h406982d0} /* (28, 15, 6) {real, imag} */,
  {32'hbf602cd0, 32'h40e03f2a} /* (28, 15, 5) {real, imag} */,
  {32'hc0a88776, 32'hbf1a8068} /* (28, 15, 4) {real, imag} */,
  {32'hc019bea8, 32'hc0825510} /* (28, 15, 3) {real, imag} */,
  {32'hc0177c88, 32'hc081293f} /* (28, 15, 2) {real, imag} */,
  {32'hbf50b3bc, 32'hbf9511d6} /* (28, 15, 1) {real, imag} */,
  {32'h40091570, 32'h3f7302c4} /* (28, 15, 0) {real, imag} */,
  {32'hbf3c7fb8, 32'hbf08a1dc} /* (28, 14, 31) {real, imag} */,
  {32'hbc994a00, 32'hbfa2aada} /* (28, 14, 30) {real, imag} */,
  {32'hc0d5ee04, 32'h3f82c692} /* (28, 14, 29) {real, imag} */,
  {32'hc13ec7ec, 32'h3f9e883c} /* (28, 14, 28) {real, imag} */,
  {32'hc08236c8, 32'hc0131745} /* (28, 14, 27) {real, imag} */,
  {32'h3fbbf828, 32'hc0802a70} /* (28, 14, 26) {real, imag} */,
  {32'hc008aa40, 32'h3e67bd20} /* (28, 14, 25) {real, imag} */,
  {32'hc02457fc, 32'h40554abc} /* (28, 14, 24) {real, imag} */,
  {32'hc02d7b18, 32'hbfe8b4ac} /* (28, 14, 23) {real, imag} */,
  {32'h40901f47, 32'hc09898fc} /* (28, 14, 22) {real, imag} */,
  {32'h40bf9c02, 32'hbfb103a8} /* (28, 14, 21) {real, imag} */,
  {32'hbe0abb80, 32'hc02575b6} /* (28, 14, 20) {real, imag} */,
  {32'hc0b0774e, 32'h3ffc9a08} /* (28, 14, 19) {real, imag} */,
  {32'hbf13aea0, 32'hbf429390} /* (28, 14, 18) {real, imag} */,
  {32'h4054e3ec, 32'hc10602b9} /* (28, 14, 17) {real, imag} */,
  {32'h40034b90, 32'hc00702a3} /* (28, 14, 16) {real, imag} */,
  {32'h401c7900, 32'h404d10f6} /* (28, 14, 15) {real, imag} */,
  {32'h40424a8c, 32'h40384120} /* (28, 14, 14) {real, imag} */,
  {32'hc097f6de, 32'hbdda7d80} /* (28, 14, 13) {real, imag} */,
  {32'hc0d65320, 32'h3fb09c6e} /* (28, 14, 12) {real, imag} */,
  {32'hc024a242, 32'hbfdead38} /* (28, 14, 11) {real, imag} */,
  {32'hc0494b32, 32'h4078d344} /* (28, 14, 10) {real, imag} */,
  {32'hc0bdb3ab, 32'h4115a46a} /* (28, 14, 9) {real, imag} */,
  {32'hc0cda7c6, 32'h40dd21b9} /* (28, 14, 8) {real, imag} */,
  {32'hc02743b0, 32'h40c078c0} /* (28, 14, 7) {real, imag} */,
  {32'hbfc3504c, 32'h40c5f61e} /* (28, 14, 6) {real, imag} */,
  {32'h403a9cdc, 32'h404d2b00} /* (28, 14, 5) {real, imag} */,
  {32'hc02435a0, 32'h3f8839b0} /* (28, 14, 4) {real, imag} */,
  {32'hc0b38694, 32'h4088cff3} /* (28, 14, 3) {real, imag} */,
  {32'hc0505e20, 32'h40ec5ff9} /* (28, 14, 2) {real, imag} */,
  {32'h40b8f16d, 32'h3f9aaede} /* (28, 14, 1) {real, imag} */,
  {32'h3fd53f00, 32'h3d8b4660} /* (28, 14, 0) {real, imag} */,
  {32'h3fe2288c, 32'hc05301a1} /* (28, 13, 31) {real, imag} */,
  {32'hc010d2e0, 32'h4048a339} /* (28, 13, 30) {real, imag} */,
  {32'hc0bb869c, 32'h402045a7} /* (28, 13, 29) {real, imag} */,
  {32'h40533cee, 32'hbe2dc630} /* (28, 13, 28) {real, imag} */,
  {32'hc025fce4, 32'h3f8c90bc} /* (28, 13, 27) {real, imag} */,
  {32'hbf5fef20, 32'hbf9ede74} /* (28, 13, 26) {real, imag} */,
  {32'h3fab6ed8, 32'hc05f86af} /* (28, 13, 25) {real, imag} */,
  {32'h400df145, 32'hc05fb924} /* (28, 13, 24) {real, imag} */,
  {32'h3f6521e0, 32'h408369fe} /* (28, 13, 23) {real, imag} */,
  {32'h3ff21910, 32'hbf851ef6} /* (28, 13, 22) {real, imag} */,
  {32'h40c2d760, 32'h3def7700} /* (28, 13, 21) {real, imag} */,
  {32'h40da115a, 32'h4056174d} /* (28, 13, 20) {real, imag} */,
  {32'h40b3e042, 32'h409930f7} /* (28, 13, 19) {real, imag} */,
  {32'h3ec18a60, 32'h403ce480} /* (28, 13, 18) {real, imag} */,
  {32'hc018c038, 32'h3f0c5194} /* (28, 13, 17) {real, imag} */,
  {32'hbf9bed00, 32'hc0ac0bdd} /* (28, 13, 16) {real, imag} */,
  {32'hc1037a2a, 32'hc07a1e54} /* (28, 13, 15) {real, imag} */,
  {32'hc11ef7df, 32'h3fd0b3cd} /* (28, 13, 14) {real, imag} */,
  {32'hbd6e2680, 32'h412e57c0} /* (28, 13, 13) {real, imag} */,
  {32'h40cc039c, 32'h3f903bf8} /* (28, 13, 12) {real, imag} */,
  {32'h40c54bd6, 32'hbfb9f1f2} /* (28, 13, 11) {real, imag} */,
  {32'h4103c4c4, 32'h3ebf5020} /* (28, 13, 10) {real, imag} */,
  {32'h40a22093, 32'hc09394b9} /* (28, 13, 9) {real, imag} */,
  {32'h40a6c15a, 32'hc0cc8d34} /* (28, 13, 8) {real, imag} */,
  {32'hbf1e6b40, 32'hbe72e6f0} /* (28, 13, 7) {real, imag} */,
  {32'h3facd7f4, 32'hbf563160} /* (28, 13, 6) {real, imag} */,
  {32'h4119025a, 32'hbe41bf50} /* (28, 13, 5) {real, imag} */,
  {32'h408e1319, 32'hbe9d3818} /* (28, 13, 4) {real, imag} */,
  {32'hbe8231e0, 32'hc0d6aa50} /* (28, 13, 3) {real, imag} */,
  {32'h402e5f84, 32'hc0b9bcea} /* (28, 13, 2) {real, imag} */,
  {32'h402daae9, 32'h3f93595e} /* (28, 13, 1) {real, imag} */,
  {32'h3f7fbc48, 32'h406e4eec} /* (28, 13, 0) {real, imag} */,
  {32'h40cbaa4b, 32'hc0b224b2} /* (28, 12, 31) {real, imag} */,
  {32'h40ca71de, 32'h3fb38190} /* (28, 12, 30) {real, imag} */,
  {32'h40b8917b, 32'h411b1c48} /* (28, 12, 29) {real, imag} */,
  {32'h3f5666c0, 32'h410b85ea} /* (28, 12, 28) {real, imag} */,
  {32'hc01843f5, 32'h409862be} /* (28, 12, 27) {real, imag} */,
  {32'hc0110cd2, 32'h3eb28410} /* (28, 12, 26) {real, imag} */,
  {32'hc02b5bcf, 32'h3ffd462c} /* (28, 12, 25) {real, imag} */,
  {32'hc0cbf84e, 32'hc09ba372} /* (28, 12, 24) {real, imag} */,
  {32'h3fad6624, 32'hc10f2538} /* (28, 12, 23) {real, imag} */,
  {32'hc09cd734, 32'hc09fe098} /* (28, 12, 22) {real, imag} */,
  {32'hc14b033f, 32'hc06f4147} /* (28, 12, 21) {real, imag} */,
  {32'hc02f2db6, 32'hc0a8cede} /* (28, 12, 20) {real, imag} */,
  {32'h40fb7206, 32'hc006ad5b} /* (28, 12, 19) {real, imag} */,
  {32'h40e41ff4, 32'hc06c6c10} /* (28, 12, 18) {real, imag} */,
  {32'h410c257a, 32'h3f5b9820} /* (28, 12, 17) {real, imag} */,
  {32'h40cbbe30, 32'h40b11115} /* (28, 12, 16) {real, imag} */,
  {32'h40173f7a, 32'hbf0deaca} /* (28, 12, 15) {real, imag} */,
  {32'h40858f73, 32'h4090933c} /* (28, 12, 14) {real, imag} */,
  {32'hc07851d4, 32'h411d11ad} /* (28, 12, 13) {real, imag} */,
  {32'h3f5494b0, 32'h4087e8d1} /* (28, 12, 12) {real, imag} */,
  {32'h41026458, 32'hbffed063} /* (28, 12, 11) {real, imag} */,
  {32'h40191cba, 32'h40e0909d} /* (28, 12, 10) {real, imag} */,
  {32'hc0f8c11b, 32'h4139e2f5} /* (28, 12, 9) {real, imag} */,
  {32'hc0a0b12e, 32'h4004813c} /* (28, 12, 8) {real, imag} */,
  {32'hc0e4c25a, 32'h401704fc} /* (28, 12, 7) {real, imag} */,
  {32'h402bc0b8, 32'hc0412102} /* (28, 12, 6) {real, imag} */,
  {32'h40efe4a4, 32'h3f30c564} /* (28, 12, 5) {real, imag} */,
  {32'h4105cecc, 32'h400a7962} /* (28, 12, 4) {real, imag} */,
  {32'h3fb7969c, 32'hc02dda74} /* (28, 12, 3) {real, imag} */,
  {32'hc01b4c40, 32'hc059bcdc} /* (28, 12, 2) {real, imag} */,
  {32'h406ecfc1, 32'hbff812f8} /* (28, 12, 1) {real, imag} */,
  {32'h4038f9f4, 32'hc025ba72} /* (28, 12, 0) {real, imag} */,
  {32'h3f9db4fa, 32'h40889132} /* (28, 11, 31) {real, imag} */,
  {32'hbf7d8558, 32'h405b9cf4} /* (28, 11, 30) {real, imag} */,
  {32'hc0f19d0d, 32'h40c42683} /* (28, 11, 29) {real, imag} */,
  {32'hc0e492b1, 32'h4145b960} /* (28, 11, 28) {real, imag} */,
  {32'hc119b646, 32'h40a4c520} /* (28, 11, 27) {real, imag} */,
  {32'hc10900b5, 32'h3faa8640} /* (28, 11, 26) {real, imag} */,
  {32'hc0f99714, 32'hbfb7a7ac} /* (28, 11, 25) {real, imag} */,
  {32'hc0c96d32, 32'h4046945c} /* (28, 11, 24) {real, imag} */,
  {32'hc13bb531, 32'h40e763c6} /* (28, 11, 23) {real, imag} */,
  {32'hc152931c, 32'h409ef7d2} /* (28, 11, 22) {real, imag} */,
  {32'hc0e65420, 32'h3f78af90} /* (28, 11, 21) {real, imag} */,
  {32'hc04810df, 32'h40923a8d} /* (28, 11, 20) {real, imag} */,
  {32'hc0f02be2, 32'h3f3b6a80} /* (28, 11, 19) {real, imag} */,
  {32'hbfd3eb80, 32'hbff88a24} /* (28, 11, 18) {real, imag} */,
  {32'h406dd9f0, 32'hbf494500} /* (28, 11, 17) {real, imag} */,
  {32'h4134472d, 32'h40b8af6f} /* (28, 11, 16) {real, imag} */,
  {32'h414b3481, 32'hbf9a0559} /* (28, 11, 15) {real, imag} */,
  {32'h413559d7, 32'hc119a135} /* (28, 11, 14) {real, imag} */,
  {32'hc02195ba, 32'hc10947b0} /* (28, 11, 13) {real, imag} */,
  {32'hc02fc332, 32'hc12e87ea} /* (28, 11, 12) {real, imag} */,
  {32'h407fa477, 32'hc0b977db} /* (28, 11, 11) {real, imag} */,
  {32'hc0f34c6b, 32'h3fb3edc8} /* (28, 11, 10) {real, imag} */,
  {32'hc191afa8, 32'h4124ee1a} /* (28, 11, 9) {real, imag} */,
  {32'hc1789cb9, 32'h40e07db5} /* (28, 11, 8) {real, imag} */,
  {32'hc16e9d4c, 32'h4098c7c1} /* (28, 11, 7) {real, imag} */,
  {32'hc01e3db5, 32'h4054ed36} /* (28, 11, 6) {real, imag} */,
  {32'h3fbc7aea, 32'hc08fc14a} /* (28, 11, 5) {real, imag} */,
  {32'hc01e7fe2, 32'h403d567a} /* (28, 11, 4) {real, imag} */,
  {32'hbf893a24, 32'h40d4dc68} /* (28, 11, 3) {real, imag} */,
  {32'h408aca15, 32'h3f05a2a0} /* (28, 11, 2) {real, imag} */,
  {32'h407e5940, 32'hc083c803} /* (28, 11, 1) {real, imag} */,
  {32'h408181d9, 32'h3fb9408e} /* (28, 11, 0) {real, imag} */,
  {32'hc067901d, 32'hbfcbc264} /* (28, 10, 31) {real, imag} */,
  {32'hbed8e180, 32'h40d20ee6} /* (28, 10, 30) {real, imag} */,
  {32'h40e31a4c, 32'hc035ce8c} /* (28, 10, 29) {real, imag} */,
  {32'h40a74f64, 32'hbf140868} /* (28, 10, 28) {real, imag} */,
  {32'h41020027, 32'hbfd7a632} /* (28, 10, 27) {real, imag} */,
  {32'hbf7dfca0, 32'hbf1f7dd4} /* (28, 10, 26) {real, imag} */,
  {32'hbe8671e8, 32'hbf7bba80} /* (28, 10, 25) {real, imag} */,
  {32'h4033dcdc, 32'hc0a46698} /* (28, 10, 24) {real, imag} */,
  {32'hc027820b, 32'hbfed9eca} /* (28, 10, 23) {real, imag} */,
  {32'h409f7e34, 32'hc07687af} /* (28, 10, 22) {real, imag} */,
  {32'h401152d4, 32'h3dce85a0} /* (28, 10, 21) {real, imag} */,
  {32'h407ced1c, 32'h4138241a} /* (28, 10, 20) {real, imag} */,
  {32'h41149639, 32'h40d5f748} /* (28, 10, 19) {real, imag} */,
  {32'h411fab8b, 32'h40cd9373} /* (28, 10, 18) {real, imag} */,
  {32'hbfbf45fc, 32'h4148d3ee} /* (28, 10, 17) {real, imag} */,
  {32'hc0b75932, 32'h41a95224} /* (28, 10, 16) {real, imag} */,
  {32'h4065b879, 32'h413221d6} /* (28, 10, 15) {real, imag} */,
  {32'hc00f74c8, 32'h413146f4} /* (28, 10, 14) {real, imag} */,
  {32'h3f90459e, 32'h415921dc} /* (28, 10, 13) {real, imag} */,
  {32'hc0bac51b, 32'h415077e4} /* (28, 10, 12) {real, imag} */,
  {32'h3fb3a65e, 32'h412335a7} /* (28, 10, 11) {real, imag} */,
  {32'h41704ce7, 32'h40439e31} /* (28, 10, 10) {real, imag} */,
  {32'h40fe0ba2, 32'hc0ea4f52} /* (28, 10, 9) {real, imag} */,
  {32'h40b33f62, 32'hc10eeb7a} /* (28, 10, 8) {real, imag} */,
  {32'h40fb3cd2, 32'hc0cde41c} /* (28, 10, 7) {real, imag} */,
  {32'h40857630, 32'h40cbab0e} /* (28, 10, 6) {real, imag} */,
  {32'h4182763c, 32'h406873a8} /* (28, 10, 5) {real, imag} */,
  {32'h4149bb1f, 32'h4029dda4} /* (28, 10, 4) {real, imag} */,
  {32'h40ae55de, 32'h401ea718} /* (28, 10, 3) {real, imag} */,
  {32'hc0ecfaa8, 32'h40e4bca8} /* (28, 10, 2) {real, imag} */,
  {32'hc119411a, 32'h40fbb7af} /* (28, 10, 1) {real, imag} */,
  {32'hc0a2417a, 32'hc062e5c8} /* (28, 10, 0) {real, imag} */,
  {32'hc00300c1, 32'h40750d87} /* (28, 9, 31) {real, imag} */,
  {32'hbf34e430, 32'h409ee20b} /* (28, 9, 30) {real, imag} */,
  {32'hbfaf13b8, 32'hc0179edb} /* (28, 9, 29) {real, imag} */,
  {32'h3fae54c4, 32'hc10ba347} /* (28, 9, 28) {real, imag} */,
  {32'h41467aa0, 32'hc1caa9c5} /* (28, 9, 27) {real, imag} */,
  {32'h41aeb01c, 32'hc10564bd} /* (28, 9, 26) {real, imag} */,
  {32'h4181b745, 32'h408cf028} /* (28, 9, 25) {real, imag} */,
  {32'h4140fad7, 32'hc10c817c} /* (28, 9, 24) {real, imag} */,
  {32'h4005329e, 32'hc03a94e0} /* (28, 9, 23) {real, imag} */,
  {32'h40a3e75f, 32'h3fbd59d4} /* (28, 9, 22) {real, imag} */,
  {32'h409de04d, 32'h3f828f90} /* (28, 9, 21) {real, imag} */,
  {32'hc0c16718, 32'h412b0998} /* (28, 9, 20) {real, imag} */,
  {32'hc1731ebd, 32'h40eedb5f} /* (28, 9, 19) {real, imag} */,
  {32'hc1acfafc, 32'h40546964} /* (28, 9, 18) {real, imag} */,
  {32'hc17e0669, 32'hbf94cfa8} /* (28, 9, 17) {real, imag} */,
  {32'h41078eee, 32'hbe0c0e40} /* (28, 9, 16) {real, imag} */,
  {32'h413e4a9a, 32'hbeb96680} /* (28, 9, 15) {real, imag} */,
  {32'hbff04310, 32'hc0c734aa} /* (28, 9, 14) {real, imag} */,
  {32'hc02366e3, 32'h3e491220} /* (28, 9, 13) {real, imag} */,
  {32'h3e5840e0, 32'h41002787} /* (28, 9, 12) {real, imag} */,
  {32'hc0ffea34, 32'hbf8fa9c6} /* (28, 9, 11) {real, imag} */,
  {32'h40844dd9, 32'hc0b118af} /* (28, 9, 10) {real, imag} */,
  {32'h41532aed, 32'hc02c8f64} /* (28, 9, 9) {real, imag} */,
  {32'h4179d391, 32'hc11a124d} /* (28, 9, 8) {real, imag} */,
  {32'h413f7f5a, 32'hc17c3055} /* (28, 9, 7) {real, imag} */,
  {32'hc0ad06c2, 32'h3e07e3a0} /* (28, 9, 6) {real, imag} */,
  {32'hc103e1c7, 32'h3ff27620} /* (28, 9, 5) {real, imag} */,
  {32'hc0d0aa7a, 32'hbf554040} /* (28, 9, 4) {real, imag} */,
  {32'h3ff89d86, 32'h40d2b558} /* (28, 9, 3) {real, imag} */,
  {32'hc069d310, 32'h40a2b18c} /* (28, 9, 2) {real, imag} */,
  {32'h3fb63970, 32'hc10b0628} /* (28, 9, 1) {real, imag} */,
  {32'h40685f4d, 32'hc0b09bd0} /* (28, 9, 0) {real, imag} */,
  {32'h3fb99f3c, 32'h40b46a33} /* (28, 8, 31) {real, imag} */,
  {32'hbfa6bcf0, 32'h417f14b4} /* (28, 8, 30) {real, imag} */,
  {32'hc0284a70, 32'h41a96c51} /* (28, 8, 29) {real, imag} */,
  {32'h4015ef0c, 32'h4136d2b1} /* (28, 8, 28) {real, imag} */,
  {32'hc13a9272, 32'h4178a52f} /* (28, 8, 27) {real, imag} */,
  {32'h3e4c6d00, 32'h41237bec} /* (28, 8, 26) {real, imag} */,
  {32'h40e47438, 32'h41596414} /* (28, 8, 25) {real, imag} */,
  {32'hc0edd9c4, 32'h41a4e2da} /* (28, 8, 24) {real, imag} */,
  {32'hc16f4c7a, 32'h40a6c792} /* (28, 8, 23) {real, imag} */,
  {32'hc082d1e0, 32'h41080be2} /* (28, 8, 22) {real, imag} */,
  {32'hc12441b9, 32'h40b54b5c} /* (28, 8, 21) {real, imag} */,
  {32'hc157f427, 32'hc12950fb} /* (28, 8, 20) {real, imag} */,
  {32'h40462fa8, 32'h4066c86e} /* (28, 8, 19) {real, imag} */,
  {32'h40eb1c40, 32'h4164a956} /* (28, 8, 18) {real, imag} */,
  {32'h40278310, 32'hc0eef661} /* (28, 8, 17) {real, imag} */,
  {32'hc0b0e2f1, 32'hc1b6a9ed} /* (28, 8, 16) {real, imag} */,
  {32'h3f4d951c, 32'hc1ec1b6c} /* (28, 8, 15) {real, imag} */,
  {32'h411615b0, 32'hc0d1c69d} /* (28, 8, 14) {real, imag} */,
  {32'h40f6a3cc, 32'hc0c397f4} /* (28, 8, 13) {real, imag} */,
  {32'h40616290, 32'hc1c485be} /* (28, 8, 12) {real, imag} */,
  {32'hbfb3dd78, 32'hc14fe77d} /* (28, 8, 11) {real, imag} */,
  {32'hbf24b6a0, 32'hbeb7f930} /* (28, 8, 10) {real, imag} */,
  {32'h3db7f640, 32'h41310208} /* (28, 8, 9) {real, imag} */,
  {32'hc08273f4, 32'h41ea7017} /* (28, 8, 8) {real, imag} */,
  {32'hc0d99600, 32'h41d5c040} /* (28, 8, 7) {real, imag} */,
  {32'h4096347d, 32'h4201eb30} /* (28, 8, 6) {real, imag} */,
  {32'hc082f92b, 32'h41f1145a} /* (28, 8, 5) {real, imag} */,
  {32'hc0edd894, 32'h412247ac} /* (28, 8, 4) {real, imag} */,
  {32'hc0fac199, 32'h4164838e} /* (28, 8, 3) {real, imag} */,
  {32'hc1a1682c, 32'h4199ea2a} /* (28, 8, 2) {real, imag} */,
  {32'hc198ae9a, 32'h41aba7ce} /* (28, 8, 1) {real, imag} */,
  {32'hc114b508, 32'h41655a56} /* (28, 8, 0) {real, imag} */,
  {32'hc0de3b8a, 32'h3ffd69a2} /* (28, 7, 31) {real, imag} */,
  {32'hc18d5c86, 32'h406f30c2} /* (28, 7, 30) {real, imag} */,
  {32'hc0b650fe, 32'hc0edc08a} /* (28, 7, 29) {real, imag} */,
  {32'h3f780bd0, 32'hc0372f88} /* (28, 7, 28) {real, imag} */,
  {32'h40bd25ef, 32'h416a7e4e} /* (28, 7, 27) {real, imag} */,
  {32'hc13b3172, 32'h415e7277} /* (28, 7, 26) {real, imag} */,
  {32'hc0b21a5b, 32'h413cee39} /* (28, 7, 25) {real, imag} */,
  {32'hbf99dbc8, 32'h413ebe5e} /* (28, 7, 24) {real, imag} */,
  {32'h41121574, 32'h405e6df0} /* (28, 7, 23) {real, imag} */,
  {32'hc0018c5c, 32'hc12ceaee} /* (28, 7, 22) {real, imag} */,
  {32'h3fa96fc0, 32'hc087f96c} /* (28, 7, 21) {real, imag} */,
  {32'h41ab0f4b, 32'hc16bacaf} /* (28, 7, 20) {real, imag} */,
  {32'h40a7285d, 32'hc1436fbc} /* (28, 7, 19) {real, imag} */,
  {32'hc0566474, 32'hc18a6272} /* (28, 7, 18) {real, imag} */,
  {32'h418d5469, 32'hc14414f7} /* (28, 7, 17) {real, imag} */,
  {32'h41471432, 32'h4099c482} /* (28, 7, 16) {real, imag} */,
  {32'h4079dda6, 32'h404faad2} /* (28, 7, 15) {real, imag} */,
  {32'hc126f450, 32'hc11a9fd3} /* (28, 7, 14) {real, imag} */,
  {32'hc13096f4, 32'hc186f3d7} /* (28, 7, 13) {real, imag} */,
  {32'hc085090c, 32'hbfbd7224} /* (28, 7, 12) {real, imag} */,
  {32'hc0c31130, 32'h41785e0d} /* (28, 7, 11) {real, imag} */,
  {32'h3ef84a41, 32'h41cb958b} /* (28, 7, 10) {real, imag} */,
  {32'h4118e2f1, 32'h419d7cf2} /* (28, 7, 9) {real, imag} */,
  {32'h40e3faee, 32'h41629ea4} /* (28, 7, 8) {real, imag} */,
  {32'h4154bf18, 32'h4085ca30} /* (28, 7, 7) {real, imag} */,
  {32'h40bdd5fa, 32'hc12ac1f2} /* (28, 7, 6) {real, imag} */,
  {32'hc0070930, 32'hc1c91c84} /* (28, 7, 5) {real, imag} */,
  {32'h3fde3a28, 32'hc13c1770} /* (28, 7, 4) {real, imag} */,
  {32'hbe7218c0, 32'h40def794} /* (28, 7, 3) {real, imag} */,
  {32'h409dfd40, 32'hc122cd56} /* (28, 7, 2) {real, imag} */,
  {32'hc0075e40, 32'hc06f0611} /* (28, 7, 1) {real, imag} */,
  {32'hc08530bb, 32'hc0a4c822} /* (28, 7, 0) {real, imag} */,
  {32'h3fe64d18, 32'hc094fb12} /* (28, 6, 31) {real, imag} */,
  {32'hbfa30400, 32'hc0eff7a5} /* (28, 6, 30) {real, imag} */,
  {32'hc0f7f208, 32'hc184cda9} /* (28, 6, 29) {real, imag} */,
  {32'h3fd72b80, 32'hc1a2033e} /* (28, 6, 28) {real, imag} */,
  {32'h417cea49, 32'hc066fd7f} /* (28, 6, 27) {real, imag} */,
  {32'h413f20a6, 32'h41b33cb9} /* (28, 6, 26) {real, imag} */,
  {32'h417bf095, 32'hc0c68d68} /* (28, 6, 25) {real, imag} */,
  {32'h41466d6b, 32'hc11fb678} /* (28, 6, 24) {real, imag} */,
  {32'hbfa09c28, 32'h40c99be8} /* (28, 6, 23) {real, imag} */,
  {32'hc197c4c7, 32'h4180eade} /* (28, 6, 22) {real, imag} */,
  {32'hc17c0204, 32'h40412658} /* (28, 6, 21) {real, imag} */,
  {32'hc0bdaa5c, 32'hc1869a00} /* (28, 6, 20) {real, imag} */,
  {32'hc0407fb5, 32'hc1102567} /* (28, 6, 19) {real, imag} */,
  {32'h416736ee, 32'h408f7b27} /* (28, 6, 18) {real, imag} */,
  {32'hc1386818, 32'h3f2c9554} /* (28, 6, 17) {real, imag} */,
  {32'hc1810c44, 32'hc0e6bcfd} /* (28, 6, 16) {real, imag} */,
  {32'hc1546d57, 32'hc1409fcc} /* (28, 6, 15) {real, imag} */,
  {32'hc18ebda0, 32'hc1acf746} /* (28, 6, 14) {real, imag} */,
  {32'hc1911cca, 32'hc1b4e106} /* (28, 6, 13) {real, imag} */,
  {32'hc16e943d, 32'hc15320cb} /* (28, 6, 12) {real, imag} */,
  {32'hc03fc0e5, 32'hbf251830} /* (28, 6, 11) {real, imag} */,
  {32'hc189f768, 32'hc0cb4c49} /* (28, 6, 10) {real, imag} */,
  {32'hc07c38e7, 32'hc12aad12} /* (28, 6, 9) {real, imag} */,
  {32'h40915f5d, 32'hc1857bfe} /* (28, 6, 8) {real, imag} */,
  {32'h40f7d80c, 32'hc02017bc} /* (28, 6, 7) {real, imag} */,
  {32'h40728e68, 32'h417fd49a} /* (28, 6, 6) {real, imag} */,
  {32'hc1355900, 32'h415453a1} /* (28, 6, 5) {real, imag} */,
  {32'hc08ce92d, 32'h4007516e} /* (28, 6, 4) {real, imag} */,
  {32'hc0dbe23a, 32'hc0c94d9c} /* (28, 6, 3) {real, imag} */,
  {32'hc13588fb, 32'hc0607074} /* (28, 6, 2) {real, imag} */,
  {32'h40874828, 32'h4193a0b2} /* (28, 6, 1) {real, imag} */,
  {32'h41345bcc, 32'h41aab954} /* (28, 6, 0) {real, imag} */,
  {32'h413a5aad, 32'h41aa379e} /* (28, 5, 31) {real, imag} */,
  {32'h3f235eb0, 32'h419a1ca0} /* (28, 5, 30) {real, imag} */,
  {32'h414fde62, 32'h41d28a42} /* (28, 5, 29) {real, imag} */,
  {32'h4109d881, 32'h422206ef} /* (28, 5, 28) {real, imag} */,
  {32'hc0a01ebe, 32'h4232fa47} /* (28, 5, 27) {real, imag} */,
  {32'hc09cce3a, 32'h4216bb4d} /* (28, 5, 26) {real, imag} */,
  {32'h3fbeda48, 32'h41d22a5e} /* (28, 5, 25) {real, imag} */,
  {32'h409ec3a6, 32'h423196b9} /* (28, 5, 24) {real, imag} */,
  {32'h4075abff, 32'h4201d1aa} /* (28, 5, 23) {real, imag} */,
  {32'hbf320dc8, 32'h4201d9a6} /* (28, 5, 22) {real, imag} */,
  {32'hc0a2ef62, 32'h41a5bdab} /* (28, 5, 21) {real, imag} */,
  {32'hbfa9f502, 32'h4104f40a} /* (28, 5, 20) {real, imag} */,
  {32'hc1a39f87, 32'h3f3e3938} /* (28, 5, 19) {real, imag} */,
  {32'hc1bdbb6b, 32'hc17c6b64} /* (28, 5, 18) {real, imag} */,
  {32'h3fa3a460, 32'hc1b1efef} /* (28, 5, 17) {real, imag} */,
  {32'h40bd0554, 32'hc19e92b1} /* (28, 5, 16) {real, imag} */,
  {32'hc185d44e, 32'hc1cc6bf8} /* (28, 5, 15) {real, imag} */,
  {32'hc1570f3e, 32'hc1e2ac0c} /* (28, 5, 14) {real, imag} */,
  {32'h4085ebc2, 32'hc20fb5ad} /* (28, 5, 13) {real, imag} */,
  {32'h415d053e, 32'hc209965a} /* (28, 5, 12) {real, imag} */,
  {32'h405881c0, 32'hc1f40ba0} /* (28, 5, 11) {real, imag} */,
  {32'hc19e3360, 32'hc181e10e} /* (28, 5, 10) {real, imag} */,
  {32'hc2154351, 32'h3f42a2fc} /* (28, 5, 9) {real, imag} */,
  {32'hc1a99657, 32'h411bd661} /* (28, 5, 8) {real, imag} */,
  {32'h403b5258, 32'h4180f149} /* (28, 5, 7) {real, imag} */,
  {32'h4111f78b, 32'h40b5a6ae} /* (28, 5, 6) {real, imag} */,
  {32'h412a69e1, 32'h4189df8c} /* (28, 5, 5) {real, imag} */,
  {32'h3f8a1564, 32'h41950eb7} /* (28, 5, 4) {real, imag} */,
  {32'hc016f87a, 32'h4181cf68} /* (28, 5, 3) {real, imag} */,
  {32'h41986171, 32'h41cd9b60} /* (28, 5, 2) {real, imag} */,
  {32'h4114b670, 32'h41be5296} /* (28, 5, 1) {real, imag} */,
  {32'hbf7aa040, 32'h41bdf476} /* (28, 5, 0) {real, imag} */,
  {32'hc0753844, 32'hc1499e1d} /* (28, 4, 31) {real, imag} */,
  {32'h41141ae6, 32'hc0625b50} /* (28, 4, 30) {real, imag} */,
  {32'h41cc533f, 32'h3fba98a0} /* (28, 4, 29) {real, imag} */,
  {32'h419838bc, 32'hc1cf3793} /* (28, 4, 28) {real, imag} */,
  {32'h41120195, 32'hc10e01ef} /* (28, 4, 27) {real, imag} */,
  {32'hc0c96614, 32'hc1a44762} /* (28, 4, 26) {real, imag} */,
  {32'hc0e5d968, 32'hc206fad4} /* (28, 4, 25) {real, imag} */,
  {32'h3fdde3f0, 32'hc1b6aac0} /* (28, 4, 24) {real, imag} */,
  {32'h41527026, 32'hc205b2a2} /* (28, 4, 23) {real, imag} */,
  {32'h409d901c, 32'hc1f67d4e} /* (28, 4, 22) {real, imag} */,
  {32'h409d38de, 32'hc1d76ba5} /* (28, 4, 21) {real, imag} */,
  {32'hc12e5216, 32'h41b23ae0} /* (28, 4, 20) {real, imag} */,
  {32'hc1576f74, 32'h41b7ad12} /* (28, 4, 19) {real, imag} */,
  {32'hc1da35b2, 32'h41cba5b6} /* (28, 4, 18) {real, imag} */,
  {32'hc201b3e8, 32'h41854982} /* (28, 4, 17) {real, imag} */,
  {32'h409d5a7e, 32'h410bcb11} /* (28, 4, 16) {real, imag} */,
  {32'h402db654, 32'h419c5093} /* (28, 4, 15) {real, imag} */,
  {32'hc0c6246a, 32'h41d48ea4} /* (28, 4, 14) {real, imag} */,
  {32'hc0a29292, 32'h41d26c43} /* (28, 4, 13) {real, imag} */,
  {32'hc0d7884f, 32'h41989431} /* (28, 4, 12) {real, imag} */,
  {32'h4082f996, 32'h41376ab1} /* (28, 4, 11) {real, imag} */,
  {32'h418b1a9a, 32'hc11931f3} /* (28, 4, 10) {real, imag} */,
  {32'h421a8a00, 32'hc204a2ee} /* (28, 4, 9) {real, imag} */,
  {32'h41eb9cf4, 32'hc218d838} /* (28, 4, 8) {real, imag} */,
  {32'h41e3094a, 32'hc1b6d3d8} /* (28, 4, 7) {real, imag} */,
  {32'h41d8b212, 32'hc1992be9} /* (28, 4, 6) {real, imag} */,
  {32'hbffbe490, 32'hc1c95dca} /* (28, 4, 5) {real, imag} */,
  {32'h410fba5f, 32'hc140d4d9} /* (28, 4, 4) {real, imag} */,
  {32'hc0ea11b3, 32'hc1f6e046} /* (28, 4, 3) {real, imag} */,
  {32'hc1436cb2, 32'hc245ce7a} /* (28, 4, 2) {real, imag} */,
  {32'hc127a924, 32'hc2005302} /* (28, 4, 1) {real, imag} */,
  {32'h3fae8078, 32'hc196a48f} /* (28, 4, 0) {real, imag} */,
  {32'hbfe03c9c, 32'hc0df2b98} /* (28, 3, 31) {real, imag} */,
  {32'h41d086ef, 32'hbd188f40} /* (28, 3, 30) {real, imag} */,
  {32'h41a63789, 32'h413b367d} /* (28, 3, 29) {real, imag} */,
  {32'hbf80d920, 32'hc0ba4516} /* (28, 3, 28) {real, imag} */,
  {32'hc1235f3d, 32'hc1725920} /* (28, 3, 27) {real, imag} */,
  {32'h40918d62, 32'h3f916c04} /* (28, 3, 26) {real, imag} */,
  {32'h41503631, 32'h4114a9f2} /* (28, 3, 25) {real, imag} */,
  {32'hbef35280, 32'hc0e1b5b1} /* (28, 3, 24) {real, imag} */,
  {32'hc115ae64, 32'hc0daeff2} /* (28, 3, 23) {real, imag} */,
  {32'hc11c185c, 32'h417548d1} /* (28, 3, 22) {real, imag} */,
  {32'h41069c07, 32'h41b3acbe} /* (28, 3, 21) {real, imag} */,
  {32'hc195997a, 32'hc0559bd0} /* (28, 3, 20) {real, imag} */,
  {32'hc23e6406, 32'h40f324f8} /* (28, 3, 19) {real, imag} */,
  {32'hc2644828, 32'h4196eab8} /* (28, 3, 18) {real, imag} */,
  {32'hc2348195, 32'h4207f0b3} /* (28, 3, 17) {real, imag} */,
  {32'hc244da40, 32'h420cf1db} /* (28, 3, 16) {real, imag} */,
  {32'hc1a18412, 32'h4168a521} /* (28, 3, 15) {real, imag} */,
  {32'hbfcd96b8, 32'h3f52d9b8} /* (28, 3, 14) {real, imag} */,
  {32'h41b984e2, 32'hc0abe1f4} /* (28, 3, 13) {real, imag} */,
  {32'h4204db8c, 32'hc016300c} /* (28, 3, 12) {real, imag} */,
  {32'h419c3a82, 32'hc1361fd2} /* (28, 3, 11) {real, imag} */,
  {32'h41c5c900, 32'hc1a7fb4e} /* (28, 3, 10) {real, imag} */,
  {32'h42229cde, 32'hc1a3a9f1} /* (28, 3, 9) {real, imag} */,
  {32'h4210ccdc, 32'hc19b31f8} /* (28, 3, 8) {real, imag} */,
  {32'h4214f64d, 32'hc1682778} /* (28, 3, 7) {real, imag} */,
  {32'h422ae55b, 32'h40761988} /* (28, 3, 6) {real, imag} */,
  {32'h41dd40bb, 32'hbf3ee620} /* (28, 3, 5) {real, imag} */,
  {32'h4117679d, 32'h3fcbdb18} /* (28, 3, 4) {real, imag} */,
  {32'h420f6e76, 32'hc1a645ee} /* (28, 3, 3) {real, imag} */,
  {32'h42474084, 32'hc1b98073} /* (28, 3, 2) {real, imag} */,
  {32'h414ee089, 32'hc170b8ae} /* (28, 3, 1) {real, imag} */,
  {32'hc0d546b0, 32'hc0984e1e} /* (28, 3, 0) {real, imag} */,
  {32'hbe317dc0, 32'h4235f564} /* (28, 2, 31) {real, imag} */,
  {32'hc05ea4a0, 32'h4257d019} /* (28, 2, 30) {real, imag} */,
  {32'hbef35b00, 32'h420f50c0} /* (28, 2, 29) {real, imag} */,
  {32'hc0bf7bbc, 32'h425b4092} /* (28, 2, 28) {real, imag} */,
  {32'h40a2cfea, 32'h4243f0ca} /* (28, 2, 27) {real, imag} */,
  {32'h41da39ab, 32'h424825fa} /* (28, 2, 26) {real, imag} */,
  {32'h41b6ab70, 32'h4257b33c} /* (28, 2, 25) {real, imag} */,
  {32'hbf090330, 32'h4283105e} /* (28, 2, 24) {real, imag} */,
  {32'h3fdac010, 32'h42505686} /* (28, 2, 23) {real, imag} */,
  {32'h410772f6, 32'h425d6064} /* (28, 2, 22) {real, imag} */,
  {32'hc1139d4a, 32'h41550012} /* (28, 2, 21) {real, imag} */,
  {32'hc25d9d18, 32'hc25a48e1} /* (28, 2, 20) {real, imag} */,
  {32'hc24cf599, 32'hc2541169} /* (28, 2, 19) {real, imag} */,
  {32'hc27d0df3, 32'hc1ed1c22} /* (28, 2, 18) {real, imag} */,
  {32'hc21b2926, 32'hc23bdaa8} /* (28, 2, 17) {real, imag} */,
  {32'hc16d06fd, 32'hc27092b3} /* (28, 2, 16) {real, imag} */,
  {32'h41b5e540, 32'hc2732d4c} /* (28, 2, 15) {real, imag} */,
  {32'h404519de, 32'hc275efb5} /* (28, 2, 14) {real, imag} */,
  {32'hc0c03716, 32'hc26dc640} /* (28, 2, 13) {real, imag} */,
  {32'hc019aec8, 32'hc24d21c2} /* (28, 2, 12) {real, imag} */,
  {32'h4094c155, 32'hc1dd6104} /* (28, 2, 11) {real, imag} */,
  {32'h4216e8e2, 32'h421dc35c} /* (28, 2, 10) {real, imag} */,
  {32'h421c08fa, 32'h42634a12} /* (28, 2, 9) {real, imag} */,
  {32'h42475486, 32'h427a66f2} /* (28, 2, 8) {real, imag} */,
  {32'h425c476b, 32'h42913eda} /* (28, 2, 7) {real, imag} */,
  {32'h41b64dc4, 32'h426f7957} /* (28, 2, 6) {real, imag} */,
  {32'hc028691c, 32'h426dfbad} /* (28, 2, 5) {real, imag} */,
  {32'hc133f7dd, 32'h424e83d8} /* (28, 2, 4) {real, imag} */,
  {32'h40433cb0, 32'h42170cb4} /* (28, 2, 3) {real, imag} */,
  {32'h40c50eae, 32'h42651907} /* (28, 2, 2) {real, imag} */,
  {32'h41b5891d, 32'h426aaed7} /* (28, 2, 1) {real, imag} */,
  {32'h418dd878, 32'h42264952} /* (28, 2, 0) {real, imag} */,
  {32'hc19c2492, 32'hc232caaf} /* (28, 1, 31) {real, imag} */,
  {32'hc1f1b4bc, 32'hc2a05302} /* (28, 1, 30) {real, imag} */,
  {32'hc1c800d2, 32'hc2c2c44f} /* (28, 1, 29) {real, imag} */,
  {32'hc17a193d, 32'hc299d1cc} /* (28, 1, 28) {real, imag} */,
  {32'hc167082e, 32'hc28e606f} /* (28, 1, 27) {real, imag} */,
  {32'hc0e7b85c, 32'hc29b7ff4} /* (28, 1, 26) {real, imag} */,
  {32'hc1040c85, 32'hc299e9bf} /* (28, 1, 25) {real, imag} */,
  {32'hc1c964ee, 32'hc2a4994e} /* (28, 1, 24) {real, imag} */,
  {32'hc1e7a2c2, 32'hc2842eac} /* (28, 1, 23) {real, imag} */,
  {32'hc1df2394, 32'hc28e9288} /* (28, 1, 22) {real, imag} */,
  {32'hc19e1bbc, 32'hc2309d3e} /* (28, 1, 21) {real, imag} */,
  {32'hc197aa90, 32'h42489ada} /* (28, 1, 20) {real, imag} */,
  {32'hc08d26bc, 32'h42816045} /* (28, 1, 19) {real, imag} */,
  {32'hc12f98f1, 32'h427b9e90} /* (28, 1, 18) {real, imag} */,
  {32'hc1e77553, 32'h4298de25} /* (28, 1, 17) {real, imag} */,
  {32'hc21e9497, 32'h42956209} /* (28, 1, 16) {real, imag} */,
  {32'h40e46c33, 32'h429a63ca} /* (28, 1, 15) {real, imag} */,
  {32'h415a08e2, 32'h42a18420} /* (28, 1, 14) {real, imag} */,
  {32'hc0810af8, 32'h42875c8a} /* (28, 1, 13) {real, imag} */,
  {32'h41cde3f7, 32'h42a61997} /* (28, 1, 12) {real, imag} */,
  {32'h41f010d8, 32'h429a9cab} /* (28, 1, 11) {real, imag} */,
  {32'h41ad29e2, 32'hc0f9ffdc} /* (28, 1, 10) {real, imag} */,
  {32'h41a62b5a, 32'hc267f40e} /* (28, 1, 9) {real, imag} */,
  {32'h4206efcd, 32'hc28262ba} /* (28, 1, 8) {real, imag} */,
  {32'h4138ce8a, 32'hc2717593} /* (28, 1, 7) {real, imag} */,
  {32'h402049a8, 32'hc2883f3c} /* (28, 1, 6) {real, imag} */,
  {32'hc0447d90, 32'hc26eade7} /* (28, 1, 5) {real, imag} */,
  {32'hc22fe324, 32'hc2975b50} /* (28, 1, 4) {real, imag} */,
  {32'hc2149f7d, 32'hc2c88606} /* (28, 1, 3) {real, imag} */,
  {32'hc21e9faa, 32'hc28c9cb8} /* (28, 1, 2) {real, imag} */,
  {32'hc12b4b11, 32'hc282919b} /* (28, 1, 1) {real, imag} */,
  {32'hc1805f94, 32'hc2311bdc} /* (28, 1, 0) {real, imag} */,
  {32'hc181d893, 32'hc24731af} /* (28, 0, 31) {real, imag} */,
  {32'hc21670eb, 32'hc29205ae} /* (28, 0, 30) {real, imag} */,
  {32'hc20ca236, 32'hc2341168} /* (28, 0, 29) {real, imag} */,
  {32'hc1bffea8, 32'hc23001bb} /* (28, 0, 28) {real, imag} */,
  {32'hc2066d12, 32'hc210303c} /* (28, 0, 27) {real, imag} */,
  {32'hc1ee0634, 32'hc2714826} /* (28, 0, 26) {real, imag} */,
  {32'hc1caae00, 32'hc24711c8} /* (28, 0, 25) {real, imag} */,
  {32'hc03aa95f, 32'hc225dc5a} /* (28, 0, 24) {real, imag} */,
  {32'hc035bc3e, 32'hc22118d5} /* (28, 0, 23) {real, imag} */,
  {32'hc190369f, 32'hc25dfbb9} /* (28, 0, 22) {real, imag} */,
  {32'hc189583c, 32'hc213c061} /* (28, 0, 21) {real, imag} */,
  {32'h40ec5eae, 32'h411f63a0} /* (28, 0, 20) {real, imag} */,
  {32'hc192b0ba, 32'hc13c1606} /* (28, 0, 19) {real, imag} */,
  {32'hc1a49a5a, 32'hc177aa72} /* (28, 0, 18) {real, imag} */,
  {32'hc08a4a61, 32'h3e5dfda0} /* (28, 0, 17) {real, imag} */,
  {32'h3f8a2d04, 32'h414dd744} /* (28, 0, 16) {real, imag} */,
  {32'h40880725, 32'h4202d910} /* (28, 0, 15) {real, imag} */,
  {32'h41c57e97, 32'h424ff9c0} /* (28, 0, 14) {real, imag} */,
  {32'h4202f5be, 32'h4245839a} /* (28, 0, 13) {real, imag} */,
  {32'h416cf63f, 32'h42260779} /* (28, 0, 12) {real, imag} */,
  {32'h41707bef, 32'h423f4df2} /* (28, 0, 11) {real, imag} */,
  {32'h40db79d8, 32'h4207bef9} /* (28, 0, 10) {real, imag} */,
  {32'hc191f85b, 32'h40e96646} /* (28, 0, 9) {real, imag} */,
  {32'hc153b788, 32'h400d5a54} /* (28, 0, 8) {real, imag} */,
  {32'hc0020614, 32'h41b12cf1} /* (28, 0, 7) {real, imag} */,
  {32'h4176f814, 32'h41aa7275} /* (28, 0, 6) {real, imag} */,
  {32'hc12c53a4, 32'hc2309369} /* (28, 0, 5) {real, imag} */,
  {32'hc1bdf2f8, 32'hc271ecd9} /* (28, 0, 4) {real, imag} */,
  {32'hc11ce23a, 32'hc25132f6} /* (28, 0, 3) {real, imag} */,
  {32'hc1ac4342, 32'hc2486bb0} /* (28, 0, 2) {real, imag} */,
  {32'hc19066ab, 32'hc2501f03} /* (28, 0, 1) {real, imag} */,
  {32'hc0cb50cc, 32'hc198b57a} /* (28, 0, 0) {real, imag} */,
  {32'h40df930c, 32'h4163d3a3} /* (27, 31, 31) {real, imag} */,
  {32'h4189082e, 32'h41d9042d} /* (27, 31, 30) {real, imag} */,
  {32'h41c3fbb6, 32'h41324fda} /* (27, 31, 29) {real, imag} */,
  {32'h41a8b04e, 32'h412e3c4c} /* (27, 31, 28) {real, imag} */,
  {32'h41fddc4d, 32'h417e9180} /* (27, 31, 27) {real, imag} */,
  {32'h422cea0e, 32'h42011e85} /* (27, 31, 26) {real, imag} */,
  {32'h421e8581, 32'h421aaa85} /* (27, 31, 25) {real, imag} */,
  {32'h41c4dc52, 32'h41ee8887} /* (27, 31, 24) {real, imag} */,
  {32'h41ff9afb, 32'h41f9b339} /* (27, 31, 23) {real, imag} */,
  {32'h41ac6653, 32'h41d0f086} /* (27, 31, 22) {real, imag} */,
  {32'h4070a612, 32'h4206c052} /* (27, 31, 21) {real, imag} */,
  {32'hc1c84adc, 32'h3f672bd8} /* (27, 31, 20) {real, imag} */,
  {32'hc2225c66, 32'h40362592} /* (27, 31, 19) {real, imag} */,
  {32'hc1df855e, 32'h40a3fc4e} /* (27, 31, 18) {real, imag} */,
  {32'hc1d240aa, 32'hc0c76aae} /* (27, 31, 17) {real, imag} */,
  {32'hc1270b4a, 32'hc121a4ed} /* (27, 31, 16) {real, imag} */,
  {32'hc1d9f06f, 32'hc15fec83} /* (27, 31, 15) {real, imag} */,
  {32'hc1d67161, 32'hc1e7ba20} /* (27, 31, 14) {real, imag} */,
  {32'hc14c5e15, 32'hc229442c} /* (27, 31, 13) {real, imag} */,
  {32'hc18db9ea, 32'hc18b1916} /* (27, 31, 12) {real, imag} */,
  {32'hc152f882, 32'hc19cfccc} /* (27, 31, 11) {real, imag} */,
  {32'h41a280f6, 32'hbeea2c80} /* (27, 31, 10) {real, imag} */,
  {32'h420eb02b, 32'hbec80340} /* (27, 31, 9) {real, imag} */,
  {32'h411c8f6f, 32'h409920e2} /* (27, 31, 8) {real, imag} */,
  {32'h4192bc75, 32'h4168f1c9} /* (27, 31, 7) {real, imag} */,
  {32'h3f8cf750, 32'h40c1bf28} /* (27, 31, 6) {real, imag} */,
  {32'h40b2e68e, 32'h41cb2c58} /* (27, 31, 5) {real, imag} */,
  {32'h412f4de0, 32'h421bf7a5} /* (27, 31, 4) {real, imag} */,
  {32'h41a0bc7f, 32'h4202645f} /* (27, 31, 3) {real, imag} */,
  {32'h41cf6378, 32'h41c30360} /* (27, 31, 2) {real, imag} */,
  {32'h41a2365c, 32'h41d45f29} /* (27, 31, 1) {real, imag} */,
  {32'h40b9758a, 32'h4188aac8} /* (27, 31, 0) {real, imag} */,
  {32'h3e5fbbe0, 32'hc169816a} /* (27, 30, 31) {real, imag} */,
  {32'hc0681f9b, 32'hc19f4347} /* (27, 30, 30) {real, imag} */,
  {32'hc1629d6e, 32'hc1105486} /* (27, 30, 29) {real, imag} */,
  {32'hc1c623ff, 32'hc18000cc} /* (27, 30, 28) {real, imag} */,
  {32'hc1b167b6, 32'hc1224fb2} /* (27, 30, 27) {real, imag} */,
  {32'h3ea47bb8, 32'h40a740b0} /* (27, 30, 26) {real, imag} */,
  {32'h40a07906, 32'hc1041f62} /* (27, 30, 25) {real, imag} */,
  {32'hc148a5af, 32'hc211a140} /* (27, 30, 24) {real, imag} */,
  {32'hc207f285, 32'hc2350611} /* (27, 30, 23) {real, imag} */,
  {32'hc23ea14d, 32'hc1d94b00} /* (27, 30, 22) {real, imag} */,
  {32'hc10a49a4, 32'hc1025db2} /* (27, 30, 21) {real, imag} */,
  {32'h40806b06, 32'h4181993b} /* (27, 30, 20) {real, imag} */,
  {32'h40951395, 32'h425175bc} /* (27, 30, 19) {real, imag} */,
  {32'h416aa445, 32'h428c5288} /* (27, 30, 18) {real, imag} */,
  {32'h41a07f2a, 32'h42711754} /* (27, 30, 17) {real, imag} */,
  {32'h3feefde0, 32'h42570ffa} /* (27, 30, 16) {real, imag} */,
  {32'h412ee58c, 32'h4222dc76} /* (27, 30, 15) {real, imag} */,
  {32'h40c06836, 32'h41a59bcc} /* (27, 30, 14) {real, imag} */,
  {32'h41f1a4c6, 32'h41df5c00} /* (27, 30, 13) {real, imag} */,
  {32'h41c825aa, 32'h41a8edcf} /* (27, 30, 12) {real, imag} */,
  {32'h40ea4f18, 32'h418fb29e} /* (27, 30, 11) {real, imag} */,
  {32'h40b1b388, 32'hc1e29658} /* (27, 30, 10) {real, imag} */,
  {32'h413b2758, 32'hc226f990} /* (27, 30, 9) {real, imag} */,
  {32'h40a1a728, 32'hc22e97c1} /* (27, 30, 8) {real, imag} */,
  {32'hbf9316c4, 32'hc1d462b0} /* (27, 30, 7) {real, imag} */,
  {32'h408b9fc8, 32'hc1d80412} /* (27, 30, 6) {real, imag} */,
  {32'h4126bfb9, 32'hc1db7409} /* (27, 30, 5) {real, imag} */,
  {32'h403ee341, 32'hc194b664} /* (27, 30, 4) {real, imag} */,
  {32'hc16690ef, 32'h40718fd6} /* (27, 30, 3) {real, imag} */,
  {32'hc1760d2d, 32'hbff98f04} /* (27, 30, 2) {real, imag} */,
  {32'hc1211b67, 32'hc0cd3e08} /* (27, 30, 1) {real, imag} */,
  {32'hbfa33eae, 32'hc0692764} /* (27, 30, 0) {real, imag} */,
  {32'hc0517df6, 32'h407f957c} /* (27, 29, 31) {real, imag} */,
  {32'hc07d3612, 32'h41366011} /* (27, 29, 30) {real, imag} */,
  {32'h411e6043, 32'h41c8507e} /* (27, 29, 29) {real, imag} */,
  {32'hc1163907, 32'hc01cffd2} /* (27, 29, 28) {real, imag} */,
  {32'hc0dba848, 32'h418b22f6} /* (27, 29, 27) {real, imag} */,
  {32'h4082ff4e, 32'h41919ca3} /* (27, 29, 26) {real, imag} */,
  {32'h41843e7f, 32'h4173198c} /* (27, 29, 25) {real, imag} */,
  {32'h40884593, 32'h4181af6c} /* (27, 29, 24) {real, imag} */,
  {32'hc122fb12, 32'h413d120f} /* (27, 29, 23) {real, imag} */,
  {32'hbee40e60, 32'h4139b466} /* (27, 29, 22) {real, imag} */,
  {32'hbf910f7c, 32'h408c69af} /* (27, 29, 21) {real, imag} */,
  {32'hc048df80, 32'h417db154} /* (27, 29, 20) {real, imag} */,
  {32'hc153391a, 32'h41a5b311} /* (27, 29, 19) {real, imag} */,
  {32'hc21201ff, 32'h4179ee39} /* (27, 29, 18) {real, imag} */,
  {32'hc22969f4, 32'hc03cd020} /* (27, 29, 17) {real, imag} */,
  {32'hc1db7651, 32'h40da0dca} /* (27, 29, 16) {real, imag} */,
  {32'hc02fd032, 32'hc088ae7c} /* (27, 29, 15) {real, imag} */,
  {32'h410280fd, 32'hc1d8fce7} /* (27, 29, 14) {real, imag} */,
  {32'h3f71945a, 32'hc18cc140} /* (27, 29, 13) {real, imag} */,
  {32'hc036bca8, 32'hc1a9b703} /* (27, 29, 12) {real, imag} */,
  {32'hc11074f1, 32'hc0ccf34a} /* (27, 29, 11) {real, imag} */,
  {32'hc05efe28, 32'hc1a0ade8} /* (27, 29, 10) {real, imag} */,
  {32'h412f6bca, 32'hc1caa346} /* (27, 29, 9) {real, imag} */,
  {32'h40945208, 32'hc1cec353} /* (27, 29, 8) {real, imag} */,
  {32'h408bc64a, 32'hc1ae207a} /* (27, 29, 7) {real, imag} */,
  {32'hbffaa410, 32'hc1663800} /* (27, 29, 6) {real, imag} */,
  {32'hc057aea5, 32'hc106afef} /* (27, 29, 5) {real, imag} */,
  {32'hc11ea0a9, 32'hc140e63e} /* (27, 29, 4) {real, imag} */,
  {32'hc05d0007, 32'hbf13f9b8} /* (27, 29, 3) {real, imag} */,
  {32'hc106a4c7, 32'hc14615be} /* (27, 29, 2) {real, imag} */,
  {32'h40b03dc6, 32'hc1c6f748} /* (27, 29, 1) {real, imag} */,
  {32'h414bd792, 32'hc14436f2} /* (27, 29, 0) {real, imag} */,
  {32'h40e7a966, 32'h406ee519} /* (27, 28, 31) {real, imag} */,
  {32'h41cb2724, 32'hc0f69caf} /* (27, 28, 30) {real, imag} */,
  {32'h41b17209, 32'h3fabb6f8} /* (27, 28, 29) {real, imag} */,
  {32'h40fc9328, 32'h416593e4} /* (27, 28, 28) {real, imag} */,
  {32'h41248584, 32'h410562e6} /* (27, 28, 27) {real, imag} */,
  {32'h41c07f3e, 32'h418d81f4} /* (27, 28, 26) {real, imag} */,
  {32'h41dbf6aa, 32'h40688b0e} /* (27, 28, 25) {real, imag} */,
  {32'h41eb6bdf, 32'hc11b4bcb} /* (27, 28, 24) {real, imag} */,
  {32'h41825b12, 32'hc105ae94} /* (27, 28, 23) {real, imag} */,
  {32'h40db5f36, 32'h408d5f6c} /* (27, 28, 22) {real, imag} */,
  {32'hc1425493, 32'h3ec99600} /* (27, 28, 21) {real, imag} */,
  {32'h40251654, 32'hc0224aa8} /* (27, 28, 20) {real, imag} */,
  {32'hbfd8c150, 32'h401f30e0} /* (27, 28, 19) {real, imag} */,
  {32'hc13c9552, 32'hbe3f7f40} /* (27, 28, 18) {real, imag} */,
  {32'hc1e711e6, 32'h41599c94} /* (27, 28, 17) {real, imag} */,
  {32'hc1bc208c, 32'h4180819a} /* (27, 28, 16) {real, imag} */,
  {32'h40e61aec, 32'h3f8833a0} /* (27, 28, 15) {real, imag} */,
  {32'h40c14dde, 32'hc06f1ea2} /* (27, 28, 14) {real, imag} */,
  {32'h40f1f1bd, 32'hc1312782} /* (27, 28, 13) {real, imag} */,
  {32'h3de6f440, 32'hbf7cfb48} /* (27, 28, 12) {real, imag} */,
  {32'h409b8aea, 32'h406629eb} /* (27, 28, 11) {real, imag} */,
  {32'h41bdd453, 32'h40e4725c} /* (27, 28, 10) {real, imag} */,
  {32'h41f57d38, 32'hc12e7a38} /* (27, 28, 9) {real, imag} */,
  {32'h41d504de, 32'hc0fbbd20} /* (27, 28, 8) {real, imag} */,
  {32'h4174ee60, 32'h41023c06} /* (27, 28, 7) {real, imag} */,
  {32'h41bc596b, 32'hbf9821a0} /* (27, 28, 6) {real, imag} */,
  {32'h41e0ec82, 32'hc1483193} /* (27, 28, 5) {real, imag} */,
  {32'h3ddb0de0, 32'hc1373116} /* (27, 28, 4) {real, imag} */,
  {32'hc12b3142, 32'hc0826fbc} /* (27, 28, 3) {real, imag} */,
  {32'hc14547b9, 32'h419237ba} /* (27, 28, 2) {real, imag} */,
  {32'hbf1bc2e0, 32'h41c333f5} /* (27, 28, 1) {real, imag} */,
  {32'hc0031804, 32'h40f5d84e} /* (27, 28, 0) {real, imag} */,
  {32'hc1601fa8, 32'hc1384704} /* (27, 27, 31) {real, imag} */,
  {32'hc20e72c2, 32'hc123789c} /* (27, 27, 30) {real, imag} */,
  {32'hc199d8ac, 32'hc1869ee3} /* (27, 27, 29) {real, imag} */,
  {32'hc082c2ec, 32'hc1e0a2b2} /* (27, 27, 28) {real, imag} */,
  {32'h4050688a, 32'hc1d4ec19} /* (27, 27, 27) {real, imag} */,
  {32'h403cb20c, 32'hc0a0143e} /* (27, 27, 26) {real, imag} */,
  {32'hc17ef3a3, 32'h40321c58} /* (27, 27, 25) {real, imag} */,
  {32'hc136960d, 32'h4087d646} /* (27, 27, 24) {real, imag} */,
  {32'h40988ea2, 32'hbfdc8cce} /* (27, 27, 23) {real, imag} */,
  {32'h40ad5b75, 32'hc11cacf0} /* (27, 27, 22) {real, imag} */,
  {32'hc10a4445, 32'hc00c485a} /* (27, 27, 21) {real, imag} */,
  {32'h4026b896, 32'h40942cf2} /* (27, 27, 20) {real, imag} */,
  {32'h40d57a88, 32'h3f482b90} /* (27, 27, 19) {real, imag} */,
  {32'h4005f84f, 32'hc05a3fd4} /* (27, 27, 18) {real, imag} */,
  {32'h3e944630, 32'h4100aae7} /* (27, 27, 17) {real, imag} */,
  {32'hc0eb0f55, 32'h411641e4} /* (27, 27, 16) {real, imag} */,
  {32'hc0ae9442, 32'h4044d3a4} /* (27, 27, 15) {real, imag} */,
  {32'hc108312e, 32'h40fd0464} /* (27, 27, 14) {real, imag} */,
  {32'hbefd8940, 32'h40c8e2e5} /* (27, 27, 13) {real, imag} */,
  {32'h404fb71b, 32'hbf0a0bc8} /* (27, 27, 12) {real, imag} */,
  {32'h40f80612, 32'hc0debc8f} /* (27, 27, 11) {real, imag} */,
  {32'hc0c42070, 32'hc18db976} /* (27, 27, 10) {real, imag} */,
  {32'hc0cf53ad, 32'hc0906aa8} /* (27, 27, 9) {real, imag} */,
  {32'hc104604e, 32'h415b01d6} /* (27, 27, 8) {real, imag} */,
  {32'hc19331df, 32'hc09913c2} /* (27, 27, 7) {real, imag} */,
  {32'hc1a22de0, 32'h40b09ee9} /* (27, 27, 6) {real, imag} */,
  {32'hc1826622, 32'h411ceff2} /* (27, 27, 5) {real, imag} */,
  {32'hc0c2276c, 32'h40daaa88} /* (27, 27, 4) {real, imag} */,
  {32'hc177dfa0, 32'hc0d94ad8} /* (27, 27, 3) {real, imag} */,
  {32'hc1aadf8c, 32'hc132c67d} /* (27, 27, 2) {real, imag} */,
  {32'hc12162e8, 32'hbf8bf43a} /* (27, 27, 1) {real, imag} */,
  {32'hc09f27dc, 32'hc13093ab} /* (27, 27, 0) {real, imag} */,
  {32'hc0bd95da, 32'h3ebbc438} /* (27, 26, 31) {real, imag} */,
  {32'hc1184339, 32'hc0e0b386} /* (27, 26, 30) {real, imag} */,
  {32'h4081069c, 32'hc08734ee} /* (27, 26, 29) {real, imag} */,
  {32'h3fc62e9a, 32'hc0f78596} /* (27, 26, 28) {real, imag} */,
  {32'hbfa4b5f0, 32'h3fc03800} /* (27, 26, 27) {real, imag} */,
  {32'hc0ab6f4e, 32'hc03191f0} /* (27, 26, 26) {real, imag} */,
  {32'hc1012930, 32'hc0bb119e} /* (27, 26, 25) {real, imag} */,
  {32'hc0f64d26, 32'hc1aeeda4} /* (27, 26, 24) {real, imag} */,
  {32'hc106ee9e, 32'hc112bc20} /* (27, 26, 23) {real, imag} */,
  {32'hc11cf703, 32'h40629e1d} /* (27, 26, 22) {real, imag} */,
  {32'hc04da3f8, 32'h4102a206} /* (27, 26, 21) {real, imag} */,
  {32'hc04f040c, 32'h410dbef2} /* (27, 26, 20) {real, imag} */,
  {32'hc013bcc0, 32'h4087dc66} /* (27, 26, 19) {real, imag} */,
  {32'hc02ec22e, 32'hc0709eb6} /* (27, 26, 18) {real, imag} */,
  {32'h40681250, 32'hc09f91e4} /* (27, 26, 17) {real, imag} */,
  {32'h419a6e21, 32'hc0c35b33} /* (27, 26, 16) {real, imag} */,
  {32'h41130794, 32'h41a8f290} /* (27, 26, 15) {real, imag} */,
  {32'h3f29264e, 32'h40ab7acd} /* (27, 26, 14) {real, imag} */,
  {32'h41104666, 32'h4127af02} /* (27, 26, 13) {real, imag} */,
  {32'h41a6d914, 32'h414452a7} /* (27, 26, 12) {real, imag} */,
  {32'h41935ffc, 32'h415c9197} /* (27, 26, 11) {real, imag} */,
  {32'h4137c715, 32'h4106adcc} /* (27, 26, 10) {real, imag} */,
  {32'hc0f8f3f7, 32'h4185a552} /* (27, 26, 9) {real, imag} */,
  {32'hc048057c, 32'hc0bc17c4} /* (27, 26, 8) {real, imag} */,
  {32'hbf58d128, 32'hc043fc9a} /* (27, 26, 7) {real, imag} */,
  {32'h4017acc2, 32'h4044432c} /* (27, 26, 6) {real, imag} */,
  {32'hc16e7789, 32'hc0087070} /* (27, 26, 5) {real, imag} */,
  {32'h402a5768, 32'h3fe57594} /* (27, 26, 4) {real, imag} */,
  {32'h416585ce, 32'h40e3bf95} /* (27, 26, 3) {real, imag} */,
  {32'hc0e2f46a, 32'hbedd9a90} /* (27, 26, 2) {real, imag} */,
  {32'hbf06aa44, 32'hc0d076ba} /* (27, 26, 1) {real, imag} */,
  {32'h3f6d2b9b, 32'h408fc658} /* (27, 26, 0) {real, imag} */,
  {32'h411cf538, 32'hbf975774} /* (27, 25, 31) {real, imag} */,
  {32'h3f8ebe10, 32'h407e8a28} /* (27, 25, 30) {real, imag} */,
  {32'h3fc395c2, 32'h41c0f264} /* (27, 25, 29) {real, imag} */,
  {32'h40bd4a55, 32'h41a5309e} /* (27, 25, 28) {real, imag} */,
  {32'h409fd205, 32'hc003c3cb} /* (27, 25, 27) {real, imag} */,
  {32'h41175d76, 32'hc1006010} /* (27, 25, 26) {real, imag} */,
  {32'hc030cd71, 32'h40d47da7} /* (27, 25, 25) {real, imag} */,
  {32'hc0e63562, 32'h4133213c} /* (27, 25, 24) {real, imag} */,
  {32'hc0422891, 32'hc12c0a1c} /* (27, 25, 23) {real, imag} */,
  {32'h3fc9e780, 32'hc0a892a3} /* (27, 25, 22) {real, imag} */,
  {32'hc0f2a942, 32'h413a4d7a} /* (27, 25, 21) {real, imag} */,
  {32'h3f36cb70, 32'h41eb1e32} /* (27, 25, 20) {real, imag} */,
  {32'h409fd626, 32'h4142accd} /* (27, 25, 19) {real, imag} */,
  {32'hc1dce7ce, 32'hc14798e8} /* (27, 25, 18) {real, imag} */,
  {32'hc1bb5d2f, 32'hc16bd4c0} /* (27, 25, 17) {real, imag} */,
  {32'hc170c69c, 32'hc187c337} /* (27, 25, 16) {real, imag} */,
  {32'h3f6ff074, 32'hc17edf13} /* (27, 25, 15) {real, imag} */,
  {32'h3f9d1a64, 32'hc07f2222} /* (27, 25, 14) {real, imag} */,
  {32'hc18b62f3, 32'hc0bbdd5b} /* (27, 25, 13) {real, imag} */,
  {32'hc15fb25d, 32'hc121a6d0} /* (27, 25, 12) {real, imag} */,
  {32'h41342d4a, 32'hc179d6e7} /* (27, 25, 11) {real, imag} */,
  {32'hc01fc134, 32'hc0c62c24} /* (27, 25, 10) {real, imag} */,
  {32'hc0c1a7c7, 32'h409490b2} /* (27, 25, 9) {real, imag} */,
  {32'h40a92102, 32'hc10a6232} /* (27, 25, 8) {real, imag} */,
  {32'h40db2cce, 32'hc0de110e} /* (27, 25, 7) {real, imag} */,
  {32'hc04b6478, 32'h3ec48638} /* (27, 25, 6) {real, imag} */,
  {32'h410dea4b, 32'h3f22accc} /* (27, 25, 5) {real, imag} */,
  {32'h3fcc047c, 32'hc11f3277} /* (27, 25, 4) {real, imag} */,
  {32'hc0def91d, 32'hc118799e} /* (27, 25, 3) {real, imag} */,
  {32'hc1584d5e, 32'h419a0c5f} /* (27, 25, 2) {real, imag} */,
  {32'hbff39ad0, 32'h414617f2} /* (27, 25, 1) {real, imag} */,
  {32'h40f70198, 32'hc0883a4e} /* (27, 25, 0) {real, imag} */,
  {32'hc09f3baa, 32'hc1301560} /* (27, 24, 31) {real, imag} */,
  {32'hc10e49dc, 32'hc1906fa5} /* (27, 24, 30) {real, imag} */,
  {32'hc17b680d, 32'hc028678a} /* (27, 24, 29) {real, imag} */,
  {32'h3f23e5a8, 32'hc00284c3} /* (27, 24, 28) {real, imag} */,
  {32'hc03d381e, 32'hc0341f0a} /* (27, 24, 27) {real, imag} */,
  {32'hc179a22b, 32'hc16bf485} /* (27, 24, 26) {real, imag} */,
  {32'hc17e5722, 32'hc0a4952c} /* (27, 24, 25) {real, imag} */,
  {32'hbf292ff8, 32'h3d4d2a80} /* (27, 24, 24) {real, imag} */,
  {32'hc054001b, 32'hbf9bf9aa} /* (27, 24, 23) {real, imag} */,
  {32'hc1594144, 32'h400037dc} /* (27, 24, 22) {real, imag} */,
  {32'hc056487a, 32'h41516f95} /* (27, 24, 21) {real, imag} */,
  {32'h41297a00, 32'h416cf2f3} /* (27, 24, 20) {real, imag} */,
  {32'h409d070c, 32'hbec9adc0} /* (27, 24, 19) {real, imag} */,
  {32'h4020ed24, 32'h40ab68e4} /* (27, 24, 18) {real, imag} */,
  {32'hc11eb83a, 32'h40f8c327} /* (27, 24, 17) {real, imag} */,
  {32'hc1416f53, 32'hc09b94df} /* (27, 24, 16) {real, imag} */,
  {32'hbf75e838, 32'h40197252} /* (27, 24, 15) {real, imag} */,
  {32'h41404e80, 32'h4093bbaa} /* (27, 24, 14) {real, imag} */,
  {32'h4000b880, 32'hbfae1ce8} /* (27, 24, 13) {real, imag} */,
  {32'hbe30d850, 32'h40689975} /* (27, 24, 12) {real, imag} */,
  {32'h40aa7fd2, 32'h40ab365a} /* (27, 24, 11) {real, imag} */,
  {32'h3ea09740, 32'hc01b888c} /* (27, 24, 10) {real, imag} */,
  {32'h40634724, 32'h4109ce8c} /* (27, 24, 9) {real, imag} */,
  {32'h40bb5057, 32'hc037089a} /* (27, 24, 8) {real, imag} */,
  {32'hc0adabe4, 32'hc145c776} /* (27, 24, 7) {real, imag} */,
  {32'hc10ec20a, 32'h3f5c91e0} /* (27, 24, 6) {real, imag} */,
  {32'h3f997014, 32'hbf3a7630} /* (27, 24, 5) {real, imag} */,
  {32'h410965f2, 32'hbff544f0} /* (27, 24, 4) {real, imag} */,
  {32'h40d2667a, 32'hbe866950} /* (27, 24, 3) {real, imag} */,
  {32'hc13c5cdc, 32'h400b703e} /* (27, 24, 2) {real, imag} */,
  {32'hc15ee81e, 32'h40e27fba} /* (27, 24, 1) {real, imag} */,
  {32'hc0d1f165, 32'hc02d0990} /* (27, 24, 0) {real, imag} */,
  {32'hc05539b2, 32'h40e9bd96} /* (27, 23, 31) {real, imag} */,
  {32'h3fb04270, 32'h41418238} /* (27, 23, 30) {real, imag} */,
  {32'hc0c132ee, 32'hbfe66bb4} /* (27, 23, 29) {real, imag} */,
  {32'hc163158e, 32'hc156501c} /* (27, 23, 28) {real, imag} */,
  {32'hc0ef58d0, 32'hc137e2d7} /* (27, 23, 27) {real, imag} */,
  {32'h404d732e, 32'hc13106ee} /* (27, 23, 26) {real, imag} */,
  {32'h3eb12108, 32'hc1045832} /* (27, 23, 25) {real, imag} */,
  {32'h40a80240, 32'hc0c190a1} /* (27, 23, 24) {real, imag} */,
  {32'h40dab4fc, 32'hbf9ea998} /* (27, 23, 23) {real, imag} */,
  {32'h405ffc82, 32'hc11dee50} /* (27, 23, 22) {real, imag} */,
  {32'hc09c73a5, 32'hc0396516} /* (27, 23, 21) {real, imag} */,
  {32'h40212519, 32'hc0980316} /* (27, 23, 20) {real, imag} */,
  {32'hc1383334, 32'hc12ee8f8} /* (27, 23, 19) {real, imag} */,
  {32'hc07dff94, 32'h3fcfc2e8} /* (27, 23, 18) {real, imag} */,
  {32'hc16b9816, 32'h40ede3ed} /* (27, 23, 17) {real, imag} */,
  {32'hc113cac5, 32'h4107ff82} /* (27, 23, 16) {real, imag} */,
  {32'hc09a263a, 32'h40e04fca} /* (27, 23, 15) {real, imag} */,
  {32'h4031d56e, 32'h40ae042f} /* (27, 23, 14) {real, imag} */,
  {32'hc039dca6, 32'h4152d1d4} /* (27, 23, 13) {real, imag} */,
  {32'hc1422fd4, 32'h40b3c99d} /* (27, 23, 12) {real, imag} */,
  {32'hc18c9253, 32'h4120966d} /* (27, 23, 11) {real, imag} */,
  {32'hc0da9574, 32'h412e0386} /* (27, 23, 10) {real, imag} */,
  {32'h40ec48dc, 32'h40fcbc1a} /* (27, 23, 9) {real, imag} */,
  {32'h3f8d9d30, 32'h4094d290} /* (27, 23, 8) {real, imag} */,
  {32'hc080f432, 32'h40ddddf6} /* (27, 23, 7) {real, imag} */,
  {32'hc0ac34d2, 32'hc0d8aede} /* (27, 23, 6) {real, imag} */,
  {32'hc00a73e4, 32'hc07b5445} /* (27, 23, 5) {real, imag} */,
  {32'h40e46545, 32'h407a6aab} /* (27, 23, 4) {real, imag} */,
  {32'h4154fcb4, 32'hc0f7d697} /* (27, 23, 3) {real, imag} */,
  {32'hbfb2839c, 32'hc120f7d4} /* (27, 23, 2) {real, imag} */,
  {32'h400bfb38, 32'hc1291a6e} /* (27, 23, 1) {real, imag} */,
  {32'hbf123a32, 32'hc08846f2} /* (27, 23, 0) {real, imag} */,
  {32'h409616a9, 32'hc0163c4d} /* (27, 22, 31) {real, imag} */,
  {32'h4105670b, 32'hc004af28} /* (27, 22, 30) {real, imag} */,
  {32'h407c47b4, 32'h402646dd} /* (27, 22, 29) {real, imag} */,
  {32'h3ffc2362, 32'h40cfa45c} /* (27, 22, 28) {real, imag} */,
  {32'h409288ac, 32'hbfa03dc0} /* (27, 22, 27) {real, imag} */,
  {32'h40208cb0, 32'h403c2657} /* (27, 22, 26) {real, imag} */,
  {32'hbf7dcbd4, 32'hc03b2ce4} /* (27, 22, 25) {real, imag} */,
  {32'h40486f3f, 32'hbf9a3458} /* (27, 22, 24) {real, imag} */,
  {32'h412da256, 32'h411c8458} /* (27, 22, 23) {real, imag} */,
  {32'hc0f46ddc, 32'h40a76dc8} /* (27, 22, 22) {real, imag} */,
  {32'hc10b6b83, 32'hc05bf782} /* (27, 22, 21) {real, imag} */,
  {32'h3f4d7684, 32'h3ff5b7c6} /* (27, 22, 20) {real, imag} */,
  {32'h40bfd3fe, 32'hc05669fe} /* (27, 22, 19) {real, imag} */,
  {32'h413c750b, 32'hc0540edd} /* (27, 22, 18) {real, imag} */,
  {32'h40e8f38c, 32'hc1210bb3} /* (27, 22, 17) {real, imag} */,
  {32'h40ffbb34, 32'h3fea1ca4} /* (27, 22, 16) {real, imag} */,
  {32'h40d31554, 32'hc05b3b39} /* (27, 22, 15) {real, imag} */,
  {32'hbf866ec3, 32'hc10c760f} /* (27, 22, 14) {real, imag} */,
  {32'hc02ef146, 32'hc120308e} /* (27, 22, 13) {real, imag} */,
  {32'h412dcb8e, 32'hbf73da28} /* (27, 22, 12) {real, imag} */,
  {32'h40c59496, 32'h404eff2a} /* (27, 22, 11) {real, imag} */,
  {32'h402341a0, 32'h3f384538} /* (27, 22, 10) {real, imag} */,
  {32'h40ee1b1d, 32'hc163645f} /* (27, 22, 9) {real, imag} */,
  {32'h416ea35d, 32'hc14fe958} /* (27, 22, 8) {real, imag} */,
  {32'h40b962ef, 32'hc17c00c3} /* (27, 22, 7) {real, imag} */,
  {32'h3f4d9148, 32'hc12edc2d} /* (27, 22, 6) {real, imag} */,
  {32'h3e1d0670, 32'hc1446659} /* (27, 22, 5) {real, imag} */,
  {32'h409b87d9, 32'hc0c53821} /* (27, 22, 4) {real, imag} */,
  {32'hbf1815dc, 32'hbf1e5a0a} /* (27, 22, 3) {real, imag} */,
  {32'h40333a68, 32'hc04a1252} /* (27, 22, 2) {real, imag} */,
  {32'h411b5de2, 32'h3f6f2154} /* (27, 22, 1) {real, imag} */,
  {32'h40c6aa16, 32'h3f799e04} /* (27, 22, 0) {real, imag} */,
  {32'hc053eee8, 32'hc037221c} /* (27, 21, 31) {real, imag} */,
  {32'hc03fa768, 32'hc0848559} /* (27, 21, 30) {real, imag} */,
  {32'hc05bfddc, 32'hc0d5f9bd} /* (27, 21, 29) {real, imag} */,
  {32'hc10a90dc, 32'hc06f5a1f} /* (27, 21, 28) {real, imag} */,
  {32'hc0a3f493, 32'hc039041a} /* (27, 21, 27) {real, imag} */,
  {32'h3fbb4147, 32'hc04ab3bb} /* (27, 21, 26) {real, imag} */,
  {32'hc05613bc, 32'hc0ec7824} /* (27, 21, 25) {real, imag} */,
  {32'hc1203c30, 32'hc148f9ab} /* (27, 21, 24) {real, imag} */,
  {32'hc12087c7, 32'hc0e23a33} /* (27, 21, 23) {real, imag} */,
  {32'h3fa26cfc, 32'h400acc76} /* (27, 21, 22) {real, imag} */,
  {32'hc067d619, 32'h4052d2d3} /* (27, 21, 21) {real, imag} */,
  {32'h409d008a, 32'h40244a3f} /* (27, 21, 20) {real, imag} */,
  {32'h402905fc, 32'hc03cbcf4} /* (27, 21, 19) {real, imag} */,
  {32'h3b2b6800, 32'hc0e66294} /* (27, 21, 18) {real, imag} */,
  {32'hbffe336c, 32'hc118ace0} /* (27, 21, 17) {real, imag} */,
  {32'hc0c26858, 32'hc0ddd028} /* (27, 21, 16) {real, imag} */,
  {32'hc07a647f, 32'hc0282cd4} /* (27, 21, 15) {real, imag} */,
  {32'hc00ccbb6, 32'h3ef84b80} /* (27, 21, 14) {real, imag} */,
  {32'hc0c9bf74, 32'hc0732456} /* (27, 21, 13) {real, imag} */,
  {32'hc00a5fa1, 32'hc10024cc} /* (27, 21, 12) {real, imag} */,
  {32'h40b630d6, 32'h40bb3399} /* (27, 21, 11) {real, imag} */,
  {32'hc108a5e0, 32'h408b7d37} /* (27, 21, 10) {real, imag} */,
  {32'hc11aca98, 32'hbff7dbd4} /* (27, 21, 9) {real, imag} */,
  {32'h3fe153b4, 32'hc00873c2} /* (27, 21, 8) {real, imag} */,
  {32'h40636622, 32'h40a9c095} /* (27, 21, 7) {real, imag} */,
  {32'h405f0e1e, 32'h3f27bf68} /* (27, 21, 6) {real, imag} */,
  {32'h40f7bfdd, 32'h40311fa4} /* (27, 21, 5) {real, imag} */,
  {32'hc0201f0a, 32'h413ebe96} /* (27, 21, 4) {real, imag} */,
  {32'hc039f5c9, 32'h3fcbf558} /* (27, 21, 3) {real, imag} */,
  {32'h4030482b, 32'hc0a08bc4} /* (27, 21, 2) {real, imag} */,
  {32'hbf9dded0, 32'hc036a19b} /* (27, 21, 1) {real, imag} */,
  {32'h3e891180, 32'h4001bf48} /* (27, 21, 0) {real, imag} */,
  {32'hbeb30594, 32'h4029cd5e} /* (27, 20, 31) {real, imag} */,
  {32'hc01c9a98, 32'h40c5bf42} /* (27, 20, 30) {real, imag} */,
  {32'h406fad2c, 32'h40972b32} /* (27, 20, 29) {real, imag} */,
  {32'h417c3519, 32'hbfd603c4} /* (27, 20, 28) {real, imag} */,
  {32'h410d0c02, 32'h3fe3abae} /* (27, 20, 27) {real, imag} */,
  {32'h3dff0880, 32'h4084cd3d} /* (27, 20, 26) {real, imag} */,
  {32'h405ba088, 32'h40d73066} /* (27, 20, 25) {real, imag} */,
  {32'h3ff22eea, 32'h3fadfbce} /* (27, 20, 24) {real, imag} */,
  {32'hbeb63c58, 32'hc047047c} /* (27, 20, 23) {real, imag} */,
  {32'h3f1da2c0, 32'h40c1190a} /* (27, 20, 22) {real, imag} */,
  {32'hbf4f91c2, 32'h4092f518} /* (27, 20, 21) {real, imag} */,
  {32'h40a15dda, 32'h3e1c3980} /* (27, 20, 20) {real, imag} */,
  {32'h3f4f2900, 32'hc012eb40} /* (27, 20, 19) {real, imag} */,
  {32'h3f9f3fb0, 32'h40382a8e} /* (27, 20, 18) {real, imag} */,
  {32'hbfb2cc94, 32'h3ebc1910} /* (27, 20, 17) {real, imag} */,
  {32'hc09ecade, 32'hbea6a300} /* (27, 20, 16) {real, imag} */,
  {32'hc0351720, 32'hbe821c40} /* (27, 20, 15) {real, imag} */,
  {32'h40bc8c54, 32'hbe7ce740} /* (27, 20, 14) {real, imag} */,
  {32'h41219d79, 32'h3f91b5c0} /* (27, 20, 13) {real, imag} */,
  {32'hbe43f240, 32'h3f7c3fc8} /* (27, 20, 12) {real, imag} */,
  {32'h3fea5559, 32'hc095a1ee} /* (27, 20, 11) {real, imag} */,
  {32'hbf04aebe, 32'hc06412d0} /* (27, 20, 10) {real, imag} */,
  {32'h4083d993, 32'h3f4a1d80} /* (27, 20, 9) {real, imag} */,
  {32'h41291800, 32'h3fdf6224} /* (27, 20, 8) {real, imag} */,
  {32'h40ee5a1a, 32'h40015bf3} /* (27, 20, 7) {real, imag} */,
  {32'hbf42cac8, 32'h3f51ff98} /* (27, 20, 6) {real, imag} */,
  {32'hbfa6f500, 32'hc105ef31} /* (27, 20, 5) {real, imag} */,
  {32'hbfaaa90c, 32'hc0dd2b1c} /* (27, 20, 4) {real, imag} */,
  {32'hc03a2784, 32'h3faa2938} /* (27, 20, 3) {real, imag} */,
  {32'hbf98dc62, 32'h400bd9a7} /* (27, 20, 2) {real, imag} */,
  {32'hc0244059, 32'h409bbbf3} /* (27, 20, 1) {real, imag} */,
  {32'h3f856516, 32'h3fd20114} /* (27, 20, 0) {real, imag} */,
  {32'h3ff83731, 32'hbf0ffa5c} /* (27, 19, 31) {real, imag} */,
  {32'h3ecca4e8, 32'hc02a75ab} /* (27, 19, 30) {real, imag} */,
  {32'hc09ba781, 32'hc07d2bfc} /* (27, 19, 29) {real, imag} */,
  {32'hc0872e98, 32'h4014c168} /* (27, 19, 28) {real, imag} */,
  {32'hc0d26ece, 32'hbfed9950} /* (27, 19, 27) {real, imag} */,
  {32'hc06b1c54, 32'hc10d4016} /* (27, 19, 26) {real, imag} */,
  {32'hc0c22148, 32'h3f7fe3b0} /* (27, 19, 25) {real, imag} */,
  {32'h402e5d83, 32'h405035b0} /* (27, 19, 24) {real, imag} */,
  {32'h40d2c282, 32'h3e66d600} /* (27, 19, 23) {real, imag} */,
  {32'h402f24ad, 32'hc0c24def} /* (27, 19, 22) {real, imag} */,
  {32'h410692cc, 32'hc1230902} /* (27, 19, 21) {real, imag} */,
  {32'h40449fb2, 32'hc0919568} /* (27, 19, 20) {real, imag} */,
  {32'h3ef151c8, 32'hc069d206} /* (27, 19, 19) {real, imag} */,
  {32'hc04cfadc, 32'h400e11b5} /* (27, 19, 18) {real, imag} */,
  {32'h40041af6, 32'h403cb2e2} /* (27, 19, 17) {real, imag} */,
  {32'hc00754da, 32'hc0457eda} /* (27, 19, 16) {real, imag} */,
  {32'hc10ca380, 32'hc0f0aa2a} /* (27, 19, 15) {real, imag} */,
  {32'hc03dcb06, 32'h3f191910} /* (27, 19, 14) {real, imag} */,
  {32'h400a30b0, 32'h3f13aac6} /* (27, 19, 13) {real, imag} */,
  {32'hc08a2caa, 32'hbe5171c0} /* (27, 19, 12) {real, imag} */,
  {32'hc0d5eb75, 32'h3ffe4b28} /* (27, 19, 11) {real, imag} */,
  {32'h40278f4b, 32'hc078ef3a} /* (27, 19, 10) {real, imag} */,
  {32'hc011faea, 32'hc0c78e58} /* (27, 19, 9) {real, imag} */,
  {32'hc0703102, 32'h3e765678} /* (27, 19, 8) {real, imag} */,
  {32'hc0a94a3e, 32'h405770fc} /* (27, 19, 7) {real, imag} */,
  {32'hc0e7a254, 32'hbeea4140} /* (27, 19, 6) {real, imag} */,
  {32'hc04206c9, 32'h400860ab} /* (27, 19, 5) {real, imag} */,
  {32'h3e8ca8f8, 32'h3f80a7d1} /* (27, 19, 4) {real, imag} */,
  {32'hc000359f, 32'hc02ebe5a} /* (27, 19, 3) {real, imag} */,
  {32'hc0e909c6, 32'hc06520dd} /* (27, 19, 2) {real, imag} */,
  {32'hbcb01e00, 32'hc02a5bb2} /* (27, 19, 1) {real, imag} */,
  {32'h40617304, 32'hbec16c00} /* (27, 19, 0) {real, imag} */,
  {32'hbf0af864, 32'h3f90e294} /* (27, 18, 31) {real, imag} */,
  {32'h403a74ad, 32'h40aeda65} /* (27, 18, 30) {real, imag} */,
  {32'h3f4c23d5, 32'hbf97a9b8} /* (27, 18, 29) {real, imag} */,
  {32'hc006d94a, 32'hc05ace28} /* (27, 18, 28) {real, imag} */,
  {32'h3f4580f0, 32'h40351102} /* (27, 18, 27) {real, imag} */,
  {32'hbfc16636, 32'h3f52c480} /* (27, 18, 26) {real, imag} */,
  {32'hbf9734f7, 32'hc0832385} /* (27, 18, 25) {real, imag} */,
  {32'h3ec9a7a8, 32'h40191f7e} /* (27, 18, 24) {real, imag} */,
  {32'hbfc74372, 32'hbda47fe0} /* (27, 18, 23) {real, imag} */,
  {32'hbec76980, 32'hc0f8f7b2} /* (27, 18, 22) {real, imag} */,
  {32'h3fddaf04, 32'hc0a708a0} /* (27, 18, 21) {real, imag} */,
  {32'hbe70c4c0, 32'hc0e2d782} /* (27, 18, 20) {real, imag} */,
  {32'h403f6d0e, 32'h3da7c340} /* (27, 18, 19) {real, imag} */,
  {32'h40b33c36, 32'h401b0f1c} /* (27, 18, 18) {real, imag} */,
  {32'h40ccfe66, 32'hc0472b38} /* (27, 18, 17) {real, imag} */,
  {32'h40c5d5c2, 32'hbdc3b4c0} /* (27, 18, 16) {real, imag} */,
  {32'h402d797e, 32'h3fe9cef4} /* (27, 18, 15) {real, imag} */,
  {32'h3fc3af48, 32'hc0a303ad} /* (27, 18, 14) {real, imag} */,
  {32'h407ff45e, 32'hbf48a06e} /* (27, 18, 13) {real, imag} */,
  {32'h41013ce5, 32'h401bbefa} /* (27, 18, 12) {real, imag} */,
  {32'h40956be8, 32'h402972d5} /* (27, 18, 11) {real, imag} */,
  {32'h3f3e2058, 32'h3f02bf8c} /* (27, 18, 10) {real, imag} */,
  {32'hc07bfcc6, 32'h411c9ebc} /* (27, 18, 9) {real, imag} */,
  {32'hc03fe5dc, 32'h4032ae52} /* (27, 18, 8) {real, imag} */,
  {32'hc06677cf, 32'hc021091a} /* (27, 18, 7) {real, imag} */,
  {32'hc0c163c4, 32'hc0882c10} /* (27, 18, 6) {real, imag} */,
  {32'hc0814ca3, 32'hbf276504} /* (27, 18, 5) {real, imag} */,
  {32'h4088db4e, 32'hbfc8888c} /* (27, 18, 4) {real, imag} */,
  {32'h40ee4f14, 32'hbf8df928} /* (27, 18, 3) {real, imag} */,
  {32'h40047b59, 32'hc09d8eed} /* (27, 18, 2) {real, imag} */,
  {32'hc1082fdc, 32'hc12bcf02} /* (27, 18, 1) {real, imag} */,
  {32'hc0b2c9a6, 32'hc08511e4} /* (27, 18, 0) {real, imag} */,
  {32'hbec8eb80, 32'hbe816a46} /* (27, 17, 31) {real, imag} */,
  {32'h3f6c7870, 32'hc02077d8} /* (27, 17, 30) {real, imag} */,
  {32'h40ae12d4, 32'hc00d09ea} /* (27, 17, 29) {real, imag} */,
  {32'hc01b489b, 32'hc085b510} /* (27, 17, 28) {real, imag} */,
  {32'hbf811ff0, 32'hc049f8a0} /* (27, 17, 27) {real, imag} */,
  {32'h409c39ce, 32'hbfbe5773} /* (27, 17, 26) {real, imag} */,
  {32'h3e70ebc0, 32'h3f93e39b} /* (27, 17, 25) {real, imag} */,
  {32'hbe924368, 32'h3fc44bbe} /* (27, 17, 24) {real, imag} */,
  {32'h40fd7052, 32'h402e2886} /* (27, 17, 23) {real, imag} */,
  {32'h40fc79df, 32'h40713f24} /* (27, 17, 22) {real, imag} */,
  {32'h409876f3, 32'hbfbed2b2} /* (27, 17, 21) {real, imag} */,
  {32'h3fa1c736, 32'hc08a6784} /* (27, 17, 20) {real, imag} */,
  {32'h4043ea9c, 32'hc034254e} /* (27, 17, 19) {real, imag} */,
  {32'h401ca15c, 32'hc0684c9d} /* (27, 17, 18) {real, imag} */,
  {32'h40a0e69a, 32'hbfad7842} /* (27, 17, 17) {real, imag} */,
  {32'h3f223d54, 32'hc0973c56} /* (27, 17, 16) {real, imag} */,
  {32'hbf4d8120, 32'hc0862dfe} /* (27, 17, 15) {real, imag} */,
  {32'hbf45de88, 32'hc0c605d1} /* (27, 17, 14) {real, imag} */,
  {32'hbf169b9e, 32'hc0831163} /* (27, 17, 13) {real, imag} */,
  {32'hc0b9bfc0, 32'hc0020d18} /* (27, 17, 12) {real, imag} */,
  {32'hbfade3c4, 32'hc02fc91e} /* (27, 17, 11) {real, imag} */,
  {32'h40356e23, 32'hc0a2fd08} /* (27, 17, 10) {real, imag} */,
  {32'hbf764410, 32'hbecafcf0} /* (27, 17, 9) {real, imag} */,
  {32'hbf0730e4, 32'hc06780f6} /* (27, 17, 8) {real, imag} */,
  {32'h40cb0e10, 32'hc03f6824} /* (27, 17, 7) {real, imag} */,
  {32'h40dfdb47, 32'hc05377ac} /* (27, 17, 6) {real, imag} */,
  {32'h3fcaafc6, 32'hbfc51cb0} /* (27, 17, 5) {real, imag} */,
  {32'h407b23c0, 32'h3f106618} /* (27, 17, 4) {real, imag} */,
  {32'h408d58e9, 32'hc06ba48e} /* (27, 17, 3) {real, imag} */,
  {32'h40c0be88, 32'hc0c28dd6} /* (27, 17, 2) {real, imag} */,
  {32'h3f3a27fc, 32'hc0c4fb71} /* (27, 17, 1) {real, imag} */,
  {32'hbf96eb90, 32'hc0ca7b7e} /* (27, 17, 0) {real, imag} */,
  {32'hbf9d8448, 32'hbf04b880} /* (27, 16, 31) {real, imag} */,
  {32'hc0139934, 32'hbff06d30} /* (27, 16, 30) {real, imag} */,
  {32'h3f85d7d6, 32'h3f8b6330} /* (27, 16, 29) {real, imag} */,
  {32'h404de2c6, 32'hbfd05ed0} /* (27, 16, 28) {real, imag} */,
  {32'hbeaea800, 32'hc080606c} /* (27, 16, 27) {real, imag} */,
  {32'h3ee4d6a0, 32'h3fb5a2a0} /* (27, 16, 26) {real, imag} */,
  {32'h3fb10334, 32'hc0e3cf0a} /* (27, 16, 25) {real, imag} */,
  {32'hbfb9ab98, 32'hc01d38e0} /* (27, 16, 24) {real, imag} */,
  {32'hc012de15, 32'h40344c04} /* (27, 16, 23) {real, imag} */,
  {32'hbd4fd2c0, 32'h3fa66a18} /* (27, 16, 22) {real, imag} */,
  {32'h4065993a, 32'hbe77af00} /* (27, 16, 21) {real, imag} */,
  {32'h40856720, 32'h3fd00d2c} /* (27, 16, 20) {real, imag} */,
  {32'h4003e0a1, 32'h3ce50400} /* (27, 16, 19) {real, imag} */,
  {32'h4086beb2, 32'hbf3b1308} /* (27, 16, 18) {real, imag} */,
  {32'h40a56cdc, 32'h4041e060} /* (27, 16, 17) {real, imag} */,
  {32'hbff23698, 32'h3fdc8f14} /* (27, 16, 16) {real, imag} */,
  {32'hc071ba7a, 32'h3f16c930} /* (27, 16, 15) {real, imag} */,
  {32'hbf7ea600, 32'h400ae93c} /* (27, 16, 14) {real, imag} */,
  {32'h3ed11f80, 32'h4008b6bc} /* (27, 16, 13) {real, imag} */,
  {32'hc00e45f4, 32'h3fa1ad38} /* (27, 16, 12) {real, imag} */,
  {32'hbff5aae8, 32'hbfa970d8} /* (27, 16, 11) {real, imag} */,
  {32'h3fd12ee0, 32'h400f4025} /* (27, 16, 10) {real, imag} */,
  {32'h40e36954, 32'hbf90c9ea} /* (27, 16, 9) {real, imag} */,
  {32'h40037454, 32'hc02dc3d5} /* (27, 16, 8) {real, imag} */,
  {32'h3f8eac04, 32'h3faae67a} /* (27, 16, 7) {real, imag} */,
  {32'h3ea9fdc8, 32'h4005b044} /* (27, 16, 6) {real, imag} */,
  {32'hbf94fb90, 32'h3ede6080} /* (27, 16, 5) {real, imag} */,
  {32'h3f9f37a0, 32'hbd194400} /* (27, 16, 4) {real, imag} */,
  {32'hbf7cc1ce, 32'h3f821670} /* (27, 16, 3) {real, imag} */,
  {32'hc00c5a4c, 32'h4077deba} /* (27, 16, 2) {real, imag} */,
  {32'h3ed93120, 32'hc069be40} /* (27, 16, 1) {real, imag} */,
  {32'hbf78424e, 32'hc03527c8} /* (27, 16, 0) {real, imag} */,
  {32'hbeeb03e0, 32'hbfe2ba76} /* (27, 15, 31) {real, imag} */,
  {32'hbfd198a8, 32'h3ffd1c00} /* (27, 15, 30) {real, imag} */,
  {32'h3f7b2384, 32'h4049113a} /* (27, 15, 29) {real, imag} */,
  {32'h3f49d79c, 32'h3ffb9e00} /* (27, 15, 28) {real, imag} */,
  {32'h3fbfb1b0, 32'hbfea3240} /* (27, 15, 27) {real, imag} */,
  {32'h40a6086e, 32'hbd1f6da0} /* (27, 15, 26) {real, imag} */,
  {32'h40a6e17a, 32'hc019c9fe} /* (27, 15, 25) {real, imag} */,
  {32'h401f871d, 32'hbfa874fe} /* (27, 15, 24) {real, imag} */,
  {32'hc00d4804, 32'hbf0ecc98} /* (27, 15, 23) {real, imag} */,
  {32'hbfe5b9dc, 32'hc02a8204} /* (27, 15, 22) {real, imag} */,
  {32'hc01040ce, 32'hbf8f809e} /* (27, 15, 21) {real, imag} */,
  {32'h40b27510, 32'h3f00d672} /* (27, 15, 20) {real, imag} */,
  {32'h4098981e, 32'hc04aaa52} /* (27, 15, 19) {real, imag} */,
  {32'h3eed5320, 32'hc084b8ba} /* (27, 15, 18) {real, imag} */,
  {32'h3d4d0ec0, 32'hc01279d3} /* (27, 15, 17) {real, imag} */,
  {32'hbea7bd98, 32'hc057c3dc} /* (27, 15, 16) {real, imag} */,
  {32'hbe7f8d00, 32'h3fc64846} /* (27, 15, 15) {real, imag} */,
  {32'hbf9bf78c, 32'h40d78665} /* (27, 15, 14) {real, imag} */,
  {32'h3fd4e497, 32'h4080bfeb} /* (27, 15, 13) {real, imag} */,
  {32'h40f4d798, 32'hbf62eaa0} /* (27, 15, 12) {real, imag} */,
  {32'h403178ea, 32'hc0a7ded1} /* (27, 15, 11) {real, imag} */,
  {32'hc08990fe, 32'hc01a76f2} /* (27, 15, 10) {real, imag} */,
  {32'hc03e0da4, 32'h40387ee2} /* (27, 15, 9) {real, imag} */,
  {32'h3fee99ce, 32'h40b87529} /* (27, 15, 8) {real, imag} */,
  {32'hbf88bb26, 32'h3ef5af20} /* (27, 15, 7) {real, imag} */,
  {32'hbf9be39c, 32'h3eb8ac60} /* (27, 15, 6) {real, imag} */,
  {32'hc09ecb22, 32'hbf31e0a0} /* (27, 15, 5) {real, imag} */,
  {32'hc0a86a08, 32'h405e00b2} /* (27, 15, 4) {real, imag} */,
  {32'hc09cf359, 32'h4084c91b} /* (27, 15, 3) {real, imag} */,
  {32'hbde0f300, 32'h401a814c} /* (27, 15, 2) {real, imag} */,
  {32'hc0120f77, 32'h4086d109} /* (27, 15, 1) {real, imag} */,
  {32'hc04311d0, 32'hbdfc7f60} /* (27, 15, 0) {real, imag} */,
  {32'hbfbc5bc2, 32'hc03bbe8a} /* (27, 14, 31) {real, imag} */,
  {32'hc0841418, 32'hc040640a} /* (27, 14, 30) {real, imag} */,
  {32'hbfc0c056, 32'hc0dc17aa} /* (27, 14, 29) {real, imag} */,
  {32'hbe750620, 32'hc0f39df0} /* (27, 14, 28) {real, imag} */,
  {32'h3fc85ed8, 32'hbfc79b24} /* (27, 14, 27) {real, imag} */,
  {32'h4006cd35, 32'hc00d03e0} /* (27, 14, 26) {real, imag} */,
  {32'h3f07c7be, 32'hc009540e} /* (27, 14, 25) {real, imag} */,
  {32'hc03224a1, 32'h40aa8759} /* (27, 14, 24) {real, imag} */,
  {32'h40591509, 32'h4023f1bf} /* (27, 14, 23) {real, imag} */,
  {32'h40eea280, 32'h3fd57328} /* (27, 14, 22) {real, imag} */,
  {32'h40def359, 32'h4097c620} /* (27, 14, 21) {real, imag} */,
  {32'h40b5bfde, 32'h401f32e8} /* (27, 14, 20) {real, imag} */,
  {32'h4123d5e8, 32'hbd513a80} /* (27, 14, 19) {real, imag} */,
  {32'h40bea684, 32'hc087ba4e} /* (27, 14, 18) {real, imag} */,
  {32'h3fa2d428, 32'hc01da808} /* (27, 14, 17) {real, imag} */,
  {32'hbf7664f0, 32'h3e9cd330} /* (27, 14, 16) {real, imag} */,
  {32'hc023bca6, 32'hbee0bad0} /* (27, 14, 15) {real, imag} */,
  {32'hc149b77f, 32'h401a8392} /* (27, 14, 14) {real, imag} */,
  {32'hc0dbc33f, 32'hbf0752b2} /* (27, 14, 13) {real, imag} */,
  {32'h3d2ad500, 32'hc103936e} /* (27, 14, 12) {real, imag} */,
  {32'hc0204570, 32'h3f4c1dbc} /* (27, 14, 11) {real, imag} */,
  {32'hbf122cc8, 32'h40f8d8ce} /* (27, 14, 10) {real, imag} */,
  {32'hc032a85e, 32'h4056b1e2} /* (27, 14, 9) {real, imag} */,
  {32'hc079f3b4, 32'h3e8617f0} /* (27, 14, 8) {real, imag} */,
  {32'hbfff51fa, 32'hc010e5de} /* (27, 14, 7) {real, imag} */,
  {32'h40c8b622, 32'hbf669a02} /* (27, 14, 6) {real, imag} */,
  {32'hbfc2df44, 32'hbfeaa07e} /* (27, 14, 5) {real, imag} */,
  {32'hc0e1c266, 32'hc108d6b6} /* (27, 14, 4) {real, imag} */,
  {32'h402fa4b5, 32'hc0b1740c} /* (27, 14, 3) {real, imag} */,
  {32'h405c4b13, 32'hbd34dd80} /* (27, 14, 2) {real, imag} */,
  {32'hbeb8a890, 32'h40253766} /* (27, 14, 1) {real, imag} */,
  {32'h4031cdd9, 32'h404e78f0} /* (27, 14, 0) {real, imag} */,
  {32'h3f8b10c9, 32'hc008e2bd} /* (27, 13, 31) {real, imag} */,
  {32'hbfd75292, 32'hbf4ab0f4} /* (27, 13, 30) {real, imag} */,
  {32'h3e96d5f0, 32'h4095d00e} /* (27, 13, 29) {real, imag} */,
  {32'h3e595a00, 32'h403938f8} /* (27, 13, 28) {real, imag} */,
  {32'hbfd42042, 32'hbfba01d0} /* (27, 13, 27) {real, imag} */,
  {32'hbf4b7cb8, 32'h3f3edbb8} /* (27, 13, 26) {real, imag} */,
  {32'hc0dad8ce, 32'h3e90ede0} /* (27, 13, 25) {real, imag} */,
  {32'hc04738bd, 32'h3fede9c0} /* (27, 13, 24) {real, imag} */,
  {32'hbe78fbd0, 32'hbf5b4f70} /* (27, 13, 23) {real, imag} */,
  {32'h3f0d6e6c, 32'h405c3af2} /* (27, 13, 22) {real, imag} */,
  {32'hc0c5e9c2, 32'h40eb0a31} /* (27, 13, 21) {real, imag} */,
  {32'hc03d8296, 32'h409fc72e} /* (27, 13, 20) {real, imag} */,
  {32'hc0b618c4, 32'hbe89b5f0} /* (27, 13, 19) {real, imag} */,
  {32'h400a15c4, 32'hc07b2f25} /* (27, 13, 18) {real, imag} */,
  {32'h40e282bb, 32'hc1458468} /* (27, 13, 17) {real, imag} */,
  {32'h4008dd7e, 32'hc06f7814} /* (27, 13, 16) {real, imag} */,
  {32'hc0b108ff, 32'h40dcd4ba} /* (27, 13, 15) {real, imag} */,
  {32'hbf45033a, 32'h40b22a42} /* (27, 13, 14) {real, imag} */,
  {32'hbd0db1a0, 32'h3fadea93} /* (27, 13, 13) {real, imag} */,
  {32'hc103dd01, 32'hc035cd20} /* (27, 13, 12) {real, imag} */,
  {32'hc12da7e2, 32'hc103f41d} /* (27, 13, 11) {real, imag} */,
  {32'hc0040d6d, 32'hc0beba15} /* (27, 13, 10) {real, imag} */,
  {32'hbed64310, 32'h401caa78} /* (27, 13, 9) {real, imag} */,
  {32'hc000ea44, 32'h3f9e890f} /* (27, 13, 8) {real, imag} */,
  {32'h3fbcacb2, 32'h3e54f1c0} /* (27, 13, 7) {real, imag} */,
  {32'h3f7743f0, 32'h404670e8} /* (27, 13, 6) {real, imag} */,
  {32'h3e909408, 32'hbfeac2d6} /* (27, 13, 5) {real, imag} */,
  {32'h3fd17b1e, 32'hbf204ce2} /* (27, 13, 4) {real, imag} */,
  {32'h407bbeff, 32'hc0a0787d} /* (27, 13, 3) {real, imag} */,
  {32'h3e8b56c8, 32'hc031b9f1} /* (27, 13, 2) {real, imag} */,
  {32'hc0be81ae, 32'h40df391b} /* (27, 13, 1) {real, imag} */,
  {32'hc010ab34, 32'h40015970} /* (27, 13, 0) {real, imag} */,
  {32'h4088ab45, 32'h40b15f85} /* (27, 12, 31) {real, imag} */,
  {32'h40dc506c, 32'hbf252640} /* (27, 12, 30) {real, imag} */,
  {32'h4132269c, 32'hbf1fb110} /* (27, 12, 29) {real, imag} */,
  {32'h41142009, 32'h4027ea36} /* (27, 12, 28) {real, imag} */,
  {32'hbf9abdec, 32'h3f331814} /* (27, 12, 27) {real, imag} */,
  {32'hc0b69d8a, 32'h4116f1ae} /* (27, 12, 26) {real, imag} */,
  {32'hc0148d78, 32'h40ddf480} /* (27, 12, 25) {real, imag} */,
  {32'h40a04122, 32'hc07185ad} /* (27, 12, 24) {real, imag} */,
  {32'h3fabdeca, 32'hc11189f9} /* (27, 12, 23) {real, imag} */,
  {32'h4037c769, 32'hc13809c1} /* (27, 12, 22) {real, imag} */,
  {32'h403ee13c, 32'hc0c43e26} /* (27, 12, 21) {real, imag} */,
  {32'hbf159f10, 32'h409ff11c} /* (27, 12, 20) {real, imag} */,
  {32'hc0279578, 32'h40d33458} /* (27, 12, 19) {real, imag} */,
  {32'hc0821f08, 32'h40aae1f9} /* (27, 12, 18) {real, imag} */,
  {32'hc09a7927, 32'h40aa9b73} /* (27, 12, 17) {real, imag} */,
  {32'hbf013170, 32'hc11590c6} /* (27, 12, 16) {real, imag} */,
  {32'h404fca66, 32'hc0d8eaf8} /* (27, 12, 15) {real, imag} */,
  {32'h40947c96, 32'hbeb105a0} /* (27, 12, 14) {real, imag} */,
  {32'hbf898480, 32'hbf734640} /* (27, 12, 13) {real, imag} */,
  {32'hbfdf4608, 32'hc0e9e643} /* (27, 12, 12) {real, imag} */,
  {32'h4059aed2, 32'hc021138d} /* (27, 12, 11) {real, imag} */,
  {32'h40048518, 32'h40d35f68} /* (27, 12, 10) {real, imag} */,
  {32'h3fe411a4, 32'h40b3c140} /* (27, 12, 9) {real, imag} */,
  {32'hbef397b0, 32'hc036dea6} /* (27, 12, 8) {real, imag} */,
  {32'hc00e261b, 32'hbeab2368} /* (27, 12, 7) {real, imag} */,
  {32'h40b0e72f, 32'h3fe8fd44} /* (27, 12, 6) {real, imag} */,
  {32'h3ff88170, 32'h400c9b44} /* (27, 12, 5) {real, imag} */,
  {32'h4049df7e, 32'h40c4e0ca} /* (27, 12, 4) {real, imag} */,
  {32'h407435e2, 32'h41026dfc} /* (27, 12, 3) {real, imag} */,
  {32'hbff4a452, 32'hc00bf4f9} /* (27, 12, 2) {real, imag} */,
  {32'h3f971b62, 32'h3f92ac94} /* (27, 12, 1) {real, imag} */,
  {32'h3f9fc666, 32'h4112f990} /* (27, 12, 0) {real, imag} */,
  {32'hc01290f4, 32'hc0fe3b8a} /* (27, 11, 31) {real, imag} */,
  {32'h4099174c, 32'hc16342c4} /* (27, 11, 30) {real, imag} */,
  {32'h3fdee278, 32'hc1047d30} /* (27, 11, 29) {real, imag} */,
  {32'hc072cd9e, 32'hc0768f61} /* (27, 11, 28) {real, imag} */,
  {32'h40c7fbbf, 32'h3fdf6bd4} /* (27, 11, 27) {real, imag} */,
  {32'h4042b050, 32'h40351833} /* (27, 11, 26) {real, imag} */,
  {32'h3f108810, 32'h406c1084} /* (27, 11, 25) {real, imag} */,
  {32'hbd3cf100, 32'hbf49f710} /* (27, 11, 24) {real, imag} */,
  {32'h4113e1e1, 32'hc1193f92} /* (27, 11, 23) {real, imag} */,
  {32'h41445c9a, 32'hc15d0454} /* (27, 11, 22) {real, imag} */,
  {32'h4129eb4e, 32'hbee99ba0} /* (27, 11, 21) {real, imag} */,
  {32'hc00a93fe, 32'h3f20143c} /* (27, 11, 20) {real, imag} */,
  {32'hc13123ed, 32'h403c92e8} /* (27, 11, 19) {real, imag} */,
  {32'hbee47f60, 32'h3f89d670} /* (27, 11, 18) {real, imag} */,
  {32'hbe2b4b40, 32'hbfea777e} /* (27, 11, 17) {real, imag} */,
  {32'hbfbbb700, 32'hbf1f5a30} /* (27, 11, 16) {real, imag} */,
  {32'h404ff841, 32'hc0bd2f56} /* (27, 11, 15) {real, imag} */,
  {32'h3ff96a33, 32'hc1221152} /* (27, 11, 14) {real, imag} */,
  {32'hc0960448, 32'hbfbdad71} /* (27, 11, 13) {real, imag} */,
  {32'hc04c6a9f, 32'h40b83bf3} /* (27, 11, 12) {real, imag} */,
  {32'hc0cffd5a, 32'h41353a44} /* (27, 11, 11) {real, imag} */,
  {32'hc055981a, 32'hc087926d} /* (27, 11, 10) {real, imag} */,
  {32'h404363ce, 32'hbf26b868} /* (27, 11, 9) {real, imag} */,
  {32'h41020c58, 32'hc0737862} /* (27, 11, 8) {real, imag} */,
  {32'h403180ee, 32'h3f3e9e38} /* (27, 11, 7) {real, imag} */,
  {32'hc100db5c, 32'hc007cc06} /* (27, 11, 6) {real, imag} */,
  {32'hc0b580d5, 32'hc05a2254} /* (27, 11, 5) {real, imag} */,
  {32'h3ff92c4d, 32'hc03a47a0} /* (27, 11, 4) {real, imag} */,
  {32'hc0093dbf, 32'hc0bfe248} /* (27, 11, 3) {real, imag} */,
  {32'h3e587d50, 32'h401e14bb} /* (27, 11, 2) {real, imag} */,
  {32'h41036968, 32'hc0fedc82} /* (27, 11, 1) {real, imag} */,
  {32'h40073ebc, 32'hc139605e} /* (27, 11, 0) {real, imag} */,
  {32'hc08033ff, 32'h40c41e82} /* (27, 10, 31) {real, imag} */,
  {32'h4035d6a9, 32'h40fe5894} /* (27, 10, 30) {real, imag} */,
  {32'h400023f0, 32'h4119ac8b} /* (27, 10, 29) {real, imag} */,
  {32'hbf8664a6, 32'h3f4d587c} /* (27, 10, 28) {real, imag} */,
  {32'h404231c5, 32'hc0d9b1da} /* (27, 10, 27) {real, imag} */,
  {32'h3f702680, 32'hc04f033f} /* (27, 10, 26) {real, imag} */,
  {32'h406c78af, 32'h400046b8} /* (27, 10, 25) {real, imag} */,
  {32'hc0b0bbf0, 32'h4023d564} /* (27, 10, 24) {real, imag} */,
  {32'h3fa6d6e0, 32'hbefb5560} /* (27, 10, 23) {real, imag} */,
  {32'h3fd83250, 32'hc0256a1f} /* (27, 10, 22) {real, imag} */,
  {32'hc0708d44, 32'h3fb4abbc} /* (27, 10, 21) {real, imag} */,
  {32'hc0d58a10, 32'hc0e01a60} /* (27, 10, 20) {real, imag} */,
  {32'h406f2a04, 32'hc120da4e} /* (27, 10, 19) {real, imag} */,
  {32'h41200505, 32'hc0503ae1} /* (27, 10, 18) {real, imag} */,
  {32'hbe25c240, 32'hc15be671} /* (27, 10, 17) {real, imag} */,
  {32'hc143507a, 32'hc1178282} /* (27, 10, 16) {real, imag} */,
  {32'hc09f723e, 32'h3fdf73ea} /* (27, 10, 15) {real, imag} */,
  {32'hbfb4632b, 32'hbfa1f49e} /* (27, 10, 14) {real, imag} */,
  {32'h401f1672, 32'hbf974754} /* (27, 10, 13) {real, imag} */,
  {32'hc0963115, 32'h40c79e57} /* (27, 10, 12) {real, imag} */,
  {32'hc1bd76f8, 32'h4103039c} /* (27, 10, 11) {real, imag} */,
  {32'hc1360576, 32'h41812e8e} /* (27, 10, 10) {real, imag} */,
  {32'h40b23de7, 32'h41492b45} /* (27, 10, 9) {real, imag} */,
  {32'h40f913fe, 32'h413f9830} /* (27, 10, 8) {real, imag} */,
  {32'h40a1e8f5, 32'h410b3285} /* (27, 10, 7) {real, imag} */,
  {32'h411e8fc6, 32'h410ff623} /* (27, 10, 6) {real, imag} */,
  {32'h3fdcf36a, 32'h41205a33} /* (27, 10, 5) {real, imag} */,
  {32'h3f9fd6e4, 32'h404051e2} /* (27, 10, 4) {real, imag} */,
  {32'hc0e135e8, 32'h3fdf2cdd} /* (27, 10, 3) {real, imag} */,
  {32'hc15207d6, 32'h3ffa2b2c} /* (27, 10, 2) {real, imag} */,
  {32'hc10bd86a, 32'h3fdce8e6} /* (27, 10, 1) {real, imag} */,
  {32'hc06353bc, 32'h4061e481} /* (27, 10, 0) {real, imag} */,
  {32'h406fb5d6, 32'h3ff126f6} /* (27, 9, 31) {real, imag} */,
  {32'h3f844380, 32'h409fba70} /* (27, 9, 30) {real, imag} */,
  {32'hbfe36066, 32'h4138daee} /* (27, 9, 29) {real, imag} */,
  {32'hc0a12519, 32'h41536450} /* (27, 9, 28) {real, imag} */,
  {32'hc15480f0, 32'h4128c191} /* (27, 9, 27) {real, imag} */,
  {32'hc127ec08, 32'hc09f5cbc} /* (27, 9, 26) {real, imag} */,
  {32'h408b73f0, 32'hc150ea98} /* (27, 9, 25) {real, imag} */,
  {32'h3f867a42, 32'hc149187a} /* (27, 9, 24) {real, imag} */,
  {32'h40484a17, 32'hc10dc733} /* (27, 9, 23) {real, imag} */,
  {32'hbfff7a60, 32'hc10e4528} /* (27, 9, 22) {real, imag} */,
  {32'hc0b393e7, 32'hbf92c214} /* (27, 9, 21) {real, imag} */,
  {32'h40858204, 32'hc103e46f} /* (27, 9, 20) {real, imag} */,
  {32'h411ceb2e, 32'hbfbef6ac} /* (27, 9, 19) {real, imag} */,
  {32'hc0ed3452, 32'h413c0036} /* (27, 9, 18) {real, imag} */,
  {32'hc07d1668, 32'h408ff051} /* (27, 9, 17) {real, imag} */,
  {32'hc14baecf, 32'hc0d01bd5} /* (27, 9, 16) {real, imag} */,
  {32'hbf1a96e8, 32'h4047b343} /* (27, 9, 15) {real, imag} */,
  {32'h40ead64b, 32'h413dd98e} /* (27, 9, 14) {real, imag} */,
  {32'h4176053a, 32'h4107c55c} /* (27, 9, 13) {real, imag} */,
  {32'h404b1ac8, 32'h401e036e} /* (27, 9, 12) {real, imag} */,
  {32'h413da4de, 32'hc1536561} /* (27, 9, 11) {real, imag} */,
  {32'hc00d4890, 32'hc041862e} /* (27, 9, 10) {real, imag} */,
  {32'hc13c1712, 32'hc0f78226} /* (27, 9, 9) {real, imag} */,
  {32'hc157fe73, 32'h40de333e} /* (27, 9, 8) {real, imag} */,
  {32'h3e1e5df0, 32'h40f9d0fa} /* (27, 9, 7) {real, imag} */,
  {32'hbf27e0a0, 32'h3fbef568} /* (27, 9, 6) {real, imag} */,
  {32'h41727633, 32'hc11f34e1} /* (27, 9, 5) {real, imag} */,
  {32'h40afab11, 32'hbfcadda6} /* (27, 9, 4) {real, imag} */,
  {32'h3fb33824, 32'h4166a6be} /* (27, 9, 3) {real, imag} */,
  {32'hc015d8c2, 32'h40f96df8} /* (27, 9, 2) {real, imag} */,
  {32'hc10029c4, 32'hc08f8b40} /* (27, 9, 1) {real, imag} */,
  {32'hbff39917, 32'hbf708d40} /* (27, 9, 0) {real, imag} */,
  {32'hc0c3294e, 32'h41174ff6} /* (27, 8, 31) {real, imag} */,
  {32'h3fe6c554, 32'h40bc73fd} /* (27, 8, 30) {real, imag} */,
  {32'h41025b9b, 32'hc14add12} /* (27, 8, 29) {real, imag} */,
  {32'h40bcf251, 32'hc057dd71} /* (27, 8, 28) {real, imag} */,
  {32'h4132fa30, 32'hc0ff323d} /* (27, 8, 27) {real, imag} */,
  {32'h4105197f, 32'hc1d422aa} /* (27, 8, 26) {real, imag} */,
  {32'hbf7c0458, 32'hc1a0304c} /* (27, 8, 25) {real, imag} */,
  {32'hc03112a6, 32'h3f9b233c} /* (27, 8, 24) {real, imag} */,
  {32'h3fd72c8a, 32'hc05ddb1f} /* (27, 8, 23) {real, imag} */,
  {32'h3e258780, 32'hbecb2e40} /* (27, 8, 22) {real, imag} */,
  {32'h413bdeec, 32'hc014aa54} /* (27, 8, 21) {real, imag} */,
  {32'h418ec457, 32'h40c0799a} /* (27, 8, 20) {real, imag} */,
  {32'h40388777, 32'h41426616} /* (27, 8, 19) {real, imag} */,
  {32'h40b37344, 32'h4190615c} /* (27, 8, 18) {real, imag} */,
  {32'h41424f26, 32'h41843bd4} /* (27, 8, 17) {real, imag} */,
  {32'hc12a5d99, 32'h40c3645d} /* (27, 8, 16) {real, imag} */,
  {32'hc153b26c, 32'hbfc163d4} /* (27, 8, 15) {real, imag} */,
  {32'hc15eaa9c, 32'hc1801d4c} /* (27, 8, 14) {real, imag} */,
  {32'hc0b36b34, 32'hc13dfb03} /* (27, 8, 13) {real, imag} */,
  {32'h41001c6f, 32'h4104e3a5} /* (27, 8, 12) {real, imag} */,
  {32'h413ac2d5, 32'h4025cb93} /* (27, 8, 11) {real, imag} */,
  {32'hc14c83f2, 32'hc0e4db18} /* (27, 8, 10) {real, imag} */,
  {32'hc16ed099, 32'hbe4ac380} /* (27, 8, 9) {real, imag} */,
  {32'hc03682aa, 32'hc0d15e53} /* (27, 8, 8) {real, imag} */,
  {32'hc0a61792, 32'hbf14cae0} /* (27, 8, 7) {real, imag} */,
  {32'hc1130c3e, 32'hc0e1078a} /* (27, 8, 6) {real, imag} */,
  {32'hbfd1ed0c, 32'hc1af30aa} /* (27, 8, 5) {real, imag} */,
  {32'hc0a10438, 32'hc1566678} /* (27, 8, 4) {real, imag} */,
  {32'hc04d5c4c, 32'hc0388aee} /* (27, 8, 3) {real, imag} */,
  {32'hbf2a90e8, 32'hc15c6e1e} /* (27, 8, 2) {real, imag} */,
  {32'h41218876, 32'hc135dca3} /* (27, 8, 1) {real, imag} */,
  {32'h4098e437, 32'hc08fc849} /* (27, 8, 0) {real, imag} */,
  {32'h40fc9850, 32'hbc0fe000} /* (27, 7, 31) {real, imag} */,
  {32'h41556d78, 32'h40f61c34} /* (27, 7, 30) {real, imag} */,
  {32'h40ed2f30, 32'hc085ad90} /* (27, 7, 29) {real, imag} */,
  {32'hc0c82619, 32'h411ae010} /* (27, 7, 28) {real, imag} */,
  {32'hc0ef584b, 32'h40f36416} /* (27, 7, 27) {real, imag} */,
  {32'hc16841ae, 32'h410995da} /* (27, 7, 26) {real, imag} */,
  {32'h40094871, 32'h413fcd6a} /* (27, 7, 25) {real, imag} */,
  {32'h3e5915b0, 32'h4084e575} /* (27, 7, 24) {real, imag} */,
  {32'hc0d632d0, 32'h40f1eb2c} /* (27, 7, 23) {real, imag} */,
  {32'hc15c1614, 32'h4113531e} /* (27, 7, 22) {real, imag} */,
  {32'h4068dc31, 32'hbf4d5e18} /* (27, 7, 21) {real, imag} */,
  {32'h4156090f, 32'h40211bdc} /* (27, 7, 20) {real, imag} */,
  {32'h41808af6, 32'h411c106f} /* (27, 7, 19) {real, imag} */,
  {32'h4153304f, 32'hbf9f4468} /* (27, 7, 18) {real, imag} */,
  {32'h419708ef, 32'h3f710ef8} /* (27, 7, 17) {real, imag} */,
  {32'h40ebb52b, 32'h3f38d9e0} /* (27, 7, 16) {real, imag} */,
  {32'hc0ff3c96, 32'hc0044a54} /* (27, 7, 15) {real, imag} */,
  {32'hc16db4ce, 32'hc0bcce8f} /* (27, 7, 14) {real, imag} */,
  {32'hc0b95935, 32'h40935811} /* (27, 7, 13) {real, imag} */,
  {32'hc0de7b7e, 32'hc081c2ed} /* (27, 7, 12) {real, imag} */,
  {32'h408cd85b, 32'h40893d66} /* (27, 7, 11) {real, imag} */,
  {32'hc18a8fd0, 32'h412b26f0} /* (27, 7, 10) {real, imag} */,
  {32'hc1406ec4, 32'h3fcb8906} /* (27, 7, 9) {real, imag} */,
  {32'hc0f64914, 32'h40c13011} /* (27, 7, 8) {real, imag} */,
  {32'hc15e30a5, 32'h410e06eb} /* (27, 7, 7) {real, imag} */,
  {32'hc1a03187, 32'h3e841e48} /* (27, 7, 6) {real, imag} */,
  {32'hc18b014e, 32'h4038efb5} /* (27, 7, 5) {real, imag} */,
  {32'hc13d2202, 32'hc077397d} /* (27, 7, 4) {real, imag} */,
  {32'h40bd19f3, 32'h4021d22e} /* (27, 7, 3) {real, imag} */,
  {32'hbee51fb0, 32'h413b155a} /* (27, 7, 2) {real, imag} */,
  {32'h4090fd50, 32'hbfb57660} /* (27, 7, 1) {real, imag} */,
  {32'h412c3982, 32'hbc39c400} /* (27, 7, 0) {real, imag} */,
  {32'hc0fb51e0, 32'hc026ab8d} /* (27, 6, 31) {real, imag} */,
  {32'hc1aac4dc, 32'hc1086ab5} /* (27, 6, 30) {real, imag} */,
  {32'hc1a9752f, 32'hc07b102d} /* (27, 6, 29) {real, imag} */,
  {32'hbf12defc, 32'hc17b4e5b} /* (27, 6, 28) {real, imag} */,
  {32'h41913bbb, 32'hc1fcc08e} /* (27, 6, 27) {real, imag} */,
  {32'h414ca3e1, 32'hc1421e12} /* (27, 6, 26) {real, imag} */,
  {32'hc0e44a3b, 32'hbf534ac0} /* (27, 6, 25) {real, imag} */,
  {32'hc102fe03, 32'h412d1a2b} /* (27, 6, 24) {real, imag} */,
  {32'h414052c8, 32'hc0db3011} /* (27, 6, 23) {real, imag} */,
  {32'h4064cb54, 32'h3dfc2a60} /* (27, 6, 22) {real, imag} */,
  {32'hbfd5a9ff, 32'h4135aeda} /* (27, 6, 21) {real, imag} */,
  {32'h41639221, 32'hbf81d9a6} /* (27, 6, 20) {real, imag} */,
  {32'h41aafc51, 32'hc170b4a5} /* (27, 6, 19) {real, imag} */,
  {32'h40253e0a, 32'hc0e09865} /* (27, 6, 18) {real, imag} */,
  {32'h412fae5f, 32'h403664f8} /* (27, 6, 17) {real, imag} */,
  {32'h41728942, 32'h40dbbb27} /* (27, 6, 16) {real, imag} */,
  {32'h40e3f997, 32'h403f13c0} /* (27, 6, 15) {real, imag} */,
  {32'h3ead96fd, 32'hc171b000} /* (27, 6, 14) {real, imag} */,
  {32'h40b2bf51, 32'h410c92f6} /* (27, 6, 13) {real, imag} */,
  {32'h418da47c, 32'h41655479} /* (27, 6, 12) {real, imag} */,
  {32'hc050426c, 32'hc08cc60a} /* (27, 6, 11) {real, imag} */,
  {32'hc0bcd05e, 32'hc133df60} /* (27, 6, 10) {real, imag} */,
  {32'hc0ddb5b1, 32'hc0d93c1a} /* (27, 6, 9) {real, imag} */,
  {32'h40ee7776, 32'hc1884967} /* (27, 6, 8) {real, imag} */,
  {32'h413f96a6, 32'hc13d6d00} /* (27, 6, 7) {real, imag} */,
  {32'h4147c0f8, 32'hc09aa947} /* (27, 6, 6) {real, imag} */,
  {32'hc11f2a63, 32'hc0094290} /* (27, 6, 5) {real, imag} */,
  {32'hc1a04c1b, 32'h40b538b3} /* (27, 6, 4) {real, imag} */,
  {32'hc15fa2bc, 32'h40e5fd45} /* (27, 6, 3) {real, imag} */,
  {32'hc106b745, 32'hc1129ee2} /* (27, 6, 2) {real, imag} */,
  {32'hc0979d6a, 32'hc184cfd8} /* (27, 6, 1) {real, imag} */,
  {32'hbe9b353a, 32'hc187f398} /* (27, 6, 0) {real, imag} */,
  {32'hc09f78d9, 32'hc0659c12} /* (27, 5, 31) {real, imag} */,
  {32'hc1178b1a, 32'h3f06ae48} /* (27, 5, 30) {real, imag} */,
  {32'hc1a47bc4, 32'h401f186e} /* (27, 5, 29) {real, imag} */,
  {32'hc1d3cde7, 32'hc188bc12} /* (27, 5, 28) {real, imag} */,
  {32'hc1539f46, 32'hc11671ea} /* (27, 5, 27) {real, imag} */,
  {32'h40d30fb6, 32'h4108220d} /* (27, 5, 26) {real, imag} */,
  {32'h40ed371a, 32'h41b122c3} /* (27, 5, 25) {real, imag} */,
  {32'h3ee0e700, 32'hc08d251e} /* (27, 5, 24) {real, imag} */,
  {32'hc1b1e3e4, 32'h405b37d9} /* (27, 5, 23) {real, imag} */,
  {32'hc1215c12, 32'h40e9f384} /* (27, 5, 22) {real, imag} */,
  {32'hc0c7d0c6, 32'h3fdbf6d6} /* (27, 5, 21) {real, imag} */,
  {32'hbfa9f030, 32'h40ef342a} /* (27, 5, 20) {real, imag} */,
  {32'h415f0b9c, 32'h40bbf28c} /* (27, 5, 19) {real, imag} */,
  {32'h40d5e884, 32'h40dd8a72} /* (27, 5, 18) {real, imag} */,
  {32'h408f2f7c, 32'h412ffe05} /* (27, 5, 17) {real, imag} */,
  {32'h40defccb, 32'h41464c4c} /* (27, 5, 16) {real, imag} */,
  {32'hbf01ddd0, 32'h41b87c60} /* (27, 5, 15) {real, imag} */,
  {32'h411fe132, 32'h41706f54} /* (27, 5, 14) {real, imag} */,
  {32'h40f91658, 32'h410c6592} /* (27, 5, 13) {real, imag} */,
  {32'h40358dd5, 32'h413eb972} /* (27, 5, 12) {real, imag} */,
  {32'hc13d048f, 32'h413b01a4} /* (27, 5, 11) {real, imag} */,
  {32'hc0fe3f6c, 32'hc0066ea4} /* (27, 5, 10) {real, imag} */,
  {32'hc0c603f7, 32'hc1a348d6} /* (27, 5, 9) {real, imag} */,
  {32'hc18a9d78, 32'hc20e6d82} /* (27, 5, 8) {real, imag} */,
  {32'hc1ac1bf7, 32'hc1ae59be} /* (27, 5, 7) {real, imag} */,
  {32'h3f9a0660, 32'hc1aad7b9} /* (27, 5, 6) {real, imag} */,
  {32'h410dbc2c, 32'hc1fc95db} /* (27, 5, 5) {real, imag} */,
  {32'hbf921c30, 32'hc19d4a1f} /* (27, 5, 4) {real, imag} */,
  {32'h3e6cfc80, 32'hc1b6cd66} /* (27, 5, 3) {real, imag} */,
  {32'hc1075ed9, 32'hc132444f} /* (27, 5, 2) {real, imag} */,
  {32'hc10abdc0, 32'hc048458b} /* (27, 5, 1) {real, imag} */,
  {32'h40a0304e, 32'hbff1d498} /* (27, 5, 0) {real, imag} */,
  {32'h4016d954, 32'hc0bc621e} /* (27, 4, 31) {real, imag} */,
  {32'hc084c748, 32'hc0f5786b} /* (27, 4, 30) {real, imag} */,
  {32'hc144af16, 32'h410a6dca} /* (27, 4, 29) {real, imag} */,
  {32'h3fc523ee, 32'h4187696c} /* (27, 4, 28) {real, imag} */,
  {32'h3ecc9d10, 32'h412e0032} /* (27, 4, 27) {real, imag} */,
  {32'h4162ae85, 32'h4171cc7f} /* (27, 4, 26) {real, imag} */,
  {32'h40d3f9ce, 32'h41109af6} /* (27, 4, 25) {real, imag} */,
  {32'h413f4262, 32'hc0ec9fe5} /* (27, 4, 24) {real, imag} */,
  {32'h3f28ffc0, 32'hc0d873e5} /* (27, 4, 23) {real, imag} */,
  {32'hbfea6c80, 32'hc0b4f4e0} /* (27, 4, 22) {real, imag} */,
  {32'h41188291, 32'hc1e30548} /* (27, 4, 21) {real, imag} */,
  {32'h41bdb69c, 32'hc22ffc86} /* (27, 4, 20) {real, imag} */,
  {32'h41dff912, 32'hc20b65d6} /* (27, 4, 19) {real, imag} */,
  {32'h4127e734, 32'hc1ab3532} /* (27, 4, 18) {real, imag} */,
  {32'h408223b8, 32'hc198b2e0} /* (27, 4, 17) {real, imag} */,
  {32'hc0311e44, 32'hc10680af} /* (27, 4, 16) {real, imag} */,
  {32'h40f44828, 32'hc15424d6} /* (27, 4, 15) {real, imag} */,
  {32'h4155ac71, 32'hc18b19a0} /* (27, 4, 14) {real, imag} */,
  {32'hc057a7e2, 32'hc1ba52cd} /* (27, 4, 13) {real, imag} */,
  {32'hc158b76e, 32'hc1147412} /* (27, 4, 12) {real, imag} */,
  {32'hc04436a8, 32'hc133f885} /* (27, 4, 11) {real, imag} */,
  {32'h4182e245, 32'h40cf4bec} /* (27, 4, 10) {real, imag} */,
  {32'hbec63460, 32'h41b2a520} /* (27, 4, 9) {real, imag} */,
  {32'hc13f965c, 32'h41d5db9c} /* (27, 4, 8) {real, imag} */,
  {32'hbfd4a940, 32'h3f308700} /* (27, 4, 7) {real, imag} */,
  {32'hc10ff796, 32'h41ac9380} /* (27, 4, 6) {real, imag} */,
  {32'hc0853586, 32'h4108a08f} /* (27, 4, 5) {real, imag} */,
  {32'h3ff176e6, 32'hc0e127d5} /* (27, 4, 4) {real, imag} */,
  {32'h408c7ecb, 32'hc0fa499a} /* (27, 4, 3) {real, imag} */,
  {32'hc025b12c, 32'hc01d3740} /* (27, 4, 2) {real, imag} */,
  {32'hc167f3c0, 32'h403b5be8} /* (27, 4, 1) {real, imag} */,
  {32'hc1081b79, 32'hc0529154} /* (27, 4, 0) {real, imag} */,
  {32'h40d1c523, 32'h41421831} /* (27, 3, 31) {real, imag} */,
  {32'h40990063, 32'h415ef639} /* (27, 3, 30) {real, imag} */,
  {32'hc0ed4d89, 32'h410a9bad} /* (27, 3, 29) {real, imag} */,
  {32'hc13748cb, 32'hc0afb0d7} /* (27, 3, 28) {real, imag} */,
  {32'hc115ed90, 32'h4195a0e4} /* (27, 3, 27) {real, imag} */,
  {32'hc0d63046, 32'hc0c3f891} /* (27, 3, 26) {real, imag} */,
  {32'hc1465bce, 32'hc1c0e272} /* (27, 3, 25) {real, imag} */,
  {32'hc0614af3, 32'hc08f5a78} /* (27, 3, 24) {real, imag} */,
  {32'h4189d1c7, 32'h416a5049} /* (27, 3, 23) {real, imag} */,
  {32'h41899770, 32'h415bff6a} /* (27, 3, 22) {real, imag} */,
  {32'h41652804, 32'hc186f1a9} /* (27, 3, 21) {real, imag} */,
  {32'h41150df2, 32'hc1a20f58} /* (27, 3, 20) {real, imag} */,
  {32'h415797fa, 32'hc0efc4fd} /* (27, 3, 19) {real, imag} */,
  {32'h424f68e3, 32'h402ad69c} /* (27, 3, 18) {real, imag} */,
  {32'h4238cff0, 32'h4108ff90} /* (27, 3, 17) {real, imag} */,
  {32'h41b0de57, 32'h3f1760ec} /* (27, 3, 16) {real, imag} */,
  {32'h41590796, 32'h3e1342e0} /* (27, 3, 15) {real, imag} */,
  {32'hc0f21222, 32'h41ad1413} /* (27, 3, 14) {real, imag} */,
  {32'h4019c142, 32'h4194b550} /* (27, 3, 13) {real, imag} */,
  {32'h415ebeec, 32'h3eed2fc0} /* (27, 3, 12) {real, imag} */,
  {32'h4185aa1e, 32'hbf9dcf78} /* (27, 3, 11) {real, imag} */,
  {32'hc12e6826, 32'h40afcff1} /* (27, 3, 10) {real, imag} */,
  {32'hc1ccadfb, 32'h41075b83} /* (27, 3, 9) {real, imag} */,
  {32'hc03002c7, 32'h41a51e1f} /* (27, 3, 8) {real, imag} */,
  {32'hc0c7dec8, 32'h41b820d2} /* (27, 3, 7) {real, imag} */,
  {32'hc1ed735d, 32'h42028119} /* (27, 3, 6) {real, imag} */,
  {32'hc0c6ecb2, 32'hc0e69752} /* (27, 3, 5) {real, imag} */,
  {32'h40c20216, 32'hc104b0de} /* (27, 3, 4) {real, imag} */,
  {32'h408db512, 32'h40e9f9dd} /* (27, 3, 3) {real, imag} */,
  {32'hbe8aea60, 32'h415b3f16} /* (27, 3, 2) {real, imag} */,
  {32'h4023be54, 32'h3f55ea70} /* (27, 3, 1) {real, imag} */,
  {32'h40935765, 32'h3fbd8bf0} /* (27, 3, 0) {real, imag} */,
  {32'hc1565358, 32'hc1906245} /* (27, 2, 31) {real, imag} */,
  {32'hc1139f17, 32'hc201c38a} /* (27, 2, 30) {real, imag} */,
  {32'h41818a1b, 32'hc25332ac} /* (27, 2, 29) {real, imag} */,
  {32'h4146b7fa, 32'hc2292426} /* (27, 2, 28) {real, imag} */,
  {32'hbf330aa0, 32'hc214f9b2} /* (27, 2, 27) {real, imag} */,
  {32'hc09d85cc, 32'hc2098e8a} /* (27, 2, 26) {real, imag} */,
  {32'hc06c9d80, 32'hc2113984} /* (27, 2, 25) {real, imag} */,
  {32'hc1712681, 32'hc1e8903f} /* (27, 2, 24) {real, imag} */,
  {32'hc1d1702a, 32'hc2110f6b} /* (27, 2, 23) {real, imag} */,
  {32'hc11db018, 32'hc23f75a0} /* (27, 2, 22) {real, imag} */,
  {32'h41386678, 32'hc1d742bf} /* (27, 2, 21) {real, imag} */,
  {32'h41f29fe8, 32'h40772e0a} /* (27, 2, 20) {real, imag} */,
  {32'h4186a597, 32'h41e13660} /* (27, 2, 19) {real, imag} */,
  {32'h41d52280, 32'h41a646a2} /* (27, 2, 18) {real, imag} */,
  {32'h423be7a7, 32'h41bb558f} /* (27, 2, 17) {real, imag} */,
  {32'h425c1097, 32'h41b11cec} /* (27, 2, 16) {real, imag} */,
  {32'h419c9259, 32'h41bb88d0} /* (27, 2, 15) {real, imag} */,
  {32'h40bf2046, 32'h42024056} /* (27, 2, 14) {real, imag} */,
  {32'h41259904, 32'h41e681c0} /* (27, 2, 13) {real, imag} */,
  {32'h41b98eb2, 32'h4124a2fe} /* (27, 2, 12) {real, imag} */,
  {32'h42085645, 32'h4090d7c6} /* (27, 2, 11) {real, imag} */,
  {32'hc092348e, 32'hc15427d1} /* (27, 2, 10) {real, imag} */,
  {32'hc1a87558, 32'hc20f8550} /* (27, 2, 9) {real, imag} */,
  {32'hc2061445, 32'hc2594513} /* (27, 2, 8) {real, imag} */,
  {32'hc1571d46, 32'hc20b96bc} /* (27, 2, 7) {real, imag} */,
  {32'hc071412b, 32'hc1c0f3a2} /* (27, 2, 6) {real, imag} */,
  {32'hc0fd6dfe, 32'hc18d61bb} /* (27, 2, 5) {real, imag} */,
  {32'hc100c96a, 32'hc1b54386} /* (27, 2, 4) {real, imag} */,
  {32'hc189cfc2, 32'hc177aa7a} /* (27, 2, 3) {real, imag} */,
  {32'hc162a41f, 32'hc0ffdf19} /* (27, 2, 2) {real, imag} */,
  {32'hc17e4a25, 32'hc1db31d2} /* (27, 2, 1) {real, imag} */,
  {32'hc06d42eb, 32'hc20500ce} /* (27, 2, 0) {real, imag} */,
  {32'h40f0b81e, 32'h413fcfa9} /* (27, 1, 31) {real, imag} */,
  {32'h41b01f16, 32'h41f22923} /* (27, 1, 30) {real, imag} */,
  {32'h41c5b21e, 32'h422e928a} /* (27, 1, 29) {real, imag} */,
  {32'h40831298, 32'h424faf03} /* (27, 1, 28) {real, imag} */,
  {32'h40f42aac, 32'h42651664} /* (27, 1, 27) {real, imag} */,
  {32'h3f1db780, 32'h420f20bf} /* (27, 1, 26) {real, imag} */,
  {32'h417d6801, 32'h420650c7} /* (27, 1, 25) {real, imag} */,
  {32'h41d1a7bc, 32'h421a0fee} /* (27, 1, 24) {real, imag} */,
  {32'h41d67649, 32'h425585b2} /* (27, 1, 23) {real, imag} */,
  {32'h42121dee, 32'h42674deb} /* (27, 1, 22) {real, imag} */,
  {32'h40d05913, 32'h41ba36b7} /* (27, 1, 21) {real, imag} */,
  {32'hc0d6f8de, 32'hc100bb60} /* (27, 1, 20) {real, imag} */,
  {32'hc17fc930, 32'hc0476842} /* (27, 1, 19) {real, imag} */,
  {32'hc0e48696, 32'h3ef30258} /* (27, 1, 18) {real, imag} */,
  {32'hc0ac8542, 32'hc1a40716} /* (27, 1, 17) {real, imag} */,
  {32'h400e0282, 32'hc1bce76e} /* (27, 1, 16) {real, imag} */,
  {32'hc0b89af4, 32'hc1e4c922} /* (27, 1, 15) {real, imag} */,
  {32'hc1321fb6, 32'hc129692f} /* (27, 1, 14) {real, imag} */,
  {32'hc184e75c, 32'hc1e785d0} /* (27, 1, 13) {real, imag} */,
  {32'hc1be54e8, 32'hc255d7a9} /* (27, 1, 12) {real, imag} */,
  {32'hc1a6f8eb, 32'hc2316608} /* (27, 1, 11) {real, imag} */,
  {32'hc0e3d9d0, 32'h40bf5cf7} /* (27, 1, 10) {real, imag} */,
  {32'hc0152810, 32'h419ab767} /* (27, 1, 9) {real, imag} */,
  {32'hc1c23328, 32'h41a2e8a2} /* (27, 1, 8) {real, imag} */,
  {32'hc194b69b, 32'h41bece02} /* (27, 1, 7) {real, imag} */,
  {32'h3e9bdec8, 32'h4234b65b} /* (27, 1, 6) {real, imag} */,
  {32'h419a0606, 32'h42513ec0} /* (27, 1, 5) {real, imag} */,
  {32'h41f734cc, 32'h41c738c6} /* (27, 1, 4) {real, imag} */,
  {32'h4186846f, 32'h41d32f87} /* (27, 1, 3) {real, imag} */,
  {32'h41f9fb38, 32'h4213d026} /* (27, 1, 2) {real, imag} */,
  {32'h41f8f920, 32'h422c04f4} /* (27, 1, 1) {real, imag} */,
  {32'h41a30c1c, 32'h41a10bd4} /* (27, 1, 0) {real, imag} */,
  {32'h41611409, 32'h4148be62} /* (27, 0, 31) {real, imag} */,
  {32'h41f8ecc2, 32'h41aa2c05} /* (27, 0, 30) {real, imag} */,
  {32'hc0b20224, 32'h421fdc14} /* (27, 0, 29) {real, imag} */,
  {32'h41433a24, 32'h4206cffa} /* (27, 0, 28) {real, imag} */,
  {32'h423bb37e, 32'h41c3ac3d} /* (27, 0, 27) {real, imag} */,
  {32'h41f8e70e, 32'h41a2ac53} /* (27, 0, 26) {real, imag} */,
  {32'h4126a142, 32'h41972bec} /* (27, 0, 25) {real, imag} */,
  {32'h412d1ae8, 32'h420d4118} /* (27, 0, 24) {real, imag} */,
  {32'h40ce80ae, 32'h415348a7} /* (27, 0, 23) {real, imag} */,
  {32'h40ebce48, 32'h41c6ffa4} /* (27, 0, 22) {real, imag} */,
  {32'h40cdcb69, 32'h42146619} /* (27, 0, 21) {real, imag} */,
  {32'h41579cba, 32'h418733a3} /* (27, 0, 20) {real, imag} */,
  {32'hbdf79c20, 32'h415150ca} /* (27, 0, 19) {real, imag} */,
  {32'h408f5bd0, 32'hbeeb50b0} /* (27, 0, 18) {real, imag} */,
  {32'hc1b8a78f, 32'h3c8ecc00} /* (27, 0, 17) {real, imag} */,
  {32'hc13ca061, 32'h3f2adec8} /* (27, 0, 16) {real, imag} */,
  {32'hc10ddb7e, 32'hc1cf7988} /* (27, 0, 15) {real, imag} */,
  {32'hc1e8499a, 32'hc1cc610e} /* (27, 0, 14) {real, imag} */,
  {32'hc20247fb, 32'hc1d24e7c} /* (27, 0, 13) {real, imag} */,
  {32'hc1aa7bac, 32'hc1ed0182} /* (27, 0, 12) {real, imag} */,
  {32'hc19d35bc, 32'hc1b6777c} /* (27, 0, 11) {real, imag} */,
  {32'hc16c6528, 32'h40b89200} /* (27, 0, 10) {real, imag} */,
  {32'hc0f64cd4, 32'h3fa2d1c6} /* (27, 0, 9) {real, imag} */,
  {32'h415ac5e8, 32'h4112afe1} /* (27, 0, 8) {real, imag} */,
  {32'h40a9de79, 32'h4005c133} /* (27, 0, 7) {real, imag} */,
  {32'hc0973804, 32'h40edb170} /* (27, 0, 6) {real, imag} */,
  {32'hc0dc60dc, 32'h420d61af} /* (27, 0, 5) {real, imag} */,
  {32'hc112d9f6, 32'h4207ed83} /* (27, 0, 4) {real, imag} */,
  {32'h40874cdd, 32'h42043b9a} /* (27, 0, 3) {real, imag} */,
  {32'h41a5f5d8, 32'h414be5d4} /* (27, 0, 2) {real, imag} */,
  {32'h3fcf4be8, 32'h40eaa5b0} /* (27, 0, 1) {real, imag} */,
  {32'hbe962a8c, 32'h415dc0dc} /* (27, 0, 0) {real, imag} */,
  {32'h411faa00, 32'hbfda2ff8} /* (26, 31, 31) {real, imag} */,
  {32'h416e7c65, 32'hbfc559ca} /* (26, 31, 30) {real, imag} */,
  {32'hc0a5221c, 32'hbefafeb0} /* (26, 31, 29) {real, imag} */,
  {32'h40a18041, 32'h419ce0d3} /* (26, 31, 28) {real, imag} */,
  {32'h41762b6e, 32'h40461fb4} /* (26, 31, 27) {real, imag} */,
  {32'h41921260, 32'hc086359e} /* (26, 31, 26) {real, imag} */,
  {32'h419ecb7a, 32'h3f18427c} /* (26, 31, 25) {real, imag} */,
  {32'h4135fd88, 32'h4056d9fc} /* (26, 31, 24) {real, imag} */,
  {32'h410122db, 32'h4138864a} /* (26, 31, 23) {real, imag} */,
  {32'hbfe11474, 32'h408d6a36} /* (26, 31, 22) {real, imag} */,
  {32'hc0871573, 32'h418a9048} /* (26, 31, 21) {real, imag} */,
  {32'hc07b0302, 32'h415c442e} /* (26, 31, 20) {real, imag} */,
  {32'h419bdd83, 32'h40d45078} /* (26, 31, 19) {real, imag} */,
  {32'hc0d2f246, 32'h404d8290} /* (26, 31, 18) {real, imag} */,
  {32'h414257ef, 32'h41368deb} /* (26, 31, 17) {real, imag} */,
  {32'h41921cef, 32'h40dee017} /* (26, 31, 16) {real, imag} */,
  {32'hc0df388c, 32'hc196147a} /* (26, 31, 15) {real, imag} */,
  {32'hbf06fd58, 32'h40691630} /* (26, 31, 14) {real, imag} */,
  {32'hc12323d7, 32'hbe9a2050} /* (26, 31, 13) {real, imag} */,
  {32'hc0d88c40, 32'h409a22b0} /* (26, 31, 12) {real, imag} */,
  {32'h40b64b3a, 32'h4144fc20} /* (26, 31, 11) {real, imag} */,
  {32'h412c8c60, 32'hbe913ac0} /* (26, 31, 10) {real, imag} */,
  {32'h416bc3aa, 32'hc09b13e9} /* (26, 31, 9) {real, imag} */,
  {32'h4092e2b7, 32'hc119b244} /* (26, 31, 8) {real, imag} */,
  {32'h41be2263, 32'h3e235840} /* (26, 31, 7) {real, imag} */,
  {32'h41183aff, 32'h3fb34ad8} /* (26, 31, 6) {real, imag} */,
  {32'hc10f34e1, 32'h3f01de46} /* (26, 31, 5) {real, imag} */,
  {32'hc149c6f9, 32'h4121cf95} /* (26, 31, 4) {real, imag} */,
  {32'hc0a1ac15, 32'h40878f76} /* (26, 31, 3) {real, imag} */,
  {32'hc0062024, 32'hc04d0478} /* (26, 31, 2) {real, imag} */,
  {32'hc005fd6c, 32'h41834d9a} /* (26, 31, 1) {real, imag} */,
  {32'h3fa126b4, 32'h40b1db62} /* (26, 31, 0) {real, imag} */,
  {32'h40d5733b, 32'h41368c98} /* (26, 30, 31) {real, imag} */,
  {32'h41457f73, 32'h41a621bc} /* (26, 30, 30) {real, imag} */,
  {32'h410eb998, 32'h40d11a74} /* (26, 30, 29) {real, imag} */,
  {32'h405cba7b, 32'hc16b536a} /* (26, 30, 28) {real, imag} */,
  {32'hc1010c17, 32'hc1c6ff32} /* (26, 30, 27) {real, imag} */,
  {32'hc0602a40, 32'hc1b6fbc4} /* (26, 30, 26) {real, imag} */,
  {32'hc0dd92c4, 32'hc1cb514e} /* (26, 30, 25) {real, imag} */,
  {32'hc1172d66, 32'hc1c49bee} /* (26, 30, 24) {real, imag} */,
  {32'h41023df4, 32'h408621fb} /* (26, 30, 23) {real, imag} */,
  {32'h4189ed30, 32'hc07d8670} /* (26, 30, 22) {real, imag} */,
  {32'h4021f8e0, 32'hc142729c} /* (26, 30, 21) {real, imag} */,
  {32'hc13b337e, 32'h4175eef3} /* (26, 30, 20) {real, imag} */,
  {32'hc14803cc, 32'h4181944c} /* (26, 30, 19) {real, imag} */,
  {32'hc19ef69f, 32'hbf3131c8} /* (26, 30, 18) {real, imag} */,
  {32'hc15113de, 32'hc0d83404} /* (26, 30, 17) {real, imag} */,
  {32'hc1281ab6, 32'h4119c9f8} /* (26, 30, 16) {real, imag} */,
  {32'hc0b26899, 32'h41e8da1d} /* (26, 30, 15) {real, imag} */,
  {32'h3f035080, 32'h416e7148} /* (26, 30, 14) {real, imag} */,
  {32'hc0cbe9b4, 32'hc1042ad6} /* (26, 30, 13) {real, imag} */,
  {32'hc0daa818, 32'hc041b27f} /* (26, 30, 12) {real, imag} */,
  {32'hc19405eb, 32'h4168e06b} /* (26, 30, 11) {real, imag} */,
  {32'hc173b69c, 32'h41d88082} /* (26, 30, 10) {real, imag} */,
  {32'hc07c5bd0, 32'h41f5e5eb} /* (26, 30, 9) {real, imag} */,
  {32'h3ecf5110, 32'h4158ee90} /* (26, 30, 8) {real, imag} */,
  {32'hc13cd110, 32'h41acb77b} /* (26, 30, 7) {real, imag} */,
  {32'hc087c48a, 32'h41afdec2} /* (26, 30, 6) {real, imag} */,
  {32'h418f83e8, 32'h40898306} /* (26, 30, 5) {real, imag} */,
  {32'h4172e22a, 32'h406c9e47} /* (26, 30, 4) {real, imag} */,
  {32'h40b13d0a, 32'h4186faa7} /* (26, 30, 3) {real, imag} */,
  {32'h40f19f10, 32'h414bbee0} /* (26, 30, 2) {real, imag} */,
  {32'hc0910ae0, 32'h40a7ab38} /* (26, 30, 1) {real, imag} */,
  {32'hc09a5679, 32'hbfe0357a} /* (26, 30, 0) {real, imag} */,
  {32'hbf1c4234, 32'hc14c8ea4} /* (26, 29, 31) {real, imag} */,
  {32'h40b9262d, 32'hc14a1181} /* (26, 29, 30) {real, imag} */,
  {32'hc0d412c1, 32'hc010fcbc} /* (26, 29, 29) {real, imag} */,
  {32'h40adc20c, 32'hbfe1d570} /* (26, 29, 28) {real, imag} */,
  {32'h40775778, 32'hbffba9e4} /* (26, 29, 27) {real, imag} */,
  {32'hc0a0995a, 32'hc038c370} /* (26, 29, 26) {real, imag} */,
  {32'hc137c16e, 32'h416a1e80} /* (26, 29, 25) {real, imag} */,
  {32'hc18bb5ed, 32'hbefd32a0} /* (26, 29, 24) {real, imag} */,
  {32'hc1cbc976, 32'h3f9ecf40} /* (26, 29, 23) {real, imag} */,
  {32'hc18da45c, 32'hc09bde83} /* (26, 29, 22) {real, imag} */,
  {32'hc1592f37, 32'hc162d853} /* (26, 29, 21) {real, imag} */,
  {32'hc194db4c, 32'hc11a697e} /* (26, 29, 20) {real, imag} */,
  {32'hc19c2555, 32'h40cd02de} /* (26, 29, 19) {real, imag} */,
  {32'h4030ec54, 32'h411a3104} /* (26, 29, 18) {real, imag} */,
  {32'h3f59953e, 32'hc12f58ac} /* (26, 29, 17) {real, imag} */,
  {32'h3f23c228, 32'hc083849e} /* (26, 29, 16) {real, imag} */,
  {32'h41157a4c, 32'hc06d09d3} /* (26, 29, 15) {real, imag} */,
  {32'hbef78b48, 32'h41283b03} /* (26, 29, 14) {real, imag} */,
  {32'hbfdbcf5e, 32'h419e20e6} /* (26, 29, 13) {real, imag} */,
  {32'h4105f7b4, 32'h3fba93b6} /* (26, 29, 12) {real, imag} */,
  {32'hc1784728, 32'hc13f5622} /* (26, 29, 11) {real, imag} */,
  {32'hbfa30d4f, 32'hc1820d70} /* (26, 29, 10) {real, imag} */,
  {32'h41271766, 32'hc1738f7c} /* (26, 29, 9) {real, imag} */,
  {32'h409842be, 32'hc18dc0cb} /* (26, 29, 8) {real, imag} */,
  {32'h414b248f, 32'h4047c4f8} /* (26, 29, 7) {real, imag} */,
  {32'h41352d41, 32'hc08c1ae0} /* (26, 29, 6) {real, imag} */,
  {32'hc1128503, 32'hbf8b91a5} /* (26, 29, 5) {real, imag} */,
  {32'h3efaa748, 32'hbed35a10} /* (26, 29, 4) {real, imag} */,
  {32'h41486f5d, 32'hc0d31e04} /* (26, 29, 3) {real, imag} */,
  {32'h4138c7ae, 32'hc13d3fa4} /* (26, 29, 2) {real, imag} */,
  {32'h41383870, 32'h40c468e5} /* (26, 29, 1) {real, imag} */,
  {32'h41177bc9, 32'h40cebf74} /* (26, 29, 0) {real, imag} */,
  {32'hbf628828, 32'h40d2f89c} /* (26, 28, 31) {real, imag} */,
  {32'h416a1673, 32'h40c178ac} /* (26, 28, 30) {real, imag} */,
  {32'h409164c4, 32'hc121fca2} /* (26, 28, 29) {real, imag} */,
  {32'hc0eab624, 32'hc11a8dd6} /* (26, 28, 28) {real, imag} */,
  {32'h412b5b4f, 32'hc127d73d} /* (26, 28, 27) {real, imag} */,
  {32'h41b5fe04, 32'hc0a91c56} /* (26, 28, 26) {real, imag} */,
  {32'h417087f5, 32'hbf3b4e8c} /* (26, 28, 25) {real, imag} */,
  {32'hc01bbeca, 32'hc09b282e} /* (26, 28, 24) {real, imag} */,
  {32'hc083ff9a, 32'h4189a918} /* (26, 28, 23) {real, imag} */,
  {32'hc15f4762, 32'h41e857b2} /* (26, 28, 22) {real, imag} */,
  {32'hc180a836, 32'h41ccf3e6} /* (26, 28, 21) {real, imag} */,
  {32'h411285d2, 32'h41ad468a} /* (26, 28, 20) {real, imag} */,
  {32'h411aa412, 32'h3ea03b60} /* (26, 28, 19) {real, imag} */,
  {32'hc092a08a, 32'hc19b75b0} /* (26, 28, 18) {real, imag} */,
  {32'hc0a03eb2, 32'hc0fc7460} /* (26, 28, 17) {real, imag} */,
  {32'h41312c8f, 32'h40b9261c} /* (26, 28, 16) {real, imag} */,
  {32'hc0d40007, 32'hc0bccd37} /* (26, 28, 15) {real, imag} */,
  {32'hc180488f, 32'h406b7e72} /* (26, 28, 14) {real, imag} */,
  {32'h3fdf6a08, 32'h40eb25d0} /* (26, 28, 13) {real, imag} */,
  {32'h412b9508, 32'h41745070} /* (26, 28, 12) {real, imag} */,
  {32'h413afc7e, 32'h41298160} /* (26, 28, 11) {real, imag} */,
  {32'h415ec53c, 32'h3eee12a0} /* (26, 28, 10) {real, imag} */,
  {32'hbfa43684, 32'h3e26e5f8} /* (26, 28, 9) {real, imag} */,
  {32'hc035ae5c, 32'hbe84dd18} /* (26, 28, 8) {real, imag} */,
  {32'h3f5a29cd, 32'hc1b0db76} /* (26, 28, 7) {real, imag} */,
  {32'h412446ee, 32'hc014558c} /* (26, 28, 6) {real, imag} */,
  {32'h40db83c4, 32'h40618e9e} /* (26, 28, 5) {real, imag} */,
  {32'h40826718, 32'hc0dd6828} /* (26, 28, 4) {real, imag} */,
  {32'h4141f036, 32'hc1908bab} /* (26, 28, 3) {real, imag} */,
  {32'h40f3c6de, 32'hbf881d48} /* (26, 28, 2) {real, imag} */,
  {32'h40a4c0c8, 32'h4134a6fc} /* (26, 28, 1) {real, imag} */,
  {32'hc0695a02, 32'h4023ba81} /* (26, 28, 0) {real, imag} */,
  {32'h40ba98b6, 32'h3fdb9239} /* (26, 27, 31) {real, imag} */,
  {32'hc134ae80, 32'h405d5a98} /* (26, 27, 30) {real, imag} */,
  {32'hc178eeb5, 32'h40e61de0} /* (26, 27, 29) {real, imag} */,
  {32'hc19a8424, 32'h40696d82} /* (26, 27, 28) {real, imag} */,
  {32'h403dd23c, 32'hbdbb5ce0} /* (26, 27, 27) {real, imag} */,
  {32'h400fbe5f, 32'h3fa00517} /* (26, 27, 26) {real, imag} */,
  {32'h40cceec5, 32'hc0ef2e74} /* (26, 27, 25) {real, imag} */,
  {32'hc1a1bfea, 32'hc1770bde} /* (26, 27, 24) {real, imag} */,
  {32'hc11c857e, 32'hc1a6afd6} /* (26, 27, 23) {real, imag} */,
  {32'hc151d7b1, 32'hc0064a10} /* (26, 27, 22) {real, imag} */,
  {32'hc1871d05, 32'h412d8e22} /* (26, 27, 21) {real, imag} */,
  {32'hc1b50858, 32'h418f8ad4} /* (26, 27, 20) {real, imag} */,
  {32'hc085e712, 32'h4146ef67} /* (26, 27, 19) {real, imag} */,
  {32'h40ddc392, 32'hbeca7598} /* (26, 27, 18) {real, imag} */,
  {32'h41120116, 32'h40c0ffe2} /* (26, 27, 17) {real, imag} */,
  {32'hc1066a59, 32'hc121cd13} /* (26, 27, 16) {real, imag} */,
  {32'hc09aa362, 32'hc174ad8d} /* (26, 27, 15) {real, imag} */,
  {32'hc103f04d, 32'h40d26dfe} /* (26, 27, 14) {real, imag} */,
  {32'hc11d7c80, 32'hc14066ab} /* (26, 27, 13) {real, imag} */,
  {32'hc094b811, 32'hc10801a2} /* (26, 27, 12) {real, imag} */,
  {32'hc12ef74e, 32'h3f39f5a0} /* (26, 27, 11) {real, imag} */,
  {32'hc159c5f7, 32'hc19d0fde} /* (26, 27, 10) {real, imag} */,
  {32'hc09e140e, 32'hc1be8526} /* (26, 27, 9) {real, imag} */,
  {32'h40014661, 32'hc02b8912} /* (26, 27, 8) {real, imag} */,
  {32'hbf13ff18, 32'h3f741340} /* (26, 27, 7) {real, imag} */,
  {32'hc06b091c, 32'h3fa2ff35} /* (26, 27, 6) {real, imag} */,
  {32'h41190ee4, 32'hbf4b6580} /* (26, 27, 5) {real, imag} */,
  {32'h40a328b3, 32'h4152e158} /* (26, 27, 4) {real, imag} */,
  {32'h40ecd88c, 32'h415f8587} /* (26, 27, 3) {real, imag} */,
  {32'h419a5463, 32'hc10de52f} /* (26, 27, 2) {real, imag} */,
  {32'hc00d9197, 32'hc16c92d2} /* (26, 27, 1) {real, imag} */,
  {32'hc10e566c, 32'h4061051e} /* (26, 27, 0) {real, imag} */,
  {32'h40021202, 32'h3f451580} /* (26, 26, 31) {real, imag} */,
  {32'hbfc602e2, 32'hc0cbf762} /* (26, 26, 30) {real, imag} */,
  {32'hc01ecca2, 32'h40adc50c} /* (26, 26, 29) {real, imag} */,
  {32'hbf0868f8, 32'h4155b336} /* (26, 26, 28) {real, imag} */,
  {32'hbeac6050, 32'h41beb212} /* (26, 26, 27) {real, imag} */,
  {32'h40d1939a, 32'h3d8de780} /* (26, 26, 26) {real, imag} */,
  {32'h41849b24, 32'hc11bcde0} /* (26, 26, 25) {real, imag} */,
  {32'h419969b2, 32'h41881d85} /* (26, 26, 24) {real, imag} */,
  {32'h40e3993f, 32'h3dd8c3e0} /* (26, 26, 23) {real, imag} */,
  {32'hc0f81279, 32'hbfa9da74} /* (26, 26, 22) {real, imag} */,
  {32'hc1062cac, 32'h4100eaee} /* (26, 26, 21) {real, imag} */,
  {32'hc126008a, 32'hbfa9dfca} /* (26, 26, 20) {real, imag} */,
  {32'h40cd9ff2, 32'hc071a5f7} /* (26, 26, 19) {real, imag} */,
  {32'h41061ad2, 32'h4094ae3b} /* (26, 26, 18) {real, imag} */,
  {32'hc0e357a6, 32'h412d1eae} /* (26, 26, 17) {real, imag} */,
  {32'hc1909b01, 32'hc11625e8} /* (26, 26, 16) {real, imag} */,
  {32'hc013fed5, 32'hc067739c} /* (26, 26, 15) {real, imag} */,
  {32'hc0e5d31b, 32'h413302da} /* (26, 26, 14) {real, imag} */,
  {32'hc11b3a04, 32'h41ab3c00} /* (26, 26, 13) {real, imag} */,
  {32'h4114d28b, 32'hc07e063c} /* (26, 26, 12) {real, imag} */,
  {32'h410aee29, 32'h4038e1cc} /* (26, 26, 11) {real, imag} */,
  {32'h4188ac4c, 32'h419d70e0} /* (26, 26, 10) {real, imag} */,
  {32'h40ed880e, 32'h4141c43e} /* (26, 26, 9) {real, imag} */,
  {32'hc109095b, 32'h3ee4eaf0} /* (26, 26, 8) {real, imag} */,
  {32'hc1965d60, 32'hc10b1937} /* (26, 26, 7) {real, imag} */,
  {32'hc102a7fe, 32'hc1a98048} /* (26, 26, 6) {real, imag} */,
  {32'h41170512, 32'hc04b1004} /* (26, 26, 5) {real, imag} */,
  {32'hc03217a2, 32'hc08ddcbb} /* (26, 26, 4) {real, imag} */,
  {32'hc17296c3, 32'hbfcfd22e} /* (26, 26, 3) {real, imag} */,
  {32'hc012a516, 32'hbf0d98e0} /* (26, 26, 2) {real, imag} */,
  {32'h3f53b158, 32'h415125c2} /* (26, 26, 1) {real, imag} */,
  {32'hc071e7ec, 32'h40dfbf14} /* (26, 26, 0) {real, imag} */,
  {32'h41483cd0, 32'hc0045fe9} /* (26, 25, 31) {real, imag} */,
  {32'h4012cf49, 32'h40b9183c} /* (26, 25, 30) {real, imag} */,
  {32'hbea4b71e, 32'h4062ceb7} /* (26, 25, 29) {real, imag} */,
  {32'hc11429e0, 32'h3fe7242c} /* (26, 25, 28) {real, imag} */,
  {32'hc19cec82, 32'hc071d218} /* (26, 25, 27) {real, imag} */,
  {32'hc0bf9979, 32'hc177b7ef} /* (26, 25, 26) {real, imag} */,
  {32'hc1238dd2, 32'h3cdd7a00} /* (26, 25, 25) {real, imag} */,
  {32'hc0655783, 32'h412bf66a} /* (26, 25, 24) {real, imag} */,
  {32'h4125ea92, 32'h408bb9b9} /* (26, 25, 23) {real, imag} */,
  {32'h40a65e84, 32'hc0feb5b0} /* (26, 25, 22) {real, imag} */,
  {32'hc1c4d270, 32'h4138eb2f} /* (26, 25, 21) {real, imag} */,
  {32'hc1c6ca62, 32'h41428c52} /* (26, 25, 20) {real, imag} */,
  {32'hc1c18400, 32'h41b14c4e} /* (26, 25, 19) {real, imag} */,
  {32'hc093ef16, 32'h41a06440} /* (26, 25, 18) {real, imag} */,
  {32'hbec68e30, 32'h410c9106} /* (26, 25, 17) {real, imag} */,
  {32'hbf0d3c20, 32'h41408919} /* (26, 25, 16) {real, imag} */,
  {32'hc0e9ec3c, 32'h4161cff4} /* (26, 25, 15) {real, imag} */,
  {32'h402b77ac, 32'h40cf37cc} /* (26, 25, 14) {real, imag} */,
  {32'hbf7d8a04, 32'h40d1adaf} /* (26, 25, 13) {real, imag} */,
  {32'h401b4d1e, 32'hc0dbe295} /* (26, 25, 12) {real, imag} */,
  {32'h409fb32b, 32'hc13e534e} /* (26, 25, 11) {real, imag} */,
  {32'h41cbfd72, 32'hc001985a} /* (26, 25, 10) {real, imag} */,
  {32'h41af0efc, 32'h4081285a} /* (26, 25, 9) {real, imag} */,
  {32'h40325828, 32'h4038581a} /* (26, 25, 8) {real, imag} */,
  {32'hbeff5d60, 32'h41819063} /* (26, 25, 7) {real, imag} */,
  {32'hc0deb3ba, 32'h41b56d31} /* (26, 25, 6) {real, imag} */,
  {32'hc14c072f, 32'h40dbacc0} /* (26, 25, 5) {real, imag} */,
  {32'hc1566b74, 32'h3fee291c} /* (26, 25, 4) {real, imag} */,
  {32'hc0878fbe, 32'h411123cb} /* (26, 25, 3) {real, imag} */,
  {32'hc0f15a76, 32'hc011b4f2} /* (26, 25, 2) {real, imag} */,
  {32'h4177f768, 32'h405cc22c} /* (26, 25, 1) {real, imag} */,
  {32'h4142cbc5, 32'h40c1fc34} /* (26, 25, 0) {real, imag} */,
  {32'hc0bae6c6, 32'hc04728be} /* (26, 24, 31) {real, imag} */,
  {32'hc01df2b3, 32'hc09d1147} /* (26, 24, 30) {real, imag} */,
  {32'h412c3616, 32'hc0c1d3ec} /* (26, 24, 29) {real, imag} */,
  {32'h4175c84f, 32'hc15e39ad} /* (26, 24, 28) {real, imag} */,
  {32'h4069c675, 32'hc1264735} /* (26, 24, 27) {real, imag} */,
  {32'hc1045ef8, 32'h3fcece14} /* (26, 24, 26) {real, imag} */,
  {32'hc0b1c018, 32'hbeac18a0} /* (26, 24, 25) {real, imag} */,
  {32'h4156bbd6, 32'h41000363} /* (26, 24, 24) {real, imag} */,
  {32'hc09d3cea, 32'h402243db} /* (26, 24, 23) {real, imag} */,
  {32'h4015e218, 32'hc0264048} /* (26, 24, 22) {real, imag} */,
  {32'h40be8654, 32'hc0305be8} /* (26, 24, 21) {real, imag} */,
  {32'hc0e71d94, 32'hc067e8e8} /* (26, 24, 20) {real, imag} */,
  {32'hc12de85b, 32'h41401ed3} /* (26, 24, 19) {real, imag} */,
  {32'hc0925376, 32'h418b8e97} /* (26, 24, 18) {real, imag} */,
  {32'h4151b1ce, 32'h40bf2d74} /* (26, 24, 17) {real, imag} */,
  {32'hbea53800, 32'h400614ee} /* (26, 24, 16) {real, imag} */,
  {32'hc0c7021a, 32'h40346608} /* (26, 24, 15) {real, imag} */,
  {32'h41685d89, 32'h413606cf} /* (26, 24, 14) {real, imag} */,
  {32'h41753108, 32'h40b00bbe} /* (26, 24, 13) {real, imag} */,
  {32'h40a3215c, 32'hbd9f2cc0} /* (26, 24, 12) {real, imag} */,
  {32'h4039b764, 32'h3c18ca00} /* (26, 24, 11) {real, imag} */,
  {32'hc05b15c0, 32'hc091d1a0} /* (26, 24, 10) {real, imag} */,
  {32'hc0cb0af1, 32'h40a1d978} /* (26, 24, 9) {real, imag} */,
  {32'hc15dcd24, 32'h4181887b} /* (26, 24, 8) {real, imag} */,
  {32'hc13f6cd4, 32'h40b02c6b} /* (26, 24, 7) {real, imag} */,
  {32'hc10b07e1, 32'hc0c4f114} /* (26, 24, 6) {real, imag} */,
  {32'h3f128888, 32'hc0ac8fdb} /* (26, 24, 5) {real, imag} */,
  {32'h418cdb01, 32'hbf3f0808} /* (26, 24, 4) {real, imag} */,
  {32'h4104f301, 32'h3f9b7fdc} /* (26, 24, 3) {real, imag} */,
  {32'h3f0c8b98, 32'hc06e4628} /* (26, 24, 2) {real, imag} */,
  {32'hc0c5747a, 32'hc0d5b2f6} /* (26, 24, 1) {real, imag} */,
  {32'hc143c704, 32'hbf26b180} /* (26, 24, 0) {real, imag} */,
  {32'hc05faf75, 32'hbfbcd916} /* (26, 23, 31) {real, imag} */,
  {32'hc107b7e6, 32'hbfac2ffc} /* (26, 23, 30) {real, imag} */,
  {32'h3ef1ac60, 32'h40c99cb6} /* (26, 23, 29) {real, imag} */,
  {32'h41495db8, 32'h40bc3a05} /* (26, 23, 28) {real, imag} */,
  {32'h3e958680, 32'hbfd66dac} /* (26, 23, 27) {real, imag} */,
  {32'hc09c5f1c, 32'hc102ee92} /* (26, 23, 26) {real, imag} */,
  {32'hbf2c1210, 32'hc0fa0d26} /* (26, 23, 25) {real, imag} */,
  {32'h3fa917b8, 32'hc18bb278} /* (26, 23, 24) {real, imag} */,
  {32'hc13a392d, 32'hc18b7348} /* (26, 23, 23) {real, imag} */,
  {32'hc15999e4, 32'hc15c0a8a} /* (26, 23, 22) {real, imag} */,
  {32'hc0d931d4, 32'hc08aeaa5} /* (26, 23, 21) {real, imag} */,
  {32'h3f792508, 32'hc1031c38} /* (26, 23, 20) {real, imag} */,
  {32'h41023b0c, 32'hc0ca9470} /* (26, 23, 19) {real, imag} */,
  {32'hbf1d8f20, 32'h40c0e2fb} /* (26, 23, 18) {real, imag} */,
  {32'hbf710a48, 32'h40d5c144} /* (26, 23, 17) {real, imag} */,
  {32'hc0b0f0d5, 32'h40a59c63} /* (26, 23, 16) {real, imag} */,
  {32'h41019b44, 32'hc025708a} /* (26, 23, 15) {real, imag} */,
  {32'h4173174c, 32'hc0789105} /* (26, 23, 14) {real, imag} */,
  {32'hbe4a25e8, 32'hc0f04fef} /* (26, 23, 13) {real, imag} */,
  {32'h40840cff, 32'hc1180784} /* (26, 23, 12) {real, imag} */,
  {32'h413688f2, 32'hc182fb08} /* (26, 23, 11) {real, imag} */,
  {32'h3fe15288, 32'hc09da81f} /* (26, 23, 10) {real, imag} */,
  {32'hc04349da, 32'h40564863} /* (26, 23, 9) {real, imag} */,
  {32'hc091209e, 32'hbff8516a} /* (26, 23, 8) {real, imag} */,
  {32'hc0be1580, 32'h3f07b7ec} /* (26, 23, 7) {real, imag} */,
  {32'hc085e746, 32'hc141fa5c} /* (26, 23, 6) {real, imag} */,
  {32'h408b3b18, 32'hc172c845} /* (26, 23, 5) {real, imag} */,
  {32'hbd750140, 32'hc15c9497} /* (26, 23, 4) {real, imag} */,
  {32'hc126f7bc, 32'hc11f48f6} /* (26, 23, 3) {real, imag} */,
  {32'hc0bcd8a0, 32'hc0e57b88} /* (26, 23, 2) {real, imag} */,
  {32'h403b2232, 32'hc185ac12} /* (26, 23, 1) {real, imag} */,
  {32'h41370c6a, 32'hc11a627a} /* (26, 23, 0) {real, imag} */,
  {32'h3ff4025a, 32'h4062c7e4} /* (26, 22, 31) {real, imag} */,
  {32'h3f71b21e, 32'h4122b6aa} /* (26, 22, 30) {real, imag} */,
  {32'h3d01e900, 32'h40892f40} /* (26, 22, 29) {real, imag} */,
  {32'hbfe9005e, 32'hc0f09a5a} /* (26, 22, 28) {real, imag} */,
  {32'hbfe1149c, 32'hc030de8b} /* (26, 22, 27) {real, imag} */,
  {32'h40e0572d, 32'h3efff810} /* (26, 22, 26) {real, imag} */,
  {32'h3fba73c4, 32'h3f04a0d6} /* (26, 22, 25) {real, imag} */,
  {32'hc08480bb, 32'h411162f4} /* (26, 22, 24) {real, imag} */,
  {32'hc087c4ec, 32'hbf9ead4e} /* (26, 22, 23) {real, imag} */,
  {32'h40e1604e, 32'h4071e5ce} /* (26, 22, 22) {real, imag} */,
  {32'hc03aeabc, 32'h4101035c} /* (26, 22, 21) {real, imag} */,
  {32'h40fb1c52, 32'h404daf60} /* (26, 22, 20) {real, imag} */,
  {32'h40082dcc, 32'h40ff4134} /* (26, 22, 19) {real, imag} */,
  {32'hc1441bed, 32'h4086cd02} /* (26, 22, 18) {real, imag} */,
  {32'hc01f7d33, 32'h4040d176} /* (26, 22, 17) {real, imag} */,
  {32'h4120948c, 32'h40e4d432} /* (26, 22, 16) {real, imag} */,
  {32'h415fa858, 32'h40f6b610} /* (26, 22, 15) {real, imag} */,
  {32'h40c038ea, 32'h40fa9f66} /* (26, 22, 14) {real, imag} */,
  {32'hc05ad7f6, 32'hbfb99658} /* (26, 22, 13) {real, imag} */,
  {32'hc100531c, 32'h3e0e4a60} /* (26, 22, 12) {real, imag} */,
  {32'hc0428b31, 32'hc0024389} /* (26, 22, 11) {real, imag} */,
  {32'hc0972c24, 32'hc033ae79} /* (26, 22, 10) {real, imag} */,
  {32'hc04fd4df, 32'hbfca6422} /* (26, 22, 9) {real, imag} */,
  {32'h40f2f3aa, 32'h40d4c8bc} /* (26, 22, 8) {real, imag} */,
  {32'h415ef1d2, 32'h40e80591} /* (26, 22, 7) {real, imag} */,
  {32'hc02d1ec1, 32'h3ecc31d0} /* (26, 22, 6) {real, imag} */,
  {32'hc0068be2, 32'h408e7d92} /* (26, 22, 5) {real, imag} */,
  {32'h404d67d1, 32'h3e6ffe80} /* (26, 22, 4) {real, imag} */,
  {32'hbfb4b34e, 32'hc03a8dc9} /* (26, 22, 3) {real, imag} */,
  {32'h3fe5f61e, 32'hc13a31ee} /* (26, 22, 2) {real, imag} */,
  {32'hbf65fbd8, 32'hc108e05e} /* (26, 22, 1) {real, imag} */,
  {32'hc0237bad, 32'hc0c00fc9} /* (26, 22, 0) {real, imag} */,
  {32'h4094a284, 32'h40842ca2} /* (26, 21, 31) {real, imag} */,
  {32'h410fb384, 32'h4023b1e7} /* (26, 21, 30) {real, imag} */,
  {32'h41295d6a, 32'h40c58f2a} /* (26, 21, 29) {real, imag} */,
  {32'h407ff1f8, 32'hbdb0ebd0} /* (26, 21, 28) {real, imag} */,
  {32'hc0179184, 32'hc0c19ae0} /* (26, 21, 27) {real, imag} */,
  {32'h401b122b, 32'h3ff011f2} /* (26, 21, 26) {real, imag} */,
  {32'h41310ad6, 32'hbf87f57a} /* (26, 21, 25) {real, imag} */,
  {32'h404e3266, 32'hc118383c} /* (26, 21, 24) {real, imag} */,
  {32'hc05367f5, 32'hbeb32370} /* (26, 21, 23) {real, imag} */,
  {32'h3d85a740, 32'hc078a4fb} /* (26, 21, 22) {real, imag} */,
  {32'h408f1410, 32'hc083d285} /* (26, 21, 21) {real, imag} */,
  {32'h4052212b, 32'hc0b2c9f1} /* (26, 21, 20) {real, imag} */,
  {32'h402e4386, 32'hc054dfe7} /* (26, 21, 19) {real, imag} */,
  {32'hc0f6e272, 32'hc098025c} /* (26, 21, 18) {real, imag} */,
  {32'hbf0ed96c, 32'h3fde5aea} /* (26, 21, 17) {real, imag} */,
  {32'h4109719e, 32'hc0c4ef7a} /* (26, 21, 16) {real, imag} */,
  {32'h410e5958, 32'hc0d23842} /* (26, 21, 15) {real, imag} */,
  {32'h402a0706, 32'hc11028f6} /* (26, 21, 14) {real, imag} */,
  {32'hc05f8384, 32'h3e7f51b4} /* (26, 21, 13) {real, imag} */,
  {32'h4047b0fe, 32'h40030abc} /* (26, 21, 12) {real, imag} */,
  {32'h4114b344, 32'h4092b708} /* (26, 21, 11) {real, imag} */,
  {32'h40cfca6e, 32'h40f92898} /* (26, 21, 10) {real, imag} */,
  {32'hc0a93215, 32'hc05b4fe0} /* (26, 21, 9) {real, imag} */,
  {32'hc14328e5, 32'hc101beb6} /* (26, 21, 8) {real, imag} */,
  {32'hc1531694, 32'hc0e5eb8c} /* (26, 21, 7) {real, imag} */,
  {32'hc11cc4ac, 32'h3f342520} /* (26, 21, 6) {real, imag} */,
  {32'hbdc72900, 32'h3f809ae8} /* (26, 21, 5) {real, imag} */,
  {32'h404e1e5a, 32'hbea3c530} /* (26, 21, 4) {real, imag} */,
  {32'hbf7b4b94, 32'hc088c4b6} /* (26, 21, 3) {real, imag} */,
  {32'h40490fc4, 32'hbff0f642} /* (26, 21, 2) {real, imag} */,
  {32'hbf289e9e, 32'h401bd9d3} /* (26, 21, 1) {real, imag} */,
  {32'h3e9cb5e0, 32'h3f2417dc} /* (26, 21, 0) {real, imag} */,
  {32'hc1083c03, 32'hbf813ca0} /* (26, 20, 31) {real, imag} */,
  {32'hc0cef22e, 32'h40066ab4} /* (26, 20, 30) {real, imag} */,
  {32'hc07c1cdc, 32'h40eede8c} /* (26, 20, 29) {real, imag} */,
  {32'hc01f5843, 32'h4094cf15} /* (26, 20, 28) {real, imag} */,
  {32'h3f9c9770, 32'hbf36b194} /* (26, 20, 27) {real, imag} */,
  {32'h409333b0, 32'h402d79e8} /* (26, 20, 26) {real, imag} */,
  {32'h403ddc0e, 32'h40491b0b} /* (26, 20, 25) {real, imag} */,
  {32'hc03f63aa, 32'hc05910fe} /* (26, 20, 24) {real, imag} */,
  {32'hc013ff3e, 32'hc08a01f0} /* (26, 20, 23) {real, imag} */,
  {32'hc0c95d21, 32'hc025c470} /* (26, 20, 22) {real, imag} */,
  {32'hc0a57f47, 32'hc0523a9c} /* (26, 20, 21) {real, imag} */,
  {32'h40bccdc1, 32'hbec5d4c8} /* (26, 20, 20) {real, imag} */,
  {32'h407f4a88, 32'hc04450a2} /* (26, 20, 19) {real, imag} */,
  {32'hbf872f6c, 32'hc0936128} /* (26, 20, 18) {real, imag} */,
  {32'hbfec448e, 32'h409ca4b2} /* (26, 20, 17) {real, imag} */,
  {32'hc0938746, 32'h40da526b} /* (26, 20, 16) {real, imag} */,
  {32'hbf912a50, 32'hbfdf3e1c} /* (26, 20, 15) {real, imag} */,
  {32'h403e126e, 32'hc0466dc2} /* (26, 20, 14) {real, imag} */,
  {32'h408f6d7e, 32'hbf83183a} /* (26, 20, 13) {real, imag} */,
  {32'h3f5fc936, 32'h40c92c38} /* (26, 20, 12) {real, imag} */,
  {32'h402bd7a0, 32'h411180ea} /* (26, 20, 11) {real, imag} */,
  {32'h40addc5a, 32'h40b1b322} /* (26, 20, 10) {real, imag} */,
  {32'hbfe70a52, 32'hc0332021} /* (26, 20, 9) {real, imag} */,
  {32'h3eb9e818, 32'hc012373d} /* (26, 20, 8) {real, imag} */,
  {32'h405dc664, 32'hbf180f78} /* (26, 20, 7) {real, imag} */,
  {32'hc056926d, 32'hbda4d1e0} /* (26, 20, 6) {real, imag} */,
  {32'hbf80c494, 32'hc01099bf} /* (26, 20, 5) {real, imag} */,
  {32'hc05a699e, 32'hc05869d8} /* (26, 20, 4) {real, imag} */,
  {32'hc01ba3e8, 32'hbfbe4f5c} /* (26, 20, 3) {real, imag} */,
  {32'hc10f34de, 32'hbf2edd9b} /* (26, 20, 2) {real, imag} */,
  {32'hc0a8fa16, 32'h40a455fb} /* (26, 20, 1) {real, imag} */,
  {32'hbf77ed88, 32'hbf81c8c0} /* (26, 20, 0) {real, imag} */,
  {32'h4014c492, 32'h3f3047d6} /* (26, 19, 31) {real, imag} */,
  {32'h406713bc, 32'hbf978e28} /* (26, 19, 30) {real, imag} */,
  {32'h3fa49bf7, 32'hc008260c} /* (26, 19, 29) {real, imag} */,
  {32'hbf8eaee4, 32'hbfbbf568} /* (26, 19, 28) {real, imag} */,
  {32'hc0404ba8, 32'h40256c43} /* (26, 19, 27) {real, imag} */,
  {32'hc00d5f80, 32'h3e460200} /* (26, 19, 26) {real, imag} */,
  {32'h40aaff0c, 32'hbe90db60} /* (26, 19, 25) {real, imag} */,
  {32'h40cd08ee, 32'h40c18b58} /* (26, 19, 24) {real, imag} */,
  {32'h3fd21f64, 32'hc08ff67d} /* (26, 19, 23) {real, imag} */,
  {32'hbfde9e58, 32'h4019e676} /* (26, 19, 22) {real, imag} */,
  {32'hbe9cf4c0, 32'h3e722d18} /* (26, 19, 21) {real, imag} */,
  {32'h3fd480dd, 32'hc03ed458} /* (26, 19, 20) {real, imag} */,
  {32'hc0559dc0, 32'hbe742508} /* (26, 19, 19) {real, imag} */,
  {32'hc0411f2d, 32'hc0f1791d} /* (26, 19, 18) {real, imag} */,
  {32'hc0c1a548, 32'hc10f6d47} /* (26, 19, 17) {real, imag} */,
  {32'hbf850268, 32'hc10fc8a7} /* (26, 19, 16) {real, imag} */,
  {32'h3ff1b6cc, 32'h3fed0daa} /* (26, 19, 15) {real, imag} */,
  {32'hc01cad28, 32'h40d96b70} /* (26, 19, 14) {real, imag} */,
  {32'hc07d3f1f, 32'h3fe674b8} /* (26, 19, 13) {real, imag} */,
  {32'hc0ce1a7b, 32'hc089cb79} /* (26, 19, 12) {real, imag} */,
  {32'hbfde463e, 32'hc090d042} /* (26, 19, 11) {real, imag} */,
  {32'hc03d5c11, 32'hbf1d9094} /* (26, 19, 10) {real, imag} */,
  {32'h4082d646, 32'hbfe46d80} /* (26, 19, 9) {real, imag} */,
  {32'h3fd90c9a, 32'h403b0216} /* (26, 19, 8) {real, imag} */,
  {32'h4065b9b8, 32'h401fdbb8} /* (26, 19, 7) {real, imag} */,
  {32'h3f8b4a04, 32'h40b49b1a} /* (26, 19, 6) {real, imag} */,
  {32'hc0506412, 32'h40923f5d} /* (26, 19, 5) {real, imag} */,
  {32'h403e6f98, 32'h40a2aa1c} /* (26, 19, 4) {real, imag} */,
  {32'h4075eda6, 32'h404a3ebe} /* (26, 19, 3) {real, imag} */,
  {32'h3ff0df0a, 32'h40c4d681} /* (26, 19, 2) {real, imag} */,
  {32'hc03b7162, 32'h4107e292} /* (26, 19, 1) {real, imag} */,
  {32'hbf9b57e7, 32'h40c90552} /* (26, 19, 0) {real, imag} */,
  {32'h3d8fb830, 32'hbf6cc6d0} /* (26, 18, 31) {real, imag} */,
  {32'hc084a5a0, 32'h3fd11a94} /* (26, 18, 30) {real, imag} */,
  {32'hc06792fa, 32'h40849995} /* (26, 18, 29) {real, imag} */,
  {32'hc022a9f2, 32'h408a04f0} /* (26, 18, 28) {real, imag} */,
  {32'hc07e1fe9, 32'h40412cca} /* (26, 18, 27) {real, imag} */,
  {32'hc0778bd0, 32'hc06a99f4} /* (26, 18, 26) {real, imag} */,
  {32'hc02a1e3e, 32'hbe152c58} /* (26, 18, 25) {real, imag} */,
  {32'h3f2701e4, 32'h40374616} /* (26, 18, 24) {real, imag} */,
  {32'h3f049280, 32'h403a267a} /* (26, 18, 23) {real, imag} */,
  {32'hbf88849d, 32'h4039b83a} /* (26, 18, 22) {real, imag} */,
  {32'hc02fd4bc, 32'hc04c7814} /* (26, 18, 21) {real, imag} */,
  {32'hc0023ab8, 32'hc0d17ba4} /* (26, 18, 20) {real, imag} */,
  {32'h4048a1a3, 32'hbf901d50} /* (26, 18, 19) {real, imag} */,
  {32'h4100f92e, 32'h4009d613} /* (26, 18, 18) {real, imag} */,
  {32'h3ed32b38, 32'hc03dfa1c} /* (26, 18, 17) {real, imag} */,
  {32'hc0402c98, 32'hc097716d} /* (26, 18, 16) {real, imag} */,
  {32'h3e283a20, 32'hc0a49ee7} /* (26, 18, 15) {real, imag} */,
  {32'h3ef11f90, 32'hc0be0b45} /* (26, 18, 14) {real, imag} */,
  {32'h3f579d28, 32'hc00f50d4} /* (26, 18, 13) {real, imag} */,
  {32'hbe143f70, 32'hc00b06ad} /* (26, 18, 12) {real, imag} */,
  {32'h3fcb33a0, 32'h3ea06150} /* (26, 18, 11) {real, imag} */,
  {32'hc00c6d0c, 32'hbef60548} /* (26, 18, 10) {real, imag} */,
  {32'hc081adcc, 32'h3f0e0158} /* (26, 18, 9) {real, imag} */,
  {32'hc0e99b0a, 32'hbee533f8} /* (26, 18, 8) {real, imag} */,
  {32'h3fa34674, 32'h3f1cb564} /* (26, 18, 7) {real, imag} */,
  {32'hbe9ea9d0, 32'hc09f4a32} /* (26, 18, 6) {real, imag} */,
  {32'hc0ca566e, 32'hc09ed998} /* (26, 18, 5) {real, imag} */,
  {32'hc00da226, 32'hbf70bce0} /* (26, 18, 4) {real, imag} */,
  {32'h3e4ff6a8, 32'h3e8efc88} /* (26, 18, 3) {real, imag} */,
  {32'h3f62fb84, 32'h3c8cd2a0} /* (26, 18, 2) {real, imag} */,
  {32'hc094b83f, 32'hc0d2b709} /* (26, 18, 1) {real, imag} */,
  {32'hc0a8aef4, 32'hc0ec117a} /* (26, 18, 0) {real, imag} */,
  {32'h40d863ca, 32'h3fa2eac0} /* (26, 17, 31) {real, imag} */,
  {32'h40927667, 32'hc032d704} /* (26, 17, 30) {real, imag} */,
  {32'h3e968a38, 32'hbf18de6b} /* (26, 17, 29) {real, imag} */,
  {32'h40884a7a, 32'h401ba7ce} /* (26, 17, 28) {real, imag} */,
  {32'h40009c80, 32'h3f0b55fc} /* (26, 17, 27) {real, imag} */,
  {32'hbfd46ce0, 32'hc04d6c8d} /* (26, 17, 26) {real, imag} */,
  {32'hc065ce60, 32'hc0748e69} /* (26, 17, 25) {real, imag} */,
  {32'hbff56a4d, 32'hbfd1dd45} /* (26, 17, 24) {real, imag} */,
  {32'h3f8f256c, 32'hbe3610f8} /* (26, 17, 23) {real, imag} */,
  {32'h410b9856, 32'hc09c03e8} /* (26, 17, 22) {real, imag} */,
  {32'h4060f088, 32'hc06c234e} /* (26, 17, 21) {real, imag} */,
  {32'h400873a8, 32'h3eb5d180} /* (26, 17, 20) {real, imag} */,
  {32'h409b470c, 32'h40d7c0fb} /* (26, 17, 19) {real, imag} */,
  {32'h40793c05, 32'h404ad3b3} /* (26, 17, 18) {real, imag} */,
  {32'h3f32fa08, 32'hc0cca910} /* (26, 17, 17) {real, imag} */,
  {32'h3e87e248, 32'hc10d7b50} /* (26, 17, 16) {real, imag} */,
  {32'hbfae06f4, 32'hc1002488} /* (26, 17, 15) {real, imag} */,
  {32'hbf7e1a88, 32'hc0b3dea7} /* (26, 17, 14) {real, imag} */,
  {32'h40164426, 32'hbf590266} /* (26, 17, 13) {real, imag} */,
  {32'hbe848148, 32'h4052888a} /* (26, 17, 12) {real, imag} */,
  {32'h3f458894, 32'h4031d568} /* (26, 17, 11) {real, imag} */,
  {32'h40da9fe6, 32'hc04213ac} /* (26, 17, 10) {real, imag} */,
  {32'h402e2eba, 32'h4035a472} /* (26, 17, 9) {real, imag} */,
  {32'hbfd1634c, 32'h407c7310} /* (26, 17, 8) {real, imag} */,
  {32'hbfb8e8b4, 32'hbdc51e20} /* (26, 17, 7) {real, imag} */,
  {32'h40357d70, 32'hbd7b2200} /* (26, 17, 6) {real, imag} */,
  {32'h3fdfd2e6, 32'h4030937c} /* (26, 17, 5) {real, imag} */,
  {32'hc003a079, 32'h4057e45c} /* (26, 17, 4) {real, imag} */,
  {32'h3f84df68, 32'hc00677d9} /* (26, 17, 3) {real, imag} */,
  {32'h4075d6b3, 32'hbeefede8} /* (26, 17, 2) {real, imag} */,
  {32'h3fa34d33, 32'h3f9ecdcc} /* (26, 17, 1) {real, imag} */,
  {32'h3e75e5e0, 32'h4012426d} /* (26, 17, 0) {real, imag} */,
  {32'hbf8b1097, 32'hc048120a} /* (26, 16, 31) {real, imag} */,
  {32'h406256c2, 32'hbdd17380} /* (26, 16, 30) {real, imag} */,
  {32'h401562ca, 32'hbfcd0f74} /* (26, 16, 29) {real, imag} */,
  {32'h3ff68010, 32'h3f57c750} /* (26, 16, 28) {real, imag} */,
  {32'hbd35b800, 32'hbcf70600} /* (26, 16, 27) {real, imag} */,
  {32'hc05b82c4, 32'hbd0ddb60} /* (26, 16, 26) {real, imag} */,
  {32'hc081def7, 32'h3fe023c5} /* (26, 16, 25) {real, imag} */,
  {32'h3f19c778, 32'hbe5d1bd0} /* (26, 16, 24) {real, imag} */,
  {32'h4066d5a6, 32'h3eba8770} /* (26, 16, 23) {real, imag} */,
  {32'h3d19fe60, 32'h3f7047e0} /* (26, 16, 22) {real, imag} */,
  {32'hbf79211c, 32'hc040806e} /* (26, 16, 21) {real, imag} */,
  {32'hbd142540, 32'hbe6661a0} /* (26, 16, 20) {real, imag} */,
  {32'hbf6338c4, 32'hbed202a0} /* (26, 16, 19) {real, imag} */,
  {32'h3f4281fd, 32'hc0073d64} /* (26, 16, 18) {real, imag} */,
  {32'h3f371d90, 32'hc031e2a7} /* (26, 16, 17) {real, imag} */,
  {32'hbfc9f872, 32'hbe812fac} /* (26, 16, 16) {real, imag} */,
  {32'hc03b2f72, 32'hc08ef44a} /* (26, 16, 15) {real, imag} */,
  {32'hbfc818b8, 32'hc01bf9c4} /* (26, 16, 14) {real, imag} */,
  {32'h405789c0, 32'hbff63d5a} /* (26, 16, 13) {real, imag} */,
  {32'h40944284, 32'hbf2ff2e0} /* (26, 16, 12) {real, imag} */,
  {32'h4076490e, 32'hbf9b1910} /* (26, 16, 11) {real, imag} */,
  {32'h3fcc7a9c, 32'hbe6f1c60} /* (26, 16, 10) {real, imag} */,
  {32'hc008a576, 32'h40786ab8} /* (26, 16, 9) {real, imag} */,
  {32'hc07a3450, 32'hbe71ec00} /* (26, 16, 8) {real, imag} */,
  {32'hbf9eea10, 32'h3f37fd78} /* (26, 16, 7) {real, imag} */,
  {32'hc01a4efa, 32'hbf79c0c0} /* (26, 16, 6) {real, imag} */,
  {32'h3f9e1557, 32'h3fc1a828} /* (26, 16, 5) {real, imag} */,
  {32'h4014b88c, 32'h403cf568} /* (26, 16, 4) {real, imag} */,
  {32'h405e15e3, 32'h3f6b6c30} /* (26, 16, 3) {real, imag} */,
  {32'h3fe21216, 32'h3f5d5240} /* (26, 16, 2) {real, imag} */,
  {32'hbf8952d8, 32'h3feabc80} /* (26, 16, 1) {real, imag} */,
  {32'h3f9d4050, 32'h3f782f18} /* (26, 16, 0) {real, imag} */,
  {32'hc04505b9, 32'hc08cf9d6} /* (26, 15, 31) {real, imag} */,
  {32'h400159b2, 32'hbfe5bb6f} /* (26, 15, 30) {real, imag} */,
  {32'h3f8af4da, 32'hbfda012e} /* (26, 15, 29) {real, imag} */,
  {32'hc05fdf71, 32'hc0b0aeaf} /* (26, 15, 28) {real, imag} */,
  {32'hc08c0a54, 32'hc0944cca} /* (26, 15, 27) {real, imag} */,
  {32'hc00420c0, 32'hc02fa39d} /* (26, 15, 26) {real, imag} */,
  {32'h3e51e400, 32'h3fbadd26} /* (26, 15, 25) {real, imag} */,
  {32'hbe968d34, 32'hbfb253ef} /* (26, 15, 24) {real, imag} */,
  {32'hbf99f308, 32'hbf652222} /* (26, 15, 23) {real, imag} */,
  {32'hc06a901e, 32'h402fb6a5} /* (26, 15, 22) {real, imag} */,
  {32'h4080fc16, 32'h408e2d65} /* (26, 15, 21) {real, imag} */,
  {32'hc00e91e8, 32'h41029d14} /* (26, 15, 20) {real, imag} */,
  {32'hbe5e6fd0, 32'h40c7e191} /* (26, 15, 19) {real, imag} */,
  {32'h3f832fc6, 32'hc00d418d} /* (26, 15, 18) {real, imag} */,
  {32'h3f169058, 32'hbeece300} /* (26, 15, 17) {real, imag} */,
  {32'hc050b9cf, 32'hbee40e50} /* (26, 15, 16) {real, imag} */,
  {32'hc058768e, 32'h3dc52440} /* (26, 15, 15) {real, imag} */,
  {32'hc0484796, 32'hc03f3182} /* (26, 15, 14) {real, imag} */,
  {32'hc07efbee, 32'hc0371dca} /* (26, 15, 13) {real, imag} */,
  {32'hc0a9f664, 32'hc09edb83} /* (26, 15, 12) {real, imag} */,
  {32'hbf59fc54, 32'hc09e9c3c} /* (26, 15, 11) {real, imag} */,
  {32'h3ec81048, 32'hc039477a} /* (26, 15, 10) {real, imag} */,
  {32'h404399fa, 32'hc03e592a} /* (26, 15, 9) {real, imag} */,
  {32'h401e7d8a, 32'h4051a8a4} /* (26, 15, 8) {real, imag} */,
  {32'hbe7c9020, 32'h40eae460} /* (26, 15, 7) {real, imag} */,
  {32'hc0be8800, 32'h41169a8c} /* (26, 15, 6) {real, imag} */,
  {32'hbf39315c, 32'h4101f266} /* (26, 15, 5) {real, imag} */,
  {32'h3fa9358a, 32'h40c6e7e0} /* (26, 15, 4) {real, imag} */,
  {32'hbda88618, 32'h3f201214} /* (26, 15, 3) {real, imag} */,
  {32'hbf4cd41c, 32'hbfc9809e} /* (26, 15, 2) {real, imag} */,
  {32'hbf67744e, 32'hbffa0274} /* (26, 15, 1) {real, imag} */,
  {32'hc0ac2a17, 32'hc02183d3} /* (26, 15, 0) {real, imag} */,
  {32'h3f78d6c2, 32'h3fa5d448} /* (26, 14, 31) {real, imag} */,
  {32'hc0a2b49c, 32'h403a686e} /* (26, 14, 30) {real, imag} */,
  {32'hc09ceafd, 32'hbe323eb8} /* (26, 14, 29) {real, imag} */,
  {32'hbfe0f83d, 32'hc042939c} /* (26, 14, 28) {real, imag} */,
  {32'h40700129, 32'h40823bfd} /* (26, 14, 27) {real, imag} */,
  {32'h3f73ef70, 32'h409216fe} /* (26, 14, 26) {real, imag} */,
  {32'h3fdbe9a4, 32'h403521ce} /* (26, 14, 25) {real, imag} */,
  {32'h40846766, 32'h3ffd9855} /* (26, 14, 24) {real, imag} */,
  {32'h404c9b56, 32'hbf5890a8} /* (26, 14, 23) {real, imag} */,
  {32'h40623f2a, 32'h40267f54} /* (26, 14, 22) {real, imag} */,
  {32'h4050fe30, 32'h406e7bcc} /* (26, 14, 21) {real, imag} */,
  {32'h40998fb2, 32'h40bc31c8} /* (26, 14, 20) {real, imag} */,
  {32'h3ff279b6, 32'h3e2efb80} /* (26, 14, 19) {real, imag} */,
  {32'hbfb0cb0c, 32'hbf16fb1c} /* (26, 14, 18) {real, imag} */,
  {32'hc0bff288, 32'h3ffeaba4} /* (26, 14, 17) {real, imag} */,
  {32'hc076a5cc, 32'hbe5a8e60} /* (26, 14, 16) {real, imag} */,
  {32'h3f872b5c, 32'hbf70e108} /* (26, 14, 15) {real, imag} */,
  {32'h4017c486, 32'h3eff7990} /* (26, 14, 14) {real, imag} */,
  {32'h409ffb0b, 32'h40098020} /* (26, 14, 13) {real, imag} */,
  {32'h40bacfc2, 32'hc05cee25} /* (26, 14, 12) {real, imag} */,
  {32'h3fa865f0, 32'h3fb82c90} /* (26, 14, 11) {real, imag} */,
  {32'h4005d51c, 32'h402ab9f9} /* (26, 14, 10) {real, imag} */,
  {32'h3e24bcf0, 32'hbf0f3c08} /* (26, 14, 9) {real, imag} */,
  {32'hc0f8acec, 32'hbfa5ef4e} /* (26, 14, 8) {real, imag} */,
  {32'hc1345e90, 32'hc08c9ed4} /* (26, 14, 7) {real, imag} */,
  {32'hc09fd25c, 32'hc0906e7c} /* (26, 14, 6) {real, imag} */,
  {32'h40048064, 32'hbf1fdc50} /* (26, 14, 5) {real, imag} */,
  {32'h4046aec2, 32'h3fabe0a4} /* (26, 14, 4) {real, imag} */,
  {32'h40560768, 32'h40312f0b} /* (26, 14, 3) {real, imag} */,
  {32'h3fc367f6, 32'h3ff41b66} /* (26, 14, 2) {real, imag} */,
  {32'hc0309372, 32'hc090d05d} /* (26, 14, 1) {real, imag} */,
  {32'hc0812158, 32'hc08dcc7a} /* (26, 14, 0) {real, imag} */,
  {32'hc0087642, 32'h40091b7e} /* (26, 13, 31) {real, imag} */,
  {32'hbfa3a790, 32'h3fe7f348} /* (26, 13, 30) {real, imag} */,
  {32'h402c8080, 32'hc0852c2a} /* (26, 13, 29) {real, imag} */,
  {32'h400a9a8e, 32'hbf067b78} /* (26, 13, 28) {real, imag} */,
  {32'hc0874711, 32'hbecd48f8} /* (26, 13, 27) {real, imag} */,
  {32'h40113fc8, 32'hc0130db8} /* (26, 13, 26) {real, imag} */,
  {32'h3d423a40, 32'h4084d7f4} /* (26, 13, 25) {real, imag} */,
  {32'hc0488a75, 32'h40acbeac} /* (26, 13, 24) {real, imag} */,
  {32'hc0a29a4f, 32'hbe399160} /* (26, 13, 23) {real, imag} */,
  {32'hc0f1fd00, 32'h3fc468b6} /* (26, 13, 22) {real, imag} */,
  {32'hc0be6230, 32'hbb3d5a00} /* (26, 13, 21) {real, imag} */,
  {32'h3eda9f34, 32'hbfa61f48} /* (26, 13, 20) {real, imag} */,
  {32'h3e8d42c0, 32'hbf21f8aa} /* (26, 13, 19) {real, imag} */,
  {32'hc06d1bcb, 32'h4094df95} /* (26, 13, 18) {real, imag} */,
  {32'h3f8d90d8, 32'h40da607a} /* (26, 13, 17) {real, imag} */,
  {32'h403c2664, 32'h404521a4} /* (26, 13, 16) {real, imag} */,
  {32'h405392d2, 32'h3fc3252e} /* (26, 13, 15) {real, imag} */,
  {32'h409c2f93, 32'h4078f8bc} /* (26, 13, 14) {real, imag} */,
  {32'h4073bc97, 32'h40ce5d64} /* (26, 13, 13) {real, imag} */,
  {32'h40d18571, 32'h3f93e764} /* (26, 13, 12) {real, imag} */,
  {32'h402ce291, 32'hbfccbf98} /* (26, 13, 11) {real, imag} */,
  {32'hbf8f245e, 32'hbecd7d78} /* (26, 13, 10) {real, imag} */,
  {32'hc08119da, 32'h404055e0} /* (26, 13, 9) {real, imag} */,
  {32'h400e4aeb, 32'h3f7c5996} /* (26, 13, 8) {real, imag} */,
  {32'h40be035a, 32'h3f4414e0} /* (26, 13, 7) {real, imag} */,
  {32'hc056cee4, 32'h3fcc15c0} /* (26, 13, 6) {real, imag} */,
  {32'hc02c82d6, 32'hbec5f1f0} /* (26, 13, 5) {real, imag} */,
  {32'h3e358d38, 32'hc091466e} /* (26, 13, 4) {real, imag} */,
  {32'h400be6fc, 32'h3fdfaedc} /* (26, 13, 3) {real, imag} */,
  {32'hbf0c2d34, 32'hc055362e} /* (26, 13, 2) {real, imag} */,
  {32'hc02105c2, 32'hc07f68e8} /* (26, 13, 1) {real, imag} */,
  {32'hc087513e, 32'h400f9fad} /* (26, 13, 0) {real, imag} */,
  {32'hbddc9880, 32'hc0a8a5e7} /* (26, 12, 31) {real, imag} */,
  {32'h400032c5, 32'hc122c306} /* (26, 12, 30) {real, imag} */,
  {32'h4099b50c, 32'h3f47db20} /* (26, 12, 29) {real, imag} */,
  {32'h400d8269, 32'h3fa93dcb} /* (26, 12, 28) {real, imag} */,
  {32'hbfa4b3f8, 32'h3d2780c0} /* (26, 12, 27) {real, imag} */,
  {32'hc0a55228, 32'hc0147cbc} /* (26, 12, 26) {real, imag} */,
  {32'hc0ff89f3, 32'h4085d484} /* (26, 12, 25) {real, imag} */,
  {32'hc13422e4, 32'h40550b5c} /* (26, 12, 24) {real, imag} */,
  {32'hc0340c6e, 32'h3f51841c} /* (26, 12, 23) {real, imag} */,
  {32'h3f1b8b38, 32'h405d6518} /* (26, 12, 22) {real, imag} */,
  {32'hbfe6b13c, 32'h3eade120} /* (26, 12, 21) {real, imag} */,
  {32'h408cca17, 32'h40289da3} /* (26, 12, 20) {real, imag} */,
  {32'h4127efe7, 32'h3f48ea58} /* (26, 12, 19) {real, imag} */,
  {32'hbf2195d8, 32'hc0c2c334} /* (26, 12, 18) {real, imag} */,
  {32'hbed88938, 32'h405c46cc} /* (26, 12, 17) {real, imag} */,
  {32'h40606935, 32'hc0359512} /* (26, 12, 16) {real, imag} */,
  {32'h411f93a2, 32'hc1231352} /* (26, 12, 15) {real, imag} */,
  {32'h40bfab77, 32'hc06a2550} /* (26, 12, 14) {real, imag} */,
  {32'hc0063ea5, 32'h3ffdb7ea} /* (26, 12, 13) {real, imag} */,
  {32'hc00785be, 32'hbf5435b0} /* (26, 12, 12) {real, imag} */,
  {32'hc0442258, 32'hc08931ca} /* (26, 12, 11) {real, imag} */,
  {32'hc029cc9f, 32'hc043df0b} /* (26, 12, 10) {real, imag} */,
  {32'hbfc53cfe, 32'hbf9c2c9e} /* (26, 12, 9) {real, imag} */,
  {32'h405c995f, 32'hbfac337e} /* (26, 12, 8) {real, imag} */,
  {32'h404924e4, 32'hc05de26e} /* (26, 12, 7) {real, imag} */,
  {32'h4015632f, 32'hbf458f04} /* (26, 12, 6) {real, imag} */,
  {32'h3faf17bc, 32'hbfb41a6a} /* (26, 12, 5) {real, imag} */,
  {32'h3e773aa0, 32'hc0365390} /* (26, 12, 4) {real, imag} */,
  {32'h408b2edc, 32'h3fbece8c} /* (26, 12, 3) {real, imag} */,
  {32'h3f778700, 32'hbfee7f52} /* (26, 12, 2) {real, imag} */,
  {32'hc063a444, 32'h3fcb9fbc} /* (26, 12, 1) {real, imag} */,
  {32'h3e082860, 32'hc00378f8} /* (26, 12, 0) {real, imag} */,
  {32'h3f097fd4, 32'h3f80c891} /* (26, 11, 31) {real, imag} */,
  {32'hbeb93150, 32'hbf5feae4} /* (26, 11, 30) {real, imag} */,
  {32'h3fdc80c0, 32'h4001d3a3} /* (26, 11, 29) {real, imag} */,
  {32'h40e30b04, 32'hbe3a7dc8} /* (26, 11, 28) {real, imag} */,
  {32'hc0333380, 32'h3d00cac0} /* (26, 11, 27) {real, imag} */,
  {32'hc1269cda, 32'hc0e96288} /* (26, 11, 26) {real, imag} */,
  {32'hbfaefe04, 32'hbf38e94b} /* (26, 11, 25) {real, imag} */,
  {32'h40febac9, 32'hbf617420} /* (26, 11, 24) {real, imag} */,
  {32'h4013d6bd, 32'hc13a9498} /* (26, 11, 23) {real, imag} */,
  {32'hc091d7b3, 32'hc0a86e37} /* (26, 11, 22) {real, imag} */,
  {32'hc0142978, 32'hc1055eaa} /* (26, 11, 21) {real, imag} */,
  {32'h40929522, 32'hc0906de3} /* (26, 11, 20) {real, imag} */,
  {32'h3f78ffde, 32'h40807dc6} /* (26, 11, 19) {real, imag} */,
  {32'h3f1c6274, 32'h3fdb4e02} /* (26, 11, 18) {real, imag} */,
  {32'h40a09d80, 32'h402bf4cb} /* (26, 11, 17) {real, imag} */,
  {32'h40c6d044, 32'h40be9b5a} /* (26, 11, 16) {real, imag} */,
  {32'h40bfe958, 32'h40b1faa2} /* (26, 11, 15) {real, imag} */,
  {32'h40af0c01, 32'h40bfe527} /* (26, 11, 14) {real, imag} */,
  {32'h407b8a90, 32'hc0013329} /* (26, 11, 13) {real, imag} */,
  {32'hbfd56723, 32'h3d4451a0} /* (26, 11, 12) {real, imag} */,
  {32'h401dc84a, 32'h3f263a64} /* (26, 11, 11) {real, imag} */,
  {32'h3fcb9020, 32'h41299124} /* (26, 11, 10) {real, imag} */,
  {32'hc03d4e06, 32'h40f9496c} /* (26, 11, 9) {real, imag} */,
  {32'hc09cb136, 32'h416357f6} /* (26, 11, 8) {real, imag} */,
  {32'h4092cc3f, 32'h40cfd8a0} /* (26, 11, 7) {real, imag} */,
  {32'h3e2cc120, 32'hc073f5dc} /* (26, 11, 6) {real, imag} */,
  {32'hc0880d3e, 32'hc0a4fbce} /* (26, 11, 5) {real, imag} */,
  {32'h407def1a, 32'hc10c740e} /* (26, 11, 4) {real, imag} */,
  {32'h40cafd96, 32'hc0a2ed94} /* (26, 11, 3) {real, imag} */,
  {32'h4082c50a, 32'hc06fbeb3} /* (26, 11, 2) {real, imag} */,
  {32'hbf3318fa, 32'h3f5f1e6c} /* (26, 11, 1) {real, imag} */,
  {32'hc0a30ada, 32'h40b77dd4} /* (26, 11, 0) {real, imag} */,
  {32'h3f4e30cc, 32'hc0252a54} /* (26, 10, 31) {real, imag} */,
  {32'hc0303d16, 32'hc09df6f2} /* (26, 10, 30) {real, imag} */,
  {32'hc0959306, 32'hc06d8a13} /* (26, 10, 29) {real, imag} */,
  {32'h402e92c5, 32'h40ba5bda} /* (26, 10, 28) {real, imag} */,
  {32'hc1348eb0, 32'h40b97e2e} /* (26, 10, 27) {real, imag} */,
  {32'hc11ecf50, 32'hbfa87c48} /* (26, 10, 26) {real, imag} */,
  {32'hbfb0ee44, 32'hc05ea486} /* (26, 10, 25) {real, imag} */,
  {32'h4106dda0, 32'h3f3e8c98} /* (26, 10, 24) {real, imag} */,
  {32'h3e2d89b0, 32'h408aa3e6} /* (26, 10, 23) {real, imag} */,
  {32'h4116eda9, 32'h40e54ac5} /* (26, 10, 22) {real, imag} */,
  {32'h41555e69, 32'h409abaf6} /* (26, 10, 21) {real, imag} */,
  {32'hbf9f6430, 32'hc0a75678} /* (26, 10, 20) {real, imag} */,
  {32'hc13cbdf1, 32'hc08c2d46} /* (26, 10, 19) {real, imag} */,
  {32'hc0eb221a, 32'hbf0621bc} /* (26, 10, 18) {real, imag} */,
  {32'hc08b34e8, 32'h40ccc949} /* (26, 10, 17) {real, imag} */,
  {32'h3f0f69a8, 32'h40c41782} /* (26, 10, 16) {real, imag} */,
  {32'hc166cfb8, 32'h4105e684} /* (26, 10, 15) {real, imag} */,
  {32'hc13666ef, 32'hc0432518} /* (26, 10, 14) {real, imag} */,
  {32'h407c594e, 32'hc0dda910} /* (26, 10, 13) {real, imag} */,
  {32'h41440804, 32'hc097e97f} /* (26, 10, 12) {real, imag} */,
  {32'h40802cc0, 32'h4099dfbc} /* (26, 10, 11) {real, imag} */,
  {32'hc0b31ce8, 32'h407accdb} /* (26, 10, 10) {real, imag} */,
  {32'hc02f595b, 32'hbf47c8fc} /* (26, 10, 9) {real, imag} */,
  {32'hc0334bfc, 32'h3fdaba72} /* (26, 10, 8) {real, imag} */,
  {32'hc0c52ee8, 32'h40ec4683} /* (26, 10, 7) {real, imag} */,
  {32'hc08c5318, 32'h411580f2} /* (26, 10, 6) {real, imag} */,
  {32'h3fbf3b04, 32'h400e98e7} /* (26, 10, 5) {real, imag} */,
  {32'hc0463cc3, 32'hc087ee8a} /* (26, 10, 4) {real, imag} */,
  {32'hc0e03b06, 32'hbfadf256} /* (26, 10, 3) {real, imag} */,
  {32'hc1049921, 32'h408ccbb0} /* (26, 10, 2) {real, imag} */,
  {32'hc03a6fb2, 32'hbf4c85dc} /* (26, 10, 1) {real, imag} */,
  {32'h4090d19e, 32'hbfce1c7c} /* (26, 10, 0) {real, imag} */,
  {32'h40ebe684, 32'hc096f642} /* (26, 9, 31) {real, imag} */,
  {32'h40c59f5e, 32'h4045203c} /* (26, 9, 30) {real, imag} */,
  {32'h40b61b00, 32'h401a40c8} /* (26, 9, 29) {real, imag} */,
  {32'hc039ce7c, 32'h40271a46} /* (26, 9, 28) {real, imag} */,
  {32'h3e5e3700, 32'hc1002da4} /* (26, 9, 27) {real, imag} */,
  {32'h3faaf062, 32'hbf2fc118} /* (26, 9, 26) {real, imag} */,
  {32'hc104f668, 32'h40be0926} /* (26, 9, 25) {real, imag} */,
  {32'hc0b30193, 32'h3fff6318} /* (26, 9, 24) {real, imag} */,
  {32'h410ed7f7, 32'hc0b0ef3b} /* (26, 9, 23) {real, imag} */,
  {32'h40c7fe6d, 32'hc03fe23a} /* (26, 9, 22) {real, imag} */,
  {32'h407b2d94, 32'hbfcd1db9} /* (26, 9, 21) {real, imag} */,
  {32'hbf9f28e4, 32'hc06e92d6} /* (26, 9, 20) {real, imag} */,
  {32'h410069a4, 32'h4103ed56} /* (26, 9, 19) {real, imag} */,
  {32'h4114f3dd, 32'h40f96d7b} /* (26, 9, 18) {real, imag} */,
  {32'h41073392, 32'h3e8ca320} /* (26, 9, 17) {real, imag} */,
  {32'hc0c1e945, 32'h41487d5e} /* (26, 9, 16) {real, imag} */,
  {32'hc1150466, 32'h40f45c47} /* (26, 9, 15) {real, imag} */,
  {32'h402f7a38, 32'hbe10eb10} /* (26, 9, 14) {real, imag} */,
  {32'hc02fd9ac, 32'hbfbcb6dc} /* (26, 9, 13) {real, imag} */,
  {32'h3f9fd564, 32'h3d94fdc0} /* (26, 9, 12) {real, imag} */,
  {32'h40a003bc, 32'hbfdb33bc} /* (26, 9, 11) {real, imag} */,
  {32'hbfb4d5f8, 32'h3feb26dd} /* (26, 9, 10) {real, imag} */,
  {32'hc105bbc0, 32'hc0aa4976} /* (26, 9, 9) {real, imag} */,
  {32'hc080a0dc, 32'hbe40d690} /* (26, 9, 8) {real, imag} */,
  {32'h410bc071, 32'hc09a5a82} /* (26, 9, 7) {real, imag} */,
  {32'h4009aeb8, 32'hc110a784} /* (26, 9, 6) {real, imag} */,
  {32'h40b528ac, 32'h4097777e} /* (26, 9, 5) {real, imag} */,
  {32'h403dbe17, 32'h410bae2d} /* (26, 9, 4) {real, imag} */,
  {32'h3ed9bf50, 32'h40bb0fec} /* (26, 9, 3) {real, imag} */,
  {32'hc1169b5a, 32'h4153501c} /* (26, 9, 2) {real, imag} */,
  {32'h40e2500f, 32'h40bac326} /* (26, 9, 1) {real, imag} */,
  {32'h410b8624, 32'h3f661a48} /* (26, 9, 0) {real, imag} */,
  {32'h408135a8, 32'hc11c83e0} /* (26, 8, 31) {real, imag} */,
  {32'h402e4563, 32'hc13f180e} /* (26, 8, 30) {real, imag} */,
  {32'h41321550, 32'h404e4071} /* (26, 8, 29) {real, imag} */,
  {32'h418c0d18, 32'hc104f3c7} /* (26, 8, 28) {real, imag} */,
  {32'h40c5340a, 32'hc1868328} /* (26, 8, 27) {real, imag} */,
  {32'hc01584f8, 32'hc0e998af} /* (26, 8, 26) {real, imag} */,
  {32'h41166bf3, 32'hc0832ac0} /* (26, 8, 25) {real, imag} */,
  {32'h408d69e1, 32'hc0a32d80} /* (26, 8, 24) {real, imag} */,
  {32'h40f9b8f2, 32'h408fd5e9} /* (26, 8, 23) {real, imag} */,
  {32'h40925626, 32'h409e457e} /* (26, 8, 22) {real, imag} */,
  {32'hc0865e46, 32'h41a3eb6d} /* (26, 8, 21) {real, imag} */,
  {32'hc1c80861, 32'h402c2c7a} /* (26, 8, 20) {real, imag} */,
  {32'hc0d56a7a, 32'h407edc4c} /* (26, 8, 19) {real, imag} */,
  {32'h409bedae, 32'h40e71f0c} /* (26, 8, 18) {real, imag} */,
  {32'hc02e8b92, 32'hbe5966f0} /* (26, 8, 17) {real, imag} */,
  {32'h40a4eb5a, 32'hc02559f0} /* (26, 8, 16) {real, imag} */,
  {32'h411681b3, 32'hc0e34396} /* (26, 8, 15) {real, imag} */,
  {32'h419f2358, 32'hc1225ec9} /* (26, 8, 14) {real, imag} */,
  {32'h4191f5fc, 32'hc1359561} /* (26, 8, 13) {real, imag} */,
  {32'h4120499e, 32'hbec53cd0} /* (26, 8, 12) {real, imag} */,
  {32'h4116f0a9, 32'h40a12d3d} /* (26, 8, 11) {real, imag} */,
  {32'h4169551a, 32'hbf7de650} /* (26, 8, 10) {real, imag} */,
  {32'h4169c8c0, 32'hbef89e78} /* (26, 8, 9) {real, imag} */,
  {32'h40f828dc, 32'hc148ebf0} /* (26, 8, 8) {real, imag} */,
  {32'h40813cec, 32'hc0e586cd} /* (26, 8, 7) {real, imag} */,
  {32'h3fb63820, 32'h40392278} /* (26, 8, 6) {real, imag} */,
  {32'hc0aa6147, 32'h40921ed7} /* (26, 8, 5) {real, imag} */,
  {32'hc13d5136, 32'hc0a3db8f} /* (26, 8, 4) {real, imag} */,
  {32'hc12f6125, 32'hbfddd158} /* (26, 8, 3) {real, imag} */,
  {32'hc0e4000d, 32'h40d85344} /* (26, 8, 2) {real, imag} */,
  {32'hc041d274, 32'h411c1d8d} /* (26, 8, 1) {real, imag} */,
  {32'h3f3632c8, 32'h411d2a28} /* (26, 8, 0) {real, imag} */,
  {32'hc017e082, 32'h3f3d5284} /* (26, 7, 31) {real, imag} */,
  {32'hc01ca7eb, 32'h405a3dd7} /* (26, 7, 30) {real, imag} */,
  {32'hc0115609, 32'h401431fd} /* (26, 7, 29) {real, imag} */,
  {32'hc1600dd0, 32'h40eb7f71} /* (26, 7, 28) {real, imag} */,
  {32'h40184380, 32'h4159cd0a} /* (26, 7, 27) {real, imag} */,
  {32'h40cc580f, 32'h411348ed} /* (26, 7, 26) {real, imag} */,
  {32'h4134c2da, 32'h410d74bb} /* (26, 7, 25) {real, imag} */,
  {32'h4077d78f, 32'hc003e762} /* (26, 7, 24) {real, imag} */,
  {32'h3faee58c, 32'hc0366492} /* (26, 7, 23) {real, imag} */,
  {32'hc093b6c0, 32'h3f1c6330} /* (26, 7, 22) {real, imag} */,
  {32'h3d797000, 32'h4027453c} /* (26, 7, 21) {real, imag} */,
  {32'hc1367e0f, 32'hc1386ee4} /* (26, 7, 20) {real, imag} */,
  {32'hc157250f, 32'hc13bc0ab} /* (26, 7, 19) {real, imag} */,
  {32'h3f9ac7af, 32'hc005b41c} /* (26, 7, 18) {real, imag} */,
  {32'hc0c690db, 32'h4163c8e6} /* (26, 7, 17) {real, imag} */,
  {32'hc1a50d35, 32'h3fc0d390} /* (26, 7, 16) {real, imag} */,
  {32'hc0f98d50, 32'hc0050276} /* (26, 7, 15) {real, imag} */,
  {32'hc0c80056, 32'hc0acb9da} /* (26, 7, 14) {real, imag} */,
  {32'h4087af16, 32'hc14503a0} /* (26, 7, 13) {real, imag} */,
  {32'h404fd7aa, 32'hc1074f2c} /* (26, 7, 12) {real, imag} */,
  {32'hc097f1bd, 32'hc097c083} /* (26, 7, 11) {real, imag} */,
  {32'hc0cd0b96, 32'h40367316} /* (26, 7, 10) {real, imag} */,
  {32'hbf1288b0, 32'h412f31f7} /* (26, 7, 9) {real, imag} */,
  {32'hc099f1bb, 32'h3fa8c2d8} /* (26, 7, 8) {real, imag} */,
  {32'hc177b182, 32'hc064f110} /* (26, 7, 7) {real, imag} */,
  {32'h403df950, 32'h40f7380b} /* (26, 7, 6) {real, imag} */,
  {32'h3fc8f348, 32'h4182634f} /* (26, 7, 5) {real, imag} */,
  {32'h415d26ec, 32'h40cf2b81} /* (26, 7, 4) {real, imag} */,
  {32'h4147ab39, 32'h41058f5d} /* (26, 7, 3) {real, imag} */,
  {32'h4113b8b9, 32'h412cc460} /* (26, 7, 2) {real, imag} */,
  {32'h40c9f12f, 32'h41273ed3} /* (26, 7, 1) {real, imag} */,
  {32'hc06eccbc, 32'h4109b830} /* (26, 7, 0) {real, imag} */,
  {32'h40a42601, 32'hbfd02962} /* (26, 6, 31) {real, imag} */,
  {32'h411446c5, 32'h40c68864} /* (26, 6, 30) {real, imag} */,
  {32'h401ba4a2, 32'h40e5653c} /* (26, 6, 29) {real, imag} */,
  {32'h3fc688ec, 32'hbf962470} /* (26, 6, 28) {real, imag} */,
  {32'hc11ab2e6, 32'hc1181b7d} /* (26, 6, 27) {real, imag} */,
  {32'h4011068f, 32'hc0d59833} /* (26, 6, 26) {real, imag} */,
  {32'h40f210ff, 32'hc0f98a3f} /* (26, 6, 25) {real, imag} */,
  {32'h410a20be, 32'hc0f3a0a9} /* (26, 6, 24) {real, imag} */,
  {32'h412be26e, 32'hc069083f} /* (26, 6, 23) {real, imag} */,
  {32'h412b183e, 32'hc158067c} /* (26, 6, 22) {real, imag} */,
  {32'h418c07e6, 32'hc18bf0ef} /* (26, 6, 21) {real, imag} */,
  {32'h3ff45b8c, 32'hc103a24e} /* (26, 6, 20) {real, imag} */,
  {32'hc19ec9a6, 32'h410e5b79} /* (26, 6, 19) {real, imag} */,
  {32'hc135e110, 32'h40ad9789} /* (26, 6, 18) {real, imag} */,
  {32'hc19e2ef0, 32'hc150d056} /* (26, 6, 17) {real, imag} */,
  {32'hc13077e0, 32'hc1375a5e} /* (26, 6, 16) {real, imag} */,
  {32'hc0740e2d, 32'hc14e54e5} /* (26, 6, 15) {real, imag} */,
  {32'h40ae15d3, 32'hc05fec1e} /* (26, 6, 14) {real, imag} */,
  {32'hc052e7c4, 32'hc14d9a4c} /* (26, 6, 13) {real, imag} */,
  {32'hc0dddac2, 32'hc1c24292} /* (26, 6, 12) {real, imag} */,
  {32'h40caff84, 32'hc179bcad} /* (26, 6, 11) {real, imag} */,
  {32'hc0184afc, 32'hc0963d32} /* (26, 6, 10) {real, imag} */,
  {32'hc0f6ba68, 32'h40eff284} /* (26, 6, 9) {real, imag} */,
  {32'hbf17c53c, 32'h3fa19fc0} /* (26, 6, 8) {real, imag} */,
  {32'hc0d5d6d4, 32'hc0ce029a} /* (26, 6, 7) {real, imag} */,
  {32'h4126538c, 32'h40e75831} /* (26, 6, 6) {real, imag} */,
  {32'h41895b51, 32'h417ef97b} /* (26, 6, 5) {real, imag} */,
  {32'h3d3dbce0, 32'h3f5e2cfa} /* (26, 6, 4) {real, imag} */,
  {32'hc11f0f6d, 32'hc10d479b} /* (26, 6, 3) {real, imag} */,
  {32'hc0983b7e, 32'hc11954c0} /* (26, 6, 2) {real, imag} */,
  {32'h417c324c, 32'hc0f1c73c} /* (26, 6, 1) {real, imag} */,
  {32'h413c8bcf, 32'hc0f50c6e} /* (26, 6, 0) {real, imag} */,
  {32'hc129723d, 32'h40952ea0} /* (26, 5, 31) {real, imag} */,
  {32'hc1266294, 32'h3fde89f4} /* (26, 5, 30) {real, imag} */,
  {32'h4140a3b9, 32'hc0431660} /* (26, 5, 29) {real, imag} */,
  {32'h3fef3b08, 32'hc0c7730f} /* (26, 5, 28) {real, imag} */,
  {32'h40afb832, 32'hc06875fd} /* (26, 5, 27) {real, imag} */,
  {32'hc00fc14d, 32'h405f77d2} /* (26, 5, 26) {real, imag} */,
  {32'hc17b50b0, 32'h40a7e908} /* (26, 5, 25) {real, imag} */,
  {32'hc1634d14, 32'h40abc93c} /* (26, 5, 24) {real, imag} */,
  {32'hc16c8ad8, 32'hc062b814} /* (26, 5, 23) {real, imag} */,
  {32'hc1192b67, 32'hc090e0c0} /* (26, 5, 22) {real, imag} */,
  {32'h40be0b89, 32'h3f7c5da0} /* (26, 5, 21) {real, imag} */,
  {32'h3fedada8, 32'h41608ffa} /* (26, 5, 20) {real, imag} */,
  {32'h4097e726, 32'hc0ef071a} /* (26, 5, 19) {real, imag} */,
  {32'hc071f4cd, 32'h40b03b96} /* (26, 5, 18) {real, imag} */,
  {32'hc059f602, 32'h418fca1c} /* (26, 5, 17) {real, imag} */,
  {32'h4131accf, 32'h40734edd} /* (26, 5, 16) {real, imag} */,
  {32'h41393c17, 32'hbfa3e838} /* (26, 5, 15) {real, imag} */,
  {32'h41480abf, 32'h405340f3} /* (26, 5, 14) {real, imag} */,
  {32'h412504c4, 32'h414579e9} /* (26, 5, 13) {real, imag} */,
  {32'h4116767a, 32'h40beadc9} /* (26, 5, 12) {real, imag} */,
  {32'h41167640, 32'hc1066590} /* (26, 5, 11) {real, imag} */,
  {32'hc04bc174, 32'hc0ba0186} /* (26, 5, 10) {real, imag} */,
  {32'hc0b75426, 32'hc168b77c} /* (26, 5, 9) {real, imag} */,
  {32'h400d1ccb, 32'h4182c698} /* (26, 5, 8) {real, imag} */,
  {32'hc0821f99, 32'h41608f62} /* (26, 5, 7) {real, imag} */,
  {32'hc117c016, 32'hbfd0d505} /* (26, 5, 6) {real, imag} */,
  {32'h4045e824, 32'h4161bc6e} /* (26, 5, 5) {real, imag} */,
  {32'h3fa00d4d, 32'h416fce8c} /* (26, 5, 4) {real, imag} */,
  {32'h409fcb70, 32'h4059fae4} /* (26, 5, 3) {real, imag} */,
  {32'h40ab8468, 32'hc02924d7} /* (26, 5, 2) {real, imag} */,
  {32'hc0256803, 32'h40ce1870} /* (26, 5, 1) {real, imag} */,
  {32'hbee12890, 32'h4141fafc} /* (26, 5, 0) {real, imag} */,
  {32'h402ff809, 32'h40bbf74c} /* (26, 4, 31) {real, imag} */,
  {32'hc0c5a772, 32'h41039e03} /* (26, 4, 30) {real, imag} */,
  {32'hbfa94e4a, 32'hc06286e8} /* (26, 4, 29) {real, imag} */,
  {32'h4192aec9, 32'hbf428b60} /* (26, 4, 28) {real, imag} */,
  {32'hbe995ac0, 32'h41a60f1a} /* (26, 4, 27) {real, imag} */,
  {32'hc1e5fa36, 32'h40fb5180} /* (26, 4, 26) {real, imag} */,
  {32'hc10a08e3, 32'h40c8b63e} /* (26, 4, 25) {real, imag} */,
  {32'h4126394c, 32'h3ff24d26} /* (26, 4, 24) {real, imag} */,
  {32'h41bbf36a, 32'hc13331fa} /* (26, 4, 23) {real, imag} */,
  {32'h40cccf9f, 32'h400e85a8} /* (26, 4, 22) {real, imag} */,
  {32'h41276c84, 32'h4123e724} /* (26, 4, 21) {real, imag} */,
  {32'h411bfc0c, 32'hc13af9d0} /* (26, 4, 20) {real, imag} */,
  {32'h41a6e897, 32'hc18fc288} /* (26, 4, 19) {real, imag} */,
  {32'h410c0c73, 32'hc1c65d28} /* (26, 4, 18) {real, imag} */,
  {32'hc14e8c9b, 32'hc162cf26} /* (26, 4, 17) {real, imag} */,
  {32'hbfd80ed8, 32'hbf192560} /* (26, 4, 16) {real, imag} */,
  {32'hc10abc8a, 32'h4017c9ce} /* (26, 4, 15) {real, imag} */,
  {32'h4127ab9e, 32'h4028d8a0} /* (26, 4, 14) {real, imag} */,
  {32'h41b2e218, 32'h411559be} /* (26, 4, 13) {real, imag} */,
  {32'hc0610fb2, 32'h40acae97} /* (26, 4, 12) {real, imag} */,
  {32'hbfdaab0c, 32'h4085b313} /* (26, 4, 11) {real, imag} */,
  {32'hc0913ee8, 32'h413ecb89} /* (26, 4, 10) {real, imag} */,
  {32'h40eca36f, 32'h4009de92} /* (26, 4, 9) {real, imag} */,
  {32'h41a7923c, 32'h40ec49e8} /* (26, 4, 8) {real, imag} */,
  {32'hbee745fa, 32'hc028fe5c} /* (26, 4, 7) {real, imag} */,
  {32'hc0e940bc, 32'hc0e531b2} /* (26, 4, 6) {real, imag} */,
  {32'hc1cdfd1f, 32'hc0a2a165} /* (26, 4, 5) {real, imag} */,
  {32'hc1f60ab2, 32'hc09cc9e4} /* (26, 4, 4) {real, imag} */,
  {32'hc1a29d2f, 32'hc177a74a} /* (26, 4, 3) {real, imag} */,
  {32'hc17dde4f, 32'hbfdeb4a8} /* (26, 4, 2) {real, imag} */,
  {32'h410d2e58, 32'hc10aa95e} /* (26, 4, 1) {real, imag} */,
  {32'h4176fe96, 32'h40db124a} /* (26, 4, 0) {real, imag} */,
  {32'h3ef98a20, 32'h40d8a513} /* (26, 3, 31) {real, imag} */,
  {32'h412c255a, 32'hc03a5914} /* (26, 3, 30) {real, imag} */,
  {32'h4194c342, 32'hc0e53c06} /* (26, 3, 29) {real, imag} */,
  {32'h4185704b, 32'h414272fe} /* (26, 3, 28) {real, imag} */,
  {32'h4190e528, 32'h417e432c} /* (26, 3, 27) {real, imag} */,
  {32'hbfd08c61, 32'h421bea0b} /* (26, 3, 26) {real, imag} */,
  {32'hc025f056, 32'h41963274} /* (26, 3, 25) {real, imag} */,
  {32'h40f53464, 32'h419e9a3a} /* (26, 3, 24) {real, imag} */,
  {32'h4095fc40, 32'h41c192c4} /* (26, 3, 23) {real, imag} */,
  {32'h40ff2b27, 32'h3ff164bd} /* (26, 3, 22) {real, imag} */,
  {32'h41c913d8, 32'h413042cb} /* (26, 3, 21) {real, imag} */,
  {32'h41d872cc, 32'h411dface} /* (26, 3, 20) {real, imag} */,
  {32'h40dedc58, 32'h3ed3f348} /* (26, 3, 19) {real, imag} */,
  {32'hbfebaa7b, 32'h416004d8} /* (26, 3, 18) {real, imag} */,
  {32'h3ff93b7f, 32'hc0661398} /* (26, 3, 17) {real, imag} */,
  {32'hbf269de8, 32'hc1c9d354} /* (26, 3, 16) {real, imag} */,
  {32'hc037bab0, 32'h3f5374ec} /* (26, 3, 15) {real, imag} */,
  {32'hc0fdcc4e, 32'h410872f5} /* (26, 3, 14) {real, imag} */,
  {32'hbfdc4be2, 32'h4028b130} /* (26, 3, 13) {real, imag} */,
  {32'h4132e710, 32'h3fd1d566} /* (26, 3, 12) {real, imag} */,
  {32'h413043ec, 32'hc10ac3d2} /* (26, 3, 11) {real, imag} */,
  {32'h4034c0e6, 32'hbfe002f8} /* (26, 3, 10) {real, imag} */,
  {32'h411aed3a, 32'hbfdeb520} /* (26, 3, 9) {real, imag} */,
  {32'h40d7972a, 32'h416f686e} /* (26, 3, 8) {real, imag} */,
  {32'hc1857ae2, 32'h41df3c33} /* (26, 3, 7) {real, imag} */,
  {32'hc06852f5, 32'h41ed0a96} /* (26, 3, 6) {real, imag} */,
  {32'hc08252c6, 32'h409e1d77} /* (26, 3, 5) {real, imag} */,
  {32'hc0a41a4c, 32'h41501f60} /* (26, 3, 4) {real, imag} */,
  {32'h4032bdfc, 32'h4205b232} /* (26, 3, 3) {real, imag} */,
  {32'h411cb164, 32'hbf9f4a44} /* (26, 3, 2) {real, imag} */,
  {32'h401eb9cc, 32'hc052fe16} /* (26, 3, 1) {real, imag} */,
  {32'h4151d805, 32'h4076e838} /* (26, 3, 0) {real, imag} */,
  {32'h40e5c77d, 32'h3fe88c50} /* (26, 2, 31) {real, imag} */,
  {32'h40fb6bde, 32'hc111ec11} /* (26, 2, 30) {real, imag} */,
  {32'hbfd3ef24, 32'hc13ba7ee} /* (26, 2, 29) {real, imag} */,
  {32'hc085443c, 32'hc11fe752} /* (26, 2, 28) {real, imag} */,
  {32'h3cc0ee00, 32'hc0864398} /* (26, 2, 27) {real, imag} */,
  {32'hc1d36fce, 32'hc026e2a8} /* (26, 2, 26) {real, imag} */,
  {32'hc198feb1, 32'hc16b8b2b} /* (26, 2, 25) {real, imag} */,
  {32'hc083e89f, 32'hc197a47a} /* (26, 2, 24) {real, imag} */,
  {32'hc119cf10, 32'hc10fe09c} /* (26, 2, 23) {real, imag} */,
  {32'hc1638bd3, 32'hc0024fce} /* (26, 2, 22) {real, imag} */,
  {32'hc104c07d, 32'hc064d072} /* (26, 2, 21) {real, imag} */,
  {32'h40fa3fa4, 32'hc12039ff} /* (26, 2, 20) {real, imag} */,
  {32'h4146f9ea, 32'hc1bc1922} /* (26, 2, 19) {real, imag} */,
  {32'h41a0ee79, 32'hc10c3dda} /* (26, 2, 18) {real, imag} */,
  {32'h41e5f4a5, 32'h406becb1} /* (26, 2, 17) {real, imag} */,
  {32'h3ec394e0, 32'h419d3b20} /* (26, 2, 16) {real, imag} */,
  {32'hc182fa44, 32'h41e7e815} /* (26, 2, 15) {real, imag} */,
  {32'hc188a04c, 32'h41de838c} /* (26, 2, 14) {real, imag} */,
  {32'hc1fe859b, 32'h418e06df} /* (26, 2, 13) {real, imag} */,
  {32'hc08388b2, 32'hc0c8b9be} /* (26, 2, 12) {real, imag} */,
  {32'hbf0fd540, 32'hbfb24248} /* (26, 2, 11) {real, imag} */,
  {32'hc0c95ac7, 32'h418caaf0} /* (26, 2, 10) {real, imag} */,
  {32'hbf74acb6, 32'hbfcf72d0} /* (26, 2, 9) {real, imag} */,
  {32'hc11de2f6, 32'hc0c36f24} /* (26, 2, 8) {real, imag} */,
  {32'hc170dfaa, 32'h4136a7ee} /* (26, 2, 7) {real, imag} */,
  {32'hc1418a0b, 32'h41074e44} /* (26, 2, 6) {real, imag} */,
  {32'hc0aa50dc, 32'h41066a40} /* (26, 2, 5) {real, imag} */,
  {32'h40dab4cc, 32'h40f18f30} /* (26, 2, 4) {real, imag} */,
  {32'h40b1a17e, 32'h413c5cf2} /* (26, 2, 3) {real, imag} */,
  {32'h4140ebfc, 32'h414e8e4a} /* (26, 2, 2) {real, imag} */,
  {32'h4193bd80, 32'hc026480c} /* (26, 2, 1) {real, imag} */,
  {32'hc0a6e75f, 32'h3ec1ff98} /* (26, 2, 0) {real, imag} */,
  {32'h3f4cb118, 32'hc0b1eeac} /* (26, 1, 31) {real, imag} */,
  {32'hbfa1a878, 32'hc056accf} /* (26, 1, 30) {real, imag} */,
  {32'hc103e3d3, 32'h3f3d058a} /* (26, 1, 29) {real, imag} */,
  {32'hc0f56ec9, 32'h41a33adb} /* (26, 1, 28) {real, imag} */,
  {32'hc1269eb8, 32'h4173d757} /* (26, 1, 27) {real, imag} */,
  {32'hc1a35916, 32'h40c76e7a} /* (26, 1, 26) {real, imag} */,
  {32'hc0e17af0, 32'h3fba1ea6} /* (26, 1, 25) {real, imag} */,
  {32'hc0403af2, 32'h409df412} /* (26, 1, 24) {real, imag} */,
  {32'hc0af60a2, 32'h4114f432} /* (26, 1, 23) {real, imag} */,
  {32'hc094e1ef, 32'hc0cf11f0} /* (26, 1, 22) {real, imag} */,
  {32'h41110236, 32'h414d2c9d} /* (26, 1, 21) {real, imag} */,
  {32'hc1609c78, 32'h408800cc} /* (26, 1, 20) {real, imag} */,
  {32'hc1467dba, 32'hc11b3568} /* (26, 1, 19) {real, imag} */,
  {32'hbf03d27c, 32'hc19155a4} /* (26, 1, 18) {real, imag} */,
  {32'hc196868e, 32'hc1cf992a} /* (26, 1, 17) {real, imag} */,
  {32'hc1b603b9, 32'hc013a06a} /* (26, 1, 16) {real, imag} */,
  {32'hc0abbe60, 32'hbf3fb340} /* (26, 1, 15) {real, imag} */,
  {32'h41676966, 32'hc18f21d8} /* (26, 1, 14) {real, imag} */,
  {32'h41bda3ae, 32'h40e3f45b} /* (26, 1, 13) {real, imag} */,
  {32'h41501e8e, 32'h41b18fea} /* (26, 1, 12) {real, imag} */,
  {32'h41378bd1, 32'h42114199} /* (26, 1, 11) {real, imag} */,
  {32'h41030f1e, 32'h41579c96} /* (26, 1, 10) {real, imag} */,
  {32'hc1df3017, 32'hc18f2879} /* (26, 1, 9) {real, imag} */,
  {32'hc189659e, 32'hc1d3290c} /* (26, 1, 8) {real, imag} */,
  {32'hc1928725, 32'hc1adca2e} /* (26, 1, 7) {real, imag} */,
  {32'hc209544b, 32'hc0de4796} /* (26, 1, 6) {real, imag} */,
  {32'hc190b8d4, 32'hbfd7285b} /* (26, 1, 5) {real, imag} */,
  {32'hc11bb85b, 32'h40cdc9dd} /* (26, 1, 4) {real, imag} */,
  {32'hc0406b4a, 32'h40ad76de} /* (26, 1, 3) {real, imag} */,
  {32'h3f8ffb88, 32'h41446024} /* (26, 1, 2) {real, imag} */,
  {32'hc0d8780e, 32'h404fa0b4} /* (26, 1, 1) {real, imag} */,
  {32'hbf4247d8, 32'hc0d7cd4e} /* (26, 1, 0) {real, imag} */,
  {32'hbf9d737d, 32'hc149dba6} /* (26, 0, 31) {real, imag} */,
  {32'h407d447e, 32'hc18e817c} /* (26, 0, 30) {real, imag} */,
  {32'h40afbca7, 32'h3fe41e28} /* (26, 0, 29) {real, imag} */,
  {32'h415fe426, 32'h40133864} /* (26, 0, 28) {real, imag} */,
  {32'h420d7cb8, 32'h41286eaf} /* (26, 0, 27) {real, imag} */,
  {32'h41690027, 32'h3c838940} /* (26, 0, 26) {real, imag} */,
  {32'hc167f54c, 32'h3f0729fa} /* (26, 0, 25) {real, imag} */,
  {32'hc16063e6, 32'h40944c26} /* (26, 0, 24) {real, imag} */,
  {32'h401c3b7c, 32'h4149156e} /* (26, 0, 23) {real, imag} */,
  {32'h3f82d9db, 32'hc0e13c16} /* (26, 0, 22) {real, imag} */,
  {32'hc0a7a5ac, 32'hc161b288} /* (26, 0, 21) {real, imag} */,
  {32'h40f52ba8, 32'hc1271d50} /* (26, 0, 20) {real, imag} */,
  {32'h40cce176, 32'hc1a9d9a6} /* (26, 0, 19) {real, imag} */,
  {32'hbfd06b9c, 32'hc14e03fb} /* (26, 0, 18) {real, imag} */,
  {32'hc1b4dac8, 32'h40e26cc0} /* (26, 0, 17) {real, imag} */,
  {32'hc0b34c12, 32'h3fedea97} /* (26, 0, 16) {real, imag} */,
  {32'h41025134, 32'h40fb4b62} /* (26, 0, 15) {real, imag} */,
  {32'h41a07ef0, 32'h3f933358} /* (26, 0, 14) {real, imag} */,
  {32'h41932ee0, 32'h4113216c} /* (26, 0, 13) {real, imag} */,
  {32'hc02e346b, 32'hc1273e9c} /* (26, 0, 12) {real, imag} */,
  {32'h40aba765, 32'hc0bd073e} /* (26, 0, 11) {real, imag} */,
  {32'h41065d94, 32'hc03cb2b6} /* (26, 0, 10) {real, imag} */,
  {32'h41816b7b, 32'h415de666} /* (26, 0, 9) {real, imag} */,
  {32'h418a2463, 32'h41c8406b} /* (26, 0, 8) {real, imag} */,
  {32'h411f867a, 32'hc10bdec6} /* (26, 0, 7) {real, imag} */,
  {32'h40bcde53, 32'hc1bbe78e} /* (26, 0, 6) {real, imag} */,
  {32'hc085a720, 32'hc1ef2474} /* (26, 0, 5) {real, imag} */,
  {32'h3faf5698, 32'hc1929fe1} /* (26, 0, 4) {real, imag} */,
  {32'h40ad4412, 32'hc110090d} /* (26, 0, 3) {real, imag} */,
  {32'h3faef542, 32'hc1c7fd6c} /* (26, 0, 2) {real, imag} */,
  {32'h41badcd6, 32'hc14664e4} /* (26, 0, 1) {real, imag} */,
  {32'h40c7a96a, 32'hc0acd8cd} /* (26, 0, 0) {real, imag} */,
  {32'hc0dd6c56, 32'hc085e26b} /* (25, 31, 31) {real, imag} */,
  {32'hc17e1f1c, 32'hc0e3e9cc} /* (25, 31, 30) {real, imag} */,
  {32'hc1838f74, 32'h414ec3e4} /* (25, 31, 29) {real, imag} */,
  {32'h4157cd14, 32'h40fa8f2e} /* (25, 31, 28) {real, imag} */,
  {32'h41c801df, 32'h407e81eb} /* (25, 31, 27) {real, imag} */,
  {32'h405191cc, 32'h41631e90} /* (25, 31, 26) {real, imag} */,
  {32'h3feb32b9, 32'h4197f9c8} /* (25, 31, 25) {real, imag} */,
  {32'h41c24048, 32'h4001a7c4} /* (25, 31, 24) {real, imag} */,
  {32'h414665b7, 32'hc0947222} /* (25, 31, 23) {real, imag} */,
  {32'h415b6d45, 32'h404abcb0} /* (25, 31, 22) {real, imag} */,
  {32'h41285945, 32'h4112b0ba} /* (25, 31, 21) {real, imag} */,
  {32'hc0bf17d4, 32'h403312c2} /* (25, 31, 20) {real, imag} */,
  {32'hc1a38c38, 32'hc20220b5} /* (25, 31, 19) {real, imag} */,
  {32'hc185b6a1, 32'hc1c03b18} /* (25, 31, 18) {real, imag} */,
  {32'hc09d2e7b, 32'hc183eab6} /* (25, 31, 17) {real, imag} */,
  {32'hc16de7a5, 32'hc1404a8e} /* (25, 31, 16) {real, imag} */,
  {32'hc044affe, 32'hc0ec838c} /* (25, 31, 15) {real, imag} */,
  {32'h410726c0, 32'hc1be0e6a} /* (25, 31, 14) {real, imag} */,
  {32'hc10654f1, 32'hc207b1c4} /* (25, 31, 13) {real, imag} */,
  {32'hc0860238, 32'hc1024fbc} /* (25, 31, 12) {real, imag} */,
  {32'hc0089aa4, 32'h40b2fa88} /* (25, 31, 11) {real, imag} */,
  {32'h40442f9c, 32'h40c8be44} /* (25, 31, 10) {real, imag} */,
  {32'hc12d11ee, 32'h409511e0} /* (25, 31, 9) {real, imag} */,
  {32'h40107b24, 32'hbf170fe0} /* (25, 31, 8) {real, imag} */,
  {32'h41927548, 32'hbfaefbd0} /* (25, 31, 7) {real, imag} */,
  {32'h40b2e4d0, 32'hc0cb3a28} /* (25, 31, 6) {real, imag} */,
  {32'h3f97980a, 32'hc1058140} /* (25, 31, 5) {real, imag} */,
  {32'hc121a2ca, 32'hc0085e59} /* (25, 31, 4) {real, imag} */,
  {32'hc1260010, 32'h3fe0e37c} /* (25, 31, 3) {real, imag} */,
  {32'h412cd605, 32'h4045e317} /* (25, 31, 2) {real, imag} */,
  {32'h419e48a2, 32'h3fbf2414} /* (25, 31, 1) {real, imag} */,
  {32'h3ef99090, 32'h4060390e} /* (25, 31, 0) {real, imag} */,
  {32'hc06ee02f, 32'h417a5afa} /* (25, 30, 31) {real, imag} */,
  {32'hbf3a7838, 32'h41449ebc} /* (25, 30, 30) {real, imag} */,
  {32'hc0b4a100, 32'h40393672} /* (25, 30, 29) {real, imag} */,
  {32'h41112b65, 32'hc13d8478} /* (25, 30, 28) {real, imag} */,
  {32'h4095f266, 32'hc1947968} /* (25, 30, 27) {real, imag} */,
  {32'hc14d19b7, 32'hc19ebbcd} /* (25, 30, 26) {real, imag} */,
  {32'h3fb7a5a8, 32'hc13e374d} /* (25, 30, 25) {real, imag} */,
  {32'h41652dbc, 32'h3fcac548} /* (25, 30, 24) {real, imag} */,
  {32'hc0a14c32, 32'hc09e9a0c} /* (25, 30, 23) {real, imag} */,
  {32'hbf8bf83c, 32'hc16e4767} /* (25, 30, 22) {real, imag} */,
  {32'hc00e3685, 32'hc06cfaa6} /* (25, 30, 21) {real, imag} */,
  {32'hc0b44f80, 32'h41629e34} /* (25, 30, 20) {real, imag} */,
  {32'h4019754b, 32'h40c453c5} /* (25, 30, 19) {real, imag} */,
  {32'h3ff9c06c, 32'h41a549d0} /* (25, 30, 18) {real, imag} */,
  {32'hc154469e, 32'h419d4085} /* (25, 30, 17) {real, imag} */,
  {32'h4034aa4e, 32'h4172f57c} /* (25, 30, 16) {real, imag} */,
  {32'h411e05ec, 32'hc10f5636} /* (25, 30, 15) {real, imag} */,
  {32'h41189106, 32'hc164f427} /* (25, 30, 14) {real, imag} */,
  {32'hbfa51eb0, 32'hc15ed72c} /* (25, 30, 13) {real, imag} */,
  {32'hc1916ef0, 32'h3e6d8de0} /* (25, 30, 12) {real, imag} */,
  {32'h40ad1403, 32'hbf5ff63c} /* (25, 30, 11) {real, imag} */,
  {32'h3f5d9978, 32'hc0408dd6} /* (25, 30, 10) {real, imag} */,
  {32'h3cc4ef00, 32'h4050ed59} /* (25, 30, 9) {real, imag} */,
  {32'h41aa578e, 32'h3e1a9ac8} /* (25, 30, 8) {real, imag} */,
  {32'h41ce4041, 32'hc03a70d5} /* (25, 30, 7) {real, imag} */,
  {32'hc08f9da6, 32'hc13c3aac} /* (25, 30, 6) {real, imag} */,
  {32'hc0cf7dc4, 32'hc19ee58f} /* (25, 30, 5) {real, imag} */,
  {32'hc0b21b4b, 32'hc1529140} /* (25, 30, 4) {real, imag} */,
  {32'hc1949b1a, 32'hc1227739} /* (25, 30, 3) {real, imag} */,
  {32'hc1713d2c, 32'hc13057f3} /* (25, 30, 2) {real, imag} */,
  {32'hc1179af2, 32'h3e88a334} /* (25, 30, 1) {real, imag} */,
  {32'hc0be5cb4, 32'h4101821f} /* (25, 30, 0) {real, imag} */,
  {32'h3ffc7d38, 32'hc0b232ca} /* (25, 29, 31) {real, imag} */,
  {32'h4095eb50, 32'h40b3cff0} /* (25, 29, 30) {real, imag} */,
  {32'h406eef68, 32'h4172f0d4} /* (25, 29, 29) {real, imag} */,
  {32'hc18b3f23, 32'h41920fda} /* (25, 29, 28) {real, imag} */,
  {32'hc14a72a4, 32'h4122db6c} /* (25, 29, 27) {real, imag} */,
  {32'h41177267, 32'h413c9c72} /* (25, 29, 26) {real, imag} */,
  {32'h40b79017, 32'h40eb484a} /* (25, 29, 25) {real, imag} */,
  {32'h4126abb7, 32'h410c43c6} /* (25, 29, 24) {real, imag} */,
  {32'h418d1ef3, 32'h403eb73a} /* (25, 29, 23) {real, imag} */,
  {32'h41817b20, 32'hc0b023ec} /* (25, 29, 22) {real, imag} */,
  {32'h4197c586, 32'h409b291e} /* (25, 29, 21) {real, imag} */,
  {32'h4138e732, 32'hc0ade5f5} /* (25, 29, 20) {real, imag} */,
  {32'h40bacc4b, 32'h415d25e3} /* (25, 29, 19) {real, imag} */,
  {32'hc0654c62, 32'hbec19074} /* (25, 29, 18) {real, imag} */,
  {32'hc09da851, 32'hc093f7b3} /* (25, 29, 17) {real, imag} */,
  {32'h40e5235e, 32'h4059fda5} /* (25, 29, 16) {real, imag} */,
  {32'h4194a004, 32'hc0f81da8} /* (25, 29, 15) {real, imag} */,
  {32'h409fcbdd, 32'h4095c5bf} /* (25, 29, 14) {real, imag} */,
  {32'h3f50f07c, 32'hc12b8a7c} /* (25, 29, 13) {real, imag} */,
  {32'hc0675630, 32'hc1885052} /* (25, 29, 12) {real, imag} */,
  {32'h40519284, 32'hc1587b90} /* (25, 29, 11) {real, imag} */,
  {32'hc0ace0f2, 32'hc1a784f0} /* (25, 29, 10) {real, imag} */,
  {32'hc11c1c0c, 32'hc167caee} /* (25, 29, 9) {real, imag} */,
  {32'h41422b2d, 32'h405e9df4} /* (25, 29, 8) {real, imag} */,
  {32'hc10754ce, 32'h40759e96} /* (25, 29, 7) {real, imag} */,
  {32'hc18d0a8c, 32'h4183ef39} /* (25, 29, 6) {real, imag} */,
  {32'hc086a66f, 32'h409e82d4} /* (25, 29, 5) {real, imag} */,
  {32'h40e06d11, 32'hc1cc4f93} /* (25, 29, 4) {real, imag} */,
  {32'h4141b68f, 32'hc19118da} /* (25, 29, 3) {real, imag} */,
  {32'h3fcd45f4, 32'hc0fa8d3e} /* (25, 29, 2) {real, imag} */,
  {32'h41291ae6, 32'h3fa4bb3c} /* (25, 29, 1) {real, imag} */,
  {32'h4113b96b, 32'h41053be0} /* (25, 29, 0) {real, imag} */,
  {32'h40cdaf06, 32'h40d48fbc} /* (25, 28, 31) {real, imag} */,
  {32'h40b66cd8, 32'h40eebd18} /* (25, 28, 30) {real, imag} */,
  {32'h4031242c, 32'h4116b1b9} /* (25, 28, 29) {real, imag} */,
  {32'h40228147, 32'hc079401c} /* (25, 28, 28) {real, imag} */,
  {32'hc0919f88, 32'hc195bfb8} /* (25, 28, 27) {real, imag} */,
  {32'h407b0b48, 32'hc17727ba} /* (25, 28, 26) {real, imag} */,
  {32'h40ad69b2, 32'hc1401461} /* (25, 28, 25) {real, imag} */,
  {32'h408ce075, 32'hc16b6e66} /* (25, 28, 24) {real, imag} */,
  {32'hc04f103c, 32'hc1666ee7} /* (25, 28, 23) {real, imag} */,
  {32'hc1aafebd, 32'hc03a4994} /* (25, 28, 22) {real, imag} */,
  {32'hc13fcb33, 32'hc052dc69} /* (25, 28, 21) {real, imag} */,
  {32'h4129aab9, 32'h4025b591} /* (25, 28, 20) {real, imag} */,
  {32'h41a7198f, 32'h40af13aa} /* (25, 28, 19) {real, imag} */,
  {32'h40b8fffc, 32'hbf2e6208} /* (25, 28, 18) {real, imag} */,
  {32'h413d66ca, 32'hc0a25db6} /* (25, 28, 17) {real, imag} */,
  {32'h417c94d8, 32'hc10785df} /* (25, 28, 16) {real, imag} */,
  {32'hc1248a43, 32'h41a66636} /* (25, 28, 15) {real, imag} */,
  {32'hc106733a, 32'h41b97982} /* (25, 28, 14) {real, imag} */,
  {32'hc135fce2, 32'h41450f2a} /* (25, 28, 13) {real, imag} */,
  {32'hc13d7055, 32'hc12bb012} /* (25, 28, 12) {real, imag} */,
  {32'h3ef95848, 32'hc0e0a2ff} /* (25, 28, 11) {real, imag} */,
  {32'hc16bde76, 32'hc152cd62} /* (25, 28, 10) {real, imag} */,
  {32'hc17f4d29, 32'hc1c449bb} /* (25, 28, 9) {real, imag} */,
  {32'h409673b2, 32'hc09c6afa} /* (25, 28, 8) {real, imag} */,
  {32'hbfa56728, 32'hc1376a13} /* (25, 28, 7) {real, imag} */,
  {32'hbf7ea3a8, 32'h3fe4a3fd} /* (25, 28, 6) {real, imag} */,
  {32'h3f1500fc, 32'h40aa24ab} /* (25, 28, 5) {real, imag} */,
  {32'h3e1a71e0, 32'hc08048fc} /* (25, 28, 4) {real, imag} */,
  {32'hc130cbc6, 32'h4039b2d1} /* (25, 28, 3) {real, imag} */,
  {32'hc0ca6772, 32'h4123434a} /* (25, 28, 2) {real, imag} */,
  {32'h411e3407, 32'h4076dbc6} /* (25, 28, 1) {real, imag} */,
  {32'h40aa6cb6, 32'hc061e914} /* (25, 28, 0) {real, imag} */,
  {32'hc00a3530, 32'hc0951402} /* (25, 27, 31) {real, imag} */,
  {32'hc0675e6f, 32'hc0826373} /* (25, 27, 30) {real, imag} */,
  {32'hc1257282, 32'hc05671f4} /* (25, 27, 29) {real, imag} */,
  {32'h4088c826, 32'hc12a6f23} /* (25, 27, 28) {real, imag} */,
  {32'hc18dd7c8, 32'h410a9953} /* (25, 27, 27) {real, imag} */,
  {32'hc18249ef, 32'h4181230e} /* (25, 27, 26) {real, imag} */,
  {32'h4121cba0, 32'hbfb197dc} /* (25, 27, 25) {real, imag} */,
  {32'h41a46093, 32'h4151b025} /* (25, 27, 24) {real, imag} */,
  {32'h415d23f0, 32'h41629ff0} /* (25, 27, 23) {real, imag} */,
  {32'hc01b9170, 32'h40f8c9e6} /* (25, 27, 22) {real, imag} */,
  {32'hc1076c1c, 32'h4180d90b} /* (25, 27, 21) {real, imag} */,
  {32'hc0895aa9, 32'h41453ab3} /* (25, 27, 20) {real, imag} */,
  {32'h41506b64, 32'h40c3f9e0} /* (25, 27, 19) {real, imag} */,
  {32'h41301176, 32'hc1426e60} /* (25, 27, 18) {real, imag} */,
  {32'hc19c26ab, 32'hc10fb753} /* (25, 27, 17) {real, imag} */,
  {32'hc115d585, 32'hc0ee5c74} /* (25, 27, 16) {real, imag} */,
  {32'h40920845, 32'h4032405c} /* (25, 27, 15) {real, imag} */,
  {32'h4132c8a4, 32'h40eb1044} /* (25, 27, 14) {real, imag} */,
  {32'h40161e49, 32'hbec3c1e0} /* (25, 27, 13) {real, imag} */,
  {32'hc009061a, 32'h414e605e} /* (25, 27, 12) {real, imag} */,
  {32'h3ec12e30, 32'h40dc060e} /* (25, 27, 11) {real, imag} */,
  {32'hc03bfe24, 32'h4091032a} /* (25, 27, 10) {real, imag} */,
  {32'h40095e04, 32'h4187c2aa} /* (25, 27, 9) {real, imag} */,
  {32'hc03c5e04, 32'h41db68ce} /* (25, 27, 8) {real, imag} */,
  {32'h411b801a, 32'h416103fe} /* (25, 27, 7) {real, imag} */,
  {32'h416ef115, 32'h410165a8} /* (25, 27, 6) {real, imag} */,
  {32'h410ecd78, 32'h41754400} /* (25, 27, 5) {real, imag} */,
  {32'h40b63274, 32'h3fd21ab6} /* (25, 27, 4) {real, imag} */,
  {32'hbf3593d0, 32'h400a6ce0} /* (25, 27, 3) {real, imag} */,
  {32'hbf79bb08, 32'h418cd436} /* (25, 27, 2) {real, imag} */,
  {32'hbe3fbcc0, 32'h408fed19} /* (25, 27, 1) {real, imag} */,
  {32'h40b23916, 32'hc10607fd} /* (25, 27, 0) {real, imag} */,
  {32'hc0a2eace, 32'hbefe9ab8} /* (25, 26, 31) {real, imag} */,
  {32'hc06e80fa, 32'hbf41f4dc} /* (25, 26, 30) {real, imag} */,
  {32'h408b1c40, 32'h4034e1e3} /* (25, 26, 29) {real, imag} */,
  {32'hc0065511, 32'h40a9734e} /* (25, 26, 28) {real, imag} */,
  {32'hbe8d48b8, 32'h40259885} /* (25, 26, 27) {real, imag} */,
  {32'h402c055a, 32'hc0adf102} /* (25, 26, 26) {real, imag} */,
  {32'hc0ad02f8, 32'h40b93150} /* (25, 26, 25) {real, imag} */,
  {32'h409c1ca8, 32'h40c1a230} /* (25, 26, 24) {real, imag} */,
  {32'h40dcfe69, 32'hbfecd0c6} /* (25, 26, 23) {real, imag} */,
  {32'h410a0400, 32'h4147216b} /* (25, 26, 22) {real, imag} */,
  {32'h404f2968, 32'h411b07b3} /* (25, 26, 21) {real, imag} */,
  {32'hc0b35c91, 32'hbf9c984e} /* (25, 26, 20) {real, imag} */,
  {32'hbf28a430, 32'h414fec91} /* (25, 26, 19) {real, imag} */,
  {32'h40808082, 32'h415e61e0} /* (25, 26, 18) {real, imag} */,
  {32'h3e949a4c, 32'hc0901bbe} /* (25, 26, 17) {real, imag} */,
  {32'hc0a65312, 32'h40a0f1e4} /* (25, 26, 16) {real, imag} */,
  {32'h40c1809d, 32'h408b32a4} /* (25, 26, 15) {real, imag} */,
  {32'h4135e316, 32'h4069573e} /* (25, 26, 14) {real, imag} */,
  {32'hc15299ea, 32'hc0b74502} /* (25, 26, 13) {real, imag} */,
  {32'hc171c5da, 32'hc167fde6} /* (25, 26, 12) {real, imag} */,
  {32'hc0cebdd6, 32'hc12ff319} /* (25, 26, 11) {real, imag} */,
  {32'hc0e03d5f, 32'hc087a1e2} /* (25, 26, 10) {real, imag} */,
  {32'hc0362c4a, 32'hc11dfd29} /* (25, 26, 9) {real, imag} */,
  {32'hc0bc425e, 32'hc1608f56} /* (25, 26, 8) {real, imag} */,
  {32'hc07e75e6, 32'hc108df83} /* (25, 26, 7) {real, imag} */,
  {32'hc130a59b, 32'h3fc2e6d0} /* (25, 26, 6) {real, imag} */,
  {32'hc0d227a2, 32'h410cbe4a} /* (25, 26, 5) {real, imag} */,
  {32'h408d3ceb, 32'h40ef6378} /* (25, 26, 4) {real, imag} */,
  {32'h40dffeb7, 32'hbe11c1e0} /* (25, 26, 3) {real, imag} */,
  {32'h41714752, 32'h40615cdc} /* (25, 26, 2) {real, imag} */,
  {32'h4121d2a2, 32'h4018dbc0} /* (25, 26, 1) {real, imag} */,
  {32'h4026f2f4, 32'hc0573253} /* (25, 26, 0) {real, imag} */,
  {32'hbfbd0a54, 32'hc0f8f8ca} /* (25, 25, 31) {real, imag} */,
  {32'h4064b7fd, 32'hc048ce4f} /* (25, 25, 30) {real, imag} */,
  {32'hbf38e764, 32'hbf9c4dbb} /* (25, 25, 29) {real, imag} */,
  {32'hc0f02b1a, 32'hbf02a108} /* (25, 25, 28) {real, imag} */,
  {32'hc0da25be, 32'h40f15485} /* (25, 25, 27) {real, imag} */,
  {32'h402a4872, 32'h40ca856a} /* (25, 25, 26) {real, imag} */,
  {32'hbfc23a42, 32'h414085f4} /* (25, 25, 25) {real, imag} */,
  {32'hc0719310, 32'h41641df9} /* (25, 25, 24) {real, imag} */,
  {32'hbf95c8b4, 32'h40f161d9} /* (25, 25, 23) {real, imag} */,
  {32'hc0a00c1a, 32'h410c6f94} /* (25, 25, 22) {real, imag} */,
  {32'hc0ce2aee, 32'hc0eec9f9} /* (25, 25, 21) {real, imag} */,
  {32'hc12c78ca, 32'hc10f31cf} /* (25, 25, 20) {real, imag} */,
  {32'h401e6344, 32'h3d9f6700} /* (25, 25, 19) {real, imag} */,
  {32'h40002fc1, 32'hc0dbfa32} /* (25, 25, 18) {real, imag} */,
  {32'hc0421be2, 32'hc00716fe} /* (25, 25, 17) {real, imag} */,
  {32'hc07ccfde, 32'h3fad1e76} /* (25, 25, 16) {real, imag} */,
  {32'hbf936de0, 32'hbf42be70} /* (25, 25, 15) {real, imag} */,
  {32'hc0c0ad34, 32'h3fc2c7a0} /* (25, 25, 14) {real, imag} */,
  {32'hbfbfdb24, 32'hbf88ccf2} /* (25, 25, 13) {real, imag} */,
  {32'h400710c4, 32'hc04aa9f4} /* (25, 25, 12) {real, imag} */,
  {32'hc129dabd, 32'hc0432e6e} /* (25, 25, 11) {real, imag} */,
  {32'hc0a94208, 32'h3fdff984} /* (25, 25, 10) {real, imag} */,
  {32'hbfe1730c, 32'h3fda0c5a} /* (25, 25, 9) {real, imag} */,
  {32'hc012bd9a, 32'h3f6134a0} /* (25, 25, 8) {real, imag} */,
  {32'hc14b09f6, 32'hbf5460b0} /* (25, 25, 7) {real, imag} */,
  {32'hc0f25b28, 32'hc0e1cc64} /* (25, 25, 6) {real, imag} */,
  {32'h405b5cc2, 32'h4010f8d4} /* (25, 25, 5) {real, imag} */,
  {32'h41184579, 32'h41a16979} /* (25, 25, 4) {real, imag} */,
  {32'h410252bf, 32'h413517fd} /* (25, 25, 3) {real, imag} */,
  {32'h3ffb722c, 32'hc075399a} /* (25, 25, 2) {real, imag} */,
  {32'h3ee30930, 32'hc0095c5a} /* (25, 25, 1) {real, imag} */,
  {32'h40b4bc54, 32'hc0b4459b} /* (25, 25, 0) {real, imag} */,
  {32'h408569ee, 32'h406f3ec2} /* (25, 24, 31) {real, imag} */,
  {32'hc1014571, 32'hc09a7319} /* (25, 24, 30) {real, imag} */,
  {32'hc138aa45, 32'hc12083c3} /* (25, 24, 29) {real, imag} */,
  {32'hc1303963, 32'h40a1acc8} /* (25, 24, 28) {real, imag} */,
  {32'hc0a7506a, 32'h401010f0} /* (25, 24, 27) {real, imag} */,
  {32'hbf7a3f40, 32'hc0af3386} /* (25, 24, 26) {real, imag} */,
  {32'hc027c562, 32'hc11af752} /* (25, 24, 25) {real, imag} */,
  {32'hbffbb900, 32'hc18b6eec} /* (25, 24, 24) {real, imag} */,
  {32'hbf842650, 32'hc08a4cd6} /* (25, 24, 23) {real, imag} */,
  {32'h3fdb86e4, 32'h40e5c6da} /* (25, 24, 22) {real, imag} */,
  {32'h4098e9c6, 32'h3e725f40} /* (25, 24, 21) {real, imag} */,
  {32'h414c51c2, 32'hc04a5dc2} /* (25, 24, 20) {real, imag} */,
  {32'hc0a195d6, 32'hc14bbc45} /* (25, 24, 19) {real, imag} */,
  {32'h3fd3596c, 32'hc1a7df2e} /* (25, 24, 18) {real, imag} */,
  {32'h3f9bd68c, 32'hc02d9970} /* (25, 24, 17) {real, imag} */,
  {32'hc0644fa2, 32'h3f9d4212} /* (25, 24, 16) {real, imag} */,
  {32'h3ff07c7c, 32'hc0d5712a} /* (25, 24, 15) {real, imag} */,
  {32'h3fca0514, 32'h40072cf8} /* (25, 24, 14) {real, imag} */,
  {32'hbf6b4998, 32'h40dcb3e2} /* (25, 24, 13) {real, imag} */,
  {32'hc007b4f2, 32'hbfaf5b4c} /* (25, 24, 12) {real, imag} */,
  {32'h3f58e174, 32'hc097b8f2} /* (25, 24, 11) {real, imag} */,
  {32'h41368e45, 32'hc040e644} /* (25, 24, 10) {real, imag} */,
  {32'h41895038, 32'hc0a5b75a} /* (25, 24, 9) {real, imag} */,
  {32'h408b5ff9, 32'hc0e211bd} /* (25, 24, 8) {real, imag} */,
  {32'h3e66ec20, 32'hc13df0a8} /* (25, 24, 7) {real, imag} */,
  {32'h4007dd98, 32'h3fdd69b3} /* (25, 24, 6) {real, imag} */,
  {32'h4006c7f2, 32'hc0673693} /* (25, 24, 5) {real, imag} */,
  {32'hbeff49b0, 32'h3f9f5fd6} /* (25, 24, 4) {real, imag} */,
  {32'h409c062a, 32'h4163ea0c} /* (25, 24, 3) {real, imag} */,
  {32'hbf008b00, 32'h406b00d0} /* (25, 24, 2) {real, imag} */,
  {32'h3bf44e00, 32'hc17f2f36} /* (25, 24, 1) {real, imag} */,
  {32'h40301758, 32'hc044c998} /* (25, 24, 0) {real, imag} */,
  {32'h40c99a76, 32'hc0a5199e} /* (25, 23, 31) {real, imag} */,
  {32'h40b8452b, 32'hc02f840f} /* (25, 23, 30) {real, imag} */,
  {32'h40ad903c, 32'h3f971ae4} /* (25, 23, 29) {real, imag} */,
  {32'h401117c3, 32'h403fce66} /* (25, 23, 28) {real, imag} */,
  {32'hbc18d700, 32'h40282df0} /* (25, 23, 27) {real, imag} */,
  {32'hc0bc4e40, 32'h404ef2ce} /* (25, 23, 26) {real, imag} */,
  {32'hc0750d4c, 32'h40e6ccde} /* (25, 23, 25) {real, imag} */,
  {32'hc0654d62, 32'h3f7b274c} /* (25, 23, 24) {real, imag} */,
  {32'h3e8e14b0, 32'hc13d535e} /* (25, 23, 23) {real, imag} */,
  {32'h4105a526, 32'hc15507d0} /* (25, 23, 22) {real, imag} */,
  {32'hc144fbde, 32'hc03f0743} /* (25, 23, 21) {real, imag} */,
  {32'hc10f13f0, 32'h3e9dd9a0} /* (25, 23, 20) {real, imag} */,
  {32'h406198d0, 32'hc0a149d2} /* (25, 23, 19) {real, imag} */,
  {32'h40c0b9b6, 32'hc01ccf6f} /* (25, 23, 18) {real, imag} */,
  {32'h3fedd585, 32'hc0915a5b} /* (25, 23, 17) {real, imag} */,
  {32'h40e01b1f, 32'hc03400b6} /* (25, 23, 16) {real, imag} */,
  {32'h3f1ba574, 32'h4073d7b8} /* (25, 23, 15) {real, imag} */,
  {32'hc0b3d790, 32'hc02ee26e} /* (25, 23, 14) {real, imag} */,
  {32'h409f0673, 32'hc15c6d97} /* (25, 23, 13) {real, imag} */,
  {32'h3f45daf6, 32'h3ff3a106} /* (25, 23, 12) {real, imag} */,
  {32'hc122feb4, 32'h413ed80a} /* (25, 23, 11) {real, imag} */,
  {32'hc14a8a9b, 32'h406d0d4e} /* (25, 23, 10) {real, imag} */,
  {32'hc129931f, 32'hc147346c} /* (25, 23, 9) {real, imag} */,
  {32'hc0e04636, 32'hc0814e95} /* (25, 23, 8) {real, imag} */,
  {32'h3f9ee368, 32'h3fbe3230} /* (25, 23, 7) {real, imag} */,
  {32'hc131641e, 32'hc023e6c0} /* (25, 23, 6) {real, imag} */,
  {32'hc0fff517, 32'hc0100bf2} /* (25, 23, 5) {real, imag} */,
  {32'h407481b7, 32'hc0eeeae1} /* (25, 23, 4) {real, imag} */,
  {32'h4088c4ea, 32'hc12699b8} /* (25, 23, 3) {real, imag} */,
  {32'h3fd2c4ce, 32'hbf0b0814} /* (25, 23, 2) {real, imag} */,
  {32'h3fb93afa, 32'hbfc33046} /* (25, 23, 1) {real, imag} */,
  {32'h410a584f, 32'hc07fecdc} /* (25, 23, 0) {real, imag} */,
  {32'hbf32cc46, 32'hbed58dc8} /* (25, 22, 31) {real, imag} */,
  {32'hbfbabd24, 32'h4002b836} /* (25, 22, 30) {real, imag} */,
  {32'h4035f85c, 32'h415c5ae6} /* (25, 22, 29) {real, imag} */,
  {32'h411aea14, 32'h410b7352} /* (25, 22, 28) {real, imag} */,
  {32'h4127916c, 32'hc0928a6a} /* (25, 22, 27) {real, imag} */,
  {32'h4098b6c6, 32'h3f8fa293} /* (25, 22, 26) {real, imag} */,
  {32'h3fc0d82c, 32'hc02b4c68} /* (25, 22, 25) {real, imag} */,
  {32'hbecb53a8, 32'hbf23733c} /* (25, 22, 24) {real, imag} */,
  {32'h401ef1ab, 32'h404f74b0} /* (25, 22, 23) {real, imag} */,
  {32'h3f13c3ba, 32'h3ec15340} /* (25, 22, 22) {real, imag} */,
  {32'hc00bc65a, 32'hc073bedc} /* (25, 22, 21) {real, imag} */,
  {32'hc104281a, 32'hc1255d07} /* (25, 22, 20) {real, imag} */,
  {32'hc04d4f9c, 32'hc0559bf8} /* (25, 22, 19) {real, imag} */,
  {32'hc0b3a77f, 32'hbd8a84e0} /* (25, 22, 18) {real, imag} */,
  {32'hc036ef55, 32'hc008504b} /* (25, 22, 17) {real, imag} */,
  {32'h4011f4b9, 32'hc0840158} /* (25, 22, 16) {real, imag} */,
  {32'hc0570bdc, 32'hc07c886c} /* (25, 22, 15) {real, imag} */,
  {32'h410c5b6e, 32'h40d684b4} /* (25, 22, 14) {real, imag} */,
  {32'h4181ce2e, 32'h40af7ad2} /* (25, 22, 13) {real, imag} */,
  {32'h411c6366, 32'hc1038120} /* (25, 22, 12) {real, imag} */,
  {32'h3f85ce1a, 32'hc096489a} /* (25, 22, 11) {real, imag} */,
  {32'h3f7f3358, 32'h40956ad8} /* (25, 22, 10) {real, imag} */,
  {32'hc006ddd2, 32'h40503338} /* (25, 22, 9) {real, imag} */,
  {32'hc0e54352, 32'h3f40c558} /* (25, 22, 8) {real, imag} */,
  {32'hc0d51af9, 32'h4090b833} /* (25, 22, 7) {real, imag} */,
  {32'hc004973c, 32'hc0d04c70} /* (25, 22, 6) {real, imag} */,
  {32'hc003ab63, 32'hc0dba40c} /* (25, 22, 5) {real, imag} */,
  {32'h40fdd8b8, 32'hbfd30234} /* (25, 22, 4) {real, imag} */,
  {32'h40add4e9, 32'hbfd53bd0} /* (25, 22, 3) {real, imag} */,
  {32'hbf389dd0, 32'h40913f38} /* (25, 22, 2) {real, imag} */,
  {32'h3f90925c, 32'hbf159224} /* (25, 22, 1) {real, imag} */,
  {32'hc0280eb3, 32'h3ee59335} /* (25, 22, 0) {real, imag} */,
  {32'hc054188a, 32'hbf97025a} /* (25, 21, 31) {real, imag} */,
  {32'hc08f6b90, 32'h3fc18730} /* (25, 21, 30) {real, imag} */,
  {32'hc1647278, 32'h41220e3c} /* (25, 21, 29) {real, imag} */,
  {32'hbea1e7e0, 32'h40ff8c85} /* (25, 21, 28) {real, imag} */,
  {32'h41197bd4, 32'h4118c3e6} /* (25, 21, 27) {real, imag} */,
  {32'hc01ac7e0, 32'h3f6d2ce8} /* (25, 21, 26) {real, imag} */,
  {32'hc0757812, 32'hc0b7f7a1} /* (25, 21, 25) {real, imag} */,
  {32'hc0ae23a2, 32'hc0b5241c} /* (25, 21, 24) {real, imag} */,
  {32'hc0821dc5, 32'hc0b5e458} /* (25, 21, 23) {real, imag} */,
  {32'hc10013fa, 32'hc06f3fa0} /* (25, 21, 22) {real, imag} */,
  {32'hc093eeb7, 32'hc1023898} /* (25, 21, 21) {real, imag} */,
  {32'h40a8c443, 32'hc0934c8d} /* (25, 21, 20) {real, imag} */,
  {32'h406f87c1, 32'hc0c16fee} /* (25, 21, 19) {real, imag} */,
  {32'h407dd8c2, 32'h3f546262} /* (25, 21, 18) {real, imag} */,
  {32'hbe2c9aa0, 32'h40474008} /* (25, 21, 17) {real, imag} */,
  {32'h3ff2367c, 32'h40952d9a} /* (25, 21, 16) {real, imag} */,
  {32'h4060446e, 32'h4091f958} /* (25, 21, 15) {real, imag} */,
  {32'h4141a75c, 32'h40b4e120} /* (25, 21, 14) {real, imag} */,
  {32'h412c961f, 32'h3ffe328e} /* (25, 21, 13) {real, imag} */,
  {32'hbfd4d00c, 32'h3fa9fdf0} /* (25, 21, 12) {real, imag} */,
  {32'hc0c719cd, 32'hbf3c49fc} /* (25, 21, 11) {real, imag} */,
  {32'hbd9dcf00, 32'hbf1c2f0c} /* (25, 21, 10) {real, imag} */,
  {32'h40855640, 32'h3fddd96a} /* (25, 21, 9) {real, imag} */,
  {32'h40b4406e, 32'h406f44e0} /* (25, 21, 8) {real, imag} */,
  {32'hc05ac5d7, 32'h40a88544} /* (25, 21, 7) {real, imag} */,
  {32'h3cbc37c0, 32'hc0b9d6cd} /* (25, 21, 6) {real, imag} */,
  {32'hc0234260, 32'hc0d76e72} /* (25, 21, 5) {real, imag} */,
  {32'hbf440474, 32'h40a9ae98} /* (25, 21, 4) {real, imag} */,
  {32'h3fb28e72, 32'h40228ce2} /* (25, 21, 3) {real, imag} */,
  {32'hc07b3b92, 32'h3f02a80e} /* (25, 21, 2) {real, imag} */,
  {32'hc0dd1e3a, 32'h404fbc90} /* (25, 21, 1) {real, imag} */,
  {32'hc0991dee, 32'h40ad8499} /* (25, 21, 0) {real, imag} */,
  {32'hbf42be04, 32'h400d5aff} /* (25, 20, 31) {real, imag} */,
  {32'h3fad309e, 32'h40942f33} /* (25, 20, 30) {real, imag} */,
  {32'h408b3f2f, 32'hc0d60b17} /* (25, 20, 29) {real, imag} */,
  {32'hc0759f4b, 32'h3fd464c4} /* (25, 20, 28) {real, imag} */,
  {32'hc01d6088, 32'h40850f58} /* (25, 20, 27) {real, imag} */,
  {32'h403b4f97, 32'hc084b7a9} /* (25, 20, 26) {real, imag} */,
  {32'h411b8656, 32'hbf7a4db8} /* (25, 20, 25) {real, imag} */,
  {32'h40a0e664, 32'h40015d2e} /* (25, 20, 24) {real, imag} */,
  {32'hc0857732, 32'h40615f92} /* (25, 20, 23) {real, imag} */,
  {32'h3fa61764, 32'hc027e490} /* (25, 20, 22) {real, imag} */,
  {32'h411b16fe, 32'hc08c88de} /* (25, 20, 21) {real, imag} */,
  {32'h4028f0f9, 32'hc093d162} /* (25, 20, 20) {real, imag} */,
  {32'hc0ce9220, 32'hbf611d28} /* (25, 20, 19) {real, imag} */,
  {32'hbf661f1c, 32'h3e4f8bf8} /* (25, 20, 18) {real, imag} */,
  {32'hbf0db1a0, 32'h40e570ce} /* (25, 20, 17) {real, imag} */,
  {32'hc0a36c84, 32'h41230889} /* (25, 20, 16) {real, imag} */,
  {32'h3ffdda79, 32'h407a1a94} /* (25, 20, 15) {real, imag} */,
  {32'h4045cc39, 32'hc07c5677} /* (25, 20, 14) {real, imag} */,
  {32'h400868da, 32'hc099f171} /* (25, 20, 13) {real, imag} */,
  {32'hbeb15d70, 32'hc05b8ee0} /* (25, 20, 12) {real, imag} */,
  {32'hc0987fd8, 32'h3e99f6d0} /* (25, 20, 11) {real, imag} */,
  {32'hbe9ddf8c, 32'h40c0daa4} /* (25, 20, 10) {real, imag} */,
  {32'hc061ff2a, 32'hbf335c60} /* (25, 20, 9) {real, imag} */,
  {32'hc0aaa36c, 32'hc00ab79a} /* (25, 20, 8) {real, imag} */,
  {32'hbf5633e8, 32'h3e7b7c40} /* (25, 20, 7) {real, imag} */,
  {32'hbe449480, 32'h3e5785bc} /* (25, 20, 6) {real, imag} */,
  {32'h3ea677f8, 32'h40a9e6c5} /* (25, 20, 5) {real, imag} */,
  {32'h3dca7770, 32'h40b0a252} /* (25, 20, 4) {real, imag} */,
  {32'hbf6ec74c, 32'hc06c12e0} /* (25, 20, 3) {real, imag} */,
  {32'hc092616a, 32'hc03fd376} /* (25, 20, 2) {real, imag} */,
  {32'hc073e3e6, 32'h3f30f834} /* (25, 20, 1) {real, imag} */,
  {32'hbe3be118, 32'h408d9371} /* (25, 20, 0) {real, imag} */,
  {32'hbea16932, 32'h408a7400} /* (25, 19, 31) {real, imag} */,
  {32'h3fcf4a1e, 32'h400df432} /* (25, 19, 30) {real, imag} */,
  {32'h404bef7a, 32'h404e99e8} /* (25, 19, 29) {real, imag} */,
  {32'h40866e14, 32'h4018e9be} /* (25, 19, 28) {real, imag} */,
  {32'hbfd32348, 32'h406751bd} /* (25, 19, 27) {real, imag} */,
  {32'hbfae9f9a, 32'h401b000d} /* (25, 19, 26) {real, imag} */,
  {32'hc04c1a9a, 32'h3f92c641} /* (25, 19, 25) {real, imag} */,
  {32'hc0958718, 32'hbf0ad3d8} /* (25, 19, 24) {real, imag} */,
  {32'hc095b6bd, 32'h401495b6} /* (25, 19, 23) {real, imag} */,
  {32'hc0a9b06c, 32'h40a003ba} /* (25, 19, 22) {real, imag} */,
  {32'hc04d3c62, 32'h410864a2} /* (25, 19, 21) {real, imag} */,
  {32'hbcc0c4c0, 32'h410aafda} /* (25, 19, 20) {real, imag} */,
  {32'h3ea33508, 32'hbfe53e6e} /* (25, 19, 19) {real, imag} */,
  {32'hc01c9084, 32'hc02e82c8} /* (25, 19, 18) {real, imag} */,
  {32'h3fcfda6d, 32'h4024794a} /* (25, 19, 17) {real, imag} */,
  {32'hc01e053b, 32'h3fa850ee} /* (25, 19, 16) {real, imag} */,
  {32'hc0b13ee6, 32'h3f0d1641} /* (25, 19, 15) {real, imag} */,
  {32'h3f2810e0, 32'hc01e419e} /* (25, 19, 14) {real, imag} */,
  {32'hbd54f640, 32'hc09afd84} /* (25, 19, 13) {real, imag} */,
  {32'h4071072b, 32'h402a2ce4} /* (25, 19, 12) {real, imag} */,
  {32'hc0b7eb99, 32'h3e976540} /* (25, 19, 11) {real, imag} */,
  {32'hc0eb8908, 32'h405cea2c} /* (25, 19, 10) {real, imag} */,
  {32'hc104216b, 32'h403824c8} /* (25, 19, 9) {real, imag} */,
  {32'h3fee2bac, 32'hbf5e8a7c} /* (25, 19, 8) {real, imag} */,
  {32'h4073dc8a, 32'hbf87e27d} /* (25, 19, 7) {real, imag} */,
  {32'h40a79574, 32'h3f95ba9a} /* (25, 19, 6) {real, imag} */,
  {32'hbeac134c, 32'h409984f8} /* (25, 19, 5) {real, imag} */,
  {32'hc00ea6c2, 32'hc091ad3f} /* (25, 19, 4) {real, imag} */,
  {32'h4014b191, 32'hc0cfca0b} /* (25, 19, 3) {real, imag} */,
  {32'hbe88b594, 32'h3eb45920} /* (25, 19, 2) {real, imag} */,
  {32'hbf9ba953, 32'h4047e104} /* (25, 19, 1) {real, imag} */,
  {32'h3f575470, 32'h3fbda01a} /* (25, 19, 0) {real, imag} */,
  {32'hbeec9218, 32'h3f5f6444} /* (25, 18, 31) {real, imag} */,
  {32'h3e91b4d0, 32'hc063a89a} /* (25, 18, 30) {real, imag} */,
  {32'hbf290d42, 32'hc0c2cb63} /* (25, 18, 29) {real, imag} */,
  {32'hc04d4c16, 32'hc05b9c5b} /* (25, 18, 28) {real, imag} */,
  {32'hc0271ced, 32'hc0332d7e} /* (25, 18, 27) {real, imag} */,
  {32'hbfafd9fa, 32'h40acf25e} /* (25, 18, 26) {real, imag} */,
  {32'hc051902c, 32'h407d1551} /* (25, 18, 25) {real, imag} */,
  {32'h3fd51130, 32'hbfcb561a} /* (25, 18, 24) {real, imag} */,
  {32'h4081aee3, 32'hc045a1bc} /* (25, 18, 23) {real, imag} */,
  {32'h4080dff7, 32'hbf5b34cc} /* (25, 18, 22) {real, imag} */,
  {32'h3ef2c318, 32'h3eb951d0} /* (25, 18, 21) {real, imag} */,
  {32'hc06ba0fb, 32'h3f8e0636} /* (25, 18, 20) {real, imag} */,
  {32'h3fc6bbdf, 32'h40092f90} /* (25, 18, 19) {real, imag} */,
  {32'h4081e288, 32'hc000b967} /* (25, 18, 18) {real, imag} */,
  {32'hbf476e6c, 32'hc09417ea} /* (25, 18, 17) {real, imag} */,
  {32'hc02b3e9b, 32'hc01b7393} /* (25, 18, 16) {real, imag} */,
  {32'hc0580f8e, 32'h40023562} /* (25, 18, 15) {real, imag} */,
  {32'h3e9863d4, 32'h4047a6b7} /* (25, 18, 14) {real, imag} */,
  {32'h40cd7f04, 32'h40464c86} /* (25, 18, 13) {real, imag} */,
  {32'h4090f1f1, 32'hc0610a9b} /* (25, 18, 12) {real, imag} */,
  {32'h3f4c1a25, 32'hc0621144} /* (25, 18, 11) {real, imag} */,
  {32'hbf218794, 32'h40049f56} /* (25, 18, 10) {real, imag} */,
  {32'hbfc663c0, 32'h408a1c28} /* (25, 18, 9) {real, imag} */,
  {32'hc093329d, 32'h40603650} /* (25, 18, 8) {real, imag} */,
  {32'hc043278e, 32'h3fcbcf80} /* (25, 18, 7) {real, imag} */,
  {32'hbeb84cf0, 32'h3ff8ef14} /* (25, 18, 6) {real, imag} */,
  {32'h3fe060cc, 32'h4084dc4b} /* (25, 18, 5) {real, imag} */,
  {32'hbfd5890a, 32'h3fdd293a} /* (25, 18, 4) {real, imag} */,
  {32'hc0e64e55, 32'h3f295814} /* (25, 18, 3) {real, imag} */,
  {32'hc0a66366, 32'hc067ec7e} /* (25, 18, 2) {real, imag} */,
  {32'hbff51bba, 32'hc03e2c1c} /* (25, 18, 1) {real, imag} */,
  {32'h3ff9942f, 32'h3f30345c} /* (25, 18, 0) {real, imag} */,
  {32'hbfe0a123, 32'h40138e60} /* (25, 17, 31) {real, imag} */,
  {32'hc0a2acce, 32'h40ecc6a6} /* (25, 17, 30) {real, imag} */,
  {32'hc0acfbfc, 32'h409bb6ea} /* (25, 17, 29) {real, imag} */,
  {32'hc019b692, 32'h4066c8a8} /* (25, 17, 28) {real, imag} */,
  {32'hbf3ecf82, 32'h3fb5e868} /* (25, 17, 27) {real, imag} */,
  {32'h3e8638d8, 32'hbf3dac48} /* (25, 17, 26) {real, imag} */,
  {32'hbeee4f72, 32'hc0430d54} /* (25, 17, 25) {real, imag} */,
  {32'hbfb06dec, 32'h3e0a0740} /* (25, 17, 24) {real, imag} */,
  {32'hc0359b66, 32'hbf2d5ea8} /* (25, 17, 23) {real, imag} */,
  {32'hc08b60e0, 32'hc0469f00} /* (25, 17, 22) {real, imag} */,
  {32'hc051f5a1, 32'hbeea34c0} /* (25, 17, 21) {real, imag} */,
  {32'hc020ce30, 32'hc0153872} /* (25, 17, 20) {real, imag} */,
  {32'hc05f7616, 32'hc06b8524} /* (25, 17, 19) {real, imag} */,
  {32'h3d4a0b80, 32'hc081b643} /* (25, 17, 18) {real, imag} */,
  {32'h401cc626, 32'h3e1d8aa8} /* (25, 17, 17) {real, imag} */,
  {32'hc0ffba54, 32'h402e1414} /* (25, 17, 16) {real, imag} */,
  {32'hc0d35823, 32'h3fe31688} /* (25, 17, 15) {real, imag} */,
  {32'h3fbce9c1, 32'hbfe0f352} /* (25, 17, 14) {real, imag} */,
  {32'hbf96045b, 32'hc0564408} /* (25, 17, 13) {real, imag} */,
  {32'hc0a1d035, 32'hbf3ae898} /* (25, 17, 12) {real, imag} */,
  {32'hbfdcaf00, 32'h3ff2f8b2} /* (25, 17, 11) {real, imag} */,
  {32'h404da3bc, 32'h3ff5ab9c} /* (25, 17, 10) {real, imag} */,
  {32'h408539ac, 32'hbf013060} /* (25, 17, 9) {real, imag} */,
  {32'hbf1dfe34, 32'hbf05eb20} /* (25, 17, 8) {real, imag} */,
  {32'hc0968822, 32'h3f8778b4} /* (25, 17, 7) {real, imag} */,
  {32'hc074e603, 32'hbed4b698} /* (25, 17, 6) {real, imag} */,
  {32'h3f5f33ac, 32'hbea2e504} /* (25, 17, 5) {real, imag} */,
  {32'h403250f0, 32'h3fb8af20} /* (25, 17, 4) {real, imag} */,
  {32'h3e91eb4c, 32'h4027669c} /* (25, 17, 3) {real, imag} */,
  {32'hbf1d3460, 32'h3fd5f42a} /* (25, 17, 2) {real, imag} */,
  {32'h3ea6beb8, 32'h404ea0a0} /* (25, 17, 1) {real, imag} */,
  {32'h3fc7b436, 32'h3f0019a0} /* (25, 17, 0) {real, imag} */,
  {32'h403a4cdd, 32'hbfe69b6a} /* (25, 16, 31) {real, imag} */,
  {32'h3f124848, 32'h3ebac510} /* (25, 16, 30) {real, imag} */,
  {32'hbfbb0d20, 32'hbfd65e58} /* (25, 16, 29) {real, imag} */,
  {32'hc0636a02, 32'hc08491f4} /* (25, 16, 28) {real, imag} */,
  {32'hc01fc1f5, 32'hbfedec80} /* (25, 16, 27) {real, imag} */,
  {32'hbf56ca90, 32'hc032ba32} /* (25, 16, 26) {real, imag} */,
  {32'h3f82930a, 32'hbea9eee0} /* (25, 16, 25) {real, imag} */,
  {32'h407e9dd6, 32'hc0077d16} /* (25, 16, 24) {real, imag} */,
  {32'h40020b0a, 32'hc019f046} /* (25, 16, 23) {real, imag} */,
  {32'hbfbce380, 32'hc05a4c62} /* (25, 16, 22) {real, imag} */,
  {32'hbf766578, 32'hc052a1e0} /* (25, 16, 21) {real, imag} */,
  {32'h3ff5ad2e, 32'h3db18200} /* (25, 16, 20) {real, imag} */,
  {32'hc037aed8, 32'h3fa456a0} /* (25, 16, 19) {real, imag} */,
  {32'hc072d9e0, 32'hbe973ec0} /* (25, 16, 18) {real, imag} */,
  {32'hbdaf3500, 32'hbff4ae08} /* (25, 16, 17) {real, imag} */,
  {32'hbf8915d4, 32'h3f5daf38} /* (25, 16, 16) {real, imag} */,
  {32'hbf81e5e4, 32'h3dd0ea40} /* (25, 16, 15) {real, imag} */,
  {32'h3e511b90, 32'hbe7b7520} /* (25, 16, 14) {real, imag} */,
  {32'h3f86f958, 32'h3fd10a28} /* (25, 16, 13) {real, imag} */,
  {32'h3f9b1f50, 32'h3df1a760} /* (25, 16, 12) {real, imag} */,
  {32'h4023c797, 32'h3fe2e1a5} /* (25, 16, 11) {real, imag} */,
  {32'h409a2380, 32'h4111db3c} /* (25, 16, 10) {real, imag} */,
  {32'h407bac3c, 32'h3ffc5d6c} /* (25, 16, 9) {real, imag} */,
  {32'h40a6c348, 32'hc05122a6} /* (25, 16, 8) {real, imag} */,
  {32'h40a6873c, 32'hc0324eda} /* (25, 16, 7) {real, imag} */,
  {32'hbd5af3e0, 32'hbf87f110} /* (25, 16, 6) {real, imag} */,
  {32'hbff33628, 32'h402fc91a} /* (25, 16, 5) {real, imag} */,
  {32'hbf6cdc5e, 32'h403b04ae} /* (25, 16, 4) {real, imag} */,
  {32'hbeb48190, 32'h3fbfe29a} /* (25, 16, 3) {real, imag} */,
  {32'hc00794ce, 32'h4085d0b5} /* (25, 16, 2) {real, imag} */,
  {32'hc04723cc, 32'h402da5cc} /* (25, 16, 1) {real, imag} */,
  {32'hbf98330e, 32'h3fb27950} /* (25, 16, 0) {real, imag} */,
  {32'hbf15766a, 32'hbf6f97e2} /* (25, 15, 31) {real, imag} */,
  {32'hbf55b788, 32'hc03f5f34} /* (25, 15, 30) {real, imag} */,
  {32'hc0c2584a, 32'h408d687a} /* (25, 15, 29) {real, imag} */,
  {32'hbf87b533, 32'h4041a69e} /* (25, 15, 28) {real, imag} */,
  {32'h3f9511c1, 32'hbf3e5fcc} /* (25, 15, 27) {real, imag} */,
  {32'hc08818a6, 32'hc07ecaca} /* (25, 15, 26) {real, imag} */,
  {32'hbf1abbb3, 32'hc097affe} /* (25, 15, 25) {real, imag} */,
  {32'hbf165198, 32'hbfc98dc4} /* (25, 15, 24) {real, imag} */,
  {32'hbe884c34, 32'hbf81b3a0} /* (25, 15, 23) {real, imag} */,
  {32'hbe9afba8, 32'hbfc0fc70} /* (25, 15, 22) {real, imag} */,
  {32'hbfb49592, 32'hc0980d9a} /* (25, 15, 21) {real, imag} */,
  {32'h3f3b5168, 32'hbf900de4} /* (25, 15, 20) {real, imag} */,
  {32'hbdc7b640, 32'h404ba7f4} /* (25, 15, 19) {real, imag} */,
  {32'h3e903050, 32'h3fe4ec34} /* (25, 15, 18) {real, imag} */,
  {32'hc01b9700, 32'h40524012} /* (25, 15, 17) {real, imag} */,
  {32'hbef624e0, 32'hbf12836e} /* (25, 15, 16) {real, imag} */,
  {32'hbff6114c, 32'hc04ee98c} /* (25, 15, 15) {real, imag} */,
  {32'hc088f659, 32'h3fd22962} /* (25, 15, 14) {real, imag} */,
  {32'hc01f69f2, 32'h3f509000} /* (25, 15, 13) {real, imag} */,
  {32'hc06a624a, 32'h40142cae} /* (25, 15, 12) {real, imag} */,
  {32'hc0685eca, 32'hc02d2157} /* (25, 15, 11) {real, imag} */,
  {32'hc03a425c, 32'hc046d51e} /* (25, 15, 10) {real, imag} */,
  {32'hc08b92fc, 32'h3f139b40} /* (25, 15, 9) {real, imag} */,
  {32'hc05e0e0d, 32'h3ff5f910} /* (25, 15, 8) {real, imag} */,
  {32'hc052e7b0, 32'hbff40ff4} /* (25, 15, 7) {real, imag} */,
  {32'hc0244429, 32'hbfcf645e} /* (25, 15, 6) {real, imag} */,
  {32'hc051b237, 32'hc0224d28} /* (25, 15, 5) {real, imag} */,
  {32'h3dace100, 32'hc04dd9c4} /* (25, 15, 4) {real, imag} */,
  {32'h3ff9b3bd, 32'hbf291b9e} /* (25, 15, 3) {real, imag} */,
  {32'h3fcb0b68, 32'h404e1edf} /* (25, 15, 2) {real, imag} */,
  {32'hc0448255, 32'h40251600} /* (25, 15, 1) {real, imag} */,
  {32'hbfd8803c, 32'hbf0b6400} /* (25, 15, 0) {real, imag} */,
  {32'hc0be353c, 32'hbf2ac57c} /* (25, 14, 31) {real, imag} */,
  {32'hc09d3623, 32'hbfc0dbe4} /* (25, 14, 30) {real, imag} */,
  {32'h4013c71e, 32'hbf6f7078} /* (25, 14, 29) {real, imag} */,
  {32'h40541c0c, 32'hc023ba93} /* (25, 14, 28) {real, imag} */,
  {32'h40779f61, 32'h3f40352a} /* (25, 14, 27) {real, imag} */,
  {32'h3fcab9b6, 32'h4063da97} /* (25, 14, 26) {real, imag} */,
  {32'h4025a818, 32'h4083b27c} /* (25, 14, 25) {real, imag} */,
  {32'h3f451da0, 32'h3fc8714e} /* (25, 14, 24) {real, imag} */,
  {32'h3f4747c2, 32'h3ea31694} /* (25, 14, 23) {real, imag} */,
  {32'h4037dcae, 32'h3f2abd84} /* (25, 14, 22) {real, imag} */,
  {32'h3f124e14, 32'hc0832d41} /* (25, 14, 21) {real, imag} */,
  {32'hc050d1e7, 32'hc06da165} /* (25, 14, 20) {real, imag} */,
  {32'hbfb562ab, 32'hc08cb614} /* (25, 14, 19) {real, imag} */,
  {32'h4056d26c, 32'hbf93b272} /* (25, 14, 18) {real, imag} */,
  {32'h3db25fa0, 32'h400bd348} /* (25, 14, 17) {real, imag} */,
  {32'h40003d83, 32'h40602d71} /* (25, 14, 16) {real, imag} */,
  {32'h4058084e, 32'h401c2cbe} /* (25, 14, 15) {real, imag} */,
  {32'h3ffe62fd, 32'hbfcb54ee} /* (25, 14, 14) {real, imag} */,
  {32'h404db888, 32'hbe2f8ab8} /* (25, 14, 13) {real, imag} */,
  {32'h40a12077, 32'h3dd51c60} /* (25, 14, 12) {real, imag} */,
  {32'hbd37be50, 32'h40aec8f2} /* (25, 14, 11) {real, imag} */,
  {32'hbda1c160, 32'h40e039bf} /* (25, 14, 10) {real, imag} */,
  {32'h40e034a8, 32'h3e0050d0} /* (25, 14, 9) {real, imag} */,
  {32'h40a5ea3b, 32'hc0f6c1d8} /* (25, 14, 8) {real, imag} */,
  {32'h3fb2287c, 32'hc072bd46} /* (25, 14, 7) {real, imag} */,
  {32'hc0979e2c, 32'hbf9ea154} /* (25, 14, 6) {real, imag} */,
  {32'hbfcbd31c, 32'hc03c79b6} /* (25, 14, 5) {real, imag} */,
  {32'hbc0addc0, 32'hbfff574a} /* (25, 14, 4) {real, imag} */,
  {32'h40d2b1c3, 32'h40559a33} /* (25, 14, 3) {real, imag} */,
  {32'h403d358c, 32'h400dabf2} /* (25, 14, 2) {real, imag} */,
  {32'hc06defaf, 32'hc0bcdbd2} /* (25, 14, 1) {real, imag} */,
  {32'hc018f1d8, 32'hc0c17534} /* (25, 14, 0) {real, imag} */,
  {32'hbec93332, 32'h401ce69c} /* (25, 13, 31) {real, imag} */,
  {32'h3fae822e, 32'h40622d52} /* (25, 13, 30) {real, imag} */,
  {32'h40f7b6b3, 32'h40465f88} /* (25, 13, 29) {real, imag} */,
  {32'h3f08eea0, 32'hbf9bebdc} /* (25, 13, 28) {real, imag} */,
  {32'hc05e71d4, 32'hbfe75d2e} /* (25, 13, 27) {real, imag} */,
  {32'h40165a97, 32'h408083ce} /* (25, 13, 26) {real, imag} */,
  {32'hbef42810, 32'hbe4c7bb8} /* (25, 13, 25) {real, imag} */,
  {32'h3b5ba400, 32'hc0539176} /* (25, 13, 24) {real, imag} */,
  {32'hc09ae92f, 32'hc0ab82ee} /* (25, 13, 23) {real, imag} */,
  {32'hc0276ffc, 32'hc091144a} /* (25, 13, 22) {real, imag} */,
  {32'hbfcfa40c, 32'h40412d1c} /* (25, 13, 21) {real, imag} */,
  {32'h4025acce, 32'h40899ce1} /* (25, 13, 20) {real, imag} */,
  {32'h409070f4, 32'h3db06120} /* (25, 13, 19) {real, imag} */,
  {32'h3f91531b, 32'h3fd65905} /* (25, 13, 18) {real, imag} */,
  {32'hbd8ac150, 32'h3ffd3130} /* (25, 13, 17) {real, imag} */,
  {32'h40b2634e, 32'h408a39fc} /* (25, 13, 16) {real, imag} */,
  {32'h406c5337, 32'h3cde8c20} /* (25, 13, 15) {real, imag} */,
  {32'h3fb09298, 32'hbfb25c4d} /* (25, 13, 14) {real, imag} */,
  {32'hc085e5a2, 32'h3f443834} /* (25, 13, 13) {real, imag} */,
  {32'hc0fa659e, 32'hbfbf5420} /* (25, 13, 12) {real, imag} */,
  {32'hbf793328, 32'hc073c4f4} /* (25, 13, 11) {real, imag} */,
  {32'hbf387e04, 32'hc0f5fed2} /* (25, 13, 10) {real, imag} */,
  {32'hc0a22376, 32'hc1155dd7} /* (25, 13, 9) {real, imag} */,
  {32'hc0af423c, 32'h3fcc1752} /* (25, 13, 8) {real, imag} */,
  {32'hc07fb78c, 32'h3fa0441d} /* (25, 13, 7) {real, imag} */,
  {32'hbfa14e5a, 32'hbf7e309c} /* (25, 13, 6) {real, imag} */,
  {32'h402589d6, 32'h402cec6f} /* (25, 13, 5) {real, imag} */,
  {32'h3fc10882, 32'h40c38ce3} /* (25, 13, 4) {real, imag} */,
  {32'h40a74990, 32'h4071734e} /* (25, 13, 3) {real, imag} */,
  {32'h40872815, 32'h40f6c142} /* (25, 13, 2) {real, imag} */,
  {32'h401f048e, 32'hbf1f8af8} /* (25, 13, 1) {real, imag} */,
  {32'h402e6e9c, 32'hc0213c0b} /* (25, 13, 0) {real, imag} */,
  {32'h3ee888f8, 32'hc02ef47f} /* (25, 12, 31) {real, imag} */,
  {32'h4078722d, 32'h4090a04b} /* (25, 12, 30) {real, imag} */,
  {32'hc02920e2, 32'hbf9fcb9c} /* (25, 12, 29) {real, imag} */,
  {32'hbf452b44, 32'hc0c9eea5} /* (25, 12, 28) {real, imag} */,
  {32'hc00aaee4, 32'h3f836560} /* (25, 12, 27) {real, imag} */,
  {32'hbf0f8514, 32'h409ab2cf} /* (25, 12, 26) {real, imag} */,
  {32'h3fceb5cc, 32'h4040e580} /* (25, 12, 25) {real, imag} */,
  {32'hc00f27c1, 32'h407156d2} /* (25, 12, 24) {real, imag} */,
  {32'hbf0f2216, 32'hbf30ee48} /* (25, 12, 23) {real, imag} */,
  {32'h3e87d310, 32'hbfa2e169} /* (25, 12, 22) {real, imag} */,
  {32'hc048d788, 32'hc00a31e0} /* (25, 12, 21) {real, imag} */,
  {32'h3fa1b49a, 32'hc12fe7eb} /* (25, 12, 20) {real, imag} */,
  {32'hbe9c4ee8, 32'hc11865fe} /* (25, 12, 19) {real, imag} */,
  {32'h3fa8aefe, 32'hc055a498} /* (25, 12, 18) {real, imag} */,
  {32'h40ee9ddc, 32'hbf307ed4} /* (25, 12, 17) {real, imag} */,
  {32'hbf63a854, 32'hc004cce0} /* (25, 12, 16) {real, imag} */,
  {32'hc0b7a987, 32'h40059964} /* (25, 12, 15) {real, imag} */,
  {32'h40ef9878, 32'hbfb799e2} /* (25, 12, 14) {real, imag} */,
  {32'h410fb072, 32'h4019e562} /* (25, 12, 13) {real, imag} */,
  {32'h408a9df6, 32'hbf833d48} /* (25, 12, 12) {real, imag} */,
  {32'hc0b60d6c, 32'hc029456e} /* (25, 12, 11) {real, imag} */,
  {32'hc02f30e6, 32'hbf680270} /* (25, 12, 10) {real, imag} */,
  {32'h407b9a06, 32'hbf8ab2e8} /* (25, 12, 9) {real, imag} */,
  {32'h4003b57b, 32'h40c82fdd} /* (25, 12, 8) {real, imag} */,
  {32'hbf4adfe8, 32'h3f3456c0} /* (25, 12, 7) {real, imag} */,
  {32'h3f8d6378, 32'hbfa29832} /* (25, 12, 6) {real, imag} */,
  {32'hc02efc11, 32'hbf76a948} /* (25, 12, 5) {real, imag} */,
  {32'h3f2c1fc2, 32'hc0976e0a} /* (25, 12, 4) {real, imag} */,
  {32'h40474c23, 32'hc0993414} /* (25, 12, 3) {real, imag} */,
  {32'h403dd7e9, 32'h4075ad52} /* (25, 12, 2) {real, imag} */,
  {32'h40b98b51, 32'h40b3e1fc} /* (25, 12, 1) {real, imag} */,
  {32'hc00360e6, 32'hc02d6d4e} /* (25, 12, 0) {real, imag} */,
  {32'hbf8ba2e1, 32'h40a079fc} /* (25, 11, 31) {real, imag} */,
  {32'hc061d3e0, 32'h40ff3d70} /* (25, 11, 30) {real, imag} */,
  {32'h40843eb9, 32'hbfe00b34} /* (25, 11, 29) {real, imag} */,
  {32'h40a7ef34, 32'hc0073162} /* (25, 11, 28) {real, imag} */,
  {32'h4083e614, 32'h3eb158e0} /* (25, 11, 27) {real, imag} */,
  {32'h40603890, 32'hbfbe1f8c} /* (25, 11, 26) {real, imag} */,
  {32'h3eff34b4, 32'h3f945fec} /* (25, 11, 25) {real, imag} */,
  {32'hbfc30ff8, 32'hc00e73eb} /* (25, 11, 24) {real, imag} */,
  {32'h40234a56, 32'hc0b91730} /* (25, 11, 23) {real, imag} */,
  {32'hbfa28d54, 32'hc0531fb0} /* (25, 11, 22) {real, imag} */,
  {32'h401d5b32, 32'h3ffba1d8} /* (25, 11, 21) {real, imag} */,
  {32'hc09f0ec3, 32'hc0a23921} /* (25, 11, 20) {real, imag} */,
  {32'hc0f47ede, 32'hc109487f} /* (25, 11, 19) {real, imag} */,
  {32'h403a8680, 32'hbfa40421} /* (25, 11, 18) {real, imag} */,
  {32'h4103a9de, 32'hc08c0784} /* (25, 11, 17) {real, imag} */,
  {32'h3f199000, 32'hc07b7ec3} /* (25, 11, 16) {real, imag} */,
  {32'h3ee18cd0, 32'hc09167d0} /* (25, 11, 15) {real, imag} */,
  {32'h3ef6f550, 32'h3e803b08} /* (25, 11, 14) {real, imag} */,
  {32'hc1125279, 32'h404307b3} /* (25, 11, 13) {real, imag} */,
  {32'hc13a3408, 32'h41287e31} /* (25, 11, 12) {real, imag} */,
  {32'hc0ec5d7b, 32'h40a2ec16} /* (25, 11, 11) {real, imag} */,
  {32'h4113b670, 32'h40a57880} /* (25, 11, 10) {real, imag} */,
  {32'hbef944e4, 32'hc0676897} /* (25, 11, 9) {real, imag} */,
  {32'hc09bb95a, 32'hc033a194} /* (25, 11, 8) {real, imag} */,
  {32'h401fd3e7, 32'h40079c5c} /* (25, 11, 7) {real, imag} */,
  {32'h3f9e8251, 32'h402d5f0e} /* (25, 11, 6) {real, imag} */,
  {32'hbf8676b7, 32'h3fe777be} /* (25, 11, 5) {real, imag} */,
  {32'hbec38bf8, 32'h40977240} /* (25, 11, 4) {real, imag} */,
  {32'hbdd56be0, 32'h40e6e5a3} /* (25, 11, 3) {real, imag} */,
  {32'hbf07c2de, 32'hc04376f4} /* (25, 11, 2) {real, imag} */,
  {32'h404f0b65, 32'hbe8b74a0} /* (25, 11, 1) {real, imag} */,
  {32'h3ec15b70, 32'h40a90f7b} /* (25, 11, 0) {real, imag} */,
  {32'h3fa29af1, 32'h404c2052} /* (25, 10, 31) {real, imag} */,
  {32'h40bc5f81, 32'hc042b4fa} /* (25, 10, 30) {real, imag} */,
  {32'h41470329, 32'hbea48a80} /* (25, 10, 29) {real, imag} */,
  {32'h410c9118, 32'h40a85baf} /* (25, 10, 28) {real, imag} */,
  {32'h40d60e20, 32'h41231c1b} /* (25, 10, 27) {real, imag} */,
  {32'h410416db, 32'h40313060} /* (25, 10, 26) {real, imag} */,
  {32'h40a6dbd0, 32'hbffc7d70} /* (25, 10, 25) {real, imag} */,
  {32'h40e16dac, 32'hbfe9ff7a} /* (25, 10, 24) {real, imag} */,
  {32'hbfdaad7a, 32'hc08e91f5} /* (25, 10, 23) {real, imag} */,
  {32'hbfd37237, 32'hc11d6992} /* (25, 10, 22) {real, imag} */,
  {32'hc100b77c, 32'h4058ffe0} /* (25, 10, 21) {real, imag} */,
  {32'hc164b93e, 32'h40de4efa} /* (25, 10, 20) {real, imag} */,
  {32'hc0a51744, 32'h3fb234b8} /* (25, 10, 19) {real, imag} */,
  {32'hc0bcefd1, 32'hbead1c98} /* (25, 10, 18) {real, imag} */,
  {32'hc061f013, 32'h408ac12c} /* (25, 10, 17) {real, imag} */,
  {32'h409dad4a, 32'hc09c07a0} /* (25, 10, 16) {real, imag} */,
  {32'h41476555, 32'hbffac540} /* (25, 10, 15) {real, imag} */,
  {32'h41489ba0, 32'hbf63eb00} /* (25, 10, 14) {real, imag} */,
  {32'hc0da29fe, 32'hc08dd52c} /* (25, 10, 13) {real, imag} */,
  {32'hbf9212d4, 32'hbfbb210c} /* (25, 10, 12) {real, imag} */,
  {32'h409c854a, 32'hbd95e780} /* (25, 10, 11) {real, imag} */,
  {32'hc0b90561, 32'h40ba83a0} /* (25, 10, 10) {real, imag} */,
  {32'hc02a9a6a, 32'h405f4546} /* (25, 10, 9) {real, imag} */,
  {32'h408ae1fc, 32'hc0476bbe} /* (25, 10, 8) {real, imag} */,
  {32'hc0aa8e19, 32'hbeec7310} /* (25, 10, 7) {real, imag} */,
  {32'hc105cd6c, 32'h408e1818} /* (25, 10, 6) {real, imag} */,
  {32'hc0a7afb6, 32'h4157122c} /* (25, 10, 5) {real, imag} */,
  {32'hc09a2e26, 32'h4162ec3e} /* (25, 10, 4) {real, imag} */,
  {32'hc1141e6c, 32'h40a693d2} /* (25, 10, 3) {real, imag} */,
  {32'hbffa79c0, 32'hc11132e8} /* (25, 10, 2) {real, imag} */,
  {32'h403dd4e6, 32'hc090567c} /* (25, 10, 1) {real, imag} */,
  {32'h3f0e6974, 32'hbfab5b91} /* (25, 10, 0) {real, imag} */,
  {32'h40b71d4a, 32'h3f8f7122} /* (25, 9, 31) {real, imag} */,
  {32'h40be77a3, 32'hc00c81f9} /* (25, 9, 30) {real, imag} */,
  {32'h408693b6, 32'hc127db24} /* (25, 9, 29) {real, imag} */,
  {32'h40b277a4, 32'hbee8eef4} /* (25, 9, 28) {real, imag} */,
  {32'hc0b4803c, 32'h4019608c} /* (25, 9, 27) {real, imag} */,
  {32'h3f968130, 32'hc02eac76} /* (25, 9, 26) {real, imag} */,
  {32'hc062bd70, 32'hc05c603b} /* (25, 9, 25) {real, imag} */,
  {32'hc04eaf82, 32'h409aa962} /* (25, 9, 24) {real, imag} */,
  {32'hc0c8471e, 32'h414a09cc} /* (25, 9, 23) {real, imag} */,
  {32'hc12db38a, 32'h40841359} /* (25, 9, 22) {real, imag} */,
  {32'hc10d1ce8, 32'h405d9167} /* (25, 9, 21) {real, imag} */,
  {32'h4048086e, 32'h4163ae29} /* (25, 9, 20) {real, imag} */,
  {32'h4114ffc4, 32'h41025256} /* (25, 9, 19) {real, imag} */,
  {32'hbfc8d6ee, 32'h411a693a} /* (25, 9, 18) {real, imag} */,
  {32'hbfae8b65, 32'h41125dc6} /* (25, 9, 17) {real, imag} */,
  {32'h4114a798, 32'h40817a21} /* (25, 9, 16) {real, imag} */,
  {32'h41076261, 32'hc09ed420} /* (25, 9, 15) {real, imag} */,
  {32'hc0433728, 32'hc03f6ef4} /* (25, 9, 14) {real, imag} */,
  {32'hc0b47447, 32'h40a586da} /* (25, 9, 13) {real, imag} */,
  {32'hbfc0a3f9, 32'hc02a72fd} /* (25, 9, 12) {real, imag} */,
  {32'hc0c2f264, 32'h4098c365} /* (25, 9, 11) {real, imag} */,
  {32'h3f101390, 32'h416184c2} /* (25, 9, 10) {real, imag} */,
  {32'h41094c4d, 32'hc051cdc8} /* (25, 9, 9) {real, imag} */,
  {32'h3f3d98fc, 32'hc11170f4} /* (25, 9, 8) {real, imag} */,
  {32'hc0a0f4a3, 32'hc179f82c} /* (25, 9, 7) {real, imag} */,
  {32'hc0fe3998, 32'hc1354882} /* (25, 9, 6) {real, imag} */,
  {32'hc0ad3ac1, 32'hbf68ec52} /* (25, 9, 5) {real, imag} */,
  {32'hc0764fab, 32'hbfa24abc} /* (25, 9, 4) {real, imag} */,
  {32'hbf63ab74, 32'hbd9ec5c0} /* (25, 9, 3) {real, imag} */,
  {32'hbfa7310c, 32'hc102f1e4} /* (25, 9, 2) {real, imag} */,
  {32'h3ead0408, 32'hbc014300} /* (25, 9, 1) {real, imag} */,
  {32'h40626463, 32'hbe2062b8} /* (25, 9, 0) {real, imag} */,
  {32'hc064292a, 32'hc172666c} /* (25, 8, 31) {real, imag} */,
  {32'hc0ba2f1e, 32'hc11d922a} /* (25, 8, 30) {real, imag} */,
  {32'hc14fb923, 32'h4119d5c9} /* (25, 8, 29) {real, imag} */,
  {32'hc115facf, 32'h4181f396} /* (25, 8, 28) {real, imag} */,
  {32'h41261351, 32'h411e9ee0} /* (25, 8, 27) {real, imag} */,
  {32'hbfc0ec98, 32'h40285bb8} /* (25, 8, 26) {real, imag} */,
  {32'hc0d36c8b, 32'h4083de99} /* (25, 8, 25) {real, imag} */,
  {32'h40f6e3b4, 32'hc0846871} /* (25, 8, 24) {real, imag} */,
  {32'h4199ff45, 32'h411595b5} /* (25, 8, 23) {real, imag} */,
  {32'h41196f0a, 32'h40d136de} /* (25, 8, 22) {real, imag} */,
  {32'h40ab6508, 32'h3fd7b398} /* (25, 8, 21) {real, imag} */,
  {32'h410da5f6, 32'h4133dffc} /* (25, 8, 20) {real, imag} */,
  {32'h4025a81b, 32'h410bd44f} /* (25, 8, 19) {real, imag} */,
  {32'h407f6cae, 32'h40be5950} /* (25, 8, 18) {real, imag} */,
  {32'hc0ecda9b, 32'h405c6cd8} /* (25, 8, 17) {real, imag} */,
  {32'hc154c7e0, 32'h3fdc2e82} /* (25, 8, 16) {real, imag} */,
  {32'h40bd6525, 32'h3ff26788} /* (25, 8, 15) {real, imag} */,
  {32'h416fccf6, 32'h3f4bf06a} /* (25, 8, 14) {real, imag} */,
  {32'h40fd8aad, 32'hc110526d} /* (25, 8, 13) {real, imag} */,
  {32'hc104ce28, 32'h3ea3eee0} /* (25, 8, 12) {real, imag} */,
  {32'hc0bcebf4, 32'hc01e0515} /* (25, 8, 11) {real, imag} */,
  {32'h40b012a2, 32'h405dffe4} /* (25, 8, 10) {real, imag} */,
  {32'h4064b714, 32'h4130879f} /* (25, 8, 9) {real, imag} */,
  {32'hbfcdb4ac, 32'h40988e25} /* (25, 8, 8) {real, imag} */,
  {32'hc1539c88, 32'h40df1541} /* (25, 8, 7) {real, imag} */,
  {32'hc0ee8bc0, 32'hbecfb98c} /* (25, 8, 6) {real, imag} */,
  {32'h40dbb1fb, 32'hbe801b78} /* (25, 8, 5) {real, imag} */,
  {32'h409ed133, 32'h40e91274} /* (25, 8, 4) {real, imag} */,
  {32'hc16c0a85, 32'h402b3790} /* (25, 8, 3) {real, imag} */,
  {32'hc0d695a2, 32'h40b6abc8} /* (25, 8, 2) {real, imag} */,
  {32'h40a2e5e6, 32'h413f5af2} /* (25, 8, 1) {real, imag} */,
  {32'h405c0dda, 32'hbf913851} /* (25, 8, 0) {real, imag} */,
  {32'h41046712, 32'hbfba8dc6} /* (25, 7, 31) {real, imag} */,
  {32'h40e8539c, 32'hc0953855} /* (25, 7, 30) {real, imag} */,
  {32'h400a9b59, 32'h405afbda} /* (25, 7, 29) {real, imag} */,
  {32'h403c0c8c, 32'hc09a0563} /* (25, 7, 28) {real, imag} */,
  {32'hc08e4f12, 32'hbff6ae64} /* (25, 7, 27) {real, imag} */,
  {32'h400597ee, 32'hc1230e9b} /* (25, 7, 26) {real, imag} */,
  {32'h3f2dbad0, 32'hc02978c8} /* (25, 7, 25) {real, imag} */,
  {32'hc025bff0, 32'hc04b00cc} /* (25, 7, 24) {real, imag} */,
  {32'hc08cd54c, 32'hbff5e4cc} /* (25, 7, 23) {real, imag} */,
  {32'h416423df, 32'h404236ee} /* (25, 7, 22) {real, imag} */,
  {32'h41aa18bc, 32'h40fceecb} /* (25, 7, 21) {real, imag} */,
  {32'h3f7367f8, 32'hc0b4b5e6} /* (25, 7, 20) {real, imag} */,
  {32'hc18e7ee2, 32'hc11fc753} /* (25, 7, 19) {real, imag} */,
  {32'hc11dfea5, 32'hc0bf1eaa} /* (25, 7, 18) {real, imag} */,
  {32'hc11f874c, 32'hc115e9c4} /* (25, 7, 17) {real, imag} */,
  {32'h40ba4b1d, 32'hbf650178} /* (25, 7, 16) {real, imag} */,
  {32'h40dc79f4, 32'h416451c5} /* (25, 7, 15) {real, imag} */,
  {32'h40399e90, 32'h413b0584} /* (25, 7, 14) {real, imag} */,
  {32'h40e79589, 32'h40593e1f} /* (25, 7, 13) {real, imag} */,
  {32'hc0964a11, 32'h41383057} /* (25, 7, 12) {real, imag} */,
  {32'hbf4f1910, 32'hc0b1fd4b} /* (25, 7, 11) {real, imag} */,
  {32'h40e85eb0, 32'hbf15dfe8} /* (25, 7, 10) {real, imag} */,
  {32'h40cb958f, 32'h40bbc6e6} /* (25, 7, 9) {real, imag} */,
  {32'h3faf8d39, 32'h41027cc4} /* (25, 7, 8) {real, imag} */,
  {32'h405ef310, 32'h4174d85f} /* (25, 7, 7) {real, imag} */,
  {32'h4125f9aa, 32'h40d3aa94} /* (25, 7, 6) {real, imag} */,
  {32'h40e5a3e3, 32'h411870fd} /* (25, 7, 5) {real, imag} */,
  {32'h40a152ac, 32'h40c72dfd} /* (25, 7, 4) {real, imag} */,
  {32'hc02abb51, 32'h4084f1b0} /* (25, 7, 3) {real, imag} */,
  {32'hbf5b333c, 32'h4099ea8f} /* (25, 7, 2) {real, imag} */,
  {32'hc12f9200, 32'hc1579a04} /* (25, 7, 1) {real, imag} */,
  {32'hbdb47920, 32'hc1269c80} /* (25, 7, 0) {real, imag} */,
  {32'h3e50f450, 32'hbef58ee0} /* (25, 6, 31) {real, imag} */,
  {32'h3eed3d0c, 32'hc0571277} /* (25, 6, 30) {real, imag} */,
  {32'hc0f1a01c, 32'h3f89aeca} /* (25, 6, 29) {real, imag} */,
  {32'hc09708a0, 32'hc18425e4} /* (25, 6, 28) {real, imag} */,
  {32'h3fc95c26, 32'hc0b50522} /* (25, 6, 27) {real, imag} */,
  {32'h40012360, 32'h400fc35a} /* (25, 6, 26) {real, imag} */,
  {32'h40ac4cc4, 32'h410e29fa} /* (25, 6, 25) {real, imag} */,
  {32'hc0dec26e, 32'h4197c51e} /* (25, 6, 24) {real, imag} */,
  {32'hc117d810, 32'hbfd0c2c2} /* (25, 6, 23) {real, imag} */,
  {32'hc0a2ebf3, 32'h409330be} /* (25, 6, 22) {real, imag} */,
  {32'hc0b430aa, 32'hc161c35d} /* (25, 6, 21) {real, imag} */,
  {32'h3f8515a4, 32'hc0644597} /* (25, 6, 20) {real, imag} */,
  {32'h41294084, 32'h413b0707} /* (25, 6, 19) {real, imag} */,
  {32'h406972ac, 32'hbf337c48} /* (25, 6, 18) {real, imag} */,
  {32'h3fbb52ff, 32'hc04b0f51} /* (25, 6, 17) {real, imag} */,
  {32'h3eb74458, 32'h410f29d0} /* (25, 6, 16) {real, imag} */,
  {32'h3f16f068, 32'h4173c02e} /* (25, 6, 15) {real, imag} */,
  {32'h3fb37ce0, 32'h4121903e} /* (25, 6, 14) {real, imag} */,
  {32'h4031d26e, 32'hc09e613e} /* (25, 6, 13) {real, imag} */,
  {32'h410cc8f6, 32'hbfce8944} /* (25, 6, 12) {real, imag} */,
  {32'h41485711, 32'h3f27c870} /* (25, 6, 11) {real, imag} */,
  {32'h3ff53664, 32'hc088025e} /* (25, 6, 10) {real, imag} */,
  {32'h402bded6, 32'hc04c408d} /* (25, 6, 9) {real, imag} */,
  {32'h40ad4f60, 32'hc11e1e7c} /* (25, 6, 8) {real, imag} */,
  {32'hc1245192, 32'hc11334cd} /* (25, 6, 7) {real, imag} */,
  {32'hc0cba20e, 32'h411d9586} /* (25, 6, 6) {real, imag} */,
  {32'h41301377, 32'h404f715f} /* (25, 6, 5) {real, imag} */,
  {32'hbfce24dc, 32'hc0a4a8b6} /* (25, 6, 4) {real, imag} */,
  {32'h40ddc653, 32'hc12bd12a} /* (25, 6, 3) {real, imag} */,
  {32'h404d403a, 32'hc0efa426} /* (25, 6, 2) {real, imag} */,
  {32'hc16b2650, 32'hc090401d} /* (25, 6, 1) {real, imag} */,
  {32'hc1463789, 32'h401ac63d} /* (25, 6, 0) {real, imag} */,
  {32'hc04c7cce, 32'hc08eae46} /* (25, 5, 31) {real, imag} */,
  {32'hbfa51fb6, 32'hc003ed84} /* (25, 5, 30) {real, imag} */,
  {32'h40214a96, 32'hc19ae5fc} /* (25, 5, 29) {real, imag} */,
  {32'h409b642c, 32'hc158b7f3} /* (25, 5, 28) {real, imag} */,
  {32'hc107c19d, 32'hc01ad848} /* (25, 5, 27) {real, imag} */,
  {32'hc189569d, 32'h40bde6c6} /* (25, 5, 26) {real, imag} */,
  {32'hc1905fff, 32'hc0ce9a07} /* (25, 5, 25) {real, imag} */,
  {32'hc19bd9c1, 32'hc17860f3} /* (25, 5, 24) {real, imag} */,
  {32'h41118e34, 32'h3e678280} /* (25, 5, 23) {real, imag} */,
  {32'h41cd80f8, 32'hc0123e7c} /* (25, 5, 22) {real, imag} */,
  {32'h41a1d816, 32'h405fd0e6} /* (25, 5, 21) {real, imag} */,
  {32'h3fbd5943, 32'h412bd755} /* (25, 5, 20) {real, imag} */,
  {32'h3ffaff74, 32'hc113e42a} /* (25, 5, 19) {real, imag} */,
  {32'h411f0a6e, 32'hc1594abc} /* (25, 5, 18) {real, imag} */,
  {32'hc01f4e18, 32'h4077cd9c} /* (25, 5, 17) {real, imag} */,
  {32'h3f8e4888, 32'h4071a4bf} /* (25, 5, 16) {real, imag} */,
  {32'h418c5b56, 32'h403296be} /* (25, 5, 15) {real, imag} */,
  {32'h4126dc7c, 32'hc085001c} /* (25, 5, 14) {real, imag} */,
  {32'hc0028743, 32'hc194d5ac} /* (25, 5, 13) {real, imag} */,
  {32'h41259a8e, 32'hc125a1ae} /* (25, 5, 12) {real, imag} */,
  {32'h416da4f2, 32'hc03bd2f4} /* (25, 5, 11) {real, imag} */,
  {32'hbfcc8bbd, 32'h4092b012} /* (25, 5, 10) {real, imag} */,
  {32'h4020cc18, 32'hc06c2d54} /* (25, 5, 9) {real, imag} */,
  {32'h414f7e67, 32'hc0e50a40} /* (25, 5, 8) {real, imag} */,
  {32'h41c5f13d, 32'hc106efd2} /* (25, 5, 7) {real, imag} */,
  {32'h4196839a, 32'hbfaebfe0} /* (25, 5, 6) {real, imag} */,
  {32'h4184439c, 32'h4060f7d2} /* (25, 5, 5) {real, imag} */,
  {32'h40bfd8e6, 32'hc03b6d8b} /* (25, 5, 4) {real, imag} */,
  {32'hc13e0cf7, 32'h4090522d} /* (25, 5, 3) {real, imag} */,
  {32'hc126964e, 32'h4110e48d} /* (25, 5, 2) {real, imag} */,
  {32'hc0d0f8a3, 32'hbf49cf48} /* (25, 5, 1) {real, imag} */,
  {32'hc0a222a2, 32'hc105a539} /* (25, 5, 0) {real, imag} */,
  {32'hc11f12cd, 32'h40bc33a4} /* (25, 4, 31) {real, imag} */,
  {32'hc0cf12ec, 32'h3f202890} /* (25, 4, 30) {real, imag} */,
  {32'h41659755, 32'h40d44dce} /* (25, 4, 29) {real, imag} */,
  {32'hc02a9783, 32'h4000fc5c} /* (25, 4, 28) {real, imag} */,
  {32'hc197c9b8, 32'hbfb25b88} /* (25, 4, 27) {real, imag} */,
  {32'hc187fdef, 32'h40f03e5f} /* (25, 4, 26) {real, imag} */,
  {32'hc0a334e0, 32'h40a263b2} /* (25, 4, 25) {real, imag} */,
  {32'h3f5385c2, 32'hc01ad332} /* (25, 4, 24) {real, imag} */,
  {32'h4088abd6, 32'h41255eb5} /* (25, 4, 23) {real, imag} */,
  {32'h41899569, 32'h406280e0} /* (25, 4, 22) {real, imag} */,
  {32'hc07902fc, 32'h4016b929} /* (25, 4, 21) {real, imag} */,
  {32'hc195a336, 32'h40b20c98} /* (25, 4, 20) {real, imag} */,
  {32'h3ee1d1c0, 32'hbe9dbcc8} /* (25, 4, 19) {real, imag} */,
  {32'h41845225, 32'h40e42273} /* (25, 4, 18) {real, imag} */,
  {32'h418ca415, 32'h4145b961} /* (25, 4, 17) {real, imag} */,
  {32'h402169d0, 32'h401a2170} /* (25, 4, 16) {real, imag} */,
  {32'h3e9f86e0, 32'h4054f15c} /* (25, 4, 15) {real, imag} */,
  {32'hc132a8ee, 32'h40ac6bbc} /* (25, 4, 14) {real, imag} */,
  {32'hc0fc658c, 32'hc023609a} /* (25, 4, 13) {real, imag} */,
  {32'hc0066fb4, 32'h3f658698} /* (25, 4, 12) {real, imag} */,
  {32'hc01419e9, 32'h41b6bf1f} /* (25, 4, 11) {real, imag} */,
  {32'h41220e02, 32'h412f418e} /* (25, 4, 10) {real, imag} */,
  {32'h4173b307, 32'hbd7f0a00} /* (25, 4, 9) {real, imag} */,
  {32'h3fe8ef22, 32'h3f88df5f} /* (25, 4, 8) {real, imag} */,
  {32'h41920fc0, 32'h4086982c} /* (25, 4, 7) {real, imag} */,
  {32'h41592718, 32'hc01730cd} /* (25, 4, 6) {real, imag} */,
  {32'hc0a8b408, 32'h401ba29e} /* (25, 4, 5) {real, imag} */,
  {32'hc0f661eb, 32'hc00388fe} /* (25, 4, 4) {real, imag} */,
  {32'hc0c158c0, 32'h4067d4b5} /* (25, 4, 3) {real, imag} */,
  {32'h4067b0d1, 32'h40cbc584} /* (25, 4, 2) {real, imag} */,
  {32'h41271691, 32'h40cc1cfb} /* (25, 4, 1) {real, imag} */,
  {32'h3fcef09a, 32'h3f6e67b0} /* (25, 4, 0) {real, imag} */,
  {32'hc0192314, 32'hc0a97ef0} /* (25, 3, 31) {real, imag} */,
  {32'hc1072cdd, 32'h40aacca6} /* (25, 3, 30) {real, imag} */,
  {32'hc0cbd474, 32'h4103ec8c} /* (25, 3, 29) {real, imag} */,
  {32'h3f899390, 32'h40aa3d99} /* (25, 3, 28) {real, imag} */,
  {32'hc11f72c6, 32'hc0a42e56} /* (25, 3, 27) {real, imag} */,
  {32'hc0390a61, 32'hc05c6800} /* (25, 3, 26) {real, imag} */,
  {32'h3f61a118, 32'hc09ae220} /* (25, 3, 25) {real, imag} */,
  {32'hc00bacec, 32'hc19ab9fb} /* (25, 3, 24) {real, imag} */,
  {32'hc033eb88, 32'hc0b3d3ab} /* (25, 3, 23) {real, imag} */,
  {32'hc069723e, 32'h408c7a04} /* (25, 3, 22) {real, imag} */,
  {32'hc116e09c, 32'hbfdcbaa0} /* (25, 3, 21) {real, imag} */,
  {32'hc113ce38, 32'hc14e0216} /* (25, 3, 20) {real, imag} */,
  {32'h406433a6, 32'hc11b333d} /* (25, 3, 19) {real, imag} */,
  {32'h410cf0ea, 32'h4037e36c} /* (25, 3, 18) {real, imag} */,
  {32'hc0ac80a5, 32'hc02ba9b8} /* (25, 3, 17) {real, imag} */,
  {32'hc14a94fb, 32'h412c7581} /* (25, 3, 16) {real, imag} */,
  {32'hc18c10fc, 32'h4082c180} /* (25, 3, 15) {real, imag} */,
  {32'hc18841cf, 32'h3f1928f8} /* (25, 3, 14) {real, imag} */,
  {32'hc04d8a05, 32'h4026e00a} /* (25, 3, 13) {real, imag} */,
  {32'h41953561, 32'h406aad7e} /* (25, 3, 12) {real, imag} */,
  {32'h402b83fc, 32'hbe48d940} /* (25, 3, 11) {real, imag} */,
  {32'hc168f3b7, 32'hc0c8de2e} /* (25, 3, 10) {real, imag} */,
  {32'hc184e911, 32'h414584b2} /* (25, 3, 9) {real, imag} */,
  {32'h4064204c, 32'h412f01d9} /* (25, 3, 8) {real, imag} */,
  {32'hbf43c7e4, 32'h414a6772} /* (25, 3, 7) {real, imag} */,
  {32'h3fccf880, 32'hc18cb043} /* (25, 3, 6) {real, imag} */,
  {32'h40f6c105, 32'hc1e2dad3} /* (25, 3, 5) {real, imag} */,
  {32'hbfd3282c, 32'hc13122c2} /* (25, 3, 4) {real, imag} */,
  {32'hc10fb241, 32'h3f7e2970} /* (25, 3, 3) {real, imag} */,
  {32'hc0c186f9, 32'h400e4bc3} /* (25, 3, 2) {real, imag} */,
  {32'hc186fc36, 32'hc045a898} /* (25, 3, 1) {real, imag} */,
  {32'hc170e8f5, 32'hc14b33ae} /* (25, 3, 0) {real, imag} */,
  {32'hc022eee5, 32'hbfd0bae0} /* (25, 2, 31) {real, imag} */,
  {32'h417e1db0, 32'hc1cca9de} /* (25, 2, 30) {real, imag} */,
  {32'h3f0d9fc4, 32'hc160e8bc} /* (25, 2, 29) {real, imag} */,
  {32'h403f19fd, 32'h40a1e30c} /* (25, 2, 28) {real, imag} */,
  {32'h41140232, 32'hc0e57b72} /* (25, 2, 27) {real, imag} */,
  {32'h40010414, 32'hc1917d8d} /* (25, 2, 26) {real, imag} */,
  {32'h408c0d68, 32'h3fd03428} /* (25, 2, 25) {real, imag} */,
  {32'hc0abe48c, 32'h40bdf110} /* (25, 2, 24) {real, imag} */,
  {32'hc0c7203e, 32'h40f51d54} /* (25, 2, 23) {real, imag} */,
  {32'hc14f7b02, 32'h416ba605} /* (25, 2, 22) {real, imag} */,
  {32'h4094360e, 32'h3f811954} /* (25, 2, 21) {real, imag} */,
  {32'h4133d41c, 32'hc12d34f0} /* (25, 2, 20) {real, imag} */,
  {32'hc089770c, 32'hc1341816} /* (25, 2, 19) {real, imag} */,
  {32'hc18185bf, 32'h40d19e78} /* (25, 2, 18) {real, imag} */,
  {32'hbfe7dad0, 32'h40b74ba5} /* (25, 2, 17) {real, imag} */,
  {32'hc0c52d8d, 32'hc1068d2c} /* (25, 2, 16) {real, imag} */,
  {32'hc1b71dcc, 32'hc1831777} /* (25, 2, 15) {real, imag} */,
  {32'hc0ff146c, 32'hc19f973b} /* (25, 2, 14) {real, imag} */,
  {32'h4099aa24, 32'hc077befa} /* (25, 2, 13) {real, imag} */,
  {32'h4116de18, 32'hbe9487d0} /* (25, 2, 12) {real, imag} */,
  {32'h40c0644d, 32'hc065a799} /* (25, 2, 11) {real, imag} */,
  {32'hc08fb7d1, 32'hc10d6a80} /* (25, 2, 10) {real, imag} */,
  {32'hc106c47a, 32'h4030a5cf} /* (25, 2, 9) {real, imag} */,
  {32'hbf4885c0, 32'h4028bcdc} /* (25, 2, 8) {real, imag} */,
  {32'h3e02ba80, 32'hbe771230} /* (25, 2, 7) {real, imag} */,
  {32'hc13e44af, 32'hc14f041c} /* (25, 2, 6) {real, imag} */,
  {32'hc1ec96eb, 32'hc1fa83d9} /* (25, 2, 5) {real, imag} */,
  {32'hbfc0ab54, 32'hc1f39280} /* (25, 2, 4) {real, imag} */,
  {32'h3d996400, 32'hc1cdd31c} /* (25, 2, 3) {real, imag} */,
  {32'hc0301b48, 32'hc0cd6eda} /* (25, 2, 2) {real, imag} */,
  {32'hc08c046e, 32'hc066575c} /* (25, 2, 1) {real, imag} */,
  {32'hbfec9580, 32'hc0aae562} /* (25, 2, 0) {real, imag} */,
  {32'hc0e0e5cc, 32'hc0a457f7} /* (25, 1, 31) {real, imag} */,
  {32'h4074efa0, 32'h40a949ec} /* (25, 1, 30) {real, imag} */,
  {32'h40d97437, 32'h3eb5fcc0} /* (25, 1, 29) {real, imag} */,
  {32'h416b33c0, 32'hbea9f2d8} /* (25, 1, 28) {real, imag} */,
  {32'h41b61037, 32'hc081b3a0} /* (25, 1, 27) {real, imag} */,
  {32'h40809787, 32'hc0f511d8} /* (25, 1, 26) {real, imag} */,
  {32'hbf92ba17, 32'h409b7c38} /* (25, 1, 25) {real, imag} */,
  {32'hc0a4d1f0, 32'h415e3fbb} /* (25, 1, 24) {real, imag} */,
  {32'hc08e7f52, 32'h4073e4c3} /* (25, 1, 23) {real, imag} */,
  {32'hc0ff81b6, 32'hc0a5ce24} /* (25, 1, 22) {real, imag} */,
  {32'hc10723f3, 32'hbf7ea398} /* (25, 1, 21) {real, imag} */,
  {32'h40c03574, 32'h411b051a} /* (25, 1, 20) {real, imag} */,
  {32'hbe319700, 32'h3e3a6f00} /* (25, 1, 19) {real, imag} */,
  {32'hc1346a69, 32'hc078b12c} /* (25, 1, 18) {real, imag} */,
  {32'h407223f3, 32'h40cdc87a} /* (25, 1, 17) {real, imag} */,
  {32'h415747bb, 32'hc0441250} /* (25, 1, 16) {real, imag} */,
  {32'h407de58a, 32'hc14f746c} /* (25, 1, 15) {real, imag} */,
  {32'hbff49380, 32'hc1123c5d} /* (25, 1, 14) {real, imag} */,
  {32'hc093d80a, 32'hc103859a} /* (25, 1, 13) {real, imag} */,
  {32'hc0271194, 32'hc1c7d66a} /* (25, 1, 12) {real, imag} */,
  {32'hc15dce3d, 32'hc1487a94} /* (25, 1, 11) {real, imag} */,
  {32'hc1b9bf70, 32'h41dcc25d} /* (25, 1, 10) {real, imag} */,
  {32'hc19cb931, 32'h4220156e} /* (25, 1, 9) {real, imag} */,
  {32'hc19b0f46, 32'h41f86cf1} /* (25, 1, 8) {real, imag} */,
  {32'hc11c8bdc, 32'h41c09a8f} /* (25, 1, 7) {real, imag} */,
  {32'hc0ca73ec, 32'h407cd1bd} /* (25, 1, 6) {real, imag} */,
  {32'hc0bb3fa8, 32'hc15bb8be} /* (25, 1, 5) {real, imag} */,
  {32'hc0531908, 32'hbf17cdfc} /* (25, 1, 4) {real, imag} */,
  {32'hc05eecf6, 32'h408215bd} /* (25, 1, 3) {real, imag} */,
  {32'h4104a093, 32'h41293bcb} /* (25, 1, 2) {real, imag} */,
  {32'hc13829f4, 32'h4161427e} /* (25, 1, 1) {real, imag} */,
  {32'hc109e4ae, 32'hc056bbae} /* (25, 1, 0) {real, imag} */,
  {32'hc0a69cc0, 32'hc061f937} /* (25, 0, 31) {real, imag} */,
  {32'hc11a8794, 32'h410fb774} /* (25, 0, 30) {real, imag} */,
  {32'hc13c3481, 32'h41851be8} /* (25, 0, 29) {real, imag} */,
  {32'hbfdecb38, 32'h419b5fb1} /* (25, 0, 28) {real, imag} */,
  {32'h40b9b022, 32'h4178125a} /* (25, 0, 27) {real, imag} */,
  {32'hc125b394, 32'hc0ab2ed9} /* (25, 0, 26) {real, imag} */,
  {32'hc0e3a228, 32'hc18ef86c} /* (25, 0, 25) {real, imag} */,
  {32'h40f1afd9, 32'hc131025c} /* (25, 0, 24) {real, imag} */,
  {32'hc103b926, 32'h3fdff23d} /* (25, 0, 23) {real, imag} */,
  {32'h4106ecec, 32'h414190fe} /* (25, 0, 22) {real, imag} */,
  {32'h4156bb78, 32'h419f55f4} /* (25, 0, 21) {real, imag} */,
  {32'h41107f02, 32'h415c8cd9} /* (25, 0, 20) {real, imag} */,
  {32'hc1348216, 32'h4133ca2e} /* (25, 0, 19) {real, imag} */,
  {32'hc1883bca, 32'h418328d8} /* (25, 0, 18) {real, imag} */,
  {32'h40be94cc, 32'hc040f3f8} /* (25, 0, 17) {real, imag} */,
  {32'h414a4cf6, 32'h41650266} /* (25, 0, 16) {real, imag} */,
  {32'hc0c6517b, 32'h4155ca9c} /* (25, 0, 15) {real, imag} */,
  {32'hc0d2c60e, 32'h4135a194} /* (25, 0, 14) {real, imag} */,
  {32'hc196ae04, 32'h412be29b} /* (25, 0, 13) {real, imag} */,
  {32'hc17809be, 32'h40a14da4} /* (25, 0, 12) {real, imag} */,
  {32'h402ff965, 32'hbf771c8e} /* (25, 0, 11) {real, imag} */,
  {32'h3ff122be, 32'hbfdb53dc} /* (25, 0, 10) {real, imag} */,
  {32'h416c8d23, 32'h3f7801c0} /* (25, 0, 9) {real, imag} */,
  {32'hbf8dca18, 32'hc0da92ff} /* (25, 0, 8) {real, imag} */,
  {32'hbeff1a60, 32'hc1217526} /* (25, 0, 7) {real, imag} */,
  {32'h3ca5cfc0, 32'h419e36d0} /* (25, 0, 6) {real, imag} */,
  {32'h4166746f, 32'h4107d14e} /* (25, 0, 5) {real, imag} */,
  {32'h3fcbe6d5, 32'h402a3e5a} /* (25, 0, 4) {real, imag} */,
  {32'h3fb61f30, 32'h40d4c4f4} /* (25, 0, 3) {real, imag} */,
  {32'h40194518, 32'hc0eb00b1} /* (25, 0, 2) {real, imag} */,
  {32'h418df6e2, 32'hc101fe1a} /* (25, 0, 1) {real, imag} */,
  {32'h40674965, 32'hc09b5f46} /* (25, 0, 0) {real, imag} */,
  {32'hc18776b6, 32'hbff98fd8} /* (24, 31, 31) {real, imag} */,
  {32'hc1e52462, 32'hc16a7df0} /* (24, 31, 30) {real, imag} */,
  {32'hc22818f8, 32'hc195aca4} /* (24, 31, 29) {real, imag} */,
  {32'hc221e600, 32'hc1df4313} /* (24, 31, 28) {real, imag} */,
  {32'hc23d944f, 32'hc1b259de} /* (24, 31, 27) {real, imag} */,
  {32'hc1d4efaf, 32'hc1bc2582} /* (24, 31, 26) {real, imag} */,
  {32'hc1556465, 32'hc1bb1037} /* (24, 31, 25) {real, imag} */,
  {32'hc20f34f7, 32'hc10402dc} /* (24, 31, 24) {real, imag} */,
  {32'hc20a9a31, 32'hc1e84aad} /* (24, 31, 23) {real, imag} */,
  {32'hc207e15a, 32'hc23d112f} /* (24, 31, 22) {real, imag} */,
  {32'hc172c596, 32'hc2176e1a} /* (24, 31, 21) {real, imag} */,
  {32'h41a583a3, 32'hc1c5259a} /* (24, 31, 20) {real, imag} */,
  {32'h41ebe5c8, 32'hc073d96d} /* (24, 31, 19) {real, imag} */,
  {32'h41be4688, 32'h3fc4c910} /* (24, 31, 18) {real, imag} */,
  {32'h41d7f516, 32'h4085e818} /* (24, 31, 17) {real, imag} */,
  {32'h421c97f4, 32'h41b96738} /* (24, 31, 16) {real, imag} */,
  {32'h420c96db, 32'h420a9f77} /* (24, 31, 15) {real, imag} */,
  {32'h41e4f6dd, 32'h42170e2c} /* (24, 31, 14) {real, imag} */,
  {32'h41bd9500, 32'h41b43b7a} /* (24, 31, 13) {real, imag} */,
  {32'h423ebe7c, 32'h41b7ad9b} /* (24, 31, 12) {real, imag} */,
  {32'h4231cf12, 32'h41a3b6c0} /* (24, 31, 11) {real, imag} */,
  {32'hc15d6eef, 32'hc0170510} /* (24, 31, 10) {real, imag} */,
  {32'hc1afd198, 32'hbeb7bb80} /* (24, 31, 9) {real, imag} */,
  {32'hc10e9e88, 32'h4118a037} /* (24, 31, 8) {real, imag} */,
  {32'hc0fb7be6, 32'hc115518a} /* (24, 31, 7) {real, imag} */,
  {32'hc1a167bb, 32'hc19f9278} /* (24, 31, 6) {real, imag} */,
  {32'hc20f5c72, 32'hc1c83815} /* (24, 31, 5) {real, imag} */,
  {32'hc206ff52, 32'hc220dd07} /* (24, 31, 4) {real, imag} */,
  {32'hc20e6312, 32'hc20088d8} /* (24, 31, 3) {real, imag} */,
  {32'hc19449da, 32'hc2251a58} /* (24, 31, 2) {real, imag} */,
  {32'hc1b7ea06, 32'hc2222905} /* (24, 31, 1) {real, imag} */,
  {32'hc1deca3f, 32'hc117a0d4} /* (24, 31, 0) {real, imag} */,
  {32'h4191debf, 32'h417fe5f8} /* (24, 30, 31) {real, imag} */,
  {32'h41a2d021, 32'h42010882} /* (24, 30, 30) {real, imag} */,
  {32'h41b12854, 32'h41e6ac6c} /* (24, 30, 29) {real, imag} */,
  {32'h41964d49, 32'h3f3b18a0} /* (24, 30, 28) {real, imag} */,
  {32'h41e30bf2, 32'h4181c38e} /* (24, 30, 27) {real, imag} */,
  {32'h41c7cc44, 32'h41bf224a} /* (24, 30, 26) {real, imag} */,
  {32'h41a6087a, 32'h41a153ea} /* (24, 30, 25) {real, imag} */,
  {32'h418ad810, 32'h4167721f} /* (24, 30, 24) {real, imag} */,
  {32'h419e3c28, 32'h4122027e} /* (24, 30, 23) {real, imag} */,
  {32'h41a089f3, 32'h412771bd} /* (24, 30, 22) {real, imag} */,
  {32'h40b4fd76, 32'h3f189ae0} /* (24, 30, 21) {real, imag} */,
  {32'hc18be2ac, 32'hc1917162} /* (24, 30, 20) {real, imag} */,
  {32'hc17b0c7c, 32'hc1d6631d} /* (24, 30, 19) {real, imag} */,
  {32'hc0f7b98a, 32'hc20bc0ba} /* (24, 30, 18) {real, imag} */,
  {32'hc1558fcc, 32'hc21e57e5} /* (24, 30, 17) {real, imag} */,
  {32'hc1841843, 32'hc214495a} /* (24, 30, 16) {real, imag} */,
  {32'hc1c881cb, 32'hc19498c0} /* (24, 30, 15) {real, imag} */,
  {32'hc200515a, 32'h3f7dbc08} /* (24, 30, 14) {real, imag} */,
  {32'hc1bf4ced, 32'hc0af8c7c} /* (24, 30, 13) {real, imag} */,
  {32'hc1d2a8ea, 32'hc0b896f2} /* (24, 30, 12) {real, imag} */,
  {32'hc157d21c, 32'hc12d8bac} /* (24, 30, 11) {real, imag} */,
  {32'h41a1b907, 32'h41a5c87d} /* (24, 30, 10) {real, imag} */,
  {32'h41c9bdea, 32'h4213dd1c} /* (24, 30, 9) {real, imag} */,
  {32'h41b28ce9, 32'h42121567} /* (24, 30, 8) {real, imag} */,
  {32'h41ad4922, 32'h41e7e40a} /* (24, 30, 7) {real, imag} */,
  {32'h41e06e3f, 32'h41e7a3c2} /* (24, 30, 6) {real, imag} */,
  {32'h41eab1a6, 32'h418ba88a} /* (24, 30, 5) {real, imag} */,
  {32'h41fbcc92, 32'h4013cb28} /* (24, 30, 4) {real, imag} */,
  {32'h41e86b3d, 32'h4057ed94} /* (24, 30, 3) {real, imag} */,
  {32'h42052300, 32'h40ae2f34} /* (24, 30, 2) {real, imag} */,
  {32'h4220b839, 32'h41c6d656} /* (24, 30, 1) {real, imag} */,
  {32'h41485167, 32'h419cf720} /* (24, 30, 0) {real, imag} */,
  {32'hc00e0d9e, 32'h409bc08a} /* (24, 29, 31) {real, imag} */,
  {32'hbfa1feba, 32'h416630a0} /* (24, 29, 30) {real, imag} */,
  {32'hbdc995c0, 32'h412e05f4} /* (24, 29, 29) {real, imag} */,
  {32'hc11018b5, 32'hc091274f} /* (24, 29, 28) {real, imag} */,
  {32'hc0f5c4bb, 32'h405fff74} /* (24, 29, 27) {real, imag} */,
  {32'hc0a38e4e, 32'hbfb62d2f} /* (24, 29, 26) {real, imag} */,
  {32'hc1a5b83f, 32'hc0268188} /* (24, 29, 25) {real, imag} */,
  {32'h411ab858, 32'h40f3609e} /* (24, 29, 24) {real, imag} */,
  {32'h4143d964, 32'h4184653c} /* (24, 29, 23) {real, imag} */,
  {32'hc110f420, 32'h40722948} /* (24, 29, 22) {real, imag} */,
  {32'hbfcf59e0, 32'hc144f4a3} /* (24, 29, 21) {real, imag} */,
  {32'h41945cde, 32'hc156aaea} /* (24, 29, 20) {real, imag} */,
  {32'h41e11a84, 32'h40332c3a} /* (24, 29, 19) {real, imag} */,
  {32'h411660ae, 32'hc193ee50} /* (24, 29, 18) {real, imag} */,
  {32'hbffd99b8, 32'hc1366f14} /* (24, 29, 17) {real, imag} */,
  {32'h415131e9, 32'hc11ae5ab} /* (24, 29, 16) {real, imag} */,
  {32'hbf3d1e2c, 32'h40226870} /* (24, 29, 15) {real, imag} */,
  {32'h3fbb62ac, 32'h4017799a} /* (24, 29, 14) {real, imag} */,
  {32'h3f8a10e4, 32'h414e646f} /* (24, 29, 13) {real, imag} */,
  {32'h4050d81c, 32'h412aab44} /* (24, 29, 12) {real, imag} */,
  {32'h4080ccd5, 32'h3fa130e6} /* (24, 29, 11) {real, imag} */,
  {32'h3f8c8526, 32'hc032933e} /* (24, 29, 10) {real, imag} */,
  {32'hc15a23e7, 32'hbeb19654} /* (24, 29, 9) {real, imag} */,
  {32'hc1c6e2b4, 32'h41357684} /* (24, 29, 8) {real, imag} */,
  {32'hc17f04f6, 32'h40e1ddf0} /* (24, 29, 7) {real, imag} */,
  {32'hc12aa348, 32'h40722c98} /* (24, 29, 6) {real, imag} */,
  {32'hc1e1810f, 32'h412b901c} /* (24, 29, 5) {real, imag} */,
  {32'hc1a118fe, 32'h40dc7054} /* (24, 29, 4) {real, imag} */,
  {32'h4112d3cf, 32'h409bda9b} /* (24, 29, 3) {real, imag} */,
  {32'hc02b6cc7, 32'hbf4de4bc} /* (24, 29, 2) {real, imag} */,
  {32'h3e428de0, 32'hbf9e2225} /* (24, 29, 1) {real, imag} */,
  {32'hbff0c0b3, 32'h401922b0} /* (24, 29, 0) {real, imag} */,
  {32'hbffb501d, 32'h3f98c608} /* (24, 28, 31) {real, imag} */,
  {32'hbfb5c300, 32'hc0ef1f2e} /* (24, 28, 30) {real, imag} */,
  {32'hc0292be6, 32'hc108603e} /* (24, 28, 29) {real, imag} */,
  {32'hc096a9d8, 32'h3f6e8d58} /* (24, 28, 28) {real, imag} */,
  {32'hc0967b98, 32'hc1291af3} /* (24, 28, 27) {real, imag} */,
  {32'hbf8e52dc, 32'hc00db913} /* (24, 28, 26) {real, imag} */,
  {32'hc15fdae0, 32'hbf640b58} /* (24, 28, 25) {real, imag} */,
  {32'hc0ada2e6, 32'h406883f8} /* (24, 28, 24) {real, imag} */,
  {32'hc1826e03, 32'h3f1e1a78} /* (24, 28, 23) {real, imag} */,
  {32'hc1592050, 32'hc18a4425} /* (24, 28, 22) {real, imag} */,
  {32'h413a3165, 32'hc0f21fdd} /* (24, 28, 21) {real, imag} */,
  {32'h41e67186, 32'h4045e92a} /* (24, 28, 20) {real, imag} */,
  {32'h419a8884, 32'hbec8fc54} /* (24, 28, 19) {real, imag} */,
  {32'h41c39719, 32'hc10bd44e} /* (24, 28, 18) {real, imag} */,
  {32'h41e69496, 32'hc0a804c4} /* (24, 28, 17) {real, imag} */,
  {32'h41cd7cba, 32'h4193a0cc} /* (24, 28, 16) {real, imag} */,
  {32'hc03dc0b3, 32'h41b24a47} /* (24, 28, 15) {real, imag} */,
  {32'hc083060e, 32'hc08543e8} /* (24, 28, 14) {real, imag} */,
  {32'h411d2a09, 32'hc137a93c} /* (24, 28, 13) {real, imag} */,
  {32'h415484ac, 32'hbeacdce0} /* (24, 28, 12) {real, imag} */,
  {32'hc0b666b4, 32'h40485ee4} /* (24, 28, 11) {real, imag} */,
  {32'hc10962dc, 32'h418165af} /* (24, 28, 10) {real, imag} */,
  {32'hc090d050, 32'h405590d7} /* (24, 28, 9) {real, imag} */,
  {32'hc1a12206, 32'hc07feeb4} /* (24, 28, 8) {real, imag} */,
  {32'hc1b1dce4, 32'hc087bd1b} /* (24, 28, 7) {real, imag} */,
  {32'hc1cf7dba, 32'h4112e52c} /* (24, 28, 6) {real, imag} */,
  {32'hc1a3dcf8, 32'h40ac37a8} /* (24, 28, 5) {real, imag} */,
  {32'hc1199b2f, 32'h3fce5390} /* (24, 28, 4) {real, imag} */,
  {32'hc1094e54, 32'hc00975b8} /* (24, 28, 3) {real, imag} */,
  {32'h40070140, 32'hc11ff2b6} /* (24, 28, 2) {real, imag} */,
  {32'h40ee86e8, 32'h41942f54} /* (24, 28, 1) {real, imag} */,
  {32'h4097d20c, 32'h4181fa65} /* (24, 28, 0) {real, imag} */,
  {32'h416fc05a, 32'h3f0cefc8} /* (24, 27, 31) {real, imag} */,
  {32'h416bcaea, 32'h40b5fe02} /* (24, 27, 30) {real, imag} */,
  {32'hc0844d9a, 32'h419c40c9} /* (24, 27, 29) {real, imag} */,
  {32'hbf082138, 32'h4163377b} /* (24, 27, 28) {real, imag} */,
  {32'h40d73eae, 32'h3f0e6f60} /* (24, 27, 27) {real, imag} */,
  {32'h4192ab5d, 32'hc097aada} /* (24, 27, 26) {real, imag} */,
  {32'h4165df89, 32'hbfa231d6} /* (24, 27, 25) {real, imag} */,
  {32'h41aa95a0, 32'hc0dcb010} /* (24, 27, 24) {real, imag} */,
  {32'h41fa97c3, 32'h40f6607a} /* (24, 27, 23) {real, imag} */,
  {32'h416a2e7d, 32'h3f9a14c8} /* (24, 27, 22) {real, imag} */,
  {32'h4171a3e4, 32'h400b6a5c} /* (24, 27, 21) {real, imag} */,
  {32'h40ed2ab4, 32'hbf90aec3} /* (24, 27, 20) {real, imag} */,
  {32'h4016d8f8, 32'hc06e9b65} /* (24, 27, 19) {real, imag} */,
  {32'hbf6bc3ac, 32'hbd88a560} /* (24, 27, 18) {real, imag} */,
  {32'hc0821a1f, 32'h3ff66c9d} /* (24, 27, 17) {real, imag} */,
  {32'hc11509b0, 32'hc0d74050} /* (24, 27, 16) {real, imag} */,
  {32'hc116be1f, 32'hc0ff1118} /* (24, 27, 15) {real, imag} */,
  {32'hc0401a34, 32'hc0b500de} /* (24, 27, 14) {real, imag} */,
  {32'hbfc1d153, 32'hc0d0567e} /* (24, 27, 13) {real, imag} */,
  {32'hc1011cbe, 32'h411a766a} /* (24, 27, 12) {real, imag} */,
  {32'hc13d0b2e, 32'h4137deaf} /* (24, 27, 11) {real, imag} */,
  {32'hc0ffae0a, 32'h40da45ed} /* (24, 27, 10) {real, imag} */,
  {32'hc0455f8e, 32'h40259fc2} /* (24, 27, 9) {real, imag} */,
  {32'h4130d43b, 32'h405d6c76} /* (24, 27, 8) {real, imag} */,
  {32'h413d122a, 32'hc0c97e68} /* (24, 27, 7) {real, imag} */,
  {32'h4136c385, 32'hc00590c6} /* (24, 27, 6) {real, imag} */,
  {32'h40649321, 32'h4162168e} /* (24, 27, 5) {real, imag} */,
  {32'h4098f022, 32'h40cd3ed8} /* (24, 27, 4) {real, imag} */,
  {32'h406c59d8, 32'h40bca82a} /* (24, 27, 3) {real, imag} */,
  {32'hc0660d1a, 32'h4144918e} /* (24, 27, 2) {real, imag} */,
  {32'h4152fa75, 32'h40c0bbdf} /* (24, 27, 1) {real, imag} */,
  {32'h41a60722, 32'h3fb5c6fa} /* (24, 27, 0) {real, imag} */,
  {32'h4035e45e, 32'hc10abf44} /* (24, 26, 31) {real, imag} */,
  {32'h41413ef3, 32'hc0975ff6} /* (24, 26, 30) {real, imag} */,
  {32'h41734d44, 32'h408d64a2} /* (24, 26, 29) {real, imag} */,
  {32'h40ba24ba, 32'h3ecbf8b8} /* (24, 26, 28) {real, imag} */,
  {32'hbfc1fe3c, 32'hc0fbc006} /* (24, 26, 27) {real, imag} */,
  {32'h4042fe3e, 32'hc0cbd6a2} /* (24, 26, 26) {real, imag} */,
  {32'hc0a17528, 32'h40dd53c2} /* (24, 26, 25) {real, imag} */,
  {32'hc1651556, 32'h4183c64e} /* (24, 26, 24) {real, imag} */,
  {32'hc1268afb, 32'h3fc16928} /* (24, 26, 23) {real, imag} */,
  {32'hbfb1e91b, 32'h3fccf4b8} /* (24, 26, 22) {real, imag} */,
  {32'h4057577e, 32'h40aaef01} /* (24, 26, 21) {real, imag} */,
  {32'h4045fa85, 32'h40b9a3da} /* (24, 26, 20) {real, imag} */,
  {32'h41300e1e, 32'hc0fb1bd1} /* (24, 26, 19) {real, imag} */,
  {32'h40c620d7, 32'hc1062d19} /* (24, 26, 18) {real, imag} */,
  {32'hc0a968d0, 32'hc0304864} /* (24, 26, 17) {real, imag} */,
  {32'hc1422c66, 32'h4105baf4} /* (24, 26, 16) {real, imag} */,
  {32'hc0e15b02, 32'h4006e91f} /* (24, 26, 15) {real, imag} */,
  {32'hc1131ede, 32'h3e9b8c80} /* (24, 26, 14) {real, imag} */,
  {32'hc0f45c07, 32'h3ebd6140} /* (24, 26, 13) {real, imag} */,
  {32'hc19d9c10, 32'h40a7a12c} /* (24, 26, 12) {real, imag} */,
  {32'hc0c77216, 32'h41735a8c} /* (24, 26, 11) {real, imag} */,
  {32'hc10d30b4, 32'h40a2398d} /* (24, 26, 10) {real, imag} */,
  {32'h4073d4bd, 32'hc12a8a9e} /* (24, 26, 9) {real, imag} */,
  {32'h40ebcb9c, 32'hc0a8783e} /* (24, 26, 8) {real, imag} */,
  {32'hc08c07e1, 32'h40a9d324} /* (24, 26, 7) {real, imag} */,
  {32'hc10e49d2, 32'h4095c59c} /* (24, 26, 6) {real, imag} */,
  {32'h3e01f000, 32'h41a9ef91} /* (24, 26, 5) {real, imag} */,
  {32'h4099b980, 32'h412caf5c} /* (24, 26, 4) {real, imag} */,
  {32'h401470d1, 32'h3f9c0f4d} /* (24, 26, 3) {real, imag} */,
  {32'h412e6732, 32'h400df2fc} /* (24, 26, 2) {real, imag} */,
  {32'h41215464, 32'h40db37a4} /* (24, 26, 1) {real, imag} */,
  {32'h4102ce3d, 32'h40fbcaa8} /* (24, 26, 0) {real, imag} */,
  {32'h3f4f64c4, 32'h3f8e4d4a} /* (24, 25, 31) {real, imag} */,
  {32'h409cac15, 32'h40d5b532} /* (24, 25, 30) {real, imag} */,
  {32'h3ffcb12e, 32'h4123d92a} /* (24, 25, 29) {real, imag} */,
  {32'hbfa96b45, 32'h4108c84f} /* (24, 25, 28) {real, imag} */,
  {32'hbdd92b80, 32'h4084169a} /* (24, 25, 27) {real, imag} */,
  {32'h402b5184, 32'h40881cc1} /* (24, 25, 26) {real, imag} */,
  {32'hbe5f84c0, 32'h40fb0ea5} /* (24, 25, 25) {real, imag} */,
  {32'hc0635212, 32'hc023cc9c} /* (24, 25, 24) {real, imag} */,
  {32'hc099e7d2, 32'h3f0d6920} /* (24, 25, 23) {real, imag} */,
  {32'hc107f919, 32'h3e0037c0} /* (24, 25, 22) {real, imag} */,
  {32'hc11ac91e, 32'hc1240961} /* (24, 25, 21) {real, imag} */,
  {32'h3e0c4830, 32'hc077e46f} /* (24, 25, 20) {real, imag} */,
  {32'h40d31794, 32'hc113f60f} /* (24, 25, 19) {real, imag} */,
  {32'h41190366, 32'hc0894235} /* (24, 25, 18) {real, imag} */,
  {32'hc0257ae6, 32'h3fe10184} /* (24, 25, 17) {real, imag} */,
  {32'h4122b376, 32'hc0afb32d} /* (24, 25, 16) {real, imag} */,
  {32'h4152d80e, 32'hc168b85a} /* (24, 25, 15) {real, imag} */,
  {32'h40152758, 32'hc14df50d} /* (24, 25, 14) {real, imag} */,
  {32'h3f57acb4, 32'hc1598d6e} /* (24, 25, 13) {real, imag} */,
  {32'hbf0d7314, 32'hc14ee014} /* (24, 25, 12) {real, imag} */,
  {32'h40b30a2e, 32'h4087c982} /* (24, 25, 11) {real, imag} */,
  {32'hbe45a500, 32'hc0b2cdec} /* (24, 25, 10) {real, imag} */,
  {32'h40535c41, 32'hc1b9d7b0} /* (24, 25, 9) {real, imag} */,
  {32'h404d7c7e, 32'hc18b889b} /* (24, 25, 8) {real, imag} */,
  {32'h41631fd0, 32'hc0a544a5} /* (24, 25, 7) {real, imag} */,
  {32'h41637206, 32'hbf274828} /* (24, 25, 6) {real, imag} */,
  {32'h405ce4bc, 32'hbe9df8a0} /* (24, 25, 5) {real, imag} */,
  {32'h40d44536, 32'hc047db1a} /* (24, 25, 4) {real, imag} */,
  {32'h4012103e, 32'h40b1409e} /* (24, 25, 3) {real, imag} */,
  {32'hc10994a3, 32'h40f5fc78} /* (24, 25, 2) {real, imag} */,
  {32'hc15be6e4, 32'hbf544e98} /* (24, 25, 1) {real, imag} */,
  {32'hc0911e94, 32'hc0aa33e2} /* (24, 25, 0) {real, imag} */,
  {32'h40b8c350, 32'h411247a5} /* (24, 24, 31) {real, imag} */,
  {32'h4010431c, 32'hc14c907f} /* (24, 24, 30) {real, imag} */,
  {32'hbfce8650, 32'hc1e50080} /* (24, 24, 29) {real, imag} */,
  {32'hc0ad7737, 32'hc153cc9e} /* (24, 24, 28) {real, imag} */,
  {32'h3fd5344c, 32'hc155f1a2} /* (24, 24, 27) {real, imag} */,
  {32'h416547ca, 32'hc1793c26} /* (24, 24, 26) {real, imag} */,
  {32'h416d9b23, 32'h401fbaf0} /* (24, 24, 25) {real, imag} */,
  {32'h410700b5, 32'h41a7aa35} /* (24, 24, 24) {real, imag} */,
  {32'h40385566, 32'h3fc11ea5} /* (24, 24, 23) {real, imag} */,
  {32'h414b5562, 32'h3fa39cd8} /* (24, 24, 22) {real, imag} */,
  {32'h40bbcefd, 32'h413b0079} /* (24, 24, 21) {real, imag} */,
  {32'hc05b71a3, 32'hbdb757c0} /* (24, 24, 20) {real, imag} */,
  {32'hc0c51a69, 32'hc05da0d8} /* (24, 24, 19) {real, imag} */,
  {32'h3fa4ddf8, 32'h409d33fc} /* (24, 24, 18) {real, imag} */,
  {32'h3f7d0244, 32'h3fa10fbc} /* (24, 24, 17) {real, imag} */,
  {32'hc0512435, 32'hc06def84} /* (24, 24, 16) {real, imag} */,
  {32'hc10ca20a, 32'h40501e14} /* (24, 24, 15) {real, imag} */,
  {32'hc133915a, 32'hc0a4fb9e} /* (24, 24, 14) {real, imag} */,
  {32'hc0dac662, 32'hc179928a} /* (24, 24, 13) {real, imag} */,
  {32'hc124db7f, 32'hc0eab084} /* (24, 24, 12) {real, imag} */,
  {32'hc02a04f2, 32'hc0de771f} /* (24, 24, 11) {real, imag} */,
  {32'h40c968df, 32'h4120702e} /* (24, 24, 10) {real, imag} */,
  {32'h4119d258, 32'h3e3286c0} /* (24, 24, 9) {real, imag} */,
  {32'h41358475, 32'h40c86173} /* (24, 24, 8) {real, imag} */,
  {32'h413f51b9, 32'h403b1a9e} /* (24, 24, 7) {real, imag} */,
  {32'h40ac8217, 32'h4098617e} /* (24, 24, 6) {real, imag} */,
  {32'hc11b77c7, 32'h404ce56c} /* (24, 24, 5) {real, imag} */,
  {32'h400c7a5d, 32'h40aee4a2} /* (24, 24, 4) {real, imag} */,
  {32'h3e819030, 32'hbfe5bb88} /* (24, 24, 3) {real, imag} */,
  {32'h3fae9838, 32'hc00a1c3c} /* (24, 24, 2) {real, imag} */,
  {32'h4086274c, 32'h411dd363} /* (24, 24, 1) {real, imag} */,
  {32'h40b1d973, 32'h4181d3b6} /* (24, 24, 0) {real, imag} */,
  {32'hc0dacb94, 32'h40dff0c2} /* (24, 23, 31) {real, imag} */,
  {32'hbfcae114, 32'h40c229ca} /* (24, 23, 30) {real, imag} */,
  {32'hbf03144c, 32'h411f45dc} /* (24, 23, 29) {real, imag} */,
  {32'h405c803a, 32'h4084973e} /* (24, 23, 28) {real, imag} */,
  {32'h3fbf4148, 32'hc06a186c} /* (24, 23, 27) {real, imag} */,
  {32'hc10470c1, 32'hc044aaaa} /* (24, 23, 26) {real, imag} */,
  {32'hc065bcd0, 32'hc0e05830} /* (24, 23, 25) {real, imag} */,
  {32'hbf01ed8c, 32'hc0500c6e} /* (24, 23, 24) {real, imag} */,
  {32'h3e9825e0, 32'h4078c00c} /* (24, 23, 23) {real, imag} */,
  {32'h40a83ec4, 32'h4046a388} /* (24, 23, 22) {real, imag} */,
  {32'h40fca6e6, 32'h401856d3} /* (24, 23, 21) {real, imag} */,
  {32'h4010f6ec, 32'h40904d00} /* (24, 23, 20) {real, imag} */,
  {32'hc0580812, 32'h401810e3} /* (24, 23, 19) {real, imag} */,
  {32'hc10e8ffe, 32'h40b94711} /* (24, 23, 18) {real, imag} */,
  {32'hc082f3c4, 32'hc0c20c56} /* (24, 23, 17) {real, imag} */,
  {32'hc0ba9104, 32'hc0a8bc0d} /* (24, 23, 16) {real, imag} */,
  {32'hbf2d1e24, 32'hbf138340} /* (24, 23, 15) {real, imag} */,
  {32'h3fc225d0, 32'h3ff6e2cc} /* (24, 23, 14) {real, imag} */,
  {32'h418d21ae, 32'hc0285bb0} /* (24, 23, 13) {real, imag} */,
  {32'h40d0aac6, 32'h40496a63} /* (24, 23, 12) {real, imag} */,
  {32'hbffe9118, 32'h40649c88} /* (24, 23, 11) {real, imag} */,
  {32'h4002e5c2, 32'hc0734bc4} /* (24, 23, 10) {real, imag} */,
  {32'hc0d60b86, 32'h3ea98f90} /* (24, 23, 9) {real, imag} */,
  {32'hc08c29b4, 32'h4051796e} /* (24, 23, 8) {real, imag} */,
  {32'hc109fa5c, 32'hbe7c0ce0} /* (24, 23, 7) {real, imag} */,
  {32'hc0981b49, 32'hc0924c7e} /* (24, 23, 6) {real, imag} */,
  {32'hc089735c, 32'hc0b3dad2} /* (24, 23, 5) {real, imag} */,
  {32'hc1340ba1, 32'hbf664356} /* (24, 23, 4) {real, imag} */,
  {32'hc0a0ff2d, 32'hbf05b0c0} /* (24, 23, 3) {real, imag} */,
  {32'hc07691b5, 32'h40f7a1b2} /* (24, 23, 2) {real, imag} */,
  {32'hc11247f2, 32'h410c7a06} /* (24, 23, 1) {real, imag} */,
  {32'hc04a3284, 32'h4052192a} /* (24, 23, 0) {real, imag} */,
  {32'hc0b8a6e3, 32'h3f279f6c} /* (24, 22, 31) {real, imag} */,
  {32'hc06e1d96, 32'hc00d9c7f} /* (24, 22, 30) {real, imag} */,
  {32'h3ef68a8c, 32'hbf9e7b20} /* (24, 22, 29) {real, imag} */,
  {32'hbf40097c, 32'h40f0ef5a} /* (24, 22, 28) {real, imag} */,
  {32'hbf95ec52, 32'h4017290f} /* (24, 22, 27) {real, imag} */,
  {32'h3e093790, 32'h407fb048} /* (24, 22, 26) {real, imag} */,
  {32'hbf0a0880, 32'h40a144d6} /* (24, 22, 25) {real, imag} */,
  {32'h3f8b4606, 32'h403bfff5} /* (24, 22, 24) {real, imag} */,
  {32'h4033bb38, 32'h40380cf4} /* (24, 22, 23) {real, imag} */,
  {32'hbf952a39, 32'h3f533df0} /* (24, 22, 22) {real, imag} */,
  {32'hc0644bee, 32'h4035aaea} /* (24, 22, 21) {real, imag} */,
  {32'h409e94da, 32'hc0abb93c} /* (24, 22, 20) {real, imag} */,
  {32'h40f9004c, 32'hc0b7cc71} /* (24, 22, 19) {real, imag} */,
  {32'h40ccf593, 32'hc06a5ec5} /* (24, 22, 18) {real, imag} */,
  {32'h4102e0c5, 32'hc0473a8a} /* (24, 22, 17) {real, imag} */,
  {32'h3f421e26, 32'hc057a1b9} /* (24, 22, 16) {real, imag} */,
  {32'h4008d877, 32'hc0926295} /* (24, 22, 15) {real, imag} */,
  {32'hbf48c618, 32'h3f86aba2} /* (24, 22, 14) {real, imag} */,
  {32'h3ef395b8, 32'h40ad0e97} /* (24, 22, 13) {real, imag} */,
  {32'hbfa81c50, 32'h4004a8f8} /* (24, 22, 12) {real, imag} */,
  {32'hc0ac96d0, 32'hbe1e9900} /* (24, 22, 11) {real, imag} */,
  {32'hc0d3760c, 32'h3e31a820} /* (24, 22, 10) {real, imag} */,
  {32'hc1155fa3, 32'h3d873dc0} /* (24, 22, 9) {real, imag} */,
  {32'hc141170e, 32'hc0c055c4} /* (24, 22, 8) {real, imag} */,
  {32'hc0c16f87, 32'hc0a9d41c} /* (24, 22, 7) {real, imag} */,
  {32'hbfd4bf02, 32'h4087c52e} /* (24, 22, 6) {real, imag} */,
  {32'hc0c635c0, 32'hbecd7ea0} /* (24, 22, 5) {real, imag} */,
  {32'hc07f9347, 32'hbfd2b27b} /* (24, 22, 4) {real, imag} */,
  {32'hbedb29b0, 32'hbfb9ae44} /* (24, 22, 3) {real, imag} */,
  {32'hbf342418, 32'hc032b28c} /* (24, 22, 2) {real, imag} */,
  {32'hc07bde91, 32'h3f025ea8} /* (24, 22, 1) {real, imag} */,
  {32'hc043d8c9, 32'h402ae403} /* (24, 22, 0) {real, imag} */,
  {32'h40945616, 32'hbfe71526} /* (24, 21, 31) {real, imag} */,
  {32'h408c21aa, 32'hbfbc2724} /* (24, 21, 30) {real, imag} */,
  {32'hc0040d5d, 32'hc109cdec} /* (24, 21, 29) {real, imag} */,
  {32'hc04c9290, 32'hc111d161} /* (24, 21, 28) {real, imag} */,
  {32'hc0c4c1fe, 32'hc0e9be5a} /* (24, 21, 27) {real, imag} */,
  {32'h3ea8efc0, 32'hc13e009e} /* (24, 21, 26) {real, imag} */,
  {32'h40bd7ff2, 32'hbfb83386} /* (24, 21, 25) {real, imag} */,
  {32'h400781ae, 32'hc063ff2b} /* (24, 21, 24) {real, imag} */,
  {32'h404d3aa2, 32'hc083a80e} /* (24, 21, 23) {real, imag} */,
  {32'h40f5ed10, 32'hc089d836} /* (24, 21, 22) {real, imag} */,
  {32'h40cda4d8, 32'hbf5c1e38} /* (24, 21, 21) {real, imag} */,
  {32'hc0be6684, 32'h400b9e2a} /* (24, 21, 20) {real, imag} */,
  {32'hc119671b, 32'hc03eed92} /* (24, 21, 19) {real, imag} */,
  {32'hc0647b24, 32'h3fb42e42} /* (24, 21, 18) {real, imag} */,
  {32'h40860bca, 32'h408797e2} /* (24, 21, 17) {real, imag} */,
  {32'h400c128a, 32'h3f5bb9e0} /* (24, 21, 16) {real, imag} */,
  {32'hc0aabedc, 32'hbebfcb90} /* (24, 21, 15) {real, imag} */,
  {32'hc09b3922, 32'h40757630} /* (24, 21, 14) {real, imag} */,
  {32'hc0ccfea4, 32'hbe092490} /* (24, 21, 13) {real, imag} */,
  {32'h3f3435e4, 32'hc0db7ec6} /* (24, 21, 12) {real, imag} */,
  {32'h3fa92adc, 32'hc052cbce} /* (24, 21, 11) {real, imag} */,
  {32'hbe910b78, 32'h3e61a790} /* (24, 21, 10) {real, imag} */,
  {32'hc0051157, 32'hc02e54e9} /* (24, 21, 9) {real, imag} */,
  {32'hbee9e4d8, 32'h401a0b9a} /* (24, 21, 8) {real, imag} */,
  {32'h3f74a4a0, 32'h4098d07c} /* (24, 21, 7) {real, imag} */,
  {32'h40bf5812, 32'hbfc4aef6} /* (24, 21, 6) {real, imag} */,
  {32'h40f72770, 32'hc02b32c4} /* (24, 21, 5) {real, imag} */,
  {32'h40a8c416, 32'hc03628fe} /* (24, 21, 4) {real, imag} */,
  {32'h40b90226, 32'hc0ca88b3} /* (24, 21, 3) {real, imag} */,
  {32'h40b2bdb6, 32'hc0237185} /* (24, 21, 2) {real, imag} */,
  {32'h40d37128, 32'h40b3a8fd} /* (24, 21, 1) {real, imag} */,
  {32'h4001b279, 32'h3fa4b0c2} /* (24, 21, 0) {real, imag} */,
  {32'h403e3ac4, 32'h3fc73a16} /* (24, 20, 31) {real, imag} */,
  {32'hc049e7a7, 32'h4081ebf0} /* (24, 20, 30) {real, imag} */,
  {32'hc0a8cd47, 32'hc01b1cdd} /* (24, 20, 29) {real, imag} */,
  {32'h4060a6ae, 32'hc1071402} /* (24, 20, 28) {real, imag} */,
  {32'h3fbcd090, 32'hc08ce835} /* (24, 20, 27) {real, imag} */,
  {32'hbf4f2958, 32'h402aaf3f} /* (24, 20, 26) {real, imag} */,
  {32'hc0a40770, 32'h3fef1091} /* (24, 20, 25) {real, imag} */,
  {32'h3f24e021, 32'hc0bed398} /* (24, 20, 24) {real, imag} */,
  {32'h3ff39034, 32'hc09f5e9f} /* (24, 20, 23) {real, imag} */,
  {32'h4057b61d, 32'hc08d4d66} /* (24, 20, 22) {real, imag} */,
  {32'hc0cace44, 32'h3d35cc40} /* (24, 20, 21) {real, imag} */,
  {32'hc062a5f2, 32'h40339827} /* (24, 20, 20) {real, imag} */,
  {32'hc02fa61e, 32'h3f83e9e7} /* (24, 20, 19) {real, imag} */,
  {32'hc02a57c8, 32'h40712631} /* (24, 20, 18) {real, imag} */,
  {32'hc02a77f6, 32'h40cd542b} /* (24, 20, 17) {real, imag} */,
  {32'hbfb45410, 32'hbf47eb74} /* (24, 20, 16) {real, imag} */,
  {32'h40927f8c, 32'hbfd32218} /* (24, 20, 15) {real, imag} */,
  {32'h40a025ec, 32'hbd712e00} /* (24, 20, 14) {real, imag} */,
  {32'h411502fb, 32'h406d4145} /* (24, 20, 13) {real, imag} */,
  {32'h40b8c94b, 32'hc09c24da} /* (24, 20, 12) {real, imag} */,
  {32'h3f8fff00, 32'hbf7253d6} /* (24, 20, 11) {real, imag} */,
  {32'hc0de9623, 32'h3b52f800} /* (24, 20, 10) {real, imag} */,
  {32'hc0aadf76, 32'hc002fd53} /* (24, 20, 9) {real, imag} */,
  {32'h409e9fa3, 32'hbf950806} /* (24, 20, 8) {real, imag} */,
  {32'h40810271, 32'h4010312e} /* (24, 20, 7) {real, imag} */,
  {32'h3efa2650, 32'hbef89bd0} /* (24, 20, 6) {real, imag} */,
  {32'h40398f78, 32'hc0339e99} /* (24, 20, 5) {real, imag} */,
  {32'h3f9d5376, 32'hc093786e} /* (24, 20, 4) {real, imag} */,
  {32'h3dfa5bf0, 32'hbfe698ed} /* (24, 20, 3) {real, imag} */,
  {32'hc041d740, 32'hbfe4e197} /* (24, 20, 2) {real, imag} */,
  {32'hc0e19584, 32'hbffb1201} /* (24, 20, 1) {real, imag} */,
  {32'hc006b0cd, 32'h405ad1d4} /* (24, 20, 0) {real, imag} */,
  {32'hc04e89c2, 32'h3efdcb74} /* (24, 19, 31) {real, imag} */,
  {32'hc028b22f, 32'h3f119360} /* (24, 19, 30) {real, imag} */,
  {32'hc02dc2ab, 32'hbff33500} /* (24, 19, 29) {real, imag} */,
  {32'hbfc51aea, 32'hbf9b939c} /* (24, 19, 28) {real, imag} */,
  {32'hc006d35e, 32'h40151869} /* (24, 19, 27) {real, imag} */,
  {32'h3fb4047e, 32'h3fcffc8c} /* (24, 19, 26) {real, imag} */,
  {32'h40a67780, 32'hbfe1821c} /* (24, 19, 25) {real, imag} */,
  {32'h40000b3a, 32'h40a1cd94} /* (24, 19, 24) {real, imag} */,
  {32'hbf851bc6, 32'h4087769e} /* (24, 19, 23) {real, imag} */,
  {32'hc05047fd, 32'hc08100cb} /* (24, 19, 22) {real, imag} */,
  {32'hbfa5bc20, 32'hbe72e730} /* (24, 19, 21) {real, imag} */,
  {32'hbfaf1338, 32'h3d438c00} /* (24, 19, 20) {real, imag} */,
  {32'h407d8c50, 32'h4029180d} /* (24, 19, 19) {real, imag} */,
  {32'h402d6535, 32'h4063ba0c} /* (24, 19, 18) {real, imag} */,
  {32'hbec3aa88, 32'h409c101c} /* (24, 19, 17) {real, imag} */,
  {32'h40321862, 32'h410d2ca8} /* (24, 19, 16) {real, imag} */,
  {32'h3f862f27, 32'h4109341c} /* (24, 19, 15) {real, imag} */,
  {32'hc02857d2, 32'h4091dea5} /* (24, 19, 14) {real, imag} */,
  {32'h3f9785cf, 32'h40745179} /* (24, 19, 13) {real, imag} */,
  {32'h3f345ea4, 32'h40498062} /* (24, 19, 12) {real, imag} */,
  {32'h40a8ba69, 32'hbf951cca} /* (24, 19, 11) {real, imag} */,
  {32'h405081f3, 32'hbf773540} /* (24, 19, 10) {real, imag} */,
  {32'h3f660e2c, 32'h403fd0bc} /* (24, 19, 9) {real, imag} */,
  {32'hbf919a44, 32'hc0503286} /* (24, 19, 8) {real, imag} */,
  {32'hbfc201ea, 32'hbfb64a6c} /* (24, 19, 7) {real, imag} */,
  {32'hc0112aee, 32'hbfa31f38} /* (24, 19, 6) {real, imag} */,
  {32'h3fd7cf48, 32'hc0b6ec0c} /* (24, 19, 5) {real, imag} */,
  {32'hc01aecee, 32'hbfcba786} /* (24, 19, 4) {real, imag} */,
  {32'hc0331cac, 32'h411296da} /* (24, 19, 3) {real, imag} */,
  {32'hbf6320f2, 32'h4059721f} /* (24, 19, 2) {real, imag} */,
  {32'h3fc3ef37, 32'hc0732477} /* (24, 19, 1) {real, imag} */,
  {32'h3f85cfee, 32'hbf803a46} /* (24, 19, 0) {real, imag} */,
  {32'hbeb574a8, 32'h3cbfb600} /* (24, 18, 31) {real, imag} */,
  {32'h3fdc6552, 32'hbf6cdb30} /* (24, 18, 30) {real, imag} */,
  {32'h40d70adf, 32'hbfb8122f} /* (24, 18, 29) {real, imag} */,
  {32'h40280be2, 32'hbea740c0} /* (24, 18, 28) {real, imag} */,
  {32'hbffd1e80, 32'hc068c4cf} /* (24, 18, 27) {real, imag} */,
  {32'hc06ef72a, 32'hbf88e6ff} /* (24, 18, 26) {real, imag} */,
  {32'h3fcdedba, 32'h4046e9a9} /* (24, 18, 25) {real, imag} */,
  {32'h400e7ec7, 32'h3e3d4258} /* (24, 18, 24) {real, imag} */,
  {32'h4010eabc, 32'hbf2c0fa0} /* (24, 18, 23) {real, imag} */,
  {32'h4052ed40, 32'h40950b54} /* (24, 18, 22) {real, imag} */,
  {32'hbfc2d898, 32'h40881b11} /* (24, 18, 21) {real, imag} */,
  {32'h3e84fb48, 32'h3f80b342} /* (24, 18, 20) {real, imag} */,
  {32'h3ef12ba0, 32'hbfc79baa} /* (24, 18, 19) {real, imag} */,
  {32'h407a636e, 32'hbff0ef11} /* (24, 18, 18) {real, imag} */,
  {32'hbff01434, 32'hc035066c} /* (24, 18, 17) {real, imag} */,
  {32'hc083d7cc, 32'h402964d8} /* (24, 18, 16) {real, imag} */,
  {32'hbfd5366a, 32'h40752f4e} /* (24, 18, 15) {real, imag} */,
  {32'h3f0a66e4, 32'h3f8be485} /* (24, 18, 14) {real, imag} */,
  {32'hbbd65600, 32'hbf0b5930} /* (24, 18, 13) {real, imag} */,
  {32'hbfb3e09a, 32'h3f3291dc} /* (24, 18, 12) {real, imag} */,
  {32'hbfcdff34, 32'hc03d8026} /* (24, 18, 11) {real, imag} */,
  {32'hc0964b65, 32'h3e66c490} /* (24, 18, 10) {real, imag} */,
  {32'h40082046, 32'h3f8333d6} /* (24, 18, 9) {real, imag} */,
  {32'h40112846, 32'h3fc0f8e9} /* (24, 18, 8) {real, imag} */,
  {32'h40a052fd, 32'h3e678c80} /* (24, 18, 7) {real, imag} */,
  {32'h40d32cbd, 32'hc0612e4c} /* (24, 18, 6) {real, imag} */,
  {32'h40b55024, 32'hc039edfe} /* (24, 18, 5) {real, imag} */,
  {32'hbfc4e2c8, 32'hc0287272} /* (24, 18, 4) {real, imag} */,
  {32'hc0a7216c, 32'hc0e2840e} /* (24, 18, 3) {real, imag} */,
  {32'hbf9f569a, 32'hc040bf74} /* (24, 18, 2) {real, imag} */,
  {32'h403792aa, 32'hbf5c5eec} /* (24, 18, 1) {real, imag} */,
  {32'h3f955f57, 32'hbe12f120} /* (24, 18, 0) {real, imag} */,
  {32'h402cad82, 32'hbf965bfe} /* (24, 17, 31) {real, imag} */,
  {32'h4020bab4, 32'hbffd13c4} /* (24, 17, 30) {real, imag} */,
  {32'hbeccc060, 32'h3fe4a458} /* (24, 17, 29) {real, imag} */,
  {32'h3ecc1180, 32'h3fcb76d4} /* (24, 17, 28) {real, imag} */,
  {32'h3f85f1e0, 32'h3fc1f46d} /* (24, 17, 27) {real, imag} */,
  {32'hbe8adb68, 32'h40113247} /* (24, 17, 26) {real, imag} */,
  {32'h3fb9053e, 32'h409314ac} /* (24, 17, 25) {real, imag} */,
  {32'h3fe80562, 32'h402ff35c} /* (24, 17, 24) {real, imag} */,
  {32'h40494ce8, 32'h3f8fa6cc} /* (24, 17, 23) {real, imag} */,
  {32'h4070a0f2, 32'h405d1e6e} /* (24, 17, 22) {real, imag} */,
  {32'h40223396, 32'h401a5712} /* (24, 17, 21) {real, imag} */,
  {32'h3db2e460, 32'h3f16d890} /* (24, 17, 20) {real, imag} */,
  {32'hbfa9a0ec, 32'h401e995f} /* (24, 17, 19) {real, imag} */,
  {32'hbf3eb240, 32'hbddf9c00} /* (24, 17, 18) {real, imag} */,
  {32'h40344178, 32'hc06627b4} /* (24, 17, 17) {real, imag} */,
  {32'h3fc811d0, 32'hc09b3507} /* (24, 17, 16) {real, imag} */,
  {32'h3f36a582, 32'hc0a0dae4} /* (24, 17, 15) {real, imag} */,
  {32'h3f080aee, 32'h3f284f2a} /* (24, 17, 14) {real, imag} */,
  {32'hc00c5e4b, 32'h400e36c0} /* (24, 17, 13) {real, imag} */,
  {32'h3f75d4b0, 32'h4019c1ac} /* (24, 17, 12) {real, imag} */,
  {32'h3f94c0f8, 32'h4020555f} /* (24, 17, 11) {real, imag} */,
  {32'hbfa37512, 32'h401b991a} /* (24, 17, 10) {real, imag} */,
  {32'hc008375a, 32'h4092243e} /* (24, 17, 9) {real, imag} */,
  {32'hc036264b, 32'h4036f62c} /* (24, 17, 8) {real, imag} */,
  {32'hc02eedfc, 32'hbf0bf038} /* (24, 17, 7) {real, imag} */,
  {32'hbfd50c40, 32'h3eed7358} /* (24, 17, 6) {real, imag} */,
  {32'hbf525f8c, 32'h3ff76fe4} /* (24, 17, 5) {real, imag} */,
  {32'h3ee681f0, 32'h4084b56e} /* (24, 17, 4) {real, imag} */,
  {32'h4019017e, 32'h40969fff} /* (24, 17, 3) {real, imag} */,
  {32'h3f5999d9, 32'h3ecc92e8} /* (24, 17, 2) {real, imag} */,
  {32'hbf194362, 32'h3e5ef0e8} /* (24, 17, 1) {real, imag} */,
  {32'hc001d0e2, 32'h3fa2d908} /* (24, 17, 0) {real, imag} */,
  {32'h3f5938e8, 32'h408e562e} /* (24, 16, 31) {real, imag} */,
  {32'h3ed579a0, 32'h40f03920} /* (24, 16, 30) {real, imag} */,
  {32'hc019c710, 32'h41065af1} /* (24, 16, 29) {real, imag} */,
  {32'hbfb44c58, 32'h40c520d8} /* (24, 16, 28) {real, imag} */,
  {32'hbfcca1c0, 32'h4080ebac} /* (24, 16, 27) {real, imag} */,
  {32'hbfc8a184, 32'h3eaefc10} /* (24, 16, 26) {real, imag} */,
  {32'hc016805f, 32'hbea7b9a0} /* (24, 16, 25) {real, imag} */,
  {32'h4059895a, 32'h401a3b73} /* (24, 16, 24) {real, imag} */,
  {32'h3f760130, 32'h3fd8efcf} /* (24, 16, 23) {real, imag} */,
  {32'hbe3bd200, 32'hbe51b240} /* (24, 16, 22) {real, imag} */,
  {32'h3e6461e0, 32'hbf996cc0} /* (24, 16, 21) {real, imag} */,
  {32'h3ffb85c6, 32'h3fd10b50} /* (24, 16, 20) {real, imag} */,
  {32'h405f7294, 32'h40881a7e} /* (24, 16, 19) {real, imag} */,
  {32'h400a02e7, 32'h408d7a20} /* (24, 16, 18) {real, imag} */,
  {32'hbfae1082, 32'h406c4b04} /* (24, 16, 17) {real, imag} */,
  {32'h3e886408, 32'h404bb336} /* (24, 16, 16) {real, imag} */,
  {32'h407fe954, 32'h3f1548d0} /* (24, 16, 15) {real, imag} */,
  {32'h3ee31d80, 32'h3de379c0} /* (24, 16, 14) {real, imag} */,
  {32'hbbcda800, 32'h401be2c8} /* (24, 16, 13) {real, imag} */,
  {32'h3f84bc90, 32'h401c80f6} /* (24, 16, 12) {real, imag} */,
  {32'h3f37cc30, 32'h405c190c} /* (24, 16, 11) {real, imag} */,
  {32'h3fad6298, 32'hc056ee1e} /* (24, 16, 10) {real, imag} */,
  {32'hbff80562, 32'hc09a304d} /* (24, 16, 9) {real, imag} */,
  {32'h3e7c8e60, 32'hbdb03e80} /* (24, 16, 8) {real, imag} */,
  {32'hbfd86a38, 32'h40b66e78} /* (24, 16, 7) {real, imag} */,
  {32'hbfe43510, 32'h40887ae4} /* (24, 16, 6) {real, imag} */,
  {32'h3f9abad2, 32'h3e491600} /* (24, 16, 5) {real, imag} */,
  {32'h3ecafa90, 32'h3d774400} /* (24, 16, 4) {real, imag} */,
  {32'hc09695a4, 32'hbfb37978} /* (24, 16, 3) {real, imag} */,
  {32'hc0b0860e, 32'hbfc9c050} /* (24, 16, 2) {real, imag} */,
  {32'hc0752c8c, 32'hc021f970} /* (24, 16, 1) {real, imag} */,
  {32'hbfc61290, 32'hbfb3fec8} /* (24, 16, 0) {real, imag} */,
  {32'hc06cb6a6, 32'h3ecda098} /* (24, 15, 31) {real, imag} */,
  {32'hbf841598, 32'h406c7d2a} /* (24, 15, 30) {real, imag} */,
  {32'h40140304, 32'hbe66f4c0} /* (24, 15, 29) {real, imag} */,
  {32'h40263c90, 32'hbf8c9e44} /* (24, 15, 28) {real, imag} */,
  {32'h3fa25ba0, 32'h3f1c6666} /* (24, 15, 27) {real, imag} */,
  {32'h4034673d, 32'hbe2ef2f0} /* (24, 15, 26) {real, imag} */,
  {32'h4010cc31, 32'h3e80afc0} /* (24, 15, 25) {real, imag} */,
  {32'hbffa81c2, 32'h409f3d66} /* (24, 15, 24) {real, imag} */,
  {32'hbf9bfe50, 32'h40147ada} /* (24, 15, 23) {real, imag} */,
  {32'h4036595e, 32'h3f52b0ca} /* (24, 15, 22) {real, imag} */,
  {32'h3e946ad0, 32'h3fe28bbc} /* (24, 15, 21) {real, imag} */,
  {32'hbfb5525a, 32'h3e22d840} /* (24, 15, 20) {real, imag} */,
  {32'hbf938c8c, 32'h3f87afe6} /* (24, 15, 19) {real, imag} */,
  {32'hbff55e30, 32'h3f8e9180} /* (24, 15, 18) {real, imag} */,
  {32'hbfeb5040, 32'hbf84d698} /* (24, 15, 17) {real, imag} */,
  {32'hc0108970, 32'hc072bcea} /* (24, 15, 16) {real, imag} */,
  {32'hbfa892a1, 32'hbfeeda32} /* (24, 15, 15) {real, imag} */,
  {32'h3f9efa79, 32'hbf25752a} /* (24, 15, 14) {real, imag} */,
  {32'h4049320b, 32'h402d7e38} /* (24, 15, 13) {real, imag} */,
  {32'hbe5781c0, 32'h3e5a1c48} /* (24, 15, 12) {real, imag} */,
  {32'hc0c3086e, 32'hc05b4fff} /* (24, 15, 11) {real, imag} */,
  {32'hc09805cc, 32'hbfb4784c} /* (24, 15, 10) {real, imag} */,
  {32'h3ed8a1b0, 32'hbfd4eba0} /* (24, 15, 9) {real, imag} */,
  {32'h3f6238d5, 32'hc019d444} /* (24, 15, 8) {real, imag} */,
  {32'h40102f9e, 32'hc0dc95dd} /* (24, 15, 7) {real, imag} */,
  {32'h3f66a9b0, 32'hc0ee17ee} /* (24, 15, 6) {real, imag} */,
  {32'h40284f83, 32'h3e7411e0} /* (24, 15, 5) {real, imag} */,
  {32'hbf141fd8, 32'h401322e5} /* (24, 15, 4) {real, imag} */,
  {32'hc057487e, 32'h3fd13845} /* (24, 15, 3) {real, imag} */,
  {32'h3cf888e0, 32'h40726933} /* (24, 15, 2) {real, imag} */,
  {32'h40572c40, 32'hc00ce1fe} /* (24, 15, 1) {real, imag} */,
  {32'hbd459980, 32'hc0610cc4} /* (24, 15, 0) {real, imag} */,
  {32'hc06a0759, 32'hbff3b510} /* (24, 14, 31) {real, imag} */,
  {32'hc0f329e4, 32'h3f82c0f8} /* (24, 14, 30) {real, imag} */,
  {32'hc048f116, 32'h400ac658} /* (24, 14, 29) {real, imag} */,
  {32'hc00fccba, 32'h40049248} /* (24, 14, 28) {real, imag} */,
  {32'hc0c58be4, 32'h40101ff7} /* (24, 14, 27) {real, imag} */,
  {32'hc0c95bd1, 32'h3fe1a22f} /* (24, 14, 26) {real, imag} */,
  {32'hc001eb53, 32'h3f965f2e} /* (24, 14, 25) {real, imag} */,
  {32'h40b6ff4c, 32'h40006b62} /* (24, 14, 24) {real, imag} */,
  {32'hbf3118f0, 32'hbfdf4878} /* (24, 14, 23) {real, imag} */,
  {32'hc0bcc7a8, 32'hbfc506a0} /* (24, 14, 22) {real, imag} */,
  {32'hc01d5f88, 32'h402299d2} /* (24, 14, 21) {real, imag} */,
  {32'hc08814ec, 32'h3ee93dd8} /* (24, 14, 20) {real, imag} */,
  {32'hc041646c, 32'hc05f74db} /* (24, 14, 19) {real, imag} */,
  {32'h3f945b0c, 32'hbe70a3f8} /* (24, 14, 18) {real, imag} */,
  {32'h3ea4cf50, 32'hbf8b80b8} /* (24, 14, 17) {real, imag} */,
  {32'h3fa39eae, 32'hbf617ee0} /* (24, 14, 16) {real, imag} */,
  {32'h3fc9fdfa, 32'h3e3331a0} /* (24, 14, 15) {real, imag} */,
  {32'h4099e55c, 32'h3f1a6f1a} /* (24, 14, 14) {real, imag} */,
  {32'h3fad1766, 32'hbfc363f8} /* (24, 14, 13) {real, imag} */,
  {32'hc013f333, 32'h3fbdfada} /* (24, 14, 12) {real, imag} */,
  {32'hc035e066, 32'h3e3c1ba0} /* (24, 14, 11) {real, imag} */,
  {32'hbf0b63d8, 32'hc089b574} /* (24, 14, 10) {real, imag} */,
  {32'hc0297b4e, 32'hc066decb} /* (24, 14, 9) {real, imag} */,
  {32'h3fe6dda4, 32'hbfa8f789} /* (24, 14, 8) {real, imag} */,
  {32'h3f6dbbf8, 32'h408a0fe0} /* (24, 14, 7) {real, imag} */,
  {32'hc08c087d, 32'h40d4b00e} /* (24, 14, 6) {real, imag} */,
  {32'hbfd29090, 32'h3fcc4804} /* (24, 14, 5) {real, imag} */,
  {32'h405392a4, 32'hbf88997c} /* (24, 14, 4) {real, imag} */,
  {32'h4076ea78, 32'h406fa86c} /* (24, 14, 3) {real, imag} */,
  {32'h3f3ae234, 32'h3ea74060} /* (24, 14, 2) {real, imag} */,
  {32'hbff01bd4, 32'hc02a9435} /* (24, 14, 1) {real, imag} */,
  {32'h3e910c44, 32'hbec517f0} /* (24, 14, 0) {real, imag} */,
  {32'hbea69c74, 32'hbf26c6e6} /* (24, 13, 31) {real, imag} */,
  {32'hc00277bf, 32'h407265cc} /* (24, 13, 30) {real, imag} */,
  {32'hc038223d, 32'h3f956854} /* (24, 13, 29) {real, imag} */,
  {32'hc056be07, 32'hc02deffe} /* (24, 13, 28) {real, imag} */,
  {32'hc04c0186, 32'hbefe3038} /* (24, 13, 27) {real, imag} */,
  {32'hc0cbc1f8, 32'hc015cfd3} /* (24, 13, 26) {real, imag} */,
  {32'hc0a748be, 32'h40263752} /* (24, 13, 25) {real, imag} */,
  {32'h3ef26354, 32'h3fc22fb2} /* (24, 13, 24) {real, imag} */,
  {32'hc033ca15, 32'hc0a04d96} /* (24, 13, 23) {real, imag} */,
  {32'hbef96fe8, 32'hc006504c} /* (24, 13, 22) {real, imag} */,
  {32'hbf7b0cc0, 32'h4049bc25} /* (24, 13, 21) {real, imag} */,
  {32'h3f68f2b0, 32'h4097db12} /* (24, 13, 20) {real, imag} */,
  {32'h400aba30, 32'h3f98f498} /* (24, 13, 19) {real, imag} */,
  {32'h400bcc6d, 32'hbf911e28} /* (24, 13, 18) {real, imag} */,
  {32'h40e818a8, 32'h3fef297f} /* (24, 13, 17) {real, imag} */,
  {32'h3f99f29c, 32'h3fbe1222} /* (24, 13, 16) {real, imag} */,
  {32'h3fe1d9ed, 32'hbe303180} /* (24, 13, 15) {real, imag} */,
  {32'h40ac1561, 32'hbfac7615} /* (24, 13, 14) {real, imag} */,
  {32'h406e5030, 32'hbff38752} /* (24, 13, 13) {real, imag} */,
  {32'h40aff528, 32'h40bb007f} /* (24, 13, 12) {real, imag} */,
  {32'hbe89aa70, 32'h409289a6} /* (24, 13, 11) {real, imag} */,
  {32'h3e6a56b0, 32'h400787e4} /* (24, 13, 10) {real, imag} */,
  {32'h405434b5, 32'h3f6d5c82} /* (24, 13, 9) {real, imag} */,
  {32'h408800d7, 32'hc0c345af} /* (24, 13, 8) {real, imag} */,
  {32'h408e7996, 32'hc0753176} /* (24, 13, 7) {real, imag} */,
  {32'h40746e7e, 32'hc00cceb4} /* (24, 13, 6) {real, imag} */,
  {32'h4015e7bc, 32'h3ec80d00} /* (24, 13, 5) {real, imag} */,
  {32'hbf9732d4, 32'h408ae4a2} /* (24, 13, 4) {real, imag} */,
  {32'h3d331620, 32'hbf040be8} /* (24, 13, 3) {real, imag} */,
  {32'h400346b6, 32'hc039d915} /* (24, 13, 2) {real, imag} */,
  {32'h409f0f8c, 32'h408d7cda} /* (24, 13, 1) {real, imag} */,
  {32'h40a5d7d0, 32'h3f3a5a78} /* (24, 13, 0) {real, imag} */,
  {32'hc0d8d290, 32'hbf2627b4} /* (24, 12, 31) {real, imag} */,
  {32'h3f8247c2, 32'h3c86a280} /* (24, 12, 30) {real, imag} */,
  {32'h40d6ca6b, 32'h3fb401ca} /* (24, 12, 29) {real, imag} */,
  {32'h40b767ad, 32'hbfa7072c} /* (24, 12, 28) {real, imag} */,
  {32'h408b4062, 32'h3df1aa40} /* (24, 12, 27) {real, imag} */,
  {32'hbead76b0, 32'hbf0b3a34} /* (24, 12, 26) {real, imag} */,
  {32'h40160abf, 32'h405bda40} /* (24, 12, 25) {real, imag} */,
  {32'hbff9b640, 32'h4053687f} /* (24, 12, 24) {real, imag} */,
  {32'hc0738116, 32'h40176912} /* (24, 12, 23) {real, imag} */,
  {32'hc08f69b6, 32'hc086b3ce} /* (24, 12, 22) {real, imag} */,
  {32'hbc965c00, 32'hbfe4d5c0} /* (24, 12, 21) {real, imag} */,
  {32'h3f833724, 32'hbf6429c8} /* (24, 12, 20) {real, imag} */,
  {32'h3b1c2600, 32'hc03891ba} /* (24, 12, 19) {real, imag} */,
  {32'hc0b76522, 32'h40361081} /* (24, 12, 18) {real, imag} */,
  {32'hc0aa38a1, 32'h40bd02bf} /* (24, 12, 17) {real, imag} */,
  {32'h3f454380, 32'h40b00f3e} /* (24, 12, 16) {real, imag} */,
  {32'h3f7668b4, 32'h40169bf4} /* (24, 12, 15) {real, imag} */,
  {32'hbd83f980, 32'h3fec12a0} /* (24, 12, 14) {real, imag} */,
  {32'hc00119a4, 32'hbf7342ec} /* (24, 12, 13) {real, imag} */,
  {32'hc0867673, 32'h3f7b81f2} /* (24, 12, 12) {real, imag} */,
  {32'hc034833e, 32'hc049d1b2} /* (24, 12, 11) {real, imag} */,
  {32'h40706bf2, 32'hc07f35c2} /* (24, 12, 10) {real, imag} */,
  {32'h400e9de1, 32'hc056ffe3} /* (24, 12, 9) {real, imag} */,
  {32'hc087cfb9, 32'h40c74a8e} /* (24, 12, 8) {real, imag} */,
  {32'hc0157e5e, 32'h412d0998} /* (24, 12, 7) {real, imag} */,
  {32'hc09b6f81, 32'h3f593eb8} /* (24, 12, 6) {real, imag} */,
  {32'hbd981a00, 32'h403db5e3} /* (24, 12, 5) {real, imag} */,
  {32'h4003d069, 32'h40a2ea6c} /* (24, 12, 4) {real, imag} */,
  {32'h3ea999f4, 32'h40a5b944} /* (24, 12, 3) {real, imag} */,
  {32'hc04d48c6, 32'h3fd68619} /* (24, 12, 2) {real, imag} */,
  {32'h3fa10388, 32'h40afbf28} /* (24, 12, 1) {real, imag} */,
  {32'hbfb702aa, 32'h4086806e} /* (24, 12, 0) {real, imag} */,
  {32'hbfc20f86, 32'h3fd317c0} /* (24, 11, 31) {real, imag} */,
  {32'hbff51c3d, 32'h3e0673b0} /* (24, 11, 30) {real, imag} */,
  {32'hbfaac232, 32'h4021b430} /* (24, 11, 29) {real, imag} */,
  {32'h3fa3f494, 32'h40b7f576} /* (24, 11, 28) {real, imag} */,
  {32'hc028558c, 32'hc0076f05} /* (24, 11, 27) {real, imag} */,
  {32'h4081d932, 32'hc062c778} /* (24, 11, 26) {real, imag} */,
  {32'h404d7804, 32'h40c0a638} /* (24, 11, 25) {real, imag} */,
  {32'hc0d4e73d, 32'h41117c30} /* (24, 11, 24) {real, imag} */,
  {32'hc0a868d9, 32'h40cf1de2} /* (24, 11, 23) {real, imag} */,
  {32'hc056a038, 32'h403f4b45} /* (24, 11, 22) {real, imag} */,
  {32'hc03450fc, 32'hbf9dcbb0} /* (24, 11, 21) {real, imag} */,
  {32'h4051db01, 32'h4006fcbe} /* (24, 11, 20) {real, imag} */,
  {32'h3fd00c18, 32'h3f5ccd10} /* (24, 11, 19) {real, imag} */,
  {32'h40a0065e, 32'hc07f5cd1} /* (24, 11, 18) {real, imag} */,
  {32'h4012f094, 32'hc10ab40f} /* (24, 11, 17) {real, imag} */,
  {32'hc09cd13f, 32'hc0b5723f} /* (24, 11, 16) {real, imag} */,
  {32'hc0263ab0, 32'hc06ac182} /* (24, 11, 15) {real, imag} */,
  {32'hbf3db66c, 32'hbf8f5b35} /* (24, 11, 14) {real, imag} */,
  {32'hc0547c7c, 32'h4091dbb8} /* (24, 11, 13) {real, imag} */,
  {32'h404ae5d8, 32'hbf827310} /* (24, 11, 12) {real, imag} */,
  {32'h40c2acc9, 32'hc0d19409} /* (24, 11, 11) {real, imag} */,
  {32'h403e5b65, 32'hc031256b} /* (24, 11, 10) {real, imag} */,
  {32'h40081853, 32'hc0a373ee} /* (24, 11, 9) {real, imag} */,
  {32'hc02cb5a5, 32'hc0ae8f9d} /* (24, 11, 8) {real, imag} */,
  {32'hc10981c8, 32'hbf7962a8} /* (24, 11, 7) {real, imag} */,
  {32'hc0a75ffa, 32'h3fdf509e} /* (24, 11, 6) {real, imag} */,
  {32'hc027eb8f, 32'h40cb8ce4} /* (24, 11, 5) {real, imag} */,
  {32'h40284441, 32'h4073aaf2} /* (24, 11, 4) {real, imag} */,
  {32'h40c660cc, 32'h3f5be068} /* (24, 11, 3) {real, imag} */,
  {32'h4083e83e, 32'h3ea827c8} /* (24, 11, 2) {real, imag} */,
  {32'hbf2fccf0, 32'hbe7e12a0} /* (24, 11, 1) {real, imag} */,
  {32'hbf702c84, 32'hbeeaa8b8} /* (24, 11, 0) {real, imag} */,
  {32'hc0721e16, 32'hc089d258} /* (24, 10, 31) {real, imag} */,
  {32'hc01a79d6, 32'hc080479e} /* (24, 10, 30) {real, imag} */,
  {32'hc0098386, 32'hc0ac9929} /* (24, 10, 29) {real, imag} */,
  {32'hc09b84e2, 32'h3f5554a4} /* (24, 10, 28) {real, imag} */,
  {32'h3f87b216, 32'hbf908316} /* (24, 10, 27) {real, imag} */,
  {32'hbe8e0ae8, 32'h3fdb133f} /* (24, 10, 26) {real, imag} */,
  {32'hc00317f4, 32'hc0b3465a} /* (24, 10, 25) {real, imag} */,
  {32'h3fc5632e, 32'hc030c8c1} /* (24, 10, 24) {real, imag} */,
  {32'h3f450a60, 32'h40c2cff8} /* (24, 10, 23) {real, imag} */,
  {32'h3fb832d7, 32'h403fed9a} /* (24, 10, 22) {real, imag} */,
  {32'h40bdf05b, 32'h3eac2610} /* (24, 10, 21) {real, imag} */,
  {32'h3f1483e4, 32'h40d42594} /* (24, 10, 20) {real, imag} */,
  {32'hc0dea034, 32'h3fe96dcc} /* (24, 10, 19) {real, imag} */,
  {32'hc1282dac, 32'hbfc8e452} /* (24, 10, 18) {real, imag} */,
  {32'h3f51d22c, 32'h3e94acf0} /* (24, 10, 17) {real, imag} */,
  {32'hbf683a16, 32'hbed01518} /* (24, 10, 16) {real, imag} */,
  {32'h3f0a1ecc, 32'hbed83b60} /* (24, 10, 15) {real, imag} */,
  {32'h40275472, 32'hbffe05fe} /* (24, 10, 14) {real, imag} */,
  {32'hc0a90f66, 32'hc040c7be} /* (24, 10, 13) {real, imag} */,
  {32'hc188c949, 32'hc0ad501f} /* (24, 10, 12) {real, imag} */,
  {32'hc15c13a8, 32'hc0712e40} /* (24, 10, 11) {real, imag} */,
  {32'hc132dac2, 32'hc0f45d8d} /* (24, 10, 10) {real, imag} */,
  {32'hc07ea183, 32'hc166d570} /* (24, 10, 9) {real, imag} */,
  {32'h4128a1c0, 32'hc166bb4c} /* (24, 10, 8) {real, imag} */,
  {32'h40dacfc5, 32'hc123c844} /* (24, 10, 7) {real, imag} */,
  {32'hc069e5fd, 32'hc0e13be0} /* (24, 10, 6) {real, imag} */,
  {32'hc129b7b2, 32'hc0cd953c} /* (24, 10, 5) {real, imag} */,
  {32'hc07a7977, 32'h40331a9a} /* (24, 10, 4) {real, imag} */,
  {32'h410d7736, 32'h3f8d8bca} /* (24, 10, 3) {real, imag} */,
  {32'h40bdf0e5, 32'h407b0164} /* (24, 10, 2) {real, imag} */,
  {32'h40ce074c, 32'h3f05ad58} /* (24, 10, 1) {real, imag} */,
  {32'h401feef9, 32'h3f41e84c} /* (24, 10, 0) {real, imag} */,
  {32'h408d3ac8, 32'hc0862d66} /* (24, 9, 31) {real, imag} */,
  {32'h40b66f2f, 32'hc0d54f3a} /* (24, 9, 30) {real, imag} */,
  {32'h40212b3b, 32'hbf805f60} /* (24, 9, 29) {real, imag} */,
  {32'h40a44c09, 32'h4123ebaf} /* (24, 9, 28) {real, imag} */,
  {32'h40bc79de, 32'h40a5a106} /* (24, 9, 27) {real, imag} */,
  {32'h40f42414, 32'h40900a55} /* (24, 9, 26) {real, imag} */,
  {32'hc00e6a96, 32'h40ce788e} /* (24, 9, 25) {real, imag} */,
  {32'h3e7d92f0, 32'hc09fb033} /* (24, 9, 24) {real, imag} */,
  {32'h40a22d72, 32'hc1144151} /* (24, 9, 23) {real, imag} */,
  {32'hbfeb43c2, 32'hc110dcc8} /* (24, 9, 22) {real, imag} */,
  {32'h40639755, 32'hc06fb3df} /* (24, 9, 21) {real, imag} */,
  {32'hc1608a9d, 32'hc108ce26} /* (24, 9, 20) {real, imag} */,
  {32'hc0ca7ef9, 32'hc0ccbba0} /* (24, 9, 19) {real, imag} */,
  {32'hc053b472, 32'hc0c5893d} /* (24, 9, 18) {real, imag} */,
  {32'h3f553338, 32'hc127174d} /* (24, 9, 17) {real, imag} */,
  {32'h4080ea3c, 32'hc04c6236} /* (24, 9, 16) {real, imag} */,
  {32'h3e2727b0, 32'hc0fd66d8} /* (24, 9, 15) {real, imag} */,
  {32'h4116c29f, 32'hbfbe1fdc} /* (24, 9, 14) {real, imag} */,
  {32'h40c27fca, 32'hc103fd37} /* (24, 9, 13) {real, imag} */,
  {32'h3f6364bc, 32'hbc3ebb00} /* (24, 9, 12) {real, imag} */,
  {32'hbf9ac2d4, 32'hc0a1c5e4} /* (24, 9, 11) {real, imag} */,
  {32'hbe633d40, 32'hc10b3eb9} /* (24, 9, 10) {real, imag} */,
  {32'h40953f66, 32'hc118fd90} /* (24, 9, 9) {real, imag} */,
  {32'h40287823, 32'hc0d9034d} /* (24, 9, 8) {real, imag} */,
  {32'hc0ce0d93, 32'h409278df} /* (24, 9, 7) {real, imag} */,
  {32'hc0a2cc6b, 32'hc0d694b0} /* (24, 9, 6) {real, imag} */,
  {32'hc0d4dec4, 32'h4030926c} /* (24, 9, 5) {real, imag} */,
  {32'hc11932a9, 32'h400734b6} /* (24, 9, 4) {real, imag} */,
  {32'hc09077eb, 32'hc0aa11ce} /* (24, 9, 3) {real, imag} */,
  {32'hc0fb75d6, 32'h3eaf1158} /* (24, 9, 2) {real, imag} */,
  {32'hc003a69c, 32'h40a090bd} /* (24, 9, 1) {real, imag} */,
  {32'hc0665314, 32'hc094977f} /* (24, 9, 0) {real, imag} */,
  {32'h401b19db, 32'hbfc9c868} /* (24, 8, 31) {real, imag} */,
  {32'h40be068e, 32'h4126d25d} /* (24, 8, 30) {real, imag} */,
  {32'h40f21d38, 32'h418da37c} /* (24, 8, 29) {real, imag} */,
  {32'hbfea34cc, 32'h4138256c} /* (24, 8, 28) {real, imag} */,
  {32'h409deacb, 32'h4006afcc} /* (24, 8, 27) {real, imag} */,
  {32'h40ea19b5, 32'hc0940453} /* (24, 8, 26) {real, imag} */,
  {32'h40d1d212, 32'hbf545610} /* (24, 8, 25) {real, imag} */,
  {32'h40f3d806, 32'hc098b59c} /* (24, 8, 24) {real, imag} */,
  {32'h40b0e449, 32'h3e399c28} /* (24, 8, 23) {real, imag} */,
  {32'h40a02b97, 32'h400df52c} /* (24, 8, 22) {real, imag} */,
  {32'h40bd4c39, 32'h416aa9ef} /* (24, 8, 21) {real, imag} */,
  {32'hc090ade0, 32'h40b86431} /* (24, 8, 20) {real, imag} */,
  {32'hc168d09a, 32'hc1116610} /* (24, 8, 19) {real, imag} */,
  {32'hc16d91e5, 32'hc115f170} /* (24, 8, 18) {real, imag} */,
  {32'hbf20e78c, 32'hc13f54e8} /* (24, 8, 17) {real, imag} */,
  {32'h40cd117e, 32'hc1caf366} /* (24, 8, 16) {real, imag} */,
  {32'h401a3b8f, 32'hc1cf4048} /* (24, 8, 15) {real, imag} */,
  {32'h403a7d02, 32'hc197c5b2} /* (24, 8, 14) {real, imag} */,
  {32'hbed34aa8, 32'hc1199654} /* (24, 8, 13) {real, imag} */,
  {32'h3dbdc700, 32'hc13abdbe} /* (24, 8, 12) {real, imag} */,
  {32'h40a139c3, 32'hc04b046e} /* (24, 8, 11) {real, imag} */,
  {32'h406f47a2, 32'h41310620} /* (24, 8, 10) {real, imag} */,
  {32'hbf334908, 32'h418a4712} /* (24, 8, 9) {real, imag} */,
  {32'h4077c545, 32'h4159be46} /* (24, 8, 8) {real, imag} */,
  {32'h41774293, 32'h40e04559} /* (24, 8, 7) {real, imag} */,
  {32'h41292ea4, 32'h4099d036} /* (24, 8, 6) {real, imag} */,
  {32'hbf136ad0, 32'h412c6eed} /* (24, 8, 5) {real, imag} */,
  {32'hc0c599da, 32'h41658163} /* (24, 8, 4) {real, imag} */,
  {32'hbfe50b2c, 32'h4144f873} /* (24, 8, 3) {real, imag} */,
  {32'h4113592d, 32'h408f9f32} /* (24, 8, 2) {real, imag} */,
  {32'hc03ce17c, 32'h402f71a1} /* (24, 8, 1) {real, imag} */,
  {32'hbfb5018c, 32'h4055f444} /* (24, 8, 0) {real, imag} */,
  {32'h4018b90d, 32'h40af3a8e} /* (24, 7, 31) {real, imag} */,
  {32'h4006faba, 32'h40aeee06} /* (24, 7, 30) {real, imag} */,
  {32'hc0087a9f, 32'hc057a9c8} /* (24, 7, 29) {real, imag} */,
  {32'hbe9c854c, 32'h3f767630} /* (24, 7, 28) {real, imag} */,
  {32'hc166628d, 32'h40e9ed7e} /* (24, 7, 27) {real, imag} */,
  {32'hc1866316, 32'hc1130cb8} /* (24, 7, 26) {real, imag} */,
  {32'hbf1ad418, 32'hc18cec39} /* (24, 7, 25) {real, imag} */,
  {32'h409511d3, 32'hc09f310a} /* (24, 7, 24) {real, imag} */,
  {32'h403c1d84, 32'hc190e464} /* (24, 7, 23) {real, imag} */,
  {32'hc0a17ea6, 32'hc1cfec8c} /* (24, 7, 22) {real, imag} */,
  {32'hc1046d60, 32'hc1048b5b} /* (24, 7, 21) {real, imag} */,
  {32'h4059e5a3, 32'hbfc38132} /* (24, 7, 20) {real, imag} */,
  {32'h4123ade2, 32'h410ec301} /* (24, 7, 19) {real, imag} */,
  {32'h41001618, 32'hbfde46ec} /* (24, 7, 18) {real, imag} */,
  {32'hbf8afce8, 32'hc06aadc6} /* (24, 7, 17) {real, imag} */,
  {32'hc08363d4, 32'hc0ba7803} /* (24, 7, 16) {real, imag} */,
  {32'hc09e4114, 32'hc0b9c0b8} /* (24, 7, 15) {real, imag} */,
  {32'hbf560130, 32'h4064373c} /* (24, 7, 14) {real, imag} */,
  {32'hc043f9e9, 32'hbfb2c568} /* (24, 7, 13) {real, imag} */,
  {32'hc0661ff7, 32'hc132fff2} /* (24, 7, 12) {real, imag} */,
  {32'hc0f575e6, 32'hc05c9a9c} /* (24, 7, 11) {real, imag} */,
  {32'hc0a57d7f, 32'hbf994390} /* (24, 7, 10) {real, imag} */,
  {32'hc05ad7bf, 32'h4096197a} /* (24, 7, 9) {real, imag} */,
  {32'hc111680c, 32'h4106318c} /* (24, 7, 8) {real, imag} */,
  {32'hbefbd050, 32'hbfa6c72b} /* (24, 7, 7) {real, imag} */,
  {32'h40f81593, 32'hc1730bf0} /* (24, 7, 6) {real, imag} */,
  {32'h413b05cb, 32'hc111c42d} /* (24, 7, 5) {real, imag} */,
  {32'h411b2cff, 32'h3e83354c} /* (24, 7, 4) {real, imag} */,
  {32'h4016a01a, 32'h406c04b0} /* (24, 7, 3) {real, imag} */,
  {32'hc15b97d9, 32'hc0de0350} /* (24, 7, 2) {real, imag} */,
  {32'hc0e35a4f, 32'hc100bba6} /* (24, 7, 1) {real, imag} */,
  {32'h3dc6ce00, 32'hc0d5dd8a} /* (24, 7, 0) {real, imag} */,
  {32'h3f9dd1cc, 32'h3e8ea170} /* (24, 6, 31) {real, imag} */,
  {32'hc13ec72d, 32'hc0de1cc4} /* (24, 6, 30) {real, imag} */,
  {32'hc1c35792, 32'hc01adf42} /* (24, 6, 29) {real, imag} */,
  {32'hc150933b, 32'hc05b51ff} /* (24, 6, 28) {real, imag} */,
  {32'hc0e3d7dd, 32'hc159e4a5} /* (24, 6, 27) {real, imag} */,
  {32'hc1051e84, 32'hc1644e9d} /* (24, 6, 26) {real, imag} */,
  {32'hbf22dc90, 32'hc11e4ae3} /* (24, 6, 25) {real, imag} */,
  {32'hc03e7f20, 32'hc04c38b6} /* (24, 6, 24) {real, imag} */,
  {32'hc0c07e6e, 32'h40d6b4ec} /* (24, 6, 23) {real, imag} */,
  {32'h408516d7, 32'h407a326e} /* (24, 6, 22) {real, imag} */,
  {32'hbf1f2de4, 32'hc19394e3} /* (24, 6, 21) {real, imag} */,
  {32'h402fc4ff, 32'hc18c30d0} /* (24, 6, 20) {real, imag} */,
  {32'h409bb3d0, 32'h3ffa6fcc} /* (24, 6, 19) {real, imag} */,
  {32'h4108ec8e, 32'h4120bb77} /* (24, 6, 18) {real, imag} */,
  {32'hbf1b22b8, 32'h41a00d60} /* (24, 6, 17) {real, imag} */,
  {32'hc0f133d4, 32'h410d99c4} /* (24, 6, 16) {real, imag} */,
  {32'h40342fd3, 32'h40f0f2d8} /* (24, 6, 15) {real, imag} */,
  {32'hc0ba9847, 32'h414ea486} /* (24, 6, 14) {real, imag} */,
  {32'h3fd6c744, 32'h3fd20448} /* (24, 6, 13) {real, imag} */,
  {32'hc0ad5b30, 32'h3fc1aede} /* (24, 6, 12) {real, imag} */,
  {32'hc0c2cb5a, 32'hc084de40} /* (24, 6, 11) {real, imag} */,
  {32'hbeb35600, 32'h3f9d6f0d} /* (24, 6, 10) {real, imag} */,
  {32'h3f215c8c, 32'h4060cc7b} /* (24, 6, 9) {real, imag} */,
  {32'h412917da, 32'h3f74cab0} /* (24, 6, 8) {real, imag} */,
  {32'h40c24a2b, 32'hc09df158} /* (24, 6, 7) {real, imag} */,
  {32'hc0aa7383, 32'hbeb83ae8} /* (24, 6, 6) {real, imag} */,
  {32'hc1109e02, 32'h412a0d52} /* (24, 6, 5) {real, imag} */,
  {32'hc1bb6bbc, 32'hc04abc9e} /* (24, 6, 4) {real, imag} */,
  {32'hc03c47ed, 32'hc0847cf5} /* (24, 6, 3) {real, imag} */,
  {32'h419b0e5f, 32'hbfabb4a8} /* (24, 6, 2) {real, imag} */,
  {32'h40c62d00, 32'h404b6c6c} /* (24, 6, 1) {real, imag} */,
  {32'h4018f575, 32'h408465b0} /* (24, 6, 0) {real, imag} */,
  {32'hbee54740, 32'hc0d7975b} /* (24, 5, 31) {real, imag} */,
  {32'hc0ab9529, 32'hbfb49d40} /* (24, 5, 30) {real, imag} */,
  {32'hc06f73ed, 32'h3fbdbd80} /* (24, 5, 29) {real, imag} */,
  {32'hbffe8558, 32'h40d51806} /* (24, 5, 28) {real, imag} */,
  {32'hc07e9f84, 32'h41857848} /* (24, 5, 27) {real, imag} */,
  {32'h40148528, 32'h4182d8ca} /* (24, 5, 26) {real, imag} */,
  {32'hc013b4fc, 32'h40896640} /* (24, 5, 25) {real, imag} */,
  {32'h411bcefd, 32'h3d6eb0c0} /* (24, 5, 24) {real, imag} */,
  {32'hbff64490, 32'h3f0da310} /* (24, 5, 23) {real, imag} */,
  {32'hc04ad884, 32'h41a560d0} /* (24, 5, 22) {real, imag} */,
  {32'h3f8b9fbc, 32'h417aaba3} /* (24, 5, 21) {real, imag} */,
  {32'hc0c04870, 32'h4082233d} /* (24, 5, 20) {real, imag} */,
  {32'hc0d6cbf8, 32'hbff0cc72} /* (24, 5, 19) {real, imag} */,
  {32'h406ad147, 32'h4082e5be} /* (24, 5, 18) {real, imag} */,
  {32'h4020d476, 32'hc0635c0a} /* (24, 5, 17) {real, imag} */,
  {32'h40c9f89c, 32'hc13c11e6} /* (24, 5, 16) {real, imag} */,
  {32'hbee3c1a0, 32'hc1c12eb8} /* (24, 5, 15) {real, imag} */,
  {32'hc00ea55e, 32'h4001fa42} /* (24, 5, 14) {real, imag} */,
  {32'hc0605b66, 32'hc0a59cfe} /* (24, 5, 13) {real, imag} */,
  {32'hbf8b6b54, 32'h3fe5ee64} /* (24, 5, 12) {real, imag} */,
  {32'h40077406, 32'hc0ec2a42} /* (24, 5, 11) {real, imag} */,
  {32'h40853e74, 32'hc0af2d8f} /* (24, 5, 10) {real, imag} */,
  {32'h411e8afc, 32'h410f7412} /* (24, 5, 9) {real, imag} */,
  {32'h41202765, 32'h4090c961} /* (24, 5, 8) {real, imag} */,
  {32'h3fd238b0, 32'h3fceb2dc} /* (24, 5, 7) {real, imag} */,
  {32'h3ff69518, 32'h41029c98} /* (24, 5, 6) {real, imag} */,
  {32'hc10acb16, 32'h40727a7a} /* (24, 5, 5) {real, imag} */,
  {32'hbdd3ba20, 32'h40dba13e} /* (24, 5, 4) {real, imag} */,
  {32'h408eca5e, 32'h407721cc} /* (24, 5, 3) {real, imag} */,
  {32'h401111fa, 32'h40908bb4} /* (24, 5, 2) {real, imag} */,
  {32'h411d354f, 32'h3fe3275c} /* (24, 5, 1) {real, imag} */,
  {32'h407b8f24, 32'h40152027} /* (24, 5, 0) {real, imag} */,
  {32'h407e25d0, 32'hc128157f} /* (24, 4, 31) {real, imag} */,
  {32'hc11f08f4, 32'h3e81cca8} /* (24, 4, 30) {real, imag} */,
  {32'hc153a248, 32'h4091393c} /* (24, 4, 29) {real, imag} */,
  {32'h3fbdba1a, 32'h41575a60} /* (24, 4, 28) {real, imag} */,
  {32'hc0e3f0b6, 32'h40cff712} /* (24, 4, 27) {real, imag} */,
  {32'hc13bf270, 32'h3f526244} /* (24, 4, 26) {real, imag} */,
  {32'h40874fb4, 32'hc11cfc70} /* (24, 4, 25) {real, imag} */,
  {32'h40d1cd0a, 32'hc1855401} /* (24, 4, 24) {real, imag} */,
  {32'hbf2e1060, 32'hc17c698c} /* (24, 4, 23) {real, imag} */,
  {32'hc0fd3390, 32'hc1c61ea7} /* (24, 4, 22) {real, imag} */,
  {32'hc1c12244, 32'hbf4fbc98} /* (24, 4, 21) {real, imag} */,
  {32'h3f448bc0, 32'h40abc039} /* (24, 4, 20) {real, imag} */,
  {32'h4127d419, 32'h402d1260} /* (24, 4, 19) {real, imag} */,
  {32'hbf994fb0, 32'h4189a476} /* (24, 4, 18) {real, imag} */,
  {32'h40c2f408, 32'h4209947c} /* (24, 4, 17) {real, imag} */,
  {32'h40c69422, 32'h41fddbc4} /* (24, 4, 16) {real, imag} */,
  {32'hc0a7dfca, 32'h419d0759} /* (24, 4, 15) {real, imag} */,
  {32'hc10bddf8, 32'h417b70fa} /* (24, 4, 14) {real, imag} */,
  {32'h3f1ced50, 32'h3f428b40} /* (24, 4, 13) {real, imag} */,
  {32'h40ce56f3, 32'hc0910d60} /* (24, 4, 12) {real, imag} */,
  {32'h414961b2, 32'h40e47d88} /* (24, 4, 11) {real, imag} */,
  {32'h41687fea, 32'hc0a22a65} /* (24, 4, 10) {real, imag} */,
  {32'h409f0782, 32'hc113d10e} /* (24, 4, 9) {real, imag} */,
  {32'hc0556234, 32'hc195fd22} /* (24, 4, 8) {real, imag} */,
  {32'hc05917b4, 32'hc145d3d2} /* (24, 4, 7) {real, imag} */,
  {32'h410fe0b7, 32'hc14e3616} /* (24, 4, 6) {real, imag} */,
  {32'h414165d0, 32'hc1600a88} /* (24, 4, 5) {real, imag} */,
  {32'hc015117d, 32'hc0d87786} /* (24, 4, 4) {real, imag} */,
  {32'hc0ab61a7, 32'h4131903a} /* (24, 4, 3) {real, imag} */,
  {32'hbe8055f0, 32'h4083ceab} /* (24, 4, 2) {real, imag} */,
  {32'hbe953c18, 32'hc1ac3502} /* (24, 4, 1) {real, imag} */,
  {32'h3ef38bb8, 32'hc1944d0b} /* (24, 4, 0) {real, imag} */,
  {32'h41374f42, 32'hbe9ac040} /* (24, 3, 31) {real, imag} */,
  {32'h4099d2b0, 32'hbe4c5240} /* (24, 3, 30) {real, imag} */,
  {32'h41022ee6, 32'hc01b4de0} /* (24, 3, 29) {real, imag} */,
  {32'hbfad3b5e, 32'hc06c5d2a} /* (24, 3, 28) {real, imag} */,
  {32'hc143d146, 32'hc179040f} /* (24, 3, 27) {real, imag} */,
  {32'h41339803, 32'hc0aa2c0c} /* (24, 3, 26) {real, imag} */,
  {32'h4173a452, 32'h40b9a710} /* (24, 3, 25) {real, imag} */,
  {32'h4021db54, 32'h41b0c090} /* (24, 3, 24) {real, imag} */,
  {32'h40319a08, 32'hbf0b7470} /* (24, 3, 23) {real, imag} */,
  {32'h40fcd790, 32'h414a9546} /* (24, 3, 22) {real, imag} */,
  {32'h410e19a4, 32'h41ba9e12} /* (24, 3, 21) {real, imag} */,
  {32'hc0b6d3ae, 32'h40a688bc} /* (24, 3, 20) {real, imag} */,
  {32'hc12aca53, 32'h4108a7c0} /* (24, 3, 19) {real, imag} */,
  {32'hc1e58c75, 32'hc0fbf034} /* (24, 3, 18) {real, imag} */,
  {32'hc17e4973, 32'hc13a53fe} /* (24, 3, 17) {real, imag} */,
  {32'h3fa4a0b8, 32'hc136ccd9} /* (24, 3, 16) {real, imag} */,
  {32'h40fe830c, 32'hc02a2820} /* (24, 3, 15) {real, imag} */,
  {32'h4112c36a, 32'hc04ebe32} /* (24, 3, 14) {real, imag} */,
  {32'h41262faa, 32'h414571f1} /* (24, 3, 13) {real, imag} */,
  {32'h3f8656a3, 32'h40eb7450} /* (24, 3, 12) {real, imag} */,
  {32'hc009881e, 32'h4072a17b} /* (24, 3, 11) {real, imag} */,
  {32'h3cbc7b80, 32'h410f9cb0} /* (24, 3, 10) {real, imag} */,
  {32'h3f66c9f0, 32'hc04e3a1e} /* (24, 3, 9) {real, imag} */,
  {32'h40df8048, 32'hc11e0046} /* (24, 3, 8) {real, imag} */,
  {32'h41797b86, 32'hc1f29fb8} /* (24, 3, 7) {real, imag} */,
  {32'h4159517c, 32'hc1e93f0d} /* (24, 3, 6) {real, imag} */,
  {32'h40740ec8, 32'hc1034088} /* (24, 3, 5) {real, imag} */,
  {32'h4083e1a6, 32'h405e41b9} /* (24, 3, 4) {real, imag} */,
  {32'hc134521d, 32'h40a444a5} /* (24, 3, 3) {real, imag} */,
  {32'hc0a1c9cc, 32'hbfbeae46} /* (24, 3, 2) {real, imag} */,
  {32'h41024992, 32'hc0915804} /* (24, 3, 1) {real, imag} */,
  {32'h40798ccc, 32'h40242904} /* (24, 3, 0) {real, imag} */,
  {32'hc0a38964, 32'h3f684348} /* (24, 2, 31) {real, imag} */,
  {32'hc0e60ea4, 32'h41312d6b} /* (24, 2, 30) {real, imag} */,
  {32'h401ecf40, 32'h41a1578e} /* (24, 2, 29) {real, imag} */,
  {32'hc1536672, 32'h41bdaef1} /* (24, 2, 28) {real, imag} */,
  {32'hc0a693a6, 32'h41cf44da} /* (24, 2, 27) {real, imag} */,
  {32'h3f11cfd0, 32'h4203482f} /* (24, 2, 26) {real, imag} */,
  {32'hc0bac26e, 32'h41d96ff2} /* (24, 2, 25) {real, imag} */,
  {32'h40f26906, 32'h4100355f} /* (24, 2, 24) {real, imag} */,
  {32'h419787bc, 32'h3fbf1128} /* (24, 2, 23) {real, imag} */,
  {32'h41c27357, 32'h41e31c6e} /* (24, 2, 22) {real, imag} */,
  {32'h412a9db1, 32'h41b29c0f} /* (24, 2, 21) {real, imag} */,
  {32'hc18d875c, 32'hc11b4a68} /* (24, 2, 20) {real, imag} */,
  {32'hc21a42df, 32'hc1f0c1a5} /* (24, 2, 19) {real, imag} */,
  {32'hc1e02b38, 32'hc1cf69ac} /* (24, 2, 18) {real, imag} */,
  {32'hc210a5d1, 32'hc18d9966} /* (24, 2, 17) {real, imag} */,
  {32'hc20265d6, 32'hc18db5d7} /* (24, 2, 16) {real, imag} */,
  {32'hc1b0a159, 32'hc151e0f2} /* (24, 2, 15) {real, imag} */,
  {32'hc1b9cfda, 32'hc0fb9291} /* (24, 2, 14) {real, imag} */,
  {32'hc1934ceb, 32'hc198f286} /* (24, 2, 13) {real, imag} */,
  {32'hc1538529, 32'hc1262d6f} /* (24, 2, 12) {real, imag} */,
  {32'hbfbed124, 32'h409f12e9} /* (24, 2, 11) {real, imag} */,
  {32'h41de84c3, 32'h41b01c37} /* (24, 2, 10) {real, imag} */,
  {32'h41fa47ea, 32'h421a7762} /* (24, 2, 9) {real, imag} */,
  {32'h42024e63, 32'h41ddf2e2} /* (24, 2, 8) {real, imag} */,
  {32'h4230021b, 32'h4155e664} /* (24, 2, 7) {real, imag} */,
  {32'h4234e0f8, 32'h41a9e560} /* (24, 2, 6) {real, imag} */,
  {32'h4214a0c5, 32'h417cb7b0} /* (24, 2, 5) {real, imag} */,
  {32'h41539b4b, 32'h41a20939} /* (24, 2, 4) {real, imag} */,
  {32'h418e947f, 32'h41a0870e} /* (24, 2, 3) {real, imag} */,
  {32'h422c7dfe, 32'h41cd44a6} /* (24, 2, 2) {real, imag} */,
  {32'h41d1526d, 32'h41940a50} /* (24, 2, 1) {real, imag} */,
  {32'h41339175, 32'hbec99180} /* (24, 2, 0) {real, imag} */,
  {32'hc0b73c8a, 32'hc14660a7} /* (24, 1, 31) {real, imag} */,
  {32'hc1236d0d, 32'hc20b36b4} /* (24, 1, 30) {real, imag} */,
  {32'hc19bfbf1, 32'hc2243d14} /* (24, 1, 29) {real, imag} */,
  {32'hc1bf8be7, 32'hc20dca63} /* (24, 1, 28) {real, imag} */,
  {32'hc1c89e92, 32'hc1eb3c58} /* (24, 1, 27) {real, imag} */,
  {32'hc19423ad, 32'hc1d6f862} /* (24, 1, 26) {real, imag} */,
  {32'hc1d7a014, 32'hc2297f28} /* (24, 1, 25) {real, imag} */,
  {32'hc20527f5, 32'hc1faf346} /* (24, 1, 24) {real, imag} */,
  {32'hc0b77598, 32'hc2375fee} /* (24, 1, 23) {real, imag} */,
  {32'hc18d457d, 32'hc2194913} /* (24, 1, 22) {real, imag} */,
  {32'hc21bfd24, 32'hc170a14e} /* (24, 1, 21) {real, imag} */,
  {32'hc18fbb23, 32'h410bb559} /* (24, 1, 20) {real, imag} */,
  {32'hc0ece4a8, 32'h41341da6} /* (24, 1, 19) {real, imag} */,
  {32'hc1352539, 32'h42075694} /* (24, 1, 18) {real, imag} */,
  {32'hc0970aac, 32'h421f833d} /* (24, 1, 17) {real, imag} */,
  {32'h40d35de0, 32'h41a02f98} /* (24, 1, 16) {real, imag} */,
  {32'h41ea5ad2, 32'h4205047d} /* (24, 1, 15) {real, imag} */,
  {32'h41e68607, 32'h4207c8e4} /* (24, 1, 14) {real, imag} */,
  {32'h420c9172, 32'h4226aac9} /* (24, 1, 13) {real, imag} */,
  {32'h4151d07e, 32'h41d22605} /* (24, 1, 12) {real, imag} */,
  {32'h418c6828, 32'h418687e8} /* (24, 1, 11) {real, imag} */,
  {32'h4057ffdc, 32'hc186c7ee} /* (24, 1, 10) {real, imag} */,
  {32'h3fbd17a8, 32'hc209ad76} /* (24, 1, 9) {real, imag} */,
  {32'h41121e02, 32'hc1f65d50} /* (24, 1, 8) {real, imag} */,
  {32'h40f3628e, 32'hc194dabc} /* (24, 1, 7) {real, imag} */,
  {32'hc0b79f6b, 32'hc228042f} /* (24, 1, 6) {real, imag} */,
  {32'hc1a0ee13, 32'hc24cb546} /* (24, 1, 5) {real, imag} */,
  {32'hc1bdcee0, 32'hc22feab9} /* (24, 1, 4) {real, imag} */,
  {32'hc1d528a0, 32'hc21bda66} /* (24, 1, 3) {real, imag} */,
  {32'hc1850802, 32'hc234c4ec} /* (24, 1, 2) {real, imag} */,
  {32'hc19ba1d6, 32'hc1f3018d} /* (24, 1, 1) {real, imag} */,
  {32'hc13b97a2, 32'hc16fb0c4} /* (24, 1, 0) {real, imag} */,
  {32'hc1118b00, 32'hc107657b} /* (24, 0, 31) {real, imag} */,
  {32'hc17b727b, 32'hc189bc94} /* (24, 0, 30) {real, imag} */,
  {32'hc1b32ad5, 32'hc14d018f} /* (24, 0, 29) {real, imag} */,
  {32'hc203628e, 32'hc1f7cd86} /* (24, 0, 28) {real, imag} */,
  {32'hc192049e, 32'hc1d104bf} /* (24, 0, 27) {real, imag} */,
  {32'hc1789628, 32'hc1585b1c} /* (24, 0, 26) {real, imag} */,
  {32'hc0962602, 32'hc096ec7b} /* (24, 0, 25) {real, imag} */,
  {32'hc19177f9, 32'hbf5f72cc} /* (24, 0, 24) {real, imag} */,
  {32'hc1940360, 32'hc0ac12d0} /* (24, 0, 23) {real, imag} */,
  {32'hc1855953, 32'hc18bdce0} /* (24, 0, 22) {real, imag} */,
  {32'h40355732, 32'hc1c3a660} /* (24, 0, 21) {real, imag} */,
  {32'h408d3f0e, 32'h41cf5e0b} /* (24, 0, 20) {real, imag} */,
  {32'hc1261695, 32'h412b6513} /* (24, 0, 19) {real, imag} */,
  {32'h3f565e64, 32'hc18138ee} /* (24, 0, 18) {real, imag} */,
  {32'hbfad1102, 32'hc1208cc8} /* (24, 0, 17) {real, imag} */,
  {32'h40745659, 32'h40ea816b} /* (24, 0, 16) {real, imag} */,
  {32'h417fc145, 32'h41a73eb4} /* (24, 0, 15) {real, imag} */,
  {32'h420be86f, 32'h413b3b00} /* (24, 0, 14) {real, imag} */,
  {32'h41e65396, 32'h415db0b8} /* (24, 0, 13) {real, imag} */,
  {32'h41d01d13, 32'h4189f413} /* (24, 0, 12) {real, imag} */,
  {32'h41e079ac, 32'h41c251f4} /* (24, 0, 11) {real, imag} */,
  {32'h417373d7, 32'h4137e11c} /* (24, 0, 10) {real, imag} */,
  {32'hc00dad29, 32'hc15d8e6a} /* (24, 0, 9) {real, imag} */,
  {32'hc132a338, 32'hc10d2dc3} /* (24, 0, 8) {real, imag} */,
  {32'hc115051c, 32'hbe08e690} /* (24, 0, 7) {real, imag} */,
  {32'hc15d7dd2, 32'hbe2c3a70} /* (24, 0, 6) {real, imag} */,
  {32'hc0baa78c, 32'hc14e7980} /* (24, 0, 5) {real, imag} */,
  {32'hbfd17c80, 32'hc1c1bd62} /* (24, 0, 4) {real, imag} */,
  {32'hc19bb871, 32'hc1b0865c} /* (24, 0, 3) {real, imag} */,
  {32'hc1966352, 32'hc1e917d2} /* (24, 0, 2) {real, imag} */,
  {32'hc17b5bdd, 32'hc1d28430} /* (24, 0, 1) {real, imag} */,
  {32'hc1a6020b, 32'hc19189cc} /* (24, 0, 0) {real, imag} */,
  {32'hc0313c12, 32'h41038813} /* (23, 31, 31) {real, imag} */,
  {32'hc18ca618, 32'h41ccef3a} /* (23, 31, 30) {real, imag} */,
  {32'hc1d186dc, 32'h3fab3c14} /* (23, 31, 29) {real, imag} */,
  {32'hc11418fd, 32'hc194b3fa} /* (23, 31, 28) {real, imag} */,
  {32'hc14a740e, 32'hc1317c87} /* (23, 31, 27) {real, imag} */,
  {32'hc1788a29, 32'hc07fb8fc} /* (23, 31, 26) {real, imag} */,
  {32'hc1649fae, 32'hc108572e} /* (23, 31, 25) {real, imag} */,
  {32'hc10ec958, 32'hc16183fe} /* (23, 31, 24) {real, imag} */,
  {32'hc0778505, 32'hc1473f13} /* (23, 31, 23) {real, imag} */,
  {32'hc0b82fa7, 32'hbf2b05a0} /* (23, 31, 22) {real, imag} */,
  {32'hc14f3236, 32'h412e4435} /* (23, 31, 21) {real, imag} */,
  {32'hc0d216b2, 32'h41333916} /* (23, 31, 20) {real, imag} */,
  {32'hc06ed5d4, 32'hbfa869b8} /* (23, 31, 19) {real, imag} */,
  {32'h4048a794, 32'h40ce975e} /* (23, 31, 18) {real, imag} */,
  {32'hbfa78718, 32'h409f396a} /* (23, 31, 17) {real, imag} */,
  {32'hc031761a, 32'h3f0909e0} /* (23, 31, 16) {real, imag} */,
  {32'h417adde6, 32'hbe8240b8} /* (23, 31, 15) {real, imag} */,
  {32'h417bbec6, 32'h41346481} /* (23, 31, 14) {real, imag} */,
  {32'h4182ae9e, 32'h4195ab4a} /* (23, 31, 13) {real, imag} */,
  {32'h41519064, 32'h4186f5f7} /* (23, 31, 12) {real, imag} */,
  {32'hbe56ef40, 32'h40e68ade} /* (23, 31, 11) {real, imag} */,
  {32'hc1234931, 32'h41b5451e} /* (23, 31, 10) {real, imag} */,
  {32'hc1a52840, 32'h40c5b639} /* (23, 31, 9) {real, imag} */,
  {32'hc196496f, 32'hc0942218} /* (23, 31, 8) {real, imag} */,
  {32'h3f5f7ad8, 32'hc11e9dda} /* (23, 31, 7) {real, imag} */,
  {32'hbfed1db8, 32'hc185001d} /* (23, 31, 6) {real, imag} */,
  {32'hc193e643, 32'hc08cf9a2} /* (23, 31, 5) {real, imag} */,
  {32'hc12134b5, 32'h3fb69c0c} /* (23, 31, 4) {real, imag} */,
  {32'h4115ec2a, 32'h40ed4ace} /* (23, 31, 3) {real, imag} */,
  {32'h413251b5, 32'h40cad6ef} /* (23, 31, 2) {real, imag} */,
  {32'hc075e1cc, 32'h40075d6c} /* (23, 31, 1) {real, imag} */,
  {32'hc080dc35, 32'h40780294} /* (23, 31, 0) {real, imag} */,
  {32'hc0bce66c, 32'h40d8916f} /* (23, 30, 31) {real, imag} */,
  {32'h40277c26, 32'h41304757} /* (23, 30, 30) {real, imag} */,
  {32'h40e01d0e, 32'h4168902f} /* (23, 30, 29) {real, imag} */,
  {32'h41a47e15, 32'h3ff553c6} /* (23, 30, 28) {real, imag} */,
  {32'h4165d33d, 32'h41815224} /* (23, 30, 27) {real, imag} */,
  {32'h41307932, 32'h41746ba3} /* (23, 30, 26) {real, imag} */,
  {32'hc0e262fc, 32'h41a82618} /* (23, 30, 25) {real, imag} */,
  {32'hc1747dec, 32'h41e06ac6} /* (23, 30, 24) {real, imag} */,
  {32'h402c2f23, 32'h411dc171} /* (23, 30, 23) {real, imag} */,
  {32'hc06c637c, 32'h40d59eb1} /* (23, 30, 22) {real, imag} */,
  {32'hc0ede350, 32'h41134662} /* (23, 30, 21) {real, imag} */,
  {32'hc184b62e, 32'hc14ebb5c} /* (23, 30, 20) {real, imag} */,
  {32'h404615fa, 32'hc191c054} /* (23, 30, 19) {real, imag} */,
  {32'h40866878, 32'hc0e8af7b} /* (23, 30, 18) {real, imag} */,
  {32'hc0d69fbe, 32'hc105885a} /* (23, 30, 17) {real, imag} */,
  {32'h4119e832, 32'hc112f74a} /* (23, 30, 16) {real, imag} */,
  {32'h404d6306, 32'hc0b9ead5} /* (23, 30, 15) {real, imag} */,
  {32'hbfee514c, 32'hbec730c8} /* (23, 30, 14) {real, imag} */,
  {32'hc0c39956, 32'hc0d87095} /* (23, 30, 13) {real, imag} */,
  {32'hc16e655d, 32'hc12ce6aa} /* (23, 30, 12) {real, imag} */,
  {32'hc1187c64, 32'hc17265a7} /* (23, 30, 11) {real, imag} */,
  {32'h410a3c56, 32'h3efc07e6} /* (23, 30, 10) {real, imag} */,
  {32'h403b781c, 32'h4177f134} /* (23, 30, 9) {real, imag} */,
  {32'hc0cd8bac, 32'h42052b86} /* (23, 30, 8) {real, imag} */,
  {32'h4043b7c2, 32'h41d3daab} /* (23, 30, 7) {real, imag} */,
  {32'h4188ce7e, 32'h4157f359} /* (23, 30, 6) {real, imag} */,
  {32'h40f9f60a, 32'hbf9464bc} /* (23, 30, 5) {real, imag} */,
  {32'h404542ec, 32'h3e344d00} /* (23, 30, 4) {real, imag} */,
  {32'h3e72a004, 32'hc090467a} /* (23, 30, 3) {real, imag} */,
  {32'hbee3897c, 32'hc0da7628} /* (23, 30, 2) {real, imag} */,
  {32'h3da6c110, 32'hc06841e4} /* (23, 30, 1) {real, imag} */,
  {32'h4076632a, 32'hc03c6936} /* (23, 30, 0) {real, imag} */,
  {32'h40d1cf94, 32'h408a8ca2} /* (23, 29, 31) {real, imag} */,
  {32'hc0c4e402, 32'h3f79984e} /* (23, 29, 30) {real, imag} */,
  {32'hc1786f35, 32'h3e28f1c0} /* (23, 29, 29) {real, imag} */,
  {32'hc0e58f1e, 32'h401b8763} /* (23, 29, 28) {real, imag} */,
  {32'hc0087e82, 32'hbf77b088} /* (23, 29, 27) {real, imag} */,
  {32'hc123a908, 32'hc0d1e9fd} /* (23, 29, 26) {real, imag} */,
  {32'hbf4a4abc, 32'hbf8717a4} /* (23, 29, 25) {real, imag} */,
  {32'h409bb579, 32'hc0e1779b} /* (23, 29, 24) {real, imag} */,
  {32'h41165d16, 32'hc15da70e} /* (23, 29, 23) {real, imag} */,
  {32'h41638c9b, 32'h408bdea6} /* (23, 29, 22) {real, imag} */,
  {32'h4180c9ac, 32'h40e9d104} /* (23, 29, 21) {real, imag} */,
  {32'h4199d65d, 32'h40ddcc13} /* (23, 29, 20) {real, imag} */,
  {32'h406cfd1f, 32'h3d16d600} /* (23, 29, 19) {real, imag} */,
  {32'hc1016940, 32'h3fdf2c17} /* (23, 29, 18) {real, imag} */,
  {32'h4026ec58, 32'hbece1a40} /* (23, 29, 17) {real, imag} */,
  {32'hc10c3b38, 32'h407f451c} /* (23, 29, 16) {real, imag} */,
  {32'hc0dae0bd, 32'h4130a6ef} /* (23, 29, 15) {real, imag} */,
  {32'hc0a75550, 32'hc0febc80} /* (23, 29, 14) {real, imag} */,
  {32'h40ab0c5c, 32'hc1168f32} /* (23, 29, 13) {real, imag} */,
  {32'h4075aa7c, 32'hbe4bbbe0} /* (23, 29, 12) {real, imag} */,
  {32'h40fd73a6, 32'h41180ca5} /* (23, 29, 11) {real, imag} */,
  {32'h406de0d0, 32'h41069c08} /* (23, 29, 10) {real, imag} */,
  {32'hc0a0cd2a, 32'hc18186c5} /* (23, 29, 9) {real, imag} */,
  {32'h414e57c2, 32'hc19b80e4} /* (23, 29, 8) {real, imag} */,
  {32'h3f17c9c8, 32'hbff3c120} /* (23, 29, 7) {real, imag} */,
  {32'h416cc88d, 32'h3fbc8af0} /* (23, 29, 6) {real, imag} */,
  {32'h413d4e54, 32'h41377717} /* (23, 29, 5) {real, imag} */,
  {32'hc0181172, 32'h403ca85b} /* (23, 29, 4) {real, imag} */,
  {32'h405f6c0b, 32'h410e6aaa} /* (23, 29, 3) {real, imag} */,
  {32'h40cf904f, 32'h40844950} /* (23, 29, 2) {real, imag} */,
  {32'h410643ae, 32'h40472ab0} /* (23, 29, 1) {real, imag} */,
  {32'h410f1f48, 32'h409a0441} /* (23, 29, 0) {real, imag} */,
  {32'hc01ca794, 32'hc0e24aa6} /* (23, 28, 31) {real, imag} */,
  {32'h3f29d508, 32'hc11fed1e} /* (23, 28, 30) {real, imag} */,
  {32'h408e4e3f, 32'h411f09c6} /* (23, 28, 29) {real, imag} */,
  {32'h40ac475b, 32'h413c1cf5} /* (23, 28, 28) {real, imag} */,
  {32'h40771626, 32'hc10e55af} /* (23, 28, 27) {real, imag} */,
  {32'hc1368fa2, 32'hc12c6e1e} /* (23, 28, 26) {real, imag} */,
  {32'hc0d15b62, 32'hc0b09036} /* (23, 28, 25) {real, imag} */,
  {32'h4040279f, 32'h3fb8e170} /* (23, 28, 24) {real, imag} */,
  {32'h41293885, 32'h40448899} /* (23, 28, 23) {real, imag} */,
  {32'h40b5d816, 32'hc111b50d} /* (23, 28, 22) {real, imag} */,
  {32'h3fb69b12, 32'hc16c7621} /* (23, 28, 21) {real, imag} */,
  {32'hc05e43bd, 32'hc0756164} /* (23, 28, 20) {real, imag} */,
  {32'hc13f749c, 32'h41310d5c} /* (23, 28, 19) {real, imag} */,
  {32'hc0b369f8, 32'h41452faa} /* (23, 28, 18) {real, imag} */,
  {32'hc0b1eb32, 32'h41210bc2} /* (23, 28, 17) {real, imag} */,
  {32'hc1298c4b, 32'h40f86870} /* (23, 28, 16) {real, imag} */,
  {32'h3f97354e, 32'hc021dbac} /* (23, 28, 15) {real, imag} */,
  {32'h41b3d1d6, 32'hc00eccc1} /* (23, 28, 14) {real, imag} */,
  {32'h406a9ab1, 32'hc0ab8a3e} /* (23, 28, 13) {real, imag} */,
  {32'hc0a8d120, 32'hc0258bd6} /* (23, 28, 12) {real, imag} */,
  {32'hc0db3a56, 32'hbd769c80} /* (23, 28, 11) {real, imag} */,
  {32'h40ba228f, 32'hbea430f0} /* (23, 28, 10) {real, imag} */,
  {32'h415c47b5, 32'h40f8782d} /* (23, 28, 9) {real, imag} */,
  {32'hc04f4208, 32'hc05b20ac} /* (23, 28, 8) {real, imag} */,
  {32'hc16778b2, 32'hbe08aee0} /* (23, 28, 7) {real, imag} */,
  {32'hc0e2ce79, 32'h413a8604} /* (23, 28, 6) {real, imag} */,
  {32'hc08e8d6a, 32'hbf52e218} /* (23, 28, 5) {real, imag} */,
  {32'hc121dad1, 32'hc0d9c58b} /* (23, 28, 4) {real, imag} */,
  {32'h4106b681, 32'h41198e23} /* (23, 28, 3) {real, imag} */,
  {32'h40f99c36, 32'h409c24a8} /* (23, 28, 2) {real, imag} */,
  {32'h41326c8e, 32'hc10442ce} /* (23, 28, 1) {real, imag} */,
  {32'h409d70ad, 32'hc15067de} /* (23, 28, 0) {real, imag} */,
  {32'hc061c053, 32'h40622e24} /* (23, 27, 31) {real, imag} */,
  {32'h409af520, 32'h401f24da} /* (23, 27, 30) {real, imag} */,
  {32'h3e1072d8, 32'h40cc6f70} /* (23, 27, 29) {real, imag} */,
  {32'h408dc626, 32'h4181b488} /* (23, 27, 28) {real, imag} */,
  {32'h414ce4d4, 32'h40df008d} /* (23, 27, 27) {real, imag} */,
  {32'hc04edb06, 32'h3f8bb588} /* (23, 27, 26) {real, imag} */,
  {32'h3f8a2e88, 32'h400b658e} /* (23, 27, 25) {real, imag} */,
  {32'h40e68ee8, 32'h40f67050} /* (23, 27, 24) {real, imag} */,
  {32'hbe009b00, 32'h40fe92eb} /* (23, 27, 23) {real, imag} */,
  {32'h40e50182, 32'hc056a8f2} /* (23, 27, 22) {real, imag} */,
  {32'hbf8d3fcc, 32'h4052c464} /* (23, 27, 21) {real, imag} */,
  {32'h40362dfa, 32'h3f3993f0} /* (23, 27, 20) {real, imag} */,
  {32'h415b0857, 32'hc12a751e} /* (23, 27, 19) {real, imag} */,
  {32'h40dd78ec, 32'hbe2bb680} /* (23, 27, 18) {real, imag} */,
  {32'hc091242c, 32'h4142b873} /* (23, 27, 17) {real, imag} */,
  {32'hc02fcadb, 32'hc0b1605a} /* (23, 27, 16) {real, imag} */,
  {32'h410e9264, 32'hc08e76c0} /* (23, 27, 15) {real, imag} */,
  {32'h4005caf0, 32'hc1109d4f} /* (23, 27, 14) {real, imag} */,
  {32'h3eda71f0, 32'h3fe56d3a} /* (23, 27, 13) {real, imag} */,
  {32'hc139fe01, 32'h4172ace7} /* (23, 27, 12) {real, imag} */,
  {32'hc173bc30, 32'h41443290} /* (23, 27, 11) {real, imag} */,
  {32'hc0755e5a, 32'h40ce894a} /* (23, 27, 10) {real, imag} */,
  {32'hc0101e8d, 32'hc08e9f86} /* (23, 27, 9) {real, imag} */,
  {32'h3f1de658, 32'h3f39e7f0} /* (23, 27, 8) {real, imag} */,
  {32'h41a9be26, 32'h4005f056} /* (23, 27, 7) {real, imag} */,
  {32'h41434ef7, 32'hc105cea5} /* (23, 27, 6) {real, imag} */,
  {32'h41077c86, 32'hc14d5fbe} /* (23, 27, 5) {real, imag} */,
  {32'h40a7bdd6, 32'h3f5e22b9} /* (23, 27, 4) {real, imag} */,
  {32'h400536e2, 32'h4126f18c} /* (23, 27, 3) {real, imag} */,
  {32'hbff2bea4, 32'h3febae9c} /* (23, 27, 2) {real, imag} */,
  {32'hc07a385c, 32'h3fce7e1b} /* (23, 27, 1) {real, imag} */,
  {32'h406ebb2e, 32'h41769b06} /* (23, 27, 0) {real, imag} */,
  {32'hc0eef87d, 32'hc0a20d74} /* (23, 26, 31) {real, imag} */,
  {32'hbfa7c31c, 32'hc131df98} /* (23, 26, 30) {real, imag} */,
  {32'h4133ff1e, 32'hbe806318} /* (23, 26, 29) {real, imag} */,
  {32'h415d1464, 32'hbf9aac96} /* (23, 26, 28) {real, imag} */,
  {32'h40459191, 32'h3f09dd9e} /* (23, 26, 27) {real, imag} */,
  {32'hc134fa24, 32'h410de181} /* (23, 26, 26) {real, imag} */,
  {32'hc125977f, 32'hbed24b0c} /* (23, 26, 25) {real, imag} */,
  {32'hc08b056e, 32'h40d7e419} /* (23, 26, 24) {real, imag} */,
  {32'hc105fce7, 32'h413e4f1c} /* (23, 26, 23) {real, imag} */,
  {32'hc02852d2, 32'h407ee9d4} /* (23, 26, 22) {real, imag} */,
  {32'hc1172bd4, 32'hc077f9ec} /* (23, 26, 21) {real, imag} */,
  {32'hc15e26f5, 32'hc0833182} /* (23, 26, 20) {real, imag} */,
  {32'hc1017a38, 32'hc0945c3c} /* (23, 26, 19) {real, imag} */,
  {32'hbfd347b0, 32'h3f561790} /* (23, 26, 18) {real, imag} */,
  {32'hbf886968, 32'hc097cfb4} /* (23, 26, 17) {real, imag} */,
  {32'hc1066f14, 32'hc115c802} /* (23, 26, 16) {real, imag} */,
  {32'hc13c0712, 32'hbeca33a0} /* (23, 26, 15) {real, imag} */,
  {32'hc12723d7, 32'hc1114c89} /* (23, 26, 14) {real, imag} */,
  {32'hbf5f2d38, 32'hc0d57d6a} /* (23, 26, 13) {real, imag} */,
  {32'h4076b39e, 32'hbd95e6d0} /* (23, 26, 12) {real, imag} */,
  {32'h3d9b0fc0, 32'hc123cce1} /* (23, 26, 11) {real, imag} */,
  {32'hc01e04ee, 32'hbfb4a3d5} /* (23, 26, 10) {real, imag} */,
  {32'hc153496a, 32'h41050b18} /* (23, 26, 9) {real, imag} */,
  {32'hc0f34ff4, 32'h416f4120} /* (23, 26, 8) {real, imag} */,
  {32'hc113c5f1, 32'h412082da} /* (23, 26, 7) {real, imag} */,
  {32'hc083fa2c, 32'h4075f21a} /* (23, 26, 6) {real, imag} */,
  {32'hc0d4f4ea, 32'hc02be704} /* (23, 26, 5) {real, imag} */,
  {32'h40032a38, 32'hc0237461} /* (23, 26, 4) {real, imag} */,
  {32'h4032ec2e, 32'hc0399398} /* (23, 26, 3) {real, imag} */,
  {32'hbffc348c, 32'h4017aee6} /* (23, 26, 2) {real, imag} */,
  {32'h4115e44c, 32'h3fbc5e62} /* (23, 26, 1) {real, imag} */,
  {32'h411043c8, 32'hc04a9890} /* (23, 26, 0) {real, imag} */,
  {32'h3f8a5466, 32'hc0289d81} /* (23, 25, 31) {real, imag} */,
  {32'hbf84bb47, 32'hc1472527} /* (23, 25, 30) {real, imag} */,
  {32'hc00ab70e, 32'hc13f0c6c} /* (23, 25, 29) {real, imag} */,
  {32'hc1976835, 32'hc02a44fd} /* (23, 25, 28) {real, imag} */,
  {32'hc1244e7c, 32'h408564d3} /* (23, 25, 27) {real, imag} */,
  {32'h4062f10b, 32'h410bedd5} /* (23, 25, 26) {real, imag} */,
  {32'hbf25a3f8, 32'h3fe6bd4c} /* (23, 25, 25) {real, imag} */,
  {32'hc118f585, 32'hc04ce628} /* (23, 25, 24) {real, imag} */,
  {32'hc12940b1, 32'hc09a114c} /* (23, 25, 23) {real, imag} */,
  {32'hc107a519, 32'hc1093d22} /* (23, 25, 22) {real, imag} */,
  {32'h407027f3, 32'hc090965b} /* (23, 25, 21) {real, imag} */,
  {32'hbfbec844, 32'h40849aec} /* (23, 25, 20) {real, imag} */,
  {32'hc0bbfaf5, 32'h41423b86} /* (23, 25, 19) {real, imag} */,
  {32'h41036d31, 32'hc0109904} /* (23, 25, 18) {real, imag} */,
  {32'h408cb4d8, 32'hc1015e85} /* (23, 25, 17) {real, imag} */,
  {32'hbf4dec42, 32'hbf03405a} /* (23, 25, 16) {real, imag} */,
  {32'hc0629bb4, 32'hc13ca7ee} /* (23, 25, 15) {real, imag} */,
  {32'h3fd6aca4, 32'hc165f60a} /* (23, 25, 14) {real, imag} */,
  {32'hc0909364, 32'hc1931cb8} /* (23, 25, 13) {real, imag} */,
  {32'hc160c9d9, 32'hc0c12f4c} /* (23, 25, 12) {real, imag} */,
  {32'hc0a38c44, 32'h40bf83d5} /* (23, 25, 11) {real, imag} */,
  {32'h4095eee7, 32'hc0f5dac9} /* (23, 25, 10) {real, imag} */,
  {32'h40c5003a, 32'hbfd73b70} /* (23, 25, 9) {real, imag} */,
  {32'h3f8c3cb4, 32'h402423a9} /* (23, 25, 8) {real, imag} */,
  {32'h40e4c3b6, 32'h3f12edd6} /* (23, 25, 7) {real, imag} */,
  {32'h40e17361, 32'h3ff52a22} /* (23, 25, 6) {real, imag} */,
  {32'h411e1955, 32'h3e3cac30} /* (23, 25, 5) {real, imag} */,
  {32'hbfabbf22, 32'h40f4460a} /* (23, 25, 4) {real, imag} */,
  {32'hc0b8d53c, 32'h40c27456} /* (23, 25, 3) {real, imag} */,
  {32'h4024eade, 32'hbf76dba0} /* (23, 25, 2) {real, imag} */,
  {32'hc1003c5e, 32'h40f9f986} /* (23, 25, 1) {real, imag} */,
  {32'hc1494644, 32'h4077e543} /* (23, 25, 0) {real, imag} */,
  {32'h40c82d04, 32'hc06e3592} /* (23, 24, 31) {real, imag} */,
  {32'h410fe3de, 32'hc08dadc9} /* (23, 24, 30) {real, imag} */,
  {32'h40a08afe, 32'h411c7bd9} /* (23, 24, 29) {real, imag} */,
  {32'hbfaf5d9c, 32'h41a5466c} /* (23, 24, 28) {real, imag} */,
  {32'hbf5dc9fb, 32'h40ed6a30} /* (23, 24, 27) {real, imag} */,
  {32'h404ccf92, 32'h408c5b37} /* (23, 24, 26) {real, imag} */,
  {32'h402f7885, 32'h4065f5e4} /* (23, 24, 25) {real, imag} */,
  {32'h407ec56a, 32'hc0006176} /* (23, 24, 24) {real, imag} */,
  {32'h41926a1c, 32'h41229f32} /* (23, 24, 23) {real, imag} */,
  {32'h41867fe6, 32'h4154cd28} /* (23, 24, 22) {real, imag} */,
  {32'h40e90433, 32'h405c5008} /* (23, 24, 21) {real, imag} */,
  {32'h4072b10c, 32'h3e9ec110} /* (23, 24, 20) {real, imag} */,
  {32'hc02e2b6c, 32'hbf9562d2} /* (23, 24, 19) {real, imag} */,
  {32'hbf316eaf, 32'hc0413e43} /* (23, 24, 18) {real, imag} */,
  {32'hc058ddf9, 32'hc04a9496} /* (23, 24, 17) {real, imag} */,
  {32'h412a394b, 32'hc03e33f8} /* (23, 24, 16) {real, imag} */,
  {32'h413cff62, 32'hc0c68228} /* (23, 24, 15) {real, imag} */,
  {32'h40ac68fc, 32'hbe898a54} /* (23, 24, 14) {real, imag} */,
  {32'h3fc012dc, 32'h3faeab38} /* (23, 24, 13) {real, imag} */,
  {32'h4046ca9a, 32'hc080dac7} /* (23, 24, 12) {real, imag} */,
  {32'h41293f46, 32'hc032bdd5} /* (23, 24, 11) {real, imag} */,
  {32'h40cf3cd6, 32'hc0c907f7} /* (23, 24, 10) {real, imag} */,
  {32'h3ee52448, 32'hc10c101d} /* (23, 24, 9) {real, imag} */,
  {32'hbf5ad8bc, 32'hbfae01ce} /* (23, 24, 8) {real, imag} */,
  {32'h40db068f, 32'h3ff787bc} /* (23, 24, 7) {real, imag} */,
  {32'h40b0afad, 32'h3dd72a00} /* (23, 24, 6) {real, imag} */,
  {32'h41221528, 32'hc1323e84} /* (23, 24, 5) {real, imag} */,
  {32'h4117721f, 32'hc07ffd52} /* (23, 24, 4) {real, imag} */,
  {32'h40a30ab9, 32'hc08c9ca8} /* (23, 24, 3) {real, imag} */,
  {32'hbf2a233c, 32'h3f6b222e} /* (23, 24, 2) {real, imag} */,
  {32'h40815afa, 32'h4064280a} /* (23, 24, 1) {real, imag} */,
  {32'h3f8148cc, 32'h40341b36} /* (23, 24, 0) {real, imag} */,
  {32'hbf992477, 32'hc055a547} /* (23, 23, 31) {real, imag} */,
  {32'hbf55ba72, 32'h3fbf2616} /* (23, 23, 30) {real, imag} */,
  {32'hbe7d27c4, 32'hc0b1f358} /* (23, 23, 29) {real, imag} */,
  {32'hc0dc7ed0, 32'hc09cba84} /* (23, 23, 28) {real, imag} */,
  {32'hc117e6ad, 32'hc05388ff} /* (23, 23, 27) {real, imag} */,
  {32'hc09ff97a, 32'hbfab4cd5} /* (23, 23, 26) {real, imag} */,
  {32'h40b840ee, 32'h4047ab4f} /* (23, 23, 25) {real, imag} */,
  {32'hc05ac194, 32'hbf4e2a90} /* (23, 23, 24) {real, imag} */,
  {32'hc13c41b1, 32'hc1110561} /* (23, 23, 23) {real, imag} */,
  {32'hc083be36, 32'hbf8d3fbb} /* (23, 23, 22) {real, imag} */,
  {32'hc1069316, 32'hbe617968} /* (23, 23, 21) {real, imag} */,
  {32'hc0163448, 32'hc02cfe7f} /* (23, 23, 20) {real, imag} */,
  {32'h40a280cc, 32'hbfd031c8} /* (23, 23, 19) {real, imag} */,
  {32'h3dae5d30, 32'hbfd94920} /* (23, 23, 18) {real, imag} */,
  {32'h400a28ea, 32'hbedfc248} /* (23, 23, 17) {real, imag} */,
  {32'h40b60fbe, 32'h3fb013f8} /* (23, 23, 16) {real, imag} */,
  {32'h40b73475, 32'h3f2a49b0} /* (23, 23, 15) {real, imag} */,
  {32'h3fe7e428, 32'hc0ea439f} /* (23, 23, 14) {real, imag} */,
  {32'hbca16cc0, 32'hc0e4c88b} /* (23, 23, 13) {real, imag} */,
  {32'h411608f4, 32'hc05f4f5f} /* (23, 23, 12) {real, imag} */,
  {32'h40c263b6, 32'hc00a5178} /* (23, 23, 11) {real, imag} */,
  {32'h3fd6c2e4, 32'h3f37271c} /* (23, 23, 10) {real, imag} */,
  {32'h408b6da0, 32'hc03bad1e} /* (23, 23, 9) {real, imag} */,
  {32'hc0043db0, 32'hc09632a0} /* (23, 23, 8) {real, imag} */,
  {32'hc0ba8b4e, 32'hc1057a06} /* (23, 23, 7) {real, imag} */,
  {32'hbf3ae626, 32'hbe8630c0} /* (23, 23, 6) {real, imag} */,
  {32'hc105af36, 32'h3f4157a4} /* (23, 23, 5) {real, imag} */,
  {32'hc14ff71e, 32'h3ea80008} /* (23, 23, 4) {real, imag} */,
  {32'hbffded70, 32'hc09344c2} /* (23, 23, 3) {real, imag} */,
  {32'h40f65490, 32'hc1208890} /* (23, 23, 2) {real, imag} */,
  {32'h400d859d, 32'hbfddb6b6} /* (23, 23, 1) {real, imag} */,
  {32'hc035e106, 32'h403a2e28} /* (23, 23, 0) {real, imag} */,
  {32'hbf1c745a, 32'hc0bef488} /* (23, 22, 31) {real, imag} */,
  {32'h3f52c5b6, 32'h3f1f6564} /* (23, 22, 30) {real, imag} */,
  {32'h40c568d1, 32'h40a3abbb} /* (23, 22, 29) {real, imag} */,
  {32'h3fb81766, 32'h4085219e} /* (23, 22, 28) {real, imag} */,
  {32'hc01de940, 32'h40e543d1} /* (23, 22, 27) {real, imag} */,
  {32'h4054d430, 32'h401bd826} /* (23, 22, 26) {real, imag} */,
  {32'hc0332e7f, 32'hbfc70701} /* (23, 22, 25) {real, imag} */,
  {32'hbfb1c337, 32'h3efc04b0} /* (23, 22, 24) {real, imag} */,
  {32'hc06f0385, 32'hbfc0d886} /* (23, 22, 23) {real, imag} */,
  {32'hc0e59e10, 32'hc0c6977e} /* (23, 22, 22) {real, imag} */,
  {32'hbf4836f8, 32'hc10335f0} /* (23, 22, 21) {real, imag} */,
  {32'hbf9df58a, 32'hc104b5ae} /* (23, 22, 20) {real, imag} */,
  {32'hbfec734a, 32'hbfa9b0fc} /* (23, 22, 19) {real, imag} */,
  {32'h40fcc059, 32'hc0f1727a} /* (23, 22, 18) {real, imag} */,
  {32'h4098274e, 32'hc1035093} /* (23, 22, 17) {real, imag} */,
  {32'hbf9c79ce, 32'hbf34407c} /* (23, 22, 16) {real, imag} */,
  {32'hc09dd13a, 32'h4081917b} /* (23, 22, 15) {real, imag} */,
  {32'hbf0164f8, 32'h40a9b994} /* (23, 22, 14) {real, imag} */,
  {32'hbfcb3871, 32'h40c7e4b6} /* (23, 22, 13) {real, imag} */,
  {32'hbf93b1b4, 32'h40583780} /* (23, 22, 12) {real, imag} */,
  {32'h3d9cfcc0, 32'h4080804a} /* (23, 22, 11) {real, imag} */,
  {32'hc0b018e3, 32'hbd9dfac0} /* (23, 22, 10) {real, imag} */,
  {32'hc0b25ebc, 32'h3f57bc6e} /* (23, 22, 9) {real, imag} */,
  {32'hc00f6f21, 32'hc075211e} /* (23, 22, 8) {real, imag} */,
  {32'h3fad8650, 32'h3b647400} /* (23, 22, 7) {real, imag} */,
  {32'h4054171c, 32'hc08e668a} /* (23, 22, 6) {real, imag} */,
  {32'h3f1fe136, 32'h3f9f041a} /* (23, 22, 5) {real, imag} */,
  {32'hc037bdd7, 32'hc0d91774} /* (23, 22, 4) {real, imag} */,
  {32'hc105513c, 32'hc0047bd2} /* (23, 22, 3) {real, imag} */,
  {32'hc0c87c7b, 32'h4088759b} /* (23, 22, 2) {real, imag} */,
  {32'h3fc6cc31, 32'hbfade9fe} /* (23, 22, 1) {real, imag} */,
  {32'h4084d93c, 32'hbe6cfbd4} /* (23, 22, 0) {real, imag} */,
  {32'h404202cc, 32'h40297ae4} /* (23, 21, 31) {real, imag} */,
  {32'hc0604ee0, 32'h4100eaeb} /* (23, 21, 30) {real, imag} */,
  {32'h4025d6ac, 32'h40ae2e0d} /* (23, 21, 29) {real, imag} */,
  {32'h410fd32c, 32'h3fe933da} /* (23, 21, 28) {real, imag} */,
  {32'h40e83356, 32'hc0a7fab8} /* (23, 21, 27) {real, imag} */,
  {32'hbfd09e0a, 32'hc0b67f89} /* (23, 21, 26) {real, imag} */,
  {32'hbfbf0ba3, 32'h3fdb005e} /* (23, 21, 25) {real, imag} */,
  {32'hbfd23cbe, 32'h41364e7c} /* (23, 21, 24) {real, imag} */,
  {32'hbfe6afac, 32'h400712e2} /* (23, 21, 23) {real, imag} */,
  {32'hc0ae15ce, 32'hc048bfa2} /* (23, 21, 22) {real, imag} */,
  {32'hc0fcd0b8, 32'hbf9dbb6e} /* (23, 21, 21) {real, imag} */,
  {32'hc0cbc32e, 32'hbff743cc} /* (23, 21, 20) {real, imag} */,
  {32'h4013db7e, 32'hc0ccf548} /* (23, 21, 19) {real, imag} */,
  {32'hbf79c571, 32'h4062fb4a} /* (23, 21, 18) {real, imag} */,
  {32'hbf212d3e, 32'h40e13243} /* (23, 21, 17) {real, imag} */,
  {32'h40319c0d, 32'h3f80601a} /* (23, 21, 16) {real, imag} */,
  {32'hc03ffe12, 32'h3dc903b8} /* (23, 21, 15) {real, imag} */,
  {32'hc0a5d01f, 32'hbfbc2e51} /* (23, 21, 14) {real, imag} */,
  {32'hc085af3e, 32'hc042d9e1} /* (23, 21, 13) {real, imag} */,
  {32'hc0733eed, 32'hc0a08858} /* (23, 21, 12) {real, imag} */,
  {32'hc085909d, 32'hbfad81a5} /* (23, 21, 11) {real, imag} */,
  {32'h3faad6a0, 32'hc04b199e} /* (23, 21, 10) {real, imag} */,
  {32'hbf2683b4, 32'hc075ee14} /* (23, 21, 9) {real, imag} */,
  {32'h3f34f318, 32'hc0824348} /* (23, 21, 8) {real, imag} */,
  {32'hbff2f510, 32'hc05545fa} /* (23, 21, 7) {real, imag} */,
  {32'hc0764d53, 32'h4032d9f5} /* (23, 21, 6) {real, imag} */,
  {32'h4052820a, 32'h3e5f2960} /* (23, 21, 5) {real, imag} */,
  {32'h3ef2c18c, 32'hc0240faa} /* (23, 21, 4) {real, imag} */,
  {32'hc0fd098c, 32'h3fc4470a} /* (23, 21, 3) {real, imag} */,
  {32'hc1013702, 32'hbe976c50} /* (23, 21, 2) {real, imag} */,
  {32'hc0f1f4a4, 32'hc10c69e4} /* (23, 21, 1) {real, imag} */,
  {32'h3fe910fb, 32'hc0f73b06} /* (23, 21, 0) {real, imag} */,
  {32'hc03e8d7f, 32'h40278e7c} /* (23, 20, 31) {real, imag} */,
  {32'h3f907d5c, 32'h40922666} /* (23, 20, 30) {real, imag} */,
  {32'h3f28967e, 32'hbf9f6433} /* (23, 20, 29) {real, imag} */,
  {32'hbfc02615, 32'hbef933a4} /* (23, 20, 28) {real, imag} */,
  {32'h4014a004, 32'hbf40614e} /* (23, 20, 27) {real, imag} */,
  {32'hbf57bfaa, 32'h406b94bf} /* (23, 20, 26) {real, imag} */,
  {32'hc01f9959, 32'h40318b86} /* (23, 20, 25) {real, imag} */,
  {32'hc0261be6, 32'h3e7d5ec0} /* (23, 20, 24) {real, imag} */,
  {32'hc0840f8a, 32'hc05cfa00} /* (23, 20, 23) {real, imag} */,
  {32'hc0bfba3a, 32'hc018c1a3} /* (23, 20, 22) {real, imag} */,
  {32'hc0d343d9, 32'hbf880f0c} /* (23, 20, 21) {real, imag} */,
  {32'hc10e7710, 32'hbebab7d4} /* (23, 20, 20) {real, imag} */,
  {32'hbff08ef6, 32'h403428be} /* (23, 20, 19) {real, imag} */,
  {32'h3f9ec190, 32'h401735f9} /* (23, 20, 18) {real, imag} */,
  {32'hbfc14904, 32'hc02291da} /* (23, 20, 17) {real, imag} */,
  {32'hc019449f, 32'hc090d874} /* (23, 20, 16) {real, imag} */,
  {32'h3fbb4969, 32'hc052a9b4} /* (23, 20, 15) {real, imag} */,
  {32'hc050527e, 32'h407602b4} /* (23, 20, 14) {real, imag} */,
  {32'hc0171edb, 32'h40c4b274} /* (23, 20, 13) {real, imag} */,
  {32'h402c6404, 32'h3f82b0f3} /* (23, 20, 12) {real, imag} */,
  {32'hc02ce888, 32'hbfdc8498} /* (23, 20, 11) {real, imag} */,
  {32'hc0dcb6ba, 32'h3f29ba0e} /* (23, 20, 10) {real, imag} */,
  {32'h3fe373df, 32'h3f779490} /* (23, 20, 9) {real, imag} */,
  {32'h401758f0, 32'hbf45ca48} /* (23, 20, 8) {real, imag} */,
  {32'h40229c35, 32'hbf42ebce} /* (23, 20, 7) {real, imag} */,
  {32'hbf3ca227, 32'hbfc211bd} /* (23, 20, 6) {real, imag} */,
  {32'h4080b8b0, 32'h3f5ea046} /* (23, 20, 5) {real, imag} */,
  {32'h40548073, 32'hbfa1b021} /* (23, 20, 4) {real, imag} */,
  {32'h4068bce4, 32'hc0310e6e} /* (23, 20, 3) {real, imag} */,
  {32'h4017f444, 32'hc078cb3b} /* (23, 20, 2) {real, imag} */,
  {32'h3f8b5e4e, 32'hc09d9d2e} /* (23, 20, 1) {real, imag} */,
  {32'h3fe40e31, 32'hc0652d8e} /* (23, 20, 0) {real, imag} */,
  {32'h4008c41f, 32'h3f831e2e} /* (23, 19, 31) {real, imag} */,
  {32'h3ea0a448, 32'hbe7a6e88} /* (23, 19, 30) {real, imag} */,
  {32'hc01e24f5, 32'h3f85bd42} /* (23, 19, 29) {real, imag} */,
  {32'hc08e8a24, 32'hbfb10002} /* (23, 19, 28) {real, imag} */,
  {32'hc08fe5b4, 32'hc0a1e735} /* (23, 19, 27) {real, imag} */,
  {32'hc049516f, 32'hbf891076} /* (23, 19, 26) {real, imag} */,
  {32'hbf46d984, 32'hc02aadd1} /* (23, 19, 25) {real, imag} */,
  {32'h40b9acb4, 32'hbfbe9a28} /* (23, 19, 24) {real, imag} */,
  {32'h40c3eee2, 32'h3edc5540} /* (23, 19, 23) {real, imag} */,
  {32'h3f1eb0a4, 32'hbe7979f0} /* (23, 19, 22) {real, imag} */,
  {32'h3e3d8450, 32'h3fcd8026} /* (23, 19, 21) {real, imag} */,
  {32'hbf7f27f8, 32'h40312864} /* (23, 19, 20) {real, imag} */,
  {32'hc067c173, 32'hbffb391c} /* (23, 19, 19) {real, imag} */,
  {32'h3f8ec740, 32'hc09f6252} /* (23, 19, 18) {real, imag} */,
  {32'h3f15a800, 32'hbfaea724} /* (23, 19, 17) {real, imag} */,
  {32'h404d79b8, 32'h402d6cc7} /* (23, 19, 16) {real, imag} */,
  {32'h40fa68bc, 32'h3fa2367c} /* (23, 19, 15) {real, imag} */,
  {32'h402631ea, 32'h4007515c} /* (23, 19, 14) {real, imag} */,
  {32'h3fb74e40, 32'hbf223160} /* (23, 19, 13) {real, imag} */,
  {32'hbf259780, 32'hc04baa38} /* (23, 19, 12) {real, imag} */,
  {32'hc05dbcec, 32'hc01397ea} /* (23, 19, 11) {real, imag} */,
  {32'hbfa2883b, 32'hc08943d1} /* (23, 19, 10) {real, imag} */,
  {32'hbe517c30, 32'h3fba4b54} /* (23, 19, 9) {real, imag} */,
  {32'hc041492a, 32'h408e3f18} /* (23, 19, 8) {real, imag} */,
  {32'hc007e5a1, 32'h3faae08a} /* (23, 19, 7) {real, imag} */,
  {32'hbe5f5f00, 32'hbf0b41c4} /* (23, 19, 6) {real, imag} */,
  {32'h3f4b9ed4, 32'h400a68ec} /* (23, 19, 5) {real, imag} */,
  {32'hbf918500, 32'h406784e4} /* (23, 19, 4) {real, imag} */,
  {32'h3fbf75ce, 32'h3f949fd1} /* (23, 19, 3) {real, imag} */,
  {32'h3f00512e, 32'h40076cca} /* (23, 19, 2) {real, imag} */,
  {32'hc08c3dda, 32'h40cd06cc} /* (23, 19, 1) {real, imag} */,
  {32'hbf7ad3d4, 32'h40475651} /* (23, 19, 0) {real, imag} */,
  {32'h4001a1ea, 32'hc0107e58} /* (23, 18, 31) {real, imag} */,
  {32'h3f542334, 32'hbfc5dace} /* (23, 18, 30) {real, imag} */,
  {32'hbde3ef80, 32'h3efcc530} /* (23, 18, 29) {real, imag} */,
  {32'hbf8c372a, 32'h402014fe} /* (23, 18, 28) {real, imag} */,
  {32'hc0303213, 32'h3f0e3b50} /* (23, 18, 27) {real, imag} */,
  {32'h3fdb6a7c, 32'hc013e2dd} /* (23, 18, 26) {real, imag} */,
  {32'h40f064df, 32'hc09650fe} /* (23, 18, 25) {real, imag} */,
  {32'h4095d2ba, 32'hc09e5cac} /* (23, 18, 24) {real, imag} */,
  {32'hbf2ac589, 32'hc081377e} /* (23, 18, 23) {real, imag} */,
  {32'hbff34bd6, 32'hc07d36de} /* (23, 18, 22) {real, imag} */,
  {32'hbd458d20, 32'hc00d0c34} /* (23, 18, 21) {real, imag} */,
  {32'hbf28ae28, 32'h403eee1a} /* (23, 18, 20) {real, imag} */,
  {32'hbfaa5058, 32'h408f14b1} /* (23, 18, 19) {real, imag} */,
  {32'hc01d687d, 32'h3e56ce38} /* (23, 18, 18) {real, imag} */,
  {32'h40145794, 32'hbfebb778} /* (23, 18, 17) {real, imag} */,
  {32'h400b0d6c, 32'hc052f64a} /* (23, 18, 16) {real, imag} */,
  {32'hbff5e230, 32'h3ee78d18} /* (23, 18, 15) {real, imag} */,
  {32'hc06955a4, 32'h3fd1b398} /* (23, 18, 14) {real, imag} */,
  {32'hc05b05fd, 32'h3f170996} /* (23, 18, 13) {real, imag} */,
  {32'h3ecd3cc8, 32'h3ff923fc} /* (23, 18, 12) {real, imag} */,
  {32'hbf18427c, 32'h401cf548} /* (23, 18, 11) {real, imag} */,
  {32'hbfb7983a, 32'hbf634401} /* (23, 18, 10) {real, imag} */,
  {32'h3fc2122e, 32'hc01c59ca} /* (23, 18, 9) {real, imag} */,
  {32'h400e4b5a, 32'hc0043ac8} /* (23, 18, 8) {real, imag} */,
  {32'h40293fe6, 32'hbede7660} /* (23, 18, 7) {real, imag} */,
  {32'h405272aa, 32'hbc282800} /* (23, 18, 6) {real, imag} */,
  {32'hbfaf48aa, 32'h40662bc9} /* (23, 18, 5) {real, imag} */,
  {32'hc092cb0e, 32'h400bd522} /* (23, 18, 4) {real, imag} */,
  {32'hc007a129, 32'hc0371941} /* (23, 18, 3) {real, imag} */,
  {32'hbe511a10, 32'hc0a44230} /* (23, 18, 2) {real, imag} */,
  {32'hc07387a6, 32'hc0b5dfd0} /* (23, 18, 1) {real, imag} */,
  {32'hc06ecc4e, 32'hc04598e9} /* (23, 18, 0) {real, imag} */,
  {32'hbfe7f57e, 32'hbfddb97f} /* (23, 17, 31) {real, imag} */,
  {32'h3dc75b60, 32'hc0861f7c} /* (23, 17, 30) {real, imag} */,
  {32'hbfad7c00, 32'hc0453d43} /* (23, 17, 29) {real, imag} */,
  {32'h3feb7430, 32'h3f7dff20} /* (23, 17, 28) {real, imag} */,
  {32'h3efa8898, 32'h4038841b} /* (23, 17, 27) {real, imag} */,
  {32'hbfe5128a, 32'hbfd0504a} /* (23, 17, 26) {real, imag} */,
  {32'h3fcd938b, 32'hbf32540e} /* (23, 17, 25) {real, imag} */,
  {32'hbd351e00, 32'h3ff0dc3b} /* (23, 17, 24) {real, imag} */,
  {32'h3fbfd109, 32'h3fded2d8} /* (23, 17, 23) {real, imag} */,
  {32'h40204488, 32'h401b600c} /* (23, 17, 22) {real, imag} */,
  {32'h407cd4cf, 32'hbdc5c790} /* (23, 17, 21) {real, imag} */,
  {32'h404fef16, 32'hc08477ea} /* (23, 17, 20) {real, imag} */,
  {32'h4005aa68, 32'hbe89de90} /* (23, 17, 19) {real, imag} */,
  {32'hbfd2a0e1, 32'h3fd5453e} /* (23, 17, 18) {real, imag} */,
  {32'hbffc299f, 32'hbf3b4f80} /* (23, 17, 17) {real, imag} */,
  {32'hbf25527c, 32'h3fe53f60} /* (23, 17, 16) {real, imag} */,
  {32'h4032ae96, 32'h3f55cf4c} /* (23, 17, 15) {real, imag} */,
  {32'h3f95a011, 32'h3f53fe08} /* (23, 17, 14) {real, imag} */,
  {32'h4059a3a7, 32'h3f263180} /* (23, 17, 13) {real, imag} */,
  {32'h406f0375, 32'h3f952d98} /* (23, 17, 12) {real, imag} */,
  {32'hbe9af488, 32'h3f360a66} /* (23, 17, 11) {real, imag} */,
  {32'hbf31f758, 32'hbe8176d8} /* (23, 17, 10) {real, imag} */,
  {32'hbf384318, 32'h3fd30509} /* (23, 17, 9) {real, imag} */,
  {32'hbf166c78, 32'h4071fbd6} /* (23, 17, 8) {real, imag} */,
  {32'hbff8f5b2, 32'h3ffcf334} /* (23, 17, 7) {real, imag} */,
  {32'hc04ef184, 32'h3ecd6c74} /* (23, 17, 6) {real, imag} */,
  {32'hbf854a96, 32'hbfa14e66} /* (23, 17, 5) {real, imag} */,
  {32'hbf24d746, 32'h3f99ae42} /* (23, 17, 4) {real, imag} */,
  {32'h3fa8d358, 32'h4004267f} /* (23, 17, 3) {real, imag} */,
  {32'h401f5cb4, 32'h3f94e7e9} /* (23, 17, 2) {real, imag} */,
  {32'hbf63bdc8, 32'hc007aeea} /* (23, 17, 1) {real, imag} */,
  {32'hbf98b91d, 32'hbfc85bff} /* (23, 17, 0) {real, imag} */,
  {32'h400bb95b, 32'h3e839990} /* (23, 16, 31) {real, imag} */,
  {32'hbf57ab40, 32'h4032b94f} /* (23, 16, 30) {real, imag} */,
  {32'hc011ff1c, 32'hbfe215b4} /* (23, 16, 29) {real, imag} */,
  {32'h3f2b4da0, 32'hbf15e240} /* (23, 16, 28) {real, imag} */,
  {32'h403a735b, 32'hbfac2836} /* (23, 16, 27) {real, imag} */,
  {32'h407d7ee6, 32'h3ec4448c} /* (23, 16, 26) {real, imag} */,
  {32'h4008ad16, 32'h40318640} /* (23, 16, 25) {real, imag} */,
  {32'hc05288bc, 32'h4026c0ec} /* (23, 16, 24) {real, imag} */,
  {32'hbf81b078, 32'h408d88dd} /* (23, 16, 23) {real, imag} */,
  {32'h3e8ac5f8, 32'h3ff931e0} /* (23, 16, 22) {real, imag} */,
  {32'hbfcb1846, 32'h3f81dbb6} /* (23, 16, 21) {real, imag} */,
  {32'h3fa885ec, 32'h3fc7c750} /* (23, 16, 20) {real, imag} */,
  {32'h4039daaa, 32'h403eba0a} /* (23, 16, 19) {real, imag} */,
  {32'h3f02beb0, 32'h408a5d6d} /* (23, 16, 18) {real, imag} */,
  {32'h3fd3e9fc, 32'h4026f82a} /* (23, 16, 17) {real, imag} */,
  {32'hbf4819a8, 32'h3e7b11e0} /* (23, 16, 16) {real, imag} */,
  {32'hbf48f880, 32'h3fc83316} /* (23, 16, 15) {real, imag} */,
  {32'h3e25b050, 32'h3fe898bc} /* (23, 16, 14) {real, imag} */,
  {32'hc01cb2f6, 32'h3fccc250} /* (23, 16, 13) {real, imag} */,
  {32'hbf78d790, 32'h401a0642} /* (23, 16, 12) {real, imag} */,
  {32'h3fa8c9e0, 32'hbd4d4400} /* (23, 16, 11) {real, imag} */,
  {32'hbf48ba32, 32'hbf5409f0} /* (23, 16, 10) {real, imag} */,
  {32'h3f4395e8, 32'hc02c93e4} /* (23, 16, 9) {real, imag} */,
  {32'h4029c2b8, 32'h3fd4fa89} /* (23, 16, 8) {real, imag} */,
  {32'h3edbb000, 32'h3eda0078} /* (23, 16, 7) {real, imag} */,
  {32'hbf2950d0, 32'hbe10af18} /* (23, 16, 6) {real, imag} */,
  {32'hc0283956, 32'hbf1d7ef0} /* (23, 16, 5) {real, imag} */,
  {32'hbe2b2e90, 32'h3ee26cd8} /* (23, 16, 4) {real, imag} */,
  {32'h3f4fae24, 32'h3f3c9668} /* (23, 16, 3) {real, imag} */,
  {32'hbf081b0e, 32'h3fea1f20} /* (23, 16, 2) {real, imag} */,
  {32'h4015bffa, 32'hbeb68d80} /* (23, 16, 1) {real, imag} */,
  {32'h4012d785, 32'hbf2bf87c} /* (23, 16, 0) {real, imag} */,
  {32'hbf8362ca, 32'h3ed1eca4} /* (23, 15, 31) {real, imag} */,
  {32'hbfbbcbf6, 32'h40420d17} /* (23, 15, 30) {real, imag} */,
  {32'h40053c20, 32'h3fb6209a} /* (23, 15, 29) {real, imag} */,
  {32'h4018a93e, 32'hbeef6b00} /* (23, 15, 28) {real, imag} */,
  {32'hbd956ee0, 32'hbf5c20ac} /* (23, 15, 27) {real, imag} */,
  {32'hc02fa0dd, 32'h3f481624} /* (23, 15, 26) {real, imag} */,
  {32'h3ff1f695, 32'hbdef4b90} /* (23, 15, 25) {real, imag} */,
  {32'h3f2bb060, 32'hbff5eb03} /* (23, 15, 24) {real, imag} */,
  {32'hbfe8f0f7, 32'h3d547800} /* (23, 15, 23) {real, imag} */,
  {32'hbf963517, 32'h3fdcdf20} /* (23, 15, 22) {real, imag} */,
  {32'h400e7691, 32'h4066b52e} /* (23, 15, 21) {real, imag} */,
  {32'h3d334880, 32'h3eccf460} /* (23, 15, 20) {real, imag} */,
  {32'h3fa3133d, 32'hc0a11058} /* (23, 15, 19) {real, imag} */,
  {32'h3fa868bd, 32'hbfa22816} /* (23, 15, 18) {real, imag} */,
  {32'hbf9dcc5f, 32'h408e19b7} /* (23, 15, 17) {real, imag} */,
  {32'h3e75e3b0, 32'h40762e78} /* (23, 15, 16) {real, imag} */,
  {32'h3f9e000c, 32'h40aaf18a} /* (23, 15, 15) {real, imag} */,
  {32'h3f0505ce, 32'h401e4eee} /* (23, 15, 14) {real, imag} */,
  {32'h402854b9, 32'hbf724240} /* (23, 15, 13) {real, imag} */,
  {32'h400a9933, 32'hbfd47368} /* (23, 15, 12) {real, imag} */,
  {32'h3e8a3608, 32'hc03afdd8} /* (23, 15, 11) {real, imag} */,
  {32'h3fd78b2c, 32'hc00ebb3b} /* (23, 15, 10) {real, imag} */,
  {32'h3faa1a64, 32'hc000b112} /* (23, 15, 9) {real, imag} */,
  {32'h40930beb, 32'hc093ec79} /* (23, 15, 8) {real, imag} */,
  {32'h405d17c5, 32'hc07ef8fa} /* (23, 15, 7) {real, imag} */,
  {32'hbfe48b38, 32'h3f948453} /* (23, 15, 6) {real, imag} */,
  {32'hbfd9e0c2, 32'h3fecb106} /* (23, 15, 5) {real, imag} */,
  {32'h3fca6d3b, 32'hbfabcae2} /* (23, 15, 4) {real, imag} */,
  {32'h40740d10, 32'hbff50812} /* (23, 15, 3) {real, imag} */,
  {32'h3ec8d31c, 32'h3f6bb892} /* (23, 15, 2) {real, imag} */,
  {32'h403cc364, 32'h4008e1fe} /* (23, 15, 1) {real, imag} */,
  {32'h400f2f02, 32'h3e9ad704} /* (23, 15, 0) {real, imag} */,
  {32'hbf07dfc0, 32'hbfc6d0dc} /* (23, 14, 31) {real, imag} */,
  {32'h40854d9c, 32'h3ee79c46} /* (23, 14, 30) {real, imag} */,
  {32'h4058647c, 32'h404e817e} /* (23, 14, 29) {real, imag} */,
  {32'hc02b7917, 32'hbef086c0} /* (23, 14, 28) {real, imag} */,
  {32'hc0157753, 32'hc08e7987} /* (23, 14, 27) {real, imag} */,
  {32'hbe1dc6e0, 32'hc05945b9} /* (23, 14, 26) {real, imag} */,
  {32'h3ebe2aa0, 32'hbf43478c} /* (23, 14, 25) {real, imag} */,
  {32'hc007e7ac, 32'hbf820d60} /* (23, 14, 24) {real, imag} */,
  {32'hbf840270, 32'hbfaf7d22} /* (23, 14, 23) {real, imag} */,
  {32'h4030732d, 32'hc016e65a} /* (23, 14, 22) {real, imag} */,
  {32'h3f08ddb2, 32'hbf3b728a} /* (23, 14, 21) {real, imag} */,
  {32'h3e9edf90, 32'h4013ec2a} /* (23, 14, 20) {real, imag} */,
  {32'h3d583b00, 32'h3faa7134} /* (23, 14, 19) {real, imag} */,
  {32'hbfe1ee3e, 32'h405419a2} /* (23, 14, 18) {real, imag} */,
  {32'hbf57f268, 32'h40df156a} /* (23, 14, 17) {real, imag} */,
  {32'h3f8563a7, 32'h40793e06} /* (23, 14, 16) {real, imag} */,
  {32'hbff42f68, 32'h4085aee8} /* (23, 14, 15) {real, imag} */,
  {32'h3ed549cc, 32'h3f5291f0} /* (23, 14, 14) {real, imag} */,
  {32'h3fd6b66e, 32'hc057a2c2} /* (23, 14, 13) {real, imag} */,
  {32'h3d2e25c0, 32'h3f096708} /* (23, 14, 12) {real, imag} */,
  {32'h404f92a7, 32'hbef18d00} /* (23, 14, 11) {real, imag} */,
  {32'h3ff0269e, 32'h3f48759f} /* (23, 14, 10) {real, imag} */,
  {32'h3da66ba0, 32'h3ccd3ec0} /* (23, 14, 9) {real, imag} */,
  {32'hc05442fa, 32'hc00b2948} /* (23, 14, 8) {real, imag} */,
  {32'hbfb7172c, 32'hbfd8fc38} /* (23, 14, 7) {real, imag} */,
  {32'h4019ebb6, 32'h3f5fe4d0} /* (23, 14, 6) {real, imag} */,
  {32'h40450061, 32'h3fec54e6} /* (23, 14, 5) {real, imag} */,
  {32'h3f0352cc, 32'h405e1cc6} /* (23, 14, 4) {real, imag} */,
  {32'hbd1c4f40, 32'h3da7d620} /* (23, 14, 3) {real, imag} */,
  {32'hc03df7ce, 32'hbf84b022} /* (23, 14, 2) {real, imag} */,
  {32'hbf95c4bb, 32'hbdc96200} /* (23, 14, 1) {real, imag} */,
  {32'h3f080202, 32'h3e85a8b8} /* (23, 14, 0) {real, imag} */,
  {32'hc055dc0d, 32'h3f0a122c} /* (23, 13, 31) {real, imag} */,
  {32'hc02a28a9, 32'h404b2424} /* (23, 13, 30) {real, imag} */,
  {32'hbe6191d0, 32'h40e37bb8} /* (23, 13, 29) {real, imag} */,
  {32'h3d277880, 32'h406492a1} /* (23, 13, 28) {real, imag} */,
  {32'h401093f1, 32'h3ffbef0b} /* (23, 13, 27) {real, imag} */,
  {32'hc0a8c3a8, 32'h3e5b989c} /* (23, 13, 26) {real, imag} */,
  {32'hc0091b3d, 32'h401d1d7b} /* (23, 13, 25) {real, imag} */,
  {32'hbf81081c, 32'h4067cae6} /* (23, 13, 24) {real, imag} */,
  {32'hc0914f7e, 32'h403eb100} /* (23, 13, 23) {real, imag} */,
  {32'hc0968328, 32'h401f7fa5} /* (23, 13, 22) {real, imag} */,
  {32'h3fc7e20e, 32'h3fea50ae} /* (23, 13, 21) {real, imag} */,
  {32'h3fc79f04, 32'hbf81d261} /* (23, 13, 20) {real, imag} */,
  {32'h3fb846aa, 32'hc02de0d8} /* (23, 13, 19) {real, imag} */,
  {32'h40260d90, 32'hbed84d28} /* (23, 13, 18) {real, imag} */,
  {32'hc00273cc, 32'h409f5940} /* (23, 13, 17) {real, imag} */,
  {32'hc09e3c58, 32'h405ac621} /* (23, 13, 16) {real, imag} */,
  {32'hc0b4e386, 32'h3fecacc4} /* (23, 13, 15) {real, imag} */,
  {32'hc09543e3, 32'h40625c1c} /* (23, 13, 14) {real, imag} */,
  {32'hbfd62290, 32'hbfa5aa30} /* (23, 13, 13) {real, imag} */,
  {32'h3f4788a0, 32'hbfdbbb64} /* (23, 13, 12) {real, imag} */,
  {32'hbf196f1e, 32'hbe813dc0} /* (23, 13, 11) {real, imag} */,
  {32'h3fecdd4b, 32'h401b989e} /* (23, 13, 10) {real, imag} */,
  {32'h3f819c8a, 32'h4017ff46} /* (23, 13, 9) {real, imag} */,
  {32'h400bdcb2, 32'h40603fe3} /* (23, 13, 8) {real, imag} */,
  {32'hbecfca58, 32'h3fb43fd6} /* (23, 13, 7) {real, imag} */,
  {32'hc0846744, 32'h402acbd7} /* (23, 13, 6) {real, imag} */,
  {32'hbe89efc8, 32'h3fa78158} /* (23, 13, 5) {real, imag} */,
  {32'h3fbbb444, 32'hbda14930} /* (23, 13, 4) {real, imag} */,
  {32'hc03011d7, 32'h403c6d44} /* (23, 13, 3) {real, imag} */,
  {32'h400c00d2, 32'h408ac110} /* (23, 13, 2) {real, imag} */,
  {32'h3d706500, 32'h40901eda} /* (23, 13, 1) {real, imag} */,
  {32'hc0030125, 32'h40575cd7} /* (23, 13, 0) {real, imag} */,
  {32'hbfbe8d02, 32'h4026d57a} /* (23, 12, 31) {real, imag} */,
  {32'hbf6760e0, 32'hbfde9bb8} /* (23, 12, 30) {real, imag} */,
  {32'h3fa4836f, 32'hc082bca5} /* (23, 12, 29) {real, imag} */,
  {32'hbfa4dfb1, 32'hc0132920} /* (23, 12, 28) {real, imag} */,
  {32'hbf867fbc, 32'hc01cff98} /* (23, 12, 27) {real, imag} */,
  {32'hbf9ca73d, 32'hc03dfe45} /* (23, 12, 26) {real, imag} */,
  {32'hbefd6f78, 32'h3ec45eb0} /* (23, 12, 25) {real, imag} */,
  {32'h3f4949ba, 32'h4039e90e} /* (23, 12, 24) {real, imag} */,
  {32'h408f8f2a, 32'hbf03e746} /* (23, 12, 23) {real, imag} */,
  {32'h3ed6f040, 32'h3fbbd662} /* (23, 12, 22) {real, imag} */,
  {32'hc066ca5e, 32'h4062c478} /* (23, 12, 21) {real, imag} */,
  {32'h3f3d9180, 32'h3f6fd9ee} /* (23, 12, 20) {real, imag} */,
  {32'hbf9189a2, 32'h40027af0} /* (23, 12, 19) {real, imag} */,
  {32'hc00a78b4, 32'hc074635f} /* (23, 12, 18) {real, imag} */,
  {32'hbec3c098, 32'hc097c365} /* (23, 12, 17) {real, imag} */,
  {32'h40bac600, 32'h3f85189e} /* (23, 12, 16) {real, imag} */,
  {32'h4022def2, 32'hbfe6320b} /* (23, 12, 15) {real, imag} */,
  {32'hc07214e6, 32'hc04693ba} /* (23, 12, 14) {real, imag} */,
  {32'h3fba87f6, 32'hc012ade8} /* (23, 12, 13) {real, imag} */,
  {32'hbfddaff8, 32'h3f9d8217} /* (23, 12, 12) {real, imag} */,
  {32'h3f1512e8, 32'h40b7bad2} /* (23, 12, 11) {real, imag} */,
  {32'h40563d80, 32'h3f2ac986} /* (23, 12, 10) {real, imag} */,
  {32'hbf3e3b32, 32'hc0959d46} /* (23, 12, 9) {real, imag} */,
  {32'h3f889cf4, 32'hc0bed81b} /* (23, 12, 8) {real, imag} */,
  {32'h3fec2aae, 32'hbfc540c9} /* (23, 12, 7) {real, imag} */,
  {32'h4025da4e, 32'h3fd10d29} /* (23, 12, 6) {real, imag} */,
  {32'h40d4b506, 32'h3fcf864b} /* (23, 12, 5) {real, imag} */,
  {32'h3ee10d08, 32'h4004a0aa} /* (23, 12, 4) {real, imag} */,
  {32'hc00faa08, 32'h40b4af39} /* (23, 12, 3) {real, imag} */,
  {32'h40d3b98a, 32'h3ff92392} /* (23, 12, 2) {real, imag} */,
  {32'h409276b8, 32'h3fb93c08} /* (23, 12, 1) {real, imag} */,
  {32'hbecf47dc, 32'h3f9e4be0} /* (23, 12, 0) {real, imag} */,
  {32'h3d4a6f80, 32'h3e458798} /* (23, 11, 31) {real, imag} */,
  {32'hbfcf7cb8, 32'hbf4c99fc} /* (23, 11, 30) {real, imag} */,
  {32'hc031e27e, 32'hc0171adc} /* (23, 11, 29) {real, imag} */,
  {32'h408b111e, 32'h3e4228b0} /* (23, 11, 28) {real, imag} */,
  {32'h40db90ee, 32'hc0112460} /* (23, 11, 27) {real, imag} */,
  {32'h40210c91, 32'h40260c5e} /* (23, 11, 26) {real, imag} */,
  {32'hc0772e4a, 32'h3d28fe10} /* (23, 11, 25) {real, imag} */,
  {32'hc0613f7f, 32'h3e899ec0} /* (23, 11, 24) {real, imag} */,
  {32'h3e273180, 32'h4087bf03} /* (23, 11, 23) {real, imag} */,
  {32'hc03186f5, 32'h3f651dc8} /* (23, 11, 22) {real, imag} */,
  {32'hbfed7950, 32'hc040ae37} /* (23, 11, 21) {real, imag} */,
  {32'h3facf76e, 32'hc0f4d451} /* (23, 11, 20) {real, imag} */,
  {32'hbfab202d, 32'hc0399027} /* (23, 11, 19) {real, imag} */,
  {32'hc0132854, 32'h406a2b18} /* (23, 11, 18) {real, imag} */,
  {32'hc0378688, 32'h40bfb899} /* (23, 11, 17) {real, imag} */,
  {32'h4005ea99, 32'h40c6a394} /* (23, 11, 16) {real, imag} */,
  {32'h4080b41f, 32'h3f62e089} /* (23, 11, 15) {real, imag} */,
  {32'h40a5ba5d, 32'hc085bbf0} /* (23, 11, 14) {real, imag} */,
  {32'h40f09e9e, 32'hc11f0dd0} /* (23, 11, 13) {real, imag} */,
  {32'h40ab87ee, 32'hc0670721} /* (23, 11, 12) {real, imag} */,
  {32'h40887889, 32'h4068b4ae} /* (23, 11, 11) {real, imag} */,
  {32'hbe418f30, 32'h3fcdd8bc} /* (23, 11, 10) {real, imag} */,
  {32'hbf12fc0c, 32'hc095e36e} /* (23, 11, 9) {real, imag} */,
  {32'hc0a3865d, 32'hc05e7f8e} /* (23, 11, 8) {real, imag} */,
  {32'hc0a0a856, 32'hbfa109b0} /* (23, 11, 7) {real, imag} */,
  {32'h4009afaf, 32'hbfba2e0a} /* (23, 11, 6) {real, imag} */,
  {32'h40a15591, 32'h403edf86} /* (23, 11, 5) {real, imag} */,
  {32'hbfb7d88b, 32'hc06cbaf0} /* (23, 11, 4) {real, imag} */,
  {32'hc054def1, 32'hc10057b5} /* (23, 11, 3) {real, imag} */,
  {32'h3e94c798, 32'hbf07f218} /* (23, 11, 2) {real, imag} */,
  {32'h40298144, 32'h40460f56} /* (23, 11, 1) {real, imag} */,
  {32'h403183b4, 32'hbf6ff310} /* (23, 11, 0) {real, imag} */,
  {32'hbf400f02, 32'h401a1d57} /* (23, 10, 31) {real, imag} */,
  {32'hc02c617e, 32'h40bc0d22} /* (23, 10, 30) {real, imag} */,
  {32'hbff6757c, 32'h40ac2765} /* (23, 10, 29) {real, imag} */,
  {32'hc035a72f, 32'hbe9f92a8} /* (23, 10, 28) {real, imag} */,
  {32'h3f6f7ef6, 32'h3fecdd4c} /* (23, 10, 27) {real, imag} */,
  {32'h40d736f8, 32'hbfe93e80} /* (23, 10, 26) {real, imag} */,
  {32'h4086bf58, 32'hbec2d82c} /* (23, 10, 25) {real, imag} */,
  {32'hbfce0fff, 32'hc0938695} /* (23, 10, 24) {real, imag} */,
  {32'hc114c7e0, 32'h3ded7068} /* (23, 10, 23) {real, imag} */,
  {32'hc11e5818, 32'h40a87a86} /* (23, 10, 22) {real, imag} */,
  {32'hbfded450, 32'hc01ec1c4} /* (23, 10, 21) {real, imag} */,
  {32'hbfdf5726, 32'hbf1a8cc0} /* (23, 10, 20) {real, imag} */,
  {32'hc05584f9, 32'h4042e2ce} /* (23, 10, 19) {real, imag} */,
  {32'hc02536b6, 32'h40525d23} /* (23, 10, 18) {real, imag} */,
  {32'h3fb5c2da, 32'h410e29e5} /* (23, 10, 17) {real, imag} */,
  {32'h403dcbd5, 32'h40a62086} /* (23, 10, 16) {real, imag} */,
  {32'hbf8d05a6, 32'hbf043390} /* (23, 10, 15) {real, imag} */,
  {32'h3fe750b0, 32'hbfae3b3e} /* (23, 10, 14) {real, imag} */,
  {32'h3fc540b1, 32'h3fc0d200} /* (23, 10, 13) {real, imag} */,
  {32'hbebc3e50, 32'hc04ec0a0} /* (23, 10, 12) {real, imag} */,
  {32'h41226df0, 32'hc08f91bc} /* (23, 10, 11) {real, imag} */,
  {32'h4165cf80, 32'hc08fd9d3} /* (23, 10, 10) {real, imag} */,
  {32'h409e0720, 32'hc01cfec8} /* (23, 10, 9) {real, imag} */,
  {32'hbd106240, 32'h4013b676} /* (23, 10, 8) {real, imag} */,
  {32'hc03bc450, 32'h3e5b4ad0} /* (23, 10, 7) {real, imag} */,
  {32'h3fa42b25, 32'hc0f545ec} /* (23, 10, 6) {real, imag} */,
  {32'hbfa1c2cf, 32'hc0c1d4c6} /* (23, 10, 5) {real, imag} */,
  {32'hc09dbe72, 32'hc0c1af38} /* (23, 10, 4) {real, imag} */,
  {32'h40773d8a, 32'h4046c71c} /* (23, 10, 3) {real, imag} */,
  {32'h40706ab2, 32'h3eb4ce10} /* (23, 10, 2) {real, imag} */,
  {32'h4000b2a4, 32'hc0a2d964} /* (23, 10, 1) {real, imag} */,
  {32'h40260a28, 32'hbe6df0d4} /* (23, 10, 0) {real, imag} */,
  {32'h405fbe96, 32'h408c3070} /* (23, 9, 31) {real, imag} */,
  {32'h3fa876e5, 32'h40ad4432} /* (23, 9, 30) {real, imag} */,
  {32'hbdf7c6d8, 32'h3fb77d3a} /* (23, 9, 29) {real, imag} */,
  {32'h40f116b0, 32'h3ff42232} /* (23, 9, 28) {real, imag} */,
  {32'h4045c8c5, 32'h4081b61c} /* (23, 9, 27) {real, imag} */,
  {32'hbf94263a, 32'h3d015460} /* (23, 9, 26) {real, imag} */,
  {32'h4055ae68, 32'hc056a911} /* (23, 9, 25) {real, imag} */,
  {32'h4110bd4f, 32'h404153f0} /* (23, 9, 24) {real, imag} */,
  {32'h40bcda42, 32'h3f159d40} /* (23, 9, 23) {real, imag} */,
  {32'h40a62e40, 32'h400c94ea} /* (23, 9, 22) {real, imag} */,
  {32'h40e99010, 32'hc011b202} /* (23, 9, 21) {real, imag} */,
  {32'h40f4fab6, 32'h406e44e3} /* (23, 9, 20) {real, imag} */,
  {32'h403d1fd9, 32'h4134ba8e} /* (23, 9, 19) {real, imag} */,
  {32'hbfb075cd, 32'h3f89a860} /* (23, 9, 18) {real, imag} */,
  {32'h3fab662c, 32'hc01b2175} /* (23, 9, 17) {real, imag} */,
  {32'h40e3ee6c, 32'hc0b09e18} /* (23, 9, 16) {real, imag} */,
  {32'h4087f243, 32'hc0ed5a72} /* (23, 9, 15) {real, imag} */,
  {32'hc0d4d4d0, 32'hc0bcb0e3} /* (23, 9, 14) {real, imag} */,
  {32'hbdc57370, 32'hc0ac960f} /* (23, 9, 13) {real, imag} */,
  {32'h402ed3df, 32'h3ee88d28} /* (23, 9, 12) {real, imag} */,
  {32'hbfed2816, 32'h4091b429} /* (23, 9, 11) {real, imag} */,
  {32'hc0d71545, 32'hc098b216} /* (23, 9, 10) {real, imag} */,
  {32'hc11810d4, 32'hc0b737cb} /* (23, 9, 9) {real, imag} */,
  {32'hc083f3e7, 32'hc0a62cf6} /* (23, 9, 8) {real, imag} */,
  {32'hc0b0f7da, 32'hc07433c2} /* (23, 9, 7) {real, imag} */,
  {32'hbfc39c53, 32'hc108b740} /* (23, 9, 6) {real, imag} */,
  {32'h3fbbc21c, 32'hc066f977} /* (23, 9, 5) {real, imag} */,
  {32'hc0ab153c, 32'h40cd7fda} /* (23, 9, 4) {real, imag} */,
  {32'hc122a92a, 32'h410d0572} /* (23, 9, 3) {real, imag} */,
  {32'hc07fda9c, 32'h4004eae6} /* (23, 9, 2) {real, imag} */,
  {32'hbf534714, 32'hc0a1b97c} /* (23, 9, 1) {real, imag} */,
  {32'hbfad2d4c, 32'hc03eace6} /* (23, 9, 0) {real, imag} */,
  {32'h3fbc8e92, 32'h401f5b68} /* (23, 8, 31) {real, imag} */,
  {32'h40309bbe, 32'h402dcc5c} /* (23, 8, 30) {real, imag} */,
  {32'hc06d9f4d, 32'h40a09c50} /* (23, 8, 29) {real, imag} */,
  {32'hc0e37a19, 32'h3e9140a0} /* (23, 8, 28) {real, imag} */,
  {32'hc0150959, 32'hc04aef81} /* (23, 8, 27) {real, imag} */,
  {32'hc0691306, 32'h40d6468f} /* (23, 8, 26) {real, imag} */,
  {32'h4114c3ce, 32'h409a7d16} /* (23, 8, 25) {real, imag} */,
  {32'h40f13a31, 32'h3f69fad6} /* (23, 8, 24) {real, imag} */,
  {32'hc093836e, 32'h404a1c2e} /* (23, 8, 23) {real, imag} */,
  {32'hc10b6c07, 32'h40c13c73} /* (23, 8, 22) {real, imag} */,
  {32'hc1645050, 32'h4184ee48} /* (23, 8, 21) {real, imag} */,
  {32'hc091c182, 32'h4095b01b} /* (23, 8, 20) {real, imag} */,
  {32'h401feac0, 32'hbff3e8aa} /* (23, 8, 19) {real, imag} */,
  {32'h3bdf3180, 32'hc0b65d74} /* (23, 8, 18) {real, imag} */,
  {32'hbf698484, 32'h3d6a5d80} /* (23, 8, 17) {real, imag} */,
  {32'h3f1756d0, 32'h3f7c65ae} /* (23, 8, 16) {real, imag} */,
  {32'hc09dbea0, 32'h3f959f16} /* (23, 8, 15) {real, imag} */,
  {32'hc0983992, 32'h40330df4} /* (23, 8, 14) {real, imag} */,
  {32'hc097ac61, 32'h410270f9} /* (23, 8, 13) {real, imag} */,
  {32'h404e2a36, 32'h40a248b1} /* (23, 8, 12) {real, imag} */,
  {32'h409ab6a3, 32'h402f8143} /* (23, 8, 11) {real, imag} */,
  {32'h40187930, 32'h3f5b5868} /* (23, 8, 10) {real, imag} */,
  {32'h40c769f8, 32'h410a61a1} /* (23, 8, 9) {real, imag} */,
  {32'hc08d76a6, 32'h3f648c50} /* (23, 8, 8) {real, imag} */,
  {32'h40c3f133, 32'h40106eb2} /* (23, 8, 7) {real, imag} */,
  {32'h40a807ad, 32'h411fb0b7} /* (23, 8, 6) {real, imag} */,
  {32'hbf0d3260, 32'h3f9ca1d4} /* (23, 8, 5) {real, imag} */,
  {32'h3f97b650, 32'hc0a0bbdb} /* (23, 8, 4) {real, imag} */,
  {32'h40882945, 32'hbfc2b33a} /* (23, 8, 3) {real, imag} */,
  {32'hc0a6fac2, 32'hc0802100} /* (23, 8, 2) {real, imag} */,
  {32'hc0ef61fa, 32'hc088db6d} /* (23, 8, 1) {real, imag} */,
  {32'h3fb24a78, 32'hc004f30e} /* (23, 8, 0) {real, imag} */,
  {32'h406b4321, 32'h40dfb3c0} /* (23, 7, 31) {real, imag} */,
  {32'h4020e20e, 32'h4130c323} /* (23, 7, 30) {real, imag} */,
  {32'hc0a0c1f5, 32'hbfec2fa4} /* (23, 7, 29) {real, imag} */,
  {32'h41358e7e, 32'hc128e16f} /* (23, 7, 28) {real, imag} */,
  {32'h4156544e, 32'hc0a3aee5} /* (23, 7, 27) {real, imag} */,
  {32'h40b44d32, 32'hc061197c} /* (23, 7, 26) {real, imag} */,
  {32'h409325b3, 32'hc084709b} /* (23, 7, 25) {real, imag} */,
  {32'h4120039f, 32'h402b9210} /* (23, 7, 24) {real, imag} */,
  {32'h408cb8e2, 32'hc09b461e} /* (23, 7, 23) {real, imag} */,
  {32'hc0220eb3, 32'hc08eef0f} /* (23, 7, 22) {real, imag} */,
  {32'h3fb394fa, 32'hc045a7ce} /* (23, 7, 21) {real, imag} */,
  {32'h40e33d79, 32'h40b6de8e} /* (23, 7, 20) {real, imag} */,
  {32'h408bb5b7, 32'h408b4f01} /* (23, 7, 19) {real, imag} */,
  {32'hc0cbcfd6, 32'h413c133f} /* (23, 7, 18) {real, imag} */,
  {32'hc0e55020, 32'h41354323} /* (23, 7, 17) {real, imag} */,
  {32'hc04aeb64, 32'h3f80ac9b} /* (23, 7, 16) {real, imag} */,
  {32'hc0151cc6, 32'h3dee6800} /* (23, 7, 15) {real, imag} */,
  {32'h40c00cdf, 32'h408be995} /* (23, 7, 14) {real, imag} */,
  {32'h401f637e, 32'h3fda9498} /* (23, 7, 13) {real, imag} */,
  {32'hc032ae54, 32'h413122f6} /* (23, 7, 12) {real, imag} */,
  {32'hc115c542, 32'h40b7f0f7} /* (23, 7, 11) {real, imag} */,
  {32'hc15a6cb4, 32'hc05641c6} /* (23, 7, 10) {real, imag} */,
  {32'hbfdfbff6, 32'hc08a851e} /* (23, 7, 9) {real, imag} */,
  {32'h4117709e, 32'hc03d2021} /* (23, 7, 8) {real, imag} */,
  {32'h3fead27a, 32'hbff09f37} /* (23, 7, 7) {real, imag} */,
  {32'hc17bab98, 32'hc04ab4f7} /* (23, 7, 6) {real, imag} */,
  {32'hc1575903, 32'h40320e53} /* (23, 7, 5) {real, imag} */,
  {32'hc10466a3, 32'hc0c159a6} /* (23, 7, 4) {real, imag} */,
  {32'hbf62f1d4, 32'hc0609b58} /* (23, 7, 3) {real, imag} */,
  {32'h4174de00, 32'hbf6a2e20} /* (23, 7, 2) {real, imag} */,
  {32'h412cdec0, 32'hc067d921} /* (23, 7, 1) {real, imag} */,
  {32'h3fbd69f4, 32'h3fb22fe2} /* (23, 7, 0) {real, imag} */,
  {32'h40932e53, 32'hc099376c} /* (23, 6, 31) {real, imag} */,
  {32'h411e848e, 32'hbf8e3060} /* (23, 6, 30) {real, imag} */,
  {32'h414c9e06, 32'h40a879f2} /* (23, 6, 29) {real, imag} */,
  {32'h3f04a478, 32'hbf886dc2} /* (23, 6, 28) {real, imag} */,
  {32'hc0baa56a, 32'hbfd21edb} /* (23, 6, 27) {real, imag} */,
  {32'hbebec180, 32'hbfcbc5aa} /* (23, 6, 26) {real, imag} */,
  {32'hc093604a, 32'h4064917c} /* (23, 6, 25) {real, imag} */,
  {32'h3f7c2522, 32'h3f298ba8} /* (23, 6, 24) {real, imag} */,
  {32'hc0176371, 32'h41647b22} /* (23, 6, 23) {real, imag} */,
  {32'h3efe666c, 32'h415bed8f} /* (23, 6, 22) {real, imag} */,
  {32'h40c6bad8, 32'h410fb92a} /* (23, 6, 21) {real, imag} */,
  {32'hc0aea31a, 32'h410078d1} /* (23, 6, 20) {real, imag} */,
  {32'hc102f3b4, 32'h40d46c9c} /* (23, 6, 19) {real, imag} */,
  {32'h40af1b8c, 32'hc1188785} /* (23, 6, 18) {real, imag} */,
  {32'h40f6dd02, 32'hc13550f0} /* (23, 6, 17) {real, imag} */,
  {32'hc02b22c6, 32'h3fe97b8a} /* (23, 6, 16) {real, imag} */,
  {32'h408fa71d, 32'hc138d3ed} /* (23, 6, 15) {real, imag} */,
  {32'hc00896cc, 32'hc103c629} /* (23, 6, 14) {real, imag} */,
  {32'hc10249cc, 32'h40f0ed28} /* (23, 6, 13) {real, imag} */,
  {32'hc199a300, 32'h400d6b6a} /* (23, 6, 12) {real, imag} */,
  {32'hc128242a, 32'hc05ce140} /* (23, 6, 11) {real, imag} */,
  {32'hbfd499ec, 32'h3ff122d5} /* (23, 6, 10) {real, imag} */,
  {32'h40b8d7a3, 32'hc151f22c} /* (23, 6, 9) {real, imag} */,
  {32'h40d7a044, 32'hc1129bc8} /* (23, 6, 8) {real, imag} */,
  {32'hbfcae9b8, 32'hc0c073e0} /* (23, 6, 7) {real, imag} */,
  {32'hc1456a62, 32'hc122310c} /* (23, 6, 6) {real, imag} */,
  {32'hc0ab21aa, 32'hc12ea869} /* (23, 6, 5) {real, imag} */,
  {32'hbd98a900, 32'h40970fd8} /* (23, 6, 4) {real, imag} */,
  {32'hc13a0e6a, 32'h405e5fca} /* (23, 6, 3) {real, imag} */,
  {32'hc1403242, 32'h417a262c} /* (23, 6, 2) {real, imag} */,
  {32'hc0a6c12d, 32'h410b9976} /* (23, 6, 1) {real, imag} */,
  {32'hc03799b8, 32'h40c39e08} /* (23, 6, 0) {real, imag} */,
  {32'h40e0a5da, 32'h4020341a} /* (23, 5, 31) {real, imag} */,
  {32'h4104dd45, 32'h3fb7e72f} /* (23, 5, 30) {real, imag} */,
  {32'h3e2277d8, 32'hc0f223ac} /* (23, 5, 29) {real, imag} */,
  {32'h3ff28fbf, 32'h4012dabc} /* (23, 5, 28) {real, imag} */,
  {32'h40feb2f3, 32'h40e78793} /* (23, 5, 27) {real, imag} */,
  {32'h4014d37c, 32'hbeaf69f0} /* (23, 5, 26) {real, imag} */,
  {32'hc086ac1e, 32'hc006c66a} /* (23, 5, 25) {real, imag} */,
  {32'h3ff4b338, 32'h413e0f8c} /* (23, 5, 24) {real, imag} */,
  {32'h4159b3f0, 32'h415a8be4} /* (23, 5, 23) {real, imag} */,
  {32'hbff525d8, 32'hc143bcd4} /* (23, 5, 22) {real, imag} */,
  {32'hc0d866a1, 32'hc1892c8c} /* (23, 5, 21) {real, imag} */,
  {32'h3f7f0f72, 32'hc189ca3a} /* (23, 5, 20) {real, imag} */,
  {32'h410d11bf, 32'hc1234d54} /* (23, 5, 19) {real, imag} */,
  {32'h40ad42b8, 32'hc14abeca} /* (23, 5, 18) {real, imag} */,
  {32'h406f83d0, 32'hc190edf3} /* (23, 5, 17) {real, imag} */,
  {32'hc0d67df2, 32'hc0e5a782} /* (23, 5, 16) {real, imag} */,
  {32'hc099c86d, 32'hbfa29858} /* (23, 5, 15) {real, imag} */,
  {32'hbf8b2f70, 32'hbf814338} /* (23, 5, 14) {real, imag} */,
  {32'h405955b6, 32'h411021ef} /* (23, 5, 13) {real, imag} */,
  {32'hc0627ccc, 32'hbf85fbe8} /* (23, 5, 12) {real, imag} */,
  {32'hc0aa5363, 32'hc10269b2} /* (23, 5, 11) {real, imag} */,
  {32'hbf9c4ce5, 32'h40a86098} /* (23, 5, 10) {real, imag} */,
  {32'hc0b08f5c, 32'h41489337} /* (23, 5, 9) {real, imag} */,
  {32'h40a91d93, 32'h403dbdda} /* (23, 5, 8) {real, imag} */,
  {32'h4118715c, 32'h3fe97fe0} /* (23, 5, 7) {real, imag} */,
  {32'hc0d6bb86, 32'hc0bf3aba} /* (23, 5, 6) {real, imag} */,
  {32'hc10c7ac0, 32'h3f05c8c8} /* (23, 5, 5) {real, imag} */,
  {32'h41371f1d, 32'hbd7b0910} /* (23, 5, 4) {real, imag} */,
  {32'h4024c67c, 32'h4127e8f2} /* (23, 5, 3) {real, imag} */,
  {32'hc16eddae, 32'h415a4886} /* (23, 5, 2) {real, imag} */,
  {32'hbf9230df, 32'hc08a3e79} /* (23, 5, 1) {real, imag} */,
  {32'h4035caec, 32'hc0bd98c0} /* (23, 5, 0) {real, imag} */,
  {32'h40216df8, 32'hc12b002d} /* (23, 4, 31) {real, imag} */,
  {32'h40868b28, 32'hc1372d96} /* (23, 4, 30) {real, imag} */,
  {32'hc0ab5371, 32'h3fdab488} /* (23, 4, 29) {real, imag} */,
  {32'hc0323c8a, 32'h404a45d8} /* (23, 4, 28) {real, imag} */,
  {32'h40be2e15, 32'h41402fad} /* (23, 4, 27) {real, imag} */,
  {32'h41845b3d, 32'h415ced7a} /* (23, 4, 26) {real, imag} */,
  {32'h41340e47, 32'h410bdaf3} /* (23, 4, 25) {real, imag} */,
  {32'h3ffed8ba, 32'hc02e1792} /* (23, 4, 24) {real, imag} */,
  {32'h408cbe06, 32'hc0f05960} /* (23, 4, 23) {real, imag} */,
  {32'h411882b6, 32'hbf503e50} /* (23, 4, 22) {real, imag} */,
  {32'h40b902de, 32'h3f7d4bb0} /* (23, 4, 21) {real, imag} */,
  {32'h40e52bd2, 32'h40a0651e} /* (23, 4, 20) {real, imag} */,
  {32'h3f8728e0, 32'h408329a0} /* (23, 4, 19) {real, imag} */,
  {32'hbfa2f462, 32'h3fcab4f0} /* (23, 4, 18) {real, imag} */,
  {32'hc0868c68, 32'h41930bd1} /* (23, 4, 17) {real, imag} */,
  {32'h405954fb, 32'h40cfd778} /* (23, 4, 16) {real, imag} */,
  {32'hc0b891f6, 32'h404ee788} /* (23, 4, 15) {real, imag} */,
  {32'hc0135ad0, 32'h40398721} /* (23, 4, 14) {real, imag} */,
  {32'hc1267452, 32'h417f2f35} /* (23, 4, 13) {real, imag} */,
  {32'hc19bb45f, 32'h40af4de1} /* (23, 4, 12) {real, imag} */,
  {32'hc039935c, 32'hc10df2d4} /* (23, 4, 11) {real, imag} */,
  {32'hc06ff89e, 32'hc105c8b2} /* (23, 4, 10) {real, imag} */,
  {32'hc0b57a8e, 32'h40c0ea23} /* (23, 4, 9) {real, imag} */,
  {32'hbfcf5fc4, 32'h40b683fc} /* (23, 4, 8) {real, imag} */,
  {32'hc063bf68, 32'hc0e0636d} /* (23, 4, 7) {real, imag} */,
  {32'h410cf2f9, 32'h4040b07e} /* (23, 4, 6) {real, imag} */,
  {32'h4119e027, 32'h40dfcda3} /* (23, 4, 5) {real, imag} */,
  {32'h40b62e1a, 32'h4116fa92} /* (23, 4, 4) {real, imag} */,
  {32'h3fb254a0, 32'hc0fc7d1e} /* (23, 4, 3) {real, imag} */,
  {32'hc0b079a2, 32'hc02d0065} /* (23, 4, 2) {real, imag} */,
  {32'hbee25a40, 32'h41ae053f} /* (23, 4, 1) {real, imag} */,
  {32'h400b886e, 32'h40c49bf4} /* (23, 4, 0) {real, imag} */,
  {32'hc127d49e, 32'hc0008f14} /* (23, 3, 31) {real, imag} */,
  {32'hc17befad, 32'h3f5af866} /* (23, 3, 30) {real, imag} */,
  {32'hc0274394, 32'h4117d82f} /* (23, 3, 29) {real, imag} */,
  {32'hc0a81daa, 32'h3ea680b8} /* (23, 3, 28) {real, imag} */,
  {32'hc10923c8, 32'hc0ab8c3d} /* (23, 3, 27) {real, imag} */,
  {32'h404f08c1, 32'hc0124a56} /* (23, 3, 26) {real, imag} */,
  {32'h41072a82, 32'hc0f9c2f3} /* (23, 3, 25) {real, imag} */,
  {32'hbbfdf000, 32'h3db1d180} /* (23, 3, 24) {real, imag} */,
  {32'hc0ef403d, 32'hc1274ad8} /* (23, 3, 23) {real, imag} */,
  {32'h3f66ca50, 32'hc11a17b8} /* (23, 3, 22) {real, imag} */,
  {32'h3e195400, 32'hc13265b2} /* (23, 3, 21) {real, imag} */,
  {32'hc08c08f5, 32'hc12383be} /* (23, 3, 20) {real, imag} */,
  {32'hbf2ad684, 32'h40b18da7} /* (23, 3, 19) {real, imag} */,
  {32'hc127e098, 32'h3fee7ebd} /* (23, 3, 18) {real, imag} */,
  {32'hc1a24ef3, 32'hbfc46584} /* (23, 3, 17) {real, imag} */,
  {32'hc11ed7f2, 32'h4151ae57} /* (23, 3, 16) {real, imag} */,
  {32'hc15c6312, 32'h41042e15} /* (23, 3, 15) {real, imag} */,
  {32'hc08fa0c0, 32'hc008ce98} /* (23, 3, 14) {real, imag} */,
  {32'h41551d02, 32'hbf8ed894} /* (23, 3, 13) {real, imag} */,
  {32'h41929498, 32'hc0d58a8c} /* (23, 3, 12) {real, imag} */,
  {32'h40c5ee0c, 32'hbda11c80} /* (23, 3, 11) {real, imag} */,
  {32'h4144c6ee, 32'hc07e55d8} /* (23, 3, 10) {real, imag} */,
  {32'h419d55f4, 32'hc165e296} /* (23, 3, 9) {real, imag} */,
  {32'h40f8dae1, 32'hc1432487} /* (23, 3, 8) {real, imag} */,
  {32'h4169e898, 32'hc1689130} /* (23, 3, 7) {real, imag} */,
  {32'h40c94f9a, 32'hc160e9c2} /* (23, 3, 6) {real, imag} */,
  {32'h41195644, 32'h3d421900} /* (23, 3, 5) {real, imag} */,
  {32'h40bcacb3, 32'h40c466e4} /* (23, 3, 4) {real, imag} */,
  {32'hc08db558, 32'h4155648a} /* (23, 3, 3) {real, imag} */,
  {32'hc0de423d, 32'h414e57a0} /* (23, 3, 2) {real, imag} */,
  {32'hbeec1180, 32'hc05ac9fc} /* (23, 3, 1) {real, imag} */,
  {32'hc0490ea9, 32'hc0c05fbf} /* (23, 3, 0) {real, imag} */,
  {32'hc07cb027, 32'hc0ae2b15} /* (23, 2, 31) {real, imag} */,
  {32'h4109af42, 32'hc1053e11} /* (23, 2, 30) {real, imag} */,
  {32'h418dc360, 32'hc135aa87} /* (23, 2, 29) {real, imag} */,
  {32'h404d8758, 32'h3f41da6b} /* (23, 2, 28) {real, imag} */,
  {32'hc125b05b, 32'h3eac20e0} /* (23, 2, 27) {real, imag} */,
  {32'hbf88fe88, 32'hbf6589d0} /* (23, 2, 26) {real, imag} */,
  {32'h4010d3f3, 32'h4171af80} /* (23, 2, 25) {real, imag} */,
  {32'h40b1a65c, 32'h417c9fc3} /* (23, 2, 24) {real, imag} */,
  {32'hc0da6856, 32'h418e5593} /* (23, 2, 23) {real, imag} */,
  {32'hc14f3279, 32'h41ae24e3} /* (23, 2, 22) {real, imag} */,
  {32'hc0f0fc04, 32'h3e971a10} /* (23, 2, 21) {real, imag} */,
  {32'hc0672a26, 32'hc0edaa00} /* (23, 2, 20) {real, imag} */,
  {32'hc065b15e, 32'h400801d4} /* (23, 2, 19) {real, imag} */,
  {32'hc0c5dd04, 32'hc0c9a0cd} /* (23, 2, 18) {real, imag} */,
  {32'hbfe86476, 32'hc1652fc0} /* (23, 2, 17) {real, imag} */,
  {32'hc1927446, 32'hc141e396} /* (23, 2, 16) {real, imag} */,
  {32'hc1799aba, 32'hc0b4d511} /* (23, 2, 15) {real, imag} */,
  {32'hbfce2726, 32'h40c2c74c} /* (23, 2, 14) {real, imag} */,
  {32'hc0bd27ca, 32'h4160eae0} /* (23, 2, 13) {real, imag} */,
  {32'hc1a9a688, 32'h410b1d2a} /* (23, 2, 12) {real, imag} */,
  {32'hc15cc4d8, 32'hc110f6e9} /* (23, 2, 11) {real, imag} */,
  {32'h409ce08c, 32'hbed4bf6a} /* (23, 2, 10) {real, imag} */,
  {32'h417ddb31, 32'h40fe8a51} /* (23, 2, 9) {real, imag} */,
  {32'h416d3cc2, 32'hc037d848} /* (23, 2, 8) {real, imag} */,
  {32'h416ba212, 32'h415d39fa} /* (23, 2, 7) {real, imag} */,
  {32'h4111a860, 32'h41584e8b} /* (23, 2, 6) {real, imag} */,
  {32'h41a77a06, 32'h416ed6b6} /* (23, 2, 5) {real, imag} */,
  {32'h41756e41, 32'h40149268} /* (23, 2, 4) {real, imag} */,
  {32'h3d827cf8, 32'hc185b188} /* (23, 2, 3) {real, imag} */,
  {32'hc0648104, 32'h40ac66e4} /* (23, 2, 2) {real, imag} */,
  {32'h403cd3cc, 32'h40e8062a} /* (23, 2, 1) {real, imag} */,
  {32'hbf8762ff, 32'hc00e8ce8} /* (23, 2, 0) {real, imag} */,
  {32'hc13b1cb6, 32'hc12f5225} /* (23, 1, 31) {real, imag} */,
  {32'hc113b850, 32'hc1400f94} /* (23, 1, 30) {real, imag} */,
  {32'hc097d0b8, 32'hc089e24d} /* (23, 1, 29) {real, imag} */,
  {32'hc0b816fa, 32'hc0136bf4} /* (23, 1, 28) {real, imag} */,
  {32'hc0124a5e, 32'hbe59a7c0} /* (23, 1, 27) {real, imag} */,
  {32'h413852bd, 32'hc15f3c11} /* (23, 1, 26) {real, imag} */,
  {32'hc18c589b, 32'hc0eda7b8} /* (23, 1, 25) {real, imag} */,
  {32'hc184bf50, 32'hc120aa9a} /* (23, 1, 24) {real, imag} */,
  {32'hc068232b, 32'hc147c085} /* (23, 1, 23) {real, imag} */,
  {32'hc09a069b, 32'hc18d6893} /* (23, 1, 22) {real, imag} */,
  {32'hc115992a, 32'h405a4acc} /* (23, 1, 21) {real, imag} */,
  {32'hc07e04e9, 32'h416603ea} /* (23, 1, 20) {real, imag} */,
  {32'h3f65a370, 32'h41238449} /* (23, 1, 19) {real, imag} */,
  {32'h40da693e, 32'h40e68004} /* (23, 1, 18) {real, imag} */,
  {32'hc107cfe0, 32'h40f262be} /* (23, 1, 17) {real, imag} */,
  {32'hc14049da, 32'h410d630c} /* (23, 1, 16) {real, imag} */,
  {32'hbc1ae600, 32'h40ed6e38} /* (23, 1, 15) {real, imag} */,
  {32'h40f5f39b, 32'hc00468a4} /* (23, 1, 14) {real, imag} */,
  {32'h40e8ab02, 32'h40b0c7b6} /* (23, 1, 13) {real, imag} */,
  {32'h40ac807c, 32'h3fe62c20} /* (23, 1, 12) {real, imag} */,
  {32'h4131f815, 32'h3fd23648} /* (23, 1, 11) {real, imag} */,
  {32'hbfaef480, 32'hc1169489} /* (23, 1, 10) {real, imag} */,
  {32'h3f1bf010, 32'hc06e9b0e} /* (23, 1, 9) {real, imag} */,
  {32'h412f5dc6, 32'hc0244400} /* (23, 1, 8) {real, imag} */,
  {32'hc0f80843, 32'hc12cde52} /* (23, 1, 7) {real, imag} */,
  {32'hc0f7480a, 32'hc1257578} /* (23, 1, 6) {real, imag} */,
  {32'hc1214b96, 32'hc0bb3776} /* (23, 1, 5) {real, imag} */,
  {32'hc149fa6b, 32'hc0e23d41} /* (23, 1, 4) {real, imag} */,
  {32'hc149f43e, 32'hc1545a7f} /* (23, 1, 3) {real, imag} */,
  {32'hc1515fb7, 32'hc1367886} /* (23, 1, 2) {real, imag} */,
  {32'hc14c30e3, 32'hc1b747a4} /* (23, 1, 1) {real, imag} */,
  {32'hc0616ee2, 32'hc13c0b17} /* (23, 1, 0) {real, imag} */,
  {32'h3f9ecd4e, 32'hc0dc2f03} /* (23, 0, 31) {real, imag} */,
  {32'hc15aed32, 32'hbfba3aca} /* (23, 0, 30) {real, imag} */,
  {32'hc167dda5, 32'hc1121fc6} /* (23, 0, 29) {real, imag} */,
  {32'hc101bb94, 32'hc12c76f5} /* (23, 0, 28) {real, imag} */,
  {32'hc0997786, 32'hc070f747} /* (23, 0, 27) {real, imag} */,
  {32'hc15d2f4a, 32'hc07a918a} /* (23, 0, 26) {real, imag} */,
  {32'hc13808cc, 32'hc182e540} /* (23, 0, 25) {real, imag} */,
  {32'hbf77322e, 32'hc1a7d3b6} /* (23, 0, 24) {real, imag} */,
  {32'hc000e8ec, 32'hc17fc7c2} /* (23, 0, 23) {real, imag} */,
  {32'h3ffcdbb6, 32'hc197d01b} /* (23, 0, 22) {real, imag} */,
  {32'hc0d0edee, 32'hc1085f3d} /* (23, 0, 21) {real, imag} */,
  {32'h3eb9fcce, 32'h41707be2} /* (23, 0, 20) {real, imag} */,
  {32'h41193eb6, 32'h40afd1e3} /* (23, 0, 19) {real, imag} */,
  {32'h40a2d21c, 32'h4109f2aa} /* (23, 0, 18) {real, imag} */,
  {32'hc13f60e2, 32'hbfbf3f64} /* (23, 0, 17) {real, imag} */,
  {32'hbfb897e0, 32'hc10c1f7a} /* (23, 0, 16) {real, imag} */,
  {32'h40eda110, 32'hc09bb642} /* (23, 0, 15) {real, imag} */,
  {32'h40d6a2c0, 32'hc13abb68} /* (23, 0, 14) {real, imag} */,
  {32'h4171c1dc, 32'hc1ae20df} /* (23, 0, 13) {real, imag} */,
  {32'h417ff84d, 32'hc184171c} /* (23, 0, 12) {real, imag} */,
  {32'h412f84b7, 32'h41260c10} /* (23, 0, 11) {real, imag} */,
  {32'h4025f914, 32'h40e7a574} /* (23, 0, 10) {real, imag} */,
  {32'hc0896b38, 32'hc1664119} /* (23, 0, 9) {real, imag} */,
  {32'h40323404, 32'hc01969cc} /* (23, 0, 8) {real, imag} */,
  {32'h41ac2df0, 32'h40983320} /* (23, 0, 7) {real, imag} */,
  {32'h40df1228, 32'h3fd3dd9b} /* (23, 0, 6) {real, imag} */,
  {32'hc18378ef, 32'hc156721d} /* (23, 0, 5) {real, imag} */,
  {32'hc0e3db82, 32'hc082c63c} /* (23, 0, 4) {real, imag} */,
  {32'h40a4d5f6, 32'hc0492d66} /* (23, 0, 3) {real, imag} */,
  {32'hbf85290d, 32'hc11f7a11} /* (23, 0, 2) {real, imag} */,
  {32'hc1525ff0, 32'hc1107a3a} /* (23, 0, 1) {real, imag} */,
  {32'hc036bd5f, 32'hc0e1cf4a} /* (23, 0, 0) {real, imag} */,
  {32'hc02cb100, 32'hc0cb1f0e} /* (22, 31, 31) {real, imag} */,
  {32'hc1871877, 32'hbfbea500} /* (22, 31, 30) {real, imag} */,
  {32'hc1553fac, 32'hc011f874} /* (22, 31, 29) {real, imag} */,
  {32'hc178e956, 32'h40bac324} /* (22, 31, 28) {real, imag} */,
  {32'hc0abbea6, 32'h400fff5d} /* (22, 31, 27) {real, imag} */,
  {32'hc109a62b, 32'hc13ed9b5} /* (22, 31, 26) {real, imag} */,
  {32'hc18edbe5, 32'hc0b263b5} /* (22, 31, 25) {real, imag} */,
  {32'hc1aed479, 32'hc0ffb03a} /* (22, 31, 24) {real, imag} */,
  {32'hc138571e, 32'hc12de024} /* (22, 31, 23) {real, imag} */,
  {32'hbf75267f, 32'hc0ec14eb} /* (22, 31, 22) {real, imag} */,
  {32'h402df548, 32'h3ef05f28} /* (22, 31, 21) {real, imag} */,
  {32'h414af31e, 32'h405e1c99} /* (22, 31, 20) {real, imag} */,
  {32'h41082f64, 32'h4115a2e4} /* (22, 31, 19) {real, imag} */,
  {32'h419fe08a, 32'h3fc872e8} /* (22, 31, 18) {real, imag} */,
  {32'h418cac86, 32'hbea264c2} /* (22, 31, 17) {real, imag} */,
  {32'hbeb0e876, 32'hc141813e} /* (22, 31, 16) {real, imag} */,
  {32'hbf2507f2, 32'hc0abdf31} /* (22, 31, 15) {real, imag} */,
  {32'h4036a13c, 32'hbfc3fda4} /* (22, 31, 14) {real, imag} */,
  {32'hbe1eff00, 32'h415f204e} /* (22, 31, 13) {real, imag} */,
  {32'h40bff168, 32'h40a7656c} /* (22, 31, 12) {real, imag} */,
  {32'h41931991, 32'hc10a0e73} /* (22, 31, 11) {real, imag} */,
  {32'h3f330228, 32'hc12531da} /* (22, 31, 10) {real, imag} */,
  {32'h3eb09148, 32'hc00d635c} /* (22, 31, 9) {real, imag} */,
  {32'hc024ff82, 32'h40270ef8} /* (22, 31, 8) {real, imag} */,
  {32'hc06fb9c0, 32'hbfa24e6c} /* (22, 31, 7) {real, imag} */,
  {32'hbeed0300, 32'h408bb020} /* (22, 31, 6) {real, imag} */,
  {32'h3e699508, 32'hbfcbfe20} /* (22, 31, 5) {real, imag} */,
  {32'hc11ca504, 32'hbec6cc40} /* (22, 31, 4) {real, imag} */,
  {32'hc129e2bf, 32'h40a075e4} /* (22, 31, 3) {real, imag} */,
  {32'hc11a2662, 32'h40ec5b22} /* (22, 31, 2) {real, imag} */,
  {32'hc0433d10, 32'h3fd212c0} /* (22, 31, 1) {real, imag} */,
  {32'h3fd97000, 32'hc15fa7e2} /* (22, 31, 0) {real, imag} */,
  {32'h3fe60cca, 32'h4051e272} /* (22, 30, 31) {real, imag} */,
  {32'h3fa358b0, 32'hbfaa25c8} /* (22, 30, 30) {real, imag} */,
  {32'h40c2d259, 32'hc005f728} /* (22, 30, 29) {real, imag} */,
  {32'h414e7734, 32'hc08eb94b} /* (22, 30, 28) {real, imag} */,
  {32'h415bb433, 32'hc0c24a30} /* (22, 30, 27) {real, imag} */,
  {32'h4141e48b, 32'h4107520c} /* (22, 30, 26) {real, imag} */,
  {32'hbfc25d93, 32'h403c58ec} /* (22, 30, 25) {real, imag} */,
  {32'h4104fdfc, 32'hc08ff359} /* (22, 30, 24) {real, imag} */,
  {32'h413392f9, 32'hbfdd8543} /* (22, 30, 23) {real, imag} */,
  {32'h3d7e1c00, 32'hc10aae0a} /* (22, 30, 22) {real, imag} */,
  {32'hc162c18f, 32'h413cecee} /* (22, 30, 21) {real, imag} */,
  {32'h3e865908, 32'hc0f53ec8} /* (22, 30, 20) {real, imag} */,
  {32'hbfeb2a40, 32'hc11c8e07} /* (22, 30, 19) {real, imag} */,
  {32'hc12767e3, 32'hbffb0a18} /* (22, 30, 18) {real, imag} */,
  {32'hc124975c, 32'h414dc3e6} /* (22, 30, 17) {real, imag} */,
  {32'h3f6fec1e, 32'h3f24bde0} /* (22, 30, 16) {real, imag} */,
  {32'hc0afd22c, 32'hc08637c7} /* (22, 30, 15) {real, imag} */,
  {32'hc196be32, 32'h411bb610} /* (22, 30, 14) {real, imag} */,
  {32'hc19b1eea, 32'hbfee88f4} /* (22, 30, 13) {real, imag} */,
  {32'hc11cc00a, 32'hc0937385} /* (22, 30, 12) {real, imag} */,
  {32'hc0200fe7, 32'hc028e213} /* (22, 30, 11) {real, imag} */,
  {32'h40dbbd05, 32'h40f3df42} /* (22, 30, 10) {real, imag} */,
  {32'h4194ba79, 32'h4154bcbe} /* (22, 30, 9) {real, imag} */,
  {32'h4141752a, 32'h41357c79} /* (22, 30, 8) {real, imag} */,
  {32'h41589aae, 32'hc0f5b4ce} /* (22, 30, 7) {real, imag} */,
  {32'h4179f959, 32'hc079caa5} /* (22, 30, 6) {real, imag} */,
  {32'h402d5c38, 32'hbfce6f0c} /* (22, 30, 5) {real, imag} */,
  {32'h414ea890, 32'h3f7d1a40} /* (22, 30, 4) {real, imag} */,
  {32'h40325650, 32'hc1198f36} /* (22, 30, 3) {real, imag} */,
  {32'hc119faca, 32'hbf92badc} /* (22, 30, 2) {real, imag} */,
  {32'hc0af9b58, 32'h4107bbad} /* (22, 30, 1) {real, imag} */,
  {32'hbea53200, 32'h40e4bb9b} /* (22, 30, 0) {real, imag} */,
  {32'h3d815400, 32'hbfdd45e0} /* (22, 29, 31) {real, imag} */,
  {32'h4103f7ad, 32'hc0c72f4a} /* (22, 29, 30) {real, imag} */,
  {32'h40930616, 32'hc101c1e6} /* (22, 29, 29) {real, imag} */,
  {32'h409669b6, 32'hc1280551} /* (22, 29, 28) {real, imag} */,
  {32'hc03b4eb6, 32'hc13f0762} /* (22, 29, 27) {real, imag} */,
  {32'hc092d474, 32'h3f8900a6} /* (22, 29, 26) {real, imag} */,
  {32'hbf4982f8, 32'hc0346ef2} /* (22, 29, 25) {real, imag} */,
  {32'hc0a8acea, 32'h3f86e87a} /* (22, 29, 24) {real, imag} */,
  {32'hc1143d8d, 32'h40ba0d8a} /* (22, 29, 23) {real, imag} */,
  {32'hc178a385, 32'h40885d41} /* (22, 29, 22) {real, imag} */,
  {32'hc13c5f7a, 32'h412a065b} /* (22, 29, 21) {real, imag} */,
  {32'hc0cc127c, 32'h4116ae33} /* (22, 29, 20) {real, imag} */,
  {32'hbfd78a7d, 32'h4012f24c} /* (22, 29, 19) {real, imag} */,
  {32'h41352002, 32'h3f391420} /* (22, 29, 18) {real, imag} */,
  {32'h41199442, 32'hc0d73da8} /* (22, 29, 17) {real, imag} */,
  {32'h4038128e, 32'hc0fb4d9c} /* (22, 29, 16) {real, imag} */,
  {32'h3f3c1038, 32'h401fd294} /* (22, 29, 15) {real, imag} */,
  {32'hc0a6bae2, 32'h40c99307} /* (22, 29, 14) {real, imag} */,
  {32'h404312da, 32'h410ff0bb} /* (22, 29, 13) {real, imag} */,
  {32'h41384d60, 32'h40651408} /* (22, 29, 12) {real, imag} */,
  {32'hc090f0b3, 32'h3fac5900} /* (22, 29, 11) {real, imag} */,
  {32'hc1724978, 32'h4105ebc0} /* (22, 29, 10) {real, imag} */,
  {32'hc0a309b2, 32'h409e323e} /* (22, 29, 9) {real, imag} */,
  {32'hc063efd6, 32'h40a2a4fa} /* (22, 29, 8) {real, imag} */,
  {32'hc1342c96, 32'hc06c5a0e} /* (22, 29, 7) {real, imag} */,
  {32'hc0f39023, 32'h3fa2d473} /* (22, 29, 6) {real, imag} */,
  {32'h3f505230, 32'hbffbf504} /* (22, 29, 5) {real, imag} */,
  {32'hc057f5e2, 32'hc0ce147b} /* (22, 29, 4) {real, imag} */,
  {32'hc0a2ac27, 32'hc042b08d} /* (22, 29, 3) {real, imag} */,
  {32'h4036af7a, 32'h3fd035d4} /* (22, 29, 2) {real, imag} */,
  {32'h41b2b66f, 32'h4004483a} /* (22, 29, 1) {real, imag} */,
  {32'h4127e8dd, 32'hbf295518} /* (22, 29, 0) {real, imag} */,
  {32'hbff7c85e, 32'hc0b841be} /* (22, 28, 31) {real, imag} */,
  {32'hc0cb7c06, 32'hc13e1e04} /* (22, 28, 30) {real, imag} */,
  {32'hc07bc6a4, 32'h40c17289} /* (22, 28, 29) {real, imag} */,
  {32'hc0386dc9, 32'h4183b096} /* (22, 28, 28) {real, imag} */,
  {32'hbfa8adcf, 32'h40389382} /* (22, 28, 27) {real, imag} */,
  {32'hc0c4d8ce, 32'h3f2e0818} /* (22, 28, 26) {real, imag} */,
  {32'hc01eeb04, 32'h412f1355} /* (22, 28, 25) {real, imag} */,
  {32'hc0e2b042, 32'h4137b368} /* (22, 28, 24) {real, imag} */,
  {32'hc17b60b4, 32'hc12acd60} /* (22, 28, 23) {real, imag} */,
  {32'hc1802174, 32'hc13b71e4} /* (22, 28, 22) {real, imag} */,
  {32'hc1afd708, 32'hc15f8f85} /* (22, 28, 21) {real, imag} */,
  {32'hc15e31f0, 32'hbf6fb5d9} /* (22, 28, 20) {real, imag} */,
  {32'h3fdf964a, 32'hbe47ccb0} /* (22, 28, 19) {real, imag} */,
  {32'h3f9d79a0, 32'hbebf4b90} /* (22, 28, 18) {real, imag} */,
  {32'h40127ca6, 32'h3f9958ad} /* (22, 28, 17) {real, imag} */,
  {32'h41345b5e, 32'hc082997e} /* (22, 28, 16) {real, imag} */,
  {32'h41558dd0, 32'h40d014e2} /* (22, 28, 15) {real, imag} */,
  {32'h40e694d3, 32'hc0c8a511} /* (22, 28, 14) {real, imag} */,
  {32'hc0c6d2ba, 32'hc11714a0} /* (22, 28, 13) {real, imag} */,
  {32'hbe8bf0c0, 32'hc0a9a03a} /* (22, 28, 12) {real, imag} */,
  {32'hc0eff002, 32'hc112e1d4} /* (22, 28, 11) {real, imag} */,
  {32'hc0f42d0a, 32'h40738744} /* (22, 28, 10) {real, imag} */,
  {32'hc00f1dac, 32'h4053fcb4} /* (22, 28, 9) {real, imag} */,
  {32'hbf48d412, 32'h408ce65a} /* (22, 28, 8) {real, imag} */,
  {32'h40978157, 32'h41269512} /* (22, 28, 7) {real, imag} */,
  {32'hbf87d14d, 32'h408318f2} /* (22, 28, 6) {real, imag} */,
  {32'hc0def4fb, 32'h406b0866} /* (22, 28, 5) {real, imag} */,
  {32'hc11f7ea4, 32'h40e42a70} /* (22, 28, 4) {real, imag} */,
  {32'h3f1f622c, 32'h41160be2} /* (22, 28, 3) {real, imag} */,
  {32'h417ce4e4, 32'h3f44c5a5} /* (22, 28, 2) {real, imag} */,
  {32'h3fee5760, 32'h40bc4994} /* (22, 28, 1) {real, imag} */,
  {32'hc0dfb17f, 32'h40ce538c} /* (22, 28, 0) {real, imag} */,
  {32'h3f95a257, 32'h40b23c62} /* (22, 27, 31) {real, imag} */,
  {32'h40d03cb4, 32'h41164678} /* (22, 27, 30) {real, imag} */,
  {32'h40a944a5, 32'h404e938b} /* (22, 27, 29) {real, imag} */,
  {32'h3e5aeb30, 32'h40cbc130} /* (22, 27, 28) {real, imag} */,
  {32'h405728bb, 32'h40fbcf90} /* (22, 27, 27) {real, imag} */,
  {32'h405dbb8d, 32'hc040799d} /* (22, 27, 26) {real, imag} */,
  {32'h402a2064, 32'h40987f52} /* (22, 27, 25) {real, imag} */,
  {32'h4110b616, 32'h417031ba} /* (22, 27, 24) {real, imag} */,
  {32'h41bacc41, 32'h415db524} /* (22, 27, 23) {real, imag} */,
  {32'h4162367c, 32'h4112d4b5} /* (22, 27, 22) {real, imag} */,
  {32'h4116be49, 32'hbe28cc20} /* (22, 27, 21) {real, imag} */,
  {32'h409f28c4, 32'h3f991e0d} /* (22, 27, 20) {real, imag} */,
  {32'h404d2da7, 32'hc0b88dea} /* (22, 27, 19) {real, imag} */,
  {32'h40d6a0d4, 32'h409721a3} /* (22, 27, 18) {real, imag} */,
  {32'h411d870d, 32'h40162db9} /* (22, 27, 17) {real, imag} */,
  {32'hbe8fc588, 32'h3ebfcd2c} /* (22, 27, 16) {real, imag} */,
  {32'hc0c6e68a, 32'hbf73f56c} /* (22, 27, 15) {real, imag} */,
  {32'h401530ba, 32'hc004a698} /* (22, 27, 14) {real, imag} */,
  {32'hc10571a8, 32'h40d72a13} /* (22, 27, 13) {real, imag} */,
  {32'hc16b5180, 32'h406f41f8} /* (22, 27, 12) {real, imag} */,
  {32'h4033ea3a, 32'hc0a9a33b} /* (22, 27, 11) {real, imag} */,
  {32'h3eb23ef4, 32'hc111b1c8} /* (22, 27, 10) {real, imag} */,
  {32'hc065c16a, 32'h3f25f4a8} /* (22, 27, 9) {real, imag} */,
  {32'hc0535cbb, 32'h40dc147e} /* (22, 27, 8) {real, imag} */,
  {32'hc11edf54, 32'h41016a60} /* (22, 27, 7) {real, imag} */,
  {32'hc1453e86, 32'hc0df9967} /* (22, 27, 6) {real, imag} */,
  {32'hbf3911ea, 32'hc0892824} /* (22, 27, 5) {real, imag} */,
  {32'h40da98e2, 32'hbeb26d20} /* (22, 27, 4) {real, imag} */,
  {32'h3efd3b30, 32'h40358cb1} /* (22, 27, 3) {real, imag} */,
  {32'hbee6afb0, 32'h40a76a5c} /* (22, 27, 2) {real, imag} */,
  {32'h40807cc5, 32'h3f3f08ec} /* (22, 27, 1) {real, imag} */,
  {32'h3f881f3c, 32'h4020ddcd} /* (22, 27, 0) {real, imag} */,
  {32'h3f548c46, 32'h3f28b0a4} /* (22, 26, 31) {real, imag} */,
  {32'hc07c90f8, 32'h3e9811f8} /* (22, 26, 30) {real, imag} */,
  {32'h3f0fcbd0, 32'hc0a0a1aa} /* (22, 26, 29) {real, imag} */,
  {32'hbfa20c54, 32'hbffa1a82} /* (22, 26, 28) {real, imag} */,
  {32'h40498430, 32'h40a978cc} /* (22, 26, 27) {real, imag} */,
  {32'hc0673d32, 32'h40084a7e} /* (22, 26, 26) {real, imag} */,
  {32'h40b0bf8e, 32'hc0458556} /* (22, 26, 25) {real, imag} */,
  {32'h412a44cb, 32'hc1021266} /* (22, 26, 24) {real, imag} */,
  {32'h4113657f, 32'hc0a5a0bc} /* (22, 26, 23) {real, imag} */,
  {32'hc0b50c56, 32'h3eb0a4b8} /* (22, 26, 22) {real, imag} */,
  {32'hc0277cac, 32'hc0284b1d} /* (22, 26, 21) {real, imag} */,
  {32'h40da7814, 32'h40e43099} /* (22, 26, 20) {real, imag} */,
  {32'hc0e53a84, 32'h41941cc2} /* (22, 26, 19) {real, imag} */,
  {32'hc04c7eb7, 32'h418e921d} /* (22, 26, 18) {real, imag} */,
  {32'h3f0aad68, 32'h403286a5} /* (22, 26, 17) {real, imag} */,
  {32'hbf8e326e, 32'hc092e514} /* (22, 26, 16) {real, imag} */,
  {32'hc0b942fa, 32'hc00fabb5} /* (22, 26, 15) {real, imag} */,
  {32'hc0d3b666, 32'h4038e9c6} /* (22, 26, 14) {real, imag} */,
  {32'hc13fc0f8, 32'hc0cb6c1f} /* (22, 26, 13) {real, imag} */,
  {32'hc1a28f47, 32'hc0a57d6a} /* (22, 26, 12) {real, imag} */,
  {32'hc0899bb6, 32'h3fec0cd9} /* (22, 26, 11) {real, imag} */,
  {32'hc0716bf8, 32'h3e6c2ff0} /* (22, 26, 10) {real, imag} */,
  {32'hc0fc7ac2, 32'h3fdfac57} /* (22, 26, 9) {real, imag} */,
  {32'h408d1cc8, 32'h40f9905e} /* (22, 26, 8) {real, imag} */,
  {32'hbf2b14e8, 32'h4135b8d2} /* (22, 26, 7) {real, imag} */,
  {32'hc086e62a, 32'hbe9695c8} /* (22, 26, 6) {real, imag} */,
  {32'h40662820, 32'h4011d808} /* (22, 26, 5) {real, imag} */,
  {32'h401da1d0, 32'h406a2942} /* (22, 26, 4) {real, imag} */,
  {32'hc0a287e0, 32'hc04aea32} /* (22, 26, 3) {real, imag} */,
  {32'hc10b31f8, 32'hc06ae030} /* (22, 26, 2) {real, imag} */,
  {32'hc07940c8, 32'h404e875f} /* (22, 26, 1) {real, imag} */,
  {32'hbfd8ab56, 32'hbf971dd7} /* (22, 26, 0) {real, imag} */,
  {32'hc0205c92, 32'hc0992508} /* (22, 25, 31) {real, imag} */,
  {32'hc171b854, 32'hc10ee91c} /* (22, 25, 30) {real, imag} */,
  {32'hc146e451, 32'h40d352f6} /* (22, 25, 29) {real, imag} */,
  {32'hc0b4e83b, 32'h4100a920} /* (22, 25, 28) {real, imag} */,
  {32'h3f9e6f58, 32'h3ff765b4} /* (22, 25, 27) {real, imag} */,
  {32'h3fd68fec, 32'h4056b33d} /* (22, 25, 26) {real, imag} */,
  {32'hc09be4f4, 32'h40692f2f} /* (22, 25, 25) {real, imag} */,
  {32'hc0b7c730, 32'h40033eba} /* (22, 25, 24) {real, imag} */,
  {32'hbfe019ab, 32'hc0495633} /* (22, 25, 23) {real, imag} */,
  {32'h3f0d1df8, 32'h401bb12c} /* (22, 25, 22) {real, imag} */,
  {32'hbf751364, 32'h3f289013} /* (22, 25, 21) {real, imag} */,
  {32'h40467958, 32'h4115fd62} /* (22, 25, 20) {real, imag} */,
  {32'h40383532, 32'h404e2199} /* (22, 25, 19) {real, imag} */,
  {32'h40e95b66, 32'h3f5e5678} /* (22, 25, 18) {real, imag} */,
  {32'h40df809d, 32'h408708d9} /* (22, 25, 17) {real, imag} */,
  {32'h3ed96f68, 32'h40e889cc} /* (22, 25, 16) {real, imag} */,
  {32'h3ffbe72a, 32'hbfe8a637} /* (22, 25, 15) {real, imag} */,
  {32'h40884ea0, 32'h3f2ec904} /* (22, 25, 14) {real, imag} */,
  {32'hc0bdee04, 32'hc0e8d56f} /* (22, 25, 13) {real, imag} */,
  {32'hc067fa32, 32'hc02359fb} /* (22, 25, 12) {real, imag} */,
  {32'h3f204488, 32'hbffa61b0} /* (22, 25, 11) {real, imag} */,
  {32'h3f692d6c, 32'h4066dc12} /* (22, 25, 10) {real, imag} */,
  {32'h4048422b, 32'hbfa65dc0} /* (22, 25, 9) {real, imag} */,
  {32'h4137c17a, 32'hc081a5b3} /* (22, 25, 8) {real, imag} */,
  {32'h418b646e, 32'h3fcc9c20} /* (22, 25, 7) {real, imag} */,
  {32'h4084738b, 32'h3e96d8a8} /* (22, 25, 6) {real, imag} */,
  {32'h40a86d2a, 32'h4024129d} /* (22, 25, 5) {real, imag} */,
  {32'h408bf24c, 32'h40c630ae} /* (22, 25, 4) {real, imag} */,
  {32'h40b2ae4b, 32'h400e3a4a} /* (22, 25, 3) {real, imag} */,
  {32'h40d88b7b, 32'hc01288c0} /* (22, 25, 2) {real, imag} */,
  {32'h40be01e9, 32'h4063263e} /* (22, 25, 1) {real, imag} */,
  {32'h408d2c6e, 32'h412b0399} /* (22, 25, 0) {real, imag} */,
  {32'h3fd07150, 32'h410c4188} /* (22, 24, 31) {real, imag} */,
  {32'h3f8e2125, 32'h40ea4bad} /* (22, 24, 30) {real, imag} */,
  {32'hc091b803, 32'hbf8a4252} /* (22, 24, 29) {real, imag} */,
  {32'hc02ebad4, 32'hc0c17309} /* (22, 24, 28) {real, imag} */,
  {32'h3ff77e18, 32'hc03e2b4e} /* (22, 24, 27) {real, imag} */,
  {32'h40304b60, 32'h409d62f6} /* (22, 24, 26) {real, imag} */,
  {32'h4029c7e5, 32'h405c82d0} /* (22, 24, 25) {real, imag} */,
  {32'h408e168c, 32'hc1431790} /* (22, 24, 24) {real, imag} */,
  {32'h4133b690, 32'hc0b473fa} /* (22, 24, 23) {real, imag} */,
  {32'h40cd68ee, 32'h409715ed} /* (22, 24, 22) {real, imag} */,
  {32'h40ea0241, 32'h40e074ba} /* (22, 24, 21) {real, imag} */,
  {32'h412a7a7b, 32'h40c17c5a} /* (22, 24, 20) {real, imag} */,
  {32'h40b220d5, 32'h40be22c8} /* (22, 24, 19) {real, imag} */,
  {32'hbfedcbf0, 32'h40917555} /* (22, 24, 18) {real, imag} */,
  {32'hc0c689bd, 32'h40480d2c} /* (22, 24, 17) {real, imag} */,
  {32'hc0626405, 32'hbfcbf757} /* (22, 24, 16) {real, imag} */,
  {32'h40c3cc34, 32'hbea58c18} /* (22, 24, 15) {real, imag} */,
  {32'h40f69a3a, 32'h40830ad8} /* (22, 24, 14) {real, imag} */,
  {32'hbd8089f8, 32'h3fedceee} /* (22, 24, 13) {real, imag} */,
  {32'h40f27e77, 32'hc00f53fd} /* (22, 24, 12) {real, imag} */,
  {32'hc02f04e0, 32'hc0837fc4} /* (22, 24, 11) {real, imag} */,
  {32'hc02b731c, 32'hc0089250} /* (22, 24, 10) {real, imag} */,
  {32'h4035e6f4, 32'h40f73a08} /* (22, 24, 9) {real, imag} */,
  {32'h402985c2, 32'h40bc978e} /* (22, 24, 8) {real, imag} */,
  {32'h40d06518, 32'h4084a931} /* (22, 24, 7) {real, imag} */,
  {32'h40e430ad, 32'hbf2335d0} /* (22, 24, 6) {real, imag} */,
  {32'h40bebcf5, 32'h402025fe} /* (22, 24, 5) {real, imag} */,
  {32'h40ddd0ae, 32'h406304e7} /* (22, 24, 4) {real, imag} */,
  {32'hbf7886a9, 32'hbfea1389} /* (22, 24, 3) {real, imag} */,
  {32'h3e2e0610, 32'hc09d3f28} /* (22, 24, 2) {real, imag} */,
  {32'hbf5a27f8, 32'hc0ef803b} /* (22, 24, 1) {real, imag} */,
  {32'h4000f882, 32'hbf84f3aa} /* (22, 24, 0) {real, imag} */,
  {32'h404217b8, 32'hbee88bbe} /* (22, 23, 31) {real, imag} */,
  {32'hbf9bf9fe, 32'hc01c6a89} /* (22, 23, 30) {real, imag} */,
  {32'hc051d1fa, 32'h3e11fde0} /* (22, 23, 29) {real, imag} */,
  {32'h3f85f5cc, 32'h4020a782} /* (22, 23, 28) {real, imag} */,
  {32'h4055040d, 32'h40edea39} /* (22, 23, 27) {real, imag} */,
  {32'h40938b57, 32'h40b333e8} /* (22, 23, 26) {real, imag} */,
  {32'hc020adf1, 32'hbfedef61} /* (22, 23, 25) {real, imag} */,
  {32'h4028c792, 32'hc059b9a8} /* (22, 23, 24) {real, imag} */,
  {32'h4090ed52, 32'h406a3da3} /* (22, 23, 23) {real, imag} */,
  {32'hbd508320, 32'h40010f8e} /* (22, 23, 22) {real, imag} */,
  {32'h3fe56753, 32'h408b354a} /* (22, 23, 21) {real, imag} */,
  {32'h402059a4, 32'h403a9b73} /* (22, 23, 20) {real, imag} */,
  {32'hc01f1563, 32'hc05a9698} /* (22, 23, 19) {real, imag} */,
  {32'hc09c219e, 32'hc07ddb4e} /* (22, 23, 18) {real, imag} */,
  {32'hbf871589, 32'hbdbb2940} /* (22, 23, 17) {real, imag} */,
  {32'hbfc15306, 32'h40cb113e} /* (22, 23, 16) {real, imag} */,
  {32'hc052ed36, 32'h40bbde31} /* (22, 23, 15) {real, imag} */,
  {32'h3f963ff8, 32'hbfa919ae} /* (22, 23, 14) {real, imag} */,
  {32'h40cc26cc, 32'h3f8e3eb4} /* (22, 23, 13) {real, imag} */,
  {32'h400438cc, 32'h40817f92} /* (22, 23, 12) {real, imag} */,
  {32'h3f85601a, 32'h409f37dd} /* (22, 23, 11) {real, imag} */,
  {32'h3f47e9c4, 32'h4081db97} /* (22, 23, 10) {real, imag} */,
  {32'h4046e6a9, 32'h40c4f8e4} /* (22, 23, 9) {real, imag} */,
  {32'h408ddfb2, 32'h410850f4} /* (22, 23, 8) {real, imag} */,
  {32'h3e494fc0, 32'h40b0f20a} /* (22, 23, 7) {real, imag} */,
  {32'hc0f31dad, 32'h40ebbf82} /* (22, 23, 6) {real, imag} */,
  {32'hc0b36cca, 32'h40c11c66} /* (22, 23, 5) {real, imag} */,
  {32'h400de5b8, 32'hbfb5f54e} /* (22, 23, 4) {real, imag} */,
  {32'hc0a715bd, 32'h3fcd7cfc} /* (22, 23, 3) {real, imag} */,
  {32'hc1025543, 32'hbfc1e938} /* (22, 23, 2) {real, imag} */,
  {32'h3fb9f0fd, 32'hc1359e54} /* (22, 23, 1) {real, imag} */,
  {32'h40188fa3, 32'hc125b7d1} /* (22, 23, 0) {real, imag} */,
  {32'h3e8c23cc, 32'hc02a644c} /* (22, 22, 31) {real, imag} */,
  {32'h3fe3ec3b, 32'h40014ca3} /* (22, 22, 30) {real, imag} */,
  {32'hbf9b49c0, 32'h405f3cfa} /* (22, 22, 29) {real, imag} */,
  {32'hc0741ed6, 32'hc04ec0a5} /* (22, 22, 28) {real, imag} */,
  {32'h3fc83ebc, 32'hbfe3a8e2} /* (22, 22, 27) {real, imag} */,
  {32'hbeef1884, 32'h405eebdc} /* (22, 22, 26) {real, imag} */,
  {32'hc061fecd, 32'h406bc657} /* (22, 22, 25) {real, imag} */,
  {32'hbfee2796, 32'h3f9883f2} /* (22, 22, 24) {real, imag} */,
  {32'hc08d10c2, 32'hc08103a2} /* (22, 22, 23) {real, imag} */,
  {32'hc130b541, 32'hc04eb213} /* (22, 22, 22) {real, imag} */,
  {32'hbfb6fade, 32'hbf35ac04} /* (22, 22, 21) {real, imag} */,
  {32'h408dfd92, 32'hbea9b100} /* (22, 22, 20) {real, imag} */,
  {32'hbf113018, 32'h400bddd2} /* (22, 22, 19) {real, imag} */,
  {32'hc01750b9, 32'h4037ff1c} /* (22, 22, 18) {real, imag} */,
  {32'hc0006be9, 32'h3eacd950} /* (22, 22, 17) {real, imag} */,
  {32'hc0ecbbc6, 32'hc07c309b} /* (22, 22, 16) {real, imag} */,
  {32'hc017d678, 32'h4074e7c7} /* (22, 22, 15) {real, imag} */,
  {32'hc09d2513, 32'h408ee7a7} /* (22, 22, 14) {real, imag} */,
  {32'hc0847c80, 32'hbf52d27f} /* (22, 22, 13) {real, imag} */,
  {32'h3c005900, 32'hc0ab0c89} /* (22, 22, 12) {real, imag} */,
  {32'h40be252e, 32'hbf8ecae7} /* (22, 22, 11) {real, imag} */,
  {32'h40745d9f, 32'hbff14ca2} /* (22, 22, 10) {real, imag} */,
  {32'hbf23083e, 32'hc04a426d} /* (22, 22, 9) {real, imag} */,
  {32'hc025b6bc, 32'h409ec1c8} /* (22, 22, 8) {real, imag} */,
  {32'hc0970830, 32'hc0174b62} /* (22, 22, 7) {real, imag} */,
  {32'hc03484b9, 32'hbfe92a40} /* (22, 22, 6) {real, imag} */,
  {32'h3f858a6d, 32'hbf6141a8} /* (22, 22, 5) {real, imag} */,
  {32'h40b5adce, 32'h3f287ca0} /* (22, 22, 4) {real, imag} */,
  {32'h4110adab, 32'hbff6b2b2} /* (22, 22, 3) {real, imag} */,
  {32'h40841d6a, 32'hbfe9bee4} /* (22, 22, 2) {real, imag} */,
  {32'h40622649, 32'h409ecec6} /* (22, 22, 1) {real, imag} */,
  {32'h40b796f8, 32'h400a603c} /* (22, 22, 0) {real, imag} */,
  {32'hbeb0555c, 32'h4019b828} /* (22, 21, 31) {real, imag} */,
  {32'h4084b20a, 32'h3fdefef9} /* (22, 21, 30) {real, imag} */,
  {32'h404fc387, 32'hc0856e3c} /* (22, 21, 29) {real, imag} */,
  {32'h40814734, 32'hc092ae16} /* (22, 21, 28) {real, imag} */,
  {32'h3f7f4bc0, 32'h3fc20710} /* (22, 21, 27) {real, imag} */,
  {32'hc084b48a, 32'h40927aba} /* (22, 21, 26) {real, imag} */,
  {32'hc0b646b3, 32'h3fb5577a} /* (22, 21, 25) {real, imag} */,
  {32'h3f675b38, 32'h40448fa6} /* (22, 21, 24) {real, imag} */,
  {32'h40561c3a, 32'h3eee1924} /* (22, 21, 23) {real, imag} */,
  {32'hbe1de240, 32'hbec3e588} /* (22, 21, 22) {real, imag} */,
  {32'hc0a3911f, 32'hc105d556} /* (22, 21, 21) {real, imag} */,
  {32'hc070d050, 32'hc12a1e00} /* (22, 21, 20) {real, imag} */,
  {32'hbf51f5d0, 32'hc084ca4d} /* (22, 21, 19) {real, imag} */,
  {32'hc050f386, 32'h401b88c4} /* (22, 21, 18) {real, imag} */,
  {32'hbf2c0bd2, 32'hbe348c88} /* (22, 21, 17) {real, imag} */,
  {32'hc0588f08, 32'hbfdb22fd} /* (22, 21, 16) {real, imag} */,
  {32'hbfc2613c, 32'h402500e9} /* (22, 21, 15) {real, imag} */,
  {32'h3f042a84, 32'h40656618} /* (22, 21, 14) {real, imag} */,
  {32'h405b56ab, 32'hc05635fe} /* (22, 21, 13) {real, imag} */,
  {32'h403761eb, 32'hc0bcfe45} /* (22, 21, 12) {real, imag} */,
  {32'h409d833f, 32'hc0018352} /* (22, 21, 11) {real, imag} */,
  {32'h3fa8e39d, 32'h4019a5a6} /* (22, 21, 10) {real, imag} */,
  {32'hc106f860, 32'hbf9e5abe} /* (22, 21, 9) {real, imag} */,
  {32'hc094565a, 32'hc0b7d25c} /* (22, 21, 8) {real, imag} */,
  {32'hbff7366c, 32'hc104f327} /* (22, 21, 7) {real, imag} */,
  {32'hbfe41b4e, 32'hbf03dda0} /* (22, 21, 6) {real, imag} */,
  {32'h40b5a131, 32'h3ff00a9a} /* (22, 21, 5) {real, imag} */,
  {32'hc040b063, 32'hbf6e3b10} /* (22, 21, 4) {real, imag} */,
  {32'hc0c66d33, 32'h40b90ed8} /* (22, 21, 3) {real, imag} */,
  {32'h3f1be60f, 32'h41474d78} /* (22, 21, 2) {real, imag} */,
  {32'hc04b5a77, 32'h40b7ceee} /* (22, 21, 1) {real, imag} */,
  {32'hc0edb373, 32'h3ee3054c} /* (22, 21, 0) {real, imag} */,
  {32'hbf65e72e, 32'hbee31c30} /* (22, 20, 31) {real, imag} */,
  {32'hbf138d02, 32'hc0c05ee6} /* (22, 20, 30) {real, imag} */,
  {32'hbf284b92, 32'hc0632322} /* (22, 20, 29) {real, imag} */,
  {32'hc0303b2d, 32'h40931938} /* (22, 20, 28) {real, imag} */,
  {32'hc080f176, 32'h40c1389e} /* (22, 20, 27) {real, imag} */,
  {32'hc13aabfe, 32'hbfe87660} /* (22, 20, 26) {real, imag} */,
  {32'hc0979d98, 32'hc0341dee} /* (22, 20, 25) {real, imag} */,
  {32'hc09f29f4, 32'hbda906d0} /* (22, 20, 24) {real, imag} */,
  {32'hc0847a6c, 32'h4047579f} /* (22, 20, 23) {real, imag} */,
  {32'hc0171f2c, 32'h3fb822a8} /* (22, 20, 22) {real, imag} */,
  {32'hbf17c260, 32'hc034df5d} /* (22, 20, 21) {real, imag} */,
  {32'hc0aa9d54, 32'hbf18d227} /* (22, 20, 20) {real, imag} */,
  {32'hc0653195, 32'hc0479c4c} /* (22, 20, 19) {real, imag} */,
  {32'hbfc6499f, 32'hbfc546ac} /* (22, 20, 18) {real, imag} */,
  {32'h3c843d00, 32'h40214c2e} /* (22, 20, 17) {real, imag} */,
  {32'h3f6f2192, 32'h40841709} /* (22, 20, 16) {real, imag} */,
  {32'h408bdf85, 32'h3fa3f789} /* (22, 20, 15) {real, imag} */,
  {32'h3ffa706c, 32'hc04e2610} /* (22, 20, 14) {real, imag} */,
  {32'hc0855e98, 32'hbfefae60} /* (22, 20, 13) {real, imag} */,
  {32'hc08927f8, 32'h40073c7b} /* (22, 20, 12) {real, imag} */,
  {32'hbfd46a5d, 32'hbf1c2958} /* (22, 20, 11) {real, imag} */,
  {32'h40512a60, 32'hc00dab07} /* (22, 20, 10) {real, imag} */,
  {32'h400a3b14, 32'h40086fea} /* (22, 20, 9) {real, imag} */,
  {32'hbfdcc20d, 32'h409adf36} /* (22, 20, 8) {real, imag} */,
  {32'hc00eb81e, 32'hc02bf2bf} /* (22, 20, 7) {real, imag} */,
  {32'hc039a38a, 32'hc0e8025a} /* (22, 20, 6) {real, imag} */,
  {32'hbf721ea4, 32'hbf0c0180} /* (22, 20, 5) {real, imag} */,
  {32'hbe2c4c28, 32'h4030ad9b} /* (22, 20, 4) {real, imag} */,
  {32'h4059dad3, 32'h4096e2e0} /* (22, 20, 3) {real, imag} */,
  {32'h40847b77, 32'h4085b536} /* (22, 20, 2) {real, imag} */,
  {32'h3ed2c6d8, 32'hbfce1c98} /* (22, 20, 1) {real, imag} */,
  {32'h3f996dbc, 32'hbfa04221} /* (22, 20, 0) {real, imag} */,
  {32'h402035dd, 32'h4002f503} /* (22, 19, 31) {real, imag} */,
  {32'h3f8b4096, 32'h3f33b6f8} /* (22, 19, 30) {real, imag} */,
  {32'h3eaf8b20, 32'hbf22ad7a} /* (22, 19, 29) {real, imag} */,
  {32'h4062a1d6, 32'h3ebd3ed0} /* (22, 19, 28) {real, imag} */,
  {32'h3f9e85f7, 32'hc03f01c1} /* (22, 19, 27) {real, imag} */,
  {32'hbeff8e66, 32'hc05a2544} /* (22, 19, 26) {real, imag} */,
  {32'hbf2796a8, 32'hc0962d2e} /* (22, 19, 25) {real, imag} */,
  {32'hc0647c32, 32'hc05517b9} /* (22, 19, 24) {real, imag} */,
  {32'hc00929dc, 32'hbfca1051} /* (22, 19, 23) {real, imag} */,
  {32'hbf983814, 32'hc005739e} /* (22, 19, 22) {real, imag} */,
  {32'hbf93193c, 32'hc0839354} /* (22, 19, 21) {real, imag} */,
  {32'hbe90e904, 32'hbfd5c714} /* (22, 19, 20) {real, imag} */,
  {32'h40086eca, 32'hc018f0f2} /* (22, 19, 19) {real, imag} */,
  {32'h3f1376b4, 32'h3f57ee12} /* (22, 19, 18) {real, imag} */,
  {32'h401f348a, 32'hc05b3849} /* (22, 19, 17) {real, imag} */,
  {32'hbf9c78f0, 32'hbf54e466} /* (22, 19, 16) {real, imag} */,
  {32'hbfed5d97, 32'hbcfdf420} /* (22, 19, 15) {real, imag} */,
  {32'h401ab059, 32'hc08830ad} /* (22, 19, 14) {real, imag} */,
  {32'h405102b6, 32'hc06af39a} /* (22, 19, 13) {real, imag} */,
  {32'h3eb83c80, 32'hbf7b2d95} /* (22, 19, 12) {real, imag} */,
  {32'hbfc7cc5a, 32'hc05a5079} /* (22, 19, 11) {real, imag} */,
  {32'hbf0b8e7e, 32'h3ea36494} /* (22, 19, 10) {real, imag} */,
  {32'hc05cacda, 32'hbdc39e20} /* (22, 19, 9) {real, imag} */,
  {32'hbfc9b668, 32'h40451905} /* (22, 19, 8) {real, imag} */,
  {32'h3f531e3c, 32'h3f7956f0} /* (22, 19, 7) {real, imag} */,
  {32'h40935df5, 32'h3d0f63e0} /* (22, 19, 6) {real, imag} */,
  {32'h40279b2a, 32'hbf86910d} /* (22, 19, 5) {real, imag} */,
  {32'h3ec1d370, 32'hbebd2850} /* (22, 19, 4) {real, imag} */,
  {32'h3faba9b0, 32'hbf374e14} /* (22, 19, 3) {real, imag} */,
  {32'hc05c8fd8, 32'h3ee91778} /* (22, 19, 2) {real, imag} */,
  {32'h3f8dda9c, 32'hbed8f534} /* (22, 19, 1) {real, imag} */,
  {32'h40264eb6, 32'hbfc53e26} /* (22, 19, 0) {real, imag} */,
  {32'hbfd27ae2, 32'hc092198c} /* (22, 18, 31) {real, imag} */,
  {32'hbf909810, 32'hc09cf03a} /* (22, 18, 30) {real, imag} */,
  {32'h3fe4cce4, 32'hc002e800} /* (22, 18, 29) {real, imag} */,
  {32'hbfe09728, 32'hbf8f8031} /* (22, 18, 28) {real, imag} */,
  {32'h3f8ee9a4, 32'hbf55678c} /* (22, 18, 27) {real, imag} */,
  {32'hbf42567e, 32'hc002eb14} /* (22, 18, 26) {real, imag} */,
  {32'hc01c3994, 32'hc0b23bc8} /* (22, 18, 25) {real, imag} */,
  {32'h3e869562, 32'hc0c2c00a} /* (22, 18, 24) {real, imag} */,
  {32'h3ff45b7e, 32'hc0341603} /* (22, 18, 23) {real, imag} */,
  {32'h3fcabcb0, 32'h4030bb55} /* (22, 18, 22) {real, imag} */,
  {32'h4034e011, 32'h400152d5} /* (22, 18, 21) {real, imag} */,
  {32'h3fc644a6, 32'h3f8e2fdb} /* (22, 18, 20) {real, imag} */,
  {32'h3d99d9e0, 32'h402518d4} /* (22, 18, 19) {real, imag} */,
  {32'hbfcf7a08, 32'h401bf550} /* (22, 18, 18) {real, imag} */,
  {32'h3e5b72d0, 32'h3fd32346} /* (22, 18, 17) {real, imag} */,
  {32'h40800cb0, 32'hbec29d60} /* (22, 18, 16) {real, imag} */,
  {32'h3f418300, 32'hbea3df84} /* (22, 18, 15) {real, imag} */,
  {32'h3f9617b8, 32'hc01d963e} /* (22, 18, 14) {real, imag} */,
  {32'h3f1dbef8, 32'hbf78a15e} /* (22, 18, 13) {real, imag} */,
  {32'hc054396a, 32'h3f76ff66} /* (22, 18, 12) {real, imag} */,
  {32'hc0690279, 32'h3f8e0586} /* (22, 18, 11) {real, imag} */,
  {32'hbed50b20, 32'h3ffbbe36} /* (22, 18, 10) {real, imag} */,
  {32'hc0078b5b, 32'h3fe6641b} /* (22, 18, 9) {real, imag} */,
  {32'h3ecfb7b0, 32'h3df2e9c0} /* (22, 18, 8) {real, imag} */,
  {32'hbf6d671d, 32'h3f8a323a} /* (22, 18, 7) {real, imag} */,
  {32'hbe602938, 32'hbda69870} /* (22, 18, 6) {real, imag} */,
  {32'hc0927851, 32'hbf28046b} /* (22, 18, 5) {real, imag} */,
  {32'hc0372571, 32'h406f7dd4} /* (22, 18, 4) {real, imag} */,
  {32'hc023a69d, 32'hbfec94a0} /* (22, 18, 3) {real, imag} */,
  {32'hc0051589, 32'hc08fcf61} /* (22, 18, 2) {real, imag} */,
  {32'hbea9d540, 32'h3f40a8e4} /* (22, 18, 1) {real, imag} */,
  {32'hbf187a3c, 32'h3f0201e3} /* (22, 18, 0) {real, imag} */,
  {32'h3f475d41, 32'hbf43ab8f} /* (22, 17, 31) {real, imag} */,
  {32'h3edea868, 32'hbe1aad60} /* (22, 17, 30) {real, imag} */,
  {32'hc009a71b, 32'hbfd8bc56} /* (22, 17, 29) {real, imag} */,
  {32'hc0716320, 32'hbfdaacd6} /* (22, 17, 28) {real, imag} */,
  {32'hbf412d2a, 32'hc00ebe81} /* (22, 17, 27) {real, imag} */,
  {32'h3f80e6ca, 32'hbf87774e} /* (22, 17, 26) {real, imag} */,
  {32'hbf5e54cc, 32'hbf80cb11} /* (22, 17, 25) {real, imag} */,
  {32'hc03e0ea0, 32'h3ff07fc4} /* (22, 17, 24) {real, imag} */,
  {32'h3f519884, 32'h400366c1} /* (22, 17, 23) {real, imag} */,
  {32'h3fe74a37, 32'hbfdc248c} /* (22, 17, 22) {real, imag} */,
  {32'hbf5326ae, 32'hbfdeace8} /* (22, 17, 21) {real, imag} */,
  {32'hbf741b60, 32'hbfd72096} /* (22, 17, 20) {real, imag} */,
  {32'hbfe09587, 32'hbf9db052} /* (22, 17, 19) {real, imag} */,
  {32'h404fb6e4, 32'hbe9c4f60} /* (22, 17, 18) {real, imag} */,
  {32'hbf94101e, 32'h3f909ff0} /* (22, 17, 17) {real, imag} */,
  {32'hbf39fe25, 32'hc02362d0} /* (22, 17, 16) {real, imag} */,
  {32'h3ed3ed90, 32'hbfdf6314} /* (22, 17, 15) {real, imag} */,
  {32'hbf97657d, 32'h3f6c04cc} /* (22, 17, 14) {real, imag} */,
  {32'h40bdac3d, 32'hbf6557c6} /* (22, 17, 13) {real, imag} */,
  {32'h402900df, 32'hc058b332} /* (22, 17, 12) {real, imag} */,
  {32'hc033cd11, 32'h3e659780} /* (22, 17, 11) {real, imag} */,
  {32'hbfbf7ad2, 32'h3f77fe3e} /* (22, 17, 10) {real, imag} */,
  {32'h3fcdc49d, 32'hc030bf26} /* (22, 17, 9) {real, imag} */,
  {32'h400dfbb0, 32'hc03ac6af} /* (22, 17, 8) {real, imag} */,
  {32'hc02ccaa6, 32'hbfa419dd} /* (22, 17, 7) {real, imag} */,
  {32'hc007e2f6, 32'h400a882d} /* (22, 17, 6) {real, imag} */,
  {32'h3edaa47a, 32'h4010bb43} /* (22, 17, 5) {real, imag} */,
  {32'h403656ec, 32'hbd1c8800} /* (22, 17, 4) {real, imag} */,
  {32'h3f6c912a, 32'hbf492a94} /* (22, 17, 3) {real, imag} */,
  {32'hbf871419, 32'hc03ebfb1} /* (22, 17, 2) {real, imag} */,
  {32'h3fb2d982, 32'hc0239b3f} /* (22, 17, 1) {real, imag} */,
  {32'h4007856a, 32'hc002b936} /* (22, 17, 0) {real, imag} */,
  {32'h3fa27a58, 32'h40114148} /* (22, 16, 31) {real, imag} */,
  {32'h3fc167e3, 32'h40880e50} /* (22, 16, 30) {real, imag} */,
  {32'h3fd6e30c, 32'h409f932b} /* (22, 16, 29) {real, imag} */,
  {32'h4048df54, 32'h40537120} /* (22, 16, 28) {real, imag} */,
  {32'h3e869b20, 32'hbff60c94} /* (22, 16, 27) {real, imag} */,
  {32'hbf570474, 32'hbe9fdf90} /* (22, 16, 26) {real, imag} */,
  {32'h3dc20fe0, 32'h3f48d922} /* (22, 16, 25) {real, imag} */,
  {32'hbfb20df7, 32'hbfcc9d78} /* (22, 16, 24) {real, imag} */,
  {32'hbf21f410, 32'h3db81900} /* (22, 16, 23) {real, imag} */,
  {32'h3f8f064c, 32'h3fd327c4} /* (22, 16, 22) {real, imag} */,
  {32'h3fb60d51, 32'h3fea63ec} /* (22, 16, 21) {real, imag} */,
  {32'h4044b690, 32'h3f4a21ec} /* (22, 16, 20) {real, imag} */,
  {32'h3fed1a9c, 32'hbe91eac0} /* (22, 16, 19) {real, imag} */,
  {32'h3f3b8220, 32'h3fba2184} /* (22, 16, 18) {real, imag} */,
  {32'hbfaa6790, 32'h3f49f844} /* (22, 16, 17) {real, imag} */,
  {32'hbe225d88, 32'h3f96b6da} /* (22, 16, 16) {real, imag} */,
  {32'h405b2283, 32'h3f4f6f20} /* (22, 16, 15) {real, imag} */,
  {32'h40419d50, 32'hbfa38f9c} /* (22, 16, 14) {real, imag} */,
  {32'hbf8374e0, 32'hbf85c602} /* (22, 16, 13) {real, imag} */,
  {32'hc085fd46, 32'hbf3285e4} /* (22, 16, 12) {real, imag} */,
  {32'h3f7cf89c, 32'hbf19f8c0} /* (22, 16, 11) {real, imag} */,
  {32'h3f46c24c, 32'hc0303b5c} /* (22, 16, 10) {real, imag} */,
  {32'h3e0a34c0, 32'hc08942f8} /* (22, 16, 9) {real, imag} */,
  {32'hbfc7243e, 32'hbf3922d8} /* (22, 16, 8) {real, imag} */,
  {32'h3fbd94bc, 32'h3fbf67c9} /* (22, 16, 7) {real, imag} */,
  {32'h3f43d8f0, 32'h3f7e4bc3} /* (22, 16, 6) {real, imag} */,
  {32'hbec059b4, 32'hbf7394ec} /* (22, 16, 5) {real, imag} */,
  {32'hbed7ee50, 32'hc038d757} /* (22, 16, 4) {real, imag} */,
  {32'hbf4b0ff3, 32'hc084400e} /* (22, 16, 3) {real, imag} */,
  {32'h3f9e54e4, 32'hc02b056c} /* (22, 16, 2) {real, imag} */,
  {32'h3f8c30c0, 32'hc007ebdc} /* (22, 16, 1) {real, imag} */,
  {32'h3f8dc855, 32'hbfdfc66c} /* (22, 16, 0) {real, imag} */,
  {32'hbf58a179, 32'hbe4a82a4} /* (22, 15, 31) {real, imag} */,
  {32'h3f079394, 32'h3f6ab1b8} /* (22, 15, 30) {real, imag} */,
  {32'h404a159d, 32'h3f57ea8c} /* (22, 15, 29) {real, imag} */,
  {32'h406da47c, 32'h3efd0708} /* (22, 15, 28) {real, imag} */,
  {32'hbe51bbf8, 32'h3ee0dd58} /* (22, 15, 27) {real, imag} */,
  {32'hc092aa8c, 32'hbe79a2f0} /* (22, 15, 26) {real, imag} */,
  {32'hbf189a04, 32'h3e8535f4} /* (22, 15, 25) {real, imag} */,
  {32'hbd047be0, 32'hc068809a} /* (22, 15, 24) {real, imag} */,
  {32'hbfe4be4a, 32'hc026b491} /* (22, 15, 23) {real, imag} */,
  {32'h3f579f0a, 32'hbfa07354} /* (22, 15, 22) {real, imag} */,
  {32'h40139e7e, 32'hbf3515c8} /* (22, 15, 21) {real, imag} */,
  {32'h3e8378c0, 32'h40161c7b} /* (22, 15, 20) {real, imag} */,
  {32'hbf623882, 32'h405cefdb} /* (22, 15, 19) {real, imag} */,
  {32'h3f8dd910, 32'h404286a0} /* (22, 15, 18) {real, imag} */,
  {32'h400d8fe7, 32'h3ff1b7b8} /* (22, 15, 17) {real, imag} */,
  {32'hbfa6575c, 32'h3f9c8958} /* (22, 15, 16) {real, imag} */,
  {32'hbdbbd1e0, 32'hbebd4810} /* (22, 15, 15) {real, imag} */,
  {32'h4031154c, 32'hbf8875c8} /* (22, 15, 14) {real, imag} */,
  {32'h3e067540, 32'h3ed2080c} /* (22, 15, 13) {real, imag} */,
  {32'h3f8a9812, 32'h402c2d92} /* (22, 15, 12) {real, imag} */,
  {32'h3fce1482, 32'h3fafe464} /* (22, 15, 11) {real, imag} */,
  {32'hbf570b54, 32'hbff73ff7} /* (22, 15, 10) {real, imag} */,
  {32'h3f61973e, 32'hc027011e} /* (22, 15, 9) {real, imag} */,
  {32'h3dc4bab0, 32'hc0289e53} /* (22, 15, 8) {real, imag} */,
  {32'h3f8e29b1, 32'hc03f4c1e} /* (22, 15, 7) {real, imag} */,
  {32'h3f9d45e8, 32'hbfe92864} /* (22, 15, 6) {real, imag} */,
  {32'h3fefbd68, 32'h3f163914} /* (22, 15, 5) {real, imag} */,
  {32'h3dbfae90, 32'h3f9e87e0} /* (22, 15, 4) {real, imag} */,
  {32'hc01ed26a, 32'hbf60aa44} /* (22, 15, 3) {real, imag} */,
  {32'hbddaded0, 32'h3fc3abae} /* (22, 15, 2) {real, imag} */,
  {32'hbe33b830, 32'h40210c71} /* (22, 15, 1) {real, imag} */,
  {32'h3f4c4708, 32'h3f354078} /* (22, 15, 0) {real, imag} */,
  {32'h3f003b14, 32'h3f1064e4} /* (22, 14, 31) {real, imag} */,
  {32'h3f170ad0, 32'h3f082b7c} /* (22, 14, 30) {real, imag} */,
  {32'hbe43971c, 32'h3ffeffb8} /* (22, 14, 29) {real, imag} */,
  {32'hbf581560, 32'hbeb182f4} /* (22, 14, 28) {real, imag} */,
  {32'hbfa51884, 32'h3fc8badc} /* (22, 14, 27) {real, imag} */,
  {32'hbe74a438, 32'h405a5dd8} /* (22, 14, 26) {real, imag} */,
  {32'h40208ca0, 32'h3ff139ce} /* (22, 14, 25) {real, imag} */,
  {32'h3f827eb0, 32'h409ff7c8} /* (22, 14, 24) {real, imag} */,
  {32'hbfd6ac06, 32'h40867f93} /* (22, 14, 23) {real, imag} */,
  {32'h3f52f3a0, 32'h3ffd7526} /* (22, 14, 22) {real, imag} */,
  {32'hbfea83ce, 32'h40236ac1} /* (22, 14, 21) {real, imag} */,
  {32'hbd85fba0, 32'h3fe4d4b5} /* (22, 14, 20) {real, imag} */,
  {32'h3fcbcd82, 32'h3f9732d4} /* (22, 14, 19) {real, imag} */,
  {32'hc057ab8e, 32'h4048080c} /* (22, 14, 18) {real, imag} */,
  {32'hc067334b, 32'hc00aed41} /* (22, 14, 17) {real, imag} */,
  {32'hc00a1dcc, 32'hc02658a2} /* (22, 14, 16) {real, imag} */,
  {32'hbf6c1710, 32'hbf163b96} /* (22, 14, 15) {real, imag} */,
  {32'h3fd69eb8, 32'hc0348028} /* (22, 14, 14) {real, imag} */,
  {32'h3e7b60e0, 32'hbfd6ff81} /* (22, 14, 13) {real, imag} */,
  {32'hc03dc8fe, 32'hbf3dc7a2} /* (22, 14, 12) {real, imag} */,
  {32'hc05f4ca5, 32'h408afd62} /* (22, 14, 11) {real, imag} */,
  {32'hc084cc10, 32'h3f346c34} /* (22, 14, 10) {real, imag} */,
  {32'h3e19e6b0, 32'h3e741b28} /* (22, 14, 9) {real, imag} */,
  {32'h3f531928, 32'h4062549a} /* (22, 14, 8) {real, imag} */,
  {32'h3f00ba0d, 32'hbf3ceec4} /* (22, 14, 7) {real, imag} */,
  {32'h3fac9707, 32'hbfb3df4f} /* (22, 14, 6) {real, imag} */,
  {32'hbf99b2e0, 32'h3fd7c01a} /* (22, 14, 5) {real, imag} */,
  {32'hbed3afb8, 32'hbef163c0} /* (22, 14, 4) {real, imag} */,
  {32'hbf08ba74, 32'hbfd31270} /* (22, 14, 3) {real, imag} */,
  {32'hbfc52da6, 32'h3edad2e0} /* (22, 14, 2) {real, imag} */,
  {32'h40949ed8, 32'hbbc4c600} /* (22, 14, 1) {real, imag} */,
  {32'h40662821, 32'hbf4365fd} /* (22, 14, 0) {real, imag} */,
  {32'hbf1328dc, 32'h3ebaf958} /* (22, 13, 31) {real, imag} */,
  {32'hc0300a55, 32'hbf482528} /* (22, 13, 30) {real, imag} */,
  {32'hbffd9118, 32'hbf3f093a} /* (22, 13, 29) {real, imag} */,
  {32'h402ff038, 32'hc00d078e} /* (22, 13, 28) {real, imag} */,
  {32'h4003f97c, 32'h3ef70818} /* (22, 13, 27) {real, imag} */,
  {32'hbf6b3d6b, 32'h41001603} /* (22, 13, 26) {real, imag} */,
  {32'hbf94d084, 32'h408e12a4} /* (22, 13, 25) {real, imag} */,
  {32'hc05a4284, 32'h4097264e} /* (22, 13, 24) {real, imag} */,
  {32'hbf5fa542, 32'hbf37251a} /* (22, 13, 23) {real, imag} */,
  {32'h3fe95f7c, 32'h3f85fd2f} /* (22, 13, 22) {real, imag} */,
  {32'hbebba270, 32'h3f0ac094} /* (22, 13, 21) {real, imag} */,
  {32'hbfcd0031, 32'hc05f2328} /* (22, 13, 20) {real, imag} */,
  {32'hc0016706, 32'hc04682c8} /* (22, 13, 19) {real, imag} */,
  {32'hc07cd7ef, 32'hbf0fdc42} /* (22, 13, 18) {real, imag} */,
  {32'h3f95dd19, 32'h3ff012f6} /* (22, 13, 17) {real, imag} */,
  {32'h40a8ad42, 32'hbfa987d1} /* (22, 13, 16) {real, imag} */,
  {32'h3f568942, 32'hbe20fa44} /* (22, 13, 15) {real, imag} */,
  {32'hc07d195d, 32'h3f17ec48} /* (22, 13, 14) {real, imag} */,
  {32'hc08164f9, 32'hbfb6e704} /* (22, 13, 13) {real, imag} */,
  {32'hbfa84d00, 32'h3f750077} /* (22, 13, 12) {real, imag} */,
  {32'hbf4f9ebc, 32'h408a8f54} /* (22, 13, 11) {real, imag} */,
  {32'h3fcc1327, 32'h4085b1c9} /* (22, 13, 10) {real, imag} */,
  {32'h3fda0944, 32'h403be550} /* (22, 13, 9) {real, imag} */,
  {32'hbff7d410, 32'hbfb2680a} /* (22, 13, 8) {real, imag} */,
  {32'hc007c2c1, 32'hc0bae044} /* (22, 13, 7) {real, imag} */,
  {32'h40afbd4b, 32'hc06ec7ce} /* (22, 13, 6) {real, imag} */,
  {32'h3f5d0048, 32'hc0685826} /* (22, 13, 5) {real, imag} */,
  {32'hc038e0a6, 32'h40073312} /* (22, 13, 4) {real, imag} */,
  {32'hc0508906, 32'h3fdc8e76} /* (22, 13, 3) {real, imag} */,
  {32'h40618776, 32'hc02fd7e1} /* (22, 13, 2) {real, imag} */,
  {32'h3f9825cc, 32'hbfccf5db} /* (22, 13, 1) {real, imag} */,
  {32'h3fe544a4, 32'hbea14bf0} /* (22, 13, 0) {real, imag} */,
  {32'h3ffbf5b9, 32'hbfde0684} /* (22, 12, 31) {real, imag} */,
  {32'h3fdcbe93, 32'hc0013df4} /* (22, 12, 30) {real, imag} */,
  {32'hc0029084, 32'hc06f9546} /* (22, 12, 29) {real, imag} */,
  {32'h40961e4e, 32'hc0dd53e8} /* (22, 12, 28) {real, imag} */,
  {32'h40c1572a, 32'hbfbc46aa} /* (22, 12, 27) {real, imag} */,
  {32'h409e5758, 32'h3f8ea73e} /* (22, 12, 26) {real, imag} */,
  {32'h3fbda064, 32'h3dadbc10} /* (22, 12, 25) {real, imag} */,
  {32'hbff9b7ad, 32'hc042d3be} /* (22, 12, 24) {real, imag} */,
  {32'hbe8901e0, 32'hc01ba885} /* (22, 12, 23) {real, imag} */,
  {32'hbf86dc98, 32'hc07953ea} /* (22, 12, 22) {real, imag} */,
  {32'hc0498174, 32'hc026fe25} /* (22, 12, 21) {real, imag} */,
  {32'hbfe20546, 32'h401071a0} /* (22, 12, 20) {real, imag} */,
  {32'hbfef410a, 32'hbf0d15f0} /* (22, 12, 19) {real, imag} */,
  {32'h4059cd78, 32'hbede4ff8} /* (22, 12, 18) {real, imag} */,
  {32'h4083ebd1, 32'hbef3eccc} /* (22, 12, 17) {real, imag} */,
  {32'h403fb040, 32'h404d0466} /* (22, 12, 16) {real, imag} */,
  {32'h3d236b80, 32'h402686d6} /* (22, 12, 15) {real, imag} */,
  {32'hbf4a2d90, 32'hbf06cc6e} /* (22, 12, 14) {real, imag} */,
  {32'hc018ca4c, 32'hc0614a38} /* (22, 12, 13) {real, imag} */,
  {32'h3fe8a7c9, 32'hbfcff7ba} /* (22, 12, 12) {real, imag} */,
  {32'hc0464d92, 32'h401a4a02} /* (22, 12, 11) {real, imag} */,
  {32'hc01d2a32, 32'h40978284} /* (22, 12, 10) {real, imag} */,
  {32'hc01a75b2, 32'h40a4f43f} /* (22, 12, 9) {real, imag} */,
  {32'h3fc76d1d, 32'hc079f87b} /* (22, 12, 8) {real, imag} */,
  {32'h3f5a68fd, 32'hc06b4cc7} /* (22, 12, 7) {real, imag} */,
  {32'hbf58aed6, 32'hc00d07eb} /* (22, 12, 6) {real, imag} */,
  {32'hbee26cc8, 32'hbfd630b0} /* (22, 12, 5) {real, imag} */,
  {32'h3f9e1353, 32'hbebc6548} /* (22, 12, 4) {real, imag} */,
  {32'h3f03bab4, 32'hc0a79bec} /* (22, 12, 3) {real, imag} */,
  {32'h3f0062d0, 32'hc0042791} /* (22, 12, 2) {real, imag} */,
  {32'hc026c023, 32'h40457244} /* (22, 12, 1) {real, imag} */,
  {32'hbf847d34, 32'h3f47e622} /* (22, 12, 0) {real, imag} */,
  {32'h3ff8bfc5, 32'h3ffd7975} /* (22, 11, 31) {real, imag} */,
  {32'h3e80e9cc, 32'h401dba0c} /* (22, 11, 30) {real, imag} */,
  {32'h3cc8ff00, 32'hbe81c898} /* (22, 11, 29) {real, imag} */,
  {32'hc083deba, 32'h407074f4} /* (22, 11, 28) {real, imag} */,
  {32'hbf5e5838, 32'h402ed0b0} /* (22, 11, 27) {real, imag} */,
  {32'h40c56f36, 32'hbf388be4} /* (22, 11, 26) {real, imag} */,
  {32'h3fd138fc, 32'h3f585d13} /* (22, 11, 25) {real, imag} */,
  {32'h406b0136, 32'hc018cfba} /* (22, 11, 24) {real, imag} */,
  {32'h405c4196, 32'hc0735a16} /* (22, 11, 23) {real, imag} */,
  {32'h40a2fdc4, 32'hbffc1466} /* (22, 11, 22) {real, imag} */,
  {32'h40b12909, 32'hbf063de8} /* (22, 11, 21) {real, imag} */,
  {32'h4099ff54, 32'hc08e95ca} /* (22, 11, 20) {real, imag} */,
  {32'h3feeb80c, 32'hc02e6182} /* (22, 11, 19) {real, imag} */,
  {32'hc00769da, 32'hbf3d2a72} /* (22, 11, 18) {real, imag} */,
  {32'hbeebe674, 32'h40484abc} /* (22, 11, 17) {real, imag} */,
  {32'hbf58fb60, 32'h3f984c7f} /* (22, 11, 16) {real, imag} */,
  {32'h40e4d429, 32'h40887be4} /* (22, 11, 15) {real, imag} */,
  {32'h40e30f26, 32'h4105aad9} /* (22, 11, 14) {real, imag} */,
  {32'hbffb019a, 32'h4006d106} /* (22, 11, 13) {real, imag} */,
  {32'h3fbf48da, 32'hc0c39b87} /* (22, 11, 12) {real, imag} */,
  {32'h3ffb0bc3, 32'hbe7ad448} /* (22, 11, 11) {real, imag} */,
  {32'h3f896f51, 32'h40b0aa81} /* (22, 11, 10) {real, imag} */,
  {32'hc01048de, 32'h40d40712} /* (22, 11, 9) {real, imag} */,
  {32'h3ff99332, 32'h4067d170} /* (22, 11, 8) {real, imag} */,
  {32'h3e949a9e, 32'hbffc94c8} /* (22, 11, 7) {real, imag} */,
  {32'hc028c581, 32'hc0458494} /* (22, 11, 6) {real, imag} */,
  {32'hc0220bf6, 32'hbf6241b4} /* (22, 11, 5) {real, imag} */,
  {32'h4029fd8d, 32'h4084925f} /* (22, 11, 4) {real, imag} */,
  {32'h404da81e, 32'h40c885fc} /* (22, 11, 3) {real, imag} */,
  {32'h3f9b66b8, 32'hbd7ae180} /* (22, 11, 2) {real, imag} */,
  {32'hc03c793b, 32'hc07ec9c9} /* (22, 11, 1) {real, imag} */,
  {32'hbe7cc9e0, 32'hc07fce72} /* (22, 11, 0) {real, imag} */,
  {32'h405b8574, 32'h3f64c0e1} /* (22, 10, 31) {real, imag} */,
  {32'h403cc43e, 32'hc00266b9} /* (22, 10, 30) {real, imag} */,
  {32'hbf1bc7b8, 32'hbff84450} /* (22, 10, 29) {real, imag} */,
  {32'h40176a5a, 32'h3ef0d1c8} /* (22, 10, 28) {real, imag} */,
  {32'hbfd5c1a0, 32'h40295a4f} /* (22, 10, 27) {real, imag} */,
  {32'h40807dd4, 32'h4082a12c} /* (22, 10, 26) {real, imag} */,
  {32'h40d0f83c, 32'h403550c9} /* (22, 10, 25) {real, imag} */,
  {32'h400dd97b, 32'h4030ba36} /* (22, 10, 24) {real, imag} */,
  {32'hbf37420c, 32'hbf1ac7ca} /* (22, 10, 23) {real, imag} */,
  {32'hc0ca9f9a, 32'hbe37d970} /* (22, 10, 22) {real, imag} */,
  {32'hc1026ece, 32'h40b49384} /* (22, 10, 21) {real, imag} */,
  {32'hc027e6da, 32'h4104049f} /* (22, 10, 20) {real, imag} */,
  {32'h404cd90e, 32'h408b2a2b} /* (22, 10, 19) {real, imag} */,
  {32'h408c693a, 32'h3ec3cb00} /* (22, 10, 18) {real, imag} */,
  {32'hbfc6a896, 32'h3f0f7940} /* (22, 10, 17) {real, imag} */,
  {32'h40218e24, 32'h409240e2} /* (22, 10, 16) {real, imag} */,
  {32'h401a0828, 32'h3fd57c9e} /* (22, 10, 15) {real, imag} */,
  {32'h3f9685ef, 32'hc028f44c} /* (22, 10, 14) {real, imag} */,
  {32'h402488b6, 32'h3e418b44} /* (22, 10, 13) {real, imag} */,
  {32'hbfb4b5de, 32'h4092c153} /* (22, 10, 12) {real, imag} */,
  {32'h3fe17db8, 32'hbf54cc46} /* (22, 10, 11) {real, imag} */,
  {32'h40235d0f, 32'h3edefba8} /* (22, 10, 10) {real, imag} */,
  {32'h40825bd8, 32'hc08030a8} /* (22, 10, 9) {real, imag} */,
  {32'h3e1b0100, 32'hc085174c} /* (22, 10, 8) {real, imag} */,
  {32'h3d771b00, 32'h408f3682} /* (22, 10, 7) {real, imag} */,
  {32'h4003b535, 32'h40896aca} /* (22, 10, 6) {real, imag} */,
  {32'h3f4dd82e, 32'h408aadff} /* (22, 10, 5) {real, imag} */,
  {32'hbe6cdb90, 32'h3ff0f7c6} /* (22, 10, 4) {real, imag} */,
  {32'hbf87b230, 32'h3fd5f7c8} /* (22, 10, 3) {real, imag} */,
  {32'hc08a1436, 32'hc03a63fa} /* (22, 10, 2) {real, imag} */,
  {32'hc005d631, 32'hc0271214} /* (22, 10, 1) {real, imag} */,
  {32'hc0308d5f, 32'h40906560} /* (22, 10, 0) {real, imag} */,
  {32'hbecef1a4, 32'hbf88bc28} /* (22, 9, 31) {real, imag} */,
  {32'h40993594, 32'h3fa9c196} /* (22, 9, 30) {real, imag} */,
  {32'hbedc77f0, 32'h4014c1d4} /* (22, 9, 29) {real, imag} */,
  {32'hc0c5b68b, 32'h409ccbab} /* (22, 9, 28) {real, imag} */,
  {32'hc0db6616, 32'h40f03bf5} /* (22, 9, 27) {real, imag} */,
  {32'hc01be1e2, 32'hc08348d2} /* (22, 9, 26) {real, imag} */,
  {32'hc0bfbe48, 32'hc08bbd77} /* (22, 9, 25) {real, imag} */,
  {32'hc0049c48, 32'h41087810} /* (22, 9, 24) {real, imag} */,
  {32'h40316a87, 32'h3fd73ffa} /* (22, 9, 23) {real, imag} */,
  {32'h3f524e62, 32'hc073bd4a} /* (22, 9, 22) {real, imag} */,
  {32'h3f88f21f, 32'h3fa4eb24} /* (22, 9, 21) {real, imag} */,
  {32'hbfef8938, 32'hc0a30830} /* (22, 9, 20) {real, imag} */,
  {32'hc0c468d2, 32'hc098ea78} /* (22, 9, 19) {real, imag} */,
  {32'h3f25e2a0, 32'hc00b1d16} /* (22, 9, 18) {real, imag} */,
  {32'h408de3e0, 32'h40a221b5} /* (22, 9, 17) {real, imag} */,
  {32'h40104b09, 32'h40de9ece} /* (22, 9, 16) {real, imag} */,
  {32'hc0c3ba49, 32'h40a14d6b} /* (22, 9, 15) {real, imag} */,
  {32'hc0ed92c6, 32'h40bfd90c} /* (22, 9, 14) {real, imag} */,
  {32'h3e8c1658, 32'h40bb0763} /* (22, 9, 13) {real, imag} */,
  {32'hbf4d9830, 32'h3f203a44} /* (22, 9, 12) {real, imag} */,
  {32'h4017a053, 32'hbf28c4d8} /* (22, 9, 11) {real, imag} */,
  {32'h3e94df18, 32'h400eb432} /* (22, 9, 10) {real, imag} */,
  {32'hbf904d56, 32'hc0f73adc} /* (22, 9, 9) {real, imag} */,
  {32'h4094dd9a, 32'hc0e35cff} /* (22, 9, 8) {real, imag} */,
  {32'h40092058, 32'h40bdf6a4} /* (22, 9, 7) {real, imag} */,
  {32'h3fcf73ec, 32'h404712a7} /* (22, 9, 6) {real, imag} */,
  {32'h4102291b, 32'h3f90c532} /* (22, 9, 5) {real, imag} */,
  {32'h402bb502, 32'hc0df91ba} /* (22, 9, 4) {real, imag} */,
  {32'h40023b36, 32'hc0bbdb29} /* (22, 9, 3) {real, imag} */,
  {32'h4045ff25, 32'hc09d24e0} /* (22, 9, 2) {real, imag} */,
  {32'hbf31f9da, 32'hbf408328} /* (22, 9, 1) {real, imag} */,
  {32'h40242761, 32'h401426a8} /* (22, 9, 0) {real, imag} */,
  {32'h3fbc36de, 32'hc0363550} /* (22, 8, 31) {real, imag} */,
  {32'h40265748, 32'h3fa5ca14} /* (22, 8, 30) {real, imag} */,
  {32'h401c16ea, 32'hc0844890} /* (22, 8, 29) {real, imag} */,
  {32'hbf009f00, 32'h3fdf7e5c} /* (22, 8, 28) {real, imag} */,
  {32'hbfd2ea94, 32'h40963445} /* (22, 8, 27) {real, imag} */,
  {32'h406bd618, 32'h3f9d7c17} /* (22, 8, 26) {real, imag} */,
  {32'hbf9c3686, 32'hc0828136} /* (22, 8, 25) {real, imag} */,
  {32'hc0d04d02, 32'hbd3fe380} /* (22, 8, 24) {real, imag} */,
  {32'hc1069f3c, 32'hc019ea0f} /* (22, 8, 23) {real, imag} */,
  {32'hc119f26d, 32'h40684636} /* (22, 8, 22) {real, imag} */,
  {32'h3f0ec7d8, 32'hc06e4e1d} /* (22, 8, 21) {real, imag} */,
  {32'h40f5672b, 32'h3d32bd40} /* (22, 8, 20) {real, imag} */,
  {32'h40ad5b3f, 32'hc06caf8c} /* (22, 8, 19) {real, imag} */,
  {32'h408e8a48, 32'hc0e00847} /* (22, 8, 18) {real, imag} */,
  {32'hc0305b86, 32'hc0e11372} /* (22, 8, 17) {real, imag} */,
  {32'hc11373cf, 32'hc089348a} /* (22, 8, 16) {real, imag} */,
  {32'hc1037dc0, 32'hbc9fae80} /* (22, 8, 15) {real, imag} */,
  {32'hbf2af760, 32'h4093a99c} /* (22, 8, 14) {real, imag} */,
  {32'hbebdb846, 32'h3febdcde} /* (22, 8, 13) {real, imag} */,
  {32'hc08a673d, 32'hc025369b} /* (22, 8, 12) {real, imag} */,
  {32'hc07aa8d2, 32'h3e552080} /* (22, 8, 11) {real, imag} */,
  {32'hbf29ac08, 32'hc05779d0} /* (22, 8, 10) {real, imag} */,
  {32'h410ff557, 32'h4129fd86} /* (22, 8, 9) {real, imag} */,
  {32'h416e483e, 32'h40f8402e} /* (22, 8, 8) {real, imag} */,
  {32'h4131c190, 32'h4002597e} /* (22, 8, 7) {real, imag} */,
  {32'hc0e33b6b, 32'hc01eb30a} /* (22, 8, 6) {real, imag} */,
  {32'hc10f3c72, 32'h3a851400} /* (22, 8, 5) {real, imag} */,
  {32'hbea07308, 32'hc043b399} /* (22, 8, 4) {real, imag} */,
  {32'h3fcc60e2, 32'h408b61ca} /* (22, 8, 3) {real, imag} */,
  {32'h40ea6fb2, 32'hbff3f8b0} /* (22, 8, 2) {real, imag} */,
  {32'h3effcd10, 32'hbfcbad4c} /* (22, 8, 1) {real, imag} */,
  {32'hc02877f4, 32'hc019eb9c} /* (22, 8, 0) {real, imag} */,
  {32'h3f3561f6, 32'hbfa31fae} /* (22, 7, 31) {real, imag} */,
  {32'hc03f8040, 32'hc0d0a01d} /* (22, 7, 30) {real, imag} */,
  {32'hc129b641, 32'hc1121deb} /* (22, 7, 29) {real, imag} */,
  {32'hc0823e1d, 32'hbf792570} /* (22, 7, 28) {real, imag} */,
  {32'h405c3216, 32'hc0f965d7} /* (22, 7, 27) {real, imag} */,
  {32'h40c4811f, 32'hc10bde66} /* (22, 7, 26) {real, imag} */,
  {32'h40cc8980, 32'hc03ec611} /* (22, 7, 25) {real, imag} */,
  {32'h40070b1e, 32'hc07454ae} /* (22, 7, 24) {real, imag} */,
  {32'h3f349e02, 32'hc093d0aa} /* (22, 7, 23) {real, imag} */,
  {32'hc0ba6e6d, 32'h40a56800} /* (22, 7, 22) {real, imag} */,
  {32'h40d88ab2, 32'h3f9d5e22} /* (22, 7, 21) {real, imag} */,
  {32'h410824a9, 32'hc0894cab} /* (22, 7, 20) {real, imag} */,
  {32'h405bc68e, 32'hc0b061c0} /* (22, 7, 19) {real, imag} */,
  {32'hc08e0cbc, 32'hc0f7fb3d} /* (22, 7, 18) {real, imag} */,
  {32'hc023222a, 32'hc089c27b} /* (22, 7, 17) {real, imag} */,
  {32'hc04ce4eb, 32'hbe333c00} /* (22, 7, 16) {real, imag} */,
  {32'hc0cad170, 32'h3e29f838} /* (22, 7, 15) {real, imag} */,
  {32'h405255a7, 32'hc0ba80d0} /* (22, 7, 14) {real, imag} */,
  {32'hbf105e14, 32'h3fb929a4} /* (22, 7, 13) {real, imag} */,
  {32'hc13cd68a, 32'h4115e1ec} /* (22, 7, 12) {real, imag} */,
  {32'hc100b846, 32'h411d4782} /* (22, 7, 11) {real, imag} */,
  {32'hc0c7a33c, 32'hc098b283} /* (22, 7, 10) {real, imag} */,
  {32'hc0e484cc, 32'hc161e458} /* (22, 7, 9) {real, imag} */,
  {32'hbfd83240, 32'hc0ac9075} /* (22, 7, 8) {real, imag} */,
  {32'h400429c2, 32'h4068abec} /* (22, 7, 7) {real, imag} */,
  {32'h3eb26dec, 32'h40e5e058} /* (22, 7, 6) {real, imag} */,
  {32'hc0948442, 32'hbffaa932} /* (22, 7, 5) {real, imag} */,
  {32'hbfe215d4, 32'hbf94d77a} /* (22, 7, 4) {real, imag} */,
  {32'hbe1ad220, 32'h40a52bc1} /* (22, 7, 3) {real, imag} */,
  {32'h404227d2, 32'h41295b8f} /* (22, 7, 2) {real, imag} */,
  {32'h4109f535, 32'h4128cdd2} /* (22, 7, 1) {real, imag} */,
  {32'h3f3fd8dc, 32'h408023e0} /* (22, 7, 0) {real, imag} */,
  {32'hc05c88cc, 32'h3e834d6c} /* (22, 6, 31) {real, imag} */,
  {32'hc10bab71, 32'h40b8b422} /* (22, 6, 30) {real, imag} */,
  {32'h40e48e1f, 32'h4085735a} /* (22, 6, 29) {real, imag} */,
  {32'h41397a76, 32'h40d1ee84} /* (22, 6, 28) {real, imag} */,
  {32'h40b5603c, 32'h41307510} /* (22, 6, 27) {real, imag} */,
  {32'hbfb46ccb, 32'h40f0dcc7} /* (22, 6, 26) {real, imag} */,
  {32'hc10c4124, 32'h3fdd485d} /* (22, 6, 25) {real, imag} */,
  {32'hbf5d7db0, 32'hbfa09434} /* (22, 6, 24) {real, imag} */,
  {32'h410ddd25, 32'hc10b3f92} /* (22, 6, 23) {real, imag} */,
  {32'h4127661d, 32'hc0db33fe} /* (22, 6, 22) {real, imag} */,
  {32'h404330ca, 32'hc0578ab5} /* (22, 6, 21) {real, imag} */,
  {32'h3fd6b482, 32'hbf85ddc4} /* (22, 6, 20) {real, imag} */,
  {32'hbfd893c0, 32'h4050fc4e} /* (22, 6, 19) {real, imag} */,
  {32'hc11ffcb7, 32'h4181042d} /* (22, 6, 18) {real, imag} */,
  {32'hc05dd3e2, 32'h41063d89} /* (22, 6, 17) {real, imag} */,
  {32'hc030a7e1, 32'hbf9dcf9c} /* (22, 6, 16) {real, imag} */,
  {32'h3f15a710, 32'hc0909f5a} /* (22, 6, 15) {real, imag} */,
  {32'h3fac1d3a, 32'h3fd691f8} /* (22, 6, 14) {real, imag} */,
  {32'h4050af1a, 32'h411962e8} /* (22, 6, 13) {real, imag} */,
  {32'h4055dbd8, 32'h40259cf5} /* (22, 6, 12) {real, imag} */,
  {32'h40ca3a04, 32'h3fc73a3d} /* (22, 6, 11) {real, imag} */,
  {32'h415e592e, 32'hbf7e15dc} /* (22, 6, 10) {real, imag} */,
  {32'h40b3f9de, 32'h3fbe690d} /* (22, 6, 9) {real, imag} */,
  {32'h40216d28, 32'h40a9fd9a} /* (22, 6, 8) {real, imag} */,
  {32'hc0825f5d, 32'h3d4f4800} /* (22, 6, 7) {real, imag} */,
  {32'hc0d3eac8, 32'hc00c5045} /* (22, 6, 6) {real, imag} */,
  {32'h40ede778, 32'h40571c4c} /* (22, 6, 5) {real, imag} */,
  {32'h4004f3d6, 32'hc0829893} /* (22, 6, 4) {real, imag} */,
  {32'h40bf9cea, 32'hc05dda62} /* (22, 6, 3) {real, imag} */,
  {32'h40d5eb78, 32'hc00d17d8} /* (22, 6, 2) {real, imag} */,
  {32'hc003bb2a, 32'h3ee4b380} /* (22, 6, 1) {real, imag} */,
  {32'h407895a5, 32'h400a4224} /* (22, 6, 0) {real, imag} */,
  {32'hbf70c65a, 32'h4051fadc} /* (22, 5, 31) {real, imag} */,
  {32'h40233be8, 32'h3fb997fc} /* (22, 5, 30) {real, imag} */,
  {32'hc055d092, 32'h4034fa13} /* (22, 5, 29) {real, imag} */,
  {32'hc00ce30a, 32'hc1051014} /* (22, 5, 28) {real, imag} */,
  {32'h4112de89, 32'hc0e1f864} /* (22, 5, 27) {real, imag} */,
  {32'h40f7ae66, 32'h4036ee87} /* (22, 5, 26) {real, imag} */,
  {32'h40c317a6, 32'h4105c489} /* (22, 5, 25) {real, imag} */,
  {32'h3f9ede84, 32'h3f5b1fa8} /* (22, 5, 24) {real, imag} */,
  {32'h3fa70c70, 32'hc0b2e690} /* (22, 5, 23) {real, imag} */,
  {32'hc0177c22, 32'hc0089164} /* (22, 5, 22) {real, imag} */,
  {32'h4128680f, 32'hbed29cd0} /* (22, 5, 21) {real, imag} */,
  {32'h41513114, 32'hbd03faa0} /* (22, 5, 20) {real, imag} */,
  {32'h409adc28, 32'h40bae45a} /* (22, 5, 19) {real, imag} */,
  {32'hbfefe068, 32'h40e9b0fd} /* (22, 5, 18) {real, imag} */,
  {32'hbfea0d48, 32'h4084124e} /* (22, 5, 17) {real, imag} */,
  {32'hc0ab611a, 32'h401e30ba} /* (22, 5, 16) {real, imag} */,
  {32'h4066958c, 32'hc077315d} /* (22, 5, 15) {real, imag} */,
  {32'h41598c54, 32'hc14d1adf} /* (22, 5, 14) {real, imag} */,
  {32'h400d8319, 32'hc1075df5} /* (22, 5, 13) {real, imag} */,
  {32'hc0e0a534, 32'h3de041b0} /* (22, 5, 12) {real, imag} */,
  {32'hc023210e, 32'h406101aa} /* (22, 5, 11) {real, imag} */,
  {32'hc0817389, 32'h40b43b67} /* (22, 5, 10) {real, imag} */,
  {32'hbe1a0fb0, 32'h4120ad78} /* (22, 5, 9) {real, imag} */,
  {32'hc0559d55, 32'hbf5cebb4} /* (22, 5, 8) {real, imag} */,
  {32'h409307c4, 32'hc13107d8} /* (22, 5, 7) {real, imag} */,
  {32'h406220e0, 32'hc1274138} /* (22, 5, 6) {real, imag} */,
  {32'h404ae150, 32'hc1764cfa} /* (22, 5, 5) {real, imag} */,
  {32'h3f92ca5e, 32'hc118e115} /* (22, 5, 4) {real, imag} */,
  {32'h40442152, 32'hbfc9d79e} /* (22, 5, 3) {real, imag} */,
  {32'hc09d0087, 32'hc050dd6b} /* (22, 5, 2) {real, imag} */,
  {32'hc045621a, 32'hc0149981} /* (22, 5, 1) {real, imag} */,
  {32'hbe770710, 32'h3fd5fbe2} /* (22, 5, 0) {real, imag} */,
  {32'hbfd61dd8, 32'hbe104f30} /* (22, 4, 31) {real, imag} */,
  {32'hbfa5c8fa, 32'h40852617} /* (22, 4, 30) {real, imag} */,
  {32'h409c5284, 32'h412d2e10} /* (22, 4, 29) {real, imag} */,
  {32'h40849867, 32'h4001c394} /* (22, 4, 28) {real, imag} */,
  {32'hbfd6f90f, 32'hc1513572} /* (22, 4, 27) {real, imag} */,
  {32'hc00746b4, 32'hc0de5261} /* (22, 4, 26) {real, imag} */,
  {32'hc0457342, 32'hc0081d5c} /* (22, 4, 25) {real, imag} */,
  {32'h3f697924, 32'hc11f0e5a} /* (22, 4, 24) {real, imag} */,
  {32'h408299df, 32'hc082f0a4} /* (22, 4, 23) {real, imag} */,
  {32'hc1287b5a, 32'h40d5fe37} /* (22, 4, 22) {real, imag} */,
  {32'hc08dee50, 32'hc052cfac} /* (22, 4, 21) {real, imag} */,
  {32'h40a0546f, 32'h3f9e9c98} /* (22, 4, 20) {real, imag} */,
  {32'hc0bdaf02, 32'h3fe2e4f6} /* (22, 4, 19) {real, imag} */,
  {32'hc115cd5e, 32'hc0e8588d} /* (22, 4, 18) {real, imag} */,
  {32'hc0dd8cd9, 32'hc071820e} /* (22, 4, 17) {real, imag} */,
  {32'hc175f102, 32'hc01e0c98} /* (22, 4, 16) {real, imag} */,
  {32'h409aa0ac, 32'h3f46e12c} /* (22, 4, 15) {real, imag} */,
  {32'h4025125a, 32'h4153f25c} /* (22, 4, 14) {real, imag} */,
  {32'h41065f5c, 32'h4150cde8} /* (22, 4, 13) {real, imag} */,
  {32'h4106b818, 32'h4113de07} /* (22, 4, 12) {real, imag} */,
  {32'hc106e1c7, 32'hbf9d4020} /* (22, 4, 11) {real, imag} */,
  {32'hbf27620c, 32'hc1689119} /* (22, 4, 10) {real, imag} */,
  {32'h4044f23e, 32'hc18403ee} /* (22, 4, 9) {real, imag} */,
  {32'hc060d008, 32'hc0e44ae6} /* (22, 4, 8) {real, imag} */,
  {32'hc0be0993, 32'h3da71b00} /* (22, 4, 7) {real, imag} */,
  {32'h3faea8ef, 32'h3fb6bfe8} /* (22, 4, 6) {real, imag} */,
  {32'h413b9612, 32'hc11fe116} /* (22, 4, 5) {real, imag} */,
  {32'h4195d70e, 32'hc0c29046} /* (22, 4, 4) {real, imag} */,
  {32'h40e444e2, 32'hbf201f98} /* (22, 4, 3) {real, imag} */,
  {32'hc03eb978, 32'hbf778673} /* (22, 4, 2) {real, imag} */,
  {32'hc0ee1eac, 32'h404a8e4f} /* (22, 4, 1) {real, imag} */,
  {32'hc0f2debd, 32'hbfbcc3d2} /* (22, 4, 0) {real, imag} */,
  {32'hc10d59ec, 32'h4143bb94} /* (22, 3, 31) {real, imag} */,
  {32'hc191dbb0, 32'h41bf1cf4} /* (22, 3, 30) {real, imag} */,
  {32'hc1383459, 32'h41357bc2} /* (22, 3, 29) {real, imag} */,
  {32'hc000c8d3, 32'h3f978d10} /* (22, 3, 28) {real, imag} */,
  {32'h408e7999, 32'hc0250a4a} /* (22, 3, 27) {real, imag} */,
  {32'h3eacc238, 32'hbffa0246} /* (22, 3, 26) {real, imag} */,
  {32'hc100a744, 32'hc0bed30b} /* (22, 3, 25) {real, imag} */,
  {32'hc0114c4d, 32'hbf2d04fd} /* (22, 3, 24) {real, imag} */,
  {32'hc0e381f6, 32'h4051ed03} /* (22, 3, 23) {real, imag} */,
  {32'h40e24a8a, 32'hbeed0674} /* (22, 3, 22) {real, imag} */,
  {32'h40a4616f, 32'hc1192f85} /* (22, 3, 21) {real, imag} */,
  {32'hbf2e1f30, 32'hbfec83b6} /* (22, 3, 20) {real, imag} */,
  {32'h3fbd638b, 32'h4050fe22} /* (22, 3, 19) {real, imag} */,
  {32'h40f76d1d, 32'h40dffdce} /* (22, 3, 18) {real, imag} */,
  {32'hbfbb2ab0, 32'h41023a5f} /* (22, 3, 17) {real, imag} */,
  {32'h40a99281, 32'h3ddea820} /* (22, 3, 16) {real, imag} */,
  {32'h40fd8d35, 32'h3e1c33c0} /* (22, 3, 15) {real, imag} */,
  {32'hbd9e1e20, 32'h41051956} /* (22, 3, 14) {real, imag} */,
  {32'hc0510f26, 32'h40116748} /* (22, 3, 13) {real, imag} */,
  {32'hc0c8a60f, 32'hc018fca0} /* (22, 3, 12) {real, imag} */,
  {32'h40ab1801, 32'hc0468754} /* (22, 3, 11) {real, imag} */,
  {32'hc0c1013f, 32'hc0109dde} /* (22, 3, 10) {real, imag} */,
  {32'hc0e8257e, 32'hbf63c440} /* (22, 3, 9) {real, imag} */,
  {32'h4120645c, 32'h3ee9f250} /* (22, 3, 8) {real, imag} */,
  {32'h40f80b94, 32'h4099913b} /* (22, 3, 7) {real, imag} */,
  {32'hc039da1a, 32'h409e94a6} /* (22, 3, 6) {real, imag} */,
  {32'hc134637a, 32'h3f70e80c} /* (22, 3, 5) {real, imag} */,
  {32'hc0f03879, 32'h410c59d6} /* (22, 3, 4) {real, imag} */,
  {32'hc0e1b805, 32'h41141bf3} /* (22, 3, 3) {real, imag} */,
  {32'h404d7d6c, 32'h4123220c} /* (22, 3, 2) {real, imag} */,
  {32'hc12cbdda, 32'h40e03891} /* (22, 3, 1) {real, imag} */,
  {32'hc144d65b, 32'h4006d46b} /* (22, 3, 0) {real, imag} */,
  {32'h410a5272, 32'h40a585db} /* (22, 2, 31) {real, imag} */,
  {32'h41bc313b, 32'h418b58aa} /* (22, 2, 30) {real, imag} */,
  {32'h404f562a, 32'h4183f0bf} /* (22, 2, 29) {real, imag} */,
  {32'h4061a2a2, 32'h4114a39e} /* (22, 2, 28) {real, imag} */,
  {32'hc0658aa4, 32'h3fcc5ee8} /* (22, 2, 27) {real, imag} */,
  {32'hc0cfd1b2, 32'h4040f922} /* (22, 2, 26) {real, imag} */,
  {32'hc00c56d6, 32'hc0d8f752} /* (22, 2, 25) {real, imag} */,
  {32'hc114c834, 32'hc1041ea7} /* (22, 2, 24) {real, imag} */,
  {32'h415b9093, 32'hbf1247c2} /* (22, 2, 23) {real, imag} */,
  {32'h41c1c920, 32'h409ca330} /* (22, 2, 22) {real, imag} */,
  {32'h412c54a7, 32'h401f4e6e} /* (22, 2, 21) {real, imag} */,
  {32'hc0eb559e, 32'hc04a5b1c} /* (22, 2, 20) {real, imag} */,
  {32'hc150ff98, 32'h405074bd} /* (22, 2, 19) {real, imag} */,
  {32'hc0e3665e, 32'h40623c5c} /* (22, 2, 18) {real, imag} */,
  {32'hbfe9f790, 32'hbfff862c} /* (22, 2, 17) {real, imag} */,
  {32'hc05e310c, 32'hc0a1c79d} /* (22, 2, 16) {real, imag} */,
  {32'hc0cd3126, 32'hc0677950} /* (22, 2, 15) {real, imag} */,
  {32'h402d9cac, 32'hbf006a80} /* (22, 2, 14) {real, imag} */,
  {32'h404dace0, 32'h3f92965a} /* (22, 2, 13) {real, imag} */,
  {32'h412eba62, 32'h404b20ac} /* (22, 2, 12) {real, imag} */,
  {32'h40272429, 32'h412a283b} /* (22, 2, 11) {real, imag} */,
  {32'h40ee0e55, 32'h416ef9d1} /* (22, 2, 10) {real, imag} */,
  {32'h419a0bed, 32'h410d2cb2} /* (22, 2, 9) {real, imag} */,
  {32'h418b4297, 32'hc115a29f} /* (22, 2, 8) {real, imag} */,
  {32'h41887059, 32'hc130fe35} /* (22, 2, 7) {real, imag} */,
  {32'h41ad3212, 32'hbfde1cf6} /* (22, 2, 6) {real, imag} */,
  {32'h4197bc1b, 32'hbf832530} /* (22, 2, 5) {real, imag} */,
  {32'h3f9b5660, 32'hc0b843d0} /* (22, 2, 4) {real, imag} */,
  {32'h3fdb5d90, 32'hc0015aba} /* (22, 2, 3) {real, imag} */,
  {32'h3cf47b00, 32'hc06fce08} /* (22, 2, 2) {real, imag} */,
  {32'h3f2708a0, 32'hc0d62e00} /* (22, 2, 1) {real, imag} */,
  {32'hbf19b18a, 32'hc04672f2} /* (22, 2, 0) {real, imag} */,
  {32'hc096c503, 32'hc0ff6152} /* (22, 1, 31) {real, imag} */,
  {32'h3e3de800, 32'hc1a252ea} /* (22, 1, 30) {real, imag} */,
  {32'h3e7e1d00, 32'hc1730991} /* (22, 1, 29) {real, imag} */,
  {32'hc06df246, 32'hc0ecede2} /* (22, 1, 28) {real, imag} */,
  {32'hc0b52976, 32'hbf1005fc} /* (22, 1, 27) {real, imag} */,
  {32'hc0c5fe48, 32'hbedf74a0} /* (22, 1, 26) {real, imag} */,
  {32'hc0ef563c, 32'hc0b34d77} /* (22, 1, 25) {real, imag} */,
  {32'hc18174c5, 32'hc1323bb1} /* (22, 1, 24) {real, imag} */,
  {32'hc114ba2a, 32'hc1c43118} /* (22, 1, 23) {real, imag} */,
  {32'hbc8fef60, 32'hc148f7f6} /* (22, 1, 22) {real, imag} */,
  {32'h4130c484, 32'hc06c2597} /* (22, 1, 21) {real, imag} */,
  {32'h419f9453, 32'h40c342e8} /* (22, 1, 20) {real, imag} */,
  {32'h41600d40, 32'hbf6c1538} /* (22, 1, 19) {real, imag} */,
  {32'h40b8d497, 32'hc123737e} /* (22, 1, 18) {real, imag} */,
  {32'h3f996c18, 32'h3fe1c7c8} /* (22, 1, 17) {real, imag} */,
  {32'hbeee9ed2, 32'h415a247e} /* (22, 1, 16) {real, imag} */,
  {32'h4093e6ee, 32'h412e274e} /* (22, 1, 15) {real, imag} */,
  {32'h40ad7c0e, 32'h40f88c43} /* (22, 1, 14) {real, imag} */,
  {32'h41625636, 32'h41635d4e} /* (22, 1, 13) {real, imag} */,
  {32'h4157d830, 32'h40f1dfe6} /* (22, 1, 12) {real, imag} */,
  {32'h403b3358, 32'hc104998b} /* (22, 1, 11) {real, imag} */,
  {32'h4122d8fe, 32'hc15ff886} /* (22, 1, 10) {real, imag} */,
  {32'h40decb58, 32'hc1ac1cba} /* (22, 1, 9) {real, imag} */,
  {32'h40812d76, 32'hc187b11b} /* (22, 1, 8) {real, imag} */,
  {32'hc034152a, 32'h405756a2} /* (22, 1, 7) {real, imag} */,
  {32'h40c1a725, 32'h3dc39500} /* (22, 1, 6) {real, imag} */,
  {32'hc065c524, 32'hc144cc22} /* (22, 1, 5) {real, imag} */,
  {32'hc13ab9ee, 32'hc1a366b1} /* (22, 1, 4) {real, imag} */,
  {32'hc0e79b0d, 32'hc10669eb} /* (22, 1, 3) {real, imag} */,
  {32'h40612136, 32'h4087107e} /* (22, 1, 2) {real, imag} */,
  {32'h415c4818, 32'h3e5ce860} /* (22, 1, 1) {real, imag} */,
  {32'h40b074ae, 32'hc01e0980} /* (22, 1, 0) {real, imag} */,
  {32'h40b1f3aa, 32'hbf792f0e} /* (22, 0, 31) {real, imag} */,
  {32'h3f9dbf1d, 32'h3da3fd00} /* (22, 0, 30) {real, imag} */,
  {32'hc11437e6, 32'hbf2e96a8} /* (22, 0, 29) {real, imag} */,
  {32'hc1a1e3b0, 32'hc10808a1} /* (22, 0, 28) {real, imag} */,
  {32'hc13ccad3, 32'h40e5ced3} /* (22, 0, 27) {real, imag} */,
  {32'h3fc8183c, 32'h4103867c} /* (22, 0, 26) {real, imag} */,
  {32'h405d4733, 32'h40013df8} /* (22, 0, 25) {real, imag} */,
  {32'h3f7ea312, 32'hc0fffddc} /* (22, 0, 24) {real, imag} */,
  {32'hc18bd9c2, 32'hc12115a7} /* (22, 0, 23) {real, imag} */,
  {32'hc13d46f4, 32'hc0e6863f} /* (22, 0, 22) {real, imag} */,
  {32'hbfba0551, 32'h40e94e65} /* (22, 0, 21) {real, imag} */,
  {32'hc13195da, 32'hbfb68874} /* (22, 0, 20) {real, imag} */,
  {32'h40039e22, 32'hc0e4b31e} /* (22, 0, 19) {real, imag} */,
  {32'h414f35f4, 32'hc13222c2} /* (22, 0, 18) {real, imag} */,
  {32'h4168f57e, 32'hbfc897a4} /* (22, 0, 17) {real, imag} */,
  {32'h3f315442, 32'h40a7b30a} /* (22, 0, 16) {real, imag} */,
  {32'h40a79cda, 32'h416da39a} /* (22, 0, 15) {real, imag} */,
  {32'h41a99bae, 32'h40c6fb5b} /* (22, 0, 14) {real, imag} */,
  {32'h4014a2f0, 32'hc0c686c8} /* (22, 0, 13) {real, imag} */,
  {32'hc0d37f5c, 32'hc07b2523} /* (22, 0, 12) {real, imag} */,
  {32'hc0bdb3e8, 32'h405f375c} /* (22, 0, 11) {real, imag} */,
  {32'hc09e03e4, 32'h40373aa8} /* (22, 0, 10) {real, imag} */,
  {32'hc10caa93, 32'h41663c62} /* (22, 0, 9) {real, imag} */,
  {32'h400cab37, 32'hbfdf1674} /* (22, 0, 8) {real, imag} */,
  {32'h4162c4c4, 32'hc0acbcea} /* (22, 0, 7) {real, imag} */,
  {32'h418664a8, 32'hbfab202e} /* (22, 0, 6) {real, imag} */,
  {32'h4003cf24, 32'hc05d5521} /* (22, 0, 5) {real, imag} */,
  {32'h4102ea60, 32'hc123a64c} /* (22, 0, 4) {real, imag} */,
  {32'hbf225487, 32'h3fbb9071} /* (22, 0, 3) {real, imag} */,
  {32'hc188f2e5, 32'h4186f244} /* (22, 0, 2) {real, imag} */,
  {32'hc1b5ffcc, 32'h41be9762} /* (22, 0, 1) {real, imag} */,
  {32'hc01e5004, 32'h413b1128} /* (22, 0, 0) {real, imag} */,
  {32'h40b6e812, 32'h3f9df060} /* (21, 31, 31) {real, imag} */,
  {32'h411a9073, 32'h40cd0f2a} /* (21, 31, 30) {real, imag} */,
  {32'h40d7956e, 32'h416711bb} /* (21, 31, 29) {real, imag} */,
  {32'h4154072c, 32'h4183d9cb} /* (21, 31, 28) {real, imag} */,
  {32'h41970e14, 32'h40e00684} /* (21, 31, 27) {real, imag} */,
  {32'h4141a288, 32'h3f050d8e} /* (21, 31, 26) {real, imag} */,
  {32'h419c184c, 32'h40f46ca8} /* (21, 31, 25) {real, imag} */,
  {32'h41857f9e, 32'h404fbb10} /* (21, 31, 24) {real, imag} */,
  {32'h41c32d49, 32'hc080032a} /* (21, 31, 23) {real, imag} */,
  {32'h41ae8eb4, 32'h40953814} /* (21, 31, 22) {real, imag} */,
  {32'h410d36ec, 32'h40f4c2f4} /* (21, 31, 21) {real, imag} */,
  {32'hc127ae8e, 32'h4196c256} /* (21, 31, 20) {real, imag} */,
  {32'hc08cd4a0, 32'h409b67c2} /* (21, 31, 19) {real, imag} */,
  {32'hc1188da8, 32'h410be21a} /* (21, 31, 18) {real, imag} */,
  {32'hc11049c5, 32'h40e91131} /* (21, 31, 17) {real, imag} */,
  {32'hc0ed3556, 32'hc028e2a2} /* (21, 31, 16) {real, imag} */,
  {32'hc101344c, 32'hc060102b} /* (21, 31, 15) {real, imag} */,
  {32'hc17df5d2, 32'hc08dd4c2} /* (21, 31, 14) {real, imag} */,
  {32'hc1cbe031, 32'hc0b28744} /* (21, 31, 13) {real, imag} */,
  {32'hc1124ea6, 32'hc12fce66} /* (21, 31, 12) {real, imag} */,
  {32'h40ed3366, 32'hc150ab38} /* (21, 31, 11) {real, imag} */,
  {32'h41509600, 32'hc08649ba} /* (21, 31, 10) {real, imag} */,
  {32'h412cb9f2, 32'h3fbf6960} /* (21, 31, 9) {real, imag} */,
  {32'h414d5a0a, 32'hc191d662} /* (21, 31, 8) {real, imag} */,
  {32'h416a98a7, 32'hc1834154} /* (21, 31, 7) {real, imag} */,
  {32'h4098e049, 32'hc0fa78fc} /* (21, 31, 6) {real, imag} */,
  {32'hbe7ca180, 32'h40d3f0b8} /* (21, 31, 5) {real, imag} */,
  {32'h41141d4f, 32'h418648b4} /* (21, 31, 4) {real, imag} */,
  {32'h41999dee, 32'h4048627c} /* (21, 31, 3) {real, imag} */,
  {32'h419e6828, 32'hc0b01672} /* (21, 31, 2) {real, imag} */,
  {32'h3f8e2f90, 32'hc0e1f811} /* (21, 31, 1) {real, imag} */,
  {32'h40823d6a, 32'h3fdb411c} /* (21, 31, 0) {real, imag} */,
  {32'hc1214fc8, 32'hc02a644c} /* (21, 30, 31) {real, imag} */,
  {32'hc140f890, 32'h3feefd78} /* (21, 30, 30) {real, imag} */,
  {32'hc16ec308, 32'hc013c624} /* (21, 30, 29) {real, imag} */,
  {32'hc128924e, 32'hc154b099} /* (21, 30, 28) {real, imag} */,
  {32'hc1182ecc, 32'hc15d2a50} /* (21, 30, 27) {real, imag} */,
  {32'hc132e0b6, 32'h409a658b} /* (21, 30, 26) {real, imag} */,
  {32'hc1aeceed, 32'h40c6c997} /* (21, 30, 25) {real, imag} */,
  {32'hc119ad65, 32'hc0973c42} /* (21, 30, 24) {real, imag} */,
  {32'hc0e02717, 32'h408e6e7b} /* (21, 30, 23) {real, imag} */,
  {32'hc07c8f40, 32'h405e21b1} /* (21, 30, 22) {real, imag} */,
  {32'hc0ca60a3, 32'h411ef3fd} /* (21, 30, 21) {real, imag} */,
  {32'h40d798b9, 32'h410504bf} /* (21, 30, 20) {real, imag} */,
  {32'h41509cb1, 32'h40926a30} /* (21, 30, 19) {real, imag} */,
  {32'h4138ff74, 32'h4161cb0c} /* (21, 30, 18) {real, imag} */,
  {32'h41147905, 32'h4193e6ba} /* (21, 30, 17) {real, imag} */,
  {32'h40cc906c, 32'h414bba2a} /* (21, 30, 16) {real, imag} */,
  {32'h413fee62, 32'h40900e28} /* (21, 30, 15) {real, imag} */,
  {32'h40cca2f4, 32'hc0d2c95c} /* (21, 30, 14) {real, imag} */,
  {32'hc09a5b23, 32'hc040cdac} /* (21, 30, 13) {real, imag} */,
  {32'hbe8a3460, 32'hc043011e} /* (21, 30, 12) {real, imag} */,
  {32'h415b96fe, 32'hc00a9438} /* (21, 30, 11) {real, imag} */,
  {32'hc12b416a, 32'hc0e292ec} /* (21, 30, 10) {real, imag} */,
  {32'hc19bed1e, 32'hc1933092} /* (21, 30, 9) {real, imag} */,
  {32'hc0a5d19f, 32'hc08074c8} /* (21, 30, 8) {real, imag} */,
  {32'hbfbabc88, 32'hc05ae6b0} /* (21, 30, 7) {real, imag} */,
  {32'hc0045c3e, 32'hc18e0739} /* (21, 30, 6) {real, imag} */,
  {32'hbfb91ec6, 32'hc0bcf517} /* (21, 30, 5) {real, imag} */,
  {32'hc12238e6, 32'h408e8657} /* (21, 30, 4) {real, imag} */,
  {32'hbec7c1c8, 32'h3f889cac} /* (21, 30, 3) {real, imag} */,
  {32'h3f4af758, 32'h4050a424} /* (21, 30, 2) {real, imag} */,
  {32'h3f075b38, 32'h407fbe64} /* (21, 30, 1) {real, imag} */,
  {32'hc09cc3e8, 32'hc0819474} /* (21, 30, 0) {real, imag} */,
  {32'h40f843d0, 32'h3fbea1f4} /* (21, 29, 31) {real, imag} */,
  {32'h3feef124, 32'hc1929c02} /* (21, 29, 30) {real, imag} */,
  {32'hbfbb0ac0, 32'hc1990817} /* (21, 29, 29) {real, imag} */,
  {32'h40ba1dfb, 32'hc141b263} /* (21, 29, 28) {real, imag} */,
  {32'h408ae664, 32'hc11f660e} /* (21, 29, 27) {real, imag} */,
  {32'h40315488, 32'h3f6a11b0} /* (21, 29, 26) {real, imag} */,
  {32'h4126c714, 32'h4029270a} /* (21, 29, 25) {real, imag} */,
  {32'h4105c153, 32'hc0f7590e} /* (21, 29, 24) {real, imag} */,
  {32'h410b1286, 32'hc10cf954} /* (21, 29, 23) {real, imag} */,
  {32'h40dda90e, 32'hbf0a4c80} /* (21, 29, 22) {real, imag} */,
  {32'hc08434f1, 32'hc0d2343b} /* (21, 29, 21) {real, imag} */,
  {32'hc1407536, 32'h40d37ed9} /* (21, 29, 20) {real, imag} */,
  {32'hc11a68b2, 32'h40ad0236} /* (21, 29, 19) {real, imag} */,
  {32'h3f8b52bc, 32'h40b7fb58} /* (21, 29, 18) {real, imag} */,
  {32'h4033f761, 32'h40e53efd} /* (21, 29, 17) {real, imag} */,
  {32'hc0ee6ab9, 32'hc04ffa8c} /* (21, 29, 16) {real, imag} */,
  {32'h3f68a41c, 32'h40a0818b} /* (21, 29, 15) {real, imag} */,
  {32'h4108b4a3, 32'h416a8f3d} /* (21, 29, 14) {real, imag} */,
  {32'h40c1d396, 32'h4139bf0d} /* (21, 29, 13) {real, imag} */,
  {32'h411ea00f, 32'h400d9e09} /* (21, 29, 12) {real, imag} */,
  {32'h419000ab, 32'hc094bc3b} /* (21, 29, 11) {real, imag} */,
  {32'h3f837f76, 32'hc0935aed} /* (21, 29, 10) {real, imag} */,
  {32'hc00a9db0, 32'hc0186831} /* (21, 29, 9) {real, imag} */,
  {32'h40cd42cd, 32'hc0a2f85a} /* (21, 29, 8) {real, imag} */,
  {32'h417a61d2, 32'hc0a1d9d6} /* (21, 29, 7) {real, imag} */,
  {32'h40881659, 32'hc0ff5c6d} /* (21, 29, 6) {real, imag} */,
  {32'h40082333, 32'hc080d552} /* (21, 29, 5) {real, imag} */,
  {32'h40452d9f, 32'h40b8c7b5} /* (21, 29, 4) {real, imag} */,
  {32'h40a5ee2d, 32'h3f6810b4} /* (21, 29, 3) {real, imag} */,
  {32'hc03c204a, 32'h408a3f3d} /* (21, 29, 2) {real, imag} */,
  {32'hc0bf6505, 32'h401dd257} /* (21, 29, 1) {real, imag} */,
  {32'hc04adb46, 32'h3fb1d90e} /* (21, 29, 0) {real, imag} */,
  {32'hbf407530, 32'h40871721} /* (21, 28, 31) {real, imag} */,
  {32'h40c93162, 32'h41019bcc} /* (21, 28, 30) {real, imag} */,
  {32'h40fdfefd, 32'h4096dfe5} /* (21, 28, 29) {real, imag} */,
  {32'h3f9de1d3, 32'h410c7090} /* (21, 28, 28) {real, imag} */,
  {32'hc0656a5f, 32'hc040bbc0} /* (21, 28, 27) {real, imag} */,
  {32'hc1169fee, 32'hc1524a57} /* (21, 28, 26) {real, imag} */,
  {32'h3ad44400, 32'hbeabbf40} /* (21, 28, 25) {real, imag} */,
  {32'h4128c649, 32'hc10ec217} /* (21, 28, 24) {real, imag} */,
  {32'h4162abd0, 32'hbf5d6ac8} /* (21, 28, 23) {real, imag} */,
  {32'h40c90202, 32'h4104c548} /* (21, 28, 22) {real, imag} */,
  {32'h4005aa08, 32'h40c40ad4} /* (21, 28, 21) {real, imag} */,
  {32'hbf8566d6, 32'hbfe1d96c} /* (21, 28, 20) {real, imag} */,
  {32'hc0aca51c, 32'h408255ee} /* (21, 28, 19) {real, imag} */,
  {32'hc15605d2, 32'h417c2cd0} /* (21, 28, 18) {real, imag} */,
  {32'hc1643016, 32'h41a7830e} /* (21, 28, 17) {real, imag} */,
  {32'hc0b41cb2, 32'h40f035a2} /* (21, 28, 16) {real, imag} */,
  {32'h40a35cb1, 32'h3f4ab5e0} /* (21, 28, 15) {real, imag} */,
  {32'h401cb1b1, 32'hc1065a2a} /* (21, 28, 14) {real, imag} */,
  {32'hc0bf15a2, 32'hc0067ab4} /* (21, 28, 13) {real, imag} */,
  {32'hc13d51f2, 32'hbf111ce2} /* (21, 28, 12) {real, imag} */,
  {32'hbf3eaed2, 32'hc0dee758} /* (21, 28, 11) {real, imag} */,
  {32'h4106a761, 32'hc12beef9} /* (21, 28, 10) {real, imag} */,
  {32'h411580fd, 32'hc1148c02} /* (21, 28, 9) {real, imag} */,
  {32'h40505d2e, 32'hc0d30156} /* (21, 28, 8) {real, imag} */,
  {32'hc0a17be4, 32'hbf9c89a2} /* (21, 28, 7) {real, imag} */,
  {32'hbce7c680, 32'hc02bdf70} /* (21, 28, 6) {real, imag} */,
  {32'h4112ee78, 32'hc127e6b7} /* (21, 28, 5) {real, imag} */,
  {32'h415f715b, 32'h3d5c0730} /* (21, 28, 4) {real, imag} */,
  {32'hbf39e3aa, 32'h4104595d} /* (21, 28, 3) {real, imag} */,
  {32'h40f68a6a, 32'hbac4e800} /* (21, 28, 2) {real, imag} */,
  {32'h4111de30, 32'h400ee224} /* (21, 28, 1) {real, imag} */,
  {32'hbf9b3ab1, 32'h40404b8b} /* (21, 28, 0) {real, imag} */,
  {32'hc0e11af3, 32'h3f820604} /* (21, 27, 31) {real, imag} */,
  {32'hc129bf86, 32'hc092bf29} /* (21, 27, 30) {real, imag} */,
  {32'hc13636c0, 32'hc11c3b20} /* (21, 27, 29) {real, imag} */,
  {32'hc12a0c0b, 32'hc0373075} /* (21, 27, 28) {real, imag} */,
  {32'hc1b996a5, 32'hc0d3b202} /* (21, 27, 27) {real, imag} */,
  {32'hc157ef38, 32'hc0f56d28} /* (21, 27, 26) {real, imag} */,
  {32'hc0946543, 32'h3ffd63dc} /* (21, 27, 25) {real, imag} */,
  {32'hbe2c0580, 32'h3ea695e0} /* (21, 27, 24) {real, imag} */,
  {32'hc098f7bc, 32'hbe01bee0} /* (21, 27, 23) {real, imag} */,
  {32'hc1168e79, 32'hbf2857a0} /* (21, 27, 22) {real, imag} */,
  {32'hc0bfe624, 32'hbfb39e42} /* (21, 27, 21) {real, imag} */,
  {32'h40bfd066, 32'hc118a626} /* (21, 27, 20) {real, imag} */,
  {32'h40920f89, 32'hc09f60b5} /* (21, 27, 19) {real, imag} */,
  {32'h40c72b2e, 32'hbf11bccd} /* (21, 27, 18) {real, imag} */,
  {32'h4105de16, 32'hbe0e5834} /* (21, 27, 17) {real, imag} */,
  {32'h40b509af, 32'h3f2515f0} /* (21, 27, 16) {real, imag} */,
  {32'h410e4ee7, 32'h402de8d3} /* (21, 27, 15) {real, imag} */,
  {32'h40c0cd95, 32'h408d8756} /* (21, 27, 14) {real, imag} */,
  {32'h4031be2d, 32'hc0d3b0ce} /* (21, 27, 13) {real, imag} */,
  {32'h41197f44, 32'hc08465a0} /* (21, 27, 12) {real, imag} */,
  {32'h413f7b0b, 32'h40f8bca0} /* (21, 27, 11) {real, imag} */,
  {32'hc0b35f6e, 32'h40d241d7} /* (21, 27, 10) {real, imag} */,
  {32'hc0f36eba, 32'h40cda7ae} /* (21, 27, 9) {real, imag} */,
  {32'hbdd98380, 32'h40f3c1ac} /* (21, 27, 8) {real, imag} */,
  {32'hc046487f, 32'h404cca78} /* (21, 27, 7) {real, imag} */,
  {32'h408d446e, 32'h4006d7c4} /* (21, 27, 6) {real, imag} */,
  {32'h3dea7320, 32'hc1111e88} /* (21, 27, 5) {real, imag} */,
  {32'hbfd96c65, 32'hc0812234} /* (21, 27, 4) {real, imag} */,
  {32'hc05d359c, 32'h3f3455e8} /* (21, 27, 3) {real, imag} */,
  {32'hbf83454d, 32'h3f3d3345} /* (21, 27, 2) {real, imag} */,
  {32'hc019106d, 32'h40515105} /* (21, 27, 1) {real, imag} */,
  {32'hc0ad6a28, 32'h3f45e874} /* (21, 27, 0) {real, imag} */,
  {32'h40aedc5d, 32'h40a2ed7a} /* (21, 26, 31) {real, imag} */,
  {32'h40a5454e, 32'h40897194} /* (21, 26, 30) {real, imag} */,
  {32'h404e8272, 32'hc0b67911} /* (21, 26, 29) {real, imag} */,
  {32'h3ea1f6e0, 32'hbfe1c682} /* (21, 26, 28) {real, imag} */,
  {32'hc0e266ba, 32'hc0c7237e} /* (21, 26, 27) {real, imag} */,
  {32'h3f175670, 32'hc0f98442} /* (21, 26, 26) {real, imag} */,
  {32'h40d53720, 32'hbfd4153c} /* (21, 26, 25) {real, imag} */,
  {32'hc01ba057, 32'h400cd348} /* (21, 26, 24) {real, imag} */,
  {32'hc154e862, 32'h407185e0} /* (21, 26, 23) {real, imag} */,
  {32'hc0beb58a, 32'h3e8f11d0} /* (21, 26, 22) {real, imag} */,
  {32'hc0432510, 32'hc09d6ccf} /* (21, 26, 21) {real, imag} */,
  {32'hc159b3b5, 32'hbf825b06} /* (21, 26, 20) {real, imag} */,
  {32'hc0e227d3, 32'h40b9028e} /* (21, 26, 19) {real, imag} */,
  {32'hc048dde7, 32'h3ff716e0} /* (21, 26, 18) {real, imag} */,
  {32'hc102b891, 32'h40cf3d6e} /* (21, 26, 17) {real, imag} */,
  {32'hc10d50ee, 32'hc095d32e} /* (21, 26, 16) {real, imag} */,
  {32'hc0d5c6c2, 32'hbf89f16f} /* (21, 26, 15) {real, imag} */,
  {32'hc0215962, 32'hbf0ead0e} /* (21, 26, 14) {real, imag} */,
  {32'hc133e037, 32'hbf55cc5e} /* (21, 26, 13) {real, imag} */,
  {32'hc16ef6d8, 32'h3da79180} /* (21, 26, 12) {real, imag} */,
  {32'hc12e2539, 32'h408d6904} /* (21, 26, 11) {real, imag} */,
  {32'hc0034f22, 32'h412af361} /* (21, 26, 10) {real, imag} */,
  {32'h40c9cab2, 32'h411a8159} /* (21, 26, 9) {real, imag} */,
  {32'h4047fda9, 32'h40a9980e} /* (21, 26, 8) {real, imag} */,
  {32'h3e246f34, 32'h40efe64c} /* (21, 26, 7) {real, imag} */,
  {32'h40674afb, 32'h4095d137} /* (21, 26, 6) {real, imag} */,
  {32'hc0a5a7e4, 32'h40547337} /* (21, 26, 5) {real, imag} */,
  {32'hc0b91275, 32'hc011860f} /* (21, 26, 4) {real, imag} */,
  {32'h4062b6e9, 32'hc0f40bed} /* (21, 26, 3) {real, imag} */,
  {32'h410c707a, 32'hc09a8553} /* (21, 26, 2) {real, imag} */,
  {32'hc0383c4e, 32'hc044c7d4} /* (21, 26, 1) {real, imag} */,
  {32'h3e9a4ad6, 32'hc0ba73aa} /* (21, 26, 0) {real, imag} */,
  {32'h3b842c00, 32'h41099545} /* (21, 25, 31) {real, imag} */,
  {32'hc033f116, 32'h4034a90b} /* (21, 25, 30) {real, imag} */,
  {32'hc09714aa, 32'hc0efbe10} /* (21, 25, 29) {real, imag} */,
  {32'hbe872724, 32'hc063f82a} /* (21, 25, 28) {real, imag} */,
  {32'h40a9e645, 32'hbd0e2da0} /* (21, 25, 27) {real, imag} */,
  {32'h3d2c4400, 32'h4048ecfa} /* (21, 25, 26) {real, imag} */,
  {32'hc039ea14, 32'h4114714d} /* (21, 25, 25) {real, imag} */,
  {32'hbec5bfa0, 32'h3f9506c4} /* (21, 25, 24) {real, imag} */,
  {32'h4104d706, 32'hc092152a} /* (21, 25, 23) {real, imag} */,
  {32'h3fa62e70, 32'hc02fb859} /* (21, 25, 22) {real, imag} */,
  {32'h3ece5994, 32'hc0169f28} /* (21, 25, 21) {real, imag} */,
  {32'hc0eefae3, 32'h40061156} /* (21, 25, 20) {real, imag} */,
  {32'hc19c9570, 32'hc0e5359f} /* (21, 25, 19) {real, imag} */,
  {32'hc1b6be44, 32'hc1122762} /* (21, 25, 18) {real, imag} */,
  {32'hc131cba4, 32'hc0861d9a} /* (21, 25, 17) {real, imag} */,
  {32'hbee36f34, 32'hc02d256a} /* (21, 25, 16) {real, imag} */,
  {32'hc096ed18, 32'hc04c3a08} /* (21, 25, 15) {real, imag} */,
  {32'hc04f4cca, 32'h40f4b0ae} /* (21, 25, 14) {real, imag} */,
  {32'hbfaa93a8, 32'h3fc00c60} /* (21, 25, 13) {real, imag} */,
  {32'hc110c9d6, 32'hc00cbf44} /* (21, 25, 12) {real, imag} */,
  {32'hc06b59ea, 32'h40240029} /* (21, 25, 11) {real, imag} */,
  {32'hc0b6fe5c, 32'hc082d0ec} /* (21, 25, 10) {real, imag} */,
  {32'hc053cf12, 32'hc092fe76} /* (21, 25, 9) {real, imag} */,
  {32'h40784234, 32'hc0841762} /* (21, 25, 8) {real, imag} */,
  {32'hc0c42fdb, 32'hc027647b} /* (21, 25, 7) {real, imag} */,
  {32'hc0ef4b55, 32'hbf945714} /* (21, 25, 6) {real, imag} */,
  {32'hbf5699dc, 32'h3fb8057c} /* (21, 25, 5) {real, imag} */,
  {32'h40b36cd1, 32'h3f272918} /* (21, 25, 4) {real, imag} */,
  {32'h412786b8, 32'h3f540940} /* (21, 25, 3) {real, imag} */,
  {32'h4004d376, 32'hc00446b8} /* (21, 25, 2) {real, imag} */,
  {32'h40b713bc, 32'hc042b8c1} /* (21, 25, 1) {real, imag} */,
  {32'h4080c3ce, 32'h3f21c325} /* (21, 25, 0) {real, imag} */,
  {32'h3f7b054c, 32'hbf51f948} /* (21, 24, 31) {real, imag} */,
  {32'h40868b5c, 32'h3f4ce984} /* (21, 24, 30) {real, imag} */,
  {32'h40c11c28, 32'hc0463344} /* (21, 24, 29) {real, imag} */,
  {32'hc0f5d494, 32'h3f811e98} /* (21, 24, 28) {real, imag} */,
  {32'hc052cfc3, 32'h410e25b6} /* (21, 24, 27) {real, imag} */,
  {32'h3fb059fc, 32'h40cc498e} /* (21, 24, 26) {real, imag} */,
  {32'h3ea76524, 32'hc1019eed} /* (21, 24, 25) {real, imag} */,
  {32'h40b6d68a, 32'hc01a5b08} /* (21, 24, 24) {real, imag} */,
  {32'h41009cab, 32'h404b9287} /* (21, 24, 23) {real, imag} */,
  {32'h3feb54e4, 32'hc06964ae} /* (21, 24, 22) {real, imag} */,
  {32'hbf1e48e2, 32'hbffa1d46} /* (21, 24, 21) {real, imag} */,
  {32'h4025c63a, 32'hc09f96d8} /* (21, 24, 20) {real, imag} */,
  {32'hbefad51a, 32'hbe5c35a0} /* (21, 24, 19) {real, imag} */,
  {32'hbfbbe5a6, 32'h4038946a} /* (21, 24, 18) {real, imag} */,
  {32'hc020fbe8, 32'h40164be6} /* (21, 24, 17) {real, imag} */,
  {32'hbda06870, 32'hbf92ed3e} /* (21, 24, 16) {real, imag} */,
  {32'hbe9d8990, 32'hc10c770c} /* (21, 24, 15) {real, imag} */,
  {32'hbf367c00, 32'hc0cffcbd} /* (21, 24, 14) {real, imag} */,
  {32'hbec88bc0, 32'hc052a03c} /* (21, 24, 13) {real, imag} */,
  {32'h4096905c, 32'h3f44139a} /* (21, 24, 12) {real, imag} */,
  {32'hbf9a140c, 32'hbfcdb066} /* (21, 24, 11) {real, imag} */,
  {32'hbfb30daf, 32'hc095f60a} /* (21, 24, 10) {real, imag} */,
  {32'h3e8d0ca8, 32'h3f4a639c} /* (21, 24, 9) {real, imag} */,
  {32'h3f7d27b8, 32'h40a8b308} /* (21, 24, 8) {real, imag} */,
  {32'h404b704c, 32'h40b0ccac} /* (21, 24, 7) {real, imag} */,
  {32'h3f2bd5b8, 32'hc0a039e8} /* (21, 24, 6) {real, imag} */,
  {32'h3fefa292, 32'hc105dabc} /* (21, 24, 5) {real, imag} */,
  {32'h40dd0458, 32'h4064a6b4} /* (21, 24, 4) {real, imag} */,
  {32'h3f420528, 32'h40870148} /* (21, 24, 3) {real, imag} */,
  {32'hc083c5c8, 32'hbfb69c54} /* (21, 24, 2) {real, imag} */,
  {32'hc0e9a86c, 32'h3fd84938} /* (21, 24, 1) {real, imag} */,
  {32'hc027a1dc, 32'hbe6ee100} /* (21, 24, 0) {real, imag} */,
  {32'h4004cfa0, 32'h40b93070} /* (21, 23, 31) {real, imag} */,
  {32'hbe47fc00, 32'h41283259} /* (21, 23, 30) {real, imag} */,
  {32'h3f70ed79, 32'h40b2e466} /* (21, 23, 29) {real, imag} */,
  {32'h3f9ab666, 32'h4045b6f7} /* (21, 23, 28) {real, imag} */,
  {32'h4086a7cf, 32'hbfc825dc} /* (21, 23, 27) {real, imag} */,
  {32'h3facf8f4, 32'h401bb164} /* (21, 23, 26) {real, imag} */,
  {32'hbd335420, 32'h3f4d1b40} /* (21, 23, 25) {real, imag} */,
  {32'h3f1088d2, 32'h40b9e81c} /* (21, 23, 24) {real, imag} */,
  {32'hbd791980, 32'h4107e7f2} /* (21, 23, 23) {real, imag} */,
  {32'h3fcda168, 32'h40cdc2a2} /* (21, 23, 22) {real, imag} */,
  {32'h4096900c, 32'h40d91e4f} /* (21, 23, 21) {real, imag} */,
  {32'h40a26cc8, 32'h40d18ce8} /* (21, 23, 20) {real, imag} */,
  {32'h40379042, 32'h4113c879} /* (21, 23, 19) {real, imag} */,
  {32'h3e006f20, 32'h4091dcf2} /* (21, 23, 18) {real, imag} */,
  {32'hc03b56eb, 32'hbfde6112} /* (21, 23, 17) {real, imag} */,
  {32'hbe378000, 32'h3f10cf88} /* (21, 23, 16) {real, imag} */,
  {32'h408db236, 32'h4018b486} /* (21, 23, 15) {real, imag} */,
  {32'h404f0f42, 32'hc0870a3d} /* (21, 23, 14) {real, imag} */,
  {32'hbed66d90, 32'hc02faa3a} /* (21, 23, 13) {real, imag} */,
  {32'hbf4c461c, 32'hbed700ee} /* (21, 23, 12) {real, imag} */,
  {32'hc0b13cb9, 32'hbd93ac80} /* (21, 23, 11) {real, imag} */,
  {32'hc02f5d43, 32'hbe9669a8} /* (21, 23, 10) {real, imag} */,
  {32'hc01b7bc4, 32'hc08b61ce} /* (21, 23, 9) {real, imag} */,
  {32'h3f44857a, 32'hc0d13924} /* (21, 23, 8) {real, imag} */,
  {32'hc0a71d97, 32'hbc6a0500} /* (21, 23, 7) {real, imag} */,
  {32'h3fd14dde, 32'h406a7710} /* (21, 23, 6) {real, imag} */,
  {32'h413341ef, 32'hc06c2564} /* (21, 23, 5) {real, imag} */,
  {32'h40d4c2ca, 32'hbeef0b40} /* (21, 23, 4) {real, imag} */,
  {32'h404ac86a, 32'h3fb58c3e} /* (21, 23, 3) {real, imag} */,
  {32'h411c7b06, 32'h3f3eed94} /* (21, 23, 2) {real, imag} */,
  {32'h40aac371, 32'hc07298ee} /* (21, 23, 1) {real, imag} */,
  {32'hbf6f2d7c, 32'hbf3ff055} /* (21, 23, 0) {real, imag} */,
  {32'hc082bda4, 32'hc09537ed} /* (21, 22, 31) {real, imag} */,
  {32'hbffbf9ec, 32'hc1248f5d} /* (21, 22, 30) {real, imag} */,
  {32'hbeb98ae4, 32'hc0c088e0} /* (21, 22, 29) {real, imag} */,
  {32'h3f1aa37a, 32'hbfdf856c} /* (21, 22, 28) {real, imag} */,
  {32'hbe0465e0, 32'hc0604e90} /* (21, 22, 27) {real, imag} */,
  {32'hbf39c4e0, 32'hc0471b7f} /* (21, 22, 26) {real, imag} */,
  {32'hbfa3c1e5, 32'hbe91dff8} /* (21, 22, 25) {real, imag} */,
  {32'h3fd00f98, 32'hc06ca932} /* (21, 22, 24) {real, imag} */,
  {32'h4049f1f6, 32'hc139ceef} /* (21, 22, 23) {real, imag} */,
  {32'hc007d549, 32'hc0c30550} /* (21, 22, 22) {real, imag} */,
  {32'h3eb6db74, 32'h405038e0} /* (21, 22, 21) {real, imag} */,
  {32'h40dc1c40, 32'h40a1a513} /* (21, 22, 20) {real, imag} */,
  {32'h4114c562, 32'hc0ecce2a} /* (21, 22, 19) {real, imag} */,
  {32'hbf3e7b2e, 32'hc072f3c4} /* (21, 22, 18) {real, imag} */,
  {32'hc0ab6d1d, 32'hbff83aea} /* (21, 22, 17) {real, imag} */,
  {32'h403f0e5a, 32'h3f00eae8} /* (21, 22, 16) {real, imag} */,
  {32'h4039674a, 32'h40107e47} /* (21, 22, 15) {real, imag} */,
  {32'hc0b102fa, 32'hc084b828} /* (21, 22, 14) {real, imag} */,
  {32'hc082d210, 32'h4043a880} /* (21, 22, 13) {real, imag} */,
  {32'h40673a99, 32'h4074faa6} /* (21, 22, 12) {real, imag} */,
  {32'h3fc8c8c0, 32'hbe491630} /* (21, 22, 11) {real, imag} */,
  {32'hc0207dcc, 32'hc04f9c82} /* (21, 22, 10) {real, imag} */,
  {32'h4083f1e0, 32'hc094da6a} /* (21, 22, 9) {real, imag} */,
  {32'h40672b36, 32'hbf1f05ee} /* (21, 22, 8) {real, imag} */,
  {32'hc0624218, 32'hc0525d4a} /* (21, 22, 7) {real, imag} */,
  {32'hc005da9d, 32'hc05772ce} /* (21, 22, 6) {real, imag} */,
  {32'h3e43b59c, 32'hbcfc73f0} /* (21, 22, 5) {real, imag} */,
  {32'hc04e758a, 32'h3fbf7721} /* (21, 22, 4) {real, imag} */,
  {32'hc0eeb519, 32'hbf325b18} /* (21, 22, 3) {real, imag} */,
  {32'hc0ad7048, 32'h3e0a9f38} /* (21, 22, 2) {real, imag} */,
  {32'hbfc78f0b, 32'hbfacec62} /* (21, 22, 1) {real, imag} */,
  {32'hbffda44c, 32'hc002b9e0} /* (21, 22, 0) {real, imag} */,
  {32'hc048ab84, 32'hc031718b} /* (21, 21, 31) {real, imag} */,
  {32'hc0a584e6, 32'hc0743bca} /* (21, 21, 30) {real, imag} */,
  {32'hbf467f7b, 32'h3f7f6558} /* (21, 21, 29) {real, imag} */,
  {32'hbf9b0108, 32'h402fda22} /* (21, 21, 28) {real, imag} */,
  {32'hc04e27e6, 32'h4101be67} /* (21, 21, 27) {real, imag} */,
  {32'h3ee1c130, 32'h40e66c4e} /* (21, 21, 26) {real, imag} */,
  {32'hc069a6e4, 32'h40a2e85a} /* (21, 21, 25) {real, imag} */,
  {32'hbfea1284, 32'h3fa8aec2} /* (21, 21, 24) {real, imag} */,
  {32'h3fbb85ba, 32'h3ff43eda} /* (21, 21, 23) {real, imag} */,
  {32'h3f3c544a, 32'h407e5f7c} /* (21, 21, 22) {real, imag} */,
  {32'h3f49f114, 32'h404f88d0} /* (21, 21, 21) {real, imag} */,
  {32'h40517bf7, 32'h3fdc385d} /* (21, 21, 20) {real, imag} */,
  {32'h3fc80643, 32'h3f5204b2} /* (21, 21, 19) {real, imag} */,
  {32'hc0037930, 32'h403c96ea} /* (21, 21, 18) {real, imag} */,
  {32'h3ea70440, 32'hbece270a} /* (21, 21, 17) {real, imag} */,
  {32'h405ef854, 32'h3f850a7a} /* (21, 21, 16) {real, imag} */,
  {32'h40192f63, 32'hc09a43a3} /* (21, 21, 15) {real, imag} */,
  {32'hbf960e55, 32'hc02e6bdd} /* (21, 21, 14) {real, imag} */,
  {32'h3f92bed6, 32'h3fdff69e} /* (21, 21, 13) {real, imag} */,
  {32'h3f05008e, 32'h401c851c} /* (21, 21, 12) {real, imag} */,
  {32'hbe1c1960, 32'h3fe7f583} /* (21, 21, 11) {real, imag} */,
  {32'hc04d46b9, 32'h40030cea} /* (21, 21, 10) {real, imag} */,
  {32'hc07eb909, 32'hbfbac5e7} /* (21, 21, 9) {real, imag} */,
  {32'h3f671ec0, 32'hbfe1ad7e} /* (21, 21, 8) {real, imag} */,
  {32'h402c494b, 32'h3ebe1760} /* (21, 21, 7) {real, imag} */,
  {32'h408373fe, 32'hbf449470} /* (21, 21, 6) {real, imag} */,
  {32'h40bb4084, 32'h400ce22e} /* (21, 21, 5) {real, imag} */,
  {32'h406eaf22, 32'h3fd92151} /* (21, 21, 4) {real, imag} */,
  {32'h3f92b894, 32'hbfcb4a15} /* (21, 21, 3) {real, imag} */,
  {32'hc072b382, 32'hbfcad03a} /* (21, 21, 2) {real, imag} */,
  {32'hc10e6b3b, 32'hbf44beb4} /* (21, 21, 1) {real, imag} */,
  {32'hc105390b, 32'h3fe52ed0} /* (21, 21, 0) {real, imag} */,
  {32'hc03c78f0, 32'hbfb0ad86} /* (21, 20, 31) {real, imag} */,
  {32'hc03ef6b1, 32'hbf2b5922} /* (21, 20, 30) {real, imag} */,
  {32'h3e51d3a8, 32'hbfa71794} /* (21, 20, 29) {real, imag} */,
  {32'h3fd7c58c, 32'hc029e554} /* (21, 20, 28) {real, imag} */,
  {32'hbee71be0, 32'h3bc0d900} /* (21, 20, 27) {real, imag} */,
  {32'hbfb80ba6, 32'h40828e82} /* (21, 20, 26) {real, imag} */,
  {32'h402f64c2, 32'h400bfd51} /* (21, 20, 25) {real, imag} */,
  {32'h3ed1ff64, 32'hbeff2c6a} /* (21, 20, 24) {real, imag} */,
  {32'h3f60cf7c, 32'hc05b0fe8} /* (21, 20, 23) {real, imag} */,
  {32'hbfb9583b, 32'hbfff9ade} /* (21, 20, 22) {real, imag} */,
  {32'hc01d84e1, 32'h3fe8a1c2} /* (21, 20, 21) {real, imag} */,
  {32'hc0257ac6, 32'hbfa8cce6} /* (21, 20, 20) {real, imag} */,
  {32'hc0999812, 32'h3f17abf4} /* (21, 20, 19) {real, imag} */,
  {32'h3f717ef4, 32'hbf2d0ede} /* (21, 20, 18) {real, imag} */,
  {32'hbf92cb85, 32'hbf665ae8} /* (21, 20, 17) {real, imag} */,
  {32'hbf39ebea, 32'hc0043dd3} /* (21, 20, 16) {real, imag} */,
  {32'hbf93142e, 32'hbf3b07f2} /* (21, 20, 15) {real, imag} */,
  {32'h3ce35200, 32'h4022c768} /* (21, 20, 14) {real, imag} */,
  {32'h4055a8bc, 32'h40967862} /* (21, 20, 13) {real, imag} */,
  {32'h3ea63b64, 32'h403e7e56} /* (21, 20, 12) {real, imag} */,
  {32'h3fd49c9d, 32'hbf564c04} /* (21, 20, 11) {real, imag} */,
  {32'h40323885, 32'h3df81230} /* (21, 20, 10) {real, imag} */,
  {32'h40960d3f, 32'h4097e3fb} /* (21, 20, 9) {real, imag} */,
  {32'h409a94f3, 32'h4073987a} /* (21, 20, 8) {real, imag} */,
  {32'h4036c74a, 32'h40307e30} /* (21, 20, 7) {real, imag} */,
  {32'h408250db, 32'h400a8e58} /* (21, 20, 6) {real, imag} */,
  {32'h40077c97, 32'h3eccbe58} /* (21, 20, 5) {real, imag} */,
  {32'hc04b8c8b, 32'h3f23d15d} /* (21, 20, 4) {real, imag} */,
  {32'hc04a7098, 32'h40798583} /* (21, 20, 3) {real, imag} */,
  {32'h3f1c74c0, 32'h400d86ff} /* (21, 20, 2) {real, imag} */,
  {32'hbdfdc050, 32'hc03567e7} /* (21, 20, 1) {real, imag} */,
  {32'hc029e119, 32'h3fb19150} /* (21, 20, 0) {real, imag} */,
  {32'hbfa31a27, 32'hc045b8f0} /* (21, 19, 31) {real, imag} */,
  {32'hc011f946, 32'hc00a4f1e} /* (21, 19, 30) {real, imag} */,
  {32'hbdf68fc8, 32'h3d769c80} /* (21, 19, 29) {real, imag} */,
  {32'h4011c4c0, 32'hc002ad6e} /* (21, 19, 28) {real, imag} */,
  {32'h401a6ee0, 32'hbff2e8ff} /* (21, 19, 27) {real, imag} */,
  {32'h40052906, 32'h3f1c15d0} /* (21, 19, 26) {real, imag} */,
  {32'h3f83aebf, 32'h3f3a9c54} /* (21, 19, 25) {real, imag} */,
  {32'hbe846bb0, 32'h3f91db97} /* (21, 19, 24) {real, imag} */,
  {32'h3f40e90c, 32'h3fe67db4} /* (21, 19, 23) {real, imag} */,
  {32'h408e6742, 32'hbcde2600} /* (21, 19, 22) {real, imag} */,
  {32'h40490543, 32'hc02ddd2b} /* (21, 19, 21) {real, imag} */,
  {32'hbf88f774, 32'hbe7e9234} /* (21, 19, 20) {real, imag} */,
  {32'h3e2a4738, 32'hbf0f3d10} /* (21, 19, 19) {real, imag} */,
  {32'hbeab5f9c, 32'hc03bd55e} /* (21, 19, 18) {real, imag} */,
  {32'hbf1b2e6c, 32'hc041e27c} /* (21, 19, 17) {real, imag} */,
  {32'h402ba615, 32'hc0363ea6} /* (21, 19, 16) {real, imag} */,
  {32'h402af9f6, 32'h3e662820} /* (21, 19, 15) {real, imag} */,
  {32'h3fc443e9, 32'hbf107098} /* (21, 19, 14) {real, imag} */,
  {32'hbeae4940, 32'hbf765f9c} /* (21, 19, 13) {real, imag} */,
  {32'h3f07e0f0, 32'h3ed3cffa} /* (21, 19, 12) {real, imag} */,
  {32'hbfdbc50e, 32'hbe08f27c} /* (21, 19, 11) {real, imag} */,
  {32'hc0199766, 32'hbe909c48} /* (21, 19, 10) {real, imag} */,
  {32'h3f7f6540, 32'hbf9ee5b6} /* (21, 19, 9) {real, imag} */,
  {32'h3f32d21a, 32'h3e809a54} /* (21, 19, 8) {real, imag} */,
  {32'hbeea4ef0, 32'h3f50ec80} /* (21, 19, 7) {real, imag} */,
  {32'hbe1d8b88, 32'h402de35e} /* (21, 19, 6) {real, imag} */,
  {32'h3f95cfd0, 32'h4054339c} /* (21, 19, 5) {real, imag} */,
  {32'h3f1f4264, 32'h4024194c} /* (21, 19, 4) {real, imag} */,
  {32'h3fe02e60, 32'h3edf1698} /* (21, 19, 3) {real, imag} */,
  {32'hbfc9b843, 32'hbf81631c} /* (21, 19, 2) {real, imag} */,
  {32'h40094126, 32'hbf918cc0} /* (21, 19, 1) {real, imag} */,
  {32'h402a7344, 32'hbf7bc868} /* (21, 19, 0) {real, imag} */,
  {32'hbf420fd8, 32'h3f3df468} /* (21, 18, 31) {real, imag} */,
  {32'h3f9b53ee, 32'h3eefbf28} /* (21, 18, 30) {real, imag} */,
  {32'hbf4b9998, 32'h3f03c8dc} /* (21, 18, 29) {real, imag} */,
  {32'hbf179372, 32'h3fd8534e} /* (21, 18, 28) {real, imag} */,
  {32'h3e983cf8, 32'hbeec8570} /* (21, 18, 27) {real, imag} */,
  {32'h3df5dd60, 32'hbf7ea0d2} /* (21, 18, 26) {real, imag} */,
  {32'h3fc482ac, 32'hbf15e786} /* (21, 18, 25) {real, imag} */,
  {32'h40038bf2, 32'h3fd56366} /* (21, 18, 24) {real, imag} */,
  {32'h3f94d912, 32'h3f631838} /* (21, 18, 23) {real, imag} */,
  {32'h3fb69b03, 32'h40114c4f} /* (21, 18, 22) {real, imag} */,
  {32'h3fa3916e, 32'h3f1aa7fe} /* (21, 18, 21) {real, imag} */,
  {32'h3fb11907, 32'h3e78c880} /* (21, 18, 20) {real, imag} */,
  {32'h40095cde, 32'h3e0dc23c} /* (21, 18, 19) {real, imag} */,
  {32'h403381b6, 32'hc0060bce} /* (21, 18, 18) {real, imag} */,
  {32'h3f96d478, 32'hc054077d} /* (21, 18, 17) {real, imag} */,
  {32'hbf95212a, 32'h3f850d8b} /* (21, 18, 16) {real, imag} */,
  {32'hbfa20323, 32'h3fc3da94} /* (21, 18, 15) {real, imag} */,
  {32'h3e1ccdd0, 32'h3eb75334} /* (21, 18, 14) {real, imag} */,
  {32'hc0445798, 32'h3e326cec} /* (21, 18, 13) {real, imag} */,
  {32'h3f555e14, 32'h406ffb37} /* (21, 18, 12) {real, imag} */,
  {32'h3fa48c80, 32'h404d4476} /* (21, 18, 11) {real, imag} */,
  {32'hbfac7f3c, 32'h403f6b0f} /* (21, 18, 10) {real, imag} */,
  {32'hc03ea9cc, 32'h40052ce2} /* (21, 18, 9) {real, imag} */,
  {32'hbfbe3a6e, 32'h400b710e} /* (21, 18, 8) {real, imag} */,
  {32'hbf8c1e20, 32'hbea00e14} /* (21, 18, 7) {real, imag} */,
  {32'hc02a8598, 32'hbfb3406b} /* (21, 18, 6) {real, imag} */,
  {32'hbf3aad92, 32'h3f1004ab} /* (21, 18, 5) {real, imag} */,
  {32'hbfe9c1b0, 32'h3ec66510} /* (21, 18, 4) {real, imag} */,
  {32'hbfeb64da, 32'hbe13b674} /* (21, 18, 3) {real, imag} */,
  {32'h3f33d824, 32'hbde18830} /* (21, 18, 2) {real, imag} */,
  {32'hbfc80323, 32'h3dcacd58} /* (21, 18, 1) {real, imag} */,
  {32'hbfaf74df, 32'h3f28d6ca} /* (21, 18, 0) {real, imag} */,
  {32'h3e4858d8, 32'h3e7a51c0} /* (21, 17, 31) {real, imag} */,
  {32'h3f866a1c, 32'h3fd40ad8} /* (21, 17, 30) {real, imag} */,
  {32'h3fb275b9, 32'h3f8fd364} /* (21, 17, 29) {real, imag} */,
  {32'hbf389a6b, 32'h3f5f6301} /* (21, 17, 28) {real, imag} */,
  {32'h40468596, 32'h3f584737} /* (21, 17, 27) {real, imag} */,
  {32'h4068a6f7, 32'h3de557f0} /* (21, 17, 26) {real, imag} */,
  {32'h3f52e9f8, 32'hbf36f1bc} /* (21, 17, 25) {real, imag} */,
  {32'h3f3af31c, 32'hbf17bda8} /* (21, 17, 24) {real, imag} */,
  {32'h3f2d4b28, 32'h3fcd69b2} /* (21, 17, 23) {real, imag} */,
  {32'hbfa1a42a, 32'h3e66d110} /* (21, 17, 22) {real, imag} */,
  {32'hbc6d8480, 32'hc045a580} /* (21, 17, 21) {real, imag} */,
  {32'h3f0da72a, 32'hc0681c84} /* (21, 17, 20) {real, imag} */,
  {32'h3ed46f0c, 32'hbfb5b5ba} /* (21, 17, 19) {real, imag} */,
  {32'h3f7946e0, 32'h3fec0be4} /* (21, 17, 18) {real, imag} */,
  {32'hbf8b5ee8, 32'h3fb6f44c} /* (21, 17, 17) {real, imag} */,
  {32'hbfee07d4, 32'h3f3c7d76} /* (21, 17, 16) {real, imag} */,
  {32'hbf35b380, 32'h3fe7b2cd} /* (21, 17, 15) {real, imag} */,
  {32'hbf0b41c0, 32'h3e77ca00} /* (21, 17, 14) {real, imag} */,
  {32'hbf428618, 32'hbf37a201} /* (21, 17, 13) {real, imag} */,
  {32'hbff41e8e, 32'hc0027bb2} /* (21, 17, 12) {real, imag} */,
  {32'hc00d30fc, 32'hbd171aa0} /* (21, 17, 11) {real, imag} */,
  {32'hbe401cf8, 32'h3fc47962} /* (21, 17, 10) {real, imag} */,
  {32'h40131bb4, 32'h3ebfccd0} /* (21, 17, 9) {real, imag} */,
  {32'hbf9f3c80, 32'h3f1cd6a2} /* (21, 17, 8) {real, imag} */,
  {32'h3a353000, 32'h3f87e1dc} /* (21, 17, 7) {real, imag} */,
  {32'h3fcfbc38, 32'h3f539a24} /* (21, 17, 6) {real, imag} */,
  {32'hbdd02bc0, 32'h3f6404a8} /* (21, 17, 5) {real, imag} */,
  {32'h3f3b36b0, 32'hbf5e7280} /* (21, 17, 4) {real, imag} */,
  {32'h3f55869a, 32'h3f631d5d} /* (21, 17, 3) {real, imag} */,
  {32'h3f0a2d28, 32'hbe9df1e8} /* (21, 17, 2) {real, imag} */,
  {32'h3f829516, 32'hc0397d0d} /* (21, 17, 1) {real, imag} */,
  {32'h3e0dff80, 32'hbf94f5bb} /* (21, 17, 0) {real, imag} */,
  {32'hbfc2988e, 32'hbe09c120} /* (21, 16, 31) {real, imag} */,
  {32'h3f121800, 32'hbea0dce0} /* (21, 16, 30) {real, imag} */,
  {32'h3ffbc850, 32'h40074ea3} /* (21, 16, 29) {real, imag} */,
  {32'h3f9faa68, 32'h3f9532ac} /* (21, 16, 28) {real, imag} */,
  {32'hbf5a67bc, 32'hbfa4d37a} /* (21, 16, 27) {real, imag} */,
  {32'hbf29fcfd, 32'hbef60e3c} /* (21, 16, 26) {real, imag} */,
  {32'h3f1fcf98, 32'hbfff1204} /* (21, 16, 25) {real, imag} */,
  {32'h3f16b140, 32'hbfb2945b} /* (21, 16, 24) {real, imag} */,
  {32'hbf564190, 32'hbcd73180} /* (21, 16, 23) {real, imag} */,
  {32'hbf212490, 32'h3fe4c6e0} /* (21, 16, 22) {real, imag} */,
  {32'h3f99176c, 32'h3f078154} /* (21, 16, 21) {real, imag} */,
  {32'h3f8635c8, 32'hbf3479a0} /* (21, 16, 20) {real, imag} */,
  {32'h3e82593c, 32'hbd32cfa0} /* (21, 16, 19) {real, imag} */,
  {32'h3f906090, 32'hbf8b62a0} /* (21, 16, 18) {real, imag} */,
  {32'hbf639d7a, 32'hbf79f590} /* (21, 16, 17) {real, imag} */,
  {32'h3ecb7810, 32'hbee3cc40} /* (21, 16, 16) {real, imag} */,
  {32'h406b50d2, 32'h3f3397f8} /* (21, 16, 15) {real, imag} */,
  {32'h3fe93a76, 32'h3e8e18c6} /* (21, 16, 14) {real, imag} */,
  {32'h3e9a7e78, 32'hbf83f5b1} /* (21, 16, 13) {real, imag} */,
  {32'h3e722e38, 32'hbf4b2ff8} /* (21, 16, 12) {real, imag} */,
  {32'h3f8d7c1e, 32'hbea15e40} /* (21, 16, 11) {real, imag} */,
  {32'h40267d4e, 32'hbea70340} /* (21, 16, 10) {real, imag} */,
  {32'h3fe6126e, 32'h400b564a} /* (21, 16, 9) {real, imag} */,
  {32'h4005a6de, 32'h403b7a7b} /* (21, 16, 8) {real, imag} */,
  {32'h3f7af8b8, 32'h3f70e845} /* (21, 16, 7) {real, imag} */,
  {32'hbff531ec, 32'hc03a32d4} /* (21, 16, 6) {real, imag} */,
  {32'h3efbb300, 32'hbd85cf00} /* (21, 16, 5) {real, imag} */,
  {32'h40146244, 32'h3fdf09b0} /* (21, 16, 4) {real, imag} */,
  {32'h3ebe2bd8, 32'hbf8958e4} /* (21, 16, 3) {real, imag} */,
  {32'hbf324a18, 32'hc0005a96} /* (21, 16, 2) {real, imag} */,
  {32'h3fe69b58, 32'hbfdb0b74} /* (21, 16, 1) {real, imag} */,
  {32'h3fb1d228, 32'h3e2331e0} /* (21, 16, 0) {real, imag} */,
  {32'h401a2be6, 32'h3ed75a00} /* (21, 15, 31) {real, imag} */,
  {32'h3f083d89, 32'h3ef3d0a0} /* (21, 15, 30) {real, imag} */,
  {32'hbe9ae3cc, 32'h3fefcb24} /* (21, 15, 29) {real, imag} */,
  {32'hbffe8dca, 32'h3f91ad98} /* (21, 15, 28) {real, imag} */,
  {32'hc02836f2, 32'hbeff261e} /* (21, 15, 27) {real, imag} */,
  {32'hbf3858e4, 32'h3e487b38} /* (21, 15, 26) {real, imag} */,
  {32'h3f514de8, 32'h3fee6526} /* (21, 15, 25) {real, imag} */,
  {32'hbfbc7c06, 32'h3f985d2c} /* (21, 15, 24) {real, imag} */,
  {32'hbdb57a40, 32'h3eaeafc8} /* (21, 15, 23) {real, imag} */,
  {32'hbfa30b9e, 32'hc00c3f59} /* (21, 15, 22) {real, imag} */,
  {32'hbfcdb9cf, 32'hc0531378} /* (21, 15, 21) {real, imag} */,
  {32'h3f55310a, 32'hc013c780} /* (21, 15, 20) {real, imag} */,
  {32'h3f2e790a, 32'hbef1a948} /* (21, 15, 19) {real, imag} */,
  {32'hbfad64d0, 32'h3f40a948} /* (21, 15, 18) {real, imag} */,
  {32'hbf591d80, 32'h3e8101e2} /* (21, 15, 17) {real, imag} */,
  {32'h402ce2a6, 32'hbed3e27c} /* (21, 15, 16) {real, imag} */,
  {32'h3fadc578, 32'h3fce7331} /* (21, 15, 15) {real, imag} */,
  {32'h403723f0, 32'h3f2329b0} /* (21, 15, 14) {real, imag} */,
  {32'h40072bf6, 32'h3e23076c} /* (21, 15, 13) {real, imag} */,
  {32'hbfc08652, 32'h3f8f7884} /* (21, 15, 12) {real, imag} */,
  {32'hbf627d52, 32'h402b693a} /* (21, 15, 11) {real, imag} */,
  {32'hbf8b2511, 32'h3feee45a} /* (21, 15, 10) {real, imag} */,
  {32'hc04217a2, 32'hbefe9010} /* (21, 15, 9) {real, imag} */,
  {32'hc05419b0, 32'h3fa39f31} /* (21, 15, 8) {real, imag} */,
  {32'hc0514db9, 32'h405ff046} /* (21, 15, 7) {real, imag} */,
  {32'hc02fd27c, 32'h402a94d1} /* (21, 15, 6) {real, imag} */,
  {32'h3d0e2f80, 32'h3e9b6b90} /* (21, 15, 5) {real, imag} */,
  {32'hbe258f40, 32'hbfff5798} /* (21, 15, 4) {real, imag} */,
  {32'h3fad782b, 32'hbf71d011} /* (21, 15, 3) {real, imag} */,
  {32'h407fec66, 32'hbfc96868} /* (21, 15, 2) {real, imag} */,
  {32'h3ffd35c6, 32'h3f00cde4} /* (21, 15, 1) {real, imag} */,
  {32'hbf45ddc8, 32'h3f84c9b1} /* (21, 15, 0) {real, imag} */,
  {32'hbfe018a8, 32'hbe140400} /* (21, 14, 31) {real, imag} */,
  {32'h3fb29136, 32'hc008656b} /* (21, 14, 30) {real, imag} */,
  {32'h3fa4830c, 32'hc00af107} /* (21, 14, 29) {real, imag} */,
  {32'h3f3cbf12, 32'hbe6e5b74} /* (21, 14, 28) {real, imag} */,
  {32'hc02b2e37, 32'h3f41af48} /* (21, 14, 27) {real, imag} */,
  {32'hbf74a64c, 32'hc02cbec4} /* (21, 14, 26) {real, imag} */,
  {32'h3ed47830, 32'hc00ea492} /* (21, 14, 25) {real, imag} */,
  {32'hc02a864a, 32'h40203e55} /* (21, 14, 24) {real, imag} */,
  {32'h3f2d4d6c, 32'h403c174e} /* (21, 14, 23) {real, imag} */,
  {32'h3fd30969, 32'h3fb3f196} /* (21, 14, 22) {real, imag} */,
  {32'hbe5d3bd0, 32'h3ff895d7} /* (21, 14, 21) {real, imag} */,
  {32'hbf8c6ed7, 32'h3fe9c210} /* (21, 14, 20) {real, imag} */,
  {32'hbed716b0, 32'h3f0dcbd3} /* (21, 14, 19) {real, imag} */,
  {32'hbee56c70, 32'h3ef8b880} /* (21, 14, 18) {real, imag} */,
  {32'hbf658bb0, 32'hbfd865d6} /* (21, 14, 17) {real, imag} */,
  {32'h3f62f154, 32'hbea2a1ec} /* (21, 14, 16) {real, imag} */,
  {32'h3f9b0133, 32'hbf0797fc} /* (21, 14, 15) {real, imag} */,
  {32'h4025c68d, 32'hbf8f8639} /* (21, 14, 14) {real, imag} */,
  {32'hbf1d56de, 32'hbf91cb54} /* (21, 14, 13) {real, imag} */,
  {32'hbff98dde, 32'hbfe4555e} /* (21, 14, 12) {real, imag} */,
  {32'hbe928860, 32'h400384c2} /* (21, 14, 11) {real, imag} */,
  {32'h3e8a8d50, 32'h4062716f} /* (21, 14, 10) {real, imag} */,
  {32'h3df13e00, 32'h3f08d488} /* (21, 14, 9) {real, imag} */,
  {32'h3ff09102, 32'h401f5286} /* (21, 14, 8) {real, imag} */,
  {32'hbe545080, 32'h3e6b92a8} /* (21, 14, 7) {real, imag} */,
  {32'hbe7c2c40, 32'h3f7cabd6} /* (21, 14, 6) {real, imag} */,
  {32'h400dfe5e, 32'h3f7e0ac5} /* (21, 14, 5) {real, imag} */,
  {32'h405a2c2c, 32'hbf4986cc} /* (21, 14, 4) {real, imag} */,
  {32'h3ff8dcde, 32'hbfa28398} /* (21, 14, 3) {real, imag} */,
  {32'h40132e53, 32'h3f652972} /* (21, 14, 2) {real, imag} */,
  {32'h40261ed6, 32'hbe2a382c} /* (21, 14, 1) {real, imag} */,
  {32'h3ff6b74d, 32'hc018b040} /* (21, 14, 0) {real, imag} */,
  {32'h4021eab4, 32'h3c54c000} /* (21, 13, 31) {real, imag} */,
  {32'h4034054e, 32'hbeeb9d50} /* (21, 13, 30) {real, imag} */,
  {32'hc003a42e, 32'hbffd3d84} /* (21, 13, 29) {real, imag} */,
  {32'hc0787a44, 32'h3e829074} /* (21, 13, 28) {real, imag} */,
  {32'hc02144d8, 32'hc01884f0} /* (21, 13, 27) {real, imag} */,
  {32'hbda46240, 32'hbfcc9868} /* (21, 13, 26) {real, imag} */,
  {32'h3ff093a5, 32'h3fe6bf68} /* (21, 13, 25) {real, imag} */,
  {32'h3fd32604, 32'h401ebada} /* (21, 13, 24) {real, imag} */,
  {32'h40597b49, 32'hbf91e854} /* (21, 13, 23) {real, imag} */,
  {32'h403f0c93, 32'hc0ad4f63} /* (21, 13, 22) {real, imag} */,
  {32'hbfb3e312, 32'hbfb8168a} /* (21, 13, 21) {real, imag} */,
  {32'hc0422ad6, 32'h3fb5f0fa} /* (21, 13, 20) {real, imag} */,
  {32'hc006890a, 32'hbf91d888} /* (21, 13, 19) {real, imag} */,
  {32'hc0124ac8, 32'hbffb5a20} /* (21, 13, 18) {real, imag} */,
  {32'h3fae1a4a, 32'h4001e358} /* (21, 13, 17) {real, imag} */,
  {32'h3fb4265e, 32'hbfce7449} /* (21, 13, 16) {real, imag} */,
  {32'hbfa546e9, 32'hbf8f0aec} /* (21, 13, 15) {real, imag} */,
  {32'hbeef4dfc, 32'h401453ba} /* (21, 13, 14) {real, imag} */,
  {32'h3fc638b0, 32'h3fa5bdba} /* (21, 13, 13) {real, imag} */,
  {32'h3f4cd350, 32'hbef0f8d6} /* (21, 13, 12) {real, imag} */,
  {32'hbf660c8c, 32'hc0006c90} /* (21, 13, 11) {real, imag} */,
  {32'hc0516e46, 32'h3fb4e042} /* (21, 13, 10) {real, imag} */,
  {32'hc088b7a0, 32'h3fbb0aca} /* (21, 13, 9) {real, imag} */,
  {32'hbd3a1b60, 32'h3fe5d6a5} /* (21, 13, 8) {real, imag} */,
  {32'hbe46bee0, 32'h3f90edd0} /* (21, 13, 7) {real, imag} */,
  {32'hbfd5cdd3, 32'h3f6e7df8} /* (21, 13, 6) {real, imag} */,
  {32'h3eb74610, 32'h3f20e556} /* (21, 13, 5) {real, imag} */,
  {32'h3fdb7b22, 32'h403c01ec} /* (21, 13, 4) {real, imag} */,
  {32'hbf40a490, 32'h409bfee8} /* (21, 13, 3) {real, imag} */,
  {32'h3f015942, 32'h40a7a609} /* (21, 13, 2) {real, imag} */,
  {32'h4061111e, 32'h3f4237ae} /* (21, 13, 1) {real, imag} */,
  {32'h40389ef4, 32'h3f00f516} /* (21, 13, 0) {real, imag} */,
  {32'h3f86be60, 32'h3f14b0a0} /* (21, 12, 31) {real, imag} */,
  {32'h4038d8d3, 32'h3fbe1e3b} /* (21, 12, 30) {real, imag} */,
  {32'hc02537f6, 32'hbe853c12} /* (21, 12, 29) {real, imag} */,
  {32'hc02a5c4a, 32'h3e881380} /* (21, 12, 28) {real, imag} */,
  {32'hc0280ca6, 32'h4031a8d8} /* (21, 12, 27) {real, imag} */,
  {32'hc083abde, 32'hbf55ea44} /* (21, 12, 26) {real, imag} */,
  {32'hbf86522b, 32'hbf9830fe} /* (21, 12, 25) {real, imag} */,
  {32'h3ffc65bb, 32'h3f5e77f5} /* (21, 12, 24) {real, imag} */,
  {32'hbe38c530, 32'hc02ee588} /* (21, 12, 23) {real, imag} */,
  {32'hc03c3c30, 32'h3fb44c8e} /* (21, 12, 22) {real, imag} */,
  {32'hc004916f, 32'h40bc55de} /* (21, 12, 21) {real, imag} */,
  {32'hbeba6c3c, 32'h3fcffaf2} /* (21, 12, 20) {real, imag} */,
  {32'hbefc9478, 32'hc00eb0dd} /* (21, 12, 19) {real, imag} */,
  {32'hbd60c740, 32'h4030c82c} /* (21, 12, 18) {real, imag} */,
  {32'hc0526db6, 32'hbf62dd18} /* (21, 12, 17) {real, imag} */,
  {32'hc08ccade, 32'hbf6866ac} /* (21, 12, 16) {real, imag} */,
  {32'hbe8b24e0, 32'h3fd5c1af} /* (21, 12, 15) {real, imag} */,
  {32'h3f02cbec, 32'h3f8b3095} /* (21, 12, 14) {real, imag} */,
  {32'h4001f238, 32'hbf5e1ea2} /* (21, 12, 13) {real, imag} */,
  {32'h3fa6a929, 32'hc0b04215} /* (21, 12, 12) {real, imag} */,
  {32'h3f2625ee, 32'hc01c91fb} /* (21, 12, 11) {real, imag} */,
  {32'h3f53b335, 32'h3f96e283} /* (21, 12, 10) {real, imag} */,
  {32'h3e8cdbf0, 32'h408fb48b} /* (21, 12, 9) {real, imag} */,
  {32'hc0108e06, 32'h40513aac} /* (21, 12, 8) {real, imag} */,
  {32'hc0664506, 32'h3f01d388} /* (21, 12, 7) {real, imag} */,
  {32'hbf9a2ef5, 32'h3fc9a89e} /* (21, 12, 6) {real, imag} */,
  {32'h4072fe9d, 32'h4078d72b} /* (21, 12, 5) {real, imag} */,
  {32'hc01a7f0b, 32'h3f5e2b4d} /* (21, 12, 4) {real, imag} */,
  {32'hbf2a83ea, 32'h3f4b9abc} /* (21, 12, 3) {real, imag} */,
  {32'hbf30bef8, 32'h4032cc3d} /* (21, 12, 2) {real, imag} */,
  {32'hbfeba18b, 32'hc00e5b09} /* (21, 12, 1) {real, imag} */,
  {32'hc004a40f, 32'hbf9563b4} /* (21, 12, 0) {real, imag} */,
  {32'h3cb135c0, 32'hbe88d8e8} /* (21, 11, 31) {real, imag} */,
  {32'h3f041164, 32'hbf9e4645} /* (21, 11, 30) {real, imag} */,
  {32'hbf1c7455, 32'hc01a7990} /* (21, 11, 29) {real, imag} */,
  {32'hbfb55d1c, 32'h3eabda10} /* (21, 11, 28) {real, imag} */,
  {32'h3e085360, 32'h3e7a8250} /* (21, 11, 27) {real, imag} */,
  {32'hbfa06914, 32'hc0a94fd2} /* (21, 11, 26) {real, imag} */,
  {32'hc0c33120, 32'hc0ab2a6a} /* (21, 11, 25) {real, imag} */,
  {32'hc0ecc271, 32'h400d49f9} /* (21, 11, 24) {real, imag} */,
  {32'hbfd0379a, 32'h4117b28a} /* (21, 11, 23) {real, imag} */,
  {32'h3f14f21e, 32'h40d7f9e4} /* (21, 11, 22) {real, imag} */,
  {32'hc00b855b, 32'h4019c916} /* (21, 11, 21) {real, imag} */,
  {32'hc0c57f14, 32'h3fd3b351} /* (21, 11, 20) {real, imag} */,
  {32'hbf54ecda, 32'h3fab3d49} /* (21, 11, 19) {real, imag} */,
  {32'h406795da, 32'hbeeaab70} /* (21, 11, 18) {real, imag} */,
  {32'h3fd6d988, 32'h3ff0b1f2} /* (21, 11, 17) {real, imag} */,
  {32'hc077b5a0, 32'hbe3fbbb0} /* (21, 11, 16) {real, imag} */,
  {32'hbf8166ba, 32'h4032ab70} /* (21, 11, 15) {real, imag} */,
  {32'h3db9c0b0, 32'h402c5593} /* (21, 11, 14) {real, imag} */,
  {32'hbf2a8c3c, 32'h40a4661c} /* (21, 11, 13) {real, imag} */,
  {32'hc00e5592, 32'h40dc1adc} /* (21, 11, 12) {real, imag} */,
  {32'hc00c7192, 32'h3fce5b43} /* (21, 11, 11) {real, imag} */,
  {32'hbfe8c76a, 32'h3f0387d8} /* (21, 11, 10) {real, imag} */,
  {32'hc04e4845, 32'hc028a6cc} /* (21, 11, 9) {real, imag} */,
  {32'hbf9acd98, 32'hc0ae32fe} /* (21, 11, 8) {real, imag} */,
  {32'h3fef62ee, 32'hc0b0c1f8} /* (21, 11, 7) {real, imag} */,
  {32'hc00516c5, 32'hc08e12b1} /* (21, 11, 6) {real, imag} */,
  {32'h3f72e940, 32'hc092e97f} /* (21, 11, 5) {real, imag} */,
  {32'hbf2c9b16, 32'hc0034224} /* (21, 11, 4) {real, imag} */,
  {32'hbfe5016c, 32'hc030f91a} /* (21, 11, 3) {real, imag} */,
  {32'hc07bb16a, 32'hc04f5ac3} /* (21, 11, 2) {real, imag} */,
  {32'hc004bfc1, 32'hbf49b74c} /* (21, 11, 1) {real, imag} */,
  {32'hbfcb962e, 32'hbf36dd28} /* (21, 11, 0) {real, imag} */,
  {32'hc00a3514, 32'h3fb0e04c} /* (21, 10, 31) {real, imag} */,
  {32'hc0c24185, 32'h3ffac538} /* (21, 10, 30) {real, imag} */,
  {32'h400ee4c4, 32'h40970820} /* (21, 10, 29) {real, imag} */,
  {32'h4081722d, 32'h408e0886} /* (21, 10, 28) {real, imag} */,
  {32'h40df6a0b, 32'hbff4d4a0} /* (21, 10, 27) {real, imag} */,
  {32'h4052969a, 32'h3f07abc4} /* (21, 10, 26) {real, imag} */,
  {32'hbf835e1f, 32'hc0526c8a} /* (21, 10, 25) {real, imag} */,
  {32'hc0ba4229, 32'hc08347eb} /* (21, 10, 24) {real, imag} */,
  {32'h406ba52a, 32'hc005d928} /* (21, 10, 23) {real, imag} */,
  {32'h4003d653, 32'hbf889a66} /* (21, 10, 22) {real, imag} */,
  {32'h3e92240c, 32'h3f8f8d0b} /* (21, 10, 21) {real, imag} */,
  {32'h408fdc60, 32'hc0043b56} /* (21, 10, 20) {real, imag} */,
  {32'h401ea696, 32'h3eae8e80} /* (21, 10, 19) {real, imag} */,
  {32'hbff72afd, 32'hc030ed16} /* (21, 10, 18) {real, imag} */,
  {32'hc092e821, 32'hc06ae60d} /* (21, 10, 17) {real, imag} */,
  {32'h3f072b86, 32'hc0198b4a} /* (21, 10, 16) {real, imag} */,
  {32'h4019b68e, 32'hbee39e70} /* (21, 10, 15) {real, imag} */,
  {32'hbfae0d08, 32'h40702bc6} /* (21, 10, 14) {real, imag} */,
  {32'hc022bda7, 32'hc04c1e1c} /* (21, 10, 13) {real, imag} */,
  {32'h408b0fb0, 32'hc02930ba} /* (21, 10, 12) {real, imag} */,
  {32'h404f1d54, 32'hc0d0e886} /* (21, 10, 11) {real, imag} */,
  {32'hc0b21194, 32'hc0801cdd} /* (21, 10, 10) {real, imag} */,
  {32'h3dfa2f20, 32'h3f9b7f58} /* (21, 10, 9) {real, imag} */,
  {32'hbf601140, 32'h401021ae} /* (21, 10, 8) {real, imag} */,
  {32'hc0a7471c, 32'hbf8cc370} /* (21, 10, 7) {real, imag} */,
  {32'hc0a4c5a4, 32'h3fdc6043} /* (21, 10, 6) {real, imag} */,
  {32'h3ff9696a, 32'h3f690888} /* (21, 10, 5) {real, imag} */,
  {32'h409f833f, 32'hc05d8dc0} /* (21, 10, 4) {real, imag} */,
  {32'hc081335d, 32'h4089222b} /* (21, 10, 3) {real, imag} */,
  {32'hbf979ef8, 32'h4076b144} /* (21, 10, 2) {real, imag} */,
  {32'h3fefbf81, 32'h3fab8a3c} /* (21, 10, 1) {real, imag} */,
  {32'h400df880, 32'hbfcf4745} /* (21, 10, 0) {real, imag} */,
  {32'hc02e71de, 32'h3e84d9c8} /* (21, 9, 31) {real, imag} */,
  {32'hc091eb70, 32'hbffb19e8} /* (21, 9, 30) {real, imag} */,
  {32'h3e2772a4, 32'hc04f420b} /* (21, 9, 29) {real, imag} */,
  {32'h404dd82b, 32'hc0a131bc} /* (21, 9, 28) {real, imag} */,
  {32'h3e9554c0, 32'h40316026} /* (21, 9, 27) {real, imag} */,
  {32'hbf9cddec, 32'h40f04380} /* (21, 9, 26) {real, imag} */,
  {32'h3fa58c2b, 32'h4087cd09} /* (21, 9, 25) {real, imag} */,
  {32'h3f82611f, 32'h3f6f94e0} /* (21, 9, 24) {real, imag} */,
  {32'hbfe3ffb4, 32'h3f01aad4} /* (21, 9, 23) {real, imag} */,
  {32'h40cd4c98, 32'h400add85} /* (21, 9, 22) {real, imag} */,
  {32'h4126d078, 32'hbfc7d6bc} /* (21, 9, 21) {real, imag} */,
  {32'h40a70fda, 32'hc0150068} /* (21, 9, 20) {real, imag} */,
  {32'h3ff86694, 32'hc08cb4bc} /* (21, 9, 19) {real, imag} */,
  {32'hc0305b2a, 32'hc00e99c7} /* (21, 9, 18) {real, imag} */,
  {32'hc03d2237, 32'h402298f5} /* (21, 9, 17) {real, imag} */,
  {32'h40207eb9, 32'hbe5d2092} /* (21, 9, 16) {real, imag} */,
  {32'hbea07760, 32'hbe51d6d0} /* (21, 9, 15) {real, imag} */,
  {32'hc0caee3f, 32'h40952ccb} /* (21, 9, 14) {real, imag} */,
  {32'hc0d9afd0, 32'h409c3d3f} /* (21, 9, 13) {real, imag} */,
  {32'hbf95b9fe, 32'h4007e3b0} /* (21, 9, 12) {real, imag} */,
  {32'h400d17b2, 32'h40950c4a} /* (21, 9, 11) {real, imag} */,
  {32'h40e1efe0, 32'hbe94e618} /* (21, 9, 10) {real, imag} */,
  {32'h40aea8a9, 32'hbf82606b} /* (21, 9, 9) {real, imag} */,
  {32'h404b7e0a, 32'h400b7d95} /* (21, 9, 8) {real, imag} */,
  {32'h4035f0f2, 32'h40d4ce6e} /* (21, 9, 7) {real, imag} */,
  {32'h400ecc0d, 32'h4044ac88} /* (21, 9, 6) {real, imag} */,
  {32'hc01ad9a4, 32'hbf790678} /* (21, 9, 5) {real, imag} */,
  {32'h408c10ce, 32'hc01d42a7} /* (21, 9, 4) {real, imag} */,
  {32'h400a08f2, 32'hbfc35684} /* (21, 9, 3) {real, imag} */,
  {32'hc0d1b0eb, 32'hbfadb872} /* (21, 9, 2) {real, imag} */,
  {32'hc0bd6deb, 32'hc048cc76} /* (21, 9, 1) {real, imag} */,
  {32'hc0035e78, 32'hc009f089} /* (21, 9, 0) {real, imag} */,
  {32'h40702827, 32'hbef9bdc8} /* (21, 8, 31) {real, imag} */,
  {32'h3f13ce04, 32'hbe508c10} /* (21, 8, 30) {real, imag} */,
  {32'hc108a282, 32'hc0b16834} /* (21, 8, 29) {real, imag} */,
  {32'hc0d6db50, 32'hc0fd14be} /* (21, 8, 28) {real, imag} */,
  {32'h3fcda112, 32'h40b02de3} /* (21, 8, 27) {real, imag} */,
  {32'h406f4cde, 32'h403808f9} /* (21, 8, 26) {real, imag} */,
  {32'h3f865f17, 32'hbf9c6f68} /* (21, 8, 25) {real, imag} */,
  {32'hbfcc6178, 32'hc04bae42} /* (21, 8, 24) {real, imag} */,
  {32'hc01e1fbc, 32'hc03acc11} /* (21, 8, 23) {real, imag} */,
  {32'h405c89ca, 32'hc080e2a5} /* (21, 8, 22) {real, imag} */,
  {32'hc012677c, 32'h3e2647b0} /* (21, 8, 21) {real, imag} */,
  {32'hbf3d87da, 32'h3f6147fc} /* (21, 8, 20) {real, imag} */,
  {32'h3fa2c828, 32'hc071b600} /* (21, 8, 19) {real, imag} */,
  {32'h405ee1c7, 32'hc133c980} /* (21, 8, 18) {real, imag} */,
  {32'h40bb6d6e, 32'hc12dc796} /* (21, 8, 17) {real, imag} */,
  {32'h3e493f88, 32'hc0a4ccb8} /* (21, 8, 16) {real, imag} */,
  {32'hc0d2175b, 32'h40534506} /* (21, 8, 15) {real, imag} */,
  {32'hc0f0b7e8, 32'h40101c5e} /* (21, 8, 14) {real, imag} */,
  {32'hbd2ef680, 32'h4027934a} /* (21, 8, 13) {real, imag} */,
  {32'h406f017c, 32'h4059c672} /* (21, 8, 12) {real, imag} */,
  {32'hc02ac672, 32'h403b4e0f} /* (21, 8, 11) {real, imag} */,
  {32'h3f231606, 32'h3e8b2bf8} /* (21, 8, 10) {real, imag} */,
  {32'h3f6450fc, 32'h3ffcb246} /* (21, 8, 9) {real, imag} */,
  {32'hc031faa8, 32'h406defa5} /* (21, 8, 8) {real, imag} */,
  {32'hc0a2f644, 32'hc036cb17} /* (21, 8, 7) {real, imag} */,
  {32'hc0b9ef43, 32'hc136a4be} /* (21, 8, 6) {real, imag} */,
  {32'hc0e59640, 32'hc086b171} /* (21, 8, 5) {real, imag} */,
  {32'hc0dea6d8, 32'hbf8d2d77} /* (21, 8, 4) {real, imag} */,
  {32'hc100f506, 32'hc0d08fc4} /* (21, 8, 3) {real, imag} */,
  {32'hc02e050b, 32'hc11ccc76} /* (21, 8, 2) {real, imag} */,
  {32'hc06d20c8, 32'hc11d83fb} /* (21, 8, 1) {real, imag} */,
  {32'hbf4a82b2, 32'hc080dd7d} /* (21, 8, 0) {real, imag} */,
  {32'hc0340779, 32'h4096f8fe} /* (21, 7, 31) {real, imag} */,
  {32'hc002570e, 32'hbedbd2d8} /* (21, 7, 30) {real, imag} */,
  {32'h40ce4774, 32'hc0369b70} /* (21, 7, 29) {real, imag} */,
  {32'h3f9e6536, 32'hc0767264} /* (21, 7, 28) {real, imag} */,
  {32'hbf3fdae0, 32'hc02f8bae} /* (21, 7, 27) {real, imag} */,
  {32'hbea4131c, 32'hbfdaab84} /* (21, 7, 26) {real, imag} */,
  {32'hbf5571e6, 32'h3f9a84f8} /* (21, 7, 25) {real, imag} */,
  {32'h40a9095c, 32'hc0d6eea9} /* (21, 7, 24) {real, imag} */,
  {32'h40d07418, 32'hc12b776c} /* (21, 7, 23) {real, imag} */,
  {32'h3da37180, 32'hc05fc1fb} /* (21, 7, 22) {real, imag} */,
  {32'h3e0a6338, 32'hc08d0f3a} /* (21, 7, 21) {real, imag} */,
  {32'h406c5e02, 32'hbfb3535f} /* (21, 7, 20) {real, imag} */,
  {32'hbe629140, 32'hbfe6fe94} /* (21, 7, 19) {real, imag} */,
  {32'h3e953420, 32'h4044153d} /* (21, 7, 18) {real, imag} */,
  {32'h40b26600, 32'hbf80b8c2} /* (21, 7, 17) {real, imag} */,
  {32'h4078d146, 32'h404da466} /* (21, 7, 16) {real, imag} */,
  {32'h3e047400, 32'h3fe4ef01} /* (21, 7, 15) {real, imag} */,
  {32'h3f4afb2e, 32'h3fd9fac6} /* (21, 7, 14) {real, imag} */,
  {32'h41208371, 32'h3f4350e0} /* (21, 7, 13) {real, imag} */,
  {32'h3febb216, 32'h405c066e} /* (21, 7, 12) {real, imag} */,
  {32'hc0b1cdeb, 32'h4042a4cf} /* (21, 7, 11) {real, imag} */,
  {32'hc05e6270, 32'hc0a16b54} /* (21, 7, 10) {real, imag} */,
  {32'hc02e1c48, 32'hc0ba7b42} /* (21, 7, 9) {real, imag} */,
  {32'h41086095, 32'hc04ad031} /* (21, 7, 8) {real, imag} */,
  {32'h40b7a485, 32'h4066a905} /* (21, 7, 7) {real, imag} */,
  {32'h3fef4c5c, 32'h40ac5249} /* (21, 7, 6) {real, imag} */,
  {32'h3fb2d782, 32'h40604f80} /* (21, 7, 5) {real, imag} */,
  {32'h3f1660b8, 32'hbff933be} /* (21, 7, 4) {real, imag} */,
  {32'h3fb59564, 32'h3e20d890} /* (21, 7, 3) {real, imag} */,
  {32'h40df899d, 32'hc0a1cef1} /* (21, 7, 2) {real, imag} */,
  {32'h40980c3c, 32'hc0034e4b} /* (21, 7, 1) {real, imag} */,
  {32'h3d92ea10, 32'h400a2949} /* (21, 7, 0) {real, imag} */,
  {32'hc01e4faa, 32'h3fcd3a08} /* (21, 6, 31) {real, imag} */,
  {32'hc10388cc, 32'hc09d0424} /* (21, 6, 30) {real, imag} */,
  {32'hbfa57744, 32'hc090e433} /* (21, 6, 29) {real, imag} */,
  {32'h410d6534, 32'h40cb4cb8} /* (21, 6, 28) {real, imag} */,
  {32'h412e482f, 32'h411b8ecd} /* (21, 6, 27) {real, imag} */,
  {32'h4113a0f5, 32'hbfdba798} /* (21, 6, 26) {real, imag} */,
  {32'h412e6ff8, 32'hc0cc5bb5} /* (21, 6, 25) {real, imag} */,
  {32'h40f07970, 32'hc084317c} /* (21, 6, 24) {real, imag} */,
  {32'h3e6771e0, 32'hc1403c51} /* (21, 6, 23) {real, imag} */,
  {32'h40771da7, 32'hc17f264a} /* (21, 6, 22) {real, imag} */,
  {32'h4090a356, 32'hc0bb2189} /* (21, 6, 21) {real, imag} */,
  {32'hc07ed2ec, 32'hbeb549fe} /* (21, 6, 20) {real, imag} */,
  {32'hc0e963a1, 32'hbf9a47d0} /* (21, 6, 19) {real, imag} */,
  {32'h3fc0c042, 32'h3f911c7c} /* (21, 6, 18) {real, imag} */,
  {32'h40d6bc3c, 32'hc072389f} /* (21, 6, 17) {real, imag} */,
  {32'h3fc54d48, 32'h40c381a0} /* (21, 6, 16) {real, imag} */,
  {32'h3d42a700, 32'h40533a9c} /* (21, 6, 15) {real, imag} */,
  {32'h3eab5a88, 32'h40499d4a} /* (21, 6, 14) {real, imag} */,
  {32'hbebbc6a0, 32'h3ffd6a69} /* (21, 6, 13) {real, imag} */,
  {32'hc018a9f6, 32'hc0a0a35a} /* (21, 6, 12) {real, imag} */,
  {32'hbf290fe0, 32'hc00f6559} /* (21, 6, 11) {real, imag} */,
  {32'h405522b2, 32'hc00263f8} /* (21, 6, 10) {real, imag} */,
  {32'h40de5bfe, 32'hbfab4638} /* (21, 6, 9) {real, imag} */,
  {32'hbecea948, 32'hc126b7c3} /* (21, 6, 8) {real, imag} */,
  {32'hbfc684ca, 32'h3f50f864} /* (21, 6, 7) {real, imag} */,
  {32'hbf63b7a4, 32'hc09ba855} /* (21, 6, 6) {real, imag} */,
  {32'hbff41176, 32'hc02adf4b} /* (21, 6, 5) {real, imag} */,
  {32'hbebb2050, 32'h3ef693a0} /* (21, 6, 4) {real, imag} */,
  {32'h3fd300d6, 32'hbfb9389c} /* (21, 6, 3) {real, imag} */,
  {32'hc087c0c9, 32'h4090e885} /* (21, 6, 2) {real, imag} */,
  {32'hbf7f1a5e, 32'h405a690c} /* (21, 6, 1) {real, imag} */,
  {32'h3fa10a2e, 32'h40044299} /* (21, 6, 0) {real, imag} */,
  {32'hc0bcff19, 32'hbf861afc} /* (21, 5, 31) {real, imag} */,
  {32'hc0eb2ef5, 32'hc02aca96} /* (21, 5, 30) {real, imag} */,
  {32'hc134157c, 32'hbfad2180} /* (21, 5, 29) {real, imag} */,
  {32'hc0d8a872, 32'hc064d21f} /* (21, 5, 28) {real, imag} */,
  {32'hc0fdf47b, 32'hc07d5ffb} /* (21, 5, 27) {real, imag} */,
  {32'hc03bbe20, 32'hbfca4a0e} /* (21, 5, 26) {real, imag} */,
  {32'h3f04d898, 32'hc10821b2} /* (21, 5, 25) {real, imag} */,
  {32'hc0882e06, 32'hc136cc97} /* (21, 5, 24) {real, imag} */,
  {32'hc169f3be, 32'hc14ca8ca} /* (21, 5, 23) {real, imag} */,
  {32'hc0578c54, 32'hc1031441} /* (21, 5, 22) {real, imag} */,
  {32'h40c46fe6, 32'hc10dd288} /* (21, 5, 21) {real, imag} */,
  {32'h40e8668e, 32'h400ad860} /* (21, 5, 20) {real, imag} */,
  {32'h4035a95a, 32'h40afd7f7} /* (21, 5, 19) {real, imag} */,
  {32'h3ff28be6, 32'h3fe6b636} /* (21, 5, 18) {real, imag} */,
  {32'h40113a9e, 32'hbfd05fc2} /* (21, 5, 17) {real, imag} */,
  {32'hc06d800e, 32'h401cbc2a} /* (21, 5, 16) {real, imag} */,
  {32'hc0d67b92, 32'h409adcd6} /* (21, 5, 15) {real, imag} */,
  {32'hc083faf7, 32'h410a98a5} /* (21, 5, 14) {real, imag} */,
  {32'h3fa8139e, 32'h41177789} /* (21, 5, 13) {real, imag} */,
  {32'h3f9f03f0, 32'hc04c6273} /* (21, 5, 12) {real, imag} */,
  {32'hc0f12cd2, 32'hc12e476c} /* (21, 5, 11) {real, imag} */,
  {32'hc116aaef, 32'hbf403e38} /* (21, 5, 10) {real, imag} */,
  {32'h404ce9a1, 32'h3dfe5380} /* (21, 5, 9) {real, imag} */,
  {32'h414b8a36, 32'hc08b3aa2} /* (21, 5, 8) {real, imag} */,
  {32'h41079499, 32'hc06423c4} /* (21, 5, 7) {real, imag} */,
  {32'hc0306da5, 32'hc17b95fd} /* (21, 5, 6) {real, imag} */,
  {32'hbd49b5c0, 32'hc16e587c} /* (21, 5, 5) {real, imag} */,
  {32'h4092c06f, 32'hc1425d02} /* (21, 5, 4) {real, imag} */,
  {32'h401c6f24, 32'hc09934b9} /* (21, 5, 3) {real, imag} */,
  {32'hc08e1933, 32'hbf8dbaea} /* (21, 5, 2) {real, imag} */,
  {32'hc0a71bb8, 32'h4093888e} /* (21, 5, 1) {real, imag} */,
  {32'hbf091f44, 32'h3e9c7a78} /* (21, 5, 0) {real, imag} */,
  {32'h40aec1cc, 32'h4023fcc6} /* (21, 4, 31) {real, imag} */,
  {32'h405d556c, 32'hc093561b} /* (21, 4, 30) {real, imag} */,
  {32'h3f3ff2c8, 32'hc0d0d005} /* (21, 4, 29) {real, imag} */,
  {32'hbfb14083, 32'hc137a60c} /* (21, 4, 28) {real, imag} */,
  {32'hbf036674, 32'hc1586d90} /* (21, 4, 27) {real, imag} */,
  {32'h40bb8c64, 32'hc0e5d65a} /* (21, 4, 26) {real, imag} */,
  {32'h40042030, 32'hc15734d8} /* (21, 4, 25) {real, imag} */,
  {32'h4053ff34, 32'hc15b668b} /* (21, 4, 24) {real, imag} */,
  {32'h3e12b580, 32'h4119550e} /* (21, 4, 23) {real, imag} */,
  {32'h3fb6758e, 32'h414778fc} /* (21, 4, 22) {real, imag} */,
  {32'hc007ea22, 32'h4128d3aa} /* (21, 4, 21) {real, imag} */,
  {32'hc0ba6f28, 32'h403cabda} /* (21, 4, 20) {real, imag} */,
  {32'hc042ed1b, 32'h40fae54e} /* (21, 4, 19) {real, imag} */,
  {32'hc0738240, 32'h40d1f61f} /* (21, 4, 18) {real, imag} */,
  {32'hc09494fb, 32'h3fa90a38} /* (21, 4, 17) {real, imag} */,
  {32'hc0849fa6, 32'hc0fcac7a} /* (21, 4, 16) {real, imag} */,
  {32'hc01e2d4e, 32'hc0d6416a} /* (21, 4, 15) {real, imag} */,
  {32'h40934fc0, 32'hc1033356} /* (21, 4, 14) {real, imag} */,
  {32'h401e46e0, 32'hc0082b2c} /* (21, 4, 13) {real, imag} */,
  {32'h40bb1f70, 32'hc009679c} /* (21, 4, 12) {real, imag} */,
  {32'h3fcdefd5, 32'h40b471e8} /* (21, 4, 11) {real, imag} */,
  {32'h40bbad8e, 32'h40da28ba} /* (21, 4, 10) {real, imag} */,
  {32'hc038e65c, 32'h3fdc79ea} /* (21, 4, 9) {real, imag} */,
  {32'hc15f2d40, 32'h40a0639e} /* (21, 4, 8) {real, imag} */,
  {32'hc12664ab, 32'h40896bec} /* (21, 4, 7) {real, imag} */,
  {32'h40859b38, 32'h403c7958} /* (21, 4, 6) {real, imag} */,
  {32'h4078a42d, 32'h3fca4e48} /* (21, 4, 5) {real, imag} */,
  {32'hc06b0a2c, 32'hbfd8b20e} /* (21, 4, 4) {real, imag} */,
  {32'hbf238166, 32'hbf94e346} /* (21, 4, 3) {real, imag} */,
  {32'h40829dbe, 32'hbfb4073f} /* (21, 4, 2) {real, imag} */,
  {32'h407f1f48, 32'h412e9407} /* (21, 4, 1) {real, imag} */,
  {32'h40497772, 32'h411c37a1} /* (21, 4, 0) {real, imag} */,
  {32'h40be7f44, 32'hc0ce6a7b} /* (21, 3, 31) {real, imag} */,
  {32'h4078140a, 32'hc03c456a} /* (21, 3, 30) {real, imag} */,
  {32'hbf17a7c1, 32'hc089ad65} /* (21, 3, 29) {real, imag} */,
  {32'hbfb0bafc, 32'hc0c55b12} /* (21, 3, 28) {real, imag} */,
  {32'h4009c984, 32'hc0343bda} /* (21, 3, 27) {real, imag} */,
  {32'h40c21664, 32'h41417587} /* (21, 3, 26) {real, imag} */,
  {32'h4055f81e, 32'h40a1b5c5} /* (21, 3, 25) {real, imag} */,
  {32'hc02c5865, 32'h3d9990a0} /* (21, 3, 24) {real, imag} */,
  {32'hbec269c0, 32'hc01e6806} /* (21, 3, 23) {real, imag} */,
  {32'h406b60db, 32'h4095b5af} /* (21, 3, 22) {real, imag} */,
  {32'hc041d7c4, 32'h40a9664d} /* (21, 3, 21) {real, imag} */,
  {32'h4079fa3c, 32'hc0fb9e63} /* (21, 3, 20) {real, imag} */,
  {32'h402a0ea0, 32'hc0cebc1a} /* (21, 3, 19) {real, imag} */,
  {32'h40953fe3, 32'hc0f62174} /* (21, 3, 18) {real, imag} */,
  {32'h4091cc12, 32'hc12dee12} /* (21, 3, 17) {real, imag} */,
  {32'h3f8b930c, 32'hc11f63bd} /* (21, 3, 16) {real, imag} */,
  {32'hc077cdb5, 32'hc145cc74} /* (21, 3, 15) {real, imag} */,
  {32'hbfca35c0, 32'hc1497db5} /* (21, 3, 14) {real, imag} */,
  {32'h41310cff, 32'hc16f2423} /* (21, 3, 13) {real, imag} */,
  {32'h409776fa, 32'hc02cbd01} /* (21, 3, 12) {real, imag} */,
  {32'hc132c205, 32'hbff85244} /* (21, 3, 11) {real, imag} */,
  {32'h3f7b76a8, 32'h3f353e60} /* (21, 3, 10) {real, imag} */,
  {32'hc08c20a0, 32'hbfb076be} /* (21, 3, 9) {real, imag} */,
  {32'hc027f83a, 32'h415cd4df} /* (21, 3, 8) {real, imag} */,
  {32'h3f8daf30, 32'h41852fa0} /* (21, 3, 7) {real, imag} */,
  {32'h4084f537, 32'h41860317} /* (21, 3, 6) {real, imag} */,
  {32'hc02fb21b, 32'h4045d9b3} /* (21, 3, 5) {real, imag} */,
  {32'hc0eee958, 32'hc0d34353} /* (21, 3, 4) {real, imag} */,
  {32'hc0b78959, 32'hc0b6912e} /* (21, 3, 3) {real, imag} */,
  {32'hbef760fc, 32'h40c00517} /* (21, 3, 2) {real, imag} */,
  {32'hbe2c8920, 32'hbff5c446} /* (21, 3, 1) {real, imag} */,
  {32'h4093859d, 32'hbf3264dc} /* (21, 3, 0) {real, imag} */,
  {32'hbecb1040, 32'hc136e077} /* (21, 2, 31) {real, imag} */,
  {32'hc0a46239, 32'hc156f001} /* (21, 2, 30) {real, imag} */,
  {32'hc1140710, 32'hc1650baf} /* (21, 2, 29) {real, imag} */,
  {32'hc0c00283, 32'hc1350b53} /* (21, 2, 28) {real, imag} */,
  {32'hc0dceb64, 32'hc04f5440} /* (21, 2, 27) {real, imag} */,
  {32'hc0bd776c, 32'hbfdf8c2d} /* (21, 2, 26) {real, imag} */,
  {32'hc0fd9f8c, 32'hc13d3a10} /* (21, 2, 25) {real, imag} */,
  {32'hc14a5f5d, 32'hc14baa85} /* (21, 2, 24) {real, imag} */,
  {32'hc125c144, 32'hc0f16801} /* (21, 2, 23) {real, imag} */,
  {32'hc1271da6, 32'hc1128198} /* (21, 2, 22) {real, imag} */,
  {32'hc1172f6c, 32'hc1158c1b} /* (21, 2, 21) {real, imag} */,
  {32'h414b470e, 32'hc0e2edba} /* (21, 2, 20) {real, imag} */,
  {32'h4169d941, 32'hc01acfe8} /* (21, 2, 19) {real, imag} */,
  {32'h41949b31, 32'h4017dcc0} /* (21, 2, 18) {real, imag} */,
  {32'h41b9cdb0, 32'h41033a85} /* (21, 2, 17) {real, imag} */,
  {32'h41aba84e, 32'h4091d42f} /* (21, 2, 16) {real, imag} */,
  {32'h418a5f60, 32'hbf839691} /* (21, 2, 15) {real, imag} */,
  {32'h40b71648, 32'h3fe8efaa} /* (21, 2, 14) {real, imag} */,
  {32'h409f5325, 32'h3dd0c810} /* (21, 2, 13) {real, imag} */,
  {32'hc113139f, 32'h4132d5ac} /* (21, 2, 12) {real, imag} */,
  {32'hc1290502, 32'h417eac26} /* (21, 2, 11) {real, imag} */,
  {32'hc0229b88, 32'hc02f347c} /* (21, 2, 10) {real, imag} */,
  {32'h3ee2e880, 32'h3ccfc000} /* (21, 2, 9) {real, imag} */,
  {32'hc0cfa109, 32'hc08dd1ca} /* (21, 2, 8) {real, imag} */,
  {32'hc0f585c2, 32'hc10297ee} /* (21, 2, 7) {real, imag} */,
  {32'hc181050c, 32'hc112fb8a} /* (21, 2, 6) {real, imag} */,
  {32'hc0d3f408, 32'hc0cd27ab} /* (21, 2, 5) {real, imag} */,
  {32'h40b9e819, 32'hc020021e} /* (21, 2, 4) {real, imag} */,
  {32'hbe3646b0, 32'hc0a673cd} /* (21, 2, 3) {real, imag} */,
  {32'hc0f79dad, 32'hc1170e19} /* (21, 2, 2) {real, imag} */,
  {32'hc10b3bf8, 32'h40c43312} /* (21, 2, 1) {real, imag} */,
  {32'h4020d9c2, 32'h40670c45} /* (21, 2, 0) {real, imag} */,
  {32'h4116738e, 32'h4123975b} /* (21, 1, 31) {real, imag} */,
  {32'h415aee21, 32'h4137d7b7} /* (21, 1, 30) {real, imag} */,
  {32'hbfb37368, 32'h41194459} /* (21, 1, 29) {real, imag} */,
  {32'h4115429c, 32'h416c40cd} /* (21, 1, 28) {real, imag} */,
  {32'h412bd7f8, 32'h41079620} /* (21, 1, 27) {real, imag} */,
  {32'h40ace5ff, 32'h4019f01e} /* (21, 1, 26) {real, imag} */,
  {32'h40246370, 32'h4193a824} /* (21, 1, 25) {real, imag} */,
  {32'h4168b894, 32'h41dc32b2} /* (21, 1, 24) {real, imag} */,
  {32'h41522d4e, 32'h419567c4} /* (21, 1, 23) {real, imag} */,
  {32'h4146cbf4, 32'h413bef54} /* (21, 1, 22) {real, imag} */,
  {32'h41268bac, 32'h3fad48b0} /* (21, 1, 21) {real, imag} */,
  {32'h40c6c578, 32'hc11c9590} /* (21, 1, 20) {real, imag} */,
  {32'hc08e2f22, 32'hc1269cea} /* (21, 1, 19) {real, imag} */,
  {32'hbf2f5a00, 32'hc137de12} /* (21, 1, 18) {real, imag} */,
  {32'h406592b8, 32'hc0df3ab7} /* (21, 1, 17) {real, imag} */,
  {32'hc123a8c5, 32'hc0fbf00f} /* (21, 1, 16) {real, imag} */,
  {32'hc0f07936, 32'hc05bec65} /* (21, 1, 15) {real, imag} */,
  {32'hc10fc69a, 32'hc01c6971} /* (21, 1, 14) {real, imag} */,
  {32'hbf0551a0, 32'h3f8866f6} /* (21, 1, 13) {real, imag} */,
  {32'hc06fc7c7, 32'hc0131b8c} /* (21, 1, 12) {real, imag} */,
  {32'hbfe7d5b8, 32'hc039b256} /* (21, 1, 11) {real, imag} */,
  {32'h410dafce, 32'h41b8af46} /* (21, 1, 10) {real, imag} */,
  {32'hc0f47920, 32'h4204ae3d} /* (21, 1, 9) {real, imag} */,
  {32'hc16eac16, 32'h41c21050} /* (21, 1, 8) {real, imag} */,
  {32'hc08168da, 32'h41953bd0} /* (21, 1, 7) {real, imag} */,
  {32'h4093f70b, 32'h41b3eff4} /* (21, 1, 6) {real, imag} */,
  {32'h418721e7, 32'h413846f4} /* (21, 1, 5) {real, imag} */,
  {32'h41a86e80, 32'hbe6fbb00} /* (21, 1, 4) {real, imag} */,
  {32'h41542364, 32'h3fbc7990} /* (21, 1, 3) {real, imag} */,
  {32'h3ff8f9c0, 32'hc00d3ff4} /* (21, 1, 2) {real, imag} */,
  {32'h413564dc, 32'h405c266e} /* (21, 1, 1) {real, imag} */,
  {32'h413879c5, 32'h4042cdfe} /* (21, 1, 0) {real, imag} */,
  {32'h40b6af40, 32'h40daf393} /* (21, 0, 31) {real, imag} */,
  {32'h41695b8a, 32'h4197efaa} /* (21, 0, 30) {real, imag} */,
  {32'h410397e6, 32'h40b71338} /* (21, 0, 29) {real, imag} */,
  {32'hc06a048a, 32'hbf6f61c8} /* (21, 0, 28) {real, imag} */,
  {32'hc0c3a028, 32'h40581343} /* (21, 0, 27) {real, imag} */,
  {32'h3ef56242, 32'h405a30bc} /* (21, 0, 26) {real, imag} */,
  {32'h40df2e81, 32'h404d919a} /* (21, 0, 25) {real, imag} */,
  {32'h4170bf0e, 32'hbf52272a} /* (21, 0, 24) {real, imag} */,
  {32'h416fcf63, 32'h40035ea3} /* (21, 0, 23) {real, imag} */,
  {32'h400fc30b, 32'h40b651bc} /* (21, 0, 22) {real, imag} */,
  {32'h407df292, 32'h3f08f7fc} /* (21, 0, 21) {real, imag} */,
  {32'hbf5f08b3, 32'hc1184886} /* (21, 0, 20) {real, imag} */,
  {32'h3f1c5070, 32'hc0783d30} /* (21, 0, 19) {real, imag} */,
  {32'h3e35b4c0, 32'h4150f8aa} /* (21, 0, 18) {real, imag} */,
  {32'hbf002f72, 32'h413415ba} /* (21, 0, 17) {real, imag} */,
  {32'h40e6bfbd, 32'hbd2ab080} /* (21, 0, 16) {real, imag} */,
  {32'hc06e929a, 32'hc1157796} /* (21, 0, 15) {real, imag} */,
  {32'hc0c486ba, 32'hbfbddb20} /* (21, 0, 14) {real, imag} */,
  {32'hc0cc025a, 32'hbf4bdb0a} /* (21, 0, 13) {real, imag} */,
  {32'h3c77c880, 32'hc1432352} /* (21, 0, 12) {real, imag} */,
  {32'hc0cff886, 32'hc187efcb} /* (21, 0, 11) {real, imag} */,
  {32'hc0ab3a82, 32'hc1062763} /* (21, 0, 10) {real, imag} */,
  {32'hbe9959d8, 32'hc0d9625b} /* (21, 0, 9) {real, imag} */,
  {32'hbe599b40, 32'hc11d53fb} /* (21, 0, 8) {real, imag} */,
  {32'hc12e8188, 32'hbfa12784} /* (21, 0, 7) {real, imag} */,
  {32'h3f85be44, 32'h41655fd7} /* (21, 0, 6) {real, imag} */,
  {32'h41811669, 32'h41a64745} /* (21, 0, 5) {real, imag} */,
  {32'h417725bb, 32'h40fdf330} /* (21, 0, 4) {real, imag} */,
  {32'h40d5cdbc, 32'h40b7fdfc} /* (21, 0, 3) {real, imag} */,
  {32'h414a9a80, 32'h415ee0d4} /* (21, 0, 2) {real, imag} */,
  {32'h41f22ace, 32'h411d23ee} /* (21, 0, 1) {real, imag} */,
  {32'h41838a36, 32'h411c4ca4} /* (21, 0, 0) {real, imag} */,
  {32'h40927f7b, 32'h3fb7458c} /* (20, 31, 31) {real, imag} */,
  {32'h41340956, 32'h40f9ab78} /* (20, 31, 30) {real, imag} */,
  {32'h410a3ee6, 32'h40e551f6} /* (20, 31, 29) {real, imag} */,
  {32'h4027451c, 32'hbfbe73ed} /* (20, 31, 28) {real, imag} */,
  {32'hbf7b9978, 32'h3f7a2252} /* (20, 31, 27) {real, imag} */,
  {32'hc0843346, 32'h3fc34b66} /* (20, 31, 26) {real, imag} */,
  {32'hc10ebee0, 32'hbf850bd0} /* (20, 31, 25) {real, imag} */,
  {32'hc01b27ba, 32'hbfa005d8} /* (20, 31, 24) {real, imag} */,
  {32'hbfe08cef, 32'hbe546400} /* (20, 31, 23) {real, imag} */,
  {32'hc0cac39c, 32'h3e083a00} /* (20, 31, 22) {real, imag} */,
  {32'h40a70144, 32'hc05f4c25} /* (20, 31, 21) {real, imag} */,
  {32'h414cbad5, 32'h400ca9c7} /* (20, 31, 20) {real, imag} */,
  {32'h40b5d20c, 32'h40d8f52d} /* (20, 31, 19) {real, imag} */,
  {32'h40e8c5de, 32'h40a156e6} /* (20, 31, 18) {real, imag} */,
  {32'h40c21526, 32'h3f4d2908} /* (20, 31, 17) {real, imag} */,
  {32'hc01c42b2, 32'h3eabd230} /* (20, 31, 16) {real, imag} */,
  {32'h3fb77579, 32'h408b5b29} /* (20, 31, 15) {real, imag} */,
  {32'h3bd88400, 32'hbf545254} /* (20, 31, 14) {real, imag} */,
  {32'h403da618, 32'hc0eda037} /* (20, 31, 13) {real, imag} */,
  {32'h40eba633, 32'hc0256502} /* (20, 31, 12) {real, imag} */,
  {32'h3ff14a9c, 32'h40338bba} /* (20, 31, 11) {real, imag} */,
  {32'h40d2f75d, 32'hbfbe7b00} /* (20, 31, 10) {real, imag} */,
  {32'hbf365db4, 32'hc0c68aa9} /* (20, 31, 9) {real, imag} */,
  {32'hc0f40855, 32'hc0fa0836} /* (20, 31, 8) {real, imag} */,
  {32'hc10afe98, 32'hc0540d06} /* (20, 31, 7) {real, imag} */,
  {32'hc105e55c, 32'hc01fd61c} /* (20, 31, 6) {real, imag} */,
  {32'h3fab213a, 32'h3f5cc390} /* (20, 31, 5) {real, imag} */,
  {32'h4185ec12, 32'h3efbd7b0} /* (20, 31, 4) {real, imag} */,
  {32'h4112a76c, 32'h4065d586} /* (20, 31, 3) {real, imag} */,
  {32'h403c3d4f, 32'h40028836} /* (20, 31, 2) {real, imag} */,
  {32'hc07b004b, 32'hc0dee045} /* (20, 31, 1) {real, imag} */,
  {32'hbf964223, 32'hc0ae111d} /* (20, 31, 0) {real, imag} */,
  {32'hc08ac7c5, 32'h3e360e46} /* (20, 30, 31) {real, imag} */,
  {32'h408713ba, 32'hc0835145} /* (20, 30, 30) {real, imag} */,
  {32'h3e59cd60, 32'hbfcc658c} /* (20, 30, 29) {real, imag} */,
  {32'h3f3500b3, 32'h3e48fe70} /* (20, 30, 28) {real, imag} */,
  {32'hbee0f4a8, 32'h3f187d5c} /* (20, 30, 27) {real, imag} */,
  {32'h41319411, 32'h3fdd6878} /* (20, 30, 26) {real, imag} */,
  {32'h413eb510, 32'h41096033} /* (20, 30, 25) {real, imag} */,
  {32'h416a6b9d, 32'h4085a184} /* (20, 30, 24) {real, imag} */,
  {32'h403717c8, 32'hc0add2fb} /* (20, 30, 23) {real, imag} */,
  {32'hc06f0114, 32'h4082d7c4} /* (20, 30, 22) {real, imag} */,
  {32'h40574885, 32'hbe88aca8} /* (20, 30, 21) {real, imag} */,
  {32'hbff65480, 32'h406e03dc} /* (20, 30, 20) {real, imag} */,
  {32'hc027bb5c, 32'h400a8c44} /* (20, 30, 19) {real, imag} */,
  {32'hbfcdb5af, 32'hc03b482d} /* (20, 30, 18) {real, imag} */,
  {32'hc09cdd4d, 32'hc0421a0d} /* (20, 30, 17) {real, imag} */,
  {32'hc0f28524, 32'hbf7235d0} /* (20, 30, 16) {real, imag} */,
  {32'h4040318c, 32'hbfe06ba4} /* (20, 30, 15) {real, imag} */,
  {32'hbf1cf88d, 32'h401395c0} /* (20, 30, 14) {real, imag} */,
  {32'hc04c88e4, 32'hc046b553} /* (20, 30, 13) {real, imag} */,
  {32'hbfac476d, 32'hc1843b3a} /* (20, 30, 12) {real, imag} */,
  {32'hc11d7d7b, 32'hc11b3de2} /* (20, 30, 11) {real, imag} */,
  {32'hbfce3dfc, 32'h40d7b43a} /* (20, 30, 10) {real, imag} */,
  {32'h3f7bac97, 32'h418ba996} /* (20, 30, 9) {real, imag} */,
  {32'hc1041e85, 32'h40a7c498} /* (20, 30, 8) {real, imag} */,
  {32'hc123c697, 32'hbf929f9c} /* (20, 30, 7) {real, imag} */,
  {32'hc0e3cf74, 32'hc0ddbb43} /* (20, 30, 6) {real, imag} */,
  {32'h404bfe89, 32'hc07b5072} /* (20, 30, 5) {real, imag} */,
  {32'hc008471f, 32'h3fea4562} /* (20, 30, 4) {real, imag} */,
  {32'hc0e47922, 32'hc020f024} /* (20, 30, 3) {real, imag} */,
  {32'hbd5db940, 32'hc0f68e96} /* (20, 30, 2) {real, imag} */,
  {32'h40b3f7ad, 32'hc0a8ad60} /* (20, 30, 1) {real, imag} */,
  {32'hc045cbcc, 32'h40257501} /* (20, 30, 0) {real, imag} */,
  {32'hc0353afb, 32'h3f0b43a5} /* (20, 29, 31) {real, imag} */,
  {32'h401d4230, 32'hc0168f76} /* (20, 29, 30) {real, imag} */,
  {32'h410c2a3c, 32'h3f818802} /* (20, 29, 29) {real, imag} */,
  {32'h4042799c, 32'h4090a6d5} /* (20, 29, 28) {real, imag} */,
  {32'h402d9d6e, 32'h40a014f6} /* (20, 29, 27) {real, imag} */,
  {32'h4045b393, 32'hc05c8966} /* (20, 29, 26) {real, imag} */,
  {32'hbf5284e0, 32'hbff0a340} /* (20, 29, 25) {real, imag} */,
  {32'hbf99e3e6, 32'hc02f8710} /* (20, 29, 24) {real, imag} */,
  {32'hbf12ec7d, 32'h3e710300} /* (20, 29, 23) {real, imag} */,
  {32'hc0944c00, 32'hbfed2c8a} /* (20, 29, 22) {real, imag} */,
  {32'hc040040f, 32'hc07faef8} /* (20, 29, 21) {real, imag} */,
  {32'hbfaa52b4, 32'hc15bc926} /* (20, 29, 20) {real, imag} */,
  {32'h404453d8, 32'hc130638a} /* (20, 29, 19) {real, imag} */,
  {32'h4102422c, 32'hc10db2e0} /* (20, 29, 18) {real, imag} */,
  {32'h40cca746, 32'hc0c35aea} /* (20, 29, 17) {real, imag} */,
  {32'h4007d55a, 32'hbf4a8760} /* (20, 29, 16) {real, imag} */,
  {32'h3ecd0020, 32'h3f0e0c9c} /* (20, 29, 15) {real, imag} */,
  {32'hc136cf14, 32'h40f046d2} /* (20, 29, 14) {real, imag} */,
  {32'hc10e5810, 32'h40ad9f6a} /* (20, 29, 13) {real, imag} */,
  {32'h40b3dbfd, 32'h40ff8f1c} /* (20, 29, 12) {real, imag} */,
  {32'h40356287, 32'h41102772} /* (20, 29, 11) {real, imag} */,
  {32'hbfef1a64, 32'h40cfdbcc} /* (20, 29, 10) {real, imag} */,
  {32'h3f2fcca2, 32'hc0c24bd4} /* (20, 29, 9) {real, imag} */,
  {32'h401647c8, 32'hc09aa186} /* (20, 29, 8) {real, imag} */,
  {32'h3f9d1c80, 32'hc0100ab6} /* (20, 29, 7) {real, imag} */,
  {32'h4090c779, 32'h3fbfe3ec} /* (20, 29, 6) {real, imag} */,
  {32'h401a278a, 32'h4109e036} /* (20, 29, 5) {real, imag} */,
  {32'h4046920a, 32'h40c9ea0b} /* (20, 29, 4) {real, imag} */,
  {32'h40c74af5, 32'h40582dbe} /* (20, 29, 3) {real, imag} */,
  {32'h3fc4d182, 32'hc07a4882} /* (20, 29, 2) {real, imag} */,
  {32'h3f93d1e4, 32'h408ce25e} /* (20, 29, 1) {real, imag} */,
  {32'h409c3bd2, 32'h3f280700} /* (20, 29, 0) {real, imag} */,
  {32'hbf4d75ba, 32'h3f9a7535} /* (20, 28, 31) {real, imag} */,
  {32'hc095d472, 32'h408675a2} /* (20, 28, 30) {real, imag} */,
  {32'h40a4d98a, 32'h40933f2f} /* (20, 28, 29) {real, imag} */,
  {32'h40fe85aa, 32'h412dfc52} /* (20, 28, 28) {real, imag} */,
  {32'h3f46d2b0, 32'h410de0b6} /* (20, 28, 27) {real, imag} */,
  {32'h4078e0e2, 32'h3f0ad014} /* (20, 28, 26) {real, imag} */,
  {32'h40884873, 32'hc097cf0f} /* (20, 28, 25) {real, imag} */,
  {32'hbfd5b34c, 32'hc0d473a1} /* (20, 28, 24) {real, imag} */,
  {32'hc0d424c6, 32'hc055d258} /* (20, 28, 23) {real, imag} */,
  {32'hc132fd9c, 32'h406d9e95} /* (20, 28, 22) {real, imag} */,
  {32'hc12d5ac4, 32'h40e3050d} /* (20, 28, 21) {real, imag} */,
  {32'hbfcda4ac, 32'hbd530180} /* (20, 28, 20) {real, imag} */,
  {32'hc0ce3859, 32'h406b00d2} /* (20, 28, 19) {real, imag} */,
  {32'hbf91d650, 32'h40ddebc0} /* (20, 28, 18) {real, imag} */,
  {32'h3d4b4980, 32'hbf9dfc08} /* (20, 28, 17) {real, imag} */,
  {32'hc08d88d5, 32'h3fb133fc} /* (20, 28, 16) {real, imag} */,
  {32'hc09ab018, 32'h4097a70b} /* (20, 28, 15) {real, imag} */,
  {32'hc0b64255, 32'hbf585248} /* (20, 28, 14) {real, imag} */,
  {32'hc02be6ef, 32'hc0c1d1ff} /* (20, 28, 13) {real, imag} */,
  {32'h40a00e4e, 32'hc07ddbb6} /* (20, 28, 12) {real, imag} */,
  {32'h4140f4e2, 32'hc00d0720} /* (20, 28, 11) {real, imag} */,
  {32'hc00c1875, 32'h3d9b62f0} /* (20, 28, 10) {real, imag} */,
  {32'hc0a6d77a, 32'h3f6f25bd} /* (20, 28, 9) {real, imag} */,
  {32'hc1043186, 32'hbed93bf8} /* (20, 28, 8) {real, imag} */,
  {32'hc118ac2f, 32'h40ad4ce0} /* (20, 28, 7) {real, imag} */,
  {32'hc093e484, 32'h3f9d6c76} /* (20, 28, 6) {real, imag} */,
  {32'hc0587568, 32'h400591d2} /* (20, 28, 5) {real, imag} */,
  {32'h3feaca17, 32'h40aad78c} /* (20, 28, 4) {real, imag} */,
  {32'hbf8eeb52, 32'hc026f99b} /* (20, 28, 3) {real, imag} */,
  {32'hc0b36a2e, 32'h3eae2988} /* (20, 28, 2) {real, imag} */,
  {32'hc02f7de1, 32'hc0c10199} /* (20, 28, 1) {real, imag} */,
  {32'h3ff244e8, 32'hc069add6} /* (20, 28, 0) {real, imag} */,
  {32'hbf848c01, 32'hbff8444a} /* (20, 27, 31) {real, imag} */,
  {32'h3fb078b4, 32'hc07833f3} /* (20, 27, 30) {real, imag} */,
  {32'hc06a7ba7, 32'hbce30b00} /* (20, 27, 29) {real, imag} */,
  {32'hc0718c37, 32'h41051cba} /* (20, 27, 28) {real, imag} */,
  {32'h400e5ea5, 32'h410da7af} /* (20, 27, 27) {real, imag} */,
  {32'h40501231, 32'h3fc24cec} /* (20, 27, 26) {real, imag} */,
  {32'hc10cfbce, 32'hc0c871a2} /* (20, 27, 25) {real, imag} */,
  {32'hbec37546, 32'hbfa16f64} /* (20, 27, 24) {real, imag} */,
  {32'h4149ebbd, 32'h40177f3f} /* (20, 27, 23) {real, imag} */,
  {32'h3f2c715e, 32'hc0c395ae} /* (20, 27, 22) {real, imag} */,
  {32'hc12a1d75, 32'hc0ba60e2} /* (20, 27, 21) {real, imag} */,
  {32'hbfb64a08, 32'hbfa3bc3c} /* (20, 27, 20) {real, imag} */,
  {32'h3fb4feba, 32'hc0cc1a48} /* (20, 27, 19) {real, imag} */,
  {32'h3fefb4a6, 32'h410f032c} /* (20, 27, 18) {real, imag} */,
  {32'hbf3dfe14, 32'h4139d50c} /* (20, 27, 17) {real, imag} */,
  {32'hc057cd20, 32'h3ea18840} /* (20, 27, 16) {real, imag} */,
  {32'hc10a5e28, 32'hc094326c} /* (20, 27, 15) {real, imag} */,
  {32'hc11950d8, 32'hc08de13e} /* (20, 27, 14) {real, imag} */,
  {32'hc08d6d52, 32'h3e13cabe} /* (20, 27, 13) {real, imag} */,
  {32'hc0d63767, 32'hc09ae66b} /* (20, 27, 12) {real, imag} */,
  {32'hc05e439c, 32'hc10d25ca} /* (20, 27, 11) {real, imag} */,
  {32'h3e430ed0, 32'hc15465d8} /* (20, 27, 10) {real, imag} */,
  {32'h400f1a28, 32'hc0efdd88} /* (20, 27, 9) {real, imag} */,
  {32'h3fb07b98, 32'hbf8e42e8} /* (20, 27, 8) {real, imag} */,
  {32'h40282010, 32'h40c76f14} /* (20, 27, 7) {real, imag} */,
  {32'hc0234632, 32'h407d79b4} /* (20, 27, 6) {real, imag} */,
  {32'h3f7d71d4, 32'h416666c0} /* (20, 27, 5) {real, imag} */,
  {32'h40d64450, 32'h40d1d160} /* (20, 27, 4) {real, imag} */,
  {32'h41071c96, 32'h41045811} /* (20, 27, 3) {real, imag} */,
  {32'h409c36e6, 32'h4183bd65} /* (20, 27, 2) {real, imag} */,
  {32'hbf4316f3, 32'h404feb88} /* (20, 27, 1) {real, imag} */,
  {32'hc01db97a, 32'h3da90f40} /* (20, 27, 0) {real, imag} */,
  {32'h3fbcdef6, 32'h3f70ce86} /* (20, 26, 31) {real, imag} */,
  {32'h4002ad94, 32'hbf06af08} /* (20, 26, 30) {real, imag} */,
  {32'h3f0f0f49, 32'hc0258ae6} /* (20, 26, 29) {real, imag} */,
  {32'hc02600c4, 32'hbf308238} /* (20, 26, 28) {real, imag} */,
  {32'h3ddc47f0, 32'h40b6fb68} /* (20, 26, 27) {real, imag} */,
  {32'hbfefe1e2, 32'h3f40ffee} /* (20, 26, 26) {real, imag} */,
  {32'hbf95c5e2, 32'hc091b656} /* (20, 26, 25) {real, imag} */,
  {32'hc0e3f0f0, 32'hc03a8217} /* (20, 26, 24) {real, imag} */,
  {32'hc0569e36, 32'hc0a059d5} /* (20, 26, 23) {real, imag} */,
  {32'h3f8fb32a, 32'hc0a9d54a} /* (20, 26, 22) {real, imag} */,
  {32'hc018c12e, 32'h3f4ce0fc} /* (20, 26, 21) {real, imag} */,
  {32'hbe34d668, 32'hbfca007e} /* (20, 26, 20) {real, imag} */,
  {32'hbff51176, 32'hc053dd5f} /* (20, 26, 19) {real, imag} */,
  {32'hbdeb7370, 32'hc1487bd0} /* (20, 26, 18) {real, imag} */,
  {32'hbf4ee500, 32'hc154df6a} /* (20, 26, 17) {real, imag} */,
  {32'h40c6fa9a, 32'hc001a23e} /* (20, 26, 16) {real, imag} */,
  {32'h40ec52b6, 32'hbed48cb0} /* (20, 26, 15) {real, imag} */,
  {32'hc02781db, 32'hc0ce5c22} /* (20, 26, 14) {real, imag} */,
  {32'hc0a17ca8, 32'hc0c05598} /* (20, 26, 13) {real, imag} */,
  {32'hc09b0f52, 32'hc0699be8} /* (20, 26, 12) {real, imag} */,
  {32'h3f7a4b0b, 32'hbefea588} /* (20, 26, 11) {real, imag} */,
  {32'h40121734, 32'h3ffbe91e} /* (20, 26, 10) {real, imag} */,
  {32'hc0b0b98d, 32'h3fcfc400} /* (20, 26, 9) {real, imag} */,
  {32'hc1115ce5, 32'h40c94733} /* (20, 26, 8) {real, imag} */,
  {32'hbf3e3750, 32'h410897bd} /* (20, 26, 7) {real, imag} */,
  {32'hbe11edb4, 32'h40ffc716} /* (20, 26, 6) {real, imag} */,
  {32'hbfeb4a90, 32'hbecf5444} /* (20, 26, 5) {real, imag} */,
  {32'h3f318f32, 32'hc04fef10} /* (20, 26, 4) {real, imag} */,
  {32'h3d44e840, 32'hc062d935} /* (20, 26, 3) {real, imag} */,
  {32'hc0413ba0, 32'hbfa2c8d1} /* (20, 26, 2) {real, imag} */,
  {32'hc08e77f4, 32'h40314047} /* (20, 26, 1) {real, imag} */,
  {32'hbfe0edff, 32'h3ec7f58c} /* (20, 26, 0) {real, imag} */,
  {32'hbfa26ad6, 32'hbfc41f34} /* (20, 25, 31) {real, imag} */,
  {32'hbdae1400, 32'h3eb033d0} /* (20, 25, 30) {real, imag} */,
  {32'h3f87dfaf, 32'hbf927818} /* (20, 25, 29) {real, imag} */,
  {32'h3fd324c3, 32'hc0b3f141} /* (20, 25, 28) {real, imag} */,
  {32'hbf7283e8, 32'hbf2f6960} /* (20, 25, 27) {real, imag} */,
  {32'h4091481e, 32'hbf629e40} /* (20, 25, 26) {real, imag} */,
  {32'h412f18c8, 32'hc0bbe836} /* (20, 25, 25) {real, imag} */,
  {32'h408b0e6c, 32'hc0334a25} /* (20, 25, 24) {real, imag} */,
  {32'hc07479fe, 32'h40ef5bfe} /* (20, 25, 23) {real, imag} */,
  {32'hbe021460, 32'h40d87e62} /* (20, 25, 22) {real, imag} */,
  {32'h40529666, 32'h3ea639a0} /* (20, 25, 21) {real, imag} */,
  {32'h3fd5f970, 32'h4047dfaa} /* (20, 25, 20) {real, imag} */,
  {32'h3fc266b0, 32'h4047612d} /* (20, 25, 19) {real, imag} */,
  {32'hbe9bd958, 32'h4103b19f} /* (20, 25, 18) {real, imag} */,
  {32'hbfd4d99a, 32'hc019a4ae} /* (20, 25, 17) {real, imag} */,
  {32'hc01aefec, 32'hbe1c23f0} /* (20, 25, 16) {real, imag} */,
  {32'hbfcbbcd4, 32'h40ce25f3} /* (20, 25, 15) {real, imag} */,
  {32'h403f244c, 32'h3fcf0a3a} /* (20, 25, 14) {real, imag} */,
  {32'h4084ad0e, 32'hbf419081} /* (20, 25, 13) {real, imag} */,
  {32'h403258b1, 32'h4049919d} /* (20, 25, 12) {real, imag} */,
  {32'h3f800eb2, 32'h40bb0080} /* (20, 25, 11) {real, imag} */,
  {32'h4064275b, 32'h4118dd3c} /* (20, 25, 10) {real, imag} */,
  {32'h406462b8, 32'h40eb9677} /* (20, 25, 9) {real, imag} */,
  {32'h411c2dd6, 32'h40e08b10} /* (20, 25, 8) {real, imag} */,
  {32'hbf4ded1b, 32'h4084547f} /* (20, 25, 7) {real, imag} */,
  {32'hc087a42a, 32'h3e438520} /* (20, 25, 6) {real, imag} */,
  {32'hc0ce2c48, 32'hbed9c552} /* (20, 25, 5) {real, imag} */,
  {32'hc0a3ba26, 32'h40d68cef} /* (20, 25, 4) {real, imag} */,
  {32'hbe9210d0, 32'h3f0c28f4} /* (20, 25, 3) {real, imag} */,
  {32'h406c9a77, 32'h402e94ba} /* (20, 25, 2) {real, imag} */,
  {32'h3fdb6b03, 32'h3f398e32} /* (20, 25, 1) {real, imag} */,
  {32'h3f33ab66, 32'h3fdc1ae4} /* (20, 25, 0) {real, imag} */,
  {32'h3fca20c2, 32'h40a8ec91} /* (20, 24, 31) {real, imag} */,
  {32'hbed01e12, 32'h4105c3a2} /* (20, 24, 30) {real, imag} */,
  {32'hc04af867, 32'h4119a730} /* (20, 24, 29) {real, imag} */,
  {32'hc09ae6e3, 32'h3f8d8506} /* (20, 24, 28) {real, imag} */,
  {32'h3f34f928, 32'hbec3c50b} /* (20, 24, 27) {real, imag} */,
  {32'hc00a52fb, 32'h4006d4ad} /* (20, 24, 26) {real, imag} */,
  {32'hc079be90, 32'hbf8c35e6} /* (20, 24, 25) {real, imag} */,
  {32'hbf6c3d50, 32'hc06fd0aa} /* (20, 24, 24) {real, imag} */,
  {32'h3fb464cf, 32'hc070ed6e} /* (20, 24, 23) {real, imag} */,
  {32'h3fb85ce8, 32'hc01ee279} /* (20, 24, 22) {real, imag} */,
  {32'hc01d0612, 32'hc0967452} /* (20, 24, 21) {real, imag} */,
  {32'hc0994ff8, 32'hc0a277cd} /* (20, 24, 20) {real, imag} */,
  {32'hbfd25452, 32'h4008f918} /* (20, 24, 19) {real, imag} */,
  {32'h405345a4, 32'h408ad3e4} /* (20, 24, 18) {real, imag} */,
  {32'h409674a4, 32'h4075d19c} /* (20, 24, 17) {real, imag} */,
  {32'h402a4b72, 32'h4049c3ef} /* (20, 24, 16) {real, imag} */,
  {32'h3f8e3be0, 32'h40980a98} /* (20, 24, 15) {real, imag} */,
  {32'hbf8f7a75, 32'h404cda79} /* (20, 24, 14) {real, imag} */,
  {32'hbf0925f0, 32'h3f991103} /* (20, 24, 13) {real, imag} */,
  {32'hbead5720, 32'h3e88d76c} /* (20, 24, 12) {real, imag} */,
  {32'h404464ff, 32'hbe5ef64c} /* (20, 24, 11) {real, imag} */,
  {32'h400991ed, 32'h3f893ec0} /* (20, 24, 10) {real, imag} */,
  {32'h409f0df7, 32'hbe0fd020} /* (20, 24, 9) {real, imag} */,
  {32'h406de8ee, 32'hc001afec} /* (20, 24, 8) {real, imag} */,
  {32'hc0513366, 32'hbfb66106} /* (20, 24, 7) {real, imag} */,
  {32'hbf8b26bf, 32'hc085f52c} /* (20, 24, 6) {real, imag} */,
  {32'h40007f96, 32'hbf94ee28} /* (20, 24, 5) {real, imag} */,
  {32'hbf54a7fa, 32'hc089cef4} /* (20, 24, 4) {real, imag} */,
  {32'hc02fa78f, 32'hc033af98} /* (20, 24, 3) {real, imag} */,
  {32'h3fc3aade, 32'hc08725c8} /* (20, 24, 2) {real, imag} */,
  {32'h409d9d7f, 32'hc08b292e} /* (20, 24, 1) {real, imag} */,
  {32'h40863e94, 32'hc043d78e} /* (20, 24, 0) {real, imag} */,
  {32'hc06962a9, 32'hbefb6d60} /* (20, 23, 31) {real, imag} */,
  {32'hc0f88169, 32'hbebae168} /* (20, 23, 30) {real, imag} */,
  {32'hc10246c6, 32'hc0795230} /* (20, 23, 29) {real, imag} */,
  {32'hc1023800, 32'hbf192392} /* (20, 23, 28) {real, imag} */,
  {32'hbfdf98d2, 32'hbea5db44} /* (20, 23, 27) {real, imag} */,
  {32'h3f7634f0, 32'h3ea48944} /* (20, 23, 26) {real, imag} */,
  {32'hbf0fedba, 32'h4035ad4d} /* (20, 23, 25) {real, imag} */,
  {32'hc047014b, 32'h408259c4} /* (20, 23, 24) {real, imag} */,
  {32'h3e1d6800, 32'h40057bc1} /* (20, 23, 23) {real, imag} */,
  {32'h4054c2dc, 32'h3d93ae60} /* (20, 23, 22) {real, imag} */,
  {32'h4053f31b, 32'h3e8e5ada} /* (20, 23, 21) {real, imag} */,
  {32'h409e5b70, 32'h3f312bd8} /* (20, 23, 20) {real, imag} */,
  {32'h3fcfe880, 32'h3edcee30} /* (20, 23, 19) {real, imag} */,
  {32'hbe7bfcf0, 32'hbf1db374} /* (20, 23, 18) {real, imag} */,
  {32'h3fc02022, 32'hbf404308} /* (20, 23, 17) {real, imag} */,
  {32'h401b8268, 32'hc07feba8} /* (20, 23, 16) {real, imag} */,
  {32'h403d8929, 32'hc094b7b1} /* (20, 23, 15) {real, imag} */,
  {32'h4030d0fe, 32'hbf452c74} /* (20, 23, 14) {real, imag} */,
  {32'h407d986d, 32'h409666cf} /* (20, 23, 13) {real, imag} */,
  {32'h40ce3294, 32'h3e233b48} /* (20, 23, 12) {real, imag} */,
  {32'h3e8d76d8, 32'h408d125a} /* (20, 23, 11) {real, imag} */,
  {32'hc09dc945, 32'h40ec0dbc} /* (20, 23, 10) {real, imag} */,
  {32'hbf7d4268, 32'h4046fe2c} /* (20, 23, 9) {real, imag} */,
  {32'h4017eabe, 32'h3f7d382a} /* (20, 23, 8) {real, imag} */,
  {32'hbea8bfe0, 32'hc012ee15} /* (20, 23, 7) {real, imag} */,
  {32'h402a12ca, 32'h4006c61c} /* (20, 23, 6) {real, imag} */,
  {32'h408cfc55, 32'h40e1257e} /* (20, 23, 5) {real, imag} */,
  {32'h3ffb0b4f, 32'h407d0b3e} /* (20, 23, 4) {real, imag} */,
  {32'hbefcc9a0, 32'h3ffc1656} /* (20, 23, 3) {real, imag} */,
  {32'h40bb0483, 32'hbf65d1b6} /* (20, 23, 2) {real, imag} */,
  {32'h3f274854, 32'h3fa8d85e} /* (20, 23, 1) {real, imag} */,
  {32'hc0996324, 32'hbf1bb53a} /* (20, 23, 0) {real, imag} */,
  {32'hc05dc376, 32'hbf24ba0a} /* (20, 22, 31) {real, imag} */,
  {32'hbf8a94c0, 32'hbd1e2bd0} /* (20, 22, 30) {real, imag} */,
  {32'hbe8c973a, 32'h4038a630} /* (20, 22, 29) {real, imag} */,
  {32'hbfbc96a7, 32'h401c7c84} /* (20, 22, 28) {real, imag} */,
  {32'hc022c970, 32'h401d6eee} /* (20, 22, 27) {real, imag} */,
  {32'hc0354f62, 32'hc07da799} /* (20, 22, 26) {real, imag} */,
  {32'hbf60b05a, 32'h3f37a19c} /* (20, 22, 25) {real, imag} */,
  {32'hbf83e9a6, 32'h3fd89872} /* (20, 22, 24) {real, imag} */,
  {32'h3fc1675b, 32'h40cc6666} /* (20, 22, 23) {real, imag} */,
  {32'hc091be62, 32'h408ba102} /* (20, 22, 22) {real, imag} */,
  {32'hc05e7d54, 32'hbeed3bfc} /* (20, 22, 21) {real, imag} */,
  {32'hc01484b0, 32'hbff6ba21} /* (20, 22, 20) {real, imag} */,
  {32'h3e039be0, 32'hc0c09b83} /* (20, 22, 19) {real, imag} */,
  {32'h40086bd0, 32'hc03d580a} /* (20, 22, 18) {real, imag} */,
  {32'h400d3eb4, 32'hc0710e98} /* (20, 22, 17) {real, imag} */,
  {32'h4022f3b1, 32'h3f2eac33} /* (20, 22, 16) {real, imag} */,
  {32'h40a16420, 32'h3faa2fb0} /* (20, 22, 15) {real, imag} */,
  {32'h403d4f8c, 32'hbe9f0e70} /* (20, 22, 14) {real, imag} */,
  {32'h401fe4fd, 32'hbfbc45c0} /* (20, 22, 13) {real, imag} */,
  {32'hbfacd0b2, 32'hbe085da0} /* (20, 22, 12) {real, imag} */,
  {32'hc07cdcc2, 32'h402ca47d} /* (20, 22, 11) {real, imag} */,
  {32'hbe819e54, 32'h3f51ee78} /* (20, 22, 10) {real, imag} */,
  {32'h40347171, 32'h3fd6afa0} /* (20, 22, 9) {real, imag} */,
  {32'h40602af4, 32'h3f7f5734} /* (20, 22, 8) {real, imag} */,
  {32'h4038eea8, 32'hbfdf7d69} /* (20, 22, 7) {real, imag} */,
  {32'hbedc3796, 32'hbfde3f9e} /* (20, 22, 6) {real, imag} */,
  {32'hc040ac2e, 32'hc025d32f} /* (20, 22, 5) {real, imag} */,
  {32'hc0043578, 32'h405d5ba0} /* (20, 22, 4) {real, imag} */,
  {32'h3fb36f2d, 32'h3d8a3600} /* (20, 22, 3) {real, imag} */,
  {32'h4065a9cc, 32'hbf82b2d0} /* (20, 22, 2) {real, imag} */,
  {32'hc048649e, 32'h404188e9} /* (20, 22, 1) {real, imag} */,
  {32'hc09e30fa, 32'h3fbd0a9d} /* (20, 22, 0) {real, imag} */,
  {32'h4007f9f4, 32'h3f59e38d} /* (20, 21, 31) {real, imag} */,
  {32'h3f1c68da, 32'h4097f131} /* (20, 21, 30) {real, imag} */,
  {32'h3f59a2dc, 32'h40a63ece} /* (20, 21, 29) {real, imag} */,
  {32'h400403eb, 32'h40d2ac35} /* (20, 21, 28) {real, imag} */,
  {32'h3fefb024, 32'h4081c487} /* (20, 21, 27) {real, imag} */,
  {32'hbfd01952, 32'hbf61bbc3} /* (20, 21, 26) {real, imag} */,
  {32'hbfb39ab9, 32'hc02de27f} /* (20, 21, 25) {real, imag} */,
  {32'h3e270e94, 32'h405942ec} /* (20, 21, 24) {real, imag} */,
  {32'h3e5febd0, 32'h408dd92e} /* (20, 21, 23) {real, imag} */,
  {32'hbf96c83f, 32'hc058a625} /* (20, 21, 22) {real, imag} */,
  {32'h3df34af0, 32'hc01efe66} /* (20, 21, 21) {real, imag} */,
  {32'h402489dd, 32'h3c610c00} /* (20, 21, 20) {real, imag} */,
  {32'h3fac8b90, 32'hc02705d4} /* (20, 21, 19) {real, imag} */,
  {32'h3f24458c, 32'hc089ac9e} /* (20, 21, 18) {real, imag} */,
  {32'hc00d13ed, 32'h3f95c150} /* (20, 21, 17) {real, imag} */,
  {32'hc04dbac8, 32'h3feb8b1d} /* (20, 21, 16) {real, imag} */,
  {32'hc09f6bfc, 32'h3f8940a4} /* (20, 21, 15) {real, imag} */,
  {32'h3f206d76, 32'h3ec86fdc} /* (20, 21, 14) {real, imag} */,
  {32'h3f98fb65, 32'h3fdbcd2e} /* (20, 21, 13) {real, imag} */,
  {32'hbf1b0b4e, 32'h3f01cf24} /* (20, 21, 12) {real, imag} */,
  {32'h407fe7dc, 32'h40576a84} /* (20, 21, 11) {real, imag} */,
  {32'h3eb22198, 32'h4051be76} /* (20, 21, 10) {real, imag} */,
  {32'h3ecdd518, 32'h3f9df813} /* (20, 21, 9) {real, imag} */,
  {32'h40137b0c, 32'hbf485142} /* (20, 21, 8) {real, imag} */,
  {32'hbfb2d4d8, 32'h404859bb} /* (20, 21, 7) {real, imag} */,
  {32'hc0700b97, 32'h408cb2c6} /* (20, 21, 6) {real, imag} */,
  {32'hc0a99564, 32'hbf4db454} /* (20, 21, 5) {real, imag} */,
  {32'hc03519dd, 32'hbff6fb0e} /* (20, 21, 4) {real, imag} */,
  {32'h3feee4d4, 32'hbf54bea0} /* (20, 21, 3) {real, imag} */,
  {32'hc02cf0aa, 32'h3fc2afbe} /* (20, 21, 2) {real, imag} */,
  {32'hc024d10b, 32'h40492eb6} /* (20, 21, 1) {real, imag} */,
  {32'h406a63a6, 32'hbecef514} /* (20, 21, 0) {real, imag} */,
  {32'h3fe2a290, 32'hbf8c8c0d} /* (20, 20, 31) {real, imag} */,
  {32'hbf325e7c, 32'hc01e609c} /* (20, 20, 30) {real, imag} */,
  {32'hbff9b1b2, 32'hc023404c} /* (20, 20, 29) {real, imag} */,
  {32'h3f61411e, 32'hbeced98c} /* (20, 20, 28) {real, imag} */,
  {32'hbff9be42, 32'h3f758df6} /* (20, 20, 27) {real, imag} */,
  {32'hbf826c30, 32'hc02c3fea} /* (20, 20, 26) {real, imag} */,
  {32'hbfcdf028, 32'hbf8d6d06} /* (20, 20, 25) {real, imag} */,
  {32'hbf7a1a11, 32'hc010ff0a} /* (20, 20, 24) {real, imag} */,
  {32'hbfd187b6, 32'hc0658f61} /* (20, 20, 23) {real, imag} */,
  {32'h40597f4d, 32'hc074ebb7} /* (20, 20, 22) {real, imag} */,
  {32'h404f6f79, 32'hbf1f4212} /* (20, 20, 21) {real, imag} */,
  {32'h3f8213dd, 32'hbf586c94} /* (20, 20, 20) {real, imag} */,
  {32'h402cc7a1, 32'hc03f70b6} /* (20, 20, 19) {real, imag} */,
  {32'h402320b5, 32'hbdfc7fc0} /* (20, 20, 18) {real, imag} */,
  {32'hbe61590c, 32'h4091cf50} /* (20, 20, 17) {real, imag} */,
  {32'hc0050fa4, 32'h3e74ae90} /* (20, 20, 16) {real, imag} */,
  {32'hbf09e54e, 32'hbfabdd6c} /* (20, 20, 15) {real, imag} */,
  {32'h3f18875a, 32'h3edec85c} /* (20, 20, 14) {real, imag} */,
  {32'h3fa3642a, 32'hbfad9c26} /* (20, 20, 13) {real, imag} */,
  {32'h40cd1a03, 32'hc03ff9f6} /* (20, 20, 12) {real, imag} */,
  {32'h4093f55e, 32'hbfc64a17} /* (20, 20, 11) {real, imag} */,
  {32'h3fee8dc5, 32'hc01f2bec} /* (20, 20, 10) {real, imag} */,
  {32'h3fe95962, 32'hc0a839fc} /* (20, 20, 9) {real, imag} */,
  {32'h3fe690e2, 32'hc0a41432} /* (20, 20, 8) {real, imag} */,
  {32'h3f9796dd, 32'hbf900301} /* (20, 20, 7) {real, imag} */,
  {32'h3fb86cc6, 32'h4006e509} /* (20, 20, 6) {real, imag} */,
  {32'hbfd19c73, 32'h3f5bf9ae} /* (20, 20, 5) {real, imag} */,
  {32'h3f842a89, 32'hbe667cd2} /* (20, 20, 4) {real, imag} */,
  {32'h400d82b2, 32'hc03ac074} /* (20, 20, 3) {real, imag} */,
  {32'h3f9332ca, 32'hc0b0b0ea} /* (20, 20, 2) {real, imag} */,
  {32'h3ff77d34, 32'hc0299707} /* (20, 20, 1) {real, imag} */,
  {32'h3f331f19, 32'h3f9f0b45} /* (20, 20, 0) {real, imag} */,
  {32'hc076af4f, 32'h400b361a} /* (20, 19, 31) {real, imag} */,
  {32'hc0bb396e, 32'h3ff0c821} /* (20, 19, 30) {real, imag} */,
  {32'hbf34f89c, 32'h3f090f83} /* (20, 19, 29) {real, imag} */,
  {32'h3ff35ea9, 32'hbfd4b4f4} /* (20, 19, 28) {real, imag} */,
  {32'h4011668c, 32'hc03fd5cc} /* (20, 19, 27) {real, imag} */,
  {32'h3ffc1c36, 32'hbfdc75af} /* (20, 19, 26) {real, imag} */,
  {32'h400d0536, 32'h3fa2e14f} /* (20, 19, 25) {real, imag} */,
  {32'h40015380, 32'h403c5f14} /* (20, 19, 24) {real, imag} */,
  {32'h3ff395fa, 32'h3fbc4767} /* (20, 19, 23) {real, imag} */,
  {32'hbe799e58, 32'hbd9e1f80} /* (20, 19, 22) {real, imag} */,
  {32'h3fb943e0, 32'hbfe9d1a2} /* (20, 19, 21) {real, imag} */,
  {32'h402ea799, 32'hbf798718} /* (20, 19, 20) {real, imag} */,
  {32'h401fbb1c, 32'h401753fa} /* (20, 19, 19) {real, imag} */,
  {32'h3fc125c8, 32'h40763d67} /* (20, 19, 18) {real, imag} */,
  {32'h405347cf, 32'h405fd123} /* (20, 19, 17) {real, imag} */,
  {32'h3f260f4c, 32'h3fa768a5} /* (20, 19, 16) {real, imag} */,
  {32'h3ffbc6d7, 32'hbf85b767} /* (20, 19, 15) {real, imag} */,
  {32'h408b8eac, 32'hc0221685} /* (20, 19, 14) {real, imag} */,
  {32'h400366be, 32'hbfed97ae} /* (20, 19, 13) {real, imag} */,
  {32'h3fedf57c, 32'hc00667f8} /* (20, 19, 12) {real, imag} */,
  {32'h3eb22150, 32'hbf90c394} /* (20, 19, 11) {real, imag} */,
  {32'hc02eaf02, 32'h3f17a964} /* (20, 19, 10) {real, imag} */,
  {32'hc015322c, 32'h3f6fd014} /* (20, 19, 9) {real, imag} */,
  {32'hbf7f18e0, 32'hbc2bb900} /* (20, 19, 8) {real, imag} */,
  {32'hbfb7c818, 32'h3e4c85a0} /* (20, 19, 7) {real, imag} */,
  {32'hbe6094b8, 32'hbe8625e8} /* (20, 19, 6) {real, imag} */,
  {32'hbfa3ba96, 32'hbf07379a} /* (20, 19, 5) {real, imag} */,
  {32'h3ee71210, 32'h3faa3b68} /* (20, 19, 4) {real, imag} */,
  {32'h404eb4e2, 32'hbecd80a8} /* (20, 19, 3) {real, imag} */,
  {32'hbd91a320, 32'hc0236fce} /* (20, 19, 2) {real, imag} */,
  {32'h402876ea, 32'hc041c33f} /* (20, 19, 1) {real, imag} */,
  {32'h3ee383b4, 32'hbfd71353} /* (20, 19, 0) {real, imag} */,
  {32'hc0290316, 32'hbf73b138} /* (20, 18, 31) {real, imag} */,
  {32'h3f183f63, 32'hbf851ad7} /* (20, 18, 30) {real, imag} */,
  {32'h3f35f6a0, 32'hc01aff7f} /* (20, 18, 29) {real, imag} */,
  {32'hbf2a5e6a, 32'h3d723780} /* (20, 18, 28) {real, imag} */,
  {32'hbf9b1810, 32'h406c552c} /* (20, 18, 27) {real, imag} */,
  {32'hbf55d91a, 32'h405f8c44} /* (20, 18, 26) {real, imag} */,
  {32'hbfc60a87, 32'h4069e91b} /* (20, 18, 25) {real, imag} */,
  {32'h3ff098da, 32'h3e2695e8} /* (20, 18, 24) {real, imag} */,
  {32'h3f96c77b, 32'hc01b2742} /* (20, 18, 23) {real, imag} */,
  {32'hbe468ce8, 32'hc06da567} /* (20, 18, 22) {real, imag} */,
  {32'h3fc14828, 32'hbfbad7b1} /* (20, 18, 21) {real, imag} */,
  {32'h3fbd9c0a, 32'h3f41a7cc} /* (20, 18, 20) {real, imag} */,
  {32'hbdb285d0, 32'h3ff4b0c8} /* (20, 18, 19) {real, imag} */,
  {32'hbf83c080, 32'hbddcd040} /* (20, 18, 18) {real, imag} */,
  {32'h3fca50cf, 32'hc04e4561} /* (20, 18, 17) {real, imag} */,
  {32'h3f191c80, 32'hc0169330} /* (20, 18, 16) {real, imag} */,
  {32'h3f5e3dd8, 32'hbf6e7cbd} /* (20, 18, 15) {real, imag} */,
  {32'hbd3f27c0, 32'hbe8e717e} /* (20, 18, 14) {real, imag} */,
  {32'hbf130c22, 32'hbecd8058} /* (20, 18, 13) {real, imag} */,
  {32'h3f0c26d6, 32'h3fc44810} /* (20, 18, 12) {real, imag} */,
  {32'hbfcc8c1e, 32'h3f0fd36c} /* (20, 18, 11) {real, imag} */,
  {32'hc0839b02, 32'hbe259e4c} /* (20, 18, 10) {real, imag} */,
  {32'hbf1f2c5b, 32'hbf348df0} /* (20, 18, 9) {real, imag} */,
  {32'h3fd6a958, 32'hbffa824c} /* (20, 18, 8) {real, imag} */,
  {32'h3fd6a349, 32'hc02f630f} /* (20, 18, 7) {real, imag} */,
  {32'hbe0ece1a, 32'h3db3a820} /* (20, 18, 6) {real, imag} */,
  {32'h3f34e2b0, 32'hbfd8dc43} /* (20, 18, 5) {real, imag} */,
  {32'hc0429cd7, 32'hbfe4ff27} /* (20, 18, 4) {real, imag} */,
  {32'h3f28f653, 32'hbfce1133} /* (20, 18, 3) {real, imag} */,
  {32'h407c01d6, 32'h3fc37d20} /* (20, 18, 2) {real, imag} */,
  {32'hbf9c6c28, 32'h3f81651b} /* (20, 18, 1) {real, imag} */,
  {32'hc021177e, 32'h3f86f131} /* (20, 18, 0) {real, imag} */,
  {32'hbf5ac7f8, 32'hbfafc919} /* (20, 17, 31) {real, imag} */,
  {32'h3e6e1fa0, 32'hbfdca98b} /* (20, 17, 30) {real, imag} */,
  {32'h3faa22e1, 32'hbebea280} /* (20, 17, 29) {real, imag} */,
  {32'h4070e164, 32'hc009b324} /* (20, 17, 28) {real, imag} */,
  {32'h3eda5852, 32'hbf9f0d13} /* (20, 17, 27) {real, imag} */,
  {32'hbfc55797, 32'h40046d8b} /* (20, 17, 26) {real, imag} */,
  {32'h3fbb7976, 32'h3f99b5bf} /* (20, 17, 25) {real, imag} */,
  {32'h3f850b0e, 32'h3ef13d08} /* (20, 17, 24) {real, imag} */,
  {32'hbcb26130, 32'h3dc996c0} /* (20, 17, 23) {real, imag} */,
  {32'h3fc3a806, 32'h3ee86160} /* (20, 17, 22) {real, imag} */,
  {32'h3eb79174, 32'h3e44c8a0} /* (20, 17, 21) {real, imag} */,
  {32'h3f3c58e0, 32'hbf5da951} /* (20, 17, 20) {real, imag} */,
  {32'hbf2b649c, 32'hbf83c554} /* (20, 17, 19) {real, imag} */,
  {32'h3ff7ed0f, 32'hbfa26779} /* (20, 17, 18) {real, imag} */,
  {32'h40635c4a, 32'h3de920c0} /* (20, 17, 17) {real, imag} */,
  {32'hbeeccc58, 32'h4011abc5} /* (20, 17, 16) {real, imag} */,
  {32'hbfd94ba4, 32'hbdfafcf8} /* (20, 17, 15) {real, imag} */,
  {32'hbfe314ce, 32'hbfebf5e9} /* (20, 17, 14) {real, imag} */,
  {32'hbeedef14, 32'hbf1bd42b} /* (20, 17, 13) {real, imag} */,
  {32'h3f8a575a, 32'hbe14d2b0} /* (20, 17, 12) {real, imag} */,
  {32'h3fbb90a6, 32'h3f688835} /* (20, 17, 11) {real, imag} */,
  {32'hbf3467a4, 32'h3fba21c5} /* (20, 17, 10) {real, imag} */,
  {32'hbe2966e4, 32'h3e0066f8} /* (20, 17, 9) {real, imag} */,
  {32'hbe8613d0, 32'h3f980759} /* (20, 17, 8) {real, imag} */,
  {32'h3d922df8, 32'h3edfecee} /* (20, 17, 7) {real, imag} */,
  {32'hbf82d0b4, 32'hc045183a} /* (20, 17, 6) {real, imag} */,
  {32'hbe004144, 32'h3f8d5b76} /* (20, 17, 5) {real, imag} */,
  {32'h3f677b00, 32'h3f617564} /* (20, 17, 4) {real, imag} */,
  {32'h3f913815, 32'h3ec86df4} /* (20, 17, 3) {real, imag} */,
  {32'h3fbf2f5d, 32'h3fc0cb3d} /* (20, 17, 2) {real, imag} */,
  {32'h4026d968, 32'h3f5ed6e4} /* (20, 17, 1) {real, imag} */,
  {32'h3f8244bc, 32'hbe883429} /* (20, 17, 0) {real, imag} */,
  {32'hbeba3b98, 32'hbf8032c6} /* (20, 16, 31) {real, imag} */,
  {32'hbed6d730, 32'hbf38bda4} /* (20, 16, 30) {real, imag} */,
  {32'h4010a3e2, 32'hbf02fd34} /* (20, 16, 29) {real, imag} */,
  {32'h4000aea1, 32'h3f961ca4} /* (20, 16, 28) {real, imag} */,
  {32'hbd100178, 32'h3f9d97b2} /* (20, 16, 27) {real, imag} */,
  {32'hbe5ffdf0, 32'hbf219e00} /* (20, 16, 26) {real, imag} */,
  {32'h3ec78a40, 32'hbfdef038} /* (20, 16, 25) {real, imag} */,
  {32'h3f4c65a4, 32'h3fbaebd2} /* (20, 16, 24) {real, imag} */,
  {32'h3e8db798, 32'h402626c8} /* (20, 16, 23) {real, imag} */,
  {32'hbf1703a8, 32'h40058bd4} /* (20, 16, 22) {real, imag} */,
  {32'h3f611362, 32'h3f577e58} /* (20, 16, 21) {real, imag} */,
  {32'h3c45da00, 32'hbe804d20} /* (20, 16, 20) {real, imag} */,
  {32'h3eeb74f0, 32'hbfa5d2e4} /* (20, 16, 19) {real, imag} */,
  {32'h3f9d7d5c, 32'hc0125a14} /* (20, 16, 18) {real, imag} */,
  {32'hbf219774, 32'hbf924115} /* (20, 16, 17) {real, imag} */,
  {32'hbf8a2376, 32'h3fb7f11a} /* (20, 16, 16) {real, imag} */,
  {32'h3f7ab6cb, 32'hbf9820aa} /* (20, 16, 15) {real, imag} */,
  {32'h4034d6d4, 32'hbfc12fd4} /* (20, 16, 14) {real, imag} */,
  {32'h3f299528, 32'hc00664aa} /* (20, 16, 13) {real, imag} */,
  {32'hc007f900, 32'hbf046360} /* (20, 16, 12) {real, imag} */,
  {32'hbfc3eef8, 32'hbe4f27c0} /* (20, 16, 11) {real, imag} */,
  {32'hc045e05c, 32'hbf7dcaf0} /* (20, 16, 10) {real, imag} */,
  {32'hbfebdaf0, 32'h3f58acd6} /* (20, 16, 9) {real, imag} */,
  {32'hbfd2abae, 32'h3d57c5a0} /* (20, 16, 8) {real, imag} */,
  {32'hbf4e0916, 32'h3f6e5106} /* (20, 16, 7) {real, imag} */,
  {32'h40075134, 32'h400ddc05} /* (20, 16, 6) {real, imag} */,
  {32'h3f831d0e, 32'h3fe50bb4} /* (20, 16, 5) {real, imag} */,
  {32'h3f6bc010, 32'h3fe734d4} /* (20, 16, 4) {real, imag} */,
  {32'h4004f2ec, 32'h3fd697d6} /* (20, 16, 3) {real, imag} */,
  {32'h3fb28338, 32'hbfd05d54} /* (20, 16, 2) {real, imag} */,
  {32'h3f0ea8dc, 32'h3ed7f904} /* (20, 16, 1) {real, imag} */,
  {32'hbf8babd8, 32'hbf7b9e0c} /* (20, 16, 0) {real, imag} */,
  {32'hbe8d19e0, 32'h3ffceb39} /* (20, 15, 31) {real, imag} */,
  {32'hbfa2562c, 32'h3ffc302b} /* (20, 15, 30) {real, imag} */,
  {32'hbfcc6379, 32'h3f0ea1b0} /* (20, 15, 29) {real, imag} */,
  {32'hbf05c462, 32'h3fada425} /* (20, 15, 28) {real, imag} */,
  {32'h3f3304e9, 32'h401b5e92} /* (20, 15, 27) {real, imag} */,
  {32'hbec24128, 32'hbe0b0590} /* (20, 15, 26) {real, imag} */,
  {32'hc003c841, 32'hbfa9bb5f} /* (20, 15, 25) {real, imag} */,
  {32'hbff6dd7a, 32'hbf3654d4} /* (20, 15, 24) {real, imag} */,
  {32'hbf402092, 32'hbf0a2c40} /* (20, 15, 23) {real, imag} */,
  {32'hbf92b206, 32'hbf3f8a98} /* (20, 15, 22) {real, imag} */,
  {32'hbfae0777, 32'h3fc6f99b} /* (20, 15, 21) {real, imag} */,
  {32'hbfe36ed8, 32'h402f2d44} /* (20, 15, 20) {real, imag} */,
  {32'hc01b0b1d, 32'h3ee06b62} /* (20, 15, 19) {real, imag} */,
  {32'hbd8c3390, 32'h3e37f548} /* (20, 15, 18) {real, imag} */,
  {32'h408d3450, 32'hbdabfd40} /* (20, 15, 17) {real, imag} */,
  {32'h4045b255, 32'hc0025589} /* (20, 15, 16) {real, imag} */,
  {32'hbff7147a, 32'hbfab97de} /* (20, 15, 15) {real, imag} */,
  {32'hbf876436, 32'hbf11e206} /* (20, 15, 14) {real, imag} */,
  {32'h3fe7aec9, 32'hbedc7f7a} /* (20, 15, 13) {real, imag} */,
  {32'h3fa6afd2, 32'hbfebe16f} /* (20, 15, 12) {real, imag} */,
  {32'h3fa34d1e, 32'hbf2ea87d} /* (20, 15, 11) {real, imag} */,
  {32'h3fc19022, 32'h3f525e76} /* (20, 15, 10) {real, imag} */,
  {32'h3f5ecd1b, 32'h40380b02} /* (20, 15, 9) {real, imag} */,
  {32'hc0008ffe, 32'h40358726} /* (20, 15, 8) {real, imag} */,
  {32'hbfc24a88, 32'hbf70782f} /* (20, 15, 7) {real, imag} */,
  {32'h3f241c98, 32'hbfdfedfb} /* (20, 15, 6) {real, imag} */,
  {32'h3f5b88d5, 32'hbd61eb40} /* (20, 15, 5) {real, imag} */,
  {32'hbf93e460, 32'h40a099fc} /* (20, 15, 4) {real, imag} */,
  {32'hbf5694e6, 32'h406140fe} /* (20, 15, 3) {real, imag} */,
  {32'h3fd482df, 32'h3f4b3086} /* (20, 15, 2) {real, imag} */,
  {32'h3fcecab8, 32'h3e9bbd29} /* (20, 15, 1) {real, imag} */,
  {32'h3fc36ee4, 32'h3e2ec212} /* (20, 15, 0) {real, imag} */,
  {32'h3fb4227c, 32'hbf67e160} /* (20, 14, 31) {real, imag} */,
  {32'hbeb57c1a, 32'hbff85125} /* (20, 14, 30) {real, imag} */,
  {32'h3ff88360, 32'hc06bc46f} /* (20, 14, 29) {real, imag} */,
  {32'h401de46c, 32'hbeb171c0} /* (20, 14, 28) {real, imag} */,
  {32'h3f9d9450, 32'hbe2848d0} /* (20, 14, 27) {real, imag} */,
  {32'hbecfc30c, 32'hbf16c3a8} /* (20, 14, 26) {real, imag} */,
  {32'h3f931c8f, 32'h3fdd68aa} /* (20, 14, 25) {real, imag} */,
  {32'hbe961568, 32'h40465fb6} /* (20, 14, 24) {real, imag} */,
  {32'hbe2a8338, 32'h3feca35d} /* (20, 14, 23) {real, imag} */,
  {32'h3ff9b907, 32'h3f6dd0d4} /* (20, 14, 22) {real, imag} */,
  {32'hbef0e860, 32'h3f834b1d} /* (20, 14, 21) {real, imag} */,
  {32'hc051f373, 32'hc0463369} /* (20, 14, 20) {real, imag} */,
  {32'hbfa250b9, 32'hc0581c20} /* (20, 14, 19) {real, imag} */,
  {32'h3fa99432, 32'hbfa244a8} /* (20, 14, 18) {real, imag} */,
  {32'hbf907437, 32'hbf991d2a} /* (20, 14, 17) {real, imag} */,
  {32'hc05c7b48, 32'h400b69c8} /* (20, 14, 16) {real, imag} */,
  {32'hbe94a430, 32'hbeb5b722} /* (20, 14, 15) {real, imag} */,
  {32'hbfcd05fb, 32'hc00d80c3} /* (20, 14, 14) {real, imag} */,
  {32'hbf164056, 32'hbfcc12b2} /* (20, 14, 13) {real, imag} */,
  {32'h40271cdc, 32'h3ec52260} /* (20, 14, 12) {real, imag} */,
  {32'h3f1c0534, 32'h3f33923c} /* (20, 14, 11) {real, imag} */,
  {32'h3faacf38, 32'hbf31557b} /* (20, 14, 10) {real, imag} */,
  {32'h4022bd17, 32'h40067e0c} /* (20, 14, 9) {real, imag} */,
  {32'h3ffc04ac, 32'hc03b41e6} /* (20, 14, 8) {real, imag} */,
  {32'h40114814, 32'hbffacee2} /* (20, 14, 7) {real, imag} */,
  {32'h3ded1b74, 32'hbee8e058} /* (20, 14, 6) {real, imag} */,
  {32'hbf2ae5e8, 32'hbf593cda} /* (20, 14, 5) {real, imag} */,
  {32'hbf9635de, 32'hbf2bdd82} /* (20, 14, 4) {real, imag} */,
  {32'hbf3b7ca3, 32'hbf655ca2} /* (20, 14, 3) {real, imag} */,
  {32'hbe5b1e00, 32'hbe064f1c} /* (20, 14, 2) {real, imag} */,
  {32'h400ea814, 32'hbfd6322f} /* (20, 14, 1) {real, imag} */,
  {32'h3fa3b64c, 32'hbecf4893} /* (20, 14, 0) {real, imag} */,
  {32'h3f86944e, 32'hbfa7437c} /* (20, 13, 31) {real, imag} */,
  {32'h3f2ac490, 32'hbfcaf625} /* (20, 13, 30) {real, imag} */,
  {32'hbf39adfc, 32'h3dc54b58} /* (20, 13, 29) {real, imag} */,
  {32'hbf3bff1e, 32'h3ff33c4c} /* (20, 13, 28) {real, imag} */,
  {32'h40039de8, 32'h404e351c} /* (20, 13, 27) {real, imag} */,
  {32'h3fecfc5e, 32'h4072c5c8} /* (20, 13, 26) {real, imag} */,
  {32'h3da8d980, 32'hbfb69cd1} /* (20, 13, 25) {real, imag} */,
  {32'hbfca3910, 32'h3e3e5478} /* (20, 13, 24) {real, imag} */,
  {32'h3b8a5a80, 32'h403a6970} /* (20, 13, 23) {real, imag} */,
  {32'h3f7e2ece, 32'h40a078f3} /* (20, 13, 22) {real, imag} */,
  {32'h3e682d60, 32'h406b1f79} /* (20, 13, 21) {real, imag} */,
  {32'hbd72df80, 32'h3ec481f0} /* (20, 13, 20) {real, imag} */,
  {32'h3fe2dba8, 32'hbff8db80} /* (20, 13, 19) {real, imag} */,
  {32'h3d60ddf0, 32'hbfa336b2} /* (20, 13, 18) {real, imag} */,
  {32'hc017f439, 32'h3f18df04} /* (20, 13, 17) {real, imag} */,
  {32'h3fd2a4a2, 32'h3e5f1958} /* (20, 13, 16) {real, imag} */,
  {32'h3fb3cf09, 32'hbfdcb773} /* (20, 13, 15) {real, imag} */,
  {32'hc006fae8, 32'hbeb51d68} /* (20, 13, 14) {real, imag} */,
  {32'hbf154630, 32'h4028e665} /* (20, 13, 13) {real, imag} */,
  {32'hc02c8a76, 32'h3ffb77b8} /* (20, 13, 12) {real, imag} */,
  {32'hc05210f2, 32'h409308af} /* (20, 13, 11) {real, imag} */,
  {32'h3cce8400, 32'h40cb8dac} /* (20, 13, 10) {real, imag} */,
  {32'h3f9ad473, 32'h3ff1a7a2} /* (20, 13, 9) {real, imag} */,
  {32'hbe68aa60, 32'hc0137c6b} /* (20, 13, 8) {real, imag} */,
  {32'hbf89febc, 32'hbe004760} /* (20, 13, 7) {real, imag} */,
  {32'hc00e744c, 32'h3ee5b918} /* (20, 13, 6) {real, imag} */,
  {32'hc06a663b, 32'hbdf8f130} /* (20, 13, 5) {real, imag} */,
  {32'hc0481920, 32'hbe96c440} /* (20, 13, 4) {real, imag} */,
  {32'h40420eac, 32'hbfcd2cce} /* (20, 13, 3) {real, imag} */,
  {32'h40875a98, 32'hbef8dbd4} /* (20, 13, 2) {real, imag} */,
  {32'h3fb1099c, 32'h3ff6fe16} /* (20, 13, 1) {real, imag} */,
  {32'h3fc0d843, 32'h3f116776} /* (20, 13, 0) {real, imag} */,
  {32'h401a6744, 32'h3f8c75b9} /* (20, 12, 31) {real, imag} */,
  {32'h40d5c5da, 32'hbe855500} /* (20, 12, 30) {real, imag} */,
  {32'h409a539e, 32'h4041fcc0} /* (20, 12, 29) {real, imag} */,
  {32'hbeb1eb3c, 32'h40727e98} /* (20, 12, 28) {real, imag} */,
  {32'h40005975, 32'hbddb3b70} /* (20, 12, 27) {real, imag} */,
  {32'h3fed4b72, 32'h3d94f740} /* (20, 12, 26) {real, imag} */,
  {32'hc0619db8, 32'hc073abbf} /* (20, 12, 25) {real, imag} */,
  {32'hc025c854, 32'hc0dd748d} /* (20, 12, 24) {real, imag} */,
  {32'hbdb25e40, 32'hbf60476c} /* (20, 12, 23) {real, imag} */,
  {32'h4021c12f, 32'h403a71db} /* (20, 12, 22) {real, imag} */,
  {32'h3f8d6836, 32'hbfbd4fb7} /* (20, 12, 21) {real, imag} */,
  {32'hc0229f7a, 32'h401193a0} /* (20, 12, 20) {real, imag} */,
  {32'hc0919c46, 32'h3dd885d0} /* (20, 12, 19) {real, imag} */,
  {32'hc00107dd, 32'hc09e1e21} /* (20, 12, 18) {real, imag} */,
  {32'hbf0963f3, 32'hc00dda60} /* (20, 12, 17) {real, imag} */,
  {32'hc024f4a0, 32'h3f411a7c} /* (20, 12, 16) {real, imag} */,
  {32'hc0118916, 32'h3f9c037c} /* (20, 12, 15) {real, imag} */,
  {32'hbee9af4c, 32'h3f350f42} /* (20, 12, 14) {real, imag} */,
  {32'h3fe1a2ca, 32'h3fa10ab8} /* (20, 12, 13) {real, imag} */,
  {32'hbfb48bc4, 32'h3f3de14a} /* (20, 12, 12) {real, imag} */,
  {32'h3e17e990, 32'hbfb0e755} /* (20, 12, 11) {real, imag} */,
  {32'h404b236c, 32'hc089babe} /* (20, 12, 10) {real, imag} */,
  {32'h3fbc8dfe, 32'hc0294da8} /* (20, 12, 9) {real, imag} */,
  {32'h3fa5d83a, 32'hbe9dcf28} /* (20, 12, 8) {real, imag} */,
  {32'hbe7d2e56, 32'h3f4ba406} /* (20, 12, 7) {real, imag} */,
  {32'hc055131b, 32'hc001cd0b} /* (20, 12, 6) {real, imag} */,
  {32'hbeb0547c, 32'hc06af824} /* (20, 12, 5) {real, imag} */,
  {32'hbfb09adb, 32'h3e656b6e} /* (20, 12, 4) {real, imag} */,
  {32'hbfd7e566, 32'h3fcfed3b} /* (20, 12, 3) {real, imag} */,
  {32'hbf9ea304, 32'h3fa39c66} /* (20, 12, 2) {real, imag} */,
  {32'hbe41c380, 32'h40384ea1} /* (20, 12, 1) {real, imag} */,
  {32'h3ef7d1ea, 32'h3f46f71a} /* (20, 12, 0) {real, imag} */,
  {32'h3f7a8b3e, 32'h3ffc6a62} /* (20, 11, 31) {real, imag} */,
  {32'h3efb66bc, 32'h403b9f64} /* (20, 11, 30) {real, imag} */,
  {32'h4015923f, 32'hbebe26a0} /* (20, 11, 29) {real, imag} */,
  {32'hbe23886c, 32'hc09814f1} /* (20, 11, 28) {real, imag} */,
  {32'hbc666bc0, 32'h3d63fc80} /* (20, 11, 27) {real, imag} */,
  {32'hbdb967a8, 32'hbea739fa} /* (20, 11, 26) {real, imag} */,
  {32'h3f5e3a1e, 32'hbf7a618c} /* (20, 11, 25) {real, imag} */,
  {32'hbe8b71e6, 32'h400f27d4} /* (20, 11, 24) {real, imag} */,
  {32'hc08dfb36, 32'h3e9a4068} /* (20, 11, 23) {real, imag} */,
  {32'hc0232236, 32'h3ea78158} /* (20, 11, 22) {real, imag} */,
  {32'h3e83a3a4, 32'h3c3a1e80} /* (20, 11, 21) {real, imag} */,
  {32'hbe8e52e8, 32'hc09ee8c0} /* (20, 11, 20) {real, imag} */,
  {32'h401339d0, 32'hbe99e504} /* (20, 11, 19) {real, imag} */,
  {32'h409331d0, 32'h40ea0584} /* (20, 11, 18) {real, imag} */,
  {32'h3e8f78c6, 32'h40e9e6ec} /* (20, 11, 17) {real, imag} */,
  {32'hbd8dd870, 32'h4023f424} /* (20, 11, 16) {real, imag} */,
  {32'h402675d8, 32'hbfd3079c} /* (20, 11, 15) {real, imag} */,
  {32'hbe6952a8, 32'h3e8ea994} /* (20, 11, 14) {real, imag} */,
  {32'hc090adb3, 32'h400e9949} /* (20, 11, 13) {real, imag} */,
  {32'hc0589d68, 32'h3fb3b388} /* (20, 11, 12) {real, imag} */,
  {32'hc04544b8, 32'hbfc1c8dd} /* (20, 11, 11) {real, imag} */,
  {32'hc000a043, 32'h3d6b2980} /* (20, 11, 10) {real, imag} */,
  {32'h4013e354, 32'hbea85aec} /* (20, 11, 9) {real, imag} */,
  {32'h402eda64, 32'h3fa4becd} /* (20, 11, 8) {real, imag} */,
  {32'h3fabaf5a, 32'hbf0ccb6c} /* (20, 11, 7) {real, imag} */,
  {32'hbfd9136a, 32'hc078b5a0} /* (20, 11, 6) {real, imag} */,
  {32'hc0016813, 32'h3f404ff4} /* (20, 11, 5) {real, imag} */,
  {32'h3fd5a932, 32'h3e97b2a6} /* (20, 11, 4) {real, imag} */,
  {32'hbe3353e0, 32'hc08bca35} /* (20, 11, 3) {real, imag} */,
  {32'h4008a2fa, 32'hbf6c02f4} /* (20, 11, 2) {real, imag} */,
  {32'h406d555d, 32'hbca70500} /* (20, 11, 1) {real, imag} */,
  {32'h4000b1d8, 32'h3f228936} /* (20, 11, 0) {real, imag} */,
  {32'h3dca06e0, 32'hbe2a0848} /* (20, 10, 31) {real, imag} */,
  {32'hbf816f4c, 32'h3fc43dbe} /* (20, 10, 30) {real, imag} */,
  {32'hbe62fda4, 32'hbed51a9c} /* (20, 10, 29) {real, imag} */,
  {32'h3f90196b, 32'hc0304064} /* (20, 10, 28) {real, imag} */,
  {32'hbfa7b635, 32'hbd840370} /* (20, 10, 27) {real, imag} */,
  {32'h3d4ef300, 32'hc04ef21b} /* (20, 10, 26) {real, imag} */,
  {32'hbf37efee, 32'h3e6d2cd0} /* (20, 10, 25) {real, imag} */,
  {32'h3ff1d3c2, 32'hbe62aa70} /* (20, 10, 24) {real, imag} */,
  {32'h3fba7fb7, 32'hc09b7b96} /* (20, 10, 23) {real, imag} */,
  {32'hbf9b7c27, 32'hc08dc7f6} /* (20, 10, 22) {real, imag} */,
  {32'hc093b660, 32'h403dfcca} /* (20, 10, 21) {real, imag} */,
  {32'h3e90e744, 32'h4090541f} /* (20, 10, 20) {real, imag} */,
  {32'h4040b6b8, 32'h40757982} /* (20, 10, 19) {real, imag} */,
  {32'h409fba87, 32'h4002a0f6} /* (20, 10, 18) {real, imag} */,
  {32'h40dc7522, 32'h40858fb4} /* (20, 10, 17) {real, imag} */,
  {32'h4072959d, 32'hbecc7322} /* (20, 10, 16) {real, imag} */,
  {32'h3fbf3a20, 32'hbfe986ce} /* (20, 10, 15) {real, imag} */,
  {32'h4013339a, 32'hc09267fc} /* (20, 10, 14) {real, imag} */,
  {32'h3eeebe68, 32'hc086df12} /* (20, 10, 13) {real, imag} */,
  {32'h3ea6889a, 32'hc0a0e59b} /* (20, 10, 12) {real, imag} */,
  {32'h3f665978, 32'h3eef5e68} /* (20, 10, 11) {real, imag} */,
  {32'hc02ad314, 32'h3fe750dc} /* (20, 10, 10) {real, imag} */,
  {32'hc0e35d1c, 32'h3fe9f0ec} /* (20, 10, 9) {real, imag} */,
  {32'hc0d6692a, 32'h3f8951da} /* (20, 10, 8) {real, imag} */,
  {32'hc000a80c, 32'hbdd3def0} /* (20, 10, 7) {real, imag} */,
  {32'h3f8d8a36, 32'hbfc6d18a} /* (20, 10, 6) {real, imag} */,
  {32'hbfba28ac, 32'hc0682725} /* (20, 10, 5) {real, imag} */,
  {32'hc02e4d0c, 32'hc0c3b1fc} /* (20, 10, 4) {real, imag} */,
  {32'hc0884b80, 32'hc12f9852} /* (20, 10, 3) {real, imag} */,
  {32'hbfb38b59, 32'hc0f751e8} /* (20, 10, 2) {real, imag} */,
  {32'h4013c256, 32'h3f8dc3be} /* (20, 10, 1) {real, imag} */,
  {32'h4010d7e8, 32'hbe820ef4} /* (20, 10, 0) {real, imag} */,
  {32'hbd5298c0, 32'hc0173a1a} /* (20, 9, 31) {real, imag} */,
  {32'h3f8608f4, 32'h3e80e500} /* (20, 9, 30) {real, imag} */,
  {32'hbfaba476, 32'h4052e5ec} /* (20, 9, 29) {real, imag} */,
  {32'hc031aa3a, 32'h405447b8} /* (20, 9, 28) {real, imag} */,
  {32'h3dc7cbb8, 32'h400147f0} /* (20, 9, 27) {real, imag} */,
  {32'hc024412e, 32'hc0076608} /* (20, 9, 26) {real, imag} */,
  {32'h3d2ca960, 32'hc018b0c5} /* (20, 9, 25) {real, imag} */,
  {32'h3ff73392, 32'hbe0047d0} /* (20, 9, 24) {real, imag} */,
  {32'h405ed828, 32'hc0390cc5} /* (20, 9, 23) {real, imag} */,
  {32'h40330da8, 32'hc0a34136} /* (20, 9, 22) {real, imag} */,
  {32'h3ef77578, 32'hbfe924ee} /* (20, 9, 21) {real, imag} */,
  {32'h40175018, 32'hc0daf999} /* (20, 9, 20) {real, imag} */,
  {32'h4084c400, 32'hc013fd2c} /* (20, 9, 19) {real, imag} */,
  {32'h403aa62b, 32'hc08d7a06} /* (20, 9, 18) {real, imag} */,
  {32'hc02b5315, 32'hc0b7e7cd} /* (20, 9, 17) {real, imag} */,
  {32'hc07ad18c, 32'hbfb73123} /* (20, 9, 16) {real, imag} */,
  {32'hbfe463e6, 32'hbfcdfbcd} /* (20, 9, 15) {real, imag} */,
  {32'h3fcb7e35, 32'h4088d8ba} /* (20, 9, 14) {real, imag} */,
  {32'h3ff113ce, 32'h400c0da0} /* (20, 9, 13) {real, imag} */,
  {32'h3fccac10, 32'hc00dbd5e} /* (20, 9, 12) {real, imag} */,
  {32'hbf06fe58, 32'hc011e142} /* (20, 9, 11) {real, imag} */,
  {32'hc0a450e1, 32'hc0d29e58} /* (20, 9, 10) {real, imag} */,
  {32'hc100b7c0, 32'h3f8184a8} /* (20, 9, 9) {real, imag} */,
  {32'hc0f2ec4f, 32'h3e17fdf8} /* (20, 9, 8) {real, imag} */,
  {32'hc0ab19c0, 32'h3fa458b2} /* (20, 9, 7) {real, imag} */,
  {32'h3f8e1d20, 32'hbe70d58c} /* (20, 9, 6) {real, imag} */,
  {32'h3f80ed6c, 32'hc0ae870c} /* (20, 9, 5) {real, imag} */,
  {32'hc07a7a2a, 32'h3d0c29a0} /* (20, 9, 4) {real, imag} */,
  {32'hc0603bfe, 32'h40bd00e2} /* (20, 9, 3) {real, imag} */,
  {32'hc097d191, 32'h3fd163d1} /* (20, 9, 2) {real, imag} */,
  {32'hc099147c, 32'hbfdb6a38} /* (20, 9, 1) {real, imag} */,
  {32'hbf108d84, 32'hbea97143} /* (20, 9, 0) {real, imag} */,
  {32'hc0749eb5, 32'hbed5c5b0} /* (20, 8, 31) {real, imag} */,
  {32'h3ffbd316, 32'h3fbcca4c} /* (20, 8, 30) {real, imag} */,
  {32'h400dd209, 32'hc075210f} /* (20, 8, 29) {real, imag} */,
  {32'hbf94eb34, 32'hbe356a14} /* (20, 8, 28) {real, imag} */,
  {32'h408ae178, 32'h3ee47893} /* (20, 8, 27) {real, imag} */,
  {32'h40507a69, 32'h3f86969c} /* (20, 8, 26) {real, imag} */,
  {32'h40e66f70, 32'h406878b5} /* (20, 8, 25) {real, imag} */,
  {32'h411ca77a, 32'h3e849000} /* (20, 8, 24) {real, imag} */,
  {32'h406a73a8, 32'h3f74fcc2} /* (20, 8, 23) {real, imag} */,
  {32'h40b4f6ec, 32'h3eeee608} /* (20, 8, 22) {real, imag} */,
  {32'hbf320834, 32'hc01fe7af} /* (20, 8, 21) {real, imag} */,
  {32'hbfd8efba, 32'hc055202e} /* (20, 8, 20) {real, imag} */,
  {32'hbffacd0a, 32'hc0c3f844} /* (20, 8, 19) {real, imag} */,
  {32'h400cfc1c, 32'h4068a373} /* (20, 8, 18) {real, imag} */,
  {32'h407e8904, 32'hbffa3038} /* (20, 8, 17) {real, imag} */,
  {32'h3fc0b4fb, 32'hc11ba5a4} /* (20, 8, 16) {real, imag} */,
  {32'h400425e1, 32'h3edb8968} /* (20, 8, 15) {real, imag} */,
  {32'hbf727aca, 32'h40e13b48} /* (20, 8, 14) {real, imag} */,
  {32'h3f90b950, 32'h407ae336} /* (20, 8, 13) {real, imag} */,
  {32'h40e8663a, 32'h402d1c22} /* (20, 8, 12) {real, imag} */,
  {32'h4122fba9, 32'hbfb51a82} /* (20, 8, 11) {real, imag} */,
  {32'h3ecc9236, 32'hc0f3f7a2} /* (20, 8, 10) {real, imag} */,
  {32'hc0bcc299, 32'hbf907cd6} /* (20, 8, 9) {real, imag} */,
  {32'hbe3c3780, 32'hbdb76f10} /* (20, 8, 8) {real, imag} */,
  {32'h3fd7f3f3, 32'h3e8f3a36} /* (20, 8, 7) {real, imag} */,
  {32'h4063ea16, 32'h410e3058} /* (20, 8, 6) {real, imag} */,
  {32'h408086eb, 32'h40c1953b} /* (20, 8, 5) {real, imag} */,
  {32'h4003bff4, 32'h3fc30056} /* (20, 8, 4) {real, imag} */,
  {32'h4008a32d, 32'h402c690e} /* (20, 8, 3) {real, imag} */,
  {32'h404e9171, 32'h3fdeb802} /* (20, 8, 2) {real, imag} */,
  {32'h3fb951dd, 32'hc08c1196} /* (20, 8, 1) {real, imag} */,
  {32'hbfa08ef6, 32'hc0ed3cd3} /* (20, 8, 0) {real, imag} */,
  {32'hbff2851a, 32'hbffb9fc0} /* (20, 7, 31) {real, imag} */,
  {32'hc0d6ac4a, 32'hc02b9853} /* (20, 7, 30) {real, imag} */,
  {32'hc07ef352, 32'h4003c6d0} /* (20, 7, 29) {real, imag} */,
  {32'hc003bde4, 32'hbf9d952c} /* (20, 7, 28) {real, imag} */,
  {32'h40543082, 32'hc11346b8} /* (20, 7, 27) {real, imag} */,
  {32'hc032f98d, 32'hc0dd23e6} /* (20, 7, 26) {real, imag} */,
  {32'hc092269d, 32'hbf760194} /* (20, 7, 25) {real, imag} */,
  {32'hc0e2b17e, 32'h3f9d9826} /* (20, 7, 24) {real, imag} */,
  {32'hc02f38be, 32'h40902c78} /* (20, 7, 23) {real, imag} */,
  {32'hc07f4e52, 32'h4000834c} /* (20, 7, 22) {real, imag} */,
  {32'hc0267546, 32'hc033ff90} /* (20, 7, 21) {real, imag} */,
  {32'hc0b4c662, 32'hbc56d580} /* (20, 7, 20) {real, imag} */,
  {32'hc0ca525c, 32'h4080ddd6} /* (20, 7, 19) {real, imag} */,
  {32'hc0ddb5b8, 32'h3f57fb84} /* (20, 7, 18) {real, imag} */,
  {32'hc0b92f64, 32'hc0dc1743} /* (20, 7, 17) {real, imag} */,
  {32'h400ab648, 32'hc0dd2750} /* (20, 7, 16) {real, imag} */,
  {32'h40ceadf5, 32'hc0288ffe} /* (20, 7, 15) {real, imag} */,
  {32'h40b71e68, 32'hc0ada03a} /* (20, 7, 14) {real, imag} */,
  {32'hc050a295, 32'hbf3cc5e7} /* (20, 7, 13) {real, imag} */,
  {32'hc01b5aab, 32'h40a61694} /* (20, 7, 12) {real, imag} */,
  {32'h3fcb0178, 32'hbfacd126} /* (20, 7, 11) {real, imag} */,
  {32'h3fbe77f2, 32'hc09adf23} /* (20, 7, 10) {real, imag} */,
  {32'hbe14ff50, 32'hbfba543c} /* (20, 7, 9) {real, imag} */,
  {32'hc0e2a41c, 32'h3f256dec} /* (20, 7, 8) {real, imag} */,
  {32'hbf7e9467, 32'hbddde440} /* (20, 7, 7) {real, imag} */,
  {32'h3fa3ff0c, 32'hc0794e92} /* (20, 7, 6) {real, imag} */,
  {32'h4095ef50, 32'hbe9b90b2} /* (20, 7, 5) {real, imag} */,
  {32'h40c66d46, 32'h40bda0ff} /* (20, 7, 4) {real, imag} */,
  {32'h40a9bdb6, 32'h40d30a36} /* (20, 7, 3) {real, imag} */,
  {32'h406d4df5, 32'hbd0330e0} /* (20, 7, 2) {real, imag} */,
  {32'h3fd43b93, 32'hc055719c} /* (20, 7, 1) {real, imag} */,
  {32'h3e14abc8, 32'h4011fe9e} /* (20, 7, 0) {real, imag} */,
  {32'hbfa2d4a8, 32'hc0397940} /* (20, 6, 31) {real, imag} */,
  {32'hbeaf8474, 32'hc0c0fac7} /* (20, 6, 30) {real, imag} */,
  {32'hc0088569, 32'hc0e1189f} /* (20, 6, 29) {real, imag} */,
  {32'hc0985c51, 32'hc09e0017} /* (20, 6, 28) {real, imag} */,
  {32'hc03e2768, 32'hc0136c90} /* (20, 6, 27) {real, imag} */,
  {32'hc0de90b8, 32'hc02b89f6} /* (20, 6, 26) {real, imag} */,
  {32'hc0af5076, 32'hc010227b} /* (20, 6, 25) {real, imag} */,
  {32'h3f8f7eca, 32'h406a6c29} /* (20, 6, 24) {real, imag} */,
  {32'h403e81d0, 32'h413062bc} /* (20, 6, 23) {real, imag} */,
  {32'h3f964b5c, 32'h40b004d6} /* (20, 6, 22) {real, imag} */,
  {32'hc035f820, 32'hc0b70498} /* (20, 6, 21) {real, imag} */,
  {32'h40681f4c, 32'hc042eb4d} /* (20, 6, 20) {real, imag} */,
  {32'h404898bb, 32'h4010630f} /* (20, 6, 19) {real, imag} */,
  {32'hbfeda2b5, 32'h3fae0684} /* (20, 6, 18) {real, imag} */,
  {32'hc0f254a0, 32'h40ce80a7} /* (20, 6, 17) {real, imag} */,
  {32'hc0b0f298, 32'h40a48015} /* (20, 6, 16) {real, imag} */,
  {32'hbf8e62e0, 32'h40938647} /* (20, 6, 15) {real, imag} */,
  {32'h408bc0d4, 32'h3dd3eb40} /* (20, 6, 14) {real, imag} */,
  {32'h411d7328, 32'hc0ed50aa} /* (20, 6, 13) {real, imag} */,
  {32'h402b38fd, 32'hbffa0689} /* (20, 6, 12) {real, imag} */,
  {32'hbfd819e6, 32'hc0993e42} /* (20, 6, 11) {real, imag} */,
  {32'h403810c2, 32'hc02149cd} /* (20, 6, 10) {real, imag} */,
  {32'h4106b5e9, 32'hc0a308c3} /* (20, 6, 9) {real, imag} */,
  {32'h40d462eb, 32'hc05c2e32} /* (20, 6, 8) {real, imag} */,
  {32'h40bdb610, 32'h40b15359} /* (20, 6, 7) {real, imag} */,
  {32'hbfaa9482, 32'h4146b319} /* (20, 6, 6) {real, imag} */,
  {32'hbce46000, 32'h402a332c} /* (20, 6, 5) {real, imag} */,
  {32'hc07db888, 32'hbf100fee} /* (20, 6, 4) {real, imag} */,
  {32'hc0e58a32, 32'hbf67f36c} /* (20, 6, 3) {real, imag} */,
  {32'hc0655abc, 32'hbf1411a6} /* (20, 6, 2) {real, imag} */,
  {32'hbffed50e, 32'hbe98b678} /* (20, 6, 1) {real, imag} */,
  {32'h3fb3d0e9, 32'hc0277f8a} /* (20, 6, 0) {real, imag} */,
  {32'hbfe5706f, 32'h4000f48d} /* (20, 5, 31) {real, imag} */,
  {32'h409a22c8, 32'h40005f11} /* (20, 5, 30) {real, imag} */,
  {32'h412f6290, 32'hc054fb72} /* (20, 5, 29) {real, imag} */,
  {32'h40e1c810, 32'hbf8e5d5c} /* (20, 5, 28) {real, imag} */,
  {32'h40821777, 32'h3ff00588} /* (20, 5, 27) {real, imag} */,
  {32'h3ffcc4f6, 32'h40989cb6} /* (20, 5, 26) {real, imag} */,
  {32'h40914435, 32'h414019ff} /* (20, 5, 25) {real, imag} */,
  {32'h3ff213d2, 32'h40bf32b5} /* (20, 5, 24) {real, imag} */,
  {32'h403d5714, 32'hc0f2fed4} /* (20, 5, 23) {real, imag} */,
  {32'h402d5f32, 32'hc08f41b2} /* (20, 5, 22) {real, imag} */,
  {32'hc02ea9e8, 32'h400bbabc} /* (20, 5, 21) {real, imag} */,
  {32'hc0305a4a, 32'hc0ebc679} /* (20, 5, 20) {real, imag} */,
  {32'h40165e65, 32'hc0aa360e} /* (20, 5, 19) {real, imag} */,
  {32'h3ef8bb1e, 32'h3eeecf60} /* (20, 5, 18) {real, imag} */,
  {32'h404b4665, 32'h3f534200} /* (20, 5, 17) {real, imag} */,
  {32'hc0ad11ee, 32'hbf58f1d8} /* (20, 5, 16) {real, imag} */,
  {32'hbf9a5228, 32'h3dc16720} /* (20, 5, 15) {real, imag} */,
  {32'h40949769, 32'h401eec61} /* (20, 5, 14) {real, imag} */,
  {32'hc00d3e18, 32'hbd88d2fc} /* (20, 5, 13) {real, imag} */,
  {32'hc09b86c9, 32'hc0697602} /* (20, 5, 12) {real, imag} */,
  {32'hc0077518, 32'h3f766288} /* (20, 5, 11) {real, imag} */,
  {32'hc0861f3a, 32'h40db84fc} /* (20, 5, 10) {real, imag} */,
  {32'hbf9e65f6, 32'hc0881820} /* (20, 5, 9) {real, imag} */,
  {32'h3ef7379a, 32'hc1118c3b} /* (20, 5, 8) {real, imag} */,
  {32'hbdf22160, 32'h40701611} /* (20, 5, 7) {real, imag} */,
  {32'h40a7d716, 32'h41149441} /* (20, 5, 6) {real, imag} */,
  {32'h40f2fb92, 32'h407e2e88} /* (20, 5, 5) {real, imag} */,
  {32'h3edc4c78, 32'hbfa9e752} /* (20, 5, 4) {real, imag} */,
  {32'hc020b792, 32'hc08fddbe} /* (20, 5, 3) {real, imag} */,
  {32'h3fa50007, 32'hbf239e20} /* (20, 5, 2) {real, imag} */,
  {32'hbf0f5b97, 32'h4072e5bc} /* (20, 5, 1) {real, imag} */,
  {32'hc0c5bdab, 32'h40b79d7f} /* (20, 5, 0) {real, imag} */,
  {32'hbcff6b50, 32'h400d7dcc} /* (20, 4, 31) {real, imag} */,
  {32'hbee3b628, 32'hbff09492} /* (20, 4, 30) {real, imag} */,
  {32'hc0a8c3c0, 32'hc0f0643b} /* (20, 4, 29) {real, imag} */,
  {32'h41152237, 32'hbfc0207c} /* (20, 4, 28) {real, imag} */,
  {32'h411f02d1, 32'h402f7e4a} /* (20, 4, 27) {real, imag} */,
  {32'h3f236782, 32'h3ec2dea8} /* (20, 4, 26) {real, imag} */,
  {32'hc06dbc2a, 32'h40f9f9c7} /* (20, 4, 25) {real, imag} */,
  {32'hc0bfdd6d, 32'h40bff2f7} /* (20, 4, 24) {real, imag} */,
  {32'hbf8431d0, 32'hc0c50d76} /* (20, 4, 23) {real, imag} */,
  {32'h40029510, 32'hbfac5fd2} /* (20, 4, 22) {real, imag} */,
  {32'h405b9df2, 32'h401f480e} /* (20, 4, 21) {real, imag} */,
  {32'hc0bde77d, 32'hc0a65ea3} /* (20, 4, 20) {real, imag} */,
  {32'hc00b518e, 32'hbe8a62ac} /* (20, 4, 19) {real, imag} */,
  {32'h4025724a, 32'h40208ce8} /* (20, 4, 18) {real, imag} */,
  {32'h4087e637, 32'hc10adbe2} /* (20, 4, 17) {real, imag} */,
  {32'h3fb54874, 32'hc117a86c} /* (20, 4, 16) {real, imag} */,
  {32'h3f35e1a4, 32'hc0bb250f} /* (20, 4, 15) {real, imag} */,
  {32'h405cd07e, 32'h4080b933} /* (20, 4, 14) {real, imag} */,
  {32'hc022d9fb, 32'h3fdef9fc} /* (20, 4, 13) {real, imag} */,
  {32'hc0f3b97a, 32'h40af81c5} /* (20, 4, 12) {real, imag} */,
  {32'h3ee9cd70, 32'h407cb508} /* (20, 4, 11) {real, imag} */,
  {32'h40a09120, 32'h3fc85f3b} /* (20, 4, 10) {real, imag} */,
  {32'hbf8d4e5a, 32'h400581be} /* (20, 4, 9) {real, imag} */,
  {32'h3f4b61d4, 32'hc0e75530} /* (20, 4, 8) {real, imag} */,
  {32'h40ea7d52, 32'hc0f8ab48} /* (20, 4, 7) {real, imag} */,
  {32'h4041c32f, 32'hc056a7b1} /* (20, 4, 6) {real, imag} */,
  {32'hbfb407cf, 32'hc01122ce} /* (20, 4, 5) {real, imag} */,
  {32'hbf800471, 32'hc08446ba} /* (20, 4, 4) {real, imag} */,
  {32'h405cb4fd, 32'hc0cf667e} /* (20, 4, 3) {real, imag} */,
  {32'h403c7df8, 32'hc0d36f56} /* (20, 4, 2) {real, imag} */,
  {32'hc0413357, 32'hc0987e5f} /* (20, 4, 1) {real, imag} */,
  {32'hc087032a, 32'hbfee9f35} /* (20, 4, 0) {real, imag} */,
  {32'h405e14cb, 32'hbf6e7679} /* (20, 3, 31) {real, imag} */,
  {32'h3fd8dc29, 32'hc0988b5c} /* (20, 3, 30) {real, imag} */,
  {32'hbf979e32, 32'hc05c1579} /* (20, 3, 29) {real, imag} */,
  {32'hbff4dd1f, 32'hc10019bf} /* (20, 3, 28) {real, imag} */,
  {32'hc122af00, 32'hbfed0752} /* (20, 3, 27) {real, imag} */,
  {32'hc12aeb8c, 32'hc053974a} /* (20, 3, 26) {real, imag} */,
  {32'hc12d3cd4, 32'hc0aca3dc} /* (20, 3, 25) {real, imag} */,
  {32'hbe02d234, 32'hbea70004} /* (20, 3, 24) {real, imag} */,
  {32'hbff7597e, 32'h409ed6ea} /* (20, 3, 23) {real, imag} */,
  {32'hc0c505c4, 32'h40fbed9a} /* (20, 3, 22) {real, imag} */,
  {32'hc05973b7, 32'h41513d0a} /* (20, 3, 21) {real, imag} */,
  {32'hc10f125e, 32'h3fbfed28} /* (20, 3, 20) {real, imag} */,
  {32'hc15fc024, 32'hbf6e94a0} /* (20, 3, 19) {real, imag} */,
  {32'hc0989c39, 32'h40043c99} /* (20, 3, 18) {real, imag} */,
  {32'hc0268ecd, 32'hc0152f71} /* (20, 3, 17) {real, imag} */,
  {32'h40868975, 32'hc0e59e26} /* (20, 3, 16) {real, imag} */,
  {32'h40c620fc, 32'hc0962620} /* (20, 3, 15) {real, imag} */,
  {32'h4133219e, 32'h40f26a2e} /* (20, 3, 14) {real, imag} */,
  {32'h4103baa2, 32'h40945e16} /* (20, 3, 13) {real, imag} */,
  {32'h3fbbee14, 32'h405241c4} /* (20, 3, 12) {real, imag} */,
  {32'h406e6819, 32'h408ec933} /* (20, 3, 11) {real, imag} */,
  {32'h4055fb78, 32'h40aa063c} /* (20, 3, 10) {real, imag} */,
  {32'h40070226, 32'h403e9b6d} /* (20, 3, 9) {real, imag} */,
  {32'h4098ae3d, 32'h3f6852ac} /* (20, 3, 8) {real, imag} */,
  {32'h40c0bd53, 32'hc11691e2} /* (20, 3, 7) {real, imag} */,
  {32'h4086f981, 32'hc13abc54} /* (20, 3, 6) {real, imag} */,
  {32'h40bb13d7, 32'h40102e82} /* (20, 3, 5) {real, imag} */,
  {32'h3f3cfcd0, 32'h3ec7b8b0} /* (20, 3, 4) {real, imag} */,
  {32'h3f600d00, 32'hc0971059} /* (20, 3, 3) {real, imag} */,
  {32'h404dcc5d, 32'h3fdaead5} /* (20, 3, 2) {real, imag} */,
  {32'h414104de, 32'h40e6ddcc} /* (20, 3, 1) {real, imag} */,
  {32'h40a56074, 32'h40a2fe2a} /* (20, 3, 0) {real, imag} */,
  {32'h3fc26014, 32'h3f8fe83f} /* (20, 2, 31) {real, imag} */,
  {32'hc0e937cc, 32'h403e1b01} /* (20, 2, 30) {real, imag} */,
  {32'hc0ee1df1, 32'hc017b7b4} /* (20, 2, 29) {real, imag} */,
  {32'h4004b112, 32'hc085055a} /* (20, 2, 28) {real, imag} */,
  {32'h40a23c3a, 32'h3d8d5a00} /* (20, 2, 27) {real, imag} */,
  {32'h407b1144, 32'h408bde15} /* (20, 2, 26) {real, imag} */,
  {32'h40e98f4f, 32'h4118942d} /* (20, 2, 25) {real, imag} */,
  {32'h415a8d8f, 32'h3fb4a596} /* (20, 2, 24) {real, imag} */,
  {32'h410e8f90, 32'h401e3606} /* (20, 2, 23) {real, imag} */,
  {32'h410771af, 32'h40ceef54} /* (20, 2, 22) {real, imag} */,
  {32'h40e00e8c, 32'h3fc421b8} /* (20, 2, 21) {real, imag} */,
  {32'h4029afd8, 32'h40aab78e} /* (20, 2, 20) {real, imag} */,
  {32'h40e7a966, 32'h409769b0} /* (20, 2, 19) {real, imag} */,
  {32'hc0428e60, 32'h4093f0e4} /* (20, 2, 18) {real, imag} */,
  {32'hc107b8bd, 32'h40e121e0} /* (20, 2, 17) {real, imag} */,
  {32'hc1055aa0, 32'h40aea38e} /* (20, 2, 16) {real, imag} */,
  {32'hc0f2bed0, 32'h40155c8a} /* (20, 2, 15) {real, imag} */,
  {32'h3fb79b60, 32'h402942b4} /* (20, 2, 14) {real, imag} */,
  {32'hbda68630, 32'h405de97f} /* (20, 2, 13) {real, imag} */,
  {32'hc0a6a894, 32'h4085d5ba} /* (20, 2, 12) {real, imag} */,
  {32'h4020f627, 32'h3f646e28} /* (20, 2, 11) {real, imag} */,
  {32'h402f9cf2, 32'hc002105b} /* (20, 2, 10) {real, imag} */,
  {32'hbdc8a088, 32'h4084ec52} /* (20, 2, 9) {real, imag} */,
  {32'hc0ca4bf9, 32'h40f0d64a} /* (20, 2, 8) {real, imag} */,
  {32'hc11ae407, 32'hbf15c0c6} /* (20, 2, 7) {real, imag} */,
  {32'hc0a0815c, 32'hc001182a} /* (20, 2, 6) {real, imag} */,
  {32'h40002aa5, 32'hc0deef63} /* (20, 2, 5) {real, imag} */,
  {32'hc062ff83, 32'hc0aa7178} /* (20, 2, 4) {real, imag} */,
  {32'hc095317e, 32'hc12cd5bd} /* (20, 2, 3) {real, imag} */,
  {32'hc07dc643, 32'hc01d5ecd} /* (20, 2, 2) {real, imag} */,
  {32'h4101cb6e, 32'hbfd5599b} /* (20, 2, 1) {real, imag} */,
  {32'h41233f2c, 32'hc00b39cb} /* (20, 2, 0) {real, imag} */,
  {32'hc092ab85, 32'h4110da72} /* (20, 1, 31) {real, imag} */,
  {32'hc0c5e65c, 32'h40d5df88} /* (20, 1, 30) {real, imag} */,
  {32'h408e7621, 32'hbff5a22e} /* (20, 1, 29) {real, imag} */,
  {32'h3f557d82, 32'hbf571132} /* (20, 1, 28) {real, imag} */,
  {32'hc022e214, 32'hc084c028} /* (20, 1, 27) {real, imag} */,
  {32'hbfbafd42, 32'h3fbd2646} /* (20, 1, 26) {real, imag} */,
  {32'h408144b2, 32'h40c68d80} /* (20, 1, 25) {real, imag} */,
  {32'hbf0d66b7, 32'h411856e5} /* (20, 1, 24) {real, imag} */,
  {32'h40061155, 32'hc0debfdb} /* (20, 1, 23) {real, imag} */,
  {32'h3fe31712, 32'hc10751e6} /* (20, 1, 22) {real, imag} */,
  {32'h4029270d, 32'hc000289f} /* (20, 1, 21) {real, imag} */,
  {32'h4112104f, 32'hc03ea1bd} /* (20, 1, 20) {real, imag} */,
  {32'h40d92cf6, 32'h40a8ac6b} /* (20, 1, 19) {real, imag} */,
  {32'h3f4fb210, 32'h3f6067a0} /* (20, 1, 18) {real, imag} */,
  {32'hc047c0ad, 32'hc10d67c0} /* (20, 1, 17) {real, imag} */,
  {32'hc01a959a, 32'h40b6c33c} /* (20, 1, 16) {real, imag} */,
  {32'h4034cc08, 32'h3f64712e} /* (20, 1, 15) {real, imag} */,
  {32'h415ded20, 32'hc0af3096} /* (20, 1, 14) {real, imag} */,
  {32'h4023a26a, 32'hc0c8b0b1} /* (20, 1, 13) {real, imag} */,
  {32'h400e859a, 32'hbfc9a684} /* (20, 1, 12) {real, imag} */,
  {32'h40422216, 32'h3f075bb8} /* (20, 1, 11) {real, imag} */,
  {32'h40839647, 32'h40d23b8a} /* (20, 1, 10) {real, imag} */,
  {32'h40a2b63c, 32'h4057abf6} /* (20, 1, 9) {real, imag} */,
  {32'h41088e7e, 32'hc09110da} /* (20, 1, 8) {real, imag} */,
  {32'h40c7d515, 32'h3f977d25} /* (20, 1, 7) {real, imag} */,
  {32'h4047ded6, 32'h3fbd83ae} /* (20, 1, 6) {real, imag} */,
  {32'h40875ac6, 32'hc128a09b} /* (20, 1, 5) {real, imag} */,
  {32'hc092a774, 32'hc120b21c} /* (20, 1, 4) {real, imag} */,
  {32'hc05dce3a, 32'hc02237fe} /* (20, 1, 3) {real, imag} */,
  {32'hc090b6d5, 32'hc09f2a6f} /* (20, 1, 2) {real, imag} */,
  {32'hc1025684, 32'hc0d96cbb} /* (20, 1, 1) {real, imag} */,
  {32'hc02695cc, 32'hc0d885e9} /* (20, 1, 0) {real, imag} */,
  {32'hc052f0f7, 32'h3f1e0acc} /* (20, 0, 31) {real, imag} */,
  {32'hc07cd8ea, 32'hc0333e1c} /* (20, 0, 30) {real, imag} */,
  {32'hbfc99eb8, 32'h3f10d7fc} /* (20, 0, 29) {real, imag} */,
  {32'hbfe991c6, 32'hbf07f09f} /* (20, 0, 28) {real, imag} */,
  {32'hbf7611d0, 32'h40b34cf6} /* (20, 0, 27) {real, imag} */,
  {32'h40be7620, 32'h40fc79c2} /* (20, 0, 26) {real, imag} */,
  {32'h412270b2, 32'h41318425} /* (20, 0, 25) {real, imag} */,
  {32'hbeff4368, 32'h3ff331ba} /* (20, 0, 24) {real, imag} */,
  {32'hc0efe8e6, 32'hc0b7a37e} /* (20, 0, 23) {real, imag} */,
  {32'hc10c558e, 32'h402dd470} /* (20, 0, 22) {real, imag} */,
  {32'hc0597b22, 32'h409f6f2f} /* (20, 0, 21) {real, imag} */,
  {32'hc09e070d, 32'h410f1b37} /* (20, 0, 20) {real, imag} */,
  {32'hc02cd8a8, 32'hc02d6636} /* (20, 0, 19) {real, imag} */,
  {32'hc1158562, 32'hc12836c9} /* (20, 0, 18) {real, imag} */,
  {32'hbfd75a3e, 32'hc09f170d} /* (20, 0, 17) {real, imag} */,
  {32'h40cc8094, 32'hc0a5b694} /* (20, 0, 16) {real, imag} */,
  {32'h3e5e0304, 32'h3f478a33} /* (20, 0, 15) {real, imag} */,
  {32'hc0da3c9a, 32'h41401628} /* (20, 0, 14) {real, imag} */,
  {32'hc11448e6, 32'h4111a106} /* (20, 0, 13) {real, imag} */,
  {32'h408304b6, 32'hc0598d2c} /* (20, 0, 12) {real, imag} */,
  {32'h40cc94d8, 32'hc09446fb} /* (20, 0, 11) {real, imag} */,
  {32'h410b4818, 32'h3f8b01fc} /* (20, 0, 10) {real, imag} */,
  {32'h402cd3bc, 32'hbfc81365} /* (20, 0, 9) {real, imag} */,
  {32'hbf4eb694, 32'h4047449c} /* (20, 0, 8) {real, imag} */,
  {32'h3f153224, 32'h40169a12} /* (20, 0, 7) {real, imag} */,
  {32'hc003b114, 32'h40c44d70} /* (20, 0, 6) {real, imag} */,
  {32'h40c867de, 32'hbead9f4e} /* (20, 0, 5) {real, imag} */,
  {32'h40efd17c, 32'hc0b188fc} /* (20, 0, 4) {real, imag} */,
  {32'hc135e443, 32'h40c4a3e8} /* (20, 0, 3) {real, imag} */,
  {32'hc17bed05, 32'h40964c08} /* (20, 0, 2) {real, imag} */,
  {32'hbf03ff18, 32'h3f8f674f} /* (20, 0, 1) {real, imag} */,
  {32'h4088863e, 32'h40cd5520} /* (20, 0, 0) {real, imag} */,
  {32'hc01be229, 32'hc13175cc} /* (19, 31, 31) {real, imag} */,
  {32'h404c6ecc, 32'hc107e90e} /* (19, 31, 30) {real, imag} */,
  {32'h40a841a0, 32'hc00019c4} /* (19, 31, 29) {real, imag} */,
  {32'hbf22d7f0, 32'hc09197d2} /* (19, 31, 28) {real, imag} */,
  {32'hc0cd3e78, 32'hc1496d94} /* (19, 31, 27) {real, imag} */,
  {32'h3e5e32f8, 32'hbff6e870} /* (19, 31, 26) {real, imag} */,
  {32'hbee74316, 32'h3fc14b0e} /* (19, 31, 25) {real, imag} */,
  {32'hc0a58f8f, 32'hc0357e64} /* (19, 31, 24) {real, imag} */,
  {32'h4088af49, 32'hbf9fe4a6} /* (19, 31, 23) {real, imag} */,
  {32'h410e24e6, 32'h401dc003} /* (19, 31, 22) {real, imag} */,
  {32'h407bba69, 32'hbf092a46} /* (19, 31, 21) {real, imag} */,
  {32'h4071fffc, 32'hc003ae3c} /* (19, 31, 20) {real, imag} */,
  {32'hc05657d6, 32'hc0d3d89a} /* (19, 31, 19) {real, imag} */,
  {32'hc0ca3583, 32'hc0414d6c} /* (19, 31, 18) {real, imag} */,
  {32'hc0a6ab6a, 32'hc0a3f3b9} /* (19, 31, 17) {real, imag} */,
  {32'h40290b52, 32'hc08738b9} /* (19, 31, 16) {real, imag} */,
  {32'h40ef1e63, 32'hc0444953} /* (19, 31, 15) {real, imag} */,
  {32'h4044b583, 32'h407eacd3} /* (19, 31, 14) {real, imag} */,
  {32'hc00bc7a8, 32'hc015a02e} /* (19, 31, 13) {real, imag} */,
  {32'h41407ae8, 32'hbe018200} /* (19, 31, 12) {real, imag} */,
  {32'h40607dfe, 32'h40e4ab08} /* (19, 31, 11) {real, imag} */,
  {32'h406960bc, 32'h411e8afa} /* (19, 31, 10) {real, imag} */,
  {32'h409b8e8b, 32'h3fc9442a} /* (19, 31, 9) {real, imag} */,
  {32'h3fc6fc2e, 32'h40a5e512} /* (19, 31, 8) {real, imag} */,
  {32'hc0622614, 32'hbf7a203c} /* (19, 31, 7) {real, imag} */,
  {32'hc02e05cc, 32'h3ff54bee} /* (19, 31, 6) {real, imag} */,
  {32'hbea406f0, 32'h4100d95f} /* (19, 31, 5) {real, imag} */,
  {32'h3f1bf438, 32'h40c69029} /* (19, 31, 4) {real, imag} */,
  {32'hc01c4d04, 32'h405787ac} /* (19, 31, 3) {real, imag} */,
  {32'h3f40a3b4, 32'h410de295} /* (19, 31, 2) {real, imag} */,
  {32'h4135dfed, 32'hbfce56e6} /* (19, 31, 1) {real, imag} */,
  {32'h40eabaf4, 32'hc0d922be} /* (19, 31, 0) {real, imag} */,
  {32'h40b4e396, 32'hc0b3f0b5} /* (19, 30, 31) {real, imag} */,
  {32'h413a69e0, 32'hc1231a28} /* (19, 30, 30) {real, imag} */,
  {32'hc04fe020, 32'hc0b88d6f} /* (19, 30, 29) {real, imag} */,
  {32'hc076fe08, 32'h3fc3aa30} /* (19, 30, 28) {real, imag} */,
  {32'hc0c1d19d, 32'h409acc92} /* (19, 30, 27) {real, imag} */,
  {32'hc10acb18, 32'h40aca317} /* (19, 30, 26) {real, imag} */,
  {32'hc0bda7fe, 32'h409b4d48} /* (19, 30, 25) {real, imag} */,
  {32'hc0cf9401, 32'h405b3d24} /* (19, 30, 24) {real, imag} */,
  {32'h4096f9dd, 32'h408eeec0} /* (19, 30, 23) {real, imag} */,
  {32'h40f010b1, 32'h411210d1} /* (19, 30, 22) {real, imag} */,
  {32'hbf3fecec, 32'h40503dc6} /* (19, 30, 21) {real, imag} */,
  {32'hbfe8c60c, 32'h3fc3c128} /* (19, 30, 20) {real, imag} */,
  {32'h3fe31c44, 32'h40c5c05a} /* (19, 30, 19) {real, imag} */,
  {32'h3f94e8f4, 32'hc0c16f09} /* (19, 30, 18) {real, imag} */,
  {32'hc0d16700, 32'hc0cf2d7b} /* (19, 30, 17) {real, imag} */,
  {32'hbf801905, 32'hc122f89a} /* (19, 30, 16) {real, imag} */,
  {32'h411a5e4a, 32'hc12b6075} /* (19, 30, 15) {real, imag} */,
  {32'h41168cbb, 32'hc137fb03} /* (19, 30, 14) {real, imag} */,
  {32'hc0000e4f, 32'hc0abcea2} /* (19, 30, 13) {real, imag} */,
  {32'hc059ac6b, 32'h3f7b1b88} /* (19, 30, 12) {real, imag} */,
  {32'h40d58512, 32'h4059f374} /* (19, 30, 11) {real, imag} */,
  {32'h40f06eed, 32'h3fa9c55d} /* (19, 30, 10) {real, imag} */,
  {32'h4134af3e, 32'hc0ba1847} /* (19, 30, 9) {real, imag} */,
  {32'h4122f18b, 32'hc092b353} /* (19, 30, 8) {real, imag} */,
  {32'h40ade14f, 32'hc0d59ec8} /* (19, 30, 7) {real, imag} */,
  {32'h3f3b1a9c, 32'h40ba818c} /* (19, 30, 6) {real, imag} */,
  {32'hc006031c, 32'h41389d5b} /* (19, 30, 5) {real, imag} */,
  {32'h3fb2d234, 32'h40634036} /* (19, 30, 4) {real, imag} */,
  {32'h409b6894, 32'hc068fa95} /* (19, 30, 3) {real, imag} */,
  {32'h412e270e, 32'h3f83ff26} /* (19, 30, 2) {real, imag} */,
  {32'h40d4fb83, 32'h4096875a} /* (19, 30, 1) {real, imag} */,
  {32'h3edc2f37, 32'h3f2a1f9e} /* (19, 30, 0) {real, imag} */,
  {32'h401f9b21, 32'h3fcb1675} /* (19, 29, 31) {real, imag} */,
  {32'hc0374076, 32'h40878e6d} /* (19, 29, 30) {real, imag} */,
  {32'hc02dbfaa, 32'h4039efb3} /* (19, 29, 29) {real, imag} */,
  {32'h4010af1b, 32'hbf605e1a} /* (19, 29, 28) {real, imag} */,
  {32'hc012fc80, 32'hc0e68b60} /* (19, 29, 27) {real, imag} */,
  {32'hc0594626, 32'hbfe65388} /* (19, 29, 26) {real, imag} */,
  {32'hbffb61e8, 32'hc02133b4} /* (19, 29, 25) {real, imag} */,
  {32'hbf4320db, 32'hbc767400} /* (19, 29, 24) {real, imag} */,
  {32'h3f8b8d9a, 32'h3fea5028} /* (19, 29, 23) {real, imag} */,
  {32'h40592a60, 32'hbf844648} /* (19, 29, 22) {real, imag} */,
  {32'hc0e401f9, 32'h40774a40} /* (19, 29, 21) {real, imag} */,
  {32'hc139b15b, 32'hbf42ef9c} /* (19, 29, 20) {real, imag} */,
  {32'h3cb9a2c0, 32'h3f9002a8} /* (19, 29, 19) {real, imag} */,
  {32'h4024b9f0, 32'h3e941a6f} /* (19, 29, 18) {real, imag} */,
  {32'h3f280246, 32'hc07ca951} /* (19, 29, 17) {real, imag} */,
  {32'hc00c48dd, 32'hc08da86e} /* (19, 29, 16) {real, imag} */,
  {32'h3fb65db6, 32'hbfcb7a93} /* (19, 29, 15) {real, imag} */,
  {32'hbfe15b62, 32'h4042ca6a} /* (19, 29, 14) {real, imag} */,
  {32'hc014793d, 32'h400b76b8} /* (19, 29, 13) {real, imag} */,
  {32'h3db13540, 32'h3ece0308} /* (19, 29, 12) {real, imag} */,
  {32'h3e0cc5d8, 32'hbee05a78} /* (19, 29, 11) {real, imag} */,
  {32'h3ff46cc9, 32'h405d316f} /* (19, 29, 10) {real, imag} */,
  {32'h3fd1dda4, 32'hbef1ccae} /* (19, 29, 9) {real, imag} */,
  {32'h40a3b69d, 32'hc016deed} /* (19, 29, 8) {real, imag} */,
  {32'h40d6ca71, 32'h3fa9b902} /* (19, 29, 7) {real, imag} */,
  {32'h40158c0a, 32'h3f899639} /* (19, 29, 6) {real, imag} */,
  {32'hc001e70a, 32'hc0ba2dc9} /* (19, 29, 5) {real, imag} */,
  {32'hc0b271e5, 32'hbfee7949} /* (19, 29, 4) {real, imag} */,
  {32'hc081140f, 32'h403aa742} /* (19, 29, 3) {real, imag} */,
  {32'hc1142aae, 32'h40b61564} /* (19, 29, 2) {real, imag} */,
  {32'hc10aad8c, 32'h40395883} /* (19, 29, 1) {real, imag} */,
  {32'hc0a3835c, 32'hc05cdc54} /* (19, 29, 0) {real, imag} */,
  {32'h405dbf14, 32'hbffd1dca} /* (19, 28, 31) {real, imag} */,
  {32'h404652c0, 32'hc0872bae} /* (19, 28, 30) {real, imag} */,
  {32'h40e03450, 32'h3fd618f9} /* (19, 28, 29) {real, imag} */,
  {32'h408eec4f, 32'h4084eb37} /* (19, 28, 28) {real, imag} */,
  {32'h3b53c400, 32'h4109af76} /* (19, 28, 27) {real, imag} */,
  {32'hc10153f6, 32'h4100db28} /* (19, 28, 26) {real, imag} */,
  {32'hc017f5d4, 32'h40f84b2c} /* (19, 28, 25) {real, imag} */,
  {32'h408cbc0c, 32'h40bd5866} /* (19, 28, 24) {real, imag} */,
  {32'h409ea6f2, 32'hbf963fac} /* (19, 28, 23) {real, imag} */,
  {32'h4132eac6, 32'hc0ef1414} /* (19, 28, 22) {real, imag} */,
  {32'h40e2e41c, 32'hbfa378e4} /* (19, 28, 21) {real, imag} */,
  {32'h40609bd7, 32'h3fa03376} /* (19, 28, 20) {real, imag} */,
  {32'hc03c13f2, 32'h4038ae23} /* (19, 28, 19) {real, imag} */,
  {32'h3f80a3ce, 32'h40888f5c} /* (19, 28, 18) {real, imag} */,
  {32'hbdfb38b0, 32'hbdb896a0} /* (19, 28, 17) {real, imag} */,
  {32'hc01d5a41, 32'hc01c3213} /* (19, 28, 16) {real, imag} */,
  {32'hbe52b070, 32'hc0986a89} /* (19, 28, 15) {real, imag} */,
  {32'h3f0167f8, 32'h400f1137} /* (19, 28, 14) {real, imag} */,
  {32'hbf1bd0b8, 32'h40b6c055} /* (19, 28, 13) {real, imag} */,
  {32'hbfe1bdd0, 32'h40f4cf81} /* (19, 28, 12) {real, imag} */,
  {32'hc10052c3, 32'h40d79374} /* (19, 28, 11) {real, imag} */,
  {32'hc0d2d28b, 32'h3fcba991} /* (19, 28, 10) {real, imag} */,
  {32'hbff4b712, 32'h3ea8a3fc} /* (19, 28, 9) {real, imag} */,
  {32'hc0346cc0, 32'h4005faed} /* (19, 28, 8) {real, imag} */,
  {32'h3fd1302d, 32'h3f9c35b6} /* (19, 28, 7) {real, imag} */,
  {32'h406c767c, 32'hbf88f4f5} /* (19, 28, 6) {real, imag} */,
  {32'h400bdf4c, 32'h4085defc} /* (19, 28, 5) {real, imag} */,
  {32'h3fc4c4c7, 32'h40aaf06e} /* (19, 28, 4) {real, imag} */,
  {32'hc01156b0, 32'h3d582e80} /* (19, 28, 3) {real, imag} */,
  {32'hbfb1cb33, 32'hc00bfba4} /* (19, 28, 2) {real, imag} */,
  {32'hbfb70b8e, 32'h3e283e8c} /* (19, 28, 1) {real, imag} */,
  {32'h404ad8c0, 32'h4023338a} /* (19, 28, 0) {real, imag} */,
  {32'h409fb883, 32'h40c17b23} /* (19, 27, 31) {real, imag} */,
  {32'h411584be, 32'h4032856f} /* (19, 27, 30) {real, imag} */,
  {32'h40217e93, 32'h405f6dd0} /* (19, 27, 29) {real, imag} */,
  {32'h40e04016, 32'hc02f5f76} /* (19, 27, 28) {real, imag} */,
  {32'h40baabd6, 32'hbed54850} /* (19, 27, 27) {real, imag} */,
  {32'h3fc8cd3c, 32'hc09c47ba} /* (19, 27, 26) {real, imag} */,
  {32'h40b606e1, 32'hc086b69a} /* (19, 27, 25) {real, imag} */,
  {32'h3f806512, 32'hc0425cdd} /* (19, 27, 24) {real, imag} */,
  {32'hc0c596ba, 32'hbf80f51f} /* (19, 27, 23) {real, imag} */,
  {32'h404e7d77, 32'h3f9ec1e6} /* (19, 27, 22) {real, imag} */,
  {32'h411ad1ed, 32'hc004d640} /* (19, 27, 21) {real, imag} */,
  {32'h4050fe77, 32'h40930240} /* (19, 27, 20) {real, imag} */,
  {32'hbfe694ea, 32'h4146230e} /* (19, 27, 19) {real, imag} */,
  {32'h3cbed600, 32'h3fb1984b} /* (19, 27, 18) {real, imag} */,
  {32'h3fe5f66e, 32'hc108851a} /* (19, 27, 17) {real, imag} */,
  {32'h4121b152, 32'hbfba5d4a} /* (19, 27, 16) {real, imag} */,
  {32'h401a1ded, 32'h4031c258} /* (19, 27, 15) {real, imag} */,
  {32'hc0922215, 32'h3f675d00} /* (19, 27, 14) {real, imag} */,
  {32'hbfca0398, 32'hc07561f5} /* (19, 27, 13) {real, imag} */,
  {32'h40e6cb05, 32'hc067c836} /* (19, 27, 12) {real, imag} */,
  {32'h41028124, 32'h3f4056ec} /* (19, 27, 11) {real, imag} */,
  {32'h40bc6e45, 32'h40ab43aa} /* (19, 27, 10) {real, imag} */,
  {32'hbf122048, 32'h40c6d2ac} /* (19, 27, 9) {real, imag} */,
  {32'hc06af1d2, 32'h4000cc2e} /* (19, 27, 8) {real, imag} */,
  {32'hc04a01b0, 32'h3f4c80cc} /* (19, 27, 7) {real, imag} */,
  {32'hc075404c, 32'h405b1a46} /* (19, 27, 6) {real, imag} */,
  {32'hc08b0848, 32'h4078858a} /* (19, 27, 5) {real, imag} */,
  {32'hc0bf5e9b, 32'h402de83a} /* (19, 27, 4) {real, imag} */,
  {32'hc12c2e8f, 32'h3eb75786} /* (19, 27, 3) {real, imag} */,
  {32'h40142189, 32'hc0a1046c} /* (19, 27, 2) {real, imag} */,
  {32'h40d26819, 32'hc0e7c435} /* (19, 27, 1) {real, imag} */,
  {32'hbf8d839f, 32'h3fcf59de} /* (19, 27, 0) {real, imag} */,
  {32'h403cb38f, 32'h3f111294} /* (19, 26, 31) {real, imag} */,
  {32'h3fe89531, 32'hbe755278} /* (19, 26, 30) {real, imag} */,
  {32'hc0cee81c, 32'h3f8ef344} /* (19, 26, 29) {real, imag} */,
  {32'hc1006d52, 32'h4049ae8f} /* (19, 26, 28) {real, imag} */,
  {32'hbf193c7a, 32'hbfe2f922} /* (19, 26, 27) {real, imag} */,
  {32'h3fe7ebf2, 32'h4011a89b} /* (19, 26, 26) {real, imag} */,
  {32'h40677de8, 32'h40fe6b04} /* (19, 26, 25) {real, imag} */,
  {32'hc08ca1c7, 32'h40abb74b} /* (19, 26, 24) {real, imag} */,
  {32'hc0b26e7e, 32'hc02dacaa} /* (19, 26, 23) {real, imag} */,
  {32'hbfcbdcbf, 32'hc0b732f3} /* (19, 26, 22) {real, imag} */,
  {32'h3d22ac40, 32'h3fc23408} /* (19, 26, 21) {real, imag} */,
  {32'h4104e626, 32'hbeda0570} /* (19, 26, 20) {real, imag} */,
  {32'h40ef05d4, 32'hbf7f57e9} /* (19, 26, 19) {real, imag} */,
  {32'h41227638, 32'hc0af606a} /* (19, 26, 18) {real, imag} */,
  {32'h3f3f5268, 32'hc0cef489} /* (19, 26, 17) {real, imag} */,
  {32'hbfebbf00, 32'h3fb06ed8} /* (19, 26, 16) {real, imag} */,
  {32'h3fd7bff3, 32'hbf37c02f} /* (19, 26, 15) {real, imag} */,
  {32'h40a29e5f, 32'hc03b5ec8} /* (19, 26, 14) {real, imag} */,
  {32'hbfdb6121, 32'h4067e0f5} /* (19, 26, 13) {real, imag} */,
  {32'hc09724b4, 32'h408c3304} /* (19, 26, 12) {real, imag} */,
  {32'h409ebe62, 32'h40bd47cb} /* (19, 26, 11) {real, imag} */,
  {32'h404e94b6, 32'hbfa35f6c} /* (19, 26, 10) {real, imag} */,
  {32'hc0880e09, 32'hc07f370e} /* (19, 26, 9) {real, imag} */,
  {32'hc0472dfe, 32'hc0454766} /* (19, 26, 8) {real, imag} */,
  {32'h406971ae, 32'hc02de260} /* (19, 26, 7) {real, imag} */,
  {32'h3f093b74, 32'hc0f247dc} /* (19, 26, 6) {real, imag} */,
  {32'h408dacb2, 32'hc0edc19c} /* (19, 26, 5) {real, imag} */,
  {32'h407a52ca, 32'h4013f13e} /* (19, 26, 4) {real, imag} */,
  {32'h40dd623c, 32'hbfe46cfe} /* (19, 26, 3) {real, imag} */,
  {32'hbea03918, 32'hc0df872e} /* (19, 26, 2) {real, imag} */,
  {32'hc06af761, 32'hc0491580} /* (19, 26, 1) {real, imag} */,
  {32'hbf37ff12, 32'h3fc3fd4d} /* (19, 26, 0) {real, imag} */,
  {32'h3e044ab0, 32'h4045f124} /* (19, 25, 31) {real, imag} */,
  {32'h3ffc63a8, 32'h3f52dc56} /* (19, 25, 30) {real, imag} */,
  {32'h3fde5a7a, 32'hc02b20fb} /* (19, 25, 29) {real, imag} */,
  {32'h406e96de, 32'hc05b0877} /* (19, 25, 28) {real, imag} */,
  {32'hbe8ec5a4, 32'h4027e0b6} /* (19, 25, 27) {real, imag} */,
  {32'hbeede4cc, 32'h3f38ad78} /* (19, 25, 26) {real, imag} */,
  {32'h40766ad0, 32'hc039a70a} /* (19, 25, 25) {real, imag} */,
  {32'h41018eda, 32'h3fa3beb4} /* (19, 25, 24) {real, imag} */,
  {32'h3f28d0e0, 32'h40aed4ae} /* (19, 25, 23) {real, imag} */,
  {32'hc0b598ee, 32'h3ffd018d} /* (19, 25, 22) {real, imag} */,
  {32'hbff1adee, 32'h404b717a} /* (19, 25, 21) {real, imag} */,
  {32'hc0923120, 32'hbf7191b4} /* (19, 25, 20) {real, imag} */,
  {32'hc0be8d91, 32'hbe4c3b38} /* (19, 25, 19) {real, imag} */,
  {32'hc050f5b3, 32'h4079b652} /* (19, 25, 18) {real, imag} */,
  {32'hc0b4a921, 32'h4086f7b9} /* (19, 25, 17) {real, imag} */,
  {32'hc02ad956, 32'h4009f039} /* (19, 25, 16) {real, imag} */,
  {32'hc04f69f8, 32'hbfe930e1} /* (19, 25, 15) {real, imag} */,
  {32'hc0827704, 32'hc024fe8f} /* (19, 25, 14) {real, imag} */,
  {32'hc0be3fdd, 32'hbf07848c} /* (19, 25, 13) {real, imag} */,
  {32'hc099a06c, 32'hbe4be400} /* (19, 25, 12) {real, imag} */,
  {32'hc082387b, 32'hc0a3dc73} /* (19, 25, 11) {real, imag} */,
  {32'h40909804, 32'hbfb6d4fa} /* (19, 25, 10) {real, imag} */,
  {32'h408918b2, 32'h40768bbc} /* (19, 25, 9) {real, imag} */,
  {32'hc0d51644, 32'hbeb6a2a0} /* (19, 25, 8) {real, imag} */,
  {32'hc092276a, 32'h3ef073b4} /* (19, 25, 7) {real, imag} */,
  {32'h40832ab2, 32'hc03cee67} /* (19, 25, 6) {real, imag} */,
  {32'h3f9a39e6, 32'h402601d3} /* (19, 25, 5) {real, imag} */,
  {32'hbf68f2e5, 32'h40cb6749} /* (19, 25, 4) {real, imag} */,
  {32'hc05b5a5c, 32'h3fb21c0b} /* (19, 25, 3) {real, imag} */,
  {32'hc08e4c91, 32'hbf4bdaa0} /* (19, 25, 2) {real, imag} */,
  {32'hc0980bfd, 32'hbf64ecd4} /* (19, 25, 1) {real, imag} */,
  {32'hbfd95b3a, 32'h3fb03952} /* (19, 25, 0) {real, imag} */,
  {32'h408ef092, 32'hc01ce60b} /* (19, 24, 31) {real, imag} */,
  {32'h408af17d, 32'hc0b2812e} /* (19, 24, 30) {real, imag} */,
  {32'h405704da, 32'hbed2e718} /* (19, 24, 29) {real, imag} */,
  {32'h3ea7fb6c, 32'h4082bd14} /* (19, 24, 28) {real, imag} */,
  {32'hbf03750c, 32'h3c0f7f80} /* (19, 24, 27) {real, imag} */,
  {32'hbf93646c, 32'h3fe2fd02} /* (19, 24, 26) {real, imag} */,
  {32'hbf2bf1a3, 32'h3fcf8543} /* (19, 24, 25) {real, imag} */,
  {32'h409cd3ea, 32'hc005168a} /* (19, 24, 24) {real, imag} */,
  {32'h404cefcd, 32'h4038249d} /* (19, 24, 23) {real, imag} */,
  {32'h401d79fc, 32'h401e9bea} /* (19, 24, 22) {real, imag} */,
  {32'h40af6eff, 32'hbf9b7116} /* (19, 24, 21) {real, imag} */,
  {32'h40251960, 32'hc0862aea} /* (19, 24, 20) {real, imag} */,
  {32'h3f9aea4e, 32'hc0bd8cc0} /* (19, 24, 19) {real, imag} */,
  {32'hc062fe24, 32'hc08c4d3d} /* (19, 24, 18) {real, imag} */,
  {32'h40184590, 32'h3f22c7f0} /* (19, 24, 17) {real, imag} */,
  {32'h406ae96d, 32'h3fa3f174} /* (19, 24, 16) {real, imag} */,
  {32'hc06e7821, 32'h401eb814} /* (19, 24, 15) {real, imag} */,
  {32'hc01548d6, 32'h4001b851} /* (19, 24, 14) {real, imag} */,
  {32'hbf92f687, 32'h4014fd41} /* (19, 24, 13) {real, imag} */,
  {32'hc09646cb, 32'h4101371b} /* (19, 24, 12) {real, imag} */,
  {32'hc08cc2ec, 32'h40a032a8} /* (19, 24, 11) {real, imag} */,
  {32'h404b8736, 32'h3f8a8ca1} /* (19, 24, 10) {real, imag} */,
  {32'h3fbc83b8, 32'hbd04ff60} /* (19, 24, 9) {real, imag} */,
  {32'h3f02a258, 32'hbfa5ac16} /* (19, 24, 8) {real, imag} */,
  {32'h41039f56, 32'hbff2be95} /* (19, 24, 7) {real, imag} */,
  {32'h4106b79e, 32'hc04e9870} /* (19, 24, 6) {real, imag} */,
  {32'h402b58f0, 32'hc007c2de} /* (19, 24, 5) {real, imag} */,
  {32'h40629588, 32'h3f842496} /* (19, 24, 4) {real, imag} */,
  {32'hbf8d48b5, 32'h40782e61} /* (19, 24, 3) {real, imag} */,
  {32'hbffb234c, 32'h40b9a542} /* (19, 24, 2) {real, imag} */,
  {32'h3f4489b0, 32'h40ae4d80} /* (19, 24, 1) {real, imag} */,
  {32'h3fc1bb46, 32'h404f3160} /* (19, 24, 0) {real, imag} */,
  {32'hc048b39c, 32'hbfc7ff70} /* (19, 23, 31) {real, imag} */,
  {32'hc076a9bc, 32'h3fbe0cbf} /* (19, 23, 30) {real, imag} */,
  {32'h3ea39808, 32'h409c94d9} /* (19, 23, 29) {real, imag} */,
  {32'h3ff922e4, 32'h40134364} /* (19, 23, 28) {real, imag} */,
  {32'h3f83c6eb, 32'h40a1da2f} /* (19, 23, 27) {real, imag} */,
  {32'h405594ef, 32'hbfbdd76a} /* (19, 23, 26) {real, imag} */,
  {32'h401e3a80, 32'hbfe50529} /* (19, 23, 25) {real, imag} */,
  {32'h40f7693a, 32'h409f0ee6} /* (19, 23, 24) {real, imag} */,
  {32'h409bb314, 32'h3fe792b2} /* (19, 23, 23) {real, imag} */,
  {32'hc017aa9f, 32'h3dc6b1f0} /* (19, 23, 22) {real, imag} */,
  {32'hbfd3639d, 32'h4029ef7d} /* (19, 23, 21) {real, imag} */,
  {32'hbfeed586, 32'h3e822496} /* (19, 23, 20) {real, imag} */,
  {32'hc084eaac, 32'hbfd8fb63} /* (19, 23, 19) {real, imag} */,
  {32'hbfe54b5b, 32'hbf125383} /* (19, 23, 18) {real, imag} */,
  {32'hbf21f53f, 32'hc00336a5} /* (19, 23, 17) {real, imag} */,
  {32'hc05b56f0, 32'h3fb5cc7e} /* (19, 23, 16) {real, imag} */,
  {32'hbc868e80, 32'h3f4e33d5} /* (19, 23, 15) {real, imag} */,
  {32'h3f2f4895, 32'h400d0685} /* (19, 23, 14) {real, imag} */,
  {32'h3dd0e9c0, 32'hc0836b8c} /* (19, 23, 13) {real, imag} */,
  {32'h3eb7fa14, 32'hc106fa88} /* (19, 23, 12) {real, imag} */,
  {32'h3e8551de, 32'hc0d06c08} /* (19, 23, 11) {real, imag} */,
  {32'hc0285c68, 32'hc0bce514} /* (19, 23, 10) {real, imag} */,
  {32'hc0be3506, 32'hc0b77f6f} /* (19, 23, 9) {real, imag} */,
  {32'hbebba250, 32'hbd81b000} /* (19, 23, 8) {real, imag} */,
  {32'hbfb1e55a, 32'hbfcd4d8e} /* (19, 23, 7) {real, imag} */,
  {32'hc0bceef4, 32'hc05fe4f5} /* (19, 23, 6) {real, imag} */,
  {32'hc0d0ed62, 32'hbf960484} /* (19, 23, 5) {real, imag} */,
  {32'h401e1b6d, 32'h409bd680} /* (19, 23, 4) {real, imag} */,
  {32'h4104f9bc, 32'h40d932f5} /* (19, 23, 3) {real, imag} */,
  {32'h3f79974c, 32'h3f9f9e24} /* (19, 23, 2) {real, imag} */,
  {32'hc0a127b0, 32'h3ed2a50c} /* (19, 23, 1) {real, imag} */,
  {32'hc07deb46, 32'h3f712ae1} /* (19, 23, 0) {real, imag} */,
  {32'hbedbaed8, 32'hbcbbb180} /* (19, 22, 31) {real, imag} */,
  {32'h3d9a3680, 32'h3ffb5839} /* (19, 22, 30) {real, imag} */,
  {32'hbfab9625, 32'h40427adb} /* (19, 22, 29) {real, imag} */,
  {32'h3fcccc09, 32'h4042edfa} /* (19, 22, 28) {real, imag} */,
  {32'h40903efe, 32'hc001a03d} /* (19, 22, 27) {real, imag} */,
  {32'h3f5fa582, 32'hc0678bf5} /* (19, 22, 26) {real, imag} */,
  {32'h3f5b5dd8, 32'h3f7774b2} /* (19, 22, 25) {real, imag} */,
  {32'h400f1ae8, 32'h3f738d1a} /* (19, 22, 24) {real, imag} */,
  {32'hbfa22996, 32'h3fb2563c} /* (19, 22, 23) {real, imag} */,
  {32'hc05c6cf2, 32'h40a9096a} /* (19, 22, 22) {real, imag} */,
  {32'hc0621986, 32'hbf4233f8} /* (19, 22, 21) {real, imag} */,
  {32'h400905be, 32'hbf94d721} /* (19, 22, 20) {real, imag} */,
  {32'h408e2f7c, 32'h3fbdb926} /* (19, 22, 19) {real, imag} */,
  {32'h3f4c794e, 32'hbfb8630c} /* (19, 22, 18) {real, imag} */,
  {32'hc0595d1e, 32'h3f432370} /* (19, 22, 17) {real, imag} */,
  {32'hc0cb602a, 32'h4004235e} /* (19, 22, 16) {real, imag} */,
  {32'hbfd3fe9d, 32'h409f4c32} /* (19, 22, 15) {real, imag} */,
  {32'hbecaadf8, 32'h404d20c7} /* (19, 22, 14) {real, imag} */,
  {32'hbdad98d0, 32'h3e213990} /* (19, 22, 13) {real, imag} */,
  {32'h40eb8146, 32'hbfa26fac} /* (19, 22, 12) {real, imag} */,
  {32'h4043f0fc, 32'hbff92a0d} /* (19, 22, 11) {real, imag} */,
  {32'h40674194, 32'h4006f054} /* (19, 22, 10) {real, imag} */,
  {32'h3fd363a8, 32'h40b32bfe} /* (19, 22, 9) {real, imag} */,
  {32'hbee3c368, 32'h4114e5d4} /* (19, 22, 8) {real, imag} */,
  {32'hbdce44a0, 32'h4108c0f2} /* (19, 22, 7) {real, imag} */,
  {32'h4077ecc6, 32'h3f630fc6} /* (19, 22, 6) {real, imag} */,
  {32'h40711af8, 32'hc05176fe} /* (19, 22, 5) {real, imag} */,
  {32'h4091685e, 32'hbef7a9df} /* (19, 22, 4) {real, imag} */,
  {32'h3fd0a13e, 32'hbe14e940} /* (19, 22, 3) {real, imag} */,
  {32'hc0623917, 32'hbf052228} /* (19, 22, 2) {real, imag} */,
  {32'hc02a082a, 32'h3f91de96} /* (19, 22, 1) {real, imag} */,
  {32'h3cfcb970, 32'h3fe1cf30} /* (19, 22, 0) {real, imag} */,
  {32'hbe360888, 32'h3ebf44a0} /* (19, 21, 31) {real, imag} */,
  {32'h406c0d40, 32'hc0095aa2} /* (19, 21, 30) {real, imag} */,
  {32'h3e464020, 32'h3e115cf0} /* (19, 21, 29) {real, imag} */,
  {32'hc0493425, 32'h4099c5b3} /* (19, 21, 28) {real, imag} */,
  {32'hbfae9f16, 32'h3f8f8bea} /* (19, 21, 27) {real, imag} */,
  {32'hc03e19ff, 32'hbfbc387c} /* (19, 21, 26) {real, imag} */,
  {32'hbff3eefe, 32'hc091b613} /* (19, 21, 25) {real, imag} */,
  {32'h3ed8b888, 32'hc01f3b38} /* (19, 21, 24) {real, imag} */,
  {32'h3dc92ba0, 32'hbdb9ae58} /* (19, 21, 23) {real, imag} */,
  {32'hbfab0bb9, 32'hbef81e8a} /* (19, 21, 22) {real, imag} */,
  {32'hbe965008, 32'hbea230b7} /* (19, 21, 21) {real, imag} */,
  {32'hc0778649, 32'h3f1b5f5e} /* (19, 21, 20) {real, imag} */,
  {32'hc067acb5, 32'hbfa13266} /* (19, 21, 19) {real, imag} */,
  {32'hbf9521d9, 32'hc0108964} /* (19, 21, 18) {real, imag} */,
  {32'hbf1d0360, 32'h3fc9dc58} /* (19, 21, 17) {real, imag} */,
  {32'h3f5c73d4, 32'hc00a43dd} /* (19, 21, 16) {real, imag} */,
  {32'hbe6511d8, 32'hc07142c7} /* (19, 21, 15) {real, imag} */,
  {32'hbd59f920, 32'hc0085356} /* (19, 21, 14) {real, imag} */,
  {32'h408c8744, 32'hbf311f24} /* (19, 21, 13) {real, imag} */,
  {32'h403ef012, 32'hbecbf90e} /* (19, 21, 12) {real, imag} */,
  {32'hbf471b3c, 32'hc00320f5} /* (19, 21, 11) {real, imag} */,
  {32'h3ee40b48, 32'hc0219062} /* (19, 21, 10) {real, imag} */,
  {32'h402bd830, 32'h405d2a00} /* (19, 21, 9) {real, imag} */,
  {32'h3df891a0, 32'h404d3ad5} /* (19, 21, 8) {real, imag} */,
  {32'hc02b448d, 32'h3f79de3c} /* (19, 21, 7) {real, imag} */,
  {32'hbfda88b8, 32'hbd98b820} /* (19, 21, 6) {real, imag} */,
  {32'h3ecb8bd0, 32'hc037e780} /* (19, 21, 5) {real, imag} */,
  {32'hbfbefaaa, 32'hc0819952} /* (19, 21, 4) {real, imag} */,
  {32'h4019b4a1, 32'h3f1e08b3} /* (19, 21, 3) {real, imag} */,
  {32'h4093ea13, 32'h40300d14} /* (19, 21, 2) {real, imag} */,
  {32'hbf56d65e, 32'h3f945e1c} /* (19, 21, 1) {real, imag} */,
  {32'hc02d774a, 32'h3f492806} /* (19, 21, 0) {real, imag} */,
  {32'hbfe30478, 32'hbf8d0d75} /* (19, 20, 31) {real, imag} */,
  {32'hbfbc4df0, 32'hbf28ae52} /* (19, 20, 30) {real, imag} */,
  {32'h3f854c50, 32'h3f85ed92} /* (19, 20, 29) {real, imag} */,
  {32'h3f0321fd, 32'h3e13a6e6} /* (19, 20, 28) {real, imag} */,
  {32'hbf33132c, 32'h3f25193a} /* (19, 20, 27) {real, imag} */,
  {32'h3f5a4404, 32'h3f3fbd9c} /* (19, 20, 26) {real, imag} */,
  {32'hbfe1c23a, 32'h3e9e9ea8} /* (19, 20, 25) {real, imag} */,
  {32'h3f5201a8, 32'h3edb7da2} /* (19, 20, 24) {real, imag} */,
  {32'h3fb9d77e, 32'h3f12d639} /* (19, 20, 23) {real, imag} */,
  {32'h3fb50200, 32'hbfa422cb} /* (19, 20, 22) {real, imag} */,
  {32'h3e51e638, 32'hbee76a6a} /* (19, 20, 21) {real, imag} */,
  {32'hbf8b52ad, 32'h401f4498} /* (19, 20, 20) {real, imag} */,
  {32'hbeaf1c28, 32'h3ee7a84f} /* (19, 20, 19) {real, imag} */,
  {32'hbeb5c51a, 32'hbfb686cb} /* (19, 20, 18) {real, imag} */,
  {32'hc0264cfa, 32'hbfd613ce} /* (19, 20, 17) {real, imag} */,
  {32'hc09af590, 32'hbfdeee00} /* (19, 20, 16) {real, imag} */,
  {32'hc000e0c8, 32'h3f991bd3} /* (19, 20, 15) {real, imag} */,
  {32'h40071670, 32'hbfa0c923} /* (19, 20, 14) {real, imag} */,
  {32'h3fd1a45f, 32'hbfc19aff} /* (19, 20, 13) {real, imag} */,
  {32'hc026f230, 32'hbe030088} /* (19, 20, 12) {real, imag} */,
  {32'hc029918b, 32'h401e3a6a} /* (19, 20, 11) {real, imag} */,
  {32'hc046e14a, 32'h40385376} /* (19, 20, 10) {real, imag} */,
  {32'hbe47fd24, 32'h3fdf5a79} /* (19, 20, 9) {real, imag} */,
  {32'hbfdacde5, 32'hbe655b14} /* (19, 20, 8) {real, imag} */,
  {32'hc0358a62, 32'hc064e69f} /* (19, 20, 7) {real, imag} */,
  {32'hbf7459b8, 32'hc0b3f9fa} /* (19, 20, 6) {real, imag} */,
  {32'h3f874a8b, 32'hc08b2fec} /* (19, 20, 5) {real, imag} */,
  {32'h3f1fdd99, 32'hbff988d5} /* (19, 20, 4) {real, imag} */,
  {32'h403212b4, 32'hbf906b56} /* (19, 20, 3) {real, imag} */,
  {32'h3f16876a, 32'h3e0f9b00} /* (19, 20, 2) {real, imag} */,
  {32'hbe43314c, 32'h3f230503} /* (19, 20, 1) {real, imag} */,
  {32'h3f8d7034, 32'h3ecf76d4} /* (19, 20, 0) {real, imag} */,
  {32'h3f4cd8b4, 32'h40335f41} /* (19, 19, 31) {real, imag} */,
  {32'h3f24c30e, 32'h402c3f88} /* (19, 19, 30) {real, imag} */,
  {32'hbf50792c, 32'h3f899f83} /* (19, 19, 29) {real, imag} */,
  {32'hbfafb519, 32'hbf80379b} /* (19, 19, 28) {real, imag} */,
  {32'h3ea89d34, 32'hbfd34a7c} /* (19, 19, 27) {real, imag} */,
  {32'hbfa607c3, 32'hbf0e2738} /* (19, 19, 26) {real, imag} */,
  {32'hc07992e7, 32'h3ffb6f91} /* (19, 19, 25) {real, imag} */,
  {32'hc048b8f2, 32'h3fceae51} /* (19, 19, 24) {real, imag} */,
  {32'hc00fdc03, 32'hbfbee54a} /* (19, 19, 23) {real, imag} */,
  {32'hbfaab6bf, 32'h3fefc7a0} /* (19, 19, 22) {real, imag} */,
  {32'hbf815ab5, 32'h4063d76f} /* (19, 19, 21) {real, imag} */,
  {32'hbfa3e940, 32'h3fff48a7} /* (19, 19, 20) {real, imag} */,
  {32'hbeb964c4, 32'h3fc7163d} /* (19, 19, 19) {real, imag} */,
  {32'h4008ac19, 32'h4016e6b7} /* (19, 19, 18) {real, imag} */,
  {32'h40832fc8, 32'h400049f9} /* (19, 19, 17) {real, imag} */,
  {32'h40050d74, 32'h3f8427c7} /* (19, 19, 16) {real, imag} */,
  {32'hc054bc9e, 32'hbf690478} /* (19, 19, 15) {real, imag} */,
  {32'hc07018ac, 32'h3f66b138} /* (19, 19, 14) {real, imag} */,
  {32'h3ec814a8, 32'hbee92f38} /* (19, 19, 13) {real, imag} */,
  {32'h3fae872a, 32'hbf40032c} /* (19, 19, 12) {real, imag} */,
  {32'hbfcfc787, 32'hc00f572c} /* (19, 19, 11) {real, imag} */,
  {32'hbf08d60a, 32'hbf126c45} /* (19, 19, 10) {real, imag} */,
  {32'hc044e640, 32'h3fc48dfa} /* (19, 19, 9) {real, imag} */,
  {32'hc00f7012, 32'h3e6fcdcc} /* (19, 19, 8) {real, imag} */,
  {32'hbeae7c8a, 32'hbda24f18} /* (19, 19, 7) {real, imag} */,
  {32'h3fb1ff4b, 32'hbf62cd47} /* (19, 19, 6) {real, imag} */,
  {32'h40166d1c, 32'hbe6ce5a0} /* (19, 19, 5) {real, imag} */,
  {32'h3e44c8b0, 32'hbfaf4b21} /* (19, 19, 4) {real, imag} */,
  {32'hc02224ba, 32'hc035cff8} /* (19, 19, 3) {real, imag} */,
  {32'hbf59f759, 32'hbfa67c20} /* (19, 19, 2) {real, imag} */,
  {32'h3edf5ae0, 32'hbf02f64a} /* (19, 19, 1) {real, imag} */,
  {32'hbe32eaa4, 32'h3fdf831c} /* (19, 19, 0) {real, imag} */,
  {32'hbf320184, 32'h3eca9fcc} /* (19, 18, 31) {real, imag} */,
  {32'hbf82d534, 32'h3ebef988} /* (19, 18, 30) {real, imag} */,
  {32'h3f9888e2, 32'h3e202d84} /* (19, 18, 29) {real, imag} */,
  {32'h3fc389f0, 32'hbfdf949a} /* (19, 18, 28) {real, imag} */,
  {32'h3e946974, 32'h3ea9e7f0} /* (19, 18, 27) {real, imag} */,
  {32'h3f4fb2a8, 32'h3ee968f0} /* (19, 18, 26) {real, imag} */,
  {32'h3ed85d32, 32'hbe8b78ac} /* (19, 18, 25) {real, imag} */,
  {32'h3ef51890, 32'h3fc33e25} /* (19, 18, 24) {real, imag} */,
  {32'h3fc12ada, 32'h400fdfed} /* (19, 18, 23) {real, imag} */,
  {32'h3fa38336, 32'h3f5fb240} /* (19, 18, 22) {real, imag} */,
  {32'h3fb0f17f, 32'hbf7031da} /* (19, 18, 21) {real, imag} */,
  {32'h3f605248, 32'h3f49c4de} /* (19, 18, 20) {real, imag} */,
  {32'hbf00e6e4, 32'h403ed926} /* (19, 18, 19) {real, imag} */,
  {32'h3ec636a7, 32'h3fa98b60} /* (19, 18, 18) {real, imag} */,
  {32'h3ef367d0, 32'h3ffc1e2a} /* (19, 18, 17) {real, imag} */,
  {32'hbd51d2e8, 32'h3f9f4fb0} /* (19, 18, 16) {real, imag} */,
  {32'hbf0d4668, 32'h3fb0e264} /* (19, 18, 15) {real, imag} */,
  {32'h3faab613, 32'h3f34e530} /* (19, 18, 14) {real, imag} */,
  {32'h402032a9, 32'h3f5c60da} /* (19, 18, 13) {real, imag} */,
  {32'h40324bfa, 32'h3db80870} /* (19, 18, 12) {real, imag} */,
  {32'h4041460c, 32'hbe97def4} /* (19, 18, 11) {real, imag} */,
  {32'h3e970068, 32'hbf9c0b88} /* (19, 18, 10) {real, imag} */,
  {32'h3cce7540, 32'hbf59af08} /* (19, 18, 9) {real, imag} */,
  {32'h3e524098, 32'hbe9693fc} /* (19, 18, 8) {real, imag} */,
  {32'hc000d3bc, 32'hbf43d9ec} /* (19, 18, 7) {real, imag} */,
  {32'hbfa293f2, 32'hbf92410f} /* (19, 18, 6) {real, imag} */,
  {32'hbf4e6c98, 32'h3f67b402} /* (19, 18, 5) {real, imag} */,
  {32'hbf161153, 32'h3fb89c9c} /* (19, 18, 4) {real, imag} */,
  {32'hbe60ba88, 32'h3f19eede} /* (19, 18, 3) {real, imag} */,
  {32'h3e9017b8, 32'hbeddd65a} /* (19, 18, 2) {real, imag} */,
  {32'h3f1ac0b2, 32'h3e3c6ca8} /* (19, 18, 1) {real, imag} */,
  {32'h3f6827f8, 32'h3fa35e30} /* (19, 18, 0) {real, imag} */,
  {32'h3d9d7818, 32'h3e4476a0} /* (19, 17, 31) {real, imag} */,
  {32'h3eda8c88, 32'hbec94cb0} /* (19, 17, 30) {real, imag} */,
  {32'hbeab1bcb, 32'hbd214600} /* (19, 17, 29) {real, imag} */,
  {32'hbf70f2f2, 32'h3fa3bcb4} /* (19, 17, 28) {real, imag} */,
  {32'hbfc3ef8a, 32'hbe6e51a0} /* (19, 17, 27) {real, imag} */,
  {32'h3f54bd6c, 32'h3f4fd1c2} /* (19, 17, 26) {real, imag} */,
  {32'h3f96c8b3, 32'h3fa6e141} /* (19, 17, 25) {real, imag} */,
  {32'h3fc2c06d, 32'h3cf007c0} /* (19, 17, 24) {real, imag} */,
  {32'h3eb6445e, 32'hbf03b0c3} /* (19, 17, 23) {real, imag} */,
  {32'hbede56c8, 32'hbe765cd0} /* (19, 17, 22) {real, imag} */,
  {32'hbd8848c0, 32'hbf93ebf5} /* (19, 17, 21) {real, imag} */,
  {32'h4030fa3a, 32'hbfbb9c95} /* (19, 17, 20) {real, imag} */,
  {32'h3fe11ab7, 32'hbdc9a0d8} /* (19, 17, 19) {real, imag} */,
  {32'h3f06c9b4, 32'h3f8a431b} /* (19, 17, 18) {real, imag} */,
  {32'h3f1d73ee, 32'hbf564fc0} /* (19, 17, 17) {real, imag} */,
  {32'h40005942, 32'h3e903f48} /* (19, 17, 16) {real, imag} */,
  {32'h400ac91c, 32'h3f931090} /* (19, 17, 15) {real, imag} */,
  {32'h3fad330e, 32'h3db5f1e4} /* (19, 17, 14) {real, imag} */,
  {32'hbd30a840, 32'h3f1dc9ce} /* (19, 17, 13) {real, imag} */,
  {32'hbe851d70, 32'h3cd44680} /* (19, 17, 12) {real, imag} */,
  {32'hbf836edc, 32'hbe9aa9c8} /* (19, 17, 11) {real, imag} */,
  {32'hbf58e878, 32'hbfabdc0e} /* (19, 17, 10) {real, imag} */,
  {32'h3fd217ba, 32'hbfb575f8} /* (19, 17, 9) {real, imag} */,
  {32'h4003c866, 32'hbf93d352} /* (19, 17, 8) {real, imag} */,
  {32'h3fed8038, 32'hbef7d674} /* (19, 17, 7) {real, imag} */,
  {32'h3fa558f5, 32'h3dcab758} /* (19, 17, 6) {real, imag} */,
  {32'h3ea10e18, 32'h3fa1f683} /* (19, 17, 5) {real, imag} */,
  {32'hbfcf22ad, 32'h3fcb997c} /* (19, 17, 4) {real, imag} */,
  {32'hbf5edbbe, 32'h3d467240} /* (19, 17, 3) {real, imag} */,
  {32'h3ec58688, 32'h3fe9fbb4} /* (19, 17, 2) {real, imag} */,
  {32'h3f3c7928, 32'h3fa3e0c0} /* (19, 17, 1) {real, imag} */,
  {32'h3ef003d4, 32'hbe85d09e} /* (19, 17, 0) {real, imag} */,
  {32'hbf730bc8, 32'hbe5c9380} /* (19, 16, 31) {real, imag} */,
  {32'hbfd79480, 32'h3f7ddda4} /* (19, 16, 30) {real, imag} */,
  {32'hbfd6d4e6, 32'hbd7297a0} /* (19, 16, 29) {real, imag} */,
  {32'h3d17d000, 32'h3e95b770} /* (19, 16, 28) {real, imag} */,
  {32'h3f21f448, 32'h3e832f34} /* (19, 16, 27) {real, imag} */,
  {32'h3f1dfc7f, 32'h3e983acc} /* (19, 16, 26) {real, imag} */,
  {32'hbf12d6b4, 32'hbf306c28} /* (19, 16, 25) {real, imag} */,
  {32'hbfc60a7e, 32'hbf17e69e} /* (19, 16, 24) {real, imag} */,
  {32'hbf972c10, 32'hbf4c9480} /* (19, 16, 23) {real, imag} */,
  {32'hbd883d80, 32'hbf17bc44} /* (19, 16, 22) {real, imag} */,
  {32'h3fb7273c, 32'h3f4cca40} /* (19, 16, 21) {real, imag} */,
  {32'h3f875d26, 32'h3fd0d81e} /* (19, 16, 20) {real, imag} */,
  {32'h3faf6830, 32'hbea774cc} /* (19, 16, 19) {real, imag} */,
  {32'h3fe031d4, 32'hbfbd9889} /* (19, 16, 18) {real, imag} */,
  {32'h3f9ee35c, 32'h3f2693c0} /* (19, 16, 17) {real, imag} */,
  {32'h3f1bc260, 32'h3feee08c} /* (19, 16, 16) {real, imag} */,
  {32'h401521a9, 32'h3f268bca} /* (19, 16, 15) {real, imag} */,
  {32'h3f31edcf, 32'hbfb276cc} /* (19, 16, 14) {real, imag} */,
  {32'hbf951414, 32'h3ec0bdd0} /* (19, 16, 13) {real, imag} */,
  {32'hbe24e290, 32'h3fb2dc5e} /* (19, 16, 12) {real, imag} */,
  {32'hbf4025d0, 32'h3ed9f9d0} /* (19, 16, 11) {real, imag} */,
  {32'hbfdb1634, 32'h3f974515} /* (19, 16, 10) {real, imag} */,
  {32'hbfed5fa8, 32'h3f96ea53} /* (19, 16, 9) {real, imag} */,
  {32'hbf425f20, 32'h3f40f7c0} /* (19, 16, 8) {real, imag} */,
  {32'h3e470af0, 32'h3f2703ea} /* (19, 16, 7) {real, imag} */,
  {32'h3de54aa0, 32'h402bb183} /* (19, 16, 6) {real, imag} */,
  {32'hbe683240, 32'hbfa5633c} /* (19, 16, 5) {real, imag} */,
  {32'hbe149230, 32'hbfbaf8c8} /* (19, 16, 4) {real, imag} */,
  {32'h3fd92332, 32'h3fb668c8} /* (19, 16, 3) {real, imag} */,
  {32'h402c4760, 32'h3ee51966} /* (19, 16, 2) {real, imag} */,
  {32'h40501649, 32'h3dc2a540} /* (19, 16, 1) {real, imag} */,
  {32'h3f8b35b4, 32'hbf1c54c8} /* (19, 16, 0) {real, imag} */,
  {32'hbf5f8d3d, 32'hbfabc7ec} /* (19, 15, 31) {real, imag} */,
  {32'hbf850a36, 32'hbfb7e91c} /* (19, 15, 30) {real, imag} */,
  {32'h3f141686, 32'hbfc5bf5a} /* (19, 15, 29) {real, imag} */,
  {32'h3f1eabee, 32'hbd986dc0} /* (19, 15, 28) {real, imag} */,
  {32'h3fc9922e, 32'h3f2eb6f8} /* (19, 15, 27) {real, imag} */,
  {32'h3fcaa34a, 32'h3fc3a615} /* (19, 15, 26) {real, imag} */,
  {32'h3f96117b, 32'h3f4ad636} /* (19, 15, 25) {real, imag} */,
  {32'h3f42b9aa, 32'h3e820f3c} /* (19, 15, 24) {real, imag} */,
  {32'h3f83820c, 32'hbdff19c8} /* (19, 15, 23) {real, imag} */,
  {32'hbec28df8, 32'hbe4fd110} /* (19, 15, 22) {real, imag} */,
  {32'hbfebde40, 32'hbed24e2c} /* (19, 15, 21) {real, imag} */,
  {32'hbf1a6066, 32'hbf86e90f} /* (19, 15, 20) {real, imag} */,
  {32'h3ed0ba2c, 32'hbf6f8eb5} /* (19, 15, 19) {real, imag} */,
  {32'hbba3c000, 32'h3f176cea} /* (19, 15, 18) {real, imag} */,
  {32'hbdfd29d0, 32'h40233510} /* (19, 15, 17) {real, imag} */,
  {32'h3f81fad4, 32'h4027ddb9} /* (19, 15, 16) {real, imag} */,
  {32'h3ffbfe0f, 32'h3fcb636c} /* (19, 15, 15) {real, imag} */,
  {32'h3fec72f6, 32'h3ebe9719} /* (19, 15, 14) {real, imag} */,
  {32'h3f109f9c, 32'h3eb65b01} /* (19, 15, 13) {real, imag} */,
  {32'h3f654888, 32'hbec0e1b0} /* (19, 15, 12) {real, imag} */,
  {32'hbd93c548, 32'hbf24ca14} /* (19, 15, 11) {real, imag} */,
  {32'hbf134f08, 32'hbf5d762c} /* (19, 15, 10) {real, imag} */,
  {32'h3daf5a08, 32'hbf9161e0} /* (19, 15, 9) {real, imag} */,
  {32'hbf2a8524, 32'hbf3f25f4} /* (19, 15, 8) {real, imag} */,
  {32'hbf1b8dd3, 32'hbedca48c} /* (19, 15, 7) {real, imag} */,
  {32'hbfc6929f, 32'hbf813a62} /* (19, 15, 6) {real, imag} */,
  {32'hbf92db82, 32'h3f2ce4b2} /* (19, 15, 5) {real, imag} */,
  {32'h3e5ac948, 32'h3ebebc32} /* (19, 15, 4) {real, imag} */,
  {32'h3fc8bf91, 32'h401f912f} /* (19, 15, 3) {real, imag} */,
  {32'h3e96b720, 32'h3f5cda48} /* (19, 15, 2) {real, imag} */,
  {32'hbdd79a00, 32'hbf385888} /* (19, 15, 1) {real, imag} */,
  {32'hbe111078, 32'hbf8f2ca8} /* (19, 15, 0) {real, imag} */,
  {32'h3fb3e836, 32'h3d9d5750} /* (19, 14, 31) {real, imag} */,
  {32'h3f047248, 32'hbdcf1460} /* (19, 14, 30) {real, imag} */,
  {32'hbfe8ec24, 32'h3f163489} /* (19, 14, 29) {real, imag} */,
  {32'h3f9bd55c, 32'h3f2ee5fc} /* (19, 14, 28) {real, imag} */,
  {32'h4003c86e, 32'hbeb5bd40} /* (19, 14, 27) {real, imag} */,
  {32'h401e90ae, 32'hbfe808ee} /* (19, 14, 26) {real, imag} */,
  {32'h3fd1f324, 32'h3fc9dc5d} /* (19, 14, 25) {real, imag} */,
  {32'hbf224014, 32'h400bf09a} /* (19, 14, 24) {real, imag} */,
  {32'hbf4b9a6c, 32'hbf25c154} /* (19, 14, 23) {real, imag} */,
  {32'hbcaf8a80, 32'hbf7edc30} /* (19, 14, 22) {real, imag} */,
  {32'hbf936d61, 32'h3f603f86} /* (19, 14, 21) {real, imag} */,
  {32'hbfc9cde8, 32'hbe0c2c4a} /* (19, 14, 20) {real, imag} */,
  {32'hbf5c2bd8, 32'h4009c8c2} /* (19, 14, 19) {real, imag} */,
  {32'h3f40bc08, 32'h3fb67c8c} /* (19, 14, 18) {real, imag} */,
  {32'h3faf126c, 32'hbf841d18} /* (19, 14, 17) {real, imag} */,
  {32'h3f16a354, 32'h3d28f080} /* (19, 14, 16) {real, imag} */,
  {32'h3ee5c9f0, 32'hbe2637c0} /* (19, 14, 15) {real, imag} */,
  {32'hbf75df3a, 32'hbf98fec4} /* (19, 14, 14) {real, imag} */,
  {32'hbfcd0abe, 32'h3d697920} /* (19, 14, 13) {real, imag} */,
  {32'hbf180558, 32'h3fd5f503} /* (19, 14, 12) {real, imag} */,
  {32'hbf22d996, 32'hbfc610a5} /* (19, 14, 11) {real, imag} */,
  {32'hbf45e56c, 32'hc05d6664} /* (19, 14, 10) {real, imag} */,
  {32'h3f36e51a, 32'hbf3951f0} /* (19, 14, 9) {real, imag} */,
  {32'h404b5c00, 32'hbdce6010} /* (19, 14, 8) {real, imag} */,
  {32'hbec90218, 32'h3f092ff4} /* (19, 14, 7) {real, imag} */,
  {32'hbf682d3c, 32'h3fc6030f} /* (19, 14, 6) {real, imag} */,
  {32'h3fa0c498, 32'h40729e9c} /* (19, 14, 5) {real, imag} */,
  {32'h3f9ba3d8, 32'h3f957808} /* (19, 14, 4) {real, imag} */,
  {32'hc02277cc, 32'hbdeabe50} /* (19, 14, 3) {real, imag} */,
  {32'hc03c3be1, 32'h3f5ef645} /* (19, 14, 2) {real, imag} */,
  {32'hc00a8940, 32'h3ff0441f} /* (19, 14, 1) {real, imag} */,
  {32'hbfaa43c0, 32'h3f80653c} /* (19, 14, 0) {real, imag} */,
  {32'hbf90d3fd, 32'h3fc0313e} /* (19, 13, 31) {real, imag} */,
  {32'hbe3c4328, 32'hbbb71e00} /* (19, 13, 30) {real, imag} */,
  {32'h3f57f6d0, 32'hbf5a84f2} /* (19, 13, 29) {real, imag} */,
  {32'h3ded2470, 32'h3f6f198e} /* (19, 13, 28) {real, imag} */,
  {32'h3cc3b940, 32'h3ec90e68} /* (19, 13, 27) {real, imag} */,
  {32'h3f9d4f8d, 32'h3fefae00} /* (19, 13, 26) {real, imag} */,
  {32'hbcab9f80, 32'h40713420} /* (19, 13, 25) {real, imag} */,
  {32'hc001b4ca, 32'h3ffe4887} /* (19, 13, 24) {real, imag} */,
  {32'hbf523d51, 32'h3f26d5e4} /* (19, 13, 23) {real, imag} */,
  {32'h3ed6809c, 32'hbdaa7bd8} /* (19, 13, 22) {real, imag} */,
  {32'hbf409822, 32'hbfe6732a} /* (19, 13, 21) {real, imag} */,
  {32'hc0016ef0, 32'hbf602576} /* (19, 13, 20) {real, imag} */,
  {32'hc0469c2e, 32'hbf63d886} /* (19, 13, 19) {real, imag} */,
  {32'hbf97f288, 32'hbf8aefd6} /* (19, 13, 18) {real, imag} */,
  {32'h40077408, 32'h3f5f60c4} /* (19, 13, 17) {real, imag} */,
  {32'h3f1e0a80, 32'h3dd06350} /* (19, 13, 16) {real, imag} */,
  {32'h3e89ebe4, 32'hc01497e7} /* (19, 13, 15) {real, imag} */,
  {32'hbfa9cb54, 32'hbfe454ca} /* (19, 13, 14) {real, imag} */,
  {32'h3db6aee0, 32'h3fb6a712} /* (19, 13, 13) {real, imag} */,
  {32'h3d7acb80, 32'h3fc5e7d2} /* (19, 13, 12) {real, imag} */,
  {32'h3f88ea89, 32'h3f2fc94e} /* (19, 13, 11) {real, imag} */,
  {32'hbf6c485e, 32'hbf75800d} /* (19, 13, 10) {real, imag} */,
  {32'hc00bfeec, 32'hbe9ca744} /* (19, 13, 9) {real, imag} */,
  {32'h3dbf2170, 32'hbc099740} /* (19, 13, 8) {real, imag} */,
  {32'hbf6d0123, 32'h3e66989c} /* (19, 13, 7) {real, imag} */,
  {32'hbfad03f3, 32'hbfd79b96} /* (19, 13, 6) {real, imag} */,
  {32'h3ece035c, 32'h3eb11008} /* (19, 13, 5) {real, imag} */,
  {32'h40151a52, 32'h3f69a6aa} /* (19, 13, 4) {real, imag} */,
  {32'h3f207e56, 32'h40014010} /* (19, 13, 3) {real, imag} */,
  {32'hbdf1be38, 32'h4003f188} /* (19, 13, 2) {real, imag} */,
  {32'hbf433190, 32'h3fc5bba7} /* (19, 13, 1) {real, imag} */,
  {32'hbfe5daa6, 32'h4003919b} /* (19, 13, 0) {real, imag} */,
  {32'hbe06c1ec, 32'hbd8ed7f0} /* (19, 12, 31) {real, imag} */,
  {32'hbf4b8ee0, 32'h3dfdf530} /* (19, 12, 30) {real, imag} */,
  {32'hbf8e8b58, 32'hbf1d9440} /* (19, 12, 29) {real, imag} */,
  {32'hbe1d7394, 32'h3e9f8833} /* (19, 12, 28) {real, imag} */,
  {32'hbf3dc918, 32'h3fd26631} /* (19, 12, 27) {real, imag} */,
  {32'h3e178610, 32'h3f94e7a6} /* (19, 12, 26) {real, imag} */,
  {32'hbf56e658, 32'hbf0a5910} /* (19, 12, 25) {real, imag} */,
  {32'hc0096b0b, 32'hbf6a119f} /* (19, 12, 24) {real, imag} */,
  {32'hbe602df0, 32'hbf397413} /* (19, 12, 23) {real, imag} */,
  {32'h4080f3ed, 32'hbf6ec776} /* (19, 12, 22) {real, imag} */,
  {32'h4040eb0e, 32'hbf14fc0d} /* (19, 12, 21) {real, imag} */,
  {32'hbf90c287, 32'h3f9d78ae} /* (19, 12, 20) {real, imag} */,
  {32'hbf85d266, 32'h3fa18b58} /* (19, 12, 19) {real, imag} */,
  {32'hc00d1426, 32'hc022a09c} /* (19, 12, 18) {real, imag} */,
  {32'hbfc90c87, 32'hc0875542} /* (19, 12, 17) {real, imag} */,
  {32'hbfa0b456, 32'hbff6db54} /* (19, 12, 16) {real, imag} */,
  {32'hbfd6857b, 32'h3fa51739} /* (19, 12, 15) {real, imag} */,
  {32'hbe1f1f68, 32'h3fa781e7} /* (19, 12, 14) {real, imag} */,
  {32'h400468c8, 32'h3e3cfec8} /* (19, 12, 13) {real, imag} */,
  {32'h4058807c, 32'hc060ab16} /* (19, 12, 12) {real, imag} */,
  {32'h3ff19446, 32'hbff3a547} /* (19, 12, 11) {real, imag} */,
  {32'h3fcbff24, 32'h3f70fa03} /* (19, 12, 10) {real, imag} */,
  {32'h3fda3160, 32'hbee17b8c} /* (19, 12, 9) {real, imag} */,
  {32'h3f787fb6, 32'h3fad6998} /* (19, 12, 8) {real, imag} */,
  {32'hbfc12863, 32'h3f49abb4} /* (19, 12, 7) {real, imag} */,
  {32'hc04b9592, 32'hbfb693fe} /* (19, 12, 6) {real, imag} */,
  {32'hbf2dbc9e, 32'hbe0da890} /* (19, 12, 5) {real, imag} */,
  {32'hbd853898, 32'h3ff8e111} /* (19, 12, 4) {real, imag} */,
  {32'hbf9f762f, 32'hbfe76b76} /* (19, 12, 3) {real, imag} */,
  {32'hbfbe6a65, 32'hbfced238} /* (19, 12, 2) {real, imag} */,
  {32'hc0080998, 32'hbec01bbe} /* (19, 12, 1) {real, imag} */,
  {32'h3e8d6082, 32'hbe0a6f08} /* (19, 12, 0) {real, imag} */,
  {32'hbf612eca, 32'hbfd95194} /* (19, 11, 31) {real, imag} */,
  {32'hc01860c8, 32'hc046b2dc} /* (19, 11, 30) {real, imag} */,
  {32'h3ea6e270, 32'hbfa87d02} /* (19, 11, 29) {real, imag} */,
  {32'hc01cbeeb, 32'h3fbbeb49} /* (19, 11, 28) {real, imag} */,
  {32'hc0d3899e, 32'h40687cff} /* (19, 11, 27) {real, imag} */,
  {32'hc08c64de, 32'h406f856a} /* (19, 11, 26) {real, imag} */,
  {32'hbff0fa1a, 32'h40248316} /* (19, 11, 25) {real, imag} */,
  {32'h3fcc9a54, 32'h405ad380} /* (19, 11, 24) {real, imag} */,
  {32'h4083bc48, 32'hbfc42174} /* (19, 11, 23) {real, imag} */,
  {32'h404bea90, 32'hc00e112c} /* (19, 11, 22) {real, imag} */,
  {32'h3f6da69c, 32'hbd45ea48} /* (19, 11, 21) {real, imag} */,
  {32'hbfb24946, 32'hbf8c70c7} /* (19, 11, 20) {real, imag} */,
  {32'hbfe09b8e, 32'h3da539a0} /* (19, 11, 19) {real, imag} */,
  {32'h3fa43af3, 32'hc05c83a0} /* (19, 11, 18) {real, imag} */,
  {32'h3fc6fea8, 32'hc0541988} /* (19, 11, 17) {real, imag} */,
  {32'hbfdada9e, 32'h3eaedb8e} /* (19, 11, 16) {real, imag} */,
  {32'hc0489650, 32'h406412ad} /* (19, 11, 15) {real, imag} */,
  {32'hbf94ff43, 32'h4000c81a} /* (19, 11, 14) {real, imag} */,
  {32'h3f4b13c0, 32'hbf93a117} /* (19, 11, 13) {real, imag} */,
  {32'h4050c19e, 32'hbf809a7c} /* (19, 11, 12) {real, imag} */,
  {32'h3ff428ba, 32'h403a26cd} /* (19, 11, 11) {real, imag} */,
  {32'hbfe7eb8c, 32'h40349886} /* (19, 11, 10) {real, imag} */,
  {32'hc0043200, 32'hbf93b060} /* (19, 11, 9) {real, imag} */,
  {32'hbea82db8, 32'hc0809900} /* (19, 11, 8) {real, imag} */,
  {32'hbfc802ea, 32'h3fb8de5a} /* (19, 11, 7) {real, imag} */,
  {32'hbf3a40bc, 32'h4011cd03} /* (19, 11, 6) {real, imag} */,
  {32'h4039e1a4, 32'h400e44c0} /* (19, 11, 5) {real, imag} */,
  {32'hbef36d8a, 32'h3f8626da} /* (19, 11, 4) {real, imag} */,
  {32'h3fbe2a7e, 32'hc002ac8c} /* (19, 11, 3) {real, imag} */,
  {32'h403da331, 32'hbfded9a4} /* (19, 11, 2) {real, imag} */,
  {32'h4030c5f0, 32'hbff3d264} /* (19, 11, 1) {real, imag} */,
  {32'h401b7b1a, 32'hbf9ac2be} /* (19, 11, 0) {real, imag} */,
  {32'h404d5a43, 32'h40269290} /* (19, 10, 31) {real, imag} */,
  {32'h3f8244c2, 32'h3f93385b} /* (19, 10, 30) {real, imag} */,
  {32'hc06ee542, 32'h3f2f7a64} /* (19, 10, 29) {real, imag} */,
  {32'hbe24df88, 32'h3fa51784} /* (19, 10, 28) {real, imag} */,
  {32'hc04020a8, 32'hc0bdd5be} /* (19, 10, 27) {real, imag} */,
  {32'hc07759d6, 32'hc06e3db7} /* (19, 10, 26) {real, imag} */,
  {32'h400ac332, 32'h4023d814} /* (19, 10, 25) {real, imag} */,
  {32'h40229672, 32'h3fb04d65} /* (19, 10, 24) {real, imag} */,
  {32'hbf3f4570, 32'h400dea35} /* (19, 10, 23) {real, imag} */,
  {32'h3dda0f30, 32'h407501d0} /* (19, 10, 22) {real, imag} */,
  {32'h3fcf4864, 32'hbf08ef0e} /* (19, 10, 21) {real, imag} */,
  {32'h3f2ad0b8, 32'hc0180990} /* (19, 10, 20) {real, imag} */,
  {32'h4032e567, 32'hbfc80e52} /* (19, 10, 19) {real, imag} */,
  {32'h3ecfdebc, 32'h403b659e} /* (19, 10, 18) {real, imag} */,
  {32'h3dbb4fa0, 32'h407e8ac0} /* (19, 10, 17) {real, imag} */,
  {32'h3efb21a0, 32'h3fcae974} /* (19, 10, 16) {real, imag} */,
  {32'hc02784da, 32'h3f3fe7d4} /* (19, 10, 15) {real, imag} */,
  {32'h3fdda218, 32'hbf1f0a4c} /* (19, 10, 14) {real, imag} */,
  {32'h403a755a, 32'h4017e319} /* (19, 10, 13) {real, imag} */,
  {32'h404d345d, 32'h3ff88dcc} /* (19, 10, 12) {real, imag} */,
  {32'h402b9f1c, 32'h3f8205dd} /* (19, 10, 11) {real, imag} */,
  {32'h40777ee4, 32'h3f629daa} /* (19, 10, 10) {real, imag} */,
  {32'h406c962c, 32'h3ff17a40} /* (19, 10, 9) {real, imag} */,
  {32'h40c05450, 32'h402a5aab} /* (19, 10, 8) {real, imag} */,
  {32'h408e6798, 32'h3fbdac8c} /* (19, 10, 7) {real, imag} */,
  {32'hbff66779, 32'h3d814e90} /* (19, 10, 6) {real, imag} */,
  {32'hbef8bd7c, 32'hbf8ca4cb} /* (19, 10, 5) {real, imag} */,
  {32'hbf7787e0, 32'h3e1f1fda} /* (19, 10, 4) {real, imag} */,
  {32'h3fb8fe7a, 32'h4013e4c8} /* (19, 10, 3) {real, imag} */,
  {32'hbfc4724e, 32'h3fd71398} /* (19, 10, 2) {real, imag} */,
  {32'hbfc0d43c, 32'h3d48f9c0} /* (19, 10, 1) {real, imag} */,
  {32'hbf283358, 32'hbd9e1a68} /* (19, 10, 0) {real, imag} */,
  {32'h3ff0798b, 32'hbfd84f04} /* (19, 9, 31) {real, imag} */,
  {32'h3eba5390, 32'hc07fde1e} /* (19, 9, 30) {real, imag} */,
  {32'hbfec023a, 32'hbfe905dc} /* (19, 9, 29) {real, imag} */,
  {32'hc10114fc, 32'hc0118d78} /* (19, 9, 28) {real, imag} */,
  {32'h3e92b314, 32'hbf853fb4} /* (19, 9, 27) {real, imag} */,
  {32'hc0003d45, 32'h407fdc9b} /* (19, 9, 26) {real, imag} */,
  {32'hc0b05f34, 32'hbfa2a323} /* (19, 9, 25) {real, imag} */,
  {32'hbf7f7340, 32'h3ff0837a} /* (19, 9, 24) {real, imag} */,
  {32'h402f5ddf, 32'h3fda811a} /* (19, 9, 23) {real, imag} */,
  {32'h3fb8e97a, 32'h40625682} /* (19, 9, 22) {real, imag} */,
  {32'hbfed4ffd, 32'h401720b7} /* (19, 9, 21) {real, imag} */,
  {32'h3feab996, 32'hbfd9293a} /* (19, 9, 20) {real, imag} */,
  {32'h4021f22b, 32'hbfcc2a25} /* (19, 9, 19) {real, imag} */,
  {32'h4039f86c, 32'hbfb06e38} /* (19, 9, 18) {real, imag} */,
  {32'hbea3c3fe, 32'h40b3e40e} /* (19, 9, 17) {real, imag} */,
  {32'h3f7fb99e, 32'h40bd8978} /* (19, 9, 16) {real, imag} */,
  {32'h4081a81a, 32'h3efd0762} /* (19, 9, 15) {real, imag} */,
  {32'hbfe8a774, 32'hc00b89b5} /* (19, 9, 14) {real, imag} */,
  {32'hc000f186, 32'hbf89db44} /* (19, 9, 13) {real, imag} */,
  {32'h3ff9d28d, 32'h40915608} /* (19, 9, 12) {real, imag} */,
  {32'hbf9cbce2, 32'h408e3c9a} /* (19, 9, 11) {real, imag} */,
  {32'hc07179f8, 32'h3facbfde} /* (19, 9, 10) {real, imag} */,
  {32'hc06fb66f, 32'hc028fff2} /* (19, 9, 9) {real, imag} */,
  {32'hbf5239fc, 32'hc08c6618} /* (19, 9, 8) {real, imag} */,
  {32'h3f841982, 32'hc0c4cf54} /* (19, 9, 7) {real, imag} */,
  {32'hc0198be1, 32'hc008f81b} /* (19, 9, 6) {real, imag} */,
  {32'hbf1cbf0c, 32'hbf7226a8} /* (19, 9, 5) {real, imag} */,
  {32'h401c4243, 32'hc063e129} /* (19, 9, 4) {real, imag} */,
  {32'h4032de40, 32'hc0b6c43b} /* (19, 9, 3) {real, imag} */,
  {32'h3e316890, 32'hc0ecd84d} /* (19, 9, 2) {real, imag} */,
  {32'h3f366144, 32'hc064f964} /* (19, 9, 1) {real, imag} */,
  {32'h3fba7007, 32'h3f003239} /* (19, 9, 0) {real, imag} */,
  {32'hbf0b8ffc, 32'h40181147} /* (19, 8, 31) {real, imag} */,
  {32'hc017c562, 32'h405a264f} /* (19, 8, 30) {real, imag} */,
  {32'h3f32e3ea, 32'h410579bc} /* (19, 8, 29) {real, imag} */,
  {32'h3fe72f11, 32'h4061afeb} /* (19, 8, 28) {real, imag} */,
  {32'hc08cafae, 32'h4019f1d2} /* (19, 8, 27) {real, imag} */,
  {32'hc075bda8, 32'hc00b1006} /* (19, 8, 26) {real, imag} */,
  {32'h400f7cac, 32'hbfb4a34d} /* (19, 8, 25) {real, imag} */,
  {32'h4065c0a8, 32'h3dfa4d70} /* (19, 8, 24) {real, imag} */,
  {32'h40349a0d, 32'hc08006c8} /* (19, 8, 23) {real, imag} */,
  {32'hc077a8fc, 32'hc07f1b30} /* (19, 8, 22) {real, imag} */,
  {32'hc0242fb2, 32'hbf4a8834} /* (19, 8, 21) {real, imag} */,
  {32'h3e8a390c, 32'h401d151f} /* (19, 8, 20) {real, imag} */,
  {32'hc05c5e23, 32'h3f225630} /* (19, 8, 19) {real, imag} */,
  {32'hbf1a01f0, 32'hc01619f6} /* (19, 8, 18) {real, imag} */,
  {32'h402d7f92, 32'hbe7ef600} /* (19, 8, 17) {real, imag} */,
  {32'h403a401b, 32'hc0895fbb} /* (19, 8, 16) {real, imag} */,
  {32'h3ff204a6, 32'h3f949f0f} /* (19, 8, 15) {real, imag} */,
  {32'hbedfe694, 32'h4083a62c} /* (19, 8, 14) {real, imag} */,
  {32'hbdfbbfd0, 32'h40a2cf8a} /* (19, 8, 13) {real, imag} */,
  {32'h40681d42, 32'h40242841} /* (19, 8, 12) {real, imag} */,
  {32'h3f812e18, 32'hc0ada5a4} /* (19, 8, 11) {real, imag} */,
  {32'hbef0db00, 32'h3ea2afc4} /* (19, 8, 10) {real, imag} */,
  {32'h3f9e3414, 32'h3e5d6508} /* (19, 8, 9) {real, imag} */,
  {32'h4042a8ba, 32'hbfa40806} /* (19, 8, 8) {real, imag} */,
  {32'h3f68fd68, 32'hc010ead4} /* (19, 8, 7) {real, imag} */,
  {32'h3ff733ae, 32'hbfe2355f} /* (19, 8, 6) {real, imag} */,
  {32'h406b6b64, 32'h3f54a94e} /* (19, 8, 5) {real, imag} */,
  {32'h3f052ed8, 32'h3ffc88d4} /* (19, 8, 4) {real, imag} */,
  {32'h3ea43c14, 32'hbed03308} /* (19, 8, 3) {real, imag} */,
  {32'hc00592ce, 32'hbfd792a0} /* (19, 8, 2) {real, imag} */,
  {32'hbff15038, 32'h3f7a1db0} /* (19, 8, 1) {real, imag} */,
  {32'hb9b9a000, 32'h402f8ee4} /* (19, 8, 0) {real, imag} */,
  {32'hc0e4923e, 32'h40318096} /* (19, 7, 31) {real, imag} */,
  {32'hc08e7f43, 32'h4040b116} /* (19, 7, 30) {real, imag} */,
  {32'h40ff88ac, 32'h3f9b95fc} /* (19, 7, 29) {real, imag} */,
  {32'h3ffe1c44, 32'h3ffb0a12} /* (19, 7, 28) {real, imag} */,
  {32'hc00d36da, 32'h3ec6e2f4} /* (19, 7, 27) {real, imag} */,
  {32'h402e42fc, 32'h3ecf8998} /* (19, 7, 26) {real, imag} */,
  {32'h4057d498, 32'h3f317402} /* (19, 7, 25) {real, imag} */,
  {32'h40c272f9, 32'h3f9b163c} /* (19, 7, 24) {real, imag} */,
  {32'h411005fa, 32'h401bf6df} /* (19, 7, 23) {real, imag} */,
  {32'h40aaf134, 32'h406ba868} /* (19, 7, 22) {real, imag} */,
  {32'hc09a599c, 32'hbf2f6c80} /* (19, 7, 21) {real, imag} */,
  {32'hc1057bd6, 32'hc09be944} /* (19, 7, 20) {real, imag} */,
  {32'hc0a9bb77, 32'hc083bcd4} /* (19, 7, 19) {real, imag} */,
  {32'hbf70fd04, 32'h3f1e1502} /* (19, 7, 18) {real, imag} */,
  {32'h3fa65c4c, 32'h3f7a5c12} /* (19, 7, 17) {real, imag} */,
  {32'h3fe6c443, 32'h3f5b501c} /* (19, 7, 16) {real, imag} */,
  {32'h3ea3f4e0, 32'hc0496d76} /* (19, 7, 15) {real, imag} */,
  {32'h3fd747a0, 32'h3eddc2d8} /* (19, 7, 14) {real, imag} */,
  {32'h409ee085, 32'h4039865b} /* (19, 7, 13) {real, imag} */,
  {32'h409b7a9a, 32'h404ada58} /* (19, 7, 12) {real, imag} */,
  {32'h40806007, 32'h406e06af} /* (19, 7, 11) {real, imag} */,
  {32'h40aefb94, 32'h4025cfd1} /* (19, 7, 10) {real, imag} */,
  {32'h3f627ebc, 32'h4121df5d} /* (19, 7, 9) {real, imag} */,
  {32'hbf8be400, 32'h40ccb0c2} /* (19, 7, 8) {real, imag} */,
  {32'h3e841148, 32'hc07b93a0} /* (19, 7, 7) {real, imag} */,
  {32'h3f853b02, 32'hc0e83d30} /* (19, 7, 6) {real, imag} */,
  {32'h3fb8e5fe, 32'hc07eeeb5} /* (19, 7, 5) {real, imag} */,
  {32'hbfed93ac, 32'hbf109220} /* (19, 7, 4) {real, imag} */,
  {32'hbfd01d88, 32'hc010a11b} /* (19, 7, 3) {real, imag} */,
  {32'hbfa8755f, 32'hc04d3344} /* (19, 7, 2) {real, imag} */,
  {32'hc0c4674f, 32'hc04764bb} /* (19, 7, 1) {real, imag} */,
  {32'hc04b7f2f, 32'hbf7ecf2d} /* (19, 7, 0) {real, imag} */,
  {32'h3f59fa64, 32'hc0243f48} /* (19, 6, 31) {real, imag} */,
  {32'h4028eba4, 32'hbe89c0c4} /* (19, 6, 30) {real, imag} */,
  {32'h4059d794, 32'hbf8809d0} /* (19, 6, 29) {real, imag} */,
  {32'hbf84398c, 32'h3f77cb24} /* (19, 6, 28) {real, imag} */,
  {32'h3f5454f6, 32'h40f70614} /* (19, 6, 27) {real, imag} */,
  {32'h40900e36, 32'h40531cf1} /* (19, 6, 26) {real, imag} */,
  {32'hbf8d7010, 32'h3f871e90} /* (19, 6, 25) {real, imag} */,
  {32'h4090a121, 32'h3e1fc060} /* (19, 6, 24) {real, imag} */,
  {32'hbf554420, 32'h3fcd0c63} /* (19, 6, 23) {real, imag} */,
  {32'hc08864b8, 32'hbeda8c50} /* (19, 6, 22) {real, imag} */,
  {32'hc095ba3e, 32'h3f82606c} /* (19, 6, 21) {real, imag} */,
  {32'h40092d96, 32'h40818ab9} /* (19, 6, 20) {real, imag} */,
  {32'h40048078, 32'h3e97dd3e} /* (19, 6, 19) {real, imag} */,
  {32'hc05aa73e, 32'h410bf982} /* (19, 6, 18) {real, imag} */,
  {32'hc10a5b92, 32'h4110a396} /* (19, 6, 17) {real, imag} */,
  {32'hc0d37558, 32'h40a7f748} /* (19, 6, 16) {real, imag} */,
  {32'h3ea77344, 32'h3f4aca8b} /* (19, 6, 15) {real, imag} */,
  {32'hbfbeb913, 32'h40b24230} /* (19, 6, 14) {real, imag} */,
  {32'hc0b5f6fc, 32'h408aeb84} /* (19, 6, 13) {real, imag} */,
  {32'hc050a5af, 32'hbf8bcb3e} /* (19, 6, 12) {real, imag} */,
  {32'h3f73aff0, 32'h3fa5e5e4} /* (19, 6, 11) {real, imag} */,
  {32'hc0596ff2, 32'h40a44ae9} /* (19, 6, 10) {real, imag} */,
  {32'hbcb56900, 32'h40ff6b5b} /* (19, 6, 9) {real, imag} */,
  {32'h40ac654d, 32'h40a8d5d1} /* (19, 6, 8) {real, imag} */,
  {32'h40146118, 32'h3fa95f88} /* (19, 6, 7) {real, imag} */,
  {32'hbf10c384, 32'h3f645e7c} /* (19, 6, 6) {real, imag} */,
  {32'h3d77cd00, 32'hc0ab387a} /* (19, 6, 5) {real, imag} */,
  {32'hbf86be0c, 32'hbfe68e21} /* (19, 6, 4) {real, imag} */,
  {32'h4080a06e, 32'hbff8255a} /* (19, 6, 3) {real, imag} */,
  {32'h40fa59ae, 32'hc0903bca} /* (19, 6, 2) {real, imag} */,
  {32'h40a1519b, 32'hc12d6450} /* (19, 6, 1) {real, imag} */,
  {32'h3e707862, 32'hc06aac38} /* (19, 6, 0) {real, imag} */,
  {32'hbfc5d729, 32'h3fa0ee40} /* (19, 5, 31) {real, imag} */,
  {32'hbe66f720, 32'hc0278779} /* (19, 5, 30) {real, imag} */,
  {32'h409e254e, 32'hc08d0554} /* (19, 5, 29) {real, imag} */,
  {32'hc06d71e4, 32'hc0885764} /* (19, 5, 28) {real, imag} */,
  {32'h3fc97246, 32'h3f5e3ea8} /* (19, 5, 27) {real, imag} */,
  {32'h4103635e, 32'h406e8584} /* (19, 5, 26) {real, imag} */,
  {32'h40565faa, 32'h40b52b28} /* (19, 5, 25) {real, imag} */,
  {32'hc0020020, 32'h403f0813} /* (19, 5, 24) {real, imag} */,
  {32'hbfb394ca, 32'h4082dd15} /* (19, 5, 23) {real, imag} */,
  {32'h40988bc2, 32'h3fa01b20} /* (19, 5, 22) {real, imag} */,
  {32'h405b4234, 32'hbfdc9bc8} /* (19, 5, 21) {real, imag} */,
  {32'h3b77f400, 32'h3fdca927} /* (19, 5, 20) {real, imag} */,
  {32'hbf8a88bc, 32'h3e584900} /* (19, 5, 19) {real, imag} */,
  {32'hbed0ab70, 32'hc06e3eda} /* (19, 5, 18) {real, imag} */,
  {32'hbfacf9ea, 32'hc03d737c} /* (19, 5, 17) {real, imag} */,
  {32'hc0b4e943, 32'hbfb67f9a} /* (19, 5, 16) {real, imag} */,
  {32'hc0a4ceec, 32'h40ed8a54} /* (19, 5, 15) {real, imag} */,
  {32'hc10a82b0, 32'h40fba09c} /* (19, 5, 14) {real, imag} */,
  {32'hc0a6a0e2, 32'hbd83d860} /* (19, 5, 13) {real, imag} */,
  {32'h3f350ed8, 32'hc03f2b22} /* (19, 5, 12) {real, imag} */,
  {32'h40013036, 32'hc0c4417a} /* (19, 5, 11) {real, imag} */,
  {32'h3fe07d34, 32'hc111f87d} /* (19, 5, 10) {real, imag} */,
  {32'hc0a0da4d, 32'hc00ab0d0} /* (19, 5, 9) {real, imag} */,
  {32'hc110e298, 32'h414d233a} /* (19, 5, 8) {real, imag} */,
  {32'hc0d3269c, 32'h40ee966c} /* (19, 5, 7) {real, imag} */,
  {32'h40235880, 32'hc04300fe} /* (19, 5, 6) {real, imag} */,
  {32'hc104f90c, 32'h3f3263d2} /* (19, 5, 5) {real, imag} */,
  {32'hc0e6af19, 32'h4053be2c} /* (19, 5, 4) {real, imag} */,
  {32'hbfad7028, 32'h3ece7fae} /* (19, 5, 3) {real, imag} */,
  {32'h405bb887, 32'h3fbd940a} /* (19, 5, 2) {real, imag} */,
  {32'hbe872ff0, 32'h40f7f28b} /* (19, 5, 1) {real, imag} */,
  {32'hc05450e0, 32'h3f87bcba} /* (19, 5, 0) {real, imag} */,
  {32'hbeaf9c5c, 32'h3fea5130} /* (19, 4, 31) {real, imag} */,
  {32'hc10c0128, 32'h40a27f7a} /* (19, 4, 30) {real, imag} */,
  {32'hc0aedc80, 32'hc0aeae64} /* (19, 4, 29) {real, imag} */,
  {32'h402a10d8, 32'hc0a93269} /* (19, 4, 28) {real, imag} */,
  {32'hc03535b4, 32'h3e253aa0} /* (19, 4, 27) {real, imag} */,
  {32'h3f7bf91c, 32'hbf454454} /* (19, 4, 26) {real, imag} */,
  {32'h3f8a2369, 32'hbead2a00} /* (19, 4, 25) {real, imag} */,
  {32'h3efe3244, 32'hc0a857b4} /* (19, 4, 24) {real, imag} */,
  {32'h4155dde3, 32'h4049dfa6} /* (19, 4, 23) {real, imag} */,
  {32'h40960780, 32'h40ced030} /* (19, 4, 22) {real, imag} */,
  {32'hc08bd31c, 32'h40ad8846} /* (19, 4, 21) {real, imag} */,
  {32'h3dcc6ba0, 32'h408b77b4} /* (19, 4, 20) {real, imag} */,
  {32'h40e3497f, 32'h4075f427} /* (19, 4, 19) {real, imag} */,
  {32'h40a51020, 32'h3e97eb18} /* (19, 4, 18) {real, imag} */,
  {32'h3f65f316, 32'hbff4c3a6} /* (19, 4, 17) {real, imag} */,
  {32'hbf2ab1b4, 32'hc0ae363a} /* (19, 4, 16) {real, imag} */,
  {32'hc0f5c81e, 32'hc1098202} /* (19, 4, 15) {real, imag} */,
  {32'hc121e5c6, 32'hc0d18566} /* (19, 4, 14) {real, imag} */,
  {32'hc1080610, 32'hc0ee1f1d} /* (19, 4, 13) {real, imag} */,
  {32'hc0b84182, 32'hbf9d0e9c} /* (19, 4, 12) {real, imag} */,
  {32'hc144d323, 32'hbeef5038} /* (19, 4, 11) {real, imag} */,
  {32'hc11372ae, 32'hc061a0d6} /* (19, 4, 10) {real, imag} */,
  {32'hc071aec1, 32'hc01bea66} /* (19, 4, 9) {real, imag} */,
  {32'h3f66e3f6, 32'h40895e3a} /* (19, 4, 8) {real, imag} */,
  {32'hbfb9f0f5, 32'hbfb13c3e} /* (19, 4, 7) {real, imag} */,
  {32'hc0238434, 32'h40101154} /* (19, 4, 6) {real, imag} */,
  {32'hc03a1420, 32'h40f8e60c} /* (19, 4, 5) {real, imag} */,
  {32'h3ff02331, 32'h3eabbca0} /* (19, 4, 4) {real, imag} */,
  {32'h3f7a751c, 32'h403ab8e0} /* (19, 4, 3) {real, imag} */,
  {32'h3e75a008, 32'h408442c0} /* (19, 4, 2) {real, imag} */,
  {32'hc02c5de3, 32'hbfe1f408} /* (19, 4, 1) {real, imag} */,
  {32'hc04df8b8, 32'h4029ed10} /* (19, 4, 0) {real, imag} */,
  {32'hbf77996d, 32'hc0ab951c} /* (19, 3, 31) {real, imag} */,
  {32'h400f4968, 32'hc0240982} /* (19, 3, 30) {real, imag} */,
  {32'h4042e056, 32'h40600fcd} /* (19, 3, 29) {real, imag} */,
  {32'h40c8f3b2, 32'h3fda9801} /* (19, 3, 28) {real, imag} */,
  {32'h40b28fc6, 32'h3f2bbea0} /* (19, 3, 27) {real, imag} */,
  {32'hc04131ba, 32'hc093f5fb} /* (19, 3, 26) {real, imag} */,
  {32'hc0c3045e, 32'hc0a38f9a} /* (19, 3, 25) {real, imag} */,
  {32'hc00beb65, 32'hc1034628} /* (19, 3, 24) {real, imag} */,
  {32'h3f851ca8, 32'hc098f2f3} /* (19, 3, 23) {real, imag} */,
  {32'h40d68ad6, 32'hc04510e8} /* (19, 3, 22) {real, imag} */,
  {32'h40c46153, 32'hc096b0f4} /* (19, 3, 21) {real, imag} */,
  {32'hbf7877b0, 32'h3fb1de78} /* (19, 3, 20) {real, imag} */,
  {32'h400c462c, 32'hc0b9607e} /* (19, 3, 19) {real, imag} */,
  {32'hc0b48dea, 32'hbeea9a81} /* (19, 3, 18) {real, imag} */,
  {32'hbfcb1f61, 32'h412ae22a} /* (19, 3, 17) {real, imag} */,
  {32'h405f0767, 32'h4047e40d} /* (19, 3, 16) {real, imag} */,
  {32'hbe948742, 32'h4037342e} /* (19, 3, 15) {real, imag} */,
  {32'hc052864d, 32'h40b177bf} /* (19, 3, 14) {real, imag} */,
  {32'hc0c668cc, 32'h4108d4e4} /* (19, 3, 13) {real, imag} */,
  {32'hc09c98c5, 32'h40d74eea} /* (19, 3, 12) {real, imag} */,
  {32'h3e71c318, 32'hc0963610} /* (19, 3, 11) {real, imag} */,
  {32'h3f76b4a6, 32'hc0a3eee8} /* (19, 3, 10) {real, imag} */,
  {32'hc0ddfd21, 32'hc00ed650} /* (19, 3, 9) {real, imag} */,
  {32'hbfbb5f44, 32'h3f18b84d} /* (19, 3, 8) {real, imag} */,
  {32'h40dcdbc7, 32'h406c28af} /* (19, 3, 7) {real, imag} */,
  {32'h409dc2e1, 32'hbfab05cf} /* (19, 3, 6) {real, imag} */,
  {32'h41069504, 32'hbfe91ba5} /* (19, 3, 5) {real, imag} */,
  {32'h401c93ba, 32'hc085d30b} /* (19, 3, 4) {real, imag} */,
  {32'hc04caa7e, 32'hc07d3036} /* (19, 3, 3) {real, imag} */,
  {32'hc0d47464, 32'hc1181540} /* (19, 3, 2) {real, imag} */,
  {32'h400cfe4f, 32'h40120329} /* (19, 3, 1) {real, imag} */,
  {32'hbe302f40, 32'hbe168ad8} /* (19, 3, 0) {real, imag} */,
  {32'hc00a3b9d, 32'h3f57ae18} /* (19, 2, 31) {real, imag} */,
  {32'h3dfdf040, 32'h3f324ed8} /* (19, 2, 30) {real, imag} */,
  {32'h40604908, 32'h40934bc1} /* (19, 2, 29) {real, imag} */,
  {32'hbed70600, 32'h41337a88} /* (19, 2, 28) {real, imag} */,
  {32'hc10e546c, 32'h411ff81f} /* (19, 2, 27) {real, imag} */,
  {32'hc12cbfb6, 32'hbfad727c} /* (19, 2, 26) {real, imag} */,
  {32'hc0c8343a, 32'hc0a2561a} /* (19, 2, 25) {real, imag} */,
  {32'h3f0a3cd8, 32'hc08977d6} /* (19, 2, 24) {real, imag} */,
  {32'h40ba0143, 32'h4080bfc0} /* (19, 2, 23) {real, imag} */,
  {32'hbfccc534, 32'h40342708} /* (19, 2, 22) {real, imag} */,
  {32'hbf1a0020, 32'hc0ee5047} /* (19, 2, 21) {real, imag} */,
  {32'h40a20754, 32'hc0711288} /* (19, 2, 20) {real, imag} */,
  {32'h40e311f7, 32'h40d8983e} /* (19, 2, 19) {real, imag} */,
  {32'h3f95afda, 32'h408fdb47} /* (19, 2, 18) {real, imag} */,
  {32'h407c237c, 32'h3f744408} /* (19, 2, 17) {real, imag} */,
  {32'h3fd10fd7, 32'hc0715777} /* (19, 2, 16) {real, imag} */,
  {32'hc088dba5, 32'hbb929800} /* (19, 2, 15) {real, imag} */,
  {32'hc0811730, 32'h3fc81ea8} /* (19, 2, 14) {real, imag} */,
  {32'hbf55adbc, 32'hc02820ff} /* (19, 2, 13) {real, imag} */,
  {32'hc0c703fe, 32'hc113d670} /* (19, 2, 12) {real, imag} */,
  {32'hc0c89d86, 32'hc02e1c64} /* (19, 2, 11) {real, imag} */,
  {32'hc0f7b93f, 32'hc07f2266} /* (19, 2, 10) {real, imag} */,
  {32'hc0d08d34, 32'h3cc94c00} /* (19, 2, 9) {real, imag} */,
  {32'hc01b9c04, 32'h402fc0d6} /* (19, 2, 8) {real, imag} */,
  {32'h3fd02073, 32'hc03546c0} /* (19, 2, 7) {real, imag} */,
  {32'h40a363ee, 32'hbf92f718} /* (19, 2, 6) {real, imag} */,
  {32'hc04c64fe, 32'h3fe4f070} /* (19, 2, 5) {real, imag} */,
  {32'hbfd8fbea, 32'hbe6b2c00} /* (19, 2, 4) {real, imag} */,
  {32'h40ebe116, 32'h40089db1} /* (19, 2, 3) {real, imag} */,
  {32'hc019d470, 32'h40abfd64} /* (19, 2, 2) {real, imag} */,
  {32'hc092f4e9, 32'h40e04e82} /* (19, 2, 1) {real, imag} */,
  {32'hbfadd526, 32'hbf0dde56} /* (19, 2, 0) {real, imag} */,
  {32'hbf176ac4, 32'h4072520e} /* (19, 1, 31) {real, imag} */,
  {32'hbf25a48a, 32'hbcfbb300} /* (19, 1, 30) {real, imag} */,
  {32'hc0516d6d, 32'hc05a04e0} /* (19, 1, 29) {real, imag} */,
  {32'h40dad0aa, 32'hbfca4808} /* (19, 1, 28) {real, imag} */,
  {32'h410994b5, 32'h40b2ee0b} /* (19, 1, 27) {real, imag} */,
  {32'hc00ea19e, 32'h410b8030} /* (19, 1, 26) {real, imag} */,
  {32'hbcf2b1f8, 32'h40bc499a} /* (19, 1, 25) {real, imag} */,
  {32'h40620e3e, 32'h408bce5b} /* (19, 1, 24) {real, imag} */,
  {32'hc04b1d8c, 32'hc0723d7d} /* (19, 1, 23) {real, imag} */,
  {32'hbf495548, 32'hc0eb7690} /* (19, 1, 22) {real, imag} */,
  {32'h4033187d, 32'hc089ba98} /* (19, 1, 21) {real, imag} */,
  {32'hbfd57a97, 32'hc0c763c2} /* (19, 1, 20) {real, imag} */,
  {32'hc003b446, 32'hc0bdcb34} /* (19, 1, 19) {real, imag} */,
  {32'hbfe282c4, 32'hc038029c} /* (19, 1, 18) {real, imag} */,
  {32'h3fe99e75, 32'h4013381a} /* (19, 1, 17) {real, imag} */,
  {32'h41359446, 32'h40c51f09} /* (19, 1, 16) {real, imag} */,
  {32'h40f4b71b, 32'hc029a1af} /* (19, 1, 15) {real, imag} */,
  {32'hc0768df9, 32'hc0c5890a} /* (19, 1, 14) {real, imag} */,
  {32'hbf111ea8, 32'hbb234a00} /* (19, 1, 13) {real, imag} */,
  {32'hc057ee1a, 32'h4031485b} /* (19, 1, 12) {real, imag} */,
  {32'hc0ae13a7, 32'h3f2e38e8} /* (19, 1, 11) {real, imag} */,
  {32'hc0ba92d0, 32'h3fd2f52c} /* (19, 1, 10) {real, imag} */,
  {32'h40380b4e, 32'hc06d2ac5} /* (19, 1, 9) {real, imag} */,
  {32'h3eb4af20, 32'hc10af86e} /* (19, 1, 8) {real, imag} */,
  {32'h406e534c, 32'hc091ffa8} /* (19, 1, 7) {real, imag} */,
  {32'h40de93d6, 32'h3d9e41d8} /* (19, 1, 6) {real, imag} */,
  {32'hc103c5e4, 32'h409853aa} /* (19, 1, 5) {real, imag} */,
  {32'hc08db177, 32'h400b76fa} /* (19, 1, 4) {real, imag} */,
  {32'h40aaa424, 32'hc0f3589e} /* (19, 1, 3) {real, imag} */,
  {32'h4095276c, 32'hc0016a14} /* (19, 1, 2) {real, imag} */,
  {32'h3fb167d8, 32'h3fb2b196} /* (19, 1, 1) {real, imag} */,
  {32'hbe5a4dd0, 32'h405d1bdb} /* (19, 1, 0) {real, imag} */,
  {32'hc09e4128, 32'h40cf58e6} /* (19, 0, 31) {real, imag} */,
  {32'hbe887e00, 32'h40a691dc} /* (19, 0, 30) {real, imag} */,
  {32'hbecaa8d0, 32'h3fe3e361} /* (19, 0, 29) {real, imag} */,
  {32'hc11d4e58, 32'hc0c05be1} /* (19, 0, 28) {real, imag} */,
  {32'hc11d9b88, 32'hbfe6dee7} /* (19, 0, 27) {real, imag} */,
  {32'hbff86b1a, 32'h403fd4b0} /* (19, 0, 26) {real, imag} */,
  {32'hc01da2a1, 32'hc0324241} /* (19, 0, 25) {real, imag} */,
  {32'hc0d89aee, 32'h3d6967a8} /* (19, 0, 24) {real, imag} */,
  {32'hc05e5a2e, 32'h40488ef0} /* (19, 0, 23) {real, imag} */,
  {32'hc0c389c1, 32'h40f8b2d6} /* (19, 0, 22) {real, imag} */,
  {32'h400662a6, 32'h4118bc0e} /* (19, 0, 21) {real, imag} */,
  {32'h3f9f7c36, 32'hbe5bd85c} /* (19, 0, 20) {real, imag} */,
  {32'h3e90fc98, 32'h40035de2} /* (19, 0, 19) {real, imag} */,
  {32'h4105d498, 32'h403b9b78} /* (19, 0, 18) {real, imag} */,
  {32'h413a31f2, 32'hc03bc680} /* (19, 0, 17) {real, imag} */,
  {32'hc0bd980c, 32'hc0fc5d55} /* (19, 0, 16) {real, imag} */,
  {32'hc06501cb, 32'hc08a2b61} /* (19, 0, 15) {real, imag} */,
  {32'h3fff5a7a, 32'hc10dc0ac} /* (19, 0, 14) {real, imag} */,
  {32'hc0934bd4, 32'hc0ce076f} /* (19, 0, 13) {real, imag} */,
  {32'hc09acd00, 32'hbf8769d6} /* (19, 0, 12) {real, imag} */,
  {32'h40b391da, 32'h40520db9} /* (19, 0, 11) {real, imag} */,
  {32'h4007840a, 32'hc00be104} /* (19, 0, 10) {real, imag} */,
  {32'h40bf0561, 32'hc05928a8} /* (19, 0, 9) {real, imag} */,
  {32'h40f01f80, 32'hc09a1d42} /* (19, 0, 8) {real, imag} */,
  {32'h40133564, 32'h4026b122} /* (19, 0, 7) {real, imag} */,
  {32'hc092b6a2, 32'hbf9b03c6} /* (19, 0, 6) {real, imag} */,
  {32'hc0b604be, 32'hbf06dc98} /* (19, 0, 5) {real, imag} */,
  {32'hbeb95cdc, 32'hbf984e6e} /* (19, 0, 4) {real, imag} */,
  {32'h40f15d34, 32'hc05c8cb0} /* (19, 0, 3) {real, imag} */,
  {32'h4104df0f, 32'h3e12b62c} /* (19, 0, 2) {real, imag} */,
  {32'h40c66c98, 32'h40e2bd79} /* (19, 0, 1) {real, imag} */,
  {32'hc0066aee, 32'h40a67c9d} /* (19, 0, 0) {real, imag} */,
  {32'hc0b3601c, 32'h3f696da2} /* (18, 31, 31) {real, imag} */,
  {32'hc0c94b0d, 32'hc001fa7d} /* (18, 31, 30) {real, imag} */,
  {32'hc0598e36, 32'hc0e327c8} /* (18, 31, 29) {real, imag} */,
  {32'hc12fe276, 32'hbe4257c2} /* (18, 31, 28) {real, imag} */,
  {32'hc18d1c5d, 32'h401ab752} /* (18, 31, 27) {real, imag} */,
  {32'hc1a2600e, 32'h3f93c39d} /* (18, 31, 26) {real, imag} */,
  {32'hc1817dfa, 32'hc099b7b7} /* (18, 31, 25) {real, imag} */,
  {32'hc1801e80, 32'hbfb42360} /* (18, 31, 24) {real, imag} */,
  {32'hc15fd288, 32'hc0cdb9f2} /* (18, 31, 23) {real, imag} */,
  {32'hc0d30420, 32'hc0530c56} /* (18, 31, 22) {real, imag} */,
  {32'hc091ee1e, 32'h40195303} /* (18, 31, 21) {real, imag} */,
  {32'hc00d5511, 32'hbfa645ba} /* (18, 31, 20) {real, imag} */,
  {32'h3fe22709, 32'hbf687440} /* (18, 31, 19) {real, imag} */,
  {32'h415adfaf, 32'hc0399064} /* (18, 31, 18) {real, imag} */,
  {32'h41269a1e, 32'hbfdccea4} /* (18, 31, 17) {real, imag} */,
  {32'h402b0054, 32'hc08a4bf4} /* (18, 31, 16) {real, imag} */,
  {32'h411ead88, 32'h405ec9d8} /* (18, 31, 15) {real, imag} */,
  {32'h416d53ea, 32'h403b4c08} /* (18, 31, 14) {real, imag} */,
  {32'h41669841, 32'h401b7e19} /* (18, 31, 13) {real, imag} */,
  {32'h411804aa, 32'h40027f7b} /* (18, 31, 12) {real, imag} */,
  {32'h4025a5ef, 32'h40941798} /* (18, 31, 11) {real, imag} */,
  {32'h4038d1b6, 32'hbd4cb000} /* (18, 31, 10) {real, imag} */,
  {32'hc098c32a, 32'hc09fdb39} /* (18, 31, 9) {real, imag} */,
  {32'hc142c806, 32'hbf139252} /* (18, 31, 8) {real, imag} */,
  {32'hc0a9603d, 32'h408d13ef} /* (18, 31, 7) {real, imag} */,
  {32'h4041c6ec, 32'h3f8f16de} /* (18, 31, 6) {real, imag} */,
  {32'hc02ef038, 32'hbffa186f} /* (18, 31, 5) {real, imag} */,
  {32'hc10d7ffc, 32'hc0a45e8b} /* (18, 31, 4) {real, imag} */,
  {32'hc12c9e2a, 32'hbf5927ec} /* (18, 31, 3) {real, imag} */,
  {32'hc15eafb2, 32'h409da974} /* (18, 31, 2) {real, imag} */,
  {32'hc1269a66, 32'h3f7fa218} /* (18, 31, 1) {real, imag} */,
  {32'hc0a6187f, 32'h402d0645} /* (18, 31, 0) {real, imag} */,
  {32'h40b0c715, 32'hbfdbae5c} /* (18, 30, 31) {real, imag} */,
  {32'h407c8e06, 32'h3ef51f14} /* (18, 30, 30) {real, imag} */,
  {32'h40a83586, 32'hc0ceda3d} /* (18, 30, 29) {real, imag} */,
  {32'h40dc5ba6, 32'hc090847d} /* (18, 30, 28) {real, imag} */,
  {32'h41005c59, 32'h4047de86} /* (18, 30, 27) {real, imag} */,
  {32'h410d2473, 32'h402e0d70} /* (18, 30, 26) {real, imag} */,
  {32'h40bb2694, 32'hc0081844} /* (18, 30, 25) {real, imag} */,
  {32'h40233bef, 32'hc0500ee7} /* (18, 30, 24) {real, imag} */,
  {32'hc046f16e, 32'h40a09ba8} /* (18, 30, 23) {real, imag} */,
  {32'h40a62172, 32'hc00a0dfc} /* (18, 30, 22) {real, imag} */,
  {32'h41148b3d, 32'hc0fa58c2} /* (18, 30, 21) {real, imag} */,
  {32'h3f19ce68, 32'hc112b4b2} /* (18, 30, 20) {real, imag} */,
  {32'hc0a47e7e, 32'hc10f7bdc} /* (18, 30, 19) {real, imag} */,
  {32'hc0e85362, 32'hc0add564} /* (18, 30, 18) {real, imag} */,
  {32'hc0d93291, 32'hbf8b3a9c} /* (18, 30, 17) {real, imag} */,
  {32'hc1478caf, 32'hc02a2e14} /* (18, 30, 16) {real, imag} */,
  {32'hc0f05bce, 32'hc10e35a8} /* (18, 30, 15) {real, imag} */,
  {32'hc0ef5d28, 32'h408db7ed} /* (18, 30, 14) {real, imag} */,
  {32'hc0d2bb22, 32'h4071903c} /* (18, 30, 13) {real, imag} */,
  {32'hc0212492, 32'h40acea64} /* (18, 30, 12) {real, imag} */,
  {32'hc0cf3457, 32'h415850be} /* (18, 30, 11) {real, imag} */,
  {32'h3fe88804, 32'h41086042} /* (18, 30, 10) {real, imag} */,
  {32'h4115ddf1, 32'h40bdb00f} /* (18, 30, 9) {real, imag} */,
  {32'h4130d0ac, 32'h408d8c50} /* (18, 30, 8) {real, imag} */,
  {32'h41762692, 32'h40b70ff6} /* (18, 30, 7) {real, imag} */,
  {32'h417041cb, 32'h408c732e} /* (18, 30, 6) {real, imag} */,
  {32'h40b1a212, 32'h3ed132ae} /* (18, 30, 5) {real, imag} */,
  {32'h407bf323, 32'hc00919c8} /* (18, 30, 4) {real, imag} */,
  {32'hc07f4554, 32'hc02d2af1} /* (18, 30, 3) {real, imag} */,
  {32'h401c1bc7, 32'hc069a341} /* (18, 30, 2) {real, imag} */,
  {32'h412260b3, 32'hc0f2067e} /* (18, 30, 1) {real, imag} */,
  {32'h41251e35, 32'hc0cc060f} /* (18, 30, 0) {real, imag} */,
  {32'h3f9ce910, 32'h40a39362} /* (18, 29, 31) {real, imag} */,
  {32'hc0670ac4, 32'h40cf841c} /* (18, 29, 30) {real, imag} */,
  {32'hbfbf7fcb, 32'h40645074} /* (18, 29, 29) {real, imag} */,
  {32'h3f96c046, 32'hc090ebbc} /* (18, 29, 28) {real, imag} */,
  {32'hbdbeb960, 32'hc09004ff} /* (18, 29, 27) {real, imag} */,
  {32'h409b0902, 32'hc01d8ea5} /* (18, 29, 26) {real, imag} */,
  {32'h409ccc24, 32'h3e893e38} /* (18, 29, 25) {real, imag} */,
  {32'h4106ec55, 32'hc0789ceb} /* (18, 29, 24) {real, imag} */,
  {32'h3ff6b100, 32'hc05cbae3} /* (18, 29, 23) {real, imag} */,
  {32'hc0e5af46, 32'hc03e4036} /* (18, 29, 22) {real, imag} */,
  {32'hc0a082d0, 32'hbf724dcc} /* (18, 29, 21) {real, imag} */,
  {32'h3f324cae, 32'hc01dfd7d} /* (18, 29, 20) {real, imag} */,
  {32'h3dd3b610, 32'h3e97afaa} /* (18, 29, 19) {real, imag} */,
  {32'hc0366eb2, 32'hbf30e448} /* (18, 29, 18) {real, imag} */,
  {32'h4006cd2e, 32'hc018fb8a} /* (18, 29, 17) {real, imag} */,
  {32'h3fa19318, 32'hbfa27649} /* (18, 29, 16) {real, imag} */,
  {32'h4080f6cd, 32'hbe6cfd10} /* (18, 29, 15) {real, imag} */,
  {32'h40a5e661, 32'hc080f006} /* (18, 29, 14) {real, imag} */,
  {32'hbfb1d904, 32'hc072954f} /* (18, 29, 13) {real, imag} */,
  {32'hc02365f2, 32'h3f529874} /* (18, 29, 12) {real, imag} */,
  {32'hc06474a5, 32'hbfe02978} /* (18, 29, 11) {real, imag} */,
  {32'h3ef1c37e, 32'hc016f2d4} /* (18, 29, 10) {real, imag} */,
  {32'hc0cc9615, 32'hbbe97800} /* (18, 29, 9) {real, imag} */,
  {32'hc06d4017, 32'h40d80a53} /* (18, 29, 8) {real, imag} */,
  {32'hbf4aecb0, 32'h40f8a827} /* (18, 29, 7) {real, imag} */,
  {32'h40040f78, 32'h41356360} /* (18, 29, 6) {real, imag} */,
  {32'h4091aca5, 32'h4083ed09} /* (18, 29, 5) {real, imag} */,
  {32'h40b10676, 32'h405c7c8e} /* (18, 29, 4) {real, imag} */,
  {32'h3d981600, 32'hbfda34eb} /* (18, 29, 3) {real, imag} */,
  {32'h4032615c, 32'hc08326fe} /* (18, 29, 2) {real, imag} */,
  {32'h40622b7f, 32'h401d36cd} /* (18, 29, 1) {real, imag} */,
  {32'h407e649e, 32'h4082c871} /* (18, 29, 0) {real, imag} */,
  {32'h3f38dc86, 32'h404e5c66} /* (18, 28, 31) {real, imag} */,
  {32'h3fbdbeee, 32'h3fdee68e} /* (18, 28, 30) {real, imag} */,
  {32'hbfc435ac, 32'hbf839b68} /* (18, 28, 29) {real, imag} */,
  {32'h3f83d89c, 32'hbfd1429e} /* (18, 28, 28) {real, imag} */,
  {32'h3ff4b570, 32'hc09d4a87} /* (18, 28, 27) {real, imag} */,
  {32'h400c4b6d, 32'hc027d2c4} /* (18, 28, 26) {real, imag} */,
  {32'h3f6c07d2, 32'hbe90834c} /* (18, 28, 25) {real, imag} */,
  {32'h3e8d5b6f, 32'h3fb4a779} /* (18, 28, 24) {real, imag} */,
  {32'h3fa75af6, 32'hbfb55dc9} /* (18, 28, 23) {real, imag} */,
  {32'h403b8726, 32'hc06038df} /* (18, 28, 22) {real, imag} */,
  {32'h40a52022, 32'hbed1202e} /* (18, 28, 21) {real, imag} */,
  {32'h409c3348, 32'hbee33ec8} /* (18, 28, 20) {real, imag} */,
  {32'h410fa0b8, 32'h4019f89e} /* (18, 28, 19) {real, imag} */,
  {32'h40cb8cd3, 32'h401bdb16} /* (18, 28, 18) {real, imag} */,
  {32'h40c324a6, 32'hbe7510c0} /* (18, 28, 17) {real, imag} */,
  {32'h41009572, 32'hc0556398} /* (18, 28, 16) {real, imag} */,
  {32'h3fb7ca18, 32'hbec29630} /* (18, 28, 15) {real, imag} */,
  {32'h3f264fcc, 32'h3e1a9330} /* (18, 28, 14) {real, imag} */,
  {32'h40b270f7, 32'h3e8e9a04} /* (18, 28, 13) {real, imag} */,
  {32'h401647bd, 32'h41094db6} /* (18, 28, 12) {real, imag} */,
  {32'h3fe13ee4, 32'h409d6b9d} /* (18, 28, 11) {real, imag} */,
  {32'h3f4732a4, 32'hbf8eee19} /* (18, 28, 10) {real, imag} */,
  {32'hc008da6e, 32'h3fcce011} /* (18, 28, 9) {real, imag} */,
  {32'hbf7ac154, 32'hbe768030} /* (18, 28, 8) {real, imag} */,
  {32'hc00952c4, 32'hbefeec10} /* (18, 28, 7) {real, imag} */,
  {32'hc10552eb, 32'h40da1211} /* (18, 28, 6) {real, imag} */,
  {32'hc1254aee, 32'h3fde359d} /* (18, 28, 5) {real, imag} */,
  {32'hc0ef151f, 32'h3fbe2632} /* (18, 28, 4) {real, imag} */,
  {32'hc0d5112c, 32'hbf938344} /* (18, 28, 3) {real, imag} */,
  {32'hc10d1a2a, 32'hbeeb4560} /* (18, 28, 2) {real, imag} */,
  {32'hc0900d80, 32'h40f79f52} /* (18, 28, 1) {real, imag} */,
  {32'hbf0f75c9, 32'h405ae599} /* (18, 28, 0) {real, imag} */,
  {32'h40342a64, 32'hbf14cdcb} /* (18, 27, 31) {real, imag} */,
  {32'h408ddf0c, 32'hc0a425e5} /* (18, 27, 30) {real, imag} */,
  {32'h40744f66, 32'h400cedbf} /* (18, 27, 29) {real, imag} */,
  {32'h402999d3, 32'hc013135d} /* (18, 27, 28) {real, imag} */,
  {32'h40476351, 32'hc1038c0f} /* (18, 27, 27) {real, imag} */,
  {32'h4098e413, 32'hc0c4024d} /* (18, 27, 26) {real, imag} */,
  {32'h411b7e48, 32'hbffe98ac} /* (18, 27, 25) {real, imag} */,
  {32'h4104ff61, 32'hc092e242} /* (18, 27, 24) {real, imag} */,
  {32'h40ea1f18, 32'hc02054fc} /* (18, 27, 23) {real, imag} */,
  {32'h41183954, 32'hc0200234} /* (18, 27, 22) {real, imag} */,
  {32'h40319eee, 32'hc0ce241b} /* (18, 27, 21) {real, imag} */,
  {32'hc0137799, 32'hc08fa540} /* (18, 27, 20) {real, imag} */,
  {32'hc00d4dc4, 32'h401a0524} /* (18, 27, 19) {real, imag} */,
  {32'h40c0df27, 32'h41112aa8} /* (18, 27, 18) {real, imag} */,
  {32'h3fbe22ca, 32'h4048390b} /* (18, 27, 17) {real, imag} */,
  {32'h3fe5ae4d, 32'hc09e68d2} /* (18, 27, 16) {real, imag} */,
  {32'h40c22e78, 32'hbe913720} /* (18, 27, 15) {real, imag} */,
  {32'h40f901c6, 32'hbde83440} /* (18, 27, 14) {real, imag} */,
  {32'h3ff83b11, 32'hc007e57e} /* (18, 27, 13) {real, imag} */,
  {32'h40305809, 32'hc09f2197} /* (18, 27, 12) {real, imag} */,
  {32'hbf8fa6ec, 32'h3f83930c} /* (18, 27, 11) {real, imag} */,
  {32'hbf53a120, 32'h3fdc86e2} /* (18, 27, 10) {real, imag} */,
  {32'hc0301a2c, 32'hc0b9efa1} /* (18, 27, 9) {real, imag} */,
  {32'h4002e26d, 32'hc10b91ea} /* (18, 27, 8) {real, imag} */,
  {32'hbf586fd0, 32'hc0f49a22} /* (18, 27, 7) {real, imag} */,
  {32'hbf58caac, 32'hc0909580} /* (18, 27, 6) {real, imag} */,
  {32'h3ff33d44, 32'hc06e79c6} /* (18, 27, 5) {real, imag} */,
  {32'hbfba6ae0, 32'hbfbd0b2e} /* (18, 27, 4) {real, imag} */,
  {32'hc034440b, 32'hbfcdebb2} /* (18, 27, 3) {real, imag} */,
  {32'hbfdf6526, 32'hc00f125c} /* (18, 27, 2) {real, imag} */,
  {32'h400a0102, 32'hc0c319ba} /* (18, 27, 1) {real, imag} */,
  {32'h4020bfc8, 32'hc0c01c40} /* (18, 27, 0) {real, imag} */,
  {32'h407c03c5, 32'hbff95b5b} /* (18, 26, 31) {real, imag} */,
  {32'h3f97701d, 32'h4007747e} /* (18, 26, 30) {real, imag} */,
  {32'hbf325694, 32'h3fe74e10} /* (18, 26, 29) {real, imag} */,
  {32'h3ef07826, 32'h3fe39046} /* (18, 26, 28) {real, imag} */,
  {32'h406927e6, 32'h3fba839a} /* (18, 26, 27) {real, imag} */,
  {32'h400b2e9a, 32'hbfd16ecf} /* (18, 26, 26) {real, imag} */,
  {32'hbf20c8a5, 32'hc0497c37} /* (18, 26, 25) {real, imag} */,
  {32'hc0964a50, 32'hc0265852} /* (18, 26, 24) {real, imag} */,
  {32'hc0deceb1, 32'h4016c714} /* (18, 26, 23) {real, imag} */,
  {32'hc01eba0d, 32'h409986be} /* (18, 26, 22) {real, imag} */,
  {32'h3ffbe7f4, 32'hbf19dda8} /* (18, 26, 21) {real, imag} */,
  {32'hbfa08c19, 32'h3e445140} /* (18, 26, 20) {real, imag} */,
  {32'h403b6b0c, 32'h40b2ccaa} /* (18, 26, 19) {real, imag} */,
  {32'h3f76faae, 32'h406988b1} /* (18, 26, 18) {real, imag} */,
  {32'h40867710, 32'hbfcec8d7} /* (18, 26, 17) {real, imag} */,
  {32'h4091c794, 32'h3f9e9531} /* (18, 26, 16) {real, imag} */,
  {32'h40a86510, 32'hc01c0bd7} /* (18, 26, 15) {real, imag} */,
  {32'hbe6c5f60, 32'hc09afb68} /* (18, 26, 14) {real, imag} */,
  {32'hbfbc16de, 32'hc03e1ec0} /* (18, 26, 13) {real, imag} */,
  {32'hc02cc9bc, 32'hbf1e53ee} /* (18, 26, 12) {real, imag} */,
  {32'hc06cd8df, 32'hc088855d} /* (18, 26, 11) {real, imag} */,
  {32'h4049c51f, 32'hbfe683cc} /* (18, 26, 10) {real, imag} */,
  {32'h40ef7d2c, 32'h41071950} /* (18, 26, 9) {real, imag} */,
  {32'h40b81260, 32'h411e46e9} /* (18, 26, 8) {real, imag} */,
  {32'h3ff19671, 32'h40303ac6} /* (18, 26, 7) {real, imag} */,
  {32'h4044b0c8, 32'h3fb971a4} /* (18, 26, 6) {real, imag} */,
  {32'h4084acd8, 32'h401b924e} /* (18, 26, 5) {real, imag} */,
  {32'h3e5a1dec, 32'h40490f6b} /* (18, 26, 4) {real, imag} */,
  {32'h3f517eaa, 32'hbfba9ef6} /* (18, 26, 3) {real, imag} */,
  {32'h40b0c5f0, 32'hc028b648} /* (18, 26, 2) {real, imag} */,
  {32'h405d76a9, 32'h4008409d} /* (18, 26, 1) {real, imag} */,
  {32'h40274eba, 32'hbf242069} /* (18, 26, 0) {real, imag} */,
  {32'h401eb7be, 32'hbe4c0460} /* (18, 25, 31) {real, imag} */,
  {32'h400e73b7, 32'h40392b28} /* (18, 25, 30) {real, imag} */,
  {32'h3f4ec283, 32'h40c53a6f} /* (18, 25, 29) {real, imag} */,
  {32'hbfa905c7, 32'h4082ddb8} /* (18, 25, 28) {real, imag} */,
  {32'hc0dc1a90, 32'hbfd3ff7c} /* (18, 25, 27) {real, imag} */,
  {32'hc08f02e0, 32'hbd86f820} /* (18, 25, 26) {real, imag} */,
  {32'hbfdefcd7, 32'h3f38dd78} /* (18, 25, 25) {real, imag} */,
  {32'hbe484724, 32'h3fe07422} /* (18, 25, 24) {real, imag} */,
  {32'h3faa16dd, 32'hc03b4a64} /* (18, 25, 23) {real, imag} */,
  {32'h40a425aa, 32'hc0de84fe} /* (18, 25, 22) {real, imag} */,
  {32'h4010d0d2, 32'hc0d090ca} /* (18, 25, 21) {real, imag} */,
  {32'hc03cd8a8, 32'hc0bdb604} /* (18, 25, 20) {real, imag} */,
  {32'hc0c66d10, 32'hc08765de} /* (18, 25, 19) {real, imag} */,
  {32'hc0e9cb5a, 32'hbff8262a} /* (18, 25, 18) {real, imag} */,
  {32'hc054ac42, 32'h3fb03cee} /* (18, 25, 17) {real, imag} */,
  {32'h4002b668, 32'hbcb724a0} /* (18, 25, 16) {real, imag} */,
  {32'h40c2fe8e, 32'hbf1ff238} /* (18, 25, 15) {real, imag} */,
  {32'hbe257cb8, 32'hbffa3633} /* (18, 25, 14) {real, imag} */,
  {32'h4008ae27, 32'hbe51622c} /* (18, 25, 13) {real, imag} */,
  {32'h40861de4, 32'h4105986f} /* (18, 25, 12) {real, imag} */,
  {32'hbfe462a2, 32'h3fe6be7d} /* (18, 25, 11) {real, imag} */,
  {32'hbf81dba2, 32'hbe662a00} /* (18, 25, 10) {real, imag} */,
  {32'h3e9d4610, 32'h40ec81b6} /* (18, 25, 9) {real, imag} */,
  {32'hbea8c738, 32'h40b2ea96} /* (18, 25, 8) {real, imag} */,
  {32'h40270af9, 32'hbfce825c} /* (18, 25, 7) {real, imag} */,
  {32'h406d3384, 32'hbf83ccc6} /* (18, 25, 6) {real, imag} */,
  {32'h3e1d3948, 32'h3f90f954} /* (18, 25, 5) {real, imag} */,
  {32'hc0fe9f76, 32'h40850be5} /* (18, 25, 4) {real, imag} */,
  {32'hc1090668, 32'h408c1cfb} /* (18, 25, 3) {real, imag} */,
  {32'hc050aea0, 32'hbee81758} /* (18, 25, 2) {real, imag} */,
  {32'hbf1407fe, 32'hc03bebf4} /* (18, 25, 1) {real, imag} */,
  {32'hbee5249c, 32'h3f3af724} /* (18, 25, 0) {real, imag} */,
  {32'h3fe4ac10, 32'hc0858935} /* (18, 24, 31) {real, imag} */,
  {32'h3f781532, 32'hc095ec15} /* (18, 24, 30) {real, imag} */,
  {32'hbe9261a8, 32'hbf16a1e0} /* (18, 24, 29) {real, imag} */,
  {32'h3f13d630, 32'h3f0fd080} /* (18, 24, 28) {real, imag} */,
  {32'h4030d910, 32'hc00cd6f1} /* (18, 24, 27) {real, imag} */,
  {32'h3d5adbc0, 32'hbf0b5ce4} /* (18, 24, 26) {real, imag} */,
  {32'hbf967eae, 32'hbe13e370} /* (18, 24, 25) {real, imag} */,
  {32'hc0861cc1, 32'hbd2445a0} /* (18, 24, 24) {real, imag} */,
  {32'hc04fcd7e, 32'hc02ea5a6} /* (18, 24, 23) {real, imag} */,
  {32'hbfe169ef, 32'h400eba58} /* (18, 24, 22) {real, imag} */,
  {32'hc03729b0, 32'h4066918e} /* (18, 24, 21) {real, imag} */,
  {32'hc09e1b8d, 32'hc06d467d} /* (18, 24, 20) {real, imag} */,
  {32'hbf04db9e, 32'h3fcfa5d8} /* (18, 24, 19) {real, imag} */,
  {32'h3fa49715, 32'h40439c70} /* (18, 24, 18) {real, imag} */,
  {32'hbf884cec, 32'hbdf86b70} /* (18, 24, 17) {real, imag} */,
  {32'hbfea1254, 32'hc0331a4e} /* (18, 24, 16) {real, imag} */,
  {32'hc0ad0d26, 32'hbff3dc42} /* (18, 24, 15) {real, imag} */,
  {32'hc08624b0, 32'h4008e937} /* (18, 24, 14) {real, imag} */,
  {32'h3f32ca72, 32'h405b5bf7} /* (18, 24, 13) {real, imag} */,
  {32'hbf4db74c, 32'h4058dc91} /* (18, 24, 12) {real, imag} */,
  {32'h3e92a54c, 32'h408b19fe} /* (18, 24, 11) {real, imag} */,
  {32'h3edb1fea, 32'h4033b20e} /* (18, 24, 10) {real, imag} */,
  {32'h4020851e, 32'h3f4e4190} /* (18, 24, 9) {real, imag} */,
  {32'h3f6280b4, 32'hc0086886} /* (18, 24, 8) {real, imag} */,
  {32'h3f2edb84, 32'hbdbc7d20} /* (18, 24, 7) {real, imag} */,
  {32'h3f192c00, 32'h403d937a} /* (18, 24, 6) {real, imag} */,
  {32'h4055bb93, 32'hc0416f8e} /* (18, 24, 5) {real, imag} */,
  {32'h40061ec1, 32'hc09b9b4c} /* (18, 24, 4) {real, imag} */,
  {32'h4018d911, 32'hc05ae00e} /* (18, 24, 3) {real, imag} */,
  {32'h40b0f4be, 32'hc0378d06} /* (18, 24, 2) {real, imag} */,
  {32'h406d34bb, 32'h406829e2} /* (18, 24, 1) {real, imag} */,
  {32'hbf63b8f4, 32'h403caa1e} /* (18, 24, 0) {real, imag} */,
  {32'h3dbc6bd8, 32'h3f82a0cd} /* (18, 23, 31) {real, imag} */,
  {32'hbc120480, 32'h401c37b0} /* (18, 23, 30) {real, imag} */,
  {32'h40518ea3, 32'h3fb20f1e} /* (18, 23, 29) {real, imag} */,
  {32'h409d14a1, 32'h3f890eb4} /* (18, 23, 28) {real, imag} */,
  {32'h3fdfbf28, 32'hc025c70a} /* (18, 23, 27) {real, imag} */,
  {32'h3f6445d4, 32'hc01a3cec} /* (18, 23, 26) {real, imag} */,
  {32'hc010f6b8, 32'hb9c75800} /* (18, 23, 25) {real, imag} */,
  {32'hc052c5a9, 32'hbfe316be} /* (18, 23, 24) {real, imag} */,
  {32'h3f12493a, 32'h401a03cc} /* (18, 23, 23) {real, imag} */,
  {32'h402863f4, 32'h401793d6} /* (18, 23, 22) {real, imag} */,
  {32'hbff275a1, 32'hc0a9775d} /* (18, 23, 21) {real, imag} */,
  {32'h3f9f2ef6, 32'hc0736b4a} /* (18, 23, 20) {real, imag} */,
  {32'h3c980280, 32'hbfc58ad7} /* (18, 23, 19) {real, imag} */,
  {32'hc02590a5, 32'h3f90ee96} /* (18, 23, 18) {real, imag} */,
  {32'hc09f4b9d, 32'h40266000} /* (18, 23, 17) {real, imag} */,
  {32'h3fcf2ad2, 32'h3fa98a9e} /* (18, 23, 16) {real, imag} */,
  {32'h402b12b6, 32'h3f97c022} /* (18, 23, 15) {real, imag} */,
  {32'h4056a0d4, 32'hbfdeee8d} /* (18, 23, 14) {real, imag} */,
  {32'h40511c5c, 32'hbd331ec0} /* (18, 23, 13) {real, imag} */,
  {32'h3f8ae374, 32'h3f075130} /* (18, 23, 12) {real, imag} */,
  {32'h3e6b2230, 32'hbee0ce28} /* (18, 23, 11) {real, imag} */,
  {32'hbf8d230d, 32'h3ee0560a} /* (18, 23, 10) {real, imag} */,
  {32'hc026709b, 32'hc04b1176} /* (18, 23, 9) {real, imag} */,
  {32'hc07604a8, 32'hbe9cc534} /* (18, 23, 8) {real, imag} */,
  {32'hbf71c594, 32'h402a7328} /* (18, 23, 7) {real, imag} */,
  {32'h3fb90b02, 32'h409c6e22} /* (18, 23, 6) {real, imag} */,
  {32'h403f56d2, 32'h40b94680} /* (18, 23, 5) {real, imag} */,
  {32'h40aa60cd, 32'h40d0da6f} /* (18, 23, 4) {real, imag} */,
  {32'h4078e968, 32'h3f6b85e9} /* (18, 23, 3) {real, imag} */,
  {32'h3f56173a, 32'h3f22af54} /* (18, 23, 2) {real, imag} */,
  {32'hc02c909c, 32'h3f530ce4} /* (18, 23, 1) {real, imag} */,
  {32'hbff6783c, 32'h3f9568bf} /* (18, 23, 0) {real, imag} */,
  {32'h3ed9f570, 32'hbff2d621} /* (18, 22, 31) {real, imag} */,
  {32'hc06487f6, 32'hc023a698} /* (18, 22, 30) {real, imag} */,
  {32'hbf8c9c6a, 32'hbfe8b24a} /* (18, 22, 29) {real, imag} */,
  {32'h3fd98dca, 32'hbf39d638} /* (18, 22, 28) {real, imag} */,
  {32'h4093c5ac, 32'hc03120da} /* (18, 22, 27) {real, imag} */,
  {32'h404fb063, 32'hc06b789c} /* (18, 22, 26) {real, imag} */,
  {32'h401ab55d, 32'h3f2b12f3} /* (18, 22, 25) {real, imag} */,
  {32'hbf970d6c, 32'hbfa8ac8c} /* (18, 22, 24) {real, imag} */,
  {32'h3f82b29a, 32'h3f9e472b} /* (18, 22, 23) {real, imag} */,
  {32'h40a785f8, 32'h40603ff8} /* (18, 22, 22) {real, imag} */,
  {32'h40125d6a, 32'h3fb12122} /* (18, 22, 21) {real, imag} */,
  {32'h4040ff51, 32'hbe2eff50} /* (18, 22, 20) {real, imag} */,
  {32'h40294d1c, 32'hbd7008c0} /* (18, 22, 19) {real, imag} */,
  {32'h40869e9d, 32'h3ffcfa59} /* (18, 22, 18) {real, imag} */,
  {32'h408fea75, 32'h40403a2a} /* (18, 22, 17) {real, imag} */,
  {32'h402fd9c3, 32'h3f64b8c2} /* (18, 22, 16) {real, imag} */,
  {32'h3fcf9df0, 32'hbc41f200} /* (18, 22, 15) {real, imag} */,
  {32'hbfc242d8, 32'hc049c5d2} /* (18, 22, 14) {real, imag} */,
  {32'hbeadc050, 32'hbfaace96} /* (18, 22, 13) {real, imag} */,
  {32'hbfa35e59, 32'h3f6af774} /* (18, 22, 12) {real, imag} */,
  {32'h3fe024de, 32'hc025dd37} /* (18, 22, 11) {real, imag} */,
  {32'h3c1b9880, 32'hbe913078} /* (18, 22, 10) {real, imag} */,
  {32'h3e6c52f8, 32'h3c620000} /* (18, 22, 9) {real, imag} */,
  {32'hc025d774, 32'h40421b0d} /* (18, 22, 8) {real, imag} */,
  {32'hc0535a64, 32'h3fcfcf2d} /* (18, 22, 7) {real, imag} */,
  {32'h3fac560a, 32'h4060b041} /* (18, 22, 6) {real, imag} */,
  {32'h3fcf837e, 32'h400c4efd} /* (18, 22, 5) {real, imag} */,
  {32'hc01a1a50, 32'hbf8176e5} /* (18, 22, 4) {real, imag} */,
  {32'hbec3e294, 32'h4011b2ab} /* (18, 22, 3) {real, imag} */,
  {32'hbf978b15, 32'h3eccb51a} /* (18, 22, 2) {real, imag} */,
  {32'h3f9c6bf2, 32'hbff97464} /* (18, 22, 1) {real, imag} */,
  {32'h3fcb125e, 32'h3e988392} /* (18, 22, 0) {real, imag} */,
  {32'hc01001e6, 32'h3fc5fac9} /* (18, 21, 31) {real, imag} */,
  {32'hc0532f8a, 32'h3e2c7c18} /* (18, 21, 30) {real, imag} */,
  {32'hc03891ca, 32'hc001f6fa} /* (18, 21, 29) {real, imag} */,
  {32'hbf52b842, 32'hc073449f} /* (18, 21, 28) {real, imag} */,
  {32'h3e2c9fb4, 32'hc0266420} /* (18, 21, 27) {real, imag} */,
  {32'hbf866aec, 32'h3fc2428f} /* (18, 21, 26) {real, imag} */,
  {32'hbd0c0980, 32'h3e1fa440} /* (18, 21, 25) {real, imag} */,
  {32'hbed0737c, 32'hc00d58c7} /* (18, 21, 24) {real, imag} */,
  {32'h400c11ba, 32'h3dfaec90} /* (18, 21, 23) {real, imag} */,
  {32'hbef02e08, 32'h3ec47d5a} /* (18, 21, 22) {real, imag} */,
  {32'h40209dd6, 32'h3e9ae42c} /* (18, 21, 21) {real, imag} */,
  {32'h402a99cb, 32'hbf87fa8a} /* (18, 21, 20) {real, imag} */,
  {32'hbf5b756d, 32'hbf69546c} /* (18, 21, 19) {real, imag} */,
  {32'hc0030720, 32'hbf919dce} /* (18, 21, 18) {real, imag} */,
  {32'hbfc2f4b9, 32'h4019c7ff} /* (18, 21, 17) {real, imag} */,
  {32'hbf30bad1, 32'h3f8568b5} /* (18, 21, 16) {real, imag} */,
  {32'h3df4e500, 32'h4064ddc4} /* (18, 21, 15) {real, imag} */,
  {32'h3f04b052, 32'h3fc7cc20} /* (18, 21, 14) {real, imag} */,
  {32'hbe21f1a8, 32'hbfe1e07b} /* (18, 21, 13) {real, imag} */,
  {32'h3eb75921, 32'hc05d94fe} /* (18, 21, 12) {real, imag} */,
  {32'h3eaff75a, 32'hbf1b8c4a} /* (18, 21, 11) {real, imag} */,
  {32'h3f41a029, 32'hbf3256eb} /* (18, 21, 10) {real, imag} */,
  {32'h3f5361de, 32'h3eea32ac} /* (18, 21, 9) {real, imag} */,
  {32'h3f0fa9ac, 32'hbfecdcb6} /* (18, 21, 8) {real, imag} */,
  {32'hbfd4bf99, 32'hbfecdb53} /* (18, 21, 7) {real, imag} */,
  {32'h3e0d2cd0, 32'hc04dd110} /* (18, 21, 6) {real, imag} */,
  {32'h3f2c6950, 32'hc07466aa} /* (18, 21, 5) {real, imag} */,
  {32'hbf071594, 32'hbf6bddc8} /* (18, 21, 4) {real, imag} */,
  {32'h406e3070, 32'h4006133a} /* (18, 21, 3) {real, imag} */,
  {32'h3db2d8f8, 32'h40390401} /* (18, 21, 2) {real, imag} */,
  {32'h3f903c2a, 32'h3eec9a38} /* (18, 21, 1) {real, imag} */,
  {32'h3f98bf3e, 32'h3e8bf856} /* (18, 21, 0) {real, imag} */,
  {32'hc011a4aa, 32'h3fa60270} /* (18, 20, 31) {real, imag} */,
  {32'hc0404609, 32'h4036ba66} /* (18, 20, 30) {real, imag} */,
  {32'hbe83a8f0, 32'h4099059c} /* (18, 20, 29) {real, imag} */,
  {32'h3f3d6582, 32'h4091fec4} /* (18, 20, 28) {real, imag} */,
  {32'hbf594d2a, 32'h401d53a4} /* (18, 20, 27) {real, imag} */,
  {32'h3ffe5550, 32'h3fb2b5a5} /* (18, 20, 26) {real, imag} */,
  {32'h3ff9d16a, 32'hbdf61260} /* (18, 20, 25) {real, imag} */,
  {32'hbf32be2c, 32'hc04077ce} /* (18, 20, 24) {real, imag} */,
  {32'h3f78fcdf, 32'hbf8612d5} /* (18, 20, 23) {real, imag} */,
  {32'h3d707b40, 32'h3f9bedc1} /* (18, 20, 22) {real, imag} */,
  {32'hc04933b8, 32'h404f9e38} /* (18, 20, 21) {real, imag} */,
  {32'hc02cbecd, 32'h403da859} /* (18, 20, 20) {real, imag} */,
  {32'h3fc71922, 32'h400b2b4c} /* (18, 20, 19) {real, imag} */,
  {32'h40085ab4, 32'h3f68847c} /* (18, 20, 18) {real, imag} */,
  {32'h3fe4f1b6, 32'hbff1ba7a} /* (18, 20, 17) {real, imag} */,
  {32'h3f305852, 32'hbe8c6c6c} /* (18, 20, 16) {real, imag} */,
  {32'hbfb46538, 32'hbd0264c0} /* (18, 20, 15) {real, imag} */,
  {32'hbed9ff78, 32'hbe888e88} /* (18, 20, 14) {real, imag} */,
  {32'hbfd88545, 32'h3fc8c6e6} /* (18, 20, 13) {real, imag} */,
  {32'hbfdd9a3e, 32'h3f4ab0d0} /* (18, 20, 12) {real, imag} */,
  {32'hbff9238e, 32'hc00ff512} /* (18, 20, 11) {real, imag} */,
  {32'h3f62606c, 32'h3e994f5f} /* (18, 20, 10) {real, imag} */,
  {32'h3fc3f227, 32'h406768d9} /* (18, 20, 9) {real, imag} */,
  {32'h3f7b37ac, 32'h3e3ddeb0} /* (18, 20, 8) {real, imag} */,
  {32'h3f63f81e, 32'hbdd4b9c8} /* (18, 20, 7) {real, imag} */,
  {32'h3fc4d392, 32'hbf86d756} /* (18, 20, 6) {real, imag} */,
  {32'h3f089870, 32'h3faf80de} /* (18, 20, 5) {real, imag} */,
  {32'hbfb28c3a, 32'h3d438100} /* (18, 20, 4) {real, imag} */,
  {32'hbe6ca250, 32'h3eace848} /* (18, 20, 3) {real, imag} */,
  {32'h3f321600, 32'h3fa97218} /* (18, 20, 2) {real, imag} */,
  {32'h3fce7df8, 32'h40084484} /* (18, 20, 1) {real, imag} */,
  {32'hbf577c3d, 32'h3fcccc8e} /* (18, 20, 0) {real, imag} */,
  {32'hbf13d383, 32'hbfc6f2ef} /* (18, 19, 31) {real, imag} */,
  {32'h3fbfcf0a, 32'hbfcd86a6} /* (18, 19, 30) {real, imag} */,
  {32'h3ee81d24, 32'hbeeeae64} /* (18, 19, 29) {real, imag} */,
  {32'hbfe982cd, 32'hbf878f7e} /* (18, 19, 28) {real, imag} */,
  {32'hbf58984a, 32'h3fdcea8a} /* (18, 19, 27) {real, imag} */,
  {32'h3cd14690, 32'h3f9c5225} /* (18, 19, 26) {real, imag} */,
  {32'hbf3b6138, 32'hbe9a3e34} /* (18, 19, 25) {real, imag} */,
  {32'hbff6d64f, 32'h3fe8d730} /* (18, 19, 24) {real, imag} */,
  {32'hc03f2231, 32'h4048d0db} /* (18, 19, 23) {real, imag} */,
  {32'hbf85a93f, 32'h3e60c930} /* (18, 19, 22) {real, imag} */,
  {32'hbf70bb9c, 32'hbf8a1ef8} /* (18, 19, 21) {real, imag} */,
  {32'hbfd54adb, 32'h3ffb0740} /* (18, 19, 20) {real, imag} */,
  {32'hbc402b80, 32'h3fb232f4} /* (18, 19, 19) {real, imag} */,
  {32'hbebe05ce, 32'hc0088969} /* (18, 19, 18) {real, imag} */,
  {32'hc01b6162, 32'hbeb6fa44} /* (18, 19, 17) {real, imag} */,
  {32'hbfb70f1c, 32'h3f6cdb3a} /* (18, 19, 16) {real, imag} */,
  {32'hbe69479c, 32'hbf7596ad} /* (18, 19, 15) {real, imag} */,
  {32'hbe5b4bac, 32'hbf762414} /* (18, 19, 14) {real, imag} */,
  {32'h3f8e7f38, 32'hbf82ac0e} /* (18, 19, 13) {real, imag} */,
  {32'hc0163b95, 32'hbed13ab2} /* (18, 19, 12) {real, imag} */,
  {32'hc056608a, 32'hbe8f8b14} /* (18, 19, 11) {real, imag} */,
  {32'hbfff4b68, 32'h40034d4a} /* (18, 19, 10) {real, imag} */,
  {32'hbfbaa655, 32'h3eb66e68} /* (18, 19, 9) {real, imag} */,
  {32'hbe6a65c4, 32'h3ee6cad8} /* (18, 19, 8) {real, imag} */,
  {32'h3cf14e00, 32'h3f440060} /* (18, 19, 7) {real, imag} */,
  {32'hbda67fb4, 32'h402326cd} /* (18, 19, 6) {real, imag} */,
  {32'hbf2d4c9b, 32'h40651635} /* (18, 19, 5) {real, imag} */,
  {32'hc01955e6, 32'h3d7092b0} /* (18, 19, 4) {real, imag} */,
  {32'hbecdd738, 32'hbfa72134} /* (18, 19, 3) {real, imag} */,
  {32'hbf0ed384, 32'h3d152790} /* (18, 19, 2) {real, imag} */,
  {32'hbfa18619, 32'h3f1c0057} /* (18, 19, 1) {real, imag} */,
  {32'hbf4e93f6, 32'hbeaf2ab4} /* (18, 19, 0) {real, imag} */,
  {32'h3f892154, 32'hbf2a8d28} /* (18, 18, 31) {real, imag} */,
  {32'hbdc03ae0, 32'hbed0c2de} /* (18, 18, 30) {real, imag} */,
  {32'hc006dc20, 32'h3ef2c9b8} /* (18, 18, 29) {real, imag} */,
  {32'h3d979a18, 32'h3f2c7a68} /* (18, 18, 28) {real, imag} */,
  {32'h3fd2869c, 32'h3f09a8ee} /* (18, 18, 27) {real, imag} */,
  {32'h3f80f833, 32'h3f11e380} /* (18, 18, 26) {real, imag} */,
  {32'hbe392b64, 32'hbc97be80} /* (18, 18, 25) {real, imag} */,
  {32'hbef35446, 32'hbd637220} /* (18, 18, 24) {real, imag} */,
  {32'hbf991d97, 32'hbfc655da} /* (18, 18, 23) {real, imag} */,
  {32'hc0136895, 32'hbed4db6b} /* (18, 18, 22) {real, imag} */,
  {32'h3f1125b0, 32'h3fb4ad84} /* (18, 18, 21) {real, imag} */,
  {32'h3f78cfe0, 32'h3f7505ae} /* (18, 18, 20) {real, imag} */,
  {32'hc00d71cd, 32'hbf071696} /* (18, 18, 19) {real, imag} */,
  {32'hc0258545, 32'hbec6c918} /* (18, 18, 18) {real, imag} */,
  {32'hbfb7664d, 32'h3e4f45a0} /* (18, 18, 17) {real, imag} */,
  {32'hbe2faedc, 32'h3ea93ec8} /* (18, 18, 16) {real, imag} */,
  {32'h3fe37d91, 32'h3d6f2ac0} /* (18, 18, 15) {real, imag} */,
  {32'h3fe99844, 32'h3f9402f0} /* (18, 18, 14) {real, imag} */,
  {32'h3fad6730, 32'h3f39da30} /* (18, 18, 13) {real, imag} */,
  {32'hbc64c780, 32'h3e082368} /* (18, 18, 12) {real, imag} */,
  {32'hbeb9c648, 32'hbf25e324} /* (18, 18, 11) {real, imag} */,
  {32'h3e8b5f88, 32'h3f6c3ca5} /* (18, 18, 10) {real, imag} */,
  {32'hbea090a4, 32'h3f83d5d1} /* (18, 18, 9) {real, imag} */,
  {32'hbf942d90, 32'hbf027616} /* (18, 18, 8) {real, imag} */,
  {32'h3f4cd7ac, 32'hc02418d1} /* (18, 18, 7) {real, imag} */,
  {32'h4009c320, 32'hbfd60aa5} /* (18, 18, 6) {real, imag} */,
  {32'h3f2063ba, 32'h3e7fa7a4} /* (18, 18, 5) {real, imag} */,
  {32'hbfb814fc, 32'hbefd3e47} /* (18, 18, 4) {real, imag} */,
  {32'h3f474310, 32'h3e6d9fca} /* (18, 18, 3) {real, imag} */,
  {32'hbce31580, 32'h3f389314} /* (18, 18, 2) {real, imag} */,
  {32'hbf058e6e, 32'hbbb9a200} /* (18, 18, 1) {real, imag} */,
  {32'h3f910cd4, 32'h3f3e826d} /* (18, 18, 0) {real, imag} */,
  {32'h3f23c0c4, 32'h3f4dd022} /* (18, 17, 31) {real, imag} */,
  {32'h3f01e37f, 32'h400aadaa} /* (18, 17, 30) {real, imag} */,
  {32'h3efed134, 32'h3f163bbc} /* (18, 17, 29) {real, imag} */,
  {32'h3f8565e1, 32'h3dde3aee} /* (18, 17, 28) {real, imag} */,
  {32'h3e519338, 32'h3fa53bc4} /* (18, 17, 27) {real, imag} */,
  {32'h3d424080, 32'h3fe79221} /* (18, 17, 26) {real, imag} */,
  {32'hbfe5ebcc, 32'h3f0e562e} /* (18, 17, 25) {real, imag} */,
  {32'hbf848b9a, 32'h3ec5478c} /* (18, 17, 24) {real, imag} */,
  {32'h3f3a7b10, 32'h3f368ba1} /* (18, 17, 23) {real, imag} */,
  {32'h3f3010c4, 32'h3fa2a7fb} /* (18, 17, 22) {real, imag} */,
  {32'hbeedb37c, 32'h4002f560} /* (18, 17, 21) {real, imag} */,
  {32'hbfd23277, 32'h3f8b35a4} /* (18, 17, 20) {real, imag} */,
  {32'h3f1bcdc3, 32'hbef703a9} /* (18, 17, 19) {real, imag} */,
  {32'hbde3c4c0, 32'hc002bfea} /* (18, 17, 18) {real, imag} */,
  {32'hc012ed34, 32'hc03b508d} /* (18, 17, 17) {real, imag} */,
  {32'hbf7658f2, 32'hbf414180} /* (18, 17, 16) {real, imag} */,
  {32'hbd78c8b0, 32'hbeea78c6} /* (18, 17, 15) {real, imag} */,
  {32'hbf4d3c31, 32'h3edbb5f1} /* (18, 17, 14) {real, imag} */,
  {32'hbeca6288, 32'hbc35a240} /* (18, 17, 13) {real, imag} */,
  {32'h3f161f9a, 32'hbf6a8078} /* (18, 17, 12) {real, imag} */,
  {32'h3e1c69e0, 32'hbf2ef2e7} /* (18, 17, 11) {real, imag} */,
  {32'hbdeaf5d0, 32'h3df377a0} /* (18, 17, 10) {real, imag} */,
  {32'hbf061b44, 32'h3bae3200} /* (18, 17, 9) {real, imag} */,
  {32'hc00960f0, 32'hbf96e2dc} /* (18, 17, 8) {real, imag} */,
  {32'h3e681e48, 32'hbe80b32a} /* (18, 17, 7) {real, imag} */,
  {32'hbe3b9320, 32'h3fc5d2ee} /* (18, 17, 6) {real, imag} */,
  {32'hc010c698, 32'hbd8bcab0} /* (18, 17, 5) {real, imag} */,
  {32'hbff0e736, 32'h3f612980} /* (18, 17, 4) {real, imag} */,
  {32'hbfb794ac, 32'h3f0b27e3} /* (18, 17, 3) {real, imag} */,
  {32'hbfcf4e30, 32'hbf05a6d7} /* (18, 17, 2) {real, imag} */,
  {32'hbea8af6c, 32'hbeffa358} /* (18, 17, 1) {real, imag} */,
  {32'h3f1dca16, 32'h3ee6ab12} /* (18, 17, 0) {real, imag} */,
  {32'hbee380f8, 32'h3cae5d80} /* (18, 16, 31) {real, imag} */,
  {32'h3e1b1a40, 32'h3f7d04dc} /* (18, 16, 30) {real, imag} */,
  {32'hbe33c43c, 32'h3fdb7328} /* (18, 16, 29) {real, imag} */,
  {32'hbf0d41ba, 32'h3f291148} /* (18, 16, 28) {real, imag} */,
  {32'hbccf1700, 32'hbf5084d8} /* (18, 16, 27) {real, imag} */,
  {32'h3f5447d0, 32'hbf00ad10} /* (18, 16, 26) {real, imag} */,
  {32'h3eb4f060, 32'hbd883ea0} /* (18, 16, 25) {real, imag} */,
  {32'hbe43f620, 32'h3d8d5fe0} /* (18, 16, 24) {real, imag} */,
  {32'h3e0517d0, 32'h3f9a36b2} /* (18, 16, 23) {real, imag} */,
  {32'hbf1b9998, 32'h3e9c3b30} /* (18, 16, 22) {real, imag} */,
  {32'hbfc9a588, 32'hbf8718b7} /* (18, 16, 21) {real, imag} */,
  {32'hbfd9f490, 32'h3ee974ec} /* (18, 16, 20) {real, imag} */,
  {32'hbeae2cac, 32'h3f1be314} /* (18, 16, 19) {real, imag} */,
  {32'h3e2f8200, 32'hbe229880} /* (18, 16, 18) {real, imag} */,
  {32'hbedd7fdc, 32'hbfbef9d8} /* (18, 16, 17) {real, imag} */,
  {32'hbf2485b7, 32'hbf92ff9c} /* (18, 16, 16) {real, imag} */,
  {32'hbe21c020, 32'hbfb0fa2c} /* (18, 16, 15) {real, imag} */,
  {32'h3f2e6dac, 32'hbfd24d24} /* (18, 16, 14) {real, imag} */,
  {32'h3f99edab, 32'hbf3a6544} /* (18, 16, 13) {real, imag} */,
  {32'h3f4f67b5, 32'hbfa71b36} /* (18, 16, 12) {real, imag} */,
  {32'h3faf6661, 32'hbeb5d698} /* (18, 16, 11) {real, imag} */,
  {32'h3fd8ed88, 32'h3f8b2e44} /* (18, 16, 10) {real, imag} */,
  {32'h3f4a7c08, 32'h3f39f63c} /* (18, 16, 9) {real, imag} */,
  {32'h40196eda, 32'hbeafc930} /* (18, 16, 8) {real, imag} */,
  {32'h3fb9ea1c, 32'hbf7499c0} /* (18, 16, 7) {real, imag} */,
  {32'hbe15bce0, 32'h3d7f3480} /* (18, 16, 6) {real, imag} */,
  {32'hbf2eed10, 32'hbe85e7a0} /* (18, 16, 5) {real, imag} */,
  {32'hbf2da678, 32'h3fa09c14} /* (18, 16, 4) {real, imag} */,
  {32'hbcf60c00, 32'h3f838bea} /* (18, 16, 3) {real, imag} */,
  {32'hbf1c5bb8, 32'hbf29a9cc} /* (18, 16, 2) {real, imag} */,
  {32'h3e2dccbc, 32'hbe3f8c20} /* (18, 16, 1) {real, imag} */,
  {32'h3e20320c, 32'h3e4dc210} /* (18, 16, 0) {real, imag} */,
  {32'h3f7303e4, 32'h3fcf3c91} /* (18, 15, 31) {real, imag} */,
  {32'h3db0f708, 32'h3fc10898} /* (18, 15, 30) {real, imag} */,
  {32'hbf13ac3a, 32'h3fc42eba} /* (18, 15, 29) {real, imag} */,
  {32'hbd03d120, 32'hbed98f4a} /* (18, 15, 28) {real, imag} */,
  {32'hbf86419f, 32'hbf95a1fe} /* (18, 15, 27) {real, imag} */,
  {32'hbe0e0120, 32'h3ef310ac} /* (18, 15, 26) {real, imag} */,
  {32'h3f92aae4, 32'h3fa96e77} /* (18, 15, 25) {real, imag} */,
  {32'h3f19e834, 32'h3f43ffee} /* (18, 15, 24) {real, imag} */,
  {32'hbfb060b8, 32'h3f7f3ff9} /* (18, 15, 23) {real, imag} */,
  {32'hbdfae560, 32'h3ebbef0d} /* (18, 15, 22) {real, imag} */,
  {32'hbd1569a0, 32'hbf040883} /* (18, 15, 21) {real, imag} */,
  {32'h3f940593, 32'h3da4eae8} /* (18, 15, 20) {real, imag} */,
  {32'h3fa626a4, 32'h3e0deb2a} /* (18, 15, 19) {real, imag} */,
  {32'hbf93cd2c, 32'hbf2def88} /* (18, 15, 18) {real, imag} */,
  {32'hbea430c0, 32'hbe8418b8} /* (18, 15, 17) {real, imag} */,
  {32'h3f26612a, 32'h3daea5c4} /* (18, 15, 16) {real, imag} */,
  {32'hbf5d140d, 32'h3f92933c} /* (18, 15, 15) {real, imag} */,
  {32'h3e665c84, 32'h3efcadd7} /* (18, 15, 14) {real, imag} */,
  {32'hbe7352b0, 32'hbe12789c} /* (18, 15, 13) {real, imag} */,
  {32'h3f9076d7, 32'hbf9c4b40} /* (18, 15, 12) {real, imag} */,
  {32'h4013d6ec, 32'hbf95aaae} /* (18, 15, 11) {real, imag} */,
  {32'h400e132c, 32'hbf0cfe64} /* (18, 15, 10) {real, imag} */,
  {32'h3f2007a8, 32'h3ee005f8} /* (18, 15, 9) {real, imag} */,
  {32'hbf9c7bd9, 32'h3f7ed8f8} /* (18, 15, 8) {real, imag} */,
  {32'h3f0087fe, 32'h3f5f62ab} /* (18, 15, 7) {real, imag} */,
  {32'hbee5bb80, 32'hbe91dc68} /* (18, 15, 6) {real, imag} */,
  {32'hc00b955c, 32'hc00c0c02} /* (18, 15, 5) {real, imag} */,
  {32'h3ec49ec8, 32'hbf5443d0} /* (18, 15, 4) {real, imag} */,
  {32'h3fa0f618, 32'hbfc81560} /* (18, 15, 3) {real, imag} */,
  {32'hbf9aec10, 32'hbf4bfa2f} /* (18, 15, 2) {real, imag} */,
  {32'h3debbe30, 32'h3ebe6304} /* (18, 15, 1) {real, imag} */,
  {32'h3e9e9f05, 32'hbe71a1a4} /* (18, 15, 0) {real, imag} */,
  {32'hbe833a30, 32'hbf29d4e0} /* (18, 14, 31) {real, imag} */,
  {32'hbf7ae61c, 32'h3ff765ae} /* (18, 14, 30) {real, imag} */,
  {32'hbfb00521, 32'h3f25168c} /* (18, 14, 29) {real, imag} */,
  {32'hbf95bee6, 32'h3fbef6f8} /* (18, 14, 28) {real, imag} */,
  {32'hbf525b58, 32'h3fa8100f} /* (18, 14, 27) {real, imag} */,
  {32'h3f43bc9a, 32'hbfa5195a} /* (18, 14, 26) {real, imag} */,
  {32'hbf4b775f, 32'hbf746184} /* (18, 14, 25) {real, imag} */,
  {32'hbf2d697d, 32'h3f8a56d2} /* (18, 14, 24) {real, imag} */,
  {32'h40060c52, 32'h3ff4e86e} /* (18, 14, 23) {real, imag} */,
  {32'hbe805198, 32'hbdfa2f54} /* (18, 14, 22) {real, imag} */,
  {32'hbfb863c4, 32'hbf5ea8af} /* (18, 14, 21) {real, imag} */,
  {32'hbe83fb40, 32'hbf574ee2} /* (18, 14, 20) {real, imag} */,
  {32'hbf4313ab, 32'hbffcb853} /* (18, 14, 19) {real, imag} */,
  {32'hbef97df8, 32'hc013a7ab} /* (18, 14, 18) {real, imag} */,
  {32'hbf319a26, 32'hbe23df70} /* (18, 14, 17) {real, imag} */,
  {32'h3f9bcd2c, 32'h3f3c8ef4} /* (18, 14, 16) {real, imag} */,
  {32'h3fdc02d7, 32'h3e1faff0} /* (18, 14, 15) {real, imag} */,
  {32'hbe4f1e60, 32'h3f26de3f} /* (18, 14, 14) {real, imag} */,
  {32'h3f2fe898, 32'h3e999850} /* (18, 14, 13) {real, imag} */,
  {32'hbe629708, 32'hbfd3ca5d} /* (18, 14, 12) {real, imag} */,
  {32'hbfc81360, 32'hbf30cbb4} /* (18, 14, 11) {real, imag} */,
  {32'hbf9d5796, 32'h3f0ffd1b} /* (18, 14, 10) {real, imag} */,
  {32'hbebc35dc, 32'hbf0a454e} /* (18, 14, 9) {real, imag} */,
  {32'h3f8e7ec0, 32'hbea014d4} /* (18, 14, 8) {real, imag} */,
  {32'hbf8c9f7e, 32'h3f1562c0} /* (18, 14, 7) {real, imag} */,
  {32'hbed4623c, 32'h3fc78da7} /* (18, 14, 6) {real, imag} */,
  {32'h3dbe8db0, 32'h3f54efff} /* (18, 14, 5) {real, imag} */,
  {32'hbc249e40, 32'h3df0dd64} /* (18, 14, 4) {real, imag} */,
  {32'h3ed0cc00, 32'hbe744666} /* (18, 14, 3) {real, imag} */,
  {32'h400403e7, 32'hbe1c61e0} /* (18, 14, 2) {real, imag} */,
  {32'h3f7a29be, 32'h402bae85} /* (18, 14, 1) {real, imag} */,
  {32'h3bcbb080, 32'h3ec01826} /* (18, 14, 0) {real, imag} */,
  {32'h3f9ab9f0, 32'h3d878890} /* (18, 13, 31) {real, imag} */,
  {32'h3db976a0, 32'h3e259570} /* (18, 13, 30) {real, imag} */,
  {32'hbf6b5d6a, 32'hbf49fc2a} /* (18, 13, 29) {real, imag} */,
  {32'hbfd352a7, 32'hbef6a418} /* (18, 13, 28) {real, imag} */,
  {32'hc0401c98, 32'hbfa9e0fe} /* (18, 13, 27) {real, imag} */,
  {32'hbf3f3904, 32'hbf0d17ee} /* (18, 13, 26) {real, imag} */,
  {32'h3fa1d096, 32'hbf9bfc24} /* (18, 13, 25) {real, imag} */,
  {32'h3cce7440, 32'hc0469f08} /* (18, 13, 24) {real, imag} */,
  {32'hbec17408, 32'hbfff0a52} /* (18, 13, 23) {real, imag} */,
  {32'hbfbe4c5f, 32'hc006ac2f} /* (18, 13, 22) {real, imag} */,
  {32'hbfd60a22, 32'h3d230ad0} /* (18, 13, 21) {real, imag} */,
  {32'hbdf675b0, 32'h3f2c9c88} /* (18, 13, 20) {real, imag} */,
  {32'h3ed09c14, 32'h3f04c7f3} /* (18, 13, 19) {real, imag} */,
  {32'hbfd0b784, 32'hbfa4ffda} /* (18, 13, 18) {real, imag} */,
  {32'hbfb8dad9, 32'hbfebe3fd} /* (18, 13, 17) {real, imag} */,
  {32'h3de79588, 32'hbf0c8052} /* (18, 13, 16) {real, imag} */,
  {32'h3f9159e0, 32'hbf5c27c9} /* (18, 13, 15) {real, imag} */,
  {32'hbf9e4e74, 32'hbf2c4af4} /* (18, 13, 14) {real, imag} */,
  {32'hbfcda936, 32'h3f3ee52c} /* (18, 13, 13) {real, imag} */,
  {32'hbf363754, 32'hbee3fb2a} /* (18, 13, 12) {real, imag} */,
  {32'h3f69cf60, 32'h3d263460} /* (18, 13, 11) {real, imag} */,
  {32'h3e984fb6, 32'h402661f6} /* (18, 13, 10) {real, imag} */,
  {32'h3ec4b7d4, 32'h402a19ea} /* (18, 13, 9) {real, imag} */,
  {32'h3efd2d52, 32'h3f9c78f2} /* (18, 13, 8) {real, imag} */,
  {32'h3fe0f374, 32'hbfdb8f64} /* (18, 13, 7) {real, imag} */,
  {32'h3e4f83ea, 32'hbfd6d016} /* (18, 13, 6) {real, imag} */,
  {32'h3e6349f4, 32'h3f3665cc} /* (18, 13, 5) {real, imag} */,
  {32'h3eee850c, 32'hbfb98596} /* (18, 13, 4) {real, imag} */,
  {32'hbf824dee, 32'hbf94b18a} /* (18, 13, 3) {real, imag} */,
  {32'hbff972b2, 32'hbfb62ccc} /* (18, 13, 2) {real, imag} */,
  {32'hc062279a, 32'hbed448fe} /* (18, 13, 1) {real, imag} */,
  {32'hbffa76f7, 32'h3f1881e6} /* (18, 13, 0) {real, imag} */,
  {32'h3f2dd11e, 32'h400fab6b} /* (18, 12, 31) {real, imag} */,
  {32'h4005be09, 32'h40083148} /* (18, 12, 30) {real, imag} */,
  {32'h404013ee, 32'hbe9f6b18} /* (18, 12, 29) {real, imag} */,
  {32'h40242788, 32'hbf146854} /* (18, 12, 28) {real, imag} */,
  {32'h3ef1313c, 32'hbea49880} /* (18, 12, 27) {real, imag} */,
  {32'hbff7e1ac, 32'hbe8586bc} /* (18, 12, 26) {real, imag} */,
  {32'hbf8ad0e4, 32'hbfb0b624} /* (18, 12, 25) {real, imag} */,
  {32'hbf2cfa28, 32'hbdc0c550} /* (18, 12, 24) {real, imag} */,
  {32'hbdf6bfc8, 32'hbd949390} /* (18, 12, 23) {real, imag} */,
  {32'h402cabdb, 32'h3f9fb8f3} /* (18, 12, 22) {real, imag} */,
  {32'h3f591ca6, 32'h3f723080} /* (18, 12, 21) {real, imag} */,
  {32'hbf9878d2, 32'h3fdfcfea} /* (18, 12, 20) {real, imag} */,
  {32'hbeca9d88, 32'h3eb1e640} /* (18, 12, 19) {real, imag} */,
  {32'hbf265c89, 32'h3fdff888} /* (18, 12, 18) {real, imag} */,
  {32'h3f571cec, 32'h404e1abb} /* (18, 12, 17) {real, imag} */,
  {32'h3fb98817, 32'hbe2bc698} /* (18, 12, 16) {real, imag} */,
  {32'h3f664728, 32'hc050e75f} /* (18, 12, 15) {real, imag} */,
  {32'h3f04d35e, 32'hc034a891} /* (18, 12, 14) {real, imag} */,
  {32'h3fd01609, 32'hc080cb86} /* (18, 12, 13) {real, imag} */,
  {32'h3e8eab18, 32'hc07b8334} /* (18, 12, 12) {real, imag} */,
  {32'h3fad704a, 32'h4005bfea} /* (18, 12, 11) {real, imag} */,
  {32'h3eb46fc4, 32'h3f23a172} /* (18, 12, 10) {real, imag} */,
  {32'h3e896f1c, 32'hbfa9e8fe} /* (18, 12, 9) {real, imag} */,
  {32'h3ffcf30a, 32'h3faff2ae} /* (18, 12, 8) {real, imag} */,
  {32'hbf87218b, 32'h3d7e4d10} /* (18, 12, 7) {real, imag} */,
  {32'hbfd9c9ae, 32'hc0333971} /* (18, 12, 6) {real, imag} */,
  {32'h3faf2f10, 32'hbf64c338} /* (18, 12, 5) {real, imag} */,
  {32'h3ff4cc6e, 32'h3fc66234} /* (18, 12, 4) {real, imag} */,
  {32'hbc542d00, 32'h404a3a41} /* (18, 12, 3) {real, imag} */,
  {32'h3f0db810, 32'h400401ee} /* (18, 12, 2) {real, imag} */,
  {32'hbfea1df4, 32'hc0090df4} /* (18, 12, 1) {real, imag} */,
  {32'hbfbf3f6c, 32'hbfa64c12} /* (18, 12, 0) {real, imag} */,
  {32'h3fa8fc89, 32'hbff8c1cf} /* (18, 11, 31) {real, imag} */,
  {32'h3f22434a, 32'hc0506056} /* (18, 11, 30) {real, imag} */,
  {32'hbebfa400, 32'hbfd0e368} /* (18, 11, 29) {real, imag} */,
  {32'hbfb80c87, 32'h40139201} /* (18, 11, 28) {real, imag} */,
  {32'hbff4742c, 32'h402110ee} /* (18, 11, 27) {real, imag} */,
  {32'hbe8282e0, 32'hbe210898} /* (18, 11, 26) {real, imag} */,
  {32'hbfd1053c, 32'h3e13e5d8} /* (18, 11, 25) {real, imag} */,
  {32'hbfc66301, 32'hbf0ccd74} /* (18, 11, 24) {real, imag} */,
  {32'h3e191118, 32'hc06dde6c} /* (18, 11, 23) {real, imag} */,
  {32'hc011b208, 32'h3f56d281} /* (18, 11, 22) {real, imag} */,
  {32'hbf50c20a, 32'h400a661e} /* (18, 11, 21) {real, imag} */,
  {32'hbf8bbe1e, 32'h4062f511} /* (18, 11, 20) {real, imag} */,
  {32'hbf88376e, 32'hbf3e5e48} /* (18, 11, 19) {real, imag} */,
  {32'hbf267b40, 32'h3f07e9e5} /* (18, 11, 18) {real, imag} */,
  {32'h3f10d636, 32'hc00128fb} /* (18, 11, 17) {real, imag} */,
  {32'hbefc943a, 32'hbf9e3243} /* (18, 11, 16) {real, imag} */,
  {32'hc095a456, 32'h4052fdfc} /* (18, 11, 15) {real, imag} */,
  {32'hc0853bfe, 32'h3f6e3918} /* (18, 11, 14) {real, imag} */,
  {32'hbfe8e16f, 32'h40a673fd} /* (18, 11, 13) {real, imag} */,
  {32'h3d013508, 32'h40a8b393} /* (18, 11, 12) {real, imag} */,
  {32'hbea498ba, 32'hbc049b80} /* (18, 11, 11) {real, imag} */,
  {32'h3e3eb694, 32'hbe8c1fce} /* (18, 11, 10) {real, imag} */,
  {32'h3ed1cafc, 32'h3f392ef6} /* (18, 11, 9) {real, imag} */,
  {32'h40605161, 32'hbfddcd6e} /* (18, 11, 8) {real, imag} */,
  {32'h401c14a4, 32'hc04892a4} /* (18, 11, 7) {real, imag} */,
  {32'h3ef7a048, 32'hbfd2d49b} /* (18, 11, 6) {real, imag} */,
  {32'h3ffb4c6a, 32'h3e934470} /* (18, 11, 5) {real, imag} */,
  {32'h3fb017c6, 32'hbf1a00a4} /* (18, 11, 4) {real, imag} */,
  {32'h3e38b5a0, 32'h3f67243a} /* (18, 11, 3) {real, imag} */,
  {32'hbf1b9755, 32'h4076b4f9} /* (18, 11, 2) {real, imag} */,
  {32'h4027a89f, 32'h404b818d} /* (18, 11, 1) {real, imag} */,
  {32'h406daddd, 32'h3fe37588} /* (18, 11, 0) {real, imag} */,
  {32'hc03f910a, 32'hbfbf7b73} /* (18, 10, 31) {real, imag} */,
  {32'h402d4ff2, 32'h3e872194} /* (18, 10, 30) {real, imag} */,
  {32'h408e6406, 32'h3dcae9c0} /* (18, 10, 29) {real, imag} */,
  {32'h40655eb3, 32'h3fe983fc} /* (18, 10, 28) {real, imag} */,
  {32'h4066a9c8, 32'h4031cb88} /* (18, 10, 27) {real, imag} */,
  {32'hbefaa9f8, 32'h3f84bc10} /* (18, 10, 26) {real, imag} */,
  {32'hc039a18f, 32'hbe9b8416} /* (18, 10, 25) {real, imag} */,
  {32'hbf26ee6f, 32'hc043cb94} /* (18, 10, 24) {real, imag} */,
  {32'hc01d7fc3, 32'hbf8f32ef} /* (18, 10, 23) {real, imag} */,
  {32'h3f2fa630, 32'h3e438028} /* (18, 10, 22) {real, imag} */,
  {32'h4022ad9e, 32'h3ff295fa} /* (18, 10, 21) {real, imag} */,
  {32'h3fa3d4e6, 32'h3fa2836e} /* (18, 10, 20) {real, imag} */,
  {32'h3fd29e85, 32'hbfe310da} /* (18, 10, 19) {real, imag} */,
  {32'h407ab512, 32'hbd944c70} /* (18, 10, 18) {real, imag} */,
  {32'hbc6eee00, 32'h3f190f22} /* (18, 10, 17) {real, imag} */,
  {32'hbfa773ee, 32'hbf93c99f} /* (18, 10, 16) {real, imag} */,
  {32'hbf0066af, 32'hc002642c} /* (18, 10, 15) {real, imag} */,
  {32'hbfeb3328, 32'h3f14ad10} /* (18, 10, 14) {real, imag} */,
  {32'hbfda65e8, 32'h404403e1} /* (18, 10, 13) {real, imag} */,
  {32'h3f14eba2, 32'hbed8cc30} /* (18, 10, 12) {real, imag} */,
  {32'h3f98c626, 32'hbfb46232} /* (18, 10, 11) {real, imag} */,
  {32'hbe491eb8, 32'hbea79dcc} /* (18, 10, 10) {real, imag} */,
  {32'hc01326ea, 32'hbf8cbc88} /* (18, 10, 9) {real, imag} */,
  {32'hc034e696, 32'hbea07928} /* (18, 10, 8) {real, imag} */,
  {32'hbd958610, 32'hc0367a04} /* (18, 10, 7) {real, imag} */,
  {32'h4018964b, 32'hc0e11380} /* (18, 10, 6) {real, imag} */,
  {32'h3fec7c9a, 32'hc099fd78} /* (18, 10, 5) {real, imag} */,
  {32'h3f3924b2, 32'hbff17eed} /* (18, 10, 4) {real, imag} */,
  {32'h400e7542, 32'hbfbec456} /* (18, 10, 3) {real, imag} */,
  {32'h3fd3d22f, 32'h3ff976ac} /* (18, 10, 2) {real, imag} */,
  {32'h3ff3582a, 32'h3fdd04c4} /* (18, 10, 1) {real, imag} */,
  {32'h3ff555ec, 32'hbfd0fb22} /* (18, 10, 0) {real, imag} */,
  {32'h3f9138d2, 32'hbfa5fae7} /* (18, 9, 31) {real, imag} */,
  {32'hbf0b57fe, 32'h3feb08a8} /* (18, 9, 30) {real, imag} */,
  {32'hbf2e2a2c, 32'h3ff5ea72} /* (18, 9, 29) {real, imag} */,
  {32'h40aa75b3, 32'hc075cf6e} /* (18, 9, 28) {real, imag} */,
  {32'h406543f8, 32'hc03eb48c} /* (18, 9, 27) {real, imag} */,
  {32'hbebd08d8, 32'h3fabd37d} /* (18, 9, 26) {real, imag} */,
  {32'hbc48b780, 32'h3febc490} /* (18, 9, 25) {real, imag} */,
  {32'h3f1efe14, 32'h406a385b} /* (18, 9, 24) {real, imag} */,
  {32'h3f93abc3, 32'h40aa6530} /* (18, 9, 23) {real, imag} */,
  {32'h3ef0db5c, 32'h4080d974} /* (18, 9, 22) {real, imag} */,
  {32'hbfbeed79, 32'hc01f48d6} /* (18, 9, 21) {real, imag} */,
  {32'hbfb82de6, 32'hc0af7e85} /* (18, 9, 20) {real, imag} */,
  {32'hbfa2e10e, 32'hc0a03874} /* (18, 9, 19) {real, imag} */,
  {32'hc06edb5d, 32'hbffc985e} /* (18, 9, 18) {real, imag} */,
  {32'hc027b4b2, 32'hbeecd224} /* (18, 9, 17) {real, imag} */,
  {32'hbef13128, 32'hbea3a24e} /* (18, 9, 16) {real, imag} */,
  {32'h3f190258, 32'hbf85cfe6} /* (18, 9, 15) {real, imag} */,
  {32'hbed2ebf4, 32'h3fe761bb} /* (18, 9, 14) {real, imag} */,
  {32'h3ee1d778, 32'h40621b35} /* (18, 9, 13) {real, imag} */,
  {32'h3f44f574, 32'hbc90bf00} /* (18, 9, 12) {real, imag} */,
  {32'h3fe006a3, 32'hc02af8e7} /* (18, 9, 11) {real, imag} */,
  {32'h3fa59c73, 32'hc009bb45} /* (18, 9, 10) {real, imag} */,
  {32'hbdc83620, 32'hc0812ad3} /* (18, 9, 9) {real, imag} */,
  {32'hc0294092, 32'hc06e0c54} /* (18, 9, 8) {real, imag} */,
  {32'hbf19a084, 32'hbe91f040} /* (18, 9, 7) {real, imag} */,
  {32'h3fa16cec, 32'h40115a4f} /* (18, 9, 6) {real, imag} */,
  {32'h3fe08334, 32'hbf0a8598} /* (18, 9, 5) {real, imag} */,
  {32'hc02dbdd2, 32'hbecfb230} /* (18, 9, 4) {real, imag} */,
  {32'hc08f662c, 32'hc006f71a} /* (18, 9, 3) {real, imag} */,
  {32'hc082b11b, 32'hc0603383} /* (18, 9, 2) {real, imag} */,
  {32'hc087f980, 32'hc0ba3d20} /* (18, 9, 1) {real, imag} */,
  {32'hbe361824, 32'hbffaf8d5} /* (18, 9, 0) {real, imag} */,
  {32'h40565c44, 32'h403b5bb4} /* (18, 8, 31) {real, imag} */,
  {32'h402e89a6, 32'hbef9f210} /* (18, 8, 30) {real, imag} */,
  {32'hc00288ff, 32'h402061f6} /* (18, 8, 29) {real, imag} */,
  {32'hbf637950, 32'h40d381c6} /* (18, 8, 28) {real, imag} */,
  {32'h3ea557f4, 32'h40607883} /* (18, 8, 27) {real, imag} */,
  {32'h3fc599e2, 32'hbf360764} /* (18, 8, 26) {real, imag} */,
  {32'h3fee3bbe, 32'hc0266b17} /* (18, 8, 25) {real, imag} */,
  {32'h3fcea4ac, 32'hc051c7b4} /* (18, 8, 24) {real, imag} */,
  {32'h409e1705, 32'hc0953677} /* (18, 8, 23) {real, imag} */,
  {32'h402f4c24, 32'hbfab66d1} /* (18, 8, 22) {real, imag} */,
  {32'h3f0812b8, 32'h3fd62803} /* (18, 8, 21) {real, imag} */,
  {32'hbf888507, 32'h3f41920c} /* (18, 8, 20) {real, imag} */,
  {32'hbfd5622f, 32'hbfefa014} /* (18, 8, 19) {real, imag} */,
  {32'h3e818694, 32'hc0aab18a} /* (18, 8, 18) {real, imag} */,
  {32'hc080f963, 32'hc01f5a7c} /* (18, 8, 17) {real, imag} */,
  {32'hc08b9647, 32'hbf294b68} /* (18, 8, 16) {real, imag} */,
  {32'h3f03960c, 32'hbded8928} /* (18, 8, 15) {real, imag} */,
  {32'h3e287ed0, 32'hbf174e7c} /* (18, 8, 14) {real, imag} */,
  {32'hc02114e0, 32'hc00d1ff1} /* (18, 8, 13) {real, imag} */,
  {32'hbf3d1544, 32'h3ff4ac2e} /* (18, 8, 12) {real, imag} */,
  {32'hbfbd5bf9, 32'hc0241d34} /* (18, 8, 11) {real, imag} */,
  {32'h3f4b5fa5, 32'hbfb32be0} /* (18, 8, 10) {real, imag} */,
  {32'hc035b004, 32'h4045bf24} /* (18, 8, 9) {real, imag} */,
  {32'h40075c91, 32'h3a840c00} /* (18, 8, 8) {real, imag} */,
  {32'h406c3411, 32'h4010214d} /* (18, 8, 7) {real, imag} */,
  {32'h408cc052, 32'h3fef75cd} /* (18, 8, 6) {real, imag} */,
  {32'h40842130, 32'h4080b453} /* (18, 8, 5) {real, imag} */,
  {32'h404e1ab3, 32'hbe91b2a8} /* (18, 8, 4) {real, imag} */,
  {32'h40554227, 32'hc0d5ca23} /* (18, 8, 3) {real, imag} */,
  {32'hc025ae21, 32'h3febbd48} /* (18, 8, 2) {real, imag} */,
  {32'hc0be3878, 32'h40851583} /* (18, 8, 1) {real, imag} */,
  {32'hc002a22f, 32'h3fdec78c} /* (18, 8, 0) {real, imag} */,
  {32'h3e6a55c0, 32'hc0aa4d4b} /* (18, 7, 31) {real, imag} */,
  {32'h3f292c80, 32'hc0c16afc} /* (18, 7, 30) {real, imag} */,
  {32'h40308dfb, 32'hc00df202} /* (18, 7, 29) {real, imag} */,
  {32'hc071922c, 32'h3f1a491e} /* (18, 7, 28) {real, imag} */,
  {32'hc08512ca, 32'h4092b820} /* (18, 7, 27) {real, imag} */,
  {32'hc00d1421, 32'h40e4be8a} /* (18, 7, 26) {real, imag} */,
  {32'hbda5da10, 32'h40961c05} /* (18, 7, 25) {real, imag} */,
  {32'hbbf4c480, 32'h40d0da60} /* (18, 7, 24) {real, imag} */,
  {32'hbfdd03f5, 32'h40a721b0} /* (18, 7, 23) {real, imag} */,
  {32'hc0923e9a, 32'h3fb99512} /* (18, 7, 22) {real, imag} */,
  {32'hc0ccc87f, 32'hbe1858c0} /* (18, 7, 21) {real, imag} */,
  {32'hc0023710, 32'h3fe8fa88} /* (18, 7, 20) {real, imag} */,
  {32'h400f772d, 32'hbf4705c2} /* (18, 7, 19) {real, imag} */,
  {32'h4069aecd, 32'hc0df2f68} /* (18, 7, 18) {real, imag} */,
  {32'h406f738e, 32'hc00e167a} /* (18, 7, 17) {real, imag} */,
  {32'h40363d54, 32'h3f9175f6} /* (18, 7, 16) {real, imag} */,
  {32'h3fc4fdb6, 32'h4040f47c} /* (18, 7, 15) {real, imag} */,
  {32'h3f878d4b, 32'h3ff69d55} /* (18, 7, 14) {real, imag} */,
  {32'h3ebb4280, 32'hbf15616d} /* (18, 7, 13) {real, imag} */,
  {32'h40a7cad6, 32'hc058a2b3} /* (18, 7, 12) {real, imag} */,
  {32'hbcdc16c0, 32'hbfc3adaf} /* (18, 7, 11) {real, imag} */,
  {32'hbed38c7e, 32'hbd0e0fa0} /* (18, 7, 10) {real, imag} */,
  {32'hc08d9c8a, 32'hbf0f7660} /* (18, 7, 9) {real, imag} */,
  {32'hc0a51034, 32'hbfec7a32} /* (18, 7, 8) {real, imag} */,
  {32'hbf8dded2, 32'hbfdcb494} /* (18, 7, 7) {real, imag} */,
  {32'h3f7d3830, 32'hbf8d2eaa} /* (18, 7, 6) {real, imag} */,
  {32'hbfec650b, 32'hbf999900} /* (18, 7, 5) {real, imag} */,
  {32'hc0369e5c, 32'hc099fa87} /* (18, 7, 4) {real, imag} */,
  {32'h3f991ec0, 32'hc0bf619d} /* (18, 7, 3) {real, imag} */,
  {32'h3f1569de, 32'hbfce943e} /* (18, 7, 2) {real, imag} */,
  {32'hbe551a18, 32'hc02f5a6c} /* (18, 7, 1) {real, imag} */,
  {32'h3ecd7118, 32'hc0b22c78} /* (18, 7, 0) {real, imag} */,
  {32'hbf2b58ac, 32'hc05c4498} /* (18, 6, 31) {real, imag} */,
  {32'hbeaad4ac, 32'hc0434a1e} /* (18, 6, 30) {real, imag} */,
  {32'h402c56eb, 32'hc0610154} /* (18, 6, 29) {real, imag} */,
  {32'h3fbbf3a0, 32'hc08b32a2} /* (18, 6, 28) {real, imag} */,
  {32'hbfda9ccd, 32'hbfe69e22} /* (18, 6, 27) {real, imag} */,
  {32'h3c300600, 32'hbfae3e41} /* (18, 6, 26) {real, imag} */,
  {32'hbf8a0a78, 32'hbfa54786} /* (18, 6, 25) {real, imag} */,
  {32'hc01f8907, 32'hbfa35900} /* (18, 6, 24) {real, imag} */,
  {32'hc0594d86, 32'h3f0a796a} /* (18, 6, 23) {real, imag} */,
  {32'h3ea442d0, 32'hc0457719} /* (18, 6, 22) {real, imag} */,
  {32'hc07521fa, 32'h3f83f0e5} /* (18, 6, 21) {real, imag} */,
  {32'h3fc78cab, 32'h3fd85f18} /* (18, 6, 20) {real, imag} */,
  {32'h408baee3, 32'h4039fd15} /* (18, 6, 19) {real, imag} */,
  {32'h403f3ad4, 32'h404d819b} /* (18, 6, 18) {real, imag} */,
  {32'hc005d564, 32'h3e2eb568} /* (18, 6, 17) {real, imag} */,
  {32'hc04630f5, 32'hbfe03017} /* (18, 6, 16) {real, imag} */,
  {32'hc0aa8b74, 32'hbfbfed7a} /* (18, 6, 15) {real, imag} */,
  {32'hc0d3f2bb, 32'hc08fc3c4} /* (18, 6, 14) {real, imag} */,
  {32'hbfa2318e, 32'hc0573ff2} /* (18, 6, 13) {real, imag} */,
  {32'hc01c4272, 32'hc07424d8} /* (18, 6, 12) {real, imag} */,
  {32'hc0e3d65c, 32'hbf659f08} /* (18, 6, 11) {real, imag} */,
  {32'hc0bd3cfe, 32'h40053b9e} /* (18, 6, 10) {real, imag} */,
  {32'h4022b8f7, 32'h4032366c} /* (18, 6, 9) {real, imag} */,
  {32'h4087360c, 32'hbf989838} /* (18, 6, 8) {real, imag} */,
  {32'hbfb89837, 32'hbfac689f} /* (18, 6, 7) {real, imag} */,
  {32'h3f05b790, 32'h3d840300} /* (18, 6, 6) {real, imag} */,
  {32'hc07683ff, 32'h3fbcc8b4} /* (18, 6, 5) {real, imag} */,
  {32'h3f223ba9, 32'h40431535} /* (18, 6, 4) {real, imag} */,
  {32'hbfb7f653, 32'hbe6d1994} /* (18, 6, 3) {real, imag} */,
  {32'hc07f8d38, 32'hc05da368} /* (18, 6, 2) {real, imag} */,
  {32'hc0325bb1, 32'hc06b9697} /* (18, 6, 1) {real, imag} */,
  {32'h3dc6d9f0, 32'hbf8da816} /* (18, 6, 0) {real, imag} */,
  {32'h4022a600, 32'hbf62ff55} /* (18, 5, 31) {real, imag} */,
  {32'h3ff97b7a, 32'hbfcfa1f4} /* (18, 5, 30) {real, imag} */,
  {32'hc0da9959, 32'h3f11118d} /* (18, 5, 29) {real, imag} */,
  {32'hc01e3425, 32'h40e811e2} /* (18, 5, 28) {real, imag} */,
  {32'hc048addb, 32'h403f0d14} /* (18, 5, 27) {real, imag} */,
  {32'h3f7e2440, 32'hc05f3f9e} /* (18, 5, 26) {real, imag} */,
  {32'h4000b4a4, 32'hbf0f71d7} /* (18, 5, 25) {real, imag} */,
  {32'h4093cbee, 32'h4035de87} /* (18, 5, 24) {real, imag} */,
  {32'h404028fc, 32'h4094e990} /* (18, 5, 23) {real, imag} */,
  {32'h3ec13830, 32'h409ef1c0} /* (18, 5, 22) {real, imag} */,
  {32'hbe7a20d8, 32'h3f0bf548} /* (18, 5, 21) {real, imag} */,
  {32'hbf52811d, 32'hc09e45cc} /* (18, 5, 20) {real, imag} */,
  {32'hc08420b1, 32'hc052de88} /* (18, 5, 19) {real, imag} */,
  {32'hc02dfd0a, 32'hc0917124} /* (18, 5, 18) {real, imag} */,
  {32'h401a3c08, 32'hbfb55e5e} /* (18, 5, 17) {real, imag} */,
  {32'h405322ba, 32'hc026553c} /* (18, 5, 16) {real, imag} */,
  {32'hbf17f590, 32'hc0aabd22} /* (18, 5, 15) {real, imag} */,
  {32'hc0ccd1d2, 32'hc0ebae3a} /* (18, 5, 14) {real, imag} */,
  {32'hbfb5fed5, 32'hc0729482} /* (18, 5, 13) {real, imag} */,
  {32'hc0460577, 32'hc1041d4c} /* (18, 5, 12) {real, imag} */,
  {32'hc0b057a4, 32'hc0bf4a87} /* (18, 5, 11) {real, imag} */,
  {32'h4079be28, 32'hc002173e} /* (18, 5, 10) {real, imag} */,
  {32'h4113bf9e, 32'hbfe2c7bc} /* (18, 5, 9) {real, imag} */,
  {32'h3f5e76ff, 32'h40a6bbf8} /* (18, 5, 8) {real, imag} */,
  {32'h3ff8fd3a, 32'h3f53a80c} /* (18, 5, 7) {real, imag} */,
  {32'h408cd43c, 32'h401f146b} /* (18, 5, 6) {real, imag} */,
  {32'h40c71147, 32'h3fa73d3c} /* (18, 5, 5) {real, imag} */,
  {32'h4133a74c, 32'hbfbfcc94} /* (18, 5, 4) {real, imag} */,
  {32'h40adf2a6, 32'h3f4e6daf} /* (18, 5, 3) {real, imag} */,
  {32'h406fca95, 32'hc073242a} /* (18, 5, 2) {real, imag} */,
  {32'h408d275f, 32'hc1220553} /* (18, 5, 1) {real, imag} */,
  {32'h3fa6c788, 32'hc013c4d0} /* (18, 5, 0) {real, imag} */,
  {32'h405a38f6, 32'hc046d552} /* (18, 4, 31) {real, imag} */,
  {32'hc09b107a, 32'hc11931ba} /* (18, 4, 30) {real, imag} */,
  {32'hc13ceb12, 32'hc1372f2d} /* (18, 4, 29) {real, imag} */,
  {32'hc0dc5cd5, 32'hc10650c7} /* (18, 4, 28) {real, imag} */,
  {32'hc10dd1a4, 32'hc081c4e5} /* (18, 4, 27) {real, imag} */,
  {32'hc0a90eda, 32'h3f89aee3} /* (18, 4, 26) {real, imag} */,
  {32'hbfcd791d, 32'h40881f8b} /* (18, 4, 25) {real, imag} */,
  {32'hbf970a72, 32'h4071d200} /* (18, 4, 24) {real, imag} */,
  {32'hc09495c2, 32'h3e4ffab8} /* (18, 4, 23) {real, imag} */,
  {32'hc095bf4e, 32'h3f114e54} /* (18, 4, 22) {real, imag} */,
  {32'h3f74f998, 32'hbf6cfa11} /* (18, 4, 21) {real, imag} */,
  {32'h4112a500, 32'h405bc9d3} /* (18, 4, 20) {real, imag} */,
  {32'h4141609c, 32'h412e4e90} /* (18, 4, 19) {real, imag} */,
  {32'hc07b2c7a, 32'h40f020b3} /* (18, 4, 18) {real, imag} */,
  {32'hc07b62e3, 32'h41166eb7} /* (18, 4, 17) {real, imag} */,
  {32'h4048f380, 32'h412908f7} /* (18, 4, 16) {real, imag} */,
  {32'h404308ea, 32'hc066011c} /* (18, 4, 15) {real, imag} */,
  {32'hc06cd05f, 32'hc0baf944} /* (18, 4, 14) {real, imag} */,
  {32'h3ef5bf90, 32'hbd9435d0} /* (18, 4, 13) {real, imag} */,
  {32'h40fb1254, 32'h40e24207} /* (18, 4, 12) {real, imag} */,
  {32'h4116763c, 32'h40d685f3} /* (18, 4, 11) {real, imag} */,
  {32'hbe0b6578, 32'h3f399aa8} /* (18, 4, 10) {real, imag} */,
  {32'hc0985371, 32'h3ff6a453} /* (18, 4, 9) {real, imag} */,
  {32'hc02b5fcf, 32'h40493cad} /* (18, 4, 8) {real, imag} */,
  {32'hc0aba1c8, 32'h3fd55588} /* (18, 4, 7) {real, imag} */,
  {32'hc04c0c34, 32'hc0823adf} /* (18, 4, 6) {real, imag} */,
  {32'hc0983e56, 32'hbf5de85a} /* (18, 4, 5) {real, imag} */,
  {32'hc0381f22, 32'hbdc18960} /* (18, 4, 4) {real, imag} */,
  {32'h40145c55, 32'hc015449c} /* (18, 4, 3) {real, imag} */,
  {32'h408552d7, 32'hc0a40af9} /* (18, 4, 2) {real, imag} */,
  {32'h4037d6aa, 32'h3e3235c0} /* (18, 4, 1) {real, imag} */,
  {32'hbf35bab3, 32'h400af1fd} /* (18, 4, 0) {real, imag} */,
  {32'hbfe705a0, 32'h3f7c4474} /* (18, 3, 31) {real, imag} */,
  {32'h3ca0bf00, 32'h3fefdcca} /* (18, 3, 30) {real, imag} */,
  {32'hc091cd0f, 32'hc01cc722} /* (18, 3, 29) {real, imag} */,
  {32'h3fd47242, 32'hc0b4ea60} /* (18, 3, 28) {real, imag} */,
  {32'h40c546b0, 32'hc0ed28b9} /* (18, 3, 27) {real, imag} */,
  {32'hc0281d3b, 32'hc081bd98} /* (18, 3, 26) {real, imag} */,
  {32'hc02e18a0, 32'h4023119d} /* (18, 3, 25) {real, imag} */,
  {32'hc103af19, 32'h40dfce4a} /* (18, 3, 24) {real, imag} */,
  {32'hbfd7b9c8, 32'h401c6d05} /* (18, 3, 23) {real, imag} */,
  {32'h3f6cb1f0, 32'hc005b1fa} /* (18, 3, 22) {real, imag} */,
  {32'h3fffe660, 32'h3fad8706} /* (18, 3, 21) {real, imag} */,
  {32'hbe3da688, 32'h40e250fa} /* (18, 3, 20) {real, imag} */,
  {32'hbfd9278d, 32'hbfd4d684} /* (18, 3, 19) {real, imag} */,
  {32'h4007f2ae, 32'hc0af4ff6} /* (18, 3, 18) {real, imag} */,
  {32'h408d090b, 32'hc089360b} /* (18, 3, 17) {real, imag} */,
  {32'h40280f66, 32'h3fdb24b9} /* (18, 3, 16) {real, imag} */,
  {32'h4080c3bb, 32'h408c633a} /* (18, 3, 15) {real, imag} */,
  {32'h4078a63d, 32'hc050ce72} /* (18, 3, 14) {real, imag} */,
  {32'h3f62a3b3, 32'hc091e916} /* (18, 3, 13) {real, imag} */,
  {32'hbe8179d0, 32'hc05e91d3} /* (18, 3, 12) {real, imag} */,
  {32'hc09a6d0a, 32'h411a95e0} /* (18, 3, 11) {real, imag} */,
  {32'hbec1757a, 32'h40858872} /* (18, 3, 10) {real, imag} */,
  {32'hbf3bf588, 32'hc0ae58b0} /* (18, 3, 9) {real, imag} */,
  {32'hc0ec5858, 32'hc0f53b41} /* (18, 3, 8) {real, imag} */,
  {32'hc0dd116f, 32'hc0a8715d} /* (18, 3, 7) {real, imag} */,
  {32'h3f47eb44, 32'hc13d9610} /* (18, 3, 6) {real, imag} */,
  {32'hbf8af950, 32'hc0e6a587} /* (18, 3, 5) {real, imag} */,
  {32'hc01702b4, 32'hbfe3d1b0} /* (18, 3, 4) {real, imag} */,
  {32'hc09a44f1, 32'h3fa0a82f} /* (18, 3, 3) {real, imag} */,
  {32'hc04ff43e, 32'h40387820} /* (18, 3, 2) {real, imag} */,
  {32'hc0ba413e, 32'h3f79704d} /* (18, 3, 1) {real, imag} */,
  {32'hc020b1c6, 32'hbf90fe4d} /* (18, 3, 0) {real, imag} */,
  {32'h40979d81, 32'h4024eb8a} /* (18, 2, 31) {real, imag} */,
  {32'h405d553c, 32'h406b1990} /* (18, 2, 30) {real, imag} */,
  {32'h40f7bd56, 32'h410a23cf} /* (18, 2, 29) {real, imag} */,
  {32'h4024b965, 32'h40a31a63} /* (18, 2, 28) {real, imag} */,
  {32'h40a01a2a, 32'hc047e1ac} /* (18, 2, 27) {real, imag} */,
  {32'h40eae32b, 32'hc0093608} /* (18, 2, 26) {real, imag} */,
  {32'h410c7c08, 32'hc07bcd2e} /* (18, 2, 25) {real, imag} */,
  {32'h40ac43d2, 32'h3f43032c} /* (18, 2, 24) {real, imag} */,
  {32'h4101183a, 32'hc0692c38} /* (18, 2, 23) {real, imag} */,
  {32'h40db5b4a, 32'hbf4b4560} /* (18, 2, 22) {real, imag} */,
  {32'hbfab867a, 32'h4058e485} /* (18, 2, 21) {real, imag} */,
  {32'hc11711c2, 32'h402ef2e4} /* (18, 2, 20) {real, imag} */,
  {32'hc1121029, 32'hbdcd3200} /* (18, 2, 19) {real, imag} */,
  {32'hc13a6f4f, 32'hc0c0aa68} /* (18, 2, 18) {real, imag} */,
  {32'hc15f3868, 32'hc0bea741} /* (18, 2, 17) {real, imag} */,
  {32'hc11571bf, 32'hbfca2ee7} /* (18, 2, 16) {real, imag} */,
  {32'hc1396a8d, 32'hc0433bd6} /* (18, 2, 15) {real, imag} */,
  {32'hc0cfad30, 32'hc05fe77b} /* (18, 2, 14) {real, imag} */,
  {32'hc0d36ad2, 32'hc0415c66} /* (18, 2, 13) {real, imag} */,
  {32'hc1272a1e, 32'hc0671dd4} /* (18, 2, 12) {real, imag} */,
  {32'h3ff5c0e4, 32'hbf0820f8} /* (18, 2, 11) {real, imag} */,
  {32'h411d0f88, 32'h408a423d} /* (18, 2, 10) {real, imag} */,
  {32'h411421e1, 32'hbf9490e4} /* (18, 2, 9) {real, imag} */,
  {32'h40c59304, 32'hc067b1dd} /* (18, 2, 8) {real, imag} */,
  {32'h411fc822, 32'h405a954c} /* (18, 2, 7) {real, imag} */,
  {32'h410ebe17, 32'h401c3527} /* (18, 2, 6) {real, imag} */,
  {32'h402f9790, 32'h3f6c7dd1} /* (18, 2, 5) {real, imag} */,
  {32'h4110b3a0, 32'h40743598} /* (18, 2, 4) {real, imag} */,
  {32'h414fee47, 32'h401c4d47} /* (18, 2, 3) {real, imag} */,
  {32'h41120ab3, 32'hbfd3e80e} /* (18, 2, 2) {real, imag} */,
  {32'h410c3dbd, 32'hc0941bf0} /* (18, 2, 1) {real, imag} */,
  {32'h40a69e3e, 32'hc039368e} /* (18, 2, 0) {real, imag} */,
  {32'hc08c5fa0, 32'h3f549b1a} /* (18, 1, 31) {real, imag} */,
  {32'hc08bae99, 32'h401cc3fd} /* (18, 1, 30) {real, imag} */,
  {32'hc0a87a8f, 32'h3ece17f8} /* (18, 1, 29) {real, imag} */,
  {32'hc14c0ac2, 32'h3f3632fa} /* (18, 1, 28) {real, imag} */,
  {32'hc1449276, 32'hbe88b3a8} /* (18, 1, 27) {real, imag} */,
  {32'hc080cb28, 32'h3e8130ef} /* (18, 1, 26) {real, imag} */,
  {32'hbfff1568, 32'hc04ae72e} /* (18, 1, 25) {real, imag} */,
  {32'hc05ba158, 32'hbfcef8a2} /* (18, 1, 24) {real, imag} */,
  {32'hbfb0980c, 32'h3fb2590a} /* (18, 1, 23) {real, imag} */,
  {32'hc0bf26fc, 32'hc046a262} /* (18, 1, 22) {real, imag} */,
  {32'h3f9c24b1, 32'hbfdbbdba} /* (18, 1, 21) {real, imag} */,
  {32'h40cff88e, 32'h4039cddb} /* (18, 1, 20) {real, imag} */,
  {32'h3eeb96ec, 32'hbf54fcd6} /* (18, 1, 19) {real, imag} */,
  {32'h40204ed4, 32'h40b80500} /* (18, 1, 18) {real, imag} */,
  {32'h405b7434, 32'h412b1fc2} /* (18, 1, 17) {real, imag} */,
  {32'h408d8947, 32'h40a2a708} /* (18, 1, 16) {real, imag} */,
  {32'h40cef308, 32'hbfc74409} /* (18, 1, 15) {real, imag} */,
  {32'h41434d46, 32'h4095ce4c} /* (18, 1, 14) {real, imag} */,
  {32'h4076203c, 32'h40a6d05a} /* (18, 1, 13) {real, imag} */,
  {32'h40b8cd3b, 32'h4091fd1c} /* (18, 1, 12) {real, imag} */,
  {32'h40f27678, 32'h3eab64d8} /* (18, 1, 11) {real, imag} */,
  {32'h40293926, 32'hc0c96651} /* (18, 1, 10) {real, imag} */,
  {32'hbf2c01c0, 32'hc102dcf6} /* (18, 1, 9) {real, imag} */,
  {32'hc0822164, 32'hbfe38d7d} /* (18, 1, 8) {real, imag} */,
  {32'hc12e00d6, 32'hc0c06649} /* (18, 1, 7) {real, imag} */,
  {32'hc135093b, 32'hc10d3821} /* (18, 1, 6) {real, imag} */,
  {32'hc1215c51, 32'hc022e088} /* (18, 1, 5) {real, imag} */,
  {32'hc0ed2760, 32'h410a24ac} /* (18, 1, 4) {real, imag} */,
  {32'hc08c4d28, 32'h40654449} /* (18, 1, 3) {real, imag} */,
  {32'hc134afa2, 32'hc10b64fc} /* (18, 1, 2) {real, imag} */,
  {32'hc13bfcee, 32'hc05f8300} /* (18, 1, 1) {real, imag} */,
  {32'hc0c45a15, 32'h40892684} /* (18, 1, 0) {real, imag} */,
  {32'hc098bd2c, 32'hc0ad4398} /* (18, 0, 31) {real, imag} */,
  {32'hc08d8a12, 32'hc0a24fc8} /* (18, 0, 30) {real, imag} */,
  {32'h3f8cb3d4, 32'h3f010668} /* (18, 0, 29) {real, imag} */,
  {32'hc08d6ef6, 32'hbbb62c00} /* (18, 0, 28) {real, imag} */,
  {32'hc121c4ca, 32'hc056d0b0} /* (18, 0, 27) {real, imag} */,
  {32'hc11ef575, 32'h3e237ee0} /* (18, 0, 26) {real, imag} */,
  {32'hc0c35cce, 32'h40fe6c66} /* (18, 0, 25) {real, imag} */,
  {32'hc109798c, 32'h40b3c3c0} /* (18, 0, 24) {real, imag} */,
  {32'hc0b781b8, 32'hc09890ea} /* (18, 0, 23) {real, imag} */,
  {32'hc1024d50, 32'hc0c4a8e3} /* (18, 0, 22) {real, imag} */,
  {32'hc1168537, 32'hbfd737c7} /* (18, 0, 21) {real, imag} */,
  {32'hc109f02a, 32'hbfe22a37} /* (18, 0, 20) {real, imag} */,
  {32'h4080e756, 32'hc0d06d4a} /* (18, 0, 19) {real, imag} */,
  {32'h4100d0bd, 32'hc08572a2} /* (18, 0, 18) {real, imag} */,
  {32'h401ff3c6, 32'hc13428cf} /* (18, 0, 17) {real, imag} */,
  {32'hc01f2a42, 32'hc0db476d} /* (18, 0, 16) {real, imag} */,
  {32'h40b251d5, 32'hbf933a58} /* (18, 0, 15) {real, imag} */,
  {32'h40efde32, 32'h3faad4e4} /* (18, 0, 14) {real, imag} */,
  {32'h3fdd5a7b, 32'hc08bc4ee} /* (18, 0, 13) {real, imag} */,
  {32'hbeffb1ea, 32'hbfb7b12a} /* (18, 0, 12) {real, imag} */,
  {32'h40664050, 32'h40f2f4e6} /* (18, 0, 11) {real, imag} */,
  {32'hc02a294e, 32'h40a86c65} /* (18, 0, 10) {real, imag} */,
  {32'hc08ad9e9, 32'hc02a307b} /* (18, 0, 9) {real, imag} */,
  {32'h40438acc, 32'h3f9f485c} /* (18, 0, 8) {real, imag} */,
  {32'h40a30ad0, 32'hbf3c4170} /* (18, 0, 7) {real, imag} */,
  {32'h40b8554d, 32'hc0f86115} /* (18, 0, 6) {real, imag} */,
  {32'hbff31a12, 32'hc11487d9} /* (18, 0, 5) {real, imag} */,
  {32'hc0b6c8e7, 32'hbf103a80} /* (18, 0, 4) {real, imag} */,
  {32'hc02e1170, 32'h4004054b} /* (18, 0, 3) {real, imag} */,
  {32'h40247f40, 32'h408deed0} /* (18, 0, 2) {real, imag} */,
  {32'h3fcc09cc, 32'h40c8b91d} /* (18, 0, 1) {real, imag} */,
  {32'hbfef930a, 32'hc00f50c9} /* (18, 0, 0) {real, imag} */,
  {32'h3f9a032e, 32'hc0a0c161} /* (17, 31, 31) {real, imag} */,
  {32'h3fe788ca, 32'h3e6bd6d0} /* (17, 31, 30) {real, imag} */,
  {32'h4099584d, 32'hc013e274} /* (17, 31, 29) {real, imag} */,
  {32'h3c10e740, 32'hc03b0f80} /* (17, 31, 28) {real, imag} */,
  {32'hbf95d45a, 32'hbfa6ce18} /* (17, 31, 27) {real, imag} */,
  {32'h3fc0af44, 32'h3f05684e} /* (17, 31, 26) {real, imag} */,
  {32'h40e2c20c, 32'h3d7e4000} /* (17, 31, 25) {real, imag} */,
  {32'h40961ba2, 32'hc0036816} /* (17, 31, 24) {real, imag} */,
  {32'h40a4282c, 32'hbf885d2d} /* (17, 31, 23) {real, imag} */,
  {32'h40d4fd58, 32'h40367412} /* (17, 31, 22) {real, imag} */,
  {32'h4049a3d8, 32'h3fe4c358} /* (17, 31, 21) {real, imag} */,
  {32'hc0aa3a01, 32'h406256ac} /* (17, 31, 20) {real, imag} */,
  {32'hc0733ce9, 32'h3fce96b0} /* (17, 31, 19) {real, imag} */,
  {32'hc068650c, 32'hc06389d9} /* (17, 31, 18) {real, imag} */,
  {32'h3ef5ce78, 32'hc02dd660} /* (17, 31, 17) {real, imag} */,
  {32'hc0f781e4, 32'h40143dbd} /* (17, 31, 16) {real, imag} */,
  {32'hc106fbbf, 32'h4013a9e4} /* (17, 31, 15) {real, imag} */,
  {32'h3ea4159c, 32'h4041a8a5} /* (17, 31, 14) {real, imag} */,
  {32'hc07ca79b, 32'h3eb26530} /* (17, 31, 13) {real, imag} */,
  {32'hc117ad99, 32'hbe2b1dd0} /* (17, 31, 12) {real, imag} */,
  {32'hc01467d9, 32'hc0ac97d1} /* (17, 31, 11) {real, imag} */,
  {32'hbf818a18, 32'hc086b014} /* (17, 31, 10) {real, imag} */,
  {32'h40025238, 32'hc00e533e} /* (17, 31, 9) {real, imag} */,
  {32'h4066f728, 32'hc05d6837} /* (17, 31, 8) {real, imag} */,
  {32'h40889873, 32'hc0a3e4fb} /* (17, 31, 7) {real, imag} */,
  {32'h408abc38, 32'hc08af81e} /* (17, 31, 6) {real, imag} */,
  {32'h40cabcae, 32'hbfe66354} /* (17, 31, 5) {real, imag} */,
  {32'h40f20255, 32'hbf74d280} /* (17, 31, 4) {real, imag} */,
  {32'h4113b644, 32'hbea134a4} /* (17, 31, 3) {real, imag} */,
  {32'h3fc66294, 32'h40b5eea4} /* (17, 31, 2) {real, imag} */,
  {32'h4043f423, 32'hbfec663c} /* (17, 31, 1) {real, imag} */,
  {32'h40c5feaf, 32'hc06fd63c} /* (17, 31, 0) {real, imag} */,
  {32'hc07433bb, 32'hc05a4a52} /* (17, 30, 31) {real, imag} */,
  {32'hc0d79ac4, 32'hc0781171} /* (17, 30, 30) {real, imag} */,
  {32'hc051fc3a, 32'hbfac09aa} /* (17, 30, 29) {real, imag} */,
  {32'h4042880d, 32'h3eedbaa0} /* (17, 30, 28) {real, imag} */,
  {32'h40244cef, 32'hc049f53d} /* (17, 30, 27) {real, imag} */,
  {32'hc072c18c, 32'h407276ee} /* (17, 30, 26) {real, imag} */,
  {32'hc08ca429, 32'hbfd53ab2} /* (17, 30, 25) {real, imag} */,
  {32'hc00766dc, 32'h3f434aa4} /* (17, 30, 24) {real, imag} */,
  {32'h3fac5eff, 32'hc008cdc4} /* (17, 30, 23) {real, imag} */,
  {32'h3f5cb1db, 32'hc1151f42} /* (17, 30, 22) {real, imag} */,
  {32'hbf92a714, 32'hc08c301e} /* (17, 30, 21) {real, imag} */,
  {32'h3ff305d3, 32'hc0eee0e5} /* (17, 30, 20) {real, imag} */,
  {32'h40929904, 32'hc1479604} /* (17, 30, 19) {real, imag} */,
  {32'h402091a5, 32'hc0cb3681} /* (17, 30, 18) {real, imag} */,
  {32'h4066e5d4, 32'hc0363dfa} /* (17, 30, 17) {real, imag} */,
  {32'h3f1cc780, 32'h3e9dbce8} /* (17, 30, 16) {real, imag} */,
  {32'hbd5dcf00, 32'hbe0d41a0} /* (17, 30, 15) {real, imag} */,
  {32'h404f76ab, 32'h400a5eda} /* (17, 30, 14) {real, imag} */,
  {32'h409ca551, 32'h3e93aca0} /* (17, 30, 13) {real, imag} */,
  {32'h409fd23c, 32'hbdae0f08} /* (17, 30, 12) {real, imag} */,
  {32'h3f8d2b5b, 32'hbf2d7998} /* (17, 30, 11) {real, imag} */,
  {32'hc00c32b8, 32'hc0a1a6b4} /* (17, 30, 10) {real, imag} */,
  {32'hc0af581f, 32'hc0971c1e} /* (17, 30, 9) {real, imag} */,
  {32'h3e2726ae, 32'hc07fb0ad} /* (17, 30, 8) {real, imag} */,
  {32'h40cb01a4, 32'hc046091a} /* (17, 30, 7) {real, imag} */,
  {32'h41314660, 32'hbffaeab2} /* (17, 30, 6) {real, imag} */,
  {32'hbf22b2c6, 32'hc09d2842} /* (17, 30, 5) {real, imag} */,
  {32'hc1098f8c, 32'hc006982b} /* (17, 30, 4) {real, imag} */,
  {32'hc029be7d, 32'h40616bc9} /* (17, 30, 3) {real, imag} */,
  {32'h4068f356, 32'h40228c4d} /* (17, 30, 2) {real, imag} */,
  {32'hbed53280, 32'hbe9da236} /* (17, 30, 1) {real, imag} */,
  {32'hc055d10c, 32'h3fd585d2} /* (17, 30, 0) {real, imag} */,
  {32'h406a8a31, 32'h404c744c} /* (17, 29, 31) {real, imag} */,
  {32'h3fa8232c, 32'h3ff7b59a} /* (17, 29, 30) {real, imag} */,
  {32'hbf86b9cf, 32'h400f9fe9} /* (17, 29, 29) {real, imag} */,
  {32'h40882e98, 32'h3f997940} /* (17, 29, 28) {real, imag} */,
  {32'h40392b1e, 32'hbf7c135e} /* (17, 29, 27) {real, imag} */,
  {32'h3f984d58, 32'hbce0c700} /* (17, 29, 26) {real, imag} */,
  {32'h405924ca, 32'hc0bd82e6} /* (17, 29, 25) {real, imag} */,
  {32'h3e3b2450, 32'h3ede28ac} /* (17, 29, 24) {real, imag} */,
  {32'hc0fe8abe, 32'h3f4bb85f} /* (17, 29, 23) {real, imag} */,
  {32'hc0519e95, 32'hc0169ffe} /* (17, 29, 22) {real, imag} */,
  {32'hc04af965, 32'hbfd9eba5} /* (17, 29, 21) {real, imag} */,
  {32'hbfa39d54, 32'hbf7619aa} /* (17, 29, 20) {real, imag} */,
  {32'h40184158, 32'h3f88535f} /* (17, 29, 19) {real, imag} */,
  {32'hc0ba62f4, 32'hbf7fbad4} /* (17, 29, 18) {real, imag} */,
  {32'hc106bc2c, 32'h3e20f5f0} /* (17, 29, 17) {real, imag} */,
  {32'hc0a0e8b3, 32'h3ff4ceea} /* (17, 29, 16) {real, imag} */,
  {32'hc086a83d, 32'hbeb0266c} /* (17, 29, 15) {real, imag} */,
  {32'hc0b3ca90, 32'h402debac} /* (17, 29, 14) {real, imag} */,
  {32'hc009bf41, 32'h3fca59ba} /* (17, 29, 13) {real, imag} */,
  {32'hc001869c, 32'h3f744f50} /* (17, 29, 12) {real, imag} */,
  {32'h3fbc7ea4, 32'h40030070} /* (17, 29, 11) {real, imag} */,
  {32'hbfd45152, 32'hc0812732} /* (17, 29, 10) {real, imag} */,
  {32'h3fae1fa5, 32'hc0a9440f} /* (17, 29, 9) {real, imag} */,
  {32'hbe712490, 32'h3fefb02c} /* (17, 29, 8) {real, imag} */,
  {32'h4067af5a, 32'h4003436d} /* (17, 29, 7) {real, imag} */,
  {32'h408c03e6, 32'hc11e4f12} /* (17, 29, 6) {real, imag} */,
  {32'hbf6bf994, 32'hc0824545} /* (17, 29, 5) {real, imag} */,
  {32'hc0b545c0, 32'hbf969828} /* (17, 29, 4) {real, imag} */,
  {32'hc11c9d21, 32'hc03d8103} /* (17, 29, 3) {real, imag} */,
  {32'hc04884a1, 32'h3f5525c0} /* (17, 29, 2) {real, imag} */,
  {32'h3f198ea7, 32'hb9544000} /* (17, 29, 1) {real, imag} */,
  {32'h3f5990d4, 32'hbff1dbb4} /* (17, 29, 0) {real, imag} */,
  {32'hbfcc9198, 32'hbfa839ed} /* (17, 28, 31) {real, imag} */,
  {32'hc03ca732, 32'h3f47d370} /* (17, 28, 30) {real, imag} */,
  {32'hc0f5678c, 32'h40301c72} /* (17, 28, 29) {real, imag} */,
  {32'hc12bebc0, 32'hc05b64bf} /* (17, 28, 28) {real, imag} */,
  {32'hc0ffbe84, 32'hc090c6b8} /* (17, 28, 27) {real, imag} */,
  {32'hc0f9a70d, 32'hbfcbb321} /* (17, 28, 26) {real, imag} */,
  {32'hc0d0f4d6, 32'hbf8b8a53} /* (17, 28, 25) {real, imag} */,
  {32'h3ec1e784, 32'h3e12f928} /* (17, 28, 24) {real, imag} */,
  {32'h402ae51e, 32'hbeb71be4} /* (17, 28, 23) {real, imag} */,
  {32'hc0aca864, 32'hbfc6fe0b} /* (17, 28, 22) {real, imag} */,
  {32'hbf5c37e0, 32'h3f80f4ca} /* (17, 28, 21) {real, imag} */,
  {32'hc0b09bcc, 32'h409fb2dd} /* (17, 28, 20) {real, imag} */,
  {32'hc086bfc0, 32'h3ed74b30} /* (17, 28, 19) {real, imag} */,
  {32'hbee4e368, 32'hc103ea42} /* (17, 28, 18) {real, imag} */,
  {32'hc0adb24f, 32'hbda63a00} /* (17, 28, 17) {real, imag} */,
  {32'hc0b04dde, 32'h3f106504} /* (17, 28, 16) {real, imag} */,
  {32'h4001a0fd, 32'h3e972cd0} /* (17, 28, 15) {real, imag} */,
  {32'h40092ec6, 32'hbf62f8ce} /* (17, 28, 14) {real, imag} */,
  {32'hbe910238, 32'hc078f57b} /* (17, 28, 13) {real, imag} */,
  {32'hbfc74b5e, 32'hbf4e31d0} /* (17, 28, 12) {real, imag} */,
  {32'hc10410ac, 32'h40c8baf7} /* (17, 28, 11) {real, imag} */,
  {32'hc03f8a7a, 32'h406fdcc6} /* (17, 28, 10) {real, imag} */,
  {32'hc043a3fc, 32'hc027c865} /* (17, 28, 9) {real, imag} */,
  {32'h3dbfd870, 32'hc0925ad4} /* (17, 28, 8) {real, imag} */,
  {32'h4069d016, 32'hbf4bdf45} /* (17, 28, 7) {real, imag} */,
  {32'h40a062e0, 32'hbdc7b440} /* (17, 28, 6) {real, imag} */,
  {32'h40b20bd6, 32'h3fa128ae} /* (17, 28, 5) {real, imag} */,
  {32'h407996a0, 32'h3f08ffbc} /* (17, 28, 4) {real, imag} */,
  {32'hbf52fbd0, 32'hc0a6412c} /* (17, 28, 3) {real, imag} */,
  {32'h3f4f6ba3, 32'hc00ae050} /* (17, 28, 2) {real, imag} */,
  {32'hbed620a8, 32'h4068e8c6} /* (17, 28, 1) {real, imag} */,
  {32'h3ede6c10, 32'h402015a5} /* (17, 28, 0) {real, imag} */,
  {32'h405981d4, 32'hc0127b3f} /* (17, 27, 31) {real, imag} */,
  {32'h3f9095cd, 32'hc03fe7e6} /* (17, 27, 30) {real, imag} */,
  {32'hbe5cb1d6, 32'hc00caaca} /* (17, 27, 29) {real, imag} */,
  {32'hbfc00a05, 32'h40cb4e74} /* (17, 27, 28) {real, imag} */,
  {32'hbdf20ac0, 32'h40d9b5f1} /* (17, 27, 27) {real, imag} */,
  {32'h4096bdb4, 32'h40825c3e} /* (17, 27, 26) {real, imag} */,
  {32'h40658f95, 32'h3fd38362} /* (17, 27, 25) {real, imag} */,
  {32'h4006ab34, 32'h3f1b6470} /* (17, 27, 24) {real, imag} */,
  {32'h40032f07, 32'h4041fc2a} /* (17, 27, 23) {real, imag} */,
  {32'hc030425a, 32'h3f92a6e0} /* (17, 27, 22) {real, imag} */,
  {32'hc00d2f31, 32'h40043338} /* (17, 27, 21) {real, imag} */,
  {32'hc02b25fe, 32'h3fa9939a} /* (17, 27, 20) {real, imag} */,
  {32'hbf5b42b0, 32'hbfca6752} /* (17, 27, 19) {real, imag} */,
  {32'hc09fefab, 32'hbffea559} /* (17, 27, 18) {real, imag} */,
  {32'hc0380f8a, 32'h3fef2094} /* (17, 27, 17) {real, imag} */,
  {32'h3b9e5c00, 32'h408cb3f4} /* (17, 27, 16) {real, imag} */,
  {32'h40320bdc, 32'h4004fd7e} /* (17, 27, 15) {real, imag} */,
  {32'h3f93608c, 32'hbf910ac2} /* (17, 27, 14) {real, imag} */,
  {32'hc0d5d119, 32'hbfe96311} /* (17, 27, 13) {real, imag} */,
  {32'hc08d59de, 32'hc02ab7aa} /* (17, 27, 12) {real, imag} */,
  {32'h3ec47e5c, 32'hc03a9245} /* (17, 27, 11) {real, imag} */,
  {32'h40363fc2, 32'hc08a2fc2} /* (17, 27, 10) {real, imag} */,
  {32'h40ca8f7c, 32'hc031cf4e} /* (17, 27, 9) {real, imag} */,
  {32'h402135a6, 32'h40901e50} /* (17, 27, 8) {real, imag} */,
  {32'hc08a59cf, 32'h41158990} /* (17, 27, 7) {real, imag} */,
  {32'h3c199600, 32'h40ce1983} /* (17, 27, 6) {real, imag} */,
  {32'h402a936f, 32'h40935e9b} /* (17, 27, 5) {real, imag} */,
  {32'h3f8e8329, 32'h3f672f0f} /* (17, 27, 4) {real, imag} */,
  {32'hbf95cdc1, 32'hbff1f6ce} /* (17, 27, 3) {real, imag} */,
  {32'h3fb6a83c, 32'hbf32700d} /* (17, 27, 2) {real, imag} */,
  {32'h4111a54a, 32'hbee93e20} /* (17, 27, 1) {real, imag} */,
  {32'h40e31082, 32'hc0128246} /* (17, 27, 0) {real, imag} */,
  {32'hbf3af3d1, 32'hc0768bb4} /* (17, 26, 31) {real, imag} */,
  {32'h3f050d84, 32'hc0392c1c} /* (17, 26, 30) {real, imag} */,
  {32'hc030e07c, 32'h3f1ef2cf} /* (17, 26, 29) {real, imag} */,
  {32'hc10a36d3, 32'h403744c6} /* (17, 26, 28) {real, imag} */,
  {32'hc0d91c51, 32'h3f5c9045} /* (17, 26, 27) {real, imag} */,
  {32'h3f97061a, 32'hc0720308} /* (17, 26, 26) {real, imag} */,
  {32'h3ec224ce, 32'h3e66c5e8} /* (17, 26, 25) {real, imag} */,
  {32'hbe8a0a38, 32'h4001bf6a} /* (17, 26, 24) {real, imag} */,
  {32'h409b532e, 32'hc002391e} /* (17, 26, 23) {real, imag} */,
  {32'h403694aa, 32'h3f0fc4a6} /* (17, 26, 22) {real, imag} */,
  {32'hbf9d180b, 32'h40848158} /* (17, 26, 21) {real, imag} */,
  {32'hc02ac17e, 32'h3ff94442} /* (17, 26, 20) {real, imag} */,
  {32'h3fa20879, 32'hc05a7362} /* (17, 26, 19) {real, imag} */,
  {32'h40384287, 32'h3f51e55c} /* (17, 26, 18) {real, imag} */,
  {32'h3ff47789, 32'h40828f8d} /* (17, 26, 17) {real, imag} */,
  {32'h3f9556f1, 32'hbf8d4df0} /* (17, 26, 16) {real, imag} */,
  {32'h3f953be1, 32'hc0a041cb} /* (17, 26, 15) {real, imag} */,
  {32'hbf0d04d2, 32'h3fea4334} /* (17, 26, 14) {real, imag} */,
  {32'hc094d251, 32'h406dc86e} /* (17, 26, 13) {real, imag} */,
  {32'hbe8e99d0, 32'h4072fb27} /* (17, 26, 12) {real, imag} */,
  {32'hbf26f164, 32'h402584da} /* (17, 26, 11) {real, imag} */,
  {32'h3f979432, 32'hc0410422} /* (17, 26, 10) {real, imag} */,
  {32'h3fa2bcdf, 32'hbffde740} /* (17, 26, 9) {real, imag} */,
  {32'hc0eef570, 32'h407ef9f8} /* (17, 26, 8) {real, imag} */,
  {32'hbfd57546, 32'h405b1156} /* (17, 26, 7) {real, imag} */,
  {32'h3ed9f7dc, 32'hbf98a53a} /* (17, 26, 6) {real, imag} */,
  {32'h3f7ebf58, 32'hbf0201a2} /* (17, 26, 5) {real, imag} */,
  {32'hc07c96c8, 32'hbfc470a2} /* (17, 26, 4) {real, imag} */,
  {32'hc029984d, 32'hc0b0735c} /* (17, 26, 3) {real, imag} */,
  {32'h3f32b3b8, 32'hbea46940} /* (17, 26, 2) {real, imag} */,
  {32'h3f86dd95, 32'h405d4f2a} /* (17, 26, 1) {real, imag} */,
  {32'h3fe21366, 32'hbdc930a0} /* (17, 26, 0) {real, imag} */,
  {32'h3f192575, 32'hbc05b140} /* (17, 25, 31) {real, imag} */,
  {32'h4069471e, 32'hbf549dc3} /* (17, 25, 30) {real, imag} */,
  {32'hbf7a5d0c, 32'hc074848f} /* (17, 25, 29) {real, imag} */,
  {32'hc03c5907, 32'hbf04c88b} /* (17, 25, 28) {real, imag} */,
  {32'hbf6a9a36, 32'hc05a2a0e} /* (17, 25, 27) {real, imag} */,
  {32'hbf8c5ec4, 32'hc03dea30} /* (17, 25, 26) {real, imag} */,
  {32'hbf056eb8, 32'h4051ee0e} /* (17, 25, 25) {real, imag} */,
  {32'hbfc93b28, 32'h404847ca} /* (17, 25, 24) {real, imag} */,
  {32'hc07b2fb2, 32'h4032f59d} /* (17, 25, 23) {real, imag} */,
  {32'hc0ba2acc, 32'h404fd2cc} /* (17, 25, 22) {real, imag} */,
  {32'hc0207622, 32'h401140a8} /* (17, 25, 21) {real, imag} */,
  {32'h3f491ce2, 32'hbf853aac} /* (17, 25, 20) {real, imag} */,
  {32'h404a65c6, 32'h402c72a8} /* (17, 25, 19) {real, imag} */,
  {32'h40cdca1c, 32'h3f94fcbe} /* (17, 25, 18) {real, imag} */,
  {32'h40b2527a, 32'h3f3dc838} /* (17, 25, 17) {real, imag} */,
  {32'hc01bfead, 32'h4022de14} /* (17, 25, 16) {real, imag} */,
  {32'hbfcb231a, 32'hbf0f1dee} /* (17, 25, 15) {real, imag} */,
  {32'h4056cec1, 32'hbf4c15c3} /* (17, 25, 14) {real, imag} */,
  {32'h408ffb28, 32'h40582141} /* (17, 25, 13) {real, imag} */,
  {32'h3f6e1cfa, 32'hbe1316b0} /* (17, 25, 12) {real, imag} */,
  {32'hc001bca2, 32'h3d35c780} /* (17, 25, 11) {real, imag} */,
  {32'hbf90e46d, 32'h3ff0d136} /* (17, 25, 10) {real, imag} */,
  {32'hbffe7d39, 32'h3fda1ea7} /* (17, 25, 9) {real, imag} */,
  {32'h3fb6e436, 32'h3ebb36f4} /* (17, 25, 8) {real, imag} */,
  {32'h3ef7f460, 32'hbff473d4} /* (17, 25, 7) {real, imag} */,
  {32'hc065711a, 32'h3dede720} /* (17, 25, 6) {real, imag} */,
  {32'hc0b10ae1, 32'hc057409b} /* (17, 25, 5) {real, imag} */,
  {32'hc00255cd, 32'hc0b5c258} /* (17, 25, 4) {real, imag} */,
  {32'h4070e4bc, 32'hc08828d2} /* (17, 25, 3) {real, imag} */,
  {32'h401d40b7, 32'hc0db89ad} /* (17, 25, 2) {real, imag} */,
  {32'h3fa11580, 32'hc0ce26a4} /* (17, 25, 1) {real, imag} */,
  {32'h3fd5854e, 32'hc02d83fa} /* (17, 25, 0) {real, imag} */,
  {32'hbff6a385, 32'hbee759bc} /* (17, 24, 31) {real, imag} */,
  {32'hc036bad0, 32'h3fff8c4e} /* (17, 24, 30) {real, imag} */,
  {32'hc0b9b3ea, 32'h3f0a882e} /* (17, 24, 29) {real, imag} */,
  {32'hc0ac274a, 32'hbe9e5f04} /* (17, 24, 28) {real, imag} */,
  {32'hbef5bbf6, 32'h3fa89096} /* (17, 24, 27) {real, imag} */,
  {32'h3fef446e, 32'hc0c1c7f2} /* (17, 24, 26) {real, imag} */,
  {32'hbf3fa50e, 32'hc0b60f4a} /* (17, 24, 25) {real, imag} */,
  {32'hc028f919, 32'hc02f724f} /* (17, 24, 24) {real, imag} */,
  {32'h3e8d6cec, 32'h3f1c739f} /* (17, 24, 23) {real, imag} */,
  {32'h3cb15580, 32'hbeae190e} /* (17, 24, 22) {real, imag} */,
  {32'hc01dae40, 32'hbfb36e9c} /* (17, 24, 21) {real, imag} */,
  {32'hbfce8eb6, 32'h3f1f7df4} /* (17, 24, 20) {real, imag} */,
  {32'h3eb81c2c, 32'hbfbd6e85} /* (17, 24, 19) {real, imag} */,
  {32'h405a36ec, 32'hc007625a} /* (17, 24, 18) {real, imag} */,
  {32'h3fde17d2, 32'h3f9f4804} /* (17, 24, 17) {real, imag} */,
  {32'h40590825, 32'hbf14510c} /* (17, 24, 16) {real, imag} */,
  {32'hbfedec5d, 32'hbee95a42} /* (17, 24, 15) {real, imag} */,
  {32'hc0d819f8, 32'h3ef76d92} /* (17, 24, 14) {real, imag} */,
  {32'hc09846aa, 32'hbf5d26fc} /* (17, 24, 13) {real, imag} */,
  {32'h3f503e34, 32'h3f6c50f6} /* (17, 24, 12) {real, imag} */,
  {32'h3ea44006, 32'h3fe9a8d1} /* (17, 24, 11) {real, imag} */,
  {32'h3d367e50, 32'hbf54db9c} /* (17, 24, 10) {real, imag} */,
  {32'h3d189e00, 32'h400afc48} /* (17, 24, 9) {real, imag} */,
  {32'h3fbaf0f9, 32'h3e160acc} /* (17, 24, 8) {real, imag} */,
  {32'h403309f6, 32'h3ef66b48} /* (17, 24, 7) {real, imag} */,
  {32'h3f141411, 32'h3fa282d0} /* (17, 24, 6) {real, imag} */,
  {32'hc0d59496, 32'h400645e2} /* (17, 24, 5) {real, imag} */,
  {32'hc0f7aea0, 32'h3fcdc95e} /* (17, 24, 4) {real, imag} */,
  {32'hbfe40a3f, 32'h3f12e90c} /* (17, 24, 3) {real, imag} */,
  {32'h3eede3d4, 32'h400f200f} /* (17, 24, 2) {real, imag} */,
  {32'hbf237d79, 32'h404d3236} /* (17, 24, 1) {real, imag} */,
  {32'h3e93f996, 32'hbfae3386} /* (17, 24, 0) {real, imag} */,
  {32'h3fd6cb8a, 32'h3ff80035} /* (17, 23, 31) {real, imag} */,
  {32'hbf04c9ca, 32'h3f5f3dbf} /* (17, 23, 30) {real, imag} */,
  {32'hbf1d92b2, 32'hbf255e2c} /* (17, 23, 29) {real, imag} */,
  {32'hbfe322cd, 32'hbd8af380} /* (17, 23, 28) {real, imag} */,
  {32'hbf80d7a4, 32'hbfe6a58c} /* (17, 23, 27) {real, imag} */,
  {32'h400941ba, 32'h3f7ebc86} /* (17, 23, 26) {real, imag} */,
  {32'h409009a2, 32'hbf85504b} /* (17, 23, 25) {real, imag} */,
  {32'hc02ea66e, 32'hbfba6fbd} /* (17, 23, 24) {real, imag} */,
  {32'hc082c316, 32'hbdcf06d0} /* (17, 23, 23) {real, imag} */,
  {32'h4043cb24, 32'h3f7aa716} /* (17, 23, 22) {real, imag} */,
  {32'h3f62f9e4, 32'hbfcbdaee} /* (17, 23, 21) {real, imag} */,
  {32'h3de01fa0, 32'h3f6fb2cc} /* (17, 23, 20) {real, imag} */,
  {32'h3fbcd752, 32'h408314f4} /* (17, 23, 19) {real, imag} */,
  {32'hbf1eb988, 32'hbdc554b0} /* (17, 23, 18) {real, imag} */,
  {32'hc01d53d6, 32'h40157e98} /* (17, 23, 17) {real, imag} */,
  {32'hbfaeeb6e, 32'h4048c8b3} /* (17, 23, 16) {real, imag} */,
  {32'hbf09fbf4, 32'h3f938b06} /* (17, 23, 15) {real, imag} */,
  {32'h3fbbb14e, 32'h3f490ffd} /* (17, 23, 14) {real, imag} */,
  {32'h4024ba33, 32'h400bc75c} /* (17, 23, 13) {real, imag} */,
  {32'hc03c74c6, 32'hbf1274cb} /* (17, 23, 12) {real, imag} */,
  {32'hc06a62a8, 32'hc08063b7} /* (17, 23, 11) {real, imag} */,
  {32'h4040c9be, 32'hbfc1ecae} /* (17, 23, 10) {real, imag} */,
  {32'h3fc72d21, 32'h403312e8} /* (17, 23, 9) {real, imag} */,
  {32'hc09ce176, 32'h3fb38af2} /* (17, 23, 8) {real, imag} */,
  {32'h3d9c5f40, 32'hbfe345a4} /* (17, 23, 7) {real, imag} */,
  {32'h401997a5, 32'hbf8af1dc} /* (17, 23, 6) {real, imag} */,
  {32'hbede7f34, 32'hc09af21f} /* (17, 23, 5) {real, imag} */,
  {32'h3f8c409d, 32'hc07f7990} /* (17, 23, 4) {real, imag} */,
  {32'h3fef565b, 32'hbecd5b5c} /* (17, 23, 3) {real, imag} */,
  {32'h3f087d10, 32'h3f23afcc} /* (17, 23, 2) {real, imag} */,
  {32'h40408bf6, 32'hbdc38850} /* (17, 23, 1) {real, imag} */,
  {32'h3fc5db50, 32'hbde924a0} /* (17, 23, 0) {real, imag} */,
  {32'h3fcec51e, 32'hbf6277fd} /* (17, 22, 31) {real, imag} */,
  {32'hbd8cdba0, 32'hbeb515d8} /* (17, 22, 30) {real, imag} */,
  {32'hc00c761e, 32'hbe850f26} /* (17, 22, 29) {real, imag} */,
  {32'h3c3c1380, 32'h3ea85f84} /* (17, 22, 28) {real, imag} */,
  {32'h3eb27024, 32'hc0054bcb} /* (17, 22, 27) {real, imag} */,
  {32'hbf468c08, 32'hc06b8bc8} /* (17, 22, 26) {real, imag} */,
  {32'hbf916c7a, 32'hbebe1070} /* (17, 22, 25) {real, imag} */,
  {32'hc035c158, 32'hbfe52e26} /* (17, 22, 24) {real, imag} */,
  {32'hc09808ac, 32'hc00ed8fb} /* (17, 22, 23) {real, imag} */,
  {32'h3f468b38, 32'h3f9a5ca5} /* (17, 22, 22) {real, imag} */,
  {32'h403d05aa, 32'h3f2488d0} /* (17, 22, 21) {real, imag} */,
  {32'hbf2891c2, 32'h3f84b00d} /* (17, 22, 20) {real, imag} */,
  {32'hc03e9396, 32'h401ffb10} /* (17, 22, 19) {real, imag} */,
  {32'h3f0ca939, 32'h40790c4d} /* (17, 22, 18) {real, imag} */,
  {32'h3ed7c7f1, 32'h3e6328d0} /* (17, 22, 17) {real, imag} */,
  {32'hbea92e2c, 32'hc038e2bc} /* (17, 22, 16) {real, imag} */,
  {32'h3fcac17d, 32'h3f32335c} /* (17, 22, 15) {real, imag} */,
  {32'h400097d4, 32'h400701db} /* (17, 22, 14) {real, imag} */,
  {32'hbcdf8840, 32'h3e61c2b8} /* (17, 22, 13) {real, imag} */,
  {32'hbe93b5a0, 32'h3f86f9b0} /* (17, 22, 12) {real, imag} */,
  {32'hbfb416be, 32'hbeba1374} /* (17, 22, 11) {real, imag} */,
  {32'hbf9c3a81, 32'h3ed8e2ae} /* (17, 22, 10) {real, imag} */,
  {32'hc02a7e5f, 32'h3f9f598f} /* (17, 22, 9) {real, imag} */,
  {32'h3f02f064, 32'hbef02d98} /* (17, 22, 8) {real, imag} */,
  {32'hbcdb4b00, 32'hbf98852e} /* (17, 22, 7) {real, imag} */,
  {32'hbe430008, 32'hbfa85cf7} /* (17, 22, 6) {real, imag} */,
  {32'hbed04f9c, 32'hbe57fd04} /* (17, 22, 5) {real, imag} */,
  {32'hc01709ae, 32'h3ff0a2bc} /* (17, 22, 4) {real, imag} */,
  {32'h3f7ff9fa, 32'h3ff4fea6} /* (17, 22, 3) {real, imag} */,
  {32'h3f036684, 32'h3f7703d8} /* (17, 22, 2) {real, imag} */,
  {32'hbf471b96, 32'hbf30f4c7} /* (17, 22, 1) {real, imag} */,
  {32'hbeca6dcb, 32'hbf78ab22} /* (17, 22, 0) {real, imag} */,
  {32'hbee9398a, 32'h3f95b987} /* (17, 21, 31) {real, imag} */,
  {32'hbea00e82, 32'hbeb69e66} /* (17, 21, 30) {real, imag} */,
  {32'hbfacd0de, 32'hc01d298b} /* (17, 21, 29) {real, imag} */,
  {32'h3f25dc9e, 32'hbf7c7746} /* (17, 21, 28) {real, imag} */,
  {32'h3fb633d4, 32'hc01127ac} /* (17, 21, 27) {real, imag} */,
  {32'h3fcf5dfc, 32'hbf334f29} /* (17, 21, 26) {real, imag} */,
  {32'h3ea968c8, 32'h400d5e55} /* (17, 21, 25) {real, imag} */,
  {32'hc0037087, 32'h401f34d3} /* (17, 21, 24) {real, imag} */,
  {32'hbf682d50, 32'hbe6b8e88} /* (17, 21, 23) {real, imag} */,
  {32'h3e9856a0, 32'hbf73c136} /* (17, 21, 22) {real, imag} */,
  {32'h3f55ba64, 32'hbf700e0c} /* (17, 21, 21) {real, imag} */,
  {32'hbf6442e2, 32'h3d50cdc0} /* (17, 21, 20) {real, imag} */,
  {32'hbf9e38bc, 32'hbe984dd6} /* (17, 21, 19) {real, imag} */,
  {32'h3fc2cbc2, 32'h3d683310} /* (17, 21, 18) {real, imag} */,
  {32'hbfbb0d55, 32'h3fa635a4} /* (17, 21, 17) {real, imag} */,
  {32'hc01aa0ce, 32'h3f60621e} /* (17, 21, 16) {real, imag} */,
  {32'hbf8603af, 32'hbe090788} /* (17, 21, 15) {real, imag} */,
  {32'h3fa73f2e, 32'h3f96d8fa} /* (17, 21, 14) {real, imag} */,
  {32'h4026fd1e, 32'h3dc00c68} /* (17, 21, 13) {real, imag} */,
  {32'h3f4ce30c, 32'hbeb8870c} /* (17, 21, 12) {real, imag} */,
  {32'h3ed6e7c6, 32'hbfb6bb54} /* (17, 21, 11) {real, imag} */,
  {32'h3fd5f291, 32'hbf827364} /* (17, 21, 10) {real, imag} */,
  {32'h3eef3660, 32'h3f0e0a50} /* (17, 21, 9) {real, imag} */,
  {32'hbe98ecc6, 32'hbff1adb1} /* (17, 21, 8) {real, imag} */,
  {32'hc0373108, 32'hc02cac5c} /* (17, 21, 7) {real, imag} */,
  {32'hbf9ddf9e, 32'h3f0ea4a0} /* (17, 21, 6) {real, imag} */,
  {32'h401c0f43, 32'hbf4316b0} /* (17, 21, 5) {real, imag} */,
  {32'h3fa09724, 32'hbf3e74cc} /* (17, 21, 4) {real, imag} */,
  {32'hbf23f1ce, 32'hbff70550} /* (17, 21, 3) {real, imag} */,
  {32'h40045981, 32'hbf9c2db5} /* (17, 21, 2) {real, imag} */,
  {32'h4012fd8b, 32'hbfefc642} /* (17, 21, 1) {real, imag} */,
  {32'h3f84727c, 32'hbece57b4} /* (17, 21, 0) {real, imag} */,
  {32'h3fa9455e, 32'hbf42b376} /* (17, 20, 31) {real, imag} */,
  {32'h3e24b9a8, 32'hbf858560} /* (17, 20, 30) {real, imag} */,
  {32'h3f074f86, 32'hbe1b4820} /* (17, 20, 29) {real, imag} */,
  {32'h3ef10fb4, 32'hbf1598b0} /* (17, 20, 28) {real, imag} */,
  {32'h3d4c5810, 32'h3f80d412} /* (17, 20, 27) {real, imag} */,
  {32'h3f0bd5cc, 32'hbed82108} /* (17, 20, 26) {real, imag} */,
  {32'hbfcd4e72, 32'hc037b2e0} /* (17, 20, 25) {real, imag} */,
  {32'hbfdb866e, 32'hc0353bb0} /* (17, 20, 24) {real, imag} */,
  {32'hc062ac14, 32'hbfa83eab} /* (17, 20, 23) {real, imag} */,
  {32'hc02b8abc, 32'hbf22e281} /* (17, 20, 22) {real, imag} */,
  {32'h3e586b60, 32'hbfbd5002} /* (17, 20, 21) {real, imag} */,
  {32'h3f2ce89a, 32'hbf1753d9} /* (17, 20, 20) {real, imag} */,
  {32'hbff1116b, 32'h3f5f771c} /* (17, 20, 19) {real, imag} */,
  {32'hbfa05422, 32'hbed142e4} /* (17, 20, 18) {real, imag} */,
  {32'hbe575820, 32'hbfb1f056} /* (17, 20, 17) {real, imag} */,
  {32'hbefa70b8, 32'hbf2b6ae2} /* (17, 20, 16) {real, imag} */,
  {32'hc000a510, 32'hbed436d4} /* (17, 20, 15) {real, imag} */,
  {32'hc0462a76, 32'h3f9231f6} /* (17, 20, 14) {real, imag} */,
  {32'hbf2be504, 32'hbebe0e9a} /* (17, 20, 13) {real, imag} */,
  {32'hc010a6c6, 32'hbfb87e56} /* (17, 20, 12) {real, imag} */,
  {32'hbfb35c81, 32'h3f1c4b04} /* (17, 20, 11) {real, imag} */,
  {32'hbf3d16ea, 32'h3f83c112} /* (17, 20, 10) {real, imag} */,
  {32'hbfca6f3c, 32'h3f1c966a} /* (17, 20, 9) {real, imag} */,
  {32'hbf8c8fca, 32'h3f99548c} /* (17, 20, 8) {real, imag} */,
  {32'hbdfff968, 32'h3f28e6aa} /* (17, 20, 7) {real, imag} */,
  {32'hbf0cddb3, 32'hbfea40a4} /* (17, 20, 6) {real, imag} */,
  {32'h3e29085c, 32'hbfd17891} /* (17, 20, 5) {real, imag} */,
  {32'hbb63c800, 32'hbf29847c} /* (17, 20, 4) {real, imag} */,
  {32'h3f3bef80, 32'h3de3ee70} /* (17, 20, 3) {real, imag} */,
  {32'h3f9cd11a, 32'h3f0e2d66} /* (17, 20, 2) {real, imag} */,
  {32'h4011c598, 32'h401f4626} /* (17, 20, 1) {real, imag} */,
  {32'h3fc3ce5f, 32'h3de74d4c} /* (17, 20, 0) {real, imag} */,
  {32'hbf2461ea, 32'h3f4bda3c} /* (17, 19, 31) {real, imag} */,
  {32'hbf7bbb06, 32'hbfef2e92} /* (17, 19, 30) {real, imag} */,
  {32'hbf8d1508, 32'hbff13264} /* (17, 19, 29) {real, imag} */,
  {32'hbdc9c570, 32'hbfdd27bf} /* (17, 19, 28) {real, imag} */,
  {32'hbf3db602, 32'hbfbe52dc} /* (17, 19, 27) {real, imag} */,
  {32'h3fb7fcea, 32'hbf2ceb86} /* (17, 19, 26) {real, imag} */,
  {32'h3f81ef19, 32'hbf686ba7} /* (17, 19, 25) {real, imag} */,
  {32'h3f925812, 32'hbfdd4d2a} /* (17, 19, 24) {real, imag} */,
  {32'h3edee60c, 32'hbf3162df} /* (17, 19, 23) {real, imag} */,
  {32'h3ec4daa2, 32'h3f336366} /* (17, 19, 22) {real, imag} */,
  {32'hbddf5ab8, 32'h3f8dc51d} /* (17, 19, 21) {real, imag} */,
  {32'hbf3f04f4, 32'h3f7f6a7b} /* (17, 19, 20) {real, imag} */,
  {32'h3b537500, 32'h3e84df96} /* (17, 19, 19) {real, imag} */,
  {32'h3f358ade, 32'h3ef136ce} /* (17, 19, 18) {real, imag} */,
  {32'h3ecc169c, 32'h402fd4f7} /* (17, 19, 17) {real, imag} */,
  {32'h3ed3e244, 32'hbef55428} /* (17, 19, 16) {real, imag} */,
  {32'h3ed93614, 32'hbf8159ad} /* (17, 19, 15) {real, imag} */,
  {32'hbf6075d9, 32'hbe31ef7c} /* (17, 19, 14) {real, imag} */,
  {32'hbf0add2c, 32'hbfd596c8} /* (17, 19, 13) {real, imag} */,
  {32'h3ff1a21e, 32'hc00e6cee} /* (17, 19, 12) {real, imag} */,
  {32'h40420b0a, 32'hbf205f31} /* (17, 19, 11) {real, imag} */,
  {32'h3fc8617c, 32'h3fbfaf37} /* (17, 19, 10) {real, imag} */,
  {32'h4006ecba, 32'hbf3b5a84} /* (17, 19, 9) {real, imag} */,
  {32'h3ed4c804, 32'hbf7cb1bf} /* (17, 19, 8) {real, imag} */,
  {32'h3f4b17af, 32'hbf5a9c48} /* (17, 19, 7) {real, imag} */,
  {32'h3f6ca6e8, 32'h3f87b434} /* (17, 19, 6) {real, imag} */,
  {32'hbf8d0d84, 32'hbf85cee0} /* (17, 19, 5) {real, imag} */,
  {32'hbfc1294b, 32'hbf1f24be} /* (17, 19, 4) {real, imag} */,
  {32'hc027ae62, 32'h3f59045f} /* (17, 19, 3) {real, imag} */,
  {32'hbf7dc69c, 32'h3f154990} /* (17, 19, 2) {real, imag} */,
  {32'hbef6f7c6, 32'h3f57c278} /* (17, 19, 1) {real, imag} */,
  {32'hbfb6b6b6, 32'h3f29436f} /* (17, 19, 0) {real, imag} */,
  {32'hbdb9c648, 32'h3f0469ad} /* (17, 18, 31) {real, imag} */,
  {32'hbf4fa73a, 32'hbf474eea} /* (17, 18, 30) {real, imag} */,
  {32'hbe804c0c, 32'hbff9ff4e} /* (17, 18, 29) {real, imag} */,
  {32'h3e58b92a, 32'hbfc6e8c4} /* (17, 18, 28) {real, imag} */,
  {32'hbd844a20, 32'h3f6cc554} /* (17, 18, 27) {real, imag} */,
  {32'h3f01877c, 32'h40291e64} /* (17, 18, 26) {real, imag} */,
  {32'h400f71e0, 32'h3f39e4c7} /* (17, 18, 25) {real, imag} */,
  {32'h3fd41f54, 32'h3fc9df0e} /* (17, 18, 24) {real, imag} */,
  {32'hbf93fcd2, 32'h3fca228e} /* (17, 18, 23) {real, imag} */,
  {32'hbe34149c, 32'h3fa80060} /* (17, 18, 22) {real, imag} */,
  {32'h3fb1ddd8, 32'h3fb9a651} /* (17, 18, 21) {real, imag} */,
  {32'h3d8949c8, 32'h3f760f95} /* (17, 18, 20) {real, imag} */,
  {32'h3eca3144, 32'h3ef31b30} /* (17, 18, 19) {real, imag} */,
  {32'h3f5346cc, 32'h3c9a5340} /* (17, 18, 18) {real, imag} */,
  {32'h3f8e1ed2, 32'hbf598f10} /* (17, 18, 17) {real, imag} */,
  {32'hbeb506f0, 32'hbf73160c} /* (17, 18, 16) {real, imag} */,
  {32'hbf0cbf3f, 32'h3e519a78} /* (17, 18, 15) {real, imag} */,
  {32'hbe5d6dac, 32'h3f923702} /* (17, 18, 14) {real, imag} */,
  {32'hbf3855bf, 32'h4000860a} /* (17, 18, 13) {real, imag} */,
  {32'hbf603533, 32'h3fa426e2} /* (17, 18, 12) {real, imag} */,
  {32'hbf0f5a74, 32'hbf511110} /* (17, 18, 11) {real, imag} */,
  {32'h3f4b0c08, 32'hbcb896c0} /* (17, 18, 10) {real, imag} */,
  {32'h3fb45846, 32'hbe9517dc} /* (17, 18, 9) {real, imag} */,
  {32'h3f65af8a, 32'h3f91a446} /* (17, 18, 8) {real, imag} */,
  {32'h3f97ea3b, 32'h3efead20} /* (17, 18, 7) {real, imag} */,
  {32'h3f1eb8d7, 32'h3fb6f7ac} /* (17, 18, 6) {real, imag} */,
  {32'h3f5fe41e, 32'h3fa2cac0} /* (17, 18, 5) {real, imag} */,
  {32'h3fa8b982, 32'h3f26a49e} /* (17, 18, 4) {real, imag} */,
  {32'h3fbf065a, 32'hbee8ce38} /* (17, 18, 3) {real, imag} */,
  {32'h3f5982b6, 32'h3f2f4ad9} /* (17, 18, 2) {real, imag} */,
  {32'h3dddde80, 32'h3efad5ed} /* (17, 18, 1) {real, imag} */,
  {32'hbed02f7c, 32'h3f81ded0} /* (17, 18, 0) {real, imag} */,
  {32'hbd2921c0, 32'hbe149060} /* (17, 17, 31) {real, imag} */,
  {32'hbf6e3183, 32'hbec98d54} /* (17, 17, 30) {real, imag} */,
  {32'hbf01a505, 32'h3cb9c2c0} /* (17, 17, 29) {real, imag} */,
  {32'h3ea16f5e, 32'hbc39bf60} /* (17, 17, 28) {real, imag} */,
  {32'h3e1ef340, 32'hbf41bff3} /* (17, 17, 27) {real, imag} */,
  {32'h3f017bf8, 32'hbeac34d1} /* (17, 17, 26) {real, imag} */,
  {32'h3fa9657a, 32'h3f8ad11e} /* (17, 17, 25) {real, imag} */,
  {32'h3efb8012, 32'h3fc07052} /* (17, 17, 24) {real, imag} */,
  {32'h3e9b9f3e, 32'h3e30f2c0} /* (17, 17, 23) {real, imag} */,
  {32'h3e1c7760, 32'hbf21a73e} /* (17, 17, 22) {real, imag} */,
  {32'h3f486d36, 32'hbe567628} /* (17, 17, 21) {real, imag} */,
  {32'h3ebb9eaa, 32'h3f361a90} /* (17, 17, 20) {real, imag} */,
  {32'h3f9a5404, 32'h3f1b443f} /* (17, 17, 19) {real, imag} */,
  {32'hbf972612, 32'h3d834560} /* (17, 17, 18) {real, imag} */,
  {32'hbff9fdce, 32'hbf4e051a} /* (17, 17, 17) {real, imag} */,
  {32'h3e2a122c, 32'h3dae4008} /* (17, 17, 16) {real, imag} */,
  {32'h3f233a10, 32'h3f5eaa0c} /* (17, 17, 15) {real, imag} */,
  {32'h3f732926, 32'h3e4e3a08} /* (17, 17, 14) {real, imag} */,
  {32'h3ebeaddc, 32'hbd94faf0} /* (17, 17, 13) {real, imag} */,
  {32'hbf54df00, 32'h3ee2d03c} /* (17, 17, 12) {real, imag} */,
  {32'hbf70ba94, 32'hbf11a536} /* (17, 17, 11) {real, imag} */,
  {32'h3deb45c0, 32'hbf70b9f4} /* (17, 17, 10) {real, imag} */,
  {32'hbf1cacac, 32'h3f549635} /* (17, 17, 9) {real, imag} */,
  {32'h3eca1d14, 32'h3f89d223} /* (17, 17, 8) {real, imag} */,
  {32'hbea6df18, 32'h3df8c2e0} /* (17, 17, 7) {real, imag} */,
  {32'hbf19dfc5, 32'h3e979d1c} /* (17, 17, 6) {real, imag} */,
  {32'h3e259a30, 32'hbd573ad0} /* (17, 17, 5) {real, imag} */,
  {32'hbfc5cdeb, 32'hbe1c019c} /* (17, 17, 4) {real, imag} */,
  {32'hbfa71340, 32'h3eb73e4c} /* (17, 17, 3) {real, imag} */,
  {32'h3e32fee8, 32'h3f4f913a} /* (17, 17, 2) {real, imag} */,
  {32'hbe92bf06, 32'h3de7f260} /* (17, 17, 1) {real, imag} */,
  {32'h3f72922e, 32'hbf89ba0a} /* (17, 17, 0) {real, imag} */,
  {32'h3f49104c, 32'h3f6420d0} /* (17, 16, 31) {real, imag} */,
  {32'h3ea25bf8, 32'h3fb4f2ce} /* (17, 16, 30) {real, imag} */,
  {32'h3f0abdbe, 32'h3ebc2a00} /* (17, 16, 29) {real, imag} */,
  {32'h3f3cfef8, 32'hbf3bc0a8} /* (17, 16, 28) {real, imag} */,
  {32'hbd851538, 32'hbf6bcc44} /* (17, 16, 27) {real, imag} */,
  {32'hbf6156b2, 32'hbf54f0d0} /* (17, 16, 26) {real, imag} */,
  {32'h3ed0b3c4, 32'hbe9d8c18} /* (17, 16, 25) {real, imag} */,
  {32'h3f6adb39, 32'h3f3d1ab4} /* (17, 16, 24) {real, imag} */,
  {32'hbe83bbb2, 32'h3fb85786} /* (17, 16, 23) {real, imag} */,
  {32'h3ef79829, 32'h3f2b6352} /* (17, 16, 22) {real, imag} */,
  {32'hbea0d540, 32'h3e36fe50} /* (17, 16, 21) {real, imag} */,
  {32'hbe12d4c0, 32'h3f85126a} /* (17, 16, 20) {real, imag} */,
  {32'h3ecdfcbc, 32'h3e437978} /* (17, 16, 19) {real, imag} */,
  {32'h3d94b440, 32'hbec69640} /* (17, 16, 18) {real, imag} */,
  {32'h3d7ec5f0, 32'hbefaf8d0} /* (17, 16, 17) {real, imag} */,
  {32'h3f621fcc, 32'hbfc1d63c} /* (17, 16, 16) {real, imag} */,
  {32'h3bc10a00, 32'h3c922000} /* (17, 16, 15) {real, imag} */,
  {32'hbf83fc50, 32'h3df890c0} /* (17, 16, 14) {real, imag} */,
  {32'h3f67a8ba, 32'hbf5ce538} /* (17, 16, 13) {real, imag} */,
  {32'h3fef7d37, 32'hbe5200a8} /* (17, 16, 12) {real, imag} */,
  {32'h3d1bbd20, 32'h3f806bbf} /* (17, 16, 11) {real, imag} */,
  {32'hbdd2a188, 32'h3eacacac} /* (17, 16, 10) {real, imag} */,
  {32'hbe8a5c98, 32'hbf1839b8} /* (17, 16, 9) {real, imag} */,
  {32'hbff4c7b0, 32'h3f0de10c} /* (17, 16, 8) {real, imag} */,
  {32'hbe8dd194, 32'hbf6367b0} /* (17, 16, 7) {real, imag} */,
  {32'h4007ceaa, 32'hbfdcd5aa} /* (17, 16, 6) {real, imag} */,
  {32'hbeb881b8, 32'hbf9667c7} /* (17, 16, 5) {real, imag} */,
  {32'hbf56fcec, 32'hbe8e9960} /* (17, 16, 4) {real, imag} */,
  {32'h3e027b88, 32'h3b7c6000} /* (17, 16, 3) {real, imag} */,
  {32'hbf62e3c2, 32'hc018e392} /* (17, 16, 2) {real, imag} */,
  {32'hbf8f97ba, 32'hbf84dc96} /* (17, 16, 1) {real, imag} */,
  {32'hbe0232bc, 32'h3f4afbb0} /* (17, 16, 0) {real, imag} */,
  {32'hbe71da70, 32'hbf30d078} /* (17, 15, 31) {real, imag} */,
  {32'h3f6e9a7d, 32'hbfb6dc2b} /* (17, 15, 30) {real, imag} */,
  {32'hbe28847c, 32'hbf45fc1a} /* (17, 15, 29) {real, imag} */,
  {32'hbf8464cc, 32'hbf13f9da} /* (17, 15, 28) {real, imag} */,
  {32'h3dc99480, 32'hbf177b63} /* (17, 15, 27) {real, imag} */,
  {32'hbd675b80, 32'hbf02e0c2} /* (17, 15, 26) {real, imag} */,
  {32'hbf6406ec, 32'hbda86c98} /* (17, 15, 25) {real, imag} */,
  {32'h3f778d2f, 32'h3f7b67ac} /* (17, 15, 24) {real, imag} */,
  {32'h3e929b92, 32'h3d64e580} /* (17, 15, 23) {real, imag} */,
  {32'h3de45bc0, 32'hbfc0d4bf} /* (17, 15, 22) {real, imag} */,
  {32'h3ec22ead, 32'h3f4f655a} /* (17, 15, 21) {real, imag} */,
  {32'h3e71922c, 32'h3fef656e} /* (17, 15, 20) {real, imag} */,
  {32'h3e0e1a60, 32'h3ee15d52} /* (17, 15, 19) {real, imag} */,
  {32'hbf4a8b27, 32'h3f8214fa} /* (17, 15, 18) {real, imag} */,
  {32'hbe2ab1d0, 32'h3f295a4e} /* (17, 15, 17) {real, imag} */,
  {32'h3f1a6135, 32'h3e8509d6} /* (17, 15, 16) {real, imag} */,
  {32'h3d059a00, 32'h3ef08b78} /* (17, 15, 15) {real, imag} */,
  {32'hbf233a8a, 32'hbd7422a0} /* (17, 15, 14) {real, imag} */,
  {32'hbe4e6d28, 32'hbe557d58} /* (17, 15, 13) {real, imag} */,
  {32'h3edc4e20, 32'hbf4c645c} /* (17, 15, 12) {real, imag} */,
  {32'h3f7314c4, 32'hbeeafc8c} /* (17, 15, 11) {real, imag} */,
  {32'h3d5ee700, 32'hbf1d14f0} /* (17, 15, 10) {real, imag} */,
  {32'hbfbfe41c, 32'hbf86e162} /* (17, 15, 9) {real, imag} */,
  {32'hbf1ac21a, 32'hbf12882c} /* (17, 15, 8) {real, imag} */,
  {32'hbd7e89c0, 32'h3dfa5ce0} /* (17, 15, 7) {real, imag} */,
  {32'h3e52c2dc, 32'hbef7ee2c} /* (17, 15, 6) {real, imag} */,
  {32'h3eebf058, 32'hbf266353} /* (17, 15, 5) {real, imag} */,
  {32'hbe59b528, 32'hbeb6497e} /* (17, 15, 4) {real, imag} */,
  {32'hbf5ed579, 32'hc00e5536} /* (17, 15, 3) {real, imag} */,
  {32'h3f73dc64, 32'hbeb938a4} /* (17, 15, 2) {real, imag} */,
  {32'h3e94df76, 32'hbf2cd354} /* (17, 15, 1) {real, imag} */,
  {32'hbe9e4514, 32'hbf8038c2} /* (17, 15, 0) {real, imag} */,
  {32'h3ee4c44a, 32'hbe3a44dc} /* (17, 14, 31) {real, imag} */,
  {32'hbfb39a7d, 32'hbfb89e67} /* (17, 14, 30) {real, imag} */,
  {32'hbf8ffe3f, 32'h3f78ddbc} /* (17, 14, 29) {real, imag} */,
  {32'h3e899e33, 32'h3f87721a} /* (17, 14, 28) {real, imag} */,
  {32'h3fe3e40a, 32'hbd02c5c0} /* (17, 14, 27) {real, imag} */,
  {32'h3ec733a0, 32'h3e6b10a8} /* (17, 14, 26) {real, imag} */,
  {32'hbf674448, 32'h3f0df8bd} /* (17, 14, 25) {real, imag} */,
  {32'h3e028614, 32'h3f61bd90} /* (17, 14, 24) {real, imag} */,
  {32'h3f14a477, 32'h3fb7a6aa} /* (17, 14, 23) {real, imag} */,
  {32'hbf9ca65c, 32'h3f318110} /* (17, 14, 22) {real, imag} */,
  {32'hbff8f48c, 32'h3f2363f2} /* (17, 14, 21) {real, imag} */,
  {32'hbf6941bd, 32'hbe1aea2c} /* (17, 14, 20) {real, imag} */,
  {32'h3f1a003a, 32'h3f2d4328} /* (17, 14, 19) {real, imag} */,
  {32'h3fe0ac82, 32'h3f41742a} /* (17, 14, 18) {real, imag} */,
  {32'h3eacda80, 32'h3f77f00c} /* (17, 14, 17) {real, imag} */,
  {32'h3ebcfa90, 32'h3f74861c} /* (17, 14, 16) {real, imag} */,
  {32'hbe6163cc, 32'hbe408860} /* (17, 14, 15) {real, imag} */,
  {32'hbee042a2, 32'hbf0fbc3d} /* (17, 14, 14) {real, imag} */,
  {32'hbf0164e3, 32'hbf49846f} /* (17, 14, 13) {real, imag} */,
  {32'hbf4ff0a5, 32'h3fbd1166} /* (17, 14, 12) {real, imag} */,
  {32'hbf3cb0dc, 32'h3e304d1e} /* (17, 14, 11) {real, imag} */,
  {32'hbfb30190, 32'h3f90d5cf} /* (17, 14, 10) {real, imag} */,
  {32'hbe9c66d6, 32'h3ebb88ec} /* (17, 14, 9) {real, imag} */,
  {32'hbfef94e7, 32'hbfaf3972} /* (17, 14, 8) {real, imag} */,
  {32'hbfdccecd, 32'hbfc04b06} /* (17, 14, 7) {real, imag} */,
  {32'h3f565cf7, 32'hbef9aa62} /* (17, 14, 6) {real, imag} */,
  {32'h3f7be5ba, 32'hbf0efcb1} /* (17, 14, 5) {real, imag} */,
  {32'h3f32e0e4, 32'h3f94cb59} /* (17, 14, 4) {real, imag} */,
  {32'hbe26fbb4, 32'h3d8b4b40} /* (17, 14, 3) {real, imag} */,
  {32'hbe8ef14c, 32'hbf7225eb} /* (17, 14, 2) {real, imag} */,
  {32'h4078d6ce, 32'h3f0ca1e4} /* (17, 14, 1) {real, imag} */,
  {32'h403e60a0, 32'h3f75cf3f} /* (17, 14, 0) {real, imag} */,
  {32'h3ef1ba54, 32'h3eba0828} /* (17, 13, 31) {real, imag} */,
  {32'hbead8a34, 32'h3f08b5cc} /* (17, 13, 30) {real, imag} */,
  {32'h3f009f7c, 32'hbf462760} /* (17, 13, 29) {real, imag} */,
  {32'h40817326, 32'h3f0127b2} /* (17, 13, 28) {real, imag} */,
  {32'h4026b21a, 32'hbef33a88} /* (17, 13, 27) {real, imag} */,
  {32'h3f063681, 32'hbfca474d} /* (17, 13, 26) {real, imag} */,
  {32'hbfb496e7, 32'hbf1302c7} /* (17, 13, 25) {real, imag} */,
  {32'hbe7c1e8c, 32'hbe55287c} /* (17, 13, 24) {real, imag} */,
  {32'hbf042156, 32'hbf85ec8c} /* (17, 13, 23) {real, imag} */,
  {32'hbf33c84b, 32'hbf2332a6} /* (17, 13, 22) {real, imag} */,
  {32'hbf664777, 32'hbf8ea571} /* (17, 13, 21) {real, imag} */,
  {32'hbf0fb47c, 32'h3fc08ac4} /* (17, 13, 20) {real, imag} */,
  {32'hbf2cdb59, 32'h3e16accb} /* (17, 13, 19) {real, imag} */,
  {32'hbf920d33, 32'h3f88ae48} /* (17, 13, 18) {real, imag} */,
  {32'hbf870779, 32'hbcd82980} /* (17, 13, 17) {real, imag} */,
  {32'hbea6fda4, 32'hc0313045} /* (17, 13, 16) {real, imag} */,
  {32'hbd0a31e0, 32'hbf76836e} /* (17, 13, 15) {real, imag} */,
  {32'hbf4bff87, 32'hbacf5a00} /* (17, 13, 14) {real, imag} */,
  {32'hbe8a3c2c, 32'h3f6aedbf} /* (17, 13, 13) {real, imag} */,
  {32'h3e8dedc0, 32'h3eb9aff0} /* (17, 13, 12) {real, imag} */,
  {32'hbf309a9e, 32'hbebd7f3a} /* (17, 13, 11) {real, imag} */,
  {32'hbf8fc0a0, 32'hbf32f5a6} /* (17, 13, 10) {real, imag} */,
  {32'hbcbe0cc0, 32'hbf797f04} /* (17, 13, 9) {real, imag} */,
  {32'h3f9c328b, 32'hbf5b215d} /* (17, 13, 8) {real, imag} */,
  {32'h3f16028d, 32'hbef1ef20} /* (17, 13, 7) {real, imag} */,
  {32'h3f16df58, 32'hbee07be0} /* (17, 13, 6) {real, imag} */,
  {32'hbf1b014d, 32'h3fb29b5e} /* (17, 13, 5) {real, imag} */,
  {32'hbf8c6635, 32'h3f6272b8} /* (17, 13, 4) {real, imag} */,
  {32'h3d2e52e0, 32'h3fed671c} /* (17, 13, 3) {real, imag} */,
  {32'hbfc3bd7c, 32'h4001f4b0} /* (17, 13, 2) {real, imag} */,
  {32'h3f2d9c09, 32'hbd23ef60} /* (17, 13, 1) {real, imag} */,
  {32'h3f236374, 32'hbf8ac56e} /* (17, 13, 0) {real, imag} */,
  {32'hbf66616b, 32'hbf838547} /* (17, 12, 31) {real, imag} */,
  {32'hbc3c8d80, 32'hbc5548c0} /* (17, 12, 30) {real, imag} */,
  {32'h3ed400ec, 32'hc003b51a} /* (17, 12, 29) {real, imag} */,
  {32'hbf87a557, 32'hc004db14} /* (17, 12, 28) {real, imag} */,
  {32'hbfd3740c, 32'hbf9be794} /* (17, 12, 27) {real, imag} */,
  {32'hbf8ec366, 32'hbf1dbce6} /* (17, 12, 26) {real, imag} */,
  {32'h3ea85378, 32'hbe34b818} /* (17, 12, 25) {real, imag} */,
  {32'hc00a1a1d, 32'hbc129600} /* (17, 12, 24) {real, imag} */,
  {32'hbf80910c, 32'h3b5fba00} /* (17, 12, 23) {real, imag} */,
  {32'h3e704768, 32'h3f88ebc7} /* (17, 12, 22) {real, imag} */,
  {32'h3e51d76c, 32'hbf475e33} /* (17, 12, 21) {real, imag} */,
  {32'h3f374d2a, 32'hbeed4a56} /* (17, 12, 20) {real, imag} */,
  {32'hbf6263ea, 32'hbe175dd0} /* (17, 12, 19) {real, imag} */,
  {32'hbec5fc1a, 32'hbf167042} /* (17, 12, 18) {real, imag} */,
  {32'h400de298, 32'h400fe3c2} /* (17, 12, 17) {real, imag} */,
  {32'h3ffb031e, 32'h3f5c349a} /* (17, 12, 16) {real, imag} */,
  {32'h3f42b17e, 32'hbe2b83e8} /* (17, 12, 15) {real, imag} */,
  {32'h3f6451ce, 32'h3ea2fb82} /* (17, 12, 14) {real, imag} */,
  {32'hbdcc0400, 32'hbfebf9b6} /* (17, 12, 13) {real, imag} */,
  {32'h400ecfb4, 32'hc02cbb0b} /* (17, 12, 12) {real, imag} */,
  {32'h3f8f1c07, 32'hc0074306} /* (17, 12, 11) {real, imag} */,
  {32'h3e65dd58, 32'hbeb95db0} /* (17, 12, 10) {real, imag} */,
  {32'h401d59c2, 32'h3ff9e8d7} /* (17, 12, 9) {real, imag} */,
  {32'h3f21c1a7, 32'hbd575b80} /* (17, 12, 8) {real, imag} */,
  {32'h3e53f57c, 32'hc049b3e4} /* (17, 12, 7) {real, imag} */,
  {32'h3f455ea5, 32'hbf5efd24} /* (17, 12, 6) {real, imag} */,
  {32'hbf0d3949, 32'h3f491c46} /* (17, 12, 5) {real, imag} */,
  {32'h3fdbf32a, 32'h3ebb99f8} /* (17, 12, 4) {real, imag} */,
  {32'hbbdb15c0, 32'hbd4a4860} /* (17, 12, 3) {real, imag} */,
  {32'hbefe1ae6, 32'h402f7cf2} /* (17, 12, 2) {real, imag} */,
  {32'hbfda46cc, 32'h4028f29e} /* (17, 12, 1) {real, imag} */,
  {32'h3e71af68, 32'hbea9ca8b} /* (17, 12, 0) {real, imag} */,
  {32'hbf912e4a, 32'h3d7a5c80} /* (17, 11, 31) {real, imag} */,
  {32'hbfae47be, 32'h3fa64088} /* (17, 11, 30) {real, imag} */,
  {32'hbf79aaac, 32'h3e23a990} /* (17, 11, 29) {real, imag} */,
  {32'hc045fa4e, 32'h3fdc3edf} /* (17, 11, 28) {real, imag} */,
  {32'hc022c224, 32'h3f6acbbe} /* (17, 11, 27) {real, imag} */,
  {32'hc00ef130, 32'h4015b612} /* (17, 11, 26) {real, imag} */,
  {32'h3eb7f328, 32'hbefc4698} /* (17, 11, 25) {real, imag} */,
  {32'h3fe5c4da, 32'hc01c0105} /* (17, 11, 24) {real, imag} */,
  {32'h3d928904, 32'hc03b45c0} /* (17, 11, 23) {real, imag} */,
  {32'hbfb2f644, 32'hbffd8b25} /* (17, 11, 22) {real, imag} */,
  {32'h3f81f313, 32'h3fc57f58} /* (17, 11, 21) {real, imag} */,
  {32'h3f934b0d, 32'h40249bcd} /* (17, 11, 20) {real, imag} */,
  {32'h402944f5, 32'h3fc37482} /* (17, 11, 19) {real, imag} */,
  {32'h404cb73b, 32'h3eb4fe52} /* (17, 11, 18) {real, imag} */,
  {32'h4009102c, 32'hc016c70e} /* (17, 11, 17) {real, imag} */,
  {32'h400b94a0, 32'hbfaa768d} /* (17, 11, 16) {real, imag} */,
  {32'hbf93585b, 32'hbfa0756b} /* (17, 11, 15) {real, imag} */,
  {32'hbfd618c2, 32'hbfbd7462} /* (17, 11, 14) {real, imag} */,
  {32'h3fa377d4, 32'h3f935078} /* (17, 11, 13) {real, imag} */,
  {32'hbfc4fb32, 32'h3fc49493} /* (17, 11, 12) {real, imag} */,
  {32'hc00ee098, 32'h3e2a0e60} /* (17, 11, 11) {real, imag} */,
  {32'hbed86afc, 32'hc0597172} /* (17, 11, 10) {real, imag} */,
  {32'hbf007e30, 32'hc04f1834} /* (17, 11, 9) {real, imag} */,
  {32'hbecafd6e, 32'hbf23e312} /* (17, 11, 8) {real, imag} */,
  {32'h402901b4, 32'hbf70517e} /* (17, 11, 7) {real, imag} */,
  {32'h3ff8dade, 32'hbf9ed49e} /* (17, 11, 6) {real, imag} */,
  {32'hbda4fba0, 32'hbf97b8ba} /* (17, 11, 5) {real, imag} */,
  {32'hbd452090, 32'hc06105a5} /* (17, 11, 4) {real, imag} */,
  {32'h3f878cc5, 32'hbf542469} /* (17, 11, 3) {real, imag} */,
  {32'h404fbcc3, 32'h3faab107} /* (17, 11, 2) {real, imag} */,
  {32'h3fb3be86, 32'h3f02cd00} /* (17, 11, 1) {real, imag} */,
  {32'hbf40e561, 32'h3f304216} /* (17, 11, 0) {real, imag} */,
  {32'hbe56809c, 32'h40371295} /* (17, 10, 31) {real, imag} */,
  {32'h3f3156b0, 32'h408e1444} /* (17, 10, 30) {real, imag} */,
  {32'hc0257dc0, 32'h3fd568b8} /* (17, 10, 29) {real, imag} */,
  {32'hc01c706c, 32'h3fd2d315} /* (17, 10, 28) {real, imag} */,
  {32'hbe9b8a74, 32'h401a33b9} /* (17, 10, 27) {real, imag} */,
  {32'h3db630e0, 32'h40357f8a} /* (17, 10, 26) {real, imag} */,
  {32'hbfefb842, 32'h4096c8c3} /* (17, 10, 25) {real, imag} */,
  {32'hbfe46ac7, 32'h40690e99} /* (17, 10, 24) {real, imag} */,
  {32'h4033ef27, 32'h40be217a} /* (17, 10, 23) {real, imag} */,
  {32'h408834a3, 32'h3fbe2f33} /* (17, 10, 22) {real, imag} */,
  {32'h3f4bf526, 32'hbf656ce8} /* (17, 10, 21) {real, imag} */,
  {32'h3fb9ba0f, 32'h3eb3f884} /* (17, 10, 20) {real, imag} */,
  {32'hbef80e0c, 32'hbf232e02} /* (17, 10, 19) {real, imag} */,
  {32'hbf0cfe6b, 32'h3ea95598} /* (17, 10, 18) {real, imag} */,
  {32'h3fabba7a, 32'h3f993496} /* (17, 10, 17) {real, imag} */,
  {32'h4006b866, 32'hbfd7e88f} /* (17, 10, 16) {real, imag} */,
  {32'h3fee24c1, 32'hc038e89f} /* (17, 10, 15) {real, imag} */,
  {32'h4085b272, 32'hc0151413} /* (17, 10, 14) {real, imag} */,
  {32'h4052b18e, 32'h390fa000} /* (17, 10, 13) {real, imag} */,
  {32'h3f5b2aa0, 32'hbe79e760} /* (17, 10, 12) {real, imag} */,
  {32'hbf18d89b, 32'hbfbcf747} /* (17, 10, 11) {real, imag} */,
  {32'hbf1d8366, 32'hbff398c6} /* (17, 10, 10) {real, imag} */,
  {32'h3ffaaee2, 32'hbec0746d} /* (17, 10, 9) {real, imag} */,
  {32'h3f83d99a, 32'h3ff60fe2} /* (17, 10, 8) {real, imag} */,
  {32'h406c3300, 32'hc0314f8c} /* (17, 10, 7) {real, imag} */,
  {32'h3fa207db, 32'hbf02d1ca} /* (17, 10, 6) {real, imag} */,
  {32'hc05d8e72, 32'h3e9eae1a} /* (17, 10, 5) {real, imag} */,
  {32'hc03c9644, 32'hbf3d81f8} /* (17, 10, 4) {real, imag} */,
  {32'hc076e614, 32'hc03320e9} /* (17, 10, 3) {real, imag} */,
  {32'hc02ae67d, 32'hbf7319fc} /* (17, 10, 2) {real, imag} */,
  {32'hc007baba, 32'hbebe1cc2} /* (17, 10, 1) {real, imag} */,
  {32'hbecf0cb3, 32'h3d981230} /* (17, 10, 0) {real, imag} */,
  {32'hc014188d, 32'h3f5359ce} /* (17, 9, 31) {real, imag} */,
  {32'hc0187b96, 32'hbf714be7} /* (17, 9, 30) {real, imag} */,
  {32'h3f88c6f7, 32'hbfd2c606} /* (17, 9, 29) {real, imag} */,
  {32'h3fae3b13, 32'h4027de5c} /* (17, 9, 28) {real, imag} */,
  {32'h3f01fc14, 32'h3fa704ec} /* (17, 9, 27) {real, imag} */,
  {32'hbf2c8720, 32'hbf15d35e} /* (17, 9, 26) {real, imag} */,
  {32'h3ed0a418, 32'h3f4cedea} /* (17, 9, 25) {real, imag} */,
  {32'h3f7d2e3f, 32'h404bec70} /* (17, 9, 24) {real, imag} */,
  {32'hbf8c07ac, 32'h40758438} /* (17, 9, 23) {real, imag} */,
  {32'hc0574ac6, 32'h408c5b63} /* (17, 9, 22) {real, imag} */,
  {32'h400889b5, 32'h404174e5} /* (17, 9, 21) {real, imag} */,
  {32'h3fb9e475, 32'h4055d239} /* (17, 9, 20) {real, imag} */,
  {32'hc072f5c3, 32'hbe7b2630} /* (17, 9, 19) {real, imag} */,
  {32'h3f2a30d8, 32'hbf9ad40d} /* (17, 9, 18) {real, imag} */,
  {32'h3f9bc783, 32'h403377e0} /* (17, 9, 17) {real, imag} */,
  {32'hbe9d1fae, 32'h404c9f1d} /* (17, 9, 16) {real, imag} */,
  {32'h3ff63816, 32'h3f09cdec} /* (17, 9, 15) {real, imag} */,
  {32'h40a935c0, 32'hbfc009b0} /* (17, 9, 14) {real, imag} */,
  {32'h40d72adc, 32'h3e198b18} /* (17, 9, 13) {real, imag} */,
  {32'h3f17cb60, 32'h3fae3bda} /* (17, 9, 12) {real, imag} */,
  {32'hbf594756, 32'h3d866d80} /* (17, 9, 11) {real, imag} */,
  {32'hc0319166, 32'hbeeee7c2} /* (17, 9, 10) {real, imag} */,
  {32'hc09d0cff, 32'h3ef6346c} /* (17, 9, 9) {real, imag} */,
  {32'hc07cace5, 32'h40596441} /* (17, 9, 8) {real, imag} */,
  {32'hc05ddc0a, 32'h3fd611fc} /* (17, 9, 7) {real, imag} */,
  {32'h3e793b10, 32'h3ac53800} /* (17, 9, 6) {real, imag} */,
  {32'h402eb922, 32'h3fb0ffdc} /* (17, 9, 5) {real, imag} */,
  {32'h404017e2, 32'h3f8e5188} /* (17, 9, 4) {real, imag} */,
  {32'h3ed7e27c, 32'h4017d6a4} /* (17, 9, 3) {real, imag} */,
  {32'hbf6267a0, 32'h3ea99c60} /* (17, 9, 2) {real, imag} */,
  {32'h3ed4f790, 32'hbf5743e2} /* (17, 9, 1) {real, imag} */,
  {32'hbfb93156, 32'h3f7f54c0} /* (17, 9, 0) {real, imag} */,
  {32'hc0018f4a, 32'h40439232} /* (17, 8, 31) {real, imag} */,
  {32'hbfc83e64, 32'hbd26c6c0} /* (17, 8, 30) {real, imag} */,
  {32'hbeb2b158, 32'hbf8a34eb} /* (17, 8, 29) {real, imag} */,
  {32'hbec43580, 32'hbe4f7628} /* (17, 8, 28) {real, imag} */,
  {32'hbf87546a, 32'hbf31791c} /* (17, 8, 27) {real, imag} */,
  {32'hbf7a59cb, 32'hbfc8f6da} /* (17, 8, 26) {real, imag} */,
  {32'h3efe3164, 32'h404f0a01} /* (17, 8, 25) {real, imag} */,
  {32'h3fb84696, 32'h402b45bf} /* (17, 8, 24) {real, imag} */,
  {32'h4012fe10, 32'h400916be} /* (17, 8, 23) {real, imag} */,
  {32'h3fddefa8, 32'h3eba0de0} /* (17, 8, 22) {real, imag} */,
  {32'h402ad772, 32'hbf68a598} /* (17, 8, 21) {real, imag} */,
  {32'h40862c4e, 32'hc0058821} /* (17, 8, 20) {real, imag} */,
  {32'h4085d2b1, 32'hbfe8b093} /* (17, 8, 19) {real, imag} */,
  {32'h3ff6f69b, 32'hbf1f0920} /* (17, 8, 18) {real, imag} */,
  {32'h3f42cfe4, 32'h40340d74} /* (17, 8, 17) {real, imag} */,
  {32'h3fa43f62, 32'h407a42c5} /* (17, 8, 16) {real, imag} */,
  {32'hbc973bc0, 32'h3f9817de} /* (17, 8, 15) {real, imag} */,
  {32'hc04763f0, 32'hbf86245c} /* (17, 8, 14) {real, imag} */,
  {32'hc07fa31f, 32'hc0ca8a22} /* (17, 8, 13) {real, imag} */,
  {32'hc0149928, 32'hc03c391e} /* (17, 8, 12) {real, imag} */,
  {32'hbe1b8de4, 32'h402e8f14} /* (17, 8, 11) {real, imag} */,
  {32'h3fb794fc, 32'h404bef81} /* (17, 8, 10) {real, imag} */,
  {32'hbef208a8, 32'h3e3af2b0} /* (17, 8, 9) {real, imag} */,
  {32'h3f72d71e, 32'hbf92b474} /* (17, 8, 8) {real, imag} */,
  {32'hc07b6d76, 32'h3f94b4b8} /* (17, 8, 7) {real, imag} */,
  {32'hbfef4b34, 32'hc0769d60} /* (17, 8, 6) {real, imag} */,
  {32'hbafeb800, 32'hbeb09c4c} /* (17, 8, 5) {real, imag} */,
  {32'hbf777724, 32'h3eda5fd8} /* (17, 8, 4) {real, imag} */,
  {32'h3e1ac068, 32'h40222c3f} /* (17, 8, 3) {real, imag} */,
  {32'hbe559288, 32'h4046f80d} /* (17, 8, 2) {real, imag} */,
  {32'hbf08b7e5, 32'h4008c2ec} /* (17, 8, 1) {real, imag} */,
  {32'h3edab2a2, 32'h3f409dbc} /* (17, 8, 0) {real, imag} */,
  {32'h3e010774, 32'hbf24eced} /* (17, 7, 31) {real, imag} */,
  {32'hc051079e, 32'hc025377b} /* (17, 7, 30) {real, imag} */,
  {32'hc0ab25e6, 32'h3fb3c492} /* (17, 7, 29) {real, imag} */,
  {32'hc0ac6ec4, 32'h3fec18ca} /* (17, 7, 28) {real, imag} */,
  {32'hc0748056, 32'hc032a1ea} /* (17, 7, 27) {real, imag} */,
  {32'hc0b9aa68, 32'hc0821e3f} /* (17, 7, 26) {real, imag} */,
  {32'hc06c41d0, 32'h3f5754f8} /* (17, 7, 25) {real, imag} */,
  {32'h3fcbd09c, 32'hbfbedb41} /* (17, 7, 24) {real, imag} */,
  {32'h3f20ef40, 32'hbfe0f17e} /* (17, 7, 23) {real, imag} */,
  {32'hbf10284c, 32'h3fdc33c1} /* (17, 7, 22) {real, imag} */,
  {32'hc04971d8, 32'hbe112c58} /* (17, 7, 21) {real, imag} */,
  {32'h3f687bc4, 32'hc085f747} /* (17, 7, 20) {real, imag} */,
  {32'h3d0583e0, 32'h3ec5fef4} /* (17, 7, 19) {real, imag} */,
  {32'hbd63b3c0, 32'hc0529fd9} /* (17, 7, 18) {real, imag} */,
  {32'h3fdd41df, 32'hc0b5cbe7} /* (17, 7, 17) {real, imag} */,
  {32'hc0249d77, 32'hc0891d6f} /* (17, 7, 16) {real, imag} */,
  {32'hc0492019, 32'hbebbd55b} /* (17, 7, 15) {real, imag} */,
  {32'hc017bd5f, 32'h3fe65f28} /* (17, 7, 14) {real, imag} */,
  {32'h3f2f610c, 32'h4002bd47} /* (17, 7, 13) {real, imag} */,
  {32'hbecf0c80, 32'hc024bff3} /* (17, 7, 12) {real, imag} */,
  {32'hc0175094, 32'h3f591ede} /* (17, 7, 11) {real, imag} */,
  {32'hbfb00e47, 32'h4010def5} /* (17, 7, 10) {real, imag} */,
  {32'hbf22b06a, 32'hc0099c40} /* (17, 7, 9) {real, imag} */,
  {32'hbe0996f0, 32'h3dc3c670} /* (17, 7, 8) {real, imag} */,
  {32'hc00740be, 32'hbdd82378} /* (17, 7, 7) {real, imag} */,
  {32'hc085535e, 32'h400e9bf0} /* (17, 7, 6) {real, imag} */,
  {32'hbf7ebee8, 32'h408d955a} /* (17, 7, 5) {real, imag} */,
  {32'hc004dcef, 32'hbf343b70} /* (17, 7, 4) {real, imag} */,
  {32'h3fca8819, 32'h3e845c1c} /* (17, 7, 3) {real, imag} */,
  {32'h3ff33f12, 32'h3eccbd10} /* (17, 7, 2) {real, imag} */,
  {32'h3f47183f, 32'h4032d980} /* (17, 7, 1) {real, imag} */,
  {32'hc0425ee5, 32'hbe537490} /* (17, 7, 0) {real, imag} */,
  {32'hbfbff6ac, 32'h3fe6cc60} /* (17, 6, 31) {real, imag} */,
  {32'hc0225a1c, 32'h3fd8738d} /* (17, 6, 30) {real, imag} */,
  {32'hc06f8e0a, 32'h4022ea19} /* (17, 6, 29) {real, imag} */,
  {32'h3ef12d20, 32'h3f062936} /* (17, 6, 28) {real, imag} */,
  {32'hc019591e, 32'h3e2e1184} /* (17, 6, 27) {real, imag} */,
  {32'hbf8816a8, 32'hc0322dac} /* (17, 6, 26) {real, imag} */,
  {32'hbf65ca23, 32'hc0859eb9} /* (17, 6, 25) {real, imag} */,
  {32'hc018863c, 32'hbfabb8e5} /* (17, 6, 24) {real, imag} */,
  {32'hc0404d5f, 32'h3ff38e5a} /* (17, 6, 23) {real, imag} */,
  {32'hbf94678b, 32'hbf1d9626} /* (17, 6, 22) {real, imag} */,
  {32'h3fce9199, 32'hc019322a} /* (17, 6, 21) {real, imag} */,
  {32'h3ffb27c7, 32'hbfc0aeb6} /* (17, 6, 20) {real, imag} */,
  {32'hc011f192, 32'hbf4d3bb6} /* (17, 6, 19) {real, imag} */,
  {32'hc0226e0d, 32'hbf2aeb1c} /* (17, 6, 18) {real, imag} */,
  {32'h4019b273, 32'h3fda0954} /* (17, 6, 17) {real, imag} */,
  {32'hc0890d88, 32'h400772cf} /* (17, 6, 16) {real, imag} */,
  {32'hc05f1ade, 32'h404e4c6a} /* (17, 6, 15) {real, imag} */,
  {32'h4033f0c0, 32'h3f4b7c83} /* (17, 6, 14) {real, imag} */,
  {32'h3fdc2b81, 32'h40bf1649} /* (17, 6, 13) {real, imag} */,
  {32'h408e0aeb, 32'h40d11a10} /* (17, 6, 12) {real, imag} */,
  {32'h40723323, 32'h4076e7a8} /* (17, 6, 11) {real, imag} */,
  {32'h3f8aaf12, 32'hbec019c4} /* (17, 6, 10) {real, imag} */,
  {32'h3f9f5b05, 32'h3f298414} /* (17, 6, 9) {real, imag} */,
  {32'h3fd8ae86, 32'h409f7bd4} /* (17, 6, 8) {real, imag} */,
  {32'hc00d9b47, 32'h402871ee} /* (17, 6, 7) {real, imag} */,
  {32'hc0854dbb, 32'h407480f3} /* (17, 6, 6) {real, imag} */,
  {32'hc0eab509, 32'h401ce888} /* (17, 6, 5) {real, imag} */,
  {32'hc02f332a, 32'h40486bfd} /* (17, 6, 4) {real, imag} */,
  {32'hc05aa607, 32'h3f2554bc} /* (17, 6, 3) {real, imag} */,
  {32'hc0bb0e0e, 32'hc0a21eea} /* (17, 6, 2) {real, imag} */,
  {32'hc02c0ef8, 32'hbde0f9c0} /* (17, 6, 1) {real, imag} */,
  {32'hc0899c30, 32'h408396ac} /* (17, 6, 0) {real, imag} */,
  {32'h3fd4262c, 32'hbf89f506} /* (17, 5, 31) {real, imag} */,
  {32'h3f48eb00, 32'hbf29a516} /* (17, 5, 30) {real, imag} */,
  {32'h3db7a55c, 32'hbf05cd61} /* (17, 5, 29) {real, imag} */,
  {32'h40999e24, 32'hc012f028} /* (17, 5, 28) {real, imag} */,
  {32'hc0709e04, 32'hbf5cd628} /* (17, 5, 27) {real, imag} */,
  {32'hc0957004, 32'h3f923b2e} /* (17, 5, 26) {real, imag} */,
  {32'hc001fccf, 32'hc0383031} /* (17, 5, 25) {real, imag} */,
  {32'hc0ac982c, 32'hc061d250} /* (17, 5, 24) {real, imag} */,
  {32'hc000e26b, 32'hbebe937c} /* (17, 5, 23) {real, imag} */,
  {32'h402b5320, 32'h401c2572} /* (17, 5, 22) {real, imag} */,
  {32'hc0379d7b, 32'h4005c134} /* (17, 5, 21) {real, imag} */,
  {32'hc0bc04fd, 32'h40389023} /* (17, 5, 20) {real, imag} */,
  {32'hc044831f, 32'h3fccc68e} /* (17, 5, 19) {real, imag} */,
  {32'hbfd17cbc, 32'hbe0a9bf8} /* (17, 5, 18) {real, imag} */,
  {32'h3fb651dd, 32'h3f1247af} /* (17, 5, 17) {real, imag} */,
  {32'h40892990, 32'h3f9fbc82} /* (17, 5, 16) {real, imag} */,
  {32'h402ffee0, 32'h40c1f2ed} /* (17, 5, 15) {real, imag} */,
  {32'h40dc6061, 32'h409f7608} /* (17, 5, 14) {real, imag} */,
  {32'h413769c0, 32'hc040d164} /* (17, 5, 13) {real, imag} */,
  {32'h412804d8, 32'hc05b64f4} /* (17, 5, 12) {real, imag} */,
  {32'h4045b9ea, 32'hc021980b} /* (17, 5, 11) {real, imag} */,
  {32'hc0246f6e, 32'hc064c0f1} /* (17, 5, 10) {real, imag} */,
  {32'hbfbf6fb2, 32'hbfdae8d0} /* (17, 5, 9) {real, imag} */,
  {32'h40091208, 32'hbfaf3cdf} /* (17, 5, 8) {real, imag} */,
  {32'h3f63a7b6, 32'hbfe2417c} /* (17, 5, 7) {real, imag} */,
  {32'hc035a47e, 32'hc03d4bf2} /* (17, 5, 6) {real, imag} */,
  {32'hc091c5f8, 32'hbff0d8c3} /* (17, 5, 5) {real, imag} */,
  {32'hbfb013cb, 32'hc01131a4} /* (17, 5, 4) {real, imag} */,
  {32'h4000e1a2, 32'h4047dcdd} /* (17, 5, 3) {real, imag} */,
  {32'h40b06955, 32'hbf8487d6} /* (17, 5, 2) {real, imag} */,
  {32'h3f051808, 32'hc09db2b8} /* (17, 5, 1) {real, imag} */,
  {32'h3fd34826, 32'hc0aab673} /* (17, 5, 0) {real, imag} */,
  {32'hbfa1ee28, 32'h40615624} /* (17, 4, 31) {real, imag} */,
  {32'hbff1b5e4, 32'h40702f6c} /* (17, 4, 30) {real, imag} */,
  {32'h3f399590, 32'h3e9ae370} /* (17, 4, 29) {real, imag} */,
  {32'h4060c14e, 32'hbfb2a7be} /* (17, 4, 28) {real, imag} */,
  {32'h408aa8c8, 32'hbf127252} /* (17, 4, 27) {real, imag} */,
  {32'h3ffb4b8c, 32'hbfc30edb} /* (17, 4, 26) {real, imag} */,
  {32'hbebc0248, 32'hbff75757} /* (17, 4, 25) {real, imag} */,
  {32'hc04ae5ec, 32'hbbc8e600} /* (17, 4, 24) {real, imag} */,
  {32'hbfafb6e0, 32'h408b3623} /* (17, 4, 23) {real, imag} */,
  {32'hc034a490, 32'h3fa9d745} /* (17, 4, 22) {real, imag} */,
  {32'h3e683312, 32'hbfb1fdee} /* (17, 4, 21) {real, imag} */,
  {32'hbf4427b4, 32'h402d26de} /* (17, 4, 20) {real, imag} */,
  {32'hbf965d99, 32'h40f4ecb5} /* (17, 4, 19) {real, imag} */,
  {32'h401029e9, 32'h413682de} /* (17, 4, 18) {real, imag} */,
  {32'h409b1a4d, 32'h40a8d0d6} /* (17, 4, 17) {real, imag} */,
  {32'h40302bbd, 32'hc0b37ff8} /* (17, 4, 16) {real, imag} */,
  {32'h3f9c3748, 32'hc0a59f8b} /* (17, 4, 15) {real, imag} */,
  {32'hbe24db08, 32'hbfbad021} /* (17, 4, 14) {real, imag} */,
  {32'hbfd13ae4, 32'hbffa363e} /* (17, 4, 13) {real, imag} */,
  {32'h3e5606b0, 32'hc0c2f473} /* (17, 4, 12) {real, imag} */,
  {32'h40a12864, 32'hc01aac32} /* (17, 4, 11) {real, imag} */,
  {32'h41110dc0, 32'h3f151db6} /* (17, 4, 10) {real, imag} */,
  {32'h4086c878, 32'h3ffe1646} /* (17, 4, 9) {real, imag} */,
  {32'h4042e884, 32'h3e36ee10} /* (17, 4, 8) {real, imag} */,
  {32'hc003a9ca, 32'h3f864ef4} /* (17, 4, 7) {real, imag} */,
  {32'hc0b63e48, 32'h40a931f3} /* (17, 4, 6) {real, imag} */,
  {32'hc06092d7, 32'h3f87d096} /* (17, 4, 5) {real, imag} */,
  {32'hbfe53a68, 32'h40731691} /* (17, 4, 4) {real, imag} */,
  {32'h3fc5d74a, 32'hbfaaacb5} /* (17, 4, 3) {real, imag} */,
  {32'h40296dab, 32'hc0efa6c0} /* (17, 4, 2) {real, imag} */,
  {32'h3e036590, 32'hc02c7b8a} /* (17, 4, 1) {real, imag} */,
  {32'h3f8cc75c, 32'h3e8d6e90} /* (17, 4, 0) {real, imag} */,
  {32'h40376a6b, 32'hc034bf02} /* (17, 3, 31) {real, imag} */,
  {32'h410271c2, 32'hbfafc43e} /* (17, 3, 30) {real, imag} */,
  {32'h403b6546, 32'h3f22011c} /* (17, 3, 29) {real, imag} */,
  {32'h4092b050, 32'hbc4b42c0} /* (17, 3, 28) {real, imag} */,
  {32'h40e49a31, 32'h4059348c} /* (17, 3, 27) {real, imag} */,
  {32'h4059a2ae, 32'h40a315c9} /* (17, 3, 26) {real, imag} */,
  {32'h3ee540a4, 32'h401dc08c} /* (17, 3, 25) {real, imag} */,
  {32'h4043c01d, 32'hc043a2e4} /* (17, 3, 24) {real, imag} */,
  {32'hc0780108, 32'h40042a1c} /* (17, 3, 23) {real, imag} */,
  {32'h3f997a9e, 32'h401874d6} /* (17, 3, 22) {real, imag} */,
  {32'h40ba694e, 32'h40593582} /* (17, 3, 21) {real, imag} */,
  {32'h410c45bc, 32'h4053d776} /* (17, 3, 20) {real, imag} */,
  {32'h3fb18686, 32'hbf5155d1} /* (17, 3, 19) {real, imag} */,
  {32'hbf9e8dda, 32'hc08e22e2} /* (17, 3, 18) {real, imag} */,
  {32'h4003bcc0, 32'hc08662b2} /* (17, 3, 17) {real, imag} */,
  {32'hbfd51f3d, 32'hbf6c911b} /* (17, 3, 16) {real, imag} */,
  {32'h3e83472c, 32'hc0116b24} /* (17, 3, 15) {real, imag} */,
  {32'hc045e41c, 32'hbf3e7a3e} /* (17, 3, 14) {real, imag} */,
  {32'hbf9f9936, 32'h3ee768f8} /* (17, 3, 13) {real, imag} */,
  {32'h40a4f892, 32'hbf389210} /* (17, 3, 12) {real, imag} */,
  {32'hc03b4fc8, 32'hc0247fd4} /* (17, 3, 11) {real, imag} */,
  {32'hc0a88b6a, 32'h3f73d9ac} /* (17, 3, 10) {real, imag} */,
  {32'h4079e408, 32'h408f3581} /* (17, 3, 9) {real, imag} */,
  {32'h40c9ea16, 32'h3eb618b6} /* (17, 3, 8) {real, imag} */,
  {32'hbea0f07c, 32'h3db7ffe0} /* (17, 3, 7) {real, imag} */,
  {32'h404b6d75, 32'h405fbc81} /* (17, 3, 6) {real, imag} */,
  {32'h400575e7, 32'h40869269} /* (17, 3, 5) {real, imag} */,
  {32'h3f835ea0, 32'h403660fa} /* (17, 3, 4) {real, imag} */,
  {32'h3f2acd10, 32'h3f3a17d4} /* (17, 3, 3) {real, imag} */,
  {32'hc03fd81f, 32'hbee0afd0} /* (17, 3, 2) {real, imag} */,
  {32'hbfde3f2e, 32'h3f2e9676} /* (17, 3, 1) {real, imag} */,
  {32'hbc96ad50, 32'h3ecad3ba} /* (17, 3, 0) {real, imag} */,
  {32'hbebc34c8, 32'hbf410150} /* (17, 2, 31) {real, imag} */,
  {32'h409c60c0, 32'hc04039c9} /* (17, 2, 30) {real, imag} */,
  {32'h40df24d7, 32'hc08e5df0} /* (17, 2, 29) {real, imag} */,
  {32'h3fa1c9ae, 32'hc0bd8ff2} /* (17, 2, 28) {real, imag} */,
  {32'hc06b83d3, 32'hc0913d80} /* (17, 2, 27) {real, imag} */,
  {32'hbff2a8a1, 32'hc0861de5} /* (17, 2, 26) {real, imag} */,
  {32'hc01ce42d, 32'hc0afaabc} /* (17, 2, 25) {real, imag} */,
  {32'hc00399d0, 32'hbfc26eb8} /* (17, 2, 24) {real, imag} */,
  {32'hbf35bb9a, 32'hc0324eae} /* (17, 2, 23) {real, imag} */,
  {32'hbf05b9fb, 32'h3f399438} /* (17, 2, 22) {real, imag} */,
  {32'hc002c83a, 32'h403874dc} /* (17, 2, 21) {real, imag} */,
  {32'hbfeb4805, 32'h40877e6f} /* (17, 2, 20) {real, imag} */,
  {32'h3edbb2c8, 32'h3fe10d04} /* (17, 2, 19) {real, imag} */,
  {32'hc0a84a2c, 32'h40acdd05} /* (17, 2, 18) {real, imag} */,
  {32'h3fe858f7, 32'h4099eab3} /* (17, 2, 17) {real, imag} */,
  {32'h410b0161, 32'h408205ba} /* (17, 2, 16) {real, imag} */,
  {32'h40480b68, 32'h3e28dd48} /* (17, 2, 15) {real, imag} */,
  {32'hbe6c09b0, 32'hc07e3c6e} /* (17, 2, 14) {real, imag} */,
  {32'hbfaef0c4, 32'hc034a5dc} /* (17, 2, 13) {real, imag} */,
  {32'h403e325f, 32'hbf76dea1} /* (17, 2, 12) {real, imag} */,
  {32'h3fd1925d, 32'h3c24cf20} /* (17, 2, 11) {real, imag} */,
  {32'hbf983c3f, 32'h3f82ecd2} /* (17, 2, 10) {real, imag} */,
  {32'hc0bcb19f, 32'h3e5ccec0} /* (17, 2, 9) {real, imag} */,
  {32'hbe95c399, 32'hbfdac70a} /* (17, 2, 8) {real, imag} */,
  {32'hc0bac8aa, 32'h4009fe02} /* (17, 2, 7) {real, imag} */,
  {32'hc0f3dd5c, 32'hbfd2ccb2} /* (17, 2, 6) {real, imag} */,
  {32'hc0229c34, 32'hc0ecfcf4} /* (17, 2, 5) {real, imag} */,
  {32'h4024cbdb, 32'hc02457a3} /* (17, 2, 4) {real, imag} */,
  {32'hbf9ac4da, 32'hc047143b} /* (17, 2, 3) {real, imag} */,
  {32'hbe585588, 32'hc0881ada} /* (17, 2, 2) {real, imag} */,
  {32'h405ddcbc, 32'h3fcdbd5c} /* (17, 2, 1) {real, imag} */,
  {32'h3fbe87e9, 32'h403766e9} /* (17, 2, 0) {real, imag} */,
  {32'hc0b04b4e, 32'h401603f2} /* (17, 1, 31) {real, imag} */,
  {32'hc0726553, 32'h40337b75} /* (17, 1, 30) {real, imag} */,
  {32'h3f9e628c, 32'h41049f92} /* (17, 1, 29) {real, imag} */,
  {32'hbfd50b90, 32'h409a088e} /* (17, 1, 28) {real, imag} */,
  {32'h4060479b, 32'h405c90d8} /* (17, 1, 27) {real, imag} */,
  {32'h41091e84, 32'h3fd1fce9} /* (17, 1, 26) {real, imag} */,
  {32'h400a3258, 32'h404a437c} /* (17, 1, 25) {real, imag} */,
  {32'h3fe6e1b2, 32'h408e3d52} /* (17, 1, 24) {real, imag} */,
  {32'h40f10b24, 32'hbec1605c} /* (17, 1, 23) {real, imag} */,
  {32'h411a52a8, 32'hc12f7a34} /* (17, 1, 22) {real, imag} */,
  {32'h4066c540, 32'hc099e164} /* (17, 1, 21) {real, imag} */,
  {32'hc06c0376, 32'h3f0251a2} /* (17, 1, 20) {real, imag} */,
  {32'hc0393acb, 32'h400b6022} /* (17, 1, 19) {real, imag} */,
  {32'hc04688dc, 32'h4108d2b6} /* (17, 1, 18) {real, imag} */,
  {32'hc097d76a, 32'h40ee50d0} /* (17, 1, 17) {real, imag} */,
  {32'hc08e1ac4, 32'h40773223} /* (17, 1, 16) {real, imag} */,
  {32'hc012310c, 32'hc0049f74} /* (17, 1, 15) {real, imag} */,
  {32'hbf4cabca, 32'h40023f45} /* (17, 1, 14) {real, imag} */,
  {32'hbfc1c8c2, 32'h4007343b} /* (17, 1, 13) {real, imag} */,
  {32'hc12e85d7, 32'h408560da} /* (17, 1, 12) {real, imag} */,
  {32'hc122b57c, 32'h3f0530e8} /* (17, 1, 11) {real, imag} */,
  {32'hc0bcad47, 32'hc09d6d0c} /* (17, 1, 10) {real, imag} */,
  {32'hbf02e02c, 32'hc0b83333} /* (17, 1, 9) {real, imag} */,
  {32'h40adf0e4, 32'h3f35bfe4} /* (17, 1, 8) {real, imag} */,
  {32'hc070b976, 32'h3d971d40} /* (17, 1, 7) {real, imag} */,
  {32'hc030ab10, 32'hbf85e86f} /* (17, 1, 6) {real, imag} */,
  {32'h4080b382, 32'h3fc66730} /* (17, 1, 5) {real, imag} */,
  {32'h40d1612b, 32'h408d16e5} /* (17, 1, 4) {real, imag} */,
  {32'h40c09228, 32'h405c6b7c} /* (17, 1, 3) {real, imag} */,
  {32'h405e8432, 32'hc0208cbf} /* (17, 1, 2) {real, imag} */,
  {32'h4069af97, 32'hc117ab48} /* (17, 1, 1) {real, imag} */,
  {32'h4008231a, 32'hc0d5d816} /* (17, 1, 0) {real, imag} */,
  {32'hc07cbe2f, 32'h40d7fcfe} /* (17, 0, 31) {real, imag} */,
  {32'hc03020af, 32'h3fafb8fa} /* (17, 0, 30) {real, imag} */,
  {32'h40150b14, 32'hc0d7ebd1} /* (17, 0, 29) {real, imag} */,
  {32'h4111c5c0, 32'hc0845697} /* (17, 0, 28) {real, imag} */,
  {32'h40029880, 32'hbf9ac18e} /* (17, 0, 27) {real, imag} */,
  {32'hbfb008a7, 32'hbfa41d64} /* (17, 0, 26) {real, imag} */,
  {32'h3f954601, 32'hc0dbfc4e} /* (17, 0, 25) {real, imag} */,
  {32'h3f3dc061, 32'h401a769d} /* (17, 0, 24) {real, imag} */,
  {32'hbfd5120e, 32'h40e463a2} /* (17, 0, 23) {real, imag} */,
  {32'h3f884994, 32'h3e967bcd} /* (17, 0, 22) {real, imag} */,
  {32'h4093120e, 32'hc0104519} /* (17, 0, 21) {real, imag} */,
  {32'h40e61a87, 32'hc076de63} /* (17, 0, 20) {real, imag} */,
  {32'h408c3ed2, 32'h3fd222f9} /* (17, 0, 19) {real, imag} */,
  {32'h3f979550, 32'hc10c4cac} /* (17, 0, 18) {real, imag} */,
  {32'hbfd27d80, 32'hc118d0be} /* (17, 0, 17) {real, imag} */,
  {32'h40264907, 32'hc0326d5c} /* (17, 0, 16) {real, imag} */,
  {32'h402eed89, 32'hc09f5c1e} /* (17, 0, 15) {real, imag} */,
  {32'h40222a68, 32'hc0379712} /* (17, 0, 14) {real, imag} */,
  {32'h3ff0c21d, 32'hc0a1e7dc} /* (17, 0, 13) {real, imag} */,
  {32'hc0669d88, 32'hbf1c0596} /* (17, 0, 12) {real, imag} */,
  {32'hc021aa68, 32'h3feaa9c9} /* (17, 0, 11) {real, imag} */,
  {32'hbf7e44a9, 32'h404db9ac} /* (17, 0, 10) {real, imag} */,
  {32'hc012630c, 32'h403b93f7} /* (17, 0, 9) {real, imag} */,
  {32'hc08f7d70, 32'h3dea9e40} /* (17, 0, 8) {real, imag} */,
  {32'hc0752d3a, 32'h3f32f214} /* (17, 0, 7) {real, imag} */,
  {32'hbf467b59, 32'hc0a47346} /* (17, 0, 6) {real, imag} */,
  {32'h40c1e3ca, 32'hbe5d6e88} /* (17, 0, 5) {real, imag} */,
  {32'h40622251, 32'h4026a102} /* (17, 0, 4) {real, imag} */,
  {32'h3fe1504d, 32'h3f98524c} /* (17, 0, 3) {real, imag} */,
  {32'hbefc18ac, 32'h3f9dd5f6} /* (17, 0, 2) {real, imag} */,
  {32'hc071c0f1, 32'h40419749} /* (17, 0, 1) {real, imag} */,
  {32'hbfbc054a, 32'h40761090} /* (17, 0, 0) {real, imag} */,
  {32'hbfef768c, 32'hc015409f} /* (16, 31, 31) {real, imag} */,
  {32'hbfabcd45, 32'hc0e576ca} /* (16, 31, 30) {real, imag} */,
  {32'hc0816088, 32'hc07d9be4} /* (16, 31, 29) {real, imag} */,
  {32'hbfbb9008, 32'hc0341764} /* (16, 31, 28) {real, imag} */,
  {32'h406344f4, 32'hbf88afeb} /* (16, 31, 27) {real, imag} */,
  {32'h3fd61d7c, 32'h40105b66} /* (16, 31, 26) {real, imag} */,
  {32'h4037e3d6, 32'h408bca2a} /* (16, 31, 25) {real, imag} */,
  {32'h406963b7, 32'h40f74906} /* (16, 31, 24) {real, imag} */,
  {32'hbe899002, 32'h4044349c} /* (16, 31, 23) {real, imag} */,
  {32'h3f83972b, 32'hc0a9ae34} /* (16, 31, 22) {real, imag} */,
  {32'h3efd86e0, 32'hbf251cfe} /* (16, 31, 21) {real, imag} */,
  {32'hbfa13818, 32'hbe26ecd0} /* (16, 31, 20) {real, imag} */,
  {32'hbed6f1aa, 32'h3ee3aa12} /* (16, 31, 19) {real, imag} */,
  {32'hbf597ed6, 32'h405e021a} /* (16, 31, 18) {real, imag} */,
  {32'hc01f2ab2, 32'h3fdbb298} /* (16, 31, 17) {real, imag} */,
  {32'hc083316e, 32'hc084ef0a} /* (16, 31, 16) {real, imag} */,
  {32'h3e915c20, 32'hc032f13c} /* (16, 31, 15) {real, imag} */,
  {32'h3f9f3290, 32'hbeb7be9c} /* (16, 31, 14) {real, imag} */,
  {32'h3ea25cb0, 32'h40048cd8} /* (16, 31, 13) {real, imag} */,
  {32'h40ff49ae, 32'h3fd2f378} /* (16, 31, 12) {real, imag} */,
  {32'h40bdb6f4, 32'h407a6260} /* (16, 31, 11) {real, imag} */,
  {32'h3fa08cc4, 32'h404e5cff} /* (16, 31, 10) {real, imag} */,
  {32'hbfc6eb1c, 32'h3fbcc556} /* (16, 31, 9) {real, imag} */,
  {32'hc01a341a, 32'h40851d50} /* (16, 31, 8) {real, imag} */,
  {32'h4045f472, 32'h40802fe7} /* (16, 31, 7) {real, imag} */,
  {32'h400082bd, 32'h3f8fdec7} /* (16, 31, 6) {real, imag} */,
  {32'h409922b9, 32'h3f7615d7} /* (16, 31, 5) {real, imag} */,
  {32'h40db3c74, 32'hbe46df34} /* (16, 31, 4) {real, imag} */,
  {32'h3fa56716, 32'h3f79d241} /* (16, 31, 3) {real, imag} */,
  {32'h40581a77, 32'hbffb1df7} /* (16, 31, 2) {real, imag} */,
  {32'h4039f0a0, 32'hc022d3d5} /* (16, 31, 1) {real, imag} */,
  {32'hbfdc126c, 32'hbf8c6f43} /* (16, 31, 0) {real, imag} */,
  {32'h3f9fd2a0, 32'h3e96e502} /* (16, 30, 31) {real, imag} */,
  {32'h3eb17bd8, 32'hbfce2d1c} /* (16, 30, 30) {real, imag} */,
  {32'hbf7b8426, 32'hbfb719da} /* (16, 30, 29) {real, imag} */,
  {32'h3eccc890, 32'hc02f138a} /* (16, 30, 28) {real, imag} */,
  {32'hbf2d0c20, 32'hc0f31997} /* (16, 30, 27) {real, imag} */,
  {32'h404026f9, 32'hc060a98f} /* (16, 30, 26) {real, imag} */,
  {32'h3e9edd54, 32'h3fedb9c4} /* (16, 30, 25) {real, imag} */,
  {32'h3db47920, 32'h3e0e09da} /* (16, 30, 24) {real, imag} */,
  {32'hbe291e70, 32'hbffcf4b8} /* (16, 30, 23) {real, imag} */,
  {32'h3e9d514c, 32'h3ff3aa82} /* (16, 30, 22) {real, imag} */,
  {32'h4049f021, 32'hbf07ecd4} /* (16, 30, 21) {real, imag} */,
  {32'h4018b6d4, 32'hc065395c} /* (16, 30, 20) {real, imag} */,
  {32'hc0510f1c, 32'h408f6d4c} /* (16, 30, 19) {real, imag} */,
  {32'h3fd3743a, 32'h40bdff28} /* (16, 30, 18) {real, imag} */,
  {32'h40182738, 32'hc05e25a4} /* (16, 30, 17) {real, imag} */,
  {32'h400cdc11, 32'hc0b19916} /* (16, 30, 16) {real, imag} */,
  {32'h404a7d6c, 32'hc0ae0ecd} /* (16, 30, 15) {real, imag} */,
  {32'h40b88aa5, 32'hbf817794} /* (16, 30, 14) {real, imag} */,
  {32'h3fadba24, 32'hbf48a415} /* (16, 30, 13) {real, imag} */,
  {32'hbff8f4b8, 32'h401e2e3a} /* (16, 30, 12) {real, imag} */,
  {32'h3eeb9d36, 32'h4058a3aa} /* (16, 30, 11) {real, imag} */,
  {32'hc0945b94, 32'h3fcf3cac} /* (16, 30, 10) {real, imag} */,
  {32'hbfd24578, 32'h408450f2} /* (16, 30, 9) {real, imag} */,
  {32'hbf611004, 32'h3f149b7c} /* (16, 30, 8) {real, imag} */,
  {32'hbf6979aa, 32'hc024484f} /* (16, 30, 7) {real, imag} */,
  {32'h400762f1, 32'h3f7fb14c} /* (16, 30, 6) {real, imag} */,
  {32'hbf3dc9c9, 32'h40a023ce} /* (16, 30, 5) {real, imag} */,
  {32'hbfcf0197, 32'h3f4186ba} /* (16, 30, 4) {real, imag} */,
  {32'hbd516180, 32'h3f8bc753} /* (16, 30, 3) {real, imag} */,
  {32'hc0c6a8d7, 32'h406d912f} /* (16, 30, 2) {real, imag} */,
  {32'hc03676b9, 32'hbfbbcd24} /* (16, 30, 1) {real, imag} */,
  {32'hbfd6c0d5, 32'hc059a6ab} /* (16, 30, 0) {real, imag} */,
  {32'hc069f49a, 32'hbd156bf8} /* (16, 29, 31) {real, imag} */,
  {32'hc09f7d2e, 32'hc05173aa} /* (16, 29, 30) {real, imag} */,
  {32'hc1037962, 32'hc00ba439} /* (16, 29, 29) {real, imag} */,
  {32'hc0c698ef, 32'h3fe72323} /* (16, 29, 28) {real, imag} */,
  {32'hbff34c8e, 32'h3fe32a7a} /* (16, 29, 27) {real, imag} */,
  {32'h4085fd8b, 32'h3df161e0} /* (16, 29, 26) {real, imag} */,
  {32'h4089b052, 32'h40206962} /* (16, 29, 25) {real, imag} */,
  {32'hbf5e976b, 32'hc07a324d} /* (16, 29, 24) {real, imag} */,
  {32'h4031e506, 32'hc087d4b2} /* (16, 29, 23) {real, imag} */,
  {32'hbe14c7bc, 32'hbf2b06a6} /* (16, 29, 22) {real, imag} */,
  {32'hc0510e50, 32'hc0a1b64d} /* (16, 29, 21) {real, imag} */,
  {32'hbf298510, 32'hbd921e68} /* (16, 29, 20) {real, imag} */,
  {32'h3ff5a25e, 32'h3fa92e93} /* (16, 29, 19) {real, imag} */,
  {32'h3fec27e8, 32'h40b6c8e7} /* (16, 29, 18) {real, imag} */,
  {32'h410263f6, 32'h40fdb19e} /* (16, 29, 17) {real, imag} */,
  {32'h40e36466, 32'h40f293c8} /* (16, 29, 16) {real, imag} */,
  {32'h40416c8c, 32'h403ae598} /* (16, 29, 15) {real, imag} */,
  {32'h3ee07330, 32'hbf8c515d} /* (16, 29, 14) {real, imag} */,
  {32'h3ff0a314, 32'h4002a08b} /* (16, 29, 13) {real, imag} */,
  {32'h40443fad, 32'h3fee4903} /* (16, 29, 12) {real, imag} */,
  {32'hbe92ce9c, 32'h4096b958} /* (16, 29, 11) {real, imag} */,
  {32'hc01f6b42, 32'hc005d2ce} /* (16, 29, 10) {real, imag} */,
  {32'hc048c97e, 32'hc0b81e08} /* (16, 29, 9) {real, imag} */,
  {32'h3f572e6a, 32'hbf5f905a} /* (16, 29, 8) {real, imag} */,
  {32'hbf79ba19, 32'h3fc372bf} /* (16, 29, 7) {real, imag} */,
  {32'h3f9014a8, 32'hc09ae079} /* (16, 29, 6) {real, imag} */,
  {32'hbf756298, 32'h3db54248} /* (16, 29, 5) {real, imag} */,
  {32'hbe53f3fc, 32'hbf120640} /* (16, 29, 4) {real, imag} */,
  {32'h3fdf9c04, 32'hbf92b1ec} /* (16, 29, 3) {real, imag} */,
  {32'hc07df846, 32'hbf81e5ae} /* (16, 29, 2) {real, imag} */,
  {32'hc0b97d2f, 32'hc07e7242} /* (16, 29, 1) {real, imag} */,
  {32'hc088a1c2, 32'h3e671ae7} /* (16, 29, 0) {real, imag} */,
  {32'h3ebd9542, 32'h3e675bb0} /* (16, 28, 31) {real, imag} */,
  {32'hc071968d, 32'h408503c1} /* (16, 28, 30) {real, imag} */,
  {32'h3eab1b79, 32'h40c398ec} /* (16, 28, 29) {real, imag} */,
  {32'h3fafabae, 32'h403ad8ee} /* (16, 28, 28) {real, imag} */,
  {32'h3fe5fb29, 32'h4030943c} /* (16, 28, 27) {real, imag} */,
  {32'h407725cf, 32'hc0a4fa02} /* (16, 28, 26) {real, imag} */,
  {32'h4044afde, 32'hc03c95b4} /* (16, 28, 25) {real, imag} */,
  {32'h4003f723, 32'h40f99c4a} /* (16, 28, 24) {real, imag} */,
  {32'hc0a2afcc, 32'h40f1d3d2} /* (16, 28, 23) {real, imag} */,
  {32'h3fbe3ab3, 32'h400293fb} /* (16, 28, 22) {real, imag} */,
  {32'h4029a040, 32'hc0018fe7} /* (16, 28, 21) {real, imag} */,
  {32'hbfdb7b5a, 32'hc0ab2025} /* (16, 28, 20) {real, imag} */,
  {32'hbfcedff9, 32'hc0c5d144} /* (16, 28, 19) {real, imag} */,
  {32'h3fe8b55a, 32'hbfdac988} /* (16, 28, 18) {real, imag} */,
  {32'hc06f3d83, 32'hc0c63df3} /* (16, 28, 17) {real, imag} */,
  {32'hc0616208, 32'hbf94ca00} /* (16, 28, 16) {real, imag} */,
  {32'hc0ba8e53, 32'hbe41e9f0} /* (16, 28, 15) {real, imag} */,
  {32'hc0298567, 32'hc0711b16} /* (16, 28, 14) {real, imag} */,
  {32'hbdf0cef0, 32'hc0c4feb4} /* (16, 28, 13) {real, imag} */,
  {32'hbec87a56, 32'hbfcf2de4} /* (16, 28, 12) {real, imag} */,
  {32'hbf69bc7d, 32'h4023278f} /* (16, 28, 11) {real, imag} */,
  {32'h3fc35b6a, 32'h3f251aca} /* (16, 28, 10) {real, imag} */,
  {32'h3fe937c8, 32'h4017982e} /* (16, 28, 9) {real, imag} */,
  {32'hc076cc8c, 32'h40e7a1aa} /* (16, 28, 8) {real, imag} */,
  {32'hc0131036, 32'h40a35826} /* (16, 28, 7) {real, imag} */,
  {32'hc0add5a2, 32'h40d30c84} /* (16, 28, 6) {real, imag} */,
  {32'hc0845f15, 32'h4081af1e} /* (16, 28, 5) {real, imag} */,
  {32'hbf7dbe6f, 32'hbd86ee28} /* (16, 28, 4) {real, imag} */,
  {32'h4064965d, 32'hc0122670} /* (16, 28, 3) {real, imag} */,
  {32'hbf8e20a5, 32'h3f888797} /* (16, 28, 2) {real, imag} */,
  {32'hbf18b514, 32'h3e93be22} /* (16, 28, 1) {real, imag} */,
  {32'hbe31580a, 32'hbf57257d} /* (16, 28, 0) {real, imag} */,
  {32'hbdbdb638, 32'hbfe4f025} /* (16, 27, 31) {real, imag} */,
  {32'hc080867e, 32'h3da8eae0} /* (16, 27, 30) {real, imag} */,
  {32'hbf1a6a71, 32'h4075a997} /* (16, 27, 29) {real, imag} */,
  {32'hbfcc907b, 32'h3efaa5ac} /* (16, 27, 28) {real, imag} */,
  {32'hc0548b48, 32'h3f937ca5} /* (16, 27, 27) {real, imag} */,
  {32'hc0169dde, 32'h3fa67515} /* (16, 27, 26) {real, imag} */,
  {32'h3def4574, 32'h404bd5c8} /* (16, 27, 25) {real, imag} */,
  {32'h3fb62f4d, 32'h408260fa} /* (16, 27, 24) {real, imag} */,
  {32'h4011b910, 32'h4084169a} /* (16, 27, 23) {real, imag} */,
  {32'hbe914cf8, 32'h3fdb1429} /* (16, 27, 22) {real, imag} */,
  {32'h3f79e72a, 32'hbff1beb8} /* (16, 27, 21) {real, imag} */,
  {32'h40a79f12, 32'hbe484148} /* (16, 27, 20) {real, imag} */,
  {32'h4013a4c7, 32'hbfeab243} /* (16, 27, 19) {real, imag} */,
  {32'h3f08cf3c, 32'hbe275c94} /* (16, 27, 18) {real, imag} */,
  {32'h4073cd62, 32'hbeb42ccc} /* (16, 27, 17) {real, imag} */,
  {32'hbfc35642, 32'h3f988d7f} /* (16, 27, 16) {real, imag} */,
  {32'hc0bc94ce, 32'h3f3b6eae} /* (16, 27, 15) {real, imag} */,
  {32'hc0aa656f, 32'hbfec82a2} /* (16, 27, 14) {real, imag} */,
  {32'hc06c3706, 32'hc06bb2be} /* (16, 27, 13) {real, imag} */,
  {32'h3ff82019, 32'hc0081454} /* (16, 27, 12) {real, imag} */,
  {32'h3f833cff, 32'hbd3827d0} /* (16, 27, 11) {real, imag} */,
  {32'h4011fa8b, 32'h401bb63c} /* (16, 27, 10) {real, imag} */,
  {32'h409dbdfa, 32'h4021d7f2} /* (16, 27, 9) {real, imag} */,
  {32'h4008ec43, 32'h4096d14e} /* (16, 27, 8) {real, imag} */,
  {32'hbf664b76, 32'h3fbfc8f8} /* (16, 27, 7) {real, imag} */,
  {32'hbfbbcd96, 32'h3f907563} /* (16, 27, 6) {real, imag} */,
  {32'hc039ba70, 32'h4040b4d5} /* (16, 27, 5) {real, imag} */,
  {32'h3d88d5dc, 32'h409026ba} /* (16, 27, 4) {real, imag} */,
  {32'h3eb299a8, 32'h40aa799e} /* (16, 27, 3) {real, imag} */,
  {32'h3f2b92a2, 32'h406b008a} /* (16, 27, 2) {real, imag} */,
  {32'hbfc3cd85, 32'hbfcd9527} /* (16, 27, 1) {real, imag} */,
  {32'hbee7d7cc, 32'hc03e49ae} /* (16, 27, 0) {real, imag} */,
  {32'hc0764708, 32'h40304cf4} /* (16, 26, 31) {real, imag} */,
  {32'hc0537c6e, 32'h4092d34a} /* (16, 26, 30) {real, imag} */,
  {32'hbffd0743, 32'h4083f259} /* (16, 26, 29) {real, imag} */,
  {32'hc08a6000, 32'h3f5d950f} /* (16, 26, 28) {real, imag} */,
  {32'hbe197b10, 32'h3f5a5ee0} /* (16, 26, 27) {real, imag} */,
  {32'hc01234fe, 32'h3e79fec4} /* (16, 26, 26) {real, imag} */,
  {32'hbf8ee2bd, 32'h3fa1d60a} /* (16, 26, 25) {real, imag} */,
  {32'hbeb0b09e, 32'h3eb730dc} /* (16, 26, 24) {real, imag} */,
  {32'hc01c7865, 32'h4049f57c} /* (16, 26, 23) {real, imag} */,
  {32'hbeca20cc, 32'hbdd6e894} /* (16, 26, 22) {real, imag} */,
  {32'h4047148e, 32'hbfc6c242} /* (16, 26, 21) {real, imag} */,
  {32'h3fa548ed, 32'hbe8aa6b5} /* (16, 26, 20) {real, imag} */,
  {32'h3f5f0f4e, 32'hc0482e3a} /* (16, 26, 19) {real, imag} */,
  {32'h3f6a3fc6, 32'hbf813d22} /* (16, 26, 18) {real, imag} */,
  {32'h40169291, 32'h402e8e5a} /* (16, 26, 17) {real, imag} */,
  {32'h402c7097, 32'h3f1a67a0} /* (16, 26, 16) {real, imag} */,
  {32'h3fde0fa8, 32'h3f7df728} /* (16, 26, 15) {real, imag} */,
  {32'hbf5038bc, 32'hbe2e79a4} /* (16, 26, 14) {real, imag} */,
  {32'h3fe10e25, 32'hc04249c7} /* (16, 26, 13) {real, imag} */,
  {32'h40a5c7dd, 32'hc04b4544} /* (16, 26, 12) {real, imag} */,
  {32'hbd2aade0, 32'hbf9152eb} /* (16, 26, 11) {real, imag} */,
  {32'hc08ccbb4, 32'h3d485c00} /* (16, 26, 10) {real, imag} */,
  {32'h3e906574, 32'hbf8c9cc9} /* (16, 26, 9) {real, imag} */,
  {32'h4096a704, 32'hbeb0c6b8} /* (16, 26, 8) {real, imag} */,
  {32'h3f94b846, 32'h40255646} /* (16, 26, 7) {real, imag} */,
  {32'h3f8ac2bf, 32'h40d1a568} /* (16, 26, 6) {real, imag} */,
  {32'hbdde4fc0, 32'h40b9b7d8} /* (16, 26, 5) {real, imag} */,
  {32'h3fdbc58b, 32'h40e50826} /* (16, 26, 4) {real, imag} */,
  {32'h4018fc20, 32'h409db47b} /* (16, 26, 3) {real, imag} */,
  {32'h3eb78688, 32'hc016ad56} /* (16, 26, 2) {real, imag} */,
  {32'hc01b5b28, 32'hc08400a2} /* (16, 26, 1) {real, imag} */,
  {32'hbf841638, 32'h400ab261} /* (16, 26, 0) {real, imag} */,
  {32'h3ec5f2da, 32'hc07a2e2b} /* (16, 25, 31) {real, imag} */,
  {32'h400e7ab6, 32'hc04e3105} /* (16, 25, 30) {real, imag} */,
  {32'h407ce3ae, 32'h40077340} /* (16, 25, 29) {real, imag} */,
  {32'h3e184290, 32'h4068b145} /* (16, 25, 28) {real, imag} */,
  {32'hbf7921c4, 32'h3f6920b2} /* (16, 25, 27) {real, imag} */,
  {32'h3fc384fc, 32'h3dbb5a24} /* (16, 25, 26) {real, imag} */,
  {32'h3fcc3793, 32'h3e9e232e} /* (16, 25, 25) {real, imag} */,
  {32'h3d25d0c0, 32'hbfb1ef0d} /* (16, 25, 24) {real, imag} */,
  {32'hbf35cdb1, 32'hbed62f0c} /* (16, 25, 23) {real, imag} */,
  {32'hbf1cd3ec, 32'h3f04bb2a} /* (16, 25, 22) {real, imag} */,
  {32'h4081420d, 32'hbd8f9e40} /* (16, 25, 21) {real, imag} */,
  {32'h40108827, 32'hc005f41a} /* (16, 25, 20) {real, imag} */,
  {32'hbeeab028, 32'hbf4742e8} /* (16, 25, 19) {real, imag} */,
  {32'h3e5332a0, 32'hbf35cdbf} /* (16, 25, 18) {real, imag} */,
  {32'hbf9385f0, 32'hbf360c12} /* (16, 25, 17) {real, imag} */,
  {32'hbf2af650, 32'hbe00767e} /* (16, 25, 16) {real, imag} */,
  {32'h3f2b9e8a, 32'h3f9342c8} /* (16, 25, 15) {real, imag} */,
  {32'hc0138f22, 32'hc0902cd9} /* (16, 25, 14) {real, imag} */,
  {32'hc0656214, 32'hc08a618d} /* (16, 25, 13) {real, imag} */,
  {32'h3f86430b, 32'hc06b1964} /* (16, 25, 12) {real, imag} */,
  {32'h40188ff9, 32'hc01082cd} /* (16, 25, 11) {real, imag} */,
  {32'hbff432b4, 32'hbfbc842c} /* (16, 25, 10) {real, imag} */,
  {32'hbffee8f8, 32'hbfc9a566} /* (16, 25, 9) {real, imag} */,
  {32'hbfc271c0, 32'hbfaf36e2} /* (16, 25, 8) {real, imag} */,
  {32'h3ee8b676, 32'hbe98b3a0} /* (16, 25, 7) {real, imag} */,
  {32'h3fec8c8a, 32'hbf02cf7b} /* (16, 25, 6) {real, imag} */,
  {32'h406d296c, 32'hbff03827} /* (16, 25, 5) {real, imag} */,
  {32'h400148e8, 32'h3fa54a2c} /* (16, 25, 4) {real, imag} */,
  {32'hbfa28b3c, 32'h40155d31} /* (16, 25, 3) {real, imag} */,
  {32'hbdd2bef0, 32'hbe9d0c20} /* (16, 25, 2) {real, imag} */,
  {32'hc0107bd4, 32'hc013732c} /* (16, 25, 1) {real, imag} */,
  {32'hc06280f6, 32'hc046a322} /* (16, 25, 0) {real, imag} */,
  {32'hbf92c480, 32'hbf33c2f6} /* (16, 24, 31) {real, imag} */,
  {32'hbfc42048, 32'hbf960228} /* (16, 24, 30) {real, imag} */,
  {32'h3ee21602, 32'hc0ade1ee} /* (16, 24, 29) {real, imag} */,
  {32'h409fe4d5, 32'hc0e726da} /* (16, 24, 28) {real, imag} */,
  {32'h40dbcc38, 32'hc0909820} /* (16, 24, 27) {real, imag} */,
  {32'h3fbeea7f, 32'h3efd8194} /* (16, 24, 26) {real, imag} */,
  {32'hbf5a94b4, 32'h3fedf14b} /* (16, 24, 25) {real, imag} */,
  {32'hbf998346, 32'hbf090778} /* (16, 24, 24) {real, imag} */,
  {32'hc07651ed, 32'hc015218b} /* (16, 24, 23) {real, imag} */,
  {32'hc08c6a44, 32'hc073a21a} /* (16, 24, 22) {real, imag} */,
  {32'hbf94d570, 32'hbe6b9570} /* (16, 24, 21) {real, imag} */,
  {32'hc03b9c16, 32'h3eae266e} /* (16, 24, 20) {real, imag} */,
  {32'hc054e0f4, 32'hbfdde60c} /* (16, 24, 19) {real, imag} */,
  {32'hbf442028, 32'h4049001b} /* (16, 24, 18) {real, imag} */,
  {32'h3f632bd3, 32'h409ea006} /* (16, 24, 17) {real, imag} */,
  {32'hbf1ceb9a, 32'h40b12c28} /* (16, 24, 16) {real, imag} */,
  {32'hbf3fc0de, 32'h4027eacd} /* (16, 24, 15) {real, imag} */,
  {32'h3f5e8268, 32'h3f592ad4} /* (16, 24, 14) {real, imag} */,
  {32'h40576de5, 32'h3e334724} /* (16, 24, 13) {real, imag} */,
  {32'hc02e88d0, 32'h3f81cc3d} /* (16, 24, 12) {real, imag} */,
  {32'hbdb12568, 32'h4011ea9e} /* (16, 24, 11) {real, imag} */,
  {32'hbe9842d0, 32'h3fa9c6a8} /* (16, 24, 10) {real, imag} */,
  {32'h3e99b858, 32'h4064daed} /* (16, 24, 9) {real, imag} */,
  {32'h3f8f74d6, 32'h3fbc385a} /* (16, 24, 8) {real, imag} */,
  {32'h3fff461a, 32'hbfa6ae4f} /* (16, 24, 7) {real, imag} */,
  {32'h3fe62333, 32'h3f400fef} /* (16, 24, 6) {real, imag} */,
  {32'hbe567b44, 32'h404e3da6} /* (16, 24, 5) {real, imag} */,
  {32'hc0337198, 32'hbf62ca9d} /* (16, 24, 4) {real, imag} */,
  {32'hbfddb6a8, 32'hc05b6d60} /* (16, 24, 3) {real, imag} */,
  {32'h3f26b76c, 32'hc0421eec} /* (16, 24, 2) {real, imag} */,
  {32'hbfde41f5, 32'hbfa93050} /* (16, 24, 1) {real, imag} */,
  {32'hc00f17f6, 32'hbf8828be} /* (16, 24, 0) {real, imag} */,
  {32'h3fc309ae, 32'hbfc101a2} /* (16, 23, 31) {real, imag} */,
  {32'h3fd13fc7, 32'hbfacc426} /* (16, 23, 30) {real, imag} */,
  {32'hc03f206e, 32'hc0448446} /* (16, 23, 29) {real, imag} */,
  {32'hbfbda444, 32'hbfb52146} /* (16, 23, 28) {real, imag} */,
  {32'h40565b53, 32'h3e587fba} /* (16, 23, 27) {real, imag} */,
  {32'h3fc2592a, 32'h3e48512e} /* (16, 23, 26) {real, imag} */,
  {32'hbf985f69, 32'hbef19a2a} /* (16, 23, 25) {real, imag} */,
  {32'hc01c3235, 32'hbfdc9ca9} /* (16, 23, 24) {real, imag} */,
  {32'hbf2176a5, 32'hc07786d0} /* (16, 23, 23) {real, imag} */,
  {32'h3d8d0000, 32'hc027ae72} /* (16, 23, 22) {real, imag} */,
  {32'hbf56fc6e, 32'hbf23f790} /* (16, 23, 21) {real, imag} */,
  {32'hbfaa4076, 32'h3ea9251c} /* (16, 23, 20) {real, imag} */,
  {32'h40343190, 32'hbef250dc} /* (16, 23, 19) {real, imag} */,
  {32'hbf00e634, 32'hbff53efa} /* (16, 23, 18) {real, imag} */,
  {32'hc03250c2, 32'hbdc874cc} /* (16, 23, 17) {real, imag} */,
  {32'hbfdcfa64, 32'hbf4e4928} /* (16, 23, 16) {real, imag} */,
  {32'hbe951d2e, 32'hbec7526a} /* (16, 23, 15) {real, imag} */,
  {32'h3fe557a8, 32'h404c88a3} /* (16, 23, 14) {real, imag} */,
  {32'hbf00f746, 32'hbed77be0} /* (16, 23, 13) {real, imag} */,
  {32'hbfda1b77, 32'h3f5355f8} /* (16, 23, 12) {real, imag} */,
  {32'h4065b601, 32'hbe785380} /* (16, 23, 11) {real, imag} */,
  {32'h401b2054, 32'h40766d4e} /* (16, 23, 10) {real, imag} */,
  {32'hbe31d650, 32'h40050dd7} /* (16, 23, 9) {real, imag} */,
  {32'hbcb04800, 32'h406f2223} /* (16, 23, 8) {real, imag} */,
  {32'h3f68530f, 32'h40a9195d} /* (16, 23, 7) {real, imag} */,
  {32'h3fe3e0fc, 32'h3f172aa1} /* (16, 23, 6) {real, imag} */,
  {32'hbd40ecc0, 32'h3ef646e4} /* (16, 23, 5) {real, imag} */,
  {32'h3f47d018, 32'hc05b6a3e} /* (16, 23, 4) {real, imag} */,
  {32'hbfaf31c2, 32'hc09a4078} /* (16, 23, 3) {real, imag} */,
  {32'hbfc91dd1, 32'hc088b52c} /* (16, 23, 2) {real, imag} */,
  {32'h3faf2af6, 32'hc089328f} /* (16, 23, 1) {real, imag} */,
  {32'hbfc775fc, 32'hc0962d39} /* (16, 23, 0) {real, imag} */,
  {32'hbf196fc8, 32'h3f7989a8} /* (16, 22, 31) {real, imag} */,
  {32'h3ebc7038, 32'h3e8c1a38} /* (16, 22, 30) {real, imag} */,
  {32'h3f3ecf12, 32'h3fbe38f9} /* (16, 22, 29) {real, imag} */,
  {32'hbf17bc44, 32'hbfa9fa40} /* (16, 22, 28) {real, imag} */,
  {32'h40086062, 32'hbf1d9db4} /* (16, 22, 27) {real, imag} */,
  {32'h40803b63, 32'h3fb2f19a} /* (16, 22, 26) {real, imag} */,
  {32'h404df57e, 32'hbfb3ad38} /* (16, 22, 25) {real, imag} */,
  {32'hbf25a602, 32'h3f47a836} /* (16, 22, 24) {real, imag} */,
  {32'hc02cb023, 32'h4035ca04} /* (16, 22, 23) {real, imag} */,
  {32'hc0119a54, 32'h3f1cc0b0} /* (16, 22, 22) {real, imag} */,
  {32'hbe5a1d38, 32'hbf36fd74} /* (16, 22, 21) {real, imag} */,
  {32'h3febfe31, 32'hbeda3715} /* (16, 22, 20) {real, imag} */,
  {32'h3fca9065, 32'h3d0efd80} /* (16, 22, 19) {real, imag} */,
  {32'hbe8da374, 32'hc0057af7} /* (16, 22, 18) {real, imag} */,
  {32'h3f28a495, 32'h3f5e3ad0} /* (16, 22, 17) {real, imag} */,
  {32'h3fd8d98e, 32'h401f8c42} /* (16, 22, 16) {real, imag} */,
  {32'h4045e130, 32'h4025df3b} /* (16, 22, 15) {real, imag} */,
  {32'h40651dad, 32'h3fba5656} /* (16, 22, 14) {real, imag} */,
  {32'h40374826, 32'h3e4735b0} /* (16, 22, 13) {real, imag} */,
  {32'h4027222c, 32'h3e592858} /* (16, 22, 12) {real, imag} */,
  {32'h400c1772, 32'h3f8c4ec5} /* (16, 22, 11) {real, imag} */,
  {32'h3fe5e43c, 32'hbff92848} /* (16, 22, 10) {real, imag} */,
  {32'h4018aa96, 32'h4029d0b2} /* (16, 22, 9) {real, imag} */,
  {32'h400feb65, 32'h40885258} /* (16, 22, 8) {real, imag} */,
  {32'hbfc3de92, 32'h3cf6ebc0} /* (16, 22, 7) {real, imag} */,
  {32'h3f9022ed, 32'h3ea873e8} /* (16, 22, 6) {real, imag} */,
  {32'h4037b196, 32'h3f283d40} /* (16, 22, 5) {real, imag} */,
  {32'h402aa83e, 32'h3fa376c0} /* (16, 22, 4) {real, imag} */,
  {32'h40379ec8, 32'h400caab4} /* (16, 22, 3) {real, imag} */,
  {32'hbf3ad014, 32'hbdf838f0} /* (16, 22, 2) {real, imag} */,
  {32'hc08dca55, 32'hbe56c4d0} /* (16, 22, 1) {real, imag} */,
  {32'hc018886f, 32'h3e2a7270} /* (16, 22, 0) {real, imag} */,
  {32'h3f9652be, 32'hbf92aecb} /* (16, 21, 31) {real, imag} */,
  {32'h3ea63698, 32'hbf168d74} /* (16, 21, 30) {real, imag} */,
  {32'h3f4b16d1, 32'h3fdf4832} /* (16, 21, 29) {real, imag} */,
  {32'h3ffa6b89, 32'h3fb2dff9} /* (16, 21, 28) {real, imag} */,
  {32'h3fa01db0, 32'h403e6aaa} /* (16, 21, 27) {real, imag} */,
  {32'hbf53058e, 32'h4035aa44} /* (16, 21, 26) {real, imag} */,
  {32'hbf68da2a, 32'h3d8554f0} /* (16, 21, 25) {real, imag} */,
  {32'hbff2d54b, 32'hbfbc4fa5} /* (16, 21, 24) {real, imag} */,
  {32'hbfe1f34c, 32'hbc972f80} /* (16, 21, 23) {real, imag} */,
  {32'hbec56108, 32'h3e3d7118} /* (16, 21, 22) {real, imag} */,
  {32'h3f68d772, 32'h3f83d970} /* (16, 21, 21) {real, imag} */,
  {32'h3ee85608, 32'h3fbb837e} /* (16, 21, 20) {real, imag} */,
  {32'h3ec3fee6, 32'hbef9c604} /* (16, 21, 19) {real, imag} */,
  {32'h40204ec3, 32'h3f8148a8} /* (16, 21, 18) {real, imag} */,
  {32'h3fd4acdc, 32'h3f150c26} /* (16, 21, 17) {real, imag} */,
  {32'h3fa029ea, 32'hbd828a70} /* (16, 21, 16) {real, imag} */,
  {32'h3f59e720, 32'h3f61e884} /* (16, 21, 15) {real, imag} */,
  {32'h3ea470e0, 32'h3f2cc7cc} /* (16, 21, 14) {real, imag} */,
  {32'hbe0cea68, 32'h40039c42} /* (16, 21, 13) {real, imag} */,
  {32'hc01ce3d4, 32'h400da9a6} /* (16, 21, 12) {real, imag} */,
  {32'hc04b2b8c, 32'h3fb8138c} /* (16, 21, 11) {real, imag} */,
  {32'hbfc05e68, 32'h3e0677f8} /* (16, 21, 10) {real, imag} */,
  {32'h400ebe64, 32'h3f0f5360} /* (16, 21, 9) {real, imag} */,
  {32'hbe8eb3c0, 32'h3fc420bf} /* (16, 21, 8) {real, imag} */,
  {32'hbe3fd1ba, 32'hbeef1daa} /* (16, 21, 7) {real, imag} */,
  {32'h3f8b619a, 32'h3fbac5cf} /* (16, 21, 6) {real, imag} */,
  {32'h3fcd0e20, 32'h3f93ce66} /* (16, 21, 5) {real, imag} */,
  {32'hbe6fabde, 32'hbdf3eae0} /* (16, 21, 4) {real, imag} */,
  {32'hc0333adb, 32'hc01acfb6} /* (16, 21, 3) {real, imag} */,
  {32'hc008a4ba, 32'hbf9776cd} /* (16, 21, 2) {real, imag} */,
  {32'hc005186c, 32'h3eb3c86c} /* (16, 21, 1) {real, imag} */,
  {32'hbe8a376c, 32'hbf9f4d7f} /* (16, 21, 0) {real, imag} */,
  {32'h3fcdc6f6, 32'h3e8e04a8} /* (16, 20, 31) {real, imag} */,
  {32'h3fe40ec6, 32'h4024b9c0} /* (16, 20, 30) {real, imag} */,
  {32'h3ea94343, 32'h3dadbde0} /* (16, 20, 29) {real, imag} */,
  {32'hbf06afcb, 32'hbfe312b4} /* (16, 20, 28) {real, imag} */,
  {32'hbee38ad4, 32'h3f9acab5} /* (16, 20, 27) {real, imag} */,
  {32'hbf99213e, 32'h4038669d} /* (16, 20, 26) {real, imag} */,
  {32'hbf928360, 32'hbf3a86d4} /* (16, 20, 25) {real, imag} */,
  {32'h3fc69a46, 32'hbee35120} /* (16, 20, 24) {real, imag} */,
  {32'h404d548d, 32'hbee7c7e0} /* (16, 20, 23) {real, imag} */,
  {32'h3fc9001b, 32'h3f9f3528} /* (16, 20, 22) {real, imag} */,
  {32'hbece7dac, 32'h403c7b4b} /* (16, 20, 21) {real, imag} */,
  {32'h3f02ad95, 32'h3d43aa80} /* (16, 20, 20) {real, imag} */,
  {32'h400c7d72, 32'h3e122740} /* (16, 20, 19) {real, imag} */,
  {32'h3f6671a3, 32'h3f1425f1} /* (16, 20, 18) {real, imag} */,
  {32'h3f6413c4, 32'hbe04a3e0} /* (16, 20, 17) {real, imag} */,
  {32'h40105858, 32'hbf1a4f73} /* (16, 20, 16) {real, imag} */,
  {32'h3fb541e4, 32'hc0585947} /* (16, 20, 15) {real, imag} */,
  {32'h3eee39d8, 32'hc035ec7c} /* (16, 20, 14) {real, imag} */,
  {32'h3f8c65ad, 32'h3f160694} /* (16, 20, 13) {real, imag} */,
  {32'h3eb9bc2e, 32'h3f28b8cb} /* (16, 20, 12) {real, imag} */,
  {32'h3df0b278, 32'h3fe3af72} /* (16, 20, 11) {real, imag} */,
  {32'h40514b9b, 32'h4009f2f0} /* (16, 20, 10) {real, imag} */,
  {32'h3fdd55d4, 32'h3fb3213c} /* (16, 20, 9) {real, imag} */,
  {32'h401de698, 32'hbec4e1a8} /* (16, 20, 8) {real, imag} */,
  {32'h3ffa8e14, 32'h3f1b2b20} /* (16, 20, 7) {real, imag} */,
  {32'hbc093800, 32'h3f41b4a0} /* (16, 20, 6) {real, imag} */,
  {32'h3fa76e04, 32'hbedf7308} /* (16, 20, 5) {real, imag} */,
  {32'hbf3d5c1d, 32'h3f7042f5} /* (16, 20, 4) {real, imag} */,
  {32'h3f57869c, 32'h403a2992} /* (16, 20, 3) {real, imag} */,
  {32'hbf6cd8a6, 32'h3fe1c28b} /* (16, 20, 2) {real, imag} */,
  {32'hbfc18218, 32'hbf92e150} /* (16, 20, 1) {real, imag} */,
  {32'hbe9d5673, 32'hc01c6506} /* (16, 20, 0) {real, imag} */,
  {32'h3ef48dac, 32'h3eb3005b} /* (16, 19, 31) {real, imag} */,
  {32'h3f68840c, 32'h3fcf30fc} /* (16, 19, 30) {real, imag} */,
  {32'h402fa71e, 32'h3e86eb76} /* (16, 19, 29) {real, imag} */,
  {32'h4017313a, 32'hbf9c2d03} /* (16, 19, 28) {real, imag} */,
  {32'hbf1d61e4, 32'hbf6d80c8} /* (16, 19, 27) {real, imag} */,
  {32'hbfb05da0, 32'h3faa078c} /* (16, 19, 26) {real, imag} */,
  {32'hc0195b98, 32'h3fc5ce71} /* (16, 19, 25) {real, imag} */,
  {32'h3f8e1db4, 32'h3fc239d2} /* (16, 19, 24) {real, imag} */,
  {32'h3fac41e4, 32'hbf532eac} /* (16, 19, 23) {real, imag} */,
  {32'h3f44c585, 32'hbfde39b9} /* (16, 19, 22) {real, imag} */,
  {32'h3fed678c, 32'h3fa59b74} /* (16, 19, 21) {real, imag} */,
  {32'h407476e6, 32'h3fe7cf54} /* (16, 19, 20) {real, imag} */,
  {32'h3fdd7fe6, 32'h3fbc02b9} /* (16, 19, 19) {real, imag} */,
  {32'h3d7ab370, 32'h3ddd8c40} /* (16, 19, 18) {real, imag} */,
  {32'hbf109228, 32'hbeeb6120} /* (16, 19, 17) {real, imag} */,
  {32'hbe83aca8, 32'h3e39f4d0} /* (16, 19, 16) {real, imag} */,
  {32'hbee46154, 32'h3f51beec} /* (16, 19, 15) {real, imag} */,
  {32'h3f182f70, 32'hbf476850} /* (16, 19, 14) {real, imag} */,
  {32'hbf1d150c, 32'hbf9fe252} /* (16, 19, 13) {real, imag} */,
  {32'hbf378dd4, 32'hbe927684} /* (16, 19, 12) {real, imag} */,
  {32'hbfa6881b, 32'h3f102f34} /* (16, 19, 11) {real, imag} */,
  {32'hbfdbb7fd, 32'hbee1a088} /* (16, 19, 10) {real, imag} */,
  {32'hc00094d6, 32'hbfb2db52} /* (16, 19, 9) {real, imag} */,
  {32'hc09188ed, 32'hc087f3ef} /* (16, 19, 8) {real, imag} */,
  {32'hc0226b91, 32'hc01a3f14} /* (16, 19, 7) {real, imag} */,
  {32'hbfc6ee66, 32'h3f2b6b70} /* (16, 19, 6) {real, imag} */,
  {32'hbebc4058, 32'hbf43b019} /* (16, 19, 5) {real, imag} */,
  {32'h3eb4c7e6, 32'hbf54ae48} /* (16, 19, 4) {real, imag} */,
  {32'hbf2727dc, 32'h3f13ca41} /* (16, 19, 3) {real, imag} */,
  {32'h3f800184, 32'hbed51dd0} /* (16, 19, 2) {real, imag} */,
  {32'h3fc711b8, 32'hbf380112} /* (16, 19, 1) {real, imag} */,
  {32'h3f60456a, 32'hbe163949} /* (16, 19, 0) {real, imag} */,
  {32'h3f650bf9, 32'hbfb223ec} /* (16, 18, 31) {real, imag} */,
  {32'h4011d02e, 32'hc031e266} /* (16, 18, 30) {real, imag} */,
  {32'h3f48a194, 32'hbf41fd74} /* (16, 18, 29) {real, imag} */,
  {32'h3f2f4f1a, 32'h3dd91c40} /* (16, 18, 28) {real, imag} */,
  {32'h3f1ef124, 32'hbd601780} /* (16, 18, 27) {real, imag} */,
  {32'h3e9cbd40, 32'hbf339044} /* (16, 18, 26) {real, imag} */,
  {32'h3faf35e8, 32'hbde97560} /* (16, 18, 25) {real, imag} */,
  {32'h3f445d4d, 32'h3ed2885d} /* (16, 18, 24) {real, imag} */,
  {32'h3fe04474, 32'hbfba71fe} /* (16, 18, 23) {real, imag} */,
  {32'h400b9dae, 32'hbf8128f2} /* (16, 18, 22) {real, imag} */,
  {32'h3ff27a3a, 32'hbf511de8} /* (16, 18, 21) {real, imag} */,
  {32'h3f207866, 32'h3f317780} /* (16, 18, 20) {real, imag} */,
  {32'h3f63a6c0, 32'h3f9cc4e2} /* (16, 18, 19) {real, imag} */,
  {32'h3dc15928, 32'h3fdbf4e8} /* (16, 18, 18) {real, imag} */,
  {32'hbee97c10, 32'h3f65f528} /* (16, 18, 17) {real, imag} */,
  {32'hbfc7bb02, 32'h3e934f18} /* (16, 18, 16) {real, imag} */,
  {32'h3db549f0, 32'hbfad459c} /* (16, 18, 15) {real, imag} */,
  {32'h4009ae30, 32'hbece17f4} /* (16, 18, 14) {real, imag} */,
  {32'h3ec2a289, 32'hbe81225e} /* (16, 18, 13) {real, imag} */,
  {32'hbf8c15ac, 32'hbf8fc132} /* (16, 18, 12) {real, imag} */,
  {32'h3f005f5f, 32'hbf9be75f} /* (16, 18, 11) {real, imag} */,
  {32'h3efccd70, 32'hbe8613a0} /* (16, 18, 10) {real, imag} */,
  {32'hbda7e580, 32'h3f34129e} /* (16, 18, 9) {real, imag} */,
  {32'h3ea15dd8, 32'h3f58c0c0} /* (16, 18, 8) {real, imag} */,
  {32'hbf0fcd56, 32'h3f156c34} /* (16, 18, 7) {real, imag} */,
  {32'h3d51cac0, 32'h3f7c5f08} /* (16, 18, 6) {real, imag} */,
  {32'h3e02d6ec, 32'h3ee1d9e0} /* (16, 18, 5) {real, imag} */,
  {32'hbf9709df, 32'hbeacee95} /* (16, 18, 4) {real, imag} */,
  {32'hbf768f70, 32'hbfa8eb45} /* (16, 18, 3) {real, imag} */,
  {32'hbe948c90, 32'hbdb861e0} /* (16, 18, 2) {real, imag} */,
  {32'hbefa5528, 32'h3f77c071} /* (16, 18, 1) {real, imag} */,
  {32'hbea50724, 32'h3f0868ac} /* (16, 18, 0) {real, imag} */,
  {32'hbf7b6d18, 32'hbd19c6c0} /* (16, 17, 31) {real, imag} */,
  {32'hbfa047e1, 32'h3f8062d6} /* (16, 17, 30) {real, imag} */,
  {32'hbfd71f07, 32'h3f86d23d} /* (16, 17, 29) {real, imag} */,
  {32'hbfba16ce, 32'h3ed3b0a4} /* (16, 17, 28) {real, imag} */,
  {32'hbeb8f910, 32'hbe32dc06} /* (16, 17, 27) {real, imag} */,
  {32'hbe61f350, 32'h3ef46044} /* (16, 17, 26) {real, imag} */,
  {32'hbf0ae676, 32'hbf5867ec} /* (16, 17, 25) {real, imag} */,
  {32'hbf1a5d64, 32'hbf8352a8} /* (16, 17, 24) {real, imag} */,
  {32'hbfa1bdbc, 32'hbf080b36} /* (16, 17, 23) {real, imag} */,
  {32'hbf8d1281, 32'hbdbf3700} /* (16, 17, 22) {real, imag} */,
  {32'hbf327e90, 32'h3f851b97} /* (16, 17, 21) {real, imag} */,
  {32'hbee0a5b6, 32'h3ecb016c} /* (16, 17, 20) {real, imag} */,
  {32'hbf29acaf, 32'h3e7bef6b} /* (16, 17, 19) {real, imag} */,
  {32'h3db2198c, 32'hbebdb8fc} /* (16, 17, 18) {real, imag} */,
  {32'hbf901198, 32'hbf136fcd} /* (16, 17, 17) {real, imag} */,
  {32'hbfce6f45, 32'h3e11bf40} /* (16, 17, 16) {real, imag} */,
  {32'hbfa7e09c, 32'h3e9457b4} /* (16, 17, 15) {real, imag} */,
  {32'hbfff4ebc, 32'h3f8b2e0b} /* (16, 17, 14) {real, imag} */,
  {32'hbf5ea558, 32'h3f8d32dd} /* (16, 17, 13) {real, imag} */,
  {32'h3f3a1fd4, 32'h3f5d7cc5} /* (16, 17, 12) {real, imag} */,
  {32'hbd566040, 32'hbec15720} /* (16, 17, 11) {real, imag} */,
  {32'h3e67bea0, 32'hbfef313a} /* (16, 17, 10) {real, imag} */,
  {32'h3e847028, 32'hbc56eb00} /* (16, 17, 9) {real, imag} */,
  {32'h3faa69e4, 32'h3fdf7c46} /* (16, 17, 8) {real, imag} */,
  {32'h3f837670, 32'h3fe3e7c4} /* (16, 17, 7) {real, imag} */,
  {32'h3ebf7ac2, 32'h3eba144c} /* (16, 17, 6) {real, imag} */,
  {32'hbf2e1e08, 32'h3ccd1da0} /* (16, 17, 5) {real, imag} */,
  {32'h3f54c74c, 32'hbdc97c88} /* (16, 17, 4) {real, imag} */,
  {32'h3fc6436c, 32'hbebf809e} /* (16, 17, 3) {real, imag} */,
  {32'hbeb96188, 32'h3ea76bc4} /* (16, 17, 2) {real, imag} */,
  {32'hbf588fda, 32'h3e68a6c0} /* (16, 17, 1) {real, imag} */,
  {32'hbf95b52c, 32'h3de81e34} /* (16, 17, 0) {real, imag} */,
  {32'hbf86b9f8, 32'h00000000} /* (16, 16, 31) {real, imag} */,
  {32'hbfa10ee8, 32'h00000000} /* (16, 16, 30) {real, imag} */,
  {32'h3d8f8968, 32'h00000000} /* (16, 16, 29) {real, imag} */,
  {32'h3f526bdc, 32'h00000000} /* (16, 16, 28) {real, imag} */,
  {32'h40039b9a, 32'h00000000} /* (16, 16, 27) {real, imag} */,
  {32'h40006dfd, 32'h00000000} /* (16, 16, 26) {real, imag} */,
  {32'h3ff45cc2, 32'h00000000} /* (16, 16, 25) {real, imag} */,
  {32'h3f1fc8a8, 32'h00000000} /* (16, 16, 24) {real, imag} */,
  {32'hbca04100, 32'h00000000} /* (16, 16, 23) {real, imag} */,
  {32'hbfd967fa, 32'h00000000} /* (16, 16, 22) {real, imag} */,
  {32'hbfded164, 32'h00000000} /* (16, 16, 21) {real, imag} */,
  {32'hbf400d21, 32'h00000000} /* (16, 16, 20) {real, imag} */,
  {32'h3ef8764c, 32'h00000000} /* (16, 16, 19) {real, imag} */,
  {32'h3ffcd282, 32'h00000000} /* (16, 16, 18) {real, imag} */,
  {32'h40192da6, 32'h00000000} /* (16, 16, 17) {real, imag} */,
  {32'h3fc7b1b3, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h402a2788, 32'h00000000} /* (16, 16, 15) {real, imag} */,
  {32'h3ef37380, 32'h00000000} /* (16, 16, 14) {real, imag} */,
  {32'h3c219000, 32'h00000000} /* (16, 16, 13) {real, imag} */,
  {32'hbf8f3295, 32'h00000000} /* (16, 16, 12) {real, imag} */,
  {32'hbf67af29, 32'h00000000} /* (16, 16, 11) {real, imag} */,
  {32'hbe4fa400, 32'h00000000} /* (16, 16, 10) {real, imag} */,
  {32'hbef423e0, 32'h00000000} /* (16, 16, 9) {real, imag} */,
  {32'hbeb40d70, 32'h00000000} /* (16, 16, 8) {real, imag} */,
  {32'hbf3a3fd4, 32'h00000000} /* (16, 16, 7) {real, imag} */,
  {32'h3e95f8e4, 32'h00000000} /* (16, 16, 6) {real, imag} */,
  {32'h3fad4bf6, 32'h00000000} /* (16, 16, 5) {real, imag} */,
  {32'h3eb6668e, 32'h00000000} /* (16, 16, 4) {real, imag} */,
  {32'hbbd85400, 32'h00000000} /* (16, 16, 3) {real, imag} */,
  {32'h3c8d5180, 32'h00000000} /* (16, 16, 2) {real, imag} */,
  {32'hbe6331a0, 32'h00000000} /* (16, 16, 1) {real, imag} */,
  {32'hbe5bf740, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'hbf7b6d18, 32'h3d19c6c0} /* (16, 15, 31) {real, imag} */,
  {32'hbfa047e1, 32'hbf8062d6} /* (16, 15, 30) {real, imag} */,
  {32'hbfd71f07, 32'hbf86d23d} /* (16, 15, 29) {real, imag} */,
  {32'hbfba16ce, 32'hbed3b0a4} /* (16, 15, 28) {real, imag} */,
  {32'hbeb8f910, 32'h3e32dc06} /* (16, 15, 27) {real, imag} */,
  {32'hbe61f350, 32'hbef46044} /* (16, 15, 26) {real, imag} */,
  {32'hbf0ae676, 32'h3f5867ec} /* (16, 15, 25) {real, imag} */,
  {32'hbf1a5d64, 32'h3f8352a8} /* (16, 15, 24) {real, imag} */,
  {32'hbfa1bdbc, 32'h3f080b36} /* (16, 15, 23) {real, imag} */,
  {32'hbf8d1281, 32'h3dbf3700} /* (16, 15, 22) {real, imag} */,
  {32'hbf327e90, 32'hbf851b97} /* (16, 15, 21) {real, imag} */,
  {32'hbee0a5b6, 32'hbecb016c} /* (16, 15, 20) {real, imag} */,
  {32'hbf29acaf, 32'hbe7bef6b} /* (16, 15, 19) {real, imag} */,
  {32'h3db2198c, 32'h3ebdb8fc} /* (16, 15, 18) {real, imag} */,
  {32'hbf901198, 32'h3f136fcd} /* (16, 15, 17) {real, imag} */,
  {32'hbfce6f45, 32'hbe11bf40} /* (16, 15, 16) {real, imag} */,
  {32'hbfa7e09c, 32'hbe9457b4} /* (16, 15, 15) {real, imag} */,
  {32'hbfff4ebc, 32'hbf8b2e0b} /* (16, 15, 14) {real, imag} */,
  {32'hbf5ea558, 32'hbf8d32dd} /* (16, 15, 13) {real, imag} */,
  {32'h3f3a1fd4, 32'hbf5d7cc5} /* (16, 15, 12) {real, imag} */,
  {32'hbd566040, 32'h3ec15720} /* (16, 15, 11) {real, imag} */,
  {32'h3e67bea0, 32'h3fef313a} /* (16, 15, 10) {real, imag} */,
  {32'h3e847028, 32'h3c56eb00} /* (16, 15, 9) {real, imag} */,
  {32'h3faa69e4, 32'hbfdf7c46} /* (16, 15, 8) {real, imag} */,
  {32'h3f837670, 32'hbfe3e7c4} /* (16, 15, 7) {real, imag} */,
  {32'h3ebf7ac2, 32'hbeba144c} /* (16, 15, 6) {real, imag} */,
  {32'hbf2e1e08, 32'hbccd1da0} /* (16, 15, 5) {real, imag} */,
  {32'h3f54c74c, 32'h3dc97c88} /* (16, 15, 4) {real, imag} */,
  {32'h3fc6436c, 32'h3ebf809e} /* (16, 15, 3) {real, imag} */,
  {32'hbeb96188, 32'hbea76bc4} /* (16, 15, 2) {real, imag} */,
  {32'hbf588fda, 32'hbe68a6c0} /* (16, 15, 1) {real, imag} */,
  {32'hbf95b52c, 32'hbde81e34} /* (16, 15, 0) {real, imag} */,
  {32'h3f650bf9, 32'h3fb223ec} /* (16, 14, 31) {real, imag} */,
  {32'h4011d02e, 32'h4031e266} /* (16, 14, 30) {real, imag} */,
  {32'h3f48a194, 32'h3f41fd74} /* (16, 14, 29) {real, imag} */,
  {32'h3f2f4f1a, 32'hbdd91c40} /* (16, 14, 28) {real, imag} */,
  {32'h3f1ef124, 32'h3d601780} /* (16, 14, 27) {real, imag} */,
  {32'h3e9cbd40, 32'h3f339044} /* (16, 14, 26) {real, imag} */,
  {32'h3faf35e8, 32'h3de97560} /* (16, 14, 25) {real, imag} */,
  {32'h3f445d4d, 32'hbed2885d} /* (16, 14, 24) {real, imag} */,
  {32'h3fe04474, 32'h3fba71fe} /* (16, 14, 23) {real, imag} */,
  {32'h400b9dae, 32'h3f8128f2} /* (16, 14, 22) {real, imag} */,
  {32'h3ff27a3a, 32'h3f511de8} /* (16, 14, 21) {real, imag} */,
  {32'h3f207866, 32'hbf317780} /* (16, 14, 20) {real, imag} */,
  {32'h3f63a6c0, 32'hbf9cc4e2} /* (16, 14, 19) {real, imag} */,
  {32'h3dc15928, 32'hbfdbf4e8} /* (16, 14, 18) {real, imag} */,
  {32'hbee97c10, 32'hbf65f528} /* (16, 14, 17) {real, imag} */,
  {32'hbfc7bb02, 32'hbe934f18} /* (16, 14, 16) {real, imag} */,
  {32'h3db549f0, 32'h3fad459c} /* (16, 14, 15) {real, imag} */,
  {32'h4009ae30, 32'h3ece17f4} /* (16, 14, 14) {real, imag} */,
  {32'h3ec2a289, 32'h3e81225e} /* (16, 14, 13) {real, imag} */,
  {32'hbf8c15ac, 32'h3f8fc132} /* (16, 14, 12) {real, imag} */,
  {32'h3f005f5f, 32'h3f9be75f} /* (16, 14, 11) {real, imag} */,
  {32'h3efccd70, 32'h3e8613a0} /* (16, 14, 10) {real, imag} */,
  {32'hbda7e580, 32'hbf34129e} /* (16, 14, 9) {real, imag} */,
  {32'h3ea15dd8, 32'hbf58c0c0} /* (16, 14, 8) {real, imag} */,
  {32'hbf0fcd56, 32'hbf156c34} /* (16, 14, 7) {real, imag} */,
  {32'h3d51cac0, 32'hbf7c5f08} /* (16, 14, 6) {real, imag} */,
  {32'h3e02d6ec, 32'hbee1d9e0} /* (16, 14, 5) {real, imag} */,
  {32'hbf9709df, 32'h3eacee95} /* (16, 14, 4) {real, imag} */,
  {32'hbf768f70, 32'h3fa8eb45} /* (16, 14, 3) {real, imag} */,
  {32'hbe948c90, 32'h3db861e0} /* (16, 14, 2) {real, imag} */,
  {32'hbefa5528, 32'hbf77c071} /* (16, 14, 1) {real, imag} */,
  {32'hbea50724, 32'hbf0868ac} /* (16, 14, 0) {real, imag} */,
  {32'h3ef48dac, 32'hbeb3005b} /* (16, 13, 31) {real, imag} */,
  {32'h3f68840c, 32'hbfcf30fc} /* (16, 13, 30) {real, imag} */,
  {32'h402fa71e, 32'hbe86eb76} /* (16, 13, 29) {real, imag} */,
  {32'h4017313a, 32'h3f9c2d03} /* (16, 13, 28) {real, imag} */,
  {32'hbf1d61e4, 32'h3f6d80c8} /* (16, 13, 27) {real, imag} */,
  {32'hbfb05da0, 32'hbfaa078c} /* (16, 13, 26) {real, imag} */,
  {32'hc0195b98, 32'hbfc5ce71} /* (16, 13, 25) {real, imag} */,
  {32'h3f8e1db4, 32'hbfc239d2} /* (16, 13, 24) {real, imag} */,
  {32'h3fac41e4, 32'h3f532eac} /* (16, 13, 23) {real, imag} */,
  {32'h3f44c585, 32'h3fde39b9} /* (16, 13, 22) {real, imag} */,
  {32'h3fed678c, 32'hbfa59b74} /* (16, 13, 21) {real, imag} */,
  {32'h407476e6, 32'hbfe7cf54} /* (16, 13, 20) {real, imag} */,
  {32'h3fdd7fe6, 32'hbfbc02b9} /* (16, 13, 19) {real, imag} */,
  {32'h3d7ab370, 32'hbddd8c40} /* (16, 13, 18) {real, imag} */,
  {32'hbf109228, 32'h3eeb6120} /* (16, 13, 17) {real, imag} */,
  {32'hbe83aca8, 32'hbe39f4d0} /* (16, 13, 16) {real, imag} */,
  {32'hbee46154, 32'hbf51beec} /* (16, 13, 15) {real, imag} */,
  {32'h3f182f70, 32'h3f476850} /* (16, 13, 14) {real, imag} */,
  {32'hbf1d150c, 32'h3f9fe252} /* (16, 13, 13) {real, imag} */,
  {32'hbf378dd4, 32'h3e927684} /* (16, 13, 12) {real, imag} */,
  {32'hbfa6881b, 32'hbf102f34} /* (16, 13, 11) {real, imag} */,
  {32'hbfdbb7fd, 32'h3ee1a088} /* (16, 13, 10) {real, imag} */,
  {32'hc00094d6, 32'h3fb2db52} /* (16, 13, 9) {real, imag} */,
  {32'hc09188ed, 32'h4087f3ef} /* (16, 13, 8) {real, imag} */,
  {32'hc0226b91, 32'h401a3f14} /* (16, 13, 7) {real, imag} */,
  {32'hbfc6ee66, 32'hbf2b6b70} /* (16, 13, 6) {real, imag} */,
  {32'hbebc4058, 32'h3f43b019} /* (16, 13, 5) {real, imag} */,
  {32'h3eb4c7e6, 32'h3f54ae48} /* (16, 13, 4) {real, imag} */,
  {32'hbf2727dc, 32'hbf13ca41} /* (16, 13, 3) {real, imag} */,
  {32'h3f800184, 32'h3ed51dd0} /* (16, 13, 2) {real, imag} */,
  {32'h3fc711b8, 32'h3f380112} /* (16, 13, 1) {real, imag} */,
  {32'h3f60456a, 32'h3e163949} /* (16, 13, 0) {real, imag} */,
  {32'h3fcdc6f6, 32'hbe8e04a8} /* (16, 12, 31) {real, imag} */,
  {32'h3fe40ec6, 32'hc024b9c0} /* (16, 12, 30) {real, imag} */,
  {32'h3ea94343, 32'hbdadbde0} /* (16, 12, 29) {real, imag} */,
  {32'hbf06afcb, 32'h3fe312b4} /* (16, 12, 28) {real, imag} */,
  {32'hbee38ad4, 32'hbf9acab5} /* (16, 12, 27) {real, imag} */,
  {32'hbf99213e, 32'hc038669d} /* (16, 12, 26) {real, imag} */,
  {32'hbf928360, 32'h3f3a86d4} /* (16, 12, 25) {real, imag} */,
  {32'h3fc69a46, 32'h3ee35120} /* (16, 12, 24) {real, imag} */,
  {32'h404d548d, 32'h3ee7c7e0} /* (16, 12, 23) {real, imag} */,
  {32'h3fc9001b, 32'hbf9f3528} /* (16, 12, 22) {real, imag} */,
  {32'hbece7dac, 32'hc03c7b4b} /* (16, 12, 21) {real, imag} */,
  {32'h3f02ad95, 32'hbd43aa80} /* (16, 12, 20) {real, imag} */,
  {32'h400c7d72, 32'hbe122740} /* (16, 12, 19) {real, imag} */,
  {32'h3f6671a3, 32'hbf1425f1} /* (16, 12, 18) {real, imag} */,
  {32'h3f6413c4, 32'h3e04a3e0} /* (16, 12, 17) {real, imag} */,
  {32'h40105858, 32'h3f1a4f73} /* (16, 12, 16) {real, imag} */,
  {32'h3fb541e4, 32'h40585947} /* (16, 12, 15) {real, imag} */,
  {32'h3eee39d8, 32'h4035ec7c} /* (16, 12, 14) {real, imag} */,
  {32'h3f8c65ad, 32'hbf160694} /* (16, 12, 13) {real, imag} */,
  {32'h3eb9bc2e, 32'hbf28b8cb} /* (16, 12, 12) {real, imag} */,
  {32'h3df0b278, 32'hbfe3af72} /* (16, 12, 11) {real, imag} */,
  {32'h40514b9b, 32'hc009f2f0} /* (16, 12, 10) {real, imag} */,
  {32'h3fdd55d4, 32'hbfb3213c} /* (16, 12, 9) {real, imag} */,
  {32'h401de698, 32'h3ec4e1a8} /* (16, 12, 8) {real, imag} */,
  {32'h3ffa8e14, 32'hbf1b2b20} /* (16, 12, 7) {real, imag} */,
  {32'hbc093800, 32'hbf41b4a0} /* (16, 12, 6) {real, imag} */,
  {32'h3fa76e04, 32'h3edf7308} /* (16, 12, 5) {real, imag} */,
  {32'hbf3d5c1d, 32'hbf7042f5} /* (16, 12, 4) {real, imag} */,
  {32'h3f57869c, 32'hc03a2992} /* (16, 12, 3) {real, imag} */,
  {32'hbf6cd8a6, 32'hbfe1c28b} /* (16, 12, 2) {real, imag} */,
  {32'hbfc18218, 32'h3f92e150} /* (16, 12, 1) {real, imag} */,
  {32'hbe9d5673, 32'h401c6506} /* (16, 12, 0) {real, imag} */,
  {32'h3f9652be, 32'h3f92aecb} /* (16, 11, 31) {real, imag} */,
  {32'h3ea63698, 32'h3f168d74} /* (16, 11, 30) {real, imag} */,
  {32'h3f4b16d1, 32'hbfdf4832} /* (16, 11, 29) {real, imag} */,
  {32'h3ffa6b89, 32'hbfb2dff9} /* (16, 11, 28) {real, imag} */,
  {32'h3fa01db0, 32'hc03e6aaa} /* (16, 11, 27) {real, imag} */,
  {32'hbf53058e, 32'hc035aa44} /* (16, 11, 26) {real, imag} */,
  {32'hbf68da2a, 32'hbd8554f0} /* (16, 11, 25) {real, imag} */,
  {32'hbff2d54b, 32'h3fbc4fa5} /* (16, 11, 24) {real, imag} */,
  {32'hbfe1f34c, 32'h3c972f80} /* (16, 11, 23) {real, imag} */,
  {32'hbec56108, 32'hbe3d7118} /* (16, 11, 22) {real, imag} */,
  {32'h3f68d772, 32'hbf83d970} /* (16, 11, 21) {real, imag} */,
  {32'h3ee85608, 32'hbfbb837e} /* (16, 11, 20) {real, imag} */,
  {32'h3ec3fee6, 32'h3ef9c604} /* (16, 11, 19) {real, imag} */,
  {32'h40204ec3, 32'hbf8148a8} /* (16, 11, 18) {real, imag} */,
  {32'h3fd4acdc, 32'hbf150c26} /* (16, 11, 17) {real, imag} */,
  {32'h3fa029ea, 32'h3d828a70} /* (16, 11, 16) {real, imag} */,
  {32'h3f59e720, 32'hbf61e884} /* (16, 11, 15) {real, imag} */,
  {32'h3ea470e0, 32'hbf2cc7cc} /* (16, 11, 14) {real, imag} */,
  {32'hbe0cea68, 32'hc0039c42} /* (16, 11, 13) {real, imag} */,
  {32'hc01ce3d4, 32'hc00da9a6} /* (16, 11, 12) {real, imag} */,
  {32'hc04b2b8c, 32'hbfb8138c} /* (16, 11, 11) {real, imag} */,
  {32'hbfc05e68, 32'hbe0677f8} /* (16, 11, 10) {real, imag} */,
  {32'h400ebe64, 32'hbf0f5360} /* (16, 11, 9) {real, imag} */,
  {32'hbe8eb3c0, 32'hbfc420bf} /* (16, 11, 8) {real, imag} */,
  {32'hbe3fd1ba, 32'h3eef1daa} /* (16, 11, 7) {real, imag} */,
  {32'h3f8b619a, 32'hbfbac5cf} /* (16, 11, 6) {real, imag} */,
  {32'h3fcd0e20, 32'hbf93ce66} /* (16, 11, 5) {real, imag} */,
  {32'hbe6fabde, 32'h3df3eae0} /* (16, 11, 4) {real, imag} */,
  {32'hc0333adb, 32'h401acfb6} /* (16, 11, 3) {real, imag} */,
  {32'hc008a4ba, 32'h3f9776cd} /* (16, 11, 2) {real, imag} */,
  {32'hc005186c, 32'hbeb3c86c} /* (16, 11, 1) {real, imag} */,
  {32'hbe8a376c, 32'h3f9f4d7f} /* (16, 11, 0) {real, imag} */,
  {32'hbf196fc8, 32'hbf7989a8} /* (16, 10, 31) {real, imag} */,
  {32'h3ebc7038, 32'hbe8c1a38} /* (16, 10, 30) {real, imag} */,
  {32'h3f3ecf12, 32'hbfbe38f9} /* (16, 10, 29) {real, imag} */,
  {32'hbf17bc44, 32'h3fa9fa40} /* (16, 10, 28) {real, imag} */,
  {32'h40086062, 32'h3f1d9db4} /* (16, 10, 27) {real, imag} */,
  {32'h40803b63, 32'hbfb2f19a} /* (16, 10, 26) {real, imag} */,
  {32'h404df57e, 32'h3fb3ad38} /* (16, 10, 25) {real, imag} */,
  {32'hbf25a602, 32'hbf47a836} /* (16, 10, 24) {real, imag} */,
  {32'hc02cb023, 32'hc035ca04} /* (16, 10, 23) {real, imag} */,
  {32'hc0119a54, 32'hbf1cc0b0} /* (16, 10, 22) {real, imag} */,
  {32'hbe5a1d38, 32'h3f36fd74} /* (16, 10, 21) {real, imag} */,
  {32'h3febfe31, 32'h3eda3715} /* (16, 10, 20) {real, imag} */,
  {32'h3fca9065, 32'hbd0efd80} /* (16, 10, 19) {real, imag} */,
  {32'hbe8da374, 32'h40057af7} /* (16, 10, 18) {real, imag} */,
  {32'h3f28a495, 32'hbf5e3ad0} /* (16, 10, 17) {real, imag} */,
  {32'h3fd8d98e, 32'hc01f8c42} /* (16, 10, 16) {real, imag} */,
  {32'h4045e130, 32'hc025df3b} /* (16, 10, 15) {real, imag} */,
  {32'h40651dad, 32'hbfba5656} /* (16, 10, 14) {real, imag} */,
  {32'h40374826, 32'hbe4735b0} /* (16, 10, 13) {real, imag} */,
  {32'h4027222c, 32'hbe592858} /* (16, 10, 12) {real, imag} */,
  {32'h400c1772, 32'hbf8c4ec5} /* (16, 10, 11) {real, imag} */,
  {32'h3fe5e43c, 32'h3ff92848} /* (16, 10, 10) {real, imag} */,
  {32'h4018aa96, 32'hc029d0b2} /* (16, 10, 9) {real, imag} */,
  {32'h400feb65, 32'hc0885258} /* (16, 10, 8) {real, imag} */,
  {32'hbfc3de92, 32'hbcf6ebc0} /* (16, 10, 7) {real, imag} */,
  {32'h3f9022ed, 32'hbea873e8} /* (16, 10, 6) {real, imag} */,
  {32'h4037b196, 32'hbf283d40} /* (16, 10, 5) {real, imag} */,
  {32'h402aa83e, 32'hbfa376c0} /* (16, 10, 4) {real, imag} */,
  {32'h40379ec8, 32'hc00caab4} /* (16, 10, 3) {real, imag} */,
  {32'hbf3ad014, 32'h3df838f0} /* (16, 10, 2) {real, imag} */,
  {32'hc08dca55, 32'h3e56c4d0} /* (16, 10, 1) {real, imag} */,
  {32'hc018886f, 32'hbe2a7270} /* (16, 10, 0) {real, imag} */,
  {32'h3fc309ae, 32'h3fc101a2} /* (16, 9, 31) {real, imag} */,
  {32'h3fd13fc7, 32'h3facc426} /* (16, 9, 30) {real, imag} */,
  {32'hc03f206e, 32'h40448446} /* (16, 9, 29) {real, imag} */,
  {32'hbfbda444, 32'h3fb52146} /* (16, 9, 28) {real, imag} */,
  {32'h40565b53, 32'hbe587fba} /* (16, 9, 27) {real, imag} */,
  {32'h3fc2592a, 32'hbe48512e} /* (16, 9, 26) {real, imag} */,
  {32'hbf985f69, 32'h3ef19a2a} /* (16, 9, 25) {real, imag} */,
  {32'hc01c3235, 32'h3fdc9ca9} /* (16, 9, 24) {real, imag} */,
  {32'hbf2176a5, 32'h407786d0} /* (16, 9, 23) {real, imag} */,
  {32'h3d8d0000, 32'h4027ae72} /* (16, 9, 22) {real, imag} */,
  {32'hbf56fc6e, 32'h3f23f790} /* (16, 9, 21) {real, imag} */,
  {32'hbfaa4076, 32'hbea9251c} /* (16, 9, 20) {real, imag} */,
  {32'h40343190, 32'h3ef250dc} /* (16, 9, 19) {real, imag} */,
  {32'hbf00e634, 32'h3ff53efa} /* (16, 9, 18) {real, imag} */,
  {32'hc03250c2, 32'h3dc874cc} /* (16, 9, 17) {real, imag} */,
  {32'hbfdcfa64, 32'h3f4e4928} /* (16, 9, 16) {real, imag} */,
  {32'hbe951d2e, 32'h3ec7526a} /* (16, 9, 15) {real, imag} */,
  {32'h3fe557a8, 32'hc04c88a3} /* (16, 9, 14) {real, imag} */,
  {32'hbf00f746, 32'h3ed77be0} /* (16, 9, 13) {real, imag} */,
  {32'hbfda1b77, 32'hbf5355f8} /* (16, 9, 12) {real, imag} */,
  {32'h4065b601, 32'h3e785380} /* (16, 9, 11) {real, imag} */,
  {32'h401b2054, 32'hc0766d4e} /* (16, 9, 10) {real, imag} */,
  {32'hbe31d650, 32'hc0050dd7} /* (16, 9, 9) {real, imag} */,
  {32'hbcb04800, 32'hc06f2223} /* (16, 9, 8) {real, imag} */,
  {32'h3f68530f, 32'hc0a9195d} /* (16, 9, 7) {real, imag} */,
  {32'h3fe3e0fc, 32'hbf172aa1} /* (16, 9, 6) {real, imag} */,
  {32'hbd40ecc0, 32'hbef646e4} /* (16, 9, 5) {real, imag} */,
  {32'h3f47d018, 32'h405b6a3e} /* (16, 9, 4) {real, imag} */,
  {32'hbfaf31c2, 32'h409a4078} /* (16, 9, 3) {real, imag} */,
  {32'hbfc91dd1, 32'h4088b52c} /* (16, 9, 2) {real, imag} */,
  {32'h3faf2af6, 32'h4089328f} /* (16, 9, 1) {real, imag} */,
  {32'hbfc775fc, 32'h40962d39} /* (16, 9, 0) {real, imag} */,
  {32'hbf92c480, 32'h3f33c2f6} /* (16, 8, 31) {real, imag} */,
  {32'hbfc42048, 32'h3f960228} /* (16, 8, 30) {real, imag} */,
  {32'h3ee21602, 32'h40ade1ee} /* (16, 8, 29) {real, imag} */,
  {32'h409fe4d5, 32'h40e726da} /* (16, 8, 28) {real, imag} */,
  {32'h40dbcc38, 32'h40909820} /* (16, 8, 27) {real, imag} */,
  {32'h3fbeea7f, 32'hbefd8194} /* (16, 8, 26) {real, imag} */,
  {32'hbf5a94b4, 32'hbfedf14b} /* (16, 8, 25) {real, imag} */,
  {32'hbf998346, 32'h3f090778} /* (16, 8, 24) {real, imag} */,
  {32'hc07651ed, 32'h4015218b} /* (16, 8, 23) {real, imag} */,
  {32'hc08c6a44, 32'h4073a21a} /* (16, 8, 22) {real, imag} */,
  {32'hbf94d570, 32'h3e6b9570} /* (16, 8, 21) {real, imag} */,
  {32'hc03b9c16, 32'hbeae266e} /* (16, 8, 20) {real, imag} */,
  {32'hc054e0f4, 32'h3fdde60c} /* (16, 8, 19) {real, imag} */,
  {32'hbf442028, 32'hc049001b} /* (16, 8, 18) {real, imag} */,
  {32'h3f632bd3, 32'hc09ea006} /* (16, 8, 17) {real, imag} */,
  {32'hbf1ceb9a, 32'hc0b12c28} /* (16, 8, 16) {real, imag} */,
  {32'hbf3fc0de, 32'hc027eacd} /* (16, 8, 15) {real, imag} */,
  {32'h3f5e8268, 32'hbf592ad4} /* (16, 8, 14) {real, imag} */,
  {32'h40576de5, 32'hbe334724} /* (16, 8, 13) {real, imag} */,
  {32'hc02e88d0, 32'hbf81cc3d} /* (16, 8, 12) {real, imag} */,
  {32'hbdb12568, 32'hc011ea9e} /* (16, 8, 11) {real, imag} */,
  {32'hbe9842d0, 32'hbfa9c6a8} /* (16, 8, 10) {real, imag} */,
  {32'h3e99b858, 32'hc064daed} /* (16, 8, 9) {real, imag} */,
  {32'h3f8f74d6, 32'hbfbc385a} /* (16, 8, 8) {real, imag} */,
  {32'h3fff461a, 32'h3fa6ae4f} /* (16, 8, 7) {real, imag} */,
  {32'h3fe62333, 32'hbf400fef} /* (16, 8, 6) {real, imag} */,
  {32'hbe567b44, 32'hc04e3da6} /* (16, 8, 5) {real, imag} */,
  {32'hc0337198, 32'h3f62ca9d} /* (16, 8, 4) {real, imag} */,
  {32'hbfddb6a8, 32'h405b6d60} /* (16, 8, 3) {real, imag} */,
  {32'h3f26b76c, 32'h40421eec} /* (16, 8, 2) {real, imag} */,
  {32'hbfde41f5, 32'h3fa93050} /* (16, 8, 1) {real, imag} */,
  {32'hc00f17f6, 32'h3f8828be} /* (16, 8, 0) {real, imag} */,
  {32'h3ec5f2da, 32'h407a2e2b} /* (16, 7, 31) {real, imag} */,
  {32'h400e7ab6, 32'h404e3105} /* (16, 7, 30) {real, imag} */,
  {32'h407ce3ae, 32'hc0077340} /* (16, 7, 29) {real, imag} */,
  {32'h3e184290, 32'hc068b145} /* (16, 7, 28) {real, imag} */,
  {32'hbf7921c4, 32'hbf6920b2} /* (16, 7, 27) {real, imag} */,
  {32'h3fc384fc, 32'hbdbb5a24} /* (16, 7, 26) {real, imag} */,
  {32'h3fcc3793, 32'hbe9e232e} /* (16, 7, 25) {real, imag} */,
  {32'h3d25d0c0, 32'h3fb1ef0d} /* (16, 7, 24) {real, imag} */,
  {32'hbf35cdb1, 32'h3ed62f0c} /* (16, 7, 23) {real, imag} */,
  {32'hbf1cd3ec, 32'hbf04bb2a} /* (16, 7, 22) {real, imag} */,
  {32'h4081420d, 32'h3d8f9e40} /* (16, 7, 21) {real, imag} */,
  {32'h40108827, 32'h4005f41a} /* (16, 7, 20) {real, imag} */,
  {32'hbeeab028, 32'h3f4742e8} /* (16, 7, 19) {real, imag} */,
  {32'h3e5332a0, 32'h3f35cdbf} /* (16, 7, 18) {real, imag} */,
  {32'hbf9385f0, 32'h3f360c12} /* (16, 7, 17) {real, imag} */,
  {32'hbf2af650, 32'h3e00767e} /* (16, 7, 16) {real, imag} */,
  {32'h3f2b9e8a, 32'hbf9342c8} /* (16, 7, 15) {real, imag} */,
  {32'hc0138f22, 32'h40902cd9} /* (16, 7, 14) {real, imag} */,
  {32'hc0656214, 32'h408a618d} /* (16, 7, 13) {real, imag} */,
  {32'h3f86430b, 32'h406b1964} /* (16, 7, 12) {real, imag} */,
  {32'h40188ff9, 32'h401082cd} /* (16, 7, 11) {real, imag} */,
  {32'hbff432b4, 32'h3fbc842c} /* (16, 7, 10) {real, imag} */,
  {32'hbffee8f8, 32'h3fc9a566} /* (16, 7, 9) {real, imag} */,
  {32'hbfc271c0, 32'h3faf36e2} /* (16, 7, 8) {real, imag} */,
  {32'h3ee8b676, 32'h3e98b3a0} /* (16, 7, 7) {real, imag} */,
  {32'h3fec8c8a, 32'h3f02cf7b} /* (16, 7, 6) {real, imag} */,
  {32'h406d296c, 32'h3ff03827} /* (16, 7, 5) {real, imag} */,
  {32'h400148e8, 32'hbfa54a2c} /* (16, 7, 4) {real, imag} */,
  {32'hbfa28b3c, 32'hc0155d31} /* (16, 7, 3) {real, imag} */,
  {32'hbdd2bef0, 32'h3e9d0c20} /* (16, 7, 2) {real, imag} */,
  {32'hc0107bd4, 32'h4013732c} /* (16, 7, 1) {real, imag} */,
  {32'hc06280f6, 32'h4046a322} /* (16, 7, 0) {real, imag} */,
  {32'hc0764708, 32'hc0304cf4} /* (16, 6, 31) {real, imag} */,
  {32'hc0537c6e, 32'hc092d34a} /* (16, 6, 30) {real, imag} */,
  {32'hbffd0743, 32'hc083f259} /* (16, 6, 29) {real, imag} */,
  {32'hc08a6000, 32'hbf5d950f} /* (16, 6, 28) {real, imag} */,
  {32'hbe197b10, 32'hbf5a5ee0} /* (16, 6, 27) {real, imag} */,
  {32'hc01234fe, 32'hbe79fec4} /* (16, 6, 26) {real, imag} */,
  {32'hbf8ee2bd, 32'hbfa1d60a} /* (16, 6, 25) {real, imag} */,
  {32'hbeb0b09e, 32'hbeb730dc} /* (16, 6, 24) {real, imag} */,
  {32'hc01c7865, 32'hc049f57c} /* (16, 6, 23) {real, imag} */,
  {32'hbeca20cc, 32'h3dd6e894} /* (16, 6, 22) {real, imag} */,
  {32'h4047148e, 32'h3fc6c242} /* (16, 6, 21) {real, imag} */,
  {32'h3fa548ed, 32'h3e8aa6b5} /* (16, 6, 20) {real, imag} */,
  {32'h3f5f0f4e, 32'h40482e3a} /* (16, 6, 19) {real, imag} */,
  {32'h3f6a3fc6, 32'h3f813d22} /* (16, 6, 18) {real, imag} */,
  {32'h40169291, 32'hc02e8e5a} /* (16, 6, 17) {real, imag} */,
  {32'h402c7097, 32'hbf1a67a0} /* (16, 6, 16) {real, imag} */,
  {32'h3fde0fa8, 32'hbf7df728} /* (16, 6, 15) {real, imag} */,
  {32'hbf5038bc, 32'h3e2e79a4} /* (16, 6, 14) {real, imag} */,
  {32'h3fe10e25, 32'h404249c7} /* (16, 6, 13) {real, imag} */,
  {32'h40a5c7dd, 32'h404b4544} /* (16, 6, 12) {real, imag} */,
  {32'hbd2aade0, 32'h3f9152eb} /* (16, 6, 11) {real, imag} */,
  {32'hc08ccbb4, 32'hbd485c00} /* (16, 6, 10) {real, imag} */,
  {32'h3e906574, 32'h3f8c9cc9} /* (16, 6, 9) {real, imag} */,
  {32'h4096a704, 32'h3eb0c6b8} /* (16, 6, 8) {real, imag} */,
  {32'h3f94b846, 32'hc0255646} /* (16, 6, 7) {real, imag} */,
  {32'h3f8ac2bf, 32'hc0d1a568} /* (16, 6, 6) {real, imag} */,
  {32'hbdde4fc0, 32'hc0b9b7d8} /* (16, 6, 5) {real, imag} */,
  {32'h3fdbc58b, 32'hc0e50826} /* (16, 6, 4) {real, imag} */,
  {32'h4018fc20, 32'hc09db47b} /* (16, 6, 3) {real, imag} */,
  {32'h3eb78688, 32'h4016ad56} /* (16, 6, 2) {real, imag} */,
  {32'hc01b5b28, 32'h408400a2} /* (16, 6, 1) {real, imag} */,
  {32'hbf841638, 32'hc00ab261} /* (16, 6, 0) {real, imag} */,
  {32'hbdbdb638, 32'h3fe4f025} /* (16, 5, 31) {real, imag} */,
  {32'hc080867e, 32'hbda8eae0} /* (16, 5, 30) {real, imag} */,
  {32'hbf1a6a71, 32'hc075a997} /* (16, 5, 29) {real, imag} */,
  {32'hbfcc907b, 32'hbefaa5ac} /* (16, 5, 28) {real, imag} */,
  {32'hc0548b48, 32'hbf937ca5} /* (16, 5, 27) {real, imag} */,
  {32'hc0169dde, 32'hbfa67515} /* (16, 5, 26) {real, imag} */,
  {32'h3def4574, 32'hc04bd5c8} /* (16, 5, 25) {real, imag} */,
  {32'h3fb62f4d, 32'hc08260fa} /* (16, 5, 24) {real, imag} */,
  {32'h4011b910, 32'hc084169a} /* (16, 5, 23) {real, imag} */,
  {32'hbe914cf8, 32'hbfdb1429} /* (16, 5, 22) {real, imag} */,
  {32'h3f79e72a, 32'h3ff1beb8} /* (16, 5, 21) {real, imag} */,
  {32'h40a79f12, 32'h3e484148} /* (16, 5, 20) {real, imag} */,
  {32'h4013a4c7, 32'h3feab243} /* (16, 5, 19) {real, imag} */,
  {32'h3f08cf3c, 32'h3e275c94} /* (16, 5, 18) {real, imag} */,
  {32'h4073cd62, 32'h3eb42ccc} /* (16, 5, 17) {real, imag} */,
  {32'hbfc35642, 32'hbf988d7f} /* (16, 5, 16) {real, imag} */,
  {32'hc0bc94ce, 32'hbf3b6eae} /* (16, 5, 15) {real, imag} */,
  {32'hc0aa656f, 32'h3fec82a2} /* (16, 5, 14) {real, imag} */,
  {32'hc06c3706, 32'h406bb2be} /* (16, 5, 13) {real, imag} */,
  {32'h3ff82019, 32'h40081454} /* (16, 5, 12) {real, imag} */,
  {32'h3f833cff, 32'h3d3827d0} /* (16, 5, 11) {real, imag} */,
  {32'h4011fa8b, 32'hc01bb63c} /* (16, 5, 10) {real, imag} */,
  {32'h409dbdfa, 32'hc021d7f2} /* (16, 5, 9) {real, imag} */,
  {32'h4008ec43, 32'hc096d14e} /* (16, 5, 8) {real, imag} */,
  {32'hbf664b76, 32'hbfbfc8f8} /* (16, 5, 7) {real, imag} */,
  {32'hbfbbcd96, 32'hbf907563} /* (16, 5, 6) {real, imag} */,
  {32'hc039ba70, 32'hc040b4d5} /* (16, 5, 5) {real, imag} */,
  {32'h3d88d5dc, 32'hc09026ba} /* (16, 5, 4) {real, imag} */,
  {32'h3eb299a8, 32'hc0aa799e} /* (16, 5, 3) {real, imag} */,
  {32'h3f2b92a2, 32'hc06b008a} /* (16, 5, 2) {real, imag} */,
  {32'hbfc3cd85, 32'h3fcd9527} /* (16, 5, 1) {real, imag} */,
  {32'hbee7d7cc, 32'h403e49ae} /* (16, 5, 0) {real, imag} */,
  {32'h3ebd9542, 32'hbe675bb0} /* (16, 4, 31) {real, imag} */,
  {32'hc071968d, 32'hc08503c1} /* (16, 4, 30) {real, imag} */,
  {32'h3eab1b79, 32'hc0c398ec} /* (16, 4, 29) {real, imag} */,
  {32'h3fafabae, 32'hc03ad8ee} /* (16, 4, 28) {real, imag} */,
  {32'h3fe5fb29, 32'hc030943c} /* (16, 4, 27) {real, imag} */,
  {32'h407725cf, 32'h40a4fa02} /* (16, 4, 26) {real, imag} */,
  {32'h4044afde, 32'h403c95b4} /* (16, 4, 25) {real, imag} */,
  {32'h4003f723, 32'hc0f99c4a} /* (16, 4, 24) {real, imag} */,
  {32'hc0a2afcc, 32'hc0f1d3d2} /* (16, 4, 23) {real, imag} */,
  {32'h3fbe3ab3, 32'hc00293fb} /* (16, 4, 22) {real, imag} */,
  {32'h4029a040, 32'h40018fe7} /* (16, 4, 21) {real, imag} */,
  {32'hbfdb7b5a, 32'h40ab2025} /* (16, 4, 20) {real, imag} */,
  {32'hbfcedff9, 32'h40c5d144} /* (16, 4, 19) {real, imag} */,
  {32'h3fe8b55a, 32'h3fdac988} /* (16, 4, 18) {real, imag} */,
  {32'hc06f3d83, 32'h40c63df3} /* (16, 4, 17) {real, imag} */,
  {32'hc0616208, 32'h3f94ca00} /* (16, 4, 16) {real, imag} */,
  {32'hc0ba8e53, 32'h3e41e9f0} /* (16, 4, 15) {real, imag} */,
  {32'hc0298567, 32'h40711b16} /* (16, 4, 14) {real, imag} */,
  {32'hbdf0cef0, 32'h40c4feb4} /* (16, 4, 13) {real, imag} */,
  {32'hbec87a56, 32'h3fcf2de4} /* (16, 4, 12) {real, imag} */,
  {32'hbf69bc7d, 32'hc023278f} /* (16, 4, 11) {real, imag} */,
  {32'h3fc35b6a, 32'hbf251aca} /* (16, 4, 10) {real, imag} */,
  {32'h3fe937c8, 32'hc017982e} /* (16, 4, 9) {real, imag} */,
  {32'hc076cc8c, 32'hc0e7a1aa} /* (16, 4, 8) {real, imag} */,
  {32'hc0131036, 32'hc0a35826} /* (16, 4, 7) {real, imag} */,
  {32'hc0add5a2, 32'hc0d30c84} /* (16, 4, 6) {real, imag} */,
  {32'hc0845f15, 32'hc081af1e} /* (16, 4, 5) {real, imag} */,
  {32'hbf7dbe6f, 32'h3d86ee28} /* (16, 4, 4) {real, imag} */,
  {32'h4064965d, 32'h40122670} /* (16, 4, 3) {real, imag} */,
  {32'hbf8e20a5, 32'hbf888797} /* (16, 4, 2) {real, imag} */,
  {32'hbf18b514, 32'hbe93be22} /* (16, 4, 1) {real, imag} */,
  {32'hbe31580a, 32'h3f57257d} /* (16, 4, 0) {real, imag} */,
  {32'hc069f49a, 32'h3d156bf8} /* (16, 3, 31) {real, imag} */,
  {32'hc09f7d2e, 32'h405173aa} /* (16, 3, 30) {real, imag} */,
  {32'hc1037962, 32'h400ba439} /* (16, 3, 29) {real, imag} */,
  {32'hc0c698ef, 32'hbfe72323} /* (16, 3, 28) {real, imag} */,
  {32'hbff34c8e, 32'hbfe32a7a} /* (16, 3, 27) {real, imag} */,
  {32'h4085fd8b, 32'hbdf161e0} /* (16, 3, 26) {real, imag} */,
  {32'h4089b052, 32'hc0206962} /* (16, 3, 25) {real, imag} */,
  {32'hbf5e976b, 32'h407a324d} /* (16, 3, 24) {real, imag} */,
  {32'h4031e506, 32'h4087d4b2} /* (16, 3, 23) {real, imag} */,
  {32'hbe14c7bc, 32'h3f2b06a6} /* (16, 3, 22) {real, imag} */,
  {32'hc0510e50, 32'h40a1b64d} /* (16, 3, 21) {real, imag} */,
  {32'hbf298510, 32'h3d921e68} /* (16, 3, 20) {real, imag} */,
  {32'h3ff5a25e, 32'hbfa92e93} /* (16, 3, 19) {real, imag} */,
  {32'h3fec27e8, 32'hc0b6c8e7} /* (16, 3, 18) {real, imag} */,
  {32'h410263f6, 32'hc0fdb19e} /* (16, 3, 17) {real, imag} */,
  {32'h40e36466, 32'hc0f293c8} /* (16, 3, 16) {real, imag} */,
  {32'h40416c8c, 32'hc03ae598} /* (16, 3, 15) {real, imag} */,
  {32'h3ee07330, 32'h3f8c515d} /* (16, 3, 14) {real, imag} */,
  {32'h3ff0a314, 32'hc002a08b} /* (16, 3, 13) {real, imag} */,
  {32'h40443fad, 32'hbfee4903} /* (16, 3, 12) {real, imag} */,
  {32'hbe92ce9c, 32'hc096b958} /* (16, 3, 11) {real, imag} */,
  {32'hc01f6b42, 32'h4005d2ce} /* (16, 3, 10) {real, imag} */,
  {32'hc048c97e, 32'h40b81e08} /* (16, 3, 9) {real, imag} */,
  {32'h3f572e6a, 32'h3f5f905a} /* (16, 3, 8) {real, imag} */,
  {32'hbf79ba19, 32'hbfc372bf} /* (16, 3, 7) {real, imag} */,
  {32'h3f9014a8, 32'h409ae079} /* (16, 3, 6) {real, imag} */,
  {32'hbf756298, 32'hbdb54248} /* (16, 3, 5) {real, imag} */,
  {32'hbe53f3fc, 32'h3f120640} /* (16, 3, 4) {real, imag} */,
  {32'h3fdf9c04, 32'h3f92b1ec} /* (16, 3, 3) {real, imag} */,
  {32'hc07df846, 32'h3f81e5ae} /* (16, 3, 2) {real, imag} */,
  {32'hc0b97d2f, 32'h407e7242} /* (16, 3, 1) {real, imag} */,
  {32'hc088a1c2, 32'hbe671ae7} /* (16, 3, 0) {real, imag} */,
  {32'h3f9fd2a0, 32'hbe96e502} /* (16, 2, 31) {real, imag} */,
  {32'h3eb17bd8, 32'h3fce2d1c} /* (16, 2, 30) {real, imag} */,
  {32'hbf7b8426, 32'h3fb719da} /* (16, 2, 29) {real, imag} */,
  {32'h3eccc890, 32'h402f138a} /* (16, 2, 28) {real, imag} */,
  {32'hbf2d0c20, 32'h40f31997} /* (16, 2, 27) {real, imag} */,
  {32'h404026f9, 32'h4060a98f} /* (16, 2, 26) {real, imag} */,
  {32'h3e9edd54, 32'hbfedb9c4} /* (16, 2, 25) {real, imag} */,
  {32'h3db47920, 32'hbe0e09da} /* (16, 2, 24) {real, imag} */,
  {32'hbe291e70, 32'h3ffcf4b8} /* (16, 2, 23) {real, imag} */,
  {32'h3e9d514c, 32'hbff3aa82} /* (16, 2, 22) {real, imag} */,
  {32'h4049f021, 32'h3f07ecd4} /* (16, 2, 21) {real, imag} */,
  {32'h4018b6d4, 32'h4065395c} /* (16, 2, 20) {real, imag} */,
  {32'hc0510f1c, 32'hc08f6d4c} /* (16, 2, 19) {real, imag} */,
  {32'h3fd3743a, 32'hc0bdff28} /* (16, 2, 18) {real, imag} */,
  {32'h40182738, 32'h405e25a4} /* (16, 2, 17) {real, imag} */,
  {32'h400cdc11, 32'h40b19916} /* (16, 2, 16) {real, imag} */,
  {32'h404a7d6c, 32'h40ae0ecd} /* (16, 2, 15) {real, imag} */,
  {32'h40b88aa5, 32'h3f817794} /* (16, 2, 14) {real, imag} */,
  {32'h3fadba24, 32'h3f48a415} /* (16, 2, 13) {real, imag} */,
  {32'hbff8f4b8, 32'hc01e2e3a} /* (16, 2, 12) {real, imag} */,
  {32'h3eeb9d36, 32'hc058a3aa} /* (16, 2, 11) {real, imag} */,
  {32'hc0945b94, 32'hbfcf3cac} /* (16, 2, 10) {real, imag} */,
  {32'hbfd24578, 32'hc08450f2} /* (16, 2, 9) {real, imag} */,
  {32'hbf611004, 32'hbf149b7c} /* (16, 2, 8) {real, imag} */,
  {32'hbf6979aa, 32'h4024484f} /* (16, 2, 7) {real, imag} */,
  {32'h400762f1, 32'hbf7fb14c} /* (16, 2, 6) {real, imag} */,
  {32'hbf3dc9c9, 32'hc0a023ce} /* (16, 2, 5) {real, imag} */,
  {32'hbfcf0197, 32'hbf4186ba} /* (16, 2, 4) {real, imag} */,
  {32'hbd516180, 32'hbf8bc753} /* (16, 2, 3) {real, imag} */,
  {32'hc0c6a8d7, 32'hc06d912f} /* (16, 2, 2) {real, imag} */,
  {32'hc03676b9, 32'h3fbbcd24} /* (16, 2, 1) {real, imag} */,
  {32'hbfd6c0d5, 32'h4059a6ab} /* (16, 2, 0) {real, imag} */,
  {32'hbfef768c, 32'h4015409f} /* (16, 1, 31) {real, imag} */,
  {32'hbfabcd45, 32'h40e576ca} /* (16, 1, 30) {real, imag} */,
  {32'hc0816088, 32'h407d9be4} /* (16, 1, 29) {real, imag} */,
  {32'hbfbb9008, 32'h40341764} /* (16, 1, 28) {real, imag} */,
  {32'h406344f4, 32'h3f88afeb} /* (16, 1, 27) {real, imag} */,
  {32'h3fd61d7c, 32'hc0105b66} /* (16, 1, 26) {real, imag} */,
  {32'h4037e3d6, 32'hc08bca2a} /* (16, 1, 25) {real, imag} */,
  {32'h406963b7, 32'hc0f74906} /* (16, 1, 24) {real, imag} */,
  {32'hbe899002, 32'hc044349c} /* (16, 1, 23) {real, imag} */,
  {32'h3f83972b, 32'h40a9ae34} /* (16, 1, 22) {real, imag} */,
  {32'h3efd86e0, 32'h3f251cfe} /* (16, 1, 21) {real, imag} */,
  {32'hbfa13818, 32'h3e26ecd0} /* (16, 1, 20) {real, imag} */,
  {32'hbed6f1aa, 32'hbee3aa12} /* (16, 1, 19) {real, imag} */,
  {32'hbf597ed6, 32'hc05e021a} /* (16, 1, 18) {real, imag} */,
  {32'hc01f2ab2, 32'hbfdbb298} /* (16, 1, 17) {real, imag} */,
  {32'hc083316e, 32'h4084ef0a} /* (16, 1, 16) {real, imag} */,
  {32'h3e915c20, 32'h4032f13c} /* (16, 1, 15) {real, imag} */,
  {32'h3f9f3290, 32'h3eb7be9c} /* (16, 1, 14) {real, imag} */,
  {32'h3ea25cb0, 32'hc0048cd8} /* (16, 1, 13) {real, imag} */,
  {32'h40ff49ae, 32'hbfd2f378} /* (16, 1, 12) {real, imag} */,
  {32'h40bdb6f4, 32'hc07a6260} /* (16, 1, 11) {real, imag} */,
  {32'h3fa08cc4, 32'hc04e5cff} /* (16, 1, 10) {real, imag} */,
  {32'hbfc6eb1c, 32'hbfbcc556} /* (16, 1, 9) {real, imag} */,
  {32'hc01a341a, 32'hc0851d50} /* (16, 1, 8) {real, imag} */,
  {32'h4045f472, 32'hc0802fe7} /* (16, 1, 7) {real, imag} */,
  {32'h400082bd, 32'hbf8fdec7} /* (16, 1, 6) {real, imag} */,
  {32'h409922b9, 32'hbf7615d7} /* (16, 1, 5) {real, imag} */,
  {32'h40db3c74, 32'h3e46df34} /* (16, 1, 4) {real, imag} */,
  {32'h3fa56716, 32'hbf79d241} /* (16, 1, 3) {real, imag} */,
  {32'h40581a77, 32'h3ffb1df7} /* (16, 1, 2) {real, imag} */,
  {32'h4039f0a0, 32'h4022d3d5} /* (16, 1, 1) {real, imag} */,
  {32'hbfdc126c, 32'h3f8c6f43} /* (16, 1, 0) {real, imag} */,
  {32'h40e4b7dc, 32'h00000000} /* (16, 0, 31) {real, imag} */,
  {32'h40a64f12, 32'h00000000} /* (16, 0, 30) {real, imag} */,
  {32'hbf8f814e, 32'h00000000} /* (16, 0, 29) {real, imag} */,
  {32'hbf7bfe4c, 32'h00000000} /* (16, 0, 28) {real, imag} */,
  {32'h4085ebaa, 32'h00000000} /* (16, 0, 27) {real, imag} */,
  {32'hbf0dedf0, 32'h00000000} /* (16, 0, 26) {real, imag} */,
  {32'hc06d84c3, 32'h00000000} /* (16, 0, 25) {real, imag} */,
  {32'h3ea8dac0, 32'h00000000} /* (16, 0, 24) {real, imag} */,
  {32'hbe5ab940, 32'h00000000} /* (16, 0, 23) {real, imag} */,
  {32'h3eb46778, 32'h00000000} /* (16, 0, 22) {real, imag} */,
  {32'h3f036c97, 32'h00000000} /* (16, 0, 21) {real, imag} */,
  {32'hbf38694f, 32'h00000000} /* (16, 0, 20) {real, imag} */,
  {32'hc08c95b9, 32'h00000000} /* (16, 0, 19) {real, imag} */,
  {32'hc0930ecc, 32'h00000000} /* (16, 0, 18) {real, imag} */,
  {32'hc01fe2de, 32'h00000000} /* (16, 0, 17) {real, imag} */,
  {32'h3fbe5a33, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h3f3be836, 32'h00000000} /* (16, 0, 15) {real, imag} */,
  {32'hc11de6fe, 32'h00000000} /* (16, 0, 14) {real, imag} */,
  {32'h400dde76, 32'h00000000} /* (16, 0, 13) {real, imag} */,
  {32'h405bd5da, 32'h00000000} /* (16, 0, 12) {real, imag} */,
  {32'h40142326, 32'h00000000} /* (16, 0, 11) {real, imag} */,
  {32'h40448cde, 32'h00000000} /* (16, 0, 10) {real, imag} */,
  {32'h40b99731, 32'h00000000} /* (16, 0, 9) {real, imag} */,
  {32'h3f8671d8, 32'h00000000} /* (16, 0, 8) {real, imag} */,
  {32'hc0e10814, 32'h00000000} /* (16, 0, 7) {real, imag} */,
  {32'hc0609d82, 32'h00000000} /* (16, 0, 6) {real, imag} */,
  {32'hbfc6b342, 32'h00000000} /* (16, 0, 5) {real, imag} */,
  {32'h3ec35bda, 32'h00000000} /* (16, 0, 4) {real, imag} */,
  {32'h40a971bf, 32'h00000000} /* (16, 0, 3) {real, imag} */,
  {32'h40a1b4f4, 32'h00000000} /* (16, 0, 2) {real, imag} */,
  {32'hc07a7d1e, 32'h00000000} /* (16, 0, 1) {real, imag} */,
  {32'hc0829220, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'hc0b04b4e, 32'hc01603f2} /* (15, 31, 31) {real, imag} */,
  {32'hc0726553, 32'hc0337b75} /* (15, 31, 30) {real, imag} */,
  {32'h3f9e628c, 32'hc1049f92} /* (15, 31, 29) {real, imag} */,
  {32'hbfd50b90, 32'hc09a088e} /* (15, 31, 28) {real, imag} */,
  {32'h4060479b, 32'hc05c90d8} /* (15, 31, 27) {real, imag} */,
  {32'h41091e84, 32'hbfd1fce9} /* (15, 31, 26) {real, imag} */,
  {32'h400a3258, 32'hc04a437c} /* (15, 31, 25) {real, imag} */,
  {32'h3fe6e1b2, 32'hc08e3d52} /* (15, 31, 24) {real, imag} */,
  {32'h40f10b24, 32'h3ec1605c} /* (15, 31, 23) {real, imag} */,
  {32'h411a52a8, 32'h412f7a34} /* (15, 31, 22) {real, imag} */,
  {32'h4066c540, 32'h4099e164} /* (15, 31, 21) {real, imag} */,
  {32'hc06c0376, 32'hbf0251a2} /* (15, 31, 20) {real, imag} */,
  {32'hc0393acb, 32'hc00b6022} /* (15, 31, 19) {real, imag} */,
  {32'hc04688dc, 32'hc108d2b6} /* (15, 31, 18) {real, imag} */,
  {32'hc097d76a, 32'hc0ee50d0} /* (15, 31, 17) {real, imag} */,
  {32'hc08e1ac4, 32'hc0773223} /* (15, 31, 16) {real, imag} */,
  {32'hc012310c, 32'h40049f74} /* (15, 31, 15) {real, imag} */,
  {32'hbf4cabca, 32'hc0023f45} /* (15, 31, 14) {real, imag} */,
  {32'hbfc1c8c2, 32'hc007343b} /* (15, 31, 13) {real, imag} */,
  {32'hc12e85d7, 32'hc08560da} /* (15, 31, 12) {real, imag} */,
  {32'hc122b57c, 32'hbf0530e8} /* (15, 31, 11) {real, imag} */,
  {32'hc0bcad47, 32'h409d6d0c} /* (15, 31, 10) {real, imag} */,
  {32'hbf02e02c, 32'h40b83333} /* (15, 31, 9) {real, imag} */,
  {32'h40adf0e4, 32'hbf35bfe4} /* (15, 31, 8) {real, imag} */,
  {32'hc070b976, 32'hbd971d40} /* (15, 31, 7) {real, imag} */,
  {32'hc030ab10, 32'h3f85e86f} /* (15, 31, 6) {real, imag} */,
  {32'h4080b382, 32'hbfc66730} /* (15, 31, 5) {real, imag} */,
  {32'h40d1612b, 32'hc08d16e5} /* (15, 31, 4) {real, imag} */,
  {32'h40c09228, 32'hc05c6b7c} /* (15, 31, 3) {real, imag} */,
  {32'h405e8432, 32'h40208cbf} /* (15, 31, 2) {real, imag} */,
  {32'h4069af97, 32'h4117ab48} /* (15, 31, 1) {real, imag} */,
  {32'h4008231a, 32'h40d5d816} /* (15, 31, 0) {real, imag} */,
  {32'hbebc34c8, 32'h3f410150} /* (15, 30, 31) {real, imag} */,
  {32'h409c60c0, 32'h404039c9} /* (15, 30, 30) {real, imag} */,
  {32'h40df24d7, 32'h408e5df0} /* (15, 30, 29) {real, imag} */,
  {32'h3fa1c9ae, 32'h40bd8ff2} /* (15, 30, 28) {real, imag} */,
  {32'hc06b83d3, 32'h40913d80} /* (15, 30, 27) {real, imag} */,
  {32'hbff2a8a1, 32'h40861de5} /* (15, 30, 26) {real, imag} */,
  {32'hc01ce42d, 32'h40afaabc} /* (15, 30, 25) {real, imag} */,
  {32'hc00399d0, 32'h3fc26eb8} /* (15, 30, 24) {real, imag} */,
  {32'hbf35bb9a, 32'h40324eae} /* (15, 30, 23) {real, imag} */,
  {32'hbf05b9fb, 32'hbf399438} /* (15, 30, 22) {real, imag} */,
  {32'hc002c83a, 32'hc03874dc} /* (15, 30, 21) {real, imag} */,
  {32'hbfeb4805, 32'hc0877e6f} /* (15, 30, 20) {real, imag} */,
  {32'h3edbb2c8, 32'hbfe10d04} /* (15, 30, 19) {real, imag} */,
  {32'hc0a84a2c, 32'hc0acdd05} /* (15, 30, 18) {real, imag} */,
  {32'h3fe858f7, 32'hc099eab3} /* (15, 30, 17) {real, imag} */,
  {32'h410b0161, 32'hc08205ba} /* (15, 30, 16) {real, imag} */,
  {32'h40480b68, 32'hbe28dd48} /* (15, 30, 15) {real, imag} */,
  {32'hbe6c09b0, 32'h407e3c6e} /* (15, 30, 14) {real, imag} */,
  {32'hbfaef0c4, 32'h4034a5dc} /* (15, 30, 13) {real, imag} */,
  {32'h403e325f, 32'h3f76dea1} /* (15, 30, 12) {real, imag} */,
  {32'h3fd1925d, 32'hbc24cf20} /* (15, 30, 11) {real, imag} */,
  {32'hbf983c3f, 32'hbf82ecd2} /* (15, 30, 10) {real, imag} */,
  {32'hc0bcb19f, 32'hbe5ccec0} /* (15, 30, 9) {real, imag} */,
  {32'hbe95c399, 32'h3fdac70a} /* (15, 30, 8) {real, imag} */,
  {32'hc0bac8aa, 32'hc009fe02} /* (15, 30, 7) {real, imag} */,
  {32'hc0f3dd5c, 32'h3fd2ccb2} /* (15, 30, 6) {real, imag} */,
  {32'hc0229c34, 32'h40ecfcf4} /* (15, 30, 5) {real, imag} */,
  {32'h4024cbdb, 32'h402457a3} /* (15, 30, 4) {real, imag} */,
  {32'hbf9ac4da, 32'h4047143b} /* (15, 30, 3) {real, imag} */,
  {32'hbe585588, 32'h40881ada} /* (15, 30, 2) {real, imag} */,
  {32'h405ddcbc, 32'hbfcdbd5c} /* (15, 30, 1) {real, imag} */,
  {32'h3fbe87e9, 32'hc03766e9} /* (15, 30, 0) {real, imag} */,
  {32'h40376a6b, 32'h4034bf02} /* (15, 29, 31) {real, imag} */,
  {32'h410271c2, 32'h3fafc43e} /* (15, 29, 30) {real, imag} */,
  {32'h403b6546, 32'hbf22011c} /* (15, 29, 29) {real, imag} */,
  {32'h4092b050, 32'h3c4b42c0} /* (15, 29, 28) {real, imag} */,
  {32'h40e49a31, 32'hc059348c} /* (15, 29, 27) {real, imag} */,
  {32'h4059a2ae, 32'hc0a315c9} /* (15, 29, 26) {real, imag} */,
  {32'h3ee540a4, 32'hc01dc08c} /* (15, 29, 25) {real, imag} */,
  {32'h4043c01d, 32'h4043a2e4} /* (15, 29, 24) {real, imag} */,
  {32'hc0780108, 32'hc0042a1c} /* (15, 29, 23) {real, imag} */,
  {32'h3f997a9e, 32'hc01874d6} /* (15, 29, 22) {real, imag} */,
  {32'h40ba694e, 32'hc0593582} /* (15, 29, 21) {real, imag} */,
  {32'h410c45bc, 32'hc053d776} /* (15, 29, 20) {real, imag} */,
  {32'h3fb18686, 32'h3f5155d1} /* (15, 29, 19) {real, imag} */,
  {32'hbf9e8dda, 32'h408e22e2} /* (15, 29, 18) {real, imag} */,
  {32'h4003bcc0, 32'h408662b2} /* (15, 29, 17) {real, imag} */,
  {32'hbfd51f3d, 32'h3f6c911b} /* (15, 29, 16) {real, imag} */,
  {32'h3e83472c, 32'h40116b24} /* (15, 29, 15) {real, imag} */,
  {32'hc045e41c, 32'h3f3e7a3e} /* (15, 29, 14) {real, imag} */,
  {32'hbf9f9936, 32'hbee768f8} /* (15, 29, 13) {real, imag} */,
  {32'h40a4f892, 32'h3f389210} /* (15, 29, 12) {real, imag} */,
  {32'hc03b4fc8, 32'h40247fd4} /* (15, 29, 11) {real, imag} */,
  {32'hc0a88b6a, 32'hbf73d9ac} /* (15, 29, 10) {real, imag} */,
  {32'h4079e408, 32'hc08f3581} /* (15, 29, 9) {real, imag} */,
  {32'h40c9ea16, 32'hbeb618b6} /* (15, 29, 8) {real, imag} */,
  {32'hbea0f07c, 32'hbdb7ffe0} /* (15, 29, 7) {real, imag} */,
  {32'h404b6d75, 32'hc05fbc81} /* (15, 29, 6) {real, imag} */,
  {32'h400575e7, 32'hc0869269} /* (15, 29, 5) {real, imag} */,
  {32'h3f835ea0, 32'hc03660fa} /* (15, 29, 4) {real, imag} */,
  {32'h3f2acd10, 32'hbf3a17d4} /* (15, 29, 3) {real, imag} */,
  {32'hc03fd81f, 32'h3ee0afd0} /* (15, 29, 2) {real, imag} */,
  {32'hbfde3f2e, 32'hbf2e9676} /* (15, 29, 1) {real, imag} */,
  {32'hbc96ad50, 32'hbecad3ba} /* (15, 29, 0) {real, imag} */,
  {32'hbfa1ee28, 32'hc0615624} /* (15, 28, 31) {real, imag} */,
  {32'hbff1b5e4, 32'hc0702f6c} /* (15, 28, 30) {real, imag} */,
  {32'h3f399590, 32'hbe9ae370} /* (15, 28, 29) {real, imag} */,
  {32'h4060c14e, 32'h3fb2a7be} /* (15, 28, 28) {real, imag} */,
  {32'h408aa8c8, 32'h3f127252} /* (15, 28, 27) {real, imag} */,
  {32'h3ffb4b8c, 32'h3fc30edb} /* (15, 28, 26) {real, imag} */,
  {32'hbebc0248, 32'h3ff75757} /* (15, 28, 25) {real, imag} */,
  {32'hc04ae5ec, 32'h3bc8e600} /* (15, 28, 24) {real, imag} */,
  {32'hbfafb6e0, 32'hc08b3623} /* (15, 28, 23) {real, imag} */,
  {32'hc034a490, 32'hbfa9d745} /* (15, 28, 22) {real, imag} */,
  {32'h3e683312, 32'h3fb1fdee} /* (15, 28, 21) {real, imag} */,
  {32'hbf4427b4, 32'hc02d26de} /* (15, 28, 20) {real, imag} */,
  {32'hbf965d99, 32'hc0f4ecb5} /* (15, 28, 19) {real, imag} */,
  {32'h401029e9, 32'hc13682de} /* (15, 28, 18) {real, imag} */,
  {32'h409b1a4d, 32'hc0a8d0d6} /* (15, 28, 17) {real, imag} */,
  {32'h40302bbd, 32'h40b37ff8} /* (15, 28, 16) {real, imag} */,
  {32'h3f9c3748, 32'h40a59f8b} /* (15, 28, 15) {real, imag} */,
  {32'hbe24db08, 32'h3fbad021} /* (15, 28, 14) {real, imag} */,
  {32'hbfd13ae4, 32'h3ffa363e} /* (15, 28, 13) {real, imag} */,
  {32'h3e5606b0, 32'h40c2f473} /* (15, 28, 12) {real, imag} */,
  {32'h40a12864, 32'h401aac32} /* (15, 28, 11) {real, imag} */,
  {32'h41110dc0, 32'hbf151db6} /* (15, 28, 10) {real, imag} */,
  {32'h4086c878, 32'hbffe1646} /* (15, 28, 9) {real, imag} */,
  {32'h4042e884, 32'hbe36ee10} /* (15, 28, 8) {real, imag} */,
  {32'hc003a9ca, 32'hbf864ef4} /* (15, 28, 7) {real, imag} */,
  {32'hc0b63e48, 32'hc0a931f3} /* (15, 28, 6) {real, imag} */,
  {32'hc06092d7, 32'hbf87d096} /* (15, 28, 5) {real, imag} */,
  {32'hbfe53a68, 32'hc0731691} /* (15, 28, 4) {real, imag} */,
  {32'h3fc5d74a, 32'h3faaacb5} /* (15, 28, 3) {real, imag} */,
  {32'h40296dab, 32'h40efa6c0} /* (15, 28, 2) {real, imag} */,
  {32'h3e036590, 32'h402c7b8a} /* (15, 28, 1) {real, imag} */,
  {32'h3f8cc75c, 32'hbe8d6e90} /* (15, 28, 0) {real, imag} */,
  {32'h3fd4262c, 32'h3f89f506} /* (15, 27, 31) {real, imag} */,
  {32'h3f48eb00, 32'h3f29a516} /* (15, 27, 30) {real, imag} */,
  {32'h3db7a55c, 32'h3f05cd61} /* (15, 27, 29) {real, imag} */,
  {32'h40999e24, 32'h4012f028} /* (15, 27, 28) {real, imag} */,
  {32'hc0709e04, 32'h3f5cd628} /* (15, 27, 27) {real, imag} */,
  {32'hc0957004, 32'hbf923b2e} /* (15, 27, 26) {real, imag} */,
  {32'hc001fccf, 32'h40383031} /* (15, 27, 25) {real, imag} */,
  {32'hc0ac982c, 32'h4061d250} /* (15, 27, 24) {real, imag} */,
  {32'hc000e26b, 32'h3ebe937c} /* (15, 27, 23) {real, imag} */,
  {32'h402b5320, 32'hc01c2572} /* (15, 27, 22) {real, imag} */,
  {32'hc0379d7b, 32'hc005c134} /* (15, 27, 21) {real, imag} */,
  {32'hc0bc04fd, 32'hc0389023} /* (15, 27, 20) {real, imag} */,
  {32'hc044831f, 32'hbfccc68e} /* (15, 27, 19) {real, imag} */,
  {32'hbfd17cbc, 32'h3e0a9bf8} /* (15, 27, 18) {real, imag} */,
  {32'h3fb651dd, 32'hbf1247af} /* (15, 27, 17) {real, imag} */,
  {32'h40892990, 32'hbf9fbc82} /* (15, 27, 16) {real, imag} */,
  {32'h402ffee0, 32'hc0c1f2ed} /* (15, 27, 15) {real, imag} */,
  {32'h40dc6061, 32'hc09f7608} /* (15, 27, 14) {real, imag} */,
  {32'h413769c0, 32'h4040d164} /* (15, 27, 13) {real, imag} */,
  {32'h412804d8, 32'h405b64f4} /* (15, 27, 12) {real, imag} */,
  {32'h4045b9ea, 32'h4021980b} /* (15, 27, 11) {real, imag} */,
  {32'hc0246f6e, 32'h4064c0f1} /* (15, 27, 10) {real, imag} */,
  {32'hbfbf6fb2, 32'h3fdae8d0} /* (15, 27, 9) {real, imag} */,
  {32'h40091208, 32'h3faf3cdf} /* (15, 27, 8) {real, imag} */,
  {32'h3f63a7b6, 32'h3fe2417c} /* (15, 27, 7) {real, imag} */,
  {32'hc035a47e, 32'h403d4bf2} /* (15, 27, 6) {real, imag} */,
  {32'hc091c5f8, 32'h3ff0d8c3} /* (15, 27, 5) {real, imag} */,
  {32'hbfb013cb, 32'h401131a4} /* (15, 27, 4) {real, imag} */,
  {32'h4000e1a2, 32'hc047dcdd} /* (15, 27, 3) {real, imag} */,
  {32'h40b06955, 32'h3f8487d6} /* (15, 27, 2) {real, imag} */,
  {32'h3f051808, 32'h409db2b8} /* (15, 27, 1) {real, imag} */,
  {32'h3fd34826, 32'h40aab673} /* (15, 27, 0) {real, imag} */,
  {32'hbfbff6ac, 32'hbfe6cc60} /* (15, 26, 31) {real, imag} */,
  {32'hc0225a1c, 32'hbfd8738d} /* (15, 26, 30) {real, imag} */,
  {32'hc06f8e0a, 32'hc022ea19} /* (15, 26, 29) {real, imag} */,
  {32'h3ef12d20, 32'hbf062936} /* (15, 26, 28) {real, imag} */,
  {32'hc019591e, 32'hbe2e1184} /* (15, 26, 27) {real, imag} */,
  {32'hbf8816a8, 32'h40322dac} /* (15, 26, 26) {real, imag} */,
  {32'hbf65ca23, 32'h40859eb9} /* (15, 26, 25) {real, imag} */,
  {32'hc018863c, 32'h3fabb8e5} /* (15, 26, 24) {real, imag} */,
  {32'hc0404d5f, 32'hbff38e5a} /* (15, 26, 23) {real, imag} */,
  {32'hbf94678b, 32'h3f1d9626} /* (15, 26, 22) {real, imag} */,
  {32'h3fce9199, 32'h4019322a} /* (15, 26, 21) {real, imag} */,
  {32'h3ffb27c7, 32'h3fc0aeb6} /* (15, 26, 20) {real, imag} */,
  {32'hc011f192, 32'h3f4d3bb6} /* (15, 26, 19) {real, imag} */,
  {32'hc0226e0d, 32'h3f2aeb1c} /* (15, 26, 18) {real, imag} */,
  {32'h4019b273, 32'hbfda0954} /* (15, 26, 17) {real, imag} */,
  {32'hc0890d88, 32'hc00772cf} /* (15, 26, 16) {real, imag} */,
  {32'hc05f1ade, 32'hc04e4c6a} /* (15, 26, 15) {real, imag} */,
  {32'h4033f0c0, 32'hbf4b7c83} /* (15, 26, 14) {real, imag} */,
  {32'h3fdc2b81, 32'hc0bf1649} /* (15, 26, 13) {real, imag} */,
  {32'h408e0aeb, 32'hc0d11a10} /* (15, 26, 12) {real, imag} */,
  {32'h40723323, 32'hc076e7a8} /* (15, 26, 11) {real, imag} */,
  {32'h3f8aaf12, 32'h3ec019c4} /* (15, 26, 10) {real, imag} */,
  {32'h3f9f5b05, 32'hbf298414} /* (15, 26, 9) {real, imag} */,
  {32'h3fd8ae86, 32'hc09f7bd4} /* (15, 26, 8) {real, imag} */,
  {32'hc00d9b47, 32'hc02871ee} /* (15, 26, 7) {real, imag} */,
  {32'hc0854dbb, 32'hc07480f3} /* (15, 26, 6) {real, imag} */,
  {32'hc0eab509, 32'hc01ce888} /* (15, 26, 5) {real, imag} */,
  {32'hc02f332a, 32'hc0486bfd} /* (15, 26, 4) {real, imag} */,
  {32'hc05aa607, 32'hbf2554bc} /* (15, 26, 3) {real, imag} */,
  {32'hc0bb0e0e, 32'h40a21eea} /* (15, 26, 2) {real, imag} */,
  {32'hc02c0ef8, 32'h3de0f9c0} /* (15, 26, 1) {real, imag} */,
  {32'hc0899c30, 32'hc08396ac} /* (15, 26, 0) {real, imag} */,
  {32'h3e010774, 32'h3f24eced} /* (15, 25, 31) {real, imag} */,
  {32'hc051079e, 32'h4025377b} /* (15, 25, 30) {real, imag} */,
  {32'hc0ab25e6, 32'hbfb3c492} /* (15, 25, 29) {real, imag} */,
  {32'hc0ac6ec4, 32'hbfec18ca} /* (15, 25, 28) {real, imag} */,
  {32'hc0748056, 32'h4032a1ea} /* (15, 25, 27) {real, imag} */,
  {32'hc0b9aa68, 32'h40821e3f} /* (15, 25, 26) {real, imag} */,
  {32'hc06c41d0, 32'hbf5754f8} /* (15, 25, 25) {real, imag} */,
  {32'h3fcbd09c, 32'h3fbedb41} /* (15, 25, 24) {real, imag} */,
  {32'h3f20ef40, 32'h3fe0f17e} /* (15, 25, 23) {real, imag} */,
  {32'hbf10284c, 32'hbfdc33c1} /* (15, 25, 22) {real, imag} */,
  {32'hc04971d8, 32'h3e112c58} /* (15, 25, 21) {real, imag} */,
  {32'h3f687bc4, 32'h4085f747} /* (15, 25, 20) {real, imag} */,
  {32'h3d0583e0, 32'hbec5fef4} /* (15, 25, 19) {real, imag} */,
  {32'hbd63b3c0, 32'h40529fd9} /* (15, 25, 18) {real, imag} */,
  {32'h3fdd41df, 32'h40b5cbe7} /* (15, 25, 17) {real, imag} */,
  {32'hc0249d77, 32'h40891d6f} /* (15, 25, 16) {real, imag} */,
  {32'hc0492019, 32'h3ebbd55b} /* (15, 25, 15) {real, imag} */,
  {32'hc017bd5f, 32'hbfe65f28} /* (15, 25, 14) {real, imag} */,
  {32'h3f2f610c, 32'hc002bd47} /* (15, 25, 13) {real, imag} */,
  {32'hbecf0c80, 32'h4024bff3} /* (15, 25, 12) {real, imag} */,
  {32'hc0175094, 32'hbf591ede} /* (15, 25, 11) {real, imag} */,
  {32'hbfb00e47, 32'hc010def5} /* (15, 25, 10) {real, imag} */,
  {32'hbf22b06a, 32'h40099c40} /* (15, 25, 9) {real, imag} */,
  {32'hbe0996f0, 32'hbdc3c670} /* (15, 25, 8) {real, imag} */,
  {32'hc00740be, 32'h3dd82378} /* (15, 25, 7) {real, imag} */,
  {32'hc085535e, 32'hc00e9bf0} /* (15, 25, 6) {real, imag} */,
  {32'hbf7ebee8, 32'hc08d955a} /* (15, 25, 5) {real, imag} */,
  {32'hc004dcef, 32'h3f343b70} /* (15, 25, 4) {real, imag} */,
  {32'h3fca8819, 32'hbe845c1c} /* (15, 25, 3) {real, imag} */,
  {32'h3ff33f12, 32'hbeccbd10} /* (15, 25, 2) {real, imag} */,
  {32'h3f47183f, 32'hc032d980} /* (15, 25, 1) {real, imag} */,
  {32'hc0425ee5, 32'h3e537490} /* (15, 25, 0) {real, imag} */,
  {32'hc0018f4a, 32'hc0439232} /* (15, 24, 31) {real, imag} */,
  {32'hbfc83e64, 32'h3d26c6c0} /* (15, 24, 30) {real, imag} */,
  {32'hbeb2b158, 32'h3f8a34eb} /* (15, 24, 29) {real, imag} */,
  {32'hbec43580, 32'h3e4f7628} /* (15, 24, 28) {real, imag} */,
  {32'hbf87546a, 32'h3f31791c} /* (15, 24, 27) {real, imag} */,
  {32'hbf7a59cb, 32'h3fc8f6da} /* (15, 24, 26) {real, imag} */,
  {32'h3efe3164, 32'hc04f0a01} /* (15, 24, 25) {real, imag} */,
  {32'h3fb84696, 32'hc02b45bf} /* (15, 24, 24) {real, imag} */,
  {32'h4012fe10, 32'hc00916be} /* (15, 24, 23) {real, imag} */,
  {32'h3fddefa8, 32'hbeba0de0} /* (15, 24, 22) {real, imag} */,
  {32'h402ad772, 32'h3f68a598} /* (15, 24, 21) {real, imag} */,
  {32'h40862c4e, 32'h40058821} /* (15, 24, 20) {real, imag} */,
  {32'h4085d2b1, 32'h3fe8b093} /* (15, 24, 19) {real, imag} */,
  {32'h3ff6f69b, 32'h3f1f0920} /* (15, 24, 18) {real, imag} */,
  {32'h3f42cfe4, 32'hc0340d74} /* (15, 24, 17) {real, imag} */,
  {32'h3fa43f62, 32'hc07a42c5} /* (15, 24, 16) {real, imag} */,
  {32'hbc973bc0, 32'hbf9817de} /* (15, 24, 15) {real, imag} */,
  {32'hc04763f0, 32'h3f86245c} /* (15, 24, 14) {real, imag} */,
  {32'hc07fa31f, 32'h40ca8a22} /* (15, 24, 13) {real, imag} */,
  {32'hc0149928, 32'h403c391e} /* (15, 24, 12) {real, imag} */,
  {32'hbe1b8de4, 32'hc02e8f14} /* (15, 24, 11) {real, imag} */,
  {32'h3fb794fc, 32'hc04bef81} /* (15, 24, 10) {real, imag} */,
  {32'hbef208a8, 32'hbe3af2b0} /* (15, 24, 9) {real, imag} */,
  {32'h3f72d71e, 32'h3f92b474} /* (15, 24, 8) {real, imag} */,
  {32'hc07b6d76, 32'hbf94b4b8} /* (15, 24, 7) {real, imag} */,
  {32'hbfef4b34, 32'h40769d60} /* (15, 24, 6) {real, imag} */,
  {32'hbafeb800, 32'h3eb09c4c} /* (15, 24, 5) {real, imag} */,
  {32'hbf777724, 32'hbeda5fd8} /* (15, 24, 4) {real, imag} */,
  {32'h3e1ac068, 32'hc0222c3f} /* (15, 24, 3) {real, imag} */,
  {32'hbe559288, 32'hc046f80d} /* (15, 24, 2) {real, imag} */,
  {32'hbf08b7e5, 32'hc008c2ec} /* (15, 24, 1) {real, imag} */,
  {32'h3edab2a2, 32'hbf409dbc} /* (15, 24, 0) {real, imag} */,
  {32'hc014188d, 32'hbf5359ce} /* (15, 23, 31) {real, imag} */,
  {32'hc0187b96, 32'h3f714be7} /* (15, 23, 30) {real, imag} */,
  {32'h3f88c6f7, 32'h3fd2c606} /* (15, 23, 29) {real, imag} */,
  {32'h3fae3b13, 32'hc027de5c} /* (15, 23, 28) {real, imag} */,
  {32'h3f01fc14, 32'hbfa704ec} /* (15, 23, 27) {real, imag} */,
  {32'hbf2c8720, 32'h3f15d35e} /* (15, 23, 26) {real, imag} */,
  {32'h3ed0a418, 32'hbf4cedea} /* (15, 23, 25) {real, imag} */,
  {32'h3f7d2e3f, 32'hc04bec70} /* (15, 23, 24) {real, imag} */,
  {32'hbf8c07ac, 32'hc0758438} /* (15, 23, 23) {real, imag} */,
  {32'hc0574ac6, 32'hc08c5b63} /* (15, 23, 22) {real, imag} */,
  {32'h400889b5, 32'hc04174e5} /* (15, 23, 21) {real, imag} */,
  {32'h3fb9e475, 32'hc055d239} /* (15, 23, 20) {real, imag} */,
  {32'hc072f5c3, 32'h3e7b2630} /* (15, 23, 19) {real, imag} */,
  {32'h3f2a30d8, 32'h3f9ad40d} /* (15, 23, 18) {real, imag} */,
  {32'h3f9bc783, 32'hc03377e0} /* (15, 23, 17) {real, imag} */,
  {32'hbe9d1fae, 32'hc04c9f1d} /* (15, 23, 16) {real, imag} */,
  {32'h3ff63816, 32'hbf09cdec} /* (15, 23, 15) {real, imag} */,
  {32'h40a935c0, 32'h3fc009b0} /* (15, 23, 14) {real, imag} */,
  {32'h40d72adc, 32'hbe198b18} /* (15, 23, 13) {real, imag} */,
  {32'h3f17cb60, 32'hbfae3bda} /* (15, 23, 12) {real, imag} */,
  {32'hbf594756, 32'hbd866d80} /* (15, 23, 11) {real, imag} */,
  {32'hc0319166, 32'h3eeee7c2} /* (15, 23, 10) {real, imag} */,
  {32'hc09d0cff, 32'hbef6346c} /* (15, 23, 9) {real, imag} */,
  {32'hc07cace5, 32'hc0596441} /* (15, 23, 8) {real, imag} */,
  {32'hc05ddc0a, 32'hbfd611fc} /* (15, 23, 7) {real, imag} */,
  {32'h3e793b10, 32'hbac53800} /* (15, 23, 6) {real, imag} */,
  {32'h402eb922, 32'hbfb0ffdc} /* (15, 23, 5) {real, imag} */,
  {32'h404017e2, 32'hbf8e5188} /* (15, 23, 4) {real, imag} */,
  {32'h3ed7e27c, 32'hc017d6a4} /* (15, 23, 3) {real, imag} */,
  {32'hbf6267a0, 32'hbea99c60} /* (15, 23, 2) {real, imag} */,
  {32'h3ed4f790, 32'h3f5743e2} /* (15, 23, 1) {real, imag} */,
  {32'hbfb93156, 32'hbf7f54c0} /* (15, 23, 0) {real, imag} */,
  {32'hbe56809c, 32'hc0371295} /* (15, 22, 31) {real, imag} */,
  {32'h3f3156b0, 32'hc08e1444} /* (15, 22, 30) {real, imag} */,
  {32'hc0257dc0, 32'hbfd568b8} /* (15, 22, 29) {real, imag} */,
  {32'hc01c706c, 32'hbfd2d315} /* (15, 22, 28) {real, imag} */,
  {32'hbe9b8a74, 32'hc01a33b9} /* (15, 22, 27) {real, imag} */,
  {32'h3db630e0, 32'hc0357f8a} /* (15, 22, 26) {real, imag} */,
  {32'hbfefb842, 32'hc096c8c3} /* (15, 22, 25) {real, imag} */,
  {32'hbfe46ac7, 32'hc0690e99} /* (15, 22, 24) {real, imag} */,
  {32'h4033ef27, 32'hc0be217a} /* (15, 22, 23) {real, imag} */,
  {32'h408834a3, 32'hbfbe2f33} /* (15, 22, 22) {real, imag} */,
  {32'h3f4bf526, 32'h3f656ce8} /* (15, 22, 21) {real, imag} */,
  {32'h3fb9ba0f, 32'hbeb3f884} /* (15, 22, 20) {real, imag} */,
  {32'hbef80e0c, 32'h3f232e02} /* (15, 22, 19) {real, imag} */,
  {32'hbf0cfe6b, 32'hbea95598} /* (15, 22, 18) {real, imag} */,
  {32'h3fabba7a, 32'hbf993496} /* (15, 22, 17) {real, imag} */,
  {32'h4006b866, 32'h3fd7e88f} /* (15, 22, 16) {real, imag} */,
  {32'h3fee24c1, 32'h4038e89f} /* (15, 22, 15) {real, imag} */,
  {32'h4085b272, 32'h40151413} /* (15, 22, 14) {real, imag} */,
  {32'h4052b18e, 32'hb90fa000} /* (15, 22, 13) {real, imag} */,
  {32'h3f5b2aa0, 32'h3e79e760} /* (15, 22, 12) {real, imag} */,
  {32'hbf18d89b, 32'h3fbcf747} /* (15, 22, 11) {real, imag} */,
  {32'hbf1d8366, 32'h3ff398c6} /* (15, 22, 10) {real, imag} */,
  {32'h3ffaaee2, 32'h3ec0746d} /* (15, 22, 9) {real, imag} */,
  {32'h3f83d99a, 32'hbff60fe2} /* (15, 22, 8) {real, imag} */,
  {32'h406c3300, 32'h40314f8c} /* (15, 22, 7) {real, imag} */,
  {32'h3fa207db, 32'h3f02d1ca} /* (15, 22, 6) {real, imag} */,
  {32'hc05d8e72, 32'hbe9eae1a} /* (15, 22, 5) {real, imag} */,
  {32'hc03c9644, 32'h3f3d81f8} /* (15, 22, 4) {real, imag} */,
  {32'hc076e614, 32'h403320e9} /* (15, 22, 3) {real, imag} */,
  {32'hc02ae67d, 32'h3f7319fc} /* (15, 22, 2) {real, imag} */,
  {32'hc007baba, 32'h3ebe1cc2} /* (15, 22, 1) {real, imag} */,
  {32'hbecf0cb3, 32'hbd981230} /* (15, 22, 0) {real, imag} */,
  {32'hbf912e4a, 32'hbd7a5c80} /* (15, 21, 31) {real, imag} */,
  {32'hbfae47be, 32'hbfa64088} /* (15, 21, 30) {real, imag} */,
  {32'hbf79aaac, 32'hbe23a990} /* (15, 21, 29) {real, imag} */,
  {32'hc045fa4e, 32'hbfdc3edf} /* (15, 21, 28) {real, imag} */,
  {32'hc022c224, 32'hbf6acbbe} /* (15, 21, 27) {real, imag} */,
  {32'hc00ef130, 32'hc015b612} /* (15, 21, 26) {real, imag} */,
  {32'h3eb7f328, 32'h3efc4698} /* (15, 21, 25) {real, imag} */,
  {32'h3fe5c4da, 32'h401c0105} /* (15, 21, 24) {real, imag} */,
  {32'h3d928904, 32'h403b45c0} /* (15, 21, 23) {real, imag} */,
  {32'hbfb2f644, 32'h3ffd8b25} /* (15, 21, 22) {real, imag} */,
  {32'h3f81f313, 32'hbfc57f58} /* (15, 21, 21) {real, imag} */,
  {32'h3f934b0d, 32'hc0249bcd} /* (15, 21, 20) {real, imag} */,
  {32'h402944f5, 32'hbfc37482} /* (15, 21, 19) {real, imag} */,
  {32'h404cb73b, 32'hbeb4fe52} /* (15, 21, 18) {real, imag} */,
  {32'h4009102c, 32'h4016c70e} /* (15, 21, 17) {real, imag} */,
  {32'h400b94a0, 32'h3faa768d} /* (15, 21, 16) {real, imag} */,
  {32'hbf93585b, 32'h3fa0756b} /* (15, 21, 15) {real, imag} */,
  {32'hbfd618c2, 32'h3fbd7462} /* (15, 21, 14) {real, imag} */,
  {32'h3fa377d4, 32'hbf935078} /* (15, 21, 13) {real, imag} */,
  {32'hbfc4fb32, 32'hbfc49493} /* (15, 21, 12) {real, imag} */,
  {32'hc00ee098, 32'hbe2a0e60} /* (15, 21, 11) {real, imag} */,
  {32'hbed86afc, 32'h40597172} /* (15, 21, 10) {real, imag} */,
  {32'hbf007e30, 32'h404f1834} /* (15, 21, 9) {real, imag} */,
  {32'hbecafd6e, 32'h3f23e312} /* (15, 21, 8) {real, imag} */,
  {32'h402901b4, 32'h3f70517e} /* (15, 21, 7) {real, imag} */,
  {32'h3ff8dade, 32'h3f9ed49e} /* (15, 21, 6) {real, imag} */,
  {32'hbda4fba0, 32'h3f97b8ba} /* (15, 21, 5) {real, imag} */,
  {32'hbd452090, 32'h406105a5} /* (15, 21, 4) {real, imag} */,
  {32'h3f878cc5, 32'h3f542469} /* (15, 21, 3) {real, imag} */,
  {32'h404fbcc3, 32'hbfaab107} /* (15, 21, 2) {real, imag} */,
  {32'h3fb3be86, 32'hbf02cd00} /* (15, 21, 1) {real, imag} */,
  {32'hbf40e561, 32'hbf304216} /* (15, 21, 0) {real, imag} */,
  {32'hbf66616b, 32'h3f838547} /* (15, 20, 31) {real, imag} */,
  {32'hbc3c8d80, 32'h3c5548c0} /* (15, 20, 30) {real, imag} */,
  {32'h3ed400ec, 32'h4003b51a} /* (15, 20, 29) {real, imag} */,
  {32'hbf87a557, 32'h4004db14} /* (15, 20, 28) {real, imag} */,
  {32'hbfd3740c, 32'h3f9be794} /* (15, 20, 27) {real, imag} */,
  {32'hbf8ec366, 32'h3f1dbce6} /* (15, 20, 26) {real, imag} */,
  {32'h3ea85378, 32'h3e34b818} /* (15, 20, 25) {real, imag} */,
  {32'hc00a1a1d, 32'h3c129600} /* (15, 20, 24) {real, imag} */,
  {32'hbf80910c, 32'hbb5fba00} /* (15, 20, 23) {real, imag} */,
  {32'h3e704768, 32'hbf88ebc7} /* (15, 20, 22) {real, imag} */,
  {32'h3e51d76c, 32'h3f475e33} /* (15, 20, 21) {real, imag} */,
  {32'h3f374d2a, 32'h3eed4a56} /* (15, 20, 20) {real, imag} */,
  {32'hbf6263ea, 32'h3e175dd0} /* (15, 20, 19) {real, imag} */,
  {32'hbec5fc1a, 32'h3f167042} /* (15, 20, 18) {real, imag} */,
  {32'h400de298, 32'hc00fe3c2} /* (15, 20, 17) {real, imag} */,
  {32'h3ffb031e, 32'hbf5c349a} /* (15, 20, 16) {real, imag} */,
  {32'h3f42b17e, 32'h3e2b83e8} /* (15, 20, 15) {real, imag} */,
  {32'h3f6451ce, 32'hbea2fb82} /* (15, 20, 14) {real, imag} */,
  {32'hbdcc0400, 32'h3febf9b6} /* (15, 20, 13) {real, imag} */,
  {32'h400ecfb4, 32'h402cbb0b} /* (15, 20, 12) {real, imag} */,
  {32'h3f8f1c07, 32'h40074306} /* (15, 20, 11) {real, imag} */,
  {32'h3e65dd58, 32'h3eb95db0} /* (15, 20, 10) {real, imag} */,
  {32'h401d59c2, 32'hbff9e8d7} /* (15, 20, 9) {real, imag} */,
  {32'h3f21c1a7, 32'h3d575b80} /* (15, 20, 8) {real, imag} */,
  {32'h3e53f57c, 32'h4049b3e4} /* (15, 20, 7) {real, imag} */,
  {32'h3f455ea5, 32'h3f5efd24} /* (15, 20, 6) {real, imag} */,
  {32'hbf0d3949, 32'hbf491c46} /* (15, 20, 5) {real, imag} */,
  {32'h3fdbf32a, 32'hbebb99f8} /* (15, 20, 4) {real, imag} */,
  {32'hbbdb15c0, 32'h3d4a4860} /* (15, 20, 3) {real, imag} */,
  {32'hbefe1ae6, 32'hc02f7cf2} /* (15, 20, 2) {real, imag} */,
  {32'hbfda46cc, 32'hc028f29e} /* (15, 20, 1) {real, imag} */,
  {32'h3e71af68, 32'h3ea9ca8b} /* (15, 20, 0) {real, imag} */,
  {32'h3ef1ba54, 32'hbeba0828} /* (15, 19, 31) {real, imag} */,
  {32'hbead8a34, 32'hbf08b5cc} /* (15, 19, 30) {real, imag} */,
  {32'h3f009f7c, 32'h3f462760} /* (15, 19, 29) {real, imag} */,
  {32'h40817326, 32'hbf0127b2} /* (15, 19, 28) {real, imag} */,
  {32'h4026b21a, 32'h3ef33a88} /* (15, 19, 27) {real, imag} */,
  {32'h3f063681, 32'h3fca474d} /* (15, 19, 26) {real, imag} */,
  {32'hbfb496e7, 32'h3f1302c7} /* (15, 19, 25) {real, imag} */,
  {32'hbe7c1e8c, 32'h3e55287c} /* (15, 19, 24) {real, imag} */,
  {32'hbf042156, 32'h3f85ec8c} /* (15, 19, 23) {real, imag} */,
  {32'hbf33c84b, 32'h3f2332a6} /* (15, 19, 22) {real, imag} */,
  {32'hbf664777, 32'h3f8ea571} /* (15, 19, 21) {real, imag} */,
  {32'hbf0fb47c, 32'hbfc08ac4} /* (15, 19, 20) {real, imag} */,
  {32'hbf2cdb59, 32'hbe16accb} /* (15, 19, 19) {real, imag} */,
  {32'hbf920d33, 32'hbf88ae48} /* (15, 19, 18) {real, imag} */,
  {32'hbf870779, 32'h3cd82980} /* (15, 19, 17) {real, imag} */,
  {32'hbea6fda4, 32'h40313045} /* (15, 19, 16) {real, imag} */,
  {32'hbd0a31e0, 32'h3f76836e} /* (15, 19, 15) {real, imag} */,
  {32'hbf4bff87, 32'h3acf5a00} /* (15, 19, 14) {real, imag} */,
  {32'hbe8a3c2c, 32'hbf6aedbf} /* (15, 19, 13) {real, imag} */,
  {32'h3e8dedc0, 32'hbeb9aff0} /* (15, 19, 12) {real, imag} */,
  {32'hbf309a9e, 32'h3ebd7f3a} /* (15, 19, 11) {real, imag} */,
  {32'hbf8fc0a0, 32'h3f32f5a6} /* (15, 19, 10) {real, imag} */,
  {32'hbcbe0cc0, 32'h3f797f04} /* (15, 19, 9) {real, imag} */,
  {32'h3f9c328b, 32'h3f5b215d} /* (15, 19, 8) {real, imag} */,
  {32'h3f16028d, 32'h3ef1ef20} /* (15, 19, 7) {real, imag} */,
  {32'h3f16df58, 32'h3ee07be0} /* (15, 19, 6) {real, imag} */,
  {32'hbf1b014d, 32'hbfb29b5e} /* (15, 19, 5) {real, imag} */,
  {32'hbf8c6635, 32'hbf6272b8} /* (15, 19, 4) {real, imag} */,
  {32'h3d2e52e0, 32'hbfed671c} /* (15, 19, 3) {real, imag} */,
  {32'hbfc3bd7c, 32'hc001f4b0} /* (15, 19, 2) {real, imag} */,
  {32'h3f2d9c09, 32'h3d23ef60} /* (15, 19, 1) {real, imag} */,
  {32'h3f236374, 32'h3f8ac56e} /* (15, 19, 0) {real, imag} */,
  {32'h3ee4c44a, 32'h3e3a44dc} /* (15, 18, 31) {real, imag} */,
  {32'hbfb39a7d, 32'h3fb89e67} /* (15, 18, 30) {real, imag} */,
  {32'hbf8ffe3f, 32'hbf78ddbc} /* (15, 18, 29) {real, imag} */,
  {32'h3e899e33, 32'hbf87721a} /* (15, 18, 28) {real, imag} */,
  {32'h3fe3e40a, 32'h3d02c5c0} /* (15, 18, 27) {real, imag} */,
  {32'h3ec733a0, 32'hbe6b10a8} /* (15, 18, 26) {real, imag} */,
  {32'hbf674448, 32'hbf0df8bd} /* (15, 18, 25) {real, imag} */,
  {32'h3e028614, 32'hbf61bd90} /* (15, 18, 24) {real, imag} */,
  {32'h3f14a477, 32'hbfb7a6aa} /* (15, 18, 23) {real, imag} */,
  {32'hbf9ca65c, 32'hbf318110} /* (15, 18, 22) {real, imag} */,
  {32'hbff8f48c, 32'hbf2363f2} /* (15, 18, 21) {real, imag} */,
  {32'hbf6941bd, 32'h3e1aea2c} /* (15, 18, 20) {real, imag} */,
  {32'h3f1a003a, 32'hbf2d4328} /* (15, 18, 19) {real, imag} */,
  {32'h3fe0ac82, 32'hbf41742a} /* (15, 18, 18) {real, imag} */,
  {32'h3eacda80, 32'hbf77f00c} /* (15, 18, 17) {real, imag} */,
  {32'h3ebcfa90, 32'hbf74861c} /* (15, 18, 16) {real, imag} */,
  {32'hbe6163cc, 32'h3e408860} /* (15, 18, 15) {real, imag} */,
  {32'hbee042a2, 32'h3f0fbc3d} /* (15, 18, 14) {real, imag} */,
  {32'hbf0164e3, 32'h3f49846f} /* (15, 18, 13) {real, imag} */,
  {32'hbf4ff0a5, 32'hbfbd1166} /* (15, 18, 12) {real, imag} */,
  {32'hbf3cb0dc, 32'hbe304d1e} /* (15, 18, 11) {real, imag} */,
  {32'hbfb30190, 32'hbf90d5cf} /* (15, 18, 10) {real, imag} */,
  {32'hbe9c66d6, 32'hbebb88ec} /* (15, 18, 9) {real, imag} */,
  {32'hbfef94e7, 32'h3faf3972} /* (15, 18, 8) {real, imag} */,
  {32'hbfdccecd, 32'h3fc04b06} /* (15, 18, 7) {real, imag} */,
  {32'h3f565cf7, 32'h3ef9aa62} /* (15, 18, 6) {real, imag} */,
  {32'h3f7be5ba, 32'h3f0efcb1} /* (15, 18, 5) {real, imag} */,
  {32'h3f32e0e4, 32'hbf94cb59} /* (15, 18, 4) {real, imag} */,
  {32'hbe26fbb4, 32'hbd8b4b40} /* (15, 18, 3) {real, imag} */,
  {32'hbe8ef14c, 32'h3f7225eb} /* (15, 18, 2) {real, imag} */,
  {32'h4078d6ce, 32'hbf0ca1e4} /* (15, 18, 1) {real, imag} */,
  {32'h403e60a0, 32'hbf75cf3f} /* (15, 18, 0) {real, imag} */,
  {32'hbe71da70, 32'h3f30d078} /* (15, 17, 31) {real, imag} */,
  {32'h3f6e9a7d, 32'h3fb6dc2b} /* (15, 17, 30) {real, imag} */,
  {32'hbe28847c, 32'h3f45fc1a} /* (15, 17, 29) {real, imag} */,
  {32'hbf8464cc, 32'h3f13f9da} /* (15, 17, 28) {real, imag} */,
  {32'h3dc99480, 32'h3f177b63} /* (15, 17, 27) {real, imag} */,
  {32'hbd675b80, 32'h3f02e0c2} /* (15, 17, 26) {real, imag} */,
  {32'hbf6406ec, 32'h3da86c98} /* (15, 17, 25) {real, imag} */,
  {32'h3f778d2f, 32'hbf7b67ac} /* (15, 17, 24) {real, imag} */,
  {32'h3e929b92, 32'hbd64e580} /* (15, 17, 23) {real, imag} */,
  {32'h3de45bc0, 32'h3fc0d4bf} /* (15, 17, 22) {real, imag} */,
  {32'h3ec22ead, 32'hbf4f655a} /* (15, 17, 21) {real, imag} */,
  {32'h3e71922c, 32'hbfef656e} /* (15, 17, 20) {real, imag} */,
  {32'h3e0e1a60, 32'hbee15d52} /* (15, 17, 19) {real, imag} */,
  {32'hbf4a8b27, 32'hbf8214fa} /* (15, 17, 18) {real, imag} */,
  {32'hbe2ab1d0, 32'hbf295a4e} /* (15, 17, 17) {real, imag} */,
  {32'h3f1a6135, 32'hbe8509d6} /* (15, 17, 16) {real, imag} */,
  {32'h3d059a00, 32'hbef08b78} /* (15, 17, 15) {real, imag} */,
  {32'hbf233a8a, 32'h3d7422a0} /* (15, 17, 14) {real, imag} */,
  {32'hbe4e6d28, 32'h3e557d58} /* (15, 17, 13) {real, imag} */,
  {32'h3edc4e20, 32'h3f4c645c} /* (15, 17, 12) {real, imag} */,
  {32'h3f7314c4, 32'h3eeafc8c} /* (15, 17, 11) {real, imag} */,
  {32'h3d5ee700, 32'h3f1d14f0} /* (15, 17, 10) {real, imag} */,
  {32'hbfbfe41c, 32'h3f86e162} /* (15, 17, 9) {real, imag} */,
  {32'hbf1ac21a, 32'h3f12882c} /* (15, 17, 8) {real, imag} */,
  {32'hbd7e89c0, 32'hbdfa5ce0} /* (15, 17, 7) {real, imag} */,
  {32'h3e52c2dc, 32'h3ef7ee2c} /* (15, 17, 6) {real, imag} */,
  {32'h3eebf058, 32'h3f266353} /* (15, 17, 5) {real, imag} */,
  {32'hbe59b528, 32'h3eb6497e} /* (15, 17, 4) {real, imag} */,
  {32'hbf5ed579, 32'h400e5536} /* (15, 17, 3) {real, imag} */,
  {32'h3f73dc64, 32'h3eb938a4} /* (15, 17, 2) {real, imag} */,
  {32'h3e94df76, 32'h3f2cd354} /* (15, 17, 1) {real, imag} */,
  {32'hbe9e4514, 32'h3f8038c2} /* (15, 17, 0) {real, imag} */,
  {32'h3f49104c, 32'hbf6420d0} /* (15, 16, 31) {real, imag} */,
  {32'h3ea25bf8, 32'hbfb4f2ce} /* (15, 16, 30) {real, imag} */,
  {32'h3f0abdbe, 32'hbebc2a00} /* (15, 16, 29) {real, imag} */,
  {32'h3f3cfef8, 32'h3f3bc0a8} /* (15, 16, 28) {real, imag} */,
  {32'hbd851538, 32'h3f6bcc44} /* (15, 16, 27) {real, imag} */,
  {32'hbf6156b2, 32'h3f54f0d0} /* (15, 16, 26) {real, imag} */,
  {32'h3ed0b3c4, 32'h3e9d8c18} /* (15, 16, 25) {real, imag} */,
  {32'h3f6adb39, 32'hbf3d1ab4} /* (15, 16, 24) {real, imag} */,
  {32'hbe83bbb2, 32'hbfb85786} /* (15, 16, 23) {real, imag} */,
  {32'h3ef79829, 32'hbf2b6352} /* (15, 16, 22) {real, imag} */,
  {32'hbea0d540, 32'hbe36fe50} /* (15, 16, 21) {real, imag} */,
  {32'hbe12d4c0, 32'hbf85126a} /* (15, 16, 20) {real, imag} */,
  {32'h3ecdfcbc, 32'hbe437978} /* (15, 16, 19) {real, imag} */,
  {32'h3d94b440, 32'h3ec69640} /* (15, 16, 18) {real, imag} */,
  {32'h3d7ec5f0, 32'h3efaf8d0} /* (15, 16, 17) {real, imag} */,
  {32'h3f621fcc, 32'h3fc1d63c} /* (15, 16, 16) {real, imag} */,
  {32'h3bc10a00, 32'hbc922000} /* (15, 16, 15) {real, imag} */,
  {32'hbf83fc50, 32'hbdf890c0} /* (15, 16, 14) {real, imag} */,
  {32'h3f67a8ba, 32'h3f5ce538} /* (15, 16, 13) {real, imag} */,
  {32'h3fef7d37, 32'h3e5200a8} /* (15, 16, 12) {real, imag} */,
  {32'h3d1bbd20, 32'hbf806bbf} /* (15, 16, 11) {real, imag} */,
  {32'hbdd2a188, 32'hbeacacac} /* (15, 16, 10) {real, imag} */,
  {32'hbe8a5c98, 32'h3f1839b8} /* (15, 16, 9) {real, imag} */,
  {32'hbff4c7b0, 32'hbf0de10c} /* (15, 16, 8) {real, imag} */,
  {32'hbe8dd194, 32'h3f6367b0} /* (15, 16, 7) {real, imag} */,
  {32'h4007ceaa, 32'h3fdcd5aa} /* (15, 16, 6) {real, imag} */,
  {32'hbeb881b8, 32'h3f9667c7} /* (15, 16, 5) {real, imag} */,
  {32'hbf56fcec, 32'h3e8e9960} /* (15, 16, 4) {real, imag} */,
  {32'h3e027b88, 32'hbb7c6000} /* (15, 16, 3) {real, imag} */,
  {32'hbf62e3c2, 32'h4018e392} /* (15, 16, 2) {real, imag} */,
  {32'hbf8f97ba, 32'h3f84dc96} /* (15, 16, 1) {real, imag} */,
  {32'hbe0232bc, 32'hbf4afbb0} /* (15, 16, 0) {real, imag} */,
  {32'hbd2921c0, 32'h3e149060} /* (15, 15, 31) {real, imag} */,
  {32'hbf6e3183, 32'h3ec98d54} /* (15, 15, 30) {real, imag} */,
  {32'hbf01a505, 32'hbcb9c2c0} /* (15, 15, 29) {real, imag} */,
  {32'h3ea16f5e, 32'h3c39bf60} /* (15, 15, 28) {real, imag} */,
  {32'h3e1ef340, 32'h3f41bff3} /* (15, 15, 27) {real, imag} */,
  {32'h3f017bf8, 32'h3eac34d1} /* (15, 15, 26) {real, imag} */,
  {32'h3fa9657a, 32'hbf8ad11e} /* (15, 15, 25) {real, imag} */,
  {32'h3efb8012, 32'hbfc07052} /* (15, 15, 24) {real, imag} */,
  {32'h3e9b9f3e, 32'hbe30f2c0} /* (15, 15, 23) {real, imag} */,
  {32'h3e1c7760, 32'h3f21a73e} /* (15, 15, 22) {real, imag} */,
  {32'h3f486d36, 32'h3e567628} /* (15, 15, 21) {real, imag} */,
  {32'h3ebb9eaa, 32'hbf361a90} /* (15, 15, 20) {real, imag} */,
  {32'h3f9a5404, 32'hbf1b443f} /* (15, 15, 19) {real, imag} */,
  {32'hbf972612, 32'hbd834560} /* (15, 15, 18) {real, imag} */,
  {32'hbff9fdce, 32'h3f4e051a} /* (15, 15, 17) {real, imag} */,
  {32'h3e2a122c, 32'hbdae4008} /* (15, 15, 16) {real, imag} */,
  {32'h3f233a10, 32'hbf5eaa0c} /* (15, 15, 15) {real, imag} */,
  {32'h3f732926, 32'hbe4e3a08} /* (15, 15, 14) {real, imag} */,
  {32'h3ebeaddc, 32'h3d94faf0} /* (15, 15, 13) {real, imag} */,
  {32'hbf54df00, 32'hbee2d03c} /* (15, 15, 12) {real, imag} */,
  {32'hbf70ba94, 32'h3f11a536} /* (15, 15, 11) {real, imag} */,
  {32'h3deb45c0, 32'h3f70b9f4} /* (15, 15, 10) {real, imag} */,
  {32'hbf1cacac, 32'hbf549635} /* (15, 15, 9) {real, imag} */,
  {32'h3eca1d14, 32'hbf89d223} /* (15, 15, 8) {real, imag} */,
  {32'hbea6df18, 32'hbdf8c2e0} /* (15, 15, 7) {real, imag} */,
  {32'hbf19dfc5, 32'hbe979d1c} /* (15, 15, 6) {real, imag} */,
  {32'h3e259a30, 32'h3d573ad0} /* (15, 15, 5) {real, imag} */,
  {32'hbfc5cdeb, 32'h3e1c019c} /* (15, 15, 4) {real, imag} */,
  {32'hbfa71340, 32'hbeb73e4c} /* (15, 15, 3) {real, imag} */,
  {32'h3e32fee8, 32'hbf4f913a} /* (15, 15, 2) {real, imag} */,
  {32'hbe92bf06, 32'hbde7f260} /* (15, 15, 1) {real, imag} */,
  {32'h3f72922e, 32'h3f89ba0a} /* (15, 15, 0) {real, imag} */,
  {32'hbdb9c648, 32'hbf0469ad} /* (15, 14, 31) {real, imag} */,
  {32'hbf4fa73a, 32'h3f474eea} /* (15, 14, 30) {real, imag} */,
  {32'hbe804c0c, 32'h3ff9ff4e} /* (15, 14, 29) {real, imag} */,
  {32'h3e58b92a, 32'h3fc6e8c4} /* (15, 14, 28) {real, imag} */,
  {32'hbd844a20, 32'hbf6cc554} /* (15, 14, 27) {real, imag} */,
  {32'h3f01877c, 32'hc0291e64} /* (15, 14, 26) {real, imag} */,
  {32'h400f71e0, 32'hbf39e4c7} /* (15, 14, 25) {real, imag} */,
  {32'h3fd41f54, 32'hbfc9df0e} /* (15, 14, 24) {real, imag} */,
  {32'hbf93fcd2, 32'hbfca228e} /* (15, 14, 23) {real, imag} */,
  {32'hbe34149c, 32'hbfa80060} /* (15, 14, 22) {real, imag} */,
  {32'h3fb1ddd8, 32'hbfb9a651} /* (15, 14, 21) {real, imag} */,
  {32'h3d8949c8, 32'hbf760f95} /* (15, 14, 20) {real, imag} */,
  {32'h3eca3144, 32'hbef31b30} /* (15, 14, 19) {real, imag} */,
  {32'h3f5346cc, 32'hbc9a5340} /* (15, 14, 18) {real, imag} */,
  {32'h3f8e1ed2, 32'h3f598f10} /* (15, 14, 17) {real, imag} */,
  {32'hbeb506f0, 32'h3f73160c} /* (15, 14, 16) {real, imag} */,
  {32'hbf0cbf3f, 32'hbe519a78} /* (15, 14, 15) {real, imag} */,
  {32'hbe5d6dac, 32'hbf923702} /* (15, 14, 14) {real, imag} */,
  {32'hbf3855bf, 32'hc000860a} /* (15, 14, 13) {real, imag} */,
  {32'hbf603533, 32'hbfa426e2} /* (15, 14, 12) {real, imag} */,
  {32'hbf0f5a74, 32'h3f511110} /* (15, 14, 11) {real, imag} */,
  {32'h3f4b0c08, 32'h3cb896c0} /* (15, 14, 10) {real, imag} */,
  {32'h3fb45846, 32'h3e9517dc} /* (15, 14, 9) {real, imag} */,
  {32'h3f65af8a, 32'hbf91a446} /* (15, 14, 8) {real, imag} */,
  {32'h3f97ea3b, 32'hbefead20} /* (15, 14, 7) {real, imag} */,
  {32'h3f1eb8d7, 32'hbfb6f7ac} /* (15, 14, 6) {real, imag} */,
  {32'h3f5fe41e, 32'hbfa2cac0} /* (15, 14, 5) {real, imag} */,
  {32'h3fa8b982, 32'hbf26a49e} /* (15, 14, 4) {real, imag} */,
  {32'h3fbf065a, 32'h3ee8ce38} /* (15, 14, 3) {real, imag} */,
  {32'h3f5982b6, 32'hbf2f4ad9} /* (15, 14, 2) {real, imag} */,
  {32'h3dddde80, 32'hbefad5ed} /* (15, 14, 1) {real, imag} */,
  {32'hbed02f7c, 32'hbf81ded0} /* (15, 14, 0) {real, imag} */,
  {32'hbf2461ea, 32'hbf4bda3c} /* (15, 13, 31) {real, imag} */,
  {32'hbf7bbb06, 32'h3fef2e92} /* (15, 13, 30) {real, imag} */,
  {32'hbf8d1508, 32'h3ff13264} /* (15, 13, 29) {real, imag} */,
  {32'hbdc9c570, 32'h3fdd27bf} /* (15, 13, 28) {real, imag} */,
  {32'hbf3db602, 32'h3fbe52dc} /* (15, 13, 27) {real, imag} */,
  {32'h3fb7fcea, 32'h3f2ceb86} /* (15, 13, 26) {real, imag} */,
  {32'h3f81ef19, 32'h3f686ba7} /* (15, 13, 25) {real, imag} */,
  {32'h3f925812, 32'h3fdd4d2a} /* (15, 13, 24) {real, imag} */,
  {32'h3edee60c, 32'h3f3162df} /* (15, 13, 23) {real, imag} */,
  {32'h3ec4daa2, 32'hbf336366} /* (15, 13, 22) {real, imag} */,
  {32'hbddf5ab8, 32'hbf8dc51d} /* (15, 13, 21) {real, imag} */,
  {32'hbf3f04f4, 32'hbf7f6a7b} /* (15, 13, 20) {real, imag} */,
  {32'h3b537500, 32'hbe84df96} /* (15, 13, 19) {real, imag} */,
  {32'h3f358ade, 32'hbef136ce} /* (15, 13, 18) {real, imag} */,
  {32'h3ecc169c, 32'hc02fd4f7} /* (15, 13, 17) {real, imag} */,
  {32'h3ed3e244, 32'h3ef55428} /* (15, 13, 16) {real, imag} */,
  {32'h3ed93614, 32'h3f8159ad} /* (15, 13, 15) {real, imag} */,
  {32'hbf6075d9, 32'h3e31ef7c} /* (15, 13, 14) {real, imag} */,
  {32'hbf0add2c, 32'h3fd596c8} /* (15, 13, 13) {real, imag} */,
  {32'h3ff1a21e, 32'h400e6cee} /* (15, 13, 12) {real, imag} */,
  {32'h40420b0a, 32'h3f205f31} /* (15, 13, 11) {real, imag} */,
  {32'h3fc8617c, 32'hbfbfaf37} /* (15, 13, 10) {real, imag} */,
  {32'h4006ecba, 32'h3f3b5a84} /* (15, 13, 9) {real, imag} */,
  {32'h3ed4c804, 32'h3f7cb1bf} /* (15, 13, 8) {real, imag} */,
  {32'h3f4b17af, 32'h3f5a9c48} /* (15, 13, 7) {real, imag} */,
  {32'h3f6ca6e8, 32'hbf87b434} /* (15, 13, 6) {real, imag} */,
  {32'hbf8d0d84, 32'h3f85cee0} /* (15, 13, 5) {real, imag} */,
  {32'hbfc1294b, 32'h3f1f24be} /* (15, 13, 4) {real, imag} */,
  {32'hc027ae62, 32'hbf59045f} /* (15, 13, 3) {real, imag} */,
  {32'hbf7dc69c, 32'hbf154990} /* (15, 13, 2) {real, imag} */,
  {32'hbef6f7c6, 32'hbf57c278} /* (15, 13, 1) {real, imag} */,
  {32'hbfb6b6b6, 32'hbf29436f} /* (15, 13, 0) {real, imag} */,
  {32'h3fa9455e, 32'h3f42b376} /* (15, 12, 31) {real, imag} */,
  {32'h3e24b9a8, 32'h3f858560} /* (15, 12, 30) {real, imag} */,
  {32'h3f074f86, 32'h3e1b4820} /* (15, 12, 29) {real, imag} */,
  {32'h3ef10fb4, 32'h3f1598b0} /* (15, 12, 28) {real, imag} */,
  {32'h3d4c5810, 32'hbf80d412} /* (15, 12, 27) {real, imag} */,
  {32'h3f0bd5cc, 32'h3ed82108} /* (15, 12, 26) {real, imag} */,
  {32'hbfcd4e72, 32'h4037b2e0} /* (15, 12, 25) {real, imag} */,
  {32'hbfdb866e, 32'h40353bb0} /* (15, 12, 24) {real, imag} */,
  {32'hc062ac14, 32'h3fa83eab} /* (15, 12, 23) {real, imag} */,
  {32'hc02b8abc, 32'h3f22e281} /* (15, 12, 22) {real, imag} */,
  {32'h3e586b60, 32'h3fbd5002} /* (15, 12, 21) {real, imag} */,
  {32'h3f2ce89a, 32'h3f1753d9} /* (15, 12, 20) {real, imag} */,
  {32'hbff1116b, 32'hbf5f771c} /* (15, 12, 19) {real, imag} */,
  {32'hbfa05422, 32'h3ed142e4} /* (15, 12, 18) {real, imag} */,
  {32'hbe575820, 32'h3fb1f056} /* (15, 12, 17) {real, imag} */,
  {32'hbefa70b8, 32'h3f2b6ae2} /* (15, 12, 16) {real, imag} */,
  {32'hc000a510, 32'h3ed436d4} /* (15, 12, 15) {real, imag} */,
  {32'hc0462a76, 32'hbf9231f6} /* (15, 12, 14) {real, imag} */,
  {32'hbf2be504, 32'h3ebe0e9a} /* (15, 12, 13) {real, imag} */,
  {32'hc010a6c6, 32'h3fb87e56} /* (15, 12, 12) {real, imag} */,
  {32'hbfb35c81, 32'hbf1c4b04} /* (15, 12, 11) {real, imag} */,
  {32'hbf3d16ea, 32'hbf83c112} /* (15, 12, 10) {real, imag} */,
  {32'hbfca6f3c, 32'hbf1c966a} /* (15, 12, 9) {real, imag} */,
  {32'hbf8c8fca, 32'hbf99548c} /* (15, 12, 8) {real, imag} */,
  {32'hbdfff968, 32'hbf28e6aa} /* (15, 12, 7) {real, imag} */,
  {32'hbf0cddb3, 32'h3fea40a4} /* (15, 12, 6) {real, imag} */,
  {32'h3e29085c, 32'h3fd17891} /* (15, 12, 5) {real, imag} */,
  {32'hbb63c800, 32'h3f29847c} /* (15, 12, 4) {real, imag} */,
  {32'h3f3bef80, 32'hbde3ee70} /* (15, 12, 3) {real, imag} */,
  {32'h3f9cd11a, 32'hbf0e2d66} /* (15, 12, 2) {real, imag} */,
  {32'h4011c598, 32'hc01f4626} /* (15, 12, 1) {real, imag} */,
  {32'h3fc3ce5f, 32'hbde74d4c} /* (15, 12, 0) {real, imag} */,
  {32'hbee9398a, 32'hbf95b987} /* (15, 11, 31) {real, imag} */,
  {32'hbea00e82, 32'h3eb69e66} /* (15, 11, 30) {real, imag} */,
  {32'hbfacd0de, 32'h401d298b} /* (15, 11, 29) {real, imag} */,
  {32'h3f25dc9e, 32'h3f7c7746} /* (15, 11, 28) {real, imag} */,
  {32'h3fb633d4, 32'h401127ac} /* (15, 11, 27) {real, imag} */,
  {32'h3fcf5dfc, 32'h3f334f29} /* (15, 11, 26) {real, imag} */,
  {32'h3ea968c8, 32'hc00d5e55} /* (15, 11, 25) {real, imag} */,
  {32'hc0037087, 32'hc01f34d3} /* (15, 11, 24) {real, imag} */,
  {32'hbf682d50, 32'h3e6b8e88} /* (15, 11, 23) {real, imag} */,
  {32'h3e9856a0, 32'h3f73c136} /* (15, 11, 22) {real, imag} */,
  {32'h3f55ba64, 32'h3f700e0c} /* (15, 11, 21) {real, imag} */,
  {32'hbf6442e2, 32'hbd50cdc0} /* (15, 11, 20) {real, imag} */,
  {32'hbf9e38bc, 32'h3e984dd6} /* (15, 11, 19) {real, imag} */,
  {32'h3fc2cbc2, 32'hbd683310} /* (15, 11, 18) {real, imag} */,
  {32'hbfbb0d55, 32'hbfa635a4} /* (15, 11, 17) {real, imag} */,
  {32'hc01aa0ce, 32'hbf60621e} /* (15, 11, 16) {real, imag} */,
  {32'hbf8603af, 32'h3e090788} /* (15, 11, 15) {real, imag} */,
  {32'h3fa73f2e, 32'hbf96d8fa} /* (15, 11, 14) {real, imag} */,
  {32'h4026fd1e, 32'hbdc00c68} /* (15, 11, 13) {real, imag} */,
  {32'h3f4ce30c, 32'h3eb8870c} /* (15, 11, 12) {real, imag} */,
  {32'h3ed6e7c6, 32'h3fb6bb54} /* (15, 11, 11) {real, imag} */,
  {32'h3fd5f291, 32'h3f827364} /* (15, 11, 10) {real, imag} */,
  {32'h3eef3660, 32'hbf0e0a50} /* (15, 11, 9) {real, imag} */,
  {32'hbe98ecc6, 32'h3ff1adb1} /* (15, 11, 8) {real, imag} */,
  {32'hc0373108, 32'h402cac5c} /* (15, 11, 7) {real, imag} */,
  {32'hbf9ddf9e, 32'hbf0ea4a0} /* (15, 11, 6) {real, imag} */,
  {32'h401c0f43, 32'h3f4316b0} /* (15, 11, 5) {real, imag} */,
  {32'h3fa09724, 32'h3f3e74cc} /* (15, 11, 4) {real, imag} */,
  {32'hbf23f1ce, 32'h3ff70550} /* (15, 11, 3) {real, imag} */,
  {32'h40045981, 32'h3f9c2db5} /* (15, 11, 2) {real, imag} */,
  {32'h4012fd8b, 32'h3fefc642} /* (15, 11, 1) {real, imag} */,
  {32'h3f84727c, 32'h3ece57b4} /* (15, 11, 0) {real, imag} */,
  {32'h3fcec51e, 32'h3f6277fd} /* (15, 10, 31) {real, imag} */,
  {32'hbd8cdba0, 32'h3eb515d8} /* (15, 10, 30) {real, imag} */,
  {32'hc00c761e, 32'h3e850f26} /* (15, 10, 29) {real, imag} */,
  {32'h3c3c1380, 32'hbea85f84} /* (15, 10, 28) {real, imag} */,
  {32'h3eb27024, 32'h40054bcb} /* (15, 10, 27) {real, imag} */,
  {32'hbf468c08, 32'h406b8bc8} /* (15, 10, 26) {real, imag} */,
  {32'hbf916c7a, 32'h3ebe1070} /* (15, 10, 25) {real, imag} */,
  {32'hc035c158, 32'h3fe52e26} /* (15, 10, 24) {real, imag} */,
  {32'hc09808ac, 32'h400ed8fb} /* (15, 10, 23) {real, imag} */,
  {32'h3f468b38, 32'hbf9a5ca5} /* (15, 10, 22) {real, imag} */,
  {32'h403d05aa, 32'hbf2488d0} /* (15, 10, 21) {real, imag} */,
  {32'hbf2891c2, 32'hbf84b00d} /* (15, 10, 20) {real, imag} */,
  {32'hc03e9396, 32'hc01ffb10} /* (15, 10, 19) {real, imag} */,
  {32'h3f0ca939, 32'hc0790c4d} /* (15, 10, 18) {real, imag} */,
  {32'h3ed7c7f1, 32'hbe6328d0} /* (15, 10, 17) {real, imag} */,
  {32'hbea92e2c, 32'h4038e2bc} /* (15, 10, 16) {real, imag} */,
  {32'h3fcac17d, 32'hbf32335c} /* (15, 10, 15) {real, imag} */,
  {32'h400097d4, 32'hc00701db} /* (15, 10, 14) {real, imag} */,
  {32'hbcdf8840, 32'hbe61c2b8} /* (15, 10, 13) {real, imag} */,
  {32'hbe93b5a0, 32'hbf86f9b0} /* (15, 10, 12) {real, imag} */,
  {32'hbfb416be, 32'h3eba1374} /* (15, 10, 11) {real, imag} */,
  {32'hbf9c3a81, 32'hbed8e2ae} /* (15, 10, 10) {real, imag} */,
  {32'hc02a7e5f, 32'hbf9f598f} /* (15, 10, 9) {real, imag} */,
  {32'h3f02f064, 32'h3ef02d98} /* (15, 10, 8) {real, imag} */,
  {32'hbcdb4b00, 32'h3f98852e} /* (15, 10, 7) {real, imag} */,
  {32'hbe430008, 32'h3fa85cf7} /* (15, 10, 6) {real, imag} */,
  {32'hbed04f9c, 32'h3e57fd04} /* (15, 10, 5) {real, imag} */,
  {32'hc01709ae, 32'hbff0a2bc} /* (15, 10, 4) {real, imag} */,
  {32'h3f7ff9fa, 32'hbff4fea6} /* (15, 10, 3) {real, imag} */,
  {32'h3f036684, 32'hbf7703d8} /* (15, 10, 2) {real, imag} */,
  {32'hbf471b96, 32'h3f30f4c7} /* (15, 10, 1) {real, imag} */,
  {32'hbeca6dcb, 32'h3f78ab22} /* (15, 10, 0) {real, imag} */,
  {32'h3fd6cb8a, 32'hbff80035} /* (15, 9, 31) {real, imag} */,
  {32'hbf04c9ca, 32'hbf5f3dbf} /* (15, 9, 30) {real, imag} */,
  {32'hbf1d92b2, 32'h3f255e2c} /* (15, 9, 29) {real, imag} */,
  {32'hbfe322cd, 32'h3d8af380} /* (15, 9, 28) {real, imag} */,
  {32'hbf80d7a4, 32'h3fe6a58c} /* (15, 9, 27) {real, imag} */,
  {32'h400941ba, 32'hbf7ebc86} /* (15, 9, 26) {real, imag} */,
  {32'h409009a2, 32'h3f85504b} /* (15, 9, 25) {real, imag} */,
  {32'hc02ea66e, 32'h3fba6fbd} /* (15, 9, 24) {real, imag} */,
  {32'hc082c316, 32'h3dcf06d0} /* (15, 9, 23) {real, imag} */,
  {32'h4043cb24, 32'hbf7aa716} /* (15, 9, 22) {real, imag} */,
  {32'h3f62f9e4, 32'h3fcbdaee} /* (15, 9, 21) {real, imag} */,
  {32'h3de01fa0, 32'hbf6fb2cc} /* (15, 9, 20) {real, imag} */,
  {32'h3fbcd752, 32'hc08314f4} /* (15, 9, 19) {real, imag} */,
  {32'hbf1eb988, 32'h3dc554b0} /* (15, 9, 18) {real, imag} */,
  {32'hc01d53d6, 32'hc0157e98} /* (15, 9, 17) {real, imag} */,
  {32'hbfaeeb6e, 32'hc048c8b3} /* (15, 9, 16) {real, imag} */,
  {32'hbf09fbf4, 32'hbf938b06} /* (15, 9, 15) {real, imag} */,
  {32'h3fbbb14e, 32'hbf490ffd} /* (15, 9, 14) {real, imag} */,
  {32'h4024ba33, 32'hc00bc75c} /* (15, 9, 13) {real, imag} */,
  {32'hc03c74c6, 32'h3f1274cb} /* (15, 9, 12) {real, imag} */,
  {32'hc06a62a8, 32'h408063b7} /* (15, 9, 11) {real, imag} */,
  {32'h4040c9be, 32'h3fc1ecae} /* (15, 9, 10) {real, imag} */,
  {32'h3fc72d21, 32'hc03312e8} /* (15, 9, 9) {real, imag} */,
  {32'hc09ce176, 32'hbfb38af2} /* (15, 9, 8) {real, imag} */,
  {32'h3d9c5f40, 32'h3fe345a4} /* (15, 9, 7) {real, imag} */,
  {32'h401997a5, 32'h3f8af1dc} /* (15, 9, 6) {real, imag} */,
  {32'hbede7f34, 32'h409af21f} /* (15, 9, 5) {real, imag} */,
  {32'h3f8c409d, 32'h407f7990} /* (15, 9, 4) {real, imag} */,
  {32'h3fef565b, 32'h3ecd5b5c} /* (15, 9, 3) {real, imag} */,
  {32'h3f087d10, 32'hbf23afcc} /* (15, 9, 2) {real, imag} */,
  {32'h40408bf6, 32'h3dc38850} /* (15, 9, 1) {real, imag} */,
  {32'h3fc5db50, 32'h3de924a0} /* (15, 9, 0) {real, imag} */,
  {32'hbff6a385, 32'h3ee759bc} /* (15, 8, 31) {real, imag} */,
  {32'hc036bad0, 32'hbfff8c4e} /* (15, 8, 30) {real, imag} */,
  {32'hc0b9b3ea, 32'hbf0a882e} /* (15, 8, 29) {real, imag} */,
  {32'hc0ac274a, 32'h3e9e5f04} /* (15, 8, 28) {real, imag} */,
  {32'hbef5bbf6, 32'hbfa89096} /* (15, 8, 27) {real, imag} */,
  {32'h3fef446e, 32'h40c1c7f2} /* (15, 8, 26) {real, imag} */,
  {32'hbf3fa50e, 32'h40b60f4a} /* (15, 8, 25) {real, imag} */,
  {32'hc028f919, 32'h402f724f} /* (15, 8, 24) {real, imag} */,
  {32'h3e8d6cec, 32'hbf1c739f} /* (15, 8, 23) {real, imag} */,
  {32'h3cb15580, 32'h3eae190e} /* (15, 8, 22) {real, imag} */,
  {32'hc01dae40, 32'h3fb36e9c} /* (15, 8, 21) {real, imag} */,
  {32'hbfce8eb6, 32'hbf1f7df4} /* (15, 8, 20) {real, imag} */,
  {32'h3eb81c2c, 32'h3fbd6e85} /* (15, 8, 19) {real, imag} */,
  {32'h405a36ec, 32'h4007625a} /* (15, 8, 18) {real, imag} */,
  {32'h3fde17d2, 32'hbf9f4804} /* (15, 8, 17) {real, imag} */,
  {32'h40590825, 32'h3f14510c} /* (15, 8, 16) {real, imag} */,
  {32'hbfedec5d, 32'h3ee95a42} /* (15, 8, 15) {real, imag} */,
  {32'hc0d819f8, 32'hbef76d92} /* (15, 8, 14) {real, imag} */,
  {32'hc09846aa, 32'h3f5d26fc} /* (15, 8, 13) {real, imag} */,
  {32'h3f503e34, 32'hbf6c50f6} /* (15, 8, 12) {real, imag} */,
  {32'h3ea44006, 32'hbfe9a8d1} /* (15, 8, 11) {real, imag} */,
  {32'h3d367e50, 32'h3f54db9c} /* (15, 8, 10) {real, imag} */,
  {32'h3d189e00, 32'hc00afc48} /* (15, 8, 9) {real, imag} */,
  {32'h3fbaf0f9, 32'hbe160acc} /* (15, 8, 8) {real, imag} */,
  {32'h403309f6, 32'hbef66b48} /* (15, 8, 7) {real, imag} */,
  {32'h3f141411, 32'hbfa282d0} /* (15, 8, 6) {real, imag} */,
  {32'hc0d59496, 32'hc00645e2} /* (15, 8, 5) {real, imag} */,
  {32'hc0f7aea0, 32'hbfcdc95e} /* (15, 8, 4) {real, imag} */,
  {32'hbfe40a3f, 32'hbf12e90c} /* (15, 8, 3) {real, imag} */,
  {32'h3eede3d4, 32'hc00f200f} /* (15, 8, 2) {real, imag} */,
  {32'hbf237d79, 32'hc04d3236} /* (15, 8, 1) {real, imag} */,
  {32'h3e93f996, 32'h3fae3386} /* (15, 8, 0) {real, imag} */,
  {32'h3f192575, 32'h3c05b140} /* (15, 7, 31) {real, imag} */,
  {32'h4069471e, 32'h3f549dc3} /* (15, 7, 30) {real, imag} */,
  {32'hbf7a5d0c, 32'h4074848f} /* (15, 7, 29) {real, imag} */,
  {32'hc03c5907, 32'h3f04c88b} /* (15, 7, 28) {real, imag} */,
  {32'hbf6a9a36, 32'h405a2a0e} /* (15, 7, 27) {real, imag} */,
  {32'hbf8c5ec4, 32'h403dea30} /* (15, 7, 26) {real, imag} */,
  {32'hbf056eb8, 32'hc051ee0e} /* (15, 7, 25) {real, imag} */,
  {32'hbfc93b28, 32'hc04847ca} /* (15, 7, 24) {real, imag} */,
  {32'hc07b2fb2, 32'hc032f59d} /* (15, 7, 23) {real, imag} */,
  {32'hc0ba2acc, 32'hc04fd2cc} /* (15, 7, 22) {real, imag} */,
  {32'hc0207622, 32'hc01140a8} /* (15, 7, 21) {real, imag} */,
  {32'h3f491ce2, 32'h3f853aac} /* (15, 7, 20) {real, imag} */,
  {32'h404a65c6, 32'hc02c72a8} /* (15, 7, 19) {real, imag} */,
  {32'h40cdca1c, 32'hbf94fcbe} /* (15, 7, 18) {real, imag} */,
  {32'h40b2527a, 32'hbf3dc838} /* (15, 7, 17) {real, imag} */,
  {32'hc01bfead, 32'hc022de14} /* (15, 7, 16) {real, imag} */,
  {32'hbfcb231a, 32'h3f0f1dee} /* (15, 7, 15) {real, imag} */,
  {32'h4056cec1, 32'h3f4c15c3} /* (15, 7, 14) {real, imag} */,
  {32'h408ffb28, 32'hc0582141} /* (15, 7, 13) {real, imag} */,
  {32'h3f6e1cfa, 32'h3e1316b0} /* (15, 7, 12) {real, imag} */,
  {32'hc001bca2, 32'hbd35c780} /* (15, 7, 11) {real, imag} */,
  {32'hbf90e46d, 32'hbff0d136} /* (15, 7, 10) {real, imag} */,
  {32'hbffe7d39, 32'hbfda1ea7} /* (15, 7, 9) {real, imag} */,
  {32'h3fb6e436, 32'hbebb36f4} /* (15, 7, 8) {real, imag} */,
  {32'h3ef7f460, 32'h3ff473d4} /* (15, 7, 7) {real, imag} */,
  {32'hc065711a, 32'hbdede720} /* (15, 7, 6) {real, imag} */,
  {32'hc0b10ae1, 32'h4057409b} /* (15, 7, 5) {real, imag} */,
  {32'hc00255cd, 32'h40b5c258} /* (15, 7, 4) {real, imag} */,
  {32'h4070e4bc, 32'h408828d2} /* (15, 7, 3) {real, imag} */,
  {32'h401d40b7, 32'h40db89ad} /* (15, 7, 2) {real, imag} */,
  {32'h3fa11580, 32'h40ce26a4} /* (15, 7, 1) {real, imag} */,
  {32'h3fd5854e, 32'h402d83fa} /* (15, 7, 0) {real, imag} */,
  {32'hbf3af3d1, 32'h40768bb4} /* (15, 6, 31) {real, imag} */,
  {32'h3f050d84, 32'h40392c1c} /* (15, 6, 30) {real, imag} */,
  {32'hc030e07c, 32'hbf1ef2cf} /* (15, 6, 29) {real, imag} */,
  {32'hc10a36d3, 32'hc03744c6} /* (15, 6, 28) {real, imag} */,
  {32'hc0d91c51, 32'hbf5c9045} /* (15, 6, 27) {real, imag} */,
  {32'h3f97061a, 32'h40720308} /* (15, 6, 26) {real, imag} */,
  {32'h3ec224ce, 32'hbe66c5e8} /* (15, 6, 25) {real, imag} */,
  {32'hbe8a0a38, 32'hc001bf6a} /* (15, 6, 24) {real, imag} */,
  {32'h409b532e, 32'h4002391e} /* (15, 6, 23) {real, imag} */,
  {32'h403694aa, 32'hbf0fc4a6} /* (15, 6, 22) {real, imag} */,
  {32'hbf9d180b, 32'hc0848158} /* (15, 6, 21) {real, imag} */,
  {32'hc02ac17e, 32'hbff94442} /* (15, 6, 20) {real, imag} */,
  {32'h3fa20879, 32'h405a7362} /* (15, 6, 19) {real, imag} */,
  {32'h40384287, 32'hbf51e55c} /* (15, 6, 18) {real, imag} */,
  {32'h3ff47789, 32'hc0828f8d} /* (15, 6, 17) {real, imag} */,
  {32'h3f9556f1, 32'h3f8d4df0} /* (15, 6, 16) {real, imag} */,
  {32'h3f953be1, 32'h40a041cb} /* (15, 6, 15) {real, imag} */,
  {32'hbf0d04d2, 32'hbfea4334} /* (15, 6, 14) {real, imag} */,
  {32'hc094d251, 32'hc06dc86e} /* (15, 6, 13) {real, imag} */,
  {32'hbe8e99d0, 32'hc072fb27} /* (15, 6, 12) {real, imag} */,
  {32'hbf26f164, 32'hc02584da} /* (15, 6, 11) {real, imag} */,
  {32'h3f979432, 32'h40410422} /* (15, 6, 10) {real, imag} */,
  {32'h3fa2bcdf, 32'h3ffde740} /* (15, 6, 9) {real, imag} */,
  {32'hc0eef570, 32'hc07ef9f8} /* (15, 6, 8) {real, imag} */,
  {32'hbfd57546, 32'hc05b1156} /* (15, 6, 7) {real, imag} */,
  {32'h3ed9f7dc, 32'h3f98a53a} /* (15, 6, 6) {real, imag} */,
  {32'h3f7ebf58, 32'h3f0201a2} /* (15, 6, 5) {real, imag} */,
  {32'hc07c96c8, 32'h3fc470a2} /* (15, 6, 4) {real, imag} */,
  {32'hc029984d, 32'h40b0735c} /* (15, 6, 3) {real, imag} */,
  {32'h3f32b3b8, 32'h3ea46940} /* (15, 6, 2) {real, imag} */,
  {32'h3f86dd95, 32'hc05d4f2a} /* (15, 6, 1) {real, imag} */,
  {32'h3fe21366, 32'h3dc930a0} /* (15, 6, 0) {real, imag} */,
  {32'h405981d4, 32'h40127b3f} /* (15, 5, 31) {real, imag} */,
  {32'h3f9095cd, 32'h403fe7e6} /* (15, 5, 30) {real, imag} */,
  {32'hbe5cb1d6, 32'h400caaca} /* (15, 5, 29) {real, imag} */,
  {32'hbfc00a05, 32'hc0cb4e74} /* (15, 5, 28) {real, imag} */,
  {32'hbdf20ac0, 32'hc0d9b5f1} /* (15, 5, 27) {real, imag} */,
  {32'h4096bdb4, 32'hc0825c3e} /* (15, 5, 26) {real, imag} */,
  {32'h40658f95, 32'hbfd38362} /* (15, 5, 25) {real, imag} */,
  {32'h4006ab34, 32'hbf1b6470} /* (15, 5, 24) {real, imag} */,
  {32'h40032f07, 32'hc041fc2a} /* (15, 5, 23) {real, imag} */,
  {32'hc030425a, 32'hbf92a6e0} /* (15, 5, 22) {real, imag} */,
  {32'hc00d2f31, 32'hc0043338} /* (15, 5, 21) {real, imag} */,
  {32'hc02b25fe, 32'hbfa9939a} /* (15, 5, 20) {real, imag} */,
  {32'hbf5b42b0, 32'h3fca6752} /* (15, 5, 19) {real, imag} */,
  {32'hc09fefab, 32'h3ffea559} /* (15, 5, 18) {real, imag} */,
  {32'hc0380f8a, 32'hbfef2094} /* (15, 5, 17) {real, imag} */,
  {32'h3b9e5c00, 32'hc08cb3f4} /* (15, 5, 16) {real, imag} */,
  {32'h40320bdc, 32'hc004fd7e} /* (15, 5, 15) {real, imag} */,
  {32'h3f93608c, 32'h3f910ac2} /* (15, 5, 14) {real, imag} */,
  {32'hc0d5d119, 32'h3fe96311} /* (15, 5, 13) {real, imag} */,
  {32'hc08d59de, 32'h402ab7aa} /* (15, 5, 12) {real, imag} */,
  {32'h3ec47e5c, 32'h403a9245} /* (15, 5, 11) {real, imag} */,
  {32'h40363fc2, 32'h408a2fc2} /* (15, 5, 10) {real, imag} */,
  {32'h40ca8f7c, 32'h4031cf4e} /* (15, 5, 9) {real, imag} */,
  {32'h402135a6, 32'hc0901e50} /* (15, 5, 8) {real, imag} */,
  {32'hc08a59cf, 32'hc1158990} /* (15, 5, 7) {real, imag} */,
  {32'h3c199600, 32'hc0ce1983} /* (15, 5, 6) {real, imag} */,
  {32'h402a936f, 32'hc0935e9b} /* (15, 5, 5) {real, imag} */,
  {32'h3f8e8329, 32'hbf672f0f} /* (15, 5, 4) {real, imag} */,
  {32'hbf95cdc1, 32'h3ff1f6ce} /* (15, 5, 3) {real, imag} */,
  {32'h3fb6a83c, 32'h3f32700d} /* (15, 5, 2) {real, imag} */,
  {32'h4111a54a, 32'h3ee93e20} /* (15, 5, 1) {real, imag} */,
  {32'h40e31082, 32'h40128246} /* (15, 5, 0) {real, imag} */,
  {32'hbfcc9198, 32'h3fa839ed} /* (15, 4, 31) {real, imag} */,
  {32'hc03ca732, 32'hbf47d370} /* (15, 4, 30) {real, imag} */,
  {32'hc0f5678c, 32'hc0301c72} /* (15, 4, 29) {real, imag} */,
  {32'hc12bebc0, 32'h405b64bf} /* (15, 4, 28) {real, imag} */,
  {32'hc0ffbe84, 32'h4090c6b8} /* (15, 4, 27) {real, imag} */,
  {32'hc0f9a70d, 32'h3fcbb321} /* (15, 4, 26) {real, imag} */,
  {32'hc0d0f4d6, 32'h3f8b8a53} /* (15, 4, 25) {real, imag} */,
  {32'h3ec1e784, 32'hbe12f928} /* (15, 4, 24) {real, imag} */,
  {32'h402ae51e, 32'h3eb71be4} /* (15, 4, 23) {real, imag} */,
  {32'hc0aca864, 32'h3fc6fe0b} /* (15, 4, 22) {real, imag} */,
  {32'hbf5c37e0, 32'hbf80f4ca} /* (15, 4, 21) {real, imag} */,
  {32'hc0b09bcc, 32'hc09fb2dd} /* (15, 4, 20) {real, imag} */,
  {32'hc086bfc0, 32'hbed74b30} /* (15, 4, 19) {real, imag} */,
  {32'hbee4e368, 32'h4103ea42} /* (15, 4, 18) {real, imag} */,
  {32'hc0adb24f, 32'h3da63a00} /* (15, 4, 17) {real, imag} */,
  {32'hc0b04dde, 32'hbf106504} /* (15, 4, 16) {real, imag} */,
  {32'h4001a0fd, 32'hbe972cd0} /* (15, 4, 15) {real, imag} */,
  {32'h40092ec6, 32'h3f62f8ce} /* (15, 4, 14) {real, imag} */,
  {32'hbe910238, 32'h4078f57b} /* (15, 4, 13) {real, imag} */,
  {32'hbfc74b5e, 32'h3f4e31d0} /* (15, 4, 12) {real, imag} */,
  {32'hc10410ac, 32'hc0c8baf7} /* (15, 4, 11) {real, imag} */,
  {32'hc03f8a7a, 32'hc06fdcc6} /* (15, 4, 10) {real, imag} */,
  {32'hc043a3fc, 32'h4027c865} /* (15, 4, 9) {real, imag} */,
  {32'h3dbfd870, 32'h40925ad4} /* (15, 4, 8) {real, imag} */,
  {32'h4069d016, 32'h3f4bdf45} /* (15, 4, 7) {real, imag} */,
  {32'h40a062e0, 32'h3dc7b440} /* (15, 4, 6) {real, imag} */,
  {32'h40b20bd6, 32'hbfa128ae} /* (15, 4, 5) {real, imag} */,
  {32'h407996a0, 32'hbf08ffbc} /* (15, 4, 4) {real, imag} */,
  {32'hbf52fbd0, 32'h40a6412c} /* (15, 4, 3) {real, imag} */,
  {32'h3f4f6ba3, 32'h400ae050} /* (15, 4, 2) {real, imag} */,
  {32'hbed620a8, 32'hc068e8c6} /* (15, 4, 1) {real, imag} */,
  {32'h3ede6c10, 32'hc02015a5} /* (15, 4, 0) {real, imag} */,
  {32'h406a8a31, 32'hc04c744c} /* (15, 3, 31) {real, imag} */,
  {32'h3fa8232c, 32'hbff7b59a} /* (15, 3, 30) {real, imag} */,
  {32'hbf86b9cf, 32'hc00f9fe9} /* (15, 3, 29) {real, imag} */,
  {32'h40882e98, 32'hbf997940} /* (15, 3, 28) {real, imag} */,
  {32'h40392b1e, 32'h3f7c135e} /* (15, 3, 27) {real, imag} */,
  {32'h3f984d58, 32'h3ce0c700} /* (15, 3, 26) {real, imag} */,
  {32'h405924ca, 32'h40bd82e6} /* (15, 3, 25) {real, imag} */,
  {32'h3e3b2450, 32'hbede28ac} /* (15, 3, 24) {real, imag} */,
  {32'hc0fe8abe, 32'hbf4bb85f} /* (15, 3, 23) {real, imag} */,
  {32'hc0519e95, 32'h40169ffe} /* (15, 3, 22) {real, imag} */,
  {32'hc04af965, 32'h3fd9eba5} /* (15, 3, 21) {real, imag} */,
  {32'hbfa39d54, 32'h3f7619aa} /* (15, 3, 20) {real, imag} */,
  {32'h40184158, 32'hbf88535f} /* (15, 3, 19) {real, imag} */,
  {32'hc0ba62f4, 32'h3f7fbad4} /* (15, 3, 18) {real, imag} */,
  {32'hc106bc2c, 32'hbe20f5f0} /* (15, 3, 17) {real, imag} */,
  {32'hc0a0e8b3, 32'hbff4ceea} /* (15, 3, 16) {real, imag} */,
  {32'hc086a83d, 32'h3eb0266c} /* (15, 3, 15) {real, imag} */,
  {32'hc0b3ca90, 32'hc02debac} /* (15, 3, 14) {real, imag} */,
  {32'hc009bf41, 32'hbfca59ba} /* (15, 3, 13) {real, imag} */,
  {32'hc001869c, 32'hbf744f50} /* (15, 3, 12) {real, imag} */,
  {32'h3fbc7ea4, 32'hc0030070} /* (15, 3, 11) {real, imag} */,
  {32'hbfd45152, 32'h40812732} /* (15, 3, 10) {real, imag} */,
  {32'h3fae1fa5, 32'h40a9440f} /* (15, 3, 9) {real, imag} */,
  {32'hbe712490, 32'hbfefb02c} /* (15, 3, 8) {real, imag} */,
  {32'h4067af5a, 32'hc003436d} /* (15, 3, 7) {real, imag} */,
  {32'h408c03e6, 32'h411e4f12} /* (15, 3, 6) {real, imag} */,
  {32'hbf6bf994, 32'h40824545} /* (15, 3, 5) {real, imag} */,
  {32'hc0b545c0, 32'h3f969828} /* (15, 3, 4) {real, imag} */,
  {32'hc11c9d21, 32'h403d8103} /* (15, 3, 3) {real, imag} */,
  {32'hc04884a1, 32'hbf5525c0} /* (15, 3, 2) {real, imag} */,
  {32'h3f198ea7, 32'h39544000} /* (15, 3, 1) {real, imag} */,
  {32'h3f5990d4, 32'h3ff1dbb4} /* (15, 3, 0) {real, imag} */,
  {32'hc07433bb, 32'h405a4a52} /* (15, 2, 31) {real, imag} */,
  {32'hc0d79ac4, 32'h40781171} /* (15, 2, 30) {real, imag} */,
  {32'hc051fc3a, 32'h3fac09aa} /* (15, 2, 29) {real, imag} */,
  {32'h4042880d, 32'hbeedbaa0} /* (15, 2, 28) {real, imag} */,
  {32'h40244cef, 32'h4049f53d} /* (15, 2, 27) {real, imag} */,
  {32'hc072c18c, 32'hc07276ee} /* (15, 2, 26) {real, imag} */,
  {32'hc08ca429, 32'h3fd53ab2} /* (15, 2, 25) {real, imag} */,
  {32'hc00766dc, 32'hbf434aa4} /* (15, 2, 24) {real, imag} */,
  {32'h3fac5eff, 32'h4008cdc4} /* (15, 2, 23) {real, imag} */,
  {32'h3f5cb1db, 32'h41151f42} /* (15, 2, 22) {real, imag} */,
  {32'hbf92a714, 32'h408c301e} /* (15, 2, 21) {real, imag} */,
  {32'h3ff305d3, 32'h40eee0e5} /* (15, 2, 20) {real, imag} */,
  {32'h40929904, 32'h41479604} /* (15, 2, 19) {real, imag} */,
  {32'h402091a5, 32'h40cb3681} /* (15, 2, 18) {real, imag} */,
  {32'h4066e5d4, 32'h40363dfa} /* (15, 2, 17) {real, imag} */,
  {32'h3f1cc780, 32'hbe9dbce8} /* (15, 2, 16) {real, imag} */,
  {32'hbd5dcf00, 32'h3e0d41a0} /* (15, 2, 15) {real, imag} */,
  {32'h404f76ab, 32'hc00a5eda} /* (15, 2, 14) {real, imag} */,
  {32'h409ca551, 32'hbe93aca0} /* (15, 2, 13) {real, imag} */,
  {32'h409fd23c, 32'h3dae0f08} /* (15, 2, 12) {real, imag} */,
  {32'h3f8d2b5b, 32'h3f2d7998} /* (15, 2, 11) {real, imag} */,
  {32'hc00c32b8, 32'h40a1a6b4} /* (15, 2, 10) {real, imag} */,
  {32'hc0af581f, 32'h40971c1e} /* (15, 2, 9) {real, imag} */,
  {32'h3e2726ae, 32'h407fb0ad} /* (15, 2, 8) {real, imag} */,
  {32'h40cb01a4, 32'h4046091a} /* (15, 2, 7) {real, imag} */,
  {32'h41314660, 32'h3ffaeab2} /* (15, 2, 6) {real, imag} */,
  {32'hbf22b2c6, 32'h409d2842} /* (15, 2, 5) {real, imag} */,
  {32'hc1098f8c, 32'h4006982b} /* (15, 2, 4) {real, imag} */,
  {32'hc029be7d, 32'hc0616bc9} /* (15, 2, 3) {real, imag} */,
  {32'h4068f356, 32'hc0228c4d} /* (15, 2, 2) {real, imag} */,
  {32'hbed53280, 32'h3e9da236} /* (15, 2, 1) {real, imag} */,
  {32'hc055d10c, 32'hbfd585d2} /* (15, 2, 0) {real, imag} */,
  {32'h3f9a032e, 32'h40a0c161} /* (15, 1, 31) {real, imag} */,
  {32'h3fe788ca, 32'hbe6bd6d0} /* (15, 1, 30) {real, imag} */,
  {32'h4099584d, 32'h4013e274} /* (15, 1, 29) {real, imag} */,
  {32'h3c10e740, 32'h403b0f80} /* (15, 1, 28) {real, imag} */,
  {32'hbf95d45a, 32'h3fa6ce18} /* (15, 1, 27) {real, imag} */,
  {32'h3fc0af44, 32'hbf05684e} /* (15, 1, 26) {real, imag} */,
  {32'h40e2c20c, 32'hbd7e4000} /* (15, 1, 25) {real, imag} */,
  {32'h40961ba2, 32'h40036816} /* (15, 1, 24) {real, imag} */,
  {32'h40a4282c, 32'h3f885d2d} /* (15, 1, 23) {real, imag} */,
  {32'h40d4fd58, 32'hc0367412} /* (15, 1, 22) {real, imag} */,
  {32'h4049a3d8, 32'hbfe4c358} /* (15, 1, 21) {real, imag} */,
  {32'hc0aa3a01, 32'hc06256ac} /* (15, 1, 20) {real, imag} */,
  {32'hc0733ce9, 32'hbfce96b0} /* (15, 1, 19) {real, imag} */,
  {32'hc068650c, 32'h406389d9} /* (15, 1, 18) {real, imag} */,
  {32'h3ef5ce78, 32'h402dd660} /* (15, 1, 17) {real, imag} */,
  {32'hc0f781e4, 32'hc0143dbd} /* (15, 1, 16) {real, imag} */,
  {32'hc106fbbf, 32'hc013a9e4} /* (15, 1, 15) {real, imag} */,
  {32'h3ea4159c, 32'hc041a8a5} /* (15, 1, 14) {real, imag} */,
  {32'hc07ca79b, 32'hbeb26530} /* (15, 1, 13) {real, imag} */,
  {32'hc117ad99, 32'h3e2b1dd0} /* (15, 1, 12) {real, imag} */,
  {32'hc01467d9, 32'h40ac97d1} /* (15, 1, 11) {real, imag} */,
  {32'hbf818a18, 32'h4086b014} /* (15, 1, 10) {real, imag} */,
  {32'h40025238, 32'h400e533e} /* (15, 1, 9) {real, imag} */,
  {32'h4066f728, 32'h405d6837} /* (15, 1, 8) {real, imag} */,
  {32'h40889873, 32'h40a3e4fb} /* (15, 1, 7) {real, imag} */,
  {32'h408abc38, 32'h408af81e} /* (15, 1, 6) {real, imag} */,
  {32'h40cabcae, 32'h3fe66354} /* (15, 1, 5) {real, imag} */,
  {32'h40f20255, 32'h3f74d280} /* (15, 1, 4) {real, imag} */,
  {32'h4113b644, 32'h3ea134a4} /* (15, 1, 3) {real, imag} */,
  {32'h3fc66294, 32'hc0b5eea4} /* (15, 1, 2) {real, imag} */,
  {32'h4043f423, 32'h3fec663c} /* (15, 1, 1) {real, imag} */,
  {32'h40c5feaf, 32'h406fd63c} /* (15, 1, 0) {real, imag} */,
  {32'hc07cbe2f, 32'hc0d7fcfe} /* (15, 0, 31) {real, imag} */,
  {32'hc03020af, 32'hbfafb8fa} /* (15, 0, 30) {real, imag} */,
  {32'h40150b14, 32'h40d7ebd1} /* (15, 0, 29) {real, imag} */,
  {32'h4111c5c0, 32'h40845697} /* (15, 0, 28) {real, imag} */,
  {32'h40029880, 32'h3f9ac18e} /* (15, 0, 27) {real, imag} */,
  {32'hbfb008a7, 32'h3fa41d64} /* (15, 0, 26) {real, imag} */,
  {32'h3f954601, 32'h40dbfc4e} /* (15, 0, 25) {real, imag} */,
  {32'h3f3dc061, 32'hc01a769d} /* (15, 0, 24) {real, imag} */,
  {32'hbfd5120e, 32'hc0e463a2} /* (15, 0, 23) {real, imag} */,
  {32'h3f884994, 32'hbe967bcd} /* (15, 0, 22) {real, imag} */,
  {32'h4093120e, 32'h40104519} /* (15, 0, 21) {real, imag} */,
  {32'h40e61a87, 32'h4076de63} /* (15, 0, 20) {real, imag} */,
  {32'h408c3ed2, 32'hbfd222f9} /* (15, 0, 19) {real, imag} */,
  {32'h3f979550, 32'h410c4cac} /* (15, 0, 18) {real, imag} */,
  {32'hbfd27d80, 32'h4118d0be} /* (15, 0, 17) {real, imag} */,
  {32'h40264907, 32'h40326d5c} /* (15, 0, 16) {real, imag} */,
  {32'h402eed89, 32'h409f5c1e} /* (15, 0, 15) {real, imag} */,
  {32'h40222a68, 32'h40379712} /* (15, 0, 14) {real, imag} */,
  {32'h3ff0c21d, 32'h40a1e7dc} /* (15, 0, 13) {real, imag} */,
  {32'hc0669d88, 32'h3f1c0596} /* (15, 0, 12) {real, imag} */,
  {32'hc021aa68, 32'hbfeaa9c9} /* (15, 0, 11) {real, imag} */,
  {32'hbf7e44a9, 32'hc04db9ac} /* (15, 0, 10) {real, imag} */,
  {32'hc012630c, 32'hc03b93f7} /* (15, 0, 9) {real, imag} */,
  {32'hc08f7d70, 32'hbdea9e40} /* (15, 0, 8) {real, imag} */,
  {32'hc0752d3a, 32'hbf32f214} /* (15, 0, 7) {real, imag} */,
  {32'hbf467b59, 32'h40a47346} /* (15, 0, 6) {real, imag} */,
  {32'h40c1e3ca, 32'h3e5d6e88} /* (15, 0, 5) {real, imag} */,
  {32'h40622251, 32'hc026a102} /* (15, 0, 4) {real, imag} */,
  {32'h3fe1504d, 32'hbf98524c} /* (15, 0, 3) {real, imag} */,
  {32'hbefc18ac, 32'hbf9dd5f6} /* (15, 0, 2) {real, imag} */,
  {32'hc071c0f1, 32'hc0419749} /* (15, 0, 1) {real, imag} */,
  {32'hbfbc054a, 32'hc0761090} /* (15, 0, 0) {real, imag} */,
  {32'hc08c5fa0, 32'hbf549b1a} /* (14, 31, 31) {real, imag} */,
  {32'hc08bae99, 32'hc01cc3fd} /* (14, 31, 30) {real, imag} */,
  {32'hc0a87a8f, 32'hbece17f8} /* (14, 31, 29) {real, imag} */,
  {32'hc14c0ac2, 32'hbf3632fa} /* (14, 31, 28) {real, imag} */,
  {32'hc1449276, 32'h3e88b3a8} /* (14, 31, 27) {real, imag} */,
  {32'hc080cb28, 32'hbe8130ef} /* (14, 31, 26) {real, imag} */,
  {32'hbfff1568, 32'h404ae72e} /* (14, 31, 25) {real, imag} */,
  {32'hc05ba158, 32'h3fcef8a2} /* (14, 31, 24) {real, imag} */,
  {32'hbfb0980c, 32'hbfb2590a} /* (14, 31, 23) {real, imag} */,
  {32'hc0bf26fc, 32'h4046a262} /* (14, 31, 22) {real, imag} */,
  {32'h3f9c24b1, 32'h3fdbbdba} /* (14, 31, 21) {real, imag} */,
  {32'h40cff88e, 32'hc039cddb} /* (14, 31, 20) {real, imag} */,
  {32'h3eeb96ec, 32'h3f54fcd6} /* (14, 31, 19) {real, imag} */,
  {32'h40204ed4, 32'hc0b80500} /* (14, 31, 18) {real, imag} */,
  {32'h405b7434, 32'hc12b1fc2} /* (14, 31, 17) {real, imag} */,
  {32'h408d8947, 32'hc0a2a708} /* (14, 31, 16) {real, imag} */,
  {32'h40cef308, 32'h3fc74409} /* (14, 31, 15) {real, imag} */,
  {32'h41434d46, 32'hc095ce4c} /* (14, 31, 14) {real, imag} */,
  {32'h4076203c, 32'hc0a6d05a} /* (14, 31, 13) {real, imag} */,
  {32'h40b8cd3b, 32'hc091fd1c} /* (14, 31, 12) {real, imag} */,
  {32'h40f27678, 32'hbeab64d8} /* (14, 31, 11) {real, imag} */,
  {32'h40293926, 32'h40c96651} /* (14, 31, 10) {real, imag} */,
  {32'hbf2c01c0, 32'h4102dcf6} /* (14, 31, 9) {real, imag} */,
  {32'hc0822164, 32'h3fe38d7d} /* (14, 31, 8) {real, imag} */,
  {32'hc12e00d6, 32'h40c06649} /* (14, 31, 7) {real, imag} */,
  {32'hc135093b, 32'h410d3821} /* (14, 31, 6) {real, imag} */,
  {32'hc1215c51, 32'h4022e088} /* (14, 31, 5) {real, imag} */,
  {32'hc0ed2760, 32'hc10a24ac} /* (14, 31, 4) {real, imag} */,
  {32'hc08c4d28, 32'hc0654449} /* (14, 31, 3) {real, imag} */,
  {32'hc134afa2, 32'h410b64fc} /* (14, 31, 2) {real, imag} */,
  {32'hc13bfcee, 32'h405f8300} /* (14, 31, 1) {real, imag} */,
  {32'hc0c45a15, 32'hc0892684} /* (14, 31, 0) {real, imag} */,
  {32'h40979d81, 32'hc024eb8a} /* (14, 30, 31) {real, imag} */,
  {32'h405d553c, 32'hc06b1990} /* (14, 30, 30) {real, imag} */,
  {32'h40f7bd56, 32'hc10a23cf} /* (14, 30, 29) {real, imag} */,
  {32'h4024b965, 32'hc0a31a63} /* (14, 30, 28) {real, imag} */,
  {32'h40a01a2a, 32'h4047e1ac} /* (14, 30, 27) {real, imag} */,
  {32'h40eae32b, 32'h40093608} /* (14, 30, 26) {real, imag} */,
  {32'h410c7c08, 32'h407bcd2e} /* (14, 30, 25) {real, imag} */,
  {32'h40ac43d2, 32'hbf43032c} /* (14, 30, 24) {real, imag} */,
  {32'h4101183a, 32'h40692c38} /* (14, 30, 23) {real, imag} */,
  {32'h40db5b4a, 32'h3f4b4560} /* (14, 30, 22) {real, imag} */,
  {32'hbfab867a, 32'hc058e485} /* (14, 30, 21) {real, imag} */,
  {32'hc11711c2, 32'hc02ef2e4} /* (14, 30, 20) {real, imag} */,
  {32'hc1121029, 32'h3dcd3200} /* (14, 30, 19) {real, imag} */,
  {32'hc13a6f4f, 32'h40c0aa68} /* (14, 30, 18) {real, imag} */,
  {32'hc15f3868, 32'h40bea741} /* (14, 30, 17) {real, imag} */,
  {32'hc11571bf, 32'h3fca2ee7} /* (14, 30, 16) {real, imag} */,
  {32'hc1396a8d, 32'h40433bd6} /* (14, 30, 15) {real, imag} */,
  {32'hc0cfad30, 32'h405fe77b} /* (14, 30, 14) {real, imag} */,
  {32'hc0d36ad2, 32'h40415c66} /* (14, 30, 13) {real, imag} */,
  {32'hc1272a1e, 32'h40671dd4} /* (14, 30, 12) {real, imag} */,
  {32'h3ff5c0e4, 32'h3f0820f8} /* (14, 30, 11) {real, imag} */,
  {32'h411d0f88, 32'hc08a423d} /* (14, 30, 10) {real, imag} */,
  {32'h411421e1, 32'h3f9490e4} /* (14, 30, 9) {real, imag} */,
  {32'h40c59304, 32'h4067b1dd} /* (14, 30, 8) {real, imag} */,
  {32'h411fc822, 32'hc05a954c} /* (14, 30, 7) {real, imag} */,
  {32'h410ebe17, 32'hc01c3527} /* (14, 30, 6) {real, imag} */,
  {32'h402f9790, 32'hbf6c7dd1} /* (14, 30, 5) {real, imag} */,
  {32'h4110b3a0, 32'hc0743598} /* (14, 30, 4) {real, imag} */,
  {32'h414fee47, 32'hc01c4d47} /* (14, 30, 3) {real, imag} */,
  {32'h41120ab3, 32'h3fd3e80e} /* (14, 30, 2) {real, imag} */,
  {32'h410c3dbd, 32'h40941bf0} /* (14, 30, 1) {real, imag} */,
  {32'h40a69e3e, 32'h4039368e} /* (14, 30, 0) {real, imag} */,
  {32'hbfe705a0, 32'hbf7c4474} /* (14, 29, 31) {real, imag} */,
  {32'h3ca0bf00, 32'hbfefdcca} /* (14, 29, 30) {real, imag} */,
  {32'hc091cd0f, 32'h401cc722} /* (14, 29, 29) {real, imag} */,
  {32'h3fd47242, 32'h40b4ea60} /* (14, 29, 28) {real, imag} */,
  {32'h40c546b0, 32'h40ed28b9} /* (14, 29, 27) {real, imag} */,
  {32'hc0281d3b, 32'h4081bd98} /* (14, 29, 26) {real, imag} */,
  {32'hc02e18a0, 32'hc023119d} /* (14, 29, 25) {real, imag} */,
  {32'hc103af19, 32'hc0dfce4a} /* (14, 29, 24) {real, imag} */,
  {32'hbfd7b9c8, 32'hc01c6d05} /* (14, 29, 23) {real, imag} */,
  {32'h3f6cb1f0, 32'h4005b1fa} /* (14, 29, 22) {real, imag} */,
  {32'h3fffe660, 32'hbfad8706} /* (14, 29, 21) {real, imag} */,
  {32'hbe3da688, 32'hc0e250fa} /* (14, 29, 20) {real, imag} */,
  {32'hbfd9278d, 32'h3fd4d684} /* (14, 29, 19) {real, imag} */,
  {32'h4007f2ae, 32'h40af4ff6} /* (14, 29, 18) {real, imag} */,
  {32'h408d090b, 32'h4089360b} /* (14, 29, 17) {real, imag} */,
  {32'h40280f66, 32'hbfdb24b9} /* (14, 29, 16) {real, imag} */,
  {32'h4080c3bb, 32'hc08c633a} /* (14, 29, 15) {real, imag} */,
  {32'h4078a63d, 32'h4050ce72} /* (14, 29, 14) {real, imag} */,
  {32'h3f62a3b3, 32'h4091e916} /* (14, 29, 13) {real, imag} */,
  {32'hbe8179d0, 32'h405e91d3} /* (14, 29, 12) {real, imag} */,
  {32'hc09a6d0a, 32'hc11a95e0} /* (14, 29, 11) {real, imag} */,
  {32'hbec1757a, 32'hc0858872} /* (14, 29, 10) {real, imag} */,
  {32'hbf3bf588, 32'h40ae58b0} /* (14, 29, 9) {real, imag} */,
  {32'hc0ec5858, 32'h40f53b41} /* (14, 29, 8) {real, imag} */,
  {32'hc0dd116f, 32'h40a8715d} /* (14, 29, 7) {real, imag} */,
  {32'h3f47eb44, 32'h413d9610} /* (14, 29, 6) {real, imag} */,
  {32'hbf8af950, 32'h40e6a587} /* (14, 29, 5) {real, imag} */,
  {32'hc01702b4, 32'h3fe3d1b0} /* (14, 29, 4) {real, imag} */,
  {32'hc09a44f1, 32'hbfa0a82f} /* (14, 29, 3) {real, imag} */,
  {32'hc04ff43e, 32'hc0387820} /* (14, 29, 2) {real, imag} */,
  {32'hc0ba413e, 32'hbf79704d} /* (14, 29, 1) {real, imag} */,
  {32'hc020b1c6, 32'h3f90fe4d} /* (14, 29, 0) {real, imag} */,
  {32'h405a38f6, 32'h4046d552} /* (14, 28, 31) {real, imag} */,
  {32'hc09b107a, 32'h411931ba} /* (14, 28, 30) {real, imag} */,
  {32'hc13ceb12, 32'h41372f2d} /* (14, 28, 29) {real, imag} */,
  {32'hc0dc5cd5, 32'h410650c7} /* (14, 28, 28) {real, imag} */,
  {32'hc10dd1a4, 32'h4081c4e5} /* (14, 28, 27) {real, imag} */,
  {32'hc0a90eda, 32'hbf89aee3} /* (14, 28, 26) {real, imag} */,
  {32'hbfcd791d, 32'hc0881f8b} /* (14, 28, 25) {real, imag} */,
  {32'hbf970a72, 32'hc071d200} /* (14, 28, 24) {real, imag} */,
  {32'hc09495c2, 32'hbe4ffab8} /* (14, 28, 23) {real, imag} */,
  {32'hc095bf4e, 32'hbf114e54} /* (14, 28, 22) {real, imag} */,
  {32'h3f74f998, 32'h3f6cfa11} /* (14, 28, 21) {real, imag} */,
  {32'h4112a500, 32'hc05bc9d3} /* (14, 28, 20) {real, imag} */,
  {32'h4141609c, 32'hc12e4e90} /* (14, 28, 19) {real, imag} */,
  {32'hc07b2c7a, 32'hc0f020b3} /* (14, 28, 18) {real, imag} */,
  {32'hc07b62e3, 32'hc1166eb7} /* (14, 28, 17) {real, imag} */,
  {32'h4048f380, 32'hc12908f7} /* (14, 28, 16) {real, imag} */,
  {32'h404308ea, 32'h4066011c} /* (14, 28, 15) {real, imag} */,
  {32'hc06cd05f, 32'h40baf944} /* (14, 28, 14) {real, imag} */,
  {32'h3ef5bf90, 32'h3d9435d0} /* (14, 28, 13) {real, imag} */,
  {32'h40fb1254, 32'hc0e24207} /* (14, 28, 12) {real, imag} */,
  {32'h4116763c, 32'hc0d685f3} /* (14, 28, 11) {real, imag} */,
  {32'hbe0b6578, 32'hbf399aa8} /* (14, 28, 10) {real, imag} */,
  {32'hc0985371, 32'hbff6a453} /* (14, 28, 9) {real, imag} */,
  {32'hc02b5fcf, 32'hc0493cad} /* (14, 28, 8) {real, imag} */,
  {32'hc0aba1c8, 32'hbfd55588} /* (14, 28, 7) {real, imag} */,
  {32'hc04c0c34, 32'h40823adf} /* (14, 28, 6) {real, imag} */,
  {32'hc0983e56, 32'h3f5de85a} /* (14, 28, 5) {real, imag} */,
  {32'hc0381f22, 32'h3dc18960} /* (14, 28, 4) {real, imag} */,
  {32'h40145c55, 32'h4015449c} /* (14, 28, 3) {real, imag} */,
  {32'h408552d7, 32'h40a40af9} /* (14, 28, 2) {real, imag} */,
  {32'h4037d6aa, 32'hbe3235c0} /* (14, 28, 1) {real, imag} */,
  {32'hbf35bab3, 32'hc00af1fd} /* (14, 28, 0) {real, imag} */,
  {32'h4022a600, 32'h3f62ff55} /* (14, 27, 31) {real, imag} */,
  {32'h3ff97b7a, 32'h3fcfa1f4} /* (14, 27, 30) {real, imag} */,
  {32'hc0da9959, 32'hbf11118d} /* (14, 27, 29) {real, imag} */,
  {32'hc01e3425, 32'hc0e811e2} /* (14, 27, 28) {real, imag} */,
  {32'hc048addb, 32'hc03f0d14} /* (14, 27, 27) {real, imag} */,
  {32'h3f7e2440, 32'h405f3f9e} /* (14, 27, 26) {real, imag} */,
  {32'h4000b4a4, 32'h3f0f71d7} /* (14, 27, 25) {real, imag} */,
  {32'h4093cbee, 32'hc035de87} /* (14, 27, 24) {real, imag} */,
  {32'h404028fc, 32'hc094e990} /* (14, 27, 23) {real, imag} */,
  {32'h3ec13830, 32'hc09ef1c0} /* (14, 27, 22) {real, imag} */,
  {32'hbe7a20d8, 32'hbf0bf548} /* (14, 27, 21) {real, imag} */,
  {32'hbf52811d, 32'h409e45cc} /* (14, 27, 20) {real, imag} */,
  {32'hc08420b1, 32'h4052de88} /* (14, 27, 19) {real, imag} */,
  {32'hc02dfd0a, 32'h40917124} /* (14, 27, 18) {real, imag} */,
  {32'h401a3c08, 32'h3fb55e5e} /* (14, 27, 17) {real, imag} */,
  {32'h405322ba, 32'h4026553c} /* (14, 27, 16) {real, imag} */,
  {32'hbf17f590, 32'h40aabd22} /* (14, 27, 15) {real, imag} */,
  {32'hc0ccd1d2, 32'h40ebae3a} /* (14, 27, 14) {real, imag} */,
  {32'hbfb5fed5, 32'h40729482} /* (14, 27, 13) {real, imag} */,
  {32'hc0460577, 32'h41041d4c} /* (14, 27, 12) {real, imag} */,
  {32'hc0b057a4, 32'h40bf4a87} /* (14, 27, 11) {real, imag} */,
  {32'h4079be28, 32'h4002173e} /* (14, 27, 10) {real, imag} */,
  {32'h4113bf9e, 32'h3fe2c7bc} /* (14, 27, 9) {real, imag} */,
  {32'h3f5e76ff, 32'hc0a6bbf8} /* (14, 27, 8) {real, imag} */,
  {32'h3ff8fd3a, 32'hbf53a80c} /* (14, 27, 7) {real, imag} */,
  {32'h408cd43c, 32'hc01f146b} /* (14, 27, 6) {real, imag} */,
  {32'h40c71147, 32'hbfa73d3c} /* (14, 27, 5) {real, imag} */,
  {32'h4133a74c, 32'h3fbfcc94} /* (14, 27, 4) {real, imag} */,
  {32'h40adf2a6, 32'hbf4e6daf} /* (14, 27, 3) {real, imag} */,
  {32'h406fca95, 32'h4073242a} /* (14, 27, 2) {real, imag} */,
  {32'h408d275f, 32'h41220553} /* (14, 27, 1) {real, imag} */,
  {32'h3fa6c788, 32'h4013c4d0} /* (14, 27, 0) {real, imag} */,
  {32'hbf2b58ac, 32'h405c4498} /* (14, 26, 31) {real, imag} */,
  {32'hbeaad4ac, 32'h40434a1e} /* (14, 26, 30) {real, imag} */,
  {32'h402c56eb, 32'h40610154} /* (14, 26, 29) {real, imag} */,
  {32'h3fbbf3a0, 32'h408b32a2} /* (14, 26, 28) {real, imag} */,
  {32'hbfda9ccd, 32'h3fe69e22} /* (14, 26, 27) {real, imag} */,
  {32'h3c300600, 32'h3fae3e41} /* (14, 26, 26) {real, imag} */,
  {32'hbf8a0a78, 32'h3fa54786} /* (14, 26, 25) {real, imag} */,
  {32'hc01f8907, 32'h3fa35900} /* (14, 26, 24) {real, imag} */,
  {32'hc0594d86, 32'hbf0a796a} /* (14, 26, 23) {real, imag} */,
  {32'h3ea442d0, 32'h40457719} /* (14, 26, 22) {real, imag} */,
  {32'hc07521fa, 32'hbf83f0e5} /* (14, 26, 21) {real, imag} */,
  {32'h3fc78cab, 32'hbfd85f18} /* (14, 26, 20) {real, imag} */,
  {32'h408baee3, 32'hc039fd15} /* (14, 26, 19) {real, imag} */,
  {32'h403f3ad4, 32'hc04d819b} /* (14, 26, 18) {real, imag} */,
  {32'hc005d564, 32'hbe2eb568} /* (14, 26, 17) {real, imag} */,
  {32'hc04630f5, 32'h3fe03017} /* (14, 26, 16) {real, imag} */,
  {32'hc0aa8b74, 32'h3fbfed7a} /* (14, 26, 15) {real, imag} */,
  {32'hc0d3f2bb, 32'h408fc3c4} /* (14, 26, 14) {real, imag} */,
  {32'hbfa2318e, 32'h40573ff2} /* (14, 26, 13) {real, imag} */,
  {32'hc01c4272, 32'h407424d8} /* (14, 26, 12) {real, imag} */,
  {32'hc0e3d65c, 32'h3f659f08} /* (14, 26, 11) {real, imag} */,
  {32'hc0bd3cfe, 32'hc0053b9e} /* (14, 26, 10) {real, imag} */,
  {32'h4022b8f7, 32'hc032366c} /* (14, 26, 9) {real, imag} */,
  {32'h4087360c, 32'h3f989838} /* (14, 26, 8) {real, imag} */,
  {32'hbfb89837, 32'h3fac689f} /* (14, 26, 7) {real, imag} */,
  {32'h3f05b790, 32'hbd840300} /* (14, 26, 6) {real, imag} */,
  {32'hc07683ff, 32'hbfbcc8b4} /* (14, 26, 5) {real, imag} */,
  {32'h3f223ba9, 32'hc0431535} /* (14, 26, 4) {real, imag} */,
  {32'hbfb7f653, 32'h3e6d1994} /* (14, 26, 3) {real, imag} */,
  {32'hc07f8d38, 32'h405da368} /* (14, 26, 2) {real, imag} */,
  {32'hc0325bb1, 32'h406b9697} /* (14, 26, 1) {real, imag} */,
  {32'h3dc6d9f0, 32'h3f8da816} /* (14, 26, 0) {real, imag} */,
  {32'h3e6a55c0, 32'h40aa4d4b} /* (14, 25, 31) {real, imag} */,
  {32'h3f292c80, 32'h40c16afc} /* (14, 25, 30) {real, imag} */,
  {32'h40308dfb, 32'h400df202} /* (14, 25, 29) {real, imag} */,
  {32'hc071922c, 32'hbf1a491e} /* (14, 25, 28) {real, imag} */,
  {32'hc08512ca, 32'hc092b820} /* (14, 25, 27) {real, imag} */,
  {32'hc00d1421, 32'hc0e4be8a} /* (14, 25, 26) {real, imag} */,
  {32'hbda5da10, 32'hc0961c05} /* (14, 25, 25) {real, imag} */,
  {32'hbbf4c480, 32'hc0d0da60} /* (14, 25, 24) {real, imag} */,
  {32'hbfdd03f5, 32'hc0a721b0} /* (14, 25, 23) {real, imag} */,
  {32'hc0923e9a, 32'hbfb99512} /* (14, 25, 22) {real, imag} */,
  {32'hc0ccc87f, 32'h3e1858c0} /* (14, 25, 21) {real, imag} */,
  {32'hc0023710, 32'hbfe8fa88} /* (14, 25, 20) {real, imag} */,
  {32'h400f772d, 32'h3f4705c2} /* (14, 25, 19) {real, imag} */,
  {32'h4069aecd, 32'h40df2f68} /* (14, 25, 18) {real, imag} */,
  {32'h406f738e, 32'h400e167a} /* (14, 25, 17) {real, imag} */,
  {32'h40363d54, 32'hbf9175f6} /* (14, 25, 16) {real, imag} */,
  {32'h3fc4fdb6, 32'hc040f47c} /* (14, 25, 15) {real, imag} */,
  {32'h3f878d4b, 32'hbff69d55} /* (14, 25, 14) {real, imag} */,
  {32'h3ebb4280, 32'h3f15616d} /* (14, 25, 13) {real, imag} */,
  {32'h40a7cad6, 32'h4058a2b3} /* (14, 25, 12) {real, imag} */,
  {32'hbcdc16c0, 32'h3fc3adaf} /* (14, 25, 11) {real, imag} */,
  {32'hbed38c7e, 32'h3d0e0fa0} /* (14, 25, 10) {real, imag} */,
  {32'hc08d9c8a, 32'h3f0f7660} /* (14, 25, 9) {real, imag} */,
  {32'hc0a51034, 32'h3fec7a32} /* (14, 25, 8) {real, imag} */,
  {32'hbf8dded2, 32'h3fdcb494} /* (14, 25, 7) {real, imag} */,
  {32'h3f7d3830, 32'h3f8d2eaa} /* (14, 25, 6) {real, imag} */,
  {32'hbfec650b, 32'h3f999900} /* (14, 25, 5) {real, imag} */,
  {32'hc0369e5c, 32'h4099fa87} /* (14, 25, 4) {real, imag} */,
  {32'h3f991ec0, 32'h40bf619d} /* (14, 25, 3) {real, imag} */,
  {32'h3f1569de, 32'h3fce943e} /* (14, 25, 2) {real, imag} */,
  {32'hbe551a18, 32'h402f5a6c} /* (14, 25, 1) {real, imag} */,
  {32'h3ecd7118, 32'h40b22c78} /* (14, 25, 0) {real, imag} */,
  {32'h40565c44, 32'hc03b5bb4} /* (14, 24, 31) {real, imag} */,
  {32'h402e89a6, 32'h3ef9f210} /* (14, 24, 30) {real, imag} */,
  {32'hc00288ff, 32'hc02061f6} /* (14, 24, 29) {real, imag} */,
  {32'hbf637950, 32'hc0d381c6} /* (14, 24, 28) {real, imag} */,
  {32'h3ea557f4, 32'hc0607883} /* (14, 24, 27) {real, imag} */,
  {32'h3fc599e2, 32'h3f360764} /* (14, 24, 26) {real, imag} */,
  {32'h3fee3bbe, 32'h40266b17} /* (14, 24, 25) {real, imag} */,
  {32'h3fcea4ac, 32'h4051c7b4} /* (14, 24, 24) {real, imag} */,
  {32'h409e1705, 32'h40953677} /* (14, 24, 23) {real, imag} */,
  {32'h402f4c24, 32'h3fab66d1} /* (14, 24, 22) {real, imag} */,
  {32'h3f0812b8, 32'hbfd62803} /* (14, 24, 21) {real, imag} */,
  {32'hbf888507, 32'hbf41920c} /* (14, 24, 20) {real, imag} */,
  {32'hbfd5622f, 32'h3fefa014} /* (14, 24, 19) {real, imag} */,
  {32'h3e818694, 32'h40aab18a} /* (14, 24, 18) {real, imag} */,
  {32'hc080f963, 32'h401f5a7c} /* (14, 24, 17) {real, imag} */,
  {32'hc08b9647, 32'h3f294b68} /* (14, 24, 16) {real, imag} */,
  {32'h3f03960c, 32'h3ded8928} /* (14, 24, 15) {real, imag} */,
  {32'h3e287ed0, 32'h3f174e7c} /* (14, 24, 14) {real, imag} */,
  {32'hc02114e0, 32'h400d1ff1} /* (14, 24, 13) {real, imag} */,
  {32'hbf3d1544, 32'hbff4ac2e} /* (14, 24, 12) {real, imag} */,
  {32'hbfbd5bf9, 32'h40241d34} /* (14, 24, 11) {real, imag} */,
  {32'h3f4b5fa5, 32'h3fb32be0} /* (14, 24, 10) {real, imag} */,
  {32'hc035b004, 32'hc045bf24} /* (14, 24, 9) {real, imag} */,
  {32'h40075c91, 32'hba840c00} /* (14, 24, 8) {real, imag} */,
  {32'h406c3411, 32'hc010214d} /* (14, 24, 7) {real, imag} */,
  {32'h408cc052, 32'hbfef75cd} /* (14, 24, 6) {real, imag} */,
  {32'h40842130, 32'hc080b453} /* (14, 24, 5) {real, imag} */,
  {32'h404e1ab3, 32'h3e91b2a8} /* (14, 24, 4) {real, imag} */,
  {32'h40554227, 32'h40d5ca23} /* (14, 24, 3) {real, imag} */,
  {32'hc025ae21, 32'hbfebbd48} /* (14, 24, 2) {real, imag} */,
  {32'hc0be3878, 32'hc0851583} /* (14, 24, 1) {real, imag} */,
  {32'hc002a22f, 32'hbfdec78c} /* (14, 24, 0) {real, imag} */,
  {32'h3f9138d2, 32'h3fa5fae7} /* (14, 23, 31) {real, imag} */,
  {32'hbf0b57fe, 32'hbfeb08a8} /* (14, 23, 30) {real, imag} */,
  {32'hbf2e2a2c, 32'hbff5ea72} /* (14, 23, 29) {real, imag} */,
  {32'h40aa75b3, 32'h4075cf6e} /* (14, 23, 28) {real, imag} */,
  {32'h406543f8, 32'h403eb48c} /* (14, 23, 27) {real, imag} */,
  {32'hbebd08d8, 32'hbfabd37d} /* (14, 23, 26) {real, imag} */,
  {32'hbc48b780, 32'hbfebc490} /* (14, 23, 25) {real, imag} */,
  {32'h3f1efe14, 32'hc06a385b} /* (14, 23, 24) {real, imag} */,
  {32'h3f93abc3, 32'hc0aa6530} /* (14, 23, 23) {real, imag} */,
  {32'h3ef0db5c, 32'hc080d974} /* (14, 23, 22) {real, imag} */,
  {32'hbfbeed79, 32'h401f48d6} /* (14, 23, 21) {real, imag} */,
  {32'hbfb82de6, 32'h40af7e85} /* (14, 23, 20) {real, imag} */,
  {32'hbfa2e10e, 32'h40a03874} /* (14, 23, 19) {real, imag} */,
  {32'hc06edb5d, 32'h3ffc985e} /* (14, 23, 18) {real, imag} */,
  {32'hc027b4b2, 32'h3eecd224} /* (14, 23, 17) {real, imag} */,
  {32'hbef13128, 32'h3ea3a24e} /* (14, 23, 16) {real, imag} */,
  {32'h3f190258, 32'h3f85cfe6} /* (14, 23, 15) {real, imag} */,
  {32'hbed2ebf4, 32'hbfe761bb} /* (14, 23, 14) {real, imag} */,
  {32'h3ee1d778, 32'hc0621b35} /* (14, 23, 13) {real, imag} */,
  {32'h3f44f574, 32'h3c90bf00} /* (14, 23, 12) {real, imag} */,
  {32'h3fe006a3, 32'h402af8e7} /* (14, 23, 11) {real, imag} */,
  {32'h3fa59c73, 32'h4009bb45} /* (14, 23, 10) {real, imag} */,
  {32'hbdc83620, 32'h40812ad3} /* (14, 23, 9) {real, imag} */,
  {32'hc0294092, 32'h406e0c54} /* (14, 23, 8) {real, imag} */,
  {32'hbf19a084, 32'h3e91f040} /* (14, 23, 7) {real, imag} */,
  {32'h3fa16cec, 32'hc0115a4f} /* (14, 23, 6) {real, imag} */,
  {32'h3fe08334, 32'h3f0a8598} /* (14, 23, 5) {real, imag} */,
  {32'hc02dbdd2, 32'h3ecfb230} /* (14, 23, 4) {real, imag} */,
  {32'hc08f662c, 32'h4006f71a} /* (14, 23, 3) {real, imag} */,
  {32'hc082b11b, 32'h40603383} /* (14, 23, 2) {real, imag} */,
  {32'hc087f980, 32'h40ba3d20} /* (14, 23, 1) {real, imag} */,
  {32'hbe361824, 32'h3ffaf8d5} /* (14, 23, 0) {real, imag} */,
  {32'hc03f910a, 32'h3fbf7b73} /* (14, 22, 31) {real, imag} */,
  {32'h402d4ff2, 32'hbe872194} /* (14, 22, 30) {real, imag} */,
  {32'h408e6406, 32'hbdcae9c0} /* (14, 22, 29) {real, imag} */,
  {32'h40655eb3, 32'hbfe983fc} /* (14, 22, 28) {real, imag} */,
  {32'h4066a9c8, 32'hc031cb88} /* (14, 22, 27) {real, imag} */,
  {32'hbefaa9f8, 32'hbf84bc10} /* (14, 22, 26) {real, imag} */,
  {32'hc039a18f, 32'h3e9b8416} /* (14, 22, 25) {real, imag} */,
  {32'hbf26ee6f, 32'h4043cb94} /* (14, 22, 24) {real, imag} */,
  {32'hc01d7fc3, 32'h3f8f32ef} /* (14, 22, 23) {real, imag} */,
  {32'h3f2fa630, 32'hbe438028} /* (14, 22, 22) {real, imag} */,
  {32'h4022ad9e, 32'hbff295fa} /* (14, 22, 21) {real, imag} */,
  {32'h3fa3d4e6, 32'hbfa2836e} /* (14, 22, 20) {real, imag} */,
  {32'h3fd29e85, 32'h3fe310da} /* (14, 22, 19) {real, imag} */,
  {32'h407ab512, 32'h3d944c70} /* (14, 22, 18) {real, imag} */,
  {32'hbc6eee00, 32'hbf190f22} /* (14, 22, 17) {real, imag} */,
  {32'hbfa773ee, 32'h3f93c99f} /* (14, 22, 16) {real, imag} */,
  {32'hbf0066af, 32'h4002642c} /* (14, 22, 15) {real, imag} */,
  {32'hbfeb3328, 32'hbf14ad10} /* (14, 22, 14) {real, imag} */,
  {32'hbfda65e8, 32'hc04403e1} /* (14, 22, 13) {real, imag} */,
  {32'h3f14eba2, 32'h3ed8cc30} /* (14, 22, 12) {real, imag} */,
  {32'h3f98c626, 32'h3fb46232} /* (14, 22, 11) {real, imag} */,
  {32'hbe491eb8, 32'h3ea79dcc} /* (14, 22, 10) {real, imag} */,
  {32'hc01326ea, 32'h3f8cbc88} /* (14, 22, 9) {real, imag} */,
  {32'hc034e696, 32'h3ea07928} /* (14, 22, 8) {real, imag} */,
  {32'hbd958610, 32'h40367a04} /* (14, 22, 7) {real, imag} */,
  {32'h4018964b, 32'h40e11380} /* (14, 22, 6) {real, imag} */,
  {32'h3fec7c9a, 32'h4099fd78} /* (14, 22, 5) {real, imag} */,
  {32'h3f3924b2, 32'h3ff17eed} /* (14, 22, 4) {real, imag} */,
  {32'h400e7542, 32'h3fbec456} /* (14, 22, 3) {real, imag} */,
  {32'h3fd3d22f, 32'hbff976ac} /* (14, 22, 2) {real, imag} */,
  {32'h3ff3582a, 32'hbfdd04c4} /* (14, 22, 1) {real, imag} */,
  {32'h3ff555ec, 32'h3fd0fb22} /* (14, 22, 0) {real, imag} */,
  {32'h3fa8fc89, 32'h3ff8c1cf} /* (14, 21, 31) {real, imag} */,
  {32'h3f22434a, 32'h40506056} /* (14, 21, 30) {real, imag} */,
  {32'hbebfa400, 32'h3fd0e368} /* (14, 21, 29) {real, imag} */,
  {32'hbfb80c87, 32'hc0139201} /* (14, 21, 28) {real, imag} */,
  {32'hbff4742c, 32'hc02110ee} /* (14, 21, 27) {real, imag} */,
  {32'hbe8282e0, 32'h3e210898} /* (14, 21, 26) {real, imag} */,
  {32'hbfd1053c, 32'hbe13e5d8} /* (14, 21, 25) {real, imag} */,
  {32'hbfc66301, 32'h3f0ccd74} /* (14, 21, 24) {real, imag} */,
  {32'h3e191118, 32'h406dde6c} /* (14, 21, 23) {real, imag} */,
  {32'hc011b208, 32'hbf56d281} /* (14, 21, 22) {real, imag} */,
  {32'hbf50c20a, 32'hc00a661e} /* (14, 21, 21) {real, imag} */,
  {32'hbf8bbe1e, 32'hc062f511} /* (14, 21, 20) {real, imag} */,
  {32'hbf88376e, 32'h3f3e5e48} /* (14, 21, 19) {real, imag} */,
  {32'hbf267b40, 32'hbf07e9e5} /* (14, 21, 18) {real, imag} */,
  {32'h3f10d636, 32'h400128fb} /* (14, 21, 17) {real, imag} */,
  {32'hbefc943a, 32'h3f9e3243} /* (14, 21, 16) {real, imag} */,
  {32'hc095a456, 32'hc052fdfc} /* (14, 21, 15) {real, imag} */,
  {32'hc0853bfe, 32'hbf6e3918} /* (14, 21, 14) {real, imag} */,
  {32'hbfe8e16f, 32'hc0a673fd} /* (14, 21, 13) {real, imag} */,
  {32'h3d013508, 32'hc0a8b393} /* (14, 21, 12) {real, imag} */,
  {32'hbea498ba, 32'h3c049b80} /* (14, 21, 11) {real, imag} */,
  {32'h3e3eb694, 32'h3e8c1fce} /* (14, 21, 10) {real, imag} */,
  {32'h3ed1cafc, 32'hbf392ef6} /* (14, 21, 9) {real, imag} */,
  {32'h40605161, 32'h3fddcd6e} /* (14, 21, 8) {real, imag} */,
  {32'h401c14a4, 32'h404892a4} /* (14, 21, 7) {real, imag} */,
  {32'h3ef7a048, 32'h3fd2d49b} /* (14, 21, 6) {real, imag} */,
  {32'h3ffb4c6a, 32'hbe934470} /* (14, 21, 5) {real, imag} */,
  {32'h3fb017c6, 32'h3f1a00a4} /* (14, 21, 4) {real, imag} */,
  {32'h3e38b5a0, 32'hbf67243a} /* (14, 21, 3) {real, imag} */,
  {32'hbf1b9755, 32'hc076b4f9} /* (14, 21, 2) {real, imag} */,
  {32'h4027a89f, 32'hc04b818d} /* (14, 21, 1) {real, imag} */,
  {32'h406daddd, 32'hbfe37588} /* (14, 21, 0) {real, imag} */,
  {32'h3f2dd11e, 32'hc00fab6b} /* (14, 20, 31) {real, imag} */,
  {32'h4005be09, 32'hc0083148} /* (14, 20, 30) {real, imag} */,
  {32'h404013ee, 32'h3e9f6b18} /* (14, 20, 29) {real, imag} */,
  {32'h40242788, 32'h3f146854} /* (14, 20, 28) {real, imag} */,
  {32'h3ef1313c, 32'h3ea49880} /* (14, 20, 27) {real, imag} */,
  {32'hbff7e1ac, 32'h3e8586bc} /* (14, 20, 26) {real, imag} */,
  {32'hbf8ad0e4, 32'h3fb0b624} /* (14, 20, 25) {real, imag} */,
  {32'hbf2cfa28, 32'h3dc0c550} /* (14, 20, 24) {real, imag} */,
  {32'hbdf6bfc8, 32'h3d949390} /* (14, 20, 23) {real, imag} */,
  {32'h402cabdb, 32'hbf9fb8f3} /* (14, 20, 22) {real, imag} */,
  {32'h3f591ca6, 32'hbf723080} /* (14, 20, 21) {real, imag} */,
  {32'hbf9878d2, 32'hbfdfcfea} /* (14, 20, 20) {real, imag} */,
  {32'hbeca9d88, 32'hbeb1e640} /* (14, 20, 19) {real, imag} */,
  {32'hbf265c89, 32'hbfdff888} /* (14, 20, 18) {real, imag} */,
  {32'h3f571cec, 32'hc04e1abb} /* (14, 20, 17) {real, imag} */,
  {32'h3fb98817, 32'h3e2bc698} /* (14, 20, 16) {real, imag} */,
  {32'h3f664728, 32'h4050e75f} /* (14, 20, 15) {real, imag} */,
  {32'h3f04d35e, 32'h4034a891} /* (14, 20, 14) {real, imag} */,
  {32'h3fd01609, 32'h4080cb86} /* (14, 20, 13) {real, imag} */,
  {32'h3e8eab18, 32'h407b8334} /* (14, 20, 12) {real, imag} */,
  {32'h3fad704a, 32'hc005bfea} /* (14, 20, 11) {real, imag} */,
  {32'h3eb46fc4, 32'hbf23a172} /* (14, 20, 10) {real, imag} */,
  {32'h3e896f1c, 32'h3fa9e8fe} /* (14, 20, 9) {real, imag} */,
  {32'h3ffcf30a, 32'hbfaff2ae} /* (14, 20, 8) {real, imag} */,
  {32'hbf87218b, 32'hbd7e4d10} /* (14, 20, 7) {real, imag} */,
  {32'hbfd9c9ae, 32'h40333971} /* (14, 20, 6) {real, imag} */,
  {32'h3faf2f10, 32'h3f64c338} /* (14, 20, 5) {real, imag} */,
  {32'h3ff4cc6e, 32'hbfc66234} /* (14, 20, 4) {real, imag} */,
  {32'hbc542d00, 32'hc04a3a41} /* (14, 20, 3) {real, imag} */,
  {32'h3f0db810, 32'hc00401ee} /* (14, 20, 2) {real, imag} */,
  {32'hbfea1df4, 32'h40090df4} /* (14, 20, 1) {real, imag} */,
  {32'hbfbf3f6c, 32'h3fa64c12} /* (14, 20, 0) {real, imag} */,
  {32'h3f9ab9f0, 32'hbd878890} /* (14, 19, 31) {real, imag} */,
  {32'h3db976a0, 32'hbe259570} /* (14, 19, 30) {real, imag} */,
  {32'hbf6b5d6a, 32'h3f49fc2a} /* (14, 19, 29) {real, imag} */,
  {32'hbfd352a7, 32'h3ef6a418} /* (14, 19, 28) {real, imag} */,
  {32'hc0401c98, 32'h3fa9e0fe} /* (14, 19, 27) {real, imag} */,
  {32'hbf3f3904, 32'h3f0d17ee} /* (14, 19, 26) {real, imag} */,
  {32'h3fa1d096, 32'h3f9bfc24} /* (14, 19, 25) {real, imag} */,
  {32'h3cce7440, 32'h40469f08} /* (14, 19, 24) {real, imag} */,
  {32'hbec17408, 32'h3fff0a52} /* (14, 19, 23) {real, imag} */,
  {32'hbfbe4c5f, 32'h4006ac2f} /* (14, 19, 22) {real, imag} */,
  {32'hbfd60a22, 32'hbd230ad0} /* (14, 19, 21) {real, imag} */,
  {32'hbdf675b0, 32'hbf2c9c88} /* (14, 19, 20) {real, imag} */,
  {32'h3ed09c14, 32'hbf04c7f3} /* (14, 19, 19) {real, imag} */,
  {32'hbfd0b784, 32'h3fa4ffda} /* (14, 19, 18) {real, imag} */,
  {32'hbfb8dad9, 32'h3febe3fd} /* (14, 19, 17) {real, imag} */,
  {32'h3de79588, 32'h3f0c8052} /* (14, 19, 16) {real, imag} */,
  {32'h3f9159e0, 32'h3f5c27c9} /* (14, 19, 15) {real, imag} */,
  {32'hbf9e4e74, 32'h3f2c4af4} /* (14, 19, 14) {real, imag} */,
  {32'hbfcda936, 32'hbf3ee52c} /* (14, 19, 13) {real, imag} */,
  {32'hbf363754, 32'h3ee3fb2a} /* (14, 19, 12) {real, imag} */,
  {32'h3f69cf60, 32'hbd263460} /* (14, 19, 11) {real, imag} */,
  {32'h3e984fb6, 32'hc02661f6} /* (14, 19, 10) {real, imag} */,
  {32'h3ec4b7d4, 32'hc02a19ea} /* (14, 19, 9) {real, imag} */,
  {32'h3efd2d52, 32'hbf9c78f2} /* (14, 19, 8) {real, imag} */,
  {32'h3fe0f374, 32'h3fdb8f64} /* (14, 19, 7) {real, imag} */,
  {32'h3e4f83ea, 32'h3fd6d016} /* (14, 19, 6) {real, imag} */,
  {32'h3e6349f4, 32'hbf3665cc} /* (14, 19, 5) {real, imag} */,
  {32'h3eee850c, 32'h3fb98596} /* (14, 19, 4) {real, imag} */,
  {32'hbf824dee, 32'h3f94b18a} /* (14, 19, 3) {real, imag} */,
  {32'hbff972b2, 32'h3fb62ccc} /* (14, 19, 2) {real, imag} */,
  {32'hc062279a, 32'h3ed448fe} /* (14, 19, 1) {real, imag} */,
  {32'hbffa76f7, 32'hbf1881e6} /* (14, 19, 0) {real, imag} */,
  {32'hbe833a30, 32'h3f29d4e0} /* (14, 18, 31) {real, imag} */,
  {32'hbf7ae61c, 32'hbff765ae} /* (14, 18, 30) {real, imag} */,
  {32'hbfb00521, 32'hbf25168c} /* (14, 18, 29) {real, imag} */,
  {32'hbf95bee6, 32'hbfbef6f8} /* (14, 18, 28) {real, imag} */,
  {32'hbf525b58, 32'hbfa8100f} /* (14, 18, 27) {real, imag} */,
  {32'h3f43bc9a, 32'h3fa5195a} /* (14, 18, 26) {real, imag} */,
  {32'hbf4b775f, 32'h3f746184} /* (14, 18, 25) {real, imag} */,
  {32'hbf2d697d, 32'hbf8a56d2} /* (14, 18, 24) {real, imag} */,
  {32'h40060c52, 32'hbff4e86e} /* (14, 18, 23) {real, imag} */,
  {32'hbe805198, 32'h3dfa2f54} /* (14, 18, 22) {real, imag} */,
  {32'hbfb863c4, 32'h3f5ea8af} /* (14, 18, 21) {real, imag} */,
  {32'hbe83fb40, 32'h3f574ee2} /* (14, 18, 20) {real, imag} */,
  {32'hbf4313ab, 32'h3ffcb853} /* (14, 18, 19) {real, imag} */,
  {32'hbef97df8, 32'h4013a7ab} /* (14, 18, 18) {real, imag} */,
  {32'hbf319a26, 32'h3e23df70} /* (14, 18, 17) {real, imag} */,
  {32'h3f9bcd2c, 32'hbf3c8ef4} /* (14, 18, 16) {real, imag} */,
  {32'h3fdc02d7, 32'hbe1faff0} /* (14, 18, 15) {real, imag} */,
  {32'hbe4f1e60, 32'hbf26de3f} /* (14, 18, 14) {real, imag} */,
  {32'h3f2fe898, 32'hbe999850} /* (14, 18, 13) {real, imag} */,
  {32'hbe629708, 32'h3fd3ca5d} /* (14, 18, 12) {real, imag} */,
  {32'hbfc81360, 32'h3f30cbb4} /* (14, 18, 11) {real, imag} */,
  {32'hbf9d5796, 32'hbf0ffd1b} /* (14, 18, 10) {real, imag} */,
  {32'hbebc35dc, 32'h3f0a454e} /* (14, 18, 9) {real, imag} */,
  {32'h3f8e7ec0, 32'h3ea014d4} /* (14, 18, 8) {real, imag} */,
  {32'hbf8c9f7e, 32'hbf1562c0} /* (14, 18, 7) {real, imag} */,
  {32'hbed4623c, 32'hbfc78da7} /* (14, 18, 6) {real, imag} */,
  {32'h3dbe8db0, 32'hbf54efff} /* (14, 18, 5) {real, imag} */,
  {32'hbc249e40, 32'hbdf0dd64} /* (14, 18, 4) {real, imag} */,
  {32'h3ed0cc00, 32'h3e744666} /* (14, 18, 3) {real, imag} */,
  {32'h400403e7, 32'h3e1c61e0} /* (14, 18, 2) {real, imag} */,
  {32'h3f7a29be, 32'hc02bae85} /* (14, 18, 1) {real, imag} */,
  {32'h3bcbb080, 32'hbec01826} /* (14, 18, 0) {real, imag} */,
  {32'h3f7303e4, 32'hbfcf3c91} /* (14, 17, 31) {real, imag} */,
  {32'h3db0f708, 32'hbfc10898} /* (14, 17, 30) {real, imag} */,
  {32'hbf13ac3a, 32'hbfc42eba} /* (14, 17, 29) {real, imag} */,
  {32'hbd03d120, 32'h3ed98f4a} /* (14, 17, 28) {real, imag} */,
  {32'hbf86419f, 32'h3f95a1fe} /* (14, 17, 27) {real, imag} */,
  {32'hbe0e0120, 32'hbef310ac} /* (14, 17, 26) {real, imag} */,
  {32'h3f92aae4, 32'hbfa96e77} /* (14, 17, 25) {real, imag} */,
  {32'h3f19e834, 32'hbf43ffee} /* (14, 17, 24) {real, imag} */,
  {32'hbfb060b8, 32'hbf7f3ff9} /* (14, 17, 23) {real, imag} */,
  {32'hbdfae560, 32'hbebbef0d} /* (14, 17, 22) {real, imag} */,
  {32'hbd1569a0, 32'h3f040883} /* (14, 17, 21) {real, imag} */,
  {32'h3f940593, 32'hbda4eae8} /* (14, 17, 20) {real, imag} */,
  {32'h3fa626a4, 32'hbe0deb2a} /* (14, 17, 19) {real, imag} */,
  {32'hbf93cd2c, 32'h3f2def88} /* (14, 17, 18) {real, imag} */,
  {32'hbea430c0, 32'h3e8418b8} /* (14, 17, 17) {real, imag} */,
  {32'h3f26612a, 32'hbdaea5c4} /* (14, 17, 16) {real, imag} */,
  {32'hbf5d140d, 32'hbf92933c} /* (14, 17, 15) {real, imag} */,
  {32'h3e665c84, 32'hbefcadd7} /* (14, 17, 14) {real, imag} */,
  {32'hbe7352b0, 32'h3e12789c} /* (14, 17, 13) {real, imag} */,
  {32'h3f9076d7, 32'h3f9c4b40} /* (14, 17, 12) {real, imag} */,
  {32'h4013d6ec, 32'h3f95aaae} /* (14, 17, 11) {real, imag} */,
  {32'h400e132c, 32'h3f0cfe64} /* (14, 17, 10) {real, imag} */,
  {32'h3f2007a8, 32'hbee005f8} /* (14, 17, 9) {real, imag} */,
  {32'hbf9c7bd9, 32'hbf7ed8f8} /* (14, 17, 8) {real, imag} */,
  {32'h3f0087fe, 32'hbf5f62ab} /* (14, 17, 7) {real, imag} */,
  {32'hbee5bb80, 32'h3e91dc68} /* (14, 17, 6) {real, imag} */,
  {32'hc00b955c, 32'h400c0c02} /* (14, 17, 5) {real, imag} */,
  {32'h3ec49ec8, 32'h3f5443d0} /* (14, 17, 4) {real, imag} */,
  {32'h3fa0f618, 32'h3fc81560} /* (14, 17, 3) {real, imag} */,
  {32'hbf9aec10, 32'h3f4bfa2f} /* (14, 17, 2) {real, imag} */,
  {32'h3debbe30, 32'hbebe6304} /* (14, 17, 1) {real, imag} */,
  {32'h3e9e9f05, 32'h3e71a1a4} /* (14, 17, 0) {real, imag} */,
  {32'hbee380f8, 32'hbcae5d80} /* (14, 16, 31) {real, imag} */,
  {32'h3e1b1a40, 32'hbf7d04dc} /* (14, 16, 30) {real, imag} */,
  {32'hbe33c43c, 32'hbfdb7328} /* (14, 16, 29) {real, imag} */,
  {32'hbf0d41ba, 32'hbf291148} /* (14, 16, 28) {real, imag} */,
  {32'hbccf1700, 32'h3f5084d8} /* (14, 16, 27) {real, imag} */,
  {32'h3f5447d0, 32'h3f00ad10} /* (14, 16, 26) {real, imag} */,
  {32'h3eb4f060, 32'h3d883ea0} /* (14, 16, 25) {real, imag} */,
  {32'hbe43f620, 32'hbd8d5fe0} /* (14, 16, 24) {real, imag} */,
  {32'h3e0517d0, 32'hbf9a36b2} /* (14, 16, 23) {real, imag} */,
  {32'hbf1b9998, 32'hbe9c3b30} /* (14, 16, 22) {real, imag} */,
  {32'hbfc9a588, 32'h3f8718b7} /* (14, 16, 21) {real, imag} */,
  {32'hbfd9f490, 32'hbee974ec} /* (14, 16, 20) {real, imag} */,
  {32'hbeae2cac, 32'hbf1be314} /* (14, 16, 19) {real, imag} */,
  {32'h3e2f8200, 32'h3e229880} /* (14, 16, 18) {real, imag} */,
  {32'hbedd7fdc, 32'h3fbef9d8} /* (14, 16, 17) {real, imag} */,
  {32'hbf2485b7, 32'h3f92ff9c} /* (14, 16, 16) {real, imag} */,
  {32'hbe21c020, 32'h3fb0fa2c} /* (14, 16, 15) {real, imag} */,
  {32'h3f2e6dac, 32'h3fd24d24} /* (14, 16, 14) {real, imag} */,
  {32'h3f99edab, 32'h3f3a6544} /* (14, 16, 13) {real, imag} */,
  {32'h3f4f67b5, 32'h3fa71b36} /* (14, 16, 12) {real, imag} */,
  {32'h3faf6661, 32'h3eb5d698} /* (14, 16, 11) {real, imag} */,
  {32'h3fd8ed88, 32'hbf8b2e44} /* (14, 16, 10) {real, imag} */,
  {32'h3f4a7c08, 32'hbf39f63c} /* (14, 16, 9) {real, imag} */,
  {32'h40196eda, 32'h3eafc930} /* (14, 16, 8) {real, imag} */,
  {32'h3fb9ea1c, 32'h3f7499c0} /* (14, 16, 7) {real, imag} */,
  {32'hbe15bce0, 32'hbd7f3480} /* (14, 16, 6) {real, imag} */,
  {32'hbf2eed10, 32'h3e85e7a0} /* (14, 16, 5) {real, imag} */,
  {32'hbf2da678, 32'hbfa09c14} /* (14, 16, 4) {real, imag} */,
  {32'hbcf60c00, 32'hbf838bea} /* (14, 16, 3) {real, imag} */,
  {32'hbf1c5bb8, 32'h3f29a9cc} /* (14, 16, 2) {real, imag} */,
  {32'h3e2dccbc, 32'h3e3f8c20} /* (14, 16, 1) {real, imag} */,
  {32'h3e20320c, 32'hbe4dc210} /* (14, 16, 0) {real, imag} */,
  {32'h3f23c0c4, 32'hbf4dd022} /* (14, 15, 31) {real, imag} */,
  {32'h3f01e37f, 32'hc00aadaa} /* (14, 15, 30) {real, imag} */,
  {32'h3efed134, 32'hbf163bbc} /* (14, 15, 29) {real, imag} */,
  {32'h3f8565e1, 32'hbdde3aee} /* (14, 15, 28) {real, imag} */,
  {32'h3e519338, 32'hbfa53bc4} /* (14, 15, 27) {real, imag} */,
  {32'h3d424080, 32'hbfe79221} /* (14, 15, 26) {real, imag} */,
  {32'hbfe5ebcc, 32'hbf0e562e} /* (14, 15, 25) {real, imag} */,
  {32'hbf848b9a, 32'hbec5478c} /* (14, 15, 24) {real, imag} */,
  {32'h3f3a7b10, 32'hbf368ba1} /* (14, 15, 23) {real, imag} */,
  {32'h3f3010c4, 32'hbfa2a7fb} /* (14, 15, 22) {real, imag} */,
  {32'hbeedb37c, 32'hc002f560} /* (14, 15, 21) {real, imag} */,
  {32'hbfd23277, 32'hbf8b35a4} /* (14, 15, 20) {real, imag} */,
  {32'h3f1bcdc3, 32'h3ef703a9} /* (14, 15, 19) {real, imag} */,
  {32'hbde3c4c0, 32'h4002bfea} /* (14, 15, 18) {real, imag} */,
  {32'hc012ed34, 32'h403b508d} /* (14, 15, 17) {real, imag} */,
  {32'hbf7658f2, 32'h3f414180} /* (14, 15, 16) {real, imag} */,
  {32'hbd78c8b0, 32'h3eea78c6} /* (14, 15, 15) {real, imag} */,
  {32'hbf4d3c31, 32'hbedbb5f1} /* (14, 15, 14) {real, imag} */,
  {32'hbeca6288, 32'h3c35a240} /* (14, 15, 13) {real, imag} */,
  {32'h3f161f9a, 32'h3f6a8078} /* (14, 15, 12) {real, imag} */,
  {32'h3e1c69e0, 32'h3f2ef2e7} /* (14, 15, 11) {real, imag} */,
  {32'hbdeaf5d0, 32'hbdf377a0} /* (14, 15, 10) {real, imag} */,
  {32'hbf061b44, 32'hbbae3200} /* (14, 15, 9) {real, imag} */,
  {32'hc00960f0, 32'h3f96e2dc} /* (14, 15, 8) {real, imag} */,
  {32'h3e681e48, 32'h3e80b32a} /* (14, 15, 7) {real, imag} */,
  {32'hbe3b9320, 32'hbfc5d2ee} /* (14, 15, 6) {real, imag} */,
  {32'hc010c698, 32'h3d8bcab0} /* (14, 15, 5) {real, imag} */,
  {32'hbff0e736, 32'hbf612980} /* (14, 15, 4) {real, imag} */,
  {32'hbfb794ac, 32'hbf0b27e3} /* (14, 15, 3) {real, imag} */,
  {32'hbfcf4e30, 32'h3f05a6d7} /* (14, 15, 2) {real, imag} */,
  {32'hbea8af6c, 32'h3effa358} /* (14, 15, 1) {real, imag} */,
  {32'h3f1dca16, 32'hbee6ab12} /* (14, 15, 0) {real, imag} */,
  {32'h3f892154, 32'h3f2a8d28} /* (14, 14, 31) {real, imag} */,
  {32'hbdc03ae0, 32'h3ed0c2de} /* (14, 14, 30) {real, imag} */,
  {32'hc006dc20, 32'hbef2c9b8} /* (14, 14, 29) {real, imag} */,
  {32'h3d979a18, 32'hbf2c7a68} /* (14, 14, 28) {real, imag} */,
  {32'h3fd2869c, 32'hbf09a8ee} /* (14, 14, 27) {real, imag} */,
  {32'h3f80f833, 32'hbf11e380} /* (14, 14, 26) {real, imag} */,
  {32'hbe392b64, 32'h3c97be80} /* (14, 14, 25) {real, imag} */,
  {32'hbef35446, 32'h3d637220} /* (14, 14, 24) {real, imag} */,
  {32'hbf991d97, 32'h3fc655da} /* (14, 14, 23) {real, imag} */,
  {32'hc0136895, 32'h3ed4db6b} /* (14, 14, 22) {real, imag} */,
  {32'h3f1125b0, 32'hbfb4ad84} /* (14, 14, 21) {real, imag} */,
  {32'h3f78cfe0, 32'hbf7505ae} /* (14, 14, 20) {real, imag} */,
  {32'hc00d71cd, 32'h3f071696} /* (14, 14, 19) {real, imag} */,
  {32'hc0258545, 32'h3ec6c918} /* (14, 14, 18) {real, imag} */,
  {32'hbfb7664d, 32'hbe4f45a0} /* (14, 14, 17) {real, imag} */,
  {32'hbe2faedc, 32'hbea93ec8} /* (14, 14, 16) {real, imag} */,
  {32'h3fe37d91, 32'hbd6f2ac0} /* (14, 14, 15) {real, imag} */,
  {32'h3fe99844, 32'hbf9402f0} /* (14, 14, 14) {real, imag} */,
  {32'h3fad6730, 32'hbf39da30} /* (14, 14, 13) {real, imag} */,
  {32'hbc64c780, 32'hbe082368} /* (14, 14, 12) {real, imag} */,
  {32'hbeb9c648, 32'h3f25e324} /* (14, 14, 11) {real, imag} */,
  {32'h3e8b5f88, 32'hbf6c3ca5} /* (14, 14, 10) {real, imag} */,
  {32'hbea090a4, 32'hbf83d5d1} /* (14, 14, 9) {real, imag} */,
  {32'hbf942d90, 32'h3f027616} /* (14, 14, 8) {real, imag} */,
  {32'h3f4cd7ac, 32'h402418d1} /* (14, 14, 7) {real, imag} */,
  {32'h4009c320, 32'h3fd60aa5} /* (14, 14, 6) {real, imag} */,
  {32'h3f2063ba, 32'hbe7fa7a4} /* (14, 14, 5) {real, imag} */,
  {32'hbfb814fc, 32'h3efd3e47} /* (14, 14, 4) {real, imag} */,
  {32'h3f474310, 32'hbe6d9fca} /* (14, 14, 3) {real, imag} */,
  {32'hbce31580, 32'hbf389314} /* (14, 14, 2) {real, imag} */,
  {32'hbf058e6e, 32'h3bb9a200} /* (14, 14, 1) {real, imag} */,
  {32'h3f910cd4, 32'hbf3e826d} /* (14, 14, 0) {real, imag} */,
  {32'hbf13d383, 32'h3fc6f2ef} /* (14, 13, 31) {real, imag} */,
  {32'h3fbfcf0a, 32'h3fcd86a6} /* (14, 13, 30) {real, imag} */,
  {32'h3ee81d24, 32'h3eeeae64} /* (14, 13, 29) {real, imag} */,
  {32'hbfe982cd, 32'h3f878f7e} /* (14, 13, 28) {real, imag} */,
  {32'hbf58984a, 32'hbfdcea8a} /* (14, 13, 27) {real, imag} */,
  {32'h3cd14690, 32'hbf9c5225} /* (14, 13, 26) {real, imag} */,
  {32'hbf3b6138, 32'h3e9a3e34} /* (14, 13, 25) {real, imag} */,
  {32'hbff6d64f, 32'hbfe8d730} /* (14, 13, 24) {real, imag} */,
  {32'hc03f2231, 32'hc048d0db} /* (14, 13, 23) {real, imag} */,
  {32'hbf85a93f, 32'hbe60c930} /* (14, 13, 22) {real, imag} */,
  {32'hbf70bb9c, 32'h3f8a1ef8} /* (14, 13, 21) {real, imag} */,
  {32'hbfd54adb, 32'hbffb0740} /* (14, 13, 20) {real, imag} */,
  {32'hbc402b80, 32'hbfb232f4} /* (14, 13, 19) {real, imag} */,
  {32'hbebe05ce, 32'h40088969} /* (14, 13, 18) {real, imag} */,
  {32'hc01b6162, 32'h3eb6fa44} /* (14, 13, 17) {real, imag} */,
  {32'hbfb70f1c, 32'hbf6cdb3a} /* (14, 13, 16) {real, imag} */,
  {32'hbe69479c, 32'h3f7596ad} /* (14, 13, 15) {real, imag} */,
  {32'hbe5b4bac, 32'h3f762414} /* (14, 13, 14) {real, imag} */,
  {32'h3f8e7f38, 32'h3f82ac0e} /* (14, 13, 13) {real, imag} */,
  {32'hc0163b95, 32'h3ed13ab2} /* (14, 13, 12) {real, imag} */,
  {32'hc056608a, 32'h3e8f8b14} /* (14, 13, 11) {real, imag} */,
  {32'hbfff4b68, 32'hc0034d4a} /* (14, 13, 10) {real, imag} */,
  {32'hbfbaa655, 32'hbeb66e68} /* (14, 13, 9) {real, imag} */,
  {32'hbe6a65c4, 32'hbee6cad8} /* (14, 13, 8) {real, imag} */,
  {32'h3cf14e00, 32'hbf440060} /* (14, 13, 7) {real, imag} */,
  {32'hbda67fb4, 32'hc02326cd} /* (14, 13, 6) {real, imag} */,
  {32'hbf2d4c9b, 32'hc0651635} /* (14, 13, 5) {real, imag} */,
  {32'hc01955e6, 32'hbd7092b0} /* (14, 13, 4) {real, imag} */,
  {32'hbecdd738, 32'h3fa72134} /* (14, 13, 3) {real, imag} */,
  {32'hbf0ed384, 32'hbd152790} /* (14, 13, 2) {real, imag} */,
  {32'hbfa18619, 32'hbf1c0057} /* (14, 13, 1) {real, imag} */,
  {32'hbf4e93f6, 32'h3eaf2ab4} /* (14, 13, 0) {real, imag} */,
  {32'hc011a4aa, 32'hbfa60270} /* (14, 12, 31) {real, imag} */,
  {32'hc0404609, 32'hc036ba66} /* (14, 12, 30) {real, imag} */,
  {32'hbe83a8f0, 32'hc099059c} /* (14, 12, 29) {real, imag} */,
  {32'h3f3d6582, 32'hc091fec4} /* (14, 12, 28) {real, imag} */,
  {32'hbf594d2a, 32'hc01d53a4} /* (14, 12, 27) {real, imag} */,
  {32'h3ffe5550, 32'hbfb2b5a5} /* (14, 12, 26) {real, imag} */,
  {32'h3ff9d16a, 32'h3df61260} /* (14, 12, 25) {real, imag} */,
  {32'hbf32be2c, 32'h404077ce} /* (14, 12, 24) {real, imag} */,
  {32'h3f78fcdf, 32'h3f8612d5} /* (14, 12, 23) {real, imag} */,
  {32'h3d707b40, 32'hbf9bedc1} /* (14, 12, 22) {real, imag} */,
  {32'hc04933b8, 32'hc04f9e38} /* (14, 12, 21) {real, imag} */,
  {32'hc02cbecd, 32'hc03da859} /* (14, 12, 20) {real, imag} */,
  {32'h3fc71922, 32'hc00b2b4c} /* (14, 12, 19) {real, imag} */,
  {32'h40085ab4, 32'hbf68847c} /* (14, 12, 18) {real, imag} */,
  {32'h3fe4f1b6, 32'h3ff1ba7a} /* (14, 12, 17) {real, imag} */,
  {32'h3f305852, 32'h3e8c6c6c} /* (14, 12, 16) {real, imag} */,
  {32'hbfb46538, 32'h3d0264c0} /* (14, 12, 15) {real, imag} */,
  {32'hbed9ff78, 32'h3e888e88} /* (14, 12, 14) {real, imag} */,
  {32'hbfd88545, 32'hbfc8c6e6} /* (14, 12, 13) {real, imag} */,
  {32'hbfdd9a3e, 32'hbf4ab0d0} /* (14, 12, 12) {real, imag} */,
  {32'hbff9238e, 32'h400ff512} /* (14, 12, 11) {real, imag} */,
  {32'h3f62606c, 32'hbe994f5f} /* (14, 12, 10) {real, imag} */,
  {32'h3fc3f227, 32'hc06768d9} /* (14, 12, 9) {real, imag} */,
  {32'h3f7b37ac, 32'hbe3ddeb0} /* (14, 12, 8) {real, imag} */,
  {32'h3f63f81e, 32'h3dd4b9c8} /* (14, 12, 7) {real, imag} */,
  {32'h3fc4d392, 32'h3f86d756} /* (14, 12, 6) {real, imag} */,
  {32'h3f089870, 32'hbfaf80de} /* (14, 12, 5) {real, imag} */,
  {32'hbfb28c3a, 32'hbd438100} /* (14, 12, 4) {real, imag} */,
  {32'hbe6ca250, 32'hbeace848} /* (14, 12, 3) {real, imag} */,
  {32'h3f321600, 32'hbfa97218} /* (14, 12, 2) {real, imag} */,
  {32'h3fce7df8, 32'hc0084484} /* (14, 12, 1) {real, imag} */,
  {32'hbf577c3d, 32'hbfcccc8e} /* (14, 12, 0) {real, imag} */,
  {32'hc01001e6, 32'hbfc5fac9} /* (14, 11, 31) {real, imag} */,
  {32'hc0532f8a, 32'hbe2c7c18} /* (14, 11, 30) {real, imag} */,
  {32'hc03891ca, 32'h4001f6fa} /* (14, 11, 29) {real, imag} */,
  {32'hbf52b842, 32'h4073449f} /* (14, 11, 28) {real, imag} */,
  {32'h3e2c9fb4, 32'h40266420} /* (14, 11, 27) {real, imag} */,
  {32'hbf866aec, 32'hbfc2428f} /* (14, 11, 26) {real, imag} */,
  {32'hbd0c0980, 32'hbe1fa440} /* (14, 11, 25) {real, imag} */,
  {32'hbed0737c, 32'h400d58c7} /* (14, 11, 24) {real, imag} */,
  {32'h400c11ba, 32'hbdfaec90} /* (14, 11, 23) {real, imag} */,
  {32'hbef02e08, 32'hbec47d5a} /* (14, 11, 22) {real, imag} */,
  {32'h40209dd6, 32'hbe9ae42c} /* (14, 11, 21) {real, imag} */,
  {32'h402a99cb, 32'h3f87fa8a} /* (14, 11, 20) {real, imag} */,
  {32'hbf5b756d, 32'h3f69546c} /* (14, 11, 19) {real, imag} */,
  {32'hc0030720, 32'h3f919dce} /* (14, 11, 18) {real, imag} */,
  {32'hbfc2f4b9, 32'hc019c7ff} /* (14, 11, 17) {real, imag} */,
  {32'hbf30bad1, 32'hbf8568b5} /* (14, 11, 16) {real, imag} */,
  {32'h3df4e500, 32'hc064ddc4} /* (14, 11, 15) {real, imag} */,
  {32'h3f04b052, 32'hbfc7cc20} /* (14, 11, 14) {real, imag} */,
  {32'hbe21f1a8, 32'h3fe1e07b} /* (14, 11, 13) {real, imag} */,
  {32'h3eb75921, 32'h405d94fe} /* (14, 11, 12) {real, imag} */,
  {32'h3eaff75a, 32'h3f1b8c4a} /* (14, 11, 11) {real, imag} */,
  {32'h3f41a029, 32'h3f3256eb} /* (14, 11, 10) {real, imag} */,
  {32'h3f5361de, 32'hbeea32ac} /* (14, 11, 9) {real, imag} */,
  {32'h3f0fa9ac, 32'h3fecdcb6} /* (14, 11, 8) {real, imag} */,
  {32'hbfd4bf99, 32'h3fecdb53} /* (14, 11, 7) {real, imag} */,
  {32'h3e0d2cd0, 32'h404dd110} /* (14, 11, 6) {real, imag} */,
  {32'h3f2c6950, 32'h407466aa} /* (14, 11, 5) {real, imag} */,
  {32'hbf071594, 32'h3f6bddc8} /* (14, 11, 4) {real, imag} */,
  {32'h406e3070, 32'hc006133a} /* (14, 11, 3) {real, imag} */,
  {32'h3db2d8f8, 32'hc0390401} /* (14, 11, 2) {real, imag} */,
  {32'h3f903c2a, 32'hbeec9a38} /* (14, 11, 1) {real, imag} */,
  {32'h3f98bf3e, 32'hbe8bf856} /* (14, 11, 0) {real, imag} */,
  {32'h3ed9f570, 32'h3ff2d621} /* (14, 10, 31) {real, imag} */,
  {32'hc06487f6, 32'h4023a698} /* (14, 10, 30) {real, imag} */,
  {32'hbf8c9c6a, 32'h3fe8b24a} /* (14, 10, 29) {real, imag} */,
  {32'h3fd98dca, 32'h3f39d638} /* (14, 10, 28) {real, imag} */,
  {32'h4093c5ac, 32'h403120da} /* (14, 10, 27) {real, imag} */,
  {32'h404fb063, 32'h406b789c} /* (14, 10, 26) {real, imag} */,
  {32'h401ab55d, 32'hbf2b12f3} /* (14, 10, 25) {real, imag} */,
  {32'hbf970d6c, 32'h3fa8ac8c} /* (14, 10, 24) {real, imag} */,
  {32'h3f82b29a, 32'hbf9e472b} /* (14, 10, 23) {real, imag} */,
  {32'h40a785f8, 32'hc0603ff8} /* (14, 10, 22) {real, imag} */,
  {32'h40125d6a, 32'hbfb12122} /* (14, 10, 21) {real, imag} */,
  {32'h4040ff51, 32'h3e2eff50} /* (14, 10, 20) {real, imag} */,
  {32'h40294d1c, 32'h3d7008c0} /* (14, 10, 19) {real, imag} */,
  {32'h40869e9d, 32'hbffcfa59} /* (14, 10, 18) {real, imag} */,
  {32'h408fea75, 32'hc0403a2a} /* (14, 10, 17) {real, imag} */,
  {32'h402fd9c3, 32'hbf64b8c2} /* (14, 10, 16) {real, imag} */,
  {32'h3fcf9df0, 32'h3c41f200} /* (14, 10, 15) {real, imag} */,
  {32'hbfc242d8, 32'h4049c5d2} /* (14, 10, 14) {real, imag} */,
  {32'hbeadc050, 32'h3faace96} /* (14, 10, 13) {real, imag} */,
  {32'hbfa35e59, 32'hbf6af774} /* (14, 10, 12) {real, imag} */,
  {32'h3fe024de, 32'h4025dd37} /* (14, 10, 11) {real, imag} */,
  {32'h3c1b9880, 32'h3e913078} /* (14, 10, 10) {real, imag} */,
  {32'h3e6c52f8, 32'hbc620000} /* (14, 10, 9) {real, imag} */,
  {32'hc025d774, 32'hc0421b0d} /* (14, 10, 8) {real, imag} */,
  {32'hc0535a64, 32'hbfcfcf2d} /* (14, 10, 7) {real, imag} */,
  {32'h3fac560a, 32'hc060b041} /* (14, 10, 6) {real, imag} */,
  {32'h3fcf837e, 32'hc00c4efd} /* (14, 10, 5) {real, imag} */,
  {32'hc01a1a50, 32'h3f8176e5} /* (14, 10, 4) {real, imag} */,
  {32'hbec3e294, 32'hc011b2ab} /* (14, 10, 3) {real, imag} */,
  {32'hbf978b15, 32'hbeccb51a} /* (14, 10, 2) {real, imag} */,
  {32'h3f9c6bf2, 32'h3ff97464} /* (14, 10, 1) {real, imag} */,
  {32'h3fcb125e, 32'hbe988392} /* (14, 10, 0) {real, imag} */,
  {32'h3dbc6bd8, 32'hbf82a0cd} /* (14, 9, 31) {real, imag} */,
  {32'hbc120480, 32'hc01c37b0} /* (14, 9, 30) {real, imag} */,
  {32'h40518ea3, 32'hbfb20f1e} /* (14, 9, 29) {real, imag} */,
  {32'h409d14a1, 32'hbf890eb4} /* (14, 9, 28) {real, imag} */,
  {32'h3fdfbf28, 32'h4025c70a} /* (14, 9, 27) {real, imag} */,
  {32'h3f6445d4, 32'h401a3cec} /* (14, 9, 26) {real, imag} */,
  {32'hc010f6b8, 32'h39c75800} /* (14, 9, 25) {real, imag} */,
  {32'hc052c5a9, 32'h3fe316be} /* (14, 9, 24) {real, imag} */,
  {32'h3f12493a, 32'hc01a03cc} /* (14, 9, 23) {real, imag} */,
  {32'h402863f4, 32'hc01793d6} /* (14, 9, 22) {real, imag} */,
  {32'hbff275a1, 32'h40a9775d} /* (14, 9, 21) {real, imag} */,
  {32'h3f9f2ef6, 32'h40736b4a} /* (14, 9, 20) {real, imag} */,
  {32'h3c980280, 32'h3fc58ad7} /* (14, 9, 19) {real, imag} */,
  {32'hc02590a5, 32'hbf90ee96} /* (14, 9, 18) {real, imag} */,
  {32'hc09f4b9d, 32'hc0266000} /* (14, 9, 17) {real, imag} */,
  {32'h3fcf2ad2, 32'hbfa98a9e} /* (14, 9, 16) {real, imag} */,
  {32'h402b12b6, 32'hbf97c022} /* (14, 9, 15) {real, imag} */,
  {32'h4056a0d4, 32'h3fdeee8d} /* (14, 9, 14) {real, imag} */,
  {32'h40511c5c, 32'h3d331ec0} /* (14, 9, 13) {real, imag} */,
  {32'h3f8ae374, 32'hbf075130} /* (14, 9, 12) {real, imag} */,
  {32'h3e6b2230, 32'h3ee0ce28} /* (14, 9, 11) {real, imag} */,
  {32'hbf8d230d, 32'hbee0560a} /* (14, 9, 10) {real, imag} */,
  {32'hc026709b, 32'h404b1176} /* (14, 9, 9) {real, imag} */,
  {32'hc07604a8, 32'h3e9cc534} /* (14, 9, 8) {real, imag} */,
  {32'hbf71c594, 32'hc02a7328} /* (14, 9, 7) {real, imag} */,
  {32'h3fb90b02, 32'hc09c6e22} /* (14, 9, 6) {real, imag} */,
  {32'h403f56d2, 32'hc0b94680} /* (14, 9, 5) {real, imag} */,
  {32'h40aa60cd, 32'hc0d0da6f} /* (14, 9, 4) {real, imag} */,
  {32'h4078e968, 32'hbf6b85e9} /* (14, 9, 3) {real, imag} */,
  {32'h3f56173a, 32'hbf22af54} /* (14, 9, 2) {real, imag} */,
  {32'hc02c909c, 32'hbf530ce4} /* (14, 9, 1) {real, imag} */,
  {32'hbff6783c, 32'hbf9568bf} /* (14, 9, 0) {real, imag} */,
  {32'h3fe4ac10, 32'h40858935} /* (14, 8, 31) {real, imag} */,
  {32'h3f781532, 32'h4095ec15} /* (14, 8, 30) {real, imag} */,
  {32'hbe9261a8, 32'h3f16a1e0} /* (14, 8, 29) {real, imag} */,
  {32'h3f13d630, 32'hbf0fd080} /* (14, 8, 28) {real, imag} */,
  {32'h4030d910, 32'h400cd6f1} /* (14, 8, 27) {real, imag} */,
  {32'h3d5adbc0, 32'h3f0b5ce4} /* (14, 8, 26) {real, imag} */,
  {32'hbf967eae, 32'h3e13e370} /* (14, 8, 25) {real, imag} */,
  {32'hc0861cc1, 32'h3d2445a0} /* (14, 8, 24) {real, imag} */,
  {32'hc04fcd7e, 32'h402ea5a6} /* (14, 8, 23) {real, imag} */,
  {32'hbfe169ef, 32'hc00eba58} /* (14, 8, 22) {real, imag} */,
  {32'hc03729b0, 32'hc066918e} /* (14, 8, 21) {real, imag} */,
  {32'hc09e1b8d, 32'h406d467d} /* (14, 8, 20) {real, imag} */,
  {32'hbf04db9e, 32'hbfcfa5d8} /* (14, 8, 19) {real, imag} */,
  {32'h3fa49715, 32'hc0439c70} /* (14, 8, 18) {real, imag} */,
  {32'hbf884cec, 32'h3df86b70} /* (14, 8, 17) {real, imag} */,
  {32'hbfea1254, 32'h40331a4e} /* (14, 8, 16) {real, imag} */,
  {32'hc0ad0d26, 32'h3ff3dc42} /* (14, 8, 15) {real, imag} */,
  {32'hc08624b0, 32'hc008e937} /* (14, 8, 14) {real, imag} */,
  {32'h3f32ca72, 32'hc05b5bf7} /* (14, 8, 13) {real, imag} */,
  {32'hbf4db74c, 32'hc058dc91} /* (14, 8, 12) {real, imag} */,
  {32'h3e92a54c, 32'hc08b19fe} /* (14, 8, 11) {real, imag} */,
  {32'h3edb1fea, 32'hc033b20e} /* (14, 8, 10) {real, imag} */,
  {32'h4020851e, 32'hbf4e4190} /* (14, 8, 9) {real, imag} */,
  {32'h3f6280b4, 32'h40086886} /* (14, 8, 8) {real, imag} */,
  {32'h3f2edb84, 32'h3dbc7d20} /* (14, 8, 7) {real, imag} */,
  {32'h3f192c00, 32'hc03d937a} /* (14, 8, 6) {real, imag} */,
  {32'h4055bb93, 32'h40416f8e} /* (14, 8, 5) {real, imag} */,
  {32'h40061ec1, 32'h409b9b4c} /* (14, 8, 4) {real, imag} */,
  {32'h4018d911, 32'h405ae00e} /* (14, 8, 3) {real, imag} */,
  {32'h40b0f4be, 32'h40378d06} /* (14, 8, 2) {real, imag} */,
  {32'h406d34bb, 32'hc06829e2} /* (14, 8, 1) {real, imag} */,
  {32'hbf63b8f4, 32'hc03caa1e} /* (14, 8, 0) {real, imag} */,
  {32'h401eb7be, 32'h3e4c0460} /* (14, 7, 31) {real, imag} */,
  {32'h400e73b7, 32'hc0392b28} /* (14, 7, 30) {real, imag} */,
  {32'h3f4ec283, 32'hc0c53a6f} /* (14, 7, 29) {real, imag} */,
  {32'hbfa905c7, 32'hc082ddb8} /* (14, 7, 28) {real, imag} */,
  {32'hc0dc1a90, 32'h3fd3ff7c} /* (14, 7, 27) {real, imag} */,
  {32'hc08f02e0, 32'h3d86f820} /* (14, 7, 26) {real, imag} */,
  {32'hbfdefcd7, 32'hbf38dd78} /* (14, 7, 25) {real, imag} */,
  {32'hbe484724, 32'hbfe07422} /* (14, 7, 24) {real, imag} */,
  {32'h3faa16dd, 32'h403b4a64} /* (14, 7, 23) {real, imag} */,
  {32'h40a425aa, 32'h40de84fe} /* (14, 7, 22) {real, imag} */,
  {32'h4010d0d2, 32'h40d090ca} /* (14, 7, 21) {real, imag} */,
  {32'hc03cd8a8, 32'h40bdb604} /* (14, 7, 20) {real, imag} */,
  {32'hc0c66d10, 32'h408765de} /* (14, 7, 19) {real, imag} */,
  {32'hc0e9cb5a, 32'h3ff8262a} /* (14, 7, 18) {real, imag} */,
  {32'hc054ac42, 32'hbfb03cee} /* (14, 7, 17) {real, imag} */,
  {32'h4002b668, 32'h3cb724a0} /* (14, 7, 16) {real, imag} */,
  {32'h40c2fe8e, 32'h3f1ff238} /* (14, 7, 15) {real, imag} */,
  {32'hbe257cb8, 32'h3ffa3633} /* (14, 7, 14) {real, imag} */,
  {32'h4008ae27, 32'h3e51622c} /* (14, 7, 13) {real, imag} */,
  {32'h40861de4, 32'hc105986f} /* (14, 7, 12) {real, imag} */,
  {32'hbfe462a2, 32'hbfe6be7d} /* (14, 7, 11) {real, imag} */,
  {32'hbf81dba2, 32'h3e662a00} /* (14, 7, 10) {real, imag} */,
  {32'h3e9d4610, 32'hc0ec81b6} /* (14, 7, 9) {real, imag} */,
  {32'hbea8c738, 32'hc0b2ea96} /* (14, 7, 8) {real, imag} */,
  {32'h40270af9, 32'h3fce825c} /* (14, 7, 7) {real, imag} */,
  {32'h406d3384, 32'h3f83ccc6} /* (14, 7, 6) {real, imag} */,
  {32'h3e1d3948, 32'hbf90f954} /* (14, 7, 5) {real, imag} */,
  {32'hc0fe9f76, 32'hc0850be5} /* (14, 7, 4) {real, imag} */,
  {32'hc1090668, 32'hc08c1cfb} /* (14, 7, 3) {real, imag} */,
  {32'hc050aea0, 32'h3ee81758} /* (14, 7, 2) {real, imag} */,
  {32'hbf1407fe, 32'h403bebf4} /* (14, 7, 1) {real, imag} */,
  {32'hbee5249c, 32'hbf3af724} /* (14, 7, 0) {real, imag} */,
  {32'h407c03c5, 32'h3ff95b5b} /* (14, 6, 31) {real, imag} */,
  {32'h3f97701d, 32'hc007747e} /* (14, 6, 30) {real, imag} */,
  {32'hbf325694, 32'hbfe74e10} /* (14, 6, 29) {real, imag} */,
  {32'h3ef07826, 32'hbfe39046} /* (14, 6, 28) {real, imag} */,
  {32'h406927e6, 32'hbfba839a} /* (14, 6, 27) {real, imag} */,
  {32'h400b2e9a, 32'h3fd16ecf} /* (14, 6, 26) {real, imag} */,
  {32'hbf20c8a5, 32'h40497c37} /* (14, 6, 25) {real, imag} */,
  {32'hc0964a50, 32'h40265852} /* (14, 6, 24) {real, imag} */,
  {32'hc0deceb1, 32'hc016c714} /* (14, 6, 23) {real, imag} */,
  {32'hc01eba0d, 32'hc09986be} /* (14, 6, 22) {real, imag} */,
  {32'h3ffbe7f4, 32'h3f19dda8} /* (14, 6, 21) {real, imag} */,
  {32'hbfa08c19, 32'hbe445140} /* (14, 6, 20) {real, imag} */,
  {32'h403b6b0c, 32'hc0b2ccaa} /* (14, 6, 19) {real, imag} */,
  {32'h3f76faae, 32'hc06988b1} /* (14, 6, 18) {real, imag} */,
  {32'h40867710, 32'h3fcec8d7} /* (14, 6, 17) {real, imag} */,
  {32'h4091c794, 32'hbf9e9531} /* (14, 6, 16) {real, imag} */,
  {32'h40a86510, 32'h401c0bd7} /* (14, 6, 15) {real, imag} */,
  {32'hbe6c5f60, 32'h409afb68} /* (14, 6, 14) {real, imag} */,
  {32'hbfbc16de, 32'h403e1ec0} /* (14, 6, 13) {real, imag} */,
  {32'hc02cc9bc, 32'h3f1e53ee} /* (14, 6, 12) {real, imag} */,
  {32'hc06cd8df, 32'h4088855d} /* (14, 6, 11) {real, imag} */,
  {32'h4049c51f, 32'h3fe683cc} /* (14, 6, 10) {real, imag} */,
  {32'h40ef7d2c, 32'hc1071950} /* (14, 6, 9) {real, imag} */,
  {32'h40b81260, 32'hc11e46e9} /* (14, 6, 8) {real, imag} */,
  {32'h3ff19671, 32'hc0303ac6} /* (14, 6, 7) {real, imag} */,
  {32'h4044b0c8, 32'hbfb971a4} /* (14, 6, 6) {real, imag} */,
  {32'h4084acd8, 32'hc01b924e} /* (14, 6, 5) {real, imag} */,
  {32'h3e5a1dec, 32'hc0490f6b} /* (14, 6, 4) {real, imag} */,
  {32'h3f517eaa, 32'h3fba9ef6} /* (14, 6, 3) {real, imag} */,
  {32'h40b0c5f0, 32'h4028b648} /* (14, 6, 2) {real, imag} */,
  {32'h405d76a9, 32'hc008409d} /* (14, 6, 1) {real, imag} */,
  {32'h40274eba, 32'h3f242069} /* (14, 6, 0) {real, imag} */,
  {32'h40342a64, 32'h3f14cdcb} /* (14, 5, 31) {real, imag} */,
  {32'h408ddf0c, 32'h40a425e5} /* (14, 5, 30) {real, imag} */,
  {32'h40744f66, 32'hc00cedbf} /* (14, 5, 29) {real, imag} */,
  {32'h402999d3, 32'h4013135d} /* (14, 5, 28) {real, imag} */,
  {32'h40476351, 32'h41038c0f} /* (14, 5, 27) {real, imag} */,
  {32'h4098e413, 32'h40c4024d} /* (14, 5, 26) {real, imag} */,
  {32'h411b7e48, 32'h3ffe98ac} /* (14, 5, 25) {real, imag} */,
  {32'h4104ff61, 32'h4092e242} /* (14, 5, 24) {real, imag} */,
  {32'h40ea1f18, 32'h402054fc} /* (14, 5, 23) {real, imag} */,
  {32'h41183954, 32'h40200234} /* (14, 5, 22) {real, imag} */,
  {32'h40319eee, 32'h40ce241b} /* (14, 5, 21) {real, imag} */,
  {32'hc0137799, 32'h408fa540} /* (14, 5, 20) {real, imag} */,
  {32'hc00d4dc4, 32'hc01a0524} /* (14, 5, 19) {real, imag} */,
  {32'h40c0df27, 32'hc1112aa8} /* (14, 5, 18) {real, imag} */,
  {32'h3fbe22ca, 32'hc048390b} /* (14, 5, 17) {real, imag} */,
  {32'h3fe5ae4d, 32'h409e68d2} /* (14, 5, 16) {real, imag} */,
  {32'h40c22e78, 32'h3e913720} /* (14, 5, 15) {real, imag} */,
  {32'h40f901c6, 32'h3de83440} /* (14, 5, 14) {real, imag} */,
  {32'h3ff83b11, 32'h4007e57e} /* (14, 5, 13) {real, imag} */,
  {32'h40305809, 32'h409f2197} /* (14, 5, 12) {real, imag} */,
  {32'hbf8fa6ec, 32'hbf83930c} /* (14, 5, 11) {real, imag} */,
  {32'hbf53a120, 32'hbfdc86e2} /* (14, 5, 10) {real, imag} */,
  {32'hc0301a2c, 32'h40b9efa1} /* (14, 5, 9) {real, imag} */,
  {32'h4002e26d, 32'h410b91ea} /* (14, 5, 8) {real, imag} */,
  {32'hbf586fd0, 32'h40f49a22} /* (14, 5, 7) {real, imag} */,
  {32'hbf58caac, 32'h40909580} /* (14, 5, 6) {real, imag} */,
  {32'h3ff33d44, 32'h406e79c6} /* (14, 5, 5) {real, imag} */,
  {32'hbfba6ae0, 32'h3fbd0b2e} /* (14, 5, 4) {real, imag} */,
  {32'hc034440b, 32'h3fcdebb2} /* (14, 5, 3) {real, imag} */,
  {32'hbfdf6526, 32'h400f125c} /* (14, 5, 2) {real, imag} */,
  {32'h400a0102, 32'h40c319ba} /* (14, 5, 1) {real, imag} */,
  {32'h4020bfc8, 32'h40c01c40} /* (14, 5, 0) {real, imag} */,
  {32'h3f38dc86, 32'hc04e5c66} /* (14, 4, 31) {real, imag} */,
  {32'h3fbdbeee, 32'hbfdee68e} /* (14, 4, 30) {real, imag} */,
  {32'hbfc435ac, 32'h3f839b68} /* (14, 4, 29) {real, imag} */,
  {32'h3f83d89c, 32'h3fd1429e} /* (14, 4, 28) {real, imag} */,
  {32'h3ff4b570, 32'h409d4a87} /* (14, 4, 27) {real, imag} */,
  {32'h400c4b6d, 32'h4027d2c4} /* (14, 4, 26) {real, imag} */,
  {32'h3f6c07d2, 32'h3e90834c} /* (14, 4, 25) {real, imag} */,
  {32'h3e8d5b6f, 32'hbfb4a779} /* (14, 4, 24) {real, imag} */,
  {32'h3fa75af6, 32'h3fb55dc9} /* (14, 4, 23) {real, imag} */,
  {32'h403b8726, 32'h406038df} /* (14, 4, 22) {real, imag} */,
  {32'h40a52022, 32'h3ed1202e} /* (14, 4, 21) {real, imag} */,
  {32'h409c3348, 32'h3ee33ec8} /* (14, 4, 20) {real, imag} */,
  {32'h410fa0b8, 32'hc019f89e} /* (14, 4, 19) {real, imag} */,
  {32'h40cb8cd3, 32'hc01bdb16} /* (14, 4, 18) {real, imag} */,
  {32'h40c324a6, 32'h3e7510c0} /* (14, 4, 17) {real, imag} */,
  {32'h41009572, 32'h40556398} /* (14, 4, 16) {real, imag} */,
  {32'h3fb7ca18, 32'h3ec29630} /* (14, 4, 15) {real, imag} */,
  {32'h3f264fcc, 32'hbe1a9330} /* (14, 4, 14) {real, imag} */,
  {32'h40b270f7, 32'hbe8e9a04} /* (14, 4, 13) {real, imag} */,
  {32'h401647bd, 32'hc1094db6} /* (14, 4, 12) {real, imag} */,
  {32'h3fe13ee4, 32'hc09d6b9d} /* (14, 4, 11) {real, imag} */,
  {32'h3f4732a4, 32'h3f8eee19} /* (14, 4, 10) {real, imag} */,
  {32'hc008da6e, 32'hbfcce011} /* (14, 4, 9) {real, imag} */,
  {32'hbf7ac154, 32'h3e768030} /* (14, 4, 8) {real, imag} */,
  {32'hc00952c4, 32'h3efeec10} /* (14, 4, 7) {real, imag} */,
  {32'hc10552eb, 32'hc0da1211} /* (14, 4, 6) {real, imag} */,
  {32'hc1254aee, 32'hbfde359d} /* (14, 4, 5) {real, imag} */,
  {32'hc0ef151f, 32'hbfbe2632} /* (14, 4, 4) {real, imag} */,
  {32'hc0d5112c, 32'h3f938344} /* (14, 4, 3) {real, imag} */,
  {32'hc10d1a2a, 32'h3eeb4560} /* (14, 4, 2) {real, imag} */,
  {32'hc0900d80, 32'hc0f79f52} /* (14, 4, 1) {real, imag} */,
  {32'hbf0f75c9, 32'hc05ae599} /* (14, 4, 0) {real, imag} */,
  {32'h3f9ce910, 32'hc0a39362} /* (14, 3, 31) {real, imag} */,
  {32'hc0670ac4, 32'hc0cf841c} /* (14, 3, 30) {real, imag} */,
  {32'hbfbf7fcb, 32'hc0645074} /* (14, 3, 29) {real, imag} */,
  {32'h3f96c046, 32'h4090ebbc} /* (14, 3, 28) {real, imag} */,
  {32'hbdbeb960, 32'h409004ff} /* (14, 3, 27) {real, imag} */,
  {32'h409b0902, 32'h401d8ea5} /* (14, 3, 26) {real, imag} */,
  {32'h409ccc24, 32'hbe893e38} /* (14, 3, 25) {real, imag} */,
  {32'h4106ec55, 32'h40789ceb} /* (14, 3, 24) {real, imag} */,
  {32'h3ff6b100, 32'h405cbae3} /* (14, 3, 23) {real, imag} */,
  {32'hc0e5af46, 32'h403e4036} /* (14, 3, 22) {real, imag} */,
  {32'hc0a082d0, 32'h3f724dcc} /* (14, 3, 21) {real, imag} */,
  {32'h3f324cae, 32'h401dfd7d} /* (14, 3, 20) {real, imag} */,
  {32'h3dd3b610, 32'hbe97afaa} /* (14, 3, 19) {real, imag} */,
  {32'hc0366eb2, 32'h3f30e448} /* (14, 3, 18) {real, imag} */,
  {32'h4006cd2e, 32'h4018fb8a} /* (14, 3, 17) {real, imag} */,
  {32'h3fa19318, 32'h3fa27649} /* (14, 3, 16) {real, imag} */,
  {32'h4080f6cd, 32'h3e6cfd10} /* (14, 3, 15) {real, imag} */,
  {32'h40a5e661, 32'h4080f006} /* (14, 3, 14) {real, imag} */,
  {32'hbfb1d904, 32'h4072954f} /* (14, 3, 13) {real, imag} */,
  {32'hc02365f2, 32'hbf529874} /* (14, 3, 12) {real, imag} */,
  {32'hc06474a5, 32'h3fe02978} /* (14, 3, 11) {real, imag} */,
  {32'h3ef1c37e, 32'h4016f2d4} /* (14, 3, 10) {real, imag} */,
  {32'hc0cc9615, 32'h3be97800} /* (14, 3, 9) {real, imag} */,
  {32'hc06d4017, 32'hc0d80a53} /* (14, 3, 8) {real, imag} */,
  {32'hbf4aecb0, 32'hc0f8a827} /* (14, 3, 7) {real, imag} */,
  {32'h40040f78, 32'hc1356360} /* (14, 3, 6) {real, imag} */,
  {32'h4091aca5, 32'hc083ed09} /* (14, 3, 5) {real, imag} */,
  {32'h40b10676, 32'hc05c7c8e} /* (14, 3, 4) {real, imag} */,
  {32'h3d981600, 32'h3fda34eb} /* (14, 3, 3) {real, imag} */,
  {32'h4032615c, 32'h408326fe} /* (14, 3, 2) {real, imag} */,
  {32'h40622b7f, 32'hc01d36cd} /* (14, 3, 1) {real, imag} */,
  {32'h407e649e, 32'hc082c871} /* (14, 3, 0) {real, imag} */,
  {32'h40b0c715, 32'h3fdbae5c} /* (14, 2, 31) {real, imag} */,
  {32'h407c8e06, 32'hbef51f14} /* (14, 2, 30) {real, imag} */,
  {32'h40a83586, 32'h40ceda3d} /* (14, 2, 29) {real, imag} */,
  {32'h40dc5ba6, 32'h4090847d} /* (14, 2, 28) {real, imag} */,
  {32'h41005c59, 32'hc047de86} /* (14, 2, 27) {real, imag} */,
  {32'h410d2473, 32'hc02e0d70} /* (14, 2, 26) {real, imag} */,
  {32'h40bb2694, 32'h40081844} /* (14, 2, 25) {real, imag} */,
  {32'h40233bef, 32'h40500ee7} /* (14, 2, 24) {real, imag} */,
  {32'hc046f16e, 32'hc0a09ba8} /* (14, 2, 23) {real, imag} */,
  {32'h40a62172, 32'h400a0dfc} /* (14, 2, 22) {real, imag} */,
  {32'h41148b3d, 32'h40fa58c2} /* (14, 2, 21) {real, imag} */,
  {32'h3f19ce68, 32'h4112b4b2} /* (14, 2, 20) {real, imag} */,
  {32'hc0a47e7e, 32'h410f7bdc} /* (14, 2, 19) {real, imag} */,
  {32'hc0e85362, 32'h40add564} /* (14, 2, 18) {real, imag} */,
  {32'hc0d93291, 32'h3f8b3a9c} /* (14, 2, 17) {real, imag} */,
  {32'hc1478caf, 32'h402a2e14} /* (14, 2, 16) {real, imag} */,
  {32'hc0f05bce, 32'h410e35a8} /* (14, 2, 15) {real, imag} */,
  {32'hc0ef5d28, 32'hc08db7ed} /* (14, 2, 14) {real, imag} */,
  {32'hc0d2bb22, 32'hc071903c} /* (14, 2, 13) {real, imag} */,
  {32'hc0212492, 32'hc0acea64} /* (14, 2, 12) {real, imag} */,
  {32'hc0cf3457, 32'hc15850be} /* (14, 2, 11) {real, imag} */,
  {32'h3fe88804, 32'hc1086042} /* (14, 2, 10) {real, imag} */,
  {32'h4115ddf1, 32'hc0bdb00f} /* (14, 2, 9) {real, imag} */,
  {32'h4130d0ac, 32'hc08d8c50} /* (14, 2, 8) {real, imag} */,
  {32'h41762692, 32'hc0b70ff6} /* (14, 2, 7) {real, imag} */,
  {32'h417041cb, 32'hc08c732e} /* (14, 2, 6) {real, imag} */,
  {32'h40b1a212, 32'hbed132ae} /* (14, 2, 5) {real, imag} */,
  {32'h407bf323, 32'h400919c8} /* (14, 2, 4) {real, imag} */,
  {32'hc07f4554, 32'h402d2af1} /* (14, 2, 3) {real, imag} */,
  {32'h401c1bc7, 32'h4069a341} /* (14, 2, 2) {real, imag} */,
  {32'h412260b3, 32'h40f2067e} /* (14, 2, 1) {real, imag} */,
  {32'h41251e35, 32'h40cc060f} /* (14, 2, 0) {real, imag} */,
  {32'hc0b3601c, 32'hbf696da2} /* (14, 1, 31) {real, imag} */,
  {32'hc0c94b0d, 32'h4001fa7d} /* (14, 1, 30) {real, imag} */,
  {32'hc0598e36, 32'h40e327c8} /* (14, 1, 29) {real, imag} */,
  {32'hc12fe276, 32'h3e4257c2} /* (14, 1, 28) {real, imag} */,
  {32'hc18d1c5d, 32'hc01ab752} /* (14, 1, 27) {real, imag} */,
  {32'hc1a2600e, 32'hbf93c39d} /* (14, 1, 26) {real, imag} */,
  {32'hc1817dfa, 32'h4099b7b7} /* (14, 1, 25) {real, imag} */,
  {32'hc1801e80, 32'h3fb42360} /* (14, 1, 24) {real, imag} */,
  {32'hc15fd288, 32'h40cdb9f2} /* (14, 1, 23) {real, imag} */,
  {32'hc0d30420, 32'h40530c56} /* (14, 1, 22) {real, imag} */,
  {32'hc091ee1e, 32'hc0195303} /* (14, 1, 21) {real, imag} */,
  {32'hc00d5511, 32'h3fa645ba} /* (14, 1, 20) {real, imag} */,
  {32'h3fe22709, 32'h3f687440} /* (14, 1, 19) {real, imag} */,
  {32'h415adfaf, 32'h40399064} /* (14, 1, 18) {real, imag} */,
  {32'h41269a1e, 32'h3fdccea4} /* (14, 1, 17) {real, imag} */,
  {32'h402b0054, 32'h408a4bf4} /* (14, 1, 16) {real, imag} */,
  {32'h411ead88, 32'hc05ec9d8} /* (14, 1, 15) {real, imag} */,
  {32'h416d53ea, 32'hc03b4c08} /* (14, 1, 14) {real, imag} */,
  {32'h41669841, 32'hc01b7e19} /* (14, 1, 13) {real, imag} */,
  {32'h411804aa, 32'hc0027f7b} /* (14, 1, 12) {real, imag} */,
  {32'h4025a5ef, 32'hc0941798} /* (14, 1, 11) {real, imag} */,
  {32'h4038d1b6, 32'h3d4cb000} /* (14, 1, 10) {real, imag} */,
  {32'hc098c32a, 32'h409fdb39} /* (14, 1, 9) {real, imag} */,
  {32'hc142c806, 32'h3f139252} /* (14, 1, 8) {real, imag} */,
  {32'hc0a9603d, 32'hc08d13ef} /* (14, 1, 7) {real, imag} */,
  {32'h4041c6ec, 32'hbf8f16de} /* (14, 1, 6) {real, imag} */,
  {32'hc02ef038, 32'h3ffa186f} /* (14, 1, 5) {real, imag} */,
  {32'hc10d7ffc, 32'h40a45e8b} /* (14, 1, 4) {real, imag} */,
  {32'hc12c9e2a, 32'h3f5927ec} /* (14, 1, 3) {real, imag} */,
  {32'hc15eafb2, 32'hc09da974} /* (14, 1, 2) {real, imag} */,
  {32'hc1269a66, 32'hbf7fa218} /* (14, 1, 1) {real, imag} */,
  {32'hc0a6187f, 32'hc02d0645} /* (14, 1, 0) {real, imag} */,
  {32'hc098bd2c, 32'h40ad4398} /* (14, 0, 31) {real, imag} */,
  {32'hc08d8a12, 32'h40a24fc8} /* (14, 0, 30) {real, imag} */,
  {32'h3f8cb3d4, 32'hbf010668} /* (14, 0, 29) {real, imag} */,
  {32'hc08d6ef6, 32'h3bb62c00} /* (14, 0, 28) {real, imag} */,
  {32'hc121c4ca, 32'h4056d0b0} /* (14, 0, 27) {real, imag} */,
  {32'hc11ef575, 32'hbe237ee0} /* (14, 0, 26) {real, imag} */,
  {32'hc0c35cce, 32'hc0fe6c66} /* (14, 0, 25) {real, imag} */,
  {32'hc109798c, 32'hc0b3c3c0} /* (14, 0, 24) {real, imag} */,
  {32'hc0b781b8, 32'h409890ea} /* (14, 0, 23) {real, imag} */,
  {32'hc1024d50, 32'h40c4a8e3} /* (14, 0, 22) {real, imag} */,
  {32'hc1168537, 32'h3fd737c7} /* (14, 0, 21) {real, imag} */,
  {32'hc109f02a, 32'h3fe22a37} /* (14, 0, 20) {real, imag} */,
  {32'h4080e756, 32'h40d06d4a} /* (14, 0, 19) {real, imag} */,
  {32'h4100d0bd, 32'h408572a2} /* (14, 0, 18) {real, imag} */,
  {32'h401ff3c6, 32'h413428cf} /* (14, 0, 17) {real, imag} */,
  {32'hc01f2a42, 32'h40db476d} /* (14, 0, 16) {real, imag} */,
  {32'h40b251d5, 32'h3f933a58} /* (14, 0, 15) {real, imag} */,
  {32'h40efde32, 32'hbfaad4e4} /* (14, 0, 14) {real, imag} */,
  {32'h3fdd5a7b, 32'h408bc4ee} /* (14, 0, 13) {real, imag} */,
  {32'hbeffb1ea, 32'h3fb7b12a} /* (14, 0, 12) {real, imag} */,
  {32'h40664050, 32'hc0f2f4e6} /* (14, 0, 11) {real, imag} */,
  {32'hc02a294e, 32'hc0a86c65} /* (14, 0, 10) {real, imag} */,
  {32'hc08ad9e9, 32'h402a307b} /* (14, 0, 9) {real, imag} */,
  {32'h40438acc, 32'hbf9f485c} /* (14, 0, 8) {real, imag} */,
  {32'h40a30ad0, 32'h3f3c4170} /* (14, 0, 7) {real, imag} */,
  {32'h40b8554d, 32'h40f86115} /* (14, 0, 6) {real, imag} */,
  {32'hbff31a12, 32'h411487d9} /* (14, 0, 5) {real, imag} */,
  {32'hc0b6c8e7, 32'h3f103a80} /* (14, 0, 4) {real, imag} */,
  {32'hc02e1170, 32'hc004054b} /* (14, 0, 3) {real, imag} */,
  {32'h40247f40, 32'hc08deed0} /* (14, 0, 2) {real, imag} */,
  {32'h3fcc09cc, 32'hc0c8b91d} /* (14, 0, 1) {real, imag} */,
  {32'hbfef930a, 32'h400f50c9} /* (14, 0, 0) {real, imag} */,
  {32'hbf176ac4, 32'hc072520e} /* (13, 31, 31) {real, imag} */,
  {32'hbf25a48a, 32'h3cfbb300} /* (13, 31, 30) {real, imag} */,
  {32'hc0516d6d, 32'h405a04e0} /* (13, 31, 29) {real, imag} */,
  {32'h40dad0aa, 32'h3fca4808} /* (13, 31, 28) {real, imag} */,
  {32'h410994b5, 32'hc0b2ee0b} /* (13, 31, 27) {real, imag} */,
  {32'hc00ea19e, 32'hc10b8030} /* (13, 31, 26) {real, imag} */,
  {32'hbcf2b1f8, 32'hc0bc499a} /* (13, 31, 25) {real, imag} */,
  {32'h40620e3e, 32'hc08bce5b} /* (13, 31, 24) {real, imag} */,
  {32'hc04b1d8c, 32'h40723d7d} /* (13, 31, 23) {real, imag} */,
  {32'hbf495548, 32'h40eb7690} /* (13, 31, 22) {real, imag} */,
  {32'h4033187d, 32'h4089ba98} /* (13, 31, 21) {real, imag} */,
  {32'hbfd57a97, 32'h40c763c2} /* (13, 31, 20) {real, imag} */,
  {32'hc003b446, 32'h40bdcb34} /* (13, 31, 19) {real, imag} */,
  {32'hbfe282c4, 32'h4038029c} /* (13, 31, 18) {real, imag} */,
  {32'h3fe99e75, 32'hc013381a} /* (13, 31, 17) {real, imag} */,
  {32'h41359446, 32'hc0c51f09} /* (13, 31, 16) {real, imag} */,
  {32'h40f4b71b, 32'h4029a1af} /* (13, 31, 15) {real, imag} */,
  {32'hc0768df9, 32'h40c5890a} /* (13, 31, 14) {real, imag} */,
  {32'hbf111ea8, 32'h3b234a00} /* (13, 31, 13) {real, imag} */,
  {32'hc057ee1a, 32'hc031485b} /* (13, 31, 12) {real, imag} */,
  {32'hc0ae13a7, 32'hbf2e38e8} /* (13, 31, 11) {real, imag} */,
  {32'hc0ba92d0, 32'hbfd2f52c} /* (13, 31, 10) {real, imag} */,
  {32'h40380b4e, 32'h406d2ac5} /* (13, 31, 9) {real, imag} */,
  {32'h3eb4af20, 32'h410af86e} /* (13, 31, 8) {real, imag} */,
  {32'h406e534c, 32'h4091ffa8} /* (13, 31, 7) {real, imag} */,
  {32'h40de93d6, 32'hbd9e41d8} /* (13, 31, 6) {real, imag} */,
  {32'hc103c5e4, 32'hc09853aa} /* (13, 31, 5) {real, imag} */,
  {32'hc08db177, 32'hc00b76fa} /* (13, 31, 4) {real, imag} */,
  {32'h40aaa424, 32'h40f3589e} /* (13, 31, 3) {real, imag} */,
  {32'h4095276c, 32'h40016a14} /* (13, 31, 2) {real, imag} */,
  {32'h3fb167d8, 32'hbfb2b196} /* (13, 31, 1) {real, imag} */,
  {32'hbe5a4dd0, 32'hc05d1bdb} /* (13, 31, 0) {real, imag} */,
  {32'hc00a3b9d, 32'hbf57ae18} /* (13, 30, 31) {real, imag} */,
  {32'h3dfdf040, 32'hbf324ed8} /* (13, 30, 30) {real, imag} */,
  {32'h40604908, 32'hc0934bc1} /* (13, 30, 29) {real, imag} */,
  {32'hbed70600, 32'hc1337a88} /* (13, 30, 28) {real, imag} */,
  {32'hc10e546c, 32'hc11ff81f} /* (13, 30, 27) {real, imag} */,
  {32'hc12cbfb6, 32'h3fad727c} /* (13, 30, 26) {real, imag} */,
  {32'hc0c8343a, 32'h40a2561a} /* (13, 30, 25) {real, imag} */,
  {32'h3f0a3cd8, 32'h408977d6} /* (13, 30, 24) {real, imag} */,
  {32'h40ba0143, 32'hc080bfc0} /* (13, 30, 23) {real, imag} */,
  {32'hbfccc534, 32'hc0342708} /* (13, 30, 22) {real, imag} */,
  {32'hbf1a0020, 32'h40ee5047} /* (13, 30, 21) {real, imag} */,
  {32'h40a20754, 32'h40711288} /* (13, 30, 20) {real, imag} */,
  {32'h40e311f7, 32'hc0d8983e} /* (13, 30, 19) {real, imag} */,
  {32'h3f95afda, 32'hc08fdb47} /* (13, 30, 18) {real, imag} */,
  {32'h407c237c, 32'hbf744408} /* (13, 30, 17) {real, imag} */,
  {32'h3fd10fd7, 32'h40715777} /* (13, 30, 16) {real, imag} */,
  {32'hc088dba5, 32'h3b929800} /* (13, 30, 15) {real, imag} */,
  {32'hc0811730, 32'hbfc81ea8} /* (13, 30, 14) {real, imag} */,
  {32'hbf55adbc, 32'h402820ff} /* (13, 30, 13) {real, imag} */,
  {32'hc0c703fe, 32'h4113d670} /* (13, 30, 12) {real, imag} */,
  {32'hc0c89d86, 32'h402e1c64} /* (13, 30, 11) {real, imag} */,
  {32'hc0f7b93f, 32'h407f2266} /* (13, 30, 10) {real, imag} */,
  {32'hc0d08d34, 32'hbcc94c00} /* (13, 30, 9) {real, imag} */,
  {32'hc01b9c04, 32'hc02fc0d6} /* (13, 30, 8) {real, imag} */,
  {32'h3fd02073, 32'h403546c0} /* (13, 30, 7) {real, imag} */,
  {32'h40a363ee, 32'h3f92f718} /* (13, 30, 6) {real, imag} */,
  {32'hc04c64fe, 32'hbfe4f070} /* (13, 30, 5) {real, imag} */,
  {32'hbfd8fbea, 32'h3e6b2c00} /* (13, 30, 4) {real, imag} */,
  {32'h40ebe116, 32'hc0089db1} /* (13, 30, 3) {real, imag} */,
  {32'hc019d470, 32'hc0abfd64} /* (13, 30, 2) {real, imag} */,
  {32'hc092f4e9, 32'hc0e04e82} /* (13, 30, 1) {real, imag} */,
  {32'hbfadd526, 32'h3f0dde56} /* (13, 30, 0) {real, imag} */,
  {32'hbf77996d, 32'h40ab951c} /* (13, 29, 31) {real, imag} */,
  {32'h400f4968, 32'h40240982} /* (13, 29, 30) {real, imag} */,
  {32'h4042e056, 32'hc0600fcd} /* (13, 29, 29) {real, imag} */,
  {32'h40c8f3b2, 32'hbfda9801} /* (13, 29, 28) {real, imag} */,
  {32'h40b28fc6, 32'hbf2bbea0} /* (13, 29, 27) {real, imag} */,
  {32'hc04131ba, 32'h4093f5fb} /* (13, 29, 26) {real, imag} */,
  {32'hc0c3045e, 32'h40a38f9a} /* (13, 29, 25) {real, imag} */,
  {32'hc00beb65, 32'h41034628} /* (13, 29, 24) {real, imag} */,
  {32'h3f851ca8, 32'h4098f2f3} /* (13, 29, 23) {real, imag} */,
  {32'h40d68ad6, 32'h404510e8} /* (13, 29, 22) {real, imag} */,
  {32'h40c46153, 32'h4096b0f4} /* (13, 29, 21) {real, imag} */,
  {32'hbf7877b0, 32'hbfb1de78} /* (13, 29, 20) {real, imag} */,
  {32'h400c462c, 32'h40b9607e} /* (13, 29, 19) {real, imag} */,
  {32'hc0b48dea, 32'h3eea9a81} /* (13, 29, 18) {real, imag} */,
  {32'hbfcb1f61, 32'hc12ae22a} /* (13, 29, 17) {real, imag} */,
  {32'h405f0767, 32'hc047e40d} /* (13, 29, 16) {real, imag} */,
  {32'hbe948742, 32'hc037342e} /* (13, 29, 15) {real, imag} */,
  {32'hc052864d, 32'hc0b177bf} /* (13, 29, 14) {real, imag} */,
  {32'hc0c668cc, 32'hc108d4e4} /* (13, 29, 13) {real, imag} */,
  {32'hc09c98c5, 32'hc0d74eea} /* (13, 29, 12) {real, imag} */,
  {32'h3e71c318, 32'h40963610} /* (13, 29, 11) {real, imag} */,
  {32'h3f76b4a6, 32'h40a3eee8} /* (13, 29, 10) {real, imag} */,
  {32'hc0ddfd21, 32'h400ed650} /* (13, 29, 9) {real, imag} */,
  {32'hbfbb5f44, 32'hbf18b84d} /* (13, 29, 8) {real, imag} */,
  {32'h40dcdbc7, 32'hc06c28af} /* (13, 29, 7) {real, imag} */,
  {32'h409dc2e1, 32'h3fab05cf} /* (13, 29, 6) {real, imag} */,
  {32'h41069504, 32'h3fe91ba5} /* (13, 29, 5) {real, imag} */,
  {32'h401c93ba, 32'h4085d30b} /* (13, 29, 4) {real, imag} */,
  {32'hc04caa7e, 32'h407d3036} /* (13, 29, 3) {real, imag} */,
  {32'hc0d47464, 32'h41181540} /* (13, 29, 2) {real, imag} */,
  {32'h400cfe4f, 32'hc0120329} /* (13, 29, 1) {real, imag} */,
  {32'hbe302f40, 32'h3e168ad8} /* (13, 29, 0) {real, imag} */,
  {32'hbeaf9c5c, 32'hbfea5130} /* (13, 28, 31) {real, imag} */,
  {32'hc10c0128, 32'hc0a27f7a} /* (13, 28, 30) {real, imag} */,
  {32'hc0aedc80, 32'h40aeae64} /* (13, 28, 29) {real, imag} */,
  {32'h402a10d8, 32'h40a93269} /* (13, 28, 28) {real, imag} */,
  {32'hc03535b4, 32'hbe253aa0} /* (13, 28, 27) {real, imag} */,
  {32'h3f7bf91c, 32'h3f454454} /* (13, 28, 26) {real, imag} */,
  {32'h3f8a2369, 32'h3ead2a00} /* (13, 28, 25) {real, imag} */,
  {32'h3efe3244, 32'h40a857b4} /* (13, 28, 24) {real, imag} */,
  {32'h4155dde3, 32'hc049dfa6} /* (13, 28, 23) {real, imag} */,
  {32'h40960780, 32'hc0ced030} /* (13, 28, 22) {real, imag} */,
  {32'hc08bd31c, 32'hc0ad8846} /* (13, 28, 21) {real, imag} */,
  {32'h3dcc6ba0, 32'hc08b77b4} /* (13, 28, 20) {real, imag} */,
  {32'h40e3497f, 32'hc075f427} /* (13, 28, 19) {real, imag} */,
  {32'h40a51020, 32'hbe97eb18} /* (13, 28, 18) {real, imag} */,
  {32'h3f65f316, 32'h3ff4c3a6} /* (13, 28, 17) {real, imag} */,
  {32'hbf2ab1b4, 32'h40ae363a} /* (13, 28, 16) {real, imag} */,
  {32'hc0f5c81e, 32'h41098202} /* (13, 28, 15) {real, imag} */,
  {32'hc121e5c6, 32'h40d18566} /* (13, 28, 14) {real, imag} */,
  {32'hc1080610, 32'h40ee1f1d} /* (13, 28, 13) {real, imag} */,
  {32'hc0b84182, 32'h3f9d0e9c} /* (13, 28, 12) {real, imag} */,
  {32'hc144d323, 32'h3eef5038} /* (13, 28, 11) {real, imag} */,
  {32'hc11372ae, 32'h4061a0d6} /* (13, 28, 10) {real, imag} */,
  {32'hc071aec1, 32'h401bea66} /* (13, 28, 9) {real, imag} */,
  {32'h3f66e3f6, 32'hc0895e3a} /* (13, 28, 8) {real, imag} */,
  {32'hbfb9f0f5, 32'h3fb13c3e} /* (13, 28, 7) {real, imag} */,
  {32'hc0238434, 32'hc0101154} /* (13, 28, 6) {real, imag} */,
  {32'hc03a1420, 32'hc0f8e60c} /* (13, 28, 5) {real, imag} */,
  {32'h3ff02331, 32'hbeabbca0} /* (13, 28, 4) {real, imag} */,
  {32'h3f7a751c, 32'hc03ab8e0} /* (13, 28, 3) {real, imag} */,
  {32'h3e75a008, 32'hc08442c0} /* (13, 28, 2) {real, imag} */,
  {32'hc02c5de3, 32'h3fe1f408} /* (13, 28, 1) {real, imag} */,
  {32'hc04df8b8, 32'hc029ed10} /* (13, 28, 0) {real, imag} */,
  {32'hbfc5d729, 32'hbfa0ee40} /* (13, 27, 31) {real, imag} */,
  {32'hbe66f720, 32'h40278779} /* (13, 27, 30) {real, imag} */,
  {32'h409e254e, 32'h408d0554} /* (13, 27, 29) {real, imag} */,
  {32'hc06d71e4, 32'h40885764} /* (13, 27, 28) {real, imag} */,
  {32'h3fc97246, 32'hbf5e3ea8} /* (13, 27, 27) {real, imag} */,
  {32'h4103635e, 32'hc06e8584} /* (13, 27, 26) {real, imag} */,
  {32'h40565faa, 32'hc0b52b28} /* (13, 27, 25) {real, imag} */,
  {32'hc0020020, 32'hc03f0813} /* (13, 27, 24) {real, imag} */,
  {32'hbfb394ca, 32'hc082dd15} /* (13, 27, 23) {real, imag} */,
  {32'h40988bc2, 32'hbfa01b20} /* (13, 27, 22) {real, imag} */,
  {32'h405b4234, 32'h3fdc9bc8} /* (13, 27, 21) {real, imag} */,
  {32'h3b77f400, 32'hbfdca927} /* (13, 27, 20) {real, imag} */,
  {32'hbf8a88bc, 32'hbe584900} /* (13, 27, 19) {real, imag} */,
  {32'hbed0ab70, 32'h406e3eda} /* (13, 27, 18) {real, imag} */,
  {32'hbfacf9ea, 32'h403d737c} /* (13, 27, 17) {real, imag} */,
  {32'hc0b4e943, 32'h3fb67f9a} /* (13, 27, 16) {real, imag} */,
  {32'hc0a4ceec, 32'hc0ed8a54} /* (13, 27, 15) {real, imag} */,
  {32'hc10a82b0, 32'hc0fba09c} /* (13, 27, 14) {real, imag} */,
  {32'hc0a6a0e2, 32'h3d83d860} /* (13, 27, 13) {real, imag} */,
  {32'h3f350ed8, 32'h403f2b22} /* (13, 27, 12) {real, imag} */,
  {32'h40013036, 32'h40c4417a} /* (13, 27, 11) {real, imag} */,
  {32'h3fe07d34, 32'h4111f87d} /* (13, 27, 10) {real, imag} */,
  {32'hc0a0da4d, 32'h400ab0d0} /* (13, 27, 9) {real, imag} */,
  {32'hc110e298, 32'hc14d233a} /* (13, 27, 8) {real, imag} */,
  {32'hc0d3269c, 32'hc0ee966c} /* (13, 27, 7) {real, imag} */,
  {32'h40235880, 32'h404300fe} /* (13, 27, 6) {real, imag} */,
  {32'hc104f90c, 32'hbf3263d2} /* (13, 27, 5) {real, imag} */,
  {32'hc0e6af19, 32'hc053be2c} /* (13, 27, 4) {real, imag} */,
  {32'hbfad7028, 32'hbece7fae} /* (13, 27, 3) {real, imag} */,
  {32'h405bb887, 32'hbfbd940a} /* (13, 27, 2) {real, imag} */,
  {32'hbe872ff0, 32'hc0f7f28b} /* (13, 27, 1) {real, imag} */,
  {32'hc05450e0, 32'hbf87bcba} /* (13, 27, 0) {real, imag} */,
  {32'h3f59fa64, 32'h40243f48} /* (13, 26, 31) {real, imag} */,
  {32'h4028eba4, 32'h3e89c0c4} /* (13, 26, 30) {real, imag} */,
  {32'h4059d794, 32'h3f8809d0} /* (13, 26, 29) {real, imag} */,
  {32'hbf84398c, 32'hbf77cb24} /* (13, 26, 28) {real, imag} */,
  {32'h3f5454f6, 32'hc0f70614} /* (13, 26, 27) {real, imag} */,
  {32'h40900e36, 32'hc0531cf1} /* (13, 26, 26) {real, imag} */,
  {32'hbf8d7010, 32'hbf871e90} /* (13, 26, 25) {real, imag} */,
  {32'h4090a121, 32'hbe1fc060} /* (13, 26, 24) {real, imag} */,
  {32'hbf554420, 32'hbfcd0c63} /* (13, 26, 23) {real, imag} */,
  {32'hc08864b8, 32'h3eda8c50} /* (13, 26, 22) {real, imag} */,
  {32'hc095ba3e, 32'hbf82606c} /* (13, 26, 21) {real, imag} */,
  {32'h40092d96, 32'hc0818ab9} /* (13, 26, 20) {real, imag} */,
  {32'h40048078, 32'hbe97dd3e} /* (13, 26, 19) {real, imag} */,
  {32'hc05aa73e, 32'hc10bf982} /* (13, 26, 18) {real, imag} */,
  {32'hc10a5b92, 32'hc110a396} /* (13, 26, 17) {real, imag} */,
  {32'hc0d37558, 32'hc0a7f748} /* (13, 26, 16) {real, imag} */,
  {32'h3ea77344, 32'hbf4aca8b} /* (13, 26, 15) {real, imag} */,
  {32'hbfbeb913, 32'hc0b24230} /* (13, 26, 14) {real, imag} */,
  {32'hc0b5f6fc, 32'hc08aeb84} /* (13, 26, 13) {real, imag} */,
  {32'hc050a5af, 32'h3f8bcb3e} /* (13, 26, 12) {real, imag} */,
  {32'h3f73aff0, 32'hbfa5e5e4} /* (13, 26, 11) {real, imag} */,
  {32'hc0596ff2, 32'hc0a44ae9} /* (13, 26, 10) {real, imag} */,
  {32'hbcb56900, 32'hc0ff6b5b} /* (13, 26, 9) {real, imag} */,
  {32'h40ac654d, 32'hc0a8d5d1} /* (13, 26, 8) {real, imag} */,
  {32'h40146118, 32'hbfa95f88} /* (13, 26, 7) {real, imag} */,
  {32'hbf10c384, 32'hbf645e7c} /* (13, 26, 6) {real, imag} */,
  {32'h3d77cd00, 32'h40ab387a} /* (13, 26, 5) {real, imag} */,
  {32'hbf86be0c, 32'h3fe68e21} /* (13, 26, 4) {real, imag} */,
  {32'h4080a06e, 32'h3ff8255a} /* (13, 26, 3) {real, imag} */,
  {32'h40fa59ae, 32'h40903bca} /* (13, 26, 2) {real, imag} */,
  {32'h40a1519b, 32'h412d6450} /* (13, 26, 1) {real, imag} */,
  {32'h3e707862, 32'h406aac38} /* (13, 26, 0) {real, imag} */,
  {32'hc0e4923e, 32'hc0318096} /* (13, 25, 31) {real, imag} */,
  {32'hc08e7f43, 32'hc040b116} /* (13, 25, 30) {real, imag} */,
  {32'h40ff88ac, 32'hbf9b95fc} /* (13, 25, 29) {real, imag} */,
  {32'h3ffe1c44, 32'hbffb0a12} /* (13, 25, 28) {real, imag} */,
  {32'hc00d36da, 32'hbec6e2f4} /* (13, 25, 27) {real, imag} */,
  {32'h402e42fc, 32'hbecf8998} /* (13, 25, 26) {real, imag} */,
  {32'h4057d498, 32'hbf317402} /* (13, 25, 25) {real, imag} */,
  {32'h40c272f9, 32'hbf9b163c} /* (13, 25, 24) {real, imag} */,
  {32'h411005fa, 32'hc01bf6df} /* (13, 25, 23) {real, imag} */,
  {32'h40aaf134, 32'hc06ba868} /* (13, 25, 22) {real, imag} */,
  {32'hc09a599c, 32'h3f2f6c80} /* (13, 25, 21) {real, imag} */,
  {32'hc1057bd6, 32'h409be944} /* (13, 25, 20) {real, imag} */,
  {32'hc0a9bb77, 32'h4083bcd4} /* (13, 25, 19) {real, imag} */,
  {32'hbf70fd04, 32'hbf1e1502} /* (13, 25, 18) {real, imag} */,
  {32'h3fa65c4c, 32'hbf7a5c12} /* (13, 25, 17) {real, imag} */,
  {32'h3fe6c443, 32'hbf5b501c} /* (13, 25, 16) {real, imag} */,
  {32'h3ea3f4e0, 32'h40496d76} /* (13, 25, 15) {real, imag} */,
  {32'h3fd747a0, 32'hbeddc2d8} /* (13, 25, 14) {real, imag} */,
  {32'h409ee085, 32'hc039865b} /* (13, 25, 13) {real, imag} */,
  {32'h409b7a9a, 32'hc04ada58} /* (13, 25, 12) {real, imag} */,
  {32'h40806007, 32'hc06e06af} /* (13, 25, 11) {real, imag} */,
  {32'h40aefb94, 32'hc025cfd1} /* (13, 25, 10) {real, imag} */,
  {32'h3f627ebc, 32'hc121df5d} /* (13, 25, 9) {real, imag} */,
  {32'hbf8be400, 32'hc0ccb0c2} /* (13, 25, 8) {real, imag} */,
  {32'h3e841148, 32'h407b93a0} /* (13, 25, 7) {real, imag} */,
  {32'h3f853b02, 32'h40e83d30} /* (13, 25, 6) {real, imag} */,
  {32'h3fb8e5fe, 32'h407eeeb5} /* (13, 25, 5) {real, imag} */,
  {32'hbfed93ac, 32'h3f109220} /* (13, 25, 4) {real, imag} */,
  {32'hbfd01d88, 32'h4010a11b} /* (13, 25, 3) {real, imag} */,
  {32'hbfa8755f, 32'h404d3344} /* (13, 25, 2) {real, imag} */,
  {32'hc0c4674f, 32'h404764bb} /* (13, 25, 1) {real, imag} */,
  {32'hc04b7f2f, 32'h3f7ecf2d} /* (13, 25, 0) {real, imag} */,
  {32'hbf0b8ffc, 32'hc0181147} /* (13, 24, 31) {real, imag} */,
  {32'hc017c562, 32'hc05a264f} /* (13, 24, 30) {real, imag} */,
  {32'h3f32e3ea, 32'hc10579bc} /* (13, 24, 29) {real, imag} */,
  {32'h3fe72f11, 32'hc061afeb} /* (13, 24, 28) {real, imag} */,
  {32'hc08cafae, 32'hc019f1d2} /* (13, 24, 27) {real, imag} */,
  {32'hc075bda8, 32'h400b1006} /* (13, 24, 26) {real, imag} */,
  {32'h400f7cac, 32'h3fb4a34d} /* (13, 24, 25) {real, imag} */,
  {32'h4065c0a8, 32'hbdfa4d70} /* (13, 24, 24) {real, imag} */,
  {32'h40349a0d, 32'h408006c8} /* (13, 24, 23) {real, imag} */,
  {32'hc077a8fc, 32'h407f1b30} /* (13, 24, 22) {real, imag} */,
  {32'hc0242fb2, 32'h3f4a8834} /* (13, 24, 21) {real, imag} */,
  {32'h3e8a390c, 32'hc01d151f} /* (13, 24, 20) {real, imag} */,
  {32'hc05c5e23, 32'hbf225630} /* (13, 24, 19) {real, imag} */,
  {32'hbf1a01f0, 32'h401619f6} /* (13, 24, 18) {real, imag} */,
  {32'h402d7f92, 32'h3e7ef600} /* (13, 24, 17) {real, imag} */,
  {32'h403a401b, 32'h40895fbb} /* (13, 24, 16) {real, imag} */,
  {32'h3ff204a6, 32'hbf949f0f} /* (13, 24, 15) {real, imag} */,
  {32'hbedfe694, 32'hc083a62c} /* (13, 24, 14) {real, imag} */,
  {32'hbdfbbfd0, 32'hc0a2cf8a} /* (13, 24, 13) {real, imag} */,
  {32'h40681d42, 32'hc0242841} /* (13, 24, 12) {real, imag} */,
  {32'h3f812e18, 32'h40ada5a4} /* (13, 24, 11) {real, imag} */,
  {32'hbef0db00, 32'hbea2afc4} /* (13, 24, 10) {real, imag} */,
  {32'h3f9e3414, 32'hbe5d6508} /* (13, 24, 9) {real, imag} */,
  {32'h4042a8ba, 32'h3fa40806} /* (13, 24, 8) {real, imag} */,
  {32'h3f68fd68, 32'h4010ead4} /* (13, 24, 7) {real, imag} */,
  {32'h3ff733ae, 32'h3fe2355f} /* (13, 24, 6) {real, imag} */,
  {32'h406b6b64, 32'hbf54a94e} /* (13, 24, 5) {real, imag} */,
  {32'h3f052ed8, 32'hbffc88d4} /* (13, 24, 4) {real, imag} */,
  {32'h3ea43c14, 32'h3ed03308} /* (13, 24, 3) {real, imag} */,
  {32'hc00592ce, 32'h3fd792a0} /* (13, 24, 2) {real, imag} */,
  {32'hbff15038, 32'hbf7a1db0} /* (13, 24, 1) {real, imag} */,
  {32'hb9b9a000, 32'hc02f8ee4} /* (13, 24, 0) {real, imag} */,
  {32'h3ff0798b, 32'h3fd84f04} /* (13, 23, 31) {real, imag} */,
  {32'h3eba5390, 32'h407fde1e} /* (13, 23, 30) {real, imag} */,
  {32'hbfec023a, 32'h3fe905dc} /* (13, 23, 29) {real, imag} */,
  {32'hc10114fc, 32'h40118d78} /* (13, 23, 28) {real, imag} */,
  {32'h3e92b314, 32'h3f853fb4} /* (13, 23, 27) {real, imag} */,
  {32'hc0003d45, 32'hc07fdc9b} /* (13, 23, 26) {real, imag} */,
  {32'hc0b05f34, 32'h3fa2a323} /* (13, 23, 25) {real, imag} */,
  {32'hbf7f7340, 32'hbff0837a} /* (13, 23, 24) {real, imag} */,
  {32'h402f5ddf, 32'hbfda811a} /* (13, 23, 23) {real, imag} */,
  {32'h3fb8e97a, 32'hc0625682} /* (13, 23, 22) {real, imag} */,
  {32'hbfed4ffd, 32'hc01720b7} /* (13, 23, 21) {real, imag} */,
  {32'h3feab996, 32'h3fd9293a} /* (13, 23, 20) {real, imag} */,
  {32'h4021f22b, 32'h3fcc2a25} /* (13, 23, 19) {real, imag} */,
  {32'h4039f86c, 32'h3fb06e38} /* (13, 23, 18) {real, imag} */,
  {32'hbea3c3fe, 32'hc0b3e40e} /* (13, 23, 17) {real, imag} */,
  {32'h3f7fb99e, 32'hc0bd8978} /* (13, 23, 16) {real, imag} */,
  {32'h4081a81a, 32'hbefd0762} /* (13, 23, 15) {real, imag} */,
  {32'hbfe8a774, 32'h400b89b5} /* (13, 23, 14) {real, imag} */,
  {32'hc000f186, 32'h3f89db44} /* (13, 23, 13) {real, imag} */,
  {32'h3ff9d28d, 32'hc0915608} /* (13, 23, 12) {real, imag} */,
  {32'hbf9cbce2, 32'hc08e3c9a} /* (13, 23, 11) {real, imag} */,
  {32'hc07179f8, 32'hbfacbfde} /* (13, 23, 10) {real, imag} */,
  {32'hc06fb66f, 32'h4028fff2} /* (13, 23, 9) {real, imag} */,
  {32'hbf5239fc, 32'h408c6618} /* (13, 23, 8) {real, imag} */,
  {32'h3f841982, 32'h40c4cf54} /* (13, 23, 7) {real, imag} */,
  {32'hc0198be1, 32'h4008f81b} /* (13, 23, 6) {real, imag} */,
  {32'hbf1cbf0c, 32'h3f7226a8} /* (13, 23, 5) {real, imag} */,
  {32'h401c4243, 32'h4063e129} /* (13, 23, 4) {real, imag} */,
  {32'h4032de40, 32'h40b6c43b} /* (13, 23, 3) {real, imag} */,
  {32'h3e316890, 32'h40ecd84d} /* (13, 23, 2) {real, imag} */,
  {32'h3f366144, 32'h4064f964} /* (13, 23, 1) {real, imag} */,
  {32'h3fba7007, 32'hbf003239} /* (13, 23, 0) {real, imag} */,
  {32'h404d5a43, 32'hc0269290} /* (13, 22, 31) {real, imag} */,
  {32'h3f8244c2, 32'hbf93385b} /* (13, 22, 30) {real, imag} */,
  {32'hc06ee542, 32'hbf2f7a64} /* (13, 22, 29) {real, imag} */,
  {32'hbe24df88, 32'hbfa51784} /* (13, 22, 28) {real, imag} */,
  {32'hc04020a8, 32'h40bdd5be} /* (13, 22, 27) {real, imag} */,
  {32'hc07759d6, 32'h406e3db7} /* (13, 22, 26) {real, imag} */,
  {32'h400ac332, 32'hc023d814} /* (13, 22, 25) {real, imag} */,
  {32'h40229672, 32'hbfb04d65} /* (13, 22, 24) {real, imag} */,
  {32'hbf3f4570, 32'hc00dea35} /* (13, 22, 23) {real, imag} */,
  {32'h3dda0f30, 32'hc07501d0} /* (13, 22, 22) {real, imag} */,
  {32'h3fcf4864, 32'h3f08ef0e} /* (13, 22, 21) {real, imag} */,
  {32'h3f2ad0b8, 32'h40180990} /* (13, 22, 20) {real, imag} */,
  {32'h4032e567, 32'h3fc80e52} /* (13, 22, 19) {real, imag} */,
  {32'h3ecfdebc, 32'hc03b659e} /* (13, 22, 18) {real, imag} */,
  {32'h3dbb4fa0, 32'hc07e8ac0} /* (13, 22, 17) {real, imag} */,
  {32'h3efb21a0, 32'hbfcae974} /* (13, 22, 16) {real, imag} */,
  {32'hc02784da, 32'hbf3fe7d4} /* (13, 22, 15) {real, imag} */,
  {32'h3fdda218, 32'h3f1f0a4c} /* (13, 22, 14) {real, imag} */,
  {32'h403a755a, 32'hc017e319} /* (13, 22, 13) {real, imag} */,
  {32'h404d345d, 32'hbff88dcc} /* (13, 22, 12) {real, imag} */,
  {32'h402b9f1c, 32'hbf8205dd} /* (13, 22, 11) {real, imag} */,
  {32'h40777ee4, 32'hbf629daa} /* (13, 22, 10) {real, imag} */,
  {32'h406c962c, 32'hbff17a40} /* (13, 22, 9) {real, imag} */,
  {32'h40c05450, 32'hc02a5aab} /* (13, 22, 8) {real, imag} */,
  {32'h408e6798, 32'hbfbdac8c} /* (13, 22, 7) {real, imag} */,
  {32'hbff66779, 32'hbd814e90} /* (13, 22, 6) {real, imag} */,
  {32'hbef8bd7c, 32'h3f8ca4cb} /* (13, 22, 5) {real, imag} */,
  {32'hbf7787e0, 32'hbe1f1fda} /* (13, 22, 4) {real, imag} */,
  {32'h3fb8fe7a, 32'hc013e4c8} /* (13, 22, 3) {real, imag} */,
  {32'hbfc4724e, 32'hbfd71398} /* (13, 22, 2) {real, imag} */,
  {32'hbfc0d43c, 32'hbd48f9c0} /* (13, 22, 1) {real, imag} */,
  {32'hbf283358, 32'h3d9e1a68} /* (13, 22, 0) {real, imag} */,
  {32'hbf612eca, 32'h3fd95194} /* (13, 21, 31) {real, imag} */,
  {32'hc01860c8, 32'h4046b2dc} /* (13, 21, 30) {real, imag} */,
  {32'h3ea6e270, 32'h3fa87d02} /* (13, 21, 29) {real, imag} */,
  {32'hc01cbeeb, 32'hbfbbeb49} /* (13, 21, 28) {real, imag} */,
  {32'hc0d3899e, 32'hc0687cff} /* (13, 21, 27) {real, imag} */,
  {32'hc08c64de, 32'hc06f856a} /* (13, 21, 26) {real, imag} */,
  {32'hbff0fa1a, 32'hc0248316} /* (13, 21, 25) {real, imag} */,
  {32'h3fcc9a54, 32'hc05ad380} /* (13, 21, 24) {real, imag} */,
  {32'h4083bc48, 32'h3fc42174} /* (13, 21, 23) {real, imag} */,
  {32'h404bea90, 32'h400e112c} /* (13, 21, 22) {real, imag} */,
  {32'h3f6da69c, 32'h3d45ea48} /* (13, 21, 21) {real, imag} */,
  {32'hbfb24946, 32'h3f8c70c7} /* (13, 21, 20) {real, imag} */,
  {32'hbfe09b8e, 32'hbda539a0} /* (13, 21, 19) {real, imag} */,
  {32'h3fa43af3, 32'h405c83a0} /* (13, 21, 18) {real, imag} */,
  {32'h3fc6fea8, 32'h40541988} /* (13, 21, 17) {real, imag} */,
  {32'hbfdada9e, 32'hbeaedb8e} /* (13, 21, 16) {real, imag} */,
  {32'hc0489650, 32'hc06412ad} /* (13, 21, 15) {real, imag} */,
  {32'hbf94ff43, 32'hc000c81a} /* (13, 21, 14) {real, imag} */,
  {32'h3f4b13c0, 32'h3f93a117} /* (13, 21, 13) {real, imag} */,
  {32'h4050c19e, 32'h3f809a7c} /* (13, 21, 12) {real, imag} */,
  {32'h3ff428ba, 32'hc03a26cd} /* (13, 21, 11) {real, imag} */,
  {32'hbfe7eb8c, 32'hc0349886} /* (13, 21, 10) {real, imag} */,
  {32'hc0043200, 32'h3f93b060} /* (13, 21, 9) {real, imag} */,
  {32'hbea82db8, 32'h40809900} /* (13, 21, 8) {real, imag} */,
  {32'hbfc802ea, 32'hbfb8de5a} /* (13, 21, 7) {real, imag} */,
  {32'hbf3a40bc, 32'hc011cd03} /* (13, 21, 6) {real, imag} */,
  {32'h4039e1a4, 32'hc00e44c0} /* (13, 21, 5) {real, imag} */,
  {32'hbef36d8a, 32'hbf8626da} /* (13, 21, 4) {real, imag} */,
  {32'h3fbe2a7e, 32'h4002ac8c} /* (13, 21, 3) {real, imag} */,
  {32'h403da331, 32'h3fded9a4} /* (13, 21, 2) {real, imag} */,
  {32'h4030c5f0, 32'h3ff3d264} /* (13, 21, 1) {real, imag} */,
  {32'h401b7b1a, 32'h3f9ac2be} /* (13, 21, 0) {real, imag} */,
  {32'hbe06c1ec, 32'h3d8ed7f0} /* (13, 20, 31) {real, imag} */,
  {32'hbf4b8ee0, 32'hbdfdf530} /* (13, 20, 30) {real, imag} */,
  {32'hbf8e8b58, 32'h3f1d9440} /* (13, 20, 29) {real, imag} */,
  {32'hbe1d7394, 32'hbe9f8833} /* (13, 20, 28) {real, imag} */,
  {32'hbf3dc918, 32'hbfd26631} /* (13, 20, 27) {real, imag} */,
  {32'h3e178610, 32'hbf94e7a6} /* (13, 20, 26) {real, imag} */,
  {32'hbf56e658, 32'h3f0a5910} /* (13, 20, 25) {real, imag} */,
  {32'hc0096b0b, 32'h3f6a119f} /* (13, 20, 24) {real, imag} */,
  {32'hbe602df0, 32'h3f397413} /* (13, 20, 23) {real, imag} */,
  {32'h4080f3ed, 32'h3f6ec776} /* (13, 20, 22) {real, imag} */,
  {32'h4040eb0e, 32'h3f14fc0d} /* (13, 20, 21) {real, imag} */,
  {32'hbf90c287, 32'hbf9d78ae} /* (13, 20, 20) {real, imag} */,
  {32'hbf85d266, 32'hbfa18b58} /* (13, 20, 19) {real, imag} */,
  {32'hc00d1426, 32'h4022a09c} /* (13, 20, 18) {real, imag} */,
  {32'hbfc90c87, 32'h40875542} /* (13, 20, 17) {real, imag} */,
  {32'hbfa0b456, 32'h3ff6db54} /* (13, 20, 16) {real, imag} */,
  {32'hbfd6857b, 32'hbfa51739} /* (13, 20, 15) {real, imag} */,
  {32'hbe1f1f68, 32'hbfa781e7} /* (13, 20, 14) {real, imag} */,
  {32'h400468c8, 32'hbe3cfec8} /* (13, 20, 13) {real, imag} */,
  {32'h4058807c, 32'h4060ab16} /* (13, 20, 12) {real, imag} */,
  {32'h3ff19446, 32'h3ff3a547} /* (13, 20, 11) {real, imag} */,
  {32'h3fcbff24, 32'hbf70fa03} /* (13, 20, 10) {real, imag} */,
  {32'h3fda3160, 32'h3ee17b8c} /* (13, 20, 9) {real, imag} */,
  {32'h3f787fb6, 32'hbfad6998} /* (13, 20, 8) {real, imag} */,
  {32'hbfc12863, 32'hbf49abb4} /* (13, 20, 7) {real, imag} */,
  {32'hc04b9592, 32'h3fb693fe} /* (13, 20, 6) {real, imag} */,
  {32'hbf2dbc9e, 32'h3e0da890} /* (13, 20, 5) {real, imag} */,
  {32'hbd853898, 32'hbff8e111} /* (13, 20, 4) {real, imag} */,
  {32'hbf9f762f, 32'h3fe76b76} /* (13, 20, 3) {real, imag} */,
  {32'hbfbe6a65, 32'h3fced238} /* (13, 20, 2) {real, imag} */,
  {32'hc0080998, 32'h3ec01bbe} /* (13, 20, 1) {real, imag} */,
  {32'h3e8d6082, 32'h3e0a6f08} /* (13, 20, 0) {real, imag} */,
  {32'hbf90d3fd, 32'hbfc0313e} /* (13, 19, 31) {real, imag} */,
  {32'hbe3c4328, 32'h3bb71e00} /* (13, 19, 30) {real, imag} */,
  {32'h3f57f6d0, 32'h3f5a84f2} /* (13, 19, 29) {real, imag} */,
  {32'h3ded2470, 32'hbf6f198e} /* (13, 19, 28) {real, imag} */,
  {32'h3cc3b940, 32'hbec90e68} /* (13, 19, 27) {real, imag} */,
  {32'h3f9d4f8d, 32'hbfefae00} /* (13, 19, 26) {real, imag} */,
  {32'hbcab9f80, 32'hc0713420} /* (13, 19, 25) {real, imag} */,
  {32'hc001b4ca, 32'hbffe4887} /* (13, 19, 24) {real, imag} */,
  {32'hbf523d51, 32'hbf26d5e4} /* (13, 19, 23) {real, imag} */,
  {32'h3ed6809c, 32'h3daa7bd8} /* (13, 19, 22) {real, imag} */,
  {32'hbf409822, 32'h3fe6732a} /* (13, 19, 21) {real, imag} */,
  {32'hc0016ef0, 32'h3f602576} /* (13, 19, 20) {real, imag} */,
  {32'hc0469c2e, 32'h3f63d886} /* (13, 19, 19) {real, imag} */,
  {32'hbf97f288, 32'h3f8aefd6} /* (13, 19, 18) {real, imag} */,
  {32'h40077408, 32'hbf5f60c4} /* (13, 19, 17) {real, imag} */,
  {32'h3f1e0a80, 32'hbdd06350} /* (13, 19, 16) {real, imag} */,
  {32'h3e89ebe4, 32'h401497e7} /* (13, 19, 15) {real, imag} */,
  {32'hbfa9cb54, 32'h3fe454ca} /* (13, 19, 14) {real, imag} */,
  {32'h3db6aee0, 32'hbfb6a712} /* (13, 19, 13) {real, imag} */,
  {32'h3d7acb80, 32'hbfc5e7d2} /* (13, 19, 12) {real, imag} */,
  {32'h3f88ea89, 32'hbf2fc94e} /* (13, 19, 11) {real, imag} */,
  {32'hbf6c485e, 32'h3f75800d} /* (13, 19, 10) {real, imag} */,
  {32'hc00bfeec, 32'h3e9ca744} /* (13, 19, 9) {real, imag} */,
  {32'h3dbf2170, 32'h3c099740} /* (13, 19, 8) {real, imag} */,
  {32'hbf6d0123, 32'hbe66989c} /* (13, 19, 7) {real, imag} */,
  {32'hbfad03f3, 32'h3fd79b96} /* (13, 19, 6) {real, imag} */,
  {32'h3ece035c, 32'hbeb11008} /* (13, 19, 5) {real, imag} */,
  {32'h40151a52, 32'hbf69a6aa} /* (13, 19, 4) {real, imag} */,
  {32'h3f207e56, 32'hc0014010} /* (13, 19, 3) {real, imag} */,
  {32'hbdf1be38, 32'hc003f188} /* (13, 19, 2) {real, imag} */,
  {32'hbf433190, 32'hbfc5bba7} /* (13, 19, 1) {real, imag} */,
  {32'hbfe5daa6, 32'hc003919b} /* (13, 19, 0) {real, imag} */,
  {32'h3fb3e836, 32'hbd9d5750} /* (13, 18, 31) {real, imag} */,
  {32'h3f047248, 32'h3dcf1460} /* (13, 18, 30) {real, imag} */,
  {32'hbfe8ec24, 32'hbf163489} /* (13, 18, 29) {real, imag} */,
  {32'h3f9bd55c, 32'hbf2ee5fc} /* (13, 18, 28) {real, imag} */,
  {32'h4003c86e, 32'h3eb5bd40} /* (13, 18, 27) {real, imag} */,
  {32'h401e90ae, 32'h3fe808ee} /* (13, 18, 26) {real, imag} */,
  {32'h3fd1f324, 32'hbfc9dc5d} /* (13, 18, 25) {real, imag} */,
  {32'hbf224014, 32'hc00bf09a} /* (13, 18, 24) {real, imag} */,
  {32'hbf4b9a6c, 32'h3f25c154} /* (13, 18, 23) {real, imag} */,
  {32'hbcaf8a80, 32'h3f7edc30} /* (13, 18, 22) {real, imag} */,
  {32'hbf936d61, 32'hbf603f86} /* (13, 18, 21) {real, imag} */,
  {32'hbfc9cde8, 32'h3e0c2c4a} /* (13, 18, 20) {real, imag} */,
  {32'hbf5c2bd8, 32'hc009c8c2} /* (13, 18, 19) {real, imag} */,
  {32'h3f40bc08, 32'hbfb67c8c} /* (13, 18, 18) {real, imag} */,
  {32'h3faf126c, 32'h3f841d18} /* (13, 18, 17) {real, imag} */,
  {32'h3f16a354, 32'hbd28f080} /* (13, 18, 16) {real, imag} */,
  {32'h3ee5c9f0, 32'h3e2637c0} /* (13, 18, 15) {real, imag} */,
  {32'hbf75df3a, 32'h3f98fec4} /* (13, 18, 14) {real, imag} */,
  {32'hbfcd0abe, 32'hbd697920} /* (13, 18, 13) {real, imag} */,
  {32'hbf180558, 32'hbfd5f503} /* (13, 18, 12) {real, imag} */,
  {32'hbf22d996, 32'h3fc610a5} /* (13, 18, 11) {real, imag} */,
  {32'hbf45e56c, 32'h405d6664} /* (13, 18, 10) {real, imag} */,
  {32'h3f36e51a, 32'h3f3951f0} /* (13, 18, 9) {real, imag} */,
  {32'h404b5c00, 32'h3dce6010} /* (13, 18, 8) {real, imag} */,
  {32'hbec90218, 32'hbf092ff4} /* (13, 18, 7) {real, imag} */,
  {32'hbf682d3c, 32'hbfc6030f} /* (13, 18, 6) {real, imag} */,
  {32'h3fa0c498, 32'hc0729e9c} /* (13, 18, 5) {real, imag} */,
  {32'h3f9ba3d8, 32'hbf957808} /* (13, 18, 4) {real, imag} */,
  {32'hc02277cc, 32'h3deabe50} /* (13, 18, 3) {real, imag} */,
  {32'hc03c3be1, 32'hbf5ef645} /* (13, 18, 2) {real, imag} */,
  {32'hc00a8940, 32'hbff0441f} /* (13, 18, 1) {real, imag} */,
  {32'hbfaa43c0, 32'hbf80653c} /* (13, 18, 0) {real, imag} */,
  {32'hbf5f8d3d, 32'h3fabc7ec} /* (13, 17, 31) {real, imag} */,
  {32'hbf850a36, 32'h3fb7e91c} /* (13, 17, 30) {real, imag} */,
  {32'h3f141686, 32'h3fc5bf5a} /* (13, 17, 29) {real, imag} */,
  {32'h3f1eabee, 32'h3d986dc0} /* (13, 17, 28) {real, imag} */,
  {32'h3fc9922e, 32'hbf2eb6f8} /* (13, 17, 27) {real, imag} */,
  {32'h3fcaa34a, 32'hbfc3a615} /* (13, 17, 26) {real, imag} */,
  {32'h3f96117b, 32'hbf4ad636} /* (13, 17, 25) {real, imag} */,
  {32'h3f42b9aa, 32'hbe820f3c} /* (13, 17, 24) {real, imag} */,
  {32'h3f83820c, 32'h3dff19c8} /* (13, 17, 23) {real, imag} */,
  {32'hbec28df8, 32'h3e4fd110} /* (13, 17, 22) {real, imag} */,
  {32'hbfebde40, 32'h3ed24e2c} /* (13, 17, 21) {real, imag} */,
  {32'hbf1a6066, 32'h3f86e90f} /* (13, 17, 20) {real, imag} */,
  {32'h3ed0ba2c, 32'h3f6f8eb5} /* (13, 17, 19) {real, imag} */,
  {32'hbba3c000, 32'hbf176cea} /* (13, 17, 18) {real, imag} */,
  {32'hbdfd29d0, 32'hc0233510} /* (13, 17, 17) {real, imag} */,
  {32'h3f81fad4, 32'hc027ddb9} /* (13, 17, 16) {real, imag} */,
  {32'h3ffbfe0f, 32'hbfcb636c} /* (13, 17, 15) {real, imag} */,
  {32'h3fec72f6, 32'hbebe9719} /* (13, 17, 14) {real, imag} */,
  {32'h3f109f9c, 32'hbeb65b01} /* (13, 17, 13) {real, imag} */,
  {32'h3f654888, 32'h3ec0e1b0} /* (13, 17, 12) {real, imag} */,
  {32'hbd93c548, 32'h3f24ca14} /* (13, 17, 11) {real, imag} */,
  {32'hbf134f08, 32'h3f5d762c} /* (13, 17, 10) {real, imag} */,
  {32'h3daf5a08, 32'h3f9161e0} /* (13, 17, 9) {real, imag} */,
  {32'hbf2a8524, 32'h3f3f25f4} /* (13, 17, 8) {real, imag} */,
  {32'hbf1b8dd3, 32'h3edca48c} /* (13, 17, 7) {real, imag} */,
  {32'hbfc6929f, 32'h3f813a62} /* (13, 17, 6) {real, imag} */,
  {32'hbf92db82, 32'hbf2ce4b2} /* (13, 17, 5) {real, imag} */,
  {32'h3e5ac948, 32'hbebebc32} /* (13, 17, 4) {real, imag} */,
  {32'h3fc8bf91, 32'hc01f912f} /* (13, 17, 3) {real, imag} */,
  {32'h3e96b720, 32'hbf5cda48} /* (13, 17, 2) {real, imag} */,
  {32'hbdd79a00, 32'h3f385888} /* (13, 17, 1) {real, imag} */,
  {32'hbe111078, 32'h3f8f2ca8} /* (13, 17, 0) {real, imag} */,
  {32'hbf730bc8, 32'h3e5c9380} /* (13, 16, 31) {real, imag} */,
  {32'hbfd79480, 32'hbf7ddda4} /* (13, 16, 30) {real, imag} */,
  {32'hbfd6d4e6, 32'h3d7297a0} /* (13, 16, 29) {real, imag} */,
  {32'h3d17d000, 32'hbe95b770} /* (13, 16, 28) {real, imag} */,
  {32'h3f21f448, 32'hbe832f34} /* (13, 16, 27) {real, imag} */,
  {32'h3f1dfc7f, 32'hbe983acc} /* (13, 16, 26) {real, imag} */,
  {32'hbf12d6b4, 32'h3f306c28} /* (13, 16, 25) {real, imag} */,
  {32'hbfc60a7e, 32'h3f17e69e} /* (13, 16, 24) {real, imag} */,
  {32'hbf972c10, 32'h3f4c9480} /* (13, 16, 23) {real, imag} */,
  {32'hbd883d80, 32'h3f17bc44} /* (13, 16, 22) {real, imag} */,
  {32'h3fb7273c, 32'hbf4cca40} /* (13, 16, 21) {real, imag} */,
  {32'h3f875d26, 32'hbfd0d81e} /* (13, 16, 20) {real, imag} */,
  {32'h3faf6830, 32'h3ea774cc} /* (13, 16, 19) {real, imag} */,
  {32'h3fe031d4, 32'h3fbd9889} /* (13, 16, 18) {real, imag} */,
  {32'h3f9ee35c, 32'hbf2693c0} /* (13, 16, 17) {real, imag} */,
  {32'h3f1bc260, 32'hbfeee08c} /* (13, 16, 16) {real, imag} */,
  {32'h401521a9, 32'hbf268bca} /* (13, 16, 15) {real, imag} */,
  {32'h3f31edcf, 32'h3fb276cc} /* (13, 16, 14) {real, imag} */,
  {32'hbf951414, 32'hbec0bdd0} /* (13, 16, 13) {real, imag} */,
  {32'hbe24e290, 32'hbfb2dc5e} /* (13, 16, 12) {real, imag} */,
  {32'hbf4025d0, 32'hbed9f9d0} /* (13, 16, 11) {real, imag} */,
  {32'hbfdb1634, 32'hbf974515} /* (13, 16, 10) {real, imag} */,
  {32'hbfed5fa8, 32'hbf96ea53} /* (13, 16, 9) {real, imag} */,
  {32'hbf425f20, 32'hbf40f7c0} /* (13, 16, 8) {real, imag} */,
  {32'h3e470af0, 32'hbf2703ea} /* (13, 16, 7) {real, imag} */,
  {32'h3de54aa0, 32'hc02bb183} /* (13, 16, 6) {real, imag} */,
  {32'hbe683240, 32'h3fa5633c} /* (13, 16, 5) {real, imag} */,
  {32'hbe149230, 32'h3fbaf8c8} /* (13, 16, 4) {real, imag} */,
  {32'h3fd92332, 32'hbfb668c8} /* (13, 16, 3) {real, imag} */,
  {32'h402c4760, 32'hbee51966} /* (13, 16, 2) {real, imag} */,
  {32'h40501649, 32'hbdc2a540} /* (13, 16, 1) {real, imag} */,
  {32'h3f8b35b4, 32'h3f1c54c8} /* (13, 16, 0) {real, imag} */,
  {32'h3d9d7818, 32'hbe4476a0} /* (13, 15, 31) {real, imag} */,
  {32'h3eda8c88, 32'h3ec94cb0} /* (13, 15, 30) {real, imag} */,
  {32'hbeab1bcb, 32'h3d214600} /* (13, 15, 29) {real, imag} */,
  {32'hbf70f2f2, 32'hbfa3bcb4} /* (13, 15, 28) {real, imag} */,
  {32'hbfc3ef8a, 32'h3e6e51a0} /* (13, 15, 27) {real, imag} */,
  {32'h3f54bd6c, 32'hbf4fd1c2} /* (13, 15, 26) {real, imag} */,
  {32'h3f96c8b3, 32'hbfa6e141} /* (13, 15, 25) {real, imag} */,
  {32'h3fc2c06d, 32'hbcf007c0} /* (13, 15, 24) {real, imag} */,
  {32'h3eb6445e, 32'h3f03b0c3} /* (13, 15, 23) {real, imag} */,
  {32'hbede56c8, 32'h3e765cd0} /* (13, 15, 22) {real, imag} */,
  {32'hbd8848c0, 32'h3f93ebf5} /* (13, 15, 21) {real, imag} */,
  {32'h4030fa3a, 32'h3fbb9c95} /* (13, 15, 20) {real, imag} */,
  {32'h3fe11ab7, 32'h3dc9a0d8} /* (13, 15, 19) {real, imag} */,
  {32'h3f06c9b4, 32'hbf8a431b} /* (13, 15, 18) {real, imag} */,
  {32'h3f1d73ee, 32'h3f564fc0} /* (13, 15, 17) {real, imag} */,
  {32'h40005942, 32'hbe903f48} /* (13, 15, 16) {real, imag} */,
  {32'h400ac91c, 32'hbf931090} /* (13, 15, 15) {real, imag} */,
  {32'h3fad330e, 32'hbdb5f1e4} /* (13, 15, 14) {real, imag} */,
  {32'hbd30a840, 32'hbf1dc9ce} /* (13, 15, 13) {real, imag} */,
  {32'hbe851d70, 32'hbcd44680} /* (13, 15, 12) {real, imag} */,
  {32'hbf836edc, 32'h3e9aa9c8} /* (13, 15, 11) {real, imag} */,
  {32'hbf58e878, 32'h3fabdc0e} /* (13, 15, 10) {real, imag} */,
  {32'h3fd217ba, 32'h3fb575f8} /* (13, 15, 9) {real, imag} */,
  {32'h4003c866, 32'h3f93d352} /* (13, 15, 8) {real, imag} */,
  {32'h3fed8038, 32'h3ef7d674} /* (13, 15, 7) {real, imag} */,
  {32'h3fa558f5, 32'hbdcab758} /* (13, 15, 6) {real, imag} */,
  {32'h3ea10e18, 32'hbfa1f683} /* (13, 15, 5) {real, imag} */,
  {32'hbfcf22ad, 32'hbfcb997c} /* (13, 15, 4) {real, imag} */,
  {32'hbf5edbbe, 32'hbd467240} /* (13, 15, 3) {real, imag} */,
  {32'h3ec58688, 32'hbfe9fbb4} /* (13, 15, 2) {real, imag} */,
  {32'h3f3c7928, 32'hbfa3e0c0} /* (13, 15, 1) {real, imag} */,
  {32'h3ef003d4, 32'h3e85d09e} /* (13, 15, 0) {real, imag} */,
  {32'hbf320184, 32'hbeca9fcc} /* (13, 14, 31) {real, imag} */,
  {32'hbf82d534, 32'hbebef988} /* (13, 14, 30) {real, imag} */,
  {32'h3f9888e2, 32'hbe202d84} /* (13, 14, 29) {real, imag} */,
  {32'h3fc389f0, 32'h3fdf949a} /* (13, 14, 28) {real, imag} */,
  {32'h3e946974, 32'hbea9e7f0} /* (13, 14, 27) {real, imag} */,
  {32'h3f4fb2a8, 32'hbee968f0} /* (13, 14, 26) {real, imag} */,
  {32'h3ed85d32, 32'h3e8b78ac} /* (13, 14, 25) {real, imag} */,
  {32'h3ef51890, 32'hbfc33e25} /* (13, 14, 24) {real, imag} */,
  {32'h3fc12ada, 32'hc00fdfed} /* (13, 14, 23) {real, imag} */,
  {32'h3fa38336, 32'hbf5fb240} /* (13, 14, 22) {real, imag} */,
  {32'h3fb0f17f, 32'h3f7031da} /* (13, 14, 21) {real, imag} */,
  {32'h3f605248, 32'hbf49c4de} /* (13, 14, 20) {real, imag} */,
  {32'hbf00e6e4, 32'hc03ed926} /* (13, 14, 19) {real, imag} */,
  {32'h3ec636a7, 32'hbfa98b60} /* (13, 14, 18) {real, imag} */,
  {32'h3ef367d0, 32'hbffc1e2a} /* (13, 14, 17) {real, imag} */,
  {32'hbd51d2e8, 32'hbf9f4fb0} /* (13, 14, 16) {real, imag} */,
  {32'hbf0d4668, 32'hbfb0e264} /* (13, 14, 15) {real, imag} */,
  {32'h3faab613, 32'hbf34e530} /* (13, 14, 14) {real, imag} */,
  {32'h402032a9, 32'hbf5c60da} /* (13, 14, 13) {real, imag} */,
  {32'h40324bfa, 32'hbdb80870} /* (13, 14, 12) {real, imag} */,
  {32'h4041460c, 32'h3e97def4} /* (13, 14, 11) {real, imag} */,
  {32'h3e970068, 32'h3f9c0b88} /* (13, 14, 10) {real, imag} */,
  {32'h3cce7540, 32'h3f59af08} /* (13, 14, 9) {real, imag} */,
  {32'h3e524098, 32'h3e9693fc} /* (13, 14, 8) {real, imag} */,
  {32'hc000d3bc, 32'h3f43d9ec} /* (13, 14, 7) {real, imag} */,
  {32'hbfa293f2, 32'h3f92410f} /* (13, 14, 6) {real, imag} */,
  {32'hbf4e6c98, 32'hbf67b402} /* (13, 14, 5) {real, imag} */,
  {32'hbf161153, 32'hbfb89c9c} /* (13, 14, 4) {real, imag} */,
  {32'hbe60ba88, 32'hbf19eede} /* (13, 14, 3) {real, imag} */,
  {32'h3e9017b8, 32'h3eddd65a} /* (13, 14, 2) {real, imag} */,
  {32'h3f1ac0b2, 32'hbe3c6ca8} /* (13, 14, 1) {real, imag} */,
  {32'h3f6827f8, 32'hbfa35e30} /* (13, 14, 0) {real, imag} */,
  {32'h3f4cd8b4, 32'hc0335f41} /* (13, 13, 31) {real, imag} */,
  {32'h3f24c30e, 32'hc02c3f88} /* (13, 13, 30) {real, imag} */,
  {32'hbf50792c, 32'hbf899f83} /* (13, 13, 29) {real, imag} */,
  {32'hbfafb519, 32'h3f80379b} /* (13, 13, 28) {real, imag} */,
  {32'h3ea89d34, 32'h3fd34a7c} /* (13, 13, 27) {real, imag} */,
  {32'hbfa607c3, 32'h3f0e2738} /* (13, 13, 26) {real, imag} */,
  {32'hc07992e7, 32'hbffb6f91} /* (13, 13, 25) {real, imag} */,
  {32'hc048b8f2, 32'hbfceae51} /* (13, 13, 24) {real, imag} */,
  {32'hc00fdc03, 32'h3fbee54a} /* (13, 13, 23) {real, imag} */,
  {32'hbfaab6bf, 32'hbfefc7a0} /* (13, 13, 22) {real, imag} */,
  {32'hbf815ab5, 32'hc063d76f} /* (13, 13, 21) {real, imag} */,
  {32'hbfa3e940, 32'hbfff48a7} /* (13, 13, 20) {real, imag} */,
  {32'hbeb964c4, 32'hbfc7163d} /* (13, 13, 19) {real, imag} */,
  {32'h4008ac19, 32'hc016e6b7} /* (13, 13, 18) {real, imag} */,
  {32'h40832fc8, 32'hc00049f9} /* (13, 13, 17) {real, imag} */,
  {32'h40050d74, 32'hbf8427c7} /* (13, 13, 16) {real, imag} */,
  {32'hc054bc9e, 32'h3f690478} /* (13, 13, 15) {real, imag} */,
  {32'hc07018ac, 32'hbf66b138} /* (13, 13, 14) {real, imag} */,
  {32'h3ec814a8, 32'h3ee92f38} /* (13, 13, 13) {real, imag} */,
  {32'h3fae872a, 32'h3f40032c} /* (13, 13, 12) {real, imag} */,
  {32'hbfcfc787, 32'h400f572c} /* (13, 13, 11) {real, imag} */,
  {32'hbf08d60a, 32'h3f126c45} /* (13, 13, 10) {real, imag} */,
  {32'hc044e640, 32'hbfc48dfa} /* (13, 13, 9) {real, imag} */,
  {32'hc00f7012, 32'hbe6fcdcc} /* (13, 13, 8) {real, imag} */,
  {32'hbeae7c8a, 32'h3da24f18} /* (13, 13, 7) {real, imag} */,
  {32'h3fb1ff4b, 32'h3f62cd47} /* (13, 13, 6) {real, imag} */,
  {32'h40166d1c, 32'h3e6ce5a0} /* (13, 13, 5) {real, imag} */,
  {32'h3e44c8b0, 32'h3faf4b21} /* (13, 13, 4) {real, imag} */,
  {32'hc02224ba, 32'h4035cff8} /* (13, 13, 3) {real, imag} */,
  {32'hbf59f759, 32'h3fa67c20} /* (13, 13, 2) {real, imag} */,
  {32'h3edf5ae0, 32'h3f02f64a} /* (13, 13, 1) {real, imag} */,
  {32'hbe32eaa4, 32'hbfdf831c} /* (13, 13, 0) {real, imag} */,
  {32'hbfe30478, 32'h3f8d0d75} /* (13, 12, 31) {real, imag} */,
  {32'hbfbc4df0, 32'h3f28ae52} /* (13, 12, 30) {real, imag} */,
  {32'h3f854c50, 32'hbf85ed92} /* (13, 12, 29) {real, imag} */,
  {32'h3f0321fd, 32'hbe13a6e6} /* (13, 12, 28) {real, imag} */,
  {32'hbf33132c, 32'hbf25193a} /* (13, 12, 27) {real, imag} */,
  {32'h3f5a4404, 32'hbf3fbd9c} /* (13, 12, 26) {real, imag} */,
  {32'hbfe1c23a, 32'hbe9e9ea8} /* (13, 12, 25) {real, imag} */,
  {32'h3f5201a8, 32'hbedb7da2} /* (13, 12, 24) {real, imag} */,
  {32'h3fb9d77e, 32'hbf12d639} /* (13, 12, 23) {real, imag} */,
  {32'h3fb50200, 32'h3fa422cb} /* (13, 12, 22) {real, imag} */,
  {32'h3e51e638, 32'h3ee76a6a} /* (13, 12, 21) {real, imag} */,
  {32'hbf8b52ad, 32'hc01f4498} /* (13, 12, 20) {real, imag} */,
  {32'hbeaf1c28, 32'hbee7a84f} /* (13, 12, 19) {real, imag} */,
  {32'hbeb5c51a, 32'h3fb686cb} /* (13, 12, 18) {real, imag} */,
  {32'hc0264cfa, 32'h3fd613ce} /* (13, 12, 17) {real, imag} */,
  {32'hc09af590, 32'h3fdeee00} /* (13, 12, 16) {real, imag} */,
  {32'hc000e0c8, 32'hbf991bd3} /* (13, 12, 15) {real, imag} */,
  {32'h40071670, 32'h3fa0c923} /* (13, 12, 14) {real, imag} */,
  {32'h3fd1a45f, 32'h3fc19aff} /* (13, 12, 13) {real, imag} */,
  {32'hc026f230, 32'h3e030088} /* (13, 12, 12) {real, imag} */,
  {32'hc029918b, 32'hc01e3a6a} /* (13, 12, 11) {real, imag} */,
  {32'hc046e14a, 32'hc0385376} /* (13, 12, 10) {real, imag} */,
  {32'hbe47fd24, 32'hbfdf5a79} /* (13, 12, 9) {real, imag} */,
  {32'hbfdacde5, 32'h3e655b14} /* (13, 12, 8) {real, imag} */,
  {32'hc0358a62, 32'h4064e69f} /* (13, 12, 7) {real, imag} */,
  {32'hbf7459b8, 32'h40b3f9fa} /* (13, 12, 6) {real, imag} */,
  {32'h3f874a8b, 32'h408b2fec} /* (13, 12, 5) {real, imag} */,
  {32'h3f1fdd99, 32'h3ff988d5} /* (13, 12, 4) {real, imag} */,
  {32'h403212b4, 32'h3f906b56} /* (13, 12, 3) {real, imag} */,
  {32'h3f16876a, 32'hbe0f9b00} /* (13, 12, 2) {real, imag} */,
  {32'hbe43314c, 32'hbf230503} /* (13, 12, 1) {real, imag} */,
  {32'h3f8d7034, 32'hbecf76d4} /* (13, 12, 0) {real, imag} */,
  {32'hbe360888, 32'hbebf44a0} /* (13, 11, 31) {real, imag} */,
  {32'h406c0d40, 32'h40095aa2} /* (13, 11, 30) {real, imag} */,
  {32'h3e464020, 32'hbe115cf0} /* (13, 11, 29) {real, imag} */,
  {32'hc0493425, 32'hc099c5b3} /* (13, 11, 28) {real, imag} */,
  {32'hbfae9f16, 32'hbf8f8bea} /* (13, 11, 27) {real, imag} */,
  {32'hc03e19ff, 32'h3fbc387c} /* (13, 11, 26) {real, imag} */,
  {32'hbff3eefe, 32'h4091b613} /* (13, 11, 25) {real, imag} */,
  {32'h3ed8b888, 32'h401f3b38} /* (13, 11, 24) {real, imag} */,
  {32'h3dc92ba0, 32'h3db9ae58} /* (13, 11, 23) {real, imag} */,
  {32'hbfab0bb9, 32'h3ef81e8a} /* (13, 11, 22) {real, imag} */,
  {32'hbe965008, 32'h3ea230b7} /* (13, 11, 21) {real, imag} */,
  {32'hc0778649, 32'hbf1b5f5e} /* (13, 11, 20) {real, imag} */,
  {32'hc067acb5, 32'h3fa13266} /* (13, 11, 19) {real, imag} */,
  {32'hbf9521d9, 32'h40108964} /* (13, 11, 18) {real, imag} */,
  {32'hbf1d0360, 32'hbfc9dc58} /* (13, 11, 17) {real, imag} */,
  {32'h3f5c73d4, 32'h400a43dd} /* (13, 11, 16) {real, imag} */,
  {32'hbe6511d8, 32'h407142c7} /* (13, 11, 15) {real, imag} */,
  {32'hbd59f920, 32'h40085356} /* (13, 11, 14) {real, imag} */,
  {32'h408c8744, 32'h3f311f24} /* (13, 11, 13) {real, imag} */,
  {32'h403ef012, 32'h3ecbf90e} /* (13, 11, 12) {real, imag} */,
  {32'hbf471b3c, 32'h400320f5} /* (13, 11, 11) {real, imag} */,
  {32'h3ee40b48, 32'h40219062} /* (13, 11, 10) {real, imag} */,
  {32'h402bd830, 32'hc05d2a00} /* (13, 11, 9) {real, imag} */,
  {32'h3df891a0, 32'hc04d3ad5} /* (13, 11, 8) {real, imag} */,
  {32'hc02b448d, 32'hbf79de3c} /* (13, 11, 7) {real, imag} */,
  {32'hbfda88b8, 32'h3d98b820} /* (13, 11, 6) {real, imag} */,
  {32'h3ecb8bd0, 32'h4037e780} /* (13, 11, 5) {real, imag} */,
  {32'hbfbefaaa, 32'h40819952} /* (13, 11, 4) {real, imag} */,
  {32'h4019b4a1, 32'hbf1e08b3} /* (13, 11, 3) {real, imag} */,
  {32'h4093ea13, 32'hc0300d14} /* (13, 11, 2) {real, imag} */,
  {32'hbf56d65e, 32'hbf945e1c} /* (13, 11, 1) {real, imag} */,
  {32'hc02d774a, 32'hbf492806} /* (13, 11, 0) {real, imag} */,
  {32'hbedbaed8, 32'h3cbbb180} /* (13, 10, 31) {real, imag} */,
  {32'h3d9a3680, 32'hbffb5839} /* (13, 10, 30) {real, imag} */,
  {32'hbfab9625, 32'hc0427adb} /* (13, 10, 29) {real, imag} */,
  {32'h3fcccc09, 32'hc042edfa} /* (13, 10, 28) {real, imag} */,
  {32'h40903efe, 32'h4001a03d} /* (13, 10, 27) {real, imag} */,
  {32'h3f5fa582, 32'h40678bf5} /* (13, 10, 26) {real, imag} */,
  {32'h3f5b5dd8, 32'hbf7774b2} /* (13, 10, 25) {real, imag} */,
  {32'h400f1ae8, 32'hbf738d1a} /* (13, 10, 24) {real, imag} */,
  {32'hbfa22996, 32'hbfb2563c} /* (13, 10, 23) {real, imag} */,
  {32'hc05c6cf2, 32'hc0a9096a} /* (13, 10, 22) {real, imag} */,
  {32'hc0621986, 32'h3f4233f8} /* (13, 10, 21) {real, imag} */,
  {32'h400905be, 32'h3f94d721} /* (13, 10, 20) {real, imag} */,
  {32'h408e2f7c, 32'hbfbdb926} /* (13, 10, 19) {real, imag} */,
  {32'h3f4c794e, 32'h3fb8630c} /* (13, 10, 18) {real, imag} */,
  {32'hc0595d1e, 32'hbf432370} /* (13, 10, 17) {real, imag} */,
  {32'hc0cb602a, 32'hc004235e} /* (13, 10, 16) {real, imag} */,
  {32'hbfd3fe9d, 32'hc09f4c32} /* (13, 10, 15) {real, imag} */,
  {32'hbecaadf8, 32'hc04d20c7} /* (13, 10, 14) {real, imag} */,
  {32'hbdad98d0, 32'hbe213990} /* (13, 10, 13) {real, imag} */,
  {32'h40eb8146, 32'h3fa26fac} /* (13, 10, 12) {real, imag} */,
  {32'h4043f0fc, 32'h3ff92a0d} /* (13, 10, 11) {real, imag} */,
  {32'h40674194, 32'hc006f054} /* (13, 10, 10) {real, imag} */,
  {32'h3fd363a8, 32'hc0b32bfe} /* (13, 10, 9) {real, imag} */,
  {32'hbee3c368, 32'hc114e5d4} /* (13, 10, 8) {real, imag} */,
  {32'hbdce44a0, 32'hc108c0f2} /* (13, 10, 7) {real, imag} */,
  {32'h4077ecc6, 32'hbf630fc6} /* (13, 10, 6) {real, imag} */,
  {32'h40711af8, 32'h405176fe} /* (13, 10, 5) {real, imag} */,
  {32'h4091685e, 32'h3ef7a9df} /* (13, 10, 4) {real, imag} */,
  {32'h3fd0a13e, 32'h3e14e940} /* (13, 10, 3) {real, imag} */,
  {32'hc0623917, 32'h3f052228} /* (13, 10, 2) {real, imag} */,
  {32'hc02a082a, 32'hbf91de96} /* (13, 10, 1) {real, imag} */,
  {32'h3cfcb970, 32'hbfe1cf30} /* (13, 10, 0) {real, imag} */,
  {32'hc048b39c, 32'h3fc7ff70} /* (13, 9, 31) {real, imag} */,
  {32'hc076a9bc, 32'hbfbe0cbf} /* (13, 9, 30) {real, imag} */,
  {32'h3ea39808, 32'hc09c94d9} /* (13, 9, 29) {real, imag} */,
  {32'h3ff922e4, 32'hc0134364} /* (13, 9, 28) {real, imag} */,
  {32'h3f83c6eb, 32'hc0a1da2f} /* (13, 9, 27) {real, imag} */,
  {32'h405594ef, 32'h3fbdd76a} /* (13, 9, 26) {real, imag} */,
  {32'h401e3a80, 32'h3fe50529} /* (13, 9, 25) {real, imag} */,
  {32'h40f7693a, 32'hc09f0ee6} /* (13, 9, 24) {real, imag} */,
  {32'h409bb314, 32'hbfe792b2} /* (13, 9, 23) {real, imag} */,
  {32'hc017aa9f, 32'hbdc6b1f0} /* (13, 9, 22) {real, imag} */,
  {32'hbfd3639d, 32'hc029ef7d} /* (13, 9, 21) {real, imag} */,
  {32'hbfeed586, 32'hbe822496} /* (13, 9, 20) {real, imag} */,
  {32'hc084eaac, 32'h3fd8fb63} /* (13, 9, 19) {real, imag} */,
  {32'hbfe54b5b, 32'h3f125383} /* (13, 9, 18) {real, imag} */,
  {32'hbf21f53f, 32'h400336a5} /* (13, 9, 17) {real, imag} */,
  {32'hc05b56f0, 32'hbfb5cc7e} /* (13, 9, 16) {real, imag} */,
  {32'hbc868e80, 32'hbf4e33d5} /* (13, 9, 15) {real, imag} */,
  {32'h3f2f4895, 32'hc00d0685} /* (13, 9, 14) {real, imag} */,
  {32'h3dd0e9c0, 32'h40836b8c} /* (13, 9, 13) {real, imag} */,
  {32'h3eb7fa14, 32'h4106fa88} /* (13, 9, 12) {real, imag} */,
  {32'h3e8551de, 32'h40d06c08} /* (13, 9, 11) {real, imag} */,
  {32'hc0285c68, 32'h40bce514} /* (13, 9, 10) {real, imag} */,
  {32'hc0be3506, 32'h40b77f6f} /* (13, 9, 9) {real, imag} */,
  {32'hbebba250, 32'h3d81b000} /* (13, 9, 8) {real, imag} */,
  {32'hbfb1e55a, 32'h3fcd4d8e} /* (13, 9, 7) {real, imag} */,
  {32'hc0bceef4, 32'h405fe4f5} /* (13, 9, 6) {real, imag} */,
  {32'hc0d0ed62, 32'h3f960484} /* (13, 9, 5) {real, imag} */,
  {32'h401e1b6d, 32'hc09bd680} /* (13, 9, 4) {real, imag} */,
  {32'h4104f9bc, 32'hc0d932f5} /* (13, 9, 3) {real, imag} */,
  {32'h3f79974c, 32'hbf9f9e24} /* (13, 9, 2) {real, imag} */,
  {32'hc0a127b0, 32'hbed2a50c} /* (13, 9, 1) {real, imag} */,
  {32'hc07deb46, 32'hbf712ae1} /* (13, 9, 0) {real, imag} */,
  {32'h408ef092, 32'h401ce60b} /* (13, 8, 31) {real, imag} */,
  {32'h408af17d, 32'h40b2812e} /* (13, 8, 30) {real, imag} */,
  {32'h405704da, 32'h3ed2e718} /* (13, 8, 29) {real, imag} */,
  {32'h3ea7fb6c, 32'hc082bd14} /* (13, 8, 28) {real, imag} */,
  {32'hbf03750c, 32'hbc0f7f80} /* (13, 8, 27) {real, imag} */,
  {32'hbf93646c, 32'hbfe2fd02} /* (13, 8, 26) {real, imag} */,
  {32'hbf2bf1a3, 32'hbfcf8543} /* (13, 8, 25) {real, imag} */,
  {32'h409cd3ea, 32'h4005168a} /* (13, 8, 24) {real, imag} */,
  {32'h404cefcd, 32'hc038249d} /* (13, 8, 23) {real, imag} */,
  {32'h401d79fc, 32'hc01e9bea} /* (13, 8, 22) {real, imag} */,
  {32'h40af6eff, 32'h3f9b7116} /* (13, 8, 21) {real, imag} */,
  {32'h40251960, 32'h40862aea} /* (13, 8, 20) {real, imag} */,
  {32'h3f9aea4e, 32'h40bd8cc0} /* (13, 8, 19) {real, imag} */,
  {32'hc062fe24, 32'h408c4d3d} /* (13, 8, 18) {real, imag} */,
  {32'h40184590, 32'hbf22c7f0} /* (13, 8, 17) {real, imag} */,
  {32'h406ae96d, 32'hbfa3f174} /* (13, 8, 16) {real, imag} */,
  {32'hc06e7821, 32'hc01eb814} /* (13, 8, 15) {real, imag} */,
  {32'hc01548d6, 32'hc001b851} /* (13, 8, 14) {real, imag} */,
  {32'hbf92f687, 32'hc014fd41} /* (13, 8, 13) {real, imag} */,
  {32'hc09646cb, 32'hc101371b} /* (13, 8, 12) {real, imag} */,
  {32'hc08cc2ec, 32'hc0a032a8} /* (13, 8, 11) {real, imag} */,
  {32'h404b8736, 32'hbf8a8ca1} /* (13, 8, 10) {real, imag} */,
  {32'h3fbc83b8, 32'h3d04ff60} /* (13, 8, 9) {real, imag} */,
  {32'h3f02a258, 32'h3fa5ac16} /* (13, 8, 8) {real, imag} */,
  {32'h41039f56, 32'h3ff2be95} /* (13, 8, 7) {real, imag} */,
  {32'h4106b79e, 32'h404e9870} /* (13, 8, 6) {real, imag} */,
  {32'h402b58f0, 32'h4007c2de} /* (13, 8, 5) {real, imag} */,
  {32'h40629588, 32'hbf842496} /* (13, 8, 4) {real, imag} */,
  {32'hbf8d48b5, 32'hc0782e61} /* (13, 8, 3) {real, imag} */,
  {32'hbffb234c, 32'hc0b9a542} /* (13, 8, 2) {real, imag} */,
  {32'h3f4489b0, 32'hc0ae4d80} /* (13, 8, 1) {real, imag} */,
  {32'h3fc1bb46, 32'hc04f3160} /* (13, 8, 0) {real, imag} */,
  {32'h3e044ab0, 32'hc045f124} /* (13, 7, 31) {real, imag} */,
  {32'h3ffc63a8, 32'hbf52dc56} /* (13, 7, 30) {real, imag} */,
  {32'h3fde5a7a, 32'h402b20fb} /* (13, 7, 29) {real, imag} */,
  {32'h406e96de, 32'h405b0877} /* (13, 7, 28) {real, imag} */,
  {32'hbe8ec5a4, 32'hc027e0b6} /* (13, 7, 27) {real, imag} */,
  {32'hbeede4cc, 32'hbf38ad78} /* (13, 7, 26) {real, imag} */,
  {32'h40766ad0, 32'h4039a70a} /* (13, 7, 25) {real, imag} */,
  {32'h41018eda, 32'hbfa3beb4} /* (13, 7, 24) {real, imag} */,
  {32'h3f28d0e0, 32'hc0aed4ae} /* (13, 7, 23) {real, imag} */,
  {32'hc0b598ee, 32'hbffd018d} /* (13, 7, 22) {real, imag} */,
  {32'hbff1adee, 32'hc04b717a} /* (13, 7, 21) {real, imag} */,
  {32'hc0923120, 32'h3f7191b4} /* (13, 7, 20) {real, imag} */,
  {32'hc0be8d91, 32'h3e4c3b38} /* (13, 7, 19) {real, imag} */,
  {32'hc050f5b3, 32'hc079b652} /* (13, 7, 18) {real, imag} */,
  {32'hc0b4a921, 32'hc086f7b9} /* (13, 7, 17) {real, imag} */,
  {32'hc02ad956, 32'hc009f039} /* (13, 7, 16) {real, imag} */,
  {32'hc04f69f8, 32'h3fe930e1} /* (13, 7, 15) {real, imag} */,
  {32'hc0827704, 32'h4024fe8f} /* (13, 7, 14) {real, imag} */,
  {32'hc0be3fdd, 32'h3f07848c} /* (13, 7, 13) {real, imag} */,
  {32'hc099a06c, 32'h3e4be400} /* (13, 7, 12) {real, imag} */,
  {32'hc082387b, 32'h40a3dc73} /* (13, 7, 11) {real, imag} */,
  {32'h40909804, 32'h3fb6d4fa} /* (13, 7, 10) {real, imag} */,
  {32'h408918b2, 32'hc0768bbc} /* (13, 7, 9) {real, imag} */,
  {32'hc0d51644, 32'h3eb6a2a0} /* (13, 7, 8) {real, imag} */,
  {32'hc092276a, 32'hbef073b4} /* (13, 7, 7) {real, imag} */,
  {32'h40832ab2, 32'h403cee67} /* (13, 7, 6) {real, imag} */,
  {32'h3f9a39e6, 32'hc02601d3} /* (13, 7, 5) {real, imag} */,
  {32'hbf68f2e5, 32'hc0cb6749} /* (13, 7, 4) {real, imag} */,
  {32'hc05b5a5c, 32'hbfb21c0b} /* (13, 7, 3) {real, imag} */,
  {32'hc08e4c91, 32'h3f4bdaa0} /* (13, 7, 2) {real, imag} */,
  {32'hc0980bfd, 32'h3f64ecd4} /* (13, 7, 1) {real, imag} */,
  {32'hbfd95b3a, 32'hbfb03952} /* (13, 7, 0) {real, imag} */,
  {32'h403cb38f, 32'hbf111294} /* (13, 6, 31) {real, imag} */,
  {32'h3fe89531, 32'h3e755278} /* (13, 6, 30) {real, imag} */,
  {32'hc0cee81c, 32'hbf8ef344} /* (13, 6, 29) {real, imag} */,
  {32'hc1006d52, 32'hc049ae8f} /* (13, 6, 28) {real, imag} */,
  {32'hbf193c7a, 32'h3fe2f922} /* (13, 6, 27) {real, imag} */,
  {32'h3fe7ebf2, 32'hc011a89b} /* (13, 6, 26) {real, imag} */,
  {32'h40677de8, 32'hc0fe6b04} /* (13, 6, 25) {real, imag} */,
  {32'hc08ca1c7, 32'hc0abb74b} /* (13, 6, 24) {real, imag} */,
  {32'hc0b26e7e, 32'h402dacaa} /* (13, 6, 23) {real, imag} */,
  {32'hbfcbdcbf, 32'h40b732f3} /* (13, 6, 22) {real, imag} */,
  {32'h3d22ac40, 32'hbfc23408} /* (13, 6, 21) {real, imag} */,
  {32'h4104e626, 32'h3eda0570} /* (13, 6, 20) {real, imag} */,
  {32'h40ef05d4, 32'h3f7f57e9} /* (13, 6, 19) {real, imag} */,
  {32'h41227638, 32'h40af606a} /* (13, 6, 18) {real, imag} */,
  {32'h3f3f5268, 32'h40cef489} /* (13, 6, 17) {real, imag} */,
  {32'hbfebbf00, 32'hbfb06ed8} /* (13, 6, 16) {real, imag} */,
  {32'h3fd7bff3, 32'h3f37c02f} /* (13, 6, 15) {real, imag} */,
  {32'h40a29e5f, 32'h403b5ec8} /* (13, 6, 14) {real, imag} */,
  {32'hbfdb6121, 32'hc067e0f5} /* (13, 6, 13) {real, imag} */,
  {32'hc09724b4, 32'hc08c3304} /* (13, 6, 12) {real, imag} */,
  {32'h409ebe62, 32'hc0bd47cb} /* (13, 6, 11) {real, imag} */,
  {32'h404e94b6, 32'h3fa35f6c} /* (13, 6, 10) {real, imag} */,
  {32'hc0880e09, 32'h407f370e} /* (13, 6, 9) {real, imag} */,
  {32'hc0472dfe, 32'h40454766} /* (13, 6, 8) {real, imag} */,
  {32'h406971ae, 32'h402de260} /* (13, 6, 7) {real, imag} */,
  {32'h3f093b74, 32'h40f247dc} /* (13, 6, 6) {real, imag} */,
  {32'h408dacb2, 32'h40edc19c} /* (13, 6, 5) {real, imag} */,
  {32'h407a52ca, 32'hc013f13e} /* (13, 6, 4) {real, imag} */,
  {32'h40dd623c, 32'h3fe46cfe} /* (13, 6, 3) {real, imag} */,
  {32'hbea03918, 32'h40df872e} /* (13, 6, 2) {real, imag} */,
  {32'hc06af761, 32'h40491580} /* (13, 6, 1) {real, imag} */,
  {32'hbf37ff12, 32'hbfc3fd4d} /* (13, 6, 0) {real, imag} */,
  {32'h409fb883, 32'hc0c17b23} /* (13, 5, 31) {real, imag} */,
  {32'h411584be, 32'hc032856f} /* (13, 5, 30) {real, imag} */,
  {32'h40217e93, 32'hc05f6dd0} /* (13, 5, 29) {real, imag} */,
  {32'h40e04016, 32'h402f5f76} /* (13, 5, 28) {real, imag} */,
  {32'h40baabd6, 32'h3ed54850} /* (13, 5, 27) {real, imag} */,
  {32'h3fc8cd3c, 32'h409c47ba} /* (13, 5, 26) {real, imag} */,
  {32'h40b606e1, 32'h4086b69a} /* (13, 5, 25) {real, imag} */,
  {32'h3f806512, 32'h40425cdd} /* (13, 5, 24) {real, imag} */,
  {32'hc0c596ba, 32'h3f80f51f} /* (13, 5, 23) {real, imag} */,
  {32'h404e7d77, 32'hbf9ec1e6} /* (13, 5, 22) {real, imag} */,
  {32'h411ad1ed, 32'h4004d640} /* (13, 5, 21) {real, imag} */,
  {32'h4050fe77, 32'hc0930240} /* (13, 5, 20) {real, imag} */,
  {32'hbfe694ea, 32'hc146230e} /* (13, 5, 19) {real, imag} */,
  {32'h3cbed600, 32'hbfb1984b} /* (13, 5, 18) {real, imag} */,
  {32'h3fe5f66e, 32'h4108851a} /* (13, 5, 17) {real, imag} */,
  {32'h4121b152, 32'h3fba5d4a} /* (13, 5, 16) {real, imag} */,
  {32'h401a1ded, 32'hc031c258} /* (13, 5, 15) {real, imag} */,
  {32'hc0922215, 32'hbf675d00} /* (13, 5, 14) {real, imag} */,
  {32'hbfca0398, 32'h407561f5} /* (13, 5, 13) {real, imag} */,
  {32'h40e6cb05, 32'h4067c836} /* (13, 5, 12) {real, imag} */,
  {32'h41028124, 32'hbf4056ec} /* (13, 5, 11) {real, imag} */,
  {32'h40bc6e45, 32'hc0ab43aa} /* (13, 5, 10) {real, imag} */,
  {32'hbf122048, 32'hc0c6d2ac} /* (13, 5, 9) {real, imag} */,
  {32'hc06af1d2, 32'hc000cc2e} /* (13, 5, 8) {real, imag} */,
  {32'hc04a01b0, 32'hbf4c80cc} /* (13, 5, 7) {real, imag} */,
  {32'hc075404c, 32'hc05b1a46} /* (13, 5, 6) {real, imag} */,
  {32'hc08b0848, 32'hc078858a} /* (13, 5, 5) {real, imag} */,
  {32'hc0bf5e9b, 32'hc02de83a} /* (13, 5, 4) {real, imag} */,
  {32'hc12c2e8f, 32'hbeb75786} /* (13, 5, 3) {real, imag} */,
  {32'h40142189, 32'h40a1046c} /* (13, 5, 2) {real, imag} */,
  {32'h40d26819, 32'h40e7c435} /* (13, 5, 1) {real, imag} */,
  {32'hbf8d839f, 32'hbfcf59de} /* (13, 5, 0) {real, imag} */,
  {32'h405dbf14, 32'h3ffd1dca} /* (13, 4, 31) {real, imag} */,
  {32'h404652c0, 32'h40872bae} /* (13, 4, 30) {real, imag} */,
  {32'h40e03450, 32'hbfd618f9} /* (13, 4, 29) {real, imag} */,
  {32'h408eec4f, 32'hc084eb37} /* (13, 4, 28) {real, imag} */,
  {32'h3b53c400, 32'hc109af76} /* (13, 4, 27) {real, imag} */,
  {32'hc10153f6, 32'hc100db28} /* (13, 4, 26) {real, imag} */,
  {32'hc017f5d4, 32'hc0f84b2c} /* (13, 4, 25) {real, imag} */,
  {32'h408cbc0c, 32'hc0bd5866} /* (13, 4, 24) {real, imag} */,
  {32'h409ea6f2, 32'h3f963fac} /* (13, 4, 23) {real, imag} */,
  {32'h4132eac6, 32'h40ef1414} /* (13, 4, 22) {real, imag} */,
  {32'h40e2e41c, 32'h3fa378e4} /* (13, 4, 21) {real, imag} */,
  {32'h40609bd7, 32'hbfa03376} /* (13, 4, 20) {real, imag} */,
  {32'hc03c13f2, 32'hc038ae23} /* (13, 4, 19) {real, imag} */,
  {32'h3f80a3ce, 32'hc0888f5c} /* (13, 4, 18) {real, imag} */,
  {32'hbdfb38b0, 32'h3db896a0} /* (13, 4, 17) {real, imag} */,
  {32'hc01d5a41, 32'h401c3213} /* (13, 4, 16) {real, imag} */,
  {32'hbe52b070, 32'h40986a89} /* (13, 4, 15) {real, imag} */,
  {32'h3f0167f8, 32'hc00f1137} /* (13, 4, 14) {real, imag} */,
  {32'hbf1bd0b8, 32'hc0b6c055} /* (13, 4, 13) {real, imag} */,
  {32'hbfe1bdd0, 32'hc0f4cf81} /* (13, 4, 12) {real, imag} */,
  {32'hc10052c3, 32'hc0d79374} /* (13, 4, 11) {real, imag} */,
  {32'hc0d2d28b, 32'hbfcba991} /* (13, 4, 10) {real, imag} */,
  {32'hbff4b712, 32'hbea8a3fc} /* (13, 4, 9) {real, imag} */,
  {32'hc0346cc0, 32'hc005faed} /* (13, 4, 8) {real, imag} */,
  {32'h3fd1302d, 32'hbf9c35b6} /* (13, 4, 7) {real, imag} */,
  {32'h406c767c, 32'h3f88f4f5} /* (13, 4, 6) {real, imag} */,
  {32'h400bdf4c, 32'hc085defc} /* (13, 4, 5) {real, imag} */,
  {32'h3fc4c4c7, 32'hc0aaf06e} /* (13, 4, 4) {real, imag} */,
  {32'hc01156b0, 32'hbd582e80} /* (13, 4, 3) {real, imag} */,
  {32'hbfb1cb33, 32'h400bfba4} /* (13, 4, 2) {real, imag} */,
  {32'hbfb70b8e, 32'hbe283e8c} /* (13, 4, 1) {real, imag} */,
  {32'h404ad8c0, 32'hc023338a} /* (13, 4, 0) {real, imag} */,
  {32'h401f9b21, 32'hbfcb1675} /* (13, 3, 31) {real, imag} */,
  {32'hc0374076, 32'hc0878e6d} /* (13, 3, 30) {real, imag} */,
  {32'hc02dbfaa, 32'hc039efb3} /* (13, 3, 29) {real, imag} */,
  {32'h4010af1b, 32'h3f605e1a} /* (13, 3, 28) {real, imag} */,
  {32'hc012fc80, 32'h40e68b60} /* (13, 3, 27) {real, imag} */,
  {32'hc0594626, 32'h3fe65388} /* (13, 3, 26) {real, imag} */,
  {32'hbffb61e8, 32'h402133b4} /* (13, 3, 25) {real, imag} */,
  {32'hbf4320db, 32'h3c767400} /* (13, 3, 24) {real, imag} */,
  {32'h3f8b8d9a, 32'hbfea5028} /* (13, 3, 23) {real, imag} */,
  {32'h40592a60, 32'h3f844648} /* (13, 3, 22) {real, imag} */,
  {32'hc0e401f9, 32'hc0774a40} /* (13, 3, 21) {real, imag} */,
  {32'hc139b15b, 32'h3f42ef9c} /* (13, 3, 20) {real, imag} */,
  {32'h3cb9a2c0, 32'hbf9002a8} /* (13, 3, 19) {real, imag} */,
  {32'h4024b9f0, 32'hbe941a6f} /* (13, 3, 18) {real, imag} */,
  {32'h3f280246, 32'h407ca951} /* (13, 3, 17) {real, imag} */,
  {32'hc00c48dd, 32'h408da86e} /* (13, 3, 16) {real, imag} */,
  {32'h3fb65db6, 32'h3fcb7a93} /* (13, 3, 15) {real, imag} */,
  {32'hbfe15b62, 32'hc042ca6a} /* (13, 3, 14) {real, imag} */,
  {32'hc014793d, 32'hc00b76b8} /* (13, 3, 13) {real, imag} */,
  {32'h3db13540, 32'hbece0308} /* (13, 3, 12) {real, imag} */,
  {32'h3e0cc5d8, 32'h3ee05a78} /* (13, 3, 11) {real, imag} */,
  {32'h3ff46cc9, 32'hc05d316f} /* (13, 3, 10) {real, imag} */,
  {32'h3fd1dda4, 32'h3ef1ccae} /* (13, 3, 9) {real, imag} */,
  {32'h40a3b69d, 32'h4016deed} /* (13, 3, 8) {real, imag} */,
  {32'h40d6ca71, 32'hbfa9b902} /* (13, 3, 7) {real, imag} */,
  {32'h40158c0a, 32'hbf899639} /* (13, 3, 6) {real, imag} */,
  {32'hc001e70a, 32'h40ba2dc9} /* (13, 3, 5) {real, imag} */,
  {32'hc0b271e5, 32'h3fee7949} /* (13, 3, 4) {real, imag} */,
  {32'hc081140f, 32'hc03aa742} /* (13, 3, 3) {real, imag} */,
  {32'hc1142aae, 32'hc0b61564} /* (13, 3, 2) {real, imag} */,
  {32'hc10aad8c, 32'hc0395883} /* (13, 3, 1) {real, imag} */,
  {32'hc0a3835c, 32'h405cdc54} /* (13, 3, 0) {real, imag} */,
  {32'h40b4e396, 32'h40b3f0b5} /* (13, 2, 31) {real, imag} */,
  {32'h413a69e0, 32'h41231a28} /* (13, 2, 30) {real, imag} */,
  {32'hc04fe020, 32'h40b88d6f} /* (13, 2, 29) {real, imag} */,
  {32'hc076fe08, 32'hbfc3aa30} /* (13, 2, 28) {real, imag} */,
  {32'hc0c1d19d, 32'hc09acc92} /* (13, 2, 27) {real, imag} */,
  {32'hc10acb18, 32'hc0aca317} /* (13, 2, 26) {real, imag} */,
  {32'hc0bda7fe, 32'hc09b4d48} /* (13, 2, 25) {real, imag} */,
  {32'hc0cf9401, 32'hc05b3d24} /* (13, 2, 24) {real, imag} */,
  {32'h4096f9dd, 32'hc08eeec0} /* (13, 2, 23) {real, imag} */,
  {32'h40f010b1, 32'hc11210d1} /* (13, 2, 22) {real, imag} */,
  {32'hbf3fecec, 32'hc0503dc6} /* (13, 2, 21) {real, imag} */,
  {32'hbfe8c60c, 32'hbfc3c128} /* (13, 2, 20) {real, imag} */,
  {32'h3fe31c44, 32'hc0c5c05a} /* (13, 2, 19) {real, imag} */,
  {32'h3f94e8f4, 32'h40c16f09} /* (13, 2, 18) {real, imag} */,
  {32'hc0d16700, 32'h40cf2d7b} /* (13, 2, 17) {real, imag} */,
  {32'hbf801905, 32'h4122f89a} /* (13, 2, 16) {real, imag} */,
  {32'h411a5e4a, 32'h412b6075} /* (13, 2, 15) {real, imag} */,
  {32'h41168cbb, 32'h4137fb03} /* (13, 2, 14) {real, imag} */,
  {32'hc0000e4f, 32'h40abcea2} /* (13, 2, 13) {real, imag} */,
  {32'hc059ac6b, 32'hbf7b1b88} /* (13, 2, 12) {real, imag} */,
  {32'h40d58512, 32'hc059f374} /* (13, 2, 11) {real, imag} */,
  {32'h40f06eed, 32'hbfa9c55d} /* (13, 2, 10) {real, imag} */,
  {32'h4134af3e, 32'h40ba1847} /* (13, 2, 9) {real, imag} */,
  {32'h4122f18b, 32'h4092b353} /* (13, 2, 8) {real, imag} */,
  {32'h40ade14f, 32'h40d59ec8} /* (13, 2, 7) {real, imag} */,
  {32'h3f3b1a9c, 32'hc0ba818c} /* (13, 2, 6) {real, imag} */,
  {32'hc006031c, 32'hc1389d5b} /* (13, 2, 5) {real, imag} */,
  {32'h3fb2d234, 32'hc0634036} /* (13, 2, 4) {real, imag} */,
  {32'h409b6894, 32'h4068fa95} /* (13, 2, 3) {real, imag} */,
  {32'h412e270e, 32'hbf83ff26} /* (13, 2, 2) {real, imag} */,
  {32'h40d4fb83, 32'hc096875a} /* (13, 2, 1) {real, imag} */,
  {32'h3edc2f37, 32'hbf2a1f9e} /* (13, 2, 0) {real, imag} */,
  {32'hc01be229, 32'h413175cc} /* (13, 1, 31) {real, imag} */,
  {32'h404c6ecc, 32'h4107e90e} /* (13, 1, 30) {real, imag} */,
  {32'h40a841a0, 32'h400019c4} /* (13, 1, 29) {real, imag} */,
  {32'hbf22d7f0, 32'h409197d2} /* (13, 1, 28) {real, imag} */,
  {32'hc0cd3e78, 32'h41496d94} /* (13, 1, 27) {real, imag} */,
  {32'h3e5e32f8, 32'h3ff6e870} /* (13, 1, 26) {real, imag} */,
  {32'hbee74316, 32'hbfc14b0e} /* (13, 1, 25) {real, imag} */,
  {32'hc0a58f8f, 32'h40357e64} /* (13, 1, 24) {real, imag} */,
  {32'h4088af49, 32'h3f9fe4a6} /* (13, 1, 23) {real, imag} */,
  {32'h410e24e6, 32'hc01dc003} /* (13, 1, 22) {real, imag} */,
  {32'h407bba69, 32'h3f092a46} /* (13, 1, 21) {real, imag} */,
  {32'h4071fffc, 32'h4003ae3c} /* (13, 1, 20) {real, imag} */,
  {32'hc05657d6, 32'h40d3d89a} /* (13, 1, 19) {real, imag} */,
  {32'hc0ca3583, 32'h40414d6c} /* (13, 1, 18) {real, imag} */,
  {32'hc0a6ab6a, 32'h40a3f3b9} /* (13, 1, 17) {real, imag} */,
  {32'h40290b52, 32'h408738b9} /* (13, 1, 16) {real, imag} */,
  {32'h40ef1e63, 32'h40444953} /* (13, 1, 15) {real, imag} */,
  {32'h4044b583, 32'hc07eacd3} /* (13, 1, 14) {real, imag} */,
  {32'hc00bc7a8, 32'h4015a02e} /* (13, 1, 13) {real, imag} */,
  {32'h41407ae8, 32'h3e018200} /* (13, 1, 12) {real, imag} */,
  {32'h40607dfe, 32'hc0e4ab08} /* (13, 1, 11) {real, imag} */,
  {32'h406960bc, 32'hc11e8afa} /* (13, 1, 10) {real, imag} */,
  {32'h409b8e8b, 32'hbfc9442a} /* (13, 1, 9) {real, imag} */,
  {32'h3fc6fc2e, 32'hc0a5e512} /* (13, 1, 8) {real, imag} */,
  {32'hc0622614, 32'h3f7a203c} /* (13, 1, 7) {real, imag} */,
  {32'hc02e05cc, 32'hbff54bee} /* (13, 1, 6) {real, imag} */,
  {32'hbea406f0, 32'hc100d95f} /* (13, 1, 5) {real, imag} */,
  {32'h3f1bf438, 32'hc0c69029} /* (13, 1, 4) {real, imag} */,
  {32'hc01c4d04, 32'hc05787ac} /* (13, 1, 3) {real, imag} */,
  {32'h3f40a3b4, 32'hc10de295} /* (13, 1, 2) {real, imag} */,
  {32'h4135dfed, 32'h3fce56e6} /* (13, 1, 1) {real, imag} */,
  {32'h40eabaf4, 32'h40d922be} /* (13, 1, 0) {real, imag} */,
  {32'hc09e4128, 32'hc0cf58e6} /* (13, 0, 31) {real, imag} */,
  {32'hbe887e00, 32'hc0a691dc} /* (13, 0, 30) {real, imag} */,
  {32'hbecaa8d0, 32'hbfe3e361} /* (13, 0, 29) {real, imag} */,
  {32'hc11d4e58, 32'h40c05be1} /* (13, 0, 28) {real, imag} */,
  {32'hc11d9b88, 32'h3fe6dee7} /* (13, 0, 27) {real, imag} */,
  {32'hbff86b1a, 32'hc03fd4b0} /* (13, 0, 26) {real, imag} */,
  {32'hc01da2a1, 32'h40324241} /* (13, 0, 25) {real, imag} */,
  {32'hc0d89aee, 32'hbd6967a8} /* (13, 0, 24) {real, imag} */,
  {32'hc05e5a2e, 32'hc0488ef0} /* (13, 0, 23) {real, imag} */,
  {32'hc0c389c1, 32'hc0f8b2d6} /* (13, 0, 22) {real, imag} */,
  {32'h400662a6, 32'hc118bc0e} /* (13, 0, 21) {real, imag} */,
  {32'h3f9f7c36, 32'h3e5bd85c} /* (13, 0, 20) {real, imag} */,
  {32'h3e90fc98, 32'hc0035de2} /* (13, 0, 19) {real, imag} */,
  {32'h4105d498, 32'hc03b9b78} /* (13, 0, 18) {real, imag} */,
  {32'h413a31f2, 32'h403bc680} /* (13, 0, 17) {real, imag} */,
  {32'hc0bd980c, 32'h40fc5d55} /* (13, 0, 16) {real, imag} */,
  {32'hc06501cb, 32'h408a2b61} /* (13, 0, 15) {real, imag} */,
  {32'h3fff5a7a, 32'h410dc0ac} /* (13, 0, 14) {real, imag} */,
  {32'hc0934bd4, 32'h40ce076f} /* (13, 0, 13) {real, imag} */,
  {32'hc09acd00, 32'h3f8769d6} /* (13, 0, 12) {real, imag} */,
  {32'h40b391da, 32'hc0520db9} /* (13, 0, 11) {real, imag} */,
  {32'h4007840a, 32'h400be104} /* (13, 0, 10) {real, imag} */,
  {32'h40bf0561, 32'h405928a8} /* (13, 0, 9) {real, imag} */,
  {32'h40f01f80, 32'h409a1d42} /* (13, 0, 8) {real, imag} */,
  {32'h40133564, 32'hc026b122} /* (13, 0, 7) {real, imag} */,
  {32'hc092b6a2, 32'h3f9b03c6} /* (13, 0, 6) {real, imag} */,
  {32'hc0b604be, 32'h3f06dc98} /* (13, 0, 5) {real, imag} */,
  {32'hbeb95cdc, 32'h3f984e6e} /* (13, 0, 4) {real, imag} */,
  {32'h40f15d34, 32'h405c8cb0} /* (13, 0, 3) {real, imag} */,
  {32'h4104df0f, 32'hbe12b62c} /* (13, 0, 2) {real, imag} */,
  {32'h40c66c98, 32'hc0e2bd79} /* (13, 0, 1) {real, imag} */,
  {32'hc0066aee, 32'hc0a67c9d} /* (13, 0, 0) {real, imag} */,
  {32'hc092ab85, 32'hc110da72} /* (12, 31, 31) {real, imag} */,
  {32'hc0c5e65c, 32'hc0d5df88} /* (12, 31, 30) {real, imag} */,
  {32'h408e7621, 32'h3ff5a22e} /* (12, 31, 29) {real, imag} */,
  {32'h3f557d82, 32'h3f571132} /* (12, 31, 28) {real, imag} */,
  {32'hc022e214, 32'h4084c028} /* (12, 31, 27) {real, imag} */,
  {32'hbfbafd42, 32'hbfbd2646} /* (12, 31, 26) {real, imag} */,
  {32'h408144b2, 32'hc0c68d80} /* (12, 31, 25) {real, imag} */,
  {32'hbf0d66b7, 32'hc11856e5} /* (12, 31, 24) {real, imag} */,
  {32'h40061155, 32'h40debfdb} /* (12, 31, 23) {real, imag} */,
  {32'h3fe31712, 32'h410751e6} /* (12, 31, 22) {real, imag} */,
  {32'h4029270d, 32'h4000289f} /* (12, 31, 21) {real, imag} */,
  {32'h4112104f, 32'h403ea1bd} /* (12, 31, 20) {real, imag} */,
  {32'h40d92cf6, 32'hc0a8ac6b} /* (12, 31, 19) {real, imag} */,
  {32'h3f4fb210, 32'hbf6067a0} /* (12, 31, 18) {real, imag} */,
  {32'hc047c0ad, 32'h410d67c0} /* (12, 31, 17) {real, imag} */,
  {32'hc01a959a, 32'hc0b6c33c} /* (12, 31, 16) {real, imag} */,
  {32'h4034cc08, 32'hbf64712e} /* (12, 31, 15) {real, imag} */,
  {32'h415ded20, 32'h40af3096} /* (12, 31, 14) {real, imag} */,
  {32'h4023a26a, 32'h40c8b0b1} /* (12, 31, 13) {real, imag} */,
  {32'h400e859a, 32'h3fc9a684} /* (12, 31, 12) {real, imag} */,
  {32'h40422216, 32'hbf075bb8} /* (12, 31, 11) {real, imag} */,
  {32'h40839647, 32'hc0d23b8a} /* (12, 31, 10) {real, imag} */,
  {32'h40a2b63c, 32'hc057abf6} /* (12, 31, 9) {real, imag} */,
  {32'h41088e7e, 32'h409110da} /* (12, 31, 8) {real, imag} */,
  {32'h40c7d515, 32'hbf977d25} /* (12, 31, 7) {real, imag} */,
  {32'h4047ded6, 32'hbfbd83ae} /* (12, 31, 6) {real, imag} */,
  {32'h40875ac6, 32'h4128a09b} /* (12, 31, 5) {real, imag} */,
  {32'hc092a774, 32'h4120b21c} /* (12, 31, 4) {real, imag} */,
  {32'hc05dce3a, 32'h402237fe} /* (12, 31, 3) {real, imag} */,
  {32'hc090b6d5, 32'h409f2a6f} /* (12, 31, 2) {real, imag} */,
  {32'hc1025684, 32'h40d96cbb} /* (12, 31, 1) {real, imag} */,
  {32'hc02695cc, 32'h40d885e9} /* (12, 31, 0) {real, imag} */,
  {32'h3fc26014, 32'hbf8fe83f} /* (12, 30, 31) {real, imag} */,
  {32'hc0e937cc, 32'hc03e1b01} /* (12, 30, 30) {real, imag} */,
  {32'hc0ee1df1, 32'h4017b7b4} /* (12, 30, 29) {real, imag} */,
  {32'h4004b112, 32'h4085055a} /* (12, 30, 28) {real, imag} */,
  {32'h40a23c3a, 32'hbd8d5a00} /* (12, 30, 27) {real, imag} */,
  {32'h407b1144, 32'hc08bde15} /* (12, 30, 26) {real, imag} */,
  {32'h40e98f4f, 32'hc118942d} /* (12, 30, 25) {real, imag} */,
  {32'h415a8d8f, 32'hbfb4a596} /* (12, 30, 24) {real, imag} */,
  {32'h410e8f90, 32'hc01e3606} /* (12, 30, 23) {real, imag} */,
  {32'h410771af, 32'hc0ceef54} /* (12, 30, 22) {real, imag} */,
  {32'h40e00e8c, 32'hbfc421b8} /* (12, 30, 21) {real, imag} */,
  {32'h4029afd8, 32'hc0aab78e} /* (12, 30, 20) {real, imag} */,
  {32'h40e7a966, 32'hc09769b0} /* (12, 30, 19) {real, imag} */,
  {32'hc0428e60, 32'hc093f0e4} /* (12, 30, 18) {real, imag} */,
  {32'hc107b8bd, 32'hc0e121e0} /* (12, 30, 17) {real, imag} */,
  {32'hc1055aa0, 32'hc0aea38e} /* (12, 30, 16) {real, imag} */,
  {32'hc0f2bed0, 32'hc0155c8a} /* (12, 30, 15) {real, imag} */,
  {32'h3fb79b60, 32'hc02942b4} /* (12, 30, 14) {real, imag} */,
  {32'hbda68630, 32'hc05de97f} /* (12, 30, 13) {real, imag} */,
  {32'hc0a6a894, 32'hc085d5ba} /* (12, 30, 12) {real, imag} */,
  {32'h4020f627, 32'hbf646e28} /* (12, 30, 11) {real, imag} */,
  {32'h402f9cf2, 32'h4002105b} /* (12, 30, 10) {real, imag} */,
  {32'hbdc8a088, 32'hc084ec52} /* (12, 30, 9) {real, imag} */,
  {32'hc0ca4bf9, 32'hc0f0d64a} /* (12, 30, 8) {real, imag} */,
  {32'hc11ae407, 32'h3f15c0c6} /* (12, 30, 7) {real, imag} */,
  {32'hc0a0815c, 32'h4001182a} /* (12, 30, 6) {real, imag} */,
  {32'h40002aa5, 32'h40deef63} /* (12, 30, 5) {real, imag} */,
  {32'hc062ff83, 32'h40aa7178} /* (12, 30, 4) {real, imag} */,
  {32'hc095317e, 32'h412cd5bd} /* (12, 30, 3) {real, imag} */,
  {32'hc07dc643, 32'h401d5ecd} /* (12, 30, 2) {real, imag} */,
  {32'h4101cb6e, 32'h3fd5599b} /* (12, 30, 1) {real, imag} */,
  {32'h41233f2c, 32'h400b39cb} /* (12, 30, 0) {real, imag} */,
  {32'h405e14cb, 32'h3f6e7679} /* (12, 29, 31) {real, imag} */,
  {32'h3fd8dc29, 32'h40988b5c} /* (12, 29, 30) {real, imag} */,
  {32'hbf979e32, 32'h405c1579} /* (12, 29, 29) {real, imag} */,
  {32'hbff4dd1f, 32'h410019bf} /* (12, 29, 28) {real, imag} */,
  {32'hc122af00, 32'h3fed0752} /* (12, 29, 27) {real, imag} */,
  {32'hc12aeb8c, 32'h4053974a} /* (12, 29, 26) {real, imag} */,
  {32'hc12d3cd4, 32'h40aca3dc} /* (12, 29, 25) {real, imag} */,
  {32'hbe02d234, 32'h3ea70004} /* (12, 29, 24) {real, imag} */,
  {32'hbff7597e, 32'hc09ed6ea} /* (12, 29, 23) {real, imag} */,
  {32'hc0c505c4, 32'hc0fbed9a} /* (12, 29, 22) {real, imag} */,
  {32'hc05973b7, 32'hc1513d0a} /* (12, 29, 21) {real, imag} */,
  {32'hc10f125e, 32'hbfbfed28} /* (12, 29, 20) {real, imag} */,
  {32'hc15fc024, 32'h3f6e94a0} /* (12, 29, 19) {real, imag} */,
  {32'hc0989c39, 32'hc0043c99} /* (12, 29, 18) {real, imag} */,
  {32'hc0268ecd, 32'h40152f71} /* (12, 29, 17) {real, imag} */,
  {32'h40868975, 32'h40e59e26} /* (12, 29, 16) {real, imag} */,
  {32'h40c620fc, 32'h40962620} /* (12, 29, 15) {real, imag} */,
  {32'h4133219e, 32'hc0f26a2e} /* (12, 29, 14) {real, imag} */,
  {32'h4103baa2, 32'hc0945e16} /* (12, 29, 13) {real, imag} */,
  {32'h3fbbee14, 32'hc05241c4} /* (12, 29, 12) {real, imag} */,
  {32'h406e6819, 32'hc08ec933} /* (12, 29, 11) {real, imag} */,
  {32'h4055fb78, 32'hc0aa063c} /* (12, 29, 10) {real, imag} */,
  {32'h40070226, 32'hc03e9b6d} /* (12, 29, 9) {real, imag} */,
  {32'h4098ae3d, 32'hbf6852ac} /* (12, 29, 8) {real, imag} */,
  {32'h40c0bd53, 32'h411691e2} /* (12, 29, 7) {real, imag} */,
  {32'h4086f981, 32'h413abc54} /* (12, 29, 6) {real, imag} */,
  {32'h40bb13d7, 32'hc0102e82} /* (12, 29, 5) {real, imag} */,
  {32'h3f3cfcd0, 32'hbec7b8b0} /* (12, 29, 4) {real, imag} */,
  {32'h3f600d00, 32'h40971059} /* (12, 29, 3) {real, imag} */,
  {32'h404dcc5d, 32'hbfdaead5} /* (12, 29, 2) {real, imag} */,
  {32'h414104de, 32'hc0e6ddcc} /* (12, 29, 1) {real, imag} */,
  {32'h40a56074, 32'hc0a2fe2a} /* (12, 29, 0) {real, imag} */,
  {32'hbcff6b50, 32'hc00d7dcc} /* (12, 28, 31) {real, imag} */,
  {32'hbee3b628, 32'h3ff09492} /* (12, 28, 30) {real, imag} */,
  {32'hc0a8c3c0, 32'h40f0643b} /* (12, 28, 29) {real, imag} */,
  {32'h41152237, 32'h3fc0207c} /* (12, 28, 28) {real, imag} */,
  {32'h411f02d1, 32'hc02f7e4a} /* (12, 28, 27) {real, imag} */,
  {32'h3f236782, 32'hbec2dea8} /* (12, 28, 26) {real, imag} */,
  {32'hc06dbc2a, 32'hc0f9f9c7} /* (12, 28, 25) {real, imag} */,
  {32'hc0bfdd6d, 32'hc0bff2f7} /* (12, 28, 24) {real, imag} */,
  {32'hbf8431d0, 32'h40c50d76} /* (12, 28, 23) {real, imag} */,
  {32'h40029510, 32'h3fac5fd2} /* (12, 28, 22) {real, imag} */,
  {32'h405b9df2, 32'hc01f480e} /* (12, 28, 21) {real, imag} */,
  {32'hc0bde77d, 32'h40a65ea3} /* (12, 28, 20) {real, imag} */,
  {32'hc00b518e, 32'h3e8a62ac} /* (12, 28, 19) {real, imag} */,
  {32'h4025724a, 32'hc0208ce8} /* (12, 28, 18) {real, imag} */,
  {32'h4087e637, 32'h410adbe2} /* (12, 28, 17) {real, imag} */,
  {32'h3fb54874, 32'h4117a86c} /* (12, 28, 16) {real, imag} */,
  {32'h3f35e1a4, 32'h40bb250f} /* (12, 28, 15) {real, imag} */,
  {32'h405cd07e, 32'hc080b933} /* (12, 28, 14) {real, imag} */,
  {32'hc022d9fb, 32'hbfdef9fc} /* (12, 28, 13) {real, imag} */,
  {32'hc0f3b97a, 32'hc0af81c5} /* (12, 28, 12) {real, imag} */,
  {32'h3ee9cd70, 32'hc07cb508} /* (12, 28, 11) {real, imag} */,
  {32'h40a09120, 32'hbfc85f3b} /* (12, 28, 10) {real, imag} */,
  {32'hbf8d4e5a, 32'hc00581be} /* (12, 28, 9) {real, imag} */,
  {32'h3f4b61d4, 32'h40e75530} /* (12, 28, 8) {real, imag} */,
  {32'h40ea7d52, 32'h40f8ab48} /* (12, 28, 7) {real, imag} */,
  {32'h4041c32f, 32'h4056a7b1} /* (12, 28, 6) {real, imag} */,
  {32'hbfb407cf, 32'h401122ce} /* (12, 28, 5) {real, imag} */,
  {32'hbf800471, 32'h408446ba} /* (12, 28, 4) {real, imag} */,
  {32'h405cb4fd, 32'h40cf667e} /* (12, 28, 3) {real, imag} */,
  {32'h403c7df8, 32'h40d36f56} /* (12, 28, 2) {real, imag} */,
  {32'hc0413357, 32'h40987e5f} /* (12, 28, 1) {real, imag} */,
  {32'hc087032a, 32'h3fee9f35} /* (12, 28, 0) {real, imag} */,
  {32'hbfe5706f, 32'hc000f48d} /* (12, 27, 31) {real, imag} */,
  {32'h409a22c8, 32'hc0005f11} /* (12, 27, 30) {real, imag} */,
  {32'h412f6290, 32'h4054fb72} /* (12, 27, 29) {real, imag} */,
  {32'h40e1c810, 32'h3f8e5d5c} /* (12, 27, 28) {real, imag} */,
  {32'h40821777, 32'hbff00588} /* (12, 27, 27) {real, imag} */,
  {32'h3ffcc4f6, 32'hc0989cb6} /* (12, 27, 26) {real, imag} */,
  {32'h40914435, 32'hc14019ff} /* (12, 27, 25) {real, imag} */,
  {32'h3ff213d2, 32'hc0bf32b5} /* (12, 27, 24) {real, imag} */,
  {32'h403d5714, 32'h40f2fed4} /* (12, 27, 23) {real, imag} */,
  {32'h402d5f32, 32'h408f41b2} /* (12, 27, 22) {real, imag} */,
  {32'hc02ea9e8, 32'hc00bbabc} /* (12, 27, 21) {real, imag} */,
  {32'hc0305a4a, 32'h40ebc679} /* (12, 27, 20) {real, imag} */,
  {32'h40165e65, 32'h40aa360e} /* (12, 27, 19) {real, imag} */,
  {32'h3ef8bb1e, 32'hbeeecf60} /* (12, 27, 18) {real, imag} */,
  {32'h404b4665, 32'hbf534200} /* (12, 27, 17) {real, imag} */,
  {32'hc0ad11ee, 32'h3f58f1d8} /* (12, 27, 16) {real, imag} */,
  {32'hbf9a5228, 32'hbdc16720} /* (12, 27, 15) {real, imag} */,
  {32'h40949769, 32'hc01eec61} /* (12, 27, 14) {real, imag} */,
  {32'hc00d3e18, 32'h3d88d2fc} /* (12, 27, 13) {real, imag} */,
  {32'hc09b86c9, 32'h40697602} /* (12, 27, 12) {real, imag} */,
  {32'hc0077518, 32'hbf766288} /* (12, 27, 11) {real, imag} */,
  {32'hc0861f3a, 32'hc0db84fc} /* (12, 27, 10) {real, imag} */,
  {32'hbf9e65f6, 32'h40881820} /* (12, 27, 9) {real, imag} */,
  {32'h3ef7379a, 32'h41118c3b} /* (12, 27, 8) {real, imag} */,
  {32'hbdf22160, 32'hc0701611} /* (12, 27, 7) {real, imag} */,
  {32'h40a7d716, 32'hc1149441} /* (12, 27, 6) {real, imag} */,
  {32'h40f2fb92, 32'hc07e2e88} /* (12, 27, 5) {real, imag} */,
  {32'h3edc4c78, 32'h3fa9e752} /* (12, 27, 4) {real, imag} */,
  {32'hc020b792, 32'h408fddbe} /* (12, 27, 3) {real, imag} */,
  {32'h3fa50007, 32'h3f239e20} /* (12, 27, 2) {real, imag} */,
  {32'hbf0f5b97, 32'hc072e5bc} /* (12, 27, 1) {real, imag} */,
  {32'hc0c5bdab, 32'hc0b79d7f} /* (12, 27, 0) {real, imag} */,
  {32'hbfa2d4a8, 32'h40397940} /* (12, 26, 31) {real, imag} */,
  {32'hbeaf8474, 32'h40c0fac7} /* (12, 26, 30) {real, imag} */,
  {32'hc0088569, 32'h40e1189f} /* (12, 26, 29) {real, imag} */,
  {32'hc0985c51, 32'h409e0017} /* (12, 26, 28) {real, imag} */,
  {32'hc03e2768, 32'h40136c90} /* (12, 26, 27) {real, imag} */,
  {32'hc0de90b8, 32'h402b89f6} /* (12, 26, 26) {real, imag} */,
  {32'hc0af5076, 32'h4010227b} /* (12, 26, 25) {real, imag} */,
  {32'h3f8f7eca, 32'hc06a6c29} /* (12, 26, 24) {real, imag} */,
  {32'h403e81d0, 32'hc13062bc} /* (12, 26, 23) {real, imag} */,
  {32'h3f964b5c, 32'hc0b004d6} /* (12, 26, 22) {real, imag} */,
  {32'hc035f820, 32'h40b70498} /* (12, 26, 21) {real, imag} */,
  {32'h40681f4c, 32'h4042eb4d} /* (12, 26, 20) {real, imag} */,
  {32'h404898bb, 32'hc010630f} /* (12, 26, 19) {real, imag} */,
  {32'hbfeda2b5, 32'hbfae0684} /* (12, 26, 18) {real, imag} */,
  {32'hc0f254a0, 32'hc0ce80a7} /* (12, 26, 17) {real, imag} */,
  {32'hc0b0f298, 32'hc0a48015} /* (12, 26, 16) {real, imag} */,
  {32'hbf8e62e0, 32'hc0938647} /* (12, 26, 15) {real, imag} */,
  {32'h408bc0d4, 32'hbdd3eb40} /* (12, 26, 14) {real, imag} */,
  {32'h411d7328, 32'h40ed50aa} /* (12, 26, 13) {real, imag} */,
  {32'h402b38fd, 32'h3ffa0689} /* (12, 26, 12) {real, imag} */,
  {32'hbfd819e6, 32'h40993e42} /* (12, 26, 11) {real, imag} */,
  {32'h403810c2, 32'h402149cd} /* (12, 26, 10) {real, imag} */,
  {32'h4106b5e9, 32'h40a308c3} /* (12, 26, 9) {real, imag} */,
  {32'h40d462eb, 32'h405c2e32} /* (12, 26, 8) {real, imag} */,
  {32'h40bdb610, 32'hc0b15359} /* (12, 26, 7) {real, imag} */,
  {32'hbfaa9482, 32'hc146b319} /* (12, 26, 6) {real, imag} */,
  {32'hbce46000, 32'hc02a332c} /* (12, 26, 5) {real, imag} */,
  {32'hc07db888, 32'h3f100fee} /* (12, 26, 4) {real, imag} */,
  {32'hc0e58a32, 32'h3f67f36c} /* (12, 26, 3) {real, imag} */,
  {32'hc0655abc, 32'h3f1411a6} /* (12, 26, 2) {real, imag} */,
  {32'hbffed50e, 32'h3e98b678} /* (12, 26, 1) {real, imag} */,
  {32'h3fb3d0e9, 32'h40277f8a} /* (12, 26, 0) {real, imag} */,
  {32'hbff2851a, 32'h3ffb9fc0} /* (12, 25, 31) {real, imag} */,
  {32'hc0d6ac4a, 32'h402b9853} /* (12, 25, 30) {real, imag} */,
  {32'hc07ef352, 32'hc003c6d0} /* (12, 25, 29) {real, imag} */,
  {32'hc003bde4, 32'h3f9d952c} /* (12, 25, 28) {real, imag} */,
  {32'h40543082, 32'h411346b8} /* (12, 25, 27) {real, imag} */,
  {32'hc032f98d, 32'h40dd23e6} /* (12, 25, 26) {real, imag} */,
  {32'hc092269d, 32'h3f760194} /* (12, 25, 25) {real, imag} */,
  {32'hc0e2b17e, 32'hbf9d9826} /* (12, 25, 24) {real, imag} */,
  {32'hc02f38be, 32'hc0902c78} /* (12, 25, 23) {real, imag} */,
  {32'hc07f4e52, 32'hc000834c} /* (12, 25, 22) {real, imag} */,
  {32'hc0267546, 32'h4033ff90} /* (12, 25, 21) {real, imag} */,
  {32'hc0b4c662, 32'h3c56d580} /* (12, 25, 20) {real, imag} */,
  {32'hc0ca525c, 32'hc080ddd6} /* (12, 25, 19) {real, imag} */,
  {32'hc0ddb5b8, 32'hbf57fb84} /* (12, 25, 18) {real, imag} */,
  {32'hc0b92f64, 32'h40dc1743} /* (12, 25, 17) {real, imag} */,
  {32'h400ab648, 32'h40dd2750} /* (12, 25, 16) {real, imag} */,
  {32'h40ceadf5, 32'h40288ffe} /* (12, 25, 15) {real, imag} */,
  {32'h40b71e68, 32'h40ada03a} /* (12, 25, 14) {real, imag} */,
  {32'hc050a295, 32'h3f3cc5e7} /* (12, 25, 13) {real, imag} */,
  {32'hc01b5aab, 32'hc0a61694} /* (12, 25, 12) {real, imag} */,
  {32'h3fcb0178, 32'h3facd126} /* (12, 25, 11) {real, imag} */,
  {32'h3fbe77f2, 32'h409adf23} /* (12, 25, 10) {real, imag} */,
  {32'hbe14ff50, 32'h3fba543c} /* (12, 25, 9) {real, imag} */,
  {32'hc0e2a41c, 32'hbf256dec} /* (12, 25, 8) {real, imag} */,
  {32'hbf7e9467, 32'h3ddde440} /* (12, 25, 7) {real, imag} */,
  {32'h3fa3ff0c, 32'h40794e92} /* (12, 25, 6) {real, imag} */,
  {32'h4095ef50, 32'h3e9b90b2} /* (12, 25, 5) {real, imag} */,
  {32'h40c66d46, 32'hc0bda0ff} /* (12, 25, 4) {real, imag} */,
  {32'h40a9bdb6, 32'hc0d30a36} /* (12, 25, 3) {real, imag} */,
  {32'h406d4df5, 32'h3d0330e0} /* (12, 25, 2) {real, imag} */,
  {32'h3fd43b93, 32'h4055719c} /* (12, 25, 1) {real, imag} */,
  {32'h3e14abc8, 32'hc011fe9e} /* (12, 25, 0) {real, imag} */,
  {32'hc0749eb5, 32'h3ed5c5b0} /* (12, 24, 31) {real, imag} */,
  {32'h3ffbd316, 32'hbfbcca4c} /* (12, 24, 30) {real, imag} */,
  {32'h400dd209, 32'h4075210f} /* (12, 24, 29) {real, imag} */,
  {32'hbf94eb34, 32'h3e356a14} /* (12, 24, 28) {real, imag} */,
  {32'h408ae178, 32'hbee47893} /* (12, 24, 27) {real, imag} */,
  {32'h40507a69, 32'hbf86969c} /* (12, 24, 26) {real, imag} */,
  {32'h40e66f70, 32'hc06878b5} /* (12, 24, 25) {real, imag} */,
  {32'h411ca77a, 32'hbe849000} /* (12, 24, 24) {real, imag} */,
  {32'h406a73a8, 32'hbf74fcc2} /* (12, 24, 23) {real, imag} */,
  {32'h40b4f6ec, 32'hbeeee608} /* (12, 24, 22) {real, imag} */,
  {32'hbf320834, 32'h401fe7af} /* (12, 24, 21) {real, imag} */,
  {32'hbfd8efba, 32'h4055202e} /* (12, 24, 20) {real, imag} */,
  {32'hbffacd0a, 32'h40c3f844} /* (12, 24, 19) {real, imag} */,
  {32'h400cfc1c, 32'hc068a373} /* (12, 24, 18) {real, imag} */,
  {32'h407e8904, 32'h3ffa3038} /* (12, 24, 17) {real, imag} */,
  {32'h3fc0b4fb, 32'h411ba5a4} /* (12, 24, 16) {real, imag} */,
  {32'h400425e1, 32'hbedb8968} /* (12, 24, 15) {real, imag} */,
  {32'hbf727aca, 32'hc0e13b48} /* (12, 24, 14) {real, imag} */,
  {32'h3f90b950, 32'hc07ae336} /* (12, 24, 13) {real, imag} */,
  {32'h40e8663a, 32'hc02d1c22} /* (12, 24, 12) {real, imag} */,
  {32'h4122fba9, 32'h3fb51a82} /* (12, 24, 11) {real, imag} */,
  {32'h3ecc9236, 32'h40f3f7a2} /* (12, 24, 10) {real, imag} */,
  {32'hc0bcc299, 32'h3f907cd6} /* (12, 24, 9) {real, imag} */,
  {32'hbe3c3780, 32'h3db76f10} /* (12, 24, 8) {real, imag} */,
  {32'h3fd7f3f3, 32'hbe8f3a36} /* (12, 24, 7) {real, imag} */,
  {32'h4063ea16, 32'hc10e3058} /* (12, 24, 6) {real, imag} */,
  {32'h408086eb, 32'hc0c1953b} /* (12, 24, 5) {real, imag} */,
  {32'h4003bff4, 32'hbfc30056} /* (12, 24, 4) {real, imag} */,
  {32'h4008a32d, 32'hc02c690e} /* (12, 24, 3) {real, imag} */,
  {32'h404e9171, 32'hbfdeb802} /* (12, 24, 2) {real, imag} */,
  {32'h3fb951dd, 32'h408c1196} /* (12, 24, 1) {real, imag} */,
  {32'hbfa08ef6, 32'h40ed3cd3} /* (12, 24, 0) {real, imag} */,
  {32'hbd5298c0, 32'h40173a1a} /* (12, 23, 31) {real, imag} */,
  {32'h3f8608f4, 32'hbe80e500} /* (12, 23, 30) {real, imag} */,
  {32'hbfaba476, 32'hc052e5ec} /* (12, 23, 29) {real, imag} */,
  {32'hc031aa3a, 32'hc05447b8} /* (12, 23, 28) {real, imag} */,
  {32'h3dc7cbb8, 32'hc00147f0} /* (12, 23, 27) {real, imag} */,
  {32'hc024412e, 32'h40076608} /* (12, 23, 26) {real, imag} */,
  {32'h3d2ca960, 32'h4018b0c5} /* (12, 23, 25) {real, imag} */,
  {32'h3ff73392, 32'h3e0047d0} /* (12, 23, 24) {real, imag} */,
  {32'h405ed828, 32'h40390cc5} /* (12, 23, 23) {real, imag} */,
  {32'h40330da8, 32'h40a34136} /* (12, 23, 22) {real, imag} */,
  {32'h3ef77578, 32'h3fe924ee} /* (12, 23, 21) {real, imag} */,
  {32'h40175018, 32'h40daf999} /* (12, 23, 20) {real, imag} */,
  {32'h4084c400, 32'h4013fd2c} /* (12, 23, 19) {real, imag} */,
  {32'h403aa62b, 32'h408d7a06} /* (12, 23, 18) {real, imag} */,
  {32'hc02b5315, 32'h40b7e7cd} /* (12, 23, 17) {real, imag} */,
  {32'hc07ad18c, 32'h3fb73123} /* (12, 23, 16) {real, imag} */,
  {32'hbfe463e6, 32'h3fcdfbcd} /* (12, 23, 15) {real, imag} */,
  {32'h3fcb7e35, 32'hc088d8ba} /* (12, 23, 14) {real, imag} */,
  {32'h3ff113ce, 32'hc00c0da0} /* (12, 23, 13) {real, imag} */,
  {32'h3fccac10, 32'h400dbd5e} /* (12, 23, 12) {real, imag} */,
  {32'hbf06fe58, 32'h4011e142} /* (12, 23, 11) {real, imag} */,
  {32'hc0a450e1, 32'h40d29e58} /* (12, 23, 10) {real, imag} */,
  {32'hc100b7c0, 32'hbf8184a8} /* (12, 23, 9) {real, imag} */,
  {32'hc0f2ec4f, 32'hbe17fdf8} /* (12, 23, 8) {real, imag} */,
  {32'hc0ab19c0, 32'hbfa458b2} /* (12, 23, 7) {real, imag} */,
  {32'h3f8e1d20, 32'h3e70d58c} /* (12, 23, 6) {real, imag} */,
  {32'h3f80ed6c, 32'h40ae870c} /* (12, 23, 5) {real, imag} */,
  {32'hc07a7a2a, 32'hbd0c29a0} /* (12, 23, 4) {real, imag} */,
  {32'hc0603bfe, 32'hc0bd00e2} /* (12, 23, 3) {real, imag} */,
  {32'hc097d191, 32'hbfd163d1} /* (12, 23, 2) {real, imag} */,
  {32'hc099147c, 32'h3fdb6a38} /* (12, 23, 1) {real, imag} */,
  {32'hbf108d84, 32'h3ea97143} /* (12, 23, 0) {real, imag} */,
  {32'h3dca06e0, 32'h3e2a0848} /* (12, 22, 31) {real, imag} */,
  {32'hbf816f4c, 32'hbfc43dbe} /* (12, 22, 30) {real, imag} */,
  {32'hbe62fda4, 32'h3ed51a9c} /* (12, 22, 29) {real, imag} */,
  {32'h3f90196b, 32'h40304064} /* (12, 22, 28) {real, imag} */,
  {32'hbfa7b635, 32'h3d840370} /* (12, 22, 27) {real, imag} */,
  {32'h3d4ef300, 32'h404ef21b} /* (12, 22, 26) {real, imag} */,
  {32'hbf37efee, 32'hbe6d2cd0} /* (12, 22, 25) {real, imag} */,
  {32'h3ff1d3c2, 32'h3e62aa70} /* (12, 22, 24) {real, imag} */,
  {32'h3fba7fb7, 32'h409b7b96} /* (12, 22, 23) {real, imag} */,
  {32'hbf9b7c27, 32'h408dc7f6} /* (12, 22, 22) {real, imag} */,
  {32'hc093b660, 32'hc03dfcca} /* (12, 22, 21) {real, imag} */,
  {32'h3e90e744, 32'hc090541f} /* (12, 22, 20) {real, imag} */,
  {32'h4040b6b8, 32'hc0757982} /* (12, 22, 19) {real, imag} */,
  {32'h409fba87, 32'hc002a0f6} /* (12, 22, 18) {real, imag} */,
  {32'h40dc7522, 32'hc0858fb4} /* (12, 22, 17) {real, imag} */,
  {32'h4072959d, 32'h3ecc7322} /* (12, 22, 16) {real, imag} */,
  {32'h3fbf3a20, 32'h3fe986ce} /* (12, 22, 15) {real, imag} */,
  {32'h4013339a, 32'h409267fc} /* (12, 22, 14) {real, imag} */,
  {32'h3eeebe68, 32'h4086df12} /* (12, 22, 13) {real, imag} */,
  {32'h3ea6889a, 32'h40a0e59b} /* (12, 22, 12) {real, imag} */,
  {32'h3f665978, 32'hbeef5e68} /* (12, 22, 11) {real, imag} */,
  {32'hc02ad314, 32'hbfe750dc} /* (12, 22, 10) {real, imag} */,
  {32'hc0e35d1c, 32'hbfe9f0ec} /* (12, 22, 9) {real, imag} */,
  {32'hc0d6692a, 32'hbf8951da} /* (12, 22, 8) {real, imag} */,
  {32'hc000a80c, 32'h3dd3def0} /* (12, 22, 7) {real, imag} */,
  {32'h3f8d8a36, 32'h3fc6d18a} /* (12, 22, 6) {real, imag} */,
  {32'hbfba28ac, 32'h40682725} /* (12, 22, 5) {real, imag} */,
  {32'hc02e4d0c, 32'h40c3b1fc} /* (12, 22, 4) {real, imag} */,
  {32'hc0884b80, 32'h412f9852} /* (12, 22, 3) {real, imag} */,
  {32'hbfb38b59, 32'h40f751e8} /* (12, 22, 2) {real, imag} */,
  {32'h4013c256, 32'hbf8dc3be} /* (12, 22, 1) {real, imag} */,
  {32'h4010d7e8, 32'h3e820ef4} /* (12, 22, 0) {real, imag} */,
  {32'h3f7a8b3e, 32'hbffc6a62} /* (12, 21, 31) {real, imag} */,
  {32'h3efb66bc, 32'hc03b9f64} /* (12, 21, 30) {real, imag} */,
  {32'h4015923f, 32'h3ebe26a0} /* (12, 21, 29) {real, imag} */,
  {32'hbe23886c, 32'h409814f1} /* (12, 21, 28) {real, imag} */,
  {32'hbc666bc0, 32'hbd63fc80} /* (12, 21, 27) {real, imag} */,
  {32'hbdb967a8, 32'h3ea739fa} /* (12, 21, 26) {real, imag} */,
  {32'h3f5e3a1e, 32'h3f7a618c} /* (12, 21, 25) {real, imag} */,
  {32'hbe8b71e6, 32'hc00f27d4} /* (12, 21, 24) {real, imag} */,
  {32'hc08dfb36, 32'hbe9a4068} /* (12, 21, 23) {real, imag} */,
  {32'hc0232236, 32'hbea78158} /* (12, 21, 22) {real, imag} */,
  {32'h3e83a3a4, 32'hbc3a1e80} /* (12, 21, 21) {real, imag} */,
  {32'hbe8e52e8, 32'h409ee8c0} /* (12, 21, 20) {real, imag} */,
  {32'h401339d0, 32'h3e99e504} /* (12, 21, 19) {real, imag} */,
  {32'h409331d0, 32'hc0ea0584} /* (12, 21, 18) {real, imag} */,
  {32'h3e8f78c6, 32'hc0e9e6ec} /* (12, 21, 17) {real, imag} */,
  {32'hbd8dd870, 32'hc023f424} /* (12, 21, 16) {real, imag} */,
  {32'h402675d8, 32'h3fd3079c} /* (12, 21, 15) {real, imag} */,
  {32'hbe6952a8, 32'hbe8ea994} /* (12, 21, 14) {real, imag} */,
  {32'hc090adb3, 32'hc00e9949} /* (12, 21, 13) {real, imag} */,
  {32'hc0589d68, 32'hbfb3b388} /* (12, 21, 12) {real, imag} */,
  {32'hc04544b8, 32'h3fc1c8dd} /* (12, 21, 11) {real, imag} */,
  {32'hc000a043, 32'hbd6b2980} /* (12, 21, 10) {real, imag} */,
  {32'h4013e354, 32'h3ea85aec} /* (12, 21, 9) {real, imag} */,
  {32'h402eda64, 32'hbfa4becd} /* (12, 21, 8) {real, imag} */,
  {32'h3fabaf5a, 32'h3f0ccb6c} /* (12, 21, 7) {real, imag} */,
  {32'hbfd9136a, 32'h4078b5a0} /* (12, 21, 6) {real, imag} */,
  {32'hc0016813, 32'hbf404ff4} /* (12, 21, 5) {real, imag} */,
  {32'h3fd5a932, 32'hbe97b2a6} /* (12, 21, 4) {real, imag} */,
  {32'hbe3353e0, 32'h408bca35} /* (12, 21, 3) {real, imag} */,
  {32'h4008a2fa, 32'h3f6c02f4} /* (12, 21, 2) {real, imag} */,
  {32'h406d555d, 32'h3ca70500} /* (12, 21, 1) {real, imag} */,
  {32'h4000b1d8, 32'hbf228936} /* (12, 21, 0) {real, imag} */,
  {32'h401a6744, 32'hbf8c75b9} /* (12, 20, 31) {real, imag} */,
  {32'h40d5c5da, 32'h3e855500} /* (12, 20, 30) {real, imag} */,
  {32'h409a539e, 32'hc041fcc0} /* (12, 20, 29) {real, imag} */,
  {32'hbeb1eb3c, 32'hc0727e98} /* (12, 20, 28) {real, imag} */,
  {32'h40005975, 32'h3ddb3b70} /* (12, 20, 27) {real, imag} */,
  {32'h3fed4b72, 32'hbd94f740} /* (12, 20, 26) {real, imag} */,
  {32'hc0619db8, 32'h4073abbf} /* (12, 20, 25) {real, imag} */,
  {32'hc025c854, 32'h40dd748d} /* (12, 20, 24) {real, imag} */,
  {32'hbdb25e40, 32'h3f60476c} /* (12, 20, 23) {real, imag} */,
  {32'h4021c12f, 32'hc03a71db} /* (12, 20, 22) {real, imag} */,
  {32'h3f8d6836, 32'h3fbd4fb7} /* (12, 20, 21) {real, imag} */,
  {32'hc0229f7a, 32'hc01193a0} /* (12, 20, 20) {real, imag} */,
  {32'hc0919c46, 32'hbdd885d0} /* (12, 20, 19) {real, imag} */,
  {32'hc00107dd, 32'h409e1e21} /* (12, 20, 18) {real, imag} */,
  {32'hbf0963f3, 32'h400dda60} /* (12, 20, 17) {real, imag} */,
  {32'hc024f4a0, 32'hbf411a7c} /* (12, 20, 16) {real, imag} */,
  {32'hc0118916, 32'hbf9c037c} /* (12, 20, 15) {real, imag} */,
  {32'hbee9af4c, 32'hbf350f42} /* (12, 20, 14) {real, imag} */,
  {32'h3fe1a2ca, 32'hbfa10ab8} /* (12, 20, 13) {real, imag} */,
  {32'hbfb48bc4, 32'hbf3de14a} /* (12, 20, 12) {real, imag} */,
  {32'h3e17e990, 32'h3fb0e755} /* (12, 20, 11) {real, imag} */,
  {32'h404b236c, 32'h4089babe} /* (12, 20, 10) {real, imag} */,
  {32'h3fbc8dfe, 32'h40294da8} /* (12, 20, 9) {real, imag} */,
  {32'h3fa5d83a, 32'h3e9dcf28} /* (12, 20, 8) {real, imag} */,
  {32'hbe7d2e56, 32'hbf4ba406} /* (12, 20, 7) {real, imag} */,
  {32'hc055131b, 32'h4001cd0b} /* (12, 20, 6) {real, imag} */,
  {32'hbeb0547c, 32'h406af824} /* (12, 20, 5) {real, imag} */,
  {32'hbfb09adb, 32'hbe656b6e} /* (12, 20, 4) {real, imag} */,
  {32'hbfd7e566, 32'hbfcfed3b} /* (12, 20, 3) {real, imag} */,
  {32'hbf9ea304, 32'hbfa39c66} /* (12, 20, 2) {real, imag} */,
  {32'hbe41c380, 32'hc0384ea1} /* (12, 20, 1) {real, imag} */,
  {32'h3ef7d1ea, 32'hbf46f71a} /* (12, 20, 0) {real, imag} */,
  {32'h3f86944e, 32'h3fa7437c} /* (12, 19, 31) {real, imag} */,
  {32'h3f2ac490, 32'h3fcaf625} /* (12, 19, 30) {real, imag} */,
  {32'hbf39adfc, 32'hbdc54b58} /* (12, 19, 29) {real, imag} */,
  {32'hbf3bff1e, 32'hbff33c4c} /* (12, 19, 28) {real, imag} */,
  {32'h40039de8, 32'hc04e351c} /* (12, 19, 27) {real, imag} */,
  {32'h3fecfc5e, 32'hc072c5c8} /* (12, 19, 26) {real, imag} */,
  {32'h3da8d980, 32'h3fb69cd1} /* (12, 19, 25) {real, imag} */,
  {32'hbfca3910, 32'hbe3e5478} /* (12, 19, 24) {real, imag} */,
  {32'h3b8a5a80, 32'hc03a6970} /* (12, 19, 23) {real, imag} */,
  {32'h3f7e2ece, 32'hc0a078f3} /* (12, 19, 22) {real, imag} */,
  {32'h3e682d60, 32'hc06b1f79} /* (12, 19, 21) {real, imag} */,
  {32'hbd72df80, 32'hbec481f0} /* (12, 19, 20) {real, imag} */,
  {32'h3fe2dba8, 32'h3ff8db80} /* (12, 19, 19) {real, imag} */,
  {32'h3d60ddf0, 32'h3fa336b2} /* (12, 19, 18) {real, imag} */,
  {32'hc017f439, 32'hbf18df04} /* (12, 19, 17) {real, imag} */,
  {32'h3fd2a4a2, 32'hbe5f1958} /* (12, 19, 16) {real, imag} */,
  {32'h3fb3cf09, 32'h3fdcb773} /* (12, 19, 15) {real, imag} */,
  {32'hc006fae8, 32'h3eb51d68} /* (12, 19, 14) {real, imag} */,
  {32'hbf154630, 32'hc028e665} /* (12, 19, 13) {real, imag} */,
  {32'hc02c8a76, 32'hbffb77b8} /* (12, 19, 12) {real, imag} */,
  {32'hc05210f2, 32'hc09308af} /* (12, 19, 11) {real, imag} */,
  {32'h3cce8400, 32'hc0cb8dac} /* (12, 19, 10) {real, imag} */,
  {32'h3f9ad473, 32'hbff1a7a2} /* (12, 19, 9) {real, imag} */,
  {32'hbe68aa60, 32'h40137c6b} /* (12, 19, 8) {real, imag} */,
  {32'hbf89febc, 32'h3e004760} /* (12, 19, 7) {real, imag} */,
  {32'hc00e744c, 32'hbee5b918} /* (12, 19, 6) {real, imag} */,
  {32'hc06a663b, 32'h3df8f130} /* (12, 19, 5) {real, imag} */,
  {32'hc0481920, 32'h3e96c440} /* (12, 19, 4) {real, imag} */,
  {32'h40420eac, 32'h3fcd2cce} /* (12, 19, 3) {real, imag} */,
  {32'h40875a98, 32'h3ef8dbd4} /* (12, 19, 2) {real, imag} */,
  {32'h3fb1099c, 32'hbff6fe16} /* (12, 19, 1) {real, imag} */,
  {32'h3fc0d843, 32'hbf116776} /* (12, 19, 0) {real, imag} */,
  {32'h3fb4227c, 32'h3f67e160} /* (12, 18, 31) {real, imag} */,
  {32'hbeb57c1a, 32'h3ff85125} /* (12, 18, 30) {real, imag} */,
  {32'h3ff88360, 32'h406bc46f} /* (12, 18, 29) {real, imag} */,
  {32'h401de46c, 32'h3eb171c0} /* (12, 18, 28) {real, imag} */,
  {32'h3f9d9450, 32'h3e2848d0} /* (12, 18, 27) {real, imag} */,
  {32'hbecfc30c, 32'h3f16c3a8} /* (12, 18, 26) {real, imag} */,
  {32'h3f931c8f, 32'hbfdd68aa} /* (12, 18, 25) {real, imag} */,
  {32'hbe961568, 32'hc0465fb6} /* (12, 18, 24) {real, imag} */,
  {32'hbe2a8338, 32'hbfeca35d} /* (12, 18, 23) {real, imag} */,
  {32'h3ff9b907, 32'hbf6dd0d4} /* (12, 18, 22) {real, imag} */,
  {32'hbef0e860, 32'hbf834b1d} /* (12, 18, 21) {real, imag} */,
  {32'hc051f373, 32'h40463369} /* (12, 18, 20) {real, imag} */,
  {32'hbfa250b9, 32'h40581c20} /* (12, 18, 19) {real, imag} */,
  {32'h3fa99432, 32'h3fa244a8} /* (12, 18, 18) {real, imag} */,
  {32'hbf907437, 32'h3f991d2a} /* (12, 18, 17) {real, imag} */,
  {32'hc05c7b48, 32'hc00b69c8} /* (12, 18, 16) {real, imag} */,
  {32'hbe94a430, 32'h3eb5b722} /* (12, 18, 15) {real, imag} */,
  {32'hbfcd05fb, 32'h400d80c3} /* (12, 18, 14) {real, imag} */,
  {32'hbf164056, 32'h3fcc12b2} /* (12, 18, 13) {real, imag} */,
  {32'h40271cdc, 32'hbec52260} /* (12, 18, 12) {real, imag} */,
  {32'h3f1c0534, 32'hbf33923c} /* (12, 18, 11) {real, imag} */,
  {32'h3faacf38, 32'h3f31557b} /* (12, 18, 10) {real, imag} */,
  {32'h4022bd17, 32'hc0067e0c} /* (12, 18, 9) {real, imag} */,
  {32'h3ffc04ac, 32'h403b41e6} /* (12, 18, 8) {real, imag} */,
  {32'h40114814, 32'h3ffacee2} /* (12, 18, 7) {real, imag} */,
  {32'h3ded1b74, 32'h3ee8e058} /* (12, 18, 6) {real, imag} */,
  {32'hbf2ae5e8, 32'h3f593cda} /* (12, 18, 5) {real, imag} */,
  {32'hbf9635de, 32'h3f2bdd82} /* (12, 18, 4) {real, imag} */,
  {32'hbf3b7ca3, 32'h3f655ca2} /* (12, 18, 3) {real, imag} */,
  {32'hbe5b1e00, 32'h3e064f1c} /* (12, 18, 2) {real, imag} */,
  {32'h400ea814, 32'h3fd6322f} /* (12, 18, 1) {real, imag} */,
  {32'h3fa3b64c, 32'h3ecf4893} /* (12, 18, 0) {real, imag} */,
  {32'hbe8d19e0, 32'hbffceb39} /* (12, 17, 31) {real, imag} */,
  {32'hbfa2562c, 32'hbffc302b} /* (12, 17, 30) {real, imag} */,
  {32'hbfcc6379, 32'hbf0ea1b0} /* (12, 17, 29) {real, imag} */,
  {32'hbf05c462, 32'hbfada425} /* (12, 17, 28) {real, imag} */,
  {32'h3f3304e9, 32'hc01b5e92} /* (12, 17, 27) {real, imag} */,
  {32'hbec24128, 32'h3e0b0590} /* (12, 17, 26) {real, imag} */,
  {32'hc003c841, 32'h3fa9bb5f} /* (12, 17, 25) {real, imag} */,
  {32'hbff6dd7a, 32'h3f3654d4} /* (12, 17, 24) {real, imag} */,
  {32'hbf402092, 32'h3f0a2c40} /* (12, 17, 23) {real, imag} */,
  {32'hbf92b206, 32'h3f3f8a98} /* (12, 17, 22) {real, imag} */,
  {32'hbfae0777, 32'hbfc6f99b} /* (12, 17, 21) {real, imag} */,
  {32'hbfe36ed8, 32'hc02f2d44} /* (12, 17, 20) {real, imag} */,
  {32'hc01b0b1d, 32'hbee06b62} /* (12, 17, 19) {real, imag} */,
  {32'hbd8c3390, 32'hbe37f548} /* (12, 17, 18) {real, imag} */,
  {32'h408d3450, 32'h3dabfd40} /* (12, 17, 17) {real, imag} */,
  {32'h4045b255, 32'h40025589} /* (12, 17, 16) {real, imag} */,
  {32'hbff7147a, 32'h3fab97de} /* (12, 17, 15) {real, imag} */,
  {32'hbf876436, 32'h3f11e206} /* (12, 17, 14) {real, imag} */,
  {32'h3fe7aec9, 32'h3edc7f7a} /* (12, 17, 13) {real, imag} */,
  {32'h3fa6afd2, 32'h3febe16f} /* (12, 17, 12) {real, imag} */,
  {32'h3fa34d1e, 32'h3f2ea87d} /* (12, 17, 11) {real, imag} */,
  {32'h3fc19022, 32'hbf525e76} /* (12, 17, 10) {real, imag} */,
  {32'h3f5ecd1b, 32'hc0380b02} /* (12, 17, 9) {real, imag} */,
  {32'hc0008ffe, 32'hc0358726} /* (12, 17, 8) {real, imag} */,
  {32'hbfc24a88, 32'h3f70782f} /* (12, 17, 7) {real, imag} */,
  {32'h3f241c98, 32'h3fdfedfb} /* (12, 17, 6) {real, imag} */,
  {32'h3f5b88d5, 32'h3d61eb40} /* (12, 17, 5) {real, imag} */,
  {32'hbf93e460, 32'hc0a099fc} /* (12, 17, 4) {real, imag} */,
  {32'hbf5694e6, 32'hc06140fe} /* (12, 17, 3) {real, imag} */,
  {32'h3fd482df, 32'hbf4b3086} /* (12, 17, 2) {real, imag} */,
  {32'h3fcecab8, 32'hbe9bbd29} /* (12, 17, 1) {real, imag} */,
  {32'h3fc36ee4, 32'hbe2ec212} /* (12, 17, 0) {real, imag} */,
  {32'hbeba3b98, 32'h3f8032c6} /* (12, 16, 31) {real, imag} */,
  {32'hbed6d730, 32'h3f38bda4} /* (12, 16, 30) {real, imag} */,
  {32'h4010a3e2, 32'h3f02fd34} /* (12, 16, 29) {real, imag} */,
  {32'h4000aea1, 32'hbf961ca4} /* (12, 16, 28) {real, imag} */,
  {32'hbd100178, 32'hbf9d97b2} /* (12, 16, 27) {real, imag} */,
  {32'hbe5ffdf0, 32'h3f219e00} /* (12, 16, 26) {real, imag} */,
  {32'h3ec78a40, 32'h3fdef038} /* (12, 16, 25) {real, imag} */,
  {32'h3f4c65a4, 32'hbfbaebd2} /* (12, 16, 24) {real, imag} */,
  {32'h3e8db798, 32'hc02626c8} /* (12, 16, 23) {real, imag} */,
  {32'hbf1703a8, 32'hc0058bd4} /* (12, 16, 22) {real, imag} */,
  {32'h3f611362, 32'hbf577e58} /* (12, 16, 21) {real, imag} */,
  {32'h3c45da00, 32'h3e804d20} /* (12, 16, 20) {real, imag} */,
  {32'h3eeb74f0, 32'h3fa5d2e4} /* (12, 16, 19) {real, imag} */,
  {32'h3f9d7d5c, 32'h40125a14} /* (12, 16, 18) {real, imag} */,
  {32'hbf219774, 32'h3f924115} /* (12, 16, 17) {real, imag} */,
  {32'hbf8a2376, 32'hbfb7f11a} /* (12, 16, 16) {real, imag} */,
  {32'h3f7ab6cb, 32'h3f9820aa} /* (12, 16, 15) {real, imag} */,
  {32'h4034d6d4, 32'h3fc12fd4} /* (12, 16, 14) {real, imag} */,
  {32'h3f299528, 32'h400664aa} /* (12, 16, 13) {real, imag} */,
  {32'hc007f900, 32'h3f046360} /* (12, 16, 12) {real, imag} */,
  {32'hbfc3eef8, 32'h3e4f27c0} /* (12, 16, 11) {real, imag} */,
  {32'hc045e05c, 32'h3f7dcaf0} /* (12, 16, 10) {real, imag} */,
  {32'hbfebdaf0, 32'hbf58acd6} /* (12, 16, 9) {real, imag} */,
  {32'hbfd2abae, 32'hbd57c5a0} /* (12, 16, 8) {real, imag} */,
  {32'hbf4e0916, 32'hbf6e5106} /* (12, 16, 7) {real, imag} */,
  {32'h40075134, 32'hc00ddc05} /* (12, 16, 6) {real, imag} */,
  {32'h3f831d0e, 32'hbfe50bb4} /* (12, 16, 5) {real, imag} */,
  {32'h3f6bc010, 32'hbfe734d4} /* (12, 16, 4) {real, imag} */,
  {32'h4004f2ec, 32'hbfd697d6} /* (12, 16, 3) {real, imag} */,
  {32'h3fb28338, 32'h3fd05d54} /* (12, 16, 2) {real, imag} */,
  {32'h3f0ea8dc, 32'hbed7f904} /* (12, 16, 1) {real, imag} */,
  {32'hbf8babd8, 32'h3f7b9e0c} /* (12, 16, 0) {real, imag} */,
  {32'hbf5ac7f8, 32'h3fafc919} /* (12, 15, 31) {real, imag} */,
  {32'h3e6e1fa0, 32'h3fdca98b} /* (12, 15, 30) {real, imag} */,
  {32'h3faa22e1, 32'h3ebea280} /* (12, 15, 29) {real, imag} */,
  {32'h4070e164, 32'h4009b324} /* (12, 15, 28) {real, imag} */,
  {32'h3eda5852, 32'h3f9f0d13} /* (12, 15, 27) {real, imag} */,
  {32'hbfc55797, 32'hc0046d8b} /* (12, 15, 26) {real, imag} */,
  {32'h3fbb7976, 32'hbf99b5bf} /* (12, 15, 25) {real, imag} */,
  {32'h3f850b0e, 32'hbef13d08} /* (12, 15, 24) {real, imag} */,
  {32'hbcb26130, 32'hbdc996c0} /* (12, 15, 23) {real, imag} */,
  {32'h3fc3a806, 32'hbee86160} /* (12, 15, 22) {real, imag} */,
  {32'h3eb79174, 32'hbe44c8a0} /* (12, 15, 21) {real, imag} */,
  {32'h3f3c58e0, 32'h3f5da951} /* (12, 15, 20) {real, imag} */,
  {32'hbf2b649c, 32'h3f83c554} /* (12, 15, 19) {real, imag} */,
  {32'h3ff7ed0f, 32'h3fa26779} /* (12, 15, 18) {real, imag} */,
  {32'h40635c4a, 32'hbde920c0} /* (12, 15, 17) {real, imag} */,
  {32'hbeeccc58, 32'hc011abc5} /* (12, 15, 16) {real, imag} */,
  {32'hbfd94ba4, 32'h3dfafcf8} /* (12, 15, 15) {real, imag} */,
  {32'hbfe314ce, 32'h3febf5e9} /* (12, 15, 14) {real, imag} */,
  {32'hbeedef14, 32'h3f1bd42b} /* (12, 15, 13) {real, imag} */,
  {32'h3f8a575a, 32'h3e14d2b0} /* (12, 15, 12) {real, imag} */,
  {32'h3fbb90a6, 32'hbf688835} /* (12, 15, 11) {real, imag} */,
  {32'hbf3467a4, 32'hbfba21c5} /* (12, 15, 10) {real, imag} */,
  {32'hbe2966e4, 32'hbe0066f8} /* (12, 15, 9) {real, imag} */,
  {32'hbe8613d0, 32'hbf980759} /* (12, 15, 8) {real, imag} */,
  {32'h3d922df8, 32'hbedfecee} /* (12, 15, 7) {real, imag} */,
  {32'hbf82d0b4, 32'h4045183a} /* (12, 15, 6) {real, imag} */,
  {32'hbe004144, 32'hbf8d5b76} /* (12, 15, 5) {real, imag} */,
  {32'h3f677b00, 32'hbf617564} /* (12, 15, 4) {real, imag} */,
  {32'h3f913815, 32'hbec86df4} /* (12, 15, 3) {real, imag} */,
  {32'h3fbf2f5d, 32'hbfc0cb3d} /* (12, 15, 2) {real, imag} */,
  {32'h4026d968, 32'hbf5ed6e4} /* (12, 15, 1) {real, imag} */,
  {32'h3f8244bc, 32'h3e883429} /* (12, 15, 0) {real, imag} */,
  {32'hc0290316, 32'h3f73b138} /* (12, 14, 31) {real, imag} */,
  {32'h3f183f63, 32'h3f851ad7} /* (12, 14, 30) {real, imag} */,
  {32'h3f35f6a0, 32'h401aff7f} /* (12, 14, 29) {real, imag} */,
  {32'hbf2a5e6a, 32'hbd723780} /* (12, 14, 28) {real, imag} */,
  {32'hbf9b1810, 32'hc06c552c} /* (12, 14, 27) {real, imag} */,
  {32'hbf55d91a, 32'hc05f8c44} /* (12, 14, 26) {real, imag} */,
  {32'hbfc60a87, 32'hc069e91b} /* (12, 14, 25) {real, imag} */,
  {32'h3ff098da, 32'hbe2695e8} /* (12, 14, 24) {real, imag} */,
  {32'h3f96c77b, 32'h401b2742} /* (12, 14, 23) {real, imag} */,
  {32'hbe468ce8, 32'h406da567} /* (12, 14, 22) {real, imag} */,
  {32'h3fc14828, 32'h3fbad7b1} /* (12, 14, 21) {real, imag} */,
  {32'h3fbd9c0a, 32'hbf41a7cc} /* (12, 14, 20) {real, imag} */,
  {32'hbdb285d0, 32'hbff4b0c8} /* (12, 14, 19) {real, imag} */,
  {32'hbf83c080, 32'h3ddcd040} /* (12, 14, 18) {real, imag} */,
  {32'h3fca50cf, 32'h404e4561} /* (12, 14, 17) {real, imag} */,
  {32'h3f191c80, 32'h40169330} /* (12, 14, 16) {real, imag} */,
  {32'h3f5e3dd8, 32'h3f6e7cbd} /* (12, 14, 15) {real, imag} */,
  {32'hbd3f27c0, 32'h3e8e717e} /* (12, 14, 14) {real, imag} */,
  {32'hbf130c22, 32'h3ecd8058} /* (12, 14, 13) {real, imag} */,
  {32'h3f0c26d6, 32'hbfc44810} /* (12, 14, 12) {real, imag} */,
  {32'hbfcc8c1e, 32'hbf0fd36c} /* (12, 14, 11) {real, imag} */,
  {32'hc0839b02, 32'h3e259e4c} /* (12, 14, 10) {real, imag} */,
  {32'hbf1f2c5b, 32'h3f348df0} /* (12, 14, 9) {real, imag} */,
  {32'h3fd6a958, 32'h3ffa824c} /* (12, 14, 8) {real, imag} */,
  {32'h3fd6a349, 32'h402f630f} /* (12, 14, 7) {real, imag} */,
  {32'hbe0ece1a, 32'hbdb3a820} /* (12, 14, 6) {real, imag} */,
  {32'h3f34e2b0, 32'h3fd8dc43} /* (12, 14, 5) {real, imag} */,
  {32'hc0429cd7, 32'h3fe4ff27} /* (12, 14, 4) {real, imag} */,
  {32'h3f28f653, 32'h3fce1133} /* (12, 14, 3) {real, imag} */,
  {32'h407c01d6, 32'hbfc37d20} /* (12, 14, 2) {real, imag} */,
  {32'hbf9c6c28, 32'hbf81651b} /* (12, 14, 1) {real, imag} */,
  {32'hc021177e, 32'hbf86f131} /* (12, 14, 0) {real, imag} */,
  {32'hc076af4f, 32'hc00b361a} /* (12, 13, 31) {real, imag} */,
  {32'hc0bb396e, 32'hbff0c821} /* (12, 13, 30) {real, imag} */,
  {32'hbf34f89c, 32'hbf090f83} /* (12, 13, 29) {real, imag} */,
  {32'h3ff35ea9, 32'h3fd4b4f4} /* (12, 13, 28) {real, imag} */,
  {32'h4011668c, 32'h403fd5cc} /* (12, 13, 27) {real, imag} */,
  {32'h3ffc1c36, 32'h3fdc75af} /* (12, 13, 26) {real, imag} */,
  {32'h400d0536, 32'hbfa2e14f} /* (12, 13, 25) {real, imag} */,
  {32'h40015380, 32'hc03c5f14} /* (12, 13, 24) {real, imag} */,
  {32'h3ff395fa, 32'hbfbc4767} /* (12, 13, 23) {real, imag} */,
  {32'hbe799e58, 32'h3d9e1f80} /* (12, 13, 22) {real, imag} */,
  {32'h3fb943e0, 32'h3fe9d1a2} /* (12, 13, 21) {real, imag} */,
  {32'h402ea799, 32'h3f798718} /* (12, 13, 20) {real, imag} */,
  {32'h401fbb1c, 32'hc01753fa} /* (12, 13, 19) {real, imag} */,
  {32'h3fc125c8, 32'hc0763d67} /* (12, 13, 18) {real, imag} */,
  {32'h405347cf, 32'hc05fd123} /* (12, 13, 17) {real, imag} */,
  {32'h3f260f4c, 32'hbfa768a5} /* (12, 13, 16) {real, imag} */,
  {32'h3ffbc6d7, 32'h3f85b767} /* (12, 13, 15) {real, imag} */,
  {32'h408b8eac, 32'h40221685} /* (12, 13, 14) {real, imag} */,
  {32'h400366be, 32'h3fed97ae} /* (12, 13, 13) {real, imag} */,
  {32'h3fedf57c, 32'h400667f8} /* (12, 13, 12) {real, imag} */,
  {32'h3eb22150, 32'h3f90c394} /* (12, 13, 11) {real, imag} */,
  {32'hc02eaf02, 32'hbf17a964} /* (12, 13, 10) {real, imag} */,
  {32'hc015322c, 32'hbf6fd014} /* (12, 13, 9) {real, imag} */,
  {32'hbf7f18e0, 32'h3c2bb900} /* (12, 13, 8) {real, imag} */,
  {32'hbfb7c818, 32'hbe4c85a0} /* (12, 13, 7) {real, imag} */,
  {32'hbe6094b8, 32'h3e8625e8} /* (12, 13, 6) {real, imag} */,
  {32'hbfa3ba96, 32'h3f07379a} /* (12, 13, 5) {real, imag} */,
  {32'h3ee71210, 32'hbfaa3b68} /* (12, 13, 4) {real, imag} */,
  {32'h404eb4e2, 32'h3ecd80a8} /* (12, 13, 3) {real, imag} */,
  {32'hbd91a320, 32'h40236fce} /* (12, 13, 2) {real, imag} */,
  {32'h402876ea, 32'h4041c33f} /* (12, 13, 1) {real, imag} */,
  {32'h3ee383b4, 32'h3fd71353} /* (12, 13, 0) {real, imag} */,
  {32'h3fe2a290, 32'h3f8c8c0d} /* (12, 12, 31) {real, imag} */,
  {32'hbf325e7c, 32'h401e609c} /* (12, 12, 30) {real, imag} */,
  {32'hbff9b1b2, 32'h4023404c} /* (12, 12, 29) {real, imag} */,
  {32'h3f61411e, 32'h3eced98c} /* (12, 12, 28) {real, imag} */,
  {32'hbff9be42, 32'hbf758df6} /* (12, 12, 27) {real, imag} */,
  {32'hbf826c30, 32'h402c3fea} /* (12, 12, 26) {real, imag} */,
  {32'hbfcdf028, 32'h3f8d6d06} /* (12, 12, 25) {real, imag} */,
  {32'hbf7a1a11, 32'h4010ff0a} /* (12, 12, 24) {real, imag} */,
  {32'hbfd187b6, 32'h40658f61} /* (12, 12, 23) {real, imag} */,
  {32'h40597f4d, 32'h4074ebb7} /* (12, 12, 22) {real, imag} */,
  {32'h404f6f79, 32'h3f1f4212} /* (12, 12, 21) {real, imag} */,
  {32'h3f8213dd, 32'h3f586c94} /* (12, 12, 20) {real, imag} */,
  {32'h402cc7a1, 32'h403f70b6} /* (12, 12, 19) {real, imag} */,
  {32'h402320b5, 32'h3dfc7fc0} /* (12, 12, 18) {real, imag} */,
  {32'hbe61590c, 32'hc091cf50} /* (12, 12, 17) {real, imag} */,
  {32'hc0050fa4, 32'hbe74ae90} /* (12, 12, 16) {real, imag} */,
  {32'hbf09e54e, 32'h3fabdd6c} /* (12, 12, 15) {real, imag} */,
  {32'h3f18875a, 32'hbedec85c} /* (12, 12, 14) {real, imag} */,
  {32'h3fa3642a, 32'h3fad9c26} /* (12, 12, 13) {real, imag} */,
  {32'h40cd1a03, 32'h403ff9f6} /* (12, 12, 12) {real, imag} */,
  {32'h4093f55e, 32'h3fc64a17} /* (12, 12, 11) {real, imag} */,
  {32'h3fee8dc5, 32'h401f2bec} /* (12, 12, 10) {real, imag} */,
  {32'h3fe95962, 32'h40a839fc} /* (12, 12, 9) {real, imag} */,
  {32'h3fe690e2, 32'h40a41432} /* (12, 12, 8) {real, imag} */,
  {32'h3f9796dd, 32'h3f900301} /* (12, 12, 7) {real, imag} */,
  {32'h3fb86cc6, 32'hc006e509} /* (12, 12, 6) {real, imag} */,
  {32'hbfd19c73, 32'hbf5bf9ae} /* (12, 12, 5) {real, imag} */,
  {32'h3f842a89, 32'h3e667cd2} /* (12, 12, 4) {real, imag} */,
  {32'h400d82b2, 32'h403ac074} /* (12, 12, 3) {real, imag} */,
  {32'h3f9332ca, 32'h40b0b0ea} /* (12, 12, 2) {real, imag} */,
  {32'h3ff77d34, 32'h40299707} /* (12, 12, 1) {real, imag} */,
  {32'h3f331f19, 32'hbf9f0b45} /* (12, 12, 0) {real, imag} */,
  {32'h4007f9f4, 32'hbf59e38d} /* (12, 11, 31) {real, imag} */,
  {32'h3f1c68da, 32'hc097f131} /* (12, 11, 30) {real, imag} */,
  {32'h3f59a2dc, 32'hc0a63ece} /* (12, 11, 29) {real, imag} */,
  {32'h400403eb, 32'hc0d2ac35} /* (12, 11, 28) {real, imag} */,
  {32'h3fefb024, 32'hc081c487} /* (12, 11, 27) {real, imag} */,
  {32'hbfd01952, 32'h3f61bbc3} /* (12, 11, 26) {real, imag} */,
  {32'hbfb39ab9, 32'h402de27f} /* (12, 11, 25) {real, imag} */,
  {32'h3e270e94, 32'hc05942ec} /* (12, 11, 24) {real, imag} */,
  {32'h3e5febd0, 32'hc08dd92e} /* (12, 11, 23) {real, imag} */,
  {32'hbf96c83f, 32'h4058a625} /* (12, 11, 22) {real, imag} */,
  {32'h3df34af0, 32'h401efe66} /* (12, 11, 21) {real, imag} */,
  {32'h402489dd, 32'hbc610c00} /* (12, 11, 20) {real, imag} */,
  {32'h3fac8b90, 32'h402705d4} /* (12, 11, 19) {real, imag} */,
  {32'h3f24458c, 32'h4089ac9e} /* (12, 11, 18) {real, imag} */,
  {32'hc00d13ed, 32'hbf95c150} /* (12, 11, 17) {real, imag} */,
  {32'hc04dbac8, 32'hbfeb8b1d} /* (12, 11, 16) {real, imag} */,
  {32'hc09f6bfc, 32'hbf8940a4} /* (12, 11, 15) {real, imag} */,
  {32'h3f206d76, 32'hbec86fdc} /* (12, 11, 14) {real, imag} */,
  {32'h3f98fb65, 32'hbfdbcd2e} /* (12, 11, 13) {real, imag} */,
  {32'hbf1b0b4e, 32'hbf01cf24} /* (12, 11, 12) {real, imag} */,
  {32'h407fe7dc, 32'hc0576a84} /* (12, 11, 11) {real, imag} */,
  {32'h3eb22198, 32'hc051be76} /* (12, 11, 10) {real, imag} */,
  {32'h3ecdd518, 32'hbf9df813} /* (12, 11, 9) {real, imag} */,
  {32'h40137b0c, 32'h3f485142} /* (12, 11, 8) {real, imag} */,
  {32'hbfb2d4d8, 32'hc04859bb} /* (12, 11, 7) {real, imag} */,
  {32'hc0700b97, 32'hc08cb2c6} /* (12, 11, 6) {real, imag} */,
  {32'hc0a99564, 32'h3f4db454} /* (12, 11, 5) {real, imag} */,
  {32'hc03519dd, 32'h3ff6fb0e} /* (12, 11, 4) {real, imag} */,
  {32'h3feee4d4, 32'h3f54bea0} /* (12, 11, 3) {real, imag} */,
  {32'hc02cf0aa, 32'hbfc2afbe} /* (12, 11, 2) {real, imag} */,
  {32'hc024d10b, 32'hc0492eb6} /* (12, 11, 1) {real, imag} */,
  {32'h406a63a6, 32'h3ecef514} /* (12, 11, 0) {real, imag} */,
  {32'hc05dc376, 32'h3f24ba0a} /* (12, 10, 31) {real, imag} */,
  {32'hbf8a94c0, 32'h3d1e2bd0} /* (12, 10, 30) {real, imag} */,
  {32'hbe8c973a, 32'hc038a630} /* (12, 10, 29) {real, imag} */,
  {32'hbfbc96a7, 32'hc01c7c84} /* (12, 10, 28) {real, imag} */,
  {32'hc022c970, 32'hc01d6eee} /* (12, 10, 27) {real, imag} */,
  {32'hc0354f62, 32'h407da799} /* (12, 10, 26) {real, imag} */,
  {32'hbf60b05a, 32'hbf37a19c} /* (12, 10, 25) {real, imag} */,
  {32'hbf83e9a6, 32'hbfd89872} /* (12, 10, 24) {real, imag} */,
  {32'h3fc1675b, 32'hc0cc6666} /* (12, 10, 23) {real, imag} */,
  {32'hc091be62, 32'hc08ba102} /* (12, 10, 22) {real, imag} */,
  {32'hc05e7d54, 32'h3eed3bfc} /* (12, 10, 21) {real, imag} */,
  {32'hc01484b0, 32'h3ff6ba21} /* (12, 10, 20) {real, imag} */,
  {32'h3e039be0, 32'h40c09b83} /* (12, 10, 19) {real, imag} */,
  {32'h40086bd0, 32'h403d580a} /* (12, 10, 18) {real, imag} */,
  {32'h400d3eb4, 32'h40710e98} /* (12, 10, 17) {real, imag} */,
  {32'h4022f3b1, 32'hbf2eac33} /* (12, 10, 16) {real, imag} */,
  {32'h40a16420, 32'hbfaa2fb0} /* (12, 10, 15) {real, imag} */,
  {32'h403d4f8c, 32'h3e9f0e70} /* (12, 10, 14) {real, imag} */,
  {32'h401fe4fd, 32'h3fbc45c0} /* (12, 10, 13) {real, imag} */,
  {32'hbfacd0b2, 32'h3e085da0} /* (12, 10, 12) {real, imag} */,
  {32'hc07cdcc2, 32'hc02ca47d} /* (12, 10, 11) {real, imag} */,
  {32'hbe819e54, 32'hbf51ee78} /* (12, 10, 10) {real, imag} */,
  {32'h40347171, 32'hbfd6afa0} /* (12, 10, 9) {real, imag} */,
  {32'h40602af4, 32'hbf7f5734} /* (12, 10, 8) {real, imag} */,
  {32'h4038eea8, 32'h3fdf7d69} /* (12, 10, 7) {real, imag} */,
  {32'hbedc3796, 32'h3fde3f9e} /* (12, 10, 6) {real, imag} */,
  {32'hc040ac2e, 32'h4025d32f} /* (12, 10, 5) {real, imag} */,
  {32'hc0043578, 32'hc05d5ba0} /* (12, 10, 4) {real, imag} */,
  {32'h3fb36f2d, 32'hbd8a3600} /* (12, 10, 3) {real, imag} */,
  {32'h4065a9cc, 32'h3f82b2d0} /* (12, 10, 2) {real, imag} */,
  {32'hc048649e, 32'hc04188e9} /* (12, 10, 1) {real, imag} */,
  {32'hc09e30fa, 32'hbfbd0a9d} /* (12, 10, 0) {real, imag} */,
  {32'hc06962a9, 32'h3efb6d60} /* (12, 9, 31) {real, imag} */,
  {32'hc0f88169, 32'h3ebae168} /* (12, 9, 30) {real, imag} */,
  {32'hc10246c6, 32'h40795230} /* (12, 9, 29) {real, imag} */,
  {32'hc1023800, 32'h3f192392} /* (12, 9, 28) {real, imag} */,
  {32'hbfdf98d2, 32'h3ea5db44} /* (12, 9, 27) {real, imag} */,
  {32'h3f7634f0, 32'hbea48944} /* (12, 9, 26) {real, imag} */,
  {32'hbf0fedba, 32'hc035ad4d} /* (12, 9, 25) {real, imag} */,
  {32'hc047014b, 32'hc08259c4} /* (12, 9, 24) {real, imag} */,
  {32'h3e1d6800, 32'hc0057bc1} /* (12, 9, 23) {real, imag} */,
  {32'h4054c2dc, 32'hbd93ae60} /* (12, 9, 22) {real, imag} */,
  {32'h4053f31b, 32'hbe8e5ada} /* (12, 9, 21) {real, imag} */,
  {32'h409e5b70, 32'hbf312bd8} /* (12, 9, 20) {real, imag} */,
  {32'h3fcfe880, 32'hbedcee30} /* (12, 9, 19) {real, imag} */,
  {32'hbe7bfcf0, 32'h3f1db374} /* (12, 9, 18) {real, imag} */,
  {32'h3fc02022, 32'h3f404308} /* (12, 9, 17) {real, imag} */,
  {32'h401b8268, 32'h407feba8} /* (12, 9, 16) {real, imag} */,
  {32'h403d8929, 32'h4094b7b1} /* (12, 9, 15) {real, imag} */,
  {32'h4030d0fe, 32'h3f452c74} /* (12, 9, 14) {real, imag} */,
  {32'h407d986d, 32'hc09666cf} /* (12, 9, 13) {real, imag} */,
  {32'h40ce3294, 32'hbe233b48} /* (12, 9, 12) {real, imag} */,
  {32'h3e8d76d8, 32'hc08d125a} /* (12, 9, 11) {real, imag} */,
  {32'hc09dc945, 32'hc0ec0dbc} /* (12, 9, 10) {real, imag} */,
  {32'hbf7d4268, 32'hc046fe2c} /* (12, 9, 9) {real, imag} */,
  {32'h4017eabe, 32'hbf7d382a} /* (12, 9, 8) {real, imag} */,
  {32'hbea8bfe0, 32'h4012ee15} /* (12, 9, 7) {real, imag} */,
  {32'h402a12ca, 32'hc006c61c} /* (12, 9, 6) {real, imag} */,
  {32'h408cfc55, 32'hc0e1257e} /* (12, 9, 5) {real, imag} */,
  {32'h3ffb0b4f, 32'hc07d0b3e} /* (12, 9, 4) {real, imag} */,
  {32'hbefcc9a0, 32'hbffc1656} /* (12, 9, 3) {real, imag} */,
  {32'h40bb0483, 32'h3f65d1b6} /* (12, 9, 2) {real, imag} */,
  {32'h3f274854, 32'hbfa8d85e} /* (12, 9, 1) {real, imag} */,
  {32'hc0996324, 32'h3f1bb53a} /* (12, 9, 0) {real, imag} */,
  {32'h3fca20c2, 32'hc0a8ec91} /* (12, 8, 31) {real, imag} */,
  {32'hbed01e12, 32'hc105c3a2} /* (12, 8, 30) {real, imag} */,
  {32'hc04af867, 32'hc119a730} /* (12, 8, 29) {real, imag} */,
  {32'hc09ae6e3, 32'hbf8d8506} /* (12, 8, 28) {real, imag} */,
  {32'h3f34f928, 32'h3ec3c50b} /* (12, 8, 27) {real, imag} */,
  {32'hc00a52fb, 32'hc006d4ad} /* (12, 8, 26) {real, imag} */,
  {32'hc079be90, 32'h3f8c35e6} /* (12, 8, 25) {real, imag} */,
  {32'hbf6c3d50, 32'h406fd0aa} /* (12, 8, 24) {real, imag} */,
  {32'h3fb464cf, 32'h4070ed6e} /* (12, 8, 23) {real, imag} */,
  {32'h3fb85ce8, 32'h401ee279} /* (12, 8, 22) {real, imag} */,
  {32'hc01d0612, 32'h40967452} /* (12, 8, 21) {real, imag} */,
  {32'hc0994ff8, 32'h40a277cd} /* (12, 8, 20) {real, imag} */,
  {32'hbfd25452, 32'hc008f918} /* (12, 8, 19) {real, imag} */,
  {32'h405345a4, 32'hc08ad3e4} /* (12, 8, 18) {real, imag} */,
  {32'h409674a4, 32'hc075d19c} /* (12, 8, 17) {real, imag} */,
  {32'h402a4b72, 32'hc049c3ef} /* (12, 8, 16) {real, imag} */,
  {32'h3f8e3be0, 32'hc0980a98} /* (12, 8, 15) {real, imag} */,
  {32'hbf8f7a75, 32'hc04cda79} /* (12, 8, 14) {real, imag} */,
  {32'hbf0925f0, 32'hbf991103} /* (12, 8, 13) {real, imag} */,
  {32'hbead5720, 32'hbe88d76c} /* (12, 8, 12) {real, imag} */,
  {32'h404464ff, 32'h3e5ef64c} /* (12, 8, 11) {real, imag} */,
  {32'h400991ed, 32'hbf893ec0} /* (12, 8, 10) {real, imag} */,
  {32'h409f0df7, 32'h3e0fd020} /* (12, 8, 9) {real, imag} */,
  {32'h406de8ee, 32'h4001afec} /* (12, 8, 8) {real, imag} */,
  {32'hc0513366, 32'h3fb66106} /* (12, 8, 7) {real, imag} */,
  {32'hbf8b26bf, 32'h4085f52c} /* (12, 8, 6) {real, imag} */,
  {32'h40007f96, 32'h3f94ee28} /* (12, 8, 5) {real, imag} */,
  {32'hbf54a7fa, 32'h4089cef4} /* (12, 8, 4) {real, imag} */,
  {32'hc02fa78f, 32'h4033af98} /* (12, 8, 3) {real, imag} */,
  {32'h3fc3aade, 32'h408725c8} /* (12, 8, 2) {real, imag} */,
  {32'h409d9d7f, 32'h408b292e} /* (12, 8, 1) {real, imag} */,
  {32'h40863e94, 32'h4043d78e} /* (12, 8, 0) {real, imag} */,
  {32'hbfa26ad6, 32'h3fc41f34} /* (12, 7, 31) {real, imag} */,
  {32'hbdae1400, 32'hbeb033d0} /* (12, 7, 30) {real, imag} */,
  {32'h3f87dfaf, 32'h3f927818} /* (12, 7, 29) {real, imag} */,
  {32'h3fd324c3, 32'h40b3f141} /* (12, 7, 28) {real, imag} */,
  {32'hbf7283e8, 32'h3f2f6960} /* (12, 7, 27) {real, imag} */,
  {32'h4091481e, 32'h3f629e40} /* (12, 7, 26) {real, imag} */,
  {32'h412f18c8, 32'h40bbe836} /* (12, 7, 25) {real, imag} */,
  {32'h408b0e6c, 32'h40334a25} /* (12, 7, 24) {real, imag} */,
  {32'hc07479fe, 32'hc0ef5bfe} /* (12, 7, 23) {real, imag} */,
  {32'hbe021460, 32'hc0d87e62} /* (12, 7, 22) {real, imag} */,
  {32'h40529666, 32'hbea639a0} /* (12, 7, 21) {real, imag} */,
  {32'h3fd5f970, 32'hc047dfaa} /* (12, 7, 20) {real, imag} */,
  {32'h3fc266b0, 32'hc047612d} /* (12, 7, 19) {real, imag} */,
  {32'hbe9bd958, 32'hc103b19f} /* (12, 7, 18) {real, imag} */,
  {32'hbfd4d99a, 32'h4019a4ae} /* (12, 7, 17) {real, imag} */,
  {32'hc01aefec, 32'h3e1c23f0} /* (12, 7, 16) {real, imag} */,
  {32'hbfcbbcd4, 32'hc0ce25f3} /* (12, 7, 15) {real, imag} */,
  {32'h403f244c, 32'hbfcf0a3a} /* (12, 7, 14) {real, imag} */,
  {32'h4084ad0e, 32'h3f419081} /* (12, 7, 13) {real, imag} */,
  {32'h403258b1, 32'hc049919d} /* (12, 7, 12) {real, imag} */,
  {32'h3f800eb2, 32'hc0bb0080} /* (12, 7, 11) {real, imag} */,
  {32'h4064275b, 32'hc118dd3c} /* (12, 7, 10) {real, imag} */,
  {32'h406462b8, 32'hc0eb9677} /* (12, 7, 9) {real, imag} */,
  {32'h411c2dd6, 32'hc0e08b10} /* (12, 7, 8) {real, imag} */,
  {32'hbf4ded1b, 32'hc084547f} /* (12, 7, 7) {real, imag} */,
  {32'hc087a42a, 32'hbe438520} /* (12, 7, 6) {real, imag} */,
  {32'hc0ce2c48, 32'h3ed9c552} /* (12, 7, 5) {real, imag} */,
  {32'hc0a3ba26, 32'hc0d68cef} /* (12, 7, 4) {real, imag} */,
  {32'hbe9210d0, 32'hbf0c28f4} /* (12, 7, 3) {real, imag} */,
  {32'h406c9a77, 32'hc02e94ba} /* (12, 7, 2) {real, imag} */,
  {32'h3fdb6b03, 32'hbf398e32} /* (12, 7, 1) {real, imag} */,
  {32'h3f33ab66, 32'hbfdc1ae4} /* (12, 7, 0) {real, imag} */,
  {32'h3fbcdef6, 32'hbf70ce86} /* (12, 6, 31) {real, imag} */,
  {32'h4002ad94, 32'h3f06af08} /* (12, 6, 30) {real, imag} */,
  {32'h3f0f0f49, 32'h40258ae6} /* (12, 6, 29) {real, imag} */,
  {32'hc02600c4, 32'h3f308238} /* (12, 6, 28) {real, imag} */,
  {32'h3ddc47f0, 32'hc0b6fb68} /* (12, 6, 27) {real, imag} */,
  {32'hbfefe1e2, 32'hbf40ffee} /* (12, 6, 26) {real, imag} */,
  {32'hbf95c5e2, 32'h4091b656} /* (12, 6, 25) {real, imag} */,
  {32'hc0e3f0f0, 32'h403a8217} /* (12, 6, 24) {real, imag} */,
  {32'hc0569e36, 32'h40a059d5} /* (12, 6, 23) {real, imag} */,
  {32'h3f8fb32a, 32'h40a9d54a} /* (12, 6, 22) {real, imag} */,
  {32'hc018c12e, 32'hbf4ce0fc} /* (12, 6, 21) {real, imag} */,
  {32'hbe34d668, 32'h3fca007e} /* (12, 6, 20) {real, imag} */,
  {32'hbff51176, 32'h4053dd5f} /* (12, 6, 19) {real, imag} */,
  {32'hbdeb7370, 32'h41487bd0} /* (12, 6, 18) {real, imag} */,
  {32'hbf4ee500, 32'h4154df6a} /* (12, 6, 17) {real, imag} */,
  {32'h40c6fa9a, 32'h4001a23e} /* (12, 6, 16) {real, imag} */,
  {32'h40ec52b6, 32'h3ed48cb0} /* (12, 6, 15) {real, imag} */,
  {32'hc02781db, 32'h40ce5c22} /* (12, 6, 14) {real, imag} */,
  {32'hc0a17ca8, 32'h40c05598} /* (12, 6, 13) {real, imag} */,
  {32'hc09b0f52, 32'h40699be8} /* (12, 6, 12) {real, imag} */,
  {32'h3f7a4b0b, 32'h3efea588} /* (12, 6, 11) {real, imag} */,
  {32'h40121734, 32'hbffbe91e} /* (12, 6, 10) {real, imag} */,
  {32'hc0b0b98d, 32'hbfcfc400} /* (12, 6, 9) {real, imag} */,
  {32'hc1115ce5, 32'hc0c94733} /* (12, 6, 8) {real, imag} */,
  {32'hbf3e3750, 32'hc10897bd} /* (12, 6, 7) {real, imag} */,
  {32'hbe11edb4, 32'hc0ffc716} /* (12, 6, 6) {real, imag} */,
  {32'hbfeb4a90, 32'h3ecf5444} /* (12, 6, 5) {real, imag} */,
  {32'h3f318f32, 32'h404fef10} /* (12, 6, 4) {real, imag} */,
  {32'h3d44e840, 32'h4062d935} /* (12, 6, 3) {real, imag} */,
  {32'hc0413ba0, 32'h3fa2c8d1} /* (12, 6, 2) {real, imag} */,
  {32'hc08e77f4, 32'hc0314047} /* (12, 6, 1) {real, imag} */,
  {32'hbfe0edff, 32'hbec7f58c} /* (12, 6, 0) {real, imag} */,
  {32'hbf848c01, 32'h3ff8444a} /* (12, 5, 31) {real, imag} */,
  {32'h3fb078b4, 32'h407833f3} /* (12, 5, 30) {real, imag} */,
  {32'hc06a7ba7, 32'h3ce30b00} /* (12, 5, 29) {real, imag} */,
  {32'hc0718c37, 32'hc1051cba} /* (12, 5, 28) {real, imag} */,
  {32'h400e5ea5, 32'hc10da7af} /* (12, 5, 27) {real, imag} */,
  {32'h40501231, 32'hbfc24cec} /* (12, 5, 26) {real, imag} */,
  {32'hc10cfbce, 32'h40c871a2} /* (12, 5, 25) {real, imag} */,
  {32'hbec37546, 32'h3fa16f64} /* (12, 5, 24) {real, imag} */,
  {32'h4149ebbd, 32'hc0177f3f} /* (12, 5, 23) {real, imag} */,
  {32'h3f2c715e, 32'h40c395ae} /* (12, 5, 22) {real, imag} */,
  {32'hc12a1d75, 32'h40ba60e2} /* (12, 5, 21) {real, imag} */,
  {32'hbfb64a08, 32'h3fa3bc3c} /* (12, 5, 20) {real, imag} */,
  {32'h3fb4feba, 32'h40cc1a48} /* (12, 5, 19) {real, imag} */,
  {32'h3fefb4a6, 32'hc10f032c} /* (12, 5, 18) {real, imag} */,
  {32'hbf3dfe14, 32'hc139d50c} /* (12, 5, 17) {real, imag} */,
  {32'hc057cd20, 32'hbea18840} /* (12, 5, 16) {real, imag} */,
  {32'hc10a5e28, 32'h4094326c} /* (12, 5, 15) {real, imag} */,
  {32'hc11950d8, 32'h408de13e} /* (12, 5, 14) {real, imag} */,
  {32'hc08d6d52, 32'hbe13cabe} /* (12, 5, 13) {real, imag} */,
  {32'hc0d63767, 32'h409ae66b} /* (12, 5, 12) {real, imag} */,
  {32'hc05e439c, 32'h410d25ca} /* (12, 5, 11) {real, imag} */,
  {32'h3e430ed0, 32'h415465d8} /* (12, 5, 10) {real, imag} */,
  {32'h400f1a28, 32'h40efdd88} /* (12, 5, 9) {real, imag} */,
  {32'h3fb07b98, 32'h3f8e42e8} /* (12, 5, 8) {real, imag} */,
  {32'h40282010, 32'hc0c76f14} /* (12, 5, 7) {real, imag} */,
  {32'hc0234632, 32'hc07d79b4} /* (12, 5, 6) {real, imag} */,
  {32'h3f7d71d4, 32'hc16666c0} /* (12, 5, 5) {real, imag} */,
  {32'h40d64450, 32'hc0d1d160} /* (12, 5, 4) {real, imag} */,
  {32'h41071c96, 32'hc1045811} /* (12, 5, 3) {real, imag} */,
  {32'h409c36e6, 32'hc183bd65} /* (12, 5, 2) {real, imag} */,
  {32'hbf4316f3, 32'hc04feb88} /* (12, 5, 1) {real, imag} */,
  {32'hc01db97a, 32'hbda90f40} /* (12, 5, 0) {real, imag} */,
  {32'hbf4d75ba, 32'hbf9a7535} /* (12, 4, 31) {real, imag} */,
  {32'hc095d472, 32'hc08675a2} /* (12, 4, 30) {real, imag} */,
  {32'h40a4d98a, 32'hc0933f2f} /* (12, 4, 29) {real, imag} */,
  {32'h40fe85aa, 32'hc12dfc52} /* (12, 4, 28) {real, imag} */,
  {32'h3f46d2b0, 32'hc10de0b6} /* (12, 4, 27) {real, imag} */,
  {32'h4078e0e2, 32'hbf0ad014} /* (12, 4, 26) {real, imag} */,
  {32'h40884873, 32'h4097cf0f} /* (12, 4, 25) {real, imag} */,
  {32'hbfd5b34c, 32'h40d473a1} /* (12, 4, 24) {real, imag} */,
  {32'hc0d424c6, 32'h4055d258} /* (12, 4, 23) {real, imag} */,
  {32'hc132fd9c, 32'hc06d9e95} /* (12, 4, 22) {real, imag} */,
  {32'hc12d5ac4, 32'hc0e3050d} /* (12, 4, 21) {real, imag} */,
  {32'hbfcda4ac, 32'h3d530180} /* (12, 4, 20) {real, imag} */,
  {32'hc0ce3859, 32'hc06b00d2} /* (12, 4, 19) {real, imag} */,
  {32'hbf91d650, 32'hc0ddebc0} /* (12, 4, 18) {real, imag} */,
  {32'h3d4b4980, 32'h3f9dfc08} /* (12, 4, 17) {real, imag} */,
  {32'hc08d88d5, 32'hbfb133fc} /* (12, 4, 16) {real, imag} */,
  {32'hc09ab018, 32'hc097a70b} /* (12, 4, 15) {real, imag} */,
  {32'hc0b64255, 32'h3f585248} /* (12, 4, 14) {real, imag} */,
  {32'hc02be6ef, 32'h40c1d1ff} /* (12, 4, 13) {real, imag} */,
  {32'h40a00e4e, 32'h407ddbb6} /* (12, 4, 12) {real, imag} */,
  {32'h4140f4e2, 32'h400d0720} /* (12, 4, 11) {real, imag} */,
  {32'hc00c1875, 32'hbd9b62f0} /* (12, 4, 10) {real, imag} */,
  {32'hc0a6d77a, 32'hbf6f25bd} /* (12, 4, 9) {real, imag} */,
  {32'hc1043186, 32'h3ed93bf8} /* (12, 4, 8) {real, imag} */,
  {32'hc118ac2f, 32'hc0ad4ce0} /* (12, 4, 7) {real, imag} */,
  {32'hc093e484, 32'hbf9d6c76} /* (12, 4, 6) {real, imag} */,
  {32'hc0587568, 32'hc00591d2} /* (12, 4, 5) {real, imag} */,
  {32'h3feaca17, 32'hc0aad78c} /* (12, 4, 4) {real, imag} */,
  {32'hbf8eeb52, 32'h4026f99b} /* (12, 4, 3) {real, imag} */,
  {32'hc0b36a2e, 32'hbeae2988} /* (12, 4, 2) {real, imag} */,
  {32'hc02f7de1, 32'h40c10199} /* (12, 4, 1) {real, imag} */,
  {32'h3ff244e8, 32'h4069add6} /* (12, 4, 0) {real, imag} */,
  {32'hc0353afb, 32'hbf0b43a5} /* (12, 3, 31) {real, imag} */,
  {32'h401d4230, 32'h40168f76} /* (12, 3, 30) {real, imag} */,
  {32'h410c2a3c, 32'hbf818802} /* (12, 3, 29) {real, imag} */,
  {32'h4042799c, 32'hc090a6d5} /* (12, 3, 28) {real, imag} */,
  {32'h402d9d6e, 32'hc0a014f6} /* (12, 3, 27) {real, imag} */,
  {32'h4045b393, 32'h405c8966} /* (12, 3, 26) {real, imag} */,
  {32'hbf5284e0, 32'h3ff0a340} /* (12, 3, 25) {real, imag} */,
  {32'hbf99e3e6, 32'h402f8710} /* (12, 3, 24) {real, imag} */,
  {32'hbf12ec7d, 32'hbe710300} /* (12, 3, 23) {real, imag} */,
  {32'hc0944c00, 32'h3fed2c8a} /* (12, 3, 22) {real, imag} */,
  {32'hc040040f, 32'h407faef8} /* (12, 3, 21) {real, imag} */,
  {32'hbfaa52b4, 32'h415bc926} /* (12, 3, 20) {real, imag} */,
  {32'h404453d8, 32'h4130638a} /* (12, 3, 19) {real, imag} */,
  {32'h4102422c, 32'h410db2e0} /* (12, 3, 18) {real, imag} */,
  {32'h40cca746, 32'h40c35aea} /* (12, 3, 17) {real, imag} */,
  {32'h4007d55a, 32'h3f4a8760} /* (12, 3, 16) {real, imag} */,
  {32'h3ecd0020, 32'hbf0e0c9c} /* (12, 3, 15) {real, imag} */,
  {32'hc136cf14, 32'hc0f046d2} /* (12, 3, 14) {real, imag} */,
  {32'hc10e5810, 32'hc0ad9f6a} /* (12, 3, 13) {real, imag} */,
  {32'h40b3dbfd, 32'hc0ff8f1c} /* (12, 3, 12) {real, imag} */,
  {32'h40356287, 32'hc1102772} /* (12, 3, 11) {real, imag} */,
  {32'hbfef1a64, 32'hc0cfdbcc} /* (12, 3, 10) {real, imag} */,
  {32'h3f2fcca2, 32'h40c24bd4} /* (12, 3, 9) {real, imag} */,
  {32'h401647c8, 32'h409aa186} /* (12, 3, 8) {real, imag} */,
  {32'h3f9d1c80, 32'h40100ab6} /* (12, 3, 7) {real, imag} */,
  {32'h4090c779, 32'hbfbfe3ec} /* (12, 3, 6) {real, imag} */,
  {32'h401a278a, 32'hc109e036} /* (12, 3, 5) {real, imag} */,
  {32'h4046920a, 32'hc0c9ea0b} /* (12, 3, 4) {real, imag} */,
  {32'h40c74af5, 32'hc0582dbe} /* (12, 3, 3) {real, imag} */,
  {32'h3fc4d182, 32'h407a4882} /* (12, 3, 2) {real, imag} */,
  {32'h3f93d1e4, 32'hc08ce25e} /* (12, 3, 1) {real, imag} */,
  {32'h409c3bd2, 32'hbf280700} /* (12, 3, 0) {real, imag} */,
  {32'hc08ac7c5, 32'hbe360e46} /* (12, 2, 31) {real, imag} */,
  {32'h408713ba, 32'h40835145} /* (12, 2, 30) {real, imag} */,
  {32'h3e59cd60, 32'h3fcc658c} /* (12, 2, 29) {real, imag} */,
  {32'h3f3500b3, 32'hbe48fe70} /* (12, 2, 28) {real, imag} */,
  {32'hbee0f4a8, 32'hbf187d5c} /* (12, 2, 27) {real, imag} */,
  {32'h41319411, 32'hbfdd6878} /* (12, 2, 26) {real, imag} */,
  {32'h413eb510, 32'hc1096033} /* (12, 2, 25) {real, imag} */,
  {32'h416a6b9d, 32'hc085a184} /* (12, 2, 24) {real, imag} */,
  {32'h403717c8, 32'h40add2fb} /* (12, 2, 23) {real, imag} */,
  {32'hc06f0114, 32'hc082d7c4} /* (12, 2, 22) {real, imag} */,
  {32'h40574885, 32'h3e88aca8} /* (12, 2, 21) {real, imag} */,
  {32'hbff65480, 32'hc06e03dc} /* (12, 2, 20) {real, imag} */,
  {32'hc027bb5c, 32'hc00a8c44} /* (12, 2, 19) {real, imag} */,
  {32'hbfcdb5af, 32'h403b482d} /* (12, 2, 18) {real, imag} */,
  {32'hc09cdd4d, 32'h40421a0d} /* (12, 2, 17) {real, imag} */,
  {32'hc0f28524, 32'h3f7235d0} /* (12, 2, 16) {real, imag} */,
  {32'h4040318c, 32'h3fe06ba4} /* (12, 2, 15) {real, imag} */,
  {32'hbf1cf88d, 32'hc01395c0} /* (12, 2, 14) {real, imag} */,
  {32'hc04c88e4, 32'h4046b553} /* (12, 2, 13) {real, imag} */,
  {32'hbfac476d, 32'h41843b3a} /* (12, 2, 12) {real, imag} */,
  {32'hc11d7d7b, 32'h411b3de2} /* (12, 2, 11) {real, imag} */,
  {32'hbfce3dfc, 32'hc0d7b43a} /* (12, 2, 10) {real, imag} */,
  {32'h3f7bac97, 32'hc18ba996} /* (12, 2, 9) {real, imag} */,
  {32'hc1041e85, 32'hc0a7c498} /* (12, 2, 8) {real, imag} */,
  {32'hc123c697, 32'h3f929f9c} /* (12, 2, 7) {real, imag} */,
  {32'hc0e3cf74, 32'h40ddbb43} /* (12, 2, 6) {real, imag} */,
  {32'h404bfe89, 32'h407b5072} /* (12, 2, 5) {real, imag} */,
  {32'hc008471f, 32'hbfea4562} /* (12, 2, 4) {real, imag} */,
  {32'hc0e47922, 32'h4020f024} /* (12, 2, 3) {real, imag} */,
  {32'hbd5db940, 32'h40f68e96} /* (12, 2, 2) {real, imag} */,
  {32'h40b3f7ad, 32'h40a8ad60} /* (12, 2, 1) {real, imag} */,
  {32'hc045cbcc, 32'hc0257501} /* (12, 2, 0) {real, imag} */,
  {32'h40927f7b, 32'hbfb7458c} /* (12, 1, 31) {real, imag} */,
  {32'h41340956, 32'hc0f9ab78} /* (12, 1, 30) {real, imag} */,
  {32'h410a3ee6, 32'hc0e551f6} /* (12, 1, 29) {real, imag} */,
  {32'h4027451c, 32'h3fbe73ed} /* (12, 1, 28) {real, imag} */,
  {32'hbf7b9978, 32'hbf7a2252} /* (12, 1, 27) {real, imag} */,
  {32'hc0843346, 32'hbfc34b66} /* (12, 1, 26) {real, imag} */,
  {32'hc10ebee0, 32'h3f850bd0} /* (12, 1, 25) {real, imag} */,
  {32'hc01b27ba, 32'h3fa005d8} /* (12, 1, 24) {real, imag} */,
  {32'hbfe08cef, 32'h3e546400} /* (12, 1, 23) {real, imag} */,
  {32'hc0cac39c, 32'hbe083a00} /* (12, 1, 22) {real, imag} */,
  {32'h40a70144, 32'h405f4c25} /* (12, 1, 21) {real, imag} */,
  {32'h414cbad5, 32'hc00ca9c7} /* (12, 1, 20) {real, imag} */,
  {32'h40b5d20c, 32'hc0d8f52d} /* (12, 1, 19) {real, imag} */,
  {32'h40e8c5de, 32'hc0a156e6} /* (12, 1, 18) {real, imag} */,
  {32'h40c21526, 32'hbf4d2908} /* (12, 1, 17) {real, imag} */,
  {32'hc01c42b2, 32'hbeabd230} /* (12, 1, 16) {real, imag} */,
  {32'h3fb77579, 32'hc08b5b29} /* (12, 1, 15) {real, imag} */,
  {32'h3bd88400, 32'h3f545254} /* (12, 1, 14) {real, imag} */,
  {32'h403da618, 32'h40eda037} /* (12, 1, 13) {real, imag} */,
  {32'h40eba633, 32'h40256502} /* (12, 1, 12) {real, imag} */,
  {32'h3ff14a9c, 32'hc0338bba} /* (12, 1, 11) {real, imag} */,
  {32'h40d2f75d, 32'h3fbe7b00} /* (12, 1, 10) {real, imag} */,
  {32'hbf365db4, 32'h40c68aa9} /* (12, 1, 9) {real, imag} */,
  {32'hc0f40855, 32'h40fa0836} /* (12, 1, 8) {real, imag} */,
  {32'hc10afe98, 32'h40540d06} /* (12, 1, 7) {real, imag} */,
  {32'hc105e55c, 32'h401fd61c} /* (12, 1, 6) {real, imag} */,
  {32'h3fab213a, 32'hbf5cc390} /* (12, 1, 5) {real, imag} */,
  {32'h4185ec12, 32'hbefbd7b0} /* (12, 1, 4) {real, imag} */,
  {32'h4112a76c, 32'hc065d586} /* (12, 1, 3) {real, imag} */,
  {32'h403c3d4f, 32'hc0028836} /* (12, 1, 2) {real, imag} */,
  {32'hc07b004b, 32'h40dee045} /* (12, 1, 1) {real, imag} */,
  {32'hbf964223, 32'h40ae111d} /* (12, 1, 0) {real, imag} */,
  {32'hc052f0f7, 32'hbf1e0acc} /* (12, 0, 31) {real, imag} */,
  {32'hc07cd8ea, 32'h40333e1c} /* (12, 0, 30) {real, imag} */,
  {32'hbfc99eb8, 32'hbf10d7fc} /* (12, 0, 29) {real, imag} */,
  {32'hbfe991c6, 32'h3f07f09f} /* (12, 0, 28) {real, imag} */,
  {32'hbf7611d0, 32'hc0b34cf6} /* (12, 0, 27) {real, imag} */,
  {32'h40be7620, 32'hc0fc79c2} /* (12, 0, 26) {real, imag} */,
  {32'h412270b2, 32'hc1318425} /* (12, 0, 25) {real, imag} */,
  {32'hbeff4368, 32'hbff331ba} /* (12, 0, 24) {real, imag} */,
  {32'hc0efe8e6, 32'h40b7a37e} /* (12, 0, 23) {real, imag} */,
  {32'hc10c558e, 32'hc02dd470} /* (12, 0, 22) {real, imag} */,
  {32'hc0597b22, 32'hc09f6f2f} /* (12, 0, 21) {real, imag} */,
  {32'hc09e070d, 32'hc10f1b37} /* (12, 0, 20) {real, imag} */,
  {32'hc02cd8a8, 32'h402d6636} /* (12, 0, 19) {real, imag} */,
  {32'hc1158562, 32'h412836c9} /* (12, 0, 18) {real, imag} */,
  {32'hbfd75a3e, 32'h409f170d} /* (12, 0, 17) {real, imag} */,
  {32'h40cc8094, 32'h40a5b694} /* (12, 0, 16) {real, imag} */,
  {32'h3e5e0304, 32'hbf478a33} /* (12, 0, 15) {real, imag} */,
  {32'hc0da3c9a, 32'hc1401628} /* (12, 0, 14) {real, imag} */,
  {32'hc11448e6, 32'hc111a106} /* (12, 0, 13) {real, imag} */,
  {32'h408304b6, 32'h40598d2c} /* (12, 0, 12) {real, imag} */,
  {32'h40cc94d8, 32'h409446fb} /* (12, 0, 11) {real, imag} */,
  {32'h410b4818, 32'hbf8b01fc} /* (12, 0, 10) {real, imag} */,
  {32'h402cd3bc, 32'h3fc81365} /* (12, 0, 9) {real, imag} */,
  {32'hbf4eb694, 32'hc047449c} /* (12, 0, 8) {real, imag} */,
  {32'h3f153224, 32'hc0169a12} /* (12, 0, 7) {real, imag} */,
  {32'hc003b114, 32'hc0c44d70} /* (12, 0, 6) {real, imag} */,
  {32'h40c867de, 32'h3ead9f4e} /* (12, 0, 5) {real, imag} */,
  {32'h40efd17c, 32'h40b188fc} /* (12, 0, 4) {real, imag} */,
  {32'hc135e443, 32'hc0c4a3e8} /* (12, 0, 3) {real, imag} */,
  {32'hc17bed05, 32'hc0964c08} /* (12, 0, 2) {real, imag} */,
  {32'hbf03ff18, 32'hbf8f674f} /* (12, 0, 1) {real, imag} */,
  {32'h4088863e, 32'hc0cd5520} /* (12, 0, 0) {real, imag} */,
  {32'h4116738e, 32'hc123975b} /* (11, 31, 31) {real, imag} */,
  {32'h415aee21, 32'hc137d7b7} /* (11, 31, 30) {real, imag} */,
  {32'hbfb37368, 32'hc1194459} /* (11, 31, 29) {real, imag} */,
  {32'h4115429c, 32'hc16c40cd} /* (11, 31, 28) {real, imag} */,
  {32'h412bd7f8, 32'hc1079620} /* (11, 31, 27) {real, imag} */,
  {32'h40ace5ff, 32'hc019f01e} /* (11, 31, 26) {real, imag} */,
  {32'h40246370, 32'hc193a824} /* (11, 31, 25) {real, imag} */,
  {32'h4168b894, 32'hc1dc32b2} /* (11, 31, 24) {real, imag} */,
  {32'h41522d4e, 32'hc19567c4} /* (11, 31, 23) {real, imag} */,
  {32'h4146cbf4, 32'hc13bef54} /* (11, 31, 22) {real, imag} */,
  {32'h41268bac, 32'hbfad48b0} /* (11, 31, 21) {real, imag} */,
  {32'h40c6c578, 32'h411c9590} /* (11, 31, 20) {real, imag} */,
  {32'hc08e2f22, 32'h41269cea} /* (11, 31, 19) {real, imag} */,
  {32'hbf2f5a00, 32'h4137de12} /* (11, 31, 18) {real, imag} */,
  {32'h406592b8, 32'h40df3ab7} /* (11, 31, 17) {real, imag} */,
  {32'hc123a8c5, 32'h40fbf00f} /* (11, 31, 16) {real, imag} */,
  {32'hc0f07936, 32'h405bec65} /* (11, 31, 15) {real, imag} */,
  {32'hc10fc69a, 32'h401c6971} /* (11, 31, 14) {real, imag} */,
  {32'hbf0551a0, 32'hbf8866f6} /* (11, 31, 13) {real, imag} */,
  {32'hc06fc7c7, 32'h40131b8c} /* (11, 31, 12) {real, imag} */,
  {32'hbfe7d5b8, 32'h4039b256} /* (11, 31, 11) {real, imag} */,
  {32'h410dafce, 32'hc1b8af46} /* (11, 31, 10) {real, imag} */,
  {32'hc0f47920, 32'hc204ae3d} /* (11, 31, 9) {real, imag} */,
  {32'hc16eac16, 32'hc1c21050} /* (11, 31, 8) {real, imag} */,
  {32'hc08168da, 32'hc1953bd0} /* (11, 31, 7) {real, imag} */,
  {32'h4093f70b, 32'hc1b3eff4} /* (11, 31, 6) {real, imag} */,
  {32'h418721e7, 32'hc13846f4} /* (11, 31, 5) {real, imag} */,
  {32'h41a86e80, 32'h3e6fbb00} /* (11, 31, 4) {real, imag} */,
  {32'h41542364, 32'hbfbc7990} /* (11, 31, 3) {real, imag} */,
  {32'h3ff8f9c0, 32'h400d3ff4} /* (11, 31, 2) {real, imag} */,
  {32'h413564dc, 32'hc05c266e} /* (11, 31, 1) {real, imag} */,
  {32'h413879c5, 32'hc042cdfe} /* (11, 31, 0) {real, imag} */,
  {32'hbecb1040, 32'h4136e077} /* (11, 30, 31) {real, imag} */,
  {32'hc0a46239, 32'h4156f001} /* (11, 30, 30) {real, imag} */,
  {32'hc1140710, 32'h41650baf} /* (11, 30, 29) {real, imag} */,
  {32'hc0c00283, 32'h41350b53} /* (11, 30, 28) {real, imag} */,
  {32'hc0dceb64, 32'h404f5440} /* (11, 30, 27) {real, imag} */,
  {32'hc0bd776c, 32'h3fdf8c2d} /* (11, 30, 26) {real, imag} */,
  {32'hc0fd9f8c, 32'h413d3a10} /* (11, 30, 25) {real, imag} */,
  {32'hc14a5f5d, 32'h414baa85} /* (11, 30, 24) {real, imag} */,
  {32'hc125c144, 32'h40f16801} /* (11, 30, 23) {real, imag} */,
  {32'hc1271da6, 32'h41128198} /* (11, 30, 22) {real, imag} */,
  {32'hc1172f6c, 32'h41158c1b} /* (11, 30, 21) {real, imag} */,
  {32'h414b470e, 32'h40e2edba} /* (11, 30, 20) {real, imag} */,
  {32'h4169d941, 32'h401acfe8} /* (11, 30, 19) {real, imag} */,
  {32'h41949b31, 32'hc017dcc0} /* (11, 30, 18) {real, imag} */,
  {32'h41b9cdb0, 32'hc1033a85} /* (11, 30, 17) {real, imag} */,
  {32'h41aba84e, 32'hc091d42f} /* (11, 30, 16) {real, imag} */,
  {32'h418a5f60, 32'h3f839691} /* (11, 30, 15) {real, imag} */,
  {32'h40b71648, 32'hbfe8efaa} /* (11, 30, 14) {real, imag} */,
  {32'h409f5325, 32'hbdd0c810} /* (11, 30, 13) {real, imag} */,
  {32'hc113139f, 32'hc132d5ac} /* (11, 30, 12) {real, imag} */,
  {32'hc1290502, 32'hc17eac26} /* (11, 30, 11) {real, imag} */,
  {32'hc0229b88, 32'h402f347c} /* (11, 30, 10) {real, imag} */,
  {32'h3ee2e880, 32'hbccfc000} /* (11, 30, 9) {real, imag} */,
  {32'hc0cfa109, 32'h408dd1ca} /* (11, 30, 8) {real, imag} */,
  {32'hc0f585c2, 32'h410297ee} /* (11, 30, 7) {real, imag} */,
  {32'hc181050c, 32'h4112fb8a} /* (11, 30, 6) {real, imag} */,
  {32'hc0d3f408, 32'h40cd27ab} /* (11, 30, 5) {real, imag} */,
  {32'h40b9e819, 32'h4020021e} /* (11, 30, 4) {real, imag} */,
  {32'hbe3646b0, 32'h40a673cd} /* (11, 30, 3) {real, imag} */,
  {32'hc0f79dad, 32'h41170e19} /* (11, 30, 2) {real, imag} */,
  {32'hc10b3bf8, 32'hc0c43312} /* (11, 30, 1) {real, imag} */,
  {32'h4020d9c2, 32'hc0670c45} /* (11, 30, 0) {real, imag} */,
  {32'h40be7f44, 32'h40ce6a7b} /* (11, 29, 31) {real, imag} */,
  {32'h4078140a, 32'h403c456a} /* (11, 29, 30) {real, imag} */,
  {32'hbf17a7c1, 32'h4089ad65} /* (11, 29, 29) {real, imag} */,
  {32'hbfb0bafc, 32'h40c55b12} /* (11, 29, 28) {real, imag} */,
  {32'h4009c984, 32'h40343bda} /* (11, 29, 27) {real, imag} */,
  {32'h40c21664, 32'hc1417587} /* (11, 29, 26) {real, imag} */,
  {32'h4055f81e, 32'hc0a1b5c5} /* (11, 29, 25) {real, imag} */,
  {32'hc02c5865, 32'hbd9990a0} /* (11, 29, 24) {real, imag} */,
  {32'hbec269c0, 32'h401e6806} /* (11, 29, 23) {real, imag} */,
  {32'h406b60db, 32'hc095b5af} /* (11, 29, 22) {real, imag} */,
  {32'hc041d7c4, 32'hc0a9664d} /* (11, 29, 21) {real, imag} */,
  {32'h4079fa3c, 32'h40fb9e63} /* (11, 29, 20) {real, imag} */,
  {32'h402a0ea0, 32'h40cebc1a} /* (11, 29, 19) {real, imag} */,
  {32'h40953fe3, 32'h40f62174} /* (11, 29, 18) {real, imag} */,
  {32'h4091cc12, 32'h412dee12} /* (11, 29, 17) {real, imag} */,
  {32'h3f8b930c, 32'h411f63bd} /* (11, 29, 16) {real, imag} */,
  {32'hc077cdb5, 32'h4145cc74} /* (11, 29, 15) {real, imag} */,
  {32'hbfca35c0, 32'h41497db5} /* (11, 29, 14) {real, imag} */,
  {32'h41310cff, 32'h416f2423} /* (11, 29, 13) {real, imag} */,
  {32'h409776fa, 32'h402cbd01} /* (11, 29, 12) {real, imag} */,
  {32'hc132c205, 32'h3ff85244} /* (11, 29, 11) {real, imag} */,
  {32'h3f7b76a8, 32'hbf353e60} /* (11, 29, 10) {real, imag} */,
  {32'hc08c20a0, 32'h3fb076be} /* (11, 29, 9) {real, imag} */,
  {32'hc027f83a, 32'hc15cd4df} /* (11, 29, 8) {real, imag} */,
  {32'h3f8daf30, 32'hc1852fa0} /* (11, 29, 7) {real, imag} */,
  {32'h4084f537, 32'hc1860317} /* (11, 29, 6) {real, imag} */,
  {32'hc02fb21b, 32'hc045d9b3} /* (11, 29, 5) {real, imag} */,
  {32'hc0eee958, 32'h40d34353} /* (11, 29, 4) {real, imag} */,
  {32'hc0b78959, 32'h40b6912e} /* (11, 29, 3) {real, imag} */,
  {32'hbef760fc, 32'hc0c00517} /* (11, 29, 2) {real, imag} */,
  {32'hbe2c8920, 32'h3ff5c446} /* (11, 29, 1) {real, imag} */,
  {32'h4093859d, 32'h3f3264dc} /* (11, 29, 0) {real, imag} */,
  {32'h40aec1cc, 32'hc023fcc6} /* (11, 28, 31) {real, imag} */,
  {32'h405d556c, 32'h4093561b} /* (11, 28, 30) {real, imag} */,
  {32'h3f3ff2c8, 32'h40d0d005} /* (11, 28, 29) {real, imag} */,
  {32'hbfb14083, 32'h4137a60c} /* (11, 28, 28) {real, imag} */,
  {32'hbf036674, 32'h41586d90} /* (11, 28, 27) {real, imag} */,
  {32'h40bb8c64, 32'h40e5d65a} /* (11, 28, 26) {real, imag} */,
  {32'h40042030, 32'h415734d8} /* (11, 28, 25) {real, imag} */,
  {32'h4053ff34, 32'h415b668b} /* (11, 28, 24) {real, imag} */,
  {32'h3e12b580, 32'hc119550e} /* (11, 28, 23) {real, imag} */,
  {32'h3fb6758e, 32'hc14778fc} /* (11, 28, 22) {real, imag} */,
  {32'hc007ea22, 32'hc128d3aa} /* (11, 28, 21) {real, imag} */,
  {32'hc0ba6f28, 32'hc03cabda} /* (11, 28, 20) {real, imag} */,
  {32'hc042ed1b, 32'hc0fae54e} /* (11, 28, 19) {real, imag} */,
  {32'hc0738240, 32'hc0d1f61f} /* (11, 28, 18) {real, imag} */,
  {32'hc09494fb, 32'hbfa90a38} /* (11, 28, 17) {real, imag} */,
  {32'hc0849fa6, 32'h40fcac7a} /* (11, 28, 16) {real, imag} */,
  {32'hc01e2d4e, 32'h40d6416a} /* (11, 28, 15) {real, imag} */,
  {32'h40934fc0, 32'h41033356} /* (11, 28, 14) {real, imag} */,
  {32'h401e46e0, 32'h40082b2c} /* (11, 28, 13) {real, imag} */,
  {32'h40bb1f70, 32'h4009679c} /* (11, 28, 12) {real, imag} */,
  {32'h3fcdefd5, 32'hc0b471e8} /* (11, 28, 11) {real, imag} */,
  {32'h40bbad8e, 32'hc0da28ba} /* (11, 28, 10) {real, imag} */,
  {32'hc038e65c, 32'hbfdc79ea} /* (11, 28, 9) {real, imag} */,
  {32'hc15f2d40, 32'hc0a0639e} /* (11, 28, 8) {real, imag} */,
  {32'hc12664ab, 32'hc0896bec} /* (11, 28, 7) {real, imag} */,
  {32'h40859b38, 32'hc03c7958} /* (11, 28, 6) {real, imag} */,
  {32'h4078a42d, 32'hbfca4e48} /* (11, 28, 5) {real, imag} */,
  {32'hc06b0a2c, 32'h3fd8b20e} /* (11, 28, 4) {real, imag} */,
  {32'hbf238166, 32'h3f94e346} /* (11, 28, 3) {real, imag} */,
  {32'h40829dbe, 32'h3fb4073f} /* (11, 28, 2) {real, imag} */,
  {32'h407f1f48, 32'hc12e9407} /* (11, 28, 1) {real, imag} */,
  {32'h40497772, 32'hc11c37a1} /* (11, 28, 0) {real, imag} */,
  {32'hc0bcff19, 32'h3f861afc} /* (11, 27, 31) {real, imag} */,
  {32'hc0eb2ef5, 32'h402aca96} /* (11, 27, 30) {real, imag} */,
  {32'hc134157c, 32'h3fad2180} /* (11, 27, 29) {real, imag} */,
  {32'hc0d8a872, 32'h4064d21f} /* (11, 27, 28) {real, imag} */,
  {32'hc0fdf47b, 32'h407d5ffb} /* (11, 27, 27) {real, imag} */,
  {32'hc03bbe20, 32'h3fca4a0e} /* (11, 27, 26) {real, imag} */,
  {32'h3f04d898, 32'h410821b2} /* (11, 27, 25) {real, imag} */,
  {32'hc0882e06, 32'h4136cc97} /* (11, 27, 24) {real, imag} */,
  {32'hc169f3be, 32'h414ca8ca} /* (11, 27, 23) {real, imag} */,
  {32'hc0578c54, 32'h41031441} /* (11, 27, 22) {real, imag} */,
  {32'h40c46fe6, 32'h410dd288} /* (11, 27, 21) {real, imag} */,
  {32'h40e8668e, 32'hc00ad860} /* (11, 27, 20) {real, imag} */,
  {32'h4035a95a, 32'hc0afd7f7} /* (11, 27, 19) {real, imag} */,
  {32'h3ff28be6, 32'hbfe6b636} /* (11, 27, 18) {real, imag} */,
  {32'h40113a9e, 32'h3fd05fc2} /* (11, 27, 17) {real, imag} */,
  {32'hc06d800e, 32'hc01cbc2a} /* (11, 27, 16) {real, imag} */,
  {32'hc0d67b92, 32'hc09adcd6} /* (11, 27, 15) {real, imag} */,
  {32'hc083faf7, 32'hc10a98a5} /* (11, 27, 14) {real, imag} */,
  {32'h3fa8139e, 32'hc1177789} /* (11, 27, 13) {real, imag} */,
  {32'h3f9f03f0, 32'h404c6273} /* (11, 27, 12) {real, imag} */,
  {32'hc0f12cd2, 32'h412e476c} /* (11, 27, 11) {real, imag} */,
  {32'hc116aaef, 32'h3f403e38} /* (11, 27, 10) {real, imag} */,
  {32'h404ce9a1, 32'hbdfe5380} /* (11, 27, 9) {real, imag} */,
  {32'h414b8a36, 32'h408b3aa2} /* (11, 27, 8) {real, imag} */,
  {32'h41079499, 32'h406423c4} /* (11, 27, 7) {real, imag} */,
  {32'hc0306da5, 32'h417b95fd} /* (11, 27, 6) {real, imag} */,
  {32'hbd49b5c0, 32'h416e587c} /* (11, 27, 5) {real, imag} */,
  {32'h4092c06f, 32'h41425d02} /* (11, 27, 4) {real, imag} */,
  {32'h401c6f24, 32'h409934b9} /* (11, 27, 3) {real, imag} */,
  {32'hc08e1933, 32'h3f8dbaea} /* (11, 27, 2) {real, imag} */,
  {32'hc0a71bb8, 32'hc093888e} /* (11, 27, 1) {real, imag} */,
  {32'hbf091f44, 32'hbe9c7a78} /* (11, 27, 0) {real, imag} */,
  {32'hc01e4faa, 32'hbfcd3a08} /* (11, 26, 31) {real, imag} */,
  {32'hc10388cc, 32'h409d0424} /* (11, 26, 30) {real, imag} */,
  {32'hbfa57744, 32'h4090e433} /* (11, 26, 29) {real, imag} */,
  {32'h410d6534, 32'hc0cb4cb8} /* (11, 26, 28) {real, imag} */,
  {32'h412e482f, 32'hc11b8ecd} /* (11, 26, 27) {real, imag} */,
  {32'h4113a0f5, 32'h3fdba798} /* (11, 26, 26) {real, imag} */,
  {32'h412e6ff8, 32'h40cc5bb5} /* (11, 26, 25) {real, imag} */,
  {32'h40f07970, 32'h4084317c} /* (11, 26, 24) {real, imag} */,
  {32'h3e6771e0, 32'h41403c51} /* (11, 26, 23) {real, imag} */,
  {32'h40771da7, 32'h417f264a} /* (11, 26, 22) {real, imag} */,
  {32'h4090a356, 32'h40bb2189} /* (11, 26, 21) {real, imag} */,
  {32'hc07ed2ec, 32'h3eb549fe} /* (11, 26, 20) {real, imag} */,
  {32'hc0e963a1, 32'h3f9a47d0} /* (11, 26, 19) {real, imag} */,
  {32'h3fc0c042, 32'hbf911c7c} /* (11, 26, 18) {real, imag} */,
  {32'h40d6bc3c, 32'h4072389f} /* (11, 26, 17) {real, imag} */,
  {32'h3fc54d48, 32'hc0c381a0} /* (11, 26, 16) {real, imag} */,
  {32'h3d42a700, 32'hc0533a9c} /* (11, 26, 15) {real, imag} */,
  {32'h3eab5a88, 32'hc0499d4a} /* (11, 26, 14) {real, imag} */,
  {32'hbebbc6a0, 32'hbffd6a69} /* (11, 26, 13) {real, imag} */,
  {32'hc018a9f6, 32'h40a0a35a} /* (11, 26, 12) {real, imag} */,
  {32'hbf290fe0, 32'h400f6559} /* (11, 26, 11) {real, imag} */,
  {32'h405522b2, 32'h400263f8} /* (11, 26, 10) {real, imag} */,
  {32'h40de5bfe, 32'h3fab4638} /* (11, 26, 9) {real, imag} */,
  {32'hbecea948, 32'h4126b7c3} /* (11, 26, 8) {real, imag} */,
  {32'hbfc684ca, 32'hbf50f864} /* (11, 26, 7) {real, imag} */,
  {32'hbf63b7a4, 32'h409ba855} /* (11, 26, 6) {real, imag} */,
  {32'hbff41176, 32'h402adf4b} /* (11, 26, 5) {real, imag} */,
  {32'hbebb2050, 32'hbef693a0} /* (11, 26, 4) {real, imag} */,
  {32'h3fd300d6, 32'h3fb9389c} /* (11, 26, 3) {real, imag} */,
  {32'hc087c0c9, 32'hc090e885} /* (11, 26, 2) {real, imag} */,
  {32'hbf7f1a5e, 32'hc05a690c} /* (11, 26, 1) {real, imag} */,
  {32'h3fa10a2e, 32'hc0044299} /* (11, 26, 0) {real, imag} */,
  {32'hc0340779, 32'hc096f8fe} /* (11, 25, 31) {real, imag} */,
  {32'hc002570e, 32'h3edbd2d8} /* (11, 25, 30) {real, imag} */,
  {32'h40ce4774, 32'h40369b70} /* (11, 25, 29) {real, imag} */,
  {32'h3f9e6536, 32'h40767264} /* (11, 25, 28) {real, imag} */,
  {32'hbf3fdae0, 32'h402f8bae} /* (11, 25, 27) {real, imag} */,
  {32'hbea4131c, 32'h3fdaab84} /* (11, 25, 26) {real, imag} */,
  {32'hbf5571e6, 32'hbf9a84f8} /* (11, 25, 25) {real, imag} */,
  {32'h40a9095c, 32'h40d6eea9} /* (11, 25, 24) {real, imag} */,
  {32'h40d07418, 32'h412b776c} /* (11, 25, 23) {real, imag} */,
  {32'h3da37180, 32'h405fc1fb} /* (11, 25, 22) {real, imag} */,
  {32'h3e0a6338, 32'h408d0f3a} /* (11, 25, 21) {real, imag} */,
  {32'h406c5e02, 32'h3fb3535f} /* (11, 25, 20) {real, imag} */,
  {32'hbe629140, 32'h3fe6fe94} /* (11, 25, 19) {real, imag} */,
  {32'h3e953420, 32'hc044153d} /* (11, 25, 18) {real, imag} */,
  {32'h40b26600, 32'h3f80b8c2} /* (11, 25, 17) {real, imag} */,
  {32'h4078d146, 32'hc04da466} /* (11, 25, 16) {real, imag} */,
  {32'h3e047400, 32'hbfe4ef01} /* (11, 25, 15) {real, imag} */,
  {32'h3f4afb2e, 32'hbfd9fac6} /* (11, 25, 14) {real, imag} */,
  {32'h41208371, 32'hbf4350e0} /* (11, 25, 13) {real, imag} */,
  {32'h3febb216, 32'hc05c066e} /* (11, 25, 12) {real, imag} */,
  {32'hc0b1cdeb, 32'hc042a4cf} /* (11, 25, 11) {real, imag} */,
  {32'hc05e6270, 32'h40a16b54} /* (11, 25, 10) {real, imag} */,
  {32'hc02e1c48, 32'h40ba7b42} /* (11, 25, 9) {real, imag} */,
  {32'h41086095, 32'h404ad031} /* (11, 25, 8) {real, imag} */,
  {32'h40b7a485, 32'hc066a905} /* (11, 25, 7) {real, imag} */,
  {32'h3fef4c5c, 32'hc0ac5249} /* (11, 25, 6) {real, imag} */,
  {32'h3fb2d782, 32'hc0604f80} /* (11, 25, 5) {real, imag} */,
  {32'h3f1660b8, 32'h3ff933be} /* (11, 25, 4) {real, imag} */,
  {32'h3fb59564, 32'hbe20d890} /* (11, 25, 3) {real, imag} */,
  {32'h40df899d, 32'h40a1cef1} /* (11, 25, 2) {real, imag} */,
  {32'h40980c3c, 32'h40034e4b} /* (11, 25, 1) {real, imag} */,
  {32'h3d92ea10, 32'hc00a2949} /* (11, 25, 0) {real, imag} */,
  {32'h40702827, 32'h3ef9bdc8} /* (11, 24, 31) {real, imag} */,
  {32'h3f13ce04, 32'h3e508c10} /* (11, 24, 30) {real, imag} */,
  {32'hc108a282, 32'h40b16834} /* (11, 24, 29) {real, imag} */,
  {32'hc0d6db50, 32'h40fd14be} /* (11, 24, 28) {real, imag} */,
  {32'h3fcda112, 32'hc0b02de3} /* (11, 24, 27) {real, imag} */,
  {32'h406f4cde, 32'hc03808f9} /* (11, 24, 26) {real, imag} */,
  {32'h3f865f17, 32'h3f9c6f68} /* (11, 24, 25) {real, imag} */,
  {32'hbfcc6178, 32'h404bae42} /* (11, 24, 24) {real, imag} */,
  {32'hc01e1fbc, 32'h403acc11} /* (11, 24, 23) {real, imag} */,
  {32'h405c89ca, 32'h4080e2a5} /* (11, 24, 22) {real, imag} */,
  {32'hc012677c, 32'hbe2647b0} /* (11, 24, 21) {real, imag} */,
  {32'hbf3d87da, 32'hbf6147fc} /* (11, 24, 20) {real, imag} */,
  {32'h3fa2c828, 32'h4071b600} /* (11, 24, 19) {real, imag} */,
  {32'h405ee1c7, 32'h4133c980} /* (11, 24, 18) {real, imag} */,
  {32'h40bb6d6e, 32'h412dc796} /* (11, 24, 17) {real, imag} */,
  {32'h3e493f88, 32'h40a4ccb8} /* (11, 24, 16) {real, imag} */,
  {32'hc0d2175b, 32'hc0534506} /* (11, 24, 15) {real, imag} */,
  {32'hc0f0b7e8, 32'hc0101c5e} /* (11, 24, 14) {real, imag} */,
  {32'hbd2ef680, 32'hc027934a} /* (11, 24, 13) {real, imag} */,
  {32'h406f017c, 32'hc059c672} /* (11, 24, 12) {real, imag} */,
  {32'hc02ac672, 32'hc03b4e0f} /* (11, 24, 11) {real, imag} */,
  {32'h3f231606, 32'hbe8b2bf8} /* (11, 24, 10) {real, imag} */,
  {32'h3f6450fc, 32'hbffcb246} /* (11, 24, 9) {real, imag} */,
  {32'hc031faa8, 32'hc06defa5} /* (11, 24, 8) {real, imag} */,
  {32'hc0a2f644, 32'h4036cb17} /* (11, 24, 7) {real, imag} */,
  {32'hc0b9ef43, 32'h4136a4be} /* (11, 24, 6) {real, imag} */,
  {32'hc0e59640, 32'h4086b171} /* (11, 24, 5) {real, imag} */,
  {32'hc0dea6d8, 32'h3f8d2d77} /* (11, 24, 4) {real, imag} */,
  {32'hc100f506, 32'h40d08fc4} /* (11, 24, 3) {real, imag} */,
  {32'hc02e050b, 32'h411ccc76} /* (11, 24, 2) {real, imag} */,
  {32'hc06d20c8, 32'h411d83fb} /* (11, 24, 1) {real, imag} */,
  {32'hbf4a82b2, 32'h4080dd7d} /* (11, 24, 0) {real, imag} */,
  {32'hc02e71de, 32'hbe84d9c8} /* (11, 23, 31) {real, imag} */,
  {32'hc091eb70, 32'h3ffb19e8} /* (11, 23, 30) {real, imag} */,
  {32'h3e2772a4, 32'h404f420b} /* (11, 23, 29) {real, imag} */,
  {32'h404dd82b, 32'h40a131bc} /* (11, 23, 28) {real, imag} */,
  {32'h3e9554c0, 32'hc0316026} /* (11, 23, 27) {real, imag} */,
  {32'hbf9cddec, 32'hc0f04380} /* (11, 23, 26) {real, imag} */,
  {32'h3fa58c2b, 32'hc087cd09} /* (11, 23, 25) {real, imag} */,
  {32'h3f82611f, 32'hbf6f94e0} /* (11, 23, 24) {real, imag} */,
  {32'hbfe3ffb4, 32'hbf01aad4} /* (11, 23, 23) {real, imag} */,
  {32'h40cd4c98, 32'hc00add85} /* (11, 23, 22) {real, imag} */,
  {32'h4126d078, 32'h3fc7d6bc} /* (11, 23, 21) {real, imag} */,
  {32'h40a70fda, 32'h40150068} /* (11, 23, 20) {real, imag} */,
  {32'h3ff86694, 32'h408cb4bc} /* (11, 23, 19) {real, imag} */,
  {32'hc0305b2a, 32'h400e99c7} /* (11, 23, 18) {real, imag} */,
  {32'hc03d2237, 32'hc02298f5} /* (11, 23, 17) {real, imag} */,
  {32'h40207eb9, 32'h3e5d2092} /* (11, 23, 16) {real, imag} */,
  {32'hbea07760, 32'h3e51d6d0} /* (11, 23, 15) {real, imag} */,
  {32'hc0caee3f, 32'hc0952ccb} /* (11, 23, 14) {real, imag} */,
  {32'hc0d9afd0, 32'hc09c3d3f} /* (11, 23, 13) {real, imag} */,
  {32'hbf95b9fe, 32'hc007e3b0} /* (11, 23, 12) {real, imag} */,
  {32'h400d17b2, 32'hc0950c4a} /* (11, 23, 11) {real, imag} */,
  {32'h40e1efe0, 32'h3e94e618} /* (11, 23, 10) {real, imag} */,
  {32'h40aea8a9, 32'h3f82606b} /* (11, 23, 9) {real, imag} */,
  {32'h404b7e0a, 32'hc00b7d95} /* (11, 23, 8) {real, imag} */,
  {32'h4035f0f2, 32'hc0d4ce6e} /* (11, 23, 7) {real, imag} */,
  {32'h400ecc0d, 32'hc044ac88} /* (11, 23, 6) {real, imag} */,
  {32'hc01ad9a4, 32'h3f790678} /* (11, 23, 5) {real, imag} */,
  {32'h408c10ce, 32'h401d42a7} /* (11, 23, 4) {real, imag} */,
  {32'h400a08f2, 32'h3fc35684} /* (11, 23, 3) {real, imag} */,
  {32'hc0d1b0eb, 32'h3fadb872} /* (11, 23, 2) {real, imag} */,
  {32'hc0bd6deb, 32'h4048cc76} /* (11, 23, 1) {real, imag} */,
  {32'hc0035e78, 32'h4009f089} /* (11, 23, 0) {real, imag} */,
  {32'hc00a3514, 32'hbfb0e04c} /* (11, 22, 31) {real, imag} */,
  {32'hc0c24185, 32'hbffac538} /* (11, 22, 30) {real, imag} */,
  {32'h400ee4c4, 32'hc0970820} /* (11, 22, 29) {real, imag} */,
  {32'h4081722d, 32'hc08e0886} /* (11, 22, 28) {real, imag} */,
  {32'h40df6a0b, 32'h3ff4d4a0} /* (11, 22, 27) {real, imag} */,
  {32'h4052969a, 32'hbf07abc4} /* (11, 22, 26) {real, imag} */,
  {32'hbf835e1f, 32'h40526c8a} /* (11, 22, 25) {real, imag} */,
  {32'hc0ba4229, 32'h408347eb} /* (11, 22, 24) {real, imag} */,
  {32'h406ba52a, 32'h4005d928} /* (11, 22, 23) {real, imag} */,
  {32'h4003d653, 32'h3f889a66} /* (11, 22, 22) {real, imag} */,
  {32'h3e92240c, 32'hbf8f8d0b} /* (11, 22, 21) {real, imag} */,
  {32'h408fdc60, 32'h40043b56} /* (11, 22, 20) {real, imag} */,
  {32'h401ea696, 32'hbeae8e80} /* (11, 22, 19) {real, imag} */,
  {32'hbff72afd, 32'h4030ed16} /* (11, 22, 18) {real, imag} */,
  {32'hc092e821, 32'h406ae60d} /* (11, 22, 17) {real, imag} */,
  {32'h3f072b86, 32'h40198b4a} /* (11, 22, 16) {real, imag} */,
  {32'h4019b68e, 32'h3ee39e70} /* (11, 22, 15) {real, imag} */,
  {32'hbfae0d08, 32'hc0702bc6} /* (11, 22, 14) {real, imag} */,
  {32'hc022bda7, 32'h404c1e1c} /* (11, 22, 13) {real, imag} */,
  {32'h408b0fb0, 32'h402930ba} /* (11, 22, 12) {real, imag} */,
  {32'h404f1d54, 32'h40d0e886} /* (11, 22, 11) {real, imag} */,
  {32'hc0b21194, 32'h40801cdd} /* (11, 22, 10) {real, imag} */,
  {32'h3dfa2f20, 32'hbf9b7f58} /* (11, 22, 9) {real, imag} */,
  {32'hbf601140, 32'hc01021ae} /* (11, 22, 8) {real, imag} */,
  {32'hc0a7471c, 32'h3f8cc370} /* (11, 22, 7) {real, imag} */,
  {32'hc0a4c5a4, 32'hbfdc6043} /* (11, 22, 6) {real, imag} */,
  {32'h3ff9696a, 32'hbf690888} /* (11, 22, 5) {real, imag} */,
  {32'h409f833f, 32'h405d8dc0} /* (11, 22, 4) {real, imag} */,
  {32'hc081335d, 32'hc089222b} /* (11, 22, 3) {real, imag} */,
  {32'hbf979ef8, 32'hc076b144} /* (11, 22, 2) {real, imag} */,
  {32'h3fefbf81, 32'hbfab8a3c} /* (11, 22, 1) {real, imag} */,
  {32'h400df880, 32'h3fcf4745} /* (11, 22, 0) {real, imag} */,
  {32'h3cb135c0, 32'h3e88d8e8} /* (11, 21, 31) {real, imag} */,
  {32'h3f041164, 32'h3f9e4645} /* (11, 21, 30) {real, imag} */,
  {32'hbf1c7455, 32'h401a7990} /* (11, 21, 29) {real, imag} */,
  {32'hbfb55d1c, 32'hbeabda10} /* (11, 21, 28) {real, imag} */,
  {32'h3e085360, 32'hbe7a8250} /* (11, 21, 27) {real, imag} */,
  {32'hbfa06914, 32'h40a94fd2} /* (11, 21, 26) {real, imag} */,
  {32'hc0c33120, 32'h40ab2a6a} /* (11, 21, 25) {real, imag} */,
  {32'hc0ecc271, 32'hc00d49f9} /* (11, 21, 24) {real, imag} */,
  {32'hbfd0379a, 32'hc117b28a} /* (11, 21, 23) {real, imag} */,
  {32'h3f14f21e, 32'hc0d7f9e4} /* (11, 21, 22) {real, imag} */,
  {32'hc00b855b, 32'hc019c916} /* (11, 21, 21) {real, imag} */,
  {32'hc0c57f14, 32'hbfd3b351} /* (11, 21, 20) {real, imag} */,
  {32'hbf54ecda, 32'hbfab3d49} /* (11, 21, 19) {real, imag} */,
  {32'h406795da, 32'h3eeaab70} /* (11, 21, 18) {real, imag} */,
  {32'h3fd6d988, 32'hbff0b1f2} /* (11, 21, 17) {real, imag} */,
  {32'hc077b5a0, 32'h3e3fbbb0} /* (11, 21, 16) {real, imag} */,
  {32'hbf8166ba, 32'hc032ab70} /* (11, 21, 15) {real, imag} */,
  {32'h3db9c0b0, 32'hc02c5593} /* (11, 21, 14) {real, imag} */,
  {32'hbf2a8c3c, 32'hc0a4661c} /* (11, 21, 13) {real, imag} */,
  {32'hc00e5592, 32'hc0dc1adc} /* (11, 21, 12) {real, imag} */,
  {32'hc00c7192, 32'hbfce5b43} /* (11, 21, 11) {real, imag} */,
  {32'hbfe8c76a, 32'hbf0387d8} /* (11, 21, 10) {real, imag} */,
  {32'hc04e4845, 32'h4028a6cc} /* (11, 21, 9) {real, imag} */,
  {32'hbf9acd98, 32'h40ae32fe} /* (11, 21, 8) {real, imag} */,
  {32'h3fef62ee, 32'h40b0c1f8} /* (11, 21, 7) {real, imag} */,
  {32'hc00516c5, 32'h408e12b1} /* (11, 21, 6) {real, imag} */,
  {32'h3f72e940, 32'h4092e97f} /* (11, 21, 5) {real, imag} */,
  {32'hbf2c9b16, 32'h40034224} /* (11, 21, 4) {real, imag} */,
  {32'hbfe5016c, 32'h4030f91a} /* (11, 21, 3) {real, imag} */,
  {32'hc07bb16a, 32'h404f5ac3} /* (11, 21, 2) {real, imag} */,
  {32'hc004bfc1, 32'h3f49b74c} /* (11, 21, 1) {real, imag} */,
  {32'hbfcb962e, 32'h3f36dd28} /* (11, 21, 0) {real, imag} */,
  {32'h3f86be60, 32'hbf14b0a0} /* (11, 20, 31) {real, imag} */,
  {32'h4038d8d3, 32'hbfbe1e3b} /* (11, 20, 30) {real, imag} */,
  {32'hc02537f6, 32'h3e853c12} /* (11, 20, 29) {real, imag} */,
  {32'hc02a5c4a, 32'hbe881380} /* (11, 20, 28) {real, imag} */,
  {32'hc0280ca6, 32'hc031a8d8} /* (11, 20, 27) {real, imag} */,
  {32'hc083abde, 32'h3f55ea44} /* (11, 20, 26) {real, imag} */,
  {32'hbf86522b, 32'h3f9830fe} /* (11, 20, 25) {real, imag} */,
  {32'h3ffc65bb, 32'hbf5e77f5} /* (11, 20, 24) {real, imag} */,
  {32'hbe38c530, 32'h402ee588} /* (11, 20, 23) {real, imag} */,
  {32'hc03c3c30, 32'hbfb44c8e} /* (11, 20, 22) {real, imag} */,
  {32'hc004916f, 32'hc0bc55de} /* (11, 20, 21) {real, imag} */,
  {32'hbeba6c3c, 32'hbfcffaf2} /* (11, 20, 20) {real, imag} */,
  {32'hbefc9478, 32'h400eb0dd} /* (11, 20, 19) {real, imag} */,
  {32'hbd60c740, 32'hc030c82c} /* (11, 20, 18) {real, imag} */,
  {32'hc0526db6, 32'h3f62dd18} /* (11, 20, 17) {real, imag} */,
  {32'hc08ccade, 32'h3f6866ac} /* (11, 20, 16) {real, imag} */,
  {32'hbe8b24e0, 32'hbfd5c1af} /* (11, 20, 15) {real, imag} */,
  {32'h3f02cbec, 32'hbf8b3095} /* (11, 20, 14) {real, imag} */,
  {32'h4001f238, 32'h3f5e1ea2} /* (11, 20, 13) {real, imag} */,
  {32'h3fa6a929, 32'h40b04215} /* (11, 20, 12) {real, imag} */,
  {32'h3f2625ee, 32'h401c91fb} /* (11, 20, 11) {real, imag} */,
  {32'h3f53b335, 32'hbf96e283} /* (11, 20, 10) {real, imag} */,
  {32'h3e8cdbf0, 32'hc08fb48b} /* (11, 20, 9) {real, imag} */,
  {32'hc0108e06, 32'hc0513aac} /* (11, 20, 8) {real, imag} */,
  {32'hc0664506, 32'hbf01d388} /* (11, 20, 7) {real, imag} */,
  {32'hbf9a2ef5, 32'hbfc9a89e} /* (11, 20, 6) {real, imag} */,
  {32'h4072fe9d, 32'hc078d72b} /* (11, 20, 5) {real, imag} */,
  {32'hc01a7f0b, 32'hbf5e2b4d} /* (11, 20, 4) {real, imag} */,
  {32'hbf2a83ea, 32'hbf4b9abc} /* (11, 20, 3) {real, imag} */,
  {32'hbf30bef8, 32'hc032cc3d} /* (11, 20, 2) {real, imag} */,
  {32'hbfeba18b, 32'h400e5b09} /* (11, 20, 1) {real, imag} */,
  {32'hc004a40f, 32'h3f9563b4} /* (11, 20, 0) {real, imag} */,
  {32'h4021eab4, 32'hbc54c000} /* (11, 19, 31) {real, imag} */,
  {32'h4034054e, 32'h3eeb9d50} /* (11, 19, 30) {real, imag} */,
  {32'hc003a42e, 32'h3ffd3d84} /* (11, 19, 29) {real, imag} */,
  {32'hc0787a44, 32'hbe829074} /* (11, 19, 28) {real, imag} */,
  {32'hc02144d8, 32'h401884f0} /* (11, 19, 27) {real, imag} */,
  {32'hbda46240, 32'h3fcc9868} /* (11, 19, 26) {real, imag} */,
  {32'h3ff093a5, 32'hbfe6bf68} /* (11, 19, 25) {real, imag} */,
  {32'h3fd32604, 32'hc01ebada} /* (11, 19, 24) {real, imag} */,
  {32'h40597b49, 32'h3f91e854} /* (11, 19, 23) {real, imag} */,
  {32'h403f0c93, 32'h40ad4f63} /* (11, 19, 22) {real, imag} */,
  {32'hbfb3e312, 32'h3fb8168a} /* (11, 19, 21) {real, imag} */,
  {32'hc0422ad6, 32'hbfb5f0fa} /* (11, 19, 20) {real, imag} */,
  {32'hc006890a, 32'h3f91d888} /* (11, 19, 19) {real, imag} */,
  {32'hc0124ac8, 32'h3ffb5a20} /* (11, 19, 18) {real, imag} */,
  {32'h3fae1a4a, 32'hc001e358} /* (11, 19, 17) {real, imag} */,
  {32'h3fb4265e, 32'h3fce7449} /* (11, 19, 16) {real, imag} */,
  {32'hbfa546e9, 32'h3f8f0aec} /* (11, 19, 15) {real, imag} */,
  {32'hbeef4dfc, 32'hc01453ba} /* (11, 19, 14) {real, imag} */,
  {32'h3fc638b0, 32'hbfa5bdba} /* (11, 19, 13) {real, imag} */,
  {32'h3f4cd350, 32'h3ef0f8d6} /* (11, 19, 12) {real, imag} */,
  {32'hbf660c8c, 32'h40006c90} /* (11, 19, 11) {real, imag} */,
  {32'hc0516e46, 32'hbfb4e042} /* (11, 19, 10) {real, imag} */,
  {32'hc088b7a0, 32'hbfbb0aca} /* (11, 19, 9) {real, imag} */,
  {32'hbd3a1b60, 32'hbfe5d6a5} /* (11, 19, 8) {real, imag} */,
  {32'hbe46bee0, 32'hbf90edd0} /* (11, 19, 7) {real, imag} */,
  {32'hbfd5cdd3, 32'hbf6e7df8} /* (11, 19, 6) {real, imag} */,
  {32'h3eb74610, 32'hbf20e556} /* (11, 19, 5) {real, imag} */,
  {32'h3fdb7b22, 32'hc03c01ec} /* (11, 19, 4) {real, imag} */,
  {32'hbf40a490, 32'hc09bfee8} /* (11, 19, 3) {real, imag} */,
  {32'h3f015942, 32'hc0a7a609} /* (11, 19, 2) {real, imag} */,
  {32'h4061111e, 32'hbf4237ae} /* (11, 19, 1) {real, imag} */,
  {32'h40389ef4, 32'hbf00f516} /* (11, 19, 0) {real, imag} */,
  {32'hbfe018a8, 32'h3e140400} /* (11, 18, 31) {real, imag} */,
  {32'h3fb29136, 32'h4008656b} /* (11, 18, 30) {real, imag} */,
  {32'h3fa4830c, 32'h400af107} /* (11, 18, 29) {real, imag} */,
  {32'h3f3cbf12, 32'h3e6e5b74} /* (11, 18, 28) {real, imag} */,
  {32'hc02b2e37, 32'hbf41af48} /* (11, 18, 27) {real, imag} */,
  {32'hbf74a64c, 32'h402cbec4} /* (11, 18, 26) {real, imag} */,
  {32'h3ed47830, 32'h400ea492} /* (11, 18, 25) {real, imag} */,
  {32'hc02a864a, 32'hc0203e55} /* (11, 18, 24) {real, imag} */,
  {32'h3f2d4d6c, 32'hc03c174e} /* (11, 18, 23) {real, imag} */,
  {32'h3fd30969, 32'hbfb3f196} /* (11, 18, 22) {real, imag} */,
  {32'hbe5d3bd0, 32'hbff895d7} /* (11, 18, 21) {real, imag} */,
  {32'hbf8c6ed7, 32'hbfe9c210} /* (11, 18, 20) {real, imag} */,
  {32'hbed716b0, 32'hbf0dcbd3} /* (11, 18, 19) {real, imag} */,
  {32'hbee56c70, 32'hbef8b880} /* (11, 18, 18) {real, imag} */,
  {32'hbf658bb0, 32'h3fd865d6} /* (11, 18, 17) {real, imag} */,
  {32'h3f62f154, 32'h3ea2a1ec} /* (11, 18, 16) {real, imag} */,
  {32'h3f9b0133, 32'h3f0797fc} /* (11, 18, 15) {real, imag} */,
  {32'h4025c68d, 32'h3f8f8639} /* (11, 18, 14) {real, imag} */,
  {32'hbf1d56de, 32'h3f91cb54} /* (11, 18, 13) {real, imag} */,
  {32'hbff98dde, 32'h3fe4555e} /* (11, 18, 12) {real, imag} */,
  {32'hbe928860, 32'hc00384c2} /* (11, 18, 11) {real, imag} */,
  {32'h3e8a8d50, 32'hc062716f} /* (11, 18, 10) {real, imag} */,
  {32'h3df13e00, 32'hbf08d488} /* (11, 18, 9) {real, imag} */,
  {32'h3ff09102, 32'hc01f5286} /* (11, 18, 8) {real, imag} */,
  {32'hbe545080, 32'hbe6b92a8} /* (11, 18, 7) {real, imag} */,
  {32'hbe7c2c40, 32'hbf7cabd6} /* (11, 18, 6) {real, imag} */,
  {32'h400dfe5e, 32'hbf7e0ac5} /* (11, 18, 5) {real, imag} */,
  {32'h405a2c2c, 32'h3f4986cc} /* (11, 18, 4) {real, imag} */,
  {32'h3ff8dcde, 32'h3fa28398} /* (11, 18, 3) {real, imag} */,
  {32'h40132e53, 32'hbf652972} /* (11, 18, 2) {real, imag} */,
  {32'h40261ed6, 32'h3e2a382c} /* (11, 18, 1) {real, imag} */,
  {32'h3ff6b74d, 32'h4018b040} /* (11, 18, 0) {real, imag} */,
  {32'h401a2be6, 32'hbed75a00} /* (11, 17, 31) {real, imag} */,
  {32'h3f083d89, 32'hbef3d0a0} /* (11, 17, 30) {real, imag} */,
  {32'hbe9ae3cc, 32'hbfefcb24} /* (11, 17, 29) {real, imag} */,
  {32'hbffe8dca, 32'hbf91ad98} /* (11, 17, 28) {real, imag} */,
  {32'hc02836f2, 32'h3eff261e} /* (11, 17, 27) {real, imag} */,
  {32'hbf3858e4, 32'hbe487b38} /* (11, 17, 26) {real, imag} */,
  {32'h3f514de8, 32'hbfee6526} /* (11, 17, 25) {real, imag} */,
  {32'hbfbc7c06, 32'hbf985d2c} /* (11, 17, 24) {real, imag} */,
  {32'hbdb57a40, 32'hbeaeafc8} /* (11, 17, 23) {real, imag} */,
  {32'hbfa30b9e, 32'h400c3f59} /* (11, 17, 22) {real, imag} */,
  {32'hbfcdb9cf, 32'h40531378} /* (11, 17, 21) {real, imag} */,
  {32'h3f55310a, 32'h4013c780} /* (11, 17, 20) {real, imag} */,
  {32'h3f2e790a, 32'h3ef1a948} /* (11, 17, 19) {real, imag} */,
  {32'hbfad64d0, 32'hbf40a948} /* (11, 17, 18) {real, imag} */,
  {32'hbf591d80, 32'hbe8101e2} /* (11, 17, 17) {real, imag} */,
  {32'h402ce2a6, 32'h3ed3e27c} /* (11, 17, 16) {real, imag} */,
  {32'h3fadc578, 32'hbfce7331} /* (11, 17, 15) {real, imag} */,
  {32'h403723f0, 32'hbf2329b0} /* (11, 17, 14) {real, imag} */,
  {32'h40072bf6, 32'hbe23076c} /* (11, 17, 13) {real, imag} */,
  {32'hbfc08652, 32'hbf8f7884} /* (11, 17, 12) {real, imag} */,
  {32'hbf627d52, 32'hc02b693a} /* (11, 17, 11) {real, imag} */,
  {32'hbf8b2511, 32'hbfeee45a} /* (11, 17, 10) {real, imag} */,
  {32'hc04217a2, 32'h3efe9010} /* (11, 17, 9) {real, imag} */,
  {32'hc05419b0, 32'hbfa39f31} /* (11, 17, 8) {real, imag} */,
  {32'hc0514db9, 32'hc05ff046} /* (11, 17, 7) {real, imag} */,
  {32'hc02fd27c, 32'hc02a94d1} /* (11, 17, 6) {real, imag} */,
  {32'h3d0e2f80, 32'hbe9b6b90} /* (11, 17, 5) {real, imag} */,
  {32'hbe258f40, 32'h3fff5798} /* (11, 17, 4) {real, imag} */,
  {32'h3fad782b, 32'h3f71d011} /* (11, 17, 3) {real, imag} */,
  {32'h407fec66, 32'h3fc96868} /* (11, 17, 2) {real, imag} */,
  {32'h3ffd35c6, 32'hbf00cde4} /* (11, 17, 1) {real, imag} */,
  {32'hbf45ddc8, 32'hbf84c9b1} /* (11, 17, 0) {real, imag} */,
  {32'hbfc2988e, 32'h3e09c120} /* (11, 16, 31) {real, imag} */,
  {32'h3f121800, 32'h3ea0dce0} /* (11, 16, 30) {real, imag} */,
  {32'h3ffbc850, 32'hc0074ea3} /* (11, 16, 29) {real, imag} */,
  {32'h3f9faa68, 32'hbf9532ac} /* (11, 16, 28) {real, imag} */,
  {32'hbf5a67bc, 32'h3fa4d37a} /* (11, 16, 27) {real, imag} */,
  {32'hbf29fcfd, 32'h3ef60e3c} /* (11, 16, 26) {real, imag} */,
  {32'h3f1fcf98, 32'h3fff1204} /* (11, 16, 25) {real, imag} */,
  {32'h3f16b140, 32'h3fb2945b} /* (11, 16, 24) {real, imag} */,
  {32'hbf564190, 32'h3cd73180} /* (11, 16, 23) {real, imag} */,
  {32'hbf212490, 32'hbfe4c6e0} /* (11, 16, 22) {real, imag} */,
  {32'h3f99176c, 32'hbf078154} /* (11, 16, 21) {real, imag} */,
  {32'h3f8635c8, 32'h3f3479a0} /* (11, 16, 20) {real, imag} */,
  {32'h3e82593c, 32'h3d32cfa0} /* (11, 16, 19) {real, imag} */,
  {32'h3f906090, 32'h3f8b62a0} /* (11, 16, 18) {real, imag} */,
  {32'hbf639d7a, 32'h3f79f590} /* (11, 16, 17) {real, imag} */,
  {32'h3ecb7810, 32'h3ee3cc40} /* (11, 16, 16) {real, imag} */,
  {32'h406b50d2, 32'hbf3397f8} /* (11, 16, 15) {real, imag} */,
  {32'h3fe93a76, 32'hbe8e18c6} /* (11, 16, 14) {real, imag} */,
  {32'h3e9a7e78, 32'h3f83f5b1} /* (11, 16, 13) {real, imag} */,
  {32'h3e722e38, 32'h3f4b2ff8} /* (11, 16, 12) {real, imag} */,
  {32'h3f8d7c1e, 32'h3ea15e40} /* (11, 16, 11) {real, imag} */,
  {32'h40267d4e, 32'h3ea70340} /* (11, 16, 10) {real, imag} */,
  {32'h3fe6126e, 32'hc00b564a} /* (11, 16, 9) {real, imag} */,
  {32'h4005a6de, 32'hc03b7a7b} /* (11, 16, 8) {real, imag} */,
  {32'h3f7af8b8, 32'hbf70e845} /* (11, 16, 7) {real, imag} */,
  {32'hbff531ec, 32'h403a32d4} /* (11, 16, 6) {real, imag} */,
  {32'h3efbb300, 32'h3d85cf00} /* (11, 16, 5) {real, imag} */,
  {32'h40146244, 32'hbfdf09b0} /* (11, 16, 4) {real, imag} */,
  {32'h3ebe2bd8, 32'h3f8958e4} /* (11, 16, 3) {real, imag} */,
  {32'hbf324a18, 32'h40005a96} /* (11, 16, 2) {real, imag} */,
  {32'h3fe69b58, 32'h3fdb0b74} /* (11, 16, 1) {real, imag} */,
  {32'h3fb1d228, 32'hbe2331e0} /* (11, 16, 0) {real, imag} */,
  {32'h3e4858d8, 32'hbe7a51c0} /* (11, 15, 31) {real, imag} */,
  {32'h3f866a1c, 32'hbfd40ad8} /* (11, 15, 30) {real, imag} */,
  {32'h3fb275b9, 32'hbf8fd364} /* (11, 15, 29) {real, imag} */,
  {32'hbf389a6b, 32'hbf5f6301} /* (11, 15, 28) {real, imag} */,
  {32'h40468596, 32'hbf584737} /* (11, 15, 27) {real, imag} */,
  {32'h4068a6f7, 32'hbde557f0} /* (11, 15, 26) {real, imag} */,
  {32'h3f52e9f8, 32'h3f36f1bc} /* (11, 15, 25) {real, imag} */,
  {32'h3f3af31c, 32'h3f17bda8} /* (11, 15, 24) {real, imag} */,
  {32'h3f2d4b28, 32'hbfcd69b2} /* (11, 15, 23) {real, imag} */,
  {32'hbfa1a42a, 32'hbe66d110} /* (11, 15, 22) {real, imag} */,
  {32'hbc6d8480, 32'h4045a580} /* (11, 15, 21) {real, imag} */,
  {32'h3f0da72a, 32'h40681c84} /* (11, 15, 20) {real, imag} */,
  {32'h3ed46f0c, 32'h3fb5b5ba} /* (11, 15, 19) {real, imag} */,
  {32'h3f7946e0, 32'hbfec0be4} /* (11, 15, 18) {real, imag} */,
  {32'hbf8b5ee8, 32'hbfb6f44c} /* (11, 15, 17) {real, imag} */,
  {32'hbfee07d4, 32'hbf3c7d76} /* (11, 15, 16) {real, imag} */,
  {32'hbf35b380, 32'hbfe7b2cd} /* (11, 15, 15) {real, imag} */,
  {32'hbf0b41c0, 32'hbe77ca00} /* (11, 15, 14) {real, imag} */,
  {32'hbf428618, 32'h3f37a201} /* (11, 15, 13) {real, imag} */,
  {32'hbff41e8e, 32'h40027bb2} /* (11, 15, 12) {real, imag} */,
  {32'hc00d30fc, 32'h3d171aa0} /* (11, 15, 11) {real, imag} */,
  {32'hbe401cf8, 32'hbfc47962} /* (11, 15, 10) {real, imag} */,
  {32'h40131bb4, 32'hbebfccd0} /* (11, 15, 9) {real, imag} */,
  {32'hbf9f3c80, 32'hbf1cd6a2} /* (11, 15, 8) {real, imag} */,
  {32'h3a353000, 32'hbf87e1dc} /* (11, 15, 7) {real, imag} */,
  {32'h3fcfbc38, 32'hbf539a24} /* (11, 15, 6) {real, imag} */,
  {32'hbdd02bc0, 32'hbf6404a8} /* (11, 15, 5) {real, imag} */,
  {32'h3f3b36b0, 32'h3f5e7280} /* (11, 15, 4) {real, imag} */,
  {32'h3f55869a, 32'hbf631d5d} /* (11, 15, 3) {real, imag} */,
  {32'h3f0a2d28, 32'h3e9df1e8} /* (11, 15, 2) {real, imag} */,
  {32'h3f829516, 32'h40397d0d} /* (11, 15, 1) {real, imag} */,
  {32'h3e0dff80, 32'h3f94f5bb} /* (11, 15, 0) {real, imag} */,
  {32'hbf420fd8, 32'hbf3df468} /* (11, 14, 31) {real, imag} */,
  {32'h3f9b53ee, 32'hbeefbf28} /* (11, 14, 30) {real, imag} */,
  {32'hbf4b9998, 32'hbf03c8dc} /* (11, 14, 29) {real, imag} */,
  {32'hbf179372, 32'hbfd8534e} /* (11, 14, 28) {real, imag} */,
  {32'h3e983cf8, 32'h3eec8570} /* (11, 14, 27) {real, imag} */,
  {32'h3df5dd60, 32'h3f7ea0d2} /* (11, 14, 26) {real, imag} */,
  {32'h3fc482ac, 32'h3f15e786} /* (11, 14, 25) {real, imag} */,
  {32'h40038bf2, 32'hbfd56366} /* (11, 14, 24) {real, imag} */,
  {32'h3f94d912, 32'hbf631838} /* (11, 14, 23) {real, imag} */,
  {32'h3fb69b03, 32'hc0114c4f} /* (11, 14, 22) {real, imag} */,
  {32'h3fa3916e, 32'hbf1aa7fe} /* (11, 14, 21) {real, imag} */,
  {32'h3fb11907, 32'hbe78c880} /* (11, 14, 20) {real, imag} */,
  {32'h40095cde, 32'hbe0dc23c} /* (11, 14, 19) {real, imag} */,
  {32'h403381b6, 32'h40060bce} /* (11, 14, 18) {real, imag} */,
  {32'h3f96d478, 32'h4054077d} /* (11, 14, 17) {real, imag} */,
  {32'hbf95212a, 32'hbf850d8b} /* (11, 14, 16) {real, imag} */,
  {32'hbfa20323, 32'hbfc3da94} /* (11, 14, 15) {real, imag} */,
  {32'h3e1ccdd0, 32'hbeb75334} /* (11, 14, 14) {real, imag} */,
  {32'hc0445798, 32'hbe326cec} /* (11, 14, 13) {real, imag} */,
  {32'h3f555e14, 32'hc06ffb37} /* (11, 14, 12) {real, imag} */,
  {32'h3fa48c80, 32'hc04d4476} /* (11, 14, 11) {real, imag} */,
  {32'hbfac7f3c, 32'hc03f6b0f} /* (11, 14, 10) {real, imag} */,
  {32'hc03ea9cc, 32'hc0052ce2} /* (11, 14, 9) {real, imag} */,
  {32'hbfbe3a6e, 32'hc00b710e} /* (11, 14, 8) {real, imag} */,
  {32'hbf8c1e20, 32'h3ea00e14} /* (11, 14, 7) {real, imag} */,
  {32'hc02a8598, 32'h3fb3406b} /* (11, 14, 6) {real, imag} */,
  {32'hbf3aad92, 32'hbf1004ab} /* (11, 14, 5) {real, imag} */,
  {32'hbfe9c1b0, 32'hbec66510} /* (11, 14, 4) {real, imag} */,
  {32'hbfeb64da, 32'h3e13b674} /* (11, 14, 3) {real, imag} */,
  {32'h3f33d824, 32'h3de18830} /* (11, 14, 2) {real, imag} */,
  {32'hbfc80323, 32'hbdcacd58} /* (11, 14, 1) {real, imag} */,
  {32'hbfaf74df, 32'hbf28d6ca} /* (11, 14, 0) {real, imag} */,
  {32'hbfa31a27, 32'h4045b8f0} /* (11, 13, 31) {real, imag} */,
  {32'hc011f946, 32'h400a4f1e} /* (11, 13, 30) {real, imag} */,
  {32'hbdf68fc8, 32'hbd769c80} /* (11, 13, 29) {real, imag} */,
  {32'h4011c4c0, 32'h4002ad6e} /* (11, 13, 28) {real, imag} */,
  {32'h401a6ee0, 32'h3ff2e8ff} /* (11, 13, 27) {real, imag} */,
  {32'h40052906, 32'hbf1c15d0} /* (11, 13, 26) {real, imag} */,
  {32'h3f83aebf, 32'hbf3a9c54} /* (11, 13, 25) {real, imag} */,
  {32'hbe846bb0, 32'hbf91db97} /* (11, 13, 24) {real, imag} */,
  {32'h3f40e90c, 32'hbfe67db4} /* (11, 13, 23) {real, imag} */,
  {32'h408e6742, 32'h3cde2600} /* (11, 13, 22) {real, imag} */,
  {32'h40490543, 32'h402ddd2b} /* (11, 13, 21) {real, imag} */,
  {32'hbf88f774, 32'h3e7e9234} /* (11, 13, 20) {real, imag} */,
  {32'h3e2a4738, 32'h3f0f3d10} /* (11, 13, 19) {real, imag} */,
  {32'hbeab5f9c, 32'h403bd55e} /* (11, 13, 18) {real, imag} */,
  {32'hbf1b2e6c, 32'h4041e27c} /* (11, 13, 17) {real, imag} */,
  {32'h402ba615, 32'h40363ea6} /* (11, 13, 16) {real, imag} */,
  {32'h402af9f6, 32'hbe662820} /* (11, 13, 15) {real, imag} */,
  {32'h3fc443e9, 32'h3f107098} /* (11, 13, 14) {real, imag} */,
  {32'hbeae4940, 32'h3f765f9c} /* (11, 13, 13) {real, imag} */,
  {32'h3f07e0f0, 32'hbed3cffa} /* (11, 13, 12) {real, imag} */,
  {32'hbfdbc50e, 32'h3e08f27c} /* (11, 13, 11) {real, imag} */,
  {32'hc0199766, 32'h3e909c48} /* (11, 13, 10) {real, imag} */,
  {32'h3f7f6540, 32'h3f9ee5b6} /* (11, 13, 9) {real, imag} */,
  {32'h3f32d21a, 32'hbe809a54} /* (11, 13, 8) {real, imag} */,
  {32'hbeea4ef0, 32'hbf50ec80} /* (11, 13, 7) {real, imag} */,
  {32'hbe1d8b88, 32'hc02de35e} /* (11, 13, 6) {real, imag} */,
  {32'h3f95cfd0, 32'hc054339c} /* (11, 13, 5) {real, imag} */,
  {32'h3f1f4264, 32'hc024194c} /* (11, 13, 4) {real, imag} */,
  {32'h3fe02e60, 32'hbedf1698} /* (11, 13, 3) {real, imag} */,
  {32'hbfc9b843, 32'h3f81631c} /* (11, 13, 2) {real, imag} */,
  {32'h40094126, 32'h3f918cc0} /* (11, 13, 1) {real, imag} */,
  {32'h402a7344, 32'h3f7bc868} /* (11, 13, 0) {real, imag} */,
  {32'hc03c78f0, 32'h3fb0ad86} /* (11, 12, 31) {real, imag} */,
  {32'hc03ef6b1, 32'h3f2b5922} /* (11, 12, 30) {real, imag} */,
  {32'h3e51d3a8, 32'h3fa71794} /* (11, 12, 29) {real, imag} */,
  {32'h3fd7c58c, 32'h4029e554} /* (11, 12, 28) {real, imag} */,
  {32'hbee71be0, 32'hbbc0d900} /* (11, 12, 27) {real, imag} */,
  {32'hbfb80ba6, 32'hc0828e82} /* (11, 12, 26) {real, imag} */,
  {32'h402f64c2, 32'hc00bfd51} /* (11, 12, 25) {real, imag} */,
  {32'h3ed1ff64, 32'h3eff2c6a} /* (11, 12, 24) {real, imag} */,
  {32'h3f60cf7c, 32'h405b0fe8} /* (11, 12, 23) {real, imag} */,
  {32'hbfb9583b, 32'h3fff9ade} /* (11, 12, 22) {real, imag} */,
  {32'hc01d84e1, 32'hbfe8a1c2} /* (11, 12, 21) {real, imag} */,
  {32'hc0257ac6, 32'h3fa8cce6} /* (11, 12, 20) {real, imag} */,
  {32'hc0999812, 32'hbf17abf4} /* (11, 12, 19) {real, imag} */,
  {32'h3f717ef4, 32'h3f2d0ede} /* (11, 12, 18) {real, imag} */,
  {32'hbf92cb85, 32'h3f665ae8} /* (11, 12, 17) {real, imag} */,
  {32'hbf39ebea, 32'h40043dd3} /* (11, 12, 16) {real, imag} */,
  {32'hbf93142e, 32'h3f3b07f2} /* (11, 12, 15) {real, imag} */,
  {32'h3ce35200, 32'hc022c768} /* (11, 12, 14) {real, imag} */,
  {32'h4055a8bc, 32'hc0967862} /* (11, 12, 13) {real, imag} */,
  {32'h3ea63b64, 32'hc03e7e56} /* (11, 12, 12) {real, imag} */,
  {32'h3fd49c9d, 32'h3f564c04} /* (11, 12, 11) {real, imag} */,
  {32'h40323885, 32'hbdf81230} /* (11, 12, 10) {real, imag} */,
  {32'h40960d3f, 32'hc097e3fb} /* (11, 12, 9) {real, imag} */,
  {32'h409a94f3, 32'hc073987a} /* (11, 12, 8) {real, imag} */,
  {32'h4036c74a, 32'hc0307e30} /* (11, 12, 7) {real, imag} */,
  {32'h408250db, 32'hc00a8e58} /* (11, 12, 6) {real, imag} */,
  {32'h40077c97, 32'hbeccbe58} /* (11, 12, 5) {real, imag} */,
  {32'hc04b8c8b, 32'hbf23d15d} /* (11, 12, 4) {real, imag} */,
  {32'hc04a7098, 32'hc0798583} /* (11, 12, 3) {real, imag} */,
  {32'h3f1c74c0, 32'hc00d86ff} /* (11, 12, 2) {real, imag} */,
  {32'hbdfdc050, 32'h403567e7} /* (11, 12, 1) {real, imag} */,
  {32'hc029e119, 32'hbfb19150} /* (11, 12, 0) {real, imag} */,
  {32'hc048ab84, 32'h4031718b} /* (11, 11, 31) {real, imag} */,
  {32'hc0a584e6, 32'h40743bca} /* (11, 11, 30) {real, imag} */,
  {32'hbf467f7b, 32'hbf7f6558} /* (11, 11, 29) {real, imag} */,
  {32'hbf9b0108, 32'hc02fda22} /* (11, 11, 28) {real, imag} */,
  {32'hc04e27e6, 32'hc101be67} /* (11, 11, 27) {real, imag} */,
  {32'h3ee1c130, 32'hc0e66c4e} /* (11, 11, 26) {real, imag} */,
  {32'hc069a6e4, 32'hc0a2e85a} /* (11, 11, 25) {real, imag} */,
  {32'hbfea1284, 32'hbfa8aec2} /* (11, 11, 24) {real, imag} */,
  {32'h3fbb85ba, 32'hbff43eda} /* (11, 11, 23) {real, imag} */,
  {32'h3f3c544a, 32'hc07e5f7c} /* (11, 11, 22) {real, imag} */,
  {32'h3f49f114, 32'hc04f88d0} /* (11, 11, 21) {real, imag} */,
  {32'h40517bf7, 32'hbfdc385d} /* (11, 11, 20) {real, imag} */,
  {32'h3fc80643, 32'hbf5204b2} /* (11, 11, 19) {real, imag} */,
  {32'hc0037930, 32'hc03c96ea} /* (11, 11, 18) {real, imag} */,
  {32'h3ea70440, 32'h3ece270a} /* (11, 11, 17) {real, imag} */,
  {32'h405ef854, 32'hbf850a7a} /* (11, 11, 16) {real, imag} */,
  {32'h40192f63, 32'h409a43a3} /* (11, 11, 15) {real, imag} */,
  {32'hbf960e55, 32'h402e6bdd} /* (11, 11, 14) {real, imag} */,
  {32'h3f92bed6, 32'hbfdff69e} /* (11, 11, 13) {real, imag} */,
  {32'h3f05008e, 32'hc01c851c} /* (11, 11, 12) {real, imag} */,
  {32'hbe1c1960, 32'hbfe7f583} /* (11, 11, 11) {real, imag} */,
  {32'hc04d46b9, 32'hc0030cea} /* (11, 11, 10) {real, imag} */,
  {32'hc07eb909, 32'h3fbac5e7} /* (11, 11, 9) {real, imag} */,
  {32'h3f671ec0, 32'h3fe1ad7e} /* (11, 11, 8) {real, imag} */,
  {32'h402c494b, 32'hbebe1760} /* (11, 11, 7) {real, imag} */,
  {32'h408373fe, 32'h3f449470} /* (11, 11, 6) {real, imag} */,
  {32'h40bb4084, 32'hc00ce22e} /* (11, 11, 5) {real, imag} */,
  {32'h406eaf22, 32'hbfd92151} /* (11, 11, 4) {real, imag} */,
  {32'h3f92b894, 32'h3fcb4a15} /* (11, 11, 3) {real, imag} */,
  {32'hc072b382, 32'h3fcad03a} /* (11, 11, 2) {real, imag} */,
  {32'hc10e6b3b, 32'h3f44beb4} /* (11, 11, 1) {real, imag} */,
  {32'hc105390b, 32'hbfe52ed0} /* (11, 11, 0) {real, imag} */,
  {32'hc082bda4, 32'h409537ed} /* (11, 10, 31) {real, imag} */,
  {32'hbffbf9ec, 32'h41248f5d} /* (11, 10, 30) {real, imag} */,
  {32'hbeb98ae4, 32'h40c088e0} /* (11, 10, 29) {real, imag} */,
  {32'h3f1aa37a, 32'h3fdf856c} /* (11, 10, 28) {real, imag} */,
  {32'hbe0465e0, 32'h40604e90} /* (11, 10, 27) {real, imag} */,
  {32'hbf39c4e0, 32'h40471b7f} /* (11, 10, 26) {real, imag} */,
  {32'hbfa3c1e5, 32'h3e91dff8} /* (11, 10, 25) {real, imag} */,
  {32'h3fd00f98, 32'h406ca932} /* (11, 10, 24) {real, imag} */,
  {32'h4049f1f6, 32'h4139ceef} /* (11, 10, 23) {real, imag} */,
  {32'hc007d549, 32'h40c30550} /* (11, 10, 22) {real, imag} */,
  {32'h3eb6db74, 32'hc05038e0} /* (11, 10, 21) {real, imag} */,
  {32'h40dc1c40, 32'hc0a1a513} /* (11, 10, 20) {real, imag} */,
  {32'h4114c562, 32'h40ecce2a} /* (11, 10, 19) {real, imag} */,
  {32'hbf3e7b2e, 32'h4072f3c4} /* (11, 10, 18) {real, imag} */,
  {32'hc0ab6d1d, 32'h3ff83aea} /* (11, 10, 17) {real, imag} */,
  {32'h403f0e5a, 32'hbf00eae8} /* (11, 10, 16) {real, imag} */,
  {32'h4039674a, 32'hc0107e47} /* (11, 10, 15) {real, imag} */,
  {32'hc0b102fa, 32'h4084b828} /* (11, 10, 14) {real, imag} */,
  {32'hc082d210, 32'hc043a880} /* (11, 10, 13) {real, imag} */,
  {32'h40673a99, 32'hc074faa6} /* (11, 10, 12) {real, imag} */,
  {32'h3fc8c8c0, 32'h3e491630} /* (11, 10, 11) {real, imag} */,
  {32'hc0207dcc, 32'h404f9c82} /* (11, 10, 10) {real, imag} */,
  {32'h4083f1e0, 32'h4094da6a} /* (11, 10, 9) {real, imag} */,
  {32'h40672b36, 32'h3f1f05ee} /* (11, 10, 8) {real, imag} */,
  {32'hc0624218, 32'h40525d4a} /* (11, 10, 7) {real, imag} */,
  {32'hc005da9d, 32'h405772ce} /* (11, 10, 6) {real, imag} */,
  {32'h3e43b59c, 32'h3cfc73f0} /* (11, 10, 5) {real, imag} */,
  {32'hc04e758a, 32'hbfbf7721} /* (11, 10, 4) {real, imag} */,
  {32'hc0eeb519, 32'h3f325b18} /* (11, 10, 3) {real, imag} */,
  {32'hc0ad7048, 32'hbe0a9f38} /* (11, 10, 2) {real, imag} */,
  {32'hbfc78f0b, 32'h3facec62} /* (11, 10, 1) {real, imag} */,
  {32'hbffda44c, 32'h4002b9e0} /* (11, 10, 0) {real, imag} */,
  {32'h4004cfa0, 32'hc0b93070} /* (11, 9, 31) {real, imag} */,
  {32'hbe47fc00, 32'hc1283259} /* (11, 9, 30) {real, imag} */,
  {32'h3f70ed79, 32'hc0b2e466} /* (11, 9, 29) {real, imag} */,
  {32'h3f9ab666, 32'hc045b6f7} /* (11, 9, 28) {real, imag} */,
  {32'h4086a7cf, 32'h3fc825dc} /* (11, 9, 27) {real, imag} */,
  {32'h3facf8f4, 32'hc01bb164} /* (11, 9, 26) {real, imag} */,
  {32'hbd335420, 32'hbf4d1b40} /* (11, 9, 25) {real, imag} */,
  {32'h3f1088d2, 32'hc0b9e81c} /* (11, 9, 24) {real, imag} */,
  {32'hbd791980, 32'hc107e7f2} /* (11, 9, 23) {real, imag} */,
  {32'h3fcda168, 32'hc0cdc2a2} /* (11, 9, 22) {real, imag} */,
  {32'h4096900c, 32'hc0d91e4f} /* (11, 9, 21) {real, imag} */,
  {32'h40a26cc8, 32'hc0d18ce8} /* (11, 9, 20) {real, imag} */,
  {32'h40379042, 32'hc113c879} /* (11, 9, 19) {real, imag} */,
  {32'h3e006f20, 32'hc091dcf2} /* (11, 9, 18) {real, imag} */,
  {32'hc03b56eb, 32'h3fde6112} /* (11, 9, 17) {real, imag} */,
  {32'hbe378000, 32'hbf10cf88} /* (11, 9, 16) {real, imag} */,
  {32'h408db236, 32'hc018b486} /* (11, 9, 15) {real, imag} */,
  {32'h404f0f42, 32'h40870a3d} /* (11, 9, 14) {real, imag} */,
  {32'hbed66d90, 32'h402faa3a} /* (11, 9, 13) {real, imag} */,
  {32'hbf4c461c, 32'h3ed700ee} /* (11, 9, 12) {real, imag} */,
  {32'hc0b13cb9, 32'h3d93ac80} /* (11, 9, 11) {real, imag} */,
  {32'hc02f5d43, 32'h3e9669a8} /* (11, 9, 10) {real, imag} */,
  {32'hc01b7bc4, 32'h408b61ce} /* (11, 9, 9) {real, imag} */,
  {32'h3f44857a, 32'h40d13924} /* (11, 9, 8) {real, imag} */,
  {32'hc0a71d97, 32'h3c6a0500} /* (11, 9, 7) {real, imag} */,
  {32'h3fd14dde, 32'hc06a7710} /* (11, 9, 6) {real, imag} */,
  {32'h413341ef, 32'h406c2564} /* (11, 9, 5) {real, imag} */,
  {32'h40d4c2ca, 32'h3eef0b40} /* (11, 9, 4) {real, imag} */,
  {32'h404ac86a, 32'hbfb58c3e} /* (11, 9, 3) {real, imag} */,
  {32'h411c7b06, 32'hbf3eed94} /* (11, 9, 2) {real, imag} */,
  {32'h40aac371, 32'h407298ee} /* (11, 9, 1) {real, imag} */,
  {32'hbf6f2d7c, 32'h3f3ff055} /* (11, 9, 0) {real, imag} */,
  {32'h3f7b054c, 32'h3f51f948} /* (11, 8, 31) {real, imag} */,
  {32'h40868b5c, 32'hbf4ce984} /* (11, 8, 30) {real, imag} */,
  {32'h40c11c28, 32'h40463344} /* (11, 8, 29) {real, imag} */,
  {32'hc0f5d494, 32'hbf811e98} /* (11, 8, 28) {real, imag} */,
  {32'hc052cfc3, 32'hc10e25b6} /* (11, 8, 27) {real, imag} */,
  {32'h3fb059fc, 32'hc0cc498e} /* (11, 8, 26) {real, imag} */,
  {32'h3ea76524, 32'h41019eed} /* (11, 8, 25) {real, imag} */,
  {32'h40b6d68a, 32'h401a5b08} /* (11, 8, 24) {real, imag} */,
  {32'h41009cab, 32'hc04b9287} /* (11, 8, 23) {real, imag} */,
  {32'h3feb54e4, 32'h406964ae} /* (11, 8, 22) {real, imag} */,
  {32'hbf1e48e2, 32'h3ffa1d46} /* (11, 8, 21) {real, imag} */,
  {32'h4025c63a, 32'h409f96d8} /* (11, 8, 20) {real, imag} */,
  {32'hbefad51a, 32'h3e5c35a0} /* (11, 8, 19) {real, imag} */,
  {32'hbfbbe5a6, 32'hc038946a} /* (11, 8, 18) {real, imag} */,
  {32'hc020fbe8, 32'hc0164be6} /* (11, 8, 17) {real, imag} */,
  {32'hbda06870, 32'h3f92ed3e} /* (11, 8, 16) {real, imag} */,
  {32'hbe9d8990, 32'h410c770c} /* (11, 8, 15) {real, imag} */,
  {32'hbf367c00, 32'h40cffcbd} /* (11, 8, 14) {real, imag} */,
  {32'hbec88bc0, 32'h4052a03c} /* (11, 8, 13) {real, imag} */,
  {32'h4096905c, 32'hbf44139a} /* (11, 8, 12) {real, imag} */,
  {32'hbf9a140c, 32'h3fcdb066} /* (11, 8, 11) {real, imag} */,
  {32'hbfb30daf, 32'h4095f60a} /* (11, 8, 10) {real, imag} */,
  {32'h3e8d0ca8, 32'hbf4a639c} /* (11, 8, 9) {real, imag} */,
  {32'h3f7d27b8, 32'hc0a8b308} /* (11, 8, 8) {real, imag} */,
  {32'h404b704c, 32'hc0b0ccac} /* (11, 8, 7) {real, imag} */,
  {32'h3f2bd5b8, 32'h40a039e8} /* (11, 8, 6) {real, imag} */,
  {32'h3fefa292, 32'h4105dabc} /* (11, 8, 5) {real, imag} */,
  {32'h40dd0458, 32'hc064a6b4} /* (11, 8, 4) {real, imag} */,
  {32'h3f420528, 32'hc0870148} /* (11, 8, 3) {real, imag} */,
  {32'hc083c5c8, 32'h3fb69c54} /* (11, 8, 2) {real, imag} */,
  {32'hc0e9a86c, 32'hbfd84938} /* (11, 8, 1) {real, imag} */,
  {32'hc027a1dc, 32'h3e6ee100} /* (11, 8, 0) {real, imag} */,
  {32'h3b842c00, 32'hc1099545} /* (11, 7, 31) {real, imag} */,
  {32'hc033f116, 32'hc034a90b} /* (11, 7, 30) {real, imag} */,
  {32'hc09714aa, 32'h40efbe10} /* (11, 7, 29) {real, imag} */,
  {32'hbe872724, 32'h4063f82a} /* (11, 7, 28) {real, imag} */,
  {32'h40a9e645, 32'h3d0e2da0} /* (11, 7, 27) {real, imag} */,
  {32'h3d2c4400, 32'hc048ecfa} /* (11, 7, 26) {real, imag} */,
  {32'hc039ea14, 32'hc114714d} /* (11, 7, 25) {real, imag} */,
  {32'hbec5bfa0, 32'hbf9506c4} /* (11, 7, 24) {real, imag} */,
  {32'h4104d706, 32'h4092152a} /* (11, 7, 23) {real, imag} */,
  {32'h3fa62e70, 32'h402fb859} /* (11, 7, 22) {real, imag} */,
  {32'h3ece5994, 32'h40169f28} /* (11, 7, 21) {real, imag} */,
  {32'hc0eefae3, 32'hc0061156} /* (11, 7, 20) {real, imag} */,
  {32'hc19c9570, 32'h40e5359f} /* (11, 7, 19) {real, imag} */,
  {32'hc1b6be44, 32'h41122762} /* (11, 7, 18) {real, imag} */,
  {32'hc131cba4, 32'h40861d9a} /* (11, 7, 17) {real, imag} */,
  {32'hbee36f34, 32'h402d256a} /* (11, 7, 16) {real, imag} */,
  {32'hc096ed18, 32'h404c3a08} /* (11, 7, 15) {real, imag} */,
  {32'hc04f4cca, 32'hc0f4b0ae} /* (11, 7, 14) {real, imag} */,
  {32'hbfaa93a8, 32'hbfc00c60} /* (11, 7, 13) {real, imag} */,
  {32'hc110c9d6, 32'h400cbf44} /* (11, 7, 12) {real, imag} */,
  {32'hc06b59ea, 32'hc0240029} /* (11, 7, 11) {real, imag} */,
  {32'hc0b6fe5c, 32'h4082d0ec} /* (11, 7, 10) {real, imag} */,
  {32'hc053cf12, 32'h4092fe76} /* (11, 7, 9) {real, imag} */,
  {32'h40784234, 32'h40841762} /* (11, 7, 8) {real, imag} */,
  {32'hc0c42fdb, 32'h4027647b} /* (11, 7, 7) {real, imag} */,
  {32'hc0ef4b55, 32'h3f945714} /* (11, 7, 6) {real, imag} */,
  {32'hbf5699dc, 32'hbfb8057c} /* (11, 7, 5) {real, imag} */,
  {32'h40b36cd1, 32'hbf272918} /* (11, 7, 4) {real, imag} */,
  {32'h412786b8, 32'hbf540940} /* (11, 7, 3) {real, imag} */,
  {32'h4004d376, 32'h400446b8} /* (11, 7, 2) {real, imag} */,
  {32'h40b713bc, 32'h4042b8c1} /* (11, 7, 1) {real, imag} */,
  {32'h4080c3ce, 32'hbf21c325} /* (11, 7, 0) {real, imag} */,
  {32'h40aedc5d, 32'hc0a2ed7a} /* (11, 6, 31) {real, imag} */,
  {32'h40a5454e, 32'hc0897194} /* (11, 6, 30) {real, imag} */,
  {32'h404e8272, 32'h40b67911} /* (11, 6, 29) {real, imag} */,
  {32'h3ea1f6e0, 32'h3fe1c682} /* (11, 6, 28) {real, imag} */,
  {32'hc0e266ba, 32'h40c7237e} /* (11, 6, 27) {real, imag} */,
  {32'h3f175670, 32'h40f98442} /* (11, 6, 26) {real, imag} */,
  {32'h40d53720, 32'h3fd4153c} /* (11, 6, 25) {real, imag} */,
  {32'hc01ba057, 32'hc00cd348} /* (11, 6, 24) {real, imag} */,
  {32'hc154e862, 32'hc07185e0} /* (11, 6, 23) {real, imag} */,
  {32'hc0beb58a, 32'hbe8f11d0} /* (11, 6, 22) {real, imag} */,
  {32'hc0432510, 32'h409d6ccf} /* (11, 6, 21) {real, imag} */,
  {32'hc159b3b5, 32'h3f825b06} /* (11, 6, 20) {real, imag} */,
  {32'hc0e227d3, 32'hc0b9028e} /* (11, 6, 19) {real, imag} */,
  {32'hc048dde7, 32'hbff716e0} /* (11, 6, 18) {real, imag} */,
  {32'hc102b891, 32'hc0cf3d6e} /* (11, 6, 17) {real, imag} */,
  {32'hc10d50ee, 32'h4095d32e} /* (11, 6, 16) {real, imag} */,
  {32'hc0d5c6c2, 32'h3f89f16f} /* (11, 6, 15) {real, imag} */,
  {32'hc0215962, 32'h3f0ead0e} /* (11, 6, 14) {real, imag} */,
  {32'hc133e037, 32'h3f55cc5e} /* (11, 6, 13) {real, imag} */,
  {32'hc16ef6d8, 32'hbda79180} /* (11, 6, 12) {real, imag} */,
  {32'hc12e2539, 32'hc08d6904} /* (11, 6, 11) {real, imag} */,
  {32'hc0034f22, 32'hc12af361} /* (11, 6, 10) {real, imag} */,
  {32'h40c9cab2, 32'hc11a8159} /* (11, 6, 9) {real, imag} */,
  {32'h4047fda9, 32'hc0a9980e} /* (11, 6, 8) {real, imag} */,
  {32'h3e246f34, 32'hc0efe64c} /* (11, 6, 7) {real, imag} */,
  {32'h40674afb, 32'hc095d137} /* (11, 6, 6) {real, imag} */,
  {32'hc0a5a7e4, 32'hc0547337} /* (11, 6, 5) {real, imag} */,
  {32'hc0b91275, 32'h4011860f} /* (11, 6, 4) {real, imag} */,
  {32'h4062b6e9, 32'h40f40bed} /* (11, 6, 3) {real, imag} */,
  {32'h410c707a, 32'h409a8553} /* (11, 6, 2) {real, imag} */,
  {32'hc0383c4e, 32'h4044c7d4} /* (11, 6, 1) {real, imag} */,
  {32'h3e9a4ad6, 32'h40ba73aa} /* (11, 6, 0) {real, imag} */,
  {32'hc0e11af3, 32'hbf820604} /* (11, 5, 31) {real, imag} */,
  {32'hc129bf86, 32'h4092bf29} /* (11, 5, 30) {real, imag} */,
  {32'hc13636c0, 32'h411c3b20} /* (11, 5, 29) {real, imag} */,
  {32'hc12a0c0b, 32'h40373075} /* (11, 5, 28) {real, imag} */,
  {32'hc1b996a5, 32'h40d3b202} /* (11, 5, 27) {real, imag} */,
  {32'hc157ef38, 32'h40f56d28} /* (11, 5, 26) {real, imag} */,
  {32'hc0946543, 32'hbffd63dc} /* (11, 5, 25) {real, imag} */,
  {32'hbe2c0580, 32'hbea695e0} /* (11, 5, 24) {real, imag} */,
  {32'hc098f7bc, 32'h3e01bee0} /* (11, 5, 23) {real, imag} */,
  {32'hc1168e79, 32'h3f2857a0} /* (11, 5, 22) {real, imag} */,
  {32'hc0bfe624, 32'h3fb39e42} /* (11, 5, 21) {real, imag} */,
  {32'h40bfd066, 32'h4118a626} /* (11, 5, 20) {real, imag} */,
  {32'h40920f89, 32'h409f60b5} /* (11, 5, 19) {real, imag} */,
  {32'h40c72b2e, 32'h3f11bccd} /* (11, 5, 18) {real, imag} */,
  {32'h4105de16, 32'h3e0e5834} /* (11, 5, 17) {real, imag} */,
  {32'h40b509af, 32'hbf2515f0} /* (11, 5, 16) {real, imag} */,
  {32'h410e4ee7, 32'hc02de8d3} /* (11, 5, 15) {real, imag} */,
  {32'h40c0cd95, 32'hc08d8756} /* (11, 5, 14) {real, imag} */,
  {32'h4031be2d, 32'h40d3b0ce} /* (11, 5, 13) {real, imag} */,
  {32'h41197f44, 32'h408465a0} /* (11, 5, 12) {real, imag} */,
  {32'h413f7b0b, 32'hc0f8bca0} /* (11, 5, 11) {real, imag} */,
  {32'hc0b35f6e, 32'hc0d241d7} /* (11, 5, 10) {real, imag} */,
  {32'hc0f36eba, 32'hc0cda7ae} /* (11, 5, 9) {real, imag} */,
  {32'hbdd98380, 32'hc0f3c1ac} /* (11, 5, 8) {real, imag} */,
  {32'hc046487f, 32'hc04cca78} /* (11, 5, 7) {real, imag} */,
  {32'h408d446e, 32'hc006d7c4} /* (11, 5, 6) {real, imag} */,
  {32'h3dea7320, 32'h41111e88} /* (11, 5, 5) {real, imag} */,
  {32'hbfd96c65, 32'h40812234} /* (11, 5, 4) {real, imag} */,
  {32'hc05d359c, 32'hbf3455e8} /* (11, 5, 3) {real, imag} */,
  {32'hbf83454d, 32'hbf3d3345} /* (11, 5, 2) {real, imag} */,
  {32'hc019106d, 32'hc0515105} /* (11, 5, 1) {real, imag} */,
  {32'hc0ad6a28, 32'hbf45e874} /* (11, 5, 0) {real, imag} */,
  {32'hbf407530, 32'hc0871721} /* (11, 4, 31) {real, imag} */,
  {32'h40c93162, 32'hc1019bcc} /* (11, 4, 30) {real, imag} */,
  {32'h40fdfefd, 32'hc096dfe5} /* (11, 4, 29) {real, imag} */,
  {32'h3f9de1d3, 32'hc10c7090} /* (11, 4, 28) {real, imag} */,
  {32'hc0656a5f, 32'h4040bbc0} /* (11, 4, 27) {real, imag} */,
  {32'hc1169fee, 32'h41524a57} /* (11, 4, 26) {real, imag} */,
  {32'h3ad44400, 32'h3eabbf40} /* (11, 4, 25) {real, imag} */,
  {32'h4128c649, 32'h410ec217} /* (11, 4, 24) {real, imag} */,
  {32'h4162abd0, 32'h3f5d6ac8} /* (11, 4, 23) {real, imag} */,
  {32'h40c90202, 32'hc104c548} /* (11, 4, 22) {real, imag} */,
  {32'h4005aa08, 32'hc0c40ad4} /* (11, 4, 21) {real, imag} */,
  {32'hbf8566d6, 32'h3fe1d96c} /* (11, 4, 20) {real, imag} */,
  {32'hc0aca51c, 32'hc08255ee} /* (11, 4, 19) {real, imag} */,
  {32'hc15605d2, 32'hc17c2cd0} /* (11, 4, 18) {real, imag} */,
  {32'hc1643016, 32'hc1a7830e} /* (11, 4, 17) {real, imag} */,
  {32'hc0b41cb2, 32'hc0f035a2} /* (11, 4, 16) {real, imag} */,
  {32'h40a35cb1, 32'hbf4ab5e0} /* (11, 4, 15) {real, imag} */,
  {32'h401cb1b1, 32'h41065a2a} /* (11, 4, 14) {real, imag} */,
  {32'hc0bf15a2, 32'h40067ab4} /* (11, 4, 13) {real, imag} */,
  {32'hc13d51f2, 32'h3f111ce2} /* (11, 4, 12) {real, imag} */,
  {32'hbf3eaed2, 32'h40dee758} /* (11, 4, 11) {real, imag} */,
  {32'h4106a761, 32'h412beef9} /* (11, 4, 10) {real, imag} */,
  {32'h411580fd, 32'h41148c02} /* (11, 4, 9) {real, imag} */,
  {32'h40505d2e, 32'h40d30156} /* (11, 4, 8) {real, imag} */,
  {32'hc0a17be4, 32'h3f9c89a2} /* (11, 4, 7) {real, imag} */,
  {32'hbce7c680, 32'h402bdf70} /* (11, 4, 6) {real, imag} */,
  {32'h4112ee78, 32'h4127e6b7} /* (11, 4, 5) {real, imag} */,
  {32'h415f715b, 32'hbd5c0730} /* (11, 4, 4) {real, imag} */,
  {32'hbf39e3aa, 32'hc104595d} /* (11, 4, 3) {real, imag} */,
  {32'h40f68a6a, 32'h3ac4e800} /* (11, 4, 2) {real, imag} */,
  {32'h4111de30, 32'hc00ee224} /* (11, 4, 1) {real, imag} */,
  {32'hbf9b3ab1, 32'hc0404b8b} /* (11, 4, 0) {real, imag} */,
  {32'h40f843d0, 32'hbfbea1f4} /* (11, 3, 31) {real, imag} */,
  {32'h3feef124, 32'h41929c02} /* (11, 3, 30) {real, imag} */,
  {32'hbfbb0ac0, 32'h41990817} /* (11, 3, 29) {real, imag} */,
  {32'h40ba1dfb, 32'h4141b263} /* (11, 3, 28) {real, imag} */,
  {32'h408ae664, 32'h411f660e} /* (11, 3, 27) {real, imag} */,
  {32'h40315488, 32'hbf6a11b0} /* (11, 3, 26) {real, imag} */,
  {32'h4126c714, 32'hc029270a} /* (11, 3, 25) {real, imag} */,
  {32'h4105c153, 32'h40f7590e} /* (11, 3, 24) {real, imag} */,
  {32'h410b1286, 32'h410cf954} /* (11, 3, 23) {real, imag} */,
  {32'h40dda90e, 32'h3f0a4c80} /* (11, 3, 22) {real, imag} */,
  {32'hc08434f1, 32'h40d2343b} /* (11, 3, 21) {real, imag} */,
  {32'hc1407536, 32'hc0d37ed9} /* (11, 3, 20) {real, imag} */,
  {32'hc11a68b2, 32'hc0ad0236} /* (11, 3, 19) {real, imag} */,
  {32'h3f8b52bc, 32'hc0b7fb58} /* (11, 3, 18) {real, imag} */,
  {32'h4033f761, 32'hc0e53efd} /* (11, 3, 17) {real, imag} */,
  {32'hc0ee6ab9, 32'h404ffa8c} /* (11, 3, 16) {real, imag} */,
  {32'h3f68a41c, 32'hc0a0818b} /* (11, 3, 15) {real, imag} */,
  {32'h4108b4a3, 32'hc16a8f3d} /* (11, 3, 14) {real, imag} */,
  {32'h40c1d396, 32'hc139bf0d} /* (11, 3, 13) {real, imag} */,
  {32'h411ea00f, 32'hc00d9e09} /* (11, 3, 12) {real, imag} */,
  {32'h419000ab, 32'h4094bc3b} /* (11, 3, 11) {real, imag} */,
  {32'h3f837f76, 32'h40935aed} /* (11, 3, 10) {real, imag} */,
  {32'hc00a9db0, 32'h40186831} /* (11, 3, 9) {real, imag} */,
  {32'h40cd42cd, 32'h40a2f85a} /* (11, 3, 8) {real, imag} */,
  {32'h417a61d2, 32'h40a1d9d6} /* (11, 3, 7) {real, imag} */,
  {32'h40881659, 32'h40ff5c6d} /* (11, 3, 6) {real, imag} */,
  {32'h40082333, 32'h4080d552} /* (11, 3, 5) {real, imag} */,
  {32'h40452d9f, 32'hc0b8c7b5} /* (11, 3, 4) {real, imag} */,
  {32'h40a5ee2d, 32'hbf6810b4} /* (11, 3, 3) {real, imag} */,
  {32'hc03c204a, 32'hc08a3f3d} /* (11, 3, 2) {real, imag} */,
  {32'hc0bf6505, 32'hc01dd257} /* (11, 3, 1) {real, imag} */,
  {32'hc04adb46, 32'hbfb1d90e} /* (11, 3, 0) {real, imag} */,
  {32'hc1214fc8, 32'h402a644c} /* (11, 2, 31) {real, imag} */,
  {32'hc140f890, 32'hbfeefd78} /* (11, 2, 30) {real, imag} */,
  {32'hc16ec308, 32'h4013c624} /* (11, 2, 29) {real, imag} */,
  {32'hc128924e, 32'h4154b099} /* (11, 2, 28) {real, imag} */,
  {32'hc1182ecc, 32'h415d2a50} /* (11, 2, 27) {real, imag} */,
  {32'hc132e0b6, 32'hc09a658b} /* (11, 2, 26) {real, imag} */,
  {32'hc1aeceed, 32'hc0c6c997} /* (11, 2, 25) {real, imag} */,
  {32'hc119ad65, 32'h40973c42} /* (11, 2, 24) {real, imag} */,
  {32'hc0e02717, 32'hc08e6e7b} /* (11, 2, 23) {real, imag} */,
  {32'hc07c8f40, 32'hc05e21b1} /* (11, 2, 22) {real, imag} */,
  {32'hc0ca60a3, 32'hc11ef3fd} /* (11, 2, 21) {real, imag} */,
  {32'h40d798b9, 32'hc10504bf} /* (11, 2, 20) {real, imag} */,
  {32'h41509cb1, 32'hc0926a30} /* (11, 2, 19) {real, imag} */,
  {32'h4138ff74, 32'hc161cb0c} /* (11, 2, 18) {real, imag} */,
  {32'h41147905, 32'hc193e6ba} /* (11, 2, 17) {real, imag} */,
  {32'h40cc906c, 32'hc14bba2a} /* (11, 2, 16) {real, imag} */,
  {32'h413fee62, 32'hc0900e28} /* (11, 2, 15) {real, imag} */,
  {32'h40cca2f4, 32'h40d2c95c} /* (11, 2, 14) {real, imag} */,
  {32'hc09a5b23, 32'h4040cdac} /* (11, 2, 13) {real, imag} */,
  {32'hbe8a3460, 32'h4043011e} /* (11, 2, 12) {real, imag} */,
  {32'h415b96fe, 32'h400a9438} /* (11, 2, 11) {real, imag} */,
  {32'hc12b416a, 32'h40e292ec} /* (11, 2, 10) {real, imag} */,
  {32'hc19bed1e, 32'h41933092} /* (11, 2, 9) {real, imag} */,
  {32'hc0a5d19f, 32'h408074c8} /* (11, 2, 8) {real, imag} */,
  {32'hbfbabc88, 32'h405ae6b0} /* (11, 2, 7) {real, imag} */,
  {32'hc0045c3e, 32'h418e0739} /* (11, 2, 6) {real, imag} */,
  {32'hbfb91ec6, 32'h40bcf517} /* (11, 2, 5) {real, imag} */,
  {32'hc12238e6, 32'hc08e8657} /* (11, 2, 4) {real, imag} */,
  {32'hbec7c1c8, 32'hbf889cac} /* (11, 2, 3) {real, imag} */,
  {32'h3f4af758, 32'hc050a424} /* (11, 2, 2) {real, imag} */,
  {32'h3f075b38, 32'hc07fbe64} /* (11, 2, 1) {real, imag} */,
  {32'hc09cc3e8, 32'h40819474} /* (11, 2, 0) {real, imag} */,
  {32'h40b6e812, 32'hbf9df060} /* (11, 1, 31) {real, imag} */,
  {32'h411a9073, 32'hc0cd0f2a} /* (11, 1, 30) {real, imag} */,
  {32'h40d7956e, 32'hc16711bb} /* (11, 1, 29) {real, imag} */,
  {32'h4154072c, 32'hc183d9cb} /* (11, 1, 28) {real, imag} */,
  {32'h41970e14, 32'hc0e00684} /* (11, 1, 27) {real, imag} */,
  {32'h4141a288, 32'hbf050d8e} /* (11, 1, 26) {real, imag} */,
  {32'h419c184c, 32'hc0f46ca8} /* (11, 1, 25) {real, imag} */,
  {32'h41857f9e, 32'hc04fbb10} /* (11, 1, 24) {real, imag} */,
  {32'h41c32d49, 32'h4080032a} /* (11, 1, 23) {real, imag} */,
  {32'h41ae8eb4, 32'hc0953814} /* (11, 1, 22) {real, imag} */,
  {32'h410d36ec, 32'hc0f4c2f4} /* (11, 1, 21) {real, imag} */,
  {32'hc127ae8e, 32'hc196c256} /* (11, 1, 20) {real, imag} */,
  {32'hc08cd4a0, 32'hc09b67c2} /* (11, 1, 19) {real, imag} */,
  {32'hc1188da8, 32'hc10be21a} /* (11, 1, 18) {real, imag} */,
  {32'hc11049c5, 32'hc0e91131} /* (11, 1, 17) {real, imag} */,
  {32'hc0ed3556, 32'h4028e2a2} /* (11, 1, 16) {real, imag} */,
  {32'hc101344c, 32'h4060102b} /* (11, 1, 15) {real, imag} */,
  {32'hc17df5d2, 32'h408dd4c2} /* (11, 1, 14) {real, imag} */,
  {32'hc1cbe031, 32'h40b28744} /* (11, 1, 13) {real, imag} */,
  {32'hc1124ea6, 32'h412fce66} /* (11, 1, 12) {real, imag} */,
  {32'h40ed3366, 32'h4150ab38} /* (11, 1, 11) {real, imag} */,
  {32'h41509600, 32'h408649ba} /* (11, 1, 10) {real, imag} */,
  {32'h412cb9f2, 32'hbfbf6960} /* (11, 1, 9) {real, imag} */,
  {32'h414d5a0a, 32'h4191d662} /* (11, 1, 8) {real, imag} */,
  {32'h416a98a7, 32'h41834154} /* (11, 1, 7) {real, imag} */,
  {32'h4098e049, 32'h40fa78fc} /* (11, 1, 6) {real, imag} */,
  {32'hbe7ca180, 32'hc0d3f0b8} /* (11, 1, 5) {real, imag} */,
  {32'h41141d4f, 32'hc18648b4} /* (11, 1, 4) {real, imag} */,
  {32'h41999dee, 32'hc048627c} /* (11, 1, 3) {real, imag} */,
  {32'h419e6828, 32'h40b01672} /* (11, 1, 2) {real, imag} */,
  {32'h3f8e2f90, 32'h40e1f811} /* (11, 1, 1) {real, imag} */,
  {32'h40823d6a, 32'hbfdb411c} /* (11, 1, 0) {real, imag} */,
  {32'h40b6af40, 32'hc0daf393} /* (11, 0, 31) {real, imag} */,
  {32'h41695b8a, 32'hc197efaa} /* (11, 0, 30) {real, imag} */,
  {32'h410397e6, 32'hc0b71338} /* (11, 0, 29) {real, imag} */,
  {32'hc06a048a, 32'h3f6f61c8} /* (11, 0, 28) {real, imag} */,
  {32'hc0c3a028, 32'hc0581343} /* (11, 0, 27) {real, imag} */,
  {32'h3ef56242, 32'hc05a30bc} /* (11, 0, 26) {real, imag} */,
  {32'h40df2e81, 32'hc04d919a} /* (11, 0, 25) {real, imag} */,
  {32'h4170bf0e, 32'h3f52272a} /* (11, 0, 24) {real, imag} */,
  {32'h416fcf63, 32'hc0035ea3} /* (11, 0, 23) {real, imag} */,
  {32'h400fc30b, 32'hc0b651bc} /* (11, 0, 22) {real, imag} */,
  {32'h407df292, 32'hbf08f7fc} /* (11, 0, 21) {real, imag} */,
  {32'hbf5f08b3, 32'h41184886} /* (11, 0, 20) {real, imag} */,
  {32'h3f1c5070, 32'h40783d30} /* (11, 0, 19) {real, imag} */,
  {32'h3e35b4c0, 32'hc150f8aa} /* (11, 0, 18) {real, imag} */,
  {32'hbf002f72, 32'hc13415ba} /* (11, 0, 17) {real, imag} */,
  {32'h40e6bfbd, 32'h3d2ab080} /* (11, 0, 16) {real, imag} */,
  {32'hc06e929a, 32'h41157796} /* (11, 0, 15) {real, imag} */,
  {32'hc0c486ba, 32'h3fbddb20} /* (11, 0, 14) {real, imag} */,
  {32'hc0cc025a, 32'h3f4bdb0a} /* (11, 0, 13) {real, imag} */,
  {32'h3c77c880, 32'h41432352} /* (11, 0, 12) {real, imag} */,
  {32'hc0cff886, 32'h4187efcb} /* (11, 0, 11) {real, imag} */,
  {32'hc0ab3a82, 32'h41062763} /* (11, 0, 10) {real, imag} */,
  {32'hbe9959d8, 32'h40d9625b} /* (11, 0, 9) {real, imag} */,
  {32'hbe599b40, 32'h411d53fb} /* (11, 0, 8) {real, imag} */,
  {32'hc12e8188, 32'h3fa12784} /* (11, 0, 7) {real, imag} */,
  {32'h3f85be44, 32'hc1655fd7} /* (11, 0, 6) {real, imag} */,
  {32'h41811669, 32'hc1a64745} /* (11, 0, 5) {real, imag} */,
  {32'h417725bb, 32'hc0fdf330} /* (11, 0, 4) {real, imag} */,
  {32'h40d5cdbc, 32'hc0b7fdfc} /* (11, 0, 3) {real, imag} */,
  {32'h414a9a80, 32'hc15ee0d4} /* (11, 0, 2) {real, imag} */,
  {32'h41f22ace, 32'hc11d23ee} /* (11, 0, 1) {real, imag} */,
  {32'h41838a36, 32'hc11c4ca4} /* (11, 0, 0) {real, imag} */,
  {32'hc096c503, 32'h40ff6152} /* (10, 31, 31) {real, imag} */,
  {32'h3e3de800, 32'h41a252ea} /* (10, 31, 30) {real, imag} */,
  {32'h3e7e1d00, 32'h41730991} /* (10, 31, 29) {real, imag} */,
  {32'hc06df246, 32'h40ecede2} /* (10, 31, 28) {real, imag} */,
  {32'hc0b52976, 32'h3f1005fc} /* (10, 31, 27) {real, imag} */,
  {32'hc0c5fe48, 32'h3edf74a0} /* (10, 31, 26) {real, imag} */,
  {32'hc0ef563c, 32'h40b34d77} /* (10, 31, 25) {real, imag} */,
  {32'hc18174c5, 32'h41323bb1} /* (10, 31, 24) {real, imag} */,
  {32'hc114ba2a, 32'h41c43118} /* (10, 31, 23) {real, imag} */,
  {32'hbc8fef60, 32'h4148f7f6} /* (10, 31, 22) {real, imag} */,
  {32'h4130c484, 32'h406c2597} /* (10, 31, 21) {real, imag} */,
  {32'h419f9453, 32'hc0c342e8} /* (10, 31, 20) {real, imag} */,
  {32'h41600d40, 32'h3f6c1538} /* (10, 31, 19) {real, imag} */,
  {32'h40b8d497, 32'h4123737e} /* (10, 31, 18) {real, imag} */,
  {32'h3f996c18, 32'hbfe1c7c8} /* (10, 31, 17) {real, imag} */,
  {32'hbeee9ed2, 32'hc15a247e} /* (10, 31, 16) {real, imag} */,
  {32'h4093e6ee, 32'hc12e274e} /* (10, 31, 15) {real, imag} */,
  {32'h40ad7c0e, 32'hc0f88c43} /* (10, 31, 14) {real, imag} */,
  {32'h41625636, 32'hc1635d4e} /* (10, 31, 13) {real, imag} */,
  {32'h4157d830, 32'hc0f1dfe6} /* (10, 31, 12) {real, imag} */,
  {32'h403b3358, 32'h4104998b} /* (10, 31, 11) {real, imag} */,
  {32'h4122d8fe, 32'h415ff886} /* (10, 31, 10) {real, imag} */,
  {32'h40decb58, 32'h41ac1cba} /* (10, 31, 9) {real, imag} */,
  {32'h40812d76, 32'h4187b11b} /* (10, 31, 8) {real, imag} */,
  {32'hc034152a, 32'hc05756a2} /* (10, 31, 7) {real, imag} */,
  {32'h40c1a725, 32'hbdc39500} /* (10, 31, 6) {real, imag} */,
  {32'hc065c524, 32'h4144cc22} /* (10, 31, 5) {real, imag} */,
  {32'hc13ab9ee, 32'h41a366b1} /* (10, 31, 4) {real, imag} */,
  {32'hc0e79b0d, 32'h410669eb} /* (10, 31, 3) {real, imag} */,
  {32'h40612136, 32'hc087107e} /* (10, 31, 2) {real, imag} */,
  {32'h415c4818, 32'hbe5ce860} /* (10, 31, 1) {real, imag} */,
  {32'h40b074ae, 32'h401e0980} /* (10, 31, 0) {real, imag} */,
  {32'h410a5272, 32'hc0a585db} /* (10, 30, 31) {real, imag} */,
  {32'h41bc313b, 32'hc18b58aa} /* (10, 30, 30) {real, imag} */,
  {32'h404f562a, 32'hc183f0bf} /* (10, 30, 29) {real, imag} */,
  {32'h4061a2a2, 32'hc114a39e} /* (10, 30, 28) {real, imag} */,
  {32'hc0658aa4, 32'hbfcc5ee8} /* (10, 30, 27) {real, imag} */,
  {32'hc0cfd1b2, 32'hc040f922} /* (10, 30, 26) {real, imag} */,
  {32'hc00c56d6, 32'h40d8f752} /* (10, 30, 25) {real, imag} */,
  {32'hc114c834, 32'h41041ea7} /* (10, 30, 24) {real, imag} */,
  {32'h415b9093, 32'h3f1247c2} /* (10, 30, 23) {real, imag} */,
  {32'h41c1c920, 32'hc09ca330} /* (10, 30, 22) {real, imag} */,
  {32'h412c54a7, 32'hc01f4e6e} /* (10, 30, 21) {real, imag} */,
  {32'hc0eb559e, 32'h404a5b1c} /* (10, 30, 20) {real, imag} */,
  {32'hc150ff98, 32'hc05074bd} /* (10, 30, 19) {real, imag} */,
  {32'hc0e3665e, 32'hc0623c5c} /* (10, 30, 18) {real, imag} */,
  {32'hbfe9f790, 32'h3fff862c} /* (10, 30, 17) {real, imag} */,
  {32'hc05e310c, 32'h40a1c79d} /* (10, 30, 16) {real, imag} */,
  {32'hc0cd3126, 32'h40677950} /* (10, 30, 15) {real, imag} */,
  {32'h402d9cac, 32'h3f006a80} /* (10, 30, 14) {real, imag} */,
  {32'h404dace0, 32'hbf92965a} /* (10, 30, 13) {real, imag} */,
  {32'h412eba62, 32'hc04b20ac} /* (10, 30, 12) {real, imag} */,
  {32'h40272429, 32'hc12a283b} /* (10, 30, 11) {real, imag} */,
  {32'h40ee0e55, 32'hc16ef9d1} /* (10, 30, 10) {real, imag} */,
  {32'h419a0bed, 32'hc10d2cb2} /* (10, 30, 9) {real, imag} */,
  {32'h418b4297, 32'h4115a29f} /* (10, 30, 8) {real, imag} */,
  {32'h41887059, 32'h4130fe35} /* (10, 30, 7) {real, imag} */,
  {32'h41ad3212, 32'h3fde1cf6} /* (10, 30, 6) {real, imag} */,
  {32'h4197bc1b, 32'h3f832530} /* (10, 30, 5) {real, imag} */,
  {32'h3f9b5660, 32'h40b843d0} /* (10, 30, 4) {real, imag} */,
  {32'h3fdb5d90, 32'h40015aba} /* (10, 30, 3) {real, imag} */,
  {32'h3cf47b00, 32'h406fce08} /* (10, 30, 2) {real, imag} */,
  {32'h3f2708a0, 32'h40d62e00} /* (10, 30, 1) {real, imag} */,
  {32'hbf19b18a, 32'h404672f2} /* (10, 30, 0) {real, imag} */,
  {32'hc10d59ec, 32'hc143bb94} /* (10, 29, 31) {real, imag} */,
  {32'hc191dbb0, 32'hc1bf1cf4} /* (10, 29, 30) {real, imag} */,
  {32'hc1383459, 32'hc1357bc2} /* (10, 29, 29) {real, imag} */,
  {32'hc000c8d3, 32'hbf978d10} /* (10, 29, 28) {real, imag} */,
  {32'h408e7999, 32'h40250a4a} /* (10, 29, 27) {real, imag} */,
  {32'h3eacc238, 32'h3ffa0246} /* (10, 29, 26) {real, imag} */,
  {32'hc100a744, 32'h40bed30b} /* (10, 29, 25) {real, imag} */,
  {32'hc0114c4d, 32'h3f2d04fd} /* (10, 29, 24) {real, imag} */,
  {32'hc0e381f6, 32'hc051ed03} /* (10, 29, 23) {real, imag} */,
  {32'h40e24a8a, 32'h3eed0674} /* (10, 29, 22) {real, imag} */,
  {32'h40a4616f, 32'h41192f85} /* (10, 29, 21) {real, imag} */,
  {32'hbf2e1f30, 32'h3fec83b6} /* (10, 29, 20) {real, imag} */,
  {32'h3fbd638b, 32'hc050fe22} /* (10, 29, 19) {real, imag} */,
  {32'h40f76d1d, 32'hc0dffdce} /* (10, 29, 18) {real, imag} */,
  {32'hbfbb2ab0, 32'hc1023a5f} /* (10, 29, 17) {real, imag} */,
  {32'h40a99281, 32'hbddea820} /* (10, 29, 16) {real, imag} */,
  {32'h40fd8d35, 32'hbe1c33c0} /* (10, 29, 15) {real, imag} */,
  {32'hbd9e1e20, 32'hc1051956} /* (10, 29, 14) {real, imag} */,
  {32'hc0510f26, 32'hc0116748} /* (10, 29, 13) {real, imag} */,
  {32'hc0c8a60f, 32'h4018fca0} /* (10, 29, 12) {real, imag} */,
  {32'h40ab1801, 32'h40468754} /* (10, 29, 11) {real, imag} */,
  {32'hc0c1013f, 32'h40109dde} /* (10, 29, 10) {real, imag} */,
  {32'hc0e8257e, 32'h3f63c440} /* (10, 29, 9) {real, imag} */,
  {32'h4120645c, 32'hbee9f250} /* (10, 29, 8) {real, imag} */,
  {32'h40f80b94, 32'hc099913b} /* (10, 29, 7) {real, imag} */,
  {32'hc039da1a, 32'hc09e94a6} /* (10, 29, 6) {real, imag} */,
  {32'hc134637a, 32'hbf70e80c} /* (10, 29, 5) {real, imag} */,
  {32'hc0f03879, 32'hc10c59d6} /* (10, 29, 4) {real, imag} */,
  {32'hc0e1b805, 32'hc1141bf3} /* (10, 29, 3) {real, imag} */,
  {32'h404d7d6c, 32'hc123220c} /* (10, 29, 2) {real, imag} */,
  {32'hc12cbdda, 32'hc0e03891} /* (10, 29, 1) {real, imag} */,
  {32'hc144d65b, 32'hc006d46b} /* (10, 29, 0) {real, imag} */,
  {32'hbfd61dd8, 32'h3e104f30} /* (10, 28, 31) {real, imag} */,
  {32'hbfa5c8fa, 32'hc0852617} /* (10, 28, 30) {real, imag} */,
  {32'h409c5284, 32'hc12d2e10} /* (10, 28, 29) {real, imag} */,
  {32'h40849867, 32'hc001c394} /* (10, 28, 28) {real, imag} */,
  {32'hbfd6f90f, 32'h41513572} /* (10, 28, 27) {real, imag} */,
  {32'hc00746b4, 32'h40de5261} /* (10, 28, 26) {real, imag} */,
  {32'hc0457342, 32'h40081d5c} /* (10, 28, 25) {real, imag} */,
  {32'h3f697924, 32'h411f0e5a} /* (10, 28, 24) {real, imag} */,
  {32'h408299df, 32'h4082f0a4} /* (10, 28, 23) {real, imag} */,
  {32'hc1287b5a, 32'hc0d5fe37} /* (10, 28, 22) {real, imag} */,
  {32'hc08dee50, 32'h4052cfac} /* (10, 28, 21) {real, imag} */,
  {32'h40a0546f, 32'hbf9e9c98} /* (10, 28, 20) {real, imag} */,
  {32'hc0bdaf02, 32'hbfe2e4f6} /* (10, 28, 19) {real, imag} */,
  {32'hc115cd5e, 32'h40e8588d} /* (10, 28, 18) {real, imag} */,
  {32'hc0dd8cd9, 32'h4071820e} /* (10, 28, 17) {real, imag} */,
  {32'hc175f102, 32'h401e0c98} /* (10, 28, 16) {real, imag} */,
  {32'h409aa0ac, 32'hbf46e12c} /* (10, 28, 15) {real, imag} */,
  {32'h4025125a, 32'hc153f25c} /* (10, 28, 14) {real, imag} */,
  {32'h41065f5c, 32'hc150cde8} /* (10, 28, 13) {real, imag} */,
  {32'h4106b818, 32'hc113de07} /* (10, 28, 12) {real, imag} */,
  {32'hc106e1c7, 32'h3f9d4020} /* (10, 28, 11) {real, imag} */,
  {32'hbf27620c, 32'h41689119} /* (10, 28, 10) {real, imag} */,
  {32'h4044f23e, 32'h418403ee} /* (10, 28, 9) {real, imag} */,
  {32'hc060d008, 32'h40e44ae6} /* (10, 28, 8) {real, imag} */,
  {32'hc0be0993, 32'hbda71b00} /* (10, 28, 7) {real, imag} */,
  {32'h3faea8ef, 32'hbfb6bfe8} /* (10, 28, 6) {real, imag} */,
  {32'h413b9612, 32'h411fe116} /* (10, 28, 5) {real, imag} */,
  {32'h4195d70e, 32'h40c29046} /* (10, 28, 4) {real, imag} */,
  {32'h40e444e2, 32'h3f201f98} /* (10, 28, 3) {real, imag} */,
  {32'hc03eb978, 32'h3f778673} /* (10, 28, 2) {real, imag} */,
  {32'hc0ee1eac, 32'hc04a8e4f} /* (10, 28, 1) {real, imag} */,
  {32'hc0f2debd, 32'h3fbcc3d2} /* (10, 28, 0) {real, imag} */,
  {32'hbf70c65a, 32'hc051fadc} /* (10, 27, 31) {real, imag} */,
  {32'h40233be8, 32'hbfb997fc} /* (10, 27, 30) {real, imag} */,
  {32'hc055d092, 32'hc034fa13} /* (10, 27, 29) {real, imag} */,
  {32'hc00ce30a, 32'h41051014} /* (10, 27, 28) {real, imag} */,
  {32'h4112de89, 32'h40e1f864} /* (10, 27, 27) {real, imag} */,
  {32'h40f7ae66, 32'hc036ee87} /* (10, 27, 26) {real, imag} */,
  {32'h40c317a6, 32'hc105c489} /* (10, 27, 25) {real, imag} */,
  {32'h3f9ede84, 32'hbf5b1fa8} /* (10, 27, 24) {real, imag} */,
  {32'h3fa70c70, 32'h40b2e690} /* (10, 27, 23) {real, imag} */,
  {32'hc0177c22, 32'h40089164} /* (10, 27, 22) {real, imag} */,
  {32'h4128680f, 32'h3ed29cd0} /* (10, 27, 21) {real, imag} */,
  {32'h41513114, 32'h3d03faa0} /* (10, 27, 20) {real, imag} */,
  {32'h409adc28, 32'hc0bae45a} /* (10, 27, 19) {real, imag} */,
  {32'hbfefe068, 32'hc0e9b0fd} /* (10, 27, 18) {real, imag} */,
  {32'hbfea0d48, 32'hc084124e} /* (10, 27, 17) {real, imag} */,
  {32'hc0ab611a, 32'hc01e30ba} /* (10, 27, 16) {real, imag} */,
  {32'h4066958c, 32'h4077315d} /* (10, 27, 15) {real, imag} */,
  {32'h41598c54, 32'h414d1adf} /* (10, 27, 14) {real, imag} */,
  {32'h400d8319, 32'h41075df5} /* (10, 27, 13) {real, imag} */,
  {32'hc0e0a534, 32'hbde041b0} /* (10, 27, 12) {real, imag} */,
  {32'hc023210e, 32'hc06101aa} /* (10, 27, 11) {real, imag} */,
  {32'hc0817389, 32'hc0b43b67} /* (10, 27, 10) {real, imag} */,
  {32'hbe1a0fb0, 32'hc120ad78} /* (10, 27, 9) {real, imag} */,
  {32'hc0559d55, 32'h3f5cebb4} /* (10, 27, 8) {real, imag} */,
  {32'h409307c4, 32'h413107d8} /* (10, 27, 7) {real, imag} */,
  {32'h406220e0, 32'h41274138} /* (10, 27, 6) {real, imag} */,
  {32'h404ae150, 32'h41764cfa} /* (10, 27, 5) {real, imag} */,
  {32'h3f92ca5e, 32'h4118e115} /* (10, 27, 4) {real, imag} */,
  {32'h40442152, 32'h3fc9d79e} /* (10, 27, 3) {real, imag} */,
  {32'hc09d0087, 32'h4050dd6b} /* (10, 27, 2) {real, imag} */,
  {32'hc045621a, 32'h40149981} /* (10, 27, 1) {real, imag} */,
  {32'hbe770710, 32'hbfd5fbe2} /* (10, 27, 0) {real, imag} */,
  {32'hc05c88cc, 32'hbe834d6c} /* (10, 26, 31) {real, imag} */,
  {32'hc10bab71, 32'hc0b8b422} /* (10, 26, 30) {real, imag} */,
  {32'h40e48e1f, 32'hc085735a} /* (10, 26, 29) {real, imag} */,
  {32'h41397a76, 32'hc0d1ee84} /* (10, 26, 28) {real, imag} */,
  {32'h40b5603c, 32'hc1307510} /* (10, 26, 27) {real, imag} */,
  {32'hbfb46ccb, 32'hc0f0dcc7} /* (10, 26, 26) {real, imag} */,
  {32'hc10c4124, 32'hbfdd485d} /* (10, 26, 25) {real, imag} */,
  {32'hbf5d7db0, 32'h3fa09434} /* (10, 26, 24) {real, imag} */,
  {32'h410ddd25, 32'h410b3f92} /* (10, 26, 23) {real, imag} */,
  {32'h4127661d, 32'h40db33fe} /* (10, 26, 22) {real, imag} */,
  {32'h404330ca, 32'h40578ab5} /* (10, 26, 21) {real, imag} */,
  {32'h3fd6b482, 32'h3f85ddc4} /* (10, 26, 20) {real, imag} */,
  {32'hbfd893c0, 32'hc050fc4e} /* (10, 26, 19) {real, imag} */,
  {32'hc11ffcb7, 32'hc181042d} /* (10, 26, 18) {real, imag} */,
  {32'hc05dd3e2, 32'hc1063d89} /* (10, 26, 17) {real, imag} */,
  {32'hc030a7e1, 32'h3f9dcf9c} /* (10, 26, 16) {real, imag} */,
  {32'h3f15a710, 32'h40909f5a} /* (10, 26, 15) {real, imag} */,
  {32'h3fac1d3a, 32'hbfd691f8} /* (10, 26, 14) {real, imag} */,
  {32'h4050af1a, 32'hc11962e8} /* (10, 26, 13) {real, imag} */,
  {32'h4055dbd8, 32'hc0259cf5} /* (10, 26, 12) {real, imag} */,
  {32'h40ca3a04, 32'hbfc73a3d} /* (10, 26, 11) {real, imag} */,
  {32'h415e592e, 32'h3f7e15dc} /* (10, 26, 10) {real, imag} */,
  {32'h40b3f9de, 32'hbfbe690d} /* (10, 26, 9) {real, imag} */,
  {32'h40216d28, 32'hc0a9fd9a} /* (10, 26, 8) {real, imag} */,
  {32'hc0825f5d, 32'hbd4f4800} /* (10, 26, 7) {real, imag} */,
  {32'hc0d3eac8, 32'h400c5045} /* (10, 26, 6) {real, imag} */,
  {32'h40ede778, 32'hc0571c4c} /* (10, 26, 5) {real, imag} */,
  {32'h4004f3d6, 32'h40829893} /* (10, 26, 4) {real, imag} */,
  {32'h40bf9cea, 32'h405dda62} /* (10, 26, 3) {real, imag} */,
  {32'h40d5eb78, 32'h400d17d8} /* (10, 26, 2) {real, imag} */,
  {32'hc003bb2a, 32'hbee4b380} /* (10, 26, 1) {real, imag} */,
  {32'h407895a5, 32'hc00a4224} /* (10, 26, 0) {real, imag} */,
  {32'h3f3561f6, 32'h3fa31fae} /* (10, 25, 31) {real, imag} */,
  {32'hc03f8040, 32'h40d0a01d} /* (10, 25, 30) {real, imag} */,
  {32'hc129b641, 32'h41121deb} /* (10, 25, 29) {real, imag} */,
  {32'hc0823e1d, 32'h3f792570} /* (10, 25, 28) {real, imag} */,
  {32'h405c3216, 32'h40f965d7} /* (10, 25, 27) {real, imag} */,
  {32'h40c4811f, 32'h410bde66} /* (10, 25, 26) {real, imag} */,
  {32'h40cc8980, 32'h403ec611} /* (10, 25, 25) {real, imag} */,
  {32'h40070b1e, 32'h407454ae} /* (10, 25, 24) {real, imag} */,
  {32'h3f349e02, 32'h4093d0aa} /* (10, 25, 23) {real, imag} */,
  {32'hc0ba6e6d, 32'hc0a56800} /* (10, 25, 22) {real, imag} */,
  {32'h40d88ab2, 32'hbf9d5e22} /* (10, 25, 21) {real, imag} */,
  {32'h410824a9, 32'h40894cab} /* (10, 25, 20) {real, imag} */,
  {32'h405bc68e, 32'h40b061c0} /* (10, 25, 19) {real, imag} */,
  {32'hc08e0cbc, 32'h40f7fb3d} /* (10, 25, 18) {real, imag} */,
  {32'hc023222a, 32'h4089c27b} /* (10, 25, 17) {real, imag} */,
  {32'hc04ce4eb, 32'h3e333c00} /* (10, 25, 16) {real, imag} */,
  {32'hc0cad170, 32'hbe29f838} /* (10, 25, 15) {real, imag} */,
  {32'h405255a7, 32'h40ba80d0} /* (10, 25, 14) {real, imag} */,
  {32'hbf105e14, 32'hbfb929a4} /* (10, 25, 13) {real, imag} */,
  {32'hc13cd68a, 32'hc115e1ec} /* (10, 25, 12) {real, imag} */,
  {32'hc100b846, 32'hc11d4782} /* (10, 25, 11) {real, imag} */,
  {32'hc0c7a33c, 32'h4098b283} /* (10, 25, 10) {real, imag} */,
  {32'hc0e484cc, 32'h4161e458} /* (10, 25, 9) {real, imag} */,
  {32'hbfd83240, 32'h40ac9075} /* (10, 25, 8) {real, imag} */,
  {32'h400429c2, 32'hc068abec} /* (10, 25, 7) {real, imag} */,
  {32'h3eb26dec, 32'hc0e5e058} /* (10, 25, 6) {real, imag} */,
  {32'hc0948442, 32'h3ffaa932} /* (10, 25, 5) {real, imag} */,
  {32'hbfe215d4, 32'h3f94d77a} /* (10, 25, 4) {real, imag} */,
  {32'hbe1ad220, 32'hc0a52bc1} /* (10, 25, 3) {real, imag} */,
  {32'h404227d2, 32'hc1295b8f} /* (10, 25, 2) {real, imag} */,
  {32'h4109f535, 32'hc128cdd2} /* (10, 25, 1) {real, imag} */,
  {32'h3f3fd8dc, 32'hc08023e0} /* (10, 25, 0) {real, imag} */,
  {32'h3fbc36de, 32'h40363550} /* (10, 24, 31) {real, imag} */,
  {32'h40265748, 32'hbfa5ca14} /* (10, 24, 30) {real, imag} */,
  {32'h401c16ea, 32'h40844890} /* (10, 24, 29) {real, imag} */,
  {32'hbf009f00, 32'hbfdf7e5c} /* (10, 24, 28) {real, imag} */,
  {32'hbfd2ea94, 32'hc0963445} /* (10, 24, 27) {real, imag} */,
  {32'h406bd618, 32'hbf9d7c17} /* (10, 24, 26) {real, imag} */,
  {32'hbf9c3686, 32'h40828136} /* (10, 24, 25) {real, imag} */,
  {32'hc0d04d02, 32'h3d3fe380} /* (10, 24, 24) {real, imag} */,
  {32'hc1069f3c, 32'h4019ea0f} /* (10, 24, 23) {real, imag} */,
  {32'hc119f26d, 32'hc0684636} /* (10, 24, 22) {real, imag} */,
  {32'h3f0ec7d8, 32'h406e4e1d} /* (10, 24, 21) {real, imag} */,
  {32'h40f5672b, 32'hbd32bd40} /* (10, 24, 20) {real, imag} */,
  {32'h40ad5b3f, 32'h406caf8c} /* (10, 24, 19) {real, imag} */,
  {32'h408e8a48, 32'h40e00847} /* (10, 24, 18) {real, imag} */,
  {32'hc0305b86, 32'h40e11372} /* (10, 24, 17) {real, imag} */,
  {32'hc11373cf, 32'h4089348a} /* (10, 24, 16) {real, imag} */,
  {32'hc1037dc0, 32'h3c9fae80} /* (10, 24, 15) {real, imag} */,
  {32'hbf2af760, 32'hc093a99c} /* (10, 24, 14) {real, imag} */,
  {32'hbebdb846, 32'hbfebdcde} /* (10, 24, 13) {real, imag} */,
  {32'hc08a673d, 32'h4025369b} /* (10, 24, 12) {real, imag} */,
  {32'hc07aa8d2, 32'hbe552080} /* (10, 24, 11) {real, imag} */,
  {32'hbf29ac08, 32'h405779d0} /* (10, 24, 10) {real, imag} */,
  {32'h410ff557, 32'hc129fd86} /* (10, 24, 9) {real, imag} */,
  {32'h416e483e, 32'hc0f8402e} /* (10, 24, 8) {real, imag} */,
  {32'h4131c190, 32'hc002597e} /* (10, 24, 7) {real, imag} */,
  {32'hc0e33b6b, 32'h401eb30a} /* (10, 24, 6) {real, imag} */,
  {32'hc10f3c72, 32'hba851400} /* (10, 24, 5) {real, imag} */,
  {32'hbea07308, 32'h4043b399} /* (10, 24, 4) {real, imag} */,
  {32'h3fcc60e2, 32'hc08b61ca} /* (10, 24, 3) {real, imag} */,
  {32'h40ea6fb2, 32'h3ff3f8b0} /* (10, 24, 2) {real, imag} */,
  {32'h3effcd10, 32'h3fcbad4c} /* (10, 24, 1) {real, imag} */,
  {32'hc02877f4, 32'h4019eb9c} /* (10, 24, 0) {real, imag} */,
  {32'hbecef1a4, 32'h3f88bc28} /* (10, 23, 31) {real, imag} */,
  {32'h40993594, 32'hbfa9c196} /* (10, 23, 30) {real, imag} */,
  {32'hbedc77f0, 32'hc014c1d4} /* (10, 23, 29) {real, imag} */,
  {32'hc0c5b68b, 32'hc09ccbab} /* (10, 23, 28) {real, imag} */,
  {32'hc0db6616, 32'hc0f03bf5} /* (10, 23, 27) {real, imag} */,
  {32'hc01be1e2, 32'h408348d2} /* (10, 23, 26) {real, imag} */,
  {32'hc0bfbe48, 32'h408bbd77} /* (10, 23, 25) {real, imag} */,
  {32'hc0049c48, 32'hc1087810} /* (10, 23, 24) {real, imag} */,
  {32'h40316a87, 32'hbfd73ffa} /* (10, 23, 23) {real, imag} */,
  {32'h3f524e62, 32'h4073bd4a} /* (10, 23, 22) {real, imag} */,
  {32'h3f88f21f, 32'hbfa4eb24} /* (10, 23, 21) {real, imag} */,
  {32'hbfef8938, 32'h40a30830} /* (10, 23, 20) {real, imag} */,
  {32'hc0c468d2, 32'h4098ea78} /* (10, 23, 19) {real, imag} */,
  {32'h3f25e2a0, 32'h400b1d16} /* (10, 23, 18) {real, imag} */,
  {32'h408de3e0, 32'hc0a221b5} /* (10, 23, 17) {real, imag} */,
  {32'h40104b09, 32'hc0de9ece} /* (10, 23, 16) {real, imag} */,
  {32'hc0c3ba49, 32'hc0a14d6b} /* (10, 23, 15) {real, imag} */,
  {32'hc0ed92c6, 32'hc0bfd90c} /* (10, 23, 14) {real, imag} */,
  {32'h3e8c1658, 32'hc0bb0763} /* (10, 23, 13) {real, imag} */,
  {32'hbf4d9830, 32'hbf203a44} /* (10, 23, 12) {real, imag} */,
  {32'h4017a053, 32'h3f28c4d8} /* (10, 23, 11) {real, imag} */,
  {32'h3e94df18, 32'hc00eb432} /* (10, 23, 10) {real, imag} */,
  {32'hbf904d56, 32'h40f73adc} /* (10, 23, 9) {real, imag} */,
  {32'h4094dd9a, 32'h40e35cff} /* (10, 23, 8) {real, imag} */,
  {32'h40092058, 32'hc0bdf6a4} /* (10, 23, 7) {real, imag} */,
  {32'h3fcf73ec, 32'hc04712a7} /* (10, 23, 6) {real, imag} */,
  {32'h4102291b, 32'hbf90c532} /* (10, 23, 5) {real, imag} */,
  {32'h402bb502, 32'h40df91ba} /* (10, 23, 4) {real, imag} */,
  {32'h40023b36, 32'h40bbdb29} /* (10, 23, 3) {real, imag} */,
  {32'h4045ff25, 32'h409d24e0} /* (10, 23, 2) {real, imag} */,
  {32'hbf31f9da, 32'h3f408328} /* (10, 23, 1) {real, imag} */,
  {32'h40242761, 32'hc01426a8} /* (10, 23, 0) {real, imag} */,
  {32'h405b8574, 32'hbf64c0e1} /* (10, 22, 31) {real, imag} */,
  {32'h403cc43e, 32'h400266b9} /* (10, 22, 30) {real, imag} */,
  {32'hbf1bc7b8, 32'h3ff84450} /* (10, 22, 29) {real, imag} */,
  {32'h40176a5a, 32'hbef0d1c8} /* (10, 22, 28) {real, imag} */,
  {32'hbfd5c1a0, 32'hc0295a4f} /* (10, 22, 27) {real, imag} */,
  {32'h40807dd4, 32'hc082a12c} /* (10, 22, 26) {real, imag} */,
  {32'h40d0f83c, 32'hc03550c9} /* (10, 22, 25) {real, imag} */,
  {32'h400dd97b, 32'hc030ba36} /* (10, 22, 24) {real, imag} */,
  {32'hbf37420c, 32'h3f1ac7ca} /* (10, 22, 23) {real, imag} */,
  {32'hc0ca9f9a, 32'h3e37d970} /* (10, 22, 22) {real, imag} */,
  {32'hc1026ece, 32'hc0b49384} /* (10, 22, 21) {real, imag} */,
  {32'hc027e6da, 32'hc104049f} /* (10, 22, 20) {real, imag} */,
  {32'h404cd90e, 32'hc08b2a2b} /* (10, 22, 19) {real, imag} */,
  {32'h408c693a, 32'hbec3cb00} /* (10, 22, 18) {real, imag} */,
  {32'hbfc6a896, 32'hbf0f7940} /* (10, 22, 17) {real, imag} */,
  {32'h40218e24, 32'hc09240e2} /* (10, 22, 16) {real, imag} */,
  {32'h401a0828, 32'hbfd57c9e} /* (10, 22, 15) {real, imag} */,
  {32'h3f9685ef, 32'h4028f44c} /* (10, 22, 14) {real, imag} */,
  {32'h402488b6, 32'hbe418b44} /* (10, 22, 13) {real, imag} */,
  {32'hbfb4b5de, 32'hc092c153} /* (10, 22, 12) {real, imag} */,
  {32'h3fe17db8, 32'h3f54cc46} /* (10, 22, 11) {real, imag} */,
  {32'h40235d0f, 32'hbedefba8} /* (10, 22, 10) {real, imag} */,
  {32'h40825bd8, 32'h408030a8} /* (10, 22, 9) {real, imag} */,
  {32'h3e1b0100, 32'h4085174c} /* (10, 22, 8) {real, imag} */,
  {32'h3d771b00, 32'hc08f3682} /* (10, 22, 7) {real, imag} */,
  {32'h4003b535, 32'hc0896aca} /* (10, 22, 6) {real, imag} */,
  {32'h3f4dd82e, 32'hc08aadff} /* (10, 22, 5) {real, imag} */,
  {32'hbe6cdb90, 32'hbff0f7c6} /* (10, 22, 4) {real, imag} */,
  {32'hbf87b230, 32'hbfd5f7c8} /* (10, 22, 3) {real, imag} */,
  {32'hc08a1436, 32'h403a63fa} /* (10, 22, 2) {real, imag} */,
  {32'hc005d631, 32'h40271214} /* (10, 22, 1) {real, imag} */,
  {32'hc0308d5f, 32'hc0906560} /* (10, 22, 0) {real, imag} */,
  {32'h3ff8bfc5, 32'hbffd7975} /* (10, 21, 31) {real, imag} */,
  {32'h3e80e9cc, 32'hc01dba0c} /* (10, 21, 30) {real, imag} */,
  {32'h3cc8ff00, 32'h3e81c898} /* (10, 21, 29) {real, imag} */,
  {32'hc083deba, 32'hc07074f4} /* (10, 21, 28) {real, imag} */,
  {32'hbf5e5838, 32'hc02ed0b0} /* (10, 21, 27) {real, imag} */,
  {32'h40c56f36, 32'h3f388be4} /* (10, 21, 26) {real, imag} */,
  {32'h3fd138fc, 32'hbf585d13} /* (10, 21, 25) {real, imag} */,
  {32'h406b0136, 32'h4018cfba} /* (10, 21, 24) {real, imag} */,
  {32'h405c4196, 32'h40735a16} /* (10, 21, 23) {real, imag} */,
  {32'h40a2fdc4, 32'h3ffc1466} /* (10, 21, 22) {real, imag} */,
  {32'h40b12909, 32'h3f063de8} /* (10, 21, 21) {real, imag} */,
  {32'h4099ff54, 32'h408e95ca} /* (10, 21, 20) {real, imag} */,
  {32'h3feeb80c, 32'h402e6182} /* (10, 21, 19) {real, imag} */,
  {32'hc00769da, 32'h3f3d2a72} /* (10, 21, 18) {real, imag} */,
  {32'hbeebe674, 32'hc0484abc} /* (10, 21, 17) {real, imag} */,
  {32'hbf58fb60, 32'hbf984c7f} /* (10, 21, 16) {real, imag} */,
  {32'h40e4d429, 32'hc0887be4} /* (10, 21, 15) {real, imag} */,
  {32'h40e30f26, 32'hc105aad9} /* (10, 21, 14) {real, imag} */,
  {32'hbffb019a, 32'hc006d106} /* (10, 21, 13) {real, imag} */,
  {32'h3fbf48da, 32'h40c39b87} /* (10, 21, 12) {real, imag} */,
  {32'h3ffb0bc3, 32'h3e7ad448} /* (10, 21, 11) {real, imag} */,
  {32'h3f896f51, 32'hc0b0aa81} /* (10, 21, 10) {real, imag} */,
  {32'hc01048de, 32'hc0d40712} /* (10, 21, 9) {real, imag} */,
  {32'h3ff99332, 32'hc067d170} /* (10, 21, 8) {real, imag} */,
  {32'h3e949a9e, 32'h3ffc94c8} /* (10, 21, 7) {real, imag} */,
  {32'hc028c581, 32'h40458494} /* (10, 21, 6) {real, imag} */,
  {32'hc0220bf6, 32'h3f6241b4} /* (10, 21, 5) {real, imag} */,
  {32'h4029fd8d, 32'hc084925f} /* (10, 21, 4) {real, imag} */,
  {32'h404da81e, 32'hc0c885fc} /* (10, 21, 3) {real, imag} */,
  {32'h3f9b66b8, 32'h3d7ae180} /* (10, 21, 2) {real, imag} */,
  {32'hc03c793b, 32'h407ec9c9} /* (10, 21, 1) {real, imag} */,
  {32'hbe7cc9e0, 32'h407fce72} /* (10, 21, 0) {real, imag} */,
  {32'h3ffbf5b9, 32'h3fde0684} /* (10, 20, 31) {real, imag} */,
  {32'h3fdcbe93, 32'h40013df4} /* (10, 20, 30) {real, imag} */,
  {32'hc0029084, 32'h406f9546} /* (10, 20, 29) {real, imag} */,
  {32'h40961e4e, 32'h40dd53e8} /* (10, 20, 28) {real, imag} */,
  {32'h40c1572a, 32'h3fbc46aa} /* (10, 20, 27) {real, imag} */,
  {32'h409e5758, 32'hbf8ea73e} /* (10, 20, 26) {real, imag} */,
  {32'h3fbda064, 32'hbdadbc10} /* (10, 20, 25) {real, imag} */,
  {32'hbff9b7ad, 32'h4042d3be} /* (10, 20, 24) {real, imag} */,
  {32'hbe8901e0, 32'h401ba885} /* (10, 20, 23) {real, imag} */,
  {32'hbf86dc98, 32'h407953ea} /* (10, 20, 22) {real, imag} */,
  {32'hc0498174, 32'h4026fe25} /* (10, 20, 21) {real, imag} */,
  {32'hbfe20546, 32'hc01071a0} /* (10, 20, 20) {real, imag} */,
  {32'hbfef410a, 32'h3f0d15f0} /* (10, 20, 19) {real, imag} */,
  {32'h4059cd78, 32'h3ede4ff8} /* (10, 20, 18) {real, imag} */,
  {32'h4083ebd1, 32'h3ef3eccc} /* (10, 20, 17) {real, imag} */,
  {32'h403fb040, 32'hc04d0466} /* (10, 20, 16) {real, imag} */,
  {32'h3d236b80, 32'hc02686d6} /* (10, 20, 15) {real, imag} */,
  {32'hbf4a2d90, 32'h3f06cc6e} /* (10, 20, 14) {real, imag} */,
  {32'hc018ca4c, 32'h40614a38} /* (10, 20, 13) {real, imag} */,
  {32'h3fe8a7c9, 32'h3fcff7ba} /* (10, 20, 12) {real, imag} */,
  {32'hc0464d92, 32'hc01a4a02} /* (10, 20, 11) {real, imag} */,
  {32'hc01d2a32, 32'hc0978284} /* (10, 20, 10) {real, imag} */,
  {32'hc01a75b2, 32'hc0a4f43f} /* (10, 20, 9) {real, imag} */,
  {32'h3fc76d1d, 32'h4079f87b} /* (10, 20, 8) {real, imag} */,
  {32'h3f5a68fd, 32'h406b4cc7} /* (10, 20, 7) {real, imag} */,
  {32'hbf58aed6, 32'h400d07eb} /* (10, 20, 6) {real, imag} */,
  {32'hbee26cc8, 32'h3fd630b0} /* (10, 20, 5) {real, imag} */,
  {32'h3f9e1353, 32'h3ebc6548} /* (10, 20, 4) {real, imag} */,
  {32'h3f03bab4, 32'h40a79bec} /* (10, 20, 3) {real, imag} */,
  {32'h3f0062d0, 32'h40042791} /* (10, 20, 2) {real, imag} */,
  {32'hc026c023, 32'hc0457244} /* (10, 20, 1) {real, imag} */,
  {32'hbf847d34, 32'hbf47e622} /* (10, 20, 0) {real, imag} */,
  {32'hbf1328dc, 32'hbebaf958} /* (10, 19, 31) {real, imag} */,
  {32'hc0300a55, 32'h3f482528} /* (10, 19, 30) {real, imag} */,
  {32'hbffd9118, 32'h3f3f093a} /* (10, 19, 29) {real, imag} */,
  {32'h402ff038, 32'h400d078e} /* (10, 19, 28) {real, imag} */,
  {32'h4003f97c, 32'hbef70818} /* (10, 19, 27) {real, imag} */,
  {32'hbf6b3d6b, 32'hc1001603} /* (10, 19, 26) {real, imag} */,
  {32'hbf94d084, 32'hc08e12a4} /* (10, 19, 25) {real, imag} */,
  {32'hc05a4284, 32'hc097264e} /* (10, 19, 24) {real, imag} */,
  {32'hbf5fa542, 32'h3f37251a} /* (10, 19, 23) {real, imag} */,
  {32'h3fe95f7c, 32'hbf85fd2f} /* (10, 19, 22) {real, imag} */,
  {32'hbebba270, 32'hbf0ac094} /* (10, 19, 21) {real, imag} */,
  {32'hbfcd0031, 32'h405f2328} /* (10, 19, 20) {real, imag} */,
  {32'hc0016706, 32'h404682c8} /* (10, 19, 19) {real, imag} */,
  {32'hc07cd7ef, 32'h3f0fdc42} /* (10, 19, 18) {real, imag} */,
  {32'h3f95dd19, 32'hbff012f6} /* (10, 19, 17) {real, imag} */,
  {32'h40a8ad42, 32'h3fa987d1} /* (10, 19, 16) {real, imag} */,
  {32'h3f568942, 32'h3e20fa44} /* (10, 19, 15) {real, imag} */,
  {32'hc07d195d, 32'hbf17ec48} /* (10, 19, 14) {real, imag} */,
  {32'hc08164f9, 32'h3fb6e704} /* (10, 19, 13) {real, imag} */,
  {32'hbfa84d00, 32'hbf750077} /* (10, 19, 12) {real, imag} */,
  {32'hbf4f9ebc, 32'hc08a8f54} /* (10, 19, 11) {real, imag} */,
  {32'h3fcc1327, 32'hc085b1c9} /* (10, 19, 10) {real, imag} */,
  {32'h3fda0944, 32'hc03be550} /* (10, 19, 9) {real, imag} */,
  {32'hbff7d410, 32'h3fb2680a} /* (10, 19, 8) {real, imag} */,
  {32'hc007c2c1, 32'h40bae044} /* (10, 19, 7) {real, imag} */,
  {32'h40afbd4b, 32'h406ec7ce} /* (10, 19, 6) {real, imag} */,
  {32'h3f5d0048, 32'h40685826} /* (10, 19, 5) {real, imag} */,
  {32'hc038e0a6, 32'hc0073312} /* (10, 19, 4) {real, imag} */,
  {32'hc0508906, 32'hbfdc8e76} /* (10, 19, 3) {real, imag} */,
  {32'h40618776, 32'h402fd7e1} /* (10, 19, 2) {real, imag} */,
  {32'h3f9825cc, 32'h3fccf5db} /* (10, 19, 1) {real, imag} */,
  {32'h3fe544a4, 32'h3ea14bf0} /* (10, 19, 0) {real, imag} */,
  {32'h3f003b14, 32'hbf1064e4} /* (10, 18, 31) {real, imag} */,
  {32'h3f170ad0, 32'hbf082b7c} /* (10, 18, 30) {real, imag} */,
  {32'hbe43971c, 32'hbffeffb8} /* (10, 18, 29) {real, imag} */,
  {32'hbf581560, 32'h3eb182f4} /* (10, 18, 28) {real, imag} */,
  {32'hbfa51884, 32'hbfc8badc} /* (10, 18, 27) {real, imag} */,
  {32'hbe74a438, 32'hc05a5dd8} /* (10, 18, 26) {real, imag} */,
  {32'h40208ca0, 32'hbff139ce} /* (10, 18, 25) {real, imag} */,
  {32'h3f827eb0, 32'hc09ff7c8} /* (10, 18, 24) {real, imag} */,
  {32'hbfd6ac06, 32'hc0867f93} /* (10, 18, 23) {real, imag} */,
  {32'h3f52f3a0, 32'hbffd7526} /* (10, 18, 22) {real, imag} */,
  {32'hbfea83ce, 32'hc0236ac1} /* (10, 18, 21) {real, imag} */,
  {32'hbd85fba0, 32'hbfe4d4b5} /* (10, 18, 20) {real, imag} */,
  {32'h3fcbcd82, 32'hbf9732d4} /* (10, 18, 19) {real, imag} */,
  {32'hc057ab8e, 32'hc048080c} /* (10, 18, 18) {real, imag} */,
  {32'hc067334b, 32'h400aed41} /* (10, 18, 17) {real, imag} */,
  {32'hc00a1dcc, 32'h402658a2} /* (10, 18, 16) {real, imag} */,
  {32'hbf6c1710, 32'h3f163b96} /* (10, 18, 15) {real, imag} */,
  {32'h3fd69eb8, 32'h40348028} /* (10, 18, 14) {real, imag} */,
  {32'h3e7b60e0, 32'h3fd6ff81} /* (10, 18, 13) {real, imag} */,
  {32'hc03dc8fe, 32'h3f3dc7a2} /* (10, 18, 12) {real, imag} */,
  {32'hc05f4ca5, 32'hc08afd62} /* (10, 18, 11) {real, imag} */,
  {32'hc084cc10, 32'hbf346c34} /* (10, 18, 10) {real, imag} */,
  {32'h3e19e6b0, 32'hbe741b28} /* (10, 18, 9) {real, imag} */,
  {32'h3f531928, 32'hc062549a} /* (10, 18, 8) {real, imag} */,
  {32'h3f00ba0d, 32'h3f3ceec4} /* (10, 18, 7) {real, imag} */,
  {32'h3fac9707, 32'h3fb3df4f} /* (10, 18, 6) {real, imag} */,
  {32'hbf99b2e0, 32'hbfd7c01a} /* (10, 18, 5) {real, imag} */,
  {32'hbed3afb8, 32'h3ef163c0} /* (10, 18, 4) {real, imag} */,
  {32'hbf08ba74, 32'h3fd31270} /* (10, 18, 3) {real, imag} */,
  {32'hbfc52da6, 32'hbedad2e0} /* (10, 18, 2) {real, imag} */,
  {32'h40949ed8, 32'h3bc4c600} /* (10, 18, 1) {real, imag} */,
  {32'h40662821, 32'h3f4365fd} /* (10, 18, 0) {real, imag} */,
  {32'hbf58a179, 32'h3e4a82a4} /* (10, 17, 31) {real, imag} */,
  {32'h3f079394, 32'hbf6ab1b8} /* (10, 17, 30) {real, imag} */,
  {32'h404a159d, 32'hbf57ea8c} /* (10, 17, 29) {real, imag} */,
  {32'h406da47c, 32'hbefd0708} /* (10, 17, 28) {real, imag} */,
  {32'hbe51bbf8, 32'hbee0dd58} /* (10, 17, 27) {real, imag} */,
  {32'hc092aa8c, 32'h3e79a2f0} /* (10, 17, 26) {real, imag} */,
  {32'hbf189a04, 32'hbe8535f4} /* (10, 17, 25) {real, imag} */,
  {32'hbd047be0, 32'h4068809a} /* (10, 17, 24) {real, imag} */,
  {32'hbfe4be4a, 32'h4026b491} /* (10, 17, 23) {real, imag} */,
  {32'h3f579f0a, 32'h3fa07354} /* (10, 17, 22) {real, imag} */,
  {32'h40139e7e, 32'h3f3515c8} /* (10, 17, 21) {real, imag} */,
  {32'h3e8378c0, 32'hc0161c7b} /* (10, 17, 20) {real, imag} */,
  {32'hbf623882, 32'hc05cefdb} /* (10, 17, 19) {real, imag} */,
  {32'h3f8dd910, 32'hc04286a0} /* (10, 17, 18) {real, imag} */,
  {32'h400d8fe7, 32'hbff1b7b8} /* (10, 17, 17) {real, imag} */,
  {32'hbfa6575c, 32'hbf9c8958} /* (10, 17, 16) {real, imag} */,
  {32'hbdbbd1e0, 32'h3ebd4810} /* (10, 17, 15) {real, imag} */,
  {32'h4031154c, 32'h3f8875c8} /* (10, 17, 14) {real, imag} */,
  {32'h3e067540, 32'hbed2080c} /* (10, 17, 13) {real, imag} */,
  {32'h3f8a9812, 32'hc02c2d92} /* (10, 17, 12) {real, imag} */,
  {32'h3fce1482, 32'hbfafe464} /* (10, 17, 11) {real, imag} */,
  {32'hbf570b54, 32'h3ff73ff7} /* (10, 17, 10) {real, imag} */,
  {32'h3f61973e, 32'h4027011e} /* (10, 17, 9) {real, imag} */,
  {32'h3dc4bab0, 32'h40289e53} /* (10, 17, 8) {real, imag} */,
  {32'h3f8e29b1, 32'h403f4c1e} /* (10, 17, 7) {real, imag} */,
  {32'h3f9d45e8, 32'h3fe92864} /* (10, 17, 6) {real, imag} */,
  {32'h3fefbd68, 32'hbf163914} /* (10, 17, 5) {real, imag} */,
  {32'h3dbfae90, 32'hbf9e87e0} /* (10, 17, 4) {real, imag} */,
  {32'hc01ed26a, 32'h3f60aa44} /* (10, 17, 3) {real, imag} */,
  {32'hbddaded0, 32'hbfc3abae} /* (10, 17, 2) {real, imag} */,
  {32'hbe33b830, 32'hc0210c71} /* (10, 17, 1) {real, imag} */,
  {32'h3f4c4708, 32'hbf354078} /* (10, 17, 0) {real, imag} */,
  {32'h3fa27a58, 32'hc0114148} /* (10, 16, 31) {real, imag} */,
  {32'h3fc167e3, 32'hc0880e50} /* (10, 16, 30) {real, imag} */,
  {32'h3fd6e30c, 32'hc09f932b} /* (10, 16, 29) {real, imag} */,
  {32'h4048df54, 32'hc0537120} /* (10, 16, 28) {real, imag} */,
  {32'h3e869b20, 32'h3ff60c94} /* (10, 16, 27) {real, imag} */,
  {32'hbf570474, 32'h3e9fdf90} /* (10, 16, 26) {real, imag} */,
  {32'h3dc20fe0, 32'hbf48d922} /* (10, 16, 25) {real, imag} */,
  {32'hbfb20df7, 32'h3fcc9d78} /* (10, 16, 24) {real, imag} */,
  {32'hbf21f410, 32'hbdb81900} /* (10, 16, 23) {real, imag} */,
  {32'h3f8f064c, 32'hbfd327c4} /* (10, 16, 22) {real, imag} */,
  {32'h3fb60d51, 32'hbfea63ec} /* (10, 16, 21) {real, imag} */,
  {32'h4044b690, 32'hbf4a21ec} /* (10, 16, 20) {real, imag} */,
  {32'h3fed1a9c, 32'h3e91eac0} /* (10, 16, 19) {real, imag} */,
  {32'h3f3b8220, 32'hbfba2184} /* (10, 16, 18) {real, imag} */,
  {32'hbfaa6790, 32'hbf49f844} /* (10, 16, 17) {real, imag} */,
  {32'hbe225d88, 32'hbf96b6da} /* (10, 16, 16) {real, imag} */,
  {32'h405b2283, 32'hbf4f6f20} /* (10, 16, 15) {real, imag} */,
  {32'h40419d50, 32'h3fa38f9c} /* (10, 16, 14) {real, imag} */,
  {32'hbf8374e0, 32'h3f85c602} /* (10, 16, 13) {real, imag} */,
  {32'hc085fd46, 32'h3f3285e4} /* (10, 16, 12) {real, imag} */,
  {32'h3f7cf89c, 32'h3f19f8c0} /* (10, 16, 11) {real, imag} */,
  {32'h3f46c24c, 32'h40303b5c} /* (10, 16, 10) {real, imag} */,
  {32'h3e0a34c0, 32'h408942f8} /* (10, 16, 9) {real, imag} */,
  {32'hbfc7243e, 32'h3f3922d8} /* (10, 16, 8) {real, imag} */,
  {32'h3fbd94bc, 32'hbfbf67c9} /* (10, 16, 7) {real, imag} */,
  {32'h3f43d8f0, 32'hbf7e4bc3} /* (10, 16, 6) {real, imag} */,
  {32'hbec059b4, 32'h3f7394ec} /* (10, 16, 5) {real, imag} */,
  {32'hbed7ee50, 32'h4038d757} /* (10, 16, 4) {real, imag} */,
  {32'hbf4b0ff3, 32'h4084400e} /* (10, 16, 3) {real, imag} */,
  {32'h3f9e54e4, 32'h402b056c} /* (10, 16, 2) {real, imag} */,
  {32'h3f8c30c0, 32'h4007ebdc} /* (10, 16, 1) {real, imag} */,
  {32'h3f8dc855, 32'h3fdfc66c} /* (10, 16, 0) {real, imag} */,
  {32'h3f475d41, 32'h3f43ab8f} /* (10, 15, 31) {real, imag} */,
  {32'h3edea868, 32'h3e1aad60} /* (10, 15, 30) {real, imag} */,
  {32'hc009a71b, 32'h3fd8bc56} /* (10, 15, 29) {real, imag} */,
  {32'hc0716320, 32'h3fdaacd6} /* (10, 15, 28) {real, imag} */,
  {32'hbf412d2a, 32'h400ebe81} /* (10, 15, 27) {real, imag} */,
  {32'h3f80e6ca, 32'h3f87774e} /* (10, 15, 26) {real, imag} */,
  {32'hbf5e54cc, 32'h3f80cb11} /* (10, 15, 25) {real, imag} */,
  {32'hc03e0ea0, 32'hbff07fc4} /* (10, 15, 24) {real, imag} */,
  {32'h3f519884, 32'hc00366c1} /* (10, 15, 23) {real, imag} */,
  {32'h3fe74a37, 32'h3fdc248c} /* (10, 15, 22) {real, imag} */,
  {32'hbf5326ae, 32'h3fdeace8} /* (10, 15, 21) {real, imag} */,
  {32'hbf741b60, 32'h3fd72096} /* (10, 15, 20) {real, imag} */,
  {32'hbfe09587, 32'h3f9db052} /* (10, 15, 19) {real, imag} */,
  {32'h404fb6e4, 32'h3e9c4f60} /* (10, 15, 18) {real, imag} */,
  {32'hbf94101e, 32'hbf909ff0} /* (10, 15, 17) {real, imag} */,
  {32'hbf39fe25, 32'h402362d0} /* (10, 15, 16) {real, imag} */,
  {32'h3ed3ed90, 32'h3fdf6314} /* (10, 15, 15) {real, imag} */,
  {32'hbf97657d, 32'hbf6c04cc} /* (10, 15, 14) {real, imag} */,
  {32'h40bdac3d, 32'h3f6557c6} /* (10, 15, 13) {real, imag} */,
  {32'h402900df, 32'h4058b332} /* (10, 15, 12) {real, imag} */,
  {32'hc033cd11, 32'hbe659780} /* (10, 15, 11) {real, imag} */,
  {32'hbfbf7ad2, 32'hbf77fe3e} /* (10, 15, 10) {real, imag} */,
  {32'h3fcdc49d, 32'h4030bf26} /* (10, 15, 9) {real, imag} */,
  {32'h400dfbb0, 32'h403ac6af} /* (10, 15, 8) {real, imag} */,
  {32'hc02ccaa6, 32'h3fa419dd} /* (10, 15, 7) {real, imag} */,
  {32'hc007e2f6, 32'hc00a882d} /* (10, 15, 6) {real, imag} */,
  {32'h3edaa47a, 32'hc010bb43} /* (10, 15, 5) {real, imag} */,
  {32'h403656ec, 32'h3d1c8800} /* (10, 15, 4) {real, imag} */,
  {32'h3f6c912a, 32'h3f492a94} /* (10, 15, 3) {real, imag} */,
  {32'hbf871419, 32'h403ebfb1} /* (10, 15, 2) {real, imag} */,
  {32'h3fb2d982, 32'h40239b3f} /* (10, 15, 1) {real, imag} */,
  {32'h4007856a, 32'h4002b936} /* (10, 15, 0) {real, imag} */,
  {32'hbfd27ae2, 32'h4092198c} /* (10, 14, 31) {real, imag} */,
  {32'hbf909810, 32'h409cf03a} /* (10, 14, 30) {real, imag} */,
  {32'h3fe4cce4, 32'h4002e800} /* (10, 14, 29) {real, imag} */,
  {32'hbfe09728, 32'h3f8f8031} /* (10, 14, 28) {real, imag} */,
  {32'h3f8ee9a4, 32'h3f55678c} /* (10, 14, 27) {real, imag} */,
  {32'hbf42567e, 32'h4002eb14} /* (10, 14, 26) {real, imag} */,
  {32'hc01c3994, 32'h40b23bc8} /* (10, 14, 25) {real, imag} */,
  {32'h3e869562, 32'h40c2c00a} /* (10, 14, 24) {real, imag} */,
  {32'h3ff45b7e, 32'h40341603} /* (10, 14, 23) {real, imag} */,
  {32'h3fcabcb0, 32'hc030bb55} /* (10, 14, 22) {real, imag} */,
  {32'h4034e011, 32'hc00152d5} /* (10, 14, 21) {real, imag} */,
  {32'h3fc644a6, 32'hbf8e2fdb} /* (10, 14, 20) {real, imag} */,
  {32'h3d99d9e0, 32'hc02518d4} /* (10, 14, 19) {real, imag} */,
  {32'hbfcf7a08, 32'hc01bf550} /* (10, 14, 18) {real, imag} */,
  {32'h3e5b72d0, 32'hbfd32346} /* (10, 14, 17) {real, imag} */,
  {32'h40800cb0, 32'h3ec29d60} /* (10, 14, 16) {real, imag} */,
  {32'h3f418300, 32'h3ea3df84} /* (10, 14, 15) {real, imag} */,
  {32'h3f9617b8, 32'h401d963e} /* (10, 14, 14) {real, imag} */,
  {32'h3f1dbef8, 32'h3f78a15e} /* (10, 14, 13) {real, imag} */,
  {32'hc054396a, 32'hbf76ff66} /* (10, 14, 12) {real, imag} */,
  {32'hc0690279, 32'hbf8e0586} /* (10, 14, 11) {real, imag} */,
  {32'hbed50b20, 32'hbffbbe36} /* (10, 14, 10) {real, imag} */,
  {32'hc0078b5b, 32'hbfe6641b} /* (10, 14, 9) {real, imag} */,
  {32'h3ecfb7b0, 32'hbdf2e9c0} /* (10, 14, 8) {real, imag} */,
  {32'hbf6d671d, 32'hbf8a323a} /* (10, 14, 7) {real, imag} */,
  {32'hbe602938, 32'h3da69870} /* (10, 14, 6) {real, imag} */,
  {32'hc0927851, 32'h3f28046b} /* (10, 14, 5) {real, imag} */,
  {32'hc0372571, 32'hc06f7dd4} /* (10, 14, 4) {real, imag} */,
  {32'hc023a69d, 32'h3fec94a0} /* (10, 14, 3) {real, imag} */,
  {32'hc0051589, 32'h408fcf61} /* (10, 14, 2) {real, imag} */,
  {32'hbea9d540, 32'hbf40a8e4} /* (10, 14, 1) {real, imag} */,
  {32'hbf187a3c, 32'hbf0201e3} /* (10, 14, 0) {real, imag} */,
  {32'h402035dd, 32'hc002f503} /* (10, 13, 31) {real, imag} */,
  {32'h3f8b4096, 32'hbf33b6f8} /* (10, 13, 30) {real, imag} */,
  {32'h3eaf8b20, 32'h3f22ad7a} /* (10, 13, 29) {real, imag} */,
  {32'h4062a1d6, 32'hbebd3ed0} /* (10, 13, 28) {real, imag} */,
  {32'h3f9e85f7, 32'h403f01c1} /* (10, 13, 27) {real, imag} */,
  {32'hbeff8e66, 32'h405a2544} /* (10, 13, 26) {real, imag} */,
  {32'hbf2796a8, 32'h40962d2e} /* (10, 13, 25) {real, imag} */,
  {32'hc0647c32, 32'h405517b9} /* (10, 13, 24) {real, imag} */,
  {32'hc00929dc, 32'h3fca1051} /* (10, 13, 23) {real, imag} */,
  {32'hbf983814, 32'h4005739e} /* (10, 13, 22) {real, imag} */,
  {32'hbf93193c, 32'h40839354} /* (10, 13, 21) {real, imag} */,
  {32'hbe90e904, 32'h3fd5c714} /* (10, 13, 20) {real, imag} */,
  {32'h40086eca, 32'h4018f0f2} /* (10, 13, 19) {real, imag} */,
  {32'h3f1376b4, 32'hbf57ee12} /* (10, 13, 18) {real, imag} */,
  {32'h401f348a, 32'h405b3849} /* (10, 13, 17) {real, imag} */,
  {32'hbf9c78f0, 32'h3f54e466} /* (10, 13, 16) {real, imag} */,
  {32'hbfed5d97, 32'h3cfdf420} /* (10, 13, 15) {real, imag} */,
  {32'h401ab059, 32'h408830ad} /* (10, 13, 14) {real, imag} */,
  {32'h405102b6, 32'h406af39a} /* (10, 13, 13) {real, imag} */,
  {32'h3eb83c80, 32'h3f7b2d95} /* (10, 13, 12) {real, imag} */,
  {32'hbfc7cc5a, 32'h405a5079} /* (10, 13, 11) {real, imag} */,
  {32'hbf0b8e7e, 32'hbea36494} /* (10, 13, 10) {real, imag} */,
  {32'hc05cacda, 32'h3dc39e20} /* (10, 13, 9) {real, imag} */,
  {32'hbfc9b668, 32'hc0451905} /* (10, 13, 8) {real, imag} */,
  {32'h3f531e3c, 32'hbf7956f0} /* (10, 13, 7) {real, imag} */,
  {32'h40935df5, 32'hbd0f63e0} /* (10, 13, 6) {real, imag} */,
  {32'h40279b2a, 32'h3f86910d} /* (10, 13, 5) {real, imag} */,
  {32'h3ec1d370, 32'h3ebd2850} /* (10, 13, 4) {real, imag} */,
  {32'h3faba9b0, 32'h3f374e14} /* (10, 13, 3) {real, imag} */,
  {32'hc05c8fd8, 32'hbee91778} /* (10, 13, 2) {real, imag} */,
  {32'h3f8dda9c, 32'h3ed8f534} /* (10, 13, 1) {real, imag} */,
  {32'h40264eb6, 32'h3fc53e26} /* (10, 13, 0) {real, imag} */,
  {32'hbf65e72e, 32'h3ee31c30} /* (10, 12, 31) {real, imag} */,
  {32'hbf138d02, 32'h40c05ee6} /* (10, 12, 30) {real, imag} */,
  {32'hbf284b92, 32'h40632322} /* (10, 12, 29) {real, imag} */,
  {32'hc0303b2d, 32'hc0931938} /* (10, 12, 28) {real, imag} */,
  {32'hc080f176, 32'hc0c1389e} /* (10, 12, 27) {real, imag} */,
  {32'hc13aabfe, 32'h3fe87660} /* (10, 12, 26) {real, imag} */,
  {32'hc0979d98, 32'h40341dee} /* (10, 12, 25) {real, imag} */,
  {32'hc09f29f4, 32'h3da906d0} /* (10, 12, 24) {real, imag} */,
  {32'hc0847a6c, 32'hc047579f} /* (10, 12, 23) {real, imag} */,
  {32'hc0171f2c, 32'hbfb822a8} /* (10, 12, 22) {real, imag} */,
  {32'hbf17c260, 32'h4034df5d} /* (10, 12, 21) {real, imag} */,
  {32'hc0aa9d54, 32'h3f18d227} /* (10, 12, 20) {real, imag} */,
  {32'hc0653195, 32'h40479c4c} /* (10, 12, 19) {real, imag} */,
  {32'hbfc6499f, 32'h3fc546ac} /* (10, 12, 18) {real, imag} */,
  {32'h3c843d00, 32'hc0214c2e} /* (10, 12, 17) {real, imag} */,
  {32'h3f6f2192, 32'hc0841709} /* (10, 12, 16) {real, imag} */,
  {32'h408bdf85, 32'hbfa3f789} /* (10, 12, 15) {real, imag} */,
  {32'h3ffa706c, 32'h404e2610} /* (10, 12, 14) {real, imag} */,
  {32'hc0855e98, 32'h3fefae60} /* (10, 12, 13) {real, imag} */,
  {32'hc08927f8, 32'hc0073c7b} /* (10, 12, 12) {real, imag} */,
  {32'hbfd46a5d, 32'h3f1c2958} /* (10, 12, 11) {real, imag} */,
  {32'h40512a60, 32'h400dab07} /* (10, 12, 10) {real, imag} */,
  {32'h400a3b14, 32'hc0086fea} /* (10, 12, 9) {real, imag} */,
  {32'hbfdcc20d, 32'hc09adf36} /* (10, 12, 8) {real, imag} */,
  {32'hc00eb81e, 32'h402bf2bf} /* (10, 12, 7) {real, imag} */,
  {32'hc039a38a, 32'h40e8025a} /* (10, 12, 6) {real, imag} */,
  {32'hbf721ea4, 32'h3f0c0180} /* (10, 12, 5) {real, imag} */,
  {32'hbe2c4c28, 32'hc030ad9b} /* (10, 12, 4) {real, imag} */,
  {32'h4059dad3, 32'hc096e2e0} /* (10, 12, 3) {real, imag} */,
  {32'h40847b77, 32'hc085b536} /* (10, 12, 2) {real, imag} */,
  {32'h3ed2c6d8, 32'h3fce1c98} /* (10, 12, 1) {real, imag} */,
  {32'h3f996dbc, 32'h3fa04221} /* (10, 12, 0) {real, imag} */,
  {32'hbeb0555c, 32'hc019b828} /* (10, 11, 31) {real, imag} */,
  {32'h4084b20a, 32'hbfdefef9} /* (10, 11, 30) {real, imag} */,
  {32'h404fc387, 32'h40856e3c} /* (10, 11, 29) {real, imag} */,
  {32'h40814734, 32'h4092ae16} /* (10, 11, 28) {real, imag} */,
  {32'h3f7f4bc0, 32'hbfc20710} /* (10, 11, 27) {real, imag} */,
  {32'hc084b48a, 32'hc0927aba} /* (10, 11, 26) {real, imag} */,
  {32'hc0b646b3, 32'hbfb5577a} /* (10, 11, 25) {real, imag} */,
  {32'h3f675b38, 32'hc0448fa6} /* (10, 11, 24) {real, imag} */,
  {32'h40561c3a, 32'hbeee1924} /* (10, 11, 23) {real, imag} */,
  {32'hbe1de240, 32'h3ec3e588} /* (10, 11, 22) {real, imag} */,
  {32'hc0a3911f, 32'h4105d556} /* (10, 11, 21) {real, imag} */,
  {32'hc070d050, 32'h412a1e00} /* (10, 11, 20) {real, imag} */,
  {32'hbf51f5d0, 32'h4084ca4d} /* (10, 11, 19) {real, imag} */,
  {32'hc050f386, 32'hc01b88c4} /* (10, 11, 18) {real, imag} */,
  {32'hbf2c0bd2, 32'h3e348c88} /* (10, 11, 17) {real, imag} */,
  {32'hc0588f08, 32'h3fdb22fd} /* (10, 11, 16) {real, imag} */,
  {32'hbfc2613c, 32'hc02500e9} /* (10, 11, 15) {real, imag} */,
  {32'h3f042a84, 32'hc0656618} /* (10, 11, 14) {real, imag} */,
  {32'h405b56ab, 32'h405635fe} /* (10, 11, 13) {real, imag} */,
  {32'h403761eb, 32'h40bcfe45} /* (10, 11, 12) {real, imag} */,
  {32'h409d833f, 32'h40018352} /* (10, 11, 11) {real, imag} */,
  {32'h3fa8e39d, 32'hc019a5a6} /* (10, 11, 10) {real, imag} */,
  {32'hc106f860, 32'h3f9e5abe} /* (10, 11, 9) {real, imag} */,
  {32'hc094565a, 32'h40b7d25c} /* (10, 11, 8) {real, imag} */,
  {32'hbff7366c, 32'h4104f327} /* (10, 11, 7) {real, imag} */,
  {32'hbfe41b4e, 32'h3f03dda0} /* (10, 11, 6) {real, imag} */,
  {32'h40b5a131, 32'hbff00a9a} /* (10, 11, 5) {real, imag} */,
  {32'hc040b063, 32'h3f6e3b10} /* (10, 11, 4) {real, imag} */,
  {32'hc0c66d33, 32'hc0b90ed8} /* (10, 11, 3) {real, imag} */,
  {32'h3f1be60f, 32'hc1474d78} /* (10, 11, 2) {real, imag} */,
  {32'hc04b5a77, 32'hc0b7ceee} /* (10, 11, 1) {real, imag} */,
  {32'hc0edb373, 32'hbee3054c} /* (10, 11, 0) {real, imag} */,
  {32'h3e8c23cc, 32'h402a644c} /* (10, 10, 31) {real, imag} */,
  {32'h3fe3ec3b, 32'hc0014ca3} /* (10, 10, 30) {real, imag} */,
  {32'hbf9b49c0, 32'hc05f3cfa} /* (10, 10, 29) {real, imag} */,
  {32'hc0741ed6, 32'h404ec0a5} /* (10, 10, 28) {real, imag} */,
  {32'h3fc83ebc, 32'h3fe3a8e2} /* (10, 10, 27) {real, imag} */,
  {32'hbeef1884, 32'hc05eebdc} /* (10, 10, 26) {real, imag} */,
  {32'hc061fecd, 32'hc06bc657} /* (10, 10, 25) {real, imag} */,
  {32'hbfee2796, 32'hbf9883f2} /* (10, 10, 24) {real, imag} */,
  {32'hc08d10c2, 32'h408103a2} /* (10, 10, 23) {real, imag} */,
  {32'hc130b541, 32'h404eb213} /* (10, 10, 22) {real, imag} */,
  {32'hbfb6fade, 32'h3f35ac04} /* (10, 10, 21) {real, imag} */,
  {32'h408dfd92, 32'h3ea9b100} /* (10, 10, 20) {real, imag} */,
  {32'hbf113018, 32'hc00bddd2} /* (10, 10, 19) {real, imag} */,
  {32'hc01750b9, 32'hc037ff1c} /* (10, 10, 18) {real, imag} */,
  {32'hc0006be9, 32'hbeacd950} /* (10, 10, 17) {real, imag} */,
  {32'hc0ecbbc6, 32'h407c309b} /* (10, 10, 16) {real, imag} */,
  {32'hc017d678, 32'hc074e7c7} /* (10, 10, 15) {real, imag} */,
  {32'hc09d2513, 32'hc08ee7a7} /* (10, 10, 14) {real, imag} */,
  {32'hc0847c80, 32'h3f52d27f} /* (10, 10, 13) {real, imag} */,
  {32'h3c005900, 32'h40ab0c89} /* (10, 10, 12) {real, imag} */,
  {32'h40be252e, 32'h3f8ecae7} /* (10, 10, 11) {real, imag} */,
  {32'h40745d9f, 32'h3ff14ca2} /* (10, 10, 10) {real, imag} */,
  {32'hbf23083e, 32'h404a426d} /* (10, 10, 9) {real, imag} */,
  {32'hc025b6bc, 32'hc09ec1c8} /* (10, 10, 8) {real, imag} */,
  {32'hc0970830, 32'h40174b62} /* (10, 10, 7) {real, imag} */,
  {32'hc03484b9, 32'h3fe92a40} /* (10, 10, 6) {real, imag} */,
  {32'h3f858a6d, 32'h3f6141a8} /* (10, 10, 5) {real, imag} */,
  {32'h40b5adce, 32'hbf287ca0} /* (10, 10, 4) {real, imag} */,
  {32'h4110adab, 32'h3ff6b2b2} /* (10, 10, 3) {real, imag} */,
  {32'h40841d6a, 32'h3fe9bee4} /* (10, 10, 2) {real, imag} */,
  {32'h40622649, 32'hc09ecec6} /* (10, 10, 1) {real, imag} */,
  {32'h40b796f8, 32'hc00a603c} /* (10, 10, 0) {real, imag} */,
  {32'h404217b8, 32'h3ee88bbe} /* (10, 9, 31) {real, imag} */,
  {32'hbf9bf9fe, 32'h401c6a89} /* (10, 9, 30) {real, imag} */,
  {32'hc051d1fa, 32'hbe11fde0} /* (10, 9, 29) {real, imag} */,
  {32'h3f85f5cc, 32'hc020a782} /* (10, 9, 28) {real, imag} */,
  {32'h4055040d, 32'hc0edea39} /* (10, 9, 27) {real, imag} */,
  {32'h40938b57, 32'hc0b333e8} /* (10, 9, 26) {real, imag} */,
  {32'hc020adf1, 32'h3fedef61} /* (10, 9, 25) {real, imag} */,
  {32'h4028c792, 32'h4059b9a8} /* (10, 9, 24) {real, imag} */,
  {32'h4090ed52, 32'hc06a3da3} /* (10, 9, 23) {real, imag} */,
  {32'hbd508320, 32'hc0010f8e} /* (10, 9, 22) {real, imag} */,
  {32'h3fe56753, 32'hc08b354a} /* (10, 9, 21) {real, imag} */,
  {32'h402059a4, 32'hc03a9b73} /* (10, 9, 20) {real, imag} */,
  {32'hc01f1563, 32'h405a9698} /* (10, 9, 19) {real, imag} */,
  {32'hc09c219e, 32'h407ddb4e} /* (10, 9, 18) {real, imag} */,
  {32'hbf871589, 32'h3dbb2940} /* (10, 9, 17) {real, imag} */,
  {32'hbfc15306, 32'hc0cb113e} /* (10, 9, 16) {real, imag} */,
  {32'hc052ed36, 32'hc0bbde31} /* (10, 9, 15) {real, imag} */,
  {32'h3f963ff8, 32'h3fa919ae} /* (10, 9, 14) {real, imag} */,
  {32'h40cc26cc, 32'hbf8e3eb4} /* (10, 9, 13) {real, imag} */,
  {32'h400438cc, 32'hc0817f92} /* (10, 9, 12) {real, imag} */,
  {32'h3f85601a, 32'hc09f37dd} /* (10, 9, 11) {real, imag} */,
  {32'h3f47e9c4, 32'hc081db97} /* (10, 9, 10) {real, imag} */,
  {32'h4046e6a9, 32'hc0c4f8e4} /* (10, 9, 9) {real, imag} */,
  {32'h408ddfb2, 32'hc10850f4} /* (10, 9, 8) {real, imag} */,
  {32'h3e494fc0, 32'hc0b0f20a} /* (10, 9, 7) {real, imag} */,
  {32'hc0f31dad, 32'hc0ebbf82} /* (10, 9, 6) {real, imag} */,
  {32'hc0b36cca, 32'hc0c11c66} /* (10, 9, 5) {real, imag} */,
  {32'h400de5b8, 32'h3fb5f54e} /* (10, 9, 4) {real, imag} */,
  {32'hc0a715bd, 32'hbfcd7cfc} /* (10, 9, 3) {real, imag} */,
  {32'hc1025543, 32'h3fc1e938} /* (10, 9, 2) {real, imag} */,
  {32'h3fb9f0fd, 32'h41359e54} /* (10, 9, 1) {real, imag} */,
  {32'h40188fa3, 32'h4125b7d1} /* (10, 9, 0) {real, imag} */,
  {32'h3fd07150, 32'hc10c4188} /* (10, 8, 31) {real, imag} */,
  {32'h3f8e2125, 32'hc0ea4bad} /* (10, 8, 30) {real, imag} */,
  {32'hc091b803, 32'h3f8a4252} /* (10, 8, 29) {real, imag} */,
  {32'hc02ebad4, 32'h40c17309} /* (10, 8, 28) {real, imag} */,
  {32'h3ff77e18, 32'h403e2b4e} /* (10, 8, 27) {real, imag} */,
  {32'h40304b60, 32'hc09d62f6} /* (10, 8, 26) {real, imag} */,
  {32'h4029c7e5, 32'hc05c82d0} /* (10, 8, 25) {real, imag} */,
  {32'h408e168c, 32'h41431790} /* (10, 8, 24) {real, imag} */,
  {32'h4133b690, 32'h40b473fa} /* (10, 8, 23) {real, imag} */,
  {32'h40cd68ee, 32'hc09715ed} /* (10, 8, 22) {real, imag} */,
  {32'h40ea0241, 32'hc0e074ba} /* (10, 8, 21) {real, imag} */,
  {32'h412a7a7b, 32'hc0c17c5a} /* (10, 8, 20) {real, imag} */,
  {32'h40b220d5, 32'hc0be22c8} /* (10, 8, 19) {real, imag} */,
  {32'hbfedcbf0, 32'hc0917555} /* (10, 8, 18) {real, imag} */,
  {32'hc0c689bd, 32'hc0480d2c} /* (10, 8, 17) {real, imag} */,
  {32'hc0626405, 32'h3fcbf757} /* (10, 8, 16) {real, imag} */,
  {32'h40c3cc34, 32'h3ea58c18} /* (10, 8, 15) {real, imag} */,
  {32'h40f69a3a, 32'hc0830ad8} /* (10, 8, 14) {real, imag} */,
  {32'hbd8089f8, 32'hbfedceee} /* (10, 8, 13) {real, imag} */,
  {32'h40f27e77, 32'h400f53fd} /* (10, 8, 12) {real, imag} */,
  {32'hc02f04e0, 32'h40837fc4} /* (10, 8, 11) {real, imag} */,
  {32'hc02b731c, 32'h40089250} /* (10, 8, 10) {real, imag} */,
  {32'h4035e6f4, 32'hc0f73a08} /* (10, 8, 9) {real, imag} */,
  {32'h402985c2, 32'hc0bc978e} /* (10, 8, 8) {real, imag} */,
  {32'h40d06518, 32'hc084a931} /* (10, 8, 7) {real, imag} */,
  {32'h40e430ad, 32'h3f2335d0} /* (10, 8, 6) {real, imag} */,
  {32'h40bebcf5, 32'hc02025fe} /* (10, 8, 5) {real, imag} */,
  {32'h40ddd0ae, 32'hc06304e7} /* (10, 8, 4) {real, imag} */,
  {32'hbf7886a9, 32'h3fea1389} /* (10, 8, 3) {real, imag} */,
  {32'h3e2e0610, 32'h409d3f28} /* (10, 8, 2) {real, imag} */,
  {32'hbf5a27f8, 32'h40ef803b} /* (10, 8, 1) {real, imag} */,
  {32'h4000f882, 32'h3f84f3aa} /* (10, 8, 0) {real, imag} */,
  {32'hc0205c92, 32'h40992508} /* (10, 7, 31) {real, imag} */,
  {32'hc171b854, 32'h410ee91c} /* (10, 7, 30) {real, imag} */,
  {32'hc146e451, 32'hc0d352f6} /* (10, 7, 29) {real, imag} */,
  {32'hc0b4e83b, 32'hc100a920} /* (10, 7, 28) {real, imag} */,
  {32'h3f9e6f58, 32'hbff765b4} /* (10, 7, 27) {real, imag} */,
  {32'h3fd68fec, 32'hc056b33d} /* (10, 7, 26) {real, imag} */,
  {32'hc09be4f4, 32'hc0692f2f} /* (10, 7, 25) {real, imag} */,
  {32'hc0b7c730, 32'hc0033eba} /* (10, 7, 24) {real, imag} */,
  {32'hbfe019ab, 32'h40495633} /* (10, 7, 23) {real, imag} */,
  {32'h3f0d1df8, 32'hc01bb12c} /* (10, 7, 22) {real, imag} */,
  {32'hbf751364, 32'hbf289013} /* (10, 7, 21) {real, imag} */,
  {32'h40467958, 32'hc115fd62} /* (10, 7, 20) {real, imag} */,
  {32'h40383532, 32'hc04e2199} /* (10, 7, 19) {real, imag} */,
  {32'h40e95b66, 32'hbf5e5678} /* (10, 7, 18) {real, imag} */,
  {32'h40df809d, 32'hc08708d9} /* (10, 7, 17) {real, imag} */,
  {32'h3ed96f68, 32'hc0e889cc} /* (10, 7, 16) {real, imag} */,
  {32'h3ffbe72a, 32'h3fe8a637} /* (10, 7, 15) {real, imag} */,
  {32'h40884ea0, 32'hbf2ec904} /* (10, 7, 14) {real, imag} */,
  {32'hc0bdee04, 32'h40e8d56f} /* (10, 7, 13) {real, imag} */,
  {32'hc067fa32, 32'h402359fb} /* (10, 7, 12) {real, imag} */,
  {32'h3f204488, 32'h3ffa61b0} /* (10, 7, 11) {real, imag} */,
  {32'h3f692d6c, 32'hc066dc12} /* (10, 7, 10) {real, imag} */,
  {32'h4048422b, 32'h3fa65dc0} /* (10, 7, 9) {real, imag} */,
  {32'h4137c17a, 32'h4081a5b3} /* (10, 7, 8) {real, imag} */,
  {32'h418b646e, 32'hbfcc9c20} /* (10, 7, 7) {real, imag} */,
  {32'h4084738b, 32'hbe96d8a8} /* (10, 7, 6) {real, imag} */,
  {32'h40a86d2a, 32'hc024129d} /* (10, 7, 5) {real, imag} */,
  {32'h408bf24c, 32'hc0c630ae} /* (10, 7, 4) {real, imag} */,
  {32'h40b2ae4b, 32'hc00e3a4a} /* (10, 7, 3) {real, imag} */,
  {32'h40d88b7b, 32'h401288c0} /* (10, 7, 2) {real, imag} */,
  {32'h40be01e9, 32'hc063263e} /* (10, 7, 1) {real, imag} */,
  {32'h408d2c6e, 32'hc12b0399} /* (10, 7, 0) {real, imag} */,
  {32'h3f548c46, 32'hbf28b0a4} /* (10, 6, 31) {real, imag} */,
  {32'hc07c90f8, 32'hbe9811f8} /* (10, 6, 30) {real, imag} */,
  {32'h3f0fcbd0, 32'h40a0a1aa} /* (10, 6, 29) {real, imag} */,
  {32'hbfa20c54, 32'h3ffa1a82} /* (10, 6, 28) {real, imag} */,
  {32'h40498430, 32'hc0a978cc} /* (10, 6, 27) {real, imag} */,
  {32'hc0673d32, 32'hc0084a7e} /* (10, 6, 26) {real, imag} */,
  {32'h40b0bf8e, 32'h40458556} /* (10, 6, 25) {real, imag} */,
  {32'h412a44cb, 32'h41021266} /* (10, 6, 24) {real, imag} */,
  {32'h4113657f, 32'h40a5a0bc} /* (10, 6, 23) {real, imag} */,
  {32'hc0b50c56, 32'hbeb0a4b8} /* (10, 6, 22) {real, imag} */,
  {32'hc0277cac, 32'h40284b1d} /* (10, 6, 21) {real, imag} */,
  {32'h40da7814, 32'hc0e43099} /* (10, 6, 20) {real, imag} */,
  {32'hc0e53a84, 32'hc1941cc2} /* (10, 6, 19) {real, imag} */,
  {32'hc04c7eb7, 32'hc18e921d} /* (10, 6, 18) {real, imag} */,
  {32'h3f0aad68, 32'hc03286a5} /* (10, 6, 17) {real, imag} */,
  {32'hbf8e326e, 32'h4092e514} /* (10, 6, 16) {real, imag} */,
  {32'hc0b942fa, 32'h400fabb5} /* (10, 6, 15) {real, imag} */,
  {32'hc0d3b666, 32'hc038e9c6} /* (10, 6, 14) {real, imag} */,
  {32'hc13fc0f8, 32'h40cb6c1f} /* (10, 6, 13) {real, imag} */,
  {32'hc1a28f47, 32'h40a57d6a} /* (10, 6, 12) {real, imag} */,
  {32'hc0899bb6, 32'hbfec0cd9} /* (10, 6, 11) {real, imag} */,
  {32'hc0716bf8, 32'hbe6c2ff0} /* (10, 6, 10) {real, imag} */,
  {32'hc0fc7ac2, 32'hbfdfac57} /* (10, 6, 9) {real, imag} */,
  {32'h408d1cc8, 32'hc0f9905e} /* (10, 6, 8) {real, imag} */,
  {32'hbf2b14e8, 32'hc135b8d2} /* (10, 6, 7) {real, imag} */,
  {32'hc086e62a, 32'h3e9695c8} /* (10, 6, 6) {real, imag} */,
  {32'h40662820, 32'hc011d808} /* (10, 6, 5) {real, imag} */,
  {32'h401da1d0, 32'hc06a2942} /* (10, 6, 4) {real, imag} */,
  {32'hc0a287e0, 32'h404aea32} /* (10, 6, 3) {real, imag} */,
  {32'hc10b31f8, 32'h406ae030} /* (10, 6, 2) {real, imag} */,
  {32'hc07940c8, 32'hc04e875f} /* (10, 6, 1) {real, imag} */,
  {32'hbfd8ab56, 32'h3f971dd7} /* (10, 6, 0) {real, imag} */,
  {32'h3f95a257, 32'hc0b23c62} /* (10, 5, 31) {real, imag} */,
  {32'h40d03cb4, 32'hc1164678} /* (10, 5, 30) {real, imag} */,
  {32'h40a944a5, 32'hc04e938b} /* (10, 5, 29) {real, imag} */,
  {32'h3e5aeb30, 32'hc0cbc130} /* (10, 5, 28) {real, imag} */,
  {32'h405728bb, 32'hc0fbcf90} /* (10, 5, 27) {real, imag} */,
  {32'h405dbb8d, 32'h4040799d} /* (10, 5, 26) {real, imag} */,
  {32'h402a2064, 32'hc0987f52} /* (10, 5, 25) {real, imag} */,
  {32'h4110b616, 32'hc17031ba} /* (10, 5, 24) {real, imag} */,
  {32'h41bacc41, 32'hc15db524} /* (10, 5, 23) {real, imag} */,
  {32'h4162367c, 32'hc112d4b5} /* (10, 5, 22) {real, imag} */,
  {32'h4116be49, 32'h3e28cc20} /* (10, 5, 21) {real, imag} */,
  {32'h409f28c4, 32'hbf991e0d} /* (10, 5, 20) {real, imag} */,
  {32'h404d2da7, 32'h40b88dea} /* (10, 5, 19) {real, imag} */,
  {32'h40d6a0d4, 32'hc09721a3} /* (10, 5, 18) {real, imag} */,
  {32'h411d870d, 32'hc0162db9} /* (10, 5, 17) {real, imag} */,
  {32'hbe8fc588, 32'hbebfcd2c} /* (10, 5, 16) {real, imag} */,
  {32'hc0c6e68a, 32'h3f73f56c} /* (10, 5, 15) {real, imag} */,
  {32'h401530ba, 32'h4004a698} /* (10, 5, 14) {real, imag} */,
  {32'hc10571a8, 32'hc0d72a13} /* (10, 5, 13) {real, imag} */,
  {32'hc16b5180, 32'hc06f41f8} /* (10, 5, 12) {real, imag} */,
  {32'h4033ea3a, 32'h40a9a33b} /* (10, 5, 11) {real, imag} */,
  {32'h3eb23ef4, 32'h4111b1c8} /* (10, 5, 10) {real, imag} */,
  {32'hc065c16a, 32'hbf25f4a8} /* (10, 5, 9) {real, imag} */,
  {32'hc0535cbb, 32'hc0dc147e} /* (10, 5, 8) {real, imag} */,
  {32'hc11edf54, 32'hc1016a60} /* (10, 5, 7) {real, imag} */,
  {32'hc1453e86, 32'h40df9967} /* (10, 5, 6) {real, imag} */,
  {32'hbf3911ea, 32'h40892824} /* (10, 5, 5) {real, imag} */,
  {32'h40da98e2, 32'h3eb26d20} /* (10, 5, 4) {real, imag} */,
  {32'h3efd3b30, 32'hc0358cb1} /* (10, 5, 3) {real, imag} */,
  {32'hbee6afb0, 32'hc0a76a5c} /* (10, 5, 2) {real, imag} */,
  {32'h40807cc5, 32'hbf3f08ec} /* (10, 5, 1) {real, imag} */,
  {32'h3f881f3c, 32'hc020ddcd} /* (10, 5, 0) {real, imag} */,
  {32'hbff7c85e, 32'h40b841be} /* (10, 4, 31) {real, imag} */,
  {32'hc0cb7c06, 32'h413e1e04} /* (10, 4, 30) {real, imag} */,
  {32'hc07bc6a4, 32'hc0c17289} /* (10, 4, 29) {real, imag} */,
  {32'hc0386dc9, 32'hc183b096} /* (10, 4, 28) {real, imag} */,
  {32'hbfa8adcf, 32'hc0389382} /* (10, 4, 27) {real, imag} */,
  {32'hc0c4d8ce, 32'hbf2e0818} /* (10, 4, 26) {real, imag} */,
  {32'hc01eeb04, 32'hc12f1355} /* (10, 4, 25) {real, imag} */,
  {32'hc0e2b042, 32'hc137b368} /* (10, 4, 24) {real, imag} */,
  {32'hc17b60b4, 32'h412acd60} /* (10, 4, 23) {real, imag} */,
  {32'hc1802174, 32'h413b71e4} /* (10, 4, 22) {real, imag} */,
  {32'hc1afd708, 32'h415f8f85} /* (10, 4, 21) {real, imag} */,
  {32'hc15e31f0, 32'h3f6fb5d9} /* (10, 4, 20) {real, imag} */,
  {32'h3fdf964a, 32'h3e47ccb0} /* (10, 4, 19) {real, imag} */,
  {32'h3f9d79a0, 32'h3ebf4b90} /* (10, 4, 18) {real, imag} */,
  {32'h40127ca6, 32'hbf9958ad} /* (10, 4, 17) {real, imag} */,
  {32'h41345b5e, 32'h4082997e} /* (10, 4, 16) {real, imag} */,
  {32'h41558dd0, 32'hc0d014e2} /* (10, 4, 15) {real, imag} */,
  {32'h40e694d3, 32'h40c8a511} /* (10, 4, 14) {real, imag} */,
  {32'hc0c6d2ba, 32'h411714a0} /* (10, 4, 13) {real, imag} */,
  {32'hbe8bf0c0, 32'h40a9a03a} /* (10, 4, 12) {real, imag} */,
  {32'hc0eff002, 32'h4112e1d4} /* (10, 4, 11) {real, imag} */,
  {32'hc0f42d0a, 32'hc0738744} /* (10, 4, 10) {real, imag} */,
  {32'hc00f1dac, 32'hc053fcb4} /* (10, 4, 9) {real, imag} */,
  {32'hbf48d412, 32'hc08ce65a} /* (10, 4, 8) {real, imag} */,
  {32'h40978157, 32'hc1269512} /* (10, 4, 7) {real, imag} */,
  {32'hbf87d14d, 32'hc08318f2} /* (10, 4, 6) {real, imag} */,
  {32'hc0def4fb, 32'hc06b0866} /* (10, 4, 5) {real, imag} */,
  {32'hc11f7ea4, 32'hc0e42a70} /* (10, 4, 4) {real, imag} */,
  {32'h3f1f622c, 32'hc1160be2} /* (10, 4, 3) {real, imag} */,
  {32'h417ce4e4, 32'hbf44c5a5} /* (10, 4, 2) {real, imag} */,
  {32'h3fee5760, 32'hc0bc4994} /* (10, 4, 1) {real, imag} */,
  {32'hc0dfb17f, 32'hc0ce538c} /* (10, 4, 0) {real, imag} */,
  {32'h3d815400, 32'h3fdd45e0} /* (10, 3, 31) {real, imag} */,
  {32'h4103f7ad, 32'h40c72f4a} /* (10, 3, 30) {real, imag} */,
  {32'h40930616, 32'h4101c1e6} /* (10, 3, 29) {real, imag} */,
  {32'h409669b6, 32'h41280551} /* (10, 3, 28) {real, imag} */,
  {32'hc03b4eb6, 32'h413f0762} /* (10, 3, 27) {real, imag} */,
  {32'hc092d474, 32'hbf8900a6} /* (10, 3, 26) {real, imag} */,
  {32'hbf4982f8, 32'h40346ef2} /* (10, 3, 25) {real, imag} */,
  {32'hc0a8acea, 32'hbf86e87a} /* (10, 3, 24) {real, imag} */,
  {32'hc1143d8d, 32'hc0ba0d8a} /* (10, 3, 23) {real, imag} */,
  {32'hc178a385, 32'hc0885d41} /* (10, 3, 22) {real, imag} */,
  {32'hc13c5f7a, 32'hc12a065b} /* (10, 3, 21) {real, imag} */,
  {32'hc0cc127c, 32'hc116ae33} /* (10, 3, 20) {real, imag} */,
  {32'hbfd78a7d, 32'hc012f24c} /* (10, 3, 19) {real, imag} */,
  {32'h41352002, 32'hbf391420} /* (10, 3, 18) {real, imag} */,
  {32'h41199442, 32'h40d73da8} /* (10, 3, 17) {real, imag} */,
  {32'h4038128e, 32'h40fb4d9c} /* (10, 3, 16) {real, imag} */,
  {32'h3f3c1038, 32'hc01fd294} /* (10, 3, 15) {real, imag} */,
  {32'hc0a6bae2, 32'hc0c99307} /* (10, 3, 14) {real, imag} */,
  {32'h404312da, 32'hc10ff0bb} /* (10, 3, 13) {real, imag} */,
  {32'h41384d60, 32'hc0651408} /* (10, 3, 12) {real, imag} */,
  {32'hc090f0b3, 32'hbfac5900} /* (10, 3, 11) {real, imag} */,
  {32'hc1724978, 32'hc105ebc0} /* (10, 3, 10) {real, imag} */,
  {32'hc0a309b2, 32'hc09e323e} /* (10, 3, 9) {real, imag} */,
  {32'hc063efd6, 32'hc0a2a4fa} /* (10, 3, 8) {real, imag} */,
  {32'hc1342c96, 32'h406c5a0e} /* (10, 3, 7) {real, imag} */,
  {32'hc0f39023, 32'hbfa2d473} /* (10, 3, 6) {real, imag} */,
  {32'h3f505230, 32'h3ffbf504} /* (10, 3, 5) {real, imag} */,
  {32'hc057f5e2, 32'h40ce147b} /* (10, 3, 4) {real, imag} */,
  {32'hc0a2ac27, 32'h4042b08d} /* (10, 3, 3) {real, imag} */,
  {32'h4036af7a, 32'hbfd035d4} /* (10, 3, 2) {real, imag} */,
  {32'h41b2b66f, 32'hc004483a} /* (10, 3, 1) {real, imag} */,
  {32'h4127e8dd, 32'h3f295518} /* (10, 3, 0) {real, imag} */,
  {32'h3fe60cca, 32'hc051e272} /* (10, 2, 31) {real, imag} */,
  {32'h3fa358b0, 32'h3faa25c8} /* (10, 2, 30) {real, imag} */,
  {32'h40c2d259, 32'h4005f728} /* (10, 2, 29) {real, imag} */,
  {32'h414e7734, 32'h408eb94b} /* (10, 2, 28) {real, imag} */,
  {32'h415bb433, 32'h40c24a30} /* (10, 2, 27) {real, imag} */,
  {32'h4141e48b, 32'hc107520c} /* (10, 2, 26) {real, imag} */,
  {32'hbfc25d93, 32'hc03c58ec} /* (10, 2, 25) {real, imag} */,
  {32'h4104fdfc, 32'h408ff359} /* (10, 2, 24) {real, imag} */,
  {32'h413392f9, 32'h3fdd8543} /* (10, 2, 23) {real, imag} */,
  {32'h3d7e1c00, 32'h410aae0a} /* (10, 2, 22) {real, imag} */,
  {32'hc162c18f, 32'hc13cecee} /* (10, 2, 21) {real, imag} */,
  {32'h3e865908, 32'h40f53ec8} /* (10, 2, 20) {real, imag} */,
  {32'hbfeb2a40, 32'h411c8e07} /* (10, 2, 19) {real, imag} */,
  {32'hc12767e3, 32'h3ffb0a18} /* (10, 2, 18) {real, imag} */,
  {32'hc124975c, 32'hc14dc3e6} /* (10, 2, 17) {real, imag} */,
  {32'h3f6fec1e, 32'hbf24bde0} /* (10, 2, 16) {real, imag} */,
  {32'hc0afd22c, 32'h408637c7} /* (10, 2, 15) {real, imag} */,
  {32'hc196be32, 32'hc11bb610} /* (10, 2, 14) {real, imag} */,
  {32'hc19b1eea, 32'h3fee88f4} /* (10, 2, 13) {real, imag} */,
  {32'hc11cc00a, 32'h40937385} /* (10, 2, 12) {real, imag} */,
  {32'hc0200fe7, 32'h4028e213} /* (10, 2, 11) {real, imag} */,
  {32'h40dbbd05, 32'hc0f3df42} /* (10, 2, 10) {real, imag} */,
  {32'h4194ba79, 32'hc154bcbe} /* (10, 2, 9) {real, imag} */,
  {32'h4141752a, 32'hc1357c79} /* (10, 2, 8) {real, imag} */,
  {32'h41589aae, 32'h40f5b4ce} /* (10, 2, 7) {real, imag} */,
  {32'h4179f959, 32'h4079caa5} /* (10, 2, 6) {real, imag} */,
  {32'h402d5c38, 32'h3fce6f0c} /* (10, 2, 5) {real, imag} */,
  {32'h414ea890, 32'hbf7d1a40} /* (10, 2, 4) {real, imag} */,
  {32'h40325650, 32'h41198f36} /* (10, 2, 3) {real, imag} */,
  {32'hc119faca, 32'h3f92badc} /* (10, 2, 2) {real, imag} */,
  {32'hc0af9b58, 32'hc107bbad} /* (10, 2, 1) {real, imag} */,
  {32'hbea53200, 32'hc0e4bb9b} /* (10, 2, 0) {real, imag} */,
  {32'hc02cb100, 32'h40cb1f0e} /* (10, 1, 31) {real, imag} */,
  {32'hc1871877, 32'h3fbea500} /* (10, 1, 30) {real, imag} */,
  {32'hc1553fac, 32'h4011f874} /* (10, 1, 29) {real, imag} */,
  {32'hc178e956, 32'hc0bac324} /* (10, 1, 28) {real, imag} */,
  {32'hc0abbea6, 32'hc00fff5d} /* (10, 1, 27) {real, imag} */,
  {32'hc109a62b, 32'h413ed9b5} /* (10, 1, 26) {real, imag} */,
  {32'hc18edbe5, 32'h40b263b5} /* (10, 1, 25) {real, imag} */,
  {32'hc1aed479, 32'h40ffb03a} /* (10, 1, 24) {real, imag} */,
  {32'hc138571e, 32'h412de024} /* (10, 1, 23) {real, imag} */,
  {32'hbf75267f, 32'h40ec14eb} /* (10, 1, 22) {real, imag} */,
  {32'h402df548, 32'hbef05f28} /* (10, 1, 21) {real, imag} */,
  {32'h414af31e, 32'hc05e1c99} /* (10, 1, 20) {real, imag} */,
  {32'h41082f64, 32'hc115a2e4} /* (10, 1, 19) {real, imag} */,
  {32'h419fe08a, 32'hbfc872e8} /* (10, 1, 18) {real, imag} */,
  {32'h418cac86, 32'h3ea264c2} /* (10, 1, 17) {real, imag} */,
  {32'hbeb0e876, 32'h4141813e} /* (10, 1, 16) {real, imag} */,
  {32'hbf2507f2, 32'h40abdf31} /* (10, 1, 15) {real, imag} */,
  {32'h4036a13c, 32'h3fc3fda4} /* (10, 1, 14) {real, imag} */,
  {32'hbe1eff00, 32'hc15f204e} /* (10, 1, 13) {real, imag} */,
  {32'h40bff168, 32'hc0a7656c} /* (10, 1, 12) {real, imag} */,
  {32'h41931991, 32'h410a0e73} /* (10, 1, 11) {real, imag} */,
  {32'h3f330228, 32'h412531da} /* (10, 1, 10) {real, imag} */,
  {32'h3eb09148, 32'h400d635c} /* (10, 1, 9) {real, imag} */,
  {32'hc024ff82, 32'hc0270ef8} /* (10, 1, 8) {real, imag} */,
  {32'hc06fb9c0, 32'h3fa24e6c} /* (10, 1, 7) {real, imag} */,
  {32'hbeed0300, 32'hc08bb020} /* (10, 1, 6) {real, imag} */,
  {32'h3e699508, 32'h3fcbfe20} /* (10, 1, 5) {real, imag} */,
  {32'hc11ca504, 32'h3ec6cc40} /* (10, 1, 4) {real, imag} */,
  {32'hc129e2bf, 32'hc0a075e4} /* (10, 1, 3) {real, imag} */,
  {32'hc11a2662, 32'hc0ec5b22} /* (10, 1, 2) {real, imag} */,
  {32'hc0433d10, 32'hbfd212c0} /* (10, 1, 1) {real, imag} */,
  {32'h3fd97000, 32'h415fa7e2} /* (10, 1, 0) {real, imag} */,
  {32'h40b1f3aa, 32'h3f792f0e} /* (10, 0, 31) {real, imag} */,
  {32'h3f9dbf1d, 32'hbda3fd00} /* (10, 0, 30) {real, imag} */,
  {32'hc11437e6, 32'h3f2e96a8} /* (10, 0, 29) {real, imag} */,
  {32'hc1a1e3b0, 32'h410808a1} /* (10, 0, 28) {real, imag} */,
  {32'hc13ccad3, 32'hc0e5ced3} /* (10, 0, 27) {real, imag} */,
  {32'h3fc8183c, 32'hc103867c} /* (10, 0, 26) {real, imag} */,
  {32'h405d4733, 32'hc0013df8} /* (10, 0, 25) {real, imag} */,
  {32'h3f7ea312, 32'h40fffddc} /* (10, 0, 24) {real, imag} */,
  {32'hc18bd9c2, 32'h412115a7} /* (10, 0, 23) {real, imag} */,
  {32'hc13d46f4, 32'h40e6863f} /* (10, 0, 22) {real, imag} */,
  {32'hbfba0551, 32'hc0e94e65} /* (10, 0, 21) {real, imag} */,
  {32'hc13195da, 32'h3fb68874} /* (10, 0, 20) {real, imag} */,
  {32'h40039e22, 32'h40e4b31e} /* (10, 0, 19) {real, imag} */,
  {32'h414f35f4, 32'h413222c2} /* (10, 0, 18) {real, imag} */,
  {32'h4168f57e, 32'h3fc897a4} /* (10, 0, 17) {real, imag} */,
  {32'h3f315442, 32'hc0a7b30a} /* (10, 0, 16) {real, imag} */,
  {32'h40a79cda, 32'hc16da39a} /* (10, 0, 15) {real, imag} */,
  {32'h41a99bae, 32'hc0c6fb5b} /* (10, 0, 14) {real, imag} */,
  {32'h4014a2f0, 32'h40c686c8} /* (10, 0, 13) {real, imag} */,
  {32'hc0d37f5c, 32'h407b2523} /* (10, 0, 12) {real, imag} */,
  {32'hc0bdb3e8, 32'hc05f375c} /* (10, 0, 11) {real, imag} */,
  {32'hc09e03e4, 32'hc0373aa8} /* (10, 0, 10) {real, imag} */,
  {32'hc10caa93, 32'hc1663c62} /* (10, 0, 9) {real, imag} */,
  {32'h400cab37, 32'h3fdf1674} /* (10, 0, 8) {real, imag} */,
  {32'h4162c4c4, 32'h40acbcea} /* (10, 0, 7) {real, imag} */,
  {32'h418664a8, 32'h3fab202e} /* (10, 0, 6) {real, imag} */,
  {32'h4003cf24, 32'h405d5521} /* (10, 0, 5) {real, imag} */,
  {32'h4102ea60, 32'h4123a64c} /* (10, 0, 4) {real, imag} */,
  {32'hbf225487, 32'hbfbb9071} /* (10, 0, 3) {real, imag} */,
  {32'hc188f2e5, 32'hc186f244} /* (10, 0, 2) {real, imag} */,
  {32'hc1b5ffcc, 32'hc1be9762} /* (10, 0, 1) {real, imag} */,
  {32'hc01e5004, 32'hc13b1128} /* (10, 0, 0) {real, imag} */,
  {32'hc13b1cb6, 32'h412f5225} /* (9, 31, 31) {real, imag} */,
  {32'hc113b850, 32'h41400f94} /* (9, 31, 30) {real, imag} */,
  {32'hc097d0b8, 32'h4089e24d} /* (9, 31, 29) {real, imag} */,
  {32'hc0b816fa, 32'h40136bf4} /* (9, 31, 28) {real, imag} */,
  {32'hc0124a5e, 32'h3e59a7c0} /* (9, 31, 27) {real, imag} */,
  {32'h413852bd, 32'h415f3c11} /* (9, 31, 26) {real, imag} */,
  {32'hc18c589b, 32'h40eda7b8} /* (9, 31, 25) {real, imag} */,
  {32'hc184bf50, 32'h4120aa9a} /* (9, 31, 24) {real, imag} */,
  {32'hc068232b, 32'h4147c085} /* (9, 31, 23) {real, imag} */,
  {32'hc09a069b, 32'h418d6893} /* (9, 31, 22) {real, imag} */,
  {32'hc115992a, 32'hc05a4acc} /* (9, 31, 21) {real, imag} */,
  {32'hc07e04e9, 32'hc16603ea} /* (9, 31, 20) {real, imag} */,
  {32'h3f65a370, 32'hc1238449} /* (9, 31, 19) {real, imag} */,
  {32'h40da693e, 32'hc0e68004} /* (9, 31, 18) {real, imag} */,
  {32'hc107cfe0, 32'hc0f262be} /* (9, 31, 17) {real, imag} */,
  {32'hc14049da, 32'hc10d630c} /* (9, 31, 16) {real, imag} */,
  {32'hbc1ae600, 32'hc0ed6e38} /* (9, 31, 15) {real, imag} */,
  {32'h40f5f39b, 32'h400468a4} /* (9, 31, 14) {real, imag} */,
  {32'h40e8ab02, 32'hc0b0c7b6} /* (9, 31, 13) {real, imag} */,
  {32'h40ac807c, 32'hbfe62c20} /* (9, 31, 12) {real, imag} */,
  {32'h4131f815, 32'hbfd23648} /* (9, 31, 11) {real, imag} */,
  {32'hbfaef480, 32'h41169489} /* (9, 31, 10) {real, imag} */,
  {32'h3f1bf010, 32'h406e9b0e} /* (9, 31, 9) {real, imag} */,
  {32'h412f5dc6, 32'h40244400} /* (9, 31, 8) {real, imag} */,
  {32'hc0f80843, 32'h412cde52} /* (9, 31, 7) {real, imag} */,
  {32'hc0f7480a, 32'h41257578} /* (9, 31, 6) {real, imag} */,
  {32'hc1214b96, 32'h40bb3776} /* (9, 31, 5) {real, imag} */,
  {32'hc149fa6b, 32'h40e23d41} /* (9, 31, 4) {real, imag} */,
  {32'hc149f43e, 32'h41545a7f} /* (9, 31, 3) {real, imag} */,
  {32'hc1515fb7, 32'h41367886} /* (9, 31, 2) {real, imag} */,
  {32'hc14c30e3, 32'h41b747a4} /* (9, 31, 1) {real, imag} */,
  {32'hc0616ee2, 32'h413c0b17} /* (9, 31, 0) {real, imag} */,
  {32'hc07cb027, 32'h40ae2b15} /* (9, 30, 31) {real, imag} */,
  {32'h4109af42, 32'h41053e11} /* (9, 30, 30) {real, imag} */,
  {32'h418dc360, 32'h4135aa87} /* (9, 30, 29) {real, imag} */,
  {32'h404d8758, 32'hbf41da6b} /* (9, 30, 28) {real, imag} */,
  {32'hc125b05b, 32'hbeac20e0} /* (9, 30, 27) {real, imag} */,
  {32'hbf88fe88, 32'h3f6589d0} /* (9, 30, 26) {real, imag} */,
  {32'h4010d3f3, 32'hc171af80} /* (9, 30, 25) {real, imag} */,
  {32'h40b1a65c, 32'hc17c9fc3} /* (9, 30, 24) {real, imag} */,
  {32'hc0da6856, 32'hc18e5593} /* (9, 30, 23) {real, imag} */,
  {32'hc14f3279, 32'hc1ae24e3} /* (9, 30, 22) {real, imag} */,
  {32'hc0f0fc04, 32'hbe971a10} /* (9, 30, 21) {real, imag} */,
  {32'hc0672a26, 32'h40edaa00} /* (9, 30, 20) {real, imag} */,
  {32'hc065b15e, 32'hc00801d4} /* (9, 30, 19) {real, imag} */,
  {32'hc0c5dd04, 32'h40c9a0cd} /* (9, 30, 18) {real, imag} */,
  {32'hbfe86476, 32'h41652fc0} /* (9, 30, 17) {real, imag} */,
  {32'hc1927446, 32'h4141e396} /* (9, 30, 16) {real, imag} */,
  {32'hc1799aba, 32'h40b4d511} /* (9, 30, 15) {real, imag} */,
  {32'hbfce2726, 32'hc0c2c74c} /* (9, 30, 14) {real, imag} */,
  {32'hc0bd27ca, 32'hc160eae0} /* (9, 30, 13) {real, imag} */,
  {32'hc1a9a688, 32'hc10b1d2a} /* (9, 30, 12) {real, imag} */,
  {32'hc15cc4d8, 32'h4110f6e9} /* (9, 30, 11) {real, imag} */,
  {32'h409ce08c, 32'h3ed4bf6a} /* (9, 30, 10) {real, imag} */,
  {32'h417ddb31, 32'hc0fe8a51} /* (9, 30, 9) {real, imag} */,
  {32'h416d3cc2, 32'h4037d848} /* (9, 30, 8) {real, imag} */,
  {32'h416ba212, 32'hc15d39fa} /* (9, 30, 7) {real, imag} */,
  {32'h4111a860, 32'hc1584e8b} /* (9, 30, 6) {real, imag} */,
  {32'h41a77a06, 32'hc16ed6b6} /* (9, 30, 5) {real, imag} */,
  {32'h41756e41, 32'hc0149268} /* (9, 30, 4) {real, imag} */,
  {32'h3d827cf8, 32'h4185b188} /* (9, 30, 3) {real, imag} */,
  {32'hc0648104, 32'hc0ac66e4} /* (9, 30, 2) {real, imag} */,
  {32'h403cd3cc, 32'hc0e8062a} /* (9, 30, 1) {real, imag} */,
  {32'hbf8762ff, 32'h400e8ce8} /* (9, 30, 0) {real, imag} */,
  {32'hc127d49e, 32'h40008f14} /* (9, 29, 31) {real, imag} */,
  {32'hc17befad, 32'hbf5af866} /* (9, 29, 30) {real, imag} */,
  {32'hc0274394, 32'hc117d82f} /* (9, 29, 29) {real, imag} */,
  {32'hc0a81daa, 32'hbea680b8} /* (9, 29, 28) {real, imag} */,
  {32'hc10923c8, 32'h40ab8c3d} /* (9, 29, 27) {real, imag} */,
  {32'h404f08c1, 32'h40124a56} /* (9, 29, 26) {real, imag} */,
  {32'h41072a82, 32'h40f9c2f3} /* (9, 29, 25) {real, imag} */,
  {32'hbbfdf000, 32'hbdb1d180} /* (9, 29, 24) {real, imag} */,
  {32'hc0ef403d, 32'h41274ad8} /* (9, 29, 23) {real, imag} */,
  {32'h3f66ca50, 32'h411a17b8} /* (9, 29, 22) {real, imag} */,
  {32'h3e195400, 32'h413265b2} /* (9, 29, 21) {real, imag} */,
  {32'hc08c08f5, 32'h412383be} /* (9, 29, 20) {real, imag} */,
  {32'hbf2ad684, 32'hc0b18da7} /* (9, 29, 19) {real, imag} */,
  {32'hc127e098, 32'hbfee7ebd} /* (9, 29, 18) {real, imag} */,
  {32'hc1a24ef3, 32'h3fc46584} /* (9, 29, 17) {real, imag} */,
  {32'hc11ed7f2, 32'hc151ae57} /* (9, 29, 16) {real, imag} */,
  {32'hc15c6312, 32'hc1042e15} /* (9, 29, 15) {real, imag} */,
  {32'hc08fa0c0, 32'h4008ce98} /* (9, 29, 14) {real, imag} */,
  {32'h41551d02, 32'h3f8ed894} /* (9, 29, 13) {real, imag} */,
  {32'h41929498, 32'h40d58a8c} /* (9, 29, 12) {real, imag} */,
  {32'h40c5ee0c, 32'h3da11c80} /* (9, 29, 11) {real, imag} */,
  {32'h4144c6ee, 32'h407e55d8} /* (9, 29, 10) {real, imag} */,
  {32'h419d55f4, 32'h4165e296} /* (9, 29, 9) {real, imag} */,
  {32'h40f8dae1, 32'h41432487} /* (9, 29, 8) {real, imag} */,
  {32'h4169e898, 32'h41689130} /* (9, 29, 7) {real, imag} */,
  {32'h40c94f9a, 32'h4160e9c2} /* (9, 29, 6) {real, imag} */,
  {32'h41195644, 32'hbd421900} /* (9, 29, 5) {real, imag} */,
  {32'h40bcacb3, 32'hc0c466e4} /* (9, 29, 4) {real, imag} */,
  {32'hc08db558, 32'hc155648a} /* (9, 29, 3) {real, imag} */,
  {32'hc0de423d, 32'hc14e57a0} /* (9, 29, 2) {real, imag} */,
  {32'hbeec1180, 32'h405ac9fc} /* (9, 29, 1) {real, imag} */,
  {32'hc0490ea9, 32'h40c05fbf} /* (9, 29, 0) {real, imag} */,
  {32'h40216df8, 32'h412b002d} /* (9, 28, 31) {real, imag} */,
  {32'h40868b28, 32'h41372d96} /* (9, 28, 30) {real, imag} */,
  {32'hc0ab5371, 32'hbfdab488} /* (9, 28, 29) {real, imag} */,
  {32'hc0323c8a, 32'hc04a45d8} /* (9, 28, 28) {real, imag} */,
  {32'h40be2e15, 32'hc1402fad} /* (9, 28, 27) {real, imag} */,
  {32'h41845b3d, 32'hc15ced7a} /* (9, 28, 26) {real, imag} */,
  {32'h41340e47, 32'hc10bdaf3} /* (9, 28, 25) {real, imag} */,
  {32'h3ffed8ba, 32'h402e1792} /* (9, 28, 24) {real, imag} */,
  {32'h408cbe06, 32'h40f05960} /* (9, 28, 23) {real, imag} */,
  {32'h411882b6, 32'h3f503e50} /* (9, 28, 22) {real, imag} */,
  {32'h40b902de, 32'hbf7d4bb0} /* (9, 28, 21) {real, imag} */,
  {32'h40e52bd2, 32'hc0a0651e} /* (9, 28, 20) {real, imag} */,
  {32'h3f8728e0, 32'hc08329a0} /* (9, 28, 19) {real, imag} */,
  {32'hbfa2f462, 32'hbfcab4f0} /* (9, 28, 18) {real, imag} */,
  {32'hc0868c68, 32'hc1930bd1} /* (9, 28, 17) {real, imag} */,
  {32'h405954fb, 32'hc0cfd778} /* (9, 28, 16) {real, imag} */,
  {32'hc0b891f6, 32'hc04ee788} /* (9, 28, 15) {real, imag} */,
  {32'hc0135ad0, 32'hc0398721} /* (9, 28, 14) {real, imag} */,
  {32'hc1267452, 32'hc17f2f35} /* (9, 28, 13) {real, imag} */,
  {32'hc19bb45f, 32'hc0af4de1} /* (9, 28, 12) {real, imag} */,
  {32'hc039935c, 32'h410df2d4} /* (9, 28, 11) {real, imag} */,
  {32'hc06ff89e, 32'h4105c8b2} /* (9, 28, 10) {real, imag} */,
  {32'hc0b57a8e, 32'hc0c0ea23} /* (9, 28, 9) {real, imag} */,
  {32'hbfcf5fc4, 32'hc0b683fc} /* (9, 28, 8) {real, imag} */,
  {32'hc063bf68, 32'h40e0636d} /* (9, 28, 7) {real, imag} */,
  {32'h410cf2f9, 32'hc040b07e} /* (9, 28, 6) {real, imag} */,
  {32'h4119e027, 32'hc0dfcda3} /* (9, 28, 5) {real, imag} */,
  {32'h40b62e1a, 32'hc116fa92} /* (9, 28, 4) {real, imag} */,
  {32'h3fb254a0, 32'h40fc7d1e} /* (9, 28, 3) {real, imag} */,
  {32'hc0b079a2, 32'h402d0065} /* (9, 28, 2) {real, imag} */,
  {32'hbee25a40, 32'hc1ae053f} /* (9, 28, 1) {real, imag} */,
  {32'h400b886e, 32'hc0c49bf4} /* (9, 28, 0) {real, imag} */,
  {32'h40e0a5da, 32'hc020341a} /* (9, 27, 31) {real, imag} */,
  {32'h4104dd45, 32'hbfb7e72f} /* (9, 27, 30) {real, imag} */,
  {32'h3e2277d8, 32'h40f223ac} /* (9, 27, 29) {real, imag} */,
  {32'h3ff28fbf, 32'hc012dabc} /* (9, 27, 28) {real, imag} */,
  {32'h40feb2f3, 32'hc0e78793} /* (9, 27, 27) {real, imag} */,
  {32'h4014d37c, 32'h3eaf69f0} /* (9, 27, 26) {real, imag} */,
  {32'hc086ac1e, 32'h4006c66a} /* (9, 27, 25) {real, imag} */,
  {32'h3ff4b338, 32'hc13e0f8c} /* (9, 27, 24) {real, imag} */,
  {32'h4159b3f0, 32'hc15a8be4} /* (9, 27, 23) {real, imag} */,
  {32'hbff525d8, 32'h4143bcd4} /* (9, 27, 22) {real, imag} */,
  {32'hc0d866a1, 32'h41892c8c} /* (9, 27, 21) {real, imag} */,
  {32'h3f7f0f72, 32'h4189ca3a} /* (9, 27, 20) {real, imag} */,
  {32'h410d11bf, 32'h41234d54} /* (9, 27, 19) {real, imag} */,
  {32'h40ad42b8, 32'h414abeca} /* (9, 27, 18) {real, imag} */,
  {32'h406f83d0, 32'h4190edf3} /* (9, 27, 17) {real, imag} */,
  {32'hc0d67df2, 32'h40e5a782} /* (9, 27, 16) {real, imag} */,
  {32'hc099c86d, 32'h3fa29858} /* (9, 27, 15) {real, imag} */,
  {32'hbf8b2f70, 32'h3f814338} /* (9, 27, 14) {real, imag} */,
  {32'h405955b6, 32'hc11021ef} /* (9, 27, 13) {real, imag} */,
  {32'hc0627ccc, 32'h3f85fbe8} /* (9, 27, 12) {real, imag} */,
  {32'hc0aa5363, 32'h410269b2} /* (9, 27, 11) {real, imag} */,
  {32'hbf9c4ce5, 32'hc0a86098} /* (9, 27, 10) {real, imag} */,
  {32'hc0b08f5c, 32'hc1489337} /* (9, 27, 9) {real, imag} */,
  {32'h40a91d93, 32'hc03dbdda} /* (9, 27, 8) {real, imag} */,
  {32'h4118715c, 32'hbfe97fe0} /* (9, 27, 7) {real, imag} */,
  {32'hc0d6bb86, 32'h40bf3aba} /* (9, 27, 6) {real, imag} */,
  {32'hc10c7ac0, 32'hbf05c8c8} /* (9, 27, 5) {real, imag} */,
  {32'h41371f1d, 32'h3d7b0910} /* (9, 27, 4) {real, imag} */,
  {32'h4024c67c, 32'hc127e8f2} /* (9, 27, 3) {real, imag} */,
  {32'hc16eddae, 32'hc15a4886} /* (9, 27, 2) {real, imag} */,
  {32'hbf9230df, 32'h408a3e79} /* (9, 27, 1) {real, imag} */,
  {32'h4035caec, 32'h40bd98c0} /* (9, 27, 0) {real, imag} */,
  {32'h40932e53, 32'h4099376c} /* (9, 26, 31) {real, imag} */,
  {32'h411e848e, 32'h3f8e3060} /* (9, 26, 30) {real, imag} */,
  {32'h414c9e06, 32'hc0a879f2} /* (9, 26, 29) {real, imag} */,
  {32'h3f04a478, 32'h3f886dc2} /* (9, 26, 28) {real, imag} */,
  {32'hc0baa56a, 32'h3fd21edb} /* (9, 26, 27) {real, imag} */,
  {32'hbebec180, 32'h3fcbc5aa} /* (9, 26, 26) {real, imag} */,
  {32'hc093604a, 32'hc064917c} /* (9, 26, 25) {real, imag} */,
  {32'h3f7c2522, 32'hbf298ba8} /* (9, 26, 24) {real, imag} */,
  {32'hc0176371, 32'hc1647b22} /* (9, 26, 23) {real, imag} */,
  {32'h3efe666c, 32'hc15bed8f} /* (9, 26, 22) {real, imag} */,
  {32'h40c6bad8, 32'hc10fb92a} /* (9, 26, 21) {real, imag} */,
  {32'hc0aea31a, 32'hc10078d1} /* (9, 26, 20) {real, imag} */,
  {32'hc102f3b4, 32'hc0d46c9c} /* (9, 26, 19) {real, imag} */,
  {32'h40af1b8c, 32'h41188785} /* (9, 26, 18) {real, imag} */,
  {32'h40f6dd02, 32'h413550f0} /* (9, 26, 17) {real, imag} */,
  {32'hc02b22c6, 32'hbfe97b8a} /* (9, 26, 16) {real, imag} */,
  {32'h408fa71d, 32'h4138d3ed} /* (9, 26, 15) {real, imag} */,
  {32'hc00896cc, 32'h4103c629} /* (9, 26, 14) {real, imag} */,
  {32'hc10249cc, 32'hc0f0ed28} /* (9, 26, 13) {real, imag} */,
  {32'hc199a300, 32'hc00d6b6a} /* (9, 26, 12) {real, imag} */,
  {32'hc128242a, 32'h405ce140} /* (9, 26, 11) {real, imag} */,
  {32'hbfd499ec, 32'hbff122d5} /* (9, 26, 10) {real, imag} */,
  {32'h40b8d7a3, 32'h4151f22c} /* (9, 26, 9) {real, imag} */,
  {32'h40d7a044, 32'h41129bc8} /* (9, 26, 8) {real, imag} */,
  {32'hbfcae9b8, 32'h40c073e0} /* (9, 26, 7) {real, imag} */,
  {32'hc1456a62, 32'h4122310c} /* (9, 26, 6) {real, imag} */,
  {32'hc0ab21aa, 32'h412ea869} /* (9, 26, 5) {real, imag} */,
  {32'hbd98a900, 32'hc0970fd8} /* (9, 26, 4) {real, imag} */,
  {32'hc13a0e6a, 32'hc05e5fca} /* (9, 26, 3) {real, imag} */,
  {32'hc1403242, 32'hc17a262c} /* (9, 26, 2) {real, imag} */,
  {32'hc0a6c12d, 32'hc10b9976} /* (9, 26, 1) {real, imag} */,
  {32'hc03799b8, 32'hc0c39e08} /* (9, 26, 0) {real, imag} */,
  {32'h406b4321, 32'hc0dfb3c0} /* (9, 25, 31) {real, imag} */,
  {32'h4020e20e, 32'hc130c323} /* (9, 25, 30) {real, imag} */,
  {32'hc0a0c1f5, 32'h3fec2fa4} /* (9, 25, 29) {real, imag} */,
  {32'h41358e7e, 32'h4128e16f} /* (9, 25, 28) {real, imag} */,
  {32'h4156544e, 32'h40a3aee5} /* (9, 25, 27) {real, imag} */,
  {32'h40b44d32, 32'h4061197c} /* (9, 25, 26) {real, imag} */,
  {32'h409325b3, 32'h4084709b} /* (9, 25, 25) {real, imag} */,
  {32'h4120039f, 32'hc02b9210} /* (9, 25, 24) {real, imag} */,
  {32'h408cb8e2, 32'h409b461e} /* (9, 25, 23) {real, imag} */,
  {32'hc0220eb3, 32'h408eef0f} /* (9, 25, 22) {real, imag} */,
  {32'h3fb394fa, 32'h4045a7ce} /* (9, 25, 21) {real, imag} */,
  {32'h40e33d79, 32'hc0b6de8e} /* (9, 25, 20) {real, imag} */,
  {32'h408bb5b7, 32'hc08b4f01} /* (9, 25, 19) {real, imag} */,
  {32'hc0cbcfd6, 32'hc13c133f} /* (9, 25, 18) {real, imag} */,
  {32'hc0e55020, 32'hc1354323} /* (9, 25, 17) {real, imag} */,
  {32'hc04aeb64, 32'hbf80ac9b} /* (9, 25, 16) {real, imag} */,
  {32'hc0151cc6, 32'hbdee6800} /* (9, 25, 15) {real, imag} */,
  {32'h40c00cdf, 32'hc08be995} /* (9, 25, 14) {real, imag} */,
  {32'h401f637e, 32'hbfda9498} /* (9, 25, 13) {real, imag} */,
  {32'hc032ae54, 32'hc13122f6} /* (9, 25, 12) {real, imag} */,
  {32'hc115c542, 32'hc0b7f0f7} /* (9, 25, 11) {real, imag} */,
  {32'hc15a6cb4, 32'h405641c6} /* (9, 25, 10) {real, imag} */,
  {32'hbfdfbff6, 32'h408a851e} /* (9, 25, 9) {real, imag} */,
  {32'h4117709e, 32'h403d2021} /* (9, 25, 8) {real, imag} */,
  {32'h3fead27a, 32'h3ff09f37} /* (9, 25, 7) {real, imag} */,
  {32'hc17bab98, 32'h404ab4f7} /* (9, 25, 6) {real, imag} */,
  {32'hc1575903, 32'hc0320e53} /* (9, 25, 5) {real, imag} */,
  {32'hc10466a3, 32'h40c159a6} /* (9, 25, 4) {real, imag} */,
  {32'hbf62f1d4, 32'h40609b58} /* (9, 25, 3) {real, imag} */,
  {32'h4174de00, 32'h3f6a2e20} /* (9, 25, 2) {real, imag} */,
  {32'h412cdec0, 32'h4067d921} /* (9, 25, 1) {real, imag} */,
  {32'h3fbd69f4, 32'hbfb22fe2} /* (9, 25, 0) {real, imag} */,
  {32'h3fbc8e92, 32'hc01f5b68} /* (9, 24, 31) {real, imag} */,
  {32'h40309bbe, 32'hc02dcc5c} /* (9, 24, 30) {real, imag} */,
  {32'hc06d9f4d, 32'hc0a09c50} /* (9, 24, 29) {real, imag} */,
  {32'hc0e37a19, 32'hbe9140a0} /* (9, 24, 28) {real, imag} */,
  {32'hc0150959, 32'h404aef81} /* (9, 24, 27) {real, imag} */,
  {32'hc0691306, 32'hc0d6468f} /* (9, 24, 26) {real, imag} */,
  {32'h4114c3ce, 32'hc09a7d16} /* (9, 24, 25) {real, imag} */,
  {32'h40f13a31, 32'hbf69fad6} /* (9, 24, 24) {real, imag} */,
  {32'hc093836e, 32'hc04a1c2e} /* (9, 24, 23) {real, imag} */,
  {32'hc10b6c07, 32'hc0c13c73} /* (9, 24, 22) {real, imag} */,
  {32'hc1645050, 32'hc184ee48} /* (9, 24, 21) {real, imag} */,
  {32'hc091c182, 32'hc095b01b} /* (9, 24, 20) {real, imag} */,
  {32'h401feac0, 32'h3ff3e8aa} /* (9, 24, 19) {real, imag} */,
  {32'h3bdf3180, 32'h40b65d74} /* (9, 24, 18) {real, imag} */,
  {32'hbf698484, 32'hbd6a5d80} /* (9, 24, 17) {real, imag} */,
  {32'h3f1756d0, 32'hbf7c65ae} /* (9, 24, 16) {real, imag} */,
  {32'hc09dbea0, 32'hbf959f16} /* (9, 24, 15) {real, imag} */,
  {32'hc0983992, 32'hc0330df4} /* (9, 24, 14) {real, imag} */,
  {32'hc097ac61, 32'hc10270f9} /* (9, 24, 13) {real, imag} */,
  {32'h404e2a36, 32'hc0a248b1} /* (9, 24, 12) {real, imag} */,
  {32'h409ab6a3, 32'hc02f8143} /* (9, 24, 11) {real, imag} */,
  {32'h40187930, 32'hbf5b5868} /* (9, 24, 10) {real, imag} */,
  {32'h40c769f8, 32'hc10a61a1} /* (9, 24, 9) {real, imag} */,
  {32'hc08d76a6, 32'hbf648c50} /* (9, 24, 8) {real, imag} */,
  {32'h40c3f133, 32'hc0106eb2} /* (9, 24, 7) {real, imag} */,
  {32'h40a807ad, 32'hc11fb0b7} /* (9, 24, 6) {real, imag} */,
  {32'hbf0d3260, 32'hbf9ca1d4} /* (9, 24, 5) {real, imag} */,
  {32'h3f97b650, 32'h40a0bbdb} /* (9, 24, 4) {real, imag} */,
  {32'h40882945, 32'h3fc2b33a} /* (9, 24, 3) {real, imag} */,
  {32'hc0a6fac2, 32'h40802100} /* (9, 24, 2) {real, imag} */,
  {32'hc0ef61fa, 32'h4088db6d} /* (9, 24, 1) {real, imag} */,
  {32'h3fb24a78, 32'h4004f30e} /* (9, 24, 0) {real, imag} */,
  {32'h405fbe96, 32'hc08c3070} /* (9, 23, 31) {real, imag} */,
  {32'h3fa876e5, 32'hc0ad4432} /* (9, 23, 30) {real, imag} */,
  {32'hbdf7c6d8, 32'hbfb77d3a} /* (9, 23, 29) {real, imag} */,
  {32'h40f116b0, 32'hbff42232} /* (9, 23, 28) {real, imag} */,
  {32'h4045c8c5, 32'hc081b61c} /* (9, 23, 27) {real, imag} */,
  {32'hbf94263a, 32'hbd015460} /* (9, 23, 26) {real, imag} */,
  {32'h4055ae68, 32'h4056a911} /* (9, 23, 25) {real, imag} */,
  {32'h4110bd4f, 32'hc04153f0} /* (9, 23, 24) {real, imag} */,
  {32'h40bcda42, 32'hbf159d40} /* (9, 23, 23) {real, imag} */,
  {32'h40a62e40, 32'hc00c94ea} /* (9, 23, 22) {real, imag} */,
  {32'h40e99010, 32'h4011b202} /* (9, 23, 21) {real, imag} */,
  {32'h40f4fab6, 32'hc06e44e3} /* (9, 23, 20) {real, imag} */,
  {32'h403d1fd9, 32'hc134ba8e} /* (9, 23, 19) {real, imag} */,
  {32'hbfb075cd, 32'hbf89a860} /* (9, 23, 18) {real, imag} */,
  {32'h3fab662c, 32'h401b2175} /* (9, 23, 17) {real, imag} */,
  {32'h40e3ee6c, 32'h40b09e18} /* (9, 23, 16) {real, imag} */,
  {32'h4087f243, 32'h40ed5a72} /* (9, 23, 15) {real, imag} */,
  {32'hc0d4d4d0, 32'h40bcb0e3} /* (9, 23, 14) {real, imag} */,
  {32'hbdc57370, 32'h40ac960f} /* (9, 23, 13) {real, imag} */,
  {32'h402ed3df, 32'hbee88d28} /* (9, 23, 12) {real, imag} */,
  {32'hbfed2816, 32'hc091b429} /* (9, 23, 11) {real, imag} */,
  {32'hc0d71545, 32'h4098b216} /* (9, 23, 10) {real, imag} */,
  {32'hc11810d4, 32'h40b737cb} /* (9, 23, 9) {real, imag} */,
  {32'hc083f3e7, 32'h40a62cf6} /* (9, 23, 8) {real, imag} */,
  {32'hc0b0f7da, 32'h407433c2} /* (9, 23, 7) {real, imag} */,
  {32'hbfc39c53, 32'h4108b740} /* (9, 23, 6) {real, imag} */,
  {32'h3fbbc21c, 32'h4066f977} /* (9, 23, 5) {real, imag} */,
  {32'hc0ab153c, 32'hc0cd7fda} /* (9, 23, 4) {real, imag} */,
  {32'hc122a92a, 32'hc10d0572} /* (9, 23, 3) {real, imag} */,
  {32'hc07fda9c, 32'hc004eae6} /* (9, 23, 2) {real, imag} */,
  {32'hbf534714, 32'h40a1b97c} /* (9, 23, 1) {real, imag} */,
  {32'hbfad2d4c, 32'h403eace6} /* (9, 23, 0) {real, imag} */,
  {32'hbf400f02, 32'hc01a1d57} /* (9, 22, 31) {real, imag} */,
  {32'hc02c617e, 32'hc0bc0d22} /* (9, 22, 30) {real, imag} */,
  {32'hbff6757c, 32'hc0ac2765} /* (9, 22, 29) {real, imag} */,
  {32'hc035a72f, 32'h3e9f92a8} /* (9, 22, 28) {real, imag} */,
  {32'h3f6f7ef6, 32'hbfecdd4c} /* (9, 22, 27) {real, imag} */,
  {32'h40d736f8, 32'h3fe93e80} /* (9, 22, 26) {real, imag} */,
  {32'h4086bf58, 32'h3ec2d82c} /* (9, 22, 25) {real, imag} */,
  {32'hbfce0fff, 32'h40938695} /* (9, 22, 24) {real, imag} */,
  {32'hc114c7e0, 32'hbded7068} /* (9, 22, 23) {real, imag} */,
  {32'hc11e5818, 32'hc0a87a86} /* (9, 22, 22) {real, imag} */,
  {32'hbfded450, 32'h401ec1c4} /* (9, 22, 21) {real, imag} */,
  {32'hbfdf5726, 32'h3f1a8cc0} /* (9, 22, 20) {real, imag} */,
  {32'hc05584f9, 32'hc042e2ce} /* (9, 22, 19) {real, imag} */,
  {32'hc02536b6, 32'hc0525d23} /* (9, 22, 18) {real, imag} */,
  {32'h3fb5c2da, 32'hc10e29e5} /* (9, 22, 17) {real, imag} */,
  {32'h403dcbd5, 32'hc0a62086} /* (9, 22, 16) {real, imag} */,
  {32'hbf8d05a6, 32'h3f043390} /* (9, 22, 15) {real, imag} */,
  {32'h3fe750b0, 32'h3fae3b3e} /* (9, 22, 14) {real, imag} */,
  {32'h3fc540b1, 32'hbfc0d200} /* (9, 22, 13) {real, imag} */,
  {32'hbebc3e50, 32'h404ec0a0} /* (9, 22, 12) {real, imag} */,
  {32'h41226df0, 32'h408f91bc} /* (9, 22, 11) {real, imag} */,
  {32'h4165cf80, 32'h408fd9d3} /* (9, 22, 10) {real, imag} */,
  {32'h409e0720, 32'h401cfec8} /* (9, 22, 9) {real, imag} */,
  {32'hbd106240, 32'hc013b676} /* (9, 22, 8) {real, imag} */,
  {32'hc03bc450, 32'hbe5b4ad0} /* (9, 22, 7) {real, imag} */,
  {32'h3fa42b25, 32'h40f545ec} /* (9, 22, 6) {real, imag} */,
  {32'hbfa1c2cf, 32'h40c1d4c6} /* (9, 22, 5) {real, imag} */,
  {32'hc09dbe72, 32'h40c1af38} /* (9, 22, 4) {real, imag} */,
  {32'h40773d8a, 32'hc046c71c} /* (9, 22, 3) {real, imag} */,
  {32'h40706ab2, 32'hbeb4ce10} /* (9, 22, 2) {real, imag} */,
  {32'h4000b2a4, 32'h40a2d964} /* (9, 22, 1) {real, imag} */,
  {32'h40260a28, 32'h3e6df0d4} /* (9, 22, 0) {real, imag} */,
  {32'h3d4a6f80, 32'hbe458798} /* (9, 21, 31) {real, imag} */,
  {32'hbfcf7cb8, 32'h3f4c99fc} /* (9, 21, 30) {real, imag} */,
  {32'hc031e27e, 32'h40171adc} /* (9, 21, 29) {real, imag} */,
  {32'h408b111e, 32'hbe4228b0} /* (9, 21, 28) {real, imag} */,
  {32'h40db90ee, 32'h40112460} /* (9, 21, 27) {real, imag} */,
  {32'h40210c91, 32'hc0260c5e} /* (9, 21, 26) {real, imag} */,
  {32'hc0772e4a, 32'hbd28fe10} /* (9, 21, 25) {real, imag} */,
  {32'hc0613f7f, 32'hbe899ec0} /* (9, 21, 24) {real, imag} */,
  {32'h3e273180, 32'hc087bf03} /* (9, 21, 23) {real, imag} */,
  {32'hc03186f5, 32'hbf651dc8} /* (9, 21, 22) {real, imag} */,
  {32'hbfed7950, 32'h4040ae37} /* (9, 21, 21) {real, imag} */,
  {32'h3facf76e, 32'h40f4d451} /* (9, 21, 20) {real, imag} */,
  {32'hbfab202d, 32'h40399027} /* (9, 21, 19) {real, imag} */,
  {32'hc0132854, 32'hc06a2b18} /* (9, 21, 18) {real, imag} */,
  {32'hc0378688, 32'hc0bfb899} /* (9, 21, 17) {real, imag} */,
  {32'h4005ea99, 32'hc0c6a394} /* (9, 21, 16) {real, imag} */,
  {32'h4080b41f, 32'hbf62e089} /* (9, 21, 15) {real, imag} */,
  {32'h40a5ba5d, 32'h4085bbf0} /* (9, 21, 14) {real, imag} */,
  {32'h40f09e9e, 32'h411f0dd0} /* (9, 21, 13) {real, imag} */,
  {32'h40ab87ee, 32'h40670721} /* (9, 21, 12) {real, imag} */,
  {32'h40887889, 32'hc068b4ae} /* (9, 21, 11) {real, imag} */,
  {32'hbe418f30, 32'hbfcdd8bc} /* (9, 21, 10) {real, imag} */,
  {32'hbf12fc0c, 32'h4095e36e} /* (9, 21, 9) {real, imag} */,
  {32'hc0a3865d, 32'h405e7f8e} /* (9, 21, 8) {real, imag} */,
  {32'hc0a0a856, 32'h3fa109b0} /* (9, 21, 7) {real, imag} */,
  {32'h4009afaf, 32'h3fba2e0a} /* (9, 21, 6) {real, imag} */,
  {32'h40a15591, 32'hc03edf86} /* (9, 21, 5) {real, imag} */,
  {32'hbfb7d88b, 32'h406cbaf0} /* (9, 21, 4) {real, imag} */,
  {32'hc054def1, 32'h410057b5} /* (9, 21, 3) {real, imag} */,
  {32'h3e94c798, 32'h3f07f218} /* (9, 21, 2) {real, imag} */,
  {32'h40298144, 32'hc0460f56} /* (9, 21, 1) {real, imag} */,
  {32'h403183b4, 32'h3f6ff310} /* (9, 21, 0) {real, imag} */,
  {32'hbfbe8d02, 32'hc026d57a} /* (9, 20, 31) {real, imag} */,
  {32'hbf6760e0, 32'h3fde9bb8} /* (9, 20, 30) {real, imag} */,
  {32'h3fa4836f, 32'h4082bca5} /* (9, 20, 29) {real, imag} */,
  {32'hbfa4dfb1, 32'h40132920} /* (9, 20, 28) {real, imag} */,
  {32'hbf867fbc, 32'h401cff98} /* (9, 20, 27) {real, imag} */,
  {32'hbf9ca73d, 32'h403dfe45} /* (9, 20, 26) {real, imag} */,
  {32'hbefd6f78, 32'hbec45eb0} /* (9, 20, 25) {real, imag} */,
  {32'h3f4949ba, 32'hc039e90e} /* (9, 20, 24) {real, imag} */,
  {32'h408f8f2a, 32'h3f03e746} /* (9, 20, 23) {real, imag} */,
  {32'h3ed6f040, 32'hbfbbd662} /* (9, 20, 22) {real, imag} */,
  {32'hc066ca5e, 32'hc062c478} /* (9, 20, 21) {real, imag} */,
  {32'h3f3d9180, 32'hbf6fd9ee} /* (9, 20, 20) {real, imag} */,
  {32'hbf9189a2, 32'hc0027af0} /* (9, 20, 19) {real, imag} */,
  {32'hc00a78b4, 32'h4074635f} /* (9, 20, 18) {real, imag} */,
  {32'hbec3c098, 32'h4097c365} /* (9, 20, 17) {real, imag} */,
  {32'h40bac600, 32'hbf85189e} /* (9, 20, 16) {real, imag} */,
  {32'h4022def2, 32'h3fe6320b} /* (9, 20, 15) {real, imag} */,
  {32'hc07214e6, 32'h404693ba} /* (9, 20, 14) {real, imag} */,
  {32'h3fba87f6, 32'h4012ade8} /* (9, 20, 13) {real, imag} */,
  {32'hbfddaff8, 32'hbf9d8217} /* (9, 20, 12) {real, imag} */,
  {32'h3f1512e8, 32'hc0b7bad2} /* (9, 20, 11) {real, imag} */,
  {32'h40563d80, 32'hbf2ac986} /* (9, 20, 10) {real, imag} */,
  {32'hbf3e3b32, 32'h40959d46} /* (9, 20, 9) {real, imag} */,
  {32'h3f889cf4, 32'h40bed81b} /* (9, 20, 8) {real, imag} */,
  {32'h3fec2aae, 32'h3fc540c9} /* (9, 20, 7) {real, imag} */,
  {32'h4025da4e, 32'hbfd10d29} /* (9, 20, 6) {real, imag} */,
  {32'h40d4b506, 32'hbfcf864b} /* (9, 20, 5) {real, imag} */,
  {32'h3ee10d08, 32'hc004a0aa} /* (9, 20, 4) {real, imag} */,
  {32'hc00faa08, 32'hc0b4af39} /* (9, 20, 3) {real, imag} */,
  {32'h40d3b98a, 32'hbff92392} /* (9, 20, 2) {real, imag} */,
  {32'h409276b8, 32'hbfb93c08} /* (9, 20, 1) {real, imag} */,
  {32'hbecf47dc, 32'hbf9e4be0} /* (9, 20, 0) {real, imag} */,
  {32'hc055dc0d, 32'hbf0a122c} /* (9, 19, 31) {real, imag} */,
  {32'hc02a28a9, 32'hc04b2424} /* (9, 19, 30) {real, imag} */,
  {32'hbe6191d0, 32'hc0e37bb8} /* (9, 19, 29) {real, imag} */,
  {32'h3d277880, 32'hc06492a1} /* (9, 19, 28) {real, imag} */,
  {32'h401093f1, 32'hbffbef0b} /* (9, 19, 27) {real, imag} */,
  {32'hc0a8c3a8, 32'hbe5b989c} /* (9, 19, 26) {real, imag} */,
  {32'hc0091b3d, 32'hc01d1d7b} /* (9, 19, 25) {real, imag} */,
  {32'hbf81081c, 32'hc067cae6} /* (9, 19, 24) {real, imag} */,
  {32'hc0914f7e, 32'hc03eb100} /* (9, 19, 23) {real, imag} */,
  {32'hc0968328, 32'hc01f7fa5} /* (9, 19, 22) {real, imag} */,
  {32'h3fc7e20e, 32'hbfea50ae} /* (9, 19, 21) {real, imag} */,
  {32'h3fc79f04, 32'h3f81d261} /* (9, 19, 20) {real, imag} */,
  {32'h3fb846aa, 32'h402de0d8} /* (9, 19, 19) {real, imag} */,
  {32'h40260d90, 32'h3ed84d28} /* (9, 19, 18) {real, imag} */,
  {32'hc00273cc, 32'hc09f5940} /* (9, 19, 17) {real, imag} */,
  {32'hc09e3c58, 32'hc05ac621} /* (9, 19, 16) {real, imag} */,
  {32'hc0b4e386, 32'hbfecacc4} /* (9, 19, 15) {real, imag} */,
  {32'hc09543e3, 32'hc0625c1c} /* (9, 19, 14) {real, imag} */,
  {32'hbfd62290, 32'h3fa5aa30} /* (9, 19, 13) {real, imag} */,
  {32'h3f4788a0, 32'h3fdbbb64} /* (9, 19, 12) {real, imag} */,
  {32'hbf196f1e, 32'h3e813dc0} /* (9, 19, 11) {real, imag} */,
  {32'h3fecdd4b, 32'hc01b989e} /* (9, 19, 10) {real, imag} */,
  {32'h3f819c8a, 32'hc017ff46} /* (9, 19, 9) {real, imag} */,
  {32'h400bdcb2, 32'hc0603fe3} /* (9, 19, 8) {real, imag} */,
  {32'hbecfca58, 32'hbfb43fd6} /* (9, 19, 7) {real, imag} */,
  {32'hc0846744, 32'hc02acbd7} /* (9, 19, 6) {real, imag} */,
  {32'hbe89efc8, 32'hbfa78158} /* (9, 19, 5) {real, imag} */,
  {32'h3fbbb444, 32'h3da14930} /* (9, 19, 4) {real, imag} */,
  {32'hc03011d7, 32'hc03c6d44} /* (9, 19, 3) {real, imag} */,
  {32'h400c00d2, 32'hc08ac110} /* (9, 19, 2) {real, imag} */,
  {32'h3d706500, 32'hc0901eda} /* (9, 19, 1) {real, imag} */,
  {32'hc0030125, 32'hc0575cd7} /* (9, 19, 0) {real, imag} */,
  {32'hbf07dfc0, 32'h3fc6d0dc} /* (9, 18, 31) {real, imag} */,
  {32'h40854d9c, 32'hbee79c46} /* (9, 18, 30) {real, imag} */,
  {32'h4058647c, 32'hc04e817e} /* (9, 18, 29) {real, imag} */,
  {32'hc02b7917, 32'h3ef086c0} /* (9, 18, 28) {real, imag} */,
  {32'hc0157753, 32'h408e7987} /* (9, 18, 27) {real, imag} */,
  {32'hbe1dc6e0, 32'h405945b9} /* (9, 18, 26) {real, imag} */,
  {32'h3ebe2aa0, 32'h3f43478c} /* (9, 18, 25) {real, imag} */,
  {32'hc007e7ac, 32'h3f820d60} /* (9, 18, 24) {real, imag} */,
  {32'hbf840270, 32'h3faf7d22} /* (9, 18, 23) {real, imag} */,
  {32'h4030732d, 32'h4016e65a} /* (9, 18, 22) {real, imag} */,
  {32'h3f08ddb2, 32'h3f3b728a} /* (9, 18, 21) {real, imag} */,
  {32'h3e9edf90, 32'hc013ec2a} /* (9, 18, 20) {real, imag} */,
  {32'h3d583b00, 32'hbfaa7134} /* (9, 18, 19) {real, imag} */,
  {32'hbfe1ee3e, 32'hc05419a2} /* (9, 18, 18) {real, imag} */,
  {32'hbf57f268, 32'hc0df156a} /* (9, 18, 17) {real, imag} */,
  {32'h3f8563a7, 32'hc0793e06} /* (9, 18, 16) {real, imag} */,
  {32'hbff42f68, 32'hc085aee8} /* (9, 18, 15) {real, imag} */,
  {32'h3ed549cc, 32'hbf5291f0} /* (9, 18, 14) {real, imag} */,
  {32'h3fd6b66e, 32'h4057a2c2} /* (9, 18, 13) {real, imag} */,
  {32'h3d2e25c0, 32'hbf096708} /* (9, 18, 12) {real, imag} */,
  {32'h404f92a7, 32'h3ef18d00} /* (9, 18, 11) {real, imag} */,
  {32'h3ff0269e, 32'hbf48759f} /* (9, 18, 10) {real, imag} */,
  {32'h3da66ba0, 32'hbccd3ec0} /* (9, 18, 9) {real, imag} */,
  {32'hc05442fa, 32'h400b2948} /* (9, 18, 8) {real, imag} */,
  {32'hbfb7172c, 32'h3fd8fc38} /* (9, 18, 7) {real, imag} */,
  {32'h4019ebb6, 32'hbf5fe4d0} /* (9, 18, 6) {real, imag} */,
  {32'h40450061, 32'hbfec54e6} /* (9, 18, 5) {real, imag} */,
  {32'h3f0352cc, 32'hc05e1cc6} /* (9, 18, 4) {real, imag} */,
  {32'hbd1c4f40, 32'hbda7d620} /* (9, 18, 3) {real, imag} */,
  {32'hc03df7ce, 32'h3f84b022} /* (9, 18, 2) {real, imag} */,
  {32'hbf95c4bb, 32'h3dc96200} /* (9, 18, 1) {real, imag} */,
  {32'h3f080202, 32'hbe85a8b8} /* (9, 18, 0) {real, imag} */,
  {32'hbf8362ca, 32'hbed1eca4} /* (9, 17, 31) {real, imag} */,
  {32'hbfbbcbf6, 32'hc0420d17} /* (9, 17, 30) {real, imag} */,
  {32'h40053c20, 32'hbfb6209a} /* (9, 17, 29) {real, imag} */,
  {32'h4018a93e, 32'h3eef6b00} /* (9, 17, 28) {real, imag} */,
  {32'hbd956ee0, 32'h3f5c20ac} /* (9, 17, 27) {real, imag} */,
  {32'hc02fa0dd, 32'hbf481624} /* (9, 17, 26) {real, imag} */,
  {32'h3ff1f695, 32'h3def4b90} /* (9, 17, 25) {real, imag} */,
  {32'h3f2bb060, 32'h3ff5eb03} /* (9, 17, 24) {real, imag} */,
  {32'hbfe8f0f7, 32'hbd547800} /* (9, 17, 23) {real, imag} */,
  {32'hbf963517, 32'hbfdcdf20} /* (9, 17, 22) {real, imag} */,
  {32'h400e7691, 32'hc066b52e} /* (9, 17, 21) {real, imag} */,
  {32'h3d334880, 32'hbeccf460} /* (9, 17, 20) {real, imag} */,
  {32'h3fa3133d, 32'h40a11058} /* (9, 17, 19) {real, imag} */,
  {32'h3fa868bd, 32'h3fa22816} /* (9, 17, 18) {real, imag} */,
  {32'hbf9dcc5f, 32'hc08e19b7} /* (9, 17, 17) {real, imag} */,
  {32'h3e75e3b0, 32'hc0762e78} /* (9, 17, 16) {real, imag} */,
  {32'h3f9e000c, 32'hc0aaf18a} /* (9, 17, 15) {real, imag} */,
  {32'h3f0505ce, 32'hc01e4eee} /* (9, 17, 14) {real, imag} */,
  {32'h402854b9, 32'h3f724240} /* (9, 17, 13) {real, imag} */,
  {32'h400a9933, 32'h3fd47368} /* (9, 17, 12) {real, imag} */,
  {32'h3e8a3608, 32'h403afdd8} /* (9, 17, 11) {real, imag} */,
  {32'h3fd78b2c, 32'h400ebb3b} /* (9, 17, 10) {real, imag} */,
  {32'h3faa1a64, 32'h4000b112} /* (9, 17, 9) {real, imag} */,
  {32'h40930beb, 32'h4093ec79} /* (9, 17, 8) {real, imag} */,
  {32'h405d17c5, 32'h407ef8fa} /* (9, 17, 7) {real, imag} */,
  {32'hbfe48b38, 32'hbf948453} /* (9, 17, 6) {real, imag} */,
  {32'hbfd9e0c2, 32'hbfecb106} /* (9, 17, 5) {real, imag} */,
  {32'h3fca6d3b, 32'h3fabcae2} /* (9, 17, 4) {real, imag} */,
  {32'h40740d10, 32'h3ff50812} /* (9, 17, 3) {real, imag} */,
  {32'h3ec8d31c, 32'hbf6bb892} /* (9, 17, 2) {real, imag} */,
  {32'h403cc364, 32'hc008e1fe} /* (9, 17, 1) {real, imag} */,
  {32'h400f2f02, 32'hbe9ad704} /* (9, 17, 0) {real, imag} */,
  {32'h400bb95b, 32'hbe839990} /* (9, 16, 31) {real, imag} */,
  {32'hbf57ab40, 32'hc032b94f} /* (9, 16, 30) {real, imag} */,
  {32'hc011ff1c, 32'h3fe215b4} /* (9, 16, 29) {real, imag} */,
  {32'h3f2b4da0, 32'h3f15e240} /* (9, 16, 28) {real, imag} */,
  {32'h403a735b, 32'h3fac2836} /* (9, 16, 27) {real, imag} */,
  {32'h407d7ee6, 32'hbec4448c} /* (9, 16, 26) {real, imag} */,
  {32'h4008ad16, 32'hc0318640} /* (9, 16, 25) {real, imag} */,
  {32'hc05288bc, 32'hc026c0ec} /* (9, 16, 24) {real, imag} */,
  {32'hbf81b078, 32'hc08d88dd} /* (9, 16, 23) {real, imag} */,
  {32'h3e8ac5f8, 32'hbff931e0} /* (9, 16, 22) {real, imag} */,
  {32'hbfcb1846, 32'hbf81dbb6} /* (9, 16, 21) {real, imag} */,
  {32'h3fa885ec, 32'hbfc7c750} /* (9, 16, 20) {real, imag} */,
  {32'h4039daaa, 32'hc03eba0a} /* (9, 16, 19) {real, imag} */,
  {32'h3f02beb0, 32'hc08a5d6d} /* (9, 16, 18) {real, imag} */,
  {32'h3fd3e9fc, 32'hc026f82a} /* (9, 16, 17) {real, imag} */,
  {32'hbf4819a8, 32'hbe7b11e0} /* (9, 16, 16) {real, imag} */,
  {32'hbf48f880, 32'hbfc83316} /* (9, 16, 15) {real, imag} */,
  {32'h3e25b050, 32'hbfe898bc} /* (9, 16, 14) {real, imag} */,
  {32'hc01cb2f6, 32'hbfccc250} /* (9, 16, 13) {real, imag} */,
  {32'hbf78d790, 32'hc01a0642} /* (9, 16, 12) {real, imag} */,
  {32'h3fa8c9e0, 32'h3d4d4400} /* (9, 16, 11) {real, imag} */,
  {32'hbf48ba32, 32'h3f5409f0} /* (9, 16, 10) {real, imag} */,
  {32'h3f4395e8, 32'h402c93e4} /* (9, 16, 9) {real, imag} */,
  {32'h4029c2b8, 32'hbfd4fa89} /* (9, 16, 8) {real, imag} */,
  {32'h3edbb000, 32'hbeda0078} /* (9, 16, 7) {real, imag} */,
  {32'hbf2950d0, 32'h3e10af18} /* (9, 16, 6) {real, imag} */,
  {32'hc0283956, 32'h3f1d7ef0} /* (9, 16, 5) {real, imag} */,
  {32'hbe2b2e90, 32'hbee26cd8} /* (9, 16, 4) {real, imag} */,
  {32'h3f4fae24, 32'hbf3c9668} /* (9, 16, 3) {real, imag} */,
  {32'hbf081b0e, 32'hbfea1f20} /* (9, 16, 2) {real, imag} */,
  {32'h4015bffa, 32'h3eb68d80} /* (9, 16, 1) {real, imag} */,
  {32'h4012d785, 32'h3f2bf87c} /* (9, 16, 0) {real, imag} */,
  {32'hbfe7f57e, 32'h3fddb97f} /* (9, 15, 31) {real, imag} */,
  {32'h3dc75b60, 32'h40861f7c} /* (9, 15, 30) {real, imag} */,
  {32'hbfad7c00, 32'h40453d43} /* (9, 15, 29) {real, imag} */,
  {32'h3feb7430, 32'hbf7dff20} /* (9, 15, 28) {real, imag} */,
  {32'h3efa8898, 32'hc038841b} /* (9, 15, 27) {real, imag} */,
  {32'hbfe5128a, 32'h3fd0504a} /* (9, 15, 26) {real, imag} */,
  {32'h3fcd938b, 32'h3f32540e} /* (9, 15, 25) {real, imag} */,
  {32'hbd351e00, 32'hbff0dc3b} /* (9, 15, 24) {real, imag} */,
  {32'h3fbfd109, 32'hbfded2d8} /* (9, 15, 23) {real, imag} */,
  {32'h40204488, 32'hc01b600c} /* (9, 15, 22) {real, imag} */,
  {32'h407cd4cf, 32'h3dc5c790} /* (9, 15, 21) {real, imag} */,
  {32'h404fef16, 32'h408477ea} /* (9, 15, 20) {real, imag} */,
  {32'h4005aa68, 32'h3e89de90} /* (9, 15, 19) {real, imag} */,
  {32'hbfd2a0e1, 32'hbfd5453e} /* (9, 15, 18) {real, imag} */,
  {32'hbffc299f, 32'h3f3b4f80} /* (9, 15, 17) {real, imag} */,
  {32'hbf25527c, 32'hbfe53f60} /* (9, 15, 16) {real, imag} */,
  {32'h4032ae96, 32'hbf55cf4c} /* (9, 15, 15) {real, imag} */,
  {32'h3f95a011, 32'hbf53fe08} /* (9, 15, 14) {real, imag} */,
  {32'h4059a3a7, 32'hbf263180} /* (9, 15, 13) {real, imag} */,
  {32'h406f0375, 32'hbf952d98} /* (9, 15, 12) {real, imag} */,
  {32'hbe9af488, 32'hbf360a66} /* (9, 15, 11) {real, imag} */,
  {32'hbf31f758, 32'h3e8176d8} /* (9, 15, 10) {real, imag} */,
  {32'hbf384318, 32'hbfd30509} /* (9, 15, 9) {real, imag} */,
  {32'hbf166c78, 32'hc071fbd6} /* (9, 15, 8) {real, imag} */,
  {32'hbff8f5b2, 32'hbffcf334} /* (9, 15, 7) {real, imag} */,
  {32'hc04ef184, 32'hbecd6c74} /* (9, 15, 6) {real, imag} */,
  {32'hbf854a96, 32'h3fa14e66} /* (9, 15, 5) {real, imag} */,
  {32'hbf24d746, 32'hbf99ae42} /* (9, 15, 4) {real, imag} */,
  {32'h3fa8d358, 32'hc004267f} /* (9, 15, 3) {real, imag} */,
  {32'h401f5cb4, 32'hbf94e7e9} /* (9, 15, 2) {real, imag} */,
  {32'hbf63bdc8, 32'h4007aeea} /* (9, 15, 1) {real, imag} */,
  {32'hbf98b91d, 32'h3fc85bff} /* (9, 15, 0) {real, imag} */,
  {32'h4001a1ea, 32'h40107e58} /* (9, 14, 31) {real, imag} */,
  {32'h3f542334, 32'h3fc5dace} /* (9, 14, 30) {real, imag} */,
  {32'hbde3ef80, 32'hbefcc530} /* (9, 14, 29) {real, imag} */,
  {32'hbf8c372a, 32'hc02014fe} /* (9, 14, 28) {real, imag} */,
  {32'hc0303213, 32'hbf0e3b50} /* (9, 14, 27) {real, imag} */,
  {32'h3fdb6a7c, 32'h4013e2dd} /* (9, 14, 26) {real, imag} */,
  {32'h40f064df, 32'h409650fe} /* (9, 14, 25) {real, imag} */,
  {32'h4095d2ba, 32'h409e5cac} /* (9, 14, 24) {real, imag} */,
  {32'hbf2ac589, 32'h4081377e} /* (9, 14, 23) {real, imag} */,
  {32'hbff34bd6, 32'h407d36de} /* (9, 14, 22) {real, imag} */,
  {32'hbd458d20, 32'h400d0c34} /* (9, 14, 21) {real, imag} */,
  {32'hbf28ae28, 32'hc03eee1a} /* (9, 14, 20) {real, imag} */,
  {32'hbfaa5058, 32'hc08f14b1} /* (9, 14, 19) {real, imag} */,
  {32'hc01d687d, 32'hbe56ce38} /* (9, 14, 18) {real, imag} */,
  {32'h40145794, 32'h3febb778} /* (9, 14, 17) {real, imag} */,
  {32'h400b0d6c, 32'h4052f64a} /* (9, 14, 16) {real, imag} */,
  {32'hbff5e230, 32'hbee78d18} /* (9, 14, 15) {real, imag} */,
  {32'hc06955a4, 32'hbfd1b398} /* (9, 14, 14) {real, imag} */,
  {32'hc05b05fd, 32'hbf170996} /* (9, 14, 13) {real, imag} */,
  {32'h3ecd3cc8, 32'hbff923fc} /* (9, 14, 12) {real, imag} */,
  {32'hbf18427c, 32'hc01cf548} /* (9, 14, 11) {real, imag} */,
  {32'hbfb7983a, 32'h3f634401} /* (9, 14, 10) {real, imag} */,
  {32'h3fc2122e, 32'h401c59ca} /* (9, 14, 9) {real, imag} */,
  {32'h400e4b5a, 32'h40043ac8} /* (9, 14, 8) {real, imag} */,
  {32'h40293fe6, 32'h3ede7660} /* (9, 14, 7) {real, imag} */,
  {32'h405272aa, 32'h3c282800} /* (9, 14, 6) {real, imag} */,
  {32'hbfaf48aa, 32'hc0662bc9} /* (9, 14, 5) {real, imag} */,
  {32'hc092cb0e, 32'hc00bd522} /* (9, 14, 4) {real, imag} */,
  {32'hc007a129, 32'h40371941} /* (9, 14, 3) {real, imag} */,
  {32'hbe511a10, 32'h40a44230} /* (9, 14, 2) {real, imag} */,
  {32'hc07387a6, 32'h40b5dfd0} /* (9, 14, 1) {real, imag} */,
  {32'hc06ecc4e, 32'h404598e9} /* (9, 14, 0) {real, imag} */,
  {32'h4008c41f, 32'hbf831e2e} /* (9, 13, 31) {real, imag} */,
  {32'h3ea0a448, 32'h3e7a6e88} /* (9, 13, 30) {real, imag} */,
  {32'hc01e24f5, 32'hbf85bd42} /* (9, 13, 29) {real, imag} */,
  {32'hc08e8a24, 32'h3fb10002} /* (9, 13, 28) {real, imag} */,
  {32'hc08fe5b4, 32'h40a1e735} /* (9, 13, 27) {real, imag} */,
  {32'hc049516f, 32'h3f891076} /* (9, 13, 26) {real, imag} */,
  {32'hbf46d984, 32'h402aadd1} /* (9, 13, 25) {real, imag} */,
  {32'h40b9acb4, 32'h3fbe9a28} /* (9, 13, 24) {real, imag} */,
  {32'h40c3eee2, 32'hbedc5540} /* (9, 13, 23) {real, imag} */,
  {32'h3f1eb0a4, 32'h3e7979f0} /* (9, 13, 22) {real, imag} */,
  {32'h3e3d8450, 32'hbfcd8026} /* (9, 13, 21) {real, imag} */,
  {32'hbf7f27f8, 32'hc0312864} /* (9, 13, 20) {real, imag} */,
  {32'hc067c173, 32'h3ffb391c} /* (9, 13, 19) {real, imag} */,
  {32'h3f8ec740, 32'h409f6252} /* (9, 13, 18) {real, imag} */,
  {32'h3f15a800, 32'h3faea724} /* (9, 13, 17) {real, imag} */,
  {32'h404d79b8, 32'hc02d6cc7} /* (9, 13, 16) {real, imag} */,
  {32'h40fa68bc, 32'hbfa2367c} /* (9, 13, 15) {real, imag} */,
  {32'h402631ea, 32'hc007515c} /* (9, 13, 14) {real, imag} */,
  {32'h3fb74e40, 32'h3f223160} /* (9, 13, 13) {real, imag} */,
  {32'hbf259780, 32'h404baa38} /* (9, 13, 12) {real, imag} */,
  {32'hc05dbcec, 32'h401397ea} /* (9, 13, 11) {real, imag} */,
  {32'hbfa2883b, 32'h408943d1} /* (9, 13, 10) {real, imag} */,
  {32'hbe517c30, 32'hbfba4b54} /* (9, 13, 9) {real, imag} */,
  {32'hc041492a, 32'hc08e3f18} /* (9, 13, 8) {real, imag} */,
  {32'hc007e5a1, 32'hbfaae08a} /* (9, 13, 7) {real, imag} */,
  {32'hbe5f5f00, 32'h3f0b41c4} /* (9, 13, 6) {real, imag} */,
  {32'h3f4b9ed4, 32'hc00a68ec} /* (9, 13, 5) {real, imag} */,
  {32'hbf918500, 32'hc06784e4} /* (9, 13, 4) {real, imag} */,
  {32'h3fbf75ce, 32'hbf949fd1} /* (9, 13, 3) {real, imag} */,
  {32'h3f00512e, 32'hc0076cca} /* (9, 13, 2) {real, imag} */,
  {32'hc08c3dda, 32'hc0cd06cc} /* (9, 13, 1) {real, imag} */,
  {32'hbf7ad3d4, 32'hc0475651} /* (9, 13, 0) {real, imag} */,
  {32'hc03e8d7f, 32'hc0278e7c} /* (9, 12, 31) {real, imag} */,
  {32'h3f907d5c, 32'hc0922666} /* (9, 12, 30) {real, imag} */,
  {32'h3f28967e, 32'h3f9f6433} /* (9, 12, 29) {real, imag} */,
  {32'hbfc02615, 32'h3ef933a4} /* (9, 12, 28) {real, imag} */,
  {32'h4014a004, 32'h3f40614e} /* (9, 12, 27) {real, imag} */,
  {32'hbf57bfaa, 32'hc06b94bf} /* (9, 12, 26) {real, imag} */,
  {32'hc01f9959, 32'hc0318b86} /* (9, 12, 25) {real, imag} */,
  {32'hc0261be6, 32'hbe7d5ec0} /* (9, 12, 24) {real, imag} */,
  {32'hc0840f8a, 32'h405cfa00} /* (9, 12, 23) {real, imag} */,
  {32'hc0bfba3a, 32'h4018c1a3} /* (9, 12, 22) {real, imag} */,
  {32'hc0d343d9, 32'h3f880f0c} /* (9, 12, 21) {real, imag} */,
  {32'hc10e7710, 32'h3ebab7d4} /* (9, 12, 20) {real, imag} */,
  {32'hbff08ef6, 32'hc03428be} /* (9, 12, 19) {real, imag} */,
  {32'h3f9ec190, 32'hc01735f9} /* (9, 12, 18) {real, imag} */,
  {32'hbfc14904, 32'h402291da} /* (9, 12, 17) {real, imag} */,
  {32'hc019449f, 32'h4090d874} /* (9, 12, 16) {real, imag} */,
  {32'h3fbb4969, 32'h4052a9b4} /* (9, 12, 15) {real, imag} */,
  {32'hc050527e, 32'hc07602b4} /* (9, 12, 14) {real, imag} */,
  {32'hc0171edb, 32'hc0c4b274} /* (9, 12, 13) {real, imag} */,
  {32'h402c6404, 32'hbf82b0f3} /* (9, 12, 12) {real, imag} */,
  {32'hc02ce888, 32'h3fdc8498} /* (9, 12, 11) {real, imag} */,
  {32'hc0dcb6ba, 32'hbf29ba0e} /* (9, 12, 10) {real, imag} */,
  {32'h3fe373df, 32'hbf779490} /* (9, 12, 9) {real, imag} */,
  {32'h401758f0, 32'h3f45ca48} /* (9, 12, 8) {real, imag} */,
  {32'h40229c35, 32'h3f42ebce} /* (9, 12, 7) {real, imag} */,
  {32'hbf3ca227, 32'h3fc211bd} /* (9, 12, 6) {real, imag} */,
  {32'h4080b8b0, 32'hbf5ea046} /* (9, 12, 5) {real, imag} */,
  {32'h40548073, 32'h3fa1b021} /* (9, 12, 4) {real, imag} */,
  {32'h4068bce4, 32'h40310e6e} /* (9, 12, 3) {real, imag} */,
  {32'h4017f444, 32'h4078cb3b} /* (9, 12, 2) {real, imag} */,
  {32'h3f8b5e4e, 32'h409d9d2e} /* (9, 12, 1) {real, imag} */,
  {32'h3fe40e31, 32'h40652d8e} /* (9, 12, 0) {real, imag} */,
  {32'h404202cc, 32'hc0297ae4} /* (9, 11, 31) {real, imag} */,
  {32'hc0604ee0, 32'hc100eaeb} /* (9, 11, 30) {real, imag} */,
  {32'h4025d6ac, 32'hc0ae2e0d} /* (9, 11, 29) {real, imag} */,
  {32'h410fd32c, 32'hbfe933da} /* (9, 11, 28) {real, imag} */,
  {32'h40e83356, 32'h40a7fab8} /* (9, 11, 27) {real, imag} */,
  {32'hbfd09e0a, 32'h40b67f89} /* (9, 11, 26) {real, imag} */,
  {32'hbfbf0ba3, 32'hbfdb005e} /* (9, 11, 25) {real, imag} */,
  {32'hbfd23cbe, 32'hc1364e7c} /* (9, 11, 24) {real, imag} */,
  {32'hbfe6afac, 32'hc00712e2} /* (9, 11, 23) {real, imag} */,
  {32'hc0ae15ce, 32'h4048bfa2} /* (9, 11, 22) {real, imag} */,
  {32'hc0fcd0b8, 32'h3f9dbb6e} /* (9, 11, 21) {real, imag} */,
  {32'hc0cbc32e, 32'h3ff743cc} /* (9, 11, 20) {real, imag} */,
  {32'h4013db7e, 32'h40ccf548} /* (9, 11, 19) {real, imag} */,
  {32'hbf79c571, 32'hc062fb4a} /* (9, 11, 18) {real, imag} */,
  {32'hbf212d3e, 32'hc0e13243} /* (9, 11, 17) {real, imag} */,
  {32'h40319c0d, 32'hbf80601a} /* (9, 11, 16) {real, imag} */,
  {32'hc03ffe12, 32'hbdc903b8} /* (9, 11, 15) {real, imag} */,
  {32'hc0a5d01f, 32'h3fbc2e51} /* (9, 11, 14) {real, imag} */,
  {32'hc085af3e, 32'h4042d9e1} /* (9, 11, 13) {real, imag} */,
  {32'hc0733eed, 32'h40a08858} /* (9, 11, 12) {real, imag} */,
  {32'hc085909d, 32'h3fad81a5} /* (9, 11, 11) {real, imag} */,
  {32'h3faad6a0, 32'h404b199e} /* (9, 11, 10) {real, imag} */,
  {32'hbf2683b4, 32'h4075ee14} /* (9, 11, 9) {real, imag} */,
  {32'h3f34f318, 32'h40824348} /* (9, 11, 8) {real, imag} */,
  {32'hbff2f510, 32'h405545fa} /* (9, 11, 7) {real, imag} */,
  {32'hc0764d53, 32'hc032d9f5} /* (9, 11, 6) {real, imag} */,
  {32'h4052820a, 32'hbe5f2960} /* (9, 11, 5) {real, imag} */,
  {32'h3ef2c18c, 32'h40240faa} /* (9, 11, 4) {real, imag} */,
  {32'hc0fd098c, 32'hbfc4470a} /* (9, 11, 3) {real, imag} */,
  {32'hc1013702, 32'h3e976c50} /* (9, 11, 2) {real, imag} */,
  {32'hc0f1f4a4, 32'h410c69e4} /* (9, 11, 1) {real, imag} */,
  {32'h3fe910fb, 32'h40f73b06} /* (9, 11, 0) {real, imag} */,
  {32'hbf1c745a, 32'h40bef488} /* (9, 10, 31) {real, imag} */,
  {32'h3f52c5b6, 32'hbf1f6564} /* (9, 10, 30) {real, imag} */,
  {32'h40c568d1, 32'hc0a3abbb} /* (9, 10, 29) {real, imag} */,
  {32'h3fb81766, 32'hc085219e} /* (9, 10, 28) {real, imag} */,
  {32'hc01de940, 32'hc0e543d1} /* (9, 10, 27) {real, imag} */,
  {32'h4054d430, 32'hc01bd826} /* (9, 10, 26) {real, imag} */,
  {32'hc0332e7f, 32'h3fc70701} /* (9, 10, 25) {real, imag} */,
  {32'hbfb1c337, 32'hbefc04b0} /* (9, 10, 24) {real, imag} */,
  {32'hc06f0385, 32'h3fc0d886} /* (9, 10, 23) {real, imag} */,
  {32'hc0e59e10, 32'h40c6977e} /* (9, 10, 22) {real, imag} */,
  {32'hbf4836f8, 32'h410335f0} /* (9, 10, 21) {real, imag} */,
  {32'hbf9df58a, 32'h4104b5ae} /* (9, 10, 20) {real, imag} */,
  {32'hbfec734a, 32'h3fa9b0fc} /* (9, 10, 19) {real, imag} */,
  {32'h40fcc059, 32'h40f1727a} /* (9, 10, 18) {real, imag} */,
  {32'h4098274e, 32'h41035093} /* (9, 10, 17) {real, imag} */,
  {32'hbf9c79ce, 32'h3f34407c} /* (9, 10, 16) {real, imag} */,
  {32'hc09dd13a, 32'hc081917b} /* (9, 10, 15) {real, imag} */,
  {32'hbf0164f8, 32'hc0a9b994} /* (9, 10, 14) {real, imag} */,
  {32'hbfcb3871, 32'hc0c7e4b6} /* (9, 10, 13) {real, imag} */,
  {32'hbf93b1b4, 32'hc0583780} /* (9, 10, 12) {real, imag} */,
  {32'h3d9cfcc0, 32'hc080804a} /* (9, 10, 11) {real, imag} */,
  {32'hc0b018e3, 32'h3d9dfac0} /* (9, 10, 10) {real, imag} */,
  {32'hc0b25ebc, 32'hbf57bc6e} /* (9, 10, 9) {real, imag} */,
  {32'hc00f6f21, 32'h4075211e} /* (9, 10, 8) {real, imag} */,
  {32'h3fad8650, 32'hbb647400} /* (9, 10, 7) {real, imag} */,
  {32'h4054171c, 32'h408e668a} /* (9, 10, 6) {real, imag} */,
  {32'h3f1fe136, 32'hbf9f041a} /* (9, 10, 5) {real, imag} */,
  {32'hc037bdd7, 32'h40d91774} /* (9, 10, 4) {real, imag} */,
  {32'hc105513c, 32'h40047bd2} /* (9, 10, 3) {real, imag} */,
  {32'hc0c87c7b, 32'hc088759b} /* (9, 10, 2) {real, imag} */,
  {32'h3fc6cc31, 32'h3fade9fe} /* (9, 10, 1) {real, imag} */,
  {32'h4084d93c, 32'h3e6cfbd4} /* (9, 10, 0) {real, imag} */,
  {32'hbf992477, 32'h4055a547} /* (9, 9, 31) {real, imag} */,
  {32'hbf55ba72, 32'hbfbf2616} /* (9, 9, 30) {real, imag} */,
  {32'hbe7d27c4, 32'h40b1f358} /* (9, 9, 29) {real, imag} */,
  {32'hc0dc7ed0, 32'h409cba84} /* (9, 9, 28) {real, imag} */,
  {32'hc117e6ad, 32'h405388ff} /* (9, 9, 27) {real, imag} */,
  {32'hc09ff97a, 32'h3fab4cd5} /* (9, 9, 26) {real, imag} */,
  {32'h40b840ee, 32'hc047ab4f} /* (9, 9, 25) {real, imag} */,
  {32'hc05ac194, 32'h3f4e2a90} /* (9, 9, 24) {real, imag} */,
  {32'hc13c41b1, 32'h41110561} /* (9, 9, 23) {real, imag} */,
  {32'hc083be36, 32'h3f8d3fbb} /* (9, 9, 22) {real, imag} */,
  {32'hc1069316, 32'h3e617968} /* (9, 9, 21) {real, imag} */,
  {32'hc0163448, 32'h402cfe7f} /* (9, 9, 20) {real, imag} */,
  {32'h40a280cc, 32'h3fd031c8} /* (9, 9, 19) {real, imag} */,
  {32'h3dae5d30, 32'h3fd94920} /* (9, 9, 18) {real, imag} */,
  {32'h400a28ea, 32'h3edfc248} /* (9, 9, 17) {real, imag} */,
  {32'h40b60fbe, 32'hbfb013f8} /* (9, 9, 16) {real, imag} */,
  {32'h40b73475, 32'hbf2a49b0} /* (9, 9, 15) {real, imag} */,
  {32'h3fe7e428, 32'h40ea439f} /* (9, 9, 14) {real, imag} */,
  {32'hbca16cc0, 32'h40e4c88b} /* (9, 9, 13) {real, imag} */,
  {32'h411608f4, 32'h405f4f5f} /* (9, 9, 12) {real, imag} */,
  {32'h40c263b6, 32'h400a5178} /* (9, 9, 11) {real, imag} */,
  {32'h3fd6c2e4, 32'hbf37271c} /* (9, 9, 10) {real, imag} */,
  {32'h408b6da0, 32'h403bad1e} /* (9, 9, 9) {real, imag} */,
  {32'hc0043db0, 32'h409632a0} /* (9, 9, 8) {real, imag} */,
  {32'hc0ba8b4e, 32'h41057a06} /* (9, 9, 7) {real, imag} */,
  {32'hbf3ae626, 32'h3e8630c0} /* (9, 9, 6) {real, imag} */,
  {32'hc105af36, 32'hbf4157a4} /* (9, 9, 5) {real, imag} */,
  {32'hc14ff71e, 32'hbea80008} /* (9, 9, 4) {real, imag} */,
  {32'hbffded70, 32'h409344c2} /* (9, 9, 3) {real, imag} */,
  {32'h40f65490, 32'h41208890} /* (9, 9, 2) {real, imag} */,
  {32'h400d859d, 32'h3fddb6b6} /* (9, 9, 1) {real, imag} */,
  {32'hc035e106, 32'hc03a2e28} /* (9, 9, 0) {real, imag} */,
  {32'h40c82d04, 32'h406e3592} /* (9, 8, 31) {real, imag} */,
  {32'h410fe3de, 32'h408dadc9} /* (9, 8, 30) {real, imag} */,
  {32'h40a08afe, 32'hc11c7bd9} /* (9, 8, 29) {real, imag} */,
  {32'hbfaf5d9c, 32'hc1a5466c} /* (9, 8, 28) {real, imag} */,
  {32'hbf5dc9fb, 32'hc0ed6a30} /* (9, 8, 27) {real, imag} */,
  {32'h404ccf92, 32'hc08c5b37} /* (9, 8, 26) {real, imag} */,
  {32'h402f7885, 32'hc065f5e4} /* (9, 8, 25) {real, imag} */,
  {32'h407ec56a, 32'h40006176} /* (9, 8, 24) {real, imag} */,
  {32'h41926a1c, 32'hc1229f32} /* (9, 8, 23) {real, imag} */,
  {32'h41867fe6, 32'hc154cd28} /* (9, 8, 22) {real, imag} */,
  {32'h40e90433, 32'hc05c5008} /* (9, 8, 21) {real, imag} */,
  {32'h4072b10c, 32'hbe9ec110} /* (9, 8, 20) {real, imag} */,
  {32'hc02e2b6c, 32'h3f9562d2} /* (9, 8, 19) {real, imag} */,
  {32'hbf316eaf, 32'h40413e43} /* (9, 8, 18) {real, imag} */,
  {32'hc058ddf9, 32'h404a9496} /* (9, 8, 17) {real, imag} */,
  {32'h412a394b, 32'h403e33f8} /* (9, 8, 16) {real, imag} */,
  {32'h413cff62, 32'h40c68228} /* (9, 8, 15) {real, imag} */,
  {32'h40ac68fc, 32'h3e898a54} /* (9, 8, 14) {real, imag} */,
  {32'h3fc012dc, 32'hbfaeab38} /* (9, 8, 13) {real, imag} */,
  {32'h4046ca9a, 32'h4080dac7} /* (9, 8, 12) {real, imag} */,
  {32'h41293f46, 32'h4032bdd5} /* (9, 8, 11) {real, imag} */,
  {32'h40cf3cd6, 32'h40c907f7} /* (9, 8, 10) {real, imag} */,
  {32'h3ee52448, 32'h410c101d} /* (9, 8, 9) {real, imag} */,
  {32'hbf5ad8bc, 32'h3fae01ce} /* (9, 8, 8) {real, imag} */,
  {32'h40db068f, 32'hbff787bc} /* (9, 8, 7) {real, imag} */,
  {32'h40b0afad, 32'hbdd72a00} /* (9, 8, 6) {real, imag} */,
  {32'h41221528, 32'h41323e84} /* (9, 8, 5) {real, imag} */,
  {32'h4117721f, 32'h407ffd52} /* (9, 8, 4) {real, imag} */,
  {32'h40a30ab9, 32'h408c9ca8} /* (9, 8, 3) {real, imag} */,
  {32'hbf2a233c, 32'hbf6b222e} /* (9, 8, 2) {real, imag} */,
  {32'h40815afa, 32'hc064280a} /* (9, 8, 1) {real, imag} */,
  {32'h3f8148cc, 32'hc0341b36} /* (9, 8, 0) {real, imag} */,
  {32'h3f8a5466, 32'h40289d81} /* (9, 7, 31) {real, imag} */,
  {32'hbf84bb47, 32'h41472527} /* (9, 7, 30) {real, imag} */,
  {32'hc00ab70e, 32'h413f0c6c} /* (9, 7, 29) {real, imag} */,
  {32'hc1976835, 32'h402a44fd} /* (9, 7, 28) {real, imag} */,
  {32'hc1244e7c, 32'hc08564d3} /* (9, 7, 27) {real, imag} */,
  {32'h4062f10b, 32'hc10bedd5} /* (9, 7, 26) {real, imag} */,
  {32'hbf25a3f8, 32'hbfe6bd4c} /* (9, 7, 25) {real, imag} */,
  {32'hc118f585, 32'h404ce628} /* (9, 7, 24) {real, imag} */,
  {32'hc12940b1, 32'h409a114c} /* (9, 7, 23) {real, imag} */,
  {32'hc107a519, 32'h41093d22} /* (9, 7, 22) {real, imag} */,
  {32'h407027f3, 32'h4090965b} /* (9, 7, 21) {real, imag} */,
  {32'hbfbec844, 32'hc0849aec} /* (9, 7, 20) {real, imag} */,
  {32'hc0bbfaf5, 32'hc1423b86} /* (9, 7, 19) {real, imag} */,
  {32'h41036d31, 32'h40109904} /* (9, 7, 18) {real, imag} */,
  {32'h408cb4d8, 32'h41015e85} /* (9, 7, 17) {real, imag} */,
  {32'hbf4dec42, 32'h3f03405a} /* (9, 7, 16) {real, imag} */,
  {32'hc0629bb4, 32'h413ca7ee} /* (9, 7, 15) {real, imag} */,
  {32'h3fd6aca4, 32'h4165f60a} /* (9, 7, 14) {real, imag} */,
  {32'hc0909364, 32'h41931cb8} /* (9, 7, 13) {real, imag} */,
  {32'hc160c9d9, 32'h40c12f4c} /* (9, 7, 12) {real, imag} */,
  {32'hc0a38c44, 32'hc0bf83d5} /* (9, 7, 11) {real, imag} */,
  {32'h4095eee7, 32'h40f5dac9} /* (9, 7, 10) {real, imag} */,
  {32'h40c5003a, 32'h3fd73b70} /* (9, 7, 9) {real, imag} */,
  {32'h3f8c3cb4, 32'hc02423a9} /* (9, 7, 8) {real, imag} */,
  {32'h40e4c3b6, 32'hbf12edd6} /* (9, 7, 7) {real, imag} */,
  {32'h40e17361, 32'hbff52a22} /* (9, 7, 6) {real, imag} */,
  {32'h411e1955, 32'hbe3cac30} /* (9, 7, 5) {real, imag} */,
  {32'hbfabbf22, 32'hc0f4460a} /* (9, 7, 4) {real, imag} */,
  {32'hc0b8d53c, 32'hc0c27456} /* (9, 7, 3) {real, imag} */,
  {32'h4024eade, 32'h3f76dba0} /* (9, 7, 2) {real, imag} */,
  {32'hc1003c5e, 32'hc0f9f986} /* (9, 7, 1) {real, imag} */,
  {32'hc1494644, 32'hc077e543} /* (9, 7, 0) {real, imag} */,
  {32'hc0eef87d, 32'h40a20d74} /* (9, 6, 31) {real, imag} */,
  {32'hbfa7c31c, 32'h4131df98} /* (9, 6, 30) {real, imag} */,
  {32'h4133ff1e, 32'h3e806318} /* (9, 6, 29) {real, imag} */,
  {32'h415d1464, 32'h3f9aac96} /* (9, 6, 28) {real, imag} */,
  {32'h40459191, 32'hbf09dd9e} /* (9, 6, 27) {real, imag} */,
  {32'hc134fa24, 32'hc10de181} /* (9, 6, 26) {real, imag} */,
  {32'hc125977f, 32'h3ed24b0c} /* (9, 6, 25) {real, imag} */,
  {32'hc08b056e, 32'hc0d7e419} /* (9, 6, 24) {real, imag} */,
  {32'hc105fce7, 32'hc13e4f1c} /* (9, 6, 23) {real, imag} */,
  {32'hc02852d2, 32'hc07ee9d4} /* (9, 6, 22) {real, imag} */,
  {32'hc1172bd4, 32'h4077f9ec} /* (9, 6, 21) {real, imag} */,
  {32'hc15e26f5, 32'h40833182} /* (9, 6, 20) {real, imag} */,
  {32'hc1017a38, 32'h40945c3c} /* (9, 6, 19) {real, imag} */,
  {32'hbfd347b0, 32'hbf561790} /* (9, 6, 18) {real, imag} */,
  {32'hbf886968, 32'h4097cfb4} /* (9, 6, 17) {real, imag} */,
  {32'hc1066f14, 32'h4115c802} /* (9, 6, 16) {real, imag} */,
  {32'hc13c0712, 32'h3eca33a0} /* (9, 6, 15) {real, imag} */,
  {32'hc12723d7, 32'h41114c89} /* (9, 6, 14) {real, imag} */,
  {32'hbf5f2d38, 32'h40d57d6a} /* (9, 6, 13) {real, imag} */,
  {32'h4076b39e, 32'h3d95e6d0} /* (9, 6, 12) {real, imag} */,
  {32'h3d9b0fc0, 32'h4123cce1} /* (9, 6, 11) {real, imag} */,
  {32'hc01e04ee, 32'h3fb4a3d5} /* (9, 6, 10) {real, imag} */,
  {32'hc153496a, 32'hc1050b18} /* (9, 6, 9) {real, imag} */,
  {32'hc0f34ff4, 32'hc16f4120} /* (9, 6, 8) {real, imag} */,
  {32'hc113c5f1, 32'hc12082da} /* (9, 6, 7) {real, imag} */,
  {32'hc083fa2c, 32'hc075f21a} /* (9, 6, 6) {real, imag} */,
  {32'hc0d4f4ea, 32'h402be704} /* (9, 6, 5) {real, imag} */,
  {32'h40032a38, 32'h40237461} /* (9, 6, 4) {real, imag} */,
  {32'h4032ec2e, 32'h40399398} /* (9, 6, 3) {real, imag} */,
  {32'hbffc348c, 32'hc017aee6} /* (9, 6, 2) {real, imag} */,
  {32'h4115e44c, 32'hbfbc5e62} /* (9, 6, 1) {real, imag} */,
  {32'h411043c8, 32'h404a9890} /* (9, 6, 0) {real, imag} */,
  {32'hc061c053, 32'hc0622e24} /* (9, 5, 31) {real, imag} */,
  {32'h409af520, 32'hc01f24da} /* (9, 5, 30) {real, imag} */,
  {32'h3e1072d8, 32'hc0cc6f70} /* (9, 5, 29) {real, imag} */,
  {32'h408dc626, 32'hc181b488} /* (9, 5, 28) {real, imag} */,
  {32'h414ce4d4, 32'hc0df008d} /* (9, 5, 27) {real, imag} */,
  {32'hc04edb06, 32'hbf8bb588} /* (9, 5, 26) {real, imag} */,
  {32'h3f8a2e88, 32'hc00b658e} /* (9, 5, 25) {real, imag} */,
  {32'h40e68ee8, 32'hc0f67050} /* (9, 5, 24) {real, imag} */,
  {32'hbe009b00, 32'hc0fe92eb} /* (9, 5, 23) {real, imag} */,
  {32'h40e50182, 32'h4056a8f2} /* (9, 5, 22) {real, imag} */,
  {32'hbf8d3fcc, 32'hc052c464} /* (9, 5, 21) {real, imag} */,
  {32'h40362dfa, 32'hbf3993f0} /* (9, 5, 20) {real, imag} */,
  {32'h415b0857, 32'h412a751e} /* (9, 5, 19) {real, imag} */,
  {32'h40dd78ec, 32'h3e2bb680} /* (9, 5, 18) {real, imag} */,
  {32'hc091242c, 32'hc142b873} /* (9, 5, 17) {real, imag} */,
  {32'hc02fcadb, 32'h40b1605a} /* (9, 5, 16) {real, imag} */,
  {32'h410e9264, 32'h408e76c0} /* (9, 5, 15) {real, imag} */,
  {32'h4005caf0, 32'h41109d4f} /* (9, 5, 14) {real, imag} */,
  {32'h3eda71f0, 32'hbfe56d3a} /* (9, 5, 13) {real, imag} */,
  {32'hc139fe01, 32'hc172ace7} /* (9, 5, 12) {real, imag} */,
  {32'hc173bc30, 32'hc1443290} /* (9, 5, 11) {real, imag} */,
  {32'hc0755e5a, 32'hc0ce894a} /* (9, 5, 10) {real, imag} */,
  {32'hc0101e8d, 32'h408e9f86} /* (9, 5, 9) {real, imag} */,
  {32'h3f1de658, 32'hbf39e7f0} /* (9, 5, 8) {real, imag} */,
  {32'h41a9be26, 32'hc005f056} /* (9, 5, 7) {real, imag} */,
  {32'h41434ef7, 32'h4105cea5} /* (9, 5, 6) {real, imag} */,
  {32'h41077c86, 32'h414d5fbe} /* (9, 5, 5) {real, imag} */,
  {32'h40a7bdd6, 32'hbf5e22b9} /* (9, 5, 4) {real, imag} */,
  {32'h400536e2, 32'hc126f18c} /* (9, 5, 3) {real, imag} */,
  {32'hbff2bea4, 32'hbfebae9c} /* (9, 5, 2) {real, imag} */,
  {32'hc07a385c, 32'hbfce7e1b} /* (9, 5, 1) {real, imag} */,
  {32'h406ebb2e, 32'hc1769b06} /* (9, 5, 0) {real, imag} */,
  {32'hc01ca794, 32'h40e24aa6} /* (9, 4, 31) {real, imag} */,
  {32'h3f29d508, 32'h411fed1e} /* (9, 4, 30) {real, imag} */,
  {32'h408e4e3f, 32'hc11f09c6} /* (9, 4, 29) {real, imag} */,
  {32'h40ac475b, 32'hc13c1cf5} /* (9, 4, 28) {real, imag} */,
  {32'h40771626, 32'h410e55af} /* (9, 4, 27) {real, imag} */,
  {32'hc1368fa2, 32'h412c6e1e} /* (9, 4, 26) {real, imag} */,
  {32'hc0d15b62, 32'h40b09036} /* (9, 4, 25) {real, imag} */,
  {32'h4040279f, 32'hbfb8e170} /* (9, 4, 24) {real, imag} */,
  {32'h41293885, 32'hc0448899} /* (9, 4, 23) {real, imag} */,
  {32'h40b5d816, 32'h4111b50d} /* (9, 4, 22) {real, imag} */,
  {32'h3fb69b12, 32'h416c7621} /* (9, 4, 21) {real, imag} */,
  {32'hc05e43bd, 32'h40756164} /* (9, 4, 20) {real, imag} */,
  {32'hc13f749c, 32'hc1310d5c} /* (9, 4, 19) {real, imag} */,
  {32'hc0b369f8, 32'hc1452faa} /* (9, 4, 18) {real, imag} */,
  {32'hc0b1eb32, 32'hc1210bc2} /* (9, 4, 17) {real, imag} */,
  {32'hc1298c4b, 32'hc0f86870} /* (9, 4, 16) {real, imag} */,
  {32'h3f97354e, 32'h4021dbac} /* (9, 4, 15) {real, imag} */,
  {32'h41b3d1d6, 32'h400eccc1} /* (9, 4, 14) {real, imag} */,
  {32'h406a9ab1, 32'h40ab8a3e} /* (9, 4, 13) {real, imag} */,
  {32'hc0a8d120, 32'h40258bd6} /* (9, 4, 12) {real, imag} */,
  {32'hc0db3a56, 32'h3d769c80} /* (9, 4, 11) {real, imag} */,
  {32'h40ba228f, 32'h3ea430f0} /* (9, 4, 10) {real, imag} */,
  {32'h415c47b5, 32'hc0f8782d} /* (9, 4, 9) {real, imag} */,
  {32'hc04f4208, 32'h405b20ac} /* (9, 4, 8) {real, imag} */,
  {32'hc16778b2, 32'h3e08aee0} /* (9, 4, 7) {real, imag} */,
  {32'hc0e2ce79, 32'hc13a8604} /* (9, 4, 6) {real, imag} */,
  {32'hc08e8d6a, 32'h3f52e218} /* (9, 4, 5) {real, imag} */,
  {32'hc121dad1, 32'h40d9c58b} /* (9, 4, 4) {real, imag} */,
  {32'h4106b681, 32'hc1198e23} /* (9, 4, 3) {real, imag} */,
  {32'h40f99c36, 32'hc09c24a8} /* (9, 4, 2) {real, imag} */,
  {32'h41326c8e, 32'h410442ce} /* (9, 4, 1) {real, imag} */,
  {32'h409d70ad, 32'h415067de} /* (9, 4, 0) {real, imag} */,
  {32'h40d1cf94, 32'hc08a8ca2} /* (9, 3, 31) {real, imag} */,
  {32'hc0c4e402, 32'hbf79984e} /* (9, 3, 30) {real, imag} */,
  {32'hc1786f35, 32'hbe28f1c0} /* (9, 3, 29) {real, imag} */,
  {32'hc0e58f1e, 32'hc01b8763} /* (9, 3, 28) {real, imag} */,
  {32'hc0087e82, 32'h3f77b088} /* (9, 3, 27) {real, imag} */,
  {32'hc123a908, 32'h40d1e9fd} /* (9, 3, 26) {real, imag} */,
  {32'hbf4a4abc, 32'h3f8717a4} /* (9, 3, 25) {real, imag} */,
  {32'h409bb579, 32'h40e1779b} /* (9, 3, 24) {real, imag} */,
  {32'h41165d16, 32'h415da70e} /* (9, 3, 23) {real, imag} */,
  {32'h41638c9b, 32'hc08bdea6} /* (9, 3, 22) {real, imag} */,
  {32'h4180c9ac, 32'hc0e9d104} /* (9, 3, 21) {real, imag} */,
  {32'h4199d65d, 32'hc0ddcc13} /* (9, 3, 20) {real, imag} */,
  {32'h406cfd1f, 32'hbd16d600} /* (9, 3, 19) {real, imag} */,
  {32'hc1016940, 32'hbfdf2c17} /* (9, 3, 18) {real, imag} */,
  {32'h4026ec58, 32'h3ece1a40} /* (9, 3, 17) {real, imag} */,
  {32'hc10c3b38, 32'hc07f451c} /* (9, 3, 16) {real, imag} */,
  {32'hc0dae0bd, 32'hc130a6ef} /* (9, 3, 15) {real, imag} */,
  {32'hc0a75550, 32'h40febc80} /* (9, 3, 14) {real, imag} */,
  {32'h40ab0c5c, 32'h41168f32} /* (9, 3, 13) {real, imag} */,
  {32'h4075aa7c, 32'h3e4bbbe0} /* (9, 3, 12) {real, imag} */,
  {32'h40fd73a6, 32'hc1180ca5} /* (9, 3, 11) {real, imag} */,
  {32'h406de0d0, 32'hc1069c08} /* (9, 3, 10) {real, imag} */,
  {32'hc0a0cd2a, 32'h418186c5} /* (9, 3, 9) {real, imag} */,
  {32'h414e57c2, 32'h419b80e4} /* (9, 3, 8) {real, imag} */,
  {32'h3f17c9c8, 32'h3ff3c120} /* (9, 3, 7) {real, imag} */,
  {32'h416cc88d, 32'hbfbc8af0} /* (9, 3, 6) {real, imag} */,
  {32'h413d4e54, 32'hc1377717} /* (9, 3, 5) {real, imag} */,
  {32'hc0181172, 32'hc03ca85b} /* (9, 3, 4) {real, imag} */,
  {32'h405f6c0b, 32'hc10e6aaa} /* (9, 3, 3) {real, imag} */,
  {32'h40cf904f, 32'hc0844950} /* (9, 3, 2) {real, imag} */,
  {32'h410643ae, 32'hc0472ab0} /* (9, 3, 1) {real, imag} */,
  {32'h410f1f48, 32'hc09a0441} /* (9, 3, 0) {real, imag} */,
  {32'hc0bce66c, 32'hc0d8916f} /* (9, 2, 31) {real, imag} */,
  {32'h40277c26, 32'hc1304757} /* (9, 2, 30) {real, imag} */,
  {32'h40e01d0e, 32'hc168902f} /* (9, 2, 29) {real, imag} */,
  {32'h41a47e15, 32'hbff553c6} /* (9, 2, 28) {real, imag} */,
  {32'h4165d33d, 32'hc1815224} /* (9, 2, 27) {real, imag} */,
  {32'h41307932, 32'hc1746ba3} /* (9, 2, 26) {real, imag} */,
  {32'hc0e262fc, 32'hc1a82618} /* (9, 2, 25) {real, imag} */,
  {32'hc1747dec, 32'hc1e06ac6} /* (9, 2, 24) {real, imag} */,
  {32'h402c2f23, 32'hc11dc171} /* (9, 2, 23) {real, imag} */,
  {32'hc06c637c, 32'hc0d59eb1} /* (9, 2, 22) {real, imag} */,
  {32'hc0ede350, 32'hc1134662} /* (9, 2, 21) {real, imag} */,
  {32'hc184b62e, 32'h414ebb5c} /* (9, 2, 20) {real, imag} */,
  {32'h404615fa, 32'h4191c054} /* (9, 2, 19) {real, imag} */,
  {32'h40866878, 32'h40e8af7b} /* (9, 2, 18) {real, imag} */,
  {32'hc0d69fbe, 32'h4105885a} /* (9, 2, 17) {real, imag} */,
  {32'h4119e832, 32'h4112f74a} /* (9, 2, 16) {real, imag} */,
  {32'h404d6306, 32'h40b9ead5} /* (9, 2, 15) {real, imag} */,
  {32'hbfee514c, 32'h3ec730c8} /* (9, 2, 14) {real, imag} */,
  {32'hc0c39956, 32'h40d87095} /* (9, 2, 13) {real, imag} */,
  {32'hc16e655d, 32'h412ce6aa} /* (9, 2, 12) {real, imag} */,
  {32'hc1187c64, 32'h417265a7} /* (9, 2, 11) {real, imag} */,
  {32'h410a3c56, 32'hbefc07e6} /* (9, 2, 10) {real, imag} */,
  {32'h403b781c, 32'hc177f134} /* (9, 2, 9) {real, imag} */,
  {32'hc0cd8bac, 32'hc2052b86} /* (9, 2, 8) {real, imag} */,
  {32'h4043b7c2, 32'hc1d3daab} /* (9, 2, 7) {real, imag} */,
  {32'h4188ce7e, 32'hc157f359} /* (9, 2, 6) {real, imag} */,
  {32'h40f9f60a, 32'h3f9464bc} /* (9, 2, 5) {real, imag} */,
  {32'h404542ec, 32'hbe344d00} /* (9, 2, 4) {real, imag} */,
  {32'h3e72a004, 32'h4090467a} /* (9, 2, 3) {real, imag} */,
  {32'hbee3897c, 32'h40da7628} /* (9, 2, 2) {real, imag} */,
  {32'h3da6c110, 32'h406841e4} /* (9, 2, 1) {real, imag} */,
  {32'h4076632a, 32'h403c6936} /* (9, 2, 0) {real, imag} */,
  {32'hc0313c12, 32'hc1038813} /* (9, 1, 31) {real, imag} */,
  {32'hc18ca618, 32'hc1ccef3a} /* (9, 1, 30) {real, imag} */,
  {32'hc1d186dc, 32'hbfab3c14} /* (9, 1, 29) {real, imag} */,
  {32'hc11418fd, 32'h4194b3fa} /* (9, 1, 28) {real, imag} */,
  {32'hc14a740e, 32'h41317c87} /* (9, 1, 27) {real, imag} */,
  {32'hc1788a29, 32'h407fb8fc} /* (9, 1, 26) {real, imag} */,
  {32'hc1649fae, 32'h4108572e} /* (9, 1, 25) {real, imag} */,
  {32'hc10ec958, 32'h416183fe} /* (9, 1, 24) {real, imag} */,
  {32'hc0778505, 32'h41473f13} /* (9, 1, 23) {real, imag} */,
  {32'hc0b82fa7, 32'h3f2b05a0} /* (9, 1, 22) {real, imag} */,
  {32'hc14f3236, 32'hc12e4435} /* (9, 1, 21) {real, imag} */,
  {32'hc0d216b2, 32'hc1333916} /* (9, 1, 20) {real, imag} */,
  {32'hc06ed5d4, 32'h3fa869b8} /* (9, 1, 19) {real, imag} */,
  {32'h4048a794, 32'hc0ce975e} /* (9, 1, 18) {real, imag} */,
  {32'hbfa78718, 32'hc09f396a} /* (9, 1, 17) {real, imag} */,
  {32'hc031761a, 32'hbf0909e0} /* (9, 1, 16) {real, imag} */,
  {32'h417adde6, 32'h3e8240b8} /* (9, 1, 15) {real, imag} */,
  {32'h417bbec6, 32'hc1346481} /* (9, 1, 14) {real, imag} */,
  {32'h4182ae9e, 32'hc195ab4a} /* (9, 1, 13) {real, imag} */,
  {32'h41519064, 32'hc186f5f7} /* (9, 1, 12) {real, imag} */,
  {32'hbe56ef40, 32'hc0e68ade} /* (9, 1, 11) {real, imag} */,
  {32'hc1234931, 32'hc1b5451e} /* (9, 1, 10) {real, imag} */,
  {32'hc1a52840, 32'hc0c5b639} /* (9, 1, 9) {real, imag} */,
  {32'hc196496f, 32'h40942218} /* (9, 1, 8) {real, imag} */,
  {32'h3f5f7ad8, 32'h411e9dda} /* (9, 1, 7) {real, imag} */,
  {32'hbfed1db8, 32'h4185001d} /* (9, 1, 6) {real, imag} */,
  {32'hc193e643, 32'h408cf9a2} /* (9, 1, 5) {real, imag} */,
  {32'hc12134b5, 32'hbfb69c0c} /* (9, 1, 4) {real, imag} */,
  {32'h4115ec2a, 32'hc0ed4ace} /* (9, 1, 3) {real, imag} */,
  {32'h413251b5, 32'hc0cad6ef} /* (9, 1, 2) {real, imag} */,
  {32'hc075e1cc, 32'hc0075d6c} /* (9, 1, 1) {real, imag} */,
  {32'hc080dc35, 32'hc0780294} /* (9, 1, 0) {real, imag} */,
  {32'h3f9ecd4e, 32'h40dc2f03} /* (9, 0, 31) {real, imag} */,
  {32'hc15aed32, 32'h3fba3aca} /* (9, 0, 30) {real, imag} */,
  {32'hc167dda5, 32'h41121fc6} /* (9, 0, 29) {real, imag} */,
  {32'hc101bb94, 32'h412c76f5} /* (9, 0, 28) {real, imag} */,
  {32'hc0997786, 32'h4070f747} /* (9, 0, 27) {real, imag} */,
  {32'hc15d2f4a, 32'h407a918a} /* (9, 0, 26) {real, imag} */,
  {32'hc13808cc, 32'h4182e540} /* (9, 0, 25) {real, imag} */,
  {32'hbf77322e, 32'h41a7d3b6} /* (9, 0, 24) {real, imag} */,
  {32'hc000e8ec, 32'h417fc7c2} /* (9, 0, 23) {real, imag} */,
  {32'h3ffcdbb6, 32'h4197d01b} /* (9, 0, 22) {real, imag} */,
  {32'hc0d0edee, 32'h41085f3d} /* (9, 0, 21) {real, imag} */,
  {32'h3eb9fcce, 32'hc1707be2} /* (9, 0, 20) {real, imag} */,
  {32'h41193eb6, 32'hc0afd1e3} /* (9, 0, 19) {real, imag} */,
  {32'h40a2d21c, 32'hc109f2aa} /* (9, 0, 18) {real, imag} */,
  {32'hc13f60e2, 32'h3fbf3f64} /* (9, 0, 17) {real, imag} */,
  {32'hbfb897e0, 32'h410c1f7a} /* (9, 0, 16) {real, imag} */,
  {32'h40eda110, 32'h409bb642} /* (9, 0, 15) {real, imag} */,
  {32'h40d6a2c0, 32'h413abb68} /* (9, 0, 14) {real, imag} */,
  {32'h4171c1dc, 32'h41ae20df} /* (9, 0, 13) {real, imag} */,
  {32'h417ff84d, 32'h4184171c} /* (9, 0, 12) {real, imag} */,
  {32'h412f84b7, 32'hc1260c10} /* (9, 0, 11) {real, imag} */,
  {32'h4025f914, 32'hc0e7a574} /* (9, 0, 10) {real, imag} */,
  {32'hc0896b38, 32'h41664119} /* (9, 0, 9) {real, imag} */,
  {32'h40323404, 32'h401969cc} /* (9, 0, 8) {real, imag} */,
  {32'h41ac2df0, 32'hc0983320} /* (9, 0, 7) {real, imag} */,
  {32'h40df1228, 32'hbfd3dd9b} /* (9, 0, 6) {real, imag} */,
  {32'hc18378ef, 32'h4156721d} /* (9, 0, 5) {real, imag} */,
  {32'hc0e3db82, 32'h4082c63c} /* (9, 0, 4) {real, imag} */,
  {32'h40a4d5f6, 32'h40492d66} /* (9, 0, 3) {real, imag} */,
  {32'hbf85290d, 32'h411f7a11} /* (9, 0, 2) {real, imag} */,
  {32'hc1525ff0, 32'h41107a3a} /* (9, 0, 1) {real, imag} */,
  {32'hc036bd5f, 32'h40e1cf4a} /* (9, 0, 0) {real, imag} */,
  {32'hc0b73c8a, 32'h414660a7} /* (8, 31, 31) {real, imag} */,
  {32'hc1236d0d, 32'h420b36b4} /* (8, 31, 30) {real, imag} */,
  {32'hc19bfbf1, 32'h42243d14} /* (8, 31, 29) {real, imag} */,
  {32'hc1bf8be7, 32'h420dca63} /* (8, 31, 28) {real, imag} */,
  {32'hc1c89e92, 32'h41eb3c58} /* (8, 31, 27) {real, imag} */,
  {32'hc19423ad, 32'h41d6f862} /* (8, 31, 26) {real, imag} */,
  {32'hc1d7a014, 32'h42297f28} /* (8, 31, 25) {real, imag} */,
  {32'hc20527f5, 32'h41faf346} /* (8, 31, 24) {real, imag} */,
  {32'hc0b77598, 32'h42375fee} /* (8, 31, 23) {real, imag} */,
  {32'hc18d457d, 32'h42194913} /* (8, 31, 22) {real, imag} */,
  {32'hc21bfd24, 32'h4170a14e} /* (8, 31, 21) {real, imag} */,
  {32'hc18fbb23, 32'hc10bb559} /* (8, 31, 20) {real, imag} */,
  {32'hc0ece4a8, 32'hc1341da6} /* (8, 31, 19) {real, imag} */,
  {32'hc1352539, 32'hc2075694} /* (8, 31, 18) {real, imag} */,
  {32'hc0970aac, 32'hc21f833d} /* (8, 31, 17) {real, imag} */,
  {32'h40d35de0, 32'hc1a02f98} /* (8, 31, 16) {real, imag} */,
  {32'h41ea5ad2, 32'hc205047d} /* (8, 31, 15) {real, imag} */,
  {32'h41e68607, 32'hc207c8e4} /* (8, 31, 14) {real, imag} */,
  {32'h420c9172, 32'hc226aac9} /* (8, 31, 13) {real, imag} */,
  {32'h4151d07e, 32'hc1d22605} /* (8, 31, 12) {real, imag} */,
  {32'h418c6828, 32'hc18687e8} /* (8, 31, 11) {real, imag} */,
  {32'h4057ffdc, 32'h4186c7ee} /* (8, 31, 10) {real, imag} */,
  {32'h3fbd17a8, 32'h4209ad76} /* (8, 31, 9) {real, imag} */,
  {32'h41121e02, 32'h41f65d50} /* (8, 31, 8) {real, imag} */,
  {32'h40f3628e, 32'h4194dabc} /* (8, 31, 7) {real, imag} */,
  {32'hc0b79f6b, 32'h4228042f} /* (8, 31, 6) {real, imag} */,
  {32'hc1a0ee13, 32'h424cb546} /* (8, 31, 5) {real, imag} */,
  {32'hc1bdcee0, 32'h422feab9} /* (8, 31, 4) {real, imag} */,
  {32'hc1d528a0, 32'h421bda66} /* (8, 31, 3) {real, imag} */,
  {32'hc1850802, 32'h4234c4ec} /* (8, 31, 2) {real, imag} */,
  {32'hc19ba1d6, 32'h41f3018d} /* (8, 31, 1) {real, imag} */,
  {32'hc13b97a2, 32'h416fb0c4} /* (8, 31, 0) {real, imag} */,
  {32'hc0a38964, 32'hbf684348} /* (8, 30, 31) {real, imag} */,
  {32'hc0e60ea4, 32'hc1312d6b} /* (8, 30, 30) {real, imag} */,
  {32'h401ecf40, 32'hc1a1578e} /* (8, 30, 29) {real, imag} */,
  {32'hc1536672, 32'hc1bdaef1} /* (8, 30, 28) {real, imag} */,
  {32'hc0a693a6, 32'hc1cf44da} /* (8, 30, 27) {real, imag} */,
  {32'h3f11cfd0, 32'hc203482f} /* (8, 30, 26) {real, imag} */,
  {32'hc0bac26e, 32'hc1d96ff2} /* (8, 30, 25) {real, imag} */,
  {32'h40f26906, 32'hc100355f} /* (8, 30, 24) {real, imag} */,
  {32'h419787bc, 32'hbfbf1128} /* (8, 30, 23) {real, imag} */,
  {32'h41c27357, 32'hc1e31c6e} /* (8, 30, 22) {real, imag} */,
  {32'h412a9db1, 32'hc1b29c0f} /* (8, 30, 21) {real, imag} */,
  {32'hc18d875c, 32'h411b4a68} /* (8, 30, 20) {real, imag} */,
  {32'hc21a42df, 32'h41f0c1a5} /* (8, 30, 19) {real, imag} */,
  {32'hc1e02b38, 32'h41cf69ac} /* (8, 30, 18) {real, imag} */,
  {32'hc210a5d1, 32'h418d9966} /* (8, 30, 17) {real, imag} */,
  {32'hc20265d6, 32'h418db5d7} /* (8, 30, 16) {real, imag} */,
  {32'hc1b0a159, 32'h4151e0f2} /* (8, 30, 15) {real, imag} */,
  {32'hc1b9cfda, 32'h40fb9291} /* (8, 30, 14) {real, imag} */,
  {32'hc1934ceb, 32'h4198f286} /* (8, 30, 13) {real, imag} */,
  {32'hc1538529, 32'h41262d6f} /* (8, 30, 12) {real, imag} */,
  {32'hbfbed124, 32'hc09f12e9} /* (8, 30, 11) {real, imag} */,
  {32'h41de84c3, 32'hc1b01c37} /* (8, 30, 10) {real, imag} */,
  {32'h41fa47ea, 32'hc21a7762} /* (8, 30, 9) {real, imag} */,
  {32'h42024e63, 32'hc1ddf2e2} /* (8, 30, 8) {real, imag} */,
  {32'h4230021b, 32'hc155e664} /* (8, 30, 7) {real, imag} */,
  {32'h4234e0f8, 32'hc1a9e560} /* (8, 30, 6) {real, imag} */,
  {32'h4214a0c5, 32'hc17cb7b0} /* (8, 30, 5) {real, imag} */,
  {32'h41539b4b, 32'hc1a20939} /* (8, 30, 4) {real, imag} */,
  {32'h418e947f, 32'hc1a0870e} /* (8, 30, 3) {real, imag} */,
  {32'h422c7dfe, 32'hc1cd44a6} /* (8, 30, 2) {real, imag} */,
  {32'h41d1526d, 32'hc1940a50} /* (8, 30, 1) {real, imag} */,
  {32'h41339175, 32'h3ec99180} /* (8, 30, 0) {real, imag} */,
  {32'h41374f42, 32'h3e9ac040} /* (8, 29, 31) {real, imag} */,
  {32'h4099d2b0, 32'h3e4c5240} /* (8, 29, 30) {real, imag} */,
  {32'h41022ee6, 32'h401b4de0} /* (8, 29, 29) {real, imag} */,
  {32'hbfad3b5e, 32'h406c5d2a} /* (8, 29, 28) {real, imag} */,
  {32'hc143d146, 32'h4179040f} /* (8, 29, 27) {real, imag} */,
  {32'h41339803, 32'h40aa2c0c} /* (8, 29, 26) {real, imag} */,
  {32'h4173a452, 32'hc0b9a710} /* (8, 29, 25) {real, imag} */,
  {32'h4021db54, 32'hc1b0c090} /* (8, 29, 24) {real, imag} */,
  {32'h40319a08, 32'h3f0b7470} /* (8, 29, 23) {real, imag} */,
  {32'h40fcd790, 32'hc14a9546} /* (8, 29, 22) {real, imag} */,
  {32'h410e19a4, 32'hc1ba9e12} /* (8, 29, 21) {real, imag} */,
  {32'hc0b6d3ae, 32'hc0a688bc} /* (8, 29, 20) {real, imag} */,
  {32'hc12aca53, 32'hc108a7c0} /* (8, 29, 19) {real, imag} */,
  {32'hc1e58c75, 32'h40fbf034} /* (8, 29, 18) {real, imag} */,
  {32'hc17e4973, 32'h413a53fe} /* (8, 29, 17) {real, imag} */,
  {32'h3fa4a0b8, 32'h4136ccd9} /* (8, 29, 16) {real, imag} */,
  {32'h40fe830c, 32'h402a2820} /* (8, 29, 15) {real, imag} */,
  {32'h4112c36a, 32'h404ebe32} /* (8, 29, 14) {real, imag} */,
  {32'h41262faa, 32'hc14571f1} /* (8, 29, 13) {real, imag} */,
  {32'h3f8656a3, 32'hc0eb7450} /* (8, 29, 12) {real, imag} */,
  {32'hc009881e, 32'hc072a17b} /* (8, 29, 11) {real, imag} */,
  {32'h3cbc7b80, 32'hc10f9cb0} /* (8, 29, 10) {real, imag} */,
  {32'h3f66c9f0, 32'h404e3a1e} /* (8, 29, 9) {real, imag} */,
  {32'h40df8048, 32'h411e0046} /* (8, 29, 8) {real, imag} */,
  {32'h41797b86, 32'h41f29fb8} /* (8, 29, 7) {real, imag} */,
  {32'h4159517c, 32'h41e93f0d} /* (8, 29, 6) {real, imag} */,
  {32'h40740ec8, 32'h41034088} /* (8, 29, 5) {real, imag} */,
  {32'h4083e1a6, 32'hc05e41b9} /* (8, 29, 4) {real, imag} */,
  {32'hc134521d, 32'hc0a444a5} /* (8, 29, 3) {real, imag} */,
  {32'hc0a1c9cc, 32'h3fbeae46} /* (8, 29, 2) {real, imag} */,
  {32'h41024992, 32'h40915804} /* (8, 29, 1) {real, imag} */,
  {32'h40798ccc, 32'hc0242904} /* (8, 29, 0) {real, imag} */,
  {32'h407e25d0, 32'h4128157f} /* (8, 28, 31) {real, imag} */,
  {32'hc11f08f4, 32'hbe81cca8} /* (8, 28, 30) {real, imag} */,
  {32'hc153a248, 32'hc091393c} /* (8, 28, 29) {real, imag} */,
  {32'h3fbdba1a, 32'hc1575a60} /* (8, 28, 28) {real, imag} */,
  {32'hc0e3f0b6, 32'hc0cff712} /* (8, 28, 27) {real, imag} */,
  {32'hc13bf270, 32'hbf526244} /* (8, 28, 26) {real, imag} */,
  {32'h40874fb4, 32'h411cfc70} /* (8, 28, 25) {real, imag} */,
  {32'h40d1cd0a, 32'h41855401} /* (8, 28, 24) {real, imag} */,
  {32'hbf2e1060, 32'h417c698c} /* (8, 28, 23) {real, imag} */,
  {32'hc0fd3390, 32'h41c61ea7} /* (8, 28, 22) {real, imag} */,
  {32'hc1c12244, 32'h3f4fbc98} /* (8, 28, 21) {real, imag} */,
  {32'h3f448bc0, 32'hc0abc039} /* (8, 28, 20) {real, imag} */,
  {32'h4127d419, 32'hc02d1260} /* (8, 28, 19) {real, imag} */,
  {32'hbf994fb0, 32'hc189a476} /* (8, 28, 18) {real, imag} */,
  {32'h40c2f408, 32'hc209947c} /* (8, 28, 17) {real, imag} */,
  {32'h40c69422, 32'hc1fddbc4} /* (8, 28, 16) {real, imag} */,
  {32'hc0a7dfca, 32'hc19d0759} /* (8, 28, 15) {real, imag} */,
  {32'hc10bddf8, 32'hc17b70fa} /* (8, 28, 14) {real, imag} */,
  {32'h3f1ced50, 32'hbf428b40} /* (8, 28, 13) {real, imag} */,
  {32'h40ce56f3, 32'h40910d60} /* (8, 28, 12) {real, imag} */,
  {32'h414961b2, 32'hc0e47d88} /* (8, 28, 11) {real, imag} */,
  {32'h41687fea, 32'h40a22a65} /* (8, 28, 10) {real, imag} */,
  {32'h409f0782, 32'h4113d10e} /* (8, 28, 9) {real, imag} */,
  {32'hc0556234, 32'h4195fd22} /* (8, 28, 8) {real, imag} */,
  {32'hc05917b4, 32'h4145d3d2} /* (8, 28, 7) {real, imag} */,
  {32'h410fe0b7, 32'h414e3616} /* (8, 28, 6) {real, imag} */,
  {32'h414165d0, 32'h41600a88} /* (8, 28, 5) {real, imag} */,
  {32'hc015117d, 32'h40d87786} /* (8, 28, 4) {real, imag} */,
  {32'hc0ab61a7, 32'hc131903a} /* (8, 28, 3) {real, imag} */,
  {32'hbe8055f0, 32'hc083ceab} /* (8, 28, 2) {real, imag} */,
  {32'hbe953c18, 32'h41ac3502} /* (8, 28, 1) {real, imag} */,
  {32'h3ef38bb8, 32'h41944d0b} /* (8, 28, 0) {real, imag} */,
  {32'hbee54740, 32'h40d7975b} /* (8, 27, 31) {real, imag} */,
  {32'hc0ab9529, 32'h3fb49d40} /* (8, 27, 30) {real, imag} */,
  {32'hc06f73ed, 32'hbfbdbd80} /* (8, 27, 29) {real, imag} */,
  {32'hbffe8558, 32'hc0d51806} /* (8, 27, 28) {real, imag} */,
  {32'hc07e9f84, 32'hc1857848} /* (8, 27, 27) {real, imag} */,
  {32'h40148528, 32'hc182d8ca} /* (8, 27, 26) {real, imag} */,
  {32'hc013b4fc, 32'hc0896640} /* (8, 27, 25) {real, imag} */,
  {32'h411bcefd, 32'hbd6eb0c0} /* (8, 27, 24) {real, imag} */,
  {32'hbff64490, 32'hbf0da310} /* (8, 27, 23) {real, imag} */,
  {32'hc04ad884, 32'hc1a560d0} /* (8, 27, 22) {real, imag} */,
  {32'h3f8b9fbc, 32'hc17aaba3} /* (8, 27, 21) {real, imag} */,
  {32'hc0c04870, 32'hc082233d} /* (8, 27, 20) {real, imag} */,
  {32'hc0d6cbf8, 32'h3ff0cc72} /* (8, 27, 19) {real, imag} */,
  {32'h406ad147, 32'hc082e5be} /* (8, 27, 18) {real, imag} */,
  {32'h4020d476, 32'h40635c0a} /* (8, 27, 17) {real, imag} */,
  {32'h40c9f89c, 32'h413c11e6} /* (8, 27, 16) {real, imag} */,
  {32'hbee3c1a0, 32'h41c12eb8} /* (8, 27, 15) {real, imag} */,
  {32'hc00ea55e, 32'hc001fa42} /* (8, 27, 14) {real, imag} */,
  {32'hc0605b66, 32'h40a59cfe} /* (8, 27, 13) {real, imag} */,
  {32'hbf8b6b54, 32'hbfe5ee64} /* (8, 27, 12) {real, imag} */,
  {32'h40077406, 32'h40ec2a42} /* (8, 27, 11) {real, imag} */,
  {32'h40853e74, 32'h40af2d8f} /* (8, 27, 10) {real, imag} */,
  {32'h411e8afc, 32'hc10f7412} /* (8, 27, 9) {real, imag} */,
  {32'h41202765, 32'hc090c961} /* (8, 27, 8) {real, imag} */,
  {32'h3fd238b0, 32'hbfceb2dc} /* (8, 27, 7) {real, imag} */,
  {32'h3ff69518, 32'hc1029c98} /* (8, 27, 6) {real, imag} */,
  {32'hc10acb16, 32'hc0727a7a} /* (8, 27, 5) {real, imag} */,
  {32'hbdd3ba20, 32'hc0dba13e} /* (8, 27, 4) {real, imag} */,
  {32'h408eca5e, 32'hc07721cc} /* (8, 27, 3) {real, imag} */,
  {32'h401111fa, 32'hc0908bb4} /* (8, 27, 2) {real, imag} */,
  {32'h411d354f, 32'hbfe3275c} /* (8, 27, 1) {real, imag} */,
  {32'h407b8f24, 32'hc0152027} /* (8, 27, 0) {real, imag} */,
  {32'h3f9dd1cc, 32'hbe8ea170} /* (8, 26, 31) {real, imag} */,
  {32'hc13ec72d, 32'h40de1cc4} /* (8, 26, 30) {real, imag} */,
  {32'hc1c35792, 32'h401adf42} /* (8, 26, 29) {real, imag} */,
  {32'hc150933b, 32'h405b51ff} /* (8, 26, 28) {real, imag} */,
  {32'hc0e3d7dd, 32'h4159e4a5} /* (8, 26, 27) {real, imag} */,
  {32'hc1051e84, 32'h41644e9d} /* (8, 26, 26) {real, imag} */,
  {32'hbf22dc90, 32'h411e4ae3} /* (8, 26, 25) {real, imag} */,
  {32'hc03e7f20, 32'h404c38b6} /* (8, 26, 24) {real, imag} */,
  {32'hc0c07e6e, 32'hc0d6b4ec} /* (8, 26, 23) {real, imag} */,
  {32'h408516d7, 32'hc07a326e} /* (8, 26, 22) {real, imag} */,
  {32'hbf1f2de4, 32'h419394e3} /* (8, 26, 21) {real, imag} */,
  {32'h402fc4ff, 32'h418c30d0} /* (8, 26, 20) {real, imag} */,
  {32'h409bb3d0, 32'hbffa6fcc} /* (8, 26, 19) {real, imag} */,
  {32'h4108ec8e, 32'hc120bb77} /* (8, 26, 18) {real, imag} */,
  {32'hbf1b22b8, 32'hc1a00d60} /* (8, 26, 17) {real, imag} */,
  {32'hc0f133d4, 32'hc10d99c4} /* (8, 26, 16) {real, imag} */,
  {32'h40342fd3, 32'hc0f0f2d8} /* (8, 26, 15) {real, imag} */,
  {32'hc0ba9847, 32'hc14ea486} /* (8, 26, 14) {real, imag} */,
  {32'h3fd6c744, 32'hbfd20448} /* (8, 26, 13) {real, imag} */,
  {32'hc0ad5b30, 32'hbfc1aede} /* (8, 26, 12) {real, imag} */,
  {32'hc0c2cb5a, 32'h4084de40} /* (8, 26, 11) {real, imag} */,
  {32'hbeb35600, 32'hbf9d6f0d} /* (8, 26, 10) {real, imag} */,
  {32'h3f215c8c, 32'hc060cc7b} /* (8, 26, 9) {real, imag} */,
  {32'h412917da, 32'hbf74cab0} /* (8, 26, 8) {real, imag} */,
  {32'h40c24a2b, 32'h409df158} /* (8, 26, 7) {real, imag} */,
  {32'hc0aa7383, 32'h3eb83ae8} /* (8, 26, 6) {real, imag} */,
  {32'hc1109e02, 32'hc12a0d52} /* (8, 26, 5) {real, imag} */,
  {32'hc1bb6bbc, 32'h404abc9e} /* (8, 26, 4) {real, imag} */,
  {32'hc03c47ed, 32'h40847cf5} /* (8, 26, 3) {real, imag} */,
  {32'h419b0e5f, 32'h3fabb4a8} /* (8, 26, 2) {real, imag} */,
  {32'h40c62d00, 32'hc04b6c6c} /* (8, 26, 1) {real, imag} */,
  {32'h4018f575, 32'hc08465b0} /* (8, 26, 0) {real, imag} */,
  {32'h4018b90d, 32'hc0af3a8e} /* (8, 25, 31) {real, imag} */,
  {32'h4006faba, 32'hc0aeee06} /* (8, 25, 30) {real, imag} */,
  {32'hc0087a9f, 32'h4057a9c8} /* (8, 25, 29) {real, imag} */,
  {32'hbe9c854c, 32'hbf767630} /* (8, 25, 28) {real, imag} */,
  {32'hc166628d, 32'hc0e9ed7e} /* (8, 25, 27) {real, imag} */,
  {32'hc1866316, 32'h41130cb8} /* (8, 25, 26) {real, imag} */,
  {32'hbf1ad418, 32'h418cec39} /* (8, 25, 25) {real, imag} */,
  {32'h409511d3, 32'h409f310a} /* (8, 25, 24) {real, imag} */,
  {32'h403c1d84, 32'h4190e464} /* (8, 25, 23) {real, imag} */,
  {32'hc0a17ea6, 32'h41cfec8c} /* (8, 25, 22) {real, imag} */,
  {32'hc1046d60, 32'h41048b5b} /* (8, 25, 21) {real, imag} */,
  {32'h4059e5a3, 32'h3fc38132} /* (8, 25, 20) {real, imag} */,
  {32'h4123ade2, 32'hc10ec301} /* (8, 25, 19) {real, imag} */,
  {32'h41001618, 32'h3fde46ec} /* (8, 25, 18) {real, imag} */,
  {32'hbf8afce8, 32'h406aadc6} /* (8, 25, 17) {real, imag} */,
  {32'hc08363d4, 32'h40ba7803} /* (8, 25, 16) {real, imag} */,
  {32'hc09e4114, 32'h40b9c0b8} /* (8, 25, 15) {real, imag} */,
  {32'hbf560130, 32'hc064373c} /* (8, 25, 14) {real, imag} */,
  {32'hc043f9e9, 32'h3fb2c568} /* (8, 25, 13) {real, imag} */,
  {32'hc0661ff7, 32'h4132fff2} /* (8, 25, 12) {real, imag} */,
  {32'hc0f575e6, 32'h405c9a9c} /* (8, 25, 11) {real, imag} */,
  {32'hc0a57d7f, 32'h3f994390} /* (8, 25, 10) {real, imag} */,
  {32'hc05ad7bf, 32'hc096197a} /* (8, 25, 9) {real, imag} */,
  {32'hc111680c, 32'hc106318c} /* (8, 25, 8) {real, imag} */,
  {32'hbefbd050, 32'h3fa6c72b} /* (8, 25, 7) {real, imag} */,
  {32'h40f81593, 32'h41730bf0} /* (8, 25, 6) {real, imag} */,
  {32'h413b05cb, 32'h4111c42d} /* (8, 25, 5) {real, imag} */,
  {32'h411b2cff, 32'hbe83354c} /* (8, 25, 4) {real, imag} */,
  {32'h4016a01a, 32'hc06c04b0} /* (8, 25, 3) {real, imag} */,
  {32'hc15b97d9, 32'h40de0350} /* (8, 25, 2) {real, imag} */,
  {32'hc0e35a4f, 32'h4100bba6} /* (8, 25, 1) {real, imag} */,
  {32'h3dc6ce00, 32'h40d5dd8a} /* (8, 25, 0) {real, imag} */,
  {32'h401b19db, 32'h3fc9c868} /* (8, 24, 31) {real, imag} */,
  {32'h40be068e, 32'hc126d25d} /* (8, 24, 30) {real, imag} */,
  {32'h40f21d38, 32'hc18da37c} /* (8, 24, 29) {real, imag} */,
  {32'hbfea34cc, 32'hc138256c} /* (8, 24, 28) {real, imag} */,
  {32'h409deacb, 32'hc006afcc} /* (8, 24, 27) {real, imag} */,
  {32'h40ea19b5, 32'h40940453} /* (8, 24, 26) {real, imag} */,
  {32'h40d1d212, 32'h3f545610} /* (8, 24, 25) {real, imag} */,
  {32'h40f3d806, 32'h4098b59c} /* (8, 24, 24) {real, imag} */,
  {32'h40b0e449, 32'hbe399c28} /* (8, 24, 23) {real, imag} */,
  {32'h40a02b97, 32'hc00df52c} /* (8, 24, 22) {real, imag} */,
  {32'h40bd4c39, 32'hc16aa9ef} /* (8, 24, 21) {real, imag} */,
  {32'hc090ade0, 32'hc0b86431} /* (8, 24, 20) {real, imag} */,
  {32'hc168d09a, 32'h41116610} /* (8, 24, 19) {real, imag} */,
  {32'hc16d91e5, 32'h4115f170} /* (8, 24, 18) {real, imag} */,
  {32'hbf20e78c, 32'h413f54e8} /* (8, 24, 17) {real, imag} */,
  {32'h40cd117e, 32'h41caf366} /* (8, 24, 16) {real, imag} */,
  {32'h401a3b8f, 32'h41cf4048} /* (8, 24, 15) {real, imag} */,
  {32'h403a7d02, 32'h4197c5b2} /* (8, 24, 14) {real, imag} */,
  {32'hbed34aa8, 32'h41199654} /* (8, 24, 13) {real, imag} */,
  {32'h3dbdc700, 32'h413abdbe} /* (8, 24, 12) {real, imag} */,
  {32'h40a139c3, 32'h404b046e} /* (8, 24, 11) {real, imag} */,
  {32'h406f47a2, 32'hc1310620} /* (8, 24, 10) {real, imag} */,
  {32'hbf334908, 32'hc18a4712} /* (8, 24, 9) {real, imag} */,
  {32'h4077c545, 32'hc159be46} /* (8, 24, 8) {real, imag} */,
  {32'h41774293, 32'hc0e04559} /* (8, 24, 7) {real, imag} */,
  {32'h41292ea4, 32'hc099d036} /* (8, 24, 6) {real, imag} */,
  {32'hbf136ad0, 32'hc12c6eed} /* (8, 24, 5) {real, imag} */,
  {32'hc0c599da, 32'hc1658163} /* (8, 24, 4) {real, imag} */,
  {32'hbfe50b2c, 32'hc144f873} /* (8, 24, 3) {real, imag} */,
  {32'h4113592d, 32'hc08f9f32} /* (8, 24, 2) {real, imag} */,
  {32'hc03ce17c, 32'hc02f71a1} /* (8, 24, 1) {real, imag} */,
  {32'hbfb5018c, 32'hc055f444} /* (8, 24, 0) {real, imag} */,
  {32'h408d3ac8, 32'h40862d66} /* (8, 23, 31) {real, imag} */,
  {32'h40b66f2f, 32'h40d54f3a} /* (8, 23, 30) {real, imag} */,
  {32'h40212b3b, 32'h3f805f60} /* (8, 23, 29) {real, imag} */,
  {32'h40a44c09, 32'hc123ebaf} /* (8, 23, 28) {real, imag} */,
  {32'h40bc79de, 32'hc0a5a106} /* (8, 23, 27) {real, imag} */,
  {32'h40f42414, 32'hc0900a55} /* (8, 23, 26) {real, imag} */,
  {32'hc00e6a96, 32'hc0ce788e} /* (8, 23, 25) {real, imag} */,
  {32'h3e7d92f0, 32'h409fb033} /* (8, 23, 24) {real, imag} */,
  {32'h40a22d72, 32'h41144151} /* (8, 23, 23) {real, imag} */,
  {32'hbfeb43c2, 32'h4110dcc8} /* (8, 23, 22) {real, imag} */,
  {32'h40639755, 32'h406fb3df} /* (8, 23, 21) {real, imag} */,
  {32'hc1608a9d, 32'h4108ce26} /* (8, 23, 20) {real, imag} */,
  {32'hc0ca7ef9, 32'h40ccbba0} /* (8, 23, 19) {real, imag} */,
  {32'hc053b472, 32'h40c5893d} /* (8, 23, 18) {real, imag} */,
  {32'h3f553338, 32'h4127174d} /* (8, 23, 17) {real, imag} */,
  {32'h4080ea3c, 32'h404c6236} /* (8, 23, 16) {real, imag} */,
  {32'h3e2727b0, 32'h40fd66d8} /* (8, 23, 15) {real, imag} */,
  {32'h4116c29f, 32'h3fbe1fdc} /* (8, 23, 14) {real, imag} */,
  {32'h40c27fca, 32'h4103fd37} /* (8, 23, 13) {real, imag} */,
  {32'h3f6364bc, 32'h3c3ebb00} /* (8, 23, 12) {real, imag} */,
  {32'hbf9ac2d4, 32'h40a1c5e4} /* (8, 23, 11) {real, imag} */,
  {32'hbe633d40, 32'h410b3eb9} /* (8, 23, 10) {real, imag} */,
  {32'h40953f66, 32'h4118fd90} /* (8, 23, 9) {real, imag} */,
  {32'h40287823, 32'h40d9034d} /* (8, 23, 8) {real, imag} */,
  {32'hc0ce0d93, 32'hc09278df} /* (8, 23, 7) {real, imag} */,
  {32'hc0a2cc6b, 32'h40d694b0} /* (8, 23, 6) {real, imag} */,
  {32'hc0d4dec4, 32'hc030926c} /* (8, 23, 5) {real, imag} */,
  {32'hc11932a9, 32'hc00734b6} /* (8, 23, 4) {real, imag} */,
  {32'hc09077eb, 32'h40aa11ce} /* (8, 23, 3) {real, imag} */,
  {32'hc0fb75d6, 32'hbeaf1158} /* (8, 23, 2) {real, imag} */,
  {32'hc003a69c, 32'hc0a090bd} /* (8, 23, 1) {real, imag} */,
  {32'hc0665314, 32'h4094977f} /* (8, 23, 0) {real, imag} */,
  {32'hc0721e16, 32'h4089d258} /* (8, 22, 31) {real, imag} */,
  {32'hc01a79d6, 32'h4080479e} /* (8, 22, 30) {real, imag} */,
  {32'hc0098386, 32'h40ac9929} /* (8, 22, 29) {real, imag} */,
  {32'hc09b84e2, 32'hbf5554a4} /* (8, 22, 28) {real, imag} */,
  {32'h3f87b216, 32'h3f908316} /* (8, 22, 27) {real, imag} */,
  {32'hbe8e0ae8, 32'hbfdb133f} /* (8, 22, 26) {real, imag} */,
  {32'hc00317f4, 32'h40b3465a} /* (8, 22, 25) {real, imag} */,
  {32'h3fc5632e, 32'h4030c8c1} /* (8, 22, 24) {real, imag} */,
  {32'h3f450a60, 32'hc0c2cff8} /* (8, 22, 23) {real, imag} */,
  {32'h3fb832d7, 32'hc03fed9a} /* (8, 22, 22) {real, imag} */,
  {32'h40bdf05b, 32'hbeac2610} /* (8, 22, 21) {real, imag} */,
  {32'h3f1483e4, 32'hc0d42594} /* (8, 22, 20) {real, imag} */,
  {32'hc0dea034, 32'hbfe96dcc} /* (8, 22, 19) {real, imag} */,
  {32'hc1282dac, 32'h3fc8e452} /* (8, 22, 18) {real, imag} */,
  {32'h3f51d22c, 32'hbe94acf0} /* (8, 22, 17) {real, imag} */,
  {32'hbf683a16, 32'h3ed01518} /* (8, 22, 16) {real, imag} */,
  {32'h3f0a1ecc, 32'h3ed83b60} /* (8, 22, 15) {real, imag} */,
  {32'h40275472, 32'h3ffe05fe} /* (8, 22, 14) {real, imag} */,
  {32'hc0a90f66, 32'h4040c7be} /* (8, 22, 13) {real, imag} */,
  {32'hc188c949, 32'h40ad501f} /* (8, 22, 12) {real, imag} */,
  {32'hc15c13a8, 32'h40712e40} /* (8, 22, 11) {real, imag} */,
  {32'hc132dac2, 32'h40f45d8d} /* (8, 22, 10) {real, imag} */,
  {32'hc07ea183, 32'h4166d570} /* (8, 22, 9) {real, imag} */,
  {32'h4128a1c0, 32'h4166bb4c} /* (8, 22, 8) {real, imag} */,
  {32'h40dacfc5, 32'h4123c844} /* (8, 22, 7) {real, imag} */,
  {32'hc069e5fd, 32'h40e13be0} /* (8, 22, 6) {real, imag} */,
  {32'hc129b7b2, 32'h40cd953c} /* (8, 22, 5) {real, imag} */,
  {32'hc07a7977, 32'hc0331a9a} /* (8, 22, 4) {real, imag} */,
  {32'h410d7736, 32'hbf8d8bca} /* (8, 22, 3) {real, imag} */,
  {32'h40bdf0e5, 32'hc07b0164} /* (8, 22, 2) {real, imag} */,
  {32'h40ce074c, 32'hbf05ad58} /* (8, 22, 1) {real, imag} */,
  {32'h401feef9, 32'hbf41e84c} /* (8, 22, 0) {real, imag} */,
  {32'hbfc20f86, 32'hbfd317c0} /* (8, 21, 31) {real, imag} */,
  {32'hbff51c3d, 32'hbe0673b0} /* (8, 21, 30) {real, imag} */,
  {32'hbfaac232, 32'hc021b430} /* (8, 21, 29) {real, imag} */,
  {32'h3fa3f494, 32'hc0b7f576} /* (8, 21, 28) {real, imag} */,
  {32'hc028558c, 32'h40076f05} /* (8, 21, 27) {real, imag} */,
  {32'h4081d932, 32'h4062c778} /* (8, 21, 26) {real, imag} */,
  {32'h404d7804, 32'hc0c0a638} /* (8, 21, 25) {real, imag} */,
  {32'hc0d4e73d, 32'hc1117c30} /* (8, 21, 24) {real, imag} */,
  {32'hc0a868d9, 32'hc0cf1de2} /* (8, 21, 23) {real, imag} */,
  {32'hc056a038, 32'hc03f4b45} /* (8, 21, 22) {real, imag} */,
  {32'hc03450fc, 32'h3f9dcbb0} /* (8, 21, 21) {real, imag} */,
  {32'h4051db01, 32'hc006fcbe} /* (8, 21, 20) {real, imag} */,
  {32'h3fd00c18, 32'hbf5ccd10} /* (8, 21, 19) {real, imag} */,
  {32'h40a0065e, 32'h407f5cd1} /* (8, 21, 18) {real, imag} */,
  {32'h4012f094, 32'h410ab40f} /* (8, 21, 17) {real, imag} */,
  {32'hc09cd13f, 32'h40b5723f} /* (8, 21, 16) {real, imag} */,
  {32'hc0263ab0, 32'h406ac182} /* (8, 21, 15) {real, imag} */,
  {32'hbf3db66c, 32'h3f8f5b35} /* (8, 21, 14) {real, imag} */,
  {32'hc0547c7c, 32'hc091dbb8} /* (8, 21, 13) {real, imag} */,
  {32'h404ae5d8, 32'h3f827310} /* (8, 21, 12) {real, imag} */,
  {32'h40c2acc9, 32'h40d19409} /* (8, 21, 11) {real, imag} */,
  {32'h403e5b65, 32'h4031256b} /* (8, 21, 10) {real, imag} */,
  {32'h40081853, 32'h40a373ee} /* (8, 21, 9) {real, imag} */,
  {32'hc02cb5a5, 32'h40ae8f9d} /* (8, 21, 8) {real, imag} */,
  {32'hc10981c8, 32'h3f7962a8} /* (8, 21, 7) {real, imag} */,
  {32'hc0a75ffa, 32'hbfdf509e} /* (8, 21, 6) {real, imag} */,
  {32'hc027eb8f, 32'hc0cb8ce4} /* (8, 21, 5) {real, imag} */,
  {32'h40284441, 32'hc073aaf2} /* (8, 21, 4) {real, imag} */,
  {32'h40c660cc, 32'hbf5be068} /* (8, 21, 3) {real, imag} */,
  {32'h4083e83e, 32'hbea827c8} /* (8, 21, 2) {real, imag} */,
  {32'hbf2fccf0, 32'h3e7e12a0} /* (8, 21, 1) {real, imag} */,
  {32'hbf702c84, 32'h3eeaa8b8} /* (8, 21, 0) {real, imag} */,
  {32'hc0d8d290, 32'h3f2627b4} /* (8, 20, 31) {real, imag} */,
  {32'h3f8247c2, 32'hbc86a280} /* (8, 20, 30) {real, imag} */,
  {32'h40d6ca6b, 32'hbfb401ca} /* (8, 20, 29) {real, imag} */,
  {32'h40b767ad, 32'h3fa7072c} /* (8, 20, 28) {real, imag} */,
  {32'h408b4062, 32'hbdf1aa40} /* (8, 20, 27) {real, imag} */,
  {32'hbead76b0, 32'h3f0b3a34} /* (8, 20, 26) {real, imag} */,
  {32'h40160abf, 32'hc05bda40} /* (8, 20, 25) {real, imag} */,
  {32'hbff9b640, 32'hc053687f} /* (8, 20, 24) {real, imag} */,
  {32'hc0738116, 32'hc0176912} /* (8, 20, 23) {real, imag} */,
  {32'hc08f69b6, 32'h4086b3ce} /* (8, 20, 22) {real, imag} */,
  {32'hbc965c00, 32'h3fe4d5c0} /* (8, 20, 21) {real, imag} */,
  {32'h3f833724, 32'h3f6429c8} /* (8, 20, 20) {real, imag} */,
  {32'h3b1c2600, 32'h403891ba} /* (8, 20, 19) {real, imag} */,
  {32'hc0b76522, 32'hc0361081} /* (8, 20, 18) {real, imag} */,
  {32'hc0aa38a1, 32'hc0bd02bf} /* (8, 20, 17) {real, imag} */,
  {32'h3f454380, 32'hc0b00f3e} /* (8, 20, 16) {real, imag} */,
  {32'h3f7668b4, 32'hc0169bf4} /* (8, 20, 15) {real, imag} */,
  {32'hbd83f980, 32'hbfec12a0} /* (8, 20, 14) {real, imag} */,
  {32'hc00119a4, 32'h3f7342ec} /* (8, 20, 13) {real, imag} */,
  {32'hc0867673, 32'hbf7b81f2} /* (8, 20, 12) {real, imag} */,
  {32'hc034833e, 32'h4049d1b2} /* (8, 20, 11) {real, imag} */,
  {32'h40706bf2, 32'h407f35c2} /* (8, 20, 10) {real, imag} */,
  {32'h400e9de1, 32'h4056ffe3} /* (8, 20, 9) {real, imag} */,
  {32'hc087cfb9, 32'hc0c74a8e} /* (8, 20, 8) {real, imag} */,
  {32'hc0157e5e, 32'hc12d0998} /* (8, 20, 7) {real, imag} */,
  {32'hc09b6f81, 32'hbf593eb8} /* (8, 20, 6) {real, imag} */,
  {32'hbd981a00, 32'hc03db5e3} /* (8, 20, 5) {real, imag} */,
  {32'h4003d069, 32'hc0a2ea6c} /* (8, 20, 4) {real, imag} */,
  {32'h3ea999f4, 32'hc0a5b944} /* (8, 20, 3) {real, imag} */,
  {32'hc04d48c6, 32'hbfd68619} /* (8, 20, 2) {real, imag} */,
  {32'h3fa10388, 32'hc0afbf28} /* (8, 20, 1) {real, imag} */,
  {32'hbfb702aa, 32'hc086806e} /* (8, 20, 0) {real, imag} */,
  {32'hbea69c74, 32'h3f26c6e6} /* (8, 19, 31) {real, imag} */,
  {32'hc00277bf, 32'hc07265cc} /* (8, 19, 30) {real, imag} */,
  {32'hc038223d, 32'hbf956854} /* (8, 19, 29) {real, imag} */,
  {32'hc056be07, 32'h402deffe} /* (8, 19, 28) {real, imag} */,
  {32'hc04c0186, 32'h3efe3038} /* (8, 19, 27) {real, imag} */,
  {32'hc0cbc1f8, 32'h4015cfd3} /* (8, 19, 26) {real, imag} */,
  {32'hc0a748be, 32'hc0263752} /* (8, 19, 25) {real, imag} */,
  {32'h3ef26354, 32'hbfc22fb2} /* (8, 19, 24) {real, imag} */,
  {32'hc033ca15, 32'h40a04d96} /* (8, 19, 23) {real, imag} */,
  {32'hbef96fe8, 32'h4006504c} /* (8, 19, 22) {real, imag} */,
  {32'hbf7b0cc0, 32'hc049bc25} /* (8, 19, 21) {real, imag} */,
  {32'h3f68f2b0, 32'hc097db12} /* (8, 19, 20) {real, imag} */,
  {32'h400aba30, 32'hbf98f498} /* (8, 19, 19) {real, imag} */,
  {32'h400bcc6d, 32'h3f911e28} /* (8, 19, 18) {real, imag} */,
  {32'h40e818a8, 32'hbfef297f} /* (8, 19, 17) {real, imag} */,
  {32'h3f99f29c, 32'hbfbe1222} /* (8, 19, 16) {real, imag} */,
  {32'h3fe1d9ed, 32'h3e303180} /* (8, 19, 15) {real, imag} */,
  {32'h40ac1561, 32'h3fac7615} /* (8, 19, 14) {real, imag} */,
  {32'h406e5030, 32'h3ff38752} /* (8, 19, 13) {real, imag} */,
  {32'h40aff528, 32'hc0bb007f} /* (8, 19, 12) {real, imag} */,
  {32'hbe89aa70, 32'hc09289a6} /* (8, 19, 11) {real, imag} */,
  {32'h3e6a56b0, 32'hc00787e4} /* (8, 19, 10) {real, imag} */,
  {32'h405434b5, 32'hbf6d5c82} /* (8, 19, 9) {real, imag} */,
  {32'h408800d7, 32'h40c345af} /* (8, 19, 8) {real, imag} */,
  {32'h408e7996, 32'h40753176} /* (8, 19, 7) {real, imag} */,
  {32'h40746e7e, 32'h400cceb4} /* (8, 19, 6) {real, imag} */,
  {32'h4015e7bc, 32'hbec80d00} /* (8, 19, 5) {real, imag} */,
  {32'hbf9732d4, 32'hc08ae4a2} /* (8, 19, 4) {real, imag} */,
  {32'h3d331620, 32'h3f040be8} /* (8, 19, 3) {real, imag} */,
  {32'h400346b6, 32'h4039d915} /* (8, 19, 2) {real, imag} */,
  {32'h409f0f8c, 32'hc08d7cda} /* (8, 19, 1) {real, imag} */,
  {32'h40a5d7d0, 32'hbf3a5a78} /* (8, 19, 0) {real, imag} */,
  {32'hc06a0759, 32'h3ff3b510} /* (8, 18, 31) {real, imag} */,
  {32'hc0f329e4, 32'hbf82c0f8} /* (8, 18, 30) {real, imag} */,
  {32'hc048f116, 32'hc00ac658} /* (8, 18, 29) {real, imag} */,
  {32'hc00fccba, 32'hc0049248} /* (8, 18, 28) {real, imag} */,
  {32'hc0c58be4, 32'hc0101ff7} /* (8, 18, 27) {real, imag} */,
  {32'hc0c95bd1, 32'hbfe1a22f} /* (8, 18, 26) {real, imag} */,
  {32'hc001eb53, 32'hbf965f2e} /* (8, 18, 25) {real, imag} */,
  {32'h40b6ff4c, 32'hc0006b62} /* (8, 18, 24) {real, imag} */,
  {32'hbf3118f0, 32'h3fdf4878} /* (8, 18, 23) {real, imag} */,
  {32'hc0bcc7a8, 32'h3fc506a0} /* (8, 18, 22) {real, imag} */,
  {32'hc01d5f88, 32'hc02299d2} /* (8, 18, 21) {real, imag} */,
  {32'hc08814ec, 32'hbee93dd8} /* (8, 18, 20) {real, imag} */,
  {32'hc041646c, 32'h405f74db} /* (8, 18, 19) {real, imag} */,
  {32'h3f945b0c, 32'h3e70a3f8} /* (8, 18, 18) {real, imag} */,
  {32'h3ea4cf50, 32'h3f8b80b8} /* (8, 18, 17) {real, imag} */,
  {32'h3fa39eae, 32'h3f617ee0} /* (8, 18, 16) {real, imag} */,
  {32'h3fc9fdfa, 32'hbe3331a0} /* (8, 18, 15) {real, imag} */,
  {32'h4099e55c, 32'hbf1a6f1a} /* (8, 18, 14) {real, imag} */,
  {32'h3fad1766, 32'h3fc363f8} /* (8, 18, 13) {real, imag} */,
  {32'hc013f333, 32'hbfbdfada} /* (8, 18, 12) {real, imag} */,
  {32'hc035e066, 32'hbe3c1ba0} /* (8, 18, 11) {real, imag} */,
  {32'hbf0b63d8, 32'h4089b574} /* (8, 18, 10) {real, imag} */,
  {32'hc0297b4e, 32'h4066decb} /* (8, 18, 9) {real, imag} */,
  {32'h3fe6dda4, 32'h3fa8f789} /* (8, 18, 8) {real, imag} */,
  {32'h3f6dbbf8, 32'hc08a0fe0} /* (8, 18, 7) {real, imag} */,
  {32'hc08c087d, 32'hc0d4b00e} /* (8, 18, 6) {real, imag} */,
  {32'hbfd29090, 32'hbfcc4804} /* (8, 18, 5) {real, imag} */,
  {32'h405392a4, 32'h3f88997c} /* (8, 18, 4) {real, imag} */,
  {32'h4076ea78, 32'hc06fa86c} /* (8, 18, 3) {real, imag} */,
  {32'h3f3ae234, 32'hbea74060} /* (8, 18, 2) {real, imag} */,
  {32'hbff01bd4, 32'h402a9435} /* (8, 18, 1) {real, imag} */,
  {32'h3e910c44, 32'h3ec517f0} /* (8, 18, 0) {real, imag} */,
  {32'hc06cb6a6, 32'hbecda098} /* (8, 17, 31) {real, imag} */,
  {32'hbf841598, 32'hc06c7d2a} /* (8, 17, 30) {real, imag} */,
  {32'h40140304, 32'h3e66f4c0} /* (8, 17, 29) {real, imag} */,
  {32'h40263c90, 32'h3f8c9e44} /* (8, 17, 28) {real, imag} */,
  {32'h3fa25ba0, 32'hbf1c6666} /* (8, 17, 27) {real, imag} */,
  {32'h4034673d, 32'h3e2ef2f0} /* (8, 17, 26) {real, imag} */,
  {32'h4010cc31, 32'hbe80afc0} /* (8, 17, 25) {real, imag} */,
  {32'hbffa81c2, 32'hc09f3d66} /* (8, 17, 24) {real, imag} */,
  {32'hbf9bfe50, 32'hc0147ada} /* (8, 17, 23) {real, imag} */,
  {32'h4036595e, 32'hbf52b0ca} /* (8, 17, 22) {real, imag} */,
  {32'h3e946ad0, 32'hbfe28bbc} /* (8, 17, 21) {real, imag} */,
  {32'hbfb5525a, 32'hbe22d840} /* (8, 17, 20) {real, imag} */,
  {32'hbf938c8c, 32'hbf87afe6} /* (8, 17, 19) {real, imag} */,
  {32'hbff55e30, 32'hbf8e9180} /* (8, 17, 18) {real, imag} */,
  {32'hbfeb5040, 32'h3f84d698} /* (8, 17, 17) {real, imag} */,
  {32'hc0108970, 32'h4072bcea} /* (8, 17, 16) {real, imag} */,
  {32'hbfa892a1, 32'h3feeda32} /* (8, 17, 15) {real, imag} */,
  {32'h3f9efa79, 32'h3f25752a} /* (8, 17, 14) {real, imag} */,
  {32'h4049320b, 32'hc02d7e38} /* (8, 17, 13) {real, imag} */,
  {32'hbe5781c0, 32'hbe5a1c48} /* (8, 17, 12) {real, imag} */,
  {32'hc0c3086e, 32'h405b4fff} /* (8, 17, 11) {real, imag} */,
  {32'hc09805cc, 32'h3fb4784c} /* (8, 17, 10) {real, imag} */,
  {32'h3ed8a1b0, 32'h3fd4eba0} /* (8, 17, 9) {real, imag} */,
  {32'h3f6238d5, 32'h4019d444} /* (8, 17, 8) {real, imag} */,
  {32'h40102f9e, 32'h40dc95dd} /* (8, 17, 7) {real, imag} */,
  {32'h3f66a9b0, 32'h40ee17ee} /* (8, 17, 6) {real, imag} */,
  {32'h40284f83, 32'hbe7411e0} /* (8, 17, 5) {real, imag} */,
  {32'hbf141fd8, 32'hc01322e5} /* (8, 17, 4) {real, imag} */,
  {32'hc057487e, 32'hbfd13845} /* (8, 17, 3) {real, imag} */,
  {32'h3cf888e0, 32'hc0726933} /* (8, 17, 2) {real, imag} */,
  {32'h40572c40, 32'h400ce1fe} /* (8, 17, 1) {real, imag} */,
  {32'hbd459980, 32'h40610cc4} /* (8, 17, 0) {real, imag} */,
  {32'h3f5938e8, 32'hc08e562e} /* (8, 16, 31) {real, imag} */,
  {32'h3ed579a0, 32'hc0f03920} /* (8, 16, 30) {real, imag} */,
  {32'hc019c710, 32'hc1065af1} /* (8, 16, 29) {real, imag} */,
  {32'hbfb44c58, 32'hc0c520d8} /* (8, 16, 28) {real, imag} */,
  {32'hbfcca1c0, 32'hc080ebac} /* (8, 16, 27) {real, imag} */,
  {32'hbfc8a184, 32'hbeaefc10} /* (8, 16, 26) {real, imag} */,
  {32'hc016805f, 32'h3ea7b9a0} /* (8, 16, 25) {real, imag} */,
  {32'h4059895a, 32'hc01a3b73} /* (8, 16, 24) {real, imag} */,
  {32'h3f760130, 32'hbfd8efcf} /* (8, 16, 23) {real, imag} */,
  {32'hbe3bd200, 32'h3e51b240} /* (8, 16, 22) {real, imag} */,
  {32'h3e6461e0, 32'h3f996cc0} /* (8, 16, 21) {real, imag} */,
  {32'h3ffb85c6, 32'hbfd10b50} /* (8, 16, 20) {real, imag} */,
  {32'h405f7294, 32'hc0881a7e} /* (8, 16, 19) {real, imag} */,
  {32'h400a02e7, 32'hc08d7a20} /* (8, 16, 18) {real, imag} */,
  {32'hbfae1082, 32'hc06c4b04} /* (8, 16, 17) {real, imag} */,
  {32'h3e886408, 32'hc04bb336} /* (8, 16, 16) {real, imag} */,
  {32'h407fe954, 32'hbf1548d0} /* (8, 16, 15) {real, imag} */,
  {32'h3ee31d80, 32'hbde379c0} /* (8, 16, 14) {real, imag} */,
  {32'hbbcda800, 32'hc01be2c8} /* (8, 16, 13) {real, imag} */,
  {32'h3f84bc90, 32'hc01c80f6} /* (8, 16, 12) {real, imag} */,
  {32'h3f37cc30, 32'hc05c190c} /* (8, 16, 11) {real, imag} */,
  {32'h3fad6298, 32'h4056ee1e} /* (8, 16, 10) {real, imag} */,
  {32'hbff80562, 32'h409a304d} /* (8, 16, 9) {real, imag} */,
  {32'h3e7c8e60, 32'h3db03e80} /* (8, 16, 8) {real, imag} */,
  {32'hbfd86a38, 32'hc0b66e78} /* (8, 16, 7) {real, imag} */,
  {32'hbfe43510, 32'hc0887ae4} /* (8, 16, 6) {real, imag} */,
  {32'h3f9abad2, 32'hbe491600} /* (8, 16, 5) {real, imag} */,
  {32'h3ecafa90, 32'hbd774400} /* (8, 16, 4) {real, imag} */,
  {32'hc09695a4, 32'h3fb37978} /* (8, 16, 3) {real, imag} */,
  {32'hc0b0860e, 32'h3fc9c050} /* (8, 16, 2) {real, imag} */,
  {32'hc0752c8c, 32'h4021f970} /* (8, 16, 1) {real, imag} */,
  {32'hbfc61290, 32'h3fb3fec8} /* (8, 16, 0) {real, imag} */,
  {32'h402cad82, 32'h3f965bfe} /* (8, 15, 31) {real, imag} */,
  {32'h4020bab4, 32'h3ffd13c4} /* (8, 15, 30) {real, imag} */,
  {32'hbeccc060, 32'hbfe4a458} /* (8, 15, 29) {real, imag} */,
  {32'h3ecc1180, 32'hbfcb76d4} /* (8, 15, 28) {real, imag} */,
  {32'h3f85f1e0, 32'hbfc1f46d} /* (8, 15, 27) {real, imag} */,
  {32'hbe8adb68, 32'hc0113247} /* (8, 15, 26) {real, imag} */,
  {32'h3fb9053e, 32'hc09314ac} /* (8, 15, 25) {real, imag} */,
  {32'h3fe80562, 32'hc02ff35c} /* (8, 15, 24) {real, imag} */,
  {32'h40494ce8, 32'hbf8fa6cc} /* (8, 15, 23) {real, imag} */,
  {32'h4070a0f2, 32'hc05d1e6e} /* (8, 15, 22) {real, imag} */,
  {32'h40223396, 32'hc01a5712} /* (8, 15, 21) {real, imag} */,
  {32'h3db2e460, 32'hbf16d890} /* (8, 15, 20) {real, imag} */,
  {32'hbfa9a0ec, 32'hc01e995f} /* (8, 15, 19) {real, imag} */,
  {32'hbf3eb240, 32'h3ddf9c00} /* (8, 15, 18) {real, imag} */,
  {32'h40344178, 32'h406627b4} /* (8, 15, 17) {real, imag} */,
  {32'h3fc811d0, 32'h409b3507} /* (8, 15, 16) {real, imag} */,
  {32'h3f36a582, 32'h40a0dae4} /* (8, 15, 15) {real, imag} */,
  {32'h3f080aee, 32'hbf284f2a} /* (8, 15, 14) {real, imag} */,
  {32'hc00c5e4b, 32'hc00e36c0} /* (8, 15, 13) {real, imag} */,
  {32'h3f75d4b0, 32'hc019c1ac} /* (8, 15, 12) {real, imag} */,
  {32'h3f94c0f8, 32'hc020555f} /* (8, 15, 11) {real, imag} */,
  {32'hbfa37512, 32'hc01b991a} /* (8, 15, 10) {real, imag} */,
  {32'hc008375a, 32'hc092243e} /* (8, 15, 9) {real, imag} */,
  {32'hc036264b, 32'hc036f62c} /* (8, 15, 8) {real, imag} */,
  {32'hc02eedfc, 32'h3f0bf038} /* (8, 15, 7) {real, imag} */,
  {32'hbfd50c40, 32'hbeed7358} /* (8, 15, 6) {real, imag} */,
  {32'hbf525f8c, 32'hbff76fe4} /* (8, 15, 5) {real, imag} */,
  {32'h3ee681f0, 32'hc084b56e} /* (8, 15, 4) {real, imag} */,
  {32'h4019017e, 32'hc0969fff} /* (8, 15, 3) {real, imag} */,
  {32'h3f5999d9, 32'hbecc92e8} /* (8, 15, 2) {real, imag} */,
  {32'hbf194362, 32'hbe5ef0e8} /* (8, 15, 1) {real, imag} */,
  {32'hc001d0e2, 32'hbfa2d908} /* (8, 15, 0) {real, imag} */,
  {32'hbeb574a8, 32'hbcbfb600} /* (8, 14, 31) {real, imag} */,
  {32'h3fdc6552, 32'h3f6cdb30} /* (8, 14, 30) {real, imag} */,
  {32'h40d70adf, 32'h3fb8122f} /* (8, 14, 29) {real, imag} */,
  {32'h40280be2, 32'h3ea740c0} /* (8, 14, 28) {real, imag} */,
  {32'hbffd1e80, 32'h4068c4cf} /* (8, 14, 27) {real, imag} */,
  {32'hc06ef72a, 32'h3f88e6ff} /* (8, 14, 26) {real, imag} */,
  {32'h3fcdedba, 32'hc046e9a9} /* (8, 14, 25) {real, imag} */,
  {32'h400e7ec7, 32'hbe3d4258} /* (8, 14, 24) {real, imag} */,
  {32'h4010eabc, 32'h3f2c0fa0} /* (8, 14, 23) {real, imag} */,
  {32'h4052ed40, 32'hc0950b54} /* (8, 14, 22) {real, imag} */,
  {32'hbfc2d898, 32'hc0881b11} /* (8, 14, 21) {real, imag} */,
  {32'h3e84fb48, 32'hbf80b342} /* (8, 14, 20) {real, imag} */,
  {32'h3ef12ba0, 32'h3fc79baa} /* (8, 14, 19) {real, imag} */,
  {32'h407a636e, 32'h3ff0ef11} /* (8, 14, 18) {real, imag} */,
  {32'hbff01434, 32'h4035066c} /* (8, 14, 17) {real, imag} */,
  {32'hc083d7cc, 32'hc02964d8} /* (8, 14, 16) {real, imag} */,
  {32'hbfd5366a, 32'hc0752f4e} /* (8, 14, 15) {real, imag} */,
  {32'h3f0a66e4, 32'hbf8be485} /* (8, 14, 14) {real, imag} */,
  {32'hbbd65600, 32'h3f0b5930} /* (8, 14, 13) {real, imag} */,
  {32'hbfb3e09a, 32'hbf3291dc} /* (8, 14, 12) {real, imag} */,
  {32'hbfcdff34, 32'h403d8026} /* (8, 14, 11) {real, imag} */,
  {32'hc0964b65, 32'hbe66c490} /* (8, 14, 10) {real, imag} */,
  {32'h40082046, 32'hbf8333d6} /* (8, 14, 9) {real, imag} */,
  {32'h40112846, 32'hbfc0f8e9} /* (8, 14, 8) {real, imag} */,
  {32'h40a052fd, 32'hbe678c80} /* (8, 14, 7) {real, imag} */,
  {32'h40d32cbd, 32'h40612e4c} /* (8, 14, 6) {real, imag} */,
  {32'h40b55024, 32'h4039edfe} /* (8, 14, 5) {real, imag} */,
  {32'hbfc4e2c8, 32'h40287272} /* (8, 14, 4) {real, imag} */,
  {32'hc0a7216c, 32'h40e2840e} /* (8, 14, 3) {real, imag} */,
  {32'hbf9f569a, 32'h4040bf74} /* (8, 14, 2) {real, imag} */,
  {32'h403792aa, 32'h3f5c5eec} /* (8, 14, 1) {real, imag} */,
  {32'h3f955f57, 32'h3e12f120} /* (8, 14, 0) {real, imag} */,
  {32'hc04e89c2, 32'hbefdcb74} /* (8, 13, 31) {real, imag} */,
  {32'hc028b22f, 32'hbf119360} /* (8, 13, 30) {real, imag} */,
  {32'hc02dc2ab, 32'h3ff33500} /* (8, 13, 29) {real, imag} */,
  {32'hbfc51aea, 32'h3f9b939c} /* (8, 13, 28) {real, imag} */,
  {32'hc006d35e, 32'hc0151869} /* (8, 13, 27) {real, imag} */,
  {32'h3fb4047e, 32'hbfcffc8c} /* (8, 13, 26) {real, imag} */,
  {32'h40a67780, 32'h3fe1821c} /* (8, 13, 25) {real, imag} */,
  {32'h40000b3a, 32'hc0a1cd94} /* (8, 13, 24) {real, imag} */,
  {32'hbf851bc6, 32'hc087769e} /* (8, 13, 23) {real, imag} */,
  {32'hc05047fd, 32'h408100cb} /* (8, 13, 22) {real, imag} */,
  {32'hbfa5bc20, 32'h3e72e730} /* (8, 13, 21) {real, imag} */,
  {32'hbfaf1338, 32'hbd438c00} /* (8, 13, 20) {real, imag} */,
  {32'h407d8c50, 32'hc029180d} /* (8, 13, 19) {real, imag} */,
  {32'h402d6535, 32'hc063ba0c} /* (8, 13, 18) {real, imag} */,
  {32'hbec3aa88, 32'hc09c101c} /* (8, 13, 17) {real, imag} */,
  {32'h40321862, 32'hc10d2ca8} /* (8, 13, 16) {real, imag} */,
  {32'h3f862f27, 32'hc109341c} /* (8, 13, 15) {real, imag} */,
  {32'hc02857d2, 32'hc091dea5} /* (8, 13, 14) {real, imag} */,
  {32'h3f9785cf, 32'hc0745179} /* (8, 13, 13) {real, imag} */,
  {32'h3f345ea4, 32'hc0498062} /* (8, 13, 12) {real, imag} */,
  {32'h40a8ba69, 32'h3f951cca} /* (8, 13, 11) {real, imag} */,
  {32'h405081f3, 32'h3f773540} /* (8, 13, 10) {real, imag} */,
  {32'h3f660e2c, 32'hc03fd0bc} /* (8, 13, 9) {real, imag} */,
  {32'hbf919a44, 32'h40503286} /* (8, 13, 8) {real, imag} */,
  {32'hbfc201ea, 32'h3fb64a6c} /* (8, 13, 7) {real, imag} */,
  {32'hc0112aee, 32'h3fa31f38} /* (8, 13, 6) {real, imag} */,
  {32'h3fd7cf48, 32'h40b6ec0c} /* (8, 13, 5) {real, imag} */,
  {32'hc01aecee, 32'h3fcba786} /* (8, 13, 4) {real, imag} */,
  {32'hc0331cac, 32'hc11296da} /* (8, 13, 3) {real, imag} */,
  {32'hbf6320f2, 32'hc059721f} /* (8, 13, 2) {real, imag} */,
  {32'h3fc3ef37, 32'h40732477} /* (8, 13, 1) {real, imag} */,
  {32'h3f85cfee, 32'h3f803a46} /* (8, 13, 0) {real, imag} */,
  {32'h403e3ac4, 32'hbfc73a16} /* (8, 12, 31) {real, imag} */,
  {32'hc049e7a7, 32'hc081ebf0} /* (8, 12, 30) {real, imag} */,
  {32'hc0a8cd47, 32'h401b1cdd} /* (8, 12, 29) {real, imag} */,
  {32'h4060a6ae, 32'h41071402} /* (8, 12, 28) {real, imag} */,
  {32'h3fbcd090, 32'h408ce835} /* (8, 12, 27) {real, imag} */,
  {32'hbf4f2958, 32'hc02aaf3f} /* (8, 12, 26) {real, imag} */,
  {32'hc0a40770, 32'hbfef1091} /* (8, 12, 25) {real, imag} */,
  {32'h3f24e021, 32'h40bed398} /* (8, 12, 24) {real, imag} */,
  {32'h3ff39034, 32'h409f5e9f} /* (8, 12, 23) {real, imag} */,
  {32'h4057b61d, 32'h408d4d66} /* (8, 12, 22) {real, imag} */,
  {32'hc0cace44, 32'hbd35cc40} /* (8, 12, 21) {real, imag} */,
  {32'hc062a5f2, 32'hc0339827} /* (8, 12, 20) {real, imag} */,
  {32'hc02fa61e, 32'hbf83e9e7} /* (8, 12, 19) {real, imag} */,
  {32'hc02a57c8, 32'hc0712631} /* (8, 12, 18) {real, imag} */,
  {32'hc02a77f6, 32'hc0cd542b} /* (8, 12, 17) {real, imag} */,
  {32'hbfb45410, 32'h3f47eb74} /* (8, 12, 16) {real, imag} */,
  {32'h40927f8c, 32'h3fd32218} /* (8, 12, 15) {real, imag} */,
  {32'h40a025ec, 32'h3d712e00} /* (8, 12, 14) {real, imag} */,
  {32'h411502fb, 32'hc06d4145} /* (8, 12, 13) {real, imag} */,
  {32'h40b8c94b, 32'h409c24da} /* (8, 12, 12) {real, imag} */,
  {32'h3f8fff00, 32'h3f7253d6} /* (8, 12, 11) {real, imag} */,
  {32'hc0de9623, 32'hbb52f800} /* (8, 12, 10) {real, imag} */,
  {32'hc0aadf76, 32'h4002fd53} /* (8, 12, 9) {real, imag} */,
  {32'h409e9fa3, 32'h3f950806} /* (8, 12, 8) {real, imag} */,
  {32'h40810271, 32'hc010312e} /* (8, 12, 7) {real, imag} */,
  {32'h3efa2650, 32'h3ef89bd0} /* (8, 12, 6) {real, imag} */,
  {32'h40398f78, 32'h40339e99} /* (8, 12, 5) {real, imag} */,
  {32'h3f9d5376, 32'h4093786e} /* (8, 12, 4) {real, imag} */,
  {32'h3dfa5bf0, 32'h3fe698ed} /* (8, 12, 3) {real, imag} */,
  {32'hc041d740, 32'h3fe4e197} /* (8, 12, 2) {real, imag} */,
  {32'hc0e19584, 32'h3ffb1201} /* (8, 12, 1) {real, imag} */,
  {32'hc006b0cd, 32'hc05ad1d4} /* (8, 12, 0) {real, imag} */,
  {32'h40945616, 32'h3fe71526} /* (8, 11, 31) {real, imag} */,
  {32'h408c21aa, 32'h3fbc2724} /* (8, 11, 30) {real, imag} */,
  {32'hc0040d5d, 32'h4109cdec} /* (8, 11, 29) {real, imag} */,
  {32'hc04c9290, 32'h4111d161} /* (8, 11, 28) {real, imag} */,
  {32'hc0c4c1fe, 32'h40e9be5a} /* (8, 11, 27) {real, imag} */,
  {32'h3ea8efc0, 32'h413e009e} /* (8, 11, 26) {real, imag} */,
  {32'h40bd7ff2, 32'h3fb83386} /* (8, 11, 25) {real, imag} */,
  {32'h400781ae, 32'h4063ff2b} /* (8, 11, 24) {real, imag} */,
  {32'h404d3aa2, 32'h4083a80e} /* (8, 11, 23) {real, imag} */,
  {32'h40f5ed10, 32'h4089d836} /* (8, 11, 22) {real, imag} */,
  {32'h40cda4d8, 32'h3f5c1e38} /* (8, 11, 21) {real, imag} */,
  {32'hc0be6684, 32'hc00b9e2a} /* (8, 11, 20) {real, imag} */,
  {32'hc119671b, 32'h403eed92} /* (8, 11, 19) {real, imag} */,
  {32'hc0647b24, 32'hbfb42e42} /* (8, 11, 18) {real, imag} */,
  {32'h40860bca, 32'hc08797e2} /* (8, 11, 17) {real, imag} */,
  {32'h400c128a, 32'hbf5bb9e0} /* (8, 11, 16) {real, imag} */,
  {32'hc0aabedc, 32'h3ebfcb90} /* (8, 11, 15) {real, imag} */,
  {32'hc09b3922, 32'hc0757630} /* (8, 11, 14) {real, imag} */,
  {32'hc0ccfea4, 32'h3e092490} /* (8, 11, 13) {real, imag} */,
  {32'h3f3435e4, 32'h40db7ec6} /* (8, 11, 12) {real, imag} */,
  {32'h3fa92adc, 32'h4052cbce} /* (8, 11, 11) {real, imag} */,
  {32'hbe910b78, 32'hbe61a790} /* (8, 11, 10) {real, imag} */,
  {32'hc0051157, 32'h402e54e9} /* (8, 11, 9) {real, imag} */,
  {32'hbee9e4d8, 32'hc01a0b9a} /* (8, 11, 8) {real, imag} */,
  {32'h3f74a4a0, 32'hc098d07c} /* (8, 11, 7) {real, imag} */,
  {32'h40bf5812, 32'h3fc4aef6} /* (8, 11, 6) {real, imag} */,
  {32'h40f72770, 32'h402b32c4} /* (8, 11, 5) {real, imag} */,
  {32'h40a8c416, 32'h403628fe} /* (8, 11, 4) {real, imag} */,
  {32'h40b90226, 32'h40ca88b3} /* (8, 11, 3) {real, imag} */,
  {32'h40b2bdb6, 32'h40237185} /* (8, 11, 2) {real, imag} */,
  {32'h40d37128, 32'hc0b3a8fd} /* (8, 11, 1) {real, imag} */,
  {32'h4001b279, 32'hbfa4b0c2} /* (8, 11, 0) {real, imag} */,
  {32'hc0b8a6e3, 32'hbf279f6c} /* (8, 10, 31) {real, imag} */,
  {32'hc06e1d96, 32'h400d9c7f} /* (8, 10, 30) {real, imag} */,
  {32'h3ef68a8c, 32'h3f9e7b20} /* (8, 10, 29) {real, imag} */,
  {32'hbf40097c, 32'hc0f0ef5a} /* (8, 10, 28) {real, imag} */,
  {32'hbf95ec52, 32'hc017290f} /* (8, 10, 27) {real, imag} */,
  {32'h3e093790, 32'hc07fb048} /* (8, 10, 26) {real, imag} */,
  {32'hbf0a0880, 32'hc0a144d6} /* (8, 10, 25) {real, imag} */,
  {32'h3f8b4606, 32'hc03bfff5} /* (8, 10, 24) {real, imag} */,
  {32'h4033bb38, 32'hc0380cf4} /* (8, 10, 23) {real, imag} */,
  {32'hbf952a39, 32'hbf533df0} /* (8, 10, 22) {real, imag} */,
  {32'hc0644bee, 32'hc035aaea} /* (8, 10, 21) {real, imag} */,
  {32'h409e94da, 32'h40abb93c} /* (8, 10, 20) {real, imag} */,
  {32'h40f9004c, 32'h40b7cc71} /* (8, 10, 19) {real, imag} */,
  {32'h40ccf593, 32'h406a5ec5} /* (8, 10, 18) {real, imag} */,
  {32'h4102e0c5, 32'h40473a8a} /* (8, 10, 17) {real, imag} */,
  {32'h3f421e26, 32'h4057a1b9} /* (8, 10, 16) {real, imag} */,
  {32'h4008d877, 32'h40926295} /* (8, 10, 15) {real, imag} */,
  {32'hbf48c618, 32'hbf86aba2} /* (8, 10, 14) {real, imag} */,
  {32'h3ef395b8, 32'hc0ad0e97} /* (8, 10, 13) {real, imag} */,
  {32'hbfa81c50, 32'hc004a8f8} /* (8, 10, 12) {real, imag} */,
  {32'hc0ac96d0, 32'h3e1e9900} /* (8, 10, 11) {real, imag} */,
  {32'hc0d3760c, 32'hbe31a820} /* (8, 10, 10) {real, imag} */,
  {32'hc1155fa3, 32'hbd873dc0} /* (8, 10, 9) {real, imag} */,
  {32'hc141170e, 32'h40c055c4} /* (8, 10, 8) {real, imag} */,
  {32'hc0c16f87, 32'h40a9d41c} /* (8, 10, 7) {real, imag} */,
  {32'hbfd4bf02, 32'hc087c52e} /* (8, 10, 6) {real, imag} */,
  {32'hc0c635c0, 32'h3ecd7ea0} /* (8, 10, 5) {real, imag} */,
  {32'hc07f9347, 32'h3fd2b27b} /* (8, 10, 4) {real, imag} */,
  {32'hbedb29b0, 32'h3fb9ae44} /* (8, 10, 3) {real, imag} */,
  {32'hbf342418, 32'h4032b28c} /* (8, 10, 2) {real, imag} */,
  {32'hc07bde91, 32'hbf025ea8} /* (8, 10, 1) {real, imag} */,
  {32'hc043d8c9, 32'hc02ae403} /* (8, 10, 0) {real, imag} */,
  {32'hc0dacb94, 32'hc0dff0c2} /* (8, 9, 31) {real, imag} */,
  {32'hbfcae114, 32'hc0c229ca} /* (8, 9, 30) {real, imag} */,
  {32'hbf03144c, 32'hc11f45dc} /* (8, 9, 29) {real, imag} */,
  {32'h405c803a, 32'hc084973e} /* (8, 9, 28) {real, imag} */,
  {32'h3fbf4148, 32'h406a186c} /* (8, 9, 27) {real, imag} */,
  {32'hc10470c1, 32'h4044aaaa} /* (8, 9, 26) {real, imag} */,
  {32'hc065bcd0, 32'h40e05830} /* (8, 9, 25) {real, imag} */,
  {32'hbf01ed8c, 32'h40500c6e} /* (8, 9, 24) {real, imag} */,
  {32'h3e9825e0, 32'hc078c00c} /* (8, 9, 23) {real, imag} */,
  {32'h40a83ec4, 32'hc046a388} /* (8, 9, 22) {real, imag} */,
  {32'h40fca6e6, 32'hc01856d3} /* (8, 9, 21) {real, imag} */,
  {32'h4010f6ec, 32'hc0904d00} /* (8, 9, 20) {real, imag} */,
  {32'hc0580812, 32'hc01810e3} /* (8, 9, 19) {real, imag} */,
  {32'hc10e8ffe, 32'hc0b94711} /* (8, 9, 18) {real, imag} */,
  {32'hc082f3c4, 32'h40c20c56} /* (8, 9, 17) {real, imag} */,
  {32'hc0ba9104, 32'h40a8bc0d} /* (8, 9, 16) {real, imag} */,
  {32'hbf2d1e24, 32'h3f138340} /* (8, 9, 15) {real, imag} */,
  {32'h3fc225d0, 32'hbff6e2cc} /* (8, 9, 14) {real, imag} */,
  {32'h418d21ae, 32'h40285bb0} /* (8, 9, 13) {real, imag} */,
  {32'h40d0aac6, 32'hc0496a63} /* (8, 9, 12) {real, imag} */,
  {32'hbffe9118, 32'hc0649c88} /* (8, 9, 11) {real, imag} */,
  {32'h4002e5c2, 32'h40734bc4} /* (8, 9, 10) {real, imag} */,
  {32'hc0d60b86, 32'hbea98f90} /* (8, 9, 9) {real, imag} */,
  {32'hc08c29b4, 32'hc051796e} /* (8, 9, 8) {real, imag} */,
  {32'hc109fa5c, 32'h3e7c0ce0} /* (8, 9, 7) {real, imag} */,
  {32'hc0981b49, 32'h40924c7e} /* (8, 9, 6) {real, imag} */,
  {32'hc089735c, 32'h40b3dad2} /* (8, 9, 5) {real, imag} */,
  {32'hc1340ba1, 32'h3f664356} /* (8, 9, 4) {real, imag} */,
  {32'hc0a0ff2d, 32'h3f05b0c0} /* (8, 9, 3) {real, imag} */,
  {32'hc07691b5, 32'hc0f7a1b2} /* (8, 9, 2) {real, imag} */,
  {32'hc11247f2, 32'hc10c7a06} /* (8, 9, 1) {real, imag} */,
  {32'hc04a3284, 32'hc052192a} /* (8, 9, 0) {real, imag} */,
  {32'h40b8c350, 32'hc11247a5} /* (8, 8, 31) {real, imag} */,
  {32'h4010431c, 32'h414c907f} /* (8, 8, 30) {real, imag} */,
  {32'hbfce8650, 32'h41e50080} /* (8, 8, 29) {real, imag} */,
  {32'hc0ad7737, 32'h4153cc9e} /* (8, 8, 28) {real, imag} */,
  {32'h3fd5344c, 32'h4155f1a2} /* (8, 8, 27) {real, imag} */,
  {32'h416547ca, 32'h41793c26} /* (8, 8, 26) {real, imag} */,
  {32'h416d9b23, 32'hc01fbaf0} /* (8, 8, 25) {real, imag} */,
  {32'h410700b5, 32'hc1a7aa35} /* (8, 8, 24) {real, imag} */,
  {32'h40385566, 32'hbfc11ea5} /* (8, 8, 23) {real, imag} */,
  {32'h414b5562, 32'hbfa39cd8} /* (8, 8, 22) {real, imag} */,
  {32'h40bbcefd, 32'hc13b0079} /* (8, 8, 21) {real, imag} */,
  {32'hc05b71a3, 32'h3db757c0} /* (8, 8, 20) {real, imag} */,
  {32'hc0c51a69, 32'h405da0d8} /* (8, 8, 19) {real, imag} */,
  {32'h3fa4ddf8, 32'hc09d33fc} /* (8, 8, 18) {real, imag} */,
  {32'h3f7d0244, 32'hbfa10fbc} /* (8, 8, 17) {real, imag} */,
  {32'hc0512435, 32'h406def84} /* (8, 8, 16) {real, imag} */,
  {32'hc10ca20a, 32'hc0501e14} /* (8, 8, 15) {real, imag} */,
  {32'hc133915a, 32'h40a4fb9e} /* (8, 8, 14) {real, imag} */,
  {32'hc0dac662, 32'h4179928a} /* (8, 8, 13) {real, imag} */,
  {32'hc124db7f, 32'h40eab084} /* (8, 8, 12) {real, imag} */,
  {32'hc02a04f2, 32'h40de771f} /* (8, 8, 11) {real, imag} */,
  {32'h40c968df, 32'hc120702e} /* (8, 8, 10) {real, imag} */,
  {32'h4119d258, 32'hbe3286c0} /* (8, 8, 9) {real, imag} */,
  {32'h41358475, 32'hc0c86173} /* (8, 8, 8) {real, imag} */,
  {32'h413f51b9, 32'hc03b1a9e} /* (8, 8, 7) {real, imag} */,
  {32'h40ac8217, 32'hc098617e} /* (8, 8, 6) {real, imag} */,
  {32'hc11b77c7, 32'hc04ce56c} /* (8, 8, 5) {real, imag} */,
  {32'h400c7a5d, 32'hc0aee4a2} /* (8, 8, 4) {real, imag} */,
  {32'h3e819030, 32'h3fe5bb88} /* (8, 8, 3) {real, imag} */,
  {32'h3fae9838, 32'h400a1c3c} /* (8, 8, 2) {real, imag} */,
  {32'h4086274c, 32'hc11dd363} /* (8, 8, 1) {real, imag} */,
  {32'h40b1d973, 32'hc181d3b6} /* (8, 8, 0) {real, imag} */,
  {32'h3f4f64c4, 32'hbf8e4d4a} /* (8, 7, 31) {real, imag} */,
  {32'h409cac15, 32'hc0d5b532} /* (8, 7, 30) {real, imag} */,
  {32'h3ffcb12e, 32'hc123d92a} /* (8, 7, 29) {real, imag} */,
  {32'hbfa96b45, 32'hc108c84f} /* (8, 7, 28) {real, imag} */,
  {32'hbdd92b80, 32'hc084169a} /* (8, 7, 27) {real, imag} */,
  {32'h402b5184, 32'hc0881cc1} /* (8, 7, 26) {real, imag} */,
  {32'hbe5f84c0, 32'hc0fb0ea5} /* (8, 7, 25) {real, imag} */,
  {32'hc0635212, 32'h4023cc9c} /* (8, 7, 24) {real, imag} */,
  {32'hc099e7d2, 32'hbf0d6920} /* (8, 7, 23) {real, imag} */,
  {32'hc107f919, 32'hbe0037c0} /* (8, 7, 22) {real, imag} */,
  {32'hc11ac91e, 32'h41240961} /* (8, 7, 21) {real, imag} */,
  {32'h3e0c4830, 32'h4077e46f} /* (8, 7, 20) {real, imag} */,
  {32'h40d31794, 32'h4113f60f} /* (8, 7, 19) {real, imag} */,
  {32'h41190366, 32'h40894235} /* (8, 7, 18) {real, imag} */,
  {32'hc0257ae6, 32'hbfe10184} /* (8, 7, 17) {real, imag} */,
  {32'h4122b376, 32'h40afb32d} /* (8, 7, 16) {real, imag} */,
  {32'h4152d80e, 32'h4168b85a} /* (8, 7, 15) {real, imag} */,
  {32'h40152758, 32'h414df50d} /* (8, 7, 14) {real, imag} */,
  {32'h3f57acb4, 32'h41598d6e} /* (8, 7, 13) {real, imag} */,
  {32'hbf0d7314, 32'h414ee014} /* (8, 7, 12) {real, imag} */,
  {32'h40b30a2e, 32'hc087c982} /* (8, 7, 11) {real, imag} */,
  {32'hbe45a500, 32'h40b2cdec} /* (8, 7, 10) {real, imag} */,
  {32'h40535c41, 32'h41b9d7b0} /* (8, 7, 9) {real, imag} */,
  {32'h404d7c7e, 32'h418b889b} /* (8, 7, 8) {real, imag} */,
  {32'h41631fd0, 32'h40a544a5} /* (8, 7, 7) {real, imag} */,
  {32'h41637206, 32'h3f274828} /* (8, 7, 6) {real, imag} */,
  {32'h405ce4bc, 32'h3e9df8a0} /* (8, 7, 5) {real, imag} */,
  {32'h40d44536, 32'h4047db1a} /* (8, 7, 4) {real, imag} */,
  {32'h4012103e, 32'hc0b1409e} /* (8, 7, 3) {real, imag} */,
  {32'hc10994a3, 32'hc0f5fc78} /* (8, 7, 2) {real, imag} */,
  {32'hc15be6e4, 32'h3f544e98} /* (8, 7, 1) {real, imag} */,
  {32'hc0911e94, 32'h40aa33e2} /* (8, 7, 0) {real, imag} */,
  {32'h4035e45e, 32'h410abf44} /* (8, 6, 31) {real, imag} */,
  {32'h41413ef3, 32'h40975ff6} /* (8, 6, 30) {real, imag} */,
  {32'h41734d44, 32'hc08d64a2} /* (8, 6, 29) {real, imag} */,
  {32'h40ba24ba, 32'hbecbf8b8} /* (8, 6, 28) {real, imag} */,
  {32'hbfc1fe3c, 32'h40fbc006} /* (8, 6, 27) {real, imag} */,
  {32'h4042fe3e, 32'h40cbd6a2} /* (8, 6, 26) {real, imag} */,
  {32'hc0a17528, 32'hc0dd53c2} /* (8, 6, 25) {real, imag} */,
  {32'hc1651556, 32'hc183c64e} /* (8, 6, 24) {real, imag} */,
  {32'hc1268afb, 32'hbfc16928} /* (8, 6, 23) {real, imag} */,
  {32'hbfb1e91b, 32'hbfccf4b8} /* (8, 6, 22) {real, imag} */,
  {32'h4057577e, 32'hc0aaef01} /* (8, 6, 21) {real, imag} */,
  {32'h4045fa85, 32'hc0b9a3da} /* (8, 6, 20) {real, imag} */,
  {32'h41300e1e, 32'h40fb1bd1} /* (8, 6, 19) {real, imag} */,
  {32'h40c620d7, 32'h41062d19} /* (8, 6, 18) {real, imag} */,
  {32'hc0a968d0, 32'h40304864} /* (8, 6, 17) {real, imag} */,
  {32'hc1422c66, 32'hc105baf4} /* (8, 6, 16) {real, imag} */,
  {32'hc0e15b02, 32'hc006e91f} /* (8, 6, 15) {real, imag} */,
  {32'hc1131ede, 32'hbe9b8c80} /* (8, 6, 14) {real, imag} */,
  {32'hc0f45c07, 32'hbebd6140} /* (8, 6, 13) {real, imag} */,
  {32'hc19d9c10, 32'hc0a7a12c} /* (8, 6, 12) {real, imag} */,
  {32'hc0c77216, 32'hc1735a8c} /* (8, 6, 11) {real, imag} */,
  {32'hc10d30b4, 32'hc0a2398d} /* (8, 6, 10) {real, imag} */,
  {32'h4073d4bd, 32'h412a8a9e} /* (8, 6, 9) {real, imag} */,
  {32'h40ebcb9c, 32'h40a8783e} /* (8, 6, 8) {real, imag} */,
  {32'hc08c07e1, 32'hc0a9d324} /* (8, 6, 7) {real, imag} */,
  {32'hc10e49d2, 32'hc095c59c} /* (8, 6, 6) {real, imag} */,
  {32'h3e01f000, 32'hc1a9ef91} /* (8, 6, 5) {real, imag} */,
  {32'h4099b980, 32'hc12caf5c} /* (8, 6, 4) {real, imag} */,
  {32'h401470d1, 32'hbf9c0f4d} /* (8, 6, 3) {real, imag} */,
  {32'h412e6732, 32'hc00df2fc} /* (8, 6, 2) {real, imag} */,
  {32'h41215464, 32'hc0db37a4} /* (8, 6, 1) {real, imag} */,
  {32'h4102ce3d, 32'hc0fbcaa8} /* (8, 6, 0) {real, imag} */,
  {32'h416fc05a, 32'hbf0cefc8} /* (8, 5, 31) {real, imag} */,
  {32'h416bcaea, 32'hc0b5fe02} /* (8, 5, 30) {real, imag} */,
  {32'hc0844d9a, 32'hc19c40c9} /* (8, 5, 29) {real, imag} */,
  {32'hbf082138, 32'hc163377b} /* (8, 5, 28) {real, imag} */,
  {32'h40d73eae, 32'hbf0e6f60} /* (8, 5, 27) {real, imag} */,
  {32'h4192ab5d, 32'h4097aada} /* (8, 5, 26) {real, imag} */,
  {32'h4165df89, 32'h3fa231d6} /* (8, 5, 25) {real, imag} */,
  {32'h41aa95a0, 32'h40dcb010} /* (8, 5, 24) {real, imag} */,
  {32'h41fa97c3, 32'hc0f6607a} /* (8, 5, 23) {real, imag} */,
  {32'h416a2e7d, 32'hbf9a14c8} /* (8, 5, 22) {real, imag} */,
  {32'h4171a3e4, 32'hc00b6a5c} /* (8, 5, 21) {real, imag} */,
  {32'h40ed2ab4, 32'h3f90aec3} /* (8, 5, 20) {real, imag} */,
  {32'h4016d8f8, 32'h406e9b65} /* (8, 5, 19) {real, imag} */,
  {32'hbf6bc3ac, 32'h3d88a560} /* (8, 5, 18) {real, imag} */,
  {32'hc0821a1f, 32'hbff66c9d} /* (8, 5, 17) {real, imag} */,
  {32'hc11509b0, 32'h40d74050} /* (8, 5, 16) {real, imag} */,
  {32'hc116be1f, 32'h40ff1118} /* (8, 5, 15) {real, imag} */,
  {32'hc0401a34, 32'h40b500de} /* (8, 5, 14) {real, imag} */,
  {32'hbfc1d153, 32'h40d0567e} /* (8, 5, 13) {real, imag} */,
  {32'hc1011cbe, 32'hc11a766a} /* (8, 5, 12) {real, imag} */,
  {32'hc13d0b2e, 32'hc137deaf} /* (8, 5, 11) {real, imag} */,
  {32'hc0ffae0a, 32'hc0da45ed} /* (8, 5, 10) {real, imag} */,
  {32'hc0455f8e, 32'hc0259fc2} /* (8, 5, 9) {real, imag} */,
  {32'h4130d43b, 32'hc05d6c76} /* (8, 5, 8) {real, imag} */,
  {32'h413d122a, 32'h40c97e68} /* (8, 5, 7) {real, imag} */,
  {32'h4136c385, 32'h400590c6} /* (8, 5, 6) {real, imag} */,
  {32'h40649321, 32'hc162168e} /* (8, 5, 5) {real, imag} */,
  {32'h4098f022, 32'hc0cd3ed8} /* (8, 5, 4) {real, imag} */,
  {32'h406c59d8, 32'hc0bca82a} /* (8, 5, 3) {real, imag} */,
  {32'hc0660d1a, 32'hc144918e} /* (8, 5, 2) {real, imag} */,
  {32'h4152fa75, 32'hc0c0bbdf} /* (8, 5, 1) {real, imag} */,
  {32'h41a60722, 32'hbfb5c6fa} /* (8, 5, 0) {real, imag} */,
  {32'hbffb501d, 32'hbf98c608} /* (8, 4, 31) {real, imag} */,
  {32'hbfb5c300, 32'h40ef1f2e} /* (8, 4, 30) {real, imag} */,
  {32'hc0292be6, 32'h4108603e} /* (8, 4, 29) {real, imag} */,
  {32'hc096a9d8, 32'hbf6e8d58} /* (8, 4, 28) {real, imag} */,
  {32'hc0967b98, 32'h41291af3} /* (8, 4, 27) {real, imag} */,
  {32'hbf8e52dc, 32'h400db913} /* (8, 4, 26) {real, imag} */,
  {32'hc15fdae0, 32'h3f640b58} /* (8, 4, 25) {real, imag} */,
  {32'hc0ada2e6, 32'hc06883f8} /* (8, 4, 24) {real, imag} */,
  {32'hc1826e03, 32'hbf1e1a78} /* (8, 4, 23) {real, imag} */,
  {32'hc1592050, 32'h418a4425} /* (8, 4, 22) {real, imag} */,
  {32'h413a3165, 32'h40f21fdd} /* (8, 4, 21) {real, imag} */,
  {32'h41e67186, 32'hc045e92a} /* (8, 4, 20) {real, imag} */,
  {32'h419a8884, 32'h3ec8fc54} /* (8, 4, 19) {real, imag} */,
  {32'h41c39719, 32'h410bd44e} /* (8, 4, 18) {real, imag} */,
  {32'h41e69496, 32'h40a804c4} /* (8, 4, 17) {real, imag} */,
  {32'h41cd7cba, 32'hc193a0cc} /* (8, 4, 16) {real, imag} */,
  {32'hc03dc0b3, 32'hc1b24a47} /* (8, 4, 15) {real, imag} */,
  {32'hc083060e, 32'h408543e8} /* (8, 4, 14) {real, imag} */,
  {32'h411d2a09, 32'h4137a93c} /* (8, 4, 13) {real, imag} */,
  {32'h415484ac, 32'h3eacdce0} /* (8, 4, 12) {real, imag} */,
  {32'hc0b666b4, 32'hc0485ee4} /* (8, 4, 11) {real, imag} */,
  {32'hc10962dc, 32'hc18165af} /* (8, 4, 10) {real, imag} */,
  {32'hc090d050, 32'hc05590d7} /* (8, 4, 9) {real, imag} */,
  {32'hc1a12206, 32'h407feeb4} /* (8, 4, 8) {real, imag} */,
  {32'hc1b1dce4, 32'h4087bd1b} /* (8, 4, 7) {real, imag} */,
  {32'hc1cf7dba, 32'hc112e52c} /* (8, 4, 6) {real, imag} */,
  {32'hc1a3dcf8, 32'hc0ac37a8} /* (8, 4, 5) {real, imag} */,
  {32'hc1199b2f, 32'hbfce5390} /* (8, 4, 4) {real, imag} */,
  {32'hc1094e54, 32'h400975b8} /* (8, 4, 3) {real, imag} */,
  {32'h40070140, 32'h411ff2b6} /* (8, 4, 2) {real, imag} */,
  {32'h40ee86e8, 32'hc1942f54} /* (8, 4, 1) {real, imag} */,
  {32'h4097d20c, 32'hc181fa65} /* (8, 4, 0) {real, imag} */,
  {32'hc00e0d9e, 32'hc09bc08a} /* (8, 3, 31) {real, imag} */,
  {32'hbfa1feba, 32'hc16630a0} /* (8, 3, 30) {real, imag} */,
  {32'hbdc995c0, 32'hc12e05f4} /* (8, 3, 29) {real, imag} */,
  {32'hc11018b5, 32'h4091274f} /* (8, 3, 28) {real, imag} */,
  {32'hc0f5c4bb, 32'hc05fff74} /* (8, 3, 27) {real, imag} */,
  {32'hc0a38e4e, 32'h3fb62d2f} /* (8, 3, 26) {real, imag} */,
  {32'hc1a5b83f, 32'h40268188} /* (8, 3, 25) {real, imag} */,
  {32'h411ab858, 32'hc0f3609e} /* (8, 3, 24) {real, imag} */,
  {32'h4143d964, 32'hc184653c} /* (8, 3, 23) {real, imag} */,
  {32'hc110f420, 32'hc0722948} /* (8, 3, 22) {real, imag} */,
  {32'hbfcf59e0, 32'h4144f4a3} /* (8, 3, 21) {real, imag} */,
  {32'h41945cde, 32'h4156aaea} /* (8, 3, 20) {real, imag} */,
  {32'h41e11a84, 32'hc0332c3a} /* (8, 3, 19) {real, imag} */,
  {32'h411660ae, 32'h4193ee50} /* (8, 3, 18) {real, imag} */,
  {32'hbffd99b8, 32'h41366f14} /* (8, 3, 17) {real, imag} */,
  {32'h415131e9, 32'h411ae5ab} /* (8, 3, 16) {real, imag} */,
  {32'hbf3d1e2c, 32'hc0226870} /* (8, 3, 15) {real, imag} */,
  {32'h3fbb62ac, 32'hc017799a} /* (8, 3, 14) {real, imag} */,
  {32'h3f8a10e4, 32'hc14e646f} /* (8, 3, 13) {real, imag} */,
  {32'h4050d81c, 32'hc12aab44} /* (8, 3, 12) {real, imag} */,
  {32'h4080ccd5, 32'hbfa130e6} /* (8, 3, 11) {real, imag} */,
  {32'h3f8c8526, 32'h4032933e} /* (8, 3, 10) {real, imag} */,
  {32'hc15a23e7, 32'h3eb19654} /* (8, 3, 9) {real, imag} */,
  {32'hc1c6e2b4, 32'hc1357684} /* (8, 3, 8) {real, imag} */,
  {32'hc17f04f6, 32'hc0e1ddf0} /* (8, 3, 7) {real, imag} */,
  {32'hc12aa348, 32'hc0722c98} /* (8, 3, 6) {real, imag} */,
  {32'hc1e1810f, 32'hc12b901c} /* (8, 3, 5) {real, imag} */,
  {32'hc1a118fe, 32'hc0dc7054} /* (8, 3, 4) {real, imag} */,
  {32'h4112d3cf, 32'hc09bda9b} /* (8, 3, 3) {real, imag} */,
  {32'hc02b6cc7, 32'h3f4de4bc} /* (8, 3, 2) {real, imag} */,
  {32'h3e428de0, 32'h3f9e2225} /* (8, 3, 1) {real, imag} */,
  {32'hbff0c0b3, 32'hc01922b0} /* (8, 3, 0) {real, imag} */,
  {32'h4191debf, 32'hc17fe5f8} /* (8, 2, 31) {real, imag} */,
  {32'h41a2d021, 32'hc2010882} /* (8, 2, 30) {real, imag} */,
  {32'h41b12854, 32'hc1e6ac6c} /* (8, 2, 29) {real, imag} */,
  {32'h41964d49, 32'hbf3b18a0} /* (8, 2, 28) {real, imag} */,
  {32'h41e30bf2, 32'hc181c38e} /* (8, 2, 27) {real, imag} */,
  {32'h41c7cc44, 32'hc1bf224a} /* (8, 2, 26) {real, imag} */,
  {32'h41a6087a, 32'hc1a153ea} /* (8, 2, 25) {real, imag} */,
  {32'h418ad810, 32'hc167721f} /* (8, 2, 24) {real, imag} */,
  {32'h419e3c28, 32'hc122027e} /* (8, 2, 23) {real, imag} */,
  {32'h41a089f3, 32'hc12771bd} /* (8, 2, 22) {real, imag} */,
  {32'h40b4fd76, 32'hbf189ae0} /* (8, 2, 21) {real, imag} */,
  {32'hc18be2ac, 32'h41917162} /* (8, 2, 20) {real, imag} */,
  {32'hc17b0c7c, 32'h41d6631d} /* (8, 2, 19) {real, imag} */,
  {32'hc0f7b98a, 32'h420bc0ba} /* (8, 2, 18) {real, imag} */,
  {32'hc1558fcc, 32'h421e57e5} /* (8, 2, 17) {real, imag} */,
  {32'hc1841843, 32'h4214495a} /* (8, 2, 16) {real, imag} */,
  {32'hc1c881cb, 32'h419498c0} /* (8, 2, 15) {real, imag} */,
  {32'hc200515a, 32'hbf7dbc08} /* (8, 2, 14) {real, imag} */,
  {32'hc1bf4ced, 32'h40af8c7c} /* (8, 2, 13) {real, imag} */,
  {32'hc1d2a8ea, 32'h40b896f2} /* (8, 2, 12) {real, imag} */,
  {32'hc157d21c, 32'h412d8bac} /* (8, 2, 11) {real, imag} */,
  {32'h41a1b907, 32'hc1a5c87d} /* (8, 2, 10) {real, imag} */,
  {32'h41c9bdea, 32'hc213dd1c} /* (8, 2, 9) {real, imag} */,
  {32'h41b28ce9, 32'hc2121567} /* (8, 2, 8) {real, imag} */,
  {32'h41ad4922, 32'hc1e7e40a} /* (8, 2, 7) {real, imag} */,
  {32'h41e06e3f, 32'hc1e7a3c2} /* (8, 2, 6) {real, imag} */,
  {32'h41eab1a6, 32'hc18ba88a} /* (8, 2, 5) {real, imag} */,
  {32'h41fbcc92, 32'hc013cb28} /* (8, 2, 4) {real, imag} */,
  {32'h41e86b3d, 32'hc057ed94} /* (8, 2, 3) {real, imag} */,
  {32'h42052300, 32'hc0ae2f34} /* (8, 2, 2) {real, imag} */,
  {32'h4220b839, 32'hc1c6d656} /* (8, 2, 1) {real, imag} */,
  {32'h41485167, 32'hc19cf720} /* (8, 2, 0) {real, imag} */,
  {32'hc18776b6, 32'h3ff98fd8} /* (8, 1, 31) {real, imag} */,
  {32'hc1e52462, 32'h416a7df0} /* (8, 1, 30) {real, imag} */,
  {32'hc22818f8, 32'h4195aca4} /* (8, 1, 29) {real, imag} */,
  {32'hc221e600, 32'h41df4313} /* (8, 1, 28) {real, imag} */,
  {32'hc23d944f, 32'h41b259de} /* (8, 1, 27) {real, imag} */,
  {32'hc1d4efaf, 32'h41bc2582} /* (8, 1, 26) {real, imag} */,
  {32'hc1556465, 32'h41bb1037} /* (8, 1, 25) {real, imag} */,
  {32'hc20f34f7, 32'h410402dc} /* (8, 1, 24) {real, imag} */,
  {32'hc20a9a31, 32'h41e84aad} /* (8, 1, 23) {real, imag} */,
  {32'hc207e15a, 32'h423d112f} /* (8, 1, 22) {real, imag} */,
  {32'hc172c596, 32'h42176e1a} /* (8, 1, 21) {real, imag} */,
  {32'h41a583a3, 32'h41c5259a} /* (8, 1, 20) {real, imag} */,
  {32'h41ebe5c8, 32'h4073d96d} /* (8, 1, 19) {real, imag} */,
  {32'h41be4688, 32'hbfc4c910} /* (8, 1, 18) {real, imag} */,
  {32'h41d7f516, 32'hc085e818} /* (8, 1, 17) {real, imag} */,
  {32'h421c97f4, 32'hc1b96738} /* (8, 1, 16) {real, imag} */,
  {32'h420c96db, 32'hc20a9f77} /* (8, 1, 15) {real, imag} */,
  {32'h41e4f6dd, 32'hc2170e2c} /* (8, 1, 14) {real, imag} */,
  {32'h41bd9500, 32'hc1b43b7a} /* (8, 1, 13) {real, imag} */,
  {32'h423ebe7c, 32'hc1b7ad9b} /* (8, 1, 12) {real, imag} */,
  {32'h4231cf12, 32'hc1a3b6c0} /* (8, 1, 11) {real, imag} */,
  {32'hc15d6eef, 32'h40170510} /* (8, 1, 10) {real, imag} */,
  {32'hc1afd198, 32'h3eb7bb80} /* (8, 1, 9) {real, imag} */,
  {32'hc10e9e88, 32'hc118a037} /* (8, 1, 8) {real, imag} */,
  {32'hc0fb7be6, 32'h4115518a} /* (8, 1, 7) {real, imag} */,
  {32'hc1a167bb, 32'h419f9278} /* (8, 1, 6) {real, imag} */,
  {32'hc20f5c72, 32'h41c83815} /* (8, 1, 5) {real, imag} */,
  {32'hc206ff52, 32'h4220dd07} /* (8, 1, 4) {real, imag} */,
  {32'hc20e6312, 32'h420088d8} /* (8, 1, 3) {real, imag} */,
  {32'hc19449da, 32'h42251a58} /* (8, 1, 2) {real, imag} */,
  {32'hc1b7ea06, 32'h42222905} /* (8, 1, 1) {real, imag} */,
  {32'hc1deca3f, 32'h4117a0d4} /* (8, 1, 0) {real, imag} */,
  {32'hc1118b00, 32'h4107657b} /* (8, 0, 31) {real, imag} */,
  {32'hc17b727b, 32'h4189bc94} /* (8, 0, 30) {real, imag} */,
  {32'hc1b32ad5, 32'h414d018f} /* (8, 0, 29) {real, imag} */,
  {32'hc203628e, 32'h41f7cd86} /* (8, 0, 28) {real, imag} */,
  {32'hc192049e, 32'h41d104bf} /* (8, 0, 27) {real, imag} */,
  {32'hc1789628, 32'h41585b1c} /* (8, 0, 26) {real, imag} */,
  {32'hc0962602, 32'h4096ec7b} /* (8, 0, 25) {real, imag} */,
  {32'hc19177f9, 32'h3f5f72cc} /* (8, 0, 24) {real, imag} */,
  {32'hc1940360, 32'h40ac12d0} /* (8, 0, 23) {real, imag} */,
  {32'hc1855953, 32'h418bdce0} /* (8, 0, 22) {real, imag} */,
  {32'h40355732, 32'h41c3a660} /* (8, 0, 21) {real, imag} */,
  {32'h408d3f0e, 32'hc1cf5e0b} /* (8, 0, 20) {real, imag} */,
  {32'hc1261695, 32'hc12b6513} /* (8, 0, 19) {real, imag} */,
  {32'h3f565e64, 32'h418138ee} /* (8, 0, 18) {real, imag} */,
  {32'hbfad1102, 32'h41208cc8} /* (8, 0, 17) {real, imag} */,
  {32'h40745659, 32'hc0ea816b} /* (8, 0, 16) {real, imag} */,
  {32'h417fc145, 32'hc1a73eb4} /* (8, 0, 15) {real, imag} */,
  {32'h420be86f, 32'hc13b3b00} /* (8, 0, 14) {real, imag} */,
  {32'h41e65396, 32'hc15db0b8} /* (8, 0, 13) {real, imag} */,
  {32'h41d01d13, 32'hc189f413} /* (8, 0, 12) {real, imag} */,
  {32'h41e079ac, 32'hc1c251f4} /* (8, 0, 11) {real, imag} */,
  {32'h417373d7, 32'hc137e11c} /* (8, 0, 10) {real, imag} */,
  {32'hc00dad29, 32'h415d8e6a} /* (8, 0, 9) {real, imag} */,
  {32'hc132a338, 32'h410d2dc3} /* (8, 0, 8) {real, imag} */,
  {32'hc115051c, 32'h3e08e690} /* (8, 0, 7) {real, imag} */,
  {32'hc15d7dd2, 32'h3e2c3a70} /* (8, 0, 6) {real, imag} */,
  {32'hc0baa78c, 32'h414e7980} /* (8, 0, 5) {real, imag} */,
  {32'hbfd17c80, 32'h41c1bd62} /* (8, 0, 4) {real, imag} */,
  {32'hc19bb871, 32'h41b0865c} /* (8, 0, 3) {real, imag} */,
  {32'hc1966352, 32'h41e917d2} /* (8, 0, 2) {real, imag} */,
  {32'hc17b5bdd, 32'h41d28430} /* (8, 0, 1) {real, imag} */,
  {32'hc1a6020b, 32'h419189cc} /* (8, 0, 0) {real, imag} */,
  {32'hc0e0e5cc, 32'h40a457f7} /* (7, 31, 31) {real, imag} */,
  {32'h4074efa0, 32'hc0a949ec} /* (7, 31, 30) {real, imag} */,
  {32'h40d97437, 32'hbeb5fcc0} /* (7, 31, 29) {real, imag} */,
  {32'h416b33c0, 32'h3ea9f2d8} /* (7, 31, 28) {real, imag} */,
  {32'h41b61037, 32'h4081b3a0} /* (7, 31, 27) {real, imag} */,
  {32'h40809787, 32'h40f511d8} /* (7, 31, 26) {real, imag} */,
  {32'hbf92ba17, 32'hc09b7c38} /* (7, 31, 25) {real, imag} */,
  {32'hc0a4d1f0, 32'hc15e3fbb} /* (7, 31, 24) {real, imag} */,
  {32'hc08e7f52, 32'hc073e4c3} /* (7, 31, 23) {real, imag} */,
  {32'hc0ff81b6, 32'h40a5ce24} /* (7, 31, 22) {real, imag} */,
  {32'hc10723f3, 32'h3f7ea398} /* (7, 31, 21) {real, imag} */,
  {32'h40c03574, 32'hc11b051a} /* (7, 31, 20) {real, imag} */,
  {32'hbe319700, 32'hbe3a6f00} /* (7, 31, 19) {real, imag} */,
  {32'hc1346a69, 32'h4078b12c} /* (7, 31, 18) {real, imag} */,
  {32'h407223f3, 32'hc0cdc87a} /* (7, 31, 17) {real, imag} */,
  {32'h415747bb, 32'h40441250} /* (7, 31, 16) {real, imag} */,
  {32'h407de58a, 32'h414f746c} /* (7, 31, 15) {real, imag} */,
  {32'hbff49380, 32'h41123c5d} /* (7, 31, 14) {real, imag} */,
  {32'hc093d80a, 32'h4103859a} /* (7, 31, 13) {real, imag} */,
  {32'hc0271194, 32'h41c7d66a} /* (7, 31, 12) {real, imag} */,
  {32'hc15dce3d, 32'h41487a94} /* (7, 31, 11) {real, imag} */,
  {32'hc1b9bf70, 32'hc1dcc25d} /* (7, 31, 10) {real, imag} */,
  {32'hc19cb931, 32'hc220156e} /* (7, 31, 9) {real, imag} */,
  {32'hc19b0f46, 32'hc1f86cf1} /* (7, 31, 8) {real, imag} */,
  {32'hc11c8bdc, 32'hc1c09a8f} /* (7, 31, 7) {real, imag} */,
  {32'hc0ca73ec, 32'hc07cd1bd} /* (7, 31, 6) {real, imag} */,
  {32'hc0bb3fa8, 32'h415bb8be} /* (7, 31, 5) {real, imag} */,
  {32'hc0531908, 32'h3f17cdfc} /* (7, 31, 4) {real, imag} */,
  {32'hc05eecf6, 32'hc08215bd} /* (7, 31, 3) {real, imag} */,
  {32'h4104a093, 32'hc1293bcb} /* (7, 31, 2) {real, imag} */,
  {32'hc13829f4, 32'hc161427e} /* (7, 31, 1) {real, imag} */,
  {32'hc109e4ae, 32'h4056bbae} /* (7, 31, 0) {real, imag} */,
  {32'hc022eee5, 32'h3fd0bae0} /* (7, 30, 31) {real, imag} */,
  {32'h417e1db0, 32'h41cca9de} /* (7, 30, 30) {real, imag} */,
  {32'h3f0d9fc4, 32'h4160e8bc} /* (7, 30, 29) {real, imag} */,
  {32'h403f19fd, 32'hc0a1e30c} /* (7, 30, 28) {real, imag} */,
  {32'h41140232, 32'h40e57b72} /* (7, 30, 27) {real, imag} */,
  {32'h40010414, 32'h41917d8d} /* (7, 30, 26) {real, imag} */,
  {32'h408c0d68, 32'hbfd03428} /* (7, 30, 25) {real, imag} */,
  {32'hc0abe48c, 32'hc0bdf110} /* (7, 30, 24) {real, imag} */,
  {32'hc0c7203e, 32'hc0f51d54} /* (7, 30, 23) {real, imag} */,
  {32'hc14f7b02, 32'hc16ba605} /* (7, 30, 22) {real, imag} */,
  {32'h4094360e, 32'hbf811954} /* (7, 30, 21) {real, imag} */,
  {32'h4133d41c, 32'h412d34f0} /* (7, 30, 20) {real, imag} */,
  {32'hc089770c, 32'h41341816} /* (7, 30, 19) {real, imag} */,
  {32'hc18185bf, 32'hc0d19e78} /* (7, 30, 18) {real, imag} */,
  {32'hbfe7dad0, 32'hc0b74ba5} /* (7, 30, 17) {real, imag} */,
  {32'hc0c52d8d, 32'h41068d2c} /* (7, 30, 16) {real, imag} */,
  {32'hc1b71dcc, 32'h41831777} /* (7, 30, 15) {real, imag} */,
  {32'hc0ff146c, 32'h419f973b} /* (7, 30, 14) {real, imag} */,
  {32'h4099aa24, 32'h4077befa} /* (7, 30, 13) {real, imag} */,
  {32'h4116de18, 32'h3e9487d0} /* (7, 30, 12) {real, imag} */,
  {32'h40c0644d, 32'h4065a799} /* (7, 30, 11) {real, imag} */,
  {32'hc08fb7d1, 32'h410d6a80} /* (7, 30, 10) {real, imag} */,
  {32'hc106c47a, 32'hc030a5cf} /* (7, 30, 9) {real, imag} */,
  {32'hbf4885c0, 32'hc028bcdc} /* (7, 30, 8) {real, imag} */,
  {32'h3e02ba80, 32'h3e771230} /* (7, 30, 7) {real, imag} */,
  {32'hc13e44af, 32'h414f041c} /* (7, 30, 6) {real, imag} */,
  {32'hc1ec96eb, 32'h41fa83d9} /* (7, 30, 5) {real, imag} */,
  {32'hbfc0ab54, 32'h41f39280} /* (7, 30, 4) {real, imag} */,
  {32'h3d996400, 32'h41cdd31c} /* (7, 30, 3) {real, imag} */,
  {32'hc0301b48, 32'h40cd6eda} /* (7, 30, 2) {real, imag} */,
  {32'hc08c046e, 32'h4066575c} /* (7, 30, 1) {real, imag} */,
  {32'hbfec9580, 32'h40aae562} /* (7, 30, 0) {real, imag} */,
  {32'hc0192314, 32'h40a97ef0} /* (7, 29, 31) {real, imag} */,
  {32'hc1072cdd, 32'hc0aacca6} /* (7, 29, 30) {real, imag} */,
  {32'hc0cbd474, 32'hc103ec8c} /* (7, 29, 29) {real, imag} */,
  {32'h3f899390, 32'hc0aa3d99} /* (7, 29, 28) {real, imag} */,
  {32'hc11f72c6, 32'h40a42e56} /* (7, 29, 27) {real, imag} */,
  {32'hc0390a61, 32'h405c6800} /* (7, 29, 26) {real, imag} */,
  {32'h3f61a118, 32'h409ae220} /* (7, 29, 25) {real, imag} */,
  {32'hc00bacec, 32'h419ab9fb} /* (7, 29, 24) {real, imag} */,
  {32'hc033eb88, 32'h40b3d3ab} /* (7, 29, 23) {real, imag} */,
  {32'hc069723e, 32'hc08c7a04} /* (7, 29, 22) {real, imag} */,
  {32'hc116e09c, 32'h3fdcbaa0} /* (7, 29, 21) {real, imag} */,
  {32'hc113ce38, 32'h414e0216} /* (7, 29, 20) {real, imag} */,
  {32'h406433a6, 32'h411b333d} /* (7, 29, 19) {real, imag} */,
  {32'h410cf0ea, 32'hc037e36c} /* (7, 29, 18) {real, imag} */,
  {32'hc0ac80a5, 32'h402ba9b8} /* (7, 29, 17) {real, imag} */,
  {32'hc14a94fb, 32'hc12c7581} /* (7, 29, 16) {real, imag} */,
  {32'hc18c10fc, 32'hc082c180} /* (7, 29, 15) {real, imag} */,
  {32'hc18841cf, 32'hbf1928f8} /* (7, 29, 14) {real, imag} */,
  {32'hc04d8a05, 32'hc026e00a} /* (7, 29, 13) {real, imag} */,
  {32'h41953561, 32'hc06aad7e} /* (7, 29, 12) {real, imag} */,
  {32'h402b83fc, 32'h3e48d940} /* (7, 29, 11) {real, imag} */,
  {32'hc168f3b7, 32'h40c8de2e} /* (7, 29, 10) {real, imag} */,
  {32'hc184e911, 32'hc14584b2} /* (7, 29, 9) {real, imag} */,
  {32'h4064204c, 32'hc12f01d9} /* (7, 29, 8) {real, imag} */,
  {32'hbf43c7e4, 32'hc14a6772} /* (7, 29, 7) {real, imag} */,
  {32'h3fccf880, 32'h418cb043} /* (7, 29, 6) {real, imag} */,
  {32'h40f6c105, 32'h41e2dad3} /* (7, 29, 5) {real, imag} */,
  {32'hbfd3282c, 32'h413122c2} /* (7, 29, 4) {real, imag} */,
  {32'hc10fb241, 32'hbf7e2970} /* (7, 29, 3) {real, imag} */,
  {32'hc0c186f9, 32'hc00e4bc3} /* (7, 29, 2) {real, imag} */,
  {32'hc186fc36, 32'h4045a898} /* (7, 29, 1) {real, imag} */,
  {32'hc170e8f5, 32'h414b33ae} /* (7, 29, 0) {real, imag} */,
  {32'hc11f12cd, 32'hc0bc33a4} /* (7, 28, 31) {real, imag} */,
  {32'hc0cf12ec, 32'hbf202890} /* (7, 28, 30) {real, imag} */,
  {32'h41659755, 32'hc0d44dce} /* (7, 28, 29) {real, imag} */,
  {32'hc02a9783, 32'hc000fc5c} /* (7, 28, 28) {real, imag} */,
  {32'hc197c9b8, 32'h3fb25b88} /* (7, 28, 27) {real, imag} */,
  {32'hc187fdef, 32'hc0f03e5f} /* (7, 28, 26) {real, imag} */,
  {32'hc0a334e0, 32'hc0a263b2} /* (7, 28, 25) {real, imag} */,
  {32'h3f5385c2, 32'h401ad332} /* (7, 28, 24) {real, imag} */,
  {32'h4088abd6, 32'hc1255eb5} /* (7, 28, 23) {real, imag} */,
  {32'h41899569, 32'hc06280e0} /* (7, 28, 22) {real, imag} */,
  {32'hc07902fc, 32'hc016b929} /* (7, 28, 21) {real, imag} */,
  {32'hc195a336, 32'hc0b20c98} /* (7, 28, 20) {real, imag} */,
  {32'h3ee1d1c0, 32'h3e9dbcc8} /* (7, 28, 19) {real, imag} */,
  {32'h41845225, 32'hc0e42273} /* (7, 28, 18) {real, imag} */,
  {32'h418ca415, 32'hc145b961} /* (7, 28, 17) {real, imag} */,
  {32'h402169d0, 32'hc01a2170} /* (7, 28, 16) {real, imag} */,
  {32'h3e9f86e0, 32'hc054f15c} /* (7, 28, 15) {real, imag} */,
  {32'hc132a8ee, 32'hc0ac6bbc} /* (7, 28, 14) {real, imag} */,
  {32'hc0fc658c, 32'h4023609a} /* (7, 28, 13) {real, imag} */,
  {32'hc0066fb4, 32'hbf658698} /* (7, 28, 12) {real, imag} */,
  {32'hc01419e9, 32'hc1b6bf1f} /* (7, 28, 11) {real, imag} */,
  {32'h41220e02, 32'hc12f418e} /* (7, 28, 10) {real, imag} */,
  {32'h4173b307, 32'h3d7f0a00} /* (7, 28, 9) {real, imag} */,
  {32'h3fe8ef22, 32'hbf88df5f} /* (7, 28, 8) {real, imag} */,
  {32'h41920fc0, 32'hc086982c} /* (7, 28, 7) {real, imag} */,
  {32'h41592718, 32'h401730cd} /* (7, 28, 6) {real, imag} */,
  {32'hc0a8b408, 32'hc01ba29e} /* (7, 28, 5) {real, imag} */,
  {32'hc0f661eb, 32'h400388fe} /* (7, 28, 4) {real, imag} */,
  {32'hc0c158c0, 32'hc067d4b5} /* (7, 28, 3) {real, imag} */,
  {32'h4067b0d1, 32'hc0cbc584} /* (7, 28, 2) {real, imag} */,
  {32'h41271691, 32'hc0cc1cfb} /* (7, 28, 1) {real, imag} */,
  {32'h3fcef09a, 32'hbf6e67b0} /* (7, 28, 0) {real, imag} */,
  {32'hc04c7cce, 32'h408eae46} /* (7, 27, 31) {real, imag} */,
  {32'hbfa51fb6, 32'h4003ed84} /* (7, 27, 30) {real, imag} */,
  {32'h40214a96, 32'h419ae5fc} /* (7, 27, 29) {real, imag} */,
  {32'h409b642c, 32'h4158b7f3} /* (7, 27, 28) {real, imag} */,
  {32'hc107c19d, 32'h401ad848} /* (7, 27, 27) {real, imag} */,
  {32'hc189569d, 32'hc0bde6c6} /* (7, 27, 26) {real, imag} */,
  {32'hc1905fff, 32'h40ce9a07} /* (7, 27, 25) {real, imag} */,
  {32'hc19bd9c1, 32'h417860f3} /* (7, 27, 24) {real, imag} */,
  {32'h41118e34, 32'hbe678280} /* (7, 27, 23) {real, imag} */,
  {32'h41cd80f8, 32'h40123e7c} /* (7, 27, 22) {real, imag} */,
  {32'h41a1d816, 32'hc05fd0e6} /* (7, 27, 21) {real, imag} */,
  {32'h3fbd5943, 32'hc12bd755} /* (7, 27, 20) {real, imag} */,
  {32'h3ffaff74, 32'h4113e42a} /* (7, 27, 19) {real, imag} */,
  {32'h411f0a6e, 32'h41594abc} /* (7, 27, 18) {real, imag} */,
  {32'hc01f4e18, 32'hc077cd9c} /* (7, 27, 17) {real, imag} */,
  {32'h3f8e4888, 32'hc071a4bf} /* (7, 27, 16) {real, imag} */,
  {32'h418c5b56, 32'hc03296be} /* (7, 27, 15) {real, imag} */,
  {32'h4126dc7c, 32'h4085001c} /* (7, 27, 14) {real, imag} */,
  {32'hc0028743, 32'h4194d5ac} /* (7, 27, 13) {real, imag} */,
  {32'h41259a8e, 32'h4125a1ae} /* (7, 27, 12) {real, imag} */,
  {32'h416da4f2, 32'h403bd2f4} /* (7, 27, 11) {real, imag} */,
  {32'hbfcc8bbd, 32'hc092b012} /* (7, 27, 10) {real, imag} */,
  {32'h4020cc18, 32'h406c2d54} /* (7, 27, 9) {real, imag} */,
  {32'h414f7e67, 32'h40e50a40} /* (7, 27, 8) {real, imag} */,
  {32'h41c5f13d, 32'h4106efd2} /* (7, 27, 7) {real, imag} */,
  {32'h4196839a, 32'h3faebfe0} /* (7, 27, 6) {real, imag} */,
  {32'h4184439c, 32'hc060f7d2} /* (7, 27, 5) {real, imag} */,
  {32'h40bfd8e6, 32'h403b6d8b} /* (7, 27, 4) {real, imag} */,
  {32'hc13e0cf7, 32'hc090522d} /* (7, 27, 3) {real, imag} */,
  {32'hc126964e, 32'hc110e48d} /* (7, 27, 2) {real, imag} */,
  {32'hc0d0f8a3, 32'h3f49cf48} /* (7, 27, 1) {real, imag} */,
  {32'hc0a222a2, 32'h4105a539} /* (7, 27, 0) {real, imag} */,
  {32'h3e50f450, 32'h3ef58ee0} /* (7, 26, 31) {real, imag} */,
  {32'h3eed3d0c, 32'h40571277} /* (7, 26, 30) {real, imag} */,
  {32'hc0f1a01c, 32'hbf89aeca} /* (7, 26, 29) {real, imag} */,
  {32'hc09708a0, 32'h418425e4} /* (7, 26, 28) {real, imag} */,
  {32'h3fc95c26, 32'h40b50522} /* (7, 26, 27) {real, imag} */,
  {32'h40012360, 32'hc00fc35a} /* (7, 26, 26) {real, imag} */,
  {32'h40ac4cc4, 32'hc10e29fa} /* (7, 26, 25) {real, imag} */,
  {32'hc0dec26e, 32'hc197c51e} /* (7, 26, 24) {real, imag} */,
  {32'hc117d810, 32'h3fd0c2c2} /* (7, 26, 23) {real, imag} */,
  {32'hc0a2ebf3, 32'hc09330be} /* (7, 26, 22) {real, imag} */,
  {32'hc0b430aa, 32'h4161c35d} /* (7, 26, 21) {real, imag} */,
  {32'h3f8515a4, 32'h40644597} /* (7, 26, 20) {real, imag} */,
  {32'h41294084, 32'hc13b0707} /* (7, 26, 19) {real, imag} */,
  {32'h406972ac, 32'h3f337c48} /* (7, 26, 18) {real, imag} */,
  {32'h3fbb52ff, 32'h404b0f51} /* (7, 26, 17) {real, imag} */,
  {32'h3eb74458, 32'hc10f29d0} /* (7, 26, 16) {real, imag} */,
  {32'h3f16f068, 32'hc173c02e} /* (7, 26, 15) {real, imag} */,
  {32'h3fb37ce0, 32'hc121903e} /* (7, 26, 14) {real, imag} */,
  {32'h4031d26e, 32'h409e613e} /* (7, 26, 13) {real, imag} */,
  {32'h410cc8f6, 32'h3fce8944} /* (7, 26, 12) {real, imag} */,
  {32'h41485711, 32'hbf27c870} /* (7, 26, 11) {real, imag} */,
  {32'h3ff53664, 32'h4088025e} /* (7, 26, 10) {real, imag} */,
  {32'h402bded6, 32'h404c408d} /* (7, 26, 9) {real, imag} */,
  {32'h40ad4f60, 32'h411e1e7c} /* (7, 26, 8) {real, imag} */,
  {32'hc1245192, 32'h411334cd} /* (7, 26, 7) {real, imag} */,
  {32'hc0cba20e, 32'hc11d9586} /* (7, 26, 6) {real, imag} */,
  {32'h41301377, 32'hc04f715f} /* (7, 26, 5) {real, imag} */,
  {32'hbfce24dc, 32'h40a4a8b6} /* (7, 26, 4) {real, imag} */,
  {32'h40ddc653, 32'h412bd12a} /* (7, 26, 3) {real, imag} */,
  {32'h404d403a, 32'h40efa426} /* (7, 26, 2) {real, imag} */,
  {32'hc16b2650, 32'h4090401d} /* (7, 26, 1) {real, imag} */,
  {32'hc1463789, 32'hc01ac63d} /* (7, 26, 0) {real, imag} */,
  {32'h41046712, 32'h3fba8dc6} /* (7, 25, 31) {real, imag} */,
  {32'h40e8539c, 32'h40953855} /* (7, 25, 30) {real, imag} */,
  {32'h400a9b59, 32'hc05afbda} /* (7, 25, 29) {real, imag} */,
  {32'h403c0c8c, 32'h409a0563} /* (7, 25, 28) {real, imag} */,
  {32'hc08e4f12, 32'h3ff6ae64} /* (7, 25, 27) {real, imag} */,
  {32'h400597ee, 32'h41230e9b} /* (7, 25, 26) {real, imag} */,
  {32'h3f2dbad0, 32'h402978c8} /* (7, 25, 25) {real, imag} */,
  {32'hc025bff0, 32'h404b00cc} /* (7, 25, 24) {real, imag} */,
  {32'hc08cd54c, 32'h3ff5e4cc} /* (7, 25, 23) {real, imag} */,
  {32'h416423df, 32'hc04236ee} /* (7, 25, 22) {real, imag} */,
  {32'h41aa18bc, 32'hc0fceecb} /* (7, 25, 21) {real, imag} */,
  {32'h3f7367f8, 32'h40b4b5e6} /* (7, 25, 20) {real, imag} */,
  {32'hc18e7ee2, 32'h411fc753} /* (7, 25, 19) {real, imag} */,
  {32'hc11dfea5, 32'h40bf1eaa} /* (7, 25, 18) {real, imag} */,
  {32'hc11f874c, 32'h4115e9c4} /* (7, 25, 17) {real, imag} */,
  {32'h40ba4b1d, 32'h3f650178} /* (7, 25, 16) {real, imag} */,
  {32'h40dc79f4, 32'hc16451c5} /* (7, 25, 15) {real, imag} */,
  {32'h40399e90, 32'hc13b0584} /* (7, 25, 14) {real, imag} */,
  {32'h40e79589, 32'hc0593e1f} /* (7, 25, 13) {real, imag} */,
  {32'hc0964a11, 32'hc1383057} /* (7, 25, 12) {real, imag} */,
  {32'hbf4f1910, 32'h40b1fd4b} /* (7, 25, 11) {real, imag} */,
  {32'h40e85eb0, 32'h3f15dfe8} /* (7, 25, 10) {real, imag} */,
  {32'h40cb958f, 32'hc0bbc6e6} /* (7, 25, 9) {real, imag} */,
  {32'h3faf8d39, 32'hc1027cc4} /* (7, 25, 8) {real, imag} */,
  {32'h405ef310, 32'hc174d85f} /* (7, 25, 7) {real, imag} */,
  {32'h4125f9aa, 32'hc0d3aa94} /* (7, 25, 6) {real, imag} */,
  {32'h40e5a3e3, 32'hc11870fd} /* (7, 25, 5) {real, imag} */,
  {32'h40a152ac, 32'hc0c72dfd} /* (7, 25, 4) {real, imag} */,
  {32'hc02abb51, 32'hc084f1b0} /* (7, 25, 3) {real, imag} */,
  {32'hbf5b333c, 32'hc099ea8f} /* (7, 25, 2) {real, imag} */,
  {32'hc12f9200, 32'h41579a04} /* (7, 25, 1) {real, imag} */,
  {32'hbdb47920, 32'h41269c80} /* (7, 25, 0) {real, imag} */,
  {32'hc064292a, 32'h4172666c} /* (7, 24, 31) {real, imag} */,
  {32'hc0ba2f1e, 32'h411d922a} /* (7, 24, 30) {real, imag} */,
  {32'hc14fb923, 32'hc119d5c9} /* (7, 24, 29) {real, imag} */,
  {32'hc115facf, 32'hc181f396} /* (7, 24, 28) {real, imag} */,
  {32'h41261351, 32'hc11e9ee0} /* (7, 24, 27) {real, imag} */,
  {32'hbfc0ec98, 32'hc0285bb8} /* (7, 24, 26) {real, imag} */,
  {32'hc0d36c8b, 32'hc083de99} /* (7, 24, 25) {real, imag} */,
  {32'h40f6e3b4, 32'h40846871} /* (7, 24, 24) {real, imag} */,
  {32'h4199ff45, 32'hc11595b5} /* (7, 24, 23) {real, imag} */,
  {32'h41196f0a, 32'hc0d136de} /* (7, 24, 22) {real, imag} */,
  {32'h40ab6508, 32'hbfd7b398} /* (7, 24, 21) {real, imag} */,
  {32'h410da5f6, 32'hc133dffc} /* (7, 24, 20) {real, imag} */,
  {32'h4025a81b, 32'hc10bd44f} /* (7, 24, 19) {real, imag} */,
  {32'h407f6cae, 32'hc0be5950} /* (7, 24, 18) {real, imag} */,
  {32'hc0ecda9b, 32'hc05c6cd8} /* (7, 24, 17) {real, imag} */,
  {32'hc154c7e0, 32'hbfdc2e82} /* (7, 24, 16) {real, imag} */,
  {32'h40bd6525, 32'hbff26788} /* (7, 24, 15) {real, imag} */,
  {32'h416fccf6, 32'hbf4bf06a} /* (7, 24, 14) {real, imag} */,
  {32'h40fd8aad, 32'h4110526d} /* (7, 24, 13) {real, imag} */,
  {32'hc104ce28, 32'hbea3eee0} /* (7, 24, 12) {real, imag} */,
  {32'hc0bcebf4, 32'h401e0515} /* (7, 24, 11) {real, imag} */,
  {32'h40b012a2, 32'hc05dffe4} /* (7, 24, 10) {real, imag} */,
  {32'h4064b714, 32'hc130879f} /* (7, 24, 9) {real, imag} */,
  {32'hbfcdb4ac, 32'hc0988e25} /* (7, 24, 8) {real, imag} */,
  {32'hc1539c88, 32'hc0df1541} /* (7, 24, 7) {real, imag} */,
  {32'hc0ee8bc0, 32'h3ecfb98c} /* (7, 24, 6) {real, imag} */,
  {32'h40dbb1fb, 32'h3e801b78} /* (7, 24, 5) {real, imag} */,
  {32'h409ed133, 32'hc0e91274} /* (7, 24, 4) {real, imag} */,
  {32'hc16c0a85, 32'hc02b3790} /* (7, 24, 3) {real, imag} */,
  {32'hc0d695a2, 32'hc0b6abc8} /* (7, 24, 2) {real, imag} */,
  {32'h40a2e5e6, 32'hc13f5af2} /* (7, 24, 1) {real, imag} */,
  {32'h405c0dda, 32'h3f913851} /* (7, 24, 0) {real, imag} */,
  {32'h40b71d4a, 32'hbf8f7122} /* (7, 23, 31) {real, imag} */,
  {32'h40be77a3, 32'h400c81f9} /* (7, 23, 30) {real, imag} */,
  {32'h408693b6, 32'h4127db24} /* (7, 23, 29) {real, imag} */,
  {32'h40b277a4, 32'h3ee8eef4} /* (7, 23, 28) {real, imag} */,
  {32'hc0b4803c, 32'hc019608c} /* (7, 23, 27) {real, imag} */,
  {32'h3f968130, 32'h402eac76} /* (7, 23, 26) {real, imag} */,
  {32'hc062bd70, 32'h405c603b} /* (7, 23, 25) {real, imag} */,
  {32'hc04eaf82, 32'hc09aa962} /* (7, 23, 24) {real, imag} */,
  {32'hc0c8471e, 32'hc14a09cc} /* (7, 23, 23) {real, imag} */,
  {32'hc12db38a, 32'hc0841359} /* (7, 23, 22) {real, imag} */,
  {32'hc10d1ce8, 32'hc05d9167} /* (7, 23, 21) {real, imag} */,
  {32'h4048086e, 32'hc163ae29} /* (7, 23, 20) {real, imag} */,
  {32'h4114ffc4, 32'hc1025256} /* (7, 23, 19) {real, imag} */,
  {32'hbfc8d6ee, 32'hc11a693a} /* (7, 23, 18) {real, imag} */,
  {32'hbfae8b65, 32'hc1125dc6} /* (7, 23, 17) {real, imag} */,
  {32'h4114a798, 32'hc0817a21} /* (7, 23, 16) {real, imag} */,
  {32'h41076261, 32'h409ed420} /* (7, 23, 15) {real, imag} */,
  {32'hc0433728, 32'h403f6ef4} /* (7, 23, 14) {real, imag} */,
  {32'hc0b47447, 32'hc0a586da} /* (7, 23, 13) {real, imag} */,
  {32'hbfc0a3f9, 32'h402a72fd} /* (7, 23, 12) {real, imag} */,
  {32'hc0c2f264, 32'hc098c365} /* (7, 23, 11) {real, imag} */,
  {32'h3f101390, 32'hc16184c2} /* (7, 23, 10) {real, imag} */,
  {32'h41094c4d, 32'h4051cdc8} /* (7, 23, 9) {real, imag} */,
  {32'h3f3d98fc, 32'h411170f4} /* (7, 23, 8) {real, imag} */,
  {32'hc0a0f4a3, 32'h4179f82c} /* (7, 23, 7) {real, imag} */,
  {32'hc0fe3998, 32'h41354882} /* (7, 23, 6) {real, imag} */,
  {32'hc0ad3ac1, 32'h3f68ec52} /* (7, 23, 5) {real, imag} */,
  {32'hc0764fab, 32'h3fa24abc} /* (7, 23, 4) {real, imag} */,
  {32'hbf63ab74, 32'h3d9ec5c0} /* (7, 23, 3) {real, imag} */,
  {32'hbfa7310c, 32'h4102f1e4} /* (7, 23, 2) {real, imag} */,
  {32'h3ead0408, 32'h3c014300} /* (7, 23, 1) {real, imag} */,
  {32'h40626463, 32'h3e2062b8} /* (7, 23, 0) {real, imag} */,
  {32'h3fa29af1, 32'hc04c2052} /* (7, 22, 31) {real, imag} */,
  {32'h40bc5f81, 32'h4042b4fa} /* (7, 22, 30) {real, imag} */,
  {32'h41470329, 32'h3ea48a80} /* (7, 22, 29) {real, imag} */,
  {32'h410c9118, 32'hc0a85baf} /* (7, 22, 28) {real, imag} */,
  {32'h40d60e20, 32'hc1231c1b} /* (7, 22, 27) {real, imag} */,
  {32'h410416db, 32'hc0313060} /* (7, 22, 26) {real, imag} */,
  {32'h40a6dbd0, 32'h3ffc7d70} /* (7, 22, 25) {real, imag} */,
  {32'h40e16dac, 32'h3fe9ff7a} /* (7, 22, 24) {real, imag} */,
  {32'hbfdaad7a, 32'h408e91f5} /* (7, 22, 23) {real, imag} */,
  {32'hbfd37237, 32'h411d6992} /* (7, 22, 22) {real, imag} */,
  {32'hc100b77c, 32'hc058ffe0} /* (7, 22, 21) {real, imag} */,
  {32'hc164b93e, 32'hc0de4efa} /* (7, 22, 20) {real, imag} */,
  {32'hc0a51744, 32'hbfb234b8} /* (7, 22, 19) {real, imag} */,
  {32'hc0bcefd1, 32'h3ead1c98} /* (7, 22, 18) {real, imag} */,
  {32'hc061f013, 32'hc08ac12c} /* (7, 22, 17) {real, imag} */,
  {32'h409dad4a, 32'h409c07a0} /* (7, 22, 16) {real, imag} */,
  {32'h41476555, 32'h3ffac540} /* (7, 22, 15) {real, imag} */,
  {32'h41489ba0, 32'h3f63eb00} /* (7, 22, 14) {real, imag} */,
  {32'hc0da29fe, 32'h408dd52c} /* (7, 22, 13) {real, imag} */,
  {32'hbf9212d4, 32'h3fbb210c} /* (7, 22, 12) {real, imag} */,
  {32'h409c854a, 32'h3d95e780} /* (7, 22, 11) {real, imag} */,
  {32'hc0b90561, 32'hc0ba83a0} /* (7, 22, 10) {real, imag} */,
  {32'hc02a9a6a, 32'hc05f4546} /* (7, 22, 9) {real, imag} */,
  {32'h408ae1fc, 32'h40476bbe} /* (7, 22, 8) {real, imag} */,
  {32'hc0aa8e19, 32'h3eec7310} /* (7, 22, 7) {real, imag} */,
  {32'hc105cd6c, 32'hc08e1818} /* (7, 22, 6) {real, imag} */,
  {32'hc0a7afb6, 32'hc157122c} /* (7, 22, 5) {real, imag} */,
  {32'hc09a2e26, 32'hc162ec3e} /* (7, 22, 4) {real, imag} */,
  {32'hc1141e6c, 32'hc0a693d2} /* (7, 22, 3) {real, imag} */,
  {32'hbffa79c0, 32'h411132e8} /* (7, 22, 2) {real, imag} */,
  {32'h403dd4e6, 32'h4090567c} /* (7, 22, 1) {real, imag} */,
  {32'h3f0e6974, 32'h3fab5b91} /* (7, 22, 0) {real, imag} */,
  {32'hbf8ba2e1, 32'hc0a079fc} /* (7, 21, 31) {real, imag} */,
  {32'hc061d3e0, 32'hc0ff3d70} /* (7, 21, 30) {real, imag} */,
  {32'h40843eb9, 32'h3fe00b34} /* (7, 21, 29) {real, imag} */,
  {32'h40a7ef34, 32'h40073162} /* (7, 21, 28) {real, imag} */,
  {32'h4083e614, 32'hbeb158e0} /* (7, 21, 27) {real, imag} */,
  {32'h40603890, 32'h3fbe1f8c} /* (7, 21, 26) {real, imag} */,
  {32'h3eff34b4, 32'hbf945fec} /* (7, 21, 25) {real, imag} */,
  {32'hbfc30ff8, 32'h400e73eb} /* (7, 21, 24) {real, imag} */,
  {32'h40234a56, 32'h40b91730} /* (7, 21, 23) {real, imag} */,
  {32'hbfa28d54, 32'h40531fb0} /* (7, 21, 22) {real, imag} */,
  {32'h401d5b32, 32'hbffba1d8} /* (7, 21, 21) {real, imag} */,
  {32'hc09f0ec3, 32'h40a23921} /* (7, 21, 20) {real, imag} */,
  {32'hc0f47ede, 32'h4109487f} /* (7, 21, 19) {real, imag} */,
  {32'h403a8680, 32'h3fa40421} /* (7, 21, 18) {real, imag} */,
  {32'h4103a9de, 32'h408c0784} /* (7, 21, 17) {real, imag} */,
  {32'h3f199000, 32'h407b7ec3} /* (7, 21, 16) {real, imag} */,
  {32'h3ee18cd0, 32'h409167d0} /* (7, 21, 15) {real, imag} */,
  {32'h3ef6f550, 32'hbe803b08} /* (7, 21, 14) {real, imag} */,
  {32'hc1125279, 32'hc04307b3} /* (7, 21, 13) {real, imag} */,
  {32'hc13a3408, 32'hc1287e31} /* (7, 21, 12) {real, imag} */,
  {32'hc0ec5d7b, 32'hc0a2ec16} /* (7, 21, 11) {real, imag} */,
  {32'h4113b670, 32'hc0a57880} /* (7, 21, 10) {real, imag} */,
  {32'hbef944e4, 32'h40676897} /* (7, 21, 9) {real, imag} */,
  {32'hc09bb95a, 32'h4033a194} /* (7, 21, 8) {real, imag} */,
  {32'h401fd3e7, 32'hc0079c5c} /* (7, 21, 7) {real, imag} */,
  {32'h3f9e8251, 32'hc02d5f0e} /* (7, 21, 6) {real, imag} */,
  {32'hbf8676b7, 32'hbfe777be} /* (7, 21, 5) {real, imag} */,
  {32'hbec38bf8, 32'hc0977240} /* (7, 21, 4) {real, imag} */,
  {32'hbdd56be0, 32'hc0e6e5a3} /* (7, 21, 3) {real, imag} */,
  {32'hbf07c2de, 32'h404376f4} /* (7, 21, 2) {real, imag} */,
  {32'h404f0b65, 32'h3e8b74a0} /* (7, 21, 1) {real, imag} */,
  {32'h3ec15b70, 32'hc0a90f7b} /* (7, 21, 0) {real, imag} */,
  {32'h3ee888f8, 32'h402ef47f} /* (7, 20, 31) {real, imag} */,
  {32'h4078722d, 32'hc090a04b} /* (7, 20, 30) {real, imag} */,
  {32'hc02920e2, 32'h3f9fcb9c} /* (7, 20, 29) {real, imag} */,
  {32'hbf452b44, 32'h40c9eea5} /* (7, 20, 28) {real, imag} */,
  {32'hc00aaee4, 32'hbf836560} /* (7, 20, 27) {real, imag} */,
  {32'hbf0f8514, 32'hc09ab2cf} /* (7, 20, 26) {real, imag} */,
  {32'h3fceb5cc, 32'hc040e580} /* (7, 20, 25) {real, imag} */,
  {32'hc00f27c1, 32'hc07156d2} /* (7, 20, 24) {real, imag} */,
  {32'hbf0f2216, 32'h3f30ee48} /* (7, 20, 23) {real, imag} */,
  {32'h3e87d310, 32'h3fa2e169} /* (7, 20, 22) {real, imag} */,
  {32'hc048d788, 32'h400a31e0} /* (7, 20, 21) {real, imag} */,
  {32'h3fa1b49a, 32'h412fe7eb} /* (7, 20, 20) {real, imag} */,
  {32'hbe9c4ee8, 32'h411865fe} /* (7, 20, 19) {real, imag} */,
  {32'h3fa8aefe, 32'h4055a498} /* (7, 20, 18) {real, imag} */,
  {32'h40ee9ddc, 32'h3f307ed4} /* (7, 20, 17) {real, imag} */,
  {32'hbf63a854, 32'h4004cce0} /* (7, 20, 16) {real, imag} */,
  {32'hc0b7a987, 32'hc0059964} /* (7, 20, 15) {real, imag} */,
  {32'h40ef9878, 32'h3fb799e2} /* (7, 20, 14) {real, imag} */,
  {32'h410fb072, 32'hc019e562} /* (7, 20, 13) {real, imag} */,
  {32'h408a9df6, 32'h3f833d48} /* (7, 20, 12) {real, imag} */,
  {32'hc0b60d6c, 32'h4029456e} /* (7, 20, 11) {real, imag} */,
  {32'hc02f30e6, 32'h3f680270} /* (7, 20, 10) {real, imag} */,
  {32'h407b9a06, 32'h3f8ab2e8} /* (7, 20, 9) {real, imag} */,
  {32'h4003b57b, 32'hc0c82fdd} /* (7, 20, 8) {real, imag} */,
  {32'hbf4adfe8, 32'hbf3456c0} /* (7, 20, 7) {real, imag} */,
  {32'h3f8d6378, 32'h3fa29832} /* (7, 20, 6) {real, imag} */,
  {32'hc02efc11, 32'h3f76a948} /* (7, 20, 5) {real, imag} */,
  {32'h3f2c1fc2, 32'h40976e0a} /* (7, 20, 4) {real, imag} */,
  {32'h40474c23, 32'h40993414} /* (7, 20, 3) {real, imag} */,
  {32'h403dd7e9, 32'hc075ad52} /* (7, 20, 2) {real, imag} */,
  {32'h40b98b51, 32'hc0b3e1fc} /* (7, 20, 1) {real, imag} */,
  {32'hc00360e6, 32'h402d6d4e} /* (7, 20, 0) {real, imag} */,
  {32'hbec93332, 32'hc01ce69c} /* (7, 19, 31) {real, imag} */,
  {32'h3fae822e, 32'hc0622d52} /* (7, 19, 30) {real, imag} */,
  {32'h40f7b6b3, 32'hc0465f88} /* (7, 19, 29) {real, imag} */,
  {32'h3f08eea0, 32'h3f9bebdc} /* (7, 19, 28) {real, imag} */,
  {32'hc05e71d4, 32'h3fe75d2e} /* (7, 19, 27) {real, imag} */,
  {32'h40165a97, 32'hc08083ce} /* (7, 19, 26) {real, imag} */,
  {32'hbef42810, 32'h3e4c7bb8} /* (7, 19, 25) {real, imag} */,
  {32'h3b5ba400, 32'h40539176} /* (7, 19, 24) {real, imag} */,
  {32'hc09ae92f, 32'h40ab82ee} /* (7, 19, 23) {real, imag} */,
  {32'hc0276ffc, 32'h4091144a} /* (7, 19, 22) {real, imag} */,
  {32'hbfcfa40c, 32'hc0412d1c} /* (7, 19, 21) {real, imag} */,
  {32'h4025acce, 32'hc0899ce1} /* (7, 19, 20) {real, imag} */,
  {32'h409070f4, 32'hbdb06120} /* (7, 19, 19) {real, imag} */,
  {32'h3f91531b, 32'hbfd65905} /* (7, 19, 18) {real, imag} */,
  {32'hbd8ac150, 32'hbffd3130} /* (7, 19, 17) {real, imag} */,
  {32'h40b2634e, 32'hc08a39fc} /* (7, 19, 16) {real, imag} */,
  {32'h406c5337, 32'hbcde8c20} /* (7, 19, 15) {real, imag} */,
  {32'h3fb09298, 32'h3fb25c4d} /* (7, 19, 14) {real, imag} */,
  {32'hc085e5a2, 32'hbf443834} /* (7, 19, 13) {real, imag} */,
  {32'hc0fa659e, 32'h3fbf5420} /* (7, 19, 12) {real, imag} */,
  {32'hbf793328, 32'h4073c4f4} /* (7, 19, 11) {real, imag} */,
  {32'hbf387e04, 32'h40f5fed2} /* (7, 19, 10) {real, imag} */,
  {32'hc0a22376, 32'h41155dd7} /* (7, 19, 9) {real, imag} */,
  {32'hc0af423c, 32'hbfcc1752} /* (7, 19, 8) {real, imag} */,
  {32'hc07fb78c, 32'hbfa0441d} /* (7, 19, 7) {real, imag} */,
  {32'hbfa14e5a, 32'h3f7e309c} /* (7, 19, 6) {real, imag} */,
  {32'h402589d6, 32'hc02cec6f} /* (7, 19, 5) {real, imag} */,
  {32'h3fc10882, 32'hc0c38ce3} /* (7, 19, 4) {real, imag} */,
  {32'h40a74990, 32'hc071734e} /* (7, 19, 3) {real, imag} */,
  {32'h40872815, 32'hc0f6c142} /* (7, 19, 2) {real, imag} */,
  {32'h401f048e, 32'h3f1f8af8} /* (7, 19, 1) {real, imag} */,
  {32'h402e6e9c, 32'h40213c0b} /* (7, 19, 0) {real, imag} */,
  {32'hc0be353c, 32'h3f2ac57c} /* (7, 18, 31) {real, imag} */,
  {32'hc09d3623, 32'h3fc0dbe4} /* (7, 18, 30) {real, imag} */,
  {32'h4013c71e, 32'h3f6f7078} /* (7, 18, 29) {real, imag} */,
  {32'h40541c0c, 32'h4023ba93} /* (7, 18, 28) {real, imag} */,
  {32'h40779f61, 32'hbf40352a} /* (7, 18, 27) {real, imag} */,
  {32'h3fcab9b6, 32'hc063da97} /* (7, 18, 26) {real, imag} */,
  {32'h4025a818, 32'hc083b27c} /* (7, 18, 25) {real, imag} */,
  {32'h3f451da0, 32'hbfc8714e} /* (7, 18, 24) {real, imag} */,
  {32'h3f4747c2, 32'hbea31694} /* (7, 18, 23) {real, imag} */,
  {32'h4037dcae, 32'hbf2abd84} /* (7, 18, 22) {real, imag} */,
  {32'h3f124e14, 32'h40832d41} /* (7, 18, 21) {real, imag} */,
  {32'hc050d1e7, 32'h406da165} /* (7, 18, 20) {real, imag} */,
  {32'hbfb562ab, 32'h408cb614} /* (7, 18, 19) {real, imag} */,
  {32'h4056d26c, 32'h3f93b272} /* (7, 18, 18) {real, imag} */,
  {32'h3db25fa0, 32'hc00bd348} /* (7, 18, 17) {real, imag} */,
  {32'h40003d83, 32'hc0602d71} /* (7, 18, 16) {real, imag} */,
  {32'h4058084e, 32'hc01c2cbe} /* (7, 18, 15) {real, imag} */,
  {32'h3ffe62fd, 32'h3fcb54ee} /* (7, 18, 14) {real, imag} */,
  {32'h404db888, 32'h3e2f8ab8} /* (7, 18, 13) {real, imag} */,
  {32'h40a12077, 32'hbdd51c60} /* (7, 18, 12) {real, imag} */,
  {32'hbd37be50, 32'hc0aec8f2} /* (7, 18, 11) {real, imag} */,
  {32'hbda1c160, 32'hc0e039bf} /* (7, 18, 10) {real, imag} */,
  {32'h40e034a8, 32'hbe0050d0} /* (7, 18, 9) {real, imag} */,
  {32'h40a5ea3b, 32'h40f6c1d8} /* (7, 18, 8) {real, imag} */,
  {32'h3fb2287c, 32'h4072bd46} /* (7, 18, 7) {real, imag} */,
  {32'hc0979e2c, 32'h3f9ea154} /* (7, 18, 6) {real, imag} */,
  {32'hbfcbd31c, 32'h403c79b6} /* (7, 18, 5) {real, imag} */,
  {32'hbc0addc0, 32'h3fff574a} /* (7, 18, 4) {real, imag} */,
  {32'h40d2b1c3, 32'hc0559a33} /* (7, 18, 3) {real, imag} */,
  {32'h403d358c, 32'hc00dabf2} /* (7, 18, 2) {real, imag} */,
  {32'hc06defaf, 32'h40bcdbd2} /* (7, 18, 1) {real, imag} */,
  {32'hc018f1d8, 32'h40c17534} /* (7, 18, 0) {real, imag} */,
  {32'hbf15766a, 32'h3f6f97e2} /* (7, 17, 31) {real, imag} */,
  {32'hbf55b788, 32'h403f5f34} /* (7, 17, 30) {real, imag} */,
  {32'hc0c2584a, 32'hc08d687a} /* (7, 17, 29) {real, imag} */,
  {32'hbf87b533, 32'hc041a69e} /* (7, 17, 28) {real, imag} */,
  {32'h3f9511c1, 32'h3f3e5fcc} /* (7, 17, 27) {real, imag} */,
  {32'hc08818a6, 32'h407ecaca} /* (7, 17, 26) {real, imag} */,
  {32'hbf1abbb3, 32'h4097affe} /* (7, 17, 25) {real, imag} */,
  {32'hbf165198, 32'h3fc98dc4} /* (7, 17, 24) {real, imag} */,
  {32'hbe884c34, 32'h3f81b3a0} /* (7, 17, 23) {real, imag} */,
  {32'hbe9afba8, 32'h3fc0fc70} /* (7, 17, 22) {real, imag} */,
  {32'hbfb49592, 32'h40980d9a} /* (7, 17, 21) {real, imag} */,
  {32'h3f3b5168, 32'h3f900de4} /* (7, 17, 20) {real, imag} */,
  {32'hbdc7b640, 32'hc04ba7f4} /* (7, 17, 19) {real, imag} */,
  {32'h3e903050, 32'hbfe4ec34} /* (7, 17, 18) {real, imag} */,
  {32'hc01b9700, 32'hc0524012} /* (7, 17, 17) {real, imag} */,
  {32'hbef624e0, 32'h3f12836e} /* (7, 17, 16) {real, imag} */,
  {32'hbff6114c, 32'h404ee98c} /* (7, 17, 15) {real, imag} */,
  {32'hc088f659, 32'hbfd22962} /* (7, 17, 14) {real, imag} */,
  {32'hc01f69f2, 32'hbf509000} /* (7, 17, 13) {real, imag} */,
  {32'hc06a624a, 32'hc0142cae} /* (7, 17, 12) {real, imag} */,
  {32'hc0685eca, 32'h402d2157} /* (7, 17, 11) {real, imag} */,
  {32'hc03a425c, 32'h4046d51e} /* (7, 17, 10) {real, imag} */,
  {32'hc08b92fc, 32'hbf139b40} /* (7, 17, 9) {real, imag} */,
  {32'hc05e0e0d, 32'hbff5f910} /* (7, 17, 8) {real, imag} */,
  {32'hc052e7b0, 32'h3ff40ff4} /* (7, 17, 7) {real, imag} */,
  {32'hc0244429, 32'h3fcf645e} /* (7, 17, 6) {real, imag} */,
  {32'hc051b237, 32'h40224d28} /* (7, 17, 5) {real, imag} */,
  {32'h3dace100, 32'h404dd9c4} /* (7, 17, 4) {real, imag} */,
  {32'h3ff9b3bd, 32'h3f291b9e} /* (7, 17, 3) {real, imag} */,
  {32'h3fcb0b68, 32'hc04e1edf} /* (7, 17, 2) {real, imag} */,
  {32'hc0448255, 32'hc0251600} /* (7, 17, 1) {real, imag} */,
  {32'hbfd8803c, 32'h3f0b6400} /* (7, 17, 0) {real, imag} */,
  {32'h403a4cdd, 32'h3fe69b6a} /* (7, 16, 31) {real, imag} */,
  {32'h3f124848, 32'hbebac510} /* (7, 16, 30) {real, imag} */,
  {32'hbfbb0d20, 32'h3fd65e58} /* (7, 16, 29) {real, imag} */,
  {32'hc0636a02, 32'h408491f4} /* (7, 16, 28) {real, imag} */,
  {32'hc01fc1f5, 32'h3fedec80} /* (7, 16, 27) {real, imag} */,
  {32'hbf56ca90, 32'h4032ba32} /* (7, 16, 26) {real, imag} */,
  {32'h3f82930a, 32'h3ea9eee0} /* (7, 16, 25) {real, imag} */,
  {32'h407e9dd6, 32'h40077d16} /* (7, 16, 24) {real, imag} */,
  {32'h40020b0a, 32'h4019f046} /* (7, 16, 23) {real, imag} */,
  {32'hbfbce380, 32'h405a4c62} /* (7, 16, 22) {real, imag} */,
  {32'hbf766578, 32'h4052a1e0} /* (7, 16, 21) {real, imag} */,
  {32'h3ff5ad2e, 32'hbdb18200} /* (7, 16, 20) {real, imag} */,
  {32'hc037aed8, 32'hbfa456a0} /* (7, 16, 19) {real, imag} */,
  {32'hc072d9e0, 32'h3e973ec0} /* (7, 16, 18) {real, imag} */,
  {32'hbdaf3500, 32'h3ff4ae08} /* (7, 16, 17) {real, imag} */,
  {32'hbf8915d4, 32'hbf5daf38} /* (7, 16, 16) {real, imag} */,
  {32'hbf81e5e4, 32'hbdd0ea40} /* (7, 16, 15) {real, imag} */,
  {32'h3e511b90, 32'h3e7b7520} /* (7, 16, 14) {real, imag} */,
  {32'h3f86f958, 32'hbfd10a28} /* (7, 16, 13) {real, imag} */,
  {32'h3f9b1f50, 32'hbdf1a760} /* (7, 16, 12) {real, imag} */,
  {32'h4023c797, 32'hbfe2e1a5} /* (7, 16, 11) {real, imag} */,
  {32'h409a2380, 32'hc111db3c} /* (7, 16, 10) {real, imag} */,
  {32'h407bac3c, 32'hbffc5d6c} /* (7, 16, 9) {real, imag} */,
  {32'h40a6c348, 32'h405122a6} /* (7, 16, 8) {real, imag} */,
  {32'h40a6873c, 32'h40324eda} /* (7, 16, 7) {real, imag} */,
  {32'hbd5af3e0, 32'h3f87f110} /* (7, 16, 6) {real, imag} */,
  {32'hbff33628, 32'hc02fc91a} /* (7, 16, 5) {real, imag} */,
  {32'hbf6cdc5e, 32'hc03b04ae} /* (7, 16, 4) {real, imag} */,
  {32'hbeb48190, 32'hbfbfe29a} /* (7, 16, 3) {real, imag} */,
  {32'hc00794ce, 32'hc085d0b5} /* (7, 16, 2) {real, imag} */,
  {32'hc04723cc, 32'hc02da5cc} /* (7, 16, 1) {real, imag} */,
  {32'hbf98330e, 32'hbfb27950} /* (7, 16, 0) {real, imag} */,
  {32'hbfe0a123, 32'hc0138e60} /* (7, 15, 31) {real, imag} */,
  {32'hc0a2acce, 32'hc0ecc6a6} /* (7, 15, 30) {real, imag} */,
  {32'hc0acfbfc, 32'hc09bb6ea} /* (7, 15, 29) {real, imag} */,
  {32'hc019b692, 32'hc066c8a8} /* (7, 15, 28) {real, imag} */,
  {32'hbf3ecf82, 32'hbfb5e868} /* (7, 15, 27) {real, imag} */,
  {32'h3e8638d8, 32'h3f3dac48} /* (7, 15, 26) {real, imag} */,
  {32'hbeee4f72, 32'h40430d54} /* (7, 15, 25) {real, imag} */,
  {32'hbfb06dec, 32'hbe0a0740} /* (7, 15, 24) {real, imag} */,
  {32'hc0359b66, 32'h3f2d5ea8} /* (7, 15, 23) {real, imag} */,
  {32'hc08b60e0, 32'h40469f00} /* (7, 15, 22) {real, imag} */,
  {32'hc051f5a1, 32'h3eea34c0} /* (7, 15, 21) {real, imag} */,
  {32'hc020ce30, 32'h40153872} /* (7, 15, 20) {real, imag} */,
  {32'hc05f7616, 32'h406b8524} /* (7, 15, 19) {real, imag} */,
  {32'h3d4a0b80, 32'h4081b643} /* (7, 15, 18) {real, imag} */,
  {32'h401cc626, 32'hbe1d8aa8} /* (7, 15, 17) {real, imag} */,
  {32'hc0ffba54, 32'hc02e1414} /* (7, 15, 16) {real, imag} */,
  {32'hc0d35823, 32'hbfe31688} /* (7, 15, 15) {real, imag} */,
  {32'h3fbce9c1, 32'h3fe0f352} /* (7, 15, 14) {real, imag} */,
  {32'hbf96045b, 32'h40564408} /* (7, 15, 13) {real, imag} */,
  {32'hc0a1d035, 32'h3f3ae898} /* (7, 15, 12) {real, imag} */,
  {32'hbfdcaf00, 32'hbff2f8b2} /* (7, 15, 11) {real, imag} */,
  {32'h404da3bc, 32'hbff5ab9c} /* (7, 15, 10) {real, imag} */,
  {32'h408539ac, 32'h3f013060} /* (7, 15, 9) {real, imag} */,
  {32'hbf1dfe34, 32'h3f05eb20} /* (7, 15, 8) {real, imag} */,
  {32'hc0968822, 32'hbf8778b4} /* (7, 15, 7) {real, imag} */,
  {32'hc074e603, 32'h3ed4b698} /* (7, 15, 6) {real, imag} */,
  {32'h3f5f33ac, 32'h3ea2e504} /* (7, 15, 5) {real, imag} */,
  {32'h403250f0, 32'hbfb8af20} /* (7, 15, 4) {real, imag} */,
  {32'h3e91eb4c, 32'hc027669c} /* (7, 15, 3) {real, imag} */,
  {32'hbf1d3460, 32'hbfd5f42a} /* (7, 15, 2) {real, imag} */,
  {32'h3ea6beb8, 32'hc04ea0a0} /* (7, 15, 1) {real, imag} */,
  {32'h3fc7b436, 32'hbf0019a0} /* (7, 15, 0) {real, imag} */,
  {32'hbeec9218, 32'hbf5f6444} /* (7, 14, 31) {real, imag} */,
  {32'h3e91b4d0, 32'h4063a89a} /* (7, 14, 30) {real, imag} */,
  {32'hbf290d42, 32'h40c2cb63} /* (7, 14, 29) {real, imag} */,
  {32'hc04d4c16, 32'h405b9c5b} /* (7, 14, 28) {real, imag} */,
  {32'hc0271ced, 32'h40332d7e} /* (7, 14, 27) {real, imag} */,
  {32'hbfafd9fa, 32'hc0acf25e} /* (7, 14, 26) {real, imag} */,
  {32'hc051902c, 32'hc07d1551} /* (7, 14, 25) {real, imag} */,
  {32'h3fd51130, 32'h3fcb561a} /* (7, 14, 24) {real, imag} */,
  {32'h4081aee3, 32'h4045a1bc} /* (7, 14, 23) {real, imag} */,
  {32'h4080dff7, 32'h3f5b34cc} /* (7, 14, 22) {real, imag} */,
  {32'h3ef2c318, 32'hbeb951d0} /* (7, 14, 21) {real, imag} */,
  {32'hc06ba0fb, 32'hbf8e0636} /* (7, 14, 20) {real, imag} */,
  {32'h3fc6bbdf, 32'hc0092f90} /* (7, 14, 19) {real, imag} */,
  {32'h4081e288, 32'h4000b967} /* (7, 14, 18) {real, imag} */,
  {32'hbf476e6c, 32'h409417ea} /* (7, 14, 17) {real, imag} */,
  {32'hc02b3e9b, 32'h401b7393} /* (7, 14, 16) {real, imag} */,
  {32'hc0580f8e, 32'hc0023562} /* (7, 14, 15) {real, imag} */,
  {32'h3e9863d4, 32'hc047a6b7} /* (7, 14, 14) {real, imag} */,
  {32'h40cd7f04, 32'hc0464c86} /* (7, 14, 13) {real, imag} */,
  {32'h4090f1f1, 32'h40610a9b} /* (7, 14, 12) {real, imag} */,
  {32'h3f4c1a25, 32'h40621144} /* (7, 14, 11) {real, imag} */,
  {32'hbf218794, 32'hc0049f56} /* (7, 14, 10) {real, imag} */,
  {32'hbfc663c0, 32'hc08a1c28} /* (7, 14, 9) {real, imag} */,
  {32'hc093329d, 32'hc0603650} /* (7, 14, 8) {real, imag} */,
  {32'hc043278e, 32'hbfcbcf80} /* (7, 14, 7) {real, imag} */,
  {32'hbeb84cf0, 32'hbff8ef14} /* (7, 14, 6) {real, imag} */,
  {32'h3fe060cc, 32'hc084dc4b} /* (7, 14, 5) {real, imag} */,
  {32'hbfd5890a, 32'hbfdd293a} /* (7, 14, 4) {real, imag} */,
  {32'hc0e64e55, 32'hbf295814} /* (7, 14, 3) {real, imag} */,
  {32'hc0a66366, 32'h4067ec7e} /* (7, 14, 2) {real, imag} */,
  {32'hbff51bba, 32'h403e2c1c} /* (7, 14, 1) {real, imag} */,
  {32'h3ff9942f, 32'hbf30345c} /* (7, 14, 0) {real, imag} */,
  {32'hbea16932, 32'hc08a7400} /* (7, 13, 31) {real, imag} */,
  {32'h3fcf4a1e, 32'hc00df432} /* (7, 13, 30) {real, imag} */,
  {32'h404bef7a, 32'hc04e99e8} /* (7, 13, 29) {real, imag} */,
  {32'h40866e14, 32'hc018e9be} /* (7, 13, 28) {real, imag} */,
  {32'hbfd32348, 32'hc06751bd} /* (7, 13, 27) {real, imag} */,
  {32'hbfae9f9a, 32'hc01b000d} /* (7, 13, 26) {real, imag} */,
  {32'hc04c1a9a, 32'hbf92c641} /* (7, 13, 25) {real, imag} */,
  {32'hc0958718, 32'h3f0ad3d8} /* (7, 13, 24) {real, imag} */,
  {32'hc095b6bd, 32'hc01495b6} /* (7, 13, 23) {real, imag} */,
  {32'hc0a9b06c, 32'hc0a003ba} /* (7, 13, 22) {real, imag} */,
  {32'hc04d3c62, 32'hc10864a2} /* (7, 13, 21) {real, imag} */,
  {32'hbcc0c4c0, 32'hc10aafda} /* (7, 13, 20) {real, imag} */,
  {32'h3ea33508, 32'h3fe53e6e} /* (7, 13, 19) {real, imag} */,
  {32'hc01c9084, 32'h402e82c8} /* (7, 13, 18) {real, imag} */,
  {32'h3fcfda6d, 32'hc024794a} /* (7, 13, 17) {real, imag} */,
  {32'hc01e053b, 32'hbfa850ee} /* (7, 13, 16) {real, imag} */,
  {32'hc0b13ee6, 32'hbf0d1641} /* (7, 13, 15) {real, imag} */,
  {32'h3f2810e0, 32'h401e419e} /* (7, 13, 14) {real, imag} */,
  {32'hbd54f640, 32'h409afd84} /* (7, 13, 13) {real, imag} */,
  {32'h4071072b, 32'hc02a2ce4} /* (7, 13, 12) {real, imag} */,
  {32'hc0b7eb99, 32'hbe976540} /* (7, 13, 11) {real, imag} */,
  {32'hc0eb8908, 32'hc05cea2c} /* (7, 13, 10) {real, imag} */,
  {32'hc104216b, 32'hc03824c8} /* (7, 13, 9) {real, imag} */,
  {32'h3fee2bac, 32'h3f5e8a7c} /* (7, 13, 8) {real, imag} */,
  {32'h4073dc8a, 32'h3f87e27d} /* (7, 13, 7) {real, imag} */,
  {32'h40a79574, 32'hbf95ba9a} /* (7, 13, 6) {real, imag} */,
  {32'hbeac134c, 32'hc09984f8} /* (7, 13, 5) {real, imag} */,
  {32'hc00ea6c2, 32'h4091ad3f} /* (7, 13, 4) {real, imag} */,
  {32'h4014b191, 32'h40cfca0b} /* (7, 13, 3) {real, imag} */,
  {32'hbe88b594, 32'hbeb45920} /* (7, 13, 2) {real, imag} */,
  {32'hbf9ba953, 32'hc047e104} /* (7, 13, 1) {real, imag} */,
  {32'h3f575470, 32'hbfbda01a} /* (7, 13, 0) {real, imag} */,
  {32'hbf42be04, 32'hc00d5aff} /* (7, 12, 31) {real, imag} */,
  {32'h3fad309e, 32'hc0942f33} /* (7, 12, 30) {real, imag} */,
  {32'h408b3f2f, 32'h40d60b17} /* (7, 12, 29) {real, imag} */,
  {32'hc0759f4b, 32'hbfd464c4} /* (7, 12, 28) {real, imag} */,
  {32'hc01d6088, 32'hc0850f58} /* (7, 12, 27) {real, imag} */,
  {32'h403b4f97, 32'h4084b7a9} /* (7, 12, 26) {real, imag} */,
  {32'h411b8656, 32'h3f7a4db8} /* (7, 12, 25) {real, imag} */,
  {32'h40a0e664, 32'hc0015d2e} /* (7, 12, 24) {real, imag} */,
  {32'hc0857732, 32'hc0615f92} /* (7, 12, 23) {real, imag} */,
  {32'h3fa61764, 32'h4027e490} /* (7, 12, 22) {real, imag} */,
  {32'h411b16fe, 32'h408c88de} /* (7, 12, 21) {real, imag} */,
  {32'h4028f0f9, 32'h4093d162} /* (7, 12, 20) {real, imag} */,
  {32'hc0ce9220, 32'h3f611d28} /* (7, 12, 19) {real, imag} */,
  {32'hbf661f1c, 32'hbe4f8bf8} /* (7, 12, 18) {real, imag} */,
  {32'hbf0db1a0, 32'hc0e570ce} /* (7, 12, 17) {real, imag} */,
  {32'hc0a36c84, 32'hc1230889} /* (7, 12, 16) {real, imag} */,
  {32'h3ffdda79, 32'hc07a1a94} /* (7, 12, 15) {real, imag} */,
  {32'h4045cc39, 32'h407c5677} /* (7, 12, 14) {real, imag} */,
  {32'h400868da, 32'h4099f171} /* (7, 12, 13) {real, imag} */,
  {32'hbeb15d70, 32'h405b8ee0} /* (7, 12, 12) {real, imag} */,
  {32'hc0987fd8, 32'hbe99f6d0} /* (7, 12, 11) {real, imag} */,
  {32'hbe9ddf8c, 32'hc0c0daa4} /* (7, 12, 10) {real, imag} */,
  {32'hc061ff2a, 32'h3f335c60} /* (7, 12, 9) {real, imag} */,
  {32'hc0aaa36c, 32'h400ab79a} /* (7, 12, 8) {real, imag} */,
  {32'hbf5633e8, 32'hbe7b7c40} /* (7, 12, 7) {real, imag} */,
  {32'hbe449480, 32'hbe5785bc} /* (7, 12, 6) {real, imag} */,
  {32'h3ea677f8, 32'hc0a9e6c5} /* (7, 12, 5) {real, imag} */,
  {32'h3dca7770, 32'hc0b0a252} /* (7, 12, 4) {real, imag} */,
  {32'hbf6ec74c, 32'h406c12e0} /* (7, 12, 3) {real, imag} */,
  {32'hc092616a, 32'h403fd376} /* (7, 12, 2) {real, imag} */,
  {32'hc073e3e6, 32'hbf30f834} /* (7, 12, 1) {real, imag} */,
  {32'hbe3be118, 32'hc08d9371} /* (7, 12, 0) {real, imag} */,
  {32'hc054188a, 32'h3f97025a} /* (7, 11, 31) {real, imag} */,
  {32'hc08f6b90, 32'hbfc18730} /* (7, 11, 30) {real, imag} */,
  {32'hc1647278, 32'hc1220e3c} /* (7, 11, 29) {real, imag} */,
  {32'hbea1e7e0, 32'hc0ff8c85} /* (7, 11, 28) {real, imag} */,
  {32'h41197bd4, 32'hc118c3e6} /* (7, 11, 27) {real, imag} */,
  {32'hc01ac7e0, 32'hbf6d2ce8} /* (7, 11, 26) {real, imag} */,
  {32'hc0757812, 32'h40b7f7a1} /* (7, 11, 25) {real, imag} */,
  {32'hc0ae23a2, 32'h40b5241c} /* (7, 11, 24) {real, imag} */,
  {32'hc0821dc5, 32'h40b5e458} /* (7, 11, 23) {real, imag} */,
  {32'hc10013fa, 32'h406f3fa0} /* (7, 11, 22) {real, imag} */,
  {32'hc093eeb7, 32'h41023898} /* (7, 11, 21) {real, imag} */,
  {32'h40a8c443, 32'h40934c8d} /* (7, 11, 20) {real, imag} */,
  {32'h406f87c1, 32'h40c16fee} /* (7, 11, 19) {real, imag} */,
  {32'h407dd8c2, 32'hbf546262} /* (7, 11, 18) {real, imag} */,
  {32'hbe2c9aa0, 32'hc0474008} /* (7, 11, 17) {real, imag} */,
  {32'h3ff2367c, 32'hc0952d9a} /* (7, 11, 16) {real, imag} */,
  {32'h4060446e, 32'hc091f958} /* (7, 11, 15) {real, imag} */,
  {32'h4141a75c, 32'hc0b4e120} /* (7, 11, 14) {real, imag} */,
  {32'h412c961f, 32'hbffe328e} /* (7, 11, 13) {real, imag} */,
  {32'hbfd4d00c, 32'hbfa9fdf0} /* (7, 11, 12) {real, imag} */,
  {32'hc0c719cd, 32'h3f3c49fc} /* (7, 11, 11) {real, imag} */,
  {32'hbd9dcf00, 32'h3f1c2f0c} /* (7, 11, 10) {real, imag} */,
  {32'h40855640, 32'hbfddd96a} /* (7, 11, 9) {real, imag} */,
  {32'h40b4406e, 32'hc06f44e0} /* (7, 11, 8) {real, imag} */,
  {32'hc05ac5d7, 32'hc0a88544} /* (7, 11, 7) {real, imag} */,
  {32'h3cbc37c0, 32'h40b9d6cd} /* (7, 11, 6) {real, imag} */,
  {32'hc0234260, 32'h40d76e72} /* (7, 11, 5) {real, imag} */,
  {32'hbf440474, 32'hc0a9ae98} /* (7, 11, 4) {real, imag} */,
  {32'h3fb28e72, 32'hc0228ce2} /* (7, 11, 3) {real, imag} */,
  {32'hc07b3b92, 32'hbf02a80e} /* (7, 11, 2) {real, imag} */,
  {32'hc0dd1e3a, 32'hc04fbc90} /* (7, 11, 1) {real, imag} */,
  {32'hc0991dee, 32'hc0ad8499} /* (7, 11, 0) {real, imag} */,
  {32'hbf32cc46, 32'h3ed58dc8} /* (7, 10, 31) {real, imag} */,
  {32'hbfbabd24, 32'hc002b836} /* (7, 10, 30) {real, imag} */,
  {32'h4035f85c, 32'hc15c5ae6} /* (7, 10, 29) {real, imag} */,
  {32'h411aea14, 32'hc10b7352} /* (7, 10, 28) {real, imag} */,
  {32'h4127916c, 32'h40928a6a} /* (7, 10, 27) {real, imag} */,
  {32'h4098b6c6, 32'hbf8fa293} /* (7, 10, 26) {real, imag} */,
  {32'h3fc0d82c, 32'h402b4c68} /* (7, 10, 25) {real, imag} */,
  {32'hbecb53a8, 32'h3f23733c} /* (7, 10, 24) {real, imag} */,
  {32'h401ef1ab, 32'hc04f74b0} /* (7, 10, 23) {real, imag} */,
  {32'h3f13c3ba, 32'hbec15340} /* (7, 10, 22) {real, imag} */,
  {32'hc00bc65a, 32'h4073bedc} /* (7, 10, 21) {real, imag} */,
  {32'hc104281a, 32'h41255d07} /* (7, 10, 20) {real, imag} */,
  {32'hc04d4f9c, 32'h40559bf8} /* (7, 10, 19) {real, imag} */,
  {32'hc0b3a77f, 32'h3d8a84e0} /* (7, 10, 18) {real, imag} */,
  {32'hc036ef55, 32'h4008504b} /* (7, 10, 17) {real, imag} */,
  {32'h4011f4b9, 32'h40840158} /* (7, 10, 16) {real, imag} */,
  {32'hc0570bdc, 32'h407c886c} /* (7, 10, 15) {real, imag} */,
  {32'h410c5b6e, 32'hc0d684b4} /* (7, 10, 14) {real, imag} */,
  {32'h4181ce2e, 32'hc0af7ad2} /* (7, 10, 13) {real, imag} */,
  {32'h411c6366, 32'h41038120} /* (7, 10, 12) {real, imag} */,
  {32'h3f85ce1a, 32'h4096489a} /* (7, 10, 11) {real, imag} */,
  {32'h3f7f3358, 32'hc0956ad8} /* (7, 10, 10) {real, imag} */,
  {32'hc006ddd2, 32'hc0503338} /* (7, 10, 9) {real, imag} */,
  {32'hc0e54352, 32'hbf40c558} /* (7, 10, 8) {real, imag} */,
  {32'hc0d51af9, 32'hc090b833} /* (7, 10, 7) {real, imag} */,
  {32'hc004973c, 32'h40d04c70} /* (7, 10, 6) {real, imag} */,
  {32'hc003ab63, 32'h40dba40c} /* (7, 10, 5) {real, imag} */,
  {32'h40fdd8b8, 32'h3fd30234} /* (7, 10, 4) {real, imag} */,
  {32'h40add4e9, 32'h3fd53bd0} /* (7, 10, 3) {real, imag} */,
  {32'hbf389dd0, 32'hc0913f38} /* (7, 10, 2) {real, imag} */,
  {32'h3f90925c, 32'h3f159224} /* (7, 10, 1) {real, imag} */,
  {32'hc0280eb3, 32'hbee59335} /* (7, 10, 0) {real, imag} */,
  {32'h40c99a76, 32'h40a5199e} /* (7, 9, 31) {real, imag} */,
  {32'h40b8452b, 32'h402f840f} /* (7, 9, 30) {real, imag} */,
  {32'h40ad903c, 32'hbf971ae4} /* (7, 9, 29) {real, imag} */,
  {32'h401117c3, 32'hc03fce66} /* (7, 9, 28) {real, imag} */,
  {32'hbc18d700, 32'hc0282df0} /* (7, 9, 27) {real, imag} */,
  {32'hc0bc4e40, 32'hc04ef2ce} /* (7, 9, 26) {real, imag} */,
  {32'hc0750d4c, 32'hc0e6ccde} /* (7, 9, 25) {real, imag} */,
  {32'hc0654d62, 32'hbf7b274c} /* (7, 9, 24) {real, imag} */,
  {32'h3e8e14b0, 32'h413d535e} /* (7, 9, 23) {real, imag} */,
  {32'h4105a526, 32'h415507d0} /* (7, 9, 22) {real, imag} */,
  {32'hc144fbde, 32'h403f0743} /* (7, 9, 21) {real, imag} */,
  {32'hc10f13f0, 32'hbe9dd9a0} /* (7, 9, 20) {real, imag} */,
  {32'h406198d0, 32'h40a149d2} /* (7, 9, 19) {real, imag} */,
  {32'h40c0b9b6, 32'h401ccf6f} /* (7, 9, 18) {real, imag} */,
  {32'h3fedd585, 32'h40915a5b} /* (7, 9, 17) {real, imag} */,
  {32'h40e01b1f, 32'h403400b6} /* (7, 9, 16) {real, imag} */,
  {32'h3f1ba574, 32'hc073d7b8} /* (7, 9, 15) {real, imag} */,
  {32'hc0b3d790, 32'h402ee26e} /* (7, 9, 14) {real, imag} */,
  {32'h409f0673, 32'h415c6d97} /* (7, 9, 13) {real, imag} */,
  {32'h3f45daf6, 32'hbff3a106} /* (7, 9, 12) {real, imag} */,
  {32'hc122feb4, 32'hc13ed80a} /* (7, 9, 11) {real, imag} */,
  {32'hc14a8a9b, 32'hc06d0d4e} /* (7, 9, 10) {real, imag} */,
  {32'hc129931f, 32'h4147346c} /* (7, 9, 9) {real, imag} */,
  {32'hc0e04636, 32'h40814e95} /* (7, 9, 8) {real, imag} */,
  {32'h3f9ee368, 32'hbfbe3230} /* (7, 9, 7) {real, imag} */,
  {32'hc131641e, 32'h4023e6c0} /* (7, 9, 6) {real, imag} */,
  {32'hc0fff517, 32'h40100bf2} /* (7, 9, 5) {real, imag} */,
  {32'h407481b7, 32'h40eeeae1} /* (7, 9, 4) {real, imag} */,
  {32'h4088c4ea, 32'h412699b8} /* (7, 9, 3) {real, imag} */,
  {32'h3fd2c4ce, 32'h3f0b0814} /* (7, 9, 2) {real, imag} */,
  {32'h3fb93afa, 32'h3fc33046} /* (7, 9, 1) {real, imag} */,
  {32'h410a584f, 32'h407fecdc} /* (7, 9, 0) {real, imag} */,
  {32'h408569ee, 32'hc06f3ec2} /* (7, 8, 31) {real, imag} */,
  {32'hc1014571, 32'h409a7319} /* (7, 8, 30) {real, imag} */,
  {32'hc138aa45, 32'h412083c3} /* (7, 8, 29) {real, imag} */,
  {32'hc1303963, 32'hc0a1acc8} /* (7, 8, 28) {real, imag} */,
  {32'hc0a7506a, 32'hc01010f0} /* (7, 8, 27) {real, imag} */,
  {32'hbf7a3f40, 32'h40af3386} /* (7, 8, 26) {real, imag} */,
  {32'hc027c562, 32'h411af752} /* (7, 8, 25) {real, imag} */,
  {32'hbffbb900, 32'h418b6eec} /* (7, 8, 24) {real, imag} */,
  {32'hbf842650, 32'h408a4cd6} /* (7, 8, 23) {real, imag} */,
  {32'h3fdb86e4, 32'hc0e5c6da} /* (7, 8, 22) {real, imag} */,
  {32'h4098e9c6, 32'hbe725f40} /* (7, 8, 21) {real, imag} */,
  {32'h414c51c2, 32'h404a5dc2} /* (7, 8, 20) {real, imag} */,
  {32'hc0a195d6, 32'h414bbc45} /* (7, 8, 19) {real, imag} */,
  {32'h3fd3596c, 32'h41a7df2e} /* (7, 8, 18) {real, imag} */,
  {32'h3f9bd68c, 32'h402d9970} /* (7, 8, 17) {real, imag} */,
  {32'hc0644fa2, 32'hbf9d4212} /* (7, 8, 16) {real, imag} */,
  {32'h3ff07c7c, 32'h40d5712a} /* (7, 8, 15) {real, imag} */,
  {32'h3fca0514, 32'hc0072cf8} /* (7, 8, 14) {real, imag} */,
  {32'hbf6b4998, 32'hc0dcb3e2} /* (7, 8, 13) {real, imag} */,
  {32'hc007b4f2, 32'h3faf5b4c} /* (7, 8, 12) {real, imag} */,
  {32'h3f58e174, 32'h4097b8f2} /* (7, 8, 11) {real, imag} */,
  {32'h41368e45, 32'h4040e644} /* (7, 8, 10) {real, imag} */,
  {32'h41895038, 32'h40a5b75a} /* (7, 8, 9) {real, imag} */,
  {32'h408b5ff9, 32'h40e211bd} /* (7, 8, 8) {real, imag} */,
  {32'h3e66ec20, 32'h413df0a8} /* (7, 8, 7) {real, imag} */,
  {32'h4007dd98, 32'hbfdd69b3} /* (7, 8, 6) {real, imag} */,
  {32'h4006c7f2, 32'h40673693} /* (7, 8, 5) {real, imag} */,
  {32'hbeff49b0, 32'hbf9f5fd6} /* (7, 8, 4) {real, imag} */,
  {32'h409c062a, 32'hc163ea0c} /* (7, 8, 3) {real, imag} */,
  {32'hbf008b00, 32'hc06b00d0} /* (7, 8, 2) {real, imag} */,
  {32'h3bf44e00, 32'h417f2f36} /* (7, 8, 1) {real, imag} */,
  {32'h40301758, 32'h4044c998} /* (7, 8, 0) {real, imag} */,
  {32'hbfbd0a54, 32'h40f8f8ca} /* (7, 7, 31) {real, imag} */,
  {32'h4064b7fd, 32'h4048ce4f} /* (7, 7, 30) {real, imag} */,
  {32'hbf38e764, 32'h3f9c4dbb} /* (7, 7, 29) {real, imag} */,
  {32'hc0f02b1a, 32'h3f02a108} /* (7, 7, 28) {real, imag} */,
  {32'hc0da25be, 32'hc0f15485} /* (7, 7, 27) {real, imag} */,
  {32'h402a4872, 32'hc0ca856a} /* (7, 7, 26) {real, imag} */,
  {32'hbfc23a42, 32'hc14085f4} /* (7, 7, 25) {real, imag} */,
  {32'hc0719310, 32'hc1641df9} /* (7, 7, 24) {real, imag} */,
  {32'hbf95c8b4, 32'hc0f161d9} /* (7, 7, 23) {real, imag} */,
  {32'hc0a00c1a, 32'hc10c6f94} /* (7, 7, 22) {real, imag} */,
  {32'hc0ce2aee, 32'h40eec9f9} /* (7, 7, 21) {real, imag} */,
  {32'hc12c78ca, 32'h410f31cf} /* (7, 7, 20) {real, imag} */,
  {32'h401e6344, 32'hbd9f6700} /* (7, 7, 19) {real, imag} */,
  {32'h40002fc1, 32'h40dbfa32} /* (7, 7, 18) {real, imag} */,
  {32'hc0421be2, 32'h400716fe} /* (7, 7, 17) {real, imag} */,
  {32'hc07ccfde, 32'hbfad1e76} /* (7, 7, 16) {real, imag} */,
  {32'hbf936de0, 32'h3f42be70} /* (7, 7, 15) {real, imag} */,
  {32'hc0c0ad34, 32'hbfc2c7a0} /* (7, 7, 14) {real, imag} */,
  {32'hbfbfdb24, 32'h3f88ccf2} /* (7, 7, 13) {real, imag} */,
  {32'h400710c4, 32'h404aa9f4} /* (7, 7, 12) {real, imag} */,
  {32'hc129dabd, 32'h40432e6e} /* (7, 7, 11) {real, imag} */,
  {32'hc0a94208, 32'hbfdff984} /* (7, 7, 10) {real, imag} */,
  {32'hbfe1730c, 32'hbfda0c5a} /* (7, 7, 9) {real, imag} */,
  {32'hc012bd9a, 32'hbf6134a0} /* (7, 7, 8) {real, imag} */,
  {32'hc14b09f6, 32'h3f5460b0} /* (7, 7, 7) {real, imag} */,
  {32'hc0f25b28, 32'h40e1cc64} /* (7, 7, 6) {real, imag} */,
  {32'h405b5cc2, 32'hc010f8d4} /* (7, 7, 5) {real, imag} */,
  {32'h41184579, 32'hc1a16979} /* (7, 7, 4) {real, imag} */,
  {32'h410252bf, 32'hc13517fd} /* (7, 7, 3) {real, imag} */,
  {32'h3ffb722c, 32'h4075399a} /* (7, 7, 2) {real, imag} */,
  {32'h3ee30930, 32'h40095c5a} /* (7, 7, 1) {real, imag} */,
  {32'h40b4bc54, 32'h40b4459b} /* (7, 7, 0) {real, imag} */,
  {32'hc0a2eace, 32'h3efe9ab8} /* (7, 6, 31) {real, imag} */,
  {32'hc06e80fa, 32'h3f41f4dc} /* (7, 6, 30) {real, imag} */,
  {32'h408b1c40, 32'hc034e1e3} /* (7, 6, 29) {real, imag} */,
  {32'hc0065511, 32'hc0a9734e} /* (7, 6, 28) {real, imag} */,
  {32'hbe8d48b8, 32'hc0259885} /* (7, 6, 27) {real, imag} */,
  {32'h402c055a, 32'h40adf102} /* (7, 6, 26) {real, imag} */,
  {32'hc0ad02f8, 32'hc0b93150} /* (7, 6, 25) {real, imag} */,
  {32'h409c1ca8, 32'hc0c1a230} /* (7, 6, 24) {real, imag} */,
  {32'h40dcfe69, 32'h3fecd0c6} /* (7, 6, 23) {real, imag} */,
  {32'h410a0400, 32'hc147216b} /* (7, 6, 22) {real, imag} */,
  {32'h404f2968, 32'hc11b07b3} /* (7, 6, 21) {real, imag} */,
  {32'hc0b35c91, 32'h3f9c984e} /* (7, 6, 20) {real, imag} */,
  {32'hbf28a430, 32'hc14fec91} /* (7, 6, 19) {real, imag} */,
  {32'h40808082, 32'hc15e61e0} /* (7, 6, 18) {real, imag} */,
  {32'h3e949a4c, 32'h40901bbe} /* (7, 6, 17) {real, imag} */,
  {32'hc0a65312, 32'hc0a0f1e4} /* (7, 6, 16) {real, imag} */,
  {32'h40c1809d, 32'hc08b32a4} /* (7, 6, 15) {real, imag} */,
  {32'h4135e316, 32'hc069573e} /* (7, 6, 14) {real, imag} */,
  {32'hc15299ea, 32'h40b74502} /* (7, 6, 13) {real, imag} */,
  {32'hc171c5da, 32'h4167fde6} /* (7, 6, 12) {real, imag} */,
  {32'hc0cebdd6, 32'h412ff319} /* (7, 6, 11) {real, imag} */,
  {32'hc0e03d5f, 32'h4087a1e2} /* (7, 6, 10) {real, imag} */,
  {32'hc0362c4a, 32'h411dfd29} /* (7, 6, 9) {real, imag} */,
  {32'hc0bc425e, 32'h41608f56} /* (7, 6, 8) {real, imag} */,
  {32'hc07e75e6, 32'h4108df83} /* (7, 6, 7) {real, imag} */,
  {32'hc130a59b, 32'hbfc2e6d0} /* (7, 6, 6) {real, imag} */,
  {32'hc0d227a2, 32'hc10cbe4a} /* (7, 6, 5) {real, imag} */,
  {32'h408d3ceb, 32'hc0ef6378} /* (7, 6, 4) {real, imag} */,
  {32'h40dffeb7, 32'h3e11c1e0} /* (7, 6, 3) {real, imag} */,
  {32'h41714752, 32'hc0615cdc} /* (7, 6, 2) {real, imag} */,
  {32'h4121d2a2, 32'hc018dbc0} /* (7, 6, 1) {real, imag} */,
  {32'h4026f2f4, 32'h40573253} /* (7, 6, 0) {real, imag} */,
  {32'hc00a3530, 32'h40951402} /* (7, 5, 31) {real, imag} */,
  {32'hc0675e6f, 32'h40826373} /* (7, 5, 30) {real, imag} */,
  {32'hc1257282, 32'h405671f4} /* (7, 5, 29) {real, imag} */,
  {32'h4088c826, 32'h412a6f23} /* (7, 5, 28) {real, imag} */,
  {32'hc18dd7c8, 32'hc10a9953} /* (7, 5, 27) {real, imag} */,
  {32'hc18249ef, 32'hc181230e} /* (7, 5, 26) {real, imag} */,
  {32'h4121cba0, 32'h3fb197dc} /* (7, 5, 25) {real, imag} */,
  {32'h41a46093, 32'hc151b025} /* (7, 5, 24) {real, imag} */,
  {32'h415d23f0, 32'hc1629ff0} /* (7, 5, 23) {real, imag} */,
  {32'hc01b9170, 32'hc0f8c9e6} /* (7, 5, 22) {real, imag} */,
  {32'hc1076c1c, 32'hc180d90b} /* (7, 5, 21) {real, imag} */,
  {32'hc0895aa9, 32'hc1453ab3} /* (7, 5, 20) {real, imag} */,
  {32'h41506b64, 32'hc0c3f9e0} /* (7, 5, 19) {real, imag} */,
  {32'h41301176, 32'h41426e60} /* (7, 5, 18) {real, imag} */,
  {32'hc19c26ab, 32'h410fb753} /* (7, 5, 17) {real, imag} */,
  {32'hc115d585, 32'h40ee5c74} /* (7, 5, 16) {real, imag} */,
  {32'h40920845, 32'hc032405c} /* (7, 5, 15) {real, imag} */,
  {32'h4132c8a4, 32'hc0eb1044} /* (7, 5, 14) {real, imag} */,
  {32'h40161e49, 32'h3ec3c1e0} /* (7, 5, 13) {real, imag} */,
  {32'hc009061a, 32'hc14e605e} /* (7, 5, 12) {real, imag} */,
  {32'h3ec12e30, 32'hc0dc060e} /* (7, 5, 11) {real, imag} */,
  {32'hc03bfe24, 32'hc091032a} /* (7, 5, 10) {real, imag} */,
  {32'h40095e04, 32'hc187c2aa} /* (7, 5, 9) {real, imag} */,
  {32'hc03c5e04, 32'hc1db68ce} /* (7, 5, 8) {real, imag} */,
  {32'h411b801a, 32'hc16103fe} /* (7, 5, 7) {real, imag} */,
  {32'h416ef115, 32'hc10165a8} /* (7, 5, 6) {real, imag} */,
  {32'h410ecd78, 32'hc1754400} /* (7, 5, 5) {real, imag} */,
  {32'h40b63274, 32'hbfd21ab6} /* (7, 5, 4) {real, imag} */,
  {32'hbf3593d0, 32'hc00a6ce0} /* (7, 5, 3) {real, imag} */,
  {32'hbf79bb08, 32'hc18cd436} /* (7, 5, 2) {real, imag} */,
  {32'hbe3fbcc0, 32'hc08fed19} /* (7, 5, 1) {real, imag} */,
  {32'h40b23916, 32'h410607fd} /* (7, 5, 0) {real, imag} */,
  {32'h40cdaf06, 32'hc0d48fbc} /* (7, 4, 31) {real, imag} */,
  {32'h40b66cd8, 32'hc0eebd18} /* (7, 4, 30) {real, imag} */,
  {32'h4031242c, 32'hc116b1b9} /* (7, 4, 29) {real, imag} */,
  {32'h40228147, 32'h4079401c} /* (7, 4, 28) {real, imag} */,
  {32'hc0919f88, 32'h4195bfb8} /* (7, 4, 27) {real, imag} */,
  {32'h407b0b48, 32'h417727ba} /* (7, 4, 26) {real, imag} */,
  {32'h40ad69b2, 32'h41401461} /* (7, 4, 25) {real, imag} */,
  {32'h408ce075, 32'h416b6e66} /* (7, 4, 24) {real, imag} */,
  {32'hc04f103c, 32'h41666ee7} /* (7, 4, 23) {real, imag} */,
  {32'hc1aafebd, 32'h403a4994} /* (7, 4, 22) {real, imag} */,
  {32'hc13fcb33, 32'h4052dc69} /* (7, 4, 21) {real, imag} */,
  {32'h4129aab9, 32'hc025b591} /* (7, 4, 20) {real, imag} */,
  {32'h41a7198f, 32'hc0af13aa} /* (7, 4, 19) {real, imag} */,
  {32'h40b8fffc, 32'h3f2e6208} /* (7, 4, 18) {real, imag} */,
  {32'h413d66ca, 32'h40a25db6} /* (7, 4, 17) {real, imag} */,
  {32'h417c94d8, 32'h410785df} /* (7, 4, 16) {real, imag} */,
  {32'hc1248a43, 32'hc1a66636} /* (7, 4, 15) {real, imag} */,
  {32'hc106733a, 32'hc1b97982} /* (7, 4, 14) {real, imag} */,
  {32'hc135fce2, 32'hc1450f2a} /* (7, 4, 13) {real, imag} */,
  {32'hc13d7055, 32'h412bb012} /* (7, 4, 12) {real, imag} */,
  {32'h3ef95848, 32'h40e0a2ff} /* (7, 4, 11) {real, imag} */,
  {32'hc16bde76, 32'h4152cd62} /* (7, 4, 10) {real, imag} */,
  {32'hc17f4d29, 32'h41c449bb} /* (7, 4, 9) {real, imag} */,
  {32'h409673b2, 32'h409c6afa} /* (7, 4, 8) {real, imag} */,
  {32'hbfa56728, 32'h41376a13} /* (7, 4, 7) {real, imag} */,
  {32'hbf7ea3a8, 32'hbfe4a3fd} /* (7, 4, 6) {real, imag} */,
  {32'h3f1500fc, 32'hc0aa24ab} /* (7, 4, 5) {real, imag} */,
  {32'h3e1a71e0, 32'h408048fc} /* (7, 4, 4) {real, imag} */,
  {32'hc130cbc6, 32'hc039b2d1} /* (7, 4, 3) {real, imag} */,
  {32'hc0ca6772, 32'hc123434a} /* (7, 4, 2) {real, imag} */,
  {32'h411e3407, 32'hc076dbc6} /* (7, 4, 1) {real, imag} */,
  {32'h40aa6cb6, 32'h4061e914} /* (7, 4, 0) {real, imag} */,
  {32'h3ffc7d38, 32'h40b232ca} /* (7, 3, 31) {real, imag} */,
  {32'h4095eb50, 32'hc0b3cff0} /* (7, 3, 30) {real, imag} */,
  {32'h406eef68, 32'hc172f0d4} /* (7, 3, 29) {real, imag} */,
  {32'hc18b3f23, 32'hc1920fda} /* (7, 3, 28) {real, imag} */,
  {32'hc14a72a4, 32'hc122db6c} /* (7, 3, 27) {real, imag} */,
  {32'h41177267, 32'hc13c9c72} /* (7, 3, 26) {real, imag} */,
  {32'h40b79017, 32'hc0eb484a} /* (7, 3, 25) {real, imag} */,
  {32'h4126abb7, 32'hc10c43c6} /* (7, 3, 24) {real, imag} */,
  {32'h418d1ef3, 32'hc03eb73a} /* (7, 3, 23) {real, imag} */,
  {32'h41817b20, 32'h40b023ec} /* (7, 3, 22) {real, imag} */,
  {32'h4197c586, 32'hc09b291e} /* (7, 3, 21) {real, imag} */,
  {32'h4138e732, 32'h40ade5f5} /* (7, 3, 20) {real, imag} */,
  {32'h40bacc4b, 32'hc15d25e3} /* (7, 3, 19) {real, imag} */,
  {32'hc0654c62, 32'h3ec19074} /* (7, 3, 18) {real, imag} */,
  {32'hc09da851, 32'h4093f7b3} /* (7, 3, 17) {real, imag} */,
  {32'h40e5235e, 32'hc059fda5} /* (7, 3, 16) {real, imag} */,
  {32'h4194a004, 32'h40f81da8} /* (7, 3, 15) {real, imag} */,
  {32'h409fcbdd, 32'hc095c5bf} /* (7, 3, 14) {real, imag} */,
  {32'h3f50f07c, 32'h412b8a7c} /* (7, 3, 13) {real, imag} */,
  {32'hc0675630, 32'h41885052} /* (7, 3, 12) {real, imag} */,
  {32'h40519284, 32'h41587b90} /* (7, 3, 11) {real, imag} */,
  {32'hc0ace0f2, 32'h41a784f0} /* (7, 3, 10) {real, imag} */,
  {32'hc11c1c0c, 32'h4167caee} /* (7, 3, 9) {real, imag} */,
  {32'h41422b2d, 32'hc05e9df4} /* (7, 3, 8) {real, imag} */,
  {32'hc10754ce, 32'hc0759e96} /* (7, 3, 7) {real, imag} */,
  {32'hc18d0a8c, 32'hc183ef39} /* (7, 3, 6) {real, imag} */,
  {32'hc086a66f, 32'hc09e82d4} /* (7, 3, 5) {real, imag} */,
  {32'h40e06d11, 32'h41cc4f93} /* (7, 3, 4) {real, imag} */,
  {32'h4141b68f, 32'h419118da} /* (7, 3, 3) {real, imag} */,
  {32'h3fcd45f4, 32'h40fa8d3e} /* (7, 3, 2) {real, imag} */,
  {32'h41291ae6, 32'hbfa4bb3c} /* (7, 3, 1) {real, imag} */,
  {32'h4113b96b, 32'hc1053be0} /* (7, 3, 0) {real, imag} */,
  {32'hc06ee02f, 32'hc17a5afa} /* (7, 2, 31) {real, imag} */,
  {32'hbf3a7838, 32'hc1449ebc} /* (7, 2, 30) {real, imag} */,
  {32'hc0b4a100, 32'hc0393672} /* (7, 2, 29) {real, imag} */,
  {32'h41112b65, 32'h413d8478} /* (7, 2, 28) {real, imag} */,
  {32'h4095f266, 32'h41947968} /* (7, 2, 27) {real, imag} */,
  {32'hc14d19b7, 32'h419ebbcd} /* (7, 2, 26) {real, imag} */,
  {32'h3fb7a5a8, 32'h413e374d} /* (7, 2, 25) {real, imag} */,
  {32'h41652dbc, 32'hbfcac548} /* (7, 2, 24) {real, imag} */,
  {32'hc0a14c32, 32'h409e9a0c} /* (7, 2, 23) {real, imag} */,
  {32'hbf8bf83c, 32'h416e4767} /* (7, 2, 22) {real, imag} */,
  {32'hc00e3685, 32'h406cfaa6} /* (7, 2, 21) {real, imag} */,
  {32'hc0b44f80, 32'hc1629e34} /* (7, 2, 20) {real, imag} */,
  {32'h4019754b, 32'hc0c453c5} /* (7, 2, 19) {real, imag} */,
  {32'h3ff9c06c, 32'hc1a549d0} /* (7, 2, 18) {real, imag} */,
  {32'hc154469e, 32'hc19d4085} /* (7, 2, 17) {real, imag} */,
  {32'h4034aa4e, 32'hc172f57c} /* (7, 2, 16) {real, imag} */,
  {32'h411e05ec, 32'h410f5636} /* (7, 2, 15) {real, imag} */,
  {32'h41189106, 32'h4164f427} /* (7, 2, 14) {real, imag} */,
  {32'hbfa51eb0, 32'h415ed72c} /* (7, 2, 13) {real, imag} */,
  {32'hc1916ef0, 32'hbe6d8de0} /* (7, 2, 12) {real, imag} */,
  {32'h40ad1403, 32'h3f5ff63c} /* (7, 2, 11) {real, imag} */,
  {32'h3f5d9978, 32'h40408dd6} /* (7, 2, 10) {real, imag} */,
  {32'h3cc4ef00, 32'hc050ed59} /* (7, 2, 9) {real, imag} */,
  {32'h41aa578e, 32'hbe1a9ac8} /* (7, 2, 8) {real, imag} */,
  {32'h41ce4041, 32'h403a70d5} /* (7, 2, 7) {real, imag} */,
  {32'hc08f9da6, 32'h413c3aac} /* (7, 2, 6) {real, imag} */,
  {32'hc0cf7dc4, 32'h419ee58f} /* (7, 2, 5) {real, imag} */,
  {32'hc0b21b4b, 32'h41529140} /* (7, 2, 4) {real, imag} */,
  {32'hc1949b1a, 32'h41227739} /* (7, 2, 3) {real, imag} */,
  {32'hc1713d2c, 32'h413057f3} /* (7, 2, 2) {real, imag} */,
  {32'hc1179af2, 32'hbe88a334} /* (7, 2, 1) {real, imag} */,
  {32'hc0be5cb4, 32'hc101821f} /* (7, 2, 0) {real, imag} */,
  {32'hc0dd6c56, 32'h4085e26b} /* (7, 1, 31) {real, imag} */,
  {32'hc17e1f1c, 32'h40e3e9cc} /* (7, 1, 30) {real, imag} */,
  {32'hc1838f74, 32'hc14ec3e4} /* (7, 1, 29) {real, imag} */,
  {32'h4157cd14, 32'hc0fa8f2e} /* (7, 1, 28) {real, imag} */,
  {32'h41c801df, 32'hc07e81eb} /* (7, 1, 27) {real, imag} */,
  {32'h405191cc, 32'hc1631e90} /* (7, 1, 26) {real, imag} */,
  {32'h3feb32b9, 32'hc197f9c8} /* (7, 1, 25) {real, imag} */,
  {32'h41c24048, 32'hc001a7c4} /* (7, 1, 24) {real, imag} */,
  {32'h414665b7, 32'h40947222} /* (7, 1, 23) {real, imag} */,
  {32'h415b6d45, 32'hc04abcb0} /* (7, 1, 22) {real, imag} */,
  {32'h41285945, 32'hc112b0ba} /* (7, 1, 21) {real, imag} */,
  {32'hc0bf17d4, 32'hc03312c2} /* (7, 1, 20) {real, imag} */,
  {32'hc1a38c38, 32'h420220b5} /* (7, 1, 19) {real, imag} */,
  {32'hc185b6a1, 32'h41c03b18} /* (7, 1, 18) {real, imag} */,
  {32'hc09d2e7b, 32'h4183eab6} /* (7, 1, 17) {real, imag} */,
  {32'hc16de7a5, 32'h41404a8e} /* (7, 1, 16) {real, imag} */,
  {32'hc044affe, 32'h40ec838c} /* (7, 1, 15) {real, imag} */,
  {32'h410726c0, 32'h41be0e6a} /* (7, 1, 14) {real, imag} */,
  {32'hc10654f1, 32'h4207b1c4} /* (7, 1, 13) {real, imag} */,
  {32'hc0860238, 32'h41024fbc} /* (7, 1, 12) {real, imag} */,
  {32'hc0089aa4, 32'hc0b2fa88} /* (7, 1, 11) {real, imag} */,
  {32'h40442f9c, 32'hc0c8be44} /* (7, 1, 10) {real, imag} */,
  {32'hc12d11ee, 32'hc09511e0} /* (7, 1, 9) {real, imag} */,
  {32'h40107b24, 32'h3f170fe0} /* (7, 1, 8) {real, imag} */,
  {32'h41927548, 32'h3faefbd0} /* (7, 1, 7) {real, imag} */,
  {32'h40b2e4d0, 32'h40cb3a28} /* (7, 1, 6) {real, imag} */,
  {32'h3f97980a, 32'h41058140} /* (7, 1, 5) {real, imag} */,
  {32'hc121a2ca, 32'h40085e59} /* (7, 1, 4) {real, imag} */,
  {32'hc1260010, 32'hbfe0e37c} /* (7, 1, 3) {real, imag} */,
  {32'h412cd605, 32'hc045e317} /* (7, 1, 2) {real, imag} */,
  {32'h419e48a2, 32'hbfbf2414} /* (7, 1, 1) {real, imag} */,
  {32'h3ef99090, 32'hc060390e} /* (7, 1, 0) {real, imag} */,
  {32'hc0a69cc0, 32'h4061f937} /* (7, 0, 31) {real, imag} */,
  {32'hc11a8794, 32'hc10fb774} /* (7, 0, 30) {real, imag} */,
  {32'hc13c3481, 32'hc1851be8} /* (7, 0, 29) {real, imag} */,
  {32'hbfdecb38, 32'hc19b5fb1} /* (7, 0, 28) {real, imag} */,
  {32'h40b9b022, 32'hc178125a} /* (7, 0, 27) {real, imag} */,
  {32'hc125b394, 32'h40ab2ed9} /* (7, 0, 26) {real, imag} */,
  {32'hc0e3a228, 32'h418ef86c} /* (7, 0, 25) {real, imag} */,
  {32'h40f1afd9, 32'h4131025c} /* (7, 0, 24) {real, imag} */,
  {32'hc103b926, 32'hbfdff23d} /* (7, 0, 23) {real, imag} */,
  {32'h4106ecec, 32'hc14190fe} /* (7, 0, 22) {real, imag} */,
  {32'h4156bb78, 32'hc19f55f4} /* (7, 0, 21) {real, imag} */,
  {32'h41107f02, 32'hc15c8cd9} /* (7, 0, 20) {real, imag} */,
  {32'hc1348216, 32'hc133ca2e} /* (7, 0, 19) {real, imag} */,
  {32'hc1883bca, 32'hc18328d8} /* (7, 0, 18) {real, imag} */,
  {32'h40be94cc, 32'h4040f3f8} /* (7, 0, 17) {real, imag} */,
  {32'h414a4cf6, 32'hc1650266} /* (7, 0, 16) {real, imag} */,
  {32'hc0c6517b, 32'hc155ca9c} /* (7, 0, 15) {real, imag} */,
  {32'hc0d2c60e, 32'hc135a194} /* (7, 0, 14) {real, imag} */,
  {32'hc196ae04, 32'hc12be29b} /* (7, 0, 13) {real, imag} */,
  {32'hc17809be, 32'hc0a14da4} /* (7, 0, 12) {real, imag} */,
  {32'h402ff965, 32'h3f771c8e} /* (7, 0, 11) {real, imag} */,
  {32'h3ff122be, 32'h3fdb53dc} /* (7, 0, 10) {real, imag} */,
  {32'h416c8d23, 32'hbf7801c0} /* (7, 0, 9) {real, imag} */,
  {32'hbf8dca18, 32'h40da92ff} /* (7, 0, 8) {real, imag} */,
  {32'hbeff1a60, 32'h41217526} /* (7, 0, 7) {real, imag} */,
  {32'h3ca5cfc0, 32'hc19e36d0} /* (7, 0, 6) {real, imag} */,
  {32'h4166746f, 32'hc107d14e} /* (7, 0, 5) {real, imag} */,
  {32'h3fcbe6d5, 32'hc02a3e5a} /* (7, 0, 4) {real, imag} */,
  {32'h3fb61f30, 32'hc0d4c4f4} /* (7, 0, 3) {real, imag} */,
  {32'h40194518, 32'h40eb00b1} /* (7, 0, 2) {real, imag} */,
  {32'h418df6e2, 32'h4101fe1a} /* (7, 0, 1) {real, imag} */,
  {32'h40674965, 32'h409b5f46} /* (7, 0, 0) {real, imag} */,
  {32'h3f4cb118, 32'h40b1eeac} /* (6, 31, 31) {real, imag} */,
  {32'hbfa1a878, 32'h4056accf} /* (6, 31, 30) {real, imag} */,
  {32'hc103e3d3, 32'hbf3d058a} /* (6, 31, 29) {real, imag} */,
  {32'hc0f56ec9, 32'hc1a33adb} /* (6, 31, 28) {real, imag} */,
  {32'hc1269eb8, 32'hc173d757} /* (6, 31, 27) {real, imag} */,
  {32'hc1a35916, 32'hc0c76e7a} /* (6, 31, 26) {real, imag} */,
  {32'hc0e17af0, 32'hbfba1ea6} /* (6, 31, 25) {real, imag} */,
  {32'hc0403af2, 32'hc09df412} /* (6, 31, 24) {real, imag} */,
  {32'hc0af60a2, 32'hc114f432} /* (6, 31, 23) {real, imag} */,
  {32'hc094e1ef, 32'h40cf11f0} /* (6, 31, 22) {real, imag} */,
  {32'h41110236, 32'hc14d2c9d} /* (6, 31, 21) {real, imag} */,
  {32'hc1609c78, 32'hc08800cc} /* (6, 31, 20) {real, imag} */,
  {32'hc1467dba, 32'h411b3568} /* (6, 31, 19) {real, imag} */,
  {32'hbf03d27c, 32'h419155a4} /* (6, 31, 18) {real, imag} */,
  {32'hc196868e, 32'h41cf992a} /* (6, 31, 17) {real, imag} */,
  {32'hc1b603b9, 32'h4013a06a} /* (6, 31, 16) {real, imag} */,
  {32'hc0abbe60, 32'h3f3fb340} /* (6, 31, 15) {real, imag} */,
  {32'h41676966, 32'h418f21d8} /* (6, 31, 14) {real, imag} */,
  {32'h41bda3ae, 32'hc0e3f45b} /* (6, 31, 13) {real, imag} */,
  {32'h41501e8e, 32'hc1b18fea} /* (6, 31, 12) {real, imag} */,
  {32'h41378bd1, 32'hc2114199} /* (6, 31, 11) {real, imag} */,
  {32'h41030f1e, 32'hc1579c96} /* (6, 31, 10) {real, imag} */,
  {32'hc1df3017, 32'h418f2879} /* (6, 31, 9) {real, imag} */,
  {32'hc189659e, 32'h41d3290c} /* (6, 31, 8) {real, imag} */,
  {32'hc1928725, 32'h41adca2e} /* (6, 31, 7) {real, imag} */,
  {32'hc209544b, 32'h40de4796} /* (6, 31, 6) {real, imag} */,
  {32'hc190b8d4, 32'h3fd7285b} /* (6, 31, 5) {real, imag} */,
  {32'hc11bb85b, 32'hc0cdc9dd} /* (6, 31, 4) {real, imag} */,
  {32'hc0406b4a, 32'hc0ad76de} /* (6, 31, 3) {real, imag} */,
  {32'h3f8ffb88, 32'hc1446024} /* (6, 31, 2) {real, imag} */,
  {32'hc0d8780e, 32'hc04fa0b4} /* (6, 31, 1) {real, imag} */,
  {32'hbf4247d8, 32'h40d7cd4e} /* (6, 31, 0) {real, imag} */,
  {32'h40e5c77d, 32'hbfe88c50} /* (6, 30, 31) {real, imag} */,
  {32'h40fb6bde, 32'h4111ec11} /* (6, 30, 30) {real, imag} */,
  {32'hbfd3ef24, 32'h413ba7ee} /* (6, 30, 29) {real, imag} */,
  {32'hc085443c, 32'h411fe752} /* (6, 30, 28) {real, imag} */,
  {32'h3cc0ee00, 32'h40864398} /* (6, 30, 27) {real, imag} */,
  {32'hc1d36fce, 32'h4026e2a8} /* (6, 30, 26) {real, imag} */,
  {32'hc198feb1, 32'h416b8b2b} /* (6, 30, 25) {real, imag} */,
  {32'hc083e89f, 32'h4197a47a} /* (6, 30, 24) {real, imag} */,
  {32'hc119cf10, 32'h410fe09c} /* (6, 30, 23) {real, imag} */,
  {32'hc1638bd3, 32'h40024fce} /* (6, 30, 22) {real, imag} */,
  {32'hc104c07d, 32'h4064d072} /* (6, 30, 21) {real, imag} */,
  {32'h40fa3fa4, 32'h412039ff} /* (6, 30, 20) {real, imag} */,
  {32'h4146f9ea, 32'h41bc1922} /* (6, 30, 19) {real, imag} */,
  {32'h41a0ee79, 32'h410c3dda} /* (6, 30, 18) {real, imag} */,
  {32'h41e5f4a5, 32'hc06becb1} /* (6, 30, 17) {real, imag} */,
  {32'h3ec394e0, 32'hc19d3b20} /* (6, 30, 16) {real, imag} */,
  {32'hc182fa44, 32'hc1e7e815} /* (6, 30, 15) {real, imag} */,
  {32'hc188a04c, 32'hc1de838c} /* (6, 30, 14) {real, imag} */,
  {32'hc1fe859b, 32'hc18e06df} /* (6, 30, 13) {real, imag} */,
  {32'hc08388b2, 32'h40c8b9be} /* (6, 30, 12) {real, imag} */,
  {32'hbf0fd540, 32'h3fb24248} /* (6, 30, 11) {real, imag} */,
  {32'hc0c95ac7, 32'hc18caaf0} /* (6, 30, 10) {real, imag} */,
  {32'hbf74acb6, 32'h3fcf72d0} /* (6, 30, 9) {real, imag} */,
  {32'hc11de2f6, 32'h40c36f24} /* (6, 30, 8) {real, imag} */,
  {32'hc170dfaa, 32'hc136a7ee} /* (6, 30, 7) {real, imag} */,
  {32'hc1418a0b, 32'hc1074e44} /* (6, 30, 6) {real, imag} */,
  {32'hc0aa50dc, 32'hc1066a40} /* (6, 30, 5) {real, imag} */,
  {32'h40dab4cc, 32'hc0f18f30} /* (6, 30, 4) {real, imag} */,
  {32'h40b1a17e, 32'hc13c5cf2} /* (6, 30, 3) {real, imag} */,
  {32'h4140ebfc, 32'hc14e8e4a} /* (6, 30, 2) {real, imag} */,
  {32'h4193bd80, 32'h4026480c} /* (6, 30, 1) {real, imag} */,
  {32'hc0a6e75f, 32'hbec1ff98} /* (6, 30, 0) {real, imag} */,
  {32'h3ef98a20, 32'hc0d8a513} /* (6, 29, 31) {real, imag} */,
  {32'h412c255a, 32'h403a5914} /* (6, 29, 30) {real, imag} */,
  {32'h4194c342, 32'h40e53c06} /* (6, 29, 29) {real, imag} */,
  {32'h4185704b, 32'hc14272fe} /* (6, 29, 28) {real, imag} */,
  {32'h4190e528, 32'hc17e432c} /* (6, 29, 27) {real, imag} */,
  {32'hbfd08c61, 32'hc21bea0b} /* (6, 29, 26) {real, imag} */,
  {32'hc025f056, 32'hc1963274} /* (6, 29, 25) {real, imag} */,
  {32'h40f53464, 32'hc19e9a3a} /* (6, 29, 24) {real, imag} */,
  {32'h4095fc40, 32'hc1c192c4} /* (6, 29, 23) {real, imag} */,
  {32'h40ff2b27, 32'hbff164bd} /* (6, 29, 22) {real, imag} */,
  {32'h41c913d8, 32'hc13042cb} /* (6, 29, 21) {real, imag} */,
  {32'h41d872cc, 32'hc11dface} /* (6, 29, 20) {real, imag} */,
  {32'h40dedc58, 32'hbed3f348} /* (6, 29, 19) {real, imag} */,
  {32'hbfebaa7b, 32'hc16004d8} /* (6, 29, 18) {real, imag} */,
  {32'h3ff93b7f, 32'h40661398} /* (6, 29, 17) {real, imag} */,
  {32'hbf269de8, 32'h41c9d354} /* (6, 29, 16) {real, imag} */,
  {32'hc037bab0, 32'hbf5374ec} /* (6, 29, 15) {real, imag} */,
  {32'hc0fdcc4e, 32'hc10872f5} /* (6, 29, 14) {real, imag} */,
  {32'hbfdc4be2, 32'hc028b130} /* (6, 29, 13) {real, imag} */,
  {32'h4132e710, 32'hbfd1d566} /* (6, 29, 12) {real, imag} */,
  {32'h413043ec, 32'h410ac3d2} /* (6, 29, 11) {real, imag} */,
  {32'h4034c0e6, 32'h3fe002f8} /* (6, 29, 10) {real, imag} */,
  {32'h411aed3a, 32'h3fdeb520} /* (6, 29, 9) {real, imag} */,
  {32'h40d7972a, 32'hc16f686e} /* (6, 29, 8) {real, imag} */,
  {32'hc1857ae2, 32'hc1df3c33} /* (6, 29, 7) {real, imag} */,
  {32'hc06852f5, 32'hc1ed0a96} /* (6, 29, 6) {real, imag} */,
  {32'hc08252c6, 32'hc09e1d77} /* (6, 29, 5) {real, imag} */,
  {32'hc0a41a4c, 32'hc1501f60} /* (6, 29, 4) {real, imag} */,
  {32'h4032bdfc, 32'hc205b232} /* (6, 29, 3) {real, imag} */,
  {32'h411cb164, 32'h3f9f4a44} /* (6, 29, 2) {real, imag} */,
  {32'h401eb9cc, 32'h4052fe16} /* (6, 29, 1) {real, imag} */,
  {32'h4151d805, 32'hc076e838} /* (6, 29, 0) {real, imag} */,
  {32'h402ff809, 32'hc0bbf74c} /* (6, 28, 31) {real, imag} */,
  {32'hc0c5a772, 32'hc1039e03} /* (6, 28, 30) {real, imag} */,
  {32'hbfa94e4a, 32'h406286e8} /* (6, 28, 29) {real, imag} */,
  {32'h4192aec9, 32'h3f428b60} /* (6, 28, 28) {real, imag} */,
  {32'hbe995ac0, 32'hc1a60f1a} /* (6, 28, 27) {real, imag} */,
  {32'hc1e5fa36, 32'hc0fb5180} /* (6, 28, 26) {real, imag} */,
  {32'hc10a08e3, 32'hc0c8b63e} /* (6, 28, 25) {real, imag} */,
  {32'h4126394c, 32'hbff24d26} /* (6, 28, 24) {real, imag} */,
  {32'h41bbf36a, 32'h413331fa} /* (6, 28, 23) {real, imag} */,
  {32'h40cccf9f, 32'hc00e85a8} /* (6, 28, 22) {real, imag} */,
  {32'h41276c84, 32'hc123e724} /* (6, 28, 21) {real, imag} */,
  {32'h411bfc0c, 32'h413af9d0} /* (6, 28, 20) {real, imag} */,
  {32'h41a6e897, 32'h418fc288} /* (6, 28, 19) {real, imag} */,
  {32'h410c0c73, 32'h41c65d28} /* (6, 28, 18) {real, imag} */,
  {32'hc14e8c9b, 32'h4162cf26} /* (6, 28, 17) {real, imag} */,
  {32'hbfd80ed8, 32'h3f192560} /* (6, 28, 16) {real, imag} */,
  {32'hc10abc8a, 32'hc017c9ce} /* (6, 28, 15) {real, imag} */,
  {32'h4127ab9e, 32'hc028d8a0} /* (6, 28, 14) {real, imag} */,
  {32'h41b2e218, 32'hc11559be} /* (6, 28, 13) {real, imag} */,
  {32'hc0610fb2, 32'hc0acae97} /* (6, 28, 12) {real, imag} */,
  {32'hbfdaab0c, 32'hc085b313} /* (6, 28, 11) {real, imag} */,
  {32'hc0913ee8, 32'hc13ecb89} /* (6, 28, 10) {real, imag} */,
  {32'h40eca36f, 32'hc009de92} /* (6, 28, 9) {real, imag} */,
  {32'h41a7923c, 32'hc0ec49e8} /* (6, 28, 8) {real, imag} */,
  {32'hbee745fa, 32'h4028fe5c} /* (6, 28, 7) {real, imag} */,
  {32'hc0e940bc, 32'h40e531b2} /* (6, 28, 6) {real, imag} */,
  {32'hc1cdfd1f, 32'h40a2a165} /* (6, 28, 5) {real, imag} */,
  {32'hc1f60ab2, 32'h409cc9e4} /* (6, 28, 4) {real, imag} */,
  {32'hc1a29d2f, 32'h4177a74a} /* (6, 28, 3) {real, imag} */,
  {32'hc17dde4f, 32'h3fdeb4a8} /* (6, 28, 2) {real, imag} */,
  {32'h410d2e58, 32'h410aa95e} /* (6, 28, 1) {real, imag} */,
  {32'h4176fe96, 32'hc0db124a} /* (6, 28, 0) {real, imag} */,
  {32'hc129723d, 32'hc0952ea0} /* (6, 27, 31) {real, imag} */,
  {32'hc1266294, 32'hbfde89f4} /* (6, 27, 30) {real, imag} */,
  {32'h4140a3b9, 32'h40431660} /* (6, 27, 29) {real, imag} */,
  {32'h3fef3b08, 32'h40c7730f} /* (6, 27, 28) {real, imag} */,
  {32'h40afb832, 32'h406875fd} /* (6, 27, 27) {real, imag} */,
  {32'hc00fc14d, 32'hc05f77d2} /* (6, 27, 26) {real, imag} */,
  {32'hc17b50b0, 32'hc0a7e908} /* (6, 27, 25) {real, imag} */,
  {32'hc1634d14, 32'hc0abc93c} /* (6, 27, 24) {real, imag} */,
  {32'hc16c8ad8, 32'h4062b814} /* (6, 27, 23) {real, imag} */,
  {32'hc1192b67, 32'h4090e0c0} /* (6, 27, 22) {real, imag} */,
  {32'h40be0b89, 32'hbf7c5da0} /* (6, 27, 21) {real, imag} */,
  {32'h3fedada8, 32'hc1608ffa} /* (6, 27, 20) {real, imag} */,
  {32'h4097e726, 32'h40ef071a} /* (6, 27, 19) {real, imag} */,
  {32'hc071f4cd, 32'hc0b03b96} /* (6, 27, 18) {real, imag} */,
  {32'hc059f602, 32'hc18fca1c} /* (6, 27, 17) {real, imag} */,
  {32'h4131accf, 32'hc0734edd} /* (6, 27, 16) {real, imag} */,
  {32'h41393c17, 32'h3fa3e838} /* (6, 27, 15) {real, imag} */,
  {32'h41480abf, 32'hc05340f3} /* (6, 27, 14) {real, imag} */,
  {32'h412504c4, 32'hc14579e9} /* (6, 27, 13) {real, imag} */,
  {32'h4116767a, 32'hc0beadc9} /* (6, 27, 12) {real, imag} */,
  {32'h41167640, 32'h41066590} /* (6, 27, 11) {real, imag} */,
  {32'hc04bc174, 32'h40ba0186} /* (6, 27, 10) {real, imag} */,
  {32'hc0b75426, 32'h4168b77c} /* (6, 27, 9) {real, imag} */,
  {32'h400d1ccb, 32'hc182c698} /* (6, 27, 8) {real, imag} */,
  {32'hc0821f99, 32'hc1608f62} /* (6, 27, 7) {real, imag} */,
  {32'hc117c016, 32'h3fd0d505} /* (6, 27, 6) {real, imag} */,
  {32'h4045e824, 32'hc161bc6e} /* (6, 27, 5) {real, imag} */,
  {32'h3fa00d4d, 32'hc16fce8c} /* (6, 27, 4) {real, imag} */,
  {32'h409fcb70, 32'hc059fae4} /* (6, 27, 3) {real, imag} */,
  {32'h40ab8468, 32'h402924d7} /* (6, 27, 2) {real, imag} */,
  {32'hc0256803, 32'hc0ce1870} /* (6, 27, 1) {real, imag} */,
  {32'hbee12890, 32'hc141fafc} /* (6, 27, 0) {real, imag} */,
  {32'h40a42601, 32'h3fd02962} /* (6, 26, 31) {real, imag} */,
  {32'h411446c5, 32'hc0c68864} /* (6, 26, 30) {real, imag} */,
  {32'h401ba4a2, 32'hc0e5653c} /* (6, 26, 29) {real, imag} */,
  {32'h3fc688ec, 32'h3f962470} /* (6, 26, 28) {real, imag} */,
  {32'hc11ab2e6, 32'h41181b7d} /* (6, 26, 27) {real, imag} */,
  {32'h4011068f, 32'h40d59833} /* (6, 26, 26) {real, imag} */,
  {32'h40f210ff, 32'h40f98a3f} /* (6, 26, 25) {real, imag} */,
  {32'h410a20be, 32'h40f3a0a9} /* (6, 26, 24) {real, imag} */,
  {32'h412be26e, 32'h4069083f} /* (6, 26, 23) {real, imag} */,
  {32'h412b183e, 32'h4158067c} /* (6, 26, 22) {real, imag} */,
  {32'h418c07e6, 32'h418bf0ef} /* (6, 26, 21) {real, imag} */,
  {32'h3ff45b8c, 32'h4103a24e} /* (6, 26, 20) {real, imag} */,
  {32'hc19ec9a6, 32'hc10e5b79} /* (6, 26, 19) {real, imag} */,
  {32'hc135e110, 32'hc0ad9789} /* (6, 26, 18) {real, imag} */,
  {32'hc19e2ef0, 32'h4150d056} /* (6, 26, 17) {real, imag} */,
  {32'hc13077e0, 32'h41375a5e} /* (6, 26, 16) {real, imag} */,
  {32'hc0740e2d, 32'h414e54e5} /* (6, 26, 15) {real, imag} */,
  {32'h40ae15d3, 32'h405fec1e} /* (6, 26, 14) {real, imag} */,
  {32'hc052e7c4, 32'h414d9a4c} /* (6, 26, 13) {real, imag} */,
  {32'hc0dddac2, 32'h41c24292} /* (6, 26, 12) {real, imag} */,
  {32'h40caff84, 32'h4179bcad} /* (6, 26, 11) {real, imag} */,
  {32'hc0184afc, 32'h40963d32} /* (6, 26, 10) {real, imag} */,
  {32'hc0f6ba68, 32'hc0eff284} /* (6, 26, 9) {real, imag} */,
  {32'hbf17c53c, 32'hbfa19fc0} /* (6, 26, 8) {real, imag} */,
  {32'hc0d5d6d4, 32'h40ce029a} /* (6, 26, 7) {real, imag} */,
  {32'h4126538c, 32'hc0e75831} /* (6, 26, 6) {real, imag} */,
  {32'h41895b51, 32'hc17ef97b} /* (6, 26, 5) {real, imag} */,
  {32'h3d3dbce0, 32'hbf5e2cfa} /* (6, 26, 4) {real, imag} */,
  {32'hc11f0f6d, 32'h410d479b} /* (6, 26, 3) {real, imag} */,
  {32'hc0983b7e, 32'h411954c0} /* (6, 26, 2) {real, imag} */,
  {32'h417c324c, 32'h40f1c73c} /* (6, 26, 1) {real, imag} */,
  {32'h413c8bcf, 32'h40f50c6e} /* (6, 26, 0) {real, imag} */,
  {32'hc017e082, 32'hbf3d5284} /* (6, 25, 31) {real, imag} */,
  {32'hc01ca7eb, 32'hc05a3dd7} /* (6, 25, 30) {real, imag} */,
  {32'hc0115609, 32'hc01431fd} /* (6, 25, 29) {real, imag} */,
  {32'hc1600dd0, 32'hc0eb7f71} /* (6, 25, 28) {real, imag} */,
  {32'h40184380, 32'hc159cd0a} /* (6, 25, 27) {real, imag} */,
  {32'h40cc580f, 32'hc11348ed} /* (6, 25, 26) {real, imag} */,
  {32'h4134c2da, 32'hc10d74bb} /* (6, 25, 25) {real, imag} */,
  {32'h4077d78f, 32'h4003e762} /* (6, 25, 24) {real, imag} */,
  {32'h3faee58c, 32'h40366492} /* (6, 25, 23) {real, imag} */,
  {32'hc093b6c0, 32'hbf1c6330} /* (6, 25, 22) {real, imag} */,
  {32'h3d797000, 32'hc027453c} /* (6, 25, 21) {real, imag} */,
  {32'hc1367e0f, 32'h41386ee4} /* (6, 25, 20) {real, imag} */,
  {32'hc157250f, 32'h413bc0ab} /* (6, 25, 19) {real, imag} */,
  {32'h3f9ac7af, 32'h4005b41c} /* (6, 25, 18) {real, imag} */,
  {32'hc0c690db, 32'hc163c8e6} /* (6, 25, 17) {real, imag} */,
  {32'hc1a50d35, 32'hbfc0d390} /* (6, 25, 16) {real, imag} */,
  {32'hc0f98d50, 32'h40050276} /* (6, 25, 15) {real, imag} */,
  {32'hc0c80056, 32'h40acb9da} /* (6, 25, 14) {real, imag} */,
  {32'h4087af16, 32'h414503a0} /* (6, 25, 13) {real, imag} */,
  {32'h404fd7aa, 32'h41074f2c} /* (6, 25, 12) {real, imag} */,
  {32'hc097f1bd, 32'h4097c083} /* (6, 25, 11) {real, imag} */,
  {32'hc0cd0b96, 32'hc0367316} /* (6, 25, 10) {real, imag} */,
  {32'hbf1288b0, 32'hc12f31f7} /* (6, 25, 9) {real, imag} */,
  {32'hc099f1bb, 32'hbfa8c2d8} /* (6, 25, 8) {real, imag} */,
  {32'hc177b182, 32'h4064f110} /* (6, 25, 7) {real, imag} */,
  {32'h403df950, 32'hc0f7380b} /* (6, 25, 6) {real, imag} */,
  {32'h3fc8f348, 32'hc182634f} /* (6, 25, 5) {real, imag} */,
  {32'h415d26ec, 32'hc0cf2b81} /* (6, 25, 4) {real, imag} */,
  {32'h4147ab39, 32'hc1058f5d} /* (6, 25, 3) {real, imag} */,
  {32'h4113b8b9, 32'hc12cc460} /* (6, 25, 2) {real, imag} */,
  {32'h40c9f12f, 32'hc1273ed3} /* (6, 25, 1) {real, imag} */,
  {32'hc06eccbc, 32'hc109b830} /* (6, 25, 0) {real, imag} */,
  {32'h408135a8, 32'h411c83e0} /* (6, 24, 31) {real, imag} */,
  {32'h402e4563, 32'h413f180e} /* (6, 24, 30) {real, imag} */,
  {32'h41321550, 32'hc04e4071} /* (6, 24, 29) {real, imag} */,
  {32'h418c0d18, 32'h4104f3c7} /* (6, 24, 28) {real, imag} */,
  {32'h40c5340a, 32'h41868328} /* (6, 24, 27) {real, imag} */,
  {32'hc01584f8, 32'h40e998af} /* (6, 24, 26) {real, imag} */,
  {32'h41166bf3, 32'h40832ac0} /* (6, 24, 25) {real, imag} */,
  {32'h408d69e1, 32'h40a32d80} /* (6, 24, 24) {real, imag} */,
  {32'h40f9b8f2, 32'hc08fd5e9} /* (6, 24, 23) {real, imag} */,
  {32'h40925626, 32'hc09e457e} /* (6, 24, 22) {real, imag} */,
  {32'hc0865e46, 32'hc1a3eb6d} /* (6, 24, 21) {real, imag} */,
  {32'hc1c80861, 32'hc02c2c7a} /* (6, 24, 20) {real, imag} */,
  {32'hc0d56a7a, 32'hc07edc4c} /* (6, 24, 19) {real, imag} */,
  {32'h409bedae, 32'hc0e71f0c} /* (6, 24, 18) {real, imag} */,
  {32'hc02e8b92, 32'h3e5966f0} /* (6, 24, 17) {real, imag} */,
  {32'h40a4eb5a, 32'h402559f0} /* (6, 24, 16) {real, imag} */,
  {32'h411681b3, 32'h40e34396} /* (6, 24, 15) {real, imag} */,
  {32'h419f2358, 32'h41225ec9} /* (6, 24, 14) {real, imag} */,
  {32'h4191f5fc, 32'h41359561} /* (6, 24, 13) {real, imag} */,
  {32'h4120499e, 32'h3ec53cd0} /* (6, 24, 12) {real, imag} */,
  {32'h4116f0a9, 32'hc0a12d3d} /* (6, 24, 11) {real, imag} */,
  {32'h4169551a, 32'h3f7de650} /* (6, 24, 10) {real, imag} */,
  {32'h4169c8c0, 32'h3ef89e78} /* (6, 24, 9) {real, imag} */,
  {32'h40f828dc, 32'h4148ebf0} /* (6, 24, 8) {real, imag} */,
  {32'h40813cec, 32'h40e586cd} /* (6, 24, 7) {real, imag} */,
  {32'h3fb63820, 32'hc0392278} /* (6, 24, 6) {real, imag} */,
  {32'hc0aa6147, 32'hc0921ed7} /* (6, 24, 5) {real, imag} */,
  {32'hc13d5136, 32'h40a3db8f} /* (6, 24, 4) {real, imag} */,
  {32'hc12f6125, 32'h3fddd158} /* (6, 24, 3) {real, imag} */,
  {32'hc0e4000d, 32'hc0d85344} /* (6, 24, 2) {real, imag} */,
  {32'hc041d274, 32'hc11c1d8d} /* (6, 24, 1) {real, imag} */,
  {32'h3f3632c8, 32'hc11d2a28} /* (6, 24, 0) {real, imag} */,
  {32'h40ebe684, 32'h4096f642} /* (6, 23, 31) {real, imag} */,
  {32'h40c59f5e, 32'hc045203c} /* (6, 23, 30) {real, imag} */,
  {32'h40b61b00, 32'hc01a40c8} /* (6, 23, 29) {real, imag} */,
  {32'hc039ce7c, 32'hc0271a46} /* (6, 23, 28) {real, imag} */,
  {32'h3e5e3700, 32'h41002da4} /* (6, 23, 27) {real, imag} */,
  {32'h3faaf062, 32'h3f2fc118} /* (6, 23, 26) {real, imag} */,
  {32'hc104f668, 32'hc0be0926} /* (6, 23, 25) {real, imag} */,
  {32'hc0b30193, 32'hbfff6318} /* (6, 23, 24) {real, imag} */,
  {32'h410ed7f7, 32'h40b0ef3b} /* (6, 23, 23) {real, imag} */,
  {32'h40c7fe6d, 32'h403fe23a} /* (6, 23, 22) {real, imag} */,
  {32'h407b2d94, 32'h3fcd1db9} /* (6, 23, 21) {real, imag} */,
  {32'hbf9f28e4, 32'h406e92d6} /* (6, 23, 20) {real, imag} */,
  {32'h410069a4, 32'hc103ed56} /* (6, 23, 19) {real, imag} */,
  {32'h4114f3dd, 32'hc0f96d7b} /* (6, 23, 18) {real, imag} */,
  {32'h41073392, 32'hbe8ca320} /* (6, 23, 17) {real, imag} */,
  {32'hc0c1e945, 32'hc1487d5e} /* (6, 23, 16) {real, imag} */,
  {32'hc1150466, 32'hc0f45c47} /* (6, 23, 15) {real, imag} */,
  {32'h402f7a38, 32'h3e10eb10} /* (6, 23, 14) {real, imag} */,
  {32'hc02fd9ac, 32'h3fbcb6dc} /* (6, 23, 13) {real, imag} */,
  {32'h3f9fd564, 32'hbd94fdc0} /* (6, 23, 12) {real, imag} */,
  {32'h40a003bc, 32'h3fdb33bc} /* (6, 23, 11) {real, imag} */,
  {32'hbfb4d5f8, 32'hbfeb26dd} /* (6, 23, 10) {real, imag} */,
  {32'hc105bbc0, 32'h40aa4976} /* (6, 23, 9) {real, imag} */,
  {32'hc080a0dc, 32'h3e40d690} /* (6, 23, 8) {real, imag} */,
  {32'h410bc071, 32'h409a5a82} /* (6, 23, 7) {real, imag} */,
  {32'h4009aeb8, 32'h4110a784} /* (6, 23, 6) {real, imag} */,
  {32'h40b528ac, 32'hc097777e} /* (6, 23, 5) {real, imag} */,
  {32'h403dbe17, 32'hc10bae2d} /* (6, 23, 4) {real, imag} */,
  {32'h3ed9bf50, 32'hc0bb0fec} /* (6, 23, 3) {real, imag} */,
  {32'hc1169b5a, 32'hc153501c} /* (6, 23, 2) {real, imag} */,
  {32'h40e2500f, 32'hc0bac326} /* (6, 23, 1) {real, imag} */,
  {32'h410b8624, 32'hbf661a48} /* (6, 23, 0) {real, imag} */,
  {32'h3f4e30cc, 32'h40252a54} /* (6, 22, 31) {real, imag} */,
  {32'hc0303d16, 32'h409df6f2} /* (6, 22, 30) {real, imag} */,
  {32'hc0959306, 32'h406d8a13} /* (6, 22, 29) {real, imag} */,
  {32'h402e92c5, 32'hc0ba5bda} /* (6, 22, 28) {real, imag} */,
  {32'hc1348eb0, 32'hc0b97e2e} /* (6, 22, 27) {real, imag} */,
  {32'hc11ecf50, 32'h3fa87c48} /* (6, 22, 26) {real, imag} */,
  {32'hbfb0ee44, 32'h405ea486} /* (6, 22, 25) {real, imag} */,
  {32'h4106dda0, 32'hbf3e8c98} /* (6, 22, 24) {real, imag} */,
  {32'h3e2d89b0, 32'hc08aa3e6} /* (6, 22, 23) {real, imag} */,
  {32'h4116eda9, 32'hc0e54ac5} /* (6, 22, 22) {real, imag} */,
  {32'h41555e69, 32'hc09abaf6} /* (6, 22, 21) {real, imag} */,
  {32'hbf9f6430, 32'h40a75678} /* (6, 22, 20) {real, imag} */,
  {32'hc13cbdf1, 32'h408c2d46} /* (6, 22, 19) {real, imag} */,
  {32'hc0eb221a, 32'h3f0621bc} /* (6, 22, 18) {real, imag} */,
  {32'hc08b34e8, 32'hc0ccc949} /* (6, 22, 17) {real, imag} */,
  {32'h3f0f69a8, 32'hc0c41782} /* (6, 22, 16) {real, imag} */,
  {32'hc166cfb8, 32'hc105e684} /* (6, 22, 15) {real, imag} */,
  {32'hc13666ef, 32'h40432518} /* (6, 22, 14) {real, imag} */,
  {32'h407c594e, 32'h40dda910} /* (6, 22, 13) {real, imag} */,
  {32'h41440804, 32'h4097e97f} /* (6, 22, 12) {real, imag} */,
  {32'h40802cc0, 32'hc099dfbc} /* (6, 22, 11) {real, imag} */,
  {32'hc0b31ce8, 32'hc07accdb} /* (6, 22, 10) {real, imag} */,
  {32'hc02f595b, 32'h3f47c8fc} /* (6, 22, 9) {real, imag} */,
  {32'hc0334bfc, 32'hbfdaba72} /* (6, 22, 8) {real, imag} */,
  {32'hc0c52ee8, 32'hc0ec4683} /* (6, 22, 7) {real, imag} */,
  {32'hc08c5318, 32'hc11580f2} /* (6, 22, 6) {real, imag} */,
  {32'h3fbf3b04, 32'hc00e98e7} /* (6, 22, 5) {real, imag} */,
  {32'hc0463cc3, 32'h4087ee8a} /* (6, 22, 4) {real, imag} */,
  {32'hc0e03b06, 32'h3fadf256} /* (6, 22, 3) {real, imag} */,
  {32'hc1049921, 32'hc08ccbb0} /* (6, 22, 2) {real, imag} */,
  {32'hc03a6fb2, 32'h3f4c85dc} /* (6, 22, 1) {real, imag} */,
  {32'h4090d19e, 32'h3fce1c7c} /* (6, 22, 0) {real, imag} */,
  {32'h3f097fd4, 32'hbf80c891} /* (6, 21, 31) {real, imag} */,
  {32'hbeb93150, 32'h3f5feae4} /* (6, 21, 30) {real, imag} */,
  {32'h3fdc80c0, 32'hc001d3a3} /* (6, 21, 29) {real, imag} */,
  {32'h40e30b04, 32'h3e3a7dc8} /* (6, 21, 28) {real, imag} */,
  {32'hc0333380, 32'hbd00cac0} /* (6, 21, 27) {real, imag} */,
  {32'hc1269cda, 32'h40e96288} /* (6, 21, 26) {real, imag} */,
  {32'hbfaefe04, 32'h3f38e94b} /* (6, 21, 25) {real, imag} */,
  {32'h40febac9, 32'h3f617420} /* (6, 21, 24) {real, imag} */,
  {32'h4013d6bd, 32'h413a9498} /* (6, 21, 23) {real, imag} */,
  {32'hc091d7b3, 32'h40a86e37} /* (6, 21, 22) {real, imag} */,
  {32'hc0142978, 32'h41055eaa} /* (6, 21, 21) {real, imag} */,
  {32'h40929522, 32'h40906de3} /* (6, 21, 20) {real, imag} */,
  {32'h3f78ffde, 32'hc0807dc6} /* (6, 21, 19) {real, imag} */,
  {32'h3f1c6274, 32'hbfdb4e02} /* (6, 21, 18) {real, imag} */,
  {32'h40a09d80, 32'hc02bf4cb} /* (6, 21, 17) {real, imag} */,
  {32'h40c6d044, 32'hc0be9b5a} /* (6, 21, 16) {real, imag} */,
  {32'h40bfe958, 32'hc0b1faa2} /* (6, 21, 15) {real, imag} */,
  {32'h40af0c01, 32'hc0bfe527} /* (6, 21, 14) {real, imag} */,
  {32'h407b8a90, 32'h40013329} /* (6, 21, 13) {real, imag} */,
  {32'hbfd56723, 32'hbd4451a0} /* (6, 21, 12) {real, imag} */,
  {32'h401dc84a, 32'hbf263a64} /* (6, 21, 11) {real, imag} */,
  {32'h3fcb9020, 32'hc1299124} /* (6, 21, 10) {real, imag} */,
  {32'hc03d4e06, 32'hc0f9496c} /* (6, 21, 9) {real, imag} */,
  {32'hc09cb136, 32'hc16357f6} /* (6, 21, 8) {real, imag} */,
  {32'h4092cc3f, 32'hc0cfd8a0} /* (6, 21, 7) {real, imag} */,
  {32'h3e2cc120, 32'h4073f5dc} /* (6, 21, 6) {real, imag} */,
  {32'hc0880d3e, 32'h40a4fbce} /* (6, 21, 5) {real, imag} */,
  {32'h407def1a, 32'h410c740e} /* (6, 21, 4) {real, imag} */,
  {32'h40cafd96, 32'h40a2ed94} /* (6, 21, 3) {real, imag} */,
  {32'h4082c50a, 32'h406fbeb3} /* (6, 21, 2) {real, imag} */,
  {32'hbf3318fa, 32'hbf5f1e6c} /* (6, 21, 1) {real, imag} */,
  {32'hc0a30ada, 32'hc0b77dd4} /* (6, 21, 0) {real, imag} */,
  {32'hbddc9880, 32'h40a8a5e7} /* (6, 20, 31) {real, imag} */,
  {32'h400032c5, 32'h4122c306} /* (6, 20, 30) {real, imag} */,
  {32'h4099b50c, 32'hbf47db20} /* (6, 20, 29) {real, imag} */,
  {32'h400d8269, 32'hbfa93dcb} /* (6, 20, 28) {real, imag} */,
  {32'hbfa4b3f8, 32'hbd2780c0} /* (6, 20, 27) {real, imag} */,
  {32'hc0a55228, 32'h40147cbc} /* (6, 20, 26) {real, imag} */,
  {32'hc0ff89f3, 32'hc085d484} /* (6, 20, 25) {real, imag} */,
  {32'hc13422e4, 32'hc0550b5c} /* (6, 20, 24) {real, imag} */,
  {32'hc0340c6e, 32'hbf51841c} /* (6, 20, 23) {real, imag} */,
  {32'h3f1b8b38, 32'hc05d6518} /* (6, 20, 22) {real, imag} */,
  {32'hbfe6b13c, 32'hbeade120} /* (6, 20, 21) {real, imag} */,
  {32'h408cca17, 32'hc0289da3} /* (6, 20, 20) {real, imag} */,
  {32'h4127efe7, 32'hbf48ea58} /* (6, 20, 19) {real, imag} */,
  {32'hbf2195d8, 32'h40c2c334} /* (6, 20, 18) {real, imag} */,
  {32'hbed88938, 32'hc05c46cc} /* (6, 20, 17) {real, imag} */,
  {32'h40606935, 32'h40359512} /* (6, 20, 16) {real, imag} */,
  {32'h411f93a2, 32'h41231352} /* (6, 20, 15) {real, imag} */,
  {32'h40bfab77, 32'h406a2550} /* (6, 20, 14) {real, imag} */,
  {32'hc0063ea5, 32'hbffdb7ea} /* (6, 20, 13) {real, imag} */,
  {32'hc00785be, 32'h3f5435b0} /* (6, 20, 12) {real, imag} */,
  {32'hc0442258, 32'h408931ca} /* (6, 20, 11) {real, imag} */,
  {32'hc029cc9f, 32'h4043df0b} /* (6, 20, 10) {real, imag} */,
  {32'hbfc53cfe, 32'h3f9c2c9e} /* (6, 20, 9) {real, imag} */,
  {32'h405c995f, 32'h3fac337e} /* (6, 20, 8) {real, imag} */,
  {32'h404924e4, 32'h405de26e} /* (6, 20, 7) {real, imag} */,
  {32'h4015632f, 32'h3f458f04} /* (6, 20, 6) {real, imag} */,
  {32'h3faf17bc, 32'h3fb41a6a} /* (6, 20, 5) {real, imag} */,
  {32'h3e773aa0, 32'h40365390} /* (6, 20, 4) {real, imag} */,
  {32'h408b2edc, 32'hbfbece8c} /* (6, 20, 3) {real, imag} */,
  {32'h3f778700, 32'h3fee7f52} /* (6, 20, 2) {real, imag} */,
  {32'hc063a444, 32'hbfcb9fbc} /* (6, 20, 1) {real, imag} */,
  {32'h3e082860, 32'h400378f8} /* (6, 20, 0) {real, imag} */,
  {32'hc0087642, 32'hc0091b7e} /* (6, 19, 31) {real, imag} */,
  {32'hbfa3a790, 32'hbfe7f348} /* (6, 19, 30) {real, imag} */,
  {32'h402c8080, 32'h40852c2a} /* (6, 19, 29) {real, imag} */,
  {32'h400a9a8e, 32'h3f067b78} /* (6, 19, 28) {real, imag} */,
  {32'hc0874711, 32'h3ecd48f8} /* (6, 19, 27) {real, imag} */,
  {32'h40113fc8, 32'h40130db8} /* (6, 19, 26) {real, imag} */,
  {32'h3d423a40, 32'hc084d7f4} /* (6, 19, 25) {real, imag} */,
  {32'hc0488a75, 32'hc0acbeac} /* (6, 19, 24) {real, imag} */,
  {32'hc0a29a4f, 32'h3e399160} /* (6, 19, 23) {real, imag} */,
  {32'hc0f1fd00, 32'hbfc468b6} /* (6, 19, 22) {real, imag} */,
  {32'hc0be6230, 32'h3b3d5a00} /* (6, 19, 21) {real, imag} */,
  {32'h3eda9f34, 32'h3fa61f48} /* (6, 19, 20) {real, imag} */,
  {32'h3e8d42c0, 32'h3f21f8aa} /* (6, 19, 19) {real, imag} */,
  {32'hc06d1bcb, 32'hc094df95} /* (6, 19, 18) {real, imag} */,
  {32'h3f8d90d8, 32'hc0da607a} /* (6, 19, 17) {real, imag} */,
  {32'h403c2664, 32'hc04521a4} /* (6, 19, 16) {real, imag} */,
  {32'h405392d2, 32'hbfc3252e} /* (6, 19, 15) {real, imag} */,
  {32'h409c2f93, 32'hc078f8bc} /* (6, 19, 14) {real, imag} */,
  {32'h4073bc97, 32'hc0ce5d64} /* (6, 19, 13) {real, imag} */,
  {32'h40d18571, 32'hbf93e764} /* (6, 19, 12) {real, imag} */,
  {32'h402ce291, 32'h3fccbf98} /* (6, 19, 11) {real, imag} */,
  {32'hbf8f245e, 32'h3ecd7d78} /* (6, 19, 10) {real, imag} */,
  {32'hc08119da, 32'hc04055e0} /* (6, 19, 9) {real, imag} */,
  {32'h400e4aeb, 32'hbf7c5996} /* (6, 19, 8) {real, imag} */,
  {32'h40be035a, 32'hbf4414e0} /* (6, 19, 7) {real, imag} */,
  {32'hc056cee4, 32'hbfcc15c0} /* (6, 19, 6) {real, imag} */,
  {32'hc02c82d6, 32'h3ec5f1f0} /* (6, 19, 5) {real, imag} */,
  {32'h3e358d38, 32'h4091466e} /* (6, 19, 4) {real, imag} */,
  {32'h400be6fc, 32'hbfdfaedc} /* (6, 19, 3) {real, imag} */,
  {32'hbf0c2d34, 32'h4055362e} /* (6, 19, 2) {real, imag} */,
  {32'hc02105c2, 32'h407f68e8} /* (6, 19, 1) {real, imag} */,
  {32'hc087513e, 32'hc00f9fad} /* (6, 19, 0) {real, imag} */,
  {32'h3f78d6c2, 32'hbfa5d448} /* (6, 18, 31) {real, imag} */,
  {32'hc0a2b49c, 32'hc03a686e} /* (6, 18, 30) {real, imag} */,
  {32'hc09ceafd, 32'h3e323eb8} /* (6, 18, 29) {real, imag} */,
  {32'hbfe0f83d, 32'h4042939c} /* (6, 18, 28) {real, imag} */,
  {32'h40700129, 32'hc0823bfd} /* (6, 18, 27) {real, imag} */,
  {32'h3f73ef70, 32'hc09216fe} /* (6, 18, 26) {real, imag} */,
  {32'h3fdbe9a4, 32'hc03521ce} /* (6, 18, 25) {real, imag} */,
  {32'h40846766, 32'hbffd9855} /* (6, 18, 24) {real, imag} */,
  {32'h404c9b56, 32'h3f5890a8} /* (6, 18, 23) {real, imag} */,
  {32'h40623f2a, 32'hc0267f54} /* (6, 18, 22) {real, imag} */,
  {32'h4050fe30, 32'hc06e7bcc} /* (6, 18, 21) {real, imag} */,
  {32'h40998fb2, 32'hc0bc31c8} /* (6, 18, 20) {real, imag} */,
  {32'h3ff279b6, 32'hbe2efb80} /* (6, 18, 19) {real, imag} */,
  {32'hbfb0cb0c, 32'h3f16fb1c} /* (6, 18, 18) {real, imag} */,
  {32'hc0bff288, 32'hbffeaba4} /* (6, 18, 17) {real, imag} */,
  {32'hc076a5cc, 32'h3e5a8e60} /* (6, 18, 16) {real, imag} */,
  {32'h3f872b5c, 32'h3f70e108} /* (6, 18, 15) {real, imag} */,
  {32'h4017c486, 32'hbeff7990} /* (6, 18, 14) {real, imag} */,
  {32'h409ffb0b, 32'hc0098020} /* (6, 18, 13) {real, imag} */,
  {32'h40bacfc2, 32'h405cee25} /* (6, 18, 12) {real, imag} */,
  {32'h3fa865f0, 32'hbfb82c90} /* (6, 18, 11) {real, imag} */,
  {32'h4005d51c, 32'hc02ab9f9} /* (6, 18, 10) {real, imag} */,
  {32'h3e24bcf0, 32'h3f0f3c08} /* (6, 18, 9) {real, imag} */,
  {32'hc0f8acec, 32'h3fa5ef4e} /* (6, 18, 8) {real, imag} */,
  {32'hc1345e90, 32'h408c9ed4} /* (6, 18, 7) {real, imag} */,
  {32'hc09fd25c, 32'h40906e7c} /* (6, 18, 6) {real, imag} */,
  {32'h40048064, 32'h3f1fdc50} /* (6, 18, 5) {real, imag} */,
  {32'h4046aec2, 32'hbfabe0a4} /* (6, 18, 4) {real, imag} */,
  {32'h40560768, 32'hc0312f0b} /* (6, 18, 3) {real, imag} */,
  {32'h3fc367f6, 32'hbff41b66} /* (6, 18, 2) {real, imag} */,
  {32'hc0309372, 32'h4090d05d} /* (6, 18, 1) {real, imag} */,
  {32'hc0812158, 32'h408dcc7a} /* (6, 18, 0) {real, imag} */,
  {32'hc04505b9, 32'h408cf9d6} /* (6, 17, 31) {real, imag} */,
  {32'h400159b2, 32'h3fe5bb6f} /* (6, 17, 30) {real, imag} */,
  {32'h3f8af4da, 32'h3fda012e} /* (6, 17, 29) {real, imag} */,
  {32'hc05fdf71, 32'h40b0aeaf} /* (6, 17, 28) {real, imag} */,
  {32'hc08c0a54, 32'h40944cca} /* (6, 17, 27) {real, imag} */,
  {32'hc00420c0, 32'h402fa39d} /* (6, 17, 26) {real, imag} */,
  {32'h3e51e400, 32'hbfbadd26} /* (6, 17, 25) {real, imag} */,
  {32'hbe968d34, 32'h3fb253ef} /* (6, 17, 24) {real, imag} */,
  {32'hbf99f308, 32'h3f652222} /* (6, 17, 23) {real, imag} */,
  {32'hc06a901e, 32'hc02fb6a5} /* (6, 17, 22) {real, imag} */,
  {32'h4080fc16, 32'hc08e2d65} /* (6, 17, 21) {real, imag} */,
  {32'hc00e91e8, 32'hc1029d14} /* (6, 17, 20) {real, imag} */,
  {32'hbe5e6fd0, 32'hc0c7e191} /* (6, 17, 19) {real, imag} */,
  {32'h3f832fc6, 32'h400d418d} /* (6, 17, 18) {real, imag} */,
  {32'h3f169058, 32'h3eece300} /* (6, 17, 17) {real, imag} */,
  {32'hc050b9cf, 32'h3ee40e50} /* (6, 17, 16) {real, imag} */,
  {32'hc058768e, 32'hbdc52440} /* (6, 17, 15) {real, imag} */,
  {32'hc0484796, 32'h403f3182} /* (6, 17, 14) {real, imag} */,
  {32'hc07efbee, 32'h40371dca} /* (6, 17, 13) {real, imag} */,
  {32'hc0a9f664, 32'h409edb83} /* (6, 17, 12) {real, imag} */,
  {32'hbf59fc54, 32'h409e9c3c} /* (6, 17, 11) {real, imag} */,
  {32'h3ec81048, 32'h4039477a} /* (6, 17, 10) {real, imag} */,
  {32'h404399fa, 32'h403e592a} /* (6, 17, 9) {real, imag} */,
  {32'h401e7d8a, 32'hc051a8a4} /* (6, 17, 8) {real, imag} */,
  {32'hbe7c9020, 32'hc0eae460} /* (6, 17, 7) {real, imag} */,
  {32'hc0be8800, 32'hc1169a8c} /* (6, 17, 6) {real, imag} */,
  {32'hbf39315c, 32'hc101f266} /* (6, 17, 5) {real, imag} */,
  {32'h3fa9358a, 32'hc0c6e7e0} /* (6, 17, 4) {real, imag} */,
  {32'hbda88618, 32'hbf201214} /* (6, 17, 3) {real, imag} */,
  {32'hbf4cd41c, 32'h3fc9809e} /* (6, 17, 2) {real, imag} */,
  {32'hbf67744e, 32'h3ffa0274} /* (6, 17, 1) {real, imag} */,
  {32'hc0ac2a17, 32'h402183d3} /* (6, 17, 0) {real, imag} */,
  {32'hbf8b1097, 32'h4048120a} /* (6, 16, 31) {real, imag} */,
  {32'h406256c2, 32'h3dd17380} /* (6, 16, 30) {real, imag} */,
  {32'h401562ca, 32'h3fcd0f74} /* (6, 16, 29) {real, imag} */,
  {32'h3ff68010, 32'hbf57c750} /* (6, 16, 28) {real, imag} */,
  {32'hbd35b800, 32'h3cf70600} /* (6, 16, 27) {real, imag} */,
  {32'hc05b82c4, 32'h3d0ddb60} /* (6, 16, 26) {real, imag} */,
  {32'hc081def7, 32'hbfe023c5} /* (6, 16, 25) {real, imag} */,
  {32'h3f19c778, 32'h3e5d1bd0} /* (6, 16, 24) {real, imag} */,
  {32'h4066d5a6, 32'hbeba8770} /* (6, 16, 23) {real, imag} */,
  {32'h3d19fe60, 32'hbf7047e0} /* (6, 16, 22) {real, imag} */,
  {32'hbf79211c, 32'h4040806e} /* (6, 16, 21) {real, imag} */,
  {32'hbd142540, 32'h3e6661a0} /* (6, 16, 20) {real, imag} */,
  {32'hbf6338c4, 32'h3ed202a0} /* (6, 16, 19) {real, imag} */,
  {32'h3f4281fd, 32'h40073d64} /* (6, 16, 18) {real, imag} */,
  {32'h3f371d90, 32'h4031e2a7} /* (6, 16, 17) {real, imag} */,
  {32'hbfc9f872, 32'h3e812fac} /* (6, 16, 16) {real, imag} */,
  {32'hc03b2f72, 32'h408ef44a} /* (6, 16, 15) {real, imag} */,
  {32'hbfc818b8, 32'h401bf9c4} /* (6, 16, 14) {real, imag} */,
  {32'h405789c0, 32'h3ff63d5a} /* (6, 16, 13) {real, imag} */,
  {32'h40944284, 32'h3f2ff2e0} /* (6, 16, 12) {real, imag} */,
  {32'h4076490e, 32'h3f9b1910} /* (6, 16, 11) {real, imag} */,
  {32'h3fcc7a9c, 32'h3e6f1c60} /* (6, 16, 10) {real, imag} */,
  {32'hc008a576, 32'hc0786ab8} /* (6, 16, 9) {real, imag} */,
  {32'hc07a3450, 32'h3e71ec00} /* (6, 16, 8) {real, imag} */,
  {32'hbf9eea10, 32'hbf37fd78} /* (6, 16, 7) {real, imag} */,
  {32'hc01a4efa, 32'h3f79c0c0} /* (6, 16, 6) {real, imag} */,
  {32'h3f9e1557, 32'hbfc1a828} /* (6, 16, 5) {real, imag} */,
  {32'h4014b88c, 32'hc03cf568} /* (6, 16, 4) {real, imag} */,
  {32'h405e15e3, 32'hbf6b6c30} /* (6, 16, 3) {real, imag} */,
  {32'h3fe21216, 32'hbf5d5240} /* (6, 16, 2) {real, imag} */,
  {32'hbf8952d8, 32'hbfeabc80} /* (6, 16, 1) {real, imag} */,
  {32'h3f9d4050, 32'hbf782f18} /* (6, 16, 0) {real, imag} */,
  {32'h40d863ca, 32'hbfa2eac0} /* (6, 15, 31) {real, imag} */,
  {32'h40927667, 32'h4032d704} /* (6, 15, 30) {real, imag} */,
  {32'h3e968a38, 32'h3f18de6b} /* (6, 15, 29) {real, imag} */,
  {32'h40884a7a, 32'hc01ba7ce} /* (6, 15, 28) {real, imag} */,
  {32'h40009c80, 32'hbf0b55fc} /* (6, 15, 27) {real, imag} */,
  {32'hbfd46ce0, 32'h404d6c8d} /* (6, 15, 26) {real, imag} */,
  {32'hc065ce60, 32'h40748e69} /* (6, 15, 25) {real, imag} */,
  {32'hbff56a4d, 32'h3fd1dd45} /* (6, 15, 24) {real, imag} */,
  {32'h3f8f256c, 32'h3e3610f8} /* (6, 15, 23) {real, imag} */,
  {32'h410b9856, 32'h409c03e8} /* (6, 15, 22) {real, imag} */,
  {32'h4060f088, 32'h406c234e} /* (6, 15, 21) {real, imag} */,
  {32'h400873a8, 32'hbeb5d180} /* (6, 15, 20) {real, imag} */,
  {32'h409b470c, 32'hc0d7c0fb} /* (6, 15, 19) {real, imag} */,
  {32'h40793c05, 32'hc04ad3b3} /* (6, 15, 18) {real, imag} */,
  {32'h3f32fa08, 32'h40cca910} /* (6, 15, 17) {real, imag} */,
  {32'h3e87e248, 32'h410d7b50} /* (6, 15, 16) {real, imag} */,
  {32'hbfae06f4, 32'h41002488} /* (6, 15, 15) {real, imag} */,
  {32'hbf7e1a88, 32'h40b3dea7} /* (6, 15, 14) {real, imag} */,
  {32'h40164426, 32'h3f590266} /* (6, 15, 13) {real, imag} */,
  {32'hbe848148, 32'hc052888a} /* (6, 15, 12) {real, imag} */,
  {32'h3f458894, 32'hc031d568} /* (6, 15, 11) {real, imag} */,
  {32'h40da9fe6, 32'h404213ac} /* (6, 15, 10) {real, imag} */,
  {32'h402e2eba, 32'hc035a472} /* (6, 15, 9) {real, imag} */,
  {32'hbfd1634c, 32'hc07c7310} /* (6, 15, 8) {real, imag} */,
  {32'hbfb8e8b4, 32'h3dc51e20} /* (6, 15, 7) {real, imag} */,
  {32'h40357d70, 32'h3d7b2200} /* (6, 15, 6) {real, imag} */,
  {32'h3fdfd2e6, 32'hc030937c} /* (6, 15, 5) {real, imag} */,
  {32'hc003a079, 32'hc057e45c} /* (6, 15, 4) {real, imag} */,
  {32'h3f84df68, 32'h400677d9} /* (6, 15, 3) {real, imag} */,
  {32'h4075d6b3, 32'h3eefede8} /* (6, 15, 2) {real, imag} */,
  {32'h3fa34d33, 32'hbf9ecdcc} /* (6, 15, 1) {real, imag} */,
  {32'h3e75e5e0, 32'hc012426d} /* (6, 15, 0) {real, imag} */,
  {32'h3d8fb830, 32'h3f6cc6d0} /* (6, 14, 31) {real, imag} */,
  {32'hc084a5a0, 32'hbfd11a94} /* (6, 14, 30) {real, imag} */,
  {32'hc06792fa, 32'hc0849995} /* (6, 14, 29) {real, imag} */,
  {32'hc022a9f2, 32'hc08a04f0} /* (6, 14, 28) {real, imag} */,
  {32'hc07e1fe9, 32'hc0412cca} /* (6, 14, 27) {real, imag} */,
  {32'hc0778bd0, 32'h406a99f4} /* (6, 14, 26) {real, imag} */,
  {32'hc02a1e3e, 32'h3e152c58} /* (6, 14, 25) {real, imag} */,
  {32'h3f2701e4, 32'hc0374616} /* (6, 14, 24) {real, imag} */,
  {32'h3f049280, 32'hc03a267a} /* (6, 14, 23) {real, imag} */,
  {32'hbf88849d, 32'hc039b83a} /* (6, 14, 22) {real, imag} */,
  {32'hc02fd4bc, 32'h404c7814} /* (6, 14, 21) {real, imag} */,
  {32'hc0023ab8, 32'h40d17ba4} /* (6, 14, 20) {real, imag} */,
  {32'h4048a1a3, 32'h3f901d50} /* (6, 14, 19) {real, imag} */,
  {32'h4100f92e, 32'hc009d613} /* (6, 14, 18) {real, imag} */,
  {32'h3ed32b38, 32'h403dfa1c} /* (6, 14, 17) {real, imag} */,
  {32'hc0402c98, 32'h4097716d} /* (6, 14, 16) {real, imag} */,
  {32'h3e283a20, 32'h40a49ee7} /* (6, 14, 15) {real, imag} */,
  {32'h3ef11f90, 32'h40be0b45} /* (6, 14, 14) {real, imag} */,
  {32'h3f579d28, 32'h400f50d4} /* (6, 14, 13) {real, imag} */,
  {32'hbe143f70, 32'h400b06ad} /* (6, 14, 12) {real, imag} */,
  {32'h3fcb33a0, 32'hbea06150} /* (6, 14, 11) {real, imag} */,
  {32'hc00c6d0c, 32'h3ef60548} /* (6, 14, 10) {real, imag} */,
  {32'hc081adcc, 32'hbf0e0158} /* (6, 14, 9) {real, imag} */,
  {32'hc0e99b0a, 32'h3ee533f8} /* (6, 14, 8) {real, imag} */,
  {32'h3fa34674, 32'hbf1cb564} /* (6, 14, 7) {real, imag} */,
  {32'hbe9ea9d0, 32'h409f4a32} /* (6, 14, 6) {real, imag} */,
  {32'hc0ca566e, 32'h409ed998} /* (6, 14, 5) {real, imag} */,
  {32'hc00da226, 32'h3f70bce0} /* (6, 14, 4) {real, imag} */,
  {32'h3e4ff6a8, 32'hbe8efc88} /* (6, 14, 3) {real, imag} */,
  {32'h3f62fb84, 32'hbc8cd2a0} /* (6, 14, 2) {real, imag} */,
  {32'hc094b83f, 32'h40d2b709} /* (6, 14, 1) {real, imag} */,
  {32'hc0a8aef4, 32'h40ec117a} /* (6, 14, 0) {real, imag} */,
  {32'h4014c492, 32'hbf3047d6} /* (6, 13, 31) {real, imag} */,
  {32'h406713bc, 32'h3f978e28} /* (6, 13, 30) {real, imag} */,
  {32'h3fa49bf7, 32'h4008260c} /* (6, 13, 29) {real, imag} */,
  {32'hbf8eaee4, 32'h3fbbf568} /* (6, 13, 28) {real, imag} */,
  {32'hc0404ba8, 32'hc0256c43} /* (6, 13, 27) {real, imag} */,
  {32'hc00d5f80, 32'hbe460200} /* (6, 13, 26) {real, imag} */,
  {32'h40aaff0c, 32'h3e90db60} /* (6, 13, 25) {real, imag} */,
  {32'h40cd08ee, 32'hc0c18b58} /* (6, 13, 24) {real, imag} */,
  {32'h3fd21f64, 32'h408ff67d} /* (6, 13, 23) {real, imag} */,
  {32'hbfde9e58, 32'hc019e676} /* (6, 13, 22) {real, imag} */,
  {32'hbe9cf4c0, 32'hbe722d18} /* (6, 13, 21) {real, imag} */,
  {32'h3fd480dd, 32'h403ed458} /* (6, 13, 20) {real, imag} */,
  {32'hc0559dc0, 32'h3e742508} /* (6, 13, 19) {real, imag} */,
  {32'hc0411f2d, 32'h40f1791d} /* (6, 13, 18) {real, imag} */,
  {32'hc0c1a548, 32'h410f6d47} /* (6, 13, 17) {real, imag} */,
  {32'hbf850268, 32'h410fc8a7} /* (6, 13, 16) {real, imag} */,
  {32'h3ff1b6cc, 32'hbfed0daa} /* (6, 13, 15) {real, imag} */,
  {32'hc01cad28, 32'hc0d96b70} /* (6, 13, 14) {real, imag} */,
  {32'hc07d3f1f, 32'hbfe674b8} /* (6, 13, 13) {real, imag} */,
  {32'hc0ce1a7b, 32'h4089cb79} /* (6, 13, 12) {real, imag} */,
  {32'hbfde463e, 32'h4090d042} /* (6, 13, 11) {real, imag} */,
  {32'hc03d5c11, 32'h3f1d9094} /* (6, 13, 10) {real, imag} */,
  {32'h4082d646, 32'h3fe46d80} /* (6, 13, 9) {real, imag} */,
  {32'h3fd90c9a, 32'hc03b0216} /* (6, 13, 8) {real, imag} */,
  {32'h4065b9b8, 32'hc01fdbb8} /* (6, 13, 7) {real, imag} */,
  {32'h3f8b4a04, 32'hc0b49b1a} /* (6, 13, 6) {real, imag} */,
  {32'hc0506412, 32'hc0923f5d} /* (6, 13, 5) {real, imag} */,
  {32'h403e6f98, 32'hc0a2aa1c} /* (6, 13, 4) {real, imag} */,
  {32'h4075eda6, 32'hc04a3ebe} /* (6, 13, 3) {real, imag} */,
  {32'h3ff0df0a, 32'hc0c4d681} /* (6, 13, 2) {real, imag} */,
  {32'hc03b7162, 32'hc107e292} /* (6, 13, 1) {real, imag} */,
  {32'hbf9b57e7, 32'hc0c90552} /* (6, 13, 0) {real, imag} */,
  {32'hc1083c03, 32'h3f813ca0} /* (6, 12, 31) {real, imag} */,
  {32'hc0cef22e, 32'hc0066ab4} /* (6, 12, 30) {real, imag} */,
  {32'hc07c1cdc, 32'hc0eede8c} /* (6, 12, 29) {real, imag} */,
  {32'hc01f5843, 32'hc094cf15} /* (6, 12, 28) {real, imag} */,
  {32'h3f9c9770, 32'h3f36b194} /* (6, 12, 27) {real, imag} */,
  {32'h409333b0, 32'hc02d79e8} /* (6, 12, 26) {real, imag} */,
  {32'h403ddc0e, 32'hc0491b0b} /* (6, 12, 25) {real, imag} */,
  {32'hc03f63aa, 32'h405910fe} /* (6, 12, 24) {real, imag} */,
  {32'hc013ff3e, 32'h408a01f0} /* (6, 12, 23) {real, imag} */,
  {32'hc0c95d21, 32'h4025c470} /* (6, 12, 22) {real, imag} */,
  {32'hc0a57f47, 32'h40523a9c} /* (6, 12, 21) {real, imag} */,
  {32'h40bccdc1, 32'h3ec5d4c8} /* (6, 12, 20) {real, imag} */,
  {32'h407f4a88, 32'h404450a2} /* (6, 12, 19) {real, imag} */,
  {32'hbf872f6c, 32'h40936128} /* (6, 12, 18) {real, imag} */,
  {32'hbfec448e, 32'hc09ca4b2} /* (6, 12, 17) {real, imag} */,
  {32'hc0938746, 32'hc0da526b} /* (6, 12, 16) {real, imag} */,
  {32'hbf912a50, 32'h3fdf3e1c} /* (6, 12, 15) {real, imag} */,
  {32'h403e126e, 32'h40466dc2} /* (6, 12, 14) {real, imag} */,
  {32'h408f6d7e, 32'h3f83183a} /* (6, 12, 13) {real, imag} */,
  {32'h3f5fc936, 32'hc0c92c38} /* (6, 12, 12) {real, imag} */,
  {32'h402bd7a0, 32'hc11180ea} /* (6, 12, 11) {real, imag} */,
  {32'h40addc5a, 32'hc0b1b322} /* (6, 12, 10) {real, imag} */,
  {32'hbfe70a52, 32'h40332021} /* (6, 12, 9) {real, imag} */,
  {32'h3eb9e818, 32'h4012373d} /* (6, 12, 8) {real, imag} */,
  {32'h405dc664, 32'h3f180f78} /* (6, 12, 7) {real, imag} */,
  {32'hc056926d, 32'h3da4d1e0} /* (6, 12, 6) {real, imag} */,
  {32'hbf80c494, 32'h401099bf} /* (6, 12, 5) {real, imag} */,
  {32'hc05a699e, 32'h405869d8} /* (6, 12, 4) {real, imag} */,
  {32'hc01ba3e8, 32'h3fbe4f5c} /* (6, 12, 3) {real, imag} */,
  {32'hc10f34de, 32'h3f2edd9b} /* (6, 12, 2) {real, imag} */,
  {32'hc0a8fa16, 32'hc0a455fb} /* (6, 12, 1) {real, imag} */,
  {32'hbf77ed88, 32'h3f81c8c0} /* (6, 12, 0) {real, imag} */,
  {32'h4094a284, 32'hc0842ca2} /* (6, 11, 31) {real, imag} */,
  {32'h410fb384, 32'hc023b1e7} /* (6, 11, 30) {real, imag} */,
  {32'h41295d6a, 32'hc0c58f2a} /* (6, 11, 29) {real, imag} */,
  {32'h407ff1f8, 32'h3db0ebd0} /* (6, 11, 28) {real, imag} */,
  {32'hc0179184, 32'h40c19ae0} /* (6, 11, 27) {real, imag} */,
  {32'h401b122b, 32'hbff011f2} /* (6, 11, 26) {real, imag} */,
  {32'h41310ad6, 32'h3f87f57a} /* (6, 11, 25) {real, imag} */,
  {32'h404e3266, 32'h4118383c} /* (6, 11, 24) {real, imag} */,
  {32'hc05367f5, 32'h3eb32370} /* (6, 11, 23) {real, imag} */,
  {32'h3d85a740, 32'h4078a4fb} /* (6, 11, 22) {real, imag} */,
  {32'h408f1410, 32'h4083d285} /* (6, 11, 21) {real, imag} */,
  {32'h4052212b, 32'h40b2c9f1} /* (6, 11, 20) {real, imag} */,
  {32'h402e4386, 32'h4054dfe7} /* (6, 11, 19) {real, imag} */,
  {32'hc0f6e272, 32'h4098025c} /* (6, 11, 18) {real, imag} */,
  {32'hbf0ed96c, 32'hbfde5aea} /* (6, 11, 17) {real, imag} */,
  {32'h4109719e, 32'h40c4ef7a} /* (6, 11, 16) {real, imag} */,
  {32'h410e5958, 32'h40d23842} /* (6, 11, 15) {real, imag} */,
  {32'h402a0706, 32'h411028f6} /* (6, 11, 14) {real, imag} */,
  {32'hc05f8384, 32'hbe7f51b4} /* (6, 11, 13) {real, imag} */,
  {32'h4047b0fe, 32'hc0030abc} /* (6, 11, 12) {real, imag} */,
  {32'h4114b344, 32'hc092b708} /* (6, 11, 11) {real, imag} */,
  {32'h40cfca6e, 32'hc0f92898} /* (6, 11, 10) {real, imag} */,
  {32'hc0a93215, 32'h405b4fe0} /* (6, 11, 9) {real, imag} */,
  {32'hc14328e5, 32'h4101beb6} /* (6, 11, 8) {real, imag} */,
  {32'hc1531694, 32'h40e5eb8c} /* (6, 11, 7) {real, imag} */,
  {32'hc11cc4ac, 32'hbf342520} /* (6, 11, 6) {real, imag} */,
  {32'hbdc72900, 32'hbf809ae8} /* (6, 11, 5) {real, imag} */,
  {32'h404e1e5a, 32'h3ea3c530} /* (6, 11, 4) {real, imag} */,
  {32'hbf7b4b94, 32'h4088c4b6} /* (6, 11, 3) {real, imag} */,
  {32'h40490fc4, 32'h3ff0f642} /* (6, 11, 2) {real, imag} */,
  {32'hbf289e9e, 32'hc01bd9d3} /* (6, 11, 1) {real, imag} */,
  {32'h3e9cb5e0, 32'hbf2417dc} /* (6, 11, 0) {real, imag} */,
  {32'h3ff4025a, 32'hc062c7e4} /* (6, 10, 31) {real, imag} */,
  {32'h3f71b21e, 32'hc122b6aa} /* (6, 10, 30) {real, imag} */,
  {32'h3d01e900, 32'hc0892f40} /* (6, 10, 29) {real, imag} */,
  {32'hbfe9005e, 32'h40f09a5a} /* (6, 10, 28) {real, imag} */,
  {32'hbfe1149c, 32'h4030de8b} /* (6, 10, 27) {real, imag} */,
  {32'h40e0572d, 32'hbefff810} /* (6, 10, 26) {real, imag} */,
  {32'h3fba73c4, 32'hbf04a0d6} /* (6, 10, 25) {real, imag} */,
  {32'hc08480bb, 32'hc11162f4} /* (6, 10, 24) {real, imag} */,
  {32'hc087c4ec, 32'h3f9ead4e} /* (6, 10, 23) {real, imag} */,
  {32'h40e1604e, 32'hc071e5ce} /* (6, 10, 22) {real, imag} */,
  {32'hc03aeabc, 32'hc101035c} /* (6, 10, 21) {real, imag} */,
  {32'h40fb1c52, 32'hc04daf60} /* (6, 10, 20) {real, imag} */,
  {32'h40082dcc, 32'hc0ff4134} /* (6, 10, 19) {real, imag} */,
  {32'hc1441bed, 32'hc086cd02} /* (6, 10, 18) {real, imag} */,
  {32'hc01f7d33, 32'hc040d176} /* (6, 10, 17) {real, imag} */,
  {32'h4120948c, 32'hc0e4d432} /* (6, 10, 16) {real, imag} */,
  {32'h415fa858, 32'hc0f6b610} /* (6, 10, 15) {real, imag} */,
  {32'h40c038ea, 32'hc0fa9f66} /* (6, 10, 14) {real, imag} */,
  {32'hc05ad7f6, 32'h3fb99658} /* (6, 10, 13) {real, imag} */,
  {32'hc100531c, 32'hbe0e4a60} /* (6, 10, 12) {real, imag} */,
  {32'hc0428b31, 32'h40024389} /* (6, 10, 11) {real, imag} */,
  {32'hc0972c24, 32'h4033ae79} /* (6, 10, 10) {real, imag} */,
  {32'hc04fd4df, 32'h3fca6422} /* (6, 10, 9) {real, imag} */,
  {32'h40f2f3aa, 32'hc0d4c8bc} /* (6, 10, 8) {real, imag} */,
  {32'h415ef1d2, 32'hc0e80591} /* (6, 10, 7) {real, imag} */,
  {32'hc02d1ec1, 32'hbecc31d0} /* (6, 10, 6) {real, imag} */,
  {32'hc0068be2, 32'hc08e7d92} /* (6, 10, 5) {real, imag} */,
  {32'h404d67d1, 32'hbe6ffe80} /* (6, 10, 4) {real, imag} */,
  {32'hbfb4b34e, 32'h403a8dc9} /* (6, 10, 3) {real, imag} */,
  {32'h3fe5f61e, 32'h413a31ee} /* (6, 10, 2) {real, imag} */,
  {32'hbf65fbd8, 32'h4108e05e} /* (6, 10, 1) {real, imag} */,
  {32'hc0237bad, 32'h40c00fc9} /* (6, 10, 0) {real, imag} */,
  {32'hc05faf75, 32'h3fbcd916} /* (6, 9, 31) {real, imag} */,
  {32'hc107b7e6, 32'h3fac2ffc} /* (6, 9, 30) {real, imag} */,
  {32'h3ef1ac60, 32'hc0c99cb6} /* (6, 9, 29) {real, imag} */,
  {32'h41495db8, 32'hc0bc3a05} /* (6, 9, 28) {real, imag} */,
  {32'h3e958680, 32'h3fd66dac} /* (6, 9, 27) {real, imag} */,
  {32'hc09c5f1c, 32'h4102ee92} /* (6, 9, 26) {real, imag} */,
  {32'hbf2c1210, 32'h40fa0d26} /* (6, 9, 25) {real, imag} */,
  {32'h3fa917b8, 32'h418bb278} /* (6, 9, 24) {real, imag} */,
  {32'hc13a392d, 32'h418b7348} /* (6, 9, 23) {real, imag} */,
  {32'hc15999e4, 32'h415c0a8a} /* (6, 9, 22) {real, imag} */,
  {32'hc0d931d4, 32'h408aeaa5} /* (6, 9, 21) {real, imag} */,
  {32'h3f792508, 32'h41031c38} /* (6, 9, 20) {real, imag} */,
  {32'h41023b0c, 32'h40ca9470} /* (6, 9, 19) {real, imag} */,
  {32'hbf1d8f20, 32'hc0c0e2fb} /* (6, 9, 18) {real, imag} */,
  {32'hbf710a48, 32'hc0d5c144} /* (6, 9, 17) {real, imag} */,
  {32'hc0b0f0d5, 32'hc0a59c63} /* (6, 9, 16) {real, imag} */,
  {32'h41019b44, 32'h4025708a} /* (6, 9, 15) {real, imag} */,
  {32'h4173174c, 32'h40789105} /* (6, 9, 14) {real, imag} */,
  {32'hbe4a25e8, 32'h40f04fef} /* (6, 9, 13) {real, imag} */,
  {32'h40840cff, 32'h41180784} /* (6, 9, 12) {real, imag} */,
  {32'h413688f2, 32'h4182fb08} /* (6, 9, 11) {real, imag} */,
  {32'h3fe15288, 32'h409da81f} /* (6, 9, 10) {real, imag} */,
  {32'hc04349da, 32'hc0564863} /* (6, 9, 9) {real, imag} */,
  {32'hc091209e, 32'h3ff8516a} /* (6, 9, 8) {real, imag} */,
  {32'hc0be1580, 32'hbf07b7ec} /* (6, 9, 7) {real, imag} */,
  {32'hc085e746, 32'h4141fa5c} /* (6, 9, 6) {real, imag} */,
  {32'h408b3b18, 32'h4172c845} /* (6, 9, 5) {real, imag} */,
  {32'hbd750140, 32'h415c9497} /* (6, 9, 4) {real, imag} */,
  {32'hc126f7bc, 32'h411f48f6} /* (6, 9, 3) {real, imag} */,
  {32'hc0bcd8a0, 32'h40e57b88} /* (6, 9, 2) {real, imag} */,
  {32'h403b2232, 32'h4185ac12} /* (6, 9, 1) {real, imag} */,
  {32'h41370c6a, 32'h411a627a} /* (6, 9, 0) {real, imag} */,
  {32'hc0bae6c6, 32'h404728be} /* (6, 8, 31) {real, imag} */,
  {32'hc01df2b3, 32'h409d1147} /* (6, 8, 30) {real, imag} */,
  {32'h412c3616, 32'h40c1d3ec} /* (6, 8, 29) {real, imag} */,
  {32'h4175c84f, 32'h415e39ad} /* (6, 8, 28) {real, imag} */,
  {32'h4069c675, 32'h41264735} /* (6, 8, 27) {real, imag} */,
  {32'hc1045ef8, 32'hbfcece14} /* (6, 8, 26) {real, imag} */,
  {32'hc0b1c018, 32'h3eac18a0} /* (6, 8, 25) {real, imag} */,
  {32'h4156bbd6, 32'hc1000363} /* (6, 8, 24) {real, imag} */,
  {32'hc09d3cea, 32'hc02243db} /* (6, 8, 23) {real, imag} */,
  {32'h4015e218, 32'h40264048} /* (6, 8, 22) {real, imag} */,
  {32'h40be8654, 32'h40305be8} /* (6, 8, 21) {real, imag} */,
  {32'hc0e71d94, 32'h4067e8e8} /* (6, 8, 20) {real, imag} */,
  {32'hc12de85b, 32'hc1401ed3} /* (6, 8, 19) {real, imag} */,
  {32'hc0925376, 32'hc18b8e97} /* (6, 8, 18) {real, imag} */,
  {32'h4151b1ce, 32'hc0bf2d74} /* (6, 8, 17) {real, imag} */,
  {32'hbea53800, 32'hc00614ee} /* (6, 8, 16) {real, imag} */,
  {32'hc0c7021a, 32'hc0346608} /* (6, 8, 15) {real, imag} */,
  {32'h41685d89, 32'hc13606cf} /* (6, 8, 14) {real, imag} */,
  {32'h41753108, 32'hc0b00bbe} /* (6, 8, 13) {real, imag} */,
  {32'h40a3215c, 32'h3d9f2cc0} /* (6, 8, 12) {real, imag} */,
  {32'h4039b764, 32'hbc18ca00} /* (6, 8, 11) {real, imag} */,
  {32'hc05b15c0, 32'h4091d1a0} /* (6, 8, 10) {real, imag} */,
  {32'hc0cb0af1, 32'hc0a1d978} /* (6, 8, 9) {real, imag} */,
  {32'hc15dcd24, 32'hc181887b} /* (6, 8, 8) {real, imag} */,
  {32'hc13f6cd4, 32'hc0b02c6b} /* (6, 8, 7) {real, imag} */,
  {32'hc10b07e1, 32'h40c4f114} /* (6, 8, 6) {real, imag} */,
  {32'h3f128888, 32'h40ac8fdb} /* (6, 8, 5) {real, imag} */,
  {32'h418cdb01, 32'h3f3f0808} /* (6, 8, 4) {real, imag} */,
  {32'h4104f301, 32'hbf9b7fdc} /* (6, 8, 3) {real, imag} */,
  {32'h3f0c8b98, 32'h406e4628} /* (6, 8, 2) {real, imag} */,
  {32'hc0c5747a, 32'h40d5b2f6} /* (6, 8, 1) {real, imag} */,
  {32'hc143c704, 32'h3f26b180} /* (6, 8, 0) {real, imag} */,
  {32'h41483cd0, 32'h40045fe9} /* (6, 7, 31) {real, imag} */,
  {32'h4012cf49, 32'hc0b9183c} /* (6, 7, 30) {real, imag} */,
  {32'hbea4b71e, 32'hc062ceb7} /* (6, 7, 29) {real, imag} */,
  {32'hc11429e0, 32'hbfe7242c} /* (6, 7, 28) {real, imag} */,
  {32'hc19cec82, 32'h4071d218} /* (6, 7, 27) {real, imag} */,
  {32'hc0bf9979, 32'h4177b7ef} /* (6, 7, 26) {real, imag} */,
  {32'hc1238dd2, 32'hbcdd7a00} /* (6, 7, 25) {real, imag} */,
  {32'hc0655783, 32'hc12bf66a} /* (6, 7, 24) {real, imag} */,
  {32'h4125ea92, 32'hc08bb9b9} /* (6, 7, 23) {real, imag} */,
  {32'h40a65e84, 32'h40feb5b0} /* (6, 7, 22) {real, imag} */,
  {32'hc1c4d270, 32'hc138eb2f} /* (6, 7, 21) {real, imag} */,
  {32'hc1c6ca62, 32'hc1428c52} /* (6, 7, 20) {real, imag} */,
  {32'hc1c18400, 32'hc1b14c4e} /* (6, 7, 19) {real, imag} */,
  {32'hc093ef16, 32'hc1a06440} /* (6, 7, 18) {real, imag} */,
  {32'hbec68e30, 32'hc10c9106} /* (6, 7, 17) {real, imag} */,
  {32'hbf0d3c20, 32'hc1408919} /* (6, 7, 16) {real, imag} */,
  {32'hc0e9ec3c, 32'hc161cff4} /* (6, 7, 15) {real, imag} */,
  {32'h402b77ac, 32'hc0cf37cc} /* (6, 7, 14) {real, imag} */,
  {32'hbf7d8a04, 32'hc0d1adaf} /* (6, 7, 13) {real, imag} */,
  {32'h401b4d1e, 32'h40dbe295} /* (6, 7, 12) {real, imag} */,
  {32'h409fb32b, 32'h413e534e} /* (6, 7, 11) {real, imag} */,
  {32'h41cbfd72, 32'h4001985a} /* (6, 7, 10) {real, imag} */,
  {32'h41af0efc, 32'hc081285a} /* (6, 7, 9) {real, imag} */,
  {32'h40325828, 32'hc038581a} /* (6, 7, 8) {real, imag} */,
  {32'hbeff5d60, 32'hc1819063} /* (6, 7, 7) {real, imag} */,
  {32'hc0deb3ba, 32'hc1b56d31} /* (6, 7, 6) {real, imag} */,
  {32'hc14c072f, 32'hc0dbacc0} /* (6, 7, 5) {real, imag} */,
  {32'hc1566b74, 32'hbfee291c} /* (6, 7, 4) {real, imag} */,
  {32'hc0878fbe, 32'hc11123cb} /* (6, 7, 3) {real, imag} */,
  {32'hc0f15a76, 32'h4011b4f2} /* (6, 7, 2) {real, imag} */,
  {32'h4177f768, 32'hc05cc22c} /* (6, 7, 1) {real, imag} */,
  {32'h4142cbc5, 32'hc0c1fc34} /* (6, 7, 0) {real, imag} */,
  {32'h40021202, 32'hbf451580} /* (6, 6, 31) {real, imag} */,
  {32'hbfc602e2, 32'h40cbf762} /* (6, 6, 30) {real, imag} */,
  {32'hc01ecca2, 32'hc0adc50c} /* (6, 6, 29) {real, imag} */,
  {32'hbf0868f8, 32'hc155b336} /* (6, 6, 28) {real, imag} */,
  {32'hbeac6050, 32'hc1beb212} /* (6, 6, 27) {real, imag} */,
  {32'h40d1939a, 32'hbd8de780} /* (6, 6, 26) {real, imag} */,
  {32'h41849b24, 32'h411bcde0} /* (6, 6, 25) {real, imag} */,
  {32'h419969b2, 32'hc1881d85} /* (6, 6, 24) {real, imag} */,
  {32'h40e3993f, 32'hbdd8c3e0} /* (6, 6, 23) {real, imag} */,
  {32'hc0f81279, 32'h3fa9da74} /* (6, 6, 22) {real, imag} */,
  {32'hc1062cac, 32'hc100eaee} /* (6, 6, 21) {real, imag} */,
  {32'hc126008a, 32'h3fa9dfca} /* (6, 6, 20) {real, imag} */,
  {32'h40cd9ff2, 32'h4071a5f7} /* (6, 6, 19) {real, imag} */,
  {32'h41061ad2, 32'hc094ae3b} /* (6, 6, 18) {real, imag} */,
  {32'hc0e357a6, 32'hc12d1eae} /* (6, 6, 17) {real, imag} */,
  {32'hc1909b01, 32'h411625e8} /* (6, 6, 16) {real, imag} */,
  {32'hc013fed5, 32'h4067739c} /* (6, 6, 15) {real, imag} */,
  {32'hc0e5d31b, 32'hc13302da} /* (6, 6, 14) {real, imag} */,
  {32'hc11b3a04, 32'hc1ab3c00} /* (6, 6, 13) {real, imag} */,
  {32'h4114d28b, 32'h407e063c} /* (6, 6, 12) {real, imag} */,
  {32'h410aee29, 32'hc038e1cc} /* (6, 6, 11) {real, imag} */,
  {32'h4188ac4c, 32'hc19d70e0} /* (6, 6, 10) {real, imag} */,
  {32'h40ed880e, 32'hc141c43e} /* (6, 6, 9) {real, imag} */,
  {32'hc109095b, 32'hbee4eaf0} /* (6, 6, 8) {real, imag} */,
  {32'hc1965d60, 32'h410b1937} /* (6, 6, 7) {real, imag} */,
  {32'hc102a7fe, 32'h41a98048} /* (6, 6, 6) {real, imag} */,
  {32'h41170512, 32'h404b1004} /* (6, 6, 5) {real, imag} */,
  {32'hc03217a2, 32'h408ddcbb} /* (6, 6, 4) {real, imag} */,
  {32'hc17296c3, 32'h3fcfd22e} /* (6, 6, 3) {real, imag} */,
  {32'hc012a516, 32'h3f0d98e0} /* (6, 6, 2) {real, imag} */,
  {32'h3f53b158, 32'hc15125c2} /* (6, 6, 1) {real, imag} */,
  {32'hc071e7ec, 32'hc0dfbf14} /* (6, 6, 0) {real, imag} */,
  {32'h40ba98b6, 32'hbfdb9239} /* (6, 5, 31) {real, imag} */,
  {32'hc134ae80, 32'hc05d5a98} /* (6, 5, 30) {real, imag} */,
  {32'hc178eeb5, 32'hc0e61de0} /* (6, 5, 29) {real, imag} */,
  {32'hc19a8424, 32'hc0696d82} /* (6, 5, 28) {real, imag} */,
  {32'h403dd23c, 32'h3dbb5ce0} /* (6, 5, 27) {real, imag} */,
  {32'h400fbe5f, 32'hbfa00517} /* (6, 5, 26) {real, imag} */,
  {32'h40cceec5, 32'h40ef2e74} /* (6, 5, 25) {real, imag} */,
  {32'hc1a1bfea, 32'h41770bde} /* (6, 5, 24) {real, imag} */,
  {32'hc11c857e, 32'h41a6afd6} /* (6, 5, 23) {real, imag} */,
  {32'hc151d7b1, 32'h40064a10} /* (6, 5, 22) {real, imag} */,
  {32'hc1871d05, 32'hc12d8e22} /* (6, 5, 21) {real, imag} */,
  {32'hc1b50858, 32'hc18f8ad4} /* (6, 5, 20) {real, imag} */,
  {32'hc085e712, 32'hc146ef67} /* (6, 5, 19) {real, imag} */,
  {32'h40ddc392, 32'h3eca7598} /* (6, 5, 18) {real, imag} */,
  {32'h41120116, 32'hc0c0ffe2} /* (6, 5, 17) {real, imag} */,
  {32'hc1066a59, 32'h4121cd13} /* (6, 5, 16) {real, imag} */,
  {32'hc09aa362, 32'h4174ad8d} /* (6, 5, 15) {real, imag} */,
  {32'hc103f04d, 32'hc0d26dfe} /* (6, 5, 14) {real, imag} */,
  {32'hc11d7c80, 32'h414066ab} /* (6, 5, 13) {real, imag} */,
  {32'hc094b811, 32'h410801a2} /* (6, 5, 12) {real, imag} */,
  {32'hc12ef74e, 32'hbf39f5a0} /* (6, 5, 11) {real, imag} */,
  {32'hc159c5f7, 32'h419d0fde} /* (6, 5, 10) {real, imag} */,
  {32'hc09e140e, 32'h41be8526} /* (6, 5, 9) {real, imag} */,
  {32'h40014661, 32'h402b8912} /* (6, 5, 8) {real, imag} */,
  {32'hbf13ff18, 32'hbf741340} /* (6, 5, 7) {real, imag} */,
  {32'hc06b091c, 32'hbfa2ff35} /* (6, 5, 6) {real, imag} */,
  {32'h41190ee4, 32'h3f4b6580} /* (6, 5, 5) {real, imag} */,
  {32'h40a328b3, 32'hc152e158} /* (6, 5, 4) {real, imag} */,
  {32'h40ecd88c, 32'hc15f8587} /* (6, 5, 3) {real, imag} */,
  {32'h419a5463, 32'h410de52f} /* (6, 5, 2) {real, imag} */,
  {32'hc00d9197, 32'h416c92d2} /* (6, 5, 1) {real, imag} */,
  {32'hc10e566c, 32'hc061051e} /* (6, 5, 0) {real, imag} */,
  {32'hbf628828, 32'hc0d2f89c} /* (6, 4, 31) {real, imag} */,
  {32'h416a1673, 32'hc0c178ac} /* (6, 4, 30) {real, imag} */,
  {32'h409164c4, 32'h4121fca2} /* (6, 4, 29) {real, imag} */,
  {32'hc0eab624, 32'h411a8dd6} /* (6, 4, 28) {real, imag} */,
  {32'h412b5b4f, 32'h4127d73d} /* (6, 4, 27) {real, imag} */,
  {32'h41b5fe04, 32'h40a91c56} /* (6, 4, 26) {real, imag} */,
  {32'h417087f5, 32'h3f3b4e8c} /* (6, 4, 25) {real, imag} */,
  {32'hc01bbeca, 32'h409b282e} /* (6, 4, 24) {real, imag} */,
  {32'hc083ff9a, 32'hc189a918} /* (6, 4, 23) {real, imag} */,
  {32'hc15f4762, 32'hc1e857b2} /* (6, 4, 22) {real, imag} */,
  {32'hc180a836, 32'hc1ccf3e6} /* (6, 4, 21) {real, imag} */,
  {32'h411285d2, 32'hc1ad468a} /* (6, 4, 20) {real, imag} */,
  {32'h411aa412, 32'hbea03b60} /* (6, 4, 19) {real, imag} */,
  {32'hc092a08a, 32'h419b75b0} /* (6, 4, 18) {real, imag} */,
  {32'hc0a03eb2, 32'h40fc7460} /* (6, 4, 17) {real, imag} */,
  {32'h41312c8f, 32'hc0b9261c} /* (6, 4, 16) {real, imag} */,
  {32'hc0d40007, 32'h40bccd37} /* (6, 4, 15) {real, imag} */,
  {32'hc180488f, 32'hc06b7e72} /* (6, 4, 14) {real, imag} */,
  {32'h3fdf6a08, 32'hc0eb25d0} /* (6, 4, 13) {real, imag} */,
  {32'h412b9508, 32'hc1745070} /* (6, 4, 12) {real, imag} */,
  {32'h413afc7e, 32'hc1298160} /* (6, 4, 11) {real, imag} */,
  {32'h415ec53c, 32'hbeee12a0} /* (6, 4, 10) {real, imag} */,
  {32'hbfa43684, 32'hbe26e5f8} /* (6, 4, 9) {real, imag} */,
  {32'hc035ae5c, 32'h3e84dd18} /* (6, 4, 8) {real, imag} */,
  {32'h3f5a29cd, 32'h41b0db76} /* (6, 4, 7) {real, imag} */,
  {32'h412446ee, 32'h4014558c} /* (6, 4, 6) {real, imag} */,
  {32'h40db83c4, 32'hc0618e9e} /* (6, 4, 5) {real, imag} */,
  {32'h40826718, 32'h40dd6828} /* (6, 4, 4) {real, imag} */,
  {32'h4141f036, 32'h41908bab} /* (6, 4, 3) {real, imag} */,
  {32'h40f3c6de, 32'h3f881d48} /* (6, 4, 2) {real, imag} */,
  {32'h40a4c0c8, 32'hc134a6fc} /* (6, 4, 1) {real, imag} */,
  {32'hc0695a02, 32'hc023ba81} /* (6, 4, 0) {real, imag} */,
  {32'hbf1c4234, 32'h414c8ea4} /* (6, 3, 31) {real, imag} */,
  {32'h40b9262d, 32'h414a1181} /* (6, 3, 30) {real, imag} */,
  {32'hc0d412c1, 32'h4010fcbc} /* (6, 3, 29) {real, imag} */,
  {32'h40adc20c, 32'h3fe1d570} /* (6, 3, 28) {real, imag} */,
  {32'h40775778, 32'h3ffba9e4} /* (6, 3, 27) {real, imag} */,
  {32'hc0a0995a, 32'h4038c370} /* (6, 3, 26) {real, imag} */,
  {32'hc137c16e, 32'hc16a1e80} /* (6, 3, 25) {real, imag} */,
  {32'hc18bb5ed, 32'h3efd32a0} /* (6, 3, 24) {real, imag} */,
  {32'hc1cbc976, 32'hbf9ecf40} /* (6, 3, 23) {real, imag} */,
  {32'hc18da45c, 32'h409bde83} /* (6, 3, 22) {real, imag} */,
  {32'hc1592f37, 32'h4162d853} /* (6, 3, 21) {real, imag} */,
  {32'hc194db4c, 32'h411a697e} /* (6, 3, 20) {real, imag} */,
  {32'hc19c2555, 32'hc0cd02de} /* (6, 3, 19) {real, imag} */,
  {32'h4030ec54, 32'hc11a3104} /* (6, 3, 18) {real, imag} */,
  {32'h3f59953e, 32'h412f58ac} /* (6, 3, 17) {real, imag} */,
  {32'h3f23c228, 32'h4083849e} /* (6, 3, 16) {real, imag} */,
  {32'h41157a4c, 32'h406d09d3} /* (6, 3, 15) {real, imag} */,
  {32'hbef78b48, 32'hc1283b03} /* (6, 3, 14) {real, imag} */,
  {32'hbfdbcf5e, 32'hc19e20e6} /* (6, 3, 13) {real, imag} */,
  {32'h4105f7b4, 32'hbfba93b6} /* (6, 3, 12) {real, imag} */,
  {32'hc1784728, 32'h413f5622} /* (6, 3, 11) {real, imag} */,
  {32'hbfa30d4f, 32'h41820d70} /* (6, 3, 10) {real, imag} */,
  {32'h41271766, 32'h41738f7c} /* (6, 3, 9) {real, imag} */,
  {32'h409842be, 32'h418dc0cb} /* (6, 3, 8) {real, imag} */,
  {32'h414b248f, 32'hc047c4f8} /* (6, 3, 7) {real, imag} */,
  {32'h41352d41, 32'h408c1ae0} /* (6, 3, 6) {real, imag} */,
  {32'hc1128503, 32'h3f8b91a5} /* (6, 3, 5) {real, imag} */,
  {32'h3efaa748, 32'h3ed35a10} /* (6, 3, 4) {real, imag} */,
  {32'h41486f5d, 32'h40d31e04} /* (6, 3, 3) {real, imag} */,
  {32'h4138c7ae, 32'h413d3fa4} /* (6, 3, 2) {real, imag} */,
  {32'h41383870, 32'hc0c468e5} /* (6, 3, 1) {real, imag} */,
  {32'h41177bc9, 32'hc0cebf74} /* (6, 3, 0) {real, imag} */,
  {32'h40d5733b, 32'hc1368c98} /* (6, 2, 31) {real, imag} */,
  {32'h41457f73, 32'hc1a621bc} /* (6, 2, 30) {real, imag} */,
  {32'h410eb998, 32'hc0d11a74} /* (6, 2, 29) {real, imag} */,
  {32'h405cba7b, 32'h416b536a} /* (6, 2, 28) {real, imag} */,
  {32'hc1010c17, 32'h41c6ff32} /* (6, 2, 27) {real, imag} */,
  {32'hc0602a40, 32'h41b6fbc4} /* (6, 2, 26) {real, imag} */,
  {32'hc0dd92c4, 32'h41cb514e} /* (6, 2, 25) {real, imag} */,
  {32'hc1172d66, 32'h41c49bee} /* (6, 2, 24) {real, imag} */,
  {32'h41023df4, 32'hc08621fb} /* (6, 2, 23) {real, imag} */,
  {32'h4189ed30, 32'h407d8670} /* (6, 2, 22) {real, imag} */,
  {32'h4021f8e0, 32'h4142729c} /* (6, 2, 21) {real, imag} */,
  {32'hc13b337e, 32'hc175eef3} /* (6, 2, 20) {real, imag} */,
  {32'hc14803cc, 32'hc181944c} /* (6, 2, 19) {real, imag} */,
  {32'hc19ef69f, 32'h3f3131c8} /* (6, 2, 18) {real, imag} */,
  {32'hc15113de, 32'h40d83404} /* (6, 2, 17) {real, imag} */,
  {32'hc1281ab6, 32'hc119c9f8} /* (6, 2, 16) {real, imag} */,
  {32'hc0b26899, 32'hc1e8da1d} /* (6, 2, 15) {real, imag} */,
  {32'h3f035080, 32'hc16e7148} /* (6, 2, 14) {real, imag} */,
  {32'hc0cbe9b4, 32'h41042ad6} /* (6, 2, 13) {real, imag} */,
  {32'hc0daa818, 32'h4041b27f} /* (6, 2, 12) {real, imag} */,
  {32'hc19405eb, 32'hc168e06b} /* (6, 2, 11) {real, imag} */,
  {32'hc173b69c, 32'hc1d88082} /* (6, 2, 10) {real, imag} */,
  {32'hc07c5bd0, 32'hc1f5e5eb} /* (6, 2, 9) {real, imag} */,
  {32'h3ecf5110, 32'hc158ee90} /* (6, 2, 8) {real, imag} */,
  {32'hc13cd110, 32'hc1acb77b} /* (6, 2, 7) {real, imag} */,
  {32'hc087c48a, 32'hc1afdec2} /* (6, 2, 6) {real, imag} */,
  {32'h418f83e8, 32'hc0898306} /* (6, 2, 5) {real, imag} */,
  {32'h4172e22a, 32'hc06c9e47} /* (6, 2, 4) {real, imag} */,
  {32'h40b13d0a, 32'hc186faa7} /* (6, 2, 3) {real, imag} */,
  {32'h40f19f10, 32'hc14bbee0} /* (6, 2, 2) {real, imag} */,
  {32'hc0910ae0, 32'hc0a7ab38} /* (6, 2, 1) {real, imag} */,
  {32'hc09a5679, 32'h3fe0357a} /* (6, 2, 0) {real, imag} */,
  {32'h411faa00, 32'h3fda2ff8} /* (6, 1, 31) {real, imag} */,
  {32'h416e7c65, 32'h3fc559ca} /* (6, 1, 30) {real, imag} */,
  {32'hc0a5221c, 32'h3efafeb0} /* (6, 1, 29) {real, imag} */,
  {32'h40a18041, 32'hc19ce0d3} /* (6, 1, 28) {real, imag} */,
  {32'h41762b6e, 32'hc0461fb4} /* (6, 1, 27) {real, imag} */,
  {32'h41921260, 32'h4086359e} /* (6, 1, 26) {real, imag} */,
  {32'h419ecb7a, 32'hbf18427c} /* (6, 1, 25) {real, imag} */,
  {32'h4135fd88, 32'hc056d9fc} /* (6, 1, 24) {real, imag} */,
  {32'h410122db, 32'hc138864a} /* (6, 1, 23) {real, imag} */,
  {32'hbfe11474, 32'hc08d6a36} /* (6, 1, 22) {real, imag} */,
  {32'hc0871573, 32'hc18a9048} /* (6, 1, 21) {real, imag} */,
  {32'hc07b0302, 32'hc15c442e} /* (6, 1, 20) {real, imag} */,
  {32'h419bdd83, 32'hc0d45078} /* (6, 1, 19) {real, imag} */,
  {32'hc0d2f246, 32'hc04d8290} /* (6, 1, 18) {real, imag} */,
  {32'h414257ef, 32'hc1368deb} /* (6, 1, 17) {real, imag} */,
  {32'h41921cef, 32'hc0dee017} /* (6, 1, 16) {real, imag} */,
  {32'hc0df388c, 32'h4196147a} /* (6, 1, 15) {real, imag} */,
  {32'hbf06fd58, 32'hc0691630} /* (6, 1, 14) {real, imag} */,
  {32'hc12323d7, 32'h3e9a2050} /* (6, 1, 13) {real, imag} */,
  {32'hc0d88c40, 32'hc09a22b0} /* (6, 1, 12) {real, imag} */,
  {32'h40b64b3a, 32'hc144fc20} /* (6, 1, 11) {real, imag} */,
  {32'h412c8c60, 32'h3e913ac0} /* (6, 1, 10) {real, imag} */,
  {32'h416bc3aa, 32'h409b13e9} /* (6, 1, 9) {real, imag} */,
  {32'h4092e2b7, 32'h4119b244} /* (6, 1, 8) {real, imag} */,
  {32'h41be2263, 32'hbe235840} /* (6, 1, 7) {real, imag} */,
  {32'h41183aff, 32'hbfb34ad8} /* (6, 1, 6) {real, imag} */,
  {32'hc10f34e1, 32'hbf01de46} /* (6, 1, 5) {real, imag} */,
  {32'hc149c6f9, 32'hc121cf95} /* (6, 1, 4) {real, imag} */,
  {32'hc0a1ac15, 32'hc0878f76} /* (6, 1, 3) {real, imag} */,
  {32'hc0062024, 32'h404d0478} /* (6, 1, 2) {real, imag} */,
  {32'hc005fd6c, 32'hc1834d9a} /* (6, 1, 1) {real, imag} */,
  {32'h3fa126b4, 32'hc0b1db62} /* (6, 1, 0) {real, imag} */,
  {32'hbf9d737d, 32'h4149dba6} /* (6, 0, 31) {real, imag} */,
  {32'h407d447e, 32'h418e817c} /* (6, 0, 30) {real, imag} */,
  {32'h40afbca7, 32'hbfe41e28} /* (6, 0, 29) {real, imag} */,
  {32'h415fe426, 32'hc0133864} /* (6, 0, 28) {real, imag} */,
  {32'h420d7cb8, 32'hc1286eaf} /* (6, 0, 27) {real, imag} */,
  {32'h41690027, 32'hbc838940} /* (6, 0, 26) {real, imag} */,
  {32'hc167f54c, 32'hbf0729fa} /* (6, 0, 25) {real, imag} */,
  {32'hc16063e6, 32'hc0944c26} /* (6, 0, 24) {real, imag} */,
  {32'h401c3b7c, 32'hc149156e} /* (6, 0, 23) {real, imag} */,
  {32'h3f82d9db, 32'h40e13c16} /* (6, 0, 22) {real, imag} */,
  {32'hc0a7a5ac, 32'h4161b288} /* (6, 0, 21) {real, imag} */,
  {32'h40f52ba8, 32'h41271d50} /* (6, 0, 20) {real, imag} */,
  {32'h40cce176, 32'h41a9d9a6} /* (6, 0, 19) {real, imag} */,
  {32'hbfd06b9c, 32'h414e03fb} /* (6, 0, 18) {real, imag} */,
  {32'hc1b4dac8, 32'hc0e26cc0} /* (6, 0, 17) {real, imag} */,
  {32'hc0b34c12, 32'hbfedea97} /* (6, 0, 16) {real, imag} */,
  {32'h41025134, 32'hc0fb4b62} /* (6, 0, 15) {real, imag} */,
  {32'h41a07ef0, 32'hbf933358} /* (6, 0, 14) {real, imag} */,
  {32'h41932ee0, 32'hc113216c} /* (6, 0, 13) {real, imag} */,
  {32'hc02e346b, 32'h41273e9c} /* (6, 0, 12) {real, imag} */,
  {32'h40aba765, 32'h40bd073e} /* (6, 0, 11) {real, imag} */,
  {32'h41065d94, 32'h403cb2b6} /* (6, 0, 10) {real, imag} */,
  {32'h41816b7b, 32'hc15de666} /* (6, 0, 9) {real, imag} */,
  {32'h418a2463, 32'hc1c8406b} /* (6, 0, 8) {real, imag} */,
  {32'h411f867a, 32'h410bdec6} /* (6, 0, 7) {real, imag} */,
  {32'h40bcde53, 32'h41bbe78e} /* (6, 0, 6) {real, imag} */,
  {32'hc085a720, 32'h41ef2474} /* (6, 0, 5) {real, imag} */,
  {32'h3faf5698, 32'h41929fe1} /* (6, 0, 4) {real, imag} */,
  {32'h40ad4412, 32'h4110090d} /* (6, 0, 3) {real, imag} */,
  {32'h3faef542, 32'h41c7fd6c} /* (6, 0, 2) {real, imag} */,
  {32'h41badcd6, 32'h414664e4} /* (6, 0, 1) {real, imag} */,
  {32'h40c7a96a, 32'h40acd8cd} /* (6, 0, 0) {real, imag} */,
  {32'h40f0b81e, 32'hc13fcfa9} /* (5, 31, 31) {real, imag} */,
  {32'h41b01f16, 32'hc1f22923} /* (5, 31, 30) {real, imag} */,
  {32'h41c5b21e, 32'hc22e928a} /* (5, 31, 29) {real, imag} */,
  {32'h40831298, 32'hc24faf03} /* (5, 31, 28) {real, imag} */,
  {32'h40f42aac, 32'hc2651664} /* (5, 31, 27) {real, imag} */,
  {32'h3f1db780, 32'hc20f20bf} /* (5, 31, 26) {real, imag} */,
  {32'h417d6801, 32'hc20650c7} /* (5, 31, 25) {real, imag} */,
  {32'h41d1a7bc, 32'hc21a0fee} /* (5, 31, 24) {real, imag} */,
  {32'h41d67649, 32'hc25585b2} /* (5, 31, 23) {real, imag} */,
  {32'h42121dee, 32'hc2674deb} /* (5, 31, 22) {real, imag} */,
  {32'h40d05913, 32'hc1ba36b7} /* (5, 31, 21) {real, imag} */,
  {32'hc0d6f8de, 32'h4100bb60} /* (5, 31, 20) {real, imag} */,
  {32'hc17fc930, 32'h40476842} /* (5, 31, 19) {real, imag} */,
  {32'hc0e48696, 32'hbef30258} /* (5, 31, 18) {real, imag} */,
  {32'hc0ac8542, 32'h41a40716} /* (5, 31, 17) {real, imag} */,
  {32'h400e0282, 32'h41bce76e} /* (5, 31, 16) {real, imag} */,
  {32'hc0b89af4, 32'h41e4c922} /* (5, 31, 15) {real, imag} */,
  {32'hc1321fb6, 32'h4129692f} /* (5, 31, 14) {real, imag} */,
  {32'hc184e75c, 32'h41e785d0} /* (5, 31, 13) {real, imag} */,
  {32'hc1be54e8, 32'h4255d7a9} /* (5, 31, 12) {real, imag} */,
  {32'hc1a6f8eb, 32'h42316608} /* (5, 31, 11) {real, imag} */,
  {32'hc0e3d9d0, 32'hc0bf5cf7} /* (5, 31, 10) {real, imag} */,
  {32'hc0152810, 32'hc19ab767} /* (5, 31, 9) {real, imag} */,
  {32'hc1c23328, 32'hc1a2e8a2} /* (5, 31, 8) {real, imag} */,
  {32'hc194b69b, 32'hc1bece02} /* (5, 31, 7) {real, imag} */,
  {32'h3e9bdec8, 32'hc234b65b} /* (5, 31, 6) {real, imag} */,
  {32'h419a0606, 32'hc2513ec0} /* (5, 31, 5) {real, imag} */,
  {32'h41f734cc, 32'hc1c738c6} /* (5, 31, 4) {real, imag} */,
  {32'h4186846f, 32'hc1d32f87} /* (5, 31, 3) {real, imag} */,
  {32'h41f9fb38, 32'hc213d026} /* (5, 31, 2) {real, imag} */,
  {32'h41f8f920, 32'hc22c04f4} /* (5, 31, 1) {real, imag} */,
  {32'h41a30c1c, 32'hc1a10bd4} /* (5, 31, 0) {real, imag} */,
  {32'hc1565358, 32'h41906245} /* (5, 30, 31) {real, imag} */,
  {32'hc1139f17, 32'h4201c38a} /* (5, 30, 30) {real, imag} */,
  {32'h41818a1b, 32'h425332ac} /* (5, 30, 29) {real, imag} */,
  {32'h4146b7fa, 32'h42292426} /* (5, 30, 28) {real, imag} */,
  {32'hbf330aa0, 32'h4214f9b2} /* (5, 30, 27) {real, imag} */,
  {32'hc09d85cc, 32'h42098e8a} /* (5, 30, 26) {real, imag} */,
  {32'hc06c9d80, 32'h42113984} /* (5, 30, 25) {real, imag} */,
  {32'hc1712681, 32'h41e8903f} /* (5, 30, 24) {real, imag} */,
  {32'hc1d1702a, 32'h42110f6b} /* (5, 30, 23) {real, imag} */,
  {32'hc11db018, 32'h423f75a0} /* (5, 30, 22) {real, imag} */,
  {32'h41386678, 32'h41d742bf} /* (5, 30, 21) {real, imag} */,
  {32'h41f29fe8, 32'hc0772e0a} /* (5, 30, 20) {real, imag} */,
  {32'h4186a597, 32'hc1e13660} /* (5, 30, 19) {real, imag} */,
  {32'h41d52280, 32'hc1a646a2} /* (5, 30, 18) {real, imag} */,
  {32'h423be7a7, 32'hc1bb558f} /* (5, 30, 17) {real, imag} */,
  {32'h425c1097, 32'hc1b11cec} /* (5, 30, 16) {real, imag} */,
  {32'h419c9259, 32'hc1bb88d0} /* (5, 30, 15) {real, imag} */,
  {32'h40bf2046, 32'hc2024056} /* (5, 30, 14) {real, imag} */,
  {32'h41259904, 32'hc1e681c0} /* (5, 30, 13) {real, imag} */,
  {32'h41b98eb2, 32'hc124a2fe} /* (5, 30, 12) {real, imag} */,
  {32'h42085645, 32'hc090d7c6} /* (5, 30, 11) {real, imag} */,
  {32'hc092348e, 32'h415427d1} /* (5, 30, 10) {real, imag} */,
  {32'hc1a87558, 32'h420f8550} /* (5, 30, 9) {real, imag} */,
  {32'hc2061445, 32'h42594513} /* (5, 30, 8) {real, imag} */,
  {32'hc1571d46, 32'h420b96bc} /* (5, 30, 7) {real, imag} */,
  {32'hc071412b, 32'h41c0f3a2} /* (5, 30, 6) {real, imag} */,
  {32'hc0fd6dfe, 32'h418d61bb} /* (5, 30, 5) {real, imag} */,
  {32'hc100c96a, 32'h41b54386} /* (5, 30, 4) {real, imag} */,
  {32'hc189cfc2, 32'h4177aa7a} /* (5, 30, 3) {real, imag} */,
  {32'hc162a41f, 32'h40ffdf19} /* (5, 30, 2) {real, imag} */,
  {32'hc17e4a25, 32'h41db31d2} /* (5, 30, 1) {real, imag} */,
  {32'hc06d42eb, 32'h420500ce} /* (5, 30, 0) {real, imag} */,
  {32'h40d1c523, 32'hc1421831} /* (5, 29, 31) {real, imag} */,
  {32'h40990063, 32'hc15ef639} /* (5, 29, 30) {real, imag} */,
  {32'hc0ed4d89, 32'hc10a9bad} /* (5, 29, 29) {real, imag} */,
  {32'hc13748cb, 32'h40afb0d7} /* (5, 29, 28) {real, imag} */,
  {32'hc115ed90, 32'hc195a0e4} /* (5, 29, 27) {real, imag} */,
  {32'hc0d63046, 32'h40c3f891} /* (5, 29, 26) {real, imag} */,
  {32'hc1465bce, 32'h41c0e272} /* (5, 29, 25) {real, imag} */,
  {32'hc0614af3, 32'h408f5a78} /* (5, 29, 24) {real, imag} */,
  {32'h4189d1c7, 32'hc16a5049} /* (5, 29, 23) {real, imag} */,
  {32'h41899770, 32'hc15bff6a} /* (5, 29, 22) {real, imag} */,
  {32'h41652804, 32'h4186f1a9} /* (5, 29, 21) {real, imag} */,
  {32'h41150df2, 32'h41a20f58} /* (5, 29, 20) {real, imag} */,
  {32'h415797fa, 32'h40efc4fd} /* (5, 29, 19) {real, imag} */,
  {32'h424f68e3, 32'hc02ad69c} /* (5, 29, 18) {real, imag} */,
  {32'h4238cff0, 32'hc108ff90} /* (5, 29, 17) {real, imag} */,
  {32'h41b0de57, 32'hbf1760ec} /* (5, 29, 16) {real, imag} */,
  {32'h41590796, 32'hbe1342e0} /* (5, 29, 15) {real, imag} */,
  {32'hc0f21222, 32'hc1ad1413} /* (5, 29, 14) {real, imag} */,
  {32'h4019c142, 32'hc194b550} /* (5, 29, 13) {real, imag} */,
  {32'h415ebeec, 32'hbeed2fc0} /* (5, 29, 12) {real, imag} */,
  {32'h4185aa1e, 32'h3f9dcf78} /* (5, 29, 11) {real, imag} */,
  {32'hc12e6826, 32'hc0afcff1} /* (5, 29, 10) {real, imag} */,
  {32'hc1ccadfb, 32'hc1075b83} /* (5, 29, 9) {real, imag} */,
  {32'hc03002c7, 32'hc1a51e1f} /* (5, 29, 8) {real, imag} */,
  {32'hc0c7dec8, 32'hc1b820d2} /* (5, 29, 7) {real, imag} */,
  {32'hc1ed735d, 32'hc2028119} /* (5, 29, 6) {real, imag} */,
  {32'hc0c6ecb2, 32'h40e69752} /* (5, 29, 5) {real, imag} */,
  {32'h40c20216, 32'h4104b0de} /* (5, 29, 4) {real, imag} */,
  {32'h408db512, 32'hc0e9f9dd} /* (5, 29, 3) {real, imag} */,
  {32'hbe8aea60, 32'hc15b3f16} /* (5, 29, 2) {real, imag} */,
  {32'h4023be54, 32'hbf55ea70} /* (5, 29, 1) {real, imag} */,
  {32'h40935765, 32'hbfbd8bf0} /* (5, 29, 0) {real, imag} */,
  {32'h4016d954, 32'h40bc621e} /* (5, 28, 31) {real, imag} */,
  {32'hc084c748, 32'h40f5786b} /* (5, 28, 30) {real, imag} */,
  {32'hc144af16, 32'hc10a6dca} /* (5, 28, 29) {real, imag} */,
  {32'h3fc523ee, 32'hc187696c} /* (5, 28, 28) {real, imag} */,
  {32'h3ecc9d10, 32'hc12e0032} /* (5, 28, 27) {real, imag} */,
  {32'h4162ae85, 32'hc171cc7f} /* (5, 28, 26) {real, imag} */,
  {32'h40d3f9ce, 32'hc1109af6} /* (5, 28, 25) {real, imag} */,
  {32'h413f4262, 32'h40ec9fe5} /* (5, 28, 24) {real, imag} */,
  {32'h3f28ffc0, 32'h40d873e5} /* (5, 28, 23) {real, imag} */,
  {32'hbfea6c80, 32'h40b4f4e0} /* (5, 28, 22) {real, imag} */,
  {32'h41188291, 32'h41e30548} /* (5, 28, 21) {real, imag} */,
  {32'h41bdb69c, 32'h422ffc86} /* (5, 28, 20) {real, imag} */,
  {32'h41dff912, 32'h420b65d6} /* (5, 28, 19) {real, imag} */,
  {32'h4127e734, 32'h41ab3532} /* (5, 28, 18) {real, imag} */,
  {32'h408223b8, 32'h4198b2e0} /* (5, 28, 17) {real, imag} */,
  {32'hc0311e44, 32'h410680af} /* (5, 28, 16) {real, imag} */,
  {32'h40f44828, 32'h415424d6} /* (5, 28, 15) {real, imag} */,
  {32'h4155ac71, 32'h418b19a0} /* (5, 28, 14) {real, imag} */,
  {32'hc057a7e2, 32'h41ba52cd} /* (5, 28, 13) {real, imag} */,
  {32'hc158b76e, 32'h41147412} /* (5, 28, 12) {real, imag} */,
  {32'hc04436a8, 32'h4133f885} /* (5, 28, 11) {real, imag} */,
  {32'h4182e245, 32'hc0cf4bec} /* (5, 28, 10) {real, imag} */,
  {32'hbec63460, 32'hc1b2a520} /* (5, 28, 9) {real, imag} */,
  {32'hc13f965c, 32'hc1d5db9c} /* (5, 28, 8) {real, imag} */,
  {32'hbfd4a940, 32'hbf308700} /* (5, 28, 7) {real, imag} */,
  {32'hc10ff796, 32'hc1ac9380} /* (5, 28, 6) {real, imag} */,
  {32'hc0853586, 32'hc108a08f} /* (5, 28, 5) {real, imag} */,
  {32'h3ff176e6, 32'h40e127d5} /* (5, 28, 4) {real, imag} */,
  {32'h408c7ecb, 32'h40fa499a} /* (5, 28, 3) {real, imag} */,
  {32'hc025b12c, 32'h401d3740} /* (5, 28, 2) {real, imag} */,
  {32'hc167f3c0, 32'hc03b5be8} /* (5, 28, 1) {real, imag} */,
  {32'hc1081b79, 32'h40529154} /* (5, 28, 0) {real, imag} */,
  {32'hc09f78d9, 32'h40659c12} /* (5, 27, 31) {real, imag} */,
  {32'hc1178b1a, 32'hbf06ae48} /* (5, 27, 30) {real, imag} */,
  {32'hc1a47bc4, 32'hc01f186e} /* (5, 27, 29) {real, imag} */,
  {32'hc1d3cde7, 32'h4188bc12} /* (5, 27, 28) {real, imag} */,
  {32'hc1539f46, 32'h411671ea} /* (5, 27, 27) {real, imag} */,
  {32'h40d30fb6, 32'hc108220d} /* (5, 27, 26) {real, imag} */,
  {32'h40ed371a, 32'hc1b122c3} /* (5, 27, 25) {real, imag} */,
  {32'h3ee0e700, 32'h408d251e} /* (5, 27, 24) {real, imag} */,
  {32'hc1b1e3e4, 32'hc05b37d9} /* (5, 27, 23) {real, imag} */,
  {32'hc1215c12, 32'hc0e9f384} /* (5, 27, 22) {real, imag} */,
  {32'hc0c7d0c6, 32'hbfdbf6d6} /* (5, 27, 21) {real, imag} */,
  {32'hbfa9f030, 32'hc0ef342a} /* (5, 27, 20) {real, imag} */,
  {32'h415f0b9c, 32'hc0bbf28c} /* (5, 27, 19) {real, imag} */,
  {32'h40d5e884, 32'hc0dd8a72} /* (5, 27, 18) {real, imag} */,
  {32'h408f2f7c, 32'hc12ffe05} /* (5, 27, 17) {real, imag} */,
  {32'h40defccb, 32'hc1464c4c} /* (5, 27, 16) {real, imag} */,
  {32'hbf01ddd0, 32'hc1b87c60} /* (5, 27, 15) {real, imag} */,
  {32'h411fe132, 32'hc1706f54} /* (5, 27, 14) {real, imag} */,
  {32'h40f91658, 32'hc10c6592} /* (5, 27, 13) {real, imag} */,
  {32'h40358dd5, 32'hc13eb972} /* (5, 27, 12) {real, imag} */,
  {32'hc13d048f, 32'hc13b01a4} /* (5, 27, 11) {real, imag} */,
  {32'hc0fe3f6c, 32'h40066ea4} /* (5, 27, 10) {real, imag} */,
  {32'hc0c603f7, 32'h41a348d6} /* (5, 27, 9) {real, imag} */,
  {32'hc18a9d78, 32'h420e6d82} /* (5, 27, 8) {real, imag} */,
  {32'hc1ac1bf7, 32'h41ae59be} /* (5, 27, 7) {real, imag} */,
  {32'h3f9a0660, 32'h41aad7b9} /* (5, 27, 6) {real, imag} */,
  {32'h410dbc2c, 32'h41fc95db} /* (5, 27, 5) {real, imag} */,
  {32'hbf921c30, 32'h419d4a1f} /* (5, 27, 4) {real, imag} */,
  {32'h3e6cfc80, 32'h41b6cd66} /* (5, 27, 3) {real, imag} */,
  {32'hc1075ed9, 32'h4132444f} /* (5, 27, 2) {real, imag} */,
  {32'hc10abdc0, 32'h4048458b} /* (5, 27, 1) {real, imag} */,
  {32'h40a0304e, 32'h3ff1d498} /* (5, 27, 0) {real, imag} */,
  {32'hc0fb51e0, 32'h4026ab8d} /* (5, 26, 31) {real, imag} */,
  {32'hc1aac4dc, 32'h41086ab5} /* (5, 26, 30) {real, imag} */,
  {32'hc1a9752f, 32'h407b102d} /* (5, 26, 29) {real, imag} */,
  {32'hbf12defc, 32'h417b4e5b} /* (5, 26, 28) {real, imag} */,
  {32'h41913bbb, 32'h41fcc08e} /* (5, 26, 27) {real, imag} */,
  {32'h414ca3e1, 32'h41421e12} /* (5, 26, 26) {real, imag} */,
  {32'hc0e44a3b, 32'h3f534ac0} /* (5, 26, 25) {real, imag} */,
  {32'hc102fe03, 32'hc12d1a2b} /* (5, 26, 24) {real, imag} */,
  {32'h414052c8, 32'h40db3011} /* (5, 26, 23) {real, imag} */,
  {32'h4064cb54, 32'hbdfc2a60} /* (5, 26, 22) {real, imag} */,
  {32'hbfd5a9ff, 32'hc135aeda} /* (5, 26, 21) {real, imag} */,
  {32'h41639221, 32'h3f81d9a6} /* (5, 26, 20) {real, imag} */,
  {32'h41aafc51, 32'h4170b4a5} /* (5, 26, 19) {real, imag} */,
  {32'h40253e0a, 32'h40e09865} /* (5, 26, 18) {real, imag} */,
  {32'h412fae5f, 32'hc03664f8} /* (5, 26, 17) {real, imag} */,
  {32'h41728942, 32'hc0dbbb27} /* (5, 26, 16) {real, imag} */,
  {32'h40e3f997, 32'hc03f13c0} /* (5, 26, 15) {real, imag} */,
  {32'h3ead96fd, 32'h4171b000} /* (5, 26, 14) {real, imag} */,
  {32'h40b2bf51, 32'hc10c92f6} /* (5, 26, 13) {real, imag} */,
  {32'h418da47c, 32'hc1655479} /* (5, 26, 12) {real, imag} */,
  {32'hc050426c, 32'h408cc60a} /* (5, 26, 11) {real, imag} */,
  {32'hc0bcd05e, 32'h4133df60} /* (5, 26, 10) {real, imag} */,
  {32'hc0ddb5b1, 32'h40d93c1a} /* (5, 26, 9) {real, imag} */,
  {32'h40ee7776, 32'h41884967} /* (5, 26, 8) {real, imag} */,
  {32'h413f96a6, 32'h413d6d00} /* (5, 26, 7) {real, imag} */,
  {32'h4147c0f8, 32'h409aa947} /* (5, 26, 6) {real, imag} */,
  {32'hc11f2a63, 32'h40094290} /* (5, 26, 5) {real, imag} */,
  {32'hc1a04c1b, 32'hc0b538b3} /* (5, 26, 4) {real, imag} */,
  {32'hc15fa2bc, 32'hc0e5fd45} /* (5, 26, 3) {real, imag} */,
  {32'hc106b745, 32'h41129ee2} /* (5, 26, 2) {real, imag} */,
  {32'hc0979d6a, 32'h4184cfd8} /* (5, 26, 1) {real, imag} */,
  {32'hbe9b353a, 32'h4187f398} /* (5, 26, 0) {real, imag} */,
  {32'h40fc9850, 32'h3c0fe000} /* (5, 25, 31) {real, imag} */,
  {32'h41556d78, 32'hc0f61c34} /* (5, 25, 30) {real, imag} */,
  {32'h40ed2f30, 32'h4085ad90} /* (5, 25, 29) {real, imag} */,
  {32'hc0c82619, 32'hc11ae010} /* (5, 25, 28) {real, imag} */,
  {32'hc0ef584b, 32'hc0f36416} /* (5, 25, 27) {real, imag} */,
  {32'hc16841ae, 32'hc10995da} /* (5, 25, 26) {real, imag} */,
  {32'h40094871, 32'hc13fcd6a} /* (5, 25, 25) {real, imag} */,
  {32'h3e5915b0, 32'hc084e575} /* (5, 25, 24) {real, imag} */,
  {32'hc0d632d0, 32'hc0f1eb2c} /* (5, 25, 23) {real, imag} */,
  {32'hc15c1614, 32'hc113531e} /* (5, 25, 22) {real, imag} */,
  {32'h4068dc31, 32'h3f4d5e18} /* (5, 25, 21) {real, imag} */,
  {32'h4156090f, 32'hc0211bdc} /* (5, 25, 20) {real, imag} */,
  {32'h41808af6, 32'hc11c106f} /* (5, 25, 19) {real, imag} */,
  {32'h4153304f, 32'h3f9f4468} /* (5, 25, 18) {real, imag} */,
  {32'h419708ef, 32'hbf710ef8} /* (5, 25, 17) {real, imag} */,
  {32'h40ebb52b, 32'hbf38d9e0} /* (5, 25, 16) {real, imag} */,
  {32'hc0ff3c96, 32'h40044a54} /* (5, 25, 15) {real, imag} */,
  {32'hc16db4ce, 32'h40bcce8f} /* (5, 25, 14) {real, imag} */,
  {32'hc0b95935, 32'hc0935811} /* (5, 25, 13) {real, imag} */,
  {32'hc0de7b7e, 32'h4081c2ed} /* (5, 25, 12) {real, imag} */,
  {32'h408cd85b, 32'hc0893d66} /* (5, 25, 11) {real, imag} */,
  {32'hc18a8fd0, 32'hc12b26f0} /* (5, 25, 10) {real, imag} */,
  {32'hc1406ec4, 32'hbfcb8906} /* (5, 25, 9) {real, imag} */,
  {32'hc0f64914, 32'hc0c13011} /* (5, 25, 8) {real, imag} */,
  {32'hc15e30a5, 32'hc10e06eb} /* (5, 25, 7) {real, imag} */,
  {32'hc1a03187, 32'hbe841e48} /* (5, 25, 6) {real, imag} */,
  {32'hc18b014e, 32'hc038efb5} /* (5, 25, 5) {real, imag} */,
  {32'hc13d2202, 32'h4077397d} /* (5, 25, 4) {real, imag} */,
  {32'h40bd19f3, 32'hc021d22e} /* (5, 25, 3) {real, imag} */,
  {32'hbee51fb0, 32'hc13b155a} /* (5, 25, 2) {real, imag} */,
  {32'h4090fd50, 32'h3fb57660} /* (5, 25, 1) {real, imag} */,
  {32'h412c3982, 32'h3c39c400} /* (5, 25, 0) {real, imag} */,
  {32'hc0c3294e, 32'hc1174ff6} /* (5, 24, 31) {real, imag} */,
  {32'h3fe6c554, 32'hc0bc73fd} /* (5, 24, 30) {real, imag} */,
  {32'h41025b9b, 32'h414add12} /* (5, 24, 29) {real, imag} */,
  {32'h40bcf251, 32'h4057dd71} /* (5, 24, 28) {real, imag} */,
  {32'h4132fa30, 32'h40ff323d} /* (5, 24, 27) {real, imag} */,
  {32'h4105197f, 32'h41d422aa} /* (5, 24, 26) {real, imag} */,
  {32'hbf7c0458, 32'h41a0304c} /* (5, 24, 25) {real, imag} */,
  {32'hc03112a6, 32'hbf9b233c} /* (5, 24, 24) {real, imag} */,
  {32'h3fd72c8a, 32'h405ddb1f} /* (5, 24, 23) {real, imag} */,
  {32'h3e258780, 32'h3ecb2e40} /* (5, 24, 22) {real, imag} */,
  {32'h413bdeec, 32'h4014aa54} /* (5, 24, 21) {real, imag} */,
  {32'h418ec457, 32'hc0c0799a} /* (5, 24, 20) {real, imag} */,
  {32'h40388777, 32'hc1426616} /* (5, 24, 19) {real, imag} */,
  {32'h40b37344, 32'hc190615c} /* (5, 24, 18) {real, imag} */,
  {32'h41424f26, 32'hc1843bd4} /* (5, 24, 17) {real, imag} */,
  {32'hc12a5d99, 32'hc0c3645d} /* (5, 24, 16) {real, imag} */,
  {32'hc153b26c, 32'h3fc163d4} /* (5, 24, 15) {real, imag} */,
  {32'hc15eaa9c, 32'h41801d4c} /* (5, 24, 14) {real, imag} */,
  {32'hc0b36b34, 32'h413dfb03} /* (5, 24, 13) {real, imag} */,
  {32'h41001c6f, 32'hc104e3a5} /* (5, 24, 12) {real, imag} */,
  {32'h413ac2d5, 32'hc025cb93} /* (5, 24, 11) {real, imag} */,
  {32'hc14c83f2, 32'h40e4db18} /* (5, 24, 10) {real, imag} */,
  {32'hc16ed099, 32'h3e4ac380} /* (5, 24, 9) {real, imag} */,
  {32'hc03682aa, 32'h40d15e53} /* (5, 24, 8) {real, imag} */,
  {32'hc0a61792, 32'h3f14cae0} /* (5, 24, 7) {real, imag} */,
  {32'hc1130c3e, 32'h40e1078a} /* (5, 24, 6) {real, imag} */,
  {32'hbfd1ed0c, 32'h41af30aa} /* (5, 24, 5) {real, imag} */,
  {32'hc0a10438, 32'h41566678} /* (5, 24, 4) {real, imag} */,
  {32'hc04d5c4c, 32'h40388aee} /* (5, 24, 3) {real, imag} */,
  {32'hbf2a90e8, 32'h415c6e1e} /* (5, 24, 2) {real, imag} */,
  {32'h41218876, 32'h4135dca3} /* (5, 24, 1) {real, imag} */,
  {32'h4098e437, 32'h408fc849} /* (5, 24, 0) {real, imag} */,
  {32'h406fb5d6, 32'hbff126f6} /* (5, 23, 31) {real, imag} */,
  {32'h3f844380, 32'hc09fba70} /* (5, 23, 30) {real, imag} */,
  {32'hbfe36066, 32'hc138daee} /* (5, 23, 29) {real, imag} */,
  {32'hc0a12519, 32'hc1536450} /* (5, 23, 28) {real, imag} */,
  {32'hc15480f0, 32'hc128c191} /* (5, 23, 27) {real, imag} */,
  {32'hc127ec08, 32'h409f5cbc} /* (5, 23, 26) {real, imag} */,
  {32'h408b73f0, 32'h4150ea98} /* (5, 23, 25) {real, imag} */,
  {32'h3f867a42, 32'h4149187a} /* (5, 23, 24) {real, imag} */,
  {32'h40484a17, 32'h410dc733} /* (5, 23, 23) {real, imag} */,
  {32'hbfff7a60, 32'h410e4528} /* (5, 23, 22) {real, imag} */,
  {32'hc0b393e7, 32'h3f92c214} /* (5, 23, 21) {real, imag} */,
  {32'h40858204, 32'h4103e46f} /* (5, 23, 20) {real, imag} */,
  {32'h411ceb2e, 32'h3fbef6ac} /* (5, 23, 19) {real, imag} */,
  {32'hc0ed3452, 32'hc13c0036} /* (5, 23, 18) {real, imag} */,
  {32'hc07d1668, 32'hc08ff051} /* (5, 23, 17) {real, imag} */,
  {32'hc14baecf, 32'h40d01bd5} /* (5, 23, 16) {real, imag} */,
  {32'hbf1a96e8, 32'hc047b343} /* (5, 23, 15) {real, imag} */,
  {32'h40ead64b, 32'hc13dd98e} /* (5, 23, 14) {real, imag} */,
  {32'h4176053a, 32'hc107c55c} /* (5, 23, 13) {real, imag} */,
  {32'h404b1ac8, 32'hc01e036e} /* (5, 23, 12) {real, imag} */,
  {32'h413da4de, 32'h41536561} /* (5, 23, 11) {real, imag} */,
  {32'hc00d4890, 32'h4041862e} /* (5, 23, 10) {real, imag} */,
  {32'hc13c1712, 32'h40f78226} /* (5, 23, 9) {real, imag} */,
  {32'hc157fe73, 32'hc0de333e} /* (5, 23, 8) {real, imag} */,
  {32'h3e1e5df0, 32'hc0f9d0fa} /* (5, 23, 7) {real, imag} */,
  {32'hbf27e0a0, 32'hbfbef568} /* (5, 23, 6) {real, imag} */,
  {32'h41727633, 32'h411f34e1} /* (5, 23, 5) {real, imag} */,
  {32'h40afab11, 32'h3fcadda6} /* (5, 23, 4) {real, imag} */,
  {32'h3fb33824, 32'hc166a6be} /* (5, 23, 3) {real, imag} */,
  {32'hc015d8c2, 32'hc0f96df8} /* (5, 23, 2) {real, imag} */,
  {32'hc10029c4, 32'h408f8b40} /* (5, 23, 1) {real, imag} */,
  {32'hbff39917, 32'h3f708d40} /* (5, 23, 0) {real, imag} */,
  {32'hc08033ff, 32'hc0c41e82} /* (5, 22, 31) {real, imag} */,
  {32'h4035d6a9, 32'hc0fe5894} /* (5, 22, 30) {real, imag} */,
  {32'h400023f0, 32'hc119ac8b} /* (5, 22, 29) {real, imag} */,
  {32'hbf8664a6, 32'hbf4d587c} /* (5, 22, 28) {real, imag} */,
  {32'h404231c5, 32'h40d9b1da} /* (5, 22, 27) {real, imag} */,
  {32'h3f702680, 32'h404f033f} /* (5, 22, 26) {real, imag} */,
  {32'h406c78af, 32'hc00046b8} /* (5, 22, 25) {real, imag} */,
  {32'hc0b0bbf0, 32'hc023d564} /* (5, 22, 24) {real, imag} */,
  {32'h3fa6d6e0, 32'h3efb5560} /* (5, 22, 23) {real, imag} */,
  {32'h3fd83250, 32'h40256a1f} /* (5, 22, 22) {real, imag} */,
  {32'hc0708d44, 32'hbfb4abbc} /* (5, 22, 21) {real, imag} */,
  {32'hc0d58a10, 32'h40e01a60} /* (5, 22, 20) {real, imag} */,
  {32'h406f2a04, 32'h4120da4e} /* (5, 22, 19) {real, imag} */,
  {32'h41200505, 32'h40503ae1} /* (5, 22, 18) {real, imag} */,
  {32'hbe25c240, 32'h415be671} /* (5, 22, 17) {real, imag} */,
  {32'hc143507a, 32'h41178282} /* (5, 22, 16) {real, imag} */,
  {32'hc09f723e, 32'hbfdf73ea} /* (5, 22, 15) {real, imag} */,
  {32'hbfb4632b, 32'h3fa1f49e} /* (5, 22, 14) {real, imag} */,
  {32'h401f1672, 32'h3f974754} /* (5, 22, 13) {real, imag} */,
  {32'hc0963115, 32'hc0c79e57} /* (5, 22, 12) {real, imag} */,
  {32'hc1bd76f8, 32'hc103039c} /* (5, 22, 11) {real, imag} */,
  {32'hc1360576, 32'hc1812e8e} /* (5, 22, 10) {real, imag} */,
  {32'h40b23de7, 32'hc1492b45} /* (5, 22, 9) {real, imag} */,
  {32'h40f913fe, 32'hc13f9830} /* (5, 22, 8) {real, imag} */,
  {32'h40a1e8f5, 32'hc10b3285} /* (5, 22, 7) {real, imag} */,
  {32'h411e8fc6, 32'hc10ff623} /* (5, 22, 6) {real, imag} */,
  {32'h3fdcf36a, 32'hc1205a33} /* (5, 22, 5) {real, imag} */,
  {32'h3f9fd6e4, 32'hc04051e2} /* (5, 22, 4) {real, imag} */,
  {32'hc0e135e8, 32'hbfdf2cdd} /* (5, 22, 3) {real, imag} */,
  {32'hc15207d6, 32'hbffa2b2c} /* (5, 22, 2) {real, imag} */,
  {32'hc10bd86a, 32'hbfdce8e6} /* (5, 22, 1) {real, imag} */,
  {32'hc06353bc, 32'hc061e481} /* (5, 22, 0) {real, imag} */,
  {32'hc01290f4, 32'h40fe3b8a} /* (5, 21, 31) {real, imag} */,
  {32'h4099174c, 32'h416342c4} /* (5, 21, 30) {real, imag} */,
  {32'h3fdee278, 32'h41047d30} /* (5, 21, 29) {real, imag} */,
  {32'hc072cd9e, 32'h40768f61} /* (5, 21, 28) {real, imag} */,
  {32'h40c7fbbf, 32'hbfdf6bd4} /* (5, 21, 27) {real, imag} */,
  {32'h4042b050, 32'hc0351833} /* (5, 21, 26) {real, imag} */,
  {32'h3f108810, 32'hc06c1084} /* (5, 21, 25) {real, imag} */,
  {32'hbd3cf100, 32'h3f49f710} /* (5, 21, 24) {real, imag} */,
  {32'h4113e1e1, 32'h41193f92} /* (5, 21, 23) {real, imag} */,
  {32'h41445c9a, 32'h415d0454} /* (5, 21, 22) {real, imag} */,
  {32'h4129eb4e, 32'h3ee99ba0} /* (5, 21, 21) {real, imag} */,
  {32'hc00a93fe, 32'hbf20143c} /* (5, 21, 20) {real, imag} */,
  {32'hc13123ed, 32'hc03c92e8} /* (5, 21, 19) {real, imag} */,
  {32'hbee47f60, 32'hbf89d670} /* (5, 21, 18) {real, imag} */,
  {32'hbe2b4b40, 32'h3fea777e} /* (5, 21, 17) {real, imag} */,
  {32'hbfbbb700, 32'h3f1f5a30} /* (5, 21, 16) {real, imag} */,
  {32'h404ff841, 32'h40bd2f56} /* (5, 21, 15) {real, imag} */,
  {32'h3ff96a33, 32'h41221152} /* (5, 21, 14) {real, imag} */,
  {32'hc0960448, 32'h3fbdad71} /* (5, 21, 13) {real, imag} */,
  {32'hc04c6a9f, 32'hc0b83bf3} /* (5, 21, 12) {real, imag} */,
  {32'hc0cffd5a, 32'hc1353a44} /* (5, 21, 11) {real, imag} */,
  {32'hc055981a, 32'h4087926d} /* (5, 21, 10) {real, imag} */,
  {32'h404363ce, 32'h3f26b868} /* (5, 21, 9) {real, imag} */,
  {32'h41020c58, 32'h40737862} /* (5, 21, 8) {real, imag} */,
  {32'h403180ee, 32'hbf3e9e38} /* (5, 21, 7) {real, imag} */,
  {32'hc100db5c, 32'h4007cc06} /* (5, 21, 6) {real, imag} */,
  {32'hc0b580d5, 32'h405a2254} /* (5, 21, 5) {real, imag} */,
  {32'h3ff92c4d, 32'h403a47a0} /* (5, 21, 4) {real, imag} */,
  {32'hc0093dbf, 32'h40bfe248} /* (5, 21, 3) {real, imag} */,
  {32'h3e587d50, 32'hc01e14bb} /* (5, 21, 2) {real, imag} */,
  {32'h41036968, 32'h40fedc82} /* (5, 21, 1) {real, imag} */,
  {32'h40073ebc, 32'h4139605e} /* (5, 21, 0) {real, imag} */,
  {32'h4088ab45, 32'hc0b15f85} /* (5, 20, 31) {real, imag} */,
  {32'h40dc506c, 32'h3f252640} /* (5, 20, 30) {real, imag} */,
  {32'h4132269c, 32'h3f1fb110} /* (5, 20, 29) {real, imag} */,
  {32'h41142009, 32'hc027ea36} /* (5, 20, 28) {real, imag} */,
  {32'hbf9abdec, 32'hbf331814} /* (5, 20, 27) {real, imag} */,
  {32'hc0b69d8a, 32'hc116f1ae} /* (5, 20, 26) {real, imag} */,
  {32'hc0148d78, 32'hc0ddf480} /* (5, 20, 25) {real, imag} */,
  {32'h40a04122, 32'h407185ad} /* (5, 20, 24) {real, imag} */,
  {32'h3fabdeca, 32'h411189f9} /* (5, 20, 23) {real, imag} */,
  {32'h4037c769, 32'h413809c1} /* (5, 20, 22) {real, imag} */,
  {32'h403ee13c, 32'h40c43e26} /* (5, 20, 21) {real, imag} */,
  {32'hbf159f10, 32'hc09ff11c} /* (5, 20, 20) {real, imag} */,
  {32'hc0279578, 32'hc0d33458} /* (5, 20, 19) {real, imag} */,
  {32'hc0821f08, 32'hc0aae1f9} /* (5, 20, 18) {real, imag} */,
  {32'hc09a7927, 32'hc0aa9b73} /* (5, 20, 17) {real, imag} */,
  {32'hbf013170, 32'h411590c6} /* (5, 20, 16) {real, imag} */,
  {32'h404fca66, 32'h40d8eaf8} /* (5, 20, 15) {real, imag} */,
  {32'h40947c96, 32'h3eb105a0} /* (5, 20, 14) {real, imag} */,
  {32'hbf898480, 32'h3f734640} /* (5, 20, 13) {real, imag} */,
  {32'hbfdf4608, 32'h40e9e643} /* (5, 20, 12) {real, imag} */,
  {32'h4059aed2, 32'h4021138d} /* (5, 20, 11) {real, imag} */,
  {32'h40048518, 32'hc0d35f68} /* (5, 20, 10) {real, imag} */,
  {32'h3fe411a4, 32'hc0b3c140} /* (5, 20, 9) {real, imag} */,
  {32'hbef397b0, 32'h4036dea6} /* (5, 20, 8) {real, imag} */,
  {32'hc00e261b, 32'h3eab2368} /* (5, 20, 7) {real, imag} */,
  {32'h40b0e72f, 32'hbfe8fd44} /* (5, 20, 6) {real, imag} */,
  {32'h3ff88170, 32'hc00c9b44} /* (5, 20, 5) {real, imag} */,
  {32'h4049df7e, 32'hc0c4e0ca} /* (5, 20, 4) {real, imag} */,
  {32'h407435e2, 32'hc1026dfc} /* (5, 20, 3) {real, imag} */,
  {32'hbff4a452, 32'h400bf4f9} /* (5, 20, 2) {real, imag} */,
  {32'h3f971b62, 32'hbf92ac94} /* (5, 20, 1) {real, imag} */,
  {32'h3f9fc666, 32'hc112f990} /* (5, 20, 0) {real, imag} */,
  {32'h3f8b10c9, 32'h4008e2bd} /* (5, 19, 31) {real, imag} */,
  {32'hbfd75292, 32'h3f4ab0f4} /* (5, 19, 30) {real, imag} */,
  {32'h3e96d5f0, 32'hc095d00e} /* (5, 19, 29) {real, imag} */,
  {32'h3e595a00, 32'hc03938f8} /* (5, 19, 28) {real, imag} */,
  {32'hbfd42042, 32'h3fba01d0} /* (5, 19, 27) {real, imag} */,
  {32'hbf4b7cb8, 32'hbf3edbb8} /* (5, 19, 26) {real, imag} */,
  {32'hc0dad8ce, 32'hbe90ede0} /* (5, 19, 25) {real, imag} */,
  {32'hc04738bd, 32'hbfede9c0} /* (5, 19, 24) {real, imag} */,
  {32'hbe78fbd0, 32'h3f5b4f70} /* (5, 19, 23) {real, imag} */,
  {32'h3f0d6e6c, 32'hc05c3af2} /* (5, 19, 22) {real, imag} */,
  {32'hc0c5e9c2, 32'hc0eb0a31} /* (5, 19, 21) {real, imag} */,
  {32'hc03d8296, 32'hc09fc72e} /* (5, 19, 20) {real, imag} */,
  {32'hc0b618c4, 32'h3e89b5f0} /* (5, 19, 19) {real, imag} */,
  {32'h400a15c4, 32'h407b2f25} /* (5, 19, 18) {real, imag} */,
  {32'h40e282bb, 32'h41458468} /* (5, 19, 17) {real, imag} */,
  {32'h4008dd7e, 32'h406f7814} /* (5, 19, 16) {real, imag} */,
  {32'hc0b108ff, 32'hc0dcd4ba} /* (5, 19, 15) {real, imag} */,
  {32'hbf45033a, 32'hc0b22a42} /* (5, 19, 14) {real, imag} */,
  {32'hbd0db1a0, 32'hbfadea93} /* (5, 19, 13) {real, imag} */,
  {32'hc103dd01, 32'h4035cd20} /* (5, 19, 12) {real, imag} */,
  {32'hc12da7e2, 32'h4103f41d} /* (5, 19, 11) {real, imag} */,
  {32'hc0040d6d, 32'h40beba15} /* (5, 19, 10) {real, imag} */,
  {32'hbed64310, 32'hc01caa78} /* (5, 19, 9) {real, imag} */,
  {32'hc000ea44, 32'hbf9e890f} /* (5, 19, 8) {real, imag} */,
  {32'h3fbcacb2, 32'hbe54f1c0} /* (5, 19, 7) {real, imag} */,
  {32'h3f7743f0, 32'hc04670e8} /* (5, 19, 6) {real, imag} */,
  {32'h3e909408, 32'h3feac2d6} /* (5, 19, 5) {real, imag} */,
  {32'h3fd17b1e, 32'h3f204ce2} /* (5, 19, 4) {real, imag} */,
  {32'h407bbeff, 32'h40a0787d} /* (5, 19, 3) {real, imag} */,
  {32'h3e8b56c8, 32'h4031b9f1} /* (5, 19, 2) {real, imag} */,
  {32'hc0be81ae, 32'hc0df391b} /* (5, 19, 1) {real, imag} */,
  {32'hc010ab34, 32'hc0015970} /* (5, 19, 0) {real, imag} */,
  {32'hbfbc5bc2, 32'h403bbe8a} /* (5, 18, 31) {real, imag} */,
  {32'hc0841418, 32'h4040640a} /* (5, 18, 30) {real, imag} */,
  {32'hbfc0c056, 32'h40dc17aa} /* (5, 18, 29) {real, imag} */,
  {32'hbe750620, 32'h40f39df0} /* (5, 18, 28) {real, imag} */,
  {32'h3fc85ed8, 32'h3fc79b24} /* (5, 18, 27) {real, imag} */,
  {32'h4006cd35, 32'h400d03e0} /* (5, 18, 26) {real, imag} */,
  {32'h3f07c7be, 32'h4009540e} /* (5, 18, 25) {real, imag} */,
  {32'hc03224a1, 32'hc0aa8759} /* (5, 18, 24) {real, imag} */,
  {32'h40591509, 32'hc023f1bf} /* (5, 18, 23) {real, imag} */,
  {32'h40eea280, 32'hbfd57328} /* (5, 18, 22) {real, imag} */,
  {32'h40def359, 32'hc097c620} /* (5, 18, 21) {real, imag} */,
  {32'h40b5bfde, 32'hc01f32e8} /* (5, 18, 20) {real, imag} */,
  {32'h4123d5e8, 32'h3d513a80} /* (5, 18, 19) {real, imag} */,
  {32'h40bea684, 32'h4087ba4e} /* (5, 18, 18) {real, imag} */,
  {32'h3fa2d428, 32'h401da808} /* (5, 18, 17) {real, imag} */,
  {32'hbf7664f0, 32'hbe9cd330} /* (5, 18, 16) {real, imag} */,
  {32'hc023bca6, 32'h3ee0bad0} /* (5, 18, 15) {real, imag} */,
  {32'hc149b77f, 32'hc01a8392} /* (5, 18, 14) {real, imag} */,
  {32'hc0dbc33f, 32'h3f0752b2} /* (5, 18, 13) {real, imag} */,
  {32'h3d2ad500, 32'h4103936e} /* (5, 18, 12) {real, imag} */,
  {32'hc0204570, 32'hbf4c1dbc} /* (5, 18, 11) {real, imag} */,
  {32'hbf122cc8, 32'hc0f8d8ce} /* (5, 18, 10) {real, imag} */,
  {32'hc032a85e, 32'hc056b1e2} /* (5, 18, 9) {real, imag} */,
  {32'hc079f3b4, 32'hbe8617f0} /* (5, 18, 8) {real, imag} */,
  {32'hbfff51fa, 32'h4010e5de} /* (5, 18, 7) {real, imag} */,
  {32'h40c8b622, 32'h3f669a02} /* (5, 18, 6) {real, imag} */,
  {32'hbfc2df44, 32'h3feaa07e} /* (5, 18, 5) {real, imag} */,
  {32'hc0e1c266, 32'h4108d6b6} /* (5, 18, 4) {real, imag} */,
  {32'h402fa4b5, 32'h40b1740c} /* (5, 18, 3) {real, imag} */,
  {32'h405c4b13, 32'h3d34dd80} /* (5, 18, 2) {real, imag} */,
  {32'hbeb8a890, 32'hc0253766} /* (5, 18, 1) {real, imag} */,
  {32'h4031cdd9, 32'hc04e78f0} /* (5, 18, 0) {real, imag} */,
  {32'hbeeb03e0, 32'h3fe2ba76} /* (5, 17, 31) {real, imag} */,
  {32'hbfd198a8, 32'hbffd1c00} /* (5, 17, 30) {real, imag} */,
  {32'h3f7b2384, 32'hc049113a} /* (5, 17, 29) {real, imag} */,
  {32'h3f49d79c, 32'hbffb9e00} /* (5, 17, 28) {real, imag} */,
  {32'h3fbfb1b0, 32'h3fea3240} /* (5, 17, 27) {real, imag} */,
  {32'h40a6086e, 32'h3d1f6da0} /* (5, 17, 26) {real, imag} */,
  {32'h40a6e17a, 32'h4019c9fe} /* (5, 17, 25) {real, imag} */,
  {32'h401f871d, 32'h3fa874fe} /* (5, 17, 24) {real, imag} */,
  {32'hc00d4804, 32'h3f0ecc98} /* (5, 17, 23) {real, imag} */,
  {32'hbfe5b9dc, 32'h402a8204} /* (5, 17, 22) {real, imag} */,
  {32'hc01040ce, 32'h3f8f809e} /* (5, 17, 21) {real, imag} */,
  {32'h40b27510, 32'hbf00d672} /* (5, 17, 20) {real, imag} */,
  {32'h4098981e, 32'h404aaa52} /* (5, 17, 19) {real, imag} */,
  {32'h3eed5320, 32'h4084b8ba} /* (5, 17, 18) {real, imag} */,
  {32'h3d4d0ec0, 32'h401279d3} /* (5, 17, 17) {real, imag} */,
  {32'hbea7bd98, 32'h4057c3dc} /* (5, 17, 16) {real, imag} */,
  {32'hbe7f8d00, 32'hbfc64846} /* (5, 17, 15) {real, imag} */,
  {32'hbf9bf78c, 32'hc0d78665} /* (5, 17, 14) {real, imag} */,
  {32'h3fd4e497, 32'hc080bfeb} /* (5, 17, 13) {real, imag} */,
  {32'h40f4d798, 32'h3f62eaa0} /* (5, 17, 12) {real, imag} */,
  {32'h403178ea, 32'h40a7ded1} /* (5, 17, 11) {real, imag} */,
  {32'hc08990fe, 32'h401a76f2} /* (5, 17, 10) {real, imag} */,
  {32'hc03e0da4, 32'hc0387ee2} /* (5, 17, 9) {real, imag} */,
  {32'h3fee99ce, 32'hc0b87529} /* (5, 17, 8) {real, imag} */,
  {32'hbf88bb26, 32'hbef5af20} /* (5, 17, 7) {real, imag} */,
  {32'hbf9be39c, 32'hbeb8ac60} /* (5, 17, 6) {real, imag} */,
  {32'hc09ecb22, 32'h3f31e0a0} /* (5, 17, 5) {real, imag} */,
  {32'hc0a86a08, 32'hc05e00b2} /* (5, 17, 4) {real, imag} */,
  {32'hc09cf359, 32'hc084c91b} /* (5, 17, 3) {real, imag} */,
  {32'hbde0f300, 32'hc01a814c} /* (5, 17, 2) {real, imag} */,
  {32'hc0120f77, 32'hc086d109} /* (5, 17, 1) {real, imag} */,
  {32'hc04311d0, 32'h3dfc7f60} /* (5, 17, 0) {real, imag} */,
  {32'hbf9d8448, 32'h3f04b880} /* (5, 16, 31) {real, imag} */,
  {32'hc0139934, 32'h3ff06d30} /* (5, 16, 30) {real, imag} */,
  {32'h3f85d7d6, 32'hbf8b6330} /* (5, 16, 29) {real, imag} */,
  {32'h404de2c6, 32'h3fd05ed0} /* (5, 16, 28) {real, imag} */,
  {32'hbeaea800, 32'h4080606c} /* (5, 16, 27) {real, imag} */,
  {32'h3ee4d6a0, 32'hbfb5a2a0} /* (5, 16, 26) {real, imag} */,
  {32'h3fb10334, 32'h40e3cf0a} /* (5, 16, 25) {real, imag} */,
  {32'hbfb9ab98, 32'h401d38e0} /* (5, 16, 24) {real, imag} */,
  {32'hc012de15, 32'hc0344c04} /* (5, 16, 23) {real, imag} */,
  {32'hbd4fd2c0, 32'hbfa66a18} /* (5, 16, 22) {real, imag} */,
  {32'h4065993a, 32'h3e77af00} /* (5, 16, 21) {real, imag} */,
  {32'h40856720, 32'hbfd00d2c} /* (5, 16, 20) {real, imag} */,
  {32'h4003e0a1, 32'hbce50400} /* (5, 16, 19) {real, imag} */,
  {32'h4086beb2, 32'h3f3b1308} /* (5, 16, 18) {real, imag} */,
  {32'h40a56cdc, 32'hc041e060} /* (5, 16, 17) {real, imag} */,
  {32'hbff23698, 32'hbfdc8f14} /* (5, 16, 16) {real, imag} */,
  {32'hc071ba7a, 32'hbf16c930} /* (5, 16, 15) {real, imag} */,
  {32'hbf7ea600, 32'hc00ae93c} /* (5, 16, 14) {real, imag} */,
  {32'h3ed11f80, 32'hc008b6bc} /* (5, 16, 13) {real, imag} */,
  {32'hc00e45f4, 32'hbfa1ad38} /* (5, 16, 12) {real, imag} */,
  {32'hbff5aae8, 32'h3fa970d8} /* (5, 16, 11) {real, imag} */,
  {32'h3fd12ee0, 32'hc00f4025} /* (5, 16, 10) {real, imag} */,
  {32'h40e36954, 32'h3f90c9ea} /* (5, 16, 9) {real, imag} */,
  {32'h40037454, 32'h402dc3d5} /* (5, 16, 8) {real, imag} */,
  {32'h3f8eac04, 32'hbfaae67a} /* (5, 16, 7) {real, imag} */,
  {32'h3ea9fdc8, 32'hc005b044} /* (5, 16, 6) {real, imag} */,
  {32'hbf94fb90, 32'hbede6080} /* (5, 16, 5) {real, imag} */,
  {32'h3f9f37a0, 32'h3d194400} /* (5, 16, 4) {real, imag} */,
  {32'hbf7cc1ce, 32'hbf821670} /* (5, 16, 3) {real, imag} */,
  {32'hc00c5a4c, 32'hc077deba} /* (5, 16, 2) {real, imag} */,
  {32'h3ed93120, 32'h4069be40} /* (5, 16, 1) {real, imag} */,
  {32'hbf78424e, 32'h403527c8} /* (5, 16, 0) {real, imag} */,
  {32'hbec8eb80, 32'h3e816a46} /* (5, 15, 31) {real, imag} */,
  {32'h3f6c7870, 32'h402077d8} /* (5, 15, 30) {real, imag} */,
  {32'h40ae12d4, 32'h400d09ea} /* (5, 15, 29) {real, imag} */,
  {32'hc01b489b, 32'h4085b510} /* (5, 15, 28) {real, imag} */,
  {32'hbf811ff0, 32'h4049f8a0} /* (5, 15, 27) {real, imag} */,
  {32'h409c39ce, 32'h3fbe5773} /* (5, 15, 26) {real, imag} */,
  {32'h3e70ebc0, 32'hbf93e39b} /* (5, 15, 25) {real, imag} */,
  {32'hbe924368, 32'hbfc44bbe} /* (5, 15, 24) {real, imag} */,
  {32'h40fd7052, 32'hc02e2886} /* (5, 15, 23) {real, imag} */,
  {32'h40fc79df, 32'hc0713f24} /* (5, 15, 22) {real, imag} */,
  {32'h409876f3, 32'h3fbed2b2} /* (5, 15, 21) {real, imag} */,
  {32'h3fa1c736, 32'h408a6784} /* (5, 15, 20) {real, imag} */,
  {32'h4043ea9c, 32'h4034254e} /* (5, 15, 19) {real, imag} */,
  {32'h401ca15c, 32'h40684c9d} /* (5, 15, 18) {real, imag} */,
  {32'h40a0e69a, 32'h3fad7842} /* (5, 15, 17) {real, imag} */,
  {32'h3f223d54, 32'h40973c56} /* (5, 15, 16) {real, imag} */,
  {32'hbf4d8120, 32'h40862dfe} /* (5, 15, 15) {real, imag} */,
  {32'hbf45de88, 32'h40c605d1} /* (5, 15, 14) {real, imag} */,
  {32'hbf169b9e, 32'h40831163} /* (5, 15, 13) {real, imag} */,
  {32'hc0b9bfc0, 32'h40020d18} /* (5, 15, 12) {real, imag} */,
  {32'hbfade3c4, 32'h402fc91e} /* (5, 15, 11) {real, imag} */,
  {32'h40356e23, 32'h40a2fd08} /* (5, 15, 10) {real, imag} */,
  {32'hbf764410, 32'h3ecafcf0} /* (5, 15, 9) {real, imag} */,
  {32'hbf0730e4, 32'h406780f6} /* (5, 15, 8) {real, imag} */,
  {32'h40cb0e10, 32'h403f6824} /* (5, 15, 7) {real, imag} */,
  {32'h40dfdb47, 32'h405377ac} /* (5, 15, 6) {real, imag} */,
  {32'h3fcaafc6, 32'h3fc51cb0} /* (5, 15, 5) {real, imag} */,
  {32'h407b23c0, 32'hbf106618} /* (5, 15, 4) {real, imag} */,
  {32'h408d58e9, 32'h406ba48e} /* (5, 15, 3) {real, imag} */,
  {32'h40c0be88, 32'h40c28dd6} /* (5, 15, 2) {real, imag} */,
  {32'h3f3a27fc, 32'h40c4fb71} /* (5, 15, 1) {real, imag} */,
  {32'hbf96eb90, 32'h40ca7b7e} /* (5, 15, 0) {real, imag} */,
  {32'hbf0af864, 32'hbf90e294} /* (5, 14, 31) {real, imag} */,
  {32'h403a74ad, 32'hc0aeda65} /* (5, 14, 30) {real, imag} */,
  {32'h3f4c23d5, 32'h3f97a9b8} /* (5, 14, 29) {real, imag} */,
  {32'hc006d94a, 32'h405ace28} /* (5, 14, 28) {real, imag} */,
  {32'h3f4580f0, 32'hc0351102} /* (5, 14, 27) {real, imag} */,
  {32'hbfc16636, 32'hbf52c480} /* (5, 14, 26) {real, imag} */,
  {32'hbf9734f7, 32'h40832385} /* (5, 14, 25) {real, imag} */,
  {32'h3ec9a7a8, 32'hc0191f7e} /* (5, 14, 24) {real, imag} */,
  {32'hbfc74372, 32'h3da47fe0} /* (5, 14, 23) {real, imag} */,
  {32'hbec76980, 32'h40f8f7b2} /* (5, 14, 22) {real, imag} */,
  {32'h3fddaf04, 32'h40a708a0} /* (5, 14, 21) {real, imag} */,
  {32'hbe70c4c0, 32'h40e2d782} /* (5, 14, 20) {real, imag} */,
  {32'h403f6d0e, 32'hbda7c340} /* (5, 14, 19) {real, imag} */,
  {32'h40b33c36, 32'hc01b0f1c} /* (5, 14, 18) {real, imag} */,
  {32'h40ccfe66, 32'h40472b38} /* (5, 14, 17) {real, imag} */,
  {32'h40c5d5c2, 32'h3dc3b4c0} /* (5, 14, 16) {real, imag} */,
  {32'h402d797e, 32'hbfe9cef4} /* (5, 14, 15) {real, imag} */,
  {32'h3fc3af48, 32'h40a303ad} /* (5, 14, 14) {real, imag} */,
  {32'h407ff45e, 32'h3f48a06e} /* (5, 14, 13) {real, imag} */,
  {32'h41013ce5, 32'hc01bbefa} /* (5, 14, 12) {real, imag} */,
  {32'h40956be8, 32'hc02972d5} /* (5, 14, 11) {real, imag} */,
  {32'h3f3e2058, 32'hbf02bf8c} /* (5, 14, 10) {real, imag} */,
  {32'hc07bfcc6, 32'hc11c9ebc} /* (5, 14, 9) {real, imag} */,
  {32'hc03fe5dc, 32'hc032ae52} /* (5, 14, 8) {real, imag} */,
  {32'hc06677cf, 32'h4021091a} /* (5, 14, 7) {real, imag} */,
  {32'hc0c163c4, 32'h40882c10} /* (5, 14, 6) {real, imag} */,
  {32'hc0814ca3, 32'h3f276504} /* (5, 14, 5) {real, imag} */,
  {32'h4088db4e, 32'h3fc8888c} /* (5, 14, 4) {real, imag} */,
  {32'h40ee4f14, 32'h3f8df928} /* (5, 14, 3) {real, imag} */,
  {32'h40047b59, 32'h409d8eed} /* (5, 14, 2) {real, imag} */,
  {32'hc1082fdc, 32'h412bcf02} /* (5, 14, 1) {real, imag} */,
  {32'hc0b2c9a6, 32'h408511e4} /* (5, 14, 0) {real, imag} */,
  {32'h3ff83731, 32'h3f0ffa5c} /* (5, 13, 31) {real, imag} */,
  {32'h3ecca4e8, 32'h402a75ab} /* (5, 13, 30) {real, imag} */,
  {32'hc09ba781, 32'h407d2bfc} /* (5, 13, 29) {real, imag} */,
  {32'hc0872e98, 32'hc014c168} /* (5, 13, 28) {real, imag} */,
  {32'hc0d26ece, 32'h3fed9950} /* (5, 13, 27) {real, imag} */,
  {32'hc06b1c54, 32'h410d4016} /* (5, 13, 26) {real, imag} */,
  {32'hc0c22148, 32'hbf7fe3b0} /* (5, 13, 25) {real, imag} */,
  {32'h402e5d83, 32'hc05035b0} /* (5, 13, 24) {real, imag} */,
  {32'h40d2c282, 32'hbe66d600} /* (5, 13, 23) {real, imag} */,
  {32'h402f24ad, 32'h40c24def} /* (5, 13, 22) {real, imag} */,
  {32'h410692cc, 32'h41230902} /* (5, 13, 21) {real, imag} */,
  {32'h40449fb2, 32'h40919568} /* (5, 13, 20) {real, imag} */,
  {32'h3ef151c8, 32'h4069d206} /* (5, 13, 19) {real, imag} */,
  {32'hc04cfadc, 32'hc00e11b5} /* (5, 13, 18) {real, imag} */,
  {32'h40041af6, 32'hc03cb2e2} /* (5, 13, 17) {real, imag} */,
  {32'hc00754da, 32'h40457eda} /* (5, 13, 16) {real, imag} */,
  {32'hc10ca380, 32'h40f0aa2a} /* (5, 13, 15) {real, imag} */,
  {32'hc03dcb06, 32'hbf191910} /* (5, 13, 14) {real, imag} */,
  {32'h400a30b0, 32'hbf13aac6} /* (5, 13, 13) {real, imag} */,
  {32'hc08a2caa, 32'h3e5171c0} /* (5, 13, 12) {real, imag} */,
  {32'hc0d5eb75, 32'hbffe4b28} /* (5, 13, 11) {real, imag} */,
  {32'h40278f4b, 32'h4078ef3a} /* (5, 13, 10) {real, imag} */,
  {32'hc011faea, 32'h40c78e58} /* (5, 13, 9) {real, imag} */,
  {32'hc0703102, 32'hbe765678} /* (5, 13, 8) {real, imag} */,
  {32'hc0a94a3e, 32'hc05770fc} /* (5, 13, 7) {real, imag} */,
  {32'hc0e7a254, 32'h3eea4140} /* (5, 13, 6) {real, imag} */,
  {32'hc04206c9, 32'hc00860ab} /* (5, 13, 5) {real, imag} */,
  {32'h3e8ca8f8, 32'hbf80a7d1} /* (5, 13, 4) {real, imag} */,
  {32'hc000359f, 32'h402ebe5a} /* (5, 13, 3) {real, imag} */,
  {32'hc0e909c6, 32'h406520dd} /* (5, 13, 2) {real, imag} */,
  {32'hbcb01e00, 32'h402a5bb2} /* (5, 13, 1) {real, imag} */,
  {32'h40617304, 32'h3ec16c00} /* (5, 13, 0) {real, imag} */,
  {32'hbeb30594, 32'hc029cd5e} /* (5, 12, 31) {real, imag} */,
  {32'hc01c9a98, 32'hc0c5bf42} /* (5, 12, 30) {real, imag} */,
  {32'h406fad2c, 32'hc0972b32} /* (5, 12, 29) {real, imag} */,
  {32'h417c3519, 32'h3fd603c4} /* (5, 12, 28) {real, imag} */,
  {32'h410d0c02, 32'hbfe3abae} /* (5, 12, 27) {real, imag} */,
  {32'h3dff0880, 32'hc084cd3d} /* (5, 12, 26) {real, imag} */,
  {32'h405ba088, 32'hc0d73066} /* (5, 12, 25) {real, imag} */,
  {32'h3ff22eea, 32'hbfadfbce} /* (5, 12, 24) {real, imag} */,
  {32'hbeb63c58, 32'h4047047c} /* (5, 12, 23) {real, imag} */,
  {32'h3f1da2c0, 32'hc0c1190a} /* (5, 12, 22) {real, imag} */,
  {32'hbf4f91c2, 32'hc092f518} /* (5, 12, 21) {real, imag} */,
  {32'h40a15dda, 32'hbe1c3980} /* (5, 12, 20) {real, imag} */,
  {32'h3f4f2900, 32'h4012eb40} /* (5, 12, 19) {real, imag} */,
  {32'h3f9f3fb0, 32'hc0382a8e} /* (5, 12, 18) {real, imag} */,
  {32'hbfb2cc94, 32'hbebc1910} /* (5, 12, 17) {real, imag} */,
  {32'hc09ecade, 32'h3ea6a300} /* (5, 12, 16) {real, imag} */,
  {32'hc0351720, 32'h3e821c40} /* (5, 12, 15) {real, imag} */,
  {32'h40bc8c54, 32'h3e7ce740} /* (5, 12, 14) {real, imag} */,
  {32'h41219d79, 32'hbf91b5c0} /* (5, 12, 13) {real, imag} */,
  {32'hbe43f240, 32'hbf7c3fc8} /* (5, 12, 12) {real, imag} */,
  {32'h3fea5559, 32'h4095a1ee} /* (5, 12, 11) {real, imag} */,
  {32'hbf04aebe, 32'h406412d0} /* (5, 12, 10) {real, imag} */,
  {32'h4083d993, 32'hbf4a1d80} /* (5, 12, 9) {real, imag} */,
  {32'h41291800, 32'hbfdf6224} /* (5, 12, 8) {real, imag} */,
  {32'h40ee5a1a, 32'hc0015bf3} /* (5, 12, 7) {real, imag} */,
  {32'hbf42cac8, 32'hbf51ff98} /* (5, 12, 6) {real, imag} */,
  {32'hbfa6f500, 32'h4105ef31} /* (5, 12, 5) {real, imag} */,
  {32'hbfaaa90c, 32'h40dd2b1c} /* (5, 12, 4) {real, imag} */,
  {32'hc03a2784, 32'hbfaa2938} /* (5, 12, 3) {real, imag} */,
  {32'hbf98dc62, 32'hc00bd9a7} /* (5, 12, 2) {real, imag} */,
  {32'hc0244059, 32'hc09bbbf3} /* (5, 12, 1) {real, imag} */,
  {32'h3f856516, 32'hbfd20114} /* (5, 12, 0) {real, imag} */,
  {32'hc053eee8, 32'h4037221c} /* (5, 11, 31) {real, imag} */,
  {32'hc03fa768, 32'h40848559} /* (5, 11, 30) {real, imag} */,
  {32'hc05bfddc, 32'h40d5f9bd} /* (5, 11, 29) {real, imag} */,
  {32'hc10a90dc, 32'h406f5a1f} /* (5, 11, 28) {real, imag} */,
  {32'hc0a3f493, 32'h4039041a} /* (5, 11, 27) {real, imag} */,
  {32'h3fbb4147, 32'h404ab3bb} /* (5, 11, 26) {real, imag} */,
  {32'hc05613bc, 32'h40ec7824} /* (5, 11, 25) {real, imag} */,
  {32'hc1203c30, 32'h4148f9ab} /* (5, 11, 24) {real, imag} */,
  {32'hc12087c7, 32'h40e23a33} /* (5, 11, 23) {real, imag} */,
  {32'h3fa26cfc, 32'hc00acc76} /* (5, 11, 22) {real, imag} */,
  {32'hc067d619, 32'hc052d2d3} /* (5, 11, 21) {real, imag} */,
  {32'h409d008a, 32'hc0244a3f} /* (5, 11, 20) {real, imag} */,
  {32'h402905fc, 32'h403cbcf4} /* (5, 11, 19) {real, imag} */,
  {32'h3b2b6800, 32'h40e66294} /* (5, 11, 18) {real, imag} */,
  {32'hbffe336c, 32'h4118ace0} /* (5, 11, 17) {real, imag} */,
  {32'hc0c26858, 32'h40ddd028} /* (5, 11, 16) {real, imag} */,
  {32'hc07a647f, 32'h40282cd4} /* (5, 11, 15) {real, imag} */,
  {32'hc00ccbb6, 32'hbef84b80} /* (5, 11, 14) {real, imag} */,
  {32'hc0c9bf74, 32'h40732456} /* (5, 11, 13) {real, imag} */,
  {32'hc00a5fa1, 32'h410024cc} /* (5, 11, 12) {real, imag} */,
  {32'h40b630d6, 32'hc0bb3399} /* (5, 11, 11) {real, imag} */,
  {32'hc108a5e0, 32'hc08b7d37} /* (5, 11, 10) {real, imag} */,
  {32'hc11aca98, 32'h3ff7dbd4} /* (5, 11, 9) {real, imag} */,
  {32'h3fe153b4, 32'h400873c2} /* (5, 11, 8) {real, imag} */,
  {32'h40636622, 32'hc0a9c095} /* (5, 11, 7) {real, imag} */,
  {32'h405f0e1e, 32'hbf27bf68} /* (5, 11, 6) {real, imag} */,
  {32'h40f7bfdd, 32'hc0311fa4} /* (5, 11, 5) {real, imag} */,
  {32'hc0201f0a, 32'hc13ebe96} /* (5, 11, 4) {real, imag} */,
  {32'hc039f5c9, 32'hbfcbf558} /* (5, 11, 3) {real, imag} */,
  {32'h4030482b, 32'h40a08bc4} /* (5, 11, 2) {real, imag} */,
  {32'hbf9dded0, 32'h4036a19b} /* (5, 11, 1) {real, imag} */,
  {32'h3e891180, 32'hc001bf48} /* (5, 11, 0) {real, imag} */,
  {32'h409616a9, 32'h40163c4d} /* (5, 10, 31) {real, imag} */,
  {32'h4105670b, 32'h4004af28} /* (5, 10, 30) {real, imag} */,
  {32'h407c47b4, 32'hc02646dd} /* (5, 10, 29) {real, imag} */,
  {32'h3ffc2362, 32'hc0cfa45c} /* (5, 10, 28) {real, imag} */,
  {32'h409288ac, 32'h3fa03dc0} /* (5, 10, 27) {real, imag} */,
  {32'h40208cb0, 32'hc03c2657} /* (5, 10, 26) {real, imag} */,
  {32'hbf7dcbd4, 32'h403b2ce4} /* (5, 10, 25) {real, imag} */,
  {32'h40486f3f, 32'h3f9a3458} /* (5, 10, 24) {real, imag} */,
  {32'h412da256, 32'hc11c8458} /* (5, 10, 23) {real, imag} */,
  {32'hc0f46ddc, 32'hc0a76dc8} /* (5, 10, 22) {real, imag} */,
  {32'hc10b6b83, 32'h405bf782} /* (5, 10, 21) {real, imag} */,
  {32'h3f4d7684, 32'hbff5b7c6} /* (5, 10, 20) {real, imag} */,
  {32'h40bfd3fe, 32'h405669fe} /* (5, 10, 19) {real, imag} */,
  {32'h413c750b, 32'h40540edd} /* (5, 10, 18) {real, imag} */,
  {32'h40e8f38c, 32'h41210bb3} /* (5, 10, 17) {real, imag} */,
  {32'h40ffbb34, 32'hbfea1ca4} /* (5, 10, 16) {real, imag} */,
  {32'h40d31554, 32'h405b3b39} /* (5, 10, 15) {real, imag} */,
  {32'hbf866ec3, 32'h410c760f} /* (5, 10, 14) {real, imag} */,
  {32'hc02ef146, 32'h4120308e} /* (5, 10, 13) {real, imag} */,
  {32'h412dcb8e, 32'h3f73da28} /* (5, 10, 12) {real, imag} */,
  {32'h40c59496, 32'hc04eff2a} /* (5, 10, 11) {real, imag} */,
  {32'h402341a0, 32'hbf384538} /* (5, 10, 10) {real, imag} */,
  {32'h40ee1b1d, 32'h4163645f} /* (5, 10, 9) {real, imag} */,
  {32'h416ea35d, 32'h414fe958} /* (5, 10, 8) {real, imag} */,
  {32'h40b962ef, 32'h417c00c3} /* (5, 10, 7) {real, imag} */,
  {32'h3f4d9148, 32'h412edc2d} /* (5, 10, 6) {real, imag} */,
  {32'h3e1d0670, 32'h41446659} /* (5, 10, 5) {real, imag} */,
  {32'h409b87d9, 32'h40c53821} /* (5, 10, 4) {real, imag} */,
  {32'hbf1815dc, 32'h3f1e5a0a} /* (5, 10, 3) {real, imag} */,
  {32'h40333a68, 32'h404a1252} /* (5, 10, 2) {real, imag} */,
  {32'h411b5de2, 32'hbf6f2154} /* (5, 10, 1) {real, imag} */,
  {32'h40c6aa16, 32'hbf799e04} /* (5, 10, 0) {real, imag} */,
  {32'hc05539b2, 32'hc0e9bd96} /* (5, 9, 31) {real, imag} */,
  {32'h3fb04270, 32'hc1418238} /* (5, 9, 30) {real, imag} */,
  {32'hc0c132ee, 32'h3fe66bb4} /* (5, 9, 29) {real, imag} */,
  {32'hc163158e, 32'h4156501c} /* (5, 9, 28) {real, imag} */,
  {32'hc0ef58d0, 32'h4137e2d7} /* (5, 9, 27) {real, imag} */,
  {32'h404d732e, 32'h413106ee} /* (5, 9, 26) {real, imag} */,
  {32'h3eb12108, 32'h41045832} /* (5, 9, 25) {real, imag} */,
  {32'h40a80240, 32'h40c190a1} /* (5, 9, 24) {real, imag} */,
  {32'h40dab4fc, 32'h3f9ea998} /* (5, 9, 23) {real, imag} */,
  {32'h405ffc82, 32'h411dee50} /* (5, 9, 22) {real, imag} */,
  {32'hc09c73a5, 32'h40396516} /* (5, 9, 21) {real, imag} */,
  {32'h40212519, 32'h40980316} /* (5, 9, 20) {real, imag} */,
  {32'hc1383334, 32'h412ee8f8} /* (5, 9, 19) {real, imag} */,
  {32'hc07dff94, 32'hbfcfc2e8} /* (5, 9, 18) {real, imag} */,
  {32'hc16b9816, 32'hc0ede3ed} /* (5, 9, 17) {real, imag} */,
  {32'hc113cac5, 32'hc107ff82} /* (5, 9, 16) {real, imag} */,
  {32'hc09a263a, 32'hc0e04fca} /* (5, 9, 15) {real, imag} */,
  {32'h4031d56e, 32'hc0ae042f} /* (5, 9, 14) {real, imag} */,
  {32'hc039dca6, 32'hc152d1d4} /* (5, 9, 13) {real, imag} */,
  {32'hc1422fd4, 32'hc0b3c99d} /* (5, 9, 12) {real, imag} */,
  {32'hc18c9253, 32'hc120966d} /* (5, 9, 11) {real, imag} */,
  {32'hc0da9574, 32'hc12e0386} /* (5, 9, 10) {real, imag} */,
  {32'h40ec48dc, 32'hc0fcbc1a} /* (5, 9, 9) {real, imag} */,
  {32'h3f8d9d30, 32'hc094d290} /* (5, 9, 8) {real, imag} */,
  {32'hc080f432, 32'hc0ddddf6} /* (5, 9, 7) {real, imag} */,
  {32'hc0ac34d2, 32'h40d8aede} /* (5, 9, 6) {real, imag} */,
  {32'hc00a73e4, 32'h407b5445} /* (5, 9, 5) {real, imag} */,
  {32'h40e46545, 32'hc07a6aab} /* (5, 9, 4) {real, imag} */,
  {32'h4154fcb4, 32'h40f7d697} /* (5, 9, 3) {real, imag} */,
  {32'hbfb2839c, 32'h4120f7d4} /* (5, 9, 2) {real, imag} */,
  {32'h400bfb38, 32'h41291a6e} /* (5, 9, 1) {real, imag} */,
  {32'hbf123a32, 32'h408846f2} /* (5, 9, 0) {real, imag} */,
  {32'hc09f3baa, 32'h41301560} /* (5, 8, 31) {real, imag} */,
  {32'hc10e49dc, 32'h41906fa5} /* (5, 8, 30) {real, imag} */,
  {32'hc17b680d, 32'h4028678a} /* (5, 8, 29) {real, imag} */,
  {32'h3f23e5a8, 32'h400284c3} /* (5, 8, 28) {real, imag} */,
  {32'hc03d381e, 32'h40341f0a} /* (5, 8, 27) {real, imag} */,
  {32'hc179a22b, 32'h416bf485} /* (5, 8, 26) {real, imag} */,
  {32'hc17e5722, 32'h40a4952c} /* (5, 8, 25) {real, imag} */,
  {32'hbf292ff8, 32'hbd4d2a80} /* (5, 8, 24) {real, imag} */,
  {32'hc054001b, 32'h3f9bf9aa} /* (5, 8, 23) {real, imag} */,
  {32'hc1594144, 32'hc00037dc} /* (5, 8, 22) {real, imag} */,
  {32'hc056487a, 32'hc1516f95} /* (5, 8, 21) {real, imag} */,
  {32'h41297a00, 32'hc16cf2f3} /* (5, 8, 20) {real, imag} */,
  {32'h409d070c, 32'h3ec9adc0} /* (5, 8, 19) {real, imag} */,
  {32'h4020ed24, 32'hc0ab68e4} /* (5, 8, 18) {real, imag} */,
  {32'hc11eb83a, 32'hc0f8c327} /* (5, 8, 17) {real, imag} */,
  {32'hc1416f53, 32'h409b94df} /* (5, 8, 16) {real, imag} */,
  {32'hbf75e838, 32'hc0197252} /* (5, 8, 15) {real, imag} */,
  {32'h41404e80, 32'hc093bbaa} /* (5, 8, 14) {real, imag} */,
  {32'h4000b880, 32'h3fae1ce8} /* (5, 8, 13) {real, imag} */,
  {32'hbe30d850, 32'hc0689975} /* (5, 8, 12) {real, imag} */,
  {32'h40aa7fd2, 32'hc0ab365a} /* (5, 8, 11) {real, imag} */,
  {32'h3ea09740, 32'h401b888c} /* (5, 8, 10) {real, imag} */,
  {32'h40634724, 32'hc109ce8c} /* (5, 8, 9) {real, imag} */,
  {32'h40bb5057, 32'h4037089a} /* (5, 8, 8) {real, imag} */,
  {32'hc0adabe4, 32'h4145c776} /* (5, 8, 7) {real, imag} */,
  {32'hc10ec20a, 32'hbf5c91e0} /* (5, 8, 6) {real, imag} */,
  {32'h3f997014, 32'h3f3a7630} /* (5, 8, 5) {real, imag} */,
  {32'h410965f2, 32'h3ff544f0} /* (5, 8, 4) {real, imag} */,
  {32'h40d2667a, 32'h3e866950} /* (5, 8, 3) {real, imag} */,
  {32'hc13c5cdc, 32'hc00b703e} /* (5, 8, 2) {real, imag} */,
  {32'hc15ee81e, 32'hc0e27fba} /* (5, 8, 1) {real, imag} */,
  {32'hc0d1f165, 32'h402d0990} /* (5, 8, 0) {real, imag} */,
  {32'h411cf538, 32'h3f975774} /* (5, 7, 31) {real, imag} */,
  {32'h3f8ebe10, 32'hc07e8a28} /* (5, 7, 30) {real, imag} */,
  {32'h3fc395c2, 32'hc1c0f264} /* (5, 7, 29) {real, imag} */,
  {32'h40bd4a55, 32'hc1a5309e} /* (5, 7, 28) {real, imag} */,
  {32'h409fd205, 32'h4003c3cb} /* (5, 7, 27) {real, imag} */,
  {32'h41175d76, 32'h41006010} /* (5, 7, 26) {real, imag} */,
  {32'hc030cd71, 32'hc0d47da7} /* (5, 7, 25) {real, imag} */,
  {32'hc0e63562, 32'hc133213c} /* (5, 7, 24) {real, imag} */,
  {32'hc0422891, 32'h412c0a1c} /* (5, 7, 23) {real, imag} */,
  {32'h3fc9e780, 32'h40a892a3} /* (5, 7, 22) {real, imag} */,
  {32'hc0f2a942, 32'hc13a4d7a} /* (5, 7, 21) {real, imag} */,
  {32'h3f36cb70, 32'hc1eb1e32} /* (5, 7, 20) {real, imag} */,
  {32'h409fd626, 32'hc142accd} /* (5, 7, 19) {real, imag} */,
  {32'hc1dce7ce, 32'h414798e8} /* (5, 7, 18) {real, imag} */,
  {32'hc1bb5d2f, 32'h416bd4c0} /* (5, 7, 17) {real, imag} */,
  {32'hc170c69c, 32'h4187c337} /* (5, 7, 16) {real, imag} */,
  {32'h3f6ff074, 32'h417edf13} /* (5, 7, 15) {real, imag} */,
  {32'h3f9d1a64, 32'h407f2222} /* (5, 7, 14) {real, imag} */,
  {32'hc18b62f3, 32'h40bbdd5b} /* (5, 7, 13) {real, imag} */,
  {32'hc15fb25d, 32'h4121a6d0} /* (5, 7, 12) {real, imag} */,
  {32'h41342d4a, 32'h4179d6e7} /* (5, 7, 11) {real, imag} */,
  {32'hc01fc134, 32'h40c62c24} /* (5, 7, 10) {real, imag} */,
  {32'hc0c1a7c7, 32'hc09490b2} /* (5, 7, 9) {real, imag} */,
  {32'h40a92102, 32'h410a6232} /* (5, 7, 8) {real, imag} */,
  {32'h40db2cce, 32'h40de110e} /* (5, 7, 7) {real, imag} */,
  {32'hc04b6478, 32'hbec48638} /* (5, 7, 6) {real, imag} */,
  {32'h410dea4b, 32'hbf22accc} /* (5, 7, 5) {real, imag} */,
  {32'h3fcc047c, 32'h411f3277} /* (5, 7, 4) {real, imag} */,
  {32'hc0def91d, 32'h4118799e} /* (5, 7, 3) {real, imag} */,
  {32'hc1584d5e, 32'hc19a0c5f} /* (5, 7, 2) {real, imag} */,
  {32'hbff39ad0, 32'hc14617f2} /* (5, 7, 1) {real, imag} */,
  {32'h40f70198, 32'h40883a4e} /* (5, 7, 0) {real, imag} */,
  {32'hc0bd95da, 32'hbebbc438} /* (5, 6, 31) {real, imag} */,
  {32'hc1184339, 32'h40e0b386} /* (5, 6, 30) {real, imag} */,
  {32'h4081069c, 32'h408734ee} /* (5, 6, 29) {real, imag} */,
  {32'h3fc62e9a, 32'h40f78596} /* (5, 6, 28) {real, imag} */,
  {32'hbfa4b5f0, 32'hbfc03800} /* (5, 6, 27) {real, imag} */,
  {32'hc0ab6f4e, 32'h403191f0} /* (5, 6, 26) {real, imag} */,
  {32'hc1012930, 32'h40bb119e} /* (5, 6, 25) {real, imag} */,
  {32'hc0f64d26, 32'h41aeeda4} /* (5, 6, 24) {real, imag} */,
  {32'hc106ee9e, 32'h4112bc20} /* (5, 6, 23) {real, imag} */,
  {32'hc11cf703, 32'hc0629e1d} /* (5, 6, 22) {real, imag} */,
  {32'hc04da3f8, 32'hc102a206} /* (5, 6, 21) {real, imag} */,
  {32'hc04f040c, 32'hc10dbef2} /* (5, 6, 20) {real, imag} */,
  {32'hc013bcc0, 32'hc087dc66} /* (5, 6, 19) {real, imag} */,
  {32'hc02ec22e, 32'h40709eb6} /* (5, 6, 18) {real, imag} */,
  {32'h40681250, 32'h409f91e4} /* (5, 6, 17) {real, imag} */,
  {32'h419a6e21, 32'h40c35b33} /* (5, 6, 16) {real, imag} */,
  {32'h41130794, 32'hc1a8f290} /* (5, 6, 15) {real, imag} */,
  {32'h3f29264e, 32'hc0ab7acd} /* (5, 6, 14) {real, imag} */,
  {32'h41104666, 32'hc127af02} /* (5, 6, 13) {real, imag} */,
  {32'h41a6d914, 32'hc14452a7} /* (5, 6, 12) {real, imag} */,
  {32'h41935ffc, 32'hc15c9197} /* (5, 6, 11) {real, imag} */,
  {32'h4137c715, 32'hc106adcc} /* (5, 6, 10) {real, imag} */,
  {32'hc0f8f3f7, 32'hc185a552} /* (5, 6, 9) {real, imag} */,
  {32'hc048057c, 32'h40bc17c4} /* (5, 6, 8) {real, imag} */,
  {32'hbf58d128, 32'h4043fc9a} /* (5, 6, 7) {real, imag} */,
  {32'h4017acc2, 32'hc044432c} /* (5, 6, 6) {real, imag} */,
  {32'hc16e7789, 32'h40087070} /* (5, 6, 5) {real, imag} */,
  {32'h402a5768, 32'hbfe57594} /* (5, 6, 4) {real, imag} */,
  {32'h416585ce, 32'hc0e3bf95} /* (5, 6, 3) {real, imag} */,
  {32'hc0e2f46a, 32'h3edd9a90} /* (5, 6, 2) {real, imag} */,
  {32'hbf06aa44, 32'h40d076ba} /* (5, 6, 1) {real, imag} */,
  {32'h3f6d2b9b, 32'hc08fc658} /* (5, 6, 0) {real, imag} */,
  {32'hc1601fa8, 32'h41384704} /* (5, 5, 31) {real, imag} */,
  {32'hc20e72c2, 32'h4123789c} /* (5, 5, 30) {real, imag} */,
  {32'hc199d8ac, 32'h41869ee3} /* (5, 5, 29) {real, imag} */,
  {32'hc082c2ec, 32'h41e0a2b2} /* (5, 5, 28) {real, imag} */,
  {32'h4050688a, 32'h41d4ec19} /* (5, 5, 27) {real, imag} */,
  {32'h403cb20c, 32'h40a0143e} /* (5, 5, 26) {real, imag} */,
  {32'hc17ef3a3, 32'hc0321c58} /* (5, 5, 25) {real, imag} */,
  {32'hc136960d, 32'hc087d646} /* (5, 5, 24) {real, imag} */,
  {32'h40988ea2, 32'h3fdc8cce} /* (5, 5, 23) {real, imag} */,
  {32'h40ad5b75, 32'h411cacf0} /* (5, 5, 22) {real, imag} */,
  {32'hc10a4445, 32'h400c485a} /* (5, 5, 21) {real, imag} */,
  {32'h4026b896, 32'hc0942cf2} /* (5, 5, 20) {real, imag} */,
  {32'h40d57a88, 32'hbf482b90} /* (5, 5, 19) {real, imag} */,
  {32'h4005f84f, 32'h405a3fd4} /* (5, 5, 18) {real, imag} */,
  {32'h3e944630, 32'hc100aae7} /* (5, 5, 17) {real, imag} */,
  {32'hc0eb0f55, 32'hc11641e4} /* (5, 5, 16) {real, imag} */,
  {32'hc0ae9442, 32'hc044d3a4} /* (5, 5, 15) {real, imag} */,
  {32'hc108312e, 32'hc0fd0464} /* (5, 5, 14) {real, imag} */,
  {32'hbefd8940, 32'hc0c8e2e5} /* (5, 5, 13) {real, imag} */,
  {32'h404fb71b, 32'h3f0a0bc8} /* (5, 5, 12) {real, imag} */,
  {32'h40f80612, 32'h40debc8f} /* (5, 5, 11) {real, imag} */,
  {32'hc0c42070, 32'h418db976} /* (5, 5, 10) {real, imag} */,
  {32'hc0cf53ad, 32'h40906aa8} /* (5, 5, 9) {real, imag} */,
  {32'hc104604e, 32'hc15b01d6} /* (5, 5, 8) {real, imag} */,
  {32'hc19331df, 32'h409913c2} /* (5, 5, 7) {real, imag} */,
  {32'hc1a22de0, 32'hc0b09ee9} /* (5, 5, 6) {real, imag} */,
  {32'hc1826622, 32'hc11ceff2} /* (5, 5, 5) {real, imag} */,
  {32'hc0c2276c, 32'hc0daaa88} /* (5, 5, 4) {real, imag} */,
  {32'hc177dfa0, 32'h40d94ad8} /* (5, 5, 3) {real, imag} */,
  {32'hc1aadf8c, 32'h4132c67d} /* (5, 5, 2) {real, imag} */,
  {32'hc12162e8, 32'h3f8bf43a} /* (5, 5, 1) {real, imag} */,
  {32'hc09f27dc, 32'h413093ab} /* (5, 5, 0) {real, imag} */,
  {32'h40e7a966, 32'hc06ee519} /* (5, 4, 31) {real, imag} */,
  {32'h41cb2724, 32'h40f69caf} /* (5, 4, 30) {real, imag} */,
  {32'h41b17209, 32'hbfabb6f8} /* (5, 4, 29) {real, imag} */,
  {32'h40fc9328, 32'hc16593e4} /* (5, 4, 28) {real, imag} */,
  {32'h41248584, 32'hc10562e6} /* (5, 4, 27) {real, imag} */,
  {32'h41c07f3e, 32'hc18d81f4} /* (5, 4, 26) {real, imag} */,
  {32'h41dbf6aa, 32'hc0688b0e} /* (5, 4, 25) {real, imag} */,
  {32'h41eb6bdf, 32'h411b4bcb} /* (5, 4, 24) {real, imag} */,
  {32'h41825b12, 32'h4105ae94} /* (5, 4, 23) {real, imag} */,
  {32'h40db5f36, 32'hc08d5f6c} /* (5, 4, 22) {real, imag} */,
  {32'hc1425493, 32'hbec99600} /* (5, 4, 21) {real, imag} */,
  {32'h40251654, 32'h40224aa8} /* (5, 4, 20) {real, imag} */,
  {32'hbfd8c150, 32'hc01f30e0} /* (5, 4, 19) {real, imag} */,
  {32'hc13c9552, 32'h3e3f7f40} /* (5, 4, 18) {real, imag} */,
  {32'hc1e711e6, 32'hc1599c94} /* (5, 4, 17) {real, imag} */,
  {32'hc1bc208c, 32'hc180819a} /* (5, 4, 16) {real, imag} */,
  {32'h40e61aec, 32'hbf8833a0} /* (5, 4, 15) {real, imag} */,
  {32'h40c14dde, 32'h406f1ea2} /* (5, 4, 14) {real, imag} */,
  {32'h40f1f1bd, 32'h41312782} /* (5, 4, 13) {real, imag} */,
  {32'h3de6f440, 32'h3f7cfb48} /* (5, 4, 12) {real, imag} */,
  {32'h409b8aea, 32'hc06629eb} /* (5, 4, 11) {real, imag} */,
  {32'h41bdd453, 32'hc0e4725c} /* (5, 4, 10) {real, imag} */,
  {32'h41f57d38, 32'h412e7a38} /* (5, 4, 9) {real, imag} */,
  {32'h41d504de, 32'h40fbbd20} /* (5, 4, 8) {real, imag} */,
  {32'h4174ee60, 32'hc1023c06} /* (5, 4, 7) {real, imag} */,
  {32'h41bc596b, 32'h3f9821a0} /* (5, 4, 6) {real, imag} */,
  {32'h41e0ec82, 32'h41483193} /* (5, 4, 5) {real, imag} */,
  {32'h3ddb0de0, 32'h41373116} /* (5, 4, 4) {real, imag} */,
  {32'hc12b3142, 32'h40826fbc} /* (5, 4, 3) {real, imag} */,
  {32'hc14547b9, 32'hc19237ba} /* (5, 4, 2) {real, imag} */,
  {32'hbf1bc2e0, 32'hc1c333f5} /* (5, 4, 1) {real, imag} */,
  {32'hc0031804, 32'hc0f5d84e} /* (5, 4, 0) {real, imag} */,
  {32'hc0517df6, 32'hc07f957c} /* (5, 3, 31) {real, imag} */,
  {32'hc07d3612, 32'hc1366011} /* (5, 3, 30) {real, imag} */,
  {32'h411e6043, 32'hc1c8507e} /* (5, 3, 29) {real, imag} */,
  {32'hc1163907, 32'h401cffd2} /* (5, 3, 28) {real, imag} */,
  {32'hc0dba848, 32'hc18b22f6} /* (5, 3, 27) {real, imag} */,
  {32'h4082ff4e, 32'hc1919ca3} /* (5, 3, 26) {real, imag} */,
  {32'h41843e7f, 32'hc173198c} /* (5, 3, 25) {real, imag} */,
  {32'h40884593, 32'hc181af6c} /* (5, 3, 24) {real, imag} */,
  {32'hc122fb12, 32'hc13d120f} /* (5, 3, 23) {real, imag} */,
  {32'hbee40e60, 32'hc139b466} /* (5, 3, 22) {real, imag} */,
  {32'hbf910f7c, 32'hc08c69af} /* (5, 3, 21) {real, imag} */,
  {32'hc048df80, 32'hc17db154} /* (5, 3, 20) {real, imag} */,
  {32'hc153391a, 32'hc1a5b311} /* (5, 3, 19) {real, imag} */,
  {32'hc21201ff, 32'hc179ee39} /* (5, 3, 18) {real, imag} */,
  {32'hc22969f4, 32'h403cd020} /* (5, 3, 17) {real, imag} */,
  {32'hc1db7651, 32'hc0da0dca} /* (5, 3, 16) {real, imag} */,
  {32'hc02fd032, 32'h4088ae7c} /* (5, 3, 15) {real, imag} */,
  {32'h410280fd, 32'h41d8fce7} /* (5, 3, 14) {real, imag} */,
  {32'h3f71945a, 32'h418cc140} /* (5, 3, 13) {real, imag} */,
  {32'hc036bca8, 32'h41a9b703} /* (5, 3, 12) {real, imag} */,
  {32'hc11074f1, 32'h40ccf34a} /* (5, 3, 11) {real, imag} */,
  {32'hc05efe28, 32'h41a0ade8} /* (5, 3, 10) {real, imag} */,
  {32'h412f6bca, 32'h41caa346} /* (5, 3, 9) {real, imag} */,
  {32'h40945208, 32'h41cec353} /* (5, 3, 8) {real, imag} */,
  {32'h408bc64a, 32'h41ae207a} /* (5, 3, 7) {real, imag} */,
  {32'hbffaa410, 32'h41663800} /* (5, 3, 6) {real, imag} */,
  {32'hc057aea5, 32'h4106afef} /* (5, 3, 5) {real, imag} */,
  {32'hc11ea0a9, 32'h4140e63e} /* (5, 3, 4) {real, imag} */,
  {32'hc05d0007, 32'h3f13f9b8} /* (5, 3, 3) {real, imag} */,
  {32'hc106a4c7, 32'h414615be} /* (5, 3, 2) {real, imag} */,
  {32'h40b03dc6, 32'h41c6f748} /* (5, 3, 1) {real, imag} */,
  {32'h414bd792, 32'h414436f2} /* (5, 3, 0) {real, imag} */,
  {32'h3e5fbbe0, 32'h4169816a} /* (5, 2, 31) {real, imag} */,
  {32'hc0681f9b, 32'h419f4347} /* (5, 2, 30) {real, imag} */,
  {32'hc1629d6e, 32'h41105486} /* (5, 2, 29) {real, imag} */,
  {32'hc1c623ff, 32'h418000cc} /* (5, 2, 28) {real, imag} */,
  {32'hc1b167b6, 32'h41224fb2} /* (5, 2, 27) {real, imag} */,
  {32'h3ea47bb8, 32'hc0a740b0} /* (5, 2, 26) {real, imag} */,
  {32'h40a07906, 32'h41041f62} /* (5, 2, 25) {real, imag} */,
  {32'hc148a5af, 32'h4211a140} /* (5, 2, 24) {real, imag} */,
  {32'hc207f285, 32'h42350611} /* (5, 2, 23) {real, imag} */,
  {32'hc23ea14d, 32'h41d94b00} /* (5, 2, 22) {real, imag} */,
  {32'hc10a49a4, 32'h41025db2} /* (5, 2, 21) {real, imag} */,
  {32'h40806b06, 32'hc181993b} /* (5, 2, 20) {real, imag} */,
  {32'h40951395, 32'hc25175bc} /* (5, 2, 19) {real, imag} */,
  {32'h416aa445, 32'hc28c5288} /* (5, 2, 18) {real, imag} */,
  {32'h41a07f2a, 32'hc2711754} /* (5, 2, 17) {real, imag} */,
  {32'h3feefde0, 32'hc2570ffa} /* (5, 2, 16) {real, imag} */,
  {32'h412ee58c, 32'hc222dc76} /* (5, 2, 15) {real, imag} */,
  {32'h40c06836, 32'hc1a59bcc} /* (5, 2, 14) {real, imag} */,
  {32'h41f1a4c6, 32'hc1df5c00} /* (5, 2, 13) {real, imag} */,
  {32'h41c825aa, 32'hc1a8edcf} /* (5, 2, 12) {real, imag} */,
  {32'h40ea4f18, 32'hc18fb29e} /* (5, 2, 11) {real, imag} */,
  {32'h40b1b388, 32'h41e29658} /* (5, 2, 10) {real, imag} */,
  {32'h413b2758, 32'h4226f990} /* (5, 2, 9) {real, imag} */,
  {32'h40a1a728, 32'h422e97c1} /* (5, 2, 8) {real, imag} */,
  {32'hbf9316c4, 32'h41d462b0} /* (5, 2, 7) {real, imag} */,
  {32'h408b9fc8, 32'h41d80412} /* (5, 2, 6) {real, imag} */,
  {32'h4126bfb9, 32'h41db7409} /* (5, 2, 5) {real, imag} */,
  {32'h403ee341, 32'h4194b664} /* (5, 2, 4) {real, imag} */,
  {32'hc16690ef, 32'hc0718fd6} /* (5, 2, 3) {real, imag} */,
  {32'hc1760d2d, 32'h3ff98f04} /* (5, 2, 2) {real, imag} */,
  {32'hc1211b67, 32'h40cd3e08} /* (5, 2, 1) {real, imag} */,
  {32'hbfa33eae, 32'h40692764} /* (5, 2, 0) {real, imag} */,
  {32'h40df930c, 32'hc163d3a3} /* (5, 1, 31) {real, imag} */,
  {32'h4189082e, 32'hc1d9042d} /* (5, 1, 30) {real, imag} */,
  {32'h41c3fbb6, 32'hc1324fda} /* (5, 1, 29) {real, imag} */,
  {32'h41a8b04e, 32'hc12e3c4c} /* (5, 1, 28) {real, imag} */,
  {32'h41fddc4d, 32'hc17e9180} /* (5, 1, 27) {real, imag} */,
  {32'h422cea0e, 32'hc2011e85} /* (5, 1, 26) {real, imag} */,
  {32'h421e8581, 32'hc21aaa85} /* (5, 1, 25) {real, imag} */,
  {32'h41c4dc52, 32'hc1ee8887} /* (5, 1, 24) {real, imag} */,
  {32'h41ff9afb, 32'hc1f9b339} /* (5, 1, 23) {real, imag} */,
  {32'h41ac6653, 32'hc1d0f086} /* (5, 1, 22) {real, imag} */,
  {32'h4070a612, 32'hc206c052} /* (5, 1, 21) {real, imag} */,
  {32'hc1c84adc, 32'hbf672bd8} /* (5, 1, 20) {real, imag} */,
  {32'hc2225c66, 32'hc0362592} /* (5, 1, 19) {real, imag} */,
  {32'hc1df855e, 32'hc0a3fc4e} /* (5, 1, 18) {real, imag} */,
  {32'hc1d240aa, 32'h40c76aae} /* (5, 1, 17) {real, imag} */,
  {32'hc1270b4a, 32'h4121a4ed} /* (5, 1, 16) {real, imag} */,
  {32'hc1d9f06f, 32'h415fec83} /* (5, 1, 15) {real, imag} */,
  {32'hc1d67161, 32'h41e7ba20} /* (5, 1, 14) {real, imag} */,
  {32'hc14c5e15, 32'h4229442c} /* (5, 1, 13) {real, imag} */,
  {32'hc18db9ea, 32'h418b1916} /* (5, 1, 12) {real, imag} */,
  {32'hc152f882, 32'h419cfccc} /* (5, 1, 11) {real, imag} */,
  {32'h41a280f6, 32'h3eea2c80} /* (5, 1, 10) {real, imag} */,
  {32'h420eb02b, 32'h3ec80340} /* (5, 1, 9) {real, imag} */,
  {32'h411c8f6f, 32'hc09920e2} /* (5, 1, 8) {real, imag} */,
  {32'h4192bc75, 32'hc168f1c9} /* (5, 1, 7) {real, imag} */,
  {32'h3f8cf750, 32'hc0c1bf28} /* (5, 1, 6) {real, imag} */,
  {32'h40b2e68e, 32'hc1cb2c58} /* (5, 1, 5) {real, imag} */,
  {32'h412f4de0, 32'hc21bf7a5} /* (5, 1, 4) {real, imag} */,
  {32'h41a0bc7f, 32'hc202645f} /* (5, 1, 3) {real, imag} */,
  {32'h41cf6378, 32'hc1c30360} /* (5, 1, 2) {real, imag} */,
  {32'h41a2365c, 32'hc1d45f29} /* (5, 1, 1) {real, imag} */,
  {32'h40b9758a, 32'hc188aac8} /* (5, 1, 0) {real, imag} */,
  {32'h41611409, 32'hc148be62} /* (5, 0, 31) {real, imag} */,
  {32'h41f8ecc2, 32'hc1aa2c05} /* (5, 0, 30) {real, imag} */,
  {32'hc0b20224, 32'hc21fdc14} /* (5, 0, 29) {real, imag} */,
  {32'h41433a24, 32'hc206cffa} /* (5, 0, 28) {real, imag} */,
  {32'h423bb37e, 32'hc1c3ac3d} /* (5, 0, 27) {real, imag} */,
  {32'h41f8e70e, 32'hc1a2ac53} /* (5, 0, 26) {real, imag} */,
  {32'h4126a142, 32'hc1972bec} /* (5, 0, 25) {real, imag} */,
  {32'h412d1ae8, 32'hc20d4118} /* (5, 0, 24) {real, imag} */,
  {32'h40ce80ae, 32'hc15348a7} /* (5, 0, 23) {real, imag} */,
  {32'h40ebce48, 32'hc1c6ffa4} /* (5, 0, 22) {real, imag} */,
  {32'h40cdcb69, 32'hc2146619} /* (5, 0, 21) {real, imag} */,
  {32'h41579cba, 32'hc18733a3} /* (5, 0, 20) {real, imag} */,
  {32'hbdf79c20, 32'hc15150ca} /* (5, 0, 19) {real, imag} */,
  {32'h408f5bd0, 32'h3eeb50b0} /* (5, 0, 18) {real, imag} */,
  {32'hc1b8a78f, 32'hbc8ecc00} /* (5, 0, 17) {real, imag} */,
  {32'hc13ca061, 32'hbf2adec8} /* (5, 0, 16) {real, imag} */,
  {32'hc10ddb7e, 32'h41cf7988} /* (5, 0, 15) {real, imag} */,
  {32'hc1e8499a, 32'h41cc610e} /* (5, 0, 14) {real, imag} */,
  {32'hc20247fb, 32'h41d24e7c} /* (5, 0, 13) {real, imag} */,
  {32'hc1aa7bac, 32'h41ed0182} /* (5, 0, 12) {real, imag} */,
  {32'hc19d35bc, 32'h41b6777c} /* (5, 0, 11) {real, imag} */,
  {32'hc16c6528, 32'hc0b89200} /* (5, 0, 10) {real, imag} */,
  {32'hc0f64cd4, 32'hbfa2d1c6} /* (5, 0, 9) {real, imag} */,
  {32'h415ac5e8, 32'hc112afe1} /* (5, 0, 8) {real, imag} */,
  {32'h40a9de79, 32'hc005c133} /* (5, 0, 7) {real, imag} */,
  {32'hc0973804, 32'hc0edb170} /* (5, 0, 6) {real, imag} */,
  {32'hc0dc60dc, 32'hc20d61af} /* (5, 0, 5) {real, imag} */,
  {32'hc112d9f6, 32'hc207ed83} /* (5, 0, 4) {real, imag} */,
  {32'h40874cdd, 32'hc2043b9a} /* (5, 0, 3) {real, imag} */,
  {32'h41a5f5d8, 32'hc14be5d4} /* (5, 0, 2) {real, imag} */,
  {32'h3fcf4be8, 32'hc0eaa5b0} /* (5, 0, 1) {real, imag} */,
  {32'hbe962a8c, 32'hc15dc0dc} /* (5, 0, 0) {real, imag} */,
  {32'hc19c2492, 32'h4232caaf} /* (4, 31, 31) {real, imag} */,
  {32'hc1f1b4bc, 32'h42a05302} /* (4, 31, 30) {real, imag} */,
  {32'hc1c800d2, 32'h42c2c44f} /* (4, 31, 29) {real, imag} */,
  {32'hc17a193d, 32'h4299d1cc} /* (4, 31, 28) {real, imag} */,
  {32'hc167082e, 32'h428e606f} /* (4, 31, 27) {real, imag} */,
  {32'hc0e7b85c, 32'h429b7ff4} /* (4, 31, 26) {real, imag} */,
  {32'hc1040c85, 32'h4299e9bf} /* (4, 31, 25) {real, imag} */,
  {32'hc1c964ee, 32'h42a4994e} /* (4, 31, 24) {real, imag} */,
  {32'hc1e7a2c2, 32'h42842eac} /* (4, 31, 23) {real, imag} */,
  {32'hc1df2394, 32'h428e9288} /* (4, 31, 22) {real, imag} */,
  {32'hc19e1bbc, 32'h42309d3e} /* (4, 31, 21) {real, imag} */,
  {32'hc197aa90, 32'hc2489ada} /* (4, 31, 20) {real, imag} */,
  {32'hc08d26bc, 32'hc2816045} /* (4, 31, 19) {real, imag} */,
  {32'hc12f98f1, 32'hc27b9e90} /* (4, 31, 18) {real, imag} */,
  {32'hc1e77553, 32'hc298de25} /* (4, 31, 17) {real, imag} */,
  {32'hc21e9497, 32'hc2956209} /* (4, 31, 16) {real, imag} */,
  {32'h40e46c33, 32'hc29a63ca} /* (4, 31, 15) {real, imag} */,
  {32'h415a08e2, 32'hc2a18420} /* (4, 31, 14) {real, imag} */,
  {32'hc0810af8, 32'hc2875c8a} /* (4, 31, 13) {real, imag} */,
  {32'h41cde3f7, 32'hc2a61997} /* (4, 31, 12) {real, imag} */,
  {32'h41f010d8, 32'hc29a9cab} /* (4, 31, 11) {real, imag} */,
  {32'h41ad29e2, 32'h40f9ffdc} /* (4, 31, 10) {real, imag} */,
  {32'h41a62b5a, 32'h4267f40e} /* (4, 31, 9) {real, imag} */,
  {32'h4206efcd, 32'h428262ba} /* (4, 31, 8) {real, imag} */,
  {32'h4138ce8a, 32'h42717593} /* (4, 31, 7) {real, imag} */,
  {32'h402049a8, 32'h42883f3c} /* (4, 31, 6) {real, imag} */,
  {32'hc0447d90, 32'h426eade7} /* (4, 31, 5) {real, imag} */,
  {32'hc22fe324, 32'h42975b50} /* (4, 31, 4) {real, imag} */,
  {32'hc2149f7d, 32'h42c88606} /* (4, 31, 3) {real, imag} */,
  {32'hc21e9faa, 32'h428c9cb8} /* (4, 31, 2) {real, imag} */,
  {32'hc12b4b11, 32'h4282919b} /* (4, 31, 1) {real, imag} */,
  {32'hc1805f94, 32'h42311bdc} /* (4, 31, 0) {real, imag} */,
  {32'hbe317dc0, 32'hc235f564} /* (4, 30, 31) {real, imag} */,
  {32'hc05ea4a0, 32'hc257d019} /* (4, 30, 30) {real, imag} */,
  {32'hbef35b00, 32'hc20f50c0} /* (4, 30, 29) {real, imag} */,
  {32'hc0bf7bbc, 32'hc25b4092} /* (4, 30, 28) {real, imag} */,
  {32'h40a2cfea, 32'hc243f0ca} /* (4, 30, 27) {real, imag} */,
  {32'h41da39ab, 32'hc24825fa} /* (4, 30, 26) {real, imag} */,
  {32'h41b6ab70, 32'hc257b33c} /* (4, 30, 25) {real, imag} */,
  {32'hbf090330, 32'hc283105e} /* (4, 30, 24) {real, imag} */,
  {32'h3fdac010, 32'hc2505686} /* (4, 30, 23) {real, imag} */,
  {32'h410772f6, 32'hc25d6064} /* (4, 30, 22) {real, imag} */,
  {32'hc1139d4a, 32'hc1550012} /* (4, 30, 21) {real, imag} */,
  {32'hc25d9d18, 32'h425a48e1} /* (4, 30, 20) {real, imag} */,
  {32'hc24cf599, 32'h42541169} /* (4, 30, 19) {real, imag} */,
  {32'hc27d0df3, 32'h41ed1c22} /* (4, 30, 18) {real, imag} */,
  {32'hc21b2926, 32'h423bdaa8} /* (4, 30, 17) {real, imag} */,
  {32'hc16d06fd, 32'h427092b3} /* (4, 30, 16) {real, imag} */,
  {32'h41b5e540, 32'h42732d4c} /* (4, 30, 15) {real, imag} */,
  {32'h404519de, 32'h4275efb5} /* (4, 30, 14) {real, imag} */,
  {32'hc0c03716, 32'h426dc640} /* (4, 30, 13) {real, imag} */,
  {32'hc019aec8, 32'h424d21c2} /* (4, 30, 12) {real, imag} */,
  {32'h4094c155, 32'h41dd6104} /* (4, 30, 11) {real, imag} */,
  {32'h4216e8e2, 32'hc21dc35c} /* (4, 30, 10) {real, imag} */,
  {32'h421c08fa, 32'hc2634a12} /* (4, 30, 9) {real, imag} */,
  {32'h42475486, 32'hc27a66f2} /* (4, 30, 8) {real, imag} */,
  {32'h425c476b, 32'hc2913eda} /* (4, 30, 7) {real, imag} */,
  {32'h41b64dc4, 32'hc26f7957} /* (4, 30, 6) {real, imag} */,
  {32'hc028691c, 32'hc26dfbad} /* (4, 30, 5) {real, imag} */,
  {32'hc133f7dd, 32'hc24e83d8} /* (4, 30, 4) {real, imag} */,
  {32'h40433cb0, 32'hc2170cb4} /* (4, 30, 3) {real, imag} */,
  {32'h40c50eae, 32'hc2651907} /* (4, 30, 2) {real, imag} */,
  {32'h41b5891d, 32'hc26aaed7} /* (4, 30, 1) {real, imag} */,
  {32'h418dd878, 32'hc2264952} /* (4, 30, 0) {real, imag} */,
  {32'hbfe03c9c, 32'h40df2b98} /* (4, 29, 31) {real, imag} */,
  {32'h41d086ef, 32'h3d188f40} /* (4, 29, 30) {real, imag} */,
  {32'h41a63789, 32'hc13b367d} /* (4, 29, 29) {real, imag} */,
  {32'hbf80d920, 32'h40ba4516} /* (4, 29, 28) {real, imag} */,
  {32'hc1235f3d, 32'h41725920} /* (4, 29, 27) {real, imag} */,
  {32'h40918d62, 32'hbf916c04} /* (4, 29, 26) {real, imag} */,
  {32'h41503631, 32'hc114a9f2} /* (4, 29, 25) {real, imag} */,
  {32'hbef35280, 32'h40e1b5b1} /* (4, 29, 24) {real, imag} */,
  {32'hc115ae64, 32'h40daeff2} /* (4, 29, 23) {real, imag} */,
  {32'hc11c185c, 32'hc17548d1} /* (4, 29, 22) {real, imag} */,
  {32'h41069c07, 32'hc1b3acbe} /* (4, 29, 21) {real, imag} */,
  {32'hc195997a, 32'h40559bd0} /* (4, 29, 20) {real, imag} */,
  {32'hc23e6406, 32'hc0f324f8} /* (4, 29, 19) {real, imag} */,
  {32'hc2644828, 32'hc196eab8} /* (4, 29, 18) {real, imag} */,
  {32'hc2348195, 32'hc207f0b3} /* (4, 29, 17) {real, imag} */,
  {32'hc244da40, 32'hc20cf1db} /* (4, 29, 16) {real, imag} */,
  {32'hc1a18412, 32'hc168a521} /* (4, 29, 15) {real, imag} */,
  {32'hbfcd96b8, 32'hbf52d9b8} /* (4, 29, 14) {real, imag} */,
  {32'h41b984e2, 32'h40abe1f4} /* (4, 29, 13) {real, imag} */,
  {32'h4204db8c, 32'h4016300c} /* (4, 29, 12) {real, imag} */,
  {32'h419c3a82, 32'h41361fd2} /* (4, 29, 11) {real, imag} */,
  {32'h41c5c900, 32'h41a7fb4e} /* (4, 29, 10) {real, imag} */,
  {32'h42229cde, 32'h41a3a9f1} /* (4, 29, 9) {real, imag} */,
  {32'h4210ccdc, 32'h419b31f8} /* (4, 29, 8) {real, imag} */,
  {32'h4214f64d, 32'h41682778} /* (4, 29, 7) {real, imag} */,
  {32'h422ae55b, 32'hc0761988} /* (4, 29, 6) {real, imag} */,
  {32'h41dd40bb, 32'h3f3ee620} /* (4, 29, 5) {real, imag} */,
  {32'h4117679d, 32'hbfcbdb18} /* (4, 29, 4) {real, imag} */,
  {32'h420f6e76, 32'h41a645ee} /* (4, 29, 3) {real, imag} */,
  {32'h42474084, 32'h41b98073} /* (4, 29, 2) {real, imag} */,
  {32'h414ee089, 32'h4170b8ae} /* (4, 29, 1) {real, imag} */,
  {32'hc0d546b0, 32'h40984e1e} /* (4, 29, 0) {real, imag} */,
  {32'hc0753844, 32'h41499e1d} /* (4, 28, 31) {real, imag} */,
  {32'h41141ae6, 32'h40625b50} /* (4, 28, 30) {real, imag} */,
  {32'h41cc533f, 32'hbfba98a0} /* (4, 28, 29) {real, imag} */,
  {32'h419838bc, 32'h41cf3793} /* (4, 28, 28) {real, imag} */,
  {32'h41120195, 32'h410e01ef} /* (4, 28, 27) {real, imag} */,
  {32'hc0c96614, 32'h41a44762} /* (4, 28, 26) {real, imag} */,
  {32'hc0e5d968, 32'h4206fad4} /* (4, 28, 25) {real, imag} */,
  {32'h3fdde3f0, 32'h41b6aac0} /* (4, 28, 24) {real, imag} */,
  {32'h41527026, 32'h4205b2a2} /* (4, 28, 23) {real, imag} */,
  {32'h409d901c, 32'h41f67d4e} /* (4, 28, 22) {real, imag} */,
  {32'h409d38de, 32'h41d76ba5} /* (4, 28, 21) {real, imag} */,
  {32'hc12e5216, 32'hc1b23ae0} /* (4, 28, 20) {real, imag} */,
  {32'hc1576f74, 32'hc1b7ad12} /* (4, 28, 19) {real, imag} */,
  {32'hc1da35b2, 32'hc1cba5b6} /* (4, 28, 18) {real, imag} */,
  {32'hc201b3e8, 32'hc1854982} /* (4, 28, 17) {real, imag} */,
  {32'h409d5a7e, 32'hc10bcb11} /* (4, 28, 16) {real, imag} */,
  {32'h402db654, 32'hc19c5093} /* (4, 28, 15) {real, imag} */,
  {32'hc0c6246a, 32'hc1d48ea4} /* (4, 28, 14) {real, imag} */,
  {32'hc0a29292, 32'hc1d26c43} /* (4, 28, 13) {real, imag} */,
  {32'hc0d7884f, 32'hc1989431} /* (4, 28, 12) {real, imag} */,
  {32'h4082f996, 32'hc1376ab1} /* (4, 28, 11) {real, imag} */,
  {32'h418b1a9a, 32'h411931f3} /* (4, 28, 10) {real, imag} */,
  {32'h421a8a00, 32'h4204a2ee} /* (4, 28, 9) {real, imag} */,
  {32'h41eb9cf4, 32'h4218d838} /* (4, 28, 8) {real, imag} */,
  {32'h41e3094a, 32'h41b6d3d8} /* (4, 28, 7) {real, imag} */,
  {32'h41d8b212, 32'h41992be9} /* (4, 28, 6) {real, imag} */,
  {32'hbffbe490, 32'h41c95dca} /* (4, 28, 5) {real, imag} */,
  {32'h410fba5f, 32'h4140d4d9} /* (4, 28, 4) {real, imag} */,
  {32'hc0ea11b3, 32'h41f6e046} /* (4, 28, 3) {real, imag} */,
  {32'hc1436cb2, 32'h4245ce7a} /* (4, 28, 2) {real, imag} */,
  {32'hc127a924, 32'h42005302} /* (4, 28, 1) {real, imag} */,
  {32'h3fae8078, 32'h4196a48f} /* (4, 28, 0) {real, imag} */,
  {32'h413a5aad, 32'hc1aa379e} /* (4, 27, 31) {real, imag} */,
  {32'h3f235eb0, 32'hc19a1ca0} /* (4, 27, 30) {real, imag} */,
  {32'h414fde62, 32'hc1d28a42} /* (4, 27, 29) {real, imag} */,
  {32'h4109d881, 32'hc22206ef} /* (4, 27, 28) {real, imag} */,
  {32'hc0a01ebe, 32'hc232fa47} /* (4, 27, 27) {real, imag} */,
  {32'hc09cce3a, 32'hc216bb4d} /* (4, 27, 26) {real, imag} */,
  {32'h3fbeda48, 32'hc1d22a5e} /* (4, 27, 25) {real, imag} */,
  {32'h409ec3a6, 32'hc23196b9} /* (4, 27, 24) {real, imag} */,
  {32'h4075abff, 32'hc201d1aa} /* (4, 27, 23) {real, imag} */,
  {32'hbf320dc8, 32'hc201d9a6} /* (4, 27, 22) {real, imag} */,
  {32'hc0a2ef62, 32'hc1a5bdab} /* (4, 27, 21) {real, imag} */,
  {32'hbfa9f502, 32'hc104f40a} /* (4, 27, 20) {real, imag} */,
  {32'hc1a39f87, 32'hbf3e3938} /* (4, 27, 19) {real, imag} */,
  {32'hc1bdbb6b, 32'h417c6b64} /* (4, 27, 18) {real, imag} */,
  {32'h3fa3a460, 32'h41b1efef} /* (4, 27, 17) {real, imag} */,
  {32'h40bd0554, 32'h419e92b1} /* (4, 27, 16) {real, imag} */,
  {32'hc185d44e, 32'h41cc6bf8} /* (4, 27, 15) {real, imag} */,
  {32'hc1570f3e, 32'h41e2ac0c} /* (4, 27, 14) {real, imag} */,
  {32'h4085ebc2, 32'h420fb5ad} /* (4, 27, 13) {real, imag} */,
  {32'h415d053e, 32'h4209965a} /* (4, 27, 12) {real, imag} */,
  {32'h405881c0, 32'h41f40ba0} /* (4, 27, 11) {real, imag} */,
  {32'hc19e3360, 32'h4181e10e} /* (4, 27, 10) {real, imag} */,
  {32'hc2154351, 32'hbf42a2fc} /* (4, 27, 9) {real, imag} */,
  {32'hc1a99657, 32'hc11bd661} /* (4, 27, 8) {real, imag} */,
  {32'h403b5258, 32'hc180f149} /* (4, 27, 7) {real, imag} */,
  {32'h4111f78b, 32'hc0b5a6ae} /* (4, 27, 6) {real, imag} */,
  {32'h412a69e1, 32'hc189df8c} /* (4, 27, 5) {real, imag} */,
  {32'h3f8a1564, 32'hc1950eb7} /* (4, 27, 4) {real, imag} */,
  {32'hc016f87a, 32'hc181cf68} /* (4, 27, 3) {real, imag} */,
  {32'h41986171, 32'hc1cd9b60} /* (4, 27, 2) {real, imag} */,
  {32'h4114b670, 32'hc1be5296} /* (4, 27, 1) {real, imag} */,
  {32'hbf7aa040, 32'hc1bdf476} /* (4, 27, 0) {real, imag} */,
  {32'h3fe64d18, 32'h4094fb12} /* (4, 26, 31) {real, imag} */,
  {32'hbfa30400, 32'h40eff7a5} /* (4, 26, 30) {real, imag} */,
  {32'hc0f7f208, 32'h4184cda9} /* (4, 26, 29) {real, imag} */,
  {32'h3fd72b80, 32'h41a2033e} /* (4, 26, 28) {real, imag} */,
  {32'h417cea49, 32'h4066fd7f} /* (4, 26, 27) {real, imag} */,
  {32'h413f20a6, 32'hc1b33cb9} /* (4, 26, 26) {real, imag} */,
  {32'h417bf095, 32'h40c68d68} /* (4, 26, 25) {real, imag} */,
  {32'h41466d6b, 32'h411fb678} /* (4, 26, 24) {real, imag} */,
  {32'hbfa09c28, 32'hc0c99be8} /* (4, 26, 23) {real, imag} */,
  {32'hc197c4c7, 32'hc180eade} /* (4, 26, 22) {real, imag} */,
  {32'hc17c0204, 32'hc0412658} /* (4, 26, 21) {real, imag} */,
  {32'hc0bdaa5c, 32'h41869a00} /* (4, 26, 20) {real, imag} */,
  {32'hc0407fb5, 32'h41102567} /* (4, 26, 19) {real, imag} */,
  {32'h416736ee, 32'hc08f7b27} /* (4, 26, 18) {real, imag} */,
  {32'hc1386818, 32'hbf2c9554} /* (4, 26, 17) {real, imag} */,
  {32'hc1810c44, 32'h40e6bcfd} /* (4, 26, 16) {real, imag} */,
  {32'hc1546d57, 32'h41409fcc} /* (4, 26, 15) {real, imag} */,
  {32'hc18ebda0, 32'h41acf746} /* (4, 26, 14) {real, imag} */,
  {32'hc1911cca, 32'h41b4e106} /* (4, 26, 13) {real, imag} */,
  {32'hc16e943d, 32'h415320cb} /* (4, 26, 12) {real, imag} */,
  {32'hc03fc0e5, 32'h3f251830} /* (4, 26, 11) {real, imag} */,
  {32'hc189f768, 32'h40cb4c49} /* (4, 26, 10) {real, imag} */,
  {32'hc07c38e7, 32'h412aad12} /* (4, 26, 9) {real, imag} */,
  {32'h40915f5d, 32'h41857bfe} /* (4, 26, 8) {real, imag} */,
  {32'h40f7d80c, 32'h402017bc} /* (4, 26, 7) {real, imag} */,
  {32'h40728e68, 32'hc17fd49a} /* (4, 26, 6) {real, imag} */,
  {32'hc1355900, 32'hc15453a1} /* (4, 26, 5) {real, imag} */,
  {32'hc08ce92d, 32'hc007516e} /* (4, 26, 4) {real, imag} */,
  {32'hc0dbe23a, 32'h40c94d9c} /* (4, 26, 3) {real, imag} */,
  {32'hc13588fb, 32'h40607074} /* (4, 26, 2) {real, imag} */,
  {32'h40874828, 32'hc193a0b2} /* (4, 26, 1) {real, imag} */,
  {32'h41345bcc, 32'hc1aab954} /* (4, 26, 0) {real, imag} */,
  {32'hc0de3b8a, 32'hbffd69a2} /* (4, 25, 31) {real, imag} */,
  {32'hc18d5c86, 32'hc06f30c2} /* (4, 25, 30) {real, imag} */,
  {32'hc0b650fe, 32'h40edc08a} /* (4, 25, 29) {real, imag} */,
  {32'h3f780bd0, 32'h40372f88} /* (4, 25, 28) {real, imag} */,
  {32'h40bd25ef, 32'hc16a7e4e} /* (4, 25, 27) {real, imag} */,
  {32'hc13b3172, 32'hc15e7277} /* (4, 25, 26) {real, imag} */,
  {32'hc0b21a5b, 32'hc13cee39} /* (4, 25, 25) {real, imag} */,
  {32'hbf99dbc8, 32'hc13ebe5e} /* (4, 25, 24) {real, imag} */,
  {32'h41121574, 32'hc05e6df0} /* (4, 25, 23) {real, imag} */,
  {32'hc0018c5c, 32'h412ceaee} /* (4, 25, 22) {real, imag} */,
  {32'h3fa96fc0, 32'h4087f96c} /* (4, 25, 21) {real, imag} */,
  {32'h41ab0f4b, 32'h416bacaf} /* (4, 25, 20) {real, imag} */,
  {32'h40a7285d, 32'h41436fbc} /* (4, 25, 19) {real, imag} */,
  {32'hc0566474, 32'h418a6272} /* (4, 25, 18) {real, imag} */,
  {32'h418d5469, 32'h414414f7} /* (4, 25, 17) {real, imag} */,
  {32'h41471432, 32'hc099c482} /* (4, 25, 16) {real, imag} */,
  {32'h4079dda6, 32'hc04faad2} /* (4, 25, 15) {real, imag} */,
  {32'hc126f450, 32'h411a9fd3} /* (4, 25, 14) {real, imag} */,
  {32'hc13096f4, 32'h4186f3d7} /* (4, 25, 13) {real, imag} */,
  {32'hc085090c, 32'h3fbd7224} /* (4, 25, 12) {real, imag} */,
  {32'hc0c31130, 32'hc1785e0d} /* (4, 25, 11) {real, imag} */,
  {32'h3ef84a41, 32'hc1cb958b} /* (4, 25, 10) {real, imag} */,
  {32'h4118e2f1, 32'hc19d7cf2} /* (4, 25, 9) {real, imag} */,
  {32'h40e3faee, 32'hc1629ea4} /* (4, 25, 8) {real, imag} */,
  {32'h4154bf18, 32'hc085ca30} /* (4, 25, 7) {real, imag} */,
  {32'h40bdd5fa, 32'h412ac1f2} /* (4, 25, 6) {real, imag} */,
  {32'hc0070930, 32'h41c91c84} /* (4, 25, 5) {real, imag} */,
  {32'h3fde3a28, 32'h413c1770} /* (4, 25, 4) {real, imag} */,
  {32'hbe7218c0, 32'hc0def794} /* (4, 25, 3) {real, imag} */,
  {32'h409dfd40, 32'h4122cd56} /* (4, 25, 2) {real, imag} */,
  {32'hc0075e40, 32'h406f0611} /* (4, 25, 1) {real, imag} */,
  {32'hc08530bb, 32'h40a4c822} /* (4, 25, 0) {real, imag} */,
  {32'h3fb99f3c, 32'hc0b46a33} /* (4, 24, 31) {real, imag} */,
  {32'hbfa6bcf0, 32'hc17f14b4} /* (4, 24, 30) {real, imag} */,
  {32'hc0284a70, 32'hc1a96c51} /* (4, 24, 29) {real, imag} */,
  {32'h4015ef0c, 32'hc136d2b1} /* (4, 24, 28) {real, imag} */,
  {32'hc13a9272, 32'hc178a52f} /* (4, 24, 27) {real, imag} */,
  {32'h3e4c6d00, 32'hc1237bec} /* (4, 24, 26) {real, imag} */,
  {32'h40e47438, 32'hc1596414} /* (4, 24, 25) {real, imag} */,
  {32'hc0edd9c4, 32'hc1a4e2da} /* (4, 24, 24) {real, imag} */,
  {32'hc16f4c7a, 32'hc0a6c792} /* (4, 24, 23) {real, imag} */,
  {32'hc082d1e0, 32'hc1080be2} /* (4, 24, 22) {real, imag} */,
  {32'hc12441b9, 32'hc0b54b5c} /* (4, 24, 21) {real, imag} */,
  {32'hc157f427, 32'h412950fb} /* (4, 24, 20) {real, imag} */,
  {32'h40462fa8, 32'hc066c86e} /* (4, 24, 19) {real, imag} */,
  {32'h40eb1c40, 32'hc164a956} /* (4, 24, 18) {real, imag} */,
  {32'h40278310, 32'h40eef661} /* (4, 24, 17) {real, imag} */,
  {32'hc0b0e2f1, 32'h41b6a9ed} /* (4, 24, 16) {real, imag} */,
  {32'h3f4d951c, 32'h41ec1b6c} /* (4, 24, 15) {real, imag} */,
  {32'h411615b0, 32'h40d1c69d} /* (4, 24, 14) {real, imag} */,
  {32'h40f6a3cc, 32'h40c397f4} /* (4, 24, 13) {real, imag} */,
  {32'h40616290, 32'h41c485be} /* (4, 24, 12) {real, imag} */,
  {32'hbfb3dd78, 32'h414fe77d} /* (4, 24, 11) {real, imag} */,
  {32'hbf24b6a0, 32'h3eb7f930} /* (4, 24, 10) {real, imag} */,
  {32'h3db7f640, 32'hc1310208} /* (4, 24, 9) {real, imag} */,
  {32'hc08273f4, 32'hc1ea7017} /* (4, 24, 8) {real, imag} */,
  {32'hc0d99600, 32'hc1d5c040} /* (4, 24, 7) {real, imag} */,
  {32'h4096347d, 32'hc201eb30} /* (4, 24, 6) {real, imag} */,
  {32'hc082f92b, 32'hc1f1145a} /* (4, 24, 5) {real, imag} */,
  {32'hc0edd894, 32'hc12247ac} /* (4, 24, 4) {real, imag} */,
  {32'hc0fac199, 32'hc164838e} /* (4, 24, 3) {real, imag} */,
  {32'hc1a1682c, 32'hc199ea2a} /* (4, 24, 2) {real, imag} */,
  {32'hc198ae9a, 32'hc1aba7ce} /* (4, 24, 1) {real, imag} */,
  {32'hc114b508, 32'hc1655a56} /* (4, 24, 0) {real, imag} */,
  {32'hc00300c1, 32'hc0750d87} /* (4, 23, 31) {real, imag} */,
  {32'hbf34e430, 32'hc09ee20b} /* (4, 23, 30) {real, imag} */,
  {32'hbfaf13b8, 32'h40179edb} /* (4, 23, 29) {real, imag} */,
  {32'h3fae54c4, 32'h410ba347} /* (4, 23, 28) {real, imag} */,
  {32'h41467aa0, 32'h41caa9c5} /* (4, 23, 27) {real, imag} */,
  {32'h41aeb01c, 32'h410564bd} /* (4, 23, 26) {real, imag} */,
  {32'h4181b745, 32'hc08cf028} /* (4, 23, 25) {real, imag} */,
  {32'h4140fad7, 32'h410c817c} /* (4, 23, 24) {real, imag} */,
  {32'h4005329e, 32'h403a94e0} /* (4, 23, 23) {real, imag} */,
  {32'h40a3e75f, 32'hbfbd59d4} /* (4, 23, 22) {real, imag} */,
  {32'h409de04d, 32'hbf828f90} /* (4, 23, 21) {real, imag} */,
  {32'hc0c16718, 32'hc12b0998} /* (4, 23, 20) {real, imag} */,
  {32'hc1731ebd, 32'hc0eedb5f} /* (4, 23, 19) {real, imag} */,
  {32'hc1acfafc, 32'hc0546964} /* (4, 23, 18) {real, imag} */,
  {32'hc17e0669, 32'h3f94cfa8} /* (4, 23, 17) {real, imag} */,
  {32'h41078eee, 32'h3e0c0e40} /* (4, 23, 16) {real, imag} */,
  {32'h413e4a9a, 32'h3eb96680} /* (4, 23, 15) {real, imag} */,
  {32'hbff04310, 32'h40c734aa} /* (4, 23, 14) {real, imag} */,
  {32'hc02366e3, 32'hbe491220} /* (4, 23, 13) {real, imag} */,
  {32'h3e5840e0, 32'hc1002787} /* (4, 23, 12) {real, imag} */,
  {32'hc0ffea34, 32'h3f8fa9c6} /* (4, 23, 11) {real, imag} */,
  {32'h40844dd9, 32'h40b118af} /* (4, 23, 10) {real, imag} */,
  {32'h41532aed, 32'h402c8f64} /* (4, 23, 9) {real, imag} */,
  {32'h4179d391, 32'h411a124d} /* (4, 23, 8) {real, imag} */,
  {32'h413f7f5a, 32'h417c3055} /* (4, 23, 7) {real, imag} */,
  {32'hc0ad06c2, 32'hbe07e3a0} /* (4, 23, 6) {real, imag} */,
  {32'hc103e1c7, 32'hbff27620} /* (4, 23, 5) {real, imag} */,
  {32'hc0d0aa7a, 32'h3f554040} /* (4, 23, 4) {real, imag} */,
  {32'h3ff89d86, 32'hc0d2b558} /* (4, 23, 3) {real, imag} */,
  {32'hc069d310, 32'hc0a2b18c} /* (4, 23, 2) {real, imag} */,
  {32'h3fb63970, 32'h410b0628} /* (4, 23, 1) {real, imag} */,
  {32'h40685f4d, 32'h40b09bd0} /* (4, 23, 0) {real, imag} */,
  {32'hc067901d, 32'h3fcbc264} /* (4, 22, 31) {real, imag} */,
  {32'hbed8e180, 32'hc0d20ee6} /* (4, 22, 30) {real, imag} */,
  {32'h40e31a4c, 32'h4035ce8c} /* (4, 22, 29) {real, imag} */,
  {32'h40a74f64, 32'h3f140868} /* (4, 22, 28) {real, imag} */,
  {32'h41020027, 32'h3fd7a632} /* (4, 22, 27) {real, imag} */,
  {32'hbf7dfca0, 32'h3f1f7dd4} /* (4, 22, 26) {real, imag} */,
  {32'hbe8671e8, 32'h3f7bba80} /* (4, 22, 25) {real, imag} */,
  {32'h4033dcdc, 32'h40a46698} /* (4, 22, 24) {real, imag} */,
  {32'hc027820b, 32'h3fed9eca} /* (4, 22, 23) {real, imag} */,
  {32'h409f7e34, 32'h407687af} /* (4, 22, 22) {real, imag} */,
  {32'h401152d4, 32'hbdce85a0} /* (4, 22, 21) {real, imag} */,
  {32'h407ced1c, 32'hc138241a} /* (4, 22, 20) {real, imag} */,
  {32'h41149639, 32'hc0d5f748} /* (4, 22, 19) {real, imag} */,
  {32'h411fab8b, 32'hc0cd9373} /* (4, 22, 18) {real, imag} */,
  {32'hbfbf45fc, 32'hc148d3ee} /* (4, 22, 17) {real, imag} */,
  {32'hc0b75932, 32'hc1a95224} /* (4, 22, 16) {real, imag} */,
  {32'h4065b879, 32'hc13221d6} /* (4, 22, 15) {real, imag} */,
  {32'hc00f74c8, 32'hc13146f4} /* (4, 22, 14) {real, imag} */,
  {32'h3f90459e, 32'hc15921dc} /* (4, 22, 13) {real, imag} */,
  {32'hc0bac51b, 32'hc15077e4} /* (4, 22, 12) {real, imag} */,
  {32'h3fb3a65e, 32'hc12335a7} /* (4, 22, 11) {real, imag} */,
  {32'h41704ce7, 32'hc0439e31} /* (4, 22, 10) {real, imag} */,
  {32'h40fe0ba2, 32'h40ea4f52} /* (4, 22, 9) {real, imag} */,
  {32'h40b33f62, 32'h410eeb7a} /* (4, 22, 8) {real, imag} */,
  {32'h40fb3cd2, 32'h40cde41c} /* (4, 22, 7) {real, imag} */,
  {32'h40857630, 32'hc0cbab0e} /* (4, 22, 6) {real, imag} */,
  {32'h4182763c, 32'hc06873a8} /* (4, 22, 5) {real, imag} */,
  {32'h4149bb1f, 32'hc029dda4} /* (4, 22, 4) {real, imag} */,
  {32'h40ae55de, 32'hc01ea718} /* (4, 22, 3) {real, imag} */,
  {32'hc0ecfaa8, 32'hc0e4bca8} /* (4, 22, 2) {real, imag} */,
  {32'hc119411a, 32'hc0fbb7af} /* (4, 22, 1) {real, imag} */,
  {32'hc0a2417a, 32'h4062e5c8} /* (4, 22, 0) {real, imag} */,
  {32'h3f9db4fa, 32'hc0889132} /* (4, 21, 31) {real, imag} */,
  {32'hbf7d8558, 32'hc05b9cf4} /* (4, 21, 30) {real, imag} */,
  {32'hc0f19d0d, 32'hc0c42683} /* (4, 21, 29) {real, imag} */,
  {32'hc0e492b1, 32'hc145b960} /* (4, 21, 28) {real, imag} */,
  {32'hc119b646, 32'hc0a4c520} /* (4, 21, 27) {real, imag} */,
  {32'hc10900b5, 32'hbfaa8640} /* (4, 21, 26) {real, imag} */,
  {32'hc0f99714, 32'h3fb7a7ac} /* (4, 21, 25) {real, imag} */,
  {32'hc0c96d32, 32'hc046945c} /* (4, 21, 24) {real, imag} */,
  {32'hc13bb531, 32'hc0e763c6} /* (4, 21, 23) {real, imag} */,
  {32'hc152931c, 32'hc09ef7d2} /* (4, 21, 22) {real, imag} */,
  {32'hc0e65420, 32'hbf78af90} /* (4, 21, 21) {real, imag} */,
  {32'hc04810df, 32'hc0923a8d} /* (4, 21, 20) {real, imag} */,
  {32'hc0f02be2, 32'hbf3b6a80} /* (4, 21, 19) {real, imag} */,
  {32'hbfd3eb80, 32'h3ff88a24} /* (4, 21, 18) {real, imag} */,
  {32'h406dd9f0, 32'h3f494500} /* (4, 21, 17) {real, imag} */,
  {32'h4134472d, 32'hc0b8af6f} /* (4, 21, 16) {real, imag} */,
  {32'h414b3481, 32'h3f9a0559} /* (4, 21, 15) {real, imag} */,
  {32'h413559d7, 32'h4119a135} /* (4, 21, 14) {real, imag} */,
  {32'hc02195ba, 32'h410947b0} /* (4, 21, 13) {real, imag} */,
  {32'hc02fc332, 32'h412e87ea} /* (4, 21, 12) {real, imag} */,
  {32'h407fa477, 32'h40b977db} /* (4, 21, 11) {real, imag} */,
  {32'hc0f34c6b, 32'hbfb3edc8} /* (4, 21, 10) {real, imag} */,
  {32'hc191afa8, 32'hc124ee1a} /* (4, 21, 9) {real, imag} */,
  {32'hc1789cb9, 32'hc0e07db5} /* (4, 21, 8) {real, imag} */,
  {32'hc16e9d4c, 32'hc098c7c1} /* (4, 21, 7) {real, imag} */,
  {32'hc01e3db5, 32'hc054ed36} /* (4, 21, 6) {real, imag} */,
  {32'h3fbc7aea, 32'h408fc14a} /* (4, 21, 5) {real, imag} */,
  {32'hc01e7fe2, 32'hc03d567a} /* (4, 21, 4) {real, imag} */,
  {32'hbf893a24, 32'hc0d4dc68} /* (4, 21, 3) {real, imag} */,
  {32'h408aca15, 32'hbf05a2a0} /* (4, 21, 2) {real, imag} */,
  {32'h407e5940, 32'h4083c803} /* (4, 21, 1) {real, imag} */,
  {32'h408181d9, 32'hbfb9408e} /* (4, 21, 0) {real, imag} */,
  {32'h40cbaa4b, 32'h40b224b2} /* (4, 20, 31) {real, imag} */,
  {32'h40ca71de, 32'hbfb38190} /* (4, 20, 30) {real, imag} */,
  {32'h40b8917b, 32'hc11b1c48} /* (4, 20, 29) {real, imag} */,
  {32'h3f5666c0, 32'hc10b85ea} /* (4, 20, 28) {real, imag} */,
  {32'hc01843f5, 32'hc09862be} /* (4, 20, 27) {real, imag} */,
  {32'hc0110cd2, 32'hbeb28410} /* (4, 20, 26) {real, imag} */,
  {32'hc02b5bcf, 32'hbffd462c} /* (4, 20, 25) {real, imag} */,
  {32'hc0cbf84e, 32'h409ba372} /* (4, 20, 24) {real, imag} */,
  {32'h3fad6624, 32'h410f2538} /* (4, 20, 23) {real, imag} */,
  {32'hc09cd734, 32'h409fe098} /* (4, 20, 22) {real, imag} */,
  {32'hc14b033f, 32'h406f4147} /* (4, 20, 21) {real, imag} */,
  {32'hc02f2db6, 32'h40a8cede} /* (4, 20, 20) {real, imag} */,
  {32'h40fb7206, 32'h4006ad5b} /* (4, 20, 19) {real, imag} */,
  {32'h40e41ff4, 32'h406c6c10} /* (4, 20, 18) {real, imag} */,
  {32'h410c257a, 32'hbf5b9820} /* (4, 20, 17) {real, imag} */,
  {32'h40cbbe30, 32'hc0b11115} /* (4, 20, 16) {real, imag} */,
  {32'h40173f7a, 32'h3f0deaca} /* (4, 20, 15) {real, imag} */,
  {32'h40858f73, 32'hc090933c} /* (4, 20, 14) {real, imag} */,
  {32'hc07851d4, 32'hc11d11ad} /* (4, 20, 13) {real, imag} */,
  {32'h3f5494b0, 32'hc087e8d1} /* (4, 20, 12) {real, imag} */,
  {32'h41026458, 32'h3ffed063} /* (4, 20, 11) {real, imag} */,
  {32'h40191cba, 32'hc0e0909d} /* (4, 20, 10) {real, imag} */,
  {32'hc0f8c11b, 32'hc139e2f5} /* (4, 20, 9) {real, imag} */,
  {32'hc0a0b12e, 32'hc004813c} /* (4, 20, 8) {real, imag} */,
  {32'hc0e4c25a, 32'hc01704fc} /* (4, 20, 7) {real, imag} */,
  {32'h402bc0b8, 32'h40412102} /* (4, 20, 6) {real, imag} */,
  {32'h40efe4a4, 32'hbf30c564} /* (4, 20, 5) {real, imag} */,
  {32'h4105cecc, 32'hc00a7962} /* (4, 20, 4) {real, imag} */,
  {32'h3fb7969c, 32'h402dda74} /* (4, 20, 3) {real, imag} */,
  {32'hc01b4c40, 32'h4059bcdc} /* (4, 20, 2) {real, imag} */,
  {32'h406ecfc1, 32'h3ff812f8} /* (4, 20, 1) {real, imag} */,
  {32'h4038f9f4, 32'h4025ba72} /* (4, 20, 0) {real, imag} */,
  {32'h3fe2288c, 32'h405301a1} /* (4, 19, 31) {real, imag} */,
  {32'hc010d2e0, 32'hc048a339} /* (4, 19, 30) {real, imag} */,
  {32'hc0bb869c, 32'hc02045a7} /* (4, 19, 29) {real, imag} */,
  {32'h40533cee, 32'h3e2dc630} /* (4, 19, 28) {real, imag} */,
  {32'hc025fce4, 32'hbf8c90bc} /* (4, 19, 27) {real, imag} */,
  {32'hbf5fef20, 32'h3f9ede74} /* (4, 19, 26) {real, imag} */,
  {32'h3fab6ed8, 32'h405f86af} /* (4, 19, 25) {real, imag} */,
  {32'h400df145, 32'h405fb924} /* (4, 19, 24) {real, imag} */,
  {32'h3f6521e0, 32'hc08369fe} /* (4, 19, 23) {real, imag} */,
  {32'h3ff21910, 32'h3f851ef6} /* (4, 19, 22) {real, imag} */,
  {32'h40c2d760, 32'hbdef7700} /* (4, 19, 21) {real, imag} */,
  {32'h40da115a, 32'hc056174d} /* (4, 19, 20) {real, imag} */,
  {32'h40b3e042, 32'hc09930f7} /* (4, 19, 19) {real, imag} */,
  {32'h3ec18a60, 32'hc03ce480} /* (4, 19, 18) {real, imag} */,
  {32'hc018c038, 32'hbf0c5194} /* (4, 19, 17) {real, imag} */,
  {32'hbf9bed00, 32'h40ac0bdd} /* (4, 19, 16) {real, imag} */,
  {32'hc1037a2a, 32'h407a1e54} /* (4, 19, 15) {real, imag} */,
  {32'hc11ef7df, 32'hbfd0b3cd} /* (4, 19, 14) {real, imag} */,
  {32'hbd6e2680, 32'hc12e57c0} /* (4, 19, 13) {real, imag} */,
  {32'h40cc039c, 32'hbf903bf8} /* (4, 19, 12) {real, imag} */,
  {32'h40c54bd6, 32'h3fb9f1f2} /* (4, 19, 11) {real, imag} */,
  {32'h4103c4c4, 32'hbebf5020} /* (4, 19, 10) {real, imag} */,
  {32'h40a22093, 32'h409394b9} /* (4, 19, 9) {real, imag} */,
  {32'h40a6c15a, 32'h40cc8d34} /* (4, 19, 8) {real, imag} */,
  {32'hbf1e6b40, 32'h3e72e6f0} /* (4, 19, 7) {real, imag} */,
  {32'h3facd7f4, 32'h3f563160} /* (4, 19, 6) {real, imag} */,
  {32'h4119025a, 32'h3e41bf50} /* (4, 19, 5) {real, imag} */,
  {32'h408e1319, 32'h3e9d3818} /* (4, 19, 4) {real, imag} */,
  {32'hbe8231e0, 32'h40d6aa50} /* (4, 19, 3) {real, imag} */,
  {32'h402e5f84, 32'h40b9bcea} /* (4, 19, 2) {real, imag} */,
  {32'h402daae9, 32'hbf93595e} /* (4, 19, 1) {real, imag} */,
  {32'h3f7fbc48, 32'hc06e4eec} /* (4, 19, 0) {real, imag} */,
  {32'hbf3c7fb8, 32'h3f08a1dc} /* (4, 18, 31) {real, imag} */,
  {32'hbc994a00, 32'h3fa2aada} /* (4, 18, 30) {real, imag} */,
  {32'hc0d5ee04, 32'hbf82c692} /* (4, 18, 29) {real, imag} */,
  {32'hc13ec7ec, 32'hbf9e883c} /* (4, 18, 28) {real, imag} */,
  {32'hc08236c8, 32'h40131745} /* (4, 18, 27) {real, imag} */,
  {32'h3fbbf828, 32'h40802a70} /* (4, 18, 26) {real, imag} */,
  {32'hc008aa40, 32'hbe67bd20} /* (4, 18, 25) {real, imag} */,
  {32'hc02457fc, 32'hc0554abc} /* (4, 18, 24) {real, imag} */,
  {32'hc02d7b18, 32'h3fe8b4ac} /* (4, 18, 23) {real, imag} */,
  {32'h40901f47, 32'h409898fc} /* (4, 18, 22) {real, imag} */,
  {32'h40bf9c02, 32'h3fb103a8} /* (4, 18, 21) {real, imag} */,
  {32'hbe0abb80, 32'h402575b6} /* (4, 18, 20) {real, imag} */,
  {32'hc0b0774e, 32'hbffc9a08} /* (4, 18, 19) {real, imag} */,
  {32'hbf13aea0, 32'h3f429390} /* (4, 18, 18) {real, imag} */,
  {32'h4054e3ec, 32'h410602b9} /* (4, 18, 17) {real, imag} */,
  {32'h40034b90, 32'h400702a3} /* (4, 18, 16) {real, imag} */,
  {32'h401c7900, 32'hc04d10f6} /* (4, 18, 15) {real, imag} */,
  {32'h40424a8c, 32'hc0384120} /* (4, 18, 14) {real, imag} */,
  {32'hc097f6de, 32'h3dda7d80} /* (4, 18, 13) {real, imag} */,
  {32'hc0d65320, 32'hbfb09c6e} /* (4, 18, 12) {real, imag} */,
  {32'hc024a242, 32'h3fdead38} /* (4, 18, 11) {real, imag} */,
  {32'hc0494b32, 32'hc078d344} /* (4, 18, 10) {real, imag} */,
  {32'hc0bdb3ab, 32'hc115a46a} /* (4, 18, 9) {real, imag} */,
  {32'hc0cda7c6, 32'hc0dd21b9} /* (4, 18, 8) {real, imag} */,
  {32'hc02743b0, 32'hc0c078c0} /* (4, 18, 7) {real, imag} */,
  {32'hbfc3504c, 32'hc0c5f61e} /* (4, 18, 6) {real, imag} */,
  {32'h403a9cdc, 32'hc04d2b00} /* (4, 18, 5) {real, imag} */,
  {32'hc02435a0, 32'hbf8839b0} /* (4, 18, 4) {real, imag} */,
  {32'hc0b38694, 32'hc088cff3} /* (4, 18, 3) {real, imag} */,
  {32'hc0505e20, 32'hc0ec5ff9} /* (4, 18, 2) {real, imag} */,
  {32'h40b8f16d, 32'hbf9aaede} /* (4, 18, 1) {real, imag} */,
  {32'h3fd53f00, 32'hbd8b4660} /* (4, 18, 0) {real, imag} */,
  {32'h4005f58f, 32'hc07576c3} /* (4, 17, 31) {real, imag} */,
  {32'h40faf4ba, 32'hbff0fa90} /* (4, 17, 30) {real, imag} */,
  {32'h40474608, 32'h40a73a9a} /* (4, 17, 29) {real, imag} */,
  {32'h3f058ce0, 32'h4084e21c} /* (4, 17, 28) {real, imag} */,
  {32'h3fae0c2c, 32'hc02789bf} /* (4, 17, 27) {real, imag} */,
  {32'hc00f1e7a, 32'hc0156328} /* (4, 17, 26) {real, imag} */,
  {32'hc013f794, 32'h3e947d28} /* (4, 17, 25) {real, imag} */,
  {32'hc09d5758, 32'h3f98aad4} /* (4, 17, 24) {real, imag} */,
  {32'hc03f9814, 32'hbfba0fe8} /* (4, 17, 23) {real, imag} */,
  {32'hc099cb3c, 32'hbf7b4768} /* (4, 17, 22) {real, imag} */,
  {32'hc02814be, 32'h3dcefb00} /* (4, 17, 21) {real, imag} */,
  {32'hc0659391, 32'h3f46d190} /* (4, 17, 20) {real, imag} */,
  {32'h3e954350, 32'h3e591a20} /* (4, 17, 19) {real, imag} */,
  {32'h40862b76, 32'hc0e7d6f8} /* (4, 17, 18) {real, imag} */,
  {32'h404d5c09, 32'hbfd7eb08} /* (4, 17, 17) {real, imag} */,
  {32'hbf7b20ec, 32'hc0004560} /* (4, 17, 16) {real, imag} */,
  {32'hc08c8de6, 32'hc0a6aac4} /* (4, 17, 15) {real, imag} */,
  {32'hc0913916, 32'hbfdb0b12} /* (4, 17, 14) {real, imag} */,
  {32'hc081ce84, 32'hc0249242} /* (4, 17, 13) {real, imag} */,
  {32'hbfcd0076, 32'hbf84f7c8} /* (4, 17, 12) {real, imag} */,
  {32'hbdf69fb0, 32'h3f9db254} /* (4, 17, 11) {real, imag} */,
  {32'hbfe4a60e, 32'hc1118eb7} /* (4, 17, 10) {real, imag} */,
  {32'h3fdfcca0, 32'hc066fb0c} /* (4, 17, 9) {real, imag} */,
  {32'h40618204, 32'h4034db74} /* (4, 17, 8) {real, imag} */,
  {32'h40859ad8, 32'hc01efbd6} /* (4, 17, 7) {real, imag} */,
  {32'h40ad7ce6, 32'hc06982d0} /* (4, 17, 6) {real, imag} */,
  {32'hbf602cd0, 32'hc0e03f2a} /* (4, 17, 5) {real, imag} */,
  {32'hc0a88776, 32'h3f1a8068} /* (4, 17, 4) {real, imag} */,
  {32'hc019bea8, 32'h40825510} /* (4, 17, 3) {real, imag} */,
  {32'hc0177c88, 32'h4081293f} /* (4, 17, 2) {real, imag} */,
  {32'hbf50b3bc, 32'h3f9511d6} /* (4, 17, 1) {real, imag} */,
  {32'h40091570, 32'hbf7302c4} /* (4, 17, 0) {real, imag} */,
  {32'hc008fd66, 32'hbf8dfea0} /* (4, 16, 31) {real, imag} */,
  {32'h40706600, 32'h3fd7c220} /* (4, 16, 30) {real, imag} */,
  {32'h40b86172, 32'h40bbaed0} /* (4, 16, 29) {real, imag} */,
  {32'h40a41d1e, 32'h410a34c4} /* (4, 16, 28) {real, imag} */,
  {32'h40410668, 32'h40347480} /* (4, 16, 27) {real, imag} */,
  {32'hbf81e4c0, 32'h3f027c00} /* (4, 16, 26) {real, imag} */,
  {32'hbfda7838, 32'h3f0bf7e0} /* (4, 16, 25) {real, imag} */,
  {32'h3fd3c3e2, 32'hc092b914} /* (4, 16, 24) {real, imag} */,
  {32'h4031017a, 32'h3eb62d80} /* (4, 16, 23) {real, imag} */,
  {32'h3fbf94b0, 32'hbf700600} /* (4, 16, 22) {real, imag} */,
  {32'hc0ae1ebc, 32'h40503770} /* (4, 16, 21) {real, imag} */,
  {32'hc09d93f2, 32'h410381a6} /* (4, 16, 20) {real, imag} */,
  {32'hc10bdb54, 32'h40a62d9c} /* (4, 16, 19) {real, imag} */,
  {32'hbfce4260, 32'h40835344} /* (4, 16, 18) {real, imag} */,
  {32'h40778792, 32'hbfda842c} /* (4, 16, 17) {real, imag} */,
  {32'h4010345a, 32'hc06f69f2} /* (4, 16, 16) {real, imag} */,
  {32'h3eb9927c, 32'h3f3593e0} /* (4, 16, 15) {real, imag} */,
  {32'hbfc33190, 32'hbe1d4680} /* (4, 16, 14) {real, imag} */,
  {32'hbfc67dd0, 32'h401c4f20} /* (4, 16, 13) {real, imag} */,
  {32'h3fe783c8, 32'h40742cf0} /* (4, 16, 12) {real, imag} */,
  {32'h3f638f30, 32'h40812390} /* (4, 16, 11) {real, imag} */,
  {32'h40409475, 32'h403bce10} /* (4, 16, 10) {real, imag} */,
  {32'hbf2bdf20, 32'h3f63dd90} /* (4, 16, 9) {real, imag} */,
  {32'hbfdd7a0c, 32'h4034fae4} /* (4, 16, 8) {real, imag} */,
  {32'hc0b18759, 32'h3f752a20} /* (4, 16, 7) {real, imag} */,
  {32'h3df7ff00, 32'h3f6d1ae0} /* (4, 16, 6) {real, imag} */,
  {32'h40909c9d, 32'h400d5230} /* (4, 16, 5) {real, imag} */,
  {32'hbe61ed00, 32'h3e505f00} /* (4, 16, 4) {real, imag} */,
  {32'h3cf98100, 32'h4001c580} /* (4, 16, 3) {real, imag} */,
  {32'h40a751ae, 32'h3f884cb0} /* (4, 16, 2) {real, imag} */,
  {32'h409018d0, 32'h3fcaf120} /* (4, 16, 1) {real, imag} */,
  {32'hbf4a57e0, 32'h405ffc9c} /* (4, 16, 0) {real, imag} */,
  {32'hbfd04726, 32'h401bdee3} /* (4, 15, 31) {real, imag} */,
  {32'hc0d4cb02, 32'h3f5b4b20} /* (4, 15, 30) {real, imag} */,
  {32'hc00389b8, 32'hc05558f4} /* (4, 15, 29) {real, imag} */,
  {32'h40d618f0, 32'hbf0f0ee4} /* (4, 15, 28) {real, imag} */,
  {32'hbf0aa858, 32'h409eb210} /* (4, 15, 27) {real, imag} */,
  {32'hc0b49b07, 32'h40644ca8} /* (4, 15, 26) {real, imag} */,
  {32'hc0291d6c, 32'hc0796ec5} /* (4, 15, 25) {real, imag} */,
  {32'hc08006b8, 32'hc0947745} /* (4, 15, 24) {real, imag} */,
  {32'hbfe333d8, 32'h3f1f41d0} /* (4, 15, 23) {real, imag} */,
  {32'h3f0224e0, 32'h401b35da} /* (4, 15, 22) {real, imag} */,
  {32'hbe43e120, 32'h403e7b48} /* (4, 15, 21) {real, imag} */,
  {32'h3f9038d6, 32'hbfa82b48} /* (4, 15, 20) {real, imag} */,
  {32'h41049afa, 32'hbff90d84} /* (4, 15, 19) {real, imag} */,
  {32'h4084e1a6, 32'h400fcb00} /* (4, 15, 18) {real, imag} */,
  {32'hbf4d911c, 32'h40027f84} /* (4, 15, 17) {real, imag} */,
  {32'h40b59d52, 32'h401b9cb0} /* (4, 15, 16) {real, imag} */,
  {32'h40aef980, 32'hbedb5a40} /* (4, 15, 15) {real, imag} */,
  {32'h405744e4, 32'hc04c2577} /* (4, 15, 14) {real, imag} */,
  {32'h403edc40, 32'hc052acfe} /* (4, 15, 13) {real, imag} */,
  {32'hc00d035d, 32'hbfebee78} /* (4, 15, 12) {real, imag} */,
  {32'hc05252aa, 32'hc06cb9ca} /* (4, 15, 11) {real, imag} */,
  {32'hc05b9a6f, 32'hbf3c2ce0} /* (4, 15, 10) {real, imag} */,
  {32'hc107d2b4, 32'hc026fdfc} /* (4, 15, 9) {real, imag} */,
  {32'hc00bf83c, 32'hc05e3514} /* (4, 15, 8) {real, imag} */,
  {32'h40ba5850, 32'hc03fb79a} /* (4, 15, 7) {real, imag} */,
  {32'h40538654, 32'hbedb5980} /* (4, 15, 6) {real, imag} */,
  {32'h3fc5bfa8, 32'hc04797fb} /* (4, 15, 5) {real, imag} */,
  {32'h3e880f58, 32'hc0a8b76d} /* (4, 15, 4) {real, imag} */,
  {32'hc0ccc4c8, 32'h409da720} /* (4, 15, 3) {real, imag} */,
  {32'hc107091e, 32'h411f8140} /* (4, 15, 2) {real, imag} */,
  {32'hc0b41efa, 32'h401b2ef5} /* (4, 15, 1) {real, imag} */,
  {32'hbf740a42, 32'h3f879462} /* (4, 15, 0) {real, imag} */,
  {32'h409d64b5, 32'h401debe9} /* (4, 14, 31) {real, imag} */,
  {32'hbecb05a0, 32'h4039fd83} /* (4, 14, 30) {real, imag} */,
  {32'h40146278, 32'hc0216a47} /* (4, 14, 29) {real, imag} */,
  {32'h40880338, 32'h4066e11e} /* (4, 14, 28) {real, imag} */,
  {32'h3f3b9da0, 32'h411edaaf} /* (4, 14, 27) {real, imag} */,
  {32'h3f9e2af8, 32'h40bbdab8} /* (4, 14, 26) {real, imag} */,
  {32'hbf813340, 32'h40496f52} /* (4, 14, 25) {real, imag} */,
  {32'h408457be, 32'h3db82d80} /* (4, 14, 24) {real, imag} */,
  {32'h40930054, 32'hbf188798} /* (4, 14, 23) {real, imag} */,
  {32'h401fbee2, 32'h3fa2f7cf} /* (4, 14, 22) {real, imag} */,
  {32'hbf6c3224, 32'h404085e0} /* (4, 14, 21) {real, imag} */,
  {32'h3cae0c00, 32'hbe16f560} /* (4, 14, 20) {real, imag} */,
  {32'h3e29ec40, 32'hbda31980} /* (4, 14, 19) {real, imag} */,
  {32'hc0b8b61c, 32'hbe2e3140} /* (4, 14, 18) {real, imag} */,
  {32'hc0b447c2, 32'hc0210d44} /* (4, 14, 17) {real, imag} */,
  {32'hbf471240, 32'hbd7654c0} /* (4, 14, 16) {real, imag} */,
  {32'h40702750, 32'hc0c73bad} /* (4, 14, 15) {real, imag} */,
  {32'hc0f963ec, 32'hbfb41c00} /* (4, 14, 14) {real, imag} */,
  {32'hc163c985, 32'hbf5912b0} /* (4, 14, 13) {real, imag} */,
  {32'hc0d9a56a, 32'h401083c7} /* (4, 14, 12) {real, imag} */,
  {32'hc0a645b9, 32'h4091cd8e} /* (4, 14, 11) {real, imag} */,
  {32'hc0725f4a, 32'h3f2c3d90} /* (4, 14, 10) {real, imag} */,
  {32'h3fa1c24c, 32'h3f9fd5d0} /* (4, 14, 9) {real, imag} */,
  {32'h3fdd61c8, 32'h3fa74ae4} /* (4, 14, 8) {real, imag} */,
  {32'h409b72f0, 32'h3f2ab184} /* (4, 14, 7) {real, imag} */,
  {32'h404c8222, 32'hbeb1d628} /* (4, 14, 6) {real, imag} */,
  {32'h409795ca, 32'hbee2107c} /* (4, 14, 5) {real, imag} */,
  {32'h408ba608, 32'h402db0c8} /* (4, 14, 4) {real, imag} */,
  {32'h4014787c, 32'hc004e69a} /* (4, 14, 3) {real, imag} */,
  {32'h40794520, 32'hbff3077c} /* (4, 14, 2) {real, imag} */,
  {32'h40a2edff, 32'hc00bc051} /* (4, 14, 1) {real, imag} */,
  {32'h40c84028, 32'hbf2e2f34} /* (4, 14, 0) {real, imag} */,
  {32'hc0728c06, 32'h40d5e8e0} /* (4, 13, 31) {real, imag} */,
  {32'hc09fb446, 32'h40082317} /* (4, 13, 30) {real, imag} */,
  {32'hbe9582d8, 32'h3fbe92ae} /* (4, 13, 29) {real, imag} */,
  {32'hbe8dbeb0, 32'hc0ec5e46} /* (4, 13, 28) {real, imag} */,
  {32'h3f4566c2, 32'hc08b50b3} /* (4, 13, 27) {real, imag} */,
  {32'h4090ffc3, 32'hbfcf1c4c} /* (4, 13, 26) {real, imag} */,
  {32'h40ad37c6, 32'hc09217ee} /* (4, 13, 25) {real, imag} */,
  {32'hc0948274, 32'h4015cd78} /* (4, 13, 24) {real, imag} */,
  {32'hc1266ac2, 32'h40844b96} /* (4, 13, 23) {real, imag} */,
  {32'hc0831be4, 32'h4003a16b} /* (4, 13, 22) {real, imag} */,
  {32'hbf1fd280, 32'h3e4fb900} /* (4, 13, 21) {real, imag} */,
  {32'hbd6b6340, 32'hc0eac59a} /* (4, 13, 20) {real, imag} */,
  {32'hc0c00656, 32'hc0dd242f} /* (4, 13, 19) {real, imag} */,
  {32'hc0d88fca, 32'hc0b2508c} /* (4, 13, 18) {real, imag} */,
  {32'h40327a48, 32'hc032edcd} /* (4, 13, 17) {real, imag} */,
  {32'hbedd7400, 32'hc0a5fe17} /* (4, 13, 16) {real, imag} */,
  {32'hbf67a938, 32'hc0d98e4a} /* (4, 13, 15) {real, imag} */,
  {32'h40570fec, 32'hbfa8892d} /* (4, 13, 14) {real, imag} */,
  {32'h4071f512, 32'hc11cd7a0} /* (4, 13, 13) {real, imag} */,
  {32'hc0938eb4, 32'hc1373e95} /* (4, 13, 12) {real, imag} */,
  {32'hbee344e8, 32'hc0849f42} /* (4, 13, 11) {real, imag} */,
  {32'h3f00ce38, 32'h4095ee0e} /* (4, 13, 10) {real, imag} */,
  {32'hc060b6ca, 32'h402adf42} /* (4, 13, 9) {real, imag} */,
  {32'hc0a6905e, 32'hc07383a0} /* (4, 13, 8) {real, imag} */,
  {32'hc0d21900, 32'hc02fb8e5} /* (4, 13, 7) {real, imag} */,
  {32'hbfcdcdac, 32'h3fbe8758} /* (4, 13, 6) {real, imag} */,
  {32'hc0bcfdaf, 32'h40c45bae} /* (4, 13, 5) {real, imag} */,
  {32'hc0f18f77, 32'h402a001b} /* (4, 13, 4) {real, imag} */,
  {32'hc0dfbd3e, 32'hc0826640} /* (4, 13, 3) {real, imag} */,
  {32'hc0d3a6ae, 32'h3f9764f8} /* (4, 13, 2) {real, imag} */,
  {32'hbf3cb054, 32'h406f3ca1} /* (4, 13, 1) {real, imag} */,
  {32'h3dd32ac0, 32'h40dd33d4} /* (4, 13, 0) {real, imag} */,
  {32'hbe8ade70, 32'h405db83f} /* (4, 12, 31) {real, imag} */,
  {32'h40c33e32, 32'hc07ebf3c} /* (4, 12, 30) {real, imag} */,
  {32'hc102239e, 32'hc0a8c9dd} /* (4, 12, 29) {real, imag} */,
  {32'hc194906c, 32'hc08050e2} /* (4, 12, 28) {real, imag} */,
  {32'hc0814262, 32'hc083914e} /* (4, 12, 27) {real, imag} */,
  {32'h408def3f, 32'hc07b6426} /* (4, 12, 26) {real, imag} */,
  {32'h3f938026, 32'hbf1bd5a8} /* (4, 12, 25) {real, imag} */,
  {32'h3e390d40, 32'hc0083db7} /* (4, 12, 24) {real, imag} */,
  {32'h4059fa22, 32'hbda2a280} /* (4, 12, 23) {real, imag} */,
  {32'hbee6cba8, 32'h40a643d4} /* (4, 12, 22) {real, imag} */,
  {32'h40aa88d2, 32'hc0964b64} /* (4, 12, 21) {real, imag} */,
  {32'h3ffe88a4, 32'hbfe503c6} /* (4, 12, 20) {real, imag} */,
  {32'hbfd56b52, 32'h4009ed9d} /* (4, 12, 19) {real, imag} */,
  {32'h3fedae90, 32'h4082a2e4} /* (4, 12, 18) {real, imag} */,
  {32'h4030bd26, 32'h40b364b0} /* (4, 12, 17) {real, imag} */,
  {32'h412664f4, 32'hbf8a3f5c} /* (4, 12, 16) {real, imag} */,
  {32'h40175a84, 32'h3f964a5b} /* (4, 12, 15) {real, imag} */,
  {32'hc058c9f4, 32'h40054cd0} /* (4, 12, 14) {real, imag} */,
  {32'hbeb41580, 32'hc03106cc} /* (4, 12, 13) {real, imag} */,
  {32'hc0d45be0, 32'hc0ad7267} /* (4, 12, 12) {real, imag} */,
  {32'hc0892148, 32'hbfde4ec3} /* (4, 12, 11) {real, imag} */,
  {32'hc01b1e56, 32'h40ff91ff} /* (4, 12, 10) {real, imag} */,
  {32'hbffe69ac, 32'h41375371} /* (4, 12, 9) {real, imag} */,
  {32'hc12805bb, 32'hbf9a3aa8} /* (4, 12, 8) {real, imag} */,
  {32'hc0ea8c1e, 32'hc00e0044} /* (4, 12, 7) {real, imag} */,
  {32'hbf011d60, 32'hbe860c70} /* (4, 12, 6) {real, imag} */,
  {32'h4049a164, 32'hc02411ff} /* (4, 12, 5) {real, imag} */,
  {32'h4076e4c0, 32'h408a629b} /* (4, 12, 4) {real, imag} */,
  {32'hc0ee972d, 32'h3ee2a260} /* (4, 12, 3) {real, imag} */,
  {32'hbfe4e338, 32'hc0cdd116} /* (4, 12, 2) {real, imag} */,
  {32'h3fdfcf3e, 32'hc144c919} /* (4, 12, 1) {real, imag} */,
  {32'hc02b22ac, 32'hc01fa8ca} /* (4, 12, 0) {real, imag} */,
  {32'h41038919, 32'hc0bb838a} /* (4, 11, 31) {real, imag} */,
  {32'h40b22d3f, 32'hc0b13a26} /* (4, 11, 30) {real, imag} */,
  {32'h404eafc6, 32'hc0f6e37b} /* (4, 11, 29) {real, imag} */,
  {32'h40b6a52b, 32'hc15c12a4} /* (4, 11, 28) {real, imag} */,
  {32'hbf8168f4, 32'hc1715efe} /* (4, 11, 27) {real, imag} */,
  {32'h4021b064, 32'hc12bc38a} /* (4, 11, 26) {real, imag} */,
  {32'h4055905f, 32'h40d9c901} /* (4, 11, 25) {real, imag} */,
  {32'h402c782b, 32'h4157a4eb} /* (4, 11, 24) {real, imag} */,
  {32'h410b258b, 32'h4096585e} /* (4, 11, 23) {real, imag} */,
  {32'h4139011a, 32'h40dc8f36} /* (4, 11, 22) {real, imag} */,
  {32'h40b1e5be, 32'h4011cb88} /* (4, 11, 21) {real, imag} */,
  {32'hc0dacbfc, 32'hc0732a1e} /* (4, 11, 20) {real, imag} */,
  {32'hc0c044c8, 32'hbeb9ca00} /* (4, 11, 19) {real, imag} */,
  {32'hc14034b4, 32'hc0b3d16f} /* (4, 11, 18) {real, imag} */,
  {32'hc0c1a044, 32'hc122629d} /* (4, 11, 17) {real, imag} */,
  {32'hbf90dbd8, 32'hbf3a3678} /* (4, 11, 16) {real, imag} */,
  {32'hc12dc5c1, 32'hbf10e072} /* (4, 11, 15) {real, imag} */,
  {32'hc11d3109, 32'hc0f6db46} /* (4, 11, 14) {real, imag} */,
  {32'hc13c565e, 32'h3f93dcc4} /* (4, 11, 13) {real, imag} */,
  {32'hbfd187b4, 32'h400aafa6} /* (4, 11, 12) {real, imag} */,
  {32'hc0bde630, 32'h40e55507} /* (4, 11, 11) {real, imag} */,
  {32'hbf150b88, 32'hbf58b520} /* (4, 11, 10) {real, imag} */,
  {32'h410df029, 32'h4082cb19} /* (4, 11, 9) {real, imag} */,
  {32'h401c3e0c, 32'h40438c1e} /* (4, 11, 8) {real, imag} */,
  {32'hbf9b4980, 32'h403f1f9e} /* (4, 11, 7) {real, imag} */,
  {32'h4126caf7, 32'h4071acc6} /* (4, 11, 6) {real, imag} */,
  {32'h403c1c0d, 32'h40363b44} /* (4, 11, 5) {real, imag} */,
  {32'h40d3a8a1, 32'h41406e10} /* (4, 11, 4) {real, imag} */,
  {32'h4117e65e, 32'h41541050} /* (4, 11, 3) {real, imag} */,
  {32'h41347a18, 32'hc085c0a0} /* (4, 11, 2) {real, imag} */,
  {32'h41200422, 32'hc121e7ac} /* (4, 11, 1) {real, imag} */,
  {32'h3fce45f4, 32'hc09ea046} /* (4, 11, 0) {real, imag} */,
  {32'h3d8c4160, 32'hc06d8754} /* (4, 10, 31) {real, imag} */,
  {32'hc0c01a92, 32'hc1077c1a} /* (4, 10, 30) {real, imag} */,
  {32'h3eb13fc8, 32'hc0b5f646} /* (4, 10, 29) {real, imag} */,
  {32'hc08b5ee4, 32'hc102c75e} /* (4, 10, 28) {real, imag} */,
  {32'hc1af5d88, 32'h40e20614} /* (4, 10, 27) {real, imag} */,
  {32'hc18be1fb, 32'h409afd92} /* (4, 10, 26) {real, imag} */,
  {32'h40160d9b, 32'hc122ccf2} /* (4, 10, 25) {real, imag} */,
  {32'h40a4754b, 32'hc1942e2f} /* (4, 10, 24) {real, imag} */,
  {32'hc0f1232e, 32'hc0b09726} /* (4, 10, 23) {real, imag} */,
  {32'hc110d37c, 32'hbfaf087e} /* (4, 10, 22) {real, imag} */,
  {32'h40ad6a1c, 32'hbf34fac4} /* (4, 10, 21) {real, imag} */,
  {32'h410ed5db, 32'h3fc9917c} /* (4, 10, 20) {real, imag} */,
  {32'h40675f7c, 32'h41072f85} /* (4, 10, 19) {real, imag} */,
  {32'h4094832e, 32'h402a96be} /* (4, 10, 18) {real, imag} */,
  {32'h40ff73af, 32'h40ca0a9c} /* (4, 10, 17) {real, imag} */,
  {32'hc0491b8c, 32'h410afa9c} /* (4, 10, 16) {real, imag} */,
  {32'hc0b2c210, 32'h4058741c} /* (4, 10, 15) {real, imag} */,
  {32'h3efd5380, 32'hbef83bb0} /* (4, 10, 14) {real, imag} */,
  {32'hc0a5f040, 32'h40b541cc} /* (4, 10, 13) {real, imag} */,
  {32'hbfdbb6b0, 32'h3f91d8d4} /* (4, 10, 12) {real, imag} */,
  {32'hc051d859, 32'hc0929818} /* (4, 10, 11) {real, imag} */,
  {32'hc0d717f6, 32'hc016c1d3} /* (4, 10, 10) {real, imag} */,
  {32'hc13016d1, 32'hc08440b0} /* (4, 10, 9) {real, imag} */,
  {32'hc0e76704, 32'hbff0436c} /* (4, 10, 8) {real, imag} */,
  {32'hc0f1a9c6, 32'hc1180973} /* (4, 10, 7) {real, imag} */,
  {32'hc1743182, 32'h40805fae} /* (4, 10, 6) {real, imag} */,
  {32'hc15a316d, 32'h417a7a1a} /* (4, 10, 5) {real, imag} */,
  {32'hc0e87cfa, 32'hc041b518} /* (4, 10, 4) {real, imag} */,
  {32'h40d300d6, 32'hc0a9cd3e} /* (4, 10, 3) {real, imag} */,
  {32'h40bbccc8, 32'h414fb552} /* (4, 10, 2) {real, imag} */,
  {32'h410b0ad8, 32'h40ddc6c1} /* (4, 10, 1) {real, imag} */,
  {32'h408031c4, 32'hbf17dd70} /* (4, 10, 0) {real, imag} */,
  {32'hc03d4ba1, 32'h3fbe64e2} /* (4, 9, 31) {real, imag} */,
  {32'hc1116785, 32'hc0b39a6f} /* (4, 9, 30) {real, imag} */,
  {32'hc08040ce, 32'h3d011540} /* (4, 9, 29) {real, imag} */,
  {32'h3f36d218, 32'h40512d8c} /* (4, 9, 28) {real, imag} */,
  {32'h40f43b7f, 32'h4072add8} /* (4, 9, 27) {real, imag} */,
  {32'h405a09f0, 32'hc0314694} /* (4, 9, 26) {real, imag} */,
  {32'hc1a1024b, 32'hc052d748} /* (4, 9, 25) {real, imag} */,
  {32'hc1980868, 32'h4118b960} /* (4, 9, 24) {real, imag} */,
  {32'hc0ad8cd5, 32'h41674c7e} /* (4, 9, 23) {real, imag} */,
  {32'h3fc1db0c, 32'hbe6fd8e0} /* (4, 9, 22) {real, imag} */,
  {32'h4093a3ed, 32'hc1574ba8} /* (4, 9, 21) {real, imag} */,
  {32'h4094dd88, 32'hbe2de280} /* (4, 9, 20) {real, imag} */,
  {32'h412410c3, 32'h4136b7cc} /* (4, 9, 19) {real, imag} */,
  {32'h41869aa8, 32'h418965fe} /* (4, 9, 18) {real, imag} */,
  {32'h4189d18e, 32'h4190d198} /* (4, 9, 17) {real, imag} */,
  {32'h40050fae, 32'h40880b5e} /* (4, 9, 16) {real, imag} */,
  {32'hc05f13fc, 32'hc128c906} /* (4, 9, 15) {real, imag} */,
  {32'hc096b50c, 32'hc12503bd} /* (4, 9, 14) {real, imag} */,
  {32'hbf4789ec, 32'hc0cc4fb7} /* (4, 9, 13) {real, imag} */,
  {32'h40bf3bd6, 32'hc11890e5} /* (4, 9, 12) {real, imag} */,
  {32'h3f22b284, 32'hbf159a2c} /* (4, 9, 11) {real, imag} */,
  {32'hc0c8c537, 32'hc09f65b9} /* (4, 9, 10) {real, imag} */,
  {32'hc18c03c6, 32'hc10f8d8f} /* (4, 9, 9) {real, imag} */,
  {32'hc15c4e27, 32'h407e5828} /* (4, 9, 8) {real, imag} */,
  {32'hc09a0a0f, 32'h3f832668} /* (4, 9, 7) {real, imag} */,
  {32'h40b2ea8e, 32'hc14e19e0} /* (4, 9, 6) {real, imag} */,
  {32'h3ffcc738, 32'hc1c64637} /* (4, 9, 5) {real, imag} */,
  {32'h40851082, 32'hc194317e} /* (4, 9, 4) {real, imag} */,
  {32'h3fe9da4a, 32'h3f49b834} /* (4, 9, 3) {real, imag} */,
  {32'hc0e5dee6, 32'hc10701af} /* (4, 9, 2) {real, imag} */,
  {32'hc18696e7, 32'hc0df3cd4} /* (4, 9, 1) {real, imag} */,
  {32'hbfc949ae, 32'h40235aab} /* (4, 9, 0) {real, imag} */,
  {32'h40d5b83b, 32'h4114914a} /* (4, 8, 31) {real, imag} */,
  {32'h3ff82ad0, 32'hbfceee04} /* (4, 8, 30) {real, imag} */,
  {32'hbf9b09b0, 32'hc12ae894} /* (4, 8, 29) {real, imag} */,
  {32'h41cbff14, 32'hc1860410} /* (4, 8, 28) {real, imag} */,
  {32'h41c21a2f, 32'hc1bb0eb4} /* (4, 8, 27) {real, imag} */,
  {32'h4180c5e6, 32'hc18f926b} /* (4, 8, 26) {real, imag} */,
  {32'h4194bc02, 32'hc1640030} /* (4, 8, 25) {real, imag} */,
  {32'h412797a2, 32'hc0868f16} /* (4, 8, 24) {real, imag} */,
  {32'h41497a26, 32'hc053323c} /* (4, 8, 23) {real, imag} */,
  {32'h41854dee, 32'hc0bbd9b5} /* (4, 8, 22) {real, imag} */,
  {32'hc088b4ba, 32'h4074cd10} /* (4, 8, 21) {real, imag} */,
  {32'hc201c9d2, 32'h4083cec6} /* (4, 8, 20) {real, imag} */,
  {32'hc1b8ebfb, 32'h40eea661} /* (4, 8, 19) {real, imag} */,
  {32'hc1a14628, 32'h4135025e} /* (4, 8, 18) {real, imag} */,
  {32'hc1a9b266, 32'h41278384} /* (4, 8, 17) {real, imag} */,
  {32'hc18afdae, 32'h40b03d2c} /* (4, 8, 16) {real, imag} */,
  {32'hc107cba4, 32'h41b39b0a} /* (4, 8, 15) {real, imag} */,
  {32'h408c7c28, 32'h414294fa} /* (4, 8, 14) {real, imag} */,
  {32'hc08b40f4, 32'h40d144e8} /* (4, 8, 13) {real, imag} */,
  {32'hc1ad904e, 32'h41966232} /* (4, 8, 12) {real, imag} */,
  {32'hc1f142c8, 32'h4177b9b3} /* (4, 8, 11) {real, imag} */,
  {32'hc1dde6b9, 32'h4122ffa2} /* (4, 8, 10) {real, imag} */,
  {32'h410d8100, 32'hbe65a4a0} /* (4, 8, 9) {real, imag} */,
  {32'h41c37670, 32'hc1a39693} /* (4, 8, 8) {real, imag} */,
  {32'h41aa609a, 32'hc1957bb0} /* (4, 8, 7) {real, imag} */,
  {32'h4088901b, 32'hc18cb965} /* (4, 8, 6) {real, imag} */,
  {32'hc0841ecf, 32'hc0bd4bd6} /* (4, 8, 5) {real, imag} */,
  {32'h41648c7e, 32'hc0bfac7d} /* (4, 8, 4) {real, imag} */,
  {32'h41223c94, 32'h40bd2a1c} /* (4, 8, 3) {real, imag} */,
  {32'h41122751, 32'hc0c8fd21} /* (4, 8, 2) {real, imag} */,
  {32'h41c64cb2, 32'hc099794c} /* (4, 8, 1) {real, imag} */,
  {32'h4193aaee, 32'h40a1e334} /* (4, 8, 0) {real, imag} */,
  {32'hc07f4864, 32'h40d62e5c} /* (4, 7, 31) {real, imag} */,
  {32'h3ffd8628, 32'h40cc18ab} /* (4, 7, 30) {real, imag} */,
  {32'hc0a8cdbe, 32'h41599c9f} /* (4, 7, 29) {real, imag} */,
  {32'hc17ae413, 32'h415580ac} /* (4, 7, 28) {real, imag} */,
  {32'hc1765a4c, 32'hc00ec34a} /* (4, 7, 27) {real, imag} */,
  {32'hc151465e, 32'h4008225c} /* (4, 7, 26) {real, imag} */,
  {32'h406b6dca, 32'h41b38270} /* (4, 7, 25) {real, imag} */,
  {32'h413ca87d, 32'h419922a9} /* (4, 7, 24) {real, imag} */,
  {32'hc171704e, 32'h414f2452} /* (4, 7, 23) {real, imag} */,
  {32'hc1a61268, 32'h4070fc3e} /* (4, 7, 22) {real, imag} */,
  {32'hc20127ef, 32'h41bf650c} /* (4, 7, 21) {real, imag} */,
  {32'hc1cb42b1, 32'h4122491f} /* (4, 7, 20) {real, imag} */,
  {32'h40ba2b2b, 32'h40ff9701} /* (4, 7, 19) {real, imag} */,
  {32'h41d75aaa, 32'hc082ab0e} /* (4, 7, 18) {real, imag} */,
  {32'h414776e0, 32'hc16c1ae3} /* (4, 7, 17) {real, imag} */,
  {32'h402c1d52, 32'h40fbb772} /* (4, 7, 16) {real, imag} */,
  {32'h416b6bea, 32'h3fb93f50} /* (4, 7, 15) {real, imag} */,
  {32'h419c3e46, 32'hc126c6cb} /* (4, 7, 14) {real, imag} */,
  {32'h3e30be80, 32'hc15d6672} /* (4, 7, 13) {real, imag} */,
  {32'h413dc062, 32'hc1366898} /* (4, 7, 12) {real, imag} */,
  {32'h4154fec6, 32'hc0ccbf92} /* (4, 7, 11) {real, imag} */,
  {32'hbf6cc7e0, 32'h40ae506c} /* (4, 7, 10) {real, imag} */,
  {32'hbeaa16e0, 32'hc1051db2} /* (4, 7, 9) {real, imag} */,
  {32'hc0ca87e2, 32'hc140ed68} /* (4, 7, 8) {real, imag} */,
  {32'hc18ccf87, 32'h400d1688} /* (4, 7, 7) {real, imag} */,
  {32'hc18060e0, 32'h4111f790} /* (4, 7, 6) {real, imag} */,
  {32'hc0a961ec, 32'h40299b48} /* (4, 7, 5) {real, imag} */,
  {32'h4165b1c7, 32'hc084c590} /* (4, 7, 4) {real, imag} */,
  {32'h40fde46a, 32'h4051348b} /* (4, 7, 3) {real, imag} */,
  {32'hc0a41f62, 32'h3ed2ced0} /* (4, 7, 2) {real, imag} */,
  {32'hc1959f9c, 32'h4085581c} /* (4, 7, 1) {real, imag} */,
  {32'hc0e15131, 32'h3eddb5f8} /* (4, 7, 0) {real, imag} */,
  {32'hc1772363, 32'hc0b40aca} /* (4, 6, 31) {real, imag} */,
  {32'hc1ffee04, 32'hc1a2f687} /* (4, 6, 30) {real, imag} */,
  {32'hc0d9bbf8, 32'hc193ad97} /* (4, 6, 29) {real, imag} */,
  {32'h410ae618, 32'hc04e4980} /* (4, 6, 28) {real, imag} */,
  {32'hc17f6f6f, 32'hc0735e8f} /* (4, 6, 27) {real, imag} */,
  {32'hc18b79ab, 32'hc08c5928} /* (4, 6, 26) {real, imag} */,
  {32'hbe469f40, 32'hc0d2bbfc} /* (4, 6, 25) {real, imag} */,
  {32'h412f47d5, 32'hc0de4f24} /* (4, 6, 24) {real, imag} */,
  {32'h40b1610f, 32'h40283d38} /* (4, 6, 23) {real, imag} */,
  {32'hbf587740, 32'hc1138a6d} /* (4, 6, 22) {real, imag} */,
  {32'h4091d641, 32'hc11c14c4} /* (4, 6, 21) {real, imag} */,
  {32'h4012f9b9, 32'hbe37c5c0} /* (4, 6, 20) {real, imag} */,
  {32'h41161529, 32'h402d5a00} /* (4, 6, 19) {real, imag} */,
  {32'h419258a9, 32'hc036a79a} /* (4, 6, 18) {real, imag} */,
  {32'hc084b977, 32'hbfcf8d92} /* (4, 6, 17) {real, imag} */,
  {32'hc119bfd7, 32'hbf9d41cc} /* (4, 6, 16) {real, imag} */,
  {32'hbea41ea0, 32'hc07ad554} /* (4, 6, 15) {real, imag} */,
  {32'hc1b8b57c, 32'h3fc0fe88} /* (4, 6, 14) {real, imag} */,
  {32'hc18d9952, 32'hc04e4dd8} /* (4, 6, 13) {real, imag} */,
  {32'h406cfc5c, 32'hc10e0019} /* (4, 6, 12) {real, imag} */,
  {32'h41023948, 32'hbfd54cd0} /* (4, 6, 11) {real, imag} */,
  {32'h4083fef6, 32'hc0cb67e7} /* (4, 6, 10) {real, imag} */,
  {32'hbf8420be, 32'h400e1814} /* (4, 6, 9) {real, imag} */,
  {32'h4161dec2, 32'h4117ea48} /* (4, 6, 8) {real, imag} */,
  {32'h4180d5a9, 32'h4066c2f8} /* (4, 6, 7) {real, imag} */,
  {32'h40b7bd60, 32'hc0ec20bc} /* (4, 6, 6) {real, imag} */,
  {32'h407133e8, 32'hc11c18e7} /* (4, 6, 5) {real, imag} */,
  {32'h3f784ac8, 32'hc0207036} /* (4, 6, 4) {real, imag} */,
  {32'hc06c7c24, 32'hc10286a9} /* (4, 6, 3) {real, imag} */,
  {32'h3fd10b68, 32'h4160af7d} /* (4, 6, 2) {real, imag} */,
  {32'hc171a45a, 32'h3e86f200} /* (4, 6, 1) {real, imag} */,
  {32'hc1282a0c, 32'hc142f25f} /* (4, 6, 0) {real, imag} */,
  {32'h4168f843, 32'h3fd065c8} /* (4, 5, 31) {real, imag} */,
  {32'h41eef078, 32'h3f5addb0} /* (4, 5, 30) {real, imag} */,
  {32'h415c993e, 32'hc114d9b0} /* (4, 5, 29) {real, imag} */,
  {32'h4022ea11, 32'hc16b82b8} /* (4, 5, 28) {real, imag} */,
  {32'h41795831, 32'hc146f4dc} /* (4, 5, 27) {real, imag} */,
  {32'h418ce592, 32'hc17d3acc} /* (4, 5, 26) {real, imag} */,
  {32'h416db7e7, 32'hc1c48166} /* (4, 5, 25) {real, imag} */,
  {32'h410b4015, 32'hc1b7b686} /* (4, 5, 24) {real, imag} */,
  {32'h3f09eebc, 32'hc1cd1282} /* (4, 5, 23) {real, imag} */,
  {32'h40ad4f6b, 32'hc18a312b} /* (4, 5, 22) {real, imag} */,
  {32'h40eb16f0, 32'h4125215e} /* (4, 5, 21) {real, imag} */,
  {32'h40a91ca2, 32'h41478f9e} /* (4, 5, 20) {real, imag} */,
  {32'hc14be6d6, 32'hc11f36de} /* (4, 5, 19) {real, imag} */,
  {32'hc193dc79, 32'hc0be8e1f} /* (4, 5, 18) {real, imag} */,
  {32'hc121510e, 32'h40e9242b} /* (4, 5, 17) {real, imag} */,
  {32'hc048add9, 32'h40c9d86c} /* (4, 5, 16) {real, imag} */,
  {32'hbece8ce0, 32'h418aacd8} /* (4, 5, 15) {real, imag} */,
  {32'hbf1dc3f8, 32'h41bc55f0} /* (4, 5, 14) {real, imag} */,
  {32'hc0279683, 32'h407fe220} /* (4, 5, 13) {real, imag} */,
  {32'hc13b44dc, 32'h40975b60} /* (4, 5, 12) {real, imag} */,
  {32'hc1a5c3b1, 32'h41437cdb} /* (4, 5, 11) {real, imag} */,
  {32'h4113694c, 32'h400400ee} /* (4, 5, 10) {real, imag} */,
  {32'h410c377d, 32'hc05da805} /* (4, 5, 9) {real, imag} */,
  {32'h4185b683, 32'hc17a87fb} /* (4, 5, 8) {real, imag} */,
  {32'h4196da05, 32'h40d6f989} /* (4, 5, 7) {real, imag} */,
  {32'hc0c609c2, 32'h419edf04} /* (4, 5, 6) {real, imag} */,
  {32'h411bee61, 32'h402a3578} /* (4, 5, 5) {real, imag} */,
  {32'h415f60b0, 32'hc1d96fb9} /* (4, 5, 4) {real, imag} */,
  {32'h4135999a, 32'hc2029c3f} /* (4, 5, 3) {real, imag} */,
  {32'h4116f89c, 32'hc138dfa7} /* (4, 5, 2) {real, imag} */,
  {32'hbefb5a70, 32'hc1021623} /* (4, 5, 1) {real, imag} */,
  {32'h4118f3da, 32'hc136652b} /* (4, 5, 0) {real, imag} */,
  {32'hc1a859b0, 32'h411a1be3} /* (4, 4, 31) {real, imag} */,
  {32'hc1656d0c, 32'h41a9b4b4} /* (4, 4, 30) {real, imag} */,
  {32'hbeadc540, 32'h417b5438} /* (4, 4, 29) {real, imag} */,
  {32'h4108ca38, 32'h418cd841} /* (4, 4, 28) {real, imag} */,
  {32'hc08434ee, 32'h414964c7} /* (4, 4, 27) {real, imag} */,
  {32'hc178035e, 32'h41129d76} /* (4, 4, 26) {real, imag} */,
  {32'hc1b131bc, 32'h417c02da} /* (4, 4, 25) {real, imag} */,
  {32'hc2088d42, 32'h40e43580} /* (4, 4, 24) {real, imag} */,
  {32'hc1e9ecf7, 32'h3fae7420} /* (4, 4, 23) {real, imag} */,
  {32'hc134c712, 32'hc0a06aa6} /* (4, 4, 22) {real, imag} */,
  {32'h419d61f6, 32'hc17e3242} /* (4, 4, 21) {real, imag} */,
  {32'h42167f26, 32'hc18b1594} /* (4, 4, 20) {real, imag} */,
  {32'h41dd7a48, 32'hc1c4ab3e} /* (4, 4, 19) {real, imag} */,
  {32'h42373c59, 32'hc1183573} /* (4, 4, 18) {real, imag} */,
  {32'h427020ea, 32'hc0ce8232} /* (4, 4, 17) {real, imag} */,
  {32'h41dc7882, 32'hc1883bbc} /* (4, 4, 16) {real, imag} */,
  {32'h4099e607, 32'hc19a5d75} /* (4, 4, 15) {real, imag} */,
  {32'h406cda5b, 32'hc1df8cbc} /* (4, 4, 14) {real, imag} */,
  {32'hc05c9a60, 32'hc1af9235} /* (4, 4, 13) {real, imag} */,
  {32'h413dbe0c, 32'hc1e74101} /* (4, 4, 12) {real, imag} */,
  {32'h417590fd, 32'hc15d9635} /* (4, 4, 11) {real, imag} */,
  {32'hc150e68c, 32'h411c49ed} /* (4, 4, 10) {real, imag} */,
  {32'hc24d6afc, 32'h40978522} /* (4, 4, 9) {real, imag} */,
  {32'hc22d990e, 32'h4101204b} /* (4, 4, 8) {real, imag} */,
  {32'hc1c6291a, 32'h40463454} /* (4, 4, 7) {real, imag} */,
  {32'hc19e1408, 32'hc04380d8} /* (4, 4, 6) {real, imag} */,
  {32'hc1b6d097, 32'h4170b49b} /* (4, 4, 5) {real, imag} */,
  {32'hc1827992, 32'h41500a07} /* (4, 4, 4) {real, imag} */,
  {32'h3fd3f624, 32'h41eb5896} /* (4, 4, 3) {real, imag} */,
  {32'hc18079c9, 32'h41e08424} /* (4, 4, 2) {real, imag} */,
  {32'hc1b3edce, 32'h420cc0f6} /* (4, 4, 1) {real, imag} */,
  {32'hc156162b, 32'h41bdd97d} /* (4, 4, 0) {real, imag} */,
  {32'h4141a3a4, 32'h408d6788} /* (4, 3, 31) {real, imag} */,
  {32'h4126198e, 32'h3e4cae90} /* (4, 3, 30) {real, imag} */,
  {32'hc12091a6, 32'hc1147fd3} /* (4, 3, 29) {real, imag} */,
  {32'hc1b59618, 32'hc0ceb472} /* (4, 3, 28) {real, imag} */,
  {32'hc04b663c, 32'h418793d4} /* (4, 3, 27) {real, imag} */,
  {32'h41251231, 32'h4147264a} /* (4, 3, 26) {real, imag} */,
  {32'h411e19ad, 32'hc02796e6} /* (4, 3, 25) {real, imag} */,
  {32'hc1896ce4, 32'hc1710de0} /* (4, 3, 24) {real, imag} */,
  {32'h3f5f1ec0, 32'hc12ed725} /* (4, 3, 23) {real, imag} */,
  {32'h40465672, 32'h41986db0} /* (4, 3, 22) {real, imag} */,
  {32'h414bb40d, 32'h40259ac4} /* (4, 3, 21) {real, imag} */,
  {32'h4200b621, 32'h4192d86a} /* (4, 3, 20) {real, imag} */,
  {32'h41621f8a, 32'h41e3d77c} /* (4, 3, 19) {real, imag} */,
  {32'h40f38e60, 32'h41d89d1c} /* (4, 3, 18) {real, imag} */,
  {32'h4208c027, 32'h4174c895} /* (4, 3, 17) {real, imag} */,
  {32'h41c89bd4, 32'h412e843c} /* (4, 3, 16) {real, imag} */,
  {32'h41346621, 32'hc1254bab} /* (4, 3, 15) {real, imag} */,
  {32'h41ca4636, 32'h40a209c5} /* (4, 3, 14) {real, imag} */,
  {32'h3fcd7a38, 32'h3fa4fa88} /* (4, 3, 13) {real, imag} */,
  {32'hbff4cb10, 32'h41a94694} /* (4, 3, 12) {real, imag} */,
  {32'hc18b8366, 32'h40c8aabc} /* (4, 3, 11) {real, imag} */,
  {32'hc212bc8c, 32'hc182fb98} /* (4, 3, 10) {real, imag} */,
  {32'hc1d5b09c, 32'hc0880d5c} /* (4, 3, 9) {real, imag} */,
  {32'hc137332b, 32'hc0cb8fbe} /* (4, 3, 8) {real, imag} */,
  {32'hc1b7f230, 32'hc179fce0} /* (4, 3, 7) {real, imag} */,
  {32'hc1916d00, 32'hc1e9740f} /* (4, 3, 6) {real, imag} */,
  {32'hc085a8f4, 32'hc187cd89} /* (4, 3, 5) {real, imag} */,
  {32'h41211723, 32'hc14932c9} /* (4, 3, 4) {real, imag} */,
  {32'h3fc27780, 32'hc2035cf5} /* (4, 3, 3) {real, imag} */,
  {32'hc04faa20, 32'hc199e17d} /* (4, 3, 2) {real, imag} */,
  {32'h4093bfb6, 32'hc0dc714c} /* (4, 3, 1) {real, imag} */,
  {32'hbf94c9f8, 32'h40df29cc} /* (4, 3, 0) {real, imag} */,
  {32'h41b992dc, 32'hc20393e2} /* (4, 2, 31) {real, imag} */,
  {32'h42107b62, 32'hc25122fb} /* (4, 2, 30) {real, imag} */,
  {32'h4206b0cb, 32'hc22f984c} /* (4, 2, 29) {real, imag} */,
  {32'h41acfbf3, 32'hc1f7af7b} /* (4, 2, 28) {real, imag} */,
  {32'h41fd9432, 32'hc23c467a} /* (4, 2, 27) {real, imag} */,
  {32'h4164c19e, 32'hc27595d2} /* (4, 2, 26) {real, imag} */,
  {32'h41868a22, 32'hc2392a20} /* (4, 2, 25) {real, imag} */,
  {32'h41eeb878, 32'hc2265370} /* (4, 2, 24) {real, imag} */,
  {32'h4204d78c, 32'hc23314be} /* (4, 2, 23) {real, imag} */,
  {32'h41f77eb5, 32'hc26e8c8e} /* (4, 2, 22) {real, imag} */,
  {32'h41cfc7f9, 32'hc120bcaa} /* (4, 2, 21) {real, imag} */,
  {32'h41b71f80, 32'h429c0db8} /* (4, 2, 20) {real, imag} */,
  {32'h4076e970, 32'h4294b741} /* (4, 2, 19) {real, imag} */,
  {32'h40bfa508, 32'h42923f16} /* (4, 2, 18) {real, imag} */,
  {32'hc1324be6, 32'h42a5c168} /* (4, 2, 17) {real, imag} */,
  {32'hc20c88aa, 32'h428a7578} /* (4, 2, 16) {real, imag} */,
  {32'hc1b5ea7e, 32'h423bd4d8} /* (4, 2, 15) {real, imag} */,
  {32'hc189dda8, 32'h42660e3d} /* (4, 2, 14) {real, imag} */,
  {32'hc15dff4d, 32'h42280ea4} /* (4, 2, 13) {real, imag} */,
  {32'hc1c67ca1, 32'h4207d746} /* (4, 2, 12) {real, imag} */,
  {32'hc1893427, 32'h3fbde688} /* (4, 2, 11) {real, imag} */,
  {32'hc131373a, 32'hc28bf1f7} /* (4, 2, 10) {real, imag} */,
  {32'h40b65478, 32'hc2c06e81} /* (4, 2, 9) {real, imag} */,
  {32'h408c5da4, 32'hc2a44507} /* (4, 2, 8) {real, imag} */,
  {32'h3e9b4e00, 32'hc28a2dd6} /* (4, 2, 7) {real, imag} */,
  {32'h40322934, 32'hc27910b9} /* (4, 2, 6) {real, imag} */,
  {32'h4190a22e, 32'hc25250ef} /* (4, 2, 5) {real, imag} */,
  {32'h41e964e8, 32'hc1ecdda8} /* (4, 2, 4) {real, imag} */,
  {32'h41c2fcac, 32'hc225729c} /* (4, 2, 3) {real, imag} */,
  {32'h418d4428, 32'hc25f6685} /* (4, 2, 2) {real, imag} */,
  {32'h41cadad7, 32'hc26a6761} /* (4, 2, 1) {real, imag} */,
  {32'h410e3698, 32'hc2034062} /* (4, 2, 0) {real, imag} */,
  {32'hc120003b, 32'h4203b8f7} /* (4, 1, 31) {real, imag} */,
  {32'hc23704da, 32'h427e6b74} /* (4, 1, 30) {real, imag} */,
  {32'hc282e3ac, 32'h4284d6a9} /* (4, 1, 29) {real, imag} */,
  {32'hc237e123, 32'h428d26d8} /* (4, 1, 28) {real, imag} */,
  {32'hc2131964, 32'h42810d89} /* (4, 1, 27) {real, imag} */,
  {32'hc218de84, 32'h426a8a88} /* (4, 1, 26) {real, imag} */,
  {32'hc20cfaab, 32'h42817cd1} /* (4, 1, 25) {real, imag} */,
  {32'hc1dc55c8, 32'h42885db2} /* (4, 1, 24) {real, imag} */,
  {32'hc25c742b, 32'h42987b26} /* (4, 1, 23) {real, imag} */,
  {32'hc24a00ce, 32'h42c1e51c} /* (4, 1, 22) {real, imag} */,
  {32'hc24d0b16, 32'h42954ce0} /* (4, 1, 21) {real, imag} */,
  {32'h3fc4f588, 32'hc1b54f73} /* (4, 1, 20) {real, imag} */,
  {32'h421b62bc, 32'hc209252e} /* (4, 1, 19) {real, imag} */,
  {32'h42222bad, 32'h40b0fd3c} /* (4, 1, 18) {real, imag} */,
  {32'h421ad2be, 32'hc15db410} /* (4, 1, 17) {real, imag} */,
  {32'h422910ff, 32'hc1a472cb} /* (4, 1, 16) {real, imag} */,
  {32'h41a6226f, 32'hc25d629f} /* (4, 1, 15) {real, imag} */,
  {32'h42461404, 32'hc2aea7cc} /* (4, 1, 14) {real, imag} */,
  {32'h42363bcb, 32'hc2a48ca8} /* (4, 1, 13) {real, imag} */,
  {32'h419e4b99, 32'hc28dc1f1} /* (4, 1, 12) {real, imag} */,
  {32'h41af5bac, 32'hc28d9ad9} /* (4, 1, 11) {real, imag} */,
  {32'hc1cc223a, 32'h3ed88360} /* (4, 1, 10) {real, imag} */,
  {32'hc29dcfa4, 32'h411d49d2} /* (4, 1, 9) {real, imag} */,
  {32'hc27487ff, 32'h40f6d478} /* (4, 1, 8) {real, imag} */,
  {32'hc2851dd1, 32'h41f7ffc2} /* (4, 1, 7) {real, imag} */,
  {32'hc2667d0c, 32'h41ddd458} /* (4, 1, 6) {real, imag} */,
  {32'hc23efa63, 32'h423d8831} /* (4, 1, 5) {real, imag} */,
  {32'hc20a69a4, 32'h4280de3c} /* (4, 1, 4) {real, imag} */,
  {32'hc2061257, 32'h42715523} /* (4, 1, 3) {real, imag} */,
  {32'hc2153b50, 32'h4289903c} /* (4, 1, 2) {real, imag} */,
  {32'hc179a4e7, 32'h4297ac21} /* (4, 1, 1) {real, imag} */,
  {32'hc111d775, 32'h421c27d4} /* (4, 1, 0) {real, imag} */,
  {32'hc181d893, 32'h424731af} /* (4, 0, 31) {real, imag} */,
  {32'hc21670eb, 32'h429205ae} /* (4, 0, 30) {real, imag} */,
  {32'hc20ca236, 32'h42341168} /* (4, 0, 29) {real, imag} */,
  {32'hc1bffea8, 32'h423001bb} /* (4, 0, 28) {real, imag} */,
  {32'hc2066d12, 32'h4210303c} /* (4, 0, 27) {real, imag} */,
  {32'hc1ee0634, 32'h42714826} /* (4, 0, 26) {real, imag} */,
  {32'hc1caae00, 32'h424711c8} /* (4, 0, 25) {real, imag} */,
  {32'hc03aa95f, 32'h4225dc5a} /* (4, 0, 24) {real, imag} */,
  {32'hc035bc3e, 32'h422118d5} /* (4, 0, 23) {real, imag} */,
  {32'hc190369f, 32'h425dfbb9} /* (4, 0, 22) {real, imag} */,
  {32'hc189583c, 32'h4213c061} /* (4, 0, 21) {real, imag} */,
  {32'h40ec5eae, 32'hc11f63a0} /* (4, 0, 20) {real, imag} */,
  {32'hc192b0ba, 32'h413c1606} /* (4, 0, 19) {real, imag} */,
  {32'hc1a49a5a, 32'h4177aa72} /* (4, 0, 18) {real, imag} */,
  {32'hc08a4a61, 32'hbe5dfda0} /* (4, 0, 17) {real, imag} */,
  {32'h3f8a2d04, 32'hc14dd744} /* (4, 0, 16) {real, imag} */,
  {32'h40880725, 32'hc202d910} /* (4, 0, 15) {real, imag} */,
  {32'h41c57e97, 32'hc24ff9c0} /* (4, 0, 14) {real, imag} */,
  {32'h4202f5be, 32'hc245839a} /* (4, 0, 13) {real, imag} */,
  {32'h416cf63f, 32'hc2260779} /* (4, 0, 12) {real, imag} */,
  {32'h41707bef, 32'hc23f4df2} /* (4, 0, 11) {real, imag} */,
  {32'h40db79d8, 32'hc207bef9} /* (4, 0, 10) {real, imag} */,
  {32'hc191f85b, 32'hc0e96646} /* (4, 0, 9) {real, imag} */,
  {32'hc153b788, 32'hc00d5a54} /* (4, 0, 8) {real, imag} */,
  {32'hc0020614, 32'hc1b12cf1} /* (4, 0, 7) {real, imag} */,
  {32'h4176f814, 32'hc1aa7275} /* (4, 0, 6) {real, imag} */,
  {32'hc12c53a4, 32'h42309369} /* (4, 0, 5) {real, imag} */,
  {32'hc1bdf2f8, 32'h4271ecd9} /* (4, 0, 4) {real, imag} */,
  {32'hc11ce23a, 32'h425132f6} /* (4, 0, 3) {real, imag} */,
  {32'hc1ac4342, 32'h42486bb0} /* (4, 0, 2) {real, imag} */,
  {32'hc19066ab, 32'h42501f03} /* (4, 0, 1) {real, imag} */,
  {32'hc0cb50cc, 32'h4198b57a} /* (4, 0, 0) {real, imag} */,
  {32'hc197be20, 32'h42440d83} /* (3, 31, 31) {real, imag} */,
  {32'hc17ed0d0, 32'h42956e72} /* (3, 31, 30) {real, imag} */,
  {32'hc183c77b, 32'h42b349ca} /* (3, 31, 29) {real, imag} */,
  {32'hc1d78f84, 32'h42e616f8} /* (3, 31, 28) {real, imag} */,
  {32'hc1b4ae41, 32'h42d10e61} /* (3, 31, 27) {real, imag} */,
  {32'hc16c0812, 32'h42af6ce7} /* (3, 31, 26) {real, imag} */,
  {32'hc1f12eb0, 32'h42af8c94} /* (3, 31, 25) {real, imag} */,
  {32'hc1d142dc, 32'h42b9acb9} /* (3, 31, 24) {real, imag} */,
  {32'hc20f53ec, 32'h429ce9a1} /* (3, 31, 23) {real, imag} */,
  {32'hc203ebc4, 32'h428df5b4} /* (3, 31, 22) {real, imag} */,
  {32'hc12fedc0, 32'h4243d83f} /* (3, 31, 21) {real, imag} */,
  {32'hc1e888ac, 32'hc1e7c688} /* (3, 31, 20) {real, imag} */,
  {32'hc1dbb601, 32'hc1bc5d6c} /* (3, 31, 19) {real, imag} */,
  {32'hc10e1dd8, 32'hc2015a68} /* (3, 31, 18) {real, imag} */,
  {32'h3ef645c0, 32'hc1ee1381} /* (3, 31, 17) {real, imag} */,
  {32'hc167631f, 32'hc2616478} /* (3, 31, 16) {real, imag} */,
  {32'hc11380aa, 32'hc28655b0} /* (3, 31, 15) {real, imag} */,
  {32'h40af4d18, 32'hc29938f1} /* (3, 31, 14) {real, imag} */,
  {32'h41e6038b, 32'hc2bfaaf7} /* (3, 31, 13) {real, imag} */,
  {32'h4210f1a7, 32'hc2eea4d1} /* (3, 31, 12) {real, imag} */,
  {32'h42085c0b, 32'hc2b923f0} /* (3, 31, 11) {real, imag} */,
  {32'h4265e188, 32'h41ded9f5} /* (3, 31, 10) {real, imag} */,
  {32'h424a2b61, 32'h42894ff9} /* (3, 31, 9) {real, imag} */,
  {32'h41bfd9fa, 32'h429e65b5} /* (3, 31, 8) {real, imag} */,
  {32'h41db475c, 32'h429017a0} /* (3, 31, 7) {real, imag} */,
  {32'h41bf19b6, 32'h42147f58} /* (3, 31, 6) {real, imag} */,
  {32'hc05b9140, 32'h42794f7c} /* (3, 31, 5) {real, imag} */,
  {32'hc06b3664, 32'h429efe36} /* (3, 31, 4) {real, imag} */,
  {32'hc154132a, 32'h429c94ce} /* (3, 31, 3) {real, imag} */,
  {32'hc1dca6de, 32'h42877dd2} /* (3, 31, 2) {real, imag} */,
  {32'hc1e332c4, 32'h429b3c63} /* (3, 31, 1) {real, imag} */,
  {32'hc0e11131, 32'h42261035} /* (3, 31, 0) {real, imag} */,
  {32'h40cf94b9, 32'hc2598893} /* (3, 30, 31) {real, imag} */,
  {32'h417c571c, 32'hc2b8785c} /* (3, 30, 30) {real, imag} */,
  {32'h3ed2d440, 32'hc270c099} /* (3, 30, 29) {real, imag} */,
  {32'hc20893a9, 32'hc2083461} /* (3, 30, 28) {real, imag} */,
  {32'hc180b9a0, 32'hc243418e} /* (3, 30, 27) {real, imag} */,
  {32'h3ebd2540, 32'hc289bb29} /* (3, 30, 26) {real, imag} */,
  {32'h4014dff0, 32'hc281431b} /* (3, 30, 25) {real, imag} */,
  {32'h40a72d2c, 32'hc280eaa4} /* (3, 30, 24) {real, imag} */,
  {32'h41a386ac, 32'hc28ffd6d} /* (3, 30, 23) {real, imag} */,
  {32'h421f5016, 32'hc24b3eec} /* (3, 30, 22) {real, imag} */,
  {32'h4185b532, 32'h416351e6} /* (3, 30, 21) {real, imag} */,
  {32'hc2311cec, 32'h426c961b} /* (3, 30, 20) {real, imag} */,
  {32'hc279306f, 32'h42264a3f} /* (3, 30, 19) {real, imag} */,
  {32'hc23dd895, 32'h4248b30c} /* (3, 30, 18) {real, imag} */,
  {32'hc25236b2, 32'h4284c3ed} /* (3, 30, 17) {real, imag} */,
  {32'hc21bce61, 32'h423d5dae} /* (3, 30, 16) {real, imag} */,
  {32'hc16fb76d, 32'h4259ea3a} /* (3, 30, 15) {real, imag} */,
  {32'hc1a5b50a, 32'h425cdc45} /* (3, 30, 14) {real, imag} */,
  {32'hc1b8e254, 32'h42637b72} /* (3, 30, 13) {real, imag} */,
  {32'hc10a9ddd, 32'h4242eabe} /* (3, 30, 12) {real, imag} */,
  {32'h408e314a, 32'h41d84077} /* (3, 30, 11) {real, imag} */,
  {32'h419f37a4, 32'hc20913b6} /* (3, 30, 10) {real, imag} */,
  {32'h4211f7ba, 32'hc28b4265} /* (3, 30, 9) {real, imag} */,
  {32'h4242aaee, 32'hc2999cdf} /* (3, 30, 8) {real, imag} */,
  {32'h4247943b, 32'hc2a68160} /* (3, 30, 7) {real, imag} */,
  {32'h423d0788, 32'hc28f344b} /* (3, 30, 6) {real, imag} */,
  {32'h415a889a, 32'hc2890675} /* (3, 30, 5) {real, imag} */,
  {32'h41a376b0, 32'hc272ec84} /* (3, 30, 4) {real, imag} */,
  {32'h4133f512, 32'hc29887de} /* (3, 30, 3) {real, imag} */,
  {32'hbe000f80, 32'hc278e085} /* (3, 30, 2) {real, imag} */,
  {32'hc19453d0, 32'hc23b7123} /* (3, 30, 1) {real, imag} */,
  {32'hc1d444be, 32'hc1e4a59a} /* (3, 30, 0) {real, imag} */,
  {32'hc14a5846, 32'h40ab71fc} /* (3, 29, 31) {real, imag} */,
  {32'hc1ff7696, 32'h41073668} /* (3, 29, 30) {real, imag} */,
  {32'hc180b228, 32'hc0925cfa} /* (3, 29, 29) {real, imag} */,
  {32'h3e540ba0, 32'hc0983262} /* (3, 29, 28) {real, imag} */,
  {32'hc068fe14, 32'hc20237fb} /* (3, 29, 27) {real, imag} */,
  {32'hc0f87d60, 32'hc200e84a} /* (3, 29, 26) {real, imag} */,
  {32'hc18b0eee, 32'hc0bf7066} /* (3, 29, 25) {real, imag} */,
  {32'h409cc251, 32'hc19d7fc8} /* (3, 29, 24) {real, imag} */,
  {32'h41461878, 32'hbff67940} /* (3, 29, 23) {real, imag} */,
  {32'h414d60cd, 32'h4125ca9f} /* (3, 29, 22) {real, imag} */,
  {32'hc05771ae, 32'h416fc0dc} /* (3, 29, 21) {real, imag} */,
  {32'hc230eb58, 32'hc1e7a094} /* (3, 29, 20) {real, imag} */,
  {32'hc2543c1b, 32'hc0bead74} /* (3, 29, 19) {real, imag} */,
  {32'hc1f9ff96, 32'h419cb30e} /* (3, 29, 18) {real, imag} */,
  {32'hc233e51a, 32'hc07f1e2a} /* (3, 29, 17) {real, imag} */,
  {32'hc2129be2, 32'hc0f280a6} /* (3, 29, 16) {real, imag} */,
  {32'h3ff61b84, 32'h41847742} /* (3, 29, 15) {real, imag} */,
  {32'h413835d4, 32'h3fc0f048} /* (3, 29, 14) {real, imag} */,
  {32'hc13df4f8, 32'hc0e302da} /* (3, 29, 13) {real, imag} */,
  {32'hc1393b08, 32'hc0d9a27a} /* (3, 29, 12) {real, imag} */,
  {32'h4105b10a, 32'hc07be7e8} /* (3, 29, 11) {real, imag} */,
  {32'h424bc962, 32'h4137bc48} /* (3, 29, 10) {real, imag} */,
  {32'h4277450a, 32'hbf741f40} /* (3, 29, 9) {real, imag} */,
  {32'h42502fdb, 32'hc054aba4} /* (3, 29, 8) {real, imag} */,
  {32'h41d0f253, 32'h408b4c4c} /* (3, 29, 7) {real, imag} */,
  {32'h41b818c1, 32'h40350fcc} /* (3, 29, 6) {real, imag} */,
  {32'h41d14ca2, 32'hbfd0ecc8} /* (3, 29, 5) {real, imag} */,
  {32'h4147cea4, 32'hc00e751e} /* (3, 29, 4) {real, imag} */,
  {32'h40ed6a9e, 32'h403e6d40} /* (3, 29, 3) {real, imag} */,
  {32'h3ec18400, 32'h4128d44f} /* (3, 29, 2) {real, imag} */,
  {32'hc19077fa, 32'h3f52cff0} /* (3, 29, 1) {real, imag} */,
  {32'hc1554892, 32'hc10e34f6} /* (3, 29, 0) {real, imag} */,
  {32'h411ae2b2, 32'h407e10fb} /* (3, 28, 31) {real, imag} */,
  {32'h3eaf5e8a, 32'hc03cd2a6} /* (3, 28, 30) {real, imag} */,
  {32'hc0e71aa5, 32'h415b9198} /* (3, 28, 29) {real, imag} */,
  {32'h41cbf048, 32'h419b7e34} /* (3, 28, 28) {real, imag} */,
  {32'h411ee156, 32'h4205d80e} /* (3, 28, 27) {real, imag} */,
  {32'hc0abda08, 32'h41b4f616} /* (3, 28, 26) {real, imag} */,
  {32'h4129dc1e, 32'h4206a81f} /* (3, 28, 25) {real, imag} */,
  {32'h40f2139c, 32'h41ee0ada} /* (3, 28, 24) {real, imag} */,
  {32'hc10ff599, 32'h41b4f345} /* (3, 28, 23) {real, imag} */,
  {32'h3f8ceb20, 32'h41686946} /* (3, 28, 22) {real, imag} */,
  {32'h40a1e0b8, 32'hc1941e62} /* (3, 28, 21) {real, imag} */,
  {32'hc1d4904f, 32'hc1f454c6} /* (3, 28, 20) {real, imag} */,
  {32'hc1cba013, 32'hc1b4ef57} /* (3, 28, 19) {real, imag} */,
  {32'hc130e852, 32'hc1af5964} /* (3, 28, 18) {real, imag} */,
  {32'hc18fb6d8, 32'hc208bfc2} /* (3, 28, 17) {real, imag} */,
  {32'hc16f4089, 32'hc2363834} /* (3, 28, 16) {real, imag} */,
  {32'hc1146aa6, 32'hc1cade76} /* (3, 28, 15) {real, imag} */,
  {32'hc18ae704, 32'hc1fa83ee} /* (3, 28, 14) {real, imag} */,
  {32'hc10c9890, 32'hc18db66b} /* (3, 28, 13) {real, imag} */,
  {32'hc024ab24, 32'hc1308f50} /* (3, 28, 12) {real, imag} */,
  {32'h4080e7ff, 32'h4003ce26} /* (3, 28, 11) {real, imag} */,
  {32'h41fad6f4, 32'h416b33ac} /* (3, 28, 10) {real, imag} */,
  {32'h42044bd0, 32'h41245ef1} /* (3, 28, 9) {real, imag} */,
  {32'h41b34eff, 32'h41a77631} /* (3, 28, 8) {real, imag} */,
  {32'h421125c5, 32'h41651c9b} /* (3, 28, 7) {real, imag} */,
  {32'h423cfd13, 32'h42060dba} /* (3, 28, 6) {real, imag} */,
  {32'h42270732, 32'h422ad2a6} /* (3, 28, 5) {real, imag} */,
  {32'h409e8468, 32'h41a34caa} /* (3, 28, 4) {real, imag} */,
  {32'hc055cd98, 32'hc11f1e0c} /* (3, 28, 3) {real, imag} */,
  {32'h4151f5ce, 32'hc1424152} /* (3, 28, 2) {real, imag} */,
  {32'h419f2590, 32'h410439da} /* (3, 28, 1) {real, imag} */,
  {32'h415c8545, 32'h41410f38} /* (3, 28, 0) {real, imag} */,
  {32'hc029653e, 32'hc16e8495} /* (3, 27, 31) {real, imag} */,
  {32'hc1440e38, 32'hc197e27a} /* (3, 27, 30) {real, imag} */,
  {32'hc14f5ad2, 32'hc19417bf} /* (3, 27, 29) {real, imag} */,
  {32'h41517313, 32'hc193293a} /* (3, 27, 28) {real, imag} */,
  {32'h40818cd4, 32'hc1964867} /* (3, 27, 27) {real, imag} */,
  {32'hc1550f24, 32'hc18b8605} /* (3, 27, 26) {real, imag} */,
  {32'h3fa63870, 32'hc197dd73} /* (3, 27, 25) {real, imag} */,
  {32'h41113e00, 32'hc15403ae} /* (3, 27, 24) {real, imag} */,
  {32'h40d41c85, 32'hc1eb80a6} /* (3, 27, 23) {real, imag} */,
  {32'hc005597a, 32'hc2246000} /* (3, 27, 22) {real, imag} */,
  {32'hc0fa9591, 32'hc1fe01c4} /* (3, 27, 21) {real, imag} */,
  {32'h40a1a86b, 32'hc10b5f98} /* (3, 27, 20) {real, imag} */,
  {32'h418d5efe, 32'h413e63a0} /* (3, 27, 19) {real, imag} */,
  {32'h417591a4, 32'h41a194df} /* (3, 27, 18) {real, imag} */,
  {32'h40801afc, 32'h41849dbe} /* (3, 27, 17) {real, imag} */,
  {32'hc0e460c4, 32'hc0f7f4c2} /* (3, 27, 16) {real, imag} */,
  {32'h41588c13, 32'hc097cc2a} /* (3, 27, 15) {real, imag} */,
  {32'h41034192, 32'hc03ab8fc} /* (3, 27, 14) {real, imag} */,
  {32'h40dd1748, 32'h41c37009} /* (3, 27, 13) {real, imag} */,
  {32'h4127c29a, 32'h420e9f9b} /* (3, 27, 12) {real, imag} */,
  {32'h41558616, 32'h41999497} /* (3, 27, 11) {real, imag} */,
  {32'h4170bcca, 32'hc11829c9} /* (3, 27, 10) {real, imag} */,
  {32'h40ea1cb0, 32'hc15060e8} /* (3, 27, 9) {real, imag} */,
  {32'h411449b6, 32'hc1ee3f0d} /* (3, 27, 8) {real, imag} */,
  {32'h415ad828, 32'hc2057b65} /* (3, 27, 7) {real, imag} */,
  {32'h4103ebbd, 32'hc13baea3} /* (3, 27, 6) {real, imag} */,
  {32'h414810e0, 32'hc0cffc77} /* (3, 27, 5) {real, imag} */,
  {32'hc0bf9aa6, 32'hc163b999} /* (3, 27, 4) {real, imag} */,
  {32'hc1428c7a, 32'hc216110a} /* (3, 27, 3) {real, imag} */,
  {32'hc128fc74, 32'hc1eb2c2e} /* (3, 27, 2) {real, imag} */,
  {32'hc1032e9e, 32'hc19ae5b8} /* (3, 27, 1) {real, imag} */,
  {32'hbf32c438, 32'hc16b9e62} /* (3, 27, 0) {real, imag} */,
  {32'h413c9235, 32'hc053895c} /* (3, 26, 31) {real, imag} */,
  {32'h40bc2338, 32'hc1c059f6} /* (3, 26, 30) {real, imag} */,
  {32'hc12115ba, 32'hc1a83e65} /* (3, 26, 29) {real, imag} */,
  {32'h404f87d8, 32'hc153acd8} /* (3, 26, 28) {real, imag} */,
  {32'h3f7d7be0, 32'hc0a151ff} /* (3, 26, 27) {real, imag} */,
  {32'hc08682b4, 32'h40c636c6} /* (3, 26, 26) {real, imag} */,
  {32'h40c9740a, 32'hc1840a71} /* (3, 26, 25) {real, imag} */,
  {32'h4161a52a, 32'h4008d036} /* (3, 26, 24) {real, imag} */,
  {32'h41436c2e, 32'h418ed3ce} /* (3, 26, 23) {real, imag} */,
  {32'h4087bd6f, 32'hc023b5e0} /* (3, 26, 22) {real, imag} */,
  {32'h40f22f3c, 32'hc139a9b8} /* (3, 26, 21) {real, imag} */,
  {32'hbfe1191c, 32'hc0241402} /* (3, 26, 20) {real, imag} */,
  {32'hc0561aa6, 32'h4117a2f6} /* (3, 26, 19) {real, imag} */,
  {32'hc031d114, 32'hc078a80e} /* (3, 26, 18) {real, imag} */,
  {32'hbf98bf54, 32'hc18b5d38} /* (3, 26, 17) {real, imag} */,
  {32'h40e0989c, 32'h404a6e7e} /* (3, 26, 16) {real, imag} */,
  {32'hc0b825e6, 32'h4199a2c2} /* (3, 26, 15) {real, imag} */,
  {32'hc155801b, 32'h402ad0bc} /* (3, 26, 14) {real, imag} */,
  {32'h416f7f4a, 32'hc163d4bf} /* (3, 26, 13) {real, imag} */,
  {32'h4137d175, 32'hc0ef6806} /* (3, 26, 12) {real, imag} */,
  {32'hc0334efe, 32'hc0d8e442} /* (3, 26, 11) {real, imag} */,
  {32'hc119723a, 32'h4038d010} /* (3, 26, 10) {real, imag} */,
  {32'h40d89c5d, 32'h411dae4d} /* (3, 26, 9) {real, imag} */,
  {32'h400e98a0, 32'hc1186c4f} /* (3, 26, 8) {real, imag} */,
  {32'h3d2b26c0, 32'hc0e34634} /* (3, 26, 7) {real, imag} */,
  {32'h4144b610, 32'h410cb380} /* (3, 26, 6) {real, imag} */,
  {32'hc11006c6, 32'h41139186} /* (3, 26, 5) {real, imag} */,
  {32'hc16c467d, 32'hc066812c} /* (3, 26, 4) {real, imag} */,
  {32'hc1168f64, 32'hc12ed178} /* (3, 26, 3) {real, imag} */,
  {32'h4083f15b, 32'hc1bb0006} /* (3, 26, 2) {real, imag} */,
  {32'h417f534b, 32'h40692b18} /* (3, 26, 1) {real, imag} */,
  {32'h41159aab, 32'h40c92ad9} /* (3, 26, 0) {real, imag} */,
  {32'hc03330fb, 32'h410e7844} /* (3, 25, 31) {real, imag} */,
  {32'hc047ac98, 32'h410326f3} /* (3, 25, 30) {real, imag} */,
  {32'h3f097b10, 32'h4132f424} /* (3, 25, 29) {real, imag} */,
  {32'hc04d27e6, 32'h40e43ffa} /* (3, 25, 28) {real, imag} */,
  {32'h402a7413, 32'h413b0d4c} /* (3, 25, 27) {real, imag} */,
  {32'hc0c9227a, 32'h4194ece6} /* (3, 25, 26) {real, imag} */,
  {32'h3ffa7cce, 32'h418fdb3e} /* (3, 25, 25) {real, imag} */,
  {32'h4199b198, 32'h3f6f8670} /* (3, 25, 24) {real, imag} */,
  {32'h4185d4c2, 32'hbe4cc340} /* (3, 25, 23) {real, imag} */,
  {32'h4000ba16, 32'h403d476c} /* (3, 25, 22) {real, imag} */,
  {32'hc16cb408, 32'h402db190} /* (3, 25, 21) {real, imag} */,
  {32'hc069dcda, 32'h40a31e1e} /* (3, 25, 20) {real, imag} */,
  {32'hc06188f9, 32'hbecbc860} /* (3, 25, 19) {real, imag} */,
  {32'hc114aafc, 32'h4150aca8} /* (3, 25, 18) {real, imag} */,
  {32'h40a7c358, 32'h40c71ab6} /* (3, 25, 17) {real, imag} */,
  {32'hc1452ecd, 32'h3fca1120} /* (3, 25, 16) {real, imag} */,
  {32'hc0818c44, 32'hc0935409} /* (3, 25, 15) {real, imag} */,
  {32'hc1048f9a, 32'h4092fdf4} /* (3, 25, 14) {real, imag} */,
  {32'hc1d03c53, 32'hc1276c20} /* (3, 25, 13) {real, imag} */,
  {32'hc10c2bcc, 32'hc0e5d0ef} /* (3, 25, 12) {real, imag} */,
  {32'h41b61bd8, 32'hc0738cd2} /* (3, 25, 11) {real, imag} */,
  {32'h412b23aa, 32'hc0b474a6} /* (3, 25, 10) {real, imag} */,
  {32'h4176b637, 32'hc1979e05} /* (3, 25, 9) {real, imag} */,
  {32'h416c5416, 32'hc15077be} /* (3, 25, 8) {real, imag} */,
  {32'h410ab180, 32'h416d698b} /* (3, 25, 7) {real, imag} */,
  {32'hc04e8ac5, 32'h41d46598} /* (3, 25, 6) {real, imag} */,
  {32'hc0e88ea3, 32'h407e9ff4} /* (3, 25, 5) {real, imag} */,
  {32'hc072caf0, 32'h40bd6cc1} /* (3, 25, 4) {real, imag} */,
  {32'h411a00fe, 32'h41d8a7ac} /* (3, 25, 3) {real, imag} */,
  {32'h418e154b, 32'h41f9e3c4} /* (3, 25, 2) {real, imag} */,
  {32'h41903968, 32'h41bddcaf} /* (3, 25, 1) {real, imag} */,
  {32'h4059ac84, 32'h40dda965} /* (3, 25, 0) {real, imag} */,
  {32'hc13fcb04, 32'h3f7cd3e0} /* (3, 24, 31) {real, imag} */,
  {32'hc146460c, 32'h4124e052} /* (3, 24, 30) {real, imag} */,
  {32'hc003293e, 32'hc16d16e8} /* (3, 24, 29) {real, imag} */,
  {32'h40d1adec, 32'hc1bde3c2} /* (3, 24, 28) {real, imag} */,
  {32'h41823c8f, 32'hc18d2504} /* (3, 24, 27) {real, imag} */,
  {32'h412b3269, 32'hc0f800ee} /* (3, 24, 26) {real, imag} */,
  {32'hc0d1ce62, 32'hc18f317a} /* (3, 24, 25) {real, imag} */,
  {32'hc18d5d3e, 32'hc1ca6200} /* (3, 24, 24) {real, imag} */,
  {32'hc116e474, 32'hc1935794} /* (3, 24, 23) {real, imag} */,
  {32'hc09d4b1c, 32'hc14c560c} /* (3, 24, 22) {real, imag} */,
  {32'hc1606655, 32'hc1379efb} /* (3, 24, 21) {real, imag} */,
  {32'hc1980ec0, 32'h418b8c71} /* (3, 24, 20) {real, imag} */,
  {32'hc0be7418, 32'h4195fe91} /* (3, 24, 19) {real, imag} */,
  {32'hbfd1048c, 32'h41a1e694} /* (3, 24, 18) {real, imag} */,
  {32'hc0fcb35a, 32'h41335966} /* (3, 24, 17) {real, imag} */,
  {32'h415a7c3f, 32'h411e8c60} /* (3, 24, 16) {real, imag} */,
  {32'h4200a23b, 32'h40cb2f78} /* (3, 24, 15) {real, imag} */,
  {32'h419f74d6, 32'h405a9e80} /* (3, 24, 14) {real, imag} */,
  {32'h4045f4bb, 32'h407064e1} /* (3, 24, 13) {real, imag} */,
  {32'h416706a2, 32'h40fb0c18} /* (3, 24, 12) {real, imag} */,
  {32'h40483478, 32'h41bfc882} /* (3, 24, 11) {real, imag} */,
  {32'hbe8cae80, 32'h40e58fb4} /* (3, 24, 10) {real, imag} */,
  {32'h41aae2b8, 32'h40553bee} /* (3, 24, 9) {real, imag} */,
  {32'h4086dec4, 32'h4146c116} /* (3, 24, 8) {real, imag} */,
  {32'hc11b4159, 32'hbfb02215} /* (3, 24, 7) {real, imag} */,
  {32'hc0c4da00, 32'hc1bd7d4c} /* (3, 24, 6) {real, imag} */,
  {32'hc11b8db7, 32'hc12a2ada} /* (3, 24, 5) {real, imag} */,
  {32'hc125a118, 32'hc1b4b82e} /* (3, 24, 4) {real, imag} */,
  {32'hc091455e, 32'hc1621ecd} /* (3, 24, 3) {real, imag} */,
  {32'hc01ffdfa, 32'hc1012713} /* (3, 24, 2) {real, imag} */,
  {32'h410cd107, 32'hc195307b} /* (3, 24, 1) {real, imag} */,
  {32'h3fb67714, 32'hc18633cd} /* (3, 24, 0) {real, imag} */,
  {32'hc0d6c3ee, 32'hc11fc18a} /* (3, 23, 31) {real, imag} */,
  {32'h40dea8b6, 32'hbf4950b8} /* (3, 23, 30) {real, imag} */,
  {32'h40411ac0, 32'hc02fdeb8} /* (3, 23, 29) {real, imag} */,
  {32'h40c92887, 32'hbf4c36e8} /* (3, 23, 28) {real, imag} */,
  {32'hbf99e2f8, 32'hc0938e50} /* (3, 23, 27) {real, imag} */,
  {32'hc0c56bcd, 32'hc0b51c78} /* (3, 23, 26) {real, imag} */,
  {32'hbf477020, 32'hbea52ae8} /* (3, 23, 25) {real, imag} */,
  {32'hc0989cea, 32'h3fc955e8} /* (3, 23, 24) {real, imag} */,
  {32'hbf9c1bb4, 32'h4029a3d8} /* (3, 23, 23) {real, imag} */,
  {32'hbf005ab8, 32'hc0bc9a83} /* (3, 23, 22) {real, imag} */,
  {32'hbfe8f480, 32'hc14d2977} /* (3, 23, 21) {real, imag} */,
  {32'hc15388dc, 32'hc1876cab} /* (3, 23, 20) {real, imag} */,
  {32'hc0039783, 32'hbfc23bf8} /* (3, 23, 19) {real, imag} */,
  {32'hbfcc202c, 32'h4122e88a} /* (3, 23, 18) {real, imag} */,
  {32'hc1117571, 32'hc02332cc} /* (3, 23, 17) {real, imag} */,
  {32'hc10c7263, 32'hc0b01b9a} /* (3, 23, 16) {real, imag} */,
  {32'h40974378, 32'hc0b3c94d} /* (3, 23, 15) {real, imag} */,
  {32'hbf53d2b0, 32'hc0a2d7c6} /* (3, 23, 14) {real, imag} */,
  {32'hbf9d9a54, 32'h411a157e} /* (3, 23, 13) {real, imag} */,
  {32'hbf7d74b0, 32'h4140e230} /* (3, 23, 12) {real, imag} */,
  {32'h4092734e, 32'h41bea00d} /* (3, 23, 11) {real, imag} */,
  {32'h41889bac, 32'h417a4f46} /* (3, 23, 10) {real, imag} */,
  {32'h408597fa, 32'h41091e6e} /* (3, 23, 9) {real, imag} */,
  {32'h40e5cd4f, 32'h414d943c} /* (3, 23, 8) {real, imag} */,
  {32'h414eb605, 32'hc0c92c7a} /* (3, 23, 7) {real, imag} */,
  {32'h410b7cef, 32'h413d21ad} /* (3, 23, 6) {real, imag} */,
  {32'hbff71174, 32'h4178818e} /* (3, 23, 5) {real, imag} */,
  {32'hbe37ce00, 32'h40e22298} /* (3, 23, 4) {real, imag} */,
  {32'h40faa0e5, 32'h40e3b23e} /* (3, 23, 3) {real, imag} */,
  {32'h414b2500, 32'h40e45ab1} /* (3, 23, 2) {real, imag} */,
  {32'h40ef8a12, 32'hc029b101} /* (3, 23, 1) {real, imag} */,
  {32'h3f4fa034, 32'h3dc35b40} /* (3, 23, 0) {real, imag} */,
  {32'h41539164, 32'h4070b998} /* (3, 22, 31) {real, imag} */,
  {32'h41a36873, 32'h40c2c334} /* (3, 22, 30) {real, imag} */,
  {32'h41be8156, 32'h413ad11a} /* (3, 22, 29) {real, imag} */,
  {32'hc039231d, 32'h40eb68f7} /* (3, 22, 28) {real, imag} */,
  {32'hc1857b61, 32'h415598b8} /* (3, 22, 27) {real, imag} */,
  {32'hc19c9326, 32'h40809dde} /* (3, 22, 26) {real, imag} */,
  {32'hc0975728, 32'hbf519238} /* (3, 22, 25) {real, imag} */,
  {32'h41296022, 32'h405c4ca6} /* (3, 22, 24) {real, imag} */,
  {32'h410ac9c6, 32'hc0db6916} /* (3, 22, 23) {real, imag} */,
  {32'h41837d14, 32'hc126f22f} /* (3, 22, 22) {real, imag} */,
  {32'h41bd41f6, 32'hc0ddb022} /* (3, 22, 21) {real, imag} */,
  {32'h412f12ce, 32'hc142f8ca} /* (3, 22, 20) {real, imag} */,
  {32'hc0a3b139, 32'hc10d660e} /* (3, 22, 19) {real, imag} */,
  {32'hc105d71d, 32'hbf3269c8} /* (3, 22, 18) {real, imag} */,
  {32'h407cc7ea, 32'hbf770e78} /* (3, 22, 17) {real, imag} */,
  {32'h40062e4d, 32'h40f73be5} /* (3, 22, 16) {real, imag} */,
  {32'hc07d57a3, 32'hc1128560} /* (3, 22, 15) {real, imag} */,
  {32'hc14e64c0, 32'hc0c5ccb0} /* (3, 22, 14) {real, imag} */,
  {32'hc10ce7b8, 32'h40d6d748} /* (3, 22, 13) {real, imag} */,
  {32'h405625b8, 32'h411eb793} /* (3, 22, 12) {real, imag} */,
  {32'hc0ac4382, 32'h4128d523} /* (3, 22, 11) {real, imag} */,
  {32'hc081d2b3, 32'h4145d4f4} /* (3, 22, 10) {real, imag} */,
  {32'h408d3569, 32'h41d8b178} /* (3, 22, 9) {real, imag} */,
  {32'h40b2ab7a, 32'h414420de} /* (3, 22, 8) {real, imag} */,
  {32'h4169d372, 32'h410dd964} /* (3, 22, 7) {real, imag} */,
  {32'h41207a00, 32'h41173fe0} /* (3, 22, 6) {real, imag} */,
  {32'hbf6f91d0, 32'hc0973ee9} /* (3, 22, 5) {real, imag} */,
  {32'hbf4840d0, 32'hc0b6bda0} /* (3, 22, 4) {real, imag} */,
  {32'h405ff8b3, 32'hc0f719a7} /* (3, 22, 3) {real, imag} */,
  {32'hc091d09e, 32'hc02fd500} /* (3, 22, 2) {real, imag} */,
  {32'hc107b3bf, 32'hc0d9e484} /* (3, 22, 1) {real, imag} */,
  {32'hbfe0ff92, 32'hbfec7bb8} /* (3, 22, 0) {real, imag} */,
  {32'hc00883c2, 32'h40de2bf9} /* (3, 21, 31) {real, imag} */,
  {32'hc0a05a03, 32'h411b3a83} /* (3, 21, 30) {real, imag} */,
  {32'h40fced40, 32'h401a133c} /* (3, 21, 29) {real, imag} */,
  {32'hbf0addc0, 32'hc119b70e} /* (3, 21, 28) {real, imag} */,
  {32'hc1614e2f, 32'hc13d80a0} /* (3, 21, 27) {real, imag} */,
  {32'hc0f7dd6a, 32'hc0eb702b} /* (3, 21, 26) {real, imag} */,
  {32'hc12bdadc, 32'hc157103e} /* (3, 21, 25) {real, imag} */,
  {32'hc0dfdfa2, 32'hc15400d6} /* (3, 21, 24) {real, imag} */,
  {32'hc0d51f31, 32'hc138bd1b} /* (3, 21, 23) {real, imag} */,
  {32'h40866a2c, 32'h4030aad8} /* (3, 21, 22) {real, imag} */,
  {32'hc03b68ba, 32'h40e4ec76} /* (3, 21, 21) {real, imag} */,
  {32'h3ee37cf0, 32'hbe15ce90} /* (3, 21, 20) {real, imag} */,
  {32'hbfa8a6b8, 32'hc0fd68de} /* (3, 21, 19) {real, imag} */,
  {32'hc06c8612, 32'hc09b633a} /* (3, 21, 18) {real, imag} */,
  {32'h40332114, 32'h40b50c1a} /* (3, 21, 17) {real, imag} */,
  {32'h40b452a8, 32'h40ffc95e} /* (3, 21, 16) {real, imag} */,
  {32'h40398278, 32'h4158c978} /* (3, 21, 15) {real, imag} */,
  {32'hc061817e, 32'h412be556} /* (3, 21, 14) {real, imag} */,
  {32'h412a2f9a, 32'hbf934a3c} /* (3, 21, 13) {real, imag} */,
  {32'h40fab607, 32'hc08456ca} /* (3, 21, 12) {real, imag} */,
  {32'h40a392fe, 32'hc112f6d7} /* (3, 21, 11) {real, imag} */,
  {32'hc0730d7a, 32'hc07542d6} /* (3, 21, 10) {real, imag} */,
  {32'hc14cbd84, 32'h40e74bb3} /* (3, 21, 9) {real, imag} */,
  {32'hc0a7f937, 32'hbd3a6980} /* (3, 21, 8) {real, imag} */,
  {32'hc064c52a, 32'hbfb70be0} /* (3, 21, 7) {real, imag} */,
  {32'hc11897c2, 32'hc00107a0} /* (3, 21, 6) {real, imag} */,
  {32'hc122caad, 32'hc0def0e5} /* (3, 21, 5) {real, imag} */,
  {32'hc14ec6ad, 32'hc1082d85} /* (3, 21, 4) {real, imag} */,
  {32'hc1782ab3, 32'hc08ae232} /* (3, 21, 3) {real, imag} */,
  {32'hc09d19bd, 32'hc03e74d0} /* (3, 21, 2) {real, imag} */,
  {32'h40835530, 32'hc04ee700} /* (3, 21, 1) {real, imag} */,
  {32'h3f1641e8, 32'hc0088bae} /* (3, 21, 0) {real, imag} */,
  {32'h3f383e88, 32'hbf1f0cf4} /* (3, 20, 31) {real, imag} */,
  {32'hbfeab158, 32'h4079068e} /* (3, 20, 30) {real, imag} */,
  {32'h3f872dd4, 32'h404df0a6} /* (3, 20, 29) {real, imag} */,
  {32'hbfda926c, 32'h40a86797} /* (3, 20, 28) {real, imag} */,
  {32'hbf085790, 32'hbf905d64} /* (3, 20, 27) {real, imag} */,
  {32'h40e8ad03, 32'h400c56f6} /* (3, 20, 26) {real, imag} */,
  {32'h40c4cea4, 32'h40f0f4d8} /* (3, 20, 25) {real, imag} */,
  {32'h40b656b9, 32'h415383ad} /* (3, 20, 24) {real, imag} */,
  {32'h40b432f2, 32'h4064dd51} /* (3, 20, 23) {real, imag} */,
  {32'h4086a333, 32'hc1122e12} /* (3, 20, 22) {real, imag} */,
  {32'h40854ec0, 32'hc0bb5caf} /* (3, 20, 21) {real, imag} */,
  {32'h3ed81e80, 32'hc062af90} /* (3, 20, 20) {real, imag} */,
  {32'hbeaf1360, 32'hbf073c46} /* (3, 20, 19) {real, imag} */,
  {32'hbf84e2d2, 32'hc1490664} /* (3, 20, 18) {real, imag} */,
  {32'hc0a9f0b7, 32'hc15751fa} /* (3, 20, 17) {real, imag} */,
  {32'h40841385, 32'h3f960510} /* (3, 20, 16) {real, imag} */,
  {32'hbdc32310, 32'h41094b9a} /* (3, 20, 15) {real, imag} */,
  {32'hc032e666, 32'hc0a103d4} /* (3, 20, 14) {real, imag} */,
  {32'h40ea4cb5, 32'hc0fd522d} /* (3, 20, 13) {real, imag} */,
  {32'h4123711c, 32'hbfdcd192} /* (3, 20, 12) {real, imag} */,
  {32'h4139ebaa, 32'h402b37df} /* (3, 20, 11) {real, imag} */,
  {32'h3ff9094c, 32'hbf9d4cf4} /* (3, 20, 10) {real, imag} */,
  {32'h3fa1b562, 32'hc0bb7471} /* (3, 20, 9) {real, imag} */,
  {32'h40293734, 32'hc15ab9d0} /* (3, 20, 8) {real, imag} */,
  {32'h3eddb418, 32'hc0b5affc} /* (3, 20, 7) {real, imag} */,
  {32'hc0bf5ac6, 32'h4013970d} /* (3, 20, 6) {real, imag} */,
  {32'hc108192e, 32'hc00dae2e} /* (3, 20, 5) {real, imag} */,
  {32'hc020f6b4, 32'hbfb4ec22} /* (3, 20, 4) {real, imag} */,
  {32'hc081d8d0, 32'hc064f2ca} /* (3, 20, 3) {real, imag} */,
  {32'hc004df3d, 32'h40d3f415} /* (3, 20, 2) {real, imag} */,
  {32'h406e25b8, 32'h407ea170} /* (3, 20, 1) {real, imag} */,
  {32'h40aa172f, 32'hc0c2f67e} /* (3, 20, 0) {real, imag} */,
  {32'hbf5914ba, 32'hc0013248} /* (3, 19, 31) {real, imag} */,
  {32'hbfd28bd8, 32'hc00bdf22} /* (3, 19, 30) {real, imag} */,
  {32'h3fc57990, 32'hc09bc5ff} /* (3, 19, 29) {real, imag} */,
  {32'h40876c36, 32'hc0b3430d} /* (3, 19, 28) {real, imag} */,
  {32'hbf6cb104, 32'hc085b80b} /* (3, 19, 27) {real, imag} */,
  {32'h3fdf89ee, 32'h3fd54ff2} /* (3, 19, 26) {real, imag} */,
  {32'h41139d4e, 32'h40225fdb} /* (3, 19, 25) {real, imag} */,
  {32'h4090b9b3, 32'hbfceeb88} /* (3, 19, 24) {real, imag} */,
  {32'hbfa43dd0, 32'hc04df1bc} /* (3, 19, 23) {real, imag} */,
  {32'h4006659d, 32'h402d2f72} /* (3, 19, 22) {real, imag} */,
  {32'h40af1cb9, 32'h408e77d6} /* (3, 19, 21) {real, imag} */,
  {32'hbfc5a410, 32'h4082f5c0} /* (3, 19, 20) {real, imag} */,
  {32'hc1295453, 32'hc07f2fa4} /* (3, 19, 19) {real, imag} */,
  {32'hc046016a, 32'hc0cde11b} /* (3, 19, 18) {real, imag} */,
  {32'h3f51e7c0, 32'hbfc92e76} /* (3, 19, 17) {real, imag} */,
  {32'hc130b367, 32'hbf951c1c} /* (3, 19, 16) {real, imag} */,
  {32'hc131c703, 32'hbdc58760} /* (3, 19, 15) {real, imag} */,
  {32'h400f4ef8, 32'hbfc63038} /* (3, 19, 14) {real, imag} */,
  {32'hbf8e2eae, 32'hbedf9860} /* (3, 19, 13) {real, imag} */,
  {32'hc09fde08, 32'h40cbf454} /* (3, 19, 12) {real, imag} */,
  {32'h3f329c68, 32'h3f80e322} /* (3, 19, 11) {real, imag} */,
  {32'h40447da8, 32'hbf0e9948} /* (3, 19, 10) {real, imag} */,
  {32'hc0564a74, 32'h3ff1cbc8} /* (3, 19, 9) {real, imag} */,
  {32'hc0ed4624, 32'h408b2578} /* (3, 19, 8) {real, imag} */,
  {32'hc04b90ac, 32'h404a9c0a} /* (3, 19, 7) {real, imag} */,
  {32'hbfbfbb1e, 32'h40987bf0} /* (3, 19, 6) {real, imag} */,
  {32'h3f5f9c38, 32'h41291cb0} /* (3, 19, 5) {real, imag} */,
  {32'h406b33fc, 32'h40e54751} /* (3, 19, 4) {real, imag} */,
  {32'h404aa205, 32'h40961670} /* (3, 19, 3) {real, imag} */,
  {32'h40375f2d, 32'h407c830d} /* (3, 19, 2) {real, imag} */,
  {32'h3e69dde0, 32'h405cb42c} /* (3, 19, 1) {real, imag} */,
  {32'hc085bd72, 32'h40e2d296} /* (3, 19, 0) {real, imag} */,
  {32'hc0bf158c, 32'h40ae247d} /* (3, 18, 31) {real, imag} */,
  {32'hc10167e2, 32'h3fe35270} /* (3, 18, 30) {real, imag} */,
  {32'hc12146a8, 32'h3f0d7d30} /* (3, 18, 29) {real, imag} */,
  {32'hc02c6570, 32'h4080e19d} /* (3, 18, 28) {real, imag} */,
  {32'hbea0ee70, 32'h3f3b3e48} /* (3, 18, 27) {real, imag} */,
  {32'hc01035a6, 32'hbfbeac00} /* (3, 18, 26) {real, imag} */,
  {32'hc0a35167, 32'hc042cce8} /* (3, 18, 25) {real, imag} */,
  {32'hc08bd3fa, 32'hbf8fc618} /* (3, 18, 24) {real, imag} */,
  {32'hc067bd42, 32'hbf7850d0} /* (3, 18, 23) {real, imag} */,
  {32'hc04dfc74, 32'hc0950919} /* (3, 18, 22) {real, imag} */,
  {32'hc126b36f, 32'hc0876543} /* (3, 18, 21) {real, imag} */,
  {32'hbf5935c0, 32'h406b3571} /* (3, 18, 20) {real, imag} */,
  {32'h40e7ca78, 32'h411e1ba0} /* (3, 18, 19) {real, imag} */,
  {32'hbe7cdc40, 32'h40ae4010} /* (3, 18, 18) {real, imag} */,
  {32'hbe20ab40, 32'h3fc79bc0} /* (3, 18, 17) {real, imag} */,
  {32'h3fcecd78, 32'h40fce143} /* (3, 18, 16) {real, imag} */,
  {32'hbd28df40, 32'h40aeb122} /* (3, 18, 15) {real, imag} */,
  {32'h4055269e, 32'h3f463b58} /* (3, 18, 14) {real, imag} */,
  {32'h40b93fec, 32'hc0191296} /* (3, 18, 13) {real, imag} */,
  {32'h409767e0, 32'h4008ebb8} /* (3, 18, 12) {real, imag} */,
  {32'hbff4e5a6, 32'h40a0e2ef} /* (3, 18, 11) {real, imag} */,
  {32'h3f87dfa0, 32'hc0ac308c} /* (3, 18, 10) {real, imag} */,
  {32'h3ddb6880, 32'hc0bd5029} /* (3, 18, 9) {real, imag} */,
  {32'h40347340, 32'h3f8a4b5e} /* (3, 18, 8) {real, imag} */,
  {32'hc02375fc, 32'hc08c2ea8} /* (3, 18, 7) {real, imag} */,
  {32'hc06bef70, 32'hc0f92d6f} /* (3, 18, 6) {real, imag} */,
  {32'hbec65570, 32'h40809c91} /* (3, 18, 5) {real, imag} */,
  {32'hc02af514, 32'h404734e2} /* (3, 18, 4) {real, imag} */,
  {32'hc052c34b, 32'hc00f3c0a} /* (3, 18, 3) {real, imag} */,
  {32'hc0fb5c98, 32'h3f6130ac} /* (3, 18, 2) {real, imag} */,
  {32'hc12a895d, 32'h3f609354} /* (3, 18, 1) {real, imag} */,
  {32'hc0e252b2, 32'hbffbb64f} /* (3, 18, 0) {real, imag} */,
  {32'h4012ee2d, 32'hbfeef05e} /* (3, 17, 31) {real, imag} */,
  {32'hc0809743, 32'h4040a5fe} /* (3, 17, 30) {real, imag} */,
  {32'hbea62084, 32'h4080ee48} /* (3, 17, 29) {real, imag} */,
  {32'h3f466cd2, 32'hbfe2e318} /* (3, 17, 28) {real, imag} */,
  {32'h409f22d8, 32'hbfd9cfd8} /* (3, 17, 27) {real, imag} */,
  {32'h3fcb77d0, 32'hc0214ba0} /* (3, 17, 26) {real, imag} */,
  {32'hc040366c, 32'hc0b263cc} /* (3, 17, 25) {real, imag} */,
  {32'hc06d0525, 32'hc08dc565} /* (3, 17, 24) {real, imag} */,
  {32'hc08ea357, 32'hc093d7ad} /* (3, 17, 23) {real, imag} */,
  {32'hc0e0a1ae, 32'h3f64e7f0} /* (3, 17, 22) {real, imag} */,
  {32'hc09aaf81, 32'h3d934d30} /* (3, 17, 21) {real, imag} */,
  {32'hc089c5e8, 32'h406bed15} /* (3, 17, 20) {real, imag} */,
  {32'hc09361b0, 32'h4079b8e0} /* (3, 17, 19) {real, imag} */,
  {32'hc0879a70, 32'h3eff3c80} /* (3, 17, 18) {real, imag} */,
  {32'hc0bdc2d0, 32'h400c2edc} /* (3, 17, 17) {real, imag} */,
  {32'hc0e3fe7e, 32'hbf8f00b0} /* (3, 17, 16) {real, imag} */,
  {32'hbffa12ec, 32'hc025ab69} /* (3, 17, 15) {real, imag} */,
  {32'hbfb2b8a0, 32'h3f7cb0ec} /* (3, 17, 14) {real, imag} */,
  {32'hbd5407c0, 32'h40cfcec0} /* (3, 17, 13) {real, imag} */,
  {32'hc0c2a656, 32'h404d5f68} /* (3, 17, 12) {real, imag} */,
  {32'hc09fe6c7, 32'h403f0028} /* (3, 17, 11) {real, imag} */,
  {32'hc04203b0, 32'h40606de6} /* (3, 17, 10) {real, imag} */,
  {32'hbfd5fb3e, 32'h3fa19d40} /* (3, 17, 9) {real, imag} */,
  {32'h3ebc9fa0, 32'h40467258} /* (3, 17, 8) {real, imag} */,
  {32'h40f307ca, 32'h4068023c} /* (3, 17, 7) {real, imag} */,
  {32'h40aa712a, 32'h3f6c07c0} /* (3, 17, 6) {real, imag} */,
  {32'h4066ef90, 32'h402627ba} /* (3, 17, 5) {real, imag} */,
  {32'h40f2687a, 32'hbf181360} /* (3, 17, 4) {real, imag} */,
  {32'hbfb864c0, 32'hc03730e8} /* (3, 17, 3) {real, imag} */,
  {32'hc04d1bb2, 32'h40510d18} /* (3, 17, 2) {real, imag} */,
  {32'hbf5d1f24, 32'h40184cd6} /* (3, 17, 1) {real, imag} */,
  {32'hbf38d1ba, 32'hbf4712f4} /* (3, 17, 0) {real, imag} */,
  {32'hbe912f00, 32'h3f293848} /* (3, 16, 31) {real, imag} */,
  {32'h3f5ccca0, 32'h3eb70180} /* (3, 16, 30) {real, imag} */,
  {32'hc04b558a, 32'h3fd401e0} /* (3, 16, 29) {real, imag} */,
  {32'h3f1b2ec0, 32'hc01ef058} /* (3, 16, 28) {real, imag} */,
  {32'hc010df60, 32'hc0694400} /* (3, 16, 27) {real, imag} */,
  {32'hbf0a7f34, 32'hc072e8f0} /* (3, 16, 26) {real, imag} */,
  {32'h4090f5b4, 32'hc0def6f8} /* (3, 16, 25) {real, imag} */,
  {32'h3faf674b, 32'hc0a3c1f8} /* (3, 16, 24) {real, imag} */,
  {32'hbff7a770, 32'hbf7e1240} /* (3, 16, 23) {real, imag} */,
  {32'hc0a5845c, 32'h4071b8c0} /* (3, 16, 22) {real, imag} */,
  {32'hbf60d220, 32'h3f1aa940} /* (3, 16, 21) {real, imag} */,
  {32'h4074736a, 32'h4025af58} /* (3, 16, 20) {real, imag} */,
  {32'h40787e24, 32'h405c9340} /* (3, 16, 19) {real, imag} */,
  {32'hbffc29c8, 32'hbe792f80} /* (3, 16, 18) {real, imag} */,
  {32'h3f7af190, 32'hc03943b0} /* (3, 16, 17) {real, imag} */,
  {32'h40867fea, 32'hc0a0b692} /* (3, 16, 16) {real, imag} */,
  {32'h3f900386, 32'hc085f13c} /* (3, 16, 15) {real, imag} */,
  {32'h3f6a5000, 32'hbf704680} /* (3, 16, 14) {real, imag} */,
  {32'hbe727840, 32'hbf2ac040} /* (3, 16, 13) {real, imag} */,
  {32'h4039d426, 32'hc04aabe0} /* (3, 16, 12) {real, imag} */,
  {32'h40abd032, 32'h3f86b720} /* (3, 16, 11) {real, imag} */,
  {32'h3fbd2550, 32'h400e54d8} /* (3, 16, 10) {real, imag} */,
  {32'hc04f57e2, 32'hbf9f2e98} /* (3, 16, 9) {real, imag} */,
  {32'hbfd20f48, 32'hc004ab79} /* (3, 16, 8) {real, imag} */,
  {32'h3f9370ef, 32'h3ef56b00} /* (3, 16, 7) {real, imag} */,
  {32'hc0313708, 32'hbf818248} /* (3, 16, 6) {real, imag} */,
  {32'h401707f0, 32'hbed25940} /* (3, 16, 5) {real, imag} */,
  {32'h40bd247a, 32'hc09eb04c} /* (3, 16, 4) {real, imag} */,
  {32'h3f6a2e40, 32'hc06bd990} /* (3, 16, 3) {real, imag} */,
  {32'h3fe4b6b4, 32'hc078c928} /* (3, 16, 2) {real, imag} */,
  {32'h40159386, 32'hc0a9d368} /* (3, 16, 1) {real, imag} */,
  {32'h3f034500, 32'hbfe579f8} /* (3, 16, 0) {real, imag} */,
  {32'h401325e3, 32'h3fd4261e} /* (3, 15, 31) {real, imag} */,
  {32'h4005cdc6, 32'h404a0482} /* (3, 15, 30) {real, imag} */,
  {32'h3fddda31, 32'hbeddca80} /* (3, 15, 29) {real, imag} */,
  {32'h3fb4fc37, 32'h3e61fec0} /* (3, 15, 28) {real, imag} */,
  {32'hc05c2240, 32'hbfd2f5a8} /* (3, 15, 27) {real, imag} */,
  {32'hc09280bc, 32'hc022e1c0} /* (3, 15, 26) {real, imag} */,
  {32'hc056f414, 32'hbf91fc10} /* (3, 15, 25) {real, imag} */,
  {32'hc06d9bbb, 32'h3e1410a0} /* (3, 15, 24) {real, imag} */,
  {32'hc0b65c59, 32'h409dd92d} /* (3, 15, 23) {real, imag} */,
  {32'hc0e2d45e, 32'hc0070bbc} /* (3, 15, 22) {real, imag} */,
  {32'h3cc38d00, 32'hbf16bc66} /* (3, 15, 21) {real, imag} */,
  {32'h40010b90, 32'h4023309b} /* (3, 15, 20) {real, imag} */,
  {32'h4017abb0, 32'hbf69e4c0} /* (3, 15, 19) {real, imag} */,
  {32'h410e9f10, 32'h40619ea0} /* (3, 15, 18) {real, imag} */,
  {32'h41218ab8, 32'h402d5f04} /* (3, 15, 17) {real, imag} */,
  {32'h408326c6, 32'hc0a6f724} /* (3, 15, 16) {real, imag} */,
  {32'h4108c21c, 32'hc0d249ec} /* (3, 15, 15) {real, imag} */,
  {32'h40cd2cf0, 32'h3f400494} /* (3, 15, 14) {real, imag} */,
  {32'h3eb055f8, 32'h3e931c08} /* (3, 15, 13) {real, imag} */,
  {32'hc0016d34, 32'h4023f658} /* (3, 15, 12) {real, imag} */,
  {32'h4083745b, 32'h403f20b8} /* (3, 15, 11) {real, imag} */,
  {32'hbef37a80, 32'hc08d1fb3} /* (3, 15, 10) {real, imag} */,
  {32'hc08b8350, 32'hc0929610} /* (3, 15, 9) {real, imag} */,
  {32'hc0eb7ef6, 32'hbf9338b0} /* (3, 15, 8) {real, imag} */,
  {32'hc120b96b, 32'hbfa5b478} /* (3, 15, 7) {real, imag} */,
  {32'hc097ecb2, 32'hbebd5400} /* (3, 15, 6) {real, imag} */,
  {32'h3eab0f40, 32'h3fbec10c} /* (3, 15, 5) {real, imag} */,
  {32'hc07fb7f4, 32'h404a2bd8} /* (3, 15, 4) {real, imag} */,
  {32'h40022340, 32'h402f49e8} /* (3, 15, 3) {real, imag} */,
  {32'h40c92651, 32'h405a7208} /* (3, 15, 2) {real, imag} */,
  {32'hbf4e075c, 32'h40bb0765} /* (3, 15, 1) {real, imag} */,
  {32'hc023ddde, 32'h409b2a66} /* (3, 15, 0) {real, imag} */,
  {32'hc08ed8f4, 32'h3ff7b40c} /* (3, 14, 31) {real, imag} */,
  {32'hc0498736, 32'h3f5c4d20} /* (3, 14, 30) {real, imag} */,
  {32'h400acbac, 32'h40b4dea2} /* (3, 14, 29) {real, imag} */,
  {32'h405e58e8, 32'h4090d9eb} /* (3, 14, 28) {real, imag} */,
  {32'h409f7ac9, 32'h3fcafb7c} /* (3, 14, 27) {real, imag} */,
  {32'h40382b3a, 32'h3fc54e80} /* (3, 14, 26) {real, imag} */,
  {32'h3fef1b24, 32'hbf648e60} /* (3, 14, 25) {real, imag} */,
  {32'h403da43c, 32'hc0407c54} /* (3, 14, 24) {real, imag} */,
  {32'h40ad0195, 32'hbebc2b60} /* (3, 14, 23) {real, imag} */,
  {32'h40c56bba, 32'h3f1de388} /* (3, 14, 22) {real, imag} */,
  {32'h40070b6c, 32'hc0ec4c2d} /* (3, 14, 21) {real, imag} */,
  {32'hc111816c, 32'hbfa7d3a2} /* (3, 14, 20) {real, imag} */,
  {32'hc0babe08, 32'h406a90c0} /* (3, 14, 19) {real, imag} */,
  {32'hc0812052, 32'h405e7c00} /* (3, 14, 18) {real, imag} */,
  {32'hc0a61442, 32'hc05cd720} /* (3, 14, 17) {real, imag} */,
  {32'h3f9a3aa8, 32'hc08ede8b} /* (3, 14, 16) {real, imag} */,
  {32'hc051c6fb, 32'h40082f9d} /* (3, 14, 15) {real, imag} */,
  {32'hc0e8263f, 32'hbf1b1058} /* (3, 14, 14) {real, imag} */,
  {32'hc0a0b970, 32'h3f58cc18} /* (3, 14, 13) {real, imag} */,
  {32'hc0422938, 32'h3f853dd0} /* (3, 14, 12) {real, imag} */,
  {32'hc042f123, 32'hc0958947} /* (3, 14, 11) {real, imag} */,
  {32'h3fa7e430, 32'hc0936ed8} /* (3, 14, 10) {real, imag} */,
  {32'h41056c8f, 32'hbf993d1c} /* (3, 14, 9) {real, imag} */,
  {32'h4104b348, 32'hc022a5ef} /* (3, 14, 8) {real, imag} */,
  {32'h3fb95fe8, 32'hc03e9c2f} /* (3, 14, 7) {real, imag} */,
  {32'h3feabec0, 32'hc0ecf771} /* (3, 14, 6) {real, imag} */,
  {32'hbfec11b4, 32'hbf681008} /* (3, 14, 5) {real, imag} */,
  {32'h4092e896, 32'h40867bef} /* (3, 14, 4) {real, imag} */,
  {32'h40ba2772, 32'h40c4f3c5} /* (3, 14, 3) {real, imag} */,
  {32'h3eeef560, 32'hc02f9f0b} /* (3, 14, 2) {real, imag} */,
  {32'h40488a7b, 32'hc0ad462a} /* (3, 14, 1) {real, imag} */,
  {32'hc0148504, 32'h3ec63a7c} /* (3, 14, 0) {real, imag} */,
  {32'h3f4e9ba6, 32'h3e4fa9b8} /* (3, 13, 31) {real, imag} */,
  {32'hc00bca6c, 32'hc0494cbe} /* (3, 13, 30) {real, imag} */,
  {32'hc0a9d9f0, 32'hc105a1c0} /* (3, 13, 29) {real, imag} */,
  {32'hc035cc31, 32'hc0759ad2} /* (3, 13, 28) {real, imag} */,
  {32'hbfef34fe, 32'hc050d9da} /* (3, 13, 27) {real, imag} */,
  {32'hbe61c410, 32'h3f7f92bc} /* (3, 13, 26) {real, imag} */,
  {32'h3f3517a8, 32'h4032fe35} /* (3, 13, 25) {real, imag} */,
  {32'hc08cae8d, 32'hbfdd7fb8} /* (3, 13, 24) {real, imag} */,
  {32'h3d001700, 32'h40e7a626} /* (3, 13, 23) {real, imag} */,
  {32'h3f1cd974, 32'h41206496} /* (3, 13, 22) {real, imag} */,
  {32'h3f4ef168, 32'h4080e41a} /* (3, 13, 21) {real, imag} */,
  {32'h3cbb4c00, 32'h40e13b94} /* (3, 13, 20) {real, imag} */,
  {32'hbf4d1fb0, 32'h40a190b6} /* (3, 13, 19) {real, imag} */,
  {32'hc0111eba, 32'h3fd8df44} /* (3, 13, 18) {real, imag} */,
  {32'hc0b329bc, 32'h402606df} /* (3, 13, 17) {real, imag} */,
  {32'h3fbc6628, 32'h403e6c62} /* (3, 13, 16) {real, imag} */,
  {32'h40c99a2a, 32'h40a20a3e} /* (3, 13, 15) {real, imag} */,
  {32'h3fa43ec0, 32'h4006ad7c} /* (3, 13, 14) {real, imag} */,
  {32'hbe90e108, 32'hc0c7e564} /* (3, 13, 13) {real, imag} */,
  {32'hc04746d8, 32'hc10de658} /* (3, 13, 12) {real, imag} */,
  {32'hc122558e, 32'hc06afbd7} /* (3, 13, 11) {real, imag} */,
  {32'hbfe48530, 32'h4099bbf9} /* (3, 13, 10) {real, imag} */,
  {32'h4005f41c, 32'hbf8a6438} /* (3, 13, 9) {real, imag} */,
  {32'h3f30da00, 32'h402e1980} /* (3, 13, 8) {real, imag} */,
  {32'h3fc7f0a8, 32'hbe7ced20} /* (3, 13, 7) {real, imag} */,
  {32'h40944950, 32'hc00941cf} /* (3, 13, 6) {real, imag} */,
  {32'h3f9f9da4, 32'h40a70625} /* (3, 13, 5) {real, imag} */,
  {32'h40b5e42a, 32'h40f78d2f} /* (3, 13, 4) {real, imag} */,
  {32'hc05f8b4b, 32'h40afa8d8} /* (3, 13, 3) {real, imag} */,
  {32'hc0c72b36, 32'h401eb571} /* (3, 13, 2) {real, imag} */,
  {32'hbeaa7270, 32'hc005951a} /* (3, 13, 1) {real, imag} */,
  {32'h3ff12f62, 32'h3f731c20} /* (3, 13, 0) {real, imag} */,
  {32'h3f1612f0, 32'hc0f1d736} /* (3, 12, 31) {real, imag} */,
  {32'h3fd1b39e, 32'hc0d32595} /* (3, 12, 30) {real, imag} */,
  {32'h40c65fab, 32'hbfa1bfcc} /* (3, 12, 29) {real, imag} */,
  {32'hc006bb32, 32'hc067b0ba} /* (3, 12, 28) {real, imag} */,
  {32'hc0cfb836, 32'h4008fb92} /* (3, 12, 27) {real, imag} */,
  {32'hc008612a, 32'h412e9f1c} /* (3, 12, 26) {real, imag} */,
  {32'hc10023ca, 32'h40fa2194} /* (3, 12, 25) {real, imag} */,
  {32'h40316316, 32'h3f8e0068} /* (3, 12, 24) {real, imag} */,
  {32'h3ff3e378, 32'hbfae1222} /* (3, 12, 23) {real, imag} */,
  {32'hc01e3ee6, 32'hc0de411b} /* (3, 12, 22) {real, imag} */,
  {32'hc1250960, 32'h3f9d995c} /* (3, 12, 21) {real, imag} */,
  {32'hc16dac56, 32'hc0cbe714} /* (3, 12, 20) {real, imag} */,
  {32'hc0c2266e, 32'hc0425b86} /* (3, 12, 19) {real, imag} */,
  {32'h40c8471c, 32'h40126ff8} /* (3, 12, 18) {real, imag} */,
  {32'h41008fee, 32'h4109c606} /* (3, 12, 17) {real, imag} */,
  {32'h40e64523, 32'h40708638} /* (3, 12, 16) {real, imag} */,
  {32'h40445888, 32'h3f2dc958} /* (3, 12, 15) {real, imag} */,
  {32'h3fc3d744, 32'hbfbe0bb0} /* (3, 12, 14) {real, imag} */,
  {32'hbf963e3c, 32'hc08729d1} /* (3, 12, 13) {real, imag} */,
  {32'hc012820e, 32'hc058c521} /* (3, 12, 12) {real, imag} */,
  {32'h407dc472, 32'h41258587} /* (3, 12, 11) {real, imag} */,
  {32'h40f45b57, 32'h40e25811} /* (3, 12, 10) {real, imag} */,
  {32'h3fa47342, 32'hbfee70b4} /* (3, 12, 9) {real, imag} */,
  {32'hc0d781c6, 32'hbfa66c74} /* (3, 12, 8) {real, imag} */,
  {32'h3ff3e326, 32'hc00fe6b8} /* (3, 12, 7) {real, imag} */,
  {32'hbc9f0e80, 32'h40214803} /* (3, 12, 6) {real, imag} */,
  {32'h405e4122, 32'hbf0052c8} /* (3, 12, 5) {real, imag} */,
  {32'h4014e6e6, 32'hbf1d733b} /* (3, 12, 4) {real, imag} */,
  {32'h3e134810, 32'h40607f16} /* (3, 12, 3) {real, imag} */,
  {32'h40e12b3c, 32'h402d4552} /* (3, 12, 2) {real, imag} */,
  {32'h3c2dd800, 32'hbf08e380} /* (3, 12, 1) {real, imag} */,
  {32'h3fbe3bdd, 32'hbffb1d86} /* (3, 12, 0) {real, imag} */,
  {32'h3df687c0, 32'hbf40b2c8} /* (3, 11, 31) {real, imag} */,
  {32'h40aaf11d, 32'hc04c91b4} /* (3, 11, 30) {real, imag} */,
  {32'hbfdc7802, 32'h40b749d4} /* (3, 11, 29) {real, imag} */,
  {32'h4106ea10, 32'h409ab5d0} /* (3, 11, 28) {real, imag} */,
  {32'h41040f89, 32'hc0245a5e} /* (3, 11, 27) {real, imag} */,
  {32'h40bebe7a, 32'hbff7ae44} /* (3, 11, 26) {real, imag} */,
  {32'h4149081c, 32'h3ff2bb54} /* (3, 11, 25) {real, imag} */,
  {32'h414dbebf, 32'hbf5a0558} /* (3, 11, 24) {real, imag} */,
  {32'h412d18b2, 32'h407a15dc} /* (3, 11, 23) {real, imag} */,
  {32'h3fefe696, 32'hc0be6d4c} /* (3, 11, 22) {real, imag} */,
  {32'hbf72d3e8, 32'hc12a65af} /* (3, 11, 21) {real, imag} */,
  {32'hc104ce94, 32'h4020dd2f} /* (3, 11, 20) {real, imag} */,
  {32'hc0e89812, 32'h40c146c2} /* (3, 11, 19) {real, imag} */,
  {32'hc047887a, 32'h3fc82128} /* (3, 11, 18) {real, imag} */,
  {32'hc13cef7f, 32'hc10a149d} /* (3, 11, 17) {real, imag} */,
  {32'hc15316f0, 32'hc1045e07} /* (3, 11, 16) {real, imag} */,
  {32'hc11054ee, 32'hbfd4568c} /* (3, 11, 15) {real, imag} */,
  {32'hc10f9d02, 32'h40f87919} /* (3, 11, 14) {real, imag} */,
  {32'hc10644de, 32'h40b092e3} /* (3, 11, 13) {real, imag} */,
  {32'h40344c36, 32'hbfb79bba} /* (3, 11, 12) {real, imag} */,
  {32'hc05d313d, 32'h40a0316a} /* (3, 11, 11) {real, imag} */,
  {32'hc0864eaf, 32'h4016e4fe} /* (3, 11, 10) {real, imag} */,
  {32'h3f3392d0, 32'hc04bf63a} /* (3, 11, 9) {real, imag} */,
  {32'h400f5a6e, 32'hc10885fc} /* (3, 11, 8) {real, imag} */,
  {32'h404bdf72, 32'hc1642397} /* (3, 11, 7) {real, imag} */,
  {32'h4076daf6, 32'hbf98e2b0} /* (3, 11, 6) {real, imag} */,
  {32'h40f74596, 32'h3fac7a24} /* (3, 11, 5) {real, imag} */,
  {32'h40062004, 32'hc12bb0b5} /* (3, 11, 4) {real, imag} */,
  {32'h41802fe2, 32'hbf7c3114} /* (3, 11, 3) {real, imag} */,
  {32'h413b7fc8, 32'h41811511} /* (3, 11, 2) {real, imag} */,
  {32'h3fffa576, 32'h40cdaa30} /* (3, 11, 1) {real, imag} */,
  {32'hbfe1c724, 32'hbfaec763} /* (3, 11, 0) {real, imag} */,
  {32'hc0cf8e07, 32'hc04026ae} /* (3, 10, 31) {real, imag} */,
  {32'hc1390f06, 32'h3ff7ed00} /* (3, 10, 30) {real, imag} */,
  {32'hc11e666c, 32'hc09b7a54} /* (3, 10, 29) {real, imag} */,
  {32'h4000fe23, 32'hc1056402} /* (3, 10, 28) {real, imag} */,
  {32'h3e62fc80, 32'h3fd092fc} /* (3, 10, 27) {real, imag} */,
  {32'hc15b6690, 32'hc0f89492} /* (3, 10, 26) {real, imag} */,
  {32'hc12d022e, 32'hc149d2d0} /* (3, 10, 25) {real, imag} */,
  {32'hc00b1360, 32'h40d58ae9} /* (3, 10, 24) {real, imag} */,
  {32'hc0ebe045, 32'h40278464} /* (3, 10, 23) {real, imag} */,
  {32'hc0004ec4, 32'hc116baa7} /* (3, 10, 22) {real, imag} */,
  {32'h40567dd0, 32'hc1644cdf} /* (3, 10, 21) {real, imag} */,
  {32'h3db99100, 32'hc138eaca} /* (3, 10, 20) {real, imag} */,
  {32'h40a94107, 32'hc044f38a} /* (3, 10, 19) {real, imag} */,
  {32'hc01edd80, 32'h3fc94e04} /* (3, 10, 18) {real, imag} */,
  {32'h4061e806, 32'hc127eae4} /* (3, 10, 17) {real, imag} */,
  {32'h40c95cc8, 32'hc008194a} /* (3, 10, 16) {real, imag} */,
  {32'h3fdd1766, 32'h411980de} /* (3, 10, 15) {real, imag} */,
  {32'h40d63d3b, 32'hc10a5b2e} /* (3, 10, 14) {real, imag} */,
  {32'h40e3fe3f, 32'hc107b940} /* (3, 10, 13) {real, imag} */,
  {32'h40df0218, 32'hc033f724} /* (3, 10, 12) {real, imag} */,
  {32'hc0b38c3c, 32'hc0cac6fe} /* (3, 10, 11) {real, imag} */,
  {32'hc0d03b33, 32'hc1b30e6c} /* (3, 10, 10) {real, imag} */,
  {32'hc0be28c7, 32'hc18aa63e} /* (3, 10, 9) {real, imag} */,
  {32'hc143301b, 32'hc1216592} /* (3, 10, 8) {real, imag} */,
  {32'hc0878703, 32'hc1483d3a} /* (3, 10, 7) {real, imag} */,
  {32'hc0833f33, 32'hc184b7cf} /* (3, 10, 6) {real, imag} */,
  {32'hc17926f7, 32'hc1399390} /* (3, 10, 5) {real, imag} */,
  {32'hc06e6fb4, 32'hc13c09d0} /* (3, 10, 4) {real, imag} */,
  {32'hc0a4a4f0, 32'h40e9ce25} /* (3, 10, 3) {real, imag} */,
  {32'h4064150f, 32'h41135ab0} /* (3, 10, 2) {real, imag} */,
  {32'h4144bfef, 32'hc0cb9238} /* (3, 10, 1) {real, imag} */,
  {32'h4019105b, 32'hc10c2f02} /* (3, 10, 0) {real, imag} */,
  {32'h40719497, 32'hbfda1bec} /* (3, 9, 31) {real, imag} */,
  {32'h40b058d6, 32'h410d2310} /* (3, 9, 30) {real, imag} */,
  {32'h415442ae, 32'h41810b00} /* (3, 9, 29) {real, imag} */,
  {32'h40055502, 32'h40216902} /* (3, 9, 28) {real, imag} */,
  {32'hc048c1aa, 32'hc137caa0} /* (3, 9, 27) {real, imag} */,
  {32'h40e172b7, 32'hc0ae8394} /* (3, 9, 26) {real, imag} */,
  {32'h412e9e0e, 32'h3fa233aa} /* (3, 9, 25) {real, imag} */,
  {32'h418c8d38, 32'h413a8bdb} /* (3, 9, 24) {real, imag} */,
  {32'h41880d37, 32'h411750bc} /* (3, 9, 23) {real, imag} */,
  {32'h41558d6a, 32'hc130a6dc} /* (3, 9, 22) {real, imag} */,
  {32'h413f34f5, 32'hc180d166} /* (3, 9, 21) {real, imag} */,
  {32'h3f884ed0, 32'hc0f1e45c} /* (3, 9, 20) {real, imag} */,
  {32'h40eeca6a, 32'hc11f85a3} /* (3, 9, 19) {real, imag} */,
  {32'h4042ab1a, 32'hc1246fd6} /* (3, 9, 18) {real, imag} */,
  {32'hbe7e7bc0, 32'hc133066d} /* (3, 9, 17) {real, imag} */,
  {32'h4134300d, 32'h3f2fd254} /* (3, 9, 16) {real, imag} */,
  {32'h4134ca9e, 32'hbf8e5a04} /* (3, 9, 15) {real, imag} */,
  {32'h412dc99d, 32'hc00e0503} /* (3, 9, 14) {real, imag} */,
  {32'h4069207e, 32'h4127372e} /* (3, 9, 13) {real, imag} */,
  {32'hc0cfd00a, 32'h413c12bc} /* (3, 9, 12) {real, imag} */,
  {32'hc1869ad4, 32'h40b86794} /* (3, 9, 11) {real, imag} */,
  {32'hc189f23e, 32'h3e2df960} /* (3, 9, 10) {real, imag} */,
  {32'hc16e0a2b, 32'h4015667a} /* (3, 9, 9) {real, imag} */,
  {32'hc15065a0, 32'hc19088c1} /* (3, 9, 8) {real, imag} */,
  {32'hc01071dc, 32'hc15a10cd} /* (3, 9, 7) {real, imag} */,
  {32'hc005a849, 32'h404b53a4} /* (3, 9, 6) {real, imag} */,
  {32'hc03c05e2, 32'hbffaae70} /* (3, 9, 5) {real, imag} */,
  {32'h3fb3ee88, 32'h41583c04} /* (3, 9, 4) {real, imag} */,
  {32'hbf7fd6f8, 32'h40ce00f6} /* (3, 9, 3) {real, imag} */,
  {32'hc11f8fda, 32'hbfe29bbc} /* (3, 9, 2) {real, imag} */,
  {32'hc13fc227, 32'hc0aab7d0} /* (3, 9, 1) {real, imag} */,
  {32'hc0a82066, 32'hc11f73fc} /* (3, 9, 0) {real, imag} */,
  {32'h41052712, 32'h41688b77} /* (3, 8, 31) {real, imag} */,
  {32'h41223358, 32'h3f012d20} /* (3, 8, 30) {real, imag} */,
  {32'h402409fa, 32'hc134fafc} /* (3, 8, 29) {real, imag} */,
  {32'h413239b2, 32'hc17989ed} /* (3, 8, 28) {real, imag} */,
  {32'h41906607, 32'hc069542e} /* (3, 8, 27) {real, imag} */,
  {32'h41353b45, 32'h3fce7b78} /* (3, 8, 26) {real, imag} */,
  {32'h418e4200, 32'hc100e819} /* (3, 8, 25) {real, imag} */,
  {32'hbf811960, 32'hc1a57444} /* (3, 8, 24) {real, imag} */,
  {32'hc0316730, 32'hc14ecc30} /* (3, 8, 23) {real, imag} */,
  {32'h418415e1, 32'h3fb8c524} /* (3, 8, 22) {real, imag} */,
  {32'h411062c3, 32'hc199f8d4} /* (3, 8, 21) {real, imag} */,
  {32'hc1516bd3, 32'hc109f2ca} /* (3, 8, 20) {real, imag} */,
  {32'hbfbdc3fa, 32'h40f4a864} /* (3, 8, 19) {real, imag} */,
  {32'hc044bbe6, 32'h3f4ec4d0} /* (3, 8, 18) {real, imag} */,
  {32'hc0ff7674, 32'h418fd2ec} /* (3, 8, 17) {real, imag} */,
  {32'h4045fbfc, 32'h41f56e1c} /* (3, 8, 16) {real, imag} */,
  {32'h40d296c6, 32'h41195008} /* (3, 8, 15) {real, imag} */,
  {32'hbf67df40, 32'h3e8f5d80} /* (3, 8, 14) {real, imag} */,
  {32'hc0f34cae, 32'hc069d0e1} /* (3, 8, 13) {real, imag} */,
  {32'hc1906b87, 32'hc0f54ec0} /* (3, 8, 12) {real, imag} */,
  {32'hc1569142, 32'hc1434084} /* (3, 8, 11) {real, imag} */,
  {32'hc0eaad24, 32'hc0112faf} /* (3, 8, 10) {real, imag} */,
  {32'hc0f18018, 32'hc06269ae} /* (3, 8, 9) {real, imag} */,
  {32'hc08687ec, 32'hc087f4c1} /* (3, 8, 8) {real, imag} */,
  {32'h403cc018, 32'hbf5eb1e6} /* (3, 8, 7) {real, imag} */,
  {32'h40aad000, 32'hc17aef4f} /* (3, 8, 6) {real, imag} */,
  {32'h4157df49, 32'hc1a42eab} /* (3, 8, 5) {real, imag} */,
  {32'h415fee8a, 32'hc0691aa0} /* (3, 8, 4) {real, imag} */,
  {32'h404d5503, 32'h4089eb4a} /* (3, 8, 3) {real, imag} */,
  {32'h400c99f6, 32'hc0b811ee} /* (3, 8, 2) {real, imag} */,
  {32'h40b15642, 32'hc18ce311} /* (3, 8, 1) {real, imag} */,
  {32'h3fe07764, 32'hc10b63a4} /* (3, 8, 0) {real, imag} */,
  {32'h40ce90e0, 32'h4092b3e7} /* (3, 7, 31) {real, imag} */,
  {32'h40f70c04, 32'h412dc7e9} /* (3, 7, 30) {real, imag} */,
  {32'hc0cb562a, 32'hc0ea439c} /* (3, 7, 29) {real, imag} */,
  {32'h4033b466, 32'hc1788ce7} /* (3, 7, 28) {real, imag} */,
  {32'hc0c2b7fe, 32'h40b75928} /* (3, 7, 27) {real, imag} */,
  {32'hbffecc7e, 32'h3fdf01c8} /* (3, 7, 26) {real, imag} */,
  {32'h40a4fc74, 32'h40a4093a} /* (3, 7, 25) {real, imag} */,
  {32'hc01b8e74, 32'h40964852} /* (3, 7, 24) {real, imag} */,
  {32'h409fdcef, 32'h417ef06f} /* (3, 7, 23) {real, imag} */,
  {32'h408f708f, 32'h4197dbd6} /* (3, 7, 22) {real, imag} */,
  {32'h3fc3b0fc, 32'h4160b5c6} /* (3, 7, 21) {real, imag} */,
  {32'h409c0fd7, 32'h41819aee} /* (3, 7, 20) {real, imag} */,
  {32'h40faa918, 32'hc18780b4} /* (3, 7, 19) {real, imag} */,
  {32'h3f8dd37c, 32'hc148c1a0} /* (3, 7, 18) {real, imag} */,
  {32'h40b406f0, 32'h41189a1d} /* (3, 7, 17) {real, imag} */,
  {32'hc0c57c62, 32'h41288934} /* (3, 7, 16) {real, imag} */,
  {32'hc1081074, 32'h3e8dba70} /* (3, 7, 15) {real, imag} */,
  {32'hc153606a, 32'h40ecae34} /* (3, 7, 14) {real, imag} */,
  {32'h4143f782, 32'h40ba8f87} /* (3, 7, 13) {real, imag} */,
  {32'h40f4991c, 32'hbfb248e4} /* (3, 7, 12) {real, imag} */,
  {32'hc098c8e2, 32'hc0a6ac2f} /* (3, 7, 11) {real, imag} */,
  {32'h40619a82, 32'hbf983362} /* (3, 7, 10) {real, imag} */,
  {32'hc14a32e1, 32'h4081d304} /* (3, 7, 9) {real, imag} */,
  {32'hc12aab3a, 32'h400a2870} /* (3, 7, 8) {real, imag} */,
  {32'hc0dd206c, 32'h41744a23} /* (3, 7, 7) {real, imag} */,
  {32'h40665527, 32'h411a6ae1} /* (3, 7, 6) {real, imag} */,
  {32'h408ca149, 32'hc04b5c84} /* (3, 7, 5) {real, imag} */,
  {32'hc0c32e7a, 32'hbfb602cc} /* (3, 7, 4) {real, imag} */,
  {32'hc0507dc2, 32'hc0a94546} /* (3, 7, 3) {real, imag} */,
  {32'h408a5d90, 32'hc019f0e0} /* (3, 7, 2) {real, imag} */,
  {32'h40c97762, 32'h412d5c1a} /* (3, 7, 1) {real, imag} */,
  {32'h412e9ff3, 32'h4185807a} /* (3, 7, 0) {real, imag} */,
  {32'h40174fc8, 32'h4032dd62} /* (3, 6, 31) {real, imag} */,
  {32'h4124b6ac, 32'hc1893bb6} /* (3, 6, 30) {real, imag} */,
  {32'h40d68a2d, 32'hc10121e2} /* (3, 6, 29) {real, imag} */,
  {32'hc17ee366, 32'hc107d362} /* (3, 6, 28) {real, imag} */,
  {32'hc1a0ed03, 32'hbf293308} /* (3, 6, 27) {real, imag} */,
  {32'hbd991560, 32'h412ad5f7} /* (3, 6, 26) {real, imag} */,
  {32'h3fcd2a96, 32'h40ff3294} /* (3, 6, 25) {real, imag} */,
  {32'hc11aa1dc, 32'h40aa4801} /* (3, 6, 24) {real, imag} */,
  {32'hc09e44bd, 32'h40ffca0a} /* (3, 6, 23) {real, imag} */,
  {32'h410eeb76, 32'h4151f62e} /* (3, 6, 22) {real, imag} */,
  {32'h412c1e96, 32'h41b7be68} /* (3, 6, 21) {real, imag} */,
  {32'hbf2419b8, 32'hc1119d0c} /* (3, 6, 20) {real, imag} */,
  {32'hbf0dc558, 32'hc179ddde} /* (3, 6, 19) {real, imag} */,
  {32'h4081192c, 32'h40fe0a5f} /* (3, 6, 18) {real, imag} */,
  {32'h414b663e, 32'h41166b8c} /* (3, 6, 17) {real, imag} */,
  {32'h41400e96, 32'hc053e05e} /* (3, 6, 16) {real, imag} */,
  {32'h40b29b16, 32'h4101c3e1} /* (3, 6, 15) {real, imag} */,
  {32'hc1935a52, 32'h4186306a} /* (3, 6, 14) {real, imag} */,
  {32'h4054468a, 32'hc09be11a} /* (3, 6, 13) {real, imag} */,
  {32'h41d8e782, 32'h40d03c3a} /* (3, 6, 12) {real, imag} */,
  {32'h41330c46, 32'h414edf35} /* (3, 6, 11) {real, imag} */,
  {32'hc148cb46, 32'h41b9e18c} /* (3, 6, 10) {real, imag} */,
  {32'hc1384e3a, 32'h4120ba89} /* (3, 6, 9) {real, imag} */,
  {32'h40d2bd90, 32'h40ba0dc4} /* (3, 6, 8) {real, imag} */,
  {32'h40da2686, 32'h401fcee0} /* (3, 6, 7) {real, imag} */,
  {32'hc08a27e0, 32'hc0ce98d4} /* (3, 6, 6) {real, imag} */,
  {32'h405fe6ce, 32'h41a848db} /* (3, 6, 5) {real, imag} */,
  {32'h40226e1c, 32'h414f9d6f} /* (3, 6, 4) {real, imag} */,
  {32'h40e6c070, 32'h3f96914c} /* (3, 6, 3) {real, imag} */,
  {32'h40cd5495, 32'hc13d91a3} /* (3, 6, 2) {real, imag} */,
  {32'h40007d34, 32'hc1c84fe4} /* (3, 6, 1) {real, imag} */,
  {32'hc110bf59, 32'hc1285a2c} /* (3, 6, 0) {real, imag} */,
  {32'h41686846, 32'hc1a3cf3e} /* (3, 5, 31) {real, imag} */,
  {32'h41075b2c, 32'hc1a9f41a} /* (3, 5, 30) {real, imag} */,
  {32'h4194ad1b, 32'hc174f1ea} /* (3, 5, 29) {real, imag} */,
  {32'h41df692c, 32'hc1afec96} /* (3, 5, 28) {real, imag} */,
  {32'h421258ca, 32'hc222c786} /* (3, 5, 27) {real, imag} */,
  {32'h4199008a, 32'hc22e4390} /* (3, 5, 26) {real, imag} */,
  {32'h412907fa, 32'hc220378e} /* (3, 5, 25) {real, imag} */,
  {32'h41d57090, 32'hc1b3b8cb} /* (3, 5, 24) {real, imag} */,
  {32'h40d03199, 32'hc198bc10} /* (3, 5, 23) {real, imag} */,
  {32'h4143c512, 32'hc17d5ef2} /* (3, 5, 22) {real, imag} */,
  {32'h41b2ada4, 32'hc177c8b3} /* (3, 5, 21) {real, imag} */,
  {32'hc03e4a3a, 32'h40d2de54} /* (3, 5, 20) {real, imag} */,
  {32'hc19d1d26, 32'h41e70520} /* (3, 5, 19) {real, imag} */,
  {32'hc1980f02, 32'h41970d7d} /* (3, 5, 18) {real, imag} */,
  {32'hc1a6f617, 32'h410c2790} /* (3, 5, 17) {real, imag} */,
  {32'hc1779e5a, 32'h41b31cb8} /* (3, 5, 16) {real, imag} */,
  {32'h41446a31, 32'h41a66eba} /* (3, 5, 15) {real, imag} */,
  {32'hc10cdf1c, 32'h418bd64a} /* (3, 5, 14) {real, imag} */,
  {32'hc1b9617e, 32'h40f4070c} /* (3, 5, 13) {real, imag} */,
  {32'hc1cb9bff, 32'h41915890} /* (3, 5, 12) {real, imag} */,
  {32'hc1cc18d9, 32'h41c6a34d} /* (3, 5, 11) {real, imag} */,
  {32'hc1265dde, 32'h40e35b46} /* (3, 5, 10) {real, imag} */,
  {32'hc0f0fa1a, 32'hc1aed73c} /* (3, 5, 9) {real, imag} */,
  {32'h41121e42, 32'hc1c20e17} /* (3, 5, 8) {real, imag} */,
  {32'h4098bf57, 32'hc0f96a80} /* (3, 5, 7) {real, imag} */,
  {32'hc11da98d, 32'h3ffadfb8} /* (3, 5, 6) {real, imag} */,
  {32'h3ebe78c0, 32'hc169b676} /* (3, 5, 5) {real, imag} */,
  {32'h418805d2, 32'hc1aa0e64} /* (3, 5, 4) {real, imag} */,
  {32'h422ed4ce, 32'hc1d5929d} /* (3, 5, 3) {real, imag} */,
  {32'h41bd1296, 32'hc10afdf3} /* (3, 5, 2) {real, imag} */,
  {32'h40d51b91, 32'hc1752900} /* (3, 5, 1) {real, imag} */,
  {32'h41276e2e, 32'hc0e37c8c} /* (3, 5, 0) {real, imag} */,
  {32'h401321d9, 32'h4107a78d} /* (3, 4, 31) {real, imag} */,
  {32'hbfd41e28, 32'h41959810} /* (3, 4, 30) {real, imag} */,
  {32'hc184c9de, 32'h41aa0498} /* (3, 4, 29) {real, imag} */,
  {32'hc0da2360, 32'h410601a1} /* (3, 4, 28) {real, imag} */,
  {32'hc179ad0c, 32'h410eefa6} /* (3, 4, 27) {real, imag} */,
  {32'hc19a5ab6, 32'h41a73204} /* (3, 4, 26) {real, imag} */,
  {32'hc139c6d6, 32'h41ac8d9e} /* (3, 4, 25) {real, imag} */,
  {32'hc1264026, 32'h41ea320a} /* (3, 4, 24) {real, imag} */,
  {32'hc1b0c792, 32'h421426d6} /* (3, 4, 23) {real, imag} */,
  {32'hc18ea860, 32'h4217a1fe} /* (3, 4, 22) {real, imag} */,
  {32'h403e6370, 32'h412d6f3b} /* (3, 4, 21) {real, imag} */,
  {32'h41d1c521, 32'hc18f80f6} /* (3, 4, 20) {real, imag} */,
  {32'h41c0e0e9, 32'hc1aaf725} /* (3, 4, 19) {real, imag} */,
  {32'h41eaa807, 32'hc1bbbe3c} /* (3, 4, 18) {real, imag} */,
  {32'h41e41264, 32'hc1a8fba3} /* (3, 4, 17) {real, imag} */,
  {32'h414da16f, 32'h4035c330} /* (3, 4, 16) {real, imag} */,
  {32'h4197d451, 32'h41467199} /* (3, 4, 15) {real, imag} */,
  {32'h422759ea, 32'hbf841a60} /* (3, 4, 14) {real, imag} */,
  {32'h4200d4b8, 32'hc06f43a8} /* (3, 4, 13) {real, imag} */,
  {32'h4158173b, 32'hc0ca6f94} /* (3, 4, 12) {real, imag} */,
  {32'h4109b47a, 32'hc169b6f6} /* (3, 4, 11) {real, imag} */,
  {32'hc1b8356c, 32'h4141136e} /* (3, 4, 10) {real, imag} */,
  {32'hc1b1775d, 32'h41b2dc60} /* (3, 4, 9) {real, imag} */,
  {32'hc1efe455, 32'h41e10d93} /* (3, 4, 8) {real, imag} */,
  {32'hc23368f3, 32'h41ff77c8} /* (3, 4, 7) {real, imag} */,
  {32'hc2232411, 32'h4201d3ba} /* (3, 4, 6) {real, imag} */,
  {32'hbfc1a510, 32'h41c43c0c} /* (3, 4, 5) {real, imag} */,
  {32'h3f197764, 32'h41a2c03a} /* (3, 4, 4) {real, imag} */,
  {32'hc127d79e, 32'h41fbc8e6} /* (3, 4, 3) {real, imag} */,
  {32'hc1ad9433, 32'h41f06e4f} /* (3, 4, 2) {real, imag} */,
  {32'hc1433e18, 32'h41e70ab9} /* (3, 4, 1) {real, imag} */,
  {32'h41387747, 32'h4107c674} /* (3, 4, 0) {real, imag} */,
  {32'h40c0f65c, 32'h3ec0f5a0} /* (3, 3, 31) {real, imag} */,
  {32'hbff2c0a0, 32'h408ce909} /* (3, 3, 30) {real, imag} */,
  {32'hc1247e5d, 32'hc137d295} /* (3, 3, 29) {real, imag} */,
  {32'h411ed09e, 32'hc1cfc2f0} /* (3, 3, 28) {real, imag} */,
  {32'h41208bb1, 32'hc0a00c58} /* (3, 3, 27) {real, imag} */,
  {32'h41a8da49, 32'hc1bbbad0} /* (3, 3, 26) {real, imag} */,
  {32'hc02211ca, 32'hc18c8d72} /* (3, 3, 25) {real, imag} */,
  {32'hc04bb6be, 32'hc1b41b44} /* (3, 3, 24) {real, imag} */,
  {32'hc14bc5a0, 32'hc0e74c1c} /* (3, 3, 23) {real, imag} */,
  {32'hc169cd1f, 32'hc15ec34d} /* (3, 3, 22) {real, imag} */,
  {32'h4147ee0a, 32'h412a1f14} /* (3, 3, 21) {real, imag} */,
  {32'h41cd4255, 32'h4204c688} /* (3, 3, 20) {real, imag} */,
  {32'h41c34176, 32'h41b4e839} /* (3, 3, 19) {real, imag} */,
  {32'h41419110, 32'h40d896da} /* (3, 3, 18) {real, imag} */,
  {32'h4199d683, 32'h40d424cb} /* (3, 3, 17) {real, imag} */,
  {32'h4240ca16, 32'h41025c49} /* (3, 3, 16) {real, imag} */,
  {32'hc113848e, 32'h40ba93f6} /* (3, 3, 15) {real, imag} */,
  {32'hc20f258b, 32'hc171bb11} /* (3, 3, 14) {real, imag} */,
  {32'hc149aed2, 32'hc04da368} /* (3, 3, 13) {real, imag} */,
  {32'h41bcc4c4, 32'h411a3c45} /* (3, 3, 12) {real, imag} */,
  {32'h415b0342, 32'h41998e3c} /* (3, 3, 11) {real, imag} */,
  {32'hc1828e7b, 32'hc190e180} /* (3, 3, 10) {real, imag} */,
  {32'hc136f8f8, 32'hc257b8fb} /* (3, 3, 9) {real, imag} */,
  {32'hc19a1d82, 32'hc1a910b0} /* (3, 3, 8) {real, imag} */,
  {32'hc21af24e, 32'hc191bdf1} /* (3, 3, 7) {real, imag} */,
  {32'hc1d14ac9, 32'hc177cb51} /* (3, 3, 6) {real, imag} */,
  {32'hc0090c00, 32'hc1a45ace} /* (3, 3, 5) {real, imag} */,
  {32'hc1101dfe, 32'hc09d2119} /* (3, 3, 4) {real, imag} */,
  {32'hc1398869, 32'h4145249c} /* (3, 3, 3) {real, imag} */,
  {32'hc130a42a, 32'hc14822a1} /* (3, 3, 2) {real, imag} */,
  {32'hc1af7efc, 32'hc1875c3a} /* (3, 3, 1) {real, imag} */,
  {32'h3f5e48c8, 32'hc0304c7c} /* (3, 3, 0) {real, imag} */,
  {32'h40e5466b, 32'hc21f15a9} /* (3, 2, 31) {real, imag} */,
  {32'h41a0dd1e, 32'hc247cc10} /* (3, 2, 30) {real, imag} */,
  {32'h41cd2eed, 32'hc25258f3} /* (3, 2, 29) {real, imag} */,
  {32'h42040ac9, 32'hc244a1ef} /* (3, 2, 28) {real, imag} */,
  {32'h42274d58, 32'hc21cbd72} /* (3, 2, 27) {real, imag} */,
  {32'h41ed5d87, 32'hc215842e} /* (3, 2, 26) {real, imag} */,
  {32'h41e9126e, 32'hc214a372} /* (3, 2, 25) {real, imag} */,
  {32'h42013942, 32'hc2063a46} /* (3, 2, 24) {real, imag} */,
  {32'h41ef9988, 32'hc25fb53c} /* (3, 2, 23) {real, imag} */,
  {32'h41fd038b, 32'hc221ba70} /* (3, 2, 22) {real, imag} */,
  {32'h41a4b18e, 32'hc0e880b4} /* (3, 2, 21) {real, imag} */,
  {32'h41ea86df, 32'h428de2d3} /* (3, 2, 20) {real, imag} */,
  {32'h416943d4, 32'h42bdcf4e} /* (3, 2, 19) {real, imag} */,
  {32'h40291f90, 32'h42c1b0ca} /* (3, 2, 18) {real, imag} */,
  {32'h411138be, 32'h42d9b40f} /* (3, 2, 17) {real, imag} */,
  {32'hc109ec03, 32'h42a806dd} /* (3, 2, 16) {real, imag} */,
  {32'hc1e2921a, 32'h425c9d64} /* (3, 2, 15) {real, imag} */,
  {32'hc192119c, 32'h42824f0a} /* (3, 2, 14) {real, imag} */,
  {32'hc1c10ec0, 32'h4211fa36} /* (3, 2, 13) {real, imag} */,
  {32'hc1becdca, 32'h41c3e797} /* (3, 2, 12) {real, imag} */,
  {32'hc1bda720, 32'h415b9a66} /* (3, 2, 11) {real, imag} */,
  {32'hc1cfcad4, 32'hc2168416} /* (3, 2, 10) {real, imag} */,
  {32'hc0cd4790, 32'hc2aa1867} /* (3, 2, 9) {real, imag} */,
  {32'hc027dd00, 32'hc299d16f} /* (3, 2, 8) {real, imag} */,
  {32'hc1637934, 32'hc2938c60} /* (3, 2, 7) {real, imag} */,
  {32'h40a935f8, 32'hc2a3d57b} /* (3, 2, 6) {real, imag} */,
  {32'h41efadbb, 32'hc2801d1f} /* (3, 2, 5) {real, imag} */,
  {32'h40e04056, 32'hc2433320} /* (3, 2, 4) {real, imag} */,
  {32'h40b2eb38, 32'hc26bef84} /* (3, 2, 3) {real, imag} */,
  {32'h418a5201, 32'hc257c6b1} /* (3, 2, 2) {real, imag} */,
  {32'h41f5ab50, 32'hc204ed19} /* (3, 2, 1) {real, imag} */,
  {32'h419b81c6, 32'hc1f475a6} /* (3, 2, 0) {real, imag} */,
  {32'hc1858fea, 32'h426d7393} /* (3, 1, 31) {real, imag} */,
  {32'hc1fe9c60, 32'h42c9b9aa} /* (3, 1, 30) {real, imag} */,
  {32'hc1a7df75, 32'h42a6d148} /* (3, 1, 29) {real, imag} */,
  {32'hc1fbd204, 32'h428eb754} /* (3, 1, 28) {real, imag} */,
  {32'hc263e570, 32'h42a5da49} /* (3, 1, 27) {real, imag} */,
  {32'hc250ffc4, 32'h42c6660d} /* (3, 1, 26) {real, imag} */,
  {32'hc27803c8, 32'h42e7d2a4} /* (3, 1, 25) {real, imag} */,
  {32'hc2230b40, 32'h42d9a8e9} /* (3, 1, 24) {real, imag} */,
  {32'hc1f10685, 32'h42990b4b} /* (3, 1, 23) {real, imag} */,
  {32'hc22ce712, 32'h42a8f8ca} /* (3, 1, 22) {real, imag} */,
  {32'hc09917e5, 32'h4227c80d} /* (3, 1, 21) {real, imag} */,
  {32'h427971d8, 32'hc2381e80} /* (3, 1, 20) {real, imag} */,
  {32'h429366bc, 32'hc238c4a2} /* (3, 1, 19) {real, imag} */,
  {32'h429c5416, 32'hc1ecc052} /* (3, 1, 18) {real, imag} */,
  {32'h4240bf38, 32'hc206dc9f} /* (3, 1, 17) {real, imag} */,
  {32'h41c61e88, 32'hc1f356ad} /* (3, 1, 16) {real, imag} */,
  {32'h41b27e12, 32'hc295273e} /* (3, 1, 15) {real, imag} */,
  {32'h423cd3b8, 32'hc2a3133b} /* (3, 1, 14) {real, imag} */,
  {32'h41c53241, 32'hc2c3af23} /* (3, 1, 13) {real, imag} */,
  {32'h409ce44a, 32'hc2a18535} /* (3, 1, 12) {real, imag} */,
  {32'h41a00da9, 32'hc28628e0} /* (3, 1, 11) {real, imag} */,
  {32'hc1906d58, 32'hc12cea9a} /* (3, 1, 10) {real, imag} */,
  {32'hc2404ab3, 32'h4217e1a6} /* (3, 1, 9) {real, imag} */,
  {32'hc21e3be5, 32'h4211abf4} /* (3, 1, 8) {real, imag} */,
  {32'hc2212910, 32'h419667ee} /* (3, 1, 7) {real, imag} */,
  {32'hc20bf3fd, 32'h4171406e} /* (3, 1, 6) {real, imag} */,
  {32'hc27394a2, 32'h4262039c} /* (3, 1, 5) {real, imag} */,
  {32'hc207620e, 32'h42b7d3ae} /* (3, 1, 4) {real, imag} */,
  {32'hc21c5808, 32'h42eb421c} /* (3, 1, 3) {real, imag} */,
  {32'hc23c1f25, 32'h42e0d402} /* (3, 1, 2) {real, imag} */,
  {32'hc18923c2, 32'h42b41fa1} /* (3, 1, 1) {real, imag} */,
  {32'hc100d2b1, 32'h4248c567} /* (3, 1, 0) {real, imag} */,
  {32'hc1d7bcb8, 32'h4140dd72} /* (3, 0, 31) {real, imag} */,
  {32'hc1da627f, 32'h41fd60d0} /* (3, 0, 30) {real, imag} */,
  {32'h415470fa, 32'h4283f754} /* (3, 0, 29) {real, imag} */,
  {32'hc189cf68, 32'h425ca8f6} /* (3, 0, 28) {real, imag} */,
  {32'hc1935af2, 32'h42894d24} /* (3, 0, 27) {real, imag} */,
  {32'h4103887b, 32'h429f7944} /* (3, 0, 26) {real, imag} */,
  {32'h420beac4, 32'h42826d1e} /* (3, 0, 25) {real, imag} */,
  {32'hbfdd9c13, 32'h42179f55} /* (3, 0, 24) {real, imag} */,
  {32'hc1ba9dc7, 32'h420e52c3} /* (3, 0, 23) {real, imag} */,
  {32'hc21c6dc0, 32'h421a4c1c} /* (3, 0, 22) {real, imag} */,
  {32'hc23eb860, 32'h423bc64f} /* (3, 0, 21) {real, imag} */,
  {32'hc06216a6, 32'h410707da} /* (3, 0, 20) {real, imag} */,
  {32'h4130e6fd, 32'hc12da657} /* (3, 0, 19) {real, imag} */,
  {32'hc10f65e1, 32'hc087a9a0} /* (3, 0, 18) {real, imag} */,
  {32'hc1c738b2, 32'h40dc9774} /* (3, 0, 17) {real, imag} */,
  {32'hc14b2c47, 32'hbf92b94a} /* (3, 0, 16) {real, imag} */,
  {32'h407da895, 32'hc22f9456} /* (3, 0, 15) {real, imag} */,
  {32'h41f502d8, 32'hc28b422b} /* (3, 0, 14) {real, imag} */,
  {32'h4193c400, 32'hc259683b} /* (3, 0, 13) {real, imag} */,
  {32'h40f7b353, 32'hc282b239} /* (3, 0, 12) {real, imag} */,
  {32'hc0f26932, 32'hc27e2a21} /* (3, 0, 11) {real, imag} */,
  {32'hc1cfc3a8, 32'hc13db1b8} /* (3, 0, 10) {real, imag} */,
  {32'hc10ca8ac, 32'hc015a57c} /* (3, 0, 9) {real, imag} */,
  {32'hc1513273, 32'hc06452cb} /* (3, 0, 8) {real, imag} */,
  {32'h3f934169, 32'hc0b37ce2} /* (3, 0, 7) {real, imag} */,
  {32'h413d23d8, 32'hc1d65bbe} /* (3, 0, 6) {real, imag} */,
  {32'hc06ff0ce, 32'h41865533} /* (3, 0, 5) {real, imag} */,
  {32'hbe1250a0, 32'h42619f80} /* (3, 0, 4) {real, imag} */,
  {32'hc178637a, 32'h42945984} /* (3, 0, 3) {real, imag} */,
  {32'hc0ff3f07, 32'h42665c6e} /* (3, 0, 2) {real, imag} */,
  {32'hc1318306, 32'h420d76db} /* (3, 0, 1) {real, imag} */,
  {32'hc189b514, 32'h41ca3030} /* (3, 0, 0) {real, imag} */,
  {32'hc18dc3a3, 32'h42fd79ed} /* (2, 31, 31) {real, imag} */,
  {32'hc1afe036, 32'h4368fe95} /* (2, 31, 30) {real, imag} */,
  {32'hc21de24e, 32'h43758503} /* (2, 31, 29) {real, imag} */,
  {32'hc1cd0438, 32'h4383130a} /* (2, 31, 28) {real, imag} */,
  {32'hc186e05e, 32'h437cb755} /* (2, 31, 27) {real, imag} */,
  {32'hc178487b, 32'h43684d5a} /* (2, 31, 26) {real, imag} */,
  {32'hc20bbb62, 32'h436e8b28} /* (2, 31, 25) {real, imag} */,
  {32'hc2332127, 32'h437b1337} /* (2, 31, 24) {real, imag} */,
  {32'hc110d5c0, 32'h43758636} /* (2, 31, 23) {real, imag} */,
  {32'hc1189e34, 32'h4360bbc7} /* (2, 31, 22) {real, imag} */,
  {32'hc22e6fd8, 32'h42f9075a} /* (2, 31, 21) {real, imag} */,
  {32'hc2a373d8, 32'hc2b90b54} /* (2, 31, 20) {real, imag} */,
  {32'hc2db814f, 32'hc30436f8} /* (2, 31, 19) {real, imag} */,
  {32'hc2dfbe5a, 32'hc2d3b782} /* (2, 31, 18) {real, imag} */,
  {32'hc2b46180, 32'hc2e076bc} /* (2, 31, 17) {real, imag} */,
  {32'hc21eb0a3, 32'hc308fdad} /* (2, 31, 16) {real, imag} */,
  {32'h41ea3934, 32'hc356f50f} /* (2, 31, 15) {real, imag} */,
  {32'h41e45cb6, 32'hc365db49} /* (2, 31, 14) {real, imag} */,
  {32'h41a3ae80, 32'hc3702677} /* (2, 31, 13) {real, imag} */,
  {32'h41ec25de, 32'hc36ea5ac} /* (2, 31, 12) {real, imag} */,
  {32'h420926f2, 32'hc343ed39} /* (2, 31, 11) {real, imag} */,
  {32'h4243e4f2, 32'h410e892c} /* (2, 31, 10) {real, imag} */,
  {32'h429fb3f5, 32'h42f32066} /* (2, 31, 9) {real, imag} */,
  {32'h42bf5452, 32'h43004c2e} /* (2, 31, 8) {real, imag} */,
  {32'h42a1c653, 32'h42f5f36b} /* (2, 31, 7) {real, imag} */,
  {32'h42942e28, 32'h43047961} /* (2, 31, 6) {real, imag} */,
  {32'hbf142aa0, 32'h4342a6e0} /* (2, 31, 5) {real, imag} */,
  {32'hc262abb6, 32'h4365e5f9} /* (2, 31, 4) {real, imag} */,
  {32'hc2523be1, 32'h43703d22} /* (2, 31, 3) {real, imag} */,
  {32'hc239e167, 32'h437cefe8} /* (2, 31, 2) {real, imag} */,
  {32'hc1c55872, 32'h43675002} /* (2, 31, 1) {real, imag} */,
  {32'hc008b730, 32'h42f71240} /* (2, 31, 0) {real, imag} */,
  {32'h411482b8, 32'hc28977e1} /* (2, 30, 31) {real, imag} */,
  {32'h40eb1dfc, 32'hc30cffec} /* (2, 30, 30) {real, imag} */,
  {32'hc1db3976, 32'hc3246107} /* (2, 30, 29) {real, imag} */,
  {32'hc0bc5fdc, 32'hc311106a} /* (2, 30, 28) {real, imag} */,
  {32'h41c0b7c0, 32'hc31fc4b2} /* (2, 30, 27) {real, imag} */,
  {32'h41e96f10, 32'hc327a7b4} /* (2, 30, 26) {real, imag} */,
  {32'h4216b22a, 32'hc31ff714} /* (2, 30, 25) {real, imag} */,
  {32'h41d67b75, 32'hc3048cd4} /* (2, 30, 24) {real, imag} */,
  {32'h41859c5e, 32'hc2f4da3c} /* (2, 30, 23) {real, imag} */,
  {32'h40418a80, 32'hc31692f1} /* (2, 30, 22) {real, imag} */,
  {32'hc2453f1e, 32'hc2b665e1} /* (2, 30, 21) {real, imag} */,
  {32'hc2e34cdd, 32'h430a972a} /* (2, 30, 20) {real, imag} */,
  {32'hc2e23ff5, 32'h4339a2f8} /* (2, 30, 19) {real, imag} */,
  {32'hc2efae82, 32'h433e660c} /* (2, 30, 18) {real, imag} */,
  {32'hc301d72c, 32'h432faa66} /* (2, 30, 17) {real, imag} */,
  {32'hc2db0be6, 32'h433006d9} /* (2, 30, 16) {real, imag} */,
  {32'hc264218a, 32'h431cc271} /* (2, 30, 15) {real, imag} */,
  {32'hc0465868, 32'h43042d65} /* (2, 30, 14) {real, imag} */,
  {32'hbf3e9a60, 32'h42dc97e7} /* (2, 30, 13) {real, imag} */,
  {32'hc181c705, 32'h430eca68} /* (2, 30, 12) {real, imag} */,
  {32'h41374892, 32'h42f729c0} /* (2, 30, 11) {real, imag} */,
  {32'h42be94ec, 32'hc2af8085} /* (2, 30, 10) {real, imag} */,
  {32'h431529be, 32'hc3470e7d} /* (2, 30, 9) {real, imag} */,
  {32'h42fd2959, 32'hc3468a9e} /* (2, 30, 8) {real, imag} */,
  {32'h42d0badc, 32'hc33b7f8b} /* (2, 30, 7) {real, imag} */,
  {32'h42cc641c, 32'hc344594e} /* (2, 30, 6) {real, imag} */,
  {32'h4257aa1e, 32'hc31b5db9} /* (2, 30, 5) {real, imag} */,
  {32'h413f7863, 32'hc2e8ab0c} /* (2, 30, 4) {real, imag} */,
  {32'hc17cd3c0, 32'hc30aeba2} /* (2, 30, 3) {real, imag} */,
  {32'h4100cf24, 32'hc3150710} /* (2, 30, 2) {real, imag} */,
  {32'hc10aee54, 32'hc31ef445} /* (2, 30, 1) {real, imag} */,
  {32'hbea11000, 32'hc2afa563} /* (2, 30, 0) {real, imag} */,
  {32'h4152e584, 32'h412c8846} /* (2, 29, 31) {real, imag} */,
  {32'hc08f3612, 32'h4076ba22} /* (2, 29, 30) {real, imag} */,
  {32'hc079c8b6, 32'h40b8c4a6} /* (2, 29, 29) {real, imag} */,
  {32'hc19e3b4e, 32'h41001367} /* (2, 29, 28) {real, imag} */,
  {32'hc20715ac, 32'h40397ef0} /* (2, 29, 27) {real, imag} */,
  {32'hbf804358, 32'hc0361e86} /* (2, 29, 26) {real, imag} */,
  {32'hbecf4e40, 32'hc21ebf28} /* (2, 29, 25) {real, imag} */,
  {32'hc10d0a5f, 32'hc1ffeac2} /* (2, 29, 24) {real, imag} */,
  {32'hc0b751f8, 32'h4117f354} /* (2, 29, 23) {real, imag} */,
  {32'h402e862b, 32'h410fb328} /* (2, 29, 22) {real, imag} */,
  {32'hc1cff6d9, 32'hc05a3a0c} /* (2, 29, 21) {real, imag} */,
  {32'hc296d72c, 32'hbfb8797e} /* (2, 29, 20) {real, imag} */,
  {32'hc2c70049, 32'hc0eadec8} /* (2, 29, 19) {real, imag} */,
  {32'hc2cb0f24, 32'hc151bd80} /* (2, 29, 18) {real, imag} */,
  {32'hc2c16c22, 32'h40360be0} /* (2, 29, 17) {real, imag} */,
  {32'hc29e7aa6, 32'hc14096de} /* (2, 29, 16) {real, imag} */,
  {32'hc21680a3, 32'hc0b20b3b} /* (2, 29, 15) {real, imag} */,
  {32'hc180134e, 32'hc089c726} /* (2, 29, 14) {real, imag} */,
  {32'h411e4e5a, 32'hc15f10c8} /* (2, 29, 13) {real, imag} */,
  {32'hc0de3792, 32'h3e604d40} /* (2, 29, 12) {real, imag} */,
  {32'h416df54c, 32'h41132662} /* (2, 29, 11) {real, imag} */,
  {32'h4261c97a, 32'h411803e0} /* (2, 29, 10) {real, imag} */,
  {32'h42b2ec5d, 32'h4150f750} /* (2, 29, 9) {real, imag} */,
  {32'h4293a825, 32'h40e6d824} /* (2, 29, 8) {real, imag} */,
  {32'h429d0c49, 32'h416e4b75} /* (2, 29, 7) {real, imag} */,
  {32'h42cbc13f, 32'hc05f0150} /* (2, 29, 6) {real, imag} */,
  {32'h4254774a, 32'hc0cb7b60} /* (2, 29, 5) {real, imag} */,
  {32'h41ae2e98, 32'h41a1b901} /* (2, 29, 4) {real, imag} */,
  {32'hc13056a5, 32'h40b4dde9} /* (2, 29, 3) {real, imag} */,
  {32'hc1c1a732, 32'hbfb46ef4} /* (2, 29, 2) {real, imag} */,
  {32'h4158a7f0, 32'hc0950484} /* (2, 29, 1) {real, imag} */,
  {32'h413be48d, 32'h4093f58e} /* (2, 29, 0) {real, imag} */,
  {32'h3ff53eee, 32'h418915d2} /* (2, 28, 31) {real, imag} */,
  {32'h3f86fc14, 32'h419d06ad} /* (2, 28, 30) {real, imag} */,
  {32'h400f0d6e, 32'h4205c36c} /* (2, 28, 29) {real, imag} */,
  {32'h411e88fb, 32'h427826d4} /* (2, 28, 28) {real, imag} */,
  {32'h416466fa, 32'h4285a008} /* (2, 28, 27) {real, imag} */,
  {32'h413d86c3, 32'h42413c0f} /* (2, 28, 26) {real, imag} */,
  {32'hc0d931bc, 32'h41fc6452} /* (2, 28, 25) {real, imag} */,
  {32'h3efb74f0, 32'h4239e3ad} /* (2, 28, 24) {real, imag} */,
  {32'h4173f118, 32'h41d5caa8} /* (2, 28, 23) {real, imag} */,
  {32'h40ca7520, 32'h4215fa30} /* (2, 28, 22) {real, imag} */,
  {32'hc0bdb5fc, 32'h419a11b6} /* (2, 28, 21) {real, imag} */,
  {32'hc2344772, 32'hc28a08eb} /* (2, 28, 20) {real, imag} */,
  {32'hc2809db4, 32'hc2951a52} /* (2, 28, 19) {real, imag} */,
  {32'hc2a862fb, 32'hc2901167} /* (2, 28, 18) {real, imag} */,
  {32'hc291e856, 32'hc2a02079} /* (2, 28, 17) {real, imag} */,
  {32'hc2574e6e, 32'hc29e7224} /* (2, 28, 16) {real, imag} */,
  {32'hc12d19bc, 32'hc28bec75} /* (2, 28, 15) {real, imag} */,
  {32'hc1ba9ea6, 32'hc2800b2e} /* (2, 28, 14) {real, imag} */,
  {32'hc1adf271, 32'hc22141f8} /* (2, 28, 13) {real, imag} */,
  {32'hc0876a75, 32'hc20feb74} /* (2, 28, 12) {real, imag} */,
  {32'hbf09ba38, 32'hc1a3e2a2} /* (2, 28, 11) {real, imag} */,
  {32'h4245fd28, 32'h4282e3f9} /* (2, 28, 10) {real, imag} */,
  {32'h425083a4, 32'h42973760} /* (2, 28, 9) {real, imag} */,
  {32'h42140978, 32'h42b55b8c} /* (2, 28, 8) {real, imag} */,
  {32'h4255f92c, 32'h42990962} /* (2, 28, 7) {real, imag} */,
  {32'h428cc774, 32'h4293b469} /* (2, 28, 6) {real, imag} */,
  {32'h41f311b4, 32'h424561ef} /* (2, 28, 5) {real, imag} */,
  {32'h41ba8afa, 32'h420fb4b0} /* (2, 28, 4) {real, imag} */,
  {32'h41a27028, 32'h425609d0} /* (2, 28, 3) {real, imag} */,
  {32'h410e7e62, 32'h427023a9} /* (2, 28, 2) {real, imag} */,
  {32'hbf440c10, 32'h41cb2ad4} /* (2, 28, 1) {real, imag} */,
  {32'hc0fdcdc6, 32'h410f1d5e} /* (2, 28, 0) {real, imag} */,
  {32'hc1746af5, 32'hc23e48f4} /* (2, 27, 31) {real, imag} */,
  {32'hc1e3ee14, 32'hc2b46ead} /* (2, 27, 30) {real, imag} */,
  {32'hc1ef82e5, 32'hc297c24f} /* (2, 27, 29) {real, imag} */,
  {32'hc1e2ff91, 32'hc295d945} /* (2, 27, 28) {real, imag} */,
  {32'hc17a6f54, 32'hc22c99d5} /* (2, 27, 27) {real, imag} */,
  {32'hc0edc5ce, 32'hc18b443b} /* (2, 27, 26) {real, imag} */,
  {32'h40aec7fc, 32'hc201dcc2} /* (2, 27, 25) {real, imag} */,
  {32'hc134f530, 32'hc299e3d5} /* (2, 27, 24) {real, imag} */,
  {32'hc1c4ffad, 32'hc29aa840} /* (2, 27, 23) {real, imag} */,
  {32'hc15f89c3, 32'hc26f37bd} /* (2, 27, 22) {real, imag} */,
  {32'hc106d877, 32'hc205ff0f} /* (2, 27, 21) {real, imag} */,
  {32'hc100dccc, 32'h415e8a8b} /* (2, 27, 20) {real, imag} */,
  {32'h41a9a4ba, 32'h41e27913} /* (2, 27, 19) {real, imag} */,
  {32'h4194b5a4, 32'h41862d7c} /* (2, 27, 18) {real, imag} */,
  {32'h41baa0a5, 32'h420b9d15} /* (2, 27, 17) {real, imag} */,
  {32'h419be238, 32'h42513f9c} /* (2, 27, 16) {real, imag} */,
  {32'h4210cf17, 32'h4265ff03} /* (2, 27, 15) {real, imag} */,
  {32'h41a6a8ab, 32'h426059cd} /* (2, 27, 14) {real, imag} */,
  {32'h4055cc0e, 32'h425b638e} /* (2, 27, 13) {real, imag} */,
  {32'h414987b0, 32'h41fe8c37} /* (2, 27, 12) {real, imag} */,
  {32'h415904c6, 32'h4209429c} /* (2, 27, 11) {real, imag} */,
  {32'hc0b1e33a, 32'h4152a706} /* (2, 27, 10) {real, imag} */,
  {32'hbf4b2248, 32'hc1503c0a} /* (2, 27, 9) {real, imag} */,
  {32'hc0315fba, 32'hc0fd088a} /* (2, 27, 8) {real, imag} */,
  {32'h411bc4f5, 32'hc1a7aece} /* (2, 27, 7) {real, imag} */,
  {32'hc040d18c, 32'hc201c6dd} /* (2, 27, 6) {real, imag} */,
  {32'hc160cb6a, 32'hc26d25c0} /* (2, 27, 5) {real, imag} */,
  {32'hc2181e10, 32'hc280e2a0} /* (2, 27, 4) {real, imag} */,
  {32'hc1c44e24, 32'hc25aa956} /* (2, 27, 3) {real, imag} */,
  {32'hc1542f14, 32'hc2379e9e} /* (2, 27, 2) {real, imag} */,
  {32'hc20727ed, 32'hc26ca5a7} /* (2, 27, 1) {real, imag} */,
  {32'hc1b453b4, 32'hc235c4be} /* (2, 27, 0) {real, imag} */,
  {32'hbef67394, 32'hc02faf86} /* (2, 26, 31) {real, imag} */,
  {32'hc0830bfd, 32'hbfbd7852} /* (2, 26, 30) {real, imag} */,
  {32'hc06ac50b, 32'h41833cc5} /* (2, 26, 29) {real, imag} */,
  {32'h4116b066, 32'h4142fff3} /* (2, 26, 28) {real, imag} */,
  {32'h40e5f4f8, 32'h3d9034c0} /* (2, 26, 27) {real, imag} */,
  {32'hc1473600, 32'hc08f0202} /* (2, 26, 26) {real, imag} */,
  {32'hc1d6f262, 32'hc18b27be} /* (2, 26, 25) {real, imag} */,
  {32'hc1857446, 32'hc1723449} /* (2, 26, 24) {real, imag} */,
  {32'hc17e05d0, 32'hc064924c} /* (2, 26, 23) {real, imag} */,
  {32'h402c8cb2, 32'hbda68200} /* (2, 26, 22) {real, imag} */,
  {32'h41a7502a, 32'h4158012c} /* (2, 26, 21) {real, imag} */,
  {32'h41fd9be0, 32'h418483e6} /* (2, 26, 20) {real, imag} */,
  {32'h408fd1b5, 32'h40bcc26d} /* (2, 26, 19) {real, imag} */,
  {32'hc04aaa3c, 32'h417cc002} /* (2, 26, 18) {real, imag} */,
  {32'h40b0bc99, 32'h419ab9a8} /* (2, 26, 17) {real, imag} */,
  {32'h4070fe1a, 32'h3edd76c0} /* (2, 26, 16) {real, imag} */,
  {32'hc070edc4, 32'h408a5e11} /* (2, 26, 15) {real, imag} */,
  {32'h409f6a25, 32'h40e025aa} /* (2, 26, 14) {real, imag} */,
  {32'h40ed42a1, 32'h4193aa60} /* (2, 26, 13) {real, imag} */,
  {32'h411ae6ec, 32'h41b8361b} /* (2, 26, 12) {real, imag} */,
  {32'h4062b24d, 32'hc00ec9cf} /* (2, 26, 11) {real, imag} */,
  {32'h414f3d81, 32'hc1a658d4} /* (2, 26, 10) {real, imag} */,
  {32'h417bfbf8, 32'hc140559c} /* (2, 26, 9) {real, imag} */,
  {32'hbfda1f00, 32'hc0d5e4dc} /* (2, 26, 8) {real, imag} */,
  {32'hc1366232, 32'h411072bc} /* (2, 26, 7) {real, imag} */,
  {32'h41486a9c, 32'hc06631fc} /* (2, 26, 6) {real, imag} */,
  {32'h40dcb014, 32'h3e841020} /* (2, 26, 5) {real, imag} */,
  {32'h40a74104, 32'hc180f3fd} /* (2, 26, 4) {real, imag} */,
  {32'h3fdabb40, 32'hc1c52243} /* (2, 26, 3) {real, imag} */,
  {32'hbfde581c, 32'hc133f938} /* (2, 26, 2) {real, imag} */,
  {32'hc1359c77, 32'h41255a99} /* (2, 26, 1) {real, imag} */,
  {32'hc053a27e, 32'h41c9ac4a} /* (2, 26, 0) {real, imag} */,
  {32'h409efb2b, 32'hc070c327} /* (2, 25, 31) {real, imag} */,
  {32'h41b7b845, 32'h409f3afb} /* (2, 25, 30) {real, imag} */,
  {32'h41a07cb4, 32'h418d1b9b} /* (2, 25, 29) {real, imag} */,
  {32'h414fea26, 32'h419babbf} /* (2, 25, 28) {real, imag} */,
  {32'h40266be0, 32'h41a3c075} /* (2, 25, 27) {real, imag} */,
  {32'h41999cce, 32'hc0120544} /* (2, 25, 26) {real, imag} */,
  {32'h40d171b6, 32'hc114586e} /* (2, 25, 25) {real, imag} */,
  {32'h4167ff7c, 32'hc0bd01fc} /* (2, 25, 24) {real, imag} */,
  {32'h3f394280, 32'h41824644} /* (2, 25, 23) {real, imag} */,
  {32'h41110ee2, 32'h419c871a} /* (2, 25, 22) {real, imag} */,
  {32'hbd394080, 32'h41380d68} /* (2, 25, 21) {real, imag} */,
  {32'hc13799e0, 32'h40f020eb} /* (2, 25, 20) {real, imag} */,
  {32'hc097ac0e, 32'hc109f95f} /* (2, 25, 19) {real, imag} */,
  {32'h3fbba2da, 32'hc1069165} /* (2, 25, 18) {real, imag} */,
  {32'hc09dc696, 32'hc05465a5} /* (2, 25, 17) {real, imag} */,
  {32'hbf529e7e, 32'hc1511f4c} /* (2, 25, 16) {real, imag} */,
  {32'hc19386e0, 32'hc099d32a} /* (2, 25, 15) {real, imag} */,
  {32'hc0d259d7, 32'hc1414aa3} /* (2, 25, 14) {real, imag} */,
  {32'hc040ec8c, 32'h3f675e28} /* (2, 25, 13) {real, imag} */,
  {32'h410a8ea7, 32'h40238978} /* (2, 25, 12) {real, imag} */,
  {32'hc142bdbc, 32'hbffd6800} /* (2, 25, 11) {real, imag} */,
  {32'h408abea9, 32'h405db6fa} /* (2, 25, 10) {real, imag} */,
  {32'h419e3920, 32'hc099172c} /* (2, 25, 9) {real, imag} */,
  {32'hbe72cc00, 32'h3fa464b8} /* (2, 25, 8) {real, imag} */,
  {32'h40b975f0, 32'hc084f97e} /* (2, 25, 7) {real, imag} */,
  {32'h41568f39, 32'hc022421c} /* (2, 25, 6) {real, imag} */,
  {32'h41b53fe7, 32'h410ea6c8} /* (2, 25, 5) {real, imag} */,
  {32'h4182de4c, 32'hc0a1dc58} /* (2, 25, 4) {real, imag} */,
  {32'h419a4a36, 32'h4140f480} /* (2, 25, 3) {real, imag} */,
  {32'h41e6d7fa, 32'h4159a448} /* (2, 25, 2) {real, imag} */,
  {32'h41377dfc, 32'h41921d18} /* (2, 25, 1) {real, imag} */,
  {32'h3fa6d82d, 32'h410c433c} /* (2, 25, 0) {real, imag} */,
  {32'hc1c42fa1, 32'hc1a85ce3} /* (2, 24, 31) {real, imag} */,
  {32'hc1b897ec, 32'hc1aec438} /* (2, 24, 30) {real, imag} */,
  {32'hc115d058, 32'hc1822b14} /* (2, 24, 29) {real, imag} */,
  {32'hc10345d7, 32'hc1d9f0a4} /* (2, 24, 28) {real, imag} */,
  {32'hc14f5dc2, 32'hc1e09a71} /* (2, 24, 27) {real, imag} */,
  {32'hc15a0bf2, 32'hc1816f3b} /* (2, 24, 26) {real, imag} */,
  {32'hc138ef38, 32'hc2150e1a} /* (2, 24, 25) {real, imag} */,
  {32'hc1b30799, 32'hc2074a56} /* (2, 24, 24) {real, imag} */,
  {32'hc1ce9212, 32'hc19e0246} /* (2, 24, 23) {real, imag} */,
  {32'hc17f3b44, 32'hc1c75d0e} /* (2, 24, 22) {real, imag} */,
  {32'h4037b2fc, 32'hc11654b3} /* (2, 24, 21) {real, imag} */,
  {32'h3ebec8c0, 32'h41f772c2} /* (2, 24, 20) {real, imag} */,
  {32'h4088fcff, 32'h4220eca3} /* (2, 24, 19) {real, imag} */,
  {32'h40facefa, 32'h41e3bc00} /* (2, 24, 18) {real, imag} */,
  {32'h40a66608, 32'h41f0a14c} /* (2, 24, 17) {real, imag} */,
  {32'h415f72b4, 32'h41fdc80d} /* (2, 24, 16) {real, imag} */,
  {32'h41db8845, 32'h41bf2100} /* (2, 24, 15) {real, imag} */,
  {32'h419a698f, 32'h41b8f8af} /* (2, 24, 14) {real, imag} */,
  {32'h41eceb43, 32'h42032bd4} /* (2, 24, 13) {real, imag} */,
  {32'h422980e7, 32'h41d5b761} /* (2, 24, 12) {real, imag} */,
  {32'h41c18fe4, 32'h4117df1d} /* (2, 24, 11) {real, imag} */,
  {32'hc0da8790, 32'hc16a06d5} /* (2, 24, 10) {real, imag} */,
  {32'hc1066a13, 32'hc1d55fca} /* (2, 24, 9) {real, imag} */,
  {32'h413ffd14, 32'hc208ac88} /* (2, 24, 8) {real, imag} */,
  {32'h419ae677, 32'hc2072d72} /* (2, 24, 7) {real, imag} */,
  {32'h418e69d3, 32'hc21691ce} /* (2, 24, 6) {real, imag} */,
  {32'h40a6e84e, 32'hc22697fc} /* (2, 24, 5) {real, imag} */,
  {32'hc1fa1054, 32'hc230f6c0} /* (2, 24, 4) {real, imag} */,
  {32'hc1f0a47c, 32'hc21c503e} /* (2, 24, 3) {real, imag} */,
  {32'hc0f7b548, 32'hc24e6827} /* (2, 24, 2) {real, imag} */,
  {32'hc1a6c993, 32'hc23a9f91} /* (2, 24, 1) {real, imag} */,
  {32'hc1b286ee, 32'hc1a2c3f4} /* (2, 24, 0) {real, imag} */,
  {32'hbf39d972, 32'hc0966f80} /* (2, 23, 31) {real, imag} */,
  {32'hc0eea73e, 32'h3f018568} /* (2, 23, 30) {real, imag} */,
  {32'hc1039d71, 32'hc0b2d30e} /* (2, 23, 29) {real, imag} */,
  {32'hc079a076, 32'hc0fcb1c3} /* (2, 23, 28) {real, imag} */,
  {32'h40e7d89f, 32'h3fb47b60} /* (2, 23, 27) {real, imag} */,
  {32'h40b754c0, 32'h3fbaaa18} /* (2, 23, 26) {real, imag} */,
  {32'hbf8e3e7c, 32'h4158465e} /* (2, 23, 25) {real, imag} */,
  {32'hbf720f48, 32'h41dac6e8} /* (2, 23, 24) {real, imag} */,
  {32'hc0823778, 32'h40fdf5f6} /* (2, 23, 23) {real, imag} */,
  {32'h40821cbd, 32'h40d34fa8} /* (2, 23, 22) {real, imag} */,
  {32'hc0f75cb5, 32'h40f02a58} /* (2, 23, 21) {real, imag} */,
  {32'hc1ec2585, 32'hc1a7bdf2} /* (2, 23, 20) {real, imag} */,
  {32'hc1e1cfe6, 32'hc182747a} /* (2, 23, 19) {real, imag} */,
  {32'hc129883a, 32'h40991ab2} /* (2, 23, 18) {real, imag} */,
  {32'hc10764c0, 32'hbff681fe} /* (2, 23, 17) {real, imag} */,
  {32'hc191a97f, 32'hc067cde8} /* (2, 23, 16) {real, imag} */,
  {32'hc0fb0831, 32'hbdcfd780} /* (2, 23, 15) {real, imag} */,
  {32'hbf42a7a8, 32'h412b3b73} /* (2, 23, 14) {real, imag} */,
  {32'hc174a62b, 32'h4130812c} /* (2, 23, 13) {real, imag} */,
  {32'hc0ecad84, 32'h40e4ca4c} /* (2, 23, 12) {real, imag} */,
  {32'hc0417d1e, 32'hbf564da0} /* (2, 23, 11) {real, imag} */,
  {32'h4188742d, 32'hc13f76ec} /* (2, 23, 10) {real, imag} */,
  {32'h41a00cd8, 32'hc16a55bf} /* (2, 23, 9) {real, imag} */,
  {32'h41bca70b, 32'hc175e497} /* (2, 23, 8) {real, imag} */,
  {32'h422df74c, 32'hbf371be0} /* (2, 23, 7) {real, imag} */,
  {32'h420c6968, 32'hc0b42722} /* (2, 23, 6) {real, imag} */,
  {32'h4193dac0, 32'h415889ac} /* (2, 23, 5) {real, imag} */,
  {32'h412e66d7, 32'h3f2fbf40} /* (2, 23, 4) {real, imag} */,
  {32'hc11a3656, 32'hc0fef825} /* (2, 23, 3) {real, imag} */,
  {32'h40f0b67c, 32'h4035fda4} /* (2, 23, 2) {real, imag} */,
  {32'h40cadfe8, 32'h401d4530} /* (2, 23, 1) {real, imag} */,
  {32'h3ff64deb, 32'hbf8dd7c0} /* (2, 23, 0) {real, imag} */,
  {32'h3fda0639, 32'h3fe962cc} /* (2, 22, 31) {real, imag} */,
  {32'h406e5132, 32'h401ffae1} /* (2, 22, 30) {real, imag} */,
  {32'h41460df4, 32'hc08dd9f9} /* (2, 22, 29) {real, imag} */,
  {32'h41ab3899, 32'hc05f67f6} /* (2, 22, 28) {real, imag} */,
  {32'h40d4ede0, 32'hc163cedf} /* (2, 22, 27) {real, imag} */,
  {32'h3f9fe3c4, 32'hc10d8ec1} /* (2, 22, 26) {real, imag} */,
  {32'h3f99c0dc, 32'h40dc504a} /* (2, 22, 25) {real, imag} */,
  {32'hc12f382b, 32'hc08c0632} /* (2, 22, 24) {real, imag} */,
  {32'hbf86e5c0, 32'h409d2742} /* (2, 22, 23) {real, imag} */,
  {32'h4025a2b6, 32'h4116684a} /* (2, 22, 22) {real, imag} */,
  {32'hc15de468, 32'h40411c79} /* (2, 22, 21) {real, imag} */,
  {32'hc1935ce5, 32'hc0d1cff8} /* (2, 22, 20) {real, imag} */,
  {32'hc17c7ede, 32'hc10e1588} /* (2, 22, 19) {real, imag} */,
  {32'hc165083b, 32'hc13aa3f2} /* (2, 22, 18) {real, imag} */,
  {32'hc18a062f, 32'hc0e2208c} /* (2, 22, 17) {real, imag} */,
  {32'hc17a7d4a, 32'hc11113ba} /* (2, 22, 16) {real, imag} */,
  {32'hc0bf2872, 32'h40088366} /* (2, 22, 15) {real, imag} */,
  {32'hbde08720, 32'h4001c065} /* (2, 22, 14) {real, imag} */,
  {32'h408b8bc2, 32'hc0adc44c} /* (2, 22, 13) {real, imag} */,
  {32'h4111f5da, 32'hc08cb624} /* (2, 22, 12) {real, imag} */,
  {32'h411f27ff, 32'h409af236} /* (2, 22, 11) {real, imag} */,
  {32'h418bff60, 32'h40d9e102} /* (2, 22, 10) {real, imag} */,
  {32'h4175b47c, 32'h40770681} /* (2, 22, 9) {real, imag} */,
  {32'h41924a6a, 32'h405fef68} /* (2, 22, 8) {real, imag} */,
  {32'h412fd430, 32'h4104be5c} /* (2, 22, 7) {real, imag} */,
  {32'h411041f0, 32'h415a4c05} /* (2, 22, 6) {real, imag} */,
  {32'hc0100ce8, 32'h4178d356} /* (2, 22, 5) {real, imag} */,
  {32'hc10431b7, 32'hc09d77c0} /* (2, 22, 4) {real, imag} */,
  {32'hc0068e04, 32'h408f6441} /* (2, 22, 3) {real, imag} */,
  {32'h41b5da63, 32'h40b2b170} /* (2, 22, 2) {real, imag} */,
  {32'h41964924, 32'h406361f4} /* (2, 22, 1) {real, imag} */,
  {32'h4102b895, 32'h401e4948} /* (2, 22, 0) {real, imag} */,
  {32'hc120d5cb, 32'hc11a1a7e} /* (2, 21, 31) {real, imag} */,
  {32'hc183a51e, 32'hc1afee3c} /* (2, 21, 30) {real, imag} */,
  {32'hc180b612, 32'hc18a65c5} /* (2, 21, 29) {real, imag} */,
  {32'hc1924c9b, 32'hc19a4cdb} /* (2, 21, 28) {real, imag} */,
  {32'hc13d0e7e, 32'hc1b7edf2} /* (2, 21, 27) {real, imag} */,
  {32'hc0988347, 32'hc1545ee6} /* (2, 21, 26) {real, imag} */,
  {32'hc12fda58, 32'hc11e142a} /* (2, 21, 25) {real, imag} */,
  {32'hc18596ef, 32'hc106b2d4} /* (2, 21, 24) {real, imag} */,
  {32'hc0f71afc, 32'hc10b4bd1} /* (2, 21, 23) {real, imag} */,
  {32'hc18adea4, 32'hc15112a8} /* (2, 21, 22) {real, imag} */,
  {32'hc1404244, 32'hc1829d58} /* (2, 21, 21) {real, imag} */,
  {32'h415f7acc, 32'h3ea509e8} /* (2, 21, 20) {real, imag} */,
  {32'h416ef3c5, 32'h415cc96e} /* (2, 21, 19) {real, imag} */,
  {32'h40d8cab5, 32'h40fbe5ee} /* (2, 21, 18) {real, imag} */,
  {32'h41b18f3a, 32'hbe00f0c0} /* (2, 21, 17) {real, imag} */,
  {32'h41919391, 32'hc1069c2e} /* (2, 21, 16) {real, imag} */,
  {32'h418794f3, 32'hbeac02e0} /* (2, 21, 15) {real, imag} */,
  {32'h4121fc70, 32'h405dea82} /* (2, 21, 14) {real, imag} */,
  {32'h412df4fe, 32'h40b20561} /* (2, 21, 13) {real, imag} */,
  {32'h41137296, 32'h41574c2a} /* (2, 21, 12) {real, imag} */,
  {32'h410472b3, 32'h40f5d728} /* (2, 21, 11) {real, imag} */,
  {32'hc0a1739e, 32'hc0780538} /* (2, 21, 10) {real, imag} */,
  {32'hc126070e, 32'h40670dac} /* (2, 21, 9) {real, imag} */,
  {32'hc1362d78, 32'hc07c5358} /* (2, 21, 8) {real, imag} */,
  {32'h40327eec, 32'hc12680d6} /* (2, 21, 7) {real, imag} */,
  {32'hc0a5accc, 32'hc1b67c9b} /* (2, 21, 6) {real, imag} */,
  {32'hc1820ff0, 32'hc1e4a0ca} /* (2, 21, 5) {real, imag} */,
  {32'hc15375aa, 32'hc1a37ae2} /* (2, 21, 4) {real, imag} */,
  {32'hc190e4d7, 32'hc12b8d2c} /* (2, 21, 3) {real, imag} */,
  {32'hc1a7aad5, 32'hc1b68fb1} /* (2, 21, 2) {real, imag} */,
  {32'hc0afb8c2, 32'hc1607589} /* (2, 21, 1) {real, imag} */,
  {32'hbfd8cec8, 32'hbf3a4cd0} /* (2, 21, 0) {real, imag} */,
  {32'hbfb92906, 32'h4098043d} /* (2, 20, 31) {real, imag} */,
  {32'hbfc6b370, 32'hbd4ec100} /* (2, 20, 30) {real, imag} */,
  {32'hbfeee82c, 32'hc0ca8d60} /* (2, 20, 29) {real, imag} */,
  {32'h3f8284ec, 32'hc08cc877} /* (2, 20, 28) {real, imag} */,
  {32'h404a9c8a, 32'hbf9d5ee0} /* (2, 20, 27) {real, imag} */,
  {32'hc0044245, 32'hbf9c1b88} /* (2, 20, 26) {real, imag} */,
  {32'hc056eea8, 32'hbf746a84} /* (2, 20, 25) {real, imag} */,
  {32'hbe522000, 32'hc09dae62} /* (2, 20, 24) {real, imag} */,
  {32'hc0353f22, 32'h4013ca5c} /* (2, 20, 23) {real, imag} */,
  {32'hc0b02bd2, 32'h40976b0c} /* (2, 20, 22) {real, imag} */,
  {32'hbf9ca4dc, 32'h4019ee06} /* (2, 20, 21) {real, imag} */,
  {32'h4099dfc0, 32'h414d079b} /* (2, 20, 20) {real, imag} */,
  {32'hc100bb23, 32'h40bd19f6} /* (2, 20, 19) {real, imag} */,
  {32'hc12b9496, 32'hc00424e8} /* (2, 20, 18) {real, imag} */,
  {32'hc0b54759, 32'h41191fca} /* (2, 20, 17) {real, imag} */,
  {32'hc0b0882e, 32'h41101479} /* (2, 20, 16) {real, imag} */,
  {32'hc1208824, 32'h40926b85} /* (2, 20, 15) {real, imag} */,
  {32'hc0ad9069, 32'hc0a7b783} /* (2, 20, 14) {real, imag} */,
  {32'h4049ca48, 32'hbfc8607a} /* (2, 20, 13) {real, imag} */,
  {32'h3f8e7e38, 32'h3fed64f0} /* (2, 20, 12) {real, imag} */,
  {32'hc0bee590, 32'hc08f2e3c} /* (2, 20, 11) {real, imag} */,
  {32'hc0cbbafb, 32'h4104bdc6} /* (2, 20, 10) {real, imag} */,
  {32'hbee37cc0, 32'h412ad5c5} /* (2, 20, 9) {real, imag} */,
  {32'hc04911a0, 32'h40419104} /* (2, 20, 8) {real, imag} */,
  {32'hc079f01c, 32'hc006d344} /* (2, 20, 7) {real, imag} */,
  {32'hc02c0b76, 32'h41522c87} /* (2, 20, 6) {real, imag} */,
  {32'hc0abff1d, 32'h40c5ff69} /* (2, 20, 5) {real, imag} */,
  {32'hbf9a7b66, 32'hbfc9dc70} /* (2, 20, 4) {real, imag} */,
  {32'h40bb7f99, 32'h3ff2f748} /* (2, 20, 3) {real, imag} */,
  {32'h40a8b263, 32'h4052bfcc} /* (2, 20, 2) {real, imag} */,
  {32'h4102e1d0, 32'h40df87c4} /* (2, 20, 1) {real, imag} */,
  {32'hbf29ec2c, 32'h3fb4c8ac} /* (2, 20, 0) {real, imag} */,
  {32'h40d1ade6, 32'h40dab16d} /* (2, 19, 31) {real, imag} */,
  {32'h41757eeb, 32'h40b7f4a6} /* (2, 19, 30) {real, imag} */,
  {32'h40be6ada, 32'hbf9ef274} /* (2, 19, 29) {real, imag} */,
  {32'h3eba0e20, 32'h3ea91160} /* (2, 19, 28) {real, imag} */,
  {32'hc12930a4, 32'h40a64220} /* (2, 19, 27) {real, imag} */,
  {32'hbeab13e0, 32'h40aae245} /* (2, 19, 26) {real, imag} */,
  {32'h4138a5f3, 32'h40c104be} /* (2, 19, 25) {real, imag} */,
  {32'h4111c2f3, 32'h40181f88} /* (2, 19, 24) {real, imag} */,
  {32'hc0b88444, 32'h406b34bb} /* (2, 19, 23) {real, imag} */,
  {32'hc11905a5, 32'h4073823a} /* (2, 19, 22) {real, imag} */,
  {32'hc0ca6e51, 32'hc00d89b0} /* (2, 19, 21) {real, imag} */,
  {32'hc094e706, 32'hc0df0822} /* (2, 19, 20) {real, imag} */,
  {32'h3f0590e8, 32'hbfe3b9f8} /* (2, 19, 19) {real, imag} */,
  {32'h3f57e558, 32'hc088faa2} /* (2, 19, 18) {real, imag} */,
  {32'hc038ac6a, 32'hbfa51060} /* (2, 19, 17) {real, imag} */,
  {32'hbe47b080, 32'h3f032128} /* (2, 19, 16) {real, imag} */,
  {32'h4075b390, 32'hc0555070} /* (2, 19, 15) {real, imag} */,
  {32'h40c7eb7f, 32'h3f510c78} /* (2, 19, 14) {real, imag} */,
  {32'hc00cda4a, 32'hc0cd946b} /* (2, 19, 13) {real, imag} */,
  {32'hc021ac19, 32'hc140ec73} /* (2, 19, 12) {real, imag} */,
  {32'h3f997d84, 32'hc1223d2e} /* (2, 19, 11) {real, imag} */,
  {32'h411a1095, 32'h3fc8352c} /* (2, 19, 10) {real, imag} */,
  {32'h40b63119, 32'h40b0f04e} /* (2, 19, 9) {real, imag} */,
  {32'h402cf81e, 32'h4012604a} /* (2, 19, 8) {real, imag} */,
  {32'h40b8d2a8, 32'h3f668ca0} /* (2, 19, 7) {real, imag} */,
  {32'h40ffc574, 32'h3f202c00} /* (2, 19, 6) {real, imag} */,
  {32'h40be9956, 32'h3fa9e596} /* (2, 19, 5) {real, imag} */,
  {32'h4055961a, 32'h3f4ab540} /* (2, 19, 4) {real, imag} */,
  {32'h40f4f646, 32'hbde4a500} /* (2, 19, 3) {real, imag} */,
  {32'h403e3b6a, 32'hbfeadc04} /* (2, 19, 2) {real, imag} */,
  {32'hc046cbce, 32'h41057ac4} /* (2, 19, 1) {real, imag} */,
  {32'h3f40f35c, 32'h414424dc} /* (2, 19, 0) {real, imag} */,
  {32'hc0ce3c73, 32'hbe836bf0} /* (2, 18, 31) {real, imag} */,
  {32'hc1117042, 32'hbfba28c6} /* (2, 18, 30) {real, imag} */,
  {32'hc1200850, 32'h402ceec3} /* (2, 18, 29) {real, imag} */,
  {32'hc10b6f01, 32'h40bca8f8} /* (2, 18, 28) {real, imag} */,
  {32'hc0a29d50, 32'hbfe04118} /* (2, 18, 27) {real, imag} */,
  {32'hc0a723b6, 32'h3f284650} /* (2, 18, 26) {real, imag} */,
  {32'hc0fe18ec, 32'hc0161a28} /* (2, 18, 25) {real, imag} */,
  {32'hc140ac6d, 32'hc0b1409a} /* (2, 18, 24) {real, imag} */,
  {32'hc0c14a82, 32'h3fd8fdd8} /* (2, 18, 23) {real, imag} */,
  {32'hc147c04f, 32'h4033ad86} /* (2, 18, 22) {real, imag} */,
  {32'hc0ded0ff, 32'h41016ca3} /* (2, 18, 21) {real, imag} */,
  {32'hc05ca230, 32'h412d4b8c} /* (2, 18, 20) {real, imag} */,
  {32'h3f9bffb0, 32'h403e1830} /* (2, 18, 19) {real, imag} */,
  {32'h3f65f1c0, 32'h40009f90} /* (2, 18, 18) {real, imag} */,
  {32'hbe2b9500, 32'h3fef7770} /* (2, 18, 17) {real, imag} */,
  {32'h40147940, 32'h40a16672} /* (2, 18, 16) {real, imag} */,
  {32'h4031fb68, 32'h401fe4bc} /* (2, 18, 15) {real, imag} */,
  {32'h3f876b98, 32'h40343e05} /* (2, 18, 14) {real, imag} */,
  {32'h40a71f5a, 32'h4125458c} /* (2, 18, 13) {real, imag} */,
  {32'h417aff28, 32'h40f03d00} /* (2, 18, 12) {real, imag} */,
  {32'h419f4e04, 32'h40294f57} /* (2, 18, 11) {real, imag} */,
  {32'h410b63bc, 32'hc02e9bbe} /* (2, 18, 10) {real, imag} */,
  {32'hbfba1680, 32'hc10318a0} /* (2, 18, 9) {real, imag} */,
  {32'hc05f5b68, 32'hc0e385ce} /* (2, 18, 8) {real, imag} */,
  {32'hc0e8ccb4, 32'hc075ea0c} /* (2, 18, 7) {real, imag} */,
  {32'hc117eed5, 32'hbf5ebcf0} /* (2, 18, 6) {real, imag} */,
  {32'hc03058ba, 32'h40c8ad21} /* (2, 18, 5) {real, imag} */,
  {32'hc0064271, 32'h41311420} /* (2, 18, 4) {real, imag} */,
  {32'hc0ba0f6e, 32'h406c3aa4} /* (2, 18, 3) {real, imag} */,
  {32'hc10cee0a, 32'hc1017d2d} /* (2, 18, 2) {real, imag} */,
  {32'hc09b3c88, 32'hc0d229e2} /* (2, 18, 1) {real, imag} */,
  {32'hbfef75e4, 32'hbed69c00} /* (2, 18, 0) {real, imag} */,
  {32'h40c43ab4, 32'hbe54d3d8} /* (2, 17, 31) {real, imag} */,
  {32'h403801e0, 32'hc049ccfc} /* (2, 17, 30) {real, imag} */,
  {32'h40d947ff, 32'hc07890ff} /* (2, 17, 29) {real, imag} */,
  {32'h408ea4d6, 32'hbe8fbc40} /* (2, 17, 28) {real, imag} */,
  {32'hbd438980, 32'hc06e3b1a} /* (2, 17, 27) {real, imag} */,
  {32'h40912772, 32'hc0882ac7} /* (2, 17, 26) {real, imag} */,
  {32'h40aa5fb8, 32'hc0a50f78} /* (2, 17, 25) {real, imag} */,
  {32'h4066d0bc, 32'hc00a64c0} /* (2, 17, 24) {real, imag} */,
  {32'h405414a8, 32'hc011c688} /* (2, 17, 23) {real, imag} */,
  {32'h40488558, 32'hc0aa50ce} /* (2, 17, 22) {real, imag} */,
  {32'h40856a26, 32'h3f65e600} /* (2, 17, 21) {real, imag} */,
  {32'h3ed6b460, 32'hbec0e680} /* (2, 17, 20) {real, imag} */,
  {32'hc06060a2, 32'hc0814496} /* (2, 17, 19) {real, imag} */,
  {32'hc13e3204, 32'hc0c838fc} /* (2, 17, 18) {real, imag} */,
  {32'hc147af68, 32'h3eebb5b0} /* (2, 17, 17) {real, imag} */,
  {32'hc06543d0, 32'hc0bb2906} /* (2, 17, 16) {real, imag} */,
  {32'h3ff70be8, 32'h3eee1484} /* (2, 17, 15) {real, imag} */,
  {32'hbfd18f58, 32'h408fb61e} /* (2, 17, 14) {real, imag} */,
  {32'hc0ba6da4, 32'h4042f81e} /* (2, 17, 13) {real, imag} */,
  {32'hc04342bc, 32'h3f6e1644} /* (2, 17, 12) {real, imag} */,
  {32'hc044670e, 32'hc06603d0} /* (2, 17, 11) {real, imag} */,
  {32'h410c10cc, 32'hc01011c6} /* (2, 17, 10) {real, imag} */,
  {32'h40af5216, 32'h4043d578} /* (2, 17, 9) {real, imag} */,
  {32'h40d8f8a4, 32'h3ffbb260} /* (2, 17, 8) {real, imag} */,
  {32'h413b865c, 32'hbf338320} /* (2, 17, 7) {real, imag} */,
  {32'h4180085b, 32'hbf087330} /* (2, 17, 6) {real, imag} */,
  {32'h414ae865, 32'h3f5ebf74} /* (2, 17, 5) {real, imag} */,
  {32'h40cb314a, 32'hc0112df4} /* (2, 17, 4) {real, imag} */,
  {32'h3fc3421c, 32'hbfc07e30} /* (2, 17, 3) {real, imag} */,
  {32'hc00387b4, 32'hc005e144} /* (2, 17, 2) {real, imag} */,
  {32'h408b6c24, 32'h3efc8160} /* (2, 17, 1) {real, imag} */,
  {32'h40bb5988, 32'h3f8c6315} /* (2, 17, 0) {real, imag} */,
  {32'hc04ae9d0, 32'hc03092b0} /* (2, 16, 31) {real, imag} */,
  {32'hc02783b0, 32'hc0c3b3c0} /* (2, 16, 30) {real, imag} */,
  {32'hbfe220b8, 32'hc02c3b40} /* (2, 16, 29) {real, imag} */,
  {32'hbe3e6c80, 32'h3fa4cc80} /* (2, 16, 28) {real, imag} */,
  {32'hbff2fb30, 32'hbfa73400} /* (2, 16, 27) {real, imag} */,
  {32'hc05e43ac, 32'h3fc9bb00} /* (2, 16, 26) {real, imag} */,
  {32'h3f20ea78, 32'hc066b5c0} /* (2, 16, 25) {real, imag} */,
  {32'h401b90a8, 32'hc0a8d770} /* (2, 16, 24) {real, imag} */,
  {32'h40bf2d08, 32'h4008b260} /* (2, 16, 23) {real, imag} */,
  {32'h3e88e440, 32'hc02aa180} /* (2, 16, 22) {real, imag} */,
  {32'h3fa340d8, 32'hc0ba0228} /* (2, 16, 21) {real, imag} */,
  {32'h4037fcdf, 32'hbfa54340} /* (2, 16, 20) {real, imag} */,
  {32'hbdef0600, 32'h400ad544} /* (2, 16, 19) {real, imag} */,
  {32'hbf993fc0, 32'hbe3406c0} /* (2, 16, 18) {real, imag} */,
  {32'hbfcbe260, 32'h3f83c818} /* (2, 16, 17) {real, imag} */,
  {32'h3fcd3230, 32'h3e46c500} /* (2, 16, 16) {real, imag} */,
  {32'hbfe2194c, 32'hc013c760} /* (2, 16, 15) {real, imag} */,
  {32'hbd93c580, 32'hbc73e000} /* (2, 16, 14) {real, imag} */,
  {32'hc03965d0, 32'hbcf85000} /* (2, 16, 13) {real, imag} */,
  {32'hc0a4b6d0, 32'hbfcf7100} /* (2, 16, 12) {real, imag} */,
  {32'hc04e3640, 32'h402a4000} /* (2, 16, 11) {real, imag} */,
  {32'hc05ed310, 32'h3fd67380} /* (2, 16, 10) {real, imag} */,
  {32'hc083b256, 32'h405a4404} /* (2, 16, 9) {real, imag} */,
  {32'h3ed5ba20, 32'h40ad9082} /* (2, 16, 8) {real, imag} */,
  {32'h409be370, 32'h40cc8d80} /* (2, 16, 7) {real, imag} */,
  {32'h3f8da4e2, 32'h403c9a16} /* (2, 16, 6) {real, imag} */,
  {32'hc10276bc, 32'hc112b8b0} /* (2, 16, 5) {real, imag} */,
  {32'hc0b50fa4, 32'hc0b4f6c0} /* (2, 16, 4) {real, imag} */,
  {32'hc01e655f, 32'hc080bb00} /* (2, 16, 3) {real, imag} */,
  {32'hc0ffeca8, 32'h3e457000} /* (2, 16, 2) {real, imag} */,
  {32'hc0134060, 32'h3f968de0} /* (2, 16, 1) {real, imag} */,
  {32'hc01ddb60, 32'h407b8020} /* (2, 16, 0) {real, imag} */,
  {32'hc0e16434, 32'hbfea6c05} /* (2, 15, 31) {real, imag} */,
  {32'hc083b4f8, 32'hc09ad8a2} /* (2, 15, 30) {real, imag} */,
  {32'h3fef65c4, 32'hc0b3b980} /* (2, 15, 29) {real, imag} */,
  {32'hc0eb8a0e, 32'hc06e8d78} /* (2, 15, 28) {real, imag} */,
  {32'hc140d9a6, 32'hc0992d33} /* (2, 15, 27) {real, imag} */,
  {32'hc0b1025a, 32'hc02e5d72} /* (2, 15, 26) {real, imag} */,
  {32'hc044bb60, 32'h40443870} /* (2, 15, 25) {real, imag} */,
  {32'h406e8cb4, 32'h409a5580} /* (2, 15, 24) {real, imag} */,
  {32'h4019cce8, 32'h4038ee08} /* (2, 15, 23) {real, imag} */,
  {32'hc0ab1e7c, 32'h3fb640b8} /* (2, 15, 22) {real, imag} */,
  {32'hc10f2297, 32'h40b81480} /* (2, 15, 21) {real, imag} */,
  {32'hc02a5fb4, 32'h4105778c} /* (2, 15, 20) {real, imag} */,
  {32'h40e7117f, 32'h40ec7e06} /* (2, 15, 19) {real, imag} */,
  {32'h40f49268, 32'h40589e78} /* (2, 15, 18) {real, imag} */,
  {32'h40285e1e, 32'hc04d81f6} /* (2, 15, 17) {real, imag} */,
  {32'hc03850d0, 32'hc02c93b4} /* (2, 15, 16) {real, imag} */,
  {32'h3ffdac78, 32'hc0047590} /* (2, 15, 15) {real, imag} */,
  {32'h40ff3766, 32'hc098185e} /* (2, 15, 14) {real, imag} */,
  {32'h40c8af64, 32'hc0cc2c4f} /* (2, 15, 13) {real, imag} */,
  {32'hc0036be4, 32'h3e972d78} /* (2, 15, 12) {real, imag} */,
  {32'hbf4f700a, 32'h4107b344} /* (2, 15, 11) {real, imag} */,
  {32'hc01ae6ae, 32'h40b324a9} /* (2, 15, 10) {real, imag} */,
  {32'hbfd607a8, 32'h40940554} /* (2, 15, 9) {real, imag} */,
  {32'h3f79daa0, 32'hbedf8380} /* (2, 15, 8) {real, imag} */,
  {32'hc04ceb10, 32'hc0041af8} /* (2, 15, 7) {real, imag} */,
  {32'hc1015a2b, 32'hc01fa4d4} /* (2, 15, 6) {real, imag} */,
  {32'hc0e3bfae, 32'hc0cff40e} /* (2, 15, 5) {real, imag} */,
  {32'hc03c03f4, 32'hc0c92146} /* (2, 15, 4) {real, imag} */,
  {32'h3e437d20, 32'hc014a328} /* (2, 15, 3) {real, imag} */,
  {32'hbf99d5d8, 32'hc0b39dde} /* (2, 15, 2) {real, imag} */,
  {32'h3f0c52a0, 32'hc08ab556} /* (2, 15, 1) {real, imag} */,
  {32'h3f463080, 32'hbfdf29d5} /* (2, 15, 0) {real, imag} */,
  {32'hbf99f014, 32'hbfadb404} /* (2, 14, 31) {real, imag} */,
  {32'h402fd5f8, 32'h3f29158c} /* (2, 14, 30) {real, imag} */,
  {32'h407c28fe, 32'hc0351d83} /* (2, 14, 29) {real, imag} */,
  {32'h41153263, 32'h40032b10} /* (2, 14, 28) {real, imag} */,
  {32'h4155b180, 32'h40673f0c} /* (2, 14, 27) {real, imag} */,
  {32'h4173aaeb, 32'h3fc0add8} /* (2, 14, 26) {real, imag} */,
  {32'h414f6554, 32'h3ec31540} /* (2, 14, 25) {real, imag} */,
  {32'h416e7c77, 32'h3e374730} /* (2, 14, 24) {real, imag} */,
  {32'h411b04ff, 32'hc0beabf6} /* (2, 14, 23) {real, imag} */,
  {32'h40b1cde2, 32'hc0a9f263} /* (2, 14, 22) {real, imag} */,
  {32'h3f754d88, 32'h3f97b5a8} /* (2, 14, 21) {real, imag} */,
  {32'hc0861b48, 32'h41163874} /* (2, 14, 20) {real, imag} */,
  {32'hc0cc1324, 32'h410e48c4} /* (2, 14, 19) {real, imag} */,
  {32'hbe820a80, 32'h3f37c3c0} /* (2, 14, 18) {real, imag} */,
  {32'hbe98a480, 32'hbfa53df0} /* (2, 14, 17) {real, imag} */,
  {32'hc0279060, 32'h4064339c} /* (2, 14, 16) {real, imag} */,
  {32'hc09e5f84, 32'h40f24b82} /* (2, 14, 15) {real, imag} */,
  {32'hc1654841, 32'h40c04d5e} /* (2, 14, 14) {real, imag} */,
  {32'hc188f502, 32'h3fdc0d9c} /* (2, 14, 13) {real, imag} */,
  {32'hc184971c, 32'hc03d8480} /* (2, 14, 12) {real, imag} */,
  {32'hc083608a, 32'hc05d5e17} /* (2, 14, 11) {real, imag} */,
  {32'h4102cecc, 32'h40a5401f} /* (2, 14, 10) {real, imag} */,
  {32'h414ad868, 32'hbfab4d82} /* (2, 14, 9) {real, imag} */,
  {32'h411676fe, 32'hc0a51732} /* (2, 14, 8) {real, imag} */,
  {32'h40837094, 32'hc09d7dba} /* (2, 14, 7) {real, imag} */,
  {32'h40c24f56, 32'hc0a3c8e2} /* (2, 14, 6) {real, imag} */,
  {32'h41145dba, 32'h4054353e} /* (2, 14, 5) {real, imag} */,
  {32'h402846e9, 32'h40aa4e80} /* (2, 14, 4) {real, imag} */,
  {32'h4048ad14, 32'h3feac2b8} /* (2, 14, 3) {real, imag} */,
  {32'h40779178, 32'hbddb4960} /* (2, 14, 2) {real, imag} */,
  {32'h40ea3d08, 32'hc0823f5e} /* (2, 14, 1) {real, imag} */,
  {32'h41127670, 32'hc090cdd0} /* (2, 14, 0) {real, imag} */,
  {32'hc029338b, 32'h3f118758} /* (2, 13, 31) {real, imag} */,
  {32'hc0657c3c, 32'h409b04e2} /* (2, 13, 30) {real, imag} */,
  {32'hbff36450, 32'h40969521} /* (2, 13, 29) {real, imag} */,
  {32'hbf980388, 32'h40afa7f6} /* (2, 13, 28) {real, imag} */,
  {32'h402575f2, 32'h40873838} /* (2, 13, 27) {real, imag} */,
  {32'h3daf6d80, 32'h401d6c4a} /* (2, 13, 26) {real, imag} */,
  {32'hbff7b0c8, 32'hbc370c00} /* (2, 13, 25) {real, imag} */,
  {32'hbfacb6ea, 32'h3edf5300} /* (2, 13, 24) {real, imag} */,
  {32'hbf5f53e0, 32'h40aa0d63} /* (2, 13, 23) {real, imag} */,
  {32'h40fe9c8e, 32'h406ba356} /* (2, 13, 22) {real, imag} */,
  {32'h3fa45cb4, 32'hbfa1d220} /* (2, 13, 21) {real, imag} */,
  {32'hbfd9319a, 32'hc05fa40b} /* (2, 13, 20) {real, imag} */,
  {32'hbf906b0c, 32'hc0076774} /* (2, 13, 19) {real, imag} */,
  {32'h40d82b2b, 32'h409b4006} /* (2, 13, 18) {real, imag} */,
  {32'h4122f9d6, 32'h4058aca0} /* (2, 13, 17) {real, imag} */,
  {32'h408427fc, 32'h3d6af680} /* (2, 13, 16) {real, imag} */,
  {32'hc06f3f60, 32'h4067d1b4} /* (2, 13, 15) {real, imag} */,
  {32'hc01a4842, 32'h40c2cefd} /* (2, 13, 14) {real, imag} */,
  {32'h3eebe2f0, 32'h40f23945} /* (2, 13, 13) {real, imag} */,
  {32'hbf0a536c, 32'h40eb3252} /* (2, 13, 12) {real, imag} */,
  {32'hbf281478, 32'h3f945d8c} /* (2, 13, 11) {real, imag} */,
  {32'hc090aa76, 32'hbfe51424} /* (2, 13, 10) {real, imag} */,
  {32'h409f3c49, 32'h3f940b28} /* (2, 13, 9) {real, imag} */,
  {32'h3d8757c0, 32'hbfe686ac} /* (2, 13, 8) {real, imag} */,
  {32'hc0fa1238, 32'hc03f30d0} /* (2, 13, 7) {real, imag} */,
  {32'hc03afe98, 32'hc0805794} /* (2, 13, 6) {real, imag} */,
  {32'h3e0619c0, 32'hbf0f1f4c} /* (2, 13, 5) {real, imag} */,
  {32'h40b33c49, 32'h3f087fc0} /* (2, 13, 4) {real, imag} */,
  {32'h4088e576, 32'hc07c2970} /* (2, 13, 3) {real, imag} */,
  {32'h404393fa, 32'hc0432ce6} /* (2, 13, 2) {real, imag} */,
  {32'hbfdc4724, 32'hbfc682a4} /* (2, 13, 1) {real, imag} */,
  {32'hc031675d, 32'h3ed9db30} /* (2, 13, 0) {real, imag} */,
  {32'hbf50629d, 32'hbf200698} /* (2, 12, 31) {real, imag} */,
  {32'hc08bfcb1, 32'h411cd82f} /* (2, 12, 30) {real, imag} */,
  {32'h3fef26c4, 32'h415d922a} /* (2, 12, 29) {real, imag} */,
  {32'h40f871f5, 32'h40c1ce7f} /* (2, 12, 28) {real, imag} */,
  {32'hbf5af5d6, 32'hc03a5bb0} /* (2, 12, 27) {real, imag} */,
  {32'hc0760445, 32'hbf7d12f0} /* (2, 12, 26) {real, imag} */,
  {32'hc0b3c426, 32'hbf98f81e} /* (2, 12, 25) {real, imag} */,
  {32'hc137899b, 32'hc0f4ed3e} /* (2, 12, 24) {real, imag} */,
  {32'hc13c3978, 32'hc062f90c} /* (2, 12, 23) {real, imag} */,
  {32'hbf993c30, 32'hc0518c38} /* (2, 12, 22) {real, imag} */,
  {32'h415c1bbe, 32'hc10069e0} /* (2, 12, 21) {real, imag} */,
  {32'h415352b8, 32'h3fde6a68} /* (2, 12, 20) {real, imag} */,
  {32'h3fe489ea, 32'h3f827808} /* (2, 12, 19) {real, imag} */,
  {32'hc00ab0b8, 32'h4002a628} /* (2, 12, 18) {real, imag} */,
  {32'h40e31897, 32'hc0c7d475} /* (2, 12, 17) {real, imag} */,
  {32'h408a7a42, 32'hc08ac372} /* (2, 12, 16) {real, imag} */,
  {32'hc027f462, 32'hc03203aa} /* (2, 12, 15) {real, imag} */,
  {32'hc106767a, 32'hbfc8f674} /* (2, 12, 14) {real, imag} */,
  {32'hc183b665, 32'h4006460d} /* (2, 12, 13) {real, imag} */,
  {32'hc098bb58, 32'hc0061d18} /* (2, 12, 12) {real, imag} */,
  {32'hc0c3486a, 32'hc0873a20} /* (2, 12, 11) {real, imag} */,
  {32'hc04b8896, 32'h40860784} /* (2, 12, 10) {real, imag} */,
  {32'h40c6267c, 32'h4010e47c} /* (2, 12, 9) {real, imag} */,
  {32'h411b5d34, 32'h3f1314f0} /* (2, 12, 8) {real, imag} */,
  {32'h3fd7fca8, 32'h40409164} /* (2, 12, 7) {real, imag} */,
  {32'hc04a91d6, 32'h406d06e4} /* (2, 12, 6) {real, imag} */,
  {32'h3f955a6c, 32'hbfb91744} /* (2, 12, 5) {real, imag} */,
  {32'hbef9be98, 32'hbf85a9d0} /* (2, 12, 4) {real, imag} */,
  {32'hc04a2efe, 32'h40d0d57a} /* (2, 12, 3) {real, imag} */,
  {32'hc0a00f79, 32'h404fd6a4} /* (2, 12, 2) {real, imag} */,
  {32'h3f9100b4, 32'h3f8634f0} /* (2, 12, 1) {real, imag} */,
  {32'hbdd05220, 32'hc0426da6} /* (2, 12, 0) {real, imag} */,
  {32'h409bd892, 32'hbfe22034} /* (2, 11, 31) {real, imag} */,
  {32'hbf8015d8, 32'hc0a3a006} /* (2, 11, 30) {real, imag} */,
  {32'h40c53711, 32'hc132dbc6} /* (2, 11, 29) {real, imag} */,
  {32'h41b519b3, 32'hc12dd85a} /* (2, 11, 28) {real, imag} */,
  {32'h41e4ef27, 32'hc156f2f0} /* (2, 11, 27) {real, imag} */,
  {32'h41712d14, 32'hc1860b78} /* (2, 11, 26) {real, imag} */,
  {32'h4192bf47, 32'hc1614b8e} /* (2, 11, 25) {real, imag} */,
  {32'h41b35199, 32'hc15dfecc} /* (2, 11, 24) {real, imag} */,
  {32'h41b37b19, 32'hc17de01f} /* (2, 11, 23) {real, imag} */,
  {32'h418ecec0, 32'hc1594608} /* (2, 11, 22) {real, imag} */,
  {32'h416c2964, 32'hc0143684} /* (2, 11, 21) {real, imag} */,
  {32'h410e4286, 32'hc09859f6} /* (2, 11, 20) {real, imag} */,
  {32'h3f9e7498, 32'hc11b7f2e} /* (2, 11, 19) {real, imag} */,
  {32'h3f20d3c8, 32'hc0aded6e} /* (2, 11, 18) {real, imag} */,
  {32'hc0e19390, 32'hbf52bc90} /* (2, 11, 17) {real, imag} */,
  {32'hc10e7472, 32'hbfa089f0} /* (2, 11, 16) {real, imag} */,
  {32'hc18064b9, 32'hc11daf5d} /* (2, 11, 15) {real, imag} */,
  {32'hc1d46534, 32'hc0b65659} /* (2, 11, 14) {real, imag} */,
  {32'hc16fa462, 32'h3fc8d7fc} /* (2, 11, 13) {real, imag} */,
  {32'hc1584664, 32'hc0ce431c} /* (2, 11, 12) {real, imag} */,
  {32'hc09a582c, 32'h4105e1a4} /* (2, 11, 11) {real, imag} */,
  {32'h4124e645, 32'h40b14da0} /* (2, 11, 10) {real, imag} */,
  {32'h4128bf20, 32'hbe9e3260} /* (2, 11, 9) {real, imag} */,
  {32'hc001c986, 32'hc078be10} /* (2, 11, 8) {real, imag} */,
  {32'h41b80f54, 32'hc10e9f8e} /* (2, 11, 7) {real, imag} */,
  {32'h420274e2, 32'hc14c46a6} /* (2, 11, 6) {real, imag} */,
  {32'h41a2f5d6, 32'hc181f654} /* (2, 11, 5) {real, imag} */,
  {32'h41eefaab, 32'hc1738e4f} /* (2, 11, 4) {real, imag} */,
  {32'h41b41f37, 32'hc129bd50} /* (2, 11, 3) {real, imag} */,
  {32'h418a33b3, 32'hc15489ee} /* (2, 11, 2) {real, imag} */,
  {32'h41379a6b, 32'hc14342ef} /* (2, 11, 1) {real, imag} */,
  {32'h4109ad12, 32'hc0d77872} /* (2, 11, 0) {real, imag} */,
  {32'hbf2b885e, 32'h40fcb211} /* (2, 10, 31) {real, imag} */,
  {32'hc15749b2, 32'h40a18f0c} /* (2, 10, 30) {real, imag} */,
  {32'hc147291a, 32'h41162f14} /* (2, 10, 29) {real, imag} */,
  {32'hc10edaea, 32'h4019af0e} /* (2, 10, 28) {real, imag} */,
  {32'hbf6cfa90, 32'hc04f6394} /* (2, 10, 27) {real, imag} */,
  {32'h3e904090, 32'hc00f20f4} /* (2, 10, 26) {real, imag} */,
  {32'hc0a587d9, 32'hc12f4a67} /* (2, 10, 25) {real, imag} */,
  {32'hc1520d57, 32'hbf6a8d70} /* (2, 10, 24) {real, imag} */,
  {32'h40b98960, 32'h415011ef} /* (2, 10, 23) {real, imag} */,
  {32'h409e6ddb, 32'h40a68118} /* (2, 10, 22) {real, imag} */,
  {32'hc124f73a, 32'hc04b7e79} /* (2, 10, 21) {real, imag} */,
  {32'h40bba09b, 32'hc10dad00} /* (2, 10, 20) {real, imag} */,
  {32'h40a676fb, 32'hc0bca113} /* (2, 10, 19) {real, imag} */,
  {32'h4181adf2, 32'hc08b985c} /* (2, 10, 18) {real, imag} */,
  {32'h41dc9df1, 32'hc1807d10} /* (2, 10, 17) {real, imag} */,
  {32'h419fe7e3, 32'hc144125e} /* (2, 10, 16) {real, imag} */,
  {32'h4081a1d6, 32'h3f9674b4} /* (2, 10, 15) {real, imag} */,
  {32'h40e04442, 32'h3d918860} /* (2, 10, 14) {real, imag} */,
  {32'h4182e0c0, 32'hc0c4eb98} /* (2, 10, 13) {real, imag} */,
  {32'h416a72d6, 32'hc0b9d400} /* (2, 10, 12) {real, imag} */,
  {32'h4063d015, 32'h40a520a6} /* (2, 10, 11) {real, imag} */,
  {32'hc0b87abe, 32'h4025c8b4} /* (2, 10, 10) {real, imag} */,
  {32'hc1b79bba, 32'hc0093ef1} /* (2, 10, 9) {real, imag} */,
  {32'hc1e88c1e, 32'h40e09990} /* (2, 10, 8) {real, imag} */,
  {32'hc113de9c, 32'h414f8808} /* (2, 10, 7) {real, imag} */,
  {32'hc1b33560, 32'h40b1667a} /* (2, 10, 6) {real, imag} */,
  {32'hc10296bc, 32'h40a275a0} /* (2, 10, 5) {real, imag} */,
  {32'hbfc3d746, 32'h41be7894} /* (2, 10, 4) {real, imag} */,
  {32'h4035e9ec, 32'h410a9d4c} /* (2, 10, 3) {real, imag} */,
  {32'hbffe33f0, 32'hc0218988} /* (2, 10, 2) {real, imag} */,
  {32'hc0220f1c, 32'h413c9b59} /* (2, 10, 1) {real, imag} */,
  {32'hbfc7fdbe, 32'h4158743e} /* (2, 10, 0) {real, imag} */,
  {32'hc033a3a6, 32'h41571a6a} /* (2, 9, 31) {real, imag} */,
  {32'h3f73456c, 32'h41563d58} /* (2, 9, 30) {real, imag} */,
  {32'h40c81f6e, 32'h41086791} /* (2, 9, 29) {real, imag} */,
  {32'h40e6c845, 32'hc0886e29} /* (2, 9, 28) {real, imag} */,
  {32'h411e7e38, 32'hc0fb2ad4} /* (2, 9, 27) {real, imag} */,
  {32'h40382a9b, 32'hc164a17b} /* (2, 9, 26) {real, imag} */,
  {32'h40f67cc5, 32'hc120d806} /* (2, 9, 25) {real, imag} */,
  {32'h40f3a3e7, 32'hc170d059} /* (2, 9, 24) {real, imag} */,
  {32'h417cb9a2, 32'hc09f5bfe} /* (2, 9, 23) {real, imag} */,
  {32'h40966723, 32'h40d606d4} /* (2, 9, 22) {real, imag} */,
  {32'h40b70beb, 32'hc13cda76} /* (2, 9, 21) {real, imag} */,
  {32'h414929f6, 32'hc1266756} /* (2, 9, 20) {real, imag} */,
  {32'h418f9bcc, 32'hc13bd6d0} /* (2, 9, 19) {real, imag} */,
  {32'h41a6e511, 32'h411572eb} /* (2, 9, 18) {real, imag} */,
  {32'h41addc3a, 32'h4098e0d0} /* (2, 9, 17) {real, imag} */,
  {32'h419374bb, 32'h4104bda2} /* (2, 9, 16) {real, imag} */,
  {32'h419a462a, 32'h41a624a0} /* (2, 9, 15) {real, imag} */,
  {32'h400caede, 32'h402c421c} /* (2, 9, 14) {real, imag} */,
  {32'hc0a7757e, 32'hc063c0a6} /* (2, 9, 13) {real, imag} */,
  {32'hbf9e78a2, 32'h40c45560} /* (2, 9, 12) {real, imag} */,
  {32'h40d73cab, 32'h4127b974} /* (2, 9, 11) {real, imag} */,
  {32'hc15758fe, 32'h4018d38e} /* (2, 9, 10) {real, imag} */,
  {32'hc20faa6d, 32'hc0e39f9a} /* (2, 9, 9) {real, imag} */,
  {32'hc1ddea7f, 32'hc0c064aa} /* (2, 9, 8) {real, imag} */,
  {32'hc1d84b78, 32'hc19e9d59} /* (2, 9, 7) {real, imag} */,
  {32'hc19eff0e, 32'hc1a05432} /* (2, 9, 6) {real, imag} */,
  {32'hbdf55000, 32'hc07b15c0} /* (2, 9, 5) {real, imag} */,
  {32'h4082619a, 32'h40d3e078} /* (2, 9, 4) {real, imag} */,
  {32'hc0d284a1, 32'h4031cd7a} /* (2, 9, 3) {real, imag} */,
  {32'h3ff65380, 32'h40d83a88} /* (2, 9, 2) {real, imag} */,
  {32'hbeeaa5a0, 32'hc09ab4c8} /* (2, 9, 1) {real, imag} */,
  {32'hc057c806, 32'hc02d5984} /* (2, 9, 0) {real, imag} */,
  {32'h41244f96, 32'hc10fa862} /* (2, 8, 31) {real, imag} */,
  {32'h41a33780, 32'hc1a63ac8} /* (2, 8, 30) {real, imag} */,
  {32'h41e96068, 32'hc16ff1f9} /* (2, 8, 29) {real, imag} */,
  {32'h41f09c4e, 32'hc1569d6f} /* (2, 8, 28) {real, imag} */,
  {32'h4199ca03, 32'hc1738422} /* (2, 8, 27) {real, imag} */,
  {32'h41cdf2a3, 32'hc1715c12} /* (2, 8, 26) {real, imag} */,
  {32'h42296144, 32'hc1eeda7c} /* (2, 8, 25) {real, imag} */,
  {32'h41f268b5, 32'hc2087536} /* (2, 8, 24) {real, imag} */,
  {32'h4181d9f8, 32'hc1eda5ae} /* (2, 8, 23) {real, imag} */,
  {32'h41756e74, 32'hc155da1c} /* (2, 8, 22) {real, imag} */,
  {32'h413aea13, 32'h40ed9956} /* (2, 8, 21) {real, imag} */,
  {32'hc07f1110, 32'h41c8edc6} /* (2, 8, 20) {real, imag} */,
  {32'hbe0fcaa0, 32'h41d730d2} /* (2, 8, 19) {real, imag} */,
  {32'h413c9193, 32'h4237f4a2} /* (2, 8, 18) {real, imag} */,
  {32'h3f5e7f5c, 32'h4257cf3c} /* (2, 8, 17) {real, imag} */,
  {32'hc1e4f81e, 32'h4204ee17} /* (2, 8, 16) {real, imag} */,
  {32'hc20f83c9, 32'h3ffb3eb8} /* (2, 8, 15) {real, imag} */,
  {32'hc21caf34, 32'h41a98fa1} /* (2, 8, 14) {real, imag} */,
  {32'hc21f159a, 32'h42076be2} /* (2, 8, 13) {real, imag} */,
  {32'hc1f95552, 32'h41bf3e61} /* (2, 8, 12) {real, imag} */,
  {32'hc190a510, 32'hc0a506ea} /* (2, 8, 11) {real, imag} */,
  {32'hc129e590, 32'hc1f96632} /* (2, 8, 10) {real, imag} */,
  {32'h41683717, 32'hc1941188} /* (2, 8, 9) {real, imag} */,
  {32'h4126fd9e, 32'hc1462982} /* (2, 8, 8) {real, imag} */,
  {32'h4168f13e, 32'hc1e5cef0} /* (2, 8, 7) {real, imag} */,
  {32'h3fe6acb4, 32'hc1f425a4} /* (2, 8, 6) {real, imag} */,
  {32'h413e0aaf, 32'hc198c8fb} /* (2, 8, 5) {real, imag} */,
  {32'h41a98e28, 32'hc18bf993} /* (2, 8, 4) {real, imag} */,
  {32'h416ee558, 32'hc1cbab3c} /* (2, 8, 3) {real, imag} */,
  {32'h416f0884, 32'hc1bb998a} /* (2, 8, 2) {real, imag} */,
  {32'h419837b5, 32'hc14ed004} /* (2, 8, 1) {real, imag} */,
  {32'h4128965c, 32'h405f1760} /* (2, 8, 0) {real, imag} */,
  {32'hc0ecd711, 32'h3f675104} /* (2, 7, 31) {real, imag} */,
  {32'hc1665fce, 32'h415c9164} /* (2, 7, 30) {real, imag} */,
  {32'hc11701b1, 32'h41789c92} /* (2, 7, 29) {real, imag} */,
  {32'hc18df5ed, 32'h41c46f0d} /* (2, 7, 28) {real, imag} */,
  {32'hc1611d10, 32'h41f652cb} /* (2, 7, 27) {real, imag} */,
  {32'h3f374570, 32'h41b2605c} /* (2, 7, 26) {real, imag} */,
  {32'h3ede6138, 32'h40f33f6b} /* (2, 7, 25) {real, imag} */,
  {32'hc15093cc, 32'h41c0c87c} /* (2, 7, 24) {real, imag} */,
  {32'hc159b606, 32'h41ccc9fe} /* (2, 7, 23) {real, imag} */,
  {32'hc079e385, 32'h407881b8} /* (2, 7, 22) {real, imag} */,
  {32'h40afd6ef, 32'hc0798776} /* (2, 7, 21) {real, imag} */,
  {32'hc0068ffe, 32'hc07957de} /* (2, 7, 20) {real, imag} */,
  {32'hc103d933, 32'hc1229c8d} /* (2, 7, 19) {real, imag} */,
  {32'h409edc5e, 32'hc0b1b14d} /* (2, 7, 18) {real, imag} */,
  {32'h40a5fa92, 32'hbefb9ed8} /* (2, 7, 17) {real, imag} */,
  {32'hbfa91fdf, 32'hc1000a1c} /* (2, 7, 16) {real, imag} */,
  {32'h415d52d4, 32'h404d0d0c} /* (2, 7, 15) {real, imag} */,
  {32'h40ef1345, 32'h4150d609} /* (2, 7, 14) {real, imag} */,
  {32'h41c3dec8, 32'hc11c81a4} /* (2, 7, 13) {real, imag} */,
  {32'h41c7bd3c, 32'hc184f01a} /* (2, 7, 12) {real, imag} */,
  {32'h402aed1a, 32'hc1792c1a} /* (2, 7, 11) {real, imag} */,
  {32'hc18eaaaa, 32'hbf82f0b3} /* (2, 7, 10) {real, imag} */,
  {32'hc1749c45, 32'h41248ee2} /* (2, 7, 9) {real, imag} */,
  {32'hc0545190, 32'hc107e613} /* (2, 7, 8) {real, imag} */,
  {32'hc18ce2f0, 32'hc109b439} /* (2, 7, 7) {real, imag} */,
  {32'hc17f24e3, 32'h414885ab} /* (2, 7, 6) {real, imag} */,
  {32'hc1830be9, 32'h4152d45c} /* (2, 7, 5) {real, imag} */,
  {32'h3f82ab08, 32'h411c7f5c} /* (2, 7, 4) {real, imag} */,
  {32'h4016d064, 32'h41cb900a} /* (2, 7, 3) {real, imag} */,
  {32'hc101f54b, 32'h40ad37b9} /* (2, 7, 2) {real, imag} */,
  {32'hc0dd0d67, 32'hbffa5f40} /* (2, 7, 1) {real, imag} */,
  {32'hbf85c79b, 32'h40c5c29a} /* (2, 7, 0) {real, imag} */,
  {32'h407dea02, 32'hbf87dd44} /* (2, 6, 31) {real, imag} */,
  {32'h419254e8, 32'hc1023a64} /* (2, 6, 30) {real, imag} */,
  {32'h40c34ed6, 32'h3fdffff4} /* (2, 6, 29) {real, imag} */,
  {32'hc00b33b6, 32'hc0f4ccd2} /* (2, 6, 28) {real, imag} */,
  {32'hbf984b58, 32'hc10d2ea4} /* (2, 6, 27) {real, imag} */,
  {32'hc0a2be58, 32'hc13418d9} /* (2, 6, 26) {real, imag} */,
  {32'hc0cd8538, 32'hc186aeee} /* (2, 6, 25) {real, imag} */,
  {32'hc119bd81, 32'hc0b908ee} /* (2, 6, 24) {real, imag} */,
  {32'hc10c5ec8, 32'hc1a8aa16} /* (2, 6, 23) {real, imag} */,
  {32'hc186b752, 32'hc126de52} /* (2, 6, 22) {real, imag} */,
  {32'hc1963fe2, 32'h40e816f0} /* (2, 6, 21) {real, imag} */,
  {32'hc182c73c, 32'h41390940} /* (2, 6, 20) {real, imag} */,
  {32'h408e2e5d, 32'h40c4fdb7} /* (2, 6, 19) {real, imag} */,
  {32'hbe7a23c0, 32'h409f181c} /* (2, 6, 18) {real, imag} */,
  {32'h3ec52fd0, 32'h418193fc} /* (2, 6, 17) {real, imag} */,
  {32'hc131b39a, 32'h41503e12} /* (2, 6, 16) {real, imag} */,
  {32'hc15f4775, 32'h4156fbf8} /* (2, 6, 15) {real, imag} */,
  {32'h40d43f27, 32'hc09544fe} /* (2, 6, 14) {real, imag} */,
  {32'hc000e556, 32'hc1d6b9d4} /* (2, 6, 13) {real, imag} */,
  {32'hc16b9d50, 32'hc0c1a208} /* (2, 6, 12) {real, imag} */,
  {32'h3f6c654c, 32'hc0f646c4} /* (2, 6, 11) {real, imag} */,
  {32'h4110afd7, 32'hc187b004} /* (2, 6, 10) {real, imag} */,
  {32'h3f21dc80, 32'hc0a0f250} /* (2, 6, 9) {real, imag} */,
  {32'hc0410148, 32'hbeac1480} /* (2, 6, 8) {real, imag} */,
  {32'h41058fca, 32'hc0d2d540} /* (2, 6, 7) {real, imag} */,
  {32'h3f92b25c, 32'hc1182ff3} /* (2, 6, 6) {real, imag} */,
  {32'hc025a611, 32'hc0c0674e} /* (2, 6, 5) {real, imag} */,
  {32'h4118ee64, 32'hbf0b27d8} /* (2, 6, 4) {real, imag} */,
  {32'h40b618b8, 32'hc0194cd8} /* (2, 6, 3) {real, imag} */,
  {32'hc0acc60f, 32'h4088ad24} /* (2, 6, 2) {real, imag} */,
  {32'hc0d235ee, 32'h419061d0} /* (2, 6, 1) {real, imag} */,
  {32'hc1147e9a, 32'h4186b8fc} /* (2, 6, 0) {real, imag} */,
  {32'h41729ebf, 32'hc1ed9571} /* (2, 5, 31) {real, imag} */,
  {32'h421ef14c, 32'hc281a0db} /* (2, 5, 30) {real, imag} */,
  {32'h41de48bd, 32'hc27365ea} /* (2, 5, 29) {real, imag} */,
  {32'h420aa974, 32'hc28f962f} /* (2, 5, 28) {real, imag} */,
  {32'h41cc0ee0, 32'hc25bf9ef} /* (2, 5, 27) {real, imag} */,
  {32'h41bc4b10, 32'hc1f0b091} /* (2, 5, 26) {real, imag} */,
  {32'h416f2180, 32'hc12fe088} /* (2, 5, 25) {real, imag} */,
  {32'h420f83a0, 32'hc1b01644} /* (2, 5, 24) {real, imag} */,
  {32'h423db920, 32'hc205f333} /* (2, 5, 23) {real, imag} */,
  {32'h41ebc59e, 32'hc281a7a8} /* (2, 5, 22) {real, imag} */,
  {32'h4187e8e4, 32'hc21467b3} /* (2, 5, 21) {real, imag} */,
  {32'hc0eef475, 32'h41ecec48} /* (2, 5, 20) {real, imag} */,
  {32'hc18ef0a6, 32'h42590142} /* (2, 5, 19) {real, imag} */,
  {32'hc139c97e, 32'h4240c42c} /* (2, 5, 18) {real, imag} */,
  {32'hc10d6e4a, 32'h41740c17} /* (2, 5, 17) {real, imag} */,
  {32'hc1829f12, 32'h4102d4f2} /* (2, 5, 16) {real, imag} */,
  {32'hc2055203, 32'h41688834} /* (2, 5, 15) {real, imag} */,
  {32'hc1f80be1, 32'h41b43ade} /* (2, 5, 14) {real, imag} */,
  {32'hc195ff86, 32'h4200185e} /* (2, 5, 13) {real, imag} */,
  {32'hc1afa5fe, 32'h42544fd4} /* (2, 5, 12) {real, imag} */,
  {32'hc1a00e73, 32'h42461752} /* (2, 5, 11) {real, imag} */,
  {32'h414a3fd7, 32'hc15096cc} /* (2, 5, 10) {real, imag} */,
  {32'h3eab2830, 32'hc2232f6c} /* (2, 5, 9) {real, imag} */,
  {32'hc11ef188, 32'hc1f2476e} /* (2, 5, 8) {real, imag} */,
  {32'h41a44b72, 32'hc25250cd} /* (2, 5, 7) {real, imag} */,
  {32'h4125ee6f, 32'hc1dcaef8} /* (2, 5, 6) {real, imag} */,
  {32'h41ba8a55, 32'hc1f25fa7} /* (2, 5, 5) {real, imag} */,
  {32'h422095be, 32'hc20a2c3d} /* (2, 5, 4) {real, imag} */,
  {32'h421e8f9a, 32'hc2260d3e} /* (2, 5, 3) {real, imag} */,
  {32'h421c0633, 32'hc271e1de} /* (2, 5, 2) {real, imag} */,
  {32'h422884f3, 32'hc26a0bdb} /* (2, 5, 1) {real, imag} */,
  {32'h418cf626, 32'hc1a9102f} /* (2, 5, 0) {real, imag} */,
  {32'hc02794ad, 32'h415a4f89} /* (2, 4, 31) {real, imag} */,
  {32'h40b55f90, 32'h41914773} /* (2, 4, 30) {real, imag} */,
  {32'h40c02283, 32'h41a0b084} /* (2, 4, 29) {real, imag} */,
  {32'hc055d921, 32'h42001de0} /* (2, 4, 28) {real, imag} */,
  {32'hc0922e4b, 32'h41815338} /* (2, 4, 27) {real, imag} */,
  {32'hc18afa2f, 32'h4195e9ea} /* (2, 4, 26) {real, imag} */,
  {32'hc1d55dbb, 32'h42237dc3} /* (2, 4, 25) {real, imag} */,
  {32'hc182e186, 32'h41f89dd2} /* (2, 4, 24) {real, imag} */,
  {32'hc1473c00, 32'h41c824c6} /* (2, 4, 23) {real, imag} */,
  {32'hc0bbf98a, 32'h4240229e} /* (2, 4, 22) {real, imag} */,
  {32'h3f9cc4da, 32'hc00dbc5c} /* (2, 4, 21) {real, imag} */,
  {32'h4257b2dc, 32'hc23ff75c} /* (2, 4, 20) {real, imag} */,
  {32'h42a7d2fc, 32'hc2403a24} /* (2, 4, 19) {real, imag} */,
  {32'h429c86cd, 32'hc240e0ec} /* (2, 4, 18) {real, imag} */,
  {32'h429ba9c2, 32'hc2621882} /* (2, 4, 17) {real, imag} */,
  {32'h428b7ad8, 32'hc241ac54} /* (2, 4, 16) {real, imag} */,
  {32'h418074b8, 32'hc21d5ca0} /* (2, 4, 15) {real, imag} */,
  {32'h41dfff8a, 32'hc2362060} /* (2, 4, 14) {real, imag} */,
  {32'h41db0d11, 32'hc2280d18} /* (2, 4, 13) {real, imag} */,
  {32'h4192532d, 32'hc233b258} /* (2, 4, 12) {real, imag} */,
  {32'h41210274, 32'hc1f0866e} /* (2, 4, 11) {real, imag} */,
  {32'hc24e6b06, 32'h417b25e2} /* (2, 4, 10) {real, imag} */,
  {32'hc2a1a9ea, 32'h42481ae0} /* (2, 4, 9) {real, imag} */,
  {32'hc26e54cc, 32'h4249537c} /* (2, 4, 8) {real, imag} */,
  {32'hc281c138, 32'h4281ccfa} /* (2, 4, 7) {real, imag} */,
  {32'hc2a26870, 32'h42298116} /* (2, 4, 6) {real, imag} */,
  {32'hc241d8ca, 32'h420ac9e1} /* (2, 4, 5) {real, imag} */,
  {32'hc20920d9, 32'h416c4e45} /* (2, 4, 4) {real, imag} */,
  {32'hc1bc31f2, 32'h413b0158} /* (2, 4, 3) {real, imag} */,
  {32'hc173725c, 32'h41d7060e} /* (2, 4, 2) {real, imag} */,
  {32'hc1a9c0ae, 32'h425ad3d6} /* (2, 4, 1) {real, imag} */,
  {32'hc10aea1d, 32'h41d3b3e7} /* (2, 4, 0) {real, imag} */,
  {32'hc0b00f34, 32'hbf248398} /* (2, 3, 31) {real, imag} */,
  {32'hbe97bae0, 32'h41075c64} /* (2, 3, 30) {real, imag} */,
  {32'h411ba2d2, 32'hc1476305} /* (2, 3, 29) {real, imag} */,
  {32'hc1391ec5, 32'hc1a647b6} /* (2, 3, 28) {real, imag} */,
  {32'hc1c725c4, 32'hc16ab6c8} /* (2, 3, 27) {real, imag} */,
  {32'hc1fa4780, 32'hc08dad8f} /* (2, 3, 26) {real, imag} */,
  {32'hc1298258, 32'hc1579ab5} /* (2, 3, 25) {real, imag} */,
  {32'h40cca29a, 32'hbfeb7868} /* (2, 3, 24) {real, imag} */,
  {32'h41b71980, 32'h412f886c} /* (2, 3, 23) {real, imag} */,
  {32'hc0db25a4, 32'hc16f2c24} /* (2, 3, 22) {real, imag} */,
  {32'h40bd19ac, 32'hc19fd47a} /* (2, 3, 21) {real, imag} */,
  {32'h428195ee, 32'hbd2c4640} /* (2, 3, 20) {real, imag} */,
  {32'h42b9dabb, 32'h41f7a2ca} /* (2, 3, 19) {real, imag} */,
  {32'h4298eff0, 32'h425e90fc} /* (2, 3, 18) {real, imag} */,
  {32'h42bcf8dc, 32'h4269786d} /* (2, 3, 17) {real, imag} */,
  {32'h4284f476, 32'h4212f5a6} /* (2, 3, 16) {real, imag} */,
  {32'h40d16338, 32'h4191de81} /* (2, 3, 15) {real, imag} */,
  {32'hc11e8df8, 32'h41ca30b2} /* (2, 3, 14) {real, imag} */,
  {32'hc0c49757, 32'h3f5241a8} /* (2, 3, 13) {real, imag} */,
  {32'hc0e25b50, 32'hc1607383} /* (2, 3, 12) {real, imag} */,
  {32'hc1a3ec74, 32'hc178e44a} /* (2, 3, 11) {real, imag} */,
  {32'hc297594d, 32'hc1ab4f9b} /* (2, 3, 10) {real, imag} */,
  {32'hc2b6e1eb, 32'hc1e2e10c} /* (2, 3, 9) {real, imag} */,
  {32'hc2a2831b, 32'hc1cc9b21} /* (2, 3, 8) {real, imag} */,
  {32'hc2a58fa1, 32'hc2160f93} /* (2, 3, 7) {real, imag} */,
  {32'hc2a6713d, 32'hc22fca81} /* (2, 3, 6) {real, imag} */,
  {32'hc0eb9de4, 32'hc183b707} /* (2, 3, 5) {real, imag} */,
  {32'h415ec089, 32'h3dfbdb00} /* (2, 3, 4) {real, imag} */,
  {32'h40661c2d, 32'hc023c9da} /* (2, 3, 3) {real, imag} */,
  {32'h41bcc45a, 32'hc0cc843f} /* (2, 3, 2) {real, imag} */,
  {32'h4136c774, 32'h41b7f559} /* (2, 3, 1) {real, imag} */,
  {32'hc1017423, 32'h4146fe19} /* (2, 3, 0) {real, imag} */,
  {32'h41c7c26c, 32'hc2ab25eb} /* (2, 2, 31) {real, imag} */,
  {32'h42450fdc, 32'hc30b2c4c} /* (2, 2, 30) {real, imag} */,
  {32'h426416a1, 32'hc3106abd} /* (2, 2, 29) {real, imag} */,
  {32'h4256483c, 32'hc311260e} /* (2, 2, 28) {real, imag} */,
  {32'h426625fe, 32'hc2f2adec} /* (2, 2, 27) {real, imag} */,
  {32'h42816e0e, 32'hc2de7070} /* (2, 2, 26) {real, imag} */,
  {32'h41cba4ac, 32'hc2e1b261} /* (2, 2, 25) {real, imag} */,
  {32'h41ea2ceb, 32'hc3176ae0} /* (2, 2, 24) {real, imag} */,
  {32'h42362e27, 32'hc3165076} /* (2, 2, 23) {real, imag} */,
  {32'h4270f4ac, 32'hc30b881f} /* (2, 2, 22) {real, imag} */,
  {32'h427fff10, 32'hc1ed41e0} /* (2, 2, 21) {real, imag} */,
  {32'h423fcb66, 32'h433c2582} /* (2, 2, 20) {real, imag} */,
  {32'h41875dfc, 32'h437107c4} /* (2, 2, 19) {real, imag} */,
  {32'h419abbe6, 32'h4379c95e} /* (2, 2, 18) {real, imag} */,
  {32'h419b0a1a, 32'h437327b2} /* (2, 2, 17) {real, imag} */,
  {32'h41d530ba, 32'h4352a4ad} /* (2, 2, 16) {real, imag} */,
  {32'hc15aa462, 32'h43298523} /* (2, 2, 15) {real, imag} */,
  {32'hc25d990e, 32'h43072567} /* (2, 2, 14) {real, imag} */,
  {32'hc24c838a, 32'h42d62f81} /* (2, 2, 13) {real, imag} */,
  {32'hc2034b30, 32'h43092818} /* (2, 2, 12) {real, imag} */,
  {32'hc22ba564, 32'h42ebe2de} /* (2, 2, 11) {real, imag} */,
  {32'hc1cd99d8, 32'hc2be6a2b} /* (2, 2, 10) {real, imag} */,
  {32'hc1867300, 32'hc3566cb3} /* (2, 2, 9) {real, imag} */,
  {32'hc18cd8ac, 32'hc375608e} /* (2, 2, 8) {real, imag} */,
  {32'hc1d15670, 32'hc36ec957} /* (2, 2, 7) {real, imag} */,
  {32'hc26ea2ad, 32'hc3505636} /* (2, 2, 6) {real, imag} */,
  {32'hc1e2b9c7, 32'hc32d8b79} /* (2, 2, 5) {real, imag} */,
  {32'h41b986b2, 32'hc320c630} /* (2, 2, 4) {real, imag} */,
  {32'h427a3594, 32'hc30af98a} /* (2, 2, 3) {real, imag} */,
  {32'h42984f2a, 32'hc3017814} /* (2, 2, 2) {real, imag} */,
  {32'h429a42e4, 32'hc2f4d5ca} /* (2, 2, 1) {real, imag} */,
  {32'h41d8d49e, 32'hc2a9b5a1} /* (2, 2, 0) {real, imag} */,
  {32'hc2147d98, 32'h42f086b3} /* (2, 1, 31) {real, imag} */,
  {32'hc29ac48c, 32'h436cda73} /* (2, 1, 30) {real, imag} */,
  {32'hc28b6680, 32'h436f9c29} /* (2, 1, 29) {real, imag} */,
  {32'hc285b8a6, 32'h43617a91} /* (2, 1, 28) {real, imag} */,
  {32'hc24a2efb, 32'h4368b315} /* (2, 1, 27) {real, imag} */,
  {32'hc22f865f, 32'h435ee4f6} /* (2, 1, 26) {real, imag} */,
  {32'hc2894b27, 32'h4372acf0} /* (2, 1, 25) {real, imag} */,
  {32'hc290e5e1, 32'h437c4021} /* (2, 1, 24) {real, imag} */,
  {32'hc2992670, 32'h4382bd82} /* (2, 1, 23) {real, imag} */,
  {32'hc2a2e42c, 32'h437d7331} /* (2, 1, 22) {real, imag} */,
  {32'h3fc66cf0, 32'h430cbe91} /* (2, 1, 21) {real, imag} */,
  {32'h42e974ee, 32'hc16c869c} /* (2, 1, 20) {real, imag} */,
  {32'h42ebafd5, 32'hc28cf800} /* (2, 1, 19) {real, imag} */,
  {32'h42a5fa56, 32'hc2bc8306} /* (2, 1, 18) {real, imag} */,
  {32'h42e083fa, 32'hc2c00546} /* (2, 1, 17) {real, imag} */,
  {32'h42e4f01e, 32'hc30eea9f} /* (2, 1, 16) {real, imag} */,
  {32'h42a1ee87, 32'hc35776e9} /* (2, 1, 15) {real, imag} */,
  {32'h42b77544, 32'hc35e4733} /* (2, 1, 14) {real, imag} */,
  {32'h42b42b4a, 32'hc36a7259} /* (2, 1, 13) {real, imag} */,
  {32'h42849470, 32'hc36f6558} /* (2, 1, 12) {real, imag} */,
  {32'h41f2134b, 32'hc347866f} /* (2, 1, 11) {real, imag} */,
  {32'hc2a6115b, 32'hc17580c6} /* (2, 1, 10) {real, imag} */,
  {32'hc30ae754, 32'h429eb7fe} /* (2, 1, 9) {real, imag} */,
  {32'hc318cb3d, 32'h42ba2547} /* (2, 1, 8) {real, imag} */,
  {32'hc305d7ea, 32'h42b4fe3b} /* (2, 1, 7) {real, imag} */,
  {32'hc2b60a20, 32'h42a267aa} /* (2, 1, 6) {real, imag} */,
  {32'hc2716cce, 32'h433726b8} /* (2, 1, 5) {real, imag} */,
  {32'hc283a34e, 32'h43628c53} /* (2, 1, 4) {real, imag} */,
  {32'hc2a93c34, 32'h435a285e} /* (2, 1, 3) {real, imag} */,
  {32'hc2bd9034, 32'h4351ea00} /* (2, 1, 2) {real, imag} */,
  {32'hc2b6aeb8, 32'h43526344} /* (2, 1, 1) {real, imag} */,
  {32'hc250013c, 32'h43020bbe} /* (2, 1, 0) {real, imag} */,
  {32'hc20a9050, 32'h4295c748} /* (2, 0, 31) {real, imag} */,
  {32'hc1c417e4, 32'h42ff62f4} /* (2, 0, 30) {real, imag} */,
  {32'hc189d400, 32'h43188fb7} /* (2, 0, 29) {real, imag} */,
  {32'hc1cde45c, 32'h4309c693} /* (2, 0, 28) {real, imag} */,
  {32'hc21da660, 32'h431c51fa} /* (2, 0, 27) {real, imag} */,
  {32'hc1fd430a, 32'h432c2c34} /* (2, 0, 26) {real, imag} */,
  {32'hc131bd66, 32'h43220fc1} /* (2, 0, 25) {real, imag} */,
  {32'hc1a8f3d7, 32'h4325a230} /* (2, 0, 24) {real, imag} */,
  {32'hc250d411, 32'h43146364} /* (2, 0, 23) {real, imag} */,
  {32'hc208b272, 32'h430b9da4} /* (2, 0, 22) {real, imag} */,
  {32'hc17eba7f, 32'h42f5a33a} /* (2, 0, 21) {real, imag} */,
  {32'h40b1c618, 32'h4210da3e} /* (2, 0, 20) {real, imag} */,
  {32'h4171b1e7, 32'h40e67e0e} /* (2, 0, 19) {real, imag} */,
  {32'hc18e002c, 32'h40bb60d6} /* (2, 0, 18) {real, imag} */,
  {32'hc1650fd8, 32'h419e04b2} /* (2, 0, 17) {real, imag} */,
  {32'h40169cfa, 32'hc1f5e61e} /* (2, 0, 16) {real, imag} */,
  {32'h416367ec, 32'hc30585c0} /* (2, 0, 15) {real, imag} */,
  {32'h41815e08, 32'hc322467c} /* (2, 0, 14) {real, imag} */,
  {32'h41e890ea, 32'hc3080118} /* (2, 0, 13) {real, imag} */,
  {32'h422a3708, 32'hc312a848} /* (2, 0, 12) {real, imag} */,
  {32'h425d8a60, 32'hc304be7c} /* (2, 0, 11) {real, imag} */,
  {32'h3b405800, 32'hc2728c2e} /* (2, 0, 10) {real, imag} */,
  {32'hc09a0322, 32'h4198e6fe} /* (2, 0, 9) {real, imag} */,
  {32'h406a8df4, 32'h4152b42b} /* (2, 0, 8) {real, imag} */,
  {32'hc17a3018, 32'hc17cbf90} /* (2, 0, 7) {real, imag} */,
  {32'hc0c9702a, 32'h4078b77a} /* (2, 0, 6) {real, imag} */,
  {32'hc1ed324a, 32'h42ba09a9} /* (2, 0, 5) {real, imag} */,
  {32'hc22a992e, 32'h4326c21e} /* (2, 0, 4) {real, imag} */,
  {32'hc1189c0d, 32'h43240dfb} /* (2, 0, 3) {real, imag} */,
  {32'hc1d5932c, 32'h4321481e} /* (2, 0, 2) {real, imag} */,
  {32'hc2241018, 32'h42f3d462} /* (2, 0, 1) {real, imag} */,
  {32'hc1f3f8bc, 32'h4289b18f} /* (2, 0, 0) {real, imag} */,
  {32'h40fe3a1e, 32'hc287bfe2} /* (1, 31, 31) {real, imag} */,
  {32'hc102f266, 32'hc2ff857e} /* (1, 31, 30) {real, imag} */,
  {32'hc0966826, 32'hc2e6925d} /* (1, 31, 29) {real, imag} */,
  {32'hc1bdb205, 32'hc3051dff} /* (1, 31, 28) {real, imag} */,
  {32'hbff75238, 32'hc31a7bed} /* (1, 31, 27) {real, imag} */,
  {32'hc13d6bb6, 32'hc3144a15} /* (1, 31, 26) {real, imag} */,
  {32'hc162884e, 32'hc30198fd} /* (1, 31, 25) {real, imag} */,
  {32'h411619c0, 32'hc321730e} /* (1, 31, 24) {real, imag} */,
  {32'hc09617be, 32'hc31b6b24} /* (1, 31, 23) {real, imag} */,
  {32'h4030c6c1, 32'hc3061403} /* (1, 31, 22) {real, imag} */,
  {32'h4220d41b, 32'hc2867dce} /* (1, 31, 21) {real, imag} */,
  {32'h424787ee, 32'h423fb45f} /* (1, 31, 20) {real, imag} */,
  {32'h4254d24b, 32'h426628ee} /* (1, 31, 19) {real, imag} */,
  {32'h42467def, 32'h4257f18f} /* (1, 31, 18) {real, imag} */,
  {32'h4275313d, 32'h421b92d1} /* (1, 31, 17) {real, imag} */,
  {32'h41dcd60e, 32'h4286046b} /* (1, 31, 16) {real, imag} */,
  {32'hc1a223cc, 32'h430143e6} /* (1, 31, 15) {real, imag} */,
  {32'hc1c9d95a, 32'h430d372c} /* (1, 31, 14) {real, imag} */,
  {32'hbda77700, 32'h42f22098} /* (1, 31, 13) {real, imag} */,
  {32'h411a68d4, 32'h430419c0} /* (1, 31, 12) {real, imag} */,
  {32'hc17be537, 32'h42b37d18} /* (1, 31, 11) {real, imag} */,
  {32'hc27136b6, 32'hc2068a5b} /* (1, 31, 10) {real, imag} */,
  {32'hc239fc61, 32'hc25fec9c} /* (1, 31, 9) {real, imag} */,
  {32'hc1b7e968, 32'hc28fdc39} /* (1, 31, 8) {real, imag} */,
  {32'hc2720c48, 32'hc292e94e} /* (1, 31, 7) {real, imag} */,
  {32'hc2733e16, 32'hc2978d5f} /* (1, 31, 6) {real, imag} */,
  {32'hc1ea5f0b, 32'hc2bc78b4} /* (1, 31, 5) {real, imag} */,
  {32'hc0f8406c, 32'hc2f10d4a} /* (1, 31, 4) {real, imag} */,
  {32'h41c6d9e8, 32'hc30e05ee} /* (1, 31, 3) {real, imag} */,
  {32'h41cd6e86, 32'hc30ca99f} /* (1, 31, 2) {real, imag} */,
  {32'h41122bee, 32'hc310d6de} /* (1, 31, 1) {real, imag} */,
  {32'h403e2692, 32'hc287f0f0} /* (1, 31, 0) {real, imag} */,
  {32'hc1555b7d, 32'h41efb520} /* (1, 30, 31) {real, imag} */,
  {32'hc1026304, 32'h42a5249a} /* (1, 30, 30) {real, imag} */,
  {32'h40106bb0, 32'h42c32d6b} /* (1, 30, 29) {real, imag} */,
  {32'h421667cc, 32'h42a9fa5e} /* (1, 30, 28) {real, imag} */,
  {32'h41d9e4a3, 32'h428c31c6} /* (1, 30, 27) {real, imag} */,
  {32'h40446620, 32'h4290ace2} /* (1, 30, 26) {real, imag} */,
  {32'h402fe302, 32'h42a7bfc5} /* (1, 30, 25) {real, imag} */,
  {32'h40646630, 32'h4276c3cc} /* (1, 30, 24) {real, imag} */,
  {32'h408ba4f0, 32'h42b1ba64} /* (1, 30, 23) {real, imag} */,
  {32'h40ff1ede, 32'h42d44bcc} /* (1, 30, 22) {real, imag} */,
  {32'h40109200, 32'h422733ca} /* (1, 30, 21) {real, imag} */,
  {32'h42195c26, 32'hc28d8a43} /* (1, 30, 20) {real, imag} */,
  {32'h426faa49, 32'hc2ec1404} /* (1, 30, 19) {real, imag} */,
  {32'h4285246f, 32'hc2cb2923} /* (1, 30, 18) {real, imag} */,
  {32'h42882762, 32'hc2d040ee} /* (1, 30, 17) {real, imag} */,
  {32'h4250cdac, 32'hc2f11320} /* (1, 30, 16) {real, imag} */,
  {32'h41aaedba, 32'hc2bd929c} /* (1, 30, 15) {real, imag} */,
  {32'h4171229a, 32'hc2a16479} /* (1, 30, 14) {real, imag} */,
  {32'h3de20300, 32'hc2986552} /* (1, 30, 13) {real, imag} */,
  {32'hc1fc7664, 32'hc292c45d} /* (1, 30, 12) {real, imag} */,
  {32'hc20531dd, 32'hc2110db5} /* (1, 30, 11) {real, imag} */,
  {32'hc22ec43e, 32'h42888c4c} /* (1, 30, 10) {real, imag} */,
  {32'hc2819f3b, 32'h42de442b} /* (1, 30, 9) {real, imag} */,
  {32'hc28a1aaa, 32'h42d347b0} /* (1, 30, 8) {real, imag} */,
  {32'hc24ba52b, 32'h42f1901c} /* (1, 30, 7) {real, imag} */,
  {32'hc20933b8, 32'h42e38978} /* (1, 30, 6) {real, imag} */,
  {32'hc120f5a0, 32'h42ca3610} /* (1, 30, 5) {real, imag} */,
  {32'hc11f66b2, 32'h42b29997} /* (1, 30, 4) {real, imag} */,
  {32'hc09065f6, 32'h42c4c7f6} /* (1, 30, 3) {real, imag} */,
  {32'h407d080c, 32'h42b7ad94} /* (1, 30, 2) {real, imag} */,
  {32'hc0abc1be, 32'h429feeb7} /* (1, 30, 1) {real, imag} */,
  {32'hc0218c68, 32'h421d1689} /* (1, 30, 0) {real, imag} */,
  {32'hc0bf43be, 32'hc07d8cfa} /* (1, 29, 31) {real, imag} */,
  {32'h403495d2, 32'hc17131c0} /* (1, 29, 30) {real, imag} */,
  {32'h416435e5, 32'hc1cad6c2} /* (1, 29, 29) {real, imag} */,
  {32'h40b14360, 32'hc1c755db} /* (1, 29, 28) {real, imag} */,
  {32'h4105b56c, 32'hc1214b18} /* (1, 29, 27) {real, imag} */,
  {32'hbf1d7464, 32'h41347230} /* (1, 29, 26) {real, imag} */,
  {32'h41aa2333, 32'hc19d4076} /* (1, 29, 25) {real, imag} */,
  {32'h414ce73c, 32'hc081866f} /* (1, 29, 24) {real, imag} */,
  {32'h40c106ca, 32'h414c546f} /* (1, 29, 23) {real, imag} */,
  {32'h3e36da80, 32'h41c77194} /* (1, 29, 22) {real, imag} */,
  {32'h40f32101, 32'h41d62784} /* (1, 29, 21) {real, imag} */,
  {32'h42085917, 32'h41bf0e20} /* (1, 29, 20) {real, imag} */,
  {32'h4200affc, 32'h40e5bbcb} /* (1, 29, 19) {real, imag} */,
  {32'h42816137, 32'h4160f246} /* (1, 29, 18) {real, imag} */,
  {32'h42517a2c, 32'h41197b03} /* (1, 29, 17) {real, imag} */,
  {32'h42023acc, 32'hc106946d} /* (1, 29, 16) {real, imag} */,
  {32'h4111983e, 32'hc0a1e3f0} /* (1, 29, 15) {real, imag} */,
  {32'h4116a37f, 32'h41864337} /* (1, 29, 14) {real, imag} */,
  {32'h419af319, 32'h41ea4759} /* (1, 29, 13) {real, imag} */,
  {32'hc165bfe5, 32'h41171d78} /* (1, 29, 12) {real, imag} */,
  {32'h40ad8ee4, 32'hc047107c} /* (1, 29, 11) {real, imag} */,
  {32'hc093eaf4, 32'h40835668} /* (1, 29, 10) {real, imag} */,
  {32'hc20f94d0, 32'hc0521108} /* (1, 29, 9) {real, imag} */,
  {32'hc2911657, 32'h3fa41eb0} /* (1, 29, 8) {real, imag} */,
  {32'hc280653d, 32'hc03bf572} /* (1, 29, 7) {real, imag} */,
  {32'hc2679371, 32'h4137049e} /* (1, 29, 6) {real, imag} */,
  {32'hc236eee4, 32'h40727c6c} /* (1, 29, 5) {real, imag} */,
  {32'h401e0aff, 32'h40663aec} /* (1, 29, 4) {real, imag} */,
  {32'h4025f814, 32'hc0d3aeb2} /* (1, 29, 3) {real, imag} */,
  {32'hbf1ad6d0, 32'h413e5b40} /* (1, 29, 2) {real, imag} */,
  {32'hbf6227e4, 32'h41290e4a} /* (1, 29, 1) {real, imag} */,
  {32'hc0635a77, 32'h3fd56966} /* (1, 29, 0) {real, imag} */,
  {32'hc0cc0e2f, 32'hc0fe323f} /* (1, 28, 31) {real, imag} */,
  {32'hc1aa9fd1, 32'hc1988e32} /* (1, 28, 30) {real, imag} */,
  {32'hc18b6b26, 32'hc22bbbe6} /* (1, 28, 29) {real, imag} */,
  {32'hc13f6e40, 32'hc22ee641} /* (1, 28, 28) {real, imag} */,
  {32'h419bc289, 32'hc1c08d2e} /* (1, 28, 27) {real, imag} */,
  {32'h41dbc56e, 32'hc1892f84} /* (1, 28, 26) {real, imag} */,
  {32'h4120a4bc, 32'hc197ce8e} /* (1, 28, 25) {real, imag} */,
  {32'hc1a7e313, 32'hc148b60f} /* (1, 28, 24) {real, imag} */,
  {32'hbecdf200, 32'hc1d8320e} /* (1, 28, 23) {real, imag} */,
  {32'h403c3578, 32'hc1aa8687} /* (1, 28, 22) {real, imag} */,
  {32'h414ec89b, 32'hc1bcc99a} /* (1, 28, 21) {real, imag} */,
  {32'h42666fce, 32'h419a728c} /* (1, 28, 20) {real, imag} */,
  {32'h423200f0, 32'h422a37cc} /* (1, 28, 19) {real, imag} */,
  {32'h424a53ed, 32'h4207da6c} /* (1, 28, 18) {real, imag} */,
  {32'h422a4b40, 32'h4256c69b} /* (1, 28, 17) {real, imag} */,
  {32'h42019c46, 32'h4246c6b6} /* (1, 28, 16) {real, imag} */,
  {32'h420c87fb, 32'h419a3233} /* (1, 28, 15) {real, imag} */,
  {32'h41cc84fb, 32'h416a43de} /* (1, 28, 14) {real, imag} */,
  {32'h416d2a71, 32'h41d42987} /* (1, 28, 13) {real, imag} */,
  {32'h41bbee7b, 32'h41310cb1} /* (1, 28, 12) {real, imag} */,
  {32'h40bf2ea0, 32'h40f5d2ce} /* (1, 28, 11) {real, imag} */,
  {32'hc1c09086, 32'hc1922510} /* (1, 28, 10) {real, imag} */,
  {32'hc14e930d, 32'hc2265950} /* (1, 28, 9) {real, imag} */,
  {32'hc2087aea, 32'hc2450105} /* (1, 28, 8) {real, imag} */,
  {32'hc2259125, 32'hc231abbe} /* (1, 28, 7) {real, imag} */,
  {32'hc1d12ec4, 32'hc238acf7} /* (1, 28, 6) {real, imag} */,
  {32'hc17dbbdd, 32'hc1cbdfab} /* (1, 28, 5) {real, imag} */,
  {32'h40f8d6ee, 32'hc15402c4} /* (1, 28, 4) {real, imag} */,
  {32'h41156b42, 32'hc1995292} /* (1, 28, 3) {real, imag} */,
  {32'hc116dbd8, 32'hc1cd425c} /* (1, 28, 2) {real, imag} */,
  {32'hc16ee546, 32'hc1cad78a} /* (1, 28, 1) {real, imag} */,
  {32'h4090c686, 32'hc1a9a3b0} /* (1, 28, 0) {real, imag} */,
  {32'h416ffafc, 32'h41d6f485} /* (1, 27, 31) {real, imag} */,
  {32'h4196caac, 32'h422007bb} /* (1, 27, 30) {real, imag} */,
  {32'h421198a8, 32'h41bb9812} /* (1, 27, 29) {real, imag} */,
  {32'h4205e088, 32'h41a020f7} /* (1, 27, 28) {real, imag} */,
  {32'h41b57afb, 32'h41f99c45} /* (1, 27, 27) {real, imag} */,
  {32'h4193f14c, 32'h41bc5a88} /* (1, 27, 26) {real, imag} */,
  {32'h41f58eb3, 32'h41edf584} /* (1, 27, 25) {real, imag} */,
  {32'h422c6785, 32'h41f30c62} /* (1, 27, 24) {real, imag} */,
  {32'h417f1560, 32'h42375c31} /* (1, 27, 23) {real, imag} */,
  {32'h3f151c50, 32'h4244cfe2} /* (1, 27, 22) {real, imag} */,
  {32'h416c88a8, 32'h42169267} /* (1, 27, 21) {real, imag} */,
  {32'h4147cd09, 32'h3deb4820} /* (1, 27, 20) {real, imag} */,
  {32'hc0448176, 32'hc0e23c03} /* (1, 27, 19) {real, imag} */,
  {32'hc0a14ca6, 32'hc18071ba} /* (1, 27, 18) {real, imag} */,
  {32'h3fbdb540, 32'hc194b069} /* (1, 27, 17) {real, imag} */,
  {32'h414fd9c1, 32'hc1dfcf78} /* (1, 27, 16) {real, imag} */,
  {32'h403fbf48, 32'hc246a5dd} /* (1, 27, 15) {real, imag} */,
  {32'hc0baaf58, 32'hc2061fac} /* (1, 27, 14) {real, imag} */,
  {32'hc0d49594, 32'hc1de3f04} /* (1, 27, 13) {real, imag} */,
  {32'hc1b3eb89, 32'hc1f3596b} /* (1, 27, 12) {real, imag} */,
  {32'hc1c27943, 32'hc1d21e5b} /* (1, 27, 11) {real, imag} */,
  {32'h414cb812, 32'hbdef7980} /* (1, 27, 10) {real, imag} */,
  {32'h40fee3f2, 32'h416de018} /* (1, 27, 9) {real, imag} */,
  {32'h40b5a96c, 32'h408d5988} /* (1, 27, 8) {real, imag} */,
  {32'h414ef312, 32'h4022b75a} /* (1, 27, 7) {real, imag} */,
  {32'h40d95d4f, 32'h40fdbf13} /* (1, 27, 6) {real, imag} */,
  {32'h41a2b97a, 32'h4190b10c} /* (1, 27, 5) {real, imag} */,
  {32'h405f07c8, 32'h41c75136} /* (1, 27, 4) {real, imag} */,
  {32'hc130bf10, 32'h41750e58} /* (1, 27, 3) {real, imag} */,
  {32'h4137f6d6, 32'h41afc943} /* (1, 27, 2) {real, imag} */,
  {32'h40d4a6e8, 32'h4242994b} /* (1, 27, 1) {real, imag} */,
  {32'hc083c717, 32'h4213d4fe} /* (1, 27, 0) {real, imag} */,
  {32'hc0ef901e, 32'hc0bb0c70} /* (1, 26, 31) {real, imag} */,
  {32'hc1e28df0, 32'hbf159670} /* (1, 26, 30) {real, imag} */,
  {32'hc1a4b393, 32'hc0d93fb3} /* (1, 26, 29) {real, imag} */,
  {32'hc16cec8c, 32'hc103a0d9} /* (1, 26, 28) {real, imag} */,
  {32'hc1e34616, 32'hc1efdb06} /* (1, 26, 27) {real, imag} */,
  {32'hc0d802f0, 32'hc1a06230} /* (1, 26, 26) {real, imag} */,
  {32'h3e276100, 32'h40c1b9b7} /* (1, 26, 25) {real, imag} */,
  {32'h411b9b81, 32'h41f20691} /* (1, 26, 24) {real, imag} */,
  {32'h41919cee, 32'h4108decb} /* (1, 26, 23) {real, imag} */,
  {32'h40213cb6, 32'h418e999e} /* (1, 26, 22) {real, imag} */,
  {32'hc0c8b210, 32'h3fffb480} /* (1, 26, 21) {real, imag} */,
  {32'h40a24012, 32'hc1814ffc} /* (1, 26, 20) {real, imag} */,
  {32'h4175c0d3, 32'hc092cb42} /* (1, 26, 19) {real, imag} */,
  {32'h411c2c13, 32'h40a4cc1e} /* (1, 26, 18) {real, imag} */,
  {32'h404b0eb8, 32'h4189cdb8} /* (1, 26, 17) {real, imag} */,
  {32'h40e821a8, 32'h414da604} /* (1, 26, 16) {real, imag} */,
  {32'hc05f5c18, 32'h415e1be3} /* (1, 26, 15) {real, imag} */,
  {32'h4115921a, 32'h4184f12c} /* (1, 26, 14) {real, imag} */,
  {32'h40ffcafc, 32'h3f6e07a0} /* (1, 26, 13) {real, imag} */,
  {32'h405485da, 32'h413454c7} /* (1, 26, 12) {real, imag} */,
  {32'hc12bfa88, 32'h4121e88a} /* (1, 26, 11) {real, imag} */,
  {32'hc11cb330, 32'h3fcbb114} /* (1, 26, 10) {real, imag} */,
  {32'h40f5fefc, 32'hc152c37f} /* (1, 26, 9) {real, imag} */,
  {32'h4138cc0c, 32'hc00b42b7} /* (1, 26, 8) {real, imag} */,
  {32'h4101a136, 32'hbf20ab78} /* (1, 26, 7) {real, imag} */,
  {32'h410d9dbf, 32'h40c9fc44} /* (1, 26, 6) {real, imag} */,
  {32'h40c0666a, 32'hc1554300} /* (1, 26, 5) {real, imag} */,
  {32'h41bec875, 32'hc136d256} /* (1, 26, 4) {real, imag} */,
  {32'h413c7d3a, 32'h415d74b8} /* (1, 26, 3) {real, imag} */,
  {32'h410d3217, 32'h41dc086a} /* (1, 26, 2) {real, imag} */,
  {32'h40b46b68, 32'hc0058b02} /* (1, 26, 1) {real, imag} */,
  {32'hc00a5391, 32'hc166bff4} /* (1, 26, 0) {real, imag} */,
  {32'hbfbf93d2, 32'h40b27d28} /* (1, 25, 31) {real, imag} */,
  {32'hc1aba056, 32'h4111b7ba} /* (1, 25, 30) {real, imag} */,
  {32'hc2002ff5, 32'h4104350e} /* (1, 25, 29) {real, imag} */,
  {32'h401b56f0, 32'h400cac42} /* (1, 25, 28) {real, imag} */,
  {32'hc10743a6, 32'hc183dcf7} /* (1, 25, 27) {real, imag} */,
  {32'hc1de3adf, 32'hc18570eb} /* (1, 25, 26) {real, imag} */,
  {32'hc16c516c, 32'h415c2a5a} /* (1, 25, 25) {real, imag} */,
  {32'hc1110923, 32'h419a6440} /* (1, 25, 24) {real, imag} */,
  {32'hc1b5130c, 32'h3ff8a5e0} /* (1, 25, 23) {real, imag} */,
  {32'hc1875ea4, 32'h3fda8850} /* (1, 25, 22) {real, imag} */,
  {32'h40837249, 32'h40609b20} /* (1, 25, 21) {real, imag} */,
  {32'h40ac1421, 32'hc141d7fe} /* (1, 25, 20) {real, imag} */,
  {32'h416b7008, 32'hc07373a4} /* (1, 25, 19) {real, imag} */,
  {32'h408af884, 32'h40bcaf00} /* (1, 25, 18) {real, imag} */,
  {32'h4091d58e, 32'h40286b16} /* (1, 25, 17) {real, imag} */,
  {32'h4104d268, 32'h411e8605} /* (1, 25, 16) {real, imag} */,
  {32'h3fc48da0, 32'h4011fff8} /* (1, 25, 15) {real, imag} */,
  {32'h4122238a, 32'hbec5cea0} /* (1, 25, 14) {real, imag} */,
  {32'h411b20b2, 32'hc104092a} /* (1, 25, 13) {real, imag} */,
  {32'h414f9da7, 32'h3f089de8} /* (1, 25, 12) {real, imag} */,
  {32'h41db2e6c, 32'h415cdc5c} /* (1, 25, 11) {real, imag} */,
  {32'h414085dc, 32'h41886a81} /* (1, 25, 10) {real, imag} */,
  {32'h4044e570, 32'h41063d26} /* (1, 25, 9) {real, imag} */,
  {32'hc0df691d, 32'h41a6c0fc} /* (1, 25, 8) {real, imag} */,
  {32'h4028a430, 32'h3f9dcfd4} /* (1, 25, 7) {real, imag} */,
  {32'h41613f49, 32'hc17dea2e} /* (1, 25, 6) {real, imag} */,
  {32'h41b2c79c, 32'hc1c587f4} /* (1, 25, 5) {real, imag} */,
  {32'h4147831b, 32'hc199a53c} /* (1, 25, 4) {real, imag} */,
  {32'h416bb510, 32'hc18c4557} /* (1, 25, 3) {real, imag} */,
  {32'hc0cb895b, 32'h4114132a} /* (1, 25, 2) {real, imag} */,
  {32'hc12a8530, 32'hbf3fe170} /* (1, 25, 1) {real, imag} */,
  {32'hc0a48e8a, 32'hc04ce9d1} /* (1, 25, 0) {real, imag} */,
  {32'h403ee065, 32'h3fdd9ad2} /* (1, 24, 31) {real, imag} */,
  {32'h41310caf, 32'h41af9dba} /* (1, 24, 30) {real, imag} */,
  {32'h41a3e692, 32'h421a9657} /* (1, 24, 29) {real, imag} */,
  {32'h41e4e46b, 32'h41b9fbd5} /* (1, 24, 28) {real, imag} */,
  {32'h417acf9b, 32'h40f2bc69} /* (1, 24, 27) {real, imag} */,
  {32'h41528f8c, 32'h410a1ae6} /* (1, 24, 26) {real, imag} */,
  {32'h4195df11, 32'h4044a504} /* (1, 24, 25) {real, imag} */,
  {32'h4047e3c2, 32'h4121e09d} /* (1, 24, 24) {real, imag} */,
  {32'hc08d2326, 32'h41afad52} /* (1, 24, 23) {real, imag} */,
  {32'hc0dcc556, 32'h4209f6d8} /* (1, 24, 22) {real, imag} */,
  {32'hbe03b640, 32'hc09c5e7c} /* (1, 24, 21) {real, imag} */,
  {32'hc0974629, 32'hc21d2f66} /* (1, 24, 20) {real, imag} */,
  {32'hc08fb7dd, 32'hc206938f} /* (1, 24, 19) {real, imag} */,
  {32'hc13aa859, 32'hc1cdc7c4} /* (1, 24, 18) {real, imag} */,
  {32'hc14910f3, 32'hc1ffd148} /* (1, 24, 17) {real, imag} */,
  {32'hc144da26, 32'hc1febf5e} /* (1, 24, 16) {real, imag} */,
  {32'h401ac7d2, 32'hc1a5a92c} /* (1, 24, 15) {real, imag} */,
  {32'hc159b440, 32'hc19f686d} /* (1, 24, 14) {real, imag} */,
  {32'hbff475f8, 32'hc1e3e422} /* (1, 24, 13) {real, imag} */,
  {32'hc10e802c, 32'hc19a0239} /* (1, 24, 12) {real, imag} */,
  {32'hc1248db0, 32'hc1423432} /* (1, 24, 11) {real, imag} */,
  {32'hbee182ec, 32'h413f308b} /* (1, 24, 10) {real, imag} */,
  {32'hbe3e94f0, 32'h41e4fccc} /* (1, 24, 9) {real, imag} */,
  {32'h3f1b5aa8, 32'h41b3288c} /* (1, 24, 8) {real, imag} */,
  {32'h4114371e, 32'h418d1a65} /* (1, 24, 7) {real, imag} */,
  {32'hbf48b138, 32'h41def9b5} /* (1, 24, 6) {real, imag} */,
  {32'hc107156a, 32'h41db696b} /* (1, 24, 5) {real, imag} */,
  {32'hc173b4ab, 32'h4193ae95} /* (1, 24, 4) {real, imag} */,
  {32'h4096aa50, 32'h4192539f} /* (1, 24, 3) {real, imag} */,
  {32'h41ba69d5, 32'h4123fa20} /* (1, 24, 2) {real, imag} */,
  {32'h417812da, 32'h40de3c24} /* (1, 24, 1) {real, imag} */,
  {32'h3fae24e6, 32'h3fa7b3fe} /* (1, 24, 0) {real, imag} */,
  {32'hc0c61236, 32'hc041407c} /* (1, 23, 31) {real, imag} */,
  {32'hc168937a, 32'hc12f1af0} /* (1, 23, 30) {real, imag} */,
  {32'hc0fb4a0a, 32'h40693bea} /* (1, 23, 29) {real, imag} */,
  {32'hc09e3cc2, 32'h40c7cb03} /* (1, 23, 28) {real, imag} */,
  {32'h4057d746, 32'hc12e5c45} /* (1, 23, 27) {real, imag} */,
  {32'h40dc64a8, 32'hc0f8227e} /* (1, 23, 26) {real, imag} */,
  {32'hc0fcd53d, 32'hc1033d96} /* (1, 23, 25) {real, imag} */,
  {32'hc13f7b36, 32'h4155b361} /* (1, 23, 24) {real, imag} */,
  {32'hc140750d, 32'h40864c78} /* (1, 23, 23) {real, imag} */,
  {32'hc1b5b352, 32'hc1152e62} /* (1, 23, 22) {real, imag} */,
  {32'hc156dd4a, 32'hc116a14e} /* (1, 23, 21) {real, imag} */,
  {32'h41391602, 32'hc13a8240} /* (1, 23, 20) {real, imag} */,
  {32'h418bad13, 32'h4154a4c6} /* (1, 23, 19) {real, imag} */,
  {32'h41d3f404, 32'h4146ee8e} /* (1, 23, 18) {real, imag} */,
  {32'h41fc8e18, 32'h40250986} /* (1, 23, 17) {real, imag} */,
  {32'h4218321a, 32'hc0a87550} /* (1, 23, 16) {real, imag} */,
  {32'h414e6a2d, 32'h40da7d1d} /* (1, 23, 15) {real, imag} */,
  {32'hbd9c7f40, 32'hc0808c54} /* (1, 23, 14) {real, imag} */,
  {32'hc1246a2c, 32'hc03fc384} /* (1, 23, 13) {real, imag} */,
  {32'hc1352227, 32'h41095420} /* (1, 23, 12) {real, imag} */,
  {32'hc1ce5b8e, 32'hc0043cec} /* (1, 23, 11) {real, imag} */,
  {32'hc1b4663a, 32'hc18837ed} /* (1, 23, 10) {real, imag} */,
  {32'hc1893638, 32'hc1557236} /* (1, 23, 9) {real, imag} */,
  {32'hc132a036, 32'h40cf2476} /* (1, 23, 8) {real, imag} */,
  {32'hc06cefc8, 32'h4130553e} /* (1, 23, 7) {real, imag} */,
  {32'h405f35fe, 32'hbfbd4994} /* (1, 23, 6) {real, imag} */,
  {32'hc0d670ec, 32'h412a0fa1} /* (1, 23, 5) {real, imag} */,
  {32'hc161e730, 32'h41a08868} /* (1, 23, 4) {real, imag} */,
  {32'hc0e70a98, 32'h40cf7d55} /* (1, 23, 3) {real, imag} */,
  {32'hc087bfdb, 32'hc0122456} /* (1, 23, 2) {real, imag} */,
  {32'h404b5974, 32'hbf7ed488} /* (1, 23, 1) {real, imag} */,
  {32'h3f95f338, 32'h41231b5a} /* (1, 23, 0) {real, imag} */,
  {32'h3f43f5e8, 32'hbf509dfc} /* (1, 22, 31) {real, imag} */,
  {32'h408c55a3, 32'hc0e32c2a} /* (1, 22, 30) {real, imag} */,
  {32'hc07dbba0, 32'hc05a7db2} /* (1, 22, 29) {real, imag} */,
  {32'hc069e63b, 32'h40d78bfa} /* (1, 22, 28) {real, imag} */,
  {32'hbfa3bae4, 32'h40ebb490} /* (1, 22, 27) {real, imag} */,
  {32'hc0dab460, 32'hbf59dc98} /* (1, 22, 26) {real, imag} */,
  {32'hbfc90380, 32'hc069a852} /* (1, 22, 25) {real, imag} */,
  {32'hc04b0b00, 32'hbf22a8a0} /* (1, 22, 24) {real, imag} */,
  {32'hc0d4167f, 32'h4130222c} /* (1, 22, 23) {real, imag} */,
  {32'hbf9fe410, 32'h40e1bcfc} /* (1, 22, 22) {real, imag} */,
  {32'hc0059de2, 32'h3fb8b330} /* (1, 22, 21) {real, imag} */,
  {32'hbf9a898c, 32'h411b8e3a} /* (1, 22, 20) {real, imag} */,
  {32'hbfff5d48, 32'h41254062} /* (1, 22, 19) {real, imag} */,
  {32'h40a0a176, 32'h411007c5} /* (1, 22, 18) {real, imag} */,
  {32'h4137a0d1, 32'h40e8d7de} /* (1, 22, 17) {real, imag} */,
  {32'h4033cd8f, 32'h40fedfa1} /* (1, 22, 16) {real, imag} */,
  {32'hc09c2b7d, 32'h3f9d25bc} /* (1, 22, 15) {real, imag} */,
  {32'h411fa5c6, 32'hc0bc04ec} /* (1, 22, 14) {real, imag} */,
  {32'h4153baa2, 32'hc04a2294} /* (1, 22, 13) {real, imag} */,
  {32'h408854c7, 32'h40ea6b12} /* (1, 22, 12) {real, imag} */,
  {32'h405ccd62, 32'hbef6c498} /* (1, 22, 11) {real, imag} */,
  {32'hc00bad1c, 32'h3f610fa8} /* (1, 22, 10) {real, imag} */,
  {32'hc133ed72, 32'h40b1df0a} /* (1, 22, 9) {real, imag} */,
  {32'hc17f81d2, 32'h3ff39fa0} /* (1, 22, 8) {real, imag} */,
  {32'hc1220b76, 32'hbf335e58} /* (1, 22, 7) {real, imag} */,
  {32'hc1288081, 32'hbf290d00} /* (1, 22, 6) {real, imag} */,
  {32'hc126fbb1, 32'h412e3d18} /* (1, 22, 5) {real, imag} */,
  {32'hc11cdd4a, 32'h415171aa} /* (1, 22, 4) {real, imag} */,
  {32'hc140f842, 32'h40cc97b0} /* (1, 22, 3) {real, imag} */,
  {32'hc1092922, 32'hbf8a2d64} /* (1, 22, 2) {real, imag} */,
  {32'hc1449d72, 32'hc13b8dba} /* (1, 22, 1) {real, imag} */,
  {32'hc044f5b1, 32'hc09c8c84} /* (1, 22, 0) {real, imag} */,
  {32'hbfd448e6, 32'h40eb6105} /* (1, 21, 31) {real, imag} */,
  {32'h4100f45c, 32'h41705c53} /* (1, 21, 30) {real, imag} */,
  {32'h41804e44, 32'h4187cde4} /* (1, 21, 29) {real, imag} */,
  {32'h416b3882, 32'h40af9f64} /* (1, 21, 28) {real, imag} */,
  {32'h41338662, 32'hbe8b7c20} /* (1, 21, 27) {real, imag} */,
  {32'h409cc61b, 32'hc07be782} /* (1, 21, 26) {real, imag} */,
  {32'h40e012ac, 32'h3f82d340} /* (1, 21, 25) {real, imag} */,
  {32'h416a733c, 32'h412955b8} /* (1, 21, 24) {real, imag} */,
  {32'h410420ee, 32'h415785e5} /* (1, 21, 23) {real, imag} */,
  {32'h41025f5f, 32'h3fffd4d8} /* (1, 21, 22) {real, imag} */,
  {32'h406f938a, 32'hbf941b9c} /* (1, 21, 21) {real, imag} */,
  {32'hc0e1b720, 32'h3f71395c} /* (1, 21, 20) {real, imag} */,
  {32'hc11aca78, 32'hbf37eefe} /* (1, 21, 19) {real, imag} */,
  {32'hc1169da1, 32'h40a2cb6f} /* (1, 21, 18) {real, imag} */,
  {32'hc058da61, 32'hbded0d00} /* (1, 21, 17) {real, imag} */,
  {32'hc1023b3f, 32'hc10fbc32} /* (1, 21, 16) {real, imag} */,
  {32'hc13fe85c, 32'hc0b88cf8} /* (1, 21, 15) {real, imag} */,
  {32'hc0e390f4, 32'hbec9cdf0} /* (1, 21, 14) {real, imag} */,
  {32'hc15fd3de, 32'h40cf0afb} /* (1, 21, 13) {real, imag} */,
  {32'hc17bd7bc, 32'hc1398843} /* (1, 21, 12) {real, imag} */,
  {32'hc0a256b8, 32'hc0f2f482} /* (1, 21, 11) {real, imag} */,
  {32'h3fdd82e4, 32'h3fcfbace} /* (1, 21, 10) {real, imag} */,
  {32'h412cfb29, 32'h4103a2da} /* (1, 21, 9) {real, imag} */,
  {32'h418f326f, 32'h40d50866} /* (1, 21, 8) {real, imag} */,
  {32'h41018209, 32'h40c87421} /* (1, 21, 7) {real, imag} */,
  {32'h412c0247, 32'h40b1a11f} /* (1, 21, 6) {real, imag} */,
  {32'h410c5352, 32'h410291f7} /* (1, 21, 5) {real, imag} */,
  {32'h40fffd4a, 32'h40bed4d0} /* (1, 21, 4) {real, imag} */,
  {32'h409022f0, 32'h40fd0ca9} /* (1, 21, 3) {real, imag} */,
  {32'h40e789a1, 32'h4112b60e} /* (1, 21, 2) {real, imag} */,
  {32'h4150ac20, 32'hc0a1b6d8} /* (1, 21, 1) {real, imag} */,
  {32'h40d2ede2, 32'hc0e8d00c} /* (1, 21, 0) {real, imag} */,
  {32'h3fc9a40b, 32'hc0358e9a} /* (1, 20, 31) {real, imag} */,
  {32'h3faa41c0, 32'h40183cb8} /* (1, 20, 30) {real, imag} */,
  {32'hc0a22656, 32'h410e123e} /* (1, 20, 29) {real, imag} */,
  {32'hc0c947c0, 32'h3fd115e8} /* (1, 20, 28) {real, imag} */,
  {32'h3fe09552, 32'hbf7416e8} /* (1, 20, 27) {real, imag} */,
  {32'h40970c87, 32'hc0820d4c} /* (1, 20, 26) {real, imag} */,
  {32'hc0d676d3, 32'hbf94e044} /* (1, 20, 25) {real, imag} */,
  {32'hc08f5e00, 32'hc0d6a04d} /* (1, 20, 24) {real, imag} */,
  {32'hc117340c, 32'hc00274fa} /* (1, 20, 23) {real, imag} */,
  {32'hc0ee753e, 32'h40f9e0f0} /* (1, 20, 22) {real, imag} */,
  {32'hbf2bcdf8, 32'h40e9750a} /* (1, 20, 21) {real, imag} */,
  {32'hbf74fe24, 32'h4113d0f9} /* (1, 20, 20) {real, imag} */,
  {32'hc09568f4, 32'h40974d7a} /* (1, 20, 19) {real, imag} */,
  {32'hc16dbcc2, 32'h405f802c} /* (1, 20, 18) {real, imag} */,
  {32'hc18cbc1c, 32'h410e150a} /* (1, 20, 17) {real, imag} */,
  {32'hc16f2fec, 32'h406bd79a} /* (1, 20, 16) {real, imag} */,
  {32'hc085037c, 32'h3e250f10} /* (1, 20, 15) {real, imag} */,
  {32'hc0bc2c2b, 32'hbfa00676} /* (1, 20, 14) {real, imag} */,
  {32'hc0ec36ad, 32'h3c73c400} /* (1, 20, 13) {real, imag} */,
  {32'hc0e7018c, 32'h40581348} /* (1, 20, 12) {real, imag} */,
  {32'hc0d87060, 32'h40ecfc0a} /* (1, 20, 11) {real, imag} */,
  {32'hc088c4e5, 32'h414191ef} /* (1, 20, 10) {real, imag} */,
  {32'hc01d2ec8, 32'h40e33b2a} /* (1, 20, 9) {real, imag} */,
  {32'hbf8afc2c, 32'hc0875a9f} /* (1, 20, 8) {real, imag} */,
  {32'hbec664e0, 32'h40e70908} /* (1, 20, 7) {real, imag} */,
  {32'hbfb430c0, 32'h40b94e58} /* (1, 20, 6) {real, imag} */,
  {32'hc0aa7a3a, 32'h40a6304c} /* (1, 20, 5) {real, imag} */,
  {32'h3f437cac, 32'h412bf204} /* (1, 20, 4) {real, imag} */,
  {32'h407dbe55, 32'h402793ee} /* (1, 20, 3) {real, imag} */,
  {32'hc0ba131a, 32'hc0c42c36} /* (1, 20, 2) {real, imag} */,
  {32'hbfbdf731, 32'h3fe0fb3d} /* (1, 20, 1) {real, imag} */,
  {32'h3fcf44b6, 32'hc01831b0} /* (1, 20, 0) {real, imag} */,
  {32'hc00dbb69, 32'hc0b5f6bb} /* (1, 19, 31) {real, imag} */,
  {32'hc0aeb5bb, 32'hbfd067fc} /* (1, 19, 30) {real, imag} */,
  {32'h408870e6, 32'h40b4c57f} /* (1, 19, 29) {real, imag} */,
  {32'h40893b34, 32'h41149622} /* (1, 19, 28) {real, imag} */,
  {32'hbf7c5d8a, 32'h402d2da4} /* (1, 19, 27) {real, imag} */,
  {32'h4027f5fc, 32'h40b74f71} /* (1, 19, 26) {real, imag} */,
  {32'h4068c326, 32'h40da0238} /* (1, 19, 25) {real, imag} */,
  {32'h40b09e7c, 32'h3f35988c} /* (1, 19, 24) {real, imag} */,
  {32'h40ad07ba, 32'h408bab04} /* (1, 19, 23) {real, imag} */,
  {32'h407f17d8, 32'h407f7706} /* (1, 19, 22) {real, imag} */,
  {32'h4075c740, 32'h40ee87ea} /* (1, 19, 21) {real, imag} */,
  {32'h3f018ec8, 32'h4075098e} /* (1, 19, 20) {real, imag} */,
  {32'hbeaf9320, 32'hbfdbdf14} /* (1, 19, 19) {real, imag} */,
  {32'hc02d617c, 32'hbf19cbd0} /* (1, 19, 18) {real, imag} */,
  {32'hc050a33f, 32'h40865942} /* (1, 19, 17) {real, imag} */,
  {32'hc051164d, 32'h406e0030} /* (1, 19, 16) {real, imag} */,
  {32'hc039cd10, 32'hc0acc34c} /* (1, 19, 15) {real, imag} */,
  {32'hc0a6e0a8, 32'hc0e79f42} /* (1, 19, 14) {real, imag} */,
  {32'hc0a641dc, 32'hc0895d01} /* (1, 19, 13) {real, imag} */,
  {32'hc0893444, 32'hc0f03804} /* (1, 19, 12) {real, imag} */,
  {32'h403caba1, 32'h3f3f8ed0} /* (1, 19, 11) {real, imag} */,
  {32'hbf02f290, 32'h40ecde01} /* (1, 19, 10) {real, imag} */,
  {32'hc1004f64, 32'hc07d6676} /* (1, 19, 9) {real, imag} */,
  {32'hc17b1ef1, 32'hc04be2fa} /* (1, 19, 8) {real, imag} */,
  {32'hc181d3f3, 32'h4080ac8d} /* (1, 19, 7) {real, imag} */,
  {32'hbfc13eb8, 32'hbfbdcafc} /* (1, 19, 6) {real, imag} */,
  {32'h409df282, 32'hc1385c3b} /* (1, 19, 5) {real, imag} */,
  {32'h4012ad51, 32'hc0e9f31f} /* (1, 19, 4) {real, imag} */,
  {32'hc1028c49, 32'hc06d8cd5} /* (1, 19, 3) {real, imag} */,
  {32'hc0ab60d5, 32'h3fc7e424} /* (1, 19, 2) {real, imag} */,
  {32'hbebe6408, 32'h3f8f9f3a} /* (1, 19, 1) {real, imag} */,
  {32'hbfb492d2, 32'h3ee7cb48} /* (1, 19, 0) {real, imag} */,
  {32'h40c508e8, 32'hbf108be8} /* (1, 18, 31) {real, imag} */,
  {32'h414cdd38, 32'h407f286c} /* (1, 18, 30) {real, imag} */,
  {32'h415b0e56, 32'h40129644} /* (1, 18, 29) {real, imag} */,
  {32'h411b9a8c, 32'h3f999a1c} /* (1, 18, 28) {real, imag} */,
  {32'h40c5f1d4, 32'h3eaaa150} /* (1, 18, 27) {real, imag} */,
  {32'h3f808fec, 32'h3f9479f2} /* (1, 18, 26) {real, imag} */,
  {32'h403daf28, 32'h40c13c30} /* (1, 18, 25) {real, imag} */,
  {32'h40b2d35b, 32'h40aac92c} /* (1, 18, 24) {real, imag} */,
  {32'h3fa909c0, 32'hbeafd480} /* (1, 18, 23) {real, imag} */,
  {32'h408f6e06, 32'hc00a8810} /* (1, 18, 22) {real, imag} */,
  {32'h411cb8ca, 32'h40ae61d2} /* (1, 18, 21) {real, imag} */,
  {32'h40863688, 32'h40aefcf3} /* (1, 18, 20) {real, imag} */,
  {32'hc09ea9a6, 32'h3f66b60a} /* (1, 18, 19) {real, imag} */,
  {32'hc0423070, 32'h3ef1b2e0} /* (1, 18, 18) {real, imag} */,
  {32'hc0899295, 32'h3e8b83a0} /* (1, 18, 17) {real, imag} */,
  {32'hc0d776b5, 32'hbfed058c} /* (1, 18, 16) {real, imag} */,
  {32'hc0b006b6, 32'hc0f1447e} /* (1, 18, 15) {real, imag} */,
  {32'hc0adb785, 32'h3fb6b584} /* (1, 18, 14) {real, imag} */,
  {32'hc03b7f18, 32'hbff49d58} /* (1, 18, 13) {real, imag} */,
  {32'hbf151b4c, 32'hc09034a7} /* (1, 18, 12) {real, imag} */,
  {32'hc12ea01c, 32'h3edefb10} /* (1, 18, 11) {real, imag} */,
  {32'h3e96a460, 32'h410fb21e} /* (1, 18, 10) {real, imag} */,
  {32'h40461c34, 32'h40aa5013} /* (1, 18, 9) {real, imag} */,
  {32'h40284508, 32'h3fb3c5a8} /* (1, 18, 8) {real, imag} */,
  {32'h3e7ccf80, 32'h402478f8} /* (1, 18, 7) {real, imag} */,
  {32'hbfd98ba8, 32'h4065ca04} /* (1, 18, 6) {real, imag} */,
  {32'h40805120, 32'hc0a9cec3} /* (1, 18, 5) {real, imag} */,
  {32'h40df3fa4, 32'hc0c86379} /* (1, 18, 4) {real, imag} */,
  {32'h40a13092, 32'h3e82c560} /* (1, 18, 3) {real, imag} */,
  {32'h40025158, 32'h404170dc} /* (1, 18, 2) {real, imag} */,
  {32'h40404364, 32'h3fd6ec3c} /* (1, 18, 1) {real, imag} */,
  {32'h3ff98236, 32'h3f50f6b0} /* (1, 18, 0) {real, imag} */,
  {32'hc05da3e3, 32'hc08d8ed2} /* (1, 17, 31) {real, imag} */,
  {32'hc0d35c78, 32'hc00fb4f0} /* (1, 17, 30) {real, imag} */,
  {32'hbf58f234, 32'h4048ebda} /* (1, 17, 29) {real, imag} */,
  {32'hbfa18c64, 32'h40a92bbf} /* (1, 17, 28) {real, imag} */,
  {32'h3fbe4940, 32'h3e1913c0} /* (1, 17, 27) {real, imag} */,
  {32'h3c81be00, 32'hbf94f518} /* (1, 17, 26) {real, imag} */,
  {32'hc0295fc2, 32'h3d06f740} /* (1, 17, 25) {real, imag} */,
  {32'hbfb748ec, 32'h40292c6d} /* (1, 17, 24) {real, imag} */,
  {32'hc050fd88, 32'h40876ae1} /* (1, 17, 23) {real, imag} */,
  {32'hbf09bdf4, 32'h406c7764} /* (1, 17, 22) {real, imag} */,
  {32'h3fd0295c, 32'h40746298} /* (1, 17, 21) {real, imag} */,
  {32'h407b2f0a, 32'h3ff2d940} /* (1, 17, 20) {real, imag} */,
  {32'hc0322bc2, 32'hc09544e7} /* (1, 17, 19) {real, imag} */,
  {32'hc069d040, 32'hbfaef194} /* (1, 17, 18) {real, imag} */,
  {32'h40c93f1a, 32'h3fe3cfc8} /* (1, 17, 17) {real, imag} */,
  {32'h4014557a, 32'hc0720cd8} /* (1, 17, 16) {real, imag} */,
  {32'hc04ca58b, 32'hc0384428} /* (1, 17, 15) {real, imag} */,
  {32'hc07697a7, 32'h40952ed9} /* (1, 17, 14) {real, imag} */,
  {32'hbeb8ada0, 32'h40922460} /* (1, 17, 13) {real, imag} */,
  {32'hbf84e0c8, 32'h3f908cbe} /* (1, 17, 12) {real, imag} */,
  {32'hc018eacf, 32'hc1028bdf} /* (1, 17, 11) {real, imag} */,
  {32'h3fdc096c, 32'hc116554a} /* (1, 17, 10) {real, imag} */,
  {32'hbed93360, 32'hbfcfcfa6} /* (1, 17, 9) {real, imag} */,
  {32'hc1176624, 32'h40458946} /* (1, 17, 8) {real, imag} */,
  {32'hc0f1bd0e, 32'h3e678540} /* (1, 17, 7) {real, imag} */,
  {32'hc008da54, 32'hbe01cad0} /* (1, 17, 6) {real, imag} */,
  {32'hc0a1c3c6, 32'h3f38b830} /* (1, 17, 5) {real, imag} */,
  {32'hc091b973, 32'h3f3cf624} /* (1, 17, 4) {real, imag} */,
  {32'hc0ae4a76, 32'h3db0dd80} /* (1, 17, 3) {real, imag} */,
  {32'hc0afda70, 32'h3e560240} /* (1, 17, 2) {real, imag} */,
  {32'hc07667d5, 32'h40ae9c35} /* (1, 17, 1) {real, imag} */,
  {32'hc021ece4, 32'h403c1e28} /* (1, 17, 0) {real, imag} */,
  {32'hbf9ec0f8, 32'h40b404b0} /* (1, 16, 31) {real, imag} */,
  {32'hbe7d4c80, 32'h411c2cd8} /* (1, 16, 30) {real, imag} */,
  {32'h3ea163b0, 32'h40c0c1f0} /* (1, 16, 29) {real, imag} */,
  {32'hbf10d568, 32'hbfb71860} /* (1, 16, 28) {real, imag} */,
  {32'hc07405bc, 32'hc086eb90} /* (1, 16, 27) {real, imag} */,
  {32'hc0876bea, 32'hbfcca700} /* (1, 16, 26) {real, imag} */,
  {32'hbf5756b8, 32'h3f2db080} /* (1, 16, 25) {real, imag} */,
  {32'h3f2673d4, 32'hc0ad1f30} /* (1, 16, 24) {real, imag} */,
  {32'hbffd10c0, 32'hc085cf60} /* (1, 16, 23) {real, imag} */,
  {32'h4076f940, 32'hc0b9d578} /* (1, 16, 22) {real, imag} */,
  {32'h40bb324b, 32'h402ff3d0} /* (1, 16, 21) {real, imag} */,
  {32'h3da4c240, 32'h3ce16c00} /* (1, 16, 20) {real, imag} */,
  {32'hc044fdfa, 32'hc0172cae} /* (1, 16, 19) {real, imag} */,
  {32'hbf2ae078, 32'h3f71c268} /* (1, 16, 18) {real, imag} */,
  {32'hbf3ab6e8, 32'hc04b06dc} /* (1, 16, 17) {real, imag} */,
  {32'hbd83b280, 32'h40843e8c} /* (1, 16, 16) {real, imag} */,
  {32'hc0b313ba, 32'h404f3be0} /* (1, 16, 15) {real, imag} */,
  {32'hc0b35530, 32'hc02d97e0} /* (1, 16, 14) {real, imag} */,
  {32'hc0742b44, 32'hc0a273b0} /* (1, 16, 13) {real, imag} */,
  {32'hbeb6a510, 32'h3f20a240} /* (1, 16, 12) {real, imag} */,
  {32'hc0a5a546, 32'hbf123780} /* (1, 16, 11) {real, imag} */,
  {32'hc08d63c6, 32'h3ff5997c} /* (1, 16, 10) {real, imag} */,
  {32'hbe8c3280, 32'h3fadb610} /* (1, 16, 9) {real, imag} */,
  {32'hbf199120, 32'h3f363728} /* (1, 16, 8) {real, imag} */,
  {32'hbf0f55a0, 32'hbffb4f80} /* (1, 16, 7) {real, imag} */,
  {32'h4031427c, 32'hc080fc25} /* (1, 16, 6) {real, imag} */,
  {32'h408fb1da, 32'hbea6bb80} /* (1, 16, 5) {real, imag} */,
  {32'h403b5e73, 32'hbf019700} /* (1, 16, 4) {real, imag} */,
  {32'h409767ef, 32'hc08658a8} /* (1, 16, 3) {real, imag} */,
  {32'h402e700c, 32'hc0ab4ae0} /* (1, 16, 2) {real, imag} */,
  {32'h40b34e31, 32'h40425690} /* (1, 16, 1) {real, imag} */,
  {32'h4016ed69, 32'h3ff46260} /* (1, 16, 0) {real, imag} */,
  {32'h3f4b651c, 32'hbf91e4b6} /* (1, 15, 31) {real, imag} */,
  {32'h40fbafc8, 32'hc03cc590} /* (1, 15, 30) {real, imag} */,
  {32'h4031e7df, 32'h3fc1944c} /* (1, 15, 29) {real, imag} */,
  {32'hc05ad182, 32'h3f966104} /* (1, 15, 28) {real, imag} */,
  {32'h4061a8e6, 32'h3f1b8810} /* (1, 15, 27) {real, imag} */,
  {32'h40d02b26, 32'h3f559830} /* (1, 15, 26) {real, imag} */,
  {32'h4025238e, 32'hc0cb870e} /* (1, 15, 25) {real, imag} */,
  {32'h40ded49f, 32'hc09c19b6} /* (1, 15, 24) {real, imag} */,
  {32'h40b58f9e, 32'hbee36c10} /* (1, 15, 23) {real, imag} */,
  {32'h3b9c2200, 32'hc0dc6332} /* (1, 15, 22) {real, imag} */,
  {32'hbf95727c, 32'hc10a0e1e} /* (1, 15, 21) {real, imag} */,
  {32'hc0454326, 32'hc0939170} /* (1, 15, 20) {real, imag} */,
  {32'hc0d716e9, 32'h3f187f78} /* (1, 15, 19) {real, imag} */,
  {32'hc04ee9f0, 32'h3fc72814} /* (1, 15, 18) {real, imag} */,
  {32'hc008985c, 32'h40540c7c} /* (1, 15, 17) {real, imag} */,
  {32'hbfd3e2cc, 32'h3fc0bff0} /* (1, 15, 16) {real, imag} */,
  {32'hc00e8495, 32'h3f0637a0} /* (1, 15, 15) {real, imag} */,
  {32'h3f8f440e, 32'h4058150e} /* (1, 15, 14) {real, imag} */,
  {32'hc03c4c64, 32'h3fa38f00} /* (1, 15, 13) {real, imag} */,
  {32'hc004214c, 32'hc07bf25f} /* (1, 15, 12) {real, imag} */,
  {32'h3f32175c, 32'h3fe765f8} /* (1, 15, 11) {real, imag} */,
  {32'hbdd9f340, 32'h3fdab04c} /* (1, 15, 10) {real, imag} */,
  {32'hbef27360, 32'h3eed5298} /* (1, 15, 9) {real, imag} */,
  {32'hbffd65c0, 32'hc0715db6} /* (1, 15, 8) {real, imag} */,
  {32'hbeb40d58, 32'hc04e8454} /* (1, 15, 7) {real, imag} */,
  {32'h41051e53, 32'h4047086d} /* (1, 15, 6) {real, imag} */,
  {32'h409a48de, 32'h409074fa} /* (1, 15, 5) {real, imag} */,
  {32'h4040d572, 32'h40736f57} /* (1, 15, 4) {real, imag} */,
  {32'hc0c590ae, 32'h3fe59e28} /* (1, 15, 3) {real, imag} */,
  {32'hc0c94520, 32'hc08bba32} /* (1, 15, 2) {real, imag} */,
  {32'h40476505, 32'hc0ea0db5} /* (1, 15, 1) {real, imag} */,
  {32'h3fd6c1f0, 32'hc01a7168} /* (1, 15, 0) {real, imag} */,
  {32'hc01ff260, 32'hc0664c46} /* (1, 14, 31) {real, imag} */,
  {32'hc0c0f420, 32'hc0e697a6} /* (1, 14, 30) {real, imag} */,
  {32'hc1216a70, 32'hc103c0f1} /* (1, 14, 29) {real, imag} */,
  {32'hc113b7dc, 32'hc02b008e} /* (1, 14, 28) {real, imag} */,
  {32'hc0a95068, 32'hc0ca56b5} /* (1, 14, 27) {real, imag} */,
  {32'h4089f825, 32'hc0759c59} /* (1, 14, 26) {real, imag} */,
  {32'hc0512a5c, 32'hc0a8e7f0} /* (1, 14, 25) {real, imag} */,
  {32'hc1103f10, 32'hc0b3925c} /* (1, 14, 24) {real, imag} */,
  {32'hc112b7ee, 32'h3f81bf60} /* (1, 14, 23) {real, imag} */,
  {32'hc0e151a4, 32'h40d29d88} /* (1, 14, 22) {real, imag} */,
  {32'h40ac53b8, 32'h403e843c} /* (1, 14, 21) {real, imag} */,
  {32'h411a2880, 32'hc04e6546} /* (1, 14, 20) {real, imag} */,
  {32'h40db1312, 32'hbf71128a} /* (1, 14, 19) {real, imag} */,
  {32'h402112c0, 32'hbead14e0} /* (1, 14, 18) {real, imag} */,
  {32'h3fd2308c, 32'hc001aef4} /* (1, 14, 17) {real, imag} */,
  {32'h4099ab63, 32'hbffb6bf4} /* (1, 14, 16) {real, imag} */,
  {32'h40a1541a, 32'hbec2ec20} /* (1, 14, 15) {real, imag} */,
  {32'h40a3ffd9, 32'h3e5b59e0} /* (1, 14, 14) {real, imag} */,
  {32'h4008f688, 32'hc0033cd4} /* (1, 14, 13) {real, imag} */,
  {32'h407734bd, 32'h3ef03470} /* (1, 14, 12) {real, imag} */,
  {32'h408dd264, 32'hc008b902} /* (1, 14, 11) {real, imag} */,
  {32'hbf6681d0, 32'hc072ec96} /* (1, 14, 10) {real, imag} */,
  {32'hbfce3018, 32'h3e5f21a0} /* (1, 14, 9) {real, imag} */,
  {32'hbe4b9680, 32'h403e9fec} /* (1, 14, 8) {real, imag} */,
  {32'hbf9ffbd0, 32'h40aca254} /* (1, 14, 7) {real, imag} */,
  {32'hc08239ca, 32'hbefb3420} /* (1, 14, 6) {real, imag} */,
  {32'hc0a1e450, 32'hc09fc49d} /* (1, 14, 5) {real, imag} */,
  {32'hc12e212e, 32'hc113898c} /* (1, 14, 4) {real, imag} */,
  {32'hc13dbc4b, 32'hc1086493} /* (1, 14, 3) {real, imag} */,
  {32'hc0d12ea4, 32'hc0e0a60e} /* (1, 14, 2) {real, imag} */,
  {32'hc12d3439, 32'hc01b871e} /* (1, 14, 1) {real, imag} */,
  {32'hc0e69828, 32'hbe8e0f60} /* (1, 14, 0) {real, imag} */,
  {32'h40b9a2a0, 32'hbf9e3d3c} /* (1, 13, 31) {real, imag} */,
  {32'h4102e7ae, 32'hbf8e3b6c} /* (1, 13, 30) {real, imag} */,
  {32'h3ec5c318, 32'hc0eb97c1} /* (1, 13, 29) {real, imag} */,
  {32'hbffdffa2, 32'hc0b39490} /* (1, 13, 28) {real, imag} */,
  {32'h4002fa44, 32'hc095d2e4} /* (1, 13, 27) {real, imag} */,
  {32'hc00a6d8a, 32'hc0b15217} /* (1, 13, 26) {real, imag} */,
  {32'hc049f3da, 32'hbec64380} /* (1, 13, 25) {real, imag} */,
  {32'hc0f2479a, 32'h3f46a8a4} /* (1, 13, 24) {real, imag} */,
  {32'hbe258640, 32'hc0bf3034} /* (1, 13, 23) {real, imag} */,
  {32'h4103e320, 32'hc1263b70} /* (1, 13, 22) {real, imag} */,
  {32'h401b1adc, 32'hbff23648} /* (1, 13, 21) {real, imag} */,
  {32'h3f98b424, 32'h3fe3e3b4} /* (1, 13, 20) {real, imag} */,
  {32'h3f06b330, 32'h3fb4c874} /* (1, 13, 19) {real, imag} */,
  {32'h40780514, 32'hc058fac0} /* (1, 13, 18) {real, imag} */,
  {32'h3f639804, 32'hc179adcb} /* (1, 13, 17) {real, imag} */,
  {32'h40a50ff2, 32'hc089bc5c} /* (1, 13, 16) {real, imag} */,
  {32'h40cb50b8, 32'h40a5b988} /* (1, 13, 15) {real, imag} */,
  {32'h40119581, 32'h417fc5b3} /* (1, 13, 14) {real, imag} */,
  {32'hbfd58752, 32'h4115b304} /* (1, 13, 13) {real, imag} */,
  {32'h4044ec3e, 32'h41016ed2} /* (1, 13, 12) {real, imag} */,
  {32'h40117d5b, 32'h4143f4f0} /* (1, 13, 11) {real, imag} */,
  {32'hc026e674, 32'h414a0da8} /* (1, 13, 10) {real, imag} */,
  {32'h40324b81, 32'h41395246} /* (1, 13, 9) {real, imag} */,
  {32'h408e606e, 32'h41800439} /* (1, 13, 8) {real, imag} */,
  {32'h3ffe06cc, 32'h411e4864} /* (1, 13, 7) {real, imag} */,
  {32'hc076935c, 32'h40a66fe9} /* (1, 13, 6) {real, imag} */,
  {32'hc09af39e, 32'hbed5f520} /* (1, 13, 5) {real, imag} */,
  {32'hc09d44de, 32'h3fe65ad4} /* (1, 13, 4) {real, imag} */,
  {32'h3f622a90, 32'h3febf586} /* (1, 13, 3) {real, imag} */,
  {32'h40efc147, 32'hc1438216} /* (1, 13, 2) {real, imag} */,
  {32'h409f625c, 32'hc1095548} /* (1, 13, 1) {real, imag} */,
  {32'h3f8eaa0a, 32'hbf22c2dc} /* (1, 13, 0) {real, imag} */,
  {32'h3f32d496, 32'hc0722b52} /* (1, 12, 31) {real, imag} */,
  {32'h40f444fc, 32'h3f49be80} /* (1, 12, 30) {real, imag} */,
  {32'h40dfeb9e, 32'hbf2c6748} /* (1, 12, 29) {real, imag} */,
  {32'hc089f33a, 32'h3f22c230} /* (1, 12, 28) {real, imag} */,
  {32'h404f4759, 32'hbfee58cc} /* (1, 12, 27) {real, imag} */,
  {32'h413f9b22, 32'hbfe0b170} /* (1, 12, 26) {real, imag} */,
  {32'h3f372450, 32'h40a9a3ad} /* (1, 12, 25) {real, imag} */,
  {32'hc1752f74, 32'h40fb1bc3} /* (1, 12, 24) {real, imag} */,
  {32'hc0968597, 32'h4101e33c} /* (1, 12, 23) {real, imag} */,
  {32'h412d8815, 32'h41276808} /* (1, 12, 22) {real, imag} */,
  {32'h410f0746, 32'h40a841ee} /* (1, 12, 21) {real, imag} */,
  {32'h40982d14, 32'h408e5ce2} /* (1, 12, 20) {real, imag} */,
  {32'h40d4e354, 32'h40dfedf6} /* (1, 12, 19) {real, imag} */,
  {32'h410e919e, 32'h409b6be6} /* (1, 12, 18) {real, imag} */,
  {32'h3fa44158, 32'h40f4fcc8} /* (1, 12, 17) {real, imag} */,
  {32'hbf692f00, 32'h40832d53} /* (1, 12, 16) {real, imag} */,
  {32'h3f0bd980, 32'h40b56eba} /* (1, 12, 15) {real, imag} */,
  {32'hbf904c8c, 32'h3cd3c180} /* (1, 12, 14) {real, imag} */,
  {32'hc097f02b, 32'hc01b3bd4} /* (1, 12, 13) {real, imag} */,
  {32'hc0013208, 32'hbf233cc0} /* (1, 12, 12) {real, imag} */,
  {32'h3d42de80, 32'h405b8b59} /* (1, 12, 11) {real, imag} */,
  {32'hc04cb722, 32'hc08649ca} /* (1, 12, 10) {real, imag} */,
  {32'hbf4daa20, 32'hc0a2010a} /* (1, 12, 9) {real, imag} */,
  {32'h40b69cfd, 32'hbf5d2746} /* (1, 12, 8) {real, imag} */,
  {32'h4138322d, 32'hc0b8bc98} /* (1, 12, 7) {real, imag} */,
  {32'hc0238e60, 32'hc02b07c0} /* (1, 12, 6) {real, imag} */,
  {32'hc101fe5f, 32'h3ea537c0} /* (1, 12, 5) {real, imag} */,
  {32'h3f25d21c, 32'hc120e318} /* (1, 12, 4) {real, imag} */,
  {32'h3e1eb630, 32'hc11d9a22} /* (1, 12, 3) {real, imag} */,
  {32'h3f7c35b0, 32'h3f238690} /* (1, 12, 2) {real, imag} */,
  {32'h40a7ecc2, 32'hc097c3e1} /* (1, 12, 1) {real, imag} */,
  {32'hbf98f426, 32'hc0aa6b18} /* (1, 12, 0) {real, imag} */,
  {32'hc039231f, 32'h410c3b6e} /* (1, 11, 31) {real, imag} */,
  {32'hbfcc77aa, 32'h40c4e8fa} /* (1, 11, 30) {real, imag} */,
  {32'hbea3dce0, 32'h4158b014} /* (1, 11, 29) {real, imag} */,
  {32'hc01ec996, 32'h40fecb96} /* (1, 11, 28) {real, imag} */,
  {32'hc161514c, 32'h3f6886b0} /* (1, 11, 27) {real, imag} */,
  {32'hc12bc0aa, 32'h40426fe6} /* (1, 11, 26) {real, imag} */,
  {32'hc1001510, 32'h3fdbb500} /* (1, 11, 25) {real, imag} */,
  {32'hc0cc4667, 32'h3f8e4680} /* (1, 11, 24) {real, imag} */,
  {32'hc112ad86, 32'h411dcd33} /* (1, 11, 23) {real, imag} */,
  {32'hc16cc1c3, 32'h41167f61} /* (1, 11, 22) {real, imag} */,
  {32'hc1623ea2, 32'h4041f86e} /* (1, 11, 21) {real, imag} */,
  {32'hc0ebdb48, 32'hbe11c450} /* (1, 11, 20) {real, imag} */,
  {32'hbf3581c8, 32'hc0751108} /* (1, 11, 19) {real, imag} */,
  {32'h4067f6d3, 32'hc1236170} /* (1, 11, 18) {real, imag} */,
  {32'h3fd1f15e, 32'hc14c0ce2} /* (1, 11, 17) {real, imag} */,
  {32'h409ae1ea, 32'hc141de3e} /* (1, 11, 16) {real, imag} */,
  {32'h40b11f30, 32'hc105d136} /* (1, 11, 15) {real, imag} */,
  {32'h410a58b6, 32'h3ffcd34c} /* (1, 11, 14) {real, imag} */,
  {32'h40cb93d5, 32'hc027d376} /* (1, 11, 13) {real, imag} */,
  {32'h4148469a, 32'hc10d1499} /* (1, 11, 12) {real, imag} */,
  {32'h41712180, 32'hc119b483} /* (1, 11, 11) {real, imag} */,
  {32'hbf62e3b8, 32'h4059f82f} /* (1, 11, 10) {real, imag} */,
  {32'hc1105981, 32'h3f0a9de8} /* (1, 11, 9) {real, imag} */,
  {32'hc111c9f6, 32'hc0a3c4c0} /* (1, 11, 8) {real, imag} */,
  {32'hc183afe6, 32'hc0a13e5f} /* (1, 11, 7) {real, imag} */,
  {32'hc0f9414b, 32'hc0801bc1} /* (1, 11, 6) {real, imag} */,
  {32'hbfa97dfe, 32'hbfb9b108} /* (1, 11, 5) {real, imag} */,
  {32'hc15278a7, 32'h4034ec89} /* (1, 11, 4) {real, imag} */,
  {32'hc16b02c8, 32'h40c2a4e7} /* (1, 11, 3) {real, imag} */,
  {32'hbf6398f8, 32'h3fd878d4} /* (1, 11, 2) {real, imag} */,
  {32'h3e809380, 32'h403d21a8} /* (1, 11, 1) {real, imag} */,
  {32'hc08fde24, 32'h40c616c4} /* (1, 11, 0) {real, imag} */,
  {32'h4056c3ea, 32'hbf9ec7ca} /* (1, 10, 31) {real, imag} */,
  {32'hc05c7946, 32'h41210e09} /* (1, 10, 30) {real, imag} */,
  {32'hc18f5d20, 32'h4091e5d1} /* (1, 10, 29) {real, imag} */,
  {32'hc073f645, 32'hc0fd0be2} /* (1, 10, 28) {real, imag} */,
  {32'h403f12a6, 32'hc1779b7a} /* (1, 10, 27) {real, imag} */,
  {32'hc09b3310, 32'hc12997d8} /* (1, 10, 26) {real, imag} */,
  {32'h41087476, 32'hbfc03f94} /* (1, 10, 25) {real, imag} */,
  {32'h41160532, 32'h40978b7a} /* (1, 10, 24) {real, imag} */,
  {32'h411550a4, 32'h3f24abe8} /* (1, 10, 23) {real, imag} */,
  {32'h41a146e9, 32'h41023690} /* (1, 10, 22) {real, imag} */,
  {32'h40d749bb, 32'hc118175c} /* (1, 10, 21) {real, imag} */,
  {32'hc009c76e, 32'hc0b87fbd} /* (1, 10, 20) {real, imag} */,
  {32'hc1033bcd, 32'h41624390} /* (1, 10, 19) {real, imag} */,
  {32'hc19d35bc, 32'h414d0b7b} /* (1, 10, 18) {real, imag} */,
  {32'hc1395b3f, 32'h3f9af798} /* (1, 10, 17) {real, imag} */,
  {32'hc0c52df8, 32'h40ec4377} /* (1, 10, 16) {real, imag} */,
  {32'hc0c7bdc5, 32'hbea2c230} /* (1, 10, 15) {real, imag} */,
  {32'hc08685d5, 32'hc00b99d0} /* (1, 10, 14) {real, imag} */,
  {32'hc0763668, 32'h4019e320} /* (1, 10, 13) {real, imag} */,
  {32'hc1101f3e, 32'h410d26cb} /* (1, 10, 12) {real, imag} */,
  {32'hc1166cce, 32'h40d1bf54} /* (1, 10, 11) {real, imag} */,
  {32'h40a62f76, 32'h40dad899} /* (1, 10, 10) {real, imag} */,
  {32'h413caaf6, 32'h3db7ae80} /* (1, 10, 9) {real, imag} */,
  {32'h412cd2d0, 32'hc169974c} /* (1, 10, 8) {real, imag} */,
  {32'h40ee5378, 32'hc139d0a8} /* (1, 10, 7) {real, imag} */,
  {32'h414972c5, 32'hc144af14} /* (1, 10, 6) {real, imag} */,
  {32'h411de349, 32'hbecc7b30} /* (1, 10, 5) {real, imag} */,
  {32'h40a43d93, 32'hc02cfbca} /* (1, 10, 4) {real, imag} */,
  {32'hbfceef44, 32'hbe29fa80} /* (1, 10, 3) {real, imag} */,
  {32'h3f80b732, 32'hbf11a538} /* (1, 10, 2) {real, imag} */,
  {32'h40f15337, 32'hc0f709b9} /* (1, 10, 1) {real, imag} */,
  {32'h412315d6, 32'hc13078b8} /* (1, 10, 0) {real, imag} */,
  {32'h3fd0a38e, 32'hc09b34a7} /* (1, 9, 31) {real, imag} */,
  {32'hc00d3efe, 32'hbfd998e4} /* (1, 9, 30) {real, imag} */,
  {32'hc1767e7d, 32'hc07a8ea6} /* (1, 9, 29) {real, imag} */,
  {32'hc121b423, 32'hc092de3b} /* (1, 9, 28) {real, imag} */,
  {32'hc12529ea, 32'h3fe7d6f8} /* (1, 9, 27) {real, imag} */,
  {32'hc0e62e30, 32'h410a4139} /* (1, 9, 26) {real, imag} */,
  {32'hc0e18df5, 32'h41b2265d} /* (1, 9, 25) {real, imag} */,
  {32'hbf94989c, 32'h410388b5} /* (1, 9, 24) {real, imag} */,
  {32'hc0da64ce, 32'h40697ac0} /* (1, 9, 23) {real, imag} */,
  {32'hc172da21, 32'hc1306ae4} /* (1, 9, 22) {real, imag} */,
  {32'hc1063fb6, 32'hc112b70e} /* (1, 9, 21) {real, imag} */,
  {32'hc126ab4a, 32'hc025df88} /* (1, 9, 20) {real, imag} */,
  {32'hc13cb772, 32'h403c5008} /* (1, 9, 19) {real, imag} */,
  {32'hc18c2780, 32'h407f3128} /* (1, 9, 18) {real, imag} */,
  {32'hc1a1df48, 32'hc0364fc6} /* (1, 9, 17) {real, imag} */,
  {32'hc11335d7, 32'hc0d9b07e} /* (1, 9, 16) {real, imag} */,
  {32'hc0836766, 32'hc0f6440b} /* (1, 9, 15) {real, imag} */,
  {32'hc052d51a, 32'hbfa657a2} /* (1, 9, 14) {real, imag} */,
  {32'hc16273cc, 32'h411e0320} /* (1, 9, 13) {real, imag} */,
  {32'hc1d5b3d2, 32'h41238b68} /* (1, 9, 12) {real, imag} */,
  {32'hc18dd168, 32'h415bd119} /* (1, 9, 11) {real, imag} */,
  {32'h40a07c16, 32'h40ca1a94} /* (1, 9, 10) {real, imag} */,
  {32'hbf80ac00, 32'hbfbe046c} /* (1, 9, 9) {real, imag} */,
  {32'h4115dcba, 32'h404d6694} /* (1, 9, 8) {real, imag} */,
  {32'hc0decd58, 32'h401db6e2} /* (1, 9, 7) {real, imag} */,
  {32'h40d946b3, 32'h4147582e} /* (1, 9, 6) {real, imag} */,
  {32'h40eeddc0, 32'h41790867} /* (1, 9, 5) {real, imag} */,
  {32'h4165a0c6, 32'h3fe85528} /* (1, 9, 4) {real, imag} */,
  {32'h4076cd7c, 32'hc1113cf8} /* (1, 9, 3) {real, imag} */,
  {32'hbec81870, 32'h410ec1a8} /* (1, 9, 2) {real, imag} */,
  {32'hc13b5add, 32'h40e5775b} /* (1, 9, 1) {real, imag} */,
  {32'hc0d1ae2a, 32'h3f5b73c0} /* (1, 9, 0) {real, imag} */,
  {32'hc0b22622, 32'h40fc9f30} /* (1, 8, 31) {real, imag} */,
  {32'hc0ff49de, 32'h415fa984} /* (1, 8, 30) {real, imag} */,
  {32'hc0a33159, 32'h417f8343} /* (1, 8, 29) {real, imag} */,
  {32'hc171a93a, 32'h418396e7} /* (1, 8, 28) {real, imag} */,
  {32'hc2067bfa, 32'h402bd71e} /* (1, 8, 27) {real, imag} */,
  {32'hc1fa6152, 32'h40572f27} /* (1, 8, 26) {real, imag} */,
  {32'hc110eaee, 32'h40f31cbe} /* (1, 8, 25) {real, imag} */,
  {32'hbf5a4cf8, 32'h410b3837} /* (1, 8, 24) {real, imag} */,
  {32'hc0adf19e, 32'h41a52f96} /* (1, 8, 23) {real, imag} */,
  {32'hbfcb84b8, 32'h41a6cbd4} /* (1, 8, 22) {real, imag} */,
  {32'hc0af8572, 32'h41366f46} /* (1, 8, 21) {real, imag} */,
  {32'h40f1f307, 32'hc0bb4244} /* (1, 8, 20) {real, imag} */,
  {32'h406e9c02, 32'hc1d9ecc0} /* (1, 8, 19) {real, imag} */,
  {32'h40e4af0e, 32'hc200ba96} /* (1, 8, 18) {real, imag} */,
  {32'h4148f087, 32'hc1896ca4} /* (1, 8, 17) {real, imag} */,
  {32'h3f8fd7d4, 32'hc1a86484} /* (1, 8, 16) {real, imag} */,
  {32'h3fb39ba4, 32'h40bfe1a6} /* (1, 8, 15) {real, imag} */,
  {32'h415db8f4, 32'hc0fb4024} /* (1, 8, 14) {real, imag} */,
  {32'h41cda8b6, 32'hc1a063f0} /* (1, 8, 13) {real, imag} */,
  {32'h40e9a008, 32'hc1e0ee97} /* (1, 8, 12) {real, imag} */,
  {32'hc060d1b8, 32'hc126f0ce} /* (1, 8, 11) {real, imag} */,
  {32'hbedac5cc, 32'h4156c0a5} /* (1, 8, 10) {real, imag} */,
  {32'hc0804604, 32'h420b2ec8} /* (1, 8, 9) {real, imag} */,
  {32'hc16d96f2, 32'h4202dac0} /* (1, 8, 8) {real, imag} */,
  {32'hc1807a0c, 32'h40ab5b68} /* (1, 8, 7) {real, imag} */,
  {32'h401ecf36, 32'h40972674} /* (1, 8, 6) {real, imag} */,
  {32'h416c2462, 32'h41bb3f4b} /* (1, 8, 5) {real, imag} */,
  {32'h411e0c91, 32'h419f52c1} /* (1, 8, 4) {real, imag} */,
  {32'hc182f87e, 32'h40cb3a04} /* (1, 8, 3) {real, imag} */,
  {32'hc1c4dc51, 32'h40c12098} /* (1, 8, 2) {real, imag} */,
  {32'hc1b8ea4b, 32'h40a9cdac} /* (1, 8, 1) {real, imag} */,
  {32'hbfa5aeda, 32'h3fbb277a} /* (1, 8, 0) {real, imag} */,
  {32'h3f3fe594, 32'hc1096c32} /* (1, 7, 31) {real, imag} */,
  {32'h3fb65908, 32'hc11002be} /* (1, 7, 30) {real, imag} */,
  {32'h411609c5, 32'hc039f47e} /* (1, 7, 29) {real, imag} */,
  {32'h40fc1e1c, 32'hc143b4e4} /* (1, 7, 28) {real, imag} */,
  {32'h413016d6, 32'hc1bbb565} /* (1, 7, 27) {real, imag} */,
  {32'h41e55aa3, 32'hc1855a49} /* (1, 7, 26) {real, imag} */,
  {32'h419c9f48, 32'hc12a3ab6} /* (1, 7, 25) {real, imag} */,
  {32'h4183b1e4, 32'hc1a65042} /* (1, 7, 24) {real, imag} */,
  {32'h41208bd0, 32'hc2002c82} /* (1, 7, 23) {real, imag} */,
  {32'h414ee53d, 32'hc1149d24} /* (1, 7, 22) {real, imag} */,
  {32'h4082eff7, 32'h4046d4f0} /* (1, 7, 21) {real, imag} */,
  {32'h404eeb92, 32'h406b9910} /* (1, 7, 20) {real, imag} */,
  {32'h40ad7530, 32'h409d1ec2} /* (1, 7, 19) {real, imag} */,
  {32'hc0c0a5b8, 32'h4099b670} /* (1, 7, 18) {real, imag} */,
  {32'hc1934b02, 32'h40ac3365} /* (1, 7, 17) {real, imag} */,
  {32'hc1aac0bb, 32'h40759cc7} /* (1, 7, 16) {real, imag} */,
  {32'hc1090eac, 32'h41c5181d} /* (1, 7, 15) {real, imag} */,
  {32'hc11c266e, 32'h411623c3} /* (1, 7, 14) {real, imag} */,
  {32'hc0f7ebbd, 32'hc128c5a6} /* (1, 7, 13) {real, imag} */,
  {32'h403165d4, 32'h4109ce48} /* (1, 7, 12) {real, imag} */,
  {32'hc01e6f2c, 32'h41b46122} /* (1, 7, 11) {real, imag} */,
  {32'h411f9d06, 32'h41582e26} /* (1, 7, 10) {real, imag} */,
  {32'h410faf94, 32'hbf2efc98} /* (1, 7, 9) {real, imag} */,
  {32'h411bf8aa, 32'h415f90a7} /* (1, 7, 8) {real, imag} */,
  {32'h41c911c5, 32'hc0cbebc9} /* (1, 7, 7) {real, imag} */,
  {32'h4178157f, 32'hc1d80063} /* (1, 7, 6) {real, imag} */,
  {32'h413461d9, 32'hc0c7bffe} /* (1, 7, 5) {real, imag} */,
  {32'h41c7177e, 32'h40087344} /* (1, 7, 4) {real, imag} */,
  {32'h40952569, 32'hc13043f4} /* (1, 7, 3) {real, imag} */,
  {32'h401a2142, 32'h407a8d4e} /* (1, 7, 2) {real, imag} */,
  {32'h4145e2da, 32'h418614ba} /* (1, 7, 1) {real, imag} */,
  {32'h4142661f, 32'h40c68f0c} /* (1, 7, 0) {real, imag} */,
  {32'h40ea4502, 32'h3dd62660} /* (1, 6, 31) {real, imag} */,
  {32'hc0a1ada8, 32'h3feea514} /* (1, 6, 30) {real, imag} */,
  {32'hc070c338, 32'hbf84d5d4} /* (1, 6, 29) {real, imag} */,
  {32'h3f17ac60, 32'hc044794d} /* (1, 6, 28) {real, imag} */,
  {32'hbf9e7198, 32'h3f65d360} /* (1, 6, 27) {real, imag} */,
  {32'hc03020c1, 32'hc0b3844a} /* (1, 6, 26) {real, imag} */,
  {32'h41437266, 32'hc08855d9} /* (1, 6, 25) {real, imag} */,
  {32'h41b67ae4, 32'h3f9519d0} /* (1, 6, 24) {real, imag} */,
  {32'hc072741e, 32'hc1135c05} /* (1, 6, 23) {real, imag} */,
  {32'hbf78e278, 32'hc0ebe304} /* (1, 6, 22) {real, imag} */,
  {32'h408d59d4, 32'hc0aa5944} /* (1, 6, 21) {real, imag} */,
  {32'h41bfbdfa, 32'hc0c73be6} /* (1, 6, 20) {real, imag} */,
  {32'h40e7dc2e, 32'h4138069f} /* (1, 6, 19) {real, imag} */,
  {32'h4016889c, 32'h408e2be2} /* (1, 6, 18) {real, imag} */,
  {32'h41051f86, 32'hc1390a53} /* (1, 6, 17) {real, imag} */,
  {32'hc11abb0c, 32'h403b2b3e} /* (1, 6, 16) {real, imag} */,
  {32'hc19b061d, 32'hc0a33bd2} /* (1, 6, 15) {real, imag} */,
  {32'h411a3b34, 32'hc174c23e} /* (1, 6, 14) {real, imag} */,
  {32'h40c257e4, 32'hc1314dcd} /* (1, 6, 13) {real, imag} */,
  {32'h41178d80, 32'hbd2d9b00} /* (1, 6, 12) {real, imag} */,
  {32'h4164af7e, 32'h4182a3a1} /* (1, 6, 11) {real, imag} */,
  {32'h421f9a50, 32'h407db4fa} /* (1, 6, 10) {real, imag} */,
  {32'h4200f6e6, 32'hc0e1c4b6} /* (1, 6, 9) {real, imag} */,
  {32'h40858d85, 32'h3f3b42dc} /* (1, 6, 8) {real, imag} */,
  {32'h410b5d34, 32'hc0edbcc5} /* (1, 6, 7) {real, imag} */,
  {32'h411b4a51, 32'hc1ad1783} /* (1, 6, 6) {real, imag} */,
  {32'h413dd7b3, 32'hbff32974} /* (1, 6, 5) {real, imag} */,
  {32'h40c64f5c, 32'h411fbb1e} /* (1, 6, 4) {real, imag} */,
  {32'hc1078c80, 32'hc143b7a6} /* (1, 6, 3) {real, imag} */,
  {32'hc1baae5c, 32'h4085bb88} /* (1, 6, 2) {real, imag} */,
  {32'hc12059d2, 32'h40e4fdfd} /* (1, 6, 1) {real, imag} */,
  {32'h405b8267, 32'hbe36b280} /* (1, 6, 0) {real, imag} */,
  {32'h400d33da, 32'h40bd5acc} /* (1, 5, 31) {real, imag} */,
  {32'h3ea409e0, 32'h41bdb412} /* (1, 5, 30) {real, imag} */,
  {32'hc1615429, 32'h41a5fc8c} /* (1, 5, 29) {real, imag} */,
  {32'hc18d6fb5, 32'h413cb47e} /* (1, 5, 28) {real, imag} */,
  {32'hc19493d1, 32'h412bee06} /* (1, 5, 27) {real, imag} */,
  {32'hc18cf76c, 32'h4110de75} /* (1, 5, 26) {real, imag} */,
  {32'hc1b64839, 32'h40ea21a8} /* (1, 5, 25) {real, imag} */,
  {32'hc23e2517, 32'h41ca3f2a} /* (1, 5, 24) {real, imag} */,
  {32'hc24dba10, 32'h424556a9} /* (1, 5, 23) {real, imag} */,
  {32'hc1a3d7fc, 32'h42349a9e} /* (1, 5, 22) {real, imag} */,
  {32'hc0cfa437, 32'h4204fc8f} /* (1, 5, 21) {real, imag} */,
  {32'hbf1ec3b0, 32'hc0e18dd0} /* (1, 5, 20) {real, imag} */,
  {32'hbf85a454, 32'hc1444050} /* (1, 5, 19) {real, imag} */,
  {32'h40f82ed6, 32'hc17fe174} /* (1, 5, 18) {real, imag} */,
  {32'h416dbf78, 32'hc16001ce} /* (1, 5, 17) {real, imag} */,
  {32'h4182ef04, 32'hc15f786d} /* (1, 5, 16) {real, imag} */,
  {32'h41aa8741, 32'hc1df378e} /* (1, 5, 15) {real, imag} */,
  {32'h41fa6eee, 32'hc1873b9d} /* (1, 5, 14) {real, imag} */,
  {32'h41f3de83, 32'hc1b61ad8} /* (1, 5, 13) {real, imag} */,
  {32'h41a7e69b, 32'hc208a722} /* (1, 5, 12) {real, imag} */,
  {32'h406d21f8, 32'hc22053a6} /* (1, 5, 11) {real, imag} */,
  {32'h410a32d2, 32'hc130f867} /* (1, 5, 10) {real, imag} */,
  {32'hc189ebfc, 32'hc03f68f0} /* (1, 5, 9) {real, imag} */,
  {32'hc1f83047, 32'h40da710e} /* (1, 5, 8) {real, imag} */,
  {32'hc17d8588, 32'h411e5f5a} /* (1, 5, 7) {real, imag} */,
  {32'hc13b96c0, 32'hbfb34134} /* (1, 5, 6) {real, imag} */,
  {32'hc11b634a, 32'h4212d4fe} /* (1, 5, 5) {real, imag} */,
  {32'hc19c34ef, 32'h42260dd3} /* (1, 5, 4) {real, imag} */,
  {32'hc0d0fa61, 32'h41d0677a} /* (1, 5, 3) {real, imag} */,
  {32'hc1972495, 32'hbfe32eb0} /* (1, 5, 2) {real, imag} */,
  {32'hc0829490, 32'h4083e708} /* (1, 5, 1) {real, imag} */,
  {32'hc0b16873, 32'h404c6af8} /* (1, 5, 0) {real, imag} */,
  {32'h417dff7e, 32'h40b7f397} /* (1, 4, 31) {real, imag} */,
  {32'h4181af8f, 32'h3fb9dd78} /* (1, 4, 30) {real, imag} */,
  {32'hc175d663, 32'hbfb9fc50} /* (1, 4, 29) {real, imag} */,
  {32'hc1ad4156, 32'hc1880d6e} /* (1, 4, 28) {real, imag} */,
  {32'h3f88beb0, 32'hc1fa3950} /* (1, 4, 27) {real, imag} */,
  {32'h40f00718, 32'hc209bbdb} /* (1, 4, 26) {real, imag} */,
  {32'hc0a4da7c, 32'h40466b54} /* (1, 4, 25) {real, imag} */,
  {32'h404ae768, 32'hc1808fb3} /* (1, 4, 24) {real, imag} */,
  {32'h41e0838e, 32'hc15c3074} /* (1, 4, 23) {real, imag} */,
  {32'h4264b70e, 32'hc17575ca} /* (1, 4, 22) {real, imag} */,
  {32'h41830f0f, 32'hbfc19d20} /* (1, 4, 21) {real, imag} */,
  {32'hc223975a, 32'h420aa884} /* (1, 4, 20) {real, imag} */,
  {32'hc22da810, 32'h41d7a294} /* (1, 4, 19) {real, imag} */,
  {32'hc215310b, 32'h406ced88} /* (1, 4, 18) {real, imag} */,
  {32'hc1a8012d, 32'h41a1d1de} /* (1, 4, 17) {real, imag} */,
  {32'hc1b55dab, 32'h41dbc16c} /* (1, 4, 16) {real, imag} */,
  {32'hc1adc1aa, 32'h416bf6c3} /* (1, 4, 15) {real, imag} */,
  {32'hc127c946, 32'h4140849e} /* (1, 4, 14) {real, imag} */,
  {32'hc12af2c3, 32'h41cbc48f} /* (1, 4, 13) {real, imag} */,
  {32'hc1c8d82f, 32'h41e0ba84} /* (1, 4, 12) {real, imag} */,
  {32'h41188ee6, 32'h3fcdcb9e} /* (1, 4, 11) {real, imag} */,
  {32'h4207f3a7, 32'hc2311cf0} /* (1, 4, 10) {real, imag} */,
  {32'h41ef0d40, 32'hc23438c8} /* (1, 4, 9) {real, imag} */,
  {32'h428a181b, 32'hc22bfbf7} /* (1, 4, 8) {real, imag} */,
  {32'h42563f2b, 32'hc276ee96} /* (1, 4, 7) {real, imag} */,
  {32'h426d91ae, 32'hc26d1409} /* (1, 4, 6) {real, imag} */,
  {32'h41ca48be, 32'hc1d28aff} /* (1, 4, 5) {real, imag} */,
  {32'hc1a0e22c, 32'hc0ff53d7} /* (1, 4, 4) {real, imag} */,
  {32'hbfd7a58c, 32'h404a9094} /* (1, 4, 3) {real, imag} */,
  {32'h41854dcc, 32'h419612d2} /* (1, 4, 2) {real, imag} */,
  {32'h41026dee, 32'h41b3bfe6} /* (1, 4, 1) {real, imag} */,
  {32'h3fd3a2ee, 32'h4187ab40} /* (1, 4, 0) {real, imag} */,
  {32'hc0ef184e, 32'h41887645} /* (1, 3, 31) {real, imag} */,
  {32'h40f9ebbf, 32'h411dcb0a} /* (1, 3, 30) {real, imag} */,
  {32'h4149c529, 32'h40706db0} /* (1, 3, 29) {real, imag} */,
  {32'h410483e0, 32'hc0ff0f34} /* (1, 3, 28) {real, imag} */,
  {32'h4082db24, 32'hc11dd578} /* (1, 3, 27) {real, imag} */,
  {32'hbfde363e, 32'h40413e52} /* (1, 3, 26) {real, imag} */,
  {32'h40381548, 32'h41d5397c} /* (1, 3, 25) {real, imag} */,
  {32'h40b5bfa1, 32'h40bf77cd} /* (1, 3, 24) {real, imag} */,
  {32'h4118829f, 32'hc108068b} /* (1, 3, 23) {real, imag} */,
  {32'h40c4a370, 32'h41377428} /* (1, 3, 22) {real, imag} */,
  {32'hc13f4ccc, 32'h413c1883} /* (1, 3, 21) {real, imag} */,
  {32'hc24d58c3, 32'h3f3b9010} /* (1, 3, 20) {real, imag} */,
  {32'hc2400e24, 32'h3f6775a8} /* (1, 3, 19) {real, imag} */,
  {32'hc25b540a, 32'hc0cf3f95} /* (1, 3, 18) {real, imag} */,
  {32'hc2166738, 32'hc1a075d6} /* (1, 3, 17) {real, imag} */,
  {32'hc248a0fc, 32'hc134872d} /* (1, 3, 16) {real, imag} */,
  {32'hc1eb8103, 32'hc1a2b421} /* (1, 3, 15) {real, imag} */,
  {32'h40a71ad6, 32'hc138d66a} /* (1, 3, 14) {real, imag} */,
  {32'h41f90dd3, 32'hc0b4693c} /* (1, 3, 13) {real, imag} */,
  {32'hbfb64978, 32'h3f85ee40} /* (1, 3, 12) {real, imag} */,
  {32'h40b2a7c2, 32'hc1264c02} /* (1, 3, 11) {real, imag} */,
  {32'h41f1a839, 32'h40b57942} /* (1, 3, 10) {real, imag} */,
  {32'h41db6d67, 32'h42041e62} /* (1, 3, 9) {real, imag} */,
  {32'h42841cd5, 32'h41fbb6c3} /* (1, 3, 8) {real, imag} */,
  {32'h429dc03b, 32'h4126d68c} /* (1, 3, 7) {real, imag} */,
  {32'h424d7ceb, 32'h40a40e34} /* (1, 3, 6) {real, imag} */,
  {32'h408101ec, 32'h41a24f00} /* (1, 3, 5) {real, imag} */,
  {32'hc10af819, 32'h41a09f9e} /* (1, 3, 4) {real, imag} */,
  {32'hc16771e1, 32'h408f6212} /* (1, 3, 3) {real, imag} */,
  {32'hc19cd39c, 32'hc12a537e} /* (1, 3, 2) {real, imag} */,
  {32'hbe76fe30, 32'hc0802b16} /* (1, 3, 1) {real, imag} */,
  {32'hc0809e1e, 32'h3f3fa12c} /* (1, 3, 0) {real, imag} */,
  {32'hc196be52, 32'h425aab34} /* (1, 2, 31) {real, imag} */,
  {32'hc1a6fa74, 32'h4290eaae} /* (1, 2, 30) {real, imag} */,
  {32'hc10b8762, 32'h42a83a69} /* (1, 2, 29) {real, imag} */,
  {32'hc1a46e1f, 32'h42d06674} /* (1, 2, 28) {real, imag} */,
  {32'hc2049e5a, 32'h42bbfb78} /* (1, 2, 27) {real, imag} */,
  {32'hc15e47d8, 32'h427dd97d} /* (1, 2, 26) {real, imag} */,
  {32'hc18ccf70, 32'h428922f7} /* (1, 2, 25) {real, imag} */,
  {32'hc2131943, 32'h42ce78d2} /* (1, 2, 24) {real, imag} */,
  {32'hc23e8b34, 32'h42d075bc} /* (1, 2, 23) {real, imag} */,
  {32'hc1a8b0fc, 32'h427db5cf} /* (1, 2, 22) {real, imag} */,
  {32'hc1b3d17b, 32'h41455c01} /* (1, 2, 21) {real, imag} */,
  {32'hc2117aca, 32'hc2bf3025} /* (1, 2, 20) {real, imag} */,
  {32'hc1da3596, 32'hc2e4cccc} /* (1, 2, 19) {real, imag} */,
  {32'hc22f2632, 32'hc30489ff} /* (1, 2, 18) {real, imag} */,
  {32'hc205e2b0, 32'hc30853db} /* (1, 2, 17) {real, imag} */,
  {32'hc1e3b001, 32'hc2e74e52} /* (1, 2, 16) {real, imag} */,
  {32'h41c7121e, 32'hc2a98dd8} /* (1, 2, 15) {real, imag} */,
  {32'h423b7a8e, 32'hc2b66c97} /* (1, 2, 14) {real, imag} */,
  {32'h422009c4, 32'hc2db15e6} /* (1, 2, 13) {real, imag} */,
  {32'h42246dba, 32'hc2c476a5} /* (1, 2, 12) {real, imag} */,
  {32'h41e283c3, 32'hc263cafb} /* (1, 2, 11) {real, imag} */,
  {32'h402a72a0, 32'h421f03eb} /* (1, 2, 10) {real, imag} */,
  {32'h412752e8, 32'h42f25087} /* (1, 2, 9) {real, imag} */,
  {32'h41e3d9a0, 32'h4313f1fb} /* (1, 2, 8) {real, imag} */,
  {32'h42202803, 32'h430df5cc} /* (1, 2, 7) {real, imag} */,
  {32'h41f848d0, 32'h42f0f6b8} /* (1, 2, 6) {real, imag} */,
  {32'hc197c372, 32'h42a8a05e} /* (1, 2, 5) {real, imag} */,
  {32'hc22649fa, 32'h42b9f17d} /* (1, 2, 4) {real, imag} */,
  {32'hc1ceea9a, 32'h42b2913a} /* (1, 2, 3) {real, imag} */,
  {32'hc1e717c2, 32'h42986ed6} /* (1, 2, 2) {real, imag} */,
  {32'hc1c09834, 32'h42bc85d9} /* (1, 2, 1) {real, imag} */,
  {32'hc0f50d38, 32'h4283c5a3} /* (1, 2, 0) {real, imag} */,
  {32'h41b84144, 32'hc29c8b2e} /* (1, 1, 31) {real, imag} */,
  {32'h421ef9aa, 32'hc3170863} /* (1, 1, 30) {real, imag} */,
  {32'h419d04cc, 32'hc3126c82} /* (1, 1, 29) {real, imag} */,
  {32'h415d2832, 32'hc303574d} /* (1, 1, 28) {real, imag} */,
  {32'h3fd8a854, 32'hc2fbc35e} /* (1, 1, 27) {real, imag} */,
  {32'h418082ad, 32'hc2df4762} /* (1, 1, 26) {real, imag} */,
  {32'h422a5a2e, 32'hc2fd44d5} /* (1, 1, 25) {real, imag} */,
  {32'h422ec80e, 32'hc31ace5e} /* (1, 1, 24) {real, imag} */,
  {32'h41420e25, 32'hc31b9a4c} /* (1, 1, 23) {real, imag} */,
  {32'h410eec99, 32'hc2fed6a2} /* (1, 1, 22) {real, imag} */,
  {32'h41061cb8, 32'hc2778c03} /* (1, 1, 21) {real, imag} */,
  {32'hc24dcc36, 32'h4229ca6d} /* (1, 1, 20) {real, imag} */,
  {32'hc28b386e, 32'h4266187a} /* (1, 1, 19) {real, imag} */,
  {32'hc2665d5d, 32'h4271c469} /* (1, 1, 18) {real, imag} */,
  {32'hc23e4527, 32'h428f2594} /* (1, 1, 17) {real, imag} */,
  {32'hc24c0b07, 32'h42bbaa91} /* (1, 1, 16) {real, imag} */,
  {32'hc190d2f4, 32'h42e51a46} /* (1, 1, 15) {real, imag} */,
  {32'hc218614d, 32'h42e61019} /* (1, 1, 14) {real, imag} */,
  {32'hc24b2984, 32'h42f9e394} /* (1, 1, 13) {real, imag} */,
  {32'hc2061259, 32'h430826b4} /* (1, 1, 12) {real, imag} */,
  {32'hc187b659, 32'h4303922a} /* (1, 1, 11) {real, imag} */,
  {32'h42287f72, 32'h41294f4c} /* (1, 1, 10) {real, imag} */,
  {32'h42ca9c10, 32'hc26a182e} /* (1, 1, 9) {real, imag} */,
  {32'h42c21df0, 32'hc218fe56} /* (1, 1, 8) {real, imag} */,
  {32'h4287b874, 32'hc21da96f} /* (1, 1, 7) {real, imag} */,
  {32'h4218ccd4, 32'hc262d55e} /* (1, 1, 6) {real, imag} */,
  {32'h41f2b67d, 32'hc2b7ac64} /* (1, 1, 5) {real, imag} */,
  {32'h4216e63a, 32'hc3067489} /* (1, 1, 4) {real, imag} */,
  {32'h42019c2c, 32'hc2ef828b} /* (1, 1, 3) {real, imag} */,
  {32'h420633a7, 32'hc2ef28d2} /* (1, 1, 2) {real, imag} */,
  {32'h41ccbd27, 32'hc3108882} /* (1, 1, 1) {real, imag} */,
  {32'h40e97085, 32'hc2b8c586} /* (1, 1, 0) {real, imag} */,
  {32'h4131d7af, 32'hc221f908} /* (1, 0, 31) {real, imag} */,
  {32'h41ade2fd, 32'hc291ba95} /* (1, 0, 30) {real, imag} */,
  {32'h4106fe6c, 32'hc2c4cd4f} /* (1, 0, 29) {real, imag} */,
  {32'hc1358670, 32'hc2bf6c40} /* (1, 0, 28) {real, imag} */,
  {32'h3fa5a3a8, 32'hc2b1ea37} /* (1, 0, 27) {real, imag} */,
  {32'h406ec97f, 32'hc294b312} /* (1, 0, 26) {real, imag} */,
  {32'h40d7c44d, 32'hc2ae4994} /* (1, 0, 25) {real, imag} */,
  {32'hc0111d99, 32'hc296804d} /* (1, 0, 24) {real, imag} */,
  {32'h41b1b26c, 32'hc293a006} /* (1, 0, 23) {real, imag} */,
  {32'h416f4f02, 32'hc2bd0aa4} /* (1, 0, 22) {real, imag} */,
  {32'h4158225e, 32'hc2ac5ade} /* (1, 0, 21) {real, imag} */,
  {32'h40fcf7fd, 32'hc1b5040d} /* (1, 0, 20) {real, imag} */,
  {32'h4117ec6a, 32'hc0889871} /* (1, 0, 19) {real, imag} */,
  {32'h40d30719, 32'h4164ad78} /* (1, 0, 18) {real, imag} */,
  {32'hbfaaba1c, 32'hc0b09712} /* (1, 0, 17) {real, imag} */,
  {32'hc1031170, 32'h41cd91ff} /* (1, 0, 16) {real, imag} */,
  {32'hc1a218fc, 32'h429c0335} /* (1, 0, 15) {real, imag} */,
  {32'hc1c0fcf2, 32'h42b73143} /* (1, 0, 14) {real, imag} */,
  {32'hc1802526, 32'h42a4a3c1} /* (1, 0, 13) {real, imag} */,
  {32'hc106f944, 32'h4297793c} /* (1, 0, 12) {real, imag} */,
  {32'hc0c83fa6, 32'h42830347} /* (1, 0, 11) {real, imag} */,
  {32'hbfa9e2f8, 32'h4186c7e6} /* (1, 0, 10) {real, imag} */,
  {32'hc15a7420, 32'h414740c4} /* (1, 0, 9) {real, imag} */,
  {32'hc18bf2f1, 32'h40bd627b} /* (1, 0, 8) {real, imag} */,
  {32'h41b78cc2, 32'h4110edda} /* (1, 0, 7) {real, imag} */,
  {32'h41c1723c, 32'h41229046} /* (1, 0, 6) {real, imag} */,
  {32'hc004e60d, 32'hc27e06d4} /* (1, 0, 5) {real, imag} */,
  {32'h40bf0006, 32'hc29f4ae0} /* (1, 0, 4) {real, imag} */,
  {32'h403ccbe8, 32'hc2a7323e} /* (1, 0, 3) {real, imag} */,
  {32'h41141feb, 32'hc29c6652} /* (1, 0, 2) {real, imag} */,
  {32'h410ee7c4, 32'hc2ae22c6} /* (1, 0, 1) {real, imag} */,
  {32'h4103450e, 32'hc2122467} /* (1, 0, 0) {real, imag} */,
  {32'hc03cbde5, 32'hc04160be} /* (0, 31, 31) {real, imag} */,
  {32'h3fbe9f02, 32'hc182326f} /* (0, 31, 30) {real, imag} */,
  {32'hc1855454, 32'hc144e5c8} /* (0, 31, 29) {real, imag} */,
  {32'hc127b75c, 32'hbfcd4dc6} /* (0, 31, 28) {real, imag} */,
  {32'h4141b6bb, 32'h414379ed} /* (0, 31, 27) {real, imag} */,
  {32'hc0efa0ea, 32'hc04a22d4} /* (0, 31, 26) {real, imag} */,
  {32'h408bf19e, 32'hc1d10244} /* (0, 31, 25) {real, imag} */,
  {32'h4136907c, 32'hc09ef32c} /* (0, 31, 24) {real, imag} */,
  {32'hc0e8f0eb, 32'h419444af} /* (0, 31, 23) {real, imag} */,
  {32'hc005942e, 32'h42195d50} /* (0, 31, 22) {real, imag} */,
  {32'h40d1e47e, 32'h40b23444} /* (0, 31, 21) {real, imag} */,
  {32'h41801916, 32'hc030fe69} /* (0, 31, 20) {real, imag} */,
  {32'h41afecac, 32'hc1cdacca} /* (0, 31, 19) {real, imag} */,
  {32'hc1161778, 32'hc1b001be} /* (0, 31, 18) {real, imag} */,
  {32'h4115cf1b, 32'h40a981f9} /* (0, 31, 17) {real, imag} */,
  {32'hc10424c2, 32'h41a3817a} /* (0, 31, 16) {real, imag} */,
  {32'hc1c87c3b, 32'hbcdf7e80} /* (0, 31, 15) {real, imag} */,
  {32'hc14854e8, 32'hc103f10c} /* (0, 31, 14) {real, imag} */,
  {32'hc057a3c1, 32'hc12b409e} /* (0, 31, 13) {real, imag} */,
  {32'h40c0fb56, 32'hc0f84b20} /* (0, 31, 12) {real, imag} */,
  {32'h4168fbd2, 32'hc0f00422} /* (0, 31, 11) {real, imag} */,
  {32'h40f23c4d, 32'h4133471a} /* (0, 31, 10) {real, imag} */,
  {32'hc15fe4aa, 32'hc17cf879} /* (0, 31, 9) {real, imag} */,
  {32'hc0938b7c, 32'h415a9780} /* (0, 31, 8) {real, imag} */,
  {32'h40970fd8, 32'h41f0396d} /* (0, 31, 7) {real, imag} */,
  {32'h4190a623, 32'hc1429bc0} /* (0, 31, 6) {real, imag} */,
  {32'h410ae361, 32'hc104233a} /* (0, 31, 5) {real, imag} */,
  {32'h3ed93a18, 32'h40a2a322} /* (0, 31, 4) {real, imag} */,
  {32'h4180b90c, 32'h3eee7f90} /* (0, 31, 3) {real, imag} */,
  {32'h400876e8, 32'h40a4c4e7} /* (0, 31, 2) {real, imag} */,
  {32'hc09d8cb4, 32'h41d62eb4} /* (0, 31, 1) {real, imag} */,
  {32'h407ea3c4, 32'h41728da4} /* (0, 31, 0) {real, imag} */,
  {32'hbdbfd7b0, 32'hc0afeae7} /* (0, 30, 31) {real, imag} */,
  {32'hc1805a84, 32'hbf44cd40} /* (0, 30, 30) {real, imag} */,
  {32'hc1087efe, 32'hc19112ec} /* (0, 30, 29) {real, imag} */,
  {32'h40afda84, 32'hc12466c3} /* (0, 30, 28) {real, imag} */,
  {32'hbeb3e640, 32'h3fa65702} /* (0, 30, 27) {real, imag} */,
  {32'h4081ace9, 32'hc0a333b0} /* (0, 30, 26) {real, imag} */,
  {32'h412df720, 32'h40e52612} /* (0, 30, 25) {real, imag} */,
  {32'h413f5fb4, 32'h41913c3c} /* (0, 30, 24) {real, imag} */,
  {32'hbeeed2b4, 32'h4055c944} /* (0, 30, 23) {real, imag} */,
  {32'hc17b7863, 32'hc0eaea8a} /* (0, 30, 22) {real, imag} */,
  {32'h41188d67, 32'h3fc928ac} /* (0, 30, 21) {real, imag} */,
  {32'hc151b16d, 32'h408d3256} /* (0, 30, 20) {real, imag} */,
  {32'hc193032c, 32'h411581e2} /* (0, 30, 19) {real, imag} */,
  {32'h3fef19c2, 32'h3fd054d0} /* (0, 30, 18) {real, imag} */,
  {32'h3f89e3e4, 32'hc06f03b0} /* (0, 30, 17) {real, imag} */,
  {32'h4164baea, 32'hc089dac0} /* (0, 30, 16) {real, imag} */,
  {32'h3f937da6, 32'h405434fa} /* (0, 30, 15) {real, imag} */,
  {32'h3e831acc, 32'h41fe050b} /* (0, 30, 14) {real, imag} */,
  {32'h400017e3, 32'h4203a35e} /* (0, 30, 13) {real, imag} */,
  {32'hc161fd96, 32'hc107b250} /* (0, 30, 12) {real, imag} */,
  {32'h401b8e9c, 32'hc1fee6d2} /* (0, 30, 11) {real, imag} */,
  {32'h419aaa82, 32'hc194d4b9} /* (0, 30, 10) {real, imag} */,
  {32'h419e8bfd, 32'h417ad3e1} /* (0, 30, 9) {real, imag} */,
  {32'hc16ee821, 32'h3ee6a150} /* (0, 30, 8) {real, imag} */,
  {32'hc24253e4, 32'h3f875007} /* (0, 30, 7) {real, imag} */,
  {32'hc1a3d3fc, 32'h40a9909b} /* (0, 30, 6) {real, imag} */,
  {32'hc12f17d2, 32'hc102efaa} /* (0, 30, 5) {real, imag} */,
  {32'hc144ac48, 32'hc13b53e6} /* (0, 30, 4) {real, imag} */,
  {32'hc113a294, 32'hc0171f79} /* (0, 30, 3) {real, imag} */,
  {32'h412ef954, 32'h41a78a2a} /* (0, 30, 2) {real, imag} */,
  {32'h418a76fb, 32'h40224890} /* (0, 30, 1) {real, imag} */,
  {32'h41742e1c, 32'hc08d7124} /* (0, 30, 0) {real, imag} */,
  {32'h3f845e4c, 32'hc14452b0} /* (0, 29, 31) {real, imag} */,
  {32'h4223fb08, 32'hc12f8dbf} /* (0, 29, 30) {real, imag} */,
  {32'h41ccc5e8, 32'h411a5b66} /* (0, 29, 29) {real, imag} */,
  {32'h40fd5c33, 32'h412384ce} /* (0, 29, 28) {real, imag} */,
  {32'h409dd54a, 32'hbea5e4f0} /* (0, 29, 27) {real, imag} */,
  {32'hc1315f28, 32'h4111cac8} /* (0, 29, 26) {real, imag} */,
  {32'h41e905a8, 32'hc08415a1} /* (0, 29, 25) {real, imag} */,
  {32'h422cfdb8, 32'hc144ae7a} /* (0, 29, 24) {real, imag} */,
  {32'h419de178, 32'hc16fc3ae} /* (0, 29, 23) {real, imag} */,
  {32'h403f4b3e, 32'h40ffa333} /* (0, 29, 22) {real, imag} */,
  {32'hc1a0628e, 32'h41ce70d0} /* (0, 29, 21) {real, imag} */,
  {32'hc1223295, 32'h4115d7af} /* (0, 29, 20) {real, imag} */,
  {32'h40a6e4e4, 32'hc1a0cfce} /* (0, 29, 19) {real, imag} */,
  {32'h40170e5d, 32'h3fc69c4b} /* (0, 29, 18) {real, imag} */,
  {32'h40027d90, 32'hc0f8310f} /* (0, 29, 17) {real, imag} */,
  {32'h419e46e6, 32'hc1acde76} /* (0, 29, 16) {real, imag} */,
  {32'h418575dd, 32'hc18b41cb} /* (0, 29, 15) {real, imag} */,
  {32'h40d18d4c, 32'h4003b8f8} /* (0, 29, 14) {real, imag} */,
  {32'h412df48a, 32'h4102cfe7} /* (0, 29, 13) {real, imag} */,
  {32'h4034f920, 32'hc11cbbc2} /* (0, 29, 12) {real, imag} */,
  {32'h41ae9522, 32'hc05f6144} /* (0, 29, 11) {real, imag} */,
  {32'hc00656fc, 32'hc0d22b4c} /* (0, 29, 10) {real, imag} */,
  {32'hc1645fd0, 32'h3fa2ef50} /* (0, 29, 9) {real, imag} */,
  {32'hc1871ce6, 32'h419d4b0a} /* (0, 29, 8) {real, imag} */,
  {32'hc0da7b3a, 32'h40601197} /* (0, 29, 7) {real, imag} */,
  {32'h41283fc5, 32'hc0748c28} /* (0, 29, 6) {real, imag} */,
  {32'hc1422ef2, 32'h3ea56470} /* (0, 29, 5) {real, imag} */,
  {32'hc10e5ad6, 32'h3cdbd180} /* (0, 29, 4) {real, imag} */,
  {32'h40f0b142, 32'h402e9b4e} /* (0, 29, 3) {real, imag} */,
  {32'h4178fa53, 32'hbf9712e1} /* (0, 29, 2) {real, imag} */,
  {32'hc0baff95, 32'hc1a5939d} /* (0, 29, 1) {real, imag} */,
  {32'hc1234a3c, 32'hc0d5e75c} /* (0, 29, 0) {real, imag} */,
  {32'h3fe4278d, 32'h418ab184} /* (0, 28, 31) {real, imag} */,
  {32'hbf9d3dfa, 32'h41281684} /* (0, 28, 30) {real, imag} */,
  {32'h41214547, 32'h41993c21} /* (0, 28, 29) {real, imag} */,
  {32'hc1050e7c, 32'h41dab762} /* (0, 28, 28) {real, imag} */,
  {32'hc11d6cd5, 32'hbfe08885} /* (0, 28, 27) {real, imag} */,
  {32'hc0a4d6c8, 32'hc112e86f} /* (0, 28, 26) {real, imag} */,
  {32'h4194035e, 32'h421724fc} /* (0, 28, 25) {real, imag} */,
  {32'h41e5961c, 32'h4200bfe7} /* (0, 28, 24) {real, imag} */,
  {32'hc0fe57af, 32'hc1b613a9} /* (0, 28, 23) {real, imag} */,
  {32'hc1f1da8a, 32'hc162fd40} /* (0, 28, 22) {real, imag} */,
  {32'hc19e793c, 32'hc0b2a095} /* (0, 28, 21) {real, imag} */,
  {32'h41bda67d, 32'h4032718e} /* (0, 28, 20) {real, imag} */,
  {32'h41bdf304, 32'hc0496e74} /* (0, 28, 19) {real, imag} */,
  {32'hc09b137a, 32'hc1f4b8a4} /* (0, 28, 18) {real, imag} */,
  {32'hc09b5a2a, 32'hc146f779} /* (0, 28, 17) {real, imag} */,
  {32'h3dd7aad0, 32'hc08a2389} /* (0, 28, 16) {real, imag} */,
  {32'h41509f16, 32'hc0bcafdb} /* (0, 28, 15) {real, imag} */,
  {32'h3e8214f9, 32'h41bc236e} /* (0, 28, 14) {real, imag} */,
  {32'hc1e63c7a, 32'h41b084bc} /* (0, 28, 13) {real, imag} */,
  {32'hc1fce31d, 32'h41569ec6} /* (0, 28, 12) {real, imag} */,
  {32'hc1a86b7c, 32'h415050ec} /* (0, 28, 11) {real, imag} */,
  {32'hc1e57d3a, 32'hc1511fcf} /* (0, 28, 10) {real, imag} */,
  {32'hbfe9fd4a, 32'hbf08e0fc} /* (0, 28, 9) {real, imag} */,
  {32'h3fefbb65, 32'h3f631dff} /* (0, 28, 8) {real, imag} */,
  {32'h40bada07, 32'h41b83ebe} /* (0, 28, 7) {real, imag} */,
  {32'hc0f97d26, 32'h414625f5} /* (0, 28, 6) {real, imag} */,
  {32'hc189b4df, 32'hc09a7fa6} /* (0, 28, 5) {real, imag} */,
  {32'hc0a95f98, 32'hc1a752a2} /* (0, 28, 4) {real, imag} */,
  {32'h4110bd5a, 32'hc1e84038} /* (0, 28, 3) {real, imag} */,
  {32'hc149a599, 32'hc1aa1d4c} /* (0, 28, 2) {real, imag} */,
  {32'hc1973a83, 32'hbfef3087} /* (0, 28, 1) {real, imag} */,
  {32'hc0a6b74e, 32'h411830ed} /* (0, 28, 0) {real, imag} */,
  {32'hc0c30ce6, 32'h3f1b5dac} /* (0, 27, 31) {real, imag} */,
  {32'hc13d8987, 32'h40b9a83d} /* (0, 27, 30) {real, imag} */,
  {32'hbfb49080, 32'h412daa16} /* (0, 27, 29) {real, imag} */,
  {32'h3f90d89c, 32'hc0c44da3} /* (0, 27, 28) {real, imag} */,
  {32'h4195ab4d, 32'hbfd4ea4e} /* (0, 27, 27) {real, imag} */,
  {32'h3f967c40, 32'hc083a7cb} /* (0, 27, 26) {real, imag} */,
  {32'h3f53d62a, 32'hc1e13382} /* (0, 27, 25) {real, imag} */,
  {32'h4080f849, 32'h3fde62d8} /* (0, 27, 24) {real, imag} */,
  {32'h40116796, 32'hc036217f} /* (0, 27, 23) {real, imag} */,
  {32'h406fe84e, 32'hc0d08268} /* (0, 27, 22) {real, imag} */,
  {32'hc0076290, 32'h3e95b120} /* (0, 27, 21) {real, imag} */,
  {32'hc112f8d8, 32'hc1826869} /* (0, 27, 20) {real, imag} */,
  {32'h3fd36e4c, 32'hc0fc6aba} /* (0, 27, 19) {real, imag} */,
  {32'hc07f3540, 32'hbfa560ac} /* (0, 27, 18) {real, imag} */,
  {32'hc1af3352, 32'h3f0f7910} /* (0, 27, 17) {real, imag} */,
  {32'hc1800734, 32'h40e9f71a} /* (0, 27, 16) {real, imag} */,
  {32'h40664d60, 32'h418a18e7} /* (0, 27, 15) {real, imag} */,
  {32'hc029825f, 32'h413ab656} /* (0, 27, 14) {real, imag} */,
  {32'hc093e746, 32'h41519122} /* (0, 27, 13) {real, imag} */,
  {32'h40ca5895, 32'h41ceb184} /* (0, 27, 12) {real, imag} */,
  {32'h409ac259, 32'h41ae493a} /* (0, 27, 11) {real, imag} */,
  {32'hc0be94f8, 32'hc11d803f} /* (0, 27, 10) {real, imag} */,
  {32'hc18995cd, 32'hc1350258} /* (0, 27, 9) {real, imag} */,
  {32'hc080a683, 32'hc11cfa76} /* (0, 27, 8) {real, imag} */,
  {32'hc128f7dc, 32'hc1c5ad94} /* (0, 27, 7) {real, imag} */,
  {32'hc147a7b1, 32'hc1527da7} /* (0, 27, 6) {real, imag} */,
  {32'hc04cc218, 32'hc1e44d2c} /* (0, 27, 5) {real, imag} */,
  {32'hc07e2748, 32'hc1988b06} /* (0, 27, 4) {real, imag} */,
  {32'hbfd615b0, 32'h41660ae4} /* (0, 27, 3) {real, imag} */,
  {32'hc052fdda, 32'hc090048d} /* (0, 27, 2) {real, imag} */,
  {32'hbf4ee854, 32'hc20f7796} /* (0, 27, 1) {real, imag} */,
  {32'hc12f7c8c, 32'hc199bd75} /* (0, 27, 0) {real, imag} */,
  {32'h40abe9f4, 32'h3fba8674} /* (0, 26, 31) {real, imag} */,
  {32'h407ea19a, 32'h41518016} /* (0, 26, 30) {real, imag} */,
  {32'h4082af13, 32'hc0457906} /* (0, 26, 29) {real, imag} */,
  {32'hc0283f44, 32'hc18a728c} /* (0, 26, 28) {real, imag} */,
  {32'hc0980bd8, 32'hc141fcf2} /* (0, 26, 27) {real, imag} */,
  {32'hc1136e22, 32'hc017e697} /* (0, 26, 26) {real, imag} */,
  {32'hbf329a58, 32'hc18a7178} /* (0, 26, 25) {real, imag} */,
  {32'hc11b68d4, 32'hc065e46e} /* (0, 26, 24) {real, imag} */,
  {32'h4124e1d4, 32'h40528798} /* (0, 26, 23) {real, imag} */,
  {32'h419d220b, 32'hbeafdaf0} /* (0, 26, 22) {real, imag} */,
  {32'h40f435b3, 32'hc06f7b10} /* (0, 26, 21) {real, imag} */,
  {32'hc1681f9d, 32'h403d4ce4} /* (0, 26, 20) {real, imag} */,
  {32'hc09a8cfe, 32'hbec24310} /* (0, 26, 19) {real, imag} */,
  {32'h41164a0c, 32'hc14682bc} /* (0, 26, 18) {real, imag} */,
  {32'h41453ce9, 32'h4191d25a} /* (0, 26, 17) {real, imag} */,
  {32'hc01b4a98, 32'h412c8247} /* (0, 26, 16) {real, imag} */,
  {32'hc130fa0c, 32'hbea32c70} /* (0, 26, 15) {real, imag} */,
  {32'h4030a1d6, 32'hc0707554} /* (0, 26, 14) {real, imag} */,
  {32'h41290fa6, 32'h411b1527} /* (0, 26, 13) {real, imag} */,
  {32'h3ff7addf, 32'h41c62d86} /* (0, 26, 12) {real, imag} */,
  {32'hc0d315f9, 32'h40fbc182} /* (0, 26, 11) {real, imag} */,
  {32'h40d4b054, 32'hc007baf0} /* (0, 26, 10) {real, imag} */,
  {32'h410f03ee, 32'hc0533bf0} /* (0, 26, 9) {real, imag} */,
  {32'h41536154, 32'h4189941e} /* (0, 26, 8) {real, imag} */,
  {32'h417693cc, 32'h412051cf} /* (0, 26, 7) {real, imag} */,
  {32'h410c9730, 32'hc156a1ba} /* (0, 26, 6) {real, imag} */,
  {32'h40ca71e0, 32'hc14432b1} /* (0, 26, 5) {real, imag} */,
  {32'hc06d1fd2, 32'hc12c7bfc} /* (0, 26, 4) {real, imag} */,
  {32'hc0b8ea3d, 32'hc117f2c6} /* (0, 26, 3) {real, imag} */,
  {32'h4054b226, 32'h40c42358} /* (0, 26, 2) {real, imag} */,
  {32'hbfb867a8, 32'h3ff8b6e4} /* (0, 26, 1) {real, imag} */,
  {32'h40aeb411, 32'h4048b6e9} /* (0, 26, 0) {real, imag} */,
  {32'hc10c2e4c, 32'h41b097d6} /* (0, 25, 31) {real, imag} */,
  {32'h3f0a8520, 32'h420a568e} /* (0, 25, 30) {real, imag} */,
  {32'h41654a90, 32'h404b5970} /* (0, 25, 29) {real, imag} */,
  {32'h4154100c, 32'h41392b48} /* (0, 25, 28) {real, imag} */,
  {32'h4131ff2a, 32'h4122ded2} /* (0, 25, 27) {real, imag} */,
  {32'h4114d3e0, 32'hc19b1c79} /* (0, 25, 26) {real, imag} */,
  {32'hc0bd8c72, 32'hc14dcd1a} /* (0, 25, 25) {real, imag} */,
  {32'hc1402f7a, 32'h41aaa542} /* (0, 25, 24) {real, imag} */,
  {32'hc10de720, 32'h410f9252} /* (0, 25, 23) {real, imag} */,
  {32'hc04c3225, 32'hc1197630} /* (0, 25, 22) {real, imag} */,
  {32'h4062d56a, 32'h411ccaa5} /* (0, 25, 21) {real, imag} */,
  {32'h40567ea2, 32'h41514985} /* (0, 25, 20) {real, imag} */,
  {32'hbf8920aa, 32'h40396832} /* (0, 25, 19) {real, imag} */,
  {32'h40cb2c4e, 32'hc0cff380} /* (0, 25, 18) {real, imag} */,
  {32'h3f9a1fe4, 32'h411fbfb9} /* (0, 25, 17) {real, imag} */,
  {32'h406b4590, 32'h420fdb11} /* (0, 25, 16) {real, imag} */,
  {32'h411edfe1, 32'h41815aaa} /* (0, 25, 15) {real, imag} */,
  {32'hbfb3edbc, 32'h40b57a41} /* (0, 25, 14) {real, imag} */,
  {32'hc08ea492, 32'hc0540e07} /* (0, 25, 13) {real, imag} */,
  {32'h402612af, 32'hc1266dfc} /* (0, 25, 12) {real, imag} */,
  {32'h40479b8c, 32'hc0c1dcc2} /* (0, 25, 11) {real, imag} */,
  {32'h3ef107a0, 32'hc119c6ae} /* (0, 25, 10) {real, imag} */,
  {32'hc0bdcb34, 32'h3e358880} /* (0, 25, 9) {real, imag} */,
  {32'h4099f20f, 32'hc110ab20} /* (0, 25, 8) {real, imag} */,
  {32'h40215a08, 32'hc179fab8} /* (0, 25, 7) {real, imag} */,
  {32'h4125822e, 32'h405e759d} /* (0, 25, 6) {real, imag} */,
  {32'hc09cc270, 32'h41ab0452} /* (0, 25, 5) {real, imag} */,
  {32'hc1342a30, 32'h415ed2a4} /* (0, 25, 4) {real, imag} */,
  {32'hc1472384, 32'hbf94ae20} /* (0, 25, 3) {real, imag} */,
  {32'hc04ae7ce, 32'hc19a039c} /* (0, 25, 2) {real, imag} */,
  {32'h3f7c2a24, 32'hc1617d04} /* (0, 25, 1) {real, imag} */,
  {32'hc13a49dc, 32'hc156df14} /* (0, 25, 0) {real, imag} */,
  {32'hc0b95eee, 32'hc0a622ca} /* (0, 24, 31) {real, imag} */,
  {32'hc10de8d4, 32'hc1ae9fbc} /* (0, 24, 30) {real, imag} */,
  {32'hc15578d0, 32'hc09ccfc5} /* (0, 24, 29) {real, imag} */,
  {32'h4027804f, 32'h412f9854} /* (0, 24, 28) {real, imag} */,
  {32'h40f9ef76, 32'h405a88b5} /* (0, 24, 27) {real, imag} */,
  {32'hc0a1e034, 32'hbfb02a84} /* (0, 24, 26) {real, imag} */,
  {32'hc18b4bde, 32'h41563683} /* (0, 24, 25) {real, imag} */,
  {32'hc14b713c, 32'h4092fc1d} /* (0, 24, 24) {real, imag} */,
  {32'hbcb5de00, 32'hbf0ff0e7} /* (0, 24, 23) {real, imag} */,
  {32'hbd63b600, 32'hc103fbb0} /* (0, 24, 22) {real, imag} */,
  {32'h416f8a40, 32'hc174680a} /* (0, 24, 21) {real, imag} */,
  {32'hc032754c, 32'h40a8584c} /* (0, 24, 20) {real, imag} */,
  {32'h409967c1, 32'h41392dda} /* (0, 24, 19) {real, imag} */,
  {32'h42112b36, 32'hbf6bdef0} /* (0, 24, 18) {real, imag} */,
  {32'h419ab9ca, 32'hc1026c22} /* (0, 24, 17) {real, imag} */,
  {32'hc021a5ac, 32'hc10e7d87} /* (0, 24, 16) {real, imag} */,
  {32'hc1363a40, 32'hbfef48ae} /* (0, 24, 15) {real, imag} */,
  {32'hc136991a, 32'hc1081baa} /* (0, 24, 14) {real, imag} */,
  {32'hc17fa5d8, 32'hc0b77d3e} /* (0, 24, 13) {real, imag} */,
  {32'hbff15816, 32'h417fe27a} /* (0, 24, 12) {real, imag} */,
  {32'hc0b59fb4, 32'h412c03b4} /* (0, 24, 11) {real, imag} */,
  {32'h40bdf59d, 32'h3fe479f8} /* (0, 24, 10) {real, imag} */,
  {32'h41a9ddfe, 32'hc0e8634c} /* (0, 24, 9) {real, imag} */,
  {32'h3f037910, 32'hc048edd2} /* (0, 24, 8) {real, imag} */,
  {32'hc0df2e74, 32'hc15abac2} /* (0, 24, 7) {real, imag} */,
  {32'h41387acf, 32'hc0c36277} /* (0, 24, 6) {real, imag} */,
  {32'hc101538a, 32'h41a3e1b6} /* (0, 24, 5) {real, imag} */,
  {32'hc16bc76f, 32'hbf477b40} /* (0, 24, 4) {real, imag} */,
  {32'h402cdfb8, 32'hc100f028} /* (0, 24, 3) {real, imag} */,
  {32'hc08d2f82, 32'h40b7f654} /* (0, 24, 2) {real, imag} */,
  {32'hc17fc9bd, 32'h4174d2d7} /* (0, 24, 1) {real, imag} */,
  {32'hc0faaac0, 32'h3f96e382} /* (0, 24, 0) {real, imag} */,
  {32'hc0fc7024, 32'hc0304360} /* (0, 23, 31) {real, imag} */,
  {32'hc10f8c4c, 32'h3db35b00} /* (0, 23, 30) {real, imag} */,
  {32'hc1aed052, 32'hc11b4b11} /* (0, 23, 29) {real, imag} */,
  {32'hc1a4bbd6, 32'hc0ecbbbc} /* (0, 23, 28) {real, imag} */,
  {32'hc1b5951f, 32'hc04e9fd0} /* (0, 23, 27) {real, imag} */,
  {32'hc1d9f7c4, 32'hc1484c96} /* (0, 23, 26) {real, imag} */,
  {32'hc1bd0a0a, 32'hc0ab0064} /* (0, 23, 25) {real, imag} */,
  {32'hc17b1402, 32'h404bc2a4} /* (0, 23, 24) {real, imag} */,
  {32'hc1950569, 32'h41517e02} /* (0, 23, 23) {real, imag} */,
  {32'hc01c0975, 32'h41355310} /* (0, 23, 22) {real, imag} */,
  {32'hc0cf54df, 32'h41825bab} /* (0, 23, 21) {real, imag} */,
  {32'h3f9f7110, 32'h413315d5} /* (0, 23, 20) {real, imag} */,
  {32'h40a7f5de, 32'h40d2e4b5} /* (0, 23, 19) {real, imag} */,
  {32'h414ae82d, 32'hc0b07548} /* (0, 23, 18) {real, imag} */,
  {32'h410166c8, 32'h410b7af3} /* (0, 23, 17) {real, imag} */,
  {32'h40ebb65e, 32'h41832ed2} /* (0, 23, 16) {real, imag} */,
  {32'hc10e9d21, 32'hc084d1af} /* (0, 23, 15) {real, imag} */,
  {32'h4052e896, 32'hc0f76aaf} /* (0, 23, 14) {real, imag} */,
  {32'h40fc2672, 32'h3fb1ef8a} /* (0, 23, 13) {real, imag} */,
  {32'h406402e7, 32'hc042a975} /* (0, 23, 12) {real, imag} */,
  {32'h41396145, 32'hc0f3d21c} /* (0, 23, 11) {real, imag} */,
  {32'h40b7f7c4, 32'hc078b9f0} /* (0, 23, 10) {real, imag} */,
  {32'hbe95f8e8, 32'h3facc8a8} /* (0, 23, 9) {real, imag} */,
  {32'h40f95a59, 32'hc0b2bafc} /* (0, 23, 8) {real, imag} */,
  {32'h406b0b54, 32'hc0fb3977} /* (0, 23, 7) {real, imag} */,
  {32'h4093b4bf, 32'h3fa0b8f6} /* (0, 23, 6) {real, imag} */,
  {32'h415d9c92, 32'hc0ac505a} /* (0, 23, 5) {real, imag} */,
  {32'h416357a0, 32'hc07e1f70} /* (0, 23, 4) {real, imag} */,
  {32'h40f67a20, 32'h418fb97d} /* (0, 23, 3) {real, imag} */,
  {32'h40b58da3, 32'h413a4a12} /* (0, 23, 2) {real, imag} */,
  {32'hc08a7a9e, 32'h40c85d1b} /* (0, 23, 1) {real, imag} */,
  {32'hc133de30, 32'hc0fc8377} /* (0, 23, 0) {real, imag} */,
  {32'h4024af10, 32'h414080f2} /* (0, 22, 31) {real, imag} */,
  {32'hc050955e, 32'h41406070} /* (0, 22, 30) {real, imag} */,
  {32'hbfc4089c, 32'hc02af6f4} /* (0, 22, 29) {real, imag} */,
  {32'h40beb112, 32'hc09a21ba} /* (0, 22, 28) {real, imag} */,
  {32'h3da8b300, 32'h408b3de3} /* (0, 22, 27) {real, imag} */,
  {32'hc039fa1c, 32'hc035ca39} /* (0, 22, 26) {real, imag} */,
  {32'hc067865a, 32'hc11965a2} /* (0, 22, 25) {real, imag} */,
  {32'hc19c89cc, 32'hc12fed4c} /* (0, 22, 24) {real, imag} */,
  {32'hc0b89ea8, 32'hc050d898} /* (0, 22, 23) {real, imag} */,
  {32'hc08070b8, 32'h40d1ab1d} /* (0, 22, 22) {real, imag} */,
  {32'hc1297acc, 32'hc04984bc} /* (0, 22, 21) {real, imag} */,
  {32'hc09bbc86, 32'hbec916a4} /* (0, 22, 20) {real, imag} */,
  {32'hbee9b528, 32'hc1577e06} /* (0, 22, 19) {real, imag} */,
  {32'h40bf6372, 32'hc0017cd8} /* (0, 22, 18) {real, imag} */,
  {32'h40a013c6, 32'h4111cec3} /* (0, 22, 17) {real, imag} */,
  {32'hc0f869c0, 32'hc0f8f71e} /* (0, 22, 16) {real, imag} */,
  {32'h412ec744, 32'hc1029aac} /* (0, 22, 15) {real, imag} */,
  {32'h411b5de8, 32'h3fa477f1} /* (0, 22, 14) {real, imag} */,
  {32'hc0699ad6, 32'hc0cb20d2} /* (0, 22, 13) {real, imag} */,
  {32'h3fbd727d, 32'hc1067b3d} /* (0, 22, 12) {real, imag} */,
  {32'hbfd943dc, 32'hc0d0827e} /* (0, 22, 11) {real, imag} */,
  {32'hc0b68bb6, 32'hc141fab8} /* (0, 22, 10) {real, imag} */,
  {32'hc0998dbf, 32'h41194f30} /* (0, 22, 9) {real, imag} */,
  {32'h407d0c98, 32'h41b682f2} /* (0, 22, 8) {real, imag} */,
  {32'h408aa9b8, 32'h418b92b2} /* (0, 22, 7) {real, imag} */,
  {32'h406b95ca, 32'h40db24b9} /* (0, 22, 6) {real, imag} */,
  {32'h41278e96, 32'hc0a9c4fe} /* (0, 22, 5) {real, imag} */,
  {32'h4029d17a, 32'hc12d3a00} /* (0, 22, 4) {real, imag} */,
  {32'h40538a66, 32'hc085805b} /* (0, 22, 3) {real, imag} */,
  {32'hc089cb0b, 32'hc1041476} /* (0, 22, 2) {real, imag} */,
  {32'hc120b477, 32'hbfb857dc} /* (0, 22, 1) {real, imag} */,
  {32'hc02a59b6, 32'h411ec35e} /* (0, 22, 0) {real, imag} */,
  {32'h40513778, 32'hc096b00e} /* (0, 21, 31) {real, imag} */,
  {32'h404969d4, 32'hc0cea429} /* (0, 21, 30) {real, imag} */,
  {32'hc05d7c94, 32'h40227eee} /* (0, 21, 29) {real, imag} */,
  {32'hbd663380, 32'h40bc7bf7} /* (0, 21, 28) {real, imag} */,
  {32'h40eab7db, 32'h402cd4b9} /* (0, 21, 27) {real, imag} */,
  {32'h4086b1fe, 32'hc1053db4} /* (0, 21, 26) {real, imag} */,
  {32'h4060947e, 32'h407945f0} /* (0, 21, 25) {real, imag} */,
  {32'h408ca9bb, 32'hc06d10f4} /* (0, 21, 24) {real, imag} */,
  {32'hc0dd9343, 32'hc013a8b9} /* (0, 21, 23) {real, imag} */,
  {32'hc10d06ee, 32'h40472849} /* (0, 21, 22) {real, imag} */,
  {32'h40f3a6ae, 32'h40a604b8} /* (0, 21, 21) {real, imag} */,
  {32'hbfac6694, 32'h4084589b} /* (0, 21, 20) {real, imag} */,
  {32'hc09704c0, 32'h3f13e414} /* (0, 21, 19) {real, imag} */,
  {32'hc07b6a62, 32'h408dcd63} /* (0, 21, 18) {real, imag} */,
  {32'hbfe6f1c8, 32'h3f3c44ec} /* (0, 21, 17) {real, imag} */,
  {32'hc0bffa46, 32'hbbf68e00} /* (0, 21, 16) {real, imag} */,
  {32'hc006a7ac, 32'hbfe8c0f4} /* (0, 21, 15) {real, imag} */,
  {32'h401edba9, 32'h40375006} /* (0, 21, 14) {real, imag} */,
  {32'hbdc394a0, 32'h3f8e3774} /* (0, 21, 13) {real, imag} */,
  {32'h410ba8b8, 32'hc0aaa3b4} /* (0, 21, 12) {real, imag} */,
  {32'h40e4e9e5, 32'h402774a8} /* (0, 21, 11) {real, imag} */,
  {32'h3ff33a62, 32'h4040c867} /* (0, 21, 10) {real, imag} */,
  {32'h40ace95c, 32'h3f93e08c} /* (0, 21, 9) {real, imag} */,
  {32'hbd8809c0, 32'h40b76019} /* (0, 21, 8) {real, imag} */,
  {32'hc0957ec0, 32'h4135ca48} /* (0, 21, 7) {real, imag} */,
  {32'hc13074f1, 32'h3fb5d438} /* (0, 21, 6) {real, imag} */,
  {32'hc0fbdc44, 32'h40152aa0} /* (0, 21, 5) {real, imag} */,
  {32'h40dd5510, 32'h3feec388} /* (0, 21, 4) {real, imag} */,
  {32'h41263c58, 32'h40b077b7} /* (0, 21, 3) {real, imag} */,
  {32'hc010c454, 32'h408da35d} /* (0, 21, 2) {real, imag} */,
  {32'hc03e7ad1, 32'h41205fee} /* (0, 21, 1) {real, imag} */,
  {32'hc0543f08, 32'h406b44a6} /* (0, 21, 0) {real, imag} */,
  {32'h3fb8e631, 32'h40b1855e} /* (0, 20, 31) {real, imag} */,
  {32'h40c4be5e, 32'hbf2d4678} /* (0, 20, 30) {real, imag} */,
  {32'h410ea9fd, 32'hc105a03a} /* (0, 20, 29) {real, imag} */,
  {32'h4117145c, 32'hc09278ca} /* (0, 20, 28) {real, imag} */,
  {32'h40ed5f86, 32'hbe026a28} /* (0, 20, 27) {real, imag} */,
  {32'h40f6e67c, 32'h40372cc5} /* (0, 20, 26) {real, imag} */,
  {32'h410282aa, 32'h4120fc30} /* (0, 20, 25) {real, imag} */,
  {32'h40de6ed6, 32'h40efa9a0} /* (0, 20, 24) {real, imag} */,
  {32'h3f859e8c, 32'h415926c2} /* (0, 20, 23) {real, imag} */,
  {32'h402f9eb0, 32'h411d7454} /* (0, 20, 22) {real, imag} */,
  {32'hbe3d1740, 32'h403adf86} /* (0, 20, 21) {real, imag} */,
  {32'hc0b930c4, 32'h41077fd2} /* (0, 20, 20) {real, imag} */,
  {32'h40bd7eb8, 32'h402131f0} /* (0, 20, 19) {real, imag} */,
  {32'h4058ac30, 32'h3fbf6b40} /* (0, 20, 18) {real, imag} */,
  {32'hbfb644ae, 32'hc0d9a5f6} /* (0, 20, 17) {real, imag} */,
  {32'hc037f726, 32'hc00c8f4c} /* (0, 20, 16) {real, imag} */,
  {32'hbec8ca10, 32'h40f1f0dd} /* (0, 20, 15) {real, imag} */,
  {32'h3d9e9a9b, 32'h4137b988} /* (0, 20, 14) {real, imag} */,
  {32'h40ec7810, 32'h40541fbc} /* (0, 20, 13) {real, imag} */,
  {32'hc0094878, 32'hbfc3b924} /* (0, 20, 12) {real, imag} */,
  {32'hc0834848, 32'h4103fe34} /* (0, 20, 11) {real, imag} */,
  {32'h3fce50a0, 32'h41040ecf} /* (0, 20, 10) {real, imag} */,
  {32'h4035aaad, 32'hc02dc31f} /* (0, 20, 9) {real, imag} */,
  {32'h40942eaf, 32'h3f8340d4} /* (0, 20, 8) {real, imag} */,
  {32'h4071ebba, 32'h3ffc0208} /* (0, 20, 7) {real, imag} */,
  {32'h40ca6826, 32'hc053c1ac} /* (0, 20, 6) {real, imag} */,
  {32'h40be4777, 32'hc000cf04} /* (0, 20, 5) {real, imag} */,
  {32'h40a451aa, 32'hc015d18c} /* (0, 20, 4) {real, imag} */,
  {32'h4077f27e, 32'hc08c11d2} /* (0, 20, 3) {real, imag} */,
  {32'h3f05a370, 32'hc04559d0} /* (0, 20, 2) {real, imag} */,
  {32'h40a10309, 32'h4090fa85} /* (0, 20, 1) {real, imag} */,
  {32'h401a04ed, 32'h403afba9} /* (0, 20, 0) {real, imag} */,
  {32'h3fc6c3f4, 32'hbf7f3c48} /* (0, 19, 31) {real, imag} */,
  {32'h3bcd0000, 32'h40b175b6} /* (0, 19, 30) {real, imag} */,
  {32'hbf066c00, 32'h405e4d6a} /* (0, 19, 29) {real, imag} */,
  {32'h4060d756, 32'h3f9033b8} /* (0, 19, 28) {real, imag} */,
  {32'h3fe9cf5a, 32'h4119c9c6} /* (0, 19, 27) {real, imag} */,
  {32'hbfb91c2c, 32'h412df5a0} /* (0, 19, 26) {real, imag} */,
  {32'h3ee027e0, 32'h40d20553} /* (0, 19, 25) {real, imag} */,
  {32'h401c0180, 32'h3fdc6eb0} /* (0, 19, 24) {real, imag} */,
  {32'h40c47402, 32'hc0c36044} /* (0, 19, 23) {real, imag} */,
  {32'h3f7dbc8a, 32'hc150dea8} /* (0, 19, 22) {real, imag} */,
  {32'h3fc0a5c0, 32'hbf9f8340} /* (0, 19, 21) {real, imag} */,
  {32'h414e4753, 32'h4052806f} /* (0, 19, 20) {real, imag} */,
  {32'h41365c68, 32'h3fe1fb30} /* (0, 19, 19) {real, imag} */,
  {32'hbe05da30, 32'h3d6b4060} /* (0, 19, 18) {real, imag} */,
  {32'hc088c2f0, 32'hc1012e32} /* (0, 19, 17) {real, imag} */,
  {32'hbfaba6a8, 32'h406d12b0} /* (0, 19, 16) {real, imag} */,
  {32'hc04efaa8, 32'h41223e66} /* (0, 19, 15) {real, imag} */,
  {32'hc1378846, 32'hbec0ed24} /* (0, 19, 14) {real, imag} */,
  {32'hc0398b18, 32'hc05ddfe7} /* (0, 19, 13) {real, imag} */,
  {32'hc03bf6e8, 32'hbef065f0} /* (0, 19, 12) {real, imag} */,
  {32'hc0a4075e, 32'h40ab780a} /* (0, 19, 11) {real, imag} */,
  {32'hc028f2cc, 32'h3ff70786} /* (0, 19, 10) {real, imag} */,
  {32'hc118b710, 32'hbfa10008} /* (0, 19, 9) {real, imag} */,
  {32'hc11bbdc8, 32'hc008ccd8} /* (0, 19, 8) {real, imag} */,
  {32'hc0f76eae, 32'hc085430a} /* (0, 19, 7) {real, imag} */,
  {32'hc108fd23, 32'hc00d47b8} /* (0, 19, 6) {real, imag} */,
  {32'hbe5b3760, 32'h3f2f62a8} /* (0, 19, 5) {real, imag} */,
  {32'hbe5d3980, 32'hbf8c56ba} /* (0, 19, 4) {real, imag} */,
  {32'hc0544f8d, 32'hc12f09a6} /* (0, 19, 3) {real, imag} */,
  {32'hc0d52176, 32'hc084b6ae} /* (0, 19, 2) {real, imag} */,
  {32'hc0c1bb37, 32'hbf1b6320} /* (0, 19, 1) {real, imag} */,
  {32'hc07fb75a, 32'h3eef52a0} /* (0, 19, 0) {real, imag} */,
  {32'hbf90a91f, 32'hc0890311} /* (0, 18, 31) {real, imag} */,
  {32'hbffa8088, 32'hc106b440} /* (0, 18, 30) {real, imag} */,
  {32'hc09f7728, 32'hc08b2828} /* (0, 18, 29) {real, imag} */,
  {32'hc0477428, 32'hbfe98328} /* (0, 18, 28) {real, imag} */,
  {32'hc10a3f57, 32'hc0114191} /* (0, 18, 27) {real, imag} */,
  {32'hc109aacc, 32'hc0de3562} /* (0, 18, 26) {real, imag} */,
  {32'hbf92efb0, 32'hc09b92a0} /* (0, 18, 25) {real, imag} */,
  {32'h3f93a274, 32'h4036bcde} /* (0, 18, 24) {real, imag} */,
  {32'h3f283ce2, 32'hc062066c} /* (0, 18, 23) {real, imag} */,
  {32'h3f4d8c50, 32'hc0fdd4fa} /* (0, 18, 22) {real, imag} */,
  {32'h40c8513d, 32'hc10cfc90} /* (0, 18, 21) {real, imag} */,
  {32'h40c34d42, 32'hc0081ef5} /* (0, 18, 20) {real, imag} */,
  {32'hbff64848, 32'hbe9d3850} /* (0, 18, 19) {real, imag} */,
  {32'hc078e33d, 32'hc08c9a29} /* (0, 18, 18) {real, imag} */,
  {32'h3ee34110, 32'hc069f7e6} /* (0, 18, 17) {real, imag} */,
  {32'h4028a330, 32'hc015ac38} /* (0, 18, 16) {real, imag} */,
  {32'hbe0b6360, 32'hbf614e28} /* (0, 18, 15) {real, imag} */,
  {32'hbff7a69f, 32'hc005ad68} /* (0, 18, 14) {real, imag} */,
  {32'h40312b09, 32'hc041b428} /* (0, 18, 13) {real, imag} */,
  {32'h40b9a0d8, 32'h3f287e38} /* (0, 18, 12) {real, imag} */,
  {32'h412af94f, 32'h3fe6d2e0} /* (0, 18, 11) {real, imag} */,
  {32'h40bee582, 32'h40e1d035} /* (0, 18, 10) {real, imag} */,
  {32'h40c62524, 32'h3fc2ace8} /* (0, 18, 9) {real, imag} */,
  {32'h40cdf5be, 32'h3f5fa3d0} /* (0, 18, 8) {real, imag} */,
  {32'h3fe776d0, 32'h3f7bb412} /* (0, 18, 7) {real, imag} */,
  {32'hbea82fe0, 32'hbfbbdb95} /* (0, 18, 6) {real, imag} */,
  {32'hc0095c9e, 32'hc0d45b34} /* (0, 18, 5) {real, imag} */,
  {32'hc03264c2, 32'hc0171aee} /* (0, 18, 4) {real, imag} */,
  {32'h4030896e, 32'h3fc659b6} /* (0, 18, 3) {real, imag} */,
  {32'hc08dd101, 32'h3fa969a8} /* (0, 18, 2) {real, imag} */,
  {32'hc0dfa5ec, 32'h4015d058} /* (0, 18, 1) {real, imag} */,
  {32'hbf96359c, 32'h3fd61fdd} /* (0, 18, 0) {real, imag} */,
  {32'hc017d501, 32'h3f2cd616} /* (0, 17, 31) {real, imag} */,
  {32'h3f58abc4, 32'h407ea980} /* (0, 17, 30) {real, imag} */,
  {32'hc073056e, 32'h4118faac} /* (0, 17, 29) {real, imag} */,
  {32'hbf9a479c, 32'h40c0c39c} /* (0, 17, 28) {real, imag} */,
  {32'h40586948, 32'h406da72c} /* (0, 17, 27) {real, imag} */,
  {32'hbd80c0e0, 32'h40ec3e96} /* (0, 17, 26) {real, imag} */,
  {32'hbfd2eb92, 32'h40dead26} /* (0, 17, 25) {real, imag} */,
  {32'h403a021a, 32'h3ef2feb8} /* (0, 17, 24) {real, imag} */,
  {32'h4057e65e, 32'hbfaa91b0} /* (0, 17, 23) {real, imag} */,
  {32'h40857cd3, 32'hc03743b8} /* (0, 17, 22) {real, imag} */,
  {32'h4080db8c, 32'hc040e50f} /* (0, 17, 21) {real, imag} */,
  {32'hbf63aea0, 32'hc09d1b1a} /* (0, 17, 20) {real, imag} */,
  {32'hc02fe21c, 32'hc017c64c} /* (0, 17, 19) {real, imag} */,
  {32'h4016a84a, 32'h40cc26b6} /* (0, 17, 18) {real, imag} */,
  {32'h4016c31f, 32'h3e32cda0} /* (0, 17, 17) {real, imag} */,
  {32'h409fbcad, 32'hc0819df2} /* (0, 17, 16) {real, imag} */,
  {32'h40ac1a2c, 32'hc09fb304} /* (0, 17, 15) {real, imag} */,
  {32'h3fcff7c4, 32'hbecf1c68} /* (0, 17, 14) {real, imag} */,
  {32'hc0819246, 32'hc0a08a13} /* (0, 17, 13) {real, imag} */,
  {32'hbfd7015e, 32'hc04c7007} /* (0, 17, 12) {real, imag} */,
  {32'h3f45be58, 32'hbef13890} /* (0, 17, 11) {real, imag} */,
  {32'hc04067d6, 32'h3e900c30} /* (0, 17, 10) {real, imag} */,
  {32'h3e60edc0, 32'h3ea3ed60} /* (0, 17, 9) {real, imag} */,
  {32'hbfac1e90, 32'h408c5188} /* (0, 17, 8) {real, imag} */,
  {32'hc0d1a1ce, 32'hbd220e00} /* (0, 17, 7) {real, imag} */,
  {32'hc08b4448, 32'hc0ffbb28} /* (0, 17, 6) {real, imag} */,
  {32'h400cb8d4, 32'hc0c6eae6} /* (0, 17, 5) {real, imag} */,
  {32'h406ed689, 32'hbfe22450} /* (0, 17, 4) {real, imag} */,
  {32'h405b7754, 32'h3fb5f914} /* (0, 17, 3) {real, imag} */,
  {32'hbf0d7c28, 32'h4064f1d6} /* (0, 17, 2) {real, imag} */,
  {32'hbf0d1ce4, 32'hbfc36568} /* (0, 17, 1) {real, imag} */,
  {32'hbfd160e8, 32'hbf67e500} /* (0, 17, 0) {real, imag} */,
  {32'hbdf5ca00, 32'h00000000} /* (0, 16, 31) {real, imag} */,
  {32'h40717c86, 32'h00000000} /* (0, 16, 30) {real, imag} */,
  {32'hbef16a80, 32'h00000000} /* (0, 16, 29) {real, imag} */,
  {32'hc0f1ad6d, 32'h00000000} /* (0, 16, 28) {real, imag} */,
  {32'hbebb0fc0, 32'h00000000} /* (0, 16, 27) {real, imag} */,
  {32'h403e45f0, 32'h00000000} /* (0, 16, 26) {real, imag} */,
  {32'h40cce096, 32'h00000000} /* (0, 16, 25) {real, imag} */,
  {32'h40769ca2, 32'h00000000} /* (0, 16, 24) {real, imag} */,
  {32'h40b3f705, 32'h00000000} /* (0, 16, 23) {real, imag} */,
  {32'h3fc68f00, 32'h00000000} /* (0, 16, 22) {real, imag} */,
  {32'hc05e8f28, 32'h00000000} /* (0, 16, 21) {real, imag} */,
  {32'hc0a357e8, 32'h00000000} /* (0, 16, 20) {real, imag} */,
  {32'hc0b482b1, 32'h00000000} /* (0, 16, 19) {real, imag} */,
  {32'hbf406020, 32'h00000000} /* (0, 16, 18) {real, imag} */,
  {32'h4057dab4, 32'h00000000} /* (0, 16, 17) {real, imag} */,
  {32'h40cc325b, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hc0416cbe, 32'h00000000} /* (0, 16, 15) {real, imag} */,
  {32'hc04cbaf0, 32'h00000000} /* (0, 16, 14) {real, imag} */,
  {32'h3f7c1e04, 32'h00000000} /* (0, 16, 13) {real, imag} */,
  {32'h3f414aec, 32'h00000000} /* (0, 16, 12) {real, imag} */,
  {32'h3fa05248, 32'h00000000} /* (0, 16, 11) {real, imag} */,
  {32'h4077dcb6, 32'h00000000} /* (0, 16, 10) {real, imag} */,
  {32'h40ac10dc, 32'h00000000} /* (0, 16, 9) {real, imag} */,
  {32'h4016fbb4, 32'h00000000} /* (0, 16, 8) {real, imag} */,
  {32'h3faea860, 32'h00000000} /* (0, 16, 7) {real, imag} */,
  {32'h411ec02f, 32'h00000000} /* (0, 16, 6) {real, imag} */,
  {32'h414fa0e4, 32'h00000000} /* (0, 16, 5) {real, imag} */,
  {32'h40cc3d92, 32'h00000000} /* (0, 16, 4) {real, imag} */,
  {32'h40823220, 32'h00000000} /* (0, 16, 3) {real, imag} */,
  {32'h40f1e7f2, 32'h00000000} /* (0, 16, 2) {real, imag} */,
  {32'h3c839c00, 32'h00000000} /* (0, 16, 1) {real, imag} */,
  {32'hc0215d55, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'hc017d501, 32'hbf2cd616} /* (0, 15, 31) {real, imag} */,
  {32'h3f58abc4, 32'hc07ea980} /* (0, 15, 30) {real, imag} */,
  {32'hc073056e, 32'hc118faac} /* (0, 15, 29) {real, imag} */,
  {32'hbf9a479c, 32'hc0c0c39c} /* (0, 15, 28) {real, imag} */,
  {32'h40586948, 32'hc06da72c} /* (0, 15, 27) {real, imag} */,
  {32'hbd80c0e0, 32'hc0ec3e96} /* (0, 15, 26) {real, imag} */,
  {32'hbfd2eb92, 32'hc0dead26} /* (0, 15, 25) {real, imag} */,
  {32'h403a021a, 32'hbef2feb8} /* (0, 15, 24) {real, imag} */,
  {32'h4057e65e, 32'h3faa91b0} /* (0, 15, 23) {real, imag} */,
  {32'h40857cd3, 32'h403743b8} /* (0, 15, 22) {real, imag} */,
  {32'h4080db8c, 32'h4040e50f} /* (0, 15, 21) {real, imag} */,
  {32'hbf63aea0, 32'h409d1b1a} /* (0, 15, 20) {real, imag} */,
  {32'hc02fe21c, 32'h4017c64c} /* (0, 15, 19) {real, imag} */,
  {32'h4016a84a, 32'hc0cc26b6} /* (0, 15, 18) {real, imag} */,
  {32'h4016c31f, 32'hbe32cda0} /* (0, 15, 17) {real, imag} */,
  {32'h409fbcad, 32'h40819df2} /* (0, 15, 16) {real, imag} */,
  {32'h40ac1a2c, 32'h409fb304} /* (0, 15, 15) {real, imag} */,
  {32'h3fcff7c4, 32'h3ecf1c68} /* (0, 15, 14) {real, imag} */,
  {32'hc0819246, 32'h40a08a13} /* (0, 15, 13) {real, imag} */,
  {32'hbfd7015e, 32'h404c7007} /* (0, 15, 12) {real, imag} */,
  {32'h3f45be58, 32'h3ef13890} /* (0, 15, 11) {real, imag} */,
  {32'hc04067d6, 32'hbe900c30} /* (0, 15, 10) {real, imag} */,
  {32'h3e60edc0, 32'hbea3ed60} /* (0, 15, 9) {real, imag} */,
  {32'hbfac1e90, 32'hc08c5188} /* (0, 15, 8) {real, imag} */,
  {32'hc0d1a1ce, 32'h3d220e00} /* (0, 15, 7) {real, imag} */,
  {32'hc08b4448, 32'h40ffbb28} /* (0, 15, 6) {real, imag} */,
  {32'h400cb8d4, 32'h40c6eae6} /* (0, 15, 5) {real, imag} */,
  {32'h406ed689, 32'h3fe22450} /* (0, 15, 4) {real, imag} */,
  {32'h405b7754, 32'hbfb5f914} /* (0, 15, 3) {real, imag} */,
  {32'hbf0d7c28, 32'hc064f1d6} /* (0, 15, 2) {real, imag} */,
  {32'hbf0d1ce4, 32'h3fc36568} /* (0, 15, 1) {real, imag} */,
  {32'hbfd160e8, 32'h3f67e500} /* (0, 15, 0) {real, imag} */,
  {32'hbf90a91f, 32'h40890311} /* (0, 14, 31) {real, imag} */,
  {32'hbffa8088, 32'h4106b440} /* (0, 14, 30) {real, imag} */,
  {32'hc09f7728, 32'h408b2828} /* (0, 14, 29) {real, imag} */,
  {32'hc0477428, 32'h3fe98328} /* (0, 14, 28) {real, imag} */,
  {32'hc10a3f57, 32'h40114191} /* (0, 14, 27) {real, imag} */,
  {32'hc109aacc, 32'h40de3562} /* (0, 14, 26) {real, imag} */,
  {32'hbf92efb0, 32'h409b92a0} /* (0, 14, 25) {real, imag} */,
  {32'h3f93a274, 32'hc036bcde} /* (0, 14, 24) {real, imag} */,
  {32'h3f283ce2, 32'h4062066c} /* (0, 14, 23) {real, imag} */,
  {32'h3f4d8c50, 32'h40fdd4fa} /* (0, 14, 22) {real, imag} */,
  {32'h40c8513d, 32'h410cfc90} /* (0, 14, 21) {real, imag} */,
  {32'h40c34d42, 32'h40081ef5} /* (0, 14, 20) {real, imag} */,
  {32'hbff64848, 32'h3e9d3850} /* (0, 14, 19) {real, imag} */,
  {32'hc078e33d, 32'h408c9a29} /* (0, 14, 18) {real, imag} */,
  {32'h3ee34110, 32'h4069f7e6} /* (0, 14, 17) {real, imag} */,
  {32'h4028a330, 32'h4015ac38} /* (0, 14, 16) {real, imag} */,
  {32'hbe0b6360, 32'h3f614e28} /* (0, 14, 15) {real, imag} */,
  {32'hbff7a69f, 32'h4005ad68} /* (0, 14, 14) {real, imag} */,
  {32'h40312b09, 32'h4041b428} /* (0, 14, 13) {real, imag} */,
  {32'h40b9a0d8, 32'hbf287e38} /* (0, 14, 12) {real, imag} */,
  {32'h412af94f, 32'hbfe6d2e0} /* (0, 14, 11) {real, imag} */,
  {32'h40bee582, 32'hc0e1d035} /* (0, 14, 10) {real, imag} */,
  {32'h40c62524, 32'hbfc2ace8} /* (0, 14, 9) {real, imag} */,
  {32'h40cdf5be, 32'hbf5fa3d0} /* (0, 14, 8) {real, imag} */,
  {32'h3fe776d0, 32'hbf7bb412} /* (0, 14, 7) {real, imag} */,
  {32'hbea82fe0, 32'h3fbbdb95} /* (0, 14, 6) {real, imag} */,
  {32'hc0095c9e, 32'h40d45b34} /* (0, 14, 5) {real, imag} */,
  {32'hc03264c2, 32'h40171aee} /* (0, 14, 4) {real, imag} */,
  {32'h4030896e, 32'hbfc659b6} /* (0, 14, 3) {real, imag} */,
  {32'hc08dd101, 32'hbfa969a8} /* (0, 14, 2) {real, imag} */,
  {32'hc0dfa5ec, 32'hc015d058} /* (0, 14, 1) {real, imag} */,
  {32'hbf96359c, 32'hbfd61fdd} /* (0, 14, 0) {real, imag} */,
  {32'h3fc6c3f4, 32'h3f7f3c48} /* (0, 13, 31) {real, imag} */,
  {32'h3bcd0000, 32'hc0b175b6} /* (0, 13, 30) {real, imag} */,
  {32'hbf066c00, 32'hc05e4d6a} /* (0, 13, 29) {real, imag} */,
  {32'h4060d756, 32'hbf9033b8} /* (0, 13, 28) {real, imag} */,
  {32'h3fe9cf5a, 32'hc119c9c6} /* (0, 13, 27) {real, imag} */,
  {32'hbfb91c2c, 32'hc12df5a0} /* (0, 13, 26) {real, imag} */,
  {32'h3ee027e0, 32'hc0d20553} /* (0, 13, 25) {real, imag} */,
  {32'h401c0180, 32'hbfdc6eb0} /* (0, 13, 24) {real, imag} */,
  {32'h40c47402, 32'h40c36044} /* (0, 13, 23) {real, imag} */,
  {32'h3f7dbc8a, 32'h4150dea8} /* (0, 13, 22) {real, imag} */,
  {32'h3fc0a5c0, 32'h3f9f8340} /* (0, 13, 21) {real, imag} */,
  {32'h414e4753, 32'hc052806f} /* (0, 13, 20) {real, imag} */,
  {32'h41365c68, 32'hbfe1fb30} /* (0, 13, 19) {real, imag} */,
  {32'hbe05da30, 32'hbd6b4060} /* (0, 13, 18) {real, imag} */,
  {32'hc088c2f0, 32'h41012e32} /* (0, 13, 17) {real, imag} */,
  {32'hbfaba6a8, 32'hc06d12b0} /* (0, 13, 16) {real, imag} */,
  {32'hc04efaa8, 32'hc1223e66} /* (0, 13, 15) {real, imag} */,
  {32'hc1378846, 32'h3ec0ed24} /* (0, 13, 14) {real, imag} */,
  {32'hc0398b18, 32'h405ddfe7} /* (0, 13, 13) {real, imag} */,
  {32'hc03bf6e8, 32'h3ef065f0} /* (0, 13, 12) {real, imag} */,
  {32'hc0a4075e, 32'hc0ab780a} /* (0, 13, 11) {real, imag} */,
  {32'hc028f2cc, 32'hbff70786} /* (0, 13, 10) {real, imag} */,
  {32'hc118b710, 32'h3fa10008} /* (0, 13, 9) {real, imag} */,
  {32'hc11bbdc8, 32'h4008ccd8} /* (0, 13, 8) {real, imag} */,
  {32'hc0f76eae, 32'h4085430a} /* (0, 13, 7) {real, imag} */,
  {32'hc108fd23, 32'h400d47b8} /* (0, 13, 6) {real, imag} */,
  {32'hbe5b3760, 32'hbf2f62a8} /* (0, 13, 5) {real, imag} */,
  {32'hbe5d3980, 32'h3f8c56ba} /* (0, 13, 4) {real, imag} */,
  {32'hc0544f8d, 32'h412f09a6} /* (0, 13, 3) {real, imag} */,
  {32'hc0d52176, 32'h4084b6ae} /* (0, 13, 2) {real, imag} */,
  {32'hc0c1bb37, 32'h3f1b6320} /* (0, 13, 1) {real, imag} */,
  {32'hc07fb75a, 32'hbeef52a0} /* (0, 13, 0) {real, imag} */,
  {32'h3fb8e631, 32'hc0b1855e} /* (0, 12, 31) {real, imag} */,
  {32'h40c4be5e, 32'h3f2d4678} /* (0, 12, 30) {real, imag} */,
  {32'h410ea9fd, 32'h4105a03a} /* (0, 12, 29) {real, imag} */,
  {32'h4117145c, 32'h409278ca} /* (0, 12, 28) {real, imag} */,
  {32'h40ed5f86, 32'h3e026a28} /* (0, 12, 27) {real, imag} */,
  {32'h40f6e67c, 32'hc0372cc5} /* (0, 12, 26) {real, imag} */,
  {32'h410282aa, 32'hc120fc30} /* (0, 12, 25) {real, imag} */,
  {32'h40de6ed6, 32'hc0efa9a0} /* (0, 12, 24) {real, imag} */,
  {32'h3f859e8c, 32'hc15926c2} /* (0, 12, 23) {real, imag} */,
  {32'h402f9eb0, 32'hc11d7454} /* (0, 12, 22) {real, imag} */,
  {32'hbe3d1740, 32'hc03adf86} /* (0, 12, 21) {real, imag} */,
  {32'hc0b930c4, 32'hc1077fd2} /* (0, 12, 20) {real, imag} */,
  {32'h40bd7eb8, 32'hc02131f0} /* (0, 12, 19) {real, imag} */,
  {32'h4058ac30, 32'hbfbf6b40} /* (0, 12, 18) {real, imag} */,
  {32'hbfb644ae, 32'h40d9a5f6} /* (0, 12, 17) {real, imag} */,
  {32'hc037f726, 32'h400c8f4c} /* (0, 12, 16) {real, imag} */,
  {32'hbec8ca10, 32'hc0f1f0dd} /* (0, 12, 15) {real, imag} */,
  {32'h3d9e9a9b, 32'hc137b988} /* (0, 12, 14) {real, imag} */,
  {32'h40ec7810, 32'hc0541fbc} /* (0, 12, 13) {real, imag} */,
  {32'hc0094878, 32'h3fc3b924} /* (0, 12, 12) {real, imag} */,
  {32'hc0834848, 32'hc103fe34} /* (0, 12, 11) {real, imag} */,
  {32'h3fce50a0, 32'hc1040ecf} /* (0, 12, 10) {real, imag} */,
  {32'h4035aaad, 32'h402dc31f} /* (0, 12, 9) {real, imag} */,
  {32'h40942eaf, 32'hbf8340d4} /* (0, 12, 8) {real, imag} */,
  {32'h4071ebba, 32'hbffc0208} /* (0, 12, 7) {real, imag} */,
  {32'h40ca6826, 32'h4053c1ac} /* (0, 12, 6) {real, imag} */,
  {32'h40be4777, 32'h4000cf04} /* (0, 12, 5) {real, imag} */,
  {32'h40a451aa, 32'h4015d18c} /* (0, 12, 4) {real, imag} */,
  {32'h4077f27e, 32'h408c11d2} /* (0, 12, 3) {real, imag} */,
  {32'h3f05a370, 32'h404559d0} /* (0, 12, 2) {real, imag} */,
  {32'h40a10309, 32'hc090fa85} /* (0, 12, 1) {real, imag} */,
  {32'h401a04ed, 32'hc03afba9} /* (0, 12, 0) {real, imag} */,
  {32'h40513778, 32'h4096b00e} /* (0, 11, 31) {real, imag} */,
  {32'h404969d4, 32'h40cea429} /* (0, 11, 30) {real, imag} */,
  {32'hc05d7c94, 32'hc0227eee} /* (0, 11, 29) {real, imag} */,
  {32'hbd663380, 32'hc0bc7bf7} /* (0, 11, 28) {real, imag} */,
  {32'h40eab7db, 32'hc02cd4b9} /* (0, 11, 27) {real, imag} */,
  {32'h4086b1fe, 32'h41053db4} /* (0, 11, 26) {real, imag} */,
  {32'h4060947e, 32'hc07945f0} /* (0, 11, 25) {real, imag} */,
  {32'h408ca9bb, 32'h406d10f4} /* (0, 11, 24) {real, imag} */,
  {32'hc0dd9343, 32'h4013a8b9} /* (0, 11, 23) {real, imag} */,
  {32'hc10d06ee, 32'hc0472849} /* (0, 11, 22) {real, imag} */,
  {32'h40f3a6ae, 32'hc0a604b8} /* (0, 11, 21) {real, imag} */,
  {32'hbfac6694, 32'hc084589b} /* (0, 11, 20) {real, imag} */,
  {32'hc09704c0, 32'hbf13e414} /* (0, 11, 19) {real, imag} */,
  {32'hc07b6a62, 32'hc08dcd63} /* (0, 11, 18) {real, imag} */,
  {32'hbfe6f1c8, 32'hbf3c44ec} /* (0, 11, 17) {real, imag} */,
  {32'hc0bffa46, 32'h3bf68e00} /* (0, 11, 16) {real, imag} */,
  {32'hc006a7ac, 32'h3fe8c0f4} /* (0, 11, 15) {real, imag} */,
  {32'h401edba9, 32'hc0375006} /* (0, 11, 14) {real, imag} */,
  {32'hbdc394a0, 32'hbf8e3774} /* (0, 11, 13) {real, imag} */,
  {32'h410ba8b8, 32'h40aaa3b4} /* (0, 11, 12) {real, imag} */,
  {32'h40e4e9e5, 32'hc02774a8} /* (0, 11, 11) {real, imag} */,
  {32'h3ff33a62, 32'hc040c867} /* (0, 11, 10) {real, imag} */,
  {32'h40ace95c, 32'hbf93e08c} /* (0, 11, 9) {real, imag} */,
  {32'hbd8809c0, 32'hc0b76019} /* (0, 11, 8) {real, imag} */,
  {32'hc0957ec0, 32'hc135ca48} /* (0, 11, 7) {real, imag} */,
  {32'hc13074f1, 32'hbfb5d438} /* (0, 11, 6) {real, imag} */,
  {32'hc0fbdc44, 32'hc0152aa0} /* (0, 11, 5) {real, imag} */,
  {32'h40dd5510, 32'hbfeec388} /* (0, 11, 4) {real, imag} */,
  {32'h41263c58, 32'hc0b077b7} /* (0, 11, 3) {real, imag} */,
  {32'hc010c454, 32'hc08da35d} /* (0, 11, 2) {real, imag} */,
  {32'hc03e7ad1, 32'hc1205fee} /* (0, 11, 1) {real, imag} */,
  {32'hc0543f08, 32'hc06b44a6} /* (0, 11, 0) {real, imag} */,
  {32'h4024af10, 32'hc14080f2} /* (0, 10, 31) {real, imag} */,
  {32'hc050955e, 32'hc1406070} /* (0, 10, 30) {real, imag} */,
  {32'hbfc4089c, 32'h402af6f4} /* (0, 10, 29) {real, imag} */,
  {32'h40beb112, 32'h409a21ba} /* (0, 10, 28) {real, imag} */,
  {32'h3da8b300, 32'hc08b3de3} /* (0, 10, 27) {real, imag} */,
  {32'hc039fa1c, 32'h4035ca39} /* (0, 10, 26) {real, imag} */,
  {32'hc067865a, 32'h411965a2} /* (0, 10, 25) {real, imag} */,
  {32'hc19c89cc, 32'h412fed4c} /* (0, 10, 24) {real, imag} */,
  {32'hc0b89ea8, 32'h4050d898} /* (0, 10, 23) {real, imag} */,
  {32'hc08070b8, 32'hc0d1ab1d} /* (0, 10, 22) {real, imag} */,
  {32'hc1297acc, 32'h404984bc} /* (0, 10, 21) {real, imag} */,
  {32'hc09bbc86, 32'h3ec916a4} /* (0, 10, 20) {real, imag} */,
  {32'hbee9b528, 32'h41577e06} /* (0, 10, 19) {real, imag} */,
  {32'h40bf6372, 32'h40017cd8} /* (0, 10, 18) {real, imag} */,
  {32'h40a013c6, 32'hc111cec3} /* (0, 10, 17) {real, imag} */,
  {32'hc0f869c0, 32'h40f8f71e} /* (0, 10, 16) {real, imag} */,
  {32'h412ec744, 32'h41029aac} /* (0, 10, 15) {real, imag} */,
  {32'h411b5de8, 32'hbfa477f1} /* (0, 10, 14) {real, imag} */,
  {32'hc0699ad6, 32'h40cb20d2} /* (0, 10, 13) {real, imag} */,
  {32'h3fbd727d, 32'h41067b3d} /* (0, 10, 12) {real, imag} */,
  {32'hbfd943dc, 32'h40d0827e} /* (0, 10, 11) {real, imag} */,
  {32'hc0b68bb6, 32'h4141fab8} /* (0, 10, 10) {real, imag} */,
  {32'hc0998dbf, 32'hc1194f30} /* (0, 10, 9) {real, imag} */,
  {32'h407d0c98, 32'hc1b682f2} /* (0, 10, 8) {real, imag} */,
  {32'h408aa9b8, 32'hc18b92b2} /* (0, 10, 7) {real, imag} */,
  {32'h406b95ca, 32'hc0db24b9} /* (0, 10, 6) {real, imag} */,
  {32'h41278e96, 32'h40a9c4fe} /* (0, 10, 5) {real, imag} */,
  {32'h4029d17a, 32'h412d3a00} /* (0, 10, 4) {real, imag} */,
  {32'h40538a66, 32'h4085805b} /* (0, 10, 3) {real, imag} */,
  {32'hc089cb0b, 32'h41041476} /* (0, 10, 2) {real, imag} */,
  {32'hc120b477, 32'h3fb857dc} /* (0, 10, 1) {real, imag} */,
  {32'hc02a59b6, 32'hc11ec35e} /* (0, 10, 0) {real, imag} */,
  {32'hc0fc7024, 32'h40304360} /* (0, 9, 31) {real, imag} */,
  {32'hc10f8c4c, 32'hbdb35b00} /* (0, 9, 30) {real, imag} */,
  {32'hc1aed052, 32'h411b4b11} /* (0, 9, 29) {real, imag} */,
  {32'hc1a4bbd6, 32'h40ecbbbc} /* (0, 9, 28) {real, imag} */,
  {32'hc1b5951f, 32'h404e9fd0} /* (0, 9, 27) {real, imag} */,
  {32'hc1d9f7c4, 32'h41484c96} /* (0, 9, 26) {real, imag} */,
  {32'hc1bd0a0a, 32'h40ab0064} /* (0, 9, 25) {real, imag} */,
  {32'hc17b1402, 32'hc04bc2a4} /* (0, 9, 24) {real, imag} */,
  {32'hc1950569, 32'hc1517e02} /* (0, 9, 23) {real, imag} */,
  {32'hc01c0975, 32'hc1355310} /* (0, 9, 22) {real, imag} */,
  {32'hc0cf54df, 32'hc1825bab} /* (0, 9, 21) {real, imag} */,
  {32'h3f9f7110, 32'hc13315d5} /* (0, 9, 20) {real, imag} */,
  {32'h40a7f5de, 32'hc0d2e4b5} /* (0, 9, 19) {real, imag} */,
  {32'h414ae82d, 32'h40b07548} /* (0, 9, 18) {real, imag} */,
  {32'h410166c8, 32'hc10b7af3} /* (0, 9, 17) {real, imag} */,
  {32'h40ebb65e, 32'hc1832ed2} /* (0, 9, 16) {real, imag} */,
  {32'hc10e9d21, 32'h4084d1af} /* (0, 9, 15) {real, imag} */,
  {32'h4052e896, 32'h40f76aaf} /* (0, 9, 14) {real, imag} */,
  {32'h40fc2672, 32'hbfb1ef8a} /* (0, 9, 13) {real, imag} */,
  {32'h406402e7, 32'h4042a975} /* (0, 9, 12) {real, imag} */,
  {32'h41396145, 32'h40f3d21c} /* (0, 9, 11) {real, imag} */,
  {32'h40b7f7c4, 32'h4078b9f0} /* (0, 9, 10) {real, imag} */,
  {32'hbe95f8e8, 32'hbfacc8a8} /* (0, 9, 9) {real, imag} */,
  {32'h40f95a59, 32'h40b2bafc} /* (0, 9, 8) {real, imag} */,
  {32'h406b0b54, 32'h40fb3977} /* (0, 9, 7) {real, imag} */,
  {32'h4093b4bf, 32'hbfa0b8f6} /* (0, 9, 6) {real, imag} */,
  {32'h415d9c92, 32'h40ac505a} /* (0, 9, 5) {real, imag} */,
  {32'h416357a0, 32'h407e1f70} /* (0, 9, 4) {real, imag} */,
  {32'h40f67a20, 32'hc18fb97d} /* (0, 9, 3) {real, imag} */,
  {32'h40b58da3, 32'hc13a4a12} /* (0, 9, 2) {real, imag} */,
  {32'hc08a7a9e, 32'hc0c85d1b} /* (0, 9, 1) {real, imag} */,
  {32'hc133de30, 32'h40fc8377} /* (0, 9, 0) {real, imag} */,
  {32'hc0b95eee, 32'h40a622ca} /* (0, 8, 31) {real, imag} */,
  {32'hc10de8d4, 32'h41ae9fbc} /* (0, 8, 30) {real, imag} */,
  {32'hc15578d0, 32'h409ccfc5} /* (0, 8, 29) {real, imag} */,
  {32'h4027804f, 32'hc12f9854} /* (0, 8, 28) {real, imag} */,
  {32'h40f9ef76, 32'hc05a88b5} /* (0, 8, 27) {real, imag} */,
  {32'hc0a1e034, 32'h3fb02a84} /* (0, 8, 26) {real, imag} */,
  {32'hc18b4bde, 32'hc1563683} /* (0, 8, 25) {real, imag} */,
  {32'hc14b713c, 32'hc092fc1d} /* (0, 8, 24) {real, imag} */,
  {32'hbcb5de00, 32'h3f0ff0e7} /* (0, 8, 23) {real, imag} */,
  {32'hbd63b600, 32'h4103fbb0} /* (0, 8, 22) {real, imag} */,
  {32'h416f8a40, 32'h4174680a} /* (0, 8, 21) {real, imag} */,
  {32'hc032754c, 32'hc0a8584c} /* (0, 8, 20) {real, imag} */,
  {32'h409967c1, 32'hc1392dda} /* (0, 8, 19) {real, imag} */,
  {32'h42112b36, 32'h3f6bdef0} /* (0, 8, 18) {real, imag} */,
  {32'h419ab9ca, 32'h41026c22} /* (0, 8, 17) {real, imag} */,
  {32'hc021a5ac, 32'h410e7d87} /* (0, 8, 16) {real, imag} */,
  {32'hc1363a40, 32'h3fef48ae} /* (0, 8, 15) {real, imag} */,
  {32'hc136991a, 32'h41081baa} /* (0, 8, 14) {real, imag} */,
  {32'hc17fa5d8, 32'h40b77d3e} /* (0, 8, 13) {real, imag} */,
  {32'hbff15816, 32'hc17fe27a} /* (0, 8, 12) {real, imag} */,
  {32'hc0b59fb4, 32'hc12c03b4} /* (0, 8, 11) {real, imag} */,
  {32'h40bdf59d, 32'hbfe479f8} /* (0, 8, 10) {real, imag} */,
  {32'h41a9ddfe, 32'h40e8634c} /* (0, 8, 9) {real, imag} */,
  {32'h3f037910, 32'h4048edd2} /* (0, 8, 8) {real, imag} */,
  {32'hc0df2e74, 32'h415abac2} /* (0, 8, 7) {real, imag} */,
  {32'h41387acf, 32'h40c36277} /* (0, 8, 6) {real, imag} */,
  {32'hc101538a, 32'hc1a3e1b6} /* (0, 8, 5) {real, imag} */,
  {32'hc16bc76f, 32'h3f477b40} /* (0, 8, 4) {real, imag} */,
  {32'h402cdfb8, 32'h4100f028} /* (0, 8, 3) {real, imag} */,
  {32'hc08d2f82, 32'hc0b7f654} /* (0, 8, 2) {real, imag} */,
  {32'hc17fc9bd, 32'hc174d2d7} /* (0, 8, 1) {real, imag} */,
  {32'hc0faaac0, 32'hbf96e382} /* (0, 8, 0) {real, imag} */,
  {32'hc10c2e4c, 32'hc1b097d6} /* (0, 7, 31) {real, imag} */,
  {32'h3f0a8520, 32'hc20a568e} /* (0, 7, 30) {real, imag} */,
  {32'h41654a90, 32'hc04b5970} /* (0, 7, 29) {real, imag} */,
  {32'h4154100c, 32'hc1392b48} /* (0, 7, 28) {real, imag} */,
  {32'h4131ff2a, 32'hc122ded2} /* (0, 7, 27) {real, imag} */,
  {32'h4114d3e0, 32'h419b1c79} /* (0, 7, 26) {real, imag} */,
  {32'hc0bd8c72, 32'h414dcd1a} /* (0, 7, 25) {real, imag} */,
  {32'hc1402f7a, 32'hc1aaa542} /* (0, 7, 24) {real, imag} */,
  {32'hc10de720, 32'hc10f9252} /* (0, 7, 23) {real, imag} */,
  {32'hc04c3225, 32'h41197630} /* (0, 7, 22) {real, imag} */,
  {32'h4062d56a, 32'hc11ccaa5} /* (0, 7, 21) {real, imag} */,
  {32'h40567ea2, 32'hc1514985} /* (0, 7, 20) {real, imag} */,
  {32'hbf8920aa, 32'hc0396832} /* (0, 7, 19) {real, imag} */,
  {32'h40cb2c4e, 32'h40cff380} /* (0, 7, 18) {real, imag} */,
  {32'h3f9a1fe4, 32'hc11fbfb9} /* (0, 7, 17) {real, imag} */,
  {32'h406b4590, 32'hc20fdb11} /* (0, 7, 16) {real, imag} */,
  {32'h411edfe1, 32'hc1815aaa} /* (0, 7, 15) {real, imag} */,
  {32'hbfb3edbc, 32'hc0b57a41} /* (0, 7, 14) {real, imag} */,
  {32'hc08ea492, 32'h40540e07} /* (0, 7, 13) {real, imag} */,
  {32'h402612af, 32'h41266dfc} /* (0, 7, 12) {real, imag} */,
  {32'h40479b8c, 32'h40c1dcc2} /* (0, 7, 11) {real, imag} */,
  {32'h3ef107a0, 32'h4119c6ae} /* (0, 7, 10) {real, imag} */,
  {32'hc0bdcb34, 32'hbe358880} /* (0, 7, 9) {real, imag} */,
  {32'h4099f20f, 32'h4110ab20} /* (0, 7, 8) {real, imag} */,
  {32'h40215a08, 32'h4179fab8} /* (0, 7, 7) {real, imag} */,
  {32'h4125822e, 32'hc05e759d} /* (0, 7, 6) {real, imag} */,
  {32'hc09cc270, 32'hc1ab0452} /* (0, 7, 5) {real, imag} */,
  {32'hc1342a30, 32'hc15ed2a4} /* (0, 7, 4) {real, imag} */,
  {32'hc1472384, 32'h3f94ae20} /* (0, 7, 3) {real, imag} */,
  {32'hc04ae7ce, 32'h419a039c} /* (0, 7, 2) {real, imag} */,
  {32'h3f7c2a24, 32'h41617d04} /* (0, 7, 1) {real, imag} */,
  {32'hc13a49dc, 32'h4156df14} /* (0, 7, 0) {real, imag} */,
  {32'h40abe9f4, 32'hbfba8674} /* (0, 6, 31) {real, imag} */,
  {32'h407ea19a, 32'hc1518016} /* (0, 6, 30) {real, imag} */,
  {32'h4082af13, 32'h40457906} /* (0, 6, 29) {real, imag} */,
  {32'hc0283f44, 32'h418a728c} /* (0, 6, 28) {real, imag} */,
  {32'hc0980bd8, 32'h4141fcf2} /* (0, 6, 27) {real, imag} */,
  {32'hc1136e22, 32'h4017e697} /* (0, 6, 26) {real, imag} */,
  {32'hbf329a58, 32'h418a7178} /* (0, 6, 25) {real, imag} */,
  {32'hc11b68d4, 32'h4065e46e} /* (0, 6, 24) {real, imag} */,
  {32'h4124e1d4, 32'hc0528798} /* (0, 6, 23) {real, imag} */,
  {32'h419d220b, 32'h3eafdaf0} /* (0, 6, 22) {real, imag} */,
  {32'h40f435b3, 32'h406f7b10} /* (0, 6, 21) {real, imag} */,
  {32'hc1681f9d, 32'hc03d4ce4} /* (0, 6, 20) {real, imag} */,
  {32'hc09a8cfe, 32'h3ec24310} /* (0, 6, 19) {real, imag} */,
  {32'h41164a0c, 32'h414682bc} /* (0, 6, 18) {real, imag} */,
  {32'h41453ce9, 32'hc191d25a} /* (0, 6, 17) {real, imag} */,
  {32'hc01b4a98, 32'hc12c8247} /* (0, 6, 16) {real, imag} */,
  {32'hc130fa0c, 32'h3ea32c70} /* (0, 6, 15) {real, imag} */,
  {32'h4030a1d6, 32'h40707554} /* (0, 6, 14) {real, imag} */,
  {32'h41290fa6, 32'hc11b1527} /* (0, 6, 13) {real, imag} */,
  {32'h3ff7addf, 32'hc1c62d86} /* (0, 6, 12) {real, imag} */,
  {32'hc0d315f9, 32'hc0fbc182} /* (0, 6, 11) {real, imag} */,
  {32'h40d4b054, 32'h4007baf0} /* (0, 6, 10) {real, imag} */,
  {32'h410f03ee, 32'h40533bf0} /* (0, 6, 9) {real, imag} */,
  {32'h41536154, 32'hc189941e} /* (0, 6, 8) {real, imag} */,
  {32'h417693cc, 32'hc12051cf} /* (0, 6, 7) {real, imag} */,
  {32'h410c9730, 32'h4156a1ba} /* (0, 6, 6) {real, imag} */,
  {32'h40ca71e0, 32'h414432b1} /* (0, 6, 5) {real, imag} */,
  {32'hc06d1fd2, 32'h412c7bfc} /* (0, 6, 4) {real, imag} */,
  {32'hc0b8ea3d, 32'h4117f2c6} /* (0, 6, 3) {real, imag} */,
  {32'h4054b226, 32'hc0c42358} /* (0, 6, 2) {real, imag} */,
  {32'hbfb867a8, 32'hbff8b6e4} /* (0, 6, 1) {real, imag} */,
  {32'h40aeb411, 32'hc048b6e9} /* (0, 6, 0) {real, imag} */,
  {32'hc0c30ce6, 32'hbf1b5dac} /* (0, 5, 31) {real, imag} */,
  {32'hc13d8987, 32'hc0b9a83d} /* (0, 5, 30) {real, imag} */,
  {32'hbfb49080, 32'hc12daa16} /* (0, 5, 29) {real, imag} */,
  {32'h3f90d89c, 32'h40c44da3} /* (0, 5, 28) {real, imag} */,
  {32'h4195ab4d, 32'h3fd4ea4e} /* (0, 5, 27) {real, imag} */,
  {32'h3f967c40, 32'h4083a7cb} /* (0, 5, 26) {real, imag} */,
  {32'h3f53d62a, 32'h41e13382} /* (0, 5, 25) {real, imag} */,
  {32'h4080f849, 32'hbfde62d8} /* (0, 5, 24) {real, imag} */,
  {32'h40116796, 32'h4036217f} /* (0, 5, 23) {real, imag} */,
  {32'h406fe84e, 32'h40d08268} /* (0, 5, 22) {real, imag} */,
  {32'hc0076290, 32'hbe95b120} /* (0, 5, 21) {real, imag} */,
  {32'hc112f8d8, 32'h41826869} /* (0, 5, 20) {real, imag} */,
  {32'h3fd36e4c, 32'h40fc6aba} /* (0, 5, 19) {real, imag} */,
  {32'hc07f3540, 32'h3fa560ac} /* (0, 5, 18) {real, imag} */,
  {32'hc1af3352, 32'hbf0f7910} /* (0, 5, 17) {real, imag} */,
  {32'hc1800734, 32'hc0e9f71a} /* (0, 5, 16) {real, imag} */,
  {32'h40664d60, 32'hc18a18e7} /* (0, 5, 15) {real, imag} */,
  {32'hc029825f, 32'hc13ab656} /* (0, 5, 14) {real, imag} */,
  {32'hc093e746, 32'hc1519122} /* (0, 5, 13) {real, imag} */,
  {32'h40ca5895, 32'hc1ceb184} /* (0, 5, 12) {real, imag} */,
  {32'h409ac259, 32'hc1ae493a} /* (0, 5, 11) {real, imag} */,
  {32'hc0be94f8, 32'h411d803f} /* (0, 5, 10) {real, imag} */,
  {32'hc18995cd, 32'h41350258} /* (0, 5, 9) {real, imag} */,
  {32'hc080a683, 32'h411cfa76} /* (0, 5, 8) {real, imag} */,
  {32'hc128f7dc, 32'h41c5ad94} /* (0, 5, 7) {real, imag} */,
  {32'hc147a7b1, 32'h41527da7} /* (0, 5, 6) {real, imag} */,
  {32'hc04cc218, 32'h41e44d2c} /* (0, 5, 5) {real, imag} */,
  {32'hc07e2748, 32'h41988b06} /* (0, 5, 4) {real, imag} */,
  {32'hbfd615b0, 32'hc1660ae4} /* (0, 5, 3) {real, imag} */,
  {32'hc052fdda, 32'h4090048d} /* (0, 5, 2) {real, imag} */,
  {32'hbf4ee854, 32'h420f7796} /* (0, 5, 1) {real, imag} */,
  {32'hc12f7c8c, 32'h4199bd75} /* (0, 5, 0) {real, imag} */,
  {32'h3fe4278d, 32'hc18ab184} /* (0, 4, 31) {real, imag} */,
  {32'hbf9d3dfa, 32'hc1281684} /* (0, 4, 30) {real, imag} */,
  {32'h41214547, 32'hc1993c21} /* (0, 4, 29) {real, imag} */,
  {32'hc1050e7c, 32'hc1dab762} /* (0, 4, 28) {real, imag} */,
  {32'hc11d6cd5, 32'h3fe08885} /* (0, 4, 27) {real, imag} */,
  {32'hc0a4d6c8, 32'h4112e86f} /* (0, 4, 26) {real, imag} */,
  {32'h4194035e, 32'hc21724fc} /* (0, 4, 25) {real, imag} */,
  {32'h41e5961c, 32'hc200bfe7} /* (0, 4, 24) {real, imag} */,
  {32'hc0fe57af, 32'h41b613a9} /* (0, 4, 23) {real, imag} */,
  {32'hc1f1da8a, 32'h4162fd40} /* (0, 4, 22) {real, imag} */,
  {32'hc19e793c, 32'h40b2a095} /* (0, 4, 21) {real, imag} */,
  {32'h41bda67d, 32'hc032718e} /* (0, 4, 20) {real, imag} */,
  {32'h41bdf304, 32'h40496e74} /* (0, 4, 19) {real, imag} */,
  {32'hc09b137a, 32'h41f4b8a4} /* (0, 4, 18) {real, imag} */,
  {32'hc09b5a2a, 32'h4146f779} /* (0, 4, 17) {real, imag} */,
  {32'h3dd7aad0, 32'h408a2389} /* (0, 4, 16) {real, imag} */,
  {32'h41509f16, 32'h40bcafdb} /* (0, 4, 15) {real, imag} */,
  {32'h3e8214f9, 32'hc1bc236e} /* (0, 4, 14) {real, imag} */,
  {32'hc1e63c7a, 32'hc1b084bc} /* (0, 4, 13) {real, imag} */,
  {32'hc1fce31d, 32'hc1569ec6} /* (0, 4, 12) {real, imag} */,
  {32'hc1a86b7c, 32'hc15050ec} /* (0, 4, 11) {real, imag} */,
  {32'hc1e57d3a, 32'h41511fcf} /* (0, 4, 10) {real, imag} */,
  {32'hbfe9fd4a, 32'h3f08e0fc} /* (0, 4, 9) {real, imag} */,
  {32'h3fefbb65, 32'hbf631dff} /* (0, 4, 8) {real, imag} */,
  {32'h40bada07, 32'hc1b83ebe} /* (0, 4, 7) {real, imag} */,
  {32'hc0f97d26, 32'hc14625f5} /* (0, 4, 6) {real, imag} */,
  {32'hc189b4df, 32'h409a7fa6} /* (0, 4, 5) {real, imag} */,
  {32'hc0a95f98, 32'h41a752a2} /* (0, 4, 4) {real, imag} */,
  {32'h4110bd5a, 32'h41e84038} /* (0, 4, 3) {real, imag} */,
  {32'hc149a599, 32'h41aa1d4c} /* (0, 4, 2) {real, imag} */,
  {32'hc1973a83, 32'h3fef3087} /* (0, 4, 1) {real, imag} */,
  {32'hc0a6b74e, 32'hc11830ed} /* (0, 4, 0) {real, imag} */,
  {32'h3f845e4c, 32'h414452b0} /* (0, 3, 31) {real, imag} */,
  {32'h4223fb08, 32'h412f8dbf} /* (0, 3, 30) {real, imag} */,
  {32'h41ccc5e8, 32'hc11a5b66} /* (0, 3, 29) {real, imag} */,
  {32'h40fd5c33, 32'hc12384ce} /* (0, 3, 28) {real, imag} */,
  {32'h409dd54a, 32'h3ea5e4f0} /* (0, 3, 27) {real, imag} */,
  {32'hc1315f28, 32'hc111cac8} /* (0, 3, 26) {real, imag} */,
  {32'h41e905a8, 32'h408415a1} /* (0, 3, 25) {real, imag} */,
  {32'h422cfdb8, 32'h4144ae7a} /* (0, 3, 24) {real, imag} */,
  {32'h419de178, 32'h416fc3ae} /* (0, 3, 23) {real, imag} */,
  {32'h403f4b3e, 32'hc0ffa333} /* (0, 3, 22) {real, imag} */,
  {32'hc1a0628e, 32'hc1ce70d0} /* (0, 3, 21) {real, imag} */,
  {32'hc1223295, 32'hc115d7af} /* (0, 3, 20) {real, imag} */,
  {32'h40a6e4e4, 32'h41a0cfce} /* (0, 3, 19) {real, imag} */,
  {32'h40170e5d, 32'hbfc69c4b} /* (0, 3, 18) {real, imag} */,
  {32'h40027d90, 32'h40f8310f} /* (0, 3, 17) {real, imag} */,
  {32'h419e46e6, 32'h41acde76} /* (0, 3, 16) {real, imag} */,
  {32'h418575dd, 32'h418b41cb} /* (0, 3, 15) {real, imag} */,
  {32'h40d18d4c, 32'hc003b8f8} /* (0, 3, 14) {real, imag} */,
  {32'h412df48a, 32'hc102cfe7} /* (0, 3, 13) {real, imag} */,
  {32'h4034f920, 32'h411cbbc2} /* (0, 3, 12) {real, imag} */,
  {32'h41ae9522, 32'h405f6144} /* (0, 3, 11) {real, imag} */,
  {32'hc00656fc, 32'h40d22b4c} /* (0, 3, 10) {real, imag} */,
  {32'hc1645fd0, 32'hbfa2ef50} /* (0, 3, 9) {real, imag} */,
  {32'hc1871ce6, 32'hc19d4b0a} /* (0, 3, 8) {real, imag} */,
  {32'hc0da7b3a, 32'hc0601197} /* (0, 3, 7) {real, imag} */,
  {32'h41283fc5, 32'h40748c28} /* (0, 3, 6) {real, imag} */,
  {32'hc1422ef2, 32'hbea56470} /* (0, 3, 5) {real, imag} */,
  {32'hc10e5ad6, 32'hbcdbd180} /* (0, 3, 4) {real, imag} */,
  {32'h40f0b142, 32'hc02e9b4e} /* (0, 3, 3) {real, imag} */,
  {32'h4178fa53, 32'h3f9712e1} /* (0, 3, 2) {real, imag} */,
  {32'hc0baff95, 32'h41a5939d} /* (0, 3, 1) {real, imag} */,
  {32'hc1234a3c, 32'h40d5e75c} /* (0, 3, 0) {real, imag} */,
  {32'hbdbfd7b0, 32'h40afeae7} /* (0, 2, 31) {real, imag} */,
  {32'hc1805a84, 32'h3f44cd40} /* (0, 2, 30) {real, imag} */,
  {32'hc1087efe, 32'h419112ec} /* (0, 2, 29) {real, imag} */,
  {32'h40afda84, 32'h412466c3} /* (0, 2, 28) {real, imag} */,
  {32'hbeb3e640, 32'hbfa65702} /* (0, 2, 27) {real, imag} */,
  {32'h4081ace9, 32'h40a333b0} /* (0, 2, 26) {real, imag} */,
  {32'h412df720, 32'hc0e52612} /* (0, 2, 25) {real, imag} */,
  {32'h413f5fb4, 32'hc1913c3c} /* (0, 2, 24) {real, imag} */,
  {32'hbeeed2b4, 32'hc055c944} /* (0, 2, 23) {real, imag} */,
  {32'hc17b7863, 32'h40eaea8a} /* (0, 2, 22) {real, imag} */,
  {32'h41188d67, 32'hbfc928ac} /* (0, 2, 21) {real, imag} */,
  {32'hc151b16d, 32'hc08d3256} /* (0, 2, 20) {real, imag} */,
  {32'hc193032c, 32'hc11581e2} /* (0, 2, 19) {real, imag} */,
  {32'h3fef19c2, 32'hbfd054d0} /* (0, 2, 18) {real, imag} */,
  {32'h3f89e3e4, 32'h406f03b0} /* (0, 2, 17) {real, imag} */,
  {32'h4164baea, 32'h4089dac0} /* (0, 2, 16) {real, imag} */,
  {32'h3f937da6, 32'hc05434fa} /* (0, 2, 15) {real, imag} */,
  {32'h3e831acc, 32'hc1fe050b} /* (0, 2, 14) {real, imag} */,
  {32'h400017e3, 32'hc203a35e} /* (0, 2, 13) {real, imag} */,
  {32'hc161fd96, 32'h4107b250} /* (0, 2, 12) {real, imag} */,
  {32'h401b8e9c, 32'h41fee6d2} /* (0, 2, 11) {real, imag} */,
  {32'h419aaa82, 32'h4194d4b9} /* (0, 2, 10) {real, imag} */,
  {32'h419e8bfd, 32'hc17ad3e1} /* (0, 2, 9) {real, imag} */,
  {32'hc16ee821, 32'hbee6a150} /* (0, 2, 8) {real, imag} */,
  {32'hc24253e4, 32'hbf875007} /* (0, 2, 7) {real, imag} */,
  {32'hc1a3d3fc, 32'hc0a9909b} /* (0, 2, 6) {real, imag} */,
  {32'hc12f17d2, 32'h4102efaa} /* (0, 2, 5) {real, imag} */,
  {32'hc144ac48, 32'h413b53e6} /* (0, 2, 4) {real, imag} */,
  {32'hc113a294, 32'h40171f79} /* (0, 2, 3) {real, imag} */,
  {32'h412ef954, 32'hc1a78a2a} /* (0, 2, 2) {real, imag} */,
  {32'h418a76fb, 32'hc0224890} /* (0, 2, 1) {real, imag} */,
  {32'h41742e1c, 32'h408d7124} /* (0, 2, 0) {real, imag} */,
  {32'hc03cbde5, 32'h404160be} /* (0, 1, 31) {real, imag} */,
  {32'h3fbe9f02, 32'h4182326f} /* (0, 1, 30) {real, imag} */,
  {32'hc1855454, 32'h4144e5c8} /* (0, 1, 29) {real, imag} */,
  {32'hc127b75c, 32'h3fcd4dc6} /* (0, 1, 28) {real, imag} */,
  {32'h4141b6bb, 32'hc14379ed} /* (0, 1, 27) {real, imag} */,
  {32'hc0efa0ea, 32'h404a22d4} /* (0, 1, 26) {real, imag} */,
  {32'h408bf19e, 32'h41d10244} /* (0, 1, 25) {real, imag} */,
  {32'h4136907c, 32'h409ef32c} /* (0, 1, 24) {real, imag} */,
  {32'hc0e8f0eb, 32'hc19444af} /* (0, 1, 23) {real, imag} */,
  {32'hc005942e, 32'hc2195d50} /* (0, 1, 22) {real, imag} */,
  {32'h40d1e47e, 32'hc0b23444} /* (0, 1, 21) {real, imag} */,
  {32'h41801916, 32'h4030fe69} /* (0, 1, 20) {real, imag} */,
  {32'h41afecac, 32'h41cdacca} /* (0, 1, 19) {real, imag} */,
  {32'hc1161778, 32'h41b001be} /* (0, 1, 18) {real, imag} */,
  {32'h4115cf1b, 32'hc0a981f9} /* (0, 1, 17) {real, imag} */,
  {32'hc10424c2, 32'hc1a3817a} /* (0, 1, 16) {real, imag} */,
  {32'hc1c87c3b, 32'h3cdf7e80} /* (0, 1, 15) {real, imag} */,
  {32'hc14854e8, 32'h4103f10c} /* (0, 1, 14) {real, imag} */,
  {32'hc057a3c1, 32'h412b409e} /* (0, 1, 13) {real, imag} */,
  {32'h40c0fb56, 32'h40f84b20} /* (0, 1, 12) {real, imag} */,
  {32'h4168fbd2, 32'h40f00422} /* (0, 1, 11) {real, imag} */,
  {32'h40f23c4d, 32'hc133471a} /* (0, 1, 10) {real, imag} */,
  {32'hc15fe4aa, 32'h417cf879} /* (0, 1, 9) {real, imag} */,
  {32'hc0938b7c, 32'hc15a9780} /* (0, 1, 8) {real, imag} */,
  {32'h40970fd8, 32'hc1f0396d} /* (0, 1, 7) {real, imag} */,
  {32'h4190a623, 32'h41429bc0} /* (0, 1, 6) {real, imag} */,
  {32'h410ae361, 32'h4104233a} /* (0, 1, 5) {real, imag} */,
  {32'h3ed93a18, 32'hc0a2a322} /* (0, 1, 4) {real, imag} */,
  {32'h4180b90c, 32'hbeee7f90} /* (0, 1, 3) {real, imag} */,
  {32'h400876e8, 32'hc0a4c4e7} /* (0, 1, 2) {real, imag} */,
  {32'hc09d8cb4, 32'hc1d62eb4} /* (0, 1, 1) {real, imag} */,
  {32'h407ea3c4, 32'hc1728da4} /* (0, 1, 0) {real, imag} */,
  {32'h41b5ede1, 32'h00000000} /* (0, 0, 31) {real, imag} */,
  {32'hbf0292e8, 32'h00000000} /* (0, 0, 30) {real, imag} */,
  {32'hc1b1ea52, 32'h00000000} /* (0, 0, 29) {real, imag} */,
  {32'hc12f63b4, 32'h00000000} /* (0, 0, 28) {real, imag} */,
  {32'hc09b9b77, 32'h00000000} /* (0, 0, 27) {real, imag} */,
  {32'hc183afc8, 32'h00000000} /* (0, 0, 26) {real, imag} */,
  {32'hc1ff37da, 32'h00000000} /* (0, 0, 25) {real, imag} */,
  {32'hc17d6010, 32'h00000000} /* (0, 0, 24) {real, imag} */,
  {32'h3f85a1bc, 32'h00000000} /* (0, 0, 23) {real, imag} */,
  {32'h42166ecf, 32'h00000000} /* (0, 0, 22) {real, imag} */,
  {32'h42320240, 32'h00000000} /* (0, 0, 21) {real, imag} */,
  {32'h4179a980, 32'h00000000} /* (0, 0, 20) {real, imag} */,
  {32'hc0bab661, 32'h00000000} /* (0, 0, 19) {real, imag} */,
  {32'hc0cea3a4, 32'h00000000} /* (0, 0, 18) {real, imag} */,
  {32'hc14fb45b, 32'h00000000} /* (0, 0, 17) {real, imag} */,
  {32'h3fd33c0c, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'h41444f40, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'h4112297b, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'hc05883c5, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h4051feab, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'hc1a49ce8, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'hc189b85a, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'hbf83fa02, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'h419c7480, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h41f8d44c, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'hc137bd11, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'h41af9456, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'h41a674cc, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'hc1e39340, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'hc1ce3fa6, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'hc1766d94, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'h4121d995, 32'h00000000} /* (0, 0, 0) {real, imag} */};
