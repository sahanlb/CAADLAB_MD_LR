-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
OFY5rzjEQ4giIUzO9t+pImmpEmtaJnEU/NqzuJMnnUho4WNF8S/keAm9Bq011pSp
kPOMqZdzDHMsBHD3oxafO/iM8UN/0cXE4zNA1zJTZ3fjpziNqzOhoA7ec03SeceP
KD2+VE68K0w961OOplUxaixgNUrwpzXoFbsdfEM+P5c=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 19728)
`protect data_block
ZWHDkwtMOTGaDRLsqPJfaOuOPglmLFQmQGVhuUFyUN4V5e9alb01P2jbbO7Svdeu
XZ/PHuxaF9+T5djgnHuZTIEp3EfAyfQBzT3pqOyrUthQteet3o8dhP8MGao9sGX5
ofTIvK1C9qAdabaVYNcRpwAyezQ8FvRt1ENYWyFmsj/ID4B/aNXGZZ6RGHBuEsPp
m/epgueezzIcyCbpG9nEA8yuzSdBctCzLAfzV944xqWQ35kIF++jxiIItwni57Sr
7b0l+nuVRUgUvz1jXZ1JpzCkS3Jjx8INrHDZYQ3N09nbOTTgRbZkWn78E0SmXBxB
YyETWDl+ckSZBg307rOHSQmDZmEhqghIH82Qx+xI84tqirE7Nw5PfrOK+9IlaPjY
/jnJD2sDNhKB886rz4EwmVQ6KCbiB51h1a6ZOjfWPsb+mLqMbhboBQ5yGSwdgSSb
fXcXbRhuZ0jBOpb2XVSUW1iJ7bvKJK9ArY/q/opBfLRpfP5bKACbsFtJFsvRa1Y7
yejM98CdObNNFsHA/b9d+ydcsz2RqLryLf4PE1z+T51lfWDuShwTbCvqfIRe78pu
vIJcfTHrzAiNxU47lBjbPDjW74tGVdCymjHKlDxYy5nx2WCAfB+lMhp5bJtWeRpA
nRt2ACrL5nQhhVr8TOZRpAv5NimbstgP8AE0kN00po7+trTT1171RUFbJ5Ut3YYV
jYAKRt23HxCY8lIKYCVSK2gxKhY68S0I70ct0o28HFVm0sF8hGZHGY5a+EUHCUcB
aswXg81dKdLP8mM41/EmPKw+N4s6uZ6OD+03CXeUi0FmikVK6w8KcuNyJQI+q7UG
uf47iAMsrIJzUIaxqQULfK9ni++jeaGalm7ywunljwI/0M7SJG215WAcCdw/pcqU
6tQ6arVDpRZAMINnrJcCwubuvtZbG9xBXak36mS2oILy9Rgm1trutjPSzVkbMWLA
8wOV8bGpmSnC4hZFlIDH1eLSwqKBK6CHDr5YM27SuUVvuLhnrAjeHYcs1kkUiwY/
6AT/hnGEWGvojBxEiWKkUGvAcNAt6Ug0Hj6zZ38HxZjEU0pJphQxveMHByuJGIPM
CW3YVQtvSd4lMxqvujHnEVUJLsW96UwcSa+RufnHBbyBsbKHOS5+54285GGS8/D+
POdj16B3P4G8UCMBjCmX1tnq7ighIA1A3UVwWWNUzjizYXvEGf7pMUMrV9ZURZEV
tg0XWZ7H8EwqZ7Kwed5tiRZ7V957VXecp3dumFBOuPybNbyLmJadOyfW5pdv3wsK
x/rTN+pju+SuwebfqkeWpFblbtDFA+TE4dQjpvfIi9CXbEk/0pvP2cfDD5+NFeQt
mBlmWwDDBeNP3uiGuAn1r67geNQhME+C0zXNnUzF/t9/lg4iE9zIkY0e1iv0wr86
hQVQ4Rgyy+G+v1cvdGQ662aDOa8EoE4I/Xm7r4gHRc80vhXUIkJrqvL8OKHIKSG0
+pga6ajOOhe8T6Ogj9gh2Zh9vWm7IanEec6syvsHrQPcHxV3RCX4HYYuR81EY3BF
kYpUWHs2BwChyk8ooOOL3WbGy2KwBCjn5MSbbP+vnS7Yq0SOQ+wKQPCGVrlCWqYM
wJusTLgWCmYd3knQRLtGdBpuxG2HV60MRWddaUldDmjvdxORtN8p/znJNYnzIj2j
U+Lj5sHENG+Fjvl6Nj18TqpzPMpaWi6mgAdALaNFkDrmWL9O9+Az9EUUAeEOzyXA
P3II8koCXbYlIh0UYItBebLz513j4CPI4seNWN5Kt4kyBGGtUIARtK6RFe2fS4NY
pMoKQTeMiYxlEjbULW74q/qMF9HAFveYsI5C9IhOiE1IMQxpvirqw6otvFyemMMi
iJfbOEKbv6BiDdbGcmkGRcAjxsEhLr93t46V61txDVHZlFluDWnkoFUjc4gza8UP
9aJB6OY3wh84bFIx6wUtcthik9zw6lCx0Y5NQR9tKKUFA6XAEtsgqDCBrGrp+RJ1
X3rKjS6UOLMDt7R4mThN0kzwV8Ztn1M86IGTaHuf2Tso+/KDmQtOGoy5pakgVpbR
40OrHOrHngXYuG5CgZPohhfnLdT2l2AVvvxvZXM1VOuL5UioqiF5BwUjYzSb0RDu
D7ebiW6hmXXVo3AL2N63GETsD+aeD3uhQhTzgM/54ecIby+6Uzu7WZRrAzOYS8+E
Qo/atgx9QFf3Ty8ED0Bm6oi2HMFJX4lkilsNYAe4VektyKL1guQIhSweiq4tBbMk
hkqgEKZ4zo5jgmUgUwjgxoNNXNfsjCjJ1bhBc0kVRgKMBQETppZgnuIbWnYxsYXI
yNwJRdak9X7yqIjelMfuoQgcIPd5LQSgxmQpCUuG/BnqMU+DhnBy+fRRZX+svxnt
4Hl1v/i7+G40Z8e9X9R7tfJtFEwSMHpcwlNdWfaku351OdeCsNFuSCPRD64efoM5
0Wof5CYkn4L+gTY2odfseQIYHj0kVVLxosBb3ERCn7dcOnKtzisqcUKM38XzzYV2
eytMwFvM36fDKYVLxvP2fJNiL6sJWf94YraPCs+eIdHQkVVEYXkttCv9828zSeIX
E/9crGeiyntOwPuEG9DWB9K5hdfRfV8KiUegd+RaY2kAPxlMg9f5HXke/HaBOtlm
9qjMRlT5T4JGoQYn/Xm472dZ3ujlcTlGFKUSTp0KmLE0kPosLGwUu04D9FnuSUMW
bgvDu1dCVV3aQ6+a9+MItmlw/fIV65B0c+Y3CWQbJgT5UDq16wVxoFlTYZf8vYth
rGQtbsk58Gwq6vShZKM6PjHeG7r3CaH9WzungQp/n36m+8kONX0DynQo9x0OxRed
PcGd2ovIFjF13xHYQVa81r7DzgxvnL7Fr0Ne6oDN+42mFr99dMMvyNHS2w+KuXsX
VAmf7oRafO8wlA6HvkgT1YzGtUTbrmWAikPeQJSEVdaJRpZiuXkcQukIdPD+kseD
hxLOPLlbHTncjJ3OAVabQoxaEfLbxxVQywMYE0XM0OQVh+l6kCNHrbEo7KBKxAW5
kSoV3WFRvcYDZN1azJk7cPOcrNV0UR6GJzbMtjv8+G1sAD4B3fJbdJtb4kkyusXp
L5vfCshNlSF9QLS3lIXeFM8+EoqzH0iMmuAN/XgmZStui1oRxrAhEMXGz1ltFbS3
TIYZnJJ6BdDSlvmn/gYqNCpVm1SdPzJRYYqqOZyH2ufqxslQDa+Hq6FxT2EVSLb/
YvLsY/hHQQqjkWWSJmg0QbWBaGPHyIwmq5XJo/jgaR84TqWc8OhyqSubOVhm5QGy
EwATJWqVfXYWmteJtDxv4RC1PwZHcFoTIrwN5UWrQS5y+Dn9TCBMgWswm08XkrLL
RVxOGhkhOt+THWvk74ReH7+7WXNCRpYqsXlGKIBl7nlyhR9uVgca6lDtZboW8xcQ
qIwdT2vnUNrWeICBcRINX+A/sDxn2Uu3soopJ6VeqqECns1WxBGcYwze4SLqJw2T
Wjdftc9BNW19I2RQ6fHU5UnkNTtcbSIiTdJEHgLtAKa5i3Lg5azGpoEqQW2X/5aV
XrkPtBfuyq+HfWBZasr5Wm42RzoOvbyjC7ukQ+EWQxGOc5GJJuf2S2C6l4AjJ8SZ
ti3yj9P8BhqpdfU/0odAIlVW4rumVgGTZO30/AXoMqT5b9JHPR4S7diSEP8qnwmY
ATd0tAmNDs1qomK7u1MRQToVCM/WVhu422hf00VgTd80OsIA3qv+z6tawr4gh+un
g+Pe6j5E6Kl5kduHFX/B/JReope44cuQfEuK9yXCa/pNlJksA10Q0gz/9KU/jOLj
7gAUTybVYyDRksNhJ1WX6Iaqa0esHGId3XutZjiqMRdHli3VYuqJXfujOWtPekbj
euVPb8g6G/EEtQRgfcROWaaSHBV6VS2mldGpKDbM0ah71+J9rnWEz8gieyLkL72u
LrkkWCuulwdtxeOWZoHnC/AdFxO4/3Jhb8N5VFMKpLE5jRItuEpm2wNQ7khHBjT2
17v78BAioIQ9/k5qJriXd1fBapZKbeZSkMCD47Hkc1KabgPf4gF2u3E9BNY+yayv
/XsqFaWfzlTN75Eix6K/3vrgI7IcW2J+4sUHmuwVVy9rno7vI431kcdHxbfNxMKJ
J8mrrMMreVR2cIcC85LptihgrXIHfgpLVq4t/rVlBqyobolqCzT8YBTgXkBxLFh9
yL8dbt+vN9mSo28QHTQ4ChYpy7X9qqbiW3jtcId4E/ajKvKqDaWYYefLESWqAo7M
20E+zcOHv7W0ZW/wmzIHZ9Bddnu6ZfLfZPu209tprzl9abwrUz0pyuZ652OtG/cf
HQnEily5d8dmTUxLUeUa4GxRjzEOYe8B2JETLFwMzzxmWoyZsCPS3F+aJX12GHFn
JZieRuwEuv3FvXAq4myNmOzl85TGAsFNP7r38Fz+nh9sG1/oKLvWTTWed4vc27Km
4nyik+XZsetP7TxJsLjvOPxgdlvhJNjNjnMFr3jkkDFUjf4WhznJCsurXDpXYn82
p5kOZOXWBXXI5WeT77ZNz0pPs5+/0quD4D+4tWLb13G9ITUlm1NlIfxotfzOBUc8
l/sSJn9DOOgim5l4ydc8YrAf6P8LYJQHG5ZSTW8suCk20mBee0nywHA+idjP51XW
JF0sEEzr7sWR+vhZqP9UieNnqTgIiek/PEh508tU8ncYHUiRjoHQTZKMupHKMmYx
W+oEbvWekn6mk96xfAZ98Lp+hjiTd27vdmtpPXosIQAcKKXcYMhvFCoYE37mN1Fj
H2G0KhhlJojPzGGcHWDRQXjJQ+O9z2g1rVhl6fwWfXw4IsNW6aTxloQBjaXqnA0w
H3E2dycHh9JYeuLvo398GFz9vgYsuS9QqSjsma0ANd4WUeIz9/oycdDnt4fEc9sv
LYyL7kWCSCCEbOybQkpzrKpSGk9xDw8bjoazAvSWFLxAVi601kz98dqMV/bpCxUk
gEnxcbZKZf0GzYBtvNCpYLbBGFJFlKvFv3TkOZ1fpbQgZd3zSR5ufj9/Sba54QVb
6hGwZsjjQFPEerrg91WxvAMG3osGNtjaKjy882gDsiaGOr8lnjvtpFo2zpGgV+M5
wAqrbIhP1AaE5LaheYgq/Zelrrg2ubfntMHvGaWcENIoTf3SVEYRjsHCeRtes6HE
kczRL1Gt2eigYJVXmA6HXRCGCD5RpQT1C1SwkwdtDgbTTXT4UjSNElfDVW62FBb2
gBbRGkL6v6K+oPd6FToICkOKK5lGfAPIxTfudouG+8O8kdR5jlDcKegq8zvNb/wQ
eiE6vGWQot+/SMTUkIVhk8RTxhAcHpI5gfxIHjyc1r7yjxE7baqC9Eh4iM/udT42
VGnI3iShiqWOBpIoZAkQYrAOEQqPOxQ4OOsiS3DlCc7qrBIQ0HV+HLnPChKJZyRY
PjpbY7j1Wd9oKJVqdxNtn1eX3nyMzVVp6NcFncDClpjy+W1vNjW5aDs7lrk9YWof
UNggtVKSqhkhy/sYq146Q3nqGaGKRLFuDoKLyzLZ08oFxOHsdSouk3XImUmj7itx
+1MJAlkcoEbX+j0ZivXn7HHyqHhgvMkbLZUNiwrDsjD0dhRg3Pls518+uwZpqQba
LkXCiXsijjoA7e0TA2gjEEg5zx4G7ofNroFExaoxP6J1mcLXD7ABwPC+Rsb+1Z0L
8o3YBTLEc1a7YfoMc7XYcvIh+TSNbm+fNFgRLZQs8j4IzKp9e/wF1YbLvFyVp+Ar
blxHckwVs70DfqfQ0ORh0vC1hW0Pi3zMXFSBH1H1dkRu2dVi1lTsL4qWY2EBA+mx
Tyth3QX8d6sYIsfVVXm1sPRJ88e+wA6WtLR9eaBcZfGH4iDL/xVCPI68aPGxFdIq
mgeTL0JS03Y3FkmhygOZdFw7/u3YronunmIb475Bx+RCvmM34eRbCnj0+McCfErI
UA4XN/qfMshw8L/Fm1OJyhVbMQbUssRB8UgecocGFZR+/k9vHUXdfD/mHOsosZwd
2r0UtH7If60UoScbf9fyPJSO2MsQZLLNLEOgT2eqok7ED9KT5xVUTxtR/ha8kg7N
qDieipm9ssfG8dVQRa9/J6UP2kOxOSzEcGBEZsDWPIF1Eny+VnI0KmipvcSehrmT
j1c+ZRI2N4UlALZ9K3GoFp3CeKP1Ury5Rrxy0etuYyWEuC74uJ3IZB2yJdjf+euM
AQoX98Ii6KlH75Tr+RFgFM1t4AMXghK8w9s1pTOXfNm89xKc91anyFuQmVTnSqrN
9TJ0+Srvr1EgWTni1kKA9M83qBfp35sxfn7Fx1a3vRuDerZaRFFrZyz7Ll+JDrTD
x2wmbeODsGc8WHVnrHj8TwJPepVJM7On90bFxe/YPSXHgm3i6uOZBRM1IEQKf43y
V6fMjTksqh1ugi2EBVWVJBOULWgA5jWCIpIsDMzlu7H18tSyAr1CxdnKgmk6ln7t
rZqWWQ1CWqoPhsQ2JFkqRZRAQ1L1aSzD12uq+3XqmIKXcJg9riSO+5m8H82WdhNz
HNabWxgY0/89JaMXtMC7rBkrns2xPT6/oGz0fj35mGqE/WdCJlsxJp+qsqcXtmii
4anmWvryzFMk7wmOyirpX6YL91XP94hglfqc7Hk02COgoV7tH0SIS34JyxLlcxC8
UE32VrT46KcHj8pWjy7yN4AIXOjQioJ+qcu4YfShZxdiNlTGX7svPOGCpwXB8MQ0
VAPAQDW7XMkox/BKviYaOSXmout8FAKKHPluCWAJNvF15XgPinEiYNTJsCimz+fZ
uFdLcBxo18ph+4QGP6Sqc5eCC1G/M7x1LxC2Qq8XuKw7qZUr18BKmRHQ2dnXzTWv
hMLjSD+SaEa9n6RAVvHE/oyvdjJYFkwvapYNFo8YL7JPDpUOBTRKsawQP7ruFI0u
lA8Fp0Wt6edw51tFJXzaUtdxphvCiEZoHY91qx/OrBJuRAaOHJ0A6+M5b0HN6Fxv
FlznMiy6BLXQrvvdsSL1GObO3tQVOJlkA7SKrQ+ZrjkqpvgA6MOxXQtRBxRPgauG
exlyzlQPHtsgCPglFS9mR89bjWv9tSCUXdkfvzuLlrFKqt1e/uOl54/JEklTH5eR
7pSTO9rE0tWf1Wrbi+wsBl0IS47uYqltCzZUonAOpkneJKWMgNgn85fI60O4VuTv
JfXeBo0ol5Sp8crDH5fcJBEsuXD0/rX7jyrBMfTZwqz7jKdbR4eVOxgWK99/lly0
c0cjCDfxSlxbLwREfkknaQisJOpDNnBLAMs+uZueA8/WEy5CkFbyP1kwxF5iLSTl
VVJn0ZfgUxAka6yHtiVAiyD7dg5E37F4YGrXs9zSMVnuXE9IpNqw4QdbXQQ6ibLe
V+CVM0unH6nw4NwKKOBRQhDjOgg1DXDpGBFjR3jFpTPW0QdPT561rbChR5PWOkyi
OvwWcTORJuZx+LShcVc/b+7VNpqaK3Ln+8P13Ijmd2a1ilkVwOGI5o5CdYjoUefA
DXScMMQ/g2tpKIxgcDNAFuphzr1zs3nwMwlNGvOndpWYCXghx2PraP0M0UfOZGEq
35m9siCq5k5O+ZJX3BWuRl3EktL3ISfkGFmKds1KvP9IYCNa/O8lYM44NmL9Wx3Z
rFZQ9+HMdY35j940QKspcHqOovPHU6j69fydN/j/4jdzmqR8m12B9J3tbqvl14pT
ilDY2C/+iMfMMj0YNCwXzQehZrSPFa1mCJTu4j3F2Hh9P8TW8ZwgeE247+Uvl/T5
DhP0mos3IXv4qGaJLJ/saUc3TdKcepG0N8y1NqZWHAUzUk+1kjmYW1/t0Fs6kyZJ
Mx1MH+C0cT2sqn9nYYd5N248+Lo/Oohosq+8I2f1F2ZQD5xpwSSFJc5C/6Lfbbaf
N1iuL7XEeIY68LI/FJdUVibmPAoaVL6jBrc3NXkby3efnTvHxorMzMgVtN34J2OX
2TqDXoKcJdl6uzkKIpzoS2a1koZ/U+/J48TH5V+FdY1qEDiJDomcAHOb1OZodsRR
OEUxBb5zM/vQC/6saycXaew5l8f8qOsfp0VeIQmP8mfJFJw3wVntIvsV0hQIuNfJ
tHruxszJnYVXRZfqsCZpxwvpDsH3SI1SzwYugNKHIKTmLFdQgIYkY73aiphk64JN
HBzNhkXfGjUHbg4hD8/15TpKQM63oN83gPvqQ4cTj2tmOpPAMP0CtkYLBCM1Pk1A
1cnxoso1dNVP5dcebUDO6RLDsVIztmtBodI39kbDDtk0ZQUP6PuC0JveeYFgO3R4
kgvzYC1W0uS5R3MB4efERl5VSQDJbTzg0lzUj70g8Fs/Ul31AJipotlc8OuORR03
PoaJW8WNGn8LtNbiZXVyybhQ1c/MZiOj81OLHjNZBWemPWq4v5WkRapkJZ6gh5gv
fozymDuYyxqXs5eCWSlbSZxnxN/u7DeD13+A1bMRgWE4DozzXpRv3Rf+oWXypW96
jD92p2D6MixSuUoklSpRGbr51JniRF/WpLsg6sQEcfC0kM+YkGHEMN+J4BuFffCK
S8ZDU8ViTni+vHczZVJe55r+lpTvO6FeQWcjJGnhK4H2sL0COZFMpR297nmyraEZ
1emTzaV4WmgPnnO4uO9L6QtkQdp8ArwXrNFpTT12ZrDe4ili33RDjtntkh4lJehl
JeEYr6tnyWF8quucINTEBkOTbCC2H6h/xHiOVUZBcr0ga+EVWy/aNrv8kIFLB7GU
fuWGfVuQzsy2NACZnlyVcLjpJySypI2K5auvMYUFY6qDhl8e/pRRVxL+TTfLdNbd
8dq/kIpfNQlGA7wzfcHLQBgGFafU2MpkoUD/2JR6IC/L2jNlkYPAlRB+HvlO5/p8
Nw+VrfuzfFVI2vt/hQNtOwB5Ho+5hZwpqMHMBvX29CmfMQQ9zaB4Zoc9AulkrpOE
SeT/AsLtlekfKeFkf6eu42u7obrgqqDm2uzBXGgbfDSpbhKAGp3tn0ROw+seuR/9
0qO+4MqSROtqs54/M1kAOPN6QLBmfkrDfJggUnrKwuHPUJCmWd8FIz43fRLf2Xyu
sgH34cP9/9ppGk5eHwYGp2AkH2sIl7mB2z1rAg3s3mVLtB+RPSVQwrVL2wdH85wC
hHk+W618Ma7YnfcRUtMvfwv+ZpamqlmOWvhyCRJe8NRXzG6o0TVmBd6j46/8I9SI
ZloqgoiWbI2NZ9K7SkKA9HnXlRiVS3cy7rzvfljCnqhfWE+FjoBKYj4ref77f/7v
kC3R7KBzjCzRfFsx1SciwQiPPCxjwkbXhyVRXMg3Fn8htzNCpxDoJjgAxKJRs6qB
DtdYQwv7OcWjt5tkrfOHQCRbk5yx+KdP3HQf8BE8Rfx60tzLCAr+DHG5bkK2EffI
SiCgbrREFvBt1GIzRxtTgckkLX/WHGWX60CZP0XbVG0Gx16lZjX+4IpAlcCpHhjA
WFA5FTfFpnEyBMm7FnYUdk0dh+mmZMxles8Ez1gUk8+xYRjfdHglXKrJQEPg2tAy
nRQjsQhS0RNYHz+5SlC+UEpycf6eVtH07S79UFWTj59aYZQ3FNh6cNZikNfPSO/M
b54vVv2CWm1HIZmBEdX9N441gq5vNb3224TGpqjt7MewBzzbEB0lL5TG2jOadR3X
fkSBMgDXzARTbqa6UH5y3hbfW2mMROIp9ypv6do4eZxmC/m60yJcBTulVTHEjfG3
2Dr0pijM4tb8gCbQ9liAv0e78e0QslCD8UtVdV3oesvNHgmZ8Bcyr4DBGRUod864
d4a2hmEOcsUnxS6989eLUL/z3M+iLaiL3HW1i3NYUr1m6xCwFi0ZgFAFbzGYAvCN
tlXZhG+3Js214afk8eNeWgcWB05xU67UATpYJHB3vdT41TGfwDzzjxS23HH01Kso
l48K0Wu2to35rseuMLomFs73lRngTDZjkTHYehVeH7t6rglvL6UR5zYpdnSzMWuK
fXEgMjpjEIVvcoj33aExKD3rCtqaYQyyNK20qNp0Gkf4VMSlDWjW04ItgdG1kW4t
v38ihHUsvoZfAXOAG0nf2MGPT4/SYtdz/Akms5nAELL6gCBu2P13YgqebUEj7SPr
qqHYtPRaovLLHdSGXicyhGD2cvEQca4wluFH9+TcJ0aE/l19xvLGsSZH88nSl7zU
qpmBSV2QDTAd9G5Ua1sO1Gr8kOIPYQRxi1uPcTfwFWZYs9l4q2ZzjFf2xB00y3i0
O4VbeDnNs7+/c68szAWyYjHw9Dn/EPfRp0rlxzNMRDZw4idc6fF3Lv/eqaSY6sFg
me7LHvKWU92HFxqQlXCyYgVY/mqFr6oNoaURyIgEEhZRLKU8hzjkJ1bp8CXRH0VK
n3f5LVD5Tkqgb7ZUCloR4kY4CzuCRopFId02NPUG+3y5+UrucLbqyA5H4Bp+0iOQ
Kco/co+lmMQpgEg+oYo2Djx/IIiAuMSaatrL/rk9lRe1qPJgIVRbhvFN3hld/E3J
zpS5adrhJiJo5mSkUe6JzigqBElucaLBX+66NO8CNM75KUkLkRtpW2V+hVwDtukW
MT8VHLJuOFeijDu/1wXjGjlAD3kqFPsBYOlP7YXjiUPETnYVppHnBudW8bLuhx7N
224EpBhgiBDvG014/QbBsw1ZZNnP/In91i4/RA9v8+9zPxKNENJQ/AmV4Fgmkd3T
/2OP3BLaVse8i+nLhnyexHhJPLQ3cbz4PdQ4CFmMl/9eUuauf3qtiUZ3dE98Lpf4
eGKeWgr6ecsMnuFfq7FL9pmgUW3D8NgPVHz2bCXGPj9Wi6svKC0MCK5+s3B97nzx
q55nLgkwMV+zBfUBX0s3NphWZI9YNFEA3VmDmaSoHb0blhs2pV/aXSwIswRjJHOp
GA5ydCeceXOTk99g/p6pSF1QL7yETuuVFtQa4VGExP1UTDUY5qq3a1qOE62i6yuf
NtvsVkYDvuHLOzqHfDBTrTdRlQhT4eulIK9LHX09qhkahu6LNd8Yv766T1uKsHHH
u3apgo6dfK2Je7dgcMraq6Cbh707vrdbKuTQuKFPzu/q0wegrbpFS1NlmtAQT0rx
ODG3XS7ZlTsNYtRysbdvSmYOI4vT28RzbP5+v8lQ4/VbpBkA/lXnvZntMXaYkoyK
Fvf40SX/EfqpmgT/R3a6snnY4XnhhmuCYur1Da/m30ptlzJnfHjarOpOuRxgFUGw
jkHruvQaphgX50XbYWNPJsS188I3YU8RNv0rnRimGB7BHhwlQWTlA2UPry0sA19e
5qD/lQFlTk5Js5uIh/tFOwxsEOQKssYtKUYh9bOUfL11D9ImLDWezsCxQP2nkxns
Yq97rKKKMUwcqDN9DbTTVIPi4zO0SxUsVoD2Tzf8dR5q5uaAtXb+G0biflF6zF5z
Yu8hJdw2piedu1UiPs0d/mNYd8SN3Zk7D2IsggNW8iYSYbak3Imw1ueHLFrp2Goz
jxZA3IMaC0i0SZDZNi7xqfJybZoFDa+hfakT4JspXp6cKoHnm3LUfVMzsRJXz1QI
2sW8HdEextIIIZnmiiujJ8nbYqlr2nFCSvCp0yuxYKZqVZxe3fczmwgrm3+VJxMi
Ir2NI9GvV18X8viwcZPks7dx4uvdfKcl4FxAuGF78m50emi59JmAWOd4ShLynso0
moJ/pTuMMCryCsu8fAhJKDnW1eSFRr3Fv6UJ0hNTms/8oiPpdZyPwL1cugbLBXLx
BKn8Qyfdlhz4fqL4hFBqyu/s9m1Kpo4Pc+irtNsZkRSoE4pSftKcCzT1UVWLL6tI
HAM9/M3xGaFR8wSIWEvrup62I0L+AAo6xol56aYeQ9U8cJfEXsrPJBbf39v2Vgj2
/L3GQ26OUgbwfubEWwcwQeO5Nd/1VfspoBd8NjLFWTyr7UXGwMqVTubniaBw4Yxg
vlg84BidJw4ST1w4pITtaEZWJyuEJOZucEOdCT0O//vokJ5uGFx+rdav7JlSuFZ5
tfw4XJcdZ2mxOMHJlNcGhVfjRZZvEzCgRunMKBSIGAGBy9AJ5MSvP54DObMJoksR
UPhhd+LJZ5WDSGSzJ2327Nk5QvLnroVCfWiYQxru5Ut7WFGop2BS/ZKOkjME/6Ow
aLV/RKZdDyxMSdNKW1n85gNE8nx8g6GpK5CK2C9GD9PaaiUa3y6mRwFkYrtZbhOQ
TAfRdmevuhpTuq+SCHbSOR2QeF2pM2B7sSNDTaVY1av9L0vYXUgzK2wee+1ZlTXn
PP645ay+KMkyB96TUSGlBYMMPFr8xeLcs5t1D4a4j1ZMqnl9oDoo0x8c47p/hBB7
0oWXtTaw9M5hER4HDJLSsTnykyU6/sFmdpuxTyoYP6LW5JyqvvP+kiR0ZK1G9ooo
2LqAheCSKfc4DxZ2PRelVEvHtNK7OrTlgo6Tc0UbDRAOe+sJVkOqS7Wp8tRWPkPg
/RofSybCak7H0ZNCH6g4HD2z0Gb2+eE2gptLd+JC6CcsoJO+7vT7PskNnusSQqHg
LlzckWECmnDfvJon0DSmUfeo/SwdyXO1BFR6K8EKzE08RNI4/MDXS1O6Zj+u4tly
FW4DX6ew8iG9nM2Om089TvF1meTaRHpcb8lWw8sXLjKlZf5AQLp1m0pKijfBurz1
b1zF/hdn+yD8/iC/6Q6w/MJTKvcaavRqkyGlZBske+sYQSfI9/+dWJFj30NH601m
PS7Ow5zmQzX46zXtQ0meP9C/V8Be6LRbNJd3aLzw9OfyoWDrTnT7VvTfB5QIonP/
dPHVzZDPmvPhifktdQ8FxuBO8V3GpzRU7QSVakyy7iZ0q3VqDMywVpNsR3GZ3M6d
Y/MlWb6uq1eRMUAA00AhsxNKDzcBSPAIfyWOmIwLj5t3LCCOrEJnI57EO0nAqaFv
Tl6NE2LEzHtFTEgMZ1CUIxaYjMz9Lm9uBCjCZIFfuPoNDqIMvMDYe4+SRAhHXK4r
je8dgs704jM7kKv1fen3+3TIS8EeT3DJ5T3zOJhOV2k/vi6YJIz0GoP/6hKi9ZRa
/66s8zgSEpIG1Ww9ne8haYIwSRxQwTnPr5i8Os4Pv1o3xpoziy7X/bYyATRQe9AJ
ktHkgv2ts8+NdR4jEZ2hBw7yY5aBG9RSCqsdtyl/tox1SYIJ+F/MO55dNzll8Uiy
V2b+EKPs8kMjuqEvFpFSID3AJhluRAIh5BkwB+Kbcngf5VMdmBgz4v98yhZfQ6ZJ
pM9wd643ethlgVSBdahqilt9hEHJw+D+aw4zDLQ/2nfy9YGwV+uJfmIVA63IRgXn
w3JHjMaP+iz8vZrhgEW6u+XZCNTvyMZ41yZP/6gd3yqRUyJgfxcsBZe+G1NXeYp0
GKWku9L37Kg3YI3RZU5tpyX9VU2zIsnBK0lRBz78Fi3KAhMZPPg3Sxs/2ghEhu6N
2ZwASLTa5IpySV1FruA5bdOD+yizUViSFKZ4KtoVFNvIqb94kZRB3/D+zKy7Jwm3
HKLl0aqugSjSFA/Isc0/1nKwABVqEkIruqqYDagCJ4HoFf93xRUTp4fqDDJcuDPo
40hWZujeoRqH+ilQPSGB/6LVODWIzw+r0H7UFGrxDAcVXq48KgIooR9wluW56D2n
bU1J/siblV7Mp6/RVy1hu5BrBqf84ybXnPQt0+upoMCn5QKhZCcfc+x+ZhY82IDH
BFGU5vQFh31T3S8eCDCmGwflfj7yd5+tTzin++gF7cffYlF5JVSTDmEK39cT+TKT
s7HFSRs7coXLyzODCzCDgI9Rr1evjESmPErH4UeKXtuaFZ0CWh0ELXkanYbTKL82
2Wd7rPMk4DfKRopKZZMwPzwjHyEZG1rTWKpBtjqnTATkEOgt3YgbaVFVcSr8QPYC
vdaBT1p2MW+BWNABWU+Bk7uvazPNzxLhf3oiGSqzkHB5lkFATkX4/IyBVAIqOkrB
fWsqK01RGFSsNO3acux04QYwNlCLysGQlwvtC8wafjYcAJXzX8u+6DlfvaqnZUvR
20HPmSUA4Ha9B0YjgbCQAVBO6XSd1O8Q/aptVvmtvNgYaqRPnZ0s41WobxSSCPtF
JPDM8hBR4hnTfu1kEBsDQSeaVB6sOkja7/D4ny7+wVKTR8EnyNP18D2sEPoAW/uA
1porVWjeynvVwqvBvWgJJOJCAGVPjbfl7XwhzXM76M+kRGt3nClwUavj9futIo/2
qHLX8IlDAb9fNndc5/l32lq8M6Nrmj/rLqItOiyBdjBd8/DMH9ktndZgrMgsJ6zA
G20dEBO8aLlXIUQDzHcFSyYWZRvvttv0oNJc1+ckAIlhHojv21XtKY25IlbMiuiD
SskmGulNLFzi8VUSOq1FPCfTwcUFCzcMsVTml7yTW2dueN+GoLjlSmy88Gx7m3RM
KVNeMQ/5je6wlvIh8D2UNVARQC8cGDFDS0HAvLmM131b7zF+VrI09ULFUiQ7UZs1
q1U9NYY4VA97+AUMC8Y5prHPvqr2b1n/s9mLEU8kJFsBBgR5pU5MN1gdj6+Re9o6
PBQRDe7xKrG2zjQbrQmUhCAcDm2601WxAN+XHwcMAO8BQ7cZRkIqRAGpAPscrWRX
GE4S2o6kmS9+aDA1R3JcYsY1FIYHGtiTgAUcEY/Bq+qbqmbZbh2gPSePD5VaJxwp
9HzdVYQFJcUrtZ9kA50BfimIMSWMqAs3vM/LkEBsWtjAzTWO2q9EylwOifhvMqai
EVEG63xWMGIkHxrlCBV/2QS3TUlgWfXAUezkWfHsxkPaTWSIz3frGS89Jq9W/VeB
gIuJy52ZnLvcoycoegEF4fI+Acnn/01BMFc+7fCGGbKdX/ZIoo2MWZ0KNV38wkQa
cRsZfTJ/4GA8qiMjfebMV+9syD16pO2Cfa/dU5JEwnt8i1tEo/AA99RtiRIcky1c
4+5Q7eWFeoC7FIn4s7CRHExgG8Gp1qjzpxHD93tEtDM7C293SIq7Vxd/PehkCKR1
a8vYd2E/JvJSgBB6t5Vuv0NItZNE43xlA5Li/aRc77adnCrbYkzCek3NJQxW6UyD
0U3nA2P6qqW5Uzlo6Gdkh1T1hoJCiV4bba48q1pOCjNxmBhp2THuYY3V3yNV/Y6i
B70BXvs41/Tkir7GIl3jiFHwZ1sgaGl6Mv9w2DZNPM09PShl+9QpRV+wsvtJjDy5
sMAtGKBIW/CH6IZbEU+LWIJnjIu67L0y6hQnh39umFHFLchq1fw8EXwZo8PkY9+9
bgoMUhJZDWeQsIh5ZKeVGoBd3OU70HNqf2AYvXvknH11wWMHApYWWK/vfioqlVWh
U9dwJP980TTZNgIEi524BY+dsOrGhKg1nCDaBpBZgfWSftKMtgI5Fegjb0j5nWCb
Jxnju0FpCtzKn29IyQlg2/IpDNsR4G0iy7rf4nHFS74wEm/OurMAmLQTQTMWe4bf
mjeOJybXim/aiq5HZW3CVElkzkH65Bx/NoU3c2B7Gm+/Mov7zUpNb/e6eHZtFhaX
XKb1YMN2LMNNf0vyBICt5lLMx1fYuc96ottvnx5HvkCfClczRgqjXNXe1fnaMIad
1euoH5SrfXyyFifnERCVWAlRcwjN32iBsFJWnPhf3Ue3aoHeP5KJjLE9PaOc+eCP
RUm9sET+GsGZ+kvb90dqvNZlsacQNotKR/dH5Zp1wKjxDwbqCcyT47vZoGSVqxcm
BQROCdOHHo5vR3v0hRpVYMpafnom0pyk9599W2Soww9hLCzWLbfGSplx/Q7jx6lm
GFzpL4+wdLJ9x1PLyFDDkNFelVz6wke/TaliSVxIX8OCHNPlsJz5SET6oxH57NVx
6EBNuhchCweP7wWoqdGFRtEXWMW78w3JCKQPLkuO/7xIrzJcjiGsEbeK/EP54f6Z
rN4TYB4VfVuW7OY6ahbhKDaCYwCWaKlyLHrlosbmKOtSpFWqEtzul8Vy17o3Hul1
UqOKDkcrXKgp25ZaZR4/spbNJlZCvMss6o2kHCGwmV/VAKdosQ+KvvjSd2e5BeL/
pZG8yvkW+m1TNx0SubXt7RiP+h7Mi9PqbiQ6xu25PSkZ4R+F9vL4DvRgJMF+FVib
iZ7oPTbgGD7O3KYwe3a6m7kdabuC9WQO20HkMNAyrSpUj6Uv3p+Ze2L35DsV+1GL
D8ZLXa02IR+1+gci8yTIRo8kY3P+pVgTUoFBB8VTGW8tvS0gFq036n8KCFoz9E+W
u/JbPDoMVILpLdndLNGQS6DfM6m1unGElotmstTMZ+ks4np4y71NbyXr+P/60dc+
GvPb8pOYBGBk/YNjIHmX8xK8YwDHxpY/4nyb2TxeRCG9yPaxVssTrNy2ZR1V2Qj5
7XK46GGo8U7km/ah40u97rL6+i067XZCINyC5QEHQMRTnu1EwZ9L4VFgAqq7Ub3T
HIzFL2wMdF+1dIUJwTlqS3nQw+EjQNz/u2oBs2V3q0tfA6nKVGJkd08Ue6y3loxN
8gdZh2DWrOE6Zh1M/o7iA8Vnd1FP7tTiWdtGZHfp9MPTwDk+TvlMw2El2pN4ZKsu
PWmZhlsIqeRqRtFdGV39etSBmezwN4xwMsiGoOlvy9meGLEPVB0PMu+sRBlN/mUA
01DAFf27OLKF/huzUMx6mzX9iMYkaUTJ4+siCJVQ0DvSzRiGorrne3zdnyF3cBp0
FuPf2R/cIJ1xJloO0du9KX0WuvK3nQ1YXBdYCvwak4iXz2VanjxYxKvkX8yRW0sk
PmFJ2v4xpH58HMTqdWO9SBcCaNpVIND0Lloi29Yyqq0+luw+gIIAPMZR9nB8XWdr
g3SucXHVFYY6XlvYd/6CsXnHcab0Hokn/FWKDcXTK2JAc2Npvmp4wQOYCh636qHv
ScpAGRQ/u6tER+l6Ionmm+V6R/s1U3VaiKlOh0P9kiV3hmZZ5aXPu/00W+yzqq6g
4R1pkir3huefv6Rc3QXdb0r/WusgijF5Ho9qMl7wxsLQzEJZCBq8WoaNHSrrN4HW
yeiqcqgc/srK1f0k7PmuMt0AUttpfI8OuFommkyRChWYz2+Uf9rRYchtU+xILvlf
V55c1C8UBai8qhCR26ZDZwz9iHXQHzAygdQ7OznhYvNLqLOVJVM14Ec4ZNnbJJlL
ThLnYHuQR4t/6ucRl3pViz1mQeJzJD+QJ1p5nD9CvyVK8LM7ziUAfC1+PcCExPVn
xGs8ohSeZELWGjQYovtUy6IE2/wqG01c3imtSCV3Kd+VSL/5PxOQfmIPTzYaz+qz
mg3yF6Bydm4zinx0oszk6rXEJQHmiHA33iYKumLGyYPZhHU+A8bnKFmS2XF7cw+u
P4NvQZ8SkptsLzBAWbv4He0+g0xYdpGNpqSD/Zn4QubpMStoK15m1upyWKaVJwA4
1Byl6DcnzHxpu4PCBPnZiQx3EKDZsjmRd2VFDy3nTcJxR/dCRwS7/t67w8KHJbY5
uWz1mDsWvH7U+W+xarU9LJT9qrIvhOSSuJZcADk6H9S8oa9LjMVwVIC+ozjXMcEG
Nfz6DtK+mwfNLMCdDrYpGx1EXlq73dU/8GpWLVIurPpZ+/ifqKrDMW6+92vQwuBU
+MpZ90/Wb5sWAzbE6MAKMuQoueOwwnL/AmEZYDi0Rx/oiVX5fyWSqYsAgh8JUhtj
5b0w8QHU0IO01GKlMXR1YLbF1K5L4ypefhgn631IpHNpJ3BavmHoMn1yy3pBUh5O
1ZUVOBm65nA7OCa66fChLqfqFFid2KTbBV6DVRQFKiawrth6EAGfqZZ1FJmE/08x
i0X535WXKd26R+fUOV0gbUAY/Cy4UziZcQtNPbLSZxHwBB8lxjNw2H/FFxg1RsZc
eKOvD75U7Qe3qDwNsCoYwpd57KvzGm566uJm7FUkz8mRN0iSJCI0KApDUeStHLbr
ahCWndTcxBEygSQSEgCRT58sTOpWnzLJLDXqGe/5MQuU5lBKYdQ1aQQRqj8/N/rc
z2+OCVWcRadyPAdLNG6a6rMILDXGbgq1mLTOpnyXXSGMf/QE5WBWNGvy66QBZUU/
yB5rmTl9eugO3h01TjP7aXAPP2ZB49JE7AJKp73RRC+rtNHG/WwASbmmPFTAwStl
o++PWELDoI8gyuSzAms2r0x/YiyqIVJMFaKqb1OVMD/VT8IwcnaRl4sA4vDrdDXD
MjKmBiCk4wqto1MHWlrJFGhGOK5nA9Ob+YtdpnurTNTsFgNbCi9kcX41osvsl4a5
zp2En7hVLkxfGP/mQ93UCQAaj/VETJ3c4TrIpv42U6VgmYj2Iyurn7eS2891dNHo
etK8lCR87yqjm1kREf8lP3V4bapoJhfSuLFl8V/2IKontJ8kUvMLs7f0Myjy+QWb
qjNxPS7LmdRd7hMLtWsxluzSEupVlzMVVZlzt8HY4yxvno+qYRhHik4Sc/G7e+LD
TsZolZ9P1eebArUxYjNUqFInCWd47N9YfH+yCOaDvA+fxlqZvgCOJduTIQbSoNlM
zabUrlv6ItsA5SdtbrsoKandFy7+yLDnkfwyl1Rk/0drlq4xcnTJ17CLQ/RT9wZi
dsy7kxX4DeKfhn4ky2Z5NYOaLge5zFPsAVeg77D1Kjd5lelLHtMYDbD8GRNkE4gg
gJJoZbx+xaWT4AVbsCSvAM5nOou8cGTGzaHDdnfk9P3N3XnoQlMGspM/XApaV6BK
teEasRZMZv26iIm9QvMwDc0dHMujZ7JwVVXZVpHrv5/kNE/StU1XSpKoqIpFke6k
wb42BZMZ/sCWQ46ThnCUCAjkzmo9cz2i4ln0gmoOpbEhKESRIwgHNTegsRPh8cbP
LTgejTZPq2UgliCbDwBiFQ9rrtdmsf59gwUQKhuEcLqFi7Z2ws/7sOzSo2aImp7i
R120h/IQUmzIenqXUDD0nthHq4U/hN5DucTB6t7TpXVgt8WwMzZOaGYYCVg0j20m
pMXv4G3umkBSAqobaruSkNR+advhkepEdNL23DkarUNXVTaWOOCXyc0MUQsSOPMk
9yKLJsIRXYKz0p2mZpP4MSDdYOytGtpGXMMugpp4y0ItceDqL4MC3omwyqFEKcNV
F4KRMequaJ9qSEAO8SirlJO4hqNC+BXy0JjCtTDvs/NgYq0BSwrHaJrvdzIZki7Z
g78Skw3TWJsPY3CmS9MCiLIgQ9TuGav+JRUPeeu5B42OUzsv9dEkR+2jTie7CtJ9
VWHH9AYDzlO3vr+AvURAAwIUQS0E/CSGNi9m3/lnOL85nI8NGZ9Y7BZg30lRq60e
eWM0wCSKa+D6wUpqW5ygdPComj4NySeGcAeW06ialI2vjWeRbuqpWj8bMEI/mU70
LQP4AA068ojOjpJZCMXRLNdMGuGuW8A3wgqpqXHrsJ4Zn9q8cxBOx6i5ypdlOR9D
4sDAQaHQx0ZqlyesKwRnj2p7oTRh2xxtiRPrS8LbVSun6ytRcw57H6gXWUj6gEge
T1ZO9xltai+XL5+HhcoqTYH5JyASmWiGY/lh7bQrQGHN6v8mc+HW4je9lOBzMZlK
KcuN8SKokBgnVbX2BpgKK12fIg/CIg0Ju89Sq38/XU/0mFEjIXs8BE3mkBxpDmJh
ZI2IQIqU297OxV4P7AVW5OPN1RoyVhOL9LUxpQhhemFaNpw8QGzmmGgC/jbg+FhJ
5cf+cBugUDOR0xEkgJUIGBMajIF9W4CDOAyu8RsIbIoTg604VCMx58B5OT/XJO4I
Wq/6NDyPtNM7opm0fSN7/GmRilvN6wuMkvKGIF3sjaQTKRsrbS4KSgzwcFSn/h2p
jafRqAmRgh+rwiFJ76d9iw+hwz0+LwIEoVqf0Uvz+d/gmAPzDk+HaqQOlWFXcGUP
mcgdfdSDi5q8Hs+//l9NPDIuZ4kS4R4uQe8fxObRvASNa0P3YdNW0pcuPHMi7CKS
Xr60Z5AM7XAHywbhJWmJtaOBstPs2HgILacX0m/f3i1pPDPFiTRsncv/zOwcYKtB
5YcQiLDasytvLUMDEAhl4WHuGaDxgYZi/KJiKhWYZlVjYlcsBuBsSdAgpFAcaqfj
W4Rm8wsJt3K2RQT2LFkuEsob/TW/AX7IDisiKVrmgwhc9W0Z3hxU38GM4ct3bBPq
Q6aNXaP0nCJSiAGltVdrNFYtY4vu71v8J2kTt5Lpw3XOfxIEIjTee2W1XoL8qOla
s/+SulmfAIRr3Zqd6ebLZ+7UuV3QQE7bQ4vvR7USF6mQ/AXQE+D/wOzgxu6WKKaW
2f6PU1RCcxpUX5LgYBq9G5r4zKysQc0Ayermsv5HfgLi0nNF51oN91T4KwypwykG
9X8bVww0cUykPTRVUBNJnpCuCv3fpi3F2N/jDU8+Tk9IrNhnLE6YPC8Iq0Xt8wxK
3mhjHbFsFoJr3cC7n7XRevIsYm1atgtqgU8XSLDN/cM99mG/Lx19oY7+h+vVHRju
495TKZ4e/9u36djFAqhQmHxTfcap33cpw4iWVNiJ5L2x0D87BWS4MiTKCTymqqGy
tbtVof0hQLtnyZbyzYfjmM7tJsutK1KG0LKnD3kjzvvolNk77hHYSXIUmWozuUEm
mizTpQy+k3vj62gqagXbBCg+REsnBISGkJ8Q7Pic7E7/cQHj7Ib1COsgcWTs77DC
inmDEv/aEh5X0jAnkKC44iwyCNzZyVgW/3B8gytrhqEy0WT3YlGwkNrDlzVHw+O+
I3x/jbZoCty9vqJZ96dry3hB3TV14dnNT1ctgzZ9/cC1wkm101BRELm/AihEVrJP
HPjgneRYD/cTgN2u6sjGzyuE7KUnOZKO2/57Ad4y9RM/W7PbvlGTYZ+uhV3vetBX
vCQs/KThnAcTnLA5bFepuh6QEAkPOckixK1a1LrA8SRB0Us6FREhWiwdKbF5gO6v
oE3w+7dA5CQZPgxANmuZ6Akz050Lx3mD+DSBKWNx1CPe9KRhxw4iAQzgQD2Bq4nC
VoiTzP06I+8BxDr4r8pALjncvu5ouDO7j7LoDgC/JUP/cxKn7EpH49hk36gqwyHd
1KaqemiDe4ZVofI2DjR+Lwd3hLpDwBs+b1J5O1xzKVuwss9Qrr/mUJg8+YIn1Hum
WvCXmnPhYCVSvsp2Vt4VepDdNs3ty5/Rw4yb/ni4R1CEDpx3qXQXGO97FqWQYX8/
O1JaujxDQGP/4jcnq6U2PhZ3/AMmA/FD5H4h85djNup/hODIaMmgywvf5aKgf2SV
0vF1wSJikJLWR6V6q8Iy4P4PixZMTL/znNz8tEcZwyqN/QYl0UbMigtkW5zFEuHs
P97RTzztH2ugQzw1nIMhh5TISnqMupK7tNBXTS2CrwgbqwGU9AH8U6FDLpxkOpH5
6LZo+MOT7Hzw7B08EwwXBbaRCR61lKNCq7dCI8K3RGVGmVjL2ZwNm7J8chao4kHN
GhO1zkU1BlrMA2AAvwe+RGQ8Xt4rylq+pQoA+3r8RvfNwYM1yGMD7bXORhPC2xKQ
4y03OTxb04ADKl/w/cyY9cOLfsDo2erkSz9UuYwomB0AkFGHeOY7lhud60zIYVHs
eTe5lqJMtEm3umABdmyrrUEE2OY4tTYGJbZCkbx98aUxfTmXMsA2q60wLZ2Agamw
7XngFiNUQEI8+GIN35gQM051SSjqtF0ZQRhiu5VZUbHk5k90dMhC9m5hg97oIKj5
+dHTk+wMpsBnVqcqItcY1QlB8APciBRyPF6oJj128dItWzwqjP/N0FSpSWWAG/C+
LTLztSBIYfVesEt58KIq5fqjJPygaWpwcrQ1i1xdfwyBLaxiZyhiKTIy6GHx6fkv
Hb23WpxZBuapaugAw/jAsiXjm6RCT5R6/KhBIcyX35HZFnkXzzRIgm5/0l8bDt2p
wvfNUNTVn7mqq9TsEfVeegCEYFXAuVxlaCD9i071xsTknMliUPYTIYQcKr1A67WN
/0m/pONMiAHK1r1fhjcJWaqkYO1E2ZMnWvd0N2I/ug8P5dicgUq/aD2yqA49/awM
Gk72vYdZpSv5LsreLT1kXCJMJTt4TbLvBb0LQ1nC6K8a6NvwjPm1Z6ZXJNPc2VXq
EyXR8EeK7iQqCPTRguTUR0n6J8Vg2zdeJz8J/Z9sEjqH7SbFTj5YQGS8+nu6zt3d
a/vu0utLYUWILXIN6iRLgCBanStOU0cUDzPanL0aorsrdvcloc/MsnymSwTWQbe9
ueQJo43JwjwADxgwuiY7UYHUZIKl8CwF3OZdZYzOfeEFxDEY/5f9mXAA/lrD7zIf
dg++Al0udYAJdQCVqcBdsCIesKDdiJsPS+t09Sz1azf2+IhNM8qaMnhLFh7BXgb2
qr7WLGp6mRSENkZVA3tf4p6lKWIQoubuTHfoQnR6x1tNVw0l+n7s+YP3qw/OFBMD
Oj+37Kp4O6plCBOQ256/2X1Ae/Po96TsPTnZQX7yWtwN82kciN3U6Ai1Zcpv/o1/
Yf1+oqYVj3UGwLf/p6Kp330Xt7FwHyOcOc4IrvIrCfzr9bNBnX3lJNqjb6QIfVpp
Yg92MIAMHFpaH+c6PZQcUWaGcMbZw7cnhFJHpER4CvC74FtWpXgz8aMeN4vOBDV5
FwyHkf49GPm4yKcBP5GLnpxRKZFX1f6MCmZ8W+ptWncRINDSqmaOiWFcjqgpJqT1
5rCK0JWmRBxLuCGxphNhruNgsloi5n9MKx06zhyDHZNE94BYxJVoKQv35J7OwV8G
hkSK2Xxpa7g8IAR8X+yy3Eq2rfKR4D7L+q+Z3O/V88opyvfa4BYe+iJUD9YXuDJY
dg3/tneDmlnJpWIq/ldVsp3c6E63fbJ15sEKvmeXIQIhykP2Bg8eXIPe77cC4SkG
qtuaXL87auzydeO3QHRKdvgx2NAJsOqnicXAwgPvQ2O9a225+YczmMS5B7SmtQct
THw6aYPJoS0beDHUv5cMuVXyqy4xbfS3q5595f5xPXW794pM2a4Ru+LAK3uVvI5U
kWS+ZsBWJoSy1LZqKREu/fhuBCY+pSuPW8rxldk9rX23ccxe2vyydC+vbtXaTUoW
sibvCLAs7jRG8sJSwnrMpne6rV5HNI5x6LWKAcKEUPQjUTGOE16GGA9d9b4Zs4Wl
8+XqHi/bQQAwi3TPwbkA1eVmxYmVVW/XZmJsE6b+T7AufGtcot+Ra+LlFkBYtesd
2QkEyvIOkSoamn3QF+bM/fBoKI/5xPQi+OV7+ll9K88/TIahBrBFryWkzQ6gCwEl
DLD9ysUxAijmgNBvfyCoRk4vc4Ak1vlKCFm1B8P6oE0COa6eloF4IfXUiDrGk8Wg
ZlTh1AxZ6gbZSfDWi5ssFvEnyYCszDCh28SYEtY7zZxH56Quew7Oxx0wqswRctdd
hfO+96yIuh+k6YydMX0KQRvZmKOSbjFNQhRFqtNvsaVi/gjFinN7b6/S23ntVGZp
VAEn/Axpg8QpKbBPjcuXc63pgZFSLql0bIrHfbeJfer92kb17ES0kvPN6hHICNqN
RFiL5fXnGnZKV5qLC0wlu07jBsgdpBN2jhFUHkjQX4dXHrbsMXvaUApdDp1M3ZQ4
s4NjtnAxYMHyQc2gNn8g6mU/BLKXb8oa+r7NxIJPSYneNPDAENpY3UBPqmvvw9Oo
A8MyE3XDRDJG3I9zWA20f/Ux0Mfa471idNks/OVjT1qCMCeR1nOnaYp1HaHXoyJB
7uET6ezMx27sRLh3qvYeM840exndo/9ez1l5W2KZBdMv6A9zrQ9DjJms0sici2EE
T0baI4bG1sqBx74AT8VmfB32WcJ1NhDqhzCg4vch22UscMfE/w8R2RzW5gtq/nD/
TnKUhtsPyBRTZTuGKye7m44Kfjj4Yy7cEcY2MycJPgXIgUkE5WOPYmWSsbJLJn6n
MSRX1mNW9IEtAUxNXM9Km2dplYD11kUiJhnW41ipO4jn4nO0xhffpuDEZjpppTjH
2b95ciceaR0Cm3Q9ykKlf0j/pvQk6FZOydXNdGovse44UKcf23cOScjji5sS7qcv
BvdO+TWgRPDHi5s/+NKObmG05L5bXmtpAckjwTXQWQKMX8+RJ+17rrudifmpADpd
np+faA3eBJx8l2e+rX8s7DrzS7A2kRJsgreuFmsZhjDqPeE56BEgVIlo4tSxqVI6
BHfjr5qdVnvldQ7N7U8liiJ3l7jJYdK2zD+rjvAraRsU1XupZ5Bb1j1S0TQ+5hRv
Rcw9/WyDgnuEo9k826O4lo730mKwEuIHyJ6TgqKVvezDYmRUyF6qllW3QC8cFGWm
nnlTuQ8EUZIrf0hhOZwBL2PaqAnC/SkK/Z1s/jKkd8dUf7JGszIJJmn6VNQiSfgZ
GQmTB7OwHiTTRLqCIbij8/bHIXXxY9X1jgHrqvFGhL36Un2jhb4OJueIgE9U9JTJ
NRPacP8NY6O12ZskGUcq/TfpVVOogSnuDjIAtVFx0f3FDJiNx0X33UstQcMmC+pS
ON0pDWCoiV/ObhCT/LQlkVJehF/A5sLDEAP0hqU9VElYNgt1X6xduR97wEptW+En
VHXwyuMcmnWz9mcgO9/oKGEZMkChzSajYySgPXgbCPNoXrEQ2mu+a73WUeCQ61Mt
9nuutjfK0IUHq0gmu5CyG4pySuQCGB491Xj9alarb103v1y2w/9tog4EuzTa1Yio
mWSPysdYSO1XORIs2EVWRrcLvz+ppH6nCo2wxyq/FuKSXwQ9i1wADyt3ks0FA7xP
nbGaYPha8UbyWJJeo0ilyOujRCeSHTfupNsRTdbwJ2cSV4xsenKAqRoD07bLRYsG
nUADVqQc+MNv19Dt1gVejKw85pUTbbyQOZgfEgSECeCpY/5AeXd3iNZyCgvq+dUr
BoY0qR1mSPtfSEcZ2Vv8iRLxuz13jbvWNafmibgku5lrPTBchkDAYOIsWc6/lIUn
9xMjewudu7dcf2tTVYoHgNH3XioM3aptukoF24leCM4EwwcjzsTkzXCRtsSKX+AV
S0twWseifm2qTgx5HyUrf0VnVcnL1ByOS8XTZaqNW8hf0aMWY9T40nQ2MSmiN4ac
RDCx4PicijS7EWVP7NidAATptobPMRcdvSAOwExbhWG+lGwEG1GSiEzeYCPqqhVT
athDTf5G77tplKpY4QUo0yPhWs24UgXOphJ1v/0qhdYAk5RITqqjyZlNb3tjmOKT
7pjJAbX2d+7dJV/QQx+2FiDgcjpRVZSvKslNU6EViJWDTQwPyyIYymKgnMRdThGH
+9htuoZzeo0+92XmSvIgOH/K+jesuBHJLVXSgKXVbWHCkOsffgzI1vPO2sDHLtmJ
9dBR/cjcubhTVRSFSDqpGewaO9aq9W2ZIDWH9GCZgqZdhG8aEQRJOxRum/Cewq4F
HpCmW85diu7j0hFIz5G+fV28t8rd/fBDn8MBtR/o05Al4/4JVOOAQ5b8ceDcIUD8
NO8ob3mCzpWIQeC/SXzz6gAnst6UPhr0vEhCVvTHHkifONGY7E60Ds4jX0ueOpAs
c9z7Gflfs/50W5QfGc6hKwBKQPmDERBSFb7F5VIaf2+AgtKAz+wXE+Ba/22vDtg5
v9zFrB1w0XDO3waChtdxZFG31wDMgwibNBLYBT7YbGEM+Rb3DGaEh5Kv1/a93uEz
qG9we9wo5mdLmWrA5fT+05S14AJ6jbNCdw/+prPyAtx8at/IHGuUGyLuH3fnVAPO
X1uUNe/RL9gfNO9W1kteUe/+bNwTTwzfU1Dx7y9GpO4FQszbK00KXNFa9w/IntqU
dapZvbue9ykAg5F1cV+1vPTjfJov6pNtrmLEjm1OlS+5uoX8y5OFjcA9KESDURVn
2e1Dfdr9fofgPsFZuOkcPL3P1xpJyuUjch06EKTCjmnSA+LmRydLqfzMGoqrb40E
UuRA+W+aaPLAnHPEhHygt/9RsfOUJYBMkEdcFRT/tciJr5sZZ82qQ9IUpaj5Dm+B
GxomMPdIz+kPWNMXAkcnpRce4k6fs6X6ory2KuhAhBqPJ+u95gdRChAdY8hXlAjj
+TB4lUU+SmtxkPG8FnpLCwT3fsbDPykDmenxeDnQOj3eiaH8ZosJRoRFalTnHW2B
LaLJuDaEJB9WMXMS1Z6nc1xLREH+T0pCUAV84nh/UpWVoKxbhaUhXSNA3I2rTl9x
iQXK7qK4yfR8pWK1dYSRveRf4PeubZQMv+AlVFfFgk0+5oDe3fKlhRzz/sEJ4w2V
PlTJYoHkvCI2nFxG+KUjwlzWwgFsZFluU4HS8Zm/9yY3wXT+slYk2B+ujp7NXyWS
pvejV+b1RK7fgw1tMr9fltxun7P62G60Gqs4A3prGejSDBM9ck9oZM34zbQJi7AU
ETpx+xjksxAoGDE2PiPzjyRThEKGpjhJuzo7aY/4JakhZpKqSd3Qu5+BIJrmLIuZ
eSX8/DQCqMwMl/nHGeCWPA8MhDWNY6HkwnafMCwni5pjnVfZL0Q34YFiyWY4GDNN
ziiCoyMNH1U7HdQ3r3G14kWbOqIDdVYLWelEdBbIwCiWeE08r3cYq6JJAY1h0R25
jb/NkO2Tn4IK6j2mm8RC4w/K6GTyxgijr1LNvyIUCmKKD090qaCA5l7m1XwvrWzN
MQZSQs1JL0SilLx5Dzma7opQOFnKNk9GQz9rz8X2/MbH0h1muDMGyjjmWUpH4CU/
`protect end_protected
