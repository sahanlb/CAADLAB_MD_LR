-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
7rO7MUzVZYSBKWMv/zS5EL0n/L7krmFLmapgFdENXVTzUCTrriYt2Y/seSehpcbb
56w+L+e5R48xnylzN0WBl5j7lWUrKvYgcyZfzjOx4rcKkcyd2qTfv0hxzFVNwiec
6HeGJnuDmAMV5pLTokqQ21qyGIzS8LA9hZ8eXfyGXXCQev1D2Jg9VA==
--pragma protect end_key_block
--pragma protect digest_block
8F7W37q+7iCNUMjeqGk4BNARUUQ=
--pragma protect end_digest_block
--pragma protect data_block
/bq5QKPY7modyrOGApCvLO/mqhOVqsg+rLknoYl/J+LySV0YzRNnGcSLbzmMZqUo
yMjfHYlgE0ttdxVyRRrE2CidE7sVr44sQtGKmtCAnOpYxq7uBH98wChlOqyZApY3
gOta5RvSQkDo/hlQvchfjsQDtFmJ6nKkMDrCkOK2eVnUcgOByqXp9wKe1Wp8r7zG
sbrTDfMnSXxeN2tsDYs4NBZbcghSUxIar6yYEQWkZ+ozYsjK+zm0vhEX1HJXgiSS
xN7xHoLvVWUFbGi5azKoP/MJ98lG8aDry97YAIPuZvnqAcMO9aFRAmWpSdHKUg7p
pB91ny21CCD5CeCX9MvvJrysrLRjtvqiolbXo9ZxM7SLBuoNMchkId8P8KMWPxX/
K3dotnO9wHBV4jcA7AjCahPD7o3a25S/KmR33aWVbRpRLDE+3Ps4m0gzB/R1i9Vd
hql6FiGOGnEKt8v67Y98XKr0ctIfYudG5e1kifwsFKkZXdnOMfoVaeNKAqfo7rK7
xeT2jIOWkXY0Kg8sOcsXeRZc468rtrGRBltCVzToBeI+0QtU413EJppVuxpm+Z2f
5gQuhiYVQtlPycRjUG16vz19/Y2jreZBkut+GQOVkygcZEm4UfzXcMzTFjS7a/hu
g6xf5vFjMIdEh1USCwmyjl84uxGN67SqcncCKhvIFo5d3YwCQhLEOKgB89smdvrW
cik0+LrSPtjr8tECasqvuYF8BmLV/Rsp9/yEt9IRnNdkxNwo7tQdzsYW3qdC0nip
5JHwy1KkRp9l2wAtX+dwg7dYDluBUORulVSMxS7roRQhoilloH+wG6vAirmqYR4D
RCRVRVggqoxcNdLyBLGILBbiDdAELXD3+kSz599b0SZa74iJVEgHEi/vyzNeuwnF
ShlVUbASetpuEr9uSV6Zk+Rk8On2SHQGkRQk7wnxqKyOQHYwkel0sKw8HYELT397
v1iIU+zObv0SbGaOyTaHkr2YeOoDpIscjbUgMWpQzN7WMDu37si73piLOSJBxGmn
gHsCKM7DSIPeMqtrpVijJzzTAYv1MrbRGLjIRglN9cMKr8A5DMu+fTr3JmL6TVEa
Q+sKZ6OQWytehG/TgAD3dRQ2ZPxzi2wL66EQVFWqMRCartAxqzF2+JAM43XNthNy
sKFOGDMoVlMCov6e4MBjAX8TUyf3xHqUeU63ySJmzslcWWNMDzjBKdHioGhQjf//
Ii/szXGnWXTC6KhWYG4o7AxCnkXr+4c42kFHnHqoK0+yyxuYssLZwzbCslJ1BhC5
kDvEv8S9rLAAHnfOkuSbEQgoZ6G/cvsNAll4UtLfkEl0n+eVdmKpgi9Wc/V9MJK1
jzOzegbm+o+tdlDCnySmUwAnk1eZauS4Hyk+E/H1D0dYBlObiIHqmqJZLi+zuLD8
0NItsZZ0C+NlqJYi3tj5b/9S+AYK8hXPHYQRjxaejn2QgHY8nYN71BiOht2RI8oh
+J4BP7AG85mZnlm9eJrFpHpvUD8tUJMiR1+m1ICy4tqzII4abDCbvLXp5OuMHbKE
Xcv4rZiExODzMBjpwm5Ajpn1izBG3oSFJVoMZ5DewfXmp+BkWTvZKZ0npIPKTAlH
TI9VTPl6uNBllYO6ASPHwPx3vBFUD3Or4UwRn4885MvkWM8YucTY24d4SumnJlu9
IlNMKdMUNPf9dTj/GedYvxZ5EdwuVr2ybiAgZWlYXQd0XQ0A8/T2heNUlAprwTVG
7amHKawDws3KgJptggZZvKqNVzJqcRHK0FV/jUPZmc6vk3UDb0CqesejnxB5U83W
ZVFnDw6N+M9TFRthWKBYWpWf6vZuKyQcnNq+a6otEo4QxYyHlLGnG0eNeaZ4/LBN
ADIoCha86feR58lAXVoEc1k+0if+UAOeXQCRYCn53UxvxOhUsfjhs3+h7utRD+ge
zai+2Ji/9eaBcZSRsJdVmy8KJTUTwVvwQ308RNm0OCYMrQVbUSs7KiiCYtARZRSa
zMU//zWNOV4df8xKlDu0ZlrSmYOztMfwihnqYsorbvjRanfc0LMEMtAuwiimTh5d
cHfKFyXdgDnP2wQ5+/jCv8wFcZvHHgOl1YYtrdhQnzHpa96OyUyJhordJA3jWeR+
OW3sxvzHTOaMAHQlc/HQG1n0DWeIPbJ8Ouri+akC9NefcHKxYzImjUfTKa7oTa50
qSvfhuQdaz3leE0OSifxKx0Zf8gdTG441haWiSkcqjjqKsp8DOL9LNCAObN4Spyb
zkXGPD6UFYaz1TcnnF5fCyCU5bSS/umnn+9bPdFg7Nus76OeIMpP/IIweL3AoBPC
XF2iwrZBw4WcaPByOPanOvKwySteiRqm0sYJBn0WvAgqw1n5aU7zKCCDVZcY4Vsc
WOA8apm1uhJ/J6xtJPZdovU7tKK+yqyscw3PVf+kWwNAAkwuQBhgeT0K+XBfL7MD
DmOS70TTLkPxZy80SVeLdBoEnKFgHL++Z6Int7CNb333llbSIPHH34lfeFB0X0t2
DMRrqpdsELpZO65EHTILoix5KKU1iFJ5/1V52nAU3tp5MRt98HxUbDrbii0SBjkM
eDKI34dL1lIqwWuzAexfqYRi3/4+JDez/O0Qxna1AqxJSERQUu5EvfnTT477RSTL
cwJ56XgpJKzFnDyMlhLm/tj7jiNeJ7km4ROSyLeGKPirto7x03+nhqkjG9T/Cgm3
d6BRp8LFkWfwqfqxAE4cZC//MI3/6hGbCSNs0vK/+J61rv9voly5AMpg52oopY1e
BQYVS2BxL8TLqHRW5t4W7p7PGoik1Q+8OqJhYfLhucGXcN81qBHPA1s4mDzUxFbS
NNpusuMJSuJe1DDwU5x1Z1btqx133GDHLUZVVRGCb5KXHwXpMl9sSh/k07G/tJFZ
JdXQA1XHGiOl917QWeddH0BZxb5SUHxDNorXAheSE53s9djwAyKko6c03fWes/t3
gHLdf7dKOTf4mJv88x8t0+04QmwTfX6HbOvvP/uoDVz8yUJbp4r4d6v8reDrTZbP
EhOI91msXdWfVPSYClNjSJLNFffAPDUSr/KYekl2N1PjOx7TIUSk6ip9N7LwiV2q
C03fFs+IlJPLMMxlTNQdYp6PxN2z1U+hx7HvzVwKrwMVK5fqnwWzniMBC55s8w/J
vAEsDEBMfOmm80/4XzOeN+rgzIIXshT4JkcIHtTgrIHzAbMwDzmxuRwf8V5poBa+
+VhtUc1xbOqbImwmYbYVQJgQzxSenkqMAMDgdjlQIzx+MXhUJsRvoM/4l2Qc9ARS
cFqSQTDZVHbIkbGO24QIrLRpnzqtWwtcoqNKDvjBOK0JQGqMfDSIO1LGAQI6UhVI
hCFe6VNw7CZnGjPiCRsWGXwaJcfikMNWVmvxUqYlWouEIKUZt2VZZ0NwEQ4cou4e
nUVIeEOJWf4J1Em7bm1dITmUQiNphYQKhbuUyJhoxrGh8EKpA7MY9ZgodRMyApfW
zIYy3BsjMliVHXAazc6qPbTUFRbp3PNghu9fZp03QSCg/A1ULBnQ04PLDelc/uld
j8nUfHSt4/NNgwcKyCwAHh/58JfxJ5jqo/ylarhxvG44t2gFCt1iwurs2PvWoqOf
QzDE4/SjfVDYqtaQ3r0jpe0/vhKkhWCIXqZUEM7Te/1oh8C77YQFT8PUxv9GkgzG
lLtCjjsiVb6VqNcOY0u6cD4mKWhUX7MpVc+H75vCrwqqi30DehVxU1TPpHVI8FVR
XR3p+uTO/6Z3QnBJzv1yPOFiuCCPos15pfjBC8S22lfW+MDVG9b57pFPf/EVdDZW
c/aXE8+XwWlCxDXr+ORTo6NMpyCZYkkxBFeC1yCOHS74FzPd3g2v6ahKXjOiTcmU
YU9ygCBPSWVf0DCisyzCRI9bPC2A/HGWICXjw9kYSSP6t7csRDTgguC04A3No9jw
VaRxCGan6t0b0ZI6zqx1Q3Bt7/dTTrljmt1mwpnB/G75LahK395l/H0lWteWow5f
ZZxVGiDpujQEIod9V1cSJ5vFpxz5RHUNp0VBy9HFltFkFFk/aOmMcbijTjYjUDuH
A6zE3ShdfJ582i9uc0LK7UA1zrUKERRB/m2q/mraWqzne8NLCWajFlmFWicn9uR8
9g6dOYnUGS9YFOOUaSMMPoLIdEsIdTnzoXkcpeReaNp8o0CYzGhGpq95ip9xKmkX
iwcXDMRgPYo1EvwNpnsWQgGXes4SUKhFaVT+vFbIynQfZPLttVe4d+GN1DDnHII0
kzuWr0Yegp6B00YES3X+wvyRGSjaM7yG+nqvt5nHBCbZAkSS9z5BFvykK3ZRulXH
hVkPgNwYtyWcM7yFOawC+mTzOt2wIVFH0UXa4wxrv72m9Cukwnc7t7YAGSEJQEoN
XslYRm7QAki01aghHDygtS1b/WhcumtQ3QHZDCkXl8RC3ts6F0P+e/xawyXgMOMl
dKBJgvdG1kb9Hpb/0ArL2kxaV3CcA28WWVTITZ/hF1qfF7eR99h4dRf2avyAjSE6
kQEC1X0Pk1Ss9bFUW+EOuYQ4L9WWBalvKzp2lRpBbJ2wv/rETxZyJE7YHrbmBzmI
MOgmWcuW4RoZ7riyePKSThrz1A+sEA2EictwQZ4Oa/+Z21GTJzTyC3zuZFYtc6fu
L4wKf8g1Jhc581ivZ0fwyFbsu0N963LHbqcB5H30aiCMpHsa2oVTTEzpakMw/oXQ
pZeymLiEyJ1WsrT+Lh/S729pDbCKgDFM+R/8kBXQ1Vd1F9M3CJdBWTKFGA7U+IMa
zxx9sSS/lt1uYcJEekkb2xtqmXComWDDOVFKQ8V4STQmMbGjzzIyxE5NBmtvh9y7
q3hoJQzAFKxg0EzyLcenJv0fMM4Ry01ORabNJ8oMlB189LNf9/3sJVqCbmoSiYc3
6Di1PY1StIaogGzT5O+/gtbKYsTAMf+9pU56QFo55bPBPoP7sheChksN2xMzqHA1
Tqni4UTrHpIvcu6JCnOYMZI8Jqu4YGjfafJDI7DotIYAJXgNmWD1IETWYQDfnsEJ
sJd5GOFVcW+QBkmBj4W0+P/4R5P2WsYqw2vqLipMpvBQ/QRra6HmxWkSANUJY0Bk
k4JA91ZIqmaOq9tc9y7TxwIxpJLly1PzHUqkixsCRwbuxY8UHgyqx8SP/hiBg6pA
uuFEDuFsRylhAf7Dz2cQN6YSdUE0yy0q9z4AImBC8DJjVJRu0HQLlePEoGX6rvGt
FryMxqEOx2l6rOlVUtFL6HCnLxH6cKkd+4VM/zPe+6oNwlZvxB/pOrVst1UI9XPX
MuqdMVM8dXRKwDYAQgYrazavuZdliPI9sOTWpn7PH1tq1LKQcbDCUgqs2YqblLNp
UTcou1E7m8PBQbuPv74iBeSJ6rIiDc0YpWTuYm444GUrZuGycPgKO9fNeshH3H4B
uBeaP/AMnhu6ciaTjRpLSh1eBDxdko9wcx7WESmxQDq63Rz5Pe+nZr3Wdd8Gx4x6
FSZNKsNTVLdsh9zcXBpwAl44diZJ89beErdp4dqiUrxfGtunIwzkrNpDKPVE4hla
qs5q5xr0Jxe+FeEJl+JCs5Ve60AGV9JrPIS0fjs8TGJwNgLr5FNWd9pjTVeP2Cg6
8Owpg12yH2dofhgh2qS5ArFBRmJQlghKsyaNsPIeCcoo6K77dHos6Q9x3Yf6I0/x
9qFh3H9rZesIMtrjr/9i66jvFeMyPRpOIft86PtFyYW4UZUYWBRCG6JYvYvPH8mQ
MzEPtxSmjCTNdJQFzBfE6yzTCYBf/qy39aMuIzCibkL8jsGll4HeWGXJfn+PoGjk
XZG1YdNWJl/cOtvpuzDa385HkfSEeMFuVikJLYApF+M/6IYA0to1f24KO2N/7z5K
+fHEqqCMVkS4aXRbeN7rytSTObZZetddS0lvFBHuRTiHDOqIIlxYOQM8hWeON9Hd
8NPrziYL1sTkMOntDFOdltv5EC94d4JzjC0JHrQtbdqJuzjm+XrjNXosDabW6e3U
9l7Wlw/8vIQQhLDNZrKs1VVYRD3Nz6S4IjlBeLzlKLD93rloHSn/T4A6aTYj4x1+
pr5pG+ZaHuW/+yilUZyt1UPWu5C4TXtg4E4E2/UdeV7dZIci2tIcMfxnIzOyzZQO
1djXNh0EM3OSUUccKWlVy/8jdRzAZszLcA3PrzRX8KiOJ2Ea/ztlVI/v1T3fPYvd
htJCqhoE4Lh+Yzeq87DQUGbjF5IdSacpeCVV1/6Gp0DnpG3lpIkg1IiNKrJNAxye
emPr5AsbpXLvUUmp6u9nsePb9N2VvCdAG7hu/pTY3YrVS49nYQrx/yqPjEQuSwe5
2X2lEHDT8G6iut+RfDqvAkYoxwF5sqSzAm7kAfBBToSZiB5hWUa1qlUDpEXXzZcu
1YfQb64Tr/TtNNO5L3FvCkdkw+EK7f8U1Y2R+byNheQ4kblP3aw0j4pjvBtb4a1k
k22M37KJlzYCn4yEVSmS0Ny/z/fClQ24lBB0Lnl3zyEoTGCTvnhMzrVLhNd664Yh
Vmi50dLahUxlrqtHV0MUAe1EIKgf5M5WiGtTiox8bQl+5cr0eH2UPS514If8zSrn
wNgQtcr+N1VNff7lk07Xn1J66ckG+2hkJ5XdRvJMHA0eqd45iYb7UevyNNeyxt0U
fO78mxUv/gC4UqMlAW2h2AiG7Kd0h88PBnHnnkQ3Xvic1gelC5Cr7nA/y5Sjkyjc
ljqXLv5dJWw3G+VQi1HUqfXkwghCNPK9Mra7nNGplLny2aZvOcDW7L2aNT5vK6yC
QA2uG8ECcSTr7rRgnIuN3AJvlGXWi4sKXDOqY9S2YooP+k3PmXczXgOIf5NgJd8G
m2fvDBq7hPJqKWq2oP6n3trNTPyq2L1iYtLTRg1Q1/kmkwAyBtjiiuWg7heRZ1Av
tiIAefowNKwGnlbvQPTpyjMpRzdZwUw+9hjdPf7NG1LgNF+/vRka96cCxhBWaURN
Vg8Vbsi/i+8Vd+piRhsZ41in1g/DiQKJe48occzwkE5oe2J4HXdyNaaf+5d9roMV
t8BVsPAnjXMIk2FhTW7JRky5SGwdyMFtyWIZMOg3TFhh6WbaFvfAQ33uXx6dV6ox
3i+wEjgNdo5dIFLe2X9v+y0++4o9wBoa9Y4OS4LP3kurFZ4+G7cBWxAZnW6Wa+OO
H/LiWko4Nzrb5z8yuBCnIO6kSTcIFQH4AO4lRdtircLn+5GLbnw9RTn97XCOEQUV
BNMWbXWWC5nEF9QbO0lFxB0Vbp6qVVvS2xx/L3MXm0RU8tLBQL6AsLQk9ojsnAwW
DO4N1uGbBuHWXZLhwRZsWOD2XlGQ+8rzcM1Sg5HTV+dute7GcRHvY9biTt2IST+F
4ve6QqtYKRUsScXMr4qdr121D4Caq9k9X3l+pqxUr9DGSiINfV1PGeMfNJj+OuHb
3yq1ctwv8wVaM1d/P0d12GJfRzq68jw/RKDxhYsQnsQddmCcOD5TKBcXYNF+0XR8
3h4EnD2PzKPGWbr7eVfRT5gVHjw8FZN6zhyJGcea84AxG+kiUPXZVfoYf0jk5X02
ukeBNjaewIT/4iemfckCbpA7OjWae/S1EUzylHhC6PYWLuIE0+fAP24pCr6rEkSY
ClvOsU5A/o7lt9PGixusIxoS7Le5ewnUaEG0hWAzBF6iKSbFV3sIY8/31PlfIIDp
Qi4Ldk5Jp4NuBOIjpOnwe+Td2zmfzi86N04pVF03q8+igvT7Bi9KjqVJvLI5iOxm
sRBxhX4783zkw9W4s++7l5Jxd6h3164D+JmsR8P6/t50gx+S2Th15FthCWNQHdzd
oLv8NioQHTD3GASMtFXSPa/Y+SKgANdY94c1kC5Wb8p+YMT1yf4yWr6sNEPofrih
/AWzH5U5rWqof8eosHA1K2zNe3hokSaajTdkc3whiXyrRkIRkZgjXn3sreARUV+q
rJ3CVdOefaOu1ygff7olYCqUNLXjWETH/mRhPQi4rX4=
--pragma protect end_data_block
--pragma protect digest_block
4Xoli5WDf5K1eu089CNGWKYp8QE=
--pragma protect end_digest_block
--pragma protect end_protected
