-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
AoUadeRmjzzBSl9wkJ7oJVANmskasxWNm7HlgMxvkQn9V0ux27tT3+y7LqAMYS1y
V3GKK+F29lyH9yAVpKHx4Qf47wclDAE1oynE5GU/jtWeXGK7JX/NaE3ZrIlrmybY
1kDXTCRBGo1oB7f5YnfCmXfsQCSkfJfyHEEBYm7oG18=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8816)

`protect DATA_BLOCK
pbZSi0g/o9KibfXkU0zurIAfK8tskJ3j2gUZ1vX6RPu+MpvaM0l9Sx4Dkcv6kFt1
v+VGub9c6qVmxjRR3eyUfmp+PwLY2CEkogXgS/4l4OeDwmVBBGbZ3b1byNvaU1tJ
IEsgyQyTjw4BkBAmt+EUZNAlg17t9ktopd8Jzz83WnIQnfG6oaOLdFdJKLTj60wm
0zhfwc/dP9IyYd2RJi1oZy7Eal6As2FmRezxxLSYhu72cafkPtDX08bEdwYCG3F7
i0E+Hsz+DOjSlIxZkowz6hdpMR/zy/irIeu/EXm+Eb0WqpH6GqD53eBU5mOqFl9G
4y2VJqOpiu9PSDZ/cMM/ribfT3dIMgQllIySXYesxb2AS7H1OqYsHwcyMvAAljHg
3BmTl6CzqiBU9ee6LJt7SpaR6SNhHoEDR5PWdepXNnqAsm1Ej2HGz20R8P3bS1dZ
aOzXB7jr7bJ4UqXNHKrzdUP0VoutNCH4eB8iisfHLFCAtf0k2WcCBFmGv91yJ/iS
0Ot77v3Yuf//D33uNcF4Uk/7ae3VFmjKFXnp3SGKieVCAU/v96sobQuow79nQY80
BKbhhcVec2Z6qyB2UDlIrRj9mihjR0Yi4m18vOwZ0QKDr6RWuss+VHaRKVluhVUs
diaCiNelkX4epAtdqygeoaozQtCDNuSQVY6nWTqOfI14lo0bZExJU2ZaO22CF1qk
RM0cwm0NgVtVt5xE2q4l3vmk/gmwLtQcx1gTLyaIvntUkVa/gWn1ujz2Fs1/stK9
knUBR4PV1JFsNlcmE9dbSQ3fesGvs9M6GJPcjS2ZiuvR7IVixYAYAbJPtLFa33do
pnNYRC+F9MHmIT+6Bx5noJaomvVBODqq7IHsO+lieUwyvvBkua59jVxBS2DTfqqS
E33tgOZ/jKjKhWAeN09Vwva9vZn/sQf+x/PxbMB2A3jhw8gROVhrN5CyTAJaUNGn
SL0IwuHWJDKlV94TgvY1ROCxRYBEuPjkZu2yXL+rjGG2L3rOG7CJK7K8Ibr3pYoY
IVprQAS1fab41Dg2iPStSCQ/fWZIDQLtBNR/Sok+k7baIlLP24fLCdfVEgYSGBUi
Yvxn2elwVgGYHNlaz5Dyy6U6zTgmzTZF9TLROdD1QXEJ2gnG+GJfCV4Ij2ckG+yZ
jqN7Jj+z0Yv8ZUd+ryVIF7LwNWhuKybtTN3i+zKJWOtyW8O9+KuHyv/PnWkPe/3l
aDh/8Az6UTL1VAMOlO/U7VPVP6XR6j2986Ii3P2WTMGd3IAu9plIlTQyqjZ/DTd1
mK4vxhuXSa3SjcEOY7GKf/j0QqS4Y+n7enM4/OcqyisQIMDA92zvpD05DZ+WzSGr
7P6coI49ws/4fUKepcM7EmH5VIj6joj3kOKI5+4qMiDTYjRYmqRED0UMgIUOTLdo
JWpoAqAVbiMar/cfW9c7rn4EAZ2S5iypkMXrt7Ri2ESRd9NKKNuZ6eguTm7l7LLs
SR1t4/1+lJKkdd34lZS16v3RlfXRcziTITLz1B9VuYGe0TSjHrfuskHVH7ZgrvPm
GmnTKz8K9GXor8l/RBTXJNZuatIYV2LGc+EJTHpq4bCH3Eg1kc32drO/iFqE6aRl
w8OpHOKc7CM8Lkk8TycAbnZ1kgNbYlSwnW/5UwsKxxshGec2XyCIge7ylRh4+K7n
GhSFxv1n6QSlx5h4KSg4l1pCYwKYM2adV0RfR9lKyQYRv1grZJcbFBNzRihHE8a8
XHPzJdEVMpqd+VVSWEaQyxjkYSn1MQtjs2qRIUUyYze3N2E+0s5r74VAHAZ6u3Gg
cRar4hwn7Eub3Ssugqq8NHhv3fED1PbdJVcdjaYA60sdmbNHTbnlsCARGSu++12V
F8+VGOqNQkU3vOJD8kir0n0H1sXjQdAmuJKlSO/mH+iDOxjy5AKvHBVL3WKpWsav
jIQGRBvS487vo6UkvT2c+vggR7zx7OBcUn0gPwKTdD0zdtteki5O7UfMzcDFgMnv
U3KX5brLONztMRm/8poMfsgmDST7JXh1Enk0kF2j1IEq9dxPeKJZOKoswUG+tWF2
B4iq+UkYkVEvi2eYNLaj/UgPk9AoS+wpWMEDug7k/FazTpyyMTBMDZP1VdKw46Cl
NCxM08bzkdf3guQsrqLzpig7HGPgN2o3bGquFPZVZWw5sTPrVAH6kONWwaH23l38
sd4ZJLI5zeMFd2hX6g3IpHza/7gQxrHGcDgabbFjryM3Swct9N/bAdrx8Nci4YPz
RyBoVw0HFcoa3VTYrsrfjKx35KsSYhDHPgoEGKbys1BK8nAdsiveiG1IzlFh/6zy
j8espKnLd4o9Shz744NjOEETWQkm/Lc90/3o+deG9WHXCk13PKZ2bY1Cq4iQnum+
2BZt1DPxtn2N/zZM6LIBsf3xFgPLk+1B1zJlBFQ+1aPz7MnkOiZTEYKJ/gOkA3Zn
ja9i7tCtL51OZvFY9RcKs7w4oCGiNhDnu6Ltzo/wxU+Svn/C2lpNcP688OpgFMHd
t+5bKc5C1M8TPldmy3W6lP5nglhqHBE6yyCI47LZtVKZ1NF84h1uWfDoeiykYwJ0
emJv4Uz7+yHTn799Ixb78fZjFyQKgLY8lcXMukRBTXZByqXGRNFSdUAauUOoP0Jk
wUrbpm7HBR/tWlpw3MGYYGVx5AihVzIuJ84FDv0ag1zt3mcG0pWbdlzqTQKY9hQa
XYFo6HAnRkOa9eAllTrLcv8oKGHPcZ990WfjscB0taXpGErSLKewMIRnpdBVWdbH
RENtG6ZQTo6RzWmusF4frsO3J67DWMaR9nyGq18+P1jXQ2ckfmC/f3YjN3u3UgR7
O1bps9YMPYMipZGNyPxWfVVwXwosc+8akBvxCuuHemFs6hp0jKK7XPQw6SLPRmGU
/ylvEYnjFDwKEk7Ms+U5znxQGqZKBnfjuOM4j88uq6zPvtNWvu6hRPhDT+3kUmpl
u0mM5NMxK6qR8tVOfzs1fg9hEI9WRgHVcXBnxG6oR3zjNXavSz85u9YbxYYY3t0v
hXCl6AqAXA92VGG73pDyYzW/jELtRX4ilkmYMZWeGaWy0YV4zIk5Uw6HTQrlDCmQ
9Z+K8arrD7wU3tWe0MG16AcbRdvDooUSFZWEtm2DEsqP+n6p7o8Z42FX6h1oukV3
Ltmcd29y7/JJKi5WBCRrVcE+N0gVsUNU/MqThwzj6ItdfHa19RNSJ7ZsoWSorrvf
6izFeu+ihj5QpPNKp18kjXTArRENWI0S+KqF9bouo84W25+Z8PqjAjOpPuzWB3Oc
1fbTwxnIgnXYZOXxpM1tez66athTni5S6qzllETN3+wjTKMy/jLkJJRi49DoDkOH
t8STkuls3d38N0PgM6dbiQkIaDBHZihjyG4bKh4BjjKrCpOItIhpkiAuvMZaBCDr
sgMrES4oG/IKhwIgwCImFtd67Dw+nFWGzaaH+8amJt0/hLqfD4Avs42lpg5iygBE
2+7Ng0g6/A67A6VZhpyUyAzuQk2BJ/u5epNIhhG74c5ljYXnr2frKByJtIx/GYs2
PyknJlP0JxlPsqcx7F+k/PGbCzhdVZnweKjfol6S+8WFUNvunbyRyX4BY7YQig/C
dDqZtHVj7pJV0e1fBLiA5tt4HuBMoWC5zLT0O5xnqIG3XGa+JJHEFnWR2q+RsYb6
7A52YitwPG3KLeii399HQHNmcz3cLr9rabMMKr+6X4h+S4GldKJQkc2Zm4tls0iY
SJzXvlX8P660tVhobwiG1WLln9QXdyAEh71GKhG0Pm0Pqjw0hIpEHHUYo1h7AIKh
dS3NLmy6+UDXsqCLw79bKD5xVqa7NdH1WVP+f2G7PID8TSXR4RQ+fubwS14BcM/e
/EPxPMBNKiv0T3UE3N/KFaz+gA3yyZgS9Qq7O0o5Tp5T7LwUJCQXYBwWU3unpBAl
LAR1bOkc3wZcjmtYbiNo/sAh9EsQiLOFsKHKBxXewVMSTgUmpyY4xoHG0HOFwxVC
H2P1fmJa8jb0dIl5o9hl1p2sbU74+dsd8RawzTsFO61dqIOxfwJSKB57rj2R+4W0
II5Op5vz1nSVigwKQdv5ppRosoi7AD4WHGK+6tBsVhqC+YJNrCKIQWZgP1jHEC6U
7X0DdV6NXm0ul5GX7jX8NsEoxW/5xYkllMnBh/mC+Unrzs/qIwy3t1AkMDHTE3xu
l+vqpYt7JGsq5VNbE1lDhkxkPioiNR8rUF1oNYAoqRTipdiebiLX2qTVSCmukKSo
mYBkFDUDH2s1vyKq9JaaqCn+BAX0y+HRzIDW/CmpaK80LP5JWIaLWs+n7gKFK/wr
SSsfoYPh65tBiImtTQJITFx/vILyignHF26ccgrtfCyoThkI/lokxLabooSPKva6
UnEyOcWl/soeGD4jQWK6Uj02lKTnFCdPbpvPy3xlRDVIVFcL2cPKu9uwEU7DOUuO
biGUrVjRYhD1f4tFwWK+b2PHzTf9KfioFdIEVnP4LUWNuOoDxWhEd2sILhdvP331
/JT0GusM/3+68EnaP8r/yu7dP5kVDQJSR+CtkER0BFAi15o74PVOBmO5AJHSwZDg
0ahSw9vxbQSE9GZ6enzYBO8M7gj55BL6OsY6gCwDwGpYR94y7JnpnWIxjV3tEiFx
LcaF1WcmHm472el0BVFoslD1gLYgaN6FHKt7zlDgAQyxolKbSU7eBfRMa1ugnDTx
0jk2G4yf17DePIvb5lkzxSTpqrwgdtR42Y4VedJebHHHbGOHqmSTRBPB7suojQkX
OSS8W9ODnw99giiVxYsdcbjmkDCN+0u6D1GQNnJG9WWg7zQF/oUPeqwKN4/UQ5eZ
V43rYOBN9kRa8gaN5BZ2uetIqPQlW8CfhfoXP9yymbRO4EGBfW9XO02ayWzyb/Xw
MmvZdrbXtG3FIW/IOd5b0V4vb+MZZHQBbwzRUXila0RrKALPnSpwgDiaqEmWUyYA
zzjmpeIJz0UwAZ5GxRIHeni+txZa+0gOhJ8PzKf5nbOnwD6Tv3kOty0S6pQDPG2R
98lKQScjs2aN54iFAYN1o4k8cxxanSxxiy4wdRBmniWWyx1zBroyL4gGR2x20V3X
KcjsCjOlTav4eUtjryEx+zsz0wfG3pkQegEi/KSADeEi8jzrbdcLWFvltVaZ4K6m
stk+axc43dfg0vwGgBpgCgq6QqYLxT7Fx21NUUgbX+VxQdIWtO9XKH5PsyO514lI
EZqf5CYYU2GP26UmKjk4RFUAeaaG+1HpiUpEAL8AkfwRSJkcBsSda0YLuL9jj8qG
VKkJraFw6Nir1GjqOv2a+SzEjHFEu2Aa0BojdUryWlwbpFGPKdk+ySa7Jr5MFNTD
PhL9zdPHtw8TZmELQrYDPQHlKJlYldcHzY1qiYDP8yQTp1J6MYKTI/Zqwh4Nsflg
SzdcYLKkaV4X24Zcro8zWP6iTS5kD+IUpR5LcSG2dUP9pcZwgdjm2PMyqMeop3IO
1V0OuifFRUjj8cdV6zFUi4eNJM0RsZVmX0Q4mfbgQU3MKuAouTFQmht0koz9E9z8
lF7eLS1bk+of4cWNNhCEsRnwnb0w7HvRT4hmKqv5ju5LygtBdiI2QbRqYT3JFGx4
aNFJT75MiKfb/c5dWVqU3YvvEHaEbNNcX34u/brioWaGndrNTneUXV8ybbYSkWMY
emPq1rqupdgJDKADayfiwkIKETVTQOSHHeBKYf+SjYJXcOiNoYgadTTpTtyVTe3T
nGVvnVgO81n4l5QoF7WRtfd4DudumGxd0gqcM2Ny18ckbec6by76MW2AnOjug6xa
YmvAhnrjSKL0/1ZPSD48XL1tnCxRV5NA8xYL0t+sMrOV7x7oHzB/2hqPsTQJlLHw
tXTyccaF2j44qAdfVbvvr2GYME2qdxbS34q65TvQppgWRd0uT7iZV+lsQRPaogKr
KYzO5bTNrfrLYKagGlBM7S3BVYxomhL3HAkbIgL57RfWKOprQkJEOt1P286sETva
l2/Yq/VSG1lxzWeqNgAONwTvB3LdJbx4nMh54QTYd9MSZHG+aI0Km1f/7Lq5JaMm
pfS75K3Pn1nuaZ0KtpHZgAFJEEMjsA+6tUzrLxmY8vmCdpO58ECqZIuUeIUcfxkI
QS7/x62pKFY031wU1X6OBLaElZYVS3D0PJjPfCTAmx1PDiDlQs1M28Ij3ZrBh8B4
uKziJlbWWAePcibwfV0UGegAxftveNucmCDK8L4kOq2UtPFa/TreVOwWrRQgMKWX
bbo07gm+v3GJqCXC2srce/5WLjinI1oKbn3W7XfNmtInl9YPjD//gkli5VOtGKw/
tSp5DSex1rJtQK4FIBTUzHFp9+eYjNTdcW82XD4Zmxi7Bx1guhLh3ln3tVtLIfJv
c1TUddV9Gtr6tx2q15OmjFGHE4nLlYWc+ADG6sFTyFkoOAbGMkVYFEJdiSmqQnJ0
DCAcfyIhm7T+WJ/GpvVNGhbG1eWFHZiUGOItK9UPIAAT9s4araShzLg+pXGlx9WR
UUlq7EtByoTr4Yt2Bn8+dTrs2XBkwYYkgP4j+CiHCkudhf9deOfribDQLcjATDR8
TfXibC1Veyp5YPs6grlUozkv3+Dp7+nc2UbKgaeneyGb5sezdMVGOpioOM9sILDK
cb81dsdqbnnSrXkr1FO1TM89d1UM61ViXr/bNhUkByA7a/v5iFJRhfAOZl+bQ1Ew
HZWHjP24FzekQurHBjkjNe0xFD01yQR5pw7ZZDvQnt7g7WUvAFhha2uBDHleQsip
Gs5bE/U/FVUqSNRf78DBg0ohLxW2/YhqVCbSWm/Cz9FUN1pmFbedzbLv7SAPIGmJ
PmdCUEUMLT2fReT+2TcCBWedm/1KvXkiYiWDMbRQBBHiD41wCvKotWWcO7GWE3Ee
v8viEXRG9lAD55zG2IYoI5NXCW2f4kRnUNTsMvtLVOIpBr1set28TROSs6fd9Ywg
ck2YG4qvLofY/Vo2/GkDJEy1Gh3MXZeiClHSefsv5Skh4SFNUTjJ64rNO/vZUbFf
5gJ5RuoMV9BOjXE/8csdkS5of3jl4P4IJPLftIvxZq7pVDqlqcVPoP8523L8bctb
2YB+Cq7UubCncEy3cK/yu6EVrQvwbHi/IgPPJ/XqpaUpVKYhwEoVKPiq7+sAugmR
jWXVE9IPatNpdttFpIAc5CDrU4KsIiGca8t0Nq4/MNBXmQhesUwOD8sw2liheViG
yMFtidzw6hSaOtPp6fro7aHbFU8z0ErZFKFMNM1qHBEmX/nQu1Uv8qdR6kP6Bxwz
ce9DYwgpiesvHRKIHcNwEDv6SX8fMhcnqDtN2PL7EcV5+EFSD7a5grb3CNXMB1w3
AiJM5qttEaPbqkA5H4z1RcV2vvsSMoZhO56Jcf9Xj9w3X0CJcV4IXQJ1B6lCF7vx
NkVREv0Hn0uko7ze0wtgk+UcDOaT2dxsuiVzU0IrlYHLncRgSicZ6ZL1kI+sKt/t
RZNHVMGJO4CigqdqyRObqsvqthc3NrYaKY7JIrp70FoEQVEtO7RBwgY+cYKjbMHl
iapOpIvzpejdMG4CVAyKjgZ7Xd+lUz/6Ze08kWckThH3BpO0OLkd8FokdTH1lKvb
vMF4oKGYZima+wha8nZoChIv4emF+zZRzh45nlYGBNnuK7BKty0jLNAJr+i9ejmV
qb4k2fTVti3SzfCOFgZVAJ6UQdjAAzG/C+ODev71tVql3HuI5q0fpX++JtB1Jw9Z
ACRpeSuRtXuCYce32GPGJxgtgVI0L3bC21r6k+jC+xbjzfkGN2ofl/QcOp6XI+yd
dKpov6i51yfkTifViaCxM8rDDo2XtI1wqjTbAmz2GNn90Rmq6auXu1h+P5Wcqs7f
6akzUtTZ+YuSKdaRgMxe/NjJVbO2wGsYA+ePBb9zPRI7Sw/sJgJGOeysS/uJZyDe
joqCpCnoKPQWSynoST6ZrOosjngxwWq1wlQM0sPGUv2atELMDVYwqwZpxKqCoEOI
NT+rQ3ROsoj0ylopRAFm48vz46R2HKda5gjIbYN4ZG+KaLwQ5X+7qQ04DqPH8PBn
VQgSyJyqFd2hWiMLsrcOFn3xaKrwANUFp26DeDVNdWEKCMiz30048CyzhxgkSO5y
uoNpJtBIMGAQgpa/d/IT9H3DcOLaNKgf+KZQWL0hxc/1UauTNC/mcNhoZ93KvMkS
lngkgAcxYQkhTLX3XK8wi38M5zwZLCrG/eOIIqUUy8zBQ/pxvpLyc5HIIrRCj9CN
2+2iWWauu0gTz+ZBj2OF/KsI1dQj4wwVEoiqDMzWk8wLvLuoCZ8RMd/c5qfBotLi
HhsU8NIQ+LeYFLBOCaANcsxlv+yjHd3GMoyhzIu33skR/rjmPcvyfYRwOxPwuu0O
sUTZFvTV+OaftNE7Y4jitF5/vPeyXpe/jNJnQWjpnFzNkPgIfapcL6DbvJR2yzhp
GlcHLmi6s1aR1LIm5MnMulGYNPmiZ6IXhGhP06x1m/OpmOe9i4VAiJUsN9Iby5jv
HsCFxxd6WQpAL5Zz8IRcF5SzRH9MUNSc1C+JD1cc9eSRFexqWh+OCtF6pk7fx+yI
iIywiknFVmz99k+ZcguT1OJQfKusFJ7ZEqiXau70vFM8iIuRWuUZmGf/kyeTv24+
7aEjs5QKYXJtig7bsdZQXlnNdvSfFFmwxGfr24gYOk+UHcUZtl+y1zf61pAHmwdh
wFoZ9GbZ0W+PThqS4+fDn2TRD48aZ6ZufwRk/Md6jaLfja3m/dX2yC+S+OQjFne1
7vNMzylVi/pQSN3NCRhEF/r7jRJTfqSk6I/6xTV22g/sYHzT+eaCpTY3xoNZ8KNN
4ufsYRdKTcSkIKvYOhM6Km8UUCrQL9E0UziHFNMnv+BXJgdSZlj/ILcXUzIYyOrP
DB33LsAlUXxXUm+YoAGFk7jJHaL7/DQmivtMNPptQ9RXn6nMVs+1Z2X00/qnexG0
ZYcqazgcDhtRLufYOwXbXOPBQXU5Ygb/UtU3VFoVeAbAUWowOmxVpM4UPel1biFK
7MWCoHUT9ZGxc2H7fHLu7DjYznEsh52J8aCXlYqzWmYvoQOP2rCUozy71+vV0uY3
9120PSNorgJpbdved+eRnxuDVIN8DW2v3MkEUhLq6oErRfztvCEX2GEbzxFn6BFk
2uxsX7O25gTqW6LgiJJLNGDXYhM4XaiazfgJGfhZ7HoDEQAtSfL+fowP9+JWAJFz
pNuAQy0T9uUb7dcrMMsDpGNj9KEoH23Atf92+TPU1hUCtrrVVvsg5F5NfQSyCbS9
vvbmJe4b3Hc6F5K2jNC2bT9KMLL2jCLUFWTYu6k6fw7P+jyirH5HsTqDOLkHFya3
d15sgDf+voXV5+8fBT9ey+EAhGqkFA9vuymMS0pgAkEdM078sTUOnPR5sI7Aragd
KEHhp0fdHhJcQ44NQMtBJ4KLzPv1kPf3eKvwzZwi2kswnQXtDnp5/j5OLFBvFrC+
GdD6SSKVgRLnC9pjup72N2Cm9q4hMFw9mpETpP3tF26hDhjtUEeoi7+y4TCLdGs+
wfvXiq/Fard5bhhO8499GVik3eiXZ9QsA1BaqN2/lEJRuWwaRKcjpUTIAyEzZ57o
KgA4XnhB3phzXs/x49vFShCP3aoiGn4B8KSxpcfi9loayu/V/bPGJoVhPZXeeb8n
44qwq7qLuwOBw9RfzBvFkqO/R0fd/9XkuJmS10keCDzMm7UGgi7Cee8JAesfczm2
57+wUgzzn5H78Mtl5+XsZATb8sCzgv5MN91JNS1tMyLFkBfD/puXrQIonSIYEw1Y
qRgk1SOROPyqWt79S67vTW5juQ8F4MBdZF6hfBhMKy0mhxy0LUbOTs3leCXPKNwn
niGI5Okq5+RwSJG/PqzXSZGiqNuUUIUCPmDh4saJClHkqLaQrT60ossWs1Nm2NN4
Vkkvqpc9OKmLDi/FXoJ7WxFgRWvB5yte7Qz4FwQGz78yB0OOx+25PMLXEqimQxps
NREsgrE5a7t4MxI5MDpyYfBlMKPhcQzVl0QNKxOoma4YWH7V9WxuHbDdDg/HmgTM
PG9iD07KXTTdp9VY34vnuYGCtUbDJOJARkuxC4etP2/XLD0yLG95BF/jLTFuGZKr
p57MNn3nNWmufT6P6es8TpX7+IGWaLlFoE900VC1WNjbuyRHFY/LNhAZqtiiNnvG
u4GQZk9j5m0KURypQhAPKvdrrz3uXE7A6EjkWWcdW0hBrMrl0mV8a0uxAutozfkg
Xt9gZsicTOwTgrrSTlY3Eg7oUOCK3vhqf0r5Cca2dybKZ//4AoM+V6Abrn9f1HD9
dEhPjAG3UDEvBNiYTR3gs1H5+9p5yWcbud5nKdV9is1lzBQg7Lxyy4oLdfbDFKRm
3v5MdqKz3cpzuLP/cvA786OM7FURvDW37ufGPuKV/WbCvbm7SPf87+cZp006SBZj
nbhi9hX43lQNulVrv9TF3BKjTr/dVPz78xd5OuQiqpbBrUngELkjPZiA5SNtLur6
907znr9uUTKqUVsjoPoWEB2AW/jONsH25HVK5AL23hqwkDEgaY2r/Qj95o0fUdqN
uz4dHpGOJ9gex4hzFkPSUqXvH7Rx1H2SB3nXhyvyLYtarXrN/8U1/ZmJOs4emL0t
d/X91WOsgZT8BYmrYVvb+gvDQORXLkYnwzxjRC1UEFFJCW34aszrCvPBh7bsMd8t
H5v/ypl3BtB5aPO8SnAk5f2RHP9EOQuXlllk3UMfPTn7OsXlZZuLLi++hShW088p
fkuuytyfmBCd2SNquG0TZ+/nQCiY3e/k2XxrWktEV9NOxy0U08/OwytCxLr+eIWK
JjI6hyxzu4YmLobvtrVJ97tIvhUBUycuu/UbctSDaxuP1/Pc1eAh65K6ouk0R8nb
5lRKhz5OlAj93NCGHChO0Q9QAyhFkif1t1JWxOzAEAn2pgXCXtH3WFsubz6R3EfI
MTrNGZZClRB5y6274Ys7pX0+q4izrlNy9eZiX4OXoHPy9PXTX1BpY043a2+g4FPO
oDUelSAsghIa0/8hTVVaUGJdz1TVpyi3JKuLE+51Sxf7WS+UWwCSnQFH7U36Q7wO
/UWQ2W0a+F2V7cwsQeGdunh62u5tX21byPPpoQgtISSWdOFeP6VfqOpIusZEXbFm
70foFqXmv95wNHdXhMkT43jm+1LgRSp1H4l1NciKbC4dizepFSoi/ID/onhGS+lV
iouCWMOXVBDwOEk+3q0oZonISGueiPXrMNu0AjfmlH7kqvoj2sMPooGflZyaIzpj
In3quI8zoObLO9f79SAozkat1tBvZT9TOYNRk9AXzO+RePEhzslDFpNfF4da1csv
gWs7H2hcqUXJJjoeuQZYfJHKQJ0/2pl4IVnxnXGNJ9QSC4Xtc8duH9jsEtBXJJmo
SqBtw9WCk2I7n6qQzr26ehv60syW2SfmtbJdPBsWRcnbAPeOtQtpBlqqqYp4EJI3
+lCwoaeOz2Ggl2Ol2F6yqCgfXBajTn+ZHZ36XgcO82Yv4WgsznlyxPvbkopt6gcU
znPbJMn2us16YOk3eA8eNWULETB/grCbXgKlcqPJIyTuHv99VexPChROU2UfpWXH
bYhO6RHglvsZe3aWD0sFRgiZ8H36CHoxWK3HHCyl2ceHmSHscPexb6ayaFl8e9lA
3Uc4CfCV1HeYOMBDp5J7FWR+9XCEdxe0Y4ukjYME0YRi5GLE2DYqnNgXPOAayUlj
b6S3Hsxm6Q/l7e3uQT5kdeOCX+N0VepjHuGqmL6NWdCkkSOIAbNW50x3TXrHiEz7
jRWtMEZx8XUC5Law+BwDU0ThE1AC6ULsplP4+4SRWrt09K5abaK/HqnRJAEZFTt1
D8gNSBswFSmODbA9nrzwWA==
`protect END_PROTECTED