-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
c3QAuS+Y192gp9fQyI9yIXnLHYm0BrR5RLxPpF6u/3u+rs35lKUyjEK3lPebouITlzOrXLVdWw5/
0JUPqzTF8I1CFOejpU9yf6AOY4GCh4/VwBfXXuYbeqL+2H1Zrkk814jq1zRDRRPg5WhPFzRCdLxK
Dybf66e9hGMYVL/dr8rTZqhoDbqMDRsdhhpb5C3wwiMGPZFiR2u8onSN/tbrz9x0CG870yOsSIW9
gbZRZQbCcwYehCt4/zYZRBq+BttjlgIAklXmVVkbCSPYrYcUIRe3KWXBIMVsZgwS0OJ8iZ1zgzcV
ji5dYpmtEB4LdacyoIjLLvQnXCS1jI0+x6CGEA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5472)
`protect data_block
XJq9CZrSJR9nwafkh8qT9O1v3cKPQPCvvLe6GxwlkJ59IONwNlWOV6eD8ff1O4smhOJABFVIuJDZ
WT/V05FzoEbvOo7uRWvFsrxX2I4t/HaJZYmdo/PbR3DH9fF5GEV6GKX0XokkrjSsL5AGTdRgk+f6
fGWnckrdVNPFXobcmy9ICyegf8GnxxV0ikmpFhA6mluNzwvbzUuehWfJ4rqXTJzgU278TLu5DveW
AJPi88NevXUwlSAnI/ULJ97THxJl3bYv0JtiX1piJ3lZ/Y10zIBZ2IgdhcSB5rEi90lvfgqx393v
nYe92Dk7slH5g/acdfBMUNcn/LAoCPNs/yVPqWkgLf1hsUeq6czZlAmoVffDYh7CQA4AEzHB8ZPd
fNI/QAWLGQjXVQlWhFXZgRu1P6U+znXvoSZ9zKDwal9OlAgcdT8O2gt2PQGeiy4AKYGN2hZoxR5p
fTwK7kLULOSMPzO6v4h+7P4qzwkuy8w6wuoP2QvYllC3pcL6XjMlcj9GkuMtevWia6hw0OHLTPXp
gBFzeIYIL0VPBgcE+v30zhF+RuR2CvmEly2ULzJAZvsp1WWSXMtbwhfa+xTGedkK0FrCLGdIYwZN
DvQ0v/fJn9U51pNVb8FiDb8rKbwGixB4jwOhMJGGu7VQlQ3ormq0KCTQ6ETlG8zeAbIs7ys+6EAU
+bTzvbsdl65h0PxIRpiAm10k9Krq/DKG+UYGp0TFNNHN06xTT0chLVlIdbLJELUFWLAHcu126hR5
OB9rvFG+iPFu6ciYRpvRniEtVUs40Pku7lklJBE83NWOiqMhb9zT2BjCDlrF7Xr2tnIB+YiGak3K
xajaBReBpBXOfa72qkhJFNnk8VCxJ7WKAMVtsvGpKmWir1c6zqaqjqdN/EYuityYeNAqcwS5ON8k
oHpqTuKCcO8K9WP7yuDCdvUn9CyspCQEU97gNAmDdpd2ms9j0RZKtxHkUhY/Tg4JVB3KFfl0ExHB
a+Yn0CpkI4YDLpvkkyeBGrGPOzVKmAh4k5F7oPuOpQqrX6Q6HHg7iqWYp0AscLjZViVA/WqjvV/k
vpXXko+pCvsIFjNstYAN5Z9rXWld/jYqd56MoHbIrnEGgkMCNysXj63pXzAoqeyKfbXvGKc+9GyY
9ppRJ3O6CPDiMXlAH7VZR0fxDLibUQjE+ncuG7QeVjtoEb75tfZ346qXfc2sE6z7AW6foaqCNJQ+
wS8sJS459qM/NV0XOaQqQzDGPSHCmWVw7mVIqXU2JfnSuezX8oFTsNwzhar71VhKfT0CJICWpk4g
fYlRet/nFcPUwKhayH3phz+KtWSkE1gDo+LWaxmeTlpEcIjQH9iSqla3aknGgWE7nieMO4n91RYq
WGLCO84P1pnDzLdZF0cbbVCdR0HC/fyTPNQMJ7re8CH18Fu969zV1/49zwLgc0DOux52CWkm8/M1
OoD6UxVzkycUGJWqsbHKeL/oH/aza27kjbrOAl6fJ1mq19nrSUHJ8CVUGnSJzxl/Wqg+hd/06CiT
BxAkcSrkcPsjEc5QONqhHHBHkT+dMXuNXkIsYhh/IrsBY/V9lqtOQdL/tUScGSeSpp0uKNkgWJES
wHKAyOKtUhmnUk7Te938n8AkwaPRCHvhAtMmnYnp6sG6WsegBuKBxIa0zpEXPKEtyZHlJnwRrh0b
p7LrcA8e55G46gB2TMp86Qx4i4JsonbbWum475abYT5VxAixCxf7q0+S+TY0iCSSvFvF0fH+qxa4
TWz+/K2InIvRW5UQayxcFwMpfq+lbyCTVusYXSZQMGvl6YvLVB6Q757PIetbm+zwJ+4LTxJiQR8b
LD9xLzHJSYWcNo16LWIEfE/qot8mZW1R83i1xl/3WKwVIRYbIekwoa2Dpr/XZZxC8xeYT0qFMQJ3
UwJzmjBCrEGBvLC4fIvNiYbGj/7jGpiqrd+dRnak0oOXyH0WqpTnLlw+kauuStEV1ut7xuFJzbai
+e4gLdV4BoN1ri7KxJrcI50qImiOjTu12+FFNrBVecRfzGjK6UO9hB2OVnSySmqWCZPCKlVyWHSe
sulD2FHFcwQ09WxksQHxQVGY9tnOB9pXlgjQmKXjnaSMjk8pXMricpJBOiGvWknIkSo+x5qx4CV8
vTLW770p66TJaQH0RtOy+2f/Tkyfr0zndskZuEDsC+K48DetsEBabrMdXA0gxdmMW8u9b1JElkbt
8gtW5feSnd42B1w/g9Kk4sHBrGm/sS+z7ocq/J79PJDxaoJHsrjb6vY7dH6KgAtUyy+056ggdsRk
IO9BLtlBpwg+fOBq1cD3SNfJR/LLunm8Hjp/qQhb3VyFU+piaQZACxjSLNQnKCW+GziGkWaRxTj4
psgrSn+ivGRwZ/LdgVu8bEaQS2ZNwyd3rxgVBsbbtBXg5E3RW7AGjV+bvC/rQd4rvGB5twZ0Oh/0
XYF8VLorBuIEyN6H9KAKjHnlZxCCkN2sae3C7QscwlS/kaA4vf3S90Cw6YGbtLYfEvH278zmIyQm
CbsQd06AwJHtefUKV4LaSkWfNYOU9daFtipGQznSqBscLel2Oev71hxoLcf+J/J7Jp/RkKAsZK9E
mkiSrtUrqG5ED0InTglQQnXY3sT2fD1fIJDJQveMzjXmLmfndoTpO/Nq5uPJ3Wa8eMLAxchRCR4+
oa6GMvO5iA70HcpOm90xTj+J456YjuiKIx3MRoCIb/b3cxmdjDOfr7Aosx5tFFv4HYfgRINjFrqW
yBa2V6RSpzu8aHfC9/xdOuXzqvBB8wee8y3KM4w/5t4AkPVD4nNi0kBUXULAUmChHWH5tqxMDvUW
PwqwRab+rs0wrCD8GY/64WzW3wB/Wz6K1Tt84Q16nJyI4FW7eSchi6JFgldD44YtMm4rgPwdwRuR
hRyGEYOEUMK2FAb44K5u+GgiaknTrKNNqeDEIhIvz+7Er41brTAw5zelVHHoSJ+ixC5FphoE8C9U
bZAzW3QGtv3RO3eppZc2cpMvoxGVJAvRLphuK/EpesH7WP4M0z3mTf4Y6bWSaV8rMDrcuRjT3eRf
S/lWO/GOIlo1RSfhfSw8LuUEIHWVdOsyOJaXLm+ZyvlOamSoz1mZatIumhzLeMKaJxcWL7aNQm0C
R0n1BIcsqmwUlLcMx3fssTip9+F2aeyNPhshnkTCmCOArpnlIOyUnpcukq9e6tf3tuQdr3owlXjv
Jozdj8ZRBzwqD0hFYY0Z/YChk7W+eZzVOH7/3Es5rnBxGNWnjmrixSxm5442R+IjgDHpkfmHNXwL
Tu03vk7jRPCGnWleQOaj5GoXB84SXPi95jdO/sdpnSnuf6NhE648sKoapAiHPw1uJfhr120/0gsU
hv60ORrLXye0kRHEDUffJLP7T3d6mIEk+q5uhd2BhOZ1ecvS7GmRzPO5MXYMAKhXDc2zbkUWhuHh
aIfQoq77fUjaZ5EtgVG6rU2GmeTC7C6LXLekOc1mrS2FCPYdNjPL6ASxsjgdIyWBEgG7AXvOG86k
OqEemgXxXwUI8sq5aT55gkbYOulMaqkOeXTH/xu0VCDSV9s5CPmIFVgmKql0iO3SyG/MkmcOto/2
bGiTAFZPTzzrKVTk6zQmdXGQzmA370u+TCRvNaaYTvkeUFrT+Q0nZj+ChgUKPdXk5JSfcn0vymmv
6TdAcC3McvuEeqt15tff1MW4XP9Mlm7eKBbWKJmb87ORyeEZPaYLMSWSGARcnX32HTqLR6EbQMO+
l6hI1bVrJ/dXK+b8YrqJ+hOXVUD70HVPZQS5Yw7+SF19/Q9gfeH35X1tYsbMcDp7gL/mXQGGzXtH
ThR15u7D8arWG09DdQp6fFi0O64TSo60SoOJMOBh0/bg3MVS5tHQtsO3oTzxVzXYcOcUd+sww4m+
9usff71ohdHOyzeIteR7zwyL4N1+5B/4gz+ZnMOpJ4/7rxfWRvSPvom4oEC4afSH3v5aG7w5ws0S
9YbfQtfdQD53OGMY9dNn0TmlZ+noAzngzAMpanIXKyGZnIvt+093Pm8RG2CuRhVNJ5Fk7H+S2Cbc
VXUkMszKxAJR5UKeeiaFfAOnfdJl6bWn7wKLXmLP/9iIwkKluZLNrS9MXdSJMHQqhApSA2Uzw4Ri
rmxq3GuqWf5hRMAfqtMps+Pabztr6otOKEE6TxEHrEDoDKbYcu7GNNjKJiL6tq5lbtarvJEGSWdN
6Ta9fVliIykHeZGe00RYJQGmREYMWkAckK1jtNDGWKqJ9MPuLrvvq/OGAGeEARyOzSnBA1952dIa
/5FynjLe0KKkfplTzTcTxFaCyHSaNm9PY6pH2wTWaao2eSA0mFHURWXcXp9esgdet5RpbrJbfT8n
lY5m+lLwHzt0xa0T7WehgwATrcWiWg0Mmhu57G0oJeYMYZXRZCPY2pBeS07DoDPbZRUIA6RoKOhJ
wyDrUoQHC7F/E/rFjySpcoqgjSMnGGXvmgE1tPwYQiW652MUWDyIJarNTkdZGmnfV4RikeFDWn7D
w7inoYyxshw3AFwZeDn9v21xC1uqlVE4a98mRNFeT+k72VxKacK0FDExar6y1p5RX+KRVh6A5d7k
jBIR9apTbR0AqjFyGQzyCER08iNWnJPvGjHlc9s1OxRgC8P+SUNvabYVpt5Lg1xQSjzeW2ENUAIA
XAY7hKtgHXcXfFAs0YonGCp0X9M5IniEENDgaBmFezW6DDSoeEOZIK7rhr9o+gFNpX+oTb37b1rq
1Gg3j/Kck5DAYhg63PsDyw3M50cOJg21RtqKrNKb6SuRZHYGCaVMojbycqClzGRJenandqLSUYxf
+IpcVW1wPqBWW9KQgyxSszh+wYyyjcIXvBB/YzHisYGi0p2JxdBTFisA+4udog6ROetoUmUDLev1
Xk7u/CKIqUtak0kUUFAAFlYhsl0LKKPbt2yVow8Drf2ENODw6KGWrvfVuZD6MCOwUMjireobRFmw
6KCNKO0PXTSCPb5i0sUJbcAtXlVUHbOxp6FXD8kr4oGzu1iu+Sn1HeaqrKpZOB+uJm64H8dsa2rC
UVzV6+mSiS3pdB9h0W/CtRnkz0Z78T39btjBAeVaKKzI1or8IRyyS6tnj9UUilJbToT36BrOEEu5
I97vEhHfgUqr313SKHYVJVB24bUoKK8Owx2FZQXQCnx7FQo9RbcWD/gGIfagQTBt+IKpTwqKnd9d
zetxBZ5KPg9AbR6uBo2BsFnqo7uhgm3EOp+6qo26n7HPV6fqQJC/SS/BZOt9U+XlNHtjJA/J3GGg
Qfy21S9ZOJD9XExJot+19nL10H8q6K9bFEkQTTOV8vkBTc72nbhcv8bauKvUe22uNXGdIDi5rTmR
i0B5+PwBaDEMVdjDoyrOHNTmKOMVat8DHZ+phtabd3M+AFGYkA/q9h/r1fMnXi0zUGPrrMrpWouJ
uKVomVP2G7CvL7ul51NcsrQM4bdnKdEW+JwU2xQKAq3IIKoezOODl38jB43ovUoiLpZ0kK9JYQgc
9WMNOTVHsG2l3j5FkUx/tBaCCsYpgnfDgYXDuQMTso4Bj9OpVAclcnRe34jwNDOdTOTH6J5uqavt
Oh0XQEj5OBevwt5TbD+B1XeUITcLiUzGbDr4I5EDrPeh2AtHaMbZRdugZsfRnap722Ougj68C9GB
QRePhiGoOUgUQBSrSwH9P90YOMJR8amBuihOeiTtUAX1kFFicqBBFbWgW95Pc/dpbqh0pyWY941h
NMco6C8YOag7FdndvSDUtt/cYapxuJA2iuPYlSoBgK835aIh2Ja/Y5AA7+R1MydFjytvuWRrK50w
vBmIR8wdkYlPUijYFzD1ZD3Zo5x/UxkVICq7Lm6BEppJqVU2hE9r/4Kk+aHaUq2ar+looelgq9fI
riKQrEaoQN7F1sGCOVRhO/qmTrBr1zaowN3diuDMcFZ+muILeOGv7S54FubkV3c6DkutcwWhz0So
ETdWqONz4o9Ck5yB4Afrn5+8Cpvc+YtMBSJzaI5DFs+E9ANna7rrSthkgGLjytvYhECNy04JikrO
6VgiK97P/kVYkhL1UFCvIzxcJiFiivnQ2256t7VKzuHqFTefC/fYESEgY9PfoPEcdIhvU+Xr7bh0
esb8ORaH7lHEobnXqKeNE9q4PRHo/ZnS1wc9dz8G/41h/U1KQTP8k5N3/dzqYiLiGrnEYDjKREct
AUC+I7YcKy3IB7mcp/MetQskumtwElU0V/isgXODgKOPlbqjb20/dWxTfOw3uWzJe9SMEdWsPYal
EAAieyVoD7Aj3rNenjSyc/OuhNlSzURUiid4dqUKF16M5G9gDkEk6DiRLqNS2cGDtRsHO1YAuVrB
fqBKYO2sfJF2kmWvlrAfrRMIPTh3miOJhm1Rk/cRJt6k/Oca0b9Ql+CiGJ44eDk8afltDHbLwheL
O4FjVZnJo4+VkV6i7KOyagSQgDbqqXceNozdIntXRXkF5EBirIutrW7hZRe1gbLez6vrHOVcXPgQ
AH+oJw+lyrh0B2HjCza1jjJNt5V0vkxUJGvL4D3cJFKhz4w/gyUu0r0DU7VrUqW2q86HK/o5kupd
u3WKbxQvvh3dYKX7PVTN0JFa4vsng9aD79Mb18LMPa9u2b3wzwftyFzvks59+ti6nvLp7xemz31a
Lzy5ggcdFf5kFn1P7qWxQG6neTB2K64w2myP3gJst+thMLj2sh3nGRUfeZAu8txXtUZn0X8N9lWF
4jxvaKmZTFPMOpAuqvK+24d/YoO+pxW4GcnhAVVYGYojFYPd7IJKsA1jDQ/NaN+MfKbfNeof4A8k
hr3x1pLY8G3Ps5WDAW88uXZvQBUKv3O8WbJXDntbLh5Gak6Guet0h3nhLN12NHHlqD7YXH1yIyFH
krC3aqgeenu/OL7Uij4b1uol1Ta9pBvC80M/5XG7zsGI55/fcrSQpGGveKdWnNExBDJBlZ4bi3dy
+kkovnSMCjNIVPowzjiPt7jAldr//Q6GHGfkb/gYNS5nDPRpFlAdliY0QInLHptI89LTM4Z/Wjjq
wwpcVG+mDzhn2IQzH/Gjwgz8YHeS7gRxeZJVYrV4Cn538bQwvME1zFphKko+9fFhCZKqpNdJuZT0
efbuJyquZ2y1ROTAV87hATL2TMTTsI40xMbG/Uyl/dCPDxcxLNWZSxYwCSHXp1X7zJuVUhBz17Cf
RArLRedfAfALPxIK66T5xYKEf2m2O+sLhVVpKc5yT09F6trBvNZFa411QWq10xwXG5lvbyLVUYGV
kBeTZG5hix/usZYV4xZduuru66pafTMVOgILWgx+AFfU+9KLwcX9wIVklN8WerrPLnhXPunjraxe
`protect end_protected
