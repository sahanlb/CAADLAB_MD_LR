-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
DDkg5k6ALuq7I76MtrmZM8ne8O+ZC2RcJ3Z7ig0Gkqow+JD+EAsRq84XAUZwhBiM
M1hPrd/ieVphP4IrPqXRRGF6kHKdQ1xqaoPEnMv8wP+DisExoAFu51Z71SfSWfWF
0h2y7EAZxkg/KaFwuXTkllm4jCDfT3t2x3LcjQS3boc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6000)
`protect data_block
0MLwXpnOn2nOqolD7Ds2LsjX848c8V2YKE8t3JsQel6KrTpjWz0E1z5p9jdOUXH1
+J07oLsVo1Nhw4VPhRuQEbJMjYsN+0sxi6gKe8/NwhVB+5e6sHhyqP+kXQLRlFSN
QnC8Vd9EY8LLF5Dw/zRccOBWkl9/EyDyWPIjABQ80MKaqPkrOQcODsiom0FHlid0
cLzFLKmEiwpIjaHvtZgX3Lbny3Yq0WoZtP42aVJKubBqYHyimoOLxzUbCsdH6ORo
ZcNKs2TTZFQSMqme+I7D7YQJu/S8aO517HSikg5oYHa8toXA2hC5BFzxzShtRPSY
PNjlFr7i+jj7H7DEOpWrIAqwCmhN5D9Rig+NWXHIP2z9jR/np8Uaqh76DmF1pvoA
w/2oakvELVclwmX0qVtyMfHPYCuYwi0rlrqdoTv9AWwIwu73+ACV2Kz1wi9f1RCy
gEO3Yj5UC2li/wYXTm+zkl7XRbwaVCJeEvqsSLBlODzNG/J6QUle9LQIi7PhAF8b
kY7u11/Z2EtD+ph0wVEwmNPpqBOn0rA/W4pgl76boWjRhY/ZF25Iur+yB+Oe47ok
dHwYh135U0n5XIGu+RBwIu1UbePJ5VqMgzbrtatZ4qTnMEpYu+yyvJ8FOd66QtZ0
JNrHqOaNZkxoloQltlY4MxbGWMSfRk2O5A8yohFA6/HzolHpApQb2F3vN/gi65Ub
5ax+7Iyrr/FqTRPQUyKVu9eVh1pdGP0b7/zygQUa5oSnKX8/raJSdjH6yy6UQYiy
M5YU1zsl8MdLAuXDJbyPZMf7uP0ZmfQq8UI3vzgtXVrN1nETyYwlS+XZ8g5MYigf
G/iUJaLBTlKt/dvJao0YrUw9q4AewK0nXQtTFniEkotAemMHkuT2PN/FTFqR4pO8
gn2esqLVuQiM2uxOtaDTfrM//1ZtU9XFOjFbl/659dLLbcT2Ffe+KFdbKwlrkNiZ
7lzRqvDm2Y/MahGZRxZcgyFd1ifQMJI/Ww8KtcquGImyENkEhP5fpPQ6vHDfCbMZ
e1OWSPu/oNDksl63NkkWhvIU0T4T3twJM+r3Iqmk91OyPtWBWvpymdm+Ny6yJOsp
7zo2iYzznJUor+ksjI4nyhvBe0M61cQGacSWm0KqYypcpnA4mxMJFW4wlbKu/hZ1
/yZqt/xhUu/5SNnezvFMbqB1BCKhApDcvqVA+6Z5Pv0fe4co6mEuLqF9uMay/9Q7
P/Osbf2sT+PNlIqnS2VX7y3Mm0G8PCxZC6NIPR0l1H2p72/6IH4vMJsC1BY65/Ef
ta8FMBwsFBDm/PRGSflAYs9cumbY35qHWjFipn/SQ+9g6USWA+APxg72maklO02w
y+s7QFEVqLQfuyBBEyfi8A5kQ8W/IOTm7gXWrebnkm+XyO3zn4tQBEtyyUbmdMLK
4w5VopSUZuAq2MRJnC68qsk9tGCfl/nj4RWvWxgYigJmhgy43Y5z61ztKh5JZLQz
L65JcmRcYyT5z4Lkm+XZ9e8wvTwPuyGujonecFaAZmkl+lC2phQBK4tvz8YS2KOQ
92pSOMbE628yvxULfCZce16dBqSFX3rYOw9OuTbu7+2eEq6m1oZlcDyux46KNThy
PrQN9UGSkQTWNkX7J+kYEPzW7JlK9MAKyjj3xX1MD87v+9iunPhOG7qSLK1BrgSf
Dc5qZzK7Nw0fndz7Fvovb6VEpzfO8Sa45zberI3LQ5EBjheZEsJc27TBTU1vSPEQ
Ee8cE07+JUHhuLVYSbVRBgDcXsdUFSjLyaUkwMNlbFmUiDXBL/YwkM35FkDUQ6/I
vTwK7mXmvtk/p48YmCFYVBwFdzafd28ghPuypFFJpFu5OkEwUxhz1cfkWDB/t0Vj
uoS/TI1pSQtSDJAT5s+dyYlWe0iR+npp8eaYmEPA8CK8mkMJ99uBi/J7eI3RwvSM
iewYmYhKOd1QaYVb4Igze+kKwpo2wtmvgCUdSqyrmWrGhTN2PiUlVGv1gcrDsn5w
mSNWbW3bIAW+IsfSMKOrcqR4m2sw0xhLQbFIjMLW3Kj3tAZdp5wCyofWlGjb0xje
vqgyC9eV1zSpoc00L8S0g4Ol5Ssjon7JwrEZ2Qj7w1fBf3Ro4xR1CKESVwbup8hD
Q+6/t6TDln7IFCgk+9p561N/hdvBxkUoe4QOXoIU8+cAnTh9rHlQ04DK45F2jXiP
e+eRVmF795lcF8NliaKqv5bBQdVuzgLHosNyVNv89J2KW+Fo5Hr/yD2NhCCyvJaT
5gx4FH+xgZxY7QLK1Vb71+eMjQWhSh+Fu63ijGBLkyFiuOe2FuEbXP11LXZXzgsm
bsu7Gbl1FbDa145/SjwZiGTqh5dxpVrzMZUMJzR9iwBrlFxhqVywK7yEWFulRTBP
oz8YWwO3i6cb+rVbV/IDXn0Zhs/icwjQoTJKxa63g9jpd+VwwBxuWykVrGrqmpJ3
+y0b2UKG4xrKJ482xI9L72VBnRZZtmsTinR1n1enDFEWpi0s428Mm9jSW1wOC3Pa
DYY8CaZdC2HWNbRliVTWZ+JSM0GoD1MCqX+A2k4nK0ppqZO8s0nL/I1UsNPpClOs
76h/4JEWACKHHbfN3vyI0YrTgU9ydq+MeYRuP9epqM99wl4MLVej/ck03pOpHp2j
2edLWa1ZZRh0HGzC4NlGrniE6zLjcWDJJObm3RiHDOVPJkTF6qfXmox4ZQ0BRxPq
o/mWGuIW+5K+6eXxdLNWnjUUDltLzOeboXOzjmE4CK3YsZhyWEHbZoCIC3BQ+nAW
hQo2KixKgumUMV8cAOqmG5JdZKTFjFR0G7LhU1pp5Wvfel38kHa/dhvzduz317qC
k1FXmCMctGoQTPIFydX0JjgWScYIjPXWLtxXA4d0BD9ZAwdhp6clcxcleMIxFdGE
t3xn4TPh/TAmUWMWtjqIJRVqnA3u/teg+M1KRPHiFqaPadHmN/4Jol4Se5HkxycY
UfjHFIknUM5UuqSp1jFh/ZqgxkMLAm/B+zFIy5dEX6Eb9IZJ1KrTO2KIJuow0+7S
wXl6JWoPvIcVpSvg0rMEqP0UNT66yUokuO1wP+XLhDLQzUPf9SSFcuZ5QfAg4f0R
Rcaohg++KPAyK2/3kOv6hMfwmSztGTgqBTtVLSP3ND4J1PL3qabCyn3VXz+o6J5H
YkHdL3neVIwnDQYJKFukZam7JNZPGEz6xMpMBdXysaEYwZiZwdJ8fZbumGcKlXwI
WQWrgWoTkgwV0EgDN2yJLSMI0G3WW/+uSIhwseQyWRZ5VGsnHSQ6nAonMcYP3yFI
f3JPvm4gzVTWtjj/AArG6ExyUzz1gz86ST3twICEVMx9QNrJsfL/T/DP93ve5zQS
ctzPsN1Wg6lht9D6jTE2MaTHQ18J2q5SwvKWEk+jMLHjq+4wlkhbdomabO4xBVkN
7f8UDGkQ0Tn2hdBwvPaB0eD96oIgXvK/CIghDPkfsGCKsM1Dupc0RgE1C4plfJwk
7heXyCwvXNEHsXwXd2gZdfwwdIyc740whRznfa5t8w5oohHEYdG3JbCgpBcTDSEW
M6Hrb51lbZuB5PhSctZd4ucDGQJM6EkRNl4BkBW17uWwL+9HXleWiVX8VJ6NA0La
IfbFHkPG2NXuc6R3ABACm9aw5Bsm9oBh5FoC+8pKBus55twJLpYuAx2P81gPC4rp
7U0hd/b7kKGqVg2kDPpEu+JYcPiljnW659tfCBQRcLtID33nCusRoelAD57y3xQ/
gttovyEeG+UeDsK8LulhexXw3SNFRkvTtCP6e6weT56K8k8AeqAjhSMSjwXyTGr/
PamW/wz27MY05cD+yboqSjy3OLVAuRhX4phIXxzg+nnX7qEGtuDcno1QqF7G2Rml
HOC4WwZAidz1kq1k5YQeOX+t/rBRUEx8sPW4yAl6hVsZpcGeQgngqDm56jITJfrM
do4reC+liZEYRHmPcCZgnwQHJBHvQm6NpLgZDOpejkvNgSdWN76F2GKz0g2OaKWg
6aBUl1rs/To4YvgRA4sejFnr9ioN7IVAclOfzp5zWM0CNbhJB52iCVPegF8Cixj9
NrREttQ0qYrB5D1mkxIcIIUQm/erHzTagv80jEWC5u9mVGrbFEtQphPVD0/9NYtz
hqrD/kd1hLgRXjOEJhBDTnePmMyNvUN44Zn0/6Be+0rvXzu7Tz9kR+zRDn8fPUti
znz1qIdsUk0/E5KkW4x43CMpngHlbiUTCcttvNzj0lfmkNP/B44Mu4NsPYRZzjL/
aFL7nh9cqe4/Z4xrmUhbBzj2VtG3Gm4OQieFadYF1PCzlHsAF8rCbRXuXtHeflCk
ykZT5DIXqwRJBxHrOuaSAd7LndFG4RaOVdT8RmnfBne5P+S3cougSc3/tpRJdpnM
V/OsiuaqzkKCgNR5txZzDDRJQcHvb3aUC1GCwsjWIIE8Maa/mRGOw/ihl1laxzl1
mVvhaNc7YV6YGZzmgAAtsa1OHXB+GzOEWrarTtYOcRaPeWLmCbfBghNGt97zKXuu
0Nf3EWigVhuqpPACndfnk0zVGmz1CttjcXjT8r9GaEjuknhZuuHlIu+IM3Frbcci
xbT22v9GgDZilnjiNfKlY/M0RFwWkJHH5GHwQ5DRIFXUKId3Hm6H1+BqAEB1JgEh
kjAT35jXXsv6ZrWVPXQvG9dfa3bQgi/FoXdkJGz1V20NnIv8y2Pv0ZMUOheiZkjE
XvpokEg2cWVe5TEO+ycv1QrlkUVGEfvaeQOix66JOHuQondmPz0Xiuu/1DLomcmL
D3M1+2tsN2rco1zCuRPmK9QeERYJzUIzmAA6xRHxUAMHrWWDAav5ey6p0yW7gjR/
zoLVogwTDR5LNauCUxe2o3oXaHwfCnHiV89n6mNnGZquZAPsGGJHGbZGWUx9jYWA
w79Fc7IqMviKfaILgxP2EhHd2ztYrwtejSiL473AfSNqs6l3KWXMvKwbqllHboy3
E8kdaaLViiWT7y2t0GU2VapdLnPSf7GM8SuaJm2QA2j+cSSTiahmizCl95/ZWYzc
qQlu5wCghzGWMJIZjq6PkxZ4bGK+8rS6AvJ+1Wu5ANNzqXHc3pWTGTIh6NbcWkwI
d0OktZ0Rmo+hNt57ahRrLFusyEXlhsnu7VC1W7FJOc5GVpf5VFH2PQj59QWuM6IA
pO7+zG/B/0UO2uf7e9JezKdakTQTITVgTn7BiyQV6LcBjLlf530bWR9g139YKHjF
P1zKbckwZAWuLDSPXxxpimxYuldLWCzRtTPrFyoONktYEZx1ohkRmDamjyRIOPJL
5lI8o7YC/nmL8k8PxvR42fMhww7Bk0wPV8CGHWohSAG8PPhVeYbGHAyDUIYv4+gD
4dI3OcypUUE5WhgutBbhHedahHAuLbv/Z26rzNjvgQUS7jBTHxojKrZN8XrBDUjY
8zIijagMvXDJK8vhy8pl68f2Rh7w0iZtXMfnrg6EGdH0xV56dTXbf7dyzFsmYEZC
2gjcCKSgT5M5vbY/UiCytpPrO/jNwbiTbtpqYHdW0niUbRcpF/o1k8h/oOoOnR/F
24KmyiNT5aW13mwQkoowM8RStfAnvkxsnJC5i2RIEh/1MV9o6+Sp1w5GJyFOGDkT
EIeZpdV9V7yQ+rxUa2AaXQVfqC8ZIIWJtCjwj4FKevCt8sGeYr+WXoLsswFT29B6
p34Z0CeGXPp+pUCw0eugbx05lRpIsZntmQSjYrSBQUbXX/r5zpzK7Pj6A5Tf8w1f
fvuIEiGQ6ZVQdbXdWezFYF6VQ4OFPLjElziUWvIpiCbyHjVJyi6e7xosrUbt//TX
8yMExnXLDsrqAUu7kqjdhR2fh6fb7F7IMlPOmEaBdz4ZCq2VwHtIJkomv3fEVD8A
pXvvTPWz+bl+G6Pc9j250iEsQG07KlfaEWomYXQAzvGdGDOwietvqaqwBEaWohWq
aG+9Y89hD44L+3iKg+OkyJS0qTN/BDK6hF66Z/mNMECgMXUcks78Ww9h7Ywxs2hv
vprTU38cGbQQBkpWeUWIQybVl8yknNpRjKpt2uIAeKcPus6b1NyXaWXDAR2YOlgo
hN857BOt/QnaP7WncCg3fx5eImk9DVsH13V39XyhxgPOuf3yH2xsiwPhKtx7DiZb
H5bVNBVE2dntXKvAafl0ycDL3RipNcIxYadxyih4GiB8IC3jg3RMXhktKn6XYtbK
a3AQTxRUV7vcgw00Xqs6h7USPwfGh7R1iXqsrj9K5LCdg3OHIxXGoT/wdb7t0bmd
f+2f/AEw2F6TAKOLjdTasLadmB129NOgc18QRTsZM8vQx4M6KwCvgtW3KTDvaRki
G32s1UyKK7Pc0VjCorZAmWQMCnbEAhgnBWv0EO0Y/DaNeKb3pyoKC4wcJDI26DOv
auCRNB8KwLWvi7EmBTuEohk195bA+TV4RsoigiyEbmkmwtWRPI3ddKzWcKkuJwzz
ebDOLMuL0cyCegolsbJpEStLwVepO+oUKJrGAGTMUzLVk7T1Xeft6y+MpYzbxntf
tFDYTnEZlZWonefoJkX4Gwba657zRbANadDVylSSoEMqsE+AKwVCWurdK8iY9Vvm
+xhRyRgEtBiLcFek8IBCpvKggWHRSgpZq5E5Qy+sz4r0Httx00mwv4MxqOdk3ILy
tI7veDGPHXLBZ0Il43l68DBJvbdjvL8N/nTju+NjvQdKKhI3/KiDSqJppcwQQbvY
BLqQsMr7p/2aNQ8jDzBGisK+KmkOvGZtVPosIZ//4MZuJKoh0G77lJ5YOyelGxv8
fVgB7vDR7xz4yV4G6KhiugY2DqA9Xa6s4eAR0alYsslSDzdIUXzTHcIkSOHL2+sg
HnvmJMXbbzJfRBKjUE/PzL+L50ODczTVTeWsQJcocO9oT1yoxi5wP4EQGR4Y15sH
Wke8nFbeEnz+vSWb6w6kX5xBy9w74z56aE5oj5xxIaOOinw7QmkOfR6fss+vzURh
ax4faQSh4Byuw1I7/6SXp+hUB9IFx7a2y4n2SSZoyQgCJaxkE8QfRyDpEEm3RDux
9ur4/rIDkJMXZ/V30qbz+nFOoCY4lZpetinECYg8S1XWbB6GL/zGLAWrOqjIKy/m
u9xtIZQxjL19bOTfyQNoFixWMwI/CSOEyjJKIlhSW3BniTJ6MmfTatbosVJcTME7
f1C+vw4J82qjkIB98qUnBOPY3P9bx69DiTd/eSXjgm441I7+pteVMQF/BTwZJP3e
s/RoO3Qp3gTd13ANq7VzrFztMJwIRHjgMmV6+l7SR9+dMvb9FkU65ogTpgqHedcv
z17E3o+DlJsXErCZAljnumcN46dBe1LvXUqinvWaYh4YSpB4WslGhak/2xFvArPs
bhD+od35tPKGUl2315nBz17iRjE3GG8jEhSjzVb++8DfLll8UH2uCcTVopkXDrcB
bS7yteSDa8FA7glnQgsxLKFlR20oS7dQV/gUvfgVyUttxZihdrtAzFWNoVuKvraA
L5vJwf5piIWNbeio91qtGz7tWJi76Q4ESi037GPjJhQtaAIrFGXquSink8+64vhQ
4WxN8ATQu+KLkFtUyRj6mR+YLs8atOBv0wFi4OK5jnYzL3XBn+l4VYf4jlQ5+Uma
xvLseDq2mp5MU1Iy+Om6ED+N3uvh643z0USyujfTQYOGNxtXtAQSaQZ3eyqSfj7r
4dNPrqCP7/cLR7wQDUX6H2nrx9ukOBcTsiXabqEV+NS0JnVrC+BezRyE9EBieKox
tNprkXXV42TwXbKi4MUQslXpd3bmOX9KAyvZwXKEkvCa7t8Lc8A4Oj6L7LhbbBSH
PKCLedsKcfTvG3mssj848cLkYdNyfpsTm+rIW/cyQgtRqLy5bfe1yywkToHcLJuH
Fmc8uadEDDDXtHqNZYOoV8FPYua1mVwEiuw5R8ui0+I4ryRTiXg/TOBL1znHO+50
SyEOOHGqdbghNhdBL66GEHJGmDZUGxwE3laeVKkcmKkqT1pcdCGAu7VyLCoHXos9
Cw/+4wXsAbz7gZTLx8jqDJ+2Ee7Z/rLj/hzEEqU1uIt7H3LaM7i424+1jeOWswHZ
`protect end_protected
