-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
M8kNbi2LeMhIglieCoud9G7TMQSfr/fpPshOtmbks/9wC/ma0RoA/16F7Y7TVEwoZsGrYwDcCQIa
YLBa2+awBkGxM9LR48qExu06q182uG26+A6qW7iVnKFb03cai9gNJonlH+giUDCTb7wdpW/EvDij
5VScC+S+rUzGl6CtBgshIhO4rj22Ds8kQtZSIO3CBW5R6S5pisxTLVHwA0qBno5r0tR+ISS2N/pp
Cc6b7hpX3LchmW3UVZQKX8E0WrpcDtVtzWWVKib7KXD8gOWJisPcie/NMxRT7LnGwDQpm0S1ljPw
JX+1Q/hm1xTE5hmsV+JCJTE2gLMYWBhkha3QcA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49792)
`protect data_block
L4zztPJK1PaC++YD8RiFJuy7owDvRG6E1JCFDPE+IkEP04zwqd6w7hT1yj1yOY3Wddv9JT2n3pJj
NQ0mZDQnDwR/sdGQEmrtz/8iuVXR6ZAq7YhBVXN3FzmDWlRvp/iNmF6lw1dRQV/2j7WMi9FQef5S
q9uPhM2bO/dBMeZA0leggQm9QtXnIAwKo19FqaW4KdKIuhJV5FejR+uMH4m26d27fLXT44UxSoUG
r3ztc9uYaBzhZHATKhhIFyCEXfkMew3Md16OGPQ1lHP607QH6/Igtk0rg4Yntc0xAYIwJoGknsRt
nhEiIWpDda83NdJfoYtHX3zOFiGGC22K3ZsqiGyuaWSpTc3t/Vb6hRfJIJYuGMwkRK1N7ECpyEL2
ID9yUHujOGMYucMSgUssBG/FBMeVi7poIDDBuduO5ZCjYi72koi8MTo3AhoShfg9wlef26Tp+Uj7
1NKDKyLxKvanfW/lLflKpVL4hSA2UeV4yPAaFcj+on0j2qzvKbVQPhy7VAA+x2j3L5nMZvjI+1ly
iAjgQIcW3uYihS+ITQ7sWs+tKaDn1eA4rKouVaKlun51c17CaQ22RY6MqjgRHlhyBnDOq77BjrXX
/olKTSu22/mKVLOBh5JKmrcQxSsUC9glE6uYEToZL/JcKyYBR+p05vtvxv5n8Y95CJv750PL8z9t
ifvCFzBx0GIn4pDititHmQU2gZY4QgSd1xK+yZUgXz1il1tXhOFisusmxYymZPSHRc2LzC/ZOtev
6awc3YB8ORja6YdwsKsr5FKwF/L+OF41B6HFK2cCMPTlP0LL0LJEKXRqdR/cC2h55mgAH7JOn4bQ
RJvMCDiQZMsG2bZxOQ51ryqa1naxpxD1v+ha2yC1wjacxF5rOZxEDv9AzxR0q7BgCt6088TemEns
kPVr52yELCzDJa5znFRMTPVza0BchqdEaYnku6DL9+jH/Azwh+CkIxOArfDeHbUVy0zpCYEfkH95
9PpQfOVjsSoNXbZcgMh4cF6xo4gwVXAUahOgX0Phgv+v7OunOMzisvreO400wRjyixWLsdOby7Te
1+JbVwkO1Eb98n9GWdBiaqWltkRsigt72CFqYuSm2XoulTS2B5+l6BH18MOjcZqN6uUZpHL0F/A8
Z8Ek5K0y2h8d0xUEDNRJAIWqv3BXIhUvl3/a2ExRFhbdWvVZFo7dIBU5fBNIGcIgDaotFOeTkRVf
KP+ZE97wHt70sCI40M/XOAi1XJ2G+Y1+Q78IbRvEmmFu72dhKvU1UxGRShp75S/KmzEh8MO+Lkea
TvQDePAHlznORGrvvfIcY7L+MK0oCBKYId+5sfi57IIS5jmP9iL8Pdm/oINZ+PKY2eq5Xzf7SCeK
ECEE2T6orsfumLnp3t6lk9F1TeI3jo5DPiegZI/76/kOuFueTmR2+8uuyBvxEbXoDehLxoZs8dzQ
OSqnS79QVoq23ScUf8fhEzzy7Ebj8wCxRGlu3GtChRGnssEGDYN2FTxzmoqJcMOZ3nvMppL9hq/W
qWJOGUk/zJaQGW2Y3diWEdG2XWCCzjhQABRdxZJ4hQk6eHOXmaWacIDwh9M11p6PRoNDB+jllFUt
I6WqUsx1x/1lT1wBV22HbW2EN1O8qQ4uuaYtOErRBizoCV9axbEZI1S51behTLClY86W5DWF6cNa
PzC9y1naeJK5Nm4Z7C0dij+5Pjk9hJSdoK3A5HqBVB5+5NNhha4uxGc9M7t/iYK+h0qv7cCnvmTL
JDpgCDMgjnS3H6JoPSGO9uAGtxYjMc10/AmAl6KF9RJdg2BsUuU32iAnhcBQHWV3Id3Zzbh2tBvS
JQZoOu5oJ8/n0b0lBdYlVLjdvLnxurVBaRvIc1IeSWnmATd3jX/ixI9MHn4TXp3/h/5U1OMT9DRj
xFvI1nM9MOVOwOA/e2Z03UAwQ4V/4v3HPOt0X+Fjzwc/b7havObBfmqySYLD//cm+UWZjBibfTO9
xLN08rv20bGRfQKaywkwV4vTTIvp31YeUpxLjwxYX4IqOd8rEpnOsNNnSiw6tnRw04h2VS4QFgM0
8QZKmJgAm/5gEYJa+hRG2Su6vmqiixApmaSqlB68XOV74mGBlq9fa1vYj8YlPVN5wnb9iaRroKdQ
aa2sEOFbNm1hg0M53/DFSq8cgNi6MlRQvosoNdjVqF63Vgp2q7sMEG0OBabRMXEIchmpTwEF3oem
Mj34WjTAC8RLWZo+2Qq1Mtuw6bf5qdRtUvv7kL6uLvayBICFnrioT9XXgYMEu2TDkqw/IgXNmb04
LkuxWWlBZLL/8CSIxX8f2rkPBghk/KRsEvMEeZNJBrVmYYtYYmMCTyugjiL53/GZ93fUZHskuV3c
635tglj0NtvrJKH3BnB4ehB+UyHXN4S7dtNEXAhmKZPjHLLWEZvPd4XyJo71fvlacNqddpiqeQqA
pjyDAtz9EZCXiDJ3x5/n0U6EWOI3Nal2hfipgKK2h02B554uAYKLvkc5Z3Zgx1wKpB89IIPFdsGB
XEjmgs6irlgZGqedUj45Bsy+4aHg9CxlkmGYzjjCkWNGc6xThVtoUNv1L8qtm+17+cTN9/ksahEj
ld3Oh40vaQo47HvYBed/P+Ocuw5C8aGoHkVVBsdhZI4Ap/5CjtC22u3Euq6biw+WNIqeC6DoymIT
c2fkyfSi4bbkqMsPJIBOc+MGhw/FA6ZDLyUisz1+BjVsooVGuFMpO1melW8AlgaKTb3ZBEgOO+r/
f33FM6ipL3MUPGZTANkJy+7YScAEkLNb2EUUsss+i8jA4hP9Dbgu0gwoNvwqtGvPd82HMz/ej73k
qLo4Xc/4TbSAaypGNZB3UvsNu5zfOxONuBlSNpV+x9LAULNYkTVTyVr3Ju1kY0EGK6MGkApN+ybC
qDhxCouPe6IfbJ3NyRgHVCYCD5lzaxVS4/9yKCfS1VsY+aS/2kBpIDfJedN4l6X0KysPVFu7frv3
BZ//GZGlVV4B9mIJ5PqlGMAqaFbk3dfENhnLH5jIBVq+t50eXOAn2AQAMEGfzECGcPo6XjRNchDn
wfwyqzxkRQbuGkx1rXRlJeMw+ftTwAexQS2BeQiIszUIsDDRmJr0XbyvKmrJpXz0mAtlQFMJFzVT
tbRjIpc9+2fUPUjSSogJb+xglqMc/4mE4U/fJ7DJq3MCu2PoDiU9MaiCiEtYvQwj41ojeLmmp31m
SARedE8J75ceGfF22q0UZObA7FWcSsc+3CAXkiBqaAXI53vqhRXSpUxfC62cBrJnDTltluRd8132
fY4Q6MYCkLpXsWLwIkgx8Z6w7AyFcDDs7l4XePmejowNL+x88KNMsQ8BLiXR2g1qPU0E/A6fPcge
SSeEQ8NQWLTroJSTtwdizUZPZiS9afSKcUkCqzD5sg+sGFYnhJ4tI5mUr7iIqubklhy4BcHZoFiY
M56tHHHDVoXi12/0fcaWoL9x6Z7nOWd4/Zj+OdGUtyYday9MYO1xKDIDrQRnlVdRc/TB9kABpEPK
4Sek5ek2OHeKI2J3ReEMy8CAhuYBNcLFSZUn7lEUVQPEUPyu4pVn5M5vUcQf7CVWr/E8eN0hw0Wk
UxRayuvuUn0NzdxVbsl3CvogZktKCc+qH7ZvPcbtE1BGQ0/S7c/HchJmRXgoQMoBKnr2mk5c0quk
jrq513exg3jJxArObJWuq4OzpxDupNhLDQmqie0WU/ys6Th5GJfR251uJB1BZf0SWlw8KiALSj2d
uXuQ97qARAWr8AINj13dzket6AO/bBpK3CLYseGCJ3jP4a95FEsz8e3PdUnGvYh0E6Fl2Ja2oGc6
/jQqdovJaGWJ1QKgduxb8bOqgLgWoeyUEFl2w20t4oL0/2g9E306/1KUFBJGg2vqQCi1VYJHyapr
5YJSlgCpJdSoG5cKO/S1EWdowuMi+N59GJZkrrMXgR/WrjsvuERr320tRiZ5mcelNhcGGl4OHihp
f7a7odJtZYFqYQlRkD4m1iAuZodSA1H1yyytMZmGHD1w8TWIs4Wlq84gSDHhIaQaCntdlNYew83T
UsCR9eDEUvImoJUk7WoClZVTXTiKt5JGxyGGpyPirqomsz0W+ihfNpoG1tXTIVLJaWVyMOvLwWoJ
0achqRf+y88M9whuqbDp67GuZQKh0fBG2lyNf/a/QemmZM/W4tRnGsuMXioPC7WZSYo4oiYitJuE
LxaiVuUxQcmCS2eE4/imbtb1TBFc71gm94QHjqAg7X56iWbvnXBmw++M9AXTdVH5Q3BXQs1xtCY1
RhHTPkqt24Scd6tpnzt7/z3f8C9+4Fdb9zHe0wf8u0XAJrkGgdY8Vu18PE4Gb+p1ACOjkFWyb2g8
R8lsnReL/K1Y8h/xP52ZRBvAF9DVJoB3ITj6TOgG1rtaCb9m0v6I8yxjTfOKEZtAyJ+6DGoLC7Ex
Y5TRvkjLKxpq0sLDSQo2NJa22fk+xmalfhL1Sy4BeorNVvgiR+3Z6lyjySA+sZHpk421SWWyG1Zx
eblk666fRQyWL5IlVWBh3qHT2xIsYL9Uv57jUWwPIBFbTm+36JEVQGnq++2UdAILEad0wlXY0mj2
1cNQO2+dHHgbRLYQsYb3zA725BqLL23PxXMgfLNBJxmrzxHFzjoTDJDutQq3cPZZFoDGAuTKzE8G
ZiaAiJ3aelz2b+WcnvJhQZ9EyvJmGVeuI3IFDFM/d++JXHgIhjXW+q0ijx+jLullH+GPOhRg4dsY
zW30coaaJATU4j9TTjPIlQdQog112gWgy6/oxNh1Er3ODlOg5IDXtMm3KSjzB/H14u9e+g/F4wAQ
BEx7HNDl6753DZB5Hnk9ucnY2HG4kgg3tHOfFv5dvs9UAepriNgGL5Boo0ktD3OaEGKZphpVlzT1
MXfD3yDX4lUhnNVQuabStZjPMOE+giz0XJiaVSxUq0AqfT7WecmG6sMxj17POHFAyhfgc8bo+3LW
NtaGAV185M5SB1FnnAWmu3qkjU9XTfoWE/LuI5knrwWOv05Qi7cJqIvLRO5s1kBvFRwJvni9qmd0
dxfTXmuCSRXlKmUDyfW6X/c0YR7HaTWcjvfr+vmYCSUFpdxvLmuvFnHSr7q5COV2KmC48KtXfzYn
e/qGo8kjRh1Pkj2xBuBpbl1d/qXdAwIXWti0yGahG0LKXuVVXo6dgocVmGXHVuapt9loOaK47e3x
NB0S7bjEqns8vo1+MnUmodkyNhohz5WPTgHKbrLw49qrqHj34cmerz4R7ZkvZvSR1TUTrsVk/9tl
gr+B1AL/O+G+FUhmN1o40Mmrz8MmWOiEoJJiOFMWJJ6Wd6DNjUJigkYz4CYl03bYVOM9gRlxATwt
A9iaO21/QNdBMuDIFOdQhKucLSLR1l6hgzouELhhe39d4fP0Chb0vxVnwI9lBl3/6e0FirnMYzU2
LpwU89MeCROJfGkzpSTuifOyIMvDGjbShP3MquhQ3aPlf53D9FMp77tCu2mIl9VWS8te4NLBO6DV
KTaS9wxMoi7w9MUDKb4T6ekUI7hVcxkX+0z8PaK0FROjWOK3RbRuap/Ezz3ulPdr2/Hz4P1TfGvx
rh7Uqw4Q0xNtLNsDGbNHzLZcP1fzj7FYJ9JqOlNHkQU/WunzFCDqOce6MoeFAWDUNPU7T1ier0dY
2JVNh3nzECWA9YmxxNWAkBFzaiX3WT25WK+HiNxtRxdKS7iF+hVCMchZt+RIM6QKj6RuhByAAPXP
q5Sv8YqWajWbEJzQlMbq00gKDPiJ/uI3n+zdSvCW/prJ6RD6roJe7cOTGEGOs+6lV/2XKtILzUfQ
QpPEUF4YdXKU90z241kwjrhAIrgwtZ5d+WMxMmBhObUx4AB+kEJjUZNiHk34IUGoD3+AKVmFoOHF
5Pir9F65ZsF6pn6C4eyMB9G18lXTCPglH/E+ILVTX1RunkRdHAW0t4bxpzKZaMqwnGUSV23RaGiR
r9Vs7Lgw/h42nd4o0QDnXjxFoPQVCL5mGtBbiHdIhSxlC5fsssobBMKwwDxSrMNT2jvH6CfJJBNN
FszKiG97oXIxV05Nr3JFN7YcLGsBZGFFUO5iQH/hzAoGJFMcRhKSLt/AUebGtxw/cN2dCo9p4Gyr
+5L9+nQ5ERS96igmSBVbW0wilaVXAB74xo5GYBGma3IrKeKtaLRLZkSxSvziXQldX6igskd9r77t
/OQpkrCOpGmEJKk+3zaKwW8Qx/g5/y5m8/vDFMNmKxFULXwpGTXyWgxd4Dddi7dDf9m5ie1UkmP4
UZhWuPiITFPo4Ps+HJ8mdKpPvjCJQ5vpFHmbRs0Ymp4hYr9Hnn/p+Ji6v0y3nvsfZ9cVd1UUrtbP
x7QLlk2setL910G/UcJBy4hUyn2iFnHN736tbve6YFvqGJLJ1jMJBbYvdA5mzY8IxCvCmsooTc+K
X7n+QOUmyk3lznu3NOUmgPUSqL4YwNAq7Gc2xY3j5ktsAJI084uoP3oyMSPb5sef/3DdozOBCcVd
lqY9zCVHoOqSe2R1ofOpTNqa3DZWwzlVrEmG1anDVOeA8LTLT9NEnxQQszxP9kkk+FoA7GvrL1hp
wDVHoWV+4doXghtR2BgFVGuxm4z+wdKb4e9Y/1gjE3s7qGjtWBb8G4PBBBrXtaLb8SxkxyjzzwvI
ohKrw8//iXFcmPJauslGAaB5GsH/XuFSX7yLuiYI6DxOzt6pDMiVP1IMqW1yZmyxNGnR87HFKAvl
K+VnuM+7Qf4dpMGo2m8cRE5A4n4CKFpFg/espadpS50SC7m4D+Y1/s+o8mFlGtOUZvs6u2hBcT0m
ezR8zHIdcodaruiHRhzrFDrmXvg8mmCELabQviYxHpa/x16dvHZMM+PCwrIhTpOV0yfUzrMeDYZN
4ekDT2anf3feTvqS/SH/CoDpA6iZ6VldDhGtY9+9WfIJ6ehfv/DfwWm0t5k7JDrzWrw/LeNqzsa9
0bDkJZhnwXvMwcdWG2pwsLkC66HLrdHVYAGWcxlShfBhriM4iVxuEW7gHz/YfZh+iAGeonLKkN/F
JVKzt7U/pwdokwj6+IHLzxDANKo8fjTurhZ7SYqX69dyYbnTZTwGAhRnIV9zD2+u+Of0Ir/JAvtd
7XxZxXQKMmLrLpNrEJjYakHbjhxVD8IJwzQ1vstJ5DdLK7sGmBn89bWs7fye1QJGyI4g6b+qMWi/
wQ+DoAipWI5Pp2TPlb28EtYNRGwaabnBVypKHw5VSAGi0s5BJq/gpgW4Fm6FLOpjWx4mpgKolN+i
WjANVNcRcgZleGpJOaAiUbKXLj7ARqm0v1guRCctLqgO6pL1q4c6a8+vdJNlB4Q2SzfK5C4VoZTE
OwW5t7A5OMi3ETckuFns1TQ3747SrxPf5k3IMZf4L/+yAswpXBbMQLEDL6D5Be/4UoP6eAPoJUPb
Bub9r3cAjijHk7RTLRQckXv0Ulylnsm5tHAtBXhfPrAk1xI4DwCimiWcWDIUy/CUYvEXqZwkrrxf
U0RU+ue4uvPwYCbgX7Z9R4df0k8BzofrRYZGx94TIBPwrNGCfBfoJT+/z0cuxsPpiv+ZclguBQiH
HX2bZHs+nEUipscEPDCuZ6OJ1bYdwh3x8pK5SB8qdUhQkOKaEjNO65SmWDio7GYWj5hkwuCrVcD/
PRZMM5pWiVfVuKlUaQ3LSEjfPznXlYJuBX3AiNiuOFVcEH5FpdTAnb2dd+5+RZ/Go5gfB4rVgDt7
Zfj7X2XtuLBFxM2gH7+SEhBtIoZNaIOnCJW20XP78uWybsMvDYPG/g4/zcB2JYhXWEL97Ibi3cMs
vxot10CdM3FXoVddW+0onldNiUwWbqSWsYK6iDL+Ym56s4ikWn01jNN3EyRnPTanl+fPNZ+/WwEm
C0RdF2AV1kvWNV28mFXTMLmCdj0ApscC6uMIfYX6ImNJzy8xlGye6b9cnUGR3rKVbsNwyWBHtTFX
5P8W7Bskt1MnfaWFm0AZVjln0F9OPPGVMDbEh/n2K+xYHB0vQoSD4TeAqzfza7WJNk2YHGlghOS+
Qf/TsjndwltkhfCO0RoUmvGcn5gLI3h0iFUJFF9p34BfX98awdIHh73Q10Z+Qezg6CkecIkWjqiG
ouasD+Y9KN6GKIm18yLK7mQ/z9pMMTgCfr9WC0oR/nPzDKaG9KL0Fxu+PqI7wKxPb8tq+7qlibhH
Q1eNqZEMxJVBel41JM8lAqQwQZQEp87T4KlxVWzOMFcjTVnV2F1jmWlbYPOhnGrY1flR3EYTmM64
mGojDzA0M08g+apqEtQzQ2ygRQaJO2iTV+mwW5ndEJDSL2HYoQnB+zTY4H9G9thYm78wfLq1EMlq
pHqalHLXyQ+Eum0Zs2HANFKO3QJh1QJ50r+bCgqP/kPgSmHH7cQrlQg6kit+B87w0g96DsYKSZnn
O+FRgLsG2dlFdcl4dU52/Ycb56/b7dY0Qdgf5tyex5zH4NhNz/ZxvBHsEex9C4KW5fd+toKHZ03p
35PmfZKDnBlNA/S72im/nmel7LU6DvwRaIHRp10Dk0+pwLrUcyx9MT8c00dDXhdFPNulN+IJJK+9
s3EZgKYJ2jV5K3rK228qW5J1ex7MiDtXINf+vMlpkfVPhZG/2KDTuOH8sc1AFtkNfmMLcqckwM+f
qow5+H5aSkyCgqSwSxZPLhCWWDTC7OIcKZJFMXMkMrHffEPgn8wWmEFjAGDFcqwPTEo+e1XN5A9O
dAWEav59d/NNBAzvDP7g9FxnZ7HgIKgl0E0Z1kpEeNIj/uKDI0OCYdgo81NBdXfV43j/wSG5mZCp
fQSQcPkZKLl2a4cUqr/dFD3sAdvxP56to/fwTUhA2W3xaEKGFO5WxcQSsIQVIDRRMO1LtuxuPeSV
GhDPvQOupO3BpxFJanUE7a/s/WBi2UGxE/Jcevh23DRf1CHFJHVSOttrgiOxjlK8tOexywZPLcX9
2ws9XENbJtmj8MF+LQgorANm9a0Ihj6WtAKXo0agAD7lqmt/SC0ItMtlXr0Xxrxy097D6rtC87iz
eFnAOsKXvTUNxE+GNI0c+z2m92nRa5RbiMY+ySQUvcGjXDnVkpsvxYVtqqI4oTIAnD59V2QJ+QCe
4I5P7/2XKzfVN8IdgLrosjgTP4D6a0s/BrSMtG3vbXv/uFeTy3Nuf6w3rAdOy+Cq/LS86cbfqPrY
Y8XjIF/2T1mlaMeCWPcP9HLMrHAfLzFElYjU47QuF0DhXZcQGYwZnSAjdQmEaTKcawIdEtn/v8MQ
AuzZUJj7PNP+zJ2+LuohMAFc2kymIXZQUU3VTvYBg1wauhVzX0TfZGPwWqY1gorxfDPf8zLLIRjz
4mAFPDE3kjh0JbVK5BG79kzhKOn0VpjTcP01RRGbjW1FAVYMQTmtaYEQJF8MmyBd9n6FfdMdD0Uu
d7k6RO6ng0GIIw5SaW5bkya1sdBIyf11ovtL42AjIU4Lzl3uJ5VzuCbg8kCWBgyFrkyM0e5vAPwe
R9ScQgmhIzFn8HLD3+SI/DNqrlWgpy74B2KFgQiJ8ypq2O2UHuVbhw7cW75svAlQVrw3WNojkCG2
ArXzbhcpOdR0IMJIlw1MWHhtr4EsznHSggp7DN/pk4K+bn8Zf7C5VkvMrEkSvlfkzFpOwkZbxtEy
u2i+NX0z7dsf2RKJYYnu7ykqVxQgyXbrggk48OMnJHMnuSuKeqet63TcJAgUkZsFD2sB0+ybkWmk
PQh5x96vAIi5KBfShwKSs2OZ66igG2fZLeNvZsC2JfIFDD6xzqkS8sJ4tCIvfAgRBy4pTci2q+im
3Mq8n4SKS/OEw7JKeq4r5oxyjpdw+1izGUG1bWIaDWSzmD6bjWUAYi7OcYUhZV2PgidVh/dc/o02
xcZ+9vNT+TntX/6eie/5pOqkC395huV4nlhY/ts2IfahGhYwmH4mg95hqVyolRgnURieVAH1lQnN
AmvsRD8ZirNA0PzRrPFDKDtlaZmvrsQnNFwXwwBO7W7A8lU3L4Z07EGnTdQAHcYzGFfHEiGSdnBH
Oa07L19dOYl2i4lvVoOEh/Xat1EWiWz3Elxdxxajv22Tpf/9W3fZyFzOq6diroOUUEceLRjCeEkG
3pLRJTguiDsffgOyhuG1Z6A5G/CVHf6H6Akek+okihNiw5pWp6rv4utTb7oH2+rVKKsK0WJtp47e
7Ju4AwZKdfRmmtcmx/VnYkHWknxPt+N3dcdxYDFO6Gp9iCYmySLK7DnvgPOQkG2Gixx4i6Ds6CKJ
EFSFaKF0RnjUJ12Wct9SmoUmfUUcgMXqHS+BO7Yw9NEtwbUAWTaY37mxfWAmF40Wr30QbTy687wm
T69aJLU934dKNEK0TIZuxfSfUsZ6Ip9s2xN+a67R6MdQf3/KGWRvDx5vu7f3C4DNPVOVJ8+gBf3v
ixLKQONDlrcZzjAxNGqCTANxOyl9FDdvKEkbmZDWwYpOnFfSYhxrpt92Ac+HROzBwSJVJXrEFIZn
QfDd04nZJlyRCkqA13OP9OzD9yh4kFY1+dE92dkksxlLiMwe7DUru8TvhqGGb1y9vjvq567xE/TD
s/55prF94eP6twIeg1EbMAvWK35v/7FcFrlSt+55mYwHjqQNKqEslz2HS8BrT6BCcvMKTM2tzRIb
qflTvBONOSSYuThaJetcNtn9I6pxQifCzoh8Fxn6J5XAVVc5S3b11gI5+Cv+GpSQl6mV1egxf8tn
olypKGSseRHXI9HSB25z24WDtG12r/G5xoXeV6+8hKtE4hWl0/C3rxalssL1ETwtSkNo2fVplGPg
vcVTbPcnsUCHblmBxUDyAXZpmTYRm6OCf9zR/qsOnBs1LPu1WO8Oi+Jb4JxAb+ryF2ymqA4LlNES
F3wpEhjt+t40pRvGQuVWW3k9rAPabKDaxpZxKByLcLP3rD2ZRZbWpMEOUHkri7bjwcL7Uol1NtDU
gOGNcl+ScfAsSnp39Ci54NDCQLQH7wXMMhFOqhscenG2vO6CYxONwsUgcYJYpIi+kgPVV2DZ8Qm3
YHsxQNznzbp2eTAExa3pDartAyvIH8XEnc3mFm5Ik+izafh3MhFka1Q7qwBibrFlX2Kfc44s02c6
5v+un+KT3o3YBVA2NpxodbQ2VpU9zEcUldFJt1p2kkB7XIPxnCiqCmFvvte/VUfF124XtA8MT+dH
vDh2UXPIdwfB710wezgrUKv6Gi6wWvhAjBLiYxpOVce9HwB3Ejk1HYY3VtHrQNR/1UTYmK1xQxni
xynypnYts2xhwqZmrcxlHD/jkJVtnuEg+UaFRioPFrATuE3e5Jrg+18EaLLO+gnWtn6VGpKai2hw
8/rpvxzyclazrjdbjhtLAxvyOQFPbLWJpntiun5oXlP3FjDGcMz7pIbJHtK3A0hHXQZ/ikEHw4/k
/sG/v/38vSCfg0M5Db4+NFk+Np6guRBuNzUvzs8aQybPPNWewD3TQrRxSd7wPp2zCQ/B0Fqoy4wr
zbAhUVQDv6j2Prj6+hYw3HfILyqCQSI4VC+NZBjcHhjGzNPjpQJy01fDiC44qydIJuksop8vrCYv
Xs5ojKlqKZRzX8eWBdlZOXpY5uzbQ5h+DxCqfkGI3emwrZ6nXPaQh1HSt3oiqL1zi2Kqvd2kkg4Z
ipYx90mrtVkrf6nPEnuOZzn/GGn0BlvZ8aI4hCrxfgREkkZZxxDTWzVtoUxNc54sFKhxS8w7UBiS
kJiRSVTcq4E10VK5UDLXsQpWA1SzukbK5sJX/homutlFfWPzvg7ZtNSpx6IrRtMgPQH6fIncOvl/
koGA9/0eSNpX30i8UeJ14qTiEfcvu5RyJnLwH3z7eEpZP3zbvxmZMFtlasnC3nsyIicQGBkWGnoW
rEpu9h7L9e0uVcXytMJJyod70UK58gEsjIt/ck533VOR9zEEgK9+rhTaeAZVLbZn9Qt2Tx6TM8di
3HKV2cPrmr+U/AqQJBx0V/AbW/7DrWEcw7Wf/y+ROONTPUEox9c7c+flNz7m+AXSU5F31BC2v7oS
s8e5T+4XwC+37r0E/9UVfTYEnrSzweIG7k5LSlvkj6PXo8vCy6w8ttqhDmGfrAMnUV9BVP8xs5Dq
5loKQmyVlYmI9Q8K73WIUzuZ8QTlJ3G3mpYOq+RXG8RMEK6PniWVDo9uGoAafRWvwIbOXI4BfmIj
22Jy5tVTADi1bmtdAktoNIjgzQXvYIClnHINAvX9d9nLZXuq86KNvMcxjeEcVO3y1GCsZUmJVle4
vBKc57tx0qkKRLwtMPYlwo7ynBXIzD/jkyQZ3x9u+MctnSGPGjRQvFgVNY++6GAMeq7bTxZF1q9V
qYZZv1sH9FnKdF079CsiSpl42pEyTjSpBwaWcnxkaODo19XMSAXimTzfGBJaF/QnaqzdSLwEgsHi
r3k2DsWtiP3nilyu9GT2vNxXA5rSrfjfPNFlLh+yA73fZVf+imRCS3BRfk5awxTeisyf2ogpurk7
kw52KX10amwUyBh4f9sefS4/dIEVRmNoYDh4gBPc9OoXByZ1Un5I3/IBHmETi1QC0js5vOCacSSy
cFHsTQ8HbCucgizR2RuG5Wk8s/qWTZTVrp3ptotyOOd8qHuYDR9nVG/b+o5Z4neVdjlFd+zT1TeX
pfOnktbespbxNrpKi00x1oD5tbYRra9/JKeWErsMDyvmzLN8ZPLyDcNOhylawIIa6MTKru8gX4WK
j+mq0rQwVgYXOcyQgGVeIqJGAumhkefa3QX0BU1vX2Ea7CI+GD4fjNqkZ8zBKaBUMsslbMiZunjz
yad5Tb/rPi4dM3lRcYPpiTt6ISk+rEQmTtlvkJtrzxnXaqJR5hWKrdNfUYoIjuPw6JfVagPt+s8X
KCtWFWjFgcd0VkjodPVlBqVuJCLe+pE4G6SMNrBElq1Y1/Zb2zWNZjbkVsQ56tIUoeUxeRbRBk5v
/aYrsu0YPTG5c8UqwybSK4lo/J0Jqh8tusbBGxnc4l34ekPPVss0Vl/+XE8I3h+MbbSQpanKSQZq
/gDoK4AvmJQjVzduCbMdtWVKJhnFRZiFx//NAyMEKH4mdIsOOLZN+0VfrmrwBRQtJvGU1RFPggae
zjN3j0BaKUZf42KLc5gZ/NKVthCNI3P0fkBkmB4NRU0emFsZgWTZYSDLX6OC2n7a1ONOQBfqPgwx
5xeAeUPEUAbaALY35WG9jmAQ989bZOO+Qjd2B+lxk4eycKcvCqG+IZJ2GDlz5D49jgPrhrw+GSRR
LzEhwPmGXgPW+wpqEcrQd4QeB+fw0zWeMHBeeqw9ZQRnTv2GA0j4Y2BTDtzsRrpUsT4TYlshoRCW
B6fIppdWSHrDqK+xk0MgCNLTa4h66SG+fv9RiyQTxdoLHYPsKs6ZajCJSEshi5INCzSE0tilqq+5
FOgy6Lx67qDE+1rXSqhcMoodI0PeAGv6mpFpRdcAkWF8K115V512VcAApS+34eEhg9YoQ64VnV4k
Jj6akJGyVo3pNibysdqenVimuigZYPFkLrLcVxajKJtHE5jh1TT7qAvfejivo15qCuQXaPGjX7Qk
VHVZHyndC5qHtIi9bz8FDjsx0/dMEYd4CVRnB93u8Yyn3KXQTaYJ3P38PyPJWLx/dV6upvj9PdMU
+h3OSTQRqTLLrnAmg9X7jYPl6xiO7TelNi5mwhzoMHu5EQTA4OVeK5WTUezg5GAOViHHV3udUwsO
YFTMkoM4rHiivHT9UlNgtZ+B4xyM/ohk2mBUG1vHohX+IdPaNxsUhycLoAacZzj/5S+MZU5vKFn9
XK4EEH6HJN6l9C30BjGlbMVKjD7JnlytrwoswnV8BaWFdF1U3z8It3nQKs7hrqnoohWvTjt5lx1P
+wkDynzGQ8r6cOPJStygHNVrJbl2Anuia9xYGmR7ZstNVEyiGg4vW02QacWsNf2ty/QHEeXakOHH
x1n5pbM1qv9y8JkpKp8My7OC2A/WMrMjjIroFKBhopHEqb+9kwdJF0iHk8oTNNwCDN2cIUL13HIf
0qonZ0Iri/HwpLfDcF7n4Bz2mThiJ2NkvvG9l1a+qx1dilC8pxoFeNLxREoSmSuszZDtm0Gg9G1X
mLU2mTfp62zj4BK86SgG+fY37PC7xv6ePyxEeCtv4PAB7Fbwup5VYDBYpvPnHu+q0eHj6V86U3k1
V4xvZ2tQrWwsTBkFqC5yOs5bmrMT7F5jZyT5BKu9RpebCpNy5pJ2tKFll6nzsRKSw1OmgC242xix
mCOGozjpsPohYZjyR02hw1MruODS93xjBLGYLM1ImVGrCxJ0Ao972EY1AN0a4hpwfbCEGYl0wPXd
F3RotHKGQQThzOHERRZeSiIm5VbF+3UpQO/jWKbI0bBVfIikIYKMeqpWam1EqM5gHwDqQ1g3dr81
55vfqn/p3F37tYzyJp7gSHpg3K7WfWnn1IYe8eautluw1+LcbJHI8YMGsiZke1Wcg/EBsncAh+Ks
hTiEiRfB2Wlm6gDMJHu4vOLKzcm73ovTaJOV1v9PwedLYcrYJ2XtEGMQ5JOgLhIlx47e1Wnh8jkV
apqMJDwS73bchUWTBT+0fJS+F8q4X81qTQG6kP0ooAZItJz8pFCfrmxznnC4ClD1jfQJgCeUKLjf
qkxzSjePoMuYc4BQdLJrqJ8zit8yBlSO7AFIQQidb20TiZYma5z03Uyc+jjJQpc7paeF+bNv5XYb
PYKr2jY9XHtr9G10VpMn/muEWFsx0HXqQJTrV1VEma1b3k8rxnGSc6Vzy+CfRJ0hMQvjTcbgGkgp
ClfI/ffTxY6UO3nkkarWPl4905Y230aWtzpEk5TqJPL1rMUARGQV0fqSN/ROIEfvZrte6oWevdIt
IOZgewYRRlc8Piqz8rmb8TFSEq4muiftQEtLz+ywlkzXrObBpqgp12bE73sM9E9HzTnH+RHZyc0P
taCcDjJrYxJp8YmJeb0dN5ZmQV4HiDUORAdAJdgQ4+CzhHddbBpcTizA0zQxlu4VXc2vpfzIr1uR
Gsd4B9WDQRMQxaA9GfS7RZEws1niG/ekP6L7OmNgwWjOzAX8S1U3hbr+e67zEoKFclQcBft5+S6i
5tsKkaPru35rZ6jHCMM5X5bK79NXcR8uApHszJrAPkrH/bBl7W8P2bqVP0RddL5UgHKsbNzmyafZ
5BhGXT3+2sqspj4ucDc0z12rHmd6m19adhYBrlSD3eMyEGbljR0F5qsaBvaeqUa61gva2MpbLd2i
MBl5J5VvQbNI6ArX7EV1ygou9bigC0f5cYX0oWN7YuTYBW7xEVOx7hCLRj0ORxYyDeS65BR6k6jT
TJLRzSi10h6js7Rx5SwG1mf8G2lqC6iTTlNI4kTPmbN3rUDtfmkcl5lxYiPAGHiCzTfBiNicTqsI
or7dPJMfEfkL8KT/xNZq30erVvOfqewXiSFPz3VCvM4SpQwAs97n2Qo5T3uUt+ZB1xnPqKGX0vAk
ojdL86CDM8sAQl7xon3eSXpG9OW8cyI6xvxS8Ch0SMBDg3DnGQUL5KzlNq1mEnMWGTWU/48PTWjL
qVg9JuLR0cN/PoKGoLzJuTVsPls/eRiq30DX7sbP7U58BEy2hfBGnOjjefNl1p8K7h7kBRGQhPPW
EaNqlh9iRxDTyguJawlILax28mdh/qcYkaL/zVcT2YCFOavGRxOFCdrk06zlVy40MFX/nDLEu059
Bhu9o41vAtgHJnqu/jFDsTaUKvpkmymhmgpK6VvZ7ny4HgVNKmO5C2eUMIzuUreZ+7OFVosAKrvY
yYtHcayQw/xcfvUTuxZ5mOKJahdVZhjzU8XV6frXlassrGA6jREDC0h+pBkXNYHSpYl4WNjBlFS7
7F1/Q9opgIxyyTQpBy6eLUZEmfYjKWrGHh0vZ1d1/I70relYUcWoMQr4afpg39A2cCLmq6hH+1F8
3XNGiygA+6qWr0lsDfthZluyYDa9XER5xk1ockOH1fQeKPpiLETY39fjwuhLvkqLWU0dWgySrwPd
uUhn+OSlbQnpVIHyg6cxQsco2fCYE9cW32oRanopzU1gr7tlDu5XQKsQNtwHTe3kFvegorH/xXGT
AdGWgg9OeqnkzWOoHJ328OgAKsBtyEqxke7kcnPWvV0eyTNf8Jekkm7haCe9f7BQvJerrgl4VeWt
ZWGiaMNVB26XC3YkBzfRsCZWloZGSnD34ripjjNgrfkvewGgPb96QExJAqnjSnLPKgXG0YkvbbxN
+6jRmx7vxrtULPOhIP30vKMiQhi8faJhVX9Fu4mPfn4wDZpGe1CH6djjtH6b8T4+gVgBXqRGH0/w
DxFkS/SF+trIJDxhCUwPez3PkYkxmYB538dukVIYoIj8yM5P0FosTWnES3UVcwgzeiGBQyG9Bvqj
oi+rmRHkatXp/NSo+cCDwqTt2ntN+h34pu6KAgcRaC3KMp4ysbxP4xIRJxf3jVOPfFDJ/sv55cSM
TWRZFXWFcRzOPuzFkWaUFTnOKW4AAPUUHl/qZWI4jApMPlZ1BRSketMsmV1SN4r9V60KJJWGYW7T
/FE93v8nO527qWRlxGg5Nx7Mauvwq+oGeEEeTAvj4an6ROywujw7dJ05xK3IqRNe9sBH8QMVfzsx
vL1/KAzUJScnM2UUarNY+dnXUYBmi3E5ZaTrQs0Nuz5UBvKDhyLSa4LwBVzX1c7X/hY/6O6n5UqF
+eZNpT1BquSuH8sQ3/RRgggc4qoSjDhz9zDnMNfDtlKQCRv173ucchBq8jlfh1p8hCa/9HrMuhLC
FelivYO4nwJWQolXeRAk08hMN6+xjubQKnPjV3OVqLC1Bl6bjucjiCTwC96HBvPIEJ08g9zHKxiL
TseH/QLapd1MHEvdLajUUN1y9qEyS7el82dER79uDcRKRfEaeMArHoyGlQFSQH0DMqaBIYA5ZAi3
3R2WnAexu6xUJfch0YTqqj1w52u9uiWH7WGPMsWbwDhn7k/WbGnPcZxLB+slITs4+DHAWcVuHakg
fdYpuE6HaLUxvGt7bETVeby6Tf1EqaVoUR9XD0eWBuTdAFQpkZA3shI9K9Fd59gsEGAKOd4shJsv
U4YF8TM2zF0W9PBZ1QYlr1Bjfh/ywsGAPX5Zmd36nkzaoDMpzTrMgvl+DzOxJ0JSTYBRHQjh/yYi
NfMAU6mZ4PVD2SjNlsPE2DuVb1YkyPefcWNJII4h59ZCrmIw3d1ZzfSAimb+1iHib5M0Kl1au8mo
Pk/YdCr25I07ikL3uHZwwB8poYuJA8u1Ob+R9278DcPwp00vuph7wAumT5C6vyaoxI1mVLntuZfX
Mz0UZQ6HVrivUkkQyjLFNMGz/DFQxagY5bi9jcHgzJfeFE7uQ9BFRN+/IICqWgOEUzyX+0YJDSCA
OiuUhSnYiAFc4EZ6WSojdfG74zOJWdYyL6JK2qWVgIfVJt8NpQZ69599Oc/URyhvrxIYKhh/JXP8
Eb9wJ6168sLJ8z3t25AEWcW03+bEreS0J48UC1XciAM6bifqLzgvgSnWsdzo2Ece5/d4AwWLlizq
Zl3eTDEp8x294atHl6G4dwGqndXzeMjM24FD/mT+DywyHpWEWpBXCAXQ3unzixtQCwnZdpsGyXE4
MSJarGYMaxK34uZWMcx7L+WljAfmk/uVXxeQ3bmXsCS36R1ld+qsMnqrYg457W3svdTkUXhhabew
j1CgDPQ+bbhd5oBCfV0DF1n5LfEqwZAunDQIPfaRWjl/bXiGOWx9FF2RsgpnEQNmo4DChvwsi/0W
WsD4CtPAtuoFWCnIxU1GD/ChVI5zcRLoslYKRCtEoMX3U5kPH3HpXC6x/b3Gu6DU8b1t0c5juC1o
RHCX6fqZI72FLZyp+qB/OProHttYFL8jc/md65gQo6icI2uG74KrflyUzXzXy1gVjRlWyI01/iHn
s2UVFCLrcjlVUtQN0YDf0UD2Igcxuu0jlJmzZ4A4xn+Teo6lFDZJPeSLZTAP4A4oKCfUamGhe3ij
6ELlYrcCsBf415K6eMg02LOTwzsPiEG2cgEQltyqTfzpB1/6r8hedrHX9e0luWMZVt26FfqZkN9s
ETlXQYwPP0aSjRSvBFyeq//Na1i/SArOWVRv/7sULvVYEd6CKCe9IZwG+tMQWgwuOzB80aAMgSJc
mA4P2Jz5yM1Iw7zIRKnx72mA/KNp29zXO7N3u5uRWuZpJxAm/9uFSJm8zkIVNwNyo8z+Hp9WhbiC
iG2TsJD3hBnU6WX6VxLH4p5O2++7jQd7VvvNaUNaN9FPgEZbZHjsgIbc+rKhaBcAbSmMYqFYf2cd
pl07xS4o+w0fgjiozpnhOF2PTzr7/FLhI/SDuA9hCr9vLH3qdKOPqedv4A8hZliWqKWgwx4WhVIk
T+xYYCOVQ3sOOHaYsSGzP85m3sOvgMqDckxcXz1lyb2+EtGxRUrdcCEW5UGGinu6hNEIdRFkvIbG
zUQ6ZtB02vkwSiibfhf5Q08DuZXu6Vob8iNjmiqmuiNMzyg+cdcoz3xZYo3d1cf2FDK9wOB/laOk
oI+6nN02i82HgtwMF4RV5/5DuXnnL419RKt2bv5ybgU+1By1bU2xx4HPfgIwwct7k2QN/lWzah47
lrk98DHJiMmqiSLnvYwBRT+Y7Yq5zSIg/ACO72zQd9P8lE6O8mL31jBH6D+MGJ2YC0sXgxaf3sUG
QOnSRvECZ9Jdc5RWRWbQQXRFVkNUUmsnU3zGGTV/TGDrsT16OOXPEuN6l9l9CLXaGKLj7cjGpjkf
7Ai4AxI/Evta3q7+fQ0QDT14NH6ztXMwTm3oqpi2F+K7tf/sw9IDP0PwspiWoS7rW+vyx9oNMVao
hwhYP3/nrdrZELo/HIqKnCOLkenBcGGM74guHviXsm071fBca2HGAgJL0i6IdnOMvgC9e3NJqZ7h
KEzufWXd6H1ZMpqoeXjueNWhkYv1M22VJcCmOsShLo85wJmqm5Zmnrm6kv1jbQPYYfGxT4DLpghN
+765BPecztJyDCcQbW7aNHPQcbequ8vqunS/tKLa8QkzAicMQE01R4k/SZY2GZrrDNBqHfJFVsJ4
8pRFUlPNDDWQDJUHQToAXeIL2MQ1u1NLMcM58CDz3QW0X53u+2TTrilHUWLvj886QMmG3qiTu0H2
SoZwHJZO815N/U2rc5HlegYifoS/YqX/2MQQjBlncJtdXeXV5tALqgZDP+lNwkkHaIL3doIZHDU3
Z9ueIZFOoXyy46od39bkyztLDWhjDTB8yJel/J6xnBYqz+lXa3N1RUtaZZMgYer7FfFgELNoko5I
vaaQdy+Kex5oJDySQzyx+ww5AQ6XZehSFAsOXzXBb2XxbMb3O06ObX6pj3Bg+5yq778YL3OISk8U
ELp/x7NQ98AJZr7Ukk9RCpFC6Kp8hrXqUtaFUsY4cwr5RrNT4iEMsj/b72qRsuGYCgtm8YgErRq/
18CgRKG+8bz8Zc1pVG4kp8OLlLYoaVvCGE+33D3dFt5eI5QhMPErCYoqeJ5WwCA+iDsx8bqk/hax
YzLHm1Ez/HTYvy2S+cSpz2hlq1Jxq/ynRCybvjH8vjGygjvhLtHGgF/HwQ7+HTQej7nSygpPZNQF
f357qumT35ZS1PtPV99NL2G9oqR/KDsZMdXn9X4q7iOfx4nnBiuLNTmPR9mtaLBXzJ4CkF4f+Wqi
SKvTUI4Sa+i4laplf4QZEFvXcJdLD1mZrrLYSFmjFinzx0JW5j1CYNjoK7yc5Y52M3UZXy83vESC
ffSIfFCsDF64+IYUvzPFG768Ua+GpGQ9lWPFG0wzj32aqcZM0H/co0C4Z5KXFByWgW+4FzeVFnxo
Nq6jDgDPYS6Pja/YieRedR4kQPsSGKzqxKLwT5f1nDPABtlkKaHLYdb7dZ98V6Q6PnzwiZAovQax
VLTU4xOIFDjr02TB5zgdh9EAtnUSRl39AS376LJMDqc0My/ty7xh7tGq6ULIOhe9NXS5wQvD8My1
JI8mrXRW7QmyJ22gWEGTMac3CpjTcCe1m7EGbBEeUpqbETpWZpSjYfx6X++CD+hG4q8FNUBESnyN
v/ytD+qIWcsuNRUIycJftFdI+wL6pZyzCfkNq0/27iM+VXkbh1I0c8X4K7MHyNdlh9W6hCwPbus1
FGMvhCC2TbtEMVFO+Tthm2l4rkPIcFlRdXMQybPEF7e77hJd5bQbYctqeTXrVINmHWtaqksb/PXM
Y7F5OwBQ9xRsKoZUUJB3GipokNIVzCQtv6FLcvWT6f9XFThqhS7nnmOj1aqoToxbhNZZO6LGaSni
r0W3i8Nb6zRuCMnxluro4j6GQL2gUQOd5SItpO3oJySEZXu4O77jH7JW+beqd2RPLn8WADza47jF
hkBDauf9q36zTL2QheydsH1YYikZ0kwq9MvXpHfuLOqXeW/nRN9Oh2qf3kZOFMCuZN1LZS8VVSxF
+ZQzWU80ofswfDvXdtuymSpNSDhjBC5WAhJI4lvVxL+57GPNJX58AZvT0cw5f2IP2RkK8E8gp/ug
hu98qmb5JQK290pZ54/ivXb08gNhASWMnYogMZC8oJCsRqX6V5hRHfarqVl5OOjGeENhbo0UbGf9
+8SDNLWPJenNiOwHxJqz4O/PdYg/SsMukITg39zOX567OD6k0yl2MxuQTYRFFyJinvWne7ziArEq
kNejnOhgM3mY1RIpuX4vHahRmB/gszJ9ISRovcDE7eNrP1UDr/v8NnHJTNp6VpOqI0b4qL2ErHub
L4TZvFksIWQmEBI4zLJGhdS2U6rtYwi80L5COEbKV/C+mvqaCMIEi8L3efZQHhelHRJiJAM21Oh/
3x3cIFeHjoVq3ysP9N4FVTpQyhVwJBg9PmAUbELCE1W7ZvCvebE8tE/utZtQ4AwvEXSEjWacjOH9
hTWsYbbq/Vtq2ODVn34g/EVrxOLV7+ENX+79FiQ2Ro7yBW2s+EAtUumfhUJrAwlZo+xaYBl2HCpp
LmQNoqk1gvLSx+VeHdu4Ve2Oz5OYER2oyKGEKqRW43g4+Oflrn3pTLIy6ZPKXqFtLBfFtZhD4UW4
cjvxZVRutR2D7Tn/xUo7HPxmtVJdB2g7Oa1MvGv/xIYxZvBRhOjaQyF9fnOU6Yb+Hm2ciCnzwVyd
4b9yIGAzRoQML9n/LhSOOjXI2rH1mDJ8y/rWamMie1/Hhc5W6ORu+MmiTe4miiL6fjO+NSS2sqwq
oi4Eblz1RM82yj7G4o9nT0r+WN84LYFaNZZRuFjpHlMLMEvomWf8RNRq3A92OQtugtMR2SGBK4Cv
1OLtHy1eKFgAC7Zh32zhDMtKAuVHpaEJrsG+0P2KkJ3liJ+l3AeMEhvHn/YrIyBwgcbQMUsJSRks
jGo9A20/RT00jMcD0SrrLw3hk8OlOyjOChGm+a2fRPYY6dH5ZOb6rbaSG+9TRilAwPqOEOI9d3e4
dei/Ik60FO+gfc1S8V6qfAGxHM6ZZjky8XfJjtQYqOPpER0AXYe5MLvxuWHl4Lp0cnL7sLiZGDuU
vQCM3dNeIBHww1JVEZDJtfcpDLAy0UVUbvFx3YBu+qLeXSiPrnhVaV7cepPpKUIX7zYvqc5Tj1fj
FN6VdpfsUffWgNvK3BU69R3kqWyF3LCpamMN7WiQKWnd8YJxBOke0kzzwu7D6ttC6qAiU5TiZP0e
YC4oHuNjsfWJO/AoI85LTfU/40i3aSXKIwWXL2PvRIDtb4h9GsjrAjLWuW5BtcwV64wLyJw6NM0v
1Kz0dGu0x73S3CZlTB/vJkaFDpC3S5W2O5qu3ikktD5molOt8PTcR/v6ZaERqVrVHx1SdmQbOA5Z
7tZI2zvZV5IZR7HpG3ItQTtUW3jzUnUfqj+WivzUaKm87d86YPtl2hjSZm2yCT2zHAR+xhOcOiLx
b0pjrkDUS+Q4s4AkNwIr/WyTxjibW3kLDNt+cK4Dm7u8WF8nXRTFQXjEXGRjY/YBY1b3FHZ4c1DC
iq7EAa+cbF4BBY4dHiKvzxgOfg7ZEpL6Ra8ohAUUNIVCgd7hnwMswlbofQP60rE3NfkGugyp48D9
5ZTNJNZrCJRoKvpicjGg4jVY53Z9o5NI84+S0MbrAgnUu6M84nizilzSesWhWm0vdqXXSZp543F4
w23XjmB5gTQFIIEBMb8+d1ThnipbOe08iNYuD7M9J0u0T7O8EwgSCP7QZp+mImzwnwMITIJ2IwzM
+zN0PsxkdZYbQ+hIPJJGQ+sk2HoamyCVDhbp4dJjS+rD/NszVS9/nbTRG6c2plX0poDfKhre1r4P
uEnVcB/lTwY6xQIMUwcjMpTdKNnPJoNVpW41+ciuMqK4qdgE5w7wGHUCqLPUim/3MGoqTucs5FSZ
C+gNluzOZZ5sHuyNRa0SGhwlFReF8+/azGKXMvEpeBidK+ZifYwv77ED8CX8h+SZd7hH1E1o682o
GJaQJMg61KIO1OzBYrdu/NYn58fA6NBOXHlkKUKb6WauFaXll61mdbeGbLNqmHPNHmXgXgPI9edp
KgpmbUtl8mNOWfIgMghKCEiWWej5mQvh+iAvt+iY9cVsOijG52QNlcTPJmkTOt6008px6QND83Q8
rq1ZWb1dyEozGJxVJsrclh78AKnFj9485+3YfkKVd5a5XMUQsbSGybwn2ztB2YTRZuj/TiKdQq2Z
6athLodUYScqcumvL9IFHi2f8o6nEFBDCJg27ORCSIs9qiLG+oMTIJmQVS6n9MaHB3PKTSVfluL9
lM4tn+S/VKRgO62NCRWQFXxrb49J99SzLLr/8o7cczO9lr/JxiuKOYbzZjcI8HgfOnNtJpgvdYeO
mcrI7sZJFEvf+GhIV13M8vf38JT0B6nH05a/J4VnnlbeNh0xAxB6OMAp1YKj1QopwpxnwO5Zl53t
OTmZ8u1Ex6HLTx42ej+9fB43vfkhrRP30P2abPlXlvjKoiKOnMyCZhhbQUxOB7WUbP8nevL51rAO
tAS70mzKrkxR3C99R5jJpYg6YaTglPCf7Z8Ys6K43LX/lDvZ6BSCv8CLR6iSdXN5C57NgV59Iwl9
7DjLJSIIQyZ/i6m+Rs3BG/njBotAk3acXsQZaIaJLmeHuVuGgXAnr5kBeOf/lrO+MKOmOQZ6oRRH
+HUHGnR0ua4Xb0ciWNxgx9k+9dalbrrEBAxAW0uU6EYOTID+Y1/2UvvAKn/t9yZqibvaIjmXf7M4
MxRwx9zyILcitYcQLNc2T/6A/y/W6x4W6UPVIYMCE93vxqsIRBQpR5zJZwGG75VofC4pBbaFQeME
ec7k26VZc2OUDtSscbC+6XqYlyYG8QltzLege/KaAm6TSRn+d6in6Hj4z6ycbwHXVKXMgwmQkkWk
Zgk+6xsWEvXeYPEOAaNtwjPng7U9GigiBp8kogRcQhzs/tC82an8JPIGlj2Z93rdC1iVHPkqc5o7
vAOMzO1/np68QDNz1lkq8TkV7EVzWLrnySkQV8DruBL8oQlatNeus+VeCxqPfmFU2V30auNuk1Dy
rcoDZhuSdjSnSZUWVR+h2w6Tf1/wtCqlDT1KM0Lqw6VmmUnwKVqhk4Vyq0esXQV3A0YjYUUXX5s3
5WIHBUgfegAqE1wn59BQaShPItj3JK3S9hqSW+6P5DIl1egkviYSlNry4lmcVJZCHq5kne8sCO22
fLA/6Sidd29X3KbuQqdi19eIphrZumXcvrgQAc8WKkuw5HBbOROd3cRlQKOz+PlO4irI7Wh9k4/F
Z/tLbjlIFEoJsBJs7+hQdv/PJokOpEtkJNBilVVvq9vNWcd5fh4uPh1mjxN1X6OCKcGBqY2cmopO
cCWwvfCINJa7eYJqLB5znccyz7FT4KMi/s6KwF1PuZMWLqX8r8GvdKwKOhqG/8qqmpvap1x8S5gX
eAUezBlgzFzP1gmnIz/adJg4Gfd6nDoiLLHehjoJKlE7DbRkiuosCGrtW+0z/Pi9Coa/KxOH+ToO
hDGgaKqeY797TCMnVmK6tZ04G+hpIhETs0IIc1rsVh+f6qeoJhmCimhrRaUBXlrzT4bQHE+2MS70
PB7rwO5pgyWEqKTpS8yL1saaqKn5qjfSLtWR26v+xT9uU/rbPZgGOE2eOqRtPv961QyuN2wW0Ydj
Vo+DpoGOu8dHTfuHcfhPt8b8EPvQZIUGqg107xHCci8BGU4dLu0vxyrWyJiOXzbNicamadp6cHZ6
aAJpSxCm6CQw+//loZvIExdLsiKwPaDr8Mso79/vQkP2e0w1Tgf4Yoq9kTIuuOpJjHO10VIUUUiv
zJr2txRtYZCidpDoccAfk0KUKjJagAyRiJWhE7ZDy/EwMCO611VU0c7RG03fIzj4IwGiUqajnyma
Y5rH9pNaQUVZehCk50X24KUxaXK6B8tk/aofblrc+aZek91MVmp2xwlvkbiaJuTp3JpZO9Mlz5Gc
dT6NJGu+rJPxmOq2Eu/kH6wf3UoCpudpmYomRshvkTQDRU7+cnKmd9gTL+MeAwhBOGwQ8rkFgnWZ
Qfwm5c9t79/4zkXhOQIA5KVT+ckPYJzH7+tMmmXzfDeLJ9JdfG3soLIa0vEB1qV717A6K1A4dHU5
i0kJmPUqeosFPno84X+4XZuQaMSbpM/m35ZnWOADbndLEz3vesl4bXiZairTiAfzwVx/oxGahyBY
ztrfxGdS2Sri7RsJgZyd+WphJslBAb9YBycJaaK6MmGv3xsgh1/7+uo3yIn8olgIM3Vu/BCIWgxU
blf00eWARRwccs1SIE2Nr4i9dQ7EZLSPzEaRH5JPYDH7imSDex387OviggifwTYvFewvLhEAzZPG
zcz+KSSrQ9SM8zAq5fKShacEOS6OAbkQUPV7tcuaEdPBEII/hOOvHHf/ww2XMpLADXKa/eolxZrh
i7BUWZagFH5fCIAuRABruo6j8L2o8O0iWmwCcqS6ghBX9udmB/W7kNlaymnIbunYltHWP2tAYNDv
KD9MhUFv/f2zBdHcIa6vAHqmQY6pcN8iFejGfgQ/O//Rg+235n9KSgqd32rXjQDBeJisfIxbzL9k
0mViU+PNl7ZMxjIYW6IR3Laqycw7NZdbQ/42NeualLnlEPKbFfH88NHueyUv/+jDSi/r+VBZx0Ku
/Tvr0p8ikB64A1dkIYFxawXNrGfik7P0S4PRkiDSKO+Vevd2Wv0dIi3X02O0nmmcNkHcOfDIyIUz
dkGQzAhSTp+fm3+X2EsfsHjtLmRZjD0gH3wrB4b4JO6HjShUQmhqN1d/uIyfK+gtbJShK0Lv5X4Z
e1az0UT8D0LUsivanJMu0paUU09jQAENqbdU4MhEC9YTuG/cOl2EcWqyAcCm6Sjk9pfH7F0m4ku7
Z46iS9uhGGjTUubsU1ywgwyqB2hXiDwoPj0ttqGGYO3Dq5e3cJRLhN4EVAtCF+IWzPiJw20s+AjG
MK++vIWMAJ4dBSVC8NcuU+uobCNtMNbIemTcYGSHqkceZPfzDjGKrhsn/B50ezrkgjReaxKR+wZs
eczwaHSRqQ/s0jmNVW+1khww+oAv/8XfniaIuEaM6WhENIL1oFLXSJzTR+2gMK0A4+os8Te6bZcJ
Q83msDJS+bR0CQU00Envxz4tZB/r/XYVzucx12aIRA8DFIMMN4voMuD43mTwVapZy5RP8vJ0/dr+
Dwf6h0MG8FptKKLTbDSuez+HVmlKs4la3yNX8Br0B77vbUdVZoAMQUYuo7auSyjSNLwC8bhD1iQD
mexkZzKu8u02KVVq6xX3CG8pj5vI66pMA9N+sw8V/Cd8e/gkVp/UVAbrAQ+aFXwa1M6lmQ/3Idg6
K8XMj/H2N3coQRmFK+7BD+5cLTFK7sd/0KFRs5D/HCV1RKyD8D+G2eqZw1O3J7eXoOHDw2v4a6rk
5HBpUL3vAuMgkepvtqWgzSrfM1IgI5QWsN51fXiLjgaczfepEnKayg8v1Vgzexh5iEuytJUskJ4i
EtRdjoKz5pkbtEGZSc1ApmNul/lSoqXdqR03+cCOkksiyhUUt1qbv+DBhXuuZfjpvwMRbT4+x9oZ
4dHtgvBYyXN6zCLEpzWRKQXnUKnDK75S7t2FOfjwJfSRD75Gx0WCtP8F+W9aMhsgIcbz/E6TZ7Bq
Q+s0E0556DYceD4KgrxvIXX7XDwNHjsk9B26S84oMetAFGMvLAQFkMfYG+G/uFFSLLRGC5itP6/W
YW4s4WX801C8Z9RukY+J0PXc1M8jLyKO+PHpktyU+SG7xOpuGtmAK8CjPSJxbELKzl0S1VXMxYYt
y6s1AsGuEXXEBHceDli2rwdi4bT9hABf79/zkIiR7um1V28kbVhTtnAkTkpWmqTWX8NnaX9iRPHc
xSP0V7TM78JaL+U9tFDk9UCByHVi20bXRtzWupc57U0scRuuwOOAQ82Cne3s/XI1XcRw7wHJ/DZ9
WArogH3JHKSNaG2hCrNgjZHMERVshJAHtn3r8nfZDGJgpzTpnrVipxc4dtjzhIpn8djomx7+iNZn
Acrdtw1OsyAvl4DyA0gFB3SQb2VgnjuQ+M2vYnLJI/2CFZiXJoCmvnpGO/B8twwNCqY3HZcA2ynP
HCCwK5CtZpMaKI4uiKCef/+RAqtGV7FnCH+MjWEBvElKPE0wybXxZFEkvGkn+3fAlw84fIrUkzDZ
KJQSj7gMBtH7L05LBlwRImrKmc1Aq1R+yN7M8+m2KToXVCnJ7Eg0guRqwICwDz4wylNOcP9m3Fd0
aKJf/DXh+U/fD1hL10780PmE4dMOg77za34jhaHXOGREtmHZgzqlS4k98S9WkkykCcwVEc2oYKkO
U66TulknjsmDKxzJWEOME55MsqXBj7OHQHcBAVBnCFVVZjKBEI29DL1B36+XC143yuAi5hNg0qov
A3T5xLGcEjvQKBYAB9ohDqTa4wcgOofcSgtgH8hIvkMyCQkihxUfaJKYN4ezpZ5S1IDovLlIgYVG
3wotkJZlURRIRImbNqFTCk8Jt1BL9IsbyYqdWCVoQIWpuD1UveZI5xXhhn353mLiWAjy5VlhkK7e
K2joy5d7OcUeRWMVTbzLY9wRTcGNytCL80zwUOA6VR91+ATJsoRjTxMjkB5jGY7ZHsMW3QcrQTn+
VPwn/c5vnp6SqKytUNWF7taYGDHYAomauFc5k744lsKo9DZ7zpzOsHm5hf39Dh/UsReXAVE9F4kc
7OSLCVQwRaH8gkcPtw8N4dn70ll1BZOv8rF83o9zxYUgaKp2DHU5Ld51AX7I34ZWF9HKn+ZkzdJJ
HohqFoyl6MItfbTUgbHSj8WKlSN4QvU7zIu55QLRXqr71CMZYCBvJU6G2HKS2raTtpmzcbcXnc4H
laQ1XIeXWm3OUqgDK+Zrm7q60t+aizDorFZ72UWJCemmu2048aUYyuQLpgM3i6V/uE0334RdF+cm
pi7XfpOpfYBoP/oHWdw57opnD2zfpLkhl/3ajJUl0sWx+rcre2bHxeuQ1LPZRESuRDTCj9AIxL1A
7mw2nGBPy9zX8DuqLNg/ntMJvXgXDkmGq1LQhp/ju5oApBHNjXwZSkiVwPh/jS/XRmhH7V7Sk3WN
hlWBOoqua7jb5cvNb0uf0HZn4xFh86AhKA67AkFCuR1wfqADCx0dLRlVOWxr42tWtZByMcxJOKmj
K3bps8tki5K/ET5bkc9DojV1s3ASXSDW/0hymb12BOwA4UuwcvGbBueaHGXRR47hq+ywMPnyGpRu
DJAVAYcPwqpDLIKo2MgyrlAaW7qJpri0ON6Jn7nJfEzZzzKlqXtouJv//iQV+Kl9XBB8T4X0Kz0w
8G2YmBiynJxP7ML21N94poK/QNEXvKXBsBfNxhr2LFKUDt+3y3ySc/ePp2GUQQSoykyBBWu0z+y9
SK6gxgID/KBov/Jvr4OlTVph3QPiOeiEKwi+Oexeo8UUcDrfqr8RHGRopP084IJ1cs/w1refweOQ
JNRExL4kaNMWSOBiBk+4gG1q+PhMFDbxJWfjw6qUgUmkYY2wiIljnhISzjhE9bPhnSyJpXK0pyNc
MycnHAxach8hNTFF5dffOf0UCRaH3W+xescCq7YbjD0r74JEHwnp/St0R/zBFvb1JNTfaB1h93Aw
ciWKcsPI8gxCo0y5A3mfgs97y4/cIVg8iylNGghQmkBFHnUr5aJNB4Led4jQmWc9tAPeupSJt5rm
9M3IRDrSQf5JdUpjlrg7HgjQZ+VKEloiN/PW9W67YONtTLPP8Q9Oij3Cq9Q2y4cO8wDLGpB9y1ay
TJAAJTy3MFrWSttnBGfXuEDYsB0qODTjAXPGYQW1BpBvgLVY9bsub8jN1+VbIz+M8PgwEKeZJMJ/
pI8RppuZkmFDySOULSwpCVrx+Eiaa+VtBwq7WBnmc4ZiV+izozErH+irCukzcSV9IeN1Xw8vtVGU
7lww5jLn2yaCgDoXReNvZy5V8IPmo/uPYFfHSwZ5pfp+6VgJvbBoQG+XN3DYCs+KjTWSzc7yn3Qv
KWALHjvaGVVqQxj8fKB1bwsGflKQsq2WOSDA8rh7YqZNgNNHiqvGaOQbANtDEtsXL68DpfksPMGH
HEQE4WkfnvkikJjjeyZDsi9os+bSPiV64J44C5NwpmA9hSS3tRU0xvcQP/xcslfPmeNMtWIoPHuQ
RDb7FJRgZnWkdQRRv0g2SyFCfiYUcQK1uikeBU+OfkNEdtU6wMwGrhBVZkhIsKKHRpFXYEso7nFl
3qQpPGaGSvs1IgILAyF2fwTaD9IcwlFb6umfB9Gy9WW/GcyLrfuCOPP9HctN0RsTTxYaaXeKQ8A9
VFcl1fihkRTjZAEfv6nQuxAV2VbhecVFkBgAl30oy3w5MFbHRHOX2d1pGCTzsaOWcQf+8YgWVKSl
UHbMwIIINGmWtiIKKLezfrRw01K8BKh/oaVpxfAT21uWWFrPwrKkVZjl0ssaOD6ytkEHWkmkJLCd
kuwiLXfk/nGLfV8T4iQGTQodlJ6pzaA8eICUGp2Q1VbdEVWk7RtXtTRB6ZY79bvxa1qi3DCA+CTF
L11hrFLkqovOtBhzrUR9MWzhNx0v9YSLoorhWcaOhqis88CEKrNrHDVsaxMZyF6QtNy6G7GC/Fb/
d3DDPbF6dL8sPdtde1Q5WfXqhHiUdfqmC/D/9Dg2LrGCJT4yByzfufhgKjqUhuokvWa+bmIjHhA0
WxK6U680beGktxlF1tZ7j+gdZfecK9nf7cp9U+Js2/PERpB/BQyTHzDCHRJP864xtg5Hm2zeL18D
XRM6dzPXpayxCqgDLTiWG4hhDzrLM3Cwev07TuVZD/t8dZpCBIUJ7hMLah+PbC4ccnRnp+2+GKj+
fJSwx7QvYft90X7Vb2xOWKO6u+rKNoQGtMfMUfy7KD52mYjFBiP5aUeJRrl/x5BdinkjhOtl7deQ
HZsWKfiVUu0fD/HnADESQZjIUr+keiWTQ8Fx/TZmr3qZB60AJnsgcZfJmyu6SB6GCOynkJurgIbS
Kq9zmCwXlxD2+i8cuWj4vuFYe/dkeDvFpwA3APjEcfMBld6FlFeeW41YQ5fPWsqwqG6lzbfPoaLS
WejMaNLFBjJ1Vrd8J+pDzrQ0lB5TQQxqsy2dONd6+IL7yTfPuRewAPRr5/XEwDe1q6HOOhPwTGLg
lfaII/auAEtanfpqPO2vBJiarbvzLi//ZLcxNVyi1LFLIRwH8ba5UF6eKUhdQ68qww9LsN+6U5mH
9oJfwbDvgWRb3I76fHpRFellg9P/meGfGrsW77TXtFXw+Iq5/XRKhAzRvmZKLEMlumluU8Y1fd5i
4uvMxqqx5zKTkrc/YC52MPlpDx+dqIWnbWIhWDudAXVP4uiNYKCprhXA3smP7MO4U9+HKM2drRo7
zHdRAPZTBZDGAFqGklzH21/gLcgs55IZE4a4EjzrVwo8y4jso32Tfl+qtDEWBN8fL1fEIx3OEyw3
0e5u3qImBP0VmZ7EDGkAVBDS+xY4DA1vx3DsCL7rBUEPcP33fz8FFkGM9l/b5H8+1PjfvGW7bBN7
+wODnyQzL9U9wAiJx8ISZIwsqPvKeRDKdH0TgLfR01bBUhbHI9k5vdgpTm5lDld+BsfD4Sxjiupz
B3G4OPkGJ7QD2H8F3EiXHWfA2KOE72MXHAcSMS8DgkC4LRQoNu8bmfzBcFAXu58Dbj8suzmvOjH7
QUVSpzwXpsjy2rdRwnbx9quhaHvVRNyMhiWJdgCQoNwW2CIvJaJIOEal/0+yINt5I5adO4dnFaSy
6/G5ZhoJEwlPZQLY930urBIRJzBQndDbJv1hYFOzvhw++xrianAQoHTHgBafIg+P39A/YOjIBbtL
+Z7pynDThycdYy6kNFSYRBpc37mqsAeVKNSdqwOQ0RbTcxeoJExjFbA39UMeTtWBJLZtJqDv2XFz
LA2vwPTIfEND5FgnCerrInehI4gzQ886xKiFhjCc3S+fuAUGqdgx48H6DOOgt6q2tdG0fFoqylV2
8HlPPDrxxoPQWL+BiCjAHx+FzeTbjB3e7BVg8SOSL6syGJVD0jlkzqhFocyA2LVq+XfA56DRn+2w
e7/INjqXQnmwDL9pnMF4F9ThlkDXNJwrf8036zRV9uT7HJbVlW7zhPXUv26s/FzeQILFsyhI+TfI
xK3Gq4uCTnPfI9G6ck0S2ZVk6CE4T4hyb/E6u6DCHucCZ5ARY8h+4kz/2cky7+3H+WYcM7AITfQr
Pj1gT1qIOLeHPc3UsSPm2vFh9tUPIia35DmiUqnzuO0xeCMWTo7oo04XVGsoOx9bgrmF3DKVAnVY
VTu2SBz8PekeLUJl2FwVXEocs/pAe9G6FSyHzDucuukH+OYv972q+fJVaU3YJTVKF3SWEynRadAF
08lmEwcXOvVMwzpJB+jwkfINZkdagztztoZlxKCgB94K653KO1uDB3tRBvSid9IcCBHjoOopu/8/
MRvW71+b78zsWTE/0GBKlrDL5CogW4YyT97oSZxy3Loa0xu29TNJ9eRudIIB14DRsoKVzmCV/jOK
Bl3nhonT6StLwKLWItxjktI6ynn5BfT66gvxYyg9WurXXM3v61LaLwqmuZyyNKQvG/ykIevEOk+t
FI5Mf369rRdmDU/iGOFtofy6jczjFh1IskjFhtWvhTfaHPQbXjJqRpSwlNMMbUo7fY/XX1jnwlzt
21KsgjRjmR1rEhWv+uxtIOQrVOAdFTFpsNDfZSkhQyhO/GT38LB7ux812TLlLgSEgT0uLjT1ZiiM
FJ5SCpFWKUExLTMK4IrmbOfBR9ufi9W0reAZXDzijkonB/jRuBq2bSk4cuyHlpKVh2VOgarmP+F2
vTFTpBtVJlaiU3zanlRTvQVWYt8vmEM3zgK2eplAPzvSCVOgoM90jtd5C/PJYJgDAfjQY/AZQnfE
4QOSSER9YTrMEqkr2rZac+lz1WCe8WHQX4wTxzfRc8tcApkla+bkgUkPdVtpQQhEVCCq9J8x+7j2
pXTG4tEMZpyy4zvwYLS/9UW/cSg0jd1pmFzYvmaUa5CJ1gfNqVMFAHdYs2I9tUgU9AE0LxuXtYMO
eBtXYoLDe0q2Vkpc16Rv1vndzxf9pEgNPIq8Ja0UlJT2CK/A69AUpUmqGqxX71xnqhWGbGX2sn/S
/gApjJ87aHzpqe5H6FEhHlLskeWj6CJlFYFoNP1yRzw4wtzsau2CmjZxpjTKDYEfqcH0v8NqSStg
aqi9yoKRUXTDfvC8CfIMllz/ruNgHX8o4U69NFPHRnTda+a3MkXUaN7SIgVWkYz1Zvm7cSmzXIqB
R8Rr7V5TE/1fka9PZABtmvXqTsANK1iiCnDUS5FEHNWZhiSu54MmdwJ6+9yulB5+IqwtKfsNANom
+RRtym5VQMDRCJIJRcssHb/UIQ9Y0VG7yITdYkTrfEIlMLlvXwXpQ6u7CtGSbtLFJkc6qxiCKv/M
Cr+AuotiX1T8ueQ6wXDc1bjt0m27lSXfuukBDl+DaarzFiVnhFAI+xY770bj7Cdtib92RYnkWW16
rb3DsP+EPdWdtGHaHxg0ahpbuvUa+uU2FfKuJYGgVFM4p0eZAmlt+LRmp+DfmaBriyIqLWkOHry6
Lcx0O1vpxmQpRLhyRHdEl6SGqKZGucx7J3z6bBr8ew1HMWzXCaKFPsJ3a3iUo7hQzMN0VkUEKOLF
GImjPRkraYzTd3FhIVrnLu3Fy5WVwJj/fA9VoENYSGdh7t4bARSpFqHReBBfDcL/fFZThazegnBN
DVxSzk5lW1swnlbpkx/JDWSmLeR4/h5wleNd8VElC1D5xWTY9pyT8N4JmfdazRT3oDMrHRE6eltg
b60dVW+8ZckXffoEoesq2mRmZcTOkmLvlZEOLKXWNm4avhfPHKkIAVyvNhgEG/bk+w2+i94LFqrD
0tyGcJMR3nLHCi5vQ6unupECDsajLqs7zSJCK3INOgFruimSzTqHgnb/1xrKek3MSO5NujypI7X/
f38Ps755RT+ju6o4haTnqK3Niv4dCuctbq2YSviI9bAaXBbjRKAI2lpBU+wjefRBxyEvCRZ4KTGP
lzT8CVwsWwk1i2o/uCHoBTwGdEfz0ouLjih3E/aLZ57wn3RJujJjuduoZm/E4gAN5IjR/vFqHDmA
h44sRUWDQXLCa65Wye7BTvo4fWrPnP4ZD2YkANq26R3RvBhSS6nUq5SKzcaRuP/nU/jNURzNNQzW
yfoJUDZBuX4jfUO3YCWG5my0jte5H13CjG4vs1ozxQsMTcMhrIqVUhqQR85oZFKVVgyu7r6WrPG6
qotmlgQQmoOuxFHLygVMZkFKPrTwyWClatNUtxi3u/98nWys2EdgsRacdzjwAlKb/eI1S6lVoFEP
bP12yVb0E4XuPwY2VmMyHizlcmxbLYc9qOkl9XxOXoZl03lL5pRU76NKdsLnsuD49tLKMg8ygKPp
o8LU49PxJYYkv7vomJBHTanfgUFGXJ1y1qJsh5tIwuXeS3nhXbsPEtdMceHUERUo9eHFUsYoYXpB
AZFCSKHpYHTikH5TlxOLBFU8zo/7NgXoRvKH5Qqa2/uiphXc/dSdtZ69/6uiwdOFMf1BttETP5Ji
6UomYXOy5VS9H7vbnrUy8FQXJ58dMtIGGmMj34td2YLpXbEIyN51jkzd2ZD1sIZllC6ldUq+b73C
6fZ2fax9FwBhGwwVufQWMfy0T3OGnlFbbbWkZEgeoWwy9pdSQnarxS+DyhsFOih8y7RwjMLhiJtf
/jEBVChSaTzXKhC+Swn3N8JXw3LcDO5gXx2XRQR3t9ktNL8JAgfcFGEATSpNrzJlAz81QhgaOgvQ
Y3wQp1wCS1NxCOPHT2CIiJ475jdZlmdXce6iGM1HEg4oxZV4vlDcWKSYyW2p5vWPatz75bdQfuiI
7NpUfHfm5QA2ejdxinC02RI39tz03SSQfMaRp9ztiI/NJDMDnMm0mryxFbRefxq/QEddDeA34hVI
E2xXiQ/JyV+l9T5rEu0IoPfaeXgqFw2kfci4l8yCbJV6e5JItjrgIa0DjBcUbI6frRsdfA7517T7
bnCOS5IRgr1zxOneE9NeYZmtvwKjjcNverMXH6h7li6vAzgtreoqYaN76YYFU7UIVlCi0HjTM6cv
jtfzkno4vr5B4CRpNqtZpKKuq/0xBOvTqV6APAp8Zk+/GyvO/7DSgKxILOB/dKpIMDtjwbIpff33
mSg0/BRCqE+fQPm7FvnF6JHleIThjRuzJVXF4LzeAQi/IMsLN72b2k7zWoX2K8l7TXTxP/Lq4qov
cpBOJuk0xfhhcfueL/Du+C6m3Q+Gxb42cbmkm+cKE3w9xwE0jkWIisVFCMrNiGWEkBbPVOhA6OMU
sGrZacJW4ICjyfa6YjWMkYhXEnXE9w8oE+AY3QYtXWcWU4hLhbNz3mvFBOJu2skXDaYsLBecVV7G
Xu2wuAGIazGAG/UqL3ECuaiZpxg6wCiK/J+WY0ah8dIE4G2w/LHwWUb2pJEdkGpS1aQrDsIc2A7e
5972YoTDn3cRSOL2qivuCrZjCbtgRY+eevHP8zq6FT3it9iKhOzbLuOG3JjbNDdf48YeRsQLYk+H
UyOyXNjI0AiZOwVCSx3QogYYOO/FSvc6L7wT8ShxR6PZF+4pIxfgO6UNE6dcyIolR2Ft0BiNNuds
GP7jIkQrw3M3OeSGBtud0OtQtm1EK9e5Np3ND9XNNqeZLtd3bSGp7O8pVTK6uoMlVFofKpIUsRzp
spi0/vsyAAptttsiHg5PuuPnESVCcGUtgSWFjzvdaVSSEDTq/rblf/q3Cwbu/abdI/NC3YyzeiXF
3aOV6NCPjQlrPLK6lKhJZ1oxxS7KxIzIb3MM9sX0aS/G9aditbY0aD0eG8VQb+xhyOzbBwFSxG5M
KVfYAwD308WeCMI4U+Nv/G+4cP+uO3uhb7lpqdq9fVyUW7YGjkzKDzcglvrCU0idE2fH/9SglIXY
899tlR5jcS1DyncvbCF/R9zcYRZjbClqDti5nWX2U0Db0dpHfYdhITTZmOFg1avg96bnLyNEOckP
fLDGIG2mdGdzyd3q8IsC/vLz8J8qjhH03PjySOhWTk9bMRoM3UFq/k/kRfBJox9yPz0l6lMYoF9q
S9VWUFC90GO7dFPnFkTrgas1/NEOSpJGvHvr4SqtUfdJARaRXh1VJwSGMQyIdPyMKq8zUi90tt56
m57D0diXfgAyYZa+b83vwee2cWbSAeoEgnglK5gttRiqujfFLDr9SPyIn8DSGMuB47wkfxx7FwxU
s7yWqG1u2NZLx08o7IUUejibZoV7LiRoK4LytSCfHag2aelntm6K1o77U5IiLSRdQBbcVW6rOEMF
lhmcw024stO4Z0IPi9s6SXrntivvMqL91ZCw/GF9Hx0m4IAI/rFU04+Gn350ZA86c++baUBjuHrk
5lY9a/X+saBnD/+o4ccO3U3YKbJbeEZX9sxr/+YIJoKRYl7Ynhb1i/8t0DuJ77K9hhWIN9/Pxqe6
jA85cDu0ZH1HZOtybt9ygN+96lH3p3X37JTJQSNrwlkBUTKWHhsSvMC6L9qjgYiaWpDBE06uruU+
nni1gEs2oQfbAhCqX7t3OoZM/m+vdbenZNLa155Pg5A20PQsQcPpCRoQGMDOflDjNFxAkn5aGULQ
4tVWC7I+DUe0ehjne/5m2ZsG0OKoMmVB27QQJgd3ESZnLGKXw6T6rwctjXICSbnfWlmWVUlBLuEI
HpECMW8bwzXsDQJ1GsFBkSJvWhkDT7QxuKXaPM82gfflpNg8YNrqOcZh4vpd2zUIFNhfNX8REmq7
2QXcQobh/0EbjuXN26atZFGa90pQE4R05w67YU4QRl16guzTqplkSm2edwlUjNovsVF3bhlK/2k9
5CKtszK8dVrIH5Yn3lRgUB478jT3uKjwFlDUAWCXddPVkFUTzmg5i1PCctBsGvmiZIxLiBep0MjT
g4AGqYnR7qogCNTLnB5Qavh3Z7dz+i/AVUftF2j895f+AExEk8qUP3rfztbSnn1el9BMfA7ccSc1
hqd+2WLMBEkvVzMCgA1H1drdeNYtC8Lq0uZifsxtlk9Q2fY6ZzGQclCXXianrSCDyBhrCeGZ5qCs
GxoJ465gnugDaOwpJCvJlPnP92xkBmeacxncUWVisycLt6aFDi0+9IFAj9LYgRkFLOZ+O1AAeU2K
3jYat9+ecs8ok5YACp18IcpUVwAIkhg1FS2z+ZJlb8ObxMQ3Bprx7cxCcPNG6qMMc+aRr5KIQx2T
arwc2mnDXtje5ZvxEsK2+eFPbbTxclwVfPL4855McduRET+jrENMyv6A0xLAgna2kFX617NE2eEy
LQvnNEVvKUy4moI48COSE5bwDHdTH9GYiOJOUbUCIjD9V+AOogQXYeEgky3GGvMdvtpLDx5r/0ub
0nKMRrE+af0dmQx64aRS0L0jz0qBPz1OE994yRlRIbavQ21iqFpHPHomv84xFh8yx1JcPa7/GB7E
gzfsQeQr63rO8JdR6xVz5XfrDVeWqEczHIvaakN1e3ACWBlPA94zMEd1i6/6fHYpQtbBdbmAn8cl
pm+VVCg6UVZgMzCVznOl/rGTaNrD/e6CZBswQ2E9XqqcxZ1686bZu4SzU3odoPPo8jSMoabtGYak
5tEDknCDtY9lpckjjgFS4K/8HkyP/oLMk2fBuAnxEZZhOtR7N2NBq6CuEtuexQAp+cozWuM3U2ck
JQf4niyxjlZZE24KXAsJ6536IRl+vuOIogIaCbDdjANWQWsRBOVSrrUEXONg+izjNNxfIvcpt+RZ
9rMqd769ux0cbAQN8SRcRBpYmq2dg74+XESfLLcAFIbPC4izecMm3sPxvBUmVWkytp8JheZpV/kS
illof85zdYqQlIFPab27u0iev0pr447Lb9Kcx5DxB3STQh7qERDU6WEzhc5LnlSR29Io2H3shXp/
fCp5md7nqHNunJB/2o5mxKFCBsmYgNcJgN2gpAyaAaciLuOHZPE3+w9nnEK32cCfVAH7H6myIcdm
kL1yb8eKNRri5nw32IsqsoAE0ftGZMZmrUBhl3wXgMwc4M+O+yDNwu3uo13qkSYmb0G1eMk7QQ3r
I3AYFEXn7pF+kadExsn9Im+vLKRr9uqpHsf3H5a+mNVlU23v/O7v63j7qPdam6dLnpViXl+gF2+V
880EtgGp4yeVxcTAIMYAT1f9VzkfO63gX56Y9JlbMX7IDiYqfcnjdMljVV94EQ1tjQ3w1v6tySaM
s7sLn+Ye6FJAuJLUzN3ztL8IQwkuTvWlp6K4Zy8fA8a50CG+dvNsHZQ6GD1xnurKgz1MSxME9cUa
LcMsjGfPUq6YIiDE7T3KI87FG7Pk9B/3hmaEmiCjJgAAafCSxvpJMwxvkhlbVm1Z5fLjBLaI2WqV
+yEPHZUQNcMmr8RVxThY9ljGpxTks6ja0QYDSz6yfquPtchbkks/cOvzo4QFsLDyik6awMPad6xZ
S6S13sdtN0Bs81uV/bQw9sekiC8oVAw86QVnagTjcZnE0GGdajFV0WJiiWU9+QwY0Wgux3T63bhz
3vJiB4iHX8djpz3k8KS8KudKJg8KvSZeHp4RF5Vqs1mA9GW4kCX9xZdJ59nIu2AB0BQDqq8aMx/1
1QUbsLa1NhcxlZKQMMyI9Qz3BLBoWe+QI/hctgtZ52gENoIAGPQyjwi7bkruA3CUSpp695UoNfe5
jEzuJit2julshz8uVbF+8dN8InSrAuVK/Mwib/PTS6ldV5i/Kx+adxa7JDz7IyUTuqzRAsC3ZI0J
4y8DGS4jkX6+hr18TGHOv0L17Mp4zK/vTHDyr6wkgmGsmwBIbyEWU+YVIs7NTqYOtg6WwIw7HKSB
AFlAMS8d2sCY3hHm4P3CN48dFc3hG2G3iqd0JIoe7HOCCqvKqP/VMAVNLvlWNb5urcCWGc4VOxmY
DM3/ajh9oQeVUTh8P5Oa881wQezxzbAQfj4bztgJdKU3FdE9YbhQCbQrZ/LyoJS7WkrIa0I1TKon
e5ARYbAz4QapxenuBSBYqgk/qpWMX/iKYM5dv1xMce8iINmtrTMyfj+oyUTiBLMI5RZNny4IsFWC
xqdGQ2fcJvc/0LbNf/zx2TSfeN2G1Hkib7wn1cz7ti0iRphDxNJe+zMNg82NDUBqOZWMP/OWH9A3
juXI+UHv9oDyXyHzyp1VKtWVI+SoMyJeXDlkfv6R7ytDkk/BePdUFYMDdAcU84ARHw3nKyjIP4Wh
jN/gq1e8eBJJ/nnwakxLV9v5CcTnjcVVWjCk/cXsJBMqZDLrTMBBwf+ypAFFXRLAesQItnMimAp3
vN0VdAcf5rwnWxckzapNQJAqUspkcRuO+W6Yew7B+VvtBGclkxsuD625IB27PivLY6Ezou6/BhO1
tsgQUk1I5i0+WCudUMN1zMzNCi4eJ/v8xRgw2QSLx0f6K/P5KPEbWhT7apw7hx1Ya5KG7ItYKau4
P0yYKTcBsnTwohyi60QUhYuI5UbSzA2le5nMKb5QW/v0HoKPVf7AjHfsaRuilbcivIDa3xZX0Vsb
T2EGjwQXesShO89Vscv6CgkTIzKnWOCZuhPxC9RHb7rTLK1Sz22mpT+yvbehCwc4ZkOXACYtvCMU
s7avbLfqIiW0i3zf8z6XmJnd93QOVKctwUrUpOCkEx33At8Zx5N8QpQKP3XbjQEfkQ7TZWKBd4LS
+fjV5erIIsdQaCIpzBhA3fbBDHXe5dX2Oyegw5dDRzcc0Yo0z4SUmC/Knrmq3sYPyptt5uR6z8a5
uV+EAZsp838d47sZ5mJXbYAuOAxszNLygLY5VhKPXw0fIzbvZiEetBeaq54CaA4Rlsu8efqvPPyT
9as+XWWLuis3QC6KA6rH0YIy+jb0xWRC8u/SzyuIqs8q4fUI67nILlMGZ4a5Hti/vplRJT1vItG2
cYakKWqxwbEiP42dAz+Cj1M5PiMp8BqwdjjvMBzyLAylA8FmYekYfl2wDo/cNBbfAOvfv/34mU0S
LVJ1+b9lGj8iCV7vzXhnqJVQqyi2SEuIsSANfV/YqWfw+AsLI4Mjztf2MPOAQslRpBvrda4HIkWJ
JSJeAB251a/RzmKOZc6xgqnz8vw8MD5FiqsTW+FKB0t5aGLxChK1+8Hy33y7j0ymlZhCA5Mivbt6
m7n0satwFlKteFpzCkLAA4JiVLgnHeURzlczZKO0+3lmpoNJi4S6noWmOQhwg88flOe6dq0Gn1vf
P4Y+JqI6DBf4t0sq8iApXmsXM2PXtOTMwaGcfsXFwm5Ecexb/XVvEOc8zdJMMJELCXEheSF80jUO
23/dAJN9FTnsDuwx9iQPZThXY53M6aG/mx88ohbQ/y8ch5YPyN6wuE2Ak7iHDjBIoW3YimQs+I75
DwMcFvaDt1wpptVh8fAfOezgpKZXYOhYvVhToARNiJ5EIBsOqzcWGaYYJikxG4IbHUGXw0oXKGBR
ZJFjOVeE8b1Ux6xR1h31h8zzCBwrJw21XK23lQ4P7P99FU0kmvZQ7PZwgZHXDwj42awtwDvoaQJd
MHKn8fT7XBqH0btdQUsAzN9DCVXAB3UcTJsN70neVkp16Iiufxo8sw7oyDdHGYt6FfbvgehOk3aE
0/LYjjvZFOxr0OFbEAg4S7SC/TgPTeSZ92D3BxgSCelrpneaVaAuFu3n30CJaRWz8/qDgeE8MbiE
ZvBcVobvwYLhrBilqv+NRbBWBgyawFo6sOrB1khfGIaf8hrYY3rQ0d8gvvPLK65HdJ6loHIY5XCl
7ncVtZ0UOpEu8jR7Yi/SOR6JbMJ2O1q3Q5XQaGz9xJ4a7xUx20WiwfzZIzn8q5r+01yVAjnUKCwM
PnHDLNokQHvWclSxYpMV7SKRImjmrNj/Z1QsQuW5aba0yrjY3Ozf+5eh1qf4gYM8Pn0gk25XRdzO
yB20jf+a+RM6VCdRRh6UK/99QEdYsbHn+EpcYCPQ+0UmsEH8z/mfCfk+H9zK9d6uXRFm8YGk6Sgg
XEM4SRhpNChwLjuFbKoge6YYPmh7GmXdSlrNa16yTMo/FLYuxlJncW+mk8tb5iTrZtUV5vQVuhHP
oZll4z3V1QyfM0hCFVyI/ovQm3BiRTK42b6aaHF8yKmVfoVGOShfgwnarye+fnhqrDp0CfPO/vOA
GORnDQSP+42IE+hhnvksQx/jHmMMpfpPatxbTNSDf7+bArJCIlzXrp5wxlF3AbQ09kGM3LeCEvIK
oBUUzIlDb+T/A+fBvvQBJJkeiHy/TUSIvRH+cdbQzCYZ942fdibpqdOSLf9yPR3W5lq2H/1VsJzK
h3McK7xG3ruGrX6mgyXzTho9iL2ttc5l74FxX8anTLZBQsHScAJYqfUem2VRFf6qiyOgPCZghUxd
aqB4Cif3lKoViE8pSDAZm2HXSazqRxpSE57IcomO/JzIkisBnVu5Mo8Gepj6IzKO5mQeUgk7kaRR
tk4bP+agBMpYz28LFGd1b2MCXoDrWV2ha9O54xUMU4K5HAFGGxZtOzIrzfzdHrTSuCje0Kxp6O2z
nNdRsAYdUMCSJx4A4DbenVvryWtI+Kg4BH17QrmkFBgfSBGlydOkC3FObxzZjaWURxWGdzl2kOYp
Az4fluiZnEqmZYLWwdjeiwgTN9ERJoL+Y8rQn1ZEgdEI8JLOSXb6HpOidf0ypNDWbWN/rFinGaCq
J7Mzm2XW8IriyTfYSaWMHRVHlXmwmz4aNn8NEXvPJud79RjW1lyV/ABr1GMvu97bZLuCO/j+3snV
Q5ASsGasEeD9o/2YXYO+vx/ENmYhY4KKuJQ2hmR6WGMx8h68wkXrCJTpOgi6KsmCG8AgWpMrGHj5
9P37XSxB4HfJvXKij3Gt4jLbwM7BZLZw2zHmzFTbS2eHnqtVxpvyL10ITBSeaCy06ylXoDW654jK
mlqF8U+IUkcFfxih1hVToBr/Nbf2I50movuknm0ScDK62oaZlbOZ3FGnmyZup5hpNFGWyuolFBDq
cw9kSGFuCKgcP/t9dqjusRgh3WduwNIn5h68NU7zOjmiifGsqQ+Bnm2CVZ1gJ8yHQwad1ZxwuiHM
8EYH5XeJTvcXPRz1vIJqIY1gZ8JB2lraqyIFgo05yO/T+sknXjTmY4Xk0EvjocALSti2tzRuKXmn
l/AXIfKjuJ2aTPuEl9tSHiHu3VewK9BZvylhPZAp0hBFABtAbVxYdinjznL3n6DALGCrQlSmQ/N2
dBHghLmWhMn/xEVNd/3WI50O8yOKDbplzp/mxY+ShA3UTUZraRI0hS9kQdfoNPQ++GOTL/lIjVMA
KHWjmO91G9h2wY3SDmT2B/X8JT/TtbjvjdSHMJ/62hVnesyde49sTcjXwbHr4FfSxArQhua+km2A
3jlFpufGN5N24Yc0Xdl8X5mS2mat61MHpBnyzC53C7umGDa+UT6qA/myWzFPJ4L6Waz3ZK0WWuju
Nqoy4TqPqkAC7jNAQwc7HJsyIcOopDWn1sPNBn7dV4dSfnDFPY6OsEKq+sHsKiXt6+YESy7SxMID
t6SLj4EbWoKNNhLYK8T/OALllr5IipMAgH+f/ICNMY5VJLyREJDiCE9DdpF8yj8Lx+2dCTSbchsb
HliiwpIbD24HwGqzCwh0Ry3YuHb3YZWQgOipWAip2uhGZKcuonpsLAj/+mub/3/+1NhrWnGOQgwU
N8AvMeoOwGNlOEsg6nbcEbS5VYHrpFtxe1/sSzZtQfiuKc7F2XAR1vVWuYP8/sK55P+XxM8uZLtk
6fdlPV7rBQC790JYOfqTikwKSIf1OYF3GfQgTqGzWre4oo+2khl5RX9HMqGefjXoWqpDm+OMse0d
jvV65QqC6Cxl/NeANye51+y58hxLBQO7cCjFB1Bf1g0ZkaAcrTYv/YU8Hs+84VxpUhYavMHstyX/
OvX4ZbSrr8cJvpSPCkxpV7Cwk9GYTpPzE7EleiLWNMSz1o6LKZGXyNY26kfX3L885Jk1eJs4yRMk
82UVDoVZHLMm6BHNoyeiOYQ80DBywsAQ/RYdJMcP4Yxrer8igWvwcecL9AmyK4djsvTkcUbjqcWW
T++WAsVaYYZREsUaVSrphhlPLAF1RKp0Lmvi/R9M47t6gdBtXnq3uAJ2AQ1wT2ffLt2bsoYv+UET
A9iiXnvzncVlRze+aSoUiTID7L71AyzkR5V40zJr+fuFjfQHD8PynUesX6RGeZoEtKPrGBI/z86r
YlGWTsDGdL8dK8p3t2KDdPdAuKCL+a/mX0NFwVAZpVN4b90g0ZaXeDN20Bp7sRgzMIHxJ0F38nxB
ZCJfiIzrwkbXt6bL4N8KThmaM3O3spC5jJEUn6xMsU91Gg6w67/0Yx2cNTVFSQBHc27NASDWNk97
toVo5q2QmgPgCLK24n+X3Xqkky6440DIufNjqIWY0kpn+uxtK8Gf7bEea8vnzgeBh0eeQ6Rs8z5S
YuTlIRdHpjKMZKXRsTaabt1c7ryppm0/UrXTPuMklpXDLbwuIuth9Y64wYit+ZWUTiqJGiVNja0/
iVnHjUNfBRctUSmuhdooglMbLbVovzrglj6pBD8o3qv6WhQn9zClWYG5yyFFGSdW10ROFazycfgc
yBmw4DZaQnMatugqzhvHP1F+dLb8mhi7T9h5oT+YRmWZK2IoLc3mtUVk238Yb3AkMjiXUfTSAgva
C85wUDE3AfdkcmXxPVNpwQSsy6L6fqe7J26cKFccmVeJuTg7Gwri31Ce1DkgYpaWRGXiv40QAWmT
+TOmd+h8I06eUW7X/RxhyM1FpVDfeNssltRDjfOg0vFZCc4fecK6iujSu3H9cxSjncwN4ntA91WD
1rbZs68tjI0+MUmDAd+idrb9ZLxIYmGI5KlLpj72CagrjZ1G9jhHQs4knbG+l5sZ//E8A5F+17Kj
bhGRtK7GZLurGws9F/vUuXNztBD9VNgjdC6W6O7qBASU959b8pSbhxLtOqZs+/WXX698Fqbl92Ep
wNwIm1HgJ8tFWHInOQJSUKhIzPTS8z1qL7rcxkNAlj1C6+7YkuTYkHCrDXsjuKmFV8GU47JG3PDV
su6jj7qL5OsF3g/N8fY1gMXfkeUs/KMxmZTmHbrrJCfMUDuCJ1UmY6NwNazsSa5t2s2BhmJ9CwU4
x9y0yGIxi0dpf/fknayy9+qPPKfBn2TqeI/ZY49qGOaliAYLvt7rzXXT5VDiiHKIJg2kyTwUDmAK
kMr2t0LEu5P+J+oBQdcdGvImbgv58WW3xlaN0XA1FOg0IwK/BH/FgaGa8pw+Uaznto979ytONVwW
VbMk3AlXBJsbjL815N1XTslxMDaENSWppbfRoTyETFPXSvKdZGF30BFmtBDYj42eUeW/PEy/PPcD
16lcL/HYALQIFDXJjn8gFKPhKUb6Zn0LKPA++S4dFXwvQKXxX7BKrn3myIbsXtpv+y5Mg5tsygeI
Z9dYjUH58GXxJdUI+BP9yq9+Vio0T/0bpVj+Y/U8e1m7YlEvIkNyDOQp+Odzhfm0wdKPxcjsqlEc
r/UX9b/xP9Z8klPKVG6UcQroQLVtIWs1pP8Pp5G5a534CGULgncF7cm11EZ6fso5P631lhHauyPe
FhcAYUUvWgc07VDpMdGb52JzpwAPEbI2yduAdabtt7p7uF8kpYIRj3yLznR7O+jch9FQ/Aa5Bqms
4z5y7ZDHaMwTh3vVbJpXsp4gzD5cjK+qNn9ud3y3kY4HBjbCx0AZMhnyPbNuKczamdTrl4WNnYtq
QBbEiORc2XVd0RKa/Y/gg4Mhz+UL85XZp4+0iIhrVlnR4auaOraspTRQmaBz3UhX7vf5aWThQ4Nh
I6OFzrfnGzmNuP4vdgpBx+7nscu+6VHNjpJcaOtndPDhP6WBoObUqUtNDK07bu2jdGXCf1V1XM4C
UlhQ0cmsk65+7LZeuo8zWQIJIkfWyomRo7LyQvOn5PxKPw2b/U0lrWVD2CHzABhXMoGe3Je9G0JT
ZxKf1c1SsoeHIeATkXTclO/8hLCtl2MpXpPRtOyuHjYYq8Ru7gaeYNYH3IutizAttU6N1H/x0iRi
t7y7KEKYG0P91Gj5eWq8KMqCXaiGXAToMjzq+2pvPqJgVOS6mz7kxXObq2axk/dAqxp0ikBoV2II
p4jT3PXziBMLv1aIGHX21ONgNS35j7Id88EL2VP7BbR2dEilBhkb8nJK20xUpS3RQVLA1isrskGF
W426g1zsXKQAfPktq18RDUWeyKp0fQ8oI74j50yf37Ho89W0W8wLXAX4bSk4fWOWV5QI+6OB/bEk
LW5dhSx+j9Qu4gTjMuyMsybsbrX0j7zRni/xrBUm7wjMvWceE6YDI5zijM+9zuISxi46IQOz5lGA
XmdHlq1iKBZg6HJ8IhRzpC82yvELoBSywr87v1yxzLjzH5I8K3FS4FKCe6K7ntf1/HOtROMXpJL1
jejOFglHdLlBLNMfvb/zjrt8SY6mnVCwXYId4urGkV67X9x5ey1DXGrbjYzKB+/OAwBIQPc6uhPJ
ji9jKS5MVDFN73anLPjRcu+L6Tw2SI1vOeqGrbQb1blJLkQzpPFABUSI1PE2qmD0joZcKRp/R+V9
yEmRHdzLY9a+0ygYpPT5MAqyHcNOFyR3YDSudaHXXj8YAMuVR/7rY3JIKFsNwLGr8q3r2yisGTWU
VVukwVsRDd37IADLNV2Of2lKy52uEpM7upEvUxJwCxQSDGAVIDBEQLvhkWwkpZl70VuJEfZnz6HI
sZ9EseNbEU+HrLi/a8pYDluJp2VPQm4uqgDb8DmTMw5cS/0+0uWm5b/MlG3EEDfYzoO4AjvruhGV
vvdn/GDCPWUw71gTqm/O6rOB0WzR4MTz/dVRQAGpAZ1GxJrPr+2M40ERdCiCORzVq6ORmqxpGZ4b
K2NlK3iRenmp7eh3j2L+yfJrVoH4m+jSIxOYA1ZklImm0gVHkbJIzQXeZhStk1aqe8L4JoVNRZDS
O6c4uiblIErXcyi3TgX2Bt++MExTv6z3uBJ5DZdAwoZzEEiYWW3t7+PGSIXcLt+yJU7iP79zupVP
xOSsUFCTZTJH+8nK1KHdEKHD0sc9ltJio8l5kw5SijFRMHaBVAGbimNCnxAR2aibj8ch3mbyVEJA
86rdY/MV9etn/+FzsfQPzTGPMfOoRB/5S4rjAqRHHF7G7T1rSKjUbs8qc/lXahLL0F9cSxpwNM+J
d6KSnaKu1jtTaYbT0/Ajs4oFGuTGHkVGvRv4pgnufoSDZLL6+2RLEv+Yurs0Ed38yw8qbhhesM6Y
dNGKY6UP3ClwAzHCZNLMT3j82aKQ1kbwwKtuH8/997khqZ9O9k575eP7BMP3dIqkNM4hFKi6c3YR
Aekb6YJgEERZ27jf/YVYoQmHfnk3safmZf2ebdXBKVrwosZZoV0uHxuJVAVrSI0z5bTEbdXp84NL
C0SkHsIncarLBEa4xm8+5Yvi7IeIwPOTGn/rP8gMRFyIu8SEyppQsy0O2uwyuxyTVc0h6BKTh4Hb
z9V3PXFf3VYe6gVjQhB8bgzDsiiRSlLbg6tnKwa7qswJo+UNqKdao9+syh3WjqhmSm1VbJ3UzqAJ
AYrmC67IOafokzXdtQurk0m9FswXZFhH57R9tbL38FVp4PMt4My0ryacaQfCzWwnY2tu8ABwsa1P
DfFMxTtjbBIlQxQSOIJ/b0Abhi1bO4R+ObbgZRGR+vdebrjFAkn9UGTt7E4Ao/K9nlYHF9nvBu4A
xD0N9d3idrbXxOkMuBa0dUPgyCNOFNM7EOCrBgdHn1Z+mlRzFdSY8lz1q8o5J/9Uy58e21Mx2GaB
9cGx+bYvefTHyYIt+lWQ9ueUxX93T7giPKu7uDiRFfJWKhUNQdFilw8ob5NT5cJSwxnosPlrMJIY
F5qZKCBTC9aBZ3Am+k4CG2Z3/3eeMFHkOBkqA0hAUaJP4A2s2GztbqWhs+BIO4azMz4N/+GGxME2
5Q3Rm82avuX0W4HJHfdQHZu0KMMrkHVVenTqIsmGAjiT4Uv1EQgL7chSHBjx7ukWcW9JOMUztX0I
WFGXOPxNAqC84RIV6GxcfEgaG+V5F8FM4mI23RyBy+1iiblW7skN7jiUBMwCCCzjP6SRf4tBUJOt
bjp5NHneo0BWrvsHyhOvwYt04+M5aTHhjq4XfOxj0PvGMpq/HJ7UBG5EnXXCv/KR7CzO4dt8kDrN
Z5ZJF8q86tPOCrFUVp8+uu2eG8FBr11Ygz4Kin04lF6/ZqnvnyLKhgwk8bwcCvZBVXKep6Llr3n0
ULblBe8gqGXqTLjMh97EIXWqKqUqKj8wkBgGrBGse+CpghZvPmpJwDp8i1hExI4yehFCZCFjIpwS
EgqrwLX2QBeqgvXZYxZsQCUflrGov68UzwFZ8eex5EDfnporJW4RNuzo/14ExwBm9bdeUL/rjll+
928jIiJVVnlSJKIpqqPEY8C4A05i2T8+M5aXgETICymKn+HnS0xzrX0rs1MMpxJPMmtXCm+UP7BY
nRtaT7QaBrcNdIUjWTcRIU/1S6O0E869o+QY0txIsOGheiRmXY1PdKxs3A0vPuv10UYNjsRNst/u
mtzLjrXqVy3yNvvZGZOjqesy1qmxtCUqY5II+GHE9Djv/oLZ1n5IAL4YDl4lBDGqux9/bAApfy/g
bx98Vfkq9ffb07tD80MktMRa6I4aGCmKfAvc9tfsUlILq/m0ev8/MzBof25KhH29Mn0aF8oK+inZ
v4ibNqf9uREYxVH428uhdPiq/qB0QtDUhdYFr+dRTLBr2gqqMuFQ/0sJM0k2Kpjx99Q0264Thb53
qMzodOG0NU7jbYfn7TbZmsAkKazCv9psB7GCVbp4ujeBRECXKAWccu7tWnUQ3c6Rz/qrAR+v6BcD
6Te4XJFNIhi83ysQfT+6vHJ5Gl87ZfI68muoLbxUytVqlcrizQzN5aRcTzSnQWZMuiBtghs6wnGP
EErOBjYKRTn1FTk6AHMyYuIssqLo+e9gGfi4oWEmxIX94T6id1dwYnLmdZp2slwwbGEj6xkq9yMQ
coVK5LtCkyLKigA0mcCVrRABNORZAo/V1Sxcu/PH79Cyuip3a2nNv4yh6xoQ9uQu8F5hVxIhHOTE
QlBkt6AM3PAEDT8q5/8OY4Q2rRdgUrUY7bWAinBB4jUnFXF8u6ix1Mohx6RWZN+yEE0z+7cYrcqk
NK26cCpDuj2Ak+UjYXPtyJsNs0Yp9pZMeDFx2yq1+34Ds9J+ZGOjCsv1zaaYGEN/aNW4Efu/pzSy
BQQ6uNpt3VJNHgs2iiw/hkJWtVGG7EpBDtIKZ8/955ioO7RMuSAIsyhIyvgY8QdFRzmLL+HVKSCj
TPCN1ASL1Vn1m+E7pQsr1ePgk1mHeVvxDsJxugEzFhEzWI6rggjLEDduJ0LN/YP6rfCUeRuw0b18
249ctycNEXbalk17ZONywKvNThLpPGZmrGZND8MQL8Hr8Br5NEofzf/BGCVS1HtU4urG9h7j7+i+
54NC/aIIij89BM+DFKBGXFb9FwOjKONJQ9vBjq1pSkekRi4Bj0TDR6sJoyWHqXTde7hItff3s+H4
daBwjTbbF26m2HtlM6ZLgjy1Mu3pTk3kAANIWYXkTDpghNjgU3gyobryv02X/+5HkTVS6Qdu0okB
9MuKQOTpJCGUlQwn3pVYnaAVpWC3wJiwlz/Pljro/8x3L+TGxhptTqVMaf11OhaF5e9VSvMrO/vG
1JQq66PC/wiyakJJBPuUUQ4hkPqx6dMr+9Rieh1ILhiqjxqlipVoH7hQX+v53QvJYF0DZUxCgzXY
LBm0/fUu0yA+ddqiXjf0QuDRPK7isV80283yC3zYyBbdJNutb4romM5IQtByOmvbco+xu3wxBFCE
udAdkuYQYIwLPxn0mjwRw4Oh4MvabZHd8HoiZ/19WE2X+RnjtOM1j7kF/s7eZQchUMzOQGryBhDj
v8+tv7uNjp/yxYWtdR4whdDOEYwvH+AycQyRufSU8pl4As2s7HR61NwT1VHXeV2SrjC8LAoEEONo
DkQfR2hSth8LT7MJvNoX4wYN8IXMk8elOtEwAAmyahgcB5ZSt/ZBbCrHU1TBLAN2SyHfVU3aU7x7
wiN/1NDcvQUEBVYnUc1CJ/j2Yovkb4CLjTtX/vRjjtATycqoIrVK/U6xLY8mBZqKUlbB/fvb+uSC
XGD0xuoAjvoUOyzFLXXsighQ+H96NM8Z2TJ0KACb9g1YwhH4L3eBUXjqihiaPK49we8zRs+kFKxg
xDK085LGAamTfZ3BgzTZ5jbLUHwH+gZfDd+QX9K+v4cFLdsAc73+sDUhTA4qJTSczZAKrz1yMiSB
c0Ax6pA+RLLwN7SQFZJ/bVWISm9O3gJjUYc+ocl8Xn7U8jZMtSymSbdQenRr9oH8a8nymrbIi9o1
2lojfw2ON+XgzzJdQyiQz7LqWYlN0osE7OnfUhaSlNgLOkzlLPU4AlnhqODhqGyA1gB+XFzBJRW+
RWdcvBgDEefjCdiG9UIJ0fLUeL5XF3I6GgHAiZqSBXWp1UAld3V97h36A4TlOUD8ir5ufXlejdap
o2qc9MUJ+IBKs4SfuOFDCcusRsvlx7F+sBMfZVXmor4BOdnTtsA131uCjAXyl1+4J3bxRXMHQCVb
2ZZivXo+FnLfOfNJ2yYdjT9w2r0OEEdwhqhIiHZzIjLShK+Z2y1zRbzI9bFaDV3J9y0NVxTexLcv
s0RjdIoo/BK04W8hlcug5eDRfnnpBWQZQ1VC5A4uDhBV6Bm9I53lNG6BmYHoWiRr6eKFgTmLdzYL
UssTDnUshL/DvaUGqP+4/dZxT5IyWeeqZ6Hs0t3NKz0ZiFTg6/2DRpJ6PhQ3U4iUVUyNQIwXN6B7
Ec13Y9VX89LBXpIuctLDyaDv7oLFcQCGJ3gSLZ273utfXG6rZkAq8V2iPLVGRWeC0EXHmEnGF/pC
/Eko9C1wc8qhrJfJagUMZa0zNXVEp7hQAn8/qY3M1P/I083tGdFe5cS07E218kfH6jUHKWyiqCgJ
y3T37zdt+l1KTueBGG3f6wuYv6pB4m0sgRMrBD+LaedptdSrvexTrrwIPYYAQ70FpouDmro183DI
vZnJr5zk20FZY3PJrjnrfSAgQodSatxEVqqKuhum/gFzAjUlFrpkodwrc+JFeE8ys/9mAU3HeF/K
hUka/P+Vz8sJW135OGzg6nptqROFGMnPgFYzmZfCmDR5oY9uKJvC/BcJuXmfzVA00+wLg3o8E0q6
ENqr2qzhGXguveSHGPYw1KibY44oE/JCVxQ28yE08I3nIt0Lo3uYRrLP1Xb0MG0D/7FYjO4JL8Tv
lggWLXUtBstJbECdFpmKmKvtu7sAfcT5oDBP9/5L/FJfAl0unu8Qv/CXhygNqx4fu/MiHiR47yb9
1wj3xdZ5V668XbcLIy7S351i49u+mjHRYJ10u+QaOAetdoQ04252j2V4LhvHP0wv90qa0+IgBNwa
KNfiBMtEVuz25UvME4aqxHmPmxGcKsRjDfYcDBDNDXwnrcFYijzL48xZd9wQq4pMK/VqgF3ychg8
YuEyRn3ZJVDMRevG8EcUm2V5aF7IH28ojA0z43+44GLxquy2yaUDGY5sb21QvnZHRXgVwF+kWkwJ
q6jpt58VLvv7SsSWw7p0BgSrKitX16Lsrgj3nO/RnemXdHSG83dm2Pz6dEkaQGV1Ep7Szjdb6L/3
/2dEce4e7L+YAxdMHRzMdAAqG1IlgzNGEEokzHsHT8nw4fz5kjF0cbTcDsGUFbJPvh6VZsEFonER
cnHsuBIDSyMRI9/sjNbYm1RRWa+bE2sBUyLntaj/0Db37KvOadeJIL7JyEFlM2uCSIpcN5tGS403
TZwh+X9wISdz07DTZS/UO69fVW8hhHliMKyM3kdlUHGqXjitA1ZmYt/hs3AAztJY1u+jRSS4I/H6
BU9Nz42YI1liSYyhcUi7DCuFnU/STHONgNW476nY9DJOPqFytKBLuLqTTTqXDgywQscSC9SQMtoX
LlHScrfa6WhjEAnwOLOqj9Ct96K1UEe7DgVSL/iAqw4TNK74s4Twz26LcHuLabpkVw34ETormNPn
GIPKEgWHCBxqvIsAjD02XB/4Q4hWwPszqX53Ld2ugfEa+M/O//6K8J7zjZada+RJsIKSo+fdGMo9
J+/4S9ALw8tz9Oze9gLhS3xSN23voehGOF96S6DG8d6gB58V2JPWwE5frpwA5gZ3Gfi9zniK2zQX
HJDbYjh23U6Z5kBquLpdnGOyJ6mjfdeJBDbRjfPrvDbO/VDganrw6kzqoFZVBz52jjTY7Yf9t5Dr
x9aWEXU9ahjBM6Zbtjrh3r7D22E5xZX1zHz7TZ6mHBdvlsKu4zXhC3euVZLlgF3YsN2iKVPe/tHG
EVjOnXPGsvA3KSH/MEfCzIGDN1fL/E+E/PFnMdEKnKeu1vhtE8nwLisYbeQHj1QPnr7IeXNVDDQ7
/cQwib3s0B16Ggt6hNkMEIJBpWGKTXrDPSJtrVsiXiBBz/2zIzCLhdDDYSWWNi1eMaE1jSblTtKp
MpTlqjtswY78XiemcWPFIAcC21EgfDyZTcT1BsvWO6sQvi3FUHfPZWUHEC3cC6dAzRbJ/iqTsbw6
kVAqhofa+so2Y5pfPzCK0KSIJc1UY3rMvW9IwNL4uMl3KGj5LA8aZImyvzCd90SuIOz07LgJ+rYS
I2Jap1AMW67Dc0dPGrFm5O/b6JYw50DyIr53PnZVz8FyirpHEwvino8voTlCVkvxvFyHCZf3CIcf
5jmLq62J8YIoWkIKj019SiySmumrykLtt37v9KLhWTfzVOUCjRWkejMCqc3nRImlSqfxDjNX6hgg
rSaW5uVSeikjBj3x30lofd1L7WZqKQu6jwkSlKc2Lx/lV5jUlEpx/rQEy1LKIs/rxg7REOgPl40o
Dg2rkEITxXjrXcemuXhB2f+y4r0LdN7Ae+X+7BSnZlOYuJQmWpOVaIY9kkrIA9b6nekqqLLxpeJw
IPuilIgUYC5uggzKlMv0V8Y6lpOIXtt9OM2ATwai+TZXRFZJCMlUETRWoihHMP4hAj8Rk9Ken6kS
eJUPD7ceu7NFfSBnlMpcoYbxWeFJ+FZ+PdSIqu9w5vPHjGrXqe0JxHlE72ZyvyY2Yb7ZzA0ab4Kv
bsvBKU3JE4pIPtFWGRHF4xFjKzpBjaahIr8B+YBMk+SGqNvZ6KZL+TRXdJgnzo6rHCeNEbMye6oA
cHmmpx3nzzM8eLiZGtGmfAM3PZDmxCjB068EeOACvZTPd6AQRuS20P5LWR2kUGs/abiqKcibI5O2
P7wqKnMzrLGw5u3Qcy8p3cwhCpq3I7FjL3oNvCrjduuRwGzMKBuDiEEt+vv12QV7UXKsZqb08JL4
AnaGpbnserkar1xyrWYZW+zeKPKf32Q9d63EN+K4Q+l1zwaRfuA1cUCQdqOKIqT9uMKddhKniCH+
dvFiqOWBpa8iPaMMfWdeREhyc4FMmd6LeogV4V+Kz9OBuwL/n9Q+YYH4aCbqBgKoulLxl30tjMlg
vH6GlgK6jrLrnoDWlbf41eQ1wYKbmC38ftg9cISYYu6xSFjem/wAe28AeKwSZr93e7baD3vhyNtv
iPvEqsZrX1dys0fs5Z0FWjPSnm1OYWgE4inO9whL6XsI3RVE01UzHPgCOnm7LQUl9ycwQWRZvib8
VT/PN1b+JmJbr6kRdgahBGXLOZergX3zeZVvIMUIE9ZTCyxZCmw3aJwY0VgRnxEEsUlqaOQJs4UK
idoc6+TZbIj59V0SFZ4r5mBSosGggYFo1cxu0lZl7/WYlCreLqu6ZnYRJluHz3DPVuNr1+roalXm
LvJ1GZP+QDZ4ubmgpByO7tK85Ha03CBEr+YqR26877rD3wsoMXCQPOfnG/O2Yw5z9aYOxmQBb/2L
0bIoEHYMokz0Jw+BKKfAHwpkDc4XtC62Uh9Q4KWbTO7YLtLqCCscgylxTjcSuyimVDSOHKhPDxHV
wmLJbYoEynnAnr8PX2OJQ+jxdVEZWmEi4FVNqYDbucWTrKSYj67RkzIZvxdKWDk/Se3ykzvDupvt
GPvqqC1lAPp43nawWj9UmguxJkAtkSAH0z6Iz81Hd9C1RTndykdiLc+Ea7MR4KW0Xoqr5RsJ6s3k
jJd2HNP2Kva1cxwmvQjslNpYs3JjEqi2k/LCoRItRo0u8TMgOrk7MgK4avYLcD/RnT0VeSak7n3w
Q+OnP2JoUefdGSeTrHkzLNGNBj3amVYNaYbLLdaqjHpM9VkZ5ZfmLhRwchQkvW1CGmt471pgHtri
XU3iZsKihnhddVkzxosLZbke+ONc2lh5AyquOmGqHgTKdXNWcGqcPfVKX9po+0pkzo40OWViLE+s
w9NKJ2A79B+CzmGxVj5vb5lNctwoxtQDrOMF3ljg1pFdy/OPfX1zzCIxTXZGbdeL13uyg1iDZcMF
xYXZZBMnacH/UcLf5OeepWx7B+z65cTvrJ7WhK4PeIAwZm3n4dj5lIz2TKAxf5d6JS6gRB1jRy9t
RaFSf3GgWYZ4kBYlDVHwWtHuUreo1YMtFwWg5b3LoBQPnSNMoD5fVWO1zM1gPswA8Du2Lyiwn8J0
jEASMJQC0BJrABq2IgGYYThqy+t3xqa7nZDfH/hCHTGn3nAHEVMMgbdsiEC206gj4epGZjLZ77Bm
VixEcpKw58BrB1fO0Rd1SHHq0jRxH9lLLbpMzFCvF4JhrnOxzu7+xHEppqPh3FD0XE09WEjqNbpN
nW2MrtW/fnUtwsuxFUBbh6iWP5dpCUPTmsDCOjE0MqKDXhdRxLZfQ3ZwATItAehE0KYFtsj8uFAv
LWhUWuwhHyxjdtX80AcK34y1411fx0LWPzuDRYST0w8lQyR1gWjHTQxCJiEiBzUnaM2+wmaGERns
YjlBF+9SxHyeTY+tzBGEKcZ4qr3B8in1eqMnIuk61dNO9TgZYuLvFWsClzJruxWJQahSLVQQBFwA
o4NSkoHx9UG5HdAZZ+bLuh8w3CbZExbanFgR49m9zCUfAVJkQSGUSTa/rGmU+MXnPkRIusVRXDsJ
poAWKjD17k/P7sYfr+PjZDiGqNoJe0Dmyy7LF1MfdAahkbJ1d4HOZgfWe6FwhDW0ma+RqDIRv76Z
SectyS82ttb/ZP1RkBwwwLorqG7jeQRkDjLBNApQ3LopwDSzfzVxhLuAOKrnXs2E00pyzknncxU5
DVx1YTp4R/t4ecnrDTgiO2hDJroawII9sWuedPbgDAX3uJM8r9YQrh/wfLHdnLh0CISpJiMZLbFA
7TKCIO2h44D7OjoW9xcLTqnJrN2TfU8r9RBFd8zAH8WBbkEIavmpwe8WCqRrwunRx0SarwksE68m
TzCdCU4ss2vD2A5uqMmf/Vk0m96dHKHUfCpAhIWwRBfwWXPPL7zKk8CYg8gtPTgeBlCWCcm4QPIw
FagcLvRgdGn9uFZGnjZXRy2CFGoQHCY6LEWlNmz8F8St6ILXzgYFdHfSzPLr1CrwxwI+iZD5g1Do
awogTfGs7rNxTQsHIRJCB0+s+9Ofr+m/IikF4zrw9dN5mkznEOQ7GSBlpXh1h/4Fp+O4pmxSQtVK
d/TL8qk4UgTET+Love/vlQ7ErLlnGBCBqJYXUzQ7rVAGOG5MAz+NXfikjXLJIvXdR8cMqUpYqNuu
E/qtO09DQ5SQBF1M7qc/jMkey032IhKD5xJHibqvUBuUG7VPxcO+kxkLjVztU3c+FaltU59uEXus
leKMdOaCMHDkbdHhg4eM3k2tQOvrE35tLBPMRQTjtl+NByRWBiyw8laJiiE3KM1wmVy3arkvNMXo
/dCiNytnpsoyPT8ZQSbU7zpi+DWeJwLs14qU0FH0nO24njlEofkMkL0u3908sWF7zg1WfIYXIvEQ
c/a06MX+KR70lGmJFo/l813nYLJQgqDj7wMnAnqpei/4H7S4vDXWn3lOxTngHNYZA8gWmj9eplZp
VyU8ezNgbNYNDwZfC+1ls+SQZmq7qGw97VpQSH5taC2IzWtb4m9U1RChM1t2WvK8xkahn6IDQ83J
oj0TVXEaRnsCOIpLiWw0xgFtHnEm5nV/IGfHlpeu4iv7wjagYpJM/XPld4SEC9fE98pI4sBNKDET
6tfq5MLXxMD9BVYxqiWPmHsL88cv9hB+SwYr0K+HUb9qLsd7EqzA0ghnqxmgNY9IKprVvrgY3UJz
Gi4wwIpDUXKOxBxUrF0aO0Mtjy2SyKLrVraEQiz6XUDpraXlPNn0VHSeqDamDASVx6ixHBwJuAI6
NIH1uGmM0nojfYN9sMqRMe9HZgEbw3HMTOsOKUXYbbbDkLrdWfwcqvWQMql2Oic82QmEPXeND48S
rleZPWBc/rT5K7FUNVenHtzhWY2V5QV0S0GR6HFY+UHkHdRAGuw9P9OtFCFgZ6jVFGFgm0Pwju4+
QzQ0MwMVm9wEC/lljeewGL+wpTv38k9Nkhx//AMQYJz2/mmD1SZ4XFSaGHnd3OTPQyt+lbYB9Jep
c3mywvYybjZfya8d/cQXvnJNGpyrWo4JEmZF8xu6ojfPXvk7jgPRUAD/HFAXwg6Ui52Sbc5g7nGt
i2uEViTYQrTpquxbci1I5qOIupOgLP6iANVu5sq88s+Do5Ah/9uTG/Vmr5OgNIar2Gkql0EQPWXz
pxTYtmdB7BQs5J477fCvAiV72jyGz3DO7CqJTn5ynNjNUKZknNzk4pWg4AuoqBXwFRBlt5o2LqNF
l+xJpfL8Nko/sdWMFrdw0yDrC6DpWmGhr9VbXIJJ6awU7U4zy3b8c23tGQXDa8LhY+zp4i+nwKCJ
iHz3bLEF8FiBaleg+s4jcgwhCdyR0wnPk35em67U/5833o1yg0BoKkeFzkoAbLqHjcZyiCJmXwy5
alrQujFNp4jpDAcYC9+mSiPrQJ8EQUPcqdQDZhrk2q4AqAexf8ieQQLvADN4T8E0s+aOPyPOgeIk
p3GBoPGIOS0io4OywzmaXpargRmR7rhPFkKDY86vT+pm3BH6Y+DbOG/gIQ+tVhCMks/9g9HI8Vc5
GgySPDufwTxBZ73t/mLhFKzB2LSXJvBVMskmx6PE3BiRDfUySCMvI4wa2adN9w/LlVegBi8W/501
R6bZxnJkQZ3D5ysyT1ip97qmLQD6nw+a+L3hiBY5xrVxs0ZxBWn5SmTbz294XXPygBSaLv2kGH/4
rKq4Hxj5DpzAj/kFDqseqFAKymk0iR/Ln0Iuqg078StjEvkH0rV3YdJkdUYOQLV4nCkxxtm8d/0w
qybFq3xdd4nKQEQzEHHdbAahS6DUSvkSoviNy4VKSxsNcHzGn7ILCRFUV3+C9nC9bYhKjNv1uoPy
3dXfCniqiEfiCi1ajBwJTVFwW3pXgJQ856tlObhPmhTPHAjntO6acbFgtHXiOJKKHvfAOOUk1RGi
BSheHKAXEohqsTipoG9aDNqy6A3Ec7PCV17ITxEzSB4ugZ84kN7RfPtvwpdWcxVnhk7vU0CHF92N
VfEKOI0TIV/sWejEDT8umEHL1oo9WmFcH4fk1E3m/vWXa8vzd4RP2GIhbo9/RkxxR/jehvcO+orV
AY9KnROJ0FqWrEQuPj1oUApaSLYn3u/kQTqctMDiB/cD1YH5geENEJJF9kr7w/aVCd2soAPTWHsO
Z1TDXCULlOUyQ1+1VtxOq+Fuo+JXEJ2khJ8C4Ru5QL69BCrL4AuEaGy/+n6I31sZoorB/f3CpCh4
EwJGFKk0WJNrvKFbBEAyxxcP/ApgoUoborp3OYdK+/ZuLpfgVw2P+bVC5KIbLEzGQbM5iDADLn/T
iKYL+RgixL+EgBinBOnXAAnIknQLzw10d/9SjZlKoIBjsytsCPgWaQjnxj6U0PwZFQJU0Zs98Zlp
R0tAD0jV9Bz0SN7RyH1dAjClXevieSNPfjmOO44QlhJVEQHdIBN3VJnrEsrXd1LI8ArfenMmrpCP
Lp0zekQ2d0n4ln0HuCoZF9zmSyH3y9iHk/Nv+O9MUMgpIFQqIv0gj9wJwddiYXlTCPZk1u03evvQ
4SRpc4s8wR7pH1DrjPK5H9EPLA15zS6K7+rAHrgt58ziussyFs3ES8DqRqQkkYfey1zUR3lfH+qT
c/D5MzJwwWlKmpp7UvmcVVyrWVo5NVbIDRmkeVSKEGvZUfK1fqTMydGpDhdRgObFP3XZvyEiIuPa
QH5LSGEVPu4re1st0jDAtiHZD4kB6ePsjVJcagaekV0nvpZERxdnADx1q/HbGkDmIrpxYJJd6vlR
zgYecALwiZNH16+Mvd4v7LDVFLe5C8OYdNVcNWkrU1CdyEUBKgCNFZTfs+7BbALUHm4xnG1rT7+P
LKQJw4Zc8DBnrpuYbETUU5jFdpY6AlDy4cWTkfUCJPFrXdKqucNWQjfbHk1S3wA8wz6Rcsb04AsW
axOjrgsnni1OJ2L0BHFbi0nLVa1pGH/p9dLe75nwR98+TYIHQvazjtJZ3G9uEExrEbCvHGf/Tm+i
KmGETNNiI4k4IXBXNlkhFNgBiAEtVYbCgByxVvQz5Genu+RVfAY+krFDKRYA1jdomTcUaO8oea/+
J3lVhshkd8vmpR7MhGU1xkML6oZie044I5yOaYtqEHRqVswg14dPGfw72/O/rzyPvGD3VTpWby4i
U9E9NStp62qYl7jbfvksJJ5fWiZR+zHz2aW6WAcmeUOi1opeVS1IUZdOZzgHld8tUx1QUnJLVEq2
sq3wryC+cwkRyFJkUvkbNNeWol8QdpbG6XbRoqt1AndzJiBU3B4XirOx++1Y7GnBfHRIYWsFkqxh
xolszbq5z3QgwOO9RdMCxnERC61uhvh5eZB7RxkBOZkv/fcDhPUW663gEUoKrmoSRGgbrEvr9Q2e
AhjxrFS5+IX1a0ih1aNT9VUTI+YKx37oBBXFDVo7KmsvuHwOVpQC9vkv0Yku+SWMPpYv1sX6Me0B
TcKCTpV0+N5S/ZdN+QlLz7GlOcmgDYyqvZ/P8gVlfMZD5YVsrMWU1dshfpN7v7tvoLW6kgOJCQV+
xdbVE3LrIzPyZXatm8SYW0M3GO/pgDoXc53QYL/x4ruWi7lsmtojvjiqv+LW/5txcum2xXCRLZie
iDK/WcQmeFSiZhdEw6STg7r15IgHLbtUoRn3KF6myqM+GgFYOfeVqYoX9YILpYVii6aszDgMjKNL
tgqFM68RFrCHZTMYE1IlLZ5bEkkXMChAhcJm31uO8YbghiuoFX2cguzGruhbYJCntuSmX8k2d2Me
raxpovFxQbLNZkvra+qi10To5mCXSLPWyJn/9HL69BVxYWzAnb9dxLZGiOiP+XHBhepruolFDaJq
UC4kHfI1nqQbnOgQunpzY/mr+J/uzgypraHL+IkoZEdRPrf2dqy3AOLT+0Yr8fTPKmCaN/Xp7gSe
pu4ecNdjMiZu/d5c6+KzEeo8tAyhFOfrDpMBOuGME2ddm+zoNARPtMUSoaQAHMWEzD3Byed175Nk
dMIHMUUXqj56Ru+kSfU4H2L/NhiilQqJYkiM7bKJxbl6OT5biVjjG/27tA50N0U6NxNGxDlC4elk
esw6UETaMnkMufs41PIJQL5NTCdsee4hyrEXJrDHZCnuYLh8qBPF/sBRz/bzlF8BiS1um4/IM82r
JAhMeIdSD5S9ipg4OPAc5hx681V8AiXIINBy4Jb/WFJxgqfdLZ1dJOFMJA9F+gx3iz6O9Y9BE8kl
TmKu7b8PFcncnG/teL0dAWK5eRgRO6vPefvjED6u3/7MN3E6QEhhHcUSen/OkFqvVJ1kgDqGSRg2
Np4JVdmwGkXUHMF3H2D/26ubagMIbFkCE3lHucOb/rsBH7KG8/tj7yundx7BpDiA1qAgo+irxfz/
6Q/rOoPrPVoVHjc94rTIaNijRr11cdJcu5QtnEJkAFsOJ7ZYj1nOO61BoW0s8QxVikn+OBko+E1b
guR3RiJD9fQ5vKgu2gzI50cf4YspsTiJNeiSO2Bn9N8IzqsauMK7IrbkSsPnaH9PfX/1GdtM86FJ
yqD8KIdPGHs+qzdxQyYfHY4WxZBV+cU+Vb4//w3GwrSJQp3rbc5AHcJC5DtQU5f8Mhzw6zT9+HJ6
yJfZSu0jl6kapy3Ay3NZO8m2sTmnVIcCFruZgAnsd+Ri53ue1mt7/qAsOmcdSFr7y+yhx+dnBGlZ
SyT0sMUQiXMJ1HzZZTIgdTIYZqyoqB34eFRb3eg80sIjdtbxkXR94wF6ueQGCkEZnYA4SuurID55
ljcq4AfrCoqx76dxm5/NCwuVAEZ4jZpA0RRXOc0SaGn9iKaklXGTJwoF4ozhLOzYBZBcotg5uHWQ
GM1bfZwWlpkeuhsD9UGLlN7qmKpBZ73/uMNBEPGdFZfpwt4PER68gzNRDvWEP+XbeJyMrg4bNf82
sFToYr0RtW5YdCqyx6y78xTC8h2jml7AXt9140Yvrf3Iei0Xz6+2WtqjN6nheDA2Gdc3WDrG91KK
WMthRENBYeh7/7dPSaEdyEsaew5uF9z4S78h0QyNmtHrVUn6CfY6u4Po2SWw7myHj/Z49B4dPlfK
C+HVEF06UqPFL7i51dpacFQF16OTGglcunWAavIm6Gq+yFvY0xlQOe29jNlkATw7mzZHxrUUt1Mo
Cj7vE5FH0gxiSn5mbM1EDgpqySFZa/dJ62a93iUG5M1688agVAede+fdNXQJUgLe1vEEVZF9N/9J
fPOzReRmSIgg/l0UC8xjXzke3NGOawEVf/LaadL3kAyKvSTXbFmrtts8lwhkDrr+4mO4h6pY6FFu
M5zQLuWwzE11PNn+7FwLq5fGljBwky/4ToCzu0DuI/KUMdJX6z0bEtBP1wP6xGid0ZGSKGQaAGAA
qoxDspCSe6sgm9J08AQyv8y3b281DoN9vz4uLULExORcrtksT97vxERyUIBVRRpoC6WD40j9DaI9
ybOmlJZNH9zj5xrCGvMQAyAWHjaFGXkTxe+9NkDZ0hir3GvsqmZCRo6HNRxPJHLdy1G8yaA8rua1
wWw27TJp5Nos5l8bq8PJdHwE/uCa7X8Rhz161Ms/QXw18NZQV4YOmuUh5phMRL4uIbwuD/ePVuY4
2+nmiJl1I4JwqdaJwYOTN1DfrL4UDYmd6S1O3dq8x0anxYdn/QNgXSGmj2B3BzifD1QuuG+qt9rM
VaTdK7m7PgoADUH3IEqhufhiKWODQXm/Y9CqIMRpa50QzzCZIrtXgw/E1ZygeFmDEN35l+65nR4C
QGFmghOFChr6x0c5yVfITmRQF2KeTzRiU3IuFk8WBk+GFMTubsbsfUx2wPidnt7kcJea0+LJZNnY
Zhtx8M6UmTpzQ3ilaKCuh7tcDYWxf6ejHVhPvUAMaX6/LfhhRXoylBgIxbbQhRsFSnEJ4fxhAYjh
WS01FjYeImOE356GmgCRbYrfnlt4FiX+nTYlZ8X0tOCV3AAxA4CGz6xHufmGQT89saYNUQhPZzFt
wV4JhHxfjFj4u5vQZSLwGlIU3l/5IqngbHr/h9qVCsZPa2m8LpCaZGYlJnmHGej+thP0l55XM04m
uD8YtB11Z/tPw3KlRx/uuURIxt0I84NOxF+KAT916i7ElMY9HLt5eF00dF6L1pA3xW4JZ5b18t1U
0uSAX92d87cR0LbOFm3DpjJuQZaRwZOzTvU4ZOF+mw8ZBq+YKQJ9+yAqPN6W3Wn2lIRLxqODwlwJ
noXqQfqYfg7UcWENLn+AmCI0Qp4pDSTNVGEtWXGbYainMzAT8WVTyI6s6KU8dSFgMVvkDRDpSkDl
EzKZZdMz6kFDT18jaifotU5CNSb5P5D7hXk7x1E9ZUUTWgZ5ICfBgd3AlF4kNCaQxEYuWJ3XNsob
dQIW8TU9crS/RvsSDG0MGKRy6PSsfjyOYKnxg96BlGZP0igI/Jcwk/+UWckHdP8LkHUrQwrmIpO6
q6c2Qybgccz0kWnKIRoG+iglqv0cat3G4wG7QMYuEhvk3chjMrwWbAxsmrs5LxA5jbIObmczvxf4
v000MPoh5zfZiAzDXap7f47GIPg/0eoii4KW1n/uVED1EvUqd00X9MuasVg9vBI032kTdrmI3gBl
BjpaMWPDJHXrPVlf8RcSXkpmLRGNqfnDRToZxSO9EgZbukmDnobdWJgXMOOB7xPCD8SUminx7XFU
AKC1E/nXL3qiyfEq7jYsxCv5AXUkuJXcJRMxx1sTBIWmvDNKfNBcjhjUqLdhW9723z0tFIW1gt+Z
pJ3heWQeB93nTDQST/O1JTw2AZMowwiMF6qRhqhOhfyv3vaGDJyJetfYUjBU1ZXuIENr2MMiXyIq
FrQM98e4EhfbT6h5AaQLrVOqF8JlkiAr454+Om1vub7Tv+NwKRE2pYeALWve940lI0OItmSuUs3y
nSQvp+YTAXcb0BqSWtQPIeEfqH8qeV9qLpq7KGDZFT37HnJmP462JTsBXmm1kUB7N3lc6tMgp64u
sw2RiEGUEcL4knhffVSUWAMFflg99MuaztnB1U327T7FsgW3ck0Xo6R3hNBiFsVFqgOnHBgY877o
PM1W4C7vkufRs+7zLWjGbPumNT8z/3Fyi7BzVhlGf91D8AN0K8lWxJGZTOCzfH3V6/fcPdlNAvnv
QkGDuM9IL8lqMDq+Zi0D7lKqIaX01IXmoWLz5GjpvYoAz6vCKcZNY9lF8heYYb0TTz+4cXgroxoi
GSVVXGevwQEvrolaLj7BmsrCDzely+Tq3frvGgA60lbsqfCPgum0SXp1C1q9uJnOevyGSmSnN7u5
ogoK/7JfdIGO8J0RMFelQz92/NsoflMvCaTYWCeLpEA5R7KBMqs5AhQg4TySYxRCZFCLdnMATrNV
kftEg+dq3z4ylx54153S12SJsjgESwNDGGCJ5PkcVn1wZsOyjFJrJfLsiqHcWtngrYaTDJI2x3CN
tFxm9BVENANPxGSVw0X4PY6NCaCnUqE9HR5WISBUWllv8mtWUfbq5WSgqafuKnu+hSw//x0TIHHq
5HMuqc7SN+BSsOSsD5E/GxPow3jQdSEsi+QNMg/bIQRMbWvs36QfuRExBqDuqHiExXAJengEKE4w
37npK+7k69LpmC0wlPgJ9bc28/9S2AZ0Crd8GHjfDEn81rbId/ZRZBFgqX0j8w7Nb7j6br1qW/jd
U2WPXTlETy/Lk9V8byQKXM1kaBTEo7KGnLhHJS6ur+iixamIYfk6PEfHuT8sn1Mos903JDnGWIUN
6vsdl4nVr8maD+oYtXCYyDJ9vrivLTv1aKbOMSbJ+ozkqgknI22fM/0l0AcVBnOAXhh8X6CAp7bB
WORzmtgkB3nyMGiKXzdh0hFyi6wUVcpavVvRS8x3j9Kj1Ov2ZPAHhl23Fju4I7ra5WHIFC4BIlVX
D6hiAm8vEaHEJNkWaxL4DUAzhFU2n3UNRBu2FZ4zQ1HI8uT54J8/c3jIHxY6lr2md7nNJJJ4icm/
+yWyvibYLEz2qMLC7VTsjA8HwFrL5DcYK8m0PGrpk760YBrA9QY4vqFajwQ+BHdXrXroUcIihrYq
hXQ/DHkZTS63ROS9qdYDd08MvDMAUY1iAOb1/cJmD8Eyo3HdWPSqnEPmE/QnYZk3ntIePCkvDeap
FdxxVrmxGhD+uwYDC8P2b83/QtOLRpI214QFJL2ctq2nTZPuH+cr4l5Z52AQjtUblktvwx5mrgPB
jsVdBjApy/IJbhleEg5c1xVw4fWTO6Fw+V8P5MhU+fxGeexwJgLchUrK5kpDw6YDw5hM/nG42xtR
BiSCL/lzjguRp2/fDdpfYs9IlxxW9ioKx0El7cjxYK33Ay/PspJSZqJlydmUrC91+pWolUr4hYeu
8sbtqT2gRf0LU7WXtSrQuUErb3Z57QI8+MqH54/AB+srCNoRfd6LnTZBL4N7NtKmG5gnOeSdSXlj
XmpwmDk7IB9ZYhiv+DF09TIt3WyBGfQ3WKwoNH6cuhC5g/j3E0KZdaPucwjzZ7FroJ0WvzIhKGm0
iStKfGsMOTRaHloMiLZAAODGRSmJ1gjnOape1zRfMys4TzNodPHS6W9PI1vUOteldtbbeEF7sUM0
laqsasTqpZNqivCi0kCjHP4qIpdMEiJ+1jbTVHKpYLntaBTCPB0M/c1dUFz7LIxRdZRtQVUjvL22
xteuNFe4IdbLuNDIN67B6pBWFCuJL8OA4IsuXPl2EzyVA1TYEHaKgNvHIMTk/XqsOyycaub90dMz
7j/qiETwdpibyCphBb4ATreM32buyM4y6Zegn/vKQAZQ61/DcFH6VosJOOuCq2H1rCjPi3fzthdx
0eANUgVYU+dNVOpy2gTBirP1wdBM0AVlabYCRhvj/g/GkqkB1oFnXfP9Zq12BoIViRSOxYtRuEHx
b9FSeFzdCzQc84NIZ0oGJE88fcAehVG9V7Gy6vcrUrtuEZrXwzoHxRavsRkNKuICNPbnQj8QnQNq
erjTMfUAQr+OV/bn5rhMy97hDVDdtt7IkmficfB5c6Zge8aB+YiG1Ac6X3YM8R8OAk6TzWlhTLfe
7tpT348X27jnN7Ly2G1RwZWGgeHpXzvyTtgngO2+79KHq08PvJHSzb06KEhK5WfWWwbHQglBepRv
s4cU8rhmxJtXBL+YDYDb9few17e9zyPjOKnXna28CaubicKndRqgYzIfDEEsVMHsb+iiGNaRb3+R
fqq5wH+giy936bGADSq8wDqHLZeOPOJPqCyBTzb2EHvHl2CghcVE4B7Ur1ogtCrSEAxoGC/jX4Of
E9TsFfNrUmqGELfRnZrCLIOR+LkHLbHIaQY3jiEx1hz7dWSObR3ovVnREnpik0m2VQI/zf4PFJZn
YAdH0WU2YB1eyHmcd4/PkrlzLlJsudj3cKJ22dlBn+yoPbpSHjUJv2yLgKxTOr44iFat9m6uS9kx
mtSGz0RpkdkkXistL0AZZrL4zREWxnrF+/ZwRLuvJkwFLmBh3E1cx1xxSwtb4Jkm3iU02+e+wZbk
dLaD7//VYkzKwWTxfQpcoxH0vFos8zX5RrrDRZjx/xTGlvMCcMf06zlouiI719GSBavizyrwckUw
JQ5zFgJSHWjwA5cFLvGPPcYdnmJZmlEnx9oOUdouF8p0fgDlArDR3eE/kuCXibabeNIb0e9Shlg/
/kKO6eyNshNRT8zmYST5IsdmbMl03HMU77XhA1AqVKhaZ2iT9fnL+ylmGuZT6twxCn2NJ+akk97u
hfJ/hENeulDUfacuirUHdzT7fjygcyNQ4XQYc/9JaiFIPYJtwuKxjWxUx9lH7/9cE5zDC1jRLE7W
nFy/GWyJrWFa9b1/OLWtoo6eDxrSJ9LPKhOUNENsY6Ki82yEqmTtc+PLjtSgOt74fJGMAeoOOKsj
ICNJhVx7E4GjbNoTHb4XeVOX5o+NZmQWczZi7+YjCkIoc7gQ/x8qSo5RzSnWK6XrRQHF0h1FkHF4
meardBu+wH+LRWCMiNmqzA2yYJbq+odPi0DTFsf4o9bImucFjKWq9bcjmy/QzKcXchMRCoD3DT+U
fkeu8WeVYBoTdc02wwfIl/qNS3mY48wcziSs/Tsw/xo4I8sHWJJrF0YYUGwrdDj+linT6h6Vln1C
UIlPlrbMkmCh9v/VZ5Q70jMkJLfacI4+qP7QNMNU1M+7iSWbk3YM1P6M4eHrzYSfAVngaamIIqdq
/KHeErrrteoyJ1+89E36FLkMTx4j1C3gsNyGg4IOnfAHQjoWmTmM7f+msZp6OT6s2nXW2qC9Pr4n
+g0WYtLB5/LlkevDFiqvzBHCbAVVxohuV3hh8RA03PxdE3x+o1NHMiND+eDoUegXhQwlhHuSWkUN
WdMW9++6F2IFH4dxviHpr7zHfd8pJAUd5X1q0uWpAJx4a2jcDD8LCxnUIEdx/2fDO/OABkVXAeyV
sjHcSU1zZF/kALcTK5SoWnhW1GBZhh/Aaq9YwmlLIgPamcRzNphC9Oan7QumEsGi/TRe06hz1zX/
aOyTJ74ggtc2RqEvah+Qx6V5OjwYcryDmw96W6TYDBG/2Mk8EPIs37mA7V7vEDzMf2UFExjPM6j2
a068B0Ex8F3ypH2PSePMVR2qTKeUcy1GrZ6yy9p8M42NAH+tB5YYCNwI23A7HJcjin9whSyeDZWd
ZH2hH2FSnWdZnhUO0GxtHnH0e16p13vJ6+axItSlsxN5aSN0lV4VziOr+1pWzh9NyIFudlEnhumE
/uO9/yizOqK36FZyYYzYzl6EzKs/XjDjcHpzKETr8gW+K56c9ivzo6eqqPNV8zcjFuUoKf1N1zFU
RV0WtnFs3fuAZhy2NSKXzJKUjOhsFxtixrxB16cHzaaHoqEIhTFm0E/bQnl9udl8I/DtiMOZqLs/
91S6WjGNf6hY+3FvjSJN/0pBO93g6u7WL3dliS8g7VU0yvoOgLOepi1B9QyNuPbZxMC1FLaJWuu1
HkukTmxx2+rTh+SoUk6bndvgZ2PdxYdhv7QamVUPXlMm7EAkn8y2v3K6dK3b3fgGAQ6k6JtYemUt
N99NVu0500XGSuyi8h0/e6op5kJ6wjwyufh462bRdVsWum7E1mdNhK6FnBcbvvLIyiK2w4VQ/LeS
Ka53cA/Oh7QMAKaWZmWOn8aVExSOf/3HTw+1RDbwT+P0kOa5Bw1/2UTNH43SEh1ixxQoJBN/WTfV
i8dLu55UhOLuYB4tl+yiH4myZc1jGJUGBPZP1kUc2novoIC1d4NugblMBmEo4F4H+5YgBfB99JG/
o2Hh3bz9legnb4xk+QU3nH+Lx0g+fsqsgjU6x1d0KtxWTbvQXHOH0aYgMElKpEoNR+cz8Ta64qhj
/Qpxty4MzjTJssbRErf4no26D0e3aXgc1Bgh4Gt8G9VzbhJpo8JaSYikfcVf2n7nnSMbo8w/5ILr
7af5IPz/opNLGyXJO7dwqyr7m485llXd2ShrKL2Y89r3gl5mMMqnS2dwNJzaFR7IfFMhiyqyTjoq
VGE0wPX56DJyCXL856eQdhCHk+TLVuOq5kKIFT9vxhWW6N/NdLYloLbJKv9TdMuRMxktsYLjSGDM
OJJhcq6nQsqq+epfq86u+MfXsUY03lQMo2PdIWhxHYDr8LTvdfDBVaSyQBCbmrgboFvJFW4PCY/L
JpXicjI9dE19cQ3w4LhhBhuD68AXFyaYm92C4I+GIkblmBVy/Hm54224FycRvB+kyAoc9Zw1GUVU
/kzOE94gzSMD6MYVbHjIoUTmnPVicNtNVVQf2CEKF25Fy9hePuqxV997uz0bbXP4d7L/uVh/nStc
Fh1tsXT4j7I1XsD1hiqB05alXeFNPXjMOSm0SOhWqOjdjL48FjPaFJePvOEDlYIB6nUrRtUikUlJ
zF226qs6w7lD2NnL5jadhbWWkguCF5dU1jkqxyWEzozjYoqHgoXaY1V8lefNLqNkwEZyQqw55Bxx
61oKyd4WE/wLPrzZyvR2tq77FGMh0Z9FoQvoybfcJMTi+XHkDJPHpBfpJ/qD3+ArVMImROrd7xtX
KU44px9uMaYJ3KFMf4aKl07M/Ar1o4TRiT6n+44vj+oje1ksgQiMSKXVZdZuavgc/M0vEzwrWc27
vg3HHtp7F7ZBASKx9iz0AvAo2YK2SaeNuVMWnSaezdcHmri4Mwu3C77B4+dB4xayAUl0YYstYDVS
mH5T2o5tnWG1rjX98ZAaxyWBuwQsHddKPT9Xvt9CqD6qTTG+zWdi5ftLEIAZjnJmeiSb3Sn8c6Oj
h8r6RNs2H89yP3AcmtR2mHIhAJIwRv538MSeELnEjIfHYdXsJiTZF8k+gWPhriSq0tY7FYf2EVYj
PGOTEln/7XtSs2lpgEsC+SVVL3xzXW5H0thDJiegKfDp+7YJxNR+oyCaELwuITUc15rLrgd8T2ES
OpdSr1pSV4brg0qJDhbPa/osnPw++XHzC+A/DDk5lSU2mDqO6ZwkPTtEcu3Fxq4F6HI8mfZIle/6
eEQO2E26hqAFT6G0I1vKclQJ99B2TaeU6G+z41CLLa//fHiNkO2GaxYWvOsOjeTVzlZVtUlAvVF7
tGo6nqdpFyqWDbGmlDg1DBxCItHhTyIUn2Kz10tRImUKgDVrDJDgY1W38t3KK1Ma+6J81EyjG9UP
tQ2s5QCkWk+ge/7cDczIT9EhAm3njnfvqg5YqbadaPHFS5T+rczR2T737/0lb+5d9P2F8VMmng26
XErZiygYTiG0vRwZDcZdmONvY/f1/pDLYaYleLclKkEb6cGY27lZaYzzbFbaH5gEIsAC7XJYGhzK
mOZWjPMyyYI94zukj7oI/JI1zg9ftpWlSnhILdiRYMXSyIkPsK8JJiWsWsHllSRnW6eVUoDTA1GJ
g18gmJudzIg5S4PbnhBO4Jp0BBYc/L0hdg6IuzIUbAiSfZvh9QLEVayRgqUNcWbFvTKucL/jqQou
pMneTIcI3PjgbS9xllZ6I0Tsc0H6F6DOw5getvhHdvNjbYBrwPMLzz5yh2TBA07LQg/QS9AoJwCC
TeJtI1cQjcG5bkK4pBwcJ0qj2DtVpTKOkTrrYpl9nBSNdBG7VgKY3A7SR5PGTLk/ShSDrKBU8yfm
Oh1C6vx4GIENvlng1o2bnaEq4BM3dO12rfaYUiFppfK4tADW6A74C5bNfbdBU3vqe3NKAOGi6ujV
GIj/x45PRulzQdTTF9UfxB249rzEX1EG2DaYE9G8tkub3DHU4eftxU5asXCKs2KDl/quPHxinLlF
uVuFRqQqvksaTu8bQnweEz06/1M9dn/qGoC91keax3N7YMOJdvsOQQqHAjKlrJ1szgye12ZNpyok
3hzYfYGCfWPrpD3ljXzsMYi46H/VkJCQauStBvwMihRhZG0aeOWec5VPwKHG0niAsHeoFYEJcmaj
vd6digh17NV/d3tNH1UUJ2JqbGyVy/6CCabYzbIqPA3X3eILu4/EzpKxwka63B2+U64xlO8LVHpt
EbCRnxnI+y8dWPvgxVw/z0V/Nkdq0HMH6q/2ScVkazTdbrTmIF1kpd2Q+F2GWenrM3Ih5feZoPqo
B0a2Nrt1XYqHCoMPxm8f1EX4CgPfvV5/ctYjxTlxFwZoiuNC2ptCt59p/AOwCyq+jqDgJxQdKrl9
PJdeLGALnAhDOE1MxTi6upE5V1nL+QkDeA8iY4LMUaoprLQaLtm7N7REebpuh0Fgrh30dmYw3CKG
3mqh9ajyv4QHcJO4WXYVvBDL+QjFl1oL9vu+CjAG4PFXO5hCbHeGoJ/+wCEzn8YDM1qjHH/5O3KM
y7GGleAnRDAMhQCZN/W/OBR1vu7I2caFIoyKcbV+ug==
`protect end_protected
