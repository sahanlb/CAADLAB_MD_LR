-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
CtZNX4qj5kTjLVTEHzTlShJuDu4rjNH0Z6qKvqPhKBO16C9fHDdoj+U15+5ze6ac
2SqHcGaZYvSRmfWB4Caty5JmY+cT5dHstkn3VAqvboHvCiXJPG8uSRjuhaYuy2e3
xj/aODYKYmsLjadDhNlFjZFuKmw3H2nkXrG51dUQBHk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9834)

`protect DATA_BLOCK
AeUL7XH6cHd0FRH35G9dxloV9BRWDMH6Tn82U2tPWIlux1QjPE+5OSxca/6Doow+
PLzGeqQKLlZHkhMTyUfdZkWkfbz+flPWm16dkclaa8nFO6/u2EVYnHqLfHtSl1fo
dBVCbGtrC7Wa0eDp3cGjc4pO+zaP51ErE0Jb/YPgQ6qUkIcMpWkzxKpR29FWpV0+
7aqfmjAn7nhokynu/GxdTtNEGIxX3rjo4pLeF3kqDv9gfZM3msUERkIvw7CuSpm5
1yOCZDuAIyDbJp5bvFk3x1p+IWLmkm7ARYS+y4oq4VCdllwyYfEqDALH+D1Dwqa7
waoUad81L4E78mv3TFAGkOQtUdkt3/vilhex7UUOaLPKQItY3zLcLEQtN8z/Q45n
5Db59FwSiV6zKDKzvPK9AzPQXWf43rUCM4uLPK9tXnbCWb0eqHDIcjHBfsbz6ivb
HcfB1w9oswlyaJ5Ai569qsVp5jbBTEaManWIokya5la+X4x8qFgkmiN1dPROeOWd
vqPOFLZZLpv45miuPaC42WKhJ4/PwKKUGJeHzr5oslk0dbZ7bsEn4RkIWn14bM5i
ppeHDwTSsoiP0zXkpKG5hpNBJP/YM6q1HDrYmnFRHg04nVD+q3+TTTCC0+FJ4kyE
NX9qPgjWKBebieBx0i+HLKeDM5URd6YFYXI6Q/Uxv26dqSgXqAZAFZ9b1WG0MYGV
Vwpec/vfi7KKhMEphsQZPJvXg0gaHuK6zyn4smKxKWOG00VtogMRVFyTYX58sGzl
9VeqJ24Z2/jFDRLjjxl/nUyIMm3qAxSJjhJ143u+RL1/XNdKZrm6KZVW3litpkgT
WZYHwhUb7GnYO0l38BoY01wBu0OIRwVchJZohgrxWpkRzM/o+4BJYqoFlU+pzY4t
8345JZoK6ZhaMvfrERyEx5jQswfNZmU5zd6hXmZJHYh5YjcqxmWrYTgmWjERz5Yd
t3i3NlRvnbdXurVNnJBdrPUNo6ctpSYZSfkCjj0576eqAuCyBb5YgO8SRL5z0nwL
Tm8aNT4JkL99+oSWg9sGTwgfPwKC/GvgVLmEynNT+HYl7qDOAmOmKjyB0gmGllVh
geUu27UAL/LQHYRJ6Wx/e5ietSyUQ71ZpB95JhDj+t7fct5Faz96inXww9VKRWoR
8Ml/RrQZoL+EHMesVRwsbs+kDThQ5ZmoAkySnRYOVCM74vQI83Hj1sp7ixWKNnSN
Kt+AOScnw5/RVASnGnCimLKOeNNq+Kfy0rv01k0zk7Iueio6O0M1Ti0fj6hkKaih
RfgbCycmOey9cVXnf9mAuY7b2DtM/XiMq5Zavp58dteR7p8t/nouqMhj1Ztfj/U5
WFc1dOjcdvGDf0BGA+UTEIxcYBS9TRWVvrq8ezwmfXWPv+kvsMjARxA3J00Of9K1
VC0VTOUBDnxA7nSRrHlbq31vSR0fSBZVM5uWo4oGuR7uDB08/uO94GXb8xKglyxL
SgGltWJGyWCVFlA559arE+XYZyW1Gan4ZTKReAlMVHhvK8GxMNsamAiutMt1QpI1
OkkuR+r1j2JCU7xhuniEPA3F8NKM6KUKqzWeuzFGp4lob33P/XBcVC6eAWYFYsE2
nk8V9nRyAOj2vMD8LnhiFr9s1tpwxHlyoWvf0wWRrSRcc7Yxqp+N/zL+6gDVgZOW
GxX8y7AKQxxgzP1Jpag1iQK7IE2vMr/MBOBqye40HaGCLjnsfctTDBoDGXNr+/se
xb3zHdGhF+Vw++fL1Qzjm57N3SXM5QDY4NsPUmsqhJqUpw2gAui7BbPAA/l1KBjN
S6eBxA8W6jHb7dKCOMpei/IJcHhRtlsyd2hq02vFEZpdExOcHR7m5yaqw90cp/pY
l7T0Ls1lJS8nDWlio0MsU+8JQkCgP3rf3x++uo4y6yUIF3ECOOhKuxiMHAa1tcWJ
l/8oTzIT2WReBfg0TAXe6afbmP0NHYjDDUBz0lhFJ4LuwTKknfwI3hgw+oKZ+tEx
KNskQ9iF8cF8iWM1ffPyt8MCPH+sVjozwyC5q8vqBU+Ypy7zl+Y3phWvbV8jlRJ3
UxOS//EA+Sn6i1Xgf6BphmdoslbjVAiZK0HtySdAVVUVAcFeTQuamb+a3YtBR8D6
nf7VsXngczhrfL8dWEZxIPxabEXgV+JrPUSiq8RRgVCD2c1WwkkXaHsPSd9ygnhT
YHGgzzITTtHZ87TXMA3NyAktdee07PfHGa43DDm0h3/3/zVA1DfdsDEZwiIXBzuR
dNrWY83nII029dQxa/SM/4z/VxLBxvGxUl1yLwUrTdPxmyo6x8AHH59LhVgv18Dj
ED0HCbdH76gviwkwSWF2dFpcKJ9MdRLNpqnTZZpomQrEmapMHlAf95v6Wo0TGcgN
CmzPF0GcOndONUmMElrR7XbA/rOirCCPpboCMPv0vx3cSjzk9jmrhhh1dTHtqOUv
ORwqLF4tj2KEaThqd4nA/BBwilrFyzvqPLWu+iPbuGp1cScrf5H5lqyaIMhoO9/Z
0rCMr0/dvz/3n3EmChvKfe7KhzbN/4f0Hm+UPTIQT2s6FEvKGwbbzyUsyLGwqHoW
A8s3YZnoCX5mOwyJBR4i1S4oXqUzKzgfNYFz+1B5vuH284xM9uzWVGJ9AZwrcjam
KFQT2cVEWkoxvp3ULw8CF7H61PMnuW8PwT2rqBuJE8j1L/bTMCQ9EcQ2D2K+Z31L
yRPX0SRImjmWIe1epIUgQRyYUfyRw9V29+6rdymfVqxVI3UBzENfS5//H8bGfVoK
pJQO1aEwiF6ijYgNaQ3CqIvcxZLBsMm0PaiZKsAYdKPQro+7auBAL/ypciLni0bf
fm2diDdSfP0iw3R5X23dBs8apPWNeeTdY+Gl7JRS5M8XjEXFHgVXPxYwE7/pKFlt
3HZnv/6DbTID3NFVUAFJgiqyHNs84g782CGowjqN/rjboSaVJK+13LUmk5se51c3
rdW3k75LiQqRYVx0lF8g6I3U4Rli98tfdArSdbaOLywQ0PqsPD+j/Ati4ZoWnKRr
04RtASlpYe415wTOjaVD7bIC2Cc9URfRMGVfLqqLYgdz029MPTBs09RbbWNXW47E
JFDtEG21Y5uFX5WFtvXqeXdt8VBvkwJYDDd4Y4qSDHDUQUoDnMXmC1AiClXWUdrH
wvVHK9gZKyBq6uLeFugSNsSVs4gH0jEJeA3ql4SU8v9t4l+9UrJow5+GD6AJtVSe
wM7IHKq6EXj62b9V48CvNtyWW2mOugaBTydKjZLXkLE0E5Nw7ZB1x/l8B7qRjTUe
Wv6P6YclfViEnivYzYR0NcS3+MjV0cC/39fRbgbKP3wkDuSX29a+r7p9XWfWtJDv
R7bFCBaUsPXsjSYZ0P+4YHS1Bp8ORqnjNigZncxp1dL/SSg+x906qZBJ0R6UMvhM
hKAUdXRdo5LwrWKhMjkc11WNky/hbdkpTDEPKHbs8ZSv/n8JOLjZX8X/TgF9YM8w
qnGnNFJub803S2WNLb8XBNqa0aPROCr+j3QvHthz+NUmNOYSowtAre0V09cMF7HO
ThFbsHIHsPCQyzdynCzXzsSAkfzdswlQ9GSjZfvP0E6n7lC3SRYO5XmjQE7ZVAe9
wQfp4JrgnYF7gW2GtMi/ktc6Zy1l+D3tRw1m2DG5R6w4Bql8R3r3cyXx1znc36it
6gizhu+/Xca7olNtFuDwai9IJH2UdT3aKS9/825WlQz7LG+EKQVSLhk3CknuNHHl
e/SqMjtgjBJqOxh9Zo7OtdIbHx5LT6fsNJ9hR/OlIDEGYejxyeMqSOzW2gpIVVXF
Pj8dmrkG5LwNSaRhcm876ebbj3yCxEj9Dsj3bw+kXaW0y+L7AoBRZ9JCCRGF5Ay3
jfCpye+4CagT5VCxGgrImzFIoLreRdPGbQApJlu2aYlZtV4wmpvrMz3MDwcw0y3U
7WfDoPqCcSNfnvPSZBgt75VVvwsE4Y3sIl60dNpLoSekAx3gkYxkI8sJvOpEnqX2
yBV/vt0kG/aaFNuRFzQJhKx2vDuvwZfz0lCN63Wu4BSPP7EjCft+CqYVI623W80x
mzj4cY304+MovcB0Hlku0y3WZRBywGMZu9KxCLZRYBD5eS2+TeQPIEPFYTO/58Eu
Fe3vMxhuhl18rhIo4Rne1hpeJeLWgQ+UQ8ZnUwO+SVVIaI6vDyl/8nR8CWp+DjiM
AN2GeNoJ3SsQaJ8I4xtgvPaKViuw5xnB5aan4OR8Ll6hVG9ysbwwoYIxtguFLlew
Y+er7lCnpt/Qf2+Oge8/7b8Z0lCR7/gyGa+QV8WmbZE7Oag//zWug63/qch93Udu
AC8ZyoHf/9DFiR4GRGffwll3W0i1CElx6QxlPMDEmRCerVohlFbMJpmd2+8xlvWn
eu5Ld0FV+BnKd6hvvadHXNmUFXKNUGDq6myBbXP/a0InKcgQACwXkUqRthikWViW
Y8LITLip47CtxtiQUGhcAfQzQXoDQ8JkNYWDQpaAnuRMZy7BKMQBZHQdKfzoxEmq
r8ipMGtOM79a2GHLZ1kgakDnp/9ahS+wbw9rd/9REWq1q/1lkwjNM5VMzeft72sB
7j4F0mew/gGHk/BrQqfARGBQdIVHxa1tcDS04lbdvh6UNyeMW+koG3KcAN+FaYrt
pK1cccH/7zG9iYdOPUZ6PypRwY3xirF6iXEEyr9vQqaxP8tfCipriWs9XlMLyl1+
8Eu/XZaJRzV4bUYn8uPqsILChIM4+TUWuHH2EjvcAdQKumIajGmGk2yu2KWF9RQK
oxMuOE4HRg9Kj6rjzRtqfhxXiu1T9Ermdy7lbyMFUe1viJIEeWMe4dicqLYpa7fl
MAywhZVqlOsle/4YoqJkOC+7PpnUZKQ0VVv+/uA3qlJ/UAtpg+ljIkhcbr97oTj6
WjH4tU4S2bbE5oybGq54P0HXLO80994bQ4Ux3TvCz++c7EA/GNmxt5SQYO2pi8nJ
5e+jtpL3kSMDfvFwkgUcYIZioPJvlhjELby7sqLa9ZX4ffzfUed2fKcfaVzh9A77
raE2tweMwIt8Z9odu1aePvfDshtX5BinZbC4i5Hm2snGS1YVdg/KekAbLcJkJEdT
zmYr9/kHNFf4x4W60pyaBh5RIUepZKOQHL1Zb03kWfX/hOtqSYt7Gcaw8HnAIoyn
w5OUPGpf+pVZTWNCyDx6c6Hn2qAJqgTO2TvDN1bnBFSNBw9GOBpca1UXsbJwqUAo
8962ZlH/eJt5tJ3Y+cNv0f1KlDmyoVROTeUjx6Werxpvu/P27Jfr4o9BSihr7x76
/xz5jCU9RblnSjfqCCK9xiXpLoLh0rVJ3n+t4FNpN0UnoG3Xewu7o7/g8lXr14+u
6oj5Wj/xzFkzJZ7OFB0bBkpjF/xTXHk+FEG2nPiAsWAzvnsThj9RnGXyYhoihInG
YHYZNBanuXAT0yym/Irl26X6J7X6u0eCdT7XPmnwFEHYhzeJKPEdNU1mu8APWVdI
WflMNsLh9WiEbSYAfc6cQttaL36Rw5iyO6hAqR8O/efHyS4Y3tPIincuvLPzAZWu
dh4Z1EFCJvbVbYiH3c1cY39XHPaSvXJtnYk0h5keVxNoPUCX5V5sUBz+Ol0iFNtd
GmrRgGLoq2ySijNF0lJlV/yHUljtzYbm6rZST9lcNBNKyw4bEouj3hvAjnHFZare
vsutuUOKgRkVS+hcQIaSI3izxYNjGIl4QApYteI/hVmt3P09ZXo3iKm0cXHrMRA2
kqVNCN9H8p+8qtfzxsIavt60JAJItCzHFlPcv+70m9iSZnMBS6JOkTlY/ZnUUZ6f
Q8Uu57W+BIUqS4eP11JjiiGRFrMCvsi5KnqZSjSev/LBZ9A0F5PA3MeDyQI3Hge8
7iecSRU4SmiutySIw6lIXGCdQU1x0xFz2QpFE0gWl5gJfB+lzfomoPyOgKyrugUc
1qwowXo+UxQeLUv3B7y88IwPvQfGVMRzuoIAztb3U3jUgJWQshcWVmCqlqIyRsWF
zdPE3WkcDS1zKeFSPKg+Gc80+XIKTLlaFKbVM/t572jKgQjlgnFeVe7kysqMYZBg
LNJ8QkqxUkPx/Kb4D2MjdHURO5N5hp6ErGnKjGO5D/AqFf2rimkO7BoQeKs1iQBe
d7Dcn5hzoRKGpXXhLkhBdmb3XWMpYztjk7L/DhlNho9qr0H3Bkj2jcr5dN5s494Z
m6QMorXovJFdvNLg8A581DIfbhWwHxbiwNM0GpDrAvr6htn8jzUdA3AFY8V1l2Rh
HJ+i6X+hgt0FQywoMY7I25QcRphI7yITW0FYqhzYy8I9i8J+nv1AnpjHE2DlKmLL
bllAFXduRa5OPYirr6jwjYIFJ5I7HhlU4hEfl8h4QQOOFhu4yBGtsu90jtf6UB9h
gGGEVTR1MZKbGh7oS37IuQqnCIaLIKH8yIC+AY50gStK3ih7nzDr2/HitdqRie+t
WE2+5bvmPSfCWqr/eSk92/d0QnjtVHKKlYOyvTET+7sIqrmORJwfdg1VcR1bU/xH
hjp9A67PSYTpVI4QHRl++luExJQCkPu8hTK8fTrMPtIB2j5v3tSfwHzdKDxUDGRn
hLaFEBXD955yvbS2496DVmlpA6+AaCbCJohHAu9xKat2exmIE6I+eOfu2c4TZ26g
SexZlJHIw/sCfENpIWOwFccZDCky3AefebZi1rho/yLE3BW/kGYZYF63f56DQMuK
4dvfDnHRiZB/rHOs87R2r9iXSpUtIrLI5rdl15uigrO7FnYMNyF7qaS8bZg8Ijse
FLE98QfHJYWi42c1yeNygVIze58OauDXyG1Iv6yHHl4j/7eyLDSvWkW1mTIlfaGL
qElJluLRIcmRTMg3tBukhYdNu3UkhERf7zn9g3c4DtVjZb8txZc+R1VP+p7CjAlN
Qbpg9HdhyzpLi1AxpNJufzT1sjEamYh1KDrG7hk+u2wuxhWXqdFfeh5JxJzyN7OZ
Lx3oil9eu4EgOAMIbijBtLPQoNLVDkZiVlHx5erOlKS7QYBJg2nsG7V+M2Ktzrn6
DTYRHkva3283DJXsZ+0NFVD3zWtbaB2TIRKYZDZejb5FFh7la3xn4NJv8ok1zgoY
dkxihRq7wHA0zG5fH5du203Kze+sKh95JvW0zZ34ks+Durh8WMMtiHoVe59cF7CH
acdnMqDV9lSOrg/0v8zz6imZoCBu5cSiPptMfGt6VL9GrGzERZma7/0tfCTHKMOp
A2CNoogxvTclnOJ1+E0z0EtVYUTftnRGiZGJzXdmlHCWkVyb1TTTSRLrX2Ouytdq
LhVWePMSoShjm/E2KmWMBdPqrTbdJ0gWIJ1GrQa29jdV6hPAAXfnn8Z+iG9j3rVq
VagujvqeEEA6pYJXtM6tsUnWnK9nEv0edUeISTjiBVSkYqHvrjCGhnyjNdTHygle
AeTejZQD8uMad7tRgdJmUTw31vVgG3IRgBfZkgyNbrAnB1WUYENwKzvtA8exb7gH
6qETJhjtWmlbvgTIb1aw57ois0f5qwMgP/vYGWCm/+yIajm3qesm+EQfO6MnPP3Y
VQm5w+xXrO6Y7erWTvyXhoJfIOfWA03W7Vn2PR9B5XyjXPSznnCgyP4ilRN7ajoh
mL05R3Sj/8KQV7vmLeL4PVCdE4ERIJbWCCU7Xz0Gbi+daaectvFjNfySbpJR5vCs
LusEOKnscAJj7gCKB6egasHhIbX1/wQF3x1VMUfxR713rGd8+ag9k6O0onIs5X4M
5WXL8ssW3bBw7buWuL+dFT9pc/r5bfpUcUrrz8Tv7Vp8zKhtmih868YklS9qSLbP
fiBhiTAk6QStlQrDSa5lZuG6okIWboI5mM8amms0BMC0EzZ1QiD+aUkd+aOz6I5h
InWUK9jgSa19ERi3F1bTqZwKm5elz4lbAtZVCFG2Fw3Zp53bGG3c9KwdiJtNfw0L
g1kzAqDaA4MgJC8t/wWFGXerpwWHbqSLCpU7zYvmzAufkQ/0h3ttFWcExf6cFRMw
iBAMbabKPmn9C4URhYjE7TcKf88ppwHZC0URwDXw6b5Vtd7xHp85bLqohG8cmbBC
kAFGW/VI8mlFTsWenjTgHpA6jpAF0uH6ZpZ+GEU1GDb5H9WuvZ+0PQIjEzQyzpgc
fNux0aYgBAPUW+pPMxCDE0dUtgC0fXnyvQZshgKPJwo1a+9KhSo/BWwEIUDkJppQ
l5oPV2K7Vgtv6jb+awUT074SoUqKK6AVgniPakXENfDmNU/7rZ/teT1nUn7L649i
xgfa8i4onnpzXmf2ZNQ1+eTgAl/sFzGQ/l6O8ZAqqafiBKQ+5Wk/+xFewFkYa/z2
Jzeu91TzoJkPGzYZ5RSZAcSged26+1s55wsLExqL14s3TXsGFC1+r9Jfk95wra0e
pnX6KsnTYdNPYDmjj7jT65usdm+pwAkQV3udzJQHVCBhuRemrvS/zwBlF9gaOS9e
Y+z/YpUJUq3W+/D3N3/RXNnpwqxt1uYKVA/G0zOCDUaALJ0wdOZZq7An2CqHLYRZ
U8aRIll9tin9vyebb7nUSm0r+XF31cZKl98MSYHk5VstUeZO1Djl/RtwRdcYrLbZ
s2Zxw3whJji5JOT41OI56AD8/4B+Jc3yrlIYR1jNgFgCrWuTzzTmFfsKE0q31QLo
X58n9F+he1Mvu+V7pfqO5kTAKOft21DBzLz9Tr4G0N6OmpcNq1KTillBxu8TOmKE
iw1Vu3ueo7YJycbZTIVoOOzP9aBacP/uziU2VhhhlBuJZVBTqwh+qBECRTX0VvYL
+3eY59Go6nsHFqsY2aDqKBD2EHp59QkkvJChM0JckkE2yeEivKkuxuvTSsNWaeJu
EcH+7lkWq0IsIQ5gw031TwXJoclBdo2INyO811+Y8EmBFSl/HxSSf0LofGpbclLl
sEQwwqhUG9imxhGgXbiU6IkIzJc3psFSGSTogE2p4xM7ykwnaEwGIqYhVMKQSbQ3
2uDczR+4bJmjxndPApn9Q9dElDG/xU7znzRKKAcDdquPzADJxIp6D9p5/59GTAtP
HTfdqP5GKZHz/cgxEizvjslRtMW9ZMxnjpDCZAUdoPT0EzPvpiSVFR1Ncnc3gnWJ
wGGoKJDpopwCR5rSigIHTkqTbFN1dVj8D9mtAbGbpTzJnQiuPiNLenlb7qw+1BmF
oWIoF2h/pUHG9zgl7aclMt9+MVP+jv4Dl601kecGkP8LwrcyLsUa5f7wZCV+O/rV
3qz9ITgFedXNjHhxnc5J/Ft9lWB6U2Tab5xQL7rgtH2+nkfPQsRxgWCwUZq3P3/P
9RvNDeUfAaD4ew3hKe5jjmfzxtlhM9AScK566cWcqwaMzi9M198bLTUooFnMDrYF
6plCZv0dBAyM6tdpilNpqseSiWhBa4WVEp4XM4nKS/hByABEIcebHWLNGCNVcT0g
dr3hir/aHFaJleph9OgsXL+p9XRmhqaPTahYr9WGLXCBzPmz5BuKEW1kywA2kfvg
v31dKg9G3UMjpr/GdsoDKsupLzgxTLbdk5ix48y15J7N23I/5NRqjiJ5VacSIibf
gnj6mncrq5c27d4nliMcu6dkZAYslJWV/dwXyZ9qkzrv7rBu1fEGJOtOvmDZ9Qtf
QjC6jBf+mG0EEx1Ak3eeA4zM1dAZTWwkSNf3Gq/8qV4T0uRdvilTZhNjyhzgIUFg
M8Z81HXb+CPZN8s+JpPtxQ8nHL4s8Y7A8vEhGpuw5rWhEvYxdRoPXymUejM4v/MU
MgxZ5IkoyVTmm7jRTvmfARqQKyznl7cKjU4MzykLhjVhCW3KeXURhH3HPHcQZGkt
2Rq0ouwXhfVsr380Nb6xbRLaqxb/8mo6+nzbFgPKYPtkDwBZFbk6Qf42bmIbElmC
kzmYJM48w0leoyNnkvKuJjod0UTdrhego7jE0PjvLwAraZ06H4djrJg5MkFQw3qo
62/HLXp+ephMVCTenEQBvxUkDj2bCzyhCStTu4Hv1jjfjNWUWzKLm4SnaBxiB+Ge
W0JBOuGxRnPL4UXWqQJGIeOXXZt0lAetmHham6KxdWjOfktYP2e2psENt2RteTLG
up9vpPOICYrHPk0xij0yHC5d2hZDEWhInQv3BftYYC6kmPO8Twbk0DDFS8pKA2G/
rfMBP+YU9ybYDJkouC1lWc6uWahSgvSG/pNkk2kI6sRvwJ/gnc21yIomHCjpwHbx
AWgub0HmE/Uf7EFYZSOf57PpNETHXKrXQVRO5rNC9sqZZdyzN53YTZsmF5F1W0Qb
ILCLxpz+227JUxfkT+brDjgLsRMB1RXWnRsHaKxsWq8aK+KOmBamiEFhNN1JNAYf
TfF1DgogWbx2CZd+giILknMrqiXGvIjEckP6KoFP57qqg7uE6xKHppfOJ7WdplPt
WlPECV5eGzsEO2inIOqy8RzxnoGi0lIlyF0Jwqq2SWC6wt/90WDM8NGaHJFfAtOg
53cBik+ji65bWVtFbG/eoWyp5/TuXWp8aqbHXs4VQujUl2dqlrtWXsMO/DdeNjB3
YFOuKerrYnumlsw0lcixuoZj3BKPDU9JC8VO0rzPSSAX+7h14N3i89N7XuV0WJgR
Lb5DCku11TU6q9aDTa8TkTu1wQTS/+exrVHqUzORqbs18pZYIQBFi33uIU3i1Ic0
2AIag71n9EhiwQlm0eeRX64ZjmJF8zsrIpPM22FW0oBJumw9gT3J4A6w8pwMh7I4
TSl0JXS7GWR1SN6eL8y21qNmqTFt1Oi+OGOuU2G+TrJLKlKVfja1jJGjmSv3P7fq
KoqEhRGfdf7yeS0vMA4MpluPzXYBmyCJYOHFbCo0qRTZcZv5KYL/Ha1zA6MyLiK0
voMAazhlT3hc9DB1YoY/+JIU8JR9E5s7HI1yjJf/yKFBeDs7jkNDwoANVyGP191A
nKkAUZG7GZfV553XBht/N4NgMxE3WdyK+IgjvgRg36KHiX0A7MEvAoRWLf9J8kJM
BteWvCWCFplH9qocXNfRN241r1n4gyP8irwAKHpcDirjiWVh4p1TWLP+oREiyYCp
Cz4d74s1KQzl8jilsXCkwPMfxzTN1hreVkDTIIE7gpR3x5tqdzMHg6rsEHBVYf/x
96GqmB2otVHR8EthuFhFiDcv4s9hN3N6+zrLWhx4A04011dqtOSK+dQDiIxcXGJX
rE6EDpnT42hePxGV9Ji9+gJAEhGwVwZsAHuFsI2j8C+pAEqUgpA5AYB82AqCU5wC
bYE5aruh4NVwNzEO8noqKLa5g+vEF7cfqNAMZx2Tq/uq4y5MSceKaipBCClC3rf9
KVDCoIh1iYdA4IDgUSgWoX0ylfNoaxPO/Z7PW9llNPdWpl87/SFfk7HfeoyfUDTd
ExuPaUUniHT8FC7DnI4Azr8gTfagp4i9riLNcup7fR455255I4TadVvGV0P403yw
8VpborTMlVneRM3fjzq8LuMWu9yOwu0C8ZA/6gzj5gGZCQYUv4ZvChGSjdXfkwtb
VJ5VR0UbgFr7QtSWNwtOHmoeF5P04yPO001fbYuKkEhmfAa8UFpCHcO7KkvQqsAd
K3ekvswz2HT/H0dD3kNlngEaXI1xz+3dby00PmBy4cyPFyojvx7K24AWl1FgrN7f
qrkpgsdVwi5wvxQAAVlpQEM7pSjCMQgwV5UAdO2/UxOp9xyQgBWKAes0ihp3+y+l
yrjukMHZENQiBOoecN9fmPWUXcrZoFCcjYjmcE7jUCM6ukWiBQ4Ab0h8EAj51oZA
eN/czKpUvyJoFc/4F2thNa5fYT9XAdDMMVWXuPlrS54VhBTx/0kdEUU0chaFysgt
FCDgOi7QSms7HBBhciTmQUdL4KFtTKGKiMnjsjDZyMrEPNhy1UpA/F1GaK5CLv2E
yM2U/MCUVDPF/XL0iDBuQ89m2OvjhBeQPqub/5M88PdDeAibYCvkecK49lEzLqBT
mpoFp/3Y7M7pUDl9gJJWfOM/M67hj7rpyBOw4yOKV5+NFl18kQbb9mSDiTqpCdOf
2lP7py3YlSP5Gn1gjXMWneCoNS0RbJVCvgxQJbalzw9RTp0ue8gJJYnVrrgdKko0
DaOx2Pr7E6Q8BKylK4CFpHMhvQhjRcigiyGLkmtfvZXduQxIDUKUSu1pOuZ6lFZP
JXV4A8bkOPtUlQezLFe7GzvLrAswNRP42xOvIrKDi12tJT4WMtkI5UcwRKEisXXV
5Tuj63bGQP1p7mecbNnu8w8jD1n9M41iAV56PX3uqko4ymymfO5OwWQ2UeseVLz8
5RdYU7wgFPDkicEOHvFMJTOD0qo0/KPv2pR073H/EOTqKgV6k6rQcuVoUoEKojic
ChrfTkI9wE8skqHqmJOS9hrMHCZyj/zFS4HAZVLCX02wQ6zx6l1d3q+SdxBlU7UI
/bsyi0b5Gfkxup45jonuE8clLI2i5L2noPbQz1/28ShKfbsx4D11v+qQOCHl6lOG
xVGX/w0eub8aFJQaZUbLnuTC8LUrzu72QLDaERn8gZ7DJvJmlEOlacoquS/sDfPO
4CpoixSftkz5Nq2qO4aTlBDc/sF97LkSNiy9idwz21hee39uprhILheYUVDoDc39
jtfWvSs5pt90YNwxAIH+bxf4NRpd8Zr7T2F1opJeCmaS6MeKdRNRjILe/v67BXIj
pCr37OmMORAYHB36AuBzR959MEqN9fEsRbpHAqeTgmHXwb3bRTiBElUKsUuJNuFy
vIOo6jtTkTRYxM1uLQbSP6aSWlQPbGx+Xhrx8J+qJKGBStGYU2F0x4QrownX6MdT
ocVV7YdwjSP4ss4rMNQhzqU2mduf7Vqjk4cuwTwTIjBOUxQrckjpoMLAzfty8vgr
qg2jAxfpK576pgCSUkjuKFOjKVDlffeY3jO7jE/XNhmfinZR50ioQT4aI9ocH5IB
0Fcr8y5cHt9iPOe7kCCKlemKza2vCm6F99OODUJbu2yLRAge33BU2W65IUFVerfk
IW1y1W7uAIKzLVqKJpFiJPRacWanySGpU96MdLEHUNctPZ0k510kdsi2a+BNp+Dn
ejlbpLtOQhdEf9XDL96i/4KUTei09JDuq8sT8UMZnPVVhD4zuS9hZu7sMTTtqQTc
CsLS9OaiKPaEBaetXFbamNaX68nYvcYzC/2cDlNrsTuy9Ry/ttMcWOYqFjFNHom1
/v+h/SPW/zKRaKDd1aJa6pcpJHqpVx7BeZnhpupJQj47uXJFyPv75a1yiUPjYrK+
7Px/dBp/E9njEz50A3aSHg==
`protect END_PROTECTED