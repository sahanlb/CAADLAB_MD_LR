-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
lJfbvGo+C3XavN4t8MpCA9j9ORHjG8e7AOCYqRnRA2imu8I149lbYm+Kuel8BGu0
dJLGntjdJjuoYwoED8AQWkKYghuXZ99ujnL8bKTJKSN5+RIKKYtPUhHTyDnIUuZS
xwg44r2lmapUBjc7B4uUtDFanM2P1Zv9+p1ZnTumh8k=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13664)
`protect data_block
6Ehrn6lRVIEUy699Zzc78b8dJRG7OVFr4QmjVgVPxEnFnC2W9AU5Xtgo0/AQEkyg
3b9rg7pfwg7QzyVB1bak6reCaEs5vUcEIk4BuMQwmOnWyl1i/ZZh8v3hNsedfsZX
3awefOQMj8tGnt36nPnJiyAHmFjt084dd0Miuymozt3DH8WwpPWbkWAUthRfqZDe
12uz6eMCfqZzssTtL6nXx1HNhnj5c0xAf8GfZ313NBBazB6ONUhT2oRy00cLo1ez
NLjJVVHCqw5Jqy7i8Xy/lwUfqNiGIhq31kMJRu3txmMkgzJWTU7aSb1RrdXtPT2s
qTaLuafYLlmteFw3U2BODjzEQMx4KxsuWhkzfeS0+OWBIEsrk45aLfohloqHM6QZ
qUPr9x+OcrMScHwPCysSkjjiTMjdZoPhOYR+Eq7X0AmdICovhXrBprb01mmBxQqk
s3yjMNApqU/dx5L05INSEUnDsmICbVwn1SBRYZGeiUBy/U9ugV991T29axIPVnnN
ENgJeJfQnggzc3Gd3XW9svyZHkpIU+iyVnF1GdCHQgNl/2JywIPKF68oQ1+PnVny
ege4pMYgKFPt2TgzAxVplC8WZOgF8zwTmrjAkkuVv/1xJcWIoYgrNK/j++VwRRWg
B+aicjW4enzy0+AuBIYHIqIVo5Nmrc7mYjRD2K1B6dEVuiW1Yao9zs6NVnSCslks
UC9/CiPd2w76x+cJo4P7sdgXfFNrb7JFWgouVQ4kcI+mcYgGT6GrBoDsamPI43Me
I5IB0RrzbjF39cVOCk3dlu6L3EwSSpDU1UNbY48C6+ebRh1jsDeCRiRum5NFGtJh
uSjKF7c2OrWYQAGGkrDrinKjTrKc64suSyT4q8ik0DIgCPWzUSWHvj3q4TpoPrmM
OeCjlA7yvyGcCTD/rkE81ROV/Yc/8EVgZlst7j8qJJ/CwBpi01gdp8OBcA7HIj4i
7gSepG7Jh0v8A4JXTakAhWxIhxCEK7eZYrmwTwqANeNxwGDPLpKrjO2XWEKwQX+m
kVokQ3vtg4UtM+eq3l5uXFS0EXQY3AZcUgV7co+yr7SHvTzHnx7wWRckh4ntYd8d
sa3bW5qm/uCU2pdQD1Xyfp9gyDGLAz1mNNqEhQfVjO9IiJUpV374jWv8IgqQtGrY
F9YUr7tSGKHexUAPaXpqbjog92iWCT5cKc0immmAGn2sPIoEq5fAs3PuCfhAA/se
NVxj15loTbGQrmyeVhS9px4+vvNTKQyQGZ0AbiCRtmtt75ih23p22C3haiRbN/pV
OtCQWS3FJquZD9AtSCM+f5xOxE36GgFPLhDdP6XqptQALdUeVij/ooGfbz21Qtxa
pVVpzOLbLf9jGUd4QDCYyWxzLqY7Guq/mvcNDKWG1wftjZZEapYp9HDf3Gi1dp5V
ZuOt37NQpuDfFX9bOvv5FGyoGjTfHSr1xYFTh0EKzxihZ68+niGb0KsoQfdGhi/p
+jWIKrYP8dtRgnvkR+GufviYpOdLJdaF9UtDqZJ1d0DjCcJqCD2DuvgU6KhMApPl
QzjXTEepwQVPs4l8wZlENRGAuUTM2PWiMOWezA9cKY953Nu4DyOZhLt6Yb24Fih0
sAzbOTqY/L9LmfQcM4LOUi9xu0LiCqB7pcKb7Vt3SfcnAbR29C5ycTwKkgdqMaLm
EQ+S1daqpdweOUQM300eroEIg+PAwWLAQ4AKCVPFYdwjY0HI/xmUdH9DOIAVw6pp
MpuX1vkK6v2LZt/bbIxSFZiImVShIshJONtA1tT32A+3379X7BeERTNwb5frEMis
UP3s2HB0kMkG3TOi3U6ketox22h9HM/1yyELOLpbNv7DA5sXwI19uH60SiLTlxUw
/UREm4QbZBh0r6WicsCGZ2fSpW24BcIu9zCxNPc1kZJM6sYrNLFmSrglA17BC3D2
TK3SSnQbsrzia2f3Wf62k4vnfik3+Sjnt594p0L7KnBz7R81twxxipSMvM3YIhgV
HPwNuzVV1C16YteZLG3jga/WIhyUsTDir2awLcKEb/iszb97ytYzye+E0rBC86j5
YZWHlYFQD5RrSlZpfap9tGh1UMuC8Ney9eehXNy23UeoMkLwrKEAFe0FCrG7yoCO
ggAcGnb/K9GVxmj+prhLBjnFNx5eHOfLxKpTsmNRkGOAwKitri9/lEAq7irMdMkT
8m80ztl+UogAyqDtCz2x4obUcYPeZlb5k4a51V14TsdBo4kXc3KA6Z4iQQ20TXpv
hhuS6Zu/chpi0GN/GXjvR8zjupnJoEXbwbgbCiWJeLK7+YoxuZzpzDSCUvbpF1QG
rpSesqLBDDf6TMM/lmMQZJjuplnhjJWYMJGHobeC1PO7Tq50QpZacFfGpVkz9y7n
sIDfkyB/dxs+6INzwZm7zSsYmFYVjXFp6mYSJ5Xua6RfSZRDT6+clgTH7l+Ou+2k
wUYdwV2CwGxcXWy7vR2ay0HZB377negyLWJWf/Kb/BPjaaBzZEJigun5z0JZeDlb
CsfjE+JcmEiKTQhURlBaHq8OL3HNdwhxFG6boKuWw1XJUfuzS9tjgidkrFE64Mww
vIeSTQI2paitEj7HC3Fs00Pvxm0FaUxcADNggDGMjxENo2KGS/h96zgETZOCRmsp
XXy7jtcgpX2ZSuG0VNaxCrJe0eiby05c/BbjH6DPws9yOd4c86FcKGz+HBSbGfle
dfqjj3g/gSDUwaThycoL1itsqY0djF5RxafNePjjPCLFQ6uGcDJzQFLHhkYlacDg
HO1htHXvnQqgNpl/NlTPdjChCTldzN2prPHndPv9Ad0a337T1SqpvGbsmtEmkGmK
gx/IytrlNuq56jT9Q9knZXeU2sZCRsIjNPb6bKZFur8Vl5/5uJ3W1EAUvqHS9zQJ
khI7li8G3vBcJ/gbhzT2aNkpjxuxRpzyCFmXnkP2dYSFws/LRDiM9YJjwAVOrs8g
NPtopxLETIuI59rputrplj2U7uhNLU/xXpT04NAFmAq78t3HSmRL6EKWppmM/uo2
R7yGVfePkc3AZiw4pq/Q2dalkc42VIHGXqFgXDaVqeQbVWIpdjVYEnEJKURptY6g
z94/zprp6waLzv6zBRjrekDlA/y7LZVccKvEmm8ZB/birX/5uRROvcQlpyZz+o2Z
GO2nwp+GMper2KZ0VJb3Arf5/taJzaaPWCy10xbZht1vG8/c/zDYZ6EecmZ5UfJN
Tl3BHtj9nhPBZMCsXKKKdQA+xhAfmtaPo5lKvUHb4eVjUaVEpqhG1Bm8eGRI+Vn7
RnJsWAyEojU0bXo3Ui/sv8GUhjCy8XwKy1CTYiEVAXGBgvYzEwRpKKXN8rEafvA8
kcUOmt7i+UPX/1fMHMbSdsoMhte7V+Fd+Q2jYncafBeFiU1dgIXrGjunW0wlHSSG
xxx+lgcpHhzzy1aWrDTUVL3MeyR0vBL8QJ3e975tWoq+vnrSAvHm25FU/i/qLLNl
Qqf9alXeD2vkRtx1kKwDUTmaPbt/wpr8/xgfBRPkaWK5oduIisyoHv7Q0NQiyayt
WWQOd2R/NDpDV8WKgisfXdhvKrbo5/O8AagUJ6Z31ugBJphLRNm41YOjlhPralPX
q5ixmI7XFOehv7RSxhW8y1JI+lO0E6CNtx2F2DUB2PjtqcxJJRGPMGWjkvBisRoA
hcaeW2pNIXc5meO2yIwofyO5c67+ShjPR/s9qEQ5lA8+8UW75OdZos/+mrdPYO4d
uLIgjNEYyP2b/jeRDJLVAf58Y6PX2lBD3MlZihepESfV8X1G+wwJQPDU7Q1xMi//
Iv5D1A53IDRR+UIga7aQLqJh1DBbk3mZ6vz9kuIgZRsOKQHPlk7/NPcvN1AF9BSp
+If7x23NP82bQKUtXAlCl72K4TZXuKB0RheLZQrVfoab7DhSzRk3gqxR4pyhzYwz
vBM4tKpGCU/itZw/cwTtnlaMQBavqpzXqblrtff6heEIGW1kC0KKhjoSAQOD3R0V
JyGAL4mSmytRFJa7BpyiQhJNGoB3teCaPahtIUzfyBPnW37+Q+0HMYWo+7Z8Lsid
3v2D8uBTYl9qlim7YK+4L8pJG30Kd8kWacOiNqR0dDgxqzo5nfsX6e5csdH5okSk
J7e4P7lF5FeymWDbo2gA3wbL6RSV4cBxBswQwclpLeFvHhbmhmpKSG9tx0LaWD/A
EbswpYeB6cNEOlxghxCxxSG/hKzNT9XCMV/AzTWBf1LmA6MjXy1WdaakdiUG4hax
qv04DA7uxckVYCuD9z7AH1rZJhvgOO8CIegwcwalNSJiA89ynGhGsMgiGd9Ln92P
oDJfOUq3aXU7lQD3Lv24urvA4u8wKdZ+Y30gp5lRdS+8/M63c2vJqJsU145mj/Go
uriTl8fDK7AQYqJGLkhM4BAJUYBf66DW+MhWjyZZeRzNgE1xF/ie0ztzfHTFBc8M
/WDYuUlOg4r8nDz5TYZjzKxg5mFC0USJjvEA6lTSjhL+fd2oo44oXczCl2mHvlqB
/oXKjvav1bFYEPIe//4Y3J/z5NxkaSTtoAH7U91iUwPyRAtk0nhbPXB4D6ir4S/5
u/5zosGinUjyDDq32BEV/ncjJUdv95PA7xAvFoARK7X1QaacCV3gtNXuiamGUMfe
1Vyvt/my8MHOgeWCOlrDmohNbKCHezPF9+ItQQ/MuqOUhq+hXM1Qse3iDeJbcQX/
OOU3CrNSpSCl5onknEpLgN2/t6K1ANTzPGIiSI8Q+kmQKN601uEywXURcvhUl0FL
GfQAycGjfhlZFPG0dQvcF9LzbfNhVhQf4w1Ls/JYX1RUInR1D1IW4620VY6zXecn
HsNIhCyaoWaXbFT9rRmmHPCwAsRN9h7PTE28+I9QiL63c9LByjS5VASaSXKEay6A
ACMDzCHmUfO7x4/CtcciDRsOodmRAvys9wl1XrQqIRRtOgv8J4nuhzhvDf/pPX7K
iQ4lNTEJA6Z/vxZpfXkdu0eLnqVVXe+V4AQzBkwoEe1kOvA8CXm8DCm7y/q81Eam
hr4uEp+W/KKCNWCPUw7Mf3WkxxNYuqppEGXs7KXdha++qtqT+y4AyCBmRDxd/w+/
R4X/KLAfq5QY0wSMmyFktKQoIpEz0GhS4TqCAT4pMVkSMBc8u6GL9KjnHW8FBgvh
dNM81caBLpLru74GKirCuC8QMEu8EPLQuVBECxZnAnH3N4EzBjJoemvkdgyPfQQi
YjHJl2zsMZ0WiE4EO63244zOpFEin5wJoo9ECSp22N1lINgZK1LhTpRXyfc0HngY
hGafF+sb+q6LGcJXfvbBV464Cc15abd4VLsFShyEGHAkmknJz06F99zw5m6gkWz2
D8SPDhsYvJTpFLCxjfoChN2VJPpWd0jtENbiAaBGPOwzxxrC0XeCvd3xAOLuDZOE
i2/bEpFvrlvTHH+AxzwZACKW6k5ynswKdNC4tqMed1+dMdNT/3wv0hKJPuWjVnaG
FzdY3PDNkn7yT/lhV9KmcFWE1eOgctr2JWjuVW9IoOK8ObOjMfTTYT9F7F8A9zza
FhZFloeTLUsPXxsvWDDR9PrUpGY9y31aEq09jYIipzmqASbIKYv5JephLIJ4anwV
kgz82VHqg57kKnGLv2s1YiAHv7nmZMtPoe2ntH5Gum/ZZIt4nlN3CGRWKhFLU4Xx
GkbvEDXpI4xF6oFJTaCY+Pgr5m4Rh7WiU2lGT5txzV7kQFD7ac+YWa34aRgkVECA
jK0mQ3ZmatN2Wo5asGRfBoSdNKgfbPFQdAub0FbWImIEZi27q2aj9NVzWi6VFDbn
D2D+qzMIFR19GKeu+B5HIV2RX0gcRL2kqVXqYBE0H+W6bTbwC91FgjqUm5LJc1MN
Bb6Ycpzwsovw0mR7uWX1Z5fx67iueUgv/4WwhJgANLRwiv0rTJiUoRWDxENCHR8r
Ch3qZDKVoBzQsELKsnv5KTU+fy+Ln/hRkDGaF6+bzLwYniiM9pXf9wq3E1LUA0fh
ymIYISzEQm7JvEH8c2UfIKUzSwenOgHrFChNPyIe76zYsx265dPcYtCHyR81xANH
9YchY8nPNxf2uuPyEIbo2lZc7z/ybQGmJ0NQ3V1QvCTMe1Q2DxlisjqH/Ynw4n3+
8UuchD+XHa6/FdFMvrV0PsEDwhZC+7MQj58Q5IE5Lj8Q04ozN92fFbpj9eKLizX2
NKK9PeUgVjfwIG0L0IlS+/jMRGIOjSlvmX+vhws3sa+G8izoIW0Q3eh8MTlvrL0b
xfTUyQx/TiEPWfn3pjdqHyd1iR3Y53u+JSbJakmNSBWZYaWOq06EGfGnukSW/OXr
hxRL8RgbFLg42WwYO+4mUZctXAf1hrImS8TQAm6c1Z9p3zS//wbVtxP7xr9md0Ex
wvy5rZeFTOJmXPtwQbGsY7Fg2pBGB/s6ztykT1K9vvMRTnnyb1hDsrF+M3V3fieZ
dv6YyA6VqlafjAPlDydvC1p1JMVXkKUG4HgzCuv84951ufSgQVfis5WSM8EIRyZ2
KHoVRG0JKIioMT3lokbFIGdPfP50vDPmh1X/nT+sOEG/6iHeSp/hasZkNVE6pG/K
peGDZKymPiOBBF8JQEYErjgfgqr1iueNJHAJ5MHFM8Znwd0Fp7FC+OVIYdvHn3vi
Ije95Eb5+44YCndeSe+k/lHDcbCKHMmQDNtmX80Hv9F91MgpDGRAK/gMO6QXB5uX
v+sDhnulAxM0mG5WFa1kLHynoLpfa7zs30aB/2/uinUdII5GX0M3LymfsTgM9sE1
Noj/Gqf21H1BYo7C9l/iOP2Jfiw8sBVeyC3RR13EyxlUgVZrcWqDE0NbJtRX0GGE
bfO63VTksDqT9LeU5bnMBAPZMkvH6oRZFPFj2lchKWLUY4uOQa4MSAVAMZ9BURHy
n2qQT5zfyskCKJl46xvWgkrynecRW5r0CJ9FrAxTnVQ2NYd0CeBYY4eicgwzJJRY
ZBr3aD3qA9zWnldeZndK80k3yjuedZZsvmolyBAbq/eC68AsxMzYXxd2qrINAWOZ
nSCO1jbeeGpLIT6G3DCjUbawlJ8UXC2mDyFpc1bOZe0v2NjRCRKQiY16EzXlMlah
Gn9AKarpJzJ0Yl3etiwwv/6Hhk9f7zVnBV5Q5LNxiofxfZNTrdP8LvpR1u8NONQr
JvKVmzuRi+3OaUP0cscVwW1m0DIv9nCtsoNktxt+D7YJl/LtlQljqSu+eWqs/MVp
VxfBmkfNu2+zGjkNid6VN+bqLmHbQYFOPvJbUMYFtlm4JxCT8pVsrMEwN8u/RqGT
VfnYGB+xu1SgCrfQvuQBzSFaof5HCI9T0YeaZi0eZtgi5RfplpL0vQAfsU3pbV2+
12wJ/T42cedh8vHTkdKdU1y/schCH8/LBrVDmhetFZ1/s9NEttgNIH51GhHcprox
uWNiWaPJjKQL4m21eqLXyk0QQmGMqwohLB0uwddVx4Q3PKFQ1iRVG62kxgGFhTcF
SvzCyavnoc9oj4OLGn/n3CavM6uSqP/LpsByRDyXo3RUpjuDDVRQxMcuZmA23zwk
ftHw4sSk4b4LTWvBLtIqJ7/mWGCit8KW8rpXP1Wua4EVAwPaQIVp1UsB8tY3eHR/
Sh7KOYR1vaUx1fTKmPT7uJvYAblvrJI61+lfFvczAWFQqXw3Vi2s5cIv/NzuUIr9
kv109Oc0wDq8J7Ze3CGsSN5yrDehDwnAKYRg+kMiFqMZ2bUaewyf+Ehi5GZbkGIE
ZIhJa5OQp86Wc/1J6PME6k5bdtz+UJHpYV0QDytSaqYEI36y+SsRZpDxMNjaRWWh
XHY6FAoCLu/VTGCVq8EAmElbA6OygdpX2iX9O8sgj7voUzbBBMOgc1jeKUiRf5Jv
2GBBGSsUMXZ5CW+tsWx6pOQyjesF+2joHLGAfqlPWoqFOKuIR74l00eLiHoOSaa3
ToZ9yLbQUFtNkW/0ApuW1765Cz24PHcH5YM7g1tvT8ZLekRPH0ZDhahDrAfMcIjy
lDFWUJekGjEp5HeP6nyIo7PrAshoJ+Ezhc5LdtOUi9UO2m/z5EMJiDIr023Kk4ex
9gYDCuPnTuMftrZN+UT+WsqUlO7zWq1o5xub0Iqp8MUsRqBlFiMVSU3GF7Xgw8pA
OcM+Tgo1o8WIi7VielvpBXxYamJRR1An086OnQysNnF3ZQ1XeIiRHfx3DH2An+1S
c+PJC3QqN5unlQtA3lsuoF1ZbjEgtQHBHmz85fsTmq8NzMEWHtjumkxKYX0MqsoZ
IXX3KQMf9z4Fk91aiE4GaZMmNSj84PAlRdtKoOIhEk/lA1Io4U1kGOgoEDIa2eqc
A0x7g6ZhtNlRZAcjbZuWRg4w61h9R6UY7PF2VCXv7zEQKMHj4aA3EuWTZysQJD92
OQTalgvSUzF+xt6oZDnIQgOh5cdMutMNWxBEoRjQJ332A0HEvepVa2wYga/159Y1
ASHdpfqVPy7DrnkGPcUWkIRrzei/xoM+QlpoMpdycmPlsWObP1F6/n7RTgHjSlV+
4S1rc3Z6q2ZsQH1CohqtFh5+5iqT3BHSMKf4XQqz+WfijT188FG+3yd1GSjgTj+O
9H5aOuxyKuNdldvOIOqoONSCZPDbB1mjvCg5UuCjX3nx+G3WHGrNhpbD81IsWuK5
oDbjdWIGbBRE12Xn4NiBDEfV+xeJlmpDoOem5cr4+1yTUoJX+1AbR97fNNn8xJck
pzuAa/fT+gvzTLtIQIOFar19ISo1ZXX5YcdFL4DjOj2EuvNuc9J9FHlAEnR/0DS2
ADbNMgOqocODsFGp7h5Kjzib8fuD25B6jAxfhZA45DU6dyb2qMdsMSlaNjkc5uSc
Jbts5zxUZ/jVpgzrLplFysP00OyozlajTi8Qq5ObWnUs0LnN8VGxpnpLlpwA2N05
bqEy4bFjfBdqNz9AqiKS+8TV/yjWholPQZuxv2dpP6PtTKmTBmrIKN+zHHAFXcru
oNRp43h/Ixw4Dua84PKgCAvoIem21uogQ/h9gL8wGkpqxMiB/VzjM7PP2tQheT9i
nKyqDRk4HzpZi4PwhCO3IUosrsGUJpW//KrY2HZUVSDTTm6ZsmBmP+oH2Rw8YxeQ
JShP8sL7VlaQ0Bvs4vIxMC4iVCqBKh/N9tIdWdGmxxbr1p55aa2cwYS0+66wrTUx
w5VfPfkOnnBPWikXVNBka4z1+BmWuLIiAJdlvQABz4c108fcASxnDosk0X6yyuyu
dz7yl2AlfP+Jd5gygdr2oPUmQSQ6HWHK56iYauVkw87clfjpVy0kRGQDF614ObSC
k2lN4M7IzuJP2rO361slftKnPao3U49al1gZBHDVuY3SS7sXktdOVqCr4cjJU7U/
upuSvbB3d/N/jBcaqF9zMZMJAGxoaa4XMpvR4cLXw+Iuvgw7TxsVrPnsF7RYK3q1
RjCKEvHJ8UzIDjRxENl7oSrmszyO4gn7kk4iud+OXP1lckRf1UwgiSftS6wj+6MG
OOlSPMIhVhWHHy0YpNO6h+67XaXIMC0nOw1SfQj8s1k404un3K+xvGNsv9HnvDRb
Hf/Cc0chvLLKLrYgLDItLwNX0fc/vnGLlZi4tCnbqyrm7TPiOWwIQEbdZzpLQb8b
gsi/pP4dbrl50qeW0ZtT5B9yYhLWIzxY9TGVwbuXtAchKoH7q3jqenq/s7KGhWRa
cNBNWgMtmCV//GTDPFjo25/1khORrSq2v81bVwxljZCaUWlPlsnUtayHJAHSr5VM
oFuW6Sd0s/YpRwW25U3Mgf0xN2tI26nbTJThlojPr/453DdNL4FNAO9pNfvEk7jm
X0ZOV4JpIRntMgwLKQoqpESpZ6rS2NiS+s0HV+hp9VQyGhrA/FMOWaIivS2aQ4Ey
INrNpKc8h7wkaM10KYQe3lKRhOFY00jl96mjuC6bwvjBS+SDMndCpWXm1JH7oB2+
5BXe2qgENwGGGk894LGcVLyJrmkwukx7Gbbb8am3aQX4q8tQplD/EKGbwvJgRB22
32OlQ99ootGZq1Wgl8o6WBYkDd1FPSRLHVvqf/LKg3K5/eB3+9LgJY5F3TMCMnAh
m974+sR6AREckL5olPppB1g1ynu7PCEuBrZgohAonheH2A2Dpjc72C0qukCodqHr
lQsjduHLP1TvXxpC/VK4I5dNTqvh6xou6d7JlJjnGhZJzGJg1ctRhsG/G/x7e6QC
x5s+e0klDNhZLc2PrF4/EvnQQfU4aDZOFvNFrApxUbbZWbpK+sZ4Whkq0gtNjao8
aoi7sbFvBX2FZ+e/EOx9RVxagYlry098KjOohYM5pP60m9d7JqaSFZx2f1kGSl0D
OgO6yG/iffKSdBBNnxuyHx7T56H8tk6GqVu90hSfBuVzzmJaV33kU9//OOvvMBZm
10cktkZj/IlLbjZsIq0a1ZNH0wrfU20aWvX2l4wIOE/gbOmNwi3a9c3z23BTO4KQ
q09UceG3MLJFqXu9H4yp/VWpyhO0uCEzz6lIXcBoWr9LCmCuwC+MVzDLtBmESaKD
68iKebgmxkGRowoKrj2L4arsW2T7fNO7fn475GROEpp5lIVSjW4vKWVTWNOC3aGa
uKKwt9fEawHcCzo686VBYeWbvSN6A/pJaQdRMrybLgW6gg3x4BnIIY4RLZtxwpFu
XmxVFNZiYFa0SjYOHo/ke6MDDex0J8iqcxHx82sl9cqWaPtZj1XZqeWW3w3eeHaN
Zzn8TcEXp1bWKXGH7p4VxS6cybLBXo+xcRC70/MkisZFHAIq2ocyBbAJ/LtPsvMn
QGuszK0bOAmIwcth0XXbwdrHb5CAO/la2m1D/iqWCekO+jn3q8uMuIniGx60ObTA
ZoqsCTQgRBRyRSuuM9fUDSzCPhc0JeUmIAM8EBVBXTRMOu9Ajf/dGPjiwh9Dfpry
0d93RzYkSg5nJ1mnMrBYWUWXfyhwgo8EhBUUeuHgELkbRg0mhbIBPG7/wYqkExXy
3gY7g3jBE6hceDVZXEIF6u2dia+45+o96Wq5wNP+PV+1D03Su5aeS2KbfIQeotjp
NFGCbIUZLAUkD6Z3wyFy8N50T9E42hBDWl2nhESKc+NE76vgy0KNhwo5oZpWZ9+L
fmqdCv/0da3fJMmaB12CJA/6oAz0Mz3LQ5Kke4FnNZ9SJRoAj0AHkFSN49it0aHL
m7cPZra2bzkIuZqEyj0b1I3g7epozY/bw7ftN3C3vdSGW0S/29uLEDQtBKYfyeD9
EHDbosmOJFbcm/PeErEgDaLag44QmU1bb0LCpDRhxTN9EN0C/RTNxtJoQt4c0bGP
xYeR6e3pfAQhTIxxBAC44hazBkTNA5zS4/DwPOuGJazSiTd9ERrNLhqLRDDvx1Eq
5xGSeaGjZ30onSxjnHcNntSuLkM8QIvLMgE3vKL7GqiKNlhu0SLROE3yLb8A1dA7
1PhpqRFtRUb9Lk7TaC2U63B1UHusqYD+LiN6xw8/bO/7DfLOjTsVTc6KA8JZ6kb7
mSQ2sMGMs+Ey0MBbiVvtjCtRvNVNBKx2N1L7S30E03KsTvuds2lKdxbCzKftnlmz
ktSipXSh9bMDY9HgWSZQ9xgqHJc6b79H4KIjMW/VbjL8R1QQ8WvnRYgQ4TxfZ/5y
cpt+7iGi9iB8EHAyvGUnp5Gq52rJ77KSKGQ5/BXOJ5hfn4FvzqPWexAjE2Dz1omy
F+9LKSgwNzuFEfS/PPatTVaC7SJbu/wzDyDA81e7oZBMeLN23MyeODYBdstQ87sy
GenMlHtk281hBzKj8blIwmmYgi/ppsLo7ZO/dMnrbucsFtqlwpN7obHv9n+ruYz7
NZA1fuIjqdjORUzpjBTz6j6Jhr+Gmg1GDUVuQgwQHwTaHQeBN7lxHw+4mxJ6DMrr
7G/K55WJgKIKsJ7XOhTkJ9BU4KIqjx+LdYOrRxBfXEJIBN6aRRmqi4VdlJEKxWaC
H2LNYn8myJcpFVlZVUsjsBGbnvlHBjfZOnl0dz0w4WM488UeKpwJI4mpG+r8vbO+
6PBn+KEfYMCzPqi2jnaTkpf1s0kW/oq1acK8seZsAiMxh60aM6Phyk/movnGDg+H
s+GK2B/UlqfuaJX2ISYpdVK8rV/9W9ofW7j/8lnNukbURJeMNcBT4N5bm1P2QbN4
vjAEsl4Gcr8npWhUBoW6xvAVPa+K9S0sUBUlvdKzPPg5i6HyUGB++TbZJBsVK2R/
hf8cqRNxgWWRSX2sae8HOy8XtX2iU79Otf7NeOBlxmtTUlXemI5xykYW+avTCYy0
P6hKv5ksaAC9EPEU4SlxLjva0kWcC7EjqRk8r1WCSB/zxYT6wahjKRskbB19VoPl
Sth6WDpBMZuXjD4XnlwV7OHhPn5PKAWN//H2xWnUo5xrEJlV2hfljmbp5zKDHaqc
tsZzh3EUzRdzVLySUN+V6hGj4GX6JWGJi/4qOz+MpK6w4AI2KZyN3/W1w/CciL4p
Hb6u/mERk3/0OgSjvR0kO0Liw8mR5UVd6yhxusLxnZSvQS/9WtqVZPWA/I9mt55j
6926uQDLvUTTjOjjURNTMhXr2FKHJwsPgwrqL6XvnojudlbkPT9vuU6WUjic5M4X
3bCYpmnPIAwUsy90lUN9ZDwUWyIuJBJreGKkt4gkLcPecusdnK5nHTNEZj98wUus
JYn7EgE8dNGRA1gV9wZ/r8Gn1xQaU/HdGK+41qEG0/z3Rfj++DiNqH+n54gGpAgu
ZYGRd9SEwR5SjlLZ2+yfUeaZmeYLOasuH2CBqSC0g7SIuI/dpH75JEGOu1NV1tLV
t4SRaAIaXrHS6jXOzfKjhTeftdIgVKOGIsp3LQbbxF75nWPnqFZfvJoDsTFaReR9
yiF0Sx28kUfZqKoaz9O0QSb5+Cw85+bWY6yTydt+xrrVNTTfDuWIUi9341iVkJY1
9kP1VwdJiALYQWh4gt/U0EqCDgwGhE8D93r3yQM+L7nfqasVlDx2TxMgRgJJG90l
cg3W1IcqPz9UN3RESs60KUjljzQn/0Q/dnQIy1sVo4Q31S5Lg2qX9GFSG1557iv+
Jw9dcm/4wfEtZIU6cj/0AC5a7d+1Ne/TJ2fGBw/LNwIjxMDHnXYysEGOVv/hxSu3
9/DPJPwwsAww9+BNH7Csb7m7kUAUAUgjeg5H7B58328nxbFBtJwDsXq5AIIgioBi
/XNWGCQ+GD4ql6XgsShHcTcGUuLckrKSt5OXH/Bg8pIFPTdt+08ZMNr8RR6/UIe0
0C5aXgdJzXexPtrhzrLtpyq668XdCE6XAkN1QglPFKt09gHdD1DVzAypixoMRAYi
piPyuNj0b62+XzsCplAnuSXKuLe+iuw0lHi/0Y7MH9HwlWbAP6TWpcJtYVc6knKM
w9PGMJK5mTRxfiFqE+og+pH82QENay75FlM4/thzV1nOQdyGmuWdDKZvBMdSym7C
Cc03yCDLCF7FNVIm+FRhS1I1kdb+V66NdPwvSz/eYHMDB2phZHKeo7iFW3TWUxXc
7XUYv6VLkhK8J+k4EOPLkhNIJFCHbwXDUpTd/Sm9B9RHR57AxQNsBMxuJU6ooxDD
NEqg/cP50GA/pFxJ71zBu2PY/2gaA/PaYHXkQXaezTEg6itZZPRow48dlDGMOL8i
xtyHCqk3HTggZvCLU+Tnf32fJQgVv0cYEAi9d1I6TNMHOShiCIyxFjNyia7VYtun
/TgZI1+MzWVXo+NYohQMvfoQTZQOt6XhkYKU5sCh5oA37harvWuMzWkKF8hjaLQh
B3XvMf4GYr3bMti7lOg7Q17vMG5UEwGqZogwJqp63wycZ8zm/VGyr+AigCn+mTdH
MmP/QDMEMWGpotSRcIfHbm5J7GrHc2eNiFS1eHt4jkX0j8UmHj+w4jr2XW3nPhU3
pXjpewLdsm+DnXtFWvMavFtBl1v7dgx4yCFDrKhmsjtMxtkSwPWgraRBE0FU8BBF
QIvsoE0BqPkrWb1+wfZuhyJGSco1h86KIfQhvqU/UJ3z1zwoCmr/eTk3BkXCpzgW
hl0c+v18p7CoV3Y8zxPjLnhF5B542rCdIkSvWiEd4afoheN98gY+nhPa5DxKL5ZO
5dWOU0pTDXH/3COEan1pFp9HOLUmrALj6/HurOyR9W990YYDAKkdCCfcXLI+UVEW
d8MUg5iWqxVZRUBJeWVNn+q7FqxatxY2JDDyss3vUEr8OaPk0yCgoGTtm0TXAaPY
F7RamUufbJ5IfTDfldM1spkoPSiJJ8JJOyDGnFIBxyoHVWyPwc43cFm2XAet8ijy
MVK4+XkbHdv/Lcg/wtHRjVgFGH/QmcWGdET7tMn17FrDVU4leMWhgzL4E3g92ZcN
VJDtCEZRk+O8MHgezswNpEgeTMtyEo7k7jRZaEsEXL3jgSsPp2yOcXfy077LSv8m
fJLYZ5Q3PCc0zVkD4yRYaMFGXKcZnPl798gtsnkcsRd8RI7SJNPXgi4GmBgcFy1n
sdhIfo/HEaHNUlNG/dOYnWtRPhWOCqm1W6eV1cHh6WguLxVLtSgyg/G5t/e+FQ7c
zbt8drmh4emd7pdG9C+CWiZHi0I11WIWKdOWqHZJyrnfCo3i0fEqqV7URvGtjKde
cUQWxvvL1XAkHu3Mewa8YmELHAUzPySK3XbZGuTmN6kWBCSI/TjNtbWhlf5gmJZL
Hxlzshi35vHC/V95/0grAN2FqSYdAeQImGVic/YskSdaDlkg6r7X0wlsSLiwHV9h
kbUdOvSb3OOE/zusVB8oqCbkyfGzVHaKDhhpr7d4u6PNbwGIzFPUPRjS01+yU8V5
F+qsoQZhMx7UFyI1d3m1mL6LEAsuFbndWSbA1UnFVPBCjDIRAtyBhwY5EPfmsbsd
vVJYoZkklXBkzkmurcvkEGuDQpTHI2XzYybY5mi1clZbWtSFW4gfWctr1h86y0NK
bJF8tYs13lvnYl14JLC7d2iQODWgrHTeMCb8S5TLWzH8S4G5A4CzEgC6ihnzSbF7
tMTbuVZDEAJbO+F6DSnHYPe3WsgC418bgnsDBvWN1LlcVxyQ76F1s9mQKZ+8YIxg
5W+nTC0joqEbVsI1cVNuTMblDue1+NRsGE/dLlJcpJegoVOdcoYJ7+IICP+OKp5u
UlPMbj57luYFZKMlC/4lILWRmOr9CXJbWxLoxgSYJCvzAlZVV67aC1UbE1SPtwUg
0cjskAETC1gbJZRccx7UKoC+jNX2UHgEA4AePKY5pWkED8A8LUPmpqRdrmtJin3p
MkCimA5Pk1A1zA/wqtv/VoNNCBE6k4hndVwBFUW+wT0ukkgwwQBsPUUo6SAF3Kz+
QjZhfDZ0RsnJFOLe0jJM4IoIW/w1UTDxFsDwbeIKooajfrjsnmtGCVAXm3xkquBw
NUXsm3hphhzhLQMbkYb2+NySQ7z3GMlEstS5ExvdNtGIjh0y7awMOLLBVL93KJIh
a6ubaS5NUZD0zZjH+dmNdKFZQddgZ7WhUL6mbZNe4L7VvBB5V7/iHJdeVg5ivhVs
8O4A4TqG0D6OlV5k5YEqn+wCZnVwUR5h0yZ3bJ6Ta+V+W7/MWMm+iEgv7lyz7rtK
m5ZfnXz59HugHVrAbYi4wWcGwt9u1SpRzv1AHc5+w7jvbjyScZED28GkOWq5adUn
tBaoa2x0iF5mwRP2iHesvuHWONRjXzsLfmmVzO7mDUl6knBuU3m8bfmXBVg036OF
o2lEL+qeyOghT5OlY/hHV2ccCqMQN85ouv5vMpwnWWvqAeuultAm1NV+oTETNuEW
UUNXgAkjFLaAxpMdkzjCmiLQ1A6tbgJqCI8nplVk65k+47oKpoVAcivmpMbmhcuU
jXDYs/fIhjYKj9UZhDcQnGyKNhkAuRIs5sE71gERfkplUnoxdebLZRDlMbxvrQIE
W/H9qOk8pr/9MJtRXDj26jojMLkZajMT+AvT+vIMBmqPyISZQQBDDd6fVeVCwDgQ
j1MDMD9WYB4uHEhNPMM09rlhZZGquLxwWzNSuOvWQJvzjtKScb9S43imGsMwe725
OiHBIdv7JJQKswy47nl31LoHH12CB2b1LgszTVgSwVpKUxfzPwWQKziQzYDg4vLv
12m7XKSo48riBfpgJOcqwMV+SM4KjEw6ZH3/6EkNW2Mr1z85MXuUbp415ScdStS/
UBGNlRVvobgSP85vNkwNrFztu5yNLX2unMqJUZE61Ty53Q+WBSf/rcs3FDZvFXEj
DS5cQhUPr0qWmY/L07jlPaS07r78FYEVC/cqZLwzgoJL5mr4+x9vNFWfXQ0zjmUi
eUu+KKFwoZhGhuAMDBLCAttco5mMfmANJ1x5ltVbYjAX5+R+O6njgj6veqzAlDR8
L1ZsjFILHTwU9SuHaX95CCQQRyFxFXnt4Vlr1tnLt8ZBfMJudDqxVjMb48CeaFxZ
jl+XE4TILxdHQBDjeR8yDjkj5igDNBDgtRpr6n++a/wIawfEziV0792iwYbg0Z/j
SIOwunR8PVbFbscEYDja8mMnAe4fdAX24r/73UAGwNNkbEPriAlYHa3sBRuQMByY
OX5SvAehlrEon99isnYshUreyY+ClONP2Z/+Q+awK7gsX57Xxy1QWHyBkUsV0Tlw
wWo0JQkJEN8ESkuD5DvX2Fs6g05cMkDw4RzqTwoTaGL2ENgkapuTZ7FmfoK4yWH1
SRKe7hfe/+eWEGQrdyDqUm2ZZX2JRbZsG9eKXv2NrAoAXzslmalwXUIONJWHYFHg
X9dCt/1x/KK/moyXNsM4h3L4K3+2I7BK0QpS2ki9H2kJPJCt3SgTq9Q9wVWvEx+u
nXLfysXw3ELmMe5iyA+LQhW/zaBp3I+LywkgosfktmMqRFCuIJfHysSyTnCD/PUr
OlMZFqgXvJaeLhHiW+T5fzC26+YkG4Nz/P/XNYag5uUGNC2w89/Y2VXy+S3MuPcz
4c8WX3FckH/PXUdNSCHzGYItos9GX/znO1icTyxU++8SvKYp3YuDbG2/3RAMq8h+
RjZL0ZBB7sQDexemyqXlKiQ88LoyS0Rc3P10QXApLvBCwLqq5ob6+4j54J4t7h2l
5DdS5eKMzkT3/Vp/UFbiypUARS9+C36bin7A3sQYZSdZVAJEEqe4tAprMP5yaefy
eSaQUTbha0qkn+kp8JlkVuQDbBAQ+vNfMVog6UoNTHDP4BZNK/YqBN6QWIrDa8Vc
tkFKGGKyTkH/lkV9qO0zg6KqI1V3mlozrkPWKckXCqddBLn96hcfrVZUmAoiiyof
2zklPW6qj0TfWKTaYL5yyb8kmptH2Qx2ILG/uZepIQFI26eDkKiLj17+TIyYVsVX
6z3AkZFbpQT3kUXHjZzMCUncjGQiJiWqeUG2pMlR90HwCdWmjLIjXkC3goQ+bWvV
i5cQLxBUzD3oZd2lyEtrYA1lBfWZMWM+l/xFCsu+DiM5yAr3nCf7vufQ7sdx2n/X
ACJbVg47H+3F5eOPZWo8viuikuyM6ax1mULQwxM38MoouRRNsFj8RK2gqkYC4f/O
QEgBav0ThuxaR59HdmILd9Wy1ZVpc+9DK/ofQH4oATZV/zs1YbVh4dJdDPJGYfU4
JIwT/htuwgfVrPVSMNFyUtD3sCvlpM5cBhqB16Bq5N4IV+ZjiEGnxvmEq33w9YSN
GbOT8OwL6cgfM1nlhEl7pys2AZEiQHaOPME1pjHZG1W7gOAEkdVn8FPJn+DKxC7H
aEDAqZGMyN1arxQVhqqZmHmoEAf1DFSQT0uZNZ/ccxyHUlpz5caaHc8PhRqrN9A7
LzTUZEnK7Vo06GM/A2zsVhCXWd4XKrubnrNp6BifkLk4W7OeTHrLZHv0SY8D5Q78
Is60vre8Zk5rPSyR4zSAeGuNb4raqbm2izSuMei98mLiNBEThJdW9P+hRxtOOSov
PS8GU4GCdb0odSbOfaI2bbg7pebLrp+YH5ga53WVgJ/ZeLpimQKNDZTs0kcl8Wfx
5DD0oaHrL/mKBqdjcyJP9Om/IkaGc2fmA4ei/0+kv/GAqjNNwmPTAq3c+mtbu0R9
YXlILTRwMoXOowDQ1U7jwXNdNdAFVJL3jW7ePNNkDRjIsp48JBFpm95SfDmQCa57
xEw0pFLIu4MjPic/kFAr2p7bMONpg5EXFo0u4TxWj3qrDNa1TRsuSEYZhEajTwmC
JScJTU+fdtkHv58m6Gbg+M1u+vRW7srAco4kdQGOKQ4my6upZzbg9qCTmqIpcPU+
3S1Re94S9ZSmSn7NOBmka1k8Zr/FUUYe8rb7tLnF2pJmCAWbHB7zOpzawsADupmL
uOPQd/dL1KEGrqD0xPaT3ieKqdxHy8b9Qp+4Z+lSd5T5KvO0msIggbXR4+XdAZZR
scoCY6pNpZBYjj6yZ7B5+EIVSG1vx5yNzRtev2vSdRU=
`protect end_protected
