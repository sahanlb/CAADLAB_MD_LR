localparam [0:65535][0:2][31:0] P_FORCE = {
  {32'hc4dc9919, 32'h41e185ff, 32'h42cce23a},
  {32'h43f7147a, 32'h420f00ce, 32'h432248b2},
  {32'hc4de52bd, 32'hc3cc86d3, 32'hc41bfbc0},
  {32'h44b97884, 32'h43570ac6, 32'h42a8140e},
  {32'hc41d0df4, 32'hc253c59f, 32'hc37635cf},
  {32'h441edfb2, 32'hc2854456, 32'h433af90b},
  {32'hc4432eb6, 32'hc307ec47, 32'h43bec45b},
  {32'h4491535c, 32'h43d43266, 32'h42312218},
  {32'hc4968825, 32'hc154db53, 32'hc2833a6b},
  {32'h44dc8771, 32'h435fd80e, 32'hc38572f0},
  {32'hc4a1f4b4, 32'h4346244f, 32'hc3403fbe},
  {32'hc39e4dd9, 32'h43240231, 32'h42cf9c67},
  {32'hc48909c4, 32'h431feeb6, 32'hc3c413f4},
  {32'h44adf11b, 32'hc237a027, 32'h4287cd26},
  {32'hc48992a4, 32'h43183204, 32'hc2b1c0b2},
  {32'h44f5fa34, 32'h436c45f7, 32'h43c1050e},
  {32'hc511e042, 32'h42ca7262, 32'h42907694},
  {32'h44a552e4, 32'h436e5cc0, 32'hc231d21c},
  {32'hc4ee69aa, 32'h43b72780, 32'h430903be},
  {32'h44eba5e9, 32'h43357067, 32'h42daedea},
  {32'hc5064d76, 32'h439a9a22, 32'hc319f91e},
  {32'h4503d068, 32'hc3912b7e, 32'h421d256c},
  {32'hc523f30a, 32'h4382890b, 32'hc212b1e4},
  {32'h43ca7b28, 32'hc2cde16e, 32'h43bd2990},
  {32'hc3a4f5ea, 32'hc3638f5b, 32'hc3689ad6},
  {32'h43c694a8, 32'h4185fd5d, 32'hc293a27e},
  {32'hc492a2c4, 32'h4389f74b, 32'hc392db4f},
  {32'h431a8db7, 32'hc21488f4, 32'h43e5887a},
  {32'hc4755e06, 32'hc3dc90a7, 32'hc3cdcf10},
  {32'h44bff9ab, 32'h41f50bd4, 32'h42653870},
  {32'hc4060784, 32'hc37a245f, 32'hc2b3e1ea},
  {32'h44c86d7c, 32'hc3297863, 32'hc34e944b},
  {32'hc50064cb, 32'h42466fbe, 32'h429b8c78},
  {32'h44e143e7, 32'hc2891612, 32'hc2a893f0},
  {32'hc45710bf, 32'h432ed082, 32'hc311588c},
  {32'h450fe831, 32'hc39d2091, 32'h426d688c},
  {32'hc41e30a6, 32'hc3cad3f6, 32'hc24b8e09},
  {32'h43d73ce2, 32'h42831049, 32'hc2ad6fef},
  {32'hc4ec8b51, 32'h42e48eeb, 32'h43426848},
  {32'h44e37e7b, 32'h43ba24b3, 32'h43844d03},
  {32'hc2764500, 32'h4314550c, 32'h43d74134},
  {32'h450bbbc9, 32'hc389625b, 32'h4305d192},
  {32'hc4fef33e, 32'hc3016fa3, 32'hc32e5cdf},
  {32'h43da3d48, 32'hc3149791, 32'h4382a567},
  {32'hc50e6c9d, 32'hc3a7dc71, 32'h4328659d},
  {32'h44a3f7ae, 32'h42a3142b, 32'h434c9bac},
  {32'hc437666e, 32'hc2ef95f7, 32'h428eb3be},
  {32'h45076ab4, 32'h43859a0a, 32'h43561d5f},
  {32'hc4b8fef6, 32'h437eb34a, 32'h42aca0da},
  {32'h4309cb10, 32'hc32207a4, 32'h4379648d},
  {32'hc306dfd0, 32'hc21a2410, 32'h42edb952},
  {32'h442c2419, 32'h435f2b70, 32'hc274908f},
  {32'hc43c923e, 32'hc3bb1f77, 32'h423b9b7b},
  {32'h44d1b36d, 32'hc32bec2f, 32'h439c111f},
  {32'hc43f1ac3, 32'h428eff12, 32'hc1e10197},
  {32'h43755e7a, 32'h43a89460, 32'hc2f51799},
  {32'hc4c3f4cf, 32'h43aeb99f, 32'h4320a22c},
  {32'h451406af, 32'h42a61c06, 32'h43797c3e},
  {32'hc4a3c1cd, 32'hc3818984, 32'hc3fd9f69},
  {32'h44f1f772, 32'hc3c0acb1, 32'h432ac929},
  {32'hc4e533ba, 32'hc3175ab3, 32'h43183ae6},
  {32'h4307ce92, 32'hc2ce6c06, 32'hc09651a8},
  {32'hc50ff094, 32'h4348e415, 32'hc3b91e91},
  {32'h44f54ab2, 32'hc2b67da4, 32'h421131a4},
  {32'hc46c9082, 32'hc3f5d795, 32'h42a4dfc0},
  {32'h449fb9a5, 32'hc2e69d7a, 32'h418c10e5},
  {32'hc50a2918, 32'h42b94a0e, 32'hc2465433},
  {32'h440b5732, 32'h432889c8, 32'hc3c9ee66},
  {32'hc4dbbf16, 32'hc24ef552, 32'hc32b0de6},
  {32'h441b7ecc, 32'h42020bb9, 32'h4219623b},
  {32'hc4d3ac25, 32'h431d3f88, 32'hc377e753},
  {32'hc2052380, 32'hc3725bc9, 32'hc168f80f},
  {32'hc4c73b7f, 32'h4280f7b9, 32'hc323d6b1},
  {32'h433c9f3c, 32'h41b075aa, 32'hc3791dd3},
  {32'hc410b71c, 32'hc2ef8f1c, 32'h437478bc},
  {32'h448564e6, 32'h4247ab74, 32'h43236874},
  {32'hc495aa86, 32'hc371297c, 32'h4348d0e2},
  {32'h4451ef92, 32'h3fd47338, 32'h4213aef3},
  {32'h438bdf10, 32'h432ea592, 32'h434cf678},
  {32'h45094ea0, 32'h4393a1de, 32'h43a220e3},
  {32'hc4010204, 32'h43343bad, 32'h42b7f8ac},
  {32'h43939afb, 32'hc2b9b1bf, 32'h438c911c},
  {32'hc4fc6bea, 32'h4347e7b9, 32'h42416e6f},
  {32'h452b7272, 32'hc30da3b3, 32'h43bf84c7},
  {32'hc5034fec, 32'hc358c7bd, 32'hc391db9e},
  {32'h44638f06, 32'h434d1167, 32'h43b778b7},
  {32'hc4978714, 32'h439150dd, 32'hc3142ebd},
  {32'h45017343, 32'hc2e6d989, 32'hc31582ec},
  {32'hc509dc7a, 32'hc3dcd59c, 32'hc165a471},
  {32'h450c6dac, 32'h41f313d8, 32'hc3ab9268},
  {32'hc421b138, 32'h41caa8f0, 32'hc30cb830},
  {32'h45023016, 32'hc373e287, 32'hc30ec84d},
  {32'hc4f44cb6, 32'hc3042273, 32'h43783fb5},
  {32'h45128a34, 32'h4310cb10, 32'h42add09a},
  {32'hc50087b1, 32'hc3982928, 32'hc37081e5},
  {32'h44433a47, 32'hc31cda93, 32'hc31b7dda},
  {32'hc3e83b24, 32'hc298b293, 32'h42e1e63b},
  {32'h441a76c3, 32'h43f5c558, 32'h4297a066},
  {32'hc38e6ee8, 32'hc310e3ae, 32'h435fbcf2},
  {32'hc322c540, 32'h4358a6f9, 32'h44074265},
  {32'hc4490450, 32'hc295cb8a, 32'hc28a8673},
  {32'h44f60d1e, 32'hc135307c, 32'hc10b6ff9},
  {32'hc408efac, 32'hc1876b40, 32'h43131763},
  {32'h433c42dd, 32'h43c1491d, 32'h43f94cd9},
  {32'hc504dc14, 32'hc31cf413, 32'hc2e90e05},
  {32'hc1f12500, 32'hc41bd357, 32'hc189e36b},
  {32'hc4ad361e, 32'hc32eb8a6, 32'h43303a8c},
  {32'h445e4264, 32'hc2cc6876, 32'h432ec745},
  {32'hc3d5c348, 32'hc35a32e2, 32'hc313ea32},
  {32'h44b4f281, 32'hc2d83944, 32'hc31bacf9},
  {32'hc4b38b5f, 32'hc36bf538, 32'hc359962d},
  {32'h44dd6b4a, 32'h42b92beb, 32'h4373f01b},
  {32'hc4e1d4c6, 32'hc3e5c86f, 32'h439d4b42},
  {32'hc18905a0, 32'h43743849, 32'h4355cb8c},
  {32'hc4f14d36, 32'h423ebc30, 32'h43f83843},
  {32'h4455dc21, 32'hc3a10ed1, 32'hc35c5413},
  {32'hc4a73342, 32'h43c167b1, 32'hc348015c},
  {32'h44241668, 32'h431ef75e, 32'hc2a384ce},
  {32'hc2f66097, 32'hc3cbb343, 32'h41594a0b},
  {32'h43fd34a1, 32'hc3a9a4c4, 32'hc331866e},
  {32'hc4c2c29c, 32'hc2a8cef4, 32'h4308a4dd},
  {32'h44c0bd3a, 32'h42352a28, 32'h40b598c0},
  {32'hc411629f, 32'h4170f270, 32'h42a8f880},
  {32'h43bdbefa, 32'h434b45b7, 32'h433e52ae},
  {32'hc4004b0e, 32'hc125c512, 32'hc3b6ed9e},
  {32'h450c53e7, 32'h43738209, 32'hc4063a39},
  {32'hc4e13860, 32'hc2a949cf, 32'hc325b774},
  {32'h44cdbefa, 32'h422560f5, 32'hc386c999},
  {32'hc4ccd7f7, 32'h4305b70b, 32'h41dd153b},
  {32'h4499a6dc, 32'hc2e8fed1, 32'hc3895fd8},
  {32'hc4bceec6, 32'hc2ab7f82, 32'h43953b00},
  {32'h4490aad1, 32'hc3db9e75, 32'hc3b8887b},
  {32'hc425b81e, 32'h431f0b92, 32'h43ced3bd},
  {32'h44d091f3, 32'h43313f2c, 32'hc38f8714},
  {32'hc373ab60, 32'hc34314e1, 32'h426497b6},
  {32'h4528d175, 32'hc259b86f, 32'hc3d0a63e},
  {32'h43c658e6, 32'h43dd23da, 32'hbf98292c},
  {32'h44670d68, 32'hc11e3fc2, 32'hc24dba4a},
  {32'hc3e18340, 32'hc31481a4, 32'h4164b614},
  {32'h4507c2a7, 32'h42136508, 32'h41b33e30},
  {32'hc481dace, 32'h43cabf7d, 32'h42399964},
  {32'h45093170, 32'h43866f18, 32'hc39ea50f},
  {32'hc4e24142, 32'hc3881b74, 32'h4403545b},
  {32'h44cbd42f, 32'hc1df9beb, 32'h436eb9a6},
  {32'hc4be9483, 32'h4328650f, 32'h42e07a36},
  {32'h4467f2cc, 32'h42c9a828, 32'h43967559},
  {32'hc4d3c32e, 32'h434ebdcd, 32'h438ff03a},
  {32'h4471e71a, 32'h4312ff82, 32'h42a7ab16},
  {32'hc4b8d1d2, 32'h4383420f, 32'h43426c8f},
  {32'h44187f88, 32'hc348b9cb, 32'hc3904585},
  {32'hc4ce4ba3, 32'hc21a757b, 32'hc1f30551},
  {32'h42f87950, 32'hc342a1b5, 32'hc39f7f5c},
  {32'hc4afec9a, 32'hc28c5421, 32'hc2ea097e},
  {32'h441dd556, 32'hc3de7317, 32'hc2a10061},
  {32'hc501dcbb, 32'hc3494bd2, 32'hc29271f6},
  {32'h43ab2924, 32'h43b0acdf, 32'h42985d3c},
  {32'hc5122d78, 32'hc2dce347, 32'hc2146dc0},
  {32'h434a678e, 32'hc375f6c0, 32'h42880f39},
  {32'hc42aefd3, 32'h43aed15a, 32'h4391c71e},
  {32'h4516532c, 32'h432e007d, 32'hc366734e},
  {32'hc26d59ec, 32'h40b52f2e, 32'hc3efc40f},
  {32'h442c2360, 32'hc240923f, 32'h4378ba39},
  {32'hc46d4ab8, 32'h42039e84, 32'hc05c0130},
  {32'h445560e8, 32'h431779f2, 32'hc343ea7a},
  {32'hc4cbfc0d, 32'hc2cb27b4, 32'hc1ab726f},
  {32'h44443ffc, 32'h4202e962, 32'hc38e2166},
  {32'hc4a068b7, 32'h43db26c9, 32'h4310b982},
  {32'h44fa3570, 32'h43ae89e5, 32'hc37f91f9},
  {32'hc427ffd0, 32'h41b7dc82, 32'hc35ed404},
  {32'h42728b80, 32'hc35a20eb, 32'h43a6bc1a},
  {32'hc3e6d5d8, 32'h425bed56, 32'h43aca1a5},
  {32'h43b7ebf2, 32'hc2833fb2, 32'h41db7bdc},
  {32'hc41b70c4, 32'h4162065a, 32'h42c68dd6},
  {32'h44a968fa, 32'hc21f2972, 32'h43c86c53},
  {32'hc50b1ad2, 32'hc3194a99, 32'hc20c78c8},
  {32'h448029e0, 32'h438a9c8e, 32'hc33e08f0},
  {32'hc500c1ab, 32'hc2727d98, 32'h4248ae9c},
  {32'h44de596c, 32'h4272505b, 32'h43a88d0a},
  {32'h43ae79a0, 32'h43bd3cd2, 32'hc2e83296},
  {32'h448038aa, 32'hc37768a1, 32'hc401534d},
  {32'h43d2ae90, 32'hc3b245ff, 32'h4101f6dc},
  {32'h4386538a, 32'h42880632, 32'hc4149959},
  {32'hc4ae145e, 32'h42acdde0, 32'hc38c981a},
  {32'hc21a37c0, 32'h43844beb, 32'hc214f27b},
  {32'hc4967888, 32'h440439fd, 32'hc3884d6f},
  {32'h4414132e, 32'h437be3be, 32'h43d4d287},
  {32'hc4dfe58e, 32'hc315bbea, 32'h439ff2ea},
  {32'h442b86b6, 32'h43fd435e, 32'hc32f6995},
  {32'hc4e214e0, 32'h43f04a0a, 32'hc332e796},
  {32'h4487b4f8, 32'hc341e8b0, 32'hc172c240},
  {32'hc4fe49f2, 32'hc3417f79, 32'h42f0d431},
  {32'h4466e609, 32'h415c0d43, 32'hc2cf4570},
  {32'hc49a7f72, 32'hc2de8b68, 32'hc08c56e6},
  {32'h44056036, 32'h4322edfa, 32'h4176bbdf},
  {32'hc4499078, 32'hc3646c6f, 32'hc368a13f},
  {32'h42c40340, 32'hc192f590, 32'h43c53d82},
  {32'hc4883e2f, 32'hc099f9e8, 32'h42d0f89b},
  {32'h44dc459f, 32'hc319daae, 32'h4293f5c1},
  {32'h4217d140, 32'hc315acf7, 32'h4349afbe},
  {32'h44e37424, 32'h41cb3e24, 32'h42be495c},
  {32'hc405e548, 32'hc385010c, 32'h430763ae},
  {32'h43c3da78, 32'h40130008, 32'hc21c2e23},
  {32'hc4b5b824, 32'hc3a3baa6, 32'h4302b15f},
  {32'h44de3808, 32'hc38d625c, 32'hc3a8c37e},
  {32'hc4be6268, 32'h42490198, 32'h4274b127},
  {32'h44f29d3a, 32'hc3c5bff0, 32'hc22bfa48},
  {32'hc42fc07e, 32'h4385ac22, 32'hc201a014},
  {32'hc1ebdf80, 32'hc3286aea, 32'h42fe0f3f},
  {32'hc4e598c1, 32'hc42c67e3, 32'hc331d67f},
  {32'h44e235ce, 32'h4237fe1f, 32'hc3100650},
  {32'hc5080247, 32'hc3544ec1, 32'hc15b99e6},
  {32'h44a93bd0, 32'h43532022, 32'hc21ebc4f},
  {32'hc462f38c, 32'h432dae40, 32'hc0ef881d},
  {32'h44a6d639, 32'h41ca6e8a, 32'hc2eecbae},
  {32'hc317cc90, 32'hc38f0f96, 32'hc25c5f22},
  {32'h449aa218, 32'h438b2dc3, 32'h42db3270},
  {32'hc412523c, 32'hc3503ee0, 32'hc38a539f},
  {32'h445c24f0, 32'hc236f671, 32'h42f3b9a0},
  {32'hc3296dc0, 32'hc2a78598, 32'hc2e2df93},
  {32'h4463f1aa, 32'h43d956d6, 32'h4359d040},
  {32'hc36e21b0, 32'hc35a9f3e, 32'h42d78a30},
  {32'h4491a762, 32'h4315ee68, 32'hc2dbe549},
  {32'hc4b00586, 32'h43c808b7, 32'hc3aa7bb5},
  {32'h4394d688, 32'h41e86f8a, 32'hc22aa8c3},
  {32'hc4c36030, 32'hc1205ffe, 32'hc3d5f182},
  {32'h444c33c6, 32'hc23369ef, 32'hc38e3e99},
  {32'hc4d0a40c, 32'h42d06fb9, 32'h43601bb0},
  {32'h44078787, 32'hc3cc4326, 32'h42e86476},
  {32'hc4bb218d, 32'hc33cab4c, 32'h429cc366},
  {32'h43b8a14a, 32'h43127d64, 32'hc38981d0},
  {32'hc4efab55, 32'h4239b102, 32'h43685a15},
  {32'h450140c0, 32'h3f2c3d60, 32'h439b2215},
  {32'hc4c14a56, 32'h42cbcb21, 32'h42f355db},
  {32'h44bbe8e7, 32'hc24b3a88, 32'hc22e42de},
  {32'hc4295554, 32'h43277a07, 32'h43297043},
  {32'h440927f8, 32'hc21e6c0b, 32'h4304538b},
  {32'hc4cab231, 32'hc374a103, 32'h430151c9},
  {32'h450466cb, 32'h437d0bdd, 32'hc34fc063},
  {32'hc4a25032, 32'hc318019a, 32'hc2b9607a},
  {32'h442cda13, 32'hc3305614, 32'h43f9604b},
  {32'hc4098382, 32'h435e83a5, 32'h42a98f5f},
  {32'h43f4896a, 32'hc1c7c053, 32'hc29bcc0b},
  {32'hc1f9ebc3, 32'hc3551b39, 32'hc2dcfecc},
  {32'h44f95dd4, 32'hc2e58919, 32'hc33aef6c},
  {32'hc4b4b6b8, 32'h43d365e4, 32'h42c3faee},
  {32'h449ab9ce, 32'hc295be2c, 32'h43a80c7d},
  {32'hc4425e0c, 32'hc118e865, 32'hc276192c},
  {32'h442c8e28, 32'h43592602, 32'hc2cf1841},
  {32'hc4859c1a, 32'h43240fa1, 32'hc39e5d89},
  {32'h447a166c, 32'h434b5ace, 32'h4335af32},
  {32'hc50540a4, 32'hc39cd430, 32'h42c6d468},
  {32'h43afaaaa, 32'h43c5f3ef, 32'hc2ead082},
  {32'hc4b2d5eb, 32'hc3469821, 32'hc3117481},
  {32'h43a534ee, 32'h4391ddec, 32'hc255029e},
  {32'hc29144e0, 32'hc3404a34, 32'hc3a51618},
  {32'h4452610c, 32'hc2c90cc7, 32'h4349a152},
  {32'hc277082e, 32'hc287b72f, 32'hc29212d7},
  {32'hc1144dc0, 32'h4388cc42, 32'hc2962694},
  {32'hc4d73f43, 32'h43801d63, 32'h43900a49},
  {32'h4500c852, 32'hc2e2295b, 32'hc2d8c5ad},
  {32'hc5298fb9, 32'hc3b93c03, 32'hc373b86c},
  {32'h450a952c, 32'h437a8e01, 32'hc3917820},
  {32'hc2c54de2, 32'hc205ec20, 32'hc3073b6a},
  {32'h44415400, 32'hc328cd1a, 32'h4374228d},
  {32'hc450ba0e, 32'hc11f3761, 32'h42d055c6},
  {32'h448e2807, 32'hc185400c, 32'h435601e9},
  {32'h425d0154, 32'hc21b52d3, 32'hc32951e8},
  {32'h4373887c, 32'h43016e0b, 32'hc2f6ae54},
  {32'hc4ca4ace, 32'hc37b2948, 32'hc2bba91e},
  {32'h44fba857, 32'hc3a6e417, 32'hc40cbd3e},
  {32'hc4a48de4, 32'h424b1bd0, 32'h441c0281},
  {32'h4517986f, 32'hc2a0b0ed, 32'h43253651},
  {32'hc480e8c8, 32'h425e2c68, 32'hc250619a},
  {32'h45103053, 32'hc3d8b2a3, 32'hc3864ab1},
  {32'hc506cbec, 32'h4288ea1e, 32'h41d6da5a},
  {32'h440d8fec, 32'h439fd2ba, 32'h4316c041},
  {32'hc4f83ca4, 32'h42ff82a4, 32'hc3870470},
  {32'h442fe3ef, 32'hc1c911b9, 32'h438e578d},
  {32'hc4dcd26f, 32'h435b5fe0, 32'hc30cb0d9},
  {32'h44321dac, 32'h43c4e06a, 32'h429dd224},
  {32'hc4977419, 32'h42e5107d, 32'hc3b6b263},
  {32'h450ba613, 32'h42661db9, 32'h43bcd1eb},
  {32'hc3eb80f9, 32'h43892279, 32'hc31d0af6},
  {32'h44b677bd, 32'hc231dd8e, 32'h438478fb},
  {32'hc47afce6, 32'h429df3df, 32'h43283249},
  {32'h44b17d79, 32'h434582fb, 32'hc3920dd5},
  {32'hc4feea1f, 32'h436f6dc6, 32'h4257c986},
  {32'h44a99e41, 32'h4277404b, 32'hc3aacbd8},
  {32'hc4c02cdd, 32'h415e395c, 32'hc2d07f75},
  {32'h44126b04, 32'h41ef233c, 32'hc2bb5112},
  {32'hc348938c, 32'hc2a6e69a, 32'hc35477f7},
  {32'h4222ed98, 32'hc35dd3a8, 32'hc3777527},
  {32'hc4876f18, 32'hc2c1d057, 32'hbff40fb0},
  {32'h448d2733, 32'hc3205bb8, 32'hc29bfa85},
  {32'hc50b601c, 32'h436e282a, 32'hc14b1744},
  {32'h44c2b478, 32'h421361a9, 32'h43990a34},
  {32'hc4f4764e, 32'hc3a94c9c, 32'h42d3643c},
  {32'h44d921a2, 32'hc0d46240, 32'h42a02bf7},
  {32'hc51de6f0, 32'h4323d4f2, 32'h4400a85f},
  {32'h4512e171, 32'h437b24d0, 32'h43a128c9},
  {32'hc28bc973, 32'h4319c846, 32'hc382bd0b},
  {32'h447689dc, 32'h4346f20c, 32'hc30ebd47},
  {32'hc3a8ee44, 32'hc2cc3c46, 32'h43605d8c},
  {32'h44f27232, 32'hc3830ae4, 32'h438dedac},
  {32'hc2e24740, 32'h42da83b3, 32'h41de71ec},
  {32'h4495374c, 32'h43425e40, 32'hc3a4b8f9},
  {32'hc44c3d46, 32'hc3468765, 32'h42463580},
  {32'h44bc5637, 32'h43d0b7ab, 32'hc1d5f07e},
  {32'hc4d00c7c, 32'hc2ec8cfb, 32'hc350507b},
  {32'h44d05d4e, 32'h43f7b791, 32'h440f5e51},
  {32'hc4ccc351, 32'h43873e4f, 32'h433d4384},
  {32'h44a2150a, 32'hc27f5116, 32'hc2d221e4},
  {32'hc4fe4205, 32'h439783ba, 32'h430e882f},
  {32'h44df75e5, 32'h43a0df54, 32'h43892f36},
  {32'hc4dd89c3, 32'hc3ae814d, 32'h4181452f},
  {32'h444e24f2, 32'h42a41bba, 32'h43f932fa},
  {32'hc4f2e202, 32'hc29a3167, 32'h422f5ed9},
  {32'h44898207, 32'hc380edb8, 32'h43c1862d},
  {32'hc4c2378a, 32'h43b08fde, 32'h434024f3},
  {32'h44fc04e5, 32'hc3d72812, 32'hc34f1119},
  {32'hc10ff200, 32'hc350d9c0, 32'hc265057d},
  {32'h440f5afe, 32'h43d64bbf, 32'hc0f42d0f},
  {32'hc41d1646, 32'h4392bf99, 32'h415eceda},
  {32'h448aabfe, 32'h437f4cf2, 32'hc340e140},
  {32'hc4d3706a, 32'hc35cbe61, 32'h423969b9},
  {32'h4352a773, 32'hc1eb0c84, 32'h43a841e7},
  {32'hc4f86d02, 32'hbfd0d378, 32'h42a5e37b},
  {32'h44b9753a, 32'h43330959, 32'hc26a9bcc},
  {32'hc4820374, 32'hc1c86444, 32'h4382c68f},
  {32'h44a40372, 32'h42c77faa, 32'hc37444e9},
  {32'hc4e9455f, 32'hc249624c, 32'h42cb65c4},
  {32'h4501c9a8, 32'h43e707ff, 32'h436bc4b7},
  {32'hc441fb54, 32'h43219a12, 32'hc226e606},
  {32'h45071e2a, 32'h43731050, 32'hc361a024},
  {32'hc517863c, 32'h4314cb43, 32'hc3700c5e},
  {32'h44e13c92, 32'hc2951378, 32'hc36082b7},
  {32'hc3a2769c, 32'hc37ffc8e, 32'hc2a78661},
  {32'h44901724, 32'h42811f45, 32'hc2733bd4},
  {32'hc410fe43, 32'h41b5a0cc, 32'hc2ac7aa7},
  {32'h443834bc, 32'hc389116b, 32'h4280ddd4},
  {32'hc4727c8a, 32'h4288d90e, 32'hc3582db7},
  {32'h43ec97d8, 32'hc289e870, 32'h428a7a6b},
  {32'hc3e267c0, 32'hc2b6abf4, 32'hc2c8cf55},
  {32'h44453494, 32'h4390dc5d, 32'hc36a004d},
  {32'hc41c4714, 32'h43b75834, 32'h4133d5e3},
  {32'h4431c270, 32'h42d4f5a3, 32'hc2f19ddd},
  {32'hc4a7f588, 32'h43023ba7, 32'hc29db7c8},
  {32'h44ae6e71, 32'h42e5bcfd, 32'h42cf26e7},
  {32'hc40dd147, 32'h43648ea8, 32'hc339ca60},
  {32'h452d4ee1, 32'hc2f4fe30, 32'h412d99a4},
  {32'hc5013cc6, 32'hc29ec1f5, 32'h439d917a},
  {32'h451f7768, 32'h40d901f0, 32'hc39222d2},
  {32'hc4b3e524, 32'hc2244427, 32'h44029990},
  {32'h44a8e478, 32'h42c9d73c, 32'h429b896b},
  {32'hc50c36a7, 32'hc30a5118, 32'hc39b4e62},
  {32'h44fd8b78, 32'hc27e12ce, 32'h426aa36c},
  {32'hc433736c, 32'h42af2fc3, 32'hc2cfab36},
  {32'h435604e8, 32'h43bb2fe3, 32'h437253c0},
  {32'hc41a2e57, 32'h43896eba, 32'hc110bfc2},
  {32'h4502be1a, 32'hc3085e94, 32'h4135d712},
  {32'hc453f3b3, 32'hc3fec50f, 32'h41b64c09},
  {32'h42f68310, 32'h439caca4, 32'hc354d02d},
  {32'hc4712bf8, 32'hc3b44003, 32'hc3817dec},
  {32'h43a7a4fd, 32'h439ad0a8, 32'h43430b96},
  {32'hc4a96842, 32'hc280bc68, 32'h43a53307},
  {32'h45010b3c, 32'hc22e6e60, 32'hc31d8f6a},
  {32'hc50228d4, 32'hc3941e92, 32'h43a48813},
  {32'h4509f928, 32'h435106e2, 32'hc3134407},
  {32'hc4de9e9e, 32'h4337ebe6, 32'hc36c3ec0},
  {32'h44359981, 32'h42d742f8, 32'hc0b4f0cc},
  {32'hc47689e9, 32'hc2b213ed, 32'h4339f296},
  {32'h448aa34a, 32'hc3479540, 32'h427c326e},
  {32'hc4821b0a, 32'h43399c7e, 32'h4312b8d4},
  {32'h44eccf50, 32'h428e9bb9, 32'h42bb0034},
  {32'hc4de077c, 32'h42b93ed7, 32'h42a8d2ac},
  {32'h44caf60a, 32'h43406c4f, 32'hc2cf3e58},
  {32'hc45279de, 32'hc2ed407e, 32'hc3453770},
  {32'h448a1b71, 32'h4392bda3, 32'h43c47155},
  {32'hc4127880, 32'h436cecef, 32'h43da8df8},
  {32'h44cac01e, 32'hc1918453, 32'h42a47579},
  {32'hc51c2151, 32'hc27a6ea6, 32'hc2b4a264},
  {32'h45115147, 32'h43b1be76, 32'h437f25b0},
  {32'hc4c693be, 32'h4422f492, 32'h432fb5f9},
  {32'h4469730d, 32'h435908cf, 32'h423436a1},
  {32'hc4f27983, 32'h4294e216, 32'h439a493b},
  {32'h45056ac0, 32'h41ce1752, 32'h42de4def},
  {32'hc4dd4ac7, 32'h433d6897, 32'hc2512de6},
  {32'h44b7532b, 32'h4314100a, 32'hc17ffabc},
  {32'hc4fb7a36, 32'h43a07cd7, 32'h4337e77e},
  {32'h44997772, 32'h43e0c658, 32'hc28a4e7f},
  {32'hc27aecf0, 32'h43177b27, 32'h42f83052},
  {32'h44112087, 32'hc2e7acb0, 32'hc310f063},
  {32'hc4290d96, 32'h42af537f, 32'hc387b5d3},
  {32'h44fca3a7, 32'hc2dcccd5, 32'hc3b2ac7c},
  {32'hc4d04b5f, 32'hc2b341c8, 32'hc393cfbc},
  {32'h44fd92ec, 32'hc19c397c, 32'hc3a8310d},
  {32'h428875f5, 32'hc2803e68, 32'hc28e65b4},
  {32'h43e83677, 32'hc23347d9, 32'h42d2b66c},
  {32'hc35fbbae, 32'h43392472, 32'hc34d0af6},
  {32'h4381722c, 32'hc0a72197, 32'hc36f55ba},
  {32'hc503565e, 32'h43734532, 32'hc3dcae61},
  {32'h4440cec9, 32'hc28dbf00, 32'hc3e8bc80},
  {32'hc4295d3c, 32'hc23fe8d2, 32'hc1d61c9b},
  {32'h44e0c87a, 32'hc2d764c7, 32'h41f54386},
  {32'hc4a1955b, 32'hc344c3ec, 32'h43ec7dde},
  {32'h43f188d8, 32'h42f1d2a9, 32'hc30c3525},
  {32'hc4b1b83d, 32'hc1bbdf1b, 32'h4310c8f5},
  {32'h447bec89, 32'h43ea6e54, 32'hc36d6975},
  {32'hc4a8732c, 32'h43864054, 32'h444195cb},
  {32'h43fd9a53, 32'h4380a069, 32'hc3dd73b2},
  {32'hc46cc484, 32'hc1b6b719, 32'h438a59a4},
  {32'h448a9af7, 32'h43a6eb14, 32'hc3cc19c0},
  {32'hc449ab94, 32'h43e142ba, 32'hc255ade8},
  {32'h4518ad88, 32'hc3337661, 32'hc169fd94},
  {32'h421a78e2, 32'hc20e6aeb, 32'h43d3c733},
  {32'h44e3993c, 32'hc220157b, 32'h424bdea2},
  {32'hc484aff3, 32'hc3e46d10, 32'h43443d8e},
  {32'h4302ea34, 32'h42e13af9, 32'h43537819},
  {32'hc4ac0e60, 32'hc2b4ee32, 32'h4296250f},
  {32'h43dc50b8, 32'h43472a67, 32'hc30623e1},
  {32'hc4ecba80, 32'hc2343234, 32'h426f1c57},
  {32'h44f6a978, 32'h424013d8, 32'h43d0827c},
  {32'hc44c30e4, 32'h433827b7, 32'h42de8f30},
  {32'h449756c3, 32'hc3100d68, 32'hc3bb4564},
  {32'hc51a57f0, 32'h43906f05, 32'h430a6023},
  {32'h44a9c51a, 32'hc2a4c8ca, 32'h43109c63},
  {32'hc4ed289c, 32'hc36ed63c, 32'hc34b1cf7},
  {32'h44c87854, 32'h42855d3b, 32'h41fdc337},
  {32'hc4dcda70, 32'h43006f99, 32'h42968667},
  {32'h44cbce4a, 32'hc383fac2, 32'hc325e74e},
  {32'hc484c4fb, 32'hc3e4a5b7, 32'h429c6cfd},
  {32'h44ca5615, 32'hc30e9d19, 32'hc347bebe},
  {32'h44d7d966, 32'hc3bb03dc, 32'h43441b02},
  {32'hc5086698, 32'hc41559a0, 32'h4307bc5e},
  {32'h44d291d1, 32'hc30d1e5a, 32'h43c00716},
  {32'hc486cb0d, 32'h43a16345, 32'hc301e174},
  {32'h4427ec46, 32'hc31086ab, 32'hc275e8e1},
  {32'hc457d640, 32'hc378af2d, 32'hc38d66b2},
  {32'h44c57444, 32'hc2a89e3c, 32'hc3563ede},
  {32'hc3faeb29, 32'h439718b0, 32'h434d9ce1},
  {32'h44d35ef5, 32'hc2a750a6, 32'h43ac4d2e},
  {32'hc4a31299, 32'h43bf6d88, 32'hc3db0f6b},
  {32'h439e9d98, 32'h41748ee0, 32'hc35a395a},
  {32'hc4969886, 32'h430d88d9, 32'hc333ba4f},
  {32'h44864cf6, 32'h43d88c99, 32'hc35e5431},
  {32'hc4676556, 32'h425cd59a, 32'hc33c2060},
  {32'h44b6c512, 32'hc3823ae8, 32'hc28032d9},
  {32'hc3b19884, 32'h438754e6, 32'hc3410a93},
  {32'h44ca074a, 32'h43aa3461, 32'h4383b0d6},
  {32'hc4b18ab1, 32'hc2f883cc, 32'h428d5801},
  {32'h44b46ed5, 32'h43ef7cda, 32'h43598387},
  {32'hc408d62c, 32'h4262ef6a, 32'h427f0046},
  {32'h445e39b2, 32'hc39ae985, 32'hc3b00c7f},
  {32'hc528481f, 32'h43f8b800, 32'hc2f7d781},
  {32'h43ea63f0, 32'hc3bb5286, 32'hc34c1101},
  {32'hc440ec88, 32'h4354401c, 32'h428799f2},
  {32'h441feaa0, 32'h42bdbd6a, 32'hc3946f92},
  {32'hc3fae99c, 32'hc3e1b3ba, 32'h43a5daa9},
  {32'h44337832, 32'h42a32b33, 32'hc23ce3eb},
  {32'hc3ca1a50, 32'h434342e1, 32'h421ca79e},
  {32'h43ba65cc, 32'hc369256e, 32'hc3c5883e},
  {32'hc47ab17a, 32'h433ff72e, 32'h429f82c9},
  {32'h44af72c7, 32'hc2f68f23, 32'h414fd553},
  {32'hc3ca6278, 32'hc3800a34, 32'h416c04ea},
  {32'h433703c8, 32'hc3a7239d, 32'h429d62fa},
  {32'hc48f3764, 32'hc36c9610, 32'h43373b50},
  {32'h449c12be, 32'hc38753d2, 32'h42b3ca6c},
  {32'hc456e903, 32'h41f6e419, 32'h42aa6732},
  {32'h4401cac2, 32'hc31a4f22, 32'hc2bae407},
  {32'hc4571e6d, 32'h439ae61f, 32'hc4088860},
  {32'h44a17325, 32'hc4035d2a, 32'h437c7fdc},
  {32'hc50128b5, 32'hc1bfedb2, 32'hc2f95453},
  {32'h44c6916f, 32'hc34259c2, 32'hc3620c01},
  {32'hc41f2ba6, 32'h43912ff9, 32'hc1804d66},
  {32'h44a39234, 32'hc2add2ea, 32'h41b39fda},
  {32'hc50ee07b, 32'hc34c3ad9, 32'h42e5c925},
  {32'h44dbc556, 32'hc28d0640, 32'h432c474e},
  {32'hc522dab1, 32'hc3d2cb1b, 32'h436fe976},
  {32'h4403d9e4, 32'h42ae83a8, 32'hc1ccc6a4},
  {32'hc5107265, 32'h430c5095, 32'h42a08a8f},
  {32'h447e4548, 32'h414ba92c, 32'h43895d14},
  {32'hc4248d70, 32'h42b5bc11, 32'h43135d9a},
  {32'h44f89e64, 32'h43510518, 32'h43d3edd9},
  {32'hc4a64271, 32'hc2aadcaa, 32'h43be54de},
  {32'h449d14ae, 32'h41db65af, 32'h42933155},
  {32'hc49519ea, 32'hc35791d3, 32'h4337a218},
  {32'h44b4b9c4, 32'h439b2d54, 32'h43080ad3},
  {32'hc4ba6277, 32'hc308f20e, 32'hc30f9db4},
  {32'h44ed9260, 32'hc22728a1, 32'hc2e2cf35},
  {32'hc4e363a7, 32'h439d0351, 32'hc44c1273},
  {32'h447b2840, 32'h437b56ac, 32'hc3bb1535},
  {32'hc3d963c8, 32'h42ba1b3d, 32'h42b881c6},
  {32'h44e1f3d7, 32'hc3c8c0e6, 32'h435904f3},
  {32'hc50ed3a0, 32'h42a3d526, 32'hc2a807ce},
  {32'h4460e406, 32'hc3b79abf, 32'hc38dcee1},
  {32'hc4f99e48, 32'hc36fc9f8, 32'h42a70538},
  {32'h44a01400, 32'h41a8be94, 32'h431a9da2},
  {32'hc49df109, 32'h43f04b47, 32'h41a67a80},
  {32'h450d5a68, 32'h41e7a3bf, 32'h423efbd4},
  {32'hc50230a7, 32'hc2c5a074, 32'hc30d994c},
  {32'h4421ac7f, 32'hc35b0a94, 32'hc26e9d5a},
  {32'hc3a73ee7, 32'h43243e8b, 32'hc303f82b},
  {32'h44b08782, 32'h41eccd19, 32'h41be22f2},
  {32'hc500f34b, 32'hc35f3542, 32'hc027a980},
  {32'h44bb2428, 32'h43836769, 32'hc3a5b5f1},
  {32'hc2b1d39f, 32'h429595e9, 32'hc31021ec},
  {32'h44339146, 32'h42991903, 32'h43a975b9},
  {32'hc5083e1e, 32'h43a50a1f, 32'hc3ce355a},
  {32'h44aaec7f, 32'h42ae28f5, 32'hc37b1692},
  {32'hc48a5dac, 32'hc2cbe411, 32'h434d6036},
  {32'h448c9266, 32'hc1ee52ff, 32'hc393dba3},
  {32'hc418c22a, 32'hc1c326cc, 32'h42a45237},
  {32'h4501e648, 32'hc3d83f19, 32'hc1d30827},
  {32'hc4f6de0d, 32'hc35cc306, 32'hc33770d2},
  {32'h44994d7d, 32'hc3a719c6, 32'hc3e75475},
  {32'hc4af0138, 32'h42b474c4, 32'hc379ee34},
  {32'h4491cf7c, 32'h422ec8db, 32'h4218d0d1},
  {32'hc39fb93e, 32'h42c364c5, 32'h4319b91b},
  {32'h44764823, 32'h4393700e, 32'hc2d97b78},
  {32'hc4d398ca, 32'hc399d870, 32'hc251fa1d},
  {32'h438f600c, 32'h4312d9ec, 32'hc210a016},
  {32'hc49f1f1c, 32'hc3d01c56, 32'hc251f86b},
  {32'h43f93e8d, 32'h41db7749, 32'hc38cc2d5},
  {32'hc4833c3a, 32'hc2dd2e3e, 32'h428323f8},
  {32'h4464a948, 32'hc06e19f0, 32'hc1daf9e2},
  {32'hc5054444, 32'hc32db514, 32'hc2f9abdf},
  {32'h449d39fa, 32'hc2477bcc, 32'h43432f96},
  {32'hc4f0b397, 32'hc30368a4, 32'h42cb9c19},
  {32'h442c1fe9, 32'hc3d01dc5, 32'hc3278eb8},
  {32'hc4f16453, 32'h4331f4a9, 32'hc2f9b9ec},
  {32'h4501e0c2, 32'hc386878f, 32'hc1b30786},
  {32'hc45ea988, 32'h43da3062, 32'h43036bb1},
  {32'h430fc7bc, 32'h43943bae, 32'h432192cb},
  {32'hc50290a8, 32'h43cb8802, 32'h43912d15},
  {32'h451264b0, 32'hc29a5128, 32'h42bf8145},
  {32'h42bcfd00, 32'hc39def45, 32'h4356c37b},
  {32'h4508742c, 32'h425ac1c0, 32'hc3a5c3b5},
  {32'hc4aea553, 32'h4335c5ee, 32'h42f797b2},
  {32'h451857a3, 32'h42a5cb07, 32'hc245f681},
  {32'hc41279c6, 32'h42f4dada, 32'h42d57aa2},
  {32'h446d0130, 32'hc397589d, 32'hc1b92fc4},
  {32'hc4a1af14, 32'h42d537ac, 32'h4315426e},
  {32'h450ea6b4, 32'h42f92d93, 32'hc34f104f},
  {32'hc36355af, 32'hc37be64b, 32'h42cf9da8},
  {32'h41a77a80, 32'h41a9223d, 32'h432da48b},
  {32'hc4e96bb0, 32'hc3820f8d, 32'hc29468e9},
  {32'h43c3c74c, 32'h43d8ad12, 32'h42e17e7b},
  {32'hc50fecdb, 32'hc33dc8df, 32'hc38cf8dc},
  {32'h45069e02, 32'h422c13eb, 32'hc1ec3b4a},
  {32'hc519c6dc, 32'h43554cdb, 32'hc2a81d8a},
  {32'h4508f4f3, 32'h43049ce5, 32'hc2c07346},
  {32'hc4a98772, 32'h41c1bf56, 32'h437dab86},
  {32'h444eb20e, 32'h43759cd7, 32'h43aea791},
  {32'hc51590e4, 32'hc1cd807e, 32'h438f6aa8},
  {32'h41d1b080, 32'hc1c3fb70, 32'h432ebd40},
  {32'hc407c687, 32'h42b44bcb, 32'hc07486b5},
  {32'h448805a8, 32'hc25fbe42, 32'h42505270},
  {32'h3f905800, 32'h42414d7d, 32'h427a8a29},
  {32'h450166d0, 32'hc3206e3c, 32'h42a1c994},
  {32'hc4ad1902, 32'h4318e438, 32'h436dcb5f},
  {32'h451f2d3d, 32'hc26187ac, 32'h4332ff0c},
  {32'hc4fb7be3, 32'hc301d371, 32'hc1c0758e},
  {32'h44ef50a0, 32'h41f0abbc, 32'h433a04f6},
  {32'hc50caf15, 32'h433dd230, 32'h420864d4},
  {32'h4315d030, 32'h44040af8, 32'hc34db3f5},
  {32'hc48811a5, 32'hc33f5681, 32'hc2db6ee7},
  {32'h44b817e8, 32'hc0355a9e, 32'h43d68cc5},
  {32'hc423903c, 32'hc2b91029, 32'h4228cf31},
  {32'h43ce83f8, 32'h42b0440c, 32'h432b7e8c},
  {32'hc2dfac20, 32'h4395d6a4, 32'hc3eb11ec},
  {32'h4504484d, 32'hc366ae3e, 32'h3f9da350},
  {32'hc46c99f4, 32'h433eba57, 32'hc372aa43},
  {32'h4463f442, 32'h426203e2, 32'h42fe7eb3},
  {32'h4317fa70, 32'hc0cb45c3, 32'h4352d8e4},
  {32'h442f910e, 32'hc3bf7393, 32'h43045cca},
  {32'hc23cc880, 32'hc3b9ba15, 32'h4344aebf},
  {32'h44eb8db1, 32'hc356432c, 32'h43d9a2d6},
  {32'hc335db04, 32'h41ba6a38, 32'hc306a91f},
  {32'h44a70d2c, 32'h43cb7558, 32'h4103c55d},
  {32'hc1f82edb, 32'h43fb8594, 32'h4369be6d},
  {32'h446d226a, 32'hc2e3c83b, 32'h4305375e},
  {32'hc34a650a, 32'h43932e91, 32'hc23e79a5},
  {32'h44f5f488, 32'h435ace8c, 32'h4352ce81},
  {32'hc4902ddb, 32'hc37e916c, 32'hc282be77},
  {32'h4421a839, 32'hc393b457, 32'hc28d4a82},
  {32'hc48cb39c, 32'hbf06cdc8, 32'hc3992b6a},
  {32'h4481e3b8, 32'h42da30a6, 32'hc305b690},
  {32'hc45458d4, 32'hc2cb282c, 32'h434bff65},
  {32'h44b6745c, 32'h43307472, 32'hc189eb8a},
  {32'hc4a3efe5, 32'hc394a472, 32'hc3567131},
  {32'h44d7fedc, 32'hc31b6770, 32'hc2aeeda5},
  {32'hc4690e33, 32'h43b2f309, 32'h43a71035},
  {32'h44f2d2cd, 32'hc1f5f68c, 32'hc3471662},
  {32'h421d2900, 32'hc39c7d24, 32'h4313766c},
  {32'h4441ba31, 32'hc329d467, 32'h43e0beee},
  {32'hc4b0d9fe, 32'hc270b609, 32'hc318a802},
  {32'h44e4bc6d, 32'hc3a5cd3f, 32'hc1609b3d},
  {32'hc463edb0, 32'h42e06a49, 32'hc30c6f46},
  {32'h44ed883e, 32'h42e5c26c, 32'hc2e3d162},
  {32'h42a28a60, 32'h42a0afb2, 32'h42f784a4},
  {32'h44838ff3, 32'hc2b40a58, 32'hc2bad00b},
  {32'hc4e61bee, 32'h429fa580, 32'hc2f73a76},
  {32'h44b91ef0, 32'hc3135d74, 32'hc210d9ef},
  {32'hc50629ec, 32'hc3a84690, 32'hc2ab6101},
  {32'h4351b6e9, 32'hc3aad3ac, 32'hc2c3bc14},
  {32'hc4dd566e, 32'h4392bbfd, 32'hc30a2d32},
  {32'h4511f31e, 32'h430c7dc7, 32'h42f7c7ed},
  {32'hc4b558c4, 32'hc28a6ddd, 32'hc302093c},
  {32'h44b7f52f, 32'hc1518a66, 32'hc1fadfb6},
  {32'hc461f531, 32'hc35d930f, 32'h438ba1b6},
  {32'h44801935, 32'hc3a222be, 32'h436b1d02},
  {32'hc386ffd8, 32'h438a4948, 32'hc3fbd7bc},
  {32'h44d08376, 32'h41604250, 32'h4268b413},
  {32'hc45369d7, 32'hc23b7e08, 32'hc3a30e1a},
  {32'h44049338, 32'h4292a514, 32'h41a8c7c9},
  {32'hc407f9ca, 32'h43d7074b, 32'hc37d2e53},
  {32'h4453d100, 32'hc30373d6, 32'h42cb70cd},
  {32'hc3a37db8, 32'hc290534b, 32'h4323d8e1},
  {32'h44b7e88b, 32'h42917c56, 32'hc3e0c80b},
  {32'hc4156900, 32'h43d23db6, 32'hc240527a},
  {32'h4502263e, 32'hc3300d2b, 32'h421db603},
  {32'hc36b4aa8, 32'h41c63096, 32'hc33f0123},
  {32'h428ecdf0, 32'h4319ccac, 32'hc2ccace8},
  {32'hc50dfd42, 32'h4322c25f, 32'hc2eeafef},
  {32'h450bcd6c, 32'h42f3d27f, 32'hc355f4d9},
  {32'hc39e181c, 32'hc33ed2b0, 32'h4308f57a},
  {32'h44ea1beb, 32'h429a7ff1, 32'h4396f8e4},
  {32'hc4f27942, 32'hc379a749, 32'hc054ca65},
  {32'h44c5aa25, 32'h42e6415e, 32'h419a4fdc},
  {32'hc505bd20, 32'hc3f48cad, 32'h4304b735},
  {32'h44779205, 32'hc2daa1c0, 32'hc22ddc63},
  {32'hc497962a, 32'hc28e0169, 32'h43eded4f},
  {32'h44cfe233, 32'hc31d0d26, 32'h43b1eed0},
  {32'hc5076a88, 32'hc3bcc2de, 32'h43ad10d6},
  {32'h447a8760, 32'h413eb9b1, 32'h431a61ae},
  {32'hc4513c4e, 32'h4220b6bc, 32'hc1197e84},
  {32'h44b6650e, 32'hc46413ff, 32'h43eda14e},
  {32'hc4a2a365, 32'h42385f75, 32'h434ff89d},
  {32'h449089c5, 32'hc3b3187d, 32'h43ad871c},
  {32'hc48cda57, 32'h428b3bce, 32'hc401ac4e},
  {32'h45191c94, 32'hc32748b5, 32'hc3ba2168},
  {32'hc30e2310, 32'h418299cb, 32'hc103bba2},
  {32'h44b49fb9, 32'hc0b85f61, 32'hc3b6288f},
  {32'hc4d39271, 32'h432e18ef, 32'h428e8dd2},
  {32'h450aff18, 32'h42bc2618, 32'h42cf98de},
  {32'hc4e848d4, 32'hc2345a3e, 32'h4315f898},
  {32'h44694825, 32'h43040334, 32'hc25b3c4f},
  {32'hc43c2cf5, 32'h431c1f97, 32'hc3059fd6},
  {32'h446759a2, 32'h42e540c8, 32'hc351a891},
  {32'hc393cc38, 32'hc16ce9ea, 32'h428af1bf},
  {32'h4444e232, 32'h42232fdc, 32'h44044208},
  {32'h4311c718, 32'h43d6ace5, 32'h43a11657},
  {32'h43aa97ee, 32'h4309b7f1, 32'h43cc97c0},
  {32'hc5137d7d, 32'hc19719e5, 32'hc37677ad},
  {32'h44c86a68, 32'hc390a27a, 32'hc29d8545},
  {32'hc2e7cce0, 32'h438b99d7, 32'h430d4928},
  {32'h4512067f, 32'h43cae73b, 32'h424073c6},
  {32'hc385f028, 32'h4200b8d4, 32'h42c96a4e},
  {32'h44a77aba, 32'h40f246e1, 32'h42b93044},
  {32'hc2ed4af0, 32'hc30c48f4, 32'hc39ce7c6},
  {32'h43bad1fc, 32'hc2dac0b7, 32'h423fa327},
  {32'h43294de0, 32'h43b69475, 32'hc397d30a},
  {32'h442501bb, 32'hc29c0139, 32'hc289b913},
  {32'hc42e466b, 32'h43e7c890, 32'hc2393ac2},
  {32'h447f5882, 32'h4211e09d, 32'h43864167},
  {32'hc44a6cb1, 32'hc36890d4, 32'hc1a0efeb},
  {32'h44be2cd5, 32'h4387a761, 32'hc3939eec},
  {32'hc4af6a04, 32'hc38b494b, 32'hc3faa4fe},
  {32'h451d5e68, 32'h43458091, 32'hc31f4a5d},
  {32'hc5068dff, 32'hc3bde1df, 32'hc34d1d71},
  {32'h44165dba, 32'hc2cd31b1, 32'h40ee2f84},
  {32'hc4a0de70, 32'hc03f32af, 32'hc1225bd9},
  {32'h44414fb0, 32'h40d5f5a4, 32'hc32de4af},
  {32'hc4907dac, 32'h437afcb1, 32'h42b56531},
  {32'h4514e7ef, 32'hc32738b3, 32'hc278ff1e},
  {32'hc47572fb, 32'h422518d0, 32'hc28272e6},
  {32'h4500d110, 32'h4354a191, 32'hc297ffac},
  {32'hc4ad77bc, 32'hc2f89790, 32'h435f4b11},
  {32'h4478f5f5, 32'h4068e072, 32'hc36a0029},
  {32'hc3a630a1, 32'h4287ce56, 32'h40a93a8e},
  {32'h44c88225, 32'h433e93d1, 32'hc23923b7},
  {32'hc4df16c4, 32'hc288bdea, 32'hc368328d},
  {32'h4497389d, 32'h42dc9be0, 32'h42a2363c},
  {32'hc41c8a74, 32'hc324bc80, 32'h43a5db99},
  {32'h43b476e8, 32'hc2ee205a, 32'hc21be612},
  {32'hc4d5b344, 32'h421c2af2, 32'h43848d02},
  {32'h438d9504, 32'h433d2873, 32'h43463873},
  {32'hc4c25d2f, 32'hc3870dbd, 32'h43125a71},
  {32'h44d78093, 32'h422db25a, 32'hc305db30},
  {32'hc413ca18, 32'h4160b740, 32'h4326ea36},
  {32'h44436540, 32'hc397076b, 32'h42b800b8},
  {32'hc49e43cf, 32'hc3501b14, 32'h43666117},
  {32'h44b883c5, 32'h43ef3284, 32'h43365e74},
  {32'hc4cbc3fc, 32'h427ba090, 32'hc2159a67},
  {32'h448c0a58, 32'h43c07086, 32'hc31bb016},
  {32'hc510a3e5, 32'hc32d6279, 32'h435517bf},
  {32'h44609734, 32'h43bf2866, 32'hc421c1c2},
  {32'hc4c685a1, 32'hc3264575, 32'h428127fd},
  {32'h443a4218, 32'hc23b901d, 32'hc4043125},
  {32'hc3f18338, 32'h44194b7b, 32'hc158bf88},
  {32'h44b01c02, 32'hc31bdb7b, 32'hc39f8098},
  {32'hc39466c0, 32'h4235a8ba, 32'hc3144608},
  {32'h43a78ac0, 32'h430252ce, 32'h4376f740},
  {32'hc395f598, 32'h430a43e4, 32'h437c9dde},
  {32'h449a40d0, 32'h430649aa, 32'hc2ced7e4},
  {32'hc3c4da94, 32'h438b32ac, 32'h42823eae},
  {32'h441ab1f8, 32'hc297ae92, 32'hc32230d5},
  {32'hc41160f4, 32'hc363f768, 32'h41eff88a},
  {32'h4517e8b5, 32'h419888b9, 32'hc3275e9d},
  {32'hc3ee5a9e, 32'hc2ab4710, 32'hc316d011},
  {32'h4418f302, 32'h4329643d, 32'hc33e427d},
  {32'hc487e2a2, 32'h4345b563, 32'h41cfe683},
  {32'h4310f420, 32'h439b2a43, 32'hc189d3db},
  {32'hc49f55c5, 32'hc3119a0f, 32'hc2c3eae0},
  {32'h438fae3e, 32'h431ecedc, 32'h42e5cbad},
  {32'hc36e8c40, 32'hc2554523, 32'h42d58090},
  {32'h44a9e7a1, 32'h434ea6ba, 32'h425be551},
  {32'hc31171a3, 32'h42d5a978, 32'h435f92b3},
  {32'h4479989c, 32'h424a7d89, 32'hc1b9cef5},
  {32'hc3948cf8, 32'hc2d723e8, 32'h3f1e6aa0},
  {32'h44935af6, 32'hc3d016d2, 32'hc23029fc},
  {32'hc4d1c938, 32'h42ed7c35, 32'hc239c71d},
  {32'h447997e7, 32'hc3f7846c, 32'hc3273727},
  {32'hc47b62df, 32'hc33ed845, 32'h43747106},
  {32'h43c103c8, 32'hc32e84de, 32'h41011d6d},
  {32'hc508c9d1, 32'h433766d4, 32'hc32b045d},
  {32'h44d43031, 32'hc2e22732, 32'h42a0eb04},
  {32'hc4ab7ee0, 32'hc1f6e2d0, 32'hc2453390},
  {32'h45156d67, 32'hc329708d, 32'h42f14a9d},
  {32'hc4b3508b, 32'h4249c621, 32'h43868a21},
  {32'h450f910b, 32'h4141f98e, 32'h4264208e},
  {32'hc3f1bee8, 32'hc2dc18b5, 32'h3ecfa118},
  {32'h43a613a8, 32'hc30a9342, 32'hc348835d},
  {32'hc2d40178, 32'h4398c5d0, 32'hc3426092},
  {32'h44190a64, 32'hc30f731e, 32'hc336bc2c},
  {32'hc4feecda, 32'h42becd92, 32'h439d9f79},
  {32'h45043424, 32'h431ea9f4, 32'hc2d53efe},
  {32'hc50f9815, 32'hc31fbae2, 32'hc408db56},
  {32'h44fe3844, 32'hc35302e7, 32'hc2b65554},
  {32'hc4984484, 32'hc3a16c36, 32'h434dc19b},
  {32'h441aac7c, 32'h42db37dd, 32'hc2ec573c},
  {32'hc4bd54d9, 32'h439ee190, 32'h432a8b4c},
  {32'h44906075, 32'h42cf8f82, 32'hc3f586e3},
  {32'hc5025c04, 32'hc2b01978, 32'h4277e5a2},
  {32'h42827f20, 32'hc32b6945, 32'h434ac58e},
  {32'hc4cfce95, 32'hc2d8e702, 32'hc267746b},
  {32'h44c0c681, 32'hc390b740, 32'h439a3e1b},
  {32'hc4f10e2f, 32'h4395b2e6, 32'hc2f1dabf},
  {32'h450f4283, 32'hc2dd9a40, 32'hc361e0a3},
  {32'hc4704706, 32'h435023fe, 32'hc2de960a},
  {32'h44a9f5a4, 32'h42fd57c9, 32'hc2876b79},
  {32'hc48cb9d7, 32'hc25e4f6d, 32'hc30beed4},
  {32'h44832ae8, 32'h421df596, 32'hc33ece6d},
  {32'hc3c4f9c0, 32'hc2a128d7, 32'h43842457},
  {32'h4382acd8, 32'h4330163c, 32'hc2b2b7c1},
  {32'hc4f5a983, 32'h42650733, 32'h43ab0dc2},
  {32'h44dfb55a, 32'h4267753f, 32'h43bdc617},
  {32'hc46b6b18, 32'hc3226e0c, 32'h4303232b},
  {32'h447f41ee, 32'hc2a3ea9e, 32'hc2376506},
  {32'hc50690f9, 32'hc1706853, 32'hc30fe96c},
  {32'h4505f08c, 32'hc30a7e89, 32'hc34e3dc9},
  {32'hc47dddfa, 32'h43adc83d, 32'hc3286b6a},
  {32'h4446fbf9, 32'hc2bc4005, 32'hc38c3515},
  {32'hc4ba99df, 32'h42c08309, 32'h42d3d0f2},
  {32'h444ad6bc, 32'h432a67d4, 32'h4304ab22},
  {32'h414ca000, 32'hc31517ce, 32'h421b6adc},
  {32'h43c6984e, 32'hc080370d, 32'h4354eb2f},
  {32'hc514f400, 32'h411e6478, 32'h4317b0b9},
  {32'h45175a97, 32'h43911689, 32'hc311c186},
  {32'hc3d9f300, 32'h43992fed, 32'hc35268a0},
  {32'h43a971f8, 32'h4349be43, 32'hc16eee70},
  {32'hc4dd6f6f, 32'h41f08d21, 32'h42d50e2b},
  {32'h43e631d0, 32'h42a55094, 32'hc30b77ab},
  {32'hc510463c, 32'h43a7952c, 32'hc2d9bb33},
  {32'h451bf5aa, 32'h4376e946, 32'hc3ca8991},
  {32'hc2973f60, 32'hc40612c9, 32'h43508504},
  {32'h4448d29c, 32'h432c8c65, 32'h42947b47},
  {32'hc44006ab, 32'h424e4ad3, 32'hc2beb4d8},
  {32'h43ca0ee4, 32'h43510899, 32'h43a6bdb6},
  {32'hc4918f95, 32'hc2e8f05a, 32'h4229b899},
  {32'hc2ee9c98, 32'h439227fd, 32'hc3de7a8a},
  {32'hc4914f08, 32'hc33516bf, 32'hc0bb22cb},
  {32'h448aef62, 32'hc23ebfd7, 32'h42c6d487},
  {32'hc4ad4e2b, 32'hc345dac7, 32'h41c83bc8},
  {32'h43ea117c, 32'hc20651b7, 32'hc31479c4},
  {32'hc3a37948, 32'hc337df08, 32'h4350f33d},
  {32'h4463d1cb, 32'h43bd2366, 32'h413d7b34},
  {32'hc4d3eb1f, 32'h4279fd78, 32'h438022dc},
  {32'h44357522, 32'hc38f67ca, 32'hc214493d},
  {32'hc49d5fc8, 32'h412e1630, 32'hc4244e2f},
  {32'h44cd2151, 32'h43ad546d, 32'h42dbbaaa},
  {32'hc5012f62, 32'h42dda8ae, 32'hc312b6cd},
  {32'h44c17e11, 32'h42df69f0, 32'hc189063a},
  {32'hc3dba714, 32'hc3dbc5ef, 32'hc225b8c2},
  {32'h44c1b051, 32'hc321002d, 32'hc33fedc1},
  {32'hc31ae180, 32'hc23f644e, 32'hc19183a4},
  {32'h43ab589b, 32'h42230877, 32'hc28310df},
  {32'hc2b8ee24, 32'h439ae4dc, 32'hc266a567},
  {32'h44cff425, 32'h43a3ef33, 32'h43159bbe},
  {32'hc500ac8b, 32'hc2da9c03, 32'h42d3b58d},
  {32'h44dd960d, 32'hc33d5541, 32'hc3a120b0},
  {32'hc3cd9b1e, 32'h42b10007, 32'hc130e770},
  {32'h43ceafe8, 32'hc3638b23, 32'h44168f30},
  {32'hc47237d4, 32'hc19e2b99, 32'h41fc94fc},
  {32'h44e5f9ee, 32'hc327b1ee, 32'h43329588},
  {32'hc4f7310a, 32'hc30a24f9, 32'hc36119f6},
  {32'h445e0c0f, 32'h42d0d1c3, 32'h43bd5f7d},
  {32'hc439fc2b, 32'h4324a739, 32'h43a6fe54},
  {32'h447d9983, 32'hc362cc33, 32'h428aa63d},
  {32'hc4e22c92, 32'hc30398ae, 32'hc3fa1a64},
  {32'h447c01e2, 32'hc1aaf50d, 32'h438ca776},
  {32'hc5004868, 32'hc12671bc, 32'hc3731976},
  {32'h44b83e88, 32'hc35d4c7f, 32'h42fbc914},
  {32'hc4bac03a, 32'hc1dcdcd7, 32'hc28328a2},
  {32'h450dd066, 32'hc38ae16e, 32'h43868b4d},
  {32'hc46724de, 32'hc245f472, 32'hc3dbe49d},
  {32'h4436f0db, 32'h427477bf, 32'hc31f3694},
  {32'hc4e4bfa3, 32'hc35723bc, 32'hc2d4f9dd},
  {32'h44e77752, 32'hc38503e4, 32'hc33b8b0a},
  {32'hc1e9e580, 32'hc337fd8f, 32'h42e248f8},
  {32'h435a7910, 32'hc3aac612, 32'h431c4373},
  {32'hc4fb8cd7, 32'hc110015e, 32'hc133a226},
  {32'h449c0103, 32'h41c57eda, 32'h41d63094},
  {32'hc49bdc3a, 32'hc33e592b, 32'hc2a63166},
  {32'h4406bb03, 32'hc2a88fc8, 32'hc31fed64},
  {32'hc4ef0e47, 32'hc1b2b231, 32'h431c5420},
  {32'h451f575b, 32'hc3333e20, 32'hc366238c},
  {32'hc4a5b164, 32'h4132d9e9, 32'hc35b44e9},
  {32'h445a4dcc, 32'h41b9993b, 32'h43bf2e28},
  {32'hc4da3fdf, 32'h43c5730c, 32'h42df2922},
  {32'h42c03258, 32'hc18bfca6, 32'hc41053c8},
  {32'hc4df257d, 32'hc3840e8e, 32'h435bebbc},
  {32'h44ac4ae1, 32'hc3a00907, 32'hc231285e},
  {32'h3f95d000, 32'h42ea4588, 32'hc3ff74c2},
  {32'h441523a1, 32'h4209c1c6, 32'h429b3e60},
  {32'hc4dde647, 32'hc25cf5b6, 32'h43819069},
  {32'h42364f50, 32'h432b395a, 32'h416551c2},
  {32'hc3ee264c, 32'h436aaf88, 32'hc38de490},
  {32'h450a0830, 32'h432ba38b, 32'hc32ecac0},
  {32'hc4025bb8, 32'h431a747e, 32'hc39babeb},
  {32'h44cbd035, 32'hc38dad1c, 32'h435d2bc6},
  {32'hc47ecd8d, 32'h437afbdb, 32'hc1ab3dc8},
  {32'hc2932be8, 32'h4296cc2c, 32'h42b53170},
  {32'h43328c0b, 32'h4323d9d8, 32'hc3312387},
  {32'h44c2a229, 32'hc35c8e85, 32'h4364c1c0},
  {32'hc1756b40, 32'hc33b5ae7, 32'h4337513c},
  {32'h44e591c6, 32'h413e34e6, 32'hc2027fcc},
  {32'hc4a799a2, 32'hc2fc807a, 32'hc201d655},
  {32'h449add4d, 32'h43a8c68a, 32'hc2309728},
  {32'hc5036f34, 32'h42e8d5e4, 32'h42f2f8c9},
  {32'h44dd9697, 32'hc2bd48fd, 32'hc2a62b41},
  {32'hc50eb592, 32'h40ccc431, 32'h42a385ff},
  {32'h45054972, 32'hc39c760a, 32'h4389e8df},
  {32'hc4d9a50b, 32'h42cef8fd, 32'hc2426007},
  {32'h43dfbb5e, 32'h42cdf9cf, 32'h4285c2e1},
  {32'hc506e354, 32'hc3e0dd28, 32'hc1c6e635},
  {32'hc1998f60, 32'hc292617f, 32'h440772bd},
  {32'hc3a1dfd1, 32'h43b43625, 32'hc204f201},
  {32'h45020b92, 32'h41eba428, 32'hc196413a},
  {32'hc4f47558, 32'hc34305e6, 32'h43107d85},
  {32'h43fef047, 32'h43aaeb49, 32'h43a054db},
  {32'h438225c8, 32'hc389bad9, 32'hc312d552},
  {32'h43ac6372, 32'h4296d406, 32'h4348ba76},
  {32'hc3ba0404, 32'hc317b87c, 32'hc352cbd7},
  {32'hc33a6af0, 32'hc2cea996, 32'hc2517f2a},
  {32'h44af0845, 32'h43064109, 32'h4322fc3b},
  {32'hc372e856, 32'h43c06f17, 32'hc401b9ee},
  {32'h4500a86f, 32'h4439152d, 32'h424f81a4},
  {32'hc48969bc, 32'hc333363d, 32'hc2eaec0f},
  {32'h43f99747, 32'h4201ad78, 32'hc360cff9},
  {32'hc51124fd, 32'hc2f25488, 32'h42b659a7},
  {32'h450da259, 32'hc39a0810, 32'h43cfe25e},
  {32'hc4bd6893, 32'hc38a7790, 32'hc2852b91},
  {32'h431ff2fc, 32'h4272c730, 32'h4319a3b9},
  {32'hc4e035fc, 32'hc34b81f5, 32'h424f5390},
  {32'h44d6d570, 32'h4304d134, 32'h43176fe1},
  {32'hc4832adf, 32'hc2b6f442, 32'h41818e79},
  {32'h44a5fdc2, 32'h435d1178, 32'hc29eb667},
  {32'hc4e3516e, 32'hc292f936, 32'hc27b8b0a},
  {32'h44c6c8a2, 32'h42fca7c0, 32'h43808df3},
  {32'hc4d87284, 32'h431cec20, 32'hc3facdee},
  {32'h438b538c, 32'hc250e46e, 32'hc21c3fcd},
  {32'hc411da76, 32'h410384c9, 32'hc349d9e1},
  {32'h44325d22, 32'hc2dda376, 32'hc313d264},
  {32'hc4d69fab, 32'h43b27c23, 32'hc1bca3da},
  {32'h4461eee4, 32'h4198de72, 32'hc2e6cae1},
  {32'hc4b4523e, 32'h434ef82d, 32'hc31921eb},
  {32'h451348a0, 32'h436197b5, 32'h42c3fb10},
  {32'hc3c2bb3a, 32'h413e7f3b, 32'hbe9a9e96},
  {32'h450f8350, 32'h3ff14244, 32'h43c5913e},
  {32'hc4ccdc73, 32'h42eb1e4e, 32'h42faa3bc},
  {32'h45123baf, 32'hc3c07952, 32'hc2dad4c4},
  {32'hc4dc350c, 32'h430fce06, 32'hc4024842},
  {32'h441a34dc, 32'hc08cd454, 32'hc1384303},
  {32'hc4f8ec9c, 32'hc389c4e5, 32'hc310dd34},
  {32'hc3b90ccc, 32'hc37d4494, 32'hc37c56ed},
  {32'hc42fd58c, 32'hc2dcfe41, 32'hc28c842e},
  {32'h44f826e6, 32'hc3145f3e, 32'hc2bdc493},
  {32'hc3d10cbf, 32'h43dab427, 32'hc40e09f4},
  {32'h448f73a6, 32'h40f39004, 32'h42c47582},
  {32'hc493a423, 32'hc2217e85, 32'hc29bb476},
  {32'h44e19e08, 32'h43e3cc43, 32'hc2ae4db8},
  {32'h42b5ba4b, 32'hc2810460, 32'h435c05f5},
  {32'h43d5c735, 32'h4247ac7a, 32'hc32247c9},
  {32'hc5181d61, 32'h43f7a675, 32'h42c7142c},
  {32'h44d5fe3c, 32'hc33c32c0, 32'hc3d5d97e},
  {32'hc471d756, 32'hc2d566f0, 32'hc2e03892},
  {32'h4494bd3b, 32'h439a2b3b, 32'h435871a1},
  {32'hc3fbd818, 32'hc3346fb2, 32'h4383bc51},
  {32'h44ce9c36, 32'hc313ede6, 32'h439e2d89},
  {32'hc47500e5, 32'h43654bdd, 32'hc31af4dc},
  {32'h4367f524, 32'hc28b1183, 32'hc3b5c9ff},
  {32'hbfd90800, 32'h43cf5b50, 32'h421caf82},
  {32'h44a2aba2, 32'h43cba9ed, 32'h42b0c9e6},
  {32'hc4dc5f98, 32'hc31e3e1b, 32'hc1fbec56},
  {32'h4471682a, 32'h441a9583, 32'h427dbfa0},
  {32'hc4e5f6ad, 32'hc3760fec, 32'hc3922e7c},
  {32'h44d7b610, 32'h4389df4f, 32'hc351486d},
  {32'hc44422c1, 32'h42c675a2, 32'h420b5e53},
  {32'h450ae4d4, 32'h4255d5ac, 32'hc3001765},
  {32'hc4d0c778, 32'h4400104b, 32'hc38788ec},
  {32'h44eeffbd, 32'h430d1846, 32'h42768d2a},
  {32'hc33f92e0, 32'h43941575, 32'hc3a3d9a2},
  {32'h44f7ad70, 32'h4403c4c8, 32'h42bf45de},
  {32'hc5105288, 32'h42f9cf53, 32'h4302ec45},
  {32'h4420c91b, 32'hc39d7473, 32'h41e338b3},
  {32'hc2bdd31e, 32'hc2a885bf, 32'hc3abb39a},
  {32'h451f578d, 32'hc31e6058, 32'h441250ad},
  {32'h434fdb51, 32'hc2cfc8d9, 32'h43a7826e},
  {32'h44613102, 32'h411f29f4, 32'h4326ff39},
  {32'h421d64e6, 32'h4384dee0, 32'hc280ca0e},
  {32'h44604e8c, 32'hc20f4469, 32'h42c4ad90},
  {32'hc4943f93, 32'h429b4395, 32'hc322ac44},
  {32'hc251be40, 32'h4392108d, 32'h41737ffc},
  {32'hc4f23b67, 32'h43953b5f, 32'h4333b758},
  {32'h44aa2f83, 32'hc3006f02, 32'hc1832fa1},
  {32'hc50fa85f, 32'h43df6923, 32'h42e15eb6},
  {32'h44422694, 32'hc1e7f920, 32'h42d16528},
  {32'hc3cd6511, 32'h42189de1, 32'h423be568},
  {32'h44ce733d, 32'h43412736, 32'h42a5afe3},
  {32'hc4ac675e, 32'hc2e7ebcf, 32'hc2fb7fcb},
  {32'h447ed0d6, 32'hc2618460, 32'h4367ab74},
  {32'hc4766336, 32'h422304cd, 32'h41ed32ad},
  {32'h4480e03a, 32'hc39ffba8, 32'h4420483f},
  {32'h430b5ce0, 32'hc1f8cf6a, 32'h438a95a6},
  {32'h43e33878, 32'hc1ac47b8, 32'h437846e8},
  {32'hc41fc180, 32'hc41672b4, 32'hc3f2050a},
  {32'h449443ce, 32'hc1fff9fe, 32'h43bc01a2},
  {32'hc4433e54, 32'h40e3150e, 32'h41c0ae10},
  {32'h44e74130, 32'h43810005, 32'hc2a52af8},
  {32'hc3660688, 32'h42f67386, 32'hc2925609},
  {32'h445e9e4e, 32'h428e3682, 32'hc2efb5a9},
  {32'hc4837fdc, 32'hc34c499a, 32'h4267db2a},
  {32'h440138d2, 32'hc2e56bf6, 32'h428b8a47},
  {32'hc3e94718, 32'h43dcb87b, 32'h4354cd00},
  {32'h43583553, 32'h420e8b88, 32'hc22342f3},
  {32'hc2025f00, 32'hc412ba44, 32'hc2d9b6f4},
  {32'h44fb5db8, 32'h4301634c, 32'h43b9b9ce},
  {32'hc5170edb, 32'hc3f1f337, 32'hc32bbfc1},
  {32'h44e88102, 32'hc2ae86ee, 32'hc3296d8a},
  {32'hc404ea78, 32'hc2d5ebc1, 32'h43b1e9d6},
  {32'h4483784c, 32'hc39dbaad, 32'hc3553e7a},
  {32'hc4c28736, 32'hc0a7f3e4, 32'hc3302390},
  {32'hc177d200, 32'h415e1190, 32'h426a9f8e},
  {32'h43603d30, 32'hc1c4b1ea, 32'hc3703fa9},
  {32'hc2b191b2, 32'h4311f733, 32'h435b5b45},
  {32'h410a4b00, 32'h43cd1737, 32'h42ee8e44},
  {32'h431e2f40, 32'h423cd873, 32'hc0f17832},
  {32'hc4169a60, 32'h439ae22f, 32'h439c594d},
  {32'h44145360, 32'hc325d742, 32'hc2acc538},
  {32'hc4d44ca2, 32'h422a83fc, 32'hc385c808},
  {32'h44e82988, 32'hc33ea30f, 32'h42b07cb3},
  {32'hc3ac0f2c, 32'h433a8409, 32'hc2ba3033},
  {32'h446a7130, 32'h43900248, 32'hc39a49eb},
  {32'hc510d719, 32'h431fa1a4, 32'hc2edcea4},
  {32'h42a57b50, 32'h4368578a, 32'h4322564e},
  {32'hc208f380, 32'h431d6bba, 32'hc293478c},
  {32'h44de6a4a, 32'h42297dd4, 32'hc1db711b},
  {32'hc403f365, 32'h438856e3, 32'h415ec3b0},
  {32'h44b44a76, 32'hc33dcb5c, 32'hc41f8879},
  {32'hc4cbf14f, 32'h43984165, 32'h43d2d520},
  {32'h431dd830, 32'h41dd0de5, 32'h43403556},
  {32'hc3f56e80, 32'hc2375806, 32'h43c21072},
  {32'h4495473a, 32'hc34fc9e4, 32'h43a852b5},
  {32'hc503b994, 32'h430b2a5e, 32'h4376b354},
  {32'h44299344, 32'h440fe23c, 32'h42b83f88},
  {32'hc4301982, 32'h41acd62e, 32'h4394bd1a},
  {32'h44b73810, 32'hbfe0c03a, 32'hc32d7dab},
  {32'hc48097b3, 32'h4210d92c, 32'h43f85ac1},
  {32'h44561448, 32'h432767df, 32'h4363facc},
  {32'h41ef7700, 32'h4391e8be, 32'hc2d46802},
  {32'h44c850cc, 32'h43a13c56, 32'h437c8da1},
  {32'hc457f69b, 32'hc348746a, 32'h42a507c7},
  {32'h44dc5983, 32'h43111f81, 32'h43801dea},
  {32'h42c50970, 32'h433fd0f2, 32'h430a6ced},
  {32'h45018916, 32'h41c54b1e, 32'h43c1a50f},
  {32'hc4a8c983, 32'hc2b5d919, 32'h439fe0cd},
  {32'h44e40224, 32'hc2a4fba6, 32'hc2b91e92},
  {32'hc4b16496, 32'h428843eb, 32'h42ab0dbf},
  {32'h4484f3f8, 32'hc394044b, 32'hc3a1244a},
  {32'hc4b8af43, 32'hc2744312, 32'h4149d3f4},
  {32'h44daaf39, 32'hc33c894a, 32'hc38081ae},
  {32'hc3be2dba, 32'h43a329c9, 32'h4305a29a},
  {32'hc32e41a8, 32'hc331c358, 32'h42d82463},
  {32'hc3efb37c, 32'h432404f7, 32'hc300b37e},
  {32'h4146a770, 32'hc087e338, 32'h4298a65a},
  {32'hc4a5c28e, 32'h41404471, 32'hc33a4954},
  {32'h44756fb4, 32'h42a9bc8b, 32'h43a9988f},
  {32'hc4075ee9, 32'h42d8759d, 32'hc3783c7f},
  {32'h44a10217, 32'h42fbebf6, 32'hc462df23},
  {32'hc500a4e2, 32'h436991b9, 32'h43609d80},
  {32'h446b900a, 32'h43eec2f7, 32'h42e089a1},
  {32'h43dfedf2, 32'hc32dea1f, 32'h439f859d},
  {32'h4489a991, 32'h42831d3e, 32'hc3990879},
  {32'hc3842018, 32'h42431515, 32'hc3aa2b49},
  {32'h44cb29bc, 32'hc398febc, 32'hc4063849},
  {32'hc44593d6, 32'hc2351ce8, 32'h42998fc1},
  {32'h441aaf00, 32'h42db3dda, 32'hc2916573},
  {32'hc444ff1c, 32'hc2d62c4f, 32'hc36ab524},
  {32'h43dc1c40, 32'hc3911270, 32'h401f9990},
  {32'hc4d5ce82, 32'h42b447c4, 32'hc280cf96},
  {32'h44d86586, 32'h4192be9f, 32'hc3432777},
  {32'hc4e4b95d, 32'hc3464d6f, 32'hc283607f},
  {32'h4501111f, 32'h43025c74, 32'h434830b2},
  {32'hc4d46625, 32'h41cbf293, 32'hc392f5d8},
  {32'h448f744a, 32'h4270a8cd, 32'hc3f05fd4},
  {32'h432d458a, 32'h42db7856, 32'hc32f84f1},
  {32'h44873702, 32'h43a6d71e, 32'h429a36d8},
  {32'hc502de7f, 32'h4296f8b9, 32'hc1cf8b9a},
  {32'h44d7aa27, 32'h43cc4e9a, 32'hc3177d49},
  {32'hc46a26f0, 32'hc17f03fc, 32'h43e465ad},
  {32'h449b15c6, 32'h420f1306, 32'h43612d47},
  {32'hc32f8ae8, 32'h4278f87d, 32'hc2c83a0f},
  {32'h44f99374, 32'hc3903377, 32'hc37cda6f},
  {32'hc431c77a, 32'h43c5066d, 32'hc297c278},
  {32'h449973f1, 32'hc2cec63b, 32'h430881c3},
  {32'hc4a38b70, 32'h43a5b444, 32'h42140568},
  {32'h43bc82c5, 32'hc36c3c89, 32'hbf1d02d8},
  {32'hc4e162ca, 32'hc306426c, 32'hc2611664},
  {32'h44623106, 32'h42629db8, 32'hc2d613ae},
  {32'hc35802a5, 32'hc2e04206, 32'hc27c71e9},
  {32'h43d62ad8, 32'hc37bfc11, 32'hc203b433},
  {32'h438bb09f, 32'hc327a0be, 32'h43da4215},
  {32'h43f2d66d, 32'hc3498eed, 32'hc380952e},
  {32'hc5035414, 32'hc1c76ece, 32'h41cfd9e0},
  {32'h443b68f3, 32'h438dafd6, 32'h43035582},
  {32'hc37a9b80, 32'h4377d0ca, 32'hc395849e},
  {32'h4422e252, 32'h4298105a, 32'h4419eca5},
  {32'hc50dfdf7, 32'h41e33774, 32'hc3aa5c09},
  {32'h445beb90, 32'h4342c149, 32'hc3320c84},
  {32'hc429e5d4, 32'h432840b8, 32'h43ace835},
  {32'h44157e66, 32'h4345bc80, 32'h4397b25e},
  {32'h42395340, 32'hc3785fba, 32'hc34334b5},
  {32'h44daf277, 32'h43b6226e, 32'hc295498b},
  {32'hc5153164, 32'h42b1d0ac, 32'hc3016375},
  {32'h449c0686, 32'hc328524f, 32'h4385ba50},
  {32'hc4186e16, 32'h413b1eca, 32'hc352cfe3},
  {32'h44f54a5d, 32'h43946cc0, 32'h420e423f},
  {32'hc50d05e9, 32'h4340a20a, 32'h3fc1e055},
  {32'h44954364, 32'hc33a92cc, 32'h42ff21c6},
  {32'hc433051f, 32'h42d00c82, 32'h436e8e2a},
  {32'h44b715fb, 32'hc227af91, 32'h4424ca5f},
  {32'hc3ffb708, 32'hc3a52e25, 32'h42f258b9},
  {32'h447741df, 32'h439c8824, 32'h4319cb90},
  {32'hc4a1b706, 32'hc34ca22c, 32'hbfcc1871},
  {32'h449b31c4, 32'h4345226c, 32'h43330ade},
  {32'hc502d3db, 32'hc33acb28, 32'h43a84cc4},
  {32'h44b3b06c, 32'hc1861770, 32'h43343cda},
  {32'hc4cb8f70, 32'h43d97671, 32'h4325c896},
  {32'h4479cb3e, 32'h437bf449, 32'h42c33f39},
  {32'hc51c52a0, 32'hc381f509, 32'hc11b14e0},
  {32'h43d1288a, 32'hc2b2c72e, 32'hc3aef7da},
  {32'hc410188b, 32'h43d785d0, 32'hc222f9fd},
  {32'h4456b2e0, 32'h4396ac3b, 32'h435d1c15},
  {32'hc49150b8, 32'hc26b8c99, 32'h4368a05e},
  {32'h44428767, 32'hc457c4c0, 32'h42a041a9},
  {32'hc36f1e8a, 32'hc1ccd808, 32'hc3536c8e},
  {32'h443b7eca, 32'hc323b88b, 32'hc389ea61},
  {32'hc4e82472, 32'h442534a6, 32'h439a1dd6},
  {32'h442a9ea4, 32'hc35fbf11, 32'hc1da5fcd},
  {32'hc504c1b2, 32'h433f0622, 32'hc41d2ea6},
  {32'h4476368c, 32'h43a18a01, 32'h439cffcf},
  {32'hc28091a0, 32'h42c5f4e2, 32'h40e9c789},
  {32'h4485ad35, 32'h42d773e3, 32'h4384d973},
  {32'h410d6900, 32'hc303c81c, 32'h421eb392},
  {32'h45050840, 32'h43058e00, 32'hc304e062},
  {32'hc42d73f1, 32'hc2e60c5c, 32'h420c457e},
  {32'h44b4af7f, 32'hc305834b, 32'hc3926088},
  {32'hc4aa2ea7, 32'hc3d78cf3, 32'hc364bb4a},
  {32'h4417e0ee, 32'h437b8145, 32'h426b00ed},
  {32'hc39aa495, 32'h430f9437, 32'hc2995b01},
  {32'h44d5997b, 32'hc345d965, 32'hc3670e51},
  {32'hc5060ac3, 32'hc34e94cc, 32'hc31f6d8b},
  {32'h4425a0d3, 32'hc35a58b2, 32'hc0885d7c},
  {32'hc49391d7, 32'h4362f844, 32'h42995461},
  {32'h43715fa0, 32'hc1350f32, 32'h4330ff90},
  {32'hc48b9a02, 32'h43c8ce6d, 32'h436a4bfa},
  {32'h443ecb80, 32'hc3afcb3e, 32'h4331fe6c},
  {32'hc4f92c50, 32'hc2773725, 32'hc1ab0c1e},
  {32'h4493937c, 32'hc3c1add6, 32'h444194eb},
  {32'hc44809b6, 32'hc379a02f, 32'h42af714a},
  {32'h43d4fe24, 32'hc29f615b, 32'h4239b1eb},
  {32'hc4ab2082, 32'hc35b2036, 32'hc2b42427},
  {32'h439469a0, 32'hc3148ce6, 32'hc1a03ab8},
  {32'hc4d27bbc, 32'h429c2d09, 32'h41ecee13},
  {32'h44ec3967, 32'hc3237d2e, 32'h42e93455},
  {32'hc50e9ccc, 32'h42823c59, 32'hc4062979},
  {32'h45053b8c, 32'hc367c6bd, 32'h42d8bcb4},
  {32'hc336c5d8, 32'hc244ea76, 32'h431c805c},
  {32'h430a3495, 32'h42f79c15, 32'hc3537245},
  {32'hc4ad652a, 32'h43c97b2b, 32'h4378d376},
  {32'h445ea734, 32'h426615a9, 32'h42f0c54e},
  {32'hc46ddb49, 32'h43ad80f6, 32'hc2ddbb3c},
  {32'h44105158, 32'hc3db0a6a, 32'h4380e187},
  {32'hc42998f2, 32'h42cb3710, 32'hc320d2e3},
  {32'h43ab2272, 32'hc3590e1b, 32'h43780e4d},
  {32'hc4676528, 32'hc293c872, 32'hc3160c7e},
  {32'h4479b378, 32'hc3a74780, 32'h43580832},
  {32'hc4e0d265, 32'hc1c11c3f, 32'h43183498},
  {32'h44f683aa, 32'hc33a8a94, 32'hc2b25da3},
  {32'hc3010c90, 32'h43d4b7eb, 32'hc35500a9},
  {32'h44d37fcf, 32'hc2277ae1, 32'hc3cad2d8},
  {32'hc4862576, 32'hc2829c3e, 32'hc38540fa},
  {32'h44cf985a, 32'hc3b852a9, 32'h435d98fa},
  {32'hc4e98633, 32'h42d5d30d, 32'hc217f216},
  {32'h44914236, 32'hc389c499, 32'h42dee8f3},
  {32'hc4d67008, 32'h437335ea, 32'hc3c132ec},
  {32'h4410cf24, 32'h430f0741, 32'h42afa01f},
  {32'h43a78400, 32'hc1bd82bc, 32'hc1d2f778},
  {32'h43ee663b, 32'hc3864057, 32'h42c610b9},
  {32'hc30ba680, 32'hc3659a70, 32'hc26e8f40},
  {32'h442bb5d0, 32'hc331be72, 32'h436fc534},
  {32'hc46ba9cc, 32'hc1601f17, 32'hc3a03796},
  {32'h44ab6268, 32'hc2a5b216, 32'h42d83b90},
  {32'hc484fa0b, 32'h431290dc, 32'hc32fd826},
  {32'h43e972fe, 32'hc3823a75, 32'h436f3e17},
  {32'hc4f80447, 32'hc38ce7e3, 32'hc3aa1275},
  {32'h44fa472a, 32'h43a05b8d, 32'hc1bc1139},
  {32'hc436e718, 32'h43d1f81e, 32'hc2c17349},
  {32'h44c8123f, 32'h43434b34, 32'hc2a7bc2a},
  {32'hc4abf8a6, 32'h41cba8b1, 32'h423fcbb5},
  {32'h43c030d4, 32'hc288233b, 32'h4359ed58},
  {32'hc4d1c555, 32'h4295ebf4, 32'hc3277d89},
  {32'h45238fc8, 32'h42041549, 32'h4311a5ed},
  {32'hc478fee9, 32'h43350e76, 32'h43a6753c},
  {32'h44eaa852, 32'hc3bc41bf, 32'hc30b1829},
  {32'hc3805b20, 32'h432578e6, 32'h42d0c93a},
  {32'h44cecc0c, 32'hc34e83cf, 32'h43065823},
  {32'hc3eefa14, 32'h436363ac, 32'hc3065047},
  {32'h4470acc5, 32'h433d000c, 32'hc3f2e553},
  {32'hc4992a16, 32'h430ee636, 32'hbfae9260},
  {32'h44a7a9f5, 32'hc13e6f2c, 32'hc3c8c186},
  {32'hc4e7787b, 32'h426ded7a, 32'h42c24ab2},
  {32'h44967048, 32'h432f914a, 32'hc1fd2f1b},
  {32'hc4f6c5fc, 32'hc1d0e950, 32'hc1bb1780},
  {32'h446a0800, 32'hc0fe5613, 32'h43092f7d},
  {32'hc320ba90, 32'h43c77e7f, 32'hc3603d33},
  {32'h44e87bb2, 32'h427ed393, 32'h4385e8e8},
  {32'hc4a55ce2, 32'h43fb5d85, 32'hc30c866e},
  {32'h44e20f55, 32'h4366cd50, 32'h4384a248},
  {32'hc44f8a76, 32'h43ec51d6, 32'h4330e65d},
  {32'h42cc2300, 32'h4326ea73, 32'hc2e3b733},
  {32'hc49adca0, 32'hc359a470, 32'h43e7be68},
  {32'h451b0b3c, 32'h43091a74, 32'h42f5c30f},
  {32'hc4870e88, 32'h43be5057, 32'hc2f5037f},
  {32'h4443f49b, 32'h42addbfc, 32'hc328c163},
  {32'hc3959ce8, 32'h42cdb814, 32'hc2c152da},
  {32'h4428f716, 32'hc3ae1b68, 32'hc224dde0},
  {32'hc4e33b9f, 32'hc26125b7, 32'hc29e7e00},
  {32'h44d0c98a, 32'hc379dfce, 32'h43569bc9},
  {32'hc5161b08, 32'h43a5dac5, 32'hc24b0782},
  {32'h44caf9dc, 32'hc302e382, 32'h42e9cca6},
  {32'h436a8b8a, 32'h434ebc8b, 32'h43e167f1},
  {32'h43d4c300, 32'hc3a608b1, 32'hc24fcc68},
  {32'hc5004b78, 32'hc3c5aa1e, 32'h43c94f73},
  {32'h44f8b3e2, 32'hc2a2d57d, 32'h43b774b7},
  {32'hc483fbd4, 32'h4102c350, 32'hc27676a4},
  {32'h43d64db0, 32'hc31aea02, 32'hc2970100},
  {32'hc408dabb, 32'h42cfdd00, 32'hc344170c},
  {32'h44cbc364, 32'h420fc1a9, 32'h43422c43},
  {32'hc4ff085e, 32'hc420d7d6, 32'h42b14d0c},
  {32'h44cd0d4e, 32'hc164887c, 32'h42b1c85f},
  {32'hc516ecac, 32'h428647ee, 32'hc35a00ac},
  {32'h44de6400, 32'h423c25d5, 32'hc31d3ce3},
  {32'hc494dcee, 32'h427debb2, 32'hc3b02ddd},
  {32'h424c35a0, 32'h42905dc5, 32'h436562e3},
  {32'hc390f0bf, 32'h43ebd915, 32'hc388f2a1},
  {32'h44b0788a, 32'hc390463a, 32'h42d929fd},
  {32'hc4a970c2, 32'hc1381456, 32'h416c0068},
  {32'h444a31b4, 32'h438171ca, 32'hc33b2b9b},
  {32'hc4cb3e8c, 32'h41b8b2b7, 32'h4350b2fd},
  {32'h44e67a8f, 32'h434798f9, 32'h4307f3f8},
  {32'hc4c311bd, 32'hc1e58821, 32'h42ace64c},
  {32'h450d4ed3, 32'hc2b96881, 32'h4326fd8f},
  {32'hc3d8ea28, 32'hc3576da8, 32'h430276b6},
  {32'h43ae17ea, 32'h42fd4414, 32'h438e3651},
  {32'h421322e0, 32'h42be71b8, 32'hc360ffcb},
  {32'h446ac5d4, 32'h43b08ab9, 32'hc3f14bb7},
  {32'hc4300e70, 32'h43508413, 32'hc2d5779d},
  {32'h450b9a87, 32'hc3c256a3, 32'hc32b04e5},
  {32'hc4136df4, 32'h408e01aa, 32'h438b2c27},
  {32'h41cccec0, 32'h43666263, 32'hc27252c0},
  {32'hc4621d00, 32'hc293f977, 32'hc1932e16},
  {32'h4501bd58, 32'h43082589, 32'hc1947e61},
  {32'hc394ded2, 32'h43ac0631, 32'h437a9afe},
  {32'h44de5e6a, 32'h432bcb2d, 32'h43927d33},
  {32'hc3774e50, 32'h42a0154b, 32'h42e09230},
  {32'h451f0e13, 32'h42cec779, 32'hc2c17bc8},
  {32'hc48f206b, 32'hc32bcdca, 32'h4305ffa0},
  {32'h44b7f0e0, 32'hc2ab3b07, 32'hc2816133},
  {32'hc4c616c3, 32'hc19ecc06, 32'hc29c0eba},
  {32'h44a62e4e, 32'hc1bad789, 32'h42ae8687},
  {32'hc4dceaa0, 32'h43219b53, 32'h4312019b},
  {32'h444ac8c8, 32'h428dea47, 32'h3f9bc108},
  {32'hc50147ff, 32'hc17a423d, 32'h42caa457},
  {32'h44eb74d2, 32'hc3d271e3, 32'hc2dafc6e},
  {32'hc0f4a200, 32'hc302e120, 32'hc31609de},
  {32'h440e4a9e, 32'hc33c1f64, 32'h43432621},
  {32'hc4f3ca4b, 32'h4318998f, 32'hc353878e},
  {32'h4502eeeb, 32'hc405bfa8, 32'h42e4f06c},
  {32'hc4fdf808, 32'h43b20f54, 32'h4296d3a6},
  {32'h423f3ec0, 32'hc344a664, 32'h42335d92},
  {32'hc49b6322, 32'hc3210c13, 32'h425ba9b1},
  {32'h442b3b29, 32'hc37c10c3, 32'h4081082a},
  {32'hc486aac4, 32'hc32b105b, 32'h437fb600},
  {32'h450c93b5, 32'h427201cf, 32'h419d4126},
  {32'hc4c45ecd, 32'hc314074c, 32'hc21d2266},
  {32'h4496e4df, 32'hc30d9070, 32'h4364dabd},
  {32'hc4e4a43d, 32'h44071b8b, 32'hc37fd490},
  {32'h44bfa851, 32'h411c1ad7, 32'hc3605bae},
  {32'hc4ad4d3a, 32'h42b63388, 32'hc36e46eb},
  {32'h44482de6, 32'h43095b33, 32'hc3c554b2},
  {32'hc4a45df0, 32'hc3dfc61c, 32'hc3577987},
  {32'h44d81bda, 32'hc0bed51b, 32'h42b2cdba},
  {32'hc4d7ef77, 32'hc3283542, 32'h438f5f72},
  {32'h450392e9, 32'h425be006, 32'hc29139f0},
  {32'hc303a660, 32'hc296b16e, 32'h424dd20f},
  {32'h450c1106, 32'hc2d2f4de, 32'hc2260996},
  {32'hc51747d2, 32'hc11cdf7b, 32'hc2c6be15},
  {32'h442e7524, 32'hc2d54342, 32'hc314e5e8},
  {32'hc4e6be0b, 32'hc2063da2, 32'hc3b42e43},
  {32'h44e0ef6d, 32'hc1cba596, 32'hc2b187d0},
  {32'hc4e0a98a, 32'hc30ba6f1, 32'h4392ac0f},
  {32'h451522b3, 32'h4224471a, 32'h41d50425},
  {32'hc48d411d, 32'h429b1d36, 32'h43065a88},
  {32'h43e63f21, 32'h4047a3ea, 32'h42d0a8d4},
  {32'hc41f2490, 32'hc197c257, 32'h42832807},
  {32'h44f92379, 32'hc2a6d818, 32'hc340c246},
  {32'hc3c41fc8, 32'hc0b8c378, 32'h43ca02cf},
  {32'h445819fd, 32'hc393c13f, 32'h41d48eae},
  {32'h4110e240, 32'h43f5d570, 32'hc284a991},
  {32'h43c801c9, 32'h42834829, 32'h429e8603},
  {32'hc4382834, 32'h42528fd2, 32'h435fd37c},
  {32'h4416a0c0, 32'h427382c6, 32'hc37c1ea0},
  {32'hc50138f7, 32'hc2e556d4, 32'h42889229},
  {32'h43bc1b91, 32'h435a2637, 32'h40cdc2ab},
  {32'hc4ce00e0, 32'hc2ed4f83, 32'hc274ccc6},
  {32'h450b7060, 32'hc3a7846c, 32'hc3c54ec3},
  {32'hc40e6ba9, 32'h43a8ca8b, 32'hc388e278},
  {32'h4514f070, 32'h43e3272c, 32'hc23b0f3a},
  {32'hc4453ae6, 32'hc2d96677, 32'h4370bed0},
  {32'h449ff44e, 32'hc113828d, 32'hc2d05ef5},
  {32'hc3820028, 32'h41fa862a, 32'hc2ebfc5c},
  {32'h447d27f4, 32'h437b2dbe, 32'hc366d839},
  {32'hc4bf23a2, 32'hc3195ea7, 32'hc3f7322e},
  {32'h4483492e, 32'hc3a186b2, 32'hc3c369cb},
  {32'hc4fdbd2a, 32'h3f2cf98c, 32'hc231e607},
  {32'h447399da, 32'h42c254f8, 32'hc3811835},
  {32'hc4b256aa, 32'h43ba8420, 32'hc2bc6d82},
  {32'h43acb9f4, 32'h435c3536, 32'h43a958ca},
  {32'hc496e69e, 32'hc35a2d5c, 32'hc2c949ff},
  {32'h44a1a29a, 32'hc2ec438d, 32'hbff2cc70},
  {32'hc43d00da, 32'h43620967, 32'h42b8e9db},
  {32'h44af96ec, 32'h43c61a85, 32'hc2af19a0},
  {32'h430698f6, 32'h427c4539, 32'h43a3b61f},
  {32'h44f207fd, 32'hc33e7488, 32'hc30a01c3},
  {32'hc4df855a, 32'hc3aaf57c, 32'hc30c7c7d},
  {32'h44ca110f, 32'hc3af33d1, 32'h41c02ec6},
  {32'hc4df0798, 32'hc22245c6, 32'hc3484c29},
  {32'h447199a4, 32'hc360c889, 32'hc2d90c61},
  {32'hc400da72, 32'h4350c46b, 32'h4383f5f2},
  {32'h44589ca4, 32'hc2f87a03, 32'h42e37f56},
  {32'hc45d5450, 32'h42e0f03b, 32'h42ce56c0},
  {32'h44aacbd3, 32'hc2771802, 32'hc3b55856},
  {32'hc46fa60d, 32'h431b3771, 32'h43f0d4e2},
  {32'h4502387e, 32'h42dbc9fd, 32'h42471521},
  {32'hc3542580, 32'h418de6f4, 32'h41efdbe6},
  {32'h441ad844, 32'h432f5a28, 32'hc39ab3c8},
  {32'hc46d09cd, 32'h4367dd06, 32'hc21b727e},
  {32'h44950b93, 32'h431ae494, 32'hc2a7fc78},
  {32'hc32cc250, 32'h43392fbe, 32'h42c07619},
  {32'h44e1397f, 32'hc1f93f0d, 32'hc35998e5},
  {32'hc4da77b6, 32'hc2d3fe5b, 32'hc30eaa90},
  {32'h449bcaa5, 32'hc3a0f7ac, 32'hc32d647d},
  {32'hc3234e16, 32'h431da478, 32'h430f2129},
  {32'h4406c6e8, 32'hc38546c2, 32'hc386d9ef},
  {32'h44c3aef0, 32'h432e59a8, 32'h435c3946},
  {32'hc4c49091, 32'hc3a34462, 32'h41d8b654},
  {32'h451467bd, 32'hc1135435, 32'h439b8f67},
  {32'hc4e6e076, 32'h42173595, 32'hc20cfb88},
  {32'h44361d24, 32'h4279d0e6, 32'hc3659637},
  {32'hc5040702, 32'h435671e2, 32'hc35218a0},
  {32'h44c94b79, 32'hc414ee12, 32'hc384ff6d},
  {32'hc4bbdb72, 32'h4282967e, 32'hc2971bbe},
  {32'h44c5a1b0, 32'hbf0c7c60, 32'hc1d71038},
  {32'hc48bb66c, 32'h42bc26b2, 32'h437a40b2},
  {32'h43a91888, 32'hc2bc5782, 32'hc2a05ecf},
  {32'hc51302a9, 32'hc2060950, 32'hc360c570},
  {32'h44ba77be, 32'hc31c91b3, 32'hc34b7fdc},
  {32'hc4b118ca, 32'h4247f841, 32'hc2d11983},
  {32'h4509dce5, 32'hc2c61df4, 32'h42d20752},
  {32'hc4bde0a4, 32'h43045bd4, 32'hc435a14a},
  {32'hc2ad42a0, 32'hc289f9dc, 32'hc39ff2f3},
  {32'hc4828f90, 32'h421843d5, 32'h4346eabc},
  {32'h44901eba, 32'hc3a1d8b4, 32'hc3cecde1},
  {32'hc4ce3aa6, 32'h4246c0dd, 32'hc402197a},
  {32'h44cc4241, 32'hc32570b1, 32'hc2a79efd},
  {32'hc4cbd02d, 32'hc3e46b89, 32'hc3060087},
  {32'h4495df34, 32'hc3391622, 32'hc3a594d9},
  {32'hc4efbe2a, 32'h430320bb, 32'h43066d97},
  {32'h44b49d5b, 32'h4372aaf5, 32'hc223815c},
  {32'hc38bc31a, 32'h41eda66c, 32'hc0ac3674},
  {32'h43a47e08, 32'hc1ab333e, 32'hc2b9fc7d},
  {32'hc4629a78, 32'h43b5acca, 32'hc35502fa},
  {32'h43d06fb8, 32'h430bbf11, 32'hc2af8d28},
  {32'hc4d377fb, 32'hc222852d, 32'h42a0c73f},
  {32'h4425ec66, 32'h41d540c8, 32'hc3a2af93},
  {32'hc45de70f, 32'hc415a58a, 32'h4313467d},
  {32'h43a5f950, 32'h43f02e48, 32'h433c2605},
  {32'hc4fdd613, 32'hc1e191aa, 32'hc2d22bff},
  {32'h42eb9236, 32'h42c53417, 32'hc3239e20},
  {32'hc433d762, 32'hc3f1bbc6, 32'hbfe3583a},
  {32'h44ae75cb, 32'h434f2bf3, 32'h42b14d37},
  {32'hc4a1425a, 32'h43549710, 32'h43c37696},
  {32'h44e587de, 32'hc1a59152, 32'hc30bfa7a},
  {32'hc3ac8277, 32'h4313122e, 32'h418c99c9},
  {32'h43b68f95, 32'hc28251d3, 32'hc3a095e3},
  {32'hc4dc9d87, 32'h4382a796, 32'h439b168d},
  {32'h44dda6d7, 32'h43173d5e, 32'h43c91b52},
  {32'hc51342ef, 32'h43490aa5, 32'h417b5880},
  {32'h445412bc, 32'h4186a4b4, 32'h43416ff7},
  {32'hc5084d1e, 32'hc31e0fc0, 32'hc3807625},
  {32'h4473c565, 32'h437f9c33, 32'h42a0e956},
  {32'hc4a82030, 32'h438c0202, 32'h434dcf42},
  {32'h4454cf6f, 32'h41d7e4f9, 32'h43178e3f},
  {32'hc50bf5d5, 32'hc3bad0b7, 32'hc2f91b5e},
  {32'h45115419, 32'hc35cc70b, 32'h43638be7},
  {32'hc4adece0, 32'h430ce8da, 32'h432b6fda},
  {32'h4451ab21, 32'hc38959ff, 32'hc2910a93},
  {32'hc4e26087, 32'hc316e2c4, 32'h4303e5bc},
  {32'h43a848d6, 32'h409c0b8b, 32'h42edbd64},
  {32'hc4bae278, 32'hc3670c3e, 32'hc342bc0e},
  {32'h44bea385, 32'h41c24e19, 32'h421f2437},
  {32'hc3433be8, 32'hc3152caf, 32'h43b1c909},
  {32'h451131b0, 32'h438ebe3e, 32'hc4037ecb},
  {32'hc3a7ffe8, 32'h432fa1d0, 32'hc3d1ec65},
  {32'h4518c133, 32'hc3b9035d, 32'h4333df34},
  {32'hc4c1518c, 32'hc3bd753f, 32'hc292673e},
  {32'h43367fc0, 32'h41c34b10, 32'hc33e74ab},
  {32'hc4de5b89, 32'h4382531b, 32'h438362fb},
  {32'h450276af, 32'h43b2e522, 32'h433add72},
  {32'hc4e54ed9, 32'h43bdcce8, 32'h43c2488c},
  {32'h430747e0, 32'hc205dbff, 32'h4228ae88},
  {32'hc4c404fe, 32'h434ada92, 32'h430f7abb},
  {32'h44f1934c, 32'h4121bfd7, 32'hc2a45586},
  {32'hc4cd437b, 32'hc39d62fa, 32'h42bddb74},
  {32'h44b35df9, 32'h43281b52, 32'hc37b906d},
  {32'hc42d48e6, 32'hc3c8d811, 32'h42ff7d6d},
  {32'h4521445c, 32'h43e15c20, 32'h42ae73b6},
  {32'hc485c72b, 32'h42821534, 32'hc3c8a997},
  {32'h44a18a62, 32'h4319e02d, 32'hc2bbc439},
  {32'hc4c2eea3, 32'h414561d0, 32'h431294e8},
  {32'h448b8bae, 32'h42388c66, 32'h3fcf8650},
  {32'hc49080b7, 32'h43790fe3, 32'h42663a2f},
  {32'h4485b876, 32'hc38f6d17, 32'h42e50da0},
  {32'hc48009f4, 32'hc28624b2, 32'hc20ee1f6},
  {32'h44eb0607, 32'hc2e2b589, 32'h4392e901},
  {32'hc395bdf0, 32'h424ebe63, 32'h40225756},
  {32'h44270a9a, 32'h42b46b48, 32'hc30c6238},
  {32'hc388ca58, 32'h430b3a09, 32'hc3ced21f},
  {32'h446fe418, 32'hc404beb2, 32'hc3728a7a},
  {32'hc5063665, 32'h416b1bec, 32'h43852583},
  {32'h44b82577, 32'h407919c6, 32'h43209e30},
  {32'hc500cc19, 32'h4346d0e5, 32'hc393f13a},
  {32'h44406ca2, 32'hc31337a8, 32'h43d9b566},
  {32'hc502f280, 32'h433fb5a5, 32'h4392302e},
  {32'h43e42b97, 32'h422fa57b, 32'h42a1afe3},
  {32'hc4e9ceba, 32'h42cf91c1, 32'h435eb9d0},
  {32'h4427499b, 32'hc3641a63, 32'hc38ab1f1},
  {32'hc44a58d4, 32'h43de372e, 32'h4330d4d7},
  {32'h4496ecc9, 32'hc339a1b9, 32'hc2975ad6},
  {32'hc44bbe4a, 32'hc3b2d96c, 32'h43a29136},
  {32'h4460d4d8, 32'hc37506aa, 32'h439e0f0e},
  {32'hc317f1b0, 32'hc2b24f0f, 32'hc2c91e4f},
  {32'h45061f05, 32'h43a721cc, 32'h4371f539},
  {32'hc3a99bce, 32'hc3103d1b, 32'h4292c1aa},
  {32'h45088bac, 32'h439e04ea, 32'h433b5ea1},
  {32'hc4d33712, 32'hc266f949, 32'hc312cf5d},
  {32'h45130217, 32'h419ef388, 32'h43177dc4},
  {32'hc43bc24e, 32'h42ec2b95, 32'h42566c46},
  {32'h42b785a8, 32'h42da65e3, 32'h429bf7bf},
  {32'hc5098fff, 32'h420abd84, 32'h438e9ef2},
  {32'h4521d682, 32'hc315bdbe, 32'hc381dbb3},
  {32'hc4f7c313, 32'h42c31248, 32'h42a06e42},
  {32'h45059496, 32'h41a2cf05, 32'hc28b1b3a},
  {32'h42c49940, 32'h425502f7, 32'hc380bf48},
  {32'h4506973f, 32'h439fabc6, 32'hc1fe71be},
  {32'hc3a79c90, 32'hc2fccf6a, 32'h43b30ff2},
  {32'h43c76453, 32'h434aff40, 32'hc3ce166f},
  {32'hc50b996e, 32'hc2d2746c, 32'h43234dee},
  {32'h44f01136, 32'hc339983a, 32'hc37e8d6a},
  {32'hc3904398, 32'h40c35944, 32'hc3b05dee},
  {32'h43fdb703, 32'hc34b27a1, 32'h43896d7b},
  {32'hc3906019, 32'hc374e25f, 32'hc32248e6},
  {32'h44a9fc30, 32'hc2293626, 32'hc364ba94},
  {32'hc4973c76, 32'h431adeef, 32'h42a3e739},
  {32'h43e05ec4, 32'h4261ab24, 32'h42a282dc},
  {32'hc497db0c, 32'h431d08fa, 32'h438fa912},
  {32'h4405b934, 32'hc37a4f9c, 32'h43799f6f},
  {32'hc4036b87, 32'hc28352cd, 32'h43a0a8bf},
  {32'h43d3d500, 32'hc30731ae, 32'h4345b280},
  {32'hc3e9e610, 32'hbf0527a3, 32'h441f7b2d},
  {32'h442c0fb2, 32'h40326224, 32'h41a51a7d},
  {32'hc4ceb1cf, 32'hc077ef26, 32'h41764414},
  {32'h44a3e162, 32'h42e457a6, 32'hc3d6403c},
  {32'hc4c2805e, 32'h43512ca3, 32'hc32a565d},
  {32'h44ce81f5, 32'hc360b918, 32'h43926f4c},
  {32'hc4bb42e5, 32'h43b33aa3, 32'h40802442},
  {32'h4512821c, 32'hc37831f4, 32'hc3b3f232},
  {32'hc4943ebb, 32'hc3853175, 32'hc34941dc},
  {32'h44f9abdc, 32'hc17e822f, 32'hc390e718},
  {32'hc4031dee, 32'hc3b27f5e, 32'hc25d06fa},
  {32'h44f7e6e0, 32'h428ab7ef, 32'h429189cf},
  {32'hc4e7d32a, 32'hc3f08bfd, 32'hc2d46c67},
  {32'h44ac846f, 32'h42ce25a9, 32'h438277f1},
  {32'hc4a76ed7, 32'hc11da6f3, 32'h431d6f71},
  {32'h43af34e7, 32'hc38c3f1e, 32'hc3ab9c68},
  {32'hc507a112, 32'hc26fadbf, 32'h4314fb17},
  {32'h44164dc4, 32'h431f4437, 32'hc33ec16b},
  {32'hc3be4090, 32'hc38fbe36, 32'hc2085a14},
  {32'h44b7b62e, 32'h41eff8c3, 32'hc2d895f1},
  {32'hc4fff0c7, 32'hc32674c1, 32'hc3b343c1},
  {32'h44d4a9fa, 32'h427e862a, 32'hc3afdfa7},
  {32'hc4d87b5c, 32'hc371818a, 32'h437c2725},
  {32'h4387303c, 32'hc329ae45, 32'hc325d72a},
  {32'hc2349f88, 32'h4369d079, 32'hc32b5ad3},
  {32'h447e599e, 32'hc1d7f1c0, 32'h41e185ad},
  {32'h41d66d50, 32'hc31a9f88, 32'hc333a56f},
  {32'h4460a829, 32'h433a4208, 32'hc356a9af},
  {32'hc402a1bc, 32'hc295ed52, 32'h43007974},
  {32'h4502a7c9, 32'hc2f932bd, 32'h4321fbe7},
  {32'hc50adee7, 32'h42ffd6b0, 32'hc2efa13f},
  {32'h44e4f097, 32'hc34f0181, 32'hc3523b23},
  {32'hc4feae2c, 32'h4289befa, 32'hc26866fe},
  {32'h44d633c9, 32'hc300b2d3, 32'hc2287439},
  {32'hc4afa6ca, 32'hc21b793e, 32'hc2c81042},
  {32'h44d18e5e, 32'hc2d2acc6, 32'hc3671099},
  {32'hc45fe75f, 32'hc0ec3e3c, 32'h42612374},
  {32'h42fdec24, 32'hc3004c64, 32'hc3706443},
  {32'hc4ab8b6f, 32'hc3d04cb0, 32'hc3883cf7},
  {32'h44b164ab, 32'h42a92034, 32'hc30d71e4},
  {32'hc4e48028, 32'h44019991, 32'h42661a4d},
  {32'h44de5c4f, 32'hc360dfb3, 32'h43968cec},
  {32'hc48a49f7, 32'h43140e84, 32'hc3ba90ae},
  {32'h44961440, 32'hc3555ff4, 32'hc2a2a722},
  {32'hc49f9628, 32'hc2ad4c1b, 32'hc20ca606},
  {32'hc34aec24, 32'hc33de362, 32'h42982000},
  {32'hc4d7a8fb, 32'h43382ee6, 32'hc2bbf696},
  {32'h44da4f53, 32'h422fa867, 32'hc2be4824},
  {32'hc4f88308, 32'hc2897a39, 32'h41f5851c},
  {32'h451775b6, 32'hc32d46d3, 32'h42941ca5},
  {32'hc49685b3, 32'h4328cd4e, 32'hc36af438},
  {32'h447179ce, 32'hc3c4faff, 32'hc27794d7},
  {32'hc3812f64, 32'hc30dc6ca, 32'hc22cc2f4},
  {32'h4459d625, 32'hc3a55faf, 32'hc30b7417},
  {32'hc3674e94, 32'hc3661ff0, 32'hc390baec},
  {32'h446f8807, 32'hc3340029, 32'hc2d59a5e},
  {32'hc4c4f5ab, 32'h4329f3f8, 32'hc30d3f2b},
  {32'h43d4e2d8, 32'h42f1e7e6, 32'hc37b9e1b},
  {32'h42d525c0, 32'h42017371, 32'h41f99d0a},
  {32'h44febef6, 32'hc37df969, 32'h4302dc1f},
  {32'hc49f2870, 32'h42f65d77, 32'hc2819856},
  {32'h43f03ee8, 32'hc369ad41, 32'h42cce5b7},
  {32'hc1ec4eb0, 32'hc31318be, 32'hc35a47ce},
  {32'h448fd644, 32'hc38c8346, 32'h43072a21},
  {32'hc32c2fc0, 32'h43559c6f, 32'h42673da9},
  {32'h42bfaaa0, 32'h430c18e5, 32'hc2b374da},
  {32'hc40a23a3, 32'hc291f850, 32'hc3a13e2e},
  {32'h44c61c1e, 32'hc364219d, 32'h43b91869},
  {32'hc501abda, 32'h435c3495, 32'h425d8dae},
  {32'h44a94391, 32'h439e416b, 32'h4224d90f},
  {32'hc4e89c4a, 32'hc323e412, 32'h43e4b27c},
  {32'h44382390, 32'h435cdb0d, 32'h42de29d3},
  {32'hc4ebebba, 32'hc345ca3f, 32'h40b8bc13},
  {32'h43bc27af, 32'hc2b27efa, 32'h4404ee0a},
  {32'hc4ce1e70, 32'hc31641e7, 32'h424631b5},
  {32'h450606b0, 32'hc333f2d0, 32'hc310b306},
  {32'hc503144c, 32'hc38d5cb8, 32'hc38bab5d},
  {32'h42f94098, 32'h4334d426, 32'hc198c63b},
  {32'hc41d57d8, 32'h43c1aca9, 32'hc3cd1be5},
  {32'h44cd9ebf, 32'h43c65972, 32'hc2c7b24c},
  {32'hc4d8e8a0, 32'h434879c6, 32'h43971029},
  {32'h451f2733, 32'hc20ed276, 32'h4145333e},
  {32'hc2369650, 32'hc3233b8a, 32'hc40534fb},
  {32'h444d5ed4, 32'hc37b974a, 32'h43a42857},
  {32'hc4eea70d, 32'hc2322bf9, 32'h4301de73},
  {32'h434f21e0, 32'hc432501a, 32'h42f24116},
  {32'hc4bfc29a, 32'h43145f17, 32'hc29b0fc5},
  {32'h445485a4, 32'hc1456141, 32'h429e7dd9},
  {32'hc49b65fc, 32'hc342a45c, 32'h429255ed},
  {32'h4401126a, 32'h43a91711, 32'hc347b613},
  {32'hc4c18c24, 32'hc1bf46c6, 32'h4385d48c},
  {32'h44139b77, 32'hc2337e3b, 32'hc31ac2f6},
  {32'hc333de80, 32'h44563356, 32'h41902e51},
  {32'h43c71fe4, 32'hc227d4da, 32'h43ee47b0},
  {32'hc401a974, 32'hc2fa9e88, 32'hc3782ab6},
  {32'h44c3f961, 32'h436367d3, 32'h439baf7e},
  {32'hc4dd75b8, 32'hc218e39a, 32'hc2ba0c8e},
  {32'h4503d2ce, 32'hc39428d2, 32'hc304c9a5},
  {32'hc3a0437c, 32'h424397ee, 32'hc3a6fdc3},
  {32'h43c28f20, 32'hc32b4e92, 32'hc1ce9c67},
  {32'hc4821ad0, 32'hc32683c5, 32'hc284b848},
  {32'h42c9acd0, 32'h4324620c, 32'h43c3b5df},
  {32'hc4666c1c, 32'h44020957, 32'h42a946e1},
  {32'h450a74fc, 32'hc36d263c, 32'hc25e184e},
  {32'h423807c0, 32'hc32b5cb5, 32'hc21d9228},
  {32'h4437ba8a, 32'hc31ef7ed, 32'hbf9c9110},
  {32'hc37dd7de, 32'hc339becc, 32'hc30c9509},
  {32'h44ca0068, 32'hc1b61e51, 32'h41f95fdd},
  {32'hc5035eeb, 32'hc228a4fa, 32'hc318d2f7},
  {32'h440ac2cc, 32'h42382863, 32'hc39077f1},
  {32'hc4c9bade, 32'hc39e4957, 32'h41808034},
  {32'h44d78e0e, 32'h4318516f, 32'h436244cd},
  {32'hc4240d88, 32'hc3138d37, 32'h43f0c48e},
  {32'h44b19b86, 32'hc3b8878a, 32'hc40aba4c},
  {32'hc4a1b237, 32'hc384b37f, 32'hc291351b},
  {32'h44fd9a5a, 32'hc24d8ec1, 32'hc3b9d3f7},
  {32'hc42c6be2, 32'h437fece4, 32'h42d49c73},
  {32'h44cbafea, 32'h43226dcf, 32'hc3052574},
  {32'hc478fc52, 32'h43230765, 32'h43a40c32},
  {32'h44c4e807, 32'h42d0fcbb, 32'h43362b45},
  {32'hc44df182, 32'hc2b688c2, 32'hc2a516b7},
  {32'h44f1c597, 32'h434dc6c4, 32'hc3216cc0},
  {32'hc3dffbb4, 32'hc1b6a4ad, 32'h4272db3e},
  {32'hc1b79080, 32'h43448157, 32'hc373d48e},
  {32'hc3814718, 32'hc354d141, 32'hc2299eb1},
  {32'h430a8040, 32'h43aad2c3, 32'h4190fffc},
  {32'hc4186f98, 32'h4307725c, 32'h43f950d3},
  {32'h44dab1b6, 32'h43d6dc89, 32'h42c978c1},
  {32'hc2365672, 32'h41e5ddb8, 32'h42cdd1ae},
  {32'h44b20265, 32'h435fd0b2, 32'hc15b8dcc},
  {32'hc5009aff, 32'hc3d59e01, 32'h436814e4},
  {32'h43ac03de, 32'h42f9154b, 32'hc3a4198f},
  {32'hc500b9aa, 32'h4338564a, 32'h428b6ec5},
  {32'h44d2036f, 32'h42f26b0c, 32'hc1838424},
  {32'hc3209730, 32'h42f6ad0a, 32'h433d2bff},
  {32'h4505f199, 32'hc3d66ee4, 32'hc334b890},
  {32'hc50c5b72, 32'hc29319a0, 32'hc2b599ff},
  {32'h449e42e6, 32'hc322a39c, 32'hc324e08c},
  {32'hc4a16437, 32'h439193cf, 32'hc304c78d},
  {32'h4509b61b, 32'h4278d812, 32'h42718a7a},
  {32'hc4f6e044, 32'hc2fcc1d9, 32'hbc7d1000},
  {32'hc3261256, 32'hc32e4f17, 32'hc1892db0},
  {32'hc24afa10, 32'hc37b0311, 32'hc2954eb0},
  {32'h44ce06c7, 32'hc2ccf1f9, 32'hc344ea9a},
  {32'hc389f1e8, 32'h42a23e09, 32'hc395a814},
  {32'h4310a430, 32'h43650b57, 32'h433a5a49},
  {32'hc500266e, 32'h438af516, 32'hc17bef6e},
  {32'h452d1f68, 32'h43721a2f, 32'hc36f41bf},
  {32'hc4fa5b24, 32'hc2a0710b, 32'hc3846aea},
  {32'h43ac9638, 32'h4391c20d, 32'hc3c4b164},
  {32'hc51479e5, 32'hc385cacf, 32'hc327e525},
  {32'h43076ba0, 32'hc33771a2, 32'h43284f3a},
  {32'hc40e22b5, 32'h43677981, 32'h428782e1},
  {32'h43ddf7b0, 32'hc3751007, 32'h4363e90c},
  {32'hc46ad5d1, 32'hc3d47e65, 32'hc375fec9},
  {32'h448cb5c6, 32'hc3b869bc, 32'hc31bf275},
  {32'hc4509276, 32'hc2a75f3e, 32'hc3a054dc},
  {32'h44f9507e, 32'h4272c629, 32'h433c21e9},
  {32'hc4f664a2, 32'hc2f5dbb8, 32'h43da2947},
  {32'h44affa13, 32'hc3ac7b8c, 32'hc2eb0031},
  {32'hc4fc942d, 32'hc3d1a284, 32'hc3af618a},
  {32'hc2645ce0, 32'hc2b55ccf, 32'hc2a4610c},
  {32'hc39a49be, 32'hc35fc3c5, 32'hc2b80376},
  {32'h44de2f3e, 32'h434c18ce, 32'hc31acd24},
  {32'hc41555c8, 32'hc24ec1fb, 32'h42596728},
  {32'h43525268, 32'h422941ec, 32'hc31d6562},
  {32'hc313a1d0, 32'hc28ba594, 32'h43ccad39},
  {32'h44cefc39, 32'hc0252e89, 32'h436c89e8},
  {32'hc4507e96, 32'h4339efe7, 32'hc3ca339f},
  {32'h44229953, 32'h4366d638, 32'hc39696ee},
  {32'hc5060071, 32'hc2ead29b, 32'h42c9abec},
  {32'h44b87922, 32'hc31dd982, 32'hc21fc9f4},
  {32'hc4f58d0c, 32'h41da5a36, 32'hc344c1d8},
  {32'h444dc918, 32'h427aaa43, 32'hc38514be},
  {32'h435b05a0, 32'hc25a90c4, 32'h43a39dbe},
  {32'h45090bf3, 32'hc2cdfcf5, 32'h42633545},
  {32'hc49e02e6, 32'h41d94a31, 32'h43a4a68c},
  {32'h451b6411, 32'h433b00da, 32'hc391e0a6},
  {32'hc52a5bb6, 32'hc3c49929, 32'h427f845b},
  {32'h451af161, 32'hc3913740, 32'h429f1971},
  {32'hc5187112, 32'h406448fa, 32'h42c50f0f},
  {32'h441b4e13, 32'hc1d6f2a8, 32'hc38b3fb1},
  {32'hc374aa84, 32'hc2c70498, 32'hc0459f39},
  {32'h452c5ce1, 32'h43020f2e, 32'h42445393},
  {32'hc4f43f11, 32'hc3e522ea, 32'h437a2737},
  {32'h44e775bf, 32'hc184d485, 32'h43d99227},
  {32'hc49d122c, 32'hc399a2c1, 32'hc2fa2e30},
  {32'hc36bae94, 32'hc3016024, 32'hc3138b0b},
  {32'hc46fae1f, 32'h4329cc0d, 32'h41c84ecc},
  {32'h4513f267, 32'h428ad7a5, 32'h42fb0b0a},
  {32'hc40ddedf, 32'hc310b5aa, 32'hc3806b22},
  {32'h44877e73, 32'hc36d395c, 32'hc2ba4ad5},
  {32'hc51130d9, 32'hc38df62b, 32'hc2f5f655},
  {32'h4443c2fa, 32'h4256f6a4, 32'hc383fd48},
  {32'hc4850bf7, 32'h4332ce70, 32'hc3af9e4e},
  {32'h43e5a170, 32'hc28c0567, 32'hc3528ca9},
  {32'hc4cfd52e, 32'hc3e0fc97, 32'hc2155c40},
  {32'h44808f42, 32'hc33e78a0, 32'h43c3227d},
  {32'hc4d57c29, 32'hc385aac9, 32'hc22905ac},
  {32'h44f45725, 32'h42a06786, 32'hc2c699c0},
  {32'hc4ac5b84, 32'hc19d4fcb, 32'h42cf9e2a},
  {32'h441826b0, 32'hc2aa8222, 32'hc3032246},
  {32'hc427d285, 32'hc3c482c3, 32'h43186fb2},
  {32'h446ee996, 32'h42502790, 32'hc2a5d033},
  {32'hc2af62f0, 32'h43850874, 32'h433701c3},
  {32'h438ea970, 32'hc3b58757, 32'h43932b36},
  {32'hc445e244, 32'hc3301540, 32'hc38b6c90},
  {32'h44033bac, 32'h43d1c16c, 32'h4169bee1},
  {32'hc4ecb3ed, 32'hc2c88819, 32'hc2e30604},
  {32'h431e8cb6, 32'h438f0577, 32'h41f0959a},
  {32'hc43510be, 32'h414ac482, 32'hc302707e},
  {32'h44c7405a, 32'hc391f5de, 32'hc322cab2},
  {32'hc46ca8fb, 32'hc292effb, 32'hc41fac7e},
  {32'h44050b6c, 32'hc27e10b4, 32'h41cd031d},
  {32'hc50c5c07, 32'h425cb311, 32'hc3d8dd92},
  {32'h4324f32e, 32'hc353f92c, 32'h437e7a61},
  {32'hc48bde9c, 32'hc3497fee, 32'hc3c3a001},
  {32'h45018420, 32'hc30c0580, 32'hc35f2f1d},
  {32'hc5087104, 32'h421fdca1, 32'h43081ae2},
  {32'h44ece01c, 32'h42bed7e9, 32'hc0a1e6bd},
  {32'hc50da816, 32'hc3491d61, 32'hc333e430},
  {32'h44c7df62, 32'h41f5f770, 32'hc3900068},
  {32'hc4e341c8, 32'h4347308b, 32'h416884a7},
  {32'h4483a286, 32'h434df625, 32'h4385e105},
  {32'hc42d08f0, 32'h41ab7cb7, 32'hc1037143},
  {32'h4510ba5d, 32'hc348d03e, 32'hc19d9eb3},
  {32'hc480af11, 32'hc3492b84, 32'h43566be5},
  {32'h44e042db, 32'hc2c528df, 32'hc2c83098},
  {32'hc4724b5e, 32'h4361d286, 32'hc2bf916b},
  {32'h452f2fc5, 32'h43486ba2, 32'hc30505d3},
  {32'hc39f6900, 32'hc30db6ca, 32'h41c3317a},
  {32'h44d5cab4, 32'h429d1e98, 32'hc35da242},
  {32'hc31063b6, 32'hc24d0590, 32'hc1f25e92},
  {32'h43c748d4, 32'h43c9694b, 32'h421c1208},
  {32'hc2e3691c, 32'hc3af6e33, 32'h4361c02f},
  {32'h44e45bc5, 32'h42cb4f76, 32'h4347782e},
  {32'hc48d5b96, 32'hc310d916, 32'h433865de},
  {32'h4517410d, 32'hc36c6708, 32'h430acbaa},
  {32'h4095a500, 32'h42324253, 32'h431d5155},
  {32'h448f8592, 32'hc265a10c, 32'h43a02f71},
  {32'hc4fce426, 32'h439d61c1, 32'h4354628a},
  {32'h44ac7c04, 32'hc3b56b7d, 32'hc379897c},
  {32'hc44f5112, 32'hc2a81ced, 32'hc0e221ae},
  {32'h44c675d8, 32'hc12e8a84, 32'hc36a0221},
  {32'hc5034f93, 32'hc2e1e14e, 32'h424a2027},
  {32'h440c1ae8, 32'hc25107c8, 32'h44053cc8},
  {32'hc40b3314, 32'hc2c18916, 32'hc3bbaca0},
  {32'h450b6c7e, 32'h42284ade, 32'h40cc3194},
  {32'h42144ea0, 32'hc3b00270, 32'h435b1b2f},
  {32'h450e1a1a, 32'hc2d9ec56, 32'h4320b494},
  {32'hc4bb9ee5, 32'h43461773, 32'h41ae1f03},
  {32'h43676d34, 32'h43ab5ac7, 32'h4350e7ba},
  {32'hc428476c, 32'h430d37f1, 32'hc2576641},
  {32'h45257f86, 32'h43cca0ce, 32'hc2baf398},
  {32'hc506cac2, 32'hc1535405, 32'hc325f9e0},
  {32'h449ff806, 32'h4310d811, 32'h43a1196a},
  {32'hc5036054, 32'hc338dada, 32'h43ddc734},
  {32'h44c7cdf0, 32'hc2d54f47, 32'h4343bc23},
  {32'hc473cb8d, 32'hc433e457, 32'hc2671072},
  {32'h44a9a4a1, 32'h43127fd8, 32'h4357e840},
  {32'hc4f90325, 32'hc2ec0ba2, 32'h42bc4d32},
  {32'h45083c19, 32'h4303a4d7, 32'h4226d500},
  {32'hc4e39df5, 32'h43b15cd9, 32'hc3c11c59},
  {32'h4480001b, 32'h4395fda6, 32'h4395bdbe},
  {32'hc50e802e, 32'h435a3921, 32'h4385bbab},
  {32'h4443d108, 32'hc325c4e5, 32'h42c1dd38},
  {32'hc4c649a4, 32'hc32de157, 32'hc1ea6a6f},
  {32'h43d34524, 32'hc3ab5977, 32'hc2d3b9fc},
  {32'hc4473a66, 32'h418ef117, 32'hc36dbb83},
  {32'h43c8e858, 32'h43aa2ddc, 32'hc38071a8},
  {32'hc503f622, 32'hc3c6e060, 32'h43b33453},
  {32'h44f73e42, 32'h434714ce, 32'hc3459a57},
  {32'hc43f17ac, 32'h425c7c84, 32'hc2412583},
  {32'h447bd4dd, 32'h43831553, 32'hc3b0f31b},
  {32'hc4f00a4a, 32'hc3bd5d86, 32'hc39cd5d2},
  {32'h442e0722, 32'hc409e660, 32'hc09a1a1d},
  {32'hc5132e5b, 32'h438808e6, 32'hc313be96},
  {32'h43d2e900, 32'hc416c04a, 32'hc3f0472b},
  {32'hc5045b9f, 32'h42f679a7, 32'hc30d96e2},
  {32'h449377d4, 32'hc4214332, 32'h41c3e6f4},
  {32'hc2d61816, 32'hc38a6a17, 32'h4338d152},
  {32'h448133c0, 32'h430174ed, 32'hc100b3e0},
  {32'hc499819b, 32'hc39905f6, 32'h419262b9},
  {32'h448bd8ab, 32'hc2b07034, 32'h42cfcb3e},
  {32'hc5225383, 32'h42bf5f54, 32'h43e7b518},
  {32'h44f39c33, 32'h424b6ab3, 32'h4232a77a},
  {32'h43ac099c, 32'hc362df80, 32'hc1db44bf},
  {32'h44022280, 32'h41b24067, 32'h435489f0},
  {32'hc4f88aec, 32'h424cd97d, 32'h43b10217},
  {32'h448f5d1f, 32'hc394fe76, 32'hc29a213b},
  {32'hc388bf38, 32'hc37d8a0b, 32'hc2131db8},
  {32'h44f7d642, 32'h418266f8, 32'hc3068c7f},
  {32'hc4f9cfbe, 32'h41523c93, 32'h43a488a4},
  {32'h44e56edd, 32'h424f9317, 32'h43b0d880},
  {32'hc482a3d1, 32'hc2b93cfc, 32'hc2140245},
  {32'h44acfd06, 32'h4345a53e, 32'h42e9eed0},
  {32'hc4b1db20, 32'h4094c0e1, 32'h42d0b4f5},
  {32'h44ec1559, 32'hc0184ab2, 32'hc20e14f7},
  {32'hc5000a60, 32'h43d8d5c5, 32'hc1e27368},
  {32'h44204885, 32'hc2b6f67d, 32'h40f2a465},
  {32'hc4b60b3f, 32'h43659352, 32'hc3bf79b4},
  {32'h450529d2, 32'hc1697fc0, 32'h419b8269},
  {32'hc4c5df76, 32'hc3d66a8b, 32'h430c4795},
  {32'h431d9b18, 32'hc370133d, 32'h436a240a},
  {32'h42168838, 32'hc2c5d875, 32'hc3127af3},
  {32'h44598af5, 32'h437f3586, 32'h4326b46a},
  {32'hc397de98, 32'hc372f15a, 32'hc2ab09b3},
  {32'hc3f087a0, 32'h43a18877, 32'hc2a07b45},
  {32'hbf347000, 32'h43d5e9b4, 32'h43826c55},
  {32'h43b49c80, 32'hc30989fe, 32'hc1683192},
  {32'h448c2a98, 32'h4322d5ac, 32'h43218fb2},
  {32'hc2cc1f5a, 32'hc3af87cb, 32'hc33c9d21},
  {32'h44d27e9f, 32'h436eec48, 32'h43869dfc},
  {32'hc49fa51c, 32'h424e8622, 32'hc3d4ff6f},
  {32'h44169f7a, 32'h4304e9a1, 32'hc37b5122},
  {32'hc3af45be, 32'h422ab7d0, 32'hc361932c},
  {32'h448880e8, 32'h42a437c6, 32'h43bf44d0},
  {32'hc4ec869d, 32'h4220adf7, 32'hc332d625},
  {32'hc1d1ea80, 32'h430925a4, 32'h42bac004},
  {32'hc389a2c0, 32'hc1adbb9d, 32'h425a79e0},
  {32'h44ad3e5f, 32'hc1972b23, 32'h4304b8c0},
  {32'hc50745c9, 32'hc29039f9, 32'h3fda523a},
  {32'h436c2ee8, 32'h42bf9d2f, 32'hc32e6795},
  {32'hc322ef88, 32'h43c3433d, 32'hc112a2e0},
  {32'h448b3565, 32'hc366b6be, 32'h4295ddca},
  {32'hc3a47dc4, 32'hc336cfcc, 32'hc33235af},
  {32'h4387d92c, 32'hc3bee98c, 32'h4283ff28},
  {32'hc4171e32, 32'hc1a11160, 32'hc3ed0e5a},
  {32'h4500291a, 32'h42543193, 32'h432a962b},
  {32'hc405b682, 32'h424dea3c, 32'h432515fc},
  {32'h44688082, 32'hc2f118cf, 32'h42f8d323},
  {32'hc33a8750, 32'hc3a141d6, 32'hc33cc1be},
  {32'h44d03945, 32'hc3dbff6d, 32'h43a18f82},
  {32'hc3b26f08, 32'hc21b7e0c, 32'h411cd8b4},
  {32'h44dad936, 32'h435610ed, 32'h43aa6ca2},
  {32'hc490e6c7, 32'h431f110e, 32'hc3271396},
  {32'h437d8dc8, 32'h439cc7d0, 32'hc20046fd},
  {32'hc39b5838, 32'hc3232835, 32'hc3395500},
  {32'h44a6bec4, 32'hc3b9e615, 32'h411b772b},
  {32'hc50e77da, 32'h437b4298, 32'hc2919043},
  {32'h43bc747c, 32'hc264cfc0, 32'h41881edd},
  {32'hc4c6fb1a, 32'hc2a3fe5f, 32'hc31d79ba},
  {32'h44da7068, 32'h43989d8c, 32'hc3436f9a},
  {32'hc34f0b98, 32'h4101552b, 32'hc33890e9},
  {32'h43fba23c, 32'h42ea91b8, 32'h42bb05e1},
  {32'hc1cebf80, 32'hc3abf4a0, 32'h431e2540},
  {32'h4440e5bc, 32'h414aa0c3, 32'hc29a5075},
  {32'hc45ba4a5, 32'hc3a107f7, 32'h43403688},
  {32'h44dd3210, 32'hc29b5fb6, 32'h435ecae8},
  {32'hc4a0b79b, 32'hc3174c26, 32'h43af77d7},
  {32'h449972e4, 32'hc3a255eb, 32'h42be5aaa},
  {32'hc462d349, 32'hc2710e4a, 32'hc185792e},
  {32'h423b8500, 32'h40e945de, 32'h4310db6f},
  {32'hc506bea7, 32'h43876dfc, 32'h42c45a1b},
  {32'h449ed59f, 32'h423a7f8a, 32'h43f16f71},
  {32'hc3a3b3d0, 32'h41a37ada, 32'h43db3f59},
  {32'h44ce3cd6, 32'h436d465e, 32'hc1eac2ef},
  {32'hc526a456, 32'hc3192d25, 32'h43e37a52},
  {32'h45053e86, 32'h433baa67, 32'h4322a150},
  {32'hc4271458, 32'h436371c9, 32'h41d240c3},
  {32'h44cf1ac8, 32'hc38642be, 32'h43be2b31},
  {32'hc4455d96, 32'h42679d9f, 32'h43490676},
  {32'h435d7edc, 32'h43083d76, 32'hbf0b3f89},
  {32'hc4ca500d, 32'hc35bd76b, 32'h419430e4},
  {32'h445cbcc3, 32'hc3fb3b7c, 32'hc377d2c2},
  {32'hc4372475, 32'h438b05ed, 32'hc3811bfc},
  {32'h45066637, 32'hc22a79ac, 32'hc33ddb16},
  {32'hc4745efe, 32'h42cf9268, 32'hc28afaf4},
  {32'h423aebce, 32'h440056ec, 32'h434353d2},
  {32'hc46cf9bf, 32'h43395eb4, 32'hc34f29d3},
  {32'h44f91ef8, 32'hc29da56e, 32'h42b2f6d0},
  {32'h43492e5a, 32'hc3994c65, 32'h42bafccb},
  {32'h451e8f7e, 32'hc3b94d13, 32'h435d378e},
  {32'hc3844833, 32'hc27ba7a7, 32'hc396bd9b},
  {32'h44d98428, 32'h436e3cd7, 32'h4325c681},
  {32'hc4b94415, 32'hc32f5c40, 32'h4231277f},
  {32'h449f6620, 32'h41ccb8e0, 32'hc2d9f254},
  {32'h43182910, 32'h42d845ce, 32'h41fe9f81},
  {32'h44896982, 32'hc27fde58, 32'hc28a7c40},
  {32'hc4a8f955, 32'h4305ea7a, 32'hc2ade2af},
  {32'h44d9f6fc, 32'h43911636, 32'hc31e92de},
  {32'hc507699a, 32'h42e5b733, 32'hc14a9f8a},
  {32'h44ab3279, 32'h431def1d, 32'hc2f5143a},
  {32'hc3b4a67b, 32'hc3426e3e, 32'hc3017046},
  {32'h44da6f1d, 32'hc2a9ba6e, 32'hc2b1ba73},
  {32'h4394de3b, 32'hc1d8e0fe, 32'hc1675a78},
  {32'h449ab2e3, 32'hc2808562, 32'h433f0734},
  {32'hc4f7e209, 32'hc329e777, 32'h43800d90},
  {32'h450361a0, 32'h416dd166, 32'h4411795f},
  {32'hc4beaa9a, 32'hc35543d0, 32'h4309c824},
  {32'h44a5c043, 32'h42be78d0, 32'h43989a8a},
  {32'hc4ff3d03, 32'h43a633f1, 32'hc158438d},
  {32'h426f3650, 32'h421097c6, 32'hc2d1eb7e},
  {32'hc447b068, 32'h4345cfb2, 32'h437cf46c},
  {32'h43731acc, 32'h434c0807, 32'hc3389e7b},
  {32'hc44f197c, 32'hc380aa09, 32'h4402363a},
  {32'h44a49534, 32'hc35766f4, 32'hc3b7cda9},
  {32'hc3718f90, 32'hc2a46655, 32'hc09619ae},
  {32'h44c811b2, 32'hc307849c, 32'h42a2ee04},
  {32'hc2a10c70, 32'h4238e2d4, 32'h43099d9b},
  {32'h44c8b66a, 32'hc2e8586c, 32'h431133bc},
  {32'h42ede945, 32'hc2e87f21, 32'h44041bf7},
  {32'h44a69905, 32'hc3918930, 32'hc3b34e3b},
  {32'hc30c1420, 32'h42c29455, 32'h43cb835c},
  {32'h450b10d3, 32'hc3900d0f, 32'h433a5524},
  {32'hc47bb404, 32'hc2a4350b, 32'hc3ce2fc8},
  {32'h44c9d1d4, 32'h4224a7bc, 32'h43a56c8a},
  {32'hc518dd79, 32'hc319a1b1, 32'h440772ba},
  {32'h43aed9f0, 32'h43766b0d, 32'h431a7021},
  {32'hc4a3a284, 32'h43c5be8a, 32'h4287320e},
  {32'h45036397, 32'hc25179de, 32'h43941083},
  {32'hc26017a0, 32'hc2d57531, 32'h431d8ea5},
  {32'h43ab4700, 32'hc35445cf, 32'h435730b9},
  {32'hc46d3181, 32'h434251f4, 32'h42e9cec9},
  {32'h44c79906, 32'hc1f2c85c, 32'h42e1d805},
  {32'hc50b0ac7, 32'hc36f5e40, 32'h434c8549},
  {32'h44ea4426, 32'h4324ccd6, 32'h42e904ea},
  {32'hc434f03f, 32'hc381b2b9, 32'h4275ce60},
  {32'h44eed66a, 32'h42dc60a3, 32'hc2d888eb},
  {32'hc4dfc7df, 32'hc205b9b8, 32'h42e67cc6},
  {32'h42854f00, 32'h41852a00, 32'h438bf1bb},
  {32'hc4fee06c, 32'h4312725d, 32'h41b541be},
  {32'h44d2c3b4, 32'hc3ee6a51, 32'hc2cdd0bd},
  {32'hc5368712, 32'h431a2d09, 32'hc2132f90},
  {32'h44d54390, 32'h42928a1a, 32'hc30364c6},
  {32'hc4bc2b6c, 32'hc2b1e125, 32'h43867c73},
  {32'h4495299e, 32'h43753691, 32'h4352ce1d},
  {32'hc4e87362, 32'h429c9bff, 32'hc1ed9c3c},
  {32'h434b284c, 32'hc2ad214f, 32'h4398037e},
  {32'hc4ac1dfe, 32'h42b4bb44, 32'h42f12953},
  {32'h44e5f82c, 32'hc3a748fd, 32'hc12032f4},
  {32'hc16a4d00, 32'h439414cf, 32'hc1d95450},
  {32'h4520e542, 32'hc172a1b8, 32'hc21ff7d2},
  {32'hc4c28ee5, 32'h3f462920, 32'h429bf456},
  {32'h44e4e14a, 32'hc32d4849, 32'hc222141d},
  {32'hc4bc713a, 32'hc2a5204c, 32'h42a9ce12},
  {32'h44ff4fcc, 32'h429fea98, 32'h41e16eef},
  {32'hc4e0325f, 32'hc299b61d, 32'h440ea9cc},
  {32'h42afd790, 32'hc319a6f4, 32'h4208a5c3},
  {32'hc24c69c2, 32'hc09935d4, 32'hc21227c5},
  {32'h448c668d, 32'hc3b44dfb, 32'hc00d1280},
  {32'hc391b236, 32'hc34ae658, 32'h4284dca1},
  {32'h44484bd2, 32'h42bb6735, 32'hc38ab15c},
  {32'hc422dd17, 32'h43931f4f, 32'hc1d90455},
  {32'h44f16a0e, 32'h43b0e12c, 32'hc39a7adf},
  {32'hc5076600, 32'hc1b43cca, 32'h43964749},
  {32'h44c6a218, 32'h417f8e4d, 32'hc1694350},
  {32'hc451c181, 32'h4371eb9e, 32'hc360adf1},
  {32'h40ea0d00, 32'h439b0be2, 32'h4328ac31},
  {32'h423c78ae, 32'hc33eea63, 32'h4305167b},
  {32'h44d844fd, 32'hc3024171, 32'h41b86a4e},
  {32'hc4d425d8, 32'h428c89b8, 32'h4378feb2},
  {32'h44dfee1b, 32'hc3b44901, 32'h439fe3c1},
  {32'hc479ac9e, 32'hc29542b3, 32'h43cc7f4d},
  {32'h4514b7e0, 32'h444ec624, 32'h429075de},
  {32'hc4b4d844, 32'h43abde01, 32'h43136316},
  {32'h4437557b, 32'h43bf6188, 32'hc32c8b82},
  {32'hc40947ea, 32'h43342d68, 32'hc1ce82db},
  {32'h44569ad2, 32'hc31c0a7d, 32'hc1252e5c},
  {32'hc306b2b8, 32'hc1b86400, 32'hc249b6d3},
  {32'h43dcb194, 32'h4329639d, 32'hc1a3b885},
  {32'hc4919584, 32'hc224cb8d, 32'hc34b9dda},
  {32'h4415cfc5, 32'hc31430e2, 32'h4237966f},
  {32'hc503afd2, 32'h42688138, 32'hc2c36205},
  {32'h44bc2265, 32'hc37def3f, 32'h436eb1cd},
  {32'hc4f6d8fd, 32'h4319612f, 32'h41dd54a1},
  {32'h4515f88f, 32'hc2b6a900, 32'h4293c613},
  {32'hc432a58c, 32'hc40fe467, 32'hc384c57c},
  {32'h4490c1ae, 32'hc34c0406, 32'hc3801a6c},
  {32'hc43656c8, 32'hc3415e59, 32'h4252962f},
  {32'h44d67bba, 32'h4307f442, 32'hc1a52c3a},
  {32'hc4e68079, 32'h41b93358, 32'h430503b0},
  {32'h43d05f44, 32'h4308e09b, 32'hc2bc81fc},
  {32'hc4cc5fdd, 32'h43c1c987, 32'hc39d73bd},
  {32'h45116535, 32'hc38193bd, 32'hc29b303f},
  {32'hc4d7b7e7, 32'h432c4806, 32'hc3637d7a},
  {32'h449ab429, 32'h435eeae6, 32'h430529b6},
  {32'hc42067f9, 32'h41612413, 32'h436b2cc8},
  {32'h44633f8e, 32'hc2e5a2eb, 32'hc36115cb},
  {32'hc3a1c20b, 32'h433cd228, 32'hc1fccdb7},
  {32'h43ee6c12, 32'hc226fd82, 32'hc3c811b3},
  {32'hc401168c, 32'hc192219a, 32'hc35668d3},
  {32'h4491de46, 32'h43cc7947, 32'h4411a600},
  {32'hc504c5a0, 32'h43d520ac, 32'hc3f93f29},
  {32'h43ceecc0, 32'h4390c71a, 32'h43903276},
  {32'hc26f37c0, 32'hc381171e, 32'h437e4fbe},
  {32'h45038ce6, 32'h430a3530, 32'hc3c19910},
  {32'hc4e08970, 32'h43911ce2, 32'h4380e576},
  {32'h44ab485c, 32'hc3510454, 32'hc10c6046},
  {32'hc439e6ac, 32'h4397bef2, 32'hc35e967c},
  {32'h443e412d, 32'h42c9146a, 32'hc2657512},
  {32'hc48368f2, 32'hc3b5ceb6, 32'h4201c4ac},
  {32'h44c15afe, 32'h433e92d2, 32'hc1d476a2},
  {32'hc497f7a7, 32'h420cb587, 32'h433e9a54},
  {32'h440f62de, 32'hc282874e, 32'h40aa1227},
  {32'hc48ac232, 32'h42e90b3c, 32'hc3ac4b99},
  {32'h43d32c38, 32'hc36e4927, 32'hc2950190},
  {32'hc527a6ba, 32'hc2c81a6f, 32'h42b1a1e7},
  {32'h44bfc2e6, 32'hc2e1ee71, 32'hc36908eb},
  {32'hc4f83dfe, 32'hc35f2d46, 32'h43528ab3},
  {32'h44b32edd, 32'h4229850c, 32'hc199726c},
  {32'hc31bc620, 32'h435aa00e, 32'hc29dab17},
  {32'h44c029f6, 32'h43194c71, 32'h42baeb2a},
  {32'hc4fde1ed, 32'hc3083b0b, 32'hc3565b67},
  {32'h41ddff00, 32'h41e0deff, 32'h43ab5b53},
  {32'hc410fe7c, 32'hc2ad0119, 32'h435bd586},
  {32'h43aa3b85, 32'h4329c1cf, 32'h4380e156},
  {32'hc43406ac, 32'h3fef9358, 32'h4133e762},
  {32'h44a1547b, 32'h43152f30, 32'h432a13d4},
  {32'hc48f5710, 32'h40bca703, 32'h427a1f56},
  {32'h446b3ac8, 32'hc2e9ccfd, 32'hc35502f5},
  {32'hc4d2b32f, 32'hc269b53d, 32'h42ce5653},
  {32'h451aa14e, 32'hc39b9587, 32'hc30f4d5d},
  {32'hc4a2f74f, 32'h43d19b40, 32'hc3809497},
  {32'h450108fe, 32'hc40391bf, 32'h426c0714},
  {32'hc178b000, 32'hc37b1ce1, 32'hc3dd7269},
  {32'h4481b76a, 32'hc22dddff, 32'hc377217c},
  {32'hc432c2ca, 32'hc2bb15dc, 32'h43d08b10},
  {32'h4452754c, 32'hc323669d, 32'h42b5e1f7},
  {32'hc33de410, 32'hc1b32e31, 32'hc40ea1b5},
  {32'h449a2a4a, 32'h4361fe3f, 32'h429847b0},
  {32'hc46fc640, 32'hc2be0ce2, 32'hc18ec610},
  {32'h44cdaf6e, 32'h431b7e7f, 32'h420a9ae8},
  {32'hc4ee31b1, 32'hc3d6f462, 32'hc389b48d},
  {32'h44d80f33, 32'h43938148, 32'h431381be},
  {32'h42ddc53c, 32'hc2ac586c, 32'h4157cc75},
  {32'h4455b845, 32'h42f97d8d, 32'h418f9161},
  {32'hc4e4f7fe, 32'hc36677de, 32'hc2383bef},
  {32'h41aef4a0, 32'h42a4b01e, 32'h43a4ee36},
  {32'hc4d8b572, 32'h439783bc, 32'hc22b1b22},
  {32'h44176806, 32'hc301b4e6, 32'hc3eaa42f},
  {32'hc4399220, 32'hc202d184, 32'hc29bc7ac},
  {32'h43cd08fb, 32'hc34090a0, 32'hc38f44c6},
  {32'hc2f22361, 32'h43933bb4, 32'h4365bd70},
  {32'h450bca4c, 32'h433f7fe8, 32'h42e8319c},
  {32'hc496ff60, 32'hc3287ee2, 32'hc2cd9cef},
  {32'h447aea3a, 32'h43abc58f, 32'hc0ef30fe},
  {32'hc48b8e85, 32'hc33e1bb7, 32'hc35bf185},
  {32'h44ac5f2d, 32'h42b5684d, 32'hc38fa611},
  {32'hc4a5e556, 32'hc2be73c6, 32'h41829516},
  {32'h445c4672, 32'h4288845d, 32'hc312724d},
  {32'hc4400f4c, 32'hc29ec317, 32'hc3c1523a},
  {32'h4446bc82, 32'hc28f7917, 32'h42dca8e8},
  {32'hc464ac6c, 32'h42a73e66, 32'h433ef59e},
  {32'h44e411f6, 32'h43098489, 32'h42b7cebf},
  {32'hc4d429f3, 32'hc3bcd347, 32'hc15ebd4e},
  {32'h448c361e, 32'h438465c4, 32'h432d776c},
  {32'hc4816fe5, 32'hc29d93ea, 32'hc3a58503},
  {32'h44a3fb67, 32'h431cc803, 32'hc28a9fa2},
  {32'h42cb22eb, 32'hc2781483, 32'h42e9bf77},
  {32'h44092e2c, 32'h435ff7a3, 32'h4325aa7e},
  {32'hc5110e31, 32'h43b4450a, 32'hc21314ff},
  {32'h442e390c, 32'h42daa0a8, 32'hc27371c0},
  {32'hc4cb1914, 32'h436cf036, 32'h42bc86da},
  {32'h448e1e6c, 32'hc3b2c178, 32'hc293a9ec},
  {32'hc5018539, 32'h42aa2bd2, 32'hc3888b98},
  {32'h43df8e50, 32'h4308b624, 32'hc36d4f8d},
  {32'hc2ce7d00, 32'hc25e8b4e, 32'h42f71200},
  {32'h45128c97, 32'hc3128b24, 32'h43164830},
  {32'hc47c73e8, 32'h436ab28c, 32'hc2dc2e2d},
  {32'h448f25c8, 32'hc2baf990, 32'hc3604ed8},
  {32'hc46055ef, 32'h4396bba2, 32'h42793163},
  {32'h447fe437, 32'h434cdcc2, 32'hc0ac8714},
  {32'hc4966c14, 32'hc33800d7, 32'hc2d86deb},
  {32'h4505c658, 32'hc251513f, 32'hc3a015bf},
  {32'hc43f71ca, 32'h44055fba, 32'hc38db20e},
  {32'h4486a363, 32'hc3bfc925, 32'h43e28aba},
  {32'hc45c1304, 32'h428f2369, 32'hc30f4a41},
  {32'h45023317, 32'h425ce878, 32'hc317baae},
  {32'hc49b0b95, 32'hc3b8edaa, 32'h43c15721},
  {32'h450a83bb, 32'hc38d941e, 32'h41994689},
  {32'hc319d706, 32'h432ea1da, 32'hc34bb8a2},
  {32'h44264d78, 32'h41971dbe, 32'h43471361},
  {32'hc4843a13, 32'h4332c05d, 32'hc384b74f},
  {32'h4506144c, 32'h43dcceca, 32'h4336a46d},
  {32'hc40f2eda, 32'h42913dae, 32'h415f1d07},
  {32'h43ee2e90, 32'hc29a5724, 32'hc2a6bb7d},
  {32'hc4e7f829, 32'h43a9106f, 32'h42e16246},
  {32'h44b462c6, 32'h4265de73, 32'hc218abe0},
  {32'hc3aea46a, 32'h437cafc5, 32'hc3efe3b9},
  {32'h443ad60f, 32'h4239f63c, 32'hc2277e7d},
  {32'hc4a55fd3, 32'hc232f085, 32'hc415f27b},
  {32'h4499512e, 32'h40f8fea1, 32'hc350074a},
  {32'hc4b16549, 32'hc1d0732b, 32'hc3ad3d67},
  {32'h450505bd, 32'h41f8b108, 32'h424ec4e4},
  {32'hc42df05a, 32'h43dd5f56, 32'h43132fe6},
  {32'h4464de3a, 32'h425dcefc, 32'h420127eb},
  {32'hc414cb06, 32'h439c462b, 32'h42cdfac5},
  {32'h43a01afa, 32'h43458f8e, 32'hc32e6cf3},
  {32'hc4d218ca, 32'hc3204fc7, 32'hc3fd3adc},
  {32'h4470bb4e, 32'h432ede13, 32'hc266eb80},
  {32'hc5019f17, 32'hc23b3767, 32'h42b95e62},
  {32'h43f54b7c, 32'hc324ff48, 32'h434bdd3d},
  {32'hc445de7f, 32'h43125127, 32'hc3ee5ad1},
  {32'h44a34bc5, 32'hc1a8da7f, 32'hc12d322c},
  {32'hc4daf8fc, 32'hc2d3c36e, 32'h4295b97e},
  {32'h44f734df, 32'h4250776a, 32'hc33d40c2},
  {32'hc4b0f26d, 32'hc39e028e, 32'hc31ea760},
  {32'h448446a1, 32'h42707cd4, 32'hc2820126},
  {32'hc3a3051c, 32'hc295413d, 32'hc364ff92},
  {32'h40f08e00, 32'hc35b840b, 32'h432fac4a},
  {32'hc4c1f9ce, 32'hc262eb12, 32'hc3dd9a2e},
  {32'h449c110e, 32'hc235e796, 32'hc1b5d1c4},
  {32'hc2a0f892, 32'hc379d53b, 32'h4267f680},
  {32'h42e00340, 32'h42ca7b4c, 32'h42e1d867},
  {32'hc50005f9, 32'h431f7a3a, 32'hc299ac3d},
  {32'h44369018, 32'hc3505964, 32'h4360ab18},
  {32'hc48409c2, 32'hc2b6128c, 32'hc4229184},
  {32'h44ad54ea, 32'h43b497c9, 32'h439cb280},
  {32'hc3449d50, 32'hc3f95a01, 32'hc1cc9814},
  {32'h434d8058, 32'hc35022bd, 32'h4398372a},
  {32'hc520206c, 32'h434679c3, 32'hc2989c82},
  {32'h44000748, 32'hc1c6cad2, 32'h43c86a08},
  {32'hc418c770, 32'hc2a02650, 32'hc2e8d036},
  {32'h44ff808e, 32'hc344108e, 32'hc3045134},
  {32'hc4e25134, 32'hc384d080, 32'h4220db77},
  {32'h43948f30, 32'h43706f51, 32'h4287ae40},
  {32'hc48129e1, 32'hc370f4ab, 32'hc1a0ee40},
  {32'h44e75bdf, 32'h41bf3feb, 32'h43757be6},
  {32'hc4f2cf29, 32'h434cfa83, 32'hc335d83d},
  {32'h445d3dda, 32'hc330b914, 32'h42ef36e6},
  {32'hc4dbcaa9, 32'hc3c6f5a4, 32'hc2c5657b},
  {32'h44f5aa59, 32'h431e20a3, 32'h43cf2bdd},
  {32'hc4df1c10, 32'hc32fd367, 32'h42f12433},
  {32'hc3124b10, 32'hc24c2224, 32'h42c89194},
  {32'hc496c028, 32'h43ca9843, 32'hc316590e},
  {32'h448d3cc0, 32'hc1c09ffc, 32'h42b52b68},
  {32'hc38b4fd2, 32'hc33d3fc8, 32'h420a8d24},
  {32'h449a6aa6, 32'hc3e51a50, 32'h43a7c8c5},
  {32'hc2e35500, 32'h425ca640, 32'hc37fe10c},
  {32'h449e28da, 32'h41586880, 32'h411d5070},
  {32'h42fc7eaa, 32'hc30c098b, 32'h417bd452},
  {32'h44e386e7, 32'h43581850, 32'h43e5b8d4},
  {32'hc4f9cbca, 32'hc38195c6, 32'h429a33a9},
  {32'h44cf90f0, 32'h43293374, 32'h43f59daa},
  {32'hc33ed550, 32'h4288ae52, 32'h43744787},
  {32'h444de8a2, 32'h432420c7, 32'h4352c6d2},
  {32'hc4dca9e1, 32'h42480e8e, 32'hc3a189f6},
  {32'h44b8062d, 32'h4398ea78, 32'h430c5440},
  {32'hc4f993b1, 32'h43b48ac0, 32'hc2b2eae8},
  {32'h44e6dd55, 32'h434be044, 32'hc3486321},
  {32'hc5006f16, 32'h4251345b, 32'h42e94763},
  {32'h44eba19a, 32'h4289590b, 32'h406b0389},
  {32'hc4497c38, 32'h4253b4ec, 32'h4205fa97},
  {32'h43da1fe4, 32'h43365842, 32'h41a84bc4},
  {32'hc2c2fc60, 32'h427ef184, 32'h431440f2},
  {32'h44686082, 32'hc39e9319, 32'hc2de4158},
  {32'hc4d3a798, 32'hc19fd714, 32'hc39616d4},
  {32'h43c02074, 32'h42bf1be6, 32'hbfeaf46c},
  {32'hc4831056, 32'hc3fc7fe2, 32'hc209a41c},
  {32'h4505062e, 32'h43002d97, 32'hc297ab40},
  {32'hc3bd4cd0, 32'hc2d87480, 32'hc344b062},
  {32'h44da724c, 32'h423dcdb7, 32'h426b5ed8},
  {32'hc5093eab, 32'h434a8505, 32'hc3914182},
  {32'hc3ac16f0, 32'h43336e65, 32'h43610a72},
  {32'hc4f9a707, 32'h43537a61, 32'h42ac7435},
  {32'h441da1b8, 32'h43003e56, 32'h421e7bf3},
  {32'hc5049308, 32'hc31a52f0, 32'h41197a86},
  {32'h44aa851c, 32'hc2562634, 32'hc2d5db35},
  {32'hc3f8e459, 32'hc2a72272, 32'hc1b31a3f},
  {32'h450097cf, 32'h42a11191, 32'h438382dc},
  {32'hc494a442, 32'h42ee11dc, 32'hc269185c},
  {32'h449b447c, 32'hc399fb71, 32'hc3467630},
  {32'hc48c5e7b, 32'h4301083c, 32'hc3cf3510},
  {32'h451bc4da, 32'hc38ecdc6, 32'h41c85b96},
  {32'hc1ebe86f, 32'h43496d2d, 32'h4375c7ba},
  {32'h44c888dd, 32'hc311ff4d, 32'hc1db8607},
  {32'hc4f7685c, 32'h42dbe2dc, 32'hc2fb4542},
  {32'h4445aa68, 32'h43a4c6e4, 32'hc36683e9},
  {32'hc4765e23, 32'h4304b977, 32'hc2579b14},
  {32'h44a5d9ce, 32'h4378bcc5, 32'hc3de9e49},
  {32'hc43f93d9, 32'hc30252be, 32'h43b50c77},
  {32'h4511f33b, 32'h420334ef, 32'hc383deb5},
  {32'hc48c276a, 32'h419037b9, 32'h43601e92},
  {32'h43a5b710, 32'h4395129c, 32'hc2ba81f0},
  {32'hc483f3b6, 32'h4273be70, 32'h43593fd8},
  {32'hc2c21690, 32'hbe866520, 32'h4304b241},
  {32'hc4dfc988, 32'h423840cc, 32'hc3bc9467},
  {32'h43e92d81, 32'hc2275d03, 32'hc35adf67},
  {32'hc4b00277, 32'hc322461a, 32'h43cadd64},
  {32'h44915fb6, 32'h4355b4ad, 32'hc15cc2d4},
  {32'hc3b9a100, 32'hc1b3ffef, 32'h400b5d5a},
  {32'h4507af10, 32'hc318b481, 32'hc38b80eb},
  {32'hc3f51890, 32'hc31b085c, 32'h43a8ccba},
  {32'h44de1fbb, 32'hc38ed9b1, 32'hc1babf44},
  {32'hc5011bb8, 32'h4359bee1, 32'h43816ef9},
  {32'h4498c097, 32'h430b65aa, 32'hc24b2f49},
  {32'h43014626, 32'hc3a28d43, 32'hc413bcdb},
  {32'h4520f0ee, 32'h43214c24, 32'hc2e6db8b},
  {32'hc41b9908, 32'h42cae885, 32'hc2e2652a},
  {32'h44b354ca, 32'h4223539f, 32'h430c1fc9},
  {32'hc4d6f229, 32'h43227c62, 32'h43fec5d0},
  {32'h440dd2a6, 32'h4151947f, 32'h41c0064d},
  {32'h41cf7480, 32'h43508a9d, 32'h42dafab9},
  {32'h430f25b0, 32'h42f19a8a, 32'h3fdee10d},
  {32'hc4135660, 32'hc3abe58a, 32'hc4032a5c},
  {32'h44ce2326, 32'h433d5687, 32'hc3db1f6e},
  {32'hc48f10a0, 32'hc30c4873, 32'h43dd2a28},
  {32'h44aa99f4, 32'hc35fc1b4, 32'hc35c17bf},
  {32'hc498f0a4, 32'h43051ff1, 32'h431b4007},
  {32'h4388ee60, 32'hc3448604, 32'h4338f405},
  {32'hc48cf787, 32'hc1bde7e0, 32'hc311c185},
  {32'h443bc104, 32'hc3944c5c, 32'hc2984dc3},
  {32'hc4757536, 32'hc2d81fcf, 32'hc30d12de},
  {32'h43e4632c, 32'h43114f69, 32'hc2d2f074},
  {32'hc328219f, 32'hc3494c34, 32'hc30bf30c},
  {32'h44b5461f, 32'h4365823f, 32'hc23e469b},
  {32'hc4acbd9e, 32'h42915ee6, 32'h433a545a},
  {32'h43ec4f33, 32'h412c9a88, 32'hc27c2120},
  {32'hc4fdf912, 32'h42446f14, 32'h4243713a},
  {32'h443a2374, 32'hc2875d6c, 32'hc36ae5a2},
  {32'hc4f61678, 32'h41ab0c88, 32'h4210dc92},
  {32'h4459aada, 32'hc2764450, 32'hc3826f8b},
  {32'hc4b6f2b7, 32'hc270f8da, 32'hc311bd67},
  {32'h440d1184, 32'hc2d37eee, 32'h429d9166},
  {32'hc498103d, 32'hc37e1971, 32'h42b84b8c},
  {32'h448abde2, 32'hc34915ed, 32'hc3015f8b},
  {32'hc374394c, 32'h41b7885e, 32'hc1578609},
  {32'h4435fa44, 32'h43a07008, 32'hc28f6d18},
  {32'hc4d3d156, 32'hc383ea48, 32'hc33a208a},
  {32'h43c94d30, 32'hc386b8f1, 32'hc2eb8563},
  {32'h431d09d0, 32'h431d0225, 32'h43e1a978},
  {32'h44f3c130, 32'h42a1e177, 32'hc34d3190},
  {32'hc406dd88, 32'hc1106e3a, 32'h430efbc5},
  {32'h432b77f7, 32'hc2a16d28, 32'hc24b39ca},
  {32'hc4939ad5, 32'h4218d7b0, 32'h431b940e},
  {32'h448aaa63, 32'hc2a91618, 32'hc3789336},
  {32'hc3d1d8c2, 32'hc3a7b7d3, 32'hc2a4ae02},
  {32'h43659e68, 32'h41419254, 32'h42cf79f7},
  {32'hc438b696, 32'h43bf21a4, 32'h4232b268},
  {32'h445998c4, 32'h4331d238, 32'hc2cdbf6c},
  {32'hc51396f9, 32'hc3553f74, 32'h43b8e8bf},
  {32'h44de388b, 32'h43820c5c, 32'h42c8c0c7},
  {32'hc3fad200, 32'hc3d6a3c0, 32'h41eadc12},
  {32'h44a8f0c5, 32'h42b77ed1, 32'hc380590d},
  {32'hc4ebcb79, 32'hc303d218, 32'h42fd3a9b},
  {32'h44ce8d60, 32'hc3d6d566, 32'hc31a98de},
  {32'hc29d7ebb, 32'hc363ba38, 32'hc268373c},
  {32'h44fb2a49, 32'h42b8baf3, 32'hc2cce550},
  {32'h44602a7d, 32'hc2f10df4, 32'h3fdcb3e4},
  {32'hc4ce1caf, 32'h42abc3d3, 32'h43db4261},
  {32'h447cd8dc, 32'hc3a40677, 32'hc2a745eb},
  {32'hc40f3aac, 32'hc34abb76, 32'hc3870e3f},
  {32'h4414c0f8, 32'h442b681d, 32'hc3259650},
  {32'hc423deba, 32'h43b5ede5, 32'hc30b0985},
  {32'h42cb6fc8, 32'h4308bd9f, 32'hc1ffdd7b},
  {32'hc49e63a2, 32'h430885e0, 32'hc3c96ed3},
  {32'h4431f3c0, 32'hc3932756, 32'hc1bd5d14},
  {32'hc41dd1cd, 32'h43cb3488, 32'hc2fd24c1},
  {32'h42461350, 32'hc2fefcbb, 32'hc3a1566e},
  {32'hc494e1f0, 32'hc2d80198, 32'hbff4d4cc},
  {32'h443a89ab, 32'h43790d9b, 32'hc39d8b6c},
  {32'hc3ebc88c, 32'hc3a8a3c7, 32'hc3da4ea9},
  {32'h4461e46e, 32'hc3b1dfb0, 32'hc3209d25},
  {32'hc45afaf6, 32'h42ae8bdc, 32'h4114473e},
  {32'h44ca1148, 32'h4391f580, 32'h420500a0},
  {32'hc4984445, 32'hc296ac37, 32'hc2cccc32},
  {32'h449c9afa, 32'h43ea606a, 32'h430d9461},
  {32'hc4e95ada, 32'h438cbf5e, 32'hc2d7cbdc},
  {32'h432d35c0, 32'hc3a5f063, 32'hc347343e},
  {32'hc48bdb29, 32'hc3b28fa9, 32'h4342fe83},
  {32'h44feee14, 32'h4367a610, 32'h4374698e},
  {32'hc465468c, 32'h4380370a, 32'hc33b07fe},
  {32'h450dd61f, 32'hc0a03273, 32'h42be37b2},
  {32'hc2dd6278, 32'h433f5f33, 32'h42b36037},
  {32'h44c2a50b, 32'h41de4360, 32'hc22ff3bb},
  {32'hc405c665, 32'hc321d274, 32'h43c76a5c},
  {32'hc1af5c80, 32'h4298c10f, 32'hc405bd30},
  {32'hc49da053, 32'hc30e4e91, 32'hc33d2985},
  {32'h4502f1ce, 32'hc20e490c, 32'hc32763c4},
  {32'hc4d7e458, 32'h42da19ff, 32'h4249eed0},
  {32'h44ef23e9, 32'h441aa5e7, 32'h4333f587},
  {32'hc42f4004, 32'hc318d51b, 32'hc23bf448},
  {32'h4477c4e2, 32'hc38c7e42, 32'hc36a9082},
  {32'hc50c1997, 32'h41c8d1af, 32'hc1772eb1},
  {32'h448bc4ec, 32'hc333f578, 32'hc386413a},
  {32'hc478e4d9, 32'h440f31c2, 32'hc33784df},
  {32'h448c9370, 32'h423c92db, 32'h43d43c61},
  {32'hc4501e16, 32'h4303a737, 32'h42985426},
  {32'h4370c484, 32'hc185b436, 32'hc2d72da5},
  {32'hc3e0933b, 32'h430e9900, 32'h42914bc1},
  {32'h45077da7, 32'hc399b4e5, 32'h43ab3119},
  {32'hc40dd2c9, 32'hc303fb4c, 32'h437de843},
  {32'h44268016, 32'h42d7f81f, 32'h432929ed},
  {32'h429d7f40, 32'h408e4b30, 32'h43c32cb2},
  {32'h44de16b3, 32'h42857d50, 32'hc2da8c8d},
  {32'hc41b6fc8, 32'h4153f262, 32'h43982208},
  {32'h446010ba, 32'h428662fe, 32'h4365df38},
  {32'hc4310108, 32'hc35956e3, 32'h4210612f},
  {32'h4498e777, 32'hc391ad2f, 32'h42e094a5},
  {32'hc41ad410, 32'hc346dd1c, 32'hc2fe1aa5},
  {32'h44a56b51, 32'hc2680923, 32'h439f97b2},
  {32'hc443f78b, 32'h4375c755, 32'h4355780c},
  {32'h4446e152, 32'h43afb0a7, 32'h41f7c914},
  {32'hc45fc47f, 32'h43cf370d, 32'hc34c0440},
  {32'h4500c09b, 32'hc30dd574, 32'hc3585e2d},
  {32'hc444b2d8, 32'hc07206d0, 32'hc34c0e88},
  {32'h448c2ba5, 32'hc26190a4, 32'hc32a0b9a},
  {32'h431907f0, 32'hc3e35e2a, 32'hc3ddb4d4},
  {32'h44171c85, 32'hc4170d3f, 32'h4316060b},
  {32'hc382fa68, 32'h42ca5e38, 32'h4327ec50},
  {32'h4507644c, 32'hc3526191, 32'h4346c31e},
  {32'hc38c2986, 32'h43365582, 32'h428c3563},
  {32'h44c42134, 32'hc36dd679, 32'hc3b4512e},
  {32'hc4a50927, 32'hc2e4fac6, 32'h44220f04},
  {32'h43537c28, 32'hc1a3e09a, 32'h3fb85a38},
  {32'hc3ddb0ae, 32'h41df20e2, 32'hc16a89d4},
  {32'h4439d119, 32'h43f6d232, 32'h429de621},
  {32'hc4bc6060, 32'hc25d1c09, 32'h43e082da},
  {32'h4508371d, 32'hc2c1cb88, 32'h43c1ae1d},
  {32'hc49d1006, 32'hc37e7574, 32'h4253cce4},
  {32'h44107805, 32'hc358d203, 32'hc39d9ac2},
  {32'hc4cbfd1a, 32'hc2fc131e, 32'h419de1e4},
  {32'h45021fac, 32'hc3397305, 32'hc3a99145},
  {32'hc40a9ad0, 32'h432b3563, 32'h42f94e6f},
  {32'h442a059d, 32'h42995e60, 32'h428327e2},
  {32'hc4cd2955, 32'h438e30c5, 32'hc3dbe916},
  {32'h445b71b8, 32'h42ebdd52, 32'hc380e85b},
  {32'hc4d9be9a, 32'hc399c5de, 32'h436c2015},
  {32'h4434e9e2, 32'hc33d10de, 32'hc2e5ec43},
  {32'hc4c8d6ce, 32'h420fa9ed, 32'hc30d467d},
  {32'h4402fc79, 32'hc3ae0bd1, 32'hc300f736},
  {32'hc3d56fa2, 32'hc2ad9062, 32'h41116282},
  {32'h44e40047, 32'h42eef481, 32'h41f88abd},
  {32'hc500463c, 32'h429e8086, 32'h439afd55},
  {32'h44492dba, 32'h430c0578, 32'h438c7342},
  {32'hc44f8784, 32'hc36673f5, 32'h430a0109},
  {32'h44a90161, 32'h3fac67c2, 32'hc2a609cb},
  {32'hc4ed5dac, 32'hc3d29c2a, 32'hc391c026},
  {32'h4523f790, 32'hc26bea30, 32'hc33ea3ba},
  {32'hc46176a4, 32'h42cf9c2a, 32'h435ad050},
  {32'h449b3d0e, 32'h42042986, 32'hc331e2c8},
  {32'hc4f76994, 32'h433616bb, 32'hc33c1186},
  {32'h4451878c, 32'h421d062b, 32'hc284fbac},
  {32'hc4d2e835, 32'hc35a9845, 32'hc2ecb623},
  {32'h44d6e4fa, 32'hc2a2d9c2, 32'hc32fde7c},
  {32'hc4c444f7, 32'h424a6fe8, 32'hc1ded870},
  {32'h452648ce, 32'hc2aeda9a, 32'h42b98694},
  {32'hc42058b6, 32'h41b4cd28, 32'h4399220c},
  {32'h436a6938, 32'h42b15fbe, 32'hc3952bd1},
  {32'hc47914ac, 32'h428ee261, 32'h4306a7fa},
  {32'h44344758, 32'hc2394fa2, 32'h43ba1f50},
  {32'hc4cd89e4, 32'hc1d66756, 32'h433fcae6},
  {32'h43c05d14, 32'hc3a8d46f, 32'hc29a6ff3},
  {32'hc4fbb578, 32'h42cbe2da, 32'hc22528d6},
  {32'h439cb782, 32'hc3e39dd1, 32'h438609bd},
  {32'hc4c50b23, 32'hc3e85f10, 32'hc3135442},
  {32'h44cc5199, 32'hc2f89af4, 32'hc3c8dc5a},
  {32'hc4898c70, 32'hc20308ba, 32'h41f41260},
  {32'h44d41e7e, 32'hc321aa81, 32'hc303eabe},
  {32'hc48b9411, 32'h42a703df, 32'h4350d507},
  {32'h44ab485a, 32'hc34608e7, 32'hc128d43f},
  {32'hc41239d8, 32'hc2bb4d7c, 32'h4339699c},
  {32'h442bbd09, 32'hc2dd40a3, 32'h436d0be9},
  {32'hc49aa9c7, 32'hc39d35d9, 32'hc258e1db},
  {32'h45076974, 32'hc1e69e28, 32'hc3936c2b},
  {32'hc4ef443b, 32'hc3032247, 32'h42251e0e},
  {32'h44454cae, 32'h42e43da7, 32'hc375ee9d},
  {32'hc4e1bc8b, 32'h43148fc8, 32'h42a3ec1b},
  {32'h42e641bf, 32'hc2509539, 32'h426cd2c6},
  {32'hc4d8ac1e, 32'h439bc759, 32'h42f8714d},
  {32'h44cf292b, 32'h42ac6a40, 32'hc1d65db5},
  {32'hc40ce641, 32'h4309cd55, 32'h438d3590},
  {32'h43fe93bf, 32'h424a860d, 32'h4326674b},
  {32'hc479fa2a, 32'h43756461, 32'h4328359c},
  {32'h4520fb02, 32'hc2d3d7bf, 32'h43438339},
  {32'hc3a20730, 32'hc32478ff, 32'hc3374d97},
  {32'h44f7bc97, 32'h4338a858, 32'h436ee93d},
  {32'hc48d9252, 32'hc341f909, 32'h43a99e61},
  {32'h44287eb6, 32'h4328db52, 32'h438d0024},
  {32'hc4887362, 32'hc2ca612a, 32'h41a46fe3},
  {32'h44f34aeb, 32'hc2a36ab0, 32'h4113452e},
  {32'hc4ef3ace, 32'h4344f09f, 32'hc27815e1},
  {32'h44ce2988, 32'hc3ad76da, 32'h421e3c70},
  {32'hc4e92240, 32'h42ca0680, 32'hc2e8cded},
  {32'h44bb4d08, 32'hc36b4e16, 32'h433e361d},
  {32'hc3bb424c, 32'hc4033c3b, 32'h4284c355},
  {32'h45018340, 32'hc185b520, 32'h438ad39f},
  {32'h425119c0, 32'h43371814, 32'h418ac208},
  {32'h44c643e3, 32'hc33793a4, 32'hc2e163bb},
  {32'hc4e09081, 32'hc2540647, 32'hc2dda9d8},
  {32'h44208c24, 32'hc2a8e585, 32'hc3852d8f},
  {32'hc4815998, 32'hc32fd39d, 32'h44289c93},
  {32'h43c4c148, 32'h4281caf5, 32'h43792350},
  {32'hc48840f8, 32'hc29fc971, 32'hc36f145c},
  {32'h44e0dc5b, 32'hc3066222, 32'h401e4c0c},
  {32'hc47013ef, 32'h4357ef0f, 32'h4250dd3c},
  {32'h44d6cbca, 32'h4297d77c, 32'h428d41c8},
  {32'hc4f2f67a, 32'h439d4c9c, 32'h437caa46},
  {32'h44842775, 32'hc211916c, 32'hc297fbdc},
  {32'hc4662738, 32'hc3aa1d15, 32'hc30c3073},
  {32'h42194380, 32'hc373f22f, 32'hc1cf49bd},
  {32'hc31bca1c, 32'h430342dc, 32'hc4093ac7},
  {32'h44ea0f63, 32'hc2c4986c, 32'h42d0abdc},
  {32'hc4bd2c4a, 32'hc31ce7de, 32'h4391bb6f},
  {32'h44ff7686, 32'hc4206e46, 32'hc2d5d49c},
  {32'hc4b9b199, 32'h43580367, 32'hc358dbcd},
  {32'h448f3cb5, 32'h437ab7a8, 32'h4265a6bd},
  {32'hc4f259df, 32'h4352d163, 32'h4330cd00},
  {32'h445bac80, 32'h43b04288, 32'hc30f8abb},
  {32'hc4e0e4ac, 32'hc3b4a0fa, 32'h40f2df34},
  {32'h44ee343f, 32'hc2ff13fe, 32'hc2e5935c},
  {32'hc4c9917b, 32'hc2ced3e6, 32'hc19bef3b},
  {32'h449ad5bb, 32'h40d50712, 32'h42ad28e2},
  {32'hc4848382, 32'hc3578b44, 32'hc350a3af},
  {32'h4507f7e4, 32'hc387046d, 32'hc322e00e},
  {32'hc4b575a0, 32'hc2f48f7e, 32'hc3875067},
  {32'h44e6ff70, 32'hc2d9feca, 32'h4267d230},
  {32'hc50ad1c8, 32'hc2d18f70, 32'hc1b3287a},
  {32'h44fee926, 32'h42643bbc, 32'h42442ec1},
  {32'hc02dc000, 32'h436a2e5c, 32'h433731c2},
  {32'h446b4964, 32'hc3e658ca, 32'h43796526},
  {32'hc484a564, 32'h4329c024, 32'h4380f740},
  {32'h446a7501, 32'h438ca515, 32'hc15d8291},
  {32'hc4960a2b, 32'hc3aa4d47, 32'hc35e74f6},
  {32'hc285c5b0, 32'h42495479, 32'h435c7142},
  {32'hc3b012cc, 32'hc38f0d22, 32'hc330d61e},
  {32'h44b044b1, 32'h43a8fab4, 32'h440bc478},
  {32'hc4d33f9c, 32'h43c692f0, 32'hc36694ea},
  {32'h44ff42db, 32'h42ffc6e5, 32'hc2ed3686},
  {32'hc4c9dfd9, 32'hc36877ac, 32'hc388137e},
  {32'h434a6a8c, 32'hc3bdf01f, 32'hc37446e1},
  {32'hc4819c69, 32'hc321761d, 32'hc1267003},
  {32'h438bc000, 32'hc385a11b, 32'hc30de653},
  {32'hc485b67d, 32'h43c25c74, 32'h4305aed7},
  {32'h441a7cb0, 32'h428b8b3d, 32'h422be482},
  {32'hc4eea721, 32'h436f17e1, 32'hc3cca495},
  {32'h43a1e04c, 32'hc35d98b9, 32'h43b8cfe0},
  {32'hc4853923, 32'h43bcde8b, 32'h41800c42},
  {32'h44cbb981, 32'h43b981a6, 32'h41a18542},
  {32'hc4292a83, 32'h4330c3a9, 32'hc3ddb586},
  {32'h440bc2d4, 32'h42cab9e3, 32'h4311f1ea},
  {32'hc4c19e8f, 32'hc1974e69, 32'hc332eeba},
  {32'h4457a63e, 32'h42a92098, 32'h4183eb48},
  {32'hc3162d68, 32'hc121410d, 32'hc358e53a},
  {32'h44c785b4, 32'h4391a0ff, 32'h419012f0},
  {32'hc5034dae, 32'hc39c7869, 32'hc394de86},
  {32'h44799820, 32'h431680b8, 32'hc04360c0},
  {32'hc47482e6, 32'hc2aad4fe, 32'h429e70f1},
  {32'h44f83468, 32'hc3596921, 32'h41e669ea},
  {32'hc4f689f0, 32'hc3058506, 32'h432aa88e},
  {32'h44b6d841, 32'hc381c20c, 32'h4300a79c},
  {32'hc4a0e12b, 32'h4304067c, 32'hc2179d9d},
  {32'h450534b0, 32'hc3505a21, 32'hc35cb6a9},
  {32'hc4be597f, 32'h43aa8d5b, 32'h4320d40e},
  {32'h4498bd8b, 32'hc38fa225, 32'h42fd93b8},
  {32'hc40ad7d3, 32'hc330ff12, 32'hc3b7df1f},
  {32'h44b4a5a8, 32'hc231f504, 32'h42a38ee0},
  {32'hc4c19877, 32'h42121ad3, 32'hc32bcca8},
  {32'h44ed7e89, 32'hc1b4e022, 32'hc3adc0ca},
  {32'hc4f34146, 32'hc2f1e756, 32'hc29672ca},
  {32'h4506b134, 32'h43d708c4, 32'hc3195ac5},
  {32'hc4047507, 32'hc360af00, 32'h4381bc67},
  {32'h42535a80, 32'h3fa7b770, 32'hc19e4182},
  {32'hc4dce896, 32'hc27286bf, 32'h431a8849},
  {32'h44ec38e8, 32'hc36ba88c, 32'hc310d8e3},
  {32'hc50a2cba, 32'h42fd614a, 32'hc2a14e52},
  {32'h43b0d5a5, 32'hc35ad226, 32'hc2fa50cb},
  {32'hc3ea6478, 32'hc269b4db, 32'hc2bf4dcc},
  {32'h45034fc1, 32'hc200d2cf, 32'hc2a428b5},
  {32'hc312a000, 32'h4348f23e, 32'h423e6fb8},
  {32'h4382c889, 32'h41c35e76, 32'h43546548},
  {32'hc4ce456f, 32'h4200d131, 32'h41f816ff},
  {32'h44ce845e, 32'hc3f3613c, 32'hc3c8fb7b},
  {32'hc3fda7bc, 32'hc30c44de, 32'h4207ffbb},
  {32'hc3461c60, 32'hc3f74c77, 32'hc417b799},
  {32'hc5071c14, 32'h43146d43, 32'hc32c68c7},
  {32'h44e11625, 32'h41a88bb9, 32'h43b6a334},
  {32'hc487a08e, 32'hc1920ea8, 32'hc38778cb},
  {32'h443c7e0d, 32'h42219630, 32'h42205155},
  {32'hc4856997, 32'hc280786e, 32'hc36ebef6},
  {32'h4424d701, 32'hc2f57806, 32'hc4064748},
  {32'hc4de43bc, 32'h42d7c107, 32'hc08093ba},
  {32'h44a205eb, 32'h430517c5, 32'hc2bf5d22},
  {32'hc3fcc404, 32'hc37ec842, 32'h4304cfa9},
  {32'h44211764, 32'h43b478bf, 32'hc132ac5e},
  {32'hc40c58e8, 32'hc0bbad0c, 32'hc1f025dc},
  {32'h440ac0ba, 32'hc36405c2, 32'h42a26d0e},
  {32'hc492c15a, 32'h42f5cd3c, 32'hc2ec420a},
  {32'h438456fe, 32'hc2d36393, 32'hc34eb04a},
  {32'hc421bedc, 32'h411733ec, 32'h4351e63d},
  {32'h44d8552e, 32'h430bae70, 32'hc3358ed0},
  {32'hc45e734a, 32'hc32eca1c, 32'h434cdbea},
  {32'h44857266, 32'h434ae306, 32'hc2bc3674},
  {32'hc3eb8a4a, 32'h42d55b05, 32'h42edb9df},
  {32'h450acfe9, 32'hc16d5013, 32'h4348b57a},
  {32'hc4845317, 32'h420ae51c, 32'hc301fa3f},
  {32'h447df295, 32'h421b3909, 32'hc3cb9c71},
  {32'hc4c36e22, 32'hc283961d, 32'h42c8dcd4},
  {32'h44c76cac, 32'h439debef, 32'hc1d6bf29},
  {32'hc4725870, 32'h4414226b, 32'hc36ae278},
  {32'h44880829, 32'hc33c8f16, 32'h4310320b},
  {32'hc4d31b14, 32'h423aad26, 32'hc15c817c},
  {32'h4486b8f7, 32'h431bfe5f, 32'h41fb7b3d},
  {32'hc4de0ac7, 32'hc3dc2868, 32'hc3f2f59c},
  {32'h44f5f2d8, 32'hc242b547, 32'h4380daf8},
  {32'hbddb8000, 32'h4389a260, 32'h43469048},
  {32'h43e09150, 32'h433bd402, 32'h43f1a587},
  {32'hc4125de4, 32'hc3df107e, 32'hc382f028},
  {32'h44e928d6, 32'h43752d49, 32'hc32b581b},
  {32'hc4d0ad4b, 32'h43975e93, 32'hc3967569},
  {32'h44a8ffdc, 32'hc2c82016, 32'hc4120098},
  {32'hc39700d6, 32'hc2a9f84b, 32'h42431952},
  {32'h45287574, 32'hc37bae58, 32'h4304c64d},
  {32'hc4f27916, 32'h434ad044, 32'h433a9bbf},
  {32'h4514b356, 32'h43376059, 32'hc297d354},
  {32'hc5036075, 32'hc2cfb1a0, 32'h4382d6b5},
  {32'h44475893, 32'h440760b0, 32'h432bfc12},
  {32'hc490abfb, 32'hc2bccfa5, 32'hc32ab338},
  {32'h42396f70, 32'h43341cb7, 32'hc3723dc3},
  {32'hc4eea6cc, 32'h426dddf5, 32'hc2505fc6},
  {32'h445dacd4, 32'hc31511ec, 32'hc2dcd786},
  {32'hc4d9cad2, 32'h407c3441, 32'hc36de7b1},
  {32'h443a94bc, 32'hc3e34601, 32'hc3e769bc},
  {32'hc4a25256, 32'h4352f31f, 32'h42fea36a},
  {32'h43b249dc, 32'hc2823268, 32'hc21904f5},
  {32'hc2863ef8, 32'hc3608f46, 32'h438388b6},
  {32'h4470d088, 32'h43811bed, 32'hc3a16fd5},
  {32'h4291e7fc, 32'hc3caeb41, 32'h429ece45},
  {32'h44109839, 32'h44169e76, 32'h43bc826e},
  {32'hc49ad8d0, 32'hc3b680d8, 32'h4355f6ee},
  {32'h4415f5c3, 32'h42092299, 32'hc2b90ad8},
  {32'hc4362efd, 32'hc1edebd7, 32'h4314d004},
  {32'h43123940, 32'h42cd78f4, 32'h425130bd},
  {32'hc1ace2c0, 32'hc3a5a0a0, 32'h41fe916f},
  {32'h43fdeb6c, 32'hc2dde652, 32'hc25f0873},
  {32'hc4b318a5, 32'h434ea6c3, 32'hc34bdcdc},
  {32'h42da7ec0, 32'hc3285f3e, 32'hc2a4a5b2},
  {32'hc4dfd673, 32'hc3016e5f, 32'hc3f5ea5c},
  {32'h449da932, 32'hc346f8b6, 32'h43257c68},
  {32'hc3894798, 32'h433f4305, 32'hc384ab7d},
  {32'h43d9eca2, 32'hc334c666, 32'hc13ff906},
  {32'hc24a4a40, 32'h43f03074, 32'h434a18b4},
  {32'h428be8e0, 32'hc3280b31, 32'hc393fecc},
  {32'hc4945bd4, 32'h43142067, 32'h434e79de},
  {32'h443774ef, 32'h43d4286a, 32'h42a677f5},
  {32'hc484e955, 32'h42884ff1, 32'h432b5e4a},
  {32'h4443f18c, 32'hc1ac1e34, 32'hc37c676c},
  {32'hc495b19c, 32'hc39c657f, 32'h4258936d},
  {32'h44309f5d, 32'h4289b186, 32'h429878e3},
  {32'hc497bd2c, 32'h4284e16f, 32'hc2f7efad},
  {32'h44e21f61, 32'hc31ecd74, 32'hc267b431},
  {32'hc2e77bb4, 32'h43995c89, 32'hc39d099e},
  {32'h44cf4a92, 32'hc1dc3963, 32'hc28d4df1},
  {32'hc51bc22f, 32'hc22b617f, 32'h43301602},
  {32'h44d0f71b, 32'hc200a43d, 32'hc361d9ad},
  {32'hc50abf62, 32'h42f7c63d, 32'h42f37f14},
  {32'h437be2b0, 32'h42cdfc48, 32'hc30c103c},
  {32'hc4299314, 32'h431b09e4, 32'h40f0cf7e},
  {32'h44d66bee, 32'hc2a4f59d, 32'hc22626ef},
  {32'hc48619f0, 32'h43d0ac5b, 32'h43849356},
  {32'h4420aa7c, 32'hc2a272bd, 32'h42120d1a},
  {32'h41cdfd5a, 32'hc297f81e, 32'h432f41f6},
  {32'h448aa616, 32'hc3efce76, 32'h430ebce7},
  {32'hc500c2d1, 32'h431ca82c, 32'h434e6aec},
  {32'h44c0d0b8, 32'hc3c2165f, 32'hc4060dc8},
  {32'hc3e439a4, 32'hc2a5e502, 32'h41e1cf26},
  {32'h45054426, 32'hc38a4c6b, 32'hc398ac2d},
  {32'hc5081a7c, 32'h42c8bc6a, 32'hc3d5d964},
  {32'h440bade6, 32'h42795819, 32'hc1dcfede},
  {32'hc4f9f2a0, 32'h435bebf0, 32'h42eef9ad},
  {32'h44e0684a, 32'hc18e22ff, 32'h4226382d},
  {32'hc4ad5876, 32'h43aa9415, 32'h43682cf9},
  {32'h450be074, 32'hc2351a8b, 32'hc3aeb514},
  {32'hc3a224fe, 32'h42b1fd6a, 32'h42e907ce},
  {32'h44afa910, 32'hc3b185b0, 32'h43660f61},
  {32'hc4a0bde6, 32'h43aed7ac, 32'h4357e77b},
  {32'h451f851e, 32'hc2b23362, 32'h430dc37e},
  {32'hc4627b76, 32'h4385c6cd, 32'h419907ea},
  {32'h4506e941, 32'hc319bb07, 32'hc38b6c71},
  {32'hc4f6d2c2, 32'h43bfdc81, 32'hc29dbbc6},
  {32'h44196294, 32'hc30faf7a, 32'hc361f2a6},
  {32'hc518ae24, 32'h4385363f, 32'h439fb313},
  {32'h43e3a6ae, 32'h43105d03, 32'hc2ee2d91},
  {32'hc5128244, 32'h425570d5, 32'hc1a4b7af},
  {32'h45176cc9, 32'h43a2d467, 32'h435c6198},
  {32'hc40c1b4c, 32'hc368f9b4, 32'h4323e69f},
  {32'h4336c228, 32'hc20c9ce3, 32'hc2d9be38},
  {32'hc34a3390, 32'h41f47717, 32'hc2920949},
  {32'h44b7b4bf, 32'hc3865734, 32'h43d4a83e},
  {32'hc3cb5258, 32'h42cd0af3, 32'hc23a0820},
  {32'h44a7a8b2, 32'h4375075b, 32'hc263e872},
  {32'hc4d28c57, 32'hc3209e0e, 32'h426f8023},
  {32'h447f6b74, 32'h434fc070, 32'h421812d5},
  {32'hc3d2d425, 32'h438633d2, 32'hc241ce04},
  {32'h44072060, 32'hc31e1140, 32'hc250e9e1},
  {32'hc51201c8, 32'h42e7a598, 32'h3f7ede5a},
  {32'h4426ed88, 32'h4320e5f3, 32'hc391b1a7},
  {32'hc4b763a7, 32'hc3d5fe14, 32'h439aa50a},
  {32'h450beeec, 32'hc3cd6dea, 32'hc2956364},
  {32'hc4dad360, 32'h43469640, 32'hbfa3b720},
  {32'h441c34f0, 32'hc3b6f712, 32'h4294603e},
  {32'hc4ba8057, 32'hc2f6c87a, 32'hc18b0d7f},
  {32'h44aa3799, 32'h436560f9, 32'h4337caad},
  {32'hc4dee058, 32'h431db405, 32'h415a3e2c},
  {32'h44dd3efc, 32'h42dfddc1, 32'hc3ba15e1},
  {32'hc50d7098, 32'h438b24c8, 32'h424399bb},
  {32'h44bfe71b, 32'h433a1463, 32'hc2dd696b},
  {32'hc414647a, 32'hc1240f76, 32'hc23ac8b8},
  {32'h4391e6c4, 32'hc1d0df6b, 32'hc35bc800},
  {32'hc41c5baf, 32'h42a17b5b, 32'h42c7ad46},
  {32'h44de20d1, 32'h4288bda3, 32'hc371d124},
  {32'hc40c491e, 32'h42e80bfc, 32'h43ad3be5},
  {32'h450aad5a, 32'hc35fa79a, 32'h435b30a2},
  {32'hc4b1c576, 32'h437bf3e9, 32'hc237f498},
  {32'h436f7398, 32'hc401a775, 32'hc386b224},
  {32'hc3ccb2ad, 32'h420150d0, 32'hc3a0101f},
  {32'h441eb500, 32'h431796ca, 32'h43f22972},
  {32'hc4ebeb06, 32'h40982fff, 32'hc38c06b6},
  {32'h44cfea3c, 32'h424d831a, 32'h4370d782},
  {32'hc4fb4afd, 32'hc3948678, 32'h431152af},
  {32'h44959219, 32'hc2a0e6ff, 32'h4332f273},
  {32'h43020f08, 32'hc397566c, 32'hc38a9aba},
  {32'h44f18593, 32'h43c18654, 32'hc23f731e},
  {32'hc4f75bb9, 32'h43cdaa47, 32'hc235749c},
  {32'h43c5dd98, 32'h422e2c0b, 32'h43b3b8f5},
  {32'hc3822e70, 32'hc2ef9d24, 32'hc382dc7b},
  {32'h45185840, 32'h438e5746, 32'h439748a7},
  {32'hc49a55e3, 32'hc3563aa8, 32'hc36b3f51},
  {32'h45258316, 32'h439f2984, 32'h43a093a3},
  {32'h43809d50, 32'hc36c759d, 32'hc3bd0e1d},
  {32'h4503d9f6, 32'h41aea095, 32'hc4171f20},
  {32'hc42a8b46, 32'h43c85c22, 32'h43a033fb},
  {32'h439c7150, 32'h436430e2, 32'hc32302a3},
  {32'hc4e2241a, 32'h43a4ef23, 32'hc3d5e608},
  {32'h42a19eb0, 32'hc1f4bfb2, 32'h42d0c0f9},
  {32'hc50dc7f1, 32'hc2517e01, 32'h43c84298},
  {32'h44e16998, 32'h40dd1810, 32'hc377ebc8},
  {32'hc4e018e9, 32'h42f3b6af, 32'h43cdb06c},
  {32'h44ea4d68, 32'hc1ee9a71, 32'h4208721b},
  {32'hc31e90a0, 32'hc302c788, 32'hc3842247},
  {32'h450ee933, 32'h43087688, 32'h43199954},
  {32'hc4c1bbe4, 32'hc3c1e65c, 32'h4415b641},
  {32'h451588fe, 32'hc331d457, 32'hc3946902},
  {32'hc4b18fe8, 32'hc3615507, 32'h43644a29},
  {32'h44cb30a8, 32'hc38b721f, 32'hc3957b5e},
  {32'hc4eee670, 32'h422bd6ab, 32'hc303619c},
  {32'h44cacbc1, 32'hc23610de, 32'h42e3f4c1},
  {32'hc4dfb3e7, 32'hc1ab250e, 32'hc354cc1a},
  {32'h43868a57, 32'hc33ffd28, 32'hc146ab08},
  {32'hc43f4d77, 32'h430da317, 32'hc40ca35d},
  {32'h43d1f5c8, 32'hc29e83bd, 32'h43c1aaeb},
  {32'hc41d819d, 32'h42e42ceb, 32'hc38eaaa5},
  {32'h448f0e10, 32'hc35176e5, 32'hc3461426},
  {32'hc3df81d0, 32'h43e0a6ea, 32'hc324e93e},
  {32'h4351d0d5, 32'h42a6246e, 32'h4373bdf2},
  {32'hc4c6f3b2, 32'hc2ce0615, 32'hc3209fe0},
  {32'h446f6c2c, 32'hc23504d3, 32'h428460f8},
  {32'hc49610c0, 32'h42318d75, 32'h42e8f198},
  {32'h45054b09, 32'hc32dac54, 32'h42ca4bbe},
  {32'hc4a013b7, 32'h414bcc98, 32'hc265d7c1},
  {32'h450184cd, 32'h4388b21f, 32'h4389e816},
  {32'hc3c3fdaf, 32'hc3535178, 32'h42808fd7},
  {32'h43700d70, 32'h43864253, 32'h42e1d8aa},
  {32'hc3b30046, 32'h41e1aba1, 32'hc30078c3},
  {32'h4487f6e9, 32'h437fc23c, 32'h43372d9b},
  {32'hc4dfeb7e, 32'hc2e98165, 32'hc2ab272c},
  {32'h44d8c309, 32'h43e2dc6d, 32'h42b32c9a},
  {32'hc2ef1167, 32'h439b11fd, 32'hc316aac7},
  {32'h4422bc47, 32'h43010c85, 32'h43003149},
  {32'hc3a53230, 32'h4298a8d2, 32'hc38fd94e},
  {32'h44589505, 32'hc3415a07, 32'h430bd6d8},
  {32'hc4c306a5, 32'hc3bc3a05, 32'hc3969fa4},
  {32'h44d0e212, 32'h4351035a, 32'h43c60f76},
  {32'hc4982702, 32'hc283362b, 32'hc3567759},
  {32'h44f190a5, 32'h42c503e8, 32'hc3daab11},
  {32'hc4b9ecee, 32'hc30440a3, 32'hc3150dab},
  {32'h44ff4419, 32'h42c5dabb, 32'hc35b810a},
  {32'hc4ae4dc0, 32'h423fcdd0, 32'hc2dc4d12},
  {32'h444dbeb3, 32'hc1d5819a, 32'h430da36a},
  {32'hc502e461, 32'h42998255, 32'hc2632cf7},
  {32'hc49ebb25, 32'hc3af4c1a, 32'h43614369},
  {32'h44f5a5ad, 32'hc26f1e56, 32'hc198fbc7},
  {32'hc471a5a2, 32'h4296ad2e, 32'h424e381d},
  {32'h451764e3, 32'hc2133a1b, 32'h434bdcdc},
  {32'hc50f0b4e, 32'hc1da570a, 32'hc18314dc},
  {32'h43bed612, 32'hc34c0833, 32'hc23200d9},
  {32'hc36ce2d8, 32'hc3f74bab, 32'hc3d78b59},
  {32'h430df0fc, 32'h43569b88, 32'hc32f2d9f},
  {32'hc457d898, 32'hc2cb9423, 32'hc31bfed6},
  {32'h44936b0d, 32'hc33e3d3a, 32'hc2ecec60},
  {32'hc4024afa, 32'h4340417c, 32'hc38cee50},
  {32'h447a74bf, 32'hc38a0ed5, 32'h4340f847},
  {32'hc4ebe658, 32'h42570511, 32'hc2360540},
  {32'h44eab71b, 32'h43198124, 32'hc29904a6},
  {32'hc4af93eb, 32'h42a83a6a, 32'hc2924eb8},
  {32'h44d1757b, 32'h42bbf6f4, 32'hc1e4da96},
  {32'hc30a4750, 32'h428f7612, 32'hc333318c},
  {32'h44871171, 32'hc20121dc, 32'hc20bc08a},
  {32'hc4f73b0a, 32'h41d62585, 32'hc2e487ea},
  {32'h4509598c, 32'hc29b2000, 32'hc186750a},
  {32'hc4cb3c46, 32'hc367e185, 32'hc3cc8812},
  {32'h44fb184d, 32'hc3a0ee62, 32'h4262d7e4},
  {32'hc4a7931a, 32'h4179da94, 32'h41ccc288},
  {32'h441cf978, 32'h434d61fc, 32'h438519cd},
  {32'hc4621acc, 32'hc1be0fd0, 32'hc3848436},
  {32'h4474dda3, 32'hc39d2917, 32'hc3d08042},
  {32'hc4b4224e, 32'h434e0527, 32'h42f31ad4},
  {32'h44255b22, 32'h42c4d7ca, 32'h4392d4a2},
  {32'hc44decb6, 32'h4386c28e, 32'hc40e3c37},
  {32'h449ea81b, 32'hc2428845, 32'h42c5ace7},
  {32'hc4d07e6d, 32'hc2c058be, 32'h4275cb60},
  {32'h443420b9, 32'hc378ecb9, 32'h42a54094},
  {32'hc502f973, 32'hc3f6353a, 32'hc22cccce},
  {32'h44d04ac0, 32'hc3463a05, 32'h43867c26},
  {32'hc463342b, 32'h42e42a38, 32'hc2337112},
  {32'h44d07ba0, 32'h4387e545, 32'hc377fe53},
  {32'hc3e8a399, 32'hc30d97ea, 32'h4375928e},
  {32'hc2cb74a0, 32'h41f90459, 32'hc3d3247c},
  {32'hc50ce63d, 32'h435f4a25, 32'h42b079b9},
  {32'h446f4e44, 32'h438069de, 32'hc3a74553},
  {32'hc4757f7e, 32'hc2161b43, 32'h40d5e586},
  {32'h450a4ea3, 32'h43bb8ea4, 32'h41f45b7a},
  {32'hc3d25bc4, 32'hc38077fa, 32'hc3710521},
  {32'h44976150, 32'hc393203e, 32'h432c4054},
  {32'hc490d914, 32'h433f71fd, 32'h423d3399},
  {32'h4502d180, 32'hc125797a, 32'h43d87e1d},
  {32'hc50b0df1, 32'h43fd9a8a, 32'hc37dbf43},
  {32'h444a30ac, 32'hc2dd3963, 32'h42730126},
  {32'hc2f24b7c, 32'h42ac8e8a, 32'h41947125},
  {32'h44209b4a, 32'hc340b810, 32'hc31a61b4},
  {32'hc2ecb8a0, 32'hc367eff0, 32'hc10b06ba},
  {32'h45226b38, 32'h43122863, 32'hc23b1cd8},
  {32'hc41bdf60, 32'h43e096c1, 32'h438c8bdd},
  {32'h44c4d709, 32'hc3ef1337, 32'h421ca9c6},
  {32'hc467781e, 32'h42a7cd50, 32'hc2dc10dd},
  {32'h44e0dc25, 32'hc2328fe8, 32'hc2cd6a05},
  {32'hc40f765c, 32'h432ea0b6, 32'hc1f3f841},
  {32'h443b9588, 32'h42ae220e, 32'h430945aa},
  {32'hc4a6c35b, 32'hc0bbc0d8, 32'h42e38116},
  {32'h44b0693c, 32'hc39cc4c9, 32'h4282209b},
  {32'hc51f7128, 32'h439450da, 32'hc2cff660},
  {32'h44af7188, 32'hc390c8dd, 32'h4396040d},
  {32'hc37455d0, 32'hc3559d82, 32'h43162d41},
  {32'h44bec6cc, 32'h42f12dc7, 32'h43b93712},
  {32'hc417518b, 32'h43a9f667, 32'hc293cbfe},
  {32'h44f6e186, 32'h43f526f6, 32'hc181b650},
  {32'hc3ab2ea4, 32'h4200ab34, 32'hc2fbd0d3},
  {32'h44d8653b, 32'hc2e391df, 32'h419e8174},
  {32'hc3a49f78, 32'h44290049, 32'h4222b303},
  {32'h44a16874, 32'h43da7e42, 32'h4367c297},
  {32'hc4b3705a, 32'h43a0e471, 32'hc1e664d4},
  {32'h44ce2b56, 32'h431d1428, 32'hc2a37d81},
  {32'hc2b92434, 32'h42704d04, 32'h41416e12},
  {32'h4515dcdd, 32'h43b7465e, 32'h43a1211a},
  {32'hc4f871cb, 32'h42c6c78a, 32'h43d3ad1f},
  {32'h446d95ac, 32'h431162bc, 32'h4398fb8a},
  {32'hc3c6be94, 32'h43816612, 32'hc31b4885},
  {32'h44b07964, 32'h42ef5bde, 32'h434347fa},
  {32'hc3c464f8, 32'h4331ff0a, 32'h420f2595},
  {32'h4416a2f4, 32'h42fc8052, 32'hc2328388},
  {32'h439616a8, 32'hc32d6fe2, 32'hc324e45d},
  {32'h4441f072, 32'h4315a34d, 32'hc4004395},
  {32'hc4b34708, 32'h43c614d2, 32'hc2a9819b},
  {32'h44a2b466, 32'hc382f5b7, 32'h431f6672},
  {32'hc2124b00, 32'h43fdc75c, 32'h437705a7},
  {32'h4514a103, 32'hc376d582, 32'h4283fa67},
  {32'hc3409aa3, 32'hc31ee00b, 32'h4276ad66},
  {32'h45110ae8, 32'hc39d4088, 32'h42020ee1},
  {32'hc49bc475, 32'h436300a8, 32'h41a40c5b},
  {32'h44c20726, 32'hc337afaf, 32'hc3256417},
  {32'hc4f2dec2, 32'h43b11356, 32'h43968eb7},
  {32'h448e9c1c, 32'hc32b5640, 32'hc328ceb6},
  {32'hc5082aba, 32'hc203edf5, 32'h4311570d},
  {32'h44a33457, 32'h4382148c, 32'h42d6058f},
  {32'hc334ccb0, 32'h423e35f4, 32'h43b48af0},
  {32'h447c0dd8, 32'hc3acc5c7, 32'h41b232e6},
  {32'hc4c0c974, 32'hc30356f2, 32'h440584db},
  {32'h443b1a44, 32'hc3455ca4, 32'hc2a048e0},
  {32'hc3695f60, 32'h42a0cade, 32'hc3aa4962},
  {32'h451d19c6, 32'hc38ee075, 32'hc2767528},
  {32'hc48f25e7, 32'hc3ae387a, 32'h428fa1f0},
  {32'h43fb8bc6, 32'h43f0a256, 32'h432be2a9},
  {32'h426c4250, 32'h43382525, 32'h4320453a},
  {32'h44a43f96, 32'h42f0131e, 32'h43b42f00},
  {32'hc3712210, 32'h430b2d25, 32'hc28525c5},
  {32'h4407a20e, 32'hc3bb5c0c, 32'hc36e2b7c},
  {32'hc2d89c40, 32'hc3855de2, 32'h419fdac0},
  {32'h4432cc88, 32'hc3ec29db, 32'h421acb68},
  {32'hc4a6aead, 32'hbfbf6d14, 32'h43d1ab19},
  {32'h443a59be, 32'h4380f495, 32'hc32ae553},
  {32'hc434fd28, 32'h40cca27c, 32'hc2a82ce2},
  {32'h44dcbd40, 32'h4310c108, 32'hc185c24d},
  {32'hc43d8fd0, 32'h43724088, 32'h43bd4738},
  {32'h45029471, 32'hc2828cf6, 32'h4001ae6e},
  {32'hc48001ae, 32'h4408a4c9, 32'h43af688b},
  {32'h439a8a81, 32'h43ad80d6, 32'hc3e33e5d},
  {32'hc2eff560, 32'hc39ab49d, 32'hc2f199a4},
  {32'h443ccc8a, 32'hc2f6ea3a, 32'hc3241553},
  {32'hc4158ff8, 32'hc3150b57, 32'h431951a9},
  {32'h42064fe0, 32'hc199c445, 32'hc28eabec},
  {32'hc46e0e9c, 32'h42db1b03, 32'h4343b7d8},
  {32'h44277830, 32'h423b5dfc, 32'h43856220},
  {32'hc488b14c, 32'h428133e1, 32'h437a6dd6},
  {32'h4504a27c, 32'h41ce3bd0, 32'h435e4322},
  {32'hc4676652, 32'h4279f398, 32'h41d8ddc2},
  {32'h4512bb44, 32'hc282c28a, 32'h438ab38e},
  {32'hc51b92d7, 32'hc27d483a, 32'h4300e0af},
  {32'h438df554, 32'h42b8ed4f, 32'hc3676676},
  {32'hc3b6c7f8, 32'h43a4f910, 32'h42380a97},
  {32'h452574b2, 32'h43580172, 32'hc3107946},
  {32'hc3c2b028, 32'h43a74a9f, 32'h43afe2af},
  {32'h44780570, 32'hc0a6c105, 32'hc3433f44},
  {32'hc50c1504, 32'h41253a01, 32'h434b4a65},
  {32'h433fe3e8, 32'hc2a8a93a, 32'hc3b8dfe0},
  {32'hc474205c, 32'hc338363f, 32'h438e47d0},
  {32'h4465f326, 32'hc2e4c31e, 32'hc3883ac3},
  {32'hc5079723, 32'hc1ad6ea0, 32'hc3e7a370},
  {32'h44cc455e, 32'h430b2686, 32'h4121fdb8},
  {32'hc4ac2aae, 32'hc38e5f3b, 32'h436c2c84},
  {32'h4438042d, 32'hc333dd50, 32'h43462a0d},
  {32'hc4f8e21c, 32'h43918937, 32'h430443e6},
  {32'h44849d82, 32'hc37682e3, 32'h434c7610},
  {32'hc4808111, 32'hc350f71e, 32'h44013bb2},
  {32'h42d404b6, 32'hc3b5be3c, 32'h42af465d},
  {32'hc4b5a721, 32'h420928a5, 32'hc1ddc3cc},
  {32'h4309ca81, 32'h43613762, 32'hc3f6ed09},
  {32'hc5079d2c, 32'hc1f82ebb, 32'hbf777d60},
  {32'h4500a5f6, 32'hc3b1a8b5, 32'h43be51cb},
  {32'hc4534973, 32'hc3dc749d, 32'h440456a6},
  {32'h44c8007f, 32'h42c5ab22, 32'hc3a7e741},
  {32'h426e0900, 32'h438bd07c, 32'hc2296cc0},
  {32'h448c56c0, 32'h42798605, 32'hc19b08db},
  {32'hc4eacf86, 32'hc29ae14d, 32'h42c1961e},
  {32'h449eb786, 32'hc33dea20, 32'h439c0cc6},
  {32'hc3e74140, 32'h438e8be1, 32'h43f95284},
  {32'h449cfba5, 32'h42c6d34a, 32'hc3026f39},
  {32'hc3e94148, 32'h430cfed6, 32'h43c2d8ec},
  {32'h44cde0dd, 32'hc25a9c40, 32'h435f9612},
  {32'hc495e87f, 32'hc28b6740, 32'hc2bc09d2},
  {32'h44c72ab2, 32'h42b99052, 32'h439f514e},
  {32'h43b07378, 32'h43bba293, 32'h41d81669},
  {32'h442601d8, 32'h4300fd14, 32'hc355bba4},
  {32'hc4067026, 32'hc1da2869, 32'hc354dbf4},
  {32'h44397342, 32'h4248f6c7, 32'hc29596ca},
  {32'hc507eeb4, 32'h423d90fd, 32'hc32869b5},
  {32'h44586b94, 32'h431f1afe, 32'hc303a492},
  {32'hc43621f0, 32'h42a7ca5c, 32'hc22cab81},
  {32'h44d67fe0, 32'hc331157f, 32'hc331783e},
  {32'hc4ae801c, 32'h433ea401, 32'hc32915ca},
  {32'h44689943, 32'hc3fb8188, 32'h43b3456e},
  {32'hc4968cd3, 32'hc2dff9d5, 32'hc22f7a02},
  {32'h43f385f3, 32'hc2c3e5ed, 32'h3f8a43d4},
  {32'hc5072dbc, 32'hc308b52f, 32'h43bc3598},
  {32'h447a274d, 32'hc2b41563, 32'hc39f3a13},
  {32'hc49c34c7, 32'h433bc7b7, 32'hc3171dc6},
  {32'h450772cd, 32'hc2475cc1, 32'hc261a4cc},
  {32'hc41afa34, 32'h421e0b65, 32'hc38b8b68},
  {32'h444fb2cc, 32'hc305fe68, 32'hc253179e},
  {32'hc3c5ec60, 32'h436e2755, 32'h42c7d9e2},
  {32'h44cd171b, 32'hc2e72b73, 32'h43af499d},
  {32'hc24efc80, 32'h41ab1638, 32'h42f3f09a},
  {32'h440a6a3e, 32'h43746130, 32'h430e50c2},
  {32'hc341db65, 32'hc2d65223, 32'h439ff364},
  {32'h443543a2, 32'h4354ab86, 32'hc34d45c8},
  {32'hc4b51c66, 32'hc33e2dba, 32'hc2004165},
  {32'h45054846, 32'h413b5d7a, 32'h430ad650},
  {32'hc4f876c6, 32'hc2d0796d, 32'hc2ce5cfc},
  {32'h44d618ad, 32'h4386c94a, 32'h431e3ece},
  {32'hc4b154ba, 32'h41ba4627, 32'h4324dfb5},
  {32'h4526ee3e, 32'h42351a1b, 32'hc325c5b3},
  {32'hc4892559, 32'h43ea91a5, 32'h428c150e},
  {32'h448ddc6f, 32'hc36cd661, 32'hc28debf0},
  {32'hc1e39944, 32'hc36ba9b7, 32'hc299bd85},
  {32'h435c8530, 32'h43b83d82, 32'h4350dad2},
  {32'hc4fe46f7, 32'h43230b83, 32'hc3f427b7},
  {32'h449c6c4a, 32'h42e2b0e0, 32'h42e8346f},
  {32'hc4ebe680, 32'h4322cde8, 32'h4344ce49},
  {32'h4523469c, 32'hc31234ae, 32'h42e32172},
  {32'hc5232b7f, 32'h43c56c6f, 32'h440aba7a},
  {32'h446ab73e, 32'h43b7b87b, 32'h433a287c},
  {32'hc43462a7, 32'h43a4c653, 32'hc33fc0f9},
  {32'h43da1a70, 32'hc3a424c2, 32'hc392a279},
  {32'hc4e17a27, 32'h426893c2, 32'hc2c5b160},
  {32'h4481da28, 32'hc3278784, 32'hc3a3f8c0},
  {32'hc4b207c1, 32'h42178561, 32'h4413ea41},
  {32'h42efa0fa, 32'hc3adffab, 32'hc332bbd3},
  {32'hc5072438, 32'hc329f403, 32'h437f3838},
  {32'h44efc702, 32'h42d91905, 32'h43926bb6},
  {32'hc44c162a, 32'hc234543c, 32'hc3804a38},
  {32'h44d696b6, 32'hc3813c3a, 32'hc3eda858},
  {32'hc44a7db0, 32'h43040c28, 32'h431aaa46},
  {32'h44d7d0e6, 32'h423badde, 32'hc4203885},
  {32'hc4443bd0, 32'hc2627ea4, 32'hc0e4abea},
  {32'h44d754b4, 32'hc37f9c36, 32'h42ca1fa6},
  {32'hc507cb19, 32'h43353bf8, 32'h44061bf0},
  {32'h433818b8, 32'h42cf6908, 32'h434a2c58},
  {32'hc4cfb7a4, 32'hc3ab9901, 32'hc258321e},
  {32'h44f63590, 32'h426f7617, 32'hc2063f44},
  {32'hc4fda3b2, 32'hc40ae697, 32'h43767d48},
  {32'h449367e9, 32'hc2f6d977, 32'hc38d7d39},
  {32'hc4273748, 32'hc38a8d3a, 32'hc35174f3},
  {32'h44b17380, 32'hc3958a8e, 32'hc334e96b},
  {32'hc4f11408, 32'hc38fd096, 32'h42b421b3},
  {32'h43074bb0, 32'hc3251097, 32'hc359395a},
  {32'hc4d4993a, 32'h42b21935, 32'h437f5f9d},
  {32'h4510ae16, 32'hc36ef403, 32'hc2f9bbe6},
  {32'hc4f4a00a, 32'h43dc5c85, 32'hc0e28353},
  {32'h449c0fc7, 32'hc38e09c3, 32'hc38585c7},
  {32'hc40e13de, 32'h4300832c, 32'h436af8e5},
  {32'h4486e2fe, 32'hc3b174e5, 32'h4328ef3c},
  {32'hc44da112, 32'hc2939dd2, 32'h4157f661},
  {32'h448bb250, 32'h433b8972, 32'hc30bc245},
  {32'hc33d34e0, 32'hc21fae4f, 32'hc22ed72b},
  {32'h4307dbb8, 32'hc1e930f3, 32'hc11a2a0b},
  {32'hc4f88cbc, 32'hc2a3bd68, 32'hc38b5e06},
  {32'h44f4e1da, 32'hc3084059, 32'hc265bc2a},
  {32'hc4ee3c12, 32'h430d0b48, 32'hc31163e8},
  {32'h445180ed, 32'hc4123266, 32'h43090fa9},
  {32'hc4761678, 32'h42a13bfe, 32'h43a8f1fc},
  {32'h450492d2, 32'h410ac0ce, 32'hc2adec2e},
  {32'hc4ef2546, 32'hbfb7ca80, 32'h423d9fba},
  {32'h44fd44de, 32'hc3747a4e, 32'h42e10d00},
  {32'hc4d6dc58, 32'h41d71549, 32'h42748d30},
  {32'h448e5a33, 32'hc3c1d711, 32'h434517f1},
  {32'hc3c3dddf, 32'hc36f553a, 32'h43731dbd},
  {32'h431574cc, 32'hc388ba1e, 32'h4314c4a4},
  {32'hc40845d8, 32'h43b85f22, 32'h423301d3},
  {32'h442794fe, 32'hc3bd969e, 32'h42b04a77},
  {32'hc40938fd, 32'h4300b9d8, 32'hc2e102ea},
  {32'h43a1d28a, 32'hc4425a72, 32'h42f6e5f1},
  {32'hc4d976ca, 32'h43a4f926, 32'hc32209bf},
  {32'h449418bf, 32'hc3359895, 32'hc2786e06},
  {32'hc28f7770, 32'hc3191452, 32'hc2db0482},
  {32'h44f63ff8, 32'h41da0bf8, 32'hc274f57b},
  {32'hc38055f8, 32'hc356c0c1, 32'hc3b43552},
  {32'h4490141a, 32'hc3efd2f1, 32'h42b7a6fc},
  {32'hc42ece80, 32'h4394ea62, 32'h41141c8a},
  {32'h446a184a, 32'h4343a8c9, 32'h42a32577},
  {32'hc5057d0f, 32'hc3831c75, 32'hc42c5296},
  {32'h448e0209, 32'h436c02e5, 32'hc3a8c9e0},
  {32'hc508f5da, 32'h43d85077, 32'h438cba9c},
  {32'h45006d8d, 32'hc0bd3736, 32'h4103f146},
  {32'h424bb180, 32'hc29895f9, 32'hc33a3458},
  {32'h44e22312, 32'h42fcc2e5, 32'hc3e57bce},
  {32'hc387bfb8, 32'hc3a5cc3a, 32'hc35d44ec},
  {32'h44a072d9, 32'hc2d18f46, 32'h41fb0dc4},
  {32'hc4c16dde, 32'hc38f279c, 32'h428d2eeb},
  {32'h44820946, 32'h43531962, 32'hc20d1b59},
  {32'hc4c044b4, 32'hc33c8e6a, 32'hc33e2e31},
  {32'h44d7226c, 32'hc3c6ef2c, 32'hc39d18a0},
  {32'hc50fc001, 32'hc38c3768, 32'h43b7cfb3},
  {32'h450b7c34, 32'hc3940c18, 32'hc233d7fa},
  {32'hc4a015e9, 32'hc3ae8ba2, 32'hc30a8194},
  {32'h443bde40, 32'h43ab1bf1, 32'hc0659e5a},
  {32'hc4bc4350, 32'h41d2dc10, 32'hc3efa76d},
  {32'h4513aac9, 32'hc3d69ec0, 32'h43219a14},
  {32'hc50885d8, 32'hc33be5ad, 32'hc253c424},
  {32'h44201783, 32'h4379256b, 32'h432dbc07},
  {32'hc487ff61, 32'h4043df03, 32'hc3b310da},
  {32'h443034d4, 32'h432eedf1, 32'h43bca090},
  {32'hc507a0c7, 32'h428419d6, 32'hc1aff618},
  {32'h4359b8b8, 32'h431bba3a, 32'hc37c5627},
  {32'hc4ec064a, 32'h4241937f, 32'hc2ac7ad9},
  {32'h44cf674d, 32'hc17185e6, 32'hc2b5c394},
  {32'hc452b035, 32'h437ba377, 32'h43b6b64c},
  {32'h4365baaa, 32'h427df567, 32'h435fe855},
  {32'hc47e1633, 32'hc307d085, 32'hc37af788},
  {32'h44ff29bc, 32'hc2a31267, 32'hc1a21918},
  {32'hc49e61a9, 32'hc394c331, 32'h42683399},
  {32'h43570444, 32'h43fff3e6, 32'hc2b84f50},
  {32'hc49ad561, 32'h4219d835, 32'hc268cd51},
  {32'h44713e52, 32'hc268d602, 32'h40e2fc22},
  {32'hc4af8df3, 32'h438ba3cc, 32'h43247714},
  {32'h44f97730, 32'h4234ae55, 32'hc1abadad},
  {32'hc2728090, 32'hc2970f46, 32'hc3a8e82f},
  {32'h442166e2, 32'hc3a4b992, 32'hc3133995},
  {32'hc447eef3, 32'h434c007c, 32'hc28279d6},
  {32'h4458aac2, 32'hc1c01233, 32'h432be230},
  {32'hc4bcb3ac, 32'h425d954d, 32'h422d8493},
  {32'h43e9df94, 32'h428f04a5, 32'hc1f1ae83},
  {32'hc495fb5f, 32'hc23a8bce, 32'h42c31db7},
  {32'h442212ae, 32'h43a71a18, 32'h4368e801},
  {32'hc4d06052, 32'h438f555c, 32'h4409297b},
  {32'h4516d44f, 32'hc2a2f70b, 32'hc2b7595e},
  {32'hc5007ca4, 32'hc24218a0, 32'h42488972},
  {32'h44c4b948, 32'hc323065e, 32'hc32ab35c},
  {32'h42a6ed60, 32'hc3143c91, 32'hc2972588},
  {32'h44055c52, 32'h421a847b, 32'hc2c15575},
  {32'hc501574b, 32'hc2c18316, 32'h42cc73fe},
  {32'h44bb96b0, 32'hc38525ca, 32'h435b36b2},
  {32'hc49705a3, 32'hc2c12aa5, 32'hc2ac68c8},
  {32'h4353dd8c, 32'hc332e488, 32'hc3911b7a},
  {32'hc4d0e7e9, 32'hc38a47b5, 32'h43cbbd84},
  {32'h4503606a, 32'hc2ead528, 32'hc216ccfe},
  {32'hc4b5be9d, 32'h4242ed1e, 32'hc2cf483c},
  {32'h44c7b91b, 32'h431887c6, 32'hc319fcf3},
  {32'hc4952fe4, 32'h439985b9, 32'hc33887b5},
  {32'h44d8983f, 32'hc3247381, 32'hc3954934},
  {32'h42a98472, 32'h42f74048, 32'hc3b122c0},
  {32'h4508f281, 32'hc31ccd4c, 32'hc3164f67},
  {32'hc481d44b, 32'h43504fb0, 32'h41cd404c},
  {32'h44c4995a, 32'hc39b3ef6, 32'hc353cc16},
  {32'hc4ac7106, 32'h42c04a36, 32'hc383195b},
  {32'h44c02b08, 32'hc35bf912, 32'h435270f2},
  {32'hc50b69ee, 32'h434b7fb1, 32'h421fbb57},
  {32'h44d389bc, 32'h439bd4af, 32'hc32fee44},
  {32'hc4a9964f, 32'h41d8a775, 32'h43495b41},
  {32'h44053532, 32'hc3828b4d, 32'hc146ccee},
  {32'hc2d60da0, 32'h429860d5, 32'h438b1c32},
  {32'h4488b7b0, 32'hc315a094, 32'h43103af3},
  {32'hc5109330, 32'h41ed8e89, 32'h422a375b},
  {32'h44537e00, 32'h420588b2, 32'h44059c57},
  {32'hc49ccf0c, 32'h441df97f, 32'h420926b6},
  {32'h450f229a, 32'h433e62c3, 32'hc365e37b},
  {32'hc4eee044, 32'h437c85fe, 32'hc30c4f8b},
  {32'h43497ac0, 32'hc30cb230, 32'hc39286f5},
  {32'hc4a964e4, 32'hc34682a5, 32'h4315815f},
  {32'h4449e2f9, 32'hc32caa19, 32'hc2cfc933},
  {32'hc4157cb7, 32'hc15bbc1f, 32'h40a1ab9b},
  {32'h45147b1c, 32'hc24f19a1, 32'h43210e05},
  {32'hc514a101, 32'hc38d1c3c, 32'h439f4a6a},
  {32'h44f8633a, 32'hc2808d5c, 32'h435be349},
  {32'hc5056a91, 32'hc2900bab, 32'h43960d15},
  {32'h44ab86be, 32'h43428b82, 32'hc3226658},
  {32'hc4b8c7b1, 32'h435efe10, 32'h43645ad8},
  {32'h443b2708, 32'h4376248d, 32'h41a3a22e},
  {32'hc4b10abc, 32'h43922707, 32'h42ee9ca5},
  {32'h45032e73, 32'h42871674, 32'hc16f1d32},
  {32'hc4807862, 32'h423aa5bf, 32'hc38c8fde},
  {32'h45038f45, 32'hc2b8e751, 32'hc286d6ca},
  {32'hc44b3cdc, 32'hc2d0c457, 32'h431ddb1b},
  {32'h43e0300a, 32'hc2a62c84, 32'h421d4c84},
  {32'hc47ff3ac, 32'h43c1ca1f, 32'h43091d47},
  {32'h42cf23fe, 32'h437daa5d, 32'h429155cd},
  {32'hc3b47460, 32'h4346f2a0, 32'h40844500},
  {32'h44f34088, 32'hc39bf67b, 32'h43309859},
  {32'hc4a19867, 32'h43d4f30e, 32'h430081a1},
  {32'h44937be9, 32'h434742fb, 32'h41f8a12d},
  {32'hc4daa220, 32'hc30d3dea, 32'hc32803ef},
  {32'h44fd2743, 32'hc2610b46, 32'h43107541},
  {32'h4226b500, 32'h420dbae3, 32'h43127d00},
  {32'h45236d96, 32'hc3acaf7a, 32'hc3d9d503},
  {32'hc23fa6c0, 32'hc2b5b082, 32'hc3e590a2},
  {32'h44c3a57f, 32'h42381ff7, 32'h43eb5f1b},
  {32'hc3cb7d96, 32'hc37af849, 32'hc1d605a8},
  {32'h4409a150, 32'h3fc13a84, 32'hc316927e},
  {32'hc4358a02, 32'hc3996211, 32'h4415c9f6},
  {32'h441de63c, 32'h4380c362, 32'hc3d52e2b},
  {32'hc5059d49, 32'hc32a56d3, 32'h431779b7},
  {32'hc3163100, 32'hc36cec65, 32'hc3a0e09c},
  {32'hc487e5e8, 32'h42f346f7, 32'h43a999a4},
  {32'h44dd0964, 32'hc22dccf7, 32'h43429fd1},
  {32'hc34e1e43, 32'h42ee0324, 32'h423e357b},
  {32'h443e2170, 32'hc39d51e1, 32'hc2ddcecc},
  {32'hc504a00d, 32'hc326219e, 32'h4351ca30},
  {32'h450b0b24, 32'hc333c3a8, 32'h42df7b41},
  {32'hc5116890, 32'h434779a7, 32'hc14c4b36},
  {32'h44aef704, 32'h431b01aa, 32'hc38169d9},
  {32'hc386b25c, 32'h43aa984e, 32'h41248819},
  {32'h447679fe, 32'hc306c152, 32'hc2b822b1},
  {32'hc4d7ee01, 32'h43342882, 32'h4312d0fe},
  {32'h44b7d53a, 32'hc30f139a, 32'h437e48f4},
  {32'hc51893b3, 32'hc38824e2, 32'hc36d6b16},
  {32'h450b76ff, 32'h42ecde8c, 32'h42f29b7d},
  {32'hc4a262e6, 32'h3f8ea97a, 32'h43847cd1},
  {32'h4461a32a, 32'hc39fbdbd, 32'hc36dd733},
  {32'hc4d75927, 32'hc3384fd9, 32'h43ba462f},
  {32'h44e54c70, 32'hc244da8a, 32'h43a186d3},
  {32'hc4a49076, 32'h43eb2f2b, 32'h43d728b2},
  {32'h451f2e9d, 32'h429b025a, 32'hc305edeb},
  {32'hc2c35980, 32'hc3223855, 32'h40610f00},
  {32'h446a1743, 32'hc24cbcd5, 32'hc35eac5b},
  {32'hc4d90f0a, 32'h438e0da4, 32'h41e58549},
  {32'h44d7a241, 32'hc3b6493a, 32'hc2801144},
  {32'hc4c712fe, 32'h42c9f82c, 32'h442d5f2a},
  {32'h44a1ac4a, 32'hc320dc8b, 32'hc287375c},
  {32'hc444407a, 32'h4383a0b4, 32'h436886c4},
  {32'h44d3d4b0, 32'h43ab2d2d, 32'hc30e6539},
  {32'hc3af38e0, 32'h436ae880, 32'h420b7dfe},
  {32'h45001a3d, 32'hc25446a6, 32'hc32c5edc},
  {32'hc4c3982e, 32'hc203e626, 32'hc28bc0f7},
  {32'h4521c35f, 32'hc265afdc, 32'hc3311296},
  {32'hc5122871, 32'h402d8e72, 32'hc2506c90},
  {32'h43e9ae04, 32'hc2de70c7, 32'h4401179e},
  {32'hc4de2b67, 32'hc3993596, 32'h41d391e0},
  {32'h44a31d8e, 32'hc3183c90, 32'h440311ba},
  {32'hc4151082, 32'h4307e955, 32'h430b598e},
  {32'h44ac6722, 32'hc40ef7f5, 32'hc3a1196f},
  {32'hc3ab542c, 32'h4342bdc2, 32'hc22c05ac},
  {32'h44338e72, 32'h433a98ed, 32'hc3972546},
  {32'hc4f62298, 32'hc3505120, 32'hc396a466},
  {32'h43851e7c, 32'h42d4bcfd, 32'h4315dc2f},
  {32'hc4ac78f0, 32'h43855edc, 32'hc2b381b7},
  {32'h44aa24d6, 32'h434158a3, 32'hc274f464},
  {32'hc413a666, 32'h4363c50f, 32'h43ce6625},
  {32'h44f34a71, 32'h42778a6d, 32'hc20527aa},
  {32'hc498802f, 32'hc358831b, 32'h43eaf254},
  {32'h43bdb2ea, 32'h42afbeab, 32'hc31320b2},
  {32'hc4e8c82a, 32'h439daf92, 32'hc32d3215},
  {32'h4428b906, 32'hc04bab8c, 32'hc356b8c2},
  {32'hc4ad6c2e, 32'hc30ce113, 32'hc3c4de45},
  {32'h44aa6a62, 32'hc292234a, 32'hc1e20163},
  {32'hc45e6db8, 32'hc2f7ce2a, 32'h4382ac56},
  {32'h442c22f8, 32'hc29fb5df, 32'hc38f795f},
  {32'hc2b35886, 32'hc337c6c7, 32'hc38229cc},
  {32'h44dc28d9, 32'hc316ba84, 32'hc2b4d01d},
  {32'hc4d035c3, 32'h422b3b00, 32'h435c7913},
  {32'h43d9472d, 32'hc1ceb15d, 32'hc3420527},
  {32'hc4e4a5f4, 32'hc18a9dc9, 32'hc28967fd},
  {32'h44a31f5e, 32'h43dc1591, 32'hc3920895},
  {32'hc43b4cd8, 32'h42dff478, 32'hc04547bf},
  {32'h44b555a8, 32'hc356a2a6, 32'h426a67ba},
  {32'h44e5e7f2, 32'h4348aa14, 32'hc0e0f200},
  {32'hc3c6e1c3, 32'h4335e3ca, 32'hc22100a6},
  {32'h438b51f4, 32'h43be84ee, 32'h420f1a7f},
  {32'hc49f833e, 32'hc22bdb6c, 32'h432f96e3},
  {32'h43e75307, 32'hc2dbf4d7, 32'hc3c80012},
  {32'hc40a33ea, 32'h43ac0c82, 32'h4342dfcc},
  {32'h44fcfb5a, 32'hc214e133, 32'h4323cf38},
  {32'hc4833446, 32'hc37d8144, 32'h43386aab},
  {32'h44556360, 32'hc1ad9d88, 32'hc3312daa},
  {32'hc3de2e24, 32'h432a5b7f, 32'hc3153f06},
  {32'h44e9d77a, 32'h434a1477, 32'hc11032ce},
  {32'hc51ca823, 32'hc34732dc, 32'hc2d526db},
  {32'h42dd6ff0, 32'hc2f6f710, 32'h4336cdf4},
  {32'hc31ed32c, 32'h43207ead, 32'hc33d3e2a},
  {32'h450af413, 32'h4334e3c2, 32'h43438a43},
  {32'hc2f3b7e0, 32'hc3b4a4cd, 32'h430ecf31},
  {32'h451360d3, 32'h439708f6, 32'hc322b5df},
  {32'hc25b4dc0, 32'hc32e0b98, 32'hc19395f6},
  {32'h44dbb104, 32'h42317b75, 32'h43429f02},
  {32'hc4ec0347, 32'h43a55b34, 32'hc363d193},
  {32'h439f8c44, 32'h4365a394, 32'hc3c0176a},
  {32'hc49ba15c, 32'hc32d4921, 32'h42309bbb},
  {32'h44bce7ec, 32'h429ab9fd, 32'hc2aa8657},
  {32'hc5109a35, 32'hc2b3531b, 32'h42d65d7c},
  {32'h43b8c9ad, 32'h42db0df5, 32'hc330ac55},
  {32'hc503098a, 32'hc1229036, 32'h438baee6},
  {32'h433bd2f0, 32'h4334de1c, 32'hc344a55d},
  {32'hc4df21e5, 32'h42f66a65, 32'hc1fa328f},
  {32'h44edd01b, 32'h43139a78, 32'h42154244},
  {32'hc3a0db94, 32'h4342fc02, 32'hc31e454b},
  {32'h450f00c3, 32'h424c8274, 32'hc38af17d},
  {32'hc23deb6a, 32'hc2c256b7, 32'h42539f77},
  {32'h4439aa3d, 32'h42bca9da, 32'hc35afa36},
  {32'hc4e213a1, 32'h43256390, 32'hc2a90f90},
  {32'h44769da2, 32'h43ca1fbc, 32'hc34fe18b},
  {32'hc4bfe098, 32'hc36d4b61, 32'hc29fd68e},
  {32'h43275f08, 32'h4308e0c9, 32'hc36cb2c2},
  {32'hc5008e6e, 32'h441bca0b, 32'hc38391fa},
  {32'h4510883e, 32'h425063dd, 32'hc392659a},
  {32'h42de39f0, 32'hc2e185b2, 32'h440dffca},
  {32'h440cf294, 32'hc35fb7fd, 32'hc3a64eb0},
  {32'hc503c512, 32'h4393eee3, 32'hc39dc7a8},
  {32'hc3219850, 32'h41d708ea, 32'h43a197ed},
  {32'hc47ee693, 32'h4224a132, 32'h432de878},
  {32'h44899bed, 32'h433ab4e8, 32'hc28b4d60},
  {32'hc3927390, 32'hc342d85d, 32'hc2908b04},
  {32'h42c1aea0, 32'hc2c89b0b, 32'h4382bd68},
  {32'hc4ecd7f6, 32'h419189c7, 32'hc3ad7ecc},
  {32'h4403c1e9, 32'h4394a039, 32'hc323d77c},
  {32'hc42e2485, 32'hc2617b0c, 32'h41cda410},
  {32'h419a58c5, 32'h42ed06b1, 32'hc329a498},
  {32'hc388b55d, 32'hc2285a3f, 32'h43b7062e},
  {32'h43da2cd4, 32'hc29870cb, 32'hc327dd1b},
  {32'hc4ba700b, 32'hc2b4d65c, 32'h42f1387f},
  {32'h448c96a3, 32'h43d2fb84, 32'hc36212ab},
  {32'hc4ecd4a6, 32'h42243924, 32'hc339fc0c},
  {32'h447c63ac, 32'hc1cd78fa, 32'h432f44cb},
  {32'h42108176, 32'hc39e237b, 32'h40325d85},
  {32'h4490c4d1, 32'h42107a58, 32'h421d566e},
  {32'hc4841f34, 32'h43c55f4f, 32'hc2d3b546},
  {32'h4512d016, 32'hc361e5de, 32'hc19d1e9b},
  {32'hc4afe45e, 32'hc226c920, 32'hc3674f6a},
  {32'hc321532a, 32'h424e8423, 32'hc320828a},
  {32'hc506a67c, 32'h43838f40, 32'h4323435a},
  {32'h448cd108, 32'h438de409, 32'hc31b0930},
  {32'hc3ad9b90, 32'h42f40729, 32'h416d61ce},
  {32'h44916ce8, 32'h438c8c7b, 32'h432f4ff8},
  {32'hc4324006, 32'hc311f122, 32'hc32a4abc},
  {32'h44c38979, 32'h42bcf061, 32'h416f646c},
  {32'hc42cc74f, 32'hc2aff040, 32'hc33a5ede},
  {32'h44ad5f78, 32'hc21eaf2d, 32'h43d02528},
  {32'hc48e312f, 32'hc33c6062, 32'hc1537e2e},
  {32'h44c9ed97, 32'h439e6839, 32'hc1b5c16a},
  {32'hc3504860, 32'h4302d886, 32'hc299607b},
  {32'h44ea5e9a, 32'h4367cbc9, 32'h42993428},
  {32'hc3d8c166, 32'h44000b99, 32'h42f7d2b1},
  {32'h44a8e878, 32'h423c1a9e, 32'hc2d64d80},
  {32'hc5035bc2, 32'h43a5cea5, 32'h42ab5687},
  {32'h4509b813, 32'hc3b704ea, 32'h43a1246c},
  {32'hc4bfd86c, 32'hc39dc214, 32'h430e78ef},
  {32'hc310c560, 32'hc352cbc9, 32'hc169d82c},
  {32'hc4d1f66a, 32'h42228f66, 32'h4396ba53},
  {32'h44bb7218, 32'h44123099, 32'h439c0692},
  {32'hc411d2fc, 32'hc0f8e536, 32'hc3b3f11a},
  {32'h450a2880, 32'hc3cbb568, 32'hc2e7d540},
  {32'hc4236cf6, 32'hc284b5d2, 32'h429f164f},
  {32'h44db031c, 32'h43a308d1, 32'hc408512e},
  {32'hc50bf6f9, 32'h431dfe16, 32'hc3888e52},
  {32'h44a0e2aa, 32'hc11097a4, 32'h42b4a44e},
  {32'hc3894b6a, 32'hc3b0826d, 32'h43c30664},
  {32'h44c4e0f9, 32'h436269be, 32'hc397bf15},
  {32'hc481cbad, 32'hc3e1c831, 32'h42b7266b},
  {32'h4501869d, 32'hc2b3cc78, 32'h429ab9fa},
  {32'hc4c4638b, 32'hc2511395, 32'hc2a1b18a},
  {32'h44dfd00f, 32'h428de94f, 32'hc2b3ce82},
  {32'hc3ff54c8, 32'h41c5f097, 32'h42c89394},
  {32'h44188092, 32'h4183e62e, 32'h43832120},
  {32'hc4091193, 32'h4250cecb, 32'hc3a53773},
  {32'h44bbe53a, 32'h43d2e36d, 32'h4225b7f8},
  {32'hc3dd5753, 32'hc38ec71b, 32'h432b84df},
  {32'h44c00dbb, 32'h4393a98c, 32'hc2bf7375},
  {32'hc4d3efd3, 32'h41a40626, 32'h43a2baea},
  {32'h4455d371, 32'h427eda62, 32'h423d35cd},
  {32'hc4fe716d, 32'h43ac82ab, 32'h41109271},
  {32'h44b16b8a, 32'hc380aa2b, 32'hc28ca107},
  {32'hc4723dfd, 32'hc2d430ea, 32'h4165f364},
  {32'h45044f91, 32'hc24200a8, 32'hc274a3d8},
  {32'hc4b0facc, 32'hc252ecc4, 32'hc28ba400},
  {32'h442a043d, 32'h434419e4, 32'hc2efd5ee},
  {32'hc4c0a097, 32'hc4087156, 32'h41a32b36},
  {32'h44b30515, 32'h42a52a4c, 32'hc23cb54f},
  {32'hc32f3974, 32'h43d3331d, 32'h439da833},
  {32'h438d5e98, 32'h43927ef0, 32'h40a6ae90},
  {32'hc4c6f8e2, 32'h4382dccf, 32'hc30f00d1},
  {32'h4504cb55, 32'h4317c8f8, 32'hc10282b0},
  {32'hc481a196, 32'hc2864b8d, 32'h3f394a38},
  {32'h43b03140, 32'hc38143a5, 32'hc28c3fd6},
  {32'hc4e130f1, 32'h42daa3d4, 32'h438519a6},
  {32'h448519fe, 32'h41f01ae8, 32'hc26983f0},
  {32'hc4ee7eb6, 32'hc2754898, 32'hc3c3933f},
  {32'h44ed8e66, 32'hc2f1f9f1, 32'h4356cc87},
  {32'hc43c0c2e, 32'hc29569cd, 32'h4340c960},
  {32'h45032275, 32'h426e44af, 32'hc207eced},
  {32'hc38ab6dd, 32'h42719ec1, 32'h423c3c1e},
  {32'h44895cac, 32'hc3dbb764, 32'h438a9091},
  {32'hc42ca654, 32'hc4125632, 32'hc39eac02},
  {32'h4440389b, 32'hc41512ac, 32'h43abd3c2},
  {32'hc4cae263, 32'h434d7902, 32'hc2de8caa},
  {32'h44eaf206, 32'hc2d98582, 32'h429d5bfa},
  {32'hc34d309e, 32'h439a9b92, 32'hc2c792ea},
  {32'h43def7de, 32'hc3b84a39, 32'hc3826c82},
  {32'hc471bfa3, 32'h43ae03ac, 32'hc3de89b5},
  {32'h44cc1b2e, 32'h4152fa68, 32'hc25151d5},
  {32'hc40f7a69, 32'hc222cdaa, 32'hc29c2d2e},
  {32'h43974978, 32'h43cb8952, 32'hc335e157},
  {32'hc2c05f48, 32'hc31cc9d4, 32'h430fd226},
  {32'h44a53e51, 32'h432c9513, 32'hc18ea8ed},
  {32'hc4122d40, 32'h41ae235e, 32'hc3d82405},
  {32'h4497257b, 32'h4353e6ec, 32'hc3a633b4},
  {32'hc4e51144, 32'h439c24f3, 32'h4394fd5a},
  {32'h44ed0c51, 32'h43dc5bc6, 32'hc2835c38},
  {32'hc425a17a, 32'hc221307d, 32'hc31d1392},
  {32'h44a36208, 32'h43c91b0d, 32'h4230e903},
  {32'h438063a0, 32'hc28e3ea7, 32'h4334c690},
  {32'h44d8a95f, 32'h43512217, 32'hc135ee6a},
  {32'hc506858f, 32'h42a1ff31, 32'hc3380f9b},
  {32'h44d5cb43, 32'h430a1c1c, 32'hc28bb48d},
  {32'hc4f6ec83, 32'hc33bfef7, 32'hc2a247ec},
  {32'h44599cea, 32'hc3971cbb, 32'h430eb177},
  {32'hc50bb9e7, 32'h429ba6f3, 32'hc30a6956},
  {32'h4488d659, 32'h4345f480, 32'hc29a9eac},
  {32'hc4d3bf6a, 32'h43d6ab59, 32'hc023d66a},
  {32'h42947c08, 32'h428967d8, 32'h4293ed95},
  {32'hc4e1e7dd, 32'hc3007e25, 32'h43b75614},
  {32'h44b071b1, 32'hc36a1310, 32'hc3007c41},
  {32'hc43ace1e, 32'hbf6be840, 32'hc31f5567},
  {32'h437f074c, 32'hc3d5cb61, 32'h439f3161},
  {32'hc4013100, 32'hc20ba11f, 32'hc3bc902f},
  {32'h43e8a1e8, 32'h427dca7d, 32'h431d8c97},
  {32'hc48c7900, 32'hc29445f0, 32'hc33b2255},
  {32'h43e0686b, 32'hc304865b, 32'h439b366c},
  {32'hc4e2063f, 32'h41beccb1, 32'hc30efc47},
  {32'h44ee77d4, 32'h4379499d, 32'h42d9515f},
  {32'hc33c598b, 32'hc39540e5, 32'hc32bb9b1},
  {32'h44ff94cc, 32'hc23e88ae, 32'hc25448db},
  {32'hc48815d0, 32'hc310813e, 32'hc38109c6},
  {32'h4458186e, 32'h429488f3, 32'hc21d6e8c},
  {32'hc4247560, 32'hc311ed32, 32'h436783c2},
  {32'h44fce2da, 32'hc31520c0, 32'h42c53a9b},
  {32'hc37713cc, 32'hc349f71a, 32'h416e2bf4},
  {32'h443595e8, 32'hc362e634, 32'hc2208bd7},
  {32'hc4bc3ac3, 32'h4397cc97, 32'h43844e12},
  {32'h448a583b, 32'h436311b0, 32'hc3c69d17},
  {32'hc3417876, 32'hc3482a67, 32'hc39588a1},
  {32'h449bdfe6, 32'h4380ea30, 32'h42e60fff},
  {32'hc4eafc68, 32'h4396e5f5, 32'hc3370cd4},
  {32'h4463ed27, 32'hc308b0d1, 32'h422e4022},
  {32'h42f723e0, 32'hc33a4339, 32'h42c672d2},
  {32'h4325e348, 32'hc2b64304, 32'h444637b2},
  {32'hc4a6d25d, 32'hc297d241, 32'h4333a617},
  {32'h44d17b48, 32'h420c3ffb, 32'h42268e07},
  {32'hc3eaab3c, 32'hc3954429, 32'h43151d8e},
  {32'h44d7b460, 32'hc37d948e, 32'h42bfcf4f},
  {32'hc508deb9, 32'hc38c5398, 32'h4205edba},
  {32'h44ccbe3b, 32'hc3114a13, 32'hc2bb9776},
  {32'h43e93be8, 32'h429f4736, 32'h428993aa},
  {32'h43c90f4f, 32'h4321470a, 32'h420e4638},
  {32'hc4bd375e, 32'hc29fce28, 32'hc3a7a082},
  {32'hc36763b0, 32'hc343968a, 32'hc2c22bc0},
  {32'hc4db0770, 32'h42fee930, 32'h43b5a855},
  {32'h450d8b1a, 32'h4360f942, 32'h43a85e3f},
  {32'hc4bc27c2, 32'h41a34e0d, 32'h41bc521a},
  {32'h44dbf3db, 32'hc2dcc831, 32'h4294ac71},
  {32'hc415b95e, 32'h4198c258, 32'h43550f18},
  {32'h451cec38, 32'hc3486fd8, 32'h43cc8044},
  {32'hc410018e, 32'hc32bb5db, 32'h4335e0a3},
  {32'h44fe99ba, 32'h41e3f3a1, 32'hc388a96c},
  {32'hc4a9a6f6, 32'hc3851789, 32'h43be7187},
  {32'h43c5a638, 32'hc38a6e35, 32'h43b3adcf},
  {32'hc42d76c8, 32'hc3c16884, 32'h43c3cea4},
  {32'h44d05b50, 32'hc31dd3a5, 32'h41e24bba},
  {32'hc3da5b72, 32'h430ef0cd, 32'hc26f3913},
  {32'h44a4d6ce, 32'h434249b2, 32'h42ad0067},
  {32'hc2a5e5a0, 32'h4365d4cb, 32'h43507657},
  {32'h4515f887, 32'hc29d972d, 32'h43b09298},
  {32'hc4df0930, 32'hc2dc6014, 32'hc39c9a08},
  {32'h445bd3b0, 32'h43933e82, 32'h424b5c1a},
  {32'hc39bfe3d, 32'h433d0fce, 32'hc38393f9},
  {32'h44982e80, 32'hc3cf48f0, 32'h4389b6d4},
  {32'hc4dcc74f, 32'hc365da35, 32'h43541da2},
  {32'h44d0fab0, 32'h4344c563, 32'h4344fd42},
  {32'hc40b6cf2, 32'hc2f7970d, 32'h43299b3d},
  {32'h44451a0a, 32'h42030182, 32'h42d2407d},
  {32'hc4f3c966, 32'h42e2e19f, 32'hc158adea},
  {32'h4419a3f2, 32'h435ef0ec, 32'hc31b42d9},
  {32'hc46b53c6, 32'hc28f99d6, 32'h4311be08},
  {32'h44fc6d13, 32'hc24bfdce, 32'hc3df316c},
  {32'hc4cfde08, 32'h4383d7b0, 32'h41291b46},
  {32'h43fc7bb8, 32'hc39e4483, 32'h43455937},
  {32'hc4725c80, 32'h42fe5f0f, 32'hc2084dbe},
  {32'h443287ac, 32'h42ccd83d, 32'h42e9f83d},
  {32'hc4d9f21a, 32'hc2f16a92, 32'h4298a34c},
  {32'h450707e1, 32'hc349f066, 32'hc435c205},
  {32'hc4e29d8e, 32'h431dd760, 32'hc3302ef1},
  {32'h44587ada, 32'h439a11a2, 32'h43c62270},
  {32'hc3f3a5bc, 32'hc28380b0, 32'hc3a77582},
  {32'h43b378c8, 32'hc2bd4b4c, 32'hc3e8d6a3},
  {32'hc4b7d3de, 32'hc383b907, 32'hc3fe0b00},
  {32'h43401d4c, 32'hc2c6b3ca, 32'hc2e7bd25},
  {32'hc383537b, 32'hc37ab00b, 32'hc1ec0446},
  {32'hc3611e64, 32'h43276f31, 32'hc362dfc1},
  {32'hc4bb2b22, 32'h43068055, 32'hc2564a49},
  {32'h44fc17a5, 32'h41ed2af2, 32'hc35c4bf9},
  {32'hc5083710, 32'hc2079295, 32'hc293f1a6},
  {32'h4400741c, 32'h429a0619, 32'h42e54841},
  {32'hc4e9c1d8, 32'hc3410fa4, 32'h42b1ce2c},
  {32'h44486082, 32'h4343d24c, 32'h431edd5c},
  {32'hc4fd762c, 32'hc3370b92, 32'hc10fb32a},
  {32'h45150240, 32'h42acb5b1, 32'h425c5fec},
  {32'hc326f360, 32'h430d9b51, 32'h42d621c4},
  {32'h449f788e, 32'hc2af6642, 32'h4257e898},
  {32'hc48dc0ac, 32'h42183869, 32'hc3b75996},
  {32'hc30c4ce6, 32'h43825fec, 32'hc31a6104},
  {32'hc4f1f193, 32'h43bd4692, 32'h43a86c17},
  {32'h4434149a, 32'h42ed80f7, 32'hc302144a},
  {32'hc36a0c94, 32'h42344ca4, 32'h4112fa0e},
  {32'h446b7c4f, 32'h43259ceb, 32'h42d2e1fe},
  {32'hc4f89f02, 32'h43279dc8, 32'h42a1cc5a},
  {32'h4473b5d6, 32'hc2a68a0c, 32'hc295043b},
  {32'hc4b9c64f, 32'h41537c6a, 32'h4378a6ef},
  {32'h447301ef, 32'h42524096, 32'hc39969e1},
  {32'hc479b6b1, 32'hc2531ae5, 32'hc3c11b6f},
  {32'h451a616f, 32'h438e7914, 32'h42fa8267},
  {32'hc4340c8a, 32'h43e0b053, 32'hc39809f6},
  {32'h436f6482, 32'hc39da695, 32'hc2449f5b},
  {32'hc4e36151, 32'hc2c52e3d, 32'h4318375c},
  {32'h43bd586a, 32'hc2ce9843, 32'hc39fc2b1},
  {32'hc4891d60, 32'h4348bdeb, 32'h42bead9d},
  {32'hc38f2dd8, 32'h41f27b06, 32'h4337b579},
  {32'hc435c2be, 32'hc308597a, 32'h421b9533},
  {32'h45154bc8, 32'hc34d28ba, 32'hc3a3d0e7},
  {32'hc50150f6, 32'h4413eb1f, 32'hc1ce62f4},
  {32'h44b0b869, 32'h42b654ba, 32'hc3bc60b9},
  {32'hc4d36720, 32'hc1822ea2, 32'hc321e80f},
  {32'h43804004, 32'h4285b030, 32'hc3ac8030},
  {32'hc40eabb4, 32'hc39a711c, 32'hc3877fa7},
  {32'h44d68254, 32'h405afd50, 32'h431e0637},
  {32'hc3b724d0, 32'hc3dfe018, 32'hc2469af1},
  {32'h44ae6638, 32'h430f5213, 32'hc253ace7},
  {32'hc4a3794f, 32'h4369a82f, 32'hc3a79cd8},
  {32'h4472cdda, 32'hc28addda, 32'hc2924507},
  {32'hc2b97f52, 32'h434b4b36, 32'h43cdabf2},
  {32'h45044e9c, 32'h43b70404, 32'h4221b1ad},
  {32'hc4d7286c, 32'h43041430, 32'hc2b3e9ab},
  {32'h45078057, 32'hc3076aac, 32'hc31f360e},
  {32'hc4f727bc, 32'hc2588f9a, 32'h430b43da},
  {32'h449f7832, 32'h43a213d4, 32'hc34fd19d},
  {32'hc3e2d598, 32'hc28c25d6, 32'h420f2a8a},
  {32'h44e957b1, 32'h435785ee, 32'h433269b8},
  {32'hc491c3dd, 32'h42f9fd50, 32'h42b0e010},
  {32'h44c74d93, 32'h42807984, 32'hc3258fee},
  {32'hc47cfd57, 32'hc2df60d5, 32'h43966d22},
  {32'h4431b594, 32'h43c4ecd3, 32'hc3007f56},
  {32'hc2113940, 32'hc3425419, 32'hc3ca4a06},
  {32'h44c886e6, 32'h436ca4f4, 32'h4270c51c},
  {32'hc48c5f6c, 32'h41af1073, 32'h43970f4d},
  {32'h44ce1d57, 32'h42900c8b, 32'hc247a946},
  {32'hc43e9d8b, 32'h419d344a, 32'h436ff328},
  {32'h447435f1, 32'hc272e85d, 32'hc2d780a5},
  {32'hc3d66dd0, 32'hc3542df2, 32'hc3e4a4ae},
  {32'h44a52748, 32'h43b3fdd3, 32'h42d70c09},
  {32'hc4c1d1f0, 32'hc2901b63, 32'hc349387e},
  {32'h44add427, 32'hc2e3cd9e, 32'h430d50bd},
  {32'hc4bcdd78, 32'h4349179b, 32'hc1bdda34},
  {32'h448d548d, 32'h434b8246, 32'hc3a437d5},
  {32'hc4855aef, 32'h4348f58a, 32'hc2a363dd},
  {32'h44d6cb88, 32'hc3603065, 32'h433b7ae4},
  {32'hc3bc7098, 32'h43399934, 32'hc3414220},
  {32'h44e9eba4, 32'h4128e656, 32'hc39a0107},
  {32'hc39ae382, 32'hc305f614, 32'h4316301d},
  {32'h450f9884, 32'h429b19f7, 32'hc302f8ba},
  {32'hc4b8a692, 32'h436d2006, 32'h42528737},
  {32'h450569b2, 32'h42cfd992, 32'h42a30200},
  {32'hc533d180, 32'hc1e851de, 32'hc26ff83b},
  {32'h44ca66e8, 32'h4277b88a, 32'hc1f3fb8a},
  {32'hc48a2ef5, 32'hc365360d, 32'h43a7b779},
  {32'h44fe8094, 32'hc3a4941a, 32'hc2213df6},
  {32'hc480ca2b, 32'h4340d39c, 32'h42907e9a},
  {32'h4390eafc, 32'hc39073ee, 32'h43ccd3aa},
  {32'hc43d6a5c, 32'h436038e5, 32'h428e9bd4},
  {32'h44aebebb, 32'h421b5b3b, 32'h43d3cada},
  {32'hc16ae6c0, 32'hc29e31e3, 32'h431528f5},
  {32'h44c73e62, 32'hc3579f8a, 32'h4389b1ad},
  {32'hc51fa875, 32'hc2def65c, 32'hc3d36f06},
  {32'h44fa4ef3, 32'hc2953b4e, 32'hc3c93d26},
  {32'hc4347db7, 32'h433e6cfa, 32'h43b3f9c5},
  {32'h44a6ca2f, 32'h439f9eb7, 32'hc236e69b},
  {32'hc42fa0e8, 32'hc18e43d1, 32'h4240b5e4},
  {32'h444489ce, 32'h4351c0ac, 32'h4390525e},
  {32'hc4e238ae, 32'hc32286e9, 32'hc2a6f0a3},
  {32'h44811eb1, 32'h42c7a3a9, 32'hc24294bb},
  {32'hc4fe3288, 32'hc38841b9, 32'h4273d925},
  {32'h44feb0be, 32'h42a2ef04, 32'hc2adb11e},
  {32'hc3b5cadc, 32'hc3d516a8, 32'hc2e20e64},
  {32'h447c7e98, 32'hc3b78a85, 32'hc34b876f},
  {32'hc3e31f82, 32'h43a96c13, 32'h4386b6ac},
  {32'h44ad9e6f, 32'hc02f52ee, 32'h42b4ac91},
  {32'hc49ee9b1, 32'hc2a8b994, 32'h427e43e4},
  {32'h43a458e1, 32'hc356889c, 32'hc3837da6},
  {32'hc4740616, 32'h4234b919, 32'h432fa9fa},
  {32'h447cf04a, 32'h42bfb71c, 32'h415a6a91},
  {32'hc442a691, 32'hc3785f11, 32'h435aeb19},
  {32'h4505f6ec, 32'h4100d275, 32'hc34e591e},
  {32'h4211c9b0, 32'hc31e4d64, 32'h43c42cd6},
  {32'h44a6653c, 32'hc3a87baa, 32'h43ec9bce},
  {32'hc508f8ae, 32'h426d10e1, 32'h4317beda},
  {32'h43c281ac, 32'h429bf306, 32'h43886012},
  {32'hc2e8d790, 32'hc27e5630, 32'hc3ecbc32},
  {32'h4460de45, 32'h430c5690, 32'h43589d49},
  {32'hc4ad4b81, 32'h43854f09, 32'h43884839},
  {32'h44b6ad93, 32'hc3855f6d, 32'hc34f708a},
  {32'hc493b80a, 32'hc24053f3, 32'h42c4d11e},
  {32'h42a84850, 32'h43a34e31, 32'h42a7537e},
  {32'hc50d6398, 32'h42dd9ca5, 32'h4120706b},
  {32'h44f3c29e, 32'h4213fc73, 32'hc307b440},
  {32'hc48a3740, 32'hc3cb1a1b, 32'hc37e4997},
  {32'h44f7a844, 32'h4302fb80, 32'hc382134b},
  {32'hc501c734, 32'h43bbd5fc, 32'hc36b92bd},
  {32'h44cc63ff, 32'h434a880b, 32'h4368da32},
  {32'hc508e1d7, 32'hc21ebca2, 32'hc316e5dc},
  {32'h44d1d24d, 32'hc3ea54d0, 32'hc1e8bacc},
  {32'hc50ed553, 32'h427fc342, 32'h4399b3f0},
  {32'h4396d4f4, 32'h43354b7e, 32'hc2f4f951},
  {32'hc4b0a95d, 32'h40bf50c0, 32'h42d0b8e6},
  {32'h44c3d752, 32'hc3b63617, 32'h4366276e},
  {32'hc483b443, 32'hc38f0959, 32'hc31cd921},
  {32'h444629be, 32'h43af373c, 32'h426dfaa0},
  {32'hc4e4539f, 32'hc3a44ff6, 32'hc306bd7a},
  {32'h44c24f5a, 32'h426e8115, 32'h426f6124},
  {32'hc3d53b65, 32'h419a055a, 32'h435b8c7d},
  {32'h44f9b1b0, 32'h4320d138, 32'h429832fc},
  {32'hc4d1a523, 32'hc2b7c51b, 32'h43de7aa9},
  {32'h44bc487c, 32'hc32a92e7, 32'hc34b38b7},
  {32'hc469ee05, 32'hc1547539, 32'h42da7e58},
  {32'h4454cb78, 32'hc321a39c, 32'h441a2dbb},
  {32'h41938550, 32'hc346bd76, 32'hc1db019e},
  {32'h449beb50, 32'h41ebef9d, 32'hc35b8f7a},
  {32'hc4be651b, 32'hc30b570a, 32'h4382afe3},
  {32'h44a82ed3, 32'h433494a9, 32'hc31bc64c},
  {32'hc496a4eb, 32'hc303b689, 32'h42ae8bf6},
  {32'h450d49ae, 32'h4228c811, 32'h428eefa0},
  {32'hc48a8f3e, 32'hc3519313, 32'hc38a5a1a},
  {32'h451f3c3e, 32'hc3359914, 32'h4404afc6},
  {32'hc4486bc6, 32'hc351e909, 32'h432b257a},
  {32'h44937a64, 32'h42fe21e2, 32'h42d9105b},
  {32'hc51791ab, 32'h435df23e, 32'hc19e9f58},
  {32'h43427b00, 32'h428e2bcf, 32'h426c837d},
  {32'hc5036f6f, 32'h43587cc9, 32'hc358d73f},
  {32'h44ca5715, 32'h429df491, 32'hc2b4a9b0},
  {32'hc4064ac0, 32'hc2ed1689, 32'hc2ae7086},
  {32'h44c38492, 32'h438ce363, 32'hc35d3029},
  {32'hc503677d, 32'h439c858e, 32'h435aafc3},
  {32'h44cd2ce0, 32'h41d967ee, 32'h43762c10},
  {32'hbf8ac800, 32'hc40a2082, 32'hc37a157e},
  {32'h44e0a130, 32'h43282544, 32'h42d233df},
  {32'hc506f3c2, 32'hc2aed32e, 32'h432ea15d},
  {32'h45090f80, 32'hc38811c1, 32'h43185b05},
  {32'hc46a70d2, 32'hc2f687d0, 32'h423c16b4},
  {32'h451cda14, 32'hc2de4f11, 32'hc2bdea73},
  {32'hc4add87d, 32'hc3348271, 32'h42ec0d82},
  {32'h4501ab7e, 32'hc2dee31e, 32'h4304fd22},
  {32'hc5012130, 32'hc3b9b01a, 32'hc2b7f1cf},
  {32'h4502f376, 32'hc2d0a203, 32'h4215f605},
  {32'hc4822826, 32'hc33dd127, 32'hc34f8580},
  {32'h43810cb8, 32'h438ef660, 32'h42bb4ccf},
  {32'hc3a51e38, 32'h42aa0307, 32'h4297a81d},
  {32'h446003c5, 32'hc2dfcdd7, 32'h43809fe1},
  {32'hc436fd62, 32'hc334da45, 32'h43063bb6},
  {32'h44a4fd61, 32'hc265752c, 32'hc3360ac3},
  {32'hc339630e, 32'hc2aa7698, 32'hc3c3e978},
  {32'hc40864ec, 32'h4330c23a, 32'h431c1729},
  {32'hc385c818, 32'h4354813b, 32'hc3a57c59},
  {32'h43971794, 32'h428364f4, 32'h4347d5c3},
  {32'hc4ccf9a4, 32'hc39c7349, 32'hc273835d},
  {32'h43a8bb92, 32'h4374dbf5, 32'hc28d8caf},
  {32'hc4c243af, 32'hc35cd2b6, 32'hc3279a47},
  {32'h448aa6c0, 32'hc413a3a7, 32'hc305710e},
  {32'hc475ba08, 32'h4300875f, 32'hc39b58d3},
  {32'h450c07f2, 32'h43b027d9, 32'hc1aec81e},
  {32'hc509c81b, 32'h420d01ee, 32'hc283beab},
  {32'h449bc806, 32'h4346b761, 32'h438a5644},
  {32'h43787bb0, 32'h4030e8b0, 32'hc364c022},
  {32'hbff67900, 32'h4308ae01, 32'h43356d98},
  {32'h42cad1e0, 32'hc32c2fa8, 32'h43cdc12e},
  {32'h4267cf80, 32'hc299458b, 32'h4354fa64},
  {32'hc3969dcc, 32'h3f84e200, 32'h4358ae34},
  {32'h4497be85, 32'h43107a61, 32'hc2f1fd13},
  {32'hc4f050de, 32'h42f52687, 32'hc30d5854},
  {32'h45042187, 32'hc3a80aa1, 32'h43910718},
  {32'hc483358d, 32'hc3a5f598, 32'h42e65c4a},
  {32'h44841f94, 32'h430bcec4, 32'h42d94048},
  {32'hc338a548, 32'hc386bb48, 32'h433eff1e},
  {32'h449738aa, 32'hc2a7e08e, 32'h43b7b418},
  {32'hc4825196, 32'hc2844c09, 32'h42f82a4c},
  {32'h44607f9a, 32'h42a1247f, 32'hc1f85720},
  {32'hc4b7c365, 32'hc369cf06, 32'hc38824c5},
  {32'h44a13c3a, 32'hc299505b, 32'hc3ab37d1},
  {32'hc4d992ac, 32'hc3f49ab1, 32'h43116ae6},
  {32'h44b78cca, 32'hc306470a, 32'hc1e7182a},
  {32'hc4555a98, 32'hc3928ce8, 32'hc3b72b8e},
  {32'h44e41114, 32'hc14ee3c1, 32'h3f95775c},
  {32'hc4ad45e3, 32'h41d03aac, 32'hc39975c8},
  {32'hc5008d26, 32'hc0bf6160, 32'h420fba2f},
  {32'h44b4556e, 32'hc3417e25, 32'h43b2de54},
  {32'hc4b39cf3, 32'hc3acd798, 32'hc2e3a303},
  {32'h434e65d2, 32'h419e56de, 32'h425748d4},
  {32'hc4acae8c, 32'hc2955fd9, 32'hc3e07ee7},
  {32'h447230a5, 32'hc1ecca7b, 32'h43d4dd2d},
  {32'hc49a7547, 32'h42c221de, 32'h4314f678},
  {32'h44e68c44, 32'h432ec636, 32'h4066d80c},
  {32'hc46b89fa, 32'h438034a9, 32'hc3c1d6fa},
  {32'h44c88758, 32'h432bcdbb, 32'hc1a51d43},
  {32'hc499d59d, 32'h435a0625, 32'hc2269f93},
  {32'h44b5289f, 32'hc3775405, 32'h43981f95},
  {32'hc503a2e9, 32'h4250745c, 32'h43057413},
  {32'h4513535f, 32'h43dc0d83, 32'hc278a4e1},
  {32'hc4fa6ed4, 32'h4318d83a, 32'hc359449a},
  {32'h448803aa, 32'hc307c749, 32'hc35e4a3f},
  {32'hc47ab55c, 32'h43297dea, 32'h432c2d70},
  {32'h451531b4, 32'h43eac5a7, 32'hc3735abf},
  {32'hc5041d14, 32'hc32b53e4, 32'hc0837b6b},
  {32'h4400f782, 32'h4005e6ac, 32'h434004a1},
  {32'hc4b7672b, 32'h4319f93f, 32'hc3cccacf},
  {32'h43dcb3f6, 32'hc3106892, 32'h42686b56},
  {32'hc3b412a4, 32'h437af9a8, 32'hc13c9fb1},
  {32'h44ff454e, 32'hc3c688fb, 32'hc1a41587},
  {32'hc4eb0d77, 32'hc2608a46, 32'h434ed90e},
  {32'h43f2d710, 32'h42e844fc, 32'h43168019},
  {32'hc43c7f40, 32'h42a1ca1d, 32'h4324c747},
  {32'h43f0c304, 32'hc373c2dc, 32'hc2fec4e1},
  {32'hc3bb991f, 32'hc37f4187, 32'hc41b35ce},
  {32'h4489c943, 32'hc3c9be57, 32'h42408334},
  {32'hc4f927da, 32'hc20efa81, 32'hc2ff4062},
  {32'h4400e538, 32'h42c52db7, 32'hc2c75830},
  {32'hc504cfdb, 32'hc393cf01, 32'hc1b7b4fc},
  {32'h44b7790c, 32'h430f4e17, 32'h438c3846},
  {32'hc47c6c04, 32'hc2dd18b8, 32'hc30bb48e},
  {32'hc3fb4dac, 32'hc324590f, 32'hc1390915},
  {32'hc40f1c0e, 32'hc3d8f3f2, 32'hc3cdc15d},
  {32'h440d38b0, 32'h4319d83f, 32'h4407d789},
  {32'hc22dad40, 32'hc294dbe9, 32'h43aaad5c},
  {32'h44c2d360, 32'h42904758, 32'h42b1632c},
  {32'hc3e7b4a2, 32'hc38566f4, 32'h4320f795},
  {32'h44ade28d, 32'h435ca91c, 32'hc31c2ef2},
  {32'hc2c8acfc, 32'hc36bf21c, 32'hc009fd79},
  {32'h443fb665, 32'hc289470d, 32'h4125389e},
  {32'hc5112c62, 32'hc1dee3ca, 32'hc407784d},
  {32'h43d59eb7, 32'h4411a7a1, 32'hc22046af},
  {32'hc4403af9, 32'hc25df579, 32'h425a3a75},
  {32'h451eebea, 32'h4291b3de, 32'h42b4efc2},
  {32'hc4e062a4, 32'h4385a866, 32'h40433600},
  {32'h450837c6, 32'h436482e4, 32'hc3b98a6d},
  {32'hc3e79ef3, 32'hc24ad67e, 32'hc2ade067},
  {32'h44bc55c1, 32'h43ac572f, 32'h43e97549},
  {32'hc50ae10e, 32'hc3dbaee8, 32'hc382d470},
  {32'h44fd39ad, 32'hc3ae697c, 32'hc31de3cd},
  {32'hc4ee5ade, 32'h43b90f7b, 32'h432d9bf6},
  {32'h44cdc65c, 32'h4306f051, 32'hc3024ee4},
  {32'hc3721b39, 32'h42c06b39, 32'h43ee6c61},
  {32'h445cf66c, 32'hc2d4109e, 32'h43ca75fe},
  {32'hc47ecb70, 32'hc3836376, 32'hc43269df},
  {32'h44c40bb3, 32'hc34d5e16, 32'h434ec925},
  {32'hc4e85cbe, 32'h422702fb, 32'h4230d3fa},
  {32'hc3a4356c, 32'h43cbbb93, 32'h439da584},
  {32'hc4fff6db, 32'hc3658540, 32'hc3a6222d},
  {32'h4327eea4, 32'h431e2923, 32'h430ea9ec},
  {32'hc4defcd8, 32'h434b4b76, 32'hc33f5bb1},
  {32'h44ad8ad5, 32'hc338efbb, 32'h422d9bdc},
  {32'hc4bbb296, 32'hc11b181a, 32'h43373c19},
  {32'h44000a42, 32'h432d3375, 32'hc3944de7},
  {32'hc4fbc5b1, 32'hc28add54, 32'hc128e882},
  {32'h44d26f8e, 32'hc1aab6af, 32'h436e5bab},
  {32'hc468d990, 32'h42a1aac0, 32'hc26f957b},
  {32'h44828524, 32'h424bdf23, 32'h434411f7},
  {32'hc4b104ff, 32'hc3ace90e, 32'h43a025de},
  {32'h444c4800, 32'h436cd6f7, 32'h427d3247},
  {32'hc24d4f00, 32'hc2ad1426, 32'hc33b9ba4},
  {32'h451875fb, 32'h43037397, 32'h4327370b},
  {32'hc42a6b08, 32'hc410cc20, 32'hc3619a54},
  {32'h44f9614b, 32'hc20d382b, 32'hc3239c2b},
  {32'hc1bb2d0e, 32'hc378bb91, 32'h42b70602},
  {32'h44bd5561, 32'h43b17ef6, 32'h431e1b8b},
  {32'h4373f2a6, 32'hc1fbfaeb, 32'h421c4f39},
  {32'h44e442fb, 32'hc036a19a, 32'hc31b35ee},
  {32'hc4053a11, 32'h430ee382, 32'hc2d3045f},
  {32'h44f6bd8e, 32'h40f335b6, 32'hc39d5d80},
  {32'hc509d506, 32'h431f9ceb, 32'hc342bc68},
  {32'h44a40538, 32'hc3b44078, 32'h438254e3},
  {32'hc4f91a20, 32'h432cdb91, 32'h431c9936},
  {32'h4492cc75, 32'hc377dc6d, 32'hc21dbdaf},
  {32'hc4713298, 32'hc32b2a2d, 32'h432eef4e},
  {32'h44e3a40a, 32'h42ebae12, 32'hc3c15a0b},
  {32'hc49d16fe, 32'hc3427030, 32'hc30b8f3b},
  {32'h448fdad3, 32'h428ac282, 32'hc3861677},
  {32'hc490911f, 32'hc28bd700, 32'hc36a5c8a},
  {32'h45092a52, 32'hc2ba2b13, 32'hc2994ff4},
  {32'hc4802d8f, 32'hc094bbd4, 32'h4416940d},
  {32'h44a7e769, 32'hc2bd5c0f, 32'h415a0d5c},
  {32'hc4f1aa6e, 32'h417faada, 32'h42d6a3cd},
  {32'h44f21a21, 32'h434a3c73, 32'hc3d44ebd},
  {32'hc487e796, 32'h43c5e966, 32'h42dc20a3},
  {32'h43b47462, 32'hc31a11d0, 32'hc33f551c},
  {32'hc42be660, 32'h43f7c963, 32'h4361d199},
  {32'h45040d00, 32'hc389a963, 32'h4207de11},
  {32'hc49739d9, 32'h427232c5, 32'h43060e8d},
  {32'h442997ea, 32'hc3ce4d80, 32'h41809e0e},
  {32'hc4cde5e8, 32'hc39a8641, 32'h433f3d4f},
  {32'h450d7db4, 32'hc1ef47c4, 32'h433197aa},
  {32'hc47dc18b, 32'hc2fecb19, 32'hc36139d5},
  {32'h447d8417, 32'hc3c29d93, 32'hc30ca4e9},
  {32'hc4a2f6b0, 32'h428c41c6, 32'h418cd414},
  {32'h444f7de4, 32'h438159c4, 32'hc2d16018},
  {32'hc2e4e059, 32'hc3188c34, 32'hc14d32ca},
  {32'h44072c7e, 32'hc31b42b4, 32'hc316f7c8},
  {32'hc4893bd4, 32'hc492ef9b, 32'hc1a4fef7},
  {32'h442a5d1e, 32'h42cf75e2, 32'hc3412d4b},
  {32'hbfc05ec0, 32'h43186f69, 32'h43519329},
  {32'h44b27bf0, 32'hc3ef820c, 32'hc3412ec6},
  {32'hc4975ecf, 32'h428c82ca, 32'hc3162a3b},
  {32'hc13aaa80, 32'hc3072903, 32'hc2f9575e},
  {32'hc46f5563, 32'hc37a1a21, 32'h41c138be},
  {32'h448cb363, 32'hc20b5d27, 32'hc3818d97},
  {32'hc44552d0, 32'hc298291c, 32'h43aaeca9},
  {32'h44bae16a, 32'hc408e4f1, 32'h42b5d08f},
  {32'hc4ecfc50, 32'hc334b556, 32'hc28f88d4},
  {32'h44a19415, 32'h4280bffa, 32'h42c46c36},
  {32'hc45a25b0, 32'h43979016, 32'h43b168dd},
  {32'h44dd4a2c, 32'h43147c85, 32'h42c3383c},
  {32'hc4398e70, 32'hc24d482e, 32'h438c16bd},
  {32'h4517c620, 32'hc2a02c87, 32'h41cd7bea},
  {32'hc49ec5ce, 32'h433f305f, 32'h43952dee},
  {32'h43bb0510, 32'h44070a0a, 32'h43696d63},
  {32'hc46ce594, 32'hc111af84, 32'h439821d5},
  {32'h44a4c874, 32'hc301cd63, 32'h4417b046},
  {32'hc4439a2c, 32'h4218ef89, 32'hc3b14d25},
  {32'h44c3310e, 32'h4235797d, 32'h42f127f3},
  {32'hc37ec26c, 32'h422a59ab, 32'h40ccb2ff},
  {32'h44921d30, 32'hc3afff2e, 32'hc444eb0e},
  {32'hc51472c7, 32'h41504f9a, 32'h41a6e0c2},
  {32'h44044a50, 32'hc356ea54, 32'hc2298a4a},
  {32'hc35f2036, 32'hc32c2cf3, 32'h430339f6},
  {32'h4386ae04, 32'hc327c0d2, 32'hc16f0a62},
  {32'hc4e3d676, 32'h415bac3e, 32'h430edaee},
  {32'h445157ff, 32'hc3965966, 32'h4336e709},
  {32'hc4b0510c, 32'hc401a242, 32'h43ab4229},
  {32'h44ed825d, 32'hc36e7998, 32'h423d15be},
  {32'hc3f72e74, 32'hc23605d8, 32'h43dff155},
  {32'h44813679, 32'h421898d0, 32'hc404ee1d},
  {32'h43eb7e2c, 32'hc39013d3, 32'hc4052274},
  {32'hc2ece1d0, 32'h438567c4, 32'hc198bc04},
  {32'hc46dbd9d, 32'h42f86c38, 32'h43a90ee8},
  {32'h42f969c0, 32'hc2d736b8, 32'h436c7a0a},
  {32'hc3f9d60c, 32'hc35cf2e3, 32'hc307a844},
  {32'h440ad11b, 32'hc40334a4, 32'hc39307b3},
  {32'hc4a6c086, 32'hc3662ebb, 32'hc280c04e},
  {32'h44d6f15a, 32'h40c103da, 32'hc201c4a6},
  {32'hc4799856, 32'h4323b96a, 32'h42021727},
  {32'h449dac41, 32'h420276fe, 32'hc331caaa},
  {32'hc47e8050, 32'h428f5b7a, 32'h42921ca2},
  {32'h44a299ad, 32'hc3556a27, 32'hc3a10734},
  {32'hc3cd1a7d, 32'h4390aeac, 32'hc316d2f0},
  {32'h446e0fac, 32'h4246dc1b, 32'hc2a2a672},
  {32'hc4f7ff0b, 32'h42fc401e, 32'h4388b435},
  {32'h44ca76dc, 32'hc202efa3, 32'h4309fed1},
  {32'hc3ebc630, 32'h42bde648, 32'hc28b9f06},
  {32'h44fa5143, 32'hc1486ca4, 32'hc32efe4e},
  {32'hc4c6b1dd, 32'hc2996d02, 32'hc2eff94d},
  {32'h44f9f5f9, 32'hc25083e4, 32'h40291d06},
  {32'hc430a1e4, 32'h420e58c2, 32'h4331d505},
  {32'h44814450, 32'hc3078fda, 32'hc13efefa},
  {32'hc507a71c, 32'h42fbaf21, 32'h42aa36af},
  {32'h4506ca58, 32'h43982e9f, 32'h435fa236},
  {32'hc35b5bb4, 32'h42b38104, 32'h42a97316},
  {32'h44f275f8, 32'hc3142db2, 32'hc30dc976},
  {32'h40df0360, 32'hc18691ed, 32'h3e80dd00},
  {32'h44bfc262, 32'hc1b2a7da, 32'h43853993},
  {32'hc50240cf, 32'hc20f9f21, 32'h43530475},
  {32'h44f96a74, 32'h43bf789c, 32'h42f250e6},
  {32'hc4c4b2fc, 32'h4375bd39, 32'h426f46fc},
  {32'h45022b6a, 32'hc33802ec, 32'hc35a9cf6},
  {32'hc4cd6992, 32'h426a73bd, 32'hc193310f},
  {32'h441cbf81, 32'hc3f8436a, 32'hc25e5b88},
  {32'hc4530b36, 32'hc24ef720, 32'h42468e7c},
  {32'h44d78fc6, 32'hc3085f5c, 32'hc21806a3},
  {32'hc4c893ee, 32'hc31806ca, 32'hc2451598},
  {32'h44b9e4d8, 32'h43a1b118, 32'h43d6960f},
  {32'hc34091c0, 32'h42495840, 32'h435b4f5e},
  {32'h44677536, 32'h433cfef0, 32'h41c54bee},
  {32'hc4388579, 32'h421d7f56, 32'hc19f51f3},
  {32'h44e79d10, 32'hc328b802, 32'h42ad5bc5},
  {32'hc4cc92b6, 32'h43c9e74c, 32'hc2009306},
  {32'h44fec82d, 32'hc36135b8, 32'h43700377},
  {32'hc3bf97d1, 32'h43ca88af, 32'h43c154c4},
  {32'h45086900, 32'h43396f50, 32'h438d8ba3},
  {32'hc4162a68, 32'h43046e9f, 32'hc3aa1785},
  {32'h4384c22c, 32'hc3d06751, 32'h43a7ebbd},
  {32'hc3b29d5b, 32'h42718530, 32'hc21585ea},
  {32'h44bd387f, 32'h43b54a32, 32'hc3bc182c},
  {32'hc50167e7, 32'h4332f959, 32'hc2a21364},
  {32'h44f75a96, 32'hc165e951, 32'h43d63b67},
  {32'hc4c2e0b1, 32'hc3311684, 32'h430d495a},
  {32'h45076763, 32'h40d2ee60, 32'h43c83248},
  {32'hc50345da, 32'h433e99f8, 32'hc1819f4c},
  {32'h44854717, 32'hc293a5d8, 32'hc3635cba},
  {32'hc433b974, 32'hc1a21ab0, 32'h4351e059},
  {32'h446ed699, 32'h410f81a2, 32'h420d83ab},
  {32'hc449a556, 32'hc22871a8, 32'h438b785b},
  {32'h443df602, 32'h42a26b4d, 32'h43a29b0d},
  {32'h424bd210, 32'h43d7c68b, 32'h4208fcb8},
  {32'h415432da, 32'hc297aabb, 32'hc1df28c4},
  {32'hc47fe534, 32'h428bb393, 32'hc1427bce},
  {32'h44ec13ee, 32'hc318b330, 32'h40edcf29},
  {32'hc324ab7b, 32'hc1db68a1, 32'h43cb1c63},
  {32'h449fad05, 32'hc26c7e81, 32'hc3609d33},
  {32'hc4e0dcfd, 32'hc2b96fed, 32'hc33c45f8},
  {32'h43624d20, 32'h43755abf, 32'hc30accf7},
  {32'hc48db602, 32'hc30a1542, 32'h42815c23},
  {32'h4501d747, 32'h42d2a8c3, 32'h432dd377},
  {32'hc4cd057c, 32'h43369c22, 32'h4231311e},
  {32'h43348e36, 32'hc2e70a28, 32'h43d259ad},
  {32'hc4c54b25, 32'h40edd8a8, 32'h42f03db6},
  {32'h450edfc5, 32'hc0ebaa30, 32'h43243181},
  {32'hc4a72090, 32'hc3031d7b, 32'hc3114b43},
  {32'h44836361, 32'h43935129, 32'h412260f0},
  {32'hc3933738, 32'hc321424e, 32'hc107f683},
  {32'h4413a080, 32'h44249dd9, 32'h41a0afa7},
  {32'hc4f2e22e, 32'hc347e855, 32'h42eccd7b},
  {32'h445bf46c, 32'hc2016253, 32'h42962b0d},
  {32'hc4c0616c, 32'h41948325, 32'h42f12730},
  {32'h44c9b57c, 32'h436f9ba7, 32'hc3ffe275},
  {32'hc4f12948, 32'hc391f878, 32'h429e1da9},
  {32'h44712a56, 32'hc1ede1d6, 32'hc38a27ad},
  {32'hc3d1a0b8, 32'h42d9a89e, 32'hc23d51bf},
  {32'h44c9c7ad, 32'hc316cab4, 32'hc1ffaadf},
  {32'hc4947558, 32'hc3148c5f, 32'h42ec6b04},
  {32'h4495ed99, 32'h43418bdd, 32'h41a1fc9f},
  {32'hc352eaa4, 32'h4311e09f, 32'h42a08201},
  {32'h44b572ea, 32'h43499c19, 32'hc12a1889},
  {32'hc353a420, 32'hc36fbd74, 32'h424b61b0},
  {32'h44c0b003, 32'h432036f4, 32'h42f42f18},
  {32'hc48fdec1, 32'hc22452b4, 32'hc2b5b180},
  {32'h450a761b, 32'h43c344c4, 32'h438089d3},
  {32'hc4ebb148, 32'hc2cf8c5c, 32'h42bca450},
  {32'h4500a996, 32'h4243ab91, 32'h40da5298},
  {32'hc4b8242b, 32'h42bbf75a, 32'h436115bc},
  {32'h43a1e9e8, 32'hc28542b6, 32'h432ba93f},
  {32'hc4bf54d4, 32'h43077b55, 32'hc24a15f4},
  {32'h43ed0f80, 32'h435f0cd0, 32'h43ec7753},
  {32'hc4046e50, 32'h4239c2be, 32'h437befaa},
  {32'h44d4c687, 32'hc3cd00ea, 32'hc3a53900},
  {32'hc4aa6f0e, 32'hc2b8cb20, 32'h42c8988a},
  {32'h438e0ba5, 32'hc391d71a, 32'hc429a376},
  {32'hc3c44a00, 32'hc384005f, 32'hc1f6cfb5},
  {32'h44199a9c, 32'h4390789c, 32'hc39dfd33},
  {32'hc4c30409, 32'h42a96d76, 32'hc3139187},
  {32'h41da4240, 32'h4373748d, 32'hc2e780b1},
  {32'hc41e1aa2, 32'h41bde443, 32'h4241f1da},
  {32'h44d78ceb, 32'hc198be20, 32'h42af6f5c},
  {32'hc4f21531, 32'hc3ee51b7, 32'hc2d8532a},
  {32'h4441e589, 32'h4383f235, 32'h42f68363},
  {32'hc4f4663e, 32'h436fa222, 32'h423259fa},
  {32'h44e60d1a, 32'h40be8020, 32'hc2603c26},
  {32'hc4f6a21a, 32'hc1be98a4, 32'h43b1494f},
  {32'h443a6688, 32'hc2e08659, 32'hc39a0759},
  {32'hc4a68223, 32'h439d1602, 32'h4338166c},
  {32'h451002ec, 32'h43888566, 32'h437fbc56},
  {32'hc3c04a9b, 32'hc34accdb, 32'h42f5de9f},
  {32'h4511c286, 32'h434d2d66, 32'hc34f8858},
  {32'h428ad7d5, 32'h3f6fd7cd, 32'hc37d50ef},
  {32'h44a3387c, 32'h4380562e, 32'hc310c7d6},
  {32'hc45503ec, 32'h4313acda, 32'h4318a2f1},
  {32'h44f68d89, 32'hc23916bb, 32'h4358ee8a},
  {32'hc4ee7b09, 32'h43ab9b20, 32'h4296c382},
  {32'h4509c8fe, 32'h4138927e, 32'hc293ef53},
  {32'hc39c21ac, 32'h43d0d12d, 32'h42fc0faa},
  {32'h44baf9a8, 32'hc3b67f43, 32'h430107db},
  {32'hc51de02a, 32'h42d2ddfd, 32'h430682fe},
  {32'h447c8480, 32'h43859d57, 32'h436574ac},
  {32'hc4de927e, 32'h437085df, 32'h42af16b6},
  {32'h44553fde, 32'hc22dec39, 32'hc2ebda44},
  {32'hc4788f8c, 32'hc18394e2, 32'h42b6c988},
  {32'h451d1436, 32'hc237622a, 32'hc30392e6},
  {32'hc465d610, 32'h4382ebc8, 32'h438281f5},
  {32'hc3702060, 32'h429aa270, 32'h428fb52a},
  {32'hc4a35447, 32'hc214b03c, 32'hc10bbc49},
  {32'h4518f228, 32'h4212dbb8, 32'h433dd161},
  {32'hc4aaeb07, 32'h42812f8d, 32'h4298fb96},
  {32'h441f108e, 32'hc3b12ace, 32'hc337259b},
  {32'hc4b5cd9f, 32'hc339e664, 32'h435f2855},
  {32'h4501e944, 32'h42b716fa, 32'hc40ebd55},
  {32'hc26e13db, 32'hc3965110, 32'hc3031d77},
  {32'h4443da1d, 32'hc298a716, 32'hc3002255},
  {32'hc4877cf1, 32'hc241087a, 32'hc3d13287},
  {32'h45206bbb, 32'h42365500, 32'h439a0a6e},
  {32'hc5079c4b, 32'hc33f464e, 32'hc3bb1cc3},
  {32'h43a94f28, 32'hc27eddce, 32'h421cacf0},
  {32'hc409d818, 32'h423ea78e, 32'h42998f06},
  {32'h440128a4, 32'h4321d8dd, 32'h424a15b4},
  {32'hc421aebc, 32'h41ae6d92, 32'hc2f4a670},
  {32'h42b297b8, 32'h4364cf6b, 32'hc394d1ea},
  {32'hc3014970, 32'h43a4f6d9, 32'h43912669},
  {32'h44c3007c, 32'hc2ecb2de, 32'h43887e61},
  {32'hc50b5448, 32'hc392ffa2, 32'hc2cc630f},
  {32'h440bfae2, 32'h4326b2dd, 32'h43aba14a},
  {32'hc3e0c710, 32'hc302bba1, 32'h438c3988},
  {32'h44f31a98, 32'h435f2914, 32'hc2344563},
  {32'hc3017540, 32'h42ba222c, 32'h432a47fa},
  {32'h451a400f, 32'hc330b914, 32'h435903b1},
  {32'hc33b9271, 32'hc2aabafa, 32'hc3ad3dfb},
  {32'h44a63468, 32'hc299485b, 32'hc2be32b2},
  {32'hc47f4d85, 32'h43b604db, 32'hc20b5a54},
  {32'h44641e38, 32'h43b49c9c, 32'h4317d4f5},
  {32'hc31d06d0, 32'hc301b31a, 32'h430ebed1},
  {32'h43eb9878, 32'hc1b702c9, 32'h430fe57a},
  {32'hc42b2db4, 32'hc33ba797, 32'h437c9d13},
  {32'h44625b43, 32'hc346e729, 32'h43767f5f},
  {32'hc408b8c6, 32'hc3014f42, 32'hc289cb96},
  {32'h4500df30, 32'h4252275e, 32'h42f88739},
  {32'hc4ef84eb, 32'h43b3666e, 32'h41d11b64},
  {32'h4503f697, 32'hc36944da, 32'h42816f18},
  {32'hc4e5c3c7, 32'h438ad91a, 32'h431b5ef1},
  {32'h44cf7cca, 32'hc3bd9bb0, 32'hc31f5513},
  {32'hc4438437, 32'h430c02ca, 32'h3ed2615c},
  {32'h44fa44ba, 32'h43161833, 32'hc389ae6f},
  {32'hc4874362, 32'h4353279f, 32'hc24089d2},
  {32'h45122e71, 32'hc18ce5a5, 32'h43a54079},
  {32'hc4da6a66, 32'hc33b258f, 32'hc26b67e7},
  {32'h428f6d70, 32'h438a8488, 32'hc3c6bc21},
  {32'hc4fd2bec, 32'hc3217d70, 32'h424f4e52},
  {32'h4301290d, 32'h42ce094c, 32'h431a8f1e},
  {32'hc4d1f448, 32'hc3942acf, 32'h44170a18},
  {32'h44dfb168, 32'h42309f0c, 32'hc2e0ad72},
  {32'hc4e46c81, 32'hc36f0eba, 32'hc31b32fe},
  {32'h43ddbd0d, 32'h43c96a6c, 32'hc21250c2},
  {32'hc3839c80, 32'hc39686db, 32'hc29b947b},
  {32'h44f5d60a, 32'hc303443c, 32'hc2d37434},
  {32'hc5020325, 32'hc2e781f6, 32'hc3a7a1af},
  {32'h44f2f7d7, 32'h42394538, 32'h433eca9a},
  {32'hc4ef226d, 32'h43b05206, 32'hc35cf21a},
  {32'h43845574, 32'hc3768b6d, 32'hc31161f6},
  {32'hc5085ccf, 32'hc35e8764, 32'hc2c967c7},
  {32'h437cb217, 32'hc37d0ae5, 32'h43a314ed},
  {32'hc4f41625, 32'h4281c15a, 32'hc34c740a},
  {32'h43826d26, 32'h4380090a, 32'hc3909c3e},
  {32'hc2940b1f, 32'hc222f015, 32'h41ca80fa},
  {32'h443318b2, 32'h4266bac8, 32'h40bad827},
  {32'hc4465c10, 32'hc33ed7c0, 32'h43139f95},
  {32'h44cdc622, 32'hc09b4e3a, 32'hc22aaf3f},
  {32'hc4132724, 32'hc354f612, 32'h436a3010},
  {32'h449b20bf, 32'h42dbbed3, 32'hc2e622bd},
  {32'hc5190d13, 32'h43140fc5, 32'hc312a65c},
  {32'h438b7da6, 32'hc2711a86, 32'h42a99d03},
  {32'hc488924a, 32'hc36361e7, 32'h43e77840},
  {32'h45060585, 32'hc2434dd7, 32'hc320bea6},
  {32'hc44070fc, 32'hc33d4593, 32'h4292802b},
  {32'h44c50a46, 32'hc2899e67, 32'h419b75d4},
  {32'hc425d1f0, 32'hc3c20409, 32'hc3460a2f},
  {32'h43720011, 32'h4193378c, 32'h42303bad},
  {32'hc4d73f58, 32'h43a97480, 32'hc169ec42},
  {32'h44f41d90, 32'h43279601, 32'hc3422ca8},
  {32'hc449586c, 32'h4358f1a5, 32'h4228ade6},
  {32'h4514fc41, 32'h4390e0fb, 32'h43a46dbb},
  {32'hc4c057f4, 32'hc3a8f705, 32'hc26e3f25},
  {32'h44c02a27, 32'hc1d532e6, 32'h4334744f},
  {32'hc39fef91, 32'hc341ef4f, 32'h4240b4f8},
  {32'h44ba68e4, 32'h43fe821e, 32'h439cc20d},
  {32'hc3fca5f5, 32'h431884de, 32'h43365f4a},
  {32'h44d2ee73, 32'h437f6460, 32'h42eb192e},
  {32'hc4f369e4, 32'hc2eb3b3b, 32'h43c0d12f},
  {32'h45282963, 32'hc3469f59, 32'h4327eb22},
  {32'hc4342314, 32'h437d81f7, 32'h43c712a0},
  {32'h44b897f3, 32'h3d66aaee, 32'h41f41ce9},
  {32'hc3d8fd3e, 32'h44067046, 32'hc342db92},
  {32'h4401833c, 32'hc33e8a0c, 32'h42a0c482},
  {32'hc39a3384, 32'h427f7d3d, 32'hc40b90d7},
  {32'h44376408, 32'hc3ebaef9, 32'h441a1860},
  {32'hc354d600, 32'h4404fd2a, 32'hc3212053},
  {32'h45142059, 32'h436075fe, 32'h42bcee41},
  {32'hc4ac1525, 32'h421a0878, 32'h437ec43d},
  {32'h447f125c, 32'hc424b429, 32'hc3b3f681},
  {32'h431ee0e0, 32'h4364158c, 32'h43745980},
  {32'h440f9d4c, 32'h434e37cc, 32'hc3cafbf7},
  {32'hc4659a1e, 32'h422fdc83, 32'hc391f9a1},
  {32'h447331e4, 32'h437ee6da, 32'h419b08b4},
  {32'hc47badee, 32'h43210704, 32'h425dc070},
  {32'h441af598, 32'hc3267f78, 32'h430f7edb},
  {32'hc4e4930c, 32'hc3ba548d, 32'hc0c48b6c},
  {32'h4489e5b4, 32'h4285188a, 32'hc189e0cc},
  {32'hc50a5900, 32'h4209e543, 32'h42888626},
  {32'h449ab9a1, 32'h422361df, 32'hc3650879},
  {32'hc2fbd260, 32'h414cf70e, 32'hc3009628},
  {32'h443c9abc, 32'hc3b1c769, 32'hc3400db2},
  {32'hc50389ae, 32'h4235a874, 32'h4209400d},
  {32'h44a1ac2d, 32'hc309aa99, 32'hc0f1c09f},
  {32'hc4d1b693, 32'hc2c00ceb, 32'h40aeb0db},
  {32'h448253aa, 32'h42befb64, 32'hc375a7d7},
  {32'hc3a6953c, 32'h433a5925, 32'h43a83f16},
  {32'h4515259d, 32'h43385868, 32'hc3a6355c},
  {32'h433554fb, 32'h424ea966, 32'h43c58534},
  {32'h44b650f7, 32'h431294c9, 32'hc2a722f4},
  {32'hc4831fba, 32'hc2a4a653, 32'hc331ffb7},
  {32'h43448990, 32'h42b964c8, 32'hc313fd9e},
  {32'hc4481c18, 32'h41bc64b8, 32'hc31c52d7},
  {32'h44f03575, 32'h42a167de, 32'hc1a2daa0},
  {32'hc3db8635, 32'hc30c0556, 32'h41a5086e},
  {32'h434717c2, 32'h439e415a, 32'hc3d6c0c4},
  {32'hc48312fa, 32'h439e6b80, 32'h41e95306},
  {32'h44ff53d4, 32'h426c83b8, 32'hc32951bd},
  {32'hc3253d2c, 32'h43105289, 32'h4376c0a4},
  {32'h445801a3, 32'h439a1ead, 32'h435224b8},
  {32'hc4ff7b1c, 32'hc1c59856, 32'h42aedd94},
  {32'h449bcfa9, 32'hc218bd28, 32'hc2ce13c2},
  {32'hc502c3a5, 32'hc2f6569d, 32'h428f1ea9},
  {32'h441407ea, 32'h41836299, 32'h4361f51d},
  {32'hc4a6d754, 32'hc3577823, 32'h43e2be6e},
  {32'h445915d4, 32'h4262ab48, 32'h426c0ff3},
  {32'hc3a91410, 32'h43cdded6, 32'hc2cdcf82},
  {32'h44ba113f, 32'h431c4544, 32'hc2c49436},
  {32'hc4fb34d8, 32'hc23910c2, 32'h43192ed5},
  {32'h449f53fb, 32'h41cb90a8, 32'h42533bf4},
  {32'hc5116e45, 32'h42febe6d, 32'h4250dbe7},
  {32'h44c9539c, 32'h42bb8450, 32'hc299b441},
  {32'hc4da4cae, 32'hc2ea7468, 32'h42eb7506},
  {32'h439f3f21, 32'h405527eb, 32'hc25c49e7},
  {32'hc481eacb, 32'hc298a6e5, 32'hc33bd94c},
  {32'h4490b41c, 32'hc12c4cb1, 32'hc3c8e34c},
  {32'hc3d202c0, 32'hc2d66ff8, 32'h43a68d4c},
  {32'h44d7cf3d, 32'hc25956f2, 32'h3e7a2e00},
  {32'hc3b6d124, 32'hc28c4e5c, 32'h43b32d63},
  {32'h450d1ed2, 32'hc282ff8a, 32'hc3813d9b},
  {32'hc4db1a86, 32'h435e7f67, 32'h42934bbb},
  {32'h43127c30, 32'hc398245a, 32'h43c5cb7c},
  {32'hc4c46f64, 32'h431af577, 32'hc318eee0},
  {32'h448e57f6, 32'h42d90dce, 32'hc3d7f857},
  {32'h44b46bee, 32'hc2e6aa6c, 32'h4335ccee},
  {32'hc4b57bf0, 32'hc1dba405, 32'h42411c02},
  {32'h44d0794f, 32'hc36d0574, 32'hbf82dc54},
  {32'hc419406e, 32'hc3a14cf2, 32'h43a0e72b},
  {32'h44c8814d, 32'hc335fe48, 32'hc29a138d},
  {32'hc4d89684, 32'h4394d3ba, 32'h438976eb},
  {32'h44c74140, 32'hc352a370, 32'h419ce1e1},
  {32'hc5188ed4, 32'hc2080712, 32'h422e8fb6},
  {32'hc15be200, 32'h42a42def, 32'h430c989b},
  {32'hc435045a, 32'h44078d60, 32'h434f1522},
  {32'h432e7880, 32'h4214a433, 32'hc39f61c5},
  {32'hc4246774, 32'h428bbf7a, 32'h438eece3},
  {32'h443fe851, 32'h41acf018, 32'hc23d08d3},
  {32'hc334ed20, 32'hc38d77a4, 32'h423f7106},
  {32'h42c64fe0, 32'hc2fab7c8, 32'hc2d17784},
  {32'hc516fc76, 32'hc34f4c9e, 32'hc29ade64},
  {32'h44afd48e, 32'hc3009ba4, 32'hc330b292},
  {32'hc448399e, 32'h432f11d2, 32'h43068974},
  {32'h4489f261, 32'hc3bfb8fd, 32'hc344724b},
  {32'hc398bd68, 32'h434a3633, 32'hc273912e},
  {32'h44c80fdf, 32'h42bf48eb, 32'hc344fd37},
  {32'hc3e12e2a, 32'h4336007f, 32'h437b6cca},
  {32'h44d90da6, 32'h435725ba, 32'hc3af9714},
  {32'hc4b49c46, 32'h430f922f, 32'hc1cc1721},
  {32'h446d1f8a, 32'hc38b4ade, 32'hc30f6fe6},
  {32'hc3807750, 32'h4381902d, 32'h43f07b8f},
  {32'h446fb8d0, 32'h433600e4, 32'h4283d789},
  {32'hc1f24980, 32'hc33ed3b7, 32'hc2b36be1},
  {32'h45066fe6, 32'hc1f44940, 32'hc3c2459d},
  {32'hc0578d00, 32'h428af8d5, 32'h42426071},
  {32'h449210ce, 32'h426a71c4, 32'hc37a8a75},
  {32'hc4f003dc, 32'h428035dd, 32'hc3348563},
  {32'h43483db4, 32'h4204702d, 32'hc1b2bfd6},
  {32'hc3cb196e, 32'hc3a3c1da, 32'h421b790d},
  {32'h42e969bb, 32'h41b770e8, 32'hc30c3703},
  {32'hc3b2aa0a, 32'h4067ef4d, 32'hc2ab82f7},
  {32'h450ac8e1, 32'hc311542d, 32'h42dcf5f1},
  {32'hc4e5c8b6, 32'hc322e28a, 32'hc297059e},
  {32'h44f4e6f3, 32'h43f34795, 32'h4337aafb},
  {32'hc4dc2243, 32'h42d67471, 32'h4344115c},
  {32'h43fe72c9, 32'h43438f7b, 32'hc26c3a1b},
  {32'hc4e78028, 32'h430ffc3c, 32'h42d4b4ba},
  {32'h43e82716, 32'hc3bad33d, 32'hc211d8c0},
  {32'hc5162f46, 32'hc148dec0, 32'hc3f544db},
  {32'h44d29c0a, 32'hc2bbc62c, 32'h433bcda8},
  {32'hc3c419de, 32'hc2d7aa8c, 32'h42d72be9},
  {32'h44bc1864, 32'h427dfc84, 32'h437c0574},
  {32'hc49bb869, 32'h4357f536, 32'hc3a87f00},
  {32'h44cfe026, 32'hc2a75939, 32'h43a8e4ff},
  {32'hc4ba5028, 32'hc342a95d, 32'h42138614},
  {32'h44054bb0, 32'h434fddf4, 32'hc3c9f6e4},
  {32'hc38a46a2, 32'hc37a6e6c, 32'h440eb372},
  {32'h4436eccc, 32'h41f8bfb2, 32'h43536521},
  {32'hc49e2c35, 32'h40b84d85, 32'h437fd97f},
  {32'h44915155, 32'hc3b2abc5, 32'hc35d56e1},
  {32'hc48e49df, 32'hc3bab678, 32'hc2863481},
  {32'h4496157e, 32'hc329c38e, 32'hc35ccb08},
  {32'hc4999cc0, 32'hc256124c, 32'hc2c7e7fa},
  {32'h44d9411e, 32'hc40b2eda, 32'h43f5536c},
  {32'h429526a0, 32'hc3468ef9, 32'hc33b8b14},
  {32'h44f3ceb0, 32'hc32e3593, 32'h4374717f},
  {32'hc4fd543c, 32'h441f6d85, 32'hc249005f},
  {32'h42ded860, 32'hc2f00b5c, 32'hc3a5aaaa},
  {32'hc3dba264, 32'hc2a3792e, 32'hc35c1e20},
  {32'h447fbc24, 32'hc2fa2d34, 32'h4294da95},
  {32'hc2debd48, 32'h4219d66e, 32'hc371799f},
  {32'h44f54866, 32'h431aec38, 32'hc4039c00},
  {32'hc4d397ff, 32'hc3b0032d, 32'h43a05d5c},
  {32'h42c67280, 32'hc34dabd9, 32'h434bb071},
  {32'hc3deb0de, 32'hc3c4932f, 32'h42a33b89},
  {32'h4513bc99, 32'h41c23120, 32'hc2c25d1e},
  {32'hc515c7bd, 32'hc28ce360, 32'h439cb053},
  {32'h42a3d0f0, 32'h43374869, 32'hc306ee69},
  {32'hc4e82a54, 32'hc305d52f, 32'h410c6fd6},
  {32'h44cfb674, 32'hc34cac42, 32'hc37242bf},
  {32'hc4f1fd58, 32'hc3ddc542, 32'h42fc9f57},
  {32'h4495e101, 32'hc3988d00, 32'hc3d9bd7c},
  {32'hc4dda7b5, 32'h43027f3b, 32'hc353a8d0},
  {32'h43cf8c88, 32'h4396c67d, 32'hc36dde3f},
  {32'hc15fa175, 32'h43bad533, 32'h423f4800},
  {32'h4512e564, 32'hc354c2c2, 32'hc2c68fb2},
  {32'hc43418b4, 32'h416d8798, 32'h426a18fe},
  {32'h43c20c44, 32'hc3d13505, 32'h42746d2f},
  {32'hc44bec97, 32'hc2884756, 32'hc286ed17},
  {32'h449f0ca9, 32'h42aac36f, 32'h421ac39b},
  {32'hc5030efc, 32'h41ea4273, 32'h43f28e0a},
  {32'h4515cc8c, 32'hc1b6c767, 32'hc2905f4e},
  {32'hc4fe0b09, 32'hc33b5ce9, 32'hc34ee4d2},
  {32'h43cd04e4, 32'hc0a2238a, 32'hc36d3f2f},
  {32'hc4b3cc6e, 32'hc2110652, 32'h440e9ee6},
  {32'h448b867a, 32'hc348271b, 32'h43998a39},
  {32'hc5089eee, 32'h434cc1b4, 32'h431e0f47},
  {32'h449bba12, 32'hc2b46304, 32'hc2f9cfe9},
  {32'hc508ffca, 32'hc353be46, 32'h4256c882},
  {32'h4462b0be, 32'h42286740, 32'h437aafdc},
  {32'hc41e1b1c, 32'hc3714d09, 32'hc13664cc},
  {32'h43b9b684, 32'h431de9ad, 32'h42f9c70e},
  {32'hc494a370, 32'h439017cf, 32'hc21a59ce},
  {32'h4460abe7, 32'h42a94326, 32'hc23ea48c},
  {32'hc44277ca, 32'hc24f2586, 32'h43c9156e},
  {32'h4372ef30, 32'h427a6350, 32'h433be020},
  {32'hc4fde67a, 32'h42ddb379, 32'h434fda18},
  {32'h451917b1, 32'hc25661e8, 32'h41ef8c7b},
  {32'hc4de8d0a, 32'hc38b3751, 32'h42d9a1d4},
  {32'h44d9f40f, 32'hc3e37b7d, 32'h43106175},
  {32'hc510a66c, 32'h43896ff9, 32'hc3428f39},
  {32'h45102d4b, 32'h42bbc9bb, 32'hc38e3702},
  {32'hc498b9f3, 32'h4262520d, 32'hc30f01f4},
  {32'h44055bc4, 32'h40c04284, 32'hc313da17},
  {32'hc4d48676, 32'hc2ce541f, 32'h432b3408},
  {32'h44a2306e, 32'h423715d8, 32'hc2cb85d0},
  {32'hc4b089f8, 32'hc3061acb, 32'hc28b824c},
  {32'h43ff80c6, 32'hc3bf5bbf, 32'h4254a713},
  {32'hc3a09ed0, 32'h4402d0d0, 32'h424c17ce},
  {32'h448c018c, 32'h42b4ad4b, 32'hbf494910},
  {32'hc4d7bde1, 32'h438d5291, 32'h41dfe986},
  {32'h4492f2be, 32'h424afa9a, 32'hc30423c9},
  {32'hc487d7a7, 32'hc183c631, 32'h4254523b},
  {32'h4507d324, 32'h438abeae, 32'h4318a91b},
  {32'hc4e19334, 32'hc2ebbba9, 32'hc3635b0e},
  {32'h44c6d7cb, 32'hc0725ce0, 32'h4365b961},
  {32'hc376e280, 32'h40d5c150, 32'h42467086},
  {32'h441c067a, 32'h43c49ca5, 32'h431fd43f},
  {32'hc424c8a9, 32'h4363e7fb, 32'hc368dddb},
  {32'h44eaddd1, 32'h43600b5c, 32'hc38b6a0a},
  {32'hc4fbca2a, 32'hc2c30ad5, 32'hc2ca6847},
  {32'h44255e96, 32'hc3369278, 32'hc359ef79},
  {32'hc4d63641, 32'h43998cbe, 32'h42968443},
  {32'h4426a598, 32'hc373e864, 32'h431b6c70},
  {32'hc4f6be63, 32'hc319fba6, 32'h43868c82},
  {32'h44c266eb, 32'h4401817b, 32'hc34dffdc},
  {32'hc429ca92, 32'h41ecab5b, 32'hc099d464},
  {32'h4464add0, 32'h43de9d53, 32'h43823a16},
  {32'hc50315f9, 32'hc32e7d6d, 32'hc363f2c6},
  {32'h451c49b4, 32'h423900b6, 32'hc3a445fc},
  {32'hc3b33bf4, 32'hc31ce5bd, 32'hc3430e4c},
  {32'h44d18c74, 32'h426939ea, 32'h43c4aead},
  {32'h422c7480, 32'hc3df765a, 32'h43cc0ac6},
  {32'h44f02bc2, 32'h4335c0ee, 32'hc2d98cdd},
  {32'hc4b604bd, 32'h3ff437d4, 32'h43d5c771},
  {32'h44faf857, 32'hc2e54762, 32'hc1833a22},
  {32'hc4b39bf2, 32'hc2778e57, 32'h42240323},
  {32'h44e12dea, 32'hc2aec942, 32'hc2894a21},
  {32'hc4624cf3, 32'hc3bd5bce, 32'hc37f12b8},
  {32'h4513176d, 32'h419a6907, 32'h4323959e},
  {32'hc4ab49e0, 32'hc39c7b7e, 32'hc348bed4},
  {32'h44d3a35d, 32'h43a64212, 32'hc33a3ae6},
  {32'hc36f9334, 32'h43b62e05, 32'h43010cf8},
  {32'h43a35950, 32'hc33f25c8, 32'hc2cef18e},
  {32'hc4a2f156, 32'h434b0c2e, 32'h42488442},
  {32'h443ca1e6, 32'h43854858, 32'h424f5fd3},
  {32'hc49ef1d3, 32'h42291651, 32'hc2982fd6},
  {32'h4502fdb7, 32'hc3b8542b, 32'hc2a702ba},
  {32'hc43b6370, 32'hc3611799, 32'h423ed054},
  {32'h43a6e114, 32'h423627f5, 32'h438bc4e8},
  {32'hc501b509, 32'hc2ca0a7f, 32'h417dc28b},
  {32'h44c7a64d, 32'h43736146, 32'hc306dc66},
  {32'hc51708c0, 32'h43654093, 32'hc3866f30},
  {32'h44c7a5af, 32'h439611fc, 32'hc31f8437},
  {32'hc461555c, 32'h43090fed, 32'h42a9e51d},
  {32'h44daae41, 32'h434dd060, 32'h42b4088d},
  {32'hc46cd2ba, 32'h42ebb7cf, 32'h43819ad7},
  {32'h448ae6d4, 32'hc28ce3d9, 32'hc38c6003},
  {32'hc3a0991c, 32'hc3824651, 32'hc1b133d2},
  {32'h448d4fec, 32'hc33f9608, 32'hc386bd49},
  {32'hc49b69c7, 32'hc265afa2, 32'hc2e85cfe},
  {32'h451986ed, 32'h4280dfd7, 32'h42b2b2b1},
  {32'hc2a6a6a0, 32'hc28d81d5, 32'hc340a7eb},
  {32'h4510e486, 32'h431eb6c8, 32'h4205bb3b},
  {32'hc49e74eb, 32'hc310eadb, 32'hc2decf34},
  {32'h44d51bb7, 32'hc3725d0b, 32'hc4115498},
  {32'hc49bab8d, 32'hc27b31f6, 32'h43adf0aa},
  {32'h441a8836, 32'h4296c13a, 32'h4352c4a6},
  {32'hc506491c, 32'h42ea708e, 32'hc3aaa9fd},
  {32'h4319d9f2, 32'hc238eeda, 32'hc342ad1b},
  {32'hc4b9547a, 32'h4353c7dc, 32'h43d168e7},
  {32'h438c8fdc, 32'hc1472d2c, 32'h430e190b},
  {32'hc4f510e8, 32'hc24a07e1, 32'hc2b1c68f},
  {32'h45120efe, 32'h42f0fb6d, 32'h42bcdd40},
  {32'hc4ccaacc, 32'hc1abda38, 32'hc2ead73b},
  {32'h44d6ca7f, 32'hc3ef1490, 32'hc29f5026},
  {32'hc311e908, 32'hc382ee8c, 32'hc377b36d},
  {32'h43128b14, 32'hc3db7e65, 32'hc3331e1d},
  {32'hc4a0a637, 32'hc2477d70, 32'h4307c9de},
  {32'h44160d17, 32'hc3aaa922, 32'h42d26246},
  {32'hc4d44898, 32'h43436dfc, 32'h43530621},
  {32'h44bd530a, 32'h424e1c53, 32'hc38f377f},
  {32'hc4fc902c, 32'h43216b8b, 32'hc3381046},
  {32'hc0b87a00, 32'hc345bd0c, 32'hc1ee76b2},
  {32'hc4de2478, 32'hc16986b3, 32'h4382283a},
  {32'h449a9e68, 32'hc35edd6d, 32'h42eadae2},
  {32'hc4917fa3, 32'h43a37a4f, 32'hbff63918},
  {32'h434b29a1, 32'hc33ba309, 32'h421b920b},
  {32'hc4b686d0, 32'hc361ee6b, 32'h42ca9b2a},
  {32'h4433e438, 32'hc3b4c8a9, 32'hc1fe5be6},
  {32'hc487cc6a, 32'h430822a1, 32'hc381509f},
  {32'h44f6c481, 32'h42acf210, 32'h430671fa},
  {32'hc487b4b5, 32'hc30678c0, 32'hc38f4c06},
  {32'h4499efb3, 32'h428223ab, 32'h4328ceeb},
  {32'hc23b3280, 32'hc3643d6a, 32'hc21a5200},
  {32'h43a0cd5a, 32'hc3078ec4, 32'hc301d8f3},
  {32'hc3bca940, 32'hc302e58a, 32'h430c8d00},
  {32'h448749b7, 32'hc368b523, 32'h434ab2b4},
  {32'hc4ff6717, 32'h427649bc, 32'h438b5180},
  {32'h44e9f352, 32'hc40ecf4c, 32'h43d54bc6},
  {32'hc51bde86, 32'h42be6e5b, 32'h42f357c7},
  {32'h41d3cb00, 32'hc33cc23c, 32'h4290b913},
  {32'hc4b091e9, 32'h434f1512, 32'hc3b2c970},
  {32'h44ba87a8, 32'hc2dfc84f, 32'h430c3d13},
  {32'hc3dddb78, 32'h420d234e, 32'hc29d3c70},
  {32'h44e088e6, 32'hc3465997, 32'hc1811b6d},
  {32'hc3a2abd4, 32'hc3bfeab2, 32'hc01437a5},
  {32'h446e40d9, 32'h435c7786, 32'h434e9148},
  {32'hc2491dc0, 32'hc3c0fed9, 32'h43957bb3},
  {32'h44ecb86e, 32'hc3ecad68, 32'h43973274},
  {32'hc46b1384, 32'hc318babd, 32'h42a9ee42},
  {32'h43806b10, 32'h4281e5fa, 32'hc2f47163},
  {32'hc4f26720, 32'hc24fdc28, 32'hc1956a0e},
  {32'h44d05ea2, 32'h4367f574, 32'hc2d21e08},
  {32'hc4f5b8bf, 32'h43b3eeab, 32'h4387f351},
  {32'h44c31bb5, 32'h431b9957, 32'h4238c5fa},
  {32'hc4bae88f, 32'h42a4fb28, 32'h4330e798},
  {32'h44689db2, 32'h435f12c3, 32'h4319d904},
  {32'hc4124c20, 32'hc384993e, 32'hc2fe856a},
  {32'h44920f0a, 32'h43f61968, 32'h417cead4},
  {32'h43361110, 32'h431d85c4, 32'hc1edceed},
  {32'h451c326a, 32'h43c67241, 32'hc14aac7d},
  {32'hc375f211, 32'hc31dee98, 32'hc2f06368},
  {32'h4405fbbf, 32'hc3945cc5, 32'hc2bb2f03},
  {32'hc47ae0a3, 32'hc0390f53, 32'hc2995b38},
  {32'h44242752, 32'h43445699, 32'hc2044f89},
  {32'hc4b2a44a, 32'h42bc0fbb, 32'hc2ffb35c},
  {32'h44e2c012, 32'h421a92ad, 32'h42a7efc5},
  {32'hc5040450, 32'hc3014626, 32'hc31dcb9f},
  {32'h4500f5ad, 32'h4155190b, 32'h42ac07eb},
  {32'hc4b8c733, 32'hc2809cd5, 32'hc353c355},
  {32'h44f4eb68, 32'hc363bd2a, 32'hc28910d4},
  {32'hc37696f5, 32'h43451c46, 32'h42d721c6},
  {32'h44801196, 32'hc2069868, 32'h430a0c44},
  {32'hc3e70311, 32'hc202f3b6, 32'h42d2639d},
  {32'h437b53d2, 32'hc21ab99a, 32'h4345856e},
  {32'hc4d83f27, 32'h430bb2db, 32'hc3a86e58},
  {32'h448c009f, 32'hc1dfce36, 32'h42331600},
  {32'hc494fd64, 32'h430b63fe, 32'h4320e7fb},
  {32'h445b12de, 32'h437d2203, 32'hc2f86620},
  {32'hc38c6420, 32'h42fa31b6, 32'hc33aecb6},
  {32'h4419ef2a, 32'hc3034ba6, 32'hc2ae32a3},
  {32'hc27bad60, 32'hc15b2bef, 32'hc33cd5da},
  {32'h42b7c7b8, 32'h42817b39, 32'h430fe27d},
  {32'hc4b1902a, 32'h42f0dd0e, 32'hc3491117},
  {32'h44839d8a, 32'hc2ae974f, 32'hc3a25547},
  {32'hc500e12f, 32'hc297f3fc, 32'h437caf04},
  {32'h43f37850, 32'h430a547f, 32'hc328756e},
  {32'hc4e5ccd6, 32'h43a1eb16, 32'hc2d79e6f},
  {32'h444c61ce, 32'h42555764, 32'hc36b1f3a},
  {32'hc4e58820, 32'h4396960b, 32'hc358934f},
  {32'hc3310147, 32'hc3305fe2, 32'h4320c940},
  {32'hc3763ee8, 32'hc1cf3c97, 32'h4324c996},
  {32'h446d389c, 32'h42b4f45e, 32'hc197422c},
  {32'hc4ab89df, 32'hc2b5dc7c, 32'h43a09ae6},
  {32'h42ed2de8, 32'h43036179, 32'hc10e8074},
  {32'hc4c0401a, 32'h4356be0a, 32'h437f92e9},
  {32'h44bc0993, 32'hc225cd6e, 32'h41d48df9},
  {32'hc2d7e23c, 32'h408b0be6, 32'h42304144},
  {32'h44f6fd2b, 32'h42d50be8, 32'hc390b71d},
  {32'hc4a819b2, 32'hc20a1b78, 32'h43a566ca},
  {32'h44e5c642, 32'h43f3d3a3, 32'h41ff2f39},
  {32'hc4e6ea80, 32'hc3437c6b, 32'h439c3214},
  {32'h44f5ce92, 32'h4337a400, 32'hc38a4c33},
  {32'hc502f6f2, 32'h43882a9f, 32'hc302cb40},
  {32'h44d9ec6e, 32'h42bd69f0, 32'h43294732},
  {32'hc4d86903, 32'h42521607, 32'h43810606},
  {32'h44fd88c9, 32'hc3044b72, 32'hc2dec287},
  {32'hc4e0fca9, 32'h430b2ba9, 32'hc20f81ae},
  {32'h44bd1116, 32'hc3c5b1c8, 32'h432579e9},
  {32'hc512be7c, 32'hc36d7ecb, 32'h430f72b0},
  {32'h44f9e626, 32'hc34c38e3, 32'h427fbbe0},
  {32'hc44e0cf2, 32'hc0dbef48, 32'h42d8e207},
  {32'h44594766, 32'h438f2df5, 32'h3fdbb1ec},
  {32'hc4759b67, 32'hc22960c2, 32'hc3af70be},
  {32'h444d32ee, 32'hc3a4e8fe, 32'h439b18c1},
  {32'hc5164f35, 32'h4326fbc5, 32'hc2c11d48},
  {32'h45066f99, 32'hc313d947, 32'hc274ae98},
  {32'hc414395a, 32'h431a378a, 32'h4319b5b4},
  {32'h44408029, 32'h42c4ebb4, 32'hc1def476},
  {32'hc4dc9072, 32'hc33776c3, 32'hc246091f},
  {32'h44a70e78, 32'h42a0341f, 32'hc1bec280},
  {32'hc3931718, 32'h4276f94d, 32'h435cc5dc},
  {32'h44bae3be, 32'hc39747b3, 32'hc3b7776a},
  {32'hc4f1cfc1, 32'hc33859a7, 32'hc3c9b42a},
  {32'h4382db6e, 32'h42bb1441, 32'h41accad3},
  {32'hc4a11583, 32'hc1725f90, 32'hc26cd98a},
  {32'h44cd7564, 32'hc2c7a582, 32'h42c6e183},
  {32'hc4f25353, 32'h4230983c, 32'h4319be9d},
  {32'h44e23f29, 32'hc34d5b22, 32'h42f1f879},
  {32'hc484a3b7, 32'hc35d2b1f, 32'h43b45092},
  {32'h43f2b0f0, 32'h42d575f8, 32'h43423f5e},
  {32'hc4127c93, 32'h43958af9, 32'h42955105},
  {32'h44ae049c, 32'hc0143168, 32'hc33f91db},
  {32'hc507c5de, 32'hc335d16d, 32'h421691c0},
  {32'h449f3edb, 32'h42dc1a7c, 32'hc2e909cf},
  {32'hc4ff432e, 32'hc3825414, 32'h4396afae},
  {32'h446ac88c, 32'h43c511fb, 32'h424948a8},
  {32'hc4b921c0, 32'h42a564ae, 32'h42874f2e},
  {32'h451989d9, 32'h431ba477, 32'hc396f52b},
  {32'hc4ef4eb2, 32'hc32d4712, 32'h43c21550},
  {32'h436057d0, 32'h4274d48a, 32'hc28db27e},
  {32'h42e38e48, 32'hc363b914, 32'h4169c3ac},
  {32'h44d55a3a, 32'hc3bc2a46, 32'hc2831b84},
  {32'hc509dee6, 32'h4106a29e, 32'h43026d04},
  {32'h44fb3e48, 32'hc397c5be, 32'hc3db459a},
  {32'hc4cff8a6, 32'h42525f38, 32'h42637577},
  {32'h450d88a5, 32'hc3a1df9f, 32'hc2a964ff},
  {32'hc509144d, 32'h4280edc2, 32'hc33cc558},
  {32'h44f950b8, 32'hc37f8a5e, 32'hc374472c},
  {32'hc487fc11, 32'hc1ffb1e4, 32'h435ddf01},
  {32'h44c83052, 32'hc087f744, 32'hc2d9c2f2},
  {32'hc52712d8, 32'h4212a9b3, 32'h42cdf8cf},
  {32'h43866f78, 32'h43c34658, 32'hc3894b89},
  {32'hc4ef60f3, 32'hc354f8d4, 32'hc3b20ae1},
  {32'h441caa84, 32'hc2c74455, 32'h4212bc3a},
  {32'hc5024faa, 32'h43420deb, 32'h42bc992d},
  {32'h44fc8a01, 32'h438dd632, 32'h4325d441},
  {32'hc49dbf64, 32'hc3a52c11, 32'hc016caea},
  {32'h44b12a83, 32'hc3c8cfbc, 32'hc33a8cd6},
  {32'hc463ea2a, 32'h40b13100, 32'h43c05744},
  {32'h44e5aac9, 32'h43e03722, 32'h437f4e70},
  {32'hc4e4455c, 32'hc3338da2, 32'h430fdbde},
  {32'h445a90de, 32'hc3fead26, 32'hc3c42b12},
  {32'hc3f24080, 32'h43e0bf4b, 32'hc2bd4a5d},
  {32'h44e29e42, 32'hc3254489, 32'h43076b70},
  {32'hc4dac4c9, 32'h43346444, 32'hc37a8776},
  {32'h44012a6e, 32'hc2ee6837, 32'hc2062765},
  {32'hc414a682, 32'h427ad9a7, 32'h43995108},
  {32'h44aa5d97, 32'h436d521b, 32'hc2df9bea},
  {32'hc51cb69b, 32'hc3760e93, 32'hc30a62fb},
  {32'h450aa4e6, 32'hc15e024a, 32'hc260aebb},
  {32'h42843a40, 32'h421fe558, 32'hc35e1be0},
  {32'h44c4707d, 32'h416f8ffc, 32'hc309cd73},
  {32'hc4db7eee, 32'hc1c8553c, 32'hc12ce0a8},
  {32'h44f8692a, 32'hc3460eb9, 32'h433c3ed2},
  {32'hc4587e56, 32'h444686b9, 32'hc385c2d6},
  {32'h451804d5, 32'h43814b60, 32'hc2edcc29},
  {32'hc4e9f1f5, 32'hc3347ff2, 32'hc3d45e7e},
  {32'h451694b6, 32'h42926b3b, 32'hc3933e47},
  {32'hc467e3c2, 32'h412a8968, 32'hc3317de8},
  {32'h4507a201, 32'hc330a0fd, 32'h434cda97},
  {32'hc4b5f4ea, 32'hc2dd6572, 32'hc29da3eb},
  {32'h445905ac, 32'hc43b3d07, 32'h42a7eef8},
  {32'hc4149b74, 32'h43c43c42, 32'hc3df12ee},
  {32'h44446c2b, 32'hc2e84462, 32'hc3e5d2cd},
  {32'hc513dc92, 32'hc3aca922, 32'hc33a2f6f},
  {32'h44dee40f, 32'h419b3674, 32'h43598787},
  {32'hc4f8d912, 32'hc2ca1080, 32'hc316abf2},
  {32'h451a29d5, 32'hc41446a2, 32'hc29ca3bc},
  {32'hc41108de, 32'hc33eaf78, 32'hc38543ee},
  {32'h4500717f, 32'h436624cb, 32'hc334e1f8},
  {32'hc4cbb7b5, 32'h43899581, 32'hc33e18c1},
  {32'h4495d6f5, 32'h420ac23f, 32'h43c76b5c},
  {32'hc4adf716, 32'hc115005d, 32'hc3a894e4},
  {32'h43c149e0, 32'hc245b966, 32'hc359ccd6},
  {32'hc48495e0, 32'h432860b2, 32'h439d90cb},
  {32'h4449ced4, 32'hc23c508c, 32'h42823765},
  {32'hc4842a6d, 32'hc298a9a1, 32'hc3a7259f},
  {32'h44c230c6, 32'hc3be0152, 32'h42b20f39},
  {32'hc4c9b4bc, 32'h42d3fd92, 32'h43337e8a},
  {32'h45040d32, 32'hc3c6e905, 32'h43f53c3c},
  {32'h431bcbe0, 32'h4327163e, 32'hc3f9ffcf},
  {32'h44deda40, 32'hc32f915f, 32'hc303dd68},
  {32'hc482e798, 32'h43e21ead, 32'h43555666},
  {32'h44d5d85c, 32'h43a781c8, 32'hc3ade275},
  {32'hc40707e8, 32'h41ff333d, 32'hc3c772c3},
  {32'h4512f564, 32'hc288b9b2, 32'h417573b2},
  {32'hc4b2059b, 32'h435442ee, 32'hc26e9c2f},
  {32'h447771d5, 32'h442c6faf, 32'hc3808121},
  {32'hc3027500, 32'hc22000c8, 32'h40592890},
  {32'h4513d57f, 32'hc24f5c7a, 32'hc2cd666b},
  {32'hc4c0bcee, 32'h4298507f, 32'h434a4d3b},
  {32'h4401ddd0, 32'h438681c6, 32'hc304a556},
  {32'hc4b6e669, 32'h4345b9bc, 32'h42c0da9e},
  {32'h44c1eb8c, 32'h43dc1228, 32'h428656d4},
  {32'hc48917b0, 32'h4291edfb, 32'hc29439c5},
  {32'h452cdbf0, 32'hc3166fa2, 32'hc2d64084},
  {32'hc443fd2e, 32'h4327c2cf, 32'hc3b51db7},
  {32'h45023174, 32'hc3167bc6, 32'h430f9f49},
  {32'hc4e48131, 32'h43120624, 32'h408952e4},
  {32'h4486af29, 32'hc305a8f4, 32'hc21bfaa3},
  {32'hc4b4fc0c, 32'hc38f709a, 32'h4398b81d},
  {32'h44b81b7d, 32'hc019de46, 32'h41ceb832},
  {32'hc4d8163b, 32'h4332b70d, 32'h4388e91f},
  {32'h44cb5dbe, 32'h43951d93, 32'hc1fe3c10},
  {32'hc4b260c6, 32'hc1939990, 32'h434de80e},
  {32'h44adee58, 32'h42d141af, 32'hc3104ee4},
  {32'hc2ec61e0, 32'h42bb373a, 32'hc3ba7671},
  {32'h45056dfe, 32'h427ede2f, 32'h439344df},
  {32'hc4a16597, 32'hc40eb622, 32'h433d88c9},
  {32'h44b4ebd6, 32'h40de3342, 32'h436cdbb3},
  {32'hc4de17a2, 32'hc39b6ead, 32'h425a23e8},
  {32'h448fab28, 32'h4297a923, 32'hc34eb939},
  {32'hc379cd9c, 32'h43947163, 32'hc38b7f3d},
  {32'h44a3deff, 32'hc2fade94, 32'h437c1aad},
  {32'hc418bab7, 32'h4402661b, 32'hc3adf7d1},
  {32'h443425e8, 32'hc2cd932c, 32'h43113aac},
  {32'hc4cd8174, 32'hc3c8cdc2, 32'h4373407e},
  {32'h4433ea74, 32'hc3818493, 32'h43aafd6a},
  {32'hc40d827a, 32'h43f75981, 32'h431cd1f9},
  {32'h44d12023, 32'hc167c84f, 32'h4335b8c8},
  {32'hc4c1000d, 32'hc2638586, 32'hc3cbc0ec},
  {32'h4403a46d, 32'h42b7078e, 32'hc1d63174},
  {32'h432360e8, 32'hc3436fea, 32'h4316b08a},
  {32'h451adba9, 32'h42edb206, 32'h41f6633c},
  {32'hc49efaa6, 32'h430fdee4, 32'h42b4cefc},
  {32'h447782a9, 32'hc3ac9fd0, 32'h42d6a1f3},
  {32'hc49c1317, 32'h43227014, 32'hc3874bfa},
  {32'h4498ac04, 32'h43ade27d, 32'h43623c9d},
  {32'hc45fba70, 32'h43836c38, 32'hc28baab4},
  {32'h44b9534f, 32'h43528a32, 32'hc24d91e4},
  {32'hc37165f0, 32'hc2381bbb, 32'h425dbace},
  {32'h44f616ca, 32'hc2c2b01b, 32'hc2eac39d},
  {32'hc4e2f314, 32'h42787883, 32'hbdaea8d0},
  {32'h44d04cef, 32'hc35dacd7, 32'hc31bf3cc},
  {32'hc4c5cf7e, 32'hc2ba737d, 32'hc2e944a3},
  {32'h445fd40f, 32'hc297cdfa, 32'h42f368b8},
  {32'hc4031990, 32'h434eb73e, 32'h42f1d579},
  {32'h4415c8bb, 32'hc0ac2d13, 32'h43a3118f},
  {32'hc4a4405d, 32'hc2564a8c, 32'hc32c2396},
  {32'h445e6774, 32'h43517da1, 32'h438fd5d0},
  {32'hc444c64b, 32'hc281995c, 32'h4286c240},
  {32'h43f80a12, 32'h43916321, 32'hc2c0c37b},
  {32'hc4dff6ca, 32'hc2bc5367, 32'hc386ca88},
  {32'h4507b9ed, 32'hc2de09e8, 32'h42210406},
  {32'hc403bea4, 32'h435c641e, 32'hc3ae25ca},
  {32'hc4688460, 32'hc39a6114, 32'hc32d0f6d},
  {32'h432e69a4, 32'hc22c669a, 32'h42c37b49},
  {32'hc3c77e50, 32'h43f33435, 32'h431cf89c},
  {32'h42096800, 32'hc30f1429, 32'h435d0f6b},
  {32'hc45257a2, 32'hc39e0cbd, 32'hc30ee00e},
  {32'h4501f876, 32'hc3e2d25f, 32'h428145d3},
  {32'hc4dff574, 32'hc3ba0a19, 32'h439a3eb3},
  {32'h44704310, 32'h4333c55b, 32'hc32e4da0},
  {32'hc49fcd98, 32'h438c3a26, 32'hc36725b8},
  {32'h44aa9248, 32'h43a830eb, 32'h41760414},
  {32'hc39f5e9e, 32'h432a8cdd, 32'hc311d538},
  {32'h450a1f44, 32'hc22d58fd, 32'hc2a66664},
  {32'hc4581fdc, 32'hc342a43a, 32'hc17117e4},
  {32'h45087503, 32'h440563d9, 32'h43a8768c},
  {32'hc4ab1d42, 32'h42a8d024, 32'h429c6ddf},
  {32'h4499293f, 32'h42973c89, 32'hc27f1c7f},
  {32'h435ad740, 32'h41ddd206, 32'hc3ab1070},
  {32'h44a69c5e, 32'hc390f11a, 32'h42ae94d0},
  {32'hc3cdaa88, 32'h434e1a5b, 32'hc32c5812},
  {32'h44f77ebe, 32'h438fd9be, 32'h43200db9},
  {32'hc4a120e1, 32'h43fe61dc, 32'hc305a238},
  {32'h44e73cd4, 32'h435c6cdc, 32'hc148a8d6},
  {32'hc493ae67, 32'h439f29eb, 32'hc3428fc6},
  {32'h44064b04, 32'hc2bc2720, 32'h42967eaa},
  {32'hc3762890, 32'h41ffffce, 32'hc3c320c6},
  {32'h4482304a, 32'h42985075, 32'h4299ce91},
  {32'hc382a650, 32'h43616a36, 32'h4233f0fe},
  {32'h43cf16e0, 32'h4388d8df, 32'h43158b1b},
  {32'hc492162e, 32'h42a3cdf0, 32'hc3a28535},
  {32'h44b5f226, 32'h438cbe1e, 32'h43a147f9},
  {32'hc3b7be30, 32'h42b26b48, 32'hc2973214},
  {32'h44d828e6, 32'h42df76bc, 32'hc2a389f8},
  {32'hc4e23df6, 32'hc32cbef1, 32'h42fa3210},
  {32'h450c5f1e, 32'hc320e292, 32'h4393f2fc},
  {32'hc50b7978, 32'h43385ae1, 32'hc355a836},
  {32'h445383f7, 32'hc329f069, 32'hc2fe4ee0},
  {32'hc39ff8b0, 32'hc300917f, 32'h42dbd1c4},
  {32'h44e7507a, 32'hc2a6a461, 32'h42df74d0},
  {32'hc43f5ae9, 32'h42b4611a, 32'h42e27ec0},
  {32'h44e95dae, 32'hc37891e7, 32'hc1c7bffc},
  {32'hc50644cd, 32'hc21ae9d0, 32'hc3065a08},
  {32'h4507de6a, 32'hc38e41c2, 32'h43cad39a},
  {32'hc4b114bb, 32'h433583ef, 32'hc2d62a5e},
  {32'h449013e8, 32'h43c83e78, 32'h4411d5c4},
  {32'hc4c77cec, 32'h4388c4e1, 32'h43ad632b},
  {32'h450dd4b2, 32'hc15afb0a, 32'h433ae095},
  {32'hc4b81310, 32'h43d197dd, 32'hc3185fb4},
  {32'h44a57bd2, 32'h435d8bc2, 32'hc295af6c},
  {32'hc5021d5c, 32'h4302f95e, 32'hc35b47e0},
  {32'h4500635f, 32'h43d7642e, 32'hc3e14f7b},
  {32'hc3f3cfc4, 32'h40ae8c56, 32'h4254f6e6},
  {32'h4505bdfa, 32'hc2a20a7b, 32'h42f9067d},
  {32'hc3a463d2, 32'h426b6e0f, 32'hc40f80d8},
  {32'h445a3a70, 32'hc2ef6770, 32'h43e33a01},
  {32'hc401b558, 32'h43823b41, 32'hc3cf1608},
  {32'h444d99e3, 32'hc22975dd, 32'hc33324e9},
  {32'hc508f54b, 32'h4395da18, 32'hc35faab4},
  {32'h438a0704, 32'h4308ba48, 32'hc3284714},
  {32'hc4e30bbd, 32'hc2b0c168, 32'h41436688},
  {32'h4517451d, 32'hc2a1027a, 32'h43867ec7},
  {32'hc51a8182, 32'h42967fe0, 32'h43aa303d},
  {32'h44dc7950, 32'hc2096db0, 32'hc2174b88},
  {32'hc4a6b59c, 32'hc2ac3fe9, 32'h423d3fc9},
  {32'h436a2d4c, 32'h43707dd0, 32'hc2a9430c},
  {32'h4343dcd8, 32'h43b11789, 32'h431656cd},
  {32'h44bbb15a, 32'h429c9d69, 32'hc33f4dcf},
  {32'hc4be46f3, 32'h4366c5a0, 32'h434945c4},
  {32'h430ed771, 32'hc15e33b5, 32'hc28a5d66},
  {32'hc4be6484, 32'h43c68509, 32'hc3949d40},
  {32'h450da68a, 32'hc3496bfc, 32'hc384b7b4},
  {32'hc430dc70, 32'h42f8a8ce, 32'h43e23f7a},
  {32'h428f0310, 32'hc3a30b86, 32'h41f29015},
  {32'hc4e7e758, 32'hc39c516d, 32'hc3a70358},
  {32'h44fe34a0, 32'h433632be, 32'h432b2a40},
  {32'hc4e4b69f, 32'hc32f6368, 32'hc37f9dd1},
  {32'h4516897b, 32'hc2e1ce21, 32'hc1123b47},
  {32'h436b0185, 32'h42cd2d3a, 32'hc312cd09},
  {32'h450eb8ef, 32'h43a4c317, 32'h43d91099},
  {32'hc4fa7ffc, 32'h436f37e3, 32'hc1eb045a},
  {32'h44c37042, 32'hc41fc3f1, 32'h4427b533},
  {32'hc44b3914, 32'hc348d701, 32'hc314f30a},
  {32'h44a04f16, 32'hc1f24818, 32'h43cdc7b0},
  {32'hc2859ce0, 32'h437fd48a, 32'hc3543e89},
  {32'h44333256, 32'hc339766b, 32'h42ff63f7},
  {32'hc50e4a00, 32'hc35cde0e, 32'h42e0b464},
  {32'h442e99d4, 32'h434b5b49, 32'h4284fbfa},
  {32'hc4bf0f23, 32'hc181c851, 32'h4307ce66},
  {32'h43b60414, 32'h4304a72a, 32'h43df09bb},
  {32'hc4d4dc4d, 32'hc2b84701, 32'hc314767d},
  {32'h445ee504, 32'h43625a20, 32'hc322f1b8},
  {32'hc4cbc9c8, 32'h42010928, 32'hc18f7e40},
  {32'h4525d850, 32'h4169c713, 32'h432702df},
  {32'hc2f86c28, 32'hc22bf017, 32'hc2e8325b},
  {32'h44298704, 32'h438ffe71, 32'hc33ce8bf},
  {32'hc395e31c, 32'h4434c32d, 32'h441036c0},
  {32'h44427273, 32'h4263fdb6, 32'hc33260e1},
  {32'h43bf3e1e, 32'h434457c5, 32'h43824029},
  {32'h44cc6c74, 32'hc36a33cc, 32'hc184a280},
  {32'hc49e0c3b, 32'h43b07c97, 32'hc1245771},
  {32'h450be245, 32'hc3fcae65, 32'hc24b778b},
  {32'hc41285d6, 32'hc317ac9e, 32'h431ce428},
  {32'h44df7b26, 32'h43f112ca, 32'hc333fde4},
  {32'h437ae958, 32'h4115fc7c, 32'h42dc128d},
  {32'h44554748, 32'hc195162d, 32'hc0ae9842},
  {32'hc4a8d208, 32'h43b919a3, 32'h4365c667},
  {32'h437ec7a8, 32'hc3a9e55e, 32'h438c0364},
  {32'h400eef4c, 32'hc14893f5, 32'hc3408f08},
  {32'h444751a4, 32'hc2a4658e, 32'h436de63b},
  {32'hc3d8877c, 32'h438975ad, 32'hc2f1c803},
  {32'h43919f90, 32'hc2cd856c, 32'h42e5d40a},
  {32'hc516ab8b, 32'hc32edb6d, 32'hc35aaaf7},
  {32'h4452aaac, 32'h44601efe, 32'h435ae302},
  {32'hc51946ec, 32'h432b6849, 32'h431901b6},
  {32'h44bdf534, 32'h42788c5b, 32'hc28e8ba7},
  {32'h437cda61, 32'h42b6f303, 32'h436f1315},
  {32'h44dca765, 32'h438ec70d, 32'hc41a1bba},
  {32'hc4cb07f3, 32'h43850e20, 32'h436c1dbc},
  {32'h446e3c8c, 32'hc32b76e6, 32'h43194b8f},
  {32'hc4fabe16, 32'h4398c994, 32'hc22327ef},
  {32'h4517d8d9, 32'hc367cf42, 32'hc3214a96},
  {32'hc40d2d50, 32'hc3927e2f, 32'h4382e083},
  {32'h44116d05, 32'h43bf780a, 32'h428f56ba},
  {32'hc4926595, 32'hc2698a60, 32'hc08a8772},
  {32'h44350099, 32'hc34a0fd7, 32'h4314fdad},
  {32'hc425efd8, 32'h41c628f0, 32'hc2e649e8},
  {32'h44f6cba8, 32'h43e624a8, 32'hc1410557},
  {32'hc4f27f16, 32'h42af6b5e, 32'hc1cb1f49},
  {32'h4484db0c, 32'h431af5f7, 32'h428e48b6},
  {32'hc4fe89e4, 32'hc37f8386, 32'h42ab385c},
  {32'h4396ca60, 32'h42c77de1, 32'h42dc879d},
  {32'hc4d3d1cd, 32'hc20d8a85, 32'hc3ec2210},
  {32'h45086895, 32'hc2fe93b1, 32'hc30de83d},
  {32'hc50e3f32, 32'h430c1065, 32'h434b99af},
  {32'h446d1fa0, 32'hc40a6161, 32'h4325d2f9},
  {32'hc4637cd6, 32'hc0a23279, 32'h430ae3db},
  {32'h435036e0, 32'h430781f3, 32'hc3c29a6a},
  {32'hc497cba0, 32'hc39b9928, 32'h43bb6459},
  {32'h44c7a3cc, 32'hc25a8e07, 32'h419e1bf2},
  {32'hc4d36b0a, 32'h439b5a88, 32'h4302ac8e},
  {32'h42bfbebc, 32'hc3f08992, 32'hc2f36a64},
  {32'hc4a66366, 32'hc23d00d6, 32'hc28c9233},
  {32'h44b5d0b5, 32'hc391e305, 32'hc344fc6b},
  {32'hc43775e0, 32'hc300f805, 32'hc31a66f9},
  {32'h44995ea6, 32'hc32bff8e, 32'hc2d6c5b5},
  {32'hc5168216, 32'h4279c1a0, 32'hc1eec4bd},
  {32'hc1923240, 32'h43534f9a, 32'hc2cd0f16},
  {32'hc4a8a2ca, 32'hc213925f, 32'h415ce346},
  {32'h44fe4c61, 32'h41431b74, 32'hc3dbf899},
  {32'hc50c24f1, 32'hc385ec2b, 32'h43466e91},
  {32'h44bc20c8, 32'h4342b3ee, 32'hc37f8cb8},
  {32'hc4965f8e, 32'hc3e78870, 32'hc2223e0f},
  {32'h44d170fc, 32'hc1c552a1, 32'hc305d088},
  {32'hc40b44d0, 32'hc23f871e, 32'h430a3094},
  {32'h44c867da, 32'h41262b9f, 32'hc3bf9829},
  {32'hc4bfd4d8, 32'h41c3c965, 32'hc21beac6},
  {32'h4484b04d, 32'hc3b5d9b9, 32'hc35e4d46},
  {32'hc4ab9344, 32'hc2ab9b4b, 32'hc3a9806f},
  {32'h44bd997e, 32'h43678eb1, 32'hc3a3df4b},
  {32'hc37707b0, 32'hc2c17372, 32'hc2a08d23},
  {32'h43b7ad2a, 32'hc3183d06, 32'h42ec085e},
  {32'hc3f09e40, 32'hc1f01a97, 32'h42d3e074},
  {32'h44f85884, 32'hc240c724, 32'hbf06c903},
  {32'hc484cf28, 32'h43812f25, 32'hc3763bf5},
  {32'h4448c25a, 32'h42c62966, 32'hc2c7468a},
  {32'hc48af889, 32'h417480fc, 32'h42c0984b},
  {32'h44ff7b4e, 32'hc2af62a4, 32'hc2c2037e},
  {32'hc5074a77, 32'hc3293bbc, 32'hc1c6e71d},
  {32'h4390c56a, 32'h42b9dbe0, 32'h41861a84},
  {32'hc4a18e2d, 32'hc3522415, 32'hc36cad8f},
  {32'h44cfa4fc, 32'hc3aa70d0, 32'hc3b66902},
  {32'hc4cf461d, 32'hc414d0df, 32'h428c3cc6},
  {32'h43ae4fe0, 32'h417279fb, 32'h4316193a},
  {32'hc4137318, 32'hc394606e, 32'h43099de9},
  {32'h44db254a, 32'h439e2323, 32'h4367be18},
  {32'h42173a7d, 32'h42aa64b3, 32'h42ea168c},
  {32'h4512ac24, 32'h410eb9a0, 32'h4330bc95},
  {32'hc4f06de9, 32'hbd89f718, 32'hc1e64bd9},
  {32'h44d2961c, 32'hc2c15087, 32'hc250fc38},
  {32'hc4fa6da7, 32'h4369d9c2, 32'hc36d0564},
  {32'h431e98e7, 32'hc2acbcc9, 32'hc32d7c10},
  {32'hc4c6491f, 32'h43528b7e, 32'h43566b93},
  {32'h450b6abd, 32'hc34b0182, 32'hc2ef99ea},
  {32'hc3901c20, 32'h433c1be3, 32'hc199cc55},
  {32'h446fe8d2, 32'h43dfe677, 32'hc19154d1},
  {32'hc3d415cc, 32'hbf8e4628, 32'hc186dcf2},
  {32'h4491c1eb, 32'h430c59ac, 32'h43e0d37e},
  {32'hc39b5874, 32'h42ef6238, 32'h427ad26b},
  {32'h4461349e, 32'h43485070, 32'h410b5ada},
  {32'hc2c29620, 32'h42fe933d, 32'hc2d7872c},
  {32'h43b4511d, 32'h43654a60, 32'hc3c78c06},
  {32'hc40992e8, 32'hc30f1db1, 32'h41c6d184},
  {32'h43921024, 32'hc33ad08c, 32'hc4058a69},
  {32'hc39253b8, 32'h426e15ec, 32'hc3c5be3c},
  {32'h45008ba6, 32'hc2845fe4, 32'hc0ddc261},
  {32'hc3d38be4, 32'hc35be41b, 32'hc2594544},
  {32'h448a6a9a, 32'hc3ec4a53, 32'hc2049814},
  {32'hc4d6dc5e, 32'h425e9b1b, 32'h435f8509},
  {32'h44b79ab6, 32'hc1cb0b47, 32'hc35897b3},
  {32'hc4575424, 32'h436394fc, 32'h431cdb3c},
  {32'h43fc458c, 32'h43249172, 32'h43a139b4},
  {32'h441e98d0, 32'hc219e692, 32'h42b54315},
  {32'h44d7b9c7, 32'h42878947, 32'h422e5c21},
  {32'hc4b5e716, 32'h42f22a24, 32'hc284c8b6},
  {32'h4221bf40, 32'h430ad430, 32'hc3491b22},
  {32'hc4879ae1, 32'h42a41baa, 32'h43beae75},
  {32'h44db3ffb, 32'hc362a7a8, 32'hc1e162d4},
  {32'hc34aaf0b, 32'hc2858eab, 32'hc2de6aee},
  {32'h449d8746, 32'hc2dd6514, 32'h42ef48b2},
  {32'hc4585896, 32'h4305dbd6, 32'hc3f74150},
  {32'h4488ad80, 32'hc1dfdc29, 32'h4342834c},
  {32'hc4f02f42, 32'h4363e098, 32'h43762180},
  {32'h4481088c, 32'h422202b7, 32'hc413bc83},
  {32'hc4fc79f5, 32'hc32e5d10, 32'hc20e030e},
  {32'h4503ebf2, 32'hc1e552c5, 32'h43cb3595},
  {32'h41696d00, 32'hc3c4fdb7, 32'h430948ee},
  {32'h446db962, 32'hc3387c15, 32'h43303e8e},
  {32'hc4e2a518, 32'hc2588836, 32'hc3cfc76a},
  {32'h4434d980, 32'h436de156, 32'h43f8cee5},
  {32'hc3da4afa, 32'hc2c21995, 32'hc271b135},
  {32'h4334aae0, 32'h421024ec, 32'h4284b848},
  {32'hc334f190, 32'hc359756e, 32'h43369da8},
  {32'h44578710, 32'hc229547b, 32'hc2da1787},
  {32'hc346f720, 32'hc298ad8e, 32'h421b12db},
  {32'h44f21f3e, 32'h42c6206e, 32'h4330a87a},
  {32'hc3eb8f86, 32'h42933865, 32'h4141ee50},
  {32'h43efb5b4, 32'h414d6b18, 32'h4335f307},
  {32'hc376fe28, 32'hc1110b31, 32'hc2c6bc9c},
  {32'h43f5f5f0, 32'h436c507e, 32'hc3b46750},
  {32'hc507ac5a, 32'hc28a0903, 32'h426434f9},
  {32'h44ef20f6, 32'h42d85fee, 32'h4370f6d6},
  {32'hc50a6f28, 32'h43689821, 32'hc3b80d41},
  {32'h44eee955, 32'h43596603, 32'h42ceded2},
  {32'hc3a7c3b8, 32'h43af3016, 32'h4210aee7},
  {32'h4489fd34, 32'h42de4017, 32'hc32128bf},
  {32'hc3d9eeb0, 32'hc2c7c8c2, 32'hc416be0d},
  {32'h43474b91, 32'hc3658dc0, 32'hc2893495},
  {32'hc3600795, 32'hc3898acc, 32'h430f32dd},
  {32'h45183c3c, 32'hc384cf70, 32'hc3a672e8},
  {32'hc49f5e7b, 32'hc36e3b00, 32'h42efdc1e},
  {32'h44fabf6a, 32'hc2ccfa4d, 32'h42edcbe3},
  {32'hc465f994, 32'hc3238f36, 32'hc36375a5},
  {32'hc3a89f2c, 32'h43923beb, 32'h4364aefc},
  {32'h43d67a64, 32'h41c7018b, 32'hc299f8b5},
  {32'h44072440, 32'hc21c956a, 32'h439480fb},
  {32'hc4d83855, 32'hc39da246, 32'hc1bd4b13},
  {32'h44215156, 32'hc3920aed, 32'h418f3a28},
  {32'hc50634f7, 32'hc2fa26aa, 32'hc202b153},
  {32'h444d6ae2, 32'hc2a7c17d, 32'hc167ca1a},
  {32'hc39a50cc, 32'h42d861ca, 32'hc2d32274},
  {32'h438ab787, 32'hc3b302ba, 32'hc3c73ad5},
  {32'hc415be84, 32'h43085d2a, 32'h43858a86},
  {32'h44c72942, 32'hc3e09e3f, 32'hc1fec8a5},
  {32'hc4bc227e, 32'hc384e161, 32'hc3845870},
  {32'h43e244f4, 32'h431066b3, 32'h42c61d3f},
  {32'hc430af68, 32'hc3d27cb9, 32'hc3279c65},
  {32'h44774ada, 32'hc397f597, 32'hc31736dd},
  {32'hc32deec8, 32'hc1947320, 32'hc4000044},
  {32'h43ccf12c, 32'h430f1f29, 32'h43163d28},
  {32'hc4af7f60, 32'hc31329f2, 32'hc3ff56e1},
  {32'h440da282, 32'hc2f1c99d, 32'h431cf770},
  {32'hc4f2023e, 32'h430ce951, 32'h42dd73e5},
  {32'h43c80517, 32'h434ed055, 32'hc2dce86d},
  {32'hc511e684, 32'hc3a39d71, 32'h432a0302},
  {32'h444ea97c, 32'h428eec28, 32'h43171645},
  {32'h42ebf5dc, 32'hc3b31f7b, 32'h439d89e1},
  {32'h44c4c3c1, 32'hc322681e, 32'h430c5897},
  {32'hc506f228, 32'h412683f6, 32'h438f5097},
  {32'h446d9652, 32'hc35c542b, 32'hc2b3d325},
  {32'hc49962ea, 32'h41658cf7, 32'hc3b6facd},
  {32'h449bd3f6, 32'h434785c3, 32'h43450e20},
  {32'hc3d33557, 32'hc1955737, 32'hc240f368},
  {32'h44863cd2, 32'h430e70c2, 32'h42d79541},
  {32'hc3d77896, 32'hc1d8b716, 32'h42aa2f0f},
  {32'h44439dd2, 32'h4302008b, 32'hc34994a5},
  {32'hc4b5c4b0, 32'hc397c7a0, 32'hc343994c},
  {32'h450aa206, 32'hc34dc876, 32'hc10edb74},
  {32'hc4426ace, 32'h43283cfd, 32'h430a8f94},
  {32'h43658026, 32'hc3065aa5, 32'hc304e3f3},
  {32'hc41bd7d4, 32'hc1a7a1b8, 32'hc3647f88},
  {32'h44f13f69, 32'h4368c9ae, 32'hc2fd1c2e},
  {32'hc2e3f860, 32'hc347a0e1, 32'hc3eb5307},
  {32'h451989bf, 32'h4307789c, 32'hc2dfa7c6},
  {32'hc2634092, 32'h43e12223, 32'hc388481d},
  {32'h44c3e2b1, 32'hc3093de0, 32'hc1d5b653},
  {32'hc35713d0, 32'h43f27b18, 32'hc3d70e58},
  {32'h44e72c0a, 32'hc30454b8, 32'hc3019867},
  {32'hc4d35174, 32'hc387b4f6, 32'h42619db6},
  {32'h447c62dc, 32'h426a770a, 32'h41a6bc66},
  {32'hc4233bee, 32'hc3b6c77a, 32'h4397149f},
  {32'h4501f679, 32'h43e0f3dc, 32'h42ce7f13},
  {32'hc3a11a88, 32'hc2383791, 32'h42727751},
  {32'h44a7a114, 32'h4388ca10, 32'h3fe2ffa0},
  {32'hc413f1fe, 32'hc30a6bfc, 32'hc2a4df54},
  {32'h44a95f41, 32'hc279b64a, 32'hc20db096},
  {32'hc5064603, 32'h431ef7d0, 32'hc196bcdf},
  {32'h44ff82b8, 32'h435b2ae0, 32'h42c86ce6},
  {32'hc513cf2a, 32'h4407817f, 32'h42361384},
  {32'h43e59f12, 32'hc3b030bf, 32'hc24182bc},
  {32'hc4b5a27a, 32'hc31059e8, 32'hc19ad194},
  {32'h44b80ab4, 32'hc2d9df6b, 32'h4335c4a6},
  {32'hc4b3aa2a, 32'h418adc84, 32'h4339ed8d},
  {32'h44aadffa, 32'hc3028a63, 32'h42c6970d},
  {32'hc453ca28, 32'h3e8a39c8, 32'hc385b31c},
  {32'h45078161, 32'h40b71d08, 32'hc1cc441d},
  {32'hc4e0e6ac, 32'hc19d763c, 32'h4381cc2b},
  {32'h44e432bb, 32'h42183f39, 32'h41312f97},
  {32'hc2988ec0, 32'h43985fa2, 32'hc383e834},
  {32'h440c6e57, 32'h4395d15d, 32'h437d51ff},
  {32'hc483c21b, 32'hc3145953, 32'h435960aa},
  {32'h4465469a, 32'h4365a6ae, 32'hc2aa8ec6},
  {32'hc48da5b4, 32'hc3429815, 32'hc3893579},
  {32'h44dbbbee, 32'hc357498b, 32'h4306c1c2},
  {32'hc4ed0fd8, 32'hc3ccf541, 32'h42f36926},
  {32'h4268d5a0, 32'hc328190a, 32'h43dabcb9},
  {32'hc5026393, 32'hc2ee35d0, 32'hc2b6835a},
  {32'h44f9ef96, 32'h42b00e9c, 32'hc31490c7},
  {32'hc4e8fa3e, 32'hc38ad86c, 32'h4335e28b},
  {32'h44c8c23c, 32'hc18aea81, 32'hc2613ddc},
  {32'hc470ba64, 32'h438daa3a, 32'hc34fa050},
  {32'h442ba4a6, 32'hc315b5ec, 32'hc2f6ca93},
  {32'hc47d1dcc, 32'h43a5421d, 32'hc345cb25},
  {32'h449495a0, 32'hc3969137, 32'h432494dc},
  {32'hc3b30be0, 32'hc391aa80, 32'hc4051af5},
  {32'h449ed069, 32'hc357ae37, 32'h438ee7df},
  {32'hc4bbef22, 32'h422ee0f6, 32'hc231b65b},
  {32'h44cc17c8, 32'h42e06a00, 32'hc1b0accd},
  {32'hc46cda70, 32'h412f52f3, 32'h412ec353},
  {32'h44a36562, 32'hc326660c, 32'h415e0842},
  {32'hc23c15a0, 32'hc307c225, 32'h43b17538},
  {32'h442b9769, 32'hc3423e40, 32'h4397c8dd},
  {32'hc45fb63a, 32'hc344ed54, 32'hc3aa0736},
  {32'h450b3052, 32'h42f658e9, 32'h439ff798},
  {32'hc3ea3180, 32'h438b4379, 32'hc288c517},
  {32'h4496cbeb, 32'h43033787, 32'h42f7a23f},
  {32'hc40241c6, 32'hc38a1bb0, 32'h4299f06f},
  {32'h44ff3b3f, 32'h43863973, 32'hc345c755},
  {32'hc51d0854, 32'h43427403, 32'hc3df2da4},
  {32'h451da98d, 32'hc3ca526f, 32'hc2cad4f4},
  {32'hc482e812, 32'hc3426ef1, 32'h42b632cf},
  {32'h423a1f00, 32'h4371e88c, 32'h4350bf2f},
  {32'hc498f76e, 32'hc0d03c10, 32'hc37174c4},
  {32'h44ec55f5, 32'hc34ec0f8, 32'hc304a8c0},
  {32'hc47c7e9f, 32'h424c4667, 32'h42758c18},
  {32'h44b184a0, 32'hc20a2b5a, 32'h42a4bab9},
  {32'hc4a7b41e, 32'hc36947c6, 32'hc2821b6e},
  {32'h450d8214, 32'hc32a360b, 32'h422d2682},
  {32'hc504fa00, 32'hc39f4d51, 32'hc3197a59},
  {32'h44ea0614, 32'hc3cbd13f, 32'h4334df9a},
  {32'hc4a6dcbf, 32'h4133a665, 32'hc219feb9},
  {32'h443ec4c0, 32'h41b7e67e, 32'h43ab10b8},
  {32'hc506533e, 32'h41c54b46, 32'h433bbdcd},
  {32'h449921bc, 32'hc3557521, 32'hc3987d00},
  {32'hc51140f7, 32'hc31444b4, 32'hc311e1e2},
  {32'h44107bee, 32'h43b51c50, 32'h43d4e3a8},
  {32'hc484fb7c, 32'h4364719e, 32'h4156b535},
  {32'h4439a4fa, 32'hc1b99e50, 32'h3fdaa210},
  {32'h43a0af98, 32'h438f11a7, 32'hc32feec1},
  {32'h44edd654, 32'hc3892317, 32'hc28a01c9},
  {32'hc3d8899b, 32'h42882e59, 32'h43364579},
  {32'h44a61cef, 32'hc39bbdf0, 32'hc37617f5},
  {32'h436349fe, 32'h4396a587, 32'hc30db112},
  {32'h44d443df, 32'h43a27820, 32'hc27a693d},
  {32'hc3e71b20, 32'h4293c974, 32'h43bbbda1},
  {32'h450ad188, 32'h432b0f45, 32'h42d077ca},
  {32'hc48d6872, 32'h42d8a988, 32'hc33ad4de},
  {32'h4514f16f, 32'h41df8bc0, 32'hc1f42b4d},
  {32'hc4442d0e, 32'h42875f33, 32'hc31b5196},
  {32'h4467d135, 32'h41c97902, 32'hc3022a42},
  {32'hc525471e, 32'hc3804dad, 32'h43488823},
  {32'h450d2b5c, 32'h42cd7d88, 32'hc19dc7a5},
  {32'hc50e8f07, 32'hc4066148, 32'hc3957ccc},
  {32'h4385afcc, 32'hc1be0abe, 32'h42ced984},
  {32'hc4c2a631, 32'hc29db43c, 32'hc38e439c},
  {32'h450f93ec, 32'h43d3fed4, 32'hc2fb4a98},
  {32'hc4ba0f63, 32'hc2e8369f, 32'h443b34bd},
  {32'h44bf04d0, 32'hc38bc83c, 32'hc36fa6a0},
  {32'hc4e98ac4, 32'h43a6647f, 32'hc40dfb8e},
  {32'h44f50965, 32'h422b9090, 32'hc297cf85},
  {32'hc49c9a5a, 32'h4331abc4, 32'hc2a28d67},
  {32'h44ff6455, 32'h4331e365, 32'hc2b4cc56},
  {32'hc4edc21c, 32'h42b1102f, 32'hc2ed26d4},
  {32'h448edeee, 32'h431f8994, 32'hc2d23385},
  {32'hc512aacf, 32'hc20b08ce, 32'h4305ed3e},
  {32'h448fd259, 32'hc388be1a, 32'h4313fd37},
  {32'hc42707b8, 32'hc2f27552, 32'h4358472e},
  {32'h44f45754, 32'hc3ea56c0, 32'hc30743e3},
  {32'hc4d07e30, 32'h43ef5156, 32'h436393f2},
  {32'h447194d0, 32'hc32b8088, 32'h42bea3e8},
  {32'hc41cfab2, 32'hc2bd68e5, 32'hc3cd0283},
  {32'h43e1302f, 32'h41a4cfda, 32'hc2b896b2},
  {32'hc411687f, 32'h42dd1f73, 32'hc2c54642},
  {32'h45081b1a, 32'h43a142de, 32'hc387dfe8},
  {32'hc43e80d4, 32'h43644144, 32'h42b041a3},
  {32'h44259ea4, 32'h42fd0841, 32'h41caab14},
  {32'hc4db709e, 32'hc32be5c4, 32'h4313e552},
  {32'h446df094, 32'hc38b4a76, 32'hc35ae40b},
  {32'hc5030a18, 32'hc3931deb, 32'hc31c8345},
  {32'h43f43a36, 32'hc2c6ac10, 32'hc351df16},
  {32'hc4f5930b, 32'h43642d12, 32'h433886f5},
  {32'h43bbacd7, 32'h42961188, 32'hc39445e6},
  {32'hc4ae02f9, 32'hc31dc5ee, 32'h43fe0997},
  {32'h444bcfcc, 32'h43019ed5, 32'hc3958342},
  {32'hc49f77dc, 32'hc2852194, 32'h434b1d0d},
  {32'h45052622, 32'h43a247aa, 32'h4276bf10},
  {32'hc418ec8d, 32'hc328fc2a, 32'h4310d208},
  {32'h44ce7d38, 32'h40b9500f, 32'hc385a072},
  {32'hc4b5023f, 32'h4320e7ef, 32'h42177bc9},
  {32'h43534cb0, 32'h428260b4, 32'h427eb2f0},
  {32'hc3e452c4, 32'h4380c9db, 32'hc22231cf},
  {32'h4507fa76, 32'hc23c161a, 32'h431c1893},
  {32'hc46c5a2d, 32'h426b8162, 32'hc2d5a091},
  {32'h438294f4, 32'h40b910bc, 32'h43e9db7d},
  {32'hc496dac4, 32'hc0629ea3, 32'h4298ef89},
  {32'h44c0fedb, 32'h42a30e4a, 32'hc3497613},
  {32'hc4bf2c31, 32'h43a3e36d, 32'hc2ff4359},
  {32'h42a952be, 32'hc3a89a85, 32'hc300fd14},
  {32'h4391256c, 32'h43620637, 32'h42e568b8},
  {32'h44c2e5cf, 32'hc2e9eb06, 32'hc32787b6},
  {32'hc4a639dc, 32'h4391df32, 32'hc2d23bc9},
  {32'h43f06534, 32'h42f15c8b, 32'hc05f2047},
  {32'hc5077c20, 32'hc345f5e5, 32'hc2f7ee9c},
  {32'h44636651, 32'h4385bc01, 32'h4223c664},
  {32'hc4bc4e1d, 32'hc38f607b, 32'h43a71a3d},
  {32'h4500a410, 32'hc31177ea, 32'h43208f64},
  {32'hc4552b7e, 32'hc37a67bc, 32'h43ff62df},
  {32'h44dec23c, 32'h42f6049c, 32'h4336f095},
  {32'hc492da23, 32'hc2c6bd23, 32'h4255af3d},
  {32'h43d60be8, 32'hc2665abf, 32'h41a7b09e},
  {32'hc411ad82, 32'h4397e1ad, 32'hc379e080},
  {32'h44ab58b0, 32'hc2ed0cc0, 32'h43507ff0},
  {32'hc2dfe7e0, 32'h4392edf7, 32'h427a6451},
  {32'h44107542, 32'hc293f7f0, 32'hc383e43f},
  {32'h43fbc401, 32'h419469c5, 32'hc3985305},
  {32'hc3ca68b8, 32'hc3c548fe, 32'h438f96f1},
  {32'h4401d7c0, 32'h431ba7b1, 32'h42833ef8},
  {32'hc4fe7fc8, 32'hc2887c97, 32'hc33800bd},
  {32'h44bbaf3e, 32'hc38d91db, 32'h421d98ab},
  {32'hc3b7b6aa, 32'h42845b5a, 32'h431df478},
  {32'h448f7ce9, 32'hc32552da, 32'hc40ef11f},
  {32'hc49ca69b, 32'hc2f76d46, 32'hc2bec71c},
  {32'h450c54f9, 32'hc347c86e, 32'hc2d17540},
  {32'hc49150bd, 32'hc2777f9e, 32'hc3ea1591},
  {32'h43d59888, 32'hc33fc294, 32'hc396757d},
  {32'hc4bb3214, 32'h437a99ed, 32'h43fafa8c},
  {32'h44e8b565, 32'hc2d8ec47, 32'hc360fd66},
  {32'hc3de0960, 32'h433c2688, 32'h42fab2ec},
  {32'h4448e976, 32'h4344edf3, 32'hc395e6e1},
  {32'hc379b3f8, 32'h43c4ddc0, 32'h4323aa6a},
  {32'h44b91d38, 32'hc33f702a, 32'hc1882ca0},
  {32'hc3e98345, 32'h42582027, 32'hc196c5eb},
  {32'h45339eb6, 32'h41f925a7, 32'hc19d9929},
  {32'hc48a29ee, 32'hc2527df2, 32'h4394e9de},
  {32'h45075622, 32'h42de4d4c, 32'h431df6c3},
  {32'hc4f68c58, 32'hc325401c, 32'hc397f0f9},
  {32'h4511c03c, 32'h428fbf86, 32'hc39fa848},
  {32'h43699640, 32'h433c41a3, 32'hc36c877f},
  {32'h448c47e6, 32'h43481951, 32'hc3a6fdd4},
  {32'hc467cf53, 32'h414ee8f2, 32'h43c331fe},
  {32'h44e47795, 32'hc356415c, 32'h4348ac41},
  {32'hc3d58d42, 32'hc300bb16, 32'hc2950c34},
  {32'h44e8bb98, 32'h43df31be, 32'hc3817012},
  {32'hc4a28e98, 32'h4357b100, 32'hc2018edd},
  {32'h442e63e0, 32'h43671d48, 32'h418e09eb},
  {32'hc48563c4, 32'h42149ad8, 32'hc2533e53},
  {32'h436d22f0, 32'h436dd687, 32'hc2e30325},
  {32'hc4bf49e9, 32'hc1cd85de, 32'hc1e7ca9d},
  {32'h44a1b0eb, 32'h4319af4c, 32'hc33149d3},
  {32'hc2aa8c40, 32'hc302479e, 32'hc231c60f},
  {32'hc3ca6840, 32'h406123c2, 32'hc3c3108c},
  {32'hc4f8db6e, 32'h43b77331, 32'hc318d291},
  {32'h45239ce5, 32'hc2edb62b, 32'h43b2c48a},
  {32'hc4cdbdf9, 32'h42a8f9f1, 32'h434ee1d1},
  {32'h4508cba0, 32'h43d2b9a3, 32'h44090df9},
  {32'hc4459e14, 32'h4314fa08, 32'h4254eb41},
  {32'h44f191d6, 32'hc2dd949c, 32'hc30dd5e5},
  {32'hc42db9f3, 32'hc42c6c59, 32'h429a8083},
  {32'h44874a1f, 32'hc30b0137, 32'h4391e31e},
  {32'hc5039b0c, 32'h430e33ef, 32'hc2aebabf},
  {32'h429b1c68, 32'h431c7228, 32'hc29b1063},
  {32'hc4dce8e9, 32'hc1fb1d13, 32'h42dfd70c},
  {32'h4496053e, 32'hc29c4b4f, 32'hc2a343d5},
  {32'hc4f59fff, 32'hc294da67, 32'h423515b6},
  {32'h439ede92, 32'h4196601d, 32'h425a7c3f},
  {32'hc33b3718, 32'hc31ed9bb, 32'h432c5d6e},
  {32'h449bba16, 32'hc2759d73, 32'hc3e2933b},
  {32'hc440c234, 32'h4176babf, 32'h42dbbbf0},
  {32'h446bcc50, 32'hc2904e35, 32'hc2d35dae},
  {32'hc48ec198, 32'h4342f6a2, 32'h420c0314},
  {32'h43afec9e, 32'h43b75bc5, 32'h4395f85e},
  {32'hc4cc703e, 32'hc2a4b8d5, 32'hc329ebf6},
  {32'h4480b52e, 32'h434b3c1c, 32'hc2920d8e},
  {32'hc34e6420, 32'h417c9364, 32'hc33f445b},
  {32'h443723e9, 32'h4391850b, 32'h430fe462},
  {32'hc4d2ffb2, 32'hc2a0301c, 32'h4372a196},
  {32'h45122818, 32'h42ae5dd2, 32'hc1d8311a},
  {32'hc3b69400, 32'h41e06ba3, 32'h42738d1f},
  {32'h436544b4, 32'h42ac1bb9, 32'h430d9bf0},
  {32'hc47be3c2, 32'h43cff1e8, 32'h436e1302},
  {32'h4507fa58, 32'hc39e8953, 32'hc34c6d9e},
  {32'hc4a19b7f, 32'h42b00b3f, 32'hc2a3288b},
  {32'h443f7948, 32'h43548c70, 32'h4340bbef},
  {32'hc4a9cee2, 32'hc3a90ec0, 32'h42e86758},
  {32'h44764e61, 32'h400bb750, 32'h4319d529},
  {32'hc413d7ae, 32'hc39c1531, 32'hc30d2530},
  {32'h43c69182, 32'hc30b99e2, 32'hc2626557},
  {32'hc415d9b8, 32'h3f22e978, 32'h432724d9},
  {32'h44c57f79, 32'hc2df7316, 32'h43c44de4},
  {32'hc507c00c, 32'hc3495153, 32'hc2a0b8cc},
  {32'h450857ca, 32'hc36300a0, 32'hc2771178},
  {32'hc45026ed, 32'hc2adbc0b, 32'h411123f1},
  {32'h44f7e3cb, 32'h435a8e7d, 32'h43975c21},
  {32'hc400958c, 32'h426f2804, 32'hc3536b80},
  {32'h450ebd44, 32'hc36b79c4, 32'h43a98b0a},
  {32'hc512454e, 32'h3fc34870, 32'hc2a9c323},
  {32'h43c8d9b7, 32'h42810e02, 32'hc1e2d7f2},
  {32'hc4bef19d, 32'hc34ce122, 32'hc37755fe},
  {32'h4441a1b0, 32'h43df9fde, 32'hc31ed002},
  {32'hc4bdbba6, 32'hc33f383d, 32'h4293d004},
  {32'h43ec8875, 32'h4205afd7, 32'hc289383e},
  {32'hc387f27c, 32'h436ffa9e, 32'hc35f5bbf},
  {32'h45078382, 32'hc3ac34d7, 32'h434f9184},
  {32'hc4310e50, 32'hc2d7bdcb, 32'h42ef3e9d},
  {32'h450c4857, 32'h438731e8, 32'h422d4c24},
  {32'hc4c1443b, 32'h42ed1334, 32'hc1fecec7},
  {32'h441e4c1b, 32'h43419f5a, 32'hbfe67fec},
  {32'hc5001f09, 32'h43d4dccd, 32'hc2e4858d},
  {32'h440721b5, 32'hc3f73533, 32'hc245fa8d},
  {32'hc43e8c83, 32'h43766d1e, 32'hc30fd9f6},
  {32'h43dd7b3a, 32'h42bb5889, 32'h43b51941},
  {32'hc4d02952, 32'hc37deb01, 32'hc2a4244f},
  {32'h44aae1be, 32'hc41d9278, 32'h41ba1aea},
  {32'hc4cbde54, 32'h429325ac, 32'h43458159},
  {32'h439439ec, 32'h43a07e4f, 32'hc3085c7c},
  {32'hc2f0b080, 32'hc13353fa, 32'h40e28b08},
  {32'h44c8fe5b, 32'h42f4b57b, 32'h43835ea5},
  {32'hc4d4b146, 32'hc328fdfc, 32'h42d147c3},
  {32'h44f8846a, 32'hc2271d53, 32'h42772dd3},
  {32'hc4ebbe8e, 32'hc317a530, 32'hc300df12},
  {32'h451cf341, 32'h41703c78, 32'h42c52ff5},
  {32'hc4ca1f07, 32'hc39ea3e6, 32'h42918297},
  {32'h439d96fa, 32'h4317db2f, 32'hc369347a},
  {32'hc46626d8, 32'hc2817ab6, 32'h41073996},
  {32'h43106218, 32'h4390598b, 32'hc268e700},
  {32'hc5097827, 32'hc2716e32, 32'h43f58d82},
  {32'h43435a30, 32'h4418d2e7, 32'h432cef65},
  {32'hc4f2920b, 32'h4374c16a, 32'hc22a781c},
  {32'h4416e076, 32'hc2fb87ad, 32'h43888200},
  {32'hc4cc028a, 32'hc36eb2a4, 32'h4194ed52},
  {32'h44e1431a, 32'hc25c767c, 32'h438a4f41},
  {32'hc4638969, 32'h41705572, 32'h436c1f3f},
  {32'h43bd8144, 32'h4301dda5, 32'h42f42d10},
  {32'hc4a2873a, 32'h43a4a35b, 32'h429a38da},
  {32'h438018a6, 32'h4391e283, 32'hc0d0a488},
  {32'hc33a18c9, 32'hc1c43595, 32'hc19ac90a},
  {32'h44393084, 32'h431185a8, 32'h43b9b9fa},
  {32'hc4cfc48e, 32'hc3114b0b, 32'h439d553f},
  {32'h44a10c18, 32'h42cb713a, 32'hc3a76cb6},
  {32'hc4234bcc, 32'hc3e1e8d2, 32'hc402cc88},
  {32'h44407517, 32'hc29890ea, 32'hc39d9013},
  {32'hc4468923, 32'h43c2a1f4, 32'h42462d70},
  {32'h44d4dfd2, 32'hc287db54, 32'h436654ac},
  {32'hc4c0bfc4, 32'h438802dd, 32'hc315ee95},
  {32'h436949b0, 32'hc3a4ebb6, 32'h439c80ce},
  {32'hc442a1ea, 32'h4286f2b3, 32'h43d4753b},
  {32'h44fa8c25, 32'hc0d1b1c2, 32'h42fcbad1},
  {32'hc4a6ea6e, 32'hc2ded2cc, 32'h4397faa7},
  {32'h44c4fdbe, 32'h43ff84ae, 32'h43850f0a},
  {32'hc3ac6131, 32'hc29ca294, 32'hc329c7f3},
  {32'h44d6a1e3, 32'hc3312d0b, 32'h429353ab},
  {32'hc512871d, 32'hc2a12c7c, 32'hc15afe9b},
  {32'h441d18bc, 32'h432eaf8e, 32'h42b3ed82},
  {32'hc4cdc0bd, 32'h43de257c, 32'h4305953a},
  {32'h4513048a, 32'hc218b6de, 32'hc30d23a4},
  {32'hc47904fa, 32'hc2af47a8, 32'hc2dd8a28},
  {32'h44ebd446, 32'h4118245f, 32'h41e471d9},
  {32'hc464ebc3, 32'hc305c7f5, 32'h4325eb57},
  {32'h4486f58d, 32'hc2911b1a, 32'h439c1fb5},
  {32'hc3d3e0da, 32'h42a15adb, 32'h4354d7e9},
  {32'h448fcd28, 32'hc2b84c3d, 32'h42af87e8},
  {32'hc38e82bb, 32'h43487a22, 32'h4183788c},
  {32'h44190f71, 32'hc19f7fa4, 32'h44017260},
  {32'hc42cd521, 32'hc1bb825f, 32'h4380bf85},
  {32'h44c4eff2, 32'hc215884f, 32'hc2f5b698},
  {32'hc45ad0b3, 32'h4307e13f, 32'hc2b015f1},
  {32'h44259922, 32'h4307aab1, 32'hc394c674},
  {32'hc4361833, 32'h4319c2e3, 32'hc1d5a3a4},
  {32'h4450ec04, 32'h42aed051, 32'h41906cd6},
  {32'hc5092abe, 32'h42e751d4, 32'h42a7e9f0},
  {32'h4492cd8f, 32'hc30365bf, 32'h419f39bf},
  {32'hc3655b39, 32'h43e49d2a, 32'h41f02de1},
  {32'h4482e2ea, 32'hc3a7ea8d, 32'hc2ef59db},
  {32'hc4bb96be, 32'h441a9578, 32'hc310d299},
  {32'h44d6f6bd, 32'hc32377dd, 32'h431b9442},
  {32'hc22b7120, 32'hc38f9060, 32'hc451b687},
  {32'h4451cf7e, 32'h429e8571, 32'h42e0b3bd},
  {32'hc33b0b00, 32'h4350abae, 32'hc3e3c5d2},
  {32'h43ada608, 32'h439d0194, 32'h4382935f},
  {32'hc4b281c1, 32'h43a190d3, 32'h4326e809},
  {32'h44352c79, 32'h429c6748, 32'hc2014934},
  {32'hc4f4758e, 32'h42c27cf8, 32'hc2b0562d},
  {32'h450e5d4a, 32'hc25f26d1, 32'hc3bd4966},
  {32'hc50a0c10, 32'hc32ec8b8, 32'h42cc4d1f},
  {32'h4425f155, 32'h436cbcd4, 32'h433c87f5},
  {32'hc3ed4766, 32'h42ecc176, 32'h43a5aef5},
  {32'h44688537, 32'h428b462d, 32'hc3eed98b},
  {32'hc478f88d, 32'hc3861d48, 32'hc18b47f3},
  {32'h43a1a8f2, 32'h43fb1c30, 32'hc32c4431},
  {32'hc48e6bf3, 32'h416ecd87, 32'hc3ed7be7},
  {32'h4502021c, 32'hc2b30658, 32'hc3a3022a},
  {32'hc482ffb4, 32'hc2d377ba, 32'hc3aed3f4},
  {32'h44f666b6, 32'h429001e8, 32'hc1ccd281},
  {32'hc468ece4, 32'h433de042, 32'hc28b7991},
  {32'h44c1420a, 32'hc1ee5e3e, 32'hc3b235ea},
  {32'hc4fe65dc, 32'hc3d5467c, 32'h42d14661},
  {32'h4503db8d, 32'h43ca99d3, 32'hc29fac8d},
  {32'hc47abefc, 32'hc2e5aa0f, 32'hc3d39a61},
  {32'h44f24785, 32'hc2bbeca9, 32'h425f2ce8},
  {32'hc50276b0, 32'h439c3cc6, 32'h43252340},
  {32'h450c46ea, 32'hc3c01f72, 32'hc31b37a3},
  {32'hc3773970, 32'h42c9d05d, 32'h42665789},
  {32'h451764f5, 32'h42c92bca, 32'hc0120ce0},
  {32'hc4b062cb, 32'h41bf5a66, 32'hc2fadc9c},
  {32'h449c6356, 32'h42acea44, 32'h440270d4},
  {32'hc418758e, 32'hc2887b29, 32'hc3da4e2d},
  {32'h44d8406e, 32'hc2789211, 32'h43a75012},
  {32'hc48126e3, 32'hc2ac7533, 32'h41fd9dda},
  {32'h449a743b, 32'hc2ebdea0, 32'hc34b7656},
  {32'hc49a1286, 32'hc3001eda, 32'h41757ba1},
  {32'h44a34863, 32'hc36cb55b, 32'hc3a62d7b},
  {32'hc4f61226, 32'hc31dd99f, 32'hc20add41},
  {32'h44a36984, 32'h4397f335, 32'hc3a3b149},
  {32'hc41de56a, 32'h43323a6b, 32'h43318243},
  {32'h445852b6, 32'hc3c86396, 32'h440758d9},
  {32'hc2e3b38d, 32'h42ae373c, 32'hc309bc62},
  {32'h45050b8e, 32'h42fb4642, 32'hc35dc892},
  {32'hc48427a0, 32'hc331e9de, 32'hc3ad8aba},
  {32'h44731c2c, 32'h41899c8a, 32'h42587343},
  {32'hc4d3231e, 32'h42c353f7, 32'h438fc06c},
  {32'h44f46800, 32'h43e17c2f, 32'h43402c31},
  {32'hc38a4f77, 32'hc379d81c, 32'h430e3556},
  {32'h450779ab, 32'h431adf27, 32'hc2bbca2f},
  {32'hc4e96402, 32'h42f7929d, 32'hc4159f97},
  {32'h4501e86d, 32'h43117496, 32'hc37f000d},
  {32'hc30ba1a6, 32'hc37782d2, 32'hc2b06847},
  {32'h447f58fb, 32'h436b0529, 32'h42a9b93a},
  {32'hc4f7025d, 32'h43b195ae, 32'h43d93149},
  {32'h44b33097, 32'h4352467b, 32'h4329b8db},
  {32'hc441c7e0, 32'h4250b38e, 32'hc3253b57},
  {32'h44f58941, 32'h41034892, 32'hc20aeba5},
  {32'hc500d3b8, 32'hc40ac937, 32'h40aa5e8e},
  {32'h44fd4c34, 32'h421f746c, 32'hc40b1530},
  {32'hc485405a, 32'hc2a964da, 32'hc2875a09},
  {32'h433b9fb0, 32'hc2d6916d, 32'hc31511f0},
  {32'hc48e6a56, 32'hc2b10a0d, 32'h427dfa7e},
  {32'h44b75c90, 32'hc22b6658, 32'h4217295d},
  {32'hc4cd320a, 32'hc37fba7a, 32'h41544806},
  {32'h439c35df, 32'hc37c57d3, 32'h43803477},
  {32'hc3a54088, 32'hc2b20200, 32'hc2cafcba},
  {32'h4514c2d1, 32'hc2966982, 32'h42e2fd11},
  {32'hc4d1d047, 32'h43224b20, 32'h42e532c4},
  {32'h45010a24, 32'h4332ecc5, 32'h42b530eb},
  {32'hc4fec2cd, 32'h43b3d2fa, 32'hc37dc46f},
  {32'h44b13d65, 32'hc1aad027, 32'hc30b821f},
  {32'hc44f0679, 32'hc269afe2, 32'h428b9afd},
  {32'h4495da0e, 32'h438b42e3, 32'hc340ca11},
  {32'hc357dcdd, 32'h419c77ac, 32'hc312cc1a},
  {32'h449ae03a, 32'hc28bc56c, 32'hc2bc2044},
  {32'hc4335f31, 32'hc2b87a15, 32'hc28005bf},
  {32'h43eddcc4, 32'hc2d90130, 32'h42e19c80},
  {32'hc447f36a, 32'hc3685e5c, 32'h4340b229},
  {32'h44a1b676, 32'h436da2df, 32'h4299e784},
  {32'hc5255a23, 32'hc2ba2204, 32'h4360140d},
  {32'h44b12c8c, 32'h42b719ba, 32'h432ebe7e},
  {32'hc4dfac7c, 32'h41b1c86b, 32'h43ba48cd},
  {32'h44e91f84, 32'h42771c23, 32'hc2962022},
  {32'hc47492fc, 32'h432bfbd5, 32'h429dfe20},
  {32'h44922742, 32'hc391995f, 32'hc33fe5b2},
  {32'hc472bf33, 32'hc31fc484, 32'hc3030f03},
  {32'h44935525, 32'h42dd39f9, 32'h4323917c},
  {32'hc4f32a37, 32'hc239b20a, 32'hc11d349c},
  {32'h45066786, 32'hc262b544, 32'h43a845f9},
  {32'hc4c1545d, 32'h42912fd4, 32'hc3093787},
  {32'h44f2b87d, 32'hc2fd6353, 32'hc2bc67dc},
  {32'hc4213cb8, 32'hc3bb7c09, 32'h438ad0de},
  {32'h43e1c75c, 32'hc35be053, 32'h43cdcb35},
  {32'hc4bf68ff, 32'h43489fec, 32'hc381663d},
  {32'h44a7e768, 32'hc3b3d506, 32'h4379c2e5},
  {32'hc410e628, 32'hc40a8184, 32'h43842885},
  {32'h43953920, 32'h41c983fa, 32'hc2be2f90},
  {32'hc4ffdba9, 32'hc140cf75, 32'h432a696b},
  {32'h4322a244, 32'h42d7471d, 32'h4357a9bc},
  {32'hc4b93e9b, 32'h4222d3bd, 32'hc1178f22},
  {32'h447f5054, 32'h425d8faa, 32'hc39b2e15},
  {32'hc347970c, 32'h4381b1bb, 32'h432f9c80},
  {32'h4430273e, 32'h428d9320, 32'h436ae883},
  {32'hc50147c5, 32'h443dd3b2, 32'h43aefc2f},
  {32'h45304a1b, 32'hc252bdf7, 32'h42bedd24},
  {32'hc4f88313, 32'hc2ab8c4f, 32'hc2c6895e},
  {32'h44418c2a, 32'h42d695cd, 32'h42b5d317},
  {32'hc50884e4, 32'hc2810e0f, 32'hc213b727},
  {32'h44e43f73, 32'hc321c6c4, 32'hc3746ac3},
  {32'hc4a7d4f4, 32'hc3c106f7, 32'h42f27f1e},
  {32'h44f1bf12, 32'hc31e860c, 32'h435762a7},
  {32'hc4e18618, 32'hc40a2f15, 32'hc41b6a67},
  {32'h44fc2f86, 32'h42154c02, 32'hc315e5ef},
  {32'hc4c96689, 32'hc23317ff, 32'h4324843b},
  {32'h440e87e4, 32'hc215cb3c, 32'hc30b7ca6},
  {32'hc47332bc, 32'hc37a5567, 32'h41d3e159},
  {32'h44a4d00e, 32'hc3ad8a26, 32'h428cf357},
  {32'hc3a141a6, 32'h435177dc, 32'hc29a8005},
  {32'h44903476, 32'h418c43dc, 32'hc30c1786},
  {32'hc4384d95, 32'h41d9227a, 32'hc36444ff},
  {32'h45215fa3, 32'hc2d5e6bd, 32'hc3480ff1},
  {32'hc4d95521, 32'h432cc2ba, 32'h4390887d},
  {32'h44bc9a6e, 32'h41f5b73f, 32'h438d3240},
  {32'hc432ebd7, 32'hc2e506bd, 32'h420ab080},
  {32'h43bb876c, 32'h42ffa7f4, 32'hc2290573},
  {32'h4291ae60, 32'h425d2184, 32'h437e1ce7},
  {32'h4481fd08, 32'h428da491, 32'hc2c6251a},
  {32'h43d132c8, 32'hc39281da, 32'hc274175f},
  {32'h44f2c966, 32'hc21c26e3, 32'h439992c0},
  {32'hc4991762, 32'h44109323, 32'h42c4d099},
  {32'h44e2d310, 32'h432ab8cf, 32'h4267be12},
  {32'hc279d7dc, 32'hc2c5c770, 32'h434769ad},
  {32'h4481dfc0, 32'h431af26a, 32'hc214ca6d},
  {32'hc4ade355, 32'h42ca6e47, 32'h43a49698},
  {32'h44fdbfb1, 32'h433aaebb, 32'hc2cbc7f4},
  {32'hc48db06c, 32'hc329eb44, 32'hc3122946},
  {32'h44929d3e, 32'hc32fafc1, 32'h40d18d1e},
  {32'hc2aef32d, 32'hc3541168, 32'h41f5eb1a},
  {32'h44406bf0, 32'hc38ffebc, 32'h42f41226},
  {32'hc446236e, 32'h42172ba5, 32'hc2603c47},
  {32'hc1854a00, 32'hc38a3855, 32'hc2e24bdf},
  {32'hc3f96be4, 32'h43181815, 32'h419f3956},
  {32'h42b63780, 32'h42bcb6a2, 32'hc3238f2e},
  {32'hc501f911, 32'hc2bb66b5, 32'hc2931ce8},
  {32'h4433eafc, 32'hc3ba7c4f, 32'h40bc909f},
  {32'hc4a884aa, 32'h436ac5da, 32'h43a4e27f},
  {32'hc2606680, 32'hc2a77471, 32'hc1b6cfa5},
  {32'hc311640c, 32'h436580d8, 32'hc3c5b1d8},
  {32'h43dc196c, 32'hc30a9ca0, 32'h43d6dd3e},
  {32'hc519fe3b, 32'h42a51db3, 32'hc0151324},
  {32'h44f50eee, 32'hc39c1b91, 32'h43d39f10},
  {32'h40532400, 32'h430ba002, 32'hc3164278},
  {32'h442bb1b4, 32'hc2ca1e69, 32'h41cfb9b8},
  {32'hc3e40f78, 32'hc38215ca, 32'h42e2ae77},
  {32'h442c9860, 32'h43587cc9, 32'hc16a1c8c},
  {32'hc43392d1, 32'hc3971cf2, 32'h43a6704f},
  {32'h450b7f3f, 32'hc3b76754, 32'h438074e1},
  {32'hc48d1535, 32'hc337d68c, 32'h432a9cda},
  {32'h4442dc7c, 32'hc2a816cd, 32'h4327654a},
  {32'hc506553a, 32'h42ecdba8, 32'hc31be6f6},
  {32'h451fe44b, 32'hc3c04483, 32'hc403cf61},
  {32'hc3993dda, 32'h42885459, 32'hc403b629},
  {32'h440a9166, 32'h42b6ca80, 32'hc2a81fe8},
  {32'hc4fde056, 32'hc326ecda, 32'h42510a73},
  {32'h451c1576, 32'hc227df57, 32'hc28a8363},
  {32'hc5055ecd, 32'h438fdd3a, 32'hc394ccb5},
  {32'h44914855, 32'h42d5705e, 32'hc344479c},
  {32'hc443ffb9, 32'hbf3efc80, 32'h41a4f900},
  {32'h44d458b6, 32'hc2b3da70, 32'hc41043f3},
  {32'hc4c1a43a, 32'hc33eadc7, 32'h43bb4ff8},
  {32'h44379850, 32'hc2b23e8b, 32'h415342e8},
  {32'hc5082936, 32'hc380b0b5, 32'h4367969a},
  {32'h44ed62bc, 32'h433b6518, 32'h420c7d44},
  {32'hc4529328, 32'hc3dab1f9, 32'hc410cbb8},
  {32'h44f017f6, 32'hc2f8548b, 32'h424c801b},
  {32'hc4eeac34, 32'hc34bcf93, 32'hc319b277},
  {32'h44c247a9, 32'hc2fd6930, 32'h435dc48d},
  {32'hc48389a9, 32'hc26fc390, 32'hc40e5887},
  {32'h43e5a4c8, 32'hc36ef67a, 32'hc30d4dbe},
  {32'hc50beb12, 32'hc29c96b6, 32'hc368653e},
  {32'h44c85d12, 32'hc2639b7c, 32'h43dbd551},
  {32'hc4fcf6fd, 32'h438ebd8c, 32'h430e0286},
  {32'h44cad934, 32'h43bd6783, 32'hc3234184},
  {32'hc4fb47fa, 32'hc33e4895, 32'hc2c77ed8},
  {32'h44b79a63, 32'h4230fdc0, 32'h42628714},
  {32'hc4e55367, 32'hc2550a96, 32'hc2bde7c5},
  {32'h4492e9d5, 32'hc4291560, 32'hc414a576},
  {32'hc47a69a4, 32'h4258cae7, 32'h42c7d16e},
  {32'h438ec93b, 32'hc2c80514, 32'h4319da66},
  {32'hc49ed576, 32'hbf829d34, 32'h4280eb49},
  {32'h439f96d5, 32'h432e3eec, 32'hc3c001c8},
  {32'hc4344180, 32'h42f1a4d8, 32'hc35e029a},
  {32'h44edf67b, 32'h433dbc3c, 32'hc29313cf},
  {32'hc4a51ecb, 32'h438b4065, 32'h435aa61d},
  {32'h43ddf291, 32'h42466927, 32'hc3568974},
  {32'hc4c5b066, 32'h42d8e230, 32'h42963d33},
  {32'h44b38fbe, 32'h40d9322e, 32'h4210e3b0},
  {32'hc508e035, 32'h42ec56f5, 32'h4319a971},
  {32'h450c2bda, 32'h42b92380, 32'hc184fd38},
  {32'hc3caaf97, 32'hc35b36e1, 32'hc38444a3},
  {32'h44de6233, 32'h3f91010d, 32'hc08a3f4b},
  {32'hc2f10923, 32'h435bbc36, 32'h432c469d},
  {32'h44157a90, 32'hc24afa04, 32'h436ab858},
  {32'hc3057470, 32'h42614264, 32'hc31225a5},
  {32'h4510ad26, 32'hc374371a, 32'h409c388c},
  {32'hc349044a, 32'h42f09865, 32'h43286408},
  {32'h450d026e, 32'h43152590, 32'hc38426b9},
  {32'hc4c1bf3e, 32'h427463ac, 32'hc31fac19},
  {32'h44b9bd8a, 32'h435509ef, 32'hc0bd2470},
  {32'hc4d63965, 32'hc328d780, 32'hc282c956},
  {32'h44d34601, 32'hc23bc990, 32'hc3146005},
  {32'hc4da8a2d, 32'hc31f60b1, 32'h4296c28b},
  {32'h44a6d531, 32'h42a50aab, 32'h42f4fb04},
  {32'hc2994e2c, 32'h4321660f, 32'h42f898d7},
  {32'h4456f9c5, 32'hc344c5e5, 32'h425b0ee6},
  {32'hc38e872a, 32'hc3ae59f0, 32'h42e89358},
  {32'h450be452, 32'h42755315, 32'hc2e3519c},
  {32'hc4b08a0a, 32'h4236c5ca, 32'hc3646b88},
  {32'h44f50123, 32'hc382d4d4, 32'hc23f88c5},
  {32'hc4b1cbf6, 32'h4050f9fa, 32'hc18f4129},
  {32'h43a05913, 32'h43dc8eca, 32'h4338f537},
  {32'hc518628b, 32'hc28f2aea, 32'h43971749},
  {32'h45177403, 32'hc3358a99, 32'h42f772da},
  {32'hc3ba4925, 32'hc2b5d8e0, 32'hc3e31364},
  {32'h450d2066, 32'h40584dc4, 32'hc300a753},
  {32'h43f6dd08, 32'h43e2130f, 32'hc410c355},
  {32'h4507e145, 32'hc25b3ac1, 32'h430c697d},
  {32'hc41f0bc4, 32'hc3073fa7, 32'h418f482f},
  {32'h423ae4d0, 32'h42839600, 32'h436f720d},
  {32'hc4e4159d, 32'hc1f9a229, 32'h420871cb},
  {32'h449994b9, 32'h42a1bf1b, 32'hc2c87922},
  {32'hc4f7f722, 32'h42d7d7d1, 32'h422c7438},
  {32'h448e48ff, 32'h43b0a317, 32'hc13b179f},
  {32'hc51c30e4, 32'h425d87df, 32'h40a5de48},
  {32'h44902329, 32'h434c5990, 32'hc2d3ca27},
  {32'hc47ee932, 32'hc2949dbf, 32'h422dd190},
  {32'h410ea240, 32'h40d37b6c, 32'h4103c7d4},
  {32'hc508bc40, 32'h438cd3dd, 32'h41cec905},
  {32'h44ae8d04, 32'h436cde8a, 32'hc2284f3b},
  {32'hc292ea6c, 32'hc323bf6b, 32'hc4010cd3},
  {32'h4512dcc3, 32'hc2ce3ab4, 32'hc2fb10b0},
  {32'hc34ad843, 32'h421b38e2, 32'hc3683537},
  {32'h4513fae9, 32'hc2fff083, 32'h4373747d},
  {32'hc5147d75, 32'hc32a628a, 32'h4304f434},
  {32'hc215c120, 32'hc26a5ce1, 32'hc1ccc320},
  {32'hc5004647, 32'hc298a7be, 32'h43331d99},
  {32'h44fa6c1e, 32'h4063f7b6, 32'hc3b94188},
  {32'hc48224b0, 32'h4352430e, 32'h42d4826b},
  {32'h44fc72e6, 32'h42fa23b5, 32'h4334427c},
  {32'hc4dad35d, 32'hc28fd67d, 32'h411a43ba},
  {32'h3eaa9600, 32'hc39f76aa, 32'h4362b00c},
  {32'hc3374748, 32'hc361f6d9, 32'h4311ca69},
  {32'h445d1398, 32'hc31e568f, 32'hc2904097},
  {32'hc4947a6c, 32'hc380bb32, 32'h424d483c},
  {32'h443604f9, 32'hc32c13e4, 32'hc2bb260c},
  {32'hc4c78686, 32'hc3a52b31, 32'hc31dc8bf},
  {32'h4502efcc, 32'h4328059a, 32'hc30d8f9b},
  {32'hc4303999, 32'h4259c1b6, 32'h420fcbfe},
  {32'h44d20226, 32'h4303dc5d, 32'hc2e8ef7c},
  {32'hc4f06fe1, 32'hc2783faa, 32'h42b84eab},
  {32'h44e73e38, 32'h43163a06, 32'h4112f788},
  {32'hc4ecce5a, 32'hc2d8a720, 32'h432b6bda},
  {32'h449f36c4, 32'hc173503f, 32'h42987232},
  {32'hc4fbd68f, 32'hc3129f09, 32'h4263eca5},
  {32'h448ef90e, 32'hc26a8415, 32'h43a49063},
  {32'hc501591e, 32'hc2fa5c6b, 32'hc37905d5},
  {32'h44535d44, 32'hc2540a63, 32'hc3cb6be7},
  {32'hc46632ed, 32'h4299a084, 32'hc36f2da9},
  {32'h44881802, 32'h43d6380a, 32'h43a5ed58},
  {32'hc301b55f, 32'h437a88d5, 32'hc2ce4dcc},
  {32'h442fe74f, 32'h428572e6, 32'h4396dee9},
  {32'hc46c89f7, 32'hc436932a, 32'hc2948f3a},
  {32'hc4fac4bd, 32'hc22b8948, 32'h422c7a15},
  {32'h44ba2270, 32'h4232552b, 32'h42e5c5bb},
  {32'hc4b45c26, 32'h441f72ba, 32'hc3baf8ae},
  {32'h448f31c0, 32'h43bc4529, 32'h4011ca3c},
  {32'h42737c16, 32'hc3c13a9e, 32'hc3437543},
  {32'h44057b17, 32'h4339455c, 32'hc32f1d4d},
  {32'hc509b47f, 32'h431222bb, 32'hc386130f},
  {32'h448b6338, 32'hc07a6738, 32'h43d45b54},
  {32'hc39ec626, 32'h429cb002, 32'h431ea982},
  {32'h445614b6, 32'h426ad878, 32'hc295b419},
  {32'hc481742d, 32'h4399e556, 32'hc3d86b10},
  {32'h4411906e, 32'hc38a611a, 32'hc2ebe899},
  {32'hc3e29aa8, 32'h43653df7, 32'hc34a4c52},
  {32'h45015e0e, 32'h417625e8, 32'h42adf6db},
  {32'hc3b073a5, 32'h43d690e2, 32'h423c1062},
  {32'h449618a6, 32'h43287b9e, 32'h43156364},
  {32'hc5090ee4, 32'hc32b0c6e, 32'h429fafa0},
  {32'h450250cc, 32'h4384a3cf, 32'h434becce},
  {32'hc4c6a912, 32'h42973c04, 32'hc2cd9cc8},
  {32'h445e8662, 32'hc30a3b2c, 32'hc36da73e},
  {32'hc4da7e82, 32'h42cbf050, 32'hc2fc6241},
  {32'h44404dc4, 32'h43398a8c, 32'h439bacea},
  {32'hc460a830, 32'hc1bcd95c, 32'h435e256e},
  {32'h43b19e9f, 32'h42261c6d, 32'hc2e71b50},
  {32'hc41e9f7e, 32'hc3dc6bbf, 32'hc3545832},
  {32'h4437a1d1, 32'h4317f71e, 32'hc316cddf},
  {32'hc49390d6, 32'hc105def8, 32'hc2f94510},
  {32'h44961c69, 32'h438d0e97, 32'h42a86969},
  {32'hc00ba8c0, 32'hc29dc939, 32'hc303b0bd},
  {32'h4426accc, 32'hc3719f3b, 32'hc3849276},
  {32'hc27e6a19, 32'h433c7115, 32'hc24a9c73},
  {32'h44ea7584, 32'h42916e20, 32'h43546907},
  {32'hc42e7be4, 32'hc36aee44, 32'h432fbae6},
  {32'h4469868e, 32'hc29c96e3, 32'hc2da488b},
  {32'hc434ec6e, 32'hc13a85d7, 32'hc36b0483},
  {32'h4513dca2, 32'hc2dfcdb7, 32'h43920a0e},
  {32'hc5032205, 32'hc3c174f1, 32'hc395e563},
  {32'h450baead, 32'hc3651f52, 32'h430be868},
  {32'hc4e90518, 32'h4223c38c, 32'h424c2c70},
  {32'h44e18aef, 32'h430401e2, 32'h435429c9},
  {32'hc4ef0cc8, 32'hc3f90d43, 32'hc2124788},
  {32'h40a68500, 32'h434620e3, 32'h423b739b},
  {32'hc502c741, 32'h429add93, 32'hc05c3c0f},
  {32'h44e69429, 32'hc33e4d81, 32'h43cba382},
  {32'hc4e87594, 32'h43a3a6ec, 32'h431f9923},
  {32'h445b786c, 32'h430d8c9e, 32'h43aceb17},
  {32'hc512fcee, 32'h42c70edd, 32'h439da8e9},
  {32'h44f31b6e, 32'h4391752c, 32'h42a14622},
  {32'hc4f303db, 32'h43575e38, 32'hc2af1595},
  {32'h450034c7, 32'h433f1352, 32'hc2883a66},
  {32'h42b8b8e0, 32'hc2eb1663, 32'h3fecbb20},
  {32'h44c418a4, 32'hc2b2b965, 32'h43712853},
  {32'hc5172878, 32'hc3da1ce5, 32'hc29f9d98},
  {32'h4502b70d, 32'hc401b58a, 32'h438ccb91},
  {32'hc4b59d8c, 32'hc394300b, 32'h42b1d1da},
  {32'h4518bc9c, 32'h40cfd1b2, 32'h427ccbb0},
  {32'hc39dd100, 32'h4284cb9a, 32'hc39af719},
  {32'h44cad91c, 32'hc0bf0ba0, 32'hc19ad9b8},
  {32'hc3d1ad90, 32'hc34548c6, 32'hc3f05ec1},
  {32'h44909f0e, 32'h431fa336, 32'h42ba5d82},
  {32'hc4695154, 32'hc3dc0350, 32'hc403661c},
  {32'h44218106, 32'h41dda2e5, 32'h438f0ec7},
  {32'hc4fc7f7a, 32'h4368e62e, 32'h438c1ded},
  {32'h45060d76, 32'h42d11d9e, 32'h42c84157},
  {32'hc4b9e378, 32'h42ba56f4, 32'h43600a19},
  {32'h44ecb226, 32'hc24bc16b, 32'hc382e7d3},
  {32'hc4a5c7b1, 32'hc309566a, 32'h42c14b90},
  {32'h4410e2a0, 32'h431112a6, 32'hc3d45f81},
  {32'hc515397b, 32'hc318cec1, 32'hc3729a41},
  {32'h444b4090, 32'h43147bbe, 32'hc33b2cdb},
  {32'h439f3512, 32'h413e6567, 32'hc138a214},
  {32'h44811242, 32'h42552d9e, 32'h42c939ea},
  {32'hc44fec00, 32'hc2003ef4, 32'h42cf2939},
  {32'h44b072f0, 32'h4185e478, 32'h439f0c7f},
  {32'hc4c9d0ab, 32'hc36bd355, 32'h4376aaad},
  {32'hc2dac0b8, 32'h418409de, 32'hc3b9a88f},
  {32'hc4372f80, 32'hc314c064, 32'h4236e439},
  {32'h44978e1e, 32'hc3cbf9aa, 32'hc3790e34},
  {32'hc4ebee9e, 32'hc3116ecd, 32'h4106bf33},
  {32'h44fdb32a, 32'h43eff0d0, 32'hc29f3b91},
  {32'hc3747b02, 32'hc35c5cb0, 32'hc2055eff},
  {32'h4514af50, 32'h4239025c, 32'h414b2077},
  {32'hc4ba737a, 32'hc312307c, 32'h4219e88a},
  {32'h45063a17, 32'h443c0db9, 32'h416ca0b2},
  {32'hc4f24c30, 32'hc2041f6e, 32'hc2db58f6},
  {32'h4492d6a9, 32'hc385a287, 32'h430a5590},
  {32'hc47e9bcc, 32'h41582268, 32'h4240cfe5},
  {32'h443ee696, 32'hc36a9b61, 32'h4328fa97},
  {32'hc4202577, 32'hc297da52, 32'h438b77e2},
  {32'h44cbdd78, 32'h4384c883, 32'hc33f308a},
  {32'hc3b63be8, 32'h43031889, 32'hc39f02ce},
  {32'h44a6f4e7, 32'hc24c5451, 32'hc21a9802},
  {32'hc3e81938, 32'h4382372c, 32'h4376e2f5},
  {32'h445e8ea2, 32'hc317d2b1, 32'hc24509d1},
  {32'hc414a60e, 32'h427db39e, 32'h4308f6f6},
  {32'h44898a71, 32'h41fd491f, 32'hc2c55def},
  {32'hc48f62f5, 32'h439d4d4a, 32'h41459c10},
  {32'h4446509f, 32'hc3629cf3, 32'hc24b7b92},
  {32'hc3958fc4, 32'h431d7749, 32'hc3140307},
  {32'h44829f74, 32'hc3bda939, 32'h435ec77f},
  {32'hc3614ee8, 32'hc2fcd65f, 32'hc32ea943},
  {32'h43d25ecc, 32'h42fd6626, 32'hc34b33c4},
  {32'hc49f3e06, 32'h43bd4721, 32'hc358db10},
  {32'h441a39dc, 32'h42da1b62, 32'h42df5551},
  {32'hc4b41466, 32'hc39e4976, 32'hc38049fd},
  {32'h444abc90, 32'h42b3dfac, 32'hc28a02a1},
  {32'h437f581e, 32'hc29696b6, 32'hc27791a2},
  {32'h44bb9870, 32'hc291f81a, 32'h42f46a2f},
  {32'hc4bc653e, 32'hc386f266, 32'hc210dc4a},
  {32'h44f9e196, 32'h4324faa3, 32'h430477a6},
  {32'hc499c323, 32'hc28de8ec, 32'h430d8e6e},
  {32'h447536d9, 32'hc333f1c1, 32'hc1b930b2},
  {32'hc4e35512, 32'h43b82729, 32'h43413a31},
  {32'hc2b1fd68, 32'hc24e276e, 32'h43e916a6},
  {32'hc5118f46, 32'hc220b7fc, 32'h437b841f},
  {32'h44ea90c0, 32'hc3379833, 32'hc2290329},
  {32'hc4b67fce, 32'hc329705d, 32'h43f7eb74},
  {32'h4506ad98, 32'h42990b18, 32'hc227ba4a},
  {32'hc4efb57b, 32'h43611fd6, 32'h42c48659},
  {32'h450c9202, 32'hc1b3ce4a, 32'h42e9fd3e},
  {32'hc4961b01, 32'h43759f15, 32'hc1d6e84e},
  {32'h44a123be, 32'h3f64b79a, 32'hc313abcc},
  {32'hc30f8b67, 32'h42539061, 32'hc230ad6b},
  {32'h428d8d10, 32'h42ffd952, 32'hc09a8708},
  {32'hc449ca9e, 32'h43870da3, 32'h4338010d},
  {32'h4491983b, 32'h42f8f2bc, 32'hc3860547},
  {32'hc404b540, 32'hc332a6c7, 32'hc276dfae},
  {32'h447349cc, 32'hc3a326a2, 32'hc1f4ff50},
  {32'hc4cfe462, 32'hc317b095, 32'h42a12ab1},
  {32'h44240a3b, 32'h44065e3e, 32'hc38b985d},
  {32'hc43d5b4e, 32'hc2a78bbb, 32'hc377d2e9},
  {32'h44c35797, 32'hc26c25f2, 32'h430d7385},
  {32'hc35d2b90, 32'h439039d0, 32'h42b029e0},
  {32'h4501e5f4, 32'h4363716a, 32'hc345f240},
  {32'hc4d47ccd, 32'hc0bc7113, 32'hc41615d8},
  {32'h443489da, 32'hc3c30bf7, 32'hc39686a5},
  {32'hc467e9e7, 32'h432fa268, 32'hc29a9402},
  {32'h44136d7d, 32'hc355f486, 32'h40d79a1b},
  {32'hc3a7fc2c, 32'hc3fe7542, 32'h42e983eb},
  {32'h4289f526, 32'h42f02c46, 32'h4268c1f1},
  {32'hc4f178c4, 32'h435ce901, 32'hc2c9470d},
  {32'h44911742, 32'h443c898a, 32'h433c7be6},
  {32'hc495d8d8, 32'h4321f12f, 32'hc2993d3d},
  {32'h44ac3591, 32'h43463e4e, 32'hc3173fb7},
  {32'hc4c3348e, 32'hc2cb30cc, 32'h3f435240},
  {32'h450bbb64, 32'hc4061eb5, 32'h4384e131},
  {32'hc414bfce, 32'hc33e1b41, 32'h4366c29e},
  {32'h43adb772, 32'h42a2da64, 32'hc2e036d1},
  {32'hc4bda354, 32'h4381d427, 32'hc3260355},
  {32'h44eb638d, 32'h4229248a, 32'hc2ae4b32},
  {32'hc4fbefb3, 32'hc3109a8b, 32'hc32beb28},
  {32'h438df419, 32'hc3bbbecb, 32'hc1a95b60},
  {32'hc506d36c, 32'hc38e65c6, 32'h42c6d5bc},
  {32'h42326562, 32'h414a7844, 32'h43333b84},
  {32'hc49cab63, 32'hc1b60a13, 32'h4335c3cb},
  {32'h43a5fbbc, 32'h41772ab7, 32'hc2e63686},
  {32'hc48cf05d, 32'hc37b976b, 32'h433242a1},
  {32'h4433f0ce, 32'h43346c5a, 32'hc1f7cda6},
  {32'hc3ce59ae, 32'h438bea59, 32'hc2135249},
  {32'h45146412, 32'hc34f29c6, 32'hc358518d},
  {32'hc3fd5a8f, 32'hc3bea22e, 32'hc3896192},
  {32'h4429e114, 32'hc2f2c593, 32'hc22a54c8},
  {32'hc49732e2, 32'hc2a7911a, 32'h43374155},
  {32'h44d5986d, 32'hc3af34ae, 32'h4378df31},
  {32'hc4b0540a, 32'hc2ff3efc, 32'h421f8bd2},
  {32'h44c24bd2, 32'hc064d275, 32'h42def935},
  {32'hc350c138, 32'h426e998c, 32'h40f80f46},
  {32'h43164030, 32'h42b5e2b0, 32'h4136cae8},
  {32'hc501a990, 32'h43bd16bc, 32'hc373ae72},
  {32'h44f48fb9, 32'hc387e75c, 32'h418b6778},
  {32'hc4a48f1d, 32'hc0bee7b2, 32'hc0af627a},
  {32'h44ebe832, 32'h43187963, 32'h436457dc},
  {32'hc4a9e8cb, 32'h437d041a, 32'hc23fcc93},
  {32'h441fedb0, 32'hc2cb2a3a, 32'hc3ea2d0f},
  {32'hc4dbf83c, 32'hc342e006, 32'h42cbf913},
  {32'h4492564e, 32'h43ab7347, 32'hc1d9bb6f},
  {32'hc4cf8014, 32'hc107af97, 32'hc0e2883a},
  {32'h44c6e7ad, 32'h412329db, 32'h42dde68e},
  {32'hc49803a2, 32'hc4082e4c, 32'h43c17e48},
  {32'h4359e32a, 32'hc20ee2be, 32'hc461be41},
  {32'hc4c5b67e, 32'hc3358870, 32'hc292a7bb},
  {32'h42a97e70, 32'h43c73d97, 32'h40658bec},
  {32'hc4df93e7, 32'h411d723f, 32'hc12d76f8},
  {32'h447c3e74, 32'h44117429, 32'h439b7945},
  {32'hc3fce8e4, 32'hc3cb924e, 32'hc2963692},
  {32'h45036f8d, 32'hc34237cb, 32'h43730626},
  {32'hc4972e0e, 32'hc3a69c64, 32'h42e113f1},
  {32'h44686790, 32'hc296cfb7, 32'hc2dbc14e},
  {32'hc45864d3, 32'h436c0eff, 32'h431dc321},
  {32'h44ff2224, 32'hc3f06209, 32'hc392e7f1},
  {32'hc498c05b, 32'h439b102a, 32'hc2de9396},
  {32'h44ad1850, 32'h40a3af8a, 32'h4369e226},
  {32'hc4b01104, 32'hc0564302, 32'hc1975d3a},
  {32'h446f61a8, 32'h42f12a64, 32'h43391e44},
  {32'hc3961fa0, 32'h4335ba3d, 32'h436bd4e0},
  {32'h449c77dd, 32'h436adec8, 32'hc3525e46},
  {32'hc4d1daca, 32'hc392e7ee, 32'h430e6541},
  {32'h448f2b2a, 32'h43baa142, 32'h42bd50fb},
  {32'hc493d106, 32'h427469a0, 32'h4139203a},
  {32'h44ed4f32, 32'hc3a53b73, 32'h4380a24f},
  {32'hc2ca25f4, 32'h41ce04a2, 32'h435dfd97},
  {32'h449bc4da, 32'hc29f3ff2, 32'h4310db24},
  {32'hc50d7643, 32'hc340b010, 32'h43bdfb81},
  {32'h44e5fe0f, 32'hc2dd1713, 32'h410cfece},
  {32'hc2a93880, 32'hc337ab48, 32'h4391a34b},
  {32'h44503dfb, 32'h42c53003, 32'hc19b9a6b},
  {32'hc3b063d0, 32'hc2ce0a4e, 32'hbf9e21b0},
  {32'h445d2e1a, 32'h4294b432, 32'hc3cfb4ba},
  {32'hc42c1150, 32'h43a26f89, 32'hc403b2a0},
  {32'h430aabff, 32'hc2a3c365, 32'h41b50216},
  {32'hc512ee76, 32'h42c04dbd, 32'h44187eb8},
  {32'h4453a37a, 32'h43610315, 32'h43c4871c},
  {32'hc49a6c43, 32'h432f5b88, 32'h42e5f71e},
  {32'h44f2e799, 32'h438d2c13, 32'h43746379},
  {32'hc41e48ec, 32'hc2cfddc5, 32'h43b28646},
  {32'h44cacefc, 32'h4381441f, 32'hc3c17dab},
  {32'hc4587424, 32'hc2dbad46, 32'hc3a2fd6a},
  {32'h450bdffa, 32'hc346deae, 32'hc2ea9f28},
  {32'hc46df3ea, 32'h418dfefc, 32'hc38f4b67},
  {32'h45117358, 32'h4321ae6e, 32'h43a6d375},
  {32'hc46a5de2, 32'hc305d35e, 32'hc29c6167},
  {32'h44cc7959, 32'h42907850, 32'hc2011a26},
  {32'hc4fe94ef, 32'hc34d6e61, 32'hc3af25b2},
  {32'h44d2e532, 32'h4331742e, 32'h4302bf8b},
  {32'hc4f57782, 32'h43697313, 32'h42576262},
  {32'h44790a96, 32'hc36ac9bf, 32'h42d30e12},
  {32'hc34c4611, 32'hc4032a44, 32'hc386b9c1},
  {32'h448d5bd8, 32'hc2abd9e2, 32'h431e1327},
  {32'hc3c7be8b, 32'hc2c4929b, 32'h4102b539},
  {32'h450889b9, 32'hc3388231, 32'h43636258},
  {32'hc4e3abaa, 32'hc1da155a, 32'h42ae6ce4},
  {32'h43fd0b32, 32'hc0a1d2b6, 32'h42fbfba4},
  {32'hc43a24c8, 32'hc364dbe4, 32'h419a739e},
  {32'h44d112f7, 32'h43520f46, 32'hc3af676c},
  {32'hc4b21a79, 32'hc2e87907, 32'h429c5bc5},
  {32'h4515a4a8, 32'hc35026d6, 32'h43acebb6},
  {32'hc49697bc, 32'hc2bf9400, 32'h42a32506},
  {32'h443d172e, 32'h4303b41e, 32'h431f4edd},
  {32'hc4e45f05, 32'h42ee52ec, 32'hc38f061e},
  {32'h4404ccee, 32'hc21bc186, 32'hc270bb4a},
  {32'hc511a79e, 32'hc324a036, 32'hc2955b96},
  {32'h440ba27a, 32'hc22d12ec, 32'hc3c5cb18},
  {32'hc4154d38, 32'h42bd8e17, 32'h41c0ceb1},
  {32'h44eb90d0, 32'hc29c0d17, 32'h43008df7},
  {32'hc4ab04ab, 32'h4308e705, 32'h416f2196},
  {32'h4472d669, 32'hc28ae4d0, 32'hc1df7df0},
  {32'hc469fff4, 32'h439c42ed, 32'hc26bd9d2},
  {32'h448188f6, 32'hc2b8be29, 32'hc315b75c},
  {32'hc4770867, 32'hc30669ee, 32'hc2ddee64},
  {32'h450c7620, 32'h433a1230, 32'h41e8e8b1},
  {32'hc48375ea, 32'hc2f3dd67, 32'h435a4122},
  {32'h43adc2bb, 32'h42512347, 32'h42650b18},
  {32'hc491b788, 32'hc349c730, 32'h430d8188},
  {32'h44c2708b, 32'hc1bdef20, 32'h428e3b95},
  {32'hc42b2c56, 32'hc3269937, 32'hc2e65f87},
  {32'h44b96af6, 32'h439dc623, 32'h428efa66},
  {32'hc467651e, 32'hc30a8447, 32'h432ab711},
  {32'h43a2c5e8, 32'h43827f98, 32'hc3bd53aa},
  {32'h44325d5d, 32'hc2841a37, 32'h41f5c02c},
  {32'h44af3e77, 32'h42b4f538, 32'h430249f9},
  {32'hc38a2664, 32'hbf968462, 32'h4371a222},
  {32'h449d2466, 32'h42cec1ce, 32'hc3264303},
  {32'hc4f63b38, 32'hc399594d, 32'h41fd0bb7},
  {32'h4513378e, 32'h432e832e, 32'h4339d6c4},
  {32'h4323d55d, 32'h42b35863, 32'hc316b774},
  {32'h44279f98, 32'h42ac2745, 32'h4395ad47},
  {32'hc40ebb0c, 32'hc1ed8ee2, 32'h40f6340a},
  {32'h4519b728, 32'h42ac391c, 32'h431405e0},
  {32'hc4e8ec5d, 32'hc2b4abe5, 32'h43af7ab1},
  {32'h42e9fa20, 32'h42864a44, 32'hc315fc51},
  {32'hc3e6cf98, 32'h42644a38, 32'hc11fa21e},
  {32'h4471b21a, 32'h42fd98c0, 32'h429d6cff},
  {32'hc51444dc, 32'h4376f9f6, 32'hc3279226},
  {32'h443ba8bc, 32'h44078f61, 32'hc2ae3eac},
  {32'hc483d015, 32'hc2b77d03, 32'hc31bd97e},
  {32'h43783687, 32'h427f4c53, 32'hc3800ecf},
  {32'hc51cd51a, 32'h4321fd9d, 32'h429f46cc},
  {32'h4351d79c, 32'h420c3b12, 32'h435c7a27},
  {32'hc4f74996, 32'h3f01339c, 32'h42429568},
  {32'h44c2f740, 32'h43790d79, 32'hc32aab54},
  {32'hc4766dd9, 32'hc336d168, 32'hc3692439},
  {32'h446dbb72, 32'h421155b2, 32'h433657d0},
  {32'hc391d3e0, 32'hc2dfc714, 32'h43588cf8},
  {32'h44c9a260, 32'hc35780f1, 32'h4312e3ac},
  {32'hc4c189c7, 32'h40384b40, 32'hc3133718},
  {32'h450c98aa, 32'h43a938cc, 32'h4285677c},
  {32'hc49fbdd6, 32'hc3484cb8, 32'hc3ea7323},
  {32'h4352fc0c, 32'h42ffe4e8, 32'h414c60f0},
  {32'hc4abbfdf, 32'hc3b0f686, 32'h43417c00},
  {32'h435282b0, 32'h43485fbb, 32'hc322e032},
  {32'hc5148a68, 32'hc33fe3ba, 32'hc3fb1de9},
  {32'h449b2a26, 32'hc3db28ff, 32'h42eed51c},
  {32'hc4bd1d13, 32'h433ba242, 32'hc2307a23},
  {32'h44fd5b0c, 32'hc2ce3362, 32'hc3cc52f2},
  {32'hc4554535, 32'h441ac9d9, 32'h43833569},
  {32'h4326d866, 32'h431bf42c, 32'h4409eb80},
  {32'hc2ce6c20, 32'hc318b271, 32'h43dd2687},
  {32'hc169fd00, 32'hc2ad7649, 32'h43378e05},
  {32'hc494f99f, 32'h41de6642, 32'hc28c22ff},
  {32'h45131a11, 32'hc2b34031, 32'h43b6e289},
  {32'hc4507886, 32'hc3a98499, 32'hc397e271},
  {32'h44985b56, 32'h43913bf5, 32'hc35f6403},
  {32'hc511e720, 32'hc3c569bd, 32'h4362a300},
  {32'h450b625b, 32'h42c70838, 32'hc37c8b33},
  {32'hc4399bae, 32'h42f66e82, 32'h430d4cbf},
  {32'h44382f3b, 32'hc30e5549, 32'hc2908b7e},
  {32'hc445793d, 32'hc296badd, 32'hc2ab0997},
  {32'h44701ede, 32'hc33db9d5, 32'hc30201d1},
  {32'hc3c4a86c, 32'h43af2e2c, 32'h43c690cb},
  {32'h43b58c16, 32'h43f9f7a2, 32'hc19ead1f},
  {32'h437c2a17, 32'hc3cd84fb, 32'hc131c398},
  {32'h450bc89c, 32'h42f5939a, 32'h3f9ef310},
  {32'hc4b2b83f, 32'h416a64b2, 32'hc328cd34},
  {32'h44f6ef8a, 32'h4315be5c, 32'h43975154},
  {32'hc4aef136, 32'hc407ec37, 32'hc4016d00},
  {32'h446a4140, 32'hc281fc98, 32'h43b3e39a},
  {32'hc3362ca6, 32'hc37b9098, 32'hc33cdb00},
  {32'h4380a5cc, 32'hc3cc09ea, 32'h42c46875},
  {32'hc45497a3, 32'h40fa2a2f, 32'h42e3bdea},
  {32'h44d6e242, 32'hc32e7954, 32'hc15f7de2},
  {32'hc4fa196b, 32'hc2f0f727, 32'hc4010c39},
  {32'h44da1e8e, 32'h42c100e8, 32'hc37eba64},
  {32'hc4675f02, 32'h4384096c, 32'hc157993a},
  {32'h44a44695, 32'h42a43311, 32'h43ad0a2d},
  {32'hc496a50d, 32'hc3680e30, 32'hc3b1170a},
  {32'h432c4e0c, 32'h43cab73c, 32'hc228d5a4},
  {32'hc30d1e0d, 32'hc4167b68, 32'hc25f1faf},
  {32'h45013421, 32'hc3a178e5, 32'h42f9e526},
  {32'hc447f17c, 32'h4308e962, 32'hc266e7e9},
  {32'h42e63f18, 32'h43ac34d5, 32'hc3df6b7e},
  {32'hc4c3095d, 32'hc1ad5d2a, 32'hc204b7b0},
  {32'h435849ac, 32'hc381b625, 32'hc1d156b7},
  {32'hc3ffb298, 32'h43415481, 32'hc3500a64},
  {32'h43c8e4d8, 32'h4194fb4e, 32'hc3065285},
  {32'hc4d78827, 32'h418458e0, 32'hc2bf753a},
  {32'h44958a6e, 32'h42f91efd, 32'hc4094b80},
  {32'hc4d69ec8, 32'hc345b600, 32'h438760d0},
  {32'h44d6c9d8, 32'hc2efa739, 32'hc143beda},
  {32'hc46ba64a, 32'hc35e724e, 32'h4293e960},
  {32'h431aeda5, 32'hc3e484f7, 32'h409de61a},
  {32'hc40aff08, 32'h43730742, 32'hc3332771},
  {32'h45009de4, 32'hc18205c6, 32'hc2ebc158},
  {32'hc506f60e, 32'hc2291f75, 32'hc277f3db},
  {32'h435d1e78, 32'h429bc2ad, 32'h43d483ac},
  {32'hc502e5a8, 32'h422c83bc, 32'hc285f432},
  {32'h44327b35, 32'h435175df, 32'h4088d88f},
  {32'h4316ceea, 32'hc38f5b6c, 32'h435da3d9},
  {32'h44a59742, 32'h4269e37b, 32'hc3aa5ab2},
  {32'hc4420974, 32'hc319c5c8, 32'hc28cd055},
  {32'h42a38570, 32'h426eb5b8, 32'hc31868c0},
  {32'hc47cdcc3, 32'h4229b059, 32'hc1f3ca90},
  {32'h44f55c48, 32'h42b592e8, 32'hc22bd2e4},
  {32'hc3b7a2d9, 32'h42839be5, 32'hc16978ea},
  {32'h44fd2ef0, 32'hc32b98f2, 32'hc35e2483},
  {32'hc3686560, 32'hc3623cec, 32'h42ee8e60},
  {32'h4489356c, 32'hc3734305, 32'hc24c2775},
  {32'h4330a311, 32'hc0291b19, 32'hc33fc692},
  {32'h44ecbced, 32'h43a862bb, 32'hc2ef5aeb},
  {32'hc424770b, 32'hc3b45067, 32'hc3100dfa},
  {32'h44905a4c, 32'h4283d942, 32'h43854eaf},
  {32'hc4e6e84e, 32'hc23dbf18, 32'hc1ee770d},
  {32'h4451b2c4, 32'hc21692c3, 32'h430e20db},
  {32'hc4a1f384, 32'h43be061d, 32'hc387413b},
  {32'h4506115e, 32'h43acea37, 32'hc425dc23},
  {32'hc4f7b82d, 32'hc35948ff, 32'h438b0dc1},
  {32'h44b60136, 32'h433f394d, 32'h42224139},
  {32'hc50b4c49, 32'hc235ee96, 32'h43521db5},
  {32'h43bec230, 32'h42f73bcc, 32'hc235e316},
  {32'hc50059ac, 32'hc275bbdd, 32'h4241ee6e},
  {32'h440343f6, 32'h432d025a, 32'h43402b46},
  {32'hc22b2940, 32'hc3964f6d, 32'h443cad3e},
  {32'h44f16094, 32'h439d51a5, 32'h42bbcb93},
  {32'hc5147be4, 32'hc2c80545, 32'hc2a659c7},
  {32'h44af384e, 32'h43617aa0, 32'hc2e5be30},
  {32'hc49db340, 32'hc1ed0578, 32'h439ba936},
  {32'h44f79e94, 32'h42ffa48a, 32'h43b11391},
  {32'hc3861650, 32'hc28044ac, 32'hc34e1076},
  {32'h44c5cfd2, 32'hc31c2ee4, 32'hc3cb865d},
  {32'hc4a19786, 32'hc3e14a51, 32'h43175e57},
  {32'h4517e3d1, 32'hc32828c9, 32'h435aa463},
  {32'hc4fc568a, 32'hc3130789, 32'hc3d0f29c},
  {32'h43fba38e, 32'h443402e4, 32'hc249686d},
  {32'hc527d4dd, 32'h43465cb6, 32'h4336bd8e},
  {32'h4379b370, 32'h441fcce9, 32'h4325eebf},
  {32'hc389cd20, 32'hc32c0ffe, 32'hc0be1eb0},
  {32'h43f805c8, 32'h43073071, 32'h422df7cc},
  {32'hc4d4a36c, 32'hc3d00dad, 32'hc388fc1a},
  {32'h44269ea4, 32'hc38c7d51, 32'hc1eb8eae},
  {32'hc50ed666, 32'h434d90b8, 32'h438da761},
  {32'h44fc2108, 32'h42a9f76c, 32'hc35c25a0},
  {32'hc48385fc, 32'hc39bf87f, 32'h43857767},
  {32'h4400284a, 32'hc36c3d1a, 32'hc290b792},
  {32'hc36a7a70, 32'h42e31d5c, 32'hc34a9f20},
  {32'h44ffc896, 32'h439b5e21, 32'h4279ebb7},
  {32'hc4f5d54d, 32'hc2f80faa, 32'h43f3208a},
  {32'h44c77f14, 32'hc3c0bef2, 32'h42af9b58},
  {32'hc3a40156, 32'hc3ce9a72, 32'h43a50ddc},
  {32'h43abc6ea, 32'h43a2ec06, 32'h43bdefe0},
  {32'hc5198e72, 32'h4308d0b4, 32'h43c2f724},
  {32'h4405814f, 32'h40ef0837, 32'hc398b832},
  {32'hc4e5363d, 32'h43043a75, 32'hc42612c1},
  {32'h447531f6, 32'hc35ddfd2, 32'h434448e3},
  {32'hc4ec5eae, 32'h4249f887, 32'hc3384d2b},
  {32'h44eed5e4, 32'h42868dec, 32'hc3801c1e},
  {32'hc4d3b3ce, 32'hc395a924, 32'h43e23f76},
  {32'h44332be0, 32'hc3b16136, 32'hc3a10f25},
  {32'hc4f30a11, 32'h4228fc31, 32'hc1e227ae},
  {32'h44f68b95, 32'h43f2f6b1, 32'h42375e71},
  {32'hc4fb8d8a, 32'h410ef599, 32'hc2bc665f},
  {32'h44efa654, 32'h4386e158, 32'hc3896a52},
  {32'hc4d350dc, 32'hc3da4f92, 32'h43e45f36},
  {32'h430bdb20, 32'h42f65175, 32'h3f8506a9},
  {32'hc50a2712, 32'hc234e299, 32'hc2dd158c},
  {32'h44e84151, 32'h438f6281, 32'hc187aa4d},
  {32'hc42a4a50, 32'hc2f498b2, 32'hc10ebe69},
  {32'h44ab00be, 32'hc25f5c60, 32'hc2da8beb},
  {32'hc3e15500, 32'h43213669, 32'hc30484c6},
  {32'h43a5e1a8, 32'h40aae1c8, 32'hc3822f6a},
  {32'hc4a6ac3f, 32'hc34250e0, 32'h42e3f746},
  {32'h44300f68, 32'hc2bdd082, 32'h421f9e33},
  {32'hc4be7849, 32'h4344eba1, 32'h43ad1d3e},
  {32'h450604aa, 32'hbf52c400, 32'hc2e4d1b9},
  {32'hc4ed49a2, 32'hc356a8e4, 32'hc30137e1},
  {32'h45069b85, 32'hc3e92f82, 32'hc37cb8f8},
  {32'hc45e3572, 32'h4326fdbc, 32'h440da213},
  {32'h449bf978, 32'h430dc50f, 32'hc2b610d5},
  {32'hc4b493fd, 32'hc357cc4a, 32'h43a10f78},
  {32'h440c1b20, 32'hc29a2f6c, 32'hc2dbf2b3},
  {32'hc492b930, 32'h43a368fb, 32'h436fdf04},
  {32'h44647387, 32'hc3fa4694, 32'h43863a79},
  {32'hc4400f67, 32'h434ca924, 32'h40ee0550},
  {32'h43a2c5ba, 32'h43ae87b2, 32'hc0bfa476},
  {32'h446b4046, 32'hc352824e, 32'h43a9bae5},
  {32'hc4d5a52f, 32'h4398fd33, 32'h43866985},
  {32'h421949f0, 32'hc3db85ab, 32'h42adfdee},
  {32'hc35da4a7, 32'h40b51e07, 32'h42edc64e},
  {32'h4481987e, 32'hc326f9da, 32'hc30bc208},
  {32'hc3ae62b4, 32'h415c1c92, 32'hc372a90e},
  {32'h4429fe32, 32'hc247e747, 32'hc42cd43e},
  {32'hc4f22805, 32'h430c1052, 32'hc384cd54},
  {32'h44311a28, 32'h429b3069, 32'h42fef240},
  {32'hc3c6ba60, 32'hc04ea860, 32'h42d05543},
  {32'h44e73e60, 32'hbff40cdc, 32'h4222eca5},
  {32'hc44fa6d0, 32'h43014891, 32'h43a2bef6},
  {32'h441bae38, 32'h43874c38, 32'hc399ee94},
  {32'hc4aff10f, 32'h42ccc524, 32'hc313c60b},
  {32'h44b01588, 32'h436eb3e9, 32'h416af5cc},
  {32'hc506c801, 32'h432ebfe1, 32'hc1df99cf},
  {32'h4513d8da, 32'hc347069a, 32'h436289d2},
  {32'hc50ff286, 32'hc2a07bbc, 32'h4213bf65},
  {32'h4420cb5e, 32'h431a0b98, 32'h42413d53},
  {32'hc405b8ac, 32'hc338372e, 32'h406c6ec0},
  {32'h4504db75, 32'hc3abd783, 32'hc2c1bae0},
  {32'hc4de4a68, 32'hc201adce, 32'hc25b915f},
  {32'h44babb18, 32'hc299db05, 32'hc2ebe852},
  {32'hc4a7f7b6, 32'h4383d634, 32'h42824fbe},
  {32'h4432427c, 32'hc2976d62, 32'hc3d6218b},
  {32'hc48adf16, 32'h41fccc34, 32'h4399d347},
  {32'h44fd13c6, 32'hc31761cd, 32'hc251bae7},
  {32'hc41382ba, 32'h43bcac46, 32'h42e95e87},
  {32'h44f7a411, 32'hc3420663, 32'h42303e5c},
  {32'hc46d3cb5, 32'hc347a0a0, 32'h43a359f8},
  {32'h4466e963, 32'hc26319a2, 32'h4382c96a},
  {32'hc44e91b4, 32'hc19720a7, 32'hc0449e0c},
  {32'h43075250, 32'hc3d1d01a, 32'h414c086e},
  {32'hc491f782, 32'hc3467f2a, 32'h4408816b},
  {32'h441e162f, 32'hc2eaffd4, 32'hc338e926},
  {32'hc43bed5c, 32'hc3521533, 32'h4254b33a},
  {32'h44c39da9, 32'hc3341146, 32'hc385e659},
  {32'hc4ebcac8, 32'h43897d0a, 32'hc272cd1e},
  {32'h450e5085, 32'hc2d7bdba, 32'h43d9b414},
  {32'hc40ee814, 32'h434fbdeb, 32'hc2c9b5f3},
  {32'h44b5ba97, 32'hc4090d74, 32'h431efc88},
  {32'hc50420a8, 32'hc114f242, 32'hc2cb47be},
  {32'h45063535, 32'hc3bb6f9f, 32'h42151d05},
  {32'hc4f4ae53, 32'h43747201, 32'hc2e10a63},
  {32'h43716820, 32'hc3795fb1, 32'h42987acc},
  {32'hc4b36958, 32'hc399aa1f, 32'hc38a0590},
  {32'h44881100, 32'hc3644515, 32'hc3aa5aa3},
  {32'hc4574cc4, 32'h432dc19d, 32'h43280431},
  {32'h44e004c9, 32'hc0eab598, 32'h43452d27},
  {32'hc41b0ab0, 32'hc2be7d9d, 32'h436b5324},
  {32'h44ec54d2, 32'h43dac280, 32'h40d968f4},
  {32'hc4faedb7, 32'hc399e6c2, 32'hc36b1796},
  {32'h44e19786, 32'hc25d21d8, 32'h43761960},
  {32'hc459354d, 32'hc08ed431, 32'h4369bd04},
  {32'h450f9d60, 32'h435a67d3, 32'h4309278c},
  {32'hc3b70668, 32'hc22c6d22, 32'hc381af59},
  {32'h443e2076, 32'h439524fd, 32'hc2ef8cd4},
  {32'hc3982883, 32'hc3899134, 32'hc3c0b426},
  {32'h44e4aedd, 32'h439f48c2, 32'hc318d74d},
  {32'hc430dbba, 32'hc3c9e18c, 32'h41eb6437},
  {32'h438a1aa8, 32'hc4505cee, 32'hc2881f23},
  {32'hc3966bec, 32'h43a4bec6, 32'hc393e109},
  {32'h44e0f707, 32'hc37c5b04, 32'h43a98851},
  {32'hc42ac15c, 32'h4280701e, 32'h4063880a},
  {32'h4504b165, 32'hc301a306, 32'h434736e1},
  {32'hc46ab920, 32'hc0d1d1b7, 32'h41df2107},
  {32'h43eaf628, 32'h41e19aba, 32'hc38cea23},
  {32'hc4c32f37, 32'hc3b95516, 32'hc3c93d38},
  {32'h44ba3951, 32'h4391926d, 32'h440e590d},
  {32'hc48f1237, 32'h4306ce68, 32'hc284e479},
  {32'h44de0a76, 32'h42d716d8, 32'hc23b23c2},
  {32'hc490574c, 32'h429db033, 32'hc32f23c9},
  {32'h44811224, 32'h437a100a, 32'h4216a4fa},
  {32'hc4ed66cc, 32'hc141aba1, 32'h436dd188},
  {32'h438ca599, 32'hc3bdadcd, 32'hc2f4576c},
  {32'hc4fd2a96, 32'hc31f5863, 32'h4331d4d3},
  {32'h44671d98, 32'h438cb469, 32'hc211b117},
  {32'hc4ddceda, 32'hc2038ed3, 32'h41a23db4},
  {32'h44e4d2de, 32'h42120aea, 32'hc2dcfa67},
  {32'hc4047f23, 32'hc2da66a3, 32'h434cd351},
  {32'h44177c3b, 32'h42c68238, 32'h42cc0b37},
  {32'hc509a40a, 32'hc3179cfe, 32'hc384999e},
  {32'h44b12076, 32'h40c286cf, 32'h431b08b9},
  {32'hc49d6ab6, 32'h412994fe, 32'hc2dce010},
  {32'h4464e1cd, 32'hc3b1231c, 32'hc2887a68},
  {32'hc438f3d8, 32'h42c2c574, 32'h42c6f379},
  {32'h44581642, 32'hc36b488d, 32'hc33b7163},
  {32'hc49dae06, 32'hc28c86c6, 32'hc3143843},
  {32'h44d46021, 32'hc3d0ec10, 32'hc3916e49},
  {32'hc492c793, 32'hc2288e2c, 32'hc31c3536},
  {32'h44f50754, 32'hc37ff49e, 32'hc33f8235},
  {32'hc4b1c712, 32'h43b6a6be, 32'hc28baa7f},
  {32'h44efb23d, 32'hc3773d8e, 32'h437695b7},
  {32'hc3fbaabc, 32'hc38db185, 32'hc38ed7a4},
  {32'h44d055c2, 32'h4319f391, 32'h43c4cd64},
  {32'hc507c705, 32'hc3b50827, 32'h41793eb2},
  {32'h44c27ac6, 32'h430afb29, 32'hc2ae3961},
  {32'hc3e83904, 32'h43a934d4, 32'hc3531726},
  {32'h44ba34e5, 32'h41ee1686, 32'hc3bf4c17},
  {32'hc496535e, 32'h4380e0e8, 32'h41399a94},
  {32'h44e74b38, 32'h4396663e, 32'h439e0188},
  {32'hc4e8ac9b, 32'h441b6a8a, 32'h43612a6b},
  {32'h43146920, 32'h42b8e185, 32'h4310034d},
  {32'hc3476b8d, 32'h42bc581b, 32'h43c33fb7},
  {32'h43d0722c, 32'h42e95008, 32'h436a6f16},
  {32'hc45f8734, 32'hc3949391, 32'hc34a70dc},
  {32'h44a744f0, 32'hc31e78b6, 32'hc3443f8f},
  {32'hc4012126, 32'h433b9a1d, 32'hc1c75350},
  {32'h44b2ce12, 32'hc34aac02, 32'h42443fd7},
  {32'hc4908cf2, 32'h439155b0, 32'h4350e5be},
  {32'h44bf6c6b, 32'hc1fbeb7d, 32'hc2709360},
  {32'hc3397056, 32'hc368a61f, 32'h43a36d99},
  {32'h441e0d63, 32'hc3620616, 32'hc33fb425},
  {32'hc519d3b1, 32'hc1bfa7e9, 32'h42565359},
  {32'h44d9a04b, 32'h4385c9be, 32'h429a4ff7},
  {32'hc3d3997c, 32'h4389fdb3, 32'hc2585006},
  {32'h450e3f8e, 32'hc15744ac, 32'h436f9fa1},
  {32'hc5010ffc, 32'h43fe0840, 32'h434387f9},
  {32'h44988f04, 32'h41809c30, 32'hc2186574},
  {32'hc4da04cd, 32'hc309971f, 32'hc2ee31ab},
  {32'h41bdf4e0, 32'h440c1d5b, 32'h4103f4b6},
  {32'hc4cf6e7a, 32'hc278fe22, 32'h4408cd8f},
  {32'h44d1b944, 32'h43d90d43, 32'h433d8fe2},
  {32'hc48e0402, 32'hc212797e, 32'hc2c03aea},
  {32'h441731b2, 32'hc349a27a, 32'hc334df4f},
  {32'hc4ed921c, 32'h422892e2, 32'hc2b1b823},
  {32'h4495dcc1, 32'h42bd7a75, 32'h41ebcf0c},
  {32'hc3aa7180, 32'hc1d78fbe, 32'hc310cf4b},
  {32'h4529179c, 32'hc2e09626, 32'hc2e4c972},
  {32'hc509d10f, 32'h43364882, 32'h4403b1df},
  {32'h429881f0, 32'h43941cee, 32'h4209ea6d},
  {32'hc3f319cc, 32'hc2213a22, 32'h42ac24ff},
  {32'h44ec6241, 32'h42ee38f0, 32'h435bec59},
  {32'hc15a0a27, 32'h4251619a, 32'h42a1e78f},
  {32'h44f79822, 32'h3ffb7460, 32'h42d5de3a},
  {32'hc4f94e09, 32'h432b6677, 32'hc2bb7936},
  {32'h4442fefe, 32'hc392104d, 32'hc3facd74},
  {32'hc487ebe4, 32'hc2d61bac, 32'hc1c6c3f2},
  {32'h44e048c0, 32'hc3757d2a, 32'h43104d56},
  {32'hc4c667be, 32'hc3098bad, 32'h43a8f1fb},
  {32'h449119bf, 32'hc0dd23ec, 32'hc306bbfb},
  {32'hc4846d89, 32'hc34e486a, 32'h432b6465},
  {32'h45056a89, 32'hc360be70, 32'hc38a9274},
  {32'hc432f18d, 32'hc31f3a48, 32'h445a218a},
  {32'h44a5b315, 32'hc166a20a, 32'h42a0e158},
  {32'hc4e58973, 32'hc24e9f84, 32'h42265347},
  {32'h44d92e61, 32'h430e6a4c, 32'hc2f99166},
  {32'hc4bd9400, 32'hc17603d1, 32'h43865454},
  {32'h44de6865, 32'h43ef14eb, 32'hc3598026},
  {32'hc48130b2, 32'h43a878b0, 32'h430e4c41},
  {32'h445e77c1, 32'hc243a644, 32'hc3000f67},
  {32'hc4dbbef2, 32'h430244b0, 32'h425c765d},
  {32'h450d35a3, 32'hc2f567de, 32'h3fec0850},
  {32'hc44c3b88, 32'h431cde43, 32'h42891a42},
  {32'h43098048, 32'hc297fc08, 32'h429ce4cb},
  {32'hc4c84f15, 32'h439ec232, 32'hc3aeb02b},
  {32'h446c94e2, 32'h424cb4da, 32'h428ea484},
  {32'hc464ef2e, 32'h4414e387, 32'hc33a85bf},
  {32'h4500fcb1, 32'hc386d118, 32'h4313a8ec},
  {32'hc4a76a93, 32'hc3d25177, 32'h438bf76f},
  {32'h444e6a79, 32'h43a4508c, 32'h413b7a18},
  {32'hc4da741c, 32'hc3477a81, 32'hc3944c0f},
  {32'h43dc4558, 32'hc2947b75, 32'hc2745ccb},
  {32'hc4b84284, 32'hc2bd5edb, 32'hc0f2b0f0},
  {32'h449ac89c, 32'hc30de6fc, 32'hc3bab1bb},
  {32'hc46451e2, 32'hc2a0fefc, 32'hc34a64b9},
  {32'h44f83b4e, 32'h43afdc9f, 32'hc1e4e43c},
  {32'hc40a5a78, 32'h40ddbc39, 32'hc252ee9a},
  {32'h44714880, 32'hc3882b7b, 32'hc2575ebc},
  {32'hc4083df4, 32'hc37ba24b, 32'h4396ffe7},
  {32'h44ec0d34, 32'hc3108708, 32'h429b4c97},
  {32'hc4a02bb4, 32'hc38280ba, 32'h43ae0086},
  {32'h44e71b04, 32'hc2b281aa, 32'h43a93f65},
  {32'hc44066de, 32'h43527cd4, 32'hc30f2220},
  {32'h45175942, 32'h439ce0fd, 32'hc2190292},
  {32'hc4d4961c, 32'hc2de73ed, 32'h431da914},
  {32'h44fcdb30, 32'hbfc49b6a, 32'h42dad519},
  {32'hc45bc3b2, 32'hc3397017, 32'h429f70ef},
  {32'h436ff6c4, 32'hc2ab512c, 32'hc1ad2cd4},
  {32'hc4d0a1af, 32'hc39914b4, 32'hc0e68b8c},
  {32'h44d53a5e, 32'h41b48eb0, 32'h41af7622},
  {32'hc4169963, 32'h425f9615, 32'hc39fe444},
  {32'h44a3c77d, 32'hc2f22ad2, 32'h42bc0110},
  {32'hc4bb331f, 32'hc3143518, 32'hc2993015},
  {32'h44867d31, 32'hc317f11c, 32'h418052ea},
  {32'hc44e7e32, 32'hc2b32488, 32'h42969ad5},
  {32'h42c0ab34, 32'hc347bdbe, 32'hc2e32895},
  {32'hc4deb983, 32'hc15edd4c, 32'h4299bef8},
  {32'h43e6305c, 32'hc25ed40e, 32'h420ad6ea},
  {32'hc5126d09, 32'h43003404, 32'h433709f4},
  {32'h442fd4c6, 32'h43890fc3, 32'hc2fbce47},
  {32'hc41b6f82, 32'h42ad88c2, 32'h4090031e},
  {32'h450abd7e, 32'hc2196303, 32'h4311ad4d},
  {32'hc4827aac, 32'hc3be1225, 32'h424c052a},
  {32'h4491b591, 32'hc38b6958, 32'h4303f446},
  {32'hc4d878b8, 32'h434a9f51, 32'h439a47c3},
  {32'h4184c260, 32'h41a17802, 32'hc383bc70},
  {32'hc44416d0, 32'hc2e387bc, 32'hc31fb1db},
  {32'h44aea962, 32'h433ed13b, 32'hc288f647},
  {32'hc3e7eb40, 32'hc3a2af3a, 32'hc2d84efc},
  {32'h444b7945, 32'hc38262b6, 32'hc236d772},
  {32'hc3116d60, 32'h435e9542, 32'h432b2818},
  {32'h44f7cd54, 32'hc344f685, 32'hc2bf1271},
  {32'hc43bc870, 32'h4353ff33, 32'hc2ebd067},
  {32'h443fe3ac, 32'hc3b2930a, 32'h441ea476},
  {32'hc508b309, 32'h41950694, 32'h4322b126},
  {32'h44ffc849, 32'h4311ccbc, 32'hc012d200},
  {32'hc42be4f9, 32'hc1da7714, 32'hc2cf32d5},
  {32'h4456991c, 32'hc15d5990, 32'h4376d35f},
  {32'hc31b7160, 32'hc39cafbf, 32'h41009269},
  {32'h44a8347d, 32'hc3054a69, 32'hc143ae02},
  {32'hc3e88902, 32'hc0e8cb4e, 32'h40309b39},
  {32'h4374d92c, 32'h43fa6f33, 32'h3fb5de69},
  {32'hc3d43570, 32'h41d1de03, 32'h42dd7c9f},
  {32'h448087ac, 32'h41e93a6f, 32'hc2d6997b},
  {32'hc46bdb66, 32'h4331377c, 32'h42000098},
  {32'h44471c90, 32'hc323b4cd, 32'hc321697d},
  {32'hc3d22d6d, 32'h430e517e, 32'h41cdca6c},
  {32'h44c91214, 32'h435895a6, 32'h434e1c8a},
  {32'hc34aae60, 32'h41a88103, 32'h432c87e2},
  {32'h44aeaeaf, 32'hc39bf056, 32'hc2c53b81},
  {32'h42fcdae7, 32'h436376cf, 32'hc28218ae},
  {32'h44494294, 32'hc3229f65, 32'h43f2d062},
  {32'hc4968a5f, 32'hbf2213f4, 32'hc32f6576},
  {32'h4342beae, 32'hc3286e88, 32'h42d9333c},
  {32'hc52293d9, 32'h4389ef33, 32'hc27cc0cc},
  {32'h44c44b19, 32'h43e87aa2, 32'h42d8cdd4},
  {32'hc4fc0cd0, 32'hc2810a4f, 32'h42ccae5e},
  {32'h436d4e36, 32'hc2bc477c, 32'hc313a3ab},
  {32'hc38e8288, 32'h43d0fa00, 32'hc3a65eb8},
  {32'hc325f124, 32'h430a332b, 32'h41b84dda},
  {32'hc331c40d, 32'h432c4642, 32'hc32cc8bb},
  {32'h44af97e3, 32'hc2269010, 32'hc195b37e},
  {32'hc4b429dc, 32'h41c8402b, 32'h4381e1a6},
  {32'h43a44e0e, 32'h43843421, 32'hc3a0a370},
  {32'hc4412ad6, 32'hc33299fc, 32'hc3817b67},
  {32'h44dc801c, 32'hc38a4dfa, 32'hc303e1ee},
  {32'hc4cc77be, 32'hc35e31dc, 32'hc3a5feeb},
  {32'h44964706, 32'hc2502584, 32'h439b3a11},
  {32'hc4e07a13, 32'hc3562492, 32'hc3c2327a},
  {32'h44d40ea7, 32'hc2a734ec, 32'hc3957a88},
  {32'hc507a585, 32'hc2fcb3e2, 32'hc26bf5dc},
  {32'h450b2083, 32'hc23e75d8, 32'hc30080d6},
  {32'hc5043277, 32'h434ee067, 32'h4331a538},
  {32'h4361fd94, 32'h43634412, 32'h432ba5f3},
  {32'h43417c30, 32'h42ce1c74, 32'hc2068e70},
  {32'h44e8892c, 32'h432d385c, 32'hc32fe81f},
  {32'hc3a1e0ae, 32'h428a5296, 32'hc384f2e3},
  {32'h448233cf, 32'h43dfe524, 32'h41d6206a},
  {32'hc3957dd8, 32'hc1a19a62, 32'hc45341b9},
  {32'h44a06d05, 32'h43a12c4e, 32'hc319a454},
  {32'hc42d55f8, 32'h437bf750, 32'h4387a312},
  {32'h44b2182d, 32'hc2414942, 32'h43bbdc29},
  {32'hc42e6482, 32'h41f764e5, 32'hc2a86c8d},
  {32'h44523fdc, 32'hc2e33900, 32'h42e2bb48},
  {32'hc4be2f1b, 32'h428cef1c, 32'hc323675b},
  {32'h448ba810, 32'hc32f4787, 32'hc38831c8},
  {32'hc4b0fa9a, 32'hc28a5e12, 32'h42a0c05d},
  {32'h449c6dce, 32'hc0d42ebe, 32'hc24f5b66},
  {32'hc3a35d08, 32'h431c0bc0, 32'h42ba7224},
  {32'h45074eb6, 32'hc30069e3, 32'h42d5d5c5},
  {32'hc4ae2f06, 32'hc387de03, 32'hc31373a2},
  {32'h4510208f, 32'hc3960084, 32'hc2de4e10},
  {32'hc4ed118c, 32'hc400bef0, 32'h42a8c924},
  {32'h4471a6b0, 32'h4312b734, 32'h417a5820},
  {32'hc4048fb5, 32'h433b3a2a, 32'hc36a23f3},
  {32'h44e2aad5, 32'h42f1312d, 32'hc2f6d256},
  {32'hc48ef8c6, 32'h4355998e, 32'h4216baae},
  {32'h44866e64, 32'hc2fbc65e, 32'h42a7500c},
  {32'hc49a3e22, 32'h40b31f13, 32'h42f51531},
  {32'h44cae7cc, 32'h4268b99e, 32'hc206a913},
  {32'hc3082780, 32'h42504e5e, 32'hc2b2ec5a},
  {32'h4402f222, 32'h41ac1e81, 32'hc26bd874},
  {32'hc5184710, 32'hc13f2605, 32'h43259133},
  {32'h44b544a0, 32'hc3b4e254, 32'h43228ff5},
  {32'hc4e0c032, 32'hc35a1c38, 32'h438c99fc},
  {32'h45070f60, 32'hc34fff2f, 32'hc2e44252},
  {32'hc4b4ad78, 32'hc28b908c, 32'h431bd2ca},
  {32'h44b3f314, 32'hc3a4656b, 32'hc393f1a6},
  {32'hc4b57362, 32'h439c471a, 32'hc38ffbd5},
  {32'h443f117c, 32'h42f5b3b0, 32'h4343eea7},
  {32'h42212440, 32'h419362ca, 32'h42bfb4e0},
  {32'h44c14b71, 32'h4323f0f7, 32'h43548dd2},
  {32'hc4c49af4, 32'hc3a63ad4, 32'h441021df},
  {32'h4420f702, 32'h41e979a8, 32'hc39e4d21},
  {32'hc45a1c52, 32'hc2b82a3b, 32'h43e060e5},
  {32'h450cfc6b, 32'h434b97a2, 32'h42ddfe91},
  {32'hc4b7b808, 32'h4340f803, 32'hc2aef3d1},
  {32'h44dd9b2c, 32'hc3e47b51, 32'hc2639241},
  {32'hc47ddbfe, 32'h4169c995, 32'hc25c3c05},
  {32'h45177a09, 32'hc364468d, 32'h43b53d4a},
  {32'hc4aae782, 32'h423555b3, 32'hc2d06939},
  {32'h443ba504, 32'h428ad72e, 32'hc2e80ccd},
  {32'hc436caee, 32'hc2b9ce24, 32'hc170e8dd},
  {32'h44854d24, 32'hc35d94f0, 32'hc30c1350},
  {32'hc22df740, 32'h408d05d0, 32'hc2998c8d},
  {32'h44a32e75, 32'hc338b477, 32'h4398da97},
  {32'hc50396e9, 32'h42fdda67, 32'h439711ec},
  {32'h45066b76, 32'h43b3cb89, 32'h412a645f},
  {32'hc365a7c0, 32'h43395f19, 32'h42b7ced7},
  {32'h44e967cb, 32'h440dcfcc, 32'hc2d22001},
  {32'hc4df94a3, 32'hc3a1eecf, 32'h4387f4cc},
  {32'h446368f4, 32'hc3e5da9f, 32'h427f1aaf},
  {32'hc408d911, 32'h4398d842, 32'h41ab4044},
  {32'h44ee9a1e, 32'h41f7856e, 32'hc31380fe},
  {32'hc3309930, 32'hc2a296fb, 32'hc2d89920},
  {32'h440322ea, 32'hc331bf6e, 32'hc374c2d6},
  {32'hc41affa0, 32'h43464ebe, 32'hc0fd754c},
  {32'h429daf90, 32'hc2e360f2, 32'h409e2398},
  {32'hc4fa7420, 32'h4397cb33, 32'h4332c6ee},
  {32'h451a823f, 32'h4315dc6d, 32'h43029c51},
  {32'hc480e3d2, 32'h43447d91, 32'h43074962},
  {32'h44ecb31c, 32'h409b1c68, 32'hc3b2f7a2},
  {32'hc48dd0c8, 32'hc3825963, 32'h42bf3e4c},
  {32'h446b899e, 32'hc2106850, 32'h4207a999},
  {32'hc491a32d, 32'h407060f2, 32'h43232cd8},
  {32'h43a0a596, 32'hc3767ca3, 32'hc3b4e834},
  {32'hc484b9d6, 32'h426b2735, 32'h43ad1222},
  {32'h44bfb8ce, 32'hc3c3de6e, 32'h42e863ba},
  {32'hc3a0bffa, 32'hc28fb150, 32'hc3cdf969},
  {32'h45049363, 32'hc2fbc618, 32'hc45a2851},
  {32'hc4dab462, 32'hc2872989, 32'h42b1246d},
  {32'h44bc0019, 32'h421ac8c5, 32'h42c3feb6},
  {32'hc45706b4, 32'hc1e0df7d, 32'hc2bc1414},
  {32'h438d7b0b, 32'h43021e19, 32'hc2ed145c},
  {32'hc4f7d634, 32'hc2bb0a8f, 32'h42aa0cce},
  {32'h4502a031, 32'h431d30be, 32'h4408986e},
  {32'hc454e754, 32'hc29e2974, 32'h42f29d6a},
  {32'h449cdb24, 32'hc2508fe8, 32'hc3192133},
  {32'hc4e0ea1b, 32'h416fa9ec, 32'h428b109b},
  {32'h44faa0f5, 32'hc38ae634, 32'hc325bce4},
  {32'hc4479d6f, 32'h432f1163, 32'h4323ca8b},
  {32'h446114e4, 32'hc2421984, 32'hc38db018},
  {32'hc5089277, 32'h4344b379, 32'hc39a4618},
  {32'h4509fd02, 32'hc3419cda, 32'hc14bdc5f},
  {32'hc44fd302, 32'hc3573ed5, 32'h43a0d882},
  {32'h448ded69, 32'h438b24f0, 32'h43178b69},
  {32'hc4411eb4, 32'hc3638348, 32'hc26963eb},
  {32'h451fe94c, 32'hc038bdee, 32'hc039f56c},
  {32'hc460cc3c, 32'h42aad362, 32'hc23c29fc},
  {32'h4465d384, 32'h42d0b52d, 32'h43ba7967},
  {32'hc509d771, 32'h440713a3, 32'hc30926b5},
  {32'h42c39968, 32'h42e59648, 32'hc13292dc},
  {32'hc4f97588, 32'h43321e1a, 32'hc28faf06},
  {32'h4377b224, 32'h43662a60, 32'h4293190c},
  {32'hc502cdc1, 32'h422d07d1, 32'hc258bad1},
  {32'h44f3909b, 32'h43cf1532, 32'h4349a6c3},
  {32'hc46123f4, 32'h43f32577, 32'h42977f16},
  {32'h44b7f87d, 32'hc35646a0, 32'hc39c57eb},
  {32'hc39a5a16, 32'h429f47f1, 32'h4101f2f9},
  {32'h44e9a343, 32'hc03990ec, 32'hc34f3220},
  {32'hc5055932, 32'hc2d5e3f3, 32'hc1763ac4},
  {32'h44b26ea5, 32'h43128ca8, 32'h43e87bad},
  {32'hc44af082, 32'h432d93c1, 32'h42eb4454},
  {32'h44b785d8, 32'hc3b47e20, 32'h43b1be59},
  {32'hc4c7b2b2, 32'h43638e56, 32'h42847109},
  {32'h451d0679, 32'h437592dd, 32'hc3bb9616},
  {32'hc4448104, 32'h439861ef, 32'hc3263c71},
  {32'h45105bc1, 32'hc3946c9d, 32'h436ba44b},
  {32'hc484af63, 32'hc336dfdd, 32'h43328815},
  {32'h44bf54c4, 32'h4306634f, 32'h434c44ab},
  {32'hc4c45a51, 32'h420fb7e2, 32'hc290fdab},
  {32'h44127f3c, 32'hc33d65d2, 32'hc40183cf},
  {32'hc45a01c5, 32'h43063f66, 32'h42d8c8fd},
  {32'h44107328, 32'h42f44f8c, 32'h439e7bef},
  {32'hc50041b5, 32'h4387f8b1, 32'h42eed152},
  {32'h450b84c3, 32'hc3343315, 32'hc2537fe9},
  {32'hc471ef64, 32'h439d6e42, 32'hc38a023f},
  {32'h44c75370, 32'h42078b27, 32'h442c7375},
  {32'hc4c34117, 32'h4386b88d, 32'h4313a210},
  {32'h446a3d00, 32'h43f0ca28, 32'hc350ac9a},
  {32'hc3fe4ba0, 32'hc1973764, 32'hc24bd3f7},
  {32'h44342b5c, 32'hc334f1ff, 32'hc400c546},
  {32'hc42bf443, 32'hc3a47cfe, 32'h42f23a9e},
  {32'h448a6425, 32'h42741410, 32'hc39f7213},
  {32'hc500fce7, 32'h437b4cdf, 32'hc3c9b94c},
  {32'h44962020, 32'hc301e03c, 32'h42c17d08},
  {32'hc50f601e, 32'hc17ea593, 32'hc31465b6},
  {32'h4482676a, 32'hc306b444, 32'h4346daff},
  {32'hc40204a9, 32'hc3a4fd69, 32'hc1de270c},
  {32'h44c8a5e0, 32'h43510a9e, 32'h40f59ea9},
  {32'hc4731dfb, 32'h4307102b, 32'h42f4248d},
  {32'h447c7dfb, 32'h40a8d745, 32'h439ae299},
  {32'hc48d27a6, 32'hc3b876e7, 32'h43a3a7b9},
  {32'h44c7a006, 32'hc197580e, 32'hc23ae35b},
  {32'hc4d99c84, 32'hc2243467, 32'hc33388d7},
  {32'h4517ebd8, 32'hc3c267cd, 32'hc323c5c7},
  {32'hc4b100c9, 32'h42ee6263, 32'h43454e49},
  {32'h44c137b4, 32'h42ab8875, 32'hc401b552},
  {32'hc416364d, 32'h42cc5293, 32'hc3b21f3c},
  {32'h43e5db08, 32'h433b1a2e, 32'h4375f428},
  {32'hc5142b84, 32'hc2df3533, 32'h437a51d6},
  {32'h441511ce, 32'hc2215d0c, 32'hc2b4a917},
  {32'hc3f3c2d9, 32'hc2d78163, 32'hc347d7a0},
  {32'h445b12c9, 32'hc2a3c24a, 32'h41b86fa9},
  {32'hc4a542ab, 32'hc314e7e4, 32'hc257ec97},
  {32'h4486f507, 32'h42ef094a, 32'h42d3743d},
  {32'hc4e54530, 32'h43061450, 32'hc3219692},
  {32'h407162c0, 32'hc3e8842f, 32'h432b02ed},
  {32'hc4bb390a, 32'h43c6e730, 32'hc39b2a81},
  {32'h4470121d, 32'hc36611f8, 32'h419c3c5c},
  {32'hc4a9d774, 32'h44160493, 32'hc3635a8d},
  {32'h45034a86, 32'hc2e566e4, 32'h432510f1},
  {32'hc50c9b9c, 32'hc3182633, 32'h42cbba6f},
  {32'h44045a1e, 32'hc224cfbd, 32'hc3e07c18},
  {32'hc4efcd28, 32'h4389b595, 32'hc2fd8c69},
  {32'h44d56c0a, 32'hc21fd726, 32'h42c73270},
  {32'hc4ec8e21, 32'hc38e81e6, 32'h4364bb9f},
  {32'h4455bae1, 32'hbffc5682, 32'h43ce605d},
  {32'hc41b3cef, 32'h430eb036, 32'hc1818745},
  {32'h4319cc00, 32'h42a92893, 32'h426e1e6d},
  {32'hc42552ad, 32'h433d6108, 32'h43b7bbb3},
  {32'h44b44cc9, 32'h43ea4758, 32'h42388a1d},
  {32'hc38f19d0, 32'hc30292ac, 32'h430583a7},
  {32'h4509280d, 32'hc37fcadb, 32'h4285c248},
  {32'hc4fb9609, 32'hc2afd6f1, 32'h41240b95},
  {32'h448e7968, 32'hc36f280a, 32'h44110f99},
  {32'hc4287977, 32'hc31aa229, 32'h412502e2},
  {32'h445864ea, 32'hc2a0ec1c, 32'hc4045c21},
  {32'hc3b97b04, 32'h4441fe32, 32'hc2685362},
  {32'h44bd3301, 32'hc41a77e8, 32'h42db18cc},
  {32'hc43ff6bb, 32'h42a86ebb, 32'hc427be9a},
  {32'h44eb8891, 32'hc41cfbe6, 32'hc31a500b},
  {32'hc4852ffc, 32'hc2a14bb6, 32'hc2b4016c},
  {32'h4464e7c2, 32'hc331ee82, 32'hc2d88642},
  {32'hc43668b0, 32'h4374cd4d, 32'hc3832421},
  {32'h42ecd540, 32'hc0812356, 32'h43bb5434},
  {32'hc47739a5, 32'hc302dc19, 32'h427f7150},
  {32'h44d3ff43, 32'h42afb757, 32'h42d71e06},
  {32'hc4395300, 32'hc37998c5, 32'h4196bcd7},
  {32'h44b37ca0, 32'h4342cade, 32'hc2f52fa6},
  {32'hc4534fa4, 32'hc36ce5c5, 32'h432a6a54},
  {32'hc49614df, 32'h43117617, 32'hc3e8c1cf},
  {32'h45021c4c, 32'h421f7fbd, 32'h43bcbbdd},
  {32'hc35a790e, 32'hc3888e1a, 32'h42ef4de0},
  {32'h44f50646, 32'h4306a2f5, 32'h4336c463},
  {32'hc5039f2d, 32'hc2c7b746, 32'hc33bf2e0},
  {32'h44f32776, 32'hc3f7d930, 32'hc33ee79b},
  {32'hc4a30d29, 32'hc2dd9eec, 32'h41d21e05},
  {32'h44a9a76c, 32'h426864ff, 32'h42b0959a},
  {32'hc442c508, 32'h41db73f3, 32'h42900294},
  {32'h44282636, 32'h432b3c4b, 32'hc2508517},
  {32'hc4e980d3, 32'h43846438, 32'hc3a45b71},
  {32'h4508398f, 32'hc3198387, 32'h4330654b},
  {32'hc4a5c361, 32'hc2fa103f, 32'h42aecd1d},
  {32'h443b8284, 32'h4386509b, 32'h43a53ad2},
  {32'hc4235647, 32'hc28b3d97, 32'hc363a565},
  {32'h432387e8, 32'hc34dad76, 32'hc3e23ec8},
  {32'hc392a574, 32'h41fcb414, 32'hc41581ec},
  {32'h43743685, 32'hc0c75d64, 32'h43ad8b80},
  {32'hc4e25bba, 32'hbf22ee60, 32'hc2b6d648},
  {32'h44808403, 32'h42bfc7d3, 32'hc2984414},
  {32'hc45567a8, 32'hc2936ac6, 32'h4236dda5},
  {32'h43359688, 32'hc383bf88, 32'h43e0cf51},
  {32'hc4ffb23c, 32'hc2fccb49, 32'hc359459e},
  {32'h449e5d31, 32'h434dec13, 32'h436bd294},
  {32'hc4f461ae, 32'h41106618, 32'hc407a166},
  {32'h44ee518d, 32'hc2d95e59, 32'hc280398d},
  {32'hc4cca552, 32'h42f52d65, 32'hc31eb8c7},
  {32'h44ee3cae, 32'hc1a770e0, 32'h42b3a3a9},
  {32'hc43c3778, 32'h43d14112, 32'hc428442c},
  {32'h43b6ebc9, 32'h428386c7, 32'hc1da3a59},
  {32'hc40f8c5e, 32'hc0a43267, 32'hc2c6b2a4},
  {32'h441f1f6b, 32'h4283284c, 32'h43ad9a05},
  {32'hc4effb12, 32'hc403b176, 32'h43a41518},
  {32'h4512958e, 32'h42ae430f, 32'h441de398},
  {32'hc50afdeb, 32'hc2c9c9bd, 32'h4302eabb},
  {32'h431dd8a0, 32'hc3616179, 32'hc39de23f},
  {32'hc4e2fc04, 32'h42a85e49, 32'h43ea703c},
  {32'h44f3d266, 32'h43610d84, 32'hc27dfb76},
  {32'hc38f3f5e, 32'hc12cf8dd, 32'hc3bc1926},
  {32'h4515cb4f, 32'h433988d5, 32'h43c028d9},
  {32'hc491524d, 32'h43925a19, 32'h43930d05},
  {32'h44f52b6c, 32'hc2d3b2c6, 32'h43a8a8c2},
  {32'hc4d257d9, 32'hc1afb06b, 32'h43a647f6},
  {32'h444f12ba, 32'h42c045c6, 32'h43e9d7de},
  {32'hc528b293, 32'hc33df340, 32'h40114238},
  {32'h40c5c880, 32'h42b93be0, 32'hc3031e9f},
  {32'hc4f507e2, 32'h4322c2d5, 32'hc339df9e},
  {32'h44183a54, 32'h4333e1bc, 32'hc3128bfd},
  {32'hc5048de7, 32'h4371b013, 32'h4306323a},
  {32'h447c3c2c, 32'h43069287, 32'h4151cb72},
  {32'hc36b4939, 32'hc20a314c, 32'hc34964c8},
  {32'h433a72c0, 32'h43400236, 32'h41ba8da0},
  {32'hc40c9d8b, 32'h43c8fc21, 32'hc24ab032},
  {32'h44fafcd2, 32'h43d0c17a, 32'h433a0e56},
  {32'hc410889f, 32'h4343fb93, 32'hc3dfc78c},
  {32'h44b076ff, 32'hc3710d06, 32'hc31f0734},
  {32'h40693900, 32'h438c5021, 32'h4259b27d},
  {32'h44fda521, 32'h433c4be0, 32'hc3049e44},
  {32'hc4cd3518, 32'h437a6935, 32'hc3b8f309},
  {32'h441593c0, 32'h42332399, 32'hc343ee06},
  {32'hc4dc4f8c, 32'h42bb5506, 32'hc372bd19},
  {32'h44bab5ee, 32'hc3588c94, 32'h42f4dd58},
  {32'hc5069f9c, 32'h41ddcd40, 32'hc28da245},
  {32'h44c7a6cc, 32'hc4109d12, 32'hc1f7a3d8},
  {32'hc4cde106, 32'h42b32609, 32'hc2b9fc60},
  {32'h44ffee47, 32'h42f3b731, 32'h43421af7},
  {32'h437b0f9e, 32'h43a7e82e, 32'hc2c0a321},
  {32'h44e71b2f, 32'hc2c9a1c7, 32'h438e9a98},
  {32'hc4894969, 32'h437276f0, 32'hc1775b03},
  {32'h44fc679e, 32'hc2806d04, 32'h431e36cb},
  {32'h43221e0f, 32'h42a5d60e, 32'h440a4e06},
  {32'h4516e517, 32'hc3044091, 32'h43891fa8},
  {32'hc40765ce, 32'hc41a69ca, 32'hc32d8f4c},
  {32'h44883de3, 32'hc2d20341, 32'hc29c123b},
  {32'hc4b64194, 32'hc2498db6, 32'h431d3a84},
  {32'h450333a4, 32'h435fd004, 32'h4216343f},
  {32'hc4ba82b8, 32'h42a2adac, 32'h4341b6d2},
  {32'h42e90280, 32'h4391cd7e, 32'hc30ef08e},
  {32'hc40ba908, 32'h4357d7fb, 32'h42d072ec},
  {32'h44bf4777, 32'hc3a6faf8, 32'h443b23d4},
  {32'hc49124a4, 32'hc3ab680b, 32'h43bd2cdc},
  {32'h4437d673, 32'hc4094e28, 32'h4322f9c6},
  {32'hc4dab726, 32'hc313bd8a, 32'h4330007b},
  {32'h431d3528, 32'h435978b4, 32'hc2bdcbe3},
  {32'hc430a836, 32'h424a8109, 32'hc3137de1},
  {32'h45144927, 32'h413d5e7d, 32'h4317c919},
  {32'hc46fbe9b, 32'hc31fcc75, 32'h437d6945},
  {32'h445835e6, 32'h42655f7a, 32'h43a3a510},
  {32'hc4a84236, 32'h43f6943e, 32'h422005b6},
  {32'h451782be, 32'hc3db5c59, 32'h43546674},
  {32'hc40dedd8, 32'h42c896a7, 32'h41e21a59},
  {32'h441ba0a1, 32'hc289b9dd, 32'h42adb477},
  {32'hc48aef15, 32'hc0c76ac2, 32'hc1bb80c8},
  {32'h44557198, 32'h42eb7735, 32'h42defaba},
  {32'hc3e21482, 32'hc41a9088, 32'h41a82519},
  {32'h432c8c90, 32'h4294218f, 32'hc30c90a5},
  {32'hc4dde2f2, 32'h438b024a, 32'h433942ea},
  {32'h44f22112, 32'h41940240, 32'hc1737b96},
  {32'hc502889a, 32'h439c4378, 32'h42554287},
  {32'h44ea6c56, 32'hc3c2a279, 32'h4378408c},
  {32'hc461d263, 32'h42e0298a, 32'h3f6abce2},
  {32'h448ce264, 32'h44062bbe, 32'h4273387b},
  {32'hc2928d35, 32'hc3b86a11, 32'hc304384d},
  {32'h44d8b585, 32'h3f291d40, 32'h4348f54c},
  {32'hc4c64419, 32'h4382a92c, 32'hc28804d0},
  {32'hc32ef358, 32'hc3811a1e, 32'h431842f8},
  {32'hc1bab500, 32'h43bfe288, 32'h43b65cb8},
  {32'h44c8e2e9, 32'hc38ca60e, 32'hc38d6374},
  {32'hc3809cf0, 32'hc367314c, 32'hc2d81a37},
  {32'h44fd5ea4, 32'hc27d58f5, 32'hc3bec018},
  {32'hc29513ce, 32'hc28dce8e, 32'hc3180708},
  {32'h44f03967, 32'h431c8e04, 32'h4243739b},
  {32'hc500d518, 32'h430ca0e3, 32'hc2f70fc3},
  {32'h43fcdfa4, 32'h415a1c8f, 32'h43d3bc24},
  {32'hc51860a1, 32'hc3124155, 32'h42d8f918},
  {32'h42d255aa, 32'hc3d923b3, 32'hc3afd4fa},
  {32'hc4410d34, 32'hc3056331, 32'h43976534},
  {32'h4506c398, 32'hc2c6700d, 32'h42eff7e8},
  {32'h43d08c28, 32'h429f5512, 32'h418364b9},
  {32'h44c99d52, 32'hc2caad46, 32'h43504048},
  {32'hc501cdb4, 32'h42948ebe, 32'hc3671a3e},
  {32'h44e06eca, 32'hc2bf906d, 32'h43d42042},
  {32'hc48edae5, 32'h4324757f, 32'h4394aef9},
  {32'h43ee888a, 32'hc2168e6b, 32'h432761f6},
  {32'hc48bf304, 32'hc215c975, 32'h4305b59b},
  {32'h43d230e6, 32'hc3c4e6e7, 32'h4225a190},
  {32'hc317c660, 32'hc2f1c442, 32'h41b5e4e1},
  {32'h45069f44, 32'h433142e1, 32'hc3b43e92},
  {32'h43aa80a4, 32'h435c7a48, 32'h42a50d92},
  {32'h445d31a6, 32'h433e62ff, 32'hc2b55576},
  {32'h438ebc14, 32'h428a17b7, 32'h432971b9},
  {32'h44d0713c, 32'hc303c02a, 32'h423552d6},
  {32'hc500d11a, 32'h4295de77, 32'h439cd326},
  {32'h43f2d7f8, 32'hc32c1a19, 32'hc2bed285},
  {32'hc3cebeb8, 32'hc2bdc34a, 32'hc2cf459e},
  {32'h44bc6b1e, 32'hc38205ca, 32'hc30877e0},
  {32'hc444f0a2, 32'h42dbe87a, 32'hc30183f2},
  {32'h45128a17, 32'h43832982, 32'hc35c8916},
  {32'hc5062478, 32'h418e2932, 32'hc33414c7},
  {32'h44c7c9cf, 32'h437b1080, 32'h43b4a0eb},
  {32'h429489a0, 32'h4097e257, 32'h4290472e},
  {32'h449503b8, 32'hc2a238e0, 32'h439df3b8},
  {32'hc3eef269, 32'h43360c40, 32'hc2f56142},
  {32'h44be0cc4, 32'h427285c6, 32'hc28e715b},
  {32'hc50d6c18, 32'h42298b02, 32'hc2e03e86},
  {32'h44759976, 32'hc2206601, 32'hc3cafaac},
  {32'hc4fcab30, 32'h41a19092, 32'h42fb9fa3},
  {32'h4507f2bd, 32'hc3ce2cb4, 32'h431f4a1a},
  {32'hc3213750, 32'h41c58db2, 32'hc386fcc7},
  {32'h449e3850, 32'h42d06956, 32'hc315c260},
  {32'hc4863a72, 32'hc395bb68, 32'h4140b664},
  {32'h43e9e4fe, 32'h414fb7f8, 32'hc37470df},
  {32'hc4903b4c, 32'h4112e7ed, 32'hc3398604},
  {32'h42ee7118, 32'h428beb71, 32'hc2f69792},
  {32'hc50b5074, 32'hc2cba5c0, 32'h43653ddc},
  {32'h443ddfc5, 32'h42b1a936, 32'hc31f033a},
  {32'hc490fbe6, 32'hc300d100, 32'h43df0e72},
  {32'h44e8f2b7, 32'h408981fb, 32'h437b1bee},
  {32'hc5127da7, 32'hc3cab19a, 32'hc3d0528f},
  {32'h44f305bf, 32'hc35d7b03, 32'hc321b74b},
  {32'hc4945cce, 32'hc3012640, 32'hc40b2c51},
  {32'h4512bf85, 32'h3febbec8, 32'hc399c694},
  {32'hc5178604, 32'h43ba2eb0, 32'h400de318},
  {32'h4501779d, 32'hc26f1ddb, 32'h42daeec6},
  {32'hc3f8c872, 32'hc3dc5d08, 32'hc288822b},
  {32'h44ea6593, 32'h424db88a, 32'hc0eb7a17},
  {32'hc4fce85c, 32'h42373eb2, 32'h40fa4334},
  {32'h448e59a8, 32'hc12a11f0, 32'h43ba2b14},
  {32'hc4e86854, 32'hc127b5f9, 32'hc31eb32a},
  {32'h44cbadf7, 32'hc37526eb, 32'h43ffdd9d},
  {32'hc43787d6, 32'hc34f0f83, 32'hc33c673f},
  {32'h43f684a4, 32'hc3713b87, 32'h4314f921},
  {32'hc4ab61d6, 32'h43b8bc79, 32'hc286257c},
  {32'h431c5cc0, 32'hc1ceaeec, 32'hc344d531},
  {32'hc498fe06, 32'hc2d4aeab, 32'h4383a32a},
  {32'h44d2d1ac, 32'hc3a50942, 32'h437c9d91},
  {32'hc41bc0bb, 32'hc20a8f32, 32'h430c7ba7},
  {32'h44b2c619, 32'hc34db58a, 32'hc2e85963},
  {32'hc44949de, 32'h428642c8, 32'h41f9dd9f},
  {32'h4507e143, 32'h4106ade3, 32'hc282550c},
  {32'hc43208d8, 32'hc259eb48, 32'h43a49d49},
  {32'h44a69751, 32'h42d1f7d4, 32'h43a35407},
  {32'hc3fedb74, 32'hc378df0f, 32'hc1da3099},
  {32'h440830ec, 32'h4388af3c, 32'h43848395},
  {32'h420fa4c0, 32'hc31d221c, 32'hc2581d40},
  {32'h4505c5b7, 32'h43a627b0, 32'hc328b148},
  {32'hc505229e, 32'h43a2f351, 32'hc3b3a1b7},
  {32'h44a9b198, 32'hc3a89cf9, 32'h4390391d},
  {32'hc5035e8a, 32'h434394a9, 32'hc252fcd7},
  {32'hc3e13b0e, 32'h42d46051, 32'hc110b92a},
  {32'hc4471ace, 32'h433935e0, 32'hc3200ab5},
  {32'h44c0f940, 32'hc3532761, 32'hc319788d},
  {32'hc41963f8, 32'hc1a8fd7c, 32'hc31c263e},
  {32'h4500e600, 32'hc3974086, 32'hc2ed4b74},
  {32'hc502c7c2, 32'hc1b91367, 32'h427615a4},
  {32'h441cb530, 32'hc3dd9b27, 32'hc251dad4},
  {32'hc40841fa, 32'hc353eab7, 32'hc2820724},
  {32'h44f9fa02, 32'hc2c318c8, 32'hc272618a},
  {32'h42afa6e0, 32'hc35050ed, 32'hc2f88152},
  {32'h44c11e55, 32'hc26d3ba0, 32'h427510a2},
  {32'hc3fdc6ae, 32'h4270b50e, 32'h43966846},
  {32'h443f01b3, 32'hc380555e, 32'h411ca6ff},
  {32'hc3a1a5e4, 32'h4212023f, 32'hc3125d0a},
  {32'h44ee085d, 32'h4334b527, 32'hc2e546ce},
  {32'hc4e29427, 32'hc354b209, 32'h43cfe7fd},
  {32'h44b6c8a2, 32'h41453ef8, 32'hc316bb86},
  {32'hc4761b08, 32'hc3f96426, 32'h42656fe7},
  {32'h4483b28d, 32'h43f99dee, 32'h4342981c},
  {32'hc3fabbb2, 32'hc2b79207, 32'hc37029fd},
  {32'h40943080, 32'h43efcdcc, 32'h429d7bc5},
  {32'hc42de70a, 32'hc19d23ec, 32'hc2af04c9},
  {32'h449e5593, 32'hc3c3e3b3, 32'hc3ad9dff},
  {32'hc4a940fa, 32'hc204fb8a, 32'hc36db9b2},
  {32'h44eaddc2, 32'hc093420c, 32'hc1d4f670},
  {32'hc49f2864, 32'hc3576e1a, 32'h429071fb},
  {32'h43d70bd0, 32'hc3122f81, 32'hc28cb899},
  {32'hc4a9b9dc, 32'hc346688b, 32'h4362bd9c},
  {32'hc139d700, 32'h4323157a, 32'h43952667},
  {32'hc4df5893, 32'hc1ccb915, 32'h43441753},
  {32'h448f6e96, 32'hc36fa921, 32'hc3bb1380},
  {32'hc4daaceb, 32'hc315715a, 32'hc36ac878},
  {32'h43e90f45, 32'h42e02fc1, 32'h42a418bf},
  {32'hc4d89986, 32'h43108714, 32'h4219e7f0},
  {32'h44a78e8e, 32'h41897aa2, 32'hc35bf228},
  {32'hc500c1ac, 32'h42854adc, 32'hc29677aa},
  {32'h449a95ac, 32'h4289c270, 32'h4123a95e},
  {32'hc4a8a426, 32'h440b1a02, 32'hc2ca802e},
  {32'h448c7755, 32'h438f13d6, 32'hc2f0d4a6},
  {32'hc483c1d8, 32'hc2fc0625, 32'h41c93589},
  {32'h44801a77, 32'hc30dd4d6, 32'hc27e6f68},
  {32'hc4a459b8, 32'h434e8d77, 32'h4372be69},
  {32'h45094cef, 32'hc36d2d6f, 32'hbfef1280},
  {32'hc4c46dc8, 32'h43765ac2, 32'hc2188bc4},
  {32'h449c2fd9, 32'hc3264545, 32'hc20866eb},
  {32'hc494c0b2, 32'h426ecfac, 32'hc21e506e},
  {32'hc3470540, 32'h42ae7ba0, 32'hc25e14be},
  {32'hc38f8347, 32'hc2f9a654, 32'h429d0bb1},
  {32'h449357d2, 32'h425b4f03, 32'hc2806e7a},
  {32'hc3aa59d0, 32'hc380eefd, 32'h4324303a},
  {32'h450a5b18, 32'hc328502b, 32'hc30c18b5},
  {32'hc43e770b, 32'hc367401e, 32'h4237ceea},
  {32'h44c5d989, 32'h4322325c, 32'hc2a0786a},
  {32'hc4261c12, 32'h41b180c3, 32'hc1867141},
  {32'h4485227f, 32'hc324b68f, 32'h437575b9},
  {32'hc4a38cc3, 32'h43c8bbc1, 32'h4309c471},
  {32'h44bb0f64, 32'hc31001af, 32'h42cece38},
  {32'hc4ad96d8, 32'hc31fb246, 32'h4258a7a8},
  {32'h44e9fffd, 32'hc15fd35a, 32'h4390b750},
  {32'hc4c7dd37, 32'hc36fd2a3, 32'h420d9d85},
  {32'h44ac1f4a, 32'hc40d0bf2, 32'h4213fa40},
  {32'hc37ab6c0, 32'h4393cb6d, 32'h4386e327},
  {32'h44c882d1, 32'h41bf76fa, 32'h42edbe42},
  {32'hc40613ef, 32'hc3f416f3, 32'h434efed0},
  {32'h44e11132, 32'h4292852d, 32'hc22feb28},
  {32'hc4764ade, 32'hc36322c0, 32'h43398071},
  {32'hbfcbe400, 32'h41bc783a, 32'hc38b59e0},
  {32'hc4986bb8, 32'hc347e80f, 32'hc274cc25},
  {32'h44c3e59e, 32'hc3170abc, 32'h42a1050f},
  {32'hc4c5eb49, 32'h431b4ab7, 32'h42651a9c},
  {32'h44ebe2b9, 32'h43ab0bfc, 32'hc3aba23e},
  {32'hc3d9248d, 32'hc20f5336, 32'hc2d02b4b},
  {32'h43df8630, 32'h41d29a80, 32'hc2db40f0},
  {32'hc4ad70ea, 32'h429d063d, 32'hc2b6aafd},
  {32'h451ea398, 32'hc2125d17, 32'hc25a56f7},
  {32'hc4a28f72, 32'h43b30e09, 32'hc3c69f96},
  {32'h4464721c, 32'hc300dcda, 32'h42ae0d7e},
  {32'hc51b8f60, 32'hc32aac8b, 32'hc221ee70},
  {32'h446bea14, 32'hc3198c51, 32'h43960e07},
  {32'hc4af08b0, 32'h43c6f2a6, 32'hc22bf820},
  {32'h4510d30a, 32'hc3b45ad8, 32'h42d4000a},
  {32'hc4a6677c, 32'hc3fdfdc0, 32'hc3573d6e},
  {32'h44881a64, 32'hc306c36c, 32'hc35d506d},
  {32'hc4424ccc, 32'hc3a90dfc, 32'hc38c223e},
  {32'h44ef86d7, 32'h434e53e7, 32'hc38b4cee},
  {32'hc4e28389, 32'hc364bd11, 32'hc38f096c},
  {32'h44bf93fa, 32'hc40dda3a, 32'h40e290ef},
  {32'hc481bd89, 32'hc36142e5, 32'hc0d8ac88},
  {32'h450bd0a7, 32'h430bdfa4, 32'hc27fc350},
  {32'hc4e679be, 32'hc05e9c90, 32'h434ecd25},
  {32'h44fc14b9, 32'hc2c83ca3, 32'h43877f2a},
  {32'hc435f87a, 32'hc208e62f, 32'h42f3b44b},
  {32'h4490459a, 32'hc07ad364, 32'hc3e107e5},
  {32'hc427d0f8, 32'h4325063d, 32'h43006f16},
  {32'h44e0dc4a, 32'h409746c2, 32'h4312f56e},
  {32'hc3ca0b6a, 32'h4407ba86, 32'h4322a0e4},
  {32'h44cddd16, 32'h410d87fc, 32'h431e5527},
  {32'hc3a29c57, 32'hc38ba950, 32'h4308d236},
  {32'h44ae314a, 32'hc32df042, 32'hc1a583e5},
  {32'hc362baff, 32'hc2a70493, 32'h43497f7d},
  {32'h44d2ea8b, 32'hc332df0a, 32'hc1786400},
  {32'hc3528c80, 32'hc28d1752, 32'hc3be76d5},
  {32'h441c7468, 32'h4259a632, 32'h42a75cc8},
  {32'hc3ae5ea0, 32'hc36350f9, 32'h40f2e090},
  {32'h43b2bb52, 32'h440ddc39, 32'h42b241b1},
  {32'hc4e2f912, 32'hc2847bcc, 32'h434ecf41},
  {32'h44fcceb2, 32'hc2ea9780, 32'hc420f0eb},
  {32'hc5156552, 32'hc310d7c9, 32'h43635904},
  {32'h4494a9ec, 32'hc38032ab, 32'h416f74e0},
  {32'hc44cca7f, 32'hc329af0f, 32'hc4037750},
  {32'h4359b0d0, 32'h431dd077, 32'h42a22dcb},
  {32'hc4f0fd4c, 32'h422bee07, 32'hc38c3dd1},
  {32'h4506a552, 32'hc36cca4b, 32'h4185cfba},
  {32'hc4d67f8c, 32'h4013556c, 32'hc3272505},
  {32'h442c0be9, 32'hc37b403b, 32'hc3cbe974},
  {32'hc5106430, 32'hc3e5b622, 32'hc33f8eb2},
  {32'h43cbc9da, 32'hc295fa96, 32'hc1eea860},
  {32'hc4b3ab84, 32'h42a324a9, 32'hc29d98e7},
  {32'h450a3f12, 32'h4307969a, 32'hc1d479d0},
  {32'hc3776a1d, 32'hc38535fd, 32'h42132de3},
  {32'h44d9d5ba, 32'h43a2f886, 32'h4365e977},
  {32'hc3452b09, 32'h42939d82, 32'hc363882d},
  {32'h43ac3882, 32'h4211941a, 32'hc3211a14},
  {32'h421bf200, 32'hc369aa75, 32'h427c3f3e},
  {32'h439e8cc0, 32'hc3110ea5, 32'hc2c11da9},
  {32'hc51397cc, 32'hc1b8146b, 32'hc312933d},
  {32'h4518ef21, 32'h438d2871, 32'h42fbf922},
  {32'hc4ef7390, 32'hc24fd203, 32'hc36965b7},
  {32'h44a1a84f, 32'h41d9ad0f, 32'h43ae2692},
  {32'hc4c7aaf5, 32'hc2ca52e0, 32'h4244771a},
  {32'hc34f6860, 32'h43916b21, 32'h42e51b5d},
  {32'hc4e811a8, 32'h4263f073, 32'hc2a95751},
  {32'h44c23e65, 32'hc28218a6, 32'h433d1ed5},
  {32'hc4893808, 32'hc35e7eca, 32'hc3bb2ba5},
  {32'h44ec4df1, 32'hc281157a, 32'h417e56ac},
  {32'hc3c634c8, 32'hc3b2b247, 32'hc3b1ed0a},
  {32'h43dd61c0, 32'h43ee66e1, 32'h430337ca},
  {32'hc4c73def, 32'h428fe84d, 32'h4359f1c5},
  {32'h44fa15bb, 32'h43fe6b2c, 32'hc27b1908},
  {32'hc1c95d00, 32'hc3ca3784, 32'hc387a152},
  {32'h44da1177, 32'hc2a53fa7, 32'h43eda26e},
  {32'hc4f29e7e, 32'hc2f29d78, 32'hc2ca90ab},
  {32'h4511b6d3, 32'h431ae6fa, 32'h4384354c},
  {32'hc49bb414, 32'h43b6f3c5, 32'hc20ea8ef},
  {32'h44e39f8c, 32'hc21d77b8, 32'hc121db08},
  {32'hc5059810, 32'hc2ed74a4, 32'hc3f34b81},
  {32'h44bae63d, 32'h43b793b1, 32'hc383b82f},
  {32'hc50483ab, 32'h412af1cc, 32'hc292dc93},
  {32'h448dd19a, 32'h42063f90, 32'hc324f858},
  {32'hc3d4c5c7, 32'h437a0cce, 32'h42672dd5},
  {32'h4482c56c, 32'hc383c003, 32'h425c7cbf},
  {32'hc345ad68, 32'h4296c031, 32'h42e279f8},
  {32'h447de3ee, 32'hc3121842, 32'hc1ef6b3a},
  {32'hc4ef2772, 32'h43c8d223, 32'h42e9e4b7},
  {32'h448042cb, 32'h43c77d90, 32'hc38842c1},
  {32'hc4c05c31, 32'hc322ac87, 32'hc312ccd6},
  {32'h44addf50, 32'hc2aed924, 32'h43121780},
  {32'hc38eed35, 32'h4399cdca, 32'h436332ce},
  {32'h44ec631a, 32'h43ceaf9a, 32'hc327f8f4},
  {32'hc4fbc589, 32'h3f194a14, 32'hc345b7ef},
  {32'h444d5bfb, 32'hc358d28d, 32'hc3990fc1},
  {32'hc466e678, 32'h41e1e8d0, 32'h424e33dc},
  {32'h44901c1c, 32'h42be1758, 32'h42f36cb8},
  {32'hc505e631, 32'h431b1961, 32'h43108a2a},
  {32'h43830aac, 32'hc050bc87, 32'hc2f105b3},
  {32'hc07f3000, 32'h43b29cde, 32'h4335dff4},
  {32'h44805f63, 32'hc33aa634, 32'h43b86af2},
  {32'hc4916f86, 32'h4279ae55, 32'hc1be3a4c},
  {32'hc28d1294, 32'hc3d259a9, 32'hc2ab0c4b},
  {32'hc4f6a7d5, 32'hc2da23c0, 32'hc306cd0d},
  {32'h43276f88, 32'hc3b4dfea, 32'h42b3389f},
  {32'hc4f5f3ba, 32'h43ccf3d6, 32'h4381a597},
  {32'h44cf9088, 32'hc2d54f8d, 32'hc35c77cf},
  {32'hc417535a, 32'hc3a06f91, 32'h441a914b},
  {32'h44f41898, 32'hc1de0517, 32'hc1ec6a9c},
  {32'hc4af8135, 32'hc38e45f6, 32'hc2c619c5},
  {32'h44f43f48, 32'hc3614355, 32'hc06d6d46},
  {32'hc5078a6e, 32'hc34a7384, 32'hc2283aab},
  {32'h4345b730, 32'hc1720060, 32'h430c0887},
  {32'hc487a0bf, 32'h4232782c, 32'h434031e0},
  {32'h449d2568, 32'h418e5f92, 32'h439a9a67},
  {32'hc444bb64, 32'hc3948d05, 32'h42fa18a0},
  {32'h442dc778, 32'hc3179f05, 32'hc2885195},
  {32'hc47f1304, 32'h431e9441, 32'h433ea74f},
  {32'h44260d8e, 32'hc29fe716, 32'hc34a949e},
  {32'hc37be4b4, 32'hc304e1d0, 32'hc2ba1965},
  {32'h43ab9b8c, 32'hc2a45168, 32'hc188eab7},
  {32'hc5273722, 32'h4398687a, 32'h42198154},
  {32'h450f0a9a, 32'h429c60cc, 32'hc35eea79},
  {32'h43988948, 32'h431d60d4, 32'hc19f8684},
  {32'h44c51470, 32'hc32b6f8b, 32'h4331c67a},
  {32'hc14fcc80, 32'h43c81a07, 32'hc3497fb3},
  {32'h44b8deaa, 32'h4321dcef, 32'hc3476d8d},
  {32'hc4d56bc0, 32'hc2460eb5, 32'hc38fc20a},
  {32'h4481dcd0, 32'hc2f4384f, 32'h432382bd},
  {32'hc514ab04, 32'h438c7eff, 32'h43314765},
  {32'h44fa52ec, 32'h4336176c, 32'h41ce445a},
  {32'hc4fe7748, 32'h4218d397, 32'hc38cd6c4},
  {32'h4480bc45, 32'hc3a8e88a, 32'h43103ba2},
  {32'hc47ba772, 32'h42496178, 32'h42d48990},
  {32'h444c625a, 32'h430d03ae, 32'h41ce445e},
  {32'hc466ccb0, 32'h43538c7b, 32'h435f1925},
  {32'h4345dec4, 32'hc3a9180f, 32'h42de70f4},
  {32'hc4efa959, 32'h4297fc2b, 32'h43ac3c46},
  {32'h44639692, 32'hc30dbcb1, 32'h42d56852},
  {32'hc2083e00, 32'h430195d6, 32'hc2812886},
  {32'h443c82b8, 32'h4362ab22, 32'hc40f5358},
  {32'hc4dc8da8, 32'hc241c1fa, 32'hc1ea3227},
  {32'h43e764f4, 32'hc3290846, 32'hc3d02069},
  {32'hc5088a9f, 32'h428beeca, 32'h435594b5},
  {32'h44a4b81c, 32'h4305c97a, 32'hc3b44b31},
  {32'hc4f600bf, 32'hc2b02dcb, 32'hc34a6a70},
  {32'h44b76e85, 32'h430ae79a, 32'h42f0a07f},
  {32'hc4afa399, 32'hc392ecbd, 32'hc3188cd3},
  {32'h425a96a0, 32'h43f87589, 32'hc2d82c8b},
  {32'hc4e66f7c, 32'hc2c296e2, 32'h4215afb6},
  {32'h450159d6, 32'hc34b0390, 32'hc2a28ee6},
  {32'hc47f3248, 32'hc366022a, 32'h4389d4f3},
  {32'h44610cd2, 32'hc3674a51, 32'hc2c0fde9},
  {32'hc478be00, 32'hc3cd34c6, 32'h43ad55e1},
  {32'h4500062c, 32'h43731fc7, 32'hc102881c},
  {32'hc461e256, 32'h43133002, 32'h4329db57},
  {32'h4485c9b8, 32'h42e0960f, 32'h410f5ea1},
  {32'hc45e726f, 32'hc24e8be8, 32'hc2b38700},
  {32'h44ec1a34, 32'hc190e8a9, 32'hc394d524},
  {32'hc4c68ee5, 32'h41a6b680, 32'hc29f0ce2},
  {32'h4429511d, 32'h438affd8, 32'h408f13f9},
  {32'hc44e7972, 32'hc1890cd0, 32'h42d467db},
  {32'h44fc0d32, 32'hc3bd2879, 32'hc3c40ae1},
  {32'hc2cef158, 32'hc32ba6da, 32'h43b524dd},
  {32'h44c52a00, 32'hc28f5d8f, 32'hc22b3826},
  {32'hc4406a1d, 32'h4312c01c, 32'h4186b3f9},
  {32'h43ca18c4, 32'h4330680e, 32'h42bfcc96},
  {32'hc4826ed2, 32'hc35be724, 32'h42e1e1eb},
  {32'h41f84220, 32'h42c5d9e0, 32'hc3a4fed9},
  {32'hc3362f48, 32'hc3134068, 32'h42a0d024},
  {32'h4461dea6, 32'hc3f1ac37, 32'h430aef55},
  {32'hc413c5e8, 32'hc2a7bb16, 32'h43df07ae},
  {32'h44aec896, 32'hc3141ae9, 32'hc3b14afb},
  {32'hc4cf8126, 32'hc2a9f4ac, 32'h42846401},
  {32'h447cc2c9, 32'hc29f997c, 32'hc2fc8109},
  {32'hc4b4e1c2, 32'hc290afad, 32'hc31b24df},
  {32'h44be9ec8, 32'h4238932e, 32'h43e814eb},
  {32'h437904e0, 32'h43596d63, 32'hc38b27fc},
  {32'hc38ccc88, 32'h41d97cba, 32'hc299c5d0},
  {32'h447a9f0f, 32'h43d1e110, 32'hc30419ec},
  {32'hc4d850c6, 32'hc2fc8851, 32'hc303ba98},
  {32'h43fe38fd, 32'hc2e42fac, 32'hc1a52ea5},
  {32'hc508de2f, 32'h433fb3a8, 32'h43e60cee},
  {32'h44f5972c, 32'hc3003e9d, 32'h4307ea9e},
  {32'hc4beb809, 32'h428cdf4a, 32'hc38449b4},
  {32'h4442278d, 32'h43eca139, 32'hc13c098c},
  {32'hc44f79e8, 32'hc390957b, 32'hc3187cf5},
  {32'h4490327f, 32'h4391d5a9, 32'hc28556dc},
  {32'hc43213d8, 32'h4144c1d0, 32'h43f9f507},
  {32'h44d54af7, 32'h43e329a4, 32'hc347cb0b},
  {32'hc4fd47c6, 32'hc3eb6de4, 32'hc3785c04},
  {32'h44ddcd23, 32'h43b5a365, 32'hc35a09a2},
  {32'hc443c276, 32'hc2d0d7ab, 32'h430a4dbc},
  {32'h451394c5, 32'hc3a06704, 32'hc2ddaecf},
  {32'hc486fb23, 32'hc29d701f, 32'h425a61bc},
  {32'h44d059b4, 32'hc3b045cc, 32'hc28a63d4},
  {32'hc41b7feb, 32'h43bca980, 32'h41f14edc},
  {32'h446a0521, 32'hc393debf, 32'h41c3b35e},
  {32'hc400932d, 32'hc370d2bd, 32'h430708a0},
  {32'h442b395e, 32'hc2744660, 32'h4239ae79},
  {32'hc483be8d, 32'h4305846c, 32'h42fb075b},
  {32'h442278ac, 32'h4390e322, 32'h429d0928},
  {32'hc4bcb376, 32'h42e73000, 32'hc26ebd01},
  {32'h4356f778, 32'hc1d735df, 32'h43082174},
  {32'hc49c369f, 32'h4282be5c, 32'hc2ad1d51},
  {32'h42241c00, 32'h42bcbe4e, 32'hc3a62f38},
  {32'hc44b2e0d, 32'hc2d6c016, 32'h415d1480},
  {32'h4413750c, 32'hc2a1f9ba, 32'h4341c98d},
  {32'hc4f32575, 32'hc4181694, 32'h430f84bf},
  {32'h448e2d5e, 32'h42bc67dc, 32'hc3f87f95},
  {32'hc445cf6a, 32'hc2f29808, 32'h42c5ded5},
  {32'h45198014, 32'h424350cc, 32'h4323f829},
  {32'hc24d4cc0, 32'h42ac56a4, 32'hc3a8304e},
  {32'h4437647f, 32'h42be2f82, 32'h41abdae9},
  {32'hc4eb9d8b, 32'hc381717d, 32'hc2dd46e5},
  {32'h44eb61f4, 32'hc2b7aec1, 32'h426d7493},
  {32'hc509a691, 32'hc1d992d3, 32'hc35597ee},
  {32'h44cc716f, 32'hc31f9b4b, 32'hc35da543},
  {32'hc0ec4a00, 32'h43ef0b00, 32'h42889e8a},
  {32'hc08fe080, 32'h3f2d2c7c, 32'h4407a2e6},
  {32'hc33dd6c0, 32'h4427f8c1, 32'h43e6bdf6},
  {32'h452314ec, 32'h4271ccf4, 32'h4303a347},
  {32'hc502c6f2, 32'h42734b4d, 32'hc2a0b59b},
  {32'h429f4b40, 32'h434a2700, 32'h42991700},
  {32'hc41fe87e, 32'h430204b1, 32'hc3857b48},
  {32'h45057e0e, 32'hc2bd6b68, 32'h428a5777},
  {32'hc50697f4, 32'hc390f9be, 32'h42b274fa},
  {32'h43ff3cb0, 32'h426c77f0, 32'h4286e0c0},
  {32'hc4f526f6, 32'hc2e53ea1, 32'h403f5b17},
  {32'h44a2842d, 32'hc37c1440, 32'h4366aec7},
  {32'hc4823ec8, 32'h4393d365, 32'hc40e9a27},
  {32'h44c4d893, 32'hc37b06e5, 32'hc37ce34d},
  {32'hc3a181c8, 32'hc2804fa2, 32'hc20a43e1},
  {32'h44be6f75, 32'hc2be70b8, 32'hc3bc4536},
  {32'hc4f985c9, 32'hc255e1a6, 32'h42d13313},
  {32'h40b608c0, 32'hc23569f1, 32'hc245a1fc},
  {32'hc4135ea6, 32'h42e277e3, 32'hc3a3e3f2},
  {32'h43ebfbf8, 32'h4331cba3, 32'hc3e71496},
  {32'hc4e5b1ec, 32'hc3c4031a, 32'hc399db71},
  {32'h441bf06b, 32'h4000c73c, 32'hc23eb12e},
  {32'hc4b65ed5, 32'hc300130d, 32'h42b7fcee},
  {32'h421100c0, 32'hc221c6b9, 32'h432656ef},
  {32'hc4e19781, 32'hc16ec9b1, 32'hc0cc623f},
  {32'h44ace483, 32'hc3969e34, 32'h424557c5},
  {32'hc40d0883, 32'hc368b884, 32'h42305037},
  {32'h442f01ae, 32'hc1ab6f27, 32'h430ef96f},
  {32'hc35f6f1a, 32'h42f5d094, 32'h4321aec3},
  {32'h44dcb4a3, 32'hc2215f85, 32'hc2777d94},
  {32'hc4ed4fdc, 32'hc1e99759, 32'h4374be50},
  {32'h44b7c385, 32'h43abd1f3, 32'h406acdf4},
  {32'hc4a73186, 32'h43f7d5ae, 32'hc31e3873},
  {32'h45035a4c, 32'h43a9755c, 32'hc233db6a},
  {32'hc479c919, 32'h439ece3e, 32'hc3b779f9},
  {32'h44e10afe, 32'h43c2b3a3, 32'hc325c071},
  {32'hc4cdfd02, 32'h439240af, 32'h43b060fd},
  {32'h44bb7e3c, 32'hc32eedd2, 32'h42f97260},
  {32'hc50ea816, 32'h432fdb4c, 32'hc37cb5c7},
  {32'h450b3b0d, 32'h4295926d, 32'hc2f34740},
  {32'hc407b671, 32'hc2cbb4dd, 32'h42f7674c},
  {32'h448fbfc6, 32'h43f12afd, 32'hc2af392d},
  {32'hc4e30103, 32'h412d3e5b, 32'h4389b92d},
  {32'h44a471e2, 32'h439d4023, 32'h43278a63},
  {32'hc4cf5650, 32'h42cb25c1, 32'hc331f593},
  {32'h429c4fc0, 32'h42d140f8, 32'hc41072f1},
  {32'h4289b419, 32'hc38631e1, 32'hc33c6efa},
  {32'h439b1eea, 32'h436c63b7, 32'h43999ea8},
  {32'hc4a47014, 32'hc3350175, 32'h4345abcb},
  {32'h4458fe61, 32'hc2879210, 32'hc3bb4e98},
  {32'hc3fd02d5, 32'h43af91da, 32'h411e5f6e},
  {32'h44af56e8, 32'hc2ab67a9, 32'hc282636d},
  {32'hc45c675a, 32'h4360f79d, 32'h42db4fde},
  {32'h44eccd63, 32'hc2aa193b, 32'hc2f42e15},
  {32'hc481eb7c, 32'h4012277a, 32'hc29c1548},
  {32'h44c80ec2, 32'hc393045f, 32'h4391ce55},
  {32'hc4c7c0de, 32'hc3513869, 32'h43451fd7},
  {32'h45143d92, 32'hc328a2a2, 32'hc2f817b5},
  {32'hc46cba88, 32'h420bd4f9, 32'hc302b37c},
  {32'h445b455d, 32'h4055d1f0, 32'hc3a45a42},
  {32'hc4fd07ec, 32'hc1c61a26, 32'hc26387ce},
  {32'h4476d5ce, 32'h43089b19, 32'hc2c1dd5f},
  {32'hc5019656, 32'h40502dac, 32'h42de89fa},
  {32'h448c3c26, 32'hbfa401b8, 32'hc399c683},
  {32'hc4148968, 32'h3f0996f4, 32'hc305e77f},
  {32'h44b177af, 32'h42d70271, 32'hc2d8eac2},
  {32'hc406c6a2, 32'hc35aa112, 32'h43b3b617},
  {32'h444eb6c6, 32'hc383a791, 32'hc115a380},
  {32'hc3d63cb6, 32'hc3076a8b, 32'hc31d674b},
  {32'h449eb3d6, 32'hc1aca191, 32'h43012303},
  {32'hc49704bb, 32'h43a25d79, 32'hc28656d3},
  {32'h449a6fc1, 32'h43f6bee5, 32'hc3bca45a},
  {32'hc4bc88a8, 32'h43a9b4e0, 32'h42384bee},
  {32'h448252f5, 32'hc16d5772, 32'hc2c8a4af},
  {32'hc4db6369, 32'hc385b25c, 32'h4364fd3b},
  {32'h43166dd0, 32'hc30a59aa, 32'h43ba6373},
  {32'hc4d5718a, 32'hc35d794a, 32'h41bdcb7c},
  {32'h44426c6a, 32'h4340464b, 32'h433d5763},
  {32'hc46de6b1, 32'h437b5766, 32'h4421447b},
  {32'h44f7b28a, 32'hc39a1615, 32'h438e5275},
  {32'hc5030f97, 32'hc2ff84bd, 32'h4417279b},
  {32'h447380e3, 32'h439897d8, 32'h431b8a4f},
  {32'hc48d06d2, 32'h41729e82, 32'h4271eace},
  {32'h44856953, 32'h42b1250e, 32'h433531ab},
  {32'hc49836ab, 32'hc26b849a, 32'hc36e8830},
  {32'h4419bc35, 32'h431ce8cd, 32'h428bbe4f},
  {32'hc48ad19a, 32'h41907654, 32'h434830f4},
  {32'h44859adb, 32'h43936d2d, 32'h433dd90d},
  {32'hc5004ad8, 32'hc23fa880, 32'hc237e92d},
  {32'h43fb4098, 32'h434ff54e, 32'hc35f24c9},
  {32'hc35966a0, 32'hc3733002, 32'hc38d1206},
  {32'h44ba3146, 32'hc1bfae52, 32'hc225d406},
  {32'hc4244a3b, 32'hc31a6089, 32'hc27bb9fe},
  {32'h44fde7d1, 32'h43bd1b99, 32'hc319c841},
  {32'hc4f5acd0, 32'h429094c9, 32'hc3484cf8},
  {32'h44be9c77, 32'h41c9f8e4, 32'h41e767e4},
  {32'hc4f4a4ff, 32'h4313aeec, 32'hc31e0223},
  {32'h45054a44, 32'h42e131dc, 32'hc22e978d},
  {32'hc4cb79ac, 32'h4345b910, 32'hc1b0231c},
  {32'h44ef6861, 32'hc2c45471, 32'h429b7dd4},
  {32'hc4893069, 32'hc2b95455, 32'h4211e999},
  {32'h43941a8c, 32'h43cc01f0, 32'h42e8261e},
  {32'hc50ebd5f, 32'hc3849324, 32'hc0e70622},
  {32'h44ddd256, 32'h42fa007b, 32'h42b82b26},
  {32'hc50ad6b9, 32'h43647aab, 32'hc182f633},
  {32'h4385bfd0, 32'hc420c918, 32'h434f5ddf},
  {32'hc4e34ea1, 32'h4169179b, 32'hc2bac80c},
  {32'h449b5554, 32'h416058d8, 32'h434578b1},
  {32'hc3c92b5c, 32'h43075c30, 32'h4327b91d},
  {32'h44eae48f, 32'hc34e38b7, 32'h431d1bc7},
  {32'hc43655a2, 32'hc39d0d88, 32'h42a6f58b},
  {32'h443cf9c1, 32'hc384f60a, 32'hc2720475},
  {32'hc4f458a4, 32'h432f5461, 32'h42da43fc},
  {32'h44c82ca0, 32'hc105620d, 32'hc2390742},
  {32'hc43c89ab, 32'hc303419a, 32'hc282823e},
  {32'h451012ed, 32'h43c477ee, 32'h41aa5da6},
  {32'hc2b8cedc, 32'hc18303a8, 32'hc2ea42f2},
  {32'h4504162c, 32'hc2dabe82, 32'hc3b7f298},
  {32'hc4135f04, 32'h41276611, 32'h428bf7bd},
  {32'hc245e160, 32'h42729380, 32'h4188d276},
  {32'hc4c73287, 32'h435257f5, 32'h432ec295},
  {32'h43a98d97, 32'h42cb29e2, 32'hc38eda0d},
  {32'hc4fddf37, 32'hc3e9ec6b, 32'hc29dd5f1},
  {32'h45171d74, 32'h43155f70, 32'h43ab5111},
  {32'hc484fd0d, 32'h43df2c5b, 32'hc2c6f1ca},
  {32'h44f85de1, 32'hc3480cb5, 32'h4375e2a3},
  {32'hc4eedb38, 32'h42c98409, 32'h41f8c15b},
  {32'h44fa41e4, 32'h4305cb6a, 32'h4127980b},
  {32'hc4fdcc7e, 32'hc3b8cddf, 32'h426f6956},
  {32'h44a70c6a, 32'h434eeb52, 32'h423df98a},
  {32'hc4347a98, 32'h41257a22, 32'h42ac37c2},
  {32'h450d5374, 32'h43123115, 32'hc3ae9635},
  {32'hc3c9fafa, 32'h410587f3, 32'hc34560d7},
  {32'h4516e583, 32'h41eeda6e, 32'hc19985dc},
  {32'hc4fb9e40, 32'h4391abaf, 32'h4381a65d},
  {32'h442b9036, 32'h42950ab4, 32'h4344b572},
  {32'hc3a291a0, 32'hc34e90cd, 32'hc2fbe8a9},
  {32'h44ca628e, 32'h425705e5, 32'h437cd513},
  {32'hc50f2dc6, 32'hc2415d1f, 32'h438a0a27},
  {32'h4404b898, 32'h432cf11d, 32'h4335bd7b},
  {32'hc45d8c98, 32'h424b10de, 32'h42ba77e1},
  {32'h44e59dff, 32'h43a7db76, 32'h403fb1ec},
  {32'hc49d62c7, 32'h4265b4f6, 32'hc3e9e9b9},
  {32'h43d4477e, 32'h430f9038, 32'h4315dcbe},
  {32'hc4647f90, 32'h420651ed, 32'hc371fe9f},
  {32'h4411c630, 32'h421fa625, 32'h430585ae},
  {32'hc50667dc, 32'h43737aa8, 32'hc2a6e2e2},
  {32'h4382ed26, 32'hc2570eea, 32'h43122341},
  {32'hc435d712, 32'h44007660, 32'h43b8d5c6},
  {32'h44477550, 32'hc39944ec, 32'h43e5edd0},
  {32'hc3109a90, 32'hc3523b7b, 32'h43448ec9},
  {32'hc1f8b140, 32'hc357f5d4, 32'h41a54a46},
  {32'hc50ae537, 32'h4328726d, 32'hc3876982},
  {32'h43852640, 32'h438e3b38, 32'hc2fa93f4},
  {32'hc4d65897, 32'h42393537, 32'h431dacf2},
  {32'h45063568, 32'h43f63574, 32'hc37d4d88},
  {32'hc4eed23f, 32'hc36a262e, 32'h438f1038},
  {32'h44e2a8c1, 32'h43097991, 32'h43a6b269},
  {32'h42af4260, 32'hc35a5558, 32'h42b28812},
  {32'h44486571, 32'hc350c5b4, 32'h4250baa5},
  {32'hc4451776, 32'hc338b737, 32'h42c3667d},
  {32'h44b5e8c9, 32'hc331833c, 32'hc0517aa4},
  {32'hc46a928e, 32'h43b5a33e, 32'h43e166f5},
  {32'h4505e7a3, 32'hc2c8ecf1, 32'h4382bd30},
  {32'hc4aeabc1, 32'hc2fa5a58, 32'hc39e1a1b},
  {32'h4401c61e, 32'hc33b9eff, 32'h42c888fe},
  {32'hc44a1366, 32'h4440e526, 32'hc28a779a},
  {32'h449e241d, 32'hc29ab5bf, 32'hc3bd5306},
  {32'hc466b41e, 32'hc20a21d3, 32'h42dc6c0f},
  {32'h44a87a25, 32'h438db0bb, 32'hc3adca7e},
  {32'hc4d15d2c, 32'hc10fb362, 32'h4354cca4},
  {32'h44ca8641, 32'hc3211d16, 32'hc2f90c09},
  {32'hc3020f64, 32'hc230ba12, 32'hc2e3d61f},
  {32'h4409278f, 32'h439a506d, 32'hc0b09b15},
  {32'hc43dccbf, 32'hc3cb3baf, 32'h43006eec},
  {32'h447908c0, 32'hc3930c65, 32'hc1f9b2eb},
  {32'hc4b7b9cc, 32'hc3221422, 32'h43b8e0ea},
  {32'h45077169, 32'hc23d4853, 32'hc3cb4255},
  {32'hc430d38d, 32'h43509275, 32'h4392c8ef},
  {32'h4504a116, 32'h430d63da, 32'h43db0843},
  {32'hc4f85ad2, 32'h42846ce6, 32'hc308813f},
  {32'h44bdd889, 32'hc307b762, 32'hc30d5f0c},
  {32'hc48cb963, 32'hc3bbd195, 32'hc2f968ad},
  {32'h443fcc5f, 32'hc2821a99, 32'h4238116e},
  {32'hc4a5d9b5, 32'h4228fa2e, 32'hc30e447e},
  {32'h43f265a0, 32'hc3f9304a, 32'hc084f53e},
  {32'hc2f49149, 32'hc1eb8223, 32'hc2c495d4},
  {32'h44e59f93, 32'h41db93f9, 32'h41054326},
  {32'hc489a9ec, 32'hc3698921, 32'hc3012b33},
  {32'hc280c198, 32'hc35e41f8, 32'h43aaffb5},
  {32'hc489239f, 32'hc3c2a244, 32'hc2e6f804},
  {32'h4409d45f, 32'h439a9f87, 32'hc3e88595},
  {32'hc500433e, 32'h420bf086, 32'h4374d99b},
  {32'h44fb370d, 32'hc3115160, 32'hc3a7e898},
  {32'hc316e510, 32'hc35240c9, 32'h42c8c0b4},
  {32'h44f1ea8c, 32'h4333deb0, 32'h41bbd237},
  {32'hc4e4a950, 32'hc35cdae8, 32'h43ad4277},
  {32'h44bea77a, 32'hc4027614, 32'h44033ca6},
  {32'hc3badfd5, 32'hc3a0c412, 32'hc29702e0},
  {32'h441cbeed, 32'h42b7d64d, 32'hc264d62a},
  {32'hc3c82eec, 32'h43157c62, 32'h439c1e1e},
  {32'h43ae7571, 32'h4296fdf2, 32'h42aa8223},
  {32'h418864e0, 32'hc3392688, 32'h41de4dca},
  {32'h44e54b2a, 32'hc3d181ef, 32'h42b13a48},
  {32'hc4863170, 32'hc3232654, 32'h41e5c136},
  {32'h44b769dc, 32'hc16c9cde, 32'h411aaa6c},
  {32'hc4ce802f, 32'h432a90fe, 32'hc3097706},
  {32'h4521700e, 32'hc41349aa, 32'hc2157c90},
  {32'hc508db29, 32'hc379980e, 32'h4017d198},
  {32'h4455bc9f, 32'h437f0544, 32'hc340521b},
  {32'h432c9060, 32'hc3705f5b, 32'hc1740708},
  {32'h44a1da06, 32'hc36fd9ce, 32'h4408f9a4},
  {32'hc4a0b759, 32'hc2e76ed3, 32'hc2faa158},
  {32'h45038beb, 32'hc3f1213c, 32'hc2ed2c77},
  {32'hc48e98e1, 32'hbf9c081e, 32'hc33557fb},
  {32'h44adc969, 32'hc2c3f022, 32'hc2afcae5},
  {32'hc4cfc5b1, 32'h426ed5eb, 32'h41dce829},
  {32'h441065c2, 32'h40b7d853, 32'h42e023b4},
  {32'hc481824b, 32'h4228730c, 32'h439cdea8},
  {32'h44a4b8bd, 32'h429d84ff, 32'hc365a6a2},
  {32'hc3f16f18, 32'h43b9252b, 32'hc34c8de3},
  {32'hc3bd3dc5, 32'h42c58537, 32'h4355c26e},
  {32'hc4d0d971, 32'h42f81928, 32'hc30f547a},
  {32'h44fa8688, 32'hc13c5d1c, 32'h42c8f083},
  {32'hc488aee4, 32'hc2e6d66f, 32'hc21238a6},
  {32'h44c4c507, 32'hc340145b, 32'hc1ab7cbf},
  {32'hc48780c7, 32'h4229f754, 32'hc2eade51},
  {32'h4510358c, 32'hc31e6731, 32'h4202a250},
  {32'hc386da48, 32'h4348424e, 32'h41e3fc49},
  {32'h451f0be4, 32'hc424216c, 32'h42da08d1},
  {32'hc4e8d480, 32'hc1cb4d0e, 32'h43df3ccf},
  {32'h450934da, 32'hc3d1292c, 32'hc407f65c},
  {32'h436b9160, 32'hc38963c6, 32'hc30d7ca4},
  {32'h44ee395a, 32'h42cff90a, 32'hc3308afa},
  {32'hc3b13418, 32'hc31d487b, 32'h438a5fc3},
  {32'h4482e98e, 32'hc246acf9, 32'h4258f3e9},
  {32'hc514dd45, 32'hc39c3b50, 32'hc3198a6e},
  {32'h4462799b, 32'h43b28265, 32'hc297bc1e},
  {32'hc3ffd888, 32'h3d866ee0, 32'h434a87de},
  {32'h4508ba99, 32'h40488ad5, 32'hc2e5a1ae},
  {32'hc4dac31c, 32'hc23f8be1, 32'hc231095a},
  {32'h44be09dd, 32'h41f9b0e8, 32'h4343e1cd},
  {32'hc3417480, 32'hc3a50be0, 32'h42987718},
  {32'h450ad81b, 32'hc1bdcc51, 32'hc338ac9d},
  {32'hc4061164, 32'hc33342d8, 32'hc30cafa2},
  {32'h44ddd46f, 32'hc2b8c088, 32'h42d2b20a},
  {32'hc4332124, 32'hc3787610, 32'h439a32dc},
  {32'h4480a594, 32'hc37e8792, 32'h438e9b81},
  {32'hc51301b6, 32'hc384ec88, 32'hc3bc97ca},
  {32'h45065c2d, 32'hc2d6dbe2, 32'h421a9522},
  {32'hc513096e, 32'h436f1acb, 32'h43870732},
  {32'h4504405e, 32'hc2deb5aa, 32'hc3483ea4},
  {32'hc451f44d, 32'h4401a0ce, 32'hc20217dd},
  {32'h44526d11, 32'h433e6904, 32'hc3f7c668},
  {32'hc4b4ce3b, 32'h41513bfa, 32'h430a05e6},
  {32'h44b839ec, 32'h432cb1c9, 32'h42bbfb9b},
  {32'hc51c4b10, 32'hc353d79c, 32'h42256de6},
  {32'h4505dccf, 32'hc3092bea, 32'h428e3eb7},
  {32'hc40f052a, 32'hc401be19, 32'h42525f01},
  {32'h450b4bd9, 32'hc33d9d74, 32'hc2bbd282},
  {32'hc4217ae4, 32'h43958a9b, 32'hc3475b1c},
  {32'h43d8409a, 32'h43743297, 32'hc2595492},
  {32'hc450fd2d, 32'hc3024dcf, 32'h42c49524},
  {32'h44b73285, 32'h424347c1, 32'hc2c58338},
  {32'hc496303e, 32'h4367986b, 32'h42638d2a},
  {32'h446cf732, 32'h42b6d6db, 32'h42a67067},
  {32'hc4c8c2ee, 32'h43dce6a9, 32'h43379b47},
  {32'h44512a40, 32'hc2e4dd3d, 32'h435e4e88},
  {32'hc42eb8b5, 32'hc2f3fac6, 32'hc35ff7bb},
  {32'h44b466f9, 32'h428243a3, 32'hc196725d},
  {32'hc447f710, 32'h4380ba2b, 32'h431b098a},
  {32'h4453fe12, 32'h425871b5, 32'h4380342c},
  {32'hc4b1439d, 32'h4213b4fd, 32'hc2f71306},
  {32'h44bb2da9, 32'h435caa3a, 32'h4334f9d2},
  {32'hc4b53867, 32'hc1486da0, 32'hc2ae1b10},
  {32'h440bb1b0, 32'h41d9c4ce, 32'h42f7d7ac},
  {32'h433ffab0, 32'h42cc8279, 32'h43163ebe},
  {32'h441d0774, 32'hc382fa89, 32'hc4157975},
  {32'hc3b1df6d, 32'hc299d4ac, 32'h42f2a7f0},
  {32'h43c0a4f4, 32'h436dc2dd, 32'hc38b5264},
  {32'hc48c0285, 32'hc39c49af, 32'hc39751ff},
  {32'h4452d886, 32'h42fd733c, 32'h42749510},
  {32'hc4ebdae0, 32'hc31b419d, 32'hc2921edf},
  {32'h44bc4e35, 32'hc1624408, 32'hc3a2c8f8},
  {32'hc4ea6e7d, 32'h4301d1da, 32'hc36ebe48},
  {32'h44314c32, 32'hc22ae74d, 32'h43248629},
  {32'hc48f5b08, 32'hc2518042, 32'h421b4604},
  {32'h44ad4efa, 32'h4318a2c3, 32'h419967ac},
  {32'hc43911a0, 32'h43b8a31e, 32'h43dc4e61},
  {32'h450bf3b2, 32'hc26fac84, 32'h43c3cdc3},
  {32'hc1c5ee40, 32'hc3adf128, 32'h421b5126},
  {32'h4471b83c, 32'h42ef71fb, 32'hc341668e},
  {32'hc41c3de8, 32'hc269f5c6, 32'hc3aabf0a},
  {32'h443adc86, 32'hc306edff, 32'hc3b6f2ca},
  {32'hc47907ca, 32'h428c1208, 32'h41b59f36},
  {32'h4498dc55, 32'h430f341b, 32'hc3dbe94c},
  {32'hc434bc38, 32'h4415cb2b, 32'hc2dba97e},
  {32'h43be5740, 32'h432948f1, 32'h43858eb5},
  {32'hc3392c6c, 32'hc2f7b88a, 32'hc3a3f42c},
  {32'h450b15b9, 32'h43b2728b, 32'hc334f2ad},
  {32'hc515ce75, 32'hc3f73c0b, 32'hc1ffdc86},
  {32'h44f7465a, 32'h43d108b7, 32'hc187a9ad},
  {32'hc4bd9f18, 32'hc2bdd7ca, 32'h408944fe},
  {32'h44ee1c21, 32'h4313c8be, 32'h4362fab2},
  {32'hc43e9e05, 32'h4257ce5f, 32'hc3b90bfd},
  {32'h44d74085, 32'h423da82c, 32'hc388e006},
  {32'hc482c6b4, 32'hc16146ac, 32'h42cc7490},
  {32'h45099b64, 32'hc34a5181, 32'hc3a96b03},
  {32'hc48fd654, 32'h43a074eb, 32'hc2fcf948},
  {32'h442cfec3, 32'h42cd0469, 32'h4322e946},
  {32'hc4efe939, 32'h422a53e3, 32'h42130cd0},
  {32'h44b996b2, 32'h4240a931, 32'h42877299},
  {32'hc4a42fd8, 32'h42d159c9, 32'h43412aef},
  {32'h44f8811b, 32'hc38d9cbc, 32'h43008a9b},
  {32'hc4bd06b9, 32'hc14c8079, 32'h428e092e},
  {32'hc2b9acb8, 32'h43984cea, 32'hc2b92a70},
  {32'hc49ccca8, 32'h42c54163, 32'h434741bd},
  {32'h41299400, 32'h4386bfcf, 32'h43254182},
  {32'hc37f0c28, 32'hc2a941df, 32'h4381ebcb},
  {32'h450c62f6, 32'hc23d1d69, 32'h437b2a8c},
  {32'hc43b0aa9, 32'hc19587b0, 32'h4386987d},
  {32'hbeaa1000, 32'hc33919d6, 32'hc213685a},
  {32'hc349a0fc, 32'h429deba5, 32'h40593853},
  {32'h44243d0c, 32'hc2f665a5, 32'hc3844bc2},
  {32'hc3b17648, 32'hc265f802, 32'h42b54fd8},
  {32'h43db6e99, 32'hc3172d3b, 32'hc3623dd9},
  {32'hc3fa0450, 32'hc33fdddc, 32'hc332649d},
  {32'hc20fa1c8, 32'hc22c68f6, 32'h4322ec68},
  {32'hc3808900, 32'hc3051601, 32'h430ecb9c},
  {32'h44cb24ee, 32'h42dc13bd, 32'h43581c51},
  {32'hc3fcd42c, 32'hc2b49a4a, 32'hc2ce4d81},
  {32'h44533564, 32'hc2b8f60f, 32'h436b6faf},
  {32'hc51fe062, 32'h42ae660c, 32'h40ccf6a1},
  {32'h4402f4fc, 32'hc2f0ddcf, 32'hc3420071},
  {32'hc37ba94e, 32'h4219f468, 32'h433d74e8},
  {32'h44dd4964, 32'h4317fb4f, 32'hc3155767},
  {32'hc4d48d09, 32'h4357bfcf, 32'hc36871e5},
  {32'h4489e01f, 32'hc188f938, 32'h43151575},
  {32'hc3ce969e, 32'h4356204a, 32'hc39a4bf8},
  {32'h44b63bea, 32'h43c56217, 32'h436b4417},
  {32'hc50758fb, 32'hc338523f, 32'h4392e862},
  {32'h436c3398, 32'h432c7181, 32'h42523e3a},
  {32'hc496dd66, 32'hc3159f59, 32'hc3b5812b},
  {32'h450e77cc, 32'h418ff722, 32'hc270dee1},
  {32'hc483a584, 32'h4343bf55, 32'h43e3b7b2},
  {32'h42e5e360, 32'hc357515a, 32'h428bbf67},
  {32'hc4c81d82, 32'h422f31da, 32'hc31c5301},
  {32'h440430b0, 32'h440a7c5d, 32'h4249a07e},
  {32'hc500bb2b, 32'hc2942ea4, 32'h4331b0bb},
  {32'h4419e13e, 32'hc3e2d0c8, 32'h422fdb8d},
  {32'hc4eb1ad0, 32'hc3055c51, 32'hc37494e9},
  {32'h43c88771, 32'h43b67b7c, 32'h428c93c4},
  {32'hc4e21027, 32'h43271739, 32'h43b5f135},
  {32'h44e4ca62, 32'h4276c163, 32'hc323b899},
  {32'hc4273524, 32'hc2e7194d, 32'hc00b3edc},
  {32'h42a142e0, 32'hc3ab7d28, 32'h43c56c7b},
  {32'hc4e08a3b, 32'h436c86f7, 32'h43b06387},
  {32'h449e5bac, 32'h43d4fd19, 32'h4378d418},
  {32'hc451e05e, 32'hc1389143, 32'hc38a0ae4},
  {32'h43ec45d4, 32'h4413931c, 32'h424e3bfc},
  {32'hc50ed52f, 32'hc3d2eba6, 32'h42e72399},
  {32'h4481760c, 32'hc423d525, 32'hc3f329a8},
  {32'hc3a3ea1e, 32'h41eb5eae, 32'hc3e915be},
  {32'h4507b397, 32'hc32843bd, 32'h437fdf7c},
  {32'hc4a39e98, 32'hc3c6a51c, 32'hc3a3a77f},
  {32'h44c43e2c, 32'hc3ffcb01, 32'h4313c800},
  {32'hc3b9afac, 32'h428ddb91, 32'hc3fcab5d},
  {32'h43901398, 32'hc30751c4, 32'h4379fdf8},
  {32'hc4537d6e, 32'hc334d281, 32'hc3c1e7d5},
  {32'h447d5242, 32'hc2c00212, 32'h421458f2},
  {32'hc31835b0, 32'h439160ff, 32'h4223657d},
  {32'h4483327a, 32'hc0f00d49, 32'h443798a0},
  {32'hc30ae9c8, 32'hc3bbb6ca, 32'h4350e5b2},
  {32'h450e60ef, 32'h42980440, 32'h42f83bdf},
  {32'hc5160958, 32'h4259447a, 32'h4335270a},
  {32'h442c5d42, 32'h41052594, 32'h43357936},
  {32'hc4dde53b, 32'h434f49ab, 32'hc2b231ff},
  {32'h450cd24f, 32'h42fb990d, 32'h42f175bf},
  {32'hc5032f17, 32'hc2fef4e8, 32'hc3993e34},
  {32'h4305fde8, 32'h41c7c2ef, 32'h43447097},
  {32'hc4e4b216, 32'h42d459ab, 32'hc3315a65},
  {32'h45079f24, 32'hc1bb5b48, 32'h438af1d7},
  {32'hc4da8eb5, 32'h43b9420f, 32'h429a7f02},
  {32'h43d28b58, 32'hc2546301, 32'h4406cc42},
  {32'hc50158e9, 32'hc3a909a8, 32'h43429744},
  {32'h44529ded, 32'h43497966, 32'h41cf61ce},
  {32'hc4d3461d, 32'h41f7dcd2, 32'h427b955d},
  {32'h44d414e7, 32'h412f36c4, 32'h4280ba50},
  {32'hc3bc0a4e, 32'hc2f6dfdf, 32'hc16f0ea0},
  {32'h43c6ff72, 32'h438439d8, 32'hc1ab17bd},
  {32'h42aac920, 32'hc3b73089, 32'hc2d48765},
  {32'hc2c02960, 32'hc225ac69, 32'hc2abbdd3},
  {32'h45079d1a, 32'hc393a561, 32'h43023d30},
  {32'hbff2bf20, 32'hc3723e86, 32'hc3929fb3},
  {32'h43f6086c, 32'h4351f13f, 32'h432360d2},
  {32'hc2487092, 32'h4305c9b9, 32'hc3dc9c81},
  {32'h44d6f9f0, 32'hc2af069c, 32'h4004d81d},
  {32'hc4a38656, 32'hc15ced2f, 32'hc393c220},
  {32'h44c83e88, 32'hc264cd54, 32'h41cc3c82},
  {32'hc502ba7d, 32'h41e5a3c4, 32'hc32c99c8},
  {32'h44be815a, 32'h43d38ebc, 32'hc29d87a4},
  {32'hc501d4f8, 32'hc359c6c7, 32'hc29ca0e0},
  {32'h44c8c0a7, 32'h430f5d41, 32'h436e299e},
  {32'hc4d13e4f, 32'h43cbb39c, 32'hc3144f0a},
  {32'h44b338a0, 32'h423f76c1, 32'h43fa4c3c},
  {32'hc3de5953, 32'h42376179, 32'h42648c6e},
  {32'h44dc61bb, 32'h4391fe63, 32'hc3898d3d},
  {32'hc3e9587e, 32'hc0b25900, 32'hc3912a20},
  {32'h44896cdb, 32'hc38b5466, 32'h433228c4},
  {32'hc4a65389, 32'h43d3b0ca, 32'hc31c3542},
  {32'h442a19a8, 32'hc1df81bc, 32'h4350a382},
  {32'h419ad800, 32'h42802064, 32'hc2ebfd7b},
  {32'h44ddfede, 32'hc218f674, 32'h4324ca42},
  {32'hc4425f66, 32'h42c64db2, 32'hc02ac508},
  {32'h43d380d8, 32'h433b4534, 32'h43462f54},
  {32'hc4090d27, 32'h41ff0082, 32'hc3b51882},
  {32'h4490a752, 32'hc3a32b92, 32'h43b2e362},
  {32'hc47ca00a, 32'hc18ae146, 32'hc397eb77},
  {32'h44a60148, 32'h432dd5d9, 32'h43af7299},
  {32'hc39fa258, 32'hc339f67f, 32'hc3c15d81},
  {32'h44f7d753, 32'hc389f37b, 32'hc231834f},
  {32'hc39667cc, 32'hc3573606, 32'h42266712},
  {32'h4421b079, 32'hc3a35b9e, 32'hc3197bd5},
  {32'hc41fd0e4, 32'hc17afcd6, 32'hc34c93fe},
  {32'h43953a8e, 32'hc3a2b55d, 32'hc38455e9},
  {32'hc40ac75e, 32'h42811543, 32'hc3a0630d},
  {32'h440f9315, 32'hc309333d, 32'h42f3b537},
  {32'hc3631882, 32'hc3589331, 32'h401dd40d},
  {32'h447dd798, 32'h4296243a, 32'hc38cc712},
  {32'hc3e1e2ee, 32'hc2fb9f64, 32'h427c46af},
  {32'h44b68b42, 32'h429c00b0, 32'h43973b1b},
  {32'hc411b10a, 32'hc37c4e8a, 32'h43c28b97},
  {32'h44f6c7ac, 32'h42bdfefb, 32'h429102c1},
  {32'hc4896540, 32'h41ffef38, 32'h4237f766},
  {32'h44786626, 32'h43169ed0, 32'h43aa74ef},
  {32'hc3ef3970, 32'h42e78846, 32'h431da590},
  {32'h44f90cf1, 32'h4289f8ad, 32'h42a190f9},
  {32'h437ea8c0, 32'h41b356d3, 32'h439cade0},
  {32'h44104fba, 32'hc38e6ca9, 32'hc3e70dbe},
  {32'hc421ee08, 32'hc2d7ad50, 32'h43015884},
  {32'h44eb7490, 32'hc3a73934, 32'h42f4c320},
  {32'hc48ebcfc, 32'h437a2730, 32'h43341b55},
  {32'h44e97d82, 32'hc3da645e, 32'hc21b7a2d},
  {32'hc50240a3, 32'hc39dfe4a, 32'hc33061b6},
  {32'hc3964458, 32'hc2f3b51f, 32'hc299e388},
  {32'hc4d93832, 32'hc1d9e605, 32'hc221d480},
  {32'h4435c90a, 32'hc2ab5c91, 32'hc405629a},
  {32'hc3afeef9, 32'hc3b19ce7, 32'h42c5b66d},
  {32'h44a9099c, 32'hc176963c, 32'hc3e2608c},
  {32'hc502d163, 32'hc422ab17, 32'h42276a22},
  {32'h450a4aa4, 32'hc373fd0e, 32'h43d2c394},
  {32'hc3bcf688, 32'hc44b7baa, 32'hc371d149},
  {32'h4418fc46, 32'h43242528, 32'hc2950055},
  {32'hc4d100ba, 32'hc2ed661a, 32'h419930b1},
  {32'h4310fc00, 32'hc366b4a3, 32'hc2b30acb},
  {32'hc524d834, 32'h436b6499, 32'hc36e647f},
  {32'h4502102b, 32'hc378e953, 32'h4370565f},
  {32'hc471f8f6, 32'hc27febd2, 32'h43b565e8},
  {32'h433858e0, 32'hc37b7d5e, 32'hc32e4c9f},
  {32'hc4c29ac6, 32'hc33da89a, 32'hc3737712},
  {32'h434babcc, 32'hc41ce07a, 32'h42e37400},
  {32'hc4173a90, 32'h43509b0f, 32'h4151c5a2},
  {32'h45099f4a, 32'h433310aa, 32'h41125e1c},
  {32'hc48bc484, 32'hc38e37f7, 32'h428790be},
  {32'h437ea83c, 32'hc1e82f10, 32'hc3b5f437},
  {32'hc4baa15f, 32'hc33dad34, 32'h43063d82},
  {32'h44a83652, 32'hc2aadc61, 32'h4389cf27},
  {32'hc497c0b5, 32'hc2e36073, 32'hc3a6da83},
  {32'h44fb8155, 32'hc37f57fe, 32'hc38fbfe5},
  {32'hc4ba1213, 32'h4313681c, 32'hc14b784c},
  {32'h45268ad1, 32'h44017c44, 32'h43b0047f},
  {32'hc4497afb, 32'h43232ff1, 32'h432776ba},
  {32'h430505b0, 32'hc27da30c, 32'hc387f50e},
  {32'hc2e8c530, 32'h42ac78a1, 32'h438333ed},
  {32'h44e889f1, 32'h41ed830a, 32'h4232b70e},
  {32'hc3b058ce, 32'h4399dd60, 32'h42eb661e},
  {32'h44bc6997, 32'hc2d1412e, 32'h41964c9e},
  {32'hc42ae222, 32'h42f782e5, 32'hc1390650},
  {32'h446dc280, 32'hc3a5fa75, 32'h4385d2d4},
  {32'hc39df390, 32'hc373f9ca, 32'h418ba334},
  {32'h44e1ed81, 32'h429c6bfd, 32'hc39363d6},
  {32'hc3158f20, 32'h4316abd4, 32'hc2c61d80},
  {32'h45177c6f, 32'hc380273a, 32'hc2958416},
  {32'hc4f75447, 32'hc39f8413, 32'hc2bef431},
  {32'h441b24d0, 32'hc39ab9ce, 32'h438954e4},
  {32'hc5094e5b, 32'hc2936126, 32'hc435ed48},
  {32'hc2c62330, 32'h42340cb6, 32'hc2cdf823},
  {32'hc5077675, 32'hc1cdf1b8, 32'hc38f43fc},
  {32'h44d16754, 32'h427a1b02, 32'h421d33bb},
  {32'hc4415455, 32'hc419e25c, 32'h439566a2},
  {32'h4294ee7c, 32'hc1dac01b, 32'hc1c236eb},
  {32'hc51abff6, 32'hc34d8edd, 32'h43e4a1ac},
  {32'h44552860, 32'h434e6583, 32'h41fbfdd0},
  {32'hc4fa82c1, 32'hc3b1d4fa, 32'hc35ca26f},
  {32'h4504b1e1, 32'hc1fb2e07, 32'h4307f2dd},
  {32'hc42a054e, 32'hc3d06bb4, 32'hc353ea3b},
  {32'h4439ca28, 32'hc3280542, 32'h42884517},
  {32'hc4a887d3, 32'h43ad6355, 32'hc247ac44},
  {32'h435c5cd8, 32'h420cf7f2, 32'hc1c90a87},
  {32'hc4e5aa72, 32'h430b9483, 32'h422e41ed},
  {32'h44b6f551, 32'h4418c7b1, 32'h43139e43},
  {32'h419dd900, 32'hc3d83c72, 32'h4323f6b2},
  {32'h43b9d5b2, 32'h41b4d7b1, 32'h422578b1},
  {32'hc45b8e62, 32'hc337e286, 32'hc381e64a},
  {32'h449b7fc2, 32'hc3222edf, 32'hc2c61770},
  {32'hc4b3a91d, 32'h438b0c9e, 32'hc30b4115},
  {32'h4285a9b0, 32'hc3c58bcd, 32'hc309b296},
  {32'hc4d53f71, 32'hc39e1b55, 32'h44495453},
  {32'h44738d7c, 32'hc30c0041, 32'hc1c5ac44},
  {32'hc4a52762, 32'h435aaf06, 32'h43248a33},
  {32'h44ffdd7e, 32'hc0fc58e2, 32'hc2597dcd},
  {32'hc32fc339, 32'hc23da3fa, 32'h4215123b},
  {32'h44126f9e, 32'h43165675, 32'h41018ef3},
  {32'hc506aa99, 32'hc232d156, 32'h433965b8},
  {32'h450916af, 32'hc4089224, 32'hc3337fd1},
  {32'hc3ebeca4, 32'hc28513ee, 32'h435147cc},
  {32'h44993044, 32'h43a8dd30, 32'hc35d26c1},
  {32'hc5061b7a, 32'hc2c86234, 32'hc263cd73},
  {32'h441fcb84, 32'hc3ec3b98, 32'hc324792b},
  {32'hc4191c4c, 32'hc3d93978, 32'hc3836fd8},
  {32'h44783f06, 32'h43a7bd49, 32'h4385d345},
  {32'hc4fd78ff, 32'hc2b2b962, 32'h43a1e0a5},
  {32'h4445538c, 32'h42ef356b, 32'hc04cc484},
  {32'hc43e8b72, 32'h42a796cc, 32'hc3b7ad6a},
  {32'h4444ffb2, 32'hc266834e, 32'hc008cc39},
  {32'hc2e9a790, 32'h4271ab62, 32'hc3715796},
  {32'h44d075ba, 32'h43589f12, 32'hc3d65b53},
  {32'hc4515c72, 32'h41b88d95, 32'hc38304e1},
  {32'h44bea148, 32'h43215841, 32'hc2acf056},
  {32'hc43b51d8, 32'hc38bd648, 32'hc313a1ae},
  {32'h450a95ca, 32'hc38a0d13, 32'h42097336},
  {32'hc4632f90, 32'h436bd789, 32'hc22d2f1f},
  {32'h44a9e3ee, 32'hc38b96ca, 32'h434ee7e8},
  {32'hc4d8a87a, 32'h4110315a, 32'hc234b15a},
  {32'h42330920, 32'h4309a2d9, 32'hc3113df0},
  {32'hc45aef8e, 32'h40e9b750, 32'hc2fa4f22},
  {32'h45032de1, 32'hc2221682, 32'h4299280d},
  {32'h43a5da3f, 32'hc36a3252, 32'h42f445fa},
  {32'h44faadcc, 32'hc3369241, 32'hc2dfb7ca},
  {32'hc44d9b36, 32'h43197699, 32'h4279460a},
  {32'h44a03258, 32'hc1d42861, 32'h42f346be},
  {32'hc48ffed7, 32'h42a2361b, 32'hc30c4c6b},
  {32'h4488c426, 32'h4279c61c, 32'hc40483c5},
  {32'hc50c9410, 32'h43b20311, 32'h42d3fd8a},
  {32'h43d49dc8, 32'hc3871aaa, 32'h439c4f4a},
  {32'hc49d3bce, 32'hc353d5e6, 32'hc38eab2a},
  {32'h447d3280, 32'h4374a8d1, 32'hc28917a2},
  {32'hc4b19508, 32'h43013333, 32'hc36fce3a},
  {32'h4474d264, 32'h41f1bb82, 32'h43fae36a},
  {32'hc4f4ae0f, 32'h43388d97, 32'hc3295d4e},
  {32'h44982edf, 32'h43675a02, 32'h430abb2a},
  {32'hc4426fc0, 32'hc3573c83, 32'hc1f14f62},
  {32'h44da94dc, 32'hc2d4d2d1, 32'hc2ea3847},
  {32'hc4e625c1, 32'hc2f55e71, 32'h430c5994},
  {32'h439844b6, 32'hc39b53f6, 32'hc324637b},
  {32'hc50708ba, 32'hc27d2bf0, 32'h42075b0f},
  {32'h43db8248, 32'h432c8d02, 32'hc37a2ab2},
  {32'hc43a4945, 32'hc31ee2df, 32'hc3dcda47},
  {32'h450d1698, 32'h42c347fb, 32'h43149517},
  {32'hc45a0f06, 32'hc2cbfa1f, 32'hc30c80f2},
  {32'h44a533c5, 32'h432363e3, 32'h4335e63b},
  {32'hc496f68f, 32'h4309862c, 32'h4395342d},
  {32'h44eec46c, 32'hc399b4dc, 32'h43205c34},
  {32'h41735984, 32'h4313f355, 32'h423aba54},
  {32'h44ad03cc, 32'h42b20da3, 32'h4352d47a},
  {32'hc504c75e, 32'hc1121fd1, 32'hc281aa13},
  {32'h45121ac1, 32'h43703f5f, 32'h42892bbc},
  {32'hc4b48a79, 32'hc3259b98, 32'h41ae4283},
  {32'h43d06f74, 32'h42b5b04c, 32'hc306e148},
  {32'hc3be392c, 32'hc3c67ca4, 32'h432532d1},
  {32'h4403f530, 32'hc3713f5c, 32'hc3ca415a},
  {32'hc495e0a8, 32'hc2dd9a28, 32'hc167a827},
  {32'h444fdc84, 32'h43018de6, 32'hc3874f3a},
  {32'hc44ef484, 32'h435090ce, 32'h4194009a},
  {32'h44a32ff2, 32'h435b0286, 32'h441869d7},
  {32'hc44ab230, 32'h4248d76c, 32'hc0ceccff},
  {32'h44dc7ac5, 32'hc334ea45, 32'h41ea600b},
  {32'hc4f80aa9, 32'hc23e320c, 32'hc3061254},
  {32'h43dd7744, 32'h435e6d5d, 32'hc3057620},
  {32'hc5043998, 32'hc323c98c, 32'hc31686ec},
  {32'h44676534, 32'hc35d6930, 32'hc2b5aeb4},
  {32'hc474b5f4, 32'hc239d149, 32'h436da61f},
  {32'h44ab11cc, 32'h436b1f08, 32'h42985f35},
  {32'hc4e64b5f, 32'h42b57d95, 32'h43a9046c},
  {32'h42ec7ce0, 32'hc38cbb5a, 32'h43ecc825},
  {32'hc41218aa, 32'hc2599fba, 32'hc30b3fbf},
  {32'h43afcecb, 32'hc36d0549, 32'h42d3cc81},
  {32'hc3d09390, 32'h43c9608a, 32'h419b9ed4},
  {32'h45091201, 32'hc2921813, 32'hc14911bb},
  {32'hc42f891f, 32'h439b297d, 32'hc31930a0},
  {32'h44aebf17, 32'h4156eae0, 32'h4384978f},
  {32'hc38dbc2b, 32'h427c02cc, 32'h42e9510c},
  {32'h44d44ccc, 32'h423f8351, 32'hc3635576},
  {32'hc4feff8f, 32'hc3302a71, 32'h43bc531d},
  {32'hc2854123, 32'hc05d59ed, 32'h406176df},
  {32'hc4f6b76e, 32'h438bf15f, 32'hc3826ffd},
  {32'h447cc048, 32'h42d3b3bb, 32'hc321223c},
  {32'hc511e55e, 32'h4316759b, 32'h43a26221},
  {32'h4505ac8c, 32'hc37dbc9b, 32'h43e4dc2a},
  {32'hc4b542fc, 32'h41c55626, 32'hc35b6fa8},
  {32'h447793ee, 32'hc3849b71, 32'hc30c9c90},
  {32'hc48de35f, 32'hc200abc8, 32'hc33c0fa7},
  {32'h44f3ea77, 32'hc2bf3168, 32'h43365708},
  {32'hc3c2aa80, 32'h42c2ba97, 32'h4118ef3f},
  {32'h43e42c9c, 32'h4383d08e, 32'h43e68bb1},
  {32'hc4e445c9, 32'hc3530124, 32'hc30aaa3f},
  {32'hc2484aa0, 32'h40ec2f35, 32'h4392fd85},
  {32'hc3125a32, 32'h42adace9, 32'hc39d74ed},
  {32'h4428d13e, 32'h4398614a, 32'h43841db2},
  {32'hc4b62db2, 32'hc3a5c446, 32'h4239e8e0},
  {32'h44093d4c, 32'hbfc6d018, 32'h4315f812},
  {32'hc3ff3dbc, 32'hc13277d7, 32'h4150947c},
  {32'h434bb459, 32'h439bb8ed, 32'h43ee4265},
  {32'hc494080a, 32'hc26df2b9, 32'hc378a016},
  {32'h4431ddac, 32'h431f60bc, 32'h43ce19df},
  {32'hc43cbc14, 32'hc3fa7cd7, 32'hc3a0037a},
  {32'h4490eb10, 32'hc40551c1, 32'h41ed8edf},
  {32'hc50a80ab, 32'h3f87e972, 32'hc3695fc7},
  {32'hc3450448, 32'hc4074955, 32'hc3090ffa},
  {32'hc50814c3, 32'hc2057795, 32'h44154f22},
  {32'h4405c0bb, 32'hc34b481d, 32'hc2b6e508},
  {32'hc41dae14, 32'h4314b71f, 32'hc3165035},
  {32'h44f2e098, 32'h42837c8d, 32'hc3939b32},
  {32'hc458db92, 32'h42350e44, 32'hc28efaca},
  {32'h4401ced4, 32'hc30386f4, 32'hc3703b06},
  {32'hc2b78fa0, 32'hc2d6b2ca, 32'h42cca8ff},
  {32'h43a5b578, 32'h43def68f, 32'h433e4aa5},
  {32'hc463f0ec, 32'hc3782330, 32'h42a7598b},
  {32'h43107df8, 32'h43898899, 32'h43574a29},
  {32'hc384f5ec, 32'hc3888bcf, 32'h437f2837},
  {32'h44327688, 32'h41d5a54b, 32'h4305b548},
  {32'hc4e5026b, 32'hc38de854, 32'hbfe4eb62},
  {32'h438d5f2f, 32'hc2de913a, 32'hc1c1db14},
  {32'hc4e6a530, 32'h43956f74, 32'h41e42063},
  {32'h443d9f51, 32'hc1f32312, 32'h429cdf5f},
  {32'hc3e7b4fc, 32'h43eca45e, 32'hc27b0819},
  {32'h44881f5a, 32'hc33cbc6e, 32'hc39f972b},
  {32'hc41042c9, 32'hc2b20ee6, 32'hc3bbc192},
  {32'h450011c4, 32'hc3627867, 32'hc31b502c},
  {32'hc5088423, 32'h420758bf, 32'h42ee09c9},
  {32'h450e793c, 32'hc269700d, 32'h438d4251},
  {32'hc348cd68, 32'hc33a338e, 32'h4314d616},
  {32'h44e0396a, 32'h42b67f2b, 32'h41d08beb},
  {32'hc493f639, 32'hc12c3258, 32'h4388ff88},
  {32'h43408dbc, 32'h43b0d9fb, 32'h42464a25},
  {32'hc337e770, 32'h4384e37c, 32'h4342735e},
  {32'h44c1a34c, 32'h42fb2ca3, 32'hc3a1daa3},
  {32'hc3ceae78, 32'hc3be338b, 32'h43d2f7ad},
  {32'h444de27c, 32'h437c2787, 32'hc1fe390e},
  {32'hc2223fbc, 32'h44526d85, 32'h40cd94d3},
  {32'h442730a2, 32'h42fb55a7, 32'h425cf3c1},
  {32'hc5010d91, 32'h42d981e3, 32'hc334af22},
  {32'h44f7d4c4, 32'h4344a40f, 32'h41cbf065},
  {32'hc495683b, 32'hc3e1beaa, 32'h43368d30},
  {32'h4392391e, 32'h42974846, 32'h42b63c8f},
  {32'hc3ee636c, 32'hc239ce95, 32'hc38d964a},
  {32'h442f3042, 32'h41b033b1, 32'hc201aa38},
  {32'hc467c7cd, 32'hc2be58d1, 32'hc20ab189},
  {32'h43c0af8c, 32'h439a26e3, 32'h43900657},
  {32'hc50b70d9, 32'h43453aa9, 32'hc368e55a},
  {32'h439116a1, 32'hc289d669, 32'h422eaa93},
  {32'hc500a26d, 32'hc2296da7, 32'hc291a18c},
  {32'h44e44f61, 32'h42287aba, 32'hc3d54ea1},
  {32'h42527463, 32'hc3662c53, 32'hc3876963},
  {32'hc0ee1700, 32'hc18b5f2a, 32'hc32c0a83},
  {32'hc4572032, 32'hc3818bf4, 32'hc2824997},
  {32'h443ea10f, 32'h42d22805, 32'h42f16f1b},
  {32'hc4e9da41, 32'h440c3db2, 32'h43f1c7b9},
  {32'h44394e48, 32'h425aba53, 32'h432f987f},
  {32'hc4d35d20, 32'hc2df8f68, 32'hc3d2b9f9},
  {32'h4438528a, 32'hc38d2f61, 32'hc2db48c6},
  {32'hc509e245, 32'h426ba855, 32'h40836f23},
  {32'h4406eb85, 32'h434ac48d, 32'hc34a54cc},
  {32'hc518d02c, 32'hc2a3fab4, 32'h431c4063},
  {32'h44fc7f7f, 32'hc3d822f8, 32'h42c2cead},
  {32'h42986660, 32'h430fa4f9, 32'hc248658f},
  {32'h44d81fb6, 32'h40f991e7, 32'hc39850ff},
  {32'hc4c92669, 32'h439268d8, 32'h42d19ecf},
  {32'h43f00dd8, 32'h43b5993f, 32'hc1e37c5a},
  {32'hc4585b8a, 32'hc392cfad, 32'hc163574f},
  {32'h4511b410, 32'h42030486, 32'hc1dc85f3},
  {32'hc3b71848, 32'hc238e65f, 32'hc3a3cd81},
  {32'h44161b05, 32'h4324829c, 32'hc3232da8},
  {32'hc4472f68, 32'hc3b540ae, 32'hc2c00809},
  {32'h4407b030, 32'h42c7a571, 32'hc21c9141},
  {32'hc4253d35, 32'h42eb3f96, 32'h43e9d422},
  {32'h450aa21d, 32'hc3fe8ecc, 32'h41dcf272},
  {32'hc4743b51, 32'hc2d8c184, 32'h42221efa},
  {32'h44f44f0a, 32'hc2121efb, 32'h425e8d1e},
  {32'hc4be5d5c, 32'hc30d4aa0, 32'h43bcee4a},
  {32'h44eb948e, 32'hc2a78dd1, 32'h42bb09d9},
  {32'hc3e5f96f, 32'hc31b4da5, 32'hc38646e9},
  {32'h4503e3ed, 32'hc15645dd, 32'hc10d3b78},
  {32'hc500d4d0, 32'h42cc0203, 32'hc307c236},
  {32'h44eca185, 32'hc30d9abf, 32'hc3194663},
  {32'hc4aa1ee6, 32'hc382e26e, 32'h43555d95},
  {32'h43d144e3, 32'h431eb838, 32'hc269f928},
  {32'hc4dace42, 32'hc2d382c9, 32'hc3a5afe3},
  {32'h450647db, 32'h43ab02c8, 32'hc3249be2},
  {32'hc506770c, 32'hc337942d, 32'h4346794c},
  {32'h44f93236, 32'hc3c147be, 32'h43853474},
  {32'hc424264e, 32'hc2f73b01, 32'h43098bb6},
  {32'h4481f524, 32'hc3614344, 32'hc30d3077},
  {32'hc4d7b3f3, 32'hc2ed06e5, 32'hc33f5eac},
  {32'h443e19bc, 32'hc196d63f, 32'h43e8cfe5},
  {32'hc41f4d6c, 32'h4298db99, 32'hc28a27ac},
  {32'h44d74b62, 32'hc3202c55, 32'h43b6be7e},
  {32'hc42d9658, 32'hc3846e3a, 32'hc4124134},
  {32'h44312a9a, 32'hc1b79158, 32'h43c20d7a},
  {32'hc50515b6, 32'h433ad437, 32'h42bf1b6b},
  {32'h44cb32e8, 32'h4385fdfd, 32'h43c97069},
  {32'hc3c15360, 32'h42e44670, 32'hc393690b},
  {32'hc2149540, 32'h42c81dc0, 32'h438aed36},
  {32'hc49aaab2, 32'h43c0e103, 32'hc38d1fe4},
  {32'h44ed439f, 32'hc37b708b, 32'hc30dfe14},
  {32'hc4b88241, 32'hc1b7841a, 32'hc1c30da2},
  {32'h44810732, 32'hc35f2ee8, 32'h43476430},
  {32'hc481e898, 32'hc3bd3ede, 32'hc3b5a742},
  {32'h443047c4, 32'h435f8954, 32'hc393d5e4},
  {32'hc4c15095, 32'h4378ea3d, 32'h44009b0a},
  {32'h44851741, 32'h42c01a8c, 32'hc31927d8},
  {32'hc4d6df40, 32'h43aae3e8, 32'hc318af97},
  {32'h44fce3e7, 32'h429b73fb, 32'hc2c94baf},
  {32'hc4e5700a, 32'h436ad0a7, 32'hc2f11456},
  {32'h442ba45c, 32'hc215f2a0, 32'h43afa34c},
  {32'hc4b3e69f, 32'h42e05cf0, 32'hc2e1b4dc},
  {32'h44895620, 32'hc397879c, 32'hc3b25b90},
  {32'hc427f11c, 32'h42f5015e, 32'h4397c205},
  {32'h450daf39, 32'h43b3bcd5, 32'hc3e6f8f0},
  {32'hc303dd40, 32'hc1cd752a, 32'h42841104},
  {32'h437bc520, 32'hc2a2882a, 32'hc4021051},
  {32'hc4b31af6, 32'h43a9483a, 32'h433483fb},
  {32'h449514fe, 32'hc3862bb1, 32'hc38d4b7f},
  {32'hc468705e, 32'hc3541685, 32'h42b928d4},
  {32'h43c52958, 32'hc153ffc7, 32'hc34681f2},
  {32'hc5196b27, 32'hc3d33cbf, 32'h42b914e2},
  {32'h449da64a, 32'h43d30068, 32'hc36755a0},
  {32'hc4c209fe, 32'h4365397e, 32'h4362e4e0},
  {32'h44da3040, 32'hc32fe673, 32'h42d0e891},
  {32'hc48e480d, 32'hc392cf94, 32'hc1df0e22},
  {32'h44586ef2, 32'h4139355c, 32'hc031d9c8},
  {32'hc4d5a5f6, 32'hc39358a0, 32'h43717fb3},
  {32'h443bb2e4, 32'hc2047a8d, 32'h4377be3c},
  {32'hc4eeb035, 32'h40e15b99, 32'h436d6879},
  {32'h43d652e8, 32'hc2a83da6, 32'hc4026ab2},
  {32'hc4d7d3b4, 32'hc1ac9f5b, 32'hc3161b26},
  {32'h4330dccc, 32'hc29cf862, 32'h424fa7d9},
  {32'h43120ecf, 32'hc1333385, 32'hc23d10d2},
  {32'h44315916, 32'h437e2f42, 32'hc3493bee},
  {32'hc2f9df00, 32'hc28ba6c0, 32'hc3948348},
  {32'h449a610d, 32'h41354393, 32'hc1a4fefe},
  {32'hc51ac1f0, 32'hc30441c0, 32'hc297144c},
  {32'h448bbb94, 32'hc2d9d3a2, 32'h436189f9},
  {32'hc3b90284, 32'hc2593a82, 32'hc323082a},
  {32'h440dec5a, 32'h4268a2ec, 32'hc2220df2},
  {32'hc4a705ae, 32'h42b1ab5f, 32'h43aba4e0},
  {32'h44cc2fe2, 32'h43370494, 32'hc1f6e54f},
  {32'hc4a42f04, 32'hc32bcacd, 32'h4387479c},
  {32'h42fea730, 32'h42b82268, 32'hc36199d4},
  {32'hc412eec5, 32'h428cabee, 32'h43b057c5},
  {32'h447b1446, 32'hc3894673, 32'h42d2e808},
  {32'hc3d7e02e, 32'hc38d5855, 32'h43e6af3a},
  {32'h44439e07, 32'h4401e54f, 32'hc0df3cda},
  {32'hc3d41adf, 32'hc3dabe3f, 32'hc3b983db},
  {32'h4386e47d, 32'hc0c41e76, 32'hc352ef85},
  {32'hc489b973, 32'hc2cfbc71, 32'hc3ae5d12},
  {32'h44eff973, 32'hc19fdc04, 32'h433a11bc},
  {32'hc48b5aaa, 32'h433b3198, 32'h4378f904},
  {32'h434b52a0, 32'hc399e3cf, 32'h43b8398f},
  {32'hc50f998e, 32'hc3827060, 32'hc34cbce3},
  {32'h4354d2a8, 32'hc388a8f0, 32'hc3415d08},
  {32'hc3224dd0, 32'hc34b93f4, 32'hc3972a6c},
  {32'h44f22f1a, 32'h42b62f26, 32'h4364754f},
  {32'hc3ece224, 32'h423f5174, 32'h4347fc14},
  {32'h43dacbec, 32'h43ee1ff2, 32'hc383e62c},
  {32'hc3f29228, 32'hc3556f65, 32'hc3355d13},
  {32'h435f323c, 32'h41caa7c3, 32'hc2dbe816},
  {32'hc4eba1d5, 32'hc39a1829, 32'hc284afbd},
  {32'h44a04bed, 32'h4352ea97, 32'h402eb9fc},
  {32'hc4703c7e, 32'hc31c366a, 32'hc3a78adf},
  {32'h448ebc5f, 32'hc3b27f55, 32'hc38ee901},
  {32'hc496bcba, 32'h400fe5b0, 32'h431fa3f3},
  {32'h44fb624f, 32'h42189776, 32'hc3153f00},
  {32'hc44f52f2, 32'h43077e31, 32'h434b29c7},
  {32'h44953b24, 32'h437bcfb8, 32'h42a17820},
  {32'hc392d7cc, 32'hc36fa165, 32'h43992087},
  {32'h451e57cc, 32'h42bd525b, 32'h42fee189},
  {32'h413b9dc0, 32'h4307db8f, 32'h43fe79fd},
  {32'h44eb5c44, 32'h4384f95b, 32'hc25324fa},
  {32'hc4a8c2d5, 32'hc3acdee7, 32'h41b077c6},
  {32'h44b5eb96, 32'hc11d157e, 32'hc2c970aa},
  {32'hc513a22e, 32'h41892bf7, 32'hc2ce39b0},
  {32'h43e5ba3b, 32'hc2896f67, 32'h412b7ba6},
  {32'hc5085efe, 32'hc056e390, 32'hc2aa08c1},
  {32'h44eade72, 32'hc1770ddf, 32'h420005ce},
  {32'hc48d365f, 32'hc28c1f7f, 32'h4357dfae},
  {32'h44c568f4, 32'h428a3f55, 32'h420b5ede},
  {32'hc43cc6f8, 32'h43b3439f, 32'h41908c60},
  {32'h44cdd6bb, 32'h4216763e, 32'hc38ed84c},
  {32'hc3adcdd2, 32'h43d63676, 32'hc2dd902b},
  {32'h44d62a10, 32'hc3bf9766, 32'hc114de2e},
  {32'hc4f438f1, 32'h4270823c, 32'h423cd05d},
  {32'h451a9342, 32'h422bb3e2, 32'hc0e731aa},
  {32'hc4f42cb9, 32'hc38ee4e8, 32'hc34c521a},
  {32'h44c266e0, 32'hc2bbd282, 32'hc38e5480},
  {32'hc4869e64, 32'h428c2e06, 32'hc2ce23bb},
  {32'h4504398c, 32'h43142184, 32'h429dbce7},
  {32'hc49ed68e, 32'hc28330cc, 32'h42d876c5},
  {32'h44e7a820, 32'h43d5094e, 32'hc3a8c595},
  {32'hc41af16a, 32'h422aa4ce, 32'hc24eb25c},
  {32'h4499ad34, 32'hc3b1919e, 32'hc3e089a6},
  {32'hc48415ec, 32'h4293a951, 32'h43345083},
  {32'h42bea1b4, 32'hc2888a40, 32'hc278a028},
  {32'h419bd2dc, 32'hc08f0f39, 32'h4378f199},
  {32'h4424cb72, 32'hc2fa42e4, 32'h42d34abf},
  {32'hc33d8610, 32'hc23ed7b2, 32'hc2cb6dc4},
  {32'h43e03672, 32'h43337998, 32'hc2cb42cf},
  {32'hc38a0132, 32'hc3176da4, 32'h41eed24c},
  {32'h44e209a2, 32'h43440875, 32'hc36f6629},
  {32'hc37bb088, 32'h43584447, 32'h43b6608c},
  {32'h45184bf2, 32'hc419cdbc, 32'hc33e6ef1},
  {32'h430fae30, 32'hc31b7788, 32'h42f23a3e},
  {32'h447587c8, 32'hc3900914, 32'h4387618b},
  {32'h44e07bf9, 32'h42958c1f, 32'h41b13644},
  {32'hc45050a6, 32'hc2e08d0e, 32'hc2d4e331},
  {32'h436f8380, 32'hc3f20d1d, 32'h4271e25e},
  {32'hc3a0089a, 32'h420b3993, 32'h44304cda},
  {32'h43c83377, 32'hc386fb26, 32'hc3c64ca3},
  {32'hc34a3f08, 32'h4317ee1e, 32'h43bebcab},
  {32'h44987bbe, 32'hc28fe71a, 32'hc3a28499},
  {32'hc4523252, 32'hc36050a3, 32'h431c030c},
  {32'h44cb9703, 32'hc25b6f72, 32'hc30a76cf},
  {32'hc41801cc, 32'h439e3719, 32'hc3e9be5a},
  {32'h44b2c8b8, 32'h42ffcb6a, 32'h42301ef7},
  {32'hc3e62758, 32'hc36c0733, 32'h420251b2},
  {32'h448fea7f, 32'h43a0066e, 32'h4260d3cc},
  {32'hc42fc447, 32'hc3b2199f, 32'hc383c5ea},
  {32'h4386eb4c, 32'h427e07ce, 32'h41e28330},
  {32'hc4eaa279, 32'hc34dba53, 32'h433129b0},
  {32'h43c7af87, 32'h43493594, 32'hc1cd647e},
  {32'hc43cd61e, 32'hc37d5ca1, 32'h411d1498},
  {32'h44a1bad9, 32'h40746298, 32'h42e0c91c},
  {32'hc4bd584d, 32'h437e081f, 32'hc34ce08c},
  {32'h44f61f17, 32'hc29af98a, 32'h4325e4f4},
  {32'hc51d0fec, 32'h43db21c0, 32'h42bb95b4},
  {32'h44ffca99, 32'hc39287c7, 32'hc3f05b78},
  {32'hc4ab425e, 32'h43425af8, 32'hc2d9de45},
  {32'h44e2b362, 32'h41afc02a, 32'hc208a2fa},
  {32'hc4b16dbe, 32'hc38d4a5b, 32'h43965019},
  {32'h43ca59d0, 32'h4381e38e, 32'hc21940b0},
  {32'hc4b1f594, 32'hc3c38ed5, 32'h432fac87},
  {32'h44e4c415, 32'h43e944aa, 32'hc33632bb},
  {32'hc50c9d2f, 32'hc41677a9, 32'h42f4f2bb},
  {32'h446979b2, 32'hc3ba0bc3, 32'hc31b2faf},
  {32'hc3fe1661, 32'hc329267a, 32'hc21d31fd},
  {32'h4388d85c, 32'hc3d03717, 32'hc39f7295},
  {32'hc3d96ec1, 32'hc2aa5e74, 32'hc1b2f769},
  {32'h443f296f, 32'hc29bdc4a, 32'h4264a997},
  {32'hc515c528, 32'hc2a78348, 32'h423660d6},
  {32'h44f9fbe2, 32'hc3d95fa2, 32'h42f4fb78},
  {32'hc49159a9, 32'hc3b0ee71, 32'hc31cf7e4},
  {32'h446d71d0, 32'hc39e0bfb, 32'h43e6abbd},
  {32'hc28f9cc5, 32'h426e8d23, 32'hc3cc9284},
  {32'h44d13d4a, 32'h4314ea23, 32'h422b7109},
  {32'hc4a0253c, 32'hc328cd1f, 32'h4324dc6c},
  {32'h451747d6, 32'h43801eeb, 32'hc3629c8e},
  {32'hc50df7b5, 32'hc343327d, 32'h4289c028},
  {32'h44899ef0, 32'hc0a3063c, 32'h43b744fb},
  {32'hc4ddb9ee, 32'h438f4faf, 32'h43ae9bb3},
  {32'h43980ae6, 32'hc336434e, 32'h414ade64},
  {32'hc4b2cf03, 32'h4400ef46, 32'h437b07c8},
  {32'h4406bd57, 32'h410a1209, 32'hc3122412},
  {32'hc50c8b8e, 32'hc2b3341f, 32'h43018909},
  {32'hc2715350, 32'h43689cfe, 32'hc284f71a},
  {32'hc4551194, 32'hc382bd21, 32'hc388f285},
  {32'h449b33ab, 32'h41339c25, 32'h43239554},
  {32'hc3cd3606, 32'hc317a3fa, 32'h4393faf2},
  {32'h44f34f21, 32'hc2c13e02, 32'hc311b140},
  {32'hc4f7968c, 32'hc361dce7, 32'h422ab9f5},
  {32'h441ccf04, 32'h40857f6a, 32'hc33d78ce},
  {32'hc49df52d, 32'h42852d1e, 32'hc41a7274},
  {32'hc19ce550, 32'h43511f84, 32'hc3c7b58f},
  {32'hc4d33979, 32'hc36a648d, 32'h42e8646d},
  {32'h450fb4ae, 32'h437b7ccc, 32'h436e6330},
  {32'hc46150c0, 32'h438a1217, 32'hc1b9cfc6},
  {32'h4418b11a, 32'hc11f2a60, 32'h42af7c61},
  {32'hc5012671, 32'h4224e80c, 32'hc35747c5},
  {32'h44913052, 32'hc30c64b0, 32'hbfe09968},
  {32'hc509233e, 32'hc35d1f96, 32'hc32199ec},
  {32'h452d7c98, 32'h4293e887, 32'hc3a42a07},
  {32'hc46b6a98, 32'hc373095c, 32'hc21fb35a},
  {32'h44d20fd1, 32'hc301a437, 32'h4302cdd8},
  {32'hc49a7389, 32'h41977283, 32'h41d2ab36},
  {32'h4448cc28, 32'hc358f06e, 32'hc302ac7e},
  {32'hc3d66a80, 32'h439e9399, 32'h439c36ec},
  {32'h44cb4c7c, 32'h4323e22a, 32'h424b4c81},
  {32'hc3f61022, 32'h43671bf1, 32'hc377ac08},
  {32'h450148d0, 32'h42886e26, 32'hc2a77ca5},
  {32'hc3c7e3db, 32'hc3b485ce, 32'h437a41ad},
  {32'h44d40e6d, 32'hc27279d5, 32'hc3a5e9d0},
  {32'hc4992d97, 32'hc259033f, 32'hc2f75a5c},
  {32'h4516c984, 32'hc30ef9a5, 32'h4340f1b4},
  {32'hc4c93b3c, 32'hc39daa82, 32'hc1f7497f},
  {32'h44c809a0, 32'hc389ae4f, 32'h42414710},
  {32'hc494bd1b, 32'hc1c128dc, 32'hc2e04ef5},
  {32'h451fb165, 32'h42f60637, 32'h410f7d8c},
  {32'hc26b0b78, 32'hc2b20919, 32'hc398f6cd},
  {32'h443785ce, 32'h435b5e3c, 32'h4223f716},
  {32'hc3cf1dac, 32'hc209490c, 32'hc33be68f},
  {32'h44b458ce, 32'h41e3c24c, 32'h403ff340},
  {32'hc511746e, 32'h4207967c, 32'h427ab35a},
  {32'h44a7cf18, 32'hc38cb33f, 32'h42f3608a},
  {32'hc30090b0, 32'hc359c791, 32'hc2ae7b0d},
  {32'h43e8ecd2, 32'hc12b6cea, 32'h435a8992},
  {32'h4325e0a3, 32'hc30267c8, 32'hc303ebd3},
  {32'h44ad65c6, 32'hc3946e8a, 32'h4268f5c9},
  {32'hc41e5274, 32'hc389948f, 32'hc3d59008},
  {32'h43934460, 32'h42a8893e, 32'h42f9d995},
  {32'hc4bcb9fe, 32'hc3978f55, 32'hc3752f89},
  {32'h4462b9fb, 32'hc35a551b, 32'h4284e0d2},
  {32'hc4e12b5e, 32'hc0e04cf0, 32'hc3424e11},
  {32'h4327dca0, 32'hc3b1cbd4, 32'hc310e6ec},
  {32'hc474a169, 32'h43b431a7, 32'h43efcde5},
  {32'h44a3b854, 32'h43791511, 32'h428fa738},
  {32'hc3466783, 32'h43bb0406, 32'h42cecde2},
  {32'h44e99588, 32'h4321a906, 32'h42c3b97e},
  {32'hc436996f, 32'hc30c75ff, 32'h43b63f94},
  {32'h44ec86b2, 32'h434c48f9, 32'hc0babc87},
  {32'hc49b69b0, 32'hc2e41c4c, 32'h41dafe6f},
  {32'h4515a862, 32'hc150be05, 32'h41003cb2},
  {32'hc462114a, 32'hc3102158, 32'hc03e8d94},
  {32'h44ddbd1f, 32'h431cb836, 32'h42d5dfad},
  {32'hc3044a98, 32'hc1cf0a6e, 32'hc30eae25},
  {32'h44e7b2d4, 32'h42b72d39, 32'hc2a92a1f},
  {32'hc4df4634, 32'hc40459ea, 32'h43d4bce9},
  {32'h44f14b0e, 32'hc2bdb4d9, 32'h42ff473e},
  {32'hc45b0698, 32'hc32e63f9, 32'h433300c4},
  {32'h449ef040, 32'h43835f72, 32'h43c60e63},
  {32'hc4af7368, 32'hc3611f5b, 32'h4327d5f8},
  {32'h43298d90, 32'hc3b9c246, 32'h43945d00},
  {32'hc51c6124, 32'h43eeb074, 32'hc363678a},
  {32'h43a78d5c, 32'hc33af50b, 32'h42823333},
  {32'hc3f9cf54, 32'hc06cbf6a, 32'hc18cd9cb},
  {32'h45084e78, 32'h432d5c0a, 32'hc3c2d8c5},
  {32'hc429c225, 32'h435b865d, 32'hc354f98f},
  {32'h426591b8, 32'h42341d67, 32'hc2e43521},
  {32'hc473f52e, 32'h41c73f1e, 32'hc3a0d95e},
  {32'h44160bdc, 32'hc3f12b93, 32'hc35dbca9},
  {32'hc46d9c4c, 32'hc3cfa14e, 32'h439b84a7},
  {32'h44fc9d93, 32'h4298cdb2, 32'h440a14da},
  {32'hc4109a63, 32'h4318310e, 32'hc3344fb7},
  {32'h449971ca, 32'hc3a40b73, 32'h43493d31},
  {32'hc4fb39ba, 32'h41d9858a, 32'h437a905c},
  {32'h44a48af1, 32'h420609cc, 32'h4413e0bd},
  {32'hc481b99e, 32'hc36344f0, 32'h4218c683},
  {32'h440baee5, 32'hc2a00592, 32'h42d30fc8},
  {32'hc317a1e7, 32'h43b533ee, 32'hc34e7029},
  {32'h453d47b4, 32'h435dea63, 32'h43034f91},
  {32'hc4cf6162, 32'h428bab21, 32'hc28012cf},
  {32'h43bbd9ea, 32'hc2953148, 32'hc2974e07},
  {32'hc4101d98, 32'h414edd7c, 32'hc0c85cf8},
  {32'h44d6aebc, 32'h436c14cd, 32'hc3ec9b4b},
  {32'hc4e3aae8, 32'h4245a0bd, 32'hc2ad12a8},
  {32'h44e21425, 32'h432b8d8e, 32'hc33c8dc6},
  {32'hc46c3ce5, 32'hc3a2b8ff, 32'h4295db08},
  {32'h4504401c, 32'hc3881cb5, 32'h432a1a00},
  {32'hc4e4c28a, 32'hc36a259a, 32'h434566b9},
  {32'h445d36be, 32'h41e3236c, 32'hc35f31ea},
  {32'hc4c5068f, 32'hc089b91c, 32'hc31743d4},
  {32'h444b5894, 32'hc3801a6f, 32'hc382b668},
  {32'hc4407806, 32'h43e5b5e3, 32'h43d89529},
  {32'h44db00fd, 32'h42e4e1fb, 32'hc3b0f36a},
  {32'hc4b8eecd, 32'hc186ee76, 32'hc2a4dd7d},
  {32'h4466689a, 32'hc308862a, 32'hc26d391d},
  {32'h42985ed0, 32'hc3f8cb72, 32'hc3815c0f},
  {32'h44153576, 32'hc3c46e05, 32'hc2fb97ba},
  {32'hc509d490, 32'hc38ba792, 32'hc2855399},
  {32'h43870035, 32'h42557efb, 32'h409221e9},
  {32'hc4ecfc1f, 32'hc268cde4, 32'hc11de627},
  {32'h448a6253, 32'hc34de720, 32'h431315ad},
  {32'hc4f04186, 32'hc2a02b12, 32'hc3945cb1},
  {32'h447d39b0, 32'hc3872ca0, 32'hc4135ea5},
  {32'hc502aaa0, 32'hc28ca3be, 32'hc30831b8},
  {32'hc25e57b8, 32'hc34f272c, 32'h44013642},
  {32'hc4f0f8cf, 32'hc331ceaf, 32'h438e21bc},
  {32'h448ccf8a, 32'h4248567c, 32'h41b4f0a0},
  {32'hc4f2e1e2, 32'hc26cdb9f, 32'hc3416280},
  {32'h44063137, 32'hc05bd05a, 32'h4237020a},
  {32'hc2d8c758, 32'hc3469d5e, 32'h424fcd3e},
  {32'h44ece5c9, 32'h43b3b982, 32'h41a29752},
  {32'hc50a0482, 32'hc328d54d, 32'h43a3af0c},
  {32'h44590eac, 32'h423a467c, 32'h4364e7a4},
  {32'hc395e8b9, 32'h432a5a8f, 32'hc3822dc5},
  {32'h44ffa70c, 32'h42b83137, 32'hc30417ce},
  {32'hc472af7a, 32'h439eac2e, 32'h4365c8cf},
  {32'h44d0b598, 32'h437fc110, 32'hc2e5b9a1},
  {32'hc50b1b36, 32'h43b0344d, 32'hc2adab12},
  {32'h43f92200, 32'hc204c94c, 32'h433273f4},
  {32'hc4f21d62, 32'h424586b8, 32'h431d0653},
  {32'h44cb3551, 32'h4301a946, 32'hc2a00b2e},
  {32'hc2b975f0, 32'hc30ad7fa, 32'h4264ac06},
  {32'h44c5c7f5, 32'hc347dd25, 32'h42cbc6c1},
  {32'hc4f2ecf2, 32'hc29efd26, 32'h42b2e44f},
  {32'h44d50d1d, 32'h40430926, 32'hc38ea172},
  {32'hc44c283d, 32'h4326a8fa, 32'hc36075f3},
  {32'h44ff59a7, 32'hc2a5f184, 32'hc0eb6f82},
  {32'hc4d1b09d, 32'h42818e2c, 32'hc3704f09},
  {32'h45031d43, 32'h42fe7cfa, 32'h4300a9b0},
  {32'hc4d78c97, 32'h439d61b0, 32'hc2a25b8e},
  {32'h45018c47, 32'hc3b39f73, 32'h43863725},
  {32'hc4b22bc3, 32'h43c45ed8, 32'h43211a6a},
  {32'h44876835, 32'h4128239d, 32'h438f43e9},
  {32'hc46f315c, 32'h42103808, 32'hc1d323d5},
  {32'h44fd3b13, 32'hc3843ffc, 32'h42c065f8},
  {32'hc409bbce, 32'hc33d906c, 32'hc31078d5},
  {32'h4385d185, 32'h42be23d3, 32'h43502238},
  {32'hc17b1600, 32'hc37b1d0e, 32'hc234c9aa},
  {32'h449ebb20, 32'h42ad9f71, 32'h43057899},
  {32'hc4f93164, 32'h4342fff5, 32'h41ebecc5},
  {32'h43a2decd, 32'hc3d9db53, 32'h4289271c},
  {32'hc4a9dafa, 32'h43c10986, 32'h433cd65c},
  {32'h44c5d3b0, 32'hc32f9ca0, 32'h43545e70},
  {32'h43341ba0, 32'hc398f8aa, 32'h430d37b8},
  {32'h44c6890d, 32'hc3d0b35a, 32'hc2893e33},
  {32'hc486ecd8, 32'hc3972412, 32'hc2369219},
  {32'h44b6b447, 32'hc32e157a, 32'hc32049cc},
  {32'hc4fcc18e, 32'h42865952, 32'hc25c7829},
  {32'h44a531ad, 32'h438e92ba, 32'hc35725f0},
  {32'hc4bd438d, 32'hc0756f52, 32'hc30f28d0},
  {32'h43852102, 32'hc36ff29c, 32'hc29c2df0},
  {32'hc4abb769, 32'hc3b75dab, 32'hc39c0f65},
  {32'h43d55e5c, 32'hc307d517, 32'h4220287a},
  {32'hc4b00eb8, 32'hc3416a16, 32'h43475534},
  {32'h44673bd6, 32'h42ee740d, 32'hc3243c86},
  {32'hc48fd85f, 32'hc18adeec, 32'h42a9d64c},
  {32'h4496bbea, 32'h438bfdec, 32'hc32eff21},
  {32'hc4894380, 32'hc3836e05, 32'hc3497338},
  {32'h4285136c, 32'hc349485f, 32'hc33cf2eb},
  {32'hc35d5214, 32'h42ffac6f, 32'h3facb6e3},
  {32'h4458ec6d, 32'hc33b0104, 32'h415e9808},
  {32'hc3c43ab2, 32'h43646505, 32'h4074b170},
  {32'h4316b9d4, 32'h421b9253, 32'h4306c0d5},
  {32'hc4d69f74, 32'hc2d77291, 32'h432faf1b},
  {32'h44d60c0e, 32'h43835ada, 32'h4203df87},
  {32'hc432a6f9, 32'h43090c23, 32'h43006fd5},
  {32'h4481e13b, 32'h43e38710, 32'hc3c7521d},
  {32'hc4f56307, 32'h4107dde1, 32'h43921b39},
  {32'h45175c2c, 32'hc1ffd170, 32'h4366c16d},
  {32'hc51014ce, 32'h434e907c, 32'hc3ad564a},
  {32'h445012b8, 32'h43a3cac4, 32'hc3c5c5c2},
  {32'h43323ce0, 32'hc0054254, 32'h43400785},
  {32'h450e2db0, 32'h439228cb, 32'h42340621},
  {32'hc50928a7, 32'h43794bae, 32'h429bd19f},
  {32'h44f1786c, 32'h4363b879, 32'hc367dd98},
  {32'hc38b8212, 32'h43af487d, 32'hc2d0d755},
  {32'h4475dbc9, 32'hc1e991e9, 32'h436f85f9},
  {32'hc488547e, 32'hc2df91b8, 32'h437ecfd5},
  {32'h447dde1e, 32'h43231c29, 32'hc3d059cf},
  {32'hc4016452, 32'hc393fcf4, 32'h42f6667e},
  {32'h44fe6c9a, 32'h4252ac47, 32'h4324cd78},
  {32'hc42ccb3e, 32'h437a7979, 32'hc1c4d32e},
  {32'h44f7ad51, 32'h43afb2a4, 32'h42e6fadb},
  {32'hc50c0d9e, 32'hc2f61623, 32'h43012234},
  {32'h44122a2c, 32'hc30d9ab0, 32'h4334c750},
  {32'hc4275adc, 32'hc2fd2184, 32'hc3e78cc2},
  {32'h42debc10, 32'hc35b872d, 32'hc2f14336},
  {32'h421bcaae, 32'hc3afc937, 32'h43bf34b0},
  {32'h450f8eb2, 32'h432ac03c, 32'h42ee3b8b},
  {32'hc5006d72, 32'hc25648ae, 32'h42322439},
  {32'h44dae2ff, 32'hc321a143, 32'hc2d00472},
  {32'hc50398e4, 32'hc35bc861, 32'hc348504a},
  {32'h44f1c894, 32'h43b608ab, 32'hc37de42d},
  {32'hc4d40ece, 32'h428ce960, 32'hc176866c},
  {32'h43d37946, 32'h42581113, 32'h439cbfdd},
  {32'hc48e8161, 32'h440acce9, 32'hc33bd5bd},
  {32'h44aa4c08, 32'hc18ea604, 32'hc18d3a40},
  {32'hc39a9666, 32'hc2483105, 32'h411b6889},
  {32'h44febf6c, 32'hc384ae7c, 32'hc35ab1e4},
  {32'hc4bbfd71, 32'hc326efc5, 32'hc3c1cf5f},
  {32'h43843c63, 32'hc3548c0a, 32'h43899133},
  {32'hc45e7c3c, 32'h430080bf, 32'h42c4af68},
  {32'h449d4c0e, 32'h43695ac2, 32'h43967f6d},
  {32'hc4030ae4, 32'h4338cb45, 32'h4307b6a2},
  {32'h44dd69e0, 32'hc156c82e, 32'h43911fda},
  {32'hc42c73e0, 32'h43ae0a8a, 32'h40ed801b},
  {32'h449e4a23, 32'hc2b86f83, 32'h40c48933},
  {32'hc5211dde, 32'hc28b99d2, 32'h408e324e},
  {32'h448f2219, 32'hc2ebb672, 32'h3e3d0e88},
  {32'hc49daf0d, 32'h43bce65e, 32'hc34890ff},
  {32'h44a35d0e, 32'h41a5be44, 32'hc398919d},
  {32'hc50de2a2, 32'h4300164e, 32'hc3c62775},
  {32'h43757ae5, 32'h42d92829, 32'hc43ac353},
  {32'hc4f5ad40, 32'hc3169be3, 32'hc1c9cbbf},
  {32'h447237cc, 32'h43f1d323, 32'h42020abc},
  {32'hc5058a1f, 32'h439cf4e5, 32'hc3cb6826},
  {32'h451a4f0c, 32'hc2941f08, 32'hc202621e},
  {32'hc5012422, 32'h3f6642c0, 32'h4295dd95},
  {32'h44a35901, 32'hc2e62275, 32'hc286979f},
  {32'hc40b2148, 32'hc392f60f, 32'h430c0fb4},
  {32'h44bfafe8, 32'hc33f70e3, 32'hc38057be},
  {32'hc515abaf, 32'h422b03e2, 32'hc35164f4},
  {32'h44e9c774, 32'h42e12071, 32'h4313a847},
  {32'hc451bd2a, 32'hc3d2c51a, 32'h424b3446},
  {32'h44fab701, 32'h43b193c0, 32'hc2dd9963},
  {32'hc4c96494, 32'h44036ff4, 32'hc1b302e2},
  {32'h449eb6d2, 32'h4239c245, 32'hc20925d3},
  {32'hc5122588, 32'h429f8b75, 32'hc314c4fa},
  {32'h450ecf2f, 32'h42e50d18, 32'h4319f554},
  {32'hc4e3ba4c, 32'hbfeb2ee1, 32'h4353a4cb},
  {32'h44e0c1a6, 32'h42e3bfe1, 32'hc3209fc4},
  {32'hc4c2de3d, 32'h42f7a1aa, 32'h426d6454},
  {32'h44caf6f8, 32'h439d15db, 32'hc3862bbc},
  {32'hc50c6d24, 32'hc2f78f03, 32'h43b52d66},
  {32'h450daf27, 32'h432b3938, 32'hc283ef9f},
  {32'hc480042f, 32'h43340c65, 32'hc2b02088},
  {32'h43a5087d, 32'hc38a36ac, 32'hc31d5ccb},
  {32'hc4cd69cb, 32'h43490a94, 32'hc22663f5},
  {32'h438931a8, 32'hc2cdceb7, 32'hc3a58439},
  {32'hc44fd6a0, 32'h428077b2, 32'h42cda6ba},
  {32'h445dca1c, 32'hc3183269, 32'h430cc308},
  {32'hc46cc9c6, 32'h43a83088, 32'h43944c4a},
  {32'h445ad334, 32'hc396d087, 32'hc3555142},
  {32'hc4ddd91c, 32'hc336394e, 32'hc32d218f},
  {32'h44c334b8, 32'hc2cd9ccf, 32'hc2e5a13c},
  {32'hc49283a2, 32'h4167efa2, 32'hc33a50a7},
  {32'h44c54904, 32'hc3c3c689, 32'h42c7e334},
  {32'hc5229f90, 32'h4330f4c2, 32'h42acfd9f},
  {32'h451a2b02, 32'h43a0d351, 32'h43a2799a},
  {32'hc487a9cd, 32'hc1a7c34c, 32'h42e7cd48},
  {32'h43de3bd8, 32'h4321a519, 32'hc1a50ac2},
  {32'hc42db09e, 32'hc2e417fc, 32'hc32e9a62},
  {32'h43e0cd58, 32'h428c73e5, 32'h435ea893},
  {32'hc4a9eed8, 32'h43a9d5e1, 32'h43a0f862},
  {32'h45279d49, 32'h441c3b74, 32'hc3071a6e},
  {32'hc43fe218, 32'h4247dbdf, 32'hc3515c7c},
  {32'h44066b0a, 32'hc283ffb3, 32'h429f5e57},
  {32'hc4f7b386, 32'hc2400cd1, 32'h434a8ae9},
  {32'h450b623e, 32'h440627a9, 32'h4350de2a},
  {32'hc4f63740, 32'hc397badf, 32'h4329e6f2},
  {32'h450b4bd4, 32'hc34078a9, 32'hc2e92d6d},
  {32'hc4c864ed, 32'hc2f31c6a, 32'h44315bfb},
  {32'h447c0408, 32'hc4209531, 32'h4312280f},
  {32'hc5038219, 32'h4349184a, 32'hc41e114a},
  {32'h44f2a76b, 32'h43008802, 32'h431710f1},
  {32'hc4961da4, 32'h43a7bdb3, 32'h43496bdc},
  {32'h442afd28, 32'hc310ae91, 32'hc1c4aff6},
  {32'hc4b8f678, 32'hc301bf0b, 32'hc309d523},
  {32'h43491340, 32'hc2abc0c5, 32'h42ba1d00},
  {32'hc44e253b, 32'hc26c18ed, 32'h43a9fa59},
  {32'h4510a071, 32'h435098d3, 32'h4338c6a0},
  {32'hc4de284c, 32'h42142738, 32'h43635afe},
  {32'h43f40278, 32'hc1cc3eba, 32'hc29e5311},
  {32'hc4f7fccb, 32'hc2937ef0, 32'h4351ec59},
  {32'h44750b08, 32'hc3dcba6d, 32'hc3311e5e},
  {32'hc3df40c6, 32'hc368f3b6, 32'h4304bdf9},
  {32'h45190539, 32'hc1b48ad0, 32'hc30bd9f3},
  {32'hc41ae6ea, 32'h4391091d, 32'hc373b69b},
  {32'h44e87f5e, 32'hc2da05c3, 32'h40d9b346},
  {32'hc40a7aa4, 32'hc3919bfa, 32'h42150dd9},
  {32'h45153708, 32'hc2f6953d, 32'h436b65f4},
  {32'hc4867e63, 32'hc3303de2, 32'h42d1128a},
  {32'h44a44fbc, 32'h4232a692, 32'h4320f14b},
  {32'hc48a81e3, 32'hc35b3228, 32'h421797b8},
  {32'h4418d9d8, 32'h4263ea40, 32'h438bf8f7},
  {32'hc46c156c, 32'hc138ddf2, 32'hc3098a34},
  {32'h44cf5431, 32'hc22a67d7, 32'hc2c2e811},
  {32'hc3f385b2, 32'h4140f9e3, 32'hc3e1e8d6},
  {32'h43a058e4, 32'hc2dc22ff, 32'h41578e88},
  {32'hc4219adc, 32'hc29d5dd1, 32'hc2caf3f9},
  {32'h44591e27, 32'h43780a2d, 32'h42a9d119},
  {32'hc50775bf, 32'hc2ee7663, 32'h431e7e88},
  {32'h445b4eea, 32'h41f7424a, 32'hc3263e23},
  {32'hc515aad1, 32'hc3b0d7b6, 32'h438a767c},
  {32'h446a1d1c, 32'h42f41ab8, 32'hc26c917a},
  {32'hc30313c9, 32'hc3a75a61, 32'hc343e78c},
  {32'h44e955dd, 32'h42b4fffc, 32'hc302d8c3},
  {32'hc5133c7f, 32'hc1ff0b98, 32'hc272bffc},
  {32'h44eb30d4, 32'hc3053624, 32'h4272026c},
  {32'hc50457a1, 32'hc30d0cd3, 32'h43f1c7de},
  {32'h44b06090, 32'hc300e5a4, 32'hc3512490},
  {32'hc4f75306, 32'h42dd1420, 32'h43cea63d},
  {32'h44fad518, 32'h439cba18, 32'h41eb5466},
  {32'hc4bfac63, 32'hc31cea45, 32'h439245ef},
  {32'h44120429, 32'hc35047ca, 32'h433fa391},
  {32'hc47a3d8c, 32'h42d90962, 32'h42dcb5f2},
  {32'h44990dc6, 32'hc3088be6, 32'hc291a5e4},
  {32'hc35f83f8, 32'h43240588, 32'hc3362648},
  {32'h44cb108c, 32'hc1e86046, 32'h43850a8a},
  {32'hc497f6ec, 32'h435167b8, 32'hc26409dd},
  {32'h44689eb3, 32'hc243bdcc, 32'hc36a55e5},
  {32'hc50b0c13, 32'h43e936ec, 32'hc14439c6},
  {32'h44689e90, 32'h434bf33a, 32'h43ee4c3a},
  {32'hc50d9000, 32'h42ca4b03, 32'h438914f3},
  {32'h44e49f97, 32'h439a8412, 32'hc31278d7},
  {32'hc43df9d0, 32'hc31da050, 32'hc24f54da},
  {32'h44fd9a2e, 32'hc03e5048, 32'hc2ba7adf},
  {32'hc4cdef00, 32'hc2c8916e, 32'hc3016051},
  {32'h45343d5f, 32'h43e1f6cd, 32'hc2b26592},
  {32'hc501970d, 32'hc2c1eedb, 32'h406ecf66},
  {32'h44c5cef2, 32'hc376c585, 32'hc32859bf},
  {32'hc42646fe, 32'h438b625b, 32'h40ff5062},
  {32'h44e89bde, 32'h431cc6ab, 32'hc2e4ef50},
  {32'hc4d481d4, 32'h428911a7, 32'h41ec5d04},
  {32'h45145fe7, 32'hc2b71af2, 32'h438401d7},
  {32'hc48469e8, 32'hc30b3c40, 32'hc3b1ebf3},
  {32'h44421886, 32'hc320bc8e, 32'h42e4184c},
  {32'hc4032ae1, 32'h438631b6, 32'hc38c5c0e},
  {32'h451c5283, 32'hc26a209f, 32'h4312056d},
  {32'hc4a029c1, 32'h4340c1b7, 32'h437ba066},
  {32'h44fa20ac, 32'h436cb94a, 32'hc3568c53},
  {32'hc52f6449, 32'h3f8ef608, 32'h437a0a5f},
  {32'h44e09a48, 32'hc150d0b1, 32'h43aa9fb0},
  {32'hc3f3c379, 32'h420d3f1a, 32'hc3caee07},
  {32'h439e3ed0, 32'hc193f432, 32'hc297b4a5},
  {32'hc4f39c5b, 32'hc31ee892, 32'h43768bb1},
  {32'h44f5d977, 32'hc39ca33b, 32'hc3c9cc86},
  {32'hc471eb1a, 32'h4241b8b6, 32'h43188878},
  {32'h450d1abe, 32'hc2e5bd35, 32'h4305f464},
  {32'hc299ff80, 32'hc3dc11f6, 32'hc1110044},
  {32'h42faffa0, 32'hc3e9db98, 32'h43ea1f1b},
  {32'hc3531f07, 32'h43822d8c, 32'hc39c685f},
  {32'h44caf767, 32'hc3066392, 32'hc0f385b4},
  {32'hc48c89bc, 32'h43968372, 32'hc28ccb5c},
  {32'h42e83d48, 32'hc2f626d5, 32'hc1b276aa},
  {32'hc51828f6, 32'h43111cef, 32'h40586f86},
  {32'h448be522, 32'h433c6d99, 32'h43e4574e},
  {32'hc4895993, 32'hc1e52392, 32'hc3af1f27},
  {32'h44f7b785, 32'hc2860bf5, 32'h439dd83c},
  {32'hc511e9b9, 32'h42f3d5cd, 32'h416e4bd5},
  {32'h43c71fdc, 32'h4302e2af, 32'hc3409796},
  {32'hc3f6da30, 32'h42abd62f, 32'hbec90420},
  {32'h44e893a6, 32'hc31b3dee, 32'hc1811978},
  {32'hc4752184, 32'h42f52723, 32'hc30b56aa},
  {32'h443d7fb4, 32'h438eeed2, 32'hc2c833c1},
  {32'hc4acbedf, 32'h43a45e33, 32'h4266c4b6},
  {32'hc1daef40, 32'hc2a25821, 32'hc2f82cab},
  {32'hc4da05f7, 32'h4149f4c6, 32'hc343c7e5},
  {32'h44140561, 32'h43d48641, 32'h42a469b5},
  {32'hc4d6a4b1, 32'h43ab13c0, 32'hc3b9ca03},
  {32'h43f41969, 32'hc397eb6f, 32'h4390104a},
  {32'hc49207ee, 32'h435ff269, 32'h42fb0754},
  {32'h44eb1f6d, 32'h41bad9da, 32'h440d4a84},
  {32'hc2e16804, 32'hc307af82, 32'hc4008b00},
  {32'h44b32372, 32'hc2bc1281, 32'h4363f66b},
  {32'hc4ea8cf8, 32'h4388364c, 32'hc302aed3},
  {32'h44020116, 32'hc093b787, 32'h43743f58},
  {32'hc40ec7fa, 32'h42062c08, 32'h42981202},
  {32'h445f88d4, 32'h422a275c, 32'h434d5f8d},
  {32'hc4744417, 32'h42d3a4fa, 32'hc2ce6fe7},
  {32'h440669ba, 32'h43da6f2e, 32'hc2d0b2a3},
  {32'hc3a61ff7, 32'h4357de6a, 32'hc29c176a},
  {32'h45019f8c, 32'hc207b316, 32'hc1fe9f4c},
  {32'hc4e38634, 32'hc2716628, 32'hc3707416},
  {32'h4489fab8, 32'h4368a397, 32'h408c2f05},
  {32'hc4f4d90e, 32'hc40534b4, 32'hc2ae4581},
  {32'hc1e8e780, 32'hc2dddb54, 32'hc1be6990},
  {32'h44d7a5d2, 32'h41ab4827, 32'hc31c309f},
  {32'hc4dc1e2a, 32'hc2704227, 32'hc39ddbbd},
  {32'h4432ad0b, 32'hc3028a0a, 32'hc38614ad},
  {32'hc4ba62fd, 32'h43a370d8, 32'h42265942},
  {32'h447e6c97, 32'h43b87186, 32'h435d1ae0},
  {32'hc432b608, 32'h428fc866, 32'hc3bf29f4},
  {32'h44d8ac0a, 32'h435265c4, 32'hc2ab2268},
  {32'hc4c5c2bd, 32'hc37e598e, 32'h417880a2},
  {32'h44b2e1fd, 32'hc21150f0, 32'h436614fe},
  {32'hc398b63e, 32'hc2bdfa8e, 32'hc28de7a8},
  {32'h44624521, 32'hc1a1c25f, 32'h43703c3a},
  {32'hc49da84f, 32'hc35c730e, 32'hc2987de2},
  {32'h44674982, 32'h424acf89, 32'hc3b6c6fa},
  {32'hc43a2e70, 32'hc38c9b99, 32'hc38b502c},
  {32'h438a2759, 32'h43d302f8, 32'h43848c81},
  {32'hc4744f4c, 32'h42109b50, 32'h432deb48},
  {32'h44f5e4b3, 32'hc3b03cc4, 32'hc1d818d8},
  {32'hc48dad4f, 32'h42d2d1c8, 32'hc2e60d67},
  {32'h4505a584, 32'h43a0bf6a, 32'h42f7c0e9},
  {32'hc3f6e1dc, 32'h43548fda, 32'hc2863296},
  {32'h4496f80d, 32'hc2c1acc0, 32'h42ef7daf},
  {32'hc41f5bec, 32'hc0d4d39c, 32'hc0d88bcc},
  {32'h444bb7ac, 32'h428b4543, 32'hc22c9488},
  {32'hc49c19eb, 32'h4307fcc6, 32'hc3a49269},
  {32'h43b0a4c8, 32'hc3829477, 32'h4341ab6d},
  {32'hc4e4465e, 32'hc2b15de6, 32'h438b98ba},
  {32'h4357ad40, 32'hc282bd6d, 32'h42fe745e},
  {32'hc3ca4390, 32'h432e93be, 32'hc4095a7b},
  {32'h43aa1e1f, 32'h432e6a96, 32'h43293055},
  {32'hc2dfcd20, 32'hc1ea69ca, 32'hc3a99c91},
  {32'h4391bfe4, 32'h4226dfd2, 32'h4426109c},
  {32'hc3f67c00, 32'hc304200e, 32'h42c3415c},
  {32'h43eb6680, 32'hc261bf26, 32'hc2a02a0a},
  {32'hc4c1f3d4, 32'h42ecc5de, 32'hc3c7f952},
  {32'h43d2d0e4, 32'hc380712a, 32'h41f41562},
  {32'hc3901ffa, 32'h431a28bf, 32'hc32be2b9},
  {32'h43799e50, 32'hc37279c4, 32'hbf107d68},
  {32'hc4184542, 32'hc2f4463e, 32'h430f689e},
  {32'h43d25640, 32'h4348c952, 32'hc20c575a},
  {32'hc406184d, 32'h41ff5e64, 32'hc3d49323},
  {32'h43df85f6, 32'hc284d0bc, 32'h42c29845},
  {32'hc41618b3, 32'hc3884dfd, 32'h431e7bc7},
  {32'h449167d7, 32'h431d7cb4, 32'hc396be70},
  {32'hc48d6b4a, 32'hc2ef79b2, 32'hc2242af8},
  {32'h442073c0, 32'h43edd80d, 32'h43a751f5},
  {32'hc4dc90fb, 32'h43bf0a33, 32'h42f7b257},
  {32'h44e08bdc, 32'hc301a1ea, 32'h42c23187},
  {32'hc4ca5a88, 32'hc40d54db, 32'hc2ffd847},
  {32'h44f94130, 32'h42293cbe, 32'hc36c0c6b},
  {32'hc4a379ee, 32'hc30446ca, 32'hc37e0f26},
  {32'hc1d89c80, 32'h43b8051a, 32'hc301e413},
  {32'hc4fa1368, 32'h41d70d06, 32'hc3244708},
  {32'h44b042c7, 32'h42c4519a, 32'h424210ed},
  {32'hc4c10f90, 32'hc1d4613e, 32'hc321096e},
  {32'h44b2d975, 32'hc3d5e284, 32'hc3b85a54},
  {32'hc43fefd4, 32'h439e9fb1, 32'hc3354994},
  {32'h44719ed4, 32'hc1064952, 32'hc2e11ca3},
  {32'hc443c3b4, 32'hc3ed3b90, 32'hc36c5b65},
  {32'h450e4ac4, 32'h439993b2, 32'h43cb23a0},
  {32'hc4bd0743, 32'h437fb238, 32'h42df8c8e},
  {32'h44dfa12f, 32'hc39dc26e, 32'h40c523f8},
  {32'hc414b7ec, 32'h42ee4b5a, 32'hc3094bca},
  {32'h450a34c9, 32'hc4113632, 32'h4136e538},
  {32'hc342e720, 32'h4391139d, 32'h423b6efa},
  {32'h44c6d804, 32'h4231e5ad, 32'h4358b193},
  {32'hc4dc105a, 32'h428cdb45, 32'h42a1765b},
  {32'h444402e2, 32'h430c6039, 32'hc39d3e4e},
  {32'hc4f4e6fc, 32'h420efd4e, 32'h41fd78ce},
  {32'h44010cb8, 32'hc30d40d7, 32'hc2496c0d},
  {32'hc39cd24a, 32'h43757bb8, 32'h428ba7f5},
  {32'h44ef4bdf, 32'h4378330c, 32'h4313e9de},
  {32'hc36ed79c, 32'h43366d7a, 32'hc3f92b9e},
  {32'h42b281e0, 32'h42a963d3, 32'hc18f0bf8},
  {32'hc504c377, 32'hc2a696a9, 32'h438f4bc6},
  {32'h43d6538a, 32'h43ef12ea, 32'h437f88b1},
  {32'hc4bdbb53, 32'hc2a5ad95, 32'h4217134e},
  {32'h44965bd3, 32'h426361c3, 32'hc0c1955a},
  {32'hc48fdaea, 32'h432d4d1e, 32'h434e9201},
  {32'h4513e311, 32'h4301936d, 32'h42f271f3},
  {32'hc4d4971a, 32'h436be3ff, 32'hc320a9dc},
  {32'h441e9bac, 32'h43244d42, 32'hc18f5934},
  {32'hc4518178, 32'h4381e2c7, 32'h41881d27},
  {32'h43e0f7b8, 32'h434a85fe, 32'hc3321fc3},
  {32'hc48d47ea, 32'h42de99fe, 32'h4371b6a1},
  {32'h443d3a32, 32'hc2659ff6, 32'h433320a6},
  {32'hc4a80280, 32'h42d57a88, 32'hc2de80c4},
  {32'h450d191c, 32'h43e1b472, 32'hc33d15a8},
  {32'hc2f81220, 32'h42c62c9c, 32'h43abd766},
  {32'h4500b703, 32'hc3d959dd, 32'hc34a2762},
  {32'hc4da6d74, 32'h43134cde, 32'h425fa35d},
  {32'h42ac9874, 32'h42eb88df, 32'hc261baa4},
  {32'hc2afa880, 32'h43d1868a, 32'h4299aef3},
  {32'h43363430, 32'hc2c94e92, 32'h439b9c7b},
  {32'hc4e459f0, 32'h434d0bd3, 32'h4361aff5},
  {32'h4512eba9, 32'hc3acd421, 32'hc11414ff},
  {32'hc49a1b02, 32'h43af731f, 32'h431ec0cf},
  {32'h42a88394, 32'hc35e8b27, 32'hc322c65f},
  {32'hc423f754, 32'h4259a89a, 32'h42c3860a},
  {32'h449afa7c, 32'hc418ee50, 32'h43937491},
  {32'hc3f4832e, 32'h43663234, 32'h41fa96fa},
  {32'h451c4ddb, 32'h4338f2b2, 32'hc28425e7},
  {32'hc4fb9e75, 32'h4138269d, 32'h43b09b4f},
  {32'h44cc0ad1, 32'hc28111d0, 32'h4322e2ad},
  {32'hc404bcd4, 32'h437e32e2, 32'h439893b9},
  {32'h44a013cd, 32'h4244375e, 32'hc2fa82e7},
  {32'hc3788ef0, 32'hc3651d9d, 32'h43abf3f9},
  {32'h4504a184, 32'h427fdba0, 32'hc382fb9a},
  {32'hc4fa2d57, 32'h4377ec8d, 32'h438be6ac},
  {32'h43fcd29d, 32'h43428ea6, 32'h43925b20},
  {32'hc50c62bb, 32'h436353d2, 32'hc302c6aa},
  {32'h44152a04, 32'h4209b9b9, 32'h428e66ac},
  {32'hc50d61a5, 32'h4395424c, 32'h436ae7a0},
  {32'h4484608d, 32'hc13cd9e0, 32'hc181fcae},
  {32'hc4e6b160, 32'hc3505e9b, 32'hc2e8b3ab},
  {32'h44b3df26, 32'hc3dfd03c, 32'hc4591b6e},
  {32'hc45c1460, 32'hc28af4d7, 32'h44012395},
  {32'h44d7ed82, 32'hc36105ca, 32'hc28c8db5},
  {32'hc3f3f37a, 32'hc386f5b9, 32'hc347274c},
  {32'h4513f96e, 32'h42138380, 32'hc2ced942},
  {32'hc4ef8c29, 32'hc2baf2f2, 32'hc30a1584},
  {32'h44e8ff96, 32'h42d14568, 32'h42d76fe4},
  {32'hc4502462, 32'h4295f408, 32'h43228334},
  {32'h44ca8622, 32'hc237d6a3, 32'h4340a253},
  {32'hc5014d1c, 32'hc3b2f23c, 32'h43b5625d},
  {32'h44b18d5d, 32'hc237601a, 32'h435a293a},
  {32'hc4cec336, 32'h4261c391, 32'h4394ea37},
  {32'hc2856958, 32'h433f82c2, 32'hc3071486},
  {32'h43048fab, 32'h42324c16, 32'h42df9ced},
  {32'h4484aaa7, 32'hc2ab6097, 32'h41cfab0e},
  {32'hc40f1204, 32'h436010b6, 32'h4171b9ce},
  {32'h450de6f6, 32'hc37ae564, 32'h444c1756},
  {32'hc495ae8b, 32'hc2bfbf9f, 32'hc2b815ce},
  {32'h44d0bc8e, 32'hc22238ef, 32'hc359a4c1},
  {32'hc4bfbf7c, 32'hc2f49059, 32'h439797ee},
  {32'h4508267b, 32'h4245520e, 32'hc30765ec},
  {32'hc3338980, 32'h427bf86e, 32'h431ce8e8},
  {32'h44011bd8, 32'h43886bd4, 32'hc35e2727},
  {32'hc44b5dea, 32'h43acc4b1, 32'h4391e308},
  {32'h4481404c, 32'h42958bad, 32'h4287337f},
  {32'hc47b3514, 32'h43bc689c, 32'h429fc68a},
  {32'h44e91d0e, 32'hc31b42a5, 32'h42059424},
  {32'h41ff1ad7, 32'h437683ca, 32'h4384d4a0},
  {32'h44df79cc, 32'hc3933fad, 32'h43655442},
  {32'hc4cb4c79, 32'h434eb608, 32'hc2d5773b},
  {32'h449b2fd1, 32'h434736a3, 32'hc19204b7},
  {32'hc4a575d7, 32'h422b4d74, 32'h43c78317},
  {32'h4488d02a, 32'h4392018d, 32'hc421ccb4},
  {32'hc423094d, 32'h44378cba, 32'hc1decb47},
  {32'h44c55f62, 32'hc3688b30, 32'h4371c4a4},
  {32'hc443599a, 32'h43203e16, 32'hc338bfd1},
  {32'h44cd0532, 32'h42cd184a, 32'hc137db24},
  {32'hc4948ba4, 32'hc35a54c7, 32'h4266f92e},
  {32'h4494f180, 32'h406e1279, 32'h42285930},
  {32'hc3b577aa, 32'h42c58751, 32'hc20ba955},
  {32'h44f8832c, 32'hc34885f2, 32'hc34ee316},
  {32'hc4b1309a, 32'hc28d3630, 32'hc2fd2e31},
  {32'h44ad87d3, 32'hc15cb38e, 32'hc1683f7e},
  {32'hc47541a6, 32'hc1810b92, 32'h40a40386},
  {32'h42de55a0, 32'h4297c53b, 32'h42c59c59},
  {32'hc4c20acf, 32'hc39b0133, 32'h4274f8a2},
  {32'h44e3e1d4, 32'h435ed581, 32'h43a69b34},
  {32'hc3908570, 32'h43347ff1, 32'hc37fe726},
  {32'h44fceaba, 32'h434b93fb, 32'h412485b9},
  {32'hc3b3356a, 32'hc2350533, 32'hc1a93a7f},
  {32'h450b50ba, 32'h42d96460, 32'h43804cc6},
  {32'hc4c014d6, 32'h4346580c, 32'h438b8254},
  {32'h44d4de52, 32'hc405d5fe, 32'hc358c983},
  {32'hc3e8f888, 32'hc27f88a6, 32'hc31904af},
  {32'h449a89dc, 32'h4425c921, 32'h42d3a559},
  {32'hc39cf41e, 32'h43ff73ba, 32'h4269ffab},
  {32'h443935a4, 32'h42f1f374, 32'hc36e1848},
  {32'hc42b04a8, 32'h42e2c803, 32'h43375ed3},
  {32'h44f460f2, 32'hc38a39e5, 32'hc3620ce7},
  {32'hc462a869, 32'hc2ac9730, 32'hc3963fcb},
  {32'h44d3f117, 32'hc3bb9a4c, 32'h43faf60e},
  {32'hc4a0e8a8, 32'h4358f2da, 32'hc336dc16},
  {32'h45003ca6, 32'hc340a62f, 32'h43b73a0a},
  {32'hc4bfc40a, 32'hc33cd6a1, 32'h4187e802},
  {32'h450f0d60, 32'h41d00838, 32'hc340302b},
  {32'hc42ae60a, 32'h428eaa2b, 32'h439228f2},
  {32'h44e75631, 32'hc37f16e1, 32'hc4404d92},
  {32'h42c903c6, 32'h4241c327, 32'h439f31b5},
  {32'h44c5672e, 32'h43c9abae, 32'hc28622f6},
  {32'hc49c72a0, 32'hc0dd6af2, 32'hc2d4c4a2},
  {32'h44c5a6d2, 32'hc25d8dba, 32'h4343da6a},
  {32'hc4eb4686, 32'h4300ce5a, 32'h431762a7},
  {32'h444b3810, 32'hc3139e77, 32'hc3164697},
  {32'hc4ac7617, 32'hc00fd6c0, 32'h4293f09e},
  {32'h44d31d28, 32'hc404d55c, 32'hc20081a8},
  {32'hc4b7ce12, 32'h4393c995, 32'h4408830d},
  {32'h44e16e16, 32'h4336f54f, 32'h420ab804},
  {32'hc50067bd, 32'hc30aadd7, 32'hc2e2435e},
  {32'h44d6d76d, 32'hc3748016, 32'h4353e377},
  {32'hc4c7812a, 32'h43b81163, 32'hc19b2ea4},
  {32'h452482d2, 32'hc3600ef3, 32'hc3372bdd},
  {32'hc4267294, 32'h43617504, 32'h43c92507},
  {32'h44d4c253, 32'hc3aa956e, 32'h4287b4b0},
  {32'hc4f2e574, 32'h4312d8f3, 32'h440fb941},
  {32'h44afad21, 32'hc2611a2c, 32'h4352a575},
  {32'hc50d8790, 32'h40eb39b4, 32'hc28bf25f},
  {32'h4437ac84, 32'h43772680, 32'h42a75469},
  {32'hc4d3aaeb, 32'hc3101ea5, 32'h42bbbc61},
  {32'h44106bc8, 32'hc2375847, 32'h432033b7},
  {32'hc47d50e0, 32'hc1baa2ee, 32'h43621895},
  {32'h450d1a8d, 32'h42da44ec, 32'h424cb945},
  {32'hc4af3065, 32'h428c563f, 32'h43308be7},
  {32'h445c36ee, 32'h43af0224, 32'hc2642445},
  {32'hc49778f9, 32'h4257a439, 32'hc314a53d},
  {32'h44f03a98, 32'hc2b54811, 32'h422f11ea},
  {32'hc4f8d9d4, 32'hc25b5932, 32'h4317c39f},
  {32'h4406754c, 32'hc4202286, 32'hc28727c0},
  {32'hc500552f, 32'hc253067a, 32'h427baaf4},
  {32'hc2851218, 32'hc32d00ee, 32'hc34d54b2},
  {32'hc4411904, 32'h43dbf7d0, 32'hc1d7774c},
  {32'h44ea3274, 32'h430495cd, 32'h4290f1b5},
  {32'hc50fe36e, 32'h42ab9fa3, 32'h42c95819},
  {32'h43174230, 32'h4115c4d0, 32'h4319fe73},
  {32'hc3bf1fd8, 32'h40d5fdb0, 32'h428b4c0f},
  {32'h4406a306, 32'hc359d6ba, 32'h42effd96},
  {32'h41b15800, 32'hc0680100, 32'h42604350},
  {32'h44e5b3ff, 32'h42cb3040, 32'hc1ec6788},
  {32'hc4920fea, 32'hc36c0cbb, 32'h3faf1270},
  {32'h431f5878, 32'hc2c2e815, 32'hc307b37f},
  {32'hc3a41c98, 32'h42e5945e, 32'h41bb6f2e},
  {32'h45119021, 32'h430cb127, 32'h436bab97},
  {32'h43836f30, 32'hc35a09d1, 32'hc34c0b5c},
  {32'h438ac230, 32'hc387e310, 32'h43b22498},
  {32'hc48b6188, 32'h439044fb, 32'h42102736},
  {32'h4481d077, 32'hc4036605, 32'hc34a5e79},
  {32'hc5044bb4, 32'h429f0db2, 32'hc2d56973},
  {32'h4513ee54, 32'hc298a12d, 32'hc30d3ac2},
  {32'hc4f1cd3c, 32'h42e98eb6, 32'h43562887},
  {32'h44f18561, 32'hc3f37654, 32'h430790d4},
  {32'hc50aa14c, 32'hbec27008, 32'hc1ddf100},
  {32'h4430fe18, 32'hc1da6a75, 32'hc30ba310},
  {32'h42d67bc0, 32'h4332683e, 32'h431cfa00},
  {32'h44bdab81, 32'hc29f3fb5, 32'hc2c9dc3d},
  {32'hc4e95caf, 32'hc28d34f7, 32'h43232f94},
  {32'h444a8c58, 32'hc324e579, 32'hc3728ccc},
  {32'hc2a6acfe, 32'hc28193bf, 32'h43a96db0},
  {32'h44db4a8b, 32'h432d15e0, 32'hc16a74d5},
  {32'h43e6dbf4, 32'h4067371e, 32'hc3916aee},
  {32'h42fa3c40, 32'h43318902, 32'h42e3afc8},
  {32'hc4e987d3, 32'h4315beb9, 32'hc313cb8f},
  {32'h44ea04d9, 32'h40f5c7a4, 32'h43a854af},
  {32'hc47927af, 32'h440c10d3, 32'h423a8377},
  {32'h44d6f55c, 32'h4255e074, 32'hc3a8a18c},
  {32'hc4da40e6, 32'hc27c1460, 32'hc3859734},
  {32'h450d691a, 32'hc3962678, 32'h42053aec},
  {32'hc3081280, 32'h41e51293, 32'hc3934b89},
  {32'h44526c87, 32'hc31cab33, 32'h4348b2cb},
  {32'hc483bb36, 32'hc31ad02e, 32'hc3512dbd},
  {32'h44f674b9, 32'hc260136e, 32'hc36cafab},
  {32'hc24ca7d2, 32'hc3b580cc, 32'hc254edce},
  {32'h45020eb1, 32'hc33a696c, 32'hc236508d},
  {32'hc50079e7, 32'hc1ff5669, 32'hc35348a6},
  {32'h43474f1a, 32'hc18814fc, 32'hc397632f},
  {32'hc50fe9c4, 32'hc3c8f88e, 32'h41ab84e4},
  {32'h4217fb80, 32'hc1b02a12, 32'h4330961a},
  {32'hc51cea94, 32'hc3857810, 32'hc1de0bd9},
  {32'h44e3fd5f, 32'h42c13bea, 32'hc3c9ce1e},
  {32'hc4d89690, 32'hc3541c4d, 32'h432b4c1a},
  {32'h442865bc, 32'h42bbfd72, 32'h43838346},
  {32'hc50d49ac, 32'hc316ff40, 32'hc35257ea},
  {32'h44ef62a4, 32'hc38db1ee, 32'hc2bce61e},
  {32'hc3e49c62, 32'h41384c84, 32'hc3112df5},
  {32'h44d2b2ba, 32'h4389c975, 32'h412ca666},
  {32'hc4798568, 32'h431d66ec, 32'hc2c5af74},
  {32'h4499ca28, 32'hc29ff9af, 32'h434dae2c},
  {32'hc49695f0, 32'h42fe1448, 32'h43894ab8},
  {32'h44eb7ac0, 32'hc3907b20, 32'h4309d8de},
  {32'hc503f8fe, 32'hc26f56a4, 32'hc37b2a03},
  {32'h44861caa, 32'hc3857a8e, 32'h41ff89d7},
  {32'hc4b83f74, 32'h431a7d0c, 32'h433d2956},
  {32'h4490fbc8, 32'hc21140f0, 32'h43975f5c},
  {32'hc40c2c96, 32'h43abffe7, 32'hc26c1436},
  {32'h444fb51c, 32'hc1c3c98c, 32'h42cfacfe},
  {32'hc38f90b0, 32'hc3a25ca2, 32'hc3091f0a},
  {32'h44808880, 32'h412464b8, 32'h421153e6},
  {32'hc497d20c, 32'hc2e5eff4, 32'hc2a6f493},
  {32'h44ba7e68, 32'hc2e53157, 32'hc3433574},
  {32'hc4c98af1, 32'h408033f4, 32'hc18fb27a},
  {32'h444bf265, 32'hc3f9c0e4, 32'hc2d6bba7},
  {32'hc4fe35dc, 32'hc206e7bd, 32'h43b550ac},
  {32'h449007fc, 32'h438f5b62, 32'hc1e2886d},
  {32'hc4ebda15, 32'h432052eb, 32'h436323e9},
  {32'h44cb9c8c, 32'hc380638d, 32'hc31fffd5},
  {32'hc34d2e2b, 32'h4263a7f3, 32'hc29e11db},
  {32'h43d8f942, 32'h421bacf7, 32'h42f3d65f},
  {32'hc48a319d, 32'hc2802944, 32'h434e5a49},
  {32'h450caa0c, 32'h43364618, 32'h41b8bfee},
  {32'hc512e16c, 32'h4375a9c0, 32'h43d3969f},
  {32'h450903a1, 32'h438042f8, 32'hc36419a8},
  {32'hc4baff94, 32'h422806aa, 32'hc3920e07},
  {32'h43815ba0, 32'hc34e319d, 32'hc2fcdfb0},
  {32'hc495a825, 32'h43b5a660, 32'h431bd977},
  {32'h43861cb0, 32'h431d530a, 32'h43861ce0},
  {32'hc44abaa6, 32'hc28a8284, 32'h43c41a5d},
  {32'h45105fec, 32'hc1dd9cff, 32'hc3853e20},
  {32'hc4791827, 32'h438b539e, 32'h42c54e3d},
  {32'h449fb799, 32'h432bd9b1, 32'h41ce0275},
  {32'hc4604018, 32'h439d937b, 32'hc33b8056},
  {32'h4519f3b9, 32'h42df0910, 32'hc2ba246b},
  {32'hc46d5968, 32'h42bc84e5, 32'hc30147e8},
  {32'h44f3bbda, 32'h42314724, 32'hc34baf60},
  {32'hc4a55517, 32'hc287c6ce, 32'hc4192118},
  {32'h43caf8c8, 32'h4300e47e, 32'hc2faf87a},
  {32'hc4d5b5dc, 32'h42735f97, 32'hc29a767e},
  {32'h44c529e5, 32'hc2d0240b, 32'h44028ef7},
  {32'hc38f0e96, 32'h40af44d0, 32'h429bd35e},
  {32'h438eb7bc, 32'hc3b5bd84, 32'h42d8807c},
  {32'hc3c25528, 32'h43542e5d, 32'h436c23f3},
  {32'h44e323d7, 32'hc370a4d9, 32'h4315ee4e},
  {32'hc4490484, 32'h420129e8, 32'h41628bbd},
  {32'h44e6dd70, 32'h433aeee4, 32'hc30deebd},
  {32'hc405a4be, 32'h439e2d89, 32'hc3481e70},
  {32'h44759f70, 32'h426338aa, 32'h43f625d5},
  {32'hc3662060, 32'hc318f704, 32'hc2bc2734},
  {32'h4311f08e, 32'h42cba1c2, 32'hc34ae8d1},
  {32'hc2f18e30, 32'hc38e9ca0, 32'hc15d41a9},
  {32'h4495fa96, 32'h43e72d98, 32'hc2ee05c1},
  {32'hc4e6c252, 32'h418925c9, 32'h42700db8},
  {32'h44f8e0fe, 32'hc1ca1a8e, 32'h437884a4},
  {32'hc50854ee, 32'hc3154e24, 32'h4352fda9},
  {32'h45183fea, 32'hc2a5c087, 32'hc3192b9e},
  {32'hc500ed2a, 32'hc3a36af5, 32'hc27d25f3},
  {32'h44fc3a5a, 32'h441d0a2f, 32'hc2aa60bd},
  {32'hc355cb00, 32'h420c4376, 32'h439e50cf},
  {32'h44c01e1d, 32'h43574626, 32'h42c0a2f3},
  {32'hc4d0109e, 32'hc383701e, 32'hc354c406},
  {32'h44ce13e2, 32'h42593c8a, 32'hc3c9d270},
  {32'hc433b714, 32'h441a464e, 32'hc2ab6759},
  {32'h450603fb, 32'h41e6325e, 32'hc3734a45},
  {32'hc4b62b87, 32'hc19bd3f2, 32'hc34d5af2},
  {32'h44fe05fd, 32'hc3118bb3, 32'h427e4f3b},
  {32'hc4fc5084, 32'h425e2377, 32'hc315e92b},
  {32'h4516a3c9, 32'hc3221845, 32'hc2e80239},
  {32'hc444d70c, 32'h430dac6f, 32'h42613f24},
  {32'h44c3bee8, 32'h440f4b32, 32'hc07b4a2b},
  {32'hc43cb408, 32'h43615fb4, 32'h41f37bdc},
  {32'hc21b8700, 32'h42785e1f, 32'hc3855f7b},
  {32'hc4b3ddb8, 32'h436c333a, 32'h43df5158},
  {32'h44005378, 32'h430c4b6d, 32'hc3465a9f},
  {32'hc42b4c1f, 32'hc3a79af0, 32'h4385869a},
  {32'h44e0a0f2, 32'h43622038, 32'hc2fb30f9},
  {32'hc294da18, 32'h436c2b57, 32'hc3977d12},
  {32'h44b3d57b, 32'h43043770, 32'hc395ddf9},
  {32'hc4b6cb94, 32'h430d08c0, 32'hc3a6ac66},
  {32'h4437166c, 32'hc1f1fab3, 32'h4243534b},
  {32'hc5107411, 32'hc284b716, 32'h43ac940b},
  {32'h44a09912, 32'h4320e009, 32'hc302f288},
  {32'hc4e49a67, 32'h4348b0c5, 32'h4361d03c},
  {32'h44a9c2c6, 32'h3fc4934e, 32'hc1b0d31f},
  {32'hc42debc6, 32'h43915d5b, 32'h431cd84a},
  {32'h44f1cd26, 32'h42a41764, 32'hc22cf0ad},
  {32'hc44af4a6, 32'h440d7b87, 32'hc2ece9ce},
  {32'h43b531e2, 32'hc393febb, 32'h42aa6345},
  {32'hc396fa48, 32'h4296027d, 32'h430c55fa},
  {32'h44ec87b8, 32'h42762fad, 32'hc354a78d},
  {32'hc3a85f1b, 32'h4363ff80, 32'h42e35ecb},
  {32'h4485c490, 32'hc3a37318, 32'hc35892e7},
  {32'hc246fdb0, 32'hc337a759, 32'hc2a257df},
  {32'h41595b80, 32'h41d15c50, 32'h43f2e3aa},
  {32'hc28d3110, 32'hc23dc61e, 32'hc28bdd44},
  {32'h43bbb9a0, 32'h4363c2da, 32'h43962e86},
  {32'hc3b6fff8, 32'hc3aaf093, 32'h43bd0ecc},
  {32'h445e3e19, 32'h4259bcf2, 32'hc190f61b},
  {32'hc518fa16, 32'h43266aec, 32'hc38372ca},
  {32'h44d1943b, 32'h429e44e2, 32'h43c4be7c},
  {32'hc49fdb70, 32'hc2f4a345, 32'hc2970157},
  {32'h43e0a760, 32'hc182acc2, 32'hc1bac55b},
  {32'hc4b85de3, 32'h43062848, 32'h43131d69},
  {32'h448cbf86, 32'h43439120, 32'hc3569b47},
  {32'hc4fb45d2, 32'h42d1acd3, 32'hc2c0caa5},
  {32'h448f8274, 32'hc2cda583, 32'hc273d2cf},
  {32'hc3ee1dae, 32'hc2f9eaba, 32'h426f91b8},
  {32'h44bd4603, 32'hc37533ff, 32'hc356d212},
  {32'hc46ef83c, 32'hc3e72147, 32'hc2fba065},
  {32'h44f854a3, 32'h44186bb8, 32'hc2bf143e},
  {32'hc4ada67a, 32'hc2963e3b, 32'hc3b7006b},
  {32'h43993592, 32'hc2dc935a, 32'hc2abd4b8},
  {32'hc391ef53, 32'hc29dc214, 32'hc186579b},
  {32'h44b6c76a, 32'hc2ce4377, 32'hc152539f},
  {32'hc4d92447, 32'h424029e2, 32'h43b36bb4},
  {32'h437698c0, 32'hc286a805, 32'hc313407f},
  {32'hc40d4df6, 32'hc305cda5, 32'hc3416ec5},
  {32'h4503d837, 32'hc34b5798, 32'h42880d81},
  {32'hc40c9499, 32'h40051caa, 32'hc35f039d},
  {32'h448f8b85, 32'hc294578e, 32'h4385b7ce},
  {32'hc31b2199, 32'h428d2d0c, 32'hc2d5fd73},
  {32'h446410f8, 32'hc36b8b6b, 32'hc0acbd60},
  {32'hc4929d5e, 32'h41ae7419, 32'hc1c920a6},
  {32'h44aa55ec, 32'hc25b2dae, 32'h43452a4e},
  {32'hc35685e8, 32'h42174654, 32'h43970763},
  {32'h44b31b8a, 32'hc3c6b831, 32'h424b56d9},
  {32'hc50fc35e, 32'h42091830, 32'h43eba645},
  {32'h44f2a4fc, 32'h43913cdd, 32'hc2d72511},
  {32'hc39c5eac, 32'h43661441, 32'hc20a35a4},
  {32'h449f0a6e, 32'h42f64175, 32'h4041fe14},
  {32'hc4c6b848, 32'h427fb48e, 32'hc2b91bb4},
  {32'h44d67c69, 32'hc3940ad1, 32'h4236e093},
  {32'hc4a553c8, 32'hc1b48c9b, 32'h43c0e6b9},
  {32'h450c0e0d, 32'h439cc92f, 32'hc3122771},
  {32'h4103dba8, 32'hc3782e1d, 32'h41051fff},
  {32'h451aab12, 32'h430a5e45, 32'h41919643},
  {32'hc4f791da, 32'h435fe0f7, 32'hc289abe7},
  {32'h44ac923e, 32'hc33d8172, 32'hc124cb10},
  {32'hc4cd6082, 32'h43b9433f, 32'h43185bed},
  {32'h441f7aa0, 32'h42272ecc, 32'hc34d2775},
  {32'hc50b3eee, 32'h434e79de, 32'h43fbd16b},
  {32'h44cf2350, 32'h412dc618, 32'hc2d30e2c},
  {32'hc4b882f6, 32'h434572d3, 32'hc33714d9},
  {32'h44b30367, 32'h433e5ae5, 32'h4414cf65},
  {32'hc51e5a1c, 32'hc322b11e, 32'h43b39028},
  {32'h43abcea2, 32'h43ead11f, 32'h422035f7},
  {32'hc503c658, 32'h41ac4890, 32'h42438f58},
  {32'h4509fa20, 32'h42b6de44, 32'hc372231e},
  {32'hc4b0d1b2, 32'hc3baeaeb, 32'h43e35fe8},
  {32'h44a63abd, 32'hc2b832b0, 32'hc2d1769f},
  {32'hc4ec140f, 32'hc0abb670, 32'h4360fcb2},
  {32'h446a0b26, 32'h4320ddbf, 32'h439884b8},
  {32'hc3aab02f, 32'hc309ae5a, 32'h43c0f424},
  {32'hc2aa4da0, 32'h43d9f1e0, 32'h43c48720},
  {32'hc4bf8fa2, 32'hc329479c, 32'h43abbdc5},
  {32'h442fff43, 32'hc219fc00, 32'hc3a8cf7b},
  {32'hc43df1d2, 32'hc23eaca8, 32'h434ba548},
  {32'h44afaa98, 32'hc3aeff4b, 32'hc262e697},
  {32'hc4fafecb, 32'hc3a755f4, 32'hc363ce00},
  {32'h44c2c1d9, 32'hc2e567c4, 32'h4293ab49},
  {32'hc4d94602, 32'h427063ed, 32'hc2e87523},
  {32'h4458e834, 32'h41257068, 32'hc2a58cc1},
  {32'h44fd3eff, 32'h4347085a, 32'hc2be12c7},
  {32'hc418184b, 32'hc295ae85, 32'hc3883f0c},
  {32'h441c8dfb, 32'h43bd2f58, 32'hc2c9e598},
  {32'hc4bcf958, 32'hc334c0d8, 32'h443f86a8},
  {32'h44d6e57c, 32'h42f7c3e0, 32'h428e668b},
  {32'hc3c75b46, 32'h44215251, 32'h43366296},
  {32'h448dfbf4, 32'h43971eee, 32'hc30f4607},
  {32'hc4f6e49c, 32'h43ec8483, 32'h42ed7b50},
  {32'h448b6ce7, 32'hc22426a6, 32'hc3340294},
  {32'hc4bf5baa, 32'h431a2082, 32'h433c7aba},
  {32'h44be96de, 32'h43584ea4, 32'hc3026562},
  {32'hc40272ce, 32'hc33a2063, 32'h42d1c71b},
  {32'h45174bd8, 32'h4324ec5b, 32'hc2a8221e},
  {32'hc4b43545, 32'hc1dedf5e, 32'hc30f08a1},
  {32'h44f10250, 32'hc214937c, 32'hc29df377},
  {32'hc483bdcc, 32'h4399c526, 32'hc40dc2ff},
  {32'h4471c43d, 32'h439ce0b7, 32'hc3c775b5},
  {32'hc4f832c9, 32'hc3773e90, 32'h42dede8b},
  {32'h44a6f89e, 32'hc320df1b, 32'hc33cedc0},
  {32'hc4e2d0d2, 32'h420d5733, 32'h43cddb53},
  {32'hc2d5b2c8, 32'h4358ffe4, 32'hc389adbd},
  {32'hc40e2d1c, 32'hc3968faa, 32'h42de30e1},
  {32'h44ebb200, 32'h432b239a, 32'hc2ff15c7},
  {32'h43d87710, 32'h43904af3, 32'h42cdd929},
  {32'h43834948, 32'h4362176c, 32'hc3c44098},
  {32'hc485eabf, 32'h42b6831c, 32'h42046ba6},
  {32'h45188240, 32'hc3ac69f4, 32'hc318d7ef},
  {32'hc496f9a5, 32'h427c8da9, 32'hc038bd7e},
  {32'h44b71b4d, 32'h43e96616, 32'hc363a29f},
  {32'hc4db8d28, 32'hc252ccb3, 32'h4396d02f},
  {32'h44b10453, 32'h4300d1ca, 32'hc36eb5a0},
  {32'hc39f1aa0, 32'h4397afc6, 32'h434eb35d},
  {32'h44ae2729, 32'hc311320d, 32'h42db2364},
  {32'hc4390a50, 32'h43d63f05, 32'hc2bac551},
  {32'h433f84f6, 32'hc299b3cd, 32'hc3c17533},
  {32'hc50ceabb, 32'h4237d42b, 32'h41595ead},
  {32'h43a8c468, 32'h43a0adbb, 32'h43419be9},
  {32'hc419a961, 32'h4392a50c, 32'hc3f62754},
  {32'h448b3cc8, 32'h42a774fa, 32'h430b6749},
  {32'hc4f4181f, 32'h43a0e0fc, 32'h430e8dcf},
  {32'h44386ecf, 32'hc3685b5a, 32'h415bf349},
  {32'hc3c65084, 32'h436ff39c, 32'h424d89c3},
  {32'h45041585, 32'h41b283ad, 32'h43862f09},
  {32'hc4b1adbd, 32'hc2b16978, 32'h43613cec},
  {32'h44ef2f90, 32'hc3147379, 32'hc313dbe0},
  {32'hc495a183, 32'h425c863a, 32'hc356961b},
  {32'h45113061, 32'h4031ce10, 32'h43404250},
  {32'hc3634e20, 32'hc3d47214, 32'hc2dcf8ec},
  {32'h447b0588, 32'h42f684a0, 32'hc2a585e5},
  {32'hc487b6c6, 32'h4206fec4, 32'h434ce6a0},
  {32'h4210b528, 32'h41e34336, 32'hc3674ca3},
  {32'hc33b8778, 32'h4328b3a4, 32'hc290de49},
  {32'h44a2b43c, 32'h426a0ac4, 32'hc3c84fc4},
  {32'hc4bd40ba, 32'h41dc9d44, 32'hc3a0e2d0},
  {32'h433d3574, 32'hc196bdc2, 32'hc2ea8cdb},
  {32'hc4db710a, 32'h4313c7ff, 32'hc39b4e74},
  {32'h440ddc70, 32'h437c8f02, 32'hc21915de},
  {32'hc4a8c2d2, 32'hc370e451, 32'h4258887b},
  {32'h433b0b00, 32'hc3483ae4, 32'hc201df87},
  {32'hc5120d05, 32'hc2ba7562, 32'hc3708eb8},
  {32'h435d8450, 32'h43f0f5a7, 32'hc31e09cb},
  {32'hc35fd070, 32'h425440ba, 32'h43606bbd},
  {32'hc2ca3520, 32'hc32090bf, 32'hc301cea4},
  {32'hc4a07377, 32'hc3ff2105, 32'hc2691eb5},
  {32'h448a979b, 32'h421a7481, 32'h43e035ff},
  {32'hc482c49e, 32'hc327919f, 32'hc35f0562},
  {32'h44e3c512, 32'h42284b7d, 32'hc2faad36},
  {32'hc3a9bdb0, 32'hc34de242, 32'hc28b1f46},
  {32'h44df1493, 32'hc3eded9d, 32'h432cd5de},
  {32'hc417efd8, 32'h41316ea0, 32'hc289ea7e},
  {32'h4352f248, 32'h4282982e, 32'hc3e54121},
  {32'hc50a4311, 32'h428e737e, 32'hc3308f43},
  {32'h444052a2, 32'hc3718638, 32'h44079e3c},
  {32'hc4a7d834, 32'hbfe90462, 32'h4377855f},
  {32'h43ccb34c, 32'h43453e12, 32'h43384524},
  {32'hc399f5d0, 32'h4344c754, 32'h4370e9b3},
  {32'h43fd742c, 32'h42e37c93, 32'hc10b5973},
  {32'hc4da5d0d, 32'h42979d9b, 32'h42a20fd2},
  {32'h44a09bf8, 32'hc3fd9ba8, 32'h43313d90},
  {32'hc4c1a520, 32'hc34bca91, 32'hc33764e2},
  {32'h44023815, 32'hc2b836a4, 32'h43284ead},
  {32'hc4f478e1, 32'h4311ff7e, 32'hc2ef6afe},
  {32'h450c3a12, 32'hc0663b7c, 32'hc34ef3b7},
  {32'hc49d2078, 32'h433633fa, 32'hc22236ae},
  {32'h44ff6039, 32'hc262e21f, 32'h42d3e226},
  {32'hc356cb0e, 32'hc19b9e24, 32'h4289dcff},
  {32'h42d54b84, 32'h43510af2, 32'hc32e9992},
  {32'hc4955fdf, 32'hc2c7c613, 32'hc3f66aa1},
  {32'h451aed10, 32'h43d5853e, 32'hc336f57a},
  {32'hc4106457, 32'h437fb7ca, 32'hc2eb5453},
  {32'h4484efe9, 32'hc38bcd86, 32'hc228ba91},
  {32'hc458014c, 32'hc2367c5b, 32'h432c8674},
  {32'h447f2473, 32'hc2fbe707, 32'h4289c91c},
  {32'hc386d230, 32'hc2e29145, 32'hc25feeb8},
  {32'h445d5602, 32'hc35fa07e, 32'h4310712e},
  {32'hc38e36b8, 32'h42abb2a8, 32'h431fb438},
  {32'h44a95aee, 32'hc2c2dde7, 32'h432ed133},
  {32'hc4ae327c, 32'h43b1c60a, 32'h43a7d406},
  {32'h43a01c64, 32'h43788266, 32'h430ff545},
  {32'hc3e1bec5, 32'hc3bfe525, 32'h431c3ae3},
  {32'h4490e142, 32'h43182c3a, 32'hbf7e8ac8},
  {32'hc41cb434, 32'hc3d38334, 32'hc2c60198},
  {32'h44f14b42, 32'hc24e4727, 32'h42ece43a},
  {32'hc4b38d62, 32'h4386fd77, 32'h415c81dc},
  {32'h44cc2306, 32'hc2b9db27, 32'hc38f2e9c},
  {32'hc4c64756, 32'hc3be7ae9, 32'hc2ecb38a},
  {32'h44e3f3fb, 32'hc31501ac, 32'hc3b07294},
  {32'hc2316e40, 32'hc31c08f6, 32'hc3abd77d},
  {32'h44c41306, 32'h436c76f0, 32'hc3debff9},
  {32'hc40795da, 32'hc35ac2f6, 32'hc2c4f40c},
  {32'h4513d713, 32'hc2aad73b, 32'h435b18b9},
  {32'hc4f10ae6, 32'h42a0813d, 32'h42a35a15},
  {32'h44d0666e, 32'hc1a91c7d, 32'h438206b8},
  {32'hc3929a76, 32'h43a0d3d3, 32'hc231d983},
  {32'h43b68629, 32'hc2a19358, 32'h40cdb200},
  {32'hc452af92, 32'hc224a21f, 32'hc0caa8d0},
  {32'h443c9560, 32'hc1c0a8e0, 32'hc39b7f05},
  {32'hc3fa1538, 32'hc1f5944d, 32'hc377b9ce},
  {32'h438b48d0, 32'h424ef196, 32'h431b49da},
  {32'hc5034b4f, 32'hc3269fd3, 32'h433cb50f},
  {32'h445ea540, 32'hc2341594, 32'hc337b4a0},
  {32'hc4f24c55, 32'hc36d9f38, 32'h43b78610},
  {32'h44d03c64, 32'h432065dc, 32'h42c2aca7},
  {32'hc316ef20, 32'hc37e4f12, 32'hc2d1aa8a},
  {32'h43cc9bb7, 32'h43825215, 32'h438995e6},
  {32'hc4026697, 32'h43d06ad9, 32'h438dbd37},
  {32'h43eb3a25, 32'hc2e153e1, 32'h41ad4c16},
  {32'hc4a9b296, 32'hc19b7a3e, 32'hc337ba0e},
  {32'h4537e59a, 32'h4357a2f1, 32'hc35488be},
  {32'hc43292ed, 32'h4379a1dd, 32'h439ba618},
  {32'h44c21e12, 32'h439813db, 32'hc26b2ad6},
  {32'hc41ffd4a, 32'h434c7cc7, 32'hc2d2955d},
  {32'h4408dfb1, 32'hc11239f7, 32'h438642e6},
  {32'hc48d3734, 32'h43c2894e, 32'h4259c495},
  {32'h441fd010, 32'h433edd3c, 32'hc23b27f1},
  {32'hc3c3c538, 32'hc3ac4327, 32'hc1b2e314},
  {32'h43c3ae7c, 32'hc2b94a66, 32'hc2a46996},
  {32'hc42955a6, 32'hc2ef98ce, 32'hc2d8864d},
  {32'h44d206bb, 32'h43c13d3f, 32'hc396cabb},
  {32'h426ef5d9, 32'h43ad29b5, 32'h428efa03},
  {32'h44e8e477, 32'hc38562f8, 32'h43700602},
  {32'hc428e803, 32'hc36c06d4, 32'hc3125fa5},
  {32'h44d9ecb2, 32'h43258293, 32'h42ef1476},
  {32'hc4b19dfe, 32'hc30eb123, 32'h413ef16b},
  {32'h436e748c, 32'h43cbbeb2, 32'h43c074f5},
  {32'hc437bf4a, 32'hc2875446, 32'h42887dac},
  {32'h4383da12, 32'h42e28f55, 32'hc2912d69},
  {32'hc4f710a2, 32'h4300abd9, 32'h41f49650},
  {32'h4501a2f6, 32'hc3002432, 32'h4233a4ed},
  {32'hc4ac93fc, 32'hc3abe651, 32'hc3fa5202},
  {32'h44af8070, 32'hc3141fb4, 32'hc2bf830b},
  {32'h42783d18, 32'hc2d6167a, 32'h42caecc9},
  {32'h44de3e55, 32'h4331a02d, 32'h4335695b},
  {32'hc4e0224a, 32'h4305c19b, 32'h4191e90d},
  {32'h4514ad12, 32'h43448ea9, 32'h42d706ae},
  {32'hc4c28340, 32'h4305462b, 32'h429557c8},
  {32'h43e0eaf8, 32'hc39060f6, 32'h42d7d221},
  {32'hc34605b6, 32'h42c65ad4, 32'h42010c2a},
  {32'h4406755d, 32'h42c8ace4, 32'hc322fde5},
  {32'hc45d4d23, 32'h435705ba, 32'hc3225310},
  {32'h447e9a65, 32'hc309627f, 32'h4413cc51},
  {32'hc4642609, 32'hc3ec9997, 32'hc3ef9246},
  {32'h44a9d3f7, 32'h42a4df2f, 32'h43ba2cd2},
  {32'hc3aba76e, 32'hc2e2f6f6, 32'hc36b9957},
  {32'h446c0fa8, 32'h42b2d058, 32'h41b45b43},
  {32'hc4fbef82, 32'h43b7699c, 32'h439cd52f},
  {32'h44bcc73d, 32'hc201e8dc, 32'h41688ab4},
  {32'hc47b8174, 32'hc2977c0c, 32'h437c0e80},
  {32'h45007b25, 32'h4303ff37, 32'hc15604c8},
  {32'hc4e90914, 32'h42f2d101, 32'h4393cfbf},
  {32'h449c7df0, 32'hc213df1c, 32'hc1d84b90},
  {32'hc42ee7cf, 32'h43b9135d, 32'hc297555b},
  {32'h45019d00, 32'hc31ff0fb, 32'h4309e9c7},
  {32'hc4abcc04, 32'h43b08da0, 32'h4177e09b},
  {32'h44fcb7ed, 32'hc265c15c, 32'h43675a98},
  {32'hc4e255d8, 32'h437a6d92, 32'hc37f2d9d},
  {32'h450e5eaa, 32'hc3a3c586, 32'h439efbbc},
  {32'hc43f4164, 32'hc2d36128, 32'h4368f084},
  {32'h44dc7a1e, 32'h42e19da4, 32'hc3ece2e4},
  {32'h434c0ea0, 32'hc3807b6e, 32'h4086ee15},
  {32'h444e0f92, 32'h4230744f, 32'hc38360e5},
  {32'hc457b41e, 32'h421f49f0, 32'h4271208c},
  {32'h438a443e, 32'hc32c994c, 32'hc3afb06c},
  {32'hc4b65041, 32'h43b392f3, 32'hc2b65145},
  {32'h44703820, 32'hc3993c2a, 32'hc33d41a3},
  {32'hc4b673ff, 32'hc2de4ada, 32'hc25995d3},
  {32'h43ca5858, 32'h42bc833b, 32'h423630f0},
  {32'hc389d5ac, 32'h41584340, 32'h428878d3},
  {32'h44e58055, 32'hc3262f5e, 32'hc11dba2a},
  {32'hc4b17b52, 32'hc362cf5e, 32'h43bd5eab},
  {32'h43c24690, 32'h4387dac7, 32'h43758351},
  {32'hc4c0a2f2, 32'h41428bd3, 32'hc2b4527c},
  {32'h44985b91, 32'h42855e21, 32'h431aca81},
  {32'hc4ab70c4, 32'h43933b73, 32'h436c73ec},
  {32'h440bf73f, 32'h4381fbfa, 32'h42f0df69},
  {32'hc4796620, 32'h429fa261, 32'hc32386e0},
  {32'h44b814bb, 32'h4204e6e0, 32'hc3783cf4},
  {32'hc3cd8672, 32'h431936ec, 32'h41767404},
  {32'h450f19b3, 32'h43f380d8, 32'h423c6df8},
  {32'hc3a4ed9a, 32'h41f249d4, 32'h4386f6ee},
  {32'h44cd65fc, 32'h43f84432, 32'hc29361ae},
  {32'hc4e0d36b, 32'hc28d1d32, 32'hc39ac861},
  {32'h4453c768, 32'hc1a9b96d, 32'hc2f3a232},
  {32'hc4a4e83b, 32'hc2a9d47e, 32'h43a34ba4},
  {32'h440bdb9c, 32'h43730d52, 32'hc187624d},
  {32'hc4889e5f, 32'hc2d613aa, 32'h427c26dc},
  {32'h450a8118, 32'hc38a63cf, 32'hc34b5a1b},
  {32'hc4dee869, 32'h43934774, 32'hc2c3f518},
  {32'h447a96a8, 32'hc38ee28f, 32'h42a4b515},
  {32'hc3b30b20, 32'h4203d839, 32'hc3e0b6c4},
  {32'h446e5684, 32'hc2b9c2d9, 32'h4427d7c3},
  {32'hc490f191, 32'h440272a2, 32'hc3b4d209},
  {32'h44955e01, 32'h434000c7, 32'h42b14507},
  {32'hc50635f4, 32'hc20f4e78, 32'h431c570b},
  {32'h44839eb2, 32'h4341947b, 32'hc33369e8},
  {32'hc4f9e849, 32'hc36e39f8, 32'hc3308770},
  {32'h43c2b280, 32'hc2ccba2a, 32'hc34fb53a},
  {32'h431f6d20, 32'h433c4517, 32'h441ee7bb},
  {32'h44d7c806, 32'hc3ae4cbb, 32'h4276bf94},
  {32'hc4b7dc7b, 32'h43a62230, 32'h43844124},
  {32'h450bed05, 32'h4334f109, 32'hc38b3745},
  {32'hc4d6d68a, 32'h43064e6a, 32'h422209f4},
  {32'h43d6c621, 32'hc2386d4e, 32'hc1a0bf4b},
  {32'hc2b5eca0, 32'h4295b566, 32'hc3ac5f08},
  {32'h45068fb4, 32'h4374057a, 32'hc3e39070},
  {32'hc3feff34, 32'h438b3aab, 32'h4287233f},
  {32'h45236f9d, 32'hc373b319, 32'hc3b2531d},
  {32'h428a6868, 32'h442023bb, 32'hc3066b12},
  {32'h42f7b430, 32'h43039f7f, 32'h42be16e8},
  {32'hc4dee1d5, 32'h428a72b9, 32'h43135826},
  {32'h44d2eba8, 32'hc32e1825, 32'h4356cb34},
  {32'hc504cbc8, 32'hc3250bd1, 32'hc2f2e328},
  {32'h44b92122, 32'h42cd0802, 32'h4388a5d4},
  {32'h42a51060, 32'hc2a3dcca, 32'h43354818},
  {32'h436b4d3e, 32'h439bae6d, 32'hc3506f78},
  {32'hc4667e71, 32'h42bf846f, 32'hc31e082b},
  {32'h43d09e5e, 32'hc28b7002, 32'h4297fbf5},
  {32'hc3fd1788, 32'h41f1a7be, 32'h42bb8e35},
  {32'h44930cb9, 32'h42f29120, 32'h43745de4},
  {32'hc4282b64, 32'hc299e5ef, 32'hc17ace7c},
  {32'h4490df80, 32'h42d0120b, 32'hc31e26f3},
  {32'hc462b99a, 32'h436778fb, 32'hc3c2fc85},
  {32'h44620e27, 32'h42b02b44, 32'h43661e4d},
  {32'hc40dfa80, 32'h42710cae, 32'h422e9788},
  {32'h44a7fd85, 32'hc3a7e461, 32'hc319d09a},
  {32'hc4c42520, 32'hc35e2ca0, 32'h4393f9c6},
  {32'h44d7bcdf, 32'h4355fc1b, 32'h434110a7},
  {32'hc4a638eb, 32'hc2800c71, 32'hc31d702d},
  {32'h447126e6, 32'hc26c1874, 32'h42954d44},
  {32'hc3db0be6, 32'hc2b5cc25, 32'h433cd315},
  {32'h4482015c, 32'h432207a4, 32'hc30e4f6b},
  {32'hc4ae0102, 32'h436dc9dd, 32'h434efb99},
  {32'h44845f14, 32'hc34f6100, 32'hc38123b0},
  {32'hc4e74d11, 32'h4308e815, 32'hc3a0eaec},
  {32'h44b66a09, 32'hc3042608, 32'h4327ed7a},
  {32'hc4fc0bde, 32'h434ef12e, 32'hc4020f95},
  {32'h4337aa98, 32'hc30b700e, 32'h422aa33a},
  {32'hc4ec948e, 32'h40f42550, 32'hc297dadb},
  {32'h44ade0fb, 32'h435e833a, 32'hc1f46d02},
  {32'hc3686802, 32'h434ed7b0, 32'h43c04167},
  {32'h44400c0c, 32'h43b3c4c3, 32'hc3115f29},
  {32'hc489aa3a, 32'h43a59257, 32'h433db086},
  {32'h4327b9a0, 32'hc3034ca6, 32'h438946d5},
  {32'hc4c5332f, 32'h42621da8, 32'hc28515e8},
  {32'h44f1167a, 32'hc343cf96, 32'hc2d584b7},
  {32'hc51a5e54, 32'hc351c8f0, 32'h422ea2dc},
  {32'h4501a4d0, 32'h42e09697, 32'hc3152596},
  {32'hc503e50f, 32'hc31099aa, 32'h42eac174},
  {32'h4404f9b6, 32'h4305ed6c, 32'hc3c109ca},
  {32'hc4aa8a15, 32'h432408ed, 32'hc33e1b61},
  {32'h43adf1ba, 32'h42b94cfe, 32'h4390eace},
  {32'hc4fb0f9b, 32'hc366b933, 32'hc2deab0e},
  {32'h446d6d92, 32'h42c1c0cc, 32'hc3832c5d},
  {32'hc4f9f9ca, 32'hc19ed057, 32'hc231cfbe},
  {32'h44c04d8c, 32'h43942a5b, 32'h42a7b611},
  {32'hc4955b4c, 32'h431a3403, 32'h434a3e8f},
  {32'h44951ece, 32'hc2061313, 32'h43364033},
  {32'hc4522c7f, 32'h43cc8e2d, 32'h4355a903},
  {32'h4337d380, 32'hc1eab230, 32'h43ae2b5b},
  {32'hc47250f4, 32'hc2867154, 32'h40bd6100},
  {32'h43b55c69, 32'hc28d9968, 32'hc28f1958},
  {32'hc4dcd19c, 32'hc276caf1, 32'hc2b6a5f1},
  {32'h4463792e, 32'h43405104, 32'h43964bd9},
  {32'hc4c8f74f, 32'hc1cf688c, 32'h40dc8e9a},
  {32'h4383e95c, 32'h4357e5c8, 32'h4398d781},
  {32'hc39b21da, 32'h433faa61, 32'h42f656dc},
  {32'h446a0f94, 32'hc2473633, 32'hc3c983ad},
  {32'h4332724c, 32'h41ef31de, 32'h425e24fb},
  {32'h445f5698, 32'hc07c6320, 32'hc37042d5},
  {32'hc46519aa, 32'hc1929272, 32'hc3e59e21},
  {32'h43286450, 32'h433b8e0c, 32'hc2382020},
  {32'h432503b0, 32'hc21c468e, 32'hc36fb14c},
  {32'h442a631a, 32'hc3d72ce8, 32'hc387c10a},
  {32'hc4bcfe09, 32'h43c95fd6, 32'hc32cbc7d},
  {32'h44dc1df0, 32'h42f13756, 32'hc3924c68},
  {32'hc5153063, 32'hc1725ffc, 32'h4374370a},
  {32'h4414e766, 32'hc3e79933, 32'h439ae815},
  {32'hc45c3026, 32'hc3b9d651, 32'h43fea063},
  {32'h4509f4de, 32'hc384bb99, 32'h3f640210},
  {32'hc4c7b032, 32'h430b6514, 32'h434190be},
  {32'h4516a9b8, 32'h420837dd, 32'h435a24e5},
  {32'hc4b3f97f, 32'h408c9fc2, 32'h437e993b},
  {32'h443d85ce, 32'h42bde485, 32'hc3424448},
  {32'hc50a6904, 32'hc3230621, 32'h43b9c201},
  {32'h440506aa, 32'h43d808ac, 32'hc12b089c},
  {32'hc43d66b2, 32'hc32c0e49, 32'h41cc41aa},
  {32'h4453bc71, 32'hc2e14239, 32'hc2f0feef},
  {32'hc4037728, 32'h4353643c, 32'hc3c2d91c},
  {32'h4443c305, 32'h4249cc2c, 32'h43bc012b},
  {32'hc502707a, 32'hc378e057, 32'hc366a46a},
  {32'h44f0aa22, 32'h437cdcad, 32'h431a7322},
  {32'hc507676d, 32'h439b7826, 32'h43fbaab3},
  {32'h44f4ab59, 32'h43bab18d, 32'h42d6f47e},
  {32'h43033488, 32'h43995680, 32'h42f6d601},
  {32'h448c2eb2, 32'h42d59687, 32'hc3551138},
  {32'hc4d7626d, 32'hc29aea30, 32'hc2aee9a3},
  {32'h4450d7bc, 32'h42ef811b, 32'hc310870e},
  {32'hc5011d5b, 32'hc31d9ebe, 32'h42001296},
  {32'h44609914, 32'h42e8ab90, 32'h43da60be},
  {32'hc40c81ce, 32'hc30b9c22, 32'hc20599d0},
  {32'h4499920b, 32'h43895324, 32'hc315daa4},
  {32'hc419dad0, 32'hc3913a50, 32'hc3f9bd86},
  {32'h42e20cc0, 32'h4383edde, 32'h43389c61},
  {32'hc3b7f718, 32'hc2dabfb6, 32'hc2d73ecb},
  {32'h44d31035, 32'hc285223e, 32'h431eca8a},
  {32'hc34ceb14, 32'h4320fd26, 32'hc1e69bf1},
  {32'h44bc399b, 32'h42c8eb33, 32'hc327a9f0},
  {32'hc43828b8, 32'h42931775, 32'hc3a26f0d},
  {32'h44124c3c, 32'h435258e9, 32'hc241d6df},
  {32'hc49a1042, 32'h42fddc5d, 32'h441d07f7},
  {32'h451cea1f, 32'h43766d04, 32'h4105ba54},
  {32'hc4f71bdd, 32'hc37df2f8, 32'h438fcd70},
  {32'h442c5b4a, 32'h4350711b, 32'hc3979f35},
  {32'h42794600, 32'h424a7649, 32'hc320f8e2},
  {32'h43d2f310, 32'h4357ecda, 32'hc3891696},
  {32'hc376cc40, 32'h42674dcd, 32'h4223fc34},
  {32'h45275a73, 32'hc3b333ba, 32'hc31696f4},
  {32'hc517c481, 32'h4368db9e, 32'hc3c9da74},
  {32'h449d88d8, 32'h43d6e61d, 32'h41fea687},
  {32'hc4c77373, 32'hc2168d30, 32'hc2a4cfdf},
  {32'h44973785, 32'h42c3f64e, 32'hc3000422},
  {32'hc510447d, 32'hc43b8490, 32'hc2dd9b1a},
  {32'h44e640c8, 32'h423ac77b, 32'h43e1df10},
  {32'hc4dc005e, 32'hc2765c33, 32'hc2ffc23d},
  {32'h43d49828, 32'hc35afd0f, 32'h41c1950a},
  {32'hc5076f98, 32'h423a6e85, 32'hc3152d62},
  {32'h44ce6827, 32'hc41c5b79, 32'hc34add40},
  {32'hc4d298e5, 32'h43138d70, 32'h425c27ac},
  {32'h44e7adce, 32'h3f3443f0, 32'hc20f9392},
  {32'hc47aa2da, 32'hc1e206d6, 32'h42ed8dcf},
  {32'h451ea3d3, 32'hc37d1da0, 32'h420a9ad9},
  {32'hc4c0552a, 32'h437353c8, 32'hc10f7bf5},
  {32'h43ad0ca0, 32'hc22d1f7b, 32'hc378dfc3},
  {32'hc46d8a8c, 32'hc295fe25, 32'hc2dfd89c},
  {32'h42871b3d, 32'h438287d4, 32'hc16336d5},
  {32'hc4ce7752, 32'hc0e8226c, 32'h43157353},
  {32'h44838538, 32'hc2c2480c, 32'h435b9bee},
  {32'hc42a369b, 32'hc395a271, 32'hc292c054},
  {32'h426c77d0, 32'h43a93ba2, 32'hc4046be6},
  {32'hc5194f83, 32'hc28b7f5a, 32'hc2090119},
  {32'h45056f9b, 32'hc3b3fe14, 32'hc2b2b1bd},
  {32'hc3f46937, 32'hc36d3b51, 32'hc2fafe25},
  {32'h4457021a, 32'h431798b7, 32'hc2ba65de},
  {32'hc4a753b6, 32'hc240ab04, 32'hc2d16d89},
  {32'h43817584, 32'hc2bfcec2, 32'h435e5670},
  {32'hc4bba649, 32'h43ee8619, 32'h428fd493},
  {32'h43052964, 32'hc394ae6f, 32'hc34c4889},
  {32'hc5394311, 32'hc28a1261, 32'hc2b0466e},
  {32'h441a4900, 32'hc2819d24, 32'hc32fb140},
  {32'hc410f5ee, 32'h42dcb608, 32'h437deeb0},
  {32'h450ac833, 32'hc38551e8, 32'hc26ff77c},
  {32'hc5055966, 32'hc375194a, 32'hc2470ada},
  {32'h449355f0, 32'hc3970838, 32'h40c6e33a},
  {32'hc4dcb793, 32'hc319bb3e, 32'hc3453ae9},
  {32'h447a9f5a, 32'hc32545c9, 32'h432c0fa0},
  {32'hc3d0b544, 32'hc31ae6d3, 32'h430441fc},
  {32'h44eb4ccc, 32'h434cd335, 32'h436a89ff},
  {32'hc4b3f283, 32'h429be1fd, 32'hc3a8202b},
  {32'h44d80080, 32'hc30e00b9, 32'h4286a1ee},
  {32'hc46680bc, 32'h4356ed9b, 32'h438e665c},
  {32'h43ef77d9, 32'hbfc32e7d, 32'hc30056d9},
  {32'hc4bf3cd2, 32'h42861d97, 32'h439656a0},
  {32'h442e4b70, 32'h42d3e13b, 32'h432016f7},
  {32'hc3416240, 32'h4131d889, 32'hc2fdbf87},
  {32'h44d9219c, 32'hc3302f38, 32'hc1b67420},
  {32'hc48f7476, 32'hc30c262d, 32'h40addc2f},
  {32'h450166d3, 32'hc275dabc, 32'h4290d323},
  {32'hc49c8533, 32'hc2ac0f99, 32'h43074936},
  {32'h44fce43a, 32'hc3f9a2e4, 32'hc38e4661},
  {32'hc512b7bb, 32'hc29023ae, 32'h417fd662},
  {32'h44b6e03e, 32'hc34cf27a, 32'h42ee05af},
  {32'hc5066245, 32'hc3c61105, 32'hc15d788a},
  {32'h44c3a624, 32'h41dcd77a, 32'hc17f7a3d},
  {32'hc49704bd, 32'h40d0f5ed, 32'hc19a1e8f},
  {32'h4462f498, 32'h4360d775, 32'h430e3993},
  {32'hc476d6c3, 32'h42e3f073, 32'hc356d7c8},
  {32'h44fdc0f3, 32'h435d842e, 32'hc045996e},
  {32'h4386e588, 32'hc3975e83, 32'hc359d3cf},
  {32'h44155aec, 32'hc2e1cbb4, 32'h3f57c6a0},
  {32'hc4437c5c, 32'hc0716af2, 32'hc4012c31},
  {32'h43ebd510, 32'h436cff3b, 32'h439d6386},
  {32'hc438c28a, 32'hc3e92dbf, 32'h438ad397},
  {32'hc30e9a5e, 32'hc3720a47, 32'h4176e45c},
  {32'h432905a8, 32'h42aeeb3f, 32'h4343edb4},
  {32'h44fcb53f, 32'h43709715, 32'h4315ed0a},
  {32'hc4071860, 32'hc30039ba, 32'hc3b9291a},
  {32'h4437e158, 32'h433d052d, 32'hc37ee6d0},
  {32'hc39c0cbc, 32'hc33f82c7, 32'hc37073ad},
  {32'h43b8e728, 32'h42426419, 32'h435e5dd2},
  {32'hc49799c5, 32'hc3094d2e, 32'hc352d1a0},
  {32'h44faa974, 32'h43193516, 32'h430abe5c},
  {32'hc389caa6, 32'hc2804f1a, 32'hc336088c},
  {32'h45103c8a, 32'hc10609ab, 32'hc2b8a15a},
  {32'hc40b03e0, 32'hc3275326, 32'h43c3e7b2},
  {32'h44040076, 32'h439dea17, 32'h4312548e},
  {32'hc4a30242, 32'hc33c0f19, 32'hc20751e4},
  {32'h4529bd03, 32'hc3526225, 32'hc40cb0c0},
  {32'hc48379b4, 32'hc3905543, 32'hc3bec6fa},
  {32'h43958268, 32'hc31f4359, 32'h42f4be40},
  {32'hc34376a8, 32'hc210ff1d, 32'hc3280159},
  {32'h43766b10, 32'h42b1e2c3, 32'h40036e80},
  {32'hc4b9edfc, 32'h42e8f4ee, 32'hc2f7e76a},
  {32'h44ac4edb, 32'hc3657cef, 32'h43237c7e},
  {32'hc4de2dae, 32'hc34e0fc8, 32'hc2b49a34},
  {32'h44bbdec1, 32'h4264dbb0, 32'h4387315e},
  {32'hc419b98c, 32'hc3306930, 32'hc3b6641d},
  {32'h44332284, 32'hc18cbe6c, 32'h43acdba4},
  {32'hc4f7fe11, 32'hc3c83cc4, 32'h42875b68},
  {32'h444e62f8, 32'h43cf224b, 32'h425287d8},
  {32'hc16e15ba, 32'hc3affe0c, 32'hc21fe604},
  {32'h44f54c5f, 32'h42352cff, 32'h4388bc3b},
  {32'hc36877e8, 32'hc4242057, 32'hc2156b04},
  {32'hc434755a, 32'hc2a49b88, 32'hc2ed7d86},
  {32'h44526a5b, 32'h43425363, 32'h439b760e},
  {32'hc3de8800, 32'hc2f926cd, 32'hc3cc2938},
  {32'h44e34256, 32'h3cb5a350, 32'hc2ca9c1a},
  {32'hc39658b0, 32'hc37c2dac, 32'hc3b5dc3d},
  {32'h44261efc, 32'hc32edfd7, 32'h43d4bede},
  {32'hc523d6cc, 32'h43b43df7, 32'hc393c977},
  {32'h45048f9e, 32'h430f1d55, 32'hc2153aea},
  {32'hc4c4850b, 32'hc324bab9, 32'hc32164ea},
  {32'h449c77d7, 32'hc1aee5a4, 32'h4342b50e},
  {32'hc362b6a8, 32'hc2bef984, 32'h42872357},
  {32'h44e81d70, 32'hc3781917, 32'hc2c4363b},
  {32'hc488bfa2, 32'h43941ade, 32'hc3602c2d},
  {32'h442efebc, 32'hc39c26b9, 32'h4320fd13},
  {32'hc4f1f25a, 32'h4363e115, 32'hc36528e1},
  {32'h44a78436, 32'h42d18f67, 32'hc345071c},
  {32'hc4546cf8, 32'hc1030689, 32'hc2ec674e},
  {32'h449da807, 32'h431f2074, 32'hc2b5b914},
  {32'hc4bbbfc4, 32'h430bce64, 32'hc36bd7c2},
  {32'h44ea42f0, 32'hc33dfdbf, 32'h42278e26},
  {32'hc4b1a0ec, 32'hc385f725, 32'hc22912a1},
  {32'h44b9febc, 32'hc2e7d3cf, 32'h4336e285},
  {32'hc4c930c8, 32'hc39e12bb, 32'hc35d053e},
  {32'h44539e23, 32'hc2981458, 32'h432a8686},
  {32'hc4f8c3d1, 32'h42538b4f, 32'h42e462d2},
  {32'hc3189554, 32'hc386763a, 32'hc189c18e},
  {32'hc3554d68, 32'hc29a70fd, 32'h4188cc08},
  {32'h4420732c, 32'hc3602be2, 32'h438f819e},
  {32'hc4a3abf6, 32'hc2add0bb, 32'hc4309f18},
  {32'h45015232, 32'hc348e0fe, 32'hc22a3203},
  {32'hc4f1e7f7, 32'hc1c3332e, 32'hc38af47f},
  {32'h440fcc72, 32'h423ddd4e, 32'hc34b5299},
  {32'hc4667ec6, 32'h4256e5d8, 32'h407d4626},
  {32'h43c5a94a, 32'hc1426710, 32'h413d2a45},
  {32'hc43bbb34, 32'hc1602e9c, 32'h425fbb7b},
  {32'h43d7ef36, 32'h42bd9f78, 32'hc2ad593e},
  {32'hc504f97e, 32'hc19e61b2, 32'h42b5b00c},
  {32'h44f930b9, 32'h4382f045, 32'h42fed229},
  {32'hc4533e3c, 32'hc3c26264, 32'h42ed8122},
  {32'h449fda52, 32'h4300051e, 32'h4299efd5},
  {32'h40eed400, 32'hc17f4380, 32'hc1d9719c},
  {32'h4472e208, 32'h430e01f7, 32'h431ef313},
  {32'hc4c24052, 32'h43168607, 32'hc333ed1a},
  {32'h449ab6e5, 32'h42c90230, 32'h434d39fd},
  {32'hc41b6e2c, 32'h42b2b524, 32'h421fbf9e},
  {32'h450a86d5, 32'hc1ed69dd, 32'h436f5b32},
  {32'h436cbad8, 32'hc294c4da, 32'hc352aa7d},
  {32'h448e7fea, 32'h43abd6e5, 32'h43d37f95},
  {32'hc3f66618, 32'h43905491, 32'hc34ca9a8},
  {32'h44bf26bc, 32'hc3966e5e, 32'hc392d9ea},
  {32'hc328114e, 32'h42f461f3, 32'hc380224e},
  {32'h4400b661, 32'h41086886, 32'h40f9ecb0},
  {32'hc4e9ed47, 32'h4212b5b8, 32'hc35148eb},
  {32'h4501af29, 32'h43918d03, 32'hc2ad4c1c},
  {32'hc5045870, 32'hc2d5721c, 32'h422dca0e},
  {32'h4395c964, 32'h4312e902, 32'hc11703c6},
  {32'hc4a40c3d, 32'hc38b05a2, 32'h4297c3fc},
  {32'h45088686, 32'hc3423c81, 32'hc3a95ac2},
  {32'hc5012342, 32'hc20fe9e8, 32'hc3756572},
  {32'h4394c69b, 32'hc323d2d8, 32'hc31696a9},
  {32'hc43d1cdc, 32'hc11edb9e, 32'hc349e56a},
  {32'h44edfc68, 32'hc22abbaf, 32'h43f0de21},
  {32'hc35e7b9c, 32'h4267d6c3, 32'hc2a6a41d},
  {32'h44b9f1d3, 32'h42facc12, 32'hc1eb7ce6},
  {32'hc504496a, 32'hc338e1b6, 32'h431c3b00},
  {32'h43840a92, 32'h4208e7ad, 32'h42f78386},
  {32'hc4f7144e, 32'h433a678f, 32'h4131478f},
  {32'hc20908e0, 32'hc1aa441a, 32'hc23d1968},
  {32'h43200aa0, 32'hc3050cb8, 32'hc3402e3f},
  {32'h44a1f027, 32'h438b16cc, 32'h43155a4d},
  {32'hc48be404, 32'hc31d0b82, 32'h43489286},
  {32'h450516c3, 32'hc3967ff1, 32'h429b72a9},
  {32'hc26c8320, 32'hc38d59fd, 32'h43cebc0e},
  {32'h43e78dd5, 32'hc28cd7d0, 32'h439f62f4},
  {32'hc4f3c6a8, 32'h4387c571, 32'hc16017a5},
  {32'h44fb2de7, 32'h4302bbe5, 32'hc27b4806},
  {32'hc4eef986, 32'hc3a396a1, 32'hc256245f},
  {32'h44e41d1b, 32'h42a88040, 32'hc369f1dd},
  {32'h422dde78, 32'hc29d8743, 32'h4318599b},
  {32'h4483cb4c, 32'h433b1ab6, 32'h439016cb},
  {32'h4383fc78, 32'hc34a29eb, 32'hc31b9d38},
  {32'h43b02f0e, 32'h436e5a96, 32'hc309c611},
  {32'hc4fe6476, 32'h41321600, 32'h4356d5df},
  {32'h44d8cebe, 32'hbf8c4ad9, 32'h43ca6c7b},
  {32'hc46483a4, 32'h434c14eb, 32'hc10b2708},
  {32'h4520fdd4, 32'h42e3602a, 32'h431e0b48},
  {32'hc49d9544, 32'h433af277, 32'hc2aea47f},
  {32'h44e48b69, 32'hc346fe9d, 32'hc3107a42},
  {32'hc487e7ae, 32'hc35666aa, 32'h430228ff},
  {32'h44fc9c7e, 32'h4330acac, 32'h43c5aa88},
  {32'hc4c46a66, 32'hc38a7597, 32'h43801f55},
  {32'h445b1502, 32'hc30d1033, 32'h4335ca72},
  {32'hc21cc880, 32'hc2349811, 32'h4271f70c},
  {32'h451ed545, 32'h42ca9b0e, 32'h43ecb727},
  {32'hc492d92e, 32'hbf9d4e88, 32'hc353d769},
  {32'h437b461d, 32'hc32485a6, 32'h438dfcb1},
  {32'hc47596f4, 32'h4385bd3d, 32'hc22956ec},
  {32'h44f57fd0, 32'h42dff36a, 32'hc1d59b32},
  {32'hc5003c82, 32'h42c3678b, 32'hc3858595},
  {32'h450f8710, 32'h4394d0a1, 32'h430f1005},
  {32'hc480070f, 32'h42697c92, 32'hc337879a},
  {32'h44a4f0d1, 32'h4284ff29, 32'hc2ff9bd0},
  {32'hc500da40, 32'h439abdd2, 32'hc207ace1},
  {32'h44432a22, 32'hc2c9a93f, 32'h42aa463b},
  {32'h435b18a8, 32'h4410cc11, 32'h434c0675},
  {32'h4482f604, 32'hc2acaecd, 32'hc29793b3},
  {32'hc4641a10, 32'h42ec0256, 32'h43643cc9},
  {32'h43b45380, 32'hc3abb87b, 32'h416ea2e8},
  {32'hc3622b30, 32'h414b9297, 32'h4113bbf0},
  {32'h44ae8aea, 32'hc1a2f8e9, 32'h4243d193},
  {32'hc3eb2ac8, 32'hc426443f, 32'h438ad773},
  {32'h43a10443, 32'hc3c9205c, 32'hc22e3d7d},
  {32'hc402e9a4, 32'hc2faf248, 32'h441af4e8},
  {32'hc38b4c6c, 32'hc396d4c9, 32'h4286f1df},
  {32'hc41db808, 32'hc3280384, 32'hc278312c},
  {32'h44bcd5c0, 32'hc328ffa2, 32'hc34288cb},
  {32'hc3b3275f, 32'hc11ceb65, 32'hc2d3f773},
  {32'h44a363d4, 32'hc3d88c3b, 32'h42e909d1},
  {32'hc2ad8b80, 32'hc3fd1b52, 32'hbfd70da0},
  {32'h42b6321c, 32'hc304df3c, 32'hc0aec9c2},
  {32'hc50ace82, 32'h42f8f975, 32'h435baa5b},
  {32'h45004ec6, 32'hc339ddd2, 32'hc383e495},
  {32'hc3233246, 32'h438a6b00, 32'h4304e449},
  {32'h442cee66, 32'hc3632b3d, 32'hc3c4ecce},
  {32'hc4e15c12, 32'h4315ea42, 32'hc3bd053f},
  {32'h4415277e, 32'h4392f632, 32'hc39a5d10},
  {32'hc4a4ebfb, 32'hc3b85fa1, 32'hc29288bc},
  {32'h44e120a2, 32'hc3d19f69, 32'hc315da4a},
  {32'h408b77a8, 32'hc3596224, 32'hc2f38314},
  {32'h4310eb90, 32'hc3428546, 32'hc37ec44f},
  {32'hc29eeae8, 32'hc266e53b, 32'hc3ae113a},
  {32'h45231763, 32'h439ed64e, 32'hc07041c0},
  {32'hc4300f4d, 32'h4375a5ae, 32'h4300ee24},
  {32'h44ae313e, 32'h43285b52, 32'h43138939},
  {32'hc43fce40, 32'h438f3681, 32'h3ffc5460},
  {32'h44f3b6fe, 32'h411eaa32, 32'hc244759b},
  {32'hc487a00f, 32'h43c65ca3, 32'h43630c78},
  {32'h44d2c426, 32'hc3817bf8, 32'h4360b425},
  {32'hc4a64f9d, 32'hc32c07a3, 32'hc34e4e40},
  {32'h4506aacc, 32'hc2631a21, 32'h43571c5a},
  {32'hc4b7ca54, 32'h4105a3ef, 32'h435adf9f},
  {32'h44d3e6c7, 32'hc2b0e2b2, 32'h413d9e0e},
  {32'hc445e1e8, 32'h4271b673, 32'h43366f55},
  {32'h4504da12, 32'hc360a7d9, 32'hc3a10c60},
  {32'hc4d34586, 32'h4322fb40, 32'h43354460},
  {32'h45037bf8, 32'h3f9492f1, 32'h439431b8},
  {32'hc4e7530a, 32'h4311a5b6, 32'hc3840ea4},
  {32'h44b3e615, 32'h41b90836, 32'hc3485500},
  {32'hc4486f78, 32'hc2d2e11f, 32'hc34b7365},
  {32'h44a4e0c7, 32'hc257a6bf, 32'h4203d08f},
  {32'hc3e2a772, 32'hc30113c7, 32'h4220e222},
  {32'h4507c5a8, 32'h42a9047a, 32'h43212c45},
  {32'hc4e31f34, 32'hc34c7a30, 32'hc16af239},
  {32'h442020ef, 32'h434a44b3, 32'hc30ac741},
  {32'hc506a346, 32'hc2cc5f8c, 32'hc2d6ac66},
  {32'h44785f4c, 32'h43d82d93, 32'h427a6e99},
  {32'h42dad1a0, 32'hc2eec0fe, 32'hc32e5180},
  {32'h44fda2cb, 32'h431351d3, 32'hc3ae45b0},
  {32'hc319e2c0, 32'hc3afb3e1, 32'hc359cef4},
  {32'h44efd5af, 32'hc2dac6fb, 32'h4314b492},
  {32'hc4cb2e8e, 32'h43668d4b, 32'h42ba8f83},
  {32'h439b6f30, 32'h42749131, 32'hc3a5606e},
  {32'hc435afba, 32'hc3731fe2, 32'hc2577be5},
  {32'h441d3f98, 32'hc327e9c2, 32'h41e4d44f},
  {32'hc49ef7d4, 32'h420153db, 32'hc21dadc9},
  {32'h44404d47, 32'h439accb8, 32'hc2f253a9},
  {32'hc4df5cc3, 32'hc362633a, 32'h43c314eb},
  {32'h442ebd03, 32'hc39530e2, 32'h4301675c},
  {32'hc38b8a00, 32'h42a87599, 32'h41e4a047},
  {32'h44edc777, 32'hc2c02068, 32'h430a6cd0},
  {32'hc3a48e08, 32'hc32cda8a, 32'hc3e20367},
  {32'h44e31ee7, 32'hc2f77350, 32'hc28f146c},
  {32'hc4d865c7, 32'h4384c759, 32'h42829553},
  {32'h43c3e7b2, 32'hc30722ee, 32'hc4007cdf},
  {32'hc45c8ea0, 32'h431c6e7d, 32'hc33986b3},
  {32'h44c685bd, 32'h43c59f2d, 32'h4194ddfd},
  {32'hc48430db, 32'h43d3bdde, 32'h4339297f},
  {32'h44034c58, 32'hc2c39459, 32'hc2e9a4a0},
  {32'hc4a442cb, 32'hc36a9891, 32'hc2b79514},
  {32'h4423ba38, 32'h4218a488, 32'hc3835ac2},
  {32'hc503ed4c, 32'hc30d14e7, 32'h4288dc7e},
  {32'h44484572, 32'hc44c41b1, 32'hc3dc3fef},
  {32'hc4957eb1, 32'h4369ccf3, 32'hc38fe672},
  {32'h43610750, 32'h4394fbca, 32'hc2e4722e},
  {32'hc39532d6, 32'hc3827c63, 32'hc2a140e8},
  {32'h440833b4, 32'h43000012, 32'h425441d6},
  {32'hc508de92, 32'h4286be81, 32'h438a8dd4},
  {32'h44bb7768, 32'hc394ae88, 32'hc3a65f1b},
  {32'hc4483f7a, 32'h42a62314, 32'hc31753eb},
  {32'h4368cfe8, 32'h4236b1a8, 32'hc3566508},
  {32'hc49139be, 32'hc34e0a76, 32'hc22ee41e},
  {32'h42e2ff20, 32'h4274047b, 32'hc2dd74bd},
  {32'hc463c19c, 32'hc3d676f5, 32'hc3a25e05},
  {32'h44d8efa6, 32'hc327c36c, 32'h43db9c61},
  {32'hc445a4dc, 32'hc272ec2b, 32'hc35a8a00},
  {32'h44b7348f, 32'h421cc5fd, 32'h42f12dce},
  {32'hc26eea87, 32'h41d1c1d0, 32'h440c8bed},
  {32'h449097ba, 32'h4217ac7a, 32'h42c69278},
  {32'hc4dc7d4a, 32'hc1b509e3, 32'h43c7def4},
  {32'h450c09dc, 32'hc223e21e, 32'h43a11358},
  {32'hc36dc790, 32'h420e8d53, 32'hc13bbf68},
  {32'h43f2cd3b, 32'hc37d70fc, 32'h42ab8781},
  {32'hc4ecab66, 32'hc2d961ed, 32'h43a02ff1},
  {32'h44a1a328, 32'hc3509a2b, 32'hc28f88c6},
  {32'hc4bee232, 32'hc345c50f, 32'h41e29eb8},
  {32'h44a859e8, 32'hc3599554, 32'hc304a7d0},
  {32'hc50e07ae, 32'h430e4b32, 32'hc3c14733},
  {32'h43c651ca, 32'h434fbd12, 32'hc39b9f94},
  {32'hc4622e91, 32'h429957ca, 32'h42c790f4},
  {32'h43cbcc02, 32'hc289cce7, 32'hc417ef4e},
  {32'hc47ab6a4, 32'h424936b1, 32'h43c70a08},
  {32'h44f818db, 32'h42b021f4, 32'h4188bf8e},
  {32'hc46674af, 32'h413b2488, 32'hc35119e4},
  {32'h4468009f, 32'hc2bd672e, 32'h410c1ef1},
  {32'hc51eb266, 32'h40df245e, 32'hc288e9aa},
  {32'h4509741a, 32'h40f8511c, 32'h418d9538},
  {32'hc4005fe4, 32'hc333bbb6, 32'hc37d4c27},
  {32'h44b9fabf, 32'hc21b3619, 32'hc27d355c},
  {32'hc3ea5ca8, 32'hc225f8da, 32'hc309996c},
  {32'h43a6c938, 32'h41e5ada8, 32'hc2c56123},
  {32'hc4374735, 32'hc2fc859b, 32'h41269bcb},
  {32'h4486a1d2, 32'h43008c6d, 32'hc22f373c},
  {32'hc507d829, 32'hc2052cf8, 32'hc2a5c869},
  {32'h448748e9, 32'hc3a03160, 32'h42ee9c44},
  {32'hc4eafb11, 32'hc2286b22, 32'hc3b8236f},
  {32'h44ca624d, 32'hc3cf3526, 32'h438e713c},
  {32'hc50709b8, 32'h423766ad, 32'hc38ed5b3},
  {32'h4489a892, 32'h42b01131, 32'hc290f6f9},
  {32'hc507b4cc, 32'hc21300a5, 32'hc35942e7},
  {32'h447bd50f, 32'hc3a40938, 32'h4203a744},
  {32'hc39e15f0, 32'h4322a8e3, 32'hc3098b44},
  {32'h44d6fc45, 32'h43a5b59f, 32'h43bd08dc},
  {32'hc4aeee00, 32'h4367e9eb, 32'h426c899e},
  {32'h44de4b65, 32'hc2cbb386, 32'hc30a5230},
  {32'hc496cf9e, 32'h43109da1, 32'h41ce6018},
  {32'h4459ec4e, 32'h42bce378, 32'h4195fe34},
  {32'hc4b291f3, 32'hc2bd9a44, 32'hc25fd454},
  {32'h44bb9c39, 32'hc3c14fae, 32'hc36af054},
  {32'hc4231247, 32'h42959407, 32'hc313b9f2},
  {32'h4360ff64, 32'hc310dbfd, 32'h43418efb},
  {32'hc464b7cc, 32'h43780608, 32'hc2cdab24},
  {32'h44cb1c2a, 32'h43087b6d, 32'hc3d95c6f},
  {32'hc34a7b74, 32'h42045a82, 32'hc2dfe54b},
  {32'h44946b01, 32'h4345f2b9, 32'hc2b4c45a},
  {32'hc50f2eaa, 32'hc32b1d27, 32'hc2e30fe2},
  {32'h43f4a510, 32'h43cd428c, 32'h428b68c1},
  {32'hc428a512, 32'hc2c8271f, 32'hc402d047},
  {32'h450ac11e, 32'hc402827a, 32'hc29c5627},
  {32'h4266d180, 32'hc30ef83f, 32'hc32a4d18},
  {32'h44c52e88, 32'h4304e54f, 32'h4354d44c},
  {32'hc4ef12e0, 32'h42c8fec0, 32'h43a2a474},
  {32'h4503a4e0, 32'h42dce29e, 32'hc309e3ab},
  {32'hc3268970, 32'hc400d654, 32'h4288b3c6},
  {32'h44967a55, 32'h4033f0a8, 32'hc309d7b9},
  {32'hc4d1427d, 32'hc27faaab, 32'h41f8e5f3},
  {32'h44d02098, 32'hc340d85d, 32'hc350bc1d},
  {32'hc4ea511a, 32'hc32d4f15, 32'hc2a98f28},
  {32'h44e11f52, 32'h4397b6e3, 32'h4337d689},
  {32'hc46b6652, 32'h439e9958, 32'hc39657aa},
  {32'h44c021f0, 32'h4232bd8e, 32'hc3433151},
  {32'hc4ae156e, 32'hc3c6ac96, 32'hc3d8032f},
  {32'h43e54f30, 32'h4232955b, 32'h40c91a1b},
  {32'hc442adc0, 32'hc3f08ac5, 32'hc3276ee1},
  {32'h44db8399, 32'hc375c893, 32'h434289c3},
  {32'hc459f647, 32'hc2ce7d31, 32'hc3c37f0b},
  {32'h447fd48a, 32'hc3c4f21a, 32'h435ac8bf},
  {32'hc4dff72d, 32'h439406d2, 32'hc2e6f0d2},
  {32'h44dcd172, 32'h4244a694, 32'h42c0c538},
  {32'hc4cb3482, 32'hc3242dd4, 32'hc336514f},
  {32'h44a08bdb, 32'h429db69e, 32'h431c7f81},
  {32'hc50a1aa3, 32'hc31a2870, 32'hc357dbbd},
  {32'h44a24e87, 32'hc2da4e23, 32'hc2d0acc2},
  {32'hc4ce7c64, 32'h4386284e, 32'h42a6ee39},
  {32'h450f97d6, 32'hc3c2c1e5, 32'hc3bca621},
  {32'hc4908391, 32'hc3bd2105, 32'h42ebe648},
  {32'h450b5a22, 32'hc31fd42c, 32'h41b82449},
  {32'hc4f043ce, 32'h434f5e51, 32'hc2f6e9f6},
  {32'h449ee3d7, 32'h419afde4, 32'hc312b344},
  {32'hc477b22a, 32'h428cf0db, 32'hc3cf81a1},
  {32'h44b8a156, 32'hc2cca1fd, 32'hc2d3f12d},
  {32'hc4bf2e86, 32'h43208c4c, 32'h42ab3fa1},
  {32'h44fce8d7, 32'hc362b844, 32'hc37122fd},
  {32'hc4699ca4, 32'h4393a968, 32'hc28dcda0},
  {32'h44ece3e8, 32'hc2f13b89, 32'hc343af43},
  {32'hc3790d98, 32'h427edbf7, 32'h43508a5f},
  {32'h44d2b516, 32'h439e796d, 32'h4378bd83},
  {32'h42c9d470, 32'h431a7d94, 32'hc2d7c5f1},
  {32'h4520504f, 32'h438ef1ec, 32'hc40cbafc},
  {32'hc4e66ea5, 32'hc3403d04, 32'h41bbe9c5},
  {32'h44d5dc73, 32'h42b94199, 32'h43001d7a},
  {32'hc4d863b4, 32'hc3ad6c4a, 32'h4296c397},
  {32'h44e07133, 32'hc39db2df, 32'hc36a61d9},
  {32'hc4d3d700, 32'hc3184fd0, 32'h423a0a2a},
  {32'h4463e54c, 32'hc39cc72d, 32'h439ed58e},
  {32'hc4f89472, 32'h421cf6a2, 32'h42cfe8c4},
  {32'h44c0c316, 32'hc2fc511c, 32'hc32d53cd},
  {32'hc4eeeaca, 32'h4352a837, 32'hc31b6f04},
  {32'hc30ca9fc, 32'h433bffc9, 32'h4252b400},
  {32'hc3f18bfa, 32'h4392803d, 32'h42f9deed},
  {32'h43a60344, 32'hc0381941, 32'h43634cef},
  {32'hc42d137e, 32'hc2c9f859, 32'hc318a115},
  {32'h45098c61, 32'h438d32bb, 32'hc28eb5c1},
  {32'hc503b344, 32'hc34b451e, 32'hc31ef90a},
  {32'h449285a1, 32'hc3b04d10, 32'h42c8b350},
  {32'h42bd36a6, 32'hc2ff6aff, 32'h438d022b},
  {32'h450b54a1, 32'h402d9d8d, 32'h431f8a6b},
  {32'hc5061bee, 32'h40ffb402, 32'h41f9398d},
  {32'h44d8a9c8, 32'h438839fa, 32'hc33c0caf},
  {32'h41858a60, 32'hc2425afd, 32'h42823ea8},
  {32'h45063c44, 32'h43b7d9df, 32'hc22b3a37},
  {32'hc4ae8a88, 32'hc2d8aace, 32'hc1d54f91},
  {32'h44b5a0a0, 32'hc2badbf6, 32'h41a97c9f},
  {32'hc4b36a69, 32'h411ccfe5, 32'h41b307a2},
  {32'h44b9fb71, 32'hc30c79a4, 32'h420c03e3},
  {32'hc4df0fe3, 32'hc2c1be3f, 32'hc360e695},
  {32'h4506e079, 32'hc28a1447, 32'hc28bced8},
  {32'hc3623bc8, 32'h438eda68, 32'hc3c2059d},
  {32'h443a0248, 32'h4329ef18, 32'h43996c16},
  {32'hc4c590dd, 32'hc11c248b, 32'hc3351434},
  {32'h44c47050, 32'hc353ec4a, 32'h43196812},
  {32'hc37e2944, 32'h43850a9f, 32'hc2dee73c},
  {32'h442199fc, 32'hc370e93f, 32'h44078673},
  {32'hc407bd0c, 32'h42069e4e, 32'h40950b0c},
  {32'h44b70819, 32'h43654236, 32'h43398db0},
  {32'hc3f9aeef, 32'h4339e70b, 32'h4310da24},
  {32'h44572ec4, 32'h3f6e3250, 32'hc39d8581},
  {32'hc4847d8a, 32'hc3057db9, 32'h43044a88},
  {32'h42fd4bb4, 32'hc1feeca5, 32'h43f09aa3},
  {32'hc4ac4dc2, 32'h4306fd39, 32'h43d9d15a},
  {32'h440d0534, 32'h42deeb31, 32'hc3fcd878},
  {32'hc513e4da, 32'hc204f3a1, 32'hc2de0966},
  {32'h45051e7b, 32'h41b34c31, 32'h436c1df3},
  {32'hc4897886, 32'hc3b2ee1c, 32'h4261c0fa},
  {32'h44b9c126, 32'hc1af7074, 32'hc396e087},
  {32'hc3acfbe8, 32'hc25fc44e, 32'h4307cff4},
  {32'h439b5457, 32'hc313ae2b, 32'h430c21ad},
  {32'hc4788170, 32'hc326b72a, 32'h432f732a},
  {32'h44978678, 32'h43ff54c3, 32'hc1a6ec4e},
  {32'hc4b76be3, 32'h422c1683, 32'hc34bcf75},
  {32'h44916f6e, 32'hc391f1ea, 32'h43e18398},
  {32'hc365c860, 32'h41397474, 32'hc33d63aa},
  {32'h445b5962, 32'h43908152, 32'hc30f7474},
  {32'hc350ae86, 32'h42d3fd95, 32'hc3297570},
  {32'h440bfb87, 32'h42347404, 32'hc35d354f},
  {32'hc4d891a1, 32'h4343cfc0, 32'hc2530028},
  {32'h45184a08, 32'hc386ad41, 32'hc3737d54},
  {32'h437dad0e, 32'h4367f35c, 32'h43c72692},
  {32'h4470ef80, 32'h4294bcc1, 32'h42fb802f},
  {32'hc50f978d, 32'hc3aac1a1, 32'hc240b74b},
  {32'h45142a44, 32'hc3707b5e, 32'h430840c1},
  {32'hc4b4cbe4, 32'hc2814754, 32'h3f15d7b8},
  {32'hc28adc50, 32'hc315f4dd, 32'h439ed726},
  {32'hc4c3913a, 32'hc411a208, 32'h4391b7c0},
  {32'h450f2ee0, 32'h41f04601, 32'h42926ef8},
  {32'hc34fdbf8, 32'hc2bc8937, 32'h426b5327},
  {32'h44d7254f, 32'hc31f4152, 32'hc34655be},
  {32'hc3e58438, 32'h431eddc0, 32'h411a7c4f},
  {32'h44e54cf1, 32'hc33f173e, 32'hc3468426},
  {32'hc51188ca, 32'h410d5d1a, 32'h41e1c15b},
  {32'h44d50fd9, 32'h40c0af4b, 32'hc2214bb0},
  {32'hc38b3b40, 32'hc2cb3cdd, 32'h433161a1},
  {32'h451b0387, 32'h438441ba, 32'h42da6bb5},
  {32'hc51838fb, 32'h420cb2a2, 32'hc20c84c0},
  {32'h45164052, 32'hc3351326, 32'h43269d57},
  {32'hc33e4e30, 32'hc31d1f45, 32'h43424acc},
  {32'h44c9046e, 32'hc262f40d, 32'h43c40268},
  {32'hc3cf63f8, 32'hc33a55a0, 32'hc362360a},
  {32'h45012f30, 32'h4302a9ed, 32'hc34da213},
  {32'hc4a172b3, 32'hc353a3fa, 32'h43ce2bd1},
  {32'h4460f1c4, 32'h43b2aec2, 32'hc349acee},
  {32'hc486b463, 32'h42c0a71e, 32'h42aa72f3},
  {32'h4533a254, 32'h43894082, 32'hc3938220},
  {32'hc48f8869, 32'h43bac070, 32'h435f43be},
  {32'h447bddc8, 32'h43258bd6, 32'h428bae84},
  {32'hc4cbe162, 32'h438138e0, 32'h439b8ff2},
  {32'h449eeaa6, 32'h42c0de17, 32'h43df86b9},
  {32'hc2bed700, 32'hc3c1b423, 32'hc32534fa},
  {32'h448a9295, 32'hc281d155, 32'hc36b0f09},
  {32'hc43046f6, 32'h42e91033, 32'h42d5354a},
  {32'h438aa864, 32'hc30e7fb7, 32'h41c42ffe},
  {32'hc47912c4, 32'hc33a5624, 32'h43ea8fa2},
  {32'h442625c1, 32'h437c03fb, 32'hc3779d8a},
  {32'hc45020a0, 32'h4314f330, 32'hc34417be},
  {32'h4484b0b6, 32'h438d1f21, 32'hc2cd7425},
  {32'hc4fd8441, 32'h439a05a3, 32'h401762c4},
  {32'h42c536bc, 32'h4354244b, 32'hc348fac1},
  {32'hc3d9d1c0, 32'hc33d7b35, 32'hc34017ed},
  {32'h43c159de, 32'h3fa27f85, 32'hc32633ed},
  {32'hc513cc0e, 32'hc3968876, 32'h414e864e},
  {32'h4525ecf8, 32'h43bb416e, 32'hc2605ac1},
  {32'hc3d55258, 32'hc38846bf, 32'h42d4c372},
  {32'h44fba906, 32'h425051f9, 32'hc3b92393},
  {32'hc4d20886, 32'h41dfe057, 32'h43848b77},
  {32'h451cb8ce, 32'h43c8c09e, 32'hc33bcfc5},
  {32'h4330b090, 32'hc2b77cf2, 32'hc28a11b6},
  {32'h450737a6, 32'h4148a6f5, 32'h4129c3d6},
  {32'hc4116850, 32'hc322e6d6, 32'h4306a2c4},
  {32'h44a22914, 32'h43bbbe68, 32'hc3e06bb6},
  {32'hc4ecdd60, 32'hc29e2b46, 32'h43286b94},
  {32'h44f86c52, 32'hc281b8fc, 32'hc366f0d9},
  {32'hc44476bd, 32'hc2e35f2a, 32'h4288db7c},
  {32'h44c9387c, 32'h43214507, 32'hc40a194b},
  {32'hc4b37ae3, 32'h437307d6, 32'hc2d34452},
  {32'h44e64d2c, 32'hc0954c69, 32'hc3a1d9d9},
  {32'hc4e00a53, 32'hc2162c63, 32'hc31b2cec},
  {32'h44b937af, 32'hc2e605fe, 32'h424be4ce},
  {32'hc3dce5c8, 32'h435f08c3, 32'h432d5a4c},
  {32'h44f6e986, 32'h43d3e79f, 32'hc37b63cd},
  {32'hc4945e0e, 32'hc0a5745b, 32'hc295e338},
  {32'h44dca55a, 32'hc396b8f5, 32'hc3c3a369},
  {32'hc4d27504, 32'hc38d84d1, 32'h4377b7a5},
  {32'h4491f37f, 32'hc27d3d1c, 32'h429c6824},
  {32'hc4f1d267, 32'hc3898ab7, 32'hc3e37e33},
  {32'h438bae90, 32'h42bb91fd, 32'hc2a8a93c},
  {32'hc4b8f274, 32'h409a580e, 32'h4351d553},
  {32'h43a16120, 32'hc2ae677e, 32'h40a9b038},
  {32'hc4f5c29d, 32'hc3decd1e, 32'h43003c83},
  {32'h43be9d88, 32'h43832e34, 32'h4314c871},
  {32'hc481251c, 32'h4335200a, 32'h4369524a},
  {32'h4426bc72, 32'h41f91d3c, 32'hc3bbc027},
  {32'hc49669ea, 32'hc38a4f3a, 32'hc2047608},
  {32'h4472f05b, 32'h435a623c, 32'h429e86fc},
  {32'hc50f3066, 32'h427b628e, 32'h4387412d},
  {32'h448a833c, 32'hc3abf548, 32'hc327df1d},
  {32'hc515873e, 32'h43331bba, 32'hc001c15a},
  {32'h44be289d, 32'h43826fdb, 32'h42ad7c53},
  {32'hc431d193, 32'h41331d4a, 32'hc349fa72},
  {32'h44128d43, 32'h4354d5a0, 32'hc32873eb},
  {32'hc356dc00, 32'hc309e10c, 32'hc216251a},
  {32'h448b3c22, 32'hc40c77ef, 32'hc3da3694},
  {32'hc429aef2, 32'h424eb6da, 32'h40d2b85b},
  {32'h4420bc60, 32'hc281aaa2, 32'hc3abec34},
  {32'h44773bc1, 32'h439747fe, 32'hc3860d33},
  {32'hc4406052, 32'h424005af, 32'hc2a926dc},
  {32'h44d5f00a, 32'hc3e0bfed, 32'h43be9a7d},
  {32'hc41ee1c4, 32'h42dd8938, 32'hc1b04b88},
  {32'h44f01ce2, 32'hc33e819b, 32'hc3b937c8},
  {32'hc48e7c4f, 32'h438d2300, 32'hc3d950c4},
  {32'h4493491a, 32'hc392d00f, 32'hc3bcd6d2},
  {32'hc412ce7e, 32'h43095bc3, 32'hc2a8153b},
  {32'h44f2005c, 32'hc313e334, 32'hc35fe6b8},
  {32'hc3d316b4, 32'h43ba6020, 32'h42d6e1b0},
  {32'h44da2472, 32'h42c378ea, 32'hc3086b47},
  {32'hc4bb2a21, 32'h426d89ac, 32'h4242da6e},
  {32'h4499e15b, 32'h4397fe51, 32'h42afb458},
  {32'hc422b0b9, 32'h41a9a6f4, 32'hc35ed4f7},
  {32'h44e573fc, 32'hc3845405, 32'h4303227b},
  {32'hc4d29c0c, 32'h42a3af7a, 32'h426df13a},
  {32'h449b7ae6, 32'h433b72b4, 32'h4236b842},
  {32'hc4ed7b35, 32'h4285cf84, 32'hc226f6bc},
  {32'h4445ce9f, 32'h42d8c91a, 32'hc334d448},
  {32'hc4d8ad9f, 32'h42a8cc31, 32'hc39ba890},
  {32'h44b94be1, 32'h40b8e7da, 32'h4309b616},
  {32'hc320603e, 32'hc3b8521d, 32'h42132109},
  {32'h44684d40, 32'h437616c9, 32'h438dc126},
  {32'hc41ffb9e, 32'h432f6155, 32'hc238a99f},
  {32'hc3c6df49, 32'hc2f501ec, 32'hc206754d},
  {32'hc441cf99, 32'h4309d815, 32'h43f1c32e},
  {32'h448e74bb, 32'h43a811bc, 32'hc21dc75e},
  {32'hc4dd5c6e, 32'h430247b6, 32'h437977ad},
  {32'h4469151c, 32'hc10b4125, 32'hc287eca1},
  {32'hc4ef1420, 32'h43a482a9, 32'hc35965ba},
  {32'h4504b425, 32'hc3c1b4a5, 32'h431daa27},
  {32'hc43d3769, 32'hc3a63feb, 32'h4396f48d},
  {32'h444e23db, 32'hc2f98518, 32'h41b1525f},
  {32'hc465c78d, 32'hc3b14e45, 32'h431e5c3a},
  {32'h44f84faa, 32'hc2640e7c, 32'hc3655cf3},
  {32'hc4fd6baa, 32'hc38db830, 32'h43adfc6f},
  {32'h44c26918, 32'hc314ad73, 32'hc41ca694},
  {32'hc3d7831f, 32'hc3489a06, 32'h42dc3eec},
  {32'h44af461c, 32'h4259dccf, 32'h431fadb2},
  {32'hc449240b, 32'hc22315bb, 32'hc3f9434c},
  {32'h44cc385e, 32'hc32eacdc, 32'h4372580f},
  {32'hc4fb936d, 32'h41e4c7de, 32'hc2ad13d2},
  {32'h442973be, 32'h436ce51f, 32'h4089afa9},
  {32'hc445a79d, 32'hc280e8eb, 32'h428d41f0},
  {32'h43d11cdc, 32'hc29c45fb, 32'hc1865a9c},
  {32'hc41aa994, 32'h4349fd5b, 32'hc38c66c8},
  {32'h450a54f9, 32'hc25f40c6, 32'hc28e583a},
  {32'hc50d9ea4, 32'h437fa23e, 32'hc368fc0a},
  {32'h44461204, 32'h446699a2, 32'hc3956177},
  {32'hc3ae7cbc, 32'hc24ae847, 32'h43d61a57},
  {32'h452e93f5, 32'h43255d1d, 32'h4304f9ae},
  {32'hc4bf5851, 32'hc3b2b1dc, 32'hc30af25c},
  {32'h43c8b348, 32'h439a3c91, 32'hc2a00082},
  {32'hc4bd9660, 32'h3febfc20, 32'hc266b267},
  {32'h451b2610, 32'hc2a37393, 32'hc2d33887},
  {32'hc4e58f21, 32'h429af24b, 32'h41aab3e3},
  {32'h441e22cb, 32'h43edff3d, 32'hc0edabee},
  {32'hc50eaac1, 32'h41f0d62d, 32'hc3b2741f},
  {32'h440307ba, 32'h42b60ee6, 32'h417f274d},
  {32'hc46f9e76, 32'h416a5bae, 32'hc34d20cc},
  {32'h450f7cca, 32'hc35c9405, 32'h43d785e4},
  {32'hc38e5631, 32'h41fbbb04, 32'hc2d6da0a},
  {32'h44cd25ed, 32'h44044fde, 32'hc393123c},
  {32'hc4da651d, 32'h437de49c, 32'hc2f29a55},
  {32'h44c2b354, 32'h43140b95, 32'h43c8e0dc},
  {32'hc370ad6c, 32'hc4245a65, 32'h43e560d7},
  {32'h44cd0152, 32'hc31c981d, 32'h42969383},
  {32'hc4f9c189, 32'hc3cc5828, 32'hc1da5e6c},
  {32'h44d852fe, 32'h430dc947, 32'h429de1ce},
  {32'hc49f1d00, 32'h42ebfa5e, 32'h4336b505},
  {32'h4300226a, 32'hc2bddc87, 32'hc2ab1232},
  {32'hc4ca6c5a, 32'h43293b5c, 32'h43454f21},
  {32'h440697d1, 32'h43720450, 32'h439f4956},
  {32'hc3f58fae, 32'h438570f5, 32'h438216b6},
  {32'h44b6e9fc, 32'hc3955f66, 32'hc2637929},
  {32'hc4376bb4, 32'hc23e3880, 32'h431e935e},
  {32'h44b66158, 32'h42ad8ef4, 32'hc391fd91},
  {32'hc4fe9e1c, 32'hc333de16, 32'h43159d10},
  {32'h449a8355, 32'h43a35396, 32'hc335cb64},
  {32'hc3bd1f3c, 32'h42493488, 32'h42833c21},
  {32'h4506c43a, 32'hc3be8ec2, 32'h430ccf06},
  {32'hc4e337f7, 32'h43376634, 32'h41d3dd36},
  {32'h44ebd1fc, 32'hc316c877, 32'hc2c6f7aa},
  {32'hc3e4e7f0, 32'hc1653e8f, 32'h43405339},
  {32'h44f419e7, 32'h430e040e, 32'h43295083},
  {32'hc4d2978c, 32'h43a05129, 32'h43814536},
  {32'h4488d71e, 32'hc3524600, 32'hc2832d46},
  {32'hc49365a5, 32'hc2f03012, 32'h41c67918},
  {32'h44c856cf, 32'hc3d52b7d, 32'h437e0167},
  {32'hc38edc0c, 32'hc222f79a, 32'h425a7dd3},
  {32'h44a3b77d, 32'h43b7164d, 32'h43012f20},
  {32'hc3c0598c, 32'hc29b92ee, 32'h437d1474},
  {32'h450e7e1f, 32'h43336d30, 32'hc33c5200},
  {32'hc45b0a43, 32'h42a7177c, 32'hc38ef300},
  {32'h4504a83c, 32'h4420c862, 32'hc2c29462},
  {32'hc317dbf0, 32'hc39082b4, 32'hc326261a},
  {32'h435a9320, 32'h4385efd4, 32'h4307a642},
  {32'hc3ae7a50, 32'hc1d55efa, 32'h430336d4},
  {32'h4458f100, 32'hc35cf619, 32'hc208499e},
  {32'hc50109c6, 32'h422345d9, 32'h42c02422},
  {32'h450d1b34, 32'h4359ebcf, 32'hc28113a8},
  {32'hc4224e9d, 32'hc307e98b, 32'h42461619},
  {32'h44bd8604, 32'hc341b23d, 32'hc117caab},
  {32'hc495c850, 32'hc28293e9, 32'h43622014},
  {32'h4486a940, 32'h409ab732, 32'h42e85a29},
  {32'hc3b52416, 32'hc3e2b5c9, 32'hc2aacbd8},
  {32'h4526459e, 32'hc3a9731b, 32'hc2b9cbc8},
  {32'hc43a4157, 32'hc103b774, 32'h42bf7b38},
  {32'h44a1bc34, 32'hc26dd6c6, 32'hc2fdd6be},
  {32'hc420a22c, 32'hc2620744, 32'hc3908485},
  {32'h448d04aa, 32'hc3513e64, 32'h429c47e8},
  {32'hc49f21ac, 32'hc310ea9a, 32'hc1cd71cb},
  {32'h44f6a6ad, 32'h429d7364, 32'h429aa2ef},
  {32'hc4b14edf, 32'hc2e5be40, 32'h4372a9d0},
  {32'h451d7a81, 32'h43d0a99c, 32'hc2deb89e},
  {32'hc4cbf25f, 32'hc1f35384, 32'h429e41f8},
  {32'h4460a1ba, 32'hc32f3100, 32'hc35d32af},
  {32'hc4bf72de, 32'hc40c495f, 32'hc2337458},
  {32'h450e5b18, 32'hc2ec6331, 32'hc24ef0a5},
  {32'hc417a213, 32'h438ca417, 32'h43b42eeb},
  {32'h4436b242, 32'h4364ae4c, 32'hc3239711},
  {32'hc3da57d8, 32'hc34daee5, 32'hc29c45e0},
  {32'h45114aec, 32'h43ad89c4, 32'h43490771},
  {32'hc207a740, 32'h423b0a6b, 32'h434fba71},
  {32'h44baf46f, 32'hc260005d, 32'hc03b26e0},
  {32'hc4a46bcd, 32'h43e8f36b, 32'hc309066f},
  {32'h44fce493, 32'h42ec9f34, 32'hc34b5510},
  {32'hc4468865, 32'h437f8eae, 32'hc30a7f33},
  {32'h4341ee58, 32'h4368c330, 32'h42f92f83},
  {32'hc5101216, 32'hc33ac160, 32'h440ec632},
  {32'h44a7dda4, 32'hc340065b, 32'h42fed563},
  {32'hc4fa64f2, 32'hc3efd4c3, 32'hc3391852},
  {32'h44e67d47, 32'h431d50ed, 32'hc32dcc9b},
  {32'hc4c1fb52, 32'h42b20d1d, 32'hc209d86e},
  {32'h441d476a, 32'hc28b773e, 32'h4005acd6},
  {32'hc3e7ff64, 32'h4361fd88, 32'hc0c2928d},
  {32'h450c8b7f, 32'h41d89697, 32'h4311211e},
  {32'h40cd2c20, 32'h428adc59, 32'hc30d2f35},
  {32'h43267cc9, 32'hc32de9af, 32'hc3057cb8},
  {32'hc27ef8c0, 32'h4308b323, 32'hc396889a},
  {32'h44a1b22f, 32'hc2279a19, 32'hc31715de},
  {32'hc1d32f70, 32'hc2e70039, 32'hc27f0c6f},
  {32'h44030c33, 32'h42f1e227, 32'hc31f62bc},
  {32'hc43c140e, 32'hc1f2a9b6, 32'h441d7975},
  {32'h43a1cde9, 32'h41a72b7f, 32'h43ab61eb},
  {32'hc494a86c, 32'h42c0c3bc, 32'h42a01f71},
  {32'h421b4eb6, 32'h41a3fc0b, 32'h438af22f},
  {32'hc4c9c2f1, 32'hc3213aa0, 32'hc3405792},
  {32'h44c13d5a, 32'hc3e78cda, 32'hc2bb17e3},
  {32'hc4c7be29, 32'h43f7a083, 32'hc35dd41b},
  {32'h45017bec, 32'h43826fa2, 32'hc3bcf746},
  {32'hc4d0e3f8, 32'h435e275d, 32'h42e9b580},
  {32'h44f374f7, 32'hc201a6d9, 32'hc33a650d},
  {32'hc497ecbc, 32'hc3e64aba, 32'h421c5e00},
  {32'h44ed9fd2, 32'h433de7cc, 32'h410a2c86},
  {32'hc509fbf6, 32'h432966ec, 32'hc2739215},
  {32'h44da5eea, 32'h42fa6b65, 32'h43903cc1},
  {32'hc1683280, 32'h432c35b8, 32'hc3004037},
  {32'h44de7977, 32'h43d2318c, 32'hc23cd4fd},
  {32'hc4d4de00, 32'h43945ae5, 32'hc2d3f685},
  {32'h4413f471, 32'hc1d06257, 32'h436cdf6a},
  {32'hc4e5b638, 32'hc3076ad5, 32'hc298caeb},
  {32'h4401fe02, 32'h43cc8442, 32'hc2af6fe8},
  {32'hc4a77c6f, 32'hc18a006a, 32'h430930f5},
  {32'h44932ab6, 32'hc321c01a, 32'h42592922},
  {32'hc4440740, 32'hc29af087, 32'h43640537},
  {32'h450a90bb, 32'h41a27e68, 32'hc39cd50a},
  {32'hc50a47a9, 32'hc34a200d, 32'h43519a84},
  {32'h44f6f70c, 32'h43747ee8, 32'h42770678},
  {32'hc49ef6d0, 32'h434ca5f0, 32'h42f1568f},
  {32'h4420cebb, 32'hc10100ed, 32'h4247cbae},
  {32'h43a4e290, 32'h434651a5, 32'hc3409758},
  {32'h4481297a, 32'h4355994b, 32'h43c5cd84},
  {32'hc4e95986, 32'hc3815d7a, 32'hc318dff4},
  {32'h44b337f3, 32'h4301d876, 32'h4344dfea},
  {32'hc365c4bd, 32'h43baef45, 32'h42927655},
  {32'h443b133e, 32'h43ec2a9a, 32'h4357b821},
  {32'hc4f7736c, 32'hc295f0ac, 32'h41141400},
  {32'h4506e3fc, 32'hc3548c76, 32'hc29bb860},
  {32'hc4f025e6, 32'hc2b5a369, 32'hc2612111},
  {32'h444d8d93, 32'hc376302d, 32'h434fe25c},
  {32'h3f0cf400, 32'h42d629e4, 32'hc3a20f7b},
  {32'h44864143, 32'hc3c765da, 32'hc290a9af},
  {32'hc30372a7, 32'h4219b418, 32'hc3b9229b},
  {32'h44b4d2de, 32'hc3a7d359, 32'h41917110},
  {32'hc3de9310, 32'h439f2f74, 32'hc3049038},
  {32'h44652636, 32'hc26bb9d4, 32'hc30aee1c},
  {32'hc4ad1d64, 32'h4347b4cd, 32'hc2d4210d},
  {32'h447f5180, 32'h436e8224, 32'hc32e095f},
  {32'hc487882a, 32'h432bc4e9, 32'hc35896b7},
  {32'hc341cfa3, 32'hc354d7b5, 32'h438528e1},
  {32'hc4ce2d5c, 32'h43877e4b, 32'h42ca6264},
  {32'h43be2ca0, 32'hc4072a4d, 32'hc3f8ccbe},
  {32'hc46b6d41, 32'hc306ae77, 32'h42f00af6},
  {32'h43b3e3f0, 32'hc37973b5, 32'h42b62999},
  {32'hc4301ac2, 32'hc30254ed, 32'h43a14444},
  {32'h44d4025d, 32'h430cbf37, 32'h4394db64},
  {32'hc48b4cd8, 32'hc3a7bae6, 32'h42eb3863},
  {32'h44a06eb2, 32'hc2e9ad06, 32'h43923348},
  {32'hc407f5ee, 32'hc37c8956, 32'hc1915010},
  {32'h449f4790, 32'h438e5705, 32'hc1e76e3f},
  {32'hc4b7c7be, 32'hc1c13e4e, 32'hc36f3f24},
  {32'h44f06d70, 32'hc1b211de, 32'h42a9236d},
  {32'hc4cbbc92, 32'hc1ae34be, 32'h41d57f70},
  {32'h4426acd8, 32'h42df08f1, 32'h429bf680},
  {32'hc4bc7a28, 32'hc147c110, 32'hc3a48c42},
  {32'h44ca125f, 32'hc32c4e70, 32'hc35e5cd2},
  {32'hc4f336f3, 32'hc2480b2d, 32'hc3aedef5},
  {32'h44149e0a, 32'h4298d757, 32'hc30b0fbd},
  {32'hc4e2f0bf, 32'h41fda71d, 32'h41bac0b0},
  {32'h4523b1d7, 32'h43581783, 32'hc366fd03},
  {32'hc4db86a5, 32'hc2d961ec, 32'h4338dd08},
  {32'h44898a8b, 32'h421841b6, 32'hc2885b03},
  {32'hc523f7a5, 32'h4309a6b9, 32'hc3656298},
  {32'h44b20b5b, 32'h42f73867, 32'h416c67a4},
  {32'hc4acecab, 32'hc0e5fc22, 32'hc2996ce5},
  {32'h43c0207c, 32'hc3a050c4, 32'hc31f1ad5},
  {32'hc4c6a471, 32'h4227e844, 32'h43eb23c2},
  {32'h430e7308, 32'hc2931f98, 32'hc2e912be},
  {32'hc4aa9c2a, 32'hc3898c34, 32'h43441204},
  {32'h44efb526, 32'hc3cb7164, 32'hc3cb1a37},
  {32'hc4d388fc, 32'h42839e9a, 32'hc3238591},
  {32'h443b4ab9, 32'hc2978f5d, 32'h438782e8},
  {32'hc4fc3eaf, 32'hc2ad9587, 32'h432705d9},
  {32'h44b11afe, 32'hc279748a, 32'hc3fed432},
  {32'hc4e9784c, 32'h42c218aa, 32'hc3834c4c},
  {32'h4238c7e0, 32'h443c99bc, 32'h43bb6f7b},
  {32'hc4dd76a8, 32'hc2fc2f09, 32'hc3a49b75},
  {32'h43aa8cc9, 32'hc40187ec, 32'h433321ae},
  {32'hc4a2c9ce, 32'h432736a3, 32'hc3075978},
  {32'h44ffee21, 32'h43b728f2, 32'hc179cc2b},
  {32'hc4d4d6ce, 32'h43703e0b, 32'h42a91893},
  {32'h44e3e552, 32'h43ca7592, 32'hc1fa0be8},
  {32'hc4938184, 32'hc35b5d02, 32'hc388df29},
  {32'h4512673e, 32'hc31acc55, 32'h4349cc2f},
  {32'hc439ce27, 32'hc083a63a, 32'hc37480e6},
  {32'hc321f3c8, 32'h43640e8c, 32'h4129b482},
  {32'hc42ebc20, 32'hc27e9c8c, 32'hc3723018},
  {32'h44ebc2d2, 32'hc309cd4b, 32'h430a0016},
  {32'hc301c3b4, 32'hc3443394, 32'h438f1816},
  {32'h4497b2b8, 32'h43388e87, 32'hc40d89df},
  {32'hc4a71401, 32'hc309bb56, 32'h422e4afc},
  {32'h4383e550, 32'h43037bcd, 32'hc38e9382},
  {32'hc451f7c7, 32'h434d8b87, 32'hc2b0373b},
  {32'h43fb81fc, 32'hc11d5c7a, 32'hc3816043},
  {32'hc49a1263, 32'hc1a8ba4d, 32'h42e19951},
  {32'h450cdab9, 32'hc3a36c55, 32'hc3c68f80},
  {32'hc4aa1fd9, 32'h43ba93b5, 32'h4380e252},
  {32'h441da38b, 32'hc3bf8ce8, 32'hc3751074},
  {32'h430d5370, 32'hc2c7eeb9, 32'h42cdbf53},
  {32'h45093978, 32'h4390a5dc, 32'h43a450ad},
  {32'hc3ebf738, 32'hc2c3825d, 32'hc282b223},
  {32'h44819aa7, 32'hc1e060a6, 32'h4346f680},
  {32'hc3e7000c, 32'h42f71d3f, 32'h42958803},
  {32'h44942b71, 32'h439d5447, 32'h42865fb5},
  {32'hc38c6900, 32'hc3c6b059, 32'h439ef7f2},
  {32'h44bf76b0, 32'hc2d14f66, 32'h43315ddc},
  {32'hc4be0743, 32'h43966e4d, 32'hc27841c0},
  {32'h4502dcf3, 32'h429d2d96, 32'h43e14c79},
  {32'hc3a3ca0c, 32'h434d5c0d, 32'hc3612ce8},
  {32'h44ecc55a, 32'h439a7869, 32'h435f7213},
  {32'hc50a538b, 32'h42656a2a, 32'h43922c86},
  {32'h451b0c26, 32'h430cfe2e, 32'h41562e8e},
  {32'hc4e20917, 32'hc2da0b82, 32'h4369ed05},
  {32'h44d37aab, 32'h4223f1de, 32'h430ac936},
  {32'hc39c4c68, 32'hc22fbd74, 32'h42e3e4c3},
  {32'h451d8987, 32'h440b7c07, 32'h41d0446c},
  {32'hc43c22b3, 32'hc2f8a9b0, 32'hc3528eea},
  {32'h44a72c16, 32'h43dbc382, 32'hc39dcc5b},
  {32'hc4cdc47c, 32'hc3b1f266, 32'hc2ba0aaf},
  {32'h44b0f09d, 32'h43b6afbc, 32'h4297fa73},
  {32'hc433b88e, 32'hc285c3b6, 32'h43417612},
  {32'h4455026c, 32'hc30bcbd1, 32'h423191c0},
  {32'hc4cafd46, 32'h42a0d48b, 32'hc3803a36},
  {32'h42b61940, 32'hc3b4625c, 32'h4300eb78},
  {32'hc4313754, 32'h430f7a8b, 32'h43f7e666},
  {32'h44225e7f, 32'hc19f14f3, 32'hc2c8bb46},
  {32'hc4b14891, 32'h425635aa, 32'hc3bf26cc},
  {32'h439f1998, 32'h43839bd3, 32'h43474c7c},
  {32'hc4a0487c, 32'h431d8063, 32'hc294b708},
  {32'h44cf39fe, 32'h430aa2e4, 32'hc3f1b626},
  {32'hc462e76e, 32'h42c9201c, 32'hc394b955},
  {32'h43735268, 32'hc1d821c6, 32'hc1c74290},
  {32'hc48a60af, 32'h430bff0d, 32'h42d1f085},
  {32'h44bbc4c2, 32'h42f3ff08, 32'h42a074af},
  {32'hc49389c6, 32'h43dcba48, 32'hc35022dc},
  {32'h44534b73, 32'h41e7ff20, 32'hc30e2276},
  {32'hc49bb116, 32'h439739c6, 32'hc270688e},
  {32'h43d27b5f, 32'hc3a708b4, 32'h432b06a1},
  {32'hc3a87a56, 32'h4294e7b1, 32'hc33ad9db},
  {32'h451d5a53, 32'h422b405a, 32'h42eb6aec},
  {32'hc406d078, 32'h4157b32a, 32'h420cab22},
  {32'h44827a27, 32'hc3193c1a, 32'hc2619e04},
  {32'hc4649880, 32'h4381e833, 32'hc219e5dc},
  {32'h440680f2, 32'hc2ab10ab, 32'h41e9d0b0},
  {32'hc4a29ecd, 32'hc0f4d688, 32'hc2ba5f40},
  {32'h44afccbd, 32'h42f2ed4b, 32'h4345d0b7},
  {32'hc4955f2d, 32'h41e2bad9, 32'h421b4cb4},
  {32'h448c4ba2, 32'hc23eb503, 32'hc2ef1cf7},
  {32'hc4ff70a3, 32'h431e128b, 32'hc2af29be},
  {32'h43cc453b, 32'h4294f894, 32'h409218a5},
  {32'hc41ff4ec, 32'h431904ce, 32'h420485f2},
  {32'h44eb799c, 32'h42bb417d, 32'hc28fd072},
  {32'hc4ffc230, 32'h42ed489d, 32'hc30b5f4e},
  {32'h43e70808, 32'h43939568, 32'h428f5519},
  {32'hc434ae71, 32'h432cf8da, 32'h43896233},
  {32'h44ee6790, 32'h43d4f359, 32'hc319fd8b},
  {32'hc3e99518, 32'hc3436ada, 32'h43812aec},
  {32'h44cba2c6, 32'h435a1b42, 32'h43b59c14},
  {32'hc4c418ba, 32'h4309d99a, 32'hc245d8f8},
  {32'h43b579d0, 32'h432ee09e, 32'h43cea5ac},
  {32'hc5091760, 32'hc26157da, 32'h429f39eb},
  {32'h44e68837, 32'h43dc74a8, 32'h438ac27a},
  {32'hc4403ace, 32'h43139efe, 32'h43240fac},
  {32'h44ed6cbc, 32'hc3571e81, 32'h420946fe},
  {32'hc50cf4b2, 32'hc3b3eac5, 32'h422d3340},
  {32'h43a9233c, 32'hc2e32e39, 32'h41408bf5},
  {32'hc5038245, 32'hc35640c8, 32'hc2be6896},
  {32'h44ecfcb8, 32'h430a0aaa, 32'hc3193f7c},
  {32'hc4238fa3, 32'hc39b80bb, 32'h42f254ad},
  {32'h45008d11, 32'h42ae7c67, 32'h434615c1},
  {32'hc46416a8, 32'hc02c4190, 32'hc262f6e6},
  {32'h44f37989, 32'h430a510f, 32'h40fb7da5},
  {32'hc508f34d, 32'h42d2bb36, 32'hc36175ab},
  {32'h44a9689e, 32'h4215b9de, 32'h41eb4d0f},
  {32'hc44f5bd2, 32'hc255a830, 32'hc336b623},
  {32'h44e7b96c, 32'hc361acd3, 32'h415ce883},
  {32'h42945c58, 32'h434ce676, 32'h43511492},
  {32'h441a1bea, 32'h4306f19a, 32'hc38f6ae4},
  {32'hc4fd9246, 32'h42ab3668, 32'hc2925b03},
  {32'h44c31658, 32'h42540f93, 32'h4324fbc1},
  {32'hc4d21bdf, 32'h4319564c, 32'h42af581d},
  {32'hc2efe44c, 32'hc33d65ef, 32'hc373259a},
  {32'hc4b8d604, 32'hc23b8ec6, 32'h42a2c7ef},
  {32'hc3040f84, 32'h431c83a6, 32'h42e93a5c},
  {32'hc4dfa3cb, 32'h42858ace, 32'hc2d8e31f},
  {32'h44d852b0, 32'h42004454, 32'hc2a1dcdc},
  {32'hc41ef045, 32'hc3786234, 32'h437689f0},
  {32'h43fd4748, 32'h431ab23b, 32'h42db0c8a},
  {32'hc50fc62c, 32'h43b7edb8, 32'hc3f65545},
  {32'h42972038, 32'h43cbf8cd, 32'hc30b7f9f},
  {32'hc3b135f2, 32'h4235f4e6, 32'hc30ee6e2},
  {32'h44dbb3ee, 32'hc04b0fc1, 32'hc34f9105},
  {32'hc4edb975, 32'h4334204c, 32'hc330ef21},
  {32'h451da90d, 32'h42e62a5e, 32'hc3f014d5},
  {32'hc49e16b7, 32'h4342b4d5, 32'h434ca86e},
  {32'h42d2a108, 32'hc350aadd, 32'h437e73b2},
  {32'hc401e6c1, 32'hc0f6f735, 32'hc3846ee7},
  {32'h446387b2, 32'h43889ab6, 32'hc3cb211a},
  {32'hc4c78a38, 32'hc3ee46bb, 32'hc316dfe0},
  {32'h4408ce24, 32'hc230e518, 32'hc2f96060},
  {32'hc4fc2ff7, 32'hc283a1bc, 32'h434641cb},
  {32'h44695ff2, 32'h42142088, 32'h4245cd3b},
  {32'hc435cdff, 32'hc2acb7be, 32'hc30386eb},
  {32'h44841413, 32'h428783cb, 32'hc33c6061},
  {32'hc4bc30c1, 32'h432964db, 32'hc23844b0},
  {32'h4516d91e, 32'h422ca6bc, 32'hc391735b},
  {32'hc3ec6231, 32'h43ad2181, 32'h43800a0d},
  {32'h44647a37, 32'h4235d09f, 32'hc317a4f1},
  {32'hc405a92c, 32'h424d0eb2, 32'h4405fd51},
  {32'h44dd4c37, 32'hc394d14e, 32'hc292f63f},
  {32'hc4d8cecc, 32'hc20a5184, 32'h437ca58f},
  {32'h441004f8, 32'hc3fd492c, 32'hc0db7baa},
  {32'h405cf600, 32'h431b70dc, 32'h4274eff4},
  {32'h44d29573, 32'hc2fc51f8, 32'hc354c544},
  {32'hc40066e0, 32'h436c32b5, 32'h431593d5},
  {32'h44fc8dbe, 32'hc2369d21, 32'hc2fa189c},
  {32'hc505c2e3, 32'h42bfc18c, 32'h437d97ac},
  {32'h4501f00e, 32'h420e1bf9, 32'h43055aaf},
  {32'hc5051fb3, 32'h4299ef90, 32'h4211c82f},
  {32'h44be5867, 32'h435e70c9, 32'h42ae0e31},
  {32'hc45f8ecc, 32'hc2e4215c, 32'hc2a48f0d},
  {32'h43c16606, 32'h42dd96b5, 32'hc2d8f297},
  {32'hc5008d03, 32'hc337af95, 32'h4398b929},
  {32'h44a35f28, 32'h4306f807, 32'hc0f6b6d4},
  {32'hc3f2e494, 32'h430d47a4, 32'h43a0a22d},
  {32'h4408876e, 32'hc2a063c4, 32'h4391d60e},
  {32'hc4fe8cf8, 32'h433b7838, 32'h43a27f22},
  {32'h44f08986, 32'h42cd3914, 32'h43a2a62f},
  {32'hc46a7b78, 32'hc3788050, 32'hc288c7a2},
  {32'h44b310ff, 32'h43429953, 32'h4148aef2},
  {32'hc50a85dd, 32'hc1fb18a9, 32'hc37f83e6},
  {32'h444bb835, 32'hc327b343, 32'hc2fb8b65},
  {32'hc45027e8, 32'hc199689c, 32'hc30053bd},
  {32'h43051198, 32'hc319a8a0, 32'h430642b2},
  {32'hc4c0d819, 32'h42a5dea0, 32'hc2cedf58},
  {32'h44123116, 32'h42fa87ba, 32'h42f1976d},
  {32'hc5017ed5, 32'hc2db1a22, 32'h42548f93},
  {32'h44ce25c8, 32'h42acd957, 32'h43184790},
  {32'hc42c08d4, 32'h43091d55, 32'hc2b42434},
  {32'h4456d8ca, 32'h43f6b4e2, 32'hc354ebbd},
  {32'hc504533e, 32'hc224872f, 32'h436e37b9},
  {32'h449bde91, 32'h43b050ef, 32'hc3621a49},
  {32'hc4c40bf0, 32'hc31b9b79, 32'h42bf2435},
  {32'h4442745b, 32'h434127d6, 32'h432b1865},
  {32'hc40fe3d6, 32'h414f1651, 32'hc34d66e6},
  {32'h4451b4d2, 32'hc2f83e89, 32'h421ab63b},
  {32'hc36e23a8, 32'hc1f96f57, 32'h43228509},
  {32'hc1026680, 32'h410ba9e3, 32'h430c4c53},
  {32'hc49ff09e, 32'h4253b8a1, 32'hc32c4659},
  {32'h4511809b, 32'hc2aa7bf8, 32'hc1c770f5},
  {32'h42ebefa0, 32'h424ce352, 32'hc3bb1fcb},
  {32'h44f6d03f, 32'hc22799cc, 32'hc2bf6f73},
  {32'hc509f70b, 32'hc2168491, 32'hc4151361},
  {32'h42df6560, 32'hc39d22d1, 32'hc2df572b},
  {32'hc506be5a, 32'hc24817ce, 32'hc32d04c0},
  {32'hc33845c8, 32'h430e4e0e, 32'h436b1eb0},
  {32'hc2adb92e, 32'h431c8460, 32'hc3429da4},
  {32'h44fae328, 32'h4240f2d7, 32'h4390da33},
  {32'hc4035099, 32'h43349e07, 32'hc33edfe0},
  {32'h440496e8, 32'hc27e8490, 32'h4301c001},
  {32'hc4eb73b6, 32'h431745cd, 32'h438602aa},
  {32'h44c4606f, 32'h42037e98, 32'h43b4ae59},
  {32'hc4b7e590, 32'h436025aa, 32'h4332735f},
  {32'h44ef96a5, 32'hc22c86ad, 32'h4349060a},
  {32'h42b5d6c4, 32'hc2c5a0fa, 32'h43d13e00},
  {32'h4518c60b, 32'hc37cab00, 32'h43009b75},
  {32'hc506ac95, 32'h43360f13, 32'h41d17d53},
  {32'h4436860e, 32'h430f5864, 32'h428caeaa},
  {32'hc4af0f6c, 32'h441a207b, 32'h4292efc1},
  {32'h44bb2aea, 32'hc29df7ac, 32'h439c0bd3},
  {32'hc48d9dc5, 32'h4415158e, 32'hc4002aac},
  {32'h44e64c2b, 32'hc2e7c676, 32'hc234a760},
  {32'hc4c64dd8, 32'h432e6c85, 32'hc2d120b6},
  {32'h44c81739, 32'h42e8b1f6, 32'h43cad7f8},
  {32'hc4dcddf2, 32'h42f94069, 32'hc2be6a19},
  {32'h440cd290, 32'h4374bd08, 32'hc26c15f5},
  {32'hc47386c0, 32'h4298abc9, 32'h435e2d18},
  {32'h43fbfe29, 32'h43ad377f, 32'h43542112},
  {32'hc4497307, 32'hc3b0408d, 32'h438ac6ef},
  {32'h4470d714, 32'hc4149393, 32'hc3653902},
  {32'hc4a2d712, 32'hc3bc1ed5, 32'h431a6d7e},
  {32'hc41b7342, 32'hc3922f05, 32'hc217416d},
  {32'h43f62330, 32'h439f186b, 32'h4382bb24},
  {32'hc4c27f02, 32'h42859c17, 32'h42ac88f2},
  {32'h445fa5c8, 32'hc39ddf18, 32'h42c74ea8},
  {32'hc4f5d9d4, 32'h42200844, 32'hc25a825a},
  {32'h44aa99ba, 32'hc1c0882c, 32'hc39ce387},
  {32'hc51a8472, 32'h435219b8, 32'hc36e6131},
  {32'h44be5fd1, 32'hc319ad6f, 32'h4321e2b6},
  {32'hc4b4f102, 32'h43fd3a39, 32'hc29f3ffc},
  {32'h45034280, 32'hc2630e3c, 32'hc38c2ce9},
  {32'hc42067f6, 32'hc20e3253, 32'hc2da8bce},
  {32'h4501a7d4, 32'hc34949e9, 32'h43b0014b},
  {32'hc24e67a0, 32'hc3288dea, 32'hc2ba1afa},
  {32'h45138bae, 32'h40344248, 32'hc38c275e},
  {32'hc4f86be4, 32'h42c624e7, 32'hc36b87be},
  {32'h43684adf, 32'h42c88bc3, 32'h422d8ddf},
  {32'hc4c39ae2, 32'hc31dc6ba, 32'h423a56f4},
  {32'h44b15535, 32'h43252f1e, 32'hc3206181},
  {32'hc48b708c, 32'hc355c1c7, 32'hc1159f08},
  {32'h445eb089, 32'h41883a7b, 32'hc3dd6a2a},
  {32'hc45103f8, 32'h4352fe12, 32'hc2ded003},
  {32'h45173b54, 32'hc3aadd9d, 32'hc29fd559},
  {32'hc4bc13cd, 32'hc329b031, 32'h42c63d0d},
  {32'h45138f04, 32'hc1e4fc2c, 32'hc31b71dd},
  {32'h437f0345, 32'h43459885, 32'hc29b0ad5},
  {32'h43a33f4a, 32'h4323c0a5, 32'h4228608c},
  {32'hc4b94380, 32'hc26388c3, 32'h428dbd69},
  {32'h4446cd48, 32'hc30312b0, 32'hc360b376},
  {32'hc4e013b1, 32'hc30461a3, 32'hc33e2b76},
  {32'h43da8aa6, 32'h43aa6dd7, 32'hc309b48c},
  {32'hc4cd07d1, 32'h42f2282b, 32'h41cca90c},
  {32'h43ecc7b5, 32'h435015d3, 32'h43f9da6c},
  {32'hc4bf1f32, 32'h424eb2e5, 32'hc3139dbf},
  {32'h45007f30, 32'h4313875b, 32'h42de21c0},
  {32'hc44ab376, 32'hc2667e64, 32'hc3b5ac95},
  {32'h450d7edb, 32'h432aa786, 32'h42b538cd},
  {32'hc4c7eda5, 32'h43a8d917, 32'h42d3774b},
  {32'h44a7940d, 32'h432e42fc, 32'hc308af1c},
  {32'hc4abbb6f, 32'hc2b5ae68, 32'h41b3dc56},
  {32'h42ff3050, 32'h4303bb43, 32'hc33a8a7f},
  {32'h41c040a4, 32'h43d44cfe, 32'h43084c5d},
  {32'h44bb5655, 32'hc325f44e, 32'h43c0f808},
  {32'hc4424ae4, 32'hc32f32c7, 32'hc2ae4a66},
  {32'h44cbb41f, 32'h4339351e, 32'h4356cb2a},
  {32'hc34a7808, 32'hc27d9ce4, 32'hc39d56e8},
  {32'h44ac74e5, 32'hc2fa4d0e, 32'hc36081f3},
  {32'hc511ae43, 32'hc38afdf3, 32'hc2d8bf95},
  {32'h4425911a, 32'h428829f2, 32'hc3da7f09},
  {32'hc50846ef, 32'h42de3415, 32'hc35da08d},
  {32'h450b8a86, 32'h4306da2a, 32'hc2b2a4bf},
  {32'hc4017fd0, 32'hc37ccff6, 32'hc399ed2c},
  {32'h444033f1, 32'h4314f192, 32'hc19f7675},
  {32'hc4f7f2d6, 32'hc2b99527, 32'hc33ea4b2},
  {32'h44845326, 32'h43e55eea, 32'h40b42943},
  {32'hc4a6dc3c, 32'h43d577e2, 32'hc38216f6},
  {32'h4457bdc0, 32'h41757f0f, 32'h4380e4d4},
  {32'hc4cc6a1a, 32'h43bdfcdb, 32'hc23f3f36},
  {32'h44aa022c, 32'hc04b32c2, 32'hc30654c5},
  {32'hc4a2543b, 32'h43484907, 32'h42346320},
  {32'h45130b5a, 32'hc361b091, 32'h4390cb76},
  {32'hc4e2719f, 32'h42d083b2, 32'h42af2cf5},
  {32'h438e03b0, 32'h41f29738, 32'hc21b79d4},
  {32'hc402d6a0, 32'h420255bb, 32'hc22eb3ac},
  {32'h44d63087, 32'h43bd68f4, 32'hc1c3862c},
  {32'hc4c3771e, 32'h42d53a18, 32'h430c82ac},
  {32'h43e6656a, 32'h43b4ab53, 32'hc3c7eb25},
  {32'hc4a482bb, 32'hc372e65c, 32'hc1901abc},
  {32'h44f82bbc, 32'hc361a1c4, 32'hc32fc2c6},
  {32'hc3cccbb0, 32'h4373c2fa, 32'h3d8e79e4},
  {32'h449b27c2, 32'hc318a6b0, 32'h432c8914},
  {32'hc471919e, 32'hc22407fe, 32'h4325dec5},
  {32'h4505b6c4, 32'h430719f4, 32'hc3aaafc9},
  {32'hc3e760d0, 32'hc3955057, 32'h43a023cf},
  {32'h450825c6, 32'hc4023be2, 32'hc2512016},
  {32'hc51d359a, 32'h435e2d6c, 32'hc3d12424},
  {32'h429aad50, 32'h43081e56, 32'h438cbb3e},
  {32'h41d16f00, 32'h435655ae, 32'h430922a9},
  {32'h450bc724, 32'h43a37652, 32'h430339d1},
  {32'hc38189f8, 32'hc2f443e7, 32'h426f8870},
  {32'h4524a9b0, 32'hc3070ae9, 32'h431dbc58},
  {32'hc4e25bd2, 32'h42ed4dfe, 32'hc375fbc6},
  {32'h44ab49c4, 32'hc2c9d000, 32'h4262dd8c},
  {32'hc4a724b1, 32'hc34df722, 32'hc36c08db},
  {32'h45024bcc, 32'hc3e716ac, 32'hc33c9f09},
  {32'hc4c08d44, 32'hc3813e82, 32'hc186180a},
  {32'h444396be, 32'h42c85b9c, 32'hc29bf31b},
  {32'hc504dbcb, 32'hc1896ef4, 32'hc045bffc},
  {32'h4478fe7e, 32'h419025d8, 32'hc337e3a3},
  {32'hc47d1c64, 32'hc335d0d5, 32'h42d1b676},
  {32'h43b2ead8, 32'hc20f9d14, 32'h42dc298d},
  {32'hc4a8b08e, 32'hc2fad2ee, 32'h43152814},
  {32'h44f784eb, 32'h433dc558, 32'hc26fa41a},
  {32'hc4ede4be, 32'h43837462, 32'h43b8c567},
  {32'h44adad45, 32'h43fece21, 32'h432924d9},
  {32'hc41a1dca, 32'hc11f2bec, 32'hc2b34d1e},
  {32'h44851c38, 32'hc358501f, 32'h4304fd3f},
  {32'hc50df1fa, 32'hc3160108, 32'h43343a4c},
  {32'h44c36f76, 32'h4344f7d4, 32'hc347a2a7},
  {32'hc3485ea6, 32'h43872bc2, 32'h430f2025},
  {32'h444b5990, 32'hc3a806e6, 32'hc0deddc4},
  {32'hc5066894, 32'hc395f165, 32'hc36e3729},
  {32'h45009706, 32'hc2fcc482, 32'hc2c28eda},
  {32'hc4dbf097, 32'h4148c92e, 32'h4169f818},
  {32'h445e3689, 32'h42b5201b, 32'h433a5163},
  {32'hc4ed70d6, 32'h43115759, 32'h43bf8036},
  {32'h447c885c, 32'h42e95ee9, 32'hc2a64677},
  {32'hc458c2a0, 32'h439ab645, 32'h432cb329},
  {32'h44ee1d08, 32'hc12cd9d6, 32'hc3d59067},
  {32'hc4b783ba, 32'hc16f5e69, 32'h43257bf2},
  {32'h4396840c, 32'hc113ad0c, 32'hc3b47237},
  {32'hc45365ea, 32'h43afde2c, 32'h43648b85},
  {32'h448ccf1b, 32'hbc5b9000, 32'h4300039d},
  {32'hc3fbb638, 32'h43aa70e6, 32'h428f951d},
  {32'h44d1948b, 32'h431198ef, 32'hc39f4ed2},
  {32'hc3b94f5f, 32'h42b8c6b1, 32'h4364ce56},
  {32'h446ac01a, 32'hc2ff824a, 32'h429990a4},
  {32'hc4400c33, 32'hc355dddf, 32'h43823703},
  {32'h44b4c305, 32'hc3dde435, 32'h43075564},
  {32'hc452b2b6, 32'h428985e9, 32'h433fc10f},
  {32'h44a7a4ef, 32'hc31354f9, 32'hc36ba1b4},
  {32'hc401deef, 32'h4323ffd3, 32'h4260517f},
  {32'h444a25a4, 32'hc298fcdf, 32'hc36d7043},
  {32'hc4c9c39e, 32'hc38235aa, 32'hc2a1e8cf},
  {32'h44ce3619, 32'h437a263e, 32'h42c009c0},
  {32'hc4d86662, 32'hc3edda29, 32'h43ed49f8},
  {32'h44a73ef9, 32'h43a8e8a2, 32'h4317169e},
  {32'hc32cf9e0, 32'hc31ea3df, 32'hc211674e},
  {32'h44b7c60a, 32'h43814070, 32'h43a37a73},
  {32'hc4bc98c6, 32'hc35d958c, 32'h4268cb0b},
  {32'h412bab00, 32'hc2e955d1, 32'hc2203833},
  {32'hc30c9f3a, 32'h43b4cd18, 32'hc3007fbe},
  {32'h44ec68da, 32'hc38ce838, 32'h43e595e7},
  {32'hc50705c1, 32'hc358b267, 32'h4378a353},
  {32'h4412d730, 32'hc30a3fb2, 32'hc2c95e57},
  {32'hc42101fa, 32'h41e008b2, 32'h4332dd1f},
  {32'h4507c556, 32'h427ca5a2, 32'hc1b32f06},
  {32'hc2681f20, 32'hc28b8d95, 32'hc36394bd},
  {32'h45005ceb, 32'h4323256f, 32'h4268348b},
  {32'hc4cb0bd2, 32'h42b0bbc7, 32'hc23d5371},
  {32'h45058e63, 32'hc0d2c9ea, 32'hc0e2e1ce},
  {32'hc4c95501, 32'h4287cfde, 32'hc2b7da40},
  {32'h44ed3845, 32'hc33169ff, 32'hc30e3e55},
  {32'hc4488dba, 32'h40eb1df3, 32'h43c7178a},
  {32'h4484e793, 32'hc10d91d9, 32'hc32c400d},
  {32'h43a15c75, 32'h430a9771, 32'h42ac7e18},
  {32'h449fe122, 32'hc25a4ba1, 32'hc395b360},
  {32'hc46e66ee, 32'hc213fda3, 32'h42ed6fc4},
  {32'h430dedd0, 32'hc3440471, 32'h4255f380},
  {32'hc4e9966e, 32'hc3a4110a, 32'h420d2a64},
  {32'h4215c5b0, 32'h42e0747d, 32'h4097bfe2},
  {32'hc5156ad3, 32'hc331489b, 32'hc20d39d2},
  {32'hc30f6d8c, 32'h4404454f, 32'hc34566da},
  {32'hc3926562, 32'h414cb46f, 32'h41c216d2},
  {32'h451a16d0, 32'h4332acfa, 32'hc25fce10},
  {32'hc48180f5, 32'hc31ee6e9, 32'h431f1ece},
  {32'h4520482c, 32'hc29bbc05, 32'h435ae26f},
  {32'hc4d167a8, 32'hc2cb68c4, 32'hc3610200},
  {32'h44d868bf, 32'h42bd5a78, 32'h431d3ee4},
  {32'hc4489e2a, 32'h430646a4, 32'hc3a9174c},
  {32'h44d1e718, 32'h43422e16, 32'h43c237d5},
  {32'hc4746258, 32'hc31e7949, 32'hc36bdaf6},
  {32'h4501ce12, 32'hc31bb1d6, 32'h4388ede1},
  {32'hc4f2f1bc, 32'h433c9404, 32'h43014f33},
  {32'h42c3d2b0, 32'hc3ef0390, 32'hc34ab336},
  {32'hc4d41626, 32'hc344f388, 32'h43a17821},
  {32'h442e4566, 32'h436f9ff2, 32'hc33e6579},
  {32'hc4a84102, 32'hc205c5d8, 32'hc22379c2},
  {32'h44938280, 32'hc25a8af2, 32'h42a9af9a},
  {32'hc44c6e1e, 32'hc2933d64, 32'hc393ff24},
  {32'h43871b16, 32'hc355f2aa, 32'hc08c9146},
  {32'hc4dcc9ec, 32'hc28990fb, 32'hc3416d90},
  {32'h4408b834, 32'h4226558b, 32'h42bab3d1},
  {32'hc40b6134, 32'hc346cc86, 32'hc35f4e7a},
  {32'h4455d188, 32'hc2f3e99f, 32'h42a58e63},
  {32'hc485aaa0, 32'h42b5ef71, 32'h436c63d0},
  {32'h44c55704, 32'hc2faf1c2, 32'h43856ec0},
  {32'hc4b438b8, 32'hc1ed1dc0, 32'h41cab890},
  {32'h4507e64a, 32'hc377d90e, 32'hc3d9dacd},
  {32'hc4249ca2, 32'h43a90e78, 32'hc402dac8},
  {32'h444093d4, 32'hc30307ef, 32'hc1fbbc88},
  {32'hc49054e1, 32'hc30e15c5, 32'h439f0af7},
  {32'h44fd69df, 32'h43d2b14a, 32'h42f1cc53},
  {32'hc4123f50, 32'h42683b02, 32'hc3a963c4},
  {32'h4400bc52, 32'h43022ee7, 32'h42a73ab6},
  {32'hc4959f9e, 32'h42f3192a, 32'h41e40109},
  {32'h4507512c, 32'h40fd6d76, 32'h42f9f8be},
  {32'hc4a0e725, 32'h439a675f, 32'h4401a300},
  {32'h4490ab78, 32'h42d56022, 32'hc22d32d3},
  {32'hc4c24650, 32'hc2af157f, 32'h4134f5e0},
  {32'h44dbaeb8, 32'hc26df888, 32'h4169130b},
  {32'hc49ada4c, 32'hc31a6a14, 32'h43444abd},
  {32'h43e2dbb8, 32'hc3728ac6, 32'hc2235822},
  {32'hc4d65e3f, 32'h42f18847, 32'h43ada885},
  {32'h44395074, 32'hc225e355, 32'h43963780},
  {32'hc397cb68, 32'hc3976013, 32'h435ab0be},
  {32'h4462ff36, 32'hc31c759c, 32'hc3b5ecfb},
  {32'hc4445389, 32'hc142791c, 32'h4301b95d},
  {32'h4479cfd8, 32'hc34075ed, 32'hc304fc5e},
  {32'hc28d2030, 32'hc3f9afe8, 32'h431987c1},
  {32'h43cc919c, 32'hc3036c1f, 32'h43c1c000},
  {32'h42ef8bde, 32'hc21722a5, 32'h433f85cc},
  {32'h44f2f246, 32'h43da3b13, 32'hc363d8bd},
  {32'hc4da6f75, 32'hc2f9ec70, 32'h434153f8},
  {32'h43547be8, 32'h437af058, 32'h420211bb},
  {32'hc3427884, 32'h42ea2244, 32'hc0ccb6d4},
  {32'h44db8d50, 32'h4375a25b, 32'hc2bb6109},
  {32'hc4f2e1d2, 32'hc323a3fb, 32'hc26162d2},
  {32'h4508d2c7, 32'h42a0fc3a, 32'hc37e0151},
  {32'hc48800f6, 32'hc32714ab, 32'h431941a3},
  {32'h44de1038, 32'hc3113e79, 32'h42273387},
  {32'hc4bf6514, 32'hc2fd1b11, 32'h41e26a0e},
  {32'h44b3be1c, 32'h434b02e6, 32'hc406daff},
  {32'hc4bdfeb0, 32'h407be609, 32'h4204b158},
  {32'h4311f380, 32'h3f46a8e0, 32'hc2b98af7},
  {32'hc498ac37, 32'hc38c4e02, 32'h4208b577},
  {32'h4511b494, 32'h41af09d6, 32'hc3454ff3},
  {32'hc49c68ae, 32'hc3887a3f, 32'hc379ba2d},
  {32'h445c8e9c, 32'h43a03da1, 32'hc25513c9},
  {32'hc5029bf3, 32'hc2e6bfe8, 32'h43aec04c},
  {32'hc2fd7800, 32'h429f6d5b, 32'hc3aa5a06},
  {32'hc50c45b9, 32'hc34d5f20, 32'hc20f325d},
  {32'hc2f04390, 32'hc26cba76, 32'hc1ccfe06},
  {32'h42b1aa4f, 32'h43324bcd, 32'hc2ffa1d4},
  {32'h448c1667, 32'hc34b0f88, 32'h4230954d},
  {32'hc3ca546a, 32'hc213c732, 32'hc3450448},
  {32'h444850ea, 32'h43b5c131, 32'hc0874dca},
  {32'hc4d59012, 32'h43846a03, 32'h42f1947d},
  {32'h44509eaa, 32'h41ce42aa, 32'h42347c11},
  {32'hc2fc6de0, 32'hc26fe866, 32'hc11de2fc},
  {32'h44e18b77, 32'h43941d4b, 32'hc36f98f5},
  {32'hc41e8bfa, 32'h435f3ab3, 32'hc352196f},
  {32'h449b4110, 32'h43949c45, 32'hc383e8ee},
  {32'hc2c76bc0, 32'h430273b4, 32'hc38274e9},
  {32'h43c96bfc, 32'hc33d608a, 32'hc2bd8d73},
  {32'hc4b72712, 32'hc37216c1, 32'h421a1c10},
  {32'h446cca80, 32'hc3744718, 32'hc39b5573},
  {32'hc4a6fd6b, 32'h42eea83e, 32'hc225935c},
  {32'h44fe0873, 32'h42dd53c2, 32'hc3aeb3e0},
  {32'h42fbeb5d, 32'hc2ba759b, 32'h43bacdfe},
  {32'h44e3c74e, 32'hc26a47c1, 32'hc2b43847},
  {32'hc44790a4, 32'h422b3c9e, 32'hc292bc76},
  {32'h44fc3737, 32'h43dd2fa5, 32'hc345c5b0},
  {32'hc4a00dba, 32'hc3b2df85, 32'hc1febfae},
  {32'h44ee8340, 32'h41acb484, 32'h42606955},
  {32'hc3aac3b0, 32'h43df55b4, 32'h4344e068},
  {32'h44c11fa2, 32'hc3aa5830, 32'h42957835},
  {32'hc4e8ab52, 32'h430bf5d2, 32'hc10d3ba1},
  {32'h4328ff8c, 32'h41dc6a4f, 32'h43843b3a},
  {32'hc427bb18, 32'hc378daa8, 32'hc3b39c22},
  {32'h449bf722, 32'hc3881d76, 32'h423908a4},
  {32'hc4124406, 32'h4298a783, 32'h43d1b2d0},
  {32'h44cb8a22, 32'hc34e39b6, 32'hc1ba742e},
  {32'hc49f7e0e, 32'hc320825d, 32'h4320bfdb},
  {32'h44f4ac1c, 32'hc2c283a3, 32'h43689fb1},
  {32'hc4abccde, 32'hc2969e7a, 32'hc36398c4},
  {32'h44d5dc74, 32'hc4046a79, 32'h4340e891},
  {32'hc4306cfb, 32'h438d8363, 32'h42e6c88e},
  {32'h44b66d62, 32'hc2cc0ff7, 32'hc3f9c09a},
  {32'hc39dbb02, 32'h42817f52, 32'h41b4bd09},
  {32'h4517deaa, 32'h43552516, 32'hc3c9a267},
  {32'hc4557fe8, 32'h429c9e42, 32'hc0b30b22},
  {32'h44f5ec1e, 32'hc3be26cd, 32'hc1061896},
  {32'hc50132c7, 32'hc38ffe8f, 32'hc250a4e2},
  {32'h44a55824, 32'hc2a8a2ad, 32'hc22cfb5c},
  {32'hc4832898, 32'hc3d20d43, 32'hc30d92db},
  {32'h44b9eb4d, 32'hc39d596f, 32'hc20c45cf},
  {32'hc436b7f6, 32'hc3814043, 32'hc170cc47},
  {32'h4499af8b, 32'hc2d49656, 32'h42fa9e8b},
  {32'hc4af2744, 32'hc2cdfa49, 32'hc2db3d93},
  {32'h43da2a58, 32'h428395aa, 32'hc2189bf2},
  {32'hc5148378, 32'hc29e8f54, 32'hc24505f4},
  {32'h44bb2911, 32'hc43bd037, 32'h42f62311},
  {32'hc493f032, 32'hc294c8c7, 32'hc388d745},
  {32'h4403400c, 32'h41511137, 32'h427624f9},
  {32'hc502a3a4, 32'hc33edb72, 32'hc341d41d},
  {32'h4511f332, 32'hc29d8b57, 32'hc384ae23},
  {32'hc4bdfc04, 32'hc30dfcf9, 32'hc19041c4},
  {32'h450ddaa5, 32'h434f7750, 32'h41c82b4a},
  {32'hc4342140, 32'h40a71ffa, 32'h42dc75a6},
  {32'h44c03e1b, 32'hc3d02672, 32'h437ab421},
  {32'hc3d21e4c, 32'hc0ae886f, 32'h43f0edfd},
  {32'h4402ea8c, 32'hc3275edd, 32'h42ed2c38},
  {32'hc5040c86, 32'hc22c09b7, 32'hbf4b2ac0},
  {32'h449aac48, 32'hc2d37d38, 32'h42145b74},
  {32'hc4f35a68, 32'hc21f06e0, 32'h43bfb4f5},
  {32'h44e64eff, 32'hc3d5d076, 32'h43841a71},
  {32'hc4d15d48, 32'h431820c1, 32'hc22f6307},
  {32'h44265969, 32'h404c86cb, 32'h41b3c614},
  {32'hc47a54e0, 32'h4126cdfc, 32'h4306ea78},
  {32'h44832b2d, 32'h424e24c4, 32'h43125acf},
  {32'hc4359e71, 32'hc3870712, 32'hc2dc790a},
  {32'h44da517d, 32'h42fe1840, 32'h43783924},
  {32'hc43b567a, 32'hc2c7b268, 32'h42ff993c},
  {32'h4504c980, 32'h428faf5c, 32'hc2f67b83},
  {32'hc45ee62c, 32'hc15f8150, 32'h42f86fa1},
  {32'h44ff3865, 32'hc3c45806, 32'h42fb4644},
  {32'hc4bc3cc4, 32'h4312b46e, 32'h42a28653},
  {32'h452062bd, 32'h43244d3e, 32'h42dcf7aa},
  {32'hc4836110, 32'hc08bf7c8, 32'h439a6b7c},
  {32'h44883e18, 32'h42d6a18d, 32'hc31ba626},
  {32'hc48e8d40, 32'h43eb8540, 32'h43346948},
  {32'h44db13d4, 32'h4211bb08, 32'hc2d0fe9d},
  {32'hc477510a, 32'h439d5686, 32'hc1c6bbfe},
  {32'h44b11f98, 32'hc2632a64, 32'hc34f06a8},
  {32'hc3c15eb4, 32'hc30edf84, 32'hc2779f49},
  {32'h44170787, 32'hc42821b0, 32'h433fba2b},
  {32'hc5004ab8, 32'hc20f2c88, 32'hc4148345},
  {32'h44066de0, 32'h42d7f6cc, 32'hc362a783},
  {32'hc4b873ae, 32'hc2916e72, 32'h436adbfc},
  {32'h44b35883, 32'hc28afcc2, 32'h438bf4b5},
  {32'hc51a053a, 32'hc31c6bca, 32'h4348d98b},
  {32'h449638b0, 32'hc330358e, 32'h3f9fffa6},
  {32'hc49d8e6b, 32'hc35a69c5, 32'h429b1aa7},
  {32'h44c93ab6, 32'h41909799, 32'h435cb7dd},
  {32'hc4e16cd5, 32'hc1d9d560, 32'hc2fe4f45},
  {32'h44f99556, 32'h4284c8ac, 32'h431984ba},
  {32'hc4b33764, 32'hc1d071e6, 32'hc399276b},
  {32'h446b7488, 32'h4398a6b5, 32'h43af8a45},
  {32'hc4075a4c, 32'h42769abd, 32'h43a62b23},
  {32'h4512d6a1, 32'h43bca91a, 32'hc198d1f1},
  {32'hc48466f4, 32'h41196264, 32'hc38fd834},
  {32'h44b00ef2, 32'hc2ddf737, 32'h43677889},
  {32'h42442160, 32'hc305a310, 32'hc2c50c63},
  {32'h449d73b2, 32'hc1caeb06, 32'h421e08d8},
  {32'hc511e539, 32'hc2c82ca3, 32'h433c26a9},
  {32'h44cccf20, 32'h439cf3d5, 32'hc1c67548},
  {32'hc40bf098, 32'hc240eab3, 32'hc290f6a6},
  {32'h444924b2, 32'hc2f354f6, 32'h43805e9f},
  {32'hc313ae7f, 32'h42c642fc, 32'h432f0b18},
  {32'h451263ef, 32'h429382d8, 32'h43fa629f},
  {32'hc4716712, 32'h425a357b, 32'h439354e8},
  {32'h45296e64, 32'h42958631, 32'h43afa5b8},
  {32'hc2dedc5a, 32'h4359dd16, 32'h4394dd19},
  {32'h4299da13, 32'h43b00752, 32'hc3f295ac},
  {32'hc3201800, 32'h4331dfd8, 32'h42f1939d},
  {32'h450fc31b, 32'hc1d30a14, 32'h432b2415},
  {32'hc4a797d5, 32'hc3808ada, 32'h4311d210},
  {32'h446513d7, 32'h432036b0, 32'hc2cfe55f},
  {32'hc4b04705, 32'hc34fc1b2, 32'hc2b105c2},
  {32'h43fbb1f8, 32'h432e8d90, 32'h42c278f1},
  {32'hc496be56, 32'h41f7c642, 32'h4323af52},
  {32'h44b5293e, 32'hc26372d2, 32'hc2f765d6},
  {32'hc4311af0, 32'h4373fb79, 32'h4342f9dc},
  {32'h43a02c9e, 32'h4320046f, 32'hc3408e75},
  {32'hc4233b62, 32'h4359c363, 32'hc399a12b},
  {32'h44af8cb4, 32'h43a5f3d3, 32'hc090d817},
  {32'hc483fd42, 32'h438b1ea3, 32'h4374eafc},
  {32'h43bb1c8f, 32'h4381b0ce, 32'hc309dca2},
  {32'hc50ef11b, 32'h431fdbe9, 32'hc3c766a5},
  {32'h42af06e0, 32'h433ef8b9, 32'hc35353be},
  {32'hc3d3bf50, 32'h42db62a8, 32'hc1db5205},
  {32'h44703446, 32'hc340ac14, 32'hc2ea180b},
  {32'hc4c459e6, 32'h43a6f07d, 32'hc1bd01f8},
  {32'h449a7fb6, 32'hc3921886, 32'h4374310f},
  {32'h4399b4f0, 32'h4311a670, 32'h42531a35},
  {32'h4486b4cb, 32'h42fc96f3, 32'hc35c8c2f},
  {32'hc4e9746e, 32'h42966092, 32'h43846a24},
  {32'h44f5396f, 32'hc34d249b, 32'hc30349c4},
  {32'hc4fd6be2, 32'hc3560d01, 32'h4308b3b1},
  {32'h44fa55e2, 32'h43659e65, 32'h43172156},
  {32'hc32a1a72, 32'h438a5293, 32'h4327f495},
  {32'h44f10046, 32'h3ffcd8b0, 32'h4266d5f7},
  {32'hc4a4bd8a, 32'hc40513e3, 32'h43243f9d},
  {32'h44fd1bf4, 32'hc30a1ea0, 32'h435f813f},
  {32'hc3ff12cd, 32'h434a0b3c, 32'hc209ea91},
  {32'h44b982a1, 32'h41b67730, 32'hc30cbb74},
  {32'hc4be6027, 32'hc36625f3, 32'h4171a097},
  {32'h44e10f3a, 32'h43ae864b, 32'hc35162cb},
  {32'hc498533f, 32'hc36e00db, 32'h4331795d},
  {32'h44c4bd09, 32'h433bebff, 32'h432a7669},
  {32'hc477f8a0, 32'h43a249cb, 32'hc32846bd},
  {32'h4394ece2, 32'hc40bfffe, 32'hc1045fbd},
  {32'hc4579ce8, 32'h43eac1dc, 32'hc1c4c5cd},
  {32'h44d27987, 32'h43afb486, 32'hc24faffe},
  {32'hc3876153, 32'h4356b543, 32'h43140869},
  {32'h4505ee21, 32'h43bc8e22, 32'hc2f614ca},
  {32'hc3e0efe0, 32'hc1b6dbf1, 32'hc325e2e9},
  {32'h44f02d6a, 32'h4262e84f, 32'h408002a1},
  {32'hc512233a, 32'hc2676d69, 32'hc3bda703},
  {32'h44a8c500, 32'h4246e170, 32'h429d1a56},
  {32'hc4ca9216, 32'h4383a102, 32'h4181e8bf},
  {32'h44892335, 32'hc2d290c6, 32'h43648397},
  {32'hc42e02f5, 32'hc3619fe9, 32'h440c8759},
  {32'h448e1a5a, 32'hc3b883a4, 32'hc34b6895},
  {32'hc461e807, 32'hc25bf0b0, 32'hc2aeeaf9},
  {32'h4484f914, 32'h4278d704, 32'h421352f4},
  {32'hc4d15796, 32'h42947fe6, 32'h435dc8b9},
  {32'h450f03ff, 32'hc40a701d, 32'h4168db90},
  {32'hc481b05c, 32'hc10217dc, 32'hc308277b},
  {32'h44767878, 32'hc2f5c297, 32'hc2d84add},
  {32'hc4ff1fc7, 32'h431b31a4, 32'h4336aced},
  {32'h4447a822, 32'hc36dcfdc, 32'h4396c593},
  {32'hc4ee943c, 32'hc37ef47d, 32'h4152d131},
  {32'h441a5122, 32'h41e33680, 32'h42c739c4},
  {32'hc40c6e1b, 32'h4359457a, 32'h42218b6e},
  {32'h4486fcc1, 32'h436339e5, 32'h4371de18},
  {32'hc30fb0c8, 32'h42ff7ac4, 32'hc1acd62e},
  {32'h44938bea, 32'h4258fcc8, 32'h43538bb8},
  {32'hc48da179, 32'h4104113d, 32'hc3296e31},
  {32'h4484cccc, 32'hc24a13c1, 32'hc3cc388e},
  {32'hc438acd6, 32'h42f03a82, 32'hc17475a4},
  {32'h4501f7d4, 32'hc3cf8b18, 32'hc3687734},
  {32'hc4972815, 32'h40d72673, 32'h434917fe},
  {32'h448d7700, 32'h437ceaae, 32'hc309c20d},
  {32'hc4e4f9a4, 32'hc34297d3, 32'hc3645a86},
  {32'h44e610aa, 32'hc35e876e, 32'h4205bf15},
  {32'hc4c5b4dc, 32'h43a1e05f, 32'hc3bdfe31},
  {32'h43a3be16, 32'hc1eb0d4c, 32'hc3285933},
  {32'hc5023dca, 32'hc32e1bd5, 32'h4186b59e},
  {32'h44d1077e, 32'hc3a8365b, 32'h42b7429f},
  {32'hc3f5251e, 32'h43180370, 32'h42a4c5ba},
  {32'h44d1c7fa, 32'h42c7975d, 32'h42cedb14},
  {32'hc4f14618, 32'hc1e303cc, 32'hc384d000},
  {32'h44a346e5, 32'h41adcec6, 32'h42ae189c},
  {32'hc3657b50, 32'h42b0bac1, 32'hc14d26b6},
  {32'h43ed9dac, 32'h431a88dd, 32'hc1979e26},
  {32'hc504559a, 32'hc2e3ba47, 32'hc30fe51e},
  {32'hc3070556, 32'hc3b44052, 32'h40ec598c},
  {32'hc49469ac, 32'h42505a56, 32'h42f1b371},
  {32'h45047856, 32'h42984bc5, 32'h4017fb36},
  {32'hc4be7ea4, 32'hc2585faa, 32'h42bcae86},
  {32'h4464156e, 32'hc2ce6243, 32'hbfd83150},
  {32'hc4d229ca, 32'h42ff91aa, 32'h4356b642},
  {32'h44fed513, 32'hc355b2e1, 32'hc2c67726},
  {32'hc4bb3d2a, 32'hc299e9f7, 32'h420ac1e6},
  {32'h44c6b910, 32'h42583196, 32'hc34fdb19},
  {32'hc30e2770, 32'h435fd857, 32'hc2669eb2},
  {32'h44e9c8e1, 32'hc31c78cc, 32'hc2343150},
  {32'hc34436a0, 32'hc394d8ef, 32'hc1d7a978},
  {32'h44b83645, 32'hc2cb21c6, 32'hc39847f1},
  {32'hc42df0f2, 32'h4310895d, 32'h4361ec7b},
  {32'h44adf65a, 32'hc35bf3c5, 32'hc2ff8ebe},
  {32'hc2bb2340, 32'hc3688569, 32'hc220cdca},
  {32'hc508fe11, 32'h43944876, 32'hc3e3c815},
  {32'h44fc291a, 32'h434aae35, 32'h43a4a58b},
  {32'hc4c5d210, 32'h41f966fe, 32'h42beaa4d},
  {32'h44294ed7, 32'hc3672ea4, 32'h43656ff4},
  {32'hc4e9bc74, 32'hc10d235b, 32'h41e05e0e},
  {32'h44d9617a, 32'h433b335b, 32'hc3e07de4},
  {32'hc46b355c, 32'hc1dca2da, 32'hc2c64bba},
  {32'h450437ce, 32'hc0896bc4, 32'h4184958b},
  {32'h4365e4cd, 32'hc37ad05a, 32'h43b1f2e2},
  {32'h44e9026c, 32'h4344067e, 32'hc3a969af},
  {32'hc4da3e55, 32'hc237c473, 32'h433989c6},
  {32'h447b6b95, 32'hc36091ad, 32'h43851b72},
  {32'hc4b72beb, 32'hc30ca474, 32'hc339dc84},
  {32'h45188f0d, 32'h4365ab33, 32'h42fb7767},
  {32'hc4fec942, 32'h42073997, 32'h4345ee40},
  {32'h42bef610, 32'h42bf3e03, 32'h4365ec15},
  {32'hc48a7afb, 32'h42bc9d20, 32'h42a10bf7},
  {32'hc306e090, 32'hc2968095, 32'hc325e4c0},
  {32'h42cc8fe0, 32'h42f57bbd, 32'hc3070f70},
  {32'h43f0b4d7, 32'h436521e6, 32'h434de1ae},
  {32'hc44bfb98, 32'h42ff36b5, 32'h41d5cca9},
  {32'h41a7e090, 32'hc2b6d5a4, 32'hc28fbd66},
  {32'hc3a8627a, 32'hc3cecc5a, 32'h43705f15},
  {32'h439f5829, 32'hc2dea0a0, 32'hc3f17928},
  {32'hc4c96295, 32'hc388f1ec, 32'h41ac4168},
  {32'h44f56bca, 32'h4374724a, 32'hc374e006},
  {32'hc4e3a8ba, 32'hc3143a49, 32'hc303c8e2},
  {32'h44a705d8, 32'h4396bd4c, 32'h43a22f1f},
  {32'hc45810a0, 32'hc29ec726, 32'hc3a8aa1e},
  {32'h44f31a23, 32'h43066dd8, 32'h42127962},
  {32'hc43f3e54, 32'hc3cb0098, 32'h43433fef},
  {32'h4406c936, 32'hc3827602, 32'h427f85de},
  {32'hc502714e, 32'h42f40ff3, 32'hc3950dc6},
  {32'h44c38846, 32'h42bfa59b, 32'hc1926f35},
  {32'hc22669c0, 32'hc2950edd, 32'h4381d9fd},
  {32'h43fd477a, 32'h40de65e5, 32'hc2e203a2},
  {32'hc4f7773a, 32'h43b52c3d, 32'h438c056b},
  {32'h443217d4, 32'h43069dd7, 32'h43454cb6},
  {32'hc504db9a, 32'h43c45925, 32'hc325f477},
  {32'h44cd394e, 32'hc1ca8f53, 32'h43aa2f4d},
  {32'hc4dc6e40, 32'h43a08bc6, 32'h40c595cf},
  {32'h44b4bf7a, 32'h42aa6e5d, 32'h43dcb429},
  {32'hc4340eae, 32'h4272d594, 32'h4359da12},
  {32'h44bade73, 32'hc302f471, 32'hc2ed4623},
  {32'hc4538dac, 32'h42ec274b, 32'hc2c7be47},
  {32'h44f2c5c4, 32'h4256e290, 32'hc1a30fb2},
  {32'hc41b5a4c, 32'h43026004, 32'h438a67f3},
  {32'h447b0140, 32'hc285c3b6, 32'hc17cfadf},
  {32'hc4239402, 32'h4296e516, 32'hc22a26a4},
  {32'h44944226, 32'h426efd07, 32'hc2912b3b},
  {32'hc4b2a2ea, 32'h43c2a686, 32'hc13dec08},
  {32'h44ba5c34, 32'hc3b75f2f, 32'hc30ab42f},
  {32'hc3984e98, 32'h428ad226, 32'hc39ce4ad},
  {32'h43ef29fa, 32'h4368ed20, 32'hc33f68fe},
  {32'hc40ebcd4, 32'h42192af0, 32'hc3bf2753},
  {32'h443ae36b, 32'h432d3eef, 32'hc2108e5a},
  {32'hc3fa277c, 32'h42f210e9, 32'hc31e43f4},
  {32'h45146fdb, 32'hc314f517, 32'hc3cefbb6},
  {32'hc48e6411, 32'hc1c076ac, 32'hc398992b},
  {32'h44927f53, 32'hc3671bfb, 32'h41db54a1},
  {32'hc4a78fca, 32'hc3851949, 32'hc3656d81},
  {32'h443b58e8, 32'hc39acef9, 32'hc2c67d89},
  {32'hc4d103f6, 32'hc05798c0, 32'hc0c8b1a0},
  {32'h43ee7d80, 32'hc3634534, 32'h41297ee4},
  {32'hc46fd6ce, 32'h4331626a, 32'h440c6f44},
  {32'h44ad28c3, 32'hc0e60c95, 32'hc12b34d0},
  {32'hc4e260c9, 32'hc35a00c4, 32'hc383673a},
  {32'h44948f28, 32'h4353aff2, 32'h42d7f5a5},
  {32'hc468c892, 32'hc3877d6c, 32'h4221a707},
  {32'h44c44f32, 32'h4406dfd4, 32'h410d7d85},
  {32'hc440446c, 32'hc3969dfc, 32'h424b4eae},
  {32'h445dbcb6, 32'h421bce38, 32'h431c4c83},
  {32'hc4a6c21d, 32'hc333ca63, 32'h43bc5782},
  {32'h44047674, 32'h43562836, 32'h43a8f2c9},
  {32'hc4e10483, 32'h42063bd5, 32'hc21473c8},
  {32'h446c2c92, 32'h42e8bd9d, 32'h4191f233},
  {32'hc4a25461, 32'h4365d50f, 32'hc2494246},
  {32'h44bb78b0, 32'h439e5b9c, 32'h430d3dbf},
  {32'hc4371f7d, 32'hc39b2a56, 32'hc1539376},
  {32'h4503acc7, 32'hc3157bcc, 32'h42a076b3},
  {32'hc4a25d1a, 32'h43ae59cd, 32'hc2baf8fa},
  {32'h44ffbe2b, 32'hc301a684, 32'h43ef683a},
  {32'hc511943c, 32'h42a3733d, 32'hc1a328c0},
  {32'h4430f23e, 32'hc32935d1, 32'hc1c95ec9},
  {32'hc485313f, 32'hc33ab78d, 32'h41bb52d4},
  {32'h44871f92, 32'h4390f7fb, 32'hc3dba4a8},
  {32'hc4e55a52, 32'hc39bce10, 32'hc405cb4d},
  {32'hc215c080, 32'hc2c5aa7e, 32'hc2abcb17},
  {32'hc4a5b124, 32'h41583c10, 32'h41d2006d},
  {32'h44c797d9, 32'h4309a2de, 32'h42fb7655},
  {32'hc476f792, 32'hc3310763, 32'h41ba6417},
  {32'h43d548dc, 32'hc2d0061a, 32'hc3a18743},
  {32'hc4ecc298, 32'h4372c19f, 32'h431d6121},
  {32'h4513e464, 32'h437a439c, 32'hc3aaef5a},
  {32'hc457065c, 32'hc174bd8a, 32'h44039487},
  {32'h4508b4bb, 32'hc2efe860, 32'h441e381c},
  {32'hc50758b5, 32'h42f3d8f3, 32'h42b6bb72},
  {32'h452017f1, 32'hc34ba1c4, 32'hc27cf0b0},
  {32'hc4f816e4, 32'hc3496c6d, 32'h43934cdd},
  {32'h450fbf16, 32'h426ac668, 32'hc2ff3c2f},
  {32'hc49623ca, 32'hc32e8300, 32'hc0fa6fc3},
  {32'h43ad1455, 32'h43f5d205, 32'hc3f780d7},
  {32'hc4ba9ef9, 32'hc286200c, 32'h420b32b1},
  {32'h44c3f985, 32'hc32abaa6, 32'h437d4874},
  {32'hc4681dc0, 32'hc1df94ec, 32'h40d40c6c},
  {32'h44060e2f, 32'h42e93958, 32'h421f12e4},
  {32'hc50f3c22, 32'hc3853ae3, 32'h42940c70},
  {32'h44f024f5, 32'h4394f4f5, 32'h431d1ac3},
  {32'hc425ba9a, 32'hc2937da8, 32'hc32d4450},
  {32'h4497b5f2, 32'h4388fa75, 32'hc1f3aed1},
  {32'hc51df835, 32'h43d6d5dc, 32'h43b16bf4},
  {32'h451a2373, 32'h433a6027, 32'h4379311a},
  {32'hc4febc30, 32'h43acc636, 32'h433fd999},
  {32'h44846844, 32'h43562166, 32'hc34fc7d2},
  {32'hc503cc2e, 32'h41242d73, 32'h422f3125},
  {32'h438f062d, 32'hc3cab64f, 32'hc3c0dac0},
  {32'hc5165bd0, 32'hc32f6d6f, 32'h4321405f},
  {32'h43f64336, 32'hc19bc2b2, 32'h42be266e},
  {32'hc3bc26bb, 32'h431456c0, 32'hc38f4469},
  {32'h4493aad6, 32'hc3133384, 32'h43ebae29},
  {32'hc4c282cb, 32'hc3a20183, 32'h43cb5e1e},
  {32'h44e05ec8, 32'hc3271e3e, 32'h42c53b10},
  {32'hc4a33a6f, 32'h4231d7fe, 32'h43aae89f},
  {32'h44a2bcae, 32'hc39ad5a3, 32'hc3927464},
  {32'hc426a9d8, 32'hc3269dc1, 32'hc33002d0},
  {32'h44a71acb, 32'h42843f66, 32'hc30c2d15},
  {32'hc4cdadf1, 32'hc3b3b502, 32'hc24fc5d7},
  {32'h431afdfe, 32'hc2b2a924, 32'hc358a75a},
  {32'hc40beaad, 32'h43e8d758, 32'h43636a1c},
  {32'h44b58b6a, 32'hc320dd09, 32'h43003ca8},
  {32'hc2fc1958, 32'h430ea429, 32'hc32782c2},
  {32'h442a4424, 32'h425a808b, 32'hc20424d2},
  {32'hc31668b0, 32'hc30fc293, 32'hc28e0b13},
  {32'h44db5460, 32'h438be474, 32'h43b679cd},
  {32'hc18c4840, 32'hc3929aaf, 32'h4190ecd7},
  {32'h44935376, 32'h436d164e, 32'h42250a40},
  {32'hc402895e, 32'h42b0c959, 32'hc2ab9641},
  {32'h452eec5c, 32'hc34e249f, 32'h429128dd},
  {32'hc4a9c5d8, 32'h42787ad5, 32'h42ad09f7},
  {32'h43f6f494, 32'h42eef661, 32'h4344ebba},
  {32'hc49d5671, 32'h433949b2, 32'h43741fe7},
  {32'h4459cf32, 32'h43a5f5eb, 32'hc30c2917},
  {32'hc4b455d9, 32'hc2bbeb8c, 32'hc2de467e},
  {32'h449042e7, 32'h4385936c, 32'h4362884a},
  {32'hc511bdc2, 32'h4325480c, 32'h4340d969},
  {32'h43181c24, 32'hc31bdb2d, 32'h4236e277},
  {32'hc4ed3685, 32'h42b8ec39, 32'hc2ca59c3},
  {32'h4448c394, 32'h42ab62b1, 32'hc27a8e7b},
  {32'hc34b4da0, 32'hc2c28838, 32'hc3e70c3f},
  {32'h45177b9c, 32'h42b9517f, 32'h42dc6824},
  {32'hc314833a, 32'hc2b58213, 32'h435104fb},
  {32'h44cb0f3a, 32'hc382ff93, 32'h42e4c8c8},
  {32'hc4a67983, 32'h43807e90, 32'h44101f74},
  {32'h45088957, 32'hc33697e7, 32'h42f6d316},
  {32'hc5094938, 32'h430b2235, 32'hc1a43e13},
  {32'h440e8a76, 32'hc3470be6, 32'h42808148},
  {32'hc474ef97, 32'h42f59daa, 32'h42c2e94c},
  {32'h44313153, 32'h41815783, 32'hc3f92bfb},
  {32'hc4494d82, 32'h42bd93ff, 32'h43af0a7a},
  {32'h44f30737, 32'hc2ba78e5, 32'h43955195},
  {32'hc412ed68, 32'hc3926b2f, 32'hc181703f},
  {32'h44cf0ee8, 32'h43485103, 32'h43e569b9},
  {32'hc3e6289e, 32'h433d0118, 32'hc3011d18},
  {32'h452228aa, 32'h433362df, 32'hc3334565},
  {32'hc4c2016a, 32'h433458a4, 32'hc285e1f6},
  {32'h4444133e, 32'hc3931880, 32'hc3155d04},
  {32'hc365e0c0, 32'hc1a3a9d3, 32'h424ead57},
  {32'h44080d07, 32'hc1b0668e, 32'hc3b6bf22},
  {32'hc49849d2, 32'hc3da57a6, 32'h42f75252},
  {32'h434f4788, 32'hc326a138, 32'hc39802ee},
  {32'hc4bf75b2, 32'hc390d578, 32'h41be2a9e},
  {32'h441994be, 32'h43798f96, 32'h42a14bfb},
  {32'hc3b504a7, 32'hc29ab28c, 32'hc35641fd},
  {32'h44efddae, 32'hc28b2c26, 32'h42998e2b},
  {32'hc4427281, 32'h42cf056b, 32'hc25732d7},
  {32'h44f4d137, 32'hc38c79c8, 32'h43984230},
  {32'hc3c43aa4, 32'h42968bdd, 32'hc24cfd43},
  {32'h44968cd2, 32'h42e38a0c, 32'hc3a0e955},
  {32'hc50092f3, 32'hc3f85820, 32'h4305b479},
  {32'h44189e4f, 32'h439b07d2, 32'hc33e0633},
  {32'h42d18ce5, 32'hc2e4ca3b, 32'hc30f34ef},
  {32'h44b8c3fe, 32'hc1f2cc50, 32'h4209be8f},
  {32'hc4fc841c, 32'h428a960c, 32'hc32d36ed},
  {32'h4410fd82, 32'hc31f6c45, 32'h432e96fb},
  {32'hc4c639ef, 32'h421d9c07, 32'hc32e4db4},
  {32'h440de4a7, 32'h42c761c0, 32'h43472f39},
  {32'hc48a2dd4, 32'h43672d11, 32'hc30603f2},
  {32'h44a86e74, 32'hc32a5067, 32'h4314c280},
  {32'hc4db11b0, 32'hc326fcbc, 32'h4346ffe3},
  {32'hc2c80990, 32'h43986251, 32'h4325f01e},
  {32'hc4b1715c, 32'hc03b2234, 32'hc33acf4a},
  {32'h44e54c66, 32'hc32db400, 32'h431e653c},
  {32'hc510a6b0, 32'hc320c559, 32'h429d921c},
  {32'h44f0f788, 32'hc31d3463, 32'hc2a90d7a},
  {32'hc50bb873, 32'h41e285e6, 32'h440aeef5},
  {32'h4488bc2f, 32'hc0f994ba, 32'hc2e46f04},
  {32'hc40f485f, 32'hc2e940e1, 32'h42439daa},
  {32'h44ce69e4, 32'h40e9d798, 32'h43817d4e},
  {32'hc4d053b2, 32'hc3224f53, 32'h42e23a16},
  {32'h44c99720, 32'hc3674826, 32'h43d0d2ad},
  {32'hc508def0, 32'hc2635036, 32'hc394ae36},
  {32'h44ec62fb, 32'h4319cace, 32'hc3573f60},
  {32'hc50ecbc1, 32'h4143af05, 32'hc317a005},
  {32'h447106b3, 32'h43db30b9, 32'h431530bc},
  {32'hc505ad77, 32'h433d6f7f, 32'hc323177e},
  {32'hc3082340, 32'h42866dfb, 32'hc124af80},
  {32'hc50647fb, 32'h41a7457e, 32'h42f18cf9},
  {32'h445b9d40, 32'hc3a80a59, 32'hc3914a5f},
  {32'hc40d78e7, 32'hc1da5fe8, 32'hc34e64ca},
  {32'h450f2aec, 32'h430055c0, 32'hc3f6bda2},
  {32'hc4eca09a, 32'h42ad97f5, 32'hc32d03e5},
  {32'h43634280, 32'h428377e7, 32'hc394750d},
  {32'hc4cfa353, 32'h4251220a, 32'hc2daf520},
  {32'h4512d27d, 32'h42a77e41, 32'h41f21f32},
  {32'hc445f507, 32'hc1d16a91, 32'hc2a1215f},
  {32'h43c9c892, 32'h43307840, 32'h41cad52c},
  {32'hc4f15e8e, 32'h418aff17, 32'h431a190c},
  {32'h43b00992, 32'hc34f22d4, 32'h42b14036},
  {32'hc40b0644, 32'h4304fc46, 32'h42f4fb8e},
  {32'h44fb1acc, 32'h43e48b6e, 32'h43a9e259},
  {32'hc4650887, 32'hc354cee4, 32'h432a4d76},
  {32'h44848e18, 32'h4305e949, 32'hc249494f},
  {32'hc3e1ea98, 32'hc29344d5, 32'h43909d64},
  {32'h44a761e4, 32'h43ae4c0e, 32'hc31d4909},
  {32'hc4f9ca63, 32'h42ee84c3, 32'hc1e359fb},
  {32'h447453ec, 32'hc255527c, 32'hc14214a6},
  {32'hc4e69891, 32'hc2642ec7, 32'hc3c282a7},
  {32'h44e3085a, 32'hc177e4d0, 32'hc29a7737},
  {32'hc428def1, 32'hc2ad4cbc, 32'h4201741c},
  {32'h44bbfa62, 32'hc1c651d3, 32'hc2543ba8},
  {32'hc4c039b6, 32'h419bdde3, 32'h4260a88f},
  {32'h447f77ad, 32'hc3cf32fa, 32'h42fee064},
  {32'hc42d1ada, 32'hc2072f4a, 32'h43c8dba5},
  {32'h4428c8db, 32'hc2e30323, 32'hc35bcafe},
  {32'hc4f3babe, 32'h42d69a97, 32'h42889567},
  {32'h44b8c12a, 32'h43419421, 32'h428c0059},
  {32'hc402324e, 32'hc19c27e1, 32'h423c9a77},
  {32'h4505ea96, 32'hc2283998, 32'hc20f3f8f},
  {32'hc2aed5ac, 32'h4331c842, 32'h4345272f},
  {32'h44308d44, 32'hc347f202, 32'h429b79cc},
  {32'hc471f598, 32'h435dbb18, 32'h431029ec},
  {32'h4484afd7, 32'hc17c8c12, 32'hc084c7ac},
  {32'hc4c619c1, 32'hc30591e4, 32'h43ae08eb},
  {32'h44ff3c9d, 32'hc2ca40ed, 32'h43745245},
  {32'hc3998ac8, 32'hc2a8dc58, 32'h43cd1b2c},
  {32'h44da6432, 32'hc317c9d8, 32'h42e762ff},
  {32'hc4bbd8a8, 32'hc31196b3, 32'h43267345},
  {32'h445f8715, 32'h425038ff, 32'hc34007ad},
  {32'hc4cc32a6, 32'hc3719388, 32'h40fe76da},
  {32'h44ce56b1, 32'hc2f9e112, 32'hc289be4d},
  {32'hc464dcea, 32'hc199ef6c, 32'h439f5eef},
  {32'h44caae5d, 32'hc2f8e32b, 32'hc3e812dc},
  {32'hc4dd5ce5, 32'h4331fb77, 32'h435983f6},
  {32'h441f70b0, 32'hc39c5d85, 32'hc30a014a},
  {32'hc4835e18, 32'hc33eaf50, 32'hc234ec11},
  {32'h44e4a3d7, 32'h432ccf05, 32'hc32d92c4},
  {32'hc4bf8f30, 32'hc102cc1c, 32'hc366a59c},
  {32'h44bf9c36, 32'h43313647, 32'hc3592591},
  {32'hc4c026fe, 32'h441273bb, 32'h42f36531},
  {32'h44a21f9d, 32'h428033da, 32'h4231c1ac},
  {32'hc4d6af41, 32'hc1cf50fb, 32'h4356696a},
  {32'h44c5a49c, 32'h4306e895, 32'h43b9463b},
  {32'hc48beb80, 32'hc3250248, 32'h43245c49},
  {32'h43f33bb8, 32'hc3671309, 32'h43a1ff3a},
  {32'hc3286a1a, 32'hc33252ab, 32'h435555af},
  {32'h443e00e0, 32'h424332cd, 32'hc34eb4ab},
  {32'hc4998253, 32'hc42f1c49, 32'h439054e3},
  {32'h44ce6eaa, 32'h439ce97a, 32'h43955bb3},
  {32'hc4ef1e27, 32'hc38c1384, 32'h41ec2c80},
  {32'h4492d560, 32'h4357040e, 32'h43248ce7},
  {32'hc4fbc9ea, 32'h41db8749, 32'h42c0a740},
  {32'h44337054, 32'h43423141, 32'hc254a14e},
  {32'hc3b75a24, 32'hc34ddf5f, 32'h43677724},
  {32'h44d7e52c, 32'h4311cb9f, 32'hc32a37d6},
  {32'hc523ea96, 32'hc387ecc2, 32'h42968fbf},
  {32'h4480afdd, 32'h42669a5d, 32'hc3bab863},
  {32'hc4c0c5e5, 32'hc1ac91ce, 32'h40aab160},
  {32'h44579aa4, 32'hc2859844, 32'h428ea48a},
  {32'hc4e98e81, 32'hc2e610be, 32'h42c3949f},
  {32'h446030e2, 32'hc3e962bc, 32'hc382afc1},
  {32'hbdcc4000, 32'hc322629d, 32'hc2d17b9c},
  {32'h44ee0a9c, 32'hc3c4aaab, 32'h422b3642},
  {32'hc45697d1, 32'hc2b1b994, 32'h43404c93},
  {32'h449f56d5, 32'h43564a5e, 32'hc2217356},
  {32'hc4f3ca60, 32'hc311c12c, 32'hc13ca661},
  {32'h44f1f58c, 32'h41eeba65, 32'hc0d98490},
  {32'hc4b37ba3, 32'h43a22547, 32'hc2c07b1d},
  {32'h44fec625, 32'hc3689bb6, 32'h4297ee1c},
  {32'hc481fb2b, 32'h437ed071, 32'hc3c7eba3},
  {32'h446d071f, 32'hc3a829e7, 32'h43906e8c},
  {32'hc4b022dd, 32'hc29f4c71, 32'hc287e60e},
  {32'h44aafe0d, 32'hc4052244, 32'h4361067a},
  {32'hc2a12e31, 32'hc3edafc9, 32'h43399ea7},
  {32'h451c1acf, 32'hc26a4de7, 32'h43a1bb64},
  {32'hc51286c6, 32'hc120585c, 32'hc3a17ac5},
  {32'h4501cc3d, 32'hc388e78b, 32'h43e3aafb},
  {32'hc505138f, 32'hc3047507, 32'h43b7836b},
  {32'h4510ead7, 32'h417bad42, 32'hc36a5f73},
  {32'hc204bcc0, 32'h43081aeb, 32'hc12533b3},
  {32'h4510078e, 32'hc36127b0, 32'h431617da},
  {32'hc406c5b9, 32'h430cc454, 32'h421764e5},
  {32'h442dbe6e, 32'hc34f95d4, 32'h42c2e798},
  {32'hc45a004a, 32'hc39b1a4f, 32'hc2e12982},
  {32'h3fc92400, 32'hc2d54d2b, 32'h4312e3d5},
  {32'hc4c90dba, 32'hc3d201db, 32'h426fda1b},
  {32'h44b77e53, 32'h436e5bda, 32'hc3130373},
  {32'hc3bcb2f8, 32'h42ce18ad, 32'hc35e79e3},
  {32'h43ff5085, 32'hc2a885a0, 32'h43da462a},
  {32'hc5161cf1, 32'hc2b1d134, 32'h43a64305},
  {32'h44a243b8, 32'h42f744ba, 32'h432358aa},
  {32'hc494c37e, 32'hc39c33c0, 32'hc2ad3063},
  {32'h4468a8fc, 32'hc2dcd665, 32'hc24da199},
  {32'hc49a17b0, 32'hc34cb9c9, 32'h42fa1d10},
  {32'h44eb931f, 32'hc31c5616, 32'h435f60d4},
  {32'hc4a58d0b, 32'h43a267db, 32'h433daa9d},
  {32'h442b6648, 32'hc28b447d, 32'hc359f768},
  {32'hc486bd1d, 32'h43249d2b, 32'h4312d5bd},
  {32'h4407b9ee, 32'h4282bdb2, 32'hc30cf2b9},
  {32'hc4e1178c, 32'h432f01b3, 32'hc3c55a1e},
  {32'h4405a3e2, 32'hc368e1ce, 32'h4212c1bb},
  {32'hc43b772a, 32'h433024f6, 32'h433594f7},
  {32'h44d090d4, 32'h42c9e75e, 32'hc2b47ab1},
  {32'hc5052ab0, 32'hc24a8223, 32'hc30a37e1},
  {32'h44028e6c, 32'hc38c8143, 32'hc3651f34},
  {32'hc4a75fc7, 32'h4240e284, 32'hc33e8f55},
  {32'h438a3250, 32'h42ada6b9, 32'h421e9110},
  {32'hc44a37a2, 32'hc1de2201, 32'h4324083c},
  {32'h44d7f7f5, 32'h4330ccb7, 32'hc332af46},
  {32'hc480ae30, 32'h3fda2129, 32'h4396504d},
  {32'h4506f15f, 32'h44117d9a, 32'h43ae059e},
  {32'hc50d2481, 32'h4309c0e2, 32'h439cf296},
  {32'h450c4eb8, 32'hc2903554, 32'hc31ca535},
  {32'hc50ada4e, 32'hc2fb56bd, 32'hc34f6617},
  {32'h44c49442, 32'hc2128cd2, 32'h4264ebd9},
  {32'h4030ec90, 32'h41b18a82, 32'hc3296b18},
  {32'h446381c0, 32'h43b64570, 32'h42d4e162},
  {32'hc49c4e3a, 32'h42c216ce, 32'hc2315722},
  {32'h44c0f4fe, 32'hc297f7e5, 32'hc32e9483},
  {32'hc44a092c, 32'hc261e6fc, 32'hc3880716},
  {32'h441e3f2b, 32'hc2acf929, 32'hc303ac15},
  {32'hc51b8be9, 32'hc3d12951, 32'h43c14fb9},
  {32'h43323f58, 32'h434e04d6, 32'hc25e189a},
  {32'hc477faf8, 32'h42d5fd0f, 32'hc39d7e1f},
  {32'h44263144, 32'hc37a6ab1, 32'h42de9b49},
  {32'hc4ad49d4, 32'hc361d726, 32'h41e37683},
  {32'h44ff766b, 32'hc1b5fcc8, 32'hc3acf799},
  {32'hc51ad2f2, 32'h438748b0, 32'h42773c9a},
  {32'h44c862a3, 32'h43449605, 32'h43acdc7f},
  {32'hc50c592e, 32'hc104a4b7, 32'h42b9fe47},
  {32'h45229047, 32'hc2a8765d, 32'hc3fcab30},
  {32'hc4c4dab1, 32'h3e7af5ae, 32'h43ab8ad7},
  {32'h451130f4, 32'hc2093419, 32'hc399012b},
  {32'hc4746ebc, 32'hc4170e3a, 32'hc2dffe14},
  {32'h4498f2f7, 32'h42d591ef, 32'h428a99db},
  {32'hc32f7ff0, 32'hc32f93f6, 32'h435dd6a7},
  {32'h451864d5, 32'hc3533d00, 32'hc3778550},
  {32'hc5031708, 32'hc3211a9e, 32'h414060b0},
  {32'h4482fff7, 32'hc3120e94, 32'h42b07ab8},
  {32'hc4ccc6a9, 32'h42e03525, 32'h42b00c20},
  {32'h44a319a8, 32'h43250cde, 32'hc317a410},
  {32'hc3ded53b, 32'hc2a365ee, 32'hc3c2dc41},
  {32'h450e0e5e, 32'hc296f714, 32'h429e3683},
  {32'hc3ad57fc, 32'hc363ea4a, 32'h43b5deea},
  {32'h444d5cdc, 32'hc33564fd, 32'hc333ae06},
  {32'hc49d0df5, 32'hc36a2e82, 32'hc2edb956},
  {32'h43d2d2c2, 32'h4253531e, 32'h437b1778},
  {32'hc3eda6e8, 32'hc214bf64, 32'hc3b9577b},
  {32'h44b202f6, 32'hc1be50a6, 32'h43c6dc57},
  {32'hc45124ca, 32'hc3b90da1, 32'h4192f399},
  {32'h450a6e1c, 32'hc28123ae, 32'hc26c0152},
  {32'hc4d199b6, 32'hc34be440, 32'h436c1e25},
  {32'h44012371, 32'hc2bf193d, 32'h4309f2e4},
  {32'hc48670ed, 32'h4291a74c, 32'h430a4aed},
  {32'h44e44dd5, 32'hc39034c1, 32'h432e0789},
  {32'hc504be74, 32'hc38fcab7, 32'hc33e1baa},
  {32'h43a56ec4, 32'h42968675, 32'hc2c0433b},
  {32'hc5150aca, 32'hc33eaf37, 32'hc2ff16c8},
  {32'h4518a17d, 32'hc38b9d87, 32'hc39727a2},
  {32'hc4bfb29f, 32'h409ed37e, 32'h42fdad1a},
  {32'h443540d4, 32'hc3b0e696, 32'h43f4f869},
  {32'hc3f0a952, 32'hc33070e3, 32'hc1dc56d0},
  {32'h4325d0b0, 32'h419007c9, 32'hc2cd25af},
  {32'hc5163948, 32'hc2f77dc5, 32'hc2b053c7},
  {32'h4505f054, 32'h42ece700, 32'h435309d5},
  {32'hc49702a2, 32'h43a0d284, 32'h438d8de9},
  {32'h4428475a, 32'h42914f46, 32'hc2292d88},
  {32'hc5010c8d, 32'h43abef80, 32'hc12de9ae},
  {32'h44c70dd9, 32'h435e3af8, 32'h436a690a},
  {32'h41ed7900, 32'h41e4e9c4, 32'hc3b5a885},
  {32'h44f857ef, 32'hc2c51103, 32'h42a2a353},
  {32'hc455e84f, 32'hc3b30c79, 32'h4252dc8e},
  {32'h4426a384, 32'hc36ef085, 32'h41f0bd82},
  {32'h40c1ce00, 32'h4354e6ee, 32'hc2bafb5a},
  {32'h44c5b7a1, 32'hc1ca4e1a, 32'hc2e67e35},
  {32'hc3f8e840, 32'hc3a28950, 32'h432de85c},
  {32'h440422cc, 32'hc1a05c58, 32'hc2b246eb},
  {32'hc31ac1fe, 32'h42469594, 32'hc2dcf9ad},
  {32'h449ccea4, 32'h42c95302, 32'hc2c1a8de},
  {32'hc495d796, 32'h418c74b2, 32'hc3a4b3e2},
  {32'h449f6f82, 32'hc3c3496a, 32'h4386c823},
  {32'hc4bd6e85, 32'hc38af1b2, 32'hc3f8be24},
  {32'h447f0834, 32'h4375cad5, 32'hc2fdd729},
  {32'hc4c0bee7, 32'hc3567976, 32'hc235efc4},
  {32'h44a776b2, 32'h4092df52, 32'h4339c3cc},
  {32'hc494a7e3, 32'hc3bbb6d4, 32'hc372be6a},
  {32'h4489d610, 32'hc301bae7, 32'hc346970a},
  {32'hc4ae5c60, 32'hc29cfc4b, 32'hc3827de6},
  {32'h442a0e1e, 32'h42131204, 32'hc1d342fc},
  {32'hc509ba65, 32'h435ef2dc, 32'h42f5d5c6},
  {32'h449574bb, 32'h4245182c, 32'h43800196},
  {32'h4381d9b0, 32'h43042298, 32'h4402c678},
  {32'h44f48160, 32'hc3832f30, 32'h422fdca1},
  {32'hc4d6c8e0, 32'hc319502b, 32'hc313d4df},
  {32'h44e1f5b7, 32'h4289f4e9, 32'hc29aaff8},
  {32'hc504f01f, 32'h42b2d812, 32'h439ae0ca},
  {32'h449cb183, 32'h43987089, 32'hc37c2f13},
  {32'hc4bcb75c, 32'h4326a7d7, 32'hc4159766},
  {32'h44a31132, 32'hc2fbedcd, 32'h44076b47},
  {32'hc4fb92cc, 32'hc36308f5, 32'h4395b52e},
  {32'h4502f886, 32'hc319595d, 32'h43a48be9},
  {32'hc4975d33, 32'h4305d24c, 32'hc4054463},
  {32'h4497b07c, 32'hc2806172, 32'h42d4a492},
  {32'hc3663c65, 32'h429bca8b, 32'hc2cd6fe5},
  {32'h43c5ad5a, 32'hc31b53c5, 32'h430720b2},
  {32'hc38c8180, 32'h40c2362e, 32'hc3a45840},
  {32'h4322e3b8, 32'h429b7c2d, 32'h42bf7962},
  {32'h40a5f800, 32'hc349905e, 32'h40e2c2fb},
  {32'h44eb60b2, 32'h4385010a, 32'hc30f56cb},
  {32'h40b35800, 32'hc36f7394, 32'hc34d07f2},
  {32'h447e5aa2, 32'hc271203a, 32'h431822d6},
  {32'hc4111e0c, 32'hc29ff6ba, 32'h4351cdea},
  {32'hc45efbee, 32'h422757a8, 32'h429248eb},
  {32'h451075ba, 32'hc3320d81, 32'h43864afc},
  {32'hc4ffe236, 32'hc328324b, 32'hc3840fc8},
  {32'h449fc324, 32'hc28b43fd, 32'hc39613cf},
  {32'hc4c76663, 32'h422f5028, 32'hc37b6d01},
  {32'h449fcd2a, 32'hc3d1a8b2, 32'h438b2fb9},
  {32'hc43f1850, 32'hc3958d69, 32'h430b467c},
  {32'h4492de72, 32'h43335d0d, 32'h438ec6a4},
  {32'hc511948b, 32'hc0d8d8e0, 32'hc3ae9754},
  {32'h448f0432, 32'h41a4445e, 32'hc356021c},
  {32'hc4bd5c0f, 32'h437f5348, 32'hc1ef7077},
  {32'h450f635b, 32'h4281a77f, 32'h43f85cb6},
  {32'hc3c4ceeb, 32'h438e2092, 32'hc3e2b3c2},
  {32'h44878194, 32'hc2bd6f42, 32'h43be66f3},
  {32'hc4b7de4c, 32'hc323e439, 32'hc2c192fd},
  {32'h44170e0e, 32'h43098d07, 32'hc2922170},
  {32'hc5015eeb, 32'h43928cba, 32'hc36d7269},
  {32'h44806331, 32'h4355d2cc, 32'h4389ea72},
  {32'hc4c7debb, 32'hc2a4ceef, 32'hc2815071},
  {32'h44a8c4d6, 32'hc3c3c3e2, 32'h431438de},
  {32'hc4f07fe8, 32'h42a0f22c, 32'hc379d447},
  {32'h44889a1b, 32'hc3303924, 32'hc38a208b},
  {32'hc429de1b, 32'h42a92845, 32'hc38eb560},
  {32'h448c1b94, 32'hc3c1ba63, 32'h439aedd2},
  {32'hc502eccf, 32'hc3044d46, 32'hc347e3a3},
  {32'h4510f9da, 32'hc394b7a8, 32'h435fa870},
  {32'hc4e75db5, 32'h4394f7b8, 32'h430764f0},
  {32'h443e6270, 32'h4322c4e1, 32'h435ccee7},
  {32'hc4a2a4be, 32'h432500c6, 32'hc3a05f11},
  {32'h44b87db4, 32'hc3e5abd3, 32'hc28c3cfb},
  {32'hc50965ff, 32'h40a23fe8, 32'hc29dcf17},
  {32'h44a58ec2, 32'hc3baeb12, 32'hc3755447},
  {32'hc4cf466b, 32'h420c9988, 32'hc3f5c69b},
  {32'h44ac2132, 32'h434f2611, 32'h431908c7},
  {32'hc4d5caf9, 32'hc22ef38b, 32'hc303b593},
  {32'h44b0a2a5, 32'hc35bef77, 32'h43683a68},
  {32'hc42067e8, 32'hc3aaf4a3, 32'h438ddfeb},
  {32'h44985168, 32'h4184b7e8, 32'hc341905a},
  {32'hc2200b60, 32'hc3a7e65c, 32'hc2ad33f0},
  {32'h42b8131d, 32'h4318c034, 32'hc352f35d},
  {32'hc50ceb12, 32'hc236d8e5, 32'hc2de5e82},
  {32'h43847bdf, 32'h4122958b, 32'hc3903701},
  {32'hc45c67f8, 32'hc3982d8a, 32'h42228a1c},
  {32'h451e9f93, 32'h438218ec, 32'h4268a789},
  {32'hc424dc6f, 32'hc3af942e, 32'h413930f8},
  {32'hc238fd00, 32'h43902a27, 32'h4345b888},
  {32'hc4265690, 32'h423ba3c2, 32'hc31bfeae},
  {32'h43ed4d48, 32'h438f9c04, 32'h4325df36},
  {32'hc49b315e, 32'h40c379a7, 32'hc292afaa},
  {32'h43dea432, 32'h435a4bd0, 32'h422839ac},
  {32'hc4101c7e, 32'h43ee1f49, 32'h43175c6a},
  {32'h44ebd8ed, 32'h424264d6, 32'hc30dd1ca},
  {32'hc44bd5ee, 32'hc3cdab72, 32'hc32e9693},
  {32'h4514585a, 32'hc395f16b, 32'h4315fac7},
  {32'hc50918c6, 32'h42a84bc1, 32'hc330a8c7},
  {32'h43fb3c9c, 32'h4315445a, 32'hc141d99d},
  {32'hc4f9f50e, 32'h431db953, 32'hc3861055},
  {32'h450146d0, 32'hc2ff19e7, 32'hc1407fe9},
  {32'hc3be4920, 32'h43be16a9, 32'h41595f30},
  {32'h45004bcc, 32'h4332e580, 32'h44007876},
  {32'hc4d3ecdb, 32'hc1a3c4e5, 32'hc3365311},
  {32'h44a76d2c, 32'hc3249c8c, 32'hc2bf820e},
  {32'hc4a77be9, 32'h42c53a1b, 32'hc39312db},
  {32'h44e40a7a, 32'hc2b7a445, 32'h42c6da7e},
  {32'hc4f054ef, 32'hc3a415de, 32'hc372c6b6},
  {32'h434da7d0, 32'hc3294b99, 32'h437acf9b},
  {32'hc2efa740, 32'h43b0ce33, 32'hc33f7fb9},
  {32'h450d1ae4, 32'h423f9210, 32'hc401768c},
  {32'hc4719223, 32'hc3351202, 32'hc37fef66},
  {32'h44d0013d, 32'h42e8658c, 32'h437f9c64},
  {32'h43460d28, 32'hc1b8325a, 32'hc3185cfb},
  {32'h433d0f70, 32'h4264761e, 32'h4390a224},
  {32'hc32862e0, 32'h4352ea74, 32'h4306a2f4},
  {32'h42e993f8, 32'hc1a00c48, 32'hc26140ee},
  {32'hc4b79c6f, 32'hc21664e9, 32'hc2855d8f},
  {32'h4464d9e0, 32'h4290ce87, 32'hc291660f},
  {32'hc3a34783, 32'h42d20dc5, 32'hc33870bf},
  {32'h4501432b, 32'h429c8639, 32'hc229ea0d},
  {32'h42259bb1, 32'hc3b1a9eb, 32'h433d7d95},
  {32'h45310224, 32'hc2ad2c90, 32'h42eb6eea},
  {32'hc47b54cf, 32'h4222e6ec, 32'hc369b3bd},
  {32'h451b186d, 32'hc37c49b3, 32'h4299c497},
  {32'hc4cafc50, 32'hc33f0c8c, 32'hc303fe6f},
  {32'h45075fed, 32'h42dea51d, 32'hc2fc2e28},
  {32'hc24eb700, 32'h438921ba, 32'h42677e08},
  {32'h44aeac29, 32'h42cfcab6, 32'h436ffdc7},
  {32'h42808ad0, 32'hc3805565, 32'h43ede964},
  {32'h4520a4a8, 32'hc2775632, 32'hc2d1cf9d},
  {32'hc20adee0, 32'hc3bcd2b4, 32'h433c9670},
  {32'h44e1cee7, 32'h426c77cc, 32'hc3677c8a},
  {32'hc4a41cf8, 32'hc2a386e4, 32'hc3217b7e},
  {32'h43e64b35, 32'hc153ed45, 32'h430183e4},
  {32'hc504f63a, 32'hc19f5153, 32'hc4189546},
  {32'h449eb446, 32'hc03a9c16, 32'h43738020},
  {32'hc39c25c4, 32'h42d0dec3, 32'h41cc2aff},
  {32'h451f27ab, 32'hc35d011d, 32'hc289e3fc},
  {32'hc3553420, 32'hc2904955, 32'hc3837c1a},
  {32'h43fd9418, 32'hc3b765bc, 32'hc3d1d92c},
  {32'hc494af5c, 32'hc40431c0, 32'h42aa3e8d},
  {32'h44b0d7eb, 32'h4352f917, 32'h43dfc98b},
  {32'hc42828b0, 32'h43a6a009, 32'h43764474},
  {32'h43e47e1c, 32'h439ce6eb, 32'hc333f5ce},
  {32'hc4f1ae24, 32'hc33acd4b, 32'hc28ee96d},
  {32'h435d6f80, 32'hc39b7d5a, 32'h43e86ab6},
  {32'hc4c7e4de, 32'h4297cbae, 32'h436f70d7},
  {32'h4512e4a1, 32'h427bf803, 32'hc39a4a2c},
  {32'h43c2179f, 32'hc2c503f1, 32'h428a4432},
  {32'h451e8774, 32'h42f66a91, 32'hc21ac920},
  {32'hc3ae5eec, 32'h418873d3, 32'hc1a529f2},
  {32'h44c716a0, 32'h43795fbe, 32'h43cd1258},
  {32'h43b5bd70, 32'hc350157f, 32'h431f3dce},
  {32'h44bc1146, 32'h435550bd, 32'hc2d6cc11},
  {32'hc4befa4e, 32'hc0b42e92, 32'h43942aee},
  {32'h44f23cb6, 32'h441329e6, 32'hc28f8c92},
  {32'hc4d37387, 32'hc3990f23, 32'h439900f0},
  {32'hc3039d98, 32'hc2db2aba, 32'hc35e05f9},
  {32'hc458cda6, 32'h43cb0aae, 32'hc348bfc6},
  {32'h447aeae0, 32'hc101897d, 32'hc3a703ec},
  {32'hc4fba9c4, 32'hc2b6433e, 32'h4326e780},
  {32'h44db9696, 32'hc3e1fff2, 32'hc38d32bb},
  {32'hc40e4dff, 32'hc3214d6d, 32'hc237eb25},
  {32'h44683910, 32'hc3669813, 32'h430f6c10},
  {32'hc4d0e311, 32'h425ae77e, 32'h42204281},
  {32'h43817266, 32'h4336bd5c, 32'hc328c219},
  {32'hc4f54ef3, 32'hc31562f6, 32'hc1be4b08},
  {32'h450e617c, 32'h40071760, 32'hc33d90ae},
  {32'hc4a3d313, 32'hc3a8c192, 32'hc33213ea},
  {32'h44073a6a, 32'h4301f968, 32'h4380f1d2},
  {32'hc50452e1, 32'hc21864a2, 32'h43134706},
  {32'h44cb83a0, 32'h42327836, 32'hc06c47a6},
  {32'h42c5e8c0, 32'h437cb818, 32'hc3b8a7a6},
  {32'h4508b52a, 32'hc28e8c7c, 32'h43606384},
  {32'hc4ddac4c, 32'hc333a190, 32'h42c95d32},
  {32'h441174f4, 32'hc292573a, 32'h42f3b4f6},
  {32'hc4e8716f, 32'hc2b57489, 32'hc40214f0},
  {32'h448128fc, 32'hc2abbdbc, 32'hc41d6f7b},
  {32'hc4f0df1c, 32'h41fc9cb0, 32'hc349cdd7},
  {32'h4400eecb, 32'h43095b02, 32'hc3fdbf15},
  {32'hc489fec3, 32'hc32efdf2, 32'h43b07105},
  {32'h44a6d890, 32'h41a6d9ac, 32'hc351669e},
  {32'hc48efa6b, 32'hc3d55ac1, 32'h42c88fda},
  {32'h40023c00, 32'hc390a9cd, 32'h431d3008},
  {32'hc42e5738, 32'hc376c336, 32'h43d62d96},
  {32'h446b2cd4, 32'hc3c27fa4, 32'hc3937312},
  {32'hc4eadc6a, 32'h42a6a17f, 32'h42f2899a},
  {32'h43bdbb0c, 32'h42adb740, 32'hc23a7a28},
  {32'hc4142fe2, 32'hc1b8dcd6, 32'h4387f75c},
  {32'h4498018d, 32'h42b4a7d6, 32'hc235ea78},
  {32'hc499a154, 32'h42ebd3a0, 32'h43886644},
  {32'h45001cfa, 32'h42644274, 32'hc35b1259},
  {32'hc4859a54, 32'h43d3f8ba, 32'hc191e91e},
  {32'h4495a843, 32'h43a0e543, 32'h434433ab},
  {32'hc3de7beb, 32'hc38dc336, 32'hc2fe5146},
  {32'h44e21cae, 32'hc3a21710, 32'hc28d05d1},
  {32'hc4e9f06a, 32'h43a56a64, 32'h42a7dc70},
  {32'h44d4f361, 32'h42c0e45c, 32'hc204243c},
  {32'hc47ae7d8, 32'hc1c1658c, 32'h42eac435},
  {32'hc27d13d8, 32'hc324a8ae, 32'hc301454f},
  {32'hc377ac78, 32'h43ab33e5, 32'hc225d0d1},
  {32'h43c61c5c, 32'h4314e182, 32'h43877dee},
  {32'hc4f265a8, 32'hc3387d6b, 32'h42c7ace2},
  {32'h44dca2a9, 32'hc38e3109, 32'hc3f5c059},
  {32'hc3804894, 32'h42f96d16, 32'hc1575ca7},
  {32'h41782800, 32'hc400afc2, 32'hc34d0614},
  {32'hc47b1b72, 32'h437bd52a, 32'h43607605},
  {32'h449ee194, 32'h434dab5c, 32'h41e15a67},
  {32'hc4d27b78, 32'h42c69709, 32'h43a9f8fc},
  {32'h444d88f2, 32'hc396231d, 32'h4223f293},
  {32'hc512e406, 32'hc334f8b6, 32'hc2434dd8},
  {32'h44b98f49, 32'hc3b80428, 32'hc2da408b},
  {32'hc4d65f3a, 32'h414089ef, 32'hc2854795},
  {32'h44cc840d, 32'h42dca142, 32'hc36869f7},
  {32'hc46f8e60, 32'h41b45ecc, 32'hc35f3d87},
  {32'h4404e2ec, 32'h43208be0, 32'h41574cef},
  {32'hc4dba40c, 32'hc349659b, 32'hc3dce6bc},
  {32'h445bddf0, 32'h431f0ce4, 32'h439b2f0e},
  {32'hc4a2dcae, 32'h43803759, 32'h43494d8a},
  {32'h44e4e028, 32'hc25d0459, 32'hc3019a61},
  {32'h40fbd000, 32'h43a397b8, 32'hc46899d1},
  {32'h44b99778, 32'hc2f12841, 32'hc3ecad6b},
  {32'hc3c238eb, 32'hc283d936, 32'hc3c0a0f3},
  {32'h44489e17, 32'h43b5e9c6, 32'hc3911566},
  {32'h438f4280, 32'hc2f69a71, 32'h43965eb8},
  {32'h447ab423, 32'hc2908e0d, 32'h41d145d9},
  {32'hc4c49f18, 32'hc1a2284e, 32'h420d38ba},
  {32'h4496fbde, 32'h43898938, 32'h437640ef},
  {32'hc404807b, 32'h4272eb55, 32'h41a415a6},
  {32'h4502d66c, 32'hc3caea8e, 32'hc313d690},
  {32'hc4946192, 32'hc3ad4f10, 32'hc349d878},
  {32'h43ace4fc, 32'hc36684a0, 32'hc3898ddd},
  {32'hc4049095, 32'hc3885dfe, 32'h438094c6},
  {32'h448caca8, 32'hc30dc271, 32'hc36494a1},
  {32'hbebaa800, 32'h438e5b3c, 32'h4318de68},
  {32'h44455510, 32'h41e25fc4, 32'h43d03253},
  {32'hc4a5f27e, 32'hc346b3ca, 32'hc384a553},
  {32'h44e716ee, 32'h43697fc6, 32'h441c09ca},
  {32'hc500a3d1, 32'hc20267e9, 32'h42cdf89e},
  {32'h451ae8a6, 32'hc30ba12d, 32'h435db69a},
  {32'hc4c09162, 32'h41de352b, 32'h420fe46d},
  {32'h44b7f11e, 32'hc3422449, 32'h42eef590},
  {32'hc471e982, 32'hc1b968c2, 32'hc35147b1},
  {32'h4499daf7, 32'hc3110a35, 32'h42ff2bf9},
  {32'hc47777be, 32'h3eab1ec0, 32'h4362c5b4},
  {32'h44a1ab8d, 32'h431cd747, 32'hc1a67f2b},
  {32'hc4854000, 32'hc3726337, 32'hc22f5967},
  {32'h4409ab24, 32'hc2c2840e, 32'hc3927bd0},
  {32'hc4b49f8c, 32'hc3452595, 32'h4205d372},
  {32'h446cf01f, 32'h4383d4f5, 32'hc2dafd1e},
  {32'hc5137cb9, 32'hc187f3be, 32'hc3127666},
  {32'h450ddcfb, 32'hc2939334, 32'hc3c16233},
  {32'hc4a1a353, 32'hc3942679, 32'h42f77d73},
  {32'h44c5e5b5, 32'h428f1e15, 32'h43271343},
  {32'hc40d27e0, 32'h43878599, 32'hc372fa5f},
  {32'h43d433e8, 32'hc345f898, 32'hc299add7},
  {32'hc343a2b0, 32'h413c2932, 32'hc3ec3867},
  {32'h4436e141, 32'h430600e2, 32'h430f14ae},
  {32'hc4cfef34, 32'hc3c0b0a2, 32'hc359bc76},
  {32'h428afce8, 32'h43933028, 32'h43f20fb4},
  {32'hc379e140, 32'hc20f2d92, 32'hc242686c},
  {32'h3f0acc00, 32'hc2f3906b, 32'h42660e70},
  {32'hc49b95b7, 32'hc2dcea19, 32'h426d2353},
  {32'h443de687, 32'h4284d574, 32'hc29d0a3c},
  {32'hc466700c, 32'h43020e34, 32'h432b4422},
  {32'h44a8de27, 32'h430ee954, 32'h43823daa},
  {32'hc0ef8c00, 32'h420ea041, 32'hc2ee20d5},
  {32'h42dde130, 32'hc308b2eb, 32'hc38466b0},
  {32'hc447b83b, 32'h4214e85c, 32'h43c7dc94},
  {32'h442ba307, 32'hc3ad2843, 32'hc428c185},
  {32'hc50ef7e0, 32'h40143612, 32'h42aa85aa},
  {32'h44d6d52e, 32'h430232be, 32'h42556d65},
  {32'hc4819f02, 32'hc26f6225, 32'h430df336},
  {32'h44f6102c, 32'hc31432c2, 32'hc393f404},
  {32'hc4a38ef6, 32'hc32c3d90, 32'hc29b72d1},
  {32'h440da615, 32'hc2f480ef, 32'h42c809f8},
  {32'hc4184dab, 32'h430fa0ac, 32'hc08210a7},
  {32'h44dadd0a, 32'h430f8db0, 32'hc3549678},
  {32'hc4b8a8ca, 32'hc377f42d, 32'h42ca5a47},
  {32'h44b660c4, 32'h42ee1c75, 32'h439a5129},
  {32'hc46e7e66, 32'hc396ed8f, 32'hc2a55fce},
  {32'h450770a4, 32'hc30f3055, 32'hc2a4802a},
  {32'hc4e0fe94, 32'h43024661, 32'h43119093},
  {32'h439fd818, 32'hc2b9aa2f, 32'hc1c78cf8},
  {32'hc4451b20, 32'h41f863c0, 32'h41cdc6ac},
  {32'h44b24876, 32'hc2212d70, 32'h42200ccf},
  {32'hc3fd76ab, 32'hc1d62638, 32'h43300960},
  {32'h4456f01a, 32'h439ebe93, 32'h42943370},
  {32'hc4bfe5c7, 32'hc22c7796, 32'hc39b1374},
  {32'h45032163, 32'h42f661dd, 32'h4365d856},
  {32'hc4f55584, 32'hc2aa761e, 32'h433d3137},
  {32'h44e183d0, 32'h43a3168c, 32'h419dcd00},
  {32'hc4278df8, 32'hc340100f, 32'hc3626b46},
  {32'h44c90387, 32'hc33d73b7, 32'h436ce30f},
  {32'hc4965e9e, 32'hc38566c5, 32'h433abcaf},
  {32'h435638ec, 32'hc3ab1ed5, 32'h43219517},
  {32'hc4c0796e, 32'hc343830c, 32'h42938b22},
  {32'h44007f7c, 32'h428bfc3e, 32'hc30728ee},
  {32'hc4e7fe50, 32'hc2d01bca, 32'hc3abc5b0},
  {32'h44f3f622, 32'h43748ea5, 32'hc25408a9},
  {32'hc4b5c8b8, 32'h428d2778, 32'h4355edf5},
  {32'h450ba1ea, 32'h42969d47, 32'hc3196856},
  {32'hc3be154e, 32'hc2d9eb43, 32'hc3e17fcc},
  {32'h450294aa, 32'h42f102cd, 32'hc364fecb},
  {32'hc499e24d, 32'h43890232, 32'hc3c4feb4},
  {32'h44c9a6aa, 32'hc3873c3c, 32'h43cc43f5},
  {32'hc40e4df0, 32'hc2ac59e3, 32'hc37316ca},
  {32'h44e57644, 32'hc2e7da11, 32'hc38da53b},
  {32'hc4cbd7de, 32'h4214509c, 32'h418d0bba},
  {32'h44d3b976, 32'h433e6b3d, 32'h431c614a},
  {32'hc34a3c21, 32'h43cba400, 32'hc4146526},
  {32'h447d7d48, 32'h42a1f36c, 32'hc221d19b},
  {32'hc50655f6, 32'h42626add, 32'h430bc508},
  {32'h438cf112, 32'h434c6a06, 32'hc26172f8},
  {32'hc4f98d22, 32'hc3a64f4d, 32'hc2e593bd},
  {32'h448b02e9, 32'h42e2134f, 32'h415472fb},
  {32'hc5178438, 32'h42f8aab3, 32'hc3a5afda},
  {32'h450b9871, 32'h439c1d88, 32'hc382318d},
  {32'hc5209598, 32'hc2fe1e0a, 32'h43c08381},
  {32'h4434065d, 32'hc345c691, 32'h41f36237},
  {32'hc443afb4, 32'h4279586f, 32'hc3da957e},
  {32'h44f49510, 32'hc287d22c, 32'h43803f3b},
  {32'hbfc16d40, 32'h43d5bcad, 32'h431bac5a},
  {32'h438aac5c, 32'h43babb54, 32'hc3bc806e},
  {32'hc44a2bb8, 32'h42aa1e0a, 32'hc2c7c11d},
  {32'h4437ad56, 32'hc16be3f3, 32'h42d9b9a7},
  {32'hc42a270c, 32'h4328d4a8, 32'hc380b29a},
  {32'h44713043, 32'hc3a8e4ba, 32'hc314e92c},
  {32'hc4941031, 32'h41bf4463, 32'h43dec276},
  {32'h442260a0, 32'h43b2e6e2, 32'h43b5eaf7},
  {32'hc480479a, 32'h4281a1e2, 32'h4314e26c},
  {32'h449af542, 32'hc2fcbc10, 32'hc3f7888a},
  {32'hc4431ee6, 32'hc3ab585b, 32'hc19e4c8e},
  {32'h42054e80, 32'h412ce274, 32'hc3925197},
  {32'hc3d93dbc, 32'hc2204464, 32'h4243f81c},
  {32'h450eb3f6, 32'hc2dd1986, 32'h41bea2b2},
  {32'hc49566ff, 32'hc2e1fbfa, 32'h420b1e15},
  {32'h44506170, 32'hc21e7ac4, 32'hc31cd5ad},
  {32'hc4bd28a3, 32'h43c317bc, 32'h42bb709f},
  {32'h448b6030, 32'hc339d92e, 32'h438d4cbf},
  {32'hc3f43890, 32'hc3d2f7d5, 32'hc36d475f},
  {32'hc1ea72c0, 32'hc3bb7c9f, 32'h438d5a8a},
  {32'hc525eef3, 32'h434431f0, 32'hc3c8c1de},
  {32'h45273bfa, 32'hc351879a, 32'hc37dcc59},
  {32'hc502ff88, 32'h42544a77, 32'h43e64ed1},
  {32'h44542159, 32'hc21746d1, 32'hc283a2ab},
  {32'hc46dfe91, 32'hc21d7c26, 32'hc3ab4f86},
  {32'h4511b09d, 32'hc2515d5d, 32'hc3a0c65a},
  {32'hc3d4e94c, 32'h4312c58a, 32'h42590b0f},
  {32'h44d541de, 32'hc2f11335, 32'hc39aab44},
  {32'hc49dd898, 32'hc38f2a3b, 32'h4277a39a},
  {32'h44bd888d, 32'hc09a3088, 32'hc3270150},
  {32'hc41053f1, 32'h41eda0d2, 32'h4346751f},
  {32'h44212d2d, 32'h43316fee, 32'h41591a6f},
  {32'hc3aab848, 32'h43beed35, 32'h430cdd44},
  {32'h43f95618, 32'hc358b158, 32'hc306111e},
  {32'hc493a7e8, 32'hc2e378b6, 32'hc3808854},
  {32'h45152972, 32'h43ee829e, 32'h43890b0a},
  {32'hc4c1a05e, 32'h41c0cc48, 32'h4390ed27},
  {32'h41c0edd0, 32'hc3a46565, 32'h43962cea},
  {32'hc3e8a79b, 32'h408995a9, 32'h3f03df21},
  {32'h451700c7, 32'hc3828e47, 32'hc3a58682},
  {32'hc3d8139c, 32'h42d65837, 32'hc3312861},
  {32'h44316e19, 32'hc412d7d3, 32'hc37fb077},
  {32'hc2a175f0, 32'hc2aaceb4, 32'hc3415fee},
  {32'h4539317c, 32'hc1b5231e, 32'hc349d0b5},
  {32'h439778f0, 32'hc3a5766d, 32'h4316e681},
  {32'h44af3afa, 32'hc37d81cc, 32'h4381bd68},
  {32'hc49e6179, 32'hc2d3e3fa, 32'h43d152e6},
  {32'h43b2c278, 32'h4218b090, 32'h43627bd6},
  {32'hc4bd80a3, 32'h4319873b, 32'hc343ccfd},
  {32'h451e356c, 32'hc3b3e7cc, 32'hc3b602bf},
  {32'hc4a473c4, 32'hc34f24ce, 32'hc3232fbf},
  {32'h42c08028, 32'hc2f4931f, 32'h4287a22e},
  {32'hc40eca18, 32'hc2f14292, 32'hc2b7f620},
  {32'h44d7a34b, 32'hc2c8d748, 32'h438b0963},
  {32'hc4d86f1e, 32'h41a57b24, 32'hc241b6c2},
  {32'h451ddf96, 32'h4385e673, 32'hc323da22},
  {32'hc50f1c18, 32'hc2fe7b64, 32'hc30e8763},
  {32'h4442edfc, 32'h42dace43, 32'hc1553512},
  {32'hc4d9e4e5, 32'h42c68a60, 32'hc3680fff},
  {32'h42d495e2, 32'h4381f1b4, 32'h41116d3b},
  {32'hc4df579c, 32'h43168271, 32'h428e6fce},
  {32'h4519022b, 32'hc356991c, 32'hc35ec68b},
  {32'hc489490f, 32'h42ed9d6c, 32'hc3e1809e},
  {32'h4489c3fd, 32'hc10d80d0, 32'hc28e7f7b},
  {32'hc42ea734, 32'h41987158, 32'h42a346c2},
  {32'h44fa7151, 32'h43c90ec4, 32'hc3a18afc},
  {32'hc3e4f2e7, 32'hc1f5049a, 32'h42b0e080},
  {32'h449d6332, 32'h438ed41b, 32'h41da271b},
  {32'hc45dd344, 32'h4383ba3a, 32'h4293d158},
  {32'h44b4009a, 32'h428f93d1, 32'h4213a20b},
  {32'hc3aa979a, 32'hc3000a37, 32'h43dd7053},
  {32'h44e9035d, 32'h42dd1a27, 32'hc197f5af},
  {32'hc4df53f5, 32'h3fd61616, 32'h42341fc3},
  {32'h450319e0, 32'hc29b1b82, 32'h42e1dbfb},
  {32'hc4db6170, 32'h40fb61b0, 32'hc2d47858},
  {32'h44fc7dae, 32'hc3ccfb0a, 32'hc3078b5e},
  {32'hc494dea3, 32'h43c9a93d, 32'hc381848f},
  {32'h44c17944, 32'hc2d1ad06, 32'hc342b296},
  {32'hc4a20346, 32'h4347caf6, 32'h43878e9c},
  {32'h43f0ff70, 32'h42cebf05, 32'h43b03eaa},
  {32'hc4eec53b, 32'hc30a5f4a, 32'hc418f1e9},
  {32'h4424a05f, 32'h43a82cff, 32'h432bc17c},
  {32'hc4f06a41, 32'h437d1cc7, 32'hc30eb64f},
  {32'h448f73c1, 32'h44420efb, 32'hc261d3e3},
  {32'hc3367280, 32'h4307a61c, 32'hc2e11c4f},
  {32'h4486b28f, 32'h43094602, 32'h4372f02d},
  {32'hc409cdd4, 32'hc1d389e2, 32'h43173b2f},
  {32'h443c3dd8, 32'h43c461e5, 32'hc40f243a},
  {32'hc4613670, 32'h437a29cc, 32'hc2347e04},
  {32'h44e6bb2d, 32'hc1dd7218, 32'h43557dae},
  {32'hc3bd19a0, 32'h43237760, 32'hc3b9a6dd},
  {32'h450955e6, 32'h42ac3569, 32'hc303431a},
  {32'hc4f96bcc, 32'h43d8981d, 32'hc3229a06},
  {32'h4518083e, 32'h428d35c0, 32'hc2c63681},
  {32'hc4c9fa3a, 32'hc3119269, 32'hc27dba70},
  {32'h4404bb91, 32'hc21b8ec3, 32'hc351f513},
  {32'hc50e1877, 32'h4392c452, 32'h42b2ed9f},
  {32'h44f66b82, 32'hc301da21, 32'h42ea1f65},
  {32'h4326dacb, 32'h432c8d11, 32'h4328bd4b},
  {32'h43cdcebc, 32'hc25de37e, 32'hc3abcb4d},
  {32'hc4cc449a, 32'h43284d40, 32'hc38bca8c},
  {32'h439598b6, 32'h433df03f, 32'hc0c939a6},
  {32'hc5079ca8, 32'hc31aac3a, 32'h42c2e600},
  {32'h44067fb0, 32'h4282c6ff, 32'hc42a716e},
  {32'hc44d8c82, 32'h42f6cefb, 32'h437e311b},
  {32'h4505d562, 32'h43116bfe, 32'h40a5b547},
  {32'hc50a41f4, 32'hc1795ccc, 32'h4381db4a},
  {32'h4397ec48, 32'hc28da900, 32'hc30bf8f4},
  {32'hc23557d0, 32'hc3ba254f, 32'h432a212a},
  {32'h447372b7, 32'h439319e8, 32'hc360de5b},
  {32'hc44a4dce, 32'h4353f3f1, 32'hc30e5e4f},
  {32'h44025ad0, 32'h4351d698, 32'hc2936c49},
  {32'hc4ec1b8e, 32'h418813ee, 32'h4262fc7f},
  {32'h45145ce1, 32'h431678c1, 32'h433de24c},
  {32'hc4c18e10, 32'h43c7806b, 32'hc18495f5},
  {32'h44a53707, 32'hc357d5f0, 32'hc30ece0b},
  {32'hc49e6d24, 32'hc16aec40, 32'hc1ece8ca},
  {32'hc3598396, 32'h43010c31, 32'hc2db24e4},
  {32'hc48929c2, 32'hc342b962, 32'h41df672f},
  {32'h44d8c333, 32'hc189ef3a, 32'h42e127a4},
  {32'hc42ebcf5, 32'h3f2ae7d8, 32'h427c9c2d},
  {32'h44702aa8, 32'h4338b219, 32'hc3f39185},
  {32'hc426d7fa, 32'hc0d94478, 32'hc2743594},
  {32'h44ae54cc, 32'h43934114, 32'hc33cce4e},
  {32'hc3574e9c, 32'hbfdc6a1c, 32'h43a6c1ce},
  {32'h447f5058, 32'h43cda1b9, 32'h43dc3084},
  {32'hc4b99c5c, 32'h4386dc5f, 32'h437be2fb},
  {32'h4507dfa6, 32'h4399d3be, 32'hc2e66384},
  {32'hc4a854ba, 32'hc310e738, 32'hc380d44d},
  {32'h450ea001, 32'h434cdb20, 32'h4310ea58},
  {32'hc41d6138, 32'hc14e6417, 32'h435da6b2},
  {32'h44d5aeea, 32'h4197bcca, 32'hc1bacad9},
  {32'hc46e175a, 32'hc42eebf5, 32'h4281964d},
  {32'h44df8a8e, 32'h43d7f19a, 32'hc2d3907a},
  {32'hc3504bf0, 32'h43557bb9, 32'h435227c3},
  {32'h44c69b81, 32'hc2a9f8fe, 32'hc2b4d4d5},
  {32'hc491f9c4, 32'hc30c9e25, 32'h426d5e3a},
  {32'h444d7cd7, 32'hc1338aa0, 32'h43467a3e},
  {32'hc45f6d7a, 32'hc3442232, 32'h42ed7bcc},
  {32'h4441ece6, 32'h439d3fb5, 32'hc391b780},
  {32'hc4d60eab, 32'h43ab0de0, 32'h435c0006},
  {32'h441960f4, 32'h4358ed08, 32'hc2b27ee3},
  {32'hc3c66faa, 32'h42af053c, 32'h43891a26},
  {32'h44501d64, 32'h42f33627, 32'hc327de90},
  {32'hc3bc32e2, 32'hc3e39225, 32'h43077a7a},
  {32'h44e383ec, 32'hc28c7a2c, 32'hc3722bc5},
  {32'hc4f6b60b, 32'h43275a00, 32'h438d6f5d},
  {32'h44da0268, 32'h43a5adce, 32'h42d0cbaf},
  {32'hc4a40749, 32'h4394d99b, 32'hc1e35fdc},
  {32'h4183eaa0, 32'hc3cae8e8, 32'h43860904},
  {32'hc4975626, 32'h431e4534, 32'h43af1a73},
  {32'h44ff9d56, 32'hc23ca08f, 32'hc39a1774},
  {32'h434060e8, 32'hc2e35478, 32'h436277cb},
  {32'hc3b623e4, 32'hc34179ce, 32'h43a6db1f},
  {32'h44179b9c, 32'h41d718da, 32'h4314fdf7},
  {32'hc48db326, 32'h42a613d3, 32'hc29d0253},
  {32'h44449abc, 32'h440c9cff, 32'hc33fb9f0},
  {32'hc1c31860, 32'hc32611f4, 32'h42e1e7ab},
  {32'h4475aa5b, 32'hc33ec940, 32'h432ee5b0},
  {32'hc4f0e5a2, 32'hc33745fb, 32'h42c470f4},
  {32'h44f8f104, 32'h42234fb3, 32'h4331264e},
  {32'hc484f326, 32'h42a50c25, 32'hc3af2248},
  {32'h4496d900, 32'h433c826f, 32'hc35681c0},
  {32'hc4d7b1cb, 32'h42aad456, 32'hc339a234},
  {32'h4457edfc, 32'hc359fa9e, 32'hc29c8826},
  {32'hc408db7b, 32'h428e3f71, 32'h43f42527},
  {32'h44e9b92c, 32'hc335d0aa, 32'h42be5f69},
  {32'hc485010d, 32'hc3c629ca, 32'hc213d967},
  {32'h44faeff9, 32'h4306349d, 32'hc3ee8b1b},
  {32'hc500a5a3, 32'h43a0b857, 32'hc39d90ec},
  {32'h4509303b, 32'h4381e279, 32'h43452455},
  {32'hc4b7ba1e, 32'hc30585bb, 32'hc38c77c0},
  {32'h446f30e9, 32'h43b41a0e, 32'hc2ea4730},
  {32'hc450e6ca, 32'hc2b6a4c9, 32'hc3b32028},
  {32'h433d193a, 32'hc2a60ab4, 32'hc3558a89},
  {32'hc47b7769, 32'hc2fba67e, 32'h426a6c7c},
  {32'h44e18486, 32'h43124ea4, 32'hc330ff32},
  {32'hc466645c, 32'h42a19988, 32'h4335bbfe},
  {32'h4504ed2e, 32'hc3f05504, 32'h42c60558},
  {32'hc493131c, 32'h436d3269, 32'h41253ce6},
  {32'h44a28310, 32'hc1b8af6d, 32'hc402b0bc},
  {32'hc4fe39aa, 32'h436e0680, 32'hc3b6a44c},
  {32'h44ac24ff, 32'h41fc2361, 32'h41b14bc6},
  {32'hc3941e68, 32'hc386fa53, 32'h4322878f},
  {32'h44ccfa65, 32'h42878407, 32'h43ae326f},
  {32'hc510b04b, 32'hc31b842a, 32'hc281510c},
  {32'h4510f740, 32'hc39ae8a8, 32'h42acd96e},
  {32'hc4dd8d05, 32'hc2b345f6, 32'hc21d5387},
  {32'h44425c48, 32'hc3fe74c0, 32'hc291e9ed},
  {32'hc3be258c, 32'h4346459d, 32'hc2a309a2},
  {32'h44eb7599, 32'hc409d592, 32'h4393b809},
  {32'hc47f403a, 32'hc1f8d8c3, 32'hc3096ba5},
  {32'h4438a6ba, 32'hc3713444, 32'h439d0007},
  {32'hc4dc6e9a, 32'h42a0fd03, 32'hc2c37b57},
  {32'h44e19603, 32'h438e9f92, 32'h43b4a148},
  {32'hc49076c5, 32'hc3d2ab26, 32'h43ecd589},
  {32'h44da8ec1, 32'hc30c2461, 32'hc3151db4},
  {32'hc483143b, 32'hc40f6ead, 32'hc34cc4cc},
  {32'h44db634e, 32'hc29a7e10, 32'hc356caff},
  {32'hc50f1cac, 32'h42981c67, 32'hc2a35339},
  {32'h43ef8a3c, 32'h4219799a, 32'hc30a445c},
  {32'hc4a564ee, 32'h40be6820, 32'h422817ca},
  {32'h44eeffd4, 32'h42fd5993, 32'h4370fe2e},
  {32'hc422a1f3, 32'hc3cd028d, 32'hc28e8ac6},
  {32'h450a2835, 32'hc28178b7, 32'h43414c21},
  {32'hc409923d, 32'hc323fcad, 32'h4305bb9f},
  {32'h448a3494, 32'hc2c40dc6, 32'hc3e391ba},
  {32'hc4cc9d3b, 32'hc31ede68, 32'hc310b14b},
  {32'h43241258, 32'hc39480eb, 32'h4371a340},
  {32'hc4c2101d, 32'h42ee99ab, 32'hc39fe66e},
  {32'h44a8fc49, 32'hc3513a94, 32'h44174624},
  {32'hc4bc9bae, 32'h42abf956, 32'hc234b949},
  {32'h447f1c90, 32'hc427d377, 32'h41970b9e},
  {32'hc5051df9, 32'h440ab3c1, 32'hc30e1c88},
  {32'h44db020b, 32'hc3eb48c1, 32'h42cbf545},
  {32'hc50a7e95, 32'h43e52c68, 32'hc3a3a08d},
  {32'h442b522e, 32'hc19ee09e, 32'hc20d7995},
  {32'hc49a1dde, 32'h43f55d3f, 32'hc3f82a7f},
  {32'h4445fe72, 32'h441e57b2, 32'hc1113d62},
  {32'hc47b2745, 32'hc34e7287, 32'hc1a78997},
  {32'h450ec3bd, 32'h43e1a001, 32'h438533c5},
  {32'hc4f3a96d, 32'h42ce4f6e, 32'h43a6e241},
  {32'h44f49e50, 32'hc3aef67e, 32'hc2746d42},
  {32'hc497445e, 32'h434a23b7, 32'hc345b264},
  {32'h447264f6, 32'hc38a2c2b, 32'h440d663b},
  {32'hc4e88eac, 32'h419c45a4, 32'hc35f2b57},
  {32'h438c2e3a, 32'h42b828aa, 32'h43a118d7},
  {32'hc4e84724, 32'hc39f71d5, 32'h416bba86},
  {32'h446cdeea, 32'h4207372d, 32'h435616a2},
  {32'hc4990549, 32'h43a56bde, 32'h42d92d9e},
  {32'h44479ae8, 32'hc3be432b, 32'hbfb79040},
  {32'hc50e2304, 32'h42814205, 32'hc30bf84a},
  {32'h448f2e04, 32'hc113fbc6, 32'h433722c0},
  {32'hc40d52fe, 32'h3f14e520, 32'hc273d48b},
  {32'h4504920c, 32'h41eaf41a, 32'hc3c0d14f},
  {32'hc4de1190, 32'hc2dd1486, 32'hc321e1a9},
  {32'h43efe33d, 32'h438c79fe, 32'h42f645af},
  {32'hc42ea13c, 32'hc0a1dd9e, 32'h43d51c8a},
  {32'h45046b73, 32'hc30367c4, 32'hc1d2b57d},
  {32'hc3862c28, 32'hc35b5806, 32'hc27936be},
  {32'h44ed2f2e, 32'hc14a820d, 32'h424367f5},
  {32'hc3d2df42, 32'hc243a220, 32'hc3014002},
  {32'h445e9de9, 32'h42ea4a49, 32'h4105f9f2},
  {32'hc469556e, 32'h4309e68d, 32'h41a6dfdb},
  {32'h45171947, 32'h4324af8e, 32'h43b1bef4},
  {32'hc47ede36, 32'h4311eb12, 32'h432d53b2},
  {32'h44036d78, 32'h438654ff, 32'h43282af0},
  {32'hc42372e8, 32'hc39ac2f7, 32'h4298ffc0},
  {32'h44a4c865, 32'hc2c75c73, 32'h43e2977d},
  {32'hc4b2b3a1, 32'hc165485f, 32'hc3075afb},
  {32'h44f59955, 32'h43770cc3, 32'hc3e87bd5},
  {32'hc51a2ea2, 32'hc35681ee, 32'h43eee614},
  {32'h43eea05a, 32'hc2da360e, 32'hc36020c2},
  {32'h432918c0, 32'h435d276c, 32'hc1f1da32},
  {32'h450792fe, 32'h42dbcb03, 32'hc2ed7868},
  {32'hc3ea6828, 32'hc3babdb8, 32'h42e51844},
  {32'h45062226, 32'hc308f25e, 32'hc363d473},
  {32'hc49af19c, 32'hc0fbe8c5, 32'hc28f5f31},
  {32'h450f1c60, 32'h43ad3c51, 32'hc14146e8},
  {32'hc4ce9677, 32'hc3bdca49, 32'hc25d6344},
  {32'h4493742a, 32'h43032dbe, 32'h42a07213},
  {32'hc3b85150, 32'h442f8023, 32'h43423de1},
  {32'h4280b058, 32'hc3879b72, 32'hc2855de5},
  {32'hc3c57950, 32'h43835294, 32'hc309a900},
  {32'h44757bce, 32'hc431be1c, 32'hc27eb1e9},
  {32'hc50a5b3a, 32'hc3076a57, 32'h43a743de},
  {32'h451e5fd9, 32'hc18ba903, 32'hc375ed1d},
  {32'hc4efa8bc, 32'hc3afa481, 32'hc17e823e},
  {32'h44f11f9d, 32'h43de91ea, 32'hc2fbea60},
  {32'hc4d43f0f, 32'hc1ebea07, 32'h427413df},
  {32'h441d9dc9, 32'h4384b071, 32'h4333f81f},
  {32'hc4557e98, 32'h40fdf9ea, 32'h43cae6cb},
  {32'h4337bf28, 32'hc20da2dc, 32'hc316d011},
  {32'hc4b9385d, 32'h433f0bf5, 32'h4361a82c},
  {32'h445ba1c8, 32'hc1f498b9, 32'h4386f040},
  {32'hc4bb769f, 32'h43c78740, 32'h4310197b},
  {32'h44e717c1, 32'hc2e2f888, 32'h4237c885},
  {32'hc502a440, 32'h439057bf, 32'h424d68ee},
  {32'h4384a0da, 32'hc3882850, 32'hc2ed4bda},
  {32'hc4035598, 32'hc3321a09, 32'hc30fc01d},
  {32'h4473d701, 32'h42d63c7a, 32'h41cc443b},
  {32'hc4892e9e, 32'hc3b4cc68, 32'h439d6f76},
  {32'h44ba4386, 32'hc27a617d, 32'hc306755b},
  {32'hc4dd5667, 32'hc35637a6, 32'h4317d7b1},
  {32'h4502e52b, 32'h439b63a5, 32'hc2381880},
  {32'hc4030ef5, 32'hc26c4647, 32'h4208bb8c},
  {32'h45012dbf, 32'h427ef084, 32'h425b8d6e},
  {32'hc4c5e6cc, 32'h40cbccd2, 32'h42df2a4a},
  {32'h450002d2, 32'hc2a3f4dc, 32'h434d6b07},
  {32'hc4b15d6b, 32'h410932ea, 32'h439650cc},
  {32'h430f52c8, 32'hc25781fe, 32'hc05f3e3c},
  {32'hc5011622, 32'h4285dfe6, 32'h431518aa},
  {32'h43890794, 32'hc310ab96, 32'h43238563},
  {32'hc475c146, 32'h42a80e68, 32'hc212d57e},
  {32'hc378c752, 32'hc31f4f5c, 32'hc345441e},
  {32'hc3bc7b08, 32'h42bf2074, 32'h43c09bee},
  {32'h44d9bfe2, 32'hc2b8ce6c, 32'h42ff5c0b},
  {32'hc49fd578, 32'hc2ac7ee3, 32'h431f94a9},
  {32'h44411a47, 32'hc23b526d, 32'hc2d44099},
  {32'hc4711ea4, 32'h438bece6, 32'h435756f4},
  {32'h44b5cbfa, 32'hc38882aa, 32'hc35385b4},
  {32'hc44eee64, 32'h43347a64, 32'h43aecb94},
  {32'h4386872c, 32'hc2c398ab, 32'hc2f1691e},
  {32'hc499c5d3, 32'h42be12fa, 32'h432c3e3c},
  {32'h44acdf57, 32'h4294d9cf, 32'hc31c4fc7},
  {32'hc517eee6, 32'hc305a357, 32'hc2e8d589},
  {32'hc221bf10, 32'hc29d8a8f, 32'h42e5fe01},
  {32'h4330e7f0, 32'hc1e7abfc, 32'h4399dbab},
  {32'h44eb7558, 32'h404b8ac0, 32'h410d2d30},
  {32'hc5125bc5, 32'hc3db2312, 32'hc406c74b},
  {32'h44cb5e95, 32'hc394c24f, 32'h436d22b1},
  {32'hc4bc17ff, 32'hc321ebfb, 32'hc30d8d6f},
  {32'h44f72c0e, 32'hc22ff537, 32'hc2e5238f},
  {32'hc4f47d47, 32'hc3a917d2, 32'h43471765},
  {32'h4469523a, 32'hc38d34bd, 32'h42e89dc1},
  {32'hc50a5761, 32'h432a9f19, 32'hc2dc2ba3},
  {32'h44e7940c, 32'hc2809a08, 32'hc3913831},
  {32'hc50f587d, 32'hc3b442de, 32'hc0926934},
  {32'h4446bc3f, 32'h41d2b2dc, 32'hc18d3a82},
  {32'hc4f9720e, 32'hc20b7d7f, 32'hc3a0f4ba},
  {32'h44e9698b, 32'hc3d17598, 32'h43284562},
  {32'hc4f09a61, 32'h432f6946, 32'hc20d098a},
  {32'h428462ec, 32'hc231cfbc, 32'hc3182d76},
  {32'hc259f885, 32'h414e40dd, 32'hc1f3923e},
  {32'h4422afd0, 32'hc1eb28aa, 32'h436b84ce},
  {32'hc4965fec, 32'hc3aee1b7, 32'hc3d9bd59},
  {32'h4440d883, 32'hc300a2e9, 32'hc22f2ebf},
  {32'hc3f22e59, 32'h432471bf, 32'hc38705f1},
  {32'h441ca07b, 32'hc2ad7b43, 32'hc006077c},
  {32'hc40db2ca, 32'hc28371ab, 32'hc3496d5e},
  {32'h4458ba73, 32'hc2e08952, 32'hc1f55d64},
  {32'hc4f3e2ad, 32'hc3870142, 32'h42fe21ba},
  {32'h4510ee17, 32'hc419057a, 32'h42792e88},
  {32'hc4ded8a0, 32'h4392ed8b, 32'h433c30e1},
  {32'h44f956e4, 32'hc3404b23, 32'hc39f2d1a},
  {32'hc4a9580a, 32'hc30c95ec, 32'hc2b8df54},
  {32'h44fc6ab0, 32'hc3da32a7, 32'h4390727b},
  {32'hc4702c08, 32'hc308afd9, 32'hc3a304af},
  {32'h448a202a, 32'h42d0ce0a, 32'hc31d7c73},
  {32'hc4f44bb2, 32'h42b3f632, 32'h42200bf4},
  {32'h44e6f0cf, 32'hc3b2495c, 32'h42779b0f},
  {32'hc473c082, 32'hc3db3ae8, 32'h41582dd3},
  {32'h44f28655, 32'h438e5094, 32'hc284f0e4},
  {32'hc4aed63a, 32'h42490300, 32'hc31e7aef},
  {32'h43f4f106, 32'h42b6758e, 32'h42d055fd},
  {32'hc4c27fc2, 32'hc292c20f, 32'hc2d435eb},
  {32'h4400d020, 32'hc33883a1, 32'h43187baa},
  {32'hc3ac54cc, 32'h42b6c8ce, 32'hc2c89142},
  {32'h441d1096, 32'h40b9bda9, 32'hc3860ff0},
  {32'h432a6f10, 32'h42cbcd60, 32'h42d10b86},
  {32'h44cfc138, 32'h4310fd4e, 32'h43a86264},
  {32'hc463e10c, 32'hc35cb85c, 32'hc2e86e59},
  {32'h44699ab4, 32'hc3ba25c9, 32'h43d88b66},
  {32'hc50660ae, 32'hc3b85e46, 32'h439b241f},
  {32'h4438587b, 32'hc3649189, 32'h4338517d},
  {32'hc466d3d5, 32'hc2b9bd60, 32'h431180b9},
  {32'h4504b0da, 32'h432b3f38, 32'hc3368400},
  {32'hc4a17645, 32'h440ecac1, 32'hc30fdf36},
  {32'h44f2cc3d, 32'hc4059e16, 32'hc149cd40},
  {32'hc518ea21, 32'hc2a5030a, 32'hc3d8734c},
  {32'h4445f3bd, 32'hc1c9702a, 32'hc39273e6},
  {32'hc50421ac, 32'hc3195640, 32'h43a77eaf},
  {32'h4372ce70, 32'h42d6d3a2, 32'h439bee26},
  {32'hc48ab483, 32'hc20707e5, 32'h4337c7cb},
  {32'h443b3554, 32'h435154ae, 32'h41869dcd},
  {32'hc501cbac, 32'h42a9074c, 32'hc1bd0852},
  {32'h44e15842, 32'h425ca90b, 32'h436f6a27},
  {32'hc4f6edc6, 32'hc31d4a60, 32'h4126b137},
  {32'h4505803f, 32'h42c3ccbe, 32'hc24da333},
  {32'hc4fb0749, 32'h4345ddc1, 32'hc2c031f5},
  {32'h44fd77a0, 32'h43635984, 32'hc3314876},
  {32'hc48da6be, 32'hc338ef04, 32'hc3653612},
  {32'h443db738, 32'hc151f817, 32'hc34ae6d6},
  {32'hc3db3718, 32'h442792d0, 32'hc2dfd9ce},
  {32'h44ce001d, 32'hc3357be1, 32'hc35645e9},
  {32'hc4415361, 32'hc29b309f, 32'h42e113a9},
  {32'h4500497f, 32'hc4151649, 32'h441aa14a},
  {32'hc4475280, 32'hc2c852de, 32'h42fb5d90},
  {32'h4378d5d4, 32'h438c0bef, 32'hc3bd7aea},
  {32'h431cd850, 32'h4261afba, 32'hc3d5f1bd},
  {32'h44cd3795, 32'hc3291cf9, 32'hc28b6c9f},
  {32'hc4409cf0, 32'h42e3df66, 32'hc30414a4},
  {32'h447e5c68, 32'h43c99921, 32'h424287e1},
  {32'hc4e42218, 32'hc2e9d5c4, 32'hc31b13d2},
  {32'h43fc99c8, 32'hc22f76c3, 32'h42f8a527},
  {32'hc484e9d0, 32'hc2ca16f9, 32'h41dcc79d},
  {32'h43bb3a18, 32'h3eb4b240, 32'hc2058ff8},
  {32'hc4c644da, 32'hc31aa3d8, 32'h437d93d6},
  {32'h44f037ef, 32'h4349136c, 32'hc2c433bc},
  {32'hc40b8d44, 32'hc23dcce6, 32'h435bc579},
  {32'h4502019e, 32'h43520a56, 32'h4371efc2},
  {32'hbe1a9400, 32'hc39355bf, 32'h4401d117},
  {32'h44e642b4, 32'h42a745b6, 32'hc3e8758f},
  {32'hc37eb884, 32'hc3375000, 32'hc2c70f28},
  {32'h442a894e, 32'hc2bb9f53, 32'hc363ada3},
  {32'hc3e21216, 32'h42a95d8f, 32'hc2a7033b},
  {32'h44909809, 32'h41748d4e, 32'h42a94d97},
  {32'hc3e0c365, 32'hc0f2ea7a, 32'hc2cec0ce},
  {32'hc246c250, 32'hc3bd23f2, 32'h4341d24b},
  {32'hc4c681ee, 32'hc38c4738, 32'h439ac20b},
  {32'hc3e84fb4, 32'h41ee5f40, 32'h436b9a38},
  {32'hc42a32c4, 32'hc34301aa, 32'hc2a3da11},
  {32'h443961e2, 32'hc0727328, 32'hc254e1e4},
  {32'hc40ade80, 32'hc20bcdfb, 32'hc37728e9},
  {32'h44ad4212, 32'hc38fb9f7, 32'hc190147f},
  {32'hc42deac4, 32'h43f4670c, 32'hc209866c},
  {32'h4418609e, 32'hc32c1390, 32'h42b7308b},
  {32'hc4327228, 32'hc35cd3a5, 32'hc3fa0571},
  {32'h44a844f1, 32'hc2ab9f29, 32'hc29db49b},
  {32'hc4f680a5, 32'hc055bc7a, 32'h432148af},
  {32'h449c8909, 32'h4407eb0b, 32'hc334f4d3},
  {32'hc4e9b483, 32'hc38333f8, 32'hc221ef11},
  {32'h45093fc9, 32'hc28d789c, 32'h433cc35a},
  {32'hc4a4c3fe, 32'hc3291386, 32'hc28ea7c6},
  {32'h4490f10c, 32'hc2e567a9, 32'hc391b0b0},
  {32'hc513dcbc, 32'hc308febe, 32'hc3161c24},
  {32'h4402f766, 32'h44038ddc, 32'hc34eaf35},
  {32'hc4caf6d1, 32'hc2fb3dc1, 32'hc119e821},
  {32'h44d060c7, 32'hc3107aad, 32'hc2485e9c},
  {32'hc50581b1, 32'hc25d199f, 32'h4333dd11},
  {32'h4513f15e, 32'h429ba942, 32'hc2586773},
  {32'hc48c9e00, 32'h4313a4b0, 32'h435ea01a},
  {32'h4470e71a, 32'h42906252, 32'hc1c5f069},
  {32'hc4afe901, 32'hc37e7b9d, 32'h4320da9a},
  {32'h44accfa9, 32'hc320719a, 32'hc31b7839},
  {32'hc50bce38, 32'h42b3c044, 32'hc3b56a2d},
  {32'h44929c4e, 32'hc380b51b, 32'hc3a56b64},
  {32'hc4ca49ec, 32'hc30b8113, 32'h43486af5},
  {32'h44e19bee, 32'hc0d6916a, 32'hc2b9c3c6},
  {32'hc35c43d0, 32'hc25c7c75, 32'h43ae3008},
  {32'h44fed130, 32'h431e1a80, 32'hc2b8b854},
  {32'hc4f8fa9a, 32'hc308ac0c, 32'h42e28460},
  {32'h432e7e1b, 32'hc35e6a5b, 32'h423acbd3},
  {32'hc497ee99, 32'hc3dd6472, 32'hc3724fc1},
  {32'h44b77432, 32'h4387105f, 32'h439c2902},
  {32'hc45e0978, 32'hc3eea3e8, 32'h4359234a},
  {32'hbfc4f400, 32'hc2220be8, 32'h432b69a3},
  {32'hc111d6a0, 32'h431311a9, 32'h43272476},
  {32'h44897f0e, 32'h432aad0a, 32'h42f84326},
  {32'hc4eb5fc2, 32'hc39acb05, 32'h422b3c2c},
  {32'h4405fff9, 32'hc3ba0f74, 32'hc33a5395},
  {32'hc17f5f80, 32'hc33e5ea0, 32'hc28f8c7b},
  {32'h43feb840, 32'hc2c2aa0e, 32'hc2c7c543},
  {32'hc39c2675, 32'hc2c6c0e9, 32'hc1a1d429},
  {32'h443ebc58, 32'hc21e3a4a, 32'hc34dc84d},
  {32'hc409c17a, 32'h43993503, 32'h43771c4d},
  {32'h442325c9, 32'hc2e1f973, 32'hc38703a7},
  {32'hc4938fc9, 32'hc214290d, 32'hc33196d3},
  {32'h44c82c7b, 32'hc1f9c1ad, 32'hc2b3bd8c},
  {32'hc202bbb8, 32'h43ad9b55, 32'hc396272b},
  {32'hc2b14ab4, 32'h41b27942, 32'h436034aa},
  {32'hc4f13fce, 32'hc19040a1, 32'h42f44ac5},
  {32'h441012c0, 32'hc2fd4032, 32'hc3ed3fe3},
  {32'hc3eb3f18, 32'h42e85607, 32'hc2de9682},
  {32'h43606e08, 32'hc38cd00a, 32'hc12d2212},
  {32'hc3db5368, 32'h429fcadf, 32'h433b68c0},
  {32'h44c874ce, 32'h423bc029, 32'hc2ea65fb},
  {32'hc516426d, 32'h439ba8b4, 32'hc4200f25},
  {32'h44110a2c, 32'h438d40be, 32'h4313734f},
  {32'hc50287bb, 32'hc293a348, 32'hc28054e6},
  {32'h4516aca2, 32'h43e96e9f, 32'h4400c352},
  {32'hc2102e54, 32'h437a5787, 32'h43663387},
  {32'h44c03fce, 32'h428a9b5b, 32'hc3237afc},
  {32'hc4f2ec67, 32'h43283ffa, 32'hc1bcaf90},
  {32'h4491dce0, 32'hc38325ab, 32'h412d3cb2},
  {32'hc3cd2b90, 32'h4340b90d, 32'hc3515958},
  {32'h44e2c9b9, 32'h43a321cc, 32'h43fb746e},
  {32'hc4c4a087, 32'hc3790c7a, 32'h437ada48},
  {32'h446637c0, 32'h43dc6879, 32'hc23594e6},
  {32'hc43d9bf0, 32'hc2dc4275, 32'hc095b812},
  {32'h4402e72a, 32'hc3c7ff54, 32'h435adc21},
  {32'hc50c937f, 32'h431a661a, 32'h43e25f9c},
  {32'h4502dde6, 32'hc30630b0, 32'h42accab3},
  {32'hc50b6431, 32'h43c2466a, 32'hc3d7af30},
  {32'h45209ef0, 32'hc3002903, 32'hc28cea3d},
  {32'hc4f8aa8d, 32'h42905cc2, 32'h417f0363},
  {32'h41558aa0, 32'h42ebb22f, 32'h4312a50c},
  {32'hc4fbc87b, 32'hc2b1b62a, 32'hc233337b},
  {32'h44d28427, 32'hc3820178, 32'hc37d4238},
  {32'hc4f030ea, 32'h422b1749, 32'h425a5a51},
  {32'h44ade913, 32'h4036bfc3, 32'h42765706},
  {32'hc4ca9bc2, 32'h435ca2ea, 32'h43687696},
  {32'h44e32830, 32'h430040f5, 32'hc3323025},
  {32'hc466061a, 32'h436050e8, 32'hc1f9694b},
  {32'h451481a1, 32'hc26d144e, 32'hc391b5d4},
  {32'hc5068da8, 32'hc29d1194, 32'h400f42b6},
  {32'h450e5b4b, 32'h431bd2d6, 32'hc392a3cc},
  {32'hc5069efa, 32'hc2d8942f, 32'h41118892},
  {32'h4448fe82, 32'h422cb01a, 32'hc3424bda},
  {32'hc49711ba, 32'hc3bf504f, 32'hc20dba3f},
  {32'h4486e07e, 32'h42172b88, 32'h42af1607},
  {32'hc2e21850, 32'hc2d4a369, 32'hc3426089},
  {32'h44a9efe4, 32'h43033751, 32'h42053a1a},
  {32'hc4d348e1, 32'h4410685e, 32'hc3fea12d},
  {32'h441743c8, 32'h436e565a, 32'hc34ca8d4},
  {32'hc4e6b93c, 32'h439ee656, 32'h43503539},
  {32'h45132d63, 32'h42a06889, 32'hc4117703},
  {32'hc488bd9c, 32'h4302366d, 32'hc38c28fe},
  {32'h449cbdd1, 32'h4377c590, 32'h439ca426},
  {32'hc505ace6, 32'hc30715d9, 32'hc29cc76d},
  {32'h4496f20e, 32'h41f289f8, 32'h43b03ec0},
  {32'hc4664ad4, 32'hc300e166, 32'hc1c971e6},
  {32'h4430d0a5, 32'h42c57ebd, 32'h429e9813},
  {32'hc43e4250, 32'h425df3cb, 32'hc3132c76},
  {32'h449355d2, 32'h4291acba, 32'hc2f8f308},
  {32'hc501c999, 32'hc3979b82, 32'h431f7036},
  {32'h44f471ab, 32'h422b9f9f, 32'h439d7c41},
  {32'hc4efd2b7, 32'hc3303091, 32'h43950a75},
  {32'h4515da1d, 32'h42b8bbaf, 32'hc36dc880},
  {32'hc5052b77, 32'h437650ad, 32'hc2af155c},
  {32'h4421ec80, 32'hc30e74f7, 32'h42760346},
  {32'hc2a88580, 32'h41828a36, 32'h433c1e11},
  {32'h41ffcc80, 32'hc3276f2e, 32'h433c16aa},
  {32'hc4acc6e4, 32'hc330c06d, 32'hc18b4806},
  {32'h449fbf93, 32'h41c36ecf, 32'h4160d408},
  {32'hc4d3ecca, 32'hc3199fcc, 32'hc3182f4d},
  {32'h441a965c, 32'hc1608712, 32'h4295c255},
  {32'hc495bf22, 32'h43a2ff2e, 32'h42aeac4f},
  {32'h44b43b7e, 32'hc18b0c0f, 32'hc28afcb2},
  {32'hc43cc91e, 32'hc2ca72ce, 32'hc2df8e5c},
  {32'h43f8c1c7, 32'h4256ed18, 32'h4416366d},
  {32'hc420077a, 32'h42ba7a01, 32'hc3600f3b},
  {32'h43bb7cfe, 32'h439ccf39, 32'h4383e006},
  {32'hc501c3e3, 32'hc3467315, 32'h42ce22e3},
  {32'h44ef39ee, 32'hc36f4247, 32'h43aa3da1},
  {32'hc50ec592, 32'h42a90e54, 32'h44045e34},
  {32'h44f01e68, 32'h44204f76, 32'hc378479f},
  {32'h42965fa0, 32'h43a5e465, 32'hc359f08a},
  {32'h4387a700, 32'h432a7398, 32'hc3821abc},
  {32'hc483d2d2, 32'hc23ffb9f, 32'h43597277},
  {32'h444f42c6, 32'h43471a1d, 32'hc23091e5},
  {32'hc50d32ea, 32'h42eb4756, 32'h437adbdd},
  {32'h439e31b6, 32'hc173de06, 32'hc1dfa28e},
  {32'hc489c391, 32'hc311222e, 32'hc2d7bf63},
  {32'h450f5017, 32'hc39744a0, 32'h4374418a},
  {32'hc4008320, 32'h440db145, 32'hc2200ef1},
  {32'h45006beb, 32'h41a4ad9d, 32'h4376bcae},
  {32'hc3d9929c, 32'h42794dc9, 32'hc33121e0},
  {32'h425a21a0, 32'hc2afe061, 32'h43082db1},
  {32'hc37610b4, 32'h431a7d6a, 32'h43262dd0},
  {32'h448d2df7, 32'h42982972, 32'hc30aa9a4},
  {32'hc411c8a4, 32'h4419063b, 32'hc21e214f},
  {32'h432d1980, 32'h4335bdf8, 32'hc3f24d1a},
  {32'hc2f0f840, 32'hc26af8f2, 32'hc1a950ee},
  {32'h45113dd6, 32'h42bfe361, 32'hc333e16b},
  {32'hc3a7ba6b, 32'hc304c4b8, 32'hc3131444},
  {32'h44bc6216, 32'hc2d91e23, 32'h436770d0},
  {32'hc5084f17, 32'h42b7f83b, 32'hc2e2c459},
  {32'h4513fb17, 32'h428fd11e, 32'h4186e450},
  {32'hc3dae524, 32'h42e66202, 32'h42e516e5},
  {32'h44fd081b, 32'hc3aca3f3, 32'hc216570b},
  {32'hc4dcb7ee, 32'h42d36e55, 32'h42523293},
  {32'h437b4658, 32'hc18b22ea, 32'hc23a58dd},
  {32'hc3c1f9e8, 32'h43cc0777, 32'hc40067dd},
  {32'h44029663, 32'h41778a11, 32'h438aaa45},
  {32'hc3a5ead8, 32'h43a10e01, 32'hc3bdd8f8},
  {32'h44f274c6, 32'h4333f5a7, 32'h41f667cd},
  {32'hc48cb6aa, 32'h43a66148, 32'hc2fa3a8e},
  {32'h44c4aa89, 32'h43b7a31b, 32'h424940a1},
  {32'hc4558e48, 32'hc2b3fcc9, 32'h42dd1923},
  {32'h44d75186, 32'h430081d6, 32'h42b0dac3},
  {32'hc4ff3e82, 32'h4272fdf3, 32'h42834674},
  {32'h45018af8, 32'hc223a750, 32'hc3a51540},
  {32'h421b1d46, 32'h43d3e548, 32'hc39e2003},
  {32'h43bf97de, 32'h4188cd06, 32'hc29b52e9},
  {32'hc3fc09c8, 32'h4394ecfb, 32'hc220c3cc},
  {32'h438bcca8, 32'h4201b58a, 32'hc322a8b3},
  {32'hc4e498f6, 32'h42b23283, 32'hc087041a},
  {32'h44fda9aa, 32'h438506e2, 32'h43beb89e},
  {32'hc48a699e, 32'h425f8bb4, 32'h422927a1},
  {32'h44c9e9e9, 32'h417474f1, 32'h429b7fa3},
  {32'hc4231ed9, 32'hc2d1f05c, 32'hc1d1c1b1},
  {32'h44fc783e, 32'h42025aff, 32'hc32f0fd8},
  {32'hc4d274b0, 32'h43ed8f27, 32'hc3b55275},
  {32'h43018c7c, 32'hc2f35029, 32'h42bff393},
  {32'hc4d6aaa4, 32'hc25c7eb7, 32'hc33e036f},
  {32'h445bd34c, 32'hc3757df5, 32'h42b72475},
  {32'hc4744648, 32'hc36b362f, 32'hc33065d1},
  {32'h4490acad, 32'hc335c1c6, 32'h42874ddc},
  {32'hc4e47765, 32'hc057493e, 32'h429a295c},
  {32'h44f03f9f, 32'h4209f792, 32'hc3726217},
  {32'hc332e070, 32'hc3952465, 32'hc42a8c92},
  {32'h44d2ec5b, 32'h419bea0a, 32'hc00a0820},
  {32'hc4b634b7, 32'hc33d0171, 32'hc2af2951},
  {32'hc4aa06f7, 32'hc363a794, 32'h4190871a},
  {32'h442ca58e, 32'hc2a8e63b, 32'h433e5dfc},
  {32'hc4bc55d8, 32'h43dee0ea, 32'h431ce145},
  {32'h44ebc762, 32'h43ac1af0, 32'h435067a1},
  {32'hc3ab2e9d, 32'hc3234b93, 32'hc25ded88},
  {32'h4455590a, 32'hc3c6a40d, 32'hc305063b},
  {32'hc4c769ec, 32'hc2941abc, 32'h428d77a3},
  {32'h442289d4, 32'h4369724e, 32'hc39dec26},
  {32'hc4247d64, 32'hc392563f, 32'hc2f4ec44},
  {32'hc2b35a53, 32'hc2a5af27, 32'hc1b22c14},
  {32'hc51cb724, 32'h41db6f46, 32'hc2f393bd},
  {32'h449f639c, 32'hc358709d, 32'h4288aed6},
  {32'hc457ccb1, 32'h42781cff, 32'hc3ace6d4},
  {32'h45025c6a, 32'h43c74b17, 32'h43320394},
  {32'hc4dd2197, 32'h3df2a730, 32'h4302e2df},
  {32'h44e394ce, 32'hc2d2ab28, 32'h42b5eb09},
  {32'hc47112d8, 32'h4103bfeb, 32'hc34e2eeb},
  {32'h4473689e, 32'hc3142920, 32'h428068da},
  {32'hc49e30d7, 32'h435eee23, 32'hc28a5bec},
  {32'h44402ed8, 32'hc36644b4, 32'hc2b527a3},
  {32'hc41c882f, 32'h438b49aa, 32'hc3c8807d},
  {32'h43e84294, 32'h42a2bd71, 32'h42621daa},
  {32'hc4ddc3c2, 32'hc40174e6, 32'h41d9a2d2},
  {32'h43e9e936, 32'h428b9af9, 32'h430821f2},
  {32'hc4f64723, 32'hc3773db2, 32'h4343604f},
  {32'h44d35c78, 32'h429805e0, 32'hc2af3bef},
  {32'hc5066d57, 32'hc2b68428, 32'h43aa71f7},
  {32'h450bda84, 32'h430f5e38, 32'h4326ad57},
  {32'hc5260bea, 32'hc4076d98, 32'hc3a0f791},
  {32'h44d90ae5, 32'h43583a4e, 32'hc2518068},
  {32'hc50a4570, 32'h432655d2, 32'hc35e1f7c},
  {32'h44a84760, 32'hc0c3694f, 32'h4248d100},
  {32'hc3a4fcd7, 32'hc2120fd8, 32'hc30a1d98},
  {32'h448b8655, 32'hc326abe3, 32'hc2a43985},
  {32'hc516a9da, 32'hc2cfa138, 32'h43498df4},
  {32'h44d143dd, 32'hc197fe7c, 32'hc1e6b859},
  {32'hc49b14b4, 32'h4358fcc1, 32'hc36e25f4},
  {32'h44e63561, 32'h4392bbd6, 32'hc287ba8f},
  {32'hc4bd11fa, 32'h4352e5a5, 32'h41975294},
  {32'h450427bf, 32'h42952aa6, 32'hc2da2ab4},
  {32'hc50d249b, 32'hc39303e4, 32'hc3857f0d},
  {32'h449a5b57, 32'hc155f9d6, 32'hc23ce41c},
  {32'hc4ede42a, 32'h41a393da, 32'hc2dbae5b},
  {32'h446d2f7c, 32'h42cb7461, 32'hc418b5b0},
  {32'hc50ab7d6, 32'hc3942e06, 32'hc3a87b83},
  {32'h44496d9e, 32'hc25d11b5, 32'h424a130e},
  {32'hc4b6df08, 32'h43397802, 32'hc31b0ab7},
  {32'h42ff9020, 32'hc16278eb, 32'h43a750f1},
  {32'hc4d41fb8, 32'h43c697fc, 32'hc31c3ac2},
  {32'h45018fe3, 32'hc33fd8f2, 32'hc31df9f6},
  {32'hc4e061ee, 32'h41c526ed, 32'hc222b3da},
  {32'h442158ca, 32'hc228040d, 32'h4291c9b1},
  {32'h43c092a0, 32'h43308b2d, 32'hc31b9ed6},
  {32'h4470e69a, 32'h409cd121, 32'h429e1b53},
  {32'hc50ed726, 32'h43131e61, 32'hc0e459b9},
  {32'h4450d30c, 32'hc39203bf, 32'hc31881f0},
  {32'hc509d8f0, 32'hc3072a29, 32'hc25f7b08},
  {32'h44876806, 32'h438842a2, 32'hc3c05397},
  {32'hc50d2a34, 32'h42f525d2, 32'h405c837d},
  {32'h4332075e, 32'h429568e9, 32'hc3e8ab07},
  {32'hc3a10788, 32'h43c5b62e, 32'hc3f60ebf},
  {32'h43adad1c, 32'hc3e8974a, 32'hc2bd389d},
  {32'hc4ed2bec, 32'h42fa3ab4, 32'hc3376cc2},
  {32'h44e3dce9, 32'h43d4a24e, 32'h42d7a704},
  {32'hc4acf632, 32'hc0e6234a, 32'h44107c25},
  {32'h44d4f0a9, 32'h4348c3e9, 32'hc2723b54},
  {32'hc4e807da, 32'h4332b9dc, 32'h42b5cb9e},
  {32'h44f3b4f6, 32'hc33a3cab, 32'hc41648f1},
  {32'hc502f551, 32'hc2d37955, 32'h430087cd},
  {32'h445a5f24, 32'hc1208c08, 32'h430c75c8},
  {32'hc40cf4a4, 32'hc323a796, 32'hc2d9ba78},
  {32'hc3965cda, 32'hc361931f, 32'hc2ed98b9},
  {32'hc4a11bf6, 32'h42f975cf, 32'hc39ca45e},
  {32'h43eaa8b0, 32'hc34bcf3c, 32'h42631efe},
  {32'hc4dd8558, 32'hc30525e4, 32'hc34af644},
  {32'h434475c2, 32'h4342e0d0, 32'h43884d7b},
  {32'hc35b58e0, 32'hc291b136, 32'h42f073fb},
  {32'h41f6cdc0, 32'h42b8152c, 32'hc3a6e103},
  {32'hc430bcf6, 32'h438a2450, 32'h42c9baee},
  {32'h43dedf2c, 32'hc33e7bc2, 32'h430a4334},
  {32'hc4784eae, 32'hc3ca9fd8, 32'hc20d68bc},
  {32'h44da5323, 32'hc203df70, 32'hbfcc0414},
  {32'hc50fc7da, 32'hc32dd9e2, 32'hc1eb55be},
  {32'h44a4a205, 32'hc3451dfb, 32'h425d1710},
  {32'hc4a08abc, 32'hc16c571c, 32'hc3471bbe},
  {32'h44c55819, 32'h421a5c56, 32'h4363a2f6},
  {32'hc4a7e0ad, 32'h420ce2c7, 32'h42cfc1aa},
  {32'h4473ac18, 32'h4352d018, 32'hc2a0f18e},
  {32'hc500444d, 32'hc251fdab, 32'h416ddd99},
  {32'h443d39c6, 32'h43181236, 32'hc34fd7b6},
  {32'hc487700d, 32'hc3079a3e, 32'h4290ecfb},
  {32'h450fc71c, 32'h43a11056, 32'hc2a4279a},
  {32'h4385f270, 32'hc2f99278, 32'hc3218a1a},
  {32'h450377f8, 32'h43431c84, 32'h425659d3},
  {32'hc447b884, 32'hc2c6d952, 32'hc367e395},
  {32'h450948c8, 32'h4337ab0a, 32'hc29deead},
  {32'h4378960c, 32'hc1848644, 32'h4414411a},
  {32'h43a3ff1e, 32'hc16bc6db, 32'h418831b4},
  {32'hc4d84823, 32'hc21f4e8a, 32'hc31a7ad9},
  {32'h44bc42f5, 32'hc2d90442, 32'hc298ca5a},
  {32'hc4e2f7bb, 32'hc38049a6, 32'h4345d041},
  {32'h429fd540, 32'h42fd1997, 32'h43c9ef84},
  {32'hc43bb9d0, 32'h438b2f16, 32'hc3a623bf},
  {32'h44073c4c, 32'h42459471, 32'h44466409},
  {32'hc4e7fd40, 32'h43210132, 32'h4377119e},
  {32'h44970f80, 32'hc25a6b0f, 32'h42e1eb98},
  {32'hc50580db, 32'h42c6ad9f, 32'hc33b48d6},
  {32'h4488b3d6, 32'hc38b4e18, 32'hc38310c9},
  {32'hc4d14bc0, 32'h41e9fb00, 32'h43a247cc},
  {32'h44f8a211, 32'h43eabaf8, 32'hc13123f0},
  {32'hc4ec05ad, 32'h42ea48fc, 32'h4294ee51},
  {32'h43566070, 32'h430dd046, 32'h432f252a},
  {32'hc4ed771c, 32'h43a4a384, 32'h43e1c4aa},
  {32'h43fce1b0, 32'h4294acef, 32'hc3a5cc71},
  {32'hc48db0e2, 32'h43ef169e, 32'h42ff7994},
  {32'h44efd07c, 32'hc3051fa7, 32'hc347abf0},
  {32'hc4c5e49e, 32'hc20269b0, 32'h434e3e5e},
  {32'h40f8e2c0, 32'h4136324c, 32'hc0fc4e31},
  {32'hc4fcad8f, 32'hc3a98650, 32'h431722c2},
  {32'h4517549a, 32'hc3a43f1d, 32'h4342bc62},
  {32'hc42c9844, 32'hc21f1b21, 32'hc215d5be},
  {32'h44c874bc, 32'h439b986d, 32'h434ee981},
  {32'hc3988dc4, 32'hc2cba4ef, 32'h43ded507},
  {32'h44d16e2c, 32'hc3ac6543, 32'h434df756},
  {32'hc4e7d054, 32'hc38493b6, 32'h42a45f70},
  {32'hc3c76940, 32'hc3dff0db, 32'hc32fdca5},
  {32'hc2aaafc0, 32'hc339736d, 32'hc28f91ee},
  {32'h448c8191, 32'h433d7f64, 32'h43ba332f},
  {32'hc3fbebc4, 32'h4368c0f8, 32'hc29953d1},
  {32'h44dedc12, 32'hc3abce1e, 32'hc22cdde6},
  {32'hc4cb397e, 32'hc2f452a8, 32'h43a531e7},
  {32'hc2bf26f0, 32'h432b3e7a, 32'h43a749af},
  {32'hc4a6fa60, 32'h3f4c59b0, 32'hc375b02f},
  {32'h44f99f04, 32'hc3735bb9, 32'hc30c5eda},
  {32'hc4a750df, 32'hc310e510, 32'h43acd496},
  {32'h44e618e6, 32'hc2a64d1c, 32'hc3cc42f0},
  {32'hc47c086f, 32'hc3c60be1, 32'hc39d8dbf},
  {32'h44df1b6b, 32'hc36a9c92, 32'hc2e020c0},
  {32'hc4723b98, 32'h41575fc0, 32'h4277d3fc},
  {32'h44582088, 32'hc287ff55, 32'hc24df13a},
  {32'hc4a5ff8c, 32'hc2de9f77, 32'h4343f41b},
  {32'h44d3a2cc, 32'hc2285566, 32'h42b59183},
  {32'hc48334e7, 32'h4379ea8e, 32'h43ad2307},
  {32'h44deb422, 32'h42a49fe6, 32'hc212fbce},
  {32'hc5017922, 32'h4053262c, 32'h434afa81},
  {32'h44bfeb99, 32'hc39f1bd9, 32'h42708623},
  {32'hc497317e, 32'hc2f7f4e0, 32'h43a33bf2},
  {32'h44bd3f17, 32'h43877014, 32'hc1ffd248},
  {32'hc0ccd500, 32'h411dc425, 32'h42338079},
  {32'h450f5f50, 32'h43bc3f91, 32'h42774634},
  {32'hc33e2560, 32'h438ce2d1, 32'h42e6aeb6},
  {32'h44d6649c, 32'h430f67e0, 32'h43822d3d},
  {32'hc3f7081c, 32'hc367b60f, 32'hc41707ae},
  {32'h43a344ec, 32'hc25de2ed, 32'hc37a0144},
  {32'hc4b18b37, 32'h433ef07c, 32'hc2dfe0fd},
  {32'h45046b92, 32'h43f1c005, 32'h42ac2cfd},
  {32'hc3815758, 32'hc1cb221a, 32'hc277e73a},
  {32'h44e5986c, 32'hc1f88314, 32'hc3c3069c},
  {32'hc4710367, 32'h4164e7c9, 32'hc362971e},
  {32'h44a26dff, 32'h441e0320, 32'h433e8d83},
  {32'h43a4d454, 32'hc304bbfb, 32'h43a4e933},
  {32'h44d998ec, 32'h43edc6e7, 32'hc204646c},
  {32'hc4b4e41c, 32'h42c93ab6, 32'h4048cd75},
  {32'h44dc817a, 32'h437d6f07, 32'h4221a6aa},
  {32'hc50f619d, 32'hc3ea03ee, 32'h434c41a1},
  {32'h4449acc8, 32'h436f3770, 32'h43800633},
  {32'hc4118bca, 32'h4367a42b, 32'h42fd4c52},
  {32'h446ae578, 32'h435ce04d, 32'h43f90db4},
  {32'hc2355606, 32'hc30a11be, 32'h430ab7ef},
  {32'h43b8b01c, 32'hc2ae7115, 32'h4368d7ba},
  {32'hc3eee9c9, 32'hc2d7e926, 32'h43585746},
  {32'h44b635a2, 32'hc3242e48, 32'hc2bf7686},
  {32'hc5033c5d, 32'hc40f17be, 32'h416e9233},
  {32'h43967830, 32'hc3c09280, 32'h421ec64c},
  {32'hc197ccbb, 32'h43862067, 32'h42adb3cd},
  {32'h44c043e3, 32'hc2d94d6f, 32'h429f04c8},
  {32'hc488e2ca, 32'h43a3a5d6, 32'h42d16568},
  {32'h433a5100, 32'hc3b4cb0d, 32'hc25171bb},
  {32'h411bca00, 32'h43b15c67, 32'hc3ec611b},
  {32'h44e4f1db, 32'hc3667705, 32'hc301c484},
  {32'hc4b9ffc3, 32'h42e8737b, 32'hc3303709},
  {32'h4417f388, 32'h4206c160, 32'h423dd2ac},
  {32'hc4577cf8, 32'hc2a22492, 32'hc3454105},
  {32'h43493ddc, 32'h43541048, 32'h41ca229c},
  {32'hc4ea320e, 32'h41ce533b, 32'hc39bd3bd},
  {32'h44787624, 32'h42cbc857, 32'h43ef435b},
  {32'h42b0bf60, 32'h42ca14d1, 32'hc383f1ac},
  {32'h44ebb47b, 32'hc30b2a7c, 32'h425c14f0},
  {32'hc36e38f8, 32'hc32795cf, 32'hc1e3d765},
  {32'h44c8be53, 32'h4360563e, 32'h435de076},
  {32'hc506ab62, 32'h431bc196, 32'h436ef005},
  {32'h43ea1358, 32'hc23041af, 32'hc285e67d},
  {32'hc493420e, 32'h42dbaf5a, 32'hc3bc6bcc},
  {32'h4450e290, 32'hc3da3c79, 32'hc302a17d},
  {32'hc40d1053, 32'h435e8529, 32'hc3390171},
  {32'h44f65fc5, 32'hc39bc4ff, 32'hc3a06979},
  {32'hc47158a1, 32'h43005c0e, 32'h43247453},
  {32'h43dc4128, 32'hc2b5b26b, 32'hc2fe412c},
  {32'hc5086dc5, 32'hc30d8f43, 32'hc2c842d8},
  {32'hc1cb5100, 32'h440323d6, 32'h43d4468f},
  {32'hc4adcb18, 32'h40dbf7e0, 32'hc253d09b},
  {32'h45009048, 32'h436fcf8d, 32'h43949175},
  {32'hc424dc40, 32'hc3037c30, 32'h430c29d5},
  {32'h416c769c, 32'h43520600, 32'hc3f3f7f1},
  {32'hc4582276, 32'h42f2dcaf, 32'h40857c78},
  {32'h44f93122, 32'hc1c88a06, 32'hc40b34f1},
  {32'hc20cbd50, 32'hc2813c0c, 32'hc2cd37cb},
  {32'h440598f4, 32'hc37d3efc, 32'hc1460118},
  {32'hc4318828, 32'hc28ef1b4, 32'hc2917496},
  {32'h44ccead0, 32'h42f4e5e6, 32'hc3d59072},
  {32'hc4f83397, 32'hc34c52f3, 32'h4381e0d6},
  {32'h43575830, 32'h437626be, 32'hc398bb64},
  {32'hc4070ba5, 32'h439ca1f2, 32'hc21d7217},
  {32'h448614cc, 32'hc3b2a293, 32'hc3437894},
  {32'hc4687bbd, 32'h43f6383b, 32'hc2d6864f},
  {32'h42c83860, 32'hc3bd43cb, 32'hc287904a},
  {32'hc3fb0db5, 32'hc2d94dc5, 32'hc32a551f},
  {32'h44975abb, 32'hc1f79686, 32'hc365ac99},
  {32'hc4c03569, 32'hc28a40b0, 32'h439238bb},
  {32'h44dadf89, 32'hc3859b57, 32'hc31ee16a},
  {32'hc4479aa8, 32'h4288d4c4, 32'h4125a942},
  {32'h450acf59, 32'hc310bbf4, 32'hc15e2d0e},
  {32'hc486b1a3, 32'h44063fc1, 32'hc36a01e2},
  {32'h433f130c, 32'hc32e6113, 32'hc22e2a20},
  {32'hc4add124, 32'h43a99b76, 32'hc3814a7a},
  {32'h44bda277, 32'h438b3b55, 32'hc33fcccc},
  {32'hc3207558, 32'h438bdf33, 32'hc1567d18},
  {32'h44b986fc, 32'h4374fe63, 32'h4286c413},
  {32'hc3594440, 32'hc29ca631, 32'h431f1f2a},
  {32'h448b72b1, 32'h436afaf7, 32'h41fa49b6},
  {32'hc410c31f, 32'hc24c8a31, 32'h42e26660},
  {32'h44c09da6, 32'hc3982d63, 32'hc348338e},
  {32'hc4a0ada6, 32'h42508d9f, 32'hc3236f84},
  {32'h4501ad41, 32'hc40a486e, 32'hc2b2c25d},
  {32'hc3f72410, 32'h42b1bd2c, 32'h4353c0c5},
  {32'h450556c9, 32'hc3f50a08, 32'h43fc07fe},
  {32'hc41afa60, 32'h435a58d8, 32'hc0b1991c},
  {32'h42f1a8e0, 32'hc2e82c50, 32'h42fb5f79},
  {32'hc506f07f, 32'h418f1904, 32'hc34e4daa},
  {32'h444f27a0, 32'hc2cd60a9, 32'h438780d5},
  {32'hc5006c03, 32'hc06403b5, 32'hc0b2057e},
  {32'h44992f30, 32'hc06fc8e6, 32'h41f3311b},
  {32'hc45cdffa, 32'h42bd0262, 32'h41df7082},
  {32'h4505941b, 32'hc356bd0c, 32'h42c33997},
  {32'hc4f6a58d, 32'h43f1cf4d, 32'h43fd34e2},
  {32'h446bff00, 32'h43d40d93, 32'h438be0c8},
  {32'hc505e327, 32'h4387e6aa, 32'hc19e42dc},
  {32'h44da5964, 32'hc144331d, 32'hc24b2c00},
  {32'hc4a72706, 32'h4314460d, 32'hc3ecca1c},
  {32'hc2a748b4, 32'h42e33db9, 32'hc363953a},
  {32'h4272dea8, 32'hc1bfd073, 32'h41b37b25},
  {32'h4504ed6a, 32'hc233e7a0, 32'hc2d7acca},
  {32'hc4c992a9, 32'hc0d33344, 32'h43a7f3e8},
  {32'h4485abf2, 32'hc0abde5c, 32'hc3e4146a},
  {32'hc5041fd4, 32'h43090e45, 32'hc2524dc9},
  {32'h44d1d17d, 32'h42a21158, 32'h43be3735},
  {32'hc43104f4, 32'h433203ba, 32'hc30ae41a},
  {32'h450b8c82, 32'hc3237a2f, 32'hc19cef97},
  {32'hc4b1d940, 32'hc3fe2d63, 32'hc307c586},
  {32'h452df762, 32'h431ad119, 32'hc1edad4e},
  {32'hc4acece0, 32'h43c5d278, 32'h419394f8},
  {32'h44075bac, 32'hc3b1157b, 32'h43132584},
  {32'hc2df7ce0, 32'hc3512b44, 32'hc1261932},
  {32'h44fd2330, 32'h43439bc6, 32'hc345795f},
  {32'hc4432795, 32'hc324d454, 32'hc38dc097},
  {32'h45060d38, 32'h43103e41, 32'hc34d90a9},
  {32'hc43de22c, 32'hc2b1cdfc, 32'hc2f114b0},
  {32'h447b7c97, 32'hc23cccec, 32'h433258d7},
  {32'hc51ad016, 32'hc2819901, 32'h4299daa2},
  {32'h442dd640, 32'hc365d070, 32'h43dfa9fc},
  {32'hc4fbdc5c, 32'hc388ad58, 32'hc2cd3670},
  {32'h4459dc8b, 32'hc387130e, 32'hc2a4dc15},
  {32'hc4dccef3, 32'hc3544d57, 32'hc367201e},
  {32'h44b12136, 32'hc35613aa, 32'h438ace6e},
  {32'hc368f950, 32'h428499c6, 32'hc364749d},
  {32'h4291e000, 32'hc398aedb, 32'hc197f6ab},
  {32'hc44a3508, 32'h43d53220, 32'h42adfff9},
  {32'h449f0445, 32'h440edc6c, 32'h41440ea8},
  {32'hc4e7761c, 32'hc2f040cd, 32'hc3582ce4},
  {32'h4510ed14, 32'hc2d5eb38, 32'h430f9aad},
  {32'hc3d38052, 32'hc3c73276, 32'hc36552bd},
  {32'h44f010ad, 32'h43965de5, 32'hc332c564},
  {32'hc449b7b8, 32'h428483de, 32'h432db83b},
  {32'h441833f6, 32'h436dccbc, 32'hc2fa9c27},
  {32'hc48464b6, 32'hc2c6bff6, 32'hc2f5b8a6},
  {32'h441df8e4, 32'h43784472, 32'hc10892a7},
  {32'hc35fd6e4, 32'hc119977e, 32'hc33c3bca},
  {32'h44568276, 32'hc3d8f9f6, 32'hc200f38a},
  {32'hc509e35f, 32'hc2ef9c62, 32'hc1c2ca4c},
  {32'h44af6ff7, 32'h42f61a93, 32'hc1933ecc},
  {32'hc4fb3c7b, 32'hc28935ec, 32'hc2b148a4},
  {32'h45000511, 32'h43713616, 32'hc256d8eb},
  {32'hc51564b8, 32'hc203f1dd, 32'h435cdb3b},
  {32'h4457fd80, 32'h43cf650b, 32'hc2b810a6},
  {32'hc3ef5ba8, 32'h4356b312, 32'hc2e751ea},
  {32'h44b18d0d, 32'hc321e8be, 32'hc26b5cc3},
  {32'hc519ac11, 32'h430e2ba0, 32'hc3464e32},
  {32'h44bba575, 32'hc3ac9a64, 32'h43501762},
  {32'hc506d523, 32'hc31529ad, 32'h42175cda},
  {32'h44faa07c, 32'h43ad878e, 32'hc360f5ac},
  {32'hc42cb220, 32'hc3359951, 32'h42d94160},
  {32'h44dc1f85, 32'hc33c4e2b, 32'hc383e935},
  {32'hc4e91409, 32'hc3b9d071, 32'hc2362c0b},
  {32'h4518e250, 32'h430928d5, 32'hc380e80c},
  {32'hc44389a2, 32'hc24730fb, 32'hc413965b},
  {32'h4483a9a5, 32'hc18fa299, 32'h4314d927},
  {32'hc4eb2658, 32'hc35a3bcc, 32'hc3f72094},
  {32'h44a39850, 32'hc3b82743, 32'h4403c2ee},
  {32'hc50960a2, 32'h4340760e, 32'h43994320},
  {32'h44e61bd9, 32'hc31b0d44, 32'h4357252a},
  {32'hc4ca6e8f, 32'hc282b18a, 32'h433c2f3c},
  {32'h451e4018, 32'hc281d451, 32'hc212ebf7},
  {32'hc4d36938, 32'hc143966c, 32'hc3e1edb5},
  {32'h4500ed0a, 32'h428d1cac, 32'h440b9035},
  {32'hc47050ec, 32'hc38409af, 32'hc1578631},
  {32'h4424ab27, 32'hc3be9dff, 32'h42033de1},
  {32'hc45eac81, 32'h4160567e, 32'hc3863c48},
  {32'h4348a768, 32'hc30f23a1, 32'hc3206187},
  {32'hc359ca18, 32'h43bc8c9d, 32'hc280a5b2},
  {32'h43d07b00, 32'hc1c2a232, 32'h41d5f57d},
  {32'hc4f01ad9, 32'h410211bf, 32'hc39e5d64},
  {32'h44385642, 32'hc39967ca, 32'hc378159a},
  {32'hc4d5fb65, 32'hc34a2c2b, 32'hc3d46266},
  {32'h43c3aea1, 32'hc3b7747c, 32'h43b8602f},
  {32'hc4e6fe31, 32'h4274531f, 32'h4206463e},
  {32'h4512ba69, 32'hc319b965, 32'hc3ae549f},
  {32'hc4b99eae, 32'hc33fdf5d, 32'h422e1eda},
  {32'h44f247c2, 32'hc2c41a32, 32'h4384315d},
  {32'hc4fbe99c, 32'hc217389c, 32'h4318dccf},
  {32'h452291f9, 32'h4287954c, 32'h429e06c1},
  {32'hc4dec057, 32'hc38f2151, 32'hc2e3560b},
  {32'h4448f854, 32'hc3be15e5, 32'h435b40a1},
  {32'hc4f23bcf, 32'hc2049e76, 32'hc396fcae},
  {32'h4500f4c8, 32'hc32f3904, 32'hc34b7d66},
  {32'hc476adc4, 32'h4385570f, 32'h434d3661},
  {32'h449d89f7, 32'h42b3801b, 32'hc1aafda7},
  {32'hc4b942f4, 32'h4410250f, 32'h42972f65},
  {32'h445b4bb3, 32'h42a64195, 32'hc3c0b2c1},
  {32'hc4c94b62, 32'h4267714f, 32'hc1d75c3c},
  {32'h445932cc, 32'hc36ecf95, 32'h425bcbd6},
  {32'hc4e692ca, 32'hc337c627, 32'h43bf4f00},
  {32'h450ad5d5, 32'hc0f66e3d, 32'h437a8d4e},
  {32'hc4b22858, 32'h40ad9959, 32'hc1b7bd9f},
  {32'h447e1714, 32'hc219a05c, 32'h42793413},
  {32'h42af7b40, 32'h4317d257, 32'hc28f2ee8},
  {32'h44029a70, 32'h42d87afa, 32'hc31bf018},
  {32'hc4c1e67c, 32'h4324d704, 32'h407a89e0},
  {32'hc13abe00, 32'hc43810bf, 32'h42edea89},
  {32'hc42ef898, 32'h430ab241, 32'h42cf2532},
  {32'h450875af, 32'h434b2cec, 32'hc39d566e},
  {32'hc48b2875, 32'h42be35c2, 32'h4304f7a8},
  {32'h44fd86fa, 32'hc39ec20b, 32'hc3d3d95c},
  {32'hc481b316, 32'h4376689f, 32'hc3c2bcd2},
  {32'h43c4fc06, 32'h4331f52b, 32'hc054ed1e},
  {32'hc4fc6820, 32'h42ccd177, 32'h433abc74},
  {32'h4484e9d6, 32'hc2c548c8, 32'hc266f5d3},
  {32'hc4d27a1c, 32'h4406e304, 32'h42b6efe7},
  {32'h44237eca, 32'hbf8d5c8f, 32'hc33bf59f},
  {32'hc4d72ed4, 32'hc353b5e1, 32'h4316a7d4},
  {32'h44a2e205, 32'hc397eaf7, 32'hc1a30f1c},
  {32'hc4deca1c, 32'h4309b6b8, 32'h42303054},
  {32'h44e1e99c, 32'hc220f1f7, 32'hc3871865},
  {32'hc46718fc, 32'hc406b6b2, 32'hc296cce0},
  {32'h43f33620, 32'hc204a214, 32'hc209811a},
  {32'hc48c76ca, 32'hc31a0155, 32'hc3027f31},
  {32'h451e7a69, 32'hc36dc360, 32'h41ee456d},
  {32'hc3be9b90, 32'hc35f1ce5, 32'hc38d8d88},
  {32'h4513119f, 32'h434ea563, 32'h432d933e},
  {32'hc4ca8024, 32'h43606b4f, 32'h420562ce},
  {32'h42dbd130, 32'h427a9896, 32'h43b30ff9},
  {32'hc50c94de, 32'h42c51c6f, 32'hc3651819},
  {32'h450fcd4c, 32'h415b7e41, 32'h439320d9},
  {32'hc32e5350, 32'hc3296688, 32'hc3378501},
  {32'h43ec533e, 32'h4296033e, 32'h439856e8},
  {32'hc478ce14, 32'h44032883, 32'hc325db4f},
  {32'hc384d69c, 32'h4397ba4d, 32'hc233f265},
  {32'hc4e603b4, 32'hc26b6bde, 32'h430c53a0},
  {32'h44cf1f7b, 32'hc081a094, 32'hc2b9d5b0},
  {32'hc5327575, 32'hc31202f5, 32'hc2f73955},
  {32'h438aa3a6, 32'hc22335f1, 32'h411d6436},
  {32'hc4dc13bd, 32'h4388bd1d, 32'hc33cad28},
  {32'h448a3238, 32'h428708cf, 32'h42887d29},
  {32'hc4bbe275, 32'hc3ae503b, 32'h4378fd32},
  {32'h44439ff8, 32'hc33fb8ef, 32'hc322bbf0},
  {32'hc389c5e8, 32'hc2baaa19, 32'h43e4e3fc},
  {32'h444b1c67, 32'h43866f64, 32'h439439d1},
  {32'hc45a44d7, 32'h4118468f, 32'h42ab6b82},
  {32'h44a77390, 32'h425070ed, 32'hc2e69825},
  {32'hc49a1099, 32'h42bc0e48, 32'hc30fb5e0},
  {32'h44aec0fe, 32'h428b72a0, 32'hc2c5754e},
  {32'hc4753b2e, 32'h43190ad6, 32'h42a87d25},
  {32'h44b58cba, 32'h41a793be, 32'hc393a93d},
  {32'hc45953a6, 32'h4351d54e, 32'h43557605},
  {32'h4524339d, 32'h42c5706c, 32'hc273ccb9},
  {32'h4343d5b8, 32'h4316b0ac, 32'h42f9efbc},
  {32'h44a43868, 32'h42395b1f, 32'hc2bead6c},
  {32'hc50a7fdd, 32'hc1fb82d4, 32'h43e10e8c},
  {32'h43327420, 32'h42a101d7, 32'h43621e55},
  {32'hc519401c, 32'hc21b31f4, 32'h43232c48},
  {32'h444741ab, 32'h43598f2e, 32'hc38be34b},
  {32'hc4fac77e, 32'hc3848e75, 32'hc3ddfb9a},
  {32'h4411471e, 32'h43237bf7, 32'hc32cf186},
  {32'hc49f26ba, 32'hc3193292, 32'h440772cd},
  {32'h44fe8f48, 32'hc3c59f52, 32'h43bced35},
  {32'hc4a2d910, 32'hc3c01b28, 32'hc24203ab},
  {32'h44d861b2, 32'hc2b054cf, 32'hc396c9ba},
  {32'hc5046322, 32'h429051e5, 32'hc353bf59},
  {32'h44e465d7, 32'h42e0fa06, 32'hc2884580},
  {32'hc4881630, 32'h43f728b4, 32'h42e9de9e},
  {32'h448f87e6, 32'hc31f612c, 32'hc3716527},
  {32'hc3750230, 32'h4289b9e4, 32'hc299b82e},
  {32'h44fa2ff0, 32'h435ae4f0, 32'h4272487d},
  {32'hc49065a7, 32'hc2f9dac8, 32'h42ca6e13},
  {32'h43d76530, 32'hc2c8b491, 32'hc180a699},
  {32'hc2e5231f, 32'hc1b4cec3, 32'h43f49a34},
  {32'h44ee6d20, 32'hc22b859d, 32'hc37dfdb7},
  {32'hc21e7968, 32'h43c231ae, 32'h42d3508e},
  {32'h442c11d6, 32'h433354da, 32'hc23ef3f1},
  {32'hc3a897d0, 32'h4305efbe, 32'h421bef9f},
  {32'h44a49d46, 32'hc3710aaa, 32'hc2eb4efb},
  {32'hc50b574b, 32'hc33dd87a, 32'h42d2e0d6},
  {32'h44b07432, 32'hc32990ee, 32'hbfad4d46},
  {32'hc3e9d920, 32'h43445fc6, 32'h43899415},
  {32'h441753c2, 32'h43657c3e, 32'hc3a7c5e7},
  {32'hc4774d5a, 32'hc327c0c7, 32'h41c179f6},
  {32'h44427322, 32'hc2e4eede, 32'h421af93f},
  {32'hc4cd98a6, 32'h4323f9b2, 32'h4251548b},
  {32'h43180188, 32'hc30180cc, 32'hc366aa71},
  {32'hc44c50aa, 32'h43335232, 32'h43580e5f},
  {32'h44d4278f, 32'h418c3fc0, 32'hc1a1b92d},
  {32'hc4bf5ba1, 32'hc2cdab3c, 32'h429bbd8f},
  {32'h44f3952a, 32'hc1d945b2, 32'hc2844f39},
  {32'h44d4b8d5, 32'hc36b0038, 32'hc1bb50e9},
  {32'hc50f449a, 32'h41bc7799, 32'hc38e2a9d},
  {32'h44366d58, 32'h43f77ed6, 32'hc3861fd2},
  {32'hc3e74a5e, 32'hc0476c70, 32'h41f9c708},
  {32'h4398c374, 32'hc31e2f69, 32'hc34fb20d},
  {32'hc4c849dd, 32'hc2d1ac1c, 32'h428b33e6},
  {32'hc1f44200, 32'h4397577c, 32'hc1cac528},
  {32'h43102b28, 32'h4349a83b, 32'hc3e4b6b2},
  {32'h44e6b939, 32'hc1c2e430, 32'hc18c1c4c},
  {32'hc51cb6de, 32'h430522ad, 32'hc2d87911},
  {32'h44dea94e, 32'hc214a364, 32'h430a17aa},
  {32'hc47f52f0, 32'h42b88cfc, 32'h43ac4447},
  {32'h449c4774, 32'h422bdcf7, 32'hc31e2c8f},
  {32'hc38bab11, 32'hc2cac1e4, 32'h42731277},
  {32'h44b6088c, 32'h4338e76e, 32'hc376320e},
  {32'hc4d9c127, 32'hc210ce30, 32'hc3591840},
  {32'h44a9f40e, 32'hc3122d8e, 32'hc3d51178},
  {32'hc4942d00, 32'hc2d9e693, 32'h44038db9},
  {32'h44e43156, 32'hc20ec591, 32'h43003625},
  {32'hc4c3f903, 32'hc33777a3, 32'h432e254b},
  {32'h44c00115, 32'hc29c4698, 32'hc315c90a},
  {32'hc3993514, 32'h438a9a4d, 32'h42709d5a},
  {32'h44bde5f9, 32'hc3646102, 32'h41da165b},
  {32'hc32ba28a, 32'hc32149fe, 32'h431429ec},
  {32'h44dca37c, 32'hc36042fa, 32'h4195d5e5},
  {32'hc446b26e, 32'h433e2c4b, 32'h435b9ce3},
  {32'h44864976, 32'hc2abcba0, 32'hc3b11983},
  {32'hc51ed1d6, 32'hc428c431, 32'hc38683e6},
  {32'h44a295a9, 32'h4352103b, 32'h428d7498},
  {32'hc48bc068, 32'h430005bc, 32'h40cd40dc},
  {32'h443d5c36, 32'hc368124c, 32'h4380b98e},
  {32'hc44bde15, 32'hc0c65a1c, 32'hc30c9de7},
  {32'h447a2e4f, 32'h42e9c481, 32'hc306571f},
  {32'hc4270249, 32'hc3cd4f3a, 32'h43929a96},
  {32'h449eb078, 32'h4395c187, 32'hc2bdc85e},
  {32'hc4e7e90d, 32'hc31c47cf, 32'h428cb0cb},
  {32'hc2eab958, 32'hc362f99d, 32'hc3688c55},
  {32'hc51856e3, 32'hc3678a7f, 32'h4350e20e},
  {32'h45106ce2, 32'h43be1a98, 32'hc2b24c0c},
  {32'hc4d9f4fa, 32'h41cc6023, 32'hc3bc3683},
  {32'h4501dfdb, 32'h43a599a3, 32'hc32c7a7c},
  {32'hc4c539e1, 32'h425c2399, 32'hc33145cd},
  {32'h444e0f88, 32'hc3f68f86, 32'h4381f638},
  {32'hc3cb823d, 32'hc2753cbd, 32'hc34f90a9},
  {32'h4524c263, 32'h4369ca28, 32'hc3475b64},
  {32'hc4b066ce, 32'h4265dce2, 32'hc3222755},
  {32'h44a5c0ef, 32'hc310800b, 32'h43bc6d41},
  {32'hc3c2ca90, 32'hc31c9caa, 32'h4367b9ba},
  {32'h4519b13c, 32'h42bb4ac4, 32'h428d34dd},
  {32'hc4318e04, 32'hc361b627, 32'hc2a49b1d},
  {32'h45104e2d, 32'hc294daa3, 32'h4214a909},
  {32'hc4409b4b, 32'h42d9f90e, 32'hc3085dcb},
  {32'h4406550c, 32'hc21cdd40, 32'hc306595b},
  {32'hc50bfb79, 32'h437937cd, 32'hc2bf3e74},
  {32'h44fb8ae3, 32'h42ef2a86, 32'hc3084293},
  {32'hc45f5336, 32'hc1fcbb96, 32'hc3510c67},
  {32'h44d98501, 32'h4360d3fd, 32'hc30531be},
  {32'hc4caacb9, 32'hc2c13dc6, 32'hc19a902e},
  {32'h44921955, 32'hc2bc6d77, 32'h436fe337},
  {32'h434f27a0, 32'hc33a3cdc, 32'h4386a179},
  {32'h443a1e90, 32'h42cedaed, 32'h430903d9},
  {32'hc50abfe9, 32'hc309fe48, 32'hc336888d},
  {32'h447a4d32, 32'h432e2788, 32'h43c908da},
  {32'hc4e424a0, 32'hc191e5f8, 32'h4404e129},
  {32'h45153449, 32'h431313d2, 32'hc35753a2},
  {32'hc3ce2ab8, 32'hc2faf760, 32'h43d12bb9},
  {32'h44bdd242, 32'h43ec8c12, 32'h43cb8a13},
  {32'hc38cb5bd, 32'h42782d42, 32'hc29a8533},
  {32'h44c5d24a, 32'hc2825247, 32'h431d54cd},
  {32'hc4adf1ce, 32'h435d6814, 32'h42c62f1a},
  {32'h44876112, 32'h42409f4b, 32'h4223e090},
  {32'hc488468d, 32'hc3d1aa51, 32'hc254f3f0},
  {32'h44310ab4, 32'h440375f0, 32'hc27beaba},
  {32'hc48095d7, 32'h437a450b, 32'h435bd1df},
  {32'h44bf60b4, 32'hc2409df1, 32'h432c689e},
  {32'hc5049812, 32'hc2790bc8, 32'hc3337477},
  {32'h44fd7e4f, 32'hc39e41a2, 32'hc2fdf603},
  {32'hc49ec5c2, 32'hc3853038, 32'hc3cbe202},
  {32'h4517d69a, 32'hc36cf190, 32'h43cd7569},
  {32'hc5000b76, 32'hc39ecc43, 32'hc39465fd},
  {32'h44c1c096, 32'h429c97a1, 32'hc2e34090},
  {32'hc5056fc3, 32'hc298b219, 32'hc35546a3},
  {32'h4533ac57, 32'hc1af67c1, 32'hc27dec43},
  {32'hc21b4300, 32'h429ba393, 32'hc362cbeb},
  {32'h449d7026, 32'hc392e9f2, 32'hc33e3ff0},
  {32'hc44dadf0, 32'hc29d0b9b, 32'hc303229c},
  {32'h43775182, 32'h4324faa8, 32'hc3c2c036},
  {32'hc3c8832f, 32'hc38f0906, 32'hc1dcec53},
  {32'h44d37a08, 32'h43999b7e, 32'h42275bb9},
  {32'hc4c2bf2c, 32'h43b6fd36, 32'h423dcedf},
  {32'h44467ef0, 32'hc3a5f39c, 32'hc3bd62bf},
  {32'hc44e1ed2, 32'h42f842e6, 32'h43c3385c},
  {32'h446c0cd7, 32'h4336e155, 32'hc2e1ce1c},
  {32'hc4da8084, 32'h435a89e5, 32'h429fe3c8},
  {32'h45062ca6, 32'h430a2b40, 32'hc378e103},
  {32'hc47d6a52, 32'hc2d0c416, 32'h43e0ae0b},
  {32'h439cfe30, 32'h4257e55e, 32'h442b1f90},
  {32'hc4fc39da, 32'h43d76498, 32'h43ae8a9f},
  {32'h4487e156, 32'h43daefd8, 32'hc386f63c},
  {32'hc49b36c7, 32'h42d64a22, 32'hc2b97a18},
  {32'h44f21964, 32'h43a3e7f0, 32'h431039d0},
  {32'hc4c0a80a, 32'hc36d95fe, 32'hc3c00ed4},
  {32'h4482d65c, 32'h43599c00, 32'hc32018cd},
  {32'hc3d728d8, 32'h4380d4cf, 32'h4325afc7},
  {32'h4454db7c, 32'hc2fb620c, 32'h433e5b57},
  {32'hc47384ff, 32'hc3a57d36, 32'h43d311d9},
  {32'h448ed865, 32'h4333cced, 32'hc3c8b576},
  {32'hc4214bb8, 32'hc3e1eb4b, 32'h43c139bd},
  {32'h451d02ff, 32'hc1b602e0, 32'hc25e5193},
  {32'hc4a3a532, 32'hc1862be9, 32'hc1d5726c},
  {32'h44cbb8f9, 32'hc322cca2, 32'hc3b779c8},
  {32'hc4893928, 32'h403de36a, 32'h43a99160},
  {32'h44005ad3, 32'h429725f8, 32'h42a4caff},
  {32'hc41ee304, 32'h43f1717b, 32'h42c8afca},
  {32'h45084351, 32'hc2873d88, 32'h42b1a992},
  {32'hc4d2e5a3, 32'h42a3f5b9, 32'h42a9eb40},
  {32'h43ef5de6, 32'hc368ab2e, 32'hc375868d},
  {32'hc4f1f480, 32'h42c009ba, 32'h430d6b45},
  {32'h450ee027, 32'h40d34e04, 32'hc2ecc23c},
  {32'hc3d91960, 32'h41bc1c71, 32'h439ab9f5},
  {32'h4457e3aa, 32'hc2cc64e9, 32'h4386d525},
  {32'hc45b771c, 32'hc3233249, 32'h4316ad85},
  {32'h4511627a, 32'h439d71cb, 32'h431efce2},
  {32'hc435deb7, 32'hc306ad89, 32'hc10b9509},
  {32'h435a2e90, 32'hc2a4310e, 32'h41c98d28},
  {32'hc49d0f47, 32'hc2ada43c, 32'h43279c43},
  {32'h444ab58e, 32'h42b1abc7, 32'hc383eb05},
  {32'hc5045859, 32'h41c6884a, 32'h42abe00a},
  {32'h4408726e, 32'hc14b2830, 32'hc350d839},
  {32'hc48128e7, 32'h438a5613, 32'h4331e4d4},
  {32'h441c4761, 32'hc402526a, 32'hc319e0f8},
  {32'hc4ec70bc, 32'hc431cd78, 32'h430d80b9},
  {32'h43112717, 32'hc3aae37b, 32'hc2bc57cb},
  {32'hc4a39d56, 32'h42528c5e, 32'hc12cc4e6},
  {32'h450df0a7, 32'h41ce7512, 32'hc382b6b5},
  {32'hc4dff3b1, 32'hc2c902f6, 32'hc324d2dc},
  {32'h43a170d1, 32'h430acab1, 32'h42b1d3e4},
  {32'hc48492e0, 32'hc292a5c6, 32'hc33c22e6},
  {32'h44062da8, 32'h436a38da, 32'hc3a25abf},
  {32'hc4170f42, 32'h41c30fe5, 32'h435c4128},
  {32'h4510a60c, 32'h43131c01, 32'hc3cca15b},
  {32'hc2842da0, 32'hc35c6b0d, 32'h4367a312},
  {32'h450816a9, 32'h432d0147, 32'hc20bf15f},
  {32'hc49db789, 32'hc3ae9d76, 32'hc2f02a5c},
  {32'h44395aee, 32'h439b6d90, 32'hc36f9977},
  {32'hc44e0f50, 32'h42c91c04, 32'hc346a887},
  {32'h43e6690f, 32'hc40301ed, 32'hc3234a81},
  {32'hc3c549c1, 32'hc309b9ca, 32'hc394fd04},
  {32'h448e7d42, 32'h4234613e, 32'hc29a1cb3},
  {32'hc4d2378e, 32'hc34daebb, 32'h439123f1},
  {32'h438f6a00, 32'h434430b1, 32'hc3a15692},
  {32'hc4fc300d, 32'hc395350c, 32'h42662294},
  {32'h43eeb6ce, 32'hc362adf1, 32'h423d1bc2},
  {32'hc4e6140f, 32'h42bf63ac, 32'h43bca078},
  {32'h44af2cb6, 32'hc2c6ad75, 32'h439284fc},
  {32'hc2886f70, 32'hc374bb10, 32'hc31a5364},
  {32'h448fba9f, 32'hc3409ba3, 32'h42a8e3a3},
  {32'hc436e376, 32'hc366d2b6, 32'hc3a612ee},
  {32'h44dffe28, 32'hc34944c3, 32'hc285fc12},
  {32'hc501d86e, 32'hc3e7b7fc, 32'h420d6252},
  {32'h442dfce8, 32'hc34c1930, 32'h43c62aee},
  {32'hc4b8e171, 32'hc2eea9da, 32'hc28488dd},
  {32'h44e243d4, 32'h423c726e, 32'h43a941f2},
  {32'hc3c21d72, 32'h42692698, 32'hc2c56c08},
  {32'h44d57c6b, 32'h439d5d24, 32'h42eb0fe2},
  {32'hc4af61ae, 32'hc3c73e3b, 32'h43b4d1ea},
  {32'h43facf40, 32'hc384df7c, 32'hc2a7f145},
  {32'hc3e5a7aa, 32'h43f56e92, 32'hc36addc7},
  {32'h44bddbab, 32'hc33fc5ba, 32'hc250bbd5},
  {32'hc4994c2b, 32'h4404c4b1, 32'h400ad8d0},
  {32'h4499f966, 32'h438327e6, 32'hc399ab42},
  {32'hc4951e66, 32'hc39762d2, 32'h438a96d4},
  {32'h4505e84b, 32'hc3e4230e, 32'hc3e50ed2},
  {32'h432512c0, 32'h43c0a872, 32'hc3b3a206},
  {32'h450800be, 32'hc3673abf, 32'h4336e442},
  {32'hc479ec59, 32'h43b279e1, 32'hc368e428},
  {32'h445bacec, 32'h430b6a70, 32'h4330dbcd},
  {32'hc4a6493c, 32'h436fe74b, 32'hc38bcbd8},
  {32'h4438d584, 32'h437bd5d5, 32'h43ab614d},
  {32'hc4872294, 32'h41e27a31, 32'hc314d406},
  {32'h44c73401, 32'h41c8fe32, 32'h41e6fded},
  {32'h43056ac8, 32'h43a4ce79, 32'hc3186b36},
  {32'h44d5f5e5, 32'h43861bcc, 32'h43241f96},
  {32'hc47cbfd8, 32'hc383fecf, 32'h4320a0a1},
  {32'h44833aac, 32'hc3821e73, 32'h423d8705},
  {32'hc3a4c2f7, 32'h4237c7b8, 32'h422f17b4},
  {32'h44d277b9, 32'h4240dca7, 32'hc313bad3},
  {32'hc4364ff8, 32'hc3427d52, 32'h4299d8be},
  {32'h43c2155e, 32'hc311bdfb, 32'hc277a4ac},
  {32'hc4e870af, 32'h432d0642, 32'h4370780a},
  {32'h45172352, 32'hc34520a8, 32'h42c93e78},
  {32'hc4f53e53, 32'hc3b33f1a, 32'hc36aa3c9},
  {32'h44bc4b26, 32'h41e43502, 32'hc304f29f},
  {32'hc4cf9a10, 32'hc303c39a, 32'hc307466d},
  {32'h44a63ea3, 32'hc35de676, 32'hc2f6833b},
  {32'hc429ebdc, 32'h434ba1d0, 32'hc2f01ed7},
  {32'h44c61e16, 32'hc2cddcf2, 32'hc3a23531},
  {32'hc3ec3db5, 32'hc381bf15, 32'h42eeaaad},
  {32'h45058b85, 32'h430bafe1, 32'hc3275d69},
  {32'hc4c1ec92, 32'h42f88c5c, 32'h42aaafae},
  {32'h44b8ab3a, 32'hc219ff61, 32'h43cb988a},
  {32'hc44da006, 32'h3d913280, 32'h429cc612},
  {32'h44ed28f0, 32'h432338f2, 32'h4317d138},
  {32'hc49f58ba, 32'hc3086035, 32'h42c90f71},
  {32'h44c89213, 32'hc4084d23, 32'h41a3c431},
  {32'hc49a4e2f, 32'hc3261b12, 32'hc2c9b1ed},
  {32'h447dce67, 32'h43d6c7f1, 32'hc38826fe},
  {32'hc4eb3946, 32'hc3cabcf5, 32'h430d0493},
  {32'h42b01ed0, 32'hc26a6afc, 32'hc2feb47b},
  {32'hc40ecff6, 32'h4043eb80, 32'hc38ca005},
  {32'h432de870, 32'hc2b43bad, 32'h43843279},
  {32'hc4dbc909, 32'hc084eaed, 32'h429c248c},
  {32'h44922354, 32'h42540fd3, 32'hc34e70a9},
  {32'hc49b695e, 32'h4274df15, 32'hc31f8ebb},
  {32'h4510403e, 32'hc0fba5ed, 32'hc38cb759},
  {32'h43c2b108, 32'hc3ca5ebb, 32'hc30b3196},
  {32'h440e60ae, 32'hc30b8421, 32'hc3b5009c},
  {32'hc413f2ef, 32'h43431830, 32'h4380ff6f},
  {32'h44ebc68b, 32'hc2f48691, 32'h4148c167},
  {32'hc447190e, 32'hc2899075, 32'h41e6535e},
  {32'h447e1d4a, 32'h43af1d90, 32'h43b49f30},
  {32'hc44292b3, 32'h43af651a, 32'h4331ffff},
  {32'h42d093e8, 32'h43295ee1, 32'h439d7e55},
  {32'hc50c0a05, 32'hc1cf4c78, 32'hc3e3795e},
  {32'h450c0cac, 32'hc363e55b, 32'h42adc647},
  {32'hc4f4b9eb, 32'h43acdbf7, 32'h43ba0a6d},
  {32'h443e5342, 32'h43afea91, 32'hc38cdd56},
  {32'hc44c8bf2, 32'h4401ba7b, 32'h4211dacd},
  {32'h4469d623, 32'h4262e707, 32'hc36e8f42},
  {32'hc4da0aed, 32'h4430f29e, 32'h42c3d170},
  {32'h44eb1c8a, 32'h43488400, 32'h42053c98},
  {32'hc4adeb5e, 32'h42ed0602, 32'hc3852172},
  {32'h45188764, 32'hc3cf9458, 32'h432f0bf2},
  {32'hc44e2098, 32'h422ef93a, 32'hc20f8b82},
  {32'h44f00bda, 32'h40c97da4, 32'hc295f337},
  {32'hc4ae61c7, 32'h4381f2f4, 32'hc24259b4},
  {32'h4507eecd, 32'h4388b36e, 32'hc30ada0a},
  {32'hc44459c5, 32'hc30d25c4, 32'h42f6fe96},
  {32'h44c79158, 32'h4391c0f8, 32'h43b71ca1},
  {32'hc440f15e, 32'hc3570335, 32'hc262634b},
  {32'h449596be, 32'hc15c2b82, 32'hc3be4b76},
  {32'hc3e964de, 32'h43249bde, 32'hc3801439},
  {32'h450821ec, 32'hc3801f23, 32'h42ff1127},
  {32'h42978760, 32'hc33172c5, 32'h435e8a78},
  {32'h44a4a043, 32'hc3374ce1, 32'hc1d03673},
  {32'hc2db4f60, 32'hc3da9275, 32'h42926214},
  {32'h44a41d8e, 32'h433a8797, 32'hc38ca56f},
  {32'hc4af32cb, 32'h427afe82, 32'hc331a68e},
  {32'h44c48454, 32'hc34fb5b6, 32'h43685ac9},
  {32'hc4ec347a, 32'h43098e41, 32'hc37fa8c0},
  {32'h44324670, 32'h42bfb0fc, 32'hc23c3b43},
  {32'hc3dd62b0, 32'h42c2300d, 32'hc2d4132c},
  {32'h43e29f54, 32'hc2f2d6e8, 32'hc29dedbf},
  {32'hc3246cf6, 32'h43885350, 32'h419d301e},
  {32'h44fba286, 32'h4315fa47, 32'h426da92b},
  {32'hc43975fc, 32'hc313e811, 32'hc38d2f2b},
  {32'h44f77e45, 32'hc3db0e93, 32'h432bb5b3},
  {32'hc42eb084, 32'h431294e0, 32'hc3067163},
  {32'hc1ab6eea, 32'hc41755c1, 32'hc31dd8f0},
  {32'hc4c3a92d, 32'h428b3ff2, 32'h428aadc1},
  {32'h44175d98, 32'hc3d518a7, 32'hc257481b},
  {32'hc4f05e70, 32'h4381e221, 32'h4367f0df},
  {32'h442099c1, 32'hc38969a4, 32'h431b800c},
  {32'hc4f65df6, 32'hc39202b1, 32'h43e418b1},
  {32'h45039443, 32'h40b803aa, 32'hc2f0d13f},
  {32'hc4c66200, 32'hc288f41a, 32'hc3339a6a},
  {32'hc29fde2c, 32'h4302bcb1, 32'hc33e401a},
  {32'hc359ec60, 32'hc39eb3a6, 32'h42fe16ab},
  {32'h44450769, 32'h4225c484, 32'hc3883460},
  {32'hc489ef82, 32'hc36b8199, 32'hc2cc21d2},
  {32'h44b6230d, 32'hc33187ee, 32'h41ab3bbb},
  {32'hc5045b87, 32'hc28a8687, 32'hc29f18bd},
  {32'h450365a1, 32'h42e233be, 32'hc40f02a1},
  {32'hc50576b4, 32'hc2654fd0, 32'hc19d8f64},
  {32'h4488e3b3, 32'h432cb6c2, 32'hc3097907},
  {32'hc4ac296e, 32'hc3ab1188, 32'h43c0a193},
  {32'h450ac58a, 32'h439b4278, 32'h42093ff8},
  {32'hc4358e6e, 32'h43b4ccb3, 32'hc2a236a5},
  {32'h44f3e705, 32'hc388ddf8, 32'h43209014},
  {32'hc4a14027, 32'h4327c0cc, 32'h4322f7a3},
  {32'h43af882b, 32'hc351bd6a, 32'hc319c700},
  {32'hc4ea3982, 32'hc1b65c58, 32'h418bf261},
  {32'h44efdc08, 32'h4221bcff, 32'h40b3996b},
  {32'hc480dcb6, 32'hc39a0c37, 32'hc1f9734d},
  {32'h450cd8f0, 32'hc32c6bbd, 32'h43b4d1df},
  {32'hc4bc029c, 32'hc32196f3, 32'hc217d76c},
  {32'h44242cbc, 32'hc2885a6a, 32'h429627f7},
  {32'hc4930043, 32'h4334f0c4, 32'h4290952d},
  {32'h4499963a, 32'hc301d31d, 32'h43a2f2c3},
  {32'hc51d2a3e, 32'hc3377173, 32'h4253a0e9},
  {32'h4498a13a, 32'hc32b1be9, 32'h427b8a99},
  {32'hc4ff4073, 32'hc3c8e9a8, 32'h43813ba7},
  {32'h447ba023, 32'hc0938ae2, 32'hc31bb9c3},
  {32'hc4d90876, 32'h424cd38e, 32'h425aa85c},
  {32'h44bd82ee, 32'h430a4efa, 32'hc3aeaef3},
  {32'hc490c1e0, 32'h438527bd, 32'hc3473ee1},
  {32'h43d9dc2c, 32'hc20fea0e, 32'h439b9331},
  {32'hc45815e5, 32'h41f266e8, 32'h43859bcf},
  {32'h442dd2fc, 32'h4317ac4d, 32'h40834eac},
  {32'hc4e3beb2, 32'h42611692, 32'h435cc437},
  {32'h437278d0, 32'h4325e3aa, 32'hc337bbb3},
  {32'hc5124d07, 32'hc2edf5e1, 32'hc36dd4c1},
  {32'h43cd4786, 32'h4097a4e7, 32'h42abf17f},
  {32'hc4dddca0, 32'hc38f6ac3, 32'h42c6f9ef},
  {32'h4507ab87, 32'hbfa295a8, 32'hc3a74aa3},
  {32'hc3cd8bf8, 32'hc196b82c, 32'h42a2b5c0},
  {32'h451a3242, 32'h437dfdad, 32'h438fba68},
  {32'hc44d63dc, 32'hc3d4fd57, 32'h43a24857},
  {32'h45107f63, 32'h4390798c, 32'h43e9d121},
  {32'hc4415d89, 32'h4337d10c, 32'h43661d84},
  {32'h44a2e523, 32'hc20ae1ad, 32'hc3921dfe},
  {32'hc4d827e2, 32'hc2b8ba40, 32'h421e9978},
  {32'h4503c42e, 32'h433d1b63, 32'h43b59ed1},
  {32'hc5039ae4, 32'hc287fb58, 32'hc39ebce2},
  {32'h441acd4b, 32'h43843447, 32'hc3869b00},
  {32'hc5088844, 32'h43a9fce5, 32'hc3a465d5},
  {32'h44ecb8da, 32'hc298067d, 32'h43887b33},
  {32'hc4f33353, 32'hc2902f88, 32'h41b2a252},
  {32'h44fe3620, 32'h4338887c, 32'hc33b29dc},
  {32'hc4a53382, 32'hc2d3f9ad, 32'hc3c29f05},
  {32'h44ba58c1, 32'hc377ab73, 32'hc3b753a6},
  {32'hc3f66bac, 32'h432f91c2, 32'hc270c120},
  {32'h4496a7cd, 32'h42d8dbd5, 32'h4374bb1f},
  {32'hc45874ab, 32'hc304d4a0, 32'h41af66d2},
  {32'h41f6d9d1, 32'hc2a93305, 32'hc3ab2780},
  {32'hc4f62c22, 32'hc29165ca, 32'hc3e26f67},
  {32'h447663a8, 32'hc35ca6a8, 32'h429b659c},
  {32'hc446e3dd, 32'h425894e0, 32'h422442a1},
  {32'h4468fbc3, 32'h43825e9a, 32'hc2f4b3d0},
  {32'hc513c29f, 32'h406e28e0, 32'h4374ddef},
  {32'h431c12a4, 32'hc3012ab2, 32'h423e2f67},
  {32'hc485c93e, 32'hc3a37a38, 32'hc33342a1},
  {32'h44d49168, 32'h41b548b3, 32'hc36340a0},
  {32'hc4717024, 32'hc324168f, 32'h411b4244},
  {32'h4514ecb4, 32'hc2491dd4, 32'hc35698f7},
  {32'hc46a92c0, 32'hc240df75, 32'hc38a51c8},
  {32'h43c6f148, 32'hc2d50765, 32'h42395216},
  {32'hc38c3d14, 32'hc2dccbe4, 32'h42afba55},
  {32'h448ee7ca, 32'hc3b0060b, 32'h43033eb6},
  {32'hc5138ce4, 32'h42eed16d, 32'h43ce80cc},
  {32'h44e37c29, 32'h43243d3e, 32'hc2e6be21},
  {32'hc48f4b72, 32'hc3b18bee, 32'hc395ddda},
  {32'h433f4a7c, 32'hc28d1d6b, 32'hc22011d7},
  {32'hc3abca28, 32'h431552d1, 32'hc386edf1},
  {32'h450c3e05, 32'h43017832, 32'h4303c6af},
  {32'hc50f3234, 32'h41b164ee, 32'hc39d808b},
  {32'h44b94f36, 32'hc37b83af, 32'h4483eb94},
  {32'hc457ad43, 32'hc2dc1e23, 32'h43259f0e},
  {32'h43ab0a75, 32'h438b5d91, 32'h413c94b0},
  {32'hc4f17662, 32'h431eb8be, 32'h436f4d7b},
  {32'h44e4c6d1, 32'hc2620c48, 32'hc3133e89},
  {32'hc48a05fe, 32'h429e28b8, 32'h431d9bc4},
  {32'h44a8b56f, 32'hc27f8391, 32'hc269c175},
  {32'hc515543e, 32'hc3a04ebc, 32'h42c9de54},
  {32'h44d4f8e2, 32'h42f58a3f, 32'h42294761},
  {32'hc3c6b3bc, 32'h425ede51, 32'hc30f5b84},
  {32'h43320908, 32'h4401cb73, 32'h432ebef8},
  {32'hc351cdea, 32'hc295a7f3, 32'h42246aae},
  {32'h44cc79af, 32'h431cec97, 32'h43262b95},
  {32'hc43b8c38, 32'hc34c26f1, 32'h42fa2e25},
  {32'h449d0864, 32'hc30c79ef, 32'h43ad93a9},
  {32'hc5057f54, 32'h43bb2231, 32'h43b0fffb},
  {32'h4397dcf8, 32'h4352f037, 32'hc2b263ef},
  {32'hc3b4ccb9, 32'hc1e3045a, 32'h432501f1},
  {32'h452a1479, 32'hc1e1da3b, 32'hc31240cc},
  {32'hc2bcd0d2, 32'hc2e700f1, 32'h430eb7ab},
  {32'h43c6c398, 32'hc3fa6399, 32'hc2d4348c},
  {32'hc4cb2fb2, 32'hc3e50135, 32'h4336babe},
  {32'h4431b2ca, 32'hc14a7229, 32'h439ab8b3},
  {32'hc47a525b, 32'hc3a49a1a, 32'h42ec9fa1},
  {32'h44170de9, 32'h421f3651, 32'hc3514b11},
  {32'hc4d3f1e4, 32'hc2d8435e, 32'hc3764f40},
  {32'h4460502d, 32'h42abedbe, 32'hbf836018},
  {32'hc4ea0e58, 32'hc2c3cdad, 32'hc30c07b0},
  {32'h42dd2580, 32'hc2a74ed5, 32'h43231bb5},
  {32'hc518370d, 32'h43d3815e, 32'hc2260308},
  {32'h44d8137e, 32'h439dc74e, 32'hc3476a5f},
  {32'hc4f018b3, 32'h439d2a57, 32'hc36d7e95},
  {32'h450e5cdf, 32'h43b81a6b, 32'h428b6c7b},
  {32'hc3ca0f88, 32'h437918f1, 32'h413db43e},
  {32'h435498c0, 32'h43c20ff3, 32'h42f88d5e},
  {32'hc33d8f90, 32'h43163f2b, 32'hc1e0d7a5},
  {32'h44d65445, 32'hc187dfd9, 32'h43cbe8e2},
  {32'hc50a22ca, 32'h43d58d1b, 32'h429328e0},
  {32'h4450a5db, 32'hc0da7bfa, 32'h43a88295},
  {32'hc440b59d, 32'hc3899a66, 32'h4342c73e},
  {32'h446a76a0, 32'h43356c74, 32'hc3ba083d},
  {32'hc4ebac80, 32'h42609967, 32'h425ed64d},
  {32'h45383e67, 32'h4311fbe4, 32'h4214250b},
  {32'hc501080b, 32'h42bf1d83, 32'h43df8361},
  {32'h450f4d5d, 32'hc32f1568, 32'h43b705d1},
  {32'hc46f4210, 32'hc387c5ef, 32'h43065c4a},
  {32'h43bdc618, 32'hc1bb622c, 32'hc3a3cca3},
  {32'hc517ee30, 32'h42cb128e, 32'h4383edf0},
  {32'h448f4c8f, 32'hc1e34593, 32'h438b9c8d},
  {32'hc4d364e4, 32'hc3587793, 32'hc3f86c46},
  {32'h4423ea5f, 32'hc34bbec0, 32'h43b5520b},
  {32'hc402440d, 32'hc29a1132, 32'hc2f7c884},
  {32'h45047b11, 32'h422769fa, 32'hc31a1495},
  {32'hc4f82759, 32'h42c7e9e2, 32'hc348d561},
  {32'h444ff064, 32'hc2a922c7, 32'h43f16a7d},
  {32'hc3a60741, 32'hc363f274, 32'hc3d280c9},
  {32'h44c61383, 32'hc3c5051b, 32'h441110d3},
  {32'hc27d4f00, 32'hc4036417, 32'h432ba960},
  {32'h450b2c3b, 32'hc3283cc0, 32'h425ee398},
  {32'hc4f1e685, 32'hc2002d24, 32'hc29dd932},
  {32'h44242cbe, 32'hc31e0c52, 32'hc3c0c16f},
  {32'hc482ff0e, 32'hc383d652, 32'h4094c22a},
  {32'h44d7994b, 32'hc2678179, 32'h43d8e244},
  {32'hc4131eb9, 32'hc24e9f77, 32'h420045b0},
  {32'h44380b85, 32'hc3a93b74, 32'h437ac3d9},
  {32'hc50dc4d2, 32'h3eb64464, 32'hc350bd7b},
  {32'h44953c84, 32'hc2e491af, 32'h434122fc},
  {32'hc06e0d10, 32'hc12650c6, 32'hc3a5209f},
  {32'h439ad96c, 32'h4082e646, 32'h43dd7c7f},
  {32'hc4bb3b76, 32'hc2b99132, 32'h420c3945},
  {32'h44ec8e81, 32'h41e328b7, 32'h43640db5},
  {32'hc3887410, 32'hc29cdd85, 32'hc357a965},
  {32'h43b7b4f9, 32'h41affcc5, 32'h430ab7d7},
  {32'hc4ec6e82, 32'hc303aa38, 32'h429928da},
  {32'h42f90990, 32'h411e008e, 32'hc2be1107},
  {32'hc5000aaf, 32'hc32d0ee6, 32'h439211a4},
  {32'h44deb2d5, 32'hc331889b, 32'hc3170bf9},
  {32'hc2487ae8, 32'hc2a2e8ea, 32'hc3acddd2},
  {32'h45102397, 32'h42b9c20a, 32'h43006dae},
  {32'hc4f9660e, 32'h434f8a3e, 32'h42c183be},
  {32'h45041e2c, 32'hc28bf9b2, 32'hc31b1cf7},
  {32'hc41ec2a2, 32'h415ed57a, 32'hc329a4bf},
  {32'h4413b163, 32'h3fbadc44, 32'h423bd178},
  {32'hc4b92b74, 32'hc3a69942, 32'h440845bb},
  {32'h4463b682, 32'h436560b2, 32'hc335a4db},
  {32'hc4ea7018, 32'hc29f7316, 32'h41960384},
  {32'hc2c245dc, 32'hc320b4e8, 32'h43680758},
  {32'h441065e6, 32'hc332f3ee, 32'h42ad93e6},
  {32'hc4358378, 32'hc41697d4, 32'hc2feb12b},
  {32'h4489f3dd, 32'h433ffb9b, 32'h42990a6c},
  {32'hc3dc9e22, 32'hc3824b86, 32'hc182fbd9},
  {32'h44a09afe, 32'hc3fa41f8, 32'h43f0d2f3},
  {32'hc4301a22, 32'hc2d51ce4, 32'h438ee613},
  {32'h4477f4d8, 32'h42af8a31, 32'h41612703},
  {32'hc384df4a, 32'h425f0899, 32'h420108ba},
  {32'h45088676, 32'h4394395d, 32'h43615559},
  {32'hc483415d, 32'h42d92652, 32'h41adf941},
  {32'h44de1a74, 32'h42c753f9, 32'h4348d5f8},
  {32'hc4dae7ce, 32'h41f1ff1e, 32'hc2b9683c},
  {32'h44c37140, 32'hc275cc56, 32'h43976689},
  {32'hc503d077, 32'h4326d048, 32'hc377a008},
  {32'h44ccf8f4, 32'h43272706, 32'hc2b64eca},
  {32'hc4ff0179, 32'hc279e61a, 32'h43a5f4dc},
  {32'h44e07c79, 32'h4280bbc6, 32'h42e7fa9f},
  {32'hc4861ad1, 32'h4280c954, 32'hc1ef90f0},
  {32'h449a1119, 32'h438d67bc, 32'h440470b0},
  {32'h42b222cb, 32'hc2452f44, 32'hc343268c},
  {32'h4455dbf5, 32'hc29d4444, 32'hc2ce988f},
  {32'hc4b590f4, 32'hc35fffc6, 32'h431f3a50},
  {32'h44df8ecc, 32'h433a2471, 32'h4310c860},
  {32'hc4ad0975, 32'h41c8ba15, 32'hc2cbd1e0},
  {32'h4303a490, 32'hc39f53af, 32'h42d07dc2},
  {32'hc50f1723, 32'hc1d7fa47, 32'h3fb3c2d2},
  {32'h45224eb3, 32'h42aa281f, 32'h435fc285},
  {32'hc4f4326a, 32'hc1a268d6, 32'h42a30f5d},
  {32'h44e757bb, 32'h434e3426, 32'hc2b50c8f},
  {32'hc38d6822, 32'hc384c998, 32'hc2ab55b3},
  {32'h44de3bb3, 32'hc1c0f52c, 32'h442ff185},
  {32'hc445d70a, 32'hc3699bf2, 32'hc391a5f4},
  {32'h449d4dc7, 32'hc336695f, 32'hc1fcf874},
  {32'hc5066b7b, 32'h4222aab8, 32'h4393736f},
  {32'h446aba8c, 32'h4203773d, 32'hc3252136},
  {32'hc44fcf00, 32'hc350ec6c, 32'hc37d14a7},
  {32'h44bbd998, 32'hc1de9e73, 32'h429151c1},
  {32'hc42866f8, 32'h4186ddae, 32'h439be96a},
  {32'h428fc830, 32'hc1e8a12c, 32'hc2b1c29e},
  {32'hc4d742b0, 32'hc307eeee, 32'h43223946},
  {32'h44c79c66, 32'h42a82615, 32'h430c78ce},
  {32'hc49bc1a8, 32'h418ef73d, 32'h43057742},
  {32'h44cec19e, 32'hc2bf43b1, 32'hc2b199bd},
  {32'hc4a2cd9c, 32'h42f37108, 32'hc34991c9},
  {32'h434f6a00, 32'h41f14543, 32'h42f5ffe5},
  {32'hc412a0d4, 32'h426af2da, 32'hc355b4ee},
  {32'h44b3f58e, 32'hc297359b, 32'h43789db5},
  {32'hc40b1d8a, 32'h43dcee97, 32'hc35dae76},
  {32'h43e7ba5c, 32'h43111af4, 32'hc3f17bdc},
  {32'hc4cf84aa, 32'hc2575703, 32'h432f97a4},
  {32'h43cd1298, 32'h41b4451e, 32'h433f283c},
  {32'hc46eea19, 32'h43752a53, 32'hc32fb960},
  {32'h436cff3e, 32'hc3c2b19b, 32'h428ed580},
  {32'hc501824f, 32'hc1a8f178, 32'hc2c0fa9e},
  {32'h43d047b8, 32'h43c86c80, 32'hc2d05200},
  {32'hc4b6cdf8, 32'hc2232a39, 32'h42940cd6},
  {32'h444f2f87, 32'hc3b89261, 32'hc32cf380},
  {32'hc4b48cac, 32'h435ca678, 32'hc32d7528},
  {32'h4506461f, 32'hc3ef00e1, 32'h43eefd6c},
  {32'hc469da10, 32'hc40d6157, 32'h4186a9b9},
  {32'h447de1f6, 32'h43b5b937, 32'h434e19fc},
  {32'hc3c51151, 32'h4342acc9, 32'h41b2ed65},
  {32'h44656ff3, 32'hc3a99dfa, 32'hc359810e},
  {32'hc51b8caa, 32'h437c4d42, 32'hc371b129},
  {32'h44a6aba4, 32'h40bb0ddd, 32'h4311bebf},
  {32'hc506e96d, 32'hc2e8bf7b, 32'h424787ab},
  {32'h444431ee, 32'hc328f2c8, 32'h438a6343},
  {32'hc3929d48, 32'hc30dc44a, 32'hc390612b},
  {32'h43eac670, 32'hc15a297a, 32'h44023382},
  {32'hc3cc6d4c, 32'h439b5b67, 32'h40e1b1d1},
  {32'h44a7706a, 32'hc2b1f8cd, 32'h420d951c},
  {32'hc4a6938c, 32'hc2414be8, 32'h41669977},
  {32'h44d691a6, 32'hc38a7429, 32'hc2bbf75d},
  {32'hc41df914, 32'hc3915102, 32'hc31a47a3},
  {32'h442d41f4, 32'hc0c335a8, 32'hc33504c3},
  {32'hc49fe67f, 32'hc4270fd7, 32'h42197c40},
  {32'h44988c7c, 32'hc33769a7, 32'hc3133bba},
  {32'hc508e3d7, 32'hc2205d8e, 32'hc268297b},
  {32'h43a5fc5d, 32'h428b5efa, 32'h437ee4c4},
  {32'hc49b3576, 32'h43296662, 32'h431816a2},
  {32'h433b0100, 32'h4397d503, 32'hc36a67bd},
  {32'hc5096b24, 32'hc30c605e, 32'hc254e375},
  {32'h446fe2ba, 32'hc2f93edc, 32'hc39327da},
  {32'hc37b1878, 32'hc3820652, 32'hc33487f6},
  {32'h44a4325e, 32'h43bb563c, 32'h4285f664},
  {32'hc4c1f76f, 32'h4335486e, 32'h435cb96e},
  {32'h44e08362, 32'h423083c1, 32'hc345474c},
  {32'hc504cabd, 32'h42b5bc77, 32'hc10ce996},
  {32'h44d885f3, 32'hc387c7d0, 32'h420ef7aa},
  {32'hc4cc1899, 32'hc2ef19e9, 32'h42b257b2},
  {32'h440e416d, 32'hc2b8a5cc, 32'h426eb1c4},
  {32'hc4aaa6ca, 32'hc28ed76a, 32'h42581754},
  {32'h445277dd, 32'h437a3070, 32'hc403675e},
  {32'hc438fcae, 32'h431c3443, 32'hc356a96b},
  {32'h45057e14, 32'hc2ab5664, 32'h425a06d7},
  {32'hc440e430, 32'hc28fb7c9, 32'h41fceeed},
  {32'h449699c7, 32'hc1101658, 32'h3f324800},
  {32'hc4822fc4, 32'h4236a666, 32'hc31b76bb},
  {32'h44a0b53b, 32'hc3952338, 32'h43bc68f8},
  {32'hc514ad61, 32'hc2efb382, 32'h43a18fae},
  {32'h447ed4d0, 32'hc2695029, 32'h436dd672},
  {32'hc4850be5, 32'h42cf91bc, 32'hc260da04},
  {32'h44d4611e, 32'hc295094c, 32'h43375567},
  {32'hc4f838f7, 32'hc3be6bd6, 32'h42b68821},
  {32'h447ac249, 32'hc199bfea, 32'h4207df25},
  {32'hc3a07aa1, 32'hc0cd16df, 32'hc3734a77},
  {32'h44de0d6d, 32'hc201511f, 32'h42300f34},
  {32'hc3b6c7e0, 32'hc38f1514, 32'hc329f7f5},
  {32'h45088065, 32'hc34111f9, 32'hc3b85a37},
  {32'hc3adc452, 32'hc2c11d6c, 32'h43093011},
  {32'h42a08330, 32'hc2f5f03a, 32'h434372a1},
  {32'hc4ebbdf9, 32'hc3b9e098, 32'h40f306ba},
  {32'h4432826a, 32'h433070ff, 32'h42d1d496},
  {32'hc38be052, 32'hc3873bea, 32'h43a2fb2e},
  {32'h43ba7e18, 32'hc40c70a8, 32'hc353732e},
  {32'hc4ddd30c, 32'hc3267bb0, 32'h43923e65},
  {32'h4504048e, 32'hc282ae5f, 32'h4369af93},
  {32'hc3a220b8, 32'h42ba0891, 32'h430a9b7d},
  {32'h450c59f7, 32'hc3bbaae8, 32'h43d67822},
  {32'hc0418400, 32'hc2c52c32, 32'hc2cab388},
  {32'h45032844, 32'hc38713b5, 32'h429a4260},
  {32'hc4c72028, 32'hc2f2aa9f, 32'hc20e6004},
  {32'h44d799f7, 32'hc3dcc313, 32'hc3a94f70},
  {32'hc4b1c4cf, 32'h42cb9f01, 32'h437a4a0d},
  {32'h43a9f678, 32'h439da555, 32'h434a3a4e},
  {32'hc4fb935e, 32'h41f3b1b1, 32'hc28f6c5e},
  {32'h43b52d2c, 32'hc4121845, 32'hc3b9715a},
  {32'hc40439d8, 32'hc2b46b3f, 32'hc3cfd59a},
  {32'h4409a88c, 32'hc3282fdf, 32'hc39ed3a9},
  {32'hc4da7bde, 32'h41a1a617, 32'hc3672e6b},
  {32'h450a5e06, 32'hc28206a0, 32'h43aea4e5},
  {32'hc492da71, 32'h4309bc79, 32'hc2a00762},
  {32'h44dae06e, 32'h43b0a3b7, 32'h421a6061},
  {32'hc49dfba4, 32'h42a131b0, 32'hc29dad83},
  {32'h4315a368, 32'hc3125718, 32'hc22443fc},
  {32'hc505944e, 32'h43804ee8, 32'hc1e21496},
  {32'h435038e0, 32'hc360bc7c, 32'h42ae7eac},
  {32'hc4f2dad2, 32'h42a0af14, 32'h439d1a8f},
  {32'h444b1b38, 32'h436a77b6, 32'hc2e4f5cf},
  {32'hc36ee2b8, 32'hc36a0213, 32'h42e58f2c},
  {32'h44e2cb88, 32'h41d5418e, 32'hc23b698d},
  {32'hc43faf98, 32'h438b0eb2, 32'h43bbcad3},
  {32'h44779db4, 32'hc37242ca, 32'hc34d26be},
  {32'hc38e7ac4, 32'hc2c0ca27, 32'h42a9ef3d},
  {32'h443eaf48, 32'h43277d4b, 32'hc2094ade},
  {32'hc4d292aa, 32'hc4073498, 32'h433963a0},
  {32'h4506ee0e, 32'h4380b21e, 32'h42fb33d8},
  {32'h42b84186, 32'h4088809c, 32'h439feb53},
  {32'h44a104bd, 32'hc23d3cdf, 32'h430ea7e8},
  {32'hc4dfd7e8, 32'h437a9216, 32'hc32947c2},
  {32'h44721790, 32'hc40c44bb, 32'hc30d944d},
  {32'hc438c96c, 32'hc1a81d6d, 32'h421915ab},
  {32'h450b64ba, 32'hc2fa6a62, 32'hc31616c2},
  {32'hc4e9a2e3, 32'h4295c5da, 32'hc3235749},
  {32'h44a24627, 32'hc305e66e, 32'h4310a90e},
  {32'hc4827360, 32'hc3806118, 32'hc2a4c7e2},
  {32'h4410cd74, 32'h42b4fd6e, 32'hc40ece22},
  {32'hc4d475b2, 32'hc3822b71, 32'hc3c48d06},
  {32'h436e0720, 32'h42d44de4, 32'hc339f39a},
  {32'hc4e3f8ae, 32'hc3822f5b, 32'h43e63ffb},
  {32'h44e6f224, 32'h42cb34f1, 32'hc38d44f6},
  {32'hc484f48e, 32'h4253dddb, 32'hc31e9010},
  {32'h44ef2909, 32'h42b5f95d, 32'h42c9eb29},
  {32'h42ee9b00, 32'h4332e035, 32'h424f79cc},
  {32'h44ff7a60, 32'hc30bb472, 32'h431d88d4},
  {32'hc5064e9e, 32'hc36d0335, 32'h4381e52a},
  {32'h444bff92, 32'h42b7fa89, 32'hc334d864},
  {32'hc504b9bc, 32'h43b66f97, 32'hc3079064},
  {32'h44c535c0, 32'h42d491e9, 32'h42ae64ee},
  {32'hc458aa92, 32'h4343aa12, 32'hc2940ca0},
  {32'h448652df, 32'h430e690b, 32'h4299c5e1},
  {32'hc406774a, 32'hc22430fb, 32'hc2d81d73},
  {32'h429682c0, 32'hc33286ae, 32'h436554f3},
  {32'hc4abab0d, 32'h4385e91e, 32'h40d2c5f4},
  {32'h44410481, 32'hc386b0aa, 32'h42d958c8},
  {32'hc4c90ed8, 32'h4190f024, 32'h43242cd3},
  {32'h448ec058, 32'h434709a8, 32'hc34d0ae6},
  {32'hc4a35380, 32'h42a9955d, 32'h431b252d},
  {32'h44d7d7cf, 32'h403400a0, 32'hc388c66e},
  {32'hc41bcf44, 32'hc39af5e4, 32'hc3eede1b},
  {32'h43a5027b, 32'hc36f0536, 32'hc1c8176e},
  {32'hc4c590f5, 32'h435f029b, 32'hc3c515ae},
  {32'h44f77558, 32'h43331301, 32'h41b38185},
  {32'hc4b943c4, 32'h4329b905, 32'hc383ad36},
  {32'h437b6dcc, 32'hc220304b, 32'h4214c434},
  {32'hc505d5f3, 32'h4376750a, 32'h40837b42},
  {32'h43e37144, 32'hc3497134, 32'hc1f92949},
  {32'hc372a658, 32'hc3803330, 32'h4343322c},
  {32'h44c011d5, 32'hc27b5176, 32'h43b692f5},
  {32'hc48f7916, 32'h42fed2f8, 32'hc3cee02e},
  {32'h4388e550, 32'h43a7181a, 32'h43da0dcd},
  {32'hc290a208, 32'h4326461c, 32'h43937eaf},
  {32'h44a817d0, 32'h42e4189c, 32'h43bd3598},
  {32'hc4ae2a21, 32'hc2beccc1, 32'h42adcdcf},
  {32'h440f9eac, 32'h42740ece, 32'h42fb51e3},
  {32'hc4854fe1, 32'hc2ff2592, 32'h40167cfb},
  {32'h44bbc4ca, 32'h42ef7644, 32'h4385b47f},
  {32'hc4cf31c5, 32'hc3df8cbe, 32'hc21461e0},
  {32'h44ffb109, 32'h42d42944, 32'h43ce767e},
  {32'hc3fb114a, 32'h43d30fc3, 32'hc3287fd2},
  {32'h4508ca4f, 32'hc3722a16, 32'h43244977},
  {32'hc41fb36e, 32'hc3dd3ca9, 32'hc3172bcb},
  {32'h4457a1e8, 32'h404c94ea, 32'hc3342dd1},
  {32'hc48b0360, 32'h432f17c6, 32'h41e7e34d},
  {32'h43e68184, 32'hc20a72b4, 32'h42b3e37f},
  {32'hc503d808, 32'h438ec69b, 32'hc39cf665},
  {32'h44a13f04, 32'hc368b319, 32'h43554736},
  {32'hc4e1f1a4, 32'h429b15df, 32'hc240ff7f},
  {32'h44ec197c, 32'h428748f3, 32'hc2b011d9},
  {32'hc47cb8b4, 32'hc21c0a96, 32'hc41aaf43},
  {32'h44ff4dd6, 32'h43503e54, 32'hc2844001},
  {32'hc458fe24, 32'h41e67efe, 32'h434a2b5d},
  {32'h449b2b5e, 32'hc2c50e60, 32'h43b226ca},
  {32'hc414b9c0, 32'hc3b924ba, 32'h42c92eda},
  {32'h450a459d, 32'hc2fdc613, 32'hc3acfa8f},
  {32'hc46176db, 32'hc39282d3, 32'hc33c0e37},
  {32'h44d59133, 32'h42e62fc8, 32'h43209458},
  {32'hc4dd332d, 32'hc315fbb9, 32'h4325064b},
  {32'h445f6f3a, 32'h43d58f40, 32'hc1c3a6c6},
  {32'hc39153a8, 32'hc28ea6cd, 32'hc2df7312},
  {32'h44e86510, 32'hc312fe1a, 32'hbf22dee8},
  {32'hc3b1d31e, 32'h430e1529, 32'hc1254def},
  {32'h44f7dbef, 32'h41d735c3, 32'hc2068d75},
  {32'hc43d7d64, 32'hc3ef108d, 32'h4388eb59},
  {32'h4515ccc5, 32'h4278dc10, 32'hc304814f},
  {32'hc4eb9621, 32'hc2f2a908, 32'h42525ae5},
  {32'h44a8adfd, 32'hc35b9338, 32'hc2ca8f4e},
  {32'hc4eb6f34, 32'hc366be33, 32'h41e684a2},
  {32'h4435d3ec, 32'h43b8b91d, 32'hc3b5dbe8},
  {32'hc48de1d2, 32'h433baeab, 32'h42e0896d},
  {32'h44f2376f, 32'h42fdc4d6, 32'hc3133ddf},
  {32'hc505de73, 32'hc2e33b51, 32'hc39d530a},
  {32'h4383f7c8, 32'hc270373a, 32'h4324fa49},
  {32'hc3d26330, 32'hc3137ed9, 32'h4266710e},
  {32'h43ddb0b0, 32'hc13e80ae, 32'h434191a9},
  {32'hc503ee9f, 32'hc3c14086, 32'hc3b77317},
  {32'h4481cdc5, 32'h42e0cfdc, 32'hc322ef3b},
  {32'hc449d93c, 32'hc37d16f6, 32'hc284aa52},
  {32'h4437ab32, 32'hc0951226, 32'h42b1940d},
  {32'hc402c9ea, 32'h439d19c0, 32'hc247a60d},
  {32'h42d250a0, 32'hc2e7226d, 32'h433894f8},
  {32'hc4a76399, 32'h42cfe374, 32'hc3087484},
  {32'h44f110d8, 32'hc2f6a3c4, 32'h437ba3d0},
  {32'hc4f1f9a6, 32'h4248d0ad, 32'h433aa6ca},
  {32'h44e0acb8, 32'hc2726957, 32'h43010972},
  {32'hc3324bce, 32'hc2078657, 32'hc281f7ce},
  {32'h4499ae16, 32'hc3ad9e8f, 32'hc3b2b683},
  {32'hc459d50c, 32'hc1101384, 32'hc2960ef6},
  {32'h4365d6dc, 32'h43811303, 32'h431affc1},
  {32'hc4cc2786, 32'hc3013bfe, 32'h4365308d},
  {32'h44add588, 32'hc2bc7400, 32'h43d04727},
  {32'hc4ab7f4b, 32'hc33f93f4, 32'h42d436ab},
  {32'h44b8f8d9, 32'h42842d19, 32'hc34e33fa},
  {32'hc4856b62, 32'hc3d90f24, 32'hc161ab80},
  {32'h4405afe4, 32'hc337b613, 32'hc38b5c42},
  {32'hc493f3c9, 32'hc3a38c1a, 32'h42c1eded},
  {32'h44969cd4, 32'h4331ca45, 32'hc1fb7cf0},
  {32'hc4f7af58, 32'h43b10862, 32'hc3331f88},
  {32'h44060af8, 32'h43402b97, 32'hc37a0719},
  {32'hc4b274d8, 32'hc1cb172d, 32'hc3cc4465},
  {32'h4517b8cf, 32'hbbd3f800, 32'hc161718d},
  {32'hc4fd459d, 32'h43e6a8ce, 32'h4390f93c},
  {32'h442943dc, 32'hc29fb93c, 32'h428fa404},
  {32'hc4988b57, 32'h42b2ce5b, 32'hc3574605},
  {32'h441faef2, 32'h439ce7ae, 32'h43775a2a},
  {32'hc2af6998, 32'hc28b1f91, 32'h41b53b55},
  {32'h44cebde2, 32'h43c6066d, 32'hc3612e85},
  {32'hc4855357, 32'hc3223247, 32'hc2dc202c},
  {32'h4433cc85, 32'h42fd978d, 32'h429cb862},
  {32'hc50b6787, 32'h42d61447, 32'hc208c239},
  {32'h447f4f74, 32'h42a98903, 32'h43668fba},
  {32'hc508fd1b, 32'hc21c4118, 32'hc211d782},
  {32'h431be62c, 32'h42e96041, 32'hc28fc110},
  {32'hc4acbe9d, 32'hc3c6fc7a, 32'h43672792},
  {32'h43c63432, 32'hc2eecb57, 32'h42f62264},
  {32'hc4eca848, 32'hc3257bc1, 32'hc238fc55},
  {32'h44b4c266, 32'h43944461, 32'hc2b6bb7c},
  {32'h42dbea40, 32'h438c49e9, 32'hc3c23209},
  {32'h44e5680a, 32'h41d5259d, 32'h419aeaad},
  {32'hc4fd99f9, 32'h43033493, 32'hc2294810},
  {32'h438af09a, 32'hc2b8fed0, 32'hc31d1aeb},
  {32'hc49e41b2, 32'h4225adbf, 32'h429978d4},
  {32'h45101612, 32'h3f8d1750, 32'h42706e07},
  {32'hc3f67f84, 32'h43879b68, 32'h419239a2},
  {32'h4507ec20, 32'h439c5ee7, 32'hc2907afa},
  {32'hc3c042dc, 32'hc3ad0e44, 32'h42aa9d3f},
  {32'h449644be, 32'hc209d007, 32'hc39b50ca},
  {32'hc4bbac37, 32'hc3708b9a, 32'h425416c6},
  {32'h44605118, 32'hc3825070, 32'hc32dfd37},
  {32'hc4b793eb, 32'hc2e90e7b, 32'hc3b3b126},
  {32'h44898033, 32'hc2d92a20, 32'hc31a18db},
  {32'hc3e418fa, 32'h4342c262, 32'hc2a2882f},
  {32'h450920dd, 32'hc3a4304d, 32'h421e4ed3},
  {32'hc4fd98ca, 32'h43abb99f, 32'h435a0bb3},
  {32'h44a3dbc5, 32'h43cc8ca8, 32'hc2fcded4},
  {32'hc513cfbd, 32'h41d157cc, 32'h415f1fca},
  {32'h45151a12, 32'hc35265bb, 32'h423c4d7d},
  {32'hc33a06e6, 32'h429eaac0, 32'h42f7df73},
  {32'h44e4e573, 32'h4336a5d0, 32'hc2f8171e},
  {32'hc3939546, 32'hc269ca2f, 32'hc3ae75d9},
  {32'h4508572b, 32'hc2d582ca, 32'hc180e70f},
  {32'hc4f4cd3d, 32'h430600b2, 32'h433e14b9},
  {32'h447c64e6, 32'h4385bfcf, 32'hc331a24d},
  {32'hc3fa5350, 32'hc3012964, 32'hc1d4a4e7},
  {32'hc2c4d650, 32'hc3547131, 32'h408aa510},
  {32'hc45e120a, 32'hc31f95ac, 32'hc215aa16},
  {32'h4510c7c0, 32'h42e3a93d, 32'hc378e6a3},
  {32'hc4c50780, 32'h3fb1ae00, 32'h40bc6874},
  {32'h44d4ab36, 32'h43387336, 32'h439d1231},
  {32'hc4034af6, 32'h4291dd70, 32'hc34666dc},
  {32'h44d9c2e8, 32'h42e16029, 32'h434a2e67},
  {32'hc4ae3c62, 32'h43c4ce82, 32'h4397b0b3},
  {32'h448bdc26, 32'h43292fb7, 32'h43f11e34},
  {32'hc51ef462, 32'hc3b363e2, 32'hc2870c39},
  {32'h44f2fcdb, 32'h424eb4fb, 32'hc1758152},
  {32'hc4d57123, 32'hc3078f05, 32'hc3e2e5b6},
  {32'h439ef3fb, 32'h41ff2f76, 32'h431e7f4a},
  {32'h431a6038, 32'hc380091f, 32'hc3dae311},
  {32'h4538de7c, 32'h4225a25a, 32'hc2249410},
  {32'hc50315fa, 32'h433445af, 32'hc401a9f8},
  {32'h434fc278, 32'hc3362c39, 32'h432a40a2},
  {32'hc4751720, 32'h42a6b503, 32'hc3202011},
  {32'h448fa841, 32'h42fceb36, 32'h41b12b6e},
  {32'hc29c2290, 32'hc2c10b01, 32'h433fb2f2},
  {32'h447f20e5, 32'h42c09a00, 32'h4351bcad},
  {32'hc5009e2b, 32'hc2a12886, 32'h43a5f096},
  {32'h44b807c2, 32'hc2aa959a, 32'h43807948},
  {32'hc4b0f11d, 32'hc30767db, 32'h4313c1e0},
  {32'h430a09e0, 32'hc25f9e86, 32'hc2856c34},
  {32'hc40a2e94, 32'hc2ac3e82, 32'h42888526},
  {32'h44a5953c, 32'hc0f77be4, 32'h40d75a78},
  {32'hc39535d8, 32'h41ef9966, 32'h4102a7a6},
  {32'h44831981, 32'h43e14a12, 32'h433c76b0},
  {32'hc4548fab, 32'h430ea2cf, 32'h4337da9c},
  {32'h44d6c492, 32'h42c7b934, 32'hc2a49a8b},
  {32'hc39f1b48, 32'h425ce77c, 32'h41e0ff88},
  {32'h44bfc61b, 32'h42a9dfef, 32'h434a7917},
  {32'h4284bd28, 32'h431d9a53, 32'h43cbf442},
  {32'h4450e656, 32'h41e54afa, 32'h4382a1da},
  {32'hc4cb7898, 32'h42de91a4, 32'hc367ffd9},
  {32'h44cadcdf, 32'h438df9ea, 32'hc38d3231},
  {32'hc47c6356, 32'h42897acc, 32'hc32a8142},
  {32'h44c3edd1, 32'hc29733b6, 32'hc32e44a2},
  {32'hc4206766, 32'hc274106a, 32'h427032c3},
  {32'h450b596a, 32'h42f0a469, 32'h4316bfdc},
  {32'hc4b26279, 32'hc33c9374, 32'hc2c7034c},
  {32'hc24fe15f, 32'h43924d24, 32'h42b1ee2f},
  {32'hc4d4025a, 32'h4399e687, 32'hc395492d},
  {32'h44584358, 32'h42dd93bc, 32'h43335544},
  {32'hc3afcaa0, 32'hc30bccad, 32'hc3396b53},
  {32'h4462aeec, 32'hc2e11978, 32'hc2d471b2},
  {32'hc49f8ce7, 32'hc3e97809, 32'h435cad03},
  {32'h43b1ebfa, 32'hc381ec3c, 32'h43485958},
  {32'hc4f15e42, 32'hc23e680f, 32'h422964a8},
  {32'h438a2630, 32'hc38810ad, 32'h42a73c91},
  {32'hc36869b0, 32'h435dcfa7, 32'hc3ad4175},
  {32'h43996c88, 32'hc2ea7ca5, 32'h4396b4dd},
  {32'hc50459dc, 32'h41877f3f, 32'h41d31c96},
  {32'h4507e9a6, 32'hc2a2875a, 32'hc35ecdc1},
  {32'hc4e34a84, 32'hc319af73, 32'hc1788b40},
  {32'h445d28f5, 32'hc331b0ed, 32'hc3c722d0},
  {32'hc41b3452, 32'hc38654e6, 32'hc2d2fc39},
  {32'h42ed86b0, 32'h43211a2f, 32'hc29393a4},
  {32'hc5096ec4, 32'h4375fa5d, 32'h43420a33},
  {32'h44b34129, 32'hc2d8ffd5, 32'h438f4a23},
  {32'hc4b71d69, 32'h433f6b5d, 32'hc1c8530b},
  {32'h449cb251, 32'h42d84d9c, 32'hc322e833},
  {32'hc52c1336, 32'h4384ee0f, 32'hc3195598},
  {32'h451bf795, 32'hc397e3bd, 32'h438cad66},
  {32'hc2e469cd, 32'h43b3d654, 32'hc2be3047},
  {32'h4506271f, 32'hc2f9d696, 32'hc289154d},
  {32'hc51c7ebb, 32'h428325a7, 32'hc2ade0d1},
  {32'h44b772d0, 32'h430c32b1, 32'h41db0328},
  {32'hc5030388, 32'h438f4f39, 32'h42c99016},
  {32'h446dcfc8, 32'h4295d2da, 32'h431a97b3},
  {32'hc4d32596, 32'hc380322d, 32'h41abcc31},
  {32'h450bf0ed, 32'hc334363b, 32'h438b2794},
  {32'hc4342f95, 32'h42ff485d, 32'h4383c2da},
  {32'h4512f250, 32'h43b4b71e, 32'h42efdec9},
  {32'hc4c30af8, 32'h43adda34, 32'hc3094060},
  {32'h44385df4, 32'h43218b02, 32'hc2beee78},
  {32'hc3fe2dac, 32'h424b49fa, 32'h40e461e1},
  {32'h43775464, 32'h42c4265f, 32'hc3c20a77},
  {32'hc4648e6c, 32'hc3877a81, 32'hc2e3d7a6},
  {32'h4507aeb5, 32'hc3c28283, 32'hc19e1501},
  {32'hc47869d6, 32'h42de5329, 32'hc261e19d},
  {32'h44ee7c88, 32'hc18ebda8, 32'h4310799a},
  {32'hc45ef2c8, 32'h421a42d3, 32'hc37aa94d},
  {32'h4385a9ac, 32'hc330cbcd, 32'hc3687614},
  {32'hc42ef8c2, 32'h42fb6d70, 32'hc31d4408},
  {32'h44ec5414, 32'h43bbf525, 32'h42588493},
  {32'hc50a98e1, 32'h43197448, 32'h432ceb6c},
  {32'h446798cc, 32'hc2020bda, 32'h42c7726e},
  {32'hc499f410, 32'hc243c4c4, 32'h42c818ca},
  {32'h44af6669, 32'h43290c96, 32'hc27b94c0},
  {32'hc490e8a4, 32'hc3b9994e, 32'h441257eb},
  {32'h44bfe30e, 32'h417236f5, 32'hc1b2128b},
  {32'hc4152f3c, 32'hc3cfd5aa, 32'h42de658f},
  {32'h44e016df, 32'h43162532, 32'hc2cdffa2},
  {32'hc5098b7e, 32'h42748d27, 32'h43923da4},
  {32'h44c65d8e, 32'h43976ec3, 32'hc3840d04},
  {32'hc34c168a, 32'hc2fad4ec, 32'h430b149d},
  {32'h44c67576, 32'hc0aa8588, 32'h43097b42},
  {32'hc3978b06, 32'h419b215e, 32'h438ba43f},
  {32'h45037139, 32'h419f943e, 32'hc274c2b8},
  {32'hc4a1099d, 32'hc2a9235a, 32'h430232a3},
  {32'h433736d8, 32'h42a344ae, 32'h42bdf397},
  {32'hc504c878, 32'hc237730e, 32'h435da852},
  {32'h44fc08e9, 32'h42470c7e, 32'hc1df988e},
  {32'h41e88680, 32'hc2e10164, 32'h43a4d932},
  {32'h4512761e, 32'h431de50e, 32'hc3b2b428},
  {32'hc37b2409, 32'hc3515153, 32'hc3061b23},
  {32'h44b64340, 32'h43758411, 32'hc2ad8644},
  {32'hc49b01a4, 32'hc2dca262, 32'h4291daa5},
  {32'h44082d96, 32'hc0eef158, 32'h42233da5},
  {32'hc4a13a75, 32'hc3fe6440, 32'h414a1762},
  {32'h450e7dfb, 32'hc377426a, 32'h42a9643a},
  {32'hc495f9df, 32'hc176ee76, 32'h4404c3d5},
  {32'h44d55676, 32'h43bd542e, 32'hc3583007},
  {32'hc4138b74, 32'h426b6620, 32'h43c31a08},
  {32'h450afc49, 32'h4086d6b3, 32'hc2deff6a},
  {32'hc4f373d8, 32'h4359c197, 32'hc38df37a},
  {32'h44f14078, 32'hc3439909, 32'hc3702f0b},
  {32'hc3f15b58, 32'hc1f8ec49, 32'hc28de82c},
  {32'h43b1a31c, 32'h43c6344c, 32'h42838f5b},
  {32'hc39e5ed0, 32'hc31d8eb8, 32'h42e5f596},
  {32'h42f7e056, 32'hc33c9504, 32'hc38597cd},
  {32'hc477a3e4, 32'h4201c49d, 32'h43a7e756},
  {32'h44d67108, 32'h433bfb81, 32'hc2cdac7f},
  {32'hc3f7c2bc, 32'hc28018df, 32'h42a8465a},
  {32'h44f67d40, 32'h43762181, 32'h42de8a0e},
  {32'h43483d3c, 32'hc3322a86, 32'h4386199a},
  {32'hc4b20ca4, 32'h43b6396b, 32'hc348ac41},
  {32'h44e1c9ee, 32'h4352d2dc, 32'hc375b882},
  {32'hc50614c1, 32'h42d6537b, 32'hc252b025},
  {32'h44963a67, 32'h42fbfdb0, 32'hc327eb2f},
  {32'hc4ced11f, 32'h438eac64, 32'h42b1999c},
  {32'h4345c840, 32'hc35d89fe, 32'hc3cacb04},
  {32'hc508e70f, 32'hc2e2d277, 32'hc3554935},
  {32'h44ab2987, 32'hc3e58031, 32'hc2900dd5},
  {32'hc4febcc5, 32'hc381607e, 32'hc38e79a1},
  {32'h4421a902, 32'h430d846d, 32'hc10fcd77},
  {32'hc50db6f6, 32'hc2fd4201, 32'h404eef58},
  {32'h44a38372, 32'h4283174a, 32'hc2d5dea8},
  {32'hc50ca7e2, 32'hc31df145, 32'hc3618336},
  {32'h429d74d5, 32'hc32344cc, 32'h43449682},
  {32'hc48d4987, 32'h4192f8c4, 32'h431d6060},
  {32'h449b6aea, 32'h42d9788d, 32'hc3d5a785},
  {32'hc50b12d4, 32'hc12654a6, 32'h428fd7db},
  {32'h446c973a, 32'h43966786, 32'h425f08fd},
  {32'hc500eb39, 32'h42c952f1, 32'hc2b4159e},
  {32'hc2e1e16c, 32'hc3265408, 32'hc38ec73a},
  {32'hc4122b14, 32'hc30fc2da, 32'h42d69d3f},
  {32'h44b10bd7, 32'hc2dbb5cd, 32'hc3a36424},
  {32'h41e3f980, 32'hc31e89ab, 32'h432b1ccc},
  {32'h44782144, 32'hc2e10bd9, 32'hc24bc2c1},
  {32'hc3b82c9d, 32'hc3d2ad6a, 32'h438ba74f},
  {32'h44b94b4f, 32'h430b4fc3, 32'hc2acb718},
  {32'hc4b44e3e, 32'hc2b6f6c4, 32'hc3309a04},
  {32'h43354380, 32'hc3c8911f, 32'h4291b5ab},
  {32'hc40294e0, 32'hc29ae240, 32'hc397694f},
  {32'h42c3a530, 32'hc2b9af39, 32'h42b3d955},
  {32'hc4e42470, 32'hc2b3c9aa, 32'hc4268c8d},
  {32'h44a89ddb, 32'h433d70b0, 32'hc287d814},
  {32'hc4e7553f, 32'h43e8dc67, 32'hc345977b},
  {32'h44940261, 32'h42f5c033, 32'hc355ab47},
  {32'hc50a5f7a, 32'h433245c8, 32'h43b45e64},
  {32'h4504fd6c, 32'hc2940088, 32'hc375c45a},
  {32'hc4f60975, 32'h4307056c, 32'h4354d41c},
  {32'h44afde44, 32'hc30d94a0, 32'h43885392},
  {32'hc4d6e256, 32'h438e6813, 32'hc36241f4},
  {32'h44b4594f, 32'hc31127cb, 32'hc2a2de8d},
  {32'hc3cf9110, 32'hc2205acc, 32'h438cd53f},
  {32'h44f51656, 32'hc3c58b25, 32'hc2201446},
  {32'hc439dfcc, 32'h42020fac, 32'h406458fe},
  {32'h449dd119, 32'hc2e0de89, 32'h41b67709},
  {32'hc4abe02d, 32'h43d15fc4, 32'h43aa59e2},
  {32'h4388fb63, 32'hc363e1cc, 32'hc13493d2},
  {32'hc2d68684, 32'h43792b8f, 32'hc3351098},
  {32'h443e4fb4, 32'h422e0c5b, 32'h43219b3a},
  {32'hc47193e6, 32'hc2ec4e07, 32'h43363a67},
  {32'h43c0f0fa, 32'h43c87e8c, 32'h420330c8},
  {32'hc43f3939, 32'h42c852b7, 32'hc33e529e},
  {32'h44da271a, 32'h441ac0c5, 32'h42d01120},
  {32'hc4a3d198, 32'h4338af86, 32'hc2a4bd7d},
  {32'h446584e1, 32'hc2fecb4f, 32'hc3b44d50},
  {32'hc4e4f4e8, 32'h42e3ccbb, 32'hc3ef714f},
  {32'h449c4a20, 32'h43dcecd0, 32'hc2891e01},
  {32'hc42de0fe, 32'h405255ac, 32'hc3ad172a},
  {32'h44d6464c, 32'hbfd75ec9, 32'hc39ce2d5},
  {32'hc45d72cd, 32'hc2d2ef47, 32'hc1c95ab0},
  {32'h43a5ce78, 32'hc3a1893b, 32'h4399b4e7},
  {32'hc31d3198, 32'h439eb583, 32'h42efa66f},
  {32'h4295c930, 32'hc389adb7, 32'h4307ea48},
  {32'hc4b8a8ea, 32'hc2318c79, 32'h43699a8e},
  {32'h43aff473, 32'h43621de5, 32'h434e8350},
  {32'hc48cd6fc, 32'hc3896aee, 32'hc209e574},
  {32'h44e87320, 32'hc1ca9c2a, 32'hc30106e9},
  {32'hc4c8aeb1, 32'hc2eb4fe7, 32'hc316f41a},
  {32'h44e73adc, 32'h42a43a3b, 32'h4035b74c},
  {32'hc407e373, 32'hc28afda3, 32'hc250fdf4},
  {32'h44cc2e98, 32'h4374ac9f, 32'h43098fc3},
  {32'hc2fe99a0, 32'h427a7651, 32'hc3a03778},
  {32'h44f8c061, 32'hc41aa9c5, 32'h438f0ec9},
  {32'hc487d456, 32'hc30b317d, 32'h42dff940},
  {32'h450112b7, 32'hc43a4db2, 32'hc29311da},
  {32'hc4a6cbaa, 32'h4293213e, 32'h426bbe21},
  {32'h4369e430, 32'hc3bd6f67, 32'h41c51782},
  {32'hc4bcfa41, 32'hc2a98192, 32'h42aed6c6},
  {32'h4509b434, 32'hc351a653, 32'h3fbfb652},
  {32'hc3c3f688, 32'h431509dc, 32'h4305d12b},
  {32'h439aa480, 32'h4366841f, 32'h430ad48d},
  {32'hc493edcf, 32'h43a2d720, 32'h43c86fef},
  {32'h44cd490f, 32'hc2a62807, 32'hc31f12b0},
  {32'hc503b3c2, 32'hc21c2096, 32'hc2c7b7a3},
  {32'h45041bdf, 32'h412eea1d, 32'h43af7c0b},
  {32'hc4991c33, 32'hc3101bc8, 32'h44355069},
  {32'h44c623e8, 32'hc2751646, 32'hc313d3c8},
  {32'hc461b9af, 32'hc3a49121, 32'hc19447d7},
  {32'h450e1487, 32'hc2662fe4, 32'h43259074},
  {32'hc4de8557, 32'h4386c27b, 32'h42ba9aec},
  {32'h4478c749, 32'h4307b917, 32'h42c96eaf},
  {32'hc51c1e90, 32'h43843158, 32'hc33869eb},
  {32'h450ae854, 32'hc34431de, 32'h43e3682e},
  {32'hc4e75a9e, 32'hc366f03c, 32'hc3bcf371},
  {32'h44e7fa0c, 32'h43ba34d4, 32'h42d2865c},
  {32'hc455ff69, 32'h42dd6df3, 32'h423e34c1},
  {32'h4499a4c6, 32'h4402ec72, 32'hc39397bc},
  {32'hc4be3e1c, 32'hc3073c2a, 32'hc2327f10},
  {32'h43ced330, 32'hc29e1fa3, 32'hc37954fe},
  {32'hc4bf9ccb, 32'h43c9b978, 32'h43e75492},
  {32'h449f4d33, 32'h43bb93f2, 32'h420e92e9},
  {32'hc4a469ed, 32'h43e98672, 32'h42e67e02},
  {32'hc2b8d47c, 32'h41bfa8c5, 32'h41dd2b52},
  {32'hc42f46c1, 32'h43de5183, 32'h43ad6676},
  {32'h44c19e4f, 32'h4303eb8d, 32'hc398e434},
  {32'hc4070065, 32'h43069888, 32'hc2b2ef58},
  {32'h439e4396, 32'hc3ea2b8b, 32'h42fac013},
  {32'hc3d3a400, 32'hc38b0d66, 32'hc398e5d3},
  {32'h44cbebc1, 32'h42561cc2, 32'h42217de5},
  {32'hc44523f2, 32'h4330617f, 32'hc33296fc},
  {32'h44832f63, 32'hc39e20b1, 32'hc2a85882},
  {32'hc4c79f9c, 32'h4381ca05, 32'h4399858b},
  {32'h44e3b258, 32'hc31d72dc, 32'h42d76171},
  {32'hc46d0626, 32'h43a59466, 32'hc1a95e3d},
  {32'h44b59417, 32'h43a207dc, 32'h4339f6d1},
  {32'hc4130736, 32'hc3def923, 32'hc1d8b75c},
  {32'h44a9bac2, 32'hc361f130, 32'hc3949a9e},
  {32'hc478acd9, 32'h43f89251, 32'hc38af62b},
  {32'h448dcd51, 32'hc38649f1, 32'hc265aaab},
  {32'hc4fbcd4d, 32'h433bae4c, 32'h43e03655},
  {32'h44ef4960, 32'hc3296228, 32'hc3eb5099},
  {32'hc4b3e5d4, 32'h42da1f93, 32'h4272b254},
  {32'h44d7088f, 32'h4354c3db, 32'h42d8898a},
  {32'hc473507a, 32'h4399e3f9, 32'hc26ea7fc},
  {32'h4488601c, 32'hc2b63423, 32'hc333f23e},
  {32'hc4cda77e, 32'hc1e0f8c7, 32'h43159864},
  {32'h44972f1c, 32'hc2589860, 32'h401a7498},
  {32'hc332cb24, 32'h42803933, 32'h431ed3f5},
  {32'h441cd4b2, 32'hc3cdb32c, 32'h421cddc1},
  {32'hc4102b56, 32'hc2254c2d, 32'hc2ecd615},
  {32'h44c7856a, 32'h430815fe, 32'h43c423f5},
  {32'hc4e77907, 32'hc381521c, 32'hc2a7bff6},
  {32'h452144af, 32'h43bae1fd, 32'hc1013a49},
  {32'hc43142b6, 32'hc3aaa5b2, 32'h435ab1aa},
  {32'h44d9a810, 32'h418a51c5, 32'h43219a02},
  {32'hc46bb49d, 32'h40e8725b, 32'hc11143b6},
  {32'h44c1fa39, 32'h419523ef, 32'hc3ea4faa},
  {32'hc408480c, 32'hc361fa2f, 32'hc306493c},
  {32'h44d08cea, 32'hc2aaa1ea, 32'hc29f7a18},
  {32'hc4d57dc4, 32'h439793bc, 32'hc3b564b8},
  {32'h43bd457c, 32'h41a9a45a, 32'h42cf7f79},
  {32'hc4153090, 32'h3fd1ccfa, 32'hc26ccc10},
  {32'h4404ab2a, 32'h423f3c85, 32'h43947b4e},
  {32'hc4e66716, 32'h401db490, 32'h435e82cf},
  {32'h44bd2f90, 32'h41817db2, 32'hc29b6fda},
  {32'hc402ebc4, 32'hc206942d, 32'hc2e3bfc8},
  {32'h443c54b4, 32'h4256db8a, 32'h436da193},
  {32'hc3e5e9b2, 32'h435fa9bb, 32'h42dcea3a},
  {32'h43ddad38, 32'hc1e0b4d9, 32'hc3cb39a8},
  {32'hc4d4eee8, 32'hc2aa38eb, 32'hc4125cc9},
  {32'h441c5302, 32'hbfd71233, 32'hc33a0bbe},
  {32'hc4674194, 32'hc383eb72, 32'h43f5c5be},
  {32'h44bbb49c, 32'hc3746f65, 32'hc146e0f6},
  {32'hc4ef543f, 32'hc3f47be5, 32'hc382a52e},
  {32'h447c5a72, 32'hc2ad8dd4, 32'h42326974},
  {32'hc4d315bc, 32'h433d5d96, 32'hc31edbd6},
  {32'h44dc2cc9, 32'h4225de19, 32'h42f6e28c},
  {32'hc4b23259, 32'h438cd2ba, 32'h424241bd},
  {32'h44e3b072, 32'hc3741839, 32'hc3dd485a},
  {32'hc508a30d, 32'h434d65a1, 32'hc239fe99},
  {32'h42505d9c, 32'hc3cd70c7, 32'hc3239427},
  {32'hc4c1525d, 32'hc3326c2a, 32'h4040dcbc},
  {32'h43833bb0, 32'hc2f435b5, 32'h438f8fd8},
  {32'hc420cf2e, 32'h4196ddac, 32'h43183cbf},
  {32'h449544bc, 32'hc3adaced, 32'hc0fc7e4e},
  {32'hc505858f, 32'hc42eaf36, 32'h43c5cf60},
  {32'h421f1a40, 32'h416e422d, 32'hc3276df4},
  {32'hc4925777, 32'hc37f85fc, 32'hc38f18c5},
  {32'h438bfb39, 32'hbf265d20, 32'hc25b5490},
  {32'hc24a03e4, 32'hc21a1dbb, 32'h43083f4a},
  {32'h44dbecdb, 32'hc2b6e125, 32'hc2d50704},
  {32'hc424774c, 32'h41b2b234, 32'h43a0af1a},
  {32'h4213b780, 32'h4369d875, 32'hc3c585e3},
  {32'hc409b74b, 32'hc33d451a, 32'h4327df73},
  {32'h43d21aac, 32'h431b4ea3, 32'hc1eea0d1},
  {32'hc42d9385, 32'hc32acde2, 32'hc3b1caaa},
  {32'hc288947c, 32'h4310cbc4, 32'h423304bd},
  {32'hc48fdf69, 32'h4336d24b, 32'h440a0958},
  {32'h44e46f8e, 32'hc2e12f98, 32'h4249d5c1},
  {32'hc2dc81bc, 32'hc3a9e725, 32'h43617b25},
  {32'h445e22da, 32'h43571185, 32'hc3168d5e},
  {32'hc47d0242, 32'h43f105ea, 32'h433fe6c1},
  {32'h44105270, 32'hc2fb9d1b, 32'hc2a9f29a},
  {32'hc43fb682, 32'h43e0f71c, 32'h413b2e2b},
  {32'h44d524f7, 32'hc383fc59, 32'h420494bd},
  {32'hc3c55913, 32'h4382258e, 32'h429d9c3a},
  {32'h4502c005, 32'h43290387, 32'hc40ac696},
  {32'hc50c33d3, 32'h440b968b, 32'hc3d48c1a},
  {32'h4507445c, 32'hc3987753, 32'hc2f9a31a},
  {32'hc4b23b89, 32'hc338d2d3, 32'h42aff2c9},
  {32'h43c595d8, 32'h440ac551, 32'h43aea380},
  {32'hc4cb20f0, 32'hc37c9e69, 32'hc362eacc},
  {32'h445406eb, 32'hc2ed3f2b, 32'hc36ee848},
  {32'hc4b437e4, 32'h428e9d22, 32'hc2f0ae0b},
  {32'h43ab1640, 32'h42e824fa, 32'h41aab658},
  {32'hc42d0cc4, 32'hc349375a, 32'h42e8f083},
  {32'h449557b8, 32'h436d5d16, 32'h439db2ba},
  {32'hc4c0ef2e, 32'hc45dccee, 32'h40e6e236},
  {32'h44ec6831, 32'hc3d3a7a6, 32'h43b09f4d},
  {32'hc440b030, 32'h43090a6c, 32'h3fba9c98},
  {32'h43c4cdd6, 32'h42c919c8, 32'h41cc978b},
  {32'hc480af78, 32'h418569d1, 32'h43997a17},
  {32'h445aa801, 32'hc34889c2, 32'h4360f956},
  {32'hc4fa5243, 32'hc38d701b, 32'hc1ac1ea0},
  {32'h44bf0a65, 32'hc289725c, 32'h43b10493},
  {32'hc3cd12c4, 32'hc32bf279, 32'h4300665b},
  {32'h450f12ce, 32'h42e1ceb5, 32'h43b54e2e},
  {32'hc464e128, 32'h4323e977, 32'hc40b0b43},
  {32'h44ca818e, 32'h429f9ded, 32'hc30d9a58},
  {32'hc48baa98, 32'hc1d8d9a6, 32'h43f732ae},
  {32'h43f070d9, 32'h42e86203, 32'h4390fe84},
  {32'hc4e254e3, 32'hc368462d, 32'h435dbd5c},
  {32'h44b11611, 32'h43e5a9ef, 32'h434a434a},
  {32'hc3e99b8e, 32'hc3b16fe0, 32'h43677fe9},
  {32'h44b18fd8, 32'hc3415a64, 32'hc27bfe71},
  {32'hc32c2d2e, 32'h3f231ef9, 32'hc291a4e4},
  {32'h44073d28, 32'hc3109ffd, 32'hc34b58e3},
  {32'hc4b442e6, 32'hc3627442, 32'h438da53e},
  {32'h44a52c45, 32'hc364049b, 32'hc3570b1b},
  {32'h43512168, 32'h43cdf45e, 32'h43de04ac},
  {32'h440b83a8, 32'hc3558d42, 32'hc339c0dd},
  {32'hc4967030, 32'h43397e85, 32'h4385ba1e},
  {32'h44bfcb60, 32'hc3517988, 32'h4355b117},
  {32'hc51dff32, 32'hc366099d, 32'h4396b3d8},
  {32'h441d293f, 32'h437f1f2d, 32'h435b94c1},
  {32'hc4bdddde, 32'h4155e1c0, 32'h4306e0af},
  {32'hc41844f5, 32'hc33ae0a1, 32'hc1282ca2},
  {32'hc4140768, 32'hc35f94c0, 32'h3f715831},
  {32'h44b54ba4, 32'hc3339953, 32'h434204e1},
  {32'hc4d716e2, 32'h42deeb52, 32'hc24b8e0e},
  {32'h41862a00, 32'h438a91c2, 32'h42d0e24e},
  {32'hc4e72a40, 32'hc2d9dcea, 32'hc3552280},
  {32'h445ad1df, 32'h43306323, 32'hc358f239},
  {32'hc38a31f2, 32'hc3686f9f, 32'h43b885fd},
  {32'h450e23e5, 32'h4371be00, 32'hc308523f},
  {32'hc5024ce8, 32'h436fe6e8, 32'hc2b5bb98},
  {32'h444f3bc5, 32'h43ac2009, 32'hc1b0499a},
  {32'hc4dbd66e, 32'hc2930016, 32'h42f04c43},
  {32'h445c8d49, 32'hc3c97ba6, 32'h410678be},
  {32'hc50072a0, 32'hc2d25ee7, 32'hc3319c39},
  {32'h44df37f9, 32'h43929bef, 32'hc3cebd34},
  {32'hc4d29ccf, 32'hc28540af, 32'h43309752},
  {32'h450dd0ac, 32'hc361409a, 32'hc3704ec6},
  {32'hc437c244, 32'hc317006a, 32'h43b2e890},
  {32'h433cfdea, 32'hc1ef97c2, 32'h432a551a},
  {32'hc39aaefa, 32'h42c74324, 32'h42d686db},
  {32'h44216296, 32'hc3f7b898, 32'h40aed7fc},
  {32'hc4b83df1, 32'hc3107226, 32'hc3b70e79},
  {32'h44a6ec31, 32'hc1cf9130, 32'hc303c5b5},
  {32'hc4ed4307, 32'hc29d8f9e, 32'hc35d32ba},
  {32'h44f0b681, 32'hc282591f, 32'h42dd7cd8},
  {32'hc442bc7c, 32'hc33df175, 32'h43aa094b},
  {32'h4449ae4a, 32'hc3f624a4, 32'hc28cf5ac},
  {32'hc30b7d60, 32'h436ffdf2, 32'h42626766},
  {32'h443c5556, 32'h439a70cc, 32'hc3624690},
  {32'hc4c4a7f1, 32'h4335a056, 32'hc31b6550},
  {32'h44934178, 32'hc38fdef9, 32'hc24b2442},
  {32'h42515b40, 32'h4291e31a, 32'h4311470e},
  {32'h4492072e, 32'hc35f0c16, 32'h43278809},
  {32'hc4c9e7ce, 32'hc355a897, 32'hc26ac32a},
  {32'h447699fc, 32'hc265c5a2, 32'h432a7bbb},
  {32'hc3f8c55a, 32'hc1af3295, 32'hc30cfbcd},
  {32'h44fce9c2, 32'hc3a3acfd, 32'hc2c1c7d3},
  {32'hc4d09cee, 32'hc3adf09e, 32'h4304bd5b},
  {32'h44b4a1fe, 32'h4320549d, 32'h439350df},
  {32'hc5028ab2, 32'hc280edd7, 32'h43671cd3},
  {32'h450a5a9d, 32'h43363a22, 32'hc1a4105d},
  {32'hc47f4204, 32'h43ba1c85, 32'h41ab57c6},
  {32'h44216da3, 32'h42a933c1, 32'hc02b71b0},
  {32'hc41b3850, 32'hc325126e, 32'hc303fdc4},
  {32'h44c357e5, 32'h42f13164, 32'h41c3d593},
  {32'hc4f69409, 32'h43d06e88, 32'h438c44e7},
  {32'h442b4f1a, 32'h43e7ad05, 32'hc39c1174},
  {32'hc41bf2fc, 32'h421f065f, 32'hc35dedda},
  {32'h447b5a44, 32'hc3255e01, 32'hc3cb95de},
  {32'hc4dcede3, 32'hc2517d68, 32'hc1e84b06},
  {32'h44004c75, 32'h42dbfe89, 32'hc33c7e00},
  {32'hc353a9a8, 32'h43c7ec0a, 32'h42f7d5aa},
  {32'h44827ddb, 32'h431a4063, 32'h416ba284},
  {32'hc4ff5c3d, 32'h43a7029b, 32'h4287077f},
  {32'h448d81a6, 32'h4352c546, 32'h43acabaf},
  {32'hc5025694, 32'h430a455b, 32'hc40d80da},
  {32'h44a3b5d6, 32'hc3813351, 32'h43a7dfc3},
  {32'hc45ad872, 32'h418a7114, 32'h438543f4},
  {32'h43b91ffc, 32'h41f3d18c, 32'h42c44cd8},
  {32'hc51050eb, 32'h43022b9e, 32'h42fe33d3},
  {32'h44ad67e2, 32'h425b5ac3, 32'hc3b6efe7},
  {32'hc39cac8c, 32'h41b03623, 32'h40a805be},
  {32'h4484004e, 32'hc1f12773, 32'h4221faa0},
  {32'hc492e61b, 32'hc204b280, 32'h42a7b53a},
  {32'h44b609a9, 32'hc3d58276, 32'hc2c2b8e4},
  {32'hc494148b, 32'h43c53fc2, 32'hc314bbcd},
  {32'h44f9c444, 32'hc31d176e, 32'hc3956039},
  {32'hc392ad2a, 32'h43def20a, 32'h40c7fdf6},
  {32'h43d7f4ce, 32'hc3580235, 32'hc38f4523},
  {32'hc45a3ffc, 32'h433050d4, 32'h433e32e1},
  {32'h43d500ae, 32'h434d4a8d, 32'h4249e1ff},
  {32'hc4643c28, 32'h4299a215, 32'h432865ff},
  {32'h452a2a9a, 32'h4302fbd4, 32'hc2bfb590},
  {32'hc4849c37, 32'h42cce15b, 32'h4311953f},
  {32'hc2766200, 32'h4241c034, 32'h42e21dcc},
  {32'hc4389cda, 32'h43fe2b11, 32'h4349d112},
  {32'h44f99aa5, 32'hc3160ddc, 32'hc24915bb},
  {32'hc5199ec1, 32'hc3a63536, 32'hc306e2d5},
  {32'h4340699c, 32'hc2c5246e, 32'hc2040fff},
  {32'hc4b74b99, 32'hc2650715, 32'h439ecddd},
  {32'h43fa00fe, 32'h421afeec, 32'hc3a19480},
  {32'hc3f46318, 32'h42e5da72, 32'h4174b4fd},
  {32'h44dbce95, 32'h42ccf8c2, 32'h44031b5d},
  {32'h431f6410, 32'hc3108c49, 32'hc304924f},
  {32'h443c0295, 32'h421c2ba2, 32'hc368a8de},
  {32'hc41d0760, 32'h42e24dcc, 32'h43729b7c},
  {32'h44bce54c, 32'hc340888a, 32'hc2288714},
  {32'hc47ee70d, 32'hc3286a4f, 32'h439eab94},
  {32'h44eb2457, 32'h4318e67e, 32'h438fbdd8},
  {32'hc38d365c, 32'hc34d4515, 32'hc37c28ee},
  {32'h442e6f6a, 32'h435169c5, 32'hc329affd},
  {32'hc4dcfd19, 32'hc38af7f0, 32'hc393dad7},
  {32'h449424fd, 32'hc35df91a, 32'hc40befb0},
  {32'hc499016e, 32'h438fb0e3, 32'h42e07f06},
  {32'h443872b5, 32'h4357ed4c, 32'h43174dc1},
  {32'hc4ec9570, 32'h43aac1e0, 32'h40f2b4c8},
  {32'h44e64a8e, 32'h43075bff, 32'h42f3b62c},
  {32'hc5087775, 32'hc3a5f60a, 32'hc38db62f},
  {32'h43503f50, 32'h4314c241, 32'h4311f7d7},
  {32'h42a59160, 32'h42f20269, 32'h43b19aeb},
  {32'h44d3435a, 32'h40ed6049, 32'hc382b95c},
  {32'hc3951be4, 32'hc16d7463, 32'hc38d79a4},
  {32'h44a41804, 32'hc2c90a95, 32'h427fba34},
  {32'hc43bd8a7, 32'h4370679e, 32'h420afcce},
  {32'h44b01872, 32'hc367663a, 32'hc25ce7ec},
  {32'hc4b04a70, 32'hc329bef9, 32'hc26cbcf4},
  {32'h42460c20, 32'hc3977f6b, 32'hc3adf66f},
  {32'hc5116221, 32'h4346c17b, 32'hc3bcfd38},
  {32'h450b0a36, 32'h43971e95, 32'h436c5c88},
  {32'hc4aa7af6, 32'hc327dbca, 32'hc3666ace},
  {32'h44a08ca0, 32'hc0865f46, 32'h433ee19a},
  {32'hc4f78fcb, 32'h43035ddd, 32'hc22765ae},
  {32'h4504543a, 32'h4314c14b, 32'hc32f6a50},
  {32'hc47a9002, 32'hc0080a46, 32'hc3701810},
  {32'h4523ce10, 32'hc3f5f55e, 32'h42dfd1b6},
  {32'hc4e9b8ba, 32'h435cb17b, 32'h40e8f7f7},
  {32'h44954180, 32'h431e2882, 32'hc0e57910},
  {32'hc4d281ca, 32'hc2d718b6, 32'hc3ae5e04},
  {32'h4521be4d, 32'h42b6bf3e, 32'hc3ccff0f},
  {32'hc49af98a, 32'h4347bd3c, 32'h431a204e},
  {32'h43113320, 32'h42104f7b, 32'h4329f6e7},
  {32'hc47c8197, 32'hc3380f7b, 32'hc2dd7209},
  {32'h451450ba, 32'hc108bd21, 32'hc34cdbc6},
  {32'hc39ebe18, 32'h43009cd9, 32'h42121411},
  {32'h44ccdfb8, 32'hc36763da, 32'hc3a90492},
  {32'hc3c4179c, 32'h4348e278, 32'h41a048cb},
  {32'h44b66d65, 32'h43b991ac, 32'hc2a73ef0},
  {32'hc4606f7a, 32'hc257466f, 32'hc30cda21},
  {32'h43d26680, 32'hc2e3f3f8, 32'hc2fefcf6},
  {32'hc51533fa, 32'hc311a57d, 32'hc35371d4},
  {32'h433a73ec, 32'h4237e9c9, 32'hc2e71658},
  {32'hc42287d0, 32'h43a432b1, 32'hc33bb23f},
  {32'h44ef3bae, 32'hc2102507, 32'h43ac8a91},
  {32'hc4b9d858, 32'hc1c97894, 32'hc3ac94f3},
  {32'h449627d6, 32'hc360b6dc, 32'hc374535a},
  {32'hc4369c37, 32'h43ca7bde, 32'h4366e1db},
  {32'h44efa6d8, 32'hc34a5f83, 32'hc1b2c8fa},
  {32'hc44d8066, 32'h424239c7, 32'h43296aa2},
  {32'h4489159a, 32'hc35e66d6, 32'h430d3d85},
  {32'hc4e44c1b, 32'h42f81476, 32'h42def8f7},
  {32'h44ba3b67, 32'hc17dab41, 32'hc42e01e0},
  {32'hc3baba0e, 32'hc308d0ad, 32'hc36ecb34},
  {32'h444af8ff, 32'h42a60ecb, 32'hc3ac350d},
  {32'hc4c87636, 32'h43c7bd5b, 32'h43873442},
  {32'h45062097, 32'h43aaefce, 32'h41925fc6},
  {32'h3ddd5900, 32'h424a5518, 32'hc3538d5a},
  {32'h42ba9b44, 32'hc34388c3, 32'h42cc0e26},
  {32'hc4d43323, 32'h41ae1376, 32'hc187993e},
  {32'h4508a724, 32'h436ec24a, 32'h43ae79f0},
  {32'hc4ae8644, 32'h41b0973e, 32'h431a968f},
  {32'hc2b14248, 32'h426fee7a, 32'h4341ff64},
  {32'hc4791d74, 32'hc36478c1, 32'hc399bd6e},
  {32'h43e21430, 32'h440ca926, 32'h439d3283},
  {32'hc3d8cfa8, 32'hc3074ba1, 32'h4350ac7e},
  {32'h4512537b, 32'h435a52f4, 32'hc352e9e1},
  {32'hc4f24453, 32'h432b7375, 32'h4288f63e},
  {32'h445b196c, 32'hc3b5255b, 32'h42e17099},
  {32'hc3816244, 32'hc37e74ee, 32'hc2c52fbc},
  {32'h430367e0, 32'hc3c27f04, 32'h435eae58},
  {32'hc3316344, 32'h43e24c8c, 32'h42a6e8dd},
  {32'h43d0b788, 32'hc35e6cd7, 32'h4331b784},
  {32'hc42d4d60, 32'hc3b8249d, 32'h41cce72c},
  {32'h4474ade7, 32'hc2894e73, 32'hc1e71aa2},
  {32'hc5055535, 32'h430543ef, 32'h43316d58},
  {32'h43bc4ce0, 32'h440ba73a, 32'h43eaef9e},
  {32'hc4dac0b6, 32'hc3051e65, 32'h42674dce},
  {32'h4406ae5b, 32'hc1f20e5f, 32'h4310f5b5},
  {32'hc48a00c7, 32'hc385580b, 32'hc2c4774e},
  {32'h4441fb62, 32'hc2775296, 32'h4372e46e},
  {32'h4362fe60, 32'hc3dcf1f0, 32'hc32e3d3f},
  {32'h436e1a68, 32'h4252fded, 32'h44264be0},
  {32'hc40ff8ad, 32'hc11cb46c, 32'hc36a5310},
  {32'h450ad9d2, 32'hc147b3cc, 32'hc3bc5d18},
  {32'hc46ca243, 32'h433c3db0, 32'h433de6d5},
  {32'h44c5a506, 32'h422285e2, 32'h429b2c69},
  {32'hc4a884fc, 32'h43d2a43e, 32'hc3ac9ec7},
  {32'hc39ac834, 32'h4327328e, 32'h42de5014},
  {32'hc509ff80, 32'h433afc03, 32'h42b17ee5},
  {32'h42d7e2a8, 32'hc2e61e60, 32'h4349ff05},
  {32'hc487cc3a, 32'h42d60c3d, 32'hc3a92c2a},
  {32'h451e1ae4, 32'hc371ac54, 32'h43d32742},
  {32'hc5061f5c, 32'hc336f4f5, 32'h422c5111},
  {32'h44feefd3, 32'hc2694f3a, 32'hc02e7d77},
  {32'hc4d2169e, 32'hc2f02826, 32'h4238ac72},
  {32'h44e997dd, 32'h42b7946d, 32'h42692b9c},
  {32'hc490ef57, 32'hc3776d3b, 32'hc3556447},
  {32'h439e0cbc, 32'h40bc569e, 32'h429c5eb7},
  {32'hc50b0195, 32'h43694ecd, 32'h42b73b27},
  {32'h450b82b9, 32'h4301a9b2, 32'hc2cb5373},
  {32'hc4914683, 32'h434b6bbf, 32'hc3edeb95},
  {32'h450d32c7, 32'hc20850ef, 32'h42ca50bb},
  {32'hc493eb72, 32'h436c4042, 32'h433c60cc},
  {32'h44c6f454, 32'h439248b8, 32'hc2f86825},
  {32'hc4900a6d, 32'h43380fc0, 32'hc2e70cb4},
  {32'h448c4862, 32'h4238f2fb, 32'hc328a0e6},
  {32'hc4ac5a1e, 32'h43205301, 32'h4388b1f6},
  {32'h43f05fd8, 32'hc28ad1b9, 32'h42e2f42e},
  {32'hc4473933, 32'hc2f297b3, 32'hc20b7f7d},
  {32'h448cddbf, 32'h43012eee, 32'h43a75524},
  {32'hc4b07f11, 32'h43632206, 32'hbf3acc5e},
  {32'h42dc8b00, 32'hc1e86b51, 32'h43575a18},
  {32'hc4b4f7c9, 32'hc2e4375b, 32'hc228f660},
  {32'h44d4205c, 32'h4115120a, 32'h43792b29},
  {32'hc40da072, 32'hc3b38517, 32'hc304ea56},
  {32'h44b1c4c5, 32'hc29a2043, 32'h41864c2b},
  {32'hc4a2e72e, 32'hc2ab8fab, 32'h3fe97f1e},
  {32'hc4b91312, 32'hc37b80b4, 32'hc3d6208c},
  {32'h44861ee6, 32'hc3823342, 32'h44063e65},
  {32'hc430261c, 32'h4271ed66, 32'h4382c757},
  {32'h445e0ac4, 32'h432cf85f, 32'h440c275d},
  {32'hc4b6d736, 32'hc349cfc9, 32'hc3240db8},
  {32'h4505adcb, 32'hc36c9a29, 32'hc286b579},
  {32'hc3805c08, 32'hc35f8582, 32'hc361af8b},
  {32'h44fd3222, 32'hc1e35edf, 32'h422e2f4b},
  {32'hc436ad44, 32'hc312923a, 32'hc1ca0e37},
  {32'h4508b09e, 32'hc32480dc, 32'hc227e600},
  {32'hc435a978, 32'h418f5ce8, 32'hc3ba7633},
  {32'h44d60a47, 32'hc35c9344, 32'h41a93ec0},
  {32'h42c00736, 32'h42c501d5, 32'hc2cf034f},
  {32'h4308ce5a, 32'h42de5cba, 32'hc3443abc},
  {32'hc4a02f18, 32'hc39dbf25, 32'h42ca451e},
  {32'h44819d03, 32'h432fc76e, 32'hc36f0edb},
  {32'hc4f470d8, 32'h4290d77a, 32'h41e09b77},
  {32'h43e8f644, 32'h4390e4f5, 32'h437bbfae},
  {32'hc5011759, 32'h424f59d4, 32'hc2124d19},
  {32'h422994c0, 32'h439f1c4d, 32'h439b787c},
  {32'hc35ea0c0, 32'h4320ac52, 32'h43174993},
  {32'h44ca1af1, 32'h4388e973, 32'h4409251b},
  {32'hc4e8e43a, 32'hc3c1ee16, 32'hc2a8c0d6},
  {32'h445d8859, 32'h42fbcff8, 32'h4347dbc3},
  {32'hc510b716, 32'h43ae970d, 32'hc2a3b280},
  {32'h4400f5f4, 32'hbfb381a0, 32'hc0a911bc},
  {32'hc515f1f0, 32'h438506bb, 32'h43502698},
  {32'h4461a79b, 32'hc3145b39, 32'hc2551d7a},
  {32'hc4c393a0, 32'h420d6e1a, 32'hc4031cc0},
  {32'h450eeee0, 32'h4301cda2, 32'hc2bc2c5d},
  {32'hc3fdf91a, 32'hc30a1301, 32'hc297ee0c},
  {32'h45046728, 32'h41b42694, 32'hc30bd9ef},
  {32'hc4e406af, 32'h4235805f, 32'h42b68ad0},
  {32'h43df8808, 32'h430cb7d8, 32'h42b2212c},
  {32'hc4c60162, 32'h4389c4c2, 32'h439ebac5},
  {32'h42a87940, 32'hc3470c5e, 32'h3eeabb80},
  {32'hc485e651, 32'hc161a24e, 32'h439b865c},
  {32'h44875bd7, 32'h438b8254, 32'h431fc28c},
  {32'hc4f606c1, 32'h4223ce9b, 32'hc1806d27},
  {32'h44182d7a, 32'h4316b978, 32'hc3152c24},
  {32'hc48ca03a, 32'h43a03a91, 32'h43bbaa2d},
  {32'h449d1bde, 32'h43915f24, 32'h430ee16e},
  {32'hc4dc6e0a, 32'h436ddd3b, 32'h43021384},
  {32'h44ceb221, 32'hc38bd63a, 32'hc20f2c46},
  {32'hc4a1f8c2, 32'hc38936c3, 32'hc2b0ad0a},
  {32'h4503e6f8, 32'h428c4fd7, 32'h434cb86a},
  {32'hc31f8b14, 32'hbfd2c622, 32'h43903887},
  {32'h4435d9f4, 32'hc28c2037, 32'h41ba2b39},
  {32'hc4ba3afa, 32'h422c77f7, 32'hc114ebf5},
  {32'h4506eb2b, 32'hc2576516, 32'h4367114a},
  {32'hc4866945, 32'hc3838def, 32'hc2ea7d7a},
  {32'h436a5c60, 32'h4314ef06, 32'h4113761f},
  {32'hc4d874c7, 32'hc0e0070e, 32'hc3233925},
  {32'h44cc5ca0, 32'h429f9cd8, 32'hc2e093e0},
  {32'hc4faa706, 32'h43292450, 32'hc3013bdb},
  {32'h44ec6935, 32'hc2425f05, 32'h42a0476a},
  {32'hc29dfb81, 32'h43861e52, 32'hc2aa0c10},
  {32'h4515d74c, 32'h43397d7f, 32'hc35bb5ce},
  {32'hc51d5772, 32'hc3797cba, 32'hc24de5af},
  {32'h44a958d8, 32'h439e0355, 32'h41ba0edb},
  {32'hc5194c6e, 32'hc2ead722, 32'hc1b7e3e5},
  {32'h43cce282, 32'h43273806, 32'h42cd8a6a},
  {32'hc50dc75b, 32'hc301dd47, 32'hc3e5e098},
  {32'hc2fe39c8, 32'h4356e399, 32'hc314ed99},
  {32'hc4d2f966, 32'h3f804e12, 32'h4264bbda},
  {32'h450473a0, 32'h4404836a, 32'h41e29aa6},
  {32'hc4ce367a, 32'h437bfcd9, 32'h4360ade3},
  {32'h44b3c6b5, 32'hc38a88ba, 32'hc33615ed},
  {32'hc49d9614, 32'h43e7d73a, 32'hc17e3e63},
  {32'h446927f1, 32'hc2890720, 32'h4347347f},
  {32'hc4c5c6e9, 32'h43ba9bb0, 32'hc2638e60},
  {32'h44a8a962, 32'h43819c07, 32'hc3073d4d},
  {32'hc39e96d0, 32'h428d3ced, 32'h43598300},
  {32'h44d48d0e, 32'h434c3bda, 32'hc14b8ad2},
  {32'hc49475cc, 32'hc326dd5b, 32'hc382b949},
  {32'h44c92bfe, 32'h42505dfe, 32'h4350f468},
  {32'hc41fb226, 32'hc35868b1, 32'hc3801903},
  {32'h450f3ddd, 32'hc3bd8258, 32'hc433a2a0},
  {32'h435c0cde, 32'h41bad16f, 32'h432d12d6},
  {32'h43e98120, 32'hc3aaf5b0, 32'h4213f0f6},
  {32'hc42632f7, 32'hc3cbb39a, 32'hc277eba5},
  {32'h44e72500, 32'hc3dc45fa, 32'h43242c12},
  {32'hc4a350c6, 32'hc3971854, 32'h42c14d87},
  {32'h44d69c3d, 32'h429aa8a9, 32'h434ae227},
  {32'hc49d9042, 32'hc3712f81, 32'h41036a5c},
  {32'hc3b8bff6, 32'hc2c63f45, 32'h434aa574},
  {32'hc40827f9, 32'h436a8346, 32'hc2815489},
  {32'h44a01714, 32'h43180813, 32'hc28e5f86},
  {32'hc41b1e32, 32'h43118a04, 32'h424efd54},
  {32'h446fd890, 32'hc3344222, 32'h43ac503b},
  {32'h414500d0, 32'h4356b789, 32'hc27e36ce},
  {32'h44b8e218, 32'h433b571f, 32'hc3af0443},
  {32'hc3e1742c, 32'h438dfcf7, 32'h42366a35},
  {32'h44f9861e, 32'h43372f28, 32'h432e2fb3},
  {32'hc3955da4, 32'h437cc346, 32'h434a0d41},
  {32'h43c762cc, 32'hc3bfd92d, 32'h44255378},
  {32'hc4ce35f7, 32'h439d2853, 32'hc2b845f1},
  {32'h42dae261, 32'hc3efd1b3, 32'hc1dac26e},
  {32'hc498ee95, 32'h42b9c9d4, 32'hc25d92e6},
  {32'h43ac22c6, 32'hc3974ad8, 32'h43768bac},
  {32'hc4943baf, 32'hc35841ae, 32'h430241a5},
  {32'h44558806, 32'h43b68981, 32'hc36387c1},
  {32'h4391d708, 32'h43266778, 32'h43419894},
  {32'h4431181a, 32'h4339c265, 32'h42b90236},
  {32'hc4d82a80, 32'h43c48706, 32'h428b186f},
  {32'h448cbfef, 32'hc30b176a, 32'h42dcfa5d},
  {32'hc49b3887, 32'h43a1a636, 32'h427355fc},
  {32'h430ddee4, 32'hc3b05049, 32'hc2952c8e},
  {32'hc49b13b8, 32'h432f7e7c, 32'h435df1c2},
  {32'h40025650, 32'hc1f0277e, 32'h43cdf238},
  {32'hc4a9116a, 32'hc24c06ec, 32'hc35427ab},
  {32'h447ebaa7, 32'h43d45bf4, 32'h4354a66d},
  {32'hc4c8556e, 32'h41ec1dd0, 32'hc28abee1},
  {32'h43dfa4ee, 32'h43b4bdde, 32'h42084e7d},
  {32'hc4ff42a0, 32'hc32ed9e0, 32'hc374a40d},
  {32'h44cca906, 32'hc202dc60, 32'hc404234c},
  {32'hc489378c, 32'h419248e5, 32'h43be0bb6},
  {32'h447f6e4b, 32'h4287e700, 32'hc37474b3},
  {32'hc4b1c71e, 32'hc27655c9, 32'h43cf2fdc},
  {32'h44dce990, 32'h4338aa34, 32'hc28bbe14},
  {32'hc49588e5, 32'hc2cda5ad, 32'h41961a27},
  {32'hc3e5af98, 32'hc3844f59, 32'h4384be50},
  {32'hc4a9b9d5, 32'hc23f2434, 32'hc1fa052c},
  {32'h43a1a94d, 32'hc300b47a, 32'hc2fdd845},
  {32'hc469c2d6, 32'hc30bd760, 32'hc30640b1},
  {32'h43bc9fd0, 32'h425e2d1c, 32'h428e1e38},
  {32'hc4d9cd23, 32'h431737c8, 32'h43131850},
  {32'h448dc2d8, 32'hc391b235, 32'h4284aac0},
  {32'hc4c05c39, 32'hc3537188, 32'h43043609},
  {32'h45079b06, 32'h43097134, 32'hc380ca17},
  {32'hc50e5293, 32'hbf263e00, 32'h436dee35},
  {32'h443bab88, 32'h42d333a9, 32'h42e38f9f},
  {32'hc4f79fdc, 32'hc30a2a0a, 32'h4383e336},
  {32'h44ce968f, 32'hc324b85d, 32'hc1bbfc59},
  {32'hc4cc1f8f, 32'hc1889db2, 32'hc30dde0c},
  {32'h44be667d, 32'hc20e179d, 32'h428c2543},
  {32'hc399e014, 32'h419bf109, 32'hc355c0c5},
  {32'h44a1875c, 32'h429e385e, 32'hc3b198bf},
  {32'hc49d83c6, 32'h42f7eaf8, 32'h438dd725},
  {32'h44811909, 32'hc2cc35ba, 32'h431961e7},
  {32'hc4f58a0b, 32'h439d212f, 32'h4357a932},
  {32'h44c60240, 32'h412e7a16, 32'h43d6d0c4},
  {32'hc2b05f94, 32'h4355750c, 32'h42b42094},
  {32'h4490b738, 32'h42a761e8, 32'h4331b2be},
  {32'hc451aaac, 32'h430ab04d, 32'h4277ceaf},
  {32'h448014a9, 32'h43dcabd0, 32'hc3b46823},
  {32'hc4c09859, 32'h425f263f, 32'h43a8cf1e},
  {32'h44e3a014, 32'h438752b4, 32'h44222024},
  {32'hc50bb1fc, 32'hbf5d879e, 32'hc11a10db},
  {32'h43fa1428, 32'hc26736c1, 32'hc27c2b08},
  {32'hc5179ad0, 32'h42ca10bc, 32'h42f01946},
  {32'h44fa512c, 32'hc338c739, 32'h4284f8e5},
  {32'hc49d2dba, 32'h41462b5f, 32'hc1b2f02a},
  {32'h45055c2e, 32'hc3a127c5, 32'hc3ec510e},
  {32'hc4ddb560, 32'h43861962, 32'h43083984},
  {32'h4505dda9, 32'hc3543bc3, 32'h437b172b},
  {32'hc3941140, 32'h41371d2b, 32'h432bd7af},
  {32'h44a700ec, 32'hc3e521a4, 32'hc06be768},
  {32'hc4b7addc, 32'hc2acc7b5, 32'hc24aee40},
  {32'h4414114a, 32'hc39d21a3, 32'h43b9090a},
  {32'hc4e9b6ec, 32'h43425eaa, 32'h437f131a},
  {32'h43ff0828, 32'h426e1d34, 32'hc395be76},
  {32'hc468870f, 32'hc300c546, 32'h424e5fd6},
  {32'h44690608, 32'hc39bf9ff, 32'h41116a48},
  {32'hc2894700, 32'h42d9f98b, 32'hc33a5e5c},
  {32'h450782f6, 32'h42eb60a6, 32'h42af8324},
  {32'hc41724b6, 32'h42e18da1, 32'h43c266c9},
  {32'h42495a29, 32'h43888b53, 32'hc3360029},
  {32'hc4d616a1, 32'hc398b009, 32'hc3302075},
  {32'h44b444ee, 32'h42d4e77e, 32'h433ddee4},
  {32'hc29e75b0, 32'h4388ff1d, 32'hc392cbc2},
  {32'h4449c897, 32'hc23c362d, 32'h43b4ccc1},
  {32'hc31536e4, 32'hc398b606, 32'h440d199e},
  {32'h44acf7b1, 32'h40bce138, 32'hc32d2dca},
  {32'hc447081a, 32'hc1f4ca85, 32'h414b232c},
  {32'h43dcd17a, 32'hc325b198, 32'h434d6cb9},
  {32'hc4c4a4de, 32'h42f07c89, 32'h4389a757},
  {32'h445a6e00, 32'hc381bff7, 32'hc28dbe5c},
  {32'hc495bd57, 32'hc36b894a, 32'hc3a60243},
  {32'h43a74bbc, 32'h435b6ea1, 32'hc32016cc},
  {32'hc3c8f7c8, 32'h410b05f9, 32'hc28c25a9},
  {32'h44403db0, 32'h4173e74e, 32'hc317a643},
  {32'hc4c28a14, 32'hc3ca8e67, 32'hc2851799},
  {32'h43d5279e, 32'h43e88489, 32'h42558318},
  {32'hc4e7a238, 32'hc30c20d3, 32'h42cdc9e2},
  {32'h43e2a9f4, 32'h42cf8ad0, 32'h44060e56},
  {32'hc4c2333a, 32'h424e477a, 32'h42c3d38e},
  {32'h44e43939, 32'hc3fd7ddf, 32'h43d7b0c2},
  {32'hc3aff198, 32'hc34505fc, 32'h433748fc},
  {32'h44901877, 32'h43ecc367, 32'hc3f79aaa},
  {32'hc4f535fe, 32'h43bc9497, 32'hc390306a},
  {32'h44382978, 32'h430d244c, 32'h439ca044},
  {32'hc3838758, 32'hc39ff307, 32'hc3585e59},
  {32'h44d2a8a5, 32'h4298f960, 32'hc08e3b6c},
  {32'hc5063a87, 32'h430889c8, 32'h42e5b174},
  {32'h4520b3ec, 32'h42ab3443, 32'hc30243d5},
  {32'hc4e4edbf, 32'hc419038e, 32'h42f6a226},
  {32'h44b62f10, 32'hc3725be7, 32'hc352e325},
  {32'hc456822c, 32'hc16d6266, 32'h4397aa10},
  {32'h44d4f67a, 32'h43353e18, 32'hc1f4097a},
  {32'hc44852d2, 32'hc40d3c69, 32'h432b34d6},
  {32'hc2b4d1a0, 32'h430a77c6, 32'h4323a333},
  {32'hc3a2d497, 32'h42a5d670, 32'h41fefb57},
  {32'h45062d62, 32'h42f4165d, 32'hc3920a3d},
  {32'hc430ed68, 32'h438fe17a, 32'h422cf118},
  {32'h443a4a60, 32'hc287c33e, 32'h4181a2df},
  {32'hc4fae19c, 32'hc03ff6b6, 32'hc1b43a69},
  {32'h446d9fa2, 32'h4176e673, 32'h431e4188},
  {32'hc4e6fa5c, 32'hc199350c, 32'hc42b34b4},
  {32'h450c15a8, 32'h4360f2c3, 32'hc344c980},
  {32'hc3c75b75, 32'h436d4785, 32'h43b48ed6},
  {32'h4510b668, 32'hc2499af1, 32'hc357e07c},
  {32'hc4fe0a52, 32'h41c3f5ef, 32'hc1835ffc},
  {32'h44dcc1cb, 32'hc399cc28, 32'hc351ea4d},
  {32'hc4b67974, 32'h4333a0e7, 32'h432793ac},
  {32'h446b60b4, 32'hc40360e7, 32'hc3406f68},
  {32'hc460e40e, 32'hc350d7cd, 32'h4277ce55},
  {32'h448abc3e, 32'h442e33cd, 32'h425d8e07},
  {32'hc4521f98, 32'hc2b2497e, 32'hc33962de},
  {32'h44adf529, 32'h416754e4, 32'h4332984c},
  {32'hc40cb9af, 32'h43466521, 32'hc355ae59},
  {32'h4410ea04, 32'hc29b6c04, 32'h425e9c58},
  {32'hc4c6c98e, 32'h425729b8, 32'h42d86aa9},
  {32'h450b8042, 32'hc15040f4, 32'hc432e65b},
  {32'hc4461e7d, 32'hc399479e, 32'h41ac734e},
  {32'h44d98dc1, 32'h424caab8, 32'h41c7c2da},
  {32'hc501f0e0, 32'h43f8a642, 32'h40b07873},
  {32'h450a80da, 32'h41f5764a, 32'h4319b849},
  {32'hc3685558, 32'hc336c0c6, 32'hc1736a52},
  {32'h4401d55e, 32'hc1266bae, 32'hc3460bcb},
  {32'hc42e2628, 32'h42fbdea3, 32'h4332670e},
  {32'h43f3a268, 32'hc303225c, 32'hc3b24299},
  {32'h43220bf4, 32'hc386d01c, 32'hc27b280c},
  {32'h4508a19c, 32'hc3806ab7, 32'hc30dd80e},
  {32'hc32f269c, 32'h4378a71a, 32'hc32fa08a},
  {32'h444be152, 32'h4294fbb4, 32'hc29ae592},
  {32'hc475dcc4, 32'h4239739e, 32'h43836327},
  {32'h448b81ab, 32'h43aa5125, 32'h43701856},
  {32'hc4cc7f9b, 32'h42af7482, 32'h3f43f800},
  {32'h448ea8c1, 32'h418ff878, 32'hc10c685a},
  {32'hc1cf778b, 32'hc23a47b4, 32'h431495de},
  {32'h43d8f390, 32'h425491a1, 32'hc31186fe},
  {32'hc41d8166, 32'hc3a4be83, 32'hc247cc03},
  {32'hc227b700, 32'hc284f741, 32'h439fe04f},
  {32'hc4ae0f64, 32'h433d6381, 32'hc2dff824},
  {32'h44ab64ec, 32'h4399f126, 32'h42e8afc1},
  {32'hc4e11cfd, 32'hc28109bf, 32'h424e4e66},
  {32'h43eae2ec, 32'hc34b3e11, 32'h44009a01},
  {32'hc4ec2d98, 32'hc395f136, 32'h43167004},
  {32'h44d410c3, 32'hc3b2f6b0, 32'hbf3bbda2},
  {32'hc4a9c0df, 32'h43195af9, 32'hc3554bbc},
  {32'h42300f80, 32'hc3ecdafc, 32'hc109c789},
  {32'hc5027780, 32'hc1a403c0, 32'h428b99f9},
  {32'h451373cf, 32'hc1ee62df, 32'hc27ccbfe},
  {32'hc461f7c4, 32'hc27235da, 32'hc35335ad},
  {32'h4450d3dc, 32'hc34c3da8, 32'hc34de976},
  {32'hc4d47b54, 32'hc1904b8c, 32'hc38fcdc5},
  {32'h44f3473a, 32'h4344d9f6, 32'h433d44ce},
  {32'hc4f79c50, 32'h436e3bac, 32'h41a297e2},
  {32'h451b26a1, 32'hc008b8fc, 32'h43240f68},
  {32'hc4a7043b, 32'hc38a2877, 32'hc35708e0},
  {32'h44818fe2, 32'h4246db5a, 32'hc35d4021},
  {32'hc3fc5ac3, 32'h43195c22, 32'hc29bcb23},
  {32'h4513acb1, 32'h42daadd0, 32'hc3bf3cef},
  {32'hc3e2c080, 32'hc36b7b73, 32'h42bb3e5c},
  {32'h450244d2, 32'h41e9a303, 32'h42dfb1f0},
  {32'hc4923609, 32'hc3152840, 32'h419c009b},
  {32'h445c0b30, 32'h42e22e59, 32'h425b006b},
  {32'hc4c499bb, 32'h42620acc, 32'h4202b5b1},
  {32'h45076f1c, 32'hc38f6062, 32'hc31dabea},
  {32'hc31a9940, 32'h429530ea, 32'h4312bfd2},
  {32'h443233a9, 32'hc33f0122, 32'h4312cae6},
  {32'hc4d3df2f, 32'hc309fb0a, 32'hc37a8003},
  {32'h43a4dfd8, 32'h42f7851c, 32'hc332bf1e},
  {32'hc3a1df60, 32'h4371e4e8, 32'hc33d3db8},
  {32'h43037cd8, 32'hc391b5d5, 32'h430caf28},
  {32'hc48017e2, 32'hc2b03dac, 32'hc2263826},
  {32'h44cfb088, 32'h419a7fe0, 32'h43bd2b81},
  {32'hc479234c, 32'hc33f8d59, 32'h4287efd7},
  {32'h4507ea45, 32'hc0c1483c, 32'h41c098b5},
  {32'hc4300386, 32'hc3c19588, 32'h4278e21c},
  {32'h450ebe8c, 32'hc218893e, 32'h4309c5ed},
  {32'hc4d9b130, 32'hc2eeb1da, 32'hc38d305b},
  {32'h4417c4bc, 32'h40ec2fa0, 32'h406eefb8},
  {32'hc4c891d0, 32'h43c9a73d, 32'h436e7f01},
  {32'h4481e7b5, 32'hc3a53852, 32'hc39b8833},
  {32'hc3d9b65e, 32'h42bdf9a6, 32'hc3414364},
  {32'h445de176, 32'hc2f80e1a, 32'h429a1496},
  {32'hc4790d80, 32'hc3076974, 32'hc2b922f0},
  {32'h44aff26d, 32'h42b44cc8, 32'h42c72e1e},
  {32'hc4e44adf, 32'hc205214a, 32'hc37b0695},
  {32'h44bc4cfa, 32'h4331e531, 32'hc28c452d},
  {32'hc3203e50, 32'h437d40c1, 32'h434e2b4a},
  {32'h436b523c, 32'h4432e644, 32'hc3612f27},
  {32'hc476f7ac, 32'hc1d44404, 32'hc3fc1fae},
  {32'h44392d6a, 32'hc3efab89, 32'hc383ac34},
  {32'hc3c6a778, 32'h41cf7515, 32'h4325d582},
  {32'h44bb5529, 32'hc32ba996, 32'h419ba369},
  {32'hc5030caf, 32'h42146971, 32'h43b66cad},
  {32'h4505b140, 32'hc28f5831, 32'h43db7474},
  {32'h4214cfc0, 32'hc37c1c98, 32'h4285854f},
  {32'h44abc2d0, 32'hc308587b, 32'hc3a21ab5},
  {32'hc414f947, 32'h43a828c0, 32'h4328f511},
  {32'h4515dcf5, 32'h42aee1af, 32'hc3299ca2},
  {32'hc515b986, 32'h4339fb79, 32'hc29a9d13},
  {32'h4411b9ba, 32'hc3b949a9, 32'h433847ca},
  {32'hc4aa1745, 32'h4165bea0, 32'h43b80270},
  {32'h4488871c, 32'hc1770f6f, 32'h42feece4},
  {32'hc3d662fc, 32'hc30bb5dd, 32'hc2b015ea},
  {32'h44c6ac42, 32'h432c58dc, 32'h433acc64},
  {32'hc3b30e91, 32'hc328449b, 32'h43b44a2c},
  {32'h449a4da4, 32'h439c3409, 32'hc20d662b},
  {32'hc454ab1a, 32'h4182a4f2, 32'h428ed857},
  {32'h44fb084d, 32'h42bf4750, 32'h439826e6},
  {32'hc34de760, 32'h42fb2f1e, 32'hc3c2bafc},
  {32'h4367d484, 32'hc3594a5e, 32'hc1bd408d},
  {32'hc50d67fe, 32'h429a158d, 32'hbf792fa0},
  {32'h4511f7c6, 32'hc3048572, 32'h4288f60e},
  {32'hc4cab42e, 32'hc284072c, 32'hc269be8f},
  {32'h44aa33b8, 32'hc346da1d, 32'hc3913ac0},
  {32'hc3bec960, 32'h4289de3e, 32'hc35eda3c},
  {32'h4458ac22, 32'h43293fd1, 32'h4290e9c0},
  {32'hc4c39d3d, 32'hc40b3e87, 32'hc335dde2},
  {32'h443be562, 32'hc37400fd, 32'h4301c745},
  {32'hc3051780, 32'hc32bd9b0, 32'hc326fd52},
  {32'h43b8dd04, 32'h43ba5134, 32'hc20b70f8},
  {32'hc385d6c9, 32'h43601771, 32'hc13e91d7},
  {32'h44e88f78, 32'hc36b9585, 32'h421c5dfa},
  {32'hc3168d56, 32'h4226af9e, 32'h44008986},
  {32'h44e5a1a4, 32'hc2bdcb32, 32'h43505ce4},
  {32'hc50cf6fa, 32'hc2eb952f, 32'hc349a841},
  {32'h43e6a06a, 32'hc383af3e, 32'h43a096b4},
  {32'hc4d60aaf, 32'hc20d36e3, 32'hc22cf46c},
  {32'h4502164c, 32'h432b0a72, 32'hc32a9f0f},
  {32'hc4b53f3e, 32'h431387c6, 32'hc23c932b},
  {32'h442804a1, 32'h42b4c3fc, 32'hc2d5b6f0},
  {32'hc4bfd272, 32'h410090b0, 32'hc22e284c},
  {32'h44b4e4e1, 32'hc34598af, 32'hc32cbef8},
  {32'hc42bc5f4, 32'h43556708, 32'hc2930c22},
  {32'h44ecdc29, 32'h43573b87, 32'hc3a14240},
  {32'hc4a0e4e8, 32'hc22ca2e7, 32'h445504ff},
  {32'h44ed8dce, 32'hc30e5c0e, 32'hc39abf19},
  {32'hc5112c10, 32'h429a1b42, 32'h43a1abf4},
  {32'h446d4b4c, 32'h42c1ee1f, 32'hc309acfe},
  {32'hc4b5bc2e, 32'hc37b38d2, 32'hc376d622},
  {32'h43fcf70c, 32'hc1d73b3f, 32'h4240f1b4},
  {32'hc428372e, 32'hc345d834, 32'hc31d99f8},
  {32'h436372f8, 32'h40c2604a, 32'h42fba4c6},
  {32'hc3620550, 32'h43cf044b, 32'hc2d68c76},
  {32'h441ed0b7, 32'hc3bae3c4, 32'hc2ed9f8a},
  {32'hc4aa34c5, 32'h427d9c5c, 32'h42165a9d},
  {32'h44871c02, 32'h42d950e1, 32'hc2bd2bc0},
  {32'h4344e912, 32'hc38016ba, 32'h4177f259},
  {32'h450d281c, 32'hc2a718ca, 32'hc30617f4},
  {32'hc49ba824, 32'hbeedd000, 32'hc2d5389e},
  {32'h4521cddb, 32'h42a1c0a2, 32'h433b61e5},
  {32'h4379af44, 32'h43c430f3, 32'h42be47ef},
  {32'h436dfdfc, 32'hc34bd926, 32'h4370fc8f},
  {32'hc4ac1948, 32'h4284205e, 32'h42c4d460},
  {32'h449c74f4, 32'hc17f952b, 32'hc0bccf1c},
  {32'hc1722400, 32'h42f71634, 32'h439f35c4},
  {32'h44b44bc6, 32'h4381e7cb, 32'h43258782},
  {32'hc4a8e2c8, 32'h4255eb28, 32'h42a2cd2f},
  {32'h44471845, 32'h42880974, 32'hc34d2afd},
  {32'hc4ac693e, 32'hc34b2499, 32'h42d2fca9},
  {32'h448f7b32, 32'h4183edf9, 32'hc37159f5},
  {32'h4199c000, 32'h42ddf7b0, 32'hc317773f},
  {32'h45030cab, 32'hc2134d1a, 32'hc4264f95},
  {32'hc517ddd3, 32'hc18402ca, 32'h411cdcaa},
  {32'h451b5fd5, 32'h422ab9ae, 32'h434e4b58},
  {32'hc500b7bb, 32'hc32ea83d, 32'h42dfd582},
  {32'h44c9d61c, 32'h430d2f0a, 32'hc3bb352d},
  {32'hc49ec7da, 32'h43987c7c, 32'h43939d57},
  {32'h44aaa09e, 32'hc39c9e3e, 32'hc1a9f984},
  {32'hc4a876e8, 32'hc231ed08, 32'hc2679241},
  {32'h44cd01f2, 32'hc3831fe1, 32'h422d9667},
  {32'hc481d393, 32'hc2b1a848, 32'hc2a45934},
  {32'h4519957a, 32'h4393dd18, 32'hc363ea37},
  {32'hc4dfc1f9, 32'hc214c2cd, 32'hc00d2c3c},
  {32'h44f86793, 32'h42c78816, 32'h42f986d9},
  {32'hc4c62906, 32'hc31c4d5a, 32'hc3c3cf59},
  {32'h44390d2c, 32'hc25e2002, 32'hc346b040},
  {32'hc4728ff2, 32'h439c14ab, 32'h43fb2628},
  {32'h4513b32f, 32'h437ae1a2, 32'hc2d461ef},
  {32'hc27601ba, 32'h43872742, 32'hc2a65504},
  {32'h44cd8f4e, 32'hc352b7a2, 32'h4226ee51},
  {32'hc3eab39c, 32'h41970f80, 32'hc385c997},
  {32'h44c5d5ae, 32'hc3345be3, 32'h42bda012},
  {32'hc379dfe2, 32'hc317ab9d, 32'h43e11061},
  {32'h4423d8ea, 32'h42b014f0, 32'hc384e96f},
  {32'hc4b40fbc, 32'h439380ab, 32'hc110d6d9},
  {32'h44bdeb92, 32'hc3e84dda, 32'hc3776de4},
  {32'hc4621264, 32'hc2d20d4d, 32'hc2383cdc},
  {32'h4514572a, 32'hc2acb86c, 32'hc16b9764},
  {32'hc4bc5998, 32'hc280facd, 32'hc3959948},
  {32'h44f85dd3, 32'h436ed6b1, 32'h4350df25},
  {32'hc5099dae, 32'h41194478, 32'hc3264749},
  {32'h45033f61, 32'h42609e5a, 32'h439eae5b},
  {32'hc47d61f4, 32'h423b2c45, 32'h42299783},
  {32'h43d5a85a, 32'hc234abc4, 32'hc3e05b90},
  {32'hc4a9b6e8, 32'hc233a918, 32'h41d24b7e},
  {32'h450f1a41, 32'hc36a1b52, 32'hc2f898c6},
  {32'hc497f4eb, 32'hc37556a5, 32'hc3ca3daa},
  {32'h443b8e49, 32'hc284c337, 32'hc2ccb193},
  {32'hc4d74c2d, 32'h4374ec90, 32'hc36b31b4},
  {32'h44a0c30b, 32'hc3a10039, 32'h43389cf6},
  {32'hc3946a0a, 32'h434d5c96, 32'h418e4dd5},
  {32'h44907790, 32'hc2d6f554, 32'hc3e0f34f},
  {32'hc4fa1dd8, 32'h4201bd1b, 32'h435fa7fc},
  {32'h440f274a, 32'h43d9274c, 32'hc32f487d},
  {32'hc4c1b687, 32'hc18454ef, 32'hc333022a},
  {32'h44eadf73, 32'hc33699a5, 32'h4270b324},
  {32'hc34fc570, 32'hc298f9fb, 32'h43fd6ed3},
  {32'h446c9166, 32'hc2bfed03, 32'hc2d079c7},
  {32'hc5130f80, 32'h43d87e6f, 32'h43d1357a},
  {32'h448242c2, 32'hc3939b01, 32'hc306c54e},
  {32'hc41e7708, 32'hc14b65e2, 32'h440222bb},
  {32'h443c90b0, 32'h421430f1, 32'hc3964567},
  {32'hc4bacbe0, 32'hc4011978, 32'h42baea05},
  {32'h44083eba, 32'hc3f3d4cf, 32'h4249af1a},
  {32'hc4e6365f, 32'hc36c3682, 32'hc15c4853},
  {32'h44fb28bf, 32'hc2ff1d23, 32'h41c089a1},
  {32'hc4e2d707, 32'h41eea9ef, 32'h4213fb8d},
  {32'h44e4ff66, 32'h43285a58, 32'h43b36c6f},
  {32'hc4d2d01a, 32'hc249bf83, 32'h43987a5e},
  {32'h431c4c10, 32'hc28cdf33, 32'h426c4669},
  {32'hc44b00d9, 32'h43e2a907, 32'hc316c46a},
  {32'h43fa652d, 32'hc3e873ae, 32'hc2babb36},
  {32'hc293eb70, 32'h43c8f46c, 32'h43d8ae97},
  {32'h44aa8791, 32'hc253c5d9, 32'h407bd464},
  {32'hc36b0bd0, 32'hc0d661ac, 32'h433b384c},
  {32'h44e4c1e0, 32'h42b8aa0a, 32'h431a58b9},
  {32'h44c145f1, 32'hc36888e5, 32'hc3daaf94},
  {32'hc4e9b8ba, 32'h43924fa6, 32'hc3c191de},
  {32'h448008f8, 32'h439e1bec, 32'h439aaf7a},
  {32'hc4f72998, 32'h433c05dc, 32'hc23124fd},
  {32'h44e2dc65, 32'h43c5a61f, 32'h437e6b8f},
  {32'hc4c8231a, 32'h423793b0, 32'h429f934f},
  {32'h43c71eb3, 32'h425cb0ab, 32'hc3c935d2},
  {32'hc43bb280, 32'h438f131c, 32'h41ee425b},
  {32'h4496b2d0, 32'h426cfd80, 32'hbdb6218d},
  {32'hc310499d, 32'h43011c46, 32'hc3a3eae1},
  {32'h4463588a, 32'hc3a55920, 32'hc3667cc9},
  {32'hc504de8b, 32'hc09aacf9, 32'h4386dd98},
  {32'h44f40e37, 32'hc1e6a59b, 32'h41b3d65b},
  {32'hc525f27a, 32'hc3e594da, 32'h43b3d918},
  {32'h44f491e0, 32'hc290b6ca, 32'hc12b7d38},
  {32'hc39b71cc, 32'h43b2bd63, 32'h4230a088},
  {32'h44c4f944, 32'h42ace6ac, 32'h4177c511},
  {32'hc4f78fd1, 32'hc30d9309, 32'hc330fa1b},
  {32'h44978578, 32'hc39ac53f, 32'hc280d083},
  {32'hc45df7ca, 32'h424e9518, 32'hc395d570},
  {32'h44d55f0c, 32'hc100d721, 32'h4332abf2},
  {32'hc4c5bfe8, 32'h409bfceb, 32'h418bd995},
  {32'h45164fa3, 32'hc29b4cba, 32'hc32e84e9},
  {32'hc42c0c02, 32'hc23b2b52, 32'hc22f7fb8},
  {32'h44858a27, 32'hc3515d87, 32'hc308073b},
  {32'hc4e370b3, 32'h421963af, 32'h433e7a99},
  {32'h4505af09, 32'hc34646dd, 32'h433fd7e5},
  {32'hc4d61608, 32'h436d69f4, 32'hc30c82e5},
  {32'h44eeabe8, 32'h4327f0ae, 32'h42a7c639},
  {32'hc5068319, 32'h42e906e0, 32'h419dc4d6},
  {32'h4416a291, 32'hc20d6ec1, 32'h42cd449c},
  {32'hc4c96914, 32'hc3669b0e, 32'h430d9739},
  {32'h44e8acf5, 32'hc38aaf0a, 32'h42a23630},
  {32'hc49e0c4c, 32'hc3921a82, 32'h42986d53},
  {32'h44d974a5, 32'hc2fa3ba5, 32'hc367a199},
  {32'hc33378be, 32'hc36f5703, 32'h43488364},
  {32'h449b0fe0, 32'hc3742e41, 32'h3ff8ac55},
  {32'hc4458674, 32'hc1c47b31, 32'h439cbd8b},
  {32'h4438e76c, 32'h430793d7, 32'hc3883c43},
  {32'hc39c61da, 32'h4347e35f, 32'h41300017},
  {32'h45085f79, 32'hc38dc5d9, 32'h43d040f6},
  {32'hc512c7ee, 32'h429ec6cc, 32'hc3871e04},
  {32'h44ec3b2b, 32'hc3809b8c, 32'h4314274c},
  {32'hc50c261e, 32'hc3442948, 32'h433c5f7d},
  {32'h448c7664, 32'hc365570b, 32'h431089bd},
  {32'hc4b1a4fa, 32'h43803479, 32'hc3681b8a},
  {32'h450789f7, 32'h438191cc, 32'h41fce8a3},
  {32'hc4e4af12, 32'hc379d6d9, 32'h42979dcb},
  {32'h4500abe1, 32'hc3440edc, 32'hc2bf0758},
  {32'hc4b22977, 32'h430102ca, 32'h421183b8},
  {32'h45151ba9, 32'h438fd386, 32'hc2bf16f2},
  {32'hc4a835da, 32'hc31411ec, 32'hc3117008},
  {32'h44e094e7, 32'hc2da321f, 32'hc3c1a2bf},
  {32'hc4179e4b, 32'h42f1ecf9, 32'h4213bf6f},
  {32'h43915082, 32'hc375ea21, 32'hc24b1d10},
  {32'hc398c018, 32'hc39b5417, 32'h42dfbef2},
  {32'h44a14a22, 32'h434c851c, 32'hc361199c},
  {32'hc31ad700, 32'h43be83c1, 32'hc329432e},
  {32'h44efcb92, 32'h4252abe3, 32'h41e6a20b},
  {32'hc46f324b, 32'h42629e76, 32'hc298be68},
  {32'h44923490, 32'h42e5cc6a, 32'hc2625026},
  {32'hc4343b2f, 32'h436e7270, 32'h422c8324},
  {32'h451085d3, 32'hc39eec42, 32'hc2d93b28},
  {32'hc424d1a4, 32'hc2a4cdba, 32'h432b72bc},
  {32'h44fc3e7a, 32'h43319433, 32'h42859cec},
  {32'hc501eb5e, 32'hc3c224e2, 32'h43c0376f},
  {32'h43df7050, 32'hc250a119, 32'h429b3a82},
  {32'hc449a61f, 32'h40e96ea9, 32'h42c5ce1f},
  {32'h44ad2c13, 32'hc27024e6, 32'h4269d2e1},
  {32'hc49ab031, 32'hc3f50b7a, 32'hc31ce7ee},
  {32'h45096e6b, 32'hc134a708, 32'h42f1d96d},
  {32'hc3b76598, 32'hc2715151, 32'h407589cd},
  {32'h450b83dd, 32'h40159e1f, 32'hc218f832},
  {32'hc470950c, 32'h43141ac7, 32'h41677a6c},
  {32'h4494f9ec, 32'hc1d655f5, 32'hc3581cf5},
  {32'hc397fcc8, 32'h436ccb07, 32'hc2005080},
  {32'h44e10ad8, 32'h42df42cb, 32'hc14589bf},
  {32'hc50f2365, 32'h42fd8ddf, 32'h4319c4f1},
  {32'h45176f76, 32'hc35b0fdd, 32'h4406030f},
  {32'hc1ab7a50, 32'hc388cb62, 32'hc350dc9b},
  {32'h45118676, 32'hc31e7b63, 32'hc2c39080},
  {32'hc5190efa, 32'hc31f7f6b, 32'hc25ca35a},
  {32'h4463feeb, 32'h43ae8ed2, 32'hc3b130f2},
  {32'hc4b61b18, 32'h416a6726, 32'h4386df16},
  {32'h45039351, 32'hc1bbd6d7, 32'hc34473d4},
  {32'hc4d7317d, 32'hc38e3d8b, 32'h42c0e9c8},
  {32'h4450ecba, 32'h428af78a, 32'h42b723af},
  {32'hc46b4532, 32'h4260b83d, 32'h42643d5e},
  {32'h439f53a2, 32'hc30dbba6, 32'hc317c7b0},
  {32'hc501c1b5, 32'h421e19d3, 32'hc2ac2320},
  {32'h44ccfc42, 32'h43bfae2c, 32'hc3d8467e},
  {32'hc40e3867, 32'hc377a4e7, 32'hc23371d6},
  {32'h439f08cc, 32'hc31d1024, 32'hc38a972f},
  {32'hc4c48296, 32'h4281bff3, 32'hc2199f20},
  {32'h4505514f, 32'hc3be76e4, 32'hc2fc1349},
  {32'hc4f33814, 32'h4251d470, 32'h41313274},
  {32'h4490435c, 32'h4282b388, 32'h4393ca68},
  {32'hc4ffa33d, 32'h42c8ab1a, 32'h431f766e},
  {32'h44ebad18, 32'h4260e161, 32'h43140d29},
  {32'hc4b4dd39, 32'h42ba0c18, 32'hc38825e1},
  {32'h431196b0, 32'hc324028b, 32'h42101813},
  {32'hc473eda8, 32'hc2e6f800, 32'h438e0570},
  {32'h44712e3b, 32'h43ad3bae, 32'hc34d2ee2},
  {32'hc4451742, 32'h436fe4d6, 32'h4304f94e},
  {32'h43c1f77c, 32'h430ac1a9, 32'hc2a027b0},
  {32'hc4a59216, 32'hc3c953a1, 32'h432f1f59},
  {32'h450df271, 32'hc2f5c29d, 32'hc406899d},
  {32'hc437cd2c, 32'hc4000df6, 32'h435f33c7},
  {32'h44e51ab8, 32'h43e44703, 32'hc3150ff6},
  {32'hc4717558, 32'h43143f13, 32'h4355cfc7},
  {32'h43ddab45, 32'hc3448cf1, 32'hc2fc57f6},
  {32'hc3a00df8, 32'hc217cb9e, 32'h4330e2bc},
  {32'h45093e14, 32'hc2b5db0e, 32'h43bbdfa4},
  {32'hc46dc464, 32'h43a4307a, 32'h432fa551},
  {32'h44251e99, 32'h42e9f305, 32'h42e1ec69},
  {32'h4084a000, 32'h4300f406, 32'h43005044},
  {32'h4503e070, 32'hc386f5e4, 32'hc1432fe4},
  {32'hc47ac981, 32'h43332d62, 32'hc26604d0},
  {32'h44928f46, 32'h436c995b, 32'h4119ad7c},
  {32'hc4febf2d, 32'h436cbe40, 32'h43b1aabf},
  {32'h44e76a74, 32'hc32c9b2a, 32'h43c78b4f},
  {32'hc43f0ba6, 32'hc2b95aa0, 32'hc30d6d41},
  {32'h44f3a217, 32'hc3375000, 32'h42d4a0c2},
  {32'hc462085a, 32'hc28d90ee, 32'hc3094e28},
  {32'h44bae336, 32'hc288cb9a, 32'h43d86abb},
  {32'hc2d08a53, 32'h43443534, 32'hc3420502},
  {32'h4502aa1b, 32'hc4050bde, 32'h4395ad2f},
  {32'hc48646bd, 32'h42ced8f5, 32'hc2a000d0},
  {32'h44e15856, 32'h43e698f7, 32'hc25cff51},
  {32'hc4af2efa, 32'h44074918, 32'h43b3c96e},
  {32'h44a1a7a5, 32'h3fb269b8, 32'h430e3803},
  {32'hc4d7a85e, 32'h438ffb88, 32'hc31b92b3},
  {32'h447718c0, 32'hc2266288, 32'h43a044a6},
  {32'hc4b09c53, 32'h426ba9a8, 32'h436a966e},
  {32'h44d0be30, 32'hc1c38d83, 32'h42edd3d7},
  {32'hc4f98acb, 32'hc34366d3, 32'hc13efa5e},
  {32'h4516e28d, 32'h435b7a9d, 32'h4122678e},
  {32'hc509a348, 32'hc3d01fb6, 32'h436c2811},
  {32'h43e199a0, 32'h43cf7f85, 32'h435e3417},
  {32'hc46c0953, 32'hc1b04531, 32'h4181026e},
  {32'h44837f39, 32'h4221fcd1, 32'h4345bd18},
  {32'hc4bae880, 32'h41bfe6ba, 32'h428d1165},
  {32'h44f2f772, 32'hc35412d0, 32'h42ee7908},
  {32'hc4dfe409, 32'h4262c599, 32'hc24fe226},
  {32'h44e08131, 32'h426584a1, 32'h4344fbcc},
  {32'hc48c0f76, 32'hc2f5eddd, 32'h4328beaa},
  {32'h44a6cf43, 32'h42dc0883, 32'hc310d79b},
  {32'hc439ad58, 32'hc332a3fa, 32'hc0b42910},
  {32'h44bf83a7, 32'h433301f8, 32'hc25cb31c},
  {32'hc4dc2024, 32'hc370de33, 32'hc3962188},
  {32'h4503697f, 32'h40ba023a, 32'h42c80c2a},
  {32'hc4d7b491, 32'hc1c104c4, 32'hc317b7bb},
  {32'h4043ed80, 32'hc31fdb62, 32'hc408eb4f},
  {32'hc3f4b3a6, 32'hc31511b7, 32'h436de5b4},
  {32'h4512e264, 32'h4288374a, 32'hc39351d1},
  {32'hc35fd790, 32'hc32a060a, 32'h422bc7ea},
  {32'h4499021a, 32'hc34c225b, 32'h426e9262},
  {32'hc3ec7bf4, 32'hc1444ed8, 32'hc3c90163},
  {32'h4524cc88, 32'h421fafad, 32'h424957bb},
  {32'hc49eeb26, 32'h433056f6, 32'h437f5871},
  {32'h44ba0fac, 32'hc3755433, 32'hc283245e},
  {32'hc4e6b32a, 32'hc2c5d020, 32'h42387a7c},
  {32'h43a5be84, 32'h42237ab4, 32'hc28216e7},
  {32'hc4214ebf, 32'h43499f60, 32'hc3199704},
  {32'h44f97668, 32'h4307dc8d, 32'h42b84aba},
  {32'hc38bb388, 32'hc305525f, 32'hc37f379a},
  {32'h44c6df68, 32'h418017cc, 32'h4233c903},
  {32'hc3ec447c, 32'hbf692efa, 32'hc1c844b8},
  {32'h44f5fac6, 32'hc25e9cc6, 32'h43158c7d},
  {32'hc4efaf28, 32'hc3837580, 32'h4234a8e4},
  {32'h44180382, 32'h43cbec94, 32'hc2891924},
  {32'hc4b2b43a, 32'hc397e794, 32'h42edc558},
  {32'h43241cf0, 32'hc28918ee, 32'h4115c1b7},
  {32'hc450e0ae, 32'h438f060e, 32'hc30fef29},
  {32'h43691b20, 32'hc433a31f, 32'hc334bb2f},
  {32'hc4a92bfb, 32'hc3962897, 32'hc2f00dda},
  {32'h44d97dd5, 32'h41ea7f3a, 32'hc1b1f60d},
  {32'hc49443ab, 32'hc325f1e3, 32'h434ccc36},
  {32'h44355adc, 32'h425539e8, 32'h43542bd4},
  {32'hc47251d7, 32'hc383d977, 32'h43a1086d},
  {32'h44b6594b, 32'h434fe1a9, 32'hc1ba694f},
  {32'hc4e76015, 32'hc368c758, 32'h43932f1a},
  {32'h44c2d71c, 32'h42b375f0, 32'h4298b625},
  {32'hc5045329, 32'h41fa5c22, 32'hc37c154d},
  {32'h445aaa48, 32'hc1cf8b24, 32'hc2a213c9},
  {32'hc461b75d, 32'hc1a76ce1, 32'h43616927},
  {32'h44f63258, 32'hc3846cb6, 32'h4364d0df},
  {32'hc4efb25d, 32'hc3392259, 32'hc31bc103},
  {32'h446371ab, 32'h42eb311d, 32'h41dc40c2},
  {32'hc4e1fe39, 32'hc378e6a8, 32'hc23a17cc},
  {32'h447cdc74, 32'hc20be265, 32'h43b0ef66},
  {32'hc4ad0a84, 32'h435a32f2, 32'hc1a87fde},
  {32'h4408d8c5, 32'h429e0d2e, 32'hc39c9a98},
  {32'hc3b80938, 32'hc0ffa106, 32'h423323b0},
  {32'h44e3d584, 32'hc30912e2, 32'h41603130},
  {32'hc3ea0ac5, 32'hc3236496, 32'h43dd4497},
  {32'h4447adbb, 32'hc2875ad1, 32'hc10ae789},
  {32'hc4141148, 32'hc2a6b44e, 32'h4230a016},
  {32'h430c2a38, 32'h4331af10, 32'h439927a6},
  {32'hc4b172de, 32'hc28a9cc6, 32'h4337f42e},
  {32'h44f084ee, 32'h43477e7d, 32'h432f592a},
  {32'hc4f7aba8, 32'h43725055, 32'hc1a25b81},
  {32'h4392152d, 32'hc2cb54a3, 32'h43190b47},
  {32'hc4d138c8, 32'hc1c0896b, 32'hc209a7e2},
  {32'h439f608c, 32'h4272d9b7, 32'hc3118b42},
  {32'hc3f88318, 32'hc2a05ba0, 32'h4392536e},
  {32'h44d3e60b, 32'h4402ad05, 32'h4296b227},
  {32'hc305cee0, 32'hc2732cd8, 32'h3f443c50},
  {32'h44916e08, 32'h433fe1c1, 32'h42d58c78},
  {32'hc392a22b, 32'hc3135759, 32'hc3b0c153},
  {32'h4480e876, 32'h43a8153c, 32'hc2da303a},
  {32'hc40c71e3, 32'hc2b7b45a, 32'hc3164e7d},
  {32'h44873413, 32'hc28055f3, 32'h43231368},
  {32'hc4716282, 32'hc385d00a, 32'hc2ce11a5},
  {32'h44b588ed, 32'hc311b91f, 32'h4269e68a},
  {32'hc4e32c1e, 32'hc29a1f99, 32'hc39894eb},
  {32'h450e9f8d, 32'h43b63426, 32'h42cff313},
  {32'hc46c9db6, 32'hc322238d, 32'h434322ca},
  {32'h44132d8a, 32'hc33a8543, 32'hc2d96a2d},
  {32'hc4ec4d07, 32'hc2956bdb, 32'h42dd6b36},
  {32'h447365c6, 32'hc1ae722a, 32'h4154873d},
  {32'h43075420, 32'hc27b3852, 32'h439936bd},
  {32'h43d42a25, 32'h429ac56e, 32'h42a10c3d},
  {32'hc3bb4374, 32'h43cd73c9, 32'hc2a95073},
  {32'h44839bab, 32'hc2b8259e, 32'hc3bd07f3},
  {32'hc500fb6a, 32'h43e5ec86, 32'hc341d121},
  {32'h448e71ec, 32'hc17aac01, 32'hc30bac03},
  {32'hc505082f, 32'h4338f4a1, 32'h4234b9ba},
  {32'h4510c0f5, 32'hc369c821, 32'h424c86ae},
  {32'hc4a15eca, 32'hc3b2eb6c, 32'hc2cdaf41},
  {32'h4502e49d, 32'h41e901b6, 32'hc2f76ca7},
  {32'hc4e132f2, 32'h43949dbe, 32'hc2a87b20},
  {32'h44bc88fe, 32'h43393bf3, 32'hc2f32955},
  {32'hc480e359, 32'hc2fda641, 32'h42962582},
  {32'h43fa7f10, 32'h42fa4ea2, 32'h4324a34a},
  {32'hc38928d0, 32'h42802a77, 32'hc1fe904e},
  {32'h44ad2d98, 32'h43abbc47, 32'hc37cfc4f},
  {32'hc157ce88, 32'hc35488ce, 32'h439e9583},
  {32'h451102fc, 32'h436fe3b7, 32'h40a9a908},
  {32'hc49dc1fb, 32'hc206f146, 32'hc24f7a6a},
  {32'h45000713, 32'h42e33169, 32'h4331d379},
  {32'hc508ee48, 32'hc1987434, 32'hc3726305},
  {32'h4403f72c, 32'h428f39eb, 32'h42e41c36},
  {32'hc4b43ae8, 32'h4102b0bd, 32'h4352562d},
  {32'h450eae69, 32'hc1de83ec, 32'h43997d79},
  {32'hc4ddaaaa, 32'hc3c4c27b, 32'hc2c00ddd},
  {32'h44e44466, 32'h4356f6e3, 32'hc3a07a8a},
  {32'hc2689c80, 32'hc3782982, 32'h422c88e4},
  {32'h43843e34, 32'h42bbe0d5, 32'hc3a8783c},
  {32'hc3bded2a, 32'hc327a614, 32'hc386fa70},
  {32'h447a953b, 32'h439bac16, 32'hc30640eb},
  {32'hc460a4c8, 32'hc3b1f13c, 32'h4194dcf0},
  {32'h401a5df8, 32'hc4170c5b, 32'hc2b0ec2c},
  {32'hc30d58c6, 32'h43f2a7e0, 32'hc33aa555},
  {32'h44b7400f, 32'hc3aab209, 32'h434f6976},
  {32'hc4bb6d93, 32'hc2a712d3, 32'hc197cd40},
  {32'h42894f5e, 32'hc369495c, 32'h432a4100},
  {32'hc4fff6e9, 32'hc2d25bac, 32'h4315206c},
  {32'h44a71b63, 32'hc2c326aa, 32'h42cc5b17},
  {32'hc489a3ea, 32'h4333c960, 32'h4390118c},
  {32'h44c5555a, 32'hc30e98db, 32'hc2cbf320},
  {32'hc4f2cc87, 32'h4310d53b, 32'h43910595},
  {32'h44409e8e, 32'hc3915952, 32'hc29f2fa0},
  {32'hc50914fb, 32'h4413329c, 32'h431ca448},
  {32'h44270cb2, 32'hc3ac3f79, 32'h43df3a3f},
  {32'hc445d08a, 32'hc31b0364, 32'h429bd94d},
  {32'h44f753c8, 32'h43a354a2, 32'h429f6cc6},
  {32'hc4722739, 32'h432fa002, 32'hc3d6fb27},
  {32'h450aac06, 32'hc2f60c8e, 32'hc384aa5e},
  {32'hc4956fa1, 32'h4366542a, 32'hc0579e50},
  {32'h45015865, 32'hc3444126, 32'h4283d348},
  {32'hc2f9657c, 32'hc269365c, 32'hc316b5fd},
  {32'h440e5d54, 32'hc317075b, 32'hc3995da6},
  {32'hc1521009, 32'h43354da8, 32'hc2b398ae},
  {32'h43f7d61e, 32'h43a3f7ca, 32'hc3a04c87},
  {32'hc47277d6, 32'hc3a96415, 32'hc3986c0d},
  {32'h44b5ab5a, 32'hc2cf30d3, 32'h42d72287},
  {32'hc45e1745, 32'hc380e85f, 32'h42166626},
  {32'h449eacd1, 32'h4291b103, 32'hc38837a3},
  {32'hc4e4a3fd, 32'h433da44d, 32'hc2906534},
  {32'h44907914, 32'hc2bfdbfc, 32'h40c7de4d},
  {32'hc504d779, 32'hc2eb1dcb, 32'h43c41588},
  {32'h44a94b8d, 32'hc39e421b, 32'h439ca1f7},
  {32'hc414a1bb, 32'hc23e8aa1, 32'hc18a6a74},
  {32'h4486a022, 32'h42d069fb, 32'h43c439ca},
  {32'hc40d1126, 32'hc2427cb1, 32'h432ad1a0},
  {32'h45260164, 32'h42e84103, 32'h42f5029d},
  {32'hc4c8f7fb, 32'hc3a8bee6, 32'h42e5ab6c},
  {32'h4507b314, 32'h43414a25, 32'hc382db14},
  {32'hc4a75aa7, 32'h4307192f, 32'hc293544d},
  {32'hc2debd50, 32'hc388c5bc, 32'hc40115f4},
  {32'hc47e9bfe, 32'h43fe94ce, 32'h442ee842},
  {32'h4511cf48, 32'h4391285c, 32'hc31c33fd},
  {32'hc4d78d86, 32'h421a48d9, 32'h43651e87},
  {32'h43747144, 32'hc2378382, 32'hc404807f},
  {32'hc4b0b971, 32'hc2fa988f, 32'h43180c00},
  {32'h43a98060, 32'hc2c46233, 32'h43115b16},
  {32'hc4c2395c, 32'h438db164, 32'hc3546a04},
  {32'h45182843, 32'h4262a27f, 32'h438d1402},
  {32'hc4970dbe, 32'h43a80f6f, 32'hc37ec61f},
  {32'h44cba950, 32'hc3baf09e, 32'hc3a86789},
  {32'hc497545c, 32'h43aa5492, 32'h43321b48},
  {32'h45186a2f, 32'h429de3db, 32'hc2653a92},
  {32'hc4e8980a, 32'hc43c1d3a, 32'h43887b50},
  {32'h44430b18, 32'hc2e40441, 32'hc31643bb},
  {32'hc5177cb7, 32'h41a41d77, 32'h4354b834},
  {32'h431cbd30, 32'h432e21a8, 32'h42513445},
  {32'hc431e77e, 32'hc380556f, 32'h43df03eb},
  {32'h450e79bb, 32'h43b605da, 32'hc1b8bc72},
  {32'hc0f54600, 32'h42939a52, 32'h4360c7dc},
  {32'h449d34ea, 32'hc2f89718, 32'h43a9e1b2},
  {32'hc3532828, 32'hc3da4dbb, 32'hc37c478e},
  {32'h45116f35, 32'hc38d334c, 32'h42f17c8b},
  {32'hc500ff3b, 32'h427a2b06, 32'hc0c6329b},
  {32'h44ab5312, 32'hc3ad834e, 32'hc214f13d},
  {32'hc50091ef, 32'h421a0575, 32'hc31b5833},
  {32'h4483ebc6, 32'hc1da3581, 32'hc1239f10},
  {32'hc46cf658, 32'h4317e1ef, 32'h432358d1},
  {32'h44463d3a, 32'h433c2efe, 32'h43e314ac},
  {32'hc4982424, 32'h4313ac25, 32'hc3408c0f},
  {32'h425b0630, 32'h4301651f, 32'hc3a6e80a},
  {32'hc517f18c, 32'hc1c14e28, 32'hc317e782},
  {32'h4484a63a, 32'h4218f40c, 32'hc35749ba},
  {32'hc4d5226c, 32'hc1bcff22, 32'h41dd90f9},
  {32'h450a3d94, 32'hc2873a04, 32'hc2f46229},
  {32'hc3914b48, 32'h430cc165, 32'hc33f4099},
  {32'h44a14b6a, 32'h4291c201, 32'h414d83e2},
  {32'hc3ebceeb, 32'h419c96e8, 32'hc283552e},
  {32'h4424048b, 32'hc2c019cb, 32'h43629aba},
  {32'hc504cac9, 32'hc3024bb3, 32'h42ed3c96},
  {32'h44b52c53, 32'hc15e9430, 32'h43151053},
  {32'hc3f2961c, 32'hc2c75d3b, 32'h43892610},
  {32'h43a041a4, 32'hc337bb12, 32'hc342cfda},
  {32'hc43faac0, 32'hc25a2584, 32'h426bf380},
  {32'h448256ee, 32'h4350accf, 32'h430c92ef},
  {32'hc4c9913e, 32'hc36ba348, 32'hc3133bfe},
  {32'h451af1c8, 32'hc3ab427b, 32'hc1e600f9},
  {32'hc45d2d60, 32'h42a56181, 32'hc2b6a1fc},
  {32'h45117b98, 32'h433a7898, 32'h4299c001},
  {32'hc4110d3e, 32'h4316b91c, 32'hc185a758},
  {32'h447ecc06, 32'h441f71aa, 32'h42fe7247},
  {32'hc3623190, 32'h42fe5757, 32'hc4170edd},
  {32'h45194487, 32'h4222e225, 32'h43dafd64},
  {32'hc5112a3c, 32'hc3d1ff1f, 32'hc2862640},
  {32'h43c04cd8, 32'hc3ee4c82, 32'hc19b9fc0},
  {32'hc4669954, 32'h439426d6, 32'h41b18eae},
  {32'h452d4e6c, 32'h430470d7, 32'hc3b64456},
  {32'hc3b0084c, 32'hc2e69ace, 32'h43056978},
  {32'h44a5d967, 32'hc2aef724, 32'hc3cfe65f},
  {32'hc472659b, 32'hc2a5ef05, 32'hc289fa7d},
  {32'h45138d6c, 32'hc331bf39, 32'hc2573c06},
  {32'hc4ae4060, 32'h43189094, 32'hc2e66770},
  {32'h44031e56, 32'h42753e18, 32'hc39a2031},
  {32'hc4a76306, 32'h4361c803, 32'h438899bb},
  {32'h44a38fad, 32'h42c51325, 32'hc2ff3de0},
  {32'hc38f30cd, 32'hc2d292db, 32'hc32961a0},
  {32'h421f2f90, 32'h41720a81, 32'h4403e8fc},
  {32'hc4867ab1, 32'hc426ff6b, 32'h431098aa},
  {32'h44376b46, 32'h4344f636, 32'hc2ac72cd},
  {32'hc4c39c73, 32'h42c2c057, 32'hc1978a72},
  {32'h444828c2, 32'h4291966f, 32'hc2dd3c01},
  {32'hc4917e06, 32'hc3059e43, 32'h42ecb976},
  {32'h448221fe, 32'hc3c9e9ca, 32'hc2349dec},
  {32'hc4c31521, 32'hc0e67882, 32'h42b6e43b},
  {32'h44fca13f, 32'hc192ae1b, 32'hc3ffa4d6},
  {32'hc4a93290, 32'h4238b5a7, 32'hc346e6c6},
  {32'h445aae4c, 32'hc394d5db, 32'h436214c5},
  {32'hc3d388df, 32'h43922b33, 32'hc33701f2},
  {32'h4442576e, 32'hc280cc9f, 32'h437f1663},
  {32'hc4868ef5, 32'hc329b1d8, 32'h4389fdc6},
  {32'h449c0e94, 32'hc267aa4d, 32'h43d1f212},
  {32'hc509a298, 32'hc22566fe, 32'hc1aa3d10},
  {32'h4427090a, 32'hc3284909, 32'hc2b5fbd7},
  {32'hc4e0faae, 32'h4342103a, 32'hc385a68a},
  {32'h44f9bb6c, 32'h439484d0, 32'h3fe98d70},
  {32'hc4ed15db, 32'hc3868712, 32'h4307ad46},
  {32'h44b6d86e, 32'h43bceb73, 32'h42aa2ddc},
  {32'hc4ed9171, 32'h41e02183, 32'hc33046e5},
  {32'h4517b756, 32'hc28f0c5f, 32'h42bbf1c9},
  {32'hc450e42c, 32'h4320b194, 32'hc306a701},
  {32'h4506f844, 32'h421d1cd4, 32'hc32da900},
  {32'h43148e90, 32'h43173f96, 32'hc2ad78b8},
  {32'h43e91e5f, 32'hc26379fa, 32'h43864aad},
  {32'hc5201866, 32'hc355778c, 32'hc3165654},
  {32'hc2bd4918, 32'hc227fabc, 32'h43a1c4d2},
  {32'hc4f226f7, 32'hc2f1677d, 32'h4389ac6e},
  {32'h44882886, 32'hc30d79f9, 32'hc2bceb02},
  {32'hc41186dc, 32'hc3292141, 32'h427fc470},
  {32'h44cc3707, 32'h43290acd, 32'h43878389},
  {32'hc5005420, 32'h43226602, 32'hc31874df},
  {32'h44e44179, 32'hc2af5c7b, 32'hc2884bcd},
  {32'hc4fd1484, 32'hc31688cd, 32'hc1c24895},
  {32'h449ef649, 32'hc34db773, 32'hc3c9ef99},
  {32'hc4a17a72, 32'h43739536, 32'hc27c0ae8},
  {32'h43f8d488, 32'h43b823aa, 32'hc318645d},
  {32'hc4804dd8, 32'hc3ed1b1a, 32'hc194500c},
  {32'h44373b98, 32'h4388528b, 32'h4380b410},
  {32'hc510a40a, 32'hc2dff6af, 32'h42b681f2},
  {32'h44703300, 32'h428ce9a9, 32'h44065f55},
  {32'hc4a4c838, 32'h42aac428, 32'h41f859a5},
  {32'h44623b39, 32'hc342a42f, 32'h433eeb95},
  {32'hc2c79ce4, 32'h42f8dc0b, 32'hc3e746dd},
  {32'h44f623fe, 32'hc399c341, 32'h439b9cf1},
  {32'hc4302171, 32'hc31264c0, 32'hc39378cf},
  {32'h4496d3e5, 32'h43963567, 32'h4399670d},
  {32'hc4cd8945, 32'hc2988d35, 32'hc25da60a},
  {32'h444d24fc, 32'h430dd02c, 32'h4206d65e},
  {32'h432e21e7, 32'hc3a04d6c, 32'hc2d7cb04},
  {32'h44a01f62, 32'h4236abea, 32'h43b075fc},
  {32'hc383f970, 32'h4343a3c4, 32'h435f60a5},
  {32'h44754944, 32'hc33b0609, 32'hc3639c13},
  {32'hc3228e10, 32'hc39e74da, 32'h43285b62},
  {32'h44f1ea49, 32'h4338c4fd, 32'hc3833016},
  {32'hc426ffc0, 32'hc208124a, 32'h440af642},
  {32'h4401bb3d, 32'hc2b3e5d3, 32'h43e157f1},
  {32'hc3fc84ac, 32'hc3d005a6, 32'hc2d18571},
  {32'h4490464b, 32'h3fd71bb8, 32'hc353a88e},
  {32'hc4306388, 32'hc37e2ccd, 32'hc3109369},
  {32'h448a0f0c, 32'hc39a4cc0, 32'h42e74fea},
  {32'hc4b1ade6, 32'hc2ce8fdf, 32'h434fa63f},
  {32'h40c8bb00, 32'h4319e62c, 32'h430fdc36},
  {32'hc4906313, 32'h41df90eb, 32'h41fb49dc},
  {32'h438ed18e, 32'hc2b93d4e, 32'h41c04878},
  {32'hc38c19a8, 32'h421b3814, 32'h41a76e97},
  {32'h44aa78b7, 32'h43a65ee0, 32'h430bdca7},
  {32'hc4d943a8, 32'hc1e6b7b9, 32'hc3024028},
  {32'h440181b0, 32'h43286cac, 32'hc3379ced},
  {32'hc3f35218, 32'hc2801251, 32'hc2a01ac2},
  {32'h44f4d4f0, 32'h42e59089, 32'hc2835755},
  {32'hc388ac94, 32'hc0732f70, 32'h4288ef66},
  {32'h43b38f86, 32'h41aef720, 32'h42fcfcb2},
  {32'hc4cd6c5a, 32'hc30b258b, 32'hc2180a16},
  {32'hc4c709dc, 32'hc13cb9ae, 32'hbf025d3e},
  {32'h44f8c4f6, 32'h4341b245, 32'hc0675b48},
  {32'hc4e9c8bc, 32'hc344cc7c, 32'h4362ac90},
  {32'h44c4f8ea, 32'hc297e2dc, 32'h43c65710},
  {32'hc4d0deeb, 32'h427ecfc6, 32'hc3b51258},
  {32'h44176ce0, 32'h434945e2, 32'h43b1e18c},
  {32'hc4eb30b6, 32'h428a18eb, 32'hc3de0c0c},
  {32'h44d74479, 32'hc2dfd805, 32'hc3d453c9},
  {32'hc4dfaecd, 32'h4331caab, 32'hc29bee62},
  {32'h43cba0eb, 32'h42baf2d6, 32'hc252ef4e},
  {32'hc417a48e, 32'h427af9ab, 32'hc11c8b2a},
  {32'h4423d029, 32'hc202fac3, 32'h425fe715},
  {32'hc41601ec, 32'h428cc410, 32'hc3dd655c},
  {32'h43eb47e8, 32'hc3d43884, 32'hc3400a2a},
  {32'hc4287539, 32'h4380f66c, 32'hc2d0d334},
  {32'h441bb301, 32'h42b2a157, 32'h432e9b36},
  {32'hc2aab5c0, 32'h4397c073, 32'h42ea724a},
  {32'h45139da1, 32'hc2b7d92e, 32'h42d1ef73},
  {32'hc42c25d9, 32'h43180951, 32'hc2227d28},
  {32'h44a97bcb, 32'hc391d2da, 32'hc2ad06b9},
  {32'hc44e266e, 32'h43913b35, 32'h412571e6},
  {32'h441bc548, 32'hc21ae220, 32'h423e7afa},
  {32'hc435dc82, 32'hbfc80470, 32'hc31bc34d},
  {32'h44e56b9f, 32'h42a3705b, 32'h42926e25},
  {32'hc4d7dec0, 32'hc3cad3d5, 32'h4208d2e6},
  {32'h44041eea, 32'hc371c5fc, 32'h436d8501},
  {32'hc3c595bf, 32'hc31b94a4, 32'hc34e2090},
  {32'h44d32c33, 32'hc227d4f6, 32'h439f70a6},
  {32'hc4e27609, 32'hc1290cb8, 32'hc42fbe11},
  {32'h44de6a30, 32'hc38aa0f7, 32'h43543e62},
  {32'h430ef973, 32'h42a3a7f9, 32'h412fc66f},
  {32'h43ae2c0e, 32'hc3914f5b, 32'h43a2553e},
  {32'hc4d84c3c, 32'hc355652f, 32'hc39d6397},
  {32'h44c31260, 32'h43646e7f, 32'h4280db2a},
  {32'hc3709530, 32'hc31c40cb, 32'hc37216b9},
  {32'h44b51c11, 32'h42c3c117, 32'hc318e48e},
  {32'hc4af496b, 32'h4392ec95, 32'h4202afc2},
  {32'h422d2ff0, 32'h439529e8, 32'hc3bb3a54},
  {32'hc4afa5dc, 32'hc230ab6d, 32'h436c8404},
  {32'h444b3674, 32'h434e8b01, 32'h40cb95e4},
  {32'hc46639c0, 32'hc2b02ccc, 32'hc2c986f7},
  {32'h436e1fb0, 32'h42f1985b, 32'h435c1c8d},
  {32'hc48b1747, 32'hc2b9a41a, 32'hc3f21c46},
  {32'h4441b832, 32'hc3e75042, 32'h432127e2},
  {32'hc49a9c88, 32'hc30071a0, 32'hc42bb752},
  {32'h44689571, 32'hc30df512, 32'h436e6f85},
  {32'h42d3b8f8, 32'hc327d5f9, 32'h434dbd4e},
  {32'h44c75898, 32'h43b3395e, 32'h4289289a},
  {32'hc4de6b25, 32'hc267aea4, 32'hc3004b3e},
  {32'h448938f3, 32'h44082dc0, 32'h42ace0bf},
  {32'hc3d94130, 32'hc3218897, 32'h40b79a6a},
  {32'h437cbc38, 32'hc393dae0, 32'h4333b50f},
  {32'hc4dfc3ba, 32'h4307a5de, 32'hc25499f7},
  {32'h450ef94a, 32'hc2b06f3f, 32'hc2ac99c0},
  {32'hc488e977, 32'hc30601de, 32'hc3af1f7b},
  {32'h44c6a67a, 32'h4226256a, 32'h4345f540},
  {32'hc39afe4a, 32'hc3dfd51c, 32'h4411ac40},
  {32'h43810049, 32'hc41f6f80, 32'hc32323af},
  {32'hc4982d71, 32'hc40f46d0, 32'hc258115e},
  {32'h4519d118, 32'hc38ebaa2, 32'h41e48deb},
  {32'hc49719be, 32'hc3101d54, 32'h43b8252a},
  {32'h4441e878, 32'hc06e4eda, 32'h43cf10cc},
  {32'hc47c7366, 32'hc2a3afb3, 32'h420a1331},
  {32'h4446baf8, 32'h427e6344, 32'hc3a72b94},
  {32'hc48cdb12, 32'h430fd8a0, 32'hc25ecaa4},
  {32'h444014e8, 32'h418a7e56, 32'hc3d54345},
  {32'hc4babdc6, 32'h427b508e, 32'hc215225c},
  {32'h45052448, 32'hc3548987, 32'h43b72397},
  {32'hc3eb5980, 32'h4292ce29, 32'h42130c7b},
  {32'h440abc8e, 32'hc30c29e4, 32'hc31d02e2},
  {32'hc4ff6c96, 32'hc24d3012, 32'hc22628f9},
  {32'h448bd7c5, 32'hc42e8ce7, 32'h4393b964},
  {32'hc2c8e690, 32'h42d99dfd, 32'h43f3e8ad},
  {32'h45087d7e, 32'h432d21aa, 32'hc360eb71},
  {32'hc4232962, 32'h410f8c2f, 32'h433e0016},
  {32'hc2ff76bc, 32'hc2f22001, 32'hc24c571d},
  {32'hc5007e8e, 32'h43b50c7d, 32'hc3da5bdb},
  {32'h449bf85c, 32'h4229d61b, 32'hc3c295e3},
  {32'hc2f7f688, 32'hc28ece90, 32'hc33f9e75},
  {32'h44a4fb52, 32'h43341dc8, 32'h43c9b784},
  {32'hc5259541, 32'hc3c95884, 32'hc3aef558},
  {32'h4466a5cb, 32'h436335f1, 32'h4261ab67},
  {32'hc387ed7e, 32'h4205e220, 32'hc2cd063c},
  {32'h43195e70, 32'h41fe09b5, 32'hc371429b},
  {32'hc3dd548e, 32'h439a27e9, 32'h433de7db},
  {32'h449ae6e8, 32'hc391d7ad, 32'hc298555c},
  {32'hc4e580cc, 32'h41d5c820, 32'h42adf152},
  {32'h4488d572, 32'h42ac4bc0, 32'hc2fbed2d},
  {32'hc50767ae, 32'h432c9ddf, 32'h422e34b5},
  {32'hc276dc00, 32'h43295f41, 32'hc292f2f7},
  {32'hc41d5a50, 32'hc3756f81, 32'h4370409a},
  {32'h4476b431, 32'h42bf9e1e, 32'h4336fe4f},
  {32'hc4e7de59, 32'h4312885c, 32'h43238eef},
  {32'h441a2b80, 32'hc36f5c53, 32'h43099468},
  {32'hc4651ca8, 32'h42c57e76, 32'hc287a152},
  {32'h4494d8c1, 32'h432260a0, 32'h42dacba4},
  {32'hc49a2c0c, 32'hc3f89efa, 32'h42aed88b},
  {32'h4502f1fe, 32'h418fc533, 32'h42323298},
  {32'hc4f9bacd, 32'hc2dd74dd, 32'h41d4063f},
  {32'h44e53446, 32'hc0138290, 32'hc2733612},
  {32'h42946346, 32'h436e1ed0, 32'h418fc9c2},
  {32'h450fba8f, 32'h43baf63e, 32'hc2fb857f},
  {32'hc4bc3edc, 32'hc2ef63cb, 32'hc283ff03},
  {32'h44481796, 32'h42ec865d, 32'hc29dad5d},
  {32'hc49748a7, 32'hc29fd0c0, 32'h438fca1e},
  {32'h44f06b2a, 32'hc39b40f7, 32'hc3169cb5},
  {32'hc4e1ad70, 32'hc2b2f677, 32'h4295cd5e},
  {32'h450075b9, 32'hc269fb16, 32'hc324cea4},
  {32'hc4a3bd67, 32'hc3a8578a, 32'h43cc4ed5},
  {32'h44971d35, 32'hc18fbbfe, 32'h4383c8d1},
  {32'hc38c86a8, 32'h42209e56, 32'hc202d20e},
  {32'h4367847f, 32'h428ab4ea, 32'h4397ec33},
  {32'hc4b57546, 32'hc32f0e0e, 32'hc38fccbf},
  {32'h446bcc49, 32'h433dc8d9, 32'hc2ca662a},
  {32'hc43e52c9, 32'hc2621a5a, 32'h43e8056a},
  {32'h44bb4989, 32'h428dce3c, 32'hc3ab7852},
  {32'hc49116fd, 32'hc3935c94, 32'hc28abb41},
  {32'h4435a71a, 32'h4211a8ab, 32'hc36e26e2},
  {32'hc517d947, 32'h4372bcbf, 32'h439ef9eb},
  {32'h45094ad0, 32'hc327b5f8, 32'hc31c5261},
  {32'hc3848cbd, 32'h42f094e1, 32'hc14a4115},
  {32'hc2ebcc50, 32'hc2fe15ef, 32'hc330e72d},
  {32'hc3f7fcc4, 32'h43ac46ac, 32'hc3592c30},
  {32'h448cda4e, 32'hc3b9e637, 32'h43543bae},
  {32'hc4fa5d21, 32'hc0a866a8, 32'h434b5dc4},
  {32'h44b2d36f, 32'hc329f8c9, 32'h43162167},
  {32'hc511ef97, 32'hc3884f76, 32'hc292e314},
  {32'h44f955b0, 32'hc42767b9, 32'hc18a012c},
  {32'hc4e37c97, 32'hc348e8d0, 32'h40b906e2},
  {32'h428f3a68, 32'hc2b42a75, 32'h41aa4325},
  {32'hc46d9f1e, 32'hc33698e1, 32'hc30b7a55},
  {32'h450e1382, 32'h41b61b1c, 32'h438e4e0f},
  {32'hc48ab70a, 32'h430d21d4, 32'h428b64a0},
  {32'h43f6ae9f, 32'h433531e3, 32'h42f3c409},
  {32'hc4f02532, 32'h4370ec04, 32'hc352b12a},
  {32'h45071b4a, 32'hc3dc5e6f, 32'hc325abd4},
  {32'hc4c62788, 32'h43188244, 32'h42876318},
  {32'h442f53a5, 32'h42fadbe1, 32'h4380dfbf},
  {32'hc4bfb0fe, 32'hc367d4da, 32'hc31a04ae},
  {32'h44439731, 32'h4347e4eb, 32'hc27b7836},
  {32'hc49a78a1, 32'h42ccb23e, 32'h43284dc9},
  {32'h44441024, 32'hc361a62b, 32'hc38d64ad},
  {32'hc433ade6, 32'hc25f588a, 32'hc3302f6a},
  {32'h444211ea, 32'h42a94a22, 32'hc3b6b6f2},
  {32'hc4d38758, 32'hc2e13e2c, 32'h421f0ad3},
  {32'h43ce1f84, 32'h43820f92, 32'hc3539a33},
  {32'h40aaba40, 32'h4372555c, 32'hc414a465},
  {32'h43cb8606, 32'h43aad558, 32'h427d7e19},
  {32'hc4e2ba48, 32'hc1e562ee, 32'hc2e5f60a},
  {32'h44e15993, 32'hc3444406, 32'hc2689935},
  {32'hc4dda40c, 32'hc3f63a67, 32'hc273de65},
  {32'h4500ff99, 32'h43928fde, 32'h434f0151},
  {32'hc50080ab, 32'h4390e38c, 32'h43bce0af},
  {32'h451c25bf, 32'hc3bbc874, 32'h433ab535},
  {32'hc49d48c5, 32'hc2cc2d06, 32'hc26831b4},
  {32'h4499197c, 32'hc2d3d801, 32'h433f8449},
  {32'hc3a7b962, 32'hc3225b55, 32'h431787f6},
  {32'h43900bd3, 32'hc0f41f89, 32'hc22eb747},
  {32'hc1dffe00, 32'h433b00ec, 32'h437aa53b},
  {32'h44348e4b, 32'h4226dfe1, 32'h423aba0e},
  {32'hc4875dc0, 32'hc2df771a, 32'h4391d81e},
  {32'h432ff448, 32'h43a3cfef, 32'hc3014092},
  {32'hc5004894, 32'hc2a4b6c5, 32'h4356f61d},
  {32'h43f66ee4, 32'hc3a97a81, 32'h42310440},
  {32'hc4666792, 32'h4155944e, 32'hc31e5c4b},
  {32'h43c6c6d3, 32'h42f6096f, 32'hc3a5b372},
  {32'hc5230b20, 32'h42ae19b1, 32'hc381cd19},
  {32'h448ff3b5, 32'h428cd1bb, 32'hc277c96e},
  {32'hc404f323, 32'hc1f4b38f, 32'h42d57288},
  {32'h4512dc47, 32'hc0d83368, 32'h43b05757},
  {32'hc4b37a40, 32'hc2f8899f, 32'hc2707623},
  {32'h45041c39, 32'h438f6021, 32'h3fe8caf0},
  {32'hc41c828c, 32'h430d57db, 32'hc33032ee},
  {32'h44adc549, 32'hc3accdc2, 32'hc3926837},
  {32'hc4d6221c, 32'hc3128847, 32'h40977798},
  {32'h44e4db2b, 32'h42c6fa49, 32'h421e8726},
  {32'hc50ad18c, 32'h41fb250a, 32'hc40a66cc},
  {32'h43aabce4, 32'h426984c2, 32'h4347666d},
  {32'hc3b8a884, 32'h43c787b1, 32'h416c9571},
  {32'h448c6ffa, 32'h43b0ba9d, 32'h42b8e542},
  {32'hc5081323, 32'hbf6f32a0, 32'h42c34656},
  {32'h43d4fb98, 32'hc404b2ef, 32'hc2833e25},
  {32'h41e6e139, 32'hc31fe31c, 32'h41391eda},
  {32'h439ab17c, 32'hc21c9bdb, 32'hc3b056f1},
  {32'hc4d81b15, 32'h43495db1, 32'h4316f158},
  {32'h44bbd837, 32'hc221d8d9, 32'h430df8fb},
  {32'hc1da0020, 32'hc3827cde, 32'h42686815},
  {32'h44db58e0, 32'h435664a0, 32'hc38b9519},
  {32'hc45ac0bf, 32'h43da7918, 32'h42014465},
  {32'h44c82316, 32'hc2f928b9, 32'h43abf1d8},
  {32'hc3e68cf0, 32'h42320e42, 32'h439e23db},
  {32'h44efdba8, 32'hc2feec2e, 32'hc0998340},
  {32'hc497135b, 32'hc381ecc1, 32'h431095ce},
  {32'h42be7c80, 32'h43166287, 32'hc25d38a5},
  {32'hc4d5a27e, 32'h4326d27f, 32'hc2ab59fc},
  {32'h44de2b36, 32'h40adac10, 32'hc22c0008},
  {32'hc3f8dfe6, 32'hc2c23aba, 32'h42d7a29b},
  {32'h44059a12, 32'h434020b4, 32'h440cb860},
  {32'hc3becc30, 32'hc39c4ed3, 32'hc33cd09e},
  {32'h44b0c1ca, 32'h4314cc5a, 32'h42829fac},
  {32'hc51aacb0, 32'h42abe6f2, 32'h43b13d2a},
  {32'h45096ffd, 32'h424fef4a, 32'h4218b15e},
  {32'hc500638c, 32'h4162da66, 32'hc391f695},
  {32'h44cfb621, 32'hc39f3efa, 32'hc3410f05},
  {32'hc47b46b2, 32'h4342b4c3, 32'h42204501},
  {32'h44b114d6, 32'hc24acce6, 32'h42a2bf75},
  {32'hc4fdbda0, 32'h43c62023, 32'hc286d695},
  {32'h4491528b, 32'hc34c8337, 32'hc209593f},
  {32'hc40f46bd, 32'h42e22270, 32'hc3736c57},
  {32'h43d2b842, 32'hc2b9ce7b, 32'hc3052819},
  {32'hc385f420, 32'hc320d5dd, 32'h42e64bd0},
  {32'h44e2ca68, 32'hc2c0fae3, 32'hc2974032},
  {32'hc4be91d9, 32'h42423c90, 32'h42a82c82},
  {32'h4377a4f4, 32'hc2c19de0, 32'h4402d4b5},
  {32'hc397d9e4, 32'hc29304cd, 32'hc15423a8},
  {32'h4502092e, 32'h430a6ad0, 32'hc3289a2f},
  {32'hc4245c38, 32'hc2916f45, 32'hc2484edf},
  {32'h43a3fc40, 32'hc39cd661, 32'h4409b212},
  {32'hc4ddc2e5, 32'hc25da2a9, 32'hc32e66ed},
  {32'h44d24f2f, 32'h4322e702, 32'hc383e5fd},
  {32'hc4af0818, 32'hc2964918, 32'h4299ed18},
  {32'h449c63a1, 32'h41a1d0bb, 32'hc2d47c4c},
  {32'hc4ba0ee2, 32'hc2817eb1, 32'hc286df9c},
  {32'h44b2f3bb, 32'h43b2aca6, 32'h42160cc7},
  {32'hc40fb2e8, 32'h42a0fba3, 32'hc34e9766},
  {32'h447eaeed, 32'hc3ce5ba9, 32'hc3cffb65},
  {32'hc4c954f3, 32'h41dd3001, 32'h429cb0bb},
  {32'h444dafb0, 32'h43055650, 32'h42bc82f4},
  {32'hc33910dc, 32'hc3addd6b, 32'h41b3a378},
  {32'h4492071d, 32'hc309e96d, 32'hc2a5f45c},
  {32'hc4d82930, 32'hc32fef76, 32'h43450748},
  {32'h447b9b5b, 32'h4405ae1a, 32'hc2ae6fb4},
  {32'hc4bcb67f, 32'h42f75785, 32'hc3db461d},
  {32'h451a671f, 32'hc383caea, 32'h4322183e},
  {32'hc48924a5, 32'h42c73e5a, 32'hc34494e2},
  {32'h442c2523, 32'hc2ae9955, 32'h42c36702},
  {32'hc4cd2029, 32'hc318927f, 32'hc298848e},
  {32'h44fa97bb, 32'h43811300, 32'h436e23e7},
  {32'hc417f3d3, 32'h41f85d6d, 32'h42ab449e},
  {32'h44a5b575, 32'h4172edbc, 32'h425a438e},
  {32'hc388a23a, 32'h429c1ed3, 32'hc3bcd1a3},
  {32'h44b518ba, 32'hc2b3e65a, 32'hc1707264},
  {32'hc4d4aaf1, 32'h42abff97, 32'h428bc367},
  {32'h44b342fe, 32'h4384456c, 32'h42df86e3},
  {32'hc405e37a, 32'hc1290846, 32'h4379af81},
  {32'hc2e3a434, 32'h42cb9929, 32'h433305f6},
  {32'hc4ed56f0, 32'h4140d166, 32'hc2fa21fb},
  {32'h440d7133, 32'hc381a2d3, 32'hc3a20dcd},
  {32'hc31df404, 32'hc2e439fd, 32'hc3178091},
  {32'h4509f9c6, 32'h43052f5c, 32'hc348bbe6},
  {32'hc410dbb4, 32'hc325df91, 32'h436f605e},
  {32'h443a0d5c, 32'h42bfb7bb, 32'h42b14bc5},
  {32'hc3ed9010, 32'hc0d6819c, 32'hc1b163b4},
  {32'h44f35af7, 32'hc344d675, 32'h430a379c},
  {32'hc48fc770, 32'hc3ae0dee, 32'h421f06ca},
  {32'h450feac6, 32'hc321aa25, 32'hc3fc34de},
  {32'hc4ede847, 32'hc3bb3c18, 32'hc393fcf3},
  {32'h44a3ce28, 32'h43d7787f, 32'h4232f7c1},
  {32'hc463e054, 32'h438f1086, 32'hc0939a11},
  {32'h45160589, 32'h423706d4, 32'hc396b958},
  {32'hc4f01047, 32'h40e81476, 32'hc2838402},
  {32'h444cde92, 32'h423d0664, 32'hc3024935},
  {32'hc43ca50a, 32'h42011e5e, 32'h43b4d09f},
  {32'h449145c3, 32'h437bfb68, 32'h42856bf2},
  {32'hc50f7056, 32'h43e075f8, 32'hc3a9e661},
  {32'h4504e821, 32'h4400dda5, 32'h434b982b},
  {32'hc485bab8, 32'h4276c87c, 32'h40aa9388},
  {32'h4437a716, 32'h4238c47d, 32'h435d3dc9},
  {32'hc49304b0, 32'h430072ec, 32'h41b957f1},
  {32'h437776d4, 32'hc2b92586, 32'hc3962a9c},
  {32'hc382120f, 32'h410fc51b, 32'h424fd110},
  {32'h431e933e, 32'h439d6e03, 32'h42845e47},
  {32'hc4fbdd36, 32'h42663d08, 32'h436a3024},
  {32'h4481aa2b, 32'hc15363bd, 32'hc2026b85},
  {32'hc457ba0c, 32'hc3e0dfc1, 32'h42c6a064},
  {32'h433a96b0, 32'h42f46352, 32'h4229129c},
  {32'hc3e44bcc, 32'h42d63f3a, 32'hc39e3e36},
  {32'h442f7b1f, 32'hc3985c9e, 32'hc28339af},
  {32'hc2dec5d8, 32'hc3a65045, 32'hc3856186},
  {32'h44e6971b, 32'h432e096b, 32'h4348dd8f},
  {32'hc5102aa0, 32'h438a05e4, 32'hc2fa5a1c},
  {32'h44f10478, 32'h42d33c89, 32'hc2e6018f},
  {32'hc318d498, 32'h437b61f2, 32'hc316f3f3},
  {32'h44bc456e, 32'hc328c84b, 32'hc39cb59b},
  {32'hc43958f4, 32'hc26f5b8f, 32'h43964e79},
  {32'h44826423, 32'h42bcd119, 32'h43d560f5},
  {32'h41a27300, 32'h43779e28, 32'h43151eec},
  {32'h44e8fd70, 32'h42479b64, 32'h43b2d45e},
  {32'hc4e25da2, 32'hc3967e99, 32'h427cfc88},
  {32'h4421adc8, 32'hc3a044c4, 32'h4236f265},
  {32'hc48b48a0, 32'hc329f166, 32'hc330d281},
  {32'h44b27186, 32'hc35e9ab2, 32'hc3102672},
  {32'hc4493e51, 32'hc3526042, 32'h4345c633},
  {32'h43c32508, 32'h442b685c, 32'h43495273},
  {32'hc29f5930, 32'hc31a4680, 32'hc33275a9},
  {32'h43a99aad, 32'hc09cf673, 32'h4369d005},
  {32'hc4fbc0ac, 32'h433ec0fe, 32'hc2e0289c},
  {32'h44fcf91b, 32'hc3122504, 32'hc23964cf},
  {32'hc26ef0a0, 32'h43838721, 32'h437a325c},
  {32'h44a26582, 32'hc33b5711, 32'h432db582},
  {32'hc4ac65ae, 32'hc3817f9a, 32'hc22b0a84},
  {32'h44fe7216, 32'h442ef12b, 32'hc34a6317},
  {32'hc44fff53, 32'h41bbdc73, 32'h438e1ab3},
  {32'h4487f540, 32'hc20ceda2, 32'h43010172},
  {32'hc40ceb94, 32'h432a690f, 32'hc17ab2e2},
  {32'h44e9397f, 32'h416e5c31, 32'h42ba38d2},
  {32'hc260b5b0, 32'hc3a24012, 32'hc3808c98},
  {32'h45062066, 32'hc24e9df6, 32'h4324c8f0},
  {32'hc45e9398, 32'h432021ae, 32'hc38a81e3},
  {32'h438b9e40, 32'hc33a9a68, 32'hc14c65c6},
  {32'hc4a9fe22, 32'h422e5c8c, 32'h42dc90bb},
  {32'h4436e11f, 32'hc32df2d1, 32'hc2bb6ba0},
  {32'hc3b613a2, 32'h432e927b, 32'h41539d51},
  {32'h43909bac, 32'h424f41bb, 32'hc2944159},
  {32'h431c7fc8, 32'hc3678991, 32'hc30c1c78},
  {32'h44785154, 32'hc1d0ee81, 32'hc357680a},
  {32'hc4aa866a, 32'h41b8bdb5, 32'hc38ff92b},
  {32'h44869e3a, 32'hc273b038, 32'h435e6f96},
  {32'hc506c613, 32'hc28ba641, 32'h43be2bde},
  {32'h44d6d04a, 32'h438b45a7, 32'hc1b2b61b},
  {32'hc3922aa8, 32'hc000c744, 32'h42315fe3},
  {32'h45097c59, 32'h40e8a6b0, 32'hc253078c},
  {32'hc499df8c, 32'hc20c8afe, 32'hc375fac6},
  {32'h4506cd98, 32'h439fb05e, 32'h4421d2a4},
  {32'hc416ab7a, 32'h42b6a27f, 32'hc2e1dc84},
  {32'h441a8d24, 32'h43b39a47, 32'hc23fee32},
  {32'hc50033ac, 32'hc36fc172, 32'hc299f9ca},
  {32'h44f4bb6c, 32'hc29c6480, 32'h42d22742},
  {32'hc46ee002, 32'hc301dc39, 32'hc30423c3},
  {32'h4437a132, 32'h43a49dae, 32'h41e9446e},
  {32'hc41845e0, 32'h41a2ac40, 32'hc390c1a8},
  {32'hc2133538, 32'hc2a83053, 32'h43aede76},
  {32'hc50fa528, 32'h43aed268, 32'h42bb1902},
  {32'h450c7fa7, 32'hc1b1d2ef, 32'hc351b6ad},
  {32'hc51d506f, 32'h42f8fb07, 32'h442133d4},
  {32'h430c9498, 32'hc404f9cd, 32'hc2db5f79},
  {32'hc50b2b90, 32'h43aa85e4, 32'h429f6e88},
  {32'h451440b8, 32'h437299db, 32'hc2eb66d0},
  {32'hc3c7ba30, 32'h42a348b0, 32'hc28129a0},
  {32'h447eae34, 32'h435db497, 32'hc3a24c91},
  {32'hc463d4d0, 32'hc28409f5, 32'hc2cdef84},
  {32'h44c01835, 32'hc387b5bc, 32'hc30e4795},
  {32'hc33407c0, 32'h4324bb8e, 32'hc30773ff},
  {32'h43e49a04, 32'hc30af182, 32'h432c07a3},
  {32'hc50737b6, 32'hc31416aa, 32'hc2c204af},
  {32'h4486a72e, 32'hc3a63bfe, 32'hc2f95737},
  {32'hc4959f7c, 32'hc2b2b912, 32'h42bd9cac},
  {32'h4501a349, 32'h41f8a308, 32'hc386c9ba},
  {32'hc4d87431, 32'h430cc1df, 32'hc320e6f7},
  {32'h44882532, 32'h431b7f20, 32'h428ee6e2},
  {32'hc4b86c64, 32'hc257397a, 32'hc2d7061b},
  {32'h44359954, 32'hc315005c, 32'hc3251c54},
  {32'hc49a3c26, 32'hc39ef579, 32'hc385b69b},
  {32'h450f28a5, 32'h4318fd36, 32'h41de6dde},
  {32'hc45f114e, 32'h4312bcd8, 32'hc1128172},
  {32'hc30010c0, 32'h42ade00c, 32'hc2eb5f7e},
  {32'hc4422518, 32'h43538dfb, 32'h4376ee44},
  {32'h44d99997, 32'h429a6a1f, 32'hc2e20877},
  {32'hc31e6950, 32'h421e4c5c, 32'h431ee759},
  {32'h44a9075e, 32'hc2ccad6f, 32'hc3805f9d},
  {32'h436b0be4, 32'hc3da182d, 32'hc403b338},
  {32'h42ec3140, 32'h41dd8402, 32'h42806b61},
  {32'hc4a82b7f, 32'h4322a7d9, 32'hc2829fc0},
  {32'h449d7b73, 32'h436cc4eb, 32'h4323a05c},
  {32'hc51061c0, 32'hc345d7f8, 32'h43b9a70b},
  {32'h44bddbf6, 32'h42ac5220, 32'hc311ceea},
  {32'hc50b0d76, 32'hc2ccb939, 32'h4332b7fd},
  {32'h445a2242, 32'hc2138832, 32'hc2900e74},
  {32'hc4bc3ec7, 32'h43995be1, 32'h43e7b8f9},
  {32'h446dc576, 32'h4311c053, 32'hc2d16424},
  {32'hc46df2d0, 32'h4383ad98, 32'hc0bf892d},
  {32'h44c29c0f, 32'hc20cc02e, 32'h4308e4ce},
  {32'hc39ba34c, 32'h43a51403, 32'h43758416},
  {32'h4523ac20, 32'h41ef842a, 32'h43104777},
  {32'hc42c2276, 32'h43540f47, 32'hc3a1b3d4},
  {32'h44205234, 32'hc3642417, 32'hc3a77d81},
  {32'hc41456e0, 32'hc2c0bd1b, 32'h4405efc4},
  {32'h44f8fd4b, 32'hc234d592, 32'h43fd0489},
  {32'hc3cdc600, 32'hc19620ef, 32'h439b34b9},
  {32'h4416047c, 32'hc1ce3882, 32'h43eedc10},
  {32'hc453b6fc, 32'h4222abe2, 32'hc2f75a46},
  {32'h45243b09, 32'h4337abad, 32'hc33f281d},
  {32'hc445b5db, 32'hc3afabd7, 32'h420067d5},
  {32'h44ca78d1, 32'h4340879d, 32'hc326b80a},
  {32'hc3f21b05, 32'hc2a81a23, 32'hc31de354},
  {32'h444ed4c4, 32'hc2b27d4f, 32'hc1eae20f},
  {32'hc4c444dc, 32'h435437db, 32'hc3751480},
  {32'h440ee190, 32'hc3538fcb, 32'hc3d1fa81},
  {32'hc5148b6c, 32'hc28faf47, 32'h40e460fc},
  {32'h4499ac2e, 32'h43d6a09a, 32'h42a68c77},
  {32'h42fd88ff, 32'hc28f22bd, 32'hc2b74241},
  {32'h4427cecb, 32'h42c648eb, 32'h43920e25},
  {32'hc4d94deb, 32'hc297681d, 32'hc28490a5},
  {32'h4521ea41, 32'hc1f2e1c9, 32'h431f41a6},
  {32'h425c5040, 32'h42dece14, 32'hc38d68e9},
  {32'h448fb85d, 32'h42f4c45e, 32'hc3a78d7b},
  {32'hc451b756, 32'h430b2f9a, 32'h43191fa3},
  {32'h42ba2178, 32'hc1ed54a5, 32'h431100ec},
  {32'hc4ae0263, 32'hc3cc60f2, 32'h40bffea6},
  {32'h44398704, 32'h43877f32, 32'hc3679592},
  {32'hc4826b26, 32'h428075ad, 32'h43926166},
  {32'h4407fda6, 32'h42d6a944, 32'hc3b3a8de},
  {32'hc4deb002, 32'hc29b1f1a, 32'hc2c2f6c9},
  {32'h44b0a98b, 32'h43d675ec, 32'h43859619},
  {32'hc4f1dc01, 32'h435440d5, 32'h41dc0862},
  {32'h43bfdf49, 32'h43105a7a, 32'hc2b57037},
  {32'hc4e97809, 32'h439b5ef1, 32'hc3203c17},
  {32'h4477bc08, 32'hc102dc37, 32'hc39b79b4},
  {32'hc4fe4734, 32'h4321382d, 32'h43ad5197},
  {32'h447e5f64, 32'hc3926576, 32'h439f33a7},
  {32'hc4a4a258, 32'hc32aea14, 32'h43292367},
  {32'h4503d204, 32'h43cfba77, 32'h42b82057},
  {32'h4120b500, 32'h42a07b11, 32'h425bce3e},
  {32'h4418f6bc, 32'h42afb801, 32'hc39164c5},
  {32'hc39e9564, 32'h43a98583, 32'hc3148e0c},
  {32'h447fc302, 32'hc2f65f21, 32'hc2dd6228},
  {32'hc49784eb, 32'h439d8eb5, 32'hc315efc5},
  {32'h44b47eb4, 32'h433d00c7, 32'h43876467},
  {32'hc443314b, 32'h430e68bd, 32'hc33b7a83},
  {32'h44fea322, 32'hc3288bd1, 32'hc382437b},
  {32'hc4ab281d, 32'h42749f64, 32'h42f537e8},
  {32'h44a8cf62, 32'hc1c6f852, 32'hc3a51d08},
  {32'hc4f09151, 32'hc28e0343, 32'hc309e74b},
  {32'h441b295e, 32'h4202d689, 32'h4281d7eb},
  {32'hc433a854, 32'h42b44426, 32'h42d9b1d2},
  {32'h44a141b0, 32'h433a6f6f, 32'h42a66790},
  {32'hc48156b3, 32'h4236ce62, 32'h43520b59},
  {32'h4400af1e, 32'hc109f3da, 32'hc340487a},
  {32'hc3a7a750, 32'hc2ecc6b3, 32'hc31dba26},
  {32'h44405e32, 32'hc3261b8e, 32'hc30a0abf},
  {32'hc4fc7a52, 32'h42cebfae, 32'hc26c2fba},
  {32'h44f5c86a, 32'hc261e480, 32'h43b70a55},
  {32'h45002d50, 32'hc266b364, 32'hc1e32eb0},
  {32'hc3fbaf58, 32'h42770f16, 32'h4397bd1c},
  {32'h449d84a7, 32'hc331b2c2, 32'hc3b0fdbd},
  {32'hc4919991, 32'h431250a5, 32'hc2c7cc2b},
  {32'h44abf7b4, 32'hc37f8a9f, 32'hc3891d59},
  {32'hc3ac6700, 32'h431a2ec7, 32'h42878c89},
  {32'h44f6e323, 32'h4311cb05, 32'hc2657d1b},
  {32'hc49a4664, 32'h426f495a, 32'hc2563a4e},
  {32'h449f7e5c, 32'h43406ad3, 32'hc33ee807},
  {32'hc4c95e44, 32'hc30c2ab8, 32'hc351a729},
  {32'h451a779d, 32'hc00450da, 32'h441edaa1},
  {32'hc449f940, 32'h422976c6, 32'h436421e5},
  {32'h44949af8, 32'hbe039650, 32'h416541f4},
  {32'hc47b370d, 32'hc380fc87, 32'hc1bf4871},
  {32'h44a47141, 32'hc23dfbe7, 32'h438e8bca},
  {32'hc49272de, 32'hc3b4ade3, 32'h4094f06a},
  {32'h44d3774e, 32'hc25be7c0, 32'h432f904a},
  {32'hc4a4caf2, 32'hc33cd87c, 32'hc2bd6078},
  {32'h44acbaf4, 32'h42c4cede, 32'hc2cacaa2},
  {32'hc4e5279f, 32'hc28a1d13, 32'hc2cbedaa},
  {32'h44eef71d, 32'h421dbb2c, 32'hc21d2337},
  {32'hc4157c1d, 32'hc1bd3e28, 32'h42d2e2f2},
  {32'h43efa421, 32'h4374eb4c, 32'h4387ff68},
  {32'hc3477cf8, 32'hc23f7714, 32'h43b5b1ad},
  {32'h44fea3f4, 32'hc2f64704, 32'h41e4ee5d},
  {32'h425ed040, 32'h42ad28c7, 32'h43044f4e},
  {32'h431e075a, 32'hc2833b7c, 32'hc391b615},
  {32'hc3ff6dba, 32'h4351e341, 32'h42e0e60a},
  {32'h449c0831, 32'hc3283744, 32'hc396933f},
  {32'hc48eff20, 32'hc3793bd1, 32'hc2c4780e},
  {32'h4491d55a, 32'h415492ba, 32'hc35165c1},
  {32'hc484251d, 32'hc2afdcf1, 32'h414ebd40},
  {32'h44f73a3b, 32'h439061d7, 32'h4394240f},
  {32'hc4f6c9a4, 32'h42054ba0, 32'hc3151d8b},
  {32'h44d545be, 32'hc404ef64, 32'hc31fa8fa},
  {32'hc49ea817, 32'hc3c110d9, 32'hc2afe610},
  {32'h43779350, 32'hc3967b9b, 32'hc24c0eca},
  {32'hc46b88be, 32'h436ee35f, 32'h43b67a56},
  {32'h450768d8, 32'h42470113, 32'h440223b2},
  {32'hc4c4ca8a, 32'hc312c041, 32'hc2afe1e6},
  {32'h447c0c6a, 32'hc2b31dae, 32'hc122d504},
  {32'hc3bd748e, 32'h43abbc4c, 32'h437ce661},
  {32'h451330e0, 32'h42d8fe92, 32'h43be2f8d},
  {32'hc1693d40, 32'hc3760c93, 32'h439f938c},
  {32'h450d7cc4, 32'h4293f0ea, 32'h434f5992},
  {32'hc430dd6a, 32'hc42d48ec, 32'h43f3110a},
  {32'h44a2ecfc, 32'hc29e4b3a, 32'hc375dade},
  {32'hc4b60ff8, 32'h4401dc2c, 32'hc394e432},
  {32'h44d1c768, 32'h437cbe16, 32'h42e14c79},
  {32'hc3fa83f7, 32'h43041223, 32'h43c134ac},
  {32'h44588676, 32'h4317e7ee, 32'h428d4ae8},
  {32'hc408976a, 32'h43452e0e, 32'h42448010},
  {32'h4447d23a, 32'hc2ac302c, 32'hc30a37b6},
  {32'hc4890afe, 32'h42ef7929, 32'h4270c799},
  {32'h4505f9f9, 32'hc3eb9931, 32'hc16dd36f},
  {32'hc4ef0151, 32'h4394e4fc, 32'hc2a92e70},
  {32'h440f5a56, 32'hc37438b1, 32'h4340cfcb},
  {32'h41cc4d80, 32'hc2211266, 32'hc346eb4e},
  {32'h4515229b, 32'hc432d1e9, 32'h43047cda},
  {32'h4359bba4, 32'hc2185449, 32'hc2396592},
  {32'h447042e4, 32'hc3801ee6, 32'hc331ceb5},
  {32'hc4c12d1c, 32'h43aa45da, 32'hc386e07f},
  {32'h44f48076, 32'hc3e7c762, 32'h4317767a},
  {32'hc4fe0f85, 32'h4263c470, 32'h440b5140},
  {32'h44a20efe, 32'hc18a29d7, 32'hc2a51ee3},
  {32'hc4b294e8, 32'hc33fb2b9, 32'h4409fa5f},
  {32'h4492c898, 32'h435d45f8, 32'hc39fd809},
  {32'hc41d1573, 32'hc20c6505, 32'hc1bdc4cc},
  {32'h4472ee0b, 32'h4401a36a, 32'hc203ba02},
  {32'hc498034b, 32'hc2df112a, 32'hc146400f},
  {32'h44425c9c, 32'h4306ac55, 32'h431f2c0b},
  {32'hc4e3c0b0, 32'h4258eac6, 32'hc1dc6435},
  {32'h4513a1d4, 32'hc405b526, 32'h43c1f0b9},
  {32'hc4def779, 32'hc320f01c, 32'h43b08f7e},
  {32'h443bdb70, 32'hc39d4085, 32'hc363b064},
  {32'hc4bb2a56, 32'h42d2be06, 32'hc3d9325c},
  {32'h444b2234, 32'hc3999149, 32'hc3e18caa},
  {32'hc4a2191c, 32'hc2ad0c28, 32'h4346b641},
  {32'h44ad89cf, 32'hc200b3c2, 32'hc31a9a77},
  {32'hc4706bcf, 32'h400fea28, 32'hc2bbeb37},
  {32'h43ebafda, 32'hc2bcbd69, 32'h430f41a6},
  {32'hc4d46cb5, 32'h435486df, 32'h4320485c},
  {32'h4317ac84, 32'hc2845abf, 32'h4368c334},
  {32'hc49816ef, 32'hc325b601, 32'hc30c6481},
  {32'h44b72946, 32'h432c9a3a, 32'hc0da187e},
  {32'hc51270c3, 32'h42edc1f5, 32'hc2beff15},
  {32'h4492b41a, 32'h4329a025, 32'h425be342},
  {32'hc4cb6f1f, 32'hc33adacc, 32'hc2907ebc},
  {32'h44f5cddd, 32'hc1cb9426, 32'hc103de67},
  {32'hc45ac4c6, 32'h4388c2d3, 32'hc23209d3},
  {32'h448df121, 32'h42c902d5, 32'hc2930a51},
  {32'hc3d3f9ac, 32'hc37ee022, 32'h428e8638},
  {32'h44d152e0, 32'hc1c1815a, 32'hc35930c9},
  {32'hc4f93594, 32'hc274f5a2, 32'hc2b664f2},
  {32'h450771f3, 32'hc394f6a8, 32'h4301d1de},
  {32'hc4593391, 32'h4247c58d, 32'hc33a36d3},
  {32'h44076428, 32'h43c08327, 32'hc3cfbe09},
  {32'hc4e282d6, 32'h42d5a20b, 32'hc388190e},
  {32'h44e5fc7c, 32'h432c9374, 32'h437c177d},
  {32'hc51312cf, 32'hc38d6b5f, 32'h43f8cf14},
  {32'h450a21e6, 32'hc11c0d80, 32'hc2304517},
  {32'hc4834858, 32'hc28f46b2, 32'h4232fbd1},
  {32'h43e61b0a, 32'h42fc390b, 32'h43b071f6},
  {32'hc4ec91a2, 32'h4296421f, 32'h4357facf},
  {32'h4363bce9, 32'hc3c798e1, 32'hc2f65133},
  {32'hc40c7468, 32'hc2c8ae82, 32'h42fd7c0a},
  {32'h445db6fc, 32'hc3121b5f, 32'h438edd5f},
  {32'hc4f89f19, 32'hc37cd5ef, 32'hc31f326d},
  {32'h43e9194e, 32'hc380f261, 32'h42a57851},
  {32'hc4bb0f60, 32'h438876d6, 32'hc2209844},
  {32'h443c7b10, 32'hc35381bc, 32'h43845060},
  {32'hc4a73530, 32'h41b743c0, 32'h4385ee60},
  {32'h4501abe6, 32'hc2567ed2, 32'hc1e20d63},
  {32'hc48ddb99, 32'h43143ef3, 32'h4334d7fe},
  {32'h4385e444, 32'h42b7190a, 32'hc282fbf0},
  {32'hc2a7dbe0, 32'hc25fcac8, 32'hc3f56dcf},
  {32'h43fd27a0, 32'hc3229a4e, 32'h43a4ffc0},
  {32'hc4785f92, 32'hc4095947, 32'h4271cfc5},
  {32'h44b6340b, 32'h436e3ebc, 32'hc10aa7bd},
  {32'hc5062687, 32'hc30438ac, 32'h43c08dea},
  {32'h433b4c2e, 32'h43640cf4, 32'h4103cd66},
  {32'hc43d6aca, 32'h4406b852, 32'h438b02d2},
  {32'h44c58a96, 32'hc3c90dff, 32'h429319de},
  {32'hc4aabecc, 32'h42bf8de0, 32'h41f8b82e},
  {32'h451033ac, 32'hc168d417, 32'hc39a6773},
  {32'hc504c565, 32'hc3a5acf2, 32'h44031bad},
  {32'h44396caa, 32'h43c77653, 32'hc25960d9},
  {32'hc46a0682, 32'hc370bafe, 32'h422af7ae},
  {32'h449700c9, 32'hc3972120, 32'h430a8b42},
  {32'hc387fc41, 32'hc189e598, 32'h430576cf},
  {32'h44816e23, 32'h4391bf1e, 32'h439e50d3},
  {32'hc513db92, 32'hc369a36e, 32'hc3fa154b},
  {32'h448ef883, 32'h43abd542, 32'h429b0536},
  {32'hc49ecc79, 32'h4236b264, 32'hc27c34b1},
  {32'h443e19f4, 32'h430ac771, 32'hc35172d3},
  {32'hc496d4b9, 32'h43208994, 32'hc32410f8},
  {32'h443b2645, 32'h43907a3b, 32'hc2ae1a39},
  {32'hc5144204, 32'h432d1dcb, 32'h43ac2006},
  {32'h438f8f5e, 32'hc2fff840, 32'hc3be2cc7},
  {32'hc503789b, 32'hc34556e5, 32'h429e948e},
  {32'h438ab255, 32'hc29f7af7, 32'h42d0db37},
  {32'hc38dd43b, 32'hc3769ac9, 32'h43add97f},
  {32'h44a555f9, 32'hc4013032, 32'hc2e8adc2},
  {32'hc4f00e92, 32'hc3dc0fff, 32'h4380ca97},
  {32'h4408d5e4, 32'hc2a78f06, 32'h42a4f66c},
  {32'hc311c5d5, 32'h43065b5c, 32'h4396d836},
  {32'h44fe9c72, 32'h41cb002e, 32'hc3054933},
  {32'hc4801a5d, 32'h432bdcae, 32'h427290c4},
  {32'h442c6956, 32'hc082a5e9, 32'h4387457f},
  {32'hc4920fce, 32'h4361cf9d, 32'hc2dfd9db},
  {32'h44356f4a, 32'h432e808b, 32'hc2fdbab0},
  {32'hc330df78, 32'hc38b42c6, 32'hc37f8d7b},
  {32'h44c58dfa, 32'hc2031f1b, 32'h42144077},
  {32'hc4d54eaa, 32'h4391fa8f, 32'hc3648d65},
  {32'h4436f239, 32'hc21d19b8, 32'hc32e70c1},
  {32'hc3ee57cc, 32'hc223945a, 32'hc3aa0230},
  {32'h43d947e6, 32'hc123ae78, 32'h432bb44a},
  {32'hc4318b54, 32'hc389ad9d, 32'h42f621a0},
  {32'h43fde0d4, 32'h42f02ef1, 32'hc3f03a59},
  {32'hc499ba1b, 32'hc314e70e, 32'h42da7422},
  {32'h43d47ab4, 32'h425d92c4, 32'h43b83bfd},
  {32'hc47efed1, 32'hc30a9306, 32'h42ffa7d4},
  {32'h4506b345, 32'h42c4c826, 32'hc2027c0b},
  {32'hc41eaa0c, 32'hc365534a, 32'hc264c453},
  {32'h44f3af26, 32'h43224057, 32'hc3c231a5},
  {32'hc4c4b9b6, 32'hc40d22fd, 32'hc2c56b02},
  {32'h44dfb2ea, 32'h43a04e79, 32'hc37abd52},
  {32'hc3f9a027, 32'hc33f0952, 32'h437ad7e6},
  {32'h449af810, 32'h43868093, 32'h412ef164},
  {32'hc4e4bf92, 32'h4273224f, 32'h429033ab},
  {32'h44cc012c, 32'h4113f88c, 32'hc3fcb82a},
  {32'hc4ec3392, 32'hc319d3f4, 32'h43764f5c},
  {32'hc3731364, 32'hc3cad6df, 32'h42518f71},
  {32'hc4aa1f14, 32'hc3758a64, 32'h4383449d},
  {32'h44f76573, 32'h43d5734e, 32'h42c5bc0e},
  {32'hc4829947, 32'h42b3b057, 32'hc38288ae},
  {32'h450232cc, 32'h43a86c1a, 32'h43df5af2},
  {32'hc4e20c61, 32'hc3dceaae, 32'hc291e14d},
  {32'h451843be, 32'hc3697860, 32'hc328f1fe},
  {32'hc453d664, 32'h440698d6, 32'hc32f79dc},
  {32'h44ec8c5c, 32'hc3c390c8, 32'h4334868b},
  {32'hc355955c, 32'hc287de20, 32'h4367ae22},
  {32'h43f26cec, 32'hc30c1061, 32'h42333385},
  {32'hc3a010a5, 32'hc128a45b, 32'h424f04c9},
  {32'h44e0864c, 32'hc344c02f, 32'hc2dd749a},
  {32'h42f98cff, 32'h4225a042, 32'hc1b605dc},
  {32'h436805b5, 32'hc32c60bd, 32'hc32fede0},
  {32'hc40a6f8e, 32'hc301bc23, 32'hc37ec9b6},
  {32'h442eebd8, 32'h43a9fae9, 32'h437475b8},
  {32'hc3fd8a85, 32'hc2f8acaa, 32'h429bc26b},
  {32'h43a59f48, 32'hc3b0df60, 32'h42f9a5a6},
  {32'hc48fe0ca, 32'h439ae2ed, 32'h435ad2c4},
  {32'h441654bc, 32'hc3b26ea0, 32'hc397e1a6},
  {32'hc50354a8, 32'h3f182bc0, 32'h4345c27f},
  {32'h4492930a, 32'h43952d45, 32'h4357d994},
  {32'hc51001f8, 32'hc2527d68, 32'h42a57015},
  {32'hc3c30b28, 32'hc29224f6, 32'h43e63df7},
  {32'hc1f04260, 32'hc32ee967, 32'hc36b0450},
  {32'h43b848de, 32'h4330e4ef, 32'h423cfb4c},
  {32'hc43a3734, 32'hc3ae3b14, 32'h4206c84d},
  {32'h44f8b180, 32'h436cc2e8, 32'h41318a7c},
  {32'hc4c2be00, 32'hc2fa730f, 32'h438fb0fb},
  {32'h41cf9480, 32'h431c4bd6, 32'h42835cb8},
  {32'hc37d0970, 32'hc3d8f436, 32'hc32f0076},
  {32'h448470b2, 32'hc3e611d3, 32'h43350594},
  {32'hc46250e0, 32'h4391e5cd, 32'h431aa218},
  {32'h44ceb58d, 32'h43694fcf, 32'h431c311c},
  {32'hc4ae9dea, 32'hc36e0224, 32'hc4273380},
  {32'h43b7ecbb, 32'h431ebf7b, 32'h41896838},
  {32'hc4f32775, 32'h4084cda8, 32'hc3b8c3ed},
  {32'h444d5ba0, 32'hc0d473be, 32'h42898ed9},
  {32'hc50a8d73, 32'h42912e3c, 32'h43bfbaaa},
  {32'h4499082e, 32'h42c784ae, 32'hc4039142},
  {32'hc51225a6, 32'hc32a7f5e, 32'h41eb53e4},
  {32'h43430f68, 32'h42ff88ae, 32'h42f7221e},
  {32'hc4804715, 32'h42e176a8, 32'hc3829f26},
  {32'h44ab631f, 32'hc2c9cdb2, 32'h41a75c40},
  {32'hc3f3c3b4, 32'hc37cf688, 32'h438af28e},
  {32'h44045bf4, 32'h436aff25, 32'h43b9f0ca},
  {32'hc489f2e0, 32'h43b80c91, 32'h432af0c7},
  {32'h44440ffa, 32'h434af5d7, 32'hc33cfda3},
  {32'hc4ed4715, 32'h428d8123, 32'h40a88701},
  {32'h44ad6969, 32'h43a8fc04, 32'hc30d49aa},
  {32'hc389243c, 32'h428c43de, 32'hc27e904a},
  {32'h442295e5, 32'h41e0efdc, 32'h4331975e},
  {32'hc5076ead, 32'h4310128b, 32'hc31678c4},
  {32'h44460e4b, 32'h433e36e2, 32'hc2b0f284},
  {32'hc50139b2, 32'hc2f57de9, 32'hc2c9a4e3},
  {32'h45022dba, 32'hc2af720a, 32'h4245aae4},
  {32'hc48e65ae, 32'hc085b310, 32'h420ec014},
  {32'h44ea98d6, 32'h43619141, 32'h4387b215},
  {32'hc4cd0d3d, 32'h40b23296, 32'h42c4d6de},
  {32'h44708c92, 32'h4330832d, 32'h43b1435b},
  {32'hc4f7e78c, 32'h4355f984, 32'h428f1eea},
  {32'hc15d6e60, 32'h4338fdee, 32'hc2b08453},
  {32'hc413d946, 32'h42ee8ac9, 32'hc287ed0c},
  {32'h446ba6e9, 32'h43830a7d, 32'hc3d191b8},
  {32'hc40efbd7, 32'hc2ba5ce7, 32'h4364514d},
  {32'h44d876c6, 32'h426f6152, 32'h3fa05980},
  {32'hc4ed95aa, 32'h42c406aa, 32'h430be2f7},
  {32'h44ad2cca, 32'hc334bcb0, 32'hc35bef32},
  {32'hc497463f, 32'hc3731e93, 32'hc34f82f4},
  {32'h44309cc0, 32'hc30e9972, 32'hc04109b0},
  {32'hc4fddcfc, 32'h4359cdd1, 32'h4277c516},
  {32'h42cdaa66, 32'h43b1ff57, 32'hc3081c50},
  {32'hc502a935, 32'hc1f155a7, 32'h4311a6d9},
  {32'h44c76de8, 32'hc3bf26fe, 32'h40db7187},
  {32'hc4f8ce55, 32'h4389b3bf, 32'h44115542},
  {32'h447b0e7a, 32'h43a05b08, 32'hc33ee084},
  {32'hc44c127d, 32'h42eefa09, 32'h434a04fe},
  {32'h4515cac1, 32'h42aa7a8a, 32'h4302b84e},
  {32'hc4844d72, 32'h436880d8, 32'hc2196c35},
  {32'h438e9c98, 32'hc2d8710c, 32'h43854799},
  {32'hc39c6f33, 32'hc3d9a206, 32'hc2dd5aa9},
  {32'h438aa6ac, 32'hc2769a3a, 32'hc3b08957},
  {32'hc4a1c56d, 32'h43912ad8, 32'hc448ac54},
  {32'h44d10a03, 32'h4357eee0, 32'h42a44589},
  {32'hc36bbca0, 32'hc2f8d0dd, 32'h42b7eaa9},
  {32'h4434e408, 32'h437eca29, 32'hc1487820},
  {32'hc4f311c6, 32'hc22ad722, 32'h42a3cead},
  {32'h44bf510b, 32'h42a77d58, 32'hc3d4f165},
  {32'hc4bd6912, 32'h436f7b64, 32'hc2894f23},
  {32'h435a67a0, 32'hc2f75f22, 32'hc2a7f336},
  {32'hc3e49c9c, 32'hc392c3d7, 32'h4314bd8d},
  {32'h445f7d29, 32'h42e51644, 32'hc3d55ce9},
  {32'h4410e17e, 32'h4331cae2, 32'h408e9290},
  {32'h4413fd9b, 32'h440b0b74, 32'hc379a5fe},
  {32'hc4c5e73e, 32'h42c8b6f0, 32'hc39a4ac7},
  {32'h43cddf64, 32'h44025219, 32'h4308f5c8},
  {32'hc4e9af8c, 32'hc296278b, 32'h40b3a868},
  {32'h44faa62a, 32'h43ae203e, 32'h43769255},
  {32'hc4a099e2, 32'h433f09c4, 32'h43c2b7f5},
  {32'h4488baa7, 32'hc22ea684, 32'h43765f6a},
  {32'hc3ecb988, 32'h41b67aad, 32'hc21f23ce},
  {32'h44d37fce, 32'hc300c968, 32'hc2b9e499},
  {32'hc38c24e0, 32'hc2ffdab4, 32'h4305e648},
  {32'h44d0603c, 32'hc3093881, 32'h433ea0bf},
  {32'hc3d2b06a, 32'hc2bab8e4, 32'h43ab0daa},
  {32'h45102a2f, 32'h43738279, 32'h4322d3b2},
  {32'hc466d25e, 32'h4377b195, 32'hc3d72879},
  {32'h44d73761, 32'h435aa15f, 32'hc2ac9931},
  {32'hc41747d4, 32'h428c3889, 32'h42443977},
  {32'h44e3f7e3, 32'h434eb1f0, 32'hc32185f9},
  {32'hc3867674, 32'h429f6214, 32'h419c87b6},
  {32'h434e6a44, 32'hc32ea828, 32'hc2228df7},
  {32'hc380c49f, 32'hc2efe9eb, 32'hc350be61},
  {32'h44cd4a56, 32'hc214bbe9, 32'h4248859e},
  {32'hc5022af2, 32'hc2a00b6f, 32'h429553ac},
  {32'h44c82939, 32'hc410140e, 32'h416c5c2d},
  {32'hc505a0cb, 32'hc2b26b71, 32'hc3918dd2},
  {32'h441f84e5, 32'h40af8cfa, 32'hc34bebe7},
  {32'hc49cb3fa, 32'h41b0ed3a, 32'h42eb6f3f},
  {32'h44562a20, 32'hc3399591, 32'h42d0ceae},
  {32'hc3c8bb58, 32'hc29a254d, 32'hc4028567},
  {32'h44dbe529, 32'h435a3766, 32'hc2e2f5d2},
  {32'hc467db9c, 32'hc2c932cf, 32'h424b7199},
  {32'h4499b482, 32'h439f9c42, 32'h4396123e},
  {32'hc37beb0b, 32'h4380c4fb, 32'h435aab9e},
  {32'h449c2a1b, 32'h43d16092, 32'hc33382ee},
  {32'hc4ee2412, 32'h43bab387, 32'h4329ae43},
  {32'h44a1d53b, 32'h439cd44b, 32'hc3388e77},
  {32'hc4b1fb9c, 32'h43b51db6, 32'hc2a4db74},
  {32'h446d4248, 32'h42eab1f8, 32'h43123cda},
  {32'hc4987453, 32'h4310dc5a, 32'hc2a951ad},
  {32'h41fd5c00, 32'hc2bc5e13, 32'hc2f99bf0},
  {32'hc4edb7e2, 32'h436d8a51, 32'h43c12aa1},
  {32'h4431db48, 32'hc395bdb8, 32'hc37b839c},
  {32'hc4b5237b, 32'hc30e7ccb, 32'h4396a32e},
  {32'h449cfcdf, 32'h43e4e641, 32'h43daeca8},
  {32'hc4f85ca9, 32'h439b1ef2, 32'h441b10a4},
  {32'h4466bc63, 32'hc2d56bcf, 32'hc31196be},
  {32'hc4e8b27e, 32'hc2cd81fd, 32'h43274acf},
  {32'h442fc678, 32'hc1f2b196, 32'h43bb8c14},
  {32'hc458799f, 32'hc3ae14c3, 32'h432a0ff8},
  {32'h447480ac, 32'h426302f2, 32'hc3db7fb9},
  {32'hc4f76bb8, 32'hc393b8a1, 32'h43cf6b22},
  {32'h442984cc, 32'h403d6100, 32'hc3b665ba},
  {32'hc484a5d0, 32'hc3125cd6, 32'h4301b86a},
  {32'h4519418e, 32'h42f10d3a, 32'hc35d3432},
  {32'hc4ea8fc1, 32'h4285bc3f, 32'hc3d72a5f},
  {32'h444013ca, 32'hc3383221, 32'h42d6f5ac},
  {32'hc502a867, 32'h43ce0ae9, 32'hc3cf841c},
  {32'h44a55a94, 32'hc2904e2a, 32'h431064a0},
  {32'hc512abe6, 32'hc38cd2a8, 32'h4366f115},
  {32'h43bf15d8, 32'hc22f5fc6, 32'h420f4e3d},
  {32'hc4bb85e9, 32'h41834f18, 32'h412bc160},
  {32'h44267b9c, 32'hc2a016dc, 32'hc2877620},
  {32'hc499d334, 32'h438f534c, 32'h43bcf174},
  {32'h44275bde, 32'hc397cf99, 32'h430b5ad4},
  {32'hc4cbde36, 32'h43e30678, 32'hc34e727f},
  {32'h450c54c8, 32'hc383913b, 32'hc3c5f1e8},
  {32'hc4a46f24, 32'h4374a495, 32'hc2cf40e4},
  {32'h44ed6344, 32'hc3cb9635, 32'hc39331b4},
  {32'hc405cb4c, 32'h43539b59, 32'hc3a350b2},
  {32'h4510f53d, 32'h423fe269, 32'h43d2c7b9},
  {32'hc3b009c3, 32'h43429ee9, 32'hc31a895a},
  {32'h440ceb89, 32'hbf22de29, 32'hc39c734a},
  {32'hc3dcd97c, 32'hc32f43f0, 32'hc11d88b8},
  {32'h44b7354d, 32'hc33cfa73, 32'h4164f934},
  {32'hc50ddc20, 32'hc35cbc14, 32'hc35fb8fb},
  {32'h42813690, 32'h420ee2cf, 32'hc34a0651},
  {32'hc462d868, 32'h41d994c1, 32'h4271d2de},
  {32'h45035a32, 32'h432eca3b, 32'hc316724f},
  {32'hc44204f2, 32'hc18ad1c3, 32'hc0809778},
  {32'h4506cb06, 32'h43c012b4, 32'hc15a679a},
  {32'hc4a61ca4, 32'h4343b4af, 32'h432bb9f2},
  {32'h450053c5, 32'h431218b8, 32'h43735c20},
  {32'h4251557b, 32'hc3d11901, 32'hc3287aae},
  {32'h4501a0a6, 32'h42d6438a, 32'hc381f16d},
  {32'hc4f2ede6, 32'h42ce0f2d, 32'h43506175},
  {32'h45192ea6, 32'h431c7279, 32'hc33d38f6},
  {32'hc464d137, 32'hc359f5ff, 32'hc30844fc},
  {32'h45168e0c, 32'h43bcd42d, 32'h4284f2bf},
  {32'hc4ca1b4b, 32'hc2b6bdc4, 32'hc335da6b},
  {32'h44d26148, 32'h4318cc31, 32'hc2c38b59},
  {32'hc5013201, 32'h43399264, 32'hc307ced9},
  {32'h449d6226, 32'h432a570e, 32'hc30f3a45},
  {32'hc2a88960, 32'hc3940f5d, 32'h42b78b04},
  {32'h445fd82e, 32'h4377ad2d, 32'hc35683b9},
  {32'hc4e14ade, 32'hc4366ccc, 32'hc35f773b},
  {32'h44c23824, 32'h42a4bf61, 32'hc00e84e4},
  {32'hc3863f99, 32'h426984df, 32'hc3d895ce},
  {32'h43947ec2, 32'h434b3f13, 32'hc31e0028},
  {32'hc436e572, 32'h4370447c, 32'hc3103f1b},
  {32'h44e6e072, 32'hc292f5e6, 32'hc38e071f},
  {32'hc383b1ac, 32'h435178a3, 32'hc2b3f0b6},
  {32'h44573768, 32'hc30ac830, 32'h44109134},
  {32'hc517a7a5, 32'h424461dd, 32'hc2af514a},
  {32'h450a545f, 32'hc303751c, 32'h431c1d74},
  {32'hc4de3a3b, 32'hc20a67d2, 32'h4218202c},
  {32'h446f2d9b, 32'h431f80ba, 32'h42c75b01},
  {32'hc41aad9b, 32'hc3e7b90f, 32'hc26ff782},
  {32'h43fd97a8, 32'hc3072984, 32'h431c0e27},
  {32'hc4d10140, 32'h43c9999b, 32'hc251aeea},
  {32'h45093790, 32'hc28d3cc0, 32'h440aaae1},
  {32'hc4f9faff, 32'hc31eb45a, 32'hc326271c},
  {32'h43c04e8d, 32'hc3a73a8c, 32'h42ed5c08},
  {32'hc45e27c4, 32'hc1f68a63, 32'hc2b7bf17},
  {32'h44870200, 32'hc3034734, 32'h434482dd},
  {32'hc4b20f64, 32'h42de7c41, 32'h4381e8be},
  {32'h43634ea0, 32'h43adc175, 32'hc3752b07},
  {32'hc5087b65, 32'h431a38aa, 32'h42d91b56},
  {32'h4502bb08, 32'hc39af010, 32'h434c3328},
  {32'hc46f9e9f, 32'hc327967e, 32'hc3a4a75f},
  {32'h44e109dd, 32'hc36232e4, 32'h41c828c5},
  {32'h41e880c0, 32'hc08cf1ec, 32'hc391b237},
  {32'h450e2158, 32'hc376628a, 32'h4238bec2},
  {32'hc31e81d0, 32'hc309eecb, 32'hc31f1d41},
  {32'h4314294a, 32'hc191ea7b, 32'hc399e60b},
  {32'hc4736402, 32'hc3234f23, 32'hc36ff847},
  {32'h44361650, 32'hc299956c, 32'h42899ed2},
  {32'hc518eddd, 32'hc2d3a145, 32'h4397b136},
  {32'h4514078e, 32'h439c32e8, 32'hc2aee0a6},
  {32'hc3bb54e0, 32'hc3324aa7, 32'h41a8c292},
  {32'h452a8321, 32'hc2e6e520, 32'h424eb49e},
  {32'hc50b65fe, 32'h41710004, 32'h43344c24},
  {32'h43c31062, 32'hc3807675, 32'h430992e5},
  {32'hc4f308b8, 32'hc3040eb9, 32'h41d7315a},
  {32'h448c0c82, 32'hc3cd81ef, 32'h431e7e66},
  {32'hc4399b6f, 32'h43515fd3, 32'h425d0137},
  {32'h4498e6e7, 32'hc364c89e, 32'h42b32ea6},
  {32'hc419825e, 32'h428c7604, 32'hc31391c8},
  {32'h449344d7, 32'hc3553c16, 32'h42f6590f},
  {32'hc50ad7a7, 32'hc2cb9345, 32'hc3069e0a},
  {32'h444ca5f4, 32'h4299181e, 32'hc0d43d08},
  {32'hc4bcbed6, 32'h42268926, 32'hc31241a6},
  {32'h44df3e69, 32'h438e10ee, 32'hc38b1757},
  {32'hc2788d98, 32'h43730baf, 32'h40102976},
  {32'h444c8ac0, 32'h425e1918, 32'hc291908b},
  {32'hc3c2a4f8, 32'h421500e7, 32'hc2d7fd9a},
  {32'h44d45fba, 32'h42923074, 32'h43ec279c},
  {32'hc5084be3, 32'hc1926374, 32'hc37fbe5a},
  {32'h449bdaa9, 32'h4356e720, 32'h43dc62f4},
  {32'hc3a0ff88, 32'h437b42b5, 32'h434b8fcc},
  {32'h449c1f5b, 32'h43448afe, 32'h4398ed1a},
  {32'hc4f2f64c, 32'h42d4e13b, 32'hc3228354},
  {32'h45048786, 32'hc2f72d08, 32'hc31c29d2},
  {32'hc4776582, 32'hc35618f3, 32'hc35988ec},
  {32'h4433ee6c, 32'h42640c47, 32'hc3d34b51},
  {32'hc50b09e9, 32'hc2d183ca, 32'h43539ccd},
  {32'h443f0b20, 32'h4256295e, 32'h42f0f540},
  {32'hc4876eca, 32'h440171b3, 32'hc327e91d},
  {32'h449623fb, 32'h41488f99, 32'hc2830e22},
  {32'hc510e6a7, 32'hc1b8aa84, 32'hc31fb175},
  {32'hc2bbcda8, 32'hc2b21dcb, 32'h41da76a0},
  {32'hc33d2400, 32'hc3024413, 32'hc33fb7f3},
  {32'h43f45684, 32'hc3b65e39, 32'h41c8acb5},
  {32'hc3774400, 32'h4287525c, 32'h43881f4f},
  {32'h4453ea22, 32'h4385b6fc, 32'h42a7f738},
  {32'hc514e4c6, 32'h43492677, 32'h43624255},
  {32'h4504220a, 32'h436aa1b2, 32'hc28e013a},
  {32'hc4ee816e, 32'hc2e4caf7, 32'h436a562f},
  {32'hc3a50968, 32'hc3102b14, 32'hc384578b},
  {32'h44d63dc3, 32'h434fe026, 32'h43b71362},
  {32'hc507a761, 32'h438a029b, 32'hc28d81a4},
  {32'h42d41350, 32'h41abc607, 32'h4264d1a4},
  {32'hc4fff648, 32'h414ebfa8, 32'hbfa34cb4},
  {32'h451e6f3c, 32'hc31b7125, 32'hc3935b1f},
  {32'hc512b6b3, 32'hc3d35447, 32'h4354f7bd},
  {32'h45114af6, 32'hc3913bb6, 32'hc38d552a},
  {32'hc4fa7d6c, 32'h428e9e9f, 32'hc1e9d2c4},
  {32'h44a968b5, 32'hc24c5d23, 32'h42bfb590},
  {32'hc4813317, 32'h438c58e7, 32'h42b02c11},
  {32'h450fa8b1, 32'h434ef081, 32'h432372b5},
  {32'hc3f229c0, 32'h430d66ca, 32'hc2ab582b},
  {32'h435f4dec, 32'hc2e758b5, 32'hc39b3ac0},
  {32'hc432d684, 32'hc2ae3913, 32'h43c33b24},
  {32'h450139d0, 32'hc302e8d0, 32'h427d5fde},
  {32'hc4248e3e, 32'hc3869ca0, 32'h43335fa7},
  {32'h44cc418f, 32'h42ae9ce2, 32'h43279094},
  {32'hc3d6b43b, 32'hc2883bbc, 32'hc38651f7},
  {32'h44d84003, 32'h42ae608f, 32'h439e6a31},
  {32'hc3feec45, 32'hc2a32be9, 32'hc2efdd5f},
  {32'h45086380, 32'hc31d5a7b, 32'h43bfcf89},
  {32'hc41d5d2f, 32'h41f2e1d1, 32'hc3fe6214},
  {32'h4503d28e, 32'h435ef71e, 32'h42a60266},
  {32'hc4b57c8c, 32'hc35ddb04, 32'hc30d7143},
  {32'h448907a0, 32'h439bacf5, 32'hc32016aa},
  {32'h4293351c, 32'hc2e0bae7, 32'h42afc657},
  {32'h44bafe8b, 32'hc41a6d73, 32'h437a9ada},
  {32'hc4873100, 32'h4298ca66, 32'hc342f354},
  {32'h44ae080b, 32'h43c7a439, 32'h4341a71e},
  {32'hc4616438, 32'h43300890, 32'hc24e058b},
  {32'h4306afc8, 32'hc0fb7762, 32'h442d9572},
  {32'hc4030924, 32'h4238bf91, 32'h3fca23da},
  {32'h45004163, 32'h439e7242, 32'h439d5541},
  {32'hc46bef89, 32'h4328947e, 32'hc40f9d58},
  {32'h43b42105, 32'h43030ecc, 32'h4212dcfa},
  {32'hc42cc648, 32'hc2d2654c, 32'hc38a47d9},
  {32'h436e4800, 32'h43f3a737, 32'h43878b7b},
  {32'hc50ff4ca, 32'hc194edd3, 32'hc1868b1a},
  {32'h449ea0f5, 32'h4317762a, 32'h42abb9c3},
  {32'hc3d01914, 32'hc33b5982, 32'hc220c034},
  {32'h4521b5dd, 32'h42e719d2, 32'h43a21229},
  {32'hc38c2898, 32'h4286cecd, 32'hc3489daa},
  {32'h4458917e, 32'hc3d70345, 32'hc3f85d88},
  {32'hc49b7b77, 32'hc3d149f8, 32'h435f317f},
  {32'h44eb3c2c, 32'h42d08987, 32'h432750c6},
  {32'hc43cead2, 32'h43a283be, 32'h4295c534},
  {32'h44f3c457, 32'h42c8ae55, 32'hc3762a70},
  {32'hc4e3ac0e, 32'hc202582c, 32'hc1f9f50c},
  {32'h445dcc64, 32'hc26f38f0, 32'hc2d54f7e},
  {32'hc4a4bbcc, 32'hc2f1d13c, 32'hc2177a97},
  {32'h4482ae00, 32'hc1fbaa2f, 32'hc2d9c0e5},
  {32'hc4540bd8, 32'hc2986af4, 32'hc27b881d},
  {32'h4501485b, 32'h41dd4719, 32'hc21e102c},
  {32'hc4c390b9, 32'h4362fc84, 32'hc232835c},
  {32'h44748d64, 32'hc21ce0c3, 32'hc3311166},
  {32'hc4ffd299, 32'h4336612e, 32'hc33fd421},
  {32'h44e7e6af, 32'h43950a68, 32'hc300e597},
  {32'hc4f682f6, 32'hc354c6a7, 32'hc3cc0a4f},
  {32'h44c05739, 32'hc3274a2c, 32'h439b1a44},
  {32'hc50d468e, 32'hc20003b0, 32'h4370ec36},
  {32'h4470f7b6, 32'hc36cbf2f, 32'h422d8f56},
  {32'hc4d5d776, 32'h404bf6d2, 32'hc3e24780},
  {32'h438ee9ae, 32'hc3a98586, 32'h4354b03e},
  {32'hc45ed37e, 32'h43019cae, 32'h437e0f85},
  {32'h44b7a32f, 32'h43ac21e1, 32'h4338c071},
  {32'hc495c9e4, 32'h426f68ac, 32'h423921b4},
  {32'h4507ec11, 32'h431c5dda, 32'hc3e04721},
  {32'hc425def7, 32'h43a8c54a, 32'h42b022db},
  {32'h4325c088, 32'hc3079914, 32'hc3633ca5},
  {32'hc4789f36, 32'hc24fe5fa, 32'h4398a3c8},
  {32'h44df6a01, 32'h4362b300, 32'h43ba278d},
  {32'hc437c389, 32'hc380a7fd, 32'h4402536f},
  {32'h44db5ff5, 32'hc3a12fef, 32'hc291deb4},
  {32'hc4fe9dcf, 32'h42d6ffb6, 32'h42e32a04},
  {32'h449c0270, 32'h43157ba2, 32'h42a8fda1},
  {32'hc49c47a2, 32'h43994d3a, 32'h408a443c},
  {32'h44fa408c, 32'h429442bc, 32'h42e0b324},
  {32'hc450126c, 32'h4304e670, 32'h42425ca4},
  {32'h45083e8c, 32'hc396f333, 32'h424a94f8},
  {32'hc3d6c844, 32'hc349601c, 32'h42479c9d},
  {32'h4512a460, 32'h42c09276, 32'hc356bc3e},
  {32'h44090043, 32'h43584af3, 32'hc39a18e9},
  {32'h42ffe380, 32'h4302e0e0, 32'hc3be2b37},
  {32'hc503eb23, 32'h439c18d3, 32'hc2622484},
  {32'h4471377d, 32'hc05da844, 32'hc2ebf346},
  {32'hc4f0773e, 32'hc2a77107, 32'h43a6ef9d},
  {32'h44bcb6d9, 32'h4239f7cf, 32'h436ae1fa},
  {32'hc491e5d6, 32'hc2e1c271, 32'hc32a7a7c},
  {32'h44ee4366, 32'hc38d8dcc, 32'h43a84381},
  {32'h42786e20, 32'h41435bd0, 32'hc1c759f7},
  {32'hc273269c, 32'h43102706, 32'h43211307},
  {32'hc4f7a9f4, 32'h4325d1c4, 32'hc3160022},
  {32'h44f5bee8, 32'h4342f8f7, 32'h438ffe36},
  {32'hc4851a70, 32'hc3dda0d4, 32'h43e1f5fa},
  {32'h441f6263, 32'h438189c9, 32'hc38a60fa},
  {32'hc45e3ab2, 32'hc3065aec, 32'h43a199ec},
  {32'h45177de1, 32'hc383c3bb, 32'h42a48373},
  {32'hc5062c28, 32'h439383e6, 32'h420b41d0},
  {32'h436a46c0, 32'h42d8e1a3, 32'h41f62186},
  {32'hc4b4618b, 32'h42ae4eb0, 32'hc343854d},
  {32'h447ce648, 32'hc3817d09, 32'h43445846},
  {32'hc434a114, 32'h43a23533, 32'h433468d1},
  {32'h43ec5f4c, 32'h4383470c, 32'hc30da039},
  {32'hc4c34718, 32'h437d0dc2, 32'h43397ee6},
  {32'h43cf7470, 32'h43016ebe, 32'hc2878e00},
  {32'hc2da5450, 32'h4359858e, 32'hc301bc69},
  {32'h447b8a1a, 32'hc3fd4ba8, 32'h432b75a9},
  {32'hc3fc295a, 32'h43346f69, 32'hc1e2a3c5},
  {32'h44ed0671, 32'h43c41de7, 32'hc21166c5},
  {32'hc457a42c, 32'hc37465d2, 32'h42cb4fe3},
  {32'h44ab6e02, 32'h43dd3b6f, 32'hc35ea5cd},
  {32'hc4cf444b, 32'hc3873244, 32'hc3843579},
  {32'h448c20cf, 32'hc2047101, 32'hc3853cca},
  {32'hc48524ee, 32'hc38678d7, 32'hc3590e22},
  {32'h432d433e, 32'h43a3fc42, 32'hc31d6d95},
  {32'hc38adcfe, 32'hc4022a6b, 32'h439aec1b},
  {32'h4483218d, 32'hc3af3930, 32'hc0f67cfc},
  {32'hc4b5bfdf, 32'hc28a3a40, 32'h42037a64},
  {32'h4497c5a3, 32'h42302c26, 32'h4267751a},
  {32'hc4bcb9bd, 32'h43344c42, 32'h431faf82},
  {32'h44c45b62, 32'hc2f294f6, 32'hc2f87f66},
  {32'hc3d25fb4, 32'h40d7d6a6, 32'hc23f5504},
  {32'h411a0ff0, 32'hc39f5f1c, 32'h42815ff5},
  {32'hc4b636ba, 32'hc2df92b9, 32'h43b19dc5},
  {32'h445869cc, 32'h435e8c61, 32'hc37ee146},
  {32'hc22292b0, 32'h422ae4a9, 32'h4295072c},
  {32'h4426be86, 32'hc39bcdfc, 32'h43039d02},
  {32'hc337f272, 32'hc34740e6, 32'hc2d2c025},
  {32'h4502e4bd, 32'hc2c1c752, 32'hc3d9e757},
  {32'hc4c1bd14, 32'hc32435b8, 32'h43fd68ee},
  {32'h441ca01a, 32'h429c42eb, 32'h4318704d},
  {32'hc4bcd71c, 32'hc2f4b82c, 32'h439fffd3},
  {32'h44442ab5, 32'hc22c4602, 32'hc29a7dd4},
  {32'hc44b64ed, 32'hc297cc7d, 32'hc37e0adb},
  {32'h445702c2, 32'h42e0b85d, 32'hc14e4acf},
  {32'hc4abfaba, 32'h42be3ef3, 32'hc23a7667},
  {32'h443bddd5, 32'h42c73e9f, 32'hc1c8d439},
  {32'hc4ea7330, 32'h40ab9656, 32'h43b67b3f},
  {32'hc3620e34, 32'h434b92da, 32'hc316503a},
  {32'h42f83af1, 32'h42b24666, 32'h439cdf45},
  {32'h442c4a53, 32'hc318cfc9, 32'h4310a588},
  {32'h4162ef00, 32'h4368bf17, 32'h41f11300},
  {32'h44cfe045, 32'hc298ae1c, 32'h438e41eb},
  {32'hc47ca13c, 32'h43a1369d, 32'hc2d3e447},
  {32'h44d38b8c, 32'hc3993edd, 32'hc3a45dcd},
  {32'hc45f1dd6, 32'h432527b0, 32'hc380ffa3},
  {32'h451d769b, 32'h4356e610, 32'h4345935b},
  {32'hc39c5b0a, 32'hc405b6d3, 32'h43f8f14f},
  {32'h450ae270, 32'h4347a75b, 32'h419b3bc1},
  {32'hc4471662, 32'hc303e614, 32'h43b8de0a},
  {32'h4511dfde, 32'h40dc1648, 32'hc2bb2b00},
  {32'hc4459869, 32'hc3d832ad, 32'h4242ad28},
  {32'h44df528f, 32'hc343ebd3, 32'h434982b2},
  {32'hc4cb6429, 32'h4337e4fc, 32'h420ae4be},
  {32'h44d01e1e, 32'hc35ed5a3, 32'hc310c64e},
  {32'hc375621d, 32'hc30e97cd, 32'h41a15165},
  {32'h445e4cbc, 32'hc2333551, 32'h42b54f51},
  {32'hc3ddd266, 32'h410999bf, 32'hc3a5b1a9},
  {32'h42a49f00, 32'h436c9962, 32'h43521e3f},
  {32'hc4958ec0, 32'hc259df65, 32'h430b49a3},
  {32'hc3385a20, 32'h43c64dfc, 32'hc4159856},
  {32'hc495be85, 32'h433a415a, 32'hc345162b},
  {32'h44c4ae9b, 32'hc1004276, 32'h4316f9f8},
  {32'hc4d3f94a, 32'hc31a9bab, 32'hc36ec882},
  {32'h44169919, 32'h4341cc42, 32'hc2efc5b1},
  {32'hc3dc2d80, 32'hc2a74013, 32'hc35ce44d},
  {32'h44c2db07, 32'h4339059d, 32'h4367a850},
  {32'hc5113c33, 32'h42b4228f, 32'hc3a990fd},
  {32'h44d7906b, 32'hc3935207, 32'h4391905b},
  {32'hc4aba7e6, 32'hc3e36b6e, 32'h42f8b738},
  {32'h451a19d8, 32'hc30193cc, 32'h431ad11f},
  {32'hc4695264, 32'hc3b2f5f8, 32'hc32c9e43},
  {32'h44d2383c, 32'h4211910a, 32'hc25d2c2d},
  {32'hc48f7e4c, 32'h4320d86f, 32'hc120f456},
  {32'h3da1c800, 32'hc380e8cf, 32'h4212aa9a},
  {32'hc4859eb4, 32'hc1cd1a0a, 32'hc2c2915a},
  {32'h44bb80cd, 32'hc243342c, 32'hc383dbe9},
  {32'hc508cccf, 32'h424f8ba3, 32'hc3629672},
  {32'h4415654e, 32'h41a9ff86, 32'h41e42d30},
  {32'h4383e700, 32'h42e25264, 32'hc33eff27},
  {32'h44e78501, 32'h43a788d5, 32'h43a98a2f},
  {32'h431ce9af, 32'hc21f9fa9, 32'hc2e3fa9a},
  {32'h44e41647, 32'h42369f2e, 32'hc3ef025a},
  {32'hc5126608, 32'hc1917e95, 32'hc3010e21},
  {32'h44a01cac, 32'hc35349c0, 32'hc1a1dded},
  {32'hc3c35633, 32'hc194693d, 32'hc24600b6},
  {32'h439663b0, 32'hc3087553, 32'h4172c3ae},
  {32'hc4d9aa1c, 32'hc28be2c2, 32'h41dbee99},
  {32'h450bfb9e, 32'hc4096370, 32'hc355b8b1},
  {32'hc3725360, 32'hc1b0465e, 32'h42fbe68e},
  {32'h449cf4e4, 32'h41fa43d8, 32'h43bd66b9},
  {32'hc5016db6, 32'hc351fd44, 32'hc30db8d2},
  {32'h445ee565, 32'hc3436581, 32'h422cfc3b},
  {32'hc4b2b4e2, 32'h421d1257, 32'h402e5386},
  {32'h448c4b3f, 32'hc1e0b635, 32'h424b10f8},
  {32'hc3e7fadc, 32'h439377d1, 32'hc2fe6bbf},
  {32'h429ebba5, 32'hc235cebd, 32'h4384588e},
  {32'hc4f5e7a8, 32'h42990f15, 32'h42ab3ada},
  {32'h4407a364, 32'h434b5a33, 32'h42cbecb4},
  {32'hc48fd0e2, 32'hc3aacfae, 32'h43a89126},
  {32'h43f7a318, 32'hc38b608b, 32'hc3840fce},
  {32'hc48b0d9a, 32'h428a98a1, 32'hc3e6c38e},
  {32'h446ee15a, 32'h43ffdaeb, 32'h42a98776},
  {32'hc5096cb4, 32'h43c175d6, 32'h4352970f},
  {32'h44a8d8d2, 32'h4360b5fb, 32'h4204ca6d},
  {32'hc4c68eea, 32'hc34a9256, 32'h43806a96},
  {32'h44dc00fd, 32'h43e6ab18, 32'hc32c8d84},
  {32'hc4ed8af7, 32'h4316b852, 32'hc3543070},
  {32'h43d076b0, 32'h40407c34, 32'h41f2a8dc},
  {32'hc4b29361, 32'hc241ab0a, 32'hc265f849},
  {32'h44ef3836, 32'hc339d7b3, 32'hc41be3ec},
  {32'hc4a83b7b, 32'hc09571de, 32'h41984a94},
  {32'h44c12c00, 32'hc39952ea, 32'h439d7564},
  {32'hc3be6252, 32'h433c16e2, 32'hc290aeb9},
  {32'h451b6e5f, 32'h431bb441, 32'hc1f42642},
  {32'hc33ee9ec, 32'h42b83d37, 32'hc365794a},
  {32'h45094644, 32'h4308b9a2, 32'h43fd0172},
  {32'hc4f7e274, 32'h42eff4a7, 32'h428d95e5},
  {32'h44da7b0b, 32'hc20c2005, 32'h42f748f8},
  {32'hc50bc3e0, 32'hc3a62745, 32'hc31233c0},
  {32'h44d68993, 32'hc269229a, 32'hc33c1e5b},
  {32'hc4a6cdcb, 32'h439d4877, 32'hc32a04b9},
  {32'h4442becb, 32'h41aa30e0, 32'h41771741},
  {32'h425e82e7, 32'h415cb7d8, 32'hc381f061},
  {32'h44edb536, 32'hc35b3e31, 32'hc3927f95},
  {32'hc4b5571c, 32'hc39e1eb7, 32'hc327fe0f},
  {32'h44a6e230, 32'hc31e4d9b, 32'h4376a7ef},
  {32'hc416bd68, 32'h43667b4b, 32'hc3a38c75},
  {32'h44c01c82, 32'h43aaf9ff, 32'h43125233},
  {32'hc3fb733c, 32'h425ac172, 32'h43b0f55f},
  {32'h44bff0da, 32'h42f2c080, 32'h43148c60},
  {32'hc500b68a, 32'h42da4c99, 32'hc3b97db4},
  {32'h44f267a7, 32'h42974a9f, 32'h43cca314},
  {32'hc43b2052, 32'h43222a66, 32'hc2ce0bc1},
  {32'h441778d6, 32'h430375cf, 32'hc27ea09a},
  {32'hc494bea4, 32'hc2cf672c, 32'h43003ac9},
  {32'h45136fc9, 32'hc34d27e6, 32'h43abbe7a},
  {32'hc44cb84c, 32'hc36a42e9, 32'h43e0b7cc},
  {32'h45069ed3, 32'h429bb626, 32'hc12ba78d},
  {32'h43919586, 32'h420d81a0, 32'hc32ba194},
  {32'h44105e00, 32'h42f4d125, 32'hc3de7e66},
  {32'hc4206103, 32'h42b3b45a, 32'hc350829a},
  {32'h4287a7e0, 32'hc2d86100, 32'hc2faad73},
  {32'hc4feb06b, 32'h43bd9b1b, 32'hc306b90b},
  {32'h44bd6308, 32'hc343d2b2, 32'h42fd7034},
  {32'hc3d37e80, 32'h439a0186, 32'hc398b6be},
  {32'h44a82d28, 32'hc3b06582, 32'h4216ff69},
  {32'hc497d8eb, 32'h42ad519b, 32'hc36ba777},
  {32'h4484036f, 32'h4272b9a1, 32'hc2c61860},
  {32'hc50c1980, 32'h44007bf2, 32'h42bfc492},
  {32'h44113276, 32'hc37c5cc6, 32'h433bcbf6},
  {32'hc4e400a4, 32'hc3b513c1, 32'hc3457b8d},
  {32'h44e8ba88, 32'h43494458, 32'hc2c2f922},
  {32'hc50a37a1, 32'h415c1d84, 32'hc3346245},
  {32'h44d9dbb5, 32'h42b02bb4, 32'h436549e4},
  {32'hc4f66bef, 32'hc02196ef, 32'hc3271366},
  {32'h44158978, 32'h429b1f28, 32'h43d2f02a},
  {32'hc36dac00, 32'hc2bb7a66, 32'hc3f1e3be},
  {32'h43300c18, 32'hc2f6123a, 32'h42d8f291},
  {32'h42fbe83b, 32'h43c1c42e, 32'hc22284ee},
  {32'h450ded38, 32'hc41ee16a, 32'hc38dc48b},
  {32'hc40cb3ba, 32'h42421663, 32'hc290929a},
  {32'h450d7668, 32'h42ad2fe8, 32'h4303bdbf},
  {32'hc41daeae, 32'hc40dab89, 32'h43b8ec0b},
  {32'h444c3dd0, 32'h42e21ee2, 32'hc2b02d91},
  {32'hc4adca6f, 32'h43fed05b, 32'h43041f86},
  {32'h44c9b874, 32'h43726ea2, 32'h42a600f9},
  {32'hc45450f5, 32'hc2d0a168, 32'hc330528a},
  {32'h43b44912, 32'hc2fbb3be, 32'hc11d3b96},
  {32'hc4e5765b, 32'h436846dc, 32'h433abc9f},
  {32'h44cc5fc1, 32'hc34716dd, 32'hc38a1c4b},
  {32'hc2ec6240, 32'hc32e9b5b, 32'hc253ebd4},
  {32'h440c7534, 32'h422da2db, 32'h41a503a2},
  {32'hc51358b4, 32'h43658898, 32'h4279da8b},
  {32'h44bba9aa, 32'hc3b908c0, 32'hc3be76c9},
  {32'hc4d778cc, 32'h412f52e6, 32'h42e5651b},
  {32'h4429fa3b, 32'h431a2393, 32'h42794548},
  {32'hc45de386, 32'hc3387f90, 32'h4390170e},
  {32'h44be73ce, 32'h42040024, 32'h4398dc28},
  {32'hc4b23065, 32'hc35cf6cc, 32'hc345becf},
  {32'h44fa6a23, 32'h4395748e, 32'hc33e4acc},
  {32'hc5043162, 32'hc1b3e88a, 32'hc38e1e6c},
  {32'h45013a3e, 32'h41ff594c, 32'h426eaa65},
  {32'hc39543b6, 32'h42e69287, 32'h438e8f04},
  {32'h443f58fc, 32'hc3d7030b, 32'h43910690},
  {32'hc50a31e9, 32'hc267a001, 32'h42c2daf8},
  {32'h45122a74, 32'hc3a19581, 32'hc26fc485},
  {32'hc4dfbb94, 32'hc3604e75, 32'h423ab408},
  {32'h43276782, 32'h43aaf6d1, 32'h438d5141},
  {32'hc487cf59, 32'hc313197e, 32'h434c6e51},
  {32'h44dae31b, 32'h43642c4c, 32'hc183fda4},
  {32'hc465aec2, 32'hc2ac6c63, 32'h438ad32d},
  {32'h439145a8, 32'hc389742e, 32'hc2e5adfa},
  {32'hc4299b64, 32'h432f61f0, 32'hc3f1f712},
  {32'h4468ddba, 32'hc3ae84c9, 32'h43393a90},
  {32'hc4759f22, 32'hc28d40c5, 32'hc27a6c5a},
  {32'h44de3ea4, 32'hc29e2cfc, 32'hc2daa933},
  {32'hc4a222c6, 32'h42cb2505, 32'hc1f17192},
  {32'h451bea50, 32'hc2b5c6f5, 32'h431afd9d},
  {32'hc505f8de, 32'h43595abb, 32'hc2c1fb98},
  {32'h44c1a27b, 32'hc39a37c7, 32'hc3751362},
  {32'hc50972ea, 32'h42d5d654, 32'h419e5972},
  {32'h4410a060, 32'h43882c54, 32'hc413e0fb},
  {32'hc416159c, 32'hc224a650, 32'hc352131a},
  {32'h4464ff4b, 32'hc3eb4a27, 32'hc33ec975},
  {32'hc3d52532, 32'h40c4d268, 32'hc3fbd451},
  {32'h43d540dc, 32'hc3d90ee4, 32'h42a550b5},
  {32'hc506d14e, 32'hc326fb3c, 32'hc331fba9},
  {32'h450fed64, 32'h43d42d73, 32'h434e44ab},
  {32'hc4f50417, 32'hc3848103, 32'h402e40e0},
  {32'h44af78a9, 32'hc3491e0d, 32'h432ecd85},
  {32'hc3fc7c8d, 32'hc3340055, 32'h4315cbf6},
  {32'h43bc99f8, 32'hc31cd02b, 32'h434a1edb},
  {32'hc3a2d7e6, 32'h42ab4d7c, 32'hc2b67c96},
  {32'h449427a3, 32'hc3522333, 32'hc382e8fe},
  {32'hc45743b0, 32'h4332b53d, 32'hc3ca2f14},
  {32'h447855d2, 32'hc39fd437, 32'hc3b83ade},
  {32'hc4e16a52, 32'h43b497b0, 32'hbff8fa42},
  {32'h44a72364, 32'hc31e2424, 32'hc1abbdca},
  {32'hc481c2e0, 32'hc3a6ced4, 32'h431703f6},
  {32'h45018bfe, 32'hc329a036, 32'h43d08b76},
  {32'hc4e1b5ee, 32'hc24aa898, 32'h41a412ea},
  {32'h44019494, 32'hc2e65808, 32'h43f2a7a5},
  {32'hc4dcfaf4, 32'h41db82e0, 32'h42d70ffc},
  {32'h4508e82f, 32'h42f77f6b, 32'hc1ae9e0c},
  {32'hc4279e8a, 32'h434d5b0e, 32'h435a8063},
  {32'h440aa93d, 32'h42d94b3a, 32'h438add06},
  {32'hc49ad0ad, 32'hc2d9c43c, 32'h43b8690a},
  {32'h43452b1c, 32'hc2e1d309, 32'hc2b02b2f},
  {32'hc3ae3132, 32'hc3124c71, 32'hc304b7be},
  {32'h4503905a, 32'h43a47671, 32'hc3827d7c},
  {32'hc500f1d7, 32'h43ad346b, 32'hc34f4e39},
  {32'h451077b4, 32'h430d1f06, 32'hc3634e53},
  {32'hc4da4de7, 32'hc29272fc, 32'h41c95be6},
  {32'h44f6a9cf, 32'hc34fec43, 32'hc3262e08},
  {32'hc20e8480, 32'h439e403d, 32'hc34ac3ec},
  {32'h433134b0, 32'hc32fab7e, 32'hbffb1931},
  {32'hc43475b2, 32'h438ae740, 32'hc39c6b82},
  {32'h4519ac70, 32'h43bb64fe, 32'h41dd6cab},
  {32'hc4babeb8, 32'hc2591657, 32'hc359fb11},
  {32'h43125350, 32'h4393582b, 32'hc43d3006},
  {32'hc43fb4c1, 32'h4356dd56, 32'h42ce5536},
  {32'h44c30cf7, 32'hc2c0121a, 32'h432aea78},
  {32'hc45e2dc8, 32'h43b66502, 32'h42c8ba1a},
  {32'hc1c7ecc0, 32'hc1227ec7, 32'hc31a1de2},
  {32'hc508dde7, 32'hc3e18806, 32'hc2cb9607},
  {32'h42a79210, 32'hc442cb07, 32'hc30e306a},
  {32'hc428279a, 32'hc3751488, 32'hc390c9a0},
  {32'h44a9da0c, 32'hc1ac8b54, 32'hc1ffcd43},
  {32'hc479d6bd, 32'hc2806c50, 32'h43f9bdd9},
  {32'h4519ef03, 32'hc32042b6, 32'hc2963182},
  {32'hc4f5ece1, 32'h430f2e17, 32'h43458d9c},
  {32'h44bc8b3c, 32'hc36959bc, 32'hc28db029},
  {32'hc49fdf66, 32'h43bd90d2, 32'hc2dfafbe},
  {32'h44a741c3, 32'hc3506a96, 32'h42fab436},
  {32'hc3b7ba7d, 32'h44065b59, 32'hc387f504},
  {32'h448770a6, 32'hc29f56fd, 32'h42176cbb},
  {32'hc463c090, 32'h431d7a2a, 32'h431822a2},
  {32'h44d5d45c, 32'hc378b7da, 32'h42352f3e},
  {32'hc5073e7f, 32'h43bedd78, 32'hc2bc206f},
  {32'h452080f8, 32'hc393c997, 32'h42e0ed50},
  {32'hc4fe0e51, 32'h433c16ae, 32'h43dffe48},
  {32'h443cba96, 32'hc3560442, 32'hc313a277},
  {32'hc46eb0e0, 32'hc383f7d1, 32'h430a23a8},
  {32'h45123447, 32'hc353af1c, 32'h42953ef3},
  {32'hc4a9a722, 32'hc31d4339, 32'h42c831bc},
  {32'h44d05d18, 32'h42893a92, 32'hc287bc36},
  {32'hc39ecc60, 32'hc36dd9ad, 32'h435fb347},
  {32'h44123fec, 32'h431d12ab, 32'hc38c14d9},
  {32'h431165c7, 32'hc399e10d, 32'hc2dded9c},
  {32'h4458cfc5, 32'hc39b8138, 32'h4415da80},
  {32'hc4dd0ca4, 32'hc3aaa20b, 32'hc3484f54},
  {32'h44d8f6be, 32'hc3668a1b, 32'h435a6ac2},
  {32'hc459e9c2, 32'h43221a53, 32'hc3b8d023},
  {32'h4448ab04, 32'hc310204e, 32'hc3b66980},
  {32'hc4a131b6, 32'h43f56db9, 32'hc33bbe42},
  {32'h44180efe, 32'h43e05cc8, 32'hc34fea95},
  {32'hc47d972c, 32'h43743db0, 32'hc30ad950},
  {32'h445159c8, 32'h42fc854d, 32'hc227462e},
  {32'hc4913baf, 32'h43d53b3a, 32'hc2a94f19},
  {32'h443bfab8, 32'hc2025bdc, 32'h425981f8},
  {32'hc4379b74, 32'h430e1e71, 32'hc3a80e33},
  {32'h43803d55, 32'hc3ed37a3, 32'hc16a1fff},
  {32'hc4e96b07, 32'hc12b60f4, 32'h4344c34d},
  {32'h44f90166, 32'h43269ab1, 32'hc1ceaf97},
  {32'hc44fcc38, 32'hc314981e, 32'h42459798},
  {32'h451d1aa6, 32'hc383f15d, 32'hc3839920},
  {32'hc47445ac, 32'h42b74a4a, 32'hc327e4e8},
  {32'h4481d9f6, 32'h42e2b1f5, 32'hc3377ad4},
  {32'hc4337cd3, 32'hc322e20e, 32'hc27411d3},
  {32'h44b245ed, 32'h422ff79f, 32'h41b86f1b},
  {32'hc46ae56a, 32'h431137af, 32'h42998c40},
  {32'h4428bc36, 32'h42849b8e, 32'h42f7cccc},
  {32'hc4d98a0d, 32'hc36ee6fd, 32'h435c1f80},
  {32'h45074a78, 32'hc223da75, 32'hc3165f4e},
  {32'hc4aa297c, 32'hc1926ca8, 32'hc167d7a0},
  {32'h43de8cc2, 32'hc392635c, 32'h42c98a96},
  {32'hc5115904, 32'h436bff67, 32'h41e02dea},
  {32'h432c1a60, 32'hc3109bba, 32'hc18a257a},
  {32'hc4cc3cfa, 32'h435dbe09, 32'hc2af74df},
  {32'h44cf07a3, 32'h431499f3, 32'hc30bce62},
  {32'hc4c79251, 32'h433c33b3, 32'hc2f778ee},
  {32'h444e70ec, 32'h43ecd28e, 32'h42b36848},
  {32'hc44a83e2, 32'h428ff520, 32'hc2142d38},
  {32'h4477dfec, 32'hc35c44a7, 32'h437351e7},
  {32'hc3fc7c98, 32'h43584e81, 32'hc1ae47d4},
  {32'h44589e68, 32'hc3609a98, 32'hc28a4568},
  {32'hc5097862, 32'hc251e068, 32'h436c8f86},
  {32'h449b2ec4, 32'h425ececc, 32'hc2576d0c},
  {32'hc4fbd32f, 32'hc3a1a843, 32'hc2aefc14},
  {32'h447691ab, 32'h414ecd93, 32'h436a4b6e},
  {32'hc446eb1e, 32'h43ba529f, 32'h43469a91},
  {32'h448e7fa2, 32'hc363fda0, 32'hc34f0406},
  {32'hc421b390, 32'hc27f5116, 32'h440abb86},
  {32'h44f0ccb1, 32'hc38bdbc4, 32'hc1146be5},
  {32'hc3db4510, 32'hc34622cc, 32'h43ee0745},
  {32'h438d1b08, 32'hc2d624a7, 32'hc36a206e},
  {32'hc4776f5e, 32'h42c90bb3, 32'h43417322},
  {32'h44932808, 32'hc2e8616d, 32'hc2ee297c},
  {32'hc4f6fde1, 32'hc2e1443d, 32'h4395add6},
  {32'h4500f93f, 32'h41e8f0b5, 32'hc327a809},
  {32'hc4edfcda, 32'h42474941, 32'h4399c712},
  {32'hc3b36e6f, 32'h43e61b13, 32'h428fbcaa},
  {32'hc4e2f8ab, 32'hc2f2df9b, 32'h42e6aedf},
  {32'h44e5b127, 32'hc29333be, 32'h42881232},
  {32'hc4c2a7a4, 32'hc2815404, 32'hc3a09e24},
  {32'h44e9803a, 32'hc3abbbf0, 32'hc348a125},
  {32'hc49619d4, 32'hc28fc8f2, 32'hc18c32fb},
  {32'h45182a04, 32'h429b2965, 32'h4207bcd7},
  {32'hc3f6b1b1, 32'h4380e6aa, 32'h42d0a827},
  {32'h4496156c, 32'hc1c62505, 32'hc37b27c4},
  {32'hc31c9418, 32'h42a41ee2, 32'hc2e0b689},
  {32'hc4a9bdf4, 32'hc3b233e9, 32'h426fb1e7},
  {32'h44d3a110, 32'hc173f153, 32'hc32f9c47},
  {32'hc4d585b0, 32'h428c86f0, 32'h429c7f5c},
  {32'h44fa9929, 32'hc1c5006a, 32'h4318e630},
  {32'hc4894fd5, 32'h4377d07d, 32'hc32cae43},
  {32'h44a793b0, 32'hc33445bf, 32'h429f2a1e},
  {32'hc3b7d457, 32'h43d326c4, 32'hc1bb3486},
  {32'h44f9949c, 32'hc3af18dd, 32'hc2815106},
  {32'hc41e2f44, 32'hc37ce50a, 32'h43b09e20},
  {32'h44735110, 32'h430c6a1a, 32'hc3ae6360},
  {32'hc50de881, 32'hc380fc21, 32'h439a5b22},
  {32'h4479b164, 32'h439466c5, 32'hc3205aa7},
  {32'hc4de1d70, 32'hc2d01bc3, 32'hc31237df},
  {32'h44dec450, 32'hc37baa07, 32'hc3cd542f},
  {32'hc4908cf6, 32'hc366eb74, 32'h438c027d},
  {32'h44d8690d, 32'hc351ed93, 32'hc2db3565},
  {32'hc3639cb0, 32'hc27e2b28, 32'h43e403fd},
  {32'h43595e98, 32'h42bda6e2, 32'h430415b8},
  {32'hc4a55870, 32'h42523206, 32'hc3e283f0},
  {32'h44c8fb5e, 32'hc2dd9614, 32'h4301f81e},
  {32'hc4c16910, 32'h42def7af, 32'hc1e65fd6},
  {32'h43155da0, 32'hc1ef94b5, 32'hc39e5ac7},
  {32'hc3605da0, 32'hc35abea1, 32'h437f8b51},
  {32'h43e255d4, 32'h43114180, 32'hc3334d61},
  {32'hc46e78b4, 32'hc2a292a7, 32'h43e2c0c9},
  {32'h4525fa52, 32'hc3fa5159, 32'hc39b2f94},
  {32'hc362a52d, 32'hc1c526ac, 32'h420291fa},
  {32'h44886bde, 32'hc284b313, 32'hc35a2e25},
  {32'hc48a482c, 32'h4270580a, 32'h43391b43},
  {32'h44ff7590, 32'hc2ae2396, 32'h42a7996e},
  {32'hc468a5ae, 32'hc39efa6c, 32'h43058e7f},
  {32'h44c8463c, 32'hc33c1df4, 32'hc3947c6d},
  {32'hc3857618, 32'hc3314a9c, 32'h4089b6d0},
  {32'h43bd7129, 32'h434bd22b, 32'hc39ed761},
  {32'hc419692a, 32'h42d7e7cd, 32'h428032ad},
  {32'h44b83bcf, 32'hc2a9d90e, 32'hc20f6192},
  {32'hc51a77b1, 32'h42467289, 32'h41aeaa97},
  {32'h44f90b78, 32'h432985e5, 32'hc25beab4},
  {32'hc50beb99, 32'hc20960de, 32'hc341b433},
  {32'h44e982da, 32'h43b20acf, 32'hc3014d2f},
  {32'hc5049877, 32'hc3f1c2e3, 32'h43552f4f},
  {32'h44aa36d2, 32'h432b9888, 32'hc28e9412},
  {32'hc45a2112, 32'h422779a8, 32'h42a4a558},
  {32'h441d6054, 32'hc3976b35, 32'h440bf53f},
  {32'hc5022173, 32'h431abf90, 32'h4217c732},
  {32'h44e25a37, 32'hc357b1a4, 32'h42ecb678},
  {32'hc4894768, 32'hc29ffb96, 32'h42cebf5c},
  {32'h44b4fb4c, 32'h41a56dab, 32'h4182bb3c},
  {32'hc4b43a9a, 32'hc1134368, 32'hc2b7e91a},
  {32'h43e037b8, 32'hc3844d05, 32'h409a301a},
  {32'hc3ab80e7, 32'h43f23355, 32'h4253346f},
  {32'h43fe94d9, 32'h4325c2fd, 32'hc3d6bb2a},
  {32'hc4e08ddd, 32'h43574398, 32'h4267d110},
  {32'h44255560, 32'hc2e9e455, 32'hc2b04b5b},
  {32'hc4967fcc, 32'hc335fb77, 32'hc2a0cadf},
  {32'h4494d6cc, 32'h439dde79, 32'hc3030201},
  {32'hc4a33150, 32'h417eed54, 32'hc2b91bd2},
  {32'h451225ce, 32'h431502e3, 32'h43ce269c},
  {32'hc4b980c2, 32'hc3713738, 32'hc360c402},
  {32'h450b49b7, 32'h43892fd1, 32'hc36f39ba},
  {32'hc394d068, 32'hc3fd6c01, 32'h43bf3a2a},
  {32'h4490a6c8, 32'hc3991976, 32'h43353aa7},
  {32'hc4908e6e, 32'hc39c582f, 32'hc2ff90d1},
  {32'h44840ea1, 32'h43a13c1a, 32'hc3026026},
  {32'hc5132399, 32'h4408c2f1, 32'hc35cf684},
  {32'h44f06f1a, 32'h43853a60, 32'hc3ab05df},
  {32'hc4cc4070, 32'hc3b9c6a4, 32'hc1f05c60},
  {32'h43b79216, 32'h43049063, 32'h435f4a82},
  {32'hc3b6bc0f, 32'hc36c6165, 32'hc38b8ad9},
  {32'h44520076, 32'h43bd4fad, 32'h42c6e5cc},
  {32'hc40c6030, 32'hc328509b, 32'hc15c8c02},
  {32'h44061c08, 32'h439384b5, 32'h41b6db1e},
  {32'hc43457b4, 32'h42e25974, 32'h436856be},
  {32'h44d27539, 32'h43d5ef30, 32'h43bb9b94},
  {32'hc42a1e78, 32'h43f7743c, 32'hc3a4542c},
  {32'h44cf59f8, 32'h43c99cd9, 32'hc3bd73f3},
  {32'hc4198886, 32'hc3b16cff, 32'h412e9574},
  {32'h45137710, 32'h433e4eb5, 32'h4390c95e},
  {32'hc4cf8acb, 32'hc29eeddf, 32'hc38e2f6d},
  {32'h447928c2, 32'hc29a64df, 32'h431950a9},
  {32'hc4e41d72, 32'h43cad850, 32'h412e2504},
  {32'h451f8c34, 32'h43ac81e1, 32'h44060254},
  {32'hc5112182, 32'h430be139, 32'hc34ce3b5},
  {32'h449aea88, 32'h42ece15a, 32'hc2df35d8},
  {32'hc4b50d0b, 32'hc3a1710b, 32'hc34357c6},
  {32'h44bc80de, 32'h42b0b591, 32'hc3bd1acb},
  {32'hc4b86d9f, 32'hc1904303, 32'hc2b10b2e},
  {32'h45062188, 32'hc2e37194, 32'hc29f3eeb},
  {32'hc4caf903, 32'h42e48957, 32'hc34e54bd},
  {32'h44fb3e63, 32'h4223e492, 32'hc363c193},
  {32'hc4a27a9c, 32'h41aca78b, 32'h42e1ef7c},
  {32'h44f461af, 32'hc3d15f35, 32'h40cffa9c},
  {32'hc45066e3, 32'hc2ab2bc2, 32'h419697f7},
  {32'h44ff97af, 32'hc1be74ce, 32'h4315552c},
  {32'hc523b18a, 32'hc2e628ef, 32'h439b9aee},
  {32'h441a5112, 32'hc3098d41, 32'h44023975},
  {32'hc4e30d99, 32'hc3278afb, 32'hc2c1b9c3},
  {32'h44c88b86, 32'hc4231a1b, 32'h4255c041},
  {32'hc42172b7, 32'h435e4992, 32'hc3d14854},
  {32'h44e78786, 32'h43759d10, 32'hc37cce4f},
  {32'hc4ef1088, 32'h425d551d, 32'h42894f1a},
  {32'h4306c950, 32'h441c1a31, 32'hc41adc61},
  {32'hc4de584a, 32'h43818695, 32'h432daf71},
  {32'h44e05f34, 32'h42c5780c, 32'h431b6f07},
  {32'hc424af1e, 32'hc382d16e, 32'h43dcd51e},
  {32'h44f78ce7, 32'h42c6bf8a, 32'hc3a1d687},
  {32'hc482a92a, 32'h422c15b6, 32'h43c70fa3},
  {32'h44cf4ea5, 32'hc2142958, 32'h43c55640},
  {32'hc4f7c0f6, 32'h41dd8d3b, 32'hc24246ce},
  {32'h44bd5b61, 32'hc3438072, 32'hc21f085d},
  {32'hc50b4512, 32'hc3034ea7, 32'h42857ddb},
  {32'h44f2643e, 32'h432127e9, 32'hc1757c7a},
  {32'hc448dca0, 32'h41de2231, 32'hc2824ede},
  {32'h44fd16df, 32'h41637f03, 32'hc1b5c053},
  {32'hc4e26d40, 32'h43809ab0, 32'hc1888d3d},
  {32'h44f7234e, 32'hc3d7e18b, 32'hc32f4abf},
  {32'hc4a51762, 32'h42a0d79f, 32'hc37a633c},
  {32'h44c34b26, 32'h421a1c93, 32'hc0d311f1},
  {32'hc4483266, 32'hc385182b, 32'hc2ffe871},
  {32'h43fedc35, 32'hc2fde0ea, 32'hc35aa81e},
  {32'hc42b0459, 32'hc3d4c7ce, 32'h4398b8d1},
  {32'h44ba9185, 32'hc2296b29, 32'h42e45e0e},
  {32'hc49f8900, 32'hc27ead4c, 32'h43b90e00},
  {32'h448bc1c2, 32'h428c806b, 32'hc31fd80f},
  {32'hc4526f2c, 32'hc290f4b6, 32'h425e8a6c},
  {32'h44e6dddf, 32'hc33b6520, 32'h43a8cbd2},
  {32'hc4351401, 32'hc3865014, 32'h43ae81e5},
  {32'h44e89520, 32'h4365ae73, 32'hc295e44c},
  {32'hc500ab43, 32'h438c4174, 32'h421842ca},
  {32'h44ede0b2, 32'hc380fd09, 32'h442813eb},
  {32'hc4da5b8f, 32'h43a0aa0e, 32'hc36234e1},
  {32'h447a12ee, 32'h42d992f0, 32'hc1ca82bc},
  {32'hc52a2397, 32'hc2b3ce06, 32'hc38ae2d4},
  {32'h44e40536, 32'hc186d6a4, 32'hc34754b6},
  {32'hc50690e6, 32'hc2862ab2, 32'hc30434f7},
  {32'h44bd3b90, 32'h4384623b, 32'hc2da90be},
  {32'hc50c641b, 32'hc3ed935a, 32'h430783ee},
  {32'h440d7134, 32'h43675e06, 32'h42bbfc40},
  {32'hc4dc3098, 32'h43cfac13, 32'hc2d295da},
  {32'h449e5157, 32'hc29dd80e, 32'h419f3e82},
  {32'hc4796ce1, 32'hc338ae41, 32'h43210d8e},
  {32'h451b9921, 32'h4398cb70, 32'hc2872ae0},
  {32'hc431a286, 32'hc2b3ff5e, 32'hc2682420},
  {32'h4467aed6, 32'hc285df38, 32'hc3665966},
  {32'hc4190d38, 32'hc381abca, 32'hc4035ffd},
  {32'h44e3ccd0, 32'h42f25827, 32'hc351a04f},
  {32'hc4dec464, 32'hc1e9c52a, 32'h4134f124},
  {32'h44187e7a, 32'hc0a9cc61, 32'hc27ac2fd},
  {32'hc496f263, 32'h43ab5124, 32'h430b89de},
  {32'h44afadad, 32'h438a47a2, 32'h4203a769},
  {32'hc3b7dc57, 32'h42eda697, 32'h40f6841d},
  {32'h4460a312, 32'hc25cb7f8, 32'hc3ad9caa},
  {32'hc4a27f6b, 32'h4323ac2d, 32'h433afe40},
  {32'h4499869c, 32'h4391bca0, 32'hc3ae87cb},
  {32'hc5087675, 32'h42c3220b, 32'h4390eee4},
  {32'h44abab8c, 32'hc31dcdcc, 32'hc398f4f0},
  {32'hc4a5f928, 32'hc3032c05, 32'hc36a2b24},
  {32'h4486a821, 32'h42b83274, 32'h432ef7c8},
  {32'hc4a586cb, 32'h438594ef, 32'h42b7395b},
  {32'h44dbac44, 32'hc34cf83f, 32'h43799ccc},
  {32'hc449ef90, 32'hc2d8057a, 32'hc37c5e15},
  {32'h44336428, 32'h4353d25b, 32'hc23072a4},
  {32'hc4a4e12a, 32'h42636230, 32'hc399d593},
  {32'h450f4b60, 32'h4320f8fb, 32'hc3787648},
  {32'hc4ab567e, 32'hc3a2ea67, 32'h42814f58},
  {32'h448ac55f, 32'hc38215b2, 32'hc2c64950},
  {32'hc504ffcf, 32'hc2213c89, 32'hc236abaa},
  {32'h444dfd98, 32'hc3545951, 32'hc21fac74},
  {32'hc1dd97fa, 32'hc11a795a, 32'h423b630a},
  {32'h4509fef6, 32'h425f2645, 32'h424b9c46},
  {32'hc48f78e8, 32'h426c49fa, 32'h4274995a},
  {32'h45111b56, 32'h432809e6, 32'h42ef9353},
  {32'hc4dfb295, 32'hc22ba564, 32'hc2e53ce5},
  {32'h4513b334, 32'hc36bec59, 32'h426cdc08},
  {32'hc3ecbb10, 32'hc25f41c1, 32'h4287567c},
  {32'h4450134c, 32'hc2049a32, 32'hc171f5d6},
  {32'hc388b40c, 32'hc3008c76, 32'h43ba9127},
  {32'h440efbfa, 32'h4390231e, 32'hc3317143},
  {32'hc4e2009a, 32'hc27b454e, 32'hc2119d1a},
  {32'h43afe2be, 32'hc2650d89, 32'hc2458d33},
  {32'hc4a56fba, 32'hc381cd83, 32'hc38b69d7},
  {32'h44ac6592, 32'hc2954e8a, 32'hc2514c46},
  {32'hc411e543, 32'h43000c90, 32'hc3b03cea},
  {32'h450ed496, 32'h4124110b, 32'h4257309f},
  {32'hc4fdd6ee, 32'hc0c57a24, 32'hc351a16c},
  {32'h43c97f04, 32'hc3a4a676, 32'h436668cb},
  {32'hc4aee952, 32'hc2862557, 32'h433603f8},
  {32'h449fb7dd, 32'h4261fa63, 32'h43610c3c},
  {32'hc3a60fa0, 32'h4391a682, 32'hc2877f87},
  {32'h44726a5c, 32'hc204d7f4, 32'h4283c5f4},
  {32'hc51c3676, 32'h43458984, 32'hc315339a},
  {32'h450d0601, 32'h439783f9, 32'h42e96654},
  {32'hc3b2d065, 32'hc374974f, 32'hc1fba291},
  {32'h4389660a, 32'hc30103a6, 32'h432cdb54},
  {32'hc50b1b95, 32'h43844b0a, 32'h40e4f988},
  {32'h44ea85b0, 32'h42fa4496, 32'h431ada79},
  {32'hc4e8d038, 32'h42935779, 32'h42c37aee},
  {32'h4424bae6, 32'h41fa621e, 32'hc2d9763e},
  {32'hc49edc1a, 32'hc39c5289, 32'h435d6da0},
  {32'h4404eab3, 32'h43102978, 32'h439d7281},
  {32'h4318aca0, 32'h436237f2, 32'h434626fb},
  {32'h4410ecd0, 32'h4306114c, 32'hc361cf05},
  {32'hc4b9f99e, 32'h43d509f3, 32'hc2f6b580},
  {32'h4494c80e, 32'h43c52166, 32'hc2a4da9c},
  {32'hc4aedeb0, 32'h4272fad2, 32'hc3bd369a},
  {32'h446ad834, 32'h423e8808, 32'hc408066f},
  {32'hc50745b4, 32'hc2bf345c, 32'h431e4a0e},
  {32'h44d0c2d4, 32'hc24134d2, 32'h43697211},
  {32'hc3b6af3d, 32'h437b120b, 32'h436dddc8},
  {32'h44d703a2, 32'h42ce5ae8, 32'h421c5553},
  {32'hc4a08444, 32'h42c402b6, 32'hc431e235},
  {32'h44ef67fd, 32'h42042caa, 32'hc2f74cbf},
  {32'hc48a4350, 32'hc2c83807, 32'h41ad41d1},
  {32'h448a0e77, 32'hc1ade838, 32'hc29f7e41},
  {32'hc49eb28a, 32'hc3b09f1f, 32'hc2c1a501},
  {32'h44d0773d, 32'hc320ac2a, 32'hc3d81af8},
  {32'hc4c59310, 32'h425af7da, 32'h43dc84f2},
  {32'h444cba58, 32'hc3172254, 32'hc38c6c55},
  {32'hc42a842c, 32'hc33fdcf4, 32'hc342bf32},
  {32'h447ee822, 32'hc292577f, 32'hc38d47a4},
  {32'hc46c5c76, 32'hc343db35, 32'hc1d3582a},
  {32'h448442aa, 32'h42f403f0, 32'hc2d32a6c},
  {32'hc4bf3010, 32'h41c63f6c, 32'hc35c64d8},
  {32'h451399d7, 32'hc2a3ec20, 32'h4315f817},
  {32'hc4bb2b11, 32'hc3a789d3, 32'h43823a00},
  {32'h44dc3829, 32'hc300f7cc, 32'h4185482e},
  {32'hc4ccfb3d, 32'h439c9131, 32'h42b0df50},
  {32'h450878ce, 32'hc2e804ec, 32'h423becb0},
  {32'hc382e356, 32'hc3573637, 32'h423f4254},
  {32'hc1810600, 32'hc382c1be, 32'h429e09c0},
  {32'hc4aa9311, 32'hc2cde1d5, 32'hc323d11c},
  {32'h44cc3bf0, 32'hc260bbe7, 32'hc107c35f},
  {32'hc3b25f4d, 32'h43d94711, 32'h421426b2},
  {32'h44d32131, 32'hc389b568, 32'hc2448031},
  {32'hc37413f4, 32'hc0386c44, 32'h4256e6f2},
  {32'h44446dfe, 32'h4315c88a, 32'h4311efdd},
  {32'hc49c3d9a, 32'hc2d8f776, 32'h43015641},
  {32'h44c9982a, 32'hc32871f9, 32'h43f8d28a},
  {32'hc50dfb09, 32'h426628d8, 32'h438e831c},
  {32'h42763104, 32'hc2dfcc75, 32'hc31271a0},
  {32'hc2457ae5, 32'h43f86ed0, 32'hc3643fbf},
  {32'h448b93d0, 32'h4306c4b5, 32'hc4001820},
  {32'hc2b84b60, 32'h42a729b4, 32'h435f93cd},
  {32'hc19dd8c0, 32'h43296ad4, 32'h4313a617},
  {32'hc43c84f0, 32'hc31edd16, 32'hc2afdc9b},
  {32'h44b1b8ea, 32'hc152bbde, 32'h402cc9ed},
  {32'hc4427718, 32'hc3108d53, 32'hc1acf52c},
  {32'h448d584d, 32'hc386e862, 32'hc3c1fb74},
  {32'hc3f3fd3a, 32'hc4134cde, 32'hc1b89ef4},
  {32'h44b117ec, 32'h432bc6c3, 32'h4108aa5b},
  {32'hc33df531, 32'h41316a75, 32'h43ace303},
  {32'h43da765f, 32'hc355efd5, 32'h4336486d},
  {32'hc2d24370, 32'h43d1a847, 32'hc15a9506},
  {32'h4412e62d, 32'hc3eb3ef6, 32'hc27c82e0},
  {32'hc38a232d, 32'h433fea1a, 32'hc38d4477},
  {32'h43f988cc, 32'h432607ef, 32'hc36d60ca},
  {32'h4241018f, 32'h43b839bd, 32'hc34277f8},
  {32'h42f16110, 32'h43889eec, 32'hc30c4245},
  {32'hc4fbac94, 32'h40c63dd0, 32'h411039e3},
  {32'h4401fd80, 32'hc28a0ed2, 32'h41d8edc7},
  {32'hc41f0e42, 32'h438c5d35, 32'h436fc40f},
  {32'h44574b13, 32'hc090c094, 32'h432d26f6},
  {32'hc2a0aea0, 32'h4341ecc9, 32'hc35e310a},
  {32'h44aeca3d, 32'hc3be4064, 32'h424adb5c},
  {32'h43a01d28, 32'h43e02447, 32'hc0e4a0d8},
  {32'h44dbcbaa, 32'hc329e297, 32'hc3468b7a},
  {32'hc30f4d40, 32'hc3a33413, 32'h420e5410},
  {32'h44e9d912, 32'h422a84a6, 32'hc24688b8},
  {32'hc4ed8712, 32'h4360d808, 32'hc2c63f80},
  {32'h44fb48ba, 32'hc2e1fdbf, 32'hc19fa986},
  {32'hc3cde859, 32'hc3b93427, 32'hc32a4710},
  {32'h446f2e5e, 32'h41d7f408, 32'hc4135e6e},
  {32'h42d888e0, 32'hc279e258, 32'hc0bab475},
  {32'h448cf6fc, 32'hc39d4088, 32'h41bd68b7},
  {32'hc4c276c7, 32'h42c71c02, 32'h4329a320},
  {32'h44779d38, 32'hc23eb332, 32'hc400151a},
  {32'hc42cdf7f, 32'h428bce94, 32'hc18fe890},
  {32'h450fa63a, 32'h431662a9, 32'h430e0c4c},
  {32'hc2e64908, 32'hc32c12b9, 32'h4394232b},
  {32'h450c6b19, 32'hc3034dc4, 32'hc1aeaf76},
  {32'hc46bf28c, 32'hc34dc698, 32'h43550103},
  {32'h44040352, 32'hc1cb33f9, 32'h43b04b66},
  {32'hc470685b, 32'hc2f6d392, 32'h42117f1c},
  {32'h43734cf8, 32'h43206b16, 32'hc33f0dd8},
  {32'hc2ca0348, 32'hc317aee8, 32'h431a505d},
  {32'h44c65fa6, 32'h42caf2ee, 32'hc322a3f3},
  {32'hc352fae0, 32'h41d5dfc4, 32'hc1ef152c},
  {32'h450e58c7, 32'hc2b6515f, 32'hc317458b},
  {32'hc465d954, 32'h432460ec, 32'hc3214c2a},
  {32'h42d67828, 32'hc4314ca9, 32'h4281bae8},
  {32'hc4218fc6, 32'hc3bf8a70, 32'h42112df0},
  {32'h4504ca48, 32'hc3e196cd, 32'h42fc1d94},
  {32'hc506b044, 32'hc0fb727e, 32'h43a058bf},
  {32'h44c5667f, 32'hc266d238, 32'hc12f5bdc},
  {32'hc3a57358, 32'hc35c85c1, 32'hc33996d8},
  {32'h441822ac, 32'hc307592f, 32'h426ba40a},
  {32'hc4b21143, 32'hc32da09d, 32'h43fe5af6},
  {32'h450f6de4, 32'hc30e9ddb, 32'hc34b72fe},
  {32'hc42ba7dc, 32'h432dfb85, 32'h426f17a1},
  {32'h4522c854, 32'hc39aa958, 32'hc1da51a2},
  {32'hc4b946bc, 32'hc2656502, 32'h4273a53f},
  {32'h44c91566, 32'h41399ffa, 32'h4231fbb4},
  {32'h43164a40, 32'hc390cfd3, 32'h42dca17c},
  {32'h44261b0e, 32'hc32f82c4, 32'hc2744863},
  {32'hc39c0713, 32'hc4075892, 32'h43e44300},
  {32'h44ac3d04, 32'h41cab5da, 32'hc35f5df3},
  {32'hc456842c, 32'h40830184, 32'hc28a6069},
  {32'h4515d141, 32'hc1f38b48, 32'h4385390b},
  {32'hc44a3470, 32'h4312aa48, 32'h43c00af3},
  {32'h43cfd634, 32'h43ab0442, 32'hc210502b},
  {32'hc3cfa7a0, 32'hc3a9e9be, 32'hc33df7b3},
  {32'h41433e00, 32'h4376abed, 32'h428e69a2},
  {32'hc4a185ed, 32'h412a95de, 32'h41a909b1},
  {32'h446244f0, 32'hc305ea3f, 32'hc3749e0d},
  {32'hc3c415c7, 32'hc24d4547, 32'h433164ac},
  {32'h44d7ab89, 32'hc19a9124, 32'hc3456194},
  {32'hc4f396fc, 32'h421d5091, 32'h43081c87},
  {32'h44e7c592, 32'hc1120672, 32'hc272a949},
  {32'hc3b2039a, 32'hc3289cbd, 32'h433535bc},
  {32'h447bfd9a, 32'hc0835fc0, 32'hc2eafe21},
  {32'hc4e19417, 32'hc402e126, 32'hc23d32b8},
  {32'h44833b1f, 32'hc29ec328, 32'hc360e37d},
  {32'hc508dace, 32'h4250a86d, 32'hc3a0ac77},
  {32'h440cde43, 32'hc254bd2d, 32'hc39d4ef1},
  {32'hc4b11d72, 32'h4384346a, 32'hc1f08e42},
  {32'h450c0681, 32'hc2fac696, 32'h42786078},
  {32'hc383c448, 32'h43379f39, 32'hc39462db},
  {32'h44c8dd6e, 32'hc1532eac, 32'hc1e38484},
  {32'hc501d5d3, 32'hc06733d1, 32'h43a7469f},
  {32'h4476ca3e, 32'h429a4d3b, 32'h43bc60c8},
  {32'hc51299cf, 32'hc310c3a6, 32'h42df2d5c},
  {32'h445d1551, 32'hc3200e5e, 32'hc29bfcd3},
  {32'hc3369754, 32'hc2c97c99, 32'h41a95fef},
  {32'h449e6ead, 32'h43267457, 32'hc2be5bf7},
  {32'hc4acd046, 32'h4220d82b, 32'h43dc595b},
  {32'h44029fd2, 32'hc3aed656, 32'hc39c2fd9},
  {32'hc49fecbe, 32'h42790666, 32'hc3c45007},
  {32'h44b2f5a0, 32'h4322bb18, 32'h439f696a},
  {32'hc4b5165d, 32'hc2b9df2a, 32'hc3009993},
  {32'h43d4c444, 32'hc28ec573, 32'hc178352c},
  {32'hc3aaae5c, 32'h4408347b, 32'hc3e5ec57},
  {32'h442c4792, 32'h433033a0, 32'h4347e7e6},
  {32'hc4a18ea3, 32'hc31de923, 32'hc30c2ebe},
  {32'h4529ca24, 32'hbe81b048, 32'h43064e6f},
  {32'hc51719be, 32'hc3c73dfa, 32'hc3329739},
  {32'h435edeb2, 32'h4414e999, 32'hc40dc38f},
  {32'hc52ec1b3, 32'h42790904, 32'hc2498b17},
  {32'h4508db3c, 32'hc1f9f395, 32'hc38279cd},
  {32'hc5081b1e, 32'hc22615d0, 32'h437c935e},
  {32'h43d2a974, 32'hc2246443, 32'hc35ff4d9},
  {32'hc4e11ca7, 32'h43aefb85, 32'h4230a6b1},
  {32'h44892608, 32'hc13a3284, 32'hc288338d},
  {32'hc4bad89c, 32'h431fe01c, 32'h4339ccc7},
  {32'h45010f77, 32'h43e90453, 32'h4387733b},
  {32'hc41aa93c, 32'hc39a5165, 32'h4187ea12},
  {32'h44ccecd8, 32'h414636ad, 32'hc35c0593},
  {32'hc4154f6f, 32'h41848c46, 32'h4344b5d9},
  {32'h439be8a6, 32'h42a6278d, 32'h42b2002a},
  {32'hc4cb25e5, 32'hc279de61, 32'hc185e6d2},
  {32'h45074a4f, 32'h42d65ac3, 32'h42cef2a8},
  {32'hc510ab91, 32'h433b5767, 32'h432ab177},
  {32'h44cfa263, 32'hc34bc5d8, 32'hc38080b9},
  {32'hc50e1cd8, 32'h42bfc2cd, 32'h42f0c05a},
  {32'h45158e1d, 32'h4312d24b, 32'hc406f484},
  {32'hc4493402, 32'h41d1f982, 32'hc39a9bf9},
  {32'h44facd62, 32'h4396905d, 32'hc300f10a},
  {32'hc4206332, 32'h42a63d7a, 32'h41571128},
  {32'h44e6a45c, 32'h41b53fe2, 32'hc3355e70},
  {32'hc51ab5ef, 32'hc3db47e1, 32'h40c124b0},
  {32'h44bda0eb, 32'h432f3a11, 32'h438037a4},
  {32'hc42ed544, 32'hc2c49afa, 32'h43a01006},
  {32'hc28557bc, 32'h43b395ea, 32'h429aa88f},
  {32'hc4672fc1, 32'h436afa86, 32'h430d31a4},
  {32'h45012ec1, 32'hc2da6c0e, 32'hc379cdde},
  {32'hc4ddd233, 32'hc3366c25, 32'h42a0fd5f},
  {32'h442c3a94, 32'h42bd4eca, 32'h436e6cd0},
  {32'hc50a281d, 32'hc2a4299f, 32'hc327272b},
  {32'h446691eb, 32'h41c3bb29, 32'h428e0753},
  {32'hc51efc2a, 32'hc14e328f, 32'hc3cf1499},
  {32'h445fe892, 32'h43a36286, 32'hc352e0c3},
  {32'hc3a5f9d8, 32'h43e4f9c3, 32'hc29c3050},
  {32'h43ef393c, 32'h41b7969d, 32'h42ab42de},
  {32'hc448b6a4, 32'hc1c19bb1, 32'hc3802996},
  {32'h44ee7946, 32'h42facab6, 32'hc23f9288},
  {32'hc4c0ed19, 32'h3f9ff678, 32'hc3274fb7},
  {32'h44791d2f, 32'h43017e8e, 32'hc348b944},
  {32'hc4384dc6, 32'hc3d5c6a4, 32'h439c3abc},
  {32'h43d9dd38, 32'h42a87f66, 32'hc39264a5},
  {32'h4353c10c, 32'hc1583db2, 32'h4294b646},
  {32'h449c0801, 32'h43b0cd7a, 32'h43277ee3},
  {32'hc50f69a7, 32'h42a2960e, 32'h43ee40b0},
  {32'h44f9a17f, 32'hc2de9511, 32'hc1afcbc7},
  {32'hc4c181b7, 32'h403edc1b, 32'hc194eea0},
  {32'h4451f28d, 32'hc1c12bd8, 32'h43232003},
  {32'hc4ef017a, 32'hc3a24ceb, 32'h4324cdb0},
  {32'h44c7791a, 32'h43206f6d, 32'hc38075ee},
  {32'hc3dcc56a, 32'h4357af04, 32'hc32d7045},
  {32'h444aa5c7, 32'hc1881362, 32'h4384452e},
  {32'hc2b8cae0, 32'hc29aa50a, 32'hc30c93b0},
  {32'h42938282, 32'h4238ce7f, 32'hc40ae43d},
  {32'hc43a329b, 32'hc18d7448, 32'hc356e00f},
  {32'h43efbc24, 32'hc3401ad3, 32'h421b29cd},
  {32'hc472b743, 32'hc28f4ae0, 32'hc338aab7},
  {32'h44559cba, 32'h43164e52, 32'h42eab75e},
  {32'hc44d4090, 32'hc26d8360, 32'hc391053b},
  {32'h44f8587d, 32'hc30f3e33, 32'h4378ee61},
  {32'hc4e50558, 32'h430b41d5, 32'h435cbe59},
  {32'h4415924d, 32'h42a8965a, 32'h42d47cbd},
  {32'hc3ef00ee, 32'h43817769, 32'hc38635d4},
  {32'h45126fb8, 32'hc322e5e5, 32'h43832197},
  {32'hc4a6e87f, 32'hc32101f1, 32'hc36e7d3e},
  {32'h445bf3a4, 32'hc29bd300, 32'h431d8962},
  {32'hc507696a, 32'hc2ad1c89, 32'hc280463d},
  {32'h43d0783e, 32'hc24550c4, 32'h43e4f8ed},
  {32'hc48d1bc0, 32'hc3054c0a, 32'hc3341a37},
  {32'h4505341c, 32'hc269585f, 32'hc37a6c55},
  {32'hc4bc058a, 32'hc14f40d8, 32'h432a08ff},
  {32'h44c94c8b, 32'h436d350e, 32'h432b5dde},
  {32'hc4c0ae9e, 32'h42a8789c, 32'h4239e63e},
  {32'h44cffe10, 32'h439e0b31, 32'h42f3345f},
  {32'hc4755c53, 32'hc3297591, 32'h424fd73f},
  {32'h4458df63, 32'hc3be8829, 32'h433ddedd},
  {32'hc502599c, 32'hc42766be, 32'h41935b76},
  {32'h44a4e248, 32'h40b41b98, 32'h42d1f7e0},
  {32'h42e2c8c8, 32'h42fa58ce, 32'hc23d5a17},
  {32'h450bf39a, 32'hc1e4f66b, 32'hc28a2afa},
  {32'hc3b113d2, 32'hc35313de, 32'hc33f7a7b},
  {32'h451375db, 32'hc2c5ee11, 32'hc3c5ced2},
  {32'hc43cc4e5, 32'h4314e00b, 32'h43003b87},
  {32'hc25c3d10, 32'h43975dc4, 32'h42247b22},
  {32'hc4d95027, 32'h4214d796, 32'hc36db1e6},
  {32'hc3f951f0, 32'hc29a2645, 32'h42db1c84},
  {32'h4474330f, 32'h43a72130, 32'h43a3a2df},
  {32'h42a31c96, 32'hc2db9693, 32'hc3747c56},
  {32'h43bab592, 32'hc31084a7, 32'h437a5065},
  {32'hc4a596dc, 32'hc3d6c070, 32'hc3801c44},
  {32'h44066f7c, 32'hc246291e, 32'h43a01cce},
  {32'hc458a9fa, 32'hc395849a, 32'h4287d416},
  {32'h445ae210, 32'hc2838481, 32'h430a4e74},
  {32'hc437a490, 32'h43bea905, 32'hc207ebd2},
  {32'h44c6e0c0, 32'h43858d43, 32'h43150904},
  {32'hc420d2b0, 32'h43764b1a, 32'h4381782c},
  {32'h447b5484, 32'hc304cf5d, 32'hc0c1c3d6},
  {32'hc4bd40b1, 32'h43387c3d, 32'hc2901538},
  {32'h45084802, 32'h43e4b4d4, 32'hc30e85f3},
  {32'hc424aa08, 32'h42ccaf7e, 32'h4392fc56},
  {32'h42d532e2, 32'hc387183c, 32'h4351ff97},
  {32'hc2f03ff8, 32'h438c517b, 32'hc3817e65},
  {32'h451124fe, 32'h4371206f, 32'h42e7eb32},
  {32'hc3665f67, 32'h424fc817, 32'hc32c2922},
  {32'h44dd65be, 32'hc2eb8dc6, 32'hc2ca92c3},
  {32'hc3e3aa08, 32'hc3003e37, 32'hc3646eec},
  {32'h446cddf4, 32'h42bae2ba, 32'hc393bed5},
  {32'hc4e9846c, 32'h434ccee0, 32'hc3fb9b21},
  {32'h44dc612a, 32'h429bd807, 32'h434dc99a},
  {32'hc515bf56, 32'hc100727d, 32'h435653c5},
  {32'h44b02a94, 32'hc2ffa163, 32'hc34b4c81},
  {32'hc38f5174, 32'h42bca66b, 32'hc35e308f},
  {32'h450eb766, 32'hc3512f7f, 32'h4253c4ba},
  {32'hc49ab39b, 32'hc34cee4f, 32'hc3aece67},
  {32'h42b0e3be, 32'hc32101f2, 32'hc2e64644},
  {32'hc5091e96, 32'hc304efa5, 32'h43ca57ba},
  {32'h44e46e30, 32'hc3874c00, 32'hc2585f7c},
  {32'hc4ae1a38, 32'h4217edc6, 32'hc29bf063},
  {32'h449bdded, 32'h42e98311, 32'h42b9a2a0},
  {32'hc4b08262, 32'h43b41ebe, 32'h4376ba4e},
  {32'h42e65fb0, 32'hc349cd9a, 32'h438373b0},
  {32'hc4482a78, 32'hc3373b87, 32'h436c1f86},
  {32'h4502b97e, 32'h423d9b40, 32'h43e53db4},
  {32'hc49bac29, 32'hc389ecde, 32'h43ae93b6},
  {32'h448cbf05, 32'h4300db8b, 32'hc2b68c75},
  {32'hc4ecbbab, 32'hc35ead75, 32'h42f94c6d},
  {32'h4488500f, 32'h421a9553, 32'hc2831131},
  {32'hc5022f35, 32'h437e8154, 32'hc3a30947},
  {32'h44c02ae5, 32'h438ebbef, 32'hc2416545},
  {32'hc4b57dfe, 32'h43094413, 32'h4365b2a2},
  {32'hc2a79b99, 32'h42b5ffef, 32'h43034ae6},
  {32'hc34a7650, 32'h42bd2925, 32'h41be2b2d},
  {32'h4514bf02, 32'h4359e5a8, 32'h438c7fca},
  {32'hc50a154c, 32'h4301cc15, 32'h43132c74},
  {32'h43f76ae2, 32'hc3a338e7, 32'h4256dbf8},
  {32'h42fa1fa0, 32'h439384c2, 32'hc38a5a45},
  {32'h43b74154, 32'hc38bed6a, 32'h42c5f417},
  {32'hc314b8f8, 32'hc296d507, 32'hc2047c1f},
  {32'h4476decb, 32'hc3d601ee, 32'hc3409f81},
  {32'hc4c9c948, 32'h42e9f912, 32'hc30d93c4},
  {32'h44caaad2, 32'h42dfd1dd, 32'h4261117c},
  {32'hc41815ac, 32'hc387b146, 32'h43a46d84},
  {32'h44b9bd74, 32'h4224f157, 32'hc3d2d914},
  {32'hc51d34e2, 32'hc4166d7f, 32'hc3598ace},
  {32'h442e320a, 32'hc2a8b43c, 32'hc2bd1cd2},
  {32'hc4cd6392, 32'hc3b2b7a1, 32'h42f0796c},
  {32'h450c16fd, 32'hc2decaa0, 32'h44058e38},
  {32'hc49f9891, 32'h43408fae, 32'h430cd4c3},
  {32'h4502fe9e, 32'hc31a5106, 32'h43ab4237},
  {32'hc4afeba3, 32'h438a1b26, 32'hc31c8d99},
  {32'h44bbd7bb, 32'hc39be0a5, 32'hc31a43e4},
  {32'hc470b887, 32'h4383baaf, 32'h41c77524},
  {32'h451960f8, 32'h436f033b, 32'hc30cf046},
  {32'hc4db59f0, 32'hc3e1cc91, 32'hc284c3d1},
  {32'h4500de0f, 32'h438d1671, 32'h42c31ce8},
  {32'hc4f5b3a9, 32'h4385cd4e, 32'h43e49f46},
  {32'h43c9a6d5, 32'h438e06ac, 32'h438282f1},
  {32'hc4dd567e, 32'h42b83c00, 32'hc36c1e42},
  {32'h44ed42b4, 32'hc35e5591, 32'hc371c246},
  {32'hc4f573a1, 32'hc28df90b, 32'h41b06912},
  {32'h44f55e16, 32'hc181c10a, 32'h43208b62},
  {32'hc453ea62, 32'hc37df731, 32'hc3ac6adc},
  {32'h44250928, 32'h4394bf7b, 32'hc3a3560b},
  {32'hc4a458ca, 32'hc305ab59, 32'hc3358f8d},
  {32'h446d977a, 32'h41be0fc6, 32'h43c2e432},
  {32'hc4166544, 32'hc31a89bb, 32'h41bfe2e9},
  {32'h43dccf70, 32'h438a29ff, 32'hc3b3e713},
  {32'hc482fd2b, 32'hc3be4e5b, 32'h4381b951},
  {32'h447cc657, 32'h42a61408, 32'h43470f4e},
  {32'hc4e5424c, 32'hc28e3a55, 32'h4339f42f},
  {32'h43fefe59, 32'h438e28b4, 32'h4356b554},
  {32'hc4b781ce, 32'h42a97730, 32'h42556186},
  {32'h44ac0ee8, 32'h41d0ecef, 32'hc1cf2552},
  {32'hc459ae40, 32'hc3f90e8e, 32'h4394a506},
  {32'hc35cb8f8, 32'h437ff66a, 32'hc34137f9},
  {32'hc50a9c1d, 32'h41e57cf8, 32'hc20df93b},
  {32'h445020ae, 32'hc236f60a, 32'h42b3322e},
  {32'hc0d93650, 32'hc232720e, 32'h43858123},
  {32'h43b30a8a, 32'h432acfdc, 32'h43ebf0c4},
  {32'hc4e1f316, 32'hc2b1109d, 32'hc38b33e3},
  {32'h44924918, 32'h41d7934e, 32'h42e754bb},
  {32'hc4f1480b, 32'h43272e9e, 32'hc3261ea1},
  {32'h44cd492a, 32'hc01f6c74, 32'hc34f1758},
  {32'hc4dee00c, 32'h41192404, 32'hc3ca964d},
  {32'h44f2d5bc, 32'h42d62ae4, 32'hc344435d},
  {32'h4304d3bf, 32'h429bba1a, 32'h4334e17e},
  {32'h449a768e, 32'hc230b448, 32'hc20b14fd},
  {32'hc50aa2a8, 32'hc2b03161, 32'h42e30f0f},
  {32'hc19d9308, 32'h437319cf, 32'h4285c717},
  {32'hc3a46f50, 32'hc3889e37, 32'hc3350317},
  {32'h4457a44c, 32'hc2ae4af4, 32'h42be5afb},
  {32'hc43d3b9d, 32'hc324bcbc, 32'hc337f11d},
  {32'h44940e74, 32'hc3f4e9ef, 32'hc36429e9},
  {32'h4363fe68, 32'h41afbab5, 32'h41fa447e},
  {32'hc1d2af00, 32'h439fafc5, 32'hc3196c53},
  {32'hc4b11d70, 32'hc41827d5, 32'hc1c798e3},
  {32'h40915440, 32'h411c5e51, 32'h4328b914},
  {32'h416a1f00, 32'hc3a3cc02, 32'h434977f1},
  {32'hc2ba8a44, 32'hc235d989, 32'h43bd62f1},
  {32'hc4e8611d, 32'hc3740647, 32'hc36f3838},
  {32'h4305fdb8, 32'hc32e2dcc, 32'hc335eb27},
  {32'hc1b9aad0, 32'h4308a102, 32'h43ab93ed},
  {32'h44b64afe, 32'h43998b49, 32'hc33b2d7e},
  {32'hc4ae66c0, 32'hc203835e, 32'h42a53526},
  {32'h43edfcc0, 32'hc2517602, 32'hc1f5c2ca},
  {32'hc3e1a330, 32'hc35eb21a, 32'h43114b52},
  {32'h43f68333, 32'h4168cb78, 32'h43685f67},
  {32'hc3b56f4a, 32'h44057283, 32'h429411f6},
  {32'h445163d6, 32'hc330d355, 32'hc2cbc0d0},
  {32'hc491cf08, 32'h4337375c, 32'hc31d6a01},
  {32'h450d4c73, 32'h431ee868, 32'h43028edc},
  {32'hc505caf9, 32'h42e0c2a5, 32'h4341648c},
  {32'h4331402a, 32'h43ac8b1e, 32'hc3483ed3},
  {32'h42a6c5b0, 32'hc39bb690, 32'hc2c60473},
  {32'h43f03c7c, 32'h43d6cd3a, 32'h43c525da},
  {32'hc5006b7d, 32'hc33599bc, 32'hc3208910},
  {32'h44b28bd2, 32'hc2292aa1, 32'h43a28b1e},
  {32'hc4fb9ff7, 32'hc3bdf722, 32'h4384ba8d},
  {32'h445555dc, 32'h4217a05f, 32'h426b9e52},
  {32'hc51432f4, 32'h43a73229, 32'hc37fd1a3},
  {32'h4409acf8, 32'h4324ecc9, 32'h437bb001},
  {32'hc4ea5f2c, 32'h43f63faa, 32'hc33db9cb},
  {32'h44a4f110, 32'hc2948c97, 32'hc1a541a1},
  {32'hc3c75898, 32'hc1c7e842, 32'h42967a88},
  {32'h442ef96d, 32'h42018c45, 32'h438f766c},
  {32'hc4c0cc0c, 32'h4332e4ad, 32'h431979be},
  {32'h44280112, 32'h41ddc6b6, 32'h4218bf6c},
  {32'hc4bf95ac, 32'h425ab1ae, 32'h42179002},
  {32'h44d7ec7a, 32'hc3647646, 32'hc22c52ec},
  {32'hc512ddd0, 32'h4307637e, 32'hc283abbb},
  {32'h439430d8, 32'hc311afc6, 32'h42d055d6},
  {32'hc4a3763c, 32'h41bda482, 32'hc21551c9},
  {32'h44b1e621, 32'h43cc584e, 32'hc27a83bc},
  {32'hc4860f81, 32'hc302ce8f, 32'hc3dac725},
  {32'h44d08635, 32'hc3979126, 32'h43a03bb4},
  {32'hc4959670, 32'h4287f03c, 32'h43139b87},
  {32'h44c7a60b, 32'hc35c3ecf, 32'h434aa4dd},
  {32'hc48a2e0b, 32'hc377d6c8, 32'hc1f9118c},
  {32'h43ecd178, 32'hc1f14459, 32'hc2a3237d},
  {32'hc3a06e20, 32'hc2b18770, 32'h4378a476},
  {32'h42624e40, 32'hc34e4961, 32'h435618c9},
  {32'hc3777363, 32'h43002cd5, 32'hc0879c76},
  {32'h4427a908, 32'h4333a4b7, 32'hc26cfcd1},
  {32'hc4ddebc8, 32'h4389e5b4, 32'hc1f8758e},
  {32'h44e23d59, 32'h4325910d, 32'hc232fe99},
  {32'hc49cc8d2, 32'hc3819a33, 32'hc28b5d9f},
  {32'h44e185c8, 32'h43569c3c, 32'h4388e5bc},
  {32'hc48d0fb0, 32'hc38a6565, 32'h4298ff35},
  {32'h44085988, 32'hc3248d36, 32'h421a2a1e},
  {32'hc4ea4c88, 32'h432f56fb, 32'hc210c0a2},
  {32'h44e77d01, 32'h41caf0e2, 32'h427f94f4},
  {32'hc519b0b6, 32'h42d1c5d5, 32'hc21b5155},
  {32'h44b392f8, 32'hc2eaa906, 32'hc2094c45},
  {32'hc3d6beca, 32'h43a4f3fa, 32'hc3be7fe8},
  {32'h44892192, 32'hc2b235f1, 32'hc3a87ea7},
  {32'hc431ac1c, 32'h4371c64b, 32'h4360fdf3},
  {32'h446b849c, 32'hc2c2791a, 32'h43df064f},
  {32'hc3816414, 32'h4298edc3, 32'h42901c0e},
  {32'h440eb25c, 32'hc304fbfd, 32'h439225c6},
  {32'hc420221e, 32'h439d0194, 32'h43351fcc},
  {32'h43aa54cc, 32'h40be2340, 32'h43d0b7b1},
  {32'hc2f31d90, 32'h42aaad55, 32'hc2afa11a},
  {32'h4427ad06, 32'hc2929c00, 32'h42b7635d},
  {32'hc4a19680, 32'hc3784083, 32'hc3c48414},
  {32'h439a256c, 32'hc3c08bbd, 32'h435eba10},
  {32'hc4ad5a0a, 32'h408abab6, 32'hc380fda9},
  {32'h44e452ad, 32'hc38412c6, 32'hc361e099},
  {32'hc509ccbf, 32'hc3202acf, 32'hc39941dd},
  {32'h4395e565, 32'h4223838c, 32'h4304d959},
  {32'hc48b240a, 32'hc3b4444c, 32'hc37af82c},
  {32'h44b29c6c, 32'h4348bbcb, 32'hc2eb274c},
  {32'hc48b7f98, 32'h4320f518, 32'hc289a9b3},
  {32'h441119ae, 32'h42cbbd55, 32'h422a1f68},
  {32'hc2bd6d46, 32'h4370a859, 32'hc2a1044d},
  {32'h449ac90e, 32'hc305916e, 32'h435fa20f},
  {32'hc41c3fa2, 32'h425f3296, 32'h43891a81},
  {32'h444df3d0, 32'h4406ab99, 32'h43eebcef},
  {32'hc41a3282, 32'hc3c3b878, 32'hc2d89102},
  {32'h44196928, 32'h436198b2, 32'hc318b284},
  {32'hc4d82258, 32'hc29ac515, 32'hc376b947},
  {32'h44dbe105, 32'hc3c39e7c, 32'h4281fac0},
  {32'hc4b499ce, 32'hc2faac0d, 32'h4191c14c},
  {32'h44752164, 32'hc286c1ac, 32'h4335d5c7},
  {32'hc4965a51, 32'hc3a3073b, 32'h43274803},
  {32'h43db2393, 32'h4366bbc2, 32'h4419eea0},
  {32'hc4b0e355, 32'hc2bf8469, 32'hc3a60a60},
  {32'h4416a4b8, 32'hc3ebb184, 32'h4311ec43},
  {32'hc44d0ceb, 32'hc4065876, 32'h4264fa44},
  {32'h440776bb, 32'h43694bbd, 32'hc38db92f},
  {32'hc46e9a79, 32'hc287082e, 32'h422ed719},
  {32'h44a368db, 32'h425ea967, 32'h42eaf5e3},
  {32'hc407f875, 32'hc3912181, 32'hc315f2c8},
  {32'h448e8920, 32'hc3754e19, 32'hc38e9281},
  {32'hc4a8d585, 32'hc37c78c8, 32'hc3cec530},
  {32'h44c998db, 32'hc3cbd4f0, 32'h41854397},
  {32'hc48e8610, 32'hc2034121, 32'h4385fb65},
  {32'h44b9561c, 32'hc341b5a5, 32'hc3efc75d},
  {32'hc4ddbb59, 32'h432dff3a, 32'hc2f939c2},
  {32'h446b6f73, 32'hc20b16f4, 32'h433c188b},
  {32'hc4f2b6d4, 32'hc1cea796, 32'h42babecc},
  {32'h450fb74f, 32'hc309cf6b, 32'hc32df211},
  {32'hc4b6f1c4, 32'h43068240, 32'h43112756},
  {32'h42f22e4c, 32'hc33f8b7a, 32'h43a54097},
  {32'hc48b990c, 32'hc34964d1, 32'hc2c22a35},
  {32'h443f0c7d, 32'hc20151b7, 32'h40f50e93},
  {32'hc491a9b7, 32'hc2d9f682, 32'h423e26c1},
  {32'h43052cbc, 32'hc257aa27, 32'h42d60cd5},
  {32'hc3ecc3f6, 32'hc22ef13c, 32'h43911713},
  {32'hc30ce8e4, 32'h4378941f, 32'hc43852ee},
  {32'hc4e156e3, 32'h430d92ae, 32'h43d1230d},
  {32'h451b5468, 32'hc40fde46, 32'h4376273f},
  {32'hc39bce28, 32'hc258eea9, 32'hc20ba106},
  {32'h4499cda9, 32'h42b4a3b3, 32'hc3891377},
  {32'hc50721b5, 32'hc3967cbc, 32'h433c8859},
  {32'h43f5f18c, 32'h434b6798, 32'hc33acd44},
  {32'hc4cd80ea, 32'hc309f708, 32'h438c7eb0},
  {32'h44caf94c, 32'h43d77925, 32'hc270a722},
  {32'hc4bad724, 32'h430164d6, 32'hc2f0d6ff},
  {32'h439a6d20, 32'hc33fed00, 32'h4182f012},
  {32'hc4171696, 32'hc2761c2f, 32'h42778504},
  {32'h44ec333c, 32'hc32b445f, 32'h432dbf00},
  {32'hc5081c6e, 32'h43176bbe, 32'h43787799},
  {32'h44a42946, 32'h420f4dfb, 32'hc341febf},
  {32'hc3bc59e8, 32'hc3224730, 32'h4354e56e},
  {32'h42ec2f60, 32'h42851e9a, 32'h420dbb6f},
  {32'hc4c34036, 32'h40432aa9, 32'hc214d069},
  {32'h442bcbb0, 32'h435b3d29, 32'hc32cc51d},
  {32'hc487f4c6, 32'h42739fb8, 32'hc11912ad},
  {32'hc32b0506, 32'h436f834a, 32'h43eb3793},
  {32'hc4ebd62a, 32'h433e44ff, 32'h424c0ce3},
  {32'h43a9abff, 32'h43199432, 32'hc2eda3c7},
  {32'hc485c9a3, 32'h437e1190, 32'hc3a1ae1c},
  {32'h4505d1db, 32'hc2c2c32f, 32'h42d367b6},
  {32'hc50a05b4, 32'h42efb73c, 32'hc3360412},
  {32'h44b537f8, 32'h43a830b6, 32'hc358dadd},
  {32'hc4d8a8cc, 32'hc21110db, 32'h4312b991},
  {32'h44b77c40, 32'h423d866e, 32'hc39a316a},
  {32'hc4ec535a, 32'h41f7893b, 32'hc2cbec63},
  {32'h448e64cb, 32'h43342a71, 32'h427475fc},
  {32'hc399a456, 32'hc39d56bf, 32'h4382a2ca},
  {32'h44788854, 32'h4294f0aa, 32'hc35bb320},
  {32'hc3f0f417, 32'hc32f079e, 32'hc288f737},
  {32'h433c11d0, 32'h439e40ea, 32'h43aa6435},
  {32'hc4897899, 32'h428c8f6d, 32'hc2c68a1a},
  {32'h441a484a, 32'h43075a7a, 32'h438455dd},
  {32'hc2ce0f4a, 32'h4347747e, 32'hc3abd610},
  {32'h4475f333, 32'h43075bfc, 32'hc3238025},
  {32'hc4c0244a, 32'h437ac9a5, 32'h4340dfd4},
  {32'hc19d2860, 32'h424c1895, 32'h431a6576},
  {32'hc3d97174, 32'hc38c6f22, 32'hc1e366f7},
  {32'h4516fa0b, 32'h405fed4c, 32'hc3e06821},
  {32'hc4e180aa, 32'hc2fdc777, 32'hc2ae11c2},
  {32'h445bdefc, 32'h424b5ff6, 32'h438ac15a},
  {32'hc4cb7c36, 32'hc3790fbb, 32'hc381eaff},
  {32'h447f915f, 32'h4314eb5f, 32'hc39c7723},
  {32'hc36ef268, 32'h439a9d5e, 32'h42efe240},
  {32'h43156fc0, 32'h432043c8, 32'h430d3ffa},
  {32'hc4952058, 32'hc2d9c3c0, 32'hc3b14b95},
  {32'h451f991f, 32'hc035d201, 32'hc22438e6},
  {32'hc495d80e, 32'h4273fb2b, 32'h429050fc},
  {32'h44e207a5, 32'hc2555591, 32'h43c8127e},
  {32'hc39f94f8, 32'h42ab1a42, 32'h4138fbc2},
  {32'h436fcad0, 32'hc3a37431, 32'hc3016410},
  {32'hc4afb0c1, 32'hc1a23922, 32'hc344523e},
  {32'h43023e6e, 32'hc313b4d2, 32'h4305016d},
  {32'hc4f7a4ea, 32'h43beba93, 32'h4200cbc8},
  {32'h44583728, 32'hc3bdb837, 32'hc3a95b24},
  {32'hc4c43c60, 32'h42f4c36f, 32'hc1fd8a4a},
  {32'h44b93c6c, 32'h42210e84, 32'h43a0d9a7},
  {32'hc522bac7, 32'hc0fbcf06, 32'hc411cea1},
  {32'h450981dc, 32'h4194de88, 32'h42b38d80},
  {32'hc474d25a, 32'h43d242e6, 32'hc386dabe},
  {32'h449b7e51, 32'h4287a66d, 32'hc32048e8},
  {32'hc4b8ecf6, 32'hc393911b, 32'hc31102c5},
  {32'h436e716f, 32'hc324b103, 32'hc33e4917},
  {32'hc4465108, 32'hc221b438, 32'hc30261ed},
  {32'h44b104a8, 32'hc2d9d511, 32'hc3a97adc},
  {32'hc48d115e, 32'hc3625112, 32'h4359a7fc},
  {32'h448858d1, 32'h438b522a, 32'h43eec84c},
  {32'hc512750a, 32'hc0af66fa, 32'h43330ab2},
  {32'h44e49f8e, 32'hbebc929a, 32'hc30b2398},
  {32'hc3fd914e, 32'h4400b8da, 32'h42233b3a},
  {32'h445ef800, 32'h4152f0bc, 32'hc385ed2e},
  {32'hc46a649e, 32'h4138b5f8, 32'h42cd4660},
  {32'h45040d3e, 32'h43a6e277, 32'hc195d829},
  {32'hc38066a0, 32'hc1d4b532, 32'hc368d0f4},
  {32'h45020fc3, 32'h40b141ea, 32'hc39248b0},
  {32'hc402ca76, 32'hc32adad4, 32'hc32da282},
  {32'h44a22ff1, 32'hc3c4660e, 32'h424a871e},
  {32'hc3fd8d28, 32'h438ab916, 32'hc30fdefb},
  {32'h4505d08a, 32'hc2fea802, 32'hc3885393},
  {32'hc507861c, 32'hc16aa1c8, 32'hc2eaf020},
  {32'h4488e5f0, 32'h43337682, 32'hc2908f17},
  {32'hc4edeab2, 32'hc2223ac1, 32'hc2eab3d0},
  {32'h446bd562, 32'hc36e9976, 32'h437cd5b3},
  {32'hc4fca03e, 32'h4028b434, 32'h4310a336},
  {32'h4461f307, 32'h41cf9ee5, 32'h4421cdf7},
  {32'hc4f853ba, 32'hc3245f4a, 32'hc1c3f506},
  {32'h4512cadb, 32'h422d9a42, 32'h4230c79a},
  {32'hc2e73231, 32'h435d4cde, 32'hc31cd44f},
  {32'h4503dc50, 32'hc29d5c76, 32'h4394c24c},
  {32'hc4e77793, 32'h41fcfa1c, 32'hc2bf0233},
  {32'h44ae683e, 32'h425d32a2, 32'hc2b0f39a},
  {32'hc50378e8, 32'h435c20e7, 32'hc3154d05},
  {32'hc2156020, 32'hc3991ef4, 32'h4402e173},
  {32'hc40af62e, 32'h431f2240, 32'h42932421},
  {32'h4474690b, 32'h43ce9f5e, 32'h4334951d},
  {32'hc49db238, 32'hc315d12a, 32'h42a7df12},
  {32'h45078d03, 32'h43cebfc6, 32'h4388bf3d},
  {32'hc4063ea4, 32'hc3c6f9cf, 32'hc368af83},
  {32'h45139276, 32'hc2915204, 32'hc3848181},
  {32'hc488f004, 32'hc38b352f, 32'h433f160b},
  {32'h44141cc6, 32'h430d30fb, 32'h430ce45c},
  {32'hc3e4acaf, 32'hc373e0b6, 32'hc320b8ae},
  {32'h443ffc5a, 32'hc2f3cfdf, 32'hc3ccd9d0},
  {32'hc5098380, 32'hc39eac61, 32'h42bfad02},
  {32'h4410198e, 32'h41d2e654, 32'h4295aae7},
  {32'hc47227d1, 32'hc14e39c9, 32'h431b2aa0},
  {32'h448b8a5b, 32'hc0cdd5db, 32'hc38cd549},
  {32'hc4b08e6b, 32'h4230060a, 32'hc3121e3f},
  {32'h450c494f, 32'hc36b922c, 32'hc32fc3f5},
  {32'hc4965c24, 32'hc2d638be, 32'hc3482765},
  {32'h44e80e04, 32'hc3228acb, 32'h430608f5},
  {32'hc4990e6f, 32'hc4118f28, 32'h429689ea},
  {32'h43ccdd68, 32'h43965c8c, 32'hc3e314b6},
  {32'hc4be7dab, 32'h415e6a90, 32'hc0d4b6c5},
  {32'h451a24c3, 32'h43a7fc03, 32'hc2d8ebae},
  {32'hc45815ae, 32'h43624db9, 32'hc3555270},
  {32'hc2a500e8, 32'h428f622d, 32'h437cf195},
  {32'hc4a67222, 32'h430a05b7, 32'h4325e496},
  {32'hbf47d800, 32'hc1a2632b, 32'h431c6fdd},
  {32'hc527dd9f, 32'hc1819c48, 32'h43350cfb},
  {32'h45253ff0, 32'h428ee712, 32'h43084d75},
  {32'hc5188ced, 32'hc3239703, 32'h4283118f},
  {32'h4322b3d6, 32'hc355ec1d, 32'h421888f2},
  {32'hc497f0ca, 32'hc3ac2f33, 32'h434f38b4},
  {32'h44251d44, 32'hc34e6b9a, 32'hc2685d75},
  {32'hc362e6b8, 32'h41324f80, 32'h435df354},
  {32'h43cf5968, 32'h43c91429, 32'h43604b02},
  {32'hc50b21f9, 32'hc32417cc, 32'hc23ada4e},
  {32'h44ca0f90, 32'hc15a5a2a, 32'h42012bec},
  {32'hc497c1de, 32'hc1b916f8, 32'hc3df55d3},
  {32'h44b4714c, 32'h43ad1397, 32'hc36e692c},
  {32'hc4bcaa35, 32'h435eb3a8, 32'h4180a089},
  {32'h44c7e524, 32'hc218530c, 32'h41bddf5e},
  {32'hc48767ca, 32'hc32ab033, 32'hc3def68c},
  {32'h42ffea78, 32'h43112916, 32'hc1f21e65},
  {32'hc49f38ee, 32'hc29d2830, 32'hc279c10f},
  {32'h44a0d8c9, 32'h43a7e775, 32'hc30bef4a},
  {32'hc4d550ca, 32'h427c2be6, 32'h43abe973},
  {32'h44acfadd, 32'h43884873, 32'h4259df74},
  {32'hc4a753da, 32'h436d6c82, 32'hc25c38e6},
  {32'h45047dda, 32'hc31c7dda, 32'hc38228c3},
  {32'hc455b3f8, 32'h43166016, 32'hc41750b7},
  {32'h44c21af6, 32'hc28714e7, 32'h42fa7070},
  {32'hc5092f4c, 32'hc3603117, 32'hc35f4b65},
  {32'h440c41e4, 32'h436aa677, 32'hc32d0e88},
  {32'hc3fc7549, 32'h428967c8, 32'h4378d399},
  {32'hc34c6c07, 32'hc312fd83, 32'h43a34936},
  {32'hc3d36642, 32'h4288483a, 32'hbe6cae34},
  {32'h44846e55, 32'h40e3f004, 32'hc321448e},
  {32'hc38809da, 32'hc292d9fd, 32'h4355c572},
  {32'h439511f8, 32'hc2b0ffba, 32'hc39687e6},
  {32'hc42f176a, 32'hc303e95c, 32'hc32f2aeb},
  {32'h449aea40, 32'h43d78cd5, 32'h43bbcb0d},
  {32'hc500ea60, 32'h4387b7ca, 32'h42d514f3},
  {32'h44a2f742, 32'h42e4c787, 32'hc229a66d},
  {32'hc4d1def5, 32'hc28237a0, 32'h423821f4},
  {32'h450bab9a, 32'hc2cbd6e0, 32'h42d7e75b},
  {32'hc4a21968, 32'h4395512c, 32'h43a764f8},
  {32'h44a414a6, 32'h4272ea5d, 32'hc30aaead},
  {32'hc4bd569b, 32'h42f3cfe8, 32'hc2c1b044},
  {32'h44f91382, 32'hc3560c92, 32'hc33df69b},
  {32'hc38b6c70, 32'hc30016ba, 32'hc2bbedee},
  {32'h45074bc8, 32'h433196be, 32'h435367af},
  {32'hc4e9110e, 32'h4329e15d, 32'h432f824c},
  {32'h44fb4334, 32'hc31902fa, 32'h438487c3},
  {32'hc4831b95, 32'h4217b9ec, 32'hc1522839},
  {32'h451e73fa, 32'h431f337f, 32'h42211c48},
  {32'hc3957054, 32'hc2d92eee, 32'h42c29e80},
  {32'h445d0786, 32'h4315fbb2, 32'hc35344e2},
  {32'hc49d8764, 32'h420ab8e9, 32'h43a9cb47},
  {32'h44851e02, 32'h41506713, 32'hc2d07276},
  {32'hc4e94101, 32'hc3a2602c, 32'h430ac1ce},
  {32'h44bec5f5, 32'h41a8159c, 32'hc3cd8f4f},
  {32'hc5034ee4, 32'h439b8802, 32'h43002f04},
  {32'h44de1242, 32'hc386dd56, 32'hc40cd706},
  {32'hc4240f97, 32'hc38698ee, 32'h4254e437},
  {32'h4324e4e6, 32'h413b5d58, 32'hc31740e6},
  {32'hc519fb39, 32'h42aef769, 32'hc3c84b13},
  {32'h44ac3f24, 32'h42fa01a2, 32'hc2a9881e},
  {32'hc4ba84c6, 32'h43061ee9, 32'hc39fb7eb},
  {32'h440aacf6, 32'h42a6af96, 32'hc2188520},
  {32'hc4e8791e, 32'h43c78b47, 32'h435dbb74},
  {32'h4433f4a9, 32'hc0f9c928, 32'hc3d43bb0},
  {32'hc40c473c, 32'h43220b31, 32'hc2852c09},
  {32'h45127132, 32'h43447042, 32'h42b4210d},
  {32'hc2ba9070, 32'h40ee725c, 32'hc2ba7c5d},
  {32'h4495cfe2, 32'hc33ff66d, 32'hc2fe63a7},
  {32'hc4c75b47, 32'hc3676c16, 32'h43f5e17d},
  {32'h43f1cd87, 32'hc2200324, 32'h42e74e9c},
  {32'hc4f914ad, 32'hc3871968, 32'hc2525064},
  {32'h4459079e, 32'hc1ac9dca, 32'hc3820212},
  {32'hc4f4161a, 32'hc3a69fea, 32'h4347dc2e},
  {32'h43bd8c43, 32'h43a5b157, 32'h429a399e},
  {32'hc42e202a, 32'hc1e1d6e7, 32'h437b5f15},
  {32'h451b8183, 32'hc3a7986a, 32'hc3c700e3},
  {32'hc25d3251, 32'hc31694ad, 32'h425b1f76},
  {32'hc27792b0, 32'h42fbd3bb, 32'hc35620be},
  {32'hc4ac1f09, 32'hc29e3730, 32'h43a80775},
  {32'h44d5899d, 32'h42862c5a, 32'h40ea417e},
  {32'hc423f74e, 32'hc2ee25ff, 32'hc2be302e},
  {32'h44ffc49b, 32'hc3b21e6f, 32'hc39ff6ed},
  {32'hc4f413a0, 32'hc1c3d246, 32'h4194a15f},
  {32'h43d5b050, 32'h42dba21a, 32'h42fcbd7a},
  {32'h43b0fab8, 32'hc30c6734, 32'h43e91790},
  {32'h4511f9fb, 32'h4318e0c3, 32'hc2d2382f},
  {32'h4428b666, 32'h432eab31, 32'h431436a1},
  {32'hc457a6f3, 32'hc2ea2be2, 32'hc33c5345},
  {32'h445ad70c, 32'hc3ef8161, 32'hc3a885f4},
  {32'h41054300, 32'h43e07d67, 32'h43678566},
  {32'h4476ae9a, 32'hc3a22b98, 32'hc3b0b9f5},
  {32'hc4e1254b, 32'h439a0631, 32'hc34dcaf3},
  {32'h41bd0980, 32'h41e6dd94, 32'h44070e91},
  {32'hc3f90000, 32'hc38c4cc5, 32'hc2815fe5},
  {32'hc384f1e2, 32'hc3afbd7e, 32'hc3204f2c},
  {32'hc4ea7273, 32'h43862144, 32'hc2b0bbc0},
  {32'h44d58e5a, 32'h43240ab0, 32'hc32a6d1e},
  {32'h439ce5d8, 32'h42b72e0f, 32'h43c622ef},
  {32'h45089e07, 32'h43be1529, 32'hc323c6c0},
  {32'hc3639993, 32'hc0db4a1c, 32'hc374ae89},
  {32'h44ceb3c0, 32'hc2682197, 32'hc3395232},
  {32'hc500511c, 32'h434cf70a, 32'hc2e5e5e3},
  {32'h44d62ea9, 32'h43bcbd88, 32'hc26774a3},
  {32'hc496ab18, 32'hc32aaa13, 32'hc2a6ec5b},
  {32'h4413c890, 32'h43939f72, 32'hc319abb7},
  {32'hc484113d, 32'hc3e0fa55, 32'h41fc5189},
  {32'h44a159cb, 32'h438ce00c, 32'hc288165e},
  {32'hc4cc5ac2, 32'hbfde1ffa, 32'hc175ae1e},
  {32'h4422e8fd, 32'hc3b037d3, 32'hc2f59956},
  {32'hc404077a, 32'hc007dab3, 32'h412e95f2},
  {32'h43c0e8cc, 32'h43a351a9, 32'h42a3df2c},
  {32'hc3b7bea0, 32'hc32495ec, 32'hc39b2324},
  {32'h4490d8e3, 32'h434716d1, 32'hc2d3efe6},
  {32'hc3c22e88, 32'hc3de3490, 32'h43719014},
  {32'h448b17da, 32'h42bcabc8, 32'h436f2a7a},
  {32'hc5003c65, 32'hc317e768, 32'h4206b2b0},
  {32'h430cfbc0, 32'h42f50f04, 32'hc379eacc},
  {32'hc0b12600, 32'h42313b28, 32'hc28510d6},
  {32'h4456a601, 32'hc3515701, 32'hc3897b83},
  {32'hc3e8c3a4, 32'h43b66f2b, 32'hc30c3b0e},
  {32'h4204c100, 32'hc2d79495, 32'hc2dc7318},
  {32'hc50d25aa, 32'hc384f320, 32'h43144454},
  {32'h44a0975f, 32'hc30055c7, 32'hc350bf83},
  {32'hc43e85d4, 32'h42374978, 32'h42aa8b2c},
  {32'h449aa55c, 32'hc3422b8e, 32'hc2181c18},
  {32'hc50739ec, 32'h42e89b1a, 32'h43954436},
  {32'h4411ecac, 32'hc322078a, 32'hc23fe5de},
  {32'hc4dc0600, 32'hc28be371, 32'hc31401ee},
  {32'h448ed953, 32'hc3560c17, 32'h4390ce80},
  {32'hc4576b6b, 32'hc3cf4b27, 32'h4388373e},
  {32'h445d553e, 32'hc29befbf, 32'h435e793c},
  {32'hc50839d6, 32'h439f9c13, 32'h41e2da84},
  {32'h44a91eb7, 32'h4313d477, 32'hc2ae34e5},
  {32'hc3045a5a, 32'h4220116d, 32'h43d2143a},
  {32'h44845294, 32'h442334a4, 32'hc415a722},
  {32'hc46368ce, 32'h4234aa0c, 32'h422a73ee},
  {32'h449e45cb, 32'h4363d5ef, 32'hc316fefb},
  {32'hc4c95cf6, 32'h42a20770, 32'hc343e589},
  {32'h4483a332, 32'h42bd7552, 32'h40e6f20f},
  {32'hc5097fbd, 32'hc3587770, 32'h43a97886},
  {32'h4469e9dd, 32'hc2d962c1, 32'hc26e6d8a},
  {32'hc3fa042e, 32'h43e7a639, 32'h41aad17b},
  {32'h44168fa3, 32'hc3beeb3a, 32'h42502e52},
  {32'hc44b8499, 32'hc3892f77, 32'hc3251e57},
  {32'h44ca0473, 32'h432b0091, 32'h42e8f9cb},
  {32'hc4ce30bf, 32'hc1996914, 32'hc32f44f8},
  {32'h4420d923, 32'hc4040172, 32'h43943cee},
  {32'hc49fa42c, 32'hc30d0f43, 32'hc329fb35},
  {32'h449467b0, 32'hc39d6fe9, 32'h429a4143},
  {32'hc4a81375, 32'h43c0f7a3, 32'hc1efde7e},
  {32'h43d53042, 32'hc2d0a748, 32'h42c9d0f4},
  {32'hc2f6d8d0, 32'h42ba680b, 32'hc3be42cd},
  {32'h44d06652, 32'h441536ed, 32'hc42cffa2},
  {32'hc422fa66, 32'hc348f2b0, 32'hc07e675f},
  {32'h45029fcc, 32'h44129398, 32'h43e28c4a},
  {32'hc495a986, 32'hc344d4b5, 32'h43a5e7ea},
  {32'h44a3a4a9, 32'h43751735, 32'hc39a9ce1},
  {32'hc40e7ac4, 32'hc33becde, 32'h4300942f},
  {32'h43f407a0, 32'hc3e3e719, 32'hc32393fc},
  {32'hc526f171, 32'h41fd9031, 32'hc2d3f542},
  {32'h45097644, 32'h43873b7d, 32'h4335e152},
  {32'hc4715974, 32'h43ae01f9, 32'h42bb4638},
  {32'h4512f0b9, 32'hc3f89111, 32'hc3969550},
  {32'hc3d607fc, 32'h42be43f6, 32'hc3bd6afc},
  {32'h437ae9a6, 32'hc2619060, 32'hc34f6551},
  {32'hc51f144f, 32'hc38b2096, 32'hc34bd45c},
  {32'h4514b0ed, 32'hc3ab108e, 32'h427ed532},
  {32'hc4d4f870, 32'h43c314fd, 32'hc26db5cd},
  {32'h438b5618, 32'hc2d93700, 32'h4299d71d},
  {32'hc4a7797e, 32'h439f7043, 32'hc2e3fddf},
  {32'h44bafb97, 32'hc31fdc4e, 32'h436572aa},
  {32'hc4c89e41, 32'hc21ed041, 32'hc3b5991d},
  {32'h4507ff37, 32'hc307c522, 32'hc30ea6a8},
  {32'hc4407132, 32'hc2ef77fd, 32'hc2f0b040},
  {32'h43c06b6a, 32'hc332f997, 32'h423a3f24},
  {32'hc498d348, 32'h43898043, 32'h434831e9},
  {32'h445b509a, 32'h43949615, 32'hc38ca359},
  {32'hc4d11b2c, 32'hc154eb56, 32'h44154c36},
  {32'h4509cf43, 32'hc3e63e45, 32'hc1590989},
  {32'hc4d90914, 32'h40f75fac, 32'hc2ed9c58},
  {32'h4489bd41, 32'h4377b2de, 32'hc1cceaaf},
  {32'hc4cc3f9e, 32'hc3a247c7, 32'hc22e134a},
  {32'h44a38730, 32'h41a0a798, 32'hc2bb4ece},
  {32'hc3fbd58a, 32'h416207a0, 32'hc3dfaba8},
  {32'h44ae2d51, 32'h4309fcb4, 32'h419f0e4a},
  {32'hc4bb80d1, 32'h43b3f5bb, 32'h42aea8e2},
  {32'h45007a57, 32'hc3b24353, 32'hc3bf7a24},
  {32'hc47110e6, 32'h441080a6, 32'hc25892e1},
  {32'h42e5ada8, 32'hc22cb8e6, 32'h43b4faf5},
  {32'hc391cbfa, 32'hc3965de0, 32'hc34ccd63},
  {32'h45186524, 32'hc3cc64bd, 32'h41bcf45a},
  {32'hc4d318d1, 32'h41176b71, 32'h438656fc},
  {32'h439d7ccc, 32'h41888cd6, 32'hc33d2919},
  {32'hc4b36e27, 32'h433fb3f9, 32'hc337ec4e},
  {32'h45153d58, 32'h437eead5, 32'hc3c16c6d},
  {32'hc338cbdf, 32'h436a6288, 32'h439b1beb},
  {32'h4383b956, 32'h436528f2, 32'h43b2d55d},
  {32'hc4a8e1f2, 32'hc31131dc, 32'hc259f3be},
  {32'h44b9d778, 32'hc33902bb, 32'h423104c5},
  {32'hc4328e58, 32'h42924475, 32'h431baefc},
  {32'h44eec64a, 32'h420e74ac, 32'h4404e02c},
  {32'hc381fb30, 32'h429f7cd8, 32'hc28f6cb8},
  {32'h45043aa0, 32'hc3858ed1, 32'h435f9746},
  {32'hc51e8595, 32'h428745a0, 32'hc19cffea},
  {32'h44c11bd0, 32'h425179c2, 32'h42170f34},
  {32'hc4d76a7b, 32'h4338cb11, 32'h4308c74d},
  {32'h4485bfac, 32'h430ecf52, 32'h438b7a55},
  {32'hc4448481, 32'h42b8c622, 32'h42bbc793},
  {32'h4504b580, 32'hc323aa60, 32'hc070674f},
  {32'hc4e2fc5a, 32'hc226b24b, 32'h42c63356},
  {32'h4308513a, 32'h42bf95b1, 32'h42b5f68e},
  {32'hc42ebe66, 32'h43996851, 32'h422174c9},
  {32'h433f0bb8, 32'h41db4b56, 32'h43b0f50e},
  {32'hc4ee1ce2, 32'hc192e414, 32'h428502ff},
  {32'h44c7e93c, 32'h4376101e, 32'hc2c12fa4},
  {32'h43469a78, 32'hc22256a0, 32'h42bd6b8a},
  {32'h450097a5, 32'hc39b1b69, 32'h43803b43},
  {32'hc4d150ed, 32'hc3950929, 32'h439563a1},
  {32'h44b45a9e, 32'hc2dda556, 32'h4347095e},
  {32'hc4b0a95c, 32'h42dbf0fb, 32'hc2b35882},
  {32'h44bb3ebf, 32'hc20af5a8, 32'h42b800ef},
  {32'hc4cfe69e, 32'hc2587dde, 32'h3f84e56a},
  {32'h4407e852, 32'hc2a25638, 32'h43a1e8cc},
  {32'hc4dbb0f0, 32'h41c8faa5, 32'h439fb989},
  {32'h441d7d26, 32'h431e7f4d, 32'hc207e709},
  {32'hc3d3668d, 32'h420fa828, 32'hc20d2c18},
  {32'h442968e2, 32'h419d67f0, 32'hc359c80e},
  {32'hc4fe9600, 32'h439f5227, 32'hc15d9016},
  {32'hc335aa76, 32'hc3df9145, 32'h41b43d8a},
  {32'hc49ba6d2, 32'h4415408f, 32'hc21a9b36},
  {32'h44a6831f, 32'hc3054126, 32'hc1e7a5b5},
  {32'hc2ba0b48, 32'h43075d7d, 32'hc3378d6e},
  {32'h44f493a2, 32'hc2f8331a, 32'hc3ab15aa},
  {32'h420a6f8c, 32'h42fa995c, 32'h419d7b17},
  {32'h433e910e, 32'hc2dc94a8, 32'h42079ed0},
  {32'hc3de7334, 32'hc31af02c, 32'hc30bc833},
  {32'h442e394a, 32'h4328e8c8, 32'h41315486},
  {32'hc4d1189f, 32'h43b385d7, 32'h40de42aa},
  {32'h44a2eb86, 32'hc2c00ae9, 32'hc39c4efa},
  {32'hc3e1a844, 32'hc22755e4, 32'hc20712b5},
  {32'h43de6f88, 32'hc287d848, 32'hc3286dfa},
  {32'hc2c42a20, 32'h42a62f95, 32'h43300ef2},
  {32'h44b9c75d, 32'h42a13dc5, 32'h42fd64e3},
  {32'hc4d1e036, 32'h435822e5, 32'hc3911d92},
  {32'h4515b5f3, 32'h42b923c2, 32'hc1e3581d},
  {32'hc48fe309, 32'h43786f92, 32'h43287622},
  {32'h44c631fa, 32'h43902cb4, 32'h43448f84},
  {32'hc49c531e, 32'hc2544606, 32'hc3014bc7},
  {32'h44f0e9db, 32'h43311625, 32'h43669830},
  {32'hc3650720, 32'hc3283501, 32'h42e78df2},
  {32'h44dc96d9, 32'hc384115f, 32'hc392e9a6},
  {32'hc514f7ac, 32'hc322a108, 32'hc326b716},
  {32'h4487c355, 32'h43d6677d, 32'hc2f56e84},
  {32'hc4a799d4, 32'h42121763, 32'h427c7bbb},
  {32'h439029fe, 32'h429661f2, 32'hc3920bcb},
  {32'hc5030a73, 32'h438bcd23, 32'h43b0215e},
  {32'h43ef05b6, 32'hc2ee3e9c, 32'hc3c1bf5d},
  {32'hc5095090, 32'hc10b5ca9, 32'h43171a85},
  {32'h4509d26c, 32'hc3d5b177, 32'h43578762},
  {32'hc4a9b3dd, 32'hc28a279a, 32'hc384a171},
  {32'h44ae2a3e, 32'hc1dcd11d, 32'h42f0f074},
  {32'hc4ea698e, 32'h418e5d8c, 32'hc3ba3ca7},
  {32'h445dfc7f, 32'h42d28fbb, 32'h4334869c},
  {32'hc4e7a4e2, 32'hc203aae8, 32'h44022a33},
  {32'h44bea939, 32'hc35944c8, 32'hc34a0ac1},
  {32'hc48a79be, 32'h4381dd4a, 32'hc38d8df4},
  {32'h447b4168, 32'hc4085a77, 32'hc22b9895},
  {32'hc3814a50, 32'h42874d07, 32'hc28c7fbe},
  {32'h4491fd36, 32'hc383c714, 32'hc3ab537b},
  {32'hc3f450ae, 32'hc3178fe5, 32'hc33e333f},
  {32'h44a7bab4, 32'hc24d2108, 32'h436e3ee2},
  {32'hc0a12a80, 32'h433564e2, 32'h411bb8bc},
  {32'h4454f9b0, 32'hc0e9402e, 32'h426d5a26},
  {32'hc50cb375, 32'h431a1860, 32'hc3c7fb9d},
  {32'h44a7285f, 32'hc20fee0c, 32'hc33a4d48},
  {32'hc45f3218, 32'h42d8a779, 32'h43747be2},
  {32'h44adaef5, 32'hc2469923, 32'h440ef536},
  {32'hc5182073, 32'h4142d1d0, 32'hc35ef08a},
  {32'h44cdac03, 32'hc0335377, 32'hc180cd57},
  {32'hc4b4895c, 32'hc24d8d69, 32'h4119102c},
  {32'h420e4fc0, 32'h43a0e793, 32'hc2df2e30},
  {32'hc3c97928, 32'h438aadea, 32'h429db9fb},
  {32'h44d2a0bd, 32'h438fe82a, 32'h42ab8961},
  {32'hc48f06f5, 32'h434601f1, 32'hc3bf1e22},
  {32'h44e5e6ad, 32'hc3c84654, 32'h43851e25},
  {32'hc515464a, 32'hc3ad7ac5, 32'h433b1634},
  {32'h44e7d467, 32'hc2fafc62, 32'h4352d558},
  {32'hc4cf1ae9, 32'hc33c0dd2, 32'h432f9ce8},
  {32'h450c89ac, 32'hc3d98b99, 32'hc323c9ed},
  {32'hc4d18d3a, 32'h43646f00, 32'h4337f8ab},
  {32'h43548790, 32'hc2ee399d, 32'h43520cd5},
  {32'hc3d194bc, 32'h43efb498, 32'hc3433f33},
  {32'h40f64230, 32'hc34fc9d7, 32'h420eee92},
  {32'hc4d64900, 32'h43780bc1, 32'h426cc718},
  {32'h44446d70, 32'h42aa667a, 32'hc2f83fae},
  {32'hc4a20418, 32'h422470e0, 32'hc3301586},
  {32'h44eefb81, 32'h437a4fe6, 32'h428615b4},
  {32'hc4c88121, 32'h418830a6, 32'h43c0821d},
  {32'h44fd7504, 32'h43a90005, 32'h42eff071},
  {32'hc4e73f7a, 32'hc3310084, 32'h43e686b8},
  {32'h44ef9858, 32'h4409ad73, 32'hc37b0cd4},
  {32'hc343f000, 32'hc270827b, 32'hc2b45542},
  {32'h43e41f24, 32'hc390506c, 32'hc363918e},
  {32'hc49f5656, 32'h43e21092, 32'hc31dc83f},
  {32'h44c03ef2, 32'h42072cb7, 32'h43dfd9bf},
  {32'hc4c19fde, 32'hc205f1dd, 32'h4396a429},
  {32'h44f00d67, 32'hc2e62a6c, 32'hc2e2fe71},
  {32'hc3f09a62, 32'h42daf7b2, 32'h4355eb16},
  {32'h44f03239, 32'hc226a369, 32'h417cd1ba},
  {32'hc4846b54, 32'hc3b60cbd, 32'h4276a6a4},
  {32'h45139658, 32'h43047b12, 32'h4401ca79},
  {32'hc517a313, 32'hc22a587a, 32'h41e0c13a},
  {32'h450956e4, 32'h431d7371, 32'h432e7f0d},
  {32'hc492ab36, 32'hc38c525e, 32'hc2df0b1f},
  {32'h451d573b, 32'h43bc6d97, 32'h42dc485e},
  {32'hc485b9a7, 32'h42bfbd44, 32'hc31d2669},
  {32'h44d6a373, 32'hc1a7fc36, 32'h4331ba96},
  {32'hc4b6d02d, 32'hc2464f12, 32'hc303a941},
  {32'h44fded2c, 32'h4349160b, 32'h42c5f927},
  {32'hc4884137, 32'h40f8002e, 32'h42badce0},
  {32'h43a76a8e, 32'hc37f4cf2, 32'hc3b11fb5},
  {32'hc4f166ca, 32'hc2dd7ca9, 32'hc39495eb},
  {32'h43a800b8, 32'hc1b778f6, 32'h422ef940},
  {32'hc37f0ae0, 32'h43c0a635, 32'hc2c472f5},
  {32'h447f4362, 32'hc2a4be86, 32'h4317aae4},
  {32'hc3955924, 32'hbebe07c0, 32'hc3eb0f49},
  {32'h4508fab0, 32'h4298e1c3, 32'hc3b8451f},
  {32'hc4fab621, 32'hc3a38dfa, 32'hc2cdfa8d},
  {32'h4462b2ac, 32'hc20094b4, 32'hc2ba5489},
  {32'hc4f1e173, 32'hc2789dca, 32'h41e0766c},
  {32'h4491758d, 32'h40cbd994, 32'hc3ca9be3},
  {32'hc5012bbd, 32'h425bdbcc, 32'h430b7203},
  {32'h44bf3b95, 32'hc139d646, 32'h43032a1b},
  {32'hc40c0cfd, 32'h4377d0b8, 32'h428c805b},
  {32'h43cf25fc, 32'h4382378f, 32'h4363b2f6},
  {32'hc4a4a1e9, 32'hc29747de, 32'h425d20ec},
  {32'h4444ac6c, 32'h4360c6df, 32'hc2d5435a},
  {32'hc28c6f3e, 32'h43dac6d0, 32'hc2f19f55},
  {32'h44a8d961, 32'hc3a0d917, 32'hc3309f01},
  {32'hc4c39bfa, 32'h4350e6fe, 32'h4332b393},
  {32'h4465175a, 32'h42a1f19c, 32'hc1eca2bb},
  {32'hc490c1c6, 32'hc2329b6c, 32'h41add618},
  {32'h4441a085, 32'hc2558186, 32'hc33290ae},
  {32'hc1559302, 32'hc394adc4, 32'hc3177a6d},
  {32'h438b3d60, 32'h43050b7a, 32'hc3807a9e},
  {32'hc500a230, 32'hc36263ed, 32'h432bde44},
  {32'h44d40836, 32'h4288fd18, 32'h420d3546},
  {32'hc46872f8, 32'h43adbd59, 32'h439d4aa3},
  {32'h4504cd19, 32'h43405a78, 32'hc346aae7},
  {32'hc42116f4, 32'hc28f2183, 32'h43bbb769},
  {32'h45195abf, 32'h42c94160, 32'h438a2531},
  {32'hc501b660, 32'h43aeeaca, 32'hc173ae14},
  {32'h4503e43b, 32'h4221b63c, 32'hc35f17dc},
  {32'hc4a436f4, 32'h42b03d4b, 32'h3f675758},
  {32'h44b4385f, 32'h44025b8c, 32'hc2e8de96},
  {32'h4366a650, 32'hc31d8d46, 32'hc2a84618},
  {32'h441a9a1c, 32'h42063193, 32'hc262aecf},
  {32'hc4a31224, 32'hc334dde9, 32'hc245b8e0},
  {32'h44bc2591, 32'hc386f9bb, 32'hc318dc96},
  {32'hc4c3dfdb, 32'hc2ec1dab, 32'h42cef705},
  {32'h4507a009, 32'h420af6bb, 32'hc2c6b73d},
  {32'hc3e0710c, 32'h427f0138, 32'h425585a2},
  {32'h444be4ce, 32'hc1b51974, 32'h41f50e42},
  {32'hc4c9096e, 32'h43e8f8ac, 32'h42ba98fb},
  {32'h43fdc1a4, 32'hc2eb818e, 32'h42099974},
  {32'hc5056e69, 32'h4336e5ac, 32'h422b7a70},
  {32'h4516f7fa, 32'h431c210c, 32'hc37b1b51},
  {32'hc4ff0f6e, 32'hc1244144, 32'hc2966e15},
  {32'h44f80dc0, 32'h42f328b0, 32'hc351e340},
  {32'hc4c41031, 32'h42516840, 32'hc3697d75},
  {32'h45080b9f, 32'hc2ed5966, 32'h4312fc3f},
  {32'hc4d23743, 32'h436f61d0, 32'hc27c23a0},
  {32'h44ca05cb, 32'hc3463bb1, 32'hc32d1e58},
  {32'hc3332dd0, 32'h438c1941, 32'h439de064},
  {32'h44aa5fae, 32'hc390bcd8, 32'hc3630173},
  {32'hc456bf8e, 32'h42e01659, 32'hc39cc8d1},
  {32'h44c45926, 32'h433737cf, 32'hc320c1cc},
  {32'hc4c80df3, 32'hc373c8f2, 32'hc123748e},
  {32'h4387be67, 32'h42ed7d99, 32'hc268693e},
  {32'hc31b6854, 32'hc31f6b3d, 32'hc2371046},
  {32'h444a00a2, 32'hc3cbb3b6, 32'hc3e7fb32},
  {32'hc4c055d7, 32'hc27cc781, 32'hc306526b},
  {32'h44c23c75, 32'h430da3d9, 32'h42a2621f},
  {32'hc4f7c282, 32'h42ddf758, 32'h43434f93},
  {32'h44e3d155, 32'h43d62845, 32'hc285176e},
  {32'hc47685e9, 32'h430cef00, 32'h4363bb4f},
  {32'h44d46207, 32'h43f93ae3, 32'h427af597},
  {32'hc424425f, 32'h43afdbde, 32'hc311140c},
  {32'h450c907b, 32'h4295fc4a, 32'h431530d5},
  {32'hc40f709f, 32'h4131305f, 32'h433da1e2},
  {32'h43be105c, 32'h4360be10, 32'hc367c4db},
  {32'hc37859a0, 32'hc31dd2ae, 32'h437230e2},
  {32'h4516eb36, 32'h4298ff3a, 32'hc3854ff2},
  {32'hc47d9600, 32'hc314f0b6, 32'hc3349277},
  {32'h44bb6477, 32'hc33a438f, 32'h434f2999},
  {32'hc35dd47c, 32'h436345ce, 32'h42dd46d9},
  {32'h4526b078, 32'h43a8da72, 32'h43dd4d7f},
  {32'hc4979292, 32'h422525c6, 32'h42cc5404},
  {32'h43d0ad46, 32'hc336e801, 32'h41c4844a},
  {32'hc3ed79e3, 32'hc28e9c6c, 32'h4340c1df},
  {32'h43f4dcf0, 32'hc3296a6b, 32'hc35f5bd8},
  {32'hc4d0323d, 32'h42fb7d34, 32'hc0d33280},
  {32'h44462a6d, 32'hc23bf48d, 32'hc3bb46ff},
  {32'hc49bf63a, 32'hc18e4881, 32'h43369b7e},
  {32'h44a24621, 32'hc1ab5f3b, 32'hc345c0d5},
  {32'hc44f9c46, 32'hc34cf16f, 32'h43971be6},
  {32'h44607b6a, 32'h41bc0b6c, 32'hc0b7d098},
  {32'hc512b91c, 32'h4286e1ee, 32'hc2ad8000},
  {32'h44c2a85c, 32'hc33382fd, 32'h4364fa36},
  {32'hc50ca2c9, 32'hc38b0dd1, 32'h42f69fd3},
  {32'h4480ad2e, 32'hc28c5122, 32'hc2e2e04b},
  {32'hc4ddd995, 32'h4286bc9a, 32'hc2521d67},
  {32'h4499893e, 32'hc29f81db, 32'h429469c0},
  {32'hc32e3454, 32'h438dba4d, 32'h441908b0},
  {32'h44439fd7, 32'hc31287ae, 32'h4392e8e1},
  {32'hc51c5147, 32'h4132aa7e, 32'h434263a5},
  {32'h44183adb, 32'h42ca1b56, 32'hc358de2a},
  {32'hc4f4e9cd, 32'hc3630a93, 32'h426686ec},
  {32'h43f7ea30, 32'hc26cc174, 32'h40f11eb0},
  {32'hc4bf01be, 32'h4346d2e2, 32'h437c9716},
  {32'h44ab4d5d, 32'hc39de8d0, 32'h43265885},
  {32'hc42bfb9c, 32'hc3690cbd, 32'hc36d980f},
  {32'h4420b5ba, 32'hc34c021b, 32'hc36d4594},
  {32'hc4b5c9f8, 32'hc2a6169b, 32'h428ebeea},
  {32'h44a57a2c, 32'hc207ff82, 32'hc3a6db73},
  {32'hc4d25186, 32'h4201ac36, 32'hc3c41778},
  {32'h45236a37, 32'h4202be74, 32'hc3bec77b},
  {32'hc45d86cf, 32'h4220eda1, 32'hc3fc0065},
  {32'h44d3dec5, 32'h43a6d4f0, 32'hc2e90648},
  {32'hc4a661c7, 32'hc3ba7bdb, 32'h425b7cea},
  {32'h439b8614, 32'h43283184, 32'h42a618bb},
  {32'hc4938170, 32'h434eb194, 32'hc22394a8},
  {32'h44dc30d5, 32'hc30d5a69, 32'h42a0e8a9},
  {32'hc42da100, 32'h41a2c552, 32'h432d3400},
  {32'h436f9690, 32'hc378e7e5, 32'h4106ea4a},
  {32'hc5018a49, 32'h413f4014, 32'hc380d42e},
  {32'h42f978ec, 32'hc30141d7, 32'h430c1431},
  {32'hc4e55c5c, 32'hc33ca610, 32'h426ff15b},
  {32'h44e14a19, 32'hc2c34e7f, 32'h42192c2e},
  {32'hc50da9e2, 32'hc200540e, 32'hc3158298},
  {32'h429d0b30, 32'h42b2f8cd, 32'h4303f8e4},
  {32'hc4771d04, 32'h43820829, 32'h421a5263},
  {32'h4514e1c5, 32'h43f6cdbe, 32'hc2041388},
  {32'hc4e5cc82, 32'h43896c1d, 32'hc3c25ad9},
  {32'h4323a878, 32'hc35c0042, 32'hc386f549},
  {32'hc453f5e6, 32'hc3dc766d, 32'hc39c5dbe},
  {32'h44c28cf8, 32'hc33990aa, 32'h437c869a},
  {32'hc50376eb, 32'h431447d9, 32'hc1799b0b},
  {32'h41d28200, 32'hc2ee9246, 32'hc4387c90},
  {32'hc3b47ade, 32'h438c475b, 32'h43482536},
  {32'h44921ce4, 32'hc32cd085, 32'hc35dc83b},
  {32'hc4756630, 32'h4403dde9, 32'hc33fc158},
  {32'h4500b97f, 32'h41059dc4, 32'h429f5f4e},
  {32'hc510201e, 32'h43af0fb0, 32'h43983ab0},
  {32'h4511809a, 32'hc3cc3535, 32'hc2046cca},
  {32'hc4d4bdad, 32'hc2c27d01, 32'h43b36714},
  {32'h444831b8, 32'h41f8041c, 32'h42d03b33},
  {32'hc18e4150, 32'hc32e186e, 32'hc1cc118b},
  {32'h450f3e7c, 32'h4344452d, 32'hc2ba696a},
  {32'hc4b18135, 32'h43e53f2c, 32'h437a8eb8},
  {32'h450a631d, 32'hc2948213, 32'hc39df909},
  {32'hc37efbb0, 32'hc418089f, 32'h434fcd60},
  {32'h44ee55e7, 32'hc3ab4d13, 32'h438a64f6},
  {32'hc4c32924, 32'hc344b0a4, 32'hc2daa06b},
  {32'h442a67bc, 32'h43e7ba17, 32'h43bc9f33},
  {32'hc3938470, 32'hc2a392bd, 32'hc28d7bd1},
  {32'h4425971a, 32'h43c2eeea, 32'hc308fe17},
  {32'hc37057ac, 32'h444a77bf, 32'h43696da9},
  {32'h4364f318, 32'hc34b00ec, 32'hc3664455},
  {32'hc4f83807, 32'h42eaa1bc, 32'h43d8c416},
  {32'h449fe2dd, 32'hc3241dc2, 32'h4345f333},
  {32'hc4c6191b, 32'h43a03919, 32'hc334bfc1},
  {32'h450ed3f2, 32'h43276892, 32'hc20b4d15},
  {32'hc4c8c410, 32'hc39cd12d, 32'h42fce557},
  {32'h451d4944, 32'h42bc8a28, 32'hc39496af},
  {32'hc41b1d27, 32'h439eea95, 32'hc3a90e81},
  {32'h44e39364, 32'h4301f329, 32'h432a9750},
  {32'hc4c85a84, 32'hc220ce98, 32'h43baa8bf},
  {32'h4495debf, 32'h41fdfaba, 32'hc38839ef},
  {32'hc4eb7e74, 32'h40b9f894, 32'hc311bd9a},
  {32'h44a81ed0, 32'hc1cb23dd, 32'h438ef7a5},
  {32'hc38225d8, 32'h43f254e2, 32'hc316433c},
  {32'h44dc1002, 32'h4290fad6, 32'h4109e6eb},
  {32'hc40361fa, 32'h42bdb475, 32'h429c3824},
  {32'h443ec0ab, 32'hc38405aa, 32'hc3830380},
  {32'hc4a3a2ef, 32'h43cb47a6, 32'h42480cb6},
  {32'h4502c536, 32'h40c4b88c, 32'hc24c0c2a},
  {32'hc16e1900, 32'h43563759, 32'hc3658a89},
  {32'h44167eca, 32'hc18d7692, 32'hc1c4bbca},
  {32'hc49618ee, 32'hc2916dc0, 32'hc374e076},
  {32'h44bfeac2, 32'hc2b452b3, 32'hc2f4c7f5},
  {32'hc4e51b0c, 32'h42d8ac59, 32'hc361bba5},
  {32'h435a00b0, 32'h43b793c4, 32'h439437ca},
  {32'hc4df2dc2, 32'hc3348552, 32'hc326e40e},
  {32'h43842a58, 32'h42236851, 32'h4273a541},
  {32'hc4f9c65b, 32'hc39d3083, 32'hc3a052cc},
  {32'h43ca2da8, 32'h43865c71, 32'h443336d2},
  {32'hc4e73e72, 32'hc3242620, 32'hc2c5cc50},
  {32'h43ad67a2, 32'h427aea80, 32'hc2e2366a},
  {32'hc4c30a66, 32'hc2a75894, 32'h437f832a},
  {32'h44bd4956, 32'h4413c26f, 32'h4397ee8f},
  {32'hc43834e6, 32'h4272961e, 32'h439501d3},
  {32'h43ba1928, 32'h435d2ff2, 32'h435f967f},
  {32'hc42ecd5d, 32'hc2f784f4, 32'h3fd63763},
  {32'h443410da, 32'h43ca8904, 32'hc250adfc},
  {32'hc4aa7167, 32'h440a7606, 32'h411a66a7},
  {32'h44eb7839, 32'h431b268b, 32'h4393c0af},
  {32'hc5074b3f, 32'h42d59214, 32'hc3430611},
  {32'h4492fd9b, 32'hc2324121, 32'hc27d79f3},
  {32'hc51f8f76, 32'hc39570b9, 32'hbd3fe300},
  {32'h43d3f3d0, 32'h4247d90e, 32'h421600ea},
  {32'hc4237448, 32'h432e690b, 32'hc2de9669},
  {32'h43c2f9d8, 32'hc2a1f64c, 32'h43c18c7e},
  {32'hc480e5b0, 32'hc2c0cc3f, 32'hc3a42ec0},
  {32'h4400f1f6, 32'h4366aa9a, 32'hc26dde49},
  {32'hc4883bf0, 32'h43a53108, 32'h42c9a270},
  {32'h44dcc976, 32'h43dd851c, 32'h42823c41},
  {32'hc441c7d9, 32'hc381ad03, 32'h4306e05e},
  {32'hc4eb2cdf, 32'hc2778876, 32'hc3028c6b},
  {32'h449168bc, 32'h42956db1, 32'h42a2f451},
  {32'hc479cf9c, 32'h424022a9, 32'hc3ebde2c},
  {32'h450324dd, 32'hc2ebca85, 32'hc2910dab},
  {32'hc4686708, 32'hc36d6ffb, 32'hc34b99a4},
  {32'h4482869b, 32'h41de5651, 32'hc3c0c099},
  {32'hc4456a5d, 32'hc35799f7, 32'hc2d0e4b6},
  {32'h44bc79be, 32'hbf8f1e10, 32'h426c2163},
  {32'hc4a47b68, 32'h43a7f454, 32'hc30e04a0},
  {32'h448afe5a, 32'h441eac9d, 32'h433e25da},
  {32'hc50729ec, 32'h43839693, 32'hc34d3e5a},
  {32'h444dec08, 32'hc2f95986, 32'h43a38e62},
  {32'hc4eb3ba0, 32'h420daaca, 32'hc3b2f283},
  {32'h44e4490e, 32'h439076ba, 32'h43005d39},
  {32'hc4c43d49, 32'h42f4a60c, 32'h43ac04ae},
  {32'h44b8bbca, 32'h41ead7e4, 32'h43db4102},
  {32'hc50e83bf, 32'h41b3589d, 32'hc382d886},
  {32'h447f5702, 32'hc3a2a60a, 32'h430b1396},
  {32'hc3dceaea, 32'h42d760d4, 32'h438115c9},
  {32'h447a171c, 32'h4259e22b, 32'h430d2ad9},
  {32'hc453cb00, 32'h42f508af, 32'hc1c47614},
  {32'h44ce94f0, 32'h422632e2, 32'h430ea8b8},
  {32'hc40e3135, 32'h4303982d, 32'hc1d968cd},
  {32'h44cc7752, 32'h42cdbf67, 32'hc2db6793},
  {32'hc4281838, 32'h43913272, 32'hc3c014bc},
  {32'h44e76f0f, 32'hc1e8998e, 32'hc29862c7},
  {32'hc4de43ec, 32'h438867b5, 32'hc2f7ece7},
  {32'h451a6123, 32'h4358e8e8, 32'h4283cc7e},
  {32'hc48596bf, 32'hc2fb374b, 32'hc3bf076c},
  {32'h450adf4c, 32'h439f0dfc, 32'hc2e2f66c},
  {32'hc4fdd83f, 32'hc095f172, 32'hc3d3260c},
  {32'h4473f3fb, 32'hc38b735e, 32'h439d93df},
  {32'hc4f97819, 32'h43d53877, 32'hc391ef66},
  {32'h43b744c8, 32'h4221728f, 32'h43591b9e},
  {32'hc4ec1ab7, 32'h435dddff, 32'hc1d6bbdc},
  {32'h449b2d42, 32'h43374396, 32'hc291fb71},
  {32'hc4e9cca4, 32'hc0156468, 32'h437dcc3e},
  {32'h447ef7f3, 32'h427df842, 32'hc300cc34},
  {32'h41ec9787, 32'h4292ae8d, 32'hc3a59805},
  {32'h44ba926f, 32'h43927356, 32'hc236eef7},
  {32'hc5126b92, 32'hc2606087, 32'h4358bf63},
  {32'h45088606, 32'hc2cbab04, 32'h43d53fe8},
  {32'hc3b753e8, 32'hc255a6b2, 32'h43816f26},
  {32'h443f0b85, 32'h437da307, 32'h4385feaf},
  {32'hc4cd1f6c, 32'hc35f72fe, 32'hc1e7ce66},
  {32'h44c13344, 32'hc1942a57, 32'hc32a9b8d},
  {32'hc47deec6, 32'h42f07dbe, 32'hc28dccab},
  {32'h45049080, 32'h4381068d, 32'h43294f7c},
  {32'hc4eaec1e, 32'hc2a169a4, 32'hc390ac15},
  {32'h450b5641, 32'h43ce9d76, 32'h40e5ff06},
  {32'hc42a40fe, 32'h425cdee3, 32'hc21f8a1d},
  {32'h44c32641, 32'hc2c4176a, 32'hc35e2c2d},
  {32'hc505fa9b, 32'h43a1fc62, 32'hc2e9659e},
  {32'h44f53d21, 32'hc1f2a2d8, 32'h43409089},
  {32'hc3684bac, 32'h4261003c, 32'h436a31eb},
  {32'h45069b9e, 32'h42ac9df3, 32'hc23d5d1c},
  {32'hc47d3598, 32'h4348079c, 32'hc3b161a3},
  {32'h448a97fa, 32'h43bf5115, 32'h430ca73e},
  {32'hc4db7c08, 32'hc3e962f8, 32'hc37ad8e3},
  {32'h45086700, 32'h43a80f89, 32'hc3e4b49b},
  {32'hc4df0cd9, 32'h429105b8, 32'hc34bb38b},
  {32'h42470880, 32'hc27e929e, 32'hc1e832bc},
  {32'hc4851c46, 32'hc2c266e5, 32'hc30b0d9b},
  {32'h44eb0e12, 32'hc3a0e8d0, 32'h437896ee},
  {32'hc3d5c2e0, 32'hc298c81e, 32'h4370a353},
  {32'h451c317c, 32'h424fcaeb, 32'h4204a15f},
  {32'hc5065e2c, 32'hc3585386, 32'h43881892},
  {32'h44984e7e, 32'hc3396342, 32'hc3e5a31c},
  {32'hc36a8470, 32'h4309b0d1, 32'hc37186c1},
  {32'h441eff36, 32'h43b5efcb, 32'h43527fba},
  {32'hc41cc2b9, 32'h43791e98, 32'h42d550c5},
  {32'hc0ec5c00, 32'hc2c5addf, 32'h431aa4cd},
  {32'hc4a1487c, 32'h42c60d3a, 32'h43a11132},
  {32'hc34365f0, 32'hc35b792b, 32'h423c647b},
  {32'hc3cae168, 32'h422c70f3, 32'h41c5e6ef},
  {32'h45020f06, 32'h439653ce, 32'h43a8c260},
  {32'hc493e5b8, 32'h43c44967, 32'hc1a08dc1},
  {32'h44b40bc8, 32'h4384a2cf, 32'h42818b23},
  {32'hc4a19507, 32'hc38ce287, 32'h43763bb4},
  {32'h42c562a8, 32'h41a70e59, 32'hc24efa6e},
  {32'hc3251350, 32'hc3321981, 32'h43c9891e},
  {32'hc2c5734a, 32'hc2fce4d6, 32'h42c57cc4},
  {32'hc48ce0ef, 32'h43699e00, 32'hc37ec607},
  {32'h44fe4eb8, 32'h41855ad4, 32'hc3b2b9d4},
  {32'hc3b9e0c0, 32'h4343c4c3, 32'h421e4aa0},
  {32'h44fba6b2, 32'hc3761fb0, 32'h43ba9c13},
  {32'hc48b71ec, 32'hc058e588, 32'hc31da924},
  {32'h44ccfc86, 32'h42933690, 32'hc2127ca4},
  {32'h4324abf0, 32'hc2d4b996, 32'h432e0587},
  {32'h45135c32, 32'h4316340b, 32'hc2b2a787},
  {32'h438572ba, 32'h4354145e, 32'h41227f02},
  {32'h43f12675, 32'h40a41696, 32'h43158230},
  {32'hc3ecae66, 32'hc4037ebb, 32'h4390cce2},
  {32'h44a7da00, 32'h43850021, 32'h43c21270},
  {32'hc3af9b1f, 32'hc379f7e3, 32'h433d7d5c},
  {32'hbf9d1600, 32'hc32dc1e4, 32'h430e4a33},
  {32'hc444e322, 32'h42004c76, 32'hc057c8ac},
  {32'h449f497f, 32'hc2a4086a, 32'h42e212e7},
  {32'hc5001ddb, 32'h42fbb4a5, 32'h43063853},
  {32'h44f5103d, 32'h43b8856c, 32'hc2fd1c74},
  {32'hc41b48ca, 32'hc1b5962d, 32'h43ab3433},
  {32'h44972e0b, 32'hc38238f4, 32'hc241aea6},
  {32'hc4960657, 32'h43987c40, 32'h424beefe},
  {32'h43b5938b, 32'h4343155d, 32'h42fd96ec},
  {32'hc4a6fab5, 32'h43dd760e, 32'h43854d6b},
  {32'hc37bae2e, 32'hc2197936, 32'hc2096474},
  {32'hc4639c4d, 32'h42e5f2eb, 32'hc3834794},
  {32'h442a56e6, 32'h43033747, 32'hc36af076},
  {32'hc20fae80, 32'h4329a0ce, 32'h439215fc},
  {32'h4451a180, 32'hc21bb0ea, 32'hc2e10801},
  {32'hc48c4cba, 32'h43c64f10, 32'h417f7423},
  {32'h453333d0, 32'hc1df3262, 32'h43abf63e},
  {32'hc50e5a14, 32'hc2273ecc, 32'h43a6fddb},
  {32'h44350d23, 32'h42c53c14, 32'hc300311a},
  {32'hc488c5df, 32'hc3b2dae4, 32'h4387120f},
  {32'h430c16a0, 32'hc333dc9d, 32'hc2fac389},
  {32'h42a8ef90, 32'hc31a2ed2, 32'hc32e9674},
  {32'hc2d9e994, 32'h42a4dc31, 32'h42a1401a},
  {32'hc4a8f21e, 32'hc3185f03, 32'h41f26726},
  {32'hc2564920, 32'hc24d1637, 32'hc2ccccd5},
  {32'hc3991fe0, 32'hc288100f, 32'hc38226c0},
  {32'h43ddb804, 32'hc24a708b, 32'hc1de066c},
  {32'hc3034e6c, 32'hc2069b9d, 32'h4340ca93},
  {32'h43565540, 32'hc2b29aec, 32'h42d656f9},
  {32'hc4cc9011, 32'hc2d2c20c, 32'h42846dd1},
  {32'h44362ccc, 32'hc3afac9b, 32'hc397270c},
  {32'hc4ff9fd1, 32'h4185b90c, 32'hc38f7cf9},
  {32'h44f4b140, 32'hc31cd628, 32'hc35c2585},
  {32'hc4d8d0be, 32'h43237660, 32'hc2342575},
  {32'h43f765b8, 32'h4396aa15, 32'hc322e3ac},
  {32'hc4afc736, 32'h43bf4a4f, 32'hc2e0bba0},
  {32'h440b154f, 32'hc0a94b66, 32'h42c67de2},
  {32'hc4f86ffa, 32'hc34f08d8, 32'hc30b8309},
  {32'h45017973, 32'hc385d7c7, 32'hc07f4e94},
  {32'hc41a87f0, 32'hc2b59c92, 32'h41eb1e26},
  {32'h4511b7e7, 32'hc362ef60, 32'hc398196f},
  {32'hc507380b, 32'hc361cefd, 32'hc38368eb},
  {32'h43563e70, 32'h430de809, 32'hc36c5077},
  {32'hc35043d4, 32'h438b200f, 32'hc349f5f9},
  {32'h449a2004, 32'hc2ed071f, 32'hc1c8cf78},
  {32'hc48b4654, 32'h42f041ac, 32'h43082cac},
  {32'h4413fc99, 32'hc287532c, 32'h42c9c8df},
  {32'hc4a9b214, 32'h432fa256, 32'h4402c6d6},
  {32'h44d9ec5a, 32'hc2f4ddf9, 32'h43ac6b17},
  {32'hc487a512, 32'h43385ec7, 32'hc280fc7c},
  {32'h43ed46e8, 32'h4381513c, 32'hc1c30eb0},
  {32'hc4e21770, 32'hc3923845, 32'h420fd286},
  {32'h44faa079, 32'h4397bd68, 32'hc395ac2a},
  {32'hc4bf1abd, 32'h43d70791, 32'h4208b6ae},
  {32'h44b883f0, 32'h430157ec, 32'hc3904902},
  {32'hc4a9cd9b, 32'h43426d07, 32'h425c272b},
  {32'h44957da5, 32'hc2a69c15, 32'hc31a8ace},
  {32'hc4adb441, 32'h4323a5ea, 32'hc3071e3a},
  {32'h446c8088, 32'h43144e96, 32'h42a09d82},
  {32'hc4a1b6ca, 32'hc3bf19da, 32'hc31a9adb},
  {32'h448d9970, 32'h4291e526, 32'h43c492d0},
  {32'hc4bc0572, 32'h424e8d8a, 32'hbf75e155},
  {32'h44f26dce, 32'hc30aa8b7, 32'h434320b0},
  {32'hc49ac446, 32'h431b4d87, 32'hc31e46e2},
  {32'hc26ec842, 32'hc3c4d0a5, 32'h42ab8df2},
  {32'hc4fd7b5d, 32'h434fd002, 32'hc339d6b8},
  {32'h44ad5e78, 32'h42d1e450, 32'hc3940eec},
  {32'hc523015d, 32'hc0d179b4, 32'hc3202672},
  {32'h437c4962, 32'h4325654d, 32'hc30f75be},
  {32'hc40f20ec, 32'h4360fe10, 32'hc33b1c94},
  {32'h44cd63e4, 32'h42b450b5, 32'hc2d1d90b},
  {32'hc4cb7d75, 32'h42df9d86, 32'h43671611},
  {32'h44f5088b, 32'h42ab6cd8, 32'h4354f2a5},
  {32'hc498ae0e, 32'h43b4e9df, 32'hc218d10a},
  {32'h4361ef31, 32'h41d4744e, 32'h43b6ef2b},
  {32'hc3c908a0, 32'hc299045a, 32'hc389ee5f},
  {32'h44b9e971, 32'h4300eb32, 32'hc2dd7ad6},
  {32'hc4ca0974, 32'h42bd04b5, 32'hc1407580},
  {32'h44f091b7, 32'hc146d8c7, 32'h43bd7d68},
  {32'hc42825af, 32'h43713d94, 32'hc27973ff},
  {32'h44f4551e, 32'hc3a6b5d4, 32'h44137ad0},
  {32'hc363f930, 32'h4315d485, 32'h42c6843f},
  {32'h4500c247, 32'hc3c7c1a6, 32'hc297871f},
  {32'hc4d4be85, 32'hc3a80a15, 32'hc396b818},
  {32'h4450fd02, 32'hc3996e62, 32'hc3362937},
  {32'hc4751591, 32'h438776a8, 32'hc349e740},
  {32'h45018633, 32'h43c4cfca, 32'hc3549e3a},
  {32'hc4c90c98, 32'hc33be20d, 32'hc3ae61fc},
  {32'h44776e57, 32'h42cfb24a, 32'h43c1926e},
  {32'hc483acb9, 32'hc35cc7fe, 32'h42ee12b0},
  {32'h44509ccc, 32'h43280873, 32'h439703e3},
  {32'hc4512d8a, 32'h43b5ab39, 32'h42c28f4b},
  {32'h450062ce, 32'hc13b306e, 32'h4373b371},
  {32'hc4e2103e, 32'hc269c729, 32'h428c3272},
  {32'h4323bc73, 32'h43837f84, 32'hc39ba2c7},
  {32'hc46f8bda, 32'h42ffc1f8, 32'hc38fdde2},
  {32'h43af0c9d, 32'hc358adae, 32'hc2c6e308},
  {32'hc4913864, 32'hc2ee80b0, 32'hc36a605c},
  {32'h439bdf83, 32'h4389d91d, 32'hc21fac25},
  {32'hc4c8338a, 32'hc2bc52d2, 32'h42944009},
  {32'hc2c35660, 32'h4048339f, 32'hc31e2fc2},
  {32'hc51200ef, 32'h435349aa, 32'h441011f0},
  {32'h44e7feba, 32'h42ba7809, 32'hc1cefe99},
  {32'hc41cf8f9, 32'h429be5a1, 32'h430fd50e},
  {32'h45022325, 32'h432b37b4, 32'h419fd643},
  {32'hc43b561e, 32'hc40319f6, 32'hc374e405},
  {32'h4470834a, 32'h43070837, 32'hc35a24b2},
  {32'h4287062c, 32'h42e1d1db, 32'h431f8e78},
  {32'h4416e544, 32'h4371b7f4, 32'hc34a4739},
  {32'hc506b554, 32'h4345989c, 32'h43fac892},
  {32'h43e70bac, 32'hc23481a1, 32'h44091163},
  {32'hc508933c, 32'hc403459c, 32'hc293cf7b},
  {32'h445e5ab9, 32'hc00c4fd1, 32'hc39d2017},
  {32'hc2d47f28, 32'h4321a6c5, 32'h429ba31e},
  {32'h4497f0b0, 32'hc38126bc, 32'h41d26089},
  {32'hc4d4db78, 32'hc3178c9b, 32'hc28efde6},
  {32'h43c74054, 32'hc354e589, 32'hc2e64a7c},
  {32'hc4ed6c8c, 32'h42fbb527, 32'h42e9fb9a},
  {32'h44c8abec, 32'hc206bc7a, 32'h43690e4a},
  {32'hc504b553, 32'h43045801, 32'h420fe121},
  {32'h444a5818, 32'hc1def844, 32'hc33b0402},
  {32'hc4b0034c, 32'h43362d2c, 32'hc38b0e2a},
  {32'h44b814cc, 32'h42998be4, 32'hc36e8193},
  {32'hc3d23ca0, 32'h425401e3, 32'hc2d4927e},
  {32'h449cb493, 32'h43a0a016, 32'h431157da},
  {32'hc46b2362, 32'hc39f956f, 32'h42ac8e3a},
  {32'h4488371e, 32'h437af556, 32'hc266bcb6},
  {32'hc4693dbc, 32'hc2170f55, 32'hc31cd7f5},
  {32'h44db08ec, 32'hc30cbd4c, 32'hc38d9228},
  {32'hc4ebdab0, 32'hc2734535, 32'h43071319},
  {32'h44cf08f5, 32'hc27165c4, 32'hc12a9354},
  {32'hc5157d13, 32'h42a2c88e, 32'h42eed71b},
  {32'h42317760, 32'h43850f6a, 32'h44291a56},
  {32'hc4e3e0fb, 32'h40c4a474, 32'hc21ca4ff},
  {32'h44e0987f, 32'hc358db80, 32'hc27e5ce2},
  {32'hc50456f3, 32'h43f163fa, 32'h429d5119},
  {32'h44538010, 32'h43868c14, 32'hc30b77a9},
  {32'hc364b58f, 32'hc290cbe6, 32'h43d23020},
  {32'h44c4b298, 32'hc2247e8e, 32'h43075fa7},
  {32'hc50158f0, 32'hc372acce, 32'h42e800e7},
  {32'h44718a8d, 32'hc43bf484, 32'h43be02ea},
  {32'hc4f6982d, 32'hc18a8044, 32'hc3739f68},
  {32'h44d5778b, 32'hc30778b9, 32'h40aa7f79},
  {32'hc3d84c78, 32'hc3755576, 32'hc3cad748},
  {32'h44ff311f, 32'hc3426f59, 32'h428cd1f2},
  {32'hc4111b88, 32'hc29086bb, 32'h42cb8128},
  {32'h4511e13c, 32'h41219584, 32'h43378f7e},
  {32'hc4d38448, 32'hc330bb79, 32'h43392117},
  {32'h444dcb20, 32'hc3b6cff9, 32'h42214764},
  {32'hc4a562d6, 32'h4262526d, 32'hc31e8f93},
  {32'h4435fa2e, 32'h43c60335, 32'hc147fc92},
  {32'hc43b44b4, 32'h435c6b05, 32'hc2883575},
  {32'h44b73d81, 32'hc3805089, 32'h43babebd},
  {32'hc4da9ef5, 32'h4290b5ac, 32'hc3e4c42c},
  {32'h4461e403, 32'hc307013b, 32'hc34ca468},
  {32'hc43ccce6, 32'hc2c87469, 32'hc1a1741a},
  {32'h43646488, 32'hc2124d80, 32'h432a4bff},
  {32'hc4140aac, 32'hc302a036, 32'h429713ac},
  {32'h44f710c0, 32'h43b3a5ce, 32'h433bc874},
  {32'hc40613f0, 32'hc35883cf, 32'hc3333678},
  {32'h43ed7141, 32'h42e13485, 32'hc12328b6},
  {32'hc3b3c4e8, 32'h42225596, 32'hc4102872},
  {32'h4492303f, 32'h4353328b, 32'h41f6c7bf},
  {32'hc4cffbf8, 32'hc38af848, 32'hc31d8b2c},
  {32'h44700873, 32'h440f8c11, 32'h43cdd608},
  {32'hc4ae555e, 32'h429e90c7, 32'hc20be95a},
  {32'h44092ac0, 32'h424178ae, 32'h433db58b},
  {32'hc41a8299, 32'hc2e84dd4, 32'hc36875f1},
  {32'h44e8057d, 32'hc308e58d, 32'h4340300e},
  {32'hc4157861, 32'hc40a922b, 32'hc260326f},
  {32'h43a626b6, 32'hc34059be, 32'h425b63c5},
  {32'hc4e4acb8, 32'hc3ca1f99, 32'hc4032067},
  {32'h449ad6d8, 32'hc3f717b1, 32'h43dc85e7},
  {32'hc36a154e, 32'hc2dc0bd2, 32'hc2fc3fbd},
  {32'h450be907, 32'h4393fa8a, 32'h438433cb},
  {32'hc452952e, 32'hc3269106, 32'hc364542b},
  {32'h4447f2fb, 32'hc3b8ee78, 32'h4386f932},
  {32'hc3cd69b8, 32'h42cdec86, 32'h43830e40},
  {32'h43361220, 32'hc2457be5, 32'hc360fc0f},
  {32'hc4cd4519, 32'h4359e33e, 32'h425925d9},
  {32'h45138db0, 32'hc2fb6f55, 32'hc38bde5a},
  {32'hc45a5d0f, 32'hc306c901, 32'hc0a34fb1},
  {32'h44e8a277, 32'h43e64424, 32'hc2996b50},
  {32'hc4f5f91a, 32'h4281081e, 32'hc2b691a0},
  {32'h44e25e6a, 32'hc27ec19a, 32'h4316cf9a},
  {32'hc4c7d546, 32'h4304b304, 32'hc0b58e72},
  {32'h44636f9d, 32'hc2e08972, 32'hc3dabff3},
  {32'hc4c940c0, 32'h43269294, 32'h4338b31f},
  {32'h44aafbec, 32'hc325c615, 32'h4303c5c3},
  {32'hc44bccc7, 32'hc34af131, 32'hc2c352b2},
  {32'h4468a5b1, 32'hc3d9b0ae, 32'h42dc5f46},
  {32'hc447caf8, 32'h4343b406, 32'h43e46893},
  {32'h433f4f1e, 32'h423f06dc, 32'hc3dbe655},
  {32'hc46e95fa, 32'h426602e1, 32'h43c458a6},
  {32'h438b99dc, 32'h43448e35, 32'h42a16a6e},
  {32'hc5173832, 32'hc355018b, 32'hc3861af2},
  {32'h44f34fc1, 32'h439b9b58, 32'hc1420a88},
  {32'hc4dc3f15, 32'h42917a52, 32'h43c64a1d},
  {32'h44867157, 32'h43402476, 32'h43a1fc54},
  {32'hc4ddf289, 32'hc0b96d74, 32'hc2cd712d},
  {32'h44f2ec78, 32'h4303fe7a, 32'hc30e9256},
  {32'hc4975652, 32'hc3598a73, 32'h43d4efd1},
  {32'h45105502, 32'h413047a7, 32'h4303de9a},
  {32'hc515e046, 32'hc23eeb7c, 32'hc25add4d},
  {32'h450d55c6, 32'hc2cf366b, 32'h43999f17},
  {32'hc4bed5dd, 32'h43008acf, 32'h43420194},
  {32'h428710d0, 32'hc40c08cb, 32'h4313e158},
  {32'hc500c867, 32'hc2a87bfb, 32'h42f4bbf8},
  {32'h44c0cca8, 32'hc3927801, 32'hc31e6e75},
  {32'hc52026b7, 32'h428e0d31, 32'hc386c547},
  {32'h437b2860, 32'h42c0492b, 32'h44229de8},
  {32'hc516f25e, 32'hc3661cb1, 32'hc2cfe479},
  {32'h4455b408, 32'hc12bab3b, 32'h43996ac7},
  {32'hc483a138, 32'h43a6d4bc, 32'h433cd205},
  {32'h42e5c7c0, 32'h42959ec0, 32'h438e132c},
  {32'hc50fa308, 32'hc21cefcd, 32'h43d91db1},
  {32'h4422a4a8, 32'h41b671ce, 32'h429ba0e2},
  {32'hc42a35a4, 32'h409552fc, 32'h43061fd7},
  {32'h4514a84d, 32'hc3974f63, 32'h43960ce5},
  {32'hc2c3b300, 32'hc3ac37b1, 32'h42cbdb2b},
  {32'h43a0597a, 32'hc2fe5924, 32'h41fdfc47},
  {32'hc5057ae1, 32'hc2c8a0be, 32'hc1fafc47},
  {32'h445ae3d0, 32'hc2e3ffcf, 32'hc40add8f},
  {32'hc4183844, 32'h42dffb40, 32'h43070129},
  {32'h44f65a7a, 32'hc3b8c082, 32'h4373ad64},
  {32'hc4a862dd, 32'hc2ed49a9, 32'hc33daa0c},
  {32'h4409d8d8, 32'h431526e5, 32'hc3ad4d08},
  {32'hc4025cac, 32'h439c8c35, 32'hc3aa4634},
  {32'h44e4988e, 32'hc2db28a8, 32'hc2e5aa06},
  {32'hc4577df2, 32'hc32267f5, 32'hc3a4564a},
  {32'h44dd0afd, 32'hc25b06cc, 32'hc3e67a13},
  {32'hc451dbc8, 32'h43019e0a, 32'hc2afec89},
  {32'h4508a457, 32'hc37dc27f, 32'hc3df4d74},
  {32'hc4f648b2, 32'hc2bd06f2, 32'hc2b33acf},
  {32'h4502d16a, 32'h42c9b0cc, 32'hc31538e9},
  {32'hc4640344, 32'hbdb14b00, 32'h42e1d27f},
  {32'h44c11e7a, 32'h42def2fb, 32'h4319219e},
  {32'hc3973aa0, 32'h43788ec6, 32'hc31a7555},
  {32'h44ece7e9, 32'h4116fe00, 32'hc39564c9},
  {32'hc4f1f265, 32'hc22f3346, 32'hc2696b72},
  {32'h43bfe86c, 32'hc2fcc671, 32'hc3ec072f},
  {32'hc4924f28, 32'h42a13020, 32'hc27de580},
  {32'h44bdd1fa, 32'hc30482a1, 32'h41f39f3b},
  {32'hc4edc7e7, 32'hc2f94cb1, 32'h41dd10f8},
  {32'h44aa08cb, 32'h42ef1d4c, 32'hc384ff7a},
  {32'hc40d61ec, 32'h42f733a6, 32'h436323a2},
  {32'h44ba4241, 32'h4292de74, 32'hc2efffda},
  {32'hc3f20db0, 32'h430048e8, 32'h43622912},
  {32'h450b59e6, 32'h43de1b58, 32'hc33dd376},
  {32'hc4416588, 32'hc317848c, 32'h43160480},
  {32'h44ea7e63, 32'hc36059ed, 32'h43c5b090},
  {32'hc3165240, 32'hc2754c9a, 32'h4262560c},
  {32'h4494f4da, 32'hc360ad09, 32'h427a5ec8},
  {32'hc45a4b7b, 32'hc2b41ad5, 32'hc0e4a730},
  {32'h44d0fbf2, 32'hc2cfb86c, 32'h4292eb8c},
  {32'hc4c3625e, 32'hc2343d77, 32'h4333b26c},
  {32'h44515e8c, 32'h42138df1, 32'h4102cf88},
  {32'hc4a51469, 32'hc316d132, 32'hc3ef939e},
  {32'h43c92878, 32'hc3620997, 32'h43bf9a51},
  {32'hc4b24855, 32'h438b34fb, 32'hc2ede153},
  {32'h44ffb6a6, 32'h43e36e8d, 32'h44004b8c},
  {32'hc4d63e98, 32'hc2e097c8, 32'h42a21754},
  {32'h4303a590, 32'hc2bb0acd, 32'hc36f41f4},
  {32'hc50c3150, 32'h42aa1039, 32'hc3a58d42},
  {32'h45088258, 32'h42e2eff8, 32'h43095496},
  {32'hc48f5528, 32'hc295f3b7, 32'h4113651e},
  {32'h449a1e2a, 32'h438168ed, 32'hc198d5d4},
  {32'hc308ced0, 32'hc403025e, 32'hc36dcb00},
  {32'h43263710, 32'hc345f4c7, 32'h425e3161},
  {32'hc4fdfa00, 32'h43b827b8, 32'hc3dedb5b},
  {32'h440be608, 32'h424dc488, 32'h439f80b2},
  {32'hc3ae424c, 32'h4254e6fd, 32'hc363f65e},
  {32'h44c6835e, 32'h430ade78, 32'h42cbe3cf},
  {32'hc50eb739, 32'hc33ad69a, 32'hc21656d1},
  {32'h4445a980, 32'hc4200ff6, 32'hc39c6f79},
  {32'hc464e572, 32'h4310cbf2, 32'h429ed75e},
  {32'h44869a3b, 32'hc305dbea, 32'h43bb038c},
  {32'hc2995cc8, 32'h431f9697, 32'hc3914b15},
  {32'h447417dc, 32'hc3695aaf, 32'h421f4eaa},
  {32'h43831ebf, 32'hc1130bab, 32'hc3643f34},
  {32'h442b5ba0, 32'hc134864b, 32'hc31e78d6},
  {32'hc4fcfc58, 32'h42a7b0cc, 32'hc38540f4},
  {32'h437f03e0, 32'hc2743f84, 32'hc274a02b},
  {32'hc49c5c0a, 32'hc209cf82, 32'h435f4943},
  {32'h44343f3c, 32'hc32bc406, 32'h428b5152},
  {32'hc4e047ae, 32'hc3a26a84, 32'hc366a303},
  {32'h450bccd1, 32'hc327cf93, 32'hc13845ba},
  {32'hc50efd9e, 32'hc2148e41, 32'h431a8ccd},
  {32'h44e4af80, 32'hc2bbbb54, 32'hc2af6df6},
  {32'hc4b2788e, 32'hc2eab15a, 32'h4304949c},
  {32'h45146184, 32'h42699ace, 32'hc33b264a},
  {32'hc502eea4, 32'h43a41038, 32'h414297e1},
  {32'h443546ae, 32'hc4218796, 32'hc33999ed},
  {32'hc48abb34, 32'h42dc347f, 32'h435ab444},
  {32'h4505588f, 32'hc352547d, 32'h4382b22d},
  {32'hc4f5c564, 32'hc344af5c, 32'hc3bc1eba},
  {32'h450be626, 32'hc2380dd5, 32'hc3a145e5},
  {32'hc4f00cb1, 32'hc33a477c, 32'h42a488b0},
  {32'h4434a06e, 32'h42792b2f, 32'h431e4433},
  {32'hc482c89b, 32'hc3c14f5b, 32'h43297b7b},
  {32'h4508b4d4, 32'hc1a41e12, 32'hc39508e3},
  {32'hc4a2f42a, 32'h43af383e, 32'hc392fcd8},
  {32'h44b61056, 32'hc2233d2d, 32'h4129b38a},
  {32'hc4e2b77c, 32'h439f04c8, 32'hc2077720},
  {32'h44b4785c, 32'h3da64d40, 32'hc3a8dc34},
  {32'hc50479d7, 32'h42d0981e, 32'hc3664910},
  {32'h44129e5e, 32'hc1eaa1b2, 32'h42977316},
  {32'hc4d2e2f7, 32'hc39369ca, 32'h43392148},
  {32'h44f47f5e, 32'hc1829161, 32'hc3084032},
  {32'hc4d3a97b, 32'h4299ee08, 32'h434e0296},
  {32'h447e0f84, 32'h405198be, 32'hc28739ac},
  {32'hc4a7349e, 32'h435f511a, 32'h43ba4a2d},
  {32'h44f0e852, 32'hc18645d4, 32'hc31b9628},
  {32'hc48ef07e, 32'h42f14729, 32'hc20d5349},
  {32'h43d12f4c, 32'h438b3cc5, 32'hc2ce71dd},
  {32'hc4278154, 32'h41d1f8b4, 32'h43050284},
  {32'h44472f0e, 32'h41493340, 32'hc29ea6a8},
  {32'hc3de614e, 32'h43b576c1, 32'hc31a6a32},
  {32'h43fdde78, 32'h423068d6, 32'hc239b5fa},
  {32'hc4e42208, 32'hc2bac29f, 32'hc249b662},
  {32'h450a0949, 32'hc2f2d230, 32'hc3962f2b},
  {32'hc432e21a, 32'h43a83ae6, 32'h42d50df3},
  {32'h44240bdb, 32'h430584e7, 32'hc39c0106},
  {32'hc4bb8825, 32'h434b3309, 32'h4430f679},
  {32'h4504ac16, 32'hc3c7486b, 32'h4362c228},
  {32'hc3c7a3ec, 32'hc28754b7, 32'h430aae69},
  {32'h44a1434f, 32'hc1ba3525, 32'hc2a4e34c},
  {32'hc495b29e, 32'hc3a045da, 32'hc28a883f},
  {32'h44ce3312, 32'hc2dce968, 32'h41a551d2},
  {32'hc42a898e, 32'hc290d4b1, 32'h42e4d9c6},
  {32'h421a3260, 32'h42264453, 32'hc3d57a8d},
  {32'hc4a54dde, 32'hc2285699, 32'hc3a92dc9},
  {32'h44a28b49, 32'hc2a8fd24, 32'hc3c1ebba},
  {32'hc4a4d212, 32'h4322acd0, 32'h439d19d6},
  {32'h4482ec4f, 32'h42452e05, 32'hc3d36976},
  {32'h42ddcbb0, 32'h441b74db, 32'hc20d4a0e},
  {32'h439756c4, 32'hc2c9a4f0, 32'hc2d1140e},
  {32'h44dccacc, 32'h439522da, 32'h429e68c8},
  {32'hc4a4ce9e, 32'hc1e57a82, 32'hc2ed8491},
  {32'h44331034, 32'h431471df, 32'hc390bae8},
  {32'hc509d984, 32'h43a49b58, 32'h439507d8},
  {32'h4420b4be, 32'hc2b1bee6, 32'hc381edf2},
  {32'hc4c7cb01, 32'hc328594b, 32'hc3541911},
  {32'h4480324c, 32'h43846119, 32'hc29e010e},
  {32'hc4047a56, 32'h433507af, 32'hc376feb3},
  {32'h44bc08b8, 32'hc3547b36, 32'hc23b5528},
  {32'hc3599e87, 32'hc3abfdba, 32'hc39c924f},
  {32'h44e73c37, 32'hc32d3cb3, 32'hc31c98e9},
  {32'hc4f96f7e, 32'h4297b85a, 32'hc1af8048},
  {32'h441a1314, 32'hc2c4121e, 32'hc2c464c7},
  {32'hc3fdf4d8, 32'hc25fa696, 32'hc377e689},
  {32'h449db684, 32'h4315a51f, 32'h4242d32c},
  {32'hc4290a32, 32'hc3b1b3a8, 32'h429c6a5d},
  {32'h437c9b98, 32'h427a8647, 32'h42c1f0d1},
  {32'h3f9ec100, 32'h434bee73, 32'hc2e421ac},
  {32'h44a73186, 32'hc395521e, 32'hc1a31b1e},
  {32'hc4decbb6, 32'hc20e99ed, 32'h43942e86},
  {32'h4426def2, 32'hc3a755c5, 32'hc2ab66f2},
  {32'hc3a8df80, 32'h4196c477, 32'hc3a2164a},
  {32'h44abd413, 32'h4324f976, 32'hc2fbc021},
  {32'hc4570bed, 32'h41b8fded, 32'h439afeb3},
  {32'h44a3ff01, 32'hc253586c, 32'h421f66ba},
  {32'hc38c7727, 32'h436791b2, 32'h438f3c89},
  {32'h45029f88, 32'h424edf84, 32'hc267f01b},
  {32'hc3b88ef4, 32'h42dba2ed, 32'h42990271},
  {32'h442d680e, 32'h43286adc, 32'hc2b0f931},
  {32'hc43668e4, 32'h4370000b, 32'hc2132c1c},
  {32'h44932495, 32'h42e85b23, 32'h437a37ee},
  {32'hc35ba3ec, 32'hc36c582a, 32'hc38885e6},
  {32'h4447b037, 32'hc21ae593, 32'h43644c1d},
  {32'hc4e4df73, 32'h41f23f5a, 32'h42879aa5},
  {32'h42199148, 32'h4227268c, 32'h40c4c1f4},
  {32'hc3f69046, 32'h436eb13d, 32'hc2113b36},
  {32'h448ea132, 32'hc26d717e, 32'h4257b03b},
  {32'hc4bd3608, 32'h4406fe14, 32'h43fd136b},
  {32'h44fcb2aa, 32'h42784ec4, 32'h43a3abe7},
  {32'hc35e5c70, 32'h4373924c, 32'hc3672a7c},
  {32'h43a6ac24, 32'hc3b2d960, 32'h4307622c},
  {32'hc32d8810, 32'h439d98fd, 32'h43e5fdaa},
  {32'h4501d656, 32'h42ccc361, 32'hc3e7e12b},
  {32'hc4b2d0a4, 32'h41d04833, 32'hc2a43670},
  {32'h44905b54, 32'hc326fb12, 32'hc33577d7},
  {32'hc438dd4c, 32'h431abbfd, 32'h42ee6044},
  {32'h436cb470, 32'hc3a7358b, 32'h4402fb43},
  {32'hc468c4ac, 32'hc3e0320f, 32'h43f47c8d},
  {32'h450d508a, 32'h42b6ae99, 32'h428c0795},
  {32'hc3eda888, 32'hc2d4ac10, 32'h4302da9c},
  {32'h44b67318, 32'hc20cd079, 32'h42abcdde},
  {32'hc4c58f5d, 32'h43d33006, 32'h4277e5ed},
  {32'h45067611, 32'hc2bcc464, 32'hc2577f1f},
  {32'hc4a64d79, 32'hc30a68fe, 32'hc156ef2d},
  {32'h4509ea67, 32'hc101e29c, 32'hc2308fda},
  {32'hc41b4010, 32'hc14ffd98, 32'h418b044e},
  {32'h449e1f4e, 32'h422bff34, 32'hc3c4d93d},
  {32'hc420d648, 32'hc30b8360, 32'h41f639a6},
  {32'hc1a56ef0, 32'hc3190b01, 32'h3ffff5aa},
  {32'hc3a271f3, 32'hc1ba1d6b, 32'hc1d7a961},
  {32'h44c7f7e8, 32'h439c40f0, 32'hc352b220},
  {32'hc3b011c6, 32'hc1d480a9, 32'h43d7dc94},
  {32'h44a79a72, 32'h426b4f83, 32'hc3b785b0},
  {32'hc3123973, 32'hc32d16d9, 32'h4337c5d9},
  {32'h44788faf, 32'h4415dd3e, 32'h43884812},
  {32'hc3b206b0, 32'h4297cffa, 32'h4313579e},
  {32'h440f9a7f, 32'h43605780, 32'h419fa1f1},
  {32'hc36ce538, 32'hc35de57a, 32'hc16b4782},
  {32'h4468a5da, 32'h4404fa6e, 32'hc2aa9945},
  {32'hc44afe15, 32'h423ca57c, 32'hc3530071},
  {32'h441c7c11, 32'h42789b01, 32'h43b4c30e},
  {32'hc511b3ea, 32'hc3a53480, 32'hc312c07f},
  {32'h45004d5d, 32'hc36de130, 32'hc1b92800},
  {32'hc5108e36, 32'hc291d055, 32'hc3b448b7},
  {32'h44ae1828, 32'h435f3c06, 32'h433ee06d},
  {32'hc4e1b13e, 32'h438ae6b6, 32'hc40759ea},
  {32'h44c7ed23, 32'h43ba0ae4, 32'hc20d2dd4},
  {32'hc3efe7b7, 32'hc3830f7e, 32'h401cccda},
  {32'h444966e0, 32'hc3470e5a, 32'h42900470},
  {32'hc4adf5b8, 32'hc37dc1d1, 32'hc2e59f2d},
  {32'h450bd3f0, 32'hc34dd7e0, 32'h42a3ec4d},
  {32'hc44086f8, 32'h4369d419, 32'hc38df376},
  {32'h44bf08c8, 32'h43296a57, 32'hc365c4f8},
  {32'hc5032b6b, 32'h438bb15a, 32'h42315acb},
  {32'h451f20ca, 32'h41a98036, 32'h432d0a8f},
  {32'h4344bbd8, 32'h43164c1e, 32'h4343b03a},
  {32'h44b78dfb, 32'h439f1159, 32'hc3769f2b},
  {32'hc48ebd37, 32'hc3000828, 32'hc25df890},
  {32'h44361b03, 32'h43223227, 32'h435417da},
  {32'hc35bcefa, 32'hc33e19b1, 32'h3f933e72},
  {32'hc24453e0, 32'hc3102cc4, 32'hc299062c},
  {32'hc50a15ef, 32'hc2c5dbca, 32'h430364b0},
  {32'h44fbaf8a, 32'hc19e3a93, 32'hc2e24881},
  {32'hc3da9c4f, 32'h43c64e41, 32'hc323e3a2},
  {32'h441d838a, 32'h420d4351, 32'h4388965e},
  {32'hc4617e26, 32'h43944e5f, 32'hc28703d4},
  {32'h44447868, 32'h42cc95e0, 32'h43367691},
  {32'hc3363e00, 32'hc2bd1f20, 32'h42362b14},
  {32'h44c43aa1, 32'h43df3ff7, 32'h42f358d2},
  {32'hc4d4073d, 32'hc30f426c, 32'h4289868a},
  {32'h44d8bce6, 32'h43fee233, 32'h433223b2},
  {32'hc4a9b77d, 32'hc3930cc9, 32'hc13b9958},
  {32'h448d568d, 32'h436f0dc2, 32'h41151744},
  {32'hc4fda998, 32'h4370900a, 32'h42336829},
  {32'h44c7aa98, 32'h434255a6, 32'hc30600f5},
  {32'hc45b657e, 32'hc3654fc1, 32'h4312cf8b},
  {32'h448410f8, 32'h434adad7, 32'hc326462b},
  {32'hc49e5476, 32'h4253c72f, 32'h422c9769},
  {32'h4448ed6e, 32'h4382e893, 32'h4391ee1f},
  {32'hc4973f8c, 32'h409cc902, 32'h43b1fe1e},
  {32'h44af810c, 32'hc3d28d0e, 32'h4007da14},
  {32'hc4916b6a, 32'h4396c946, 32'h43ead6ef},
  {32'hc38c1f54, 32'h42a608f8, 32'hc286aef1},
  {32'hc4d46f08, 32'h43e7aea6, 32'h4374d794},
  {32'h44212bd1, 32'h4352b4eb, 32'h43bb4459},
  {32'hc4b446b0, 32'h438b722b, 32'h439cb79a},
  {32'h42f0d710, 32'hc31309f8, 32'h4239d95d},
  {32'hc4a1549c, 32'hc3306f06, 32'h427108c9},
  {32'h4484f72c, 32'h432407e0, 32'h43205d8b},
  {32'hc4d0b684, 32'h416ec314, 32'h438ef182},
  {32'h44105e5c, 32'hc3e88a17, 32'h4397ec75},
  {32'hc42ee02a, 32'h4165cf94, 32'h432eb7ad},
  {32'h43a07065, 32'h434f8ad4, 32'h4298f2cc},
  {32'hc3ccf6d8, 32'hc2360c84, 32'h4321a997},
  {32'h44eafc60, 32'hc2349a24, 32'h43ca814e},
  {32'hc4e9245c, 32'h42889a5b, 32'h4277380a},
  {32'h44a8dc7e, 32'h42029e7e, 32'h427daac9},
  {32'hc4141eec, 32'hc3bab7fe, 32'hc1257bf2},
  {32'h44cce6b2, 32'h4387de4f, 32'hc2b86a51},
  {32'hc4620c28, 32'hc26e4aff, 32'h4352be94},
  {32'h44acfe2a, 32'hc346f07e, 32'h42995b7e},
  {32'hc4d5d7d6, 32'hc29e613f, 32'hc3a745ef},
  {32'h44f87dd1, 32'hc32f310c, 32'h429fdafc},
  {32'hc4de1852, 32'hc2ea3f43, 32'hc29147d0},
  {32'h44181cde, 32'h431d8025, 32'h43901595},
  {32'hc4994b41, 32'hc39b5818, 32'hc3ba82ac},
  {32'h45130b0f, 32'h4336cea2, 32'h4288b57f},
  {32'hc42ffb05, 32'h428b367d, 32'h438fd290},
  {32'h4382c39f, 32'hc1c37b74, 32'h41be2820},
  {32'hc4aca07d, 32'hc3b2b8cb, 32'h428b4871},
  {32'h437cd2b0, 32'h420f3095, 32'hc20151a5},
  {32'hc205d83a, 32'h434a1ccd, 32'hc3743bf0},
  {32'h44ddd331, 32'hc2849b67, 32'h429a1800},
  {32'hc483000e, 32'hc3a224f4, 32'hc317e378},
  {32'h44a91ee4, 32'h436acd8d, 32'hc2cdccec},
  {32'hc4c74223, 32'h412b6d30, 32'hc1f22b94},
  {32'h450e540a, 32'h436b725b, 32'hc22c201a},
  {32'hc48e0cfc, 32'hc2521706, 32'h42ca1531},
  {32'h44ce4fd1, 32'hc28175f2, 32'hc19a3e58},
  {32'hc2f96f75, 32'h430c470c, 32'hc28b5308},
  {32'h44601808, 32'h3d20ae00, 32'h43b8d476},
  {32'hc45feb63, 32'h438f832e, 32'h432e6993},
  {32'h4499c2df, 32'hc1908638, 32'h42ccdf7b},
  {32'hc49c1806, 32'hc3353361, 32'h439d1d62},
  {32'h43e112a2, 32'h44177d46, 32'h42486b63},
  {32'hc439d439, 32'hc311c9c0, 32'h428f2ef5},
  {32'h4495abf5, 32'hc36884f5, 32'hc1e8603d},
  {32'hc460bd45, 32'hc2735266, 32'hc3504f29},
  {32'h44dcd824, 32'hc34f1ae9, 32'hc30ac599},
  {32'hc3e0b1d4, 32'h4375b88f, 32'h429ae8a1},
  {32'h44fc2ac4, 32'h41aa096e, 32'hc356e785},
  {32'hc516e500, 32'h43660acd, 32'hc30e4ad2},
  {32'h4511041d, 32'h425e9487, 32'h43a3bd83},
  {32'hc5075a58, 32'hc356b643, 32'hc333fc9d},
  {32'h43671710, 32'hc0da1b18, 32'h43bcc08e},
  {32'hc45403f4, 32'h434a50f4, 32'hc317718f},
  {32'h4355dc5c, 32'hc36975bf, 32'hc3ef1065},
  {32'hc4f47fca, 32'h424dd056, 32'h43b71136},
  {32'h4449abf8, 32'hc2d3d885, 32'h42de76f5},
  {32'hc4017480, 32'hc17581b0, 32'h43b12542},
  {32'h44b1c1f8, 32'h43486a34, 32'hc13f9e65},
  {32'hc423bafd, 32'h43048bc8, 32'h4355a636},
  {32'h43eedd71, 32'h428e22de, 32'hc2f1a297},
  {32'hc4e21f62, 32'h4299e3c5, 32'hc2b71a9d},
  {32'h4503ea59, 32'hc302c705, 32'h42f2ef0b},
  {32'hc4a69339, 32'h4380d456, 32'hc29d28a3},
  {32'h442f148c, 32'h42d1bf88, 32'hc311a173},
  {32'hc4c66989, 32'hc2fa98ab, 32'h42e3aa6e},
  {32'h445bbe74, 32'h438e8a1b, 32'h438f3025},
  {32'hc4a957b1, 32'h43037301, 32'h43c8929e},
  {32'h447972c0, 32'h43569a01, 32'hc35ca0db},
  {32'hc48557c6, 32'hc3b21c89, 32'h437197a8},
  {32'h43a42c98, 32'hc2bd9bc6, 32'hc390f9df},
  {32'hc504fe6e, 32'hc3d9f1bc, 32'h437bcc06},
  {32'h44cb59ba, 32'hc1a1145f, 32'hc30aea98},
  {32'hc4dffdf9, 32'hc398d307, 32'hc1c57403},
  {32'h44dee192, 32'h434c0bdf, 32'h434791d6},
  {32'hc48bb351, 32'h419d8982, 32'hc36968f5},
  {32'h45099ff0, 32'hc32c85a0, 32'h43522c07},
  {32'hc37b4db0, 32'h430af311, 32'h4369756b},
  {32'h42f0769e, 32'h42e57d62, 32'h4286abc0},
  {32'hc40acd0c, 32'h42791b33, 32'h424563b0},
  {32'h4432e6f8, 32'hc348f149, 32'hc2505c96},
  {32'hc506225e, 32'hc2628695, 32'hc28b71ce},
  {32'h4438aef2, 32'h42fe29e9, 32'h42b4db34},
  {32'hc4e07b23, 32'hc34d2919, 32'h43fe9706},
  {32'h4478c411, 32'h42f7db3b, 32'hc2a195d2},
  {32'hc4e6cc15, 32'h4343cd10, 32'hc1fad0e7},
  {32'h446a0280, 32'h431a24e4, 32'h43f06664},
  {32'hc4c67a78, 32'hc38d5845, 32'h43562067},
  {32'h45186e3d, 32'h43525afb, 32'h438d5f3f},
  {32'hc4a8bf70, 32'h42a50fd8, 32'h4325cb8d},
  {32'h44713f94, 32'h433eb83f, 32'hc264ad89},
  {32'hc4314d42, 32'h42da236b, 32'hc30087b3},
  {32'h4518c2a4, 32'h4378f771, 32'hc2a8db96},
  {32'h436f6ff8, 32'hc3594585, 32'h43995092},
  {32'h44c6a71a, 32'h433b4e33, 32'h432c6ba4},
  {32'hc3e243c1, 32'h44119e2e, 32'h42136563},
  {32'h4513a9b1, 32'hc242b7d5, 32'hc3a69d49},
  {32'hc4aa134e, 32'hc336cce8, 32'h434c9c78},
  {32'h4500f11e, 32'h4109ada8, 32'h421df0fa},
  {32'hc4bfe6a9, 32'hc3165ac4, 32'h430fe501},
  {32'h44d52e7d, 32'h42bd65c4, 32'h431dc5a6},
  {32'hc4d55cb4, 32'hc2a8dc02, 32'hc2ba244e},
  {32'h444b9060, 32'hc1ddd6e0, 32'h42c81209},
  {32'hc4c919c8, 32'hc365f50e, 32'h4151b6e3},
  {32'h44ee836a, 32'h4292c6be, 32'hc33cf3ea},
  {32'hc4a6549f, 32'h438e96c6, 32'h433255f1},
  {32'h44ff89c2, 32'h42e54221, 32'h43a9a5d6},
  {32'hc489f9fa, 32'hc18c51ee, 32'h43b784ff},
  {32'h43bb282c, 32'hc4085ed2, 32'hc300b0b9},
  {32'hc4cc60ff, 32'hc23ae3d3, 32'h4307f549},
  {32'h44dc103d, 32'h424da129, 32'hc334b234},
  {32'hc4f13aea, 32'hc30cd433, 32'hc32ec156},
  {32'h43296928, 32'h42a79d9f, 32'h418b5dae},
  {32'hc3c0f9f8, 32'h43aecd87, 32'hc1b7570f},
  {32'h44dc1d5b, 32'hc25d21f4, 32'h4306acdb},
  {32'hc43a30fc, 32'h43394362, 32'h438d1773},
  {32'h445661f7, 32'hc28668a0, 32'h429e1d59},
  {32'hc4787bfe, 32'h40877af0, 32'hc3b7e264},
  {32'h448feb29, 32'hc36e323a, 32'hc33fd91f},
  {32'hc2c759a0, 32'hc37c6dba, 32'hc3eca1e9},
  {32'h4516ef5a, 32'hc3a17277, 32'h42e4db32},
  {32'hc46a3553, 32'h429a595b, 32'hc3b560c0},
  {32'h43fb63ad, 32'h440cea10, 32'hc34ce2b2},
  {32'hc49a682d, 32'h4219d2b4, 32'hc206524a},
  {32'h45010514, 32'hc0f34386, 32'hc364f86d},
  {32'hc446d456, 32'hc1b5515e, 32'h419e3a18},
  {32'h4508379f, 32'hc375eacd, 32'hc345c394},
  {32'hc4e05070, 32'h432eb9fe, 32'h42e213a0},
  {32'h44b17199, 32'hc3041aad, 32'hc3c7d538},
  {32'hc4de3b5c, 32'h43aee7a8, 32'h430f7f6b},
  {32'h449dd82f, 32'hc2c0ef84, 32'h44174154},
  {32'hc505f782, 32'h423b0ded, 32'hc23005e5},
  {32'h450a7b48, 32'hc3a98999, 32'h42d17e9a},
  {32'hc4d058cc, 32'hc2d1ca08, 32'hc3fa065e},
  {32'h43d87fe1, 32'hc34ba698, 32'hc3f23699},
  {32'hc4dd7c90, 32'hc352ca38, 32'h41823537},
  {32'h43cee8a8, 32'h4396dbaa, 32'hc2508046},
  {32'hc45a0254, 32'hc33a7308, 32'h4344fe2f},
  {32'h44f64587, 32'h41f183f3, 32'hc302d782},
  {32'hc4e86210, 32'hc2e1ec10, 32'hc340638c},
  {32'h452715b8, 32'h41d94da1, 32'hc2eda53f},
  {32'hc4e9892c, 32'h4308da9f, 32'hc34b81cf},
  {32'h44c2610d, 32'hc32d1e40, 32'h4377d56d},
  {32'hc4b5f9fd, 32'hc2881fd6, 32'hc2cafd98},
  {32'h440c6692, 32'hc31222ce, 32'hc38ae5d7},
  {32'hc467f19e, 32'h422010a3, 32'h42f9988a},
  {32'h44b2fa44, 32'h43703678, 32'hc3759f1b},
  {32'hc508823a, 32'h4384c849, 32'h42aa9706},
  {32'hc32d4520, 32'h42bfea71, 32'h40f2a22a},
  {32'hc4f5b6ec, 32'hc39ea08b, 32'hc3564e45},
  {32'h44774842, 32'h435a3fc6, 32'hc425468e},
  {32'hc4f8c025, 32'h429cd0c4, 32'hc343781a},
  {32'h45035171, 32'hc3755e3f, 32'h42c1bc42},
  {32'hc4a92bdd, 32'hc1f2bca1, 32'h42d3fa51},
  {32'h4436de4e, 32'hc2619048, 32'h41a56ca1},
  {32'hc4944852, 32'hc33e5441, 32'h441117c2},
  {32'h43f40344, 32'h42889c7c, 32'h4290dc78},
  {32'hc432f6f8, 32'hc3517b18, 32'h428655c6},
  {32'h44be6df5, 32'h42dc1ca5, 32'h42cfe6be},
  {32'hc48a668e, 32'hc25970a5, 32'h43b3e8d6},
  {32'h449fbbff, 32'hc24aa7c5, 32'hc2bf7ff8},
  {32'hc4a1c3cc, 32'hc3fc5deb, 32'hc2505427},
  {32'h450b19f5, 32'h42605315, 32'hc29f5db0},
  {32'hc493fe36, 32'hc3aefb25, 32'h410f29c9},
  {32'h43fbf4cc, 32'h43d80970, 32'hc12f3a3c},
  {32'hc4c92ae6, 32'h4315f4c5, 32'hc336c324},
  {32'h44978815, 32'h4301a1be, 32'h4374cca4},
  {32'hc4840982, 32'hc33bf388, 32'hc20e1fdb},
  {32'h44cd378d, 32'hc3aa7180, 32'h4262026a},
  {32'hc40ab484, 32'hc2900ca6, 32'h41d3a116},
  {32'h42bee4f0, 32'h42fc086a, 32'h4381fb55},
  {32'hc4fcbdea, 32'h42f9ca69, 32'h438a1bf5},
  {32'h44acd7d1, 32'h430adf98, 32'h41fe67cb},
  {32'h4265f940, 32'hc3a1fdad, 32'h4082615c},
  {32'h43025608, 32'h43419f8c, 32'h433f6421},
  {32'hc4e91294, 32'hc3d1e0de, 32'h4316393f},
  {32'h450f433e, 32'h43071c04, 32'h43dd112d},
  {32'hc400c403, 32'h431c194f, 32'h4226e63e},
  {32'h43c299e4, 32'hc2a61fe8, 32'h43f96d7b},
  {32'hc49c2941, 32'h3ff1ed4d, 32'h4438cd09},
  {32'h4402280a, 32'hc35c43d9, 32'h43d667c2},
  {32'hc42b0760, 32'h43d8a8ae, 32'hc324965c},
  {32'h4510f755, 32'h4197ba7c, 32'hc394c549},
  {32'hc38f484a, 32'hc1b8584a, 32'h433251ea},
  {32'h450360e7, 32'h41809967, 32'hc3146926},
  {32'hc50c505e, 32'hc36272fb, 32'h412a351e},
  {32'h4474aedf, 32'h4338e6c2, 32'h436c734a},
  {32'hc3bc5904, 32'h41035026, 32'hc27d6dc7},
  {32'h44af2a05, 32'hc360a74b, 32'h42c96504},
  {32'hc4656c26, 32'h43b9fbfb, 32'hc30a0ce8},
  {32'h44bdaae6, 32'h430c3482, 32'hc214d673},
  {32'hc49428a2, 32'h42f1e7b9, 32'hc3a20f5d},
  {32'h44743250, 32'hc384bfd4, 32'h436cddcc},
  {32'h43710cc0, 32'h43d34d89, 32'h43cc3c1c},
  {32'h448f6fd2, 32'h433531d8, 32'h42516d54},
  {32'hc476d541, 32'h429d9247, 32'hc1fda2c5},
  {32'h4515f574, 32'hc2482bd6, 32'h43ca773f},
  {32'hc4d9ab03, 32'hc13ef6ef, 32'h43fe180c},
  {32'h44906176, 32'hc25041c5, 32'h43a93bd8},
  {32'hc3dd7a00, 32'h42f1aeac, 32'hc3344db1},
  {32'hc358ff70, 32'h41362236, 32'h439bfdf4},
  {32'hc4279a0b, 32'hc3229a1f, 32'hc318698b},
  {32'h44c6977c, 32'h43114c61, 32'hc3916e38},
  {32'hc4b11993, 32'hc2f5c9cf, 32'hc3ad3e63},
  {32'h4447fa2a, 32'hc234e86e, 32'hc2cd7bea},
  {32'hc41e1483, 32'h42f58040, 32'h439c5a29},
  {32'h44cdb2ea, 32'h42794d70, 32'hc3910405},
  {32'hc48e9dc5, 32'hc38bf1cb, 32'hc3b6a287},
  {32'h4504a187, 32'hc3232e46, 32'h42fd846f},
  {32'h42bd85a0, 32'hc3baafc3, 32'h42a3eb23},
  {32'h44f0c052, 32'h42d7cec2, 32'h42bd796f},
  {32'hc41b4ab8, 32'hc31a08ca, 32'hc3cbdaf0},
  {32'h4490ee68, 32'hc208eb73, 32'hc2c75d3d},
  {32'hc41a3c82, 32'h41be210b, 32'h440f7e0b},
  {32'h448fef81, 32'h42bacc26, 32'hc2eb2cad},
  {32'hc4ce0f24, 32'hc330cb07, 32'hc29de732},
  {32'h44fff22c, 32'hc2b17ffb, 32'h43cabc2a},
  {32'hc4ce15ba, 32'hc28b7390, 32'h433c9f05},
  {32'h448fac4d, 32'h41c9bab2, 32'h439bf604},
  {32'hc48dba0c, 32'hc2743974, 32'h42da526d},
  {32'h45186896, 32'h433356e7, 32'hc269703f},
  {32'hc2da8950, 32'hc3a0f2a6, 32'h427af5da},
  {32'h43c4021f, 32'hc293cfab, 32'hc3dae17e},
  {32'hc361f962, 32'hc3e65527, 32'h4311c5d1},
  {32'h45047c44, 32'h4300d9fc, 32'hc38d3101},
  {32'hc3624190, 32'hc3d84f95, 32'hc39f7b0e},
  {32'h44dca6bb, 32'hc3716939, 32'h430e7355},
  {32'hc50849de, 32'h430aa4a7, 32'hc3887122},
  {32'h422bc2a0, 32'hc3d5ddaa, 32'h43226545},
  {32'hc4d5d064, 32'hc3d17476, 32'hc395f9b9},
  {32'h4511ec9a, 32'h43ac82c1, 32'hc3254aa6},
  {32'hc3e18660, 32'h4362bbf9, 32'h42eac18a},
  {32'h450da1f6, 32'h42fa4a16, 32'h42be7cfd},
  {32'hc4daade2, 32'hc3a14e71, 32'hc3124069},
  {32'h44e785e0, 32'hc1e867f9, 32'hc2157f83},
  {32'hc42bd0b4, 32'hc3758de8, 32'h437aa30d},
  {32'h44992776, 32'h4301d2de, 32'hc2bca175},
  {32'hc5133344, 32'hc3c73513, 32'h42c7931e},
  {32'h451080a6, 32'hc36c7bf8, 32'hc195cd77},
  {32'hc4edd4e5, 32'h4082963c, 32'h424826c0},
  {32'h44f53091, 32'hc3016e97, 32'h43057f4f},
  {32'hc2337522, 32'h43022138, 32'h4364dd80},
  {32'h430a5be0, 32'hc290be45, 32'h42dd25d8},
  {32'hc50475d1, 32'h427ab1ae, 32'hc3b87d46},
  {32'h44522eb9, 32'hc308e5de, 32'h42985b9b},
  {32'hc4836f46, 32'hc386caa1, 32'h4277c9f7},
  {32'h441677ba, 32'hc2a7e22a, 32'hc33eabfb},
  {32'hc4da6ec6, 32'hc2a9c5f1, 32'h42e08524},
  {32'h44dfca6e, 32'hc2df9e81, 32'hc28b1cca},
  {32'hc4c459b7, 32'h41e8cc3b, 32'h417d9454},
  {32'h44b313ff, 32'h439d7c5e, 32'h4380e20f},
  {32'hc4a01122, 32'hc2eb71e5, 32'hc2cd9a74},
  {32'h44b1357d, 32'h43935a02, 32'hc41c737d},
  {32'hc5151944, 32'h4381411f, 32'hc2f1d16a},
  {32'h451ee242, 32'h409c6435, 32'hc36553ac},
  {32'hc4dcdfe0, 32'hc2370cf3, 32'h42d4614d},
  {32'h42d51ab0, 32'hc3ed9976, 32'h43bc7ce5},
  {32'hc50c8893, 32'h42b0d3b6, 32'h42c7d6e1},
  {32'hc26d3c28, 32'h436dc3bb, 32'h42dc4ba0},
  {32'hc502ab69, 32'hc1940757, 32'h42c40ecc},
  {32'h439ab334, 32'h41a29803, 32'hc31754e0},
  {32'hc51c3c40, 32'h42685589, 32'h437f22b7},
  {32'h4211b5c0, 32'h42b678bc, 32'hc311a76d},
  {32'hc410a918, 32'hc34cfdd8, 32'hc279cce4},
  {32'h43472318, 32'h43b2eaef, 32'hc2809d0b},
  {32'hc4b48c4a, 32'hc1de4053, 32'hc150a242},
  {32'h44c23bd8, 32'h43a8ebec, 32'hc0f3c028},
  {32'hc4e88b57, 32'h42c514d6, 32'hc2c7edba},
  {32'h4417e14c, 32'hc2c9919a, 32'hc33a8c87},
  {32'hc429cc46, 32'hc39e3ba8, 32'hc25bd786},
  {32'h426d487c, 32'hc2415e1b, 32'h431c6c3a},
  {32'hc4c5f2f8, 32'h433cd235, 32'hc40b5c75},
  {32'h44d73a10, 32'h42a144ce, 32'hc35d1266},
  {32'hc3f446d8, 32'hc24fb108, 32'hc3349773},
  {32'h442fa4b3, 32'hc38bbfcc, 32'h40d7cfc9},
  {32'hc3895b08, 32'h43932849, 32'h435622fc},
  {32'h44be69f9, 32'h3e8240b3, 32'hc32581c5},
  {32'hc5018616, 32'hc3bf72ad, 32'h43138cbb},
  {32'h450b327a, 32'hc320a958, 32'h430bdeb9},
  {32'hc4f4a0e1, 32'hc39e37f8, 32'hc378b249},
  {32'h43ae7244, 32'hc385e046, 32'hc2ed2f08},
  {32'hc325232b, 32'h417c7900, 32'hc374702c},
  {32'h442ed160, 32'h42ed00f5, 32'hc24d7200},
  {32'hc4cf2815, 32'h43039c73, 32'hc42bbf88},
  {32'h44f28a16, 32'h4237de37, 32'hc27298f3},
  {32'hc4f5ed9e, 32'h433b0f8d, 32'hc3152ad8},
  {32'h44abed98, 32'h43073b72, 32'h42f74e6b},
  {32'hc4b64a75, 32'hc2e4566b, 32'hc34e6e50},
  {32'h44c5aaa2, 32'h43186cd3, 32'h4320943f},
  {32'hc4c4ba9e, 32'hc30bb1ac, 32'hc36c437d},
  {32'h451af86d, 32'h41be2056, 32'h42be9e1d},
  {32'hc4a5829f, 32'hc31ad54a, 32'h433e29c1},
  {32'h44c4e7a4, 32'hc21b04fc, 32'h43ecc8dc},
  {32'hc3e286c4, 32'h41895c79, 32'hc309ea44},
  {32'h445690a1, 32'h427d80f6, 32'h41b79a43},
  {32'h42ccfec0, 32'hc3b09893, 32'hc348494f},
  {32'h43adf390, 32'h43695bd4, 32'h43a5964f},
  {32'hc5031b1b, 32'h433a2cbf, 32'h42efe3a8},
  {32'h43649bc9, 32'h415a8d0d, 32'h43c762ea},
  {32'hc48ee1c6, 32'hc365d0d3, 32'h429637e0},
  {32'h4425304c, 32'hc2657edc, 32'hc33b9fc3},
  {32'hc3fe5624, 32'h4149b089, 32'h439b836a},
  {32'h44d4d706, 32'hc2e1ef3c, 32'h42dcd6d0},
  {32'hc4d04728, 32'hc3107d2b, 32'h439b07d3},
  {32'h442a4216, 32'h43927bd2, 32'h423b7479},
  {32'hc4016a5b, 32'hc39a73ff, 32'h42380c52},
  {32'h44dccf57, 32'hc369654f, 32'h431e8ee5},
  {32'hc4656155, 32'hc3b6a5b4, 32'h42ef2a3b},
  {32'h4466801c, 32'hc186fb1a, 32'h438e2e43},
  {32'hc51a808f, 32'h43704b9b, 32'hc2ddb432},
  {32'h44875b33, 32'hc1603409, 32'h43c377db},
  {32'hc43909d2, 32'hc3322b60, 32'hc3d116d2},
  {32'h445089a2, 32'hc2696f6e, 32'h432c9e78},
  {32'hc4e1263d, 32'hc3b89372, 32'hc3427888},
  {32'h43390c88, 32'hc22133df, 32'h418bbce1},
  {32'hc4dd4353, 32'hc345e4ad, 32'hc28b8047},
  {32'h427f17d0, 32'hc307e6f2, 32'h4373a226},
  {32'hc3f6c6e4, 32'hc3977acd, 32'hbf1aa868},
  {32'h43ddb7bf, 32'h420edf8b, 32'h4303d708},
  {32'hc4fd79a8, 32'h42ef2e18, 32'hc2b84b72},
  {32'hc3aee200, 32'h4250c1b9, 32'hc390ac1b},
  {32'h44940ce6, 32'h436fe941, 32'hc28baf67},
  {32'hc47fd094, 32'h443243d2, 32'hc10a4f62},
  {32'h40c08b00, 32'h43313ab0, 32'h438c905f},
  {32'hc402b027, 32'h434712e3, 32'h4291ac02},
  {32'h44f82a2f, 32'hc3d6dbbc, 32'h434f50a7},
  {32'hc3d3c2ea, 32'hc3c3f530, 32'hc421b2ca},
  {32'h421040b0, 32'hc302daef, 32'h4343f1c6},
  {32'hc5150c28, 32'hc33b47cd, 32'hc299b19d},
  {32'h43ceb950, 32'h42b72822, 32'h429d8fb0},
  {32'hc21ef920, 32'h43ab3a77, 32'h423a95f2},
  {32'h4506d54f, 32'h42b319d3, 32'h423993d8},
  {32'h42259e80, 32'h437e1af4, 32'hc33428d3},
  {32'hc2c50080, 32'h4331cf90, 32'h438b23fb},
  {32'hc47f6614, 32'h4328f40e, 32'h432ff8f4},
  {32'h449b8c5c, 32'h41c9fe54, 32'h43aa7555},
  {32'hc4463310, 32'h424a382d, 32'h4164709f},
  {32'h448c893a, 32'h43314f26, 32'h43a89c61},
  {32'hc36d172c, 32'h41a20337, 32'hc2b253fa},
  {32'h44ebcbfc, 32'h43c189e2, 32'h43455bab},
  {32'hc4a629e4, 32'h4315d5df, 32'hc3907803},
  {32'h44c2c18c, 32'h43b34cb8, 32'h42c26c16},
  {32'hc4d69a42, 32'h4365ad85, 32'hc2672c6e},
  {32'h450fd21b, 32'hc37898f7, 32'hbf62c770},
  {32'hc4d0e0a3, 32'h42a7ed0c, 32'hc2c2057e},
  {32'h44ea1a9e, 32'hc3b887ff, 32'h43808073},
  {32'hc3f9f6e0, 32'h438109f8, 32'hc1d6f239},
  {32'h44c9de3a, 32'hc37d72bd, 32'hc2fd030c},
  {32'hc40b91e4, 32'hc3aa639d, 32'hc29b8c5e},
  {32'h44a8ad6e, 32'h4154542c, 32'hc2cfd2f2},
  {32'hc50b7213, 32'hc31a6825, 32'h4298395b},
  {32'h4505bdc1, 32'hc3132d87, 32'hc3ba9729},
  {32'hc32649c8, 32'h41064600, 32'h41ca5f6b},
  {32'h44fe59ae, 32'h43f6f8dc, 32'hc2ec4fda},
  {32'hc32f55d8, 32'hc3aca87b, 32'hc3e54b51},
  {32'h4422b2d7, 32'hc2ff4157, 32'h43d04c47},
  {32'hc4f068d9, 32'hc2bdb005, 32'hc38297e0},
  {32'h44039f3c, 32'h43595fd8, 32'h41fa2096},
  {32'hc5065fb2, 32'hc31d7d38, 32'h42dd33b2},
  {32'h43bc84c0, 32'h4389c8fe, 32'hc31acf14},
  {32'hc4cb8b47, 32'hc307b16f, 32'hc32507f0},
  {32'h443a0bcc, 32'h4235c0a0, 32'hc22cc8aa},
  {32'hc4fddd78, 32'h43883860, 32'hc3773bde},
  {32'h45170002, 32'h436ac730, 32'h438f96a2},
  {32'hc3fb2deb, 32'hc335ac9d, 32'hc341e66a},
  {32'h44b4c577, 32'hc242245a, 32'hc32e819b},
  {32'hc5132fb8, 32'hc3168e6e, 32'h4338c787},
  {32'h44b03fad, 32'h436c5aa8, 32'hc3c15868},
  {32'hc4f1decd, 32'h429b62c1, 32'h4322cd0e},
  {32'h44ae8c65, 32'hc35b9159, 32'hc1b88824},
  {32'hc4c37a2d, 32'h419b32d1, 32'hc41c27f0},
  {32'h44307838, 32'hc40759be, 32'h43412310},
  {32'hc4c334dd, 32'hc3a4836c, 32'h43852ac8},
  {32'h448b5348, 32'h4395fe89, 32'h43a65398},
  {32'hc47cfeb0, 32'h42d150b1, 32'hc30478cb},
  {32'h43d0f93d, 32'hc03dd279, 32'hc3de1478},
  {32'hc392be30, 32'h43937b1f, 32'h432e8493},
  {32'h4497d2c1, 32'hc2ecd807, 32'hc451fe14},
  {32'hc4d65abb, 32'h41ba694c, 32'hc4314dc0},
  {32'h44cc482c, 32'hc320246a, 32'hc187dfca},
  {32'hc445e46c, 32'h429f80c0, 32'hc3c37987},
  {32'h44b443f0, 32'h43279419, 32'hc1d96b84},
  {32'hc44caf22, 32'h43ad0f62, 32'hc3d771db},
  {32'h440caf9e, 32'hc2f57cc5, 32'hc368c6e1},
  {32'hc4b3aa25, 32'h4387dc2d, 32'hc19f3010},
  {32'h44862376, 32'hc20e6da0, 32'h425a845f},
  {32'hc3268750, 32'h41dec7de, 32'hc2b96cf8},
  {32'h45118d52, 32'h43a68e58, 32'hc3328c1e},
  {32'hc468f28c, 32'hc3033d6a, 32'h404f2cea},
  {32'h44d199b4, 32'hc24b0479, 32'hc33f64aa},
  {32'hc4f224dc, 32'hc22527c6, 32'h43afe3b0},
  {32'h44eb56b4, 32'hc388458e, 32'h42984658},
  {32'hc4567d38, 32'hc3c0ad3d, 32'hc42ae338},
  {32'h444e4574, 32'hc20bdf77, 32'hc183058f},
  {32'h42ae6ff6, 32'hc386aa10, 32'h435848ca},
  {32'h43a00364, 32'h43724a3b, 32'h429586c8},
  {32'hc26e5a80, 32'hc382f244, 32'hc0d6e2c4},
  {32'hc2bd1828, 32'hc3012933, 32'hc2e90358},
  {32'hc49e58da, 32'hc2940ee6, 32'hc2d7402d},
  {32'h45095501, 32'hc29b7d07, 32'hc321e5a5},
  {32'hc50b1680, 32'h4318e7dd, 32'hc370beda},
  {32'h44e21b70, 32'h4360045a, 32'hc3d8930e},
  {32'hc4eeb021, 32'hc33dc154, 32'h41c73e57},
  {32'h44888659, 32'h421e118d, 32'h42ddc7cd},
  {32'hc4ff67b9, 32'hc3756c7f, 32'hc39862d8},
  {32'h44f10ff7, 32'h4328e17a, 32'hc229ca0c},
  {32'hc42c3442, 32'h43f001ca, 32'hc38ed6f3},
  {32'h42a6a994, 32'hc33f87b1, 32'h436609d5},
  {32'hc21d81ec, 32'h42c109d4, 32'h43611cd0},
  {32'h425fe1a0, 32'hc3ab150c, 32'hc30524c6},
  {32'hc2d5420e, 32'hc3c65dc6, 32'hc329aea1},
  {32'hc349505c, 32'hc348505f, 32'h41a628e9},
  {32'h4244d820, 32'hc367cc0d, 32'hc3384349},
  {32'h4502e378, 32'hc1e24829, 32'h42db8216},
  {32'hc4c042bc, 32'hc37884ac, 32'hc22c5322},
  {32'h447c1983, 32'hc231f40c, 32'hc375cca1},
  {32'hc3fa036c, 32'hc3830d96, 32'h43faa792},
  {32'h44b4afb8, 32'hc2b9d5bb, 32'h40cba26a},
  {32'hc4311f48, 32'hc3037e6c, 32'hc35a14d6},
  {32'h4503a556, 32'hc3ac12a6, 32'h43837fb3},
  {32'hc492cd24, 32'h41d2b049, 32'hc37bd71e},
  {32'h433eb3b0, 32'h4340ecf1, 32'h428145e7},
  {32'hc45b14c3, 32'h410543fe, 32'h43c8d73f},
  {32'h452328a7, 32'hc31bff37, 32'h41b1afcc},
  {32'hc50c5125, 32'hc2821679, 32'hc282fe82},
  {32'h43c92518, 32'h42178af3, 32'h40d92306},
  {32'hc42f1956, 32'h41f6c179, 32'h43c186c4},
  {32'h44cd2c9a, 32'hc21149d8, 32'h4337ea43},
  {32'hc49be0e9, 32'hc3b9395c, 32'h431615a4},
  {32'h44efa106, 32'hc27dc66f, 32'hc2d470a9},
  {32'hc4408a40, 32'h42f9ef93, 32'hc33aae6a},
  {32'h44fc0a56, 32'h43331191, 32'hc329b74b},
  {32'hc4116f6b, 32'h42af3e13, 32'h42835ab3},
  {32'h44b83142, 32'hc3ca1302, 32'h41af1654},
  {32'hc50134d0, 32'h42751063, 32'h44454c77},
  {32'h433a8f60, 32'h44006def, 32'hc10dfacd},
  {32'hc4b4ca78, 32'h4400ee0b, 32'h435af00d},
  {32'h44b72958, 32'hc308c93d, 32'h42e6ef26},
  {32'hc3c5dabc, 32'h43d7bfb4, 32'h4306a037},
  {32'h4483ff0e, 32'h42c351ae, 32'h42afcef4},
  {32'hc400a5d2, 32'h43500c58, 32'h426d3ac8},
  {32'h443bb740, 32'h42923b90, 32'h43524b73},
  {32'hc4ebfb4f, 32'hc2a73dcb, 32'h436f335a},
  {32'h42fe35d8, 32'h421e98dc, 32'hc1729cc2},
  {32'hc42b11fe, 32'h43a3f722, 32'h43054420},
  {32'h44656584, 32'h432c0970, 32'h43063740},
  {32'hc486d81c, 32'h42ab46d7, 32'h426695fe},
  {32'h44e6e4b8, 32'hc39daf7c, 32'h4309cfcc},
  {32'hc4093848, 32'hc169ccb7, 32'h416ffd4d},
  {32'h444f3074, 32'h433304d1, 32'hc2a9f973},
  {32'hc4f0f8d9, 32'hc219f34b, 32'h43d80b4c},
  {32'h44e7cfbc, 32'hc249016e, 32'hc311034c},
  {32'hc44fd38c, 32'h43c11da3, 32'h42b9cb57},
  {32'h4454ea7f, 32'h42f62690, 32'h436874b1},
  {32'hc4d96027, 32'h42ad883e, 32'h441e6619},
  {32'h44a27e16, 32'hc3399c43, 32'hc30e5976},
  {32'hc486c650, 32'h43bde743, 32'h439493a1},
  {32'h442dfe1e, 32'h41331105, 32'h4246d688},
  {32'hc433180c, 32'hc26ef030, 32'h42670c91},
  {32'h44c4014d, 32'h41f16643, 32'h42cebb0f},
  {32'hc506615f, 32'hc30200f6, 32'h43854242},
  {32'h44d61276, 32'hc18365e5, 32'hc342832f},
  {32'hc394fbe4, 32'hc288a2a6, 32'h43c001e7},
  {32'h4390e81c, 32'h429af405, 32'h433ece12},
  {32'hc31dd120, 32'hc3bb1ff1, 32'h4344a2cd},
  {32'h43e17ec0, 32'hc3418eb4, 32'h43361bc3},
  {32'hc4835e6c, 32'h4390662c, 32'h431e53d8},
  {32'h447bf9e4, 32'h440145b7, 32'hc167b236},
  {32'hc4c47891, 32'hc344be76, 32'h43c3438b},
  {32'h4502a3bc, 32'hc3754247, 32'h43d8b0f8},
  {32'hc430c00c, 32'hc38c0496, 32'h43a8106a},
  {32'h450d2abf, 32'hc3c7a078, 32'h42971907},
  {32'hc502bcad, 32'h43cdba25, 32'h434b6c1d},
  {32'h4353f820, 32'hc20504fc, 32'h42e2aa22},
  {32'hc4703b0a, 32'hc3145987, 32'hc32c72d1},
  {32'h448865a2, 32'h4242cc52, 32'h438461f5},
  {32'hc42add93, 32'h42ca59ea, 32'h42575b33},
  {32'h44e12c34, 32'hc2a54c67, 32'h42cb2236},
  {32'hc4ca6415, 32'hc260f117, 32'hc3a82910},
  {32'h44c45301, 32'hc375a93e, 32'hc334c040},
  {32'hc484f6ca, 32'h42e9c738, 32'h43d80a3d},
  {32'h44f2d32e, 32'hc290695e, 32'hc329131d},
  {32'hc45e19de, 32'h41571e28, 32'h43018555},
  {32'h446d5af2, 32'hc3be28d5, 32'hc30bff6c},
  {32'hc434357d, 32'h41a9786b, 32'h4312f0e6},
  {32'h4501b4e2, 32'hc3a4c81a, 32'hc318eda1},
  {32'hc45e77be, 32'h4325f892, 32'h43c80409},
  {32'h4506b19a, 32'h41ab5285, 32'hc33f357e},
  {32'hc3a33628, 32'h438e7a1f, 32'hc30a6226},
  {32'h44af997a, 32'h433498e0, 32'hc15e3049},
  {32'hc4c5c204, 32'hc3279d4e, 32'hc3608fd5},
  {32'hc2160880, 32'h433f4399, 32'h43d5573a},
  {32'hc4ddba06, 32'h4391a121, 32'h4087efcb},
  {32'h43088a60, 32'hc2d97f18, 32'h41f63047},
  {32'hc301e9a0, 32'h3e9808c4, 32'hc2900106},
  {32'h451696a6, 32'h438fce32, 32'h430ed130},
  {32'hc3d095f4, 32'h42f8635f, 32'hc38aa7ad},
  {32'h44933f09, 32'hc37f484b, 32'hc384b23b},
  {32'hc4665c20, 32'h4365ac0e, 32'h432f0a71},
  {32'h443319cf, 32'h4244059a, 32'hc3bf1fcd},
  {32'hc3d065b8, 32'hc3c831b6, 32'h43769832},
  {32'h44e37598, 32'hc356bced, 32'h42a91b89},
  {32'hc4c9174a, 32'h42ccfca7, 32'h44062da0},
  {32'h4395c988, 32'hc3556270, 32'hc23609c3},
  {32'hc4b6e378, 32'h4390d39d, 32'hc2add97c},
  {32'h436b90c0, 32'h432562c1, 32'h42d9c4e6},
  {32'hc4ab4562, 32'hc31316bc, 32'hc3b4d3e5},
  {32'h44a20b02, 32'hc2261a92, 32'hc311053f},
  {32'hc4a92626, 32'hc3837ad4, 32'h42e71405},
  {32'h4401ebb3, 32'h431f1ddd, 32'hc35c9bcc},
  {32'hc51719dc, 32'hc2cc8e95, 32'hc2164181},
  {32'h44a2deee, 32'h41d50a59, 32'hc2b87f67},
  {32'hc4c81028, 32'hc3c1b642, 32'hc1b5c4de},
  {32'h43aa4104, 32'h43a46180, 32'hc24685e7},
  {32'hc4fc03e4, 32'h435a74ec, 32'h41a4209f},
  {32'h44aeeaf2, 32'h41432237, 32'hc319eee2},
  {32'hc319ccac, 32'hc33b86a8, 32'hc31e90b9},
  {32'h45013a60, 32'h42d63f3c, 32'h40a80689},
  {32'hc4475e98, 32'h431b04e2, 32'h422526e2},
  {32'h43a4fdf8, 32'hc24b7763, 32'h4314acea},
  {32'hc5107313, 32'hc3037792, 32'h43d29aa8},
  {32'h44c35c54, 32'h42b0210a, 32'h43b04305},
  {32'hc32301b5, 32'hc3702141, 32'h436cd88b},
  {32'h44bcc7b1, 32'h42ea03aa, 32'h43284c75},
  {32'hc2b8fa70, 32'hc27007fc, 32'h4383983b},
  {32'h4508ad8b, 32'h434ef6e1, 32'h42a85133},
  {32'hc4822e3a, 32'hc3a722a4, 32'h43233f87},
  {32'h45039fc1, 32'hc3d9572f, 32'h43faf40f},
  {32'h429c5faf, 32'h42abf219, 32'h42fcf13f},
  {32'h44ecd992, 32'hc2fbc6b0, 32'h424c85bb},
  {32'hc4dd44c1, 32'hc21a89db, 32'hc33ddc29},
  {32'h4419f8f5, 32'h431dae30, 32'h4320e91e},
  {32'hc4e3c6df, 32'h42cdae47, 32'h42d143d8},
  {32'h4501b5be, 32'hc23fd657, 32'hc31fb38c},
  {32'hc30c1d18, 32'hc38d23a8, 32'h4233eafc},
  {32'h44103ea8, 32'h434872aa, 32'hc183ce32},
  {32'hc4c56186, 32'hc370b2ce, 32'hc3c68a82},
  {32'h447c9b98, 32'hc35e59f0, 32'h43d8d503},
  {32'hc45810aa, 32'h4209a9d2, 32'hc31e8f5f},
  {32'h43b1864c, 32'h43e73eac, 32'h43872d8c},
  {32'h43882277, 32'h437fc5b9, 32'hc2e25cfa},
  {32'h440d4cf8, 32'hc2d8c5ff, 32'hc31c25b8},
  {32'hc3a86133, 32'hc3675ade, 32'hc3104a42},
  {32'h44590eb4, 32'h42b9b32d, 32'hc35005f1},
  {32'hc50ef45c, 32'h43a097eb, 32'hc2a6db49},
  {32'h450bfd22, 32'h432fe4cf, 32'hc32a02d0},
  {32'hc4a4dc57, 32'h439d16b9, 32'h43114eb8},
  {32'h44f83147, 32'h434cdf95, 32'h42738a6b},
  {32'hc50a79e9, 32'hc1e882b9, 32'h42c2a02d},
  {32'h43bdbefc, 32'hc308dd9d, 32'hc3421705},
  {32'hc4e717ce, 32'h43ae742d, 32'h43495bc1},
  {32'h445e9734, 32'h4190594d, 32'hc36037b4},
  {32'hc35cc0e2, 32'hc2520158, 32'hc2b2fd1e},
  {32'h4472724c, 32'hc316ea68, 32'hc3243478},
  {32'hc4914921, 32'h433d1b8d, 32'h4193ccd2},
  {32'hc37ac65c, 32'h433cee2f, 32'hc3075d8e},
  {32'hc3e81610, 32'h42cf6ae7, 32'h437de91a},
  {32'h4306bfa0, 32'h430b348a, 32'h42a93241},
  {32'hc0fd56e0, 32'hc355fe5d, 32'hc298553f},
  {32'h42d5bcf0, 32'h41a93131, 32'h433575e6},
  {32'hc5116d42, 32'h42a53898, 32'h424e8d83},
  {32'h44cdc91a, 32'hc4104a7f, 32'hc3f31d2d},
  {32'hc514483a, 32'hc3e1ae1e, 32'h43cbf877},
  {32'h41d464f0, 32'h42bc0d06, 32'hc33693bd},
  {32'hc506d2b9, 32'h43e35e0a, 32'h41cc9a0f},
  {32'h44c763e4, 32'h43b79e6c, 32'h43645e37},
  {32'hc37032b8, 32'h42ba496b, 32'hc39b81fa},
  {32'h449a39d6, 32'hc2b2227c, 32'h437acf54},
  {32'hc4586c7e, 32'h42ca6661, 32'h4301c333},
  {32'h449587e8, 32'h4381e5e3, 32'hc18ef96e},
  {32'hc4f510a8, 32'hc3b5727a, 32'hc3505ed3},
  {32'h43f58608, 32'h430403d7, 32'hc28e3da1},
  {32'h42827460, 32'hc3dc2a5a, 32'h4311ad7f},
  {32'h4336d6b0, 32'hc38b81e0, 32'hc323255e},
  {32'hc401d11b, 32'h420f7ac3, 32'h43309173},
  {32'h44fb97e2, 32'h432c43df, 32'hc2eb0a1d},
  {32'hc4ca414e, 32'h432cdbd7, 32'hc3c701e3},
  {32'h438dbd74, 32'h43423210, 32'h420ff06e},
  {32'hc3a8c4ad, 32'h4404bc20, 32'h427c2d4a},
  {32'h4467fcc4, 32'h43085324, 32'hc2d25b87},
  {32'hc43eb408, 32'h4364b819, 32'h4382c25e},
  {32'h448c391d, 32'h43001459, 32'hc38344ee},
  {32'hc49c5efd, 32'h438d51df, 32'hc29b5ee9},
  {32'h4479d7b0, 32'hc3d8755b, 32'h431bb87f},
  {32'hc4500e3e, 32'hc351d5ca, 32'hc3b4269e},
  {32'h45134ee6, 32'hc3618038, 32'h43b8b1dd},
  {32'hc47a141a, 32'h421e8327, 32'hc2de2a51},
  {32'h44b710cd, 32'hc2c3c6b5, 32'hc3b5f366},
  {32'hc33f5b97, 32'h41525121, 32'hc3019147},
  {32'h44b0054a, 32'hc316fc76, 32'h4388f392},
  {32'hc45cde1c, 32'h43386e57, 32'hc2129b11},
  {32'h44d19ff0, 32'hc3071b3d, 32'h4190cfb7},
  {32'hc3c3e6a0, 32'h434ab9a6, 32'hc36bbb7a},
  {32'h44847062, 32'h42ca56e0, 32'h43a35f6a},
  {32'hc396ca63, 32'hc3849031, 32'hc34813ba},
  {32'h44811e85, 32'hc33bfaee, 32'hc2afe2a8},
  {32'hc273e330, 32'h42f90a10, 32'hc3312175},
  {32'h448aebb9, 32'h420ce847, 32'h42a35793},
  {32'hc4f290b4, 32'hc3804f13, 32'hc30a73e7},
  {32'h43aa941c, 32'h42fc0fe9, 32'h423ebaab},
  {32'hc3d7daf0, 32'h4425663f, 32'h43035f5c},
  {32'h440a8aeb, 32'h432f275f, 32'hc39de626},
  {32'hc4f094c9, 32'h438cde62, 32'h431c0728},
  {32'h442130b6, 32'h435f552c, 32'hc1b511fc},
  {32'hc4ebb321, 32'hc358c9d5, 32'h42138abe},
  {32'h448d308c, 32'hc244d20e, 32'h43afefdd},
  {32'hc50aede4, 32'h433148a0, 32'hc2f20eca},
  {32'h44330784, 32'h42cc2b3d, 32'hc2825e07},
  {32'hc463e3a0, 32'h42b7ccdb, 32'hc1cce693},
  {32'h45047e76, 32'hc254885a, 32'h430be8e6},
  {32'hc4b4d577, 32'hc1e5dbd5, 32'hc3a0b6eb},
  {32'h450d95e3, 32'hc2aeb599, 32'h438557cb},
  {32'hc4f0eae8, 32'h42816923, 32'h438f09e8},
  {32'h444d856e, 32'hc2f1f1b7, 32'h41ff1730},
  {32'hc4411b9c, 32'hc1a2cc16, 32'h43acdaa1},
  {32'h4482f7d6, 32'h4385ee7a, 32'h42aa2ce0},
  {32'hc4878ee0, 32'h4389b1ab, 32'hc35cc7ae},
  {32'h44eb8b43, 32'h4151e5c1, 32'h430bae44},
  {32'hc450f484, 32'hc336b246, 32'h42ddfdfc},
  {32'h44a33467, 32'h429b3d20, 32'h437f8176},
  {32'hc5019d33, 32'h4311302f, 32'hc2b83931},
  {32'h4501e70c, 32'h43e2c07d, 32'h42780c3b},
  {32'hc4bdb263, 32'hc3bd920f, 32'h43ad78e8},
  {32'h4520888f, 32'h4274de21, 32'hc25ad40f},
  {32'hc504859c, 32'hc3dfa596, 32'hc22746b6},
  {32'h44a29e08, 32'h4404f9a8, 32'hc2224d5b},
  {32'hc515d570, 32'hc2b886ef, 32'hc3a2c1fc},
  {32'h4493e145, 32'hc365f6ed, 32'hc3bcbaee},
  {32'hc3b27aa8, 32'h42db81f0, 32'hc2976747},
  {32'h446f5090, 32'hc3192b55, 32'h42c8851c},
  {32'hc410e50a, 32'hc2bbfd47, 32'hc355ccae},
  {32'h45360b04, 32'h43e6efd8, 32'h42be3672},
  {32'hc41f04c2, 32'h42cf055f, 32'h42173fea},
  {32'h450b40de, 32'hc29735e6, 32'h424cff26},
  {32'hc503c3bd, 32'h42250838, 32'h424e721a},
  {32'h44eb4aa6, 32'h42df3b79, 32'h43969f54},
  {32'hc500a655, 32'h43059bbe, 32'hc2e440bc},
  {32'h45021e40, 32'hc2b969ba, 32'h418ea150},
  {32'hc43514be, 32'h429710e8, 32'h4297be52},
  {32'h44a71a73, 32'h429cd87c, 32'h43badc13},
  {32'hc4c699fe, 32'h43a421b2, 32'hbf9113f0},
  {32'h44ce8995, 32'hc2cd54e1, 32'h424fafe0},
  {32'h42d4f070, 32'hc19b8b6c, 32'h41370a2e},
  {32'h44e21778, 32'h435a88b8, 32'h43be0894},
  {32'hc4ac0840, 32'hc386da62, 32'hc38d9af6},
  {32'h44d94159, 32'h43c89257, 32'hc2fb2bc6},
  {32'hc49acb47, 32'hc3c35108, 32'hc3a3b135},
  {32'h4491f5f4, 32'h435fac13, 32'hc252bc5a},
  {32'hc32025a6, 32'h4385b8d6, 32'h42beaa4b},
  {32'h450ffd15, 32'hc39de572, 32'h4338f4f6},
  {32'hc4a98617, 32'hc39e21d2, 32'h418f6f54},
  {32'h4302beb8, 32'hc1ea99fa, 32'h4345e52e},
  {32'hc451ec14, 32'hc3bcc6be, 32'hc31f10b0},
  {32'h44cf03f2, 32'h4316b636, 32'hc3989d04},
  {32'hc503c4dc, 32'hc24338c5, 32'h4121bbb0},
  {32'h44f90f16, 32'h426f1976, 32'hc2cde6f9},
  {32'hc4ec1a7c, 32'h438f3c1c, 32'h43a1a679},
  {32'h4505a877, 32'hc2a23a3b, 32'hc31477bd},
  {32'h43ad3e86, 32'hc35c8fef, 32'h42819b8f},
  {32'h447c2b9e, 32'hc3ce32d6, 32'hc3156a61},
  {32'hc464d62b, 32'h42b6d364, 32'hc358c847},
  {32'h44064b00, 32'hc233ee96, 32'hc3913315},
  {32'hc393ffe0, 32'hc3928463, 32'hc3a7cff5},
  {32'h44b0d100, 32'hc3953203, 32'hc2a30307},
  {32'hc49b85c2, 32'hc3105864, 32'h436dd581},
  {32'h42ad639c, 32'h4320cdbc, 32'h418d152c},
  {32'hc44ebe4e, 32'hc2abd1d8, 32'h43c12d4b},
  {32'h44f374a1, 32'h4395d9d6, 32'h4285fee9},
  {32'hc427bd59, 32'h42be2e99, 32'hc387c9dd},
  {32'h44df02c2, 32'hc2af6868, 32'hc377c931},
  {32'hc3fae392, 32'hc1a2cc44, 32'h43243a08},
  {32'h45086b7a, 32'hc2b87cda, 32'h4353775a},
  {32'hc47df4ec, 32'h42446e2e, 32'h42956221},
  {32'h447e0b1e, 32'h4404c628, 32'h43439bc4},
  {32'hc4864768, 32'h4382644f, 32'hc38a8392},
  {32'h4464507c, 32'hc26020f0, 32'hc36064c5},
  {32'hc3e62830, 32'hc30f951d, 32'h41bacb43},
  {32'h4519a434, 32'h4340884f, 32'hc320d4c8},
  {32'hc4e08405, 32'h4330de6a, 32'h43603d8c},
  {32'h441d33e8, 32'h435ee3ff, 32'h42bed0fa},
  {32'hc4c75fdf, 32'hc405ab83, 32'h440db84d},
  {32'h4430816b, 32'hc3c0de4a, 32'h42572eb2},
  {32'hc4c80e8c, 32'hc409a006, 32'h43715cb7},
  {32'h442e2684, 32'h43194eb0, 32'h438b1ffa},
  {32'hc48d6806, 32'h43869ccf, 32'h436234cc},
  {32'h3fe38f00, 32'h43ae1d3f, 32'h41a64914},
  {32'hc5090728, 32'hc37ba646, 32'h431b2e94},
  {32'h44b9d629, 32'hc2e2ea44, 32'hc048f154},
  {32'hc4460392, 32'h43b3487c, 32'h4328ae76},
  {32'h450a7011, 32'h43522a4b, 32'h42bfcabe},
  {32'hc5050591, 32'hc2cc4f08, 32'h43cc270c},
  {32'h45344847, 32'h43cb0fb2, 32'hc337d2b8},
  {32'hc514c502, 32'hc38bf608, 32'h3dba8b40},
  {32'h447d5368, 32'h43b94e85, 32'hc3457489},
  {32'hc4c3e2d7, 32'h41370c74, 32'hc3b7fb6c},
  {32'h4499014c, 32'hc3618713, 32'hc2f92954},
  {32'hc4943d30, 32'hc314e0fe, 32'hc3400ddb},
  {32'h44c6e74d, 32'h42c067c8, 32'hc2415aa3},
  {32'hc4fbb7da, 32'h430be44f, 32'hc33d1232},
  {32'h4508d777, 32'h42eedc73, 32'h42b46ceb},
  {32'hc3f0d210, 32'hc35d15a1, 32'hc3d0404e},
  {32'h45135332, 32'hc2e162f6, 32'hc36d4fe0},
  {32'hc43be076, 32'hc3addbb2, 32'hc286705d},
  {32'h4516d23a, 32'h42aebb85, 32'hc2b86088},
  {32'h429f7454, 32'h436d0312, 32'h43753c1c},
  {32'h4474c9f4, 32'h437ddc0e, 32'h43372632},
  {32'hc4abc98b, 32'hc3d16d5a, 32'hc329b81d},
  {32'h45004fdc, 32'h438a9588, 32'hc275cf06},
  {32'hc30d4280, 32'hc379d15c, 32'hc34d3e2c},
  {32'h4485322a, 32'h42db803c, 32'h430fa291},
  {32'hc3c66bec, 32'h4396ae04, 32'h43d00821},
  {32'h4514cc29, 32'h42b1fafd, 32'hc3801c50},
  {32'hc501f91f, 32'h43697b5c, 32'h42eede3d},
  {32'h44bacad6, 32'h435331cc, 32'h4363b447},
  {32'hc34dbfa0, 32'h435f6266, 32'hc34c7caa},
  {32'h44ae6b58, 32'hc34d1038, 32'hc307f4a7},
  {32'hc4d1f383, 32'h433b63e6, 32'hc3ce979a},
  {32'h44a15b06, 32'hc38cf0c1, 32'hc35df638},
  {32'hc3b45110, 32'hc2cb4f08, 32'hc2336d56},
  {32'h440c6611, 32'h42aba45f, 32'hc311732c},
  {32'hc4b0680a, 32'hc38abdad, 32'hc1cca25c},
  {32'h42a1544c, 32'h42386d74, 32'hc2de05a8},
  {32'hc4ff4a4b, 32'h42478f64, 32'hc310d648},
  {32'h44f94939, 32'hc2150de4, 32'h400c5578},
  {32'hc519107e, 32'hc21f7ad6, 32'h421eb9e8},
  {32'h43c9097a, 32'h413cfbf4, 32'hc3ad72a7},
  {32'hc3ccdd72, 32'h436b25c1, 32'h4188766d},
  {32'h451159d5, 32'h4243f14d, 32'h4260f39c},
  {32'hc4ac578c, 32'h43a6b5dd, 32'h43966b81},
  {32'h437c8e00, 32'hc328bb34, 32'hc3427d36},
  {32'hc3ecb9be, 32'h40d299f5, 32'h436efc14},
  {32'h448ba9f8, 32'hc326a273, 32'h4267724f},
  {32'hc4b0c441, 32'hc40391c3, 32'hc4157da5},
  {32'h448dc223, 32'h43e0f43b, 32'hc28830df},
  {32'hc4c92f22, 32'hc2ebce85, 32'h42b9f270},
  {32'h44e5237d, 32'h429b1cec, 32'h42857d73},
  {32'hc405f822, 32'h43495091, 32'h43b7924b},
  {32'h44f18468, 32'h42fd982d, 32'h43af2303},
  {32'hc19b8c00, 32'hc32886a3, 32'h42c973a7},
  {32'h43bb2df2, 32'h439c88fb, 32'hc33084c0},
  {32'hc4a5b2ce, 32'h43729f71, 32'h4308d633},
  {32'h4474895c, 32'hc36b0dce, 32'hc3bb3130},
  {32'hc39883e5, 32'hc2474957, 32'hc200ed96},
  {32'h4500e710, 32'h4300308e, 32'h432bc3c5},
  {32'hc515bfb7, 32'hc1ebc9e6, 32'h434720be},
  {32'h44f20a24, 32'h4383678f, 32'hc378b52b},
  {32'hc3d4d2ca, 32'hc274ab14, 32'hc2a66148},
  {32'h43febb3a, 32'h429ee09a, 32'h42c36f93},
  {32'hc462599a, 32'h4329a30d, 32'h43ca9d04},
  {32'h44ff1a7b, 32'hc207288e, 32'hc390b140},
  {32'hc4fe2313, 32'h4359a006, 32'hc374937b},
  {32'h44c3a1a4, 32'h43e2f3d8, 32'h42b1af2a},
  {32'h45114a81, 32'hc2204b8a, 32'h43fcdee2},
  {32'hc35272b6, 32'hc1e6dfd5, 32'h42d77233},
  {32'h44ad91e1, 32'hc34067ce, 32'hc2d8919f},
  {32'hc40f671c, 32'hc269ecf5, 32'h41053959},
  {32'h44f05c0b, 32'hc363fb99, 32'hc39536f8},
  {32'hc4e1a6b8, 32'h42972e14, 32'h42507032},
  {32'h4428bfaa, 32'hc2bb899a, 32'hc39cbf75},
  {32'h43a96084, 32'hc3d08db8, 32'hc2a73510},
  {32'h447a3792, 32'hc36b7750, 32'hc2367b31},
  {32'hc46bff22, 32'h431fbba3, 32'hc208cd66},
  {32'h44c24c7b, 32'h42ee926c, 32'hc29a7598},
  {32'hc4e59ce1, 32'hc24e8012, 32'h42bdff6f},
  {32'h447ef834, 32'h43547809, 32'h42b30a13},
  {32'hc50cd910, 32'hc3996f56, 32'hc3821355},
  {32'h44dd8aa1, 32'hc2e016e3, 32'h4397166b},
  {32'hc498830f, 32'hc3e1cbf8, 32'h42c1604e},
  {32'h412e3780, 32'hc328f0ba, 32'hc38b7cee},
  {32'hc3c0b9fe, 32'hc1f674d7, 32'h4384af6a},
  {32'h45004a53, 32'hc3458a91, 32'hc37f635c},
  {32'hc4169a5c, 32'h43438f26, 32'hc2d1fded},
  {32'h4446048a, 32'hc2e47290, 32'hc37e80dc},
  {32'hc4ec5bd0, 32'hc1f1fa5d, 32'h4114c195},
  {32'h44a5323a, 32'hc2e82e01, 32'hc1905f61},
  {32'hc4e7c6a5, 32'h43230075, 32'hc35182e2},
  {32'h4410cb5c, 32'hc20679f7, 32'hc368a976},
  {32'hc484fd77, 32'hc179ea91, 32'hc38af3bf},
  {32'h436badf2, 32'hc37ee895, 32'hc367d47a},
  {32'hc4f8fdf2, 32'hc3a1d883, 32'hc33c327f},
  {32'h449f09c1, 32'hc1e138ec, 32'hc32a2301},
  {32'hc43420ce, 32'hc287bb96, 32'h42d71156},
  {32'h44bf9597, 32'hc36f3b76, 32'h4403379f},
  {32'hc4b1ba3b, 32'hc317ceda, 32'hc2bf5f81},
  {32'h44abdcb3, 32'h42f01304, 32'hc39b6377},
  {32'hc503ce32, 32'h432c7ff9, 32'hc3300267},
  {32'h44b522ef, 32'h42ad64d4, 32'hc29f46f6},
  {32'hc3cc5ec0, 32'hc378f8d4, 32'hc30cebaa},
  {32'h44c41ef5, 32'hc28f2c91, 32'hc2c88189},
  {32'hc4a5c60b, 32'h440fd3b3, 32'h42605a2f},
  {32'h43f82bee, 32'hc3a52413, 32'h43b2faca},
  {32'hc48a641c, 32'h41f3b4f7, 32'h4386773a},
  {32'h43ceb75a, 32'hc385597f, 32'hc23c8037},
  {32'hc4cc2da4, 32'h430ca9fc, 32'hc3c713a2},
  {32'h448c1d20, 32'hc3b7c530, 32'h43817c85},
  {32'hc4cd1b67, 32'h4381c0fc, 32'h43b859ae},
  {32'h44dc1422, 32'hc1a7c60c, 32'h42c9daf4},
  {32'hc4eb9837, 32'hc3978b38, 32'hc2dcbe59},
  {32'h450ebc31, 32'h432e7955, 32'h43ca5366},
  {32'hc50eb8c8, 32'h42df8774, 32'hc2984e7b},
  {32'h4463280e, 32'h441cb225, 32'h42d7f159},
  {32'hc35ecb22, 32'hc31eea20, 32'h42a822d3},
  {32'h4462a03e, 32'h4280563b, 32'hc3514a63},
  {32'hc3efd774, 32'h422e994d, 32'h44002ec8},
  {32'h450e6533, 32'h444d4c21, 32'hc30b0c5d},
  {32'hc247d958, 32'hc344af55, 32'h42cdf371},
  {32'h44aa5f82, 32'hc30465b1, 32'h43b88e4c},
  {32'hc4c4a546, 32'hc31c8921, 32'hc2e94146},
  {32'h42e8f479, 32'hc20010b7, 32'h432b476d},
  {32'hc4993588, 32'hc3684302, 32'hc32ab15c},
  {32'h4519c6e3, 32'hc3abde72, 32'hc29bfa4f},
  {32'hc4c0dd45, 32'h43156b1b, 32'hc0d4508c},
  {32'h44ed9642, 32'hc3acd5f0, 32'h43a1a914},
  {32'hc43b4de2, 32'h43c7e662, 32'h43580e0d},
  {32'h4351357a, 32'h429f055e, 32'hc36b79bb},
  {32'hc5103f11, 32'h41c936ed, 32'h4398ed50},
  {32'h44ec43a6, 32'hc3199595, 32'h43221ead},
  {32'hc4f8e859, 32'hc29c9ac5, 32'h42848d19},
  {32'h4477c0f8, 32'h436aace5, 32'hc4056b79},
  {32'hc4e4997d, 32'h42e90ed3, 32'hc2e1b2f5},
  {32'h443e32b8, 32'hc382beac, 32'h4328893f},
  {32'h41c10bd6, 32'hc2c0808d, 32'h440d1499},
  {32'h451b4f77, 32'hc310c150, 32'h43342706},
  {32'hc516570b, 32'hc21dac34, 32'hc25016b6},
  {32'h4483223f, 32'h42761d9a, 32'h4425fb7b},
  {32'hc43ce6d8, 32'hc3442ec9, 32'hc3c0c1c3},
  {32'h44d0a24e, 32'hc1e3b5e9, 32'h439653e4},
  {32'hc4a7d8f8, 32'h427d1e9a, 32'hc34043c7},
  {32'h45009c11, 32'hc3fc1c20, 32'h4260c48d},
  {32'hc438a865, 32'h4409c59f, 32'hc3c9aade},
  {32'h4504ac0b, 32'hc287c8ab, 32'h44026a82},
  {32'hc4f74916, 32'hc3879fce, 32'h43359cc2},
  {32'h43d9a598, 32'hc30e63d4, 32'hc398e619},
  {32'hc4a4a9a9, 32'h428598b9, 32'h438b3451},
  {32'h44575466, 32'h423bd23f, 32'hc2bc3e77},
  {32'hc4bd8259, 32'h42cea46b, 32'hc2ea6b96},
  {32'h45056385, 32'h4285969e, 32'hc0d25010},
  {32'hc506c373, 32'h4384b49e, 32'h40bebc4a},
  {32'h44c710f5, 32'h42a7d6f7, 32'h430e8e78},
  {32'hc4c109cd, 32'hc32a9c28, 32'h42895890},
  {32'h44d3d515, 32'h42e7acf6, 32'h43674437},
  {32'hc4fd0acd, 32'hc3a4027c, 32'hc38c48d3},
  {32'h449cc106, 32'hc2d14ed7, 32'hc421164d},
  {32'hc4202fc6, 32'h42abea25, 32'h42a39d51},
  {32'h44df0639, 32'h430c3186, 32'h441bc7ee},
  {32'hc4abd582, 32'hc1a29d0b, 32'hc3839991},
  {32'h43d1e4cc, 32'h43046b45, 32'h42c367e9},
  {32'hc4ea79d0, 32'h4331f23c, 32'h43ee2bbe},
  {32'h449a0e1d, 32'h43a3bd86, 32'h423e7522},
  {32'hc487112d, 32'h4367ba7e, 32'hc3a47a16},
  {32'h43bc18a0, 32'hc3663284, 32'h42d36243},
  {32'hc41ce438, 32'h435423e0, 32'h436f2772},
  {32'h447e91cb, 32'h4253addd, 32'h43044031},
  {32'hc3109750, 32'h43f792a5, 32'hc0bc3d98},
  {32'h446a8be2, 32'hc3a29197, 32'h43974257},
  {32'hc420b274, 32'hc3bb48e2, 32'hc3765ad2},
  {32'h43da0ec6, 32'hc3a61205, 32'h431d7499},
  {32'hc4da291b, 32'hc18885be, 32'hc341edc1},
  {32'h43bb11af, 32'hc29a2344, 32'hc36b6614},
  {32'hc4bffd6f, 32'h44216711, 32'h42bbd111},
  {32'h4506fe28, 32'h3fedfd08, 32'hc2425666},
  {32'hc4cc341f, 32'hc2f91b3c, 32'hc38b3489},
  {32'h4445d01b, 32'h42becb43, 32'h42a1f166},
  {32'hc457035f, 32'hc393bbe5, 32'h42a54afc},
  {32'h44ebbdbf, 32'h435be6e2, 32'hc260f8fd},
  {32'hc3d6ce77, 32'h43925335, 32'h42f40f5b},
  {32'h44035299, 32'hc2ef4f81, 32'hc138daac},
  {32'hc4f7c11c, 32'h434b81e4, 32'hc1dcbc1f},
  {32'h44e99208, 32'h439613b3, 32'hc257eacc},
  {32'hc4956201, 32'hc34b5ae7, 32'hc405db59},
  {32'h44cbd05f, 32'h440f155c, 32'h423ab55c},
  {32'hc4cbcad0, 32'hc3d121f0, 32'hc29308ba},
  {32'h44330458, 32'h42d2e733, 32'hc3099010},
  {32'hc46df110, 32'h43b88f94, 32'h4396a9b7},
  {32'h43fbb220, 32'h43642eb9, 32'hc33ff4dd},
  {32'hc393d45b, 32'h437f7f1d, 32'hc26d996b},
  {32'h44c582d0, 32'h43952da4, 32'hc3041ec4},
  {32'hc438c144, 32'hc383282f, 32'h4210e4d8},
  {32'h45064bbe, 32'h42d8054e, 32'hc31cce4a},
  {32'hc4aad7ef, 32'h437d3220, 32'h43cb9fa0},
  {32'h44b482d4, 32'hc3c54d53, 32'hc332fd18},
  {32'hc503b81b, 32'hc36d31c5, 32'h439f645f},
  {32'h446d40d6, 32'h42a973f4, 32'h43a044b0},
  {32'h431bbd60, 32'hc2f9cc68, 32'hc1b94e9e},
  {32'h44e61f4c, 32'h41965c44, 32'hc287d449},
  {32'hc46ddb8c, 32'h4343a4b2, 32'h43081695},
  {32'h4520c6fa, 32'h43a19fef, 32'h4344f638},
  {32'hc3a966e0, 32'h42a8089c, 32'hc355b95f},
  {32'h451313e2, 32'h436f4698, 32'hc307024e},
  {32'hc4f4fc52, 32'h43773a62, 32'h43a3d787},
  {32'h44441ab1, 32'h4186b2bd, 32'hc2da65c3},
  {32'hc39d2750, 32'h42402632, 32'h43643b81},
  {32'h44392e34, 32'hc30610cd, 32'h42a319f3},
  {32'hc4847f1f, 32'h4339beed, 32'h438d137f},
  {32'h439c48f6, 32'hc3cf7207, 32'h43053351},
  {32'hc4abcd8c, 32'hc239590c, 32'hc1f92d5f},
  {32'h446cedc8, 32'hc245931f, 32'hc15a197a},
  {32'hc4bb5560, 32'hc2a9a30e, 32'hc33e2051},
  {32'h44a88938, 32'h43dd930e, 32'h43347382},
  {32'hc4c1d99e, 32'h41cc7fce, 32'h4339c2e1},
  {32'h448d5b58, 32'hc38a2d28, 32'hc292262f},
  {32'hc50221e8, 32'h439a94dd, 32'h436e5d89},
  {32'h44fd3a87, 32'hc32aa640, 32'h41bc70a5},
  {32'hc4dc7eed, 32'hc381862f, 32'hc3313f22},
  {32'h43ea9b44, 32'hc2a54118, 32'hc36a7708},
  {32'hc50c6976, 32'hc3d35f50, 32'hc27c034c},
  {32'h44e8dfa0, 32'h4353464c, 32'h42886914},
  {32'hc4c72195, 32'h424bc9be, 32'hc2deadd5},
  {32'h44e95fdf, 32'h4184eca1, 32'h4213dc4a},
  {32'hc50e9c00, 32'h4393a9d8, 32'h403137d0},
  {32'h44d5317c, 32'hc34e36f9, 32'hc316843e},
  {32'hc4a1db93, 32'h43aa7d77, 32'h43204b83},
  {32'h44ba0083, 32'h41f927d5, 32'hc383381a},
  {32'hc419cdb5, 32'h42afa345, 32'h435c3180},
  {32'h44126a42, 32'h43cdae36, 32'h42da554c},
  {32'hc4156f6a, 32'h435cbe01, 32'h43916a74},
  {32'h45073e87, 32'h42c5f2e1, 32'h436e6187},
  {32'hc3b5f6c0, 32'h418e3e04, 32'hc387dda0},
  {32'h4385467c, 32'hc34525a0, 32'h42c52f0d},
  {32'hc4bec1c7, 32'hc347a7f5, 32'hc1a56172},
  {32'h44b58916, 32'hc2e92471, 32'h4311e494},
  {32'hc3d77776, 32'h432e809c, 32'h429b8fce},
  {32'h44b9c58f, 32'hc3767e86, 32'h431bdf14},
  {32'hc41f992f, 32'h430be2ae, 32'h421414a5},
  {32'h4469d0d3, 32'h42c8cc54, 32'hc3a3a64b},
  {32'hc4c02949, 32'hc3445799, 32'h432654e8},
  {32'h45027e19, 32'h43a7b223, 32'hc238ba87},
  {32'hc3325bfa, 32'h4250f282, 32'h425a5269},
  {32'h44603ec3, 32'hc2643b37, 32'hc2d04803},
  {32'hc486f8d7, 32'hc25be227, 32'hc2884f6b},
  {32'h4497a345, 32'hc0916397, 32'hc3661267},
  {32'hc3c8dc3c, 32'h432383e0, 32'h42dedc3a},
  {32'h43c2226c, 32'hc2c6306e, 32'hc3c9eb1f},
  {32'hc3e47484, 32'h4363a5e2, 32'hc383b478},
  {32'h44c442d3, 32'hc3c29239, 32'h42047fd7},
  {32'hc5007933, 32'hc38cdf7f, 32'hc34ac2d5},
  {32'h442922b0, 32'h43aca49d, 32'h431f2e42},
  {32'hc2cd4292, 32'h42d9b1e7, 32'h429d68ec},
  {32'h44acc0d2, 32'hc29e160f, 32'hc34228d2},
  {32'hc4c399f5, 32'h44031bde, 32'hc371c44f},
  {32'h45001d3e, 32'h43fa6d17, 32'hc348a3c3},
  {32'hc255fd20, 32'h41af3dd5, 32'h42c86c2c},
  {32'h450bf05f, 32'h42b0ff27, 32'h4247027c},
  {32'hc3a2394a, 32'h423237a3, 32'hc1fe01d9},
  {32'h44b5f81b, 32'hc3690bfc, 32'hc2b429f9},
  {32'hc4631fd8, 32'h43127406, 32'h4125f788},
  {32'h43c6f93c, 32'h42d24f11, 32'h425be65e},
  {32'h42912d00, 32'hc1623948, 32'hc2228f7c},
  {32'h447ef597, 32'hc34e1c99, 32'hc3297dc0},
  {32'hc4833909, 32'hc3550b8c, 32'h43643d27},
  {32'h4506fcb9, 32'h420e8026, 32'h43ab51da},
  {32'hc42052d2, 32'hc3ae0e32, 32'h44024b58},
  {32'h445dea73, 32'h435275a5, 32'h442406c3},
  {32'hc3289db0, 32'hc36d9a98, 32'h42abac6f},
  {32'h446562f0, 32'hc31aba11, 32'hc31d734f},
  {32'hc44598d7, 32'hc2c098b4, 32'h440396fd},
  {32'h443e6ff8, 32'hc401bee1, 32'h44045765},
  {32'hc40adc5a, 32'h40cd8018, 32'h4346c07d},
  {32'h44ae6512, 32'hc3d1f832, 32'h430d42d7},
  {32'hc4f6d562, 32'hc1071620, 32'hc4355195},
  {32'h433d6230, 32'hc3161e00, 32'hc37059a6},
  {32'hc47670fc, 32'hc2e6d22f, 32'hc3132744},
  {32'h450fdbc2, 32'hc3953eee, 32'hc398a160},
  {32'hc5044ee1, 32'h43949c59, 32'h42d856b9},
  {32'h44fbe2ec, 32'h429166a5, 32'h438a34a3},
  {32'hc48a7522, 32'h42ce62b8, 32'h42ecf041},
  {32'h44efaf1e, 32'h429a2df8, 32'hc3015814},
  {32'hc4bb00f2, 32'hc32f57d2, 32'hc335ab25},
  {32'h438caa08, 32'hc3692d61, 32'h431790cd},
  {32'hc4baa0f7, 32'h430cda85, 32'hc2872e9a},
  {32'hc13aad00, 32'hc35b91ba, 32'h42fb31be},
  {32'hc4d5d024, 32'h437b3160, 32'hc31aebee},
  {32'h434a2f28, 32'hc1ef2bf4, 32'h42098b73},
  {32'hc48b47e2, 32'h43d2f4f2, 32'h43b995e9},
  {32'h43a78ddf, 32'hc2b5557c, 32'hc3da5232},
  {32'hc4c76c0c, 32'hc26d4667, 32'h43ce5a40},
  {32'h448b8d67, 32'hc3c2cbd5, 32'hc3282836},
  {32'hc498a4df, 32'hc328daed, 32'h436283a9},
  {32'h43c86bcc, 32'h4399f917, 32'h440f3349},
  {32'hc3f8b3c0, 32'hc37f4688, 32'hc2848c94},
  {32'h4432e1a9, 32'hc27f44b1, 32'h43acb7b9},
  {32'hc1aa43c0, 32'hc0ee3d0b, 32'hc19c76aa},
  {32'h44f8b1ca, 32'h4405b830, 32'hc30bf45e},
  {32'hc50a6f19, 32'hc2991508, 32'h414519a7},
  {32'h44b8c9d1, 32'h418ff56b, 32'h4288a54a},
  {32'hc4a9a42d, 32'hc319b363, 32'hc3163af0},
  {32'h44b9db17, 32'hc3608604, 32'hc2a391a7},
  {32'hc515f649, 32'hc4163d7c, 32'hc2aa56f9},
  {32'h44e31bd6, 32'hc3051c9b, 32'hc2c25147},
  {32'hc4ce43be, 32'hc378150c, 32'hc0f17135},
  {32'h44b4f137, 32'hbef04560, 32'h43682d42},
  {32'hc4a74384, 32'hc2879435, 32'hc3e52527},
  {32'h44c5cc43, 32'hc2c55bb1, 32'hc351de84},
  {32'hc4e258aa, 32'h42bfbf08, 32'h41185d8e},
  {32'h445c5d72, 32'hc31669aa, 32'hc32e5296},
  {32'hc4f8bbf3, 32'h431357ac, 32'hc200fc16},
  {32'hc29508b8, 32'h43015bf0, 32'h437ad3ca},
  {32'hc50e0638, 32'h4312014d, 32'h41e657f6},
  {32'h44a71fca, 32'hc3a1900c, 32'hc376c9a2},
  {32'hc4ba2337, 32'hc40ed6d6, 32'h414e894c},
  {32'h44fc2b80, 32'h41bf4ad9, 32'h435cb350},
  {32'hc4b78b0b, 32'hc37cf11a, 32'hc398b52a},
  {32'h43499140, 32'h434d11b6, 32'h41e085ca},
  {32'hc4ca02be, 32'h43145f68, 32'hc281530d},
  {32'h44a93de8, 32'hc380ccd9, 32'h431eda74},
  {32'hc500aea9, 32'h4386ccdd, 32'hc2a15dba},
  {32'h44c3af32, 32'hc340e8fb, 32'hc3ae8bf8},
  {32'hc4fcbab2, 32'hc3a44c34, 32'hc3e850c2},
  {32'h44c4b6b4, 32'hc2c3761d, 32'hc2359fba},
  {32'hc48ba4ed, 32'h4385ed8c, 32'hc3c2a8d8},
  {32'h451ecbec, 32'hc2ed1fc8, 32'hc381893f},
  {32'hc4fe8556, 32'hc2b2ce76, 32'hc304d47a},
  {32'h4519f34a, 32'h43bb6797, 32'hc3eb3f58},
  {32'hc2e53e53, 32'h43c5ceab, 32'h43020d50},
  {32'h44b3e159, 32'hc1a6ce7d, 32'h42f8f230},
  {32'hc41cec15, 32'hc383a77c, 32'h4294f2d6},
  {32'h43dfee78, 32'hc337120b, 32'hc36b66e0},
  {32'hc424a2ff, 32'h42ac929f, 32'h42d38d4b},
  {32'hc2fb2148, 32'h433f6591, 32'hc2a27945},
  {32'hc4e3532d, 32'hc30834d9, 32'h42be608a},
  {32'h44705c14, 32'h43fdbccb, 32'hc29bda66},
  {32'hc3a97ee5, 32'hc39aa253, 32'h429a5a63},
  {32'h44a1ccd3, 32'h4390b034, 32'h425e8293},
  {32'hc4ee9f0e, 32'h42b721fa, 32'h43131f47},
  {32'h44b96b1d, 32'hc3d7ab6f, 32'h4234858f},
  {32'hc4b1cb40, 32'h42d02bb6, 32'hc2df1285},
  {32'h44dac86f, 32'h42dc856f, 32'hc3284abd},
  {32'hc4a6f0fa, 32'hc329cb99, 32'hc330a273},
  {32'h4485f36b, 32'h4282289c, 32'hc16a71e0},
  {32'hc4d8af1c, 32'h4368f4de, 32'h4301a4d3},
  {32'h450b0502, 32'h42348618, 32'h4388eca6},
  {32'hc4aae225, 32'hc219bcc0, 32'h42931860},
  {32'h4420d152, 32'h43ed2ace, 32'h43a2204b},
  {32'hc43cc958, 32'h43864a17, 32'hc2f64b3f},
  {32'h45076451, 32'h41b135ec, 32'h42c26556},
  {32'hc4936be3, 32'hbea02498, 32'hc2425e47},
  {32'h450430ba, 32'h4393ffea, 32'hc29eda96},
  {32'hc43c0474, 32'h43835b28, 32'hc32e4510},
  {32'h4478615b, 32'hc30ea210, 32'hc3937b61},
  {32'hc4cd0f8f, 32'hc38ca122, 32'h432f6233},
  {32'h44e3f0db, 32'h43b2de12, 32'h41e0ef2e},
  {32'hc4090c12, 32'h4298fffe, 32'hc3af1b2d},
  {32'h4418e020, 32'hc35db512, 32'hc3371c28},
  {32'hc4b5cd89, 32'h438fe9c8, 32'hc2a6bbeb},
  {32'h4515e7fc, 32'hc38e72ac, 32'h43ce00a0},
  {32'hc4ded819, 32'h4245df95, 32'h42849e09},
  {32'h4416d6b8, 32'hc39d05be, 32'h4286ae97},
  {32'hc504e3ef, 32'hc38a40da, 32'h4385a03e},
  {32'h45142d22, 32'hc2a424c1, 32'hc353ada6},
  {32'hc4c4e38c, 32'h4400d893, 32'hc333c70f},
  {32'h44d06231, 32'h4108f9a2, 32'hc2c1a6e0},
  {32'hc3941b72, 32'h436816e2, 32'h4322e3a1},
  {32'h44d86e43, 32'hc29281fe, 32'hc29bdd69},
  {32'hc500c265, 32'hc403119f, 32'h43599a10},
  {32'h43861b92, 32'h40d15741, 32'hc3238c01},
  {32'hc4d9433a, 32'h42d86873, 32'hc2c22b7e},
  {32'h44f20a3f, 32'h43368c69, 32'h43230590},
  {32'hc3930fee, 32'h4320c793, 32'h425df1bb},
  {32'h42f67dc0, 32'h437f9dab, 32'h43067405},
  {32'hc50a43af, 32'hc33fd3ce, 32'h4316a245},
  {32'h45043929, 32'h439330b0, 32'h4258120f},
  {32'hc4c4d2e2, 32'h42999dc9, 32'h42f4bc1e},
  {32'h45059997, 32'h44391a17, 32'h42c53915},
  {32'hc38cef72, 32'h43597bfd, 32'h40701416},
  {32'h44de0c09, 32'h4139ad24, 32'hc2835f5d},
  {32'hc4a1d434, 32'hc3a7a8e7, 32'hc30ed26a},
  {32'h445dc7c8, 32'hc1bf8b91, 32'hc34ad99f},
  {32'hc3f019a0, 32'h428af546, 32'hc34356df},
  {32'h45001688, 32'hc3da46b0, 32'h431e5982},
  {32'hc385a096, 32'hc39cfb64, 32'h42cfbe3f},
  {32'h44182c5a, 32'h438b2a1d, 32'hc2869646},
  {32'hc4e8c8cc, 32'h43459f9e, 32'h4253878e},
  {32'h44e28d9c, 32'h43ce27a2, 32'h4390ef4d},
  {32'hc377d0d0, 32'h43356026, 32'hc36e8a41},
  {32'h44018d88, 32'h42003d47, 32'hc235fc24},
  {32'hc45984b0, 32'hc387ec58, 32'hc36925d8},
  {32'h44a35223, 32'h40a19074, 32'h4344eb2f},
  {32'hc45cf2ae, 32'hc2bbf7d5, 32'hc22e7c28},
  {32'h444323b0, 32'hc393923b, 32'h43138444},
  {32'hc4e6bc38, 32'h42310c54, 32'h41c5fde1},
  {32'h4507fc1c, 32'hc1b57d1b, 32'h43a46704},
  {32'hc4b95c6e, 32'h42cb09e3, 32'hc323cae1},
  {32'h4502279b, 32'h44118bb1, 32'h43c4e957},
  {32'hc486347b, 32'h43035746, 32'h4370d4bf},
  {32'h44060921, 32'h4333b8b9, 32'hc31b4fd8},
  {32'hc4099368, 32'h4391fc28, 32'h422daa51},
  {32'h445a1762, 32'h438e5a90, 32'hc28cae77},
  {32'hc4e9fc6c, 32'hc421489c, 32'hc3a894cf},
  {32'h440f040b, 32'h41e04440, 32'hc29ec742},
  {32'hc4e62ff0, 32'hc397b650, 32'hc20ab703},
  {32'h44dc1f2c, 32'h433cf5dd, 32'hc1e8eb06},
  {32'hc48e1f54, 32'hc2b94324, 32'h44012926},
  {32'h44c2cf2a, 32'h436fbeb6, 32'h4363fb7d},
  {32'hc44314ac, 32'hc31b2dc9, 32'hc17e3bed},
  {32'h44cce65a, 32'h43ae1a45, 32'hc2b950b7},
  {32'hc4478b8c, 32'hc2474664, 32'hc3557b17},
  {32'h449ab351, 32'hc356037c, 32'hc329c0ef},
  {32'hc38a7c70, 32'hc26b549b, 32'hc123beea},
  {32'h44a83608, 32'h43765070, 32'hc233758c},
  {32'hc4a77916, 32'h43adea20, 32'hc2c33008},
  {32'h43e37b25, 32'hc33da50c, 32'h437f4285},
  {32'hc3c3a63c, 32'hc27da5dc, 32'hc39f13d6},
  {32'h44b6f200, 32'hc33a3a4e, 32'h42c3eaa4},
  {32'hc414a490, 32'hc3a60c2a, 32'hc26678e0},
  {32'h4519e9c2, 32'h4301b280, 32'hc3a3f28b},
  {32'hc51214d2, 32'hc29975b1, 32'h43022e4a},
  {32'h44a4d2e9, 32'h42abd908, 32'h4362d39c},
  {32'hc354eaa4, 32'h4333297e, 32'h426ebcd0},
  {32'h44bb37ff, 32'hc397f921, 32'h42ef1d56},
  {32'hc47718a1, 32'h43cac752, 32'hc2694b7e},
  {32'h439d110a, 32'hc267e29e, 32'h4393d27e},
  {32'hc5235a62, 32'h430e9844, 32'hc2edfe55},
  {32'h44ed97bf, 32'hc387a217, 32'h429490e5},
  {32'hc35759c0, 32'h439561ee, 32'hc38280e2},
  {32'h436f2fa8, 32'hc36aa192, 32'hc27bed2c},
  {32'hc486a05f, 32'h432d0bf2, 32'h43221028},
  {32'h44f411d1, 32'h431ec2e1, 32'hc26b6e54},
  {32'hc4c64aa8, 32'h43e266e0, 32'hc32449ba},
  {32'h4504f44a, 32'h43781bea, 32'hc3ae36fe},
  {32'hc5213729, 32'h42e5dcb8, 32'h438e3702},
  {32'h44c2b3ba, 32'hc3952386, 32'h43d56067},
  {32'hc4fffcba, 32'hc2395ad4, 32'h431f7208},
  {32'h44d6ff16, 32'h42030053, 32'h440fbfe0},
  {32'hc3819ae8, 32'h408259c8, 32'hc3920731},
  {32'h43e8e708, 32'hc2f73da3, 32'hc251999b},
  {32'hc4bdce8a, 32'h42df1ba4, 32'hc2badaed},
  {32'h43116024, 32'h432e6784, 32'hc3674f9e},
  {32'hc48833b9, 32'h419fd2ee, 32'hc10820ef},
  {32'h44aeebd9, 32'h41afb700, 32'hc1efd677},
  {32'hc5050388, 32'hc285b53c, 32'hc2a93a54},
  {32'hc2b47b30, 32'h43c22ba2, 32'hc2172b92},
  {32'hc3d8977f, 32'h41db172d, 32'hc2a8f63d},
  {32'h451f0e08, 32'h4402fe9d, 32'h4383b2a2},
  {32'hc50cebbc, 32'hc2f59465, 32'h43554506},
  {32'h44e2eff0, 32'hc3c5a9e8, 32'h43dd7dbc},
  {32'hc4938d95, 32'h44209b16, 32'h43bd66b3},
  {32'h451f0ece, 32'hc28ad0bf, 32'h432ae810},
  {32'hc2ab4b40, 32'h439a8646, 32'hc1d297d0},
  {32'h43eac2a8, 32'h42fb145f, 32'hc2d15ae1},
  {32'hc4388449, 32'h418c7521, 32'h41f8eb30},
  {32'h44aa1322, 32'hc2d7f772, 32'h42003928},
  {32'hc4b4dd4d, 32'hc2d5b887, 32'hc35454bc},
  {32'h44e05f2e, 32'h4297b9e5, 32'h42210699},
  {32'h42cb4580, 32'h436b85cc, 32'hc1b413d2},
  {32'h44a44eb9, 32'hc1a593a8, 32'hc155c974},
  {32'hc384bcb8, 32'hc386146a, 32'h419e477c},
  {32'h451cd5f6, 32'hc2e07bde, 32'hc334a50e},
  {32'h41f40800, 32'h43aaa33b, 32'hc339c89a},
  {32'h44953c84, 32'h4232adb3, 32'hc3022ae8},
  {32'hc4dd3c77, 32'hc2c10f29, 32'hc35c1280},
  {32'h441cd884, 32'h41c9d288, 32'hc1f26ae4},
  {32'hc4fc5d15, 32'h43a0aaa5, 32'hc2e67243},
  {32'h4274a440, 32'h41a3baa3, 32'h439f916e},
  {32'hc511aa48, 32'h433a2a9a, 32'hc2cffbcf},
  {32'h45268bdf, 32'h43110873, 32'hc3acd20a},
  {32'hc3c66850, 32'h428a2aa4, 32'hc36c9916},
  {32'h451ebc4a, 32'h432ae5b6, 32'hc28577f9},
  {32'hc418041e, 32'h43ebcd80, 32'hc3b4b26a},
  {32'h443d4640, 32'h4367b70e, 32'hc319095e},
  {32'hc4bed7f5, 32'hc3dacd97, 32'h4121ba5b},
  {32'h44c10c94, 32'h42c06282, 32'h4350c0f7},
  {32'hc4db5db1, 32'h42ab1c46, 32'h43a15a6d},
  {32'h43b4fd28, 32'h4338a0f6, 32'h435fa6de},
  {32'hc39272b8, 32'h43414242, 32'h4319f3e7},
  {32'h44f660c5, 32'h43a75c17, 32'hc3b429bd},
  {32'hc502bc7c, 32'h42ad25d5, 32'hc2b02dd3},
  {32'h44c42f76, 32'h4329cd46, 32'h42c27b64},
  {32'hc48e177a, 32'hc29c93d1, 32'h4277ab62},
  {32'h445fb4d2, 32'h42577cc7, 32'hc120967a},
  {32'hc4abb654, 32'hc3524dfa, 32'hc191458e},
  {32'h448b7987, 32'h42fa5f5d, 32'h42d7abff},
  {32'hc50c5e4b, 32'h43411dce, 32'hc3100ec2},
  {32'h450a3cd9, 32'hc3856a29, 32'hc29c8331},
  {32'hc4be9e4d, 32'h422021f2, 32'hc31eae0a},
  {32'h44f30c6d, 32'h42fa9370, 32'h415761ec},
  {32'h40b3061c, 32'h43a149d2, 32'hc3cba18c},
  {32'h45033b3f, 32'hc1ed1538, 32'hc383ebd0},
  {32'hc38986d0, 32'h430b7933, 32'hc30a1248},
  {32'h44c0c8b0, 32'h42e43f12, 32'h411c2030},
  {32'hc5098c5a, 32'hc2fd5225, 32'h4397451d},
  {32'h44915a30, 32'h42a3d7d7, 32'hc28ff714},
  {32'hc47b8247, 32'hc3529093, 32'hc28682c8},
  {32'h44861be6, 32'hc22a30a1, 32'hc3d3291c},
  {32'hc462a5f2, 32'h4330f524, 32'h431921a7},
  {32'hc4038478, 32'hc2a0db9d, 32'hc2288435},
  {32'h449f7d1c, 32'hc3366fd4, 32'h43a998a6},
  {32'hc46c59bb, 32'h43bfcf59, 32'h434d8bdb},
  {32'h44da3404, 32'h42fd0032, 32'h4318e1ac},
  {32'hc281dd94, 32'hc3c19373, 32'h42faedf8},
  {32'h44540ad0, 32'hc30a0734, 32'h4307ade5},
  {32'hc4ff0bf9, 32'hc377705b, 32'h42d783bd},
  {32'h45051ebf, 32'h437adac4, 32'h410adf2b},
  {32'hc4d7d409, 32'h425c0bb8, 32'hc2f5f863},
  {32'h4453a858, 32'h424140e6, 32'hc3685168},
  {32'hc4b8ed04, 32'hc32923d4, 32'hc34ac473},
  {32'hc06a5c00, 32'hc33eb25e, 32'h43896f8f},
  {32'hc4c2b53a, 32'h4321a3bf, 32'h4294c534},
  {32'h4411c51f, 32'h42b4b37d, 32'h4344b4e1},
  {32'hc43f68a6, 32'hc3c6dae5, 32'h437f41cd},
  {32'h4432bdd2, 32'h4280eb8d, 32'h4386c253},
  {32'hc4a7711a, 32'hc0c2bbaa, 32'hc32f59eb},
  {32'h4493006f, 32'h424c64f3, 32'hc3674620},
  {32'hc4115efe, 32'h439b7757, 32'hc35c2ca2},
  {32'h441cfa31, 32'h433d2a47, 32'h4314cb23},
  {32'h4329087e, 32'h432a61e2, 32'hc2b6f729},
  {32'h43bfc49e, 32'hc23fb050, 32'hc12595ef},
  {32'hc4509892, 32'hc30536e4, 32'hc383719b},
  {32'h4484efdc, 32'hc3805093, 32'h42dd4473},
  {32'hc4ccbb15, 32'h43b1dd1d, 32'hc25874b3},
  {32'h44e67391, 32'hc0e4befb, 32'hc32fdf60},
  {32'hc49a8731, 32'hc123ed32, 32'h43497ff4},
  {32'h4510adb5, 32'hc3e50ff5, 32'hc36fa5bd},
  {32'h43f5aaf3, 32'h4406ce49, 32'h42819a99},
  {32'h445cbf42, 32'h4378bbaf, 32'h42b26b00},
  {32'hc43974e7, 32'h4359974a, 32'hc0ad5ca5},
  {32'h43c717b1, 32'hc321e5c0, 32'h432d798b},
  {32'h432886c2, 32'h431830cb, 32'h429b803c},
  {32'h44a53986, 32'hc364f912, 32'h438b746e},
  {32'hc4697e1f, 32'h4407b074, 32'h41afea14},
  {32'h4501c59d, 32'h425c420a, 32'h42b1ae5d},
  {32'hc3924680, 32'hc3232e86, 32'hc31cff96},
  {32'h44851d34, 32'h4400b676, 32'h4307e914},
  {32'hc480c6fd, 32'h43acbdb0, 32'h4285a5ad},
  {32'h452676ca, 32'h419c77a0, 32'h43bd218e},
  {32'hc4871d4e, 32'h4286b88a, 32'h43ab6d71},
  {32'h4502bae3, 32'h43b34d5c, 32'h43a681a4},
  {32'hc49a338e, 32'hc3e8b5c2, 32'hc3028c6a},
  {32'h4518f12d, 32'h433706c8, 32'h436ce0ef},
  {32'hc458a4d4, 32'hc35eef65, 32'hc34dafe8},
  {32'h44eb870a, 32'h430b280c, 32'h438ba44d},
  {32'hc35dafec, 32'hc2ba9d45, 32'h423f64c1},
  {32'h45008cea, 32'h43099590, 32'hc3b19fbb},
  {32'hc507d7d4, 32'hc1438aa5, 32'hc0bee038},
  {32'h44e8db3a, 32'hc27f84bd, 32'hc41d520f},
  {32'hc4b572da, 32'hc2420fe4, 32'hc389ded5},
  {32'h42e20cca, 32'h44071557, 32'hc280d868},
  {32'hc4241f28, 32'hc2283435, 32'hc38fc713},
  {32'h44ab7a31, 32'h427dac21, 32'hc3a1d559},
  {32'hc49ae7b7, 32'hc1df2577, 32'hc42b74dd},
  {32'h4436181e, 32'h420edb7f, 32'hc373654f},
  {32'hc4ea891b, 32'h439553da, 32'h4211350f},
  {32'h4467ea24, 32'hc3344b58, 32'hc287b9ff},
  {32'hc4977dd8, 32'hc3597e7c, 32'hc3275444},
  {32'h45034af3, 32'hc2c5ad60, 32'hc24c9d41},
  {32'hc3b5f220, 32'h4369bb08, 32'h43584fda},
  {32'h45083bce, 32'h41eec0c0, 32'h42f2b069},
  {32'hc493bce6, 32'hc2cd1a8e, 32'hc3bbf407},
  {32'h44330dd2, 32'h3f894266, 32'h43507582},
  {32'hc500c50b, 32'hc2be50df, 32'h438d1409},
  {32'h445f6206, 32'h43cd7ad2, 32'hc11ff681},
  {32'hc340d940, 32'h43846a37, 32'h40dbad90},
  {32'h44f94c17, 32'hc32d33ec, 32'hc3b0ee5e},
  {32'hc4f006fa, 32'h422108e4, 32'hc1cbaad2},
  {32'h43badfe9, 32'h42a89353, 32'hc2d58d62},
  {32'hc426d16e, 32'h43ed79ed, 32'h43021a6a},
  {32'h4371bd82, 32'hc24874de, 32'h434dcace},
  {32'hc49d23cd, 32'hc4291883, 32'h422af1ac},
  {32'h4401feff, 32'h4392f78b, 32'hc0e84872},
  {32'h43b18df8, 32'hc2596f09, 32'h4389c7a0},
  {32'h42fd2420, 32'h424e536f, 32'hc380d6e9},
  {32'hc5067608, 32'hc10096f5, 32'hc39defaa},
  {32'h44c87871, 32'hc2d8dc41, 32'h4328ca31},
  {32'hc409d1b5, 32'h439e83fd, 32'h43930a91},
  {32'h44b23e5d, 32'hc450b96e, 32'h43dcb698},
  {32'hc48dd43a, 32'hc415f669, 32'hc33e66ea},
  {32'h44f09fea, 32'h42beb685, 32'h4205c356},
  {32'hc50f7ff2, 32'h43e948bd, 32'hc10d10a7},
  {32'h43df9210, 32'h43d16d96, 32'hc3e9227e},
  {32'hc2a00840, 32'hc1fcbb98, 32'hc3beaf01},
  {32'h44b84989, 32'hc3037cd9, 32'hc32ce556},
  {32'hc4ee225c, 32'h4214cc4d, 32'h435f2a52},
  {32'h43cfd5d6, 32'h43ae806f, 32'h4324175e},
  {32'hc1f3c020, 32'h43026bcb, 32'hbfb73464},
  {32'h443bfb73, 32'hc36d3798, 32'hc3289020},
  {32'hc3e1d350, 32'hc208bf42, 32'hc33abf16},
  {32'h450cc120, 32'h4231036c, 32'h42744ecf},
  {32'hc3014cc0, 32'h41890352, 32'h4369c3d0},
  {32'h42e33430, 32'h42ef91e5, 32'h434b7177},
  {32'h43fc2098, 32'h43bdc5bf, 32'hc2a5ece4},
  {32'h44308746, 32'hc20b0480, 32'h42a03d2c},
  {32'hc44d0c65, 32'hc3d32436, 32'h4340b34f},
  {32'h44be1199, 32'h3fe87c6c, 32'h431ebb7a},
  {32'hc4cf6fc7, 32'hc2ff5272, 32'h433d0216},
  {32'h44b6f20e, 32'hc3ef3d28, 32'h4235e5be},
  {32'h43208ae8, 32'h43662410, 32'hc3adb898},
  {32'h450ab5cc, 32'h43afbeee, 32'hc27117cb},
  {32'hc4aa64e5, 32'h430c7917, 32'h4103a034},
  {32'h4428bb31, 32'h4364d315, 32'h43fd5e26},
  {32'hc50177bf, 32'h41c7f7c6, 32'h431f99e5},
  {32'h42ac360c, 32'h427635af, 32'hc3314359},
  {32'hc487ae1a, 32'hc2c4cecb, 32'hc3802d6f},
  {32'h4502550b, 32'hc2a7aa38, 32'hc390d5a6},
  {32'hc3ba8520, 32'h436805ec, 32'hc12b3c0e},
  {32'h44774f52, 32'h43b0a60d, 32'hc252978a},
  {32'hc3a4f068, 32'h43fe29e0, 32'hc2ed19e0},
  {32'h452dbae6, 32'h43b26596, 32'hc15443eb},
  {32'hc501b99f, 32'h435a7167, 32'hc3842cce},
  {32'h4447a270, 32'hc2f21b8e, 32'h42801a0c},
  {32'hc36351dd, 32'hbea66bea, 32'hc308a060},
  {32'h44fd4f5c, 32'hc2038096, 32'hc3bddfab},
  {32'hc482c8d8, 32'h41f7cf6f, 32'h43867fa7},
  {32'h43723e40, 32'h4383dce3, 32'hc2947d4c},
  {32'hc49a997c, 32'h4390e0b0, 32'h436a45b5},
  {32'h447e7b8e, 32'hc32f19e7, 32'h421a5778},
  {32'h42c07738, 32'h435b6658, 32'h43589163},
  {32'h43cd927e, 32'h4214a40e, 32'hc2604bad},
  {32'hc4eacb8b, 32'h42fd6c89, 32'h43faf74a},
  {32'h44aeab34, 32'h43bb2c46, 32'h431c6011},
  {32'hc497db45, 32'h43731cfb, 32'h4360b81f},
  {32'h43cb1805, 32'hc3c14ab3, 32'h43020845},
  {32'hc4f40525, 32'h4272bb10, 32'h439e7dd0},
  {32'h444fa1b2, 32'hc2c6e20e, 32'hc32d5eea},
  {32'hc4f65e1e, 32'hc32b22c2, 32'h40fc11c8},
  {32'h44645242, 32'h402adb38, 32'hc0c7cd03},
  {32'hc4e66a69, 32'h436f3a60, 32'hc21a483f},
  {32'h44dffb39, 32'hc330e266, 32'h430b112c},
  {32'hc381563c, 32'hc3184c42, 32'hc31ca593},
  {32'h451b7a56, 32'h43255564, 32'h42317fb3},
  {32'hc430c1e8, 32'h4347e206, 32'h439869b0},
  {32'h44e10e09, 32'hc315de04, 32'h43725e9d},
  {32'hc507c743, 32'hc2b03b9a, 32'h4220fffd},
  {32'h442024df, 32'h431dbfc5, 32'h3fd7f88c},
  {32'h4325a1cc, 32'h4355c31e, 32'h42a5fd7f},
  {32'h43db9808, 32'hc3144f39, 32'h4395cab7},
  {32'hc3f51aa7, 32'hc28c1395, 32'h43c2e5ba},
  {32'h44e21a2a, 32'h42499c7e, 32'h416f01a6},
  {32'hc408d449, 32'h434c10bb, 32'h42b7296d},
  {32'h4385994c, 32'hc39625bd, 32'h4287bcb9},
  {32'hc4901c87, 32'h43277f5b, 32'h438a58ed},
  {32'h44e428d4, 32'hc2c28655, 32'h4285ad4a},
  {32'hc5115d41, 32'h43c876ce, 32'h42fe75fe},
  {32'h44ce27ca, 32'h42ab34d4, 32'h417f6cda},
  {32'hc48063a6, 32'hc3a80d4a, 32'hc0113714},
  {32'h44a74af7, 32'hc2ccfeb4, 32'hc37dee18},
  {32'hc4ca9151, 32'h413ce5ce, 32'h42cd6af3},
  {32'h44cd9066, 32'h43a0d280, 32'h43a2913e},
  {32'hc4c6aa14, 32'h43453d2d, 32'hc333d6a8},
  {32'h4453bb20, 32'h426dd853, 32'hc2b6f635},
  {32'hc39ffc18, 32'hc2d75931, 32'h4300ff37},
  {32'h4401ead0, 32'h42580a87, 32'h42a7640a},
  {32'hc4f1a2ff, 32'hc39f42e9, 32'hc237c099},
  {32'h44990f1c, 32'hc33c59dc, 32'hc1d59363},
  {32'hc518b50c, 32'h42a6c94c, 32'hc252e477},
  {32'h449db779, 32'h427c4508, 32'h43b3ce75},
  {32'hc43138c2, 32'h439bf04c, 32'hc2c0ea47},
  {32'h44a2a699, 32'h4239bb7e, 32'hc30f97bf},
  {32'hc4bb778c, 32'h4349a3a5, 32'hc35a079d},
  {32'h438985e8, 32'h4353e20f, 32'hc33ad2b1},
  {32'hc50bf7ec, 32'hc0e60aa4, 32'hc2f25ff5},
  {32'h44cce45c, 32'h42ad0eb6, 32'h41b9adf4},
  {32'hc4cffd48, 32'hc10f3616, 32'h43bfbe7b},
  {32'h4370f620, 32'hc290db24, 32'h438cc8af},
  {32'hc3e7ebc0, 32'h42f6b566, 32'h41a355ae},
  {32'h4221c9a0, 32'hc30c0626, 32'h436a79b5},
  {32'hc39755b8, 32'h43ed1aa5, 32'hc2c07f55},
  {32'h440aa35b, 32'hc3974a63, 32'h42b867b5},
  {32'hc4cb101e, 32'hc38aa41a, 32'h43cae68b},
  {32'h44f0615e, 32'hc3a540fc, 32'h4387227a},
  {32'hc4e3d2ae, 32'h420d0fe9, 32'h419e51fc},
  {32'h4446b6e7, 32'h431d9aec, 32'h440e7dcb},
  {32'hc4949965, 32'hc2416214, 32'hc35bc2b5},
  {32'h44a1c596, 32'h42efd7e9, 32'hc303469a},
  {32'hc4a58722, 32'hc2c93b05, 32'hc33bd4a4},
  {32'h4480f7be, 32'hc3161a2a, 32'h434a96bc},
  {32'hc40c30d8, 32'h4228d738, 32'hc2dd4d58},
  {32'h450e92fc, 32'h4348dd6e, 32'h430fd2f0},
  {32'hc49e543d, 32'h41f11ea5, 32'h4144ce3b},
  {32'h450b48ad, 32'h43d3eb89, 32'h4381c168},
  {32'hc451f338, 32'h4224480a, 32'h42d0ec65},
  {32'h44173e66, 32'hc23a939a, 32'h43891ab4},
  {32'hc3677e76, 32'h432c0b11, 32'h4205ae2d},
  {32'h448fe1fe, 32'h432d637c, 32'hc20bbee8},
  {32'hc44712f8, 32'hc39cb866, 32'h4269209a},
  {32'h44284b54, 32'h43c51cb5, 32'hc2873e5a},
  {32'hc498d008, 32'h42091302, 32'h431ae875},
  {32'h44440e78, 32'hc3d2600b, 32'hc3130464},
  {32'hc3cdf444, 32'h41ac7ee0, 32'hc17db3a8},
  {32'h44ef96a0, 32'hc38fb60d, 32'h428da08d},
  {32'hc432603d, 32'h42ab0c7c, 32'h42ffcd6a},
  {32'h450bb245, 32'hc337f00c, 32'h431e4f55},
  {32'hc1afe0ff, 32'hc33fb276, 32'h42fb8252},
  {32'h43f24bb8, 32'hc209faf6, 32'h435bcea6},
  {32'hc4afed33, 32'h42142708, 32'h420c64f7},
  {32'h435163e8, 32'hc3479307, 32'h42cb2282},
  {32'hc45a76d7, 32'hc311da97, 32'hc3182149},
  {32'h45027a32, 32'h43ea3ee8, 32'h43febd77},
  {32'hc3bb3e69, 32'hc2a39778, 32'hc349c961},
  {32'h44cd1332, 32'h43c795b0, 32'h42aa801a},
  {32'hc3ea0cd4, 32'h42dcda6c, 32'h42403872},
  {32'h44542364, 32'hc34389e3, 32'hc350cc3a},
  {32'hc4a1cb28, 32'hc40544c9, 32'hc2c54455},
  {32'h44f69f75, 32'h438134d0, 32'h4287a317},
  {32'h432bf4e4, 32'h42beea69, 32'hc3320ca6},
  {32'h44bcd66c, 32'h43ea6cc1, 32'hc2e3d7a4},
  {32'hc4e1d8f6, 32'h42c06c4f, 32'h428ab9e4},
  {32'h4523227d, 32'hc3961ebc, 32'hc3b3c4ec},
  {32'hc4e4ae66, 32'h43850e81, 32'h43b14ff4},
  {32'h44353bd0, 32'h437b512c, 32'hc26666ec},
  {32'hc4de4578, 32'h4356d67f, 32'h4312b26f},
  {32'h444f90bf, 32'h430286f2, 32'h423d2115},
  {32'hc5013fe4, 32'h425480f8, 32'hc2ed392f},
  {32'h44bb3e50, 32'h4325f533, 32'h42f39f08},
  {32'hc48bfef8, 32'hc326ee26, 32'h43936211},
  {32'h43c5b9fc, 32'h439c9b42, 32'hc3393f2c},
  {32'hc441fb5c, 32'h43087c8f, 32'h4243e524},
  {32'h448264c3, 32'h41eb2bd5, 32'hc3ae2276},
  {32'hc4eaf686, 32'h43325340, 32'h41d205ce},
  {32'h4509c76e, 32'hc2867d86, 32'hc3330234},
  {32'hc4715c24, 32'h41e30936, 32'h41f3efe0},
  {32'h4501fe28, 32'h42911ed8, 32'h42446ba6},
  {32'hc367d778, 32'h4396ac1b, 32'hc31b5551},
  {32'h43fddf5a, 32'hc057bac2, 32'h4316f59d},
  {32'hc4989222, 32'h42c337a2, 32'h438fb067},
  {32'h449c4423, 32'h4358d38f, 32'hc3227af9},
  {32'hc384fad7, 32'h42d17b75, 32'h42a9edd4},
  {32'h448d4edc, 32'hc34c3918, 32'h42a97f89},
  {32'hc42a058c, 32'h4391aa94, 32'h43e8ecfe},
  {32'hc2c81210, 32'hc3563922, 32'hc27ee287},
  {32'hc4939afe, 32'hc37e5a65, 32'hc3bbc817},
  {32'h44ca79bf, 32'hc327f53f, 32'hc3602f0f},
  {32'hc4a81dd3, 32'hbfbda1c0, 32'h430478af},
  {32'h439d1b38, 32'h433755b0, 32'h4327f33c},
  {32'hc4a2aa05, 32'hc32e2474, 32'h43ccf916},
  {32'h4450bb03, 32'hc2576e75, 32'hc1875d01},
  {32'hc4edb7ea, 32'hc3463f8e, 32'hc3c9be8f},
  {32'h437fd8a8, 32'h435e456c, 32'hc383b147},
  {32'hc39b6a1f, 32'h438b3f2b, 32'h42ddfb8c},
  {32'h44fd334a, 32'hc38c51d8, 32'h4306c601},
  {32'hc468a693, 32'hc16b6872, 32'h43364bf0},
  {32'h449f9442, 32'h43deb623, 32'h4305943c},
  {32'hc4faaf1e, 32'hc2cc675a, 32'h43b367ca},
  {32'h44245710, 32'hc3131c35, 32'hc13edce8},
  {32'hc48e53b9, 32'h43fec5db, 32'h43f01719},
  {32'h44c4f63e, 32'hc31c4669, 32'hc3515119},
  {32'hc4a5607a, 32'h42a7560c, 32'h41ac2405},
  {32'h44afeeff, 32'h43223cb8, 32'hc1c32f96},
  {32'hc448130b, 32'h42c557c5, 32'hc30efd12},
  {32'h44fc29bc, 32'hc2861faf, 32'h43dc46c7},
  {32'hc3331103, 32'hc24243bc, 32'hc31d241e},
  {32'h448c1666, 32'hc2945a21, 32'hc2d198b4},
  {32'hc424986b, 32'hc286894e, 32'hc2bbb1f0},
  {32'h440d59ba, 32'h4316d942, 32'h423fdbec},
  {32'hc4ab37de, 32'hc315aa48, 32'hc3eea582},
  {32'h4500be43, 32'h43a40c07, 32'h43b427e0},
  {32'hc38aee60, 32'h43144df6, 32'hc3a1141b},
  {32'h44b8d1fd, 32'hc39201ad, 32'h4380f312},
  {32'hc4d772db, 32'hc325dade, 32'h43618614},
  {32'h4408d04f, 32'h43a4c0e4, 32'h43cb030f},
  {32'hc424f77c, 32'hc382af3c, 32'h4374f2af},
  {32'h44155b3c, 32'hc3656113, 32'hc30e5654},
  {32'hc4dea81b, 32'hc1bdec33, 32'h430511f4},
  {32'h43f1f2cb, 32'h417260f6, 32'h430a1cdf},
  {32'hc4ee9e90, 32'h431c331c, 32'h41b548ce},
  {32'h45000c68, 32'h4207aa17, 32'hc29478fb},
  {32'hc479c836, 32'h42e7fa32, 32'hc29ab61e},
  {32'h44d468c0, 32'hc25a5188, 32'hc1da282f},
  {32'hc43e84fc, 32'hc38e94c8, 32'h3df43a80},
  {32'h43dccb0e, 32'h420859e4, 32'hc383f1e9},
  {32'hc3eb79b8, 32'h42082d44, 32'hc36cf773},
  {32'h44d6747b, 32'hc3990669, 32'hc40efe9a},
  {32'hc46826bc, 32'hc373a311, 32'hc30645f6},
  {32'h4442fa83, 32'h43898140, 32'h41759ea8},
  {32'hc4b5a0f1, 32'h41d71a58, 32'hc447ff20},
  {32'h4486fc91, 32'hc31f313e, 32'hc28bee4c},
  {32'hc31ae9c0, 32'hc35dd212, 32'hc2e82ed7},
  {32'h44fea278, 32'h42fe940f, 32'hc2fa0a2b},
  {32'hc4e546e0, 32'hbf30a215, 32'h431a63e5},
  {32'h44093b7c, 32'h42d22ebf, 32'hc30f6f4a},
  {32'hc45b55b8, 32'h42b54b78, 32'h43608284},
  {32'h451f1dfa, 32'hc350d979, 32'h436a75d2},
  {32'hc4c06042, 32'hc380c65b, 32'h439551d2},
  {32'h44f7b3de, 32'hc311fc41, 32'h41c8f245},
  {32'hc3bd7b9e, 32'hc0abdacb, 32'hc166cde4},
  {32'h4514538b, 32'hc235f78e, 32'h43c8fbbe},
  {32'hc41d08c1, 32'hc2b1acbb, 32'hc34faa29},
  {32'h442bb744, 32'h42b9c7d0, 32'hc3941996},
  {32'hc4f1c924, 32'h42373376, 32'h41ac9957},
  {32'h451434c8, 32'h438bb6e8, 32'hc220dbcc},
  {32'hc3acad80, 32'h4392f5e3, 32'h428f4f62},
  {32'h451253a4, 32'h439595ea, 32'h4343e412},
  {32'hc397dd14, 32'h424315cd, 32'hc0d49e91},
  {32'h450a2fcc, 32'hc35fbef3, 32'h43f34af1},
  {32'hc4c17a00, 32'hc2f073d0, 32'hc252cf1e},
  {32'h4521ebb3, 32'hc3886178, 32'h432397ed},
  {32'hc41be196, 32'hc167302b, 32'h42e65a94},
  {32'h444b8d07, 32'h42dc1179, 32'hc18d09a2},
  {32'hc464199c, 32'hc18f0bd0, 32'h42add9d3},
  {32'h44be1090, 32'h423fa840, 32'hc3b2640b},
  {32'hc37c77a6, 32'hc322649a, 32'hc1b04b6e},
  {32'h45067afa, 32'h430a6b13, 32'h42e75a31},
  {32'hc4910c1b, 32'h4392c21e, 32'hc42725aa},
  {32'h448e9306, 32'hc3f3ca4b, 32'h42f4525f},
  {32'hc4988622, 32'hc385bb1c, 32'h43bc84ce},
  {32'h450f01ce, 32'h42339127, 32'h437b949a},
  {32'h42fb999e, 32'h4327afb9, 32'h406643de},
  {32'h451e325f, 32'hc30edee7, 32'hc38025e5},
  {32'hc49b6e0c, 32'h41e4773b, 32'h43cc8656},
  {32'h44b8ae7f, 32'h4349f740, 32'h4350a2eb},
  {32'h40ee7a00, 32'h43a9d400, 32'hc33c3c38},
  {32'hc30e0e3e, 32'hc30b053e, 32'hc409a13e},
  {32'hc4c9bbd3, 32'hc2d32324, 32'hc3b53ce9},
  {32'h44074881, 32'h4283d926, 32'h432cfad2},
  {32'hc4c5ceff, 32'h43e29003, 32'hc3f1dfaf},
  {32'h4321a381, 32'hc33ef7c2, 32'h420a43b2},
  {32'hc47da69a, 32'hc40474cf, 32'h42d04def},
  {32'h42fa0980, 32'h434d41fb, 32'hc355bafe},
  {32'hc489f60c, 32'h43430c56, 32'hc3bbb24e},
  {32'h44d26bc0, 32'hc1768cf8, 32'h405618ca},
  {32'hc5141808, 32'hc2fef6a7, 32'hc28ecdd4},
  {32'h44d6da76, 32'hc25914e8, 32'h42e2952b},
  {32'hc4d695ca, 32'hc3928ab9, 32'hc3b098c9},
  {32'h449fbd28, 32'h438bc644, 32'hc20d76b0},
  {32'hc51096c5, 32'h43cf0481, 32'h4391583c},
  {32'h450d80fc, 32'h42346fdb, 32'hc1fe8a4d},
  {32'hc3c700b8, 32'hc3246b28, 32'hc31aa40a},
  {32'h44aed93a, 32'hc1755a32, 32'hc387b6c6},
  {32'hc50ea4d2, 32'h433f420c, 32'hc22cff07},
  {32'h45139dec, 32'hc2c9f83d, 32'hc3ce4835},
  {32'hc4776d44, 32'hc3e17475, 32'hc3c9c4ab},
  {32'h44ae178c, 32'hc1a67152, 32'hc29f9508},
  {32'hc3802e53, 32'h42fc9d8c, 32'hc316c12f},
  {32'h44ed287c, 32'hc35dc7c8, 32'hc385b5cf},
  {32'hc4a9e537, 32'h43f262a7, 32'hc3a8f443},
  {32'h42a50340, 32'h42cadfcc, 32'hc30262e6},
  {32'hc3b12d0e, 32'h4379e1e6, 32'hc3c5c782},
  {32'h4505f829, 32'hc25199f2, 32'h42992fb2},
  {32'hc49ad47c, 32'h4211f0e1, 32'h4345f945},
  {32'h4431225e, 32'h43a10c7e, 32'hc2be904f},
  {32'hc507dc86, 32'hc3677c1e, 32'h4349ccee},
  {32'h44e66f94, 32'h420609cb, 32'hc352dccd},
  {32'h436fbf90, 32'h42cf1946, 32'hc28ac39a},
  {32'h441306e5, 32'h4343f862, 32'h40cb75fa},
  {32'hc4121a5c, 32'h41752b8a, 32'hc2b2eb08},
  {32'h4498a8a7, 32'hc35d63ae, 32'hc198f1c0},
  {32'hc2de0384, 32'h431d767c, 32'hc2fefda2},
  {32'h44a91b6b, 32'h432a20d1, 32'hc3a07e63},
  {32'hc4ee99fc, 32'h43d04ed5, 32'h43612d0b},
  {32'h44e00391, 32'hc3f62079, 32'h43d72425},
  {32'hc477c35c, 32'h432ea166, 32'h42d87de9},
  {32'h4344e5b4, 32'hc3b87771, 32'h428636cc},
  {32'hc44da924, 32'h43141830, 32'hc31a802c},
  {32'h44e68893, 32'hc2d4ab9a, 32'h43477b06},
  {32'hc28d81da, 32'hc16c37d2, 32'h435fc9ab},
  {32'h44054578, 32'h41e0489c, 32'hc1f0c3fa},
  {32'hc3b2657e, 32'h425ad51f, 32'hc3c6a43f},
  {32'h44b6cb30, 32'h436bd598, 32'h4298560c},
  {32'hc3414e72, 32'hc296a3f3, 32'hc3ca9068},
  {32'h44dfb8f7, 32'hc383967a, 32'hc2ca0fea},
  {32'hc4e2d0b1, 32'h4318df58, 32'h4344d366},
  {32'h43ce75e0, 32'h4299dfd1, 32'hc2b9846a},
  {32'hc467cafa, 32'h4313797c, 32'hc3068e8c},
  {32'h44d910b0, 32'hc368512d, 32'h43404565},
  {32'hc4b397f6, 32'h42dccfe4, 32'h42bb3e23},
  {32'h45186d3b, 32'hc34445a4, 32'h439ae677},
  {32'hc4224386, 32'h42fa4548, 32'h436a3fc2},
  {32'h4508fd30, 32'h41852aa1, 32'hc2dc307b},
  {32'hc40d4930, 32'hc1df8c0c, 32'h42ed73f2},
  {32'h44bdda34, 32'hc2919a11, 32'h431af1f1},
  {32'hc3cea878, 32'hbe152f40, 32'h4292f980},
  {32'h449f3785, 32'h418ce402, 32'h42890bf4},
  {32'hc4d7a3ae, 32'h4407cfdd, 32'h4344fb5b},
  {32'h45233579, 32'h4389259f, 32'hc341beb3},
  {32'hc4488120, 32'h43c6feac, 32'h428a4d94},
  {32'h43f5fabb, 32'h43b6f21f, 32'h42078253},
  {32'hc389a1d4, 32'h3fd1ab2d, 32'h4201332b},
  {32'h4500d290, 32'h4238092d, 32'hc3f3c3f6},
  {32'hc5227640, 32'hc3b870ea, 32'hc38562d2},
  {32'h44d1ed50, 32'h40d43092, 32'hc32a1094},
  {32'hc484933e, 32'hc225d068, 32'h43c734dd},
  {32'h45052fc3, 32'hc314ebcb, 32'h42c57170},
  {32'hc2db2cce, 32'hc3813e0b, 32'hc2a28ce1},
  {32'h451bc10f, 32'hc32aa666, 32'h438700ab},
  {32'hc3a8c5f4, 32'h438c6012, 32'h42c08086},
  {32'h44916823, 32'h422466a9, 32'h439a5c01},
  {32'hc4be1db4, 32'hc2fdc2d4, 32'hc388a9af},
  {32'h43aa8bf4, 32'hc3063c08, 32'hc2d7a474},
  {32'hc48131fa, 32'hc116d5a4, 32'hc399abe5},
  {32'h44c01771, 32'h4315b6b6, 32'hc40585b1},
  {32'hc3f1d940, 32'h408320c0, 32'hc30ee1cc},
  {32'h44b79e30, 32'hc14ade42, 32'hc1b69b55},
  {32'hc52c8c13, 32'hc1202358, 32'hc20ffe00},
  {32'h4258b580, 32'hc3ec3a58, 32'hc3088327},
  {32'hc4840d16, 32'h43d93d8a, 32'h43609ec7},
  {32'h426bc3d0, 32'h433bff98, 32'hc34c8700},
  {32'hc4f6be70, 32'hc39b3bf7, 32'hc37f684c},
  {32'h43ff5b70, 32'h43259fba, 32'hc330d844},
  {32'hc4615ba6, 32'h42eb284a, 32'h43286f2a},
  {32'h44e905ca, 32'hc38c570e, 32'hc3254648},
  {32'hc3382584, 32'hc38548c3, 32'h41d29234},
  {32'h44e3fb22, 32'hc31f9a65, 32'hc1578a92},
  {32'hc494f0c7, 32'h4394eaad, 32'hc366ef1e},
  {32'h4442d196, 32'hc2e8479f, 32'hc2c22787},
  {32'hc4ef3ac4, 32'h43c72d50, 32'h43235530},
  {32'h436dc34c, 32'h4313a3ae, 32'h430eedf3},
  {32'hc508b819, 32'hc30263c1, 32'hc2d75a8d},
  {32'h44aa00e8, 32'hc2f052a9, 32'h42dd825a},
  {32'hc509d4b0, 32'hc3c557c8, 32'hc00a317c},
  {32'h44ff33c0, 32'hc2943f79, 32'hc28ebb1a},
  {32'hc39086f0, 32'h3ff65918, 32'hc18e5270},
  {32'h44261114, 32'h4070dacf, 32'h423f43c0},
  {32'hc42f811c, 32'hc393b4d1, 32'h43b4025c},
  {32'h44b4719a, 32'hc30f141d, 32'hc322cd0f},
  {32'hc46d59b1, 32'h438db122, 32'h43e1c46f},
  {32'h41e62f40, 32'hc3db3adb, 32'h43474699},
  {32'hc4bf12d0, 32'hc2805dc1, 32'h42f3f00d},
  {32'h44235bd0, 32'hc2ab2f82, 32'h439cc0c8},
  {32'hc49c8d90, 32'hc296f3f1, 32'h43cb34b2},
  {32'h449e6e04, 32'h437a8a1f, 32'hc45d1849},
  {32'hc4b3a110, 32'h41ca0712, 32'hc308ff8b},
  {32'h44e51860, 32'h432446f5, 32'h42a012cd},
  {32'hc4b22d1b, 32'hc2e4b119, 32'h42ecfc3f},
  {32'h432797d0, 32'hc3231666, 32'hc39348b4},
  {32'hc3d100e7, 32'h4278cd12, 32'h44053e8f},
  {32'h44cf00d7, 32'hc282d82d, 32'hc23825ec},
  {32'hc49adc3e, 32'h4213be92, 32'h42bddb88},
  {32'h43a02e08, 32'h434c5ee6, 32'h42500701},
  {32'h44f84f19, 32'hc30175e5, 32'h422270b8},
  {32'hc4be3784, 32'hc3397fdb, 32'h42735508},
  {32'h4401e214, 32'h4433c480, 32'h429d2cdb},
  {32'hc458d744, 32'hc315da35, 32'h427c436f},
  {32'h416fcc20, 32'hc3773693, 32'hc38575ed},
  {32'h41b315e0, 32'h438d55e4, 32'h43235160},
  {32'h43e8ef39, 32'hc1ae0e8c, 32'hc1b399e4},
  {32'hc4bd8a81, 32'h43a712ef, 32'hc2f7848d},
  {32'h44084cd0, 32'h41c9a5e0, 32'hc38b0c08},
  {32'hc48e0f62, 32'hc27e3092, 32'h4393e425},
  {32'h448f7243, 32'hc38f1c88, 32'hc1816008},
  {32'hc47ea212, 32'hc2775e83, 32'hc10512d9},
  {32'h449c169d, 32'h420114b6, 32'hc10662a0},
  {32'hc448d1c0, 32'hc3b0dea5, 32'hc3842e00},
  {32'h4412a243, 32'h432115be, 32'h43830c61},
  {32'hc4ddaf38, 32'h42acbf1e, 32'hc25549c6},
  {32'h42fecc48, 32'h4384ad0a, 32'hc3b9e750},
  {32'hc29b4d94, 32'hc3e06ade, 32'h428a0fbe},
  {32'h43f3b942, 32'h43116630, 32'hc262c7e0},
  {32'hc418a4e2, 32'hc3bbbecd, 32'h42b84533},
  {32'h4431b394, 32'h432b6f9b, 32'hc39ad527},
  {32'hc4d095f9, 32'hc3c5c571, 32'h436524c1},
  {32'h4495eca9, 32'h4325015c, 32'hc37b3a30},
  {32'hc500bd2b, 32'hc18c67c2, 32'h42a6974a},
  {32'h43dd12b0, 32'hc21b6d0f, 32'hc3e128d8},
  {32'hc50717b0, 32'h4318a47a, 32'h402a85f8},
  {32'h441e7862, 32'hc38f0b02, 32'h436eb02f},
  {32'hc3ec2c48, 32'h42e6b5db, 32'hc258efc8},
  {32'h44b6855d, 32'h430b0d06, 32'hc31a8b69},
  {32'hc383da55, 32'hc211a2f7, 32'hc05baa7b},
  {32'h43a45868, 32'hc35bd127, 32'h42cc6e2a},
  {32'hc457ba98, 32'hc33bda23, 32'hc28a0056},
  {32'hc32c2b4a, 32'h43b1a986, 32'hc3f4e516},
  {32'hc4f4902a, 32'hc3c1e353, 32'hc1eba74b},
  {32'h4351da80, 32'h43cee63c, 32'hc3178a47},
  {32'hc380a137, 32'h430f3083, 32'h41600b58},
  {32'h44fd2332, 32'h43517680, 32'h436e02d6},
  {32'hc4d407a4, 32'hc319fbca, 32'h430840e7},
  {32'h44c8b1de, 32'h43b39cb7, 32'h43619145},
  {32'hc40ba35a, 32'hc2936472, 32'h44117421},
  {32'h44fc8cdf, 32'h43bee25e, 32'hc34e15b9},
  {32'hc49c0aef, 32'hc2f79ffb, 32'h42bdc874},
  {32'h451b7587, 32'hc19016d4, 32'h43bb16d4},
  {32'hc3b07120, 32'h4289c9b2, 32'hc1bb5234},
  {32'h4506d306, 32'hc311f951, 32'h41f248a0},
  {32'hc40f4254, 32'h42bd8e6d, 32'hc3c62211},
  {32'h450a5486, 32'h415ef7d1, 32'hc3da2c38},
  {32'hc1d98400, 32'hc2b5abe2, 32'hc3956b14},
  {32'h44c025e2, 32'h4283c5b3, 32'h4389ba24},
  {32'hc42a00a4, 32'h42aeb83e, 32'h42aa14e2},
  {32'h430bfd92, 32'hc2811a05, 32'h43485924},
  {32'hc5046d24, 32'h43fb90ca, 32'h42d1cebc},
  {32'hc31e712c, 32'hc2d5920f, 32'hc2e37b46},
  {32'hc40b740e, 32'h43ee2859, 32'hc303a01f},
  {32'h44e10bb4, 32'h42b60171, 32'h42df7706},
  {32'hc4fa0215, 32'h4330b6b9, 32'h42f0350b},
  {32'h44db2b25, 32'hc33ce94b, 32'hc23e4e8c},
  {32'hc3a804f0, 32'h436c65e5, 32'h3f486950},
  {32'h440a13d8, 32'hc3133811, 32'h4348c92a},
  {32'hc430293a, 32'h432409ab, 32'hc39d699b},
  {32'h438b2060, 32'hc2b3a62b, 32'h41724249},
  {32'hc4c98dc6, 32'hc2eafa37, 32'hc3ad5d14},
  {32'h45101955, 32'hc31dc914, 32'h433a9af0},
  {32'hc4484683, 32'hc323eade, 32'h44169e6e},
  {32'h452681a5, 32'h43a90d91, 32'h43563531},
  {32'hc4c07b3c, 32'hc39df3ab, 32'hc1947a4c},
  {32'h44589135, 32'h43720cf8, 32'hc2180158},
  {32'hc41c4704, 32'hc353228e, 32'hc3b81b05},
  {32'h449298f8, 32'h439fde06, 32'h42aabe8a},
  {32'hc4930d5f, 32'hc26ddeb8, 32'hc32e3e5e},
  {32'h44f78938, 32'h4332b9f9, 32'h4376e9d8},
  {32'hc4e1bdae, 32'hc2b5a2b9, 32'h42ffc024},
  {32'h43fb4e18, 32'hc1e50f9a, 32'h4381670a},
  {32'hc49d87b5, 32'h43396ce5, 32'h439dd7c6},
  {32'h44644dd2, 32'h43acfeff, 32'h439218ff},
  {32'hc523bc4a, 32'h43afe38e, 32'hc3bfe3a1},
  {32'h4451c41e, 32'h3f91c240, 32'hc04128e0},
  {32'hc3e7381f, 32'h43702936, 32'hc2e154f6},
  {32'h43b1634b, 32'hc3dbc6da, 32'h43803d82},
  {32'hc4c23997, 32'hc31f3899, 32'hc2967e57},
  {32'h44c5641a, 32'hc28e4233, 32'h428f6e00},
  {32'hc30adf80, 32'h43623d50, 32'hc30b6b5a},
  {32'h442d2518, 32'h42454e50, 32'h429437d5},
  {32'hc4962225, 32'hc29d4ea0, 32'hc3a0c447},
  {32'h44f6b153, 32'hc3110713, 32'h43aaab26},
  {32'hc28b2ab0, 32'hc2e94fde, 32'hbd3eff00},
  {32'h42810e10, 32'h42285291, 32'h42af3d43},
  {32'hc49483c3, 32'hc2a35e36, 32'hc3002d6a},
  {32'h451cb0b9, 32'h42b13f88, 32'hc30c7f99},
  {32'hc3aa0e92, 32'hc39fba3d, 32'hc1dfa6f7},
  {32'h43e9c0f0, 32'h42fd3e4a, 32'h43151854},
  {32'hc47dae1a, 32'h42d8e070, 32'h438e8c93},
  {32'h44486c21, 32'h42be31d7, 32'h42a22832},
  {32'hc40e039a, 32'h428c43c6, 32'hc391d303},
  {32'h4392003c, 32'hc3820544, 32'h4312d997},
  {32'hc50428cb, 32'h43a3d747, 32'hc281f61f},
  {32'h44d61a00, 32'hc3400044, 32'h431fa1e4},
  {32'hc4160fbd, 32'hc04f5ac1, 32'hc3a6d474},
  {32'h44fe9ff2, 32'h4289e380, 32'hc2d77068},
  {32'hc44aabd0, 32'hc196f4d0, 32'h433a05b2},
  {32'h4488b54d, 32'h429d0ea4, 32'hc3f64306},
  {32'hc4f42f3e, 32'hc2e5adcc, 32'hc39320a9},
  {32'h43ac554a, 32'hc2ae92b7, 32'hc39a08cb},
  {32'hc4d813b0, 32'h42ccd25d, 32'hc2646b73},
  {32'h44f547f4, 32'hc395b6d1, 32'h41ad6713},
  {32'hc4a8ff8e, 32'hc3d7f111, 32'h4350ec15},
  {32'h44747b01, 32'hc2f1ba93, 32'hc28d4748},
  {32'hc4948612, 32'hc324e01c, 32'h42997952},
  {32'h44e7754d, 32'h42aa0ec9, 32'hc254e15c},
  {32'hc4769d88, 32'hc389d535, 32'h43b8bcb8},
  {32'h45134668, 32'h43beb1c3, 32'hc2fa4a4e},
  {32'hc49acca0, 32'h43a91e58, 32'h42cc82b8},
  {32'hc2c3cd0c, 32'h42160f23, 32'h4362f2be},
  {32'hc44a05d4, 32'h43ea7011, 32'hc2b58b0a},
  {32'h4474b610, 32'hc3999063, 32'h42937e18},
  {32'hc3bd6a20, 32'h429288b5, 32'hc3905f39},
  {32'h442eac4e, 32'hc39d5e3e, 32'hc20e522a},
  {32'hc4a9629e, 32'hc2fc9a79, 32'hc2b9ed82},
  {32'h451d3dad, 32'hc4105a4d, 32'h41d56e22},
  {32'hc46dc166, 32'h434ee855, 32'h4385520a},
  {32'h44e02bce, 32'hc3a29997, 32'h434733b3},
  {32'hc498fc6c, 32'hc3920f43, 32'hc191abc8},
  {32'h451352c8, 32'h434295f3, 32'hc29d8eb4},
  {32'hc344d35a, 32'h431da68d, 32'h4128e2fc},
  {32'hc3077980, 32'h42a0c506, 32'hc2861c59},
  {32'hc503822a, 32'h42809a30, 32'hc39fb375},
  {32'h45080d4b, 32'h432212ae, 32'hc26054d1},
  {32'hc4c02ec9, 32'h4182b9a4, 32'hc402024a},
  {32'h444b89fe, 32'h431a4a7e, 32'h4327e473},
  {32'hc46fc86e, 32'h432476ce, 32'h42ab334f},
  {32'h44375df0, 32'hc32a8c60, 32'h41ce733a},
  {32'hc40ed9c3, 32'h4377d7ad, 32'hc3979ef0},
  {32'h448121f3, 32'hc3993c5a, 32'hc26a99ce},
  {32'hc47cc51c, 32'hc1fc89ba, 32'hc3240b64},
  {32'h44099109, 32'h427ac1a2, 32'hc32be6c7},
  {32'hc508df14, 32'hc3682bc3, 32'h424354f0},
  {32'h4491afcb, 32'h429534ef, 32'h4308d988},
  {32'h42073d00, 32'h42b4b14c, 32'h43334394},
  {32'h4419e87b, 32'hc2e1df1d, 32'h41be9a2f},
  {32'hc383be08, 32'h43f568ae, 32'hc26c10aa},
  {32'h440bae42, 32'hc1e71f91, 32'hc38c922d},
  {32'hc43148bc, 32'hc2aac29f, 32'hc1c79d94},
  {32'h44919a6f, 32'h40d49b20, 32'h43fc946b},
  {32'hc5073eba, 32'h41556673, 32'h43020aa8},
  {32'h43b41450, 32'h43a9887b, 32'hc3077747},
  {32'hc48861c3, 32'h431cc525, 32'h42ac497a},
  {32'hc1d7bb80, 32'hc3ff608d, 32'h42122974},
  {32'hc5061bff, 32'h43cfc96a, 32'h43bfcc1c},
  {32'h44b089d1, 32'h428eaea8, 32'hc203e298},
  {32'hc40c12a9, 32'hc1ffbe61, 32'h430367f5},
  {32'h432d6b44, 32'h43eceaa1, 32'hc308e9b2},
  {32'hc44bf552, 32'hc24dd9f9, 32'hc29f935a},
  {32'h44afba5b, 32'h4406bd11, 32'hc3610903},
  {32'hc4fe8112, 32'h43876d2c, 32'h40f236c1},
  {32'h445c250c, 32'h4360c1f8, 32'hc14af2d2},
  {32'hc4ff6024, 32'hc2a4bcd7, 32'h42835f01},
  {32'h431fec50, 32'hc35c4dd8, 32'hc1b56e00},
  {32'hc35e890e, 32'hc35c7c3d, 32'h431d71cd},
  {32'h44bcad0a, 32'h418fe958, 32'hc1da3d50},
  {32'hc5077f12, 32'hc2be12a4, 32'hc2d19c6e},
  {32'h443d5544, 32'hc314bfaa, 32'h432ad7f6},
  {32'hc506ba70, 32'hc2d8037c, 32'hc2de0947},
  {32'h3f8df000, 32'h42be4c1d, 32'hc31d526f},
  {32'hc5054b2c, 32'h404965a8, 32'h43b4c6b6},
  {32'h43bb1ea9, 32'h435b65df, 32'h42ea46ff},
  {32'hc3fb18d8, 32'hc39ebf90, 32'h417f1c88},
  {32'h44e1d588, 32'hc088b2e5, 32'hc39fd6a5},
  {32'hc49e925a, 32'h4328beb5, 32'h4319b3a9},
  {32'h44058d66, 32'hc3233e00, 32'hc3a70482},
  {32'hc3b8adb0, 32'h437b6e3b, 32'h4345789a},
  {32'h447ac468, 32'hc27cd8eb, 32'hc3807327},
  {32'hc3a99e50, 32'hc2de9eb0, 32'h440ff737},
  {32'h437cee44, 32'hc28fabdb, 32'hc36974ff},
  {32'hc4be6717, 32'hc34518fa, 32'hc393c75b},
  {32'h44c8d184, 32'hc335e565, 32'hc2936d40},
  {32'hc44f8ba9, 32'h438ebc72, 32'hc15a9178},
  {32'h44a573b9, 32'hc3521bed, 32'h41521b27},
  {32'hc4e42b10, 32'hc2ff794c, 32'hc2111df3},
  {32'h44210206, 32'hc31a773a, 32'hc3d231e6},
  {32'hc490f1e2, 32'h4231e118, 32'h432e7cd2},
  {32'h450028bd, 32'h43c5b75c, 32'hc31a9eb4},
  {32'hc45f07c8, 32'h42a9c75f, 32'hc31ca179},
  {32'h450fbb16, 32'hc1c2fc43, 32'hc39fb638},
  {32'hc514dd70, 32'h436b79e0, 32'h432eab89},
  {32'h449618b6, 32'hc1bdaff8, 32'hc2efe4e0},
  {32'hc513b6aa, 32'h42e6b5af, 32'hc2d5961c},
  {32'h44cffb10, 32'hc24bdad6, 32'h4313d4da},
  {32'hc30e2f38, 32'hc32b1240, 32'hc309e13d},
  {32'h4432291a, 32'h43075073, 32'hc3366b99},
  {32'hc50439bb, 32'hc3805afe, 32'hc2357552},
  {32'h4410e2c6, 32'h42fdecb2, 32'h430e8ac7},
  {32'hc33f26b8, 32'hc35d2253, 32'h4300a982},
  {32'h44ac853e, 32'hc3028490, 32'hc2a15d5e},
  {32'hc4f23bc6, 32'h428fd5d4, 32'h430c03c4},
  {32'h447972a6, 32'h42864f9c, 32'hc199e65e},
  {32'hc46f7c98, 32'hc35b58bb, 32'h416eb00a},
  {32'h43b07a88, 32'hc3101768, 32'hc3504950},
  {32'hc49322c3, 32'hc3d5d47f, 32'h426d07e0},
  {32'h44b3846a, 32'h43805c33, 32'h434e3d3a},
  {32'hc4f8fca8, 32'hc2cd152c, 32'h429862ed},
  {32'h44929aff, 32'h4328f469, 32'hc28874fd},
  {32'hc38fd2dc, 32'h4304f934, 32'h435b3d8c},
  {32'h4502251c, 32'h433508cf, 32'hc3d9424d},
  {32'hc4be0bf0, 32'hc3426bd6, 32'h43b8bfbe},
  {32'h44baa8be, 32'h4393916d, 32'hc3aff78c},
  {32'hc4968196, 32'hc3392765, 32'h4140f052},
  {32'h449e614b, 32'hc36701c5, 32'hc22b5a4f},
  {32'hc50e088e, 32'h43be1fa9, 32'hc1f01fb6},
  {32'h44ea13fd, 32'hc3ff079c, 32'hc3ae13fb},
  {32'hc4e9c1e9, 32'hc268b6a4, 32'hc349b9f8},
  {32'h44f551e4, 32'hc39635ef, 32'hc37a0fb7},
  {32'hc49aa160, 32'h425b84d4, 32'hc1f05270},
  {32'h44e6e78f, 32'hc3965c3b, 32'h43fcfe0e},
  {32'hc482bcdb, 32'hc35ff3b7, 32'hc2a119ce},
  {32'h445e2b91, 32'h41d7bb3c, 32'h43207f62},
  {32'hc4bd1553, 32'hc3809cad, 32'hc20dd05b},
  {32'h44c251f6, 32'hc299de30, 32'hc279390b},
  {32'hc4e8b904, 32'hc335a2ae, 32'h43b4a84e},
  {32'h449b32e7, 32'hc28ddc9c, 32'hc300d340},
  {32'hc4e5171c, 32'h4302a9b0, 32'hc2bf6e2a},
  {32'h43fcdab2, 32'hc381d38f, 32'hc1563eaf},
  {32'h43c81a6e, 32'h437baeea, 32'h43151f49},
  {32'h42af7ba0, 32'h4363f907, 32'h415c1aa0},
  {32'hc4e28f20, 32'hc1960dd9, 32'hc39d1959},
  {32'h44ab499e, 32'hc251afa0, 32'h42e07b96},
  {32'hc4989fc4, 32'h438943f4, 32'h4206b0aa},
  {32'h44079f72, 32'hc29fc859, 32'h42dd7692},
  {32'hc3bd6578, 32'h438f696c, 32'hc228334e},
  {32'h44bf9e4e, 32'hc30e0bbb, 32'h429c64db},
  {32'hc4e1b3ba, 32'h439611c0, 32'hc2be149d},
  {32'hc31819e8, 32'h438bd29b, 32'hc33db746},
  {32'hc4184830, 32'hc34dc849, 32'hc3425f39},
  {32'h442ee0b0, 32'h43606646, 32'h435163e8},
  {32'h435d4390, 32'hc2dba550, 32'h429e6fa5},
  {32'h44f04ebf, 32'h42d7a9a6, 32'h4222ac90},
  {32'hc373a31b, 32'h43b59f66, 32'h43595432},
  {32'h43c2aa70, 32'h42e45a24, 32'hc2ee2985},
  {32'hc4c3b4e6, 32'h43505e3f, 32'h4324078e},
  {32'h4450fe89, 32'h43f73019, 32'h438493a2},
  {32'hc3dd88e5, 32'hc3096394, 32'h43846e8e},
  {32'h44c32348, 32'h41823b13, 32'hc2fa419f},
  {32'hc4aa4db8, 32'hc1667bad, 32'h42e1cae7},
  {32'h44a9208a, 32'hc3c7788e, 32'h4404f756},
  {32'hc48b6e59, 32'h4241d324, 32'h42e7cdda},
  {32'h451226a3, 32'h4321a19f, 32'h4397d365},
  {32'hc452f2b8, 32'h41ae2cd0, 32'h4226dc00},
  {32'h436fc830, 32'h441f7a28, 32'hc3714519},
  {32'hc49a3d64, 32'hc4138924, 32'h43eae6cd},
  {32'h4428d69b, 32'h43ec1c6e, 32'hc3480237},
  {32'hc41a428c, 32'h43504a12, 32'h42e7a439},
  {32'h4505a6fe, 32'hc276b935, 32'h42f5cc03},
  {32'hc4cc388c, 32'hc3cf4bb6, 32'h430e7607},
  {32'h4472eb98, 32'hc38c32bd, 32'hc21acb4e},
  {32'hc4b99e9b, 32'h4272f1d7, 32'h412766b4},
  {32'h450fcf05, 32'hc3a92f82, 32'h43a20e25},
  {32'hc43a2504, 32'h42a79839, 32'h41f54d37},
  {32'h445579c7, 32'h43532949, 32'h42eb3000},
  {32'hc406f9fe, 32'h438aa174, 32'hc254c323},
  {32'h43f2feba, 32'hc3a3f29f, 32'hc18160cf},
  {32'hc4fa2397, 32'h437f2965, 32'h4394e7c1},
  {32'h44ac93cc, 32'h42f2b1cc, 32'hc3223a5c},
  {32'hc43272b8, 32'hc39463fa, 32'h426f9375},
  {32'h4515c427, 32'h43652cef, 32'h43934d34},
  {32'hc4b551d1, 32'h438d1a14, 32'hc2184307},
  {32'h4493609e, 32'h419cea1e, 32'h436fe672},
  {32'hc509e799, 32'h439af89d, 32'hc197fefa},
  {32'h4497f02d, 32'h432847f6, 32'h41b043d6},
  {32'hc4a1205b, 32'hc4008951, 32'hc3a03df6},
  {32'h44964487, 32'hc1d63334, 32'hc3794c6e},
  {32'hc4d10c24, 32'h408a49bd, 32'hc3db8e4c},
  {32'hc0fc9100, 32'hc2c333b8, 32'h42808b07},
  {32'hc4b15613, 32'hc38efac7, 32'h42835f5e},
  {32'h44d78f27, 32'hc364e433, 32'h4373dcc1},
  {32'hc5059a93, 32'hc2a0fa0f, 32'hc32f28a2},
  {32'h430dc010, 32'h434a2c00, 32'h430238ed},
  {32'hc3f197f3, 32'hc316506e, 32'h42a3576d},
  {32'hc39c64f1, 32'h43e0022c, 32'hc3612555},
  {32'hc50f8214, 32'hc322a969, 32'h428f9b27},
  {32'h451701f9, 32'hc38f1011, 32'h41daa3a2},
  {32'hc4c4b3be, 32'hc3ab2689, 32'hc3f61361},
  {32'h4496949b, 32'hc33ce615, 32'hc38313bf},
  {32'h4202208f, 32'hc3012ac7, 32'hc2dcc8d1},
  {32'h435bbce0, 32'hc3e2b12a, 32'h43952314},
  {32'hc4faaafa, 32'hc3785f78, 32'h436d8704},
  {32'h44d1a773, 32'h42cbaabc, 32'hc34c7bc6},
  {32'hc47e531b, 32'hc3602267, 32'h42443c87},
  {32'h44b225c3, 32'hc366e81b, 32'h438b8b8e},
  {32'hc3c6ea75, 32'hc38ad46a, 32'hc3073971},
  {32'h4516c9b6, 32'h4399310b, 32'h4304758e},
  {32'hc4cd630f, 32'h4403e84d, 32'hc2aae7ed},
  {32'h4403626c, 32'hc385a817, 32'hc39d845c},
  {32'hc4b92f78, 32'h43a968a5, 32'hc32caaa1},
  {32'h44c5df71, 32'hc3ab9d58, 32'hc2717658},
  {32'hc4094857, 32'h4285db0a, 32'hc3d15845},
  {32'h4463642a, 32'h42ca824d, 32'hc417786c},
  {32'hc497bd36, 32'hc17dafab, 32'h430b809f},
  {32'h44e14e6c, 32'hc1b62552, 32'h42c9cc5f},
  {32'hc49bf431, 32'h43887bbb, 32'h433eaf98},
  {32'h449ce8ad, 32'h406de392, 32'hc1f0a774},
  {32'hc45eaa92, 32'hc3e65003, 32'hc2cccc96},
  {32'h450c0891, 32'hc273f83f, 32'hc291ad30},
  {32'hc5018595, 32'h43834061, 32'h43bed587},
  {32'h452182fd, 32'h43092b2f, 32'h42d4d344},
  {32'h42b7c080, 32'h43d6fdf6, 32'hc30a1711},
  {32'h4501c76a, 32'h41030184, 32'h4265ff43},
  {32'hc506dfe7, 32'hc28fd5b3, 32'h428f17ea},
  {32'h4505b9d7, 32'hc2b1bf50, 32'h431e2eba},
  {32'hc4dd8a44, 32'h4232be17, 32'hc28d1d95},
  {32'h4497aa3c, 32'h43270414, 32'h41f22104},
  {32'hc4cc2824, 32'hc3d44d1b, 32'h4391dace},
  {32'h44cdb5f1, 32'hbf8d0a4f, 32'h43e0c57c},
  {32'hc4b60844, 32'hc2b9a1d4, 32'hc1b9acc0},
  {32'h44b6fe5a, 32'hc3299224, 32'h42464c51},
  {32'hc51abb58, 32'hc1f67677, 32'hc1621fee},
  {32'h442a084e, 32'h42f2f8e2, 32'hc3a94380},
  {32'hc3ef17d0, 32'hc2fb903d, 32'h4138e2b8},
  {32'h44e2bb17, 32'hc1e328e6, 32'h43ca54a8},
  {32'hc4c38e77, 32'hc1ce0b43, 32'hc2a97b19},
  {32'h450278b9, 32'hc3f04421, 32'hc1e0294a},
  {32'hc50305ec, 32'hc1f885a3, 32'hc3935bf1},
  {32'h446aa660, 32'h43ac391b, 32'hc2e2526d},
  {32'hc4085c06, 32'hc2315f5c, 32'hc3201735},
  {32'h44eeb55f, 32'h43a3fef8, 32'h4285b366},
  {32'hc481f892, 32'hc3a63751, 32'h430239ad},
  {32'h44d929f7, 32'hc0bdf73e, 32'h41c6e90c},
  {32'hc50195c5, 32'hc14a1b04, 32'hc38c52eb},
  {32'h44e13d6c, 32'hc172395d, 32'h431501a4},
  {32'hc42077f5, 32'h42d8fc0a, 32'h42a6db3c},
  {32'h4484743e, 32'hc3b340c4, 32'hc2430f59},
  {32'hc400fb24, 32'hc23f733f, 32'h43bcd7b1},
  {32'h43cfa798, 32'h41f630e1, 32'h431d7a22},
  {32'hc4c80e8d, 32'hc3466d57, 32'h42edcabb},
  {32'h4422ace4, 32'hbfffae30, 32'h42c4be2c},
  {32'hc50510af, 32'hc2d2bd81, 32'hc2a8b9c5},
  {32'h44832d64, 32'h42a11886, 32'hc1980b7d},
  {32'hc483fefa, 32'hc1500b46, 32'hc359bb6b},
  {32'h44d170d6, 32'hc38ce124, 32'h422cd7fc},
  {32'hc48310f4, 32'h4384fa18, 32'hc3e5dd6a},
  {32'h44e91d56, 32'h4385696c, 32'hc29b3601},
  {32'hc3e739f2, 32'hc2e61a1b, 32'h41ecc958},
  {32'h44e65d67, 32'hc33a5795, 32'hc3174e9a},
  {32'hc4b46eaa, 32'hc40061a5, 32'hc3d90b4f},
  {32'h44fb5598, 32'h435d4909, 32'h41f184e2},
  {32'hc43957ca, 32'h432f52d7, 32'hbf6e2f00},
  {32'h44f9eb70, 32'hc31f5e67, 32'hc28daf67},
  {32'hc50ac645, 32'hc319f04b, 32'h42ff612b},
  {32'hc2d9c784, 32'hc3d59a09, 32'hc41de79a},
  {32'hc529c626, 32'h43efce86, 32'h436b44fc},
  {32'h437b84d8, 32'hc27f0673, 32'hc356f056},
  {32'hc2fe721f, 32'hc31f8821, 32'hc365cef0},
  {32'h444c1506, 32'h42c59992, 32'h42109275},
  {32'hc516cb03, 32'h438b65fd, 32'h428cafde},
  {32'h42f79440, 32'hc37e58db, 32'hc30bff09},
  {32'hc4255bf0, 32'h4383bcca, 32'h43946d2e},
  {32'h44b8c0ac, 32'h42783f50, 32'h432933fe},
  {32'hc4b38246, 32'hc2abdb03, 32'hc28f63e8},
  {32'h450a15b6, 32'h40dbadd4, 32'hc359051f},
  {32'hc43eec50, 32'hc3c8a035, 32'h42d38b87},
  {32'h44d6f3ff, 32'h439d25fb, 32'hc3e0e0fa},
  {32'hc5165577, 32'hc252e750, 32'h43e96cef},
  {32'h4506cfb7, 32'h4296ddf6, 32'h437159aa},
  {32'hc410ee88, 32'h438e9420, 32'h43497aef},
  {32'h44a74f9c, 32'hc35552b1, 32'hc339c797},
  {32'hc50c93eb, 32'hc33250ad, 32'h43a92c11},
  {32'h440f6670, 32'hc336855f, 32'hc31de7bd},
  {32'hc502c41c, 32'hc346df2c, 32'hc2340ec8},
  {32'h4332fde0, 32'hc20e808c, 32'h42024573},
  {32'hc4a7c61f, 32'hc3a1b97b, 32'hc308acc6},
  {32'h430fc318, 32'hc3ba89f1, 32'hc2bbdbf3},
  {32'hc4dc6aa7, 32'h419c45f8, 32'h4326d543},
  {32'h45091d26, 32'hc2175fc0, 32'h4346f85d},
  {32'hc3661bb0, 32'h42a2e7e5, 32'h4339f923},
  {32'hc237d200, 32'h42bd721d, 32'h4123c319},
  {32'hc3a591e4, 32'h4338a0e6, 32'h4270e205},
  {32'h449b1f61, 32'h43656b76, 32'h42ed284e},
  {32'hc485c56e, 32'h434ee370, 32'hc0555e80},
  {32'h44f46f42, 32'h41bd27f5, 32'h43349fc4},
  {32'hc3160b5f, 32'h4317c637, 32'hc18c59d9},
  {32'h435beccc, 32'h431dd784, 32'h41f00ec2},
  {32'hc30d9f00, 32'hc232671e, 32'h42d489ea},
  {32'h4342ddfe, 32'hc28cdbcd, 32'h4292b8a4},
  {32'hc48095dc, 32'h4355adff, 32'h4330e33e},
  {32'h45031ff5, 32'hc083c30a, 32'hc1ed22be},
  {32'hc49ff5d8, 32'hc357ef6a, 32'hc3e263b1},
  {32'h43064830, 32'h42a27ee9, 32'h401d6460},
  {32'hc425a2dc, 32'hc2bc499a, 32'hc1bdd4a4},
  {32'h4474b289, 32'hc3d4b39a, 32'hc3a45e24},
  {32'h4316ddf8, 32'hc3b9f2db, 32'h42f12984},
  {32'h438b50be, 32'h43199a61, 32'h436dae0e},
  {32'hc43d90e2, 32'h4204dd07, 32'h430df60b},
  {32'h44ca57be, 32'h41a4a931, 32'h4369a4b9},
  {32'hc50be20b, 32'hc35f5141, 32'h433a8142},
  {32'h44d44a6a, 32'h421027a0, 32'hc33c75c4},
  {32'hc4f19c3c, 32'hc28c2bd4, 32'hc3275f76},
  {32'h44ec22d7, 32'h43936d6c, 32'h4259063e},
  {32'hc4e0dd14, 32'h43c9fe1b, 32'hc3b20d6d},
  {32'h44bb6baa, 32'h43045b58, 32'h439a8596},
  {32'hc501ee4e, 32'h423ba6cc, 32'h42421c71},
  {32'h44a53b2e, 32'hc2bd0bba, 32'hc3a34691},
  {32'hc48ad1f7, 32'h434cb11d, 32'hc3771a30},
  {32'h44fd48ff, 32'hc3bec36e, 32'hc2468278},
  {32'hc436430e, 32'h4396cf08, 32'hc3a831d6},
  {32'h4491fa6c, 32'h43a2a1c4, 32'h44742b4f},
  {32'hc382a06a, 32'h431792c5, 32'h426e07f5},
  {32'h44c2bd28, 32'hc3b71fb5, 32'hc2e613dd},
  {32'hc32eaa81, 32'hc30e5aeb, 32'h433dda8f},
  {32'h41fa8b50, 32'hc346a223, 32'hc31937a1},
  {32'hc4d14f90, 32'h431ccdee, 32'h42fcd80c},
  {32'h42e52674, 32'h42868574, 32'h435a2c1a},
  {32'hc4e40232, 32'hc27d875b, 32'hc2bed323},
  {32'h450949f0, 32'hc341ba21, 32'h428306d9},
  {32'hc4344268, 32'hc34e7084, 32'h43c50c8c},
  {32'h4487a67d, 32'hc3da1a2f, 32'h433a4644},
  {32'hc4ec4430, 32'hc3619d5d, 32'hc38d6773},
  {32'h449521d5, 32'h431fa33a, 32'h43536f9c},
  {32'hc3261a3f, 32'h42a1952b, 32'h42fdd996},
  {32'h44b6c41e, 32'h42a497e6, 32'h4337e523},
  {32'hc45e7064, 32'h4247d32c, 32'hc3d58393},
  {32'h43d83dd0, 32'hc2665b6c, 32'hc32880c5},
  {32'hc3db9e1a, 32'hc3b8020b, 32'hc3663f5a},
  {32'h4507a16f, 32'h4266f0e5, 32'h4317766a},
  {32'hc49ec4ba, 32'hc33b5d49, 32'hc200adf5},
  {32'h44c28fc9, 32'hc2f2fbcb, 32'h423f5738},
  {32'hc43e39b3, 32'h43a4552c, 32'hc20e6e14},
  {32'h44b1ee00, 32'h4388bab3, 32'h433d95e1},
  {32'hc301a148, 32'hc30a2b70, 32'h436d49d1},
  {32'h438200e4, 32'hc3300bb5, 32'h426f855a},
  {32'hc43447df, 32'h4195045d, 32'hc33055f8},
  {32'h44d77621, 32'h43a7ffaf, 32'h433ced87},
  {32'hc4f2bc9f, 32'hc40fc671, 32'hc319f0d9},
  {32'h4320bbe4, 32'hc1d2ac3d, 32'hc2183910},
  {32'hc3dae9cb, 32'hc31c6d27, 32'hc37228e7},
  {32'hc348a4b7, 32'hc3597cac, 32'hc3c3ac05},
  {32'h442bbbba, 32'h439ecbbf, 32'h4399c9d8},
  {32'hc392ed48, 32'h42a3f101, 32'h42cb15d8},
  {32'h4478f08a, 32'h4331085b, 32'h436b3d11},
  {32'hc4417df8, 32'hc2aaf21e, 32'hc29b61c9},
  {32'h43a97d0e, 32'h409c5c6a, 32'h434edd79},
  {32'hc481644c, 32'hc3375922, 32'hc3bbe307},
  {32'h447564a4, 32'h43618e5f, 32'h431676b1},
  {32'hc4905eb9, 32'h43359a04, 32'hc1c52580},
  {32'h439165d0, 32'hc288edc6, 32'hc2d7c34e},
  {32'hc498bb64, 32'h431fb752, 32'hc3a5564a},
  {32'h44cbfdf0, 32'hc38315a7, 32'hc2a01068},
  {32'hc486eeea, 32'h4312a637, 32'hc3614433},
  {32'h43c0503c, 32'hc373ec0d, 32'h434dd902},
  {32'h432f3ab4, 32'h42b63736, 32'h43007d9a},
  {32'h449d03a4, 32'hc30c9e1d, 32'h411be6fd},
  {32'hc479a977, 32'h42d4b27f, 32'hc2e521f1},
  {32'h4501ed3d, 32'h430c1500, 32'h437534d7},
  {32'h4370c052, 32'h439fc314, 32'hc3588dd6},
  {32'h44498fa3, 32'h43257aa3, 32'h4269752c},
  {32'hc4225118, 32'h43a28524, 32'hc34236fb},
  {32'h44edbd0c, 32'hc2c26d27, 32'h431bcfea},
  {32'hc4b9474f, 32'hc2d188db, 32'h434b1d63},
  {32'h435c0a98, 32'h43519397, 32'hc2f630b7},
  {32'hc4c133c1, 32'h4207c2ad, 32'hc302cad6},
  {32'h43b071cc, 32'hc42979da, 32'hc1114719},
  {32'hc4e53833, 32'hc39ff8e9, 32'hc164db5f},
  {32'h434cf54f, 32'hc2eb2349, 32'h438f8d1e},
  {32'hc4ffa8f2, 32'hc38a7528, 32'hc3a0e178},
  {32'h4454f7b6, 32'hc34bdf06, 32'h439d7709},
  {32'hc491a73b, 32'hc301ed34, 32'hc3801a91},
  {32'h45064727, 32'hc39675ca, 32'hc0f7d1ca},
  {32'hc4cf3281, 32'hc355ad83, 32'hc3a13853},
  {32'h44835785, 32'h43096181, 32'h42ad4756},
  {32'hc498f910, 32'h43e18f29, 32'hc3835f7e},
  {32'h4505060e, 32'hc32d8353, 32'h42a75af5},
  {32'hc4b80976, 32'hc3cd399c, 32'hc2ce36e3},
  {32'h449b6596, 32'h422ffee2, 32'h4340c704},
  {32'hc4a943c6, 32'h3cfdc65e, 32'h4390119d},
  {32'h450ae7b6, 32'h42848e51, 32'h4336ecd8},
  {32'hc4055544, 32'hc2dd9ae4, 32'h412f6f8e},
  {32'h44f500fa, 32'hc1faeb56, 32'hc1e7224e},
  {32'hc482dd17, 32'hc2c5a72e, 32'h40cf1fd0},
  {32'h439b9439, 32'hc212be74, 32'h43c59397},
  {32'hc4dd0606, 32'h422c50d3, 32'hc1923b83},
  {32'h44f96e71, 32'h4265d83a, 32'h43a711df},
  {32'hc4cb4004, 32'hc2dbf744, 32'h4181b290},
  {32'h4376f3e2, 32'h4367d027, 32'h43f3da1f},
  {32'hc4f66286, 32'hc229d76a, 32'hc2988bfe},
  {32'h445e02ed, 32'hc3d1a93a, 32'h401267d0},
  {32'hc4e790f4, 32'h439b69fc, 32'h43f386b5},
  {32'h449f2735, 32'h434faf13, 32'h43320b4a},
  {32'hc48dd95a, 32'hc2771215, 32'h431dfd88},
  {32'h450667d5, 32'hc3ac1cd8, 32'h43911fff},
  {32'h42993858, 32'hc22bcb98, 32'hc19394f9},
  {32'h448b9cc9, 32'h4236380b, 32'hc3893fdc},
  {32'hc484f205, 32'hc272430c, 32'hc3397f4f},
  {32'h4500d68e, 32'hc2a35f81, 32'hc39b654e},
  {32'hc465a33c, 32'h434e9d19, 32'hc30e8984},
  {32'h4398b4b8, 32'h425221dc, 32'h43aa8044},
  {32'hc49031d8, 32'hc2d3e9f4, 32'h431a5c5a},
  {32'h4474f848, 32'h4345c824, 32'hc2aa5cf2},
  {32'hc2314f80, 32'hc288aa62, 32'hc29477a2},
  {32'h4443faf9, 32'h42abddbc, 32'hc3339ade},
  {32'hc4cfbebb, 32'hc3b90d22, 32'h4383cff2},
  {32'h44db05ff, 32'h416b0dba, 32'h422a032d},
  {32'hc4566010, 32'h42f4eefa, 32'h4357e166},
  {32'h44d9888d, 32'h439d893e, 32'hc2f0a7fa},
  {32'hc4a383bf, 32'hc2d288f3, 32'hc2ad6326},
  {32'h44c69e61, 32'hc2febf7a, 32'hc2e41715},
  {32'hc5076440, 32'hc2609bf8, 32'h42e268be},
  {32'h442a3de4, 32'h43cbe631, 32'h43397d73},
  {32'hc4d9cae1, 32'h43018572, 32'h421c089d},
  {32'h43de7580, 32'h42646742, 32'h42929fae},
  {32'hc492611a, 32'h4265ff7d, 32'hc2d39f43},
  {32'h45023e07, 32'h43147e18, 32'hc27043d4},
  {32'hc3115c25, 32'hc2ad9dc7, 32'h43f26faf},
  {32'h44e1ee7a, 32'h4283bd03, 32'hc3a973e2},
  {32'hc4d2463f, 32'hc2a350b9, 32'hc212d244},
  {32'h44a8c731, 32'h433cb812, 32'h433a9b94},
  {32'hc4bb4976, 32'h4206fafc, 32'hc3405dfe},
  {32'h44c909b4, 32'hc35848cd, 32'h41f142b8},
  {32'h43c91f9a, 32'h406b7577, 32'h4337d85c},
  {32'h44ca75b2, 32'h41709fad, 32'h43a868e8},
  {32'hc48ee9ae, 32'hc38015f2, 32'h41e4da5b},
  {32'h444a44fc, 32'hc387fd07, 32'hc2b8b747},
  {32'hc38d71b8, 32'h43747803, 32'h437f740c},
  {32'h44f1f004, 32'h43206065, 32'hc31ae9ba},
  {32'hc2c45c48, 32'hc2d3c48b, 32'h431e200e},
  {32'h44a4210d, 32'h42d7b1ca, 32'hc2f9697d},
  {32'hc47e40f8, 32'hc325c415, 32'hc34c576e},
  {32'h440b7ce9, 32'hc39ea64e, 32'h4324e8c6},
  {32'hc505188f, 32'hc352f979, 32'h42a7612f},
  {32'h44c54e34, 32'hc37c6aca, 32'h43c60a61},
  {32'hc4cbf76b, 32'hc2d57bc8, 32'hc4081158},
  {32'h44ad4542, 32'h430e49e8, 32'h42905d71},
  {32'hc433d3b0, 32'h43134788, 32'hc3afcd70},
  {32'h44746ada, 32'hc2d4ed8c, 32'hc351bcb7},
  {32'hc3d2a2a7, 32'hc383e905, 32'hc1348b1f},
  {32'h44e198ab, 32'hc15d24b5, 32'hc310c89d},
  {32'hc4909ef5, 32'hc2971c8b, 32'hc27b5834},
  {32'h44938151, 32'h43bef1f4, 32'hc1ff3370},
  {32'hc429c164, 32'h41403666, 32'h433e1ea0},
  {32'h44867837, 32'h439b33d6, 32'h41a85c94},
  {32'h42d9d080, 32'hc2b513da, 32'h41a67ff3},
  {32'h44d51fb6, 32'hc27c59c5, 32'h42129e2f},
  {32'h4340b68c, 32'hc34016f7, 32'h43703508},
  {32'h44a69490, 32'hc1f9f19c, 32'hc158906c},
  {32'hc4fbd046, 32'h43a00bb8, 32'h415cf22d},
  {32'h44f7bb39, 32'hc298a589, 32'hc1eda92e},
  {32'hc479ad9b, 32'hc3c1883e, 32'h438b7069},
  {32'h44b22fb7, 32'hc2d17ce5, 32'hc2a6eb69},
  {32'hc3389e98, 32'hc2d12b93, 32'hc1fc6998},
  {32'h446f4676, 32'h437caa75, 32'hc2a822cb},
  {32'hc3893138, 32'hc2c53dbb, 32'h43907efd},
  {32'h44d14819, 32'hc282544a, 32'hc416df1b},
  {32'hc472e4c5, 32'h42c815c1, 32'h43456dbe},
  {32'h44a97480, 32'hc2e56eeb, 32'hc3b506a6},
  {32'hc4bae95e, 32'h430cda30, 32'hc276ede4},
  {32'h44f91227, 32'hc17f55ed, 32'hc3777386},
  {32'hc4c178cf, 32'hc02da89c, 32'h438d4d10},
  {32'h44bc029d, 32'hc3c93a0b, 32'h4367ea26},
  {32'hc3183c20, 32'h424b5b98, 32'h4340325f},
  {32'hc22b4500, 32'hc30bef90, 32'h420715f4},
  {32'hc4ce251e, 32'hc34a5076, 32'h43de3ad2},
  {32'h44ce038f, 32'h430f9601, 32'h42d20327},
  {32'hc4d759f1, 32'h4338f50f, 32'h41ee6b97},
  {32'h44975391, 32'h42957195, 32'hc37facbe},
  {32'hc3371ca8, 32'hc3dc4986, 32'hc280b4e3},
  {32'h4408dd6d, 32'h419139fa, 32'h43ac87d2},
  {32'hc3805d98, 32'h4215a397, 32'h42935f07},
  {32'h45008b86, 32'hc350a151, 32'hc3348ae4},
  {32'hc5155a5a, 32'h4278e0cc, 32'hc206e04d},
  {32'h44c792d1, 32'h42136e42, 32'h43f372b0},
  {32'hc42e2939, 32'hc21f57b1, 32'h4305e11d},
  {32'h450433fc, 32'hc32ffabc, 32'hc39233f1},
  {32'hc43d022c, 32'h422e2b51, 32'h43462ab8},
  {32'h448814a7, 32'hc37074d0, 32'h4397b9c1},
  {32'hc4e229a7, 32'hc0aa6f08, 32'h43f134fb},
  {32'h4489de38, 32'h41b9a6ce, 32'hc12f0916},
  {32'hc459dd86, 32'h429f56e2, 32'hc3d25112},
  {32'h44b7e1fc, 32'h41e8a7bf, 32'h4393bf3c},
  {32'hc4d25a90, 32'h4341991e, 32'h43b0bd23},
  {32'h44d19656, 32'hc365dab3, 32'h432c9ff1},
  {32'hc4e6dce8, 32'hc20a8052, 32'hc333f77b},
  {32'h4484fba2, 32'hc2f0b725, 32'hc23a6e02},
  {32'hc4b06b33, 32'h4364c515, 32'hc3618f35},
  {32'h450c2f43, 32'h43579fcb, 32'h434b828e},
  {32'hc4da38ae, 32'h4331d29c, 32'h439fdb1c},
  {32'h44e6a284, 32'hc28cafb0, 32'h43b95d1c},
  {32'hc49988c3, 32'hc28be916, 32'h422bab04},
  {32'hc2899620, 32'h4333e6b4, 32'h438dc874},
  {32'hc4b0749d, 32'h4138764a, 32'h4366d984},
  {32'h45041244, 32'h434502ed, 32'hc28421d8},
  {32'hc3cc07d4, 32'hc39fe2ac, 32'h439ac8a2},
  {32'h44727836, 32'h43bb22d4, 32'hc3f34ddd},
  {32'h4209d218, 32'hc3748232, 32'hc30c0c24},
  {32'h4494a32e, 32'hc2c2c36d, 32'h415c9fa8},
  {32'hc3e4410c, 32'h43753541, 32'h438715aa},
  {32'hc2331c30, 32'hc1e190b7, 32'hc3ac08e8},
  {32'hc4797c37, 32'hc159ed44, 32'h3fad67b0},
  {32'h44566220, 32'hc389ba46, 32'hc409d7d3},
  {32'hc3bb6a10, 32'hc3527092, 32'h40946660},
  {32'h44a1fa75, 32'hc2df9295, 32'hc31c80e3},
  {32'hc3e11f22, 32'hc364e266, 32'hc3c52cba},
  {32'h4430e8ba, 32'hc3c19555, 32'hc302e424},
  {32'hc4380cd8, 32'h4314ad55, 32'hc36a7809},
  {32'h440f5be4, 32'hc3842020, 32'h41fbd8e6},
  {32'hc396780b, 32'h433f6cad, 32'hc2c01790},
  {32'h4464dadd, 32'h4366b167, 32'h43a0815a},
  {32'hc50cc8af, 32'h432f5dd0, 32'h42a2de10},
  {32'h450717b1, 32'hc1f235ac, 32'hc2c6d2c5},
  {32'hc46ec4dc, 32'hc3415786, 32'h432b82f7},
  {32'h44f697fc, 32'h41536d96, 32'hc3264f53},
  {32'hc3a80b28, 32'hc28e0074, 32'h42adfd57},
  {32'h44de90b3, 32'h43ad7984, 32'h433cb4f6},
  {32'hc3271a1e, 32'h440163e5, 32'h419ca05f},
  {32'h448982d6, 32'hc352ece3, 32'h4242bc75},
  {32'h435aa3f0, 32'h42f4c73c, 32'hc2b409ce},
  {32'h4501b447, 32'h42b53277, 32'hc3668b2b},
  {32'hc490da33, 32'hc24b3a36, 32'h43c168c8},
  {32'h44b88df4, 32'hbf9087e4, 32'hc36f10d8},
  {32'hc4e34286, 32'h42e53d83, 32'h436c2484},
  {32'h4515d789, 32'hc252ea94, 32'hc21d3faa},
  {32'hc367f670, 32'h43302bb7, 32'h42b7fc58},
  {32'h44b95b86, 32'h43e495f0, 32'h41600ad4},
  {32'hc44c33e4, 32'hc2e972ea, 32'h408aeb43},
  {32'h43a9b4c4, 32'h433db73c, 32'h438d434e},
  {32'hc48c281a, 32'h43b465dd, 32'h430081b2},
  {32'h44d5c76d, 32'hc3dfb53f, 32'hc2900772},
  {32'hc493c5db, 32'hc2941b58, 32'h4313c5eb},
  {32'h450550a3, 32'hc1c73dd5, 32'h439079c5},
  {32'hc4cb9496, 32'hc3d0fb03, 32'h42c441f3},
  {32'h45152aae, 32'h43b2cdb3, 32'h44070956},
  {32'hc4eace83, 32'h436da5b3, 32'hc2ec3f3f},
  {32'h4500952a, 32'hc323a4ba, 32'h43a07b3b},
  {32'hc41e3586, 32'hc2382f2a, 32'hc26516ca},
  {32'h42b44bf0, 32'h42edda3b, 32'h4340c740},
  {32'h416a8d7c, 32'hc109bd06, 32'hc2a7f7f3},
  {32'h4442f893, 32'hc3cf85a6, 32'h435ba022},
  {32'hc4d8ecdf, 32'hc3c701a5, 32'hc2f49fb9},
  {32'h44be69ee, 32'h43178e75, 32'h4311b51b},
  {32'hc4edb5ac, 32'h417c5006, 32'h42728797},
  {32'h44405e84, 32'hc38cd133, 32'h42bf2efe},
  {32'hc483e872, 32'h42fc22f9, 32'h4165db49},
  {32'h445f7bb1, 32'hc282900d, 32'hc3ec09bf},
  {32'hc4114bfa, 32'hc1f96a6e, 32'h425a19d8},
  {32'h450cf864, 32'hc33cfb1d, 32'hc0d2a159},
  {32'hc33da668, 32'hc28fa6b1, 32'hc3a7dac3},
  {32'h44ee6b30, 32'hc29c1cfd, 32'h42c6e996},
  {32'hc29ef0d1, 32'h423d9383, 32'hc40c1c67},
  {32'h4435af44, 32'h41881bc6, 32'h428e3e81},
  {32'hc3adfd78, 32'h438d73f6, 32'hc008d634},
  {32'h44c6ad70, 32'hc2fd78fe, 32'hc28078f1},
  {32'hc4446b14, 32'h429c31ac, 32'h438101ea},
  {32'h44d09127, 32'hc3677c46, 32'h42cd5efb},
  {32'h415dfc28, 32'hc2c4b32e, 32'hc408fc5a},
  {32'h44992b09, 32'h436405fe, 32'h4321dd56},
  {32'hc3c56050, 32'hc1c3873f, 32'hc3851dea},
  {32'h4462467d, 32'h413cd0e4, 32'hc1c15cd3},
  {32'hc50420c5, 32'hc365e3e6, 32'hc304500a},
  {32'h440dc996, 32'h43501294, 32'hc3319b07},
  {32'hc49105ef, 32'hc2180ddb, 32'h4324d5da},
  {32'h44f3a95a, 32'h43a38295, 32'hc3a6cf9c},
  {32'hc37cd820, 32'hc3a4417f, 32'hc249d229},
  {32'h442017d0, 32'h43d8d490, 32'h42104e1b},
  {32'hc43bf90c, 32'hc235e74f, 32'hc31c03d1},
  {32'h44f892eb, 32'h438036c3, 32'h4245eb19},
  {32'h42c86e1b, 32'hc33e4840, 32'hc13e1de5},
  {32'h450a753c, 32'h439260e4, 32'hc24db9f1},
  {32'hc4fc1797, 32'hc245d42e, 32'h43030c1e},
  {32'h435cfc28, 32'h43cdc7df, 32'hc35cce1f},
  {32'hc432a68a, 32'h434edc0d, 32'h42046bf8},
  {32'h44eebc25, 32'hc35b220e, 32'h435adc92},
  {32'hc49f59fc, 32'hc385782a, 32'hc2bc266b},
  {32'h44f6c476, 32'h439d1032, 32'h4386ac88},
  {32'h42887d2e, 32'h434708af, 32'h420ddc81},
  {32'h444c9d48, 32'h41d03eb6, 32'hc2ae877d},
  {32'h426120a8, 32'h431fe9e2, 32'h431dbbfb},
  {32'h44f8e2a2, 32'h431a7d48, 32'hc2ade4af},
  {32'hc4ffe2ce, 32'h423fbe67, 32'hc2bbc884},
  {32'h44fbc92b, 32'hc384b5d1, 32'hc2062343},
  {32'hc4eac37a, 32'h43c2e971, 32'h4276c4e6},
  {32'h44f77956, 32'hc3c118f3, 32'hc28b6583},
  {32'hc50a8f32, 32'hc228f033, 32'h435da700},
  {32'h43af0170, 32'hc1611025, 32'h43ba24bf},
  {32'hc4a9d4dd, 32'hc32dcd3d, 32'h44012672},
  {32'h44da8fa7, 32'hc3a59d8a, 32'hc2189c8a},
  {32'hc4ca368b, 32'h4221bf99, 32'h427f9f0f},
  {32'h44ec8432, 32'h42a523e4, 32'h41b48e00},
  {32'hc5047303, 32'hc2b594b6, 32'hc3db56b5},
  {32'h44c4520f, 32'hc2eef910, 32'h42ad5044},
  {32'hc34a4eb8, 32'h4236acb2, 32'hc3561435},
  {32'h44a7ac32, 32'h42bca764, 32'h417153ce},
  {32'hc45a1871, 32'hc2340d37, 32'h439a088b},
  {32'h44527734, 32'h43edf2d3, 32'hc324585a},
  {32'hc4229339, 32'hc23085ea, 32'h428cc4c0},
  {32'h444b5aa4, 32'h439af157, 32'h43a9ab06},
  {32'hc514c424, 32'h4379526c, 32'hc186f3c6},
  {32'h4401a2be, 32'hc21143a8, 32'h42b70d25},
  {32'hc194a8c0, 32'hc39b6994, 32'hc1eb9fa4},
  {32'h430a76bb, 32'h43649245, 32'h43245d0b},
  {32'hc3f7b6b4, 32'hc3a4a869, 32'h43121bcb},
  {32'h44ee863a, 32'hc21e653b, 32'h4382578f},
  {32'hc2bd99d8, 32'h43360d6c, 32'hc0f9effb},
  {32'h44d45ee6, 32'h4339f84c, 32'h4371d59a},
  {32'h41f22b42, 32'h4340d35c, 32'h421ff5be},
  {32'h44cbe42a, 32'hc30cf2cf, 32'hc2ef2172},
  {32'hc50331ea, 32'hc353e112, 32'h42e2690f},
  {32'h44656af4, 32'hc20ec93f, 32'h4202f56f},
  {32'hc48bffda, 32'h4333e989, 32'hc3b9d759},
  {32'h44b1f60f, 32'h40c57084, 32'h428a6048},
  {32'hc3e814e4, 32'h43bab5c4, 32'h4100af6f},
  {32'h44fc2f90, 32'hc3604995, 32'h422c3b57},
  {32'hc4de789e, 32'h42e9fed9, 32'hc37f35de},
  {32'h448ae712, 32'h4388b49e, 32'hc3a0f855},
  {32'hc4cfe88e, 32'h4302e194, 32'h43012cb4},
  {32'h450ed1e6, 32'h430e6e76, 32'hc2b43987},
  {32'hc47dfda4, 32'h42c17bf6, 32'hc320e599},
  {32'h445fce22, 32'h41a84073, 32'hc2cec411},
  {32'hc411ec66, 32'h43b52fd2, 32'h42282706},
  {32'h411b0500, 32'hc32fc22a, 32'h4371019a},
  {32'hc4347ee8, 32'hc391656b, 32'h4297b701},
  {32'h44ac44b6, 32'h42d6012f, 32'h43454db4},
  {32'hc46cedec, 32'hc3423bb9, 32'hc179b558},
  {32'h43b7ebcc, 32'h4060bf6c, 32'hc274de27},
  {32'hc3544888, 32'h422edb81, 32'h4363ef14},
  {32'h44cec29f, 32'hc2cefd5b, 32'hc3414c59},
  {32'hc48656f6, 32'hc3e619cb, 32'h427532f9},
  {32'h44b0c9e6, 32'h4399de6f, 32'h4336c50f},
  {32'hc4c80934, 32'hc2a7c476, 32'hc3301ad1},
  {32'h4518e054, 32'h41e2c974, 32'h4300a2d8},
  {32'hc3eb0922, 32'hc3826c2c, 32'hc3adc2e7},
  {32'h4267e0e0, 32'h42f59658, 32'hc1ea9296},
  {32'hc4220aef, 32'h43e1b19e, 32'h42f383d1},
  {32'h44d49a46, 32'hc38b4db5, 32'h42feccf2},
  {32'hc50129aa, 32'hc31daa3c, 32'hc2fc3a6f},
  {32'h444c6b80, 32'hc1ee4ab4, 32'h43a4c2f8},
  {32'hc49c3f2c, 32'hc256092a, 32'h439e653e},
  {32'h439a20c3, 32'h43bb1ac7, 32'h43c09e1b},
  {32'hc45ab46e, 32'hc2b3c074, 32'hc36345df},
  {32'h43dd0230, 32'h430c5371, 32'hc2ad6843},
  {32'hc4f786cc, 32'h4225ad09, 32'h4217a06f},
  {32'h44b39343, 32'hc2a42966, 32'h43452ce5},
  {32'hc4832e63, 32'h437f284e, 32'h4395dddf},
  {32'h44100d90, 32'hc2e288e5, 32'h4239cf08},
  {32'hc4ef1210, 32'hc1d96194, 32'h4244012a},
  {32'h44e9b6f8, 32'h41b9e486, 32'hc3b0c911},
  {32'hc5097cd8, 32'hc3863186, 32'hc2fdc823},
  {32'h44759958, 32'h43a7d021, 32'hc34bcca5},
  {32'hc50e70f9, 32'h4394d7d8, 32'h434e99ff},
  {32'h44c5c2e3, 32'h4380e80a, 32'h421f4d01},
  {32'hc43bffd6, 32'h4310b75a, 32'h43a59768},
  {32'h44bb7373, 32'h421ab31e, 32'h4330fd0f},
  {32'hc29d4f21, 32'hc246b69f, 32'hc3073fe1},
  {32'h435ae862, 32'h43dad1bb, 32'hc1d2ed6a},
  {32'hc49d3f97, 32'hc190bf79, 32'hc36cd485},
  {32'h45148d2d, 32'h440e09e6, 32'h427d5e74},
  {32'hc4fb68d0, 32'h43740130, 32'hc2f2ccab},
  {32'h445ea049, 32'h439b9b66, 32'h433749a0},
  {32'hc5013005, 32'hc3c68ecf, 32'h43743e27},
  {32'h44d8ae90, 32'hc2b38a88, 32'h43af71f7},
  {32'hc43342e8, 32'hc23e4b4a, 32'hc2127d9a},
  {32'h44cad13e, 32'h43975d1f, 32'h4341a9d9},
  {32'hc4071314, 32'hc314b14a, 32'h424be723},
  {32'h4485ee79, 32'hc3449fea, 32'h42b7f119},
  {32'hc4daeb37, 32'hc34253d9, 32'h41e22e9e},
  {32'h43c2edc8, 32'h433ca409, 32'h4399c977},
  {32'hc4883856, 32'h4315f371, 32'h437ee478},
  {32'h44e18ca3, 32'h4374ebc1, 32'h433c5f9e},
  {32'hc4300020, 32'hc3b820f5, 32'h42f361d7},
  {32'h43d8e2e0, 32'h437e15f9, 32'hc1fa91be},
  {32'hc46c2238, 32'hc360a727, 32'hc32181d9},
  {32'h445730a0, 32'hc3515340, 32'hc327ea8f},
  {32'hc4adb3dd, 32'h426a39ff, 32'hc3a63471},
  {32'h44d4dc20, 32'hc3a27fe7, 32'hc2a2ada1},
  {32'hc4adbf0c, 32'hc229762e, 32'hc374f5fd},
  {32'h447dd2b6, 32'hc2ac4520, 32'h3dbcf000},
  {32'hc43d7584, 32'hc2334308, 32'h439547d1},
  {32'h44f73cce, 32'h430712e0, 32'h43286c4a},
  {32'hc241cec0, 32'hc2c9fac8, 32'h41347236},
  {32'h450d943f, 32'hc33f3efd, 32'hc27b8ed4},
  {32'hc472ac3a, 32'hc2d381cc, 32'hc29c4b21},
  {32'h43c067a4, 32'hc3565c59, 32'h4220d17f},
  {32'hc3aecb30, 32'h41c3b500, 32'h409986e1},
  {32'h4322141f, 32'hc2aa246e, 32'hc32296b8},
  {32'hc48c855c, 32'hc3108653, 32'h43f234bc},
  {32'h43ca9545, 32'h42b41d3f, 32'hc29a7ad9},
  {32'hc39f0bd4, 32'h43882ba2, 32'hc320c8fc},
  {32'h450bebde, 32'hc3f6ed29, 32'hc1cb9514},
  {32'hc4c38db8, 32'hc373c710, 32'hc37b529e},
  {32'h44e42489, 32'h435b2727, 32'h420d39b8},
  {32'hc502d700, 32'hc34ec1b5, 32'hc1dca548},
  {32'h44507ae4, 32'hc34b6ec8, 32'hc3de90f6},
  {32'hc3846b93, 32'h428c087b, 32'hc38b05a4},
  {32'h45041740, 32'hc2a9d6a4, 32'h4382f3c6},
  {32'hc4619f40, 32'h42978186, 32'hc2cbb894},
  {32'h43f70112, 32'hc3364234, 32'h420d14b6},
  {32'hc4ef9038, 32'h420bc4aa, 32'h4362cdd5},
  {32'h451682a2, 32'h42ee40d1, 32'hc3487ccf},
  {32'hc4d48177, 32'hc29273eb, 32'hc41cc628},
  {32'h44dedf4c, 32'hc2fcda3e, 32'h430c739f},
  {32'hc3b5a018, 32'h43831bbf, 32'hc34d780c},
  {32'h444fbb33, 32'h428abc18, 32'h42acd4a7},
  {32'hc4413a8b, 32'hc333fd2a, 32'hc35404f6},
  {32'hc25dfb60, 32'h4291a30c, 32'h42514421},
  {32'hc30cd9f8, 32'h427faf12, 32'h43a8db1c},
  {32'h448a509d, 32'h42f0c0bd, 32'h43213438},
  {32'hc4c05b97, 32'hc38ef5ec, 32'hc1d9e247},
  {32'h44e72965, 32'hc381780e, 32'hc197b7e9},
  {32'hc30e49d0, 32'h431a34d7, 32'h438bfbf0},
  {32'h43902100, 32'hc2596f8c, 32'h427083ad},
  {32'hc4fac5af, 32'h43392d16, 32'h423ef4f0},
  {32'hc21b9020, 32'hc3a0bc4e, 32'hc31e98c6},
  {32'hc3a5f750, 32'h4375352e, 32'hc313a439},
  {32'h4504aa9e, 32'h40addefc, 32'h42098d48},
  {32'hc4cc4500, 32'h428f7d4e, 32'h4313cebd},
  {32'h450b0249, 32'h42933a71, 32'hc3927bcc},
  {32'hc48165ec, 32'hc3220386, 32'h439b602f},
  {32'h45026a5f, 32'h43e989c7, 32'h43646f01},
  {32'hc4b4da43, 32'h42979456, 32'hc3097977},
  {32'h44e63997, 32'h42d3f207, 32'hc2b20bfe},
  {32'hc5298fea, 32'hc3879d79, 32'h4330e3c8},
  {32'h44a52fbf, 32'h41503060, 32'hc277a500},
  {32'hc418a6bc, 32'hc36075c0, 32'h419c8903},
  {32'h44f13f59, 32'hc28a8c11, 32'h439edce3},
  {32'h431576d5, 32'h42e46ecf, 32'h42acbbed},
  {32'h4511f4e4, 32'h43869c3c, 32'hc32ff5a5},
  {32'hc52227a1, 32'h41f93578, 32'h43b408f2},
  {32'h44e3210f, 32'hc3764d09, 32'hc2c0e176},
  {32'hc4972e90, 32'hc3acd6fc, 32'h43a8e94f},
  {32'h446e7cc8, 32'h435147b3, 32'h43789323},
  {32'hc4f863ea, 32'hc1bb0bf0, 32'h4384cccd},
  {32'h4385f623, 32'h4208b7ab, 32'h435a8d69},
  {32'hc4e2b9f9, 32'hc2a0706d, 32'h439689aa},
  {32'h450bff0c, 32'h439048ee, 32'hc31edf7c},
  {32'hc40afb6b, 32'h4329605e, 32'h42e56098},
  {32'h44d0c4c1, 32'hc1aa82b4, 32'hc2d0a291},
  {32'hc485e11a, 32'hc33a864b, 32'hc2f7bb9c},
  {32'h448b3f68, 32'h434f786a, 32'hc41ddd66},
  {32'hc4a1d292, 32'h41801e19, 32'hc326bf81},
  {32'h43e1bd68, 32'h42673f40, 32'hc3f00838},
  {32'hc4ecd58b, 32'hc2b1a4cd, 32'hc2bbac7d},
  {32'h4495df2c, 32'hc305784d, 32'h421922fa},
  {32'hc4bead3e, 32'hc1f57bc9, 32'h43c59965},
  {32'h44fbe3ca, 32'hc2388fd6, 32'h42bc9b06},
  {32'hc404fa5e, 32'hc382eb75, 32'hc1cb0429},
  {32'h446be172, 32'h43c870eb, 32'h43165384},
  {32'hc4d3b847, 32'hc29350e4, 32'h42ae7dd6},
  {32'h44eba9d6, 32'hc32d3a6a, 32'hc2d927b6},
  {32'hc5031d0d, 32'hc354834c, 32'h43d4d5f1},
  {32'h4510c524, 32'h42e4166e, 32'h41ddb1be},
  {32'hc50caa6d, 32'hc1cb31d6, 32'hc3009668},
  {32'h43e996d4, 32'h43613400, 32'h4299c65c},
  {32'hc3bdf790, 32'hc23df682, 32'h435892ee},
  {32'h43a8e4b4, 32'h433b368b, 32'hc3124bb2},
  {32'hc400193d, 32'h43ac063c, 32'h4382e79f},
  {32'h442aaa86, 32'h43952907, 32'h43a3a603},
  {32'hc5061011, 32'h43a2a97d, 32'hc31f135e},
  {32'h4399baf0, 32'h43a2779e, 32'hc3bfc957},
  {32'hc300aed8, 32'h40a43581, 32'hc18d42ae},
  {32'h44e6de40, 32'hc20683a2, 32'hc2c09861},
  {32'hc4bb8f94, 32'hc2d08f56, 32'h42320db9},
  {32'h43ee8995, 32'hc36e4825, 32'hc34d7a67},
  {32'hc49ee7e1, 32'hc3461ca5, 32'h43c019ce},
  {32'h439402ec, 32'h42a8f731, 32'hc340cec5},
  {32'hc46394b3, 32'hc3218300, 32'h429d9eb1},
  {32'h44a8fbdd, 32'h42c0f0b4, 32'hc3ad29ae},
  {32'hc30eca60, 32'h43b578f0, 32'h4384ddfe},
  {32'h44518a0e, 32'h4252ad27, 32'h431099c1},
  {32'hc46e61ce, 32'hc1b4859f, 32'h42b4cbea},
  {32'h44b34423, 32'hc350bc20, 32'h42d00484},
  {32'h43e5cac0, 32'hc349faa2, 32'hc30ae014},
  {32'hc508937a, 32'hc33ea3a1, 32'hc142bc69},
  {32'h445ea80b, 32'hc3ab0a00, 32'h43da6516},
  {32'hc4ac31e3, 32'hc3de64b3, 32'h4283bf41},
  {32'h44917087, 32'h43808b4f, 32'hc2e81b80},
  {32'hc3b8a5b2, 32'hc35790b5, 32'h43393909},
  {32'h447bf541, 32'hc3665773, 32'h4287435c},
  {32'hc4078f9c, 32'hc38075e7, 32'h432d2a5b},
  {32'h443dc6f4, 32'hc3cb74a2, 32'hc1144d76},
  {32'hc3174c44, 32'h43feddde, 32'h43bc5bd0},
  {32'h44ebe158, 32'hc2049f4b, 32'h4177f446},
  {32'hc503c1c6, 32'h4288d684, 32'h428eb858},
  {32'h44355f7c, 32'h42f10192, 32'hc3a45354},
  {32'hc496aeca, 32'hc305759f, 32'h42f54e9a},
  {32'h4438ca70, 32'hc345459b, 32'hc20e72c2},
  {32'hc4d804b0, 32'h429ef9e5, 32'h43297f26},
  {32'h43cf3209, 32'h43688bb7, 32'hc3c89ff6},
  {32'hc49b3cd1, 32'h410efc15, 32'h42e523c3},
  {32'h4489b6f9, 32'h42a49b89, 32'hc3848f1c},
  {32'hc48d522e, 32'hc24b1c0a, 32'hc38653ac},
  {32'h44832110, 32'h427c4860, 32'hc35c9b4b},
  {32'hc45c6a8a, 32'h42ada25e, 32'h4248c082},
  {32'h435b9ec8, 32'hc3b73d4e, 32'hc1e93db9},
  {32'hc291d3a0, 32'h429442ff, 32'h42a8e7f1},
  {32'h44e5acbc, 32'hc2ee8546, 32'hc31a6815},
  {32'h42055f0e, 32'h439e983e, 32'hc335c657},
  {32'h4515f788, 32'hc23e4cf1, 32'h43a0737a},
  {32'hc4e3c1e4, 32'hc3f49b1c, 32'hc2fed218},
  {32'h4335e054, 32'hc384e6f4, 32'hc35a2b7a},
  {32'hc3f9a020, 32'h42b94ae3, 32'h40ec6b60},
  {32'h44ec7338, 32'h41559370, 32'hc373d763},
  {32'hc43da48a, 32'h4260b086, 32'hc1bd47c3},
  {32'h44e48d0c, 32'h43f15219, 32'h42e5ce95},
  {32'hc44d9708, 32'h43b66eb2, 32'h428cf457},
  {32'h44527447, 32'h4302a354, 32'hc4099f21},
  {32'hc4a98a63, 32'h42b47dba, 32'h42baa742},
  {32'h4387d7e4, 32'h43090937, 32'hc2e7ab2e},
  {32'hc4b862ea, 32'hc3ce857e, 32'hc30ed450},
  {32'h44c32d6b, 32'hc29e7018, 32'h4220402f},
  {32'hc32fe899, 32'h4035e12b, 32'hc3b2fe53},
  {32'h43c8abf6, 32'hc3bb3d7f, 32'h43b680af},
  {32'hc4c6de05, 32'h432d39d7, 32'hc1cd24c4},
  {32'h440aad14, 32'h420aacdf, 32'h43903b07},
  {32'hc37dbce0, 32'hc37aa914, 32'h42750e39},
  {32'h434c56d8, 32'hc35129a1, 32'h42455bc9},
  {32'hc2078940, 32'hc34ee68a, 32'hc3314a2b},
  {32'h449314e1, 32'hc000f7a4, 32'h43614949},
  {32'hc2f0e320, 32'h43836ef4, 32'h43896b30},
  {32'h43bd38f5, 32'h44237888, 32'hc3b621e4},
  {32'hc402344b, 32'hc1e5f5bb, 32'h4302adcd},
  {32'h44c3f5c1, 32'h4305118f, 32'hc3063f4d},
  {32'hc4db00f5, 32'hc2a06288, 32'h43243cdd},
  {32'h43f5b980, 32'h4229275d, 32'h42c1917c},
  {32'hc43f3181, 32'hc326fa85, 32'h439ef023},
  {32'h4433a39f, 32'h40ff6d3e, 32'h41f7a841},
  {32'hc477e0fc, 32'hc1fd9531, 32'hc3348086},
  {32'h44d4b385, 32'h42251970, 32'hc399fa4c},
  {32'hc4b295ed, 32'hc21db45b, 32'hc337088f},
  {32'h45090cbd, 32'h42f17ee9, 32'h4402b63c},
  {32'hc470875b, 32'hc31ff0ea, 32'hc2cd7ac7},
  {32'h4494bf81, 32'hc37a7191, 32'h4352bdf5},
  {32'hc3ff4966, 32'h429bfd9d, 32'h4224dab5},
  {32'h44df9c38, 32'hc36f5106, 32'h42338407},
  {32'hc420e270, 32'h43745fae, 32'hc36d4388},
  {32'h44e5ffb9, 32'hc2230052, 32'h41e26346},
  {32'hc50cbb4f, 32'h43eb483c, 32'hc3b04346},
  {32'h449d83d6, 32'h436a7de5, 32'hc34cb1b8},
  {32'hc4819a09, 32'hc28ce711, 32'hc4139c9a},
  {32'h44b37084, 32'hc0e92807, 32'h43410514},
  {32'hc401bb0d, 32'hc0e3e134, 32'h43b50c0e},
  {32'h4500e318, 32'h42a35187, 32'hc2fe9076},
  {32'hc504f73c, 32'hc370bac8, 32'hc32ff981},
  {32'h450372c4, 32'h43bc1cea, 32'hc2fef1fc},
  {32'hc4d36709, 32'h4336051a, 32'h4309bd6b},
  {32'h442ac004, 32'hc2f2bba1, 32'h4243fe56},
  {32'hc4a4227a, 32'h432f009b, 32'hc2fe4077},
  {32'h4502b357, 32'h421eafcc, 32'hc283270e},
  {32'hc28122e0, 32'h43243d15, 32'h431be52c},
  {32'h44b92f27, 32'h42fdc063, 32'h411a96b1},
  {32'hc51aef66, 32'hc36e0ccf, 32'hc3bd838f},
  {32'h43782d20, 32'h4308a21d, 32'h43171471},
  {32'hc4672229, 32'hc3bb5073, 32'h43774ffc},
  {32'h4464b7a2, 32'hc1dbfe55, 32'h43c8d8d7},
  {32'hc413cac4, 32'hc3dd7302, 32'h42b8889c},
  {32'h44931f5c, 32'h4380e208, 32'hc347cb34},
  {32'hc43a4af4, 32'h420b6903, 32'h437c1d5d},
  {32'h43b74860, 32'h43d0332d, 32'hbf976d32},
  {32'hc44ef2c0, 32'h431cf33e, 32'hc39b6596},
  {32'h44eadf12, 32'hc2883fd0, 32'hc39007d2},
  {32'hc4e1a0e3, 32'hc3acf427, 32'hc376ab21},
  {32'h43bd8a34, 32'h430e6855, 32'hc3069034},
  {32'hc4e9198d, 32'h43563b0c, 32'h44395ae3},
  {32'h451ac51e, 32'h42f322fc, 32'h41ac4574},
  {32'hc5154d4f, 32'hc2876994, 32'hc3e69d15},
  {32'h4397874c, 32'hc30cb2f0, 32'h431707a2},
  {32'hc4926daa, 32'hc0f2e41a, 32'h429e4144},
  {32'h4478af00, 32'h4188107c, 32'hc298f726},
  {32'hc4ab63d6, 32'h4323e8ad, 32'hc29d03d9},
  {32'h43d4258c, 32'hc3606112, 32'h433c70ca},
  {32'hc507b601, 32'h426c5420, 32'h4390a5b9},
  {32'h442e477a, 32'h42b278de, 32'hc3861726},
  {32'hc435f2cc, 32'h43b4c792, 32'h42f1d947},
  {32'h450e4660, 32'hc347af0a, 32'h4276d8c0},
  {32'hc49d2d20, 32'h439822cd, 32'h42e88743},
  {32'h4330ede6, 32'hc3bea94b, 32'h434dde53},
  {32'hc4ff8489, 32'h42e6ec71, 32'hc3192f77},
  {32'h44308d2b, 32'hc20b6c4c, 32'h425899d1},
  {32'hc5058ba2, 32'h425a201c, 32'hc3373455},
  {32'h44bd5c8e, 32'h4229ac4d, 32'hc3940906},
  {32'hc4a09bd2, 32'hc2f3250f, 32'hc30b13fa},
  {32'h443f1ebc, 32'hc215f466, 32'hc314b989},
  {32'hc3f199c4, 32'hc328213d, 32'hc352df6d},
  {32'h4483f9aa, 32'hc39eed73, 32'hc330a129},
  {32'hc3ef86bf, 32'h4249144b, 32'h438f0c2a},
  {32'h4340ff50, 32'h42ccdc91, 32'h42b7b7ae},
  {32'hc4e943da, 32'hc2839328, 32'hc33163f8},
  {32'h450045cb, 32'h42840d96, 32'h40622e12},
  {32'hc37d6e23, 32'hc2f6955d, 32'h43b0329f},
  {32'h44ad379e, 32'h42d2b142, 32'h434c5adc},
  {32'hc505087b, 32'h4331f180, 32'h43e062a0},
  {32'h4254a470, 32'h43a54fe3, 32'hc41f4e8d},
  {32'hc50c08a0, 32'hc33a13ba, 32'h43ad3478},
  {32'h44de8b86, 32'hc27a18e7, 32'h43933b0a},
  {32'hc38588b4, 32'hc28e2e91, 32'hc2d34ad6},
  {32'h449fa2fa, 32'hc2c28e66, 32'hc3195c5f},
  {32'hc4430b6a, 32'hc3c43c13, 32'h42ae7b3c},
  {32'h44e41584, 32'hc3c61e9e, 32'h434b1e8d},
  {32'hc5028203, 32'h436ac72e, 32'h43c1a886},
  {32'h44c936a2, 32'h4387eb13, 32'h43773204},
  {32'hc4781be2, 32'h42dbf800, 32'hc28674ae},
  {32'hc2dfee6c, 32'h42be73f5, 32'h42ad968d},
  {32'hc51c2c24, 32'hc368eafd, 32'hc2105a50},
  {32'h44783148, 32'h427d6362, 32'hc34ca928},
  {32'hc38fa8ec, 32'h42a64692, 32'hc32165f5},
  {32'h450fe1fe, 32'h4306a9ec, 32'hc38fae93},
  {32'hc4d14df0, 32'h431a47de, 32'hc3aa1422},
  {32'h44cad4c9, 32'h41f78f39, 32'hc37583aa},
  {32'hc4d05b9d, 32'h4241bdc1, 32'h41d13af2},
  {32'h44a5fa5e, 32'hc27d92df, 32'hc380c5b8},
  {32'hc42b88da, 32'h422cd3a3, 32'hc2ddbcf5},
  {32'h44ac569b, 32'hc2d0e9b4, 32'hc313ee10},
  {32'hc4af030f, 32'h43c8f8c3, 32'hc3616245},
  {32'h441b205f, 32'h4384a648, 32'h436b59fe},
  {32'hc44dc8d8, 32'hc4307792, 32'hc38f7cfc},
  {32'h44ff20c8, 32'hc282649b, 32'h435e47e8},
  {32'hc46114a1, 32'h43a00547, 32'hc300cdf1},
  {32'h444d7291, 32'hc286b70b, 32'h438d2611},
  {32'hc4860924, 32'hc39ce74b, 32'h4335edcf},
  {32'h4414ba54, 32'hc3573793, 32'h431890d0},
  {32'h4163da00, 32'hc1b8cb9e, 32'hc33164a8},
  {32'h435005c8, 32'h42152d96, 32'h423c3970},
  {32'hc398d2a6, 32'h4341e6ec, 32'h432afdc9},
  {32'h44d45ee5, 32'hc206fca3, 32'hbfa1dfcf},
  {32'hc421c074, 32'h435f9249, 32'h412ba236},
  {32'h45021fc3, 32'h435506ea, 32'hc370c020},
  {32'hc4f7ac3e, 32'h42f86be8, 32'h437e6ce6},
  {32'h442cf4fe, 32'h421acb37, 32'hc2852106},
  {32'h41ba4e80, 32'h421c19ca, 32'hc2b0b9e2},
  {32'h45069314, 32'hc3c5007c, 32'hc338ca12},
  {32'hc31ed890, 32'hc33d8233, 32'h43ac19e8},
  {32'h44379efe, 32'h41d2f52c, 32'h43790f7e},
  {32'hc4e1045b, 32'h429506fe, 32'hc1462204},
  {32'h44ef1ab2, 32'h41cc2287, 32'hc302d49b},
  {32'hc506aaf9, 32'hc08381c0, 32'h4370e1eb},
  {32'h43ec89c4, 32'h420fc058, 32'hc363cad0},
  {32'hc4f4a1a0, 32'hc286b850, 32'hc18ac1c3},
  {32'h4416194b, 32'hc32de870, 32'h42a06404},
  {32'hc4e3e6aa, 32'h431fb6bf, 32'hc2d34f6d},
  {32'h44e94753, 32'h436b0846, 32'h4248e1b0},
  {32'hc340b06c, 32'h43b8dbb2, 32'hc2a318cf},
  {32'h44a2d554, 32'h43281fb1, 32'h42ba7267},
  {32'hc4e74d37, 32'h4376c23a, 32'hc2c584e6},
  {32'h44e3063b, 32'hc3071f76, 32'h4306f2ab},
  {32'hc5063498, 32'h42131af4, 32'hc1cbb00c},
  {32'h421ed080, 32'h4182e582, 32'h42b20230},
  {32'hc3d241d2, 32'hc3077c23, 32'hc3273e3f},
  {32'hc31ec6bc, 32'h42bc7e34, 32'hc08f6c19},
  {32'hc40c29d4, 32'h434e6ae3, 32'hc339f465},
  {32'h44ef76c5, 32'hc3516f07, 32'hc06b1440},
  {32'hc4a13ea9, 32'h434f5754, 32'hc3901f32},
  {32'h44dc83ac, 32'hc3f62eac, 32'hc39b173c},
  {32'h43259fb0, 32'h4348aee1, 32'hc09876f8},
  {32'h44de475b, 32'h4173efc6, 32'h43a818ad},
  {32'hc450cac5, 32'h432e3344, 32'hc3a35006},
  {32'h44c658ce, 32'hc3801079, 32'h43696ed6},
  {32'hc4f0c13f, 32'h434c9a05, 32'h42d0cad4},
  {32'h432429c4, 32'hc2b7b4d4, 32'hc2d8d46d},
  {32'hc49574ca, 32'hc23ead13, 32'hc2d7a7b4},
  {32'h43f93b22, 32'h42f3c62a, 32'h43b43c21},
  {32'hc32ae4c0, 32'h434c5bda, 32'hc3109405},
  {32'h4506b803, 32'h41564269, 32'h431b0262},
  {32'hc410781a, 32'hc1cb8d04, 32'hc1c20a0d},
  {32'h44b647bc, 32'h435ed85a, 32'h42c33d01},
  {32'hc4cbb1e4, 32'hc3bb7aef, 32'h42b379d7},
  {32'h44b401ed, 32'h43016ad5, 32'h42ad8b8d},
  {32'h431d2860, 32'h40442318, 32'h433e6279},
  {32'h44ddced4, 32'h4338b4c3, 32'h43077ba9},
  {32'hc4c9a289, 32'hc30703f2, 32'h41789d6a},
  {32'h448a81c8, 32'h4011c3a8, 32'h4317541a},
  {32'hc4a4f838, 32'h431b26ee, 32'hc22f5725},
  {32'h4496a64d, 32'hc1920784, 32'h420864e0},
  {32'hc48e626e, 32'hc129a065, 32'h4387df17},
  {32'h44bc3d04, 32'h4321d669, 32'hc307697b},
  {32'hc503fe94, 32'hc2dafa69, 32'h42ed20e2},
  {32'h440a6c5c, 32'hc3010290, 32'h434f0234},
  {32'hc4ace986, 32'h439281d5, 32'h43524d17},
  {32'h44625b67, 32'hc443d4b3, 32'h438333b3},
  {32'hc51b1f1d, 32'h43bfc4dc, 32'hc360bcdc},
  {32'h448d45c1, 32'hc3b353bb, 32'hc2db648d},
  {32'hc2c1d680, 32'hc388cb54, 32'hc3269a20},
  {32'h44f0c63f, 32'hc3ee82a6, 32'hc2a0f7e7},
  {32'hc4b4d3f2, 32'h43161783, 32'hc2b90926},
  {32'h448b3640, 32'h4331694e, 32'h42105dee},
  {32'hc500931d, 32'hc3341255, 32'h42ff3737},
  {32'h448fccf6, 32'hc32ee637, 32'hc24cc246},
  {32'hc2ac3c18, 32'h43566a35, 32'h436c4b8f},
  {32'h447ddd99, 32'hc34e2072, 32'hc23089bb},
  {32'hc4124673, 32'h43ee8601, 32'hc314ca09},
  {32'h436d4fa4, 32'hc295d959, 32'h3fe7bc1c},
  {32'hc4237c63, 32'h41b4b169, 32'h431c862a},
  {32'h44bc3b10, 32'h412a0ca8, 32'hc31943c6},
  {32'hc49cf139, 32'hc311cc95, 32'hc2b632d8},
  {32'h43e586d4, 32'hc390ee09, 32'hc3241056},
  {32'hc478b981, 32'h42fcd65b, 32'h4340e636},
  {32'h44943735, 32'h42be9aeb, 32'hc418413f},
  {32'hc42be080, 32'h43023379, 32'h43f46dcf},
  {32'h44654f4e, 32'h430f60a9, 32'h43200f55},
  {32'hc499abf6, 32'hc2f5a33d, 32'hc3c41e64},
  {32'h44d281cd, 32'hc3117379, 32'hc3289ec1},
  {32'h42f1fee0, 32'h413b644a, 32'h431964f0},
  {32'h44b9c88a, 32'hc2c0d95a, 32'hc1a007d4},
  {32'hc4d3ff22, 32'hc2fecb14, 32'h43b0b539},
  {32'h44ae7158, 32'hc34b098e, 32'hc3bfa72b},
  {32'hc4cbacce, 32'h41079664, 32'hc2fdee82},
  {32'h44bccca4, 32'h4337029d, 32'h4289f346},
  {32'hc4cacde6, 32'hc2c63a2a, 32'hc311ad8e},
  {32'h44162ee9, 32'hc1d9f7b9, 32'h435cdcca},
  {32'hc4d6ef7d, 32'hc35f67ff, 32'hc3d02c00},
  {32'h43d1fb7e, 32'hc317f888, 32'h4303f216},
  {32'hc45a72bc, 32'h42c7d1b9, 32'h42ad4883},
  {32'h44fe92c5, 32'hc3873044, 32'hc3ef1738},
  {32'hc490e088, 32'h4187c5a8, 32'hc3d16efa},
  {32'h45114708, 32'h432e09ac, 32'hc2f69431},
  {32'hc4f07533, 32'hc27b1412, 32'h4303cb6a},
  {32'h450bd637, 32'hc270c248, 32'h416b7232},
  {32'hc5154384, 32'hc3923be7, 32'h433ce6bb},
  {32'h44d757ad, 32'hc3fd1b29, 32'hc2664b3d},
  {32'hc45ff80d, 32'hc3677025, 32'hc2a35d0e},
  {32'h4506d762, 32'h42941bc1, 32'hc3636f5b},
  {32'hc5003fe7, 32'hc31dc870, 32'hc2568386},
  {32'h44fdfb6a, 32'hc28f364f, 32'hc143c93a},
  {32'hc4969ee1, 32'hc32ab00d, 32'hc1ffaa20},
  {32'h44b4c5b0, 32'hc296aaa0, 32'hc3c58578},
  {32'hc48388a4, 32'h438b739d, 32'hc2968612},
  {32'h440d5816, 32'h41a66de9, 32'h43130c79},
  {32'hc48e81ae, 32'h432e65c4, 32'hc3216e57},
  {32'h44b7ef50, 32'hc389b884, 32'h42936dad},
  {32'hc4a71e85, 32'h41dc6060, 32'h433d5400},
  {32'h4486c29d, 32'hc2bc17a3, 32'hc3214a0d},
  {32'hc4eef1dc, 32'hc250d8b5, 32'hc29beffd},
  {32'h44a04762, 32'hc2dbe71c, 32'hc31f2f1b},
  {32'hc4b4b26a, 32'h420c6ec4, 32'h43391383},
  {32'h441b54ae, 32'h43439100, 32'hc2f3c02b},
  {32'hc3c7fda6, 32'h4282f311, 32'h425badfe},
  {32'h44b87fa6, 32'h435ac585, 32'hc248a5df},
  {32'hc4c1924a, 32'hc31fb8a8, 32'hc1b2de28},
  {32'h450d3870, 32'h43060c27, 32'h4376bbc5},
  {32'hc4eaa9a1, 32'h4321cc62, 32'h42178897},
  {32'h445559ee, 32'h43d16c0d, 32'hc37ec4e7},
  {32'hc47ebc4c, 32'hc2591c5c, 32'hc361c926},
  {32'h450e76b7, 32'h428923fa, 32'h40d96a62},
  {32'hc4872602, 32'hc2b1e62f, 32'h42a8dc7e},
  {32'h44ee3be0, 32'h422ee903, 32'hc32a9326},
  {32'hc441cf23, 32'h432a978f, 32'hc2d08f42},
  {32'h451cb7db, 32'h42916157, 32'h426b3085},
  {32'hc41b1819, 32'hc224b6bc, 32'hc2bf2143},
  {32'h43c9c378, 32'hc3a0cf33, 32'hc35c9768},
  {32'hc48b45ae, 32'h431ca69a, 32'h428c1f97},
  {32'h44c9da7b, 32'hc3284db5, 32'hc2630e87},
  {32'hc3968fdd, 32'h41d74ba5, 32'h42b247b9},
  {32'h44be2ccf, 32'h4221c0d6, 32'h4292d1c7},
  {32'hc505a834, 32'hc3420f2d, 32'hc39ec03d},
  {32'h44c10b69, 32'hc1f29a0e, 32'hc2d4ed2b},
  {32'hc4ed5274, 32'hc380a7d8, 32'hc3996115},
  {32'h44454176, 32'hc211d1d5, 32'h427da476},
  {32'h429c4db3, 32'hc21f9406, 32'h4218d5e8},
  {32'h43dfb6c8, 32'h424ecbc8, 32'hc314c1e4},
  {32'hc4d981e5, 32'h43050441, 32'hc2a397be},
  {32'hc2c74260, 32'hc33e7ce3, 32'h4349dfd9},
  {32'h4295b9c0, 32'h43994b87, 32'hc351305b},
  {32'h448fcff5, 32'hc345f44b, 32'hc2488293},
  {32'hc434212c, 32'h433671d1, 32'hc3c11d17},
  {32'h44d7b030, 32'hc2d5f673, 32'hc1b934d5},
  {32'hc47d7869, 32'hc22dfd06, 32'h3f0aec54},
  {32'h442e3dc4, 32'hc355e7a7, 32'hc264b946},
  {32'hc51d44a1, 32'h41e02c88, 32'hc3007495},
  {32'h4421a89a, 32'h4339d956, 32'h40452bd2},
  {32'hc495eef0, 32'h435ce010, 32'h432ff5ca},
  {32'h4506a489, 32'h43ad8d46, 32'h43f5b70f},
  {32'hc4134e5e, 32'h43620d89, 32'h4310db3c},
  {32'h4490c18e, 32'h43393ddd, 32'hc28a5c38},
  {32'hc448fb94, 32'hc3811ba0, 32'h43843bc3},
  {32'h4499ce30, 32'hc323409f, 32'hc2ee13fb},
  {32'h43386c30, 32'hc3f34969, 32'h4360b660},
  {32'h44f00d05, 32'hc358e46a, 32'hc2f0203a},
  {32'hc455be4a, 32'hc2ec58e4, 32'hc20c0ce5},
  {32'h43830be3, 32'hc34433b7, 32'hc3ca0ab2},
  {32'hc4a08df7, 32'hc3c34f5c, 32'hc06abfe9},
  {32'h44576c19, 32'hc320514e, 32'h41b5c38a},
  {32'hc4bbd263, 32'h43fc2df1, 32'hc34466f8},
  {32'h44bc286d, 32'h43b3cf7d, 32'hc2b4169b},
  {32'hc2e4a9ac, 32'hc36a243d, 32'h4343fe1f},
  {32'h44106d56, 32'hc2bc5487, 32'hc1d63c13},
  {32'hc4c8a8df, 32'h43c4af09, 32'hc366e296},
  {32'hc15eae80, 32'h420e1adc, 32'hc3083187},
  {32'hc4c367d7, 32'h4239539c, 32'hc389f57a},
  {32'h44f77b2c, 32'hc31ab0cc, 32'hc26d40c1},
  {32'hc50aab24, 32'hc3b81066, 32'h43607d37},
  {32'h44ce9d5e, 32'hc3423017, 32'h4283661e},
  {32'hc49bd407, 32'h417751db, 32'hc3d71635},
  {32'h440d4abc, 32'h439bd7a5, 32'hc26b1eb8},
  {32'hc411dd28, 32'h42fdd0fe, 32'h42adab83},
  {32'h430826de, 32'hc38ed15f, 32'hc2171a65},
  {32'hc49f59ce, 32'hc23fe63e, 32'h43d4bd4a},
  {32'h446a08fe, 32'hc3a062d6, 32'h4347c879},
  {32'h42056cd4, 32'hc33fc811, 32'h439c0a86},
  {32'h44825275, 32'h4294ff45, 32'h42bd2f91},
  {32'hc3b28257, 32'h43255e48, 32'h437bbab2},
  {32'h44d20c1d, 32'hc415db20, 32'hc1288138},
  {32'hc482dcd7, 32'h43cd16c7, 32'h42c4de7c},
  {32'h450442ae, 32'h43f2ab40, 32'h434cb284},
  {32'hc424785e, 32'h42da62c7, 32'hc268b30e},
  {32'h44688640, 32'hc38d21da, 32'hc3a447d7},
  {32'hc4c9845c, 32'h4382a546, 32'hc3ff0674},
  {32'h450d4e2f, 32'h42ee3cd1, 32'h420ae764},
  {32'hc4e42834, 32'h432aea78, 32'h42f46806},
  {32'h451297b8, 32'hc2c514c3, 32'hc36266c2},
  {32'hc4a94c15, 32'hc37cb494, 32'hc3c4e2fd},
  {32'h44ff37f9, 32'hc3c76786, 32'hc35fe20f},
  {32'hc514c9c7, 32'hc196a582, 32'hc1f6f4b0},
  {32'h4526175c, 32'h4399b0a7, 32'hc2bc926c},
  {32'hc5142b73, 32'h438cf990, 32'hc37bb111},
  {32'h434ad1f2, 32'h4316bc1d, 32'hc25876d4},
  {32'hc4fbce9a, 32'hc255af08, 32'h4360fe63},
  {32'h44a60d5e, 32'h43b50cdc, 32'hc31b001b},
  {32'hc51903e8, 32'h416a9f07, 32'h43187e18},
  {32'h44427bf6, 32'hc387f8ea, 32'h41cf9e81},
  {32'hc506c320, 32'hc2dc390c, 32'h412e57a7},
  {32'h436f6334, 32'h43b2f3e5, 32'hc38647da},
  {32'hc4a1ee82, 32'hc30ecdf8, 32'h4326a82a},
  {32'h4403eb18, 32'hc275873d, 32'hc22fce1e},
  {32'hc4939c8f, 32'h3f19dcd3, 32'h4347a007},
  {32'h4510fd72, 32'h435e9781, 32'hc2908f5c},
  {32'hc4b52e22, 32'h42e5c320, 32'hc3862de4},
  {32'h44a5b11b, 32'h43435996, 32'h41939019},
  {32'hc468d8c3, 32'h430a5ecc, 32'hc306c25d},
  {32'h44334f70, 32'h438ff3de, 32'hc356d066},
  {32'hc494ec9e, 32'h42bf5e4b, 32'hc33da806},
  {32'h44aa025e, 32'h42802496, 32'h43435b07},
  {32'hc330ef6b, 32'hc389646c, 32'h42277f3e},
  {32'h4491bafc, 32'hc2527cfa, 32'h43409b0d},
  {32'hc482300e, 32'h435cecd5, 32'hc300edc1},
  {32'h44b130c3, 32'hc3d48482, 32'h42388f45},
  {32'hc4e23f32, 32'h43bf5015, 32'hc1930796},
  {32'h4444d55f, 32'h43266fc2, 32'hc2739afc},
  {32'hc46f813e, 32'h43c4c632, 32'hc3543900},
  {32'h4428accc, 32'h42bba273, 32'hc354604c},
  {32'hc484c3e4, 32'h435d6847, 32'hc3dfc669},
  {32'h450a301e, 32'hc3a69330, 32'hc353d17e},
  {32'hc5129e10, 32'hc32098e7, 32'hc3521ce8},
  {32'h43cf671f, 32'h42eaeb2d, 32'h438c0c5e},
  {32'hc1f5fde8, 32'hc2dd9def, 32'hc324afd1},
  {32'h44906abf, 32'hc2e36359, 32'hc21d0b19},
  {32'hc2fb33c0, 32'h42f510e4, 32'h439e4487},
  {32'h4432f6f6, 32'h435d5f53, 32'h42be4970},
  {32'hc4788408, 32'h420ebd0e, 32'hc29ca18a},
  {32'h42396990, 32'h4371c566, 32'h43ca7bf5},
  {32'hc4c7d240, 32'h430e9627, 32'hc3876b20},
  {32'h44f3ec34, 32'h440a9e61, 32'h434f6417},
  {32'hc41b6002, 32'hc244b5e1, 32'h439cd1b4},
  {32'h44e1d94f, 32'h44090698, 32'h432a547e},
  {32'hc2c68e7a, 32'h4306ffb4, 32'hc27b4f84},
  {32'h449de656, 32'hc3627abe, 32'h420e5900},
  {32'hc4ea2b0a, 32'h42acd5d1, 32'h4240e426},
  {32'h4483d1c5, 32'h42e23543, 32'hc2d28570},
  {32'hc440b088, 32'h43909394, 32'hc344e067},
  {32'h44b8f00d, 32'hc1c405ee, 32'h42f2d695},
  {32'hc4d8f976, 32'hc2fe2e8f, 32'h42ac5abd},
  {32'h4524faae, 32'h42b75daa, 32'hc283679a},
  {32'hc46e3c5e, 32'h43a292fa, 32'hc30e9cf2},
  {32'h450daa83, 32'hc22463e2, 32'hc2d16938},
  {32'hc38da418, 32'hc0734c40, 32'h43a31dc3},
  {32'h449fdf7e, 32'h437d0674, 32'hc3a5a21a},
  {32'hc513677f, 32'hc30d0cd0, 32'hc1c6a945},
  {32'h44d0a34b, 32'h425225de, 32'h43dbd6d3},
  {32'hc46ff0bd, 32'h4299eb81, 32'h418bb66c},
  {32'h4507b1d1, 32'h42d987ad, 32'h42ab5e85},
  {32'hc51072ee, 32'h430ab236, 32'h436afed3},
  {32'h44925097, 32'hc3904f53, 32'h43adbf18},
  {32'hc4f5dcd4, 32'h4249aeec, 32'h42597a30},
  {32'h4419cd58, 32'h41d306b6, 32'h4358ef5b},
  {32'hc4c4ba51, 32'h44194497, 32'h426e3994},
  {32'h44bf38fa, 32'h43fde2a9, 32'hc39fc067},
  {32'hc3063945, 32'h41b3e397, 32'h433536f8},
  {32'h44b61681, 32'hc14cdcd6, 32'hc3ba4903},
  {32'hc503f712, 32'h437b478e, 32'hc2d1db50},
  {32'h44341974, 32'h439478e7, 32'h421e2e60},
  {32'hc49d8e42, 32'hbf4c9980, 32'hc36a9fb8},
  {32'h44fa7752, 32'hc20559a2, 32'h43c098b4},
  {32'hc5041fe9, 32'h43acb0c3, 32'h4281b94a},
  {32'h44aa22bd, 32'hc2df6af5, 32'h43b1768a},
  {32'h431d1df0, 32'h43f2af1b, 32'hc2bfc5dc},
  {32'h44c12f4a, 32'hc2f055da, 32'h4218f82c},
  {32'hc4e0f0ba, 32'h4018fabe, 32'hc36ca838},
  {32'h45077267, 32'hc21ff97c, 32'hc329a246},
  {32'hc4c83748, 32'hc27672ef, 32'hc301d75e},
  {32'h44244c84, 32'h431147b8, 32'h43890681},
  {32'hc4d4d005, 32'h43183f4d, 32'h433d64ce},
  {32'h432b561c, 32'h4395ee6d, 32'hc327e8c5},
  {32'hc4199f4e, 32'h43dbfc6a, 32'h429b5893},
  {32'h442f381f, 32'hc2b07b77, 32'hc3aed9fa},
  {32'hc4a7c2ba, 32'h43c19b0e, 32'h4362a073},
  {32'h44f3e192, 32'hc2d5ff09, 32'h4301de8f},
  {32'h4275e2c0, 32'h42ee3d07, 32'hc370c2e3},
  {32'h428f62b4, 32'hc36fb164, 32'h43bbf34f},
  {32'hc4d3f26c, 32'h429be07c, 32'hc264c19b},
  {32'h446fadea, 32'h43c06030, 32'hc1cf4ab9},
  {32'hc4d19157, 32'h42fd8302, 32'hc19a83c8},
  {32'h44b94930, 32'hc3a44b50, 32'hc2be4d2c},
  {32'hc4027b6d, 32'h42ae1ebe, 32'h42463d87},
  {32'h44991f38, 32'h439dd767, 32'h42d6cda9},
  {32'hc496f970, 32'h4172e1fa, 32'hc2576f13},
  {32'hc4a7b9c9, 32'h438eab34, 32'h431ec22e},
  {32'h44d4bd44, 32'h42874e91, 32'h4204daab},
  {32'hc2d0c1ec, 32'h4308037a, 32'h43cc2d54},
  {32'h43f0fb4e, 32'hc35b4364, 32'hc2bbdb58},
  {32'hc4b900db, 32'h43b7ce08, 32'hc2f1e6f1},
  {32'h4413baa8, 32'h43b51a71, 32'h43249126},
  {32'hc518de99, 32'h4356e8c1, 32'h430d4bde},
  {32'h44e32ef0, 32'hc2a0deae, 32'h43cb9793},
  {32'hc5016363, 32'h43031ce5, 32'h41ae89ee},
  {32'h447bd592, 32'hc2e6b009, 32'hc2ceff79},
  {32'hc4cefb71, 32'h435f20e9, 32'hc3b5caf8},
  {32'h44dbd578, 32'h42e4396f, 32'hc281c6ab},
  {32'hc46a4509, 32'h43925015, 32'hc2b09d52},
  {32'h443cecdc, 32'h42a5a90f, 32'h42d7a19a},
  {32'hc48f5ab4, 32'h4292e87a, 32'hc3a0a5ec},
  {32'h44aaf5fd, 32'hc31ff032, 32'h42d8b97e},
  {32'hc47d5571, 32'h429fcbda, 32'h428c77e0},
  {32'h45096fad, 32'hc2914e7e, 32'hc31442bd},
  {32'hc5073187, 32'hc33abec2, 32'hc148efdc},
  {32'h44d6242a, 32'hc2b7f024, 32'h43080d3f},
  {32'hc505b779, 32'h43b85a69, 32'hc3f246ea},
  {32'h444e88e4, 32'h42791731, 32'h42967903},
  {32'hc4cb59d6, 32'hc2cc38f7, 32'hc3db42ad},
  {32'h44e3ceb2, 32'hc2a3383f, 32'h42bf96c6},
  {32'hc3440258, 32'h428cd8f1, 32'hc3bbb07b},
  {32'h44c2bd81, 32'h435c77b6, 32'h4312cbb9},
  {32'hc4ade582, 32'h432220e8, 32'h4270603a},
  {32'h4414d0f4, 32'hc40a5ff3, 32'hc3c174e3},
  {32'hc4858c8e, 32'h423cd2aa, 32'hc3121f94},
  {32'h449e796a, 32'h42f1673d, 32'hc271ae88},
  {32'hc48828be, 32'hc32a29b5, 32'h42d515ce},
  {32'h4448c408, 32'h4332e716, 32'h4366e7a8},
  {32'hc4c71ad5, 32'hc318f1c7, 32'hc2d18368},
  {32'h43a491d4, 32'hc2bb3218, 32'h435a0fde},
  {32'hc346e2f1, 32'h431d58cc, 32'hc38ab4ff},
  {32'h44cd6afe, 32'h4386473f, 32'h41f4f190},
  {32'hc4f22c5e, 32'hc28eeb07, 32'hc38c1e84},
  {32'h44d1a1d9, 32'hc38c5fee, 32'h43f6c818},
  {32'hc3b79a26, 32'h43968718, 32'hc311f8d5},
  {32'h44dd54e7, 32'hc1d0eab3, 32'h41bb3c21},
  {32'hc485bc32, 32'h44079b45, 32'h42d282e9},
  {32'h44bb2c81, 32'h428c8c28, 32'hc3d2916e},
  {32'h431794c6, 32'h42248bb6, 32'hc2acb92d},
  {32'h442bc5ee, 32'h43239274, 32'h431c7217},
  {32'hc4a6f017, 32'hc2af990b, 32'h429e670a},
  {32'h44801baf, 32'hc2e2ef14, 32'h4326f74b},
  {32'hc44f4ba8, 32'hc2bc9fd0, 32'h4323865e},
  {32'h44e878b9, 32'hc2fdb5c1, 32'hc391c71a},
  {32'hc48500ea, 32'hc21e9c5c, 32'h42978a95},
  {32'h44e38fa1, 32'h41f5ea15, 32'hc3be16d7},
  {32'hc502b653, 32'hc3d9fc23, 32'h43940fcd},
  {32'hc312eba0, 32'h437d8b86, 32'hc0bec69b},
  {32'hc4f03a46, 32'h437381e0, 32'hc3765120},
  {32'h434df4dc, 32'hc30a26c2, 32'h4031bcc3},
  {32'hc4c9e108, 32'h432cce44, 32'hc311ffc4},
  {32'h44c60a12, 32'h432600c0, 32'hc30f5b99},
  {32'hc47b9464, 32'h43c20bad, 32'hc35f4c06},
  {32'h443e94c4, 32'h42b2ca42, 32'hc347ff1f},
  {32'hc48c90cb, 32'hc3311e97, 32'h42cf739c},
  {32'h4499bb0f, 32'h428aafad, 32'hc2e99ab4},
  {32'h4290da1c, 32'h43b2ee2a, 32'hc36d205d},
  {32'h4511c5a1, 32'h425d7b12, 32'hc390a6bc},
  {32'hc482a48d, 32'hc31e4eb5, 32'hc3225ca0},
  {32'h450a8117, 32'h425de617, 32'h43016fdc},
  {32'hc4e2a61d, 32'hc2fe2cdb, 32'hc33aaa61},
  {32'h44e97fb6, 32'h43a552c4, 32'h421b40a5},
  {32'hc512e0f4, 32'hc40193ce, 32'hc23f7e0a},
  {32'h44ba8f2c, 32'hc29e065c, 32'hc41158d1},
  {32'hc49c7aa8, 32'h43c38629, 32'hc392351a},
  {32'h448d9efe, 32'h42764db6, 32'h43a3e05d},
  {32'hc4d6d35e, 32'h42e8a1d9, 32'h4259c9fe},
  {32'h443add14, 32'hc2c12f22, 32'h43bbf52a},
  {32'hc448d7ba, 32'h4305af53, 32'hc2845cb5},
  {32'h43652fe4, 32'h432a9e6c, 32'hc1b639c1},
  {32'hc4e258f3, 32'hc36026a3, 32'h428384d1},
  {32'h44dcc6e1, 32'h435d49d0, 32'hc2e5e1be},
  {32'hc451e5fb, 32'hc364064a, 32'hc32972fa},
  {32'h4421ffb0, 32'h43fd5243, 32'hc200c241},
  {32'hc3e2a798, 32'hc19c5166, 32'hc22e92dd},
  {32'h44ac98b6, 32'hc33614b4, 32'h43f8f2a7},
  {32'hc4469d98, 32'hc3986f0d, 32'h4330f74e},
  {32'h4509dcf7, 32'hc3da6ca8, 32'hc326b8a4},
  {32'hc4f20f5c, 32'h43c0a6f9, 32'hc387d88b},
  {32'h4497d556, 32'h43a65698, 32'h42735c29},
  {32'hc47c8e56, 32'h43b6c096, 32'hc31cf8cd},
  {32'h443bf974, 32'hc29ff62c, 32'hc131c060},
  {32'hc3be8a5c, 32'hc23f75f4, 32'h42930da0},
  {32'h44cf0206, 32'hc27aa484, 32'hc325b37a},
  {32'hc52e784e, 32'hc30f6f12, 32'hc3eb3400},
  {32'h451c765a, 32'hc33d0773, 32'hc31ede77},
  {32'hc47054c1, 32'h431cc540, 32'hc31bc9d4},
  {32'h4413bcbd, 32'h42e586f3, 32'hc19c1746},
  {32'hc473cf2a, 32'hc3cb5d72, 32'hc301f866},
  {32'h4510999c, 32'hc01be490, 32'h43e22f49},
  {32'hc4fae038, 32'hc331f381, 32'hc3d38c36},
  {32'h44996d33, 32'hc38f4b94, 32'hc3103b4d},
  {32'hc47ed9d2, 32'hc1c9cc59, 32'h43a0a67d},
  {32'h44cf3158, 32'hc3236390, 32'hc2ed9c02},
  {32'hc4eaa0b8, 32'h43b2e2c7, 32'hc3bcee4a},
  {32'h450c4f8a, 32'h438402e9, 32'h422ca770},
  {32'hc437a432, 32'hc38cf339, 32'hc3144660},
  {32'h45074f46, 32'h430e4c67, 32'hc3146c11},
  {32'hc47fea99, 32'hc2e392a2, 32'hc3992524},
  {32'h43e93320, 32'h4325fb4f, 32'hc273a000},
  {32'hc50d9807, 32'h4355cff0, 32'h4329e683},
  {32'h445a85e6, 32'hc3c0dc38, 32'h42822b23},
  {32'hc49266e7, 32'h3f75fd2d, 32'hc3ea32e3},
  {32'h41d8e9a0, 32'hc42546c0, 32'h435c3ffc},
  {32'hc4f293d2, 32'hc2703266, 32'h43736a36},
  {32'h44d0b21c, 32'hc2c32874, 32'hc3d63c53},
  {32'hc4a62add, 32'h435aa9d0, 32'hc35b774c},
  {32'h44afe08a, 32'hc23f13f8, 32'h4345df4b},
  {32'hc4e206c7, 32'hc266bf86, 32'h428d6b77},
  {32'h44a71d7a, 32'h4331c237, 32'h41a50d73},
  {32'hc4087890, 32'h43ef5e0a, 32'h438d70e7},
  {32'h44fc641d, 32'hc3debc55, 32'hc42072a9},
  {32'hc4fc8674, 32'h42ad2634, 32'h4237a86b},
  {32'h4502dec7, 32'h42fa71c0, 32'h4380f86d},
  {32'hc50254a2, 32'hc3a1baf9, 32'h43bb2967},
  {32'h44497b74, 32'hc313a781, 32'h428fe186},
  {32'hc50098aa, 32'h436f56be, 32'h4327819b},
  {32'h44a8494e, 32'h42f14320, 32'h4332b628},
  {32'hc3cc5a31, 32'h42837b7f, 32'h433570de},
  {32'h44840412, 32'hc33c94e1, 32'hc2c3235f},
  {32'hc414ef15, 32'h418d686e, 32'h43220ecd},
  {32'h44735763, 32'hc2a6ed1d, 32'hc3340663},
  {32'hc4d460a7, 32'hc2809083, 32'h4305c60a},
  {32'h44c2d090, 32'hc26dda4d, 32'hc3488c2c},
  {32'hc4d21d8d, 32'hc35f7f60, 32'hc25f5671},
  {32'h4538a3d8, 32'h436728a9, 32'hc37a379d},
  {32'hc391ec55, 32'h4304596a, 32'h42c4c3b2},
  {32'h43a81dfb, 32'h43943bcf, 32'h4328af5e},
  {32'hc4af7124, 32'hc2967a44, 32'h4338653e},
  {32'h44f5cd37, 32'h43611bc8, 32'hc29659ed},
  {32'hc5079c08, 32'hc38755c0, 32'h43ecfc0f},
  {32'h4433d43e, 32'hc3894e35, 32'hc3c0b1fa},
  {32'hc4a2fcf2, 32'hc2539d7f, 32'hc3398f0a},
  {32'h43b09650, 32'h43810001, 32'hc2c14841},
  {32'hc50433a4, 32'hc28a3704, 32'h42c5e80a},
  {32'h44ec0335, 32'hc384d249, 32'h429366f5},
  {32'hc39542e8, 32'hc29f1ef2, 32'hc22718ba},
  {32'h44f9093e, 32'hc08e01be, 32'h428b5746},
  {32'hc4eef20a, 32'h431ce3fd, 32'h436c06e5},
  {32'h44b5fa0c, 32'h435cb75d, 32'h3ec9d9e0},
  {32'hc4b7e800, 32'hc2ad3b2e, 32'h4319c22a},
  {32'h44a26bab, 32'h41c6a75f, 32'hc3d647b7},
  {32'hc3f1c964, 32'h43c3989d, 32'h434c27ba},
  {32'h440161d0, 32'h43e9b908, 32'hc259297e},
  {32'hc500feeb, 32'h429bb161, 32'h4372aba2},
  {32'h43e4a538, 32'hc2ae9dd3, 32'h432a6cff},
  {32'hc4221b7a, 32'h434c37e3, 32'h437ed60b},
  {32'h45073d5e, 32'hc3696ab5, 32'hc34b9587},
  {32'hc50202be, 32'hc340f012, 32'hc242f9dc},
  {32'h44d64d80, 32'hc3231974, 32'h42b3506e},
  {32'hc3d45606, 32'h43befd8c, 32'h42ef5c75},
  {32'h449a45a3, 32'hc3ac4565, 32'hc32cd7e5},
  {32'hc50187e3, 32'hc37b9910, 32'hc26d3d18},
  {32'h4360ed20, 32'hc2379d54, 32'h433fb27e},
  {32'hc49a4e01, 32'hc259fe8b, 32'hc351bb22},
  {32'h449591c8, 32'hc351c434, 32'h42bd338f},
  {32'h42c087d0, 32'h41d4b223, 32'hc3fb9748},
  {32'h44b9577a, 32'h433d6850, 32'hc39ee113},
  {32'hc462abbe, 32'hc1cc093a, 32'hc1b099ff},
  {32'h4446404d, 32'h4295ab19, 32'h43016ca2},
  {32'hc4ae51d4, 32'h437b5df2, 32'hc384b520},
  {32'h446ea3c4, 32'hc3d7a767, 32'hc12f273a},
  {32'hc46016b7, 32'h43d37214, 32'h4306a5c7},
  {32'h449d39c6, 32'h41dfe3ae, 32'hc2e0d618},
  {32'hc3b96140, 32'hc316861c, 32'hc2241bf8},
  {32'h44f41729, 32'h437428dc, 32'hc23d0c64},
  {32'hc4cf3fd1, 32'hc208d77d, 32'hc1c4b8d8},
  {32'h439348a8, 32'h426d4086, 32'h4126ef6e},
  {32'hc47d7fbd, 32'h42492892, 32'h4335661c},
  {32'h441b3144, 32'hc342e142, 32'hc2e14082},
  {32'hc40332c4, 32'h4375d01f, 32'hc30fd329},
  {32'h42116d00, 32'hc30fff5c, 32'hc325a2e0},
  {32'hc4f64ebe, 32'h43a80e57, 32'h419a28e1},
  {32'h44aa4f33, 32'hc3822d5b, 32'hc33f2b39},
  {32'hc396b58b, 32'hc3cadd70, 32'hc371a01f},
  {32'h449b3467, 32'hc32e7cdf, 32'h431369c9},
  {32'hc460e594, 32'h42ab0dd5, 32'hc2f86cea},
  {32'h44bb19e3, 32'hc1f94e95, 32'h43a020c9},
  {32'hc4909ea0, 32'hc1b19c41, 32'h430f03dd},
  {32'h440801f6, 32'hc0ee57da, 32'h42984d94},
  {32'hc4ff214d, 32'hc33a9a95, 32'h43554c0e},
  {32'h44fa5b2e, 32'hc33cf4b0, 32'h437063f0},
  {32'hc50db737, 32'h42a211d0, 32'hc10d8c83},
  {32'h43c7a06a, 32'hc3b1614e, 32'h421a50c1},
  {32'hc44e1e00, 32'hc43488f4, 32'hc2e81178},
  {32'h44220204, 32'hc36579a3, 32'h42b5ef88},
  {32'hc411ceba, 32'h43af593e, 32'h43a92b01},
  {32'h4464ef33, 32'hc262c72d, 32'h4308a08b},
  {32'hc4864387, 32'hc2175282, 32'h43115ad2},
  {32'h44724cf0, 32'hc3c698ca, 32'h42a04f07},
  {32'hc31e1a20, 32'hc2161b38, 32'h4309399c},
  {32'h44ccf97b, 32'hc38a41b3, 32'hc2eb1b09},
  {32'hc4d2d23d, 32'hc136202e, 32'h41a0fcf1},
  {32'h44e21271, 32'h42a9edb1, 32'h439b8737},
  {32'hc49abaf3, 32'h4391d621, 32'h43c529c7},
  {32'h432b2538, 32'hc326c873, 32'h41bc2721},
  {32'hc50b1985, 32'hc1ccabdc, 32'h42fcbcb3},
  {32'h448ff607, 32'h438f3ebd, 32'hc24ce843},
  {32'h4331e893, 32'h43fe75ef, 32'h41a2720e},
  {32'h424e8040, 32'hc300e478, 32'hc36a638f},
  {32'hc3c31d98, 32'hc3201f6c, 32'h43ad2806},
  {32'h4479ecf8, 32'h432e89d6, 32'hc3df7019},
  {32'hc517833d, 32'h41c78f34, 32'hbe53d8bc},
  {32'h43ec3887, 32'h4130f4f4, 32'h4315a1b9},
  {32'hc3d0dc60, 32'hc2f3b8cd, 32'hc231bd45},
  {32'h44b41ae4, 32'h40e9f32c, 32'h4416848c},
  {32'hc3cc0092, 32'h4365a3aa, 32'hc2bad89a},
  {32'h445796f6, 32'hc33b253a, 32'h43f08a53},
  {32'hc406bb78, 32'h429dc5ff, 32'h41d66e36},
  {32'h438e8488, 32'hc2b0fa69, 32'h43b8ea00},
  {32'h4018c800, 32'h43d3c3f1, 32'h41c463fd},
  {32'h44c8b39b, 32'h4348db30, 32'hc21bf405},
  {32'hc485a5af, 32'h404abed8, 32'hc38ad124},
  {32'h441e92fa, 32'h423f6768, 32'hc39d4b43},
  {32'hc49eeab6, 32'hc38c8173, 32'hc0e58b5a},
  {32'h44e8e378, 32'h4218aa28, 32'hc2ba1308},
  {32'hc4bd13d8, 32'h41382852, 32'h438695d5},
  {32'h440eab6e, 32'h434c7375, 32'h439e0419},
  {32'hc3b3d876, 32'h439c2c8d, 32'h42c2cc94},
  {32'h45033b9e, 32'hc2cbc553, 32'h432de090},
  {32'hc1b58180, 32'hc353c8c5, 32'hc39ca4b7},
  {32'h44fba775, 32'h42a9f487, 32'hc3dfb9eb},
  {32'hc4f10b2a, 32'h42820f78, 32'hc33ad6ac},
  {32'h44a0d3f4, 32'hc340586f, 32'h43626cdd},
  {32'hc48e4354, 32'hc28b4996, 32'h435baae8},
  {32'h4461b330, 32'h436a5a01, 32'hc3b33110},
  {32'hc506e842, 32'h4223c004, 32'hc34fe659},
  {32'h4493c594, 32'hc26ce334, 32'h43211404},
  {32'hc4ef530a, 32'h43820fec, 32'h41cc170b},
  {32'h44dc3ffb, 32'hc22680f8, 32'hc2a73afe},
  {32'hc4bc42ff, 32'hc17322d3, 32'hc37ee646},
  {32'h44927a29, 32'hc407fa90, 32'h42c35ba6},
  {32'hc4aa0f84, 32'hc2c1d7e9, 32'hc26f2fe7},
  {32'h44ca4279, 32'hc2f57787, 32'h4281cd14},
  {32'hc3f2ec70, 32'hc31c56ee, 32'hc30a7ebb},
  {32'h44a5ad82, 32'hc26b21f1, 32'h4411d61b},
  {32'h410639d8, 32'h43d32374, 32'hc0eb7bab},
  {32'h44620315, 32'h427b361d, 32'hc2288a4d},
  {32'hc499f495, 32'h430c1268, 32'hc2cdfa47},
  {32'h4518af21, 32'h43560f2c, 32'hc3440c84},
  {32'hc4a3e11d, 32'h438694a3, 32'hc3275288},
  {32'h443732dc, 32'hc2d6df72, 32'h42c3bc9a},
  {32'hc4555444, 32'h4225b8ce, 32'h41152380},
  {32'h44a38a6f, 32'h439aa817, 32'hc3109339},
  {32'hc4121624, 32'h43c15bd9, 32'hc2e66e92},
  {32'h449a55f0, 32'h429f68e0, 32'h434dcdce},
  {32'hc4af8954, 32'hc2bf5609, 32'hc3829863},
  {32'h4471a61e, 32'hc3847909, 32'hc33b98aa},
  {32'hc4385b61, 32'hc45190e5, 32'h42e85624},
  {32'h451ec192, 32'h4290695b, 32'hc387f05f},
  {32'hc4bba8a1, 32'hc3ac3dbc, 32'hc1955b62},
  {32'h451ba1d3, 32'hc3993f4b, 32'h4355f5a2},
  {32'hc4f1fb4f, 32'hc11a3790, 32'hc3fc43e1},
  {32'h44ee15ac, 32'hc385d937, 32'h42c2294d},
  {32'hc3de0e22, 32'h43b9a04e, 32'h431af520},
  {32'h44576ae7, 32'h43a6a3c4, 32'h43ead925},
  {32'hc4b3f988, 32'h43154753, 32'h4323fbb4},
  {32'h449b1112, 32'h41193729, 32'hc39a9d02},
  {32'hc4b1aac4, 32'hc2bac6d1, 32'hc3bd79d4},
  {32'h4425f90c, 32'hc208b700, 32'h43a547cc},
  {32'hc48eab1c, 32'hc3b17207, 32'h439806f7},
  {32'h43aec128, 32'h4332a45e, 32'h4411ff7e},
  {32'hc4b5d369, 32'h43530848, 32'hc079ecc5},
  {32'h449f3efa, 32'hc3687edb, 32'hc2523e82},
  {32'hc48db848, 32'h42be15d6, 32'h42b6a1de},
  {32'h43b6c0ab, 32'h434a7e5b, 32'hc19ea636},
  {32'hc4cf9466, 32'h43bdea6e, 32'h43efb546},
  {32'hc2e67e2f, 32'h417a0a56, 32'h4318c5c5},
  {32'hc49ebd10, 32'hc349dfad, 32'hc2965c9c},
  {32'h451aba09, 32'hc2253b5e, 32'hc3dacc8e},
  {32'hc4daf01e, 32'h4306f4e4, 32'h43b691e8},
  {32'h44e184d8, 32'hc2fce8e6, 32'hc3d394d1},
  {32'hc4bf3dc3, 32'h42129362, 32'hc275a327},
  {32'h44d0a77f, 32'h42949c50, 32'hc39d957b},
  {32'hc401d296, 32'hc3a113c0, 32'h436670e9},
  {32'h43dc2a41, 32'hc17c9a06, 32'h427f05bf},
  {32'hc518483e, 32'hc3064a09, 32'hc3184d8d},
  {32'h444bb1e4, 32'hc3a40f90, 32'h42be99fe},
  {32'hc401f3f3, 32'h43996b76, 32'h42a4266f},
  {32'h44d171ec, 32'hc340231e, 32'hc2b0f70f},
  {32'hc4a1e141, 32'h4309e56e, 32'hc2b86022},
  {32'h44868211, 32'h4311eca5, 32'h4287c260},
  {32'hc4fa153d, 32'h429d1be7, 32'h421bac2f},
  {32'h4502ab31, 32'h416438dc, 32'hc35e06f7},
  {32'hc505d182, 32'h42d1fffa, 32'h420d43db},
  {32'h44d9d3b0, 32'h43636b0d, 32'h4287e87d},
  {32'hc40f205d, 32'h429a0dfb, 32'hc1d19ba2},
  {32'h44ba5b25, 32'h42cd6601, 32'h43aaa6bc},
  {32'hc4b96bd8, 32'h439f652c, 32'h42bc9c33},
  {32'h44bfcc87, 32'h438838c6, 32'hc213810d},
  {32'hc4693765, 32'h4082534c, 32'h430dfae1},
  {32'h4346bad2, 32'h42af0faa, 32'h4210d5bd},
  {32'hc4f03b90, 32'h4352868f, 32'hc326efd7},
  {32'h450543e7, 32'hc28cad16, 32'h4309d333},
  {32'hc45314e2, 32'hc1b61ca2, 32'hc2fe4996},
  {32'h449c7e4e, 32'h439ad01b, 32'h42b323d8},
  {32'hc42d2e76, 32'h43a681a8, 32'hc239f8bd},
  {32'h44142efc, 32'hc3332780, 32'hc34e228c},
  {32'hc36d88f9, 32'hc2a10233, 32'h42915cdd},
  {32'h45036c94, 32'h43678d4b, 32'hc3a90bd1},
  {32'hc4cf15da, 32'hc301bb26, 32'hc33869fe},
  {32'h44a6fa74, 32'hc2aed250, 32'hc32d89e2},
  {32'h43041274, 32'hc1c52dd1, 32'hc2d47c68},
  {32'h446ee878, 32'h43ee547d, 32'hc3551ad3},
  {32'h42fcf580, 32'hc2e1eb69, 32'h414c66f2},
  {32'h44cda5b3, 32'hc33de2a7, 32'h4346abb5},
  {32'hc419aeda, 32'hc38eb532, 32'h439a4728},
  {32'h4506a78d, 32'hc2ed7141, 32'h42d7c57d},
  {32'hc3fcc100, 32'h42ceddc0, 32'h43d40886},
  {32'h450452c2, 32'hc23fecbd, 32'h42d8d17c},
  {32'hc4d0becf, 32'h43c67cb8, 32'hc2e87b0f},
  {32'h44d88e01, 32'h42befa04, 32'h42b35fd0},
  {32'h430564ec, 32'h41ad3f10, 32'hc105c2c1},
  {32'h45062b3a, 32'hc3d05c2a, 32'h434a7cfe},
  {32'hc5028725, 32'hc2fce4cf, 32'hc2db0669},
  {32'h44c5e3fb, 32'hc37cc327, 32'hc30b85d1},
  {32'hc33e12e8, 32'h43ad2119, 32'hc3163181},
  {32'h44be0ce8, 32'hc2a52af1, 32'h42eb3caa},
  {32'hc4ccac39, 32'hc1567c64, 32'h4319d1d6},
  {32'h4457e42e, 32'hc3b5ac41, 32'hc3491afb},
  {32'hc49c328c, 32'h4014314b, 32'hc338008e},
  {32'h44d0f590, 32'h4288e300, 32'hc3d69b24},
  {32'hc489ec35, 32'h4301c54f, 32'hc19c9582},
  {32'h44b13822, 32'h42baa6cc, 32'h429f8812},
  {32'hc4984e1b, 32'hc2ee1dc1, 32'h43182abe},
  {32'h44f34206, 32'h4336aaf4, 32'h4346fdc8},
  {32'hc50d1f87, 32'hc2a6a93a, 32'h42c075a0},
  {32'h44cb0492, 32'h413e4007, 32'h4365a92c},
  {32'hc5216d3d, 32'h43055852, 32'h3fa63b8c},
  {32'h44054cb8, 32'h4228e702, 32'hc20c88ce},
  {32'hc4a7611f, 32'h41bd3564, 32'hc38517b5},
  {32'h449859f4, 32'h4383ea6d, 32'hc3bd9115},
  {32'hc51e38e8, 32'hc31592b1, 32'hc35f36b5},
  {32'h4424e528, 32'h434f1b9c, 32'hc3674fcd},
  {32'hc415d16c, 32'h433c9fcc, 32'hc2de1104},
  {32'h4411e7f1, 32'hc1aa91ee, 32'h42ea4293},
  {32'hc49dba42, 32'hc36dfbd5, 32'h4279cf87},
  {32'h45077ba7, 32'h433b0e6d, 32'hc398ff27},
  {32'hc4de2e85, 32'h42ba241e, 32'h43a88749},
  {32'h43b12e08, 32'hc2fa53a0, 32'h4390ea02},
  {32'hc52249eb, 32'h431b2eb4, 32'hc2956216},
  {32'h44898b09, 32'h43910de1, 32'hc3b72de5},
  {32'h40cce836, 32'hc29d55f5, 32'hc127483d},
  {32'h449eb35a, 32'h43782158, 32'hc27570e0},
  {32'hc519e2d3, 32'h4317b31b, 32'hc2d15722},
  {32'h44d231bb, 32'h435298b1, 32'hc3d6a5fc},
  {32'hc4d99ccd, 32'hc266cb5d, 32'h429db655},
  {32'h44f74f4b, 32'hc3139519, 32'hc3488edf},
  {32'hc4cffbbc, 32'h42d82944, 32'h43c0857b},
  {32'h44d2751b, 32'hc299e227, 32'h42bbb042},
  {32'hc507f574, 32'h412df910, 32'h424fed9d},
  {32'h4519fe0a, 32'h4373163b, 32'h4361bc80},
  {32'hc42429b8, 32'h43cdcc08, 32'hc34f61d6},
  {32'h43cb9a40, 32'hc36f3c3e, 32'hc3837636},
  {32'hc4a5665c, 32'h42ba8db5, 32'hc351ac0e},
  {32'h44dc2b2d, 32'hc38cb47d, 32'h4379abcf},
  {32'hc4cdc50d, 32'h43ca37ad, 32'hc2c94d6e},
  {32'h4512f6a8, 32'h42e3c25f, 32'h42fae574},
  {32'hc344bf63, 32'hc332f3b1, 32'h4359d79b},
  {32'h443c17b4, 32'hc3030edb, 32'h435bd944},
  {32'hc4a0bd45, 32'hc39efece, 32'hc326cdc7},
  {32'hc20e22c0, 32'hc2c0a2af, 32'hc3601b43},
  {32'hc46e102c, 32'hc35bd8c3, 32'hc351e219},
  {32'h45071dc3, 32'h429ba6ea, 32'hc37e60b6},
  {32'hc50c6b5d, 32'h426cda8c, 32'h42d6420a},
  {32'h43f79dea, 32'hc3ba7a79, 32'h42d75c87},
  {32'hc37e8bf0, 32'hc29fc66d, 32'h430348a5},
  {32'h4447e206, 32'hc3792484, 32'h431f150c},
  {32'hc49a4d99, 32'h43a76f89, 32'h43049255},
  {32'h45257ced, 32'h433604bc, 32'h423f79f0},
  {32'hc4e9197a, 32'h431e24a4, 32'hc3c4b1e5},
  {32'h44273d90, 32'hc34f2001, 32'hc3aa7087},
  {32'hc2cd09c2, 32'h439b2c1b, 32'hc38fae32},
  {32'h4382fc20, 32'h4301babb, 32'h404e4a76},
  {32'hc4d9e45c, 32'hc3a3f6d9, 32'hc3898717},
  {32'h44943aea, 32'hc0c96409, 32'hc247823e},
  {32'hc511a393, 32'h404ebc29, 32'hc301ffb1},
  {32'h4430634c, 32'h433e65b4, 32'h41aaac99},
  {32'hc51fd0e0, 32'hc2d81688, 32'hc25e8c4f},
  {32'h449316b5, 32'hc2605f87, 32'hc0dee34e},
  {32'hc473a70a, 32'hc34513c0, 32'hc228cff1},
  {32'h45065019, 32'h43c280a7, 32'h428353a3},
  {32'hc2f76460, 32'h43dc9ca4, 32'h42d4359e},
  {32'h4400e1fe, 32'h436d0060, 32'hc34a3372},
  {32'hc4dba2fd, 32'hc109d6d6, 32'hc27eeb68},
  {32'h44b5a45b, 32'h42dcb869, 32'hc3290c97},
  {32'hc50ab6e5, 32'hc25c8796, 32'h425ce0e7},
  {32'h451809e0, 32'hc2081a4d, 32'h41e8846c},
  {32'hc38b2f4c, 32'h42ed6f8d, 32'h41622a24},
  {32'h44f81348, 32'h40fa3f08, 32'h432d5085},
  {32'hc4f005e6, 32'h42cc2968, 32'h43cb464f},
  {32'h43b5dd90, 32'h428bfece, 32'h42fe8ef9},
  {32'hc4cb4d58, 32'h420f56fc, 32'hc2cde39a},
  {32'h44e9233a, 32'hc3978fec, 32'h42d45e0f},
  {32'hc4e44986, 32'h4411e873, 32'h422b374c},
  {32'h4504712a, 32'hc2ea5d32, 32'hc395bf6b},
  {32'hc48a4530, 32'hc3b2f0cc, 32'h4397bf63},
  {32'h44328430, 32'hc3a7ed32, 32'hc419fcdb},
  {32'hc41367a8, 32'hc2c78c3e, 32'hc322b9b8},
  {32'h44aab389, 32'h42ae1fbc, 32'hc3b75e2c},
  {32'hc5027854, 32'hc284e4d8, 32'hc3a90302},
  {32'h44bc29f4, 32'hc43aca2f, 32'h4327bbf7},
  {32'hc47cbd88, 32'h4111f108, 32'h43d96ab9},
  {32'h4406cf90, 32'hc37e6699, 32'hc3f88947},
  {32'hc4fe4028, 32'hc285fb2a, 32'h4318535a},
  {32'h44c40b82, 32'h4227d226, 32'h408ad5a6},
  {32'hc38c196c, 32'h420ca2be, 32'h439734ea},
  {32'h44e863fe, 32'hc3555410, 32'h42607050},
  {32'hc4c75b74, 32'h4150a0e5, 32'hc306cc4a},
  {32'h4439f1ea, 32'hc1cb0628, 32'h4289d944},
  {32'hc4b72ee9, 32'hc1b55538, 32'h4340c502},
  {32'h44368a4c, 32'hc2fea555, 32'hc2a5eff6},
  {32'hc4a2f4b6, 32'h43838263, 32'hc16870c2},
  {32'h44fb73d0, 32'hc3b2b9ee, 32'h42e56a65},
  {32'hc3b2f82c, 32'h428e1b15, 32'h4356ed0e},
  {32'h44c76be1, 32'hc24e1701, 32'h4314e862},
  {32'hc333d4a0, 32'h436d20c1, 32'h42d390ab},
  {32'h441a9270, 32'h4280ff7f, 32'hc3c85397},
  {32'hc321ece0, 32'hc3f90616, 32'h43d1fb06},
  {32'h44efb59a, 32'hc2ce9c11, 32'hc369df6d},
  {32'h428d3a73, 32'h435d5687, 32'hc340cb9f},
  {32'h43b2936c, 32'h435a14ff, 32'hc2c50806},
  {32'hc48b37ad, 32'h43a88af1, 32'h433fba84},
  {32'h43fe3c40, 32'hc334458a, 32'h423b8e08},
  {32'hc3516d80, 32'h42e14631, 32'hc27d1d7d},
  {32'h449c65d4, 32'hc29524ba, 32'h428d55fb},
  {32'hc4688d66, 32'h4235688e, 32'h43084105},
  {32'h44affed4, 32'hc3013e46, 32'hc285542a},
  {32'h44d1d0f8, 32'h436e12f7, 32'hc3d4132e},
  {32'hc4e13ffc, 32'h40b6e635, 32'hc30bcfa7},
  {32'h44b0ba58, 32'h418afaf4, 32'h4345fa85},
  {32'hc3c93592, 32'h4276c694, 32'h43156481},
  {32'h45278eda, 32'h43bf3861, 32'hc3e90e7a},
  {32'hc509845f, 32'hc374e7aa, 32'h422d247d},
  {32'h450f97d7, 32'h428de07b, 32'hc3371045},
  {32'hc484cb60, 32'hc2b94465, 32'hc3285dd6},
  {32'h44126c44, 32'h438530e8, 32'hc30f90ae},
  {32'hc485f089, 32'hc3532d45, 32'hc3e7ae55},
  {32'h44f56e23, 32'h41b83a73, 32'hc180738d},
  {32'hc463069e, 32'h4391e4b1, 32'h42c90135},
  {32'h44a8a06e, 32'h422bf3cb, 32'hc2a2a91f},
  {32'hc4705939, 32'h40e1733b, 32'h42981004},
  {32'h4501ab7c, 32'hc38a81a9, 32'h42fd9708},
  {32'hc4a3fb0d, 32'hc2d4cf47, 32'h4203698c},
  {32'h43cb76b6, 32'hc390bb1f, 32'hc3f223ce},
  {32'hc4daa658, 32'hc2975bb6, 32'h42647dcf},
  {32'h4444b116, 32'h42ed589e, 32'h43e61870},
  {32'hc4bbc9ee, 32'h43c8afbb, 32'hc38ecd08},
  {32'hc232e680, 32'h4314adda, 32'h4230e0f1},
  {32'hc46f37ed, 32'hc34808ff, 32'h425686a5},
  {32'h44c9bfc5, 32'hc29c14b0, 32'h420cd543},
  {32'hc500972c, 32'h43330a0e, 32'h43103b95},
  {32'h44ec116b, 32'h4359afba, 32'hc319cafd},
  {32'hc48cc96f, 32'hc2ddf129, 32'h42d9dcf6},
  {32'h43a417c0, 32'hc3875531, 32'h432977ef},
  {32'hc43ab932, 32'h42f7ae2c, 32'hc3ae683d},
  {32'h44b295f9, 32'h4353ba28, 32'h43af7db3},
  {32'hc4a8f75f, 32'h435d6044, 32'hc25bb572},
  {32'h450168ad, 32'h43ab8ca6, 32'h438f7d5f},
  {32'hc4dd1853, 32'hc3974ea6, 32'hc4128290},
  {32'h43d59080, 32'hc27eb9f4, 32'hc3b59aee},
  {32'hc3b6fa1d, 32'hc1bd4a82, 32'hc3fbf80f},
  {32'h44dcc97a, 32'h43440c40, 32'hc2be1464},
  {32'hc4e22191, 32'hc1e1317b, 32'h436154ce},
  {32'h44b0c80d, 32'h439faa99, 32'h42a62fb6},
  {32'hc4856a62, 32'hc305e56b, 32'h42cd57f4},
  {32'h44c6bcde, 32'h42887f59, 32'h416b846e},
  {32'hc4ad73e0, 32'h43079692, 32'hc30470c8},
  {32'h4460fcd7, 32'hc276631e, 32'hc2917cf5},
  {32'hc49d36ec, 32'h4390e838, 32'h43a1cefe},
  {32'h448884f1, 32'hc395179d, 32'h440a7714},
  {32'hc3bde218, 32'h42b3b954, 32'hc35f4c1f},
  {32'h44a4be6a, 32'h42fbce07, 32'h4367f1c8},
  {32'hc5059fdb, 32'h41ec1008, 32'h4179eb1e},
  {32'h44f2228c, 32'hc2e031cf, 32'h43503e1c},
  {32'hc4d77ec8, 32'hc3810728, 32'hc32e615e},
  {32'h44019215, 32'hc361ffbd, 32'h43947991},
  {32'hc4ec57bc, 32'h424e49c9, 32'hc26b904a},
  {32'h4412ac61, 32'hc3a2fe75, 32'h4390438c},
  {32'hc43625ca, 32'h4402fa5c, 32'hc37901b5},
  {32'h44ccb162, 32'h41ff75be, 32'hc2fe9e46},
  {32'hc49546c3, 32'h430acfaa, 32'hc2831d94},
  {32'h44447c26, 32'h434ca0af, 32'h4374f351},
  {32'hc500dfe4, 32'h434c20b5, 32'hc000685a},
  {32'h45205b17, 32'h4335d474, 32'hc34a7f8b},
  {32'hc4d17a80, 32'h41ce1fe8, 32'hc3138c44},
  {32'h4464f310, 32'h43ad08f5, 32'hc2b15fc5},
  {32'hc3b39fd8, 32'h425b269d, 32'hc3d0ff8a},
  {32'h45121b9f, 32'hc1cb932d, 32'h43a2a7a6},
  {32'hc3e1ee86, 32'h437c8d2d, 32'hc0409930},
  {32'h438ae7b8, 32'hc27fa7cd, 32'hc310a773},
  {32'hc3ce9de2, 32'hc312f2ea, 32'h42e511a9},
  {32'h4480fee1, 32'h439ce07f, 32'h43091738},
  {32'hc4e6eed8, 32'hc2d36a59, 32'h4185b377},
  {32'h45037f1e, 32'h438b7448, 32'hc35cafd4},
  {32'hc4cbca22, 32'h3fb8429c, 32'hc2373c1d},
  {32'h442ce44c, 32'h42809458, 32'hc282170b},
  {32'hc4bdfeae, 32'hc2921935, 32'hc31349bc},
  {32'h44f41970, 32'hc269f679, 32'h40495eec},
  {32'hc423726e, 32'hc3d6effa, 32'h43112304},
  {32'h449f3cbc, 32'hc2e2bd14, 32'hc3403fa6},
  {32'hc4b7fb70, 32'h401bfa98, 32'h433a6f7e},
  {32'h4418cea0, 32'h435ab7a2, 32'hc1dbf5ed},
  {32'hc40a0980, 32'h431fec30, 32'h4365f5c8},
  {32'h44b6fdd5, 32'hc36ab962, 32'hc1860ef3},
  {32'hc4e57b98, 32'h42a109f0, 32'hc2c6e93a},
  {32'h44f37a76, 32'hc3c6ba74, 32'h43c245f9},
  {32'hc509761b, 32'hc38949e6, 32'hc03615eb},
  {32'h44b2ff10, 32'h43078b36, 32'h4345faa0},
  {32'hc48891a7, 32'hc2c37241, 32'hc21987c3},
  {32'h44e78312, 32'h43b070be, 32'hc3a50ce8},
  {32'hc436d13a, 32'h43b6b982, 32'hc4071424},
  {32'h4421e771, 32'hc04d3d8b, 32'hc31bedb5},
  {32'hc4ce7279, 32'hc364f666, 32'h41ccd127},
  {32'h4496a765, 32'hc3905b10, 32'hc2d18a61},
  {32'hc5193d47, 32'hc347d74d, 32'hc3df8f23},
  {32'h447d9082, 32'hc30531d2, 32'hc28c03cd},
  {32'hc5055507, 32'h435f97e9, 32'h43920482},
  {32'h443944b1, 32'hc1000e2f, 32'hc244b5a6},
  {32'hc4d14d14, 32'hc0cc51ba, 32'hc26b5cb6},
  {32'h44947490, 32'hc2a3b4bd, 32'h42c16e20},
  {32'hc3e44d40, 32'h43b4e7eb, 32'hc406def1},
  {32'h44a47d86, 32'hc2f42b8b, 32'h4354f806},
  {32'hc4d8fffa, 32'hc2956d37, 32'h43ab88a2},
  {32'h44bac9c0, 32'hc206add7, 32'h43e2c742},
  {32'hc3c38c2c, 32'hc3317170, 32'hc2a407cb},
  {32'h4445199c, 32'h41a07300, 32'h43921f41},
  {32'hc49aa9b0, 32'hc3bc3c01, 32'h438c63da},
  {32'h44e40b8f, 32'hc1dcddc0, 32'h420f72d6},
  {32'hc4269e09, 32'h429c2b27, 32'h4417cf1d},
  {32'h447e43bc, 32'h432ed320, 32'hc2c4572a},
  {32'hc405976c, 32'hc29ede75, 32'h42c86196},
  {32'h44e6adf1, 32'hc112aa71, 32'hc3700a88},
  {32'hc2d561e4, 32'hc32dd3f6, 32'hc2cb5152},
  {32'h446f81dd, 32'hc36d1dfe, 32'h434411ff},
  {32'hc4796304, 32'hc38c78ac, 32'hc2f2b880},
  {32'h44c1af7f, 32'hc3b02e87, 32'hc35d197f},
  {32'hc5055009, 32'hc1f8b7ff, 32'hc38a43e9},
  {32'h4506ee4e, 32'hc3aa9664, 32'hc2dfc248},
  {32'hc49dc609, 32'h43da9556, 32'h41c41e06},
  {32'h44c5b39c, 32'h4365d1c8, 32'h43b2b5c9},
  {32'hc501a6d6, 32'h4401d241, 32'h44186648},
  {32'h42a39e5a, 32'hc1a03d5e, 32'hc3665f28},
  {32'hc4fc424e, 32'hc230e24f, 32'hc2d3ef30},
  {32'h43722500, 32'h43e6b92c, 32'h42bd51d7},
  {32'hc50ca937, 32'h437a5703, 32'h433e6899},
  {32'h44587554, 32'hc2ade465, 32'hc34e21c4},
  {32'hc49df24e, 32'h4229eff0, 32'h42cb5663},
  {32'h4515e112, 32'hc3b6757e, 32'h43b5d5f0},
  {32'hc510b7a7, 32'hc34c60c3, 32'hc35f9e50},
  {32'h44646c3b, 32'h43534f8e, 32'hc2d6d4f9},
  {32'hc4f5118c, 32'hc20bca3c, 32'h43fc86aa},
  {32'h45048fd9, 32'hc317e031, 32'h4399441c},
  {32'hc4479a3b, 32'hbf86f3f2, 32'h4281e5c8},
  {32'h44b5f101, 32'hc1bd136e, 32'h433ae91e},
  {32'hc48e6e2f, 32'hc3402058, 32'hc345f45c},
  {32'h43ad5cb8, 32'h4314c4e7, 32'hc3c8b9b0},
  {32'hc4e6e7ad, 32'hc0f7accc, 32'hc23e0a17},
  {32'h448da829, 32'hc2c16c63, 32'h43c57b46},
  {32'hc39082de, 32'h4366dd6c, 32'hc300e955},
  {32'h44799761, 32'hc1944a30, 32'hc2f9cb96},
  {32'hc52b1a12, 32'h43953fa6, 32'hc3618917},
  {32'h44ada0e4, 32'h4149edf8, 32'h42865e9d},
  {32'hc43a95a0, 32'h42ffb0c6, 32'hc3e8c7de},
  {32'h44b3ef1d, 32'h42ab955e, 32'hc20798ed},
  {32'hc4f31abe, 32'hc3bf1983, 32'h43200dea},
  {32'h447d777a, 32'h43b34302, 32'h4098250b},
  {32'hc4772ce6, 32'h43e9d6f5, 32'hc238dc2c},
  {32'h44b30a70, 32'hc384ab67, 32'hc1a25730},
  {32'hc39317ae, 32'hc31cd65a, 32'h431ce681},
  {32'h432938a0, 32'h429ea26c, 32'h43aecfdd},
  {32'hc44a1381, 32'hc3bcc2b3, 32'hc2a7619d},
  {32'h44c9ad60, 32'hc32f1b51, 32'h42b6e12e},
  {32'hc49d0d5d, 32'h42bce2f9, 32'hc1886411},
  {32'h44f4c5db, 32'h4319d55d, 32'h4307bd52},
  {32'hc4888737, 32'hc386f360, 32'hc3cdf769},
  {32'h44f61215, 32'hc2e92073, 32'hc34a5496},
  {32'hc31efc04, 32'h4327341d, 32'h433f9e80},
  {32'h43bbbfa6, 32'hc19513fc, 32'hc3d582d8},
  {32'hc5018b5f, 32'h42fff8b7, 32'h436b46bf},
  {32'h45038dbc, 32'hc2dc47fb, 32'h41c9e341},
  {32'hc433fb0a, 32'hc2dcf770, 32'h434f5449},
  {32'h450e4008, 32'hc385a076, 32'hc21211ff},
  {32'hc28345e0, 32'hc29033da, 32'h418f9c46},
  {32'h4400e988, 32'hc36c2a6a, 32'h430eaa90},
  {32'hc5082410, 32'hc3cebc93, 32'hc38ea001},
  {32'h44912ebf, 32'hc24371bd, 32'hc2d7b289},
  {32'h432d1a90, 32'h42c81452, 32'h4289f8bc},
  {32'h4485c1ff, 32'hc35a6c6d, 32'h43a1101f},
  {32'hc3cac93c, 32'hc2433dfb, 32'hc18cc520},
  {32'h44e61766, 32'h43310e2e, 32'hc30c8a17},
  {32'hc4c27115, 32'hc3d05b6d, 32'h433ebc70},
  {32'h4508b71e, 32'h42d4cc83, 32'hc1b5c7cb},
  {32'hc400c22e, 32'h418a5fd3, 32'h41e7637d},
  {32'h443e756b, 32'hc3253bc6, 32'hc3cc6755},
  {32'hc448cad2, 32'h42c57658, 32'h43e0a8c5},
  {32'h44bb0694, 32'hc322d3c7, 32'hc3683cc1},
  {32'hc41564e8, 32'hc383f69e, 32'h4381140f},
  {32'h4493befc, 32'hc03f9452, 32'h4392dfef},
  {32'hc4ab919a, 32'h436bce78, 32'h4406c49a},
  {32'h44ba3e5a, 32'hc2f67937, 32'hc3c30248},
  {32'hc4b5f2fc, 32'h42968650, 32'h42dbf9a8},
  {32'h44441f31, 32'h438ab07c, 32'h416c0de0},
  {32'hc47683aa, 32'hc32d1266, 32'h42518ce8},
  {32'h438b78a2, 32'hc284aaf4, 32'h414fd44a},
  {32'hc33878d0, 32'hc4048d52, 32'h42a124d8},
  {32'h44d7ed5d, 32'hc2b6879c, 32'h42c5fe0a},
  {32'h430c6250, 32'h43d7e192, 32'h43942d10},
  {32'h44423560, 32'h40239200, 32'hc20abd4a},
  {32'hc419c6b0, 32'hc370f156, 32'hc2a44348},
  {32'h450f3e73, 32'h43a9210f, 32'hc231e4b9},
  {32'hc3ec3004, 32'hc3141c9b, 32'h42f24f49},
  {32'h44e26fef, 32'h412e757f, 32'h42aa9499},
  {32'hc3c1a032, 32'h419267d7, 32'h432cac14},
  {32'h449b0380, 32'hc22ffbb0, 32'h43027f1f},
  {32'hc4f73d94, 32'h43a20dd2, 32'hc368f633},
  {32'h449b5c9f, 32'h4353e94d, 32'h43158707},
  {32'hc34d5f33, 32'h440edaef, 32'h43752579},
  {32'h449d62fe, 32'h42eaec61, 32'hc31127b6},
  {32'hc4bc93ae, 32'h42d93c87, 32'hc3a998dc},
  {32'h4331c8c0, 32'h412bd700, 32'hc3f20d4d},
  {32'hc4aa6c00, 32'h4313af66, 32'h43ced7be},
  {32'h44f3e6b7, 32'hc224b83c, 32'h43f61461},
  {32'hc4a501e5, 32'h439d5743, 32'h42d1b8cb},
  {32'h44bf91c4, 32'hc239c88d, 32'h430787d9},
  {32'hc4b07fe4, 32'hc274df74, 32'h42728707},
  {32'h43b35e83, 32'h4230fd1a, 32'hc34737a0},
  {32'hc3813837, 32'h43376251, 32'h43724767},
  {32'h45099f48, 32'h41be20fb, 32'h4310f6d4},
  {32'hc4eb58fa, 32'h40e7ee7c, 32'h43006d92},
  {32'h43890310, 32'h4390f309, 32'hc32b35ec},
  {32'hc504ea6b, 32'hc2a753fd, 32'hc2bdeba7},
  {32'h44e470eb, 32'h432602e5, 32'hc2ca2497},
  {32'hc3d42ec8, 32'hc2c4b75f, 32'hc35a7a02},
  {32'h439d027a, 32'hc38b0524, 32'hc2cf0b37},
  {32'hc4439963, 32'hc3845f4d, 32'hc396e472},
  {32'h44d8a1a4, 32'hc2c6ccc8, 32'hc3aa91b1},
  {32'hc4ebee56, 32'h42e0fd78, 32'h42a787c7},
  {32'h44ea4920, 32'h439c1283, 32'hc3a19bac},
  {32'hc4e2e1b3, 32'hc20c3d57, 32'hc2049ac1},
  {32'h44a43bc4, 32'hc2c95b4e, 32'h4420c140},
  {32'hc500db78, 32'h4214fbac, 32'h4382254e},
  {32'h45123cb9, 32'h43bf2757, 32'hc335ecb2},
  {32'h419383d0, 32'hc3691eea, 32'hc37435a8},
  {32'h448832ce, 32'hc328ac16, 32'hc31064a8},
  {32'hc408c3ce, 32'h43c50eb4, 32'hc1fad5d0},
  {32'h44955643, 32'h42bbf4f4, 32'h42bf2d9c},
  {32'hc4d4bd3e, 32'hc391a656, 32'h4331b49b},
  {32'h44b989d4, 32'hc2bb8ec3, 32'hc24f44ea},
  {32'hc2cba8b8, 32'h4296ced5, 32'h4311591a},
  {32'h45066a7d, 32'h43871952, 32'h433e4e82},
  {32'hc4ea1dfa, 32'h432d1216, 32'h430c2a9e},
  {32'h43225578, 32'hc261c162, 32'hc30db394},
  {32'hc490425f, 32'hc2c8fd26, 32'hc29b9b3c},
  {32'h44e616e4, 32'h424e6763, 32'hc2409df6},
  {32'hc4ed6a06, 32'h4300d65a, 32'hc3823976},
  {32'h45028142, 32'h42ade99f, 32'h42aaff0e},
  {32'hc33bc430, 32'h42963375, 32'h43309188},
  {32'h44b42e95, 32'hc2821a0a, 32'h42957051},
  {32'hc4f7d240, 32'h42aeecda, 32'hc38ecb91},
  {32'h4511a3d4, 32'h42b4db47, 32'h43b56c63},
  {32'hc4cd2847, 32'h425b5690, 32'h420d38bf},
  {32'h44c2328a, 32'h43609f44, 32'hc345f210},
  {32'hc3eec3d0, 32'h41cd513b, 32'h43141708},
  {32'h449f3d97, 32'h42bfeb88, 32'hc24d828a},
  {32'hc4d4d4a1, 32'hc35d0030, 32'h433782ca},
  {32'h449669e6, 32'hc1b10f0d, 32'hc3d49b17},
  {32'hc5208645, 32'hc3a61b3b, 32'h434d8cf2},
  {32'h44804624, 32'h421615cf, 32'hc32e9509},
  {32'hc367af63, 32'hc20a4fa9, 32'hc3ab2288},
  {32'h432791e0, 32'hc348896d, 32'hc3536698},
  {32'hc4452f46, 32'h42b91ca9, 32'h42eb2293},
  {32'h43824c6a, 32'h42e4f380, 32'hc1a7c28e},
  {32'hc421f0e3, 32'h4347b539, 32'h4321c40a},
  {32'h44abd1a2, 32'h4248074f, 32'h40a667ce},
  {32'hc3fe6082, 32'hc38c5704, 32'h431493e1},
  {32'h43912684, 32'hc2458982, 32'h43a054fd},
  {32'hc48445a6, 32'h42857ea9, 32'hc2da3828},
  {32'h450642a7, 32'h4302c7a7, 32'h43c7a69f},
  {32'hc4a741de, 32'hc395ad3e, 32'h43c506ac},
  {32'h4486d320, 32'h43927706, 32'h43016b6a},
  {32'hc494c007, 32'h42d9fcee, 32'h4216efab},
  {32'h450926a2, 32'hc33495bb, 32'h4380167d},
  {32'hc4db973b, 32'hc36c270b, 32'hc39e2102},
  {32'h448209b4, 32'hc31cd6c6, 32'hc1951d77},
  {32'hc4c17cd0, 32'h43410e7d, 32'h40a1abfe},
  {32'hc2141b74, 32'hc2c1ecb0, 32'hc2ee593e},
  {32'hc4ed503d, 32'h43a35b8b, 32'h438e85a4},
  {32'h44e86e6f, 32'hc2934912, 32'h436ee23a},
  {32'hc4d6a26c, 32'h438243ee, 32'h42aa91c3},
  {32'h445c947f, 32'h42f6c04c, 32'hc28bad8a},
  {32'hc468f014, 32'h429ce879, 32'h4381d5a8},
  {32'h44deaec2, 32'h43873534, 32'h436dab0b},
  {32'hc4a85c22, 32'h4372e262, 32'h43043a7c},
  {32'h44f732fc, 32'h4353fb2a, 32'hc0fa2b82},
  {32'h43e13548, 32'hc3cf4f2d, 32'h441a42b4},
  {32'h44129ba2, 32'h43546dab, 32'h42bbf7f1},
  {32'hc48d6826, 32'h423c60f3, 32'h4380d3b6},
  {32'h44917553, 32'hc3444279, 32'h43399413},
  {32'hc48122ad, 32'hc165ecdb, 32'h44175164},
  {32'h44f950a2, 32'hc201505b, 32'hc39f2704},
  {32'hc441adfa, 32'h42fac629, 32'hc128f566},
  {32'h45151419, 32'hc3330c3c, 32'h42be09cb},
  {32'hc40f9d2e, 32'hc36a608e, 32'h421eacf9},
  {32'h45063305, 32'h433e8547, 32'h42a0ae68},
  {32'hc46312df, 32'h434f25ac, 32'hc27880e2},
  {32'h44f6bca8, 32'hc1a96eab, 32'hc2220309},
  {32'hc4a327a4, 32'h4202ec75, 32'hc30686cd},
  {32'h44a7157d, 32'hc159833a, 32'hc3470bee},
  {32'hc5064ba9, 32'hc1bb6cce, 32'h43066122},
  {32'h42160d38, 32'h43afc90a, 32'h434e9a66},
  {32'hc5013d5e, 32'h42b66641, 32'h41e35a36},
  {32'h449251db, 32'h4115d98d, 32'hc306891c},
  {32'hc4d3aabf, 32'h432876f8, 32'hc26f8886},
  {32'h451386ce, 32'hc3253db7, 32'hc3597570},
  {32'hc4513af2, 32'h43a8b6be, 32'h43057292},
  {32'h44b67ca1, 32'h434a94de, 32'h43b4a723},
  {32'hc5084c1b, 32'h42733084, 32'hc3822217},
  {32'h4505d3a2, 32'h4383b605, 32'hc2f627c6},
  {32'hc4c30a55, 32'hc4111f95, 32'h430ccde9},
  {32'h41161200, 32'h434d9c5d, 32'h430edcfd},
  {32'hc511fef1, 32'h430f85ce, 32'h41902ccc},
  {32'h44e89ed6, 32'h4238c555, 32'hc38d833e},
  {32'hc40ddb8f, 32'hc3a267bc, 32'h4359acaa},
  {32'h43a9c698, 32'h42c209d2, 32'h43afff0d},
  {32'hc4e5d9ee, 32'hc3934236, 32'hc2ef4917},
  {32'h44955c88, 32'hc360d425, 32'h4293a256},
  {32'hc50ccd7b, 32'h420ef4c2, 32'h42a22bb3},
  {32'h43e57e34, 32'hc3724eb2, 32'hc3960d72},
  {32'hc49ffed5, 32'hc3ea4fbe, 32'h43a5b2e7},
  {32'h44bd1e2f, 32'h42d9e4d5, 32'hc1ee0ed9},
  {32'h4307a6c0, 32'h436fa652, 32'hc399c4aa},
  {32'h44a4a97f, 32'hc24adbe2, 32'hc3a69a24},
  {32'hc3ebafa0, 32'h4409c7f8, 32'h43b5f8a8},
  {32'h4505f672, 32'hc3998f94, 32'h41bb2752},
  {32'hc507da94, 32'h4111b57c, 32'h439f4ab1},
  {32'h44bbda8a, 32'h437f79b6, 32'h43f9c1cb},
  {32'hc508499b, 32'hc3bb25a1, 32'hc23e7f41},
  {32'h4507f64a, 32'h4293e762, 32'hc161f572},
  {32'hc4341b8a, 32'hc1880db8, 32'hc1fc68af},
  {32'h44c2eb11, 32'h424b17da, 32'h4305f571},
  {32'hc47753d6, 32'hc23db213, 32'h416b14f7},
  {32'h44d2b2cc, 32'hc1a8dc28, 32'h43d6226d},
  {32'hc4df6e6c, 32'h42c5a1ea, 32'hc2c75531},
  {32'h44d74bca, 32'h4219e59a, 32'h42f1e6ee},
  {32'hc487996a, 32'h42ade756, 32'hc2a0466e},
  {32'h4460a322, 32'h434420df, 32'hc402a683},
  {32'hc48aa830, 32'h43569ddb, 32'hc31f9b41},
  {32'h44f6cc10, 32'hc32d07dc, 32'h41ec31ce},
  {32'hc2c22ba0, 32'hc2e150cd, 32'hc3635346},
  {32'h44acaafd, 32'h43baae14, 32'h4307c77a},
  {32'hc4f3afc1, 32'h4350be15, 32'hc310bff8},
  {32'h440e6b8a, 32'hc38918ba, 32'hc2ddbdbb},
  {32'hc4a29bfe, 32'h3f3d6b0e, 32'h431fde73},
  {32'h43cd4d88, 32'hc23bb64c, 32'hc38f1369},
  {32'hc4acb1c1, 32'hc316ba1d, 32'h41cb0b2a},
  {32'h438f71c4, 32'h43033719, 32'h436b8a12},
  {32'hc4f97e59, 32'hc2a4d1c4, 32'hc3dc85fc},
  {32'h44eb16a3, 32'h42b92f0d, 32'hc330d35a},
  {32'hc49e4cdc, 32'h4355ff3f, 32'hc081fe78},
  {32'h44c9d483, 32'h422fc483, 32'hc2efee61},
  {32'hc51494b5, 32'h438ed3f4, 32'h4359e10f},
  {32'h4503b891, 32'h43684922, 32'h43115bd9},
  {32'hc4fd8c78, 32'h41ee478f, 32'hc383cc85},
  {32'h45066d6b, 32'hc29a1e5e, 32'hc2dd7503},
  {32'hc4a2e00b, 32'h42e64d77, 32'hc404f687},
  {32'h44fe62b5, 32'h43429aff, 32'hc2563763},
  {32'hc50da55c, 32'h42ef627c, 32'h43494b27},
  {32'h44da9140, 32'h4327ad8d, 32'h42050c51},
  {32'hc51dc93a, 32'hc2b2c836, 32'hc323aa2d},
  {32'h4402f54b, 32'h40468464, 32'hc32b8379},
  {32'hc50ddf23, 32'h4226fca9, 32'h4321d9b5},
  {32'h4490014f, 32'hc3864b81, 32'hc3523156},
  {32'hc4db932f, 32'h43411232, 32'hc3050bd7},
  {32'h44b0ba0f, 32'h43d89c37, 32'h44156204},
  {32'h421edf00, 32'hc301c82b, 32'h43a177b5},
  {32'h45002da2, 32'h43833c4e, 32'h4341fa46},
  {32'hc45cae74, 32'h43071f38, 32'h43b6fd5a},
  {32'h44ba03c9, 32'hc3e54e9e, 32'hc35dfcf0},
  {32'hc394ec9c, 32'h43359580, 32'hc206aba6},
  {32'h44abb108, 32'hc3465bab, 32'h41b1227b},
  {32'hc42cfe9c, 32'h42d07dda, 32'h43a5bd74},
  {32'h44079b20, 32'hc143c92a, 32'h41cc2b47},
  {32'hc3fd4c18, 32'h416a81d6, 32'h4366b955},
  {32'h44920820, 32'hc33edd70, 32'hc187bfd4},
  {32'hc326bb6c, 32'hc2d08cac, 32'h4191f816},
  {32'h44b06805, 32'h43aac76a, 32'hc1cf7859},
  {32'hc46d3c74, 32'hc4048424, 32'h434ea020},
  {32'h44cb6bb4, 32'h41df2d2b, 32'h41750e80},
  {32'hc4c1dd88, 32'h4337cb0c, 32'h43f4c4a8},
  {32'h43bb4416, 32'h43120033, 32'hc2efeecc},
  {32'hc50a5e13, 32'hc21520a4, 32'h439edaf3},
  {32'h43de0818, 32'hc3843b75, 32'h4329cc8a},
  {32'hc4acabc2, 32'hc31bcaf2, 32'hc28ad996},
  {32'h44e3ad5f, 32'h438d5915, 32'hc3491de2},
  {32'hc502a0fa, 32'hc2d94b91, 32'hc35779e8},
  {32'h4420963b, 32'hc35ae8c3, 32'h4277d342},
  {32'hc4be5ffe, 32'h42fdf355, 32'h43db5569},
  {32'h43871f66, 32'hc34345d5, 32'h42cfcbe3},
  {32'hc2a418f7, 32'hc3a5b16b, 32'h428a286d},
  {32'h44bc46f0, 32'hc397f0f6, 32'h42be63da},
  {32'hc4f9904b, 32'hc2c2f6f9, 32'h428dfed0},
  {32'h4522d17a, 32'hc3b09931, 32'h439e07a1},
  {32'hc4156096, 32'hc33df95e, 32'h424e3dd8},
  {32'h44e37c94, 32'hc31076db, 32'h43c0b62c},
  {32'hc4a7b5a8, 32'h439271fc, 32'hc3874001},
  {32'h45036864, 32'h4221f324, 32'hc2a838d0},
  {32'hc4f90950, 32'hc3243507, 32'h41bc1fd3},
  {32'h43bc3250, 32'h43739516, 32'hc3ae0d24},
  {32'hc50dadaa, 32'h4333397d, 32'hc2971bcf},
  {32'h452b70b1, 32'hc3ac5ad1, 32'h4305a260},
  {32'hc27c8380, 32'h43937195, 32'hc385c0bc},
  {32'h43562266, 32'h4112679e, 32'h440c65bf},
  {32'hc484f46a, 32'hc35848d6, 32'hc1b1e686},
  {32'h4509aa6e, 32'hc272d49b, 32'hc269a9ea},
  {32'hc4ac4504, 32'h4427d4aa, 32'h43ae00a5},
  {32'h4516c779, 32'h42984520, 32'h41a40ac8},
  {32'hc51864cc, 32'hc3077ea7, 32'h43efad9b},
  {32'h44807b8e, 32'hc3989838, 32'hc3edbb74},
  {32'h43102f50, 32'hc355d455, 32'h41f5283d},
  {32'h451e5ec4, 32'hc365f1de, 32'hc3f64ad8},
  {32'h43d42080, 32'hc1f11347, 32'hc3465f50},
  {32'h44f283c7, 32'h436af5e9, 32'h43261e18},
  {32'hc3bb508c, 32'hc3a02e41, 32'hc202e087},
  {32'h44d00c41, 32'hc2197cb9, 32'h4336e80b},
  {32'hc31e3582, 32'h42ac81a1, 32'hc386269f},
  {32'h44ebe6fc, 32'h43255d7a, 32'h43215019},
  {32'hc43214c6, 32'hc2eeae6c, 32'hc3823dea},
  {32'h43c94770, 32'hc4312420, 32'hc3336d25},
  {32'hc31a26cc, 32'h436ea772, 32'hc3ab1b24},
  {32'h44d6eadd, 32'hc3308dec, 32'hc314abc2},
  {32'hc49b4f70, 32'h413008c4, 32'hc3e3e4d9},
  {32'h44846737, 32'hc38bd3ba, 32'h4302ce30},
  {32'hc4ed2d15, 32'hc30c4b80, 32'hc30c597c},
  {32'h4408ce2a, 32'h4350227b, 32'hc3448e14},
  {32'hc50ac528, 32'h4342dfde, 32'h419e521b},
  {32'h449a8c76, 32'h43221e92, 32'h428de2de},
  {32'h439d7e68, 32'hc3537d5f, 32'h42c64acc},
  {32'h43a2319b, 32'h435b2a2b, 32'hc3c26c47},
  {32'hc4ea689b, 32'hc2505782, 32'h43a0e403},
  {32'h4408eff8, 32'h438298f5, 32'h43797d6d},
  {32'hc4f36951, 32'h43209e84, 32'h43681b16},
  {32'h4512d062, 32'h42702286, 32'h43832e08},
  {32'hc4c62d1e, 32'hc3719ef2, 32'h4391f2ba},
  {32'h44d818d0, 32'h41a4bd44, 32'h43c80aeb},
  {32'hc348fdbc, 32'hc2124d9f, 32'hc1eb319b},
  {32'h4454a81b, 32'hc341900f, 32'h436b2516},
  {32'hc502fb6e, 32'h42b108fe, 32'h42d989c8},
  {32'h4404a7b0, 32'h427d191d, 32'hc24626b5},
  {32'hc48cb738, 32'hc3297a6e, 32'h42371483},
  {32'h44427884, 32'hc2f3a86d, 32'h42e19f16},
  {32'hc4935027, 32'h41e60544, 32'hc39c3e52},
  {32'h44e002c7, 32'h4294e078, 32'hc2977c47},
  {32'hc4def612, 32'h43a492ea, 32'hc371617f},
  {32'h4493e72f, 32'h432b73df, 32'h43092910},
  {32'h40401c00, 32'hc39c1b8e, 32'h425f6bab},
  {32'h4492082f, 32'h439c9a63, 32'hc2985beb},
  {32'hc4614b86, 32'hc2bd5c85, 32'h4173366e},
  {32'h44ba257b, 32'hc3114458, 32'h42a5a5dc},
  {32'hc4f9b7af, 32'h425f887b, 32'h42cf6c17},
  {32'hc4b8f7a7, 32'hc14a5c46, 32'h4285f989},
  {32'h43cece3c, 32'h41eadef3, 32'h43d418d9},
  {32'hc3af5d49, 32'hc414696a, 32'hc32b8b42},
  {32'h44d92f73, 32'h4389bb66, 32'h430aaeb9},
  {32'hc491739e, 32'hc3562ebb, 32'hc3934fef},
  {32'h4499fc81, 32'h4322e68d, 32'hc2ff6a0e},
  {32'hc4ea4fd6, 32'hc213b87f, 32'h4333df4d},
  {32'h45228d7a, 32'hc2678c4b, 32'hc321d3b4},
  {32'hc430b322, 32'hbfb34c68, 32'hc3a2a1ee},
  {32'h44b19448, 32'h4290423d, 32'hc1853679},
  {32'hc4f12c3f, 32'hc3733f4f, 32'hc3e5f2ca},
  {32'h44f6a665, 32'h42d65237, 32'h43f990d9},
  {32'hc357ff44, 32'h43427787, 32'hc2435dc0},
  {32'h44a419f0, 32'h43ace677, 32'h438ca84b},
  {32'hc24b8d10, 32'h43769caa, 32'hc308c588},
  {32'h44d4bbfa, 32'h42d8db21, 32'hc2f8fbc1},
  {32'hc50f94ee, 32'hc3d6e080, 32'hc2370b84},
  {32'h43eb5e74, 32'hc3918d6e, 32'hc1e90dba},
  {32'hc32cdfdc, 32'hc355d686, 32'hc20e958b},
  {32'h4421e4f8, 32'h430dcca6, 32'h429e75ee},
  {32'hc4eb640e, 32'h433d5ae7, 32'hc3c36097},
  {32'h44b08ea0, 32'h438a9364, 32'h43c82109},
  {32'hc48c1a1e, 32'h43500acf, 32'h42f26cac},
  {32'h45056c86, 32'h43357c35, 32'h428b5d64},
  {32'hc4a6a66f, 32'hc31a4a34, 32'hc2f9d6f4},
  {32'h446bd068, 32'hc2f151be, 32'hc1d86618},
  {32'hc4d8774f, 32'h439504fa, 32'h42680af9},
  {32'h4400ef90, 32'hc334bf73, 32'hc3b021d8},
  {32'hc4ec8df2, 32'h43380646, 32'h422b1620},
  {32'h4504118e, 32'hc22dc07d, 32'h41c89252},
  {32'hc5086ea2, 32'hc34d892e, 32'h42b7455e},
  {32'h44d67b5a, 32'h42ed07a3, 32'hc3238b52},
  {32'hc417544e, 32'hc305e812, 32'hc379ff71},
  {32'h448a0832, 32'hc27e7b8d, 32'h42c86c22},
  {32'hc5057abd, 32'hc3474091, 32'h43a5a78b},
  {32'h44604809, 32'hc38a793a, 32'hc311a8a1},
  {32'h42c8fe6c, 32'hc341b45e, 32'h4127bc9a},
  {32'h44a6820b, 32'h42e01914, 32'h4245f335},
  {32'hc3f66f38, 32'hc3745e46, 32'h435df12f},
  {32'h44b0d263, 32'hc360b6a1, 32'hc2aee2d9},
  {32'hc4816da1, 32'hc323cd96, 32'hc3883719},
  {32'h44e1d158, 32'hc3461d68, 32'h4274e8ba},
  {32'hc50616df, 32'hc2c4be8a, 32'h4295c932},
  {32'h4502d88f, 32'hc42efbf2, 32'h44203b52},
  {32'hc510096e, 32'h43434cd1, 32'h43efedb7},
  {32'h44b938e6, 32'h41b1f59e, 32'hc28027a9},
  {32'hc4fb4014, 32'hc22870b0, 32'h42cfbed8},
  {32'h44e62900, 32'hc2ed9724, 32'h4323b7ae},
  {32'hc44867ea, 32'hc2dc4e8e, 32'hc371200c},
  {32'h4444fdaa, 32'hc36157d5, 32'h435d913b},
  {32'hc48906eb, 32'h442a4f28, 32'hc4190c18},
  {32'h4441a1d8, 32'hc24b64ea, 32'h42eab3a2},
  {32'hc49624ac, 32'hc3506aa3, 32'hc2f4aad7},
  {32'h4352a404, 32'h42c9e924, 32'h4327cbbe},
  {32'hc4cfec86, 32'hc2245f75, 32'hc2cc706f},
  {32'h450f2d18, 32'h42f93d35, 32'hc370ad0d},
  {32'hc4cee722, 32'hc3a870aa, 32'h432f23ef},
  {32'h4503bd54, 32'hc3b92371, 32'hc3f938a1},
  {32'hc4ea347a, 32'h411c2e0f, 32'h4352d987},
  {32'h449f2578, 32'hc40a808e, 32'h429d1fb1},
  {32'hc4756e6f, 32'hc3898ef9, 32'hc3b02fde},
  {32'h450b8ede, 32'hc1630ef7, 32'h43e96bc9},
  {32'hc4306426, 32'h42035162, 32'h43019b7e},
  {32'h43d607b2, 32'h43cdb5f5, 32'h430b5305},
  {32'hc410dc60, 32'h4312ed96, 32'hc2f20cc7},
  {32'h4463455a, 32'hc413e5b5, 32'h44026806},
  {32'hc4266c34, 32'hc304d384, 32'hc338a693},
  {32'h4396fff8, 32'hc2ac2968, 32'hc2b42ffe},
  {32'hc3c2b911, 32'hc3980e73, 32'hc340da90},
  {32'h44f7d428, 32'h43edb085, 32'h43a86303},
  {32'hc4fc9663, 32'hc394ce5f, 32'h438e82b6},
  {32'hc3720770, 32'h438d9031, 32'h413680b4},
  {32'hc43a289e, 32'h43a49b14, 32'h4272eec2},
  {32'h43b53e82, 32'h43c55a09, 32'h42739d10},
  {32'hc43cbe64, 32'hc374f311, 32'hc36aa340},
  {32'h42a824f8, 32'hc21ed2c5, 32'hc27a33ff},
  {32'hc5013159, 32'hc3a3e288, 32'h424b2677},
  {32'h44c190b2, 32'hc1daebab, 32'h438f7b75},
  {32'hc4c8531d, 32'hc327044e, 32'h429d480e},
  {32'h44098df0, 32'h43259078, 32'h438ed66a},
  {32'hc4d6f9b0, 32'h40d45e2f, 32'hc3edb024},
  {32'h4445d516, 32'hc40338dd, 32'h42becdfb},
  {32'hc5071e1c, 32'h41d7d5f8, 32'hc32ab6e8},
  {32'h4445642f, 32'hc312e9ed, 32'hc31d336e},
  {32'hc51dec19, 32'h4289b215, 32'hc3739184},
  {32'h4502ff88, 32'hc1cde040, 32'h44119b2c},
  {32'h4399f02b, 32'h440ae244, 32'h43948562},
  {32'h4401d1a0, 32'hc37bc8b5, 32'h41d97bed},
  {32'hc4db9e50, 32'h41eaf52e, 32'h433c162b},
  {32'h4291f2a0, 32'h43520553, 32'h4374f527},
  {32'hc4c36048, 32'hc3b69fec, 32'h42ea51dc},
  {32'h450b937e, 32'h41cb1899, 32'hc2b0ea48},
  {32'hc4cab6a5, 32'h438051aa, 32'h440947b6},
  {32'h445a8a5d, 32'hc3244f65, 32'hc20218ad},
  {32'hc4f3d026, 32'h431e631f, 32'hc283ae6f},
  {32'h44893090, 32'h41891e97, 32'hc3684581},
  {32'hc4dede46, 32'h419c645a, 32'hc33a3f1c},
  {32'h4426d2b8, 32'hc1a6dc75, 32'hc283ae26},
  {32'hc3a14a94, 32'h41ff946c, 32'hc23bcad0},
  {32'h441c03b8, 32'h439a062e, 32'h42ea011d},
  {32'hc43d3572, 32'hc22334b2, 32'h429263a1},
  {32'h44ffdb8e, 32'h4380102b, 32'h42ef120c},
  {32'hc5151de6, 32'hc344270a, 32'hc31974d9},
  {32'h44f1ac68, 32'hc23f7f26, 32'hc354afb3},
  {32'hc50d284b, 32'hc1ecccdd, 32'h438b401e},
  {32'h443b5b16, 32'h4160abda, 32'h42e9f1d1},
  {32'hc4773358, 32'hc313be9b, 32'h433a890a},
  {32'h44641980, 32'hc314419a, 32'hc0dbe3cb},
  {32'hc4afa61a, 32'hc3784589, 32'h435e1ea4},
  {32'h44ecb0b2, 32'h43816430, 32'h43799675},
  {32'hc2946ac0, 32'hc1c93dd8, 32'h42112b42},
  {32'h44ac713c, 32'hc2a93cab, 32'hc19b85e1},
  {32'hc4936c50, 32'hc30d3298, 32'h42350a4b},
  {32'h4483195a, 32'hc39ce7ec, 32'h43e2e4a2},
  {32'hc33ff5e2, 32'hc2b708c7, 32'h4325a76c},
  {32'h4438727c, 32'h43f91660, 32'hc1801a02},
  {32'hc4eaabbe, 32'hc31302f3, 32'h435ad361},
  {32'h442bef86, 32'hc35076fb, 32'hc2c91fa7},
  {32'hc48ff6f2, 32'h43b5c5ee, 32'h42bf39f4},
  {32'h4504013c, 32'h43c325a7, 32'hc11c4da6},
  {32'hc50766b9, 32'h426e5d8a, 32'hc1f0bb72},
  {32'h447439c0, 32'h43afafbb, 32'h43b466d1},
  {32'hc3d714bc, 32'h439c0944, 32'h431a1406},
  {32'h43706938, 32'h4339a62f, 32'h432f16fa},
  {32'hc4d71562, 32'h43787126, 32'hc35c0075},
  {32'hc18ef200, 32'h4375959b, 32'hc3b056b2},
  {32'hc468c016, 32'hc3121b05, 32'h42b3ca18},
  {32'h44ae7020, 32'hc395662c, 32'h422635f4},
  {32'hc4f0b64a, 32'hc2ca36c2, 32'h428895ea},
  {32'h44b3b468, 32'h4362141d, 32'h43450205},
  {32'hc3aac970, 32'h431b1b41, 32'hc2e20896},
  {32'h43b10370, 32'hc38b4abc, 32'hc3a55232},
  {32'hc4740317, 32'hbff48030, 32'hc3671f84},
  {32'h45138ec4, 32'h433afb23, 32'h439a9eb8},
  {32'hc4105723, 32'hc1d361e0, 32'hc3177dde},
  {32'h4500f184, 32'hc34cd810, 32'hc33818fb},
  {32'hc322b3a2, 32'h416b777b, 32'h433a40e1},
  {32'h448e14a1, 32'h429aeb6d, 32'h42841973},
  {32'hc40989de, 32'hc1a995b3, 32'hc3089947},
  {32'h450aa61c, 32'h4323e95a, 32'h42a91169},
  {32'hc41e701f, 32'hc1bb0d8e, 32'hc383a2c5},
  {32'h4221c280, 32'h4377162e, 32'hc38ae6ba},
  {32'hc5014190, 32'hc312d48c, 32'h4182f5d6},
  {32'h4419e53d, 32'hc3ccf9de, 32'hc2f06d1f},
  {32'hc4b5a00a, 32'hc2d7f65e, 32'h4375fba6},
  {32'h44e496f4, 32'h433e63df, 32'h4221968f},
  {32'hc4d7d996, 32'h41210df8, 32'hc299b0e7},
  {32'h44f5b068, 32'hc30aef57, 32'h4299eb8d},
  {32'hc384a00a, 32'hc3970e96, 32'hc3c03fa1},
  {32'h43d22660, 32'hc3f4fa03, 32'hc34e77f4},
  {32'hc4760f2c, 32'hc308976d, 32'hc385ae77},
  {32'h44421b72, 32'h430e33fa, 32'hc3c8a4b7},
  {32'hc4264898, 32'hc2e47109, 32'h4370e6f0},
  {32'h44edef52, 32'h4374894a, 32'h42c601e2},
  {32'hc4a4ddd2, 32'h432a7185, 32'h42e3147e},
  {32'h4501347c, 32'hc301bb19, 32'h42a28860},
  {32'hc429e9c5, 32'hc281f8c7, 32'hc337087f},
  {32'h44be504b, 32'h42e0aafa, 32'h438e7e68},
  {32'hc4c63b8b, 32'hc3d93319, 32'hc1cb8d70},
  {32'h4406e97d, 32'hc38585f5, 32'hc1993eb6},
  {32'hc4ab15fe, 32'hc3884554, 32'h43906d95},
  {32'h44d7a9b3, 32'hc34aed3f, 32'hc39294ae},
  {32'hc4e4ec5a, 32'h436d40f4, 32'hc283d3ae},
  {32'h45035269, 32'h4279831d, 32'hc31ca3ab},
  {32'hc50801db, 32'h4315e97c, 32'h41f2af0f},
  {32'h432bc9e0, 32'h4285709b, 32'h43344a0a},
  {32'hc4a2aed6, 32'hc31d8b27, 32'h43b3602b},
  {32'h4314d210, 32'hc310a2ad, 32'hc2d26047},
  {32'hc4a84958, 32'hc29addc3, 32'hc30112bb},
  {32'h43c9fcb2, 32'hc1a6b641, 32'hc3405c1e},
  {32'hc4afd95e, 32'h43978c11, 32'h3f2500e8},
  {32'h43f4b034, 32'hc3373988, 32'h4433e4e3},
  {32'h4303a448, 32'hc39d67ce, 32'hc30b4a73},
  {32'h44d9c956, 32'hc37e0e1a, 32'hc4246d13},
  {32'hc4d56bc5, 32'h42925848, 32'hc26fac48},
  {32'h44485914, 32'h43bb4d1e, 32'h4308d156},
  {32'hc367b8d8, 32'hc357d157, 32'hc2483974},
  {32'h44fc44d5, 32'h4359bf95, 32'hc1c0711c},
  {32'hc457d1c2, 32'hc2ddfc60, 32'hc40040f6},
  {32'h44aaef64, 32'hc243350f, 32'hc388b0fd},
  {32'hc307431a, 32'hc3b79739, 32'h43ccc9a0},
  {32'h43e04062, 32'hc4465d3b, 32'h42a4b060},
  {32'hc3ffb494, 32'hc22262ee, 32'hc2e3f665},
  {32'h4505d573, 32'h436314cd, 32'h43c6c455},
  {32'hc47fe42c, 32'hc39c7550, 32'h437c87b9},
  {32'h44cd76f0, 32'h431d4e61, 32'hc3036fee},
  {32'hc5065248, 32'h42ae1b39, 32'h43a54f7a},
  {32'h45061858, 32'hc22e86d6, 32'h422f315c},
  {32'hc500fe8d, 32'h42a174ad, 32'hc3e48c7f},
  {32'h4492ef2a, 32'h3ffb18c0, 32'h421538cd},
  {32'hc4239df0, 32'h42810a84, 32'h43f7ed53},
  {32'h450b0f7a, 32'h41376ede, 32'h43373054},
  {32'hc48d1765, 32'hc3b03810, 32'h42ac752e},
  {32'h44d46afc, 32'hc0382a14, 32'hc343fed9},
  {32'hc4073b15, 32'hc3961df3, 32'hc37e6e24},
  {32'h43c744fc, 32'hc2c77f50, 32'hc223aea4},
  {32'hc408692a, 32'hc2b0abac, 32'h4377189e},
  {32'h42a11a60, 32'h42abec2b, 32'h42a7e25b},
  {32'hc4299b94, 32'hc36fd78e, 32'hc33a7e14},
  {32'h44698960, 32'hc3075f47, 32'h436491ec},
  {32'hc4e14f22, 32'h43ee6841, 32'h4339aa46},
  {32'h4460b65e, 32'hc349dd56, 32'h42cf9464},
  {32'hc497d958, 32'hc31bca40, 32'h432b3f24},
  {32'h44996dc1, 32'h42dce322, 32'hc208e394},
  {32'hc45460e6, 32'hc3571839, 32'h43b75bf7},
  {32'h44520c16, 32'h43710a47, 32'h42344532},
  {32'hc5123c90, 32'h439f48f9, 32'h4389b06e},
  {32'h44f8e806, 32'hc3abd500, 32'h4314aeee},
  {32'hc4dc82fb, 32'h427810ae, 32'hc31f2447},
  {32'h43c3bad5, 32'hc3a661e5, 32'hc3704d4f},
  {32'hc33c6cd0, 32'h43f1fd1e, 32'hc3d70dfb},
  {32'h44f9064a, 32'hc29579ea, 32'hc3f07c9e},
  {32'hc3f8ac8c, 32'h426e3f10, 32'hc3e27ff7},
  {32'h44e1ffa4, 32'hc3f7389f, 32'h425c51f0},
  {32'hc4d42daa, 32'h42252759, 32'h42d4e694},
  {32'h44b41dbd, 32'h42a301e1, 32'hc3a7441b},
  {32'hc505de4f, 32'hc384e133, 32'h417febfc},
  {32'h4500b4dc, 32'hc2547e49, 32'h41f6cd9c},
  {32'hc32d3250, 32'h411dc82e, 32'h4376e710},
  {32'h4461ba94, 32'h4395bfc8, 32'h429c3d61},
  {32'hc4e96c7d, 32'h43203eb7, 32'hc31ac9d8},
  {32'h44e7b90b, 32'h43d7ecf3, 32'hc294599c},
  {32'hc364b8f8, 32'h42b3b7f7, 32'hc219ce90},
  {32'h45120553, 32'h43cffaa4, 32'hc37f9752},
  {32'hc48d3103, 32'h43a8022c, 32'h42e998b8},
  {32'h44dcabf8, 32'hc3873220, 32'hc3a2d1e8},
  {32'hc487822c, 32'h42cb0966, 32'h43298783},
  {32'h43c60150, 32'h411083dc, 32'h4412521b},
  {32'hc4a9ca88, 32'hc3a43df6, 32'hc2a12db2},
  {32'h44a19b38, 32'h43dbd953, 32'hc38edbe3},
  {32'hc3bb8dc4, 32'h438b3ab6, 32'h435e49ad},
  {32'h44d05e3f, 32'h43533fed, 32'h43f26898},
  {32'hc4f8e727, 32'h4316a9a8, 32'h43902f2e},
  {32'h4509da97, 32'h42df3228, 32'h430f2655},
  {32'hc4d49434, 32'h423e7672, 32'h4265e325},
  {32'h442f718a, 32'hc2b9f941, 32'hc20fc08b},
  {32'hc3fc4521, 32'h438b145e, 32'hc3d2878c},
  {32'h445ea511, 32'h42f3d517, 32'h43473a45},
  {32'hc48fef91, 32'hc2e062bb, 32'hc361651b},
  {32'h44b70282, 32'hbf4c8200, 32'h441c5ede},
  {32'h43756c58, 32'h433bce01, 32'hc396fc2d},
  {32'h44b89e8a, 32'hc1606f43, 32'hc3a4e523},
  {32'hc38a7860, 32'hc3227798, 32'hc2a30a06},
  {32'h4304b2b2, 32'hc1a6e445, 32'h42f3c8e1},
  {32'hc3da9dff, 32'h438c19f5, 32'hc3160300},
  {32'h44a22262, 32'h43ba1c9a, 32'h4308c904},
  {32'hc4f8eb4a, 32'hc23ec735, 32'hc371e5aa},
  {32'h427e8cc0, 32'hc26b861b, 32'h42356910},
  {32'hc4ce8abc, 32'hc272539e, 32'h43b0bfae},
  {32'h44a9f903, 32'h4343f657, 32'hc410fd54},
  {32'hc4cbfa04, 32'h430e3b30, 32'h411e5c1a},
  {32'h43dffd52, 32'h42ecf01a, 32'h42905357},
  {32'hc505a5d2, 32'hc27c3b13, 32'h42f4bc13},
  {32'h44c2d6bf, 32'h43080558, 32'h434283db},
  {32'hc4bb0a8e, 32'hc375a5f0, 32'h41545fc2},
  {32'h4240a6cc, 32'h410cbece, 32'h438c15e2},
  {32'hc4658a06, 32'hc392aab0, 32'hc23032d6},
  {32'h44c71061, 32'hc34dfd93, 32'hc2cbaa3c},
  {32'hc46e88f4, 32'h4380a7c6, 32'hc3394330},
  {32'h449299af, 32'hc38e0f84, 32'hc2554d2a},
  {32'hc5192355, 32'hc343ac36, 32'hc3b2edb5},
  {32'h4322c972, 32'h43d86685, 32'h41824b2d},
  {32'hc472ee7c, 32'hc3663e51, 32'h42aeb869},
  {32'h44b3850e, 32'hc3158669, 32'hc324d1b9},
  {32'hc467f8ee, 32'hc317a8e7, 32'h432885e1},
  {32'h44aca4cb, 32'h435dcb6b, 32'h43a44962},
  {32'hc45e4b66, 32'h42c4f5b4, 32'hc3083f1d},
  {32'h4427df38, 32'h4361b8f6, 32'hc0a20d1e},
  {32'hc4aa4184, 32'h4251532e, 32'hc2908fb9},
  {32'h4507a408, 32'hbfabfea0, 32'hc34a82c2},
  {32'hc4bdc61b, 32'hc39a3a47, 32'hc26ee4ad},
  {32'hc1992860, 32'h43068974, 32'h4387cdce},
  {32'hc4fa6f6c, 32'hc16a2850, 32'h43cd46ad},
  {32'h451016e1, 32'hc187ddec, 32'hc2d1c31c},
  {32'hc2cb87e0, 32'hc31656fe, 32'hc412a682},
  {32'h44eb87c4, 32'h43bb81c8, 32'hc220e5ad},
  {32'h40690758, 32'h43bddf4b, 32'hc3378a46},
  {32'h44c66b5e, 32'h41d7aff0, 32'h43b7b5cc},
  {32'hc3a25c10, 32'h43226887, 32'hc3197e02},
  {32'h439efe3d, 32'hc35687e3, 32'hc2af1838},
  {32'hc4a1c68d, 32'h44037b2c, 32'h42c1a4ab},
  {32'h44dc5b0f, 32'h41c89f3c, 32'hc3b4915d},
  {32'h434cd2a9, 32'hc119c7d9, 32'h42c1e662},
  {32'h44a45eb6, 32'hc0a506ed, 32'h415f48d1},
  {32'hc4e690a9, 32'h41c53960, 32'hc069cf8d},
  {32'h445ae3b2, 32'hc308fc0a, 32'h439137f3},
  {32'hc41dbd9f, 32'h4351bfec, 32'h42d96e15},
  {32'h44db8fa1, 32'h427e3804, 32'hc295f366},
  {32'hc43264e9, 32'h43959100, 32'hc1e4894e},
  {32'h448d9422, 32'h43fffb23, 32'hc28329b6},
  {32'hc461dd26, 32'hc1c71828, 32'hc39f49ef},
  {32'h4491dbcc, 32'hc314e242, 32'h4302c56e},
  {32'hc38cdee6, 32'h42b08333, 32'h42f69dcf},
  {32'h44ec612f, 32'h415d39e6, 32'hc362d96c},
  {32'hc4a82dc2, 32'hc35d5211, 32'hc2de8027},
  {32'h451616b0, 32'hc2d9d9f4, 32'h4315d9df},
  {32'hc43ec154, 32'h439cd82e, 32'hc30f5f02},
  {32'h449c30a7, 32'h42ac3a5f, 32'h43e59d01},
  {32'h43078042, 32'h4388f8f8, 32'hc38ce87e},
  {32'h44de693e, 32'h43d309f4, 32'hc2e3ec60},
  {32'hc515231f, 32'hc30e796b, 32'h41931820},
  {32'h44846ed3, 32'h430cf2ab, 32'hc35ab35b},
  {32'hc4dcb144, 32'h42c28f3b, 32'h43ccb4f4},
  {32'h44dbdca1, 32'hc4072501, 32'h41cc9d97},
  {32'hc4ca969e, 32'hc166ad28, 32'h42a8a6b9},
  {32'h44d8d979, 32'h4361513d, 32'hc300094f},
  {32'hc4deed98, 32'hc362b21f, 32'hc421bce3},
  {32'h448dac9c, 32'h42e4c151, 32'h4217cef7},
  {32'hc4c1825e, 32'hc330584a, 32'h4182d926},
  {32'h4517a860, 32'hc38f91dd, 32'hc3e3af10},
  {32'hc45463b2, 32'hc39b814b, 32'hc3581900},
  {32'h44f25c22, 32'h4369ace7, 32'h435151e9},
  {32'hc44de322, 32'hc32594d2, 32'h42118e1e},
  {32'h44cac025, 32'hc386fd05, 32'h4399e89f},
  {32'hc4d1b89c, 32'hc3915e50, 32'h4300e9aa},
  {32'h44816590, 32'h4223a780, 32'hc2dca3d8},
  {32'hc49f4bbc, 32'h4431428b, 32'hc1e1a604},
  {32'h44a57c99, 32'hc2952eef, 32'h430d3775},
  {32'hc440ac19, 32'h4267f9d4, 32'h435f0c0a},
  {32'h45006f1d, 32'h4257e6c2, 32'h43264026},
  {32'hc503f1e7, 32'h43191aec, 32'h4408a979},
  {32'h442192ce, 32'hc2e41cb4, 32'h4403f475},
  {32'hc3376090, 32'h436d85d6, 32'hc322c3ae},
  {32'h435efa08, 32'h438cbdd9, 32'hc39a9ad4},
  {32'hc485a835, 32'h42d50c6c, 32'hc1e0c8e8},
  {32'h448a3312, 32'h42b1d356, 32'hc24ce825},
  {32'hc49eb0f8, 32'hc26616fa, 32'hc1595115},
  {32'h4481ff04, 32'h43b39371, 32'h423a34a5},
  {32'hc49b8574, 32'h42d4c846, 32'hc3849411},
  {32'h4507b130, 32'hc3c65cda, 32'h437996cb},
  {32'hc4d3adfc, 32'h4301edd2, 32'h432c94e4},
  {32'h44d20465, 32'hc35c4745, 32'hc29c162b},
  {32'hc3b25d78, 32'hc34e97a8, 32'h42f4e044},
  {32'h44f0b666, 32'h43a88cfd, 32'hc378eab7},
  {32'hc4015bc0, 32'hc4190e0e, 32'h43261d3e},
  {32'h434f17d4, 32'hc3948a22, 32'hc37bdc15},
  {32'hc4259874, 32'h42bd9b2e, 32'h42d43b27},
  {32'h44927ca3, 32'hc3519732, 32'h428bb66d},
  {32'hc50b9830, 32'hc039bb98, 32'hc3333810},
  {32'h44819f8d, 32'h43ea7f1f, 32'hc29ddc73},
  {32'hc485bf53, 32'h42a07465, 32'hc240b110},
  {32'h4466bf28, 32'h427f69bc, 32'hc3e820a1},
  {32'hc4adfc87, 32'hc2f99d66, 32'h41c523eb},
  {32'h43d6fc2a, 32'hc21164d9, 32'hc2a024a5},
  {32'hc4d32f8e, 32'h43260d37, 32'h4284c5d2},
  {32'h452413fe, 32'hc2ac874b, 32'hc38b0d68},
  {32'hc4cf52f8, 32'hc3ea10aa, 32'h431bbbe8},
  {32'h4524dd4a, 32'h428ee443, 32'hc35e8dd2},
  {32'hc40d0198, 32'hc24fc89a, 32'hc399913b},
  {32'h448a61d1, 32'h41647351, 32'h43381b0a},
  {32'hc41da610, 32'h428dca82, 32'h420f1630},
  {32'h44a2c5ce, 32'hc388377a, 32'h42edc030},
  {32'hc5074d77, 32'hc3d7cf1d, 32'hc29f800d},
  {32'h448e9cba, 32'h42a4b376, 32'h42d2e6ad},
  {32'hc411bc9c, 32'h40faf978, 32'hc3582d2e},
  {32'h4492dcf6, 32'hc3bd4fb9, 32'h4200f3e5},
  {32'h43c98498, 32'h42d04c64, 32'h43ab55d1},
  {32'h443cda26, 32'h4396993a, 32'hc3ce8fab},
  {32'hc51675b5, 32'h439d1771, 32'h3f991747},
  {32'h44c6de51, 32'h4317c2d6, 32'h43b33439},
  {32'hc41a0058, 32'hc3e9ccd3, 32'hc3475af0},
  {32'h44bc2c74, 32'h4293a9d8, 32'hc2fbe6f3},
  {32'hc507f09a, 32'hc237fc0d, 32'h4376a831},
  {32'h443df6a2, 32'hc22fd3c8, 32'h42379ae7},
  {32'hc4b0983f, 32'h4267b014, 32'h43f7e302},
  {32'h450fb7a0, 32'h439c07e3, 32'hc33e5cfb},
  {32'hc47f9388, 32'hc1256e14, 32'hc30a344a},
  {32'h44588a6e, 32'h42c642af, 32'hc3a23216},
  {32'hc4e8934a, 32'hc2c42810, 32'hc21c9f87},
  {32'h450d9671, 32'h419ff86b, 32'hc0df1f76},
  {32'hc4f8eb4e, 32'h43902bda, 32'h43912a37},
  {32'h44dbd1ce, 32'hc373c68d, 32'hc280fddc},
  {32'h4261f0e4, 32'h433b8fa8, 32'h431976e9},
  {32'h449ea67f, 32'hc2868a49, 32'h41f26d08},
  {32'hc50cb542, 32'hc215416f, 32'h42252648},
  {32'h450d2dd2, 32'h43ace916, 32'h4275478d},
  {32'hc3ad8db1, 32'hc30f2641, 32'h42ea6e1a},
  {32'h439e9a04, 32'hc2613907, 32'h42299eea},
  {32'hc490baaa, 32'h439b1077, 32'h4383a9ec},
  {32'h44459306, 32'h40be1731, 32'hc36e5dcb},
  {32'hc52e128e, 32'h4391ebd4, 32'hc285c52e},
  {32'h44b8d7ab, 32'h425e937b, 32'hc331548c},
  {32'hc4a902b9, 32'hc34a0010, 32'h43ae8153},
  {32'h44f24686, 32'hc3686d7f, 32'hc3a2da29},
  {32'hc4af9068, 32'hc32fa235, 32'hc14a6cc3},
  {32'h44f069be, 32'hc4481ee9, 32'h41ab9584},
  {32'hc4872854, 32'hc3b2bd81, 32'h417ec6be},
  {32'h45038dc5, 32'hc33bf12a, 32'hc2db28d6},
  {32'hc4604ce2, 32'hc391b744, 32'hc36402ef},
  {32'h44a568b5, 32'hc34c30f4, 32'hc3184616},
  {32'hc4a8007c, 32'hc18e764c, 32'hc35a6774},
  {32'h449c6532, 32'h4350dcb4, 32'hc10e6cfd},
  {32'hc41b8903, 32'hc300b465, 32'h43802a9b},
  {32'h44800d6a, 32'hc35d770e, 32'hc2c9e1f6},
  {32'hc482822a, 32'hc27687e8, 32'hc353a507},
  {32'h4519bda7, 32'h43da3865, 32'hc3ce3c59},
  {32'hc2ec64b5, 32'h42a7da2b, 32'h438e8b39},
  {32'h44344354, 32'h411c58be, 32'hc39f3e9c},
  {32'hc4ff1f67, 32'h4282ad91, 32'h439356e2},
  {32'h44f93db3, 32'h434a3be0, 32'hc3838d7f},
  {32'hc4f1c36c, 32'hc1ba313b, 32'hc31cfdfe},
  {32'h442ff5ec, 32'hc3698c0b, 32'hc3d00608},
  {32'hc4652b9c, 32'h43083f30, 32'hc1c18642},
  {32'h44f70c08, 32'h435e901b, 32'h432ad9c7},
  {32'hc4f85488, 32'hc3301d76, 32'h4360f741},
  {32'h44821479, 32'hc16e27d6, 32'hc352d6aa},
  {32'hc4738c6e, 32'h42c2475e, 32'h420066a1},
  {32'h44b38d86, 32'hc242cca3, 32'hc3cdb850},
  {32'h432fb3fb, 32'h414ea7d2, 32'h433ac3c5},
  {32'h4470fdc3, 32'h42a2a127, 32'hc3d4a7d5},
  {32'hc4f9fa72, 32'h4300f1d0, 32'h4108425a},
  {32'h43b191f4, 32'h42f30aa6, 32'hc2da5622},
  {32'hc4acf082, 32'hc32ee667, 32'hc361e553},
  {32'h44f27991, 32'h42fd6b47, 32'hc3790773},
  {32'hc3bf8340, 32'h4291e748, 32'h42ad560c},
  {32'h45228920, 32'h43174ada, 32'hc1e25f7b},
  {32'hc36105fa, 32'h434a411b, 32'h43d5966b},
  {32'h44c68633, 32'hc34bab5e, 32'hc309ac89},
  {32'hc3a3c6fa, 32'h42e7ba21, 32'h421e9e6c},
  {32'h44971a36, 32'h429670d7, 32'hc39a460f},
  {32'hc3641ccc, 32'h42d3690f, 32'hc2fbabe0},
  {32'h44e5fbb9, 32'hc3955f55, 32'hc283c5dc},
  {32'hc4f8de4b, 32'h43c6fb63, 32'hc2b7667e},
  {32'h43d18234, 32'h41d978ec, 32'hc2b1da0e},
  {32'hc49c6dbf, 32'h424219e9, 32'h434dfb80},
  {32'h43b01a3c, 32'hc3aacd9d, 32'hc2ad51d2},
  {32'hc4945cbe, 32'h4324ab58, 32'h4371e55b},
  {32'h44192db0, 32'h4328d3f7, 32'hc353033c},
  {32'hc4c6cc33, 32'hc33309a6, 32'h43a0539a},
  {32'h446107d0, 32'hc409d4eb, 32'hc4268e92},
  {32'hc49dbed4, 32'h436a78ba, 32'hc39afe07},
  {32'h435532a0, 32'hc353e860, 32'hc37d8cd7},
  {32'h44bff379, 32'hc2b794a4, 32'hc381c9bd},
  {32'hc4e0d20d, 32'h434e65b6, 32'hc3a1568e},
  {32'h44fa7bfb, 32'hc360df37, 32'hc30d7f21},
  {32'hc4a6b286, 32'hc384de26, 32'h42776a18},
  {32'h44317b7c, 32'hc38d979a, 32'hc30a02a2},
  {32'hc4bddc0f, 32'h431c9f3a, 32'h438ac720},
  {32'h4505fbaa, 32'hc39a4c09, 32'hc37b9565},
  {32'hc5029845, 32'hc1115166, 32'hc1ce650c},
  {32'h4376c760, 32'hc34631b6, 32'h4323ae7c},
  {32'hc4cf9056, 32'hc31f9afa, 32'hc2a6efe0},
  {32'h43f35da8, 32'hc3609565, 32'hc2d0c534},
  {32'hc506d40e, 32'h4086bfb2, 32'h430510c2},
  {32'h41ae8820, 32'h43a7c049, 32'h4342f239},
  {32'hc4c469bb, 32'h429e199d, 32'hc2cfaed3},
  {32'h43eaf6c0, 32'hc368fc37, 32'h41a2ad4c},
  {32'hc4b43757, 32'hc3e34df6, 32'h4272ce73},
  {32'h4455490a, 32'hc2137682, 32'h4353b4d6},
  {32'hc4cab5d0, 32'h41db3f8c, 32'h41612e5c},
  {32'h44f913eb, 32'h435013dd, 32'hc370f4cb},
  {32'hc3df10b9, 32'hc3a29aa3, 32'h42a030b7},
  {32'h44da1771, 32'h43ad6bfd, 32'h436e0618},
  {32'hc4e0e3c9, 32'h4343260b, 32'hc2a1eb2f},
  {32'h43c9e61c, 32'h420a21ef, 32'hc3099841},
  {32'hc4dd87e6, 32'hc23b1161, 32'h42623809},
  {32'h4509e396, 32'h426191a7, 32'hc3350ff0},
  {32'hc42d2ed2, 32'hc3727e14, 32'h4322cb8a},
  {32'h42f8be38, 32'h43754f7b, 32'hc3127517},
  {32'hc4f5f532, 32'hbfaaf048, 32'hc3307e86},
  {32'h42da75d0, 32'hc1a8cbf8, 32'h43835738},
  {32'hc50e5f4a, 32'h4309c233, 32'h43de07e1},
  {32'h43cdf9be, 32'h43872686, 32'hc3b9e230},
  {32'hc3fb9cf0, 32'h439f433e, 32'hc3a0818e},
  {32'h45029650, 32'h441d84de, 32'hc1d33550},
  {32'hc515ef59, 32'h433aec7c, 32'hc2826fc9},
  {32'h434b6e50, 32'hc313b8f1, 32'h421ae5cc},
  {32'hc50f9ce3, 32'hc3ad8b95, 32'h427fca4e},
  {32'h445af199, 32'hc39b5825, 32'hc201b8cc},
  {32'h432e18a0, 32'hc3e63761, 32'hc392e8ea},
  {32'h440e6c77, 32'h435fc81c, 32'h43bb5d29},
  {32'hc3b9b608, 32'h43065842, 32'h42ca119e},
  {32'h44b3d054, 32'hc3edb3ed, 32'h43777d9b},
  {32'hc3fe6625, 32'h4407a916, 32'h4404fa34},
  {32'h44b6de60, 32'hc243f9a3, 32'h40f82d21},
  {32'hc44edf7e, 32'hc33cae0f, 32'h4312e4d8},
  {32'h4505958a, 32'hc319eaab, 32'h439c24b0},
  {32'hc4dc5fb5, 32'hc425a271, 32'h43972b6a},
  {32'h449a7a8d, 32'h42cafbf9, 32'h404eb15e},
  {32'hc49ee123, 32'h430b035e, 32'hc2f17373},
  {32'h450a074d, 32'h425edee6, 32'hc3294765},
  {32'hc307c690, 32'h425ea1cf, 32'h4311cb44},
  {32'h44ac1eca, 32'h43e39327, 32'h436fecc8},
  {32'hc48509d0, 32'h40a5c10a, 32'h43cd9770},
  {32'h4480dcd4, 32'hc327f4e0, 32'h42b5fc22},
  {32'hc3df3008, 32'hc3493865, 32'hc1e80b85},
  {32'h44d1ca20, 32'hc394f0b8, 32'hc1d40f34},
  {32'hc3282190, 32'h437b9acc, 32'hc308c1d4},
  {32'h44eca360, 32'h41aa6f8f, 32'hc32eba2b},
  {32'hc44205ae, 32'hc32d5d28, 32'hc3384aa1},
  {32'h4501d346, 32'h4305f204, 32'hc1bd327e},
  {32'hc4f7a6c1, 32'h42b6aa19, 32'hc32a28f7},
  {32'h44aaa307, 32'hc37c7ec5, 32'hc22621e3},
  {32'hc4422f65, 32'h43d7f019, 32'h43af7e94},
  {32'h44f795a7, 32'h4147116e, 32'h435e8bfc},
  {32'hc483f0d8, 32'h41cc800d, 32'hc28e8cf9},
  {32'h4516c31b, 32'hc3ab6d2a, 32'h4385fde3},
  {32'hc4a3d02f, 32'hc39ede71, 32'h440d7778},
  {32'h44d27394, 32'h43887f7f, 32'h43ee82fa},
  {32'hc3dd330a, 32'hc307e854, 32'hc40a3493},
  {32'h42ca3970, 32'h41a5028f, 32'hc2657ae9},
  {32'hc41d62bb, 32'hc2075a5f, 32'h44085218},
  {32'h43eb3874, 32'hc3a0c073, 32'h4338992b},
  {32'hc4222e32, 32'hc308715f, 32'h4325e9d2},
  {32'h4527ecde, 32'hc31f0c64, 32'h4359faa9},
  {32'hc31a09c1, 32'h435c72c9, 32'h42115ef5},
  {32'h451441d2, 32'h4369b4fd, 32'hc1dd1edf},
  {32'hc4b603ac, 32'hc2f318c0, 32'h4290f659},
  {32'h4486475a, 32'hc3ac420e, 32'hc0bde84e},
  {32'hc4e118ab, 32'h438952a4, 32'hc38d7d6e},
  {32'h451d3858, 32'h440f13ba, 32'h431ca6d1},
  {32'hc4482120, 32'hc34445b8, 32'h43bc87fc},
  {32'h4427da37, 32'h42df3c76, 32'hc332631e},
  {32'hc3cfe03f, 32'hc3f9b7b3, 32'h437efe31},
  {32'h42b25c34, 32'h439351ed, 32'hc29b1c00},
  {32'hc4b87081, 32'hc2990811, 32'h4383efd0},
  {32'h446b564f, 32'hc2bf14a3, 32'h42ac5a63},
  {32'hc4e564fd, 32'hc1a29f12, 32'hc28fca6e},
  {32'h45142fbc, 32'h4346aaa9, 32'hc35375de},
  {32'hc4e34a1a, 32'hc0ea7c58, 32'hc32eb571},
  {32'h44fcb7c8, 32'hc2bfdc9f, 32'hc37bdf83},
  {32'hc5231274, 32'hc2cae2a6, 32'hc28b8010},
  {32'h4497290d, 32'h43e9a64a, 32'hc32fb23b},
  {32'hc3b17ee4, 32'h43c6fe7d, 32'h42b5b32d},
  {32'h4383884f, 32'hc374ab51, 32'h43a8c0c1},
  {32'hc3071b80, 32'hc16b904d, 32'h434e8400},
  {32'h44f8af20, 32'h413bdf5c, 32'hc34fc5b6},
  {32'hc4a49610, 32'h42b87425, 32'hc2baa8d5},
  {32'h4494c466, 32'hc287791d, 32'h43f8f5e4},
  {32'hc400182a, 32'h433c5ec8, 32'hc27b50e3},
  {32'h451d52af, 32'hc288584b, 32'hc27ceb9c},
  {32'hc4a418ed, 32'hc3370b53, 32'h4301ffad},
  {32'h451a442a, 32'hc385f898, 32'h435f17d9},
  {32'hc4af5dc9, 32'h43ff9a98, 32'h42e792be},
  {32'h45062ac5, 32'h43681435, 32'h44112c46},
  {32'hc4bed18f, 32'h4149ac19, 32'h43664d1a},
  {32'h445c5d4a, 32'h42f15ff5, 32'h410a896d},
  {32'hc4ba13bc, 32'h434f4131, 32'hc2eb5aea},
  {32'h449322ba, 32'hc3690b42, 32'h42fac530},
  {32'hc4182764, 32'hc2e985d9, 32'hc3074e60},
  {32'h44cef956, 32'h4210a2e2, 32'h429ae0e9},
  {32'hc3179510, 32'h431ec687, 32'hc3bc7e03},
  {32'h44864996, 32'h416b2e67, 32'hc2540235},
  {32'hc4b252fb, 32'hc3801401, 32'hc2690d73},
  {32'h4311c913, 32'hc42f30a2, 32'hbf367403},
  {32'hc506e50e, 32'hc363518c, 32'h42ae3d73},
  {32'h44ca55e3, 32'h41df63c4, 32'hc30b2d29},
  {32'hc202e440, 32'hc341938c, 32'hc2551b70},
  {32'h44ed2348, 32'hc2c82db6, 32'h43817e00},
  {32'hc49f9ff8, 32'h432c89a8, 32'h43e88381},
  {32'h45073771, 32'hc322baa5, 32'h438b7649},
  {32'hc5035269, 32'hc3be29e6, 32'h4228e5e8},
  {32'h43147b10, 32'hc3cffed1, 32'h438f71ba},
  {32'hc48531a9, 32'hc3adaeb8, 32'hc2501eb6},
  {32'h4485063c, 32'hc325cc66, 32'hc3902de7},
  {32'hc491c45a, 32'hbf97dea0, 32'hc05d9950},
  {32'h44832be0, 32'hc29b9677, 32'hc2a64ba6},
  {32'hc47b4c18, 32'h42fb9877, 32'hc30b8982},
  {32'h44a31c22, 32'h438351d6, 32'h43a7cea3},
  {32'hc32327a0, 32'hc187ca57, 32'h4240fc03},
  {32'hc2d96608, 32'h43bfcee3, 32'h43333780},
  {32'hc494cf9d, 32'h41a401e5, 32'h4379b90d},
  {32'h4506f261, 32'hc3b0ddd1, 32'hc2a5a27c},
  {32'hc4884a5c, 32'hc2da4ca7, 32'hc1a23cf5},
  {32'h44d94268, 32'h43f41970, 32'h433996ed},
  {32'hc41936fa, 32'h43090d0c, 32'h41a9bd5e},
  {32'h44b2bea2, 32'hc22c080f, 32'h42b7a094},
  {32'hc4e23cf9, 32'h431d1d3d, 32'h4357ee38},
  {32'h44ba5779, 32'h4395ef14, 32'h430392aa},
  {32'hc4f24e0c, 32'h4399ec6d, 32'h437b56c2},
  {32'h44efc9ca, 32'hc1c7f758, 32'hc28d4b17},
  {32'hc48348a0, 32'hc2ab1d63, 32'hc09703f4},
  {32'h44ca4af3, 32'h433f50f4, 32'hc31bb63c},
  {32'hc43da643, 32'h4400bafa, 32'hc39fe625},
  {32'h44cd131e, 32'hc3562d64, 32'h42bf967a},
  {32'hc46940ce, 32'h4382ae52, 32'hc3267abd},
  {32'h44ad93ca, 32'hc309bd56, 32'hc30222e7},
  {32'hc45b2c69, 32'h4284ce56, 32'h42a25e4e},
  {32'h44c5badc, 32'hc29ec360, 32'hc17cc77a},
  {32'hc4c00b87, 32'h43b2ef62, 32'hbff99bb0},
  {32'h449a0082, 32'h41e748ac, 32'h4241c805},
  {32'hc47b1870, 32'hc287ee68, 32'h426f5df5},
  {32'h44aa64a9, 32'hc1b8ec7d, 32'hc2e147fc},
  {32'hc50afdf8, 32'h43a7ce2f, 32'h43c427e3},
  {32'h4426b23b, 32'h435ab23e, 32'hc22a087f},
  {32'hc4fe4f38, 32'hc2ba2249, 32'hc3a7e33c},
  {32'h43fb498c, 32'hc3516084, 32'hc319846e},
  {32'hc43a3068, 32'h431d9cf5, 32'h42a66aac},
  {32'h4488edf3, 32'hc26fdd81, 32'h41f79148},
  {32'hc42ff83e, 32'h43abce85, 32'h43018a51},
  {32'h45065690, 32'hc3ae222a, 32'hc4096076},
  {32'hc49bbd3d, 32'hc2f03109, 32'h42ad8050},
  {32'h45005fcf, 32'h43d82ce7, 32'hc228d258},
  {32'hc46da30c, 32'hc3e713ee, 32'h42d25ef7},
  {32'h43f03f80, 32'hc35df37e, 32'hc308ee1e},
  {32'hc25f5650, 32'hc1c6122c, 32'h4283e0dc},
  {32'h44de4116, 32'h4156ef47, 32'h41016c72},
  {32'hc4bc0b47, 32'hc3fc24fe, 32'hc1c4426e},
  {32'h44ee3d5c, 32'hc26ca606, 32'hc2ad4e9a},
  {32'hc3502200, 32'hc2fed6d7, 32'hc309f918},
  {32'h45115c86, 32'hc38c97b1, 32'h428d3907},
  {32'hc473c9f4, 32'h4235abe5, 32'hc25ea7a6},
  {32'h443c947d, 32'hc28b6bd3, 32'h408be75c},
  {32'hc4893dc2, 32'h43a07070, 32'h438255f4},
  {32'h441f025a, 32'h4290c0f0, 32'hc1b99ce6},
  {32'hc41afc3e, 32'hc329999c, 32'h43708d41},
  {32'hc38f9a74, 32'h43395f3b, 32'h42b6c668},
  {32'hc4dd0e80, 32'hc33c124d, 32'hc1844935},
  {32'h43a9c0c0, 32'hc0d15902, 32'hc37e9381},
  {32'hc4e9fea2, 32'h43241cd3, 32'h43327155},
  {32'h450dfc4b, 32'hc39b070d, 32'h41444f33},
  {32'hc40f622c, 32'hc2330929, 32'hc0c080f2},
  {32'h43a96668, 32'h429676c9, 32'h426a94ca},
  {32'hc4452aae, 32'h416dc693, 32'h4314ea07},
  {32'h444c42c9, 32'h428c5137, 32'hc38fbaf2},
  {32'hc432196c, 32'h439c3bce, 32'h42f0db5f},
  {32'h4442f38a, 32'h41ee886d, 32'h4234664b},
  {32'hc43ebb0a, 32'h42cdf22b, 32'h42c61746},
  {32'h4473dca3, 32'h430ab17c, 32'hc235111f},
  {32'hc4a7143b, 32'hc32836b9, 32'hbfcbb602},
  {32'h44d18b83, 32'hc0f50dd4, 32'hc351e922},
  {32'h428803be, 32'hc1ee1fb4, 32'h430decbf},
  {32'h451ab0cc, 32'hc2ce9781, 32'h43a945f4},
  {32'hc4bad9af, 32'h43dff944, 32'h437acfc2},
  {32'h45042bfd, 32'h43277d8c, 32'h416330e8},
  {32'hc50673a0, 32'h420d7801, 32'hc31d14a4},
  {32'h43bf7e5c, 32'hc37244ca, 32'h42c3de0e},
  {32'hc4e0d356, 32'hc1d2058d, 32'hc311731a},
  {32'h44a1c27f, 32'hc299277a, 32'hc2a16660},
  {32'hc4f3a2d1, 32'hc299fa9b, 32'hc20a2dac},
  {32'h44234519, 32'hc126db91, 32'h429bf22f},
  {32'hc47de25b, 32'h429fc2eb, 32'hc27aa4cd},
  {32'hc223da80, 32'h434a2c19, 32'h42c5087c},
  {32'hc4e47617, 32'h42ab8e88, 32'h427ec122},
  {32'h42a1311c, 32'hc3873663, 32'h42694469},
  {32'hc45bc030, 32'hc3046857, 32'h422c91b8},
  {32'h447d22bc, 32'hc341a732, 32'hc377062b},
  {32'hc4e6c397, 32'h4423cf45, 32'h433d5ca4},
  {32'h44c66c5b, 32'hc3ccdb06, 32'h43259767},
  {32'hc4bcc6af, 32'hc334fe0d, 32'h42c3a3d2},
  {32'h44def70c, 32'hc398e92c, 32'h41a6de3a},
  {32'hc4d20df2, 32'h42b293cd, 32'h4401bdbf},
  {32'h442a0516, 32'hc2a71d04, 32'hc20782d0},
  {32'hc34bf697, 32'hc2634fba, 32'h4334a9ee},
  {32'h450a7cb9, 32'h433905de, 32'hc2dbdf72},
  {32'hc43414d8, 32'hc40ec90d, 32'hc2a35ba1},
  {32'h448dd35d, 32'h4343d6ec, 32'h424dd562},
  {32'hc4861790, 32'h43ab48e6, 32'h4215a0b5},
  {32'h44ae097c, 32'hc34904c5, 32'h427fec47},
  {32'hc50b1a3d, 32'h427172ea, 32'h433c868a},
  {32'h447df473, 32'hc40e6b7f, 32'h438b7920},
  {32'hc469b6f7, 32'h42842d24, 32'h437a61ba},
  {32'h44ee71ca, 32'h401b8262, 32'hc38d7c11},
  {32'hc48022ad, 32'h435ab541, 32'hc2fd38e7},
  {32'h43563b08, 32'hc1a8be0a, 32'hc34da801},
  {32'hc4dc9896, 32'hc24aaea7, 32'hc3baaa4c},
  {32'h43bcbc10, 32'hc38038f6, 32'hc3a51975},
  {32'hc430b28a, 32'h42e6babd, 32'h413a6c1b},
  {32'h44827dfc, 32'hc3773c53, 32'h41bf91fb},
  {32'hc4960cca, 32'h43b4638e, 32'hc3182917},
  {32'h44b40a9a, 32'h4283d80a, 32'hc3819379},
  {32'hc4057e9e, 32'h43542a40, 32'hc2837daf},
  {32'h44dadcf9, 32'h428394e5, 32'hc3a71df4},
  {32'hc507dd1a, 32'hc2971f6d, 32'h4350b586},
  {32'h44c794b7, 32'hc2f8819f, 32'h4269e6df},
  {32'hc4a5cc3e, 32'hc2b82bc9, 32'h433333e5},
  {32'h45087cfc, 32'h4337af64, 32'h4310b9b7},
  {32'hc41656a7, 32'hc372b922, 32'hc3179a19},
  {32'h442994b6, 32'h43be0a0d, 32'hc2eafa23},
  {32'hc40529e8, 32'hc1fa94a5, 32'h42d4a6f0},
  {32'h44837b0f, 32'hc229cbc7, 32'h43d34a02},
  {32'hc49e699a, 32'hc2cbbf85, 32'h423d335d},
  {32'h441f6998, 32'h426e3b4c, 32'hc2d65f96},
  {32'h4391ea58, 32'h42a709c9, 32'hc30b6306},
  {32'h44ac699d, 32'h419f39b5, 32'h42f21eba},
  {32'hc4b916bd, 32'h42e9a78e, 32'h43bbd921},
  {32'h44e8178e, 32'hc3a2e8f4, 32'hc256308c},
  {32'hc506c0b7, 32'h43537993, 32'hc2389b50},
  {32'h4412eecc, 32'hc2b759fb, 32'h4381cd70},
  {32'hc4a0c9e4, 32'hc3b02ba0, 32'h42b1e9b8},
  {32'h44b1a78d, 32'hc2353f59, 32'hc35f2e6c},
  {32'hc3ab6e4c, 32'h42cb3a2a, 32'hc3414b39},
  {32'h44c01da4, 32'h42c82b2e, 32'hc18c36e6},
  {32'hc4e782ba, 32'hc241934c, 32'hc3579fdf},
  {32'h44fe3e52, 32'hc3558ad4, 32'h4081993c},
  {32'hc4afe1d0, 32'hc2df899a, 32'hc2d62d43},
  {32'hc335d8a8, 32'h42fe1a62, 32'hc2ab7398},
  {32'hc3bcfcc0, 32'h42253a16, 32'hc400b24f},
  {32'h44d4e66f, 32'hc310e326, 32'h438d3c97},
  {32'hc1f17480, 32'h438aca3c, 32'h43ed5f8b},
  {32'h4442824a, 32'h43299baf, 32'h43291599},
  {32'hc4ef5358, 32'h420e846a, 32'hc3009109},
  {32'h447ab400, 32'h43df3cbd, 32'hc32ccb9a},
  {32'hc475ab11, 32'hc35af773, 32'hc344d78a},
  {32'h45163514, 32'h42a31640, 32'hc3abeca7},
  {32'hc45aa306, 32'hc3e36df3, 32'h44117f24},
  {32'h4516ef50, 32'h42a494b3, 32'hc3dbb724},
  {32'hc3eed3d4, 32'hc0522504, 32'h43466e77},
  {32'h4481c16d, 32'hc375d74e, 32'hc39f8a21},
  {32'hc3c276f0, 32'h442d1414, 32'hc26d54d0},
  {32'h44f78262, 32'h4372c819, 32'h42995c96},
  {32'hc4311820, 32'hc343463a, 32'hc2eb4d4c},
  {32'h451e85b8, 32'h42d2bdd1, 32'h4303caa8},
  {32'hc3fec0e0, 32'h42ee01b3, 32'hc225ed3b},
  {32'h452c19f0, 32'hc403af61, 32'hc373f2e5},
  {32'hc4950f67, 32'hc3591f9c, 32'hc3c8aa09},
  {32'h44b922f8, 32'hc3760277, 32'h430f75e4},
  {32'hc4fa7f37, 32'hc349c3cc, 32'h4368e643},
  {32'h4303700c, 32'hc389d8b9, 32'hc3aa38b9},
  {32'hc3341701, 32'hc245c8a8, 32'hc2a552fc},
  {32'h44ee9375, 32'hc32626c1, 32'h41e4ca1a},
  {32'hc45cae22, 32'h42ea6c9a, 32'h418fd7a2},
  {32'h44e84054, 32'h4174d4e4, 32'hc3528877},
  {32'hc4b3e6f8, 32'h43d3dbf8, 32'hc3a94795},
  {32'h44bdab94, 32'hc2558f90, 32'h42f82148},
  {32'hc508e35d, 32'h43cb0023, 32'hc290c2e4},
  {32'h449d3849, 32'hc2a30f1a, 32'h41cb1328},
  {32'hc4c15847, 32'hc32bb95b, 32'hc34a8f96},
  {32'h43da1e56, 32'hc282dfb5, 32'h432c532d},
  {32'h4327a98e, 32'hc2bf3cf1, 32'hc1a7e4a7},
  {32'h43b17c70, 32'hc2f183b2, 32'hc296450a},
  {32'hc4bb8d5f, 32'h422236b7, 32'hc3b5ba8b},
  {32'h44db6dce, 32'hc3bd419b, 32'h436b0f11},
  {32'hc48c585d, 32'hc2901ef8, 32'h43a85ab0},
  {32'h448e70c5, 32'h430844e5, 32'h42b8b298},
  {32'hc43de6dd, 32'h43979db4, 32'hc2831a4c},
  {32'h44d5d3c9, 32'hc3182f86, 32'hc33edbbb},
  {32'hc508fb90, 32'h434ed151, 32'hc2386cc8},
  {32'h4505a21b, 32'h439c3b5a, 32'h43a8b0c4},
  {32'hc3f93958, 32'h43b1d7fc, 32'h4316c864},
  {32'h43469698, 32'hc1b91b2f, 32'hc3801c1b},
  {32'hc3ec7d34, 32'hc3993066, 32'hc32f5416},
  {32'h450575b2, 32'hc3739696, 32'h426772e4},
  {32'hc3c75f57, 32'h43114379, 32'hc39abb79},
  {32'h42f63010, 32'hc34bb722, 32'h4346cf23},
  {32'hc4072a14, 32'h42134f91, 32'hc25f136f},
  {32'h45171897, 32'hc30812dc, 32'hc113d0bc},
  {32'hc501e788, 32'hc401e6fb, 32'h429e34a3},
  {32'h445ca51e, 32'h425623c0, 32'h4157afbb},
  {32'hc3310c5c, 32'hc32d67f6, 32'h43497f58},
  {32'h451bc9d5, 32'hc28990bd, 32'h42afde4a},
  {32'hc3edd7fc, 32'h4331256c, 32'h42d01a0a},
  {32'h43d4db4d, 32'hc3ba596c, 32'hc21260b4},
  {32'hc5016ab0, 32'h421c8aea, 32'hc3109d50},
  {32'h44bcde94, 32'h43880e87, 32'h42eeb96f},
  {32'hc47dff8e, 32'hc2c93eb7, 32'hc301bca6},
  {32'h44c57021, 32'hc260c8f4, 32'hc36cf17d},
  {32'hc4919103, 32'h431c3f3f, 32'hc27f1db9},
  {32'h44fd4a1f, 32'h435092d2, 32'hc34a286b},
  {32'hc4b95dc2, 32'hc1caddd1, 32'hc3da4178},
  {32'h440fd21a, 32'hc110f4c1, 32'h431ef1e2},
  {32'hc501ba44, 32'h43b8baea, 32'hc3c4338e},
  {32'h44fa813b, 32'h4374d0d0, 32'h42ad7384},
  {32'hc29b3140, 32'hc31992d4, 32'h42e4e070},
  {32'h450ddddd, 32'hc20a8448, 32'hc2eb6f39},
  {32'h42b65320, 32'hc310b4fb, 32'h43a88cc7},
  {32'h44d25752, 32'hc317df9b, 32'hc2639e8c},
  {32'hc4a9bb29, 32'hc2ea093c, 32'h4307695a},
  {32'h45087ad8, 32'h41ef8ec9, 32'h43bf83ce},
  {32'hc5210a77, 32'hc2bc0949, 32'h43d0e6b2},
  {32'h44b25e01, 32'hc36853a4, 32'h4340f8ef},
  {32'hc4c99399, 32'hc28e1ed6, 32'h4318ee22},
  {32'h44a6e416, 32'h4294cc9c, 32'hc313e5ed},
  {32'hc4862c33, 32'h431e6791, 32'h42b7015d},
  {32'h4406fc3a, 32'hc34050c8, 32'hc2a9acdc},
  {32'hc4d9e519, 32'h42d4ed8f, 32'h43b9647f},
  {32'h44aa7c0d, 32'hc23ccf5f, 32'h4327840a},
  {32'hc47a71d0, 32'h42dd5316, 32'hc3051413},
  {32'h440864d7, 32'hc3087085, 32'h43947c99},
  {32'hc4d0273c, 32'h42bd91a0, 32'hc30a27f0},
  {32'h44d35a0e, 32'hc339df2d, 32'h430fef20},
  {32'hc456e02b, 32'hc3186f30, 32'h42246dd7},
  {32'h44b5c4b2, 32'h4374d802, 32'hc20eb739},
  {32'hc35e88e4, 32'hc32df265, 32'hc3befa9e},
  {32'h43b53ef0, 32'h42213311, 32'hc2b7675b},
  {32'h43041530, 32'h41b3e940, 32'hc1fa502a},
  {32'h449cb285, 32'h420087b6, 32'hc3708a49},
  {32'hc4fed9d3, 32'h436220d4, 32'hc3af64d8},
  {32'h43e4d0d8, 32'h42e98422, 32'hc2c0e953},
  {32'hc51030b8, 32'hc269ba97, 32'hc304d62f},
  {32'h44f61a03, 32'hc14648a0, 32'h4406778a},
  {32'h41e76f80, 32'h41e75592, 32'h426cc83e},
  {32'h448a60b8, 32'hc28ca8ae, 32'hc3488a45},
  {32'hc428586f, 32'hc3adaefe, 32'h434079f6},
  {32'h449a2f6c, 32'h41bfec33, 32'hc33acbfa},
  {32'hc3cd9308, 32'hc3ad0ee6, 32'hc30cf654},
  {32'h441a9312, 32'hc3a4e45f, 32'hc2e7ac63},
  {32'hc4660d24, 32'hc2cb1f40, 32'h429bca8b},
  {32'h43ec058c, 32'hc35dffb5, 32'h42d9d831},
  {32'hc4285232, 32'hc3befb5d, 32'h438f6273},
  {32'h44bc4479, 32'hc3107399, 32'hc1ce4aca},
  {32'hc4166cf9, 32'hc29cd16c, 32'h431c3189},
  {32'h44764c7d, 32'hc2cd9fae, 32'hc2d0e7f9},
  {32'hc50f3843, 32'h439c2df9, 32'h438bba50},
  {32'h44c239bc, 32'hc1af1d81, 32'h42b2e8bb},
  {32'hc4bc69c8, 32'h42123c5f, 32'h43daf2f0},
  {32'h43f384d4, 32'hc4198a7e, 32'hc33d2f44},
  {32'hc3d17218, 32'h43dfe5e4, 32'hc35573eb},
  {32'h44125f21, 32'h42cc1673, 32'hc40ca592},
  {32'hc4ceb083, 32'h43481daf, 32'h44217f91},
  {32'h45200db7, 32'h4188be32, 32'hc3394831},
  {32'hc50880e9, 32'hc31c2a32, 32'hc3092f8a},
  {32'h4412fe2a, 32'h43461f1e, 32'hc357eb98},
  {32'hc481c0c4, 32'h4294f11e, 32'h43c005ca},
  {32'h4431b914, 32'h4297bbdc, 32'h43b92b3e},
  {32'hc4ba52b2, 32'hc3e791a4, 32'h4390b97f},
  {32'h441b4a34, 32'h438b82c2, 32'hc34bd88c},
  {32'hc512221c, 32'h431d6d71, 32'h431851d1},
  {32'h448488aa, 32'hc21d95d9, 32'hc21ea17d},
  {32'hc490a4db, 32'hc36b9bb9, 32'h432efe59},
  {32'h448b127c, 32'h4333b9ad, 32'h42c70732},
  {32'hc507b542, 32'hbf959a8e, 32'hc272c8bf},
  {32'h4474f63f, 32'h426e6db6, 32'hc304c1a8},
  {32'hc4547bed, 32'h4327e5e4, 32'h43a4c655},
  {32'h4238a2b0, 32'h43bc9f01, 32'h430b82d2},
  {32'hc50ec16b, 32'hc3106eed, 32'hc28b6f8c},
  {32'h449bae53, 32'hc2a8f5ac, 32'h432614b0},
  {32'hc50cf425, 32'h43303e4d, 32'hc3c4e7ca},
  {32'h448b682d, 32'hc2861efb, 32'h4349603a},
  {32'hc5102341, 32'hc39f8671, 32'h4356ca5d},
  {32'h4466256d, 32'h42907fb8, 32'hbdd9f660},
  {32'hc4b950af, 32'h43c0b99b, 32'hbfc0a0b0},
  {32'hc2817470, 32'hc366b488, 32'h43b1e350},
  {32'hc3e38a18, 32'h40426eb0, 32'h4257b0bd},
  {32'h4411f9a8, 32'hc366f254, 32'hc3b6c174},
  {32'hc4a1f9f1, 32'h429d866c, 32'hc08a35a8},
  {32'h44b509a7, 32'h428d18f5, 32'h4395e148},
  {32'hc4166850, 32'hc3d9d5ae, 32'h43821646},
  {32'h44ab322e, 32'h41a2042f, 32'h42e607f9},
  {32'h42d087c4, 32'h4337667c, 32'hc183d750},
  {32'h43965b30, 32'hc30ae8aa, 32'h429604b1},
  {32'hc519fc9a, 32'h438f9a37, 32'hc3e43590},
  {32'h44b55cc7, 32'hc2d58bc5, 32'h419c3f2a},
  {32'hc296c860, 32'h438a82c2, 32'hc3544840},
  {32'h44e16cb1, 32'hc0dd173a, 32'h42a0e672},
  {32'hc4a23ef4, 32'h432890fd, 32'h43c79e30},
  {32'h4312d020, 32'hc2d2a94a, 32'h436464d2},
  {32'hc347ae3e, 32'h432fb4e5, 32'hc2b7e368},
  {32'h4516e7dd, 32'h40b6372d, 32'hc32345f1},
  {32'h4325b71e, 32'h4189f193, 32'hc21add26},
  {32'h44b267ef, 32'h4339781e, 32'h41f8b824},
  {32'hc2dceee0, 32'h418d6750, 32'h42c29c4c},
  {32'h44ee6da8, 32'h431571ce, 32'hc2c8ad21},
  {32'hc438e01e, 32'h43fa7067, 32'hc37155a8},
  {32'h4449b488, 32'hc2bbde7a, 32'hc3bb60c1},
  {32'hc4c81746, 32'h439cc05e, 32'h42ee14de},
  {32'h451576ad, 32'h418bcb66, 32'h43020a0b},
  {32'hc40c04cc, 32'h420bf3f3, 32'h438a44b8},
  {32'h44ad411e, 32'h42beba17, 32'hc2327381},
  {32'hc49e643c, 32'hc29b896d, 32'h4238c21a},
  {32'h44013dcc, 32'h43b256ea, 32'h43138f26},
  {32'hc49af78d, 32'h41ed39fc, 32'hc24e4bfb},
  {32'h44fb3f3a, 32'hc3a518a4, 32'h439917b3},
  {32'hc4384116, 32'h416382e4, 32'hc1d81eb8},
  {32'h44de31d8, 32'hc28c886b, 32'hc22e40a1},
  {32'hc48fb598, 32'h41e488e1, 32'hc418703b},
  {32'h44690e5c, 32'h43605559, 32'hc2e72c3c},
  {32'hc34b0c28, 32'hc01b7ced, 32'hc318f8e7},
  {32'h44f14bb8, 32'h4200ca4e, 32'hc332e9c2},
  {32'hc411034f, 32'h42467617, 32'hc35aa78b},
  {32'h439b5160, 32'hc2b05245, 32'h4323a792},
  {32'hc4da0aac, 32'h43939a8e, 32'hc3a90b69},
  {32'h450ce50a, 32'h438da4ee, 32'h43abe23a},
  {32'hc4e7300e, 32'hc3dc27f9, 32'hc3abb3c8},
  {32'hc3375c00, 32'h43069fdf, 32'hc32a3393},
  {32'h450b3502, 32'h42c605b7, 32'h434fecc0},
  {32'hc4714121, 32'hc2e8f6d1, 32'hc40c7233},
  {32'h43755100, 32'h42fe0d37, 32'h42b12a18},
  {32'h42868d38, 32'h429d3164, 32'h42d60f91},
  {32'h450b0f24, 32'hc3bb5271, 32'h430df470},
  {32'hc459c93a, 32'hc2250b72, 32'hc39c0aa4},
  {32'h451983a8, 32'h423270df, 32'h432b6d85},
  {32'hc49bc9f8, 32'hc36a37e2, 32'hc382385b},
  {32'h44eca243, 32'hc3895c73, 32'h426e8cbd},
  {32'hc4b82970, 32'h41738b7d, 32'hc11ac9aa},
  {32'h44b32a24, 32'hc38e1bad, 32'h43cccca2},
  {32'hc50d1896, 32'h43060e21, 32'h41c1beea},
  {32'h44674998, 32'h43dc0c51, 32'hc313d79b},
  {32'hc49efb59, 32'hc3a9b628, 32'h43902657},
  {32'h44c2f6d1, 32'h431ad8ee, 32'h43530d80},
  {32'hc43be0e1, 32'h42f9a5b7, 32'hc2c7873b},
  {32'h4504e4dd, 32'hc173212f, 32'hc32ef76d},
  {32'hc4603736, 32'hc371b125, 32'hc2a8b856},
  {32'h4382bb5e, 32'hc373cd6b, 32'h42ec1b60},
  {32'hc4ac42f0, 32'h43847a09, 32'hc3c1ac86},
  {32'h44892fbf, 32'hc1b10670, 32'h433cd077},
  {32'hc50268b2, 32'h42cd26c6, 32'h4323dd3c},
  {32'h44de24d0, 32'h438302d9, 32'h4238e51d},
  {32'hc3abe160, 32'hc2c60a9c, 32'hc310ae99},
  {32'h449950e6, 32'h438f1251, 32'h43321b77},
  {32'hc4bde94a, 32'hc1f23796, 32'h42781ce1},
  {32'h449536fd, 32'h432c613e, 32'h439ecb78},
  {32'hc4385de5, 32'h435198e8, 32'hc3943fde},
  {32'h4488f995, 32'h43a56e91, 32'h43769a76},
  {32'hc4f0d178, 32'h434d79fc, 32'hc2203422},
  {32'h444bdb49, 32'hc3092115, 32'h42f73edb},
  {32'hc3b40c27, 32'h4344c965, 32'h42f2e67b},
  {32'h44b1b885, 32'hc2822f06, 32'h43bcffd5},
  {32'hc4e7afd4, 32'h42f8dd6b, 32'hc23c139d},
  {32'h44f78ae7, 32'h41ca1fea, 32'hc2a0dd24},
  {32'hc4bc8116, 32'hc15e4c4d, 32'h4294ee55},
  {32'h44658484, 32'h43baddc7, 32'h432598b2},
  {32'hc428e944, 32'hc2500075, 32'hc23c5015},
  {32'h44cc7d27, 32'hc26fa37c, 32'h420d7c9c},
  {32'hc48eae17, 32'hc36886e3, 32'hc374e413},
  {32'h43f2369c, 32'hc2e5c19f, 32'hc1ce8f79},
  {32'hc3e2c127, 32'h42756f6b, 32'h42b5870e},
  {32'h43aa6fbf, 32'h43b5cd03, 32'h43c89c29},
  {32'hc4a29287, 32'h4328b57e, 32'hc3b260ba},
  {32'h4519ec1c, 32'h43202e32, 32'h436444d2},
  {32'hc3ae561e, 32'h42617732, 32'h4234e68e},
  {32'h44d75051, 32'hc28dee50, 32'h42f55422},
  {32'hc3aed7a4, 32'h44059b1b, 32'h436b8f34},
  {32'hc38ca77c, 32'h42cbfb4d, 32'h43fd629f},
  {32'hc4ad2066, 32'hc2e82b45, 32'h40ba162e},
  {32'h44f0de88, 32'hc05ba020, 32'h42e26778},
  {32'hc4940940, 32'h435c7e7d, 32'hc3b9823c},
  {32'h440ba67c, 32'h42b107a0, 32'h42e35134},
  {32'h43061455, 32'hc1ebe77c, 32'h41c13b2c},
  {32'h450dcb15, 32'hc2a20f3a, 32'hc3775d8e},
  {32'hc24a6a80, 32'h43bf4f36, 32'h41590bfc},
  {32'h4452d93e, 32'h4311a0d6, 32'hc2fa8736},
  {32'hc499951e, 32'h4387ea2c, 32'hc38a7adf},
  {32'h45059fa1, 32'h42259879, 32'h424cc3d9},
  {32'hc4e1bccc, 32'hc284b22c, 32'h435476a7},
  {32'h44151426, 32'h42b1bf30, 32'hc3d11551},
  {32'hc4ba712e, 32'h4292d598, 32'h41e0a74c},
  {32'h446124b5, 32'hc38e034b, 32'hc25cf3cf},
  {32'hc42df5c8, 32'h4352ac52, 32'h439a91ec},
  {32'h4437f740, 32'h438c4be4, 32'h43a1f423},
  {32'hc47e3f96, 32'h42fc688b, 32'hc101ee5e},
  {32'h4411f938, 32'hc2edf022, 32'hc3ac07e8},
  {32'hc41dae18, 32'h420aad9d, 32'h4361da79},
  {32'h4481c18b, 32'hc3831605, 32'hc3d7b007},
  {32'hc4a12bfb, 32'h4403631a, 32'h4283761c},
  {32'h417e6e80, 32'hc3477d9c, 32'h432a9690},
  {32'h42cdc651, 32'hc3bd34f2, 32'hc38f66f5},
  {32'h451b49af, 32'hc1e7cb13, 32'h41ef6352},
  {32'h4136b980, 32'hc1c7fbc9, 32'h43275264},
  {32'h44cb6154, 32'h437b7c41, 32'h434f17e5},
  {32'hc47b2da6, 32'hc3abb82e, 32'hc294a994},
  {32'h44f840fc, 32'h43e9ccea, 32'h43753084},
  {32'hc512bc6a, 32'hc1c19707, 32'hc34f0b45},
  {32'h440a90e2, 32'h436f4bc5, 32'h43241fb0},
  {32'hc3ef434a, 32'hc401ca7b, 32'hc2ceb571},
  {32'h44709e6a, 32'hc37b768a, 32'hc22ff6b5},
  {32'hc4a2371b, 32'h43685fe2, 32'h433efd50},
  {32'h44df06d5, 32'h42c5265f, 32'h409e1cce},
  {32'hc3e72050, 32'hc2a9ccd4, 32'hc3988e90},
  {32'h451f3a2d, 32'hc365e41a, 32'hc2600da3},
  {32'hc5088137, 32'hc24c6f9a, 32'hc36dce50},
  {32'h43e02d00, 32'h43c17a16, 32'hc27c404a},
  {32'hc50e5ab6, 32'h44076d11, 32'hc20e9901},
  {32'h44b97983, 32'hc2907293, 32'h43650f1b},
  {32'hc4a5c962, 32'h430fd389, 32'hc3a88e6f},
  {32'h446348f5, 32'h426177ed, 32'hc3096289},
  {32'hc345bdd6, 32'h438bfc41, 32'hc3edd8be},
  {32'h42919380, 32'hc0b71348, 32'h42e79662},
  {32'hc4a46037, 32'h43ad796d, 32'h438b0f57},
  {32'h428ef185, 32'hc3b331a2, 32'h43a5b79d},
  {32'hc2a3a000, 32'hc2ac9b15, 32'h430e73f6},
  {32'h444eabb4, 32'hc3127ada, 32'hc3e3bb57},
  {32'hc4aac485, 32'hc3080f00, 32'h4201412f},
  {32'h4522b0c4, 32'hc2dddf6e, 32'h42a8fcdc},
  {32'hc50281d6, 32'h433b9e1e, 32'h42c7e2ae},
  {32'h40afd800, 32'h42f4d347, 32'hc18f060e},
  {32'hc470d8f3, 32'hc3cd8c30, 32'hc397c3c1},
  {32'h43929fc4, 32'hc267ebbc, 32'h44034724},
  {32'hc4bdaf19, 32'h42c4b8ec, 32'h43f0b39e},
  {32'hc33acfb6, 32'hc39d2140, 32'hc31a6a67},
  {32'hc4a079ae, 32'h4392858c, 32'h4219d083},
  {32'h4369b360, 32'hc3a51fb2, 32'h43a371e1},
  {32'hc4a7340e, 32'h438cb683, 32'h42a4caca},
  {32'h45128354, 32'h436ea5be, 32'hc38a1ae2},
  {32'hc3f12336, 32'hc32dec74, 32'hc1d97c6a},
  {32'hc2913c88, 32'h43cc1684, 32'hc35af260},
  {32'hc488f353, 32'h42ce6ed3, 32'h43332ddc},
  {32'h44fdf1e8, 32'hc261f00e, 32'hc3335914},
  {32'hc45d6ca2, 32'h43d1a3e5, 32'h436a56da},
  {32'h4509c5b5, 32'hc1fe3e08, 32'hc407dabf},
  {32'hc405f780, 32'hc40b3945, 32'h4322fff9},
  {32'h44c9d298, 32'hc3934491, 32'h42828ea3},
  {32'hc4b1efa6, 32'h42ed0451, 32'h41ac9bc9},
  {32'hbead5000, 32'hc3427a99, 32'h439627aa},
  {32'hc40de530, 32'h42dda617, 32'hc1da8c19},
  {32'h444ff162, 32'h42904484, 32'hc19c3cbc},
  {32'h41e3ee00, 32'h414457c1, 32'h432696b5},
  {32'h4401d300, 32'hc3752293, 32'hc2bd861b},
  {32'hc4195002, 32'h42d5428d, 32'h3ebc70a0},
  {32'h43b7b438, 32'h422431d0, 32'h440d6522},
  {32'hc3e60890, 32'hc3447b3e, 32'h432b878a},
  {32'h450c0d7a, 32'h4157da92, 32'h433d1e2e},
  {32'hc50ab025, 32'hc28a6ba9, 32'hc3a6c632},
  {32'h445e6f2a, 32'h433aab94, 32'hc2c88550},
  {32'hc4dfa06e, 32'h4395f0c1, 32'h4304dea9},
  {32'h449052a6, 32'h43aca45a, 32'h438a4ddb},
  {32'hc5091c0f, 32'hc299c16e, 32'hc3c2c48d},
  {32'h44c7e3de, 32'h42749462, 32'hc319736e},
  {32'hc5050ec2, 32'hc3a9f0c8, 32'h430b4d86},
  {32'h44ad4af2, 32'h4407cd7f, 32'hc1947857},
  {32'hc4b9be4e, 32'h41fc4652, 32'h438d483a},
  {32'h4509ccfc, 32'h435064d3, 32'h43602e2b},
  {32'hc3b4b2a4, 32'h4384100a, 32'hc21e6f63},
  {32'h450ea091, 32'h434d30a1, 32'h43005e9e},
  {32'hc3c0a374, 32'h42c115f1, 32'h420a2c55},
  {32'h45120ff4, 32'h4319f52d, 32'hc36acf7d},
  {32'hc50f7977, 32'h427d64d4, 32'hc237c7b4},
  {32'h4405cc89, 32'hc28bdcbd, 32'hc1c4da2a},
  {32'hc4d1278a, 32'hc23a5ff7, 32'h4291bb74},
  {32'h44f86279, 32'h43617a13, 32'hc306dbfe},
  {32'hc4c396ff, 32'hc2c21fc9, 32'h4358f615},
  {32'h43ee760c, 32'h43426783, 32'hc41be72b},
  {32'hc50befbe, 32'h43e57c66, 32'h43cc0c26},
  {32'h435c9140, 32'h42da3d69, 32'h43206d36},
  {32'hc4d440ae, 32'hc3ba6342, 32'hc2bb981c},
  {32'h4473d044, 32'h437411b9, 32'h42104c8d},
  {32'hc4a0c342, 32'hc316f8bf, 32'h43699fef},
  {32'h44f09fd5, 32'hc1c7b01a, 32'h43667d56},
  {32'h424d8380, 32'h434f664d, 32'h43d90db2},
  {32'h451b789f, 32'hc2da5d84, 32'hc398ac49},
  {32'h42287600, 32'hc35eec82, 32'h431653c9},
  {32'h440e9174, 32'h42913cce, 32'h4115070a},
  {32'hc4ff1700, 32'h42d1e487, 32'h43ab77a3},
  {32'h44972dd5, 32'h42b3c71d, 32'hc33cf6e9},
  {32'h430807d6, 32'h42e850bf, 32'h426d8dd8},
  {32'h43a99735, 32'h425422e2, 32'hc2925fac},
  {32'hc4317d27, 32'hc342cc69, 32'hc39876d0},
  {32'h44f764f5, 32'h4385a812, 32'h42b62f08},
  {32'hc483b9e4, 32'hc387f5cb, 32'h429d2ff4},
  {32'h4469f9fa, 32'hc2bb0a04, 32'h43e5b04c},
  {32'hc4e3e4c7, 32'hc30731c5, 32'h439b2ef7},
  {32'h44db4219, 32'h41626524, 32'h43de7bdc},
  {32'hc4b3e252, 32'h43b1ab2a, 32'hc2c46b67},
  {32'h44ff2c5d, 32'hc23db3d4, 32'h43f4d587},
  {32'hc502f073, 32'hc3de07c6, 32'hc19f0b35},
  {32'h449bc0a8, 32'hc38410ac, 32'h439f9952},
  {32'hc43a31ca, 32'h430f6a4d, 32'hc348ebd9},
  {32'h44a843d4, 32'h42f04503, 32'h408cd772},
  {32'hc45312a0, 32'hc2d371f9, 32'h4017668e},
  {32'h44a35c40, 32'hc301f014, 32'h4280aa2b},
  {32'hc4c6fe6b, 32'h438045c9, 32'h4208d181},
  {32'h42525c60, 32'hc3f6d564, 32'hc169f93a},
  {32'h409c9280, 32'h438607ab, 32'hc333de77},
  {32'h44831360, 32'h43ae1230, 32'h42861653},
  {32'hc4a51f0d, 32'h4289b462, 32'h420058a9},
  {32'h43d3dc2d, 32'hbfffdffd, 32'h423d5a47},
  {32'hc4d984e5, 32'h42aafaf2, 32'hc21d7156},
  {32'h451daf12, 32'h43b03ee3, 32'hc3cfd78a},
  {32'hc4feaf35, 32'hc34a1f5b, 32'h42ca6118},
  {32'h449e874c, 32'hc327d712, 32'h42efba8a},
  {32'hc45947d4, 32'h42b25e07, 32'hc25cb503},
  {32'h44e480f4, 32'hc2af03cb, 32'h42870ac2},
  {32'hc4a8d40e, 32'hc3732485, 32'h42c07004},
  {32'h44b258b6, 32'h42c21028, 32'hc413e5e1},
  {32'hc4b6c0b1, 32'h43aa49d8, 32'hc324bc44},
  {32'h446fe952, 32'h42bd8678, 32'h429a4c2e},
  {32'hc4cf11d7, 32'h410a58a3, 32'h4226f5a8},
  {32'h44908ce7, 32'hc35285a4, 32'h4316d345},
  {32'hc3fd3c05, 32'h4311a5d5, 32'hc16df21b},
  {32'h425f0de8, 32'hc33402d8, 32'h42e86d43},
  {32'hc4739ed2, 32'h426a5ac4, 32'hc3684e52},
  {32'h4459917d, 32'h4274b4c7, 32'h44148700},
  {32'hc4eecc8f, 32'h43641f83, 32'h42947c45},
  {32'h4503a4ae, 32'h4330d3bb, 32'hc28a5557},
  {32'hc46f546a, 32'hc310edd1, 32'h4308531c},
  {32'h44c29571, 32'h43983b2e, 32'h42de79a6},
  {32'hc4f3fbc6, 32'hc3872429, 32'hc3fdbe68},
  {32'h44da37a8, 32'h4320bc0e, 32'hc21f3a76},
  {32'hc42d95dc, 32'h431bd75b, 32'hc30dc5d0},
  {32'h43c23300, 32'h43321f77, 32'h4312c793},
  {32'hc3d544c4, 32'hc3e4b74e, 32'h4347e3ee},
  {32'h4413bf31, 32'h426b56da, 32'hc3c8aac5},
  {32'hc4cda050, 32'hc30cc37b, 32'h4304034e},
  {32'h4497b917, 32'h438dd15a, 32'h432287aa},
  {32'hc4f37f0c, 32'hc2408e7a, 32'h438604eb},
  {32'h441560ff, 32'hc488ce76, 32'hc3c850bf},
  {32'hc416a2d0, 32'hc31d8a25, 32'hc2715978},
  {32'h43cbe7a0, 32'hc00a8acc, 32'hc288cb4b},
  {32'hc47041fe, 32'h43a14fe4, 32'hc2cf48a0},
  {32'h442a344c, 32'h42c34869, 32'hc289c642},
  {32'hc49fc64d, 32'h432924d3, 32'hc2ffefe7},
  {32'h449f86f4, 32'hc2db8cd5, 32'hc2c769b9},
  {32'hc431ad60, 32'h42c4401a, 32'hc28f1382},
  {32'h44bd6daa, 32'hc2d41b73, 32'hc3f7fae3},
  {32'hc467cba3, 32'hc388ebb9, 32'h43a7b709},
  {32'h4431d3f1, 32'hc33c157b, 32'hc20fc209},
  {32'hc4d8e786, 32'hc2ea5aba, 32'h430098a5},
  {32'h436e84b8, 32'hc2b13ecf, 32'hc21b35b5},
  {32'hc4d15d4e, 32'h42a30bdb, 32'hc2a005b6},
  {32'h44e6e9e8, 32'hc242da31, 32'h4304cdab},
  {32'hc50f14d0, 32'hc2bd6672, 32'hc30573ab},
  {32'h44b8238e, 32'hc305dbf8, 32'h42e9979d},
  {32'hc4ef382e, 32'h4312cb3e, 32'hc2ae5319},
  {32'h44d94ecc, 32'h41fcdbd8, 32'h4212dcfa},
  {32'hc3efa870, 32'hc2f0b43a, 32'h43301aa3},
  {32'h44b98426, 32'h43db1074, 32'hc367b1b4},
  {32'hc48d0472, 32'h437cf1b8, 32'hc3030e1f},
  {32'h443deb05, 32'hc37165d5, 32'hc35962ab},
  {32'hc4e0a5b5, 32'h42b2ece4, 32'h42dbce88},
  {32'h44254596, 32'h43556dd2, 32'hc3555862},
  {32'hc499b6c2, 32'hc1505322, 32'h433a75c9},
  {32'h44908b6a, 32'hc39f7d7c, 32'h42a5fec8},
  {32'hc4a094ae, 32'hc3cebba2, 32'h42d5f76c},
  {32'h4410045c, 32'hc1d43ab4, 32'h439cc708},
  {32'hc48f9e49, 32'h43110343, 32'hc31b498e},
  {32'h44c3a3cf, 32'h41a751a1, 32'hc31a5a11},
  {32'hc49541a4, 32'hc3058fff, 32'hc33a76a9},
  {32'h43b82db4, 32'hc3a846b2, 32'h426ff288},
  {32'hc4fa20e0, 32'hc2a08549, 32'h4244e7b0},
  {32'h44f57c1d, 32'h42a79e97, 32'hc2839bf0},
  {32'hc3a3111a, 32'hc30e83cf, 32'hc38ebb6b},
  {32'h44a8ef2f, 32'h439ff9bb, 32'h435250fb},
  {32'hc47a92bb, 32'hc3145a7f, 32'h4393e2d5},
  {32'h44967d8e, 32'hc36cf192, 32'hc1e0abe2},
  {32'hc4a86cf9, 32'h434ebc23, 32'hc3af726c},
  {32'h447021e0, 32'hc39ac02b, 32'hc372865e},
  {32'hc4e5381a, 32'hc2e792e2, 32'hc2b4bb03},
  {32'h43a17058, 32'h43261497, 32'h439dcbe6},
  {32'hc474604c, 32'hc264f0a7, 32'hc36d68d6},
  {32'h450371aa, 32'h42a258f0, 32'hc1b5683d},
  {32'hc4800932, 32'hc2acef1a, 32'hc2a4ea26},
  {32'h44c2d5ea, 32'hc231921c, 32'h420e1702},
  {32'hc426f6ae, 32'h42703d69, 32'hc36fa586},
  {32'h42d0fc7c, 32'h42b7e6a0, 32'h43e37a68},
  {32'hc4df078c, 32'hc1bed105, 32'h43b720be},
  {32'h4488b2a8, 32'h43ca788f, 32'h41a58b13},
  {32'hc49117de, 32'h42f67a38, 32'hc381594c},
  {32'h43dd914c, 32'h4374b4e8, 32'h43a88ca6},
  {32'hc48ee5e7, 32'h42cc4f6d, 32'hc3e41cf1},
  {32'h4347ca94, 32'hc2bd29bf, 32'hc325afef},
  {32'hc45771a0, 32'hc2116b2f, 32'hc2bf6c0d},
  {32'h449786fa, 32'hc1ce2920, 32'h425f30b3},
  {32'hc44ec2a8, 32'hc2094f90, 32'hc38e277f},
  {32'h4487146e, 32'h42fbe7fe, 32'h424901ff},
  {32'hc397ff04, 32'hc2a804f9, 32'hc22a7465},
  {32'h44c2b8a2, 32'hc337d452, 32'hc39d6501},
  {32'hc27b68e7, 32'h429c3eeb, 32'h4358ab25},
  {32'h44ac524e, 32'hc2d1f49c, 32'hc23f1ec2},
  {32'hc44390dc, 32'h4232952b, 32'hc1e8737b},
  {32'h44eb123d, 32'h420e986b, 32'hc338694e},
  {32'hc48312b6, 32'hc42110a6, 32'h439a5384},
  {32'h4502bd20, 32'h4273c3f6, 32'hc2ec0bce},
  {32'hc4f5153b, 32'hc21a8b98, 32'hc2bbaf6d},
  {32'h44b7d6f0, 32'h4230dce7, 32'hc201e2a1},
  {32'hc32da284, 32'hc32ff481, 32'hc118c375},
  {32'h43bae7b0, 32'hc1f3492b, 32'h425a65a2},
  {32'hc4c14e97, 32'h435ccf95, 32'hc2c9c601},
  {32'h443dadd4, 32'hc28921da, 32'h438caec4},
  {32'hc46fb0a3, 32'h440fcc04, 32'h4382ca16},
  {32'h44852a10, 32'hc3ab2377, 32'h43b5756e},
  {32'hc49959f3, 32'h42c45966, 32'h4305d287},
  {32'h45133417, 32'h41310cbd, 32'h4150aa2f},
  {32'hc4c5191a, 32'hc3777172, 32'h4207c998},
  {32'h4385cb7c, 32'h439f5b6b, 32'hc3661e70},
  {32'hc3926298, 32'h42c1065a, 32'h43200075},
  {32'h4394a148, 32'hc383c80a, 32'h41f0afd2},
  {32'hc4ee1748, 32'hc31bec26, 32'h43f48f13},
  {32'h447393c4, 32'h429c702d, 32'hc30f428a},
  {32'h4373edb6, 32'h43810159, 32'h4301ad67},
  {32'h4350b818, 32'hc2664b04, 32'hc31754ab},
  {32'hc3b11f90, 32'h4325bf90, 32'h438012fb},
  {32'h44ab02fa, 32'hc2a4574a, 32'h43a5138b},
  {32'hc4408b28, 32'h43d3eed8, 32'hc3914586},
  {32'h44d252aa, 32'hc3698bba, 32'h43d8fd9b},
  {32'hc5092a1d, 32'h41655248, 32'h4285df68},
  {32'h451df118, 32'hc2f33fda, 32'h433d0786},
  {32'hc50d8aba, 32'h42f43204, 32'h4382964c},
  {32'h44c54ed7, 32'h432e2660, 32'hc2efa484},
  {32'hc4d2a639, 32'hc2347278, 32'h430ea77b},
  {32'h4508f5e2, 32'hc2f51afa, 32'hc307e76f},
  {32'hc484401e, 32'hc3a78b4b, 32'hc3c60a71},
  {32'h43a92d4c, 32'h405fdbe4, 32'h435ec6f4},
  {32'hc4d9c0de, 32'hc2dc001c, 32'h434e9017},
  {32'h4527e198, 32'hc38b23eb, 32'h439b009b},
  {32'hc3e5f1ca, 32'h43335c80, 32'h41e3577b},
  {32'h438934c8, 32'hc3f0767b, 32'h434f496a},
  {32'hc496518e, 32'hc177bd28, 32'h418ff23c},
  {32'h449f19a0, 32'hc303c888, 32'h4325fd19},
  {32'hc433b404, 32'h43b9af14, 32'hc3566d8a},
  {32'hc382872f, 32'h43c37125, 32'hc33ec534},
  {32'hc50903d4, 32'h436cd5e2, 32'hc3cd68c9},
  {32'h443e3af8, 32'hc2c8faa2, 32'h43f92de7},
  {32'hbfb64b80, 32'h433b33a1, 32'hc1ab7061},
  {32'h44481528, 32'hc2c6e25c, 32'h42c869d7},
  {32'hc47a8072, 32'h437dbdbd, 32'h4308c562},
  {32'h44e62a72, 32'h4390c71f, 32'hc2588809},
  {32'hc4a88ba2, 32'hc2813168, 32'hc422d93b},
  {32'h44ee208f, 32'hc31db92f, 32'h4222605e},
  {32'hc41c9cb3, 32'hc34d427b, 32'hc371e87c},
  {32'h4400f7b3, 32'h4348a844, 32'hc1af682a},
  {32'hc49723e8, 32'hc2a79dbe, 32'hc33eaea1},
  {32'h44fca736, 32'h43525c25, 32'h433e86c6},
  {32'hc4b2621c, 32'h43b9ff12, 32'h438fbb0f},
  {32'h449814da, 32'hc1fe9114, 32'h43a56bbe},
  {32'hc4c61650, 32'hc2f9027f, 32'h432990c9},
  {32'h442d46dc, 32'h439894ec, 32'hc2d07e92},
  {32'hc4348812, 32'hc2976e73, 32'hc4239697},
  {32'h44d1262e, 32'hc3445b95, 32'hc262e9b5},
  {32'h42274098, 32'h43a91797, 32'h4345d33d},
  {32'h44c1e56a, 32'hc3c9fd53, 32'h42d6600e},
  {32'hc4c98486, 32'h428a3206, 32'h41f1034a},
  {32'h44f9d546, 32'hc3111360, 32'h429ade3d},
  {32'hc505849a, 32'hc308ce80, 32'h4264fe36},
  {32'h44b302e9, 32'hc3ecd66a, 32'h4359cbf3},
  {32'hc4dc8069, 32'h424331a3, 32'hc29e7f22},
  {32'h45082b30, 32'h4360fcbc, 32'hc313bb30},
  {32'hc4ecfbfe, 32'h418f3350, 32'h4391ff77},
  {32'h4514a05e, 32'hc31519ce, 32'hc3881326},
  {32'hc4c20cb8, 32'hc0ff24e0, 32'h432a515a},
  {32'h450fff00, 32'hc31a957a, 32'hc3a62694},
  {32'hc4411e2e, 32'h4383b32d, 32'h43c921b6},
  {32'h44204468, 32'hc3bdec0d, 32'hc2d5131f},
  {32'hc49b9f04, 32'hc310811d, 32'hc31bc8e3},
  {32'h45006edf, 32'h43c4ce0b, 32'h42633b72},
  {32'hc3d55ce0, 32'hc3187a8a, 32'h438ac9c0},
  {32'h451a016c, 32'hc309ff83, 32'h42d47c43},
  {32'hc48395ca, 32'h43861262, 32'hc1d6833b},
  {32'hc2e5b18e, 32'h42b91339, 32'hc1fe95dc},
  {32'hc3f8dec0, 32'h43665bce, 32'hc2153dcc},
  {32'h44893c4c, 32'hc38f7ca2, 32'h4380e9ee},
  {32'hc4658610, 32'hc3a9c23c, 32'hc2090487},
  {32'h446c0bf7, 32'hc31eb5c7, 32'hc3eb96eb},
  {32'hc50297b6, 32'h43204e26, 32'h42ee9948},
  {32'h44ba4c7c, 32'h42dad8fc, 32'hc31460f3},
  {32'hc498f3b1, 32'h4390109e, 32'h41b869a2},
  {32'h44657afc, 32'h436574d3, 32'h4383f6c2},
  {32'hc4d6952f, 32'hc301ff5e, 32'h4306265d},
  {32'h438b6570, 32'h431fca49, 32'h43c49e71},
  {32'hc520834e, 32'h4325b54e, 32'hc2df42c4},
  {32'h451511eb, 32'h437b6347, 32'h42d8eeee},
  {32'hc4cc6d6e, 32'h433d61c3, 32'hc2d5424a},
  {32'h438bc220, 32'h43b608b4, 32'hc39747d4},
  {32'hc4ada514, 32'hc2301b90, 32'h4394a506},
  {32'h440bf8d7, 32'h4324e6df, 32'h438dee4e},
  {32'hc4b49f33, 32'hc3566aa7, 32'h41664362},
  {32'h450a765f, 32'h436eb0ec, 32'h42bea1bb},
  {32'hc39807e8, 32'hc3525775, 32'hc033ea84},
  {32'h44b709f0, 32'h40cc5e24, 32'hc1bf87d8},
  {32'hc444ba42, 32'hc3fbf625, 32'hc2c3b281},
  {32'h44d09c5b, 32'hc3100f58, 32'h43089ea0},
  {32'hc4bda89d, 32'h43908dd8, 32'h437f9f7d},
  {32'h444dff64, 32'hc331c474, 32'hc32b8c78},
  {32'hc2837078, 32'hc314aaef, 32'h428da354},
  {32'h431cbc3c, 32'hc384e3b0, 32'h42979637},
  {32'hc52a428a, 32'hc1c53704, 32'hc34684ef},
  {32'h45008748, 32'hc37deaef, 32'hc3a9593b},
  {32'hc34ae120, 32'hc31e380d, 32'hc2fb9193},
  {32'h44a98a4e, 32'hc24223a8, 32'h42ed9b94},
  {32'hc4bf327d, 32'hc2c5937c, 32'h4341f417},
  {32'h43fe3133, 32'h43860702, 32'hc294d3ce},
  {32'hc3c355d8, 32'hc3c45c43, 32'h43a0666c},
  {32'h4474a196, 32'h439891cd, 32'hc3281d47},
  {32'hc4bcb9f7, 32'h43d1f180, 32'hc30d0fd6},
  {32'h44abed08, 32'hc31fe524, 32'h41de442c},
  {32'hc4bb26f5, 32'h4303fff4, 32'h439dcf28},
  {32'h44ace826, 32'hc33e31f8, 32'h432ce64c},
  {32'hc49cb439, 32'hc23b0cbf, 32'hc3b59b29},
  {32'h450a73cb, 32'hc1e9121e, 32'h429fd105},
  {32'hc49b6515, 32'h43917fe4, 32'h43eb6e69},
  {32'h4496a449, 32'h421d8820, 32'h42333637},
  {32'hc380d790, 32'h4314eccf, 32'h431d4bb4},
  {32'h44c09e8d, 32'h42504833, 32'hc2af6c14},
  {32'hc4a81865, 32'h43361989, 32'h43869648},
  {32'h446235a4, 32'h43a887ba, 32'hc402de80},
  {32'hc3b12785, 32'hc365f56b, 32'hbfbc2ef4},
  {32'h450bc804, 32'hc3459049, 32'hc3bdd01b},
  {32'hc4437e44, 32'h4330112a, 32'hc2e3b714},
  {32'h4490da1e, 32'h4315234c, 32'hc39ba58d},
  {32'hc49f6a00, 32'h43ba1cf8, 32'h43027f94},
  {32'h450c69ee, 32'h428ff4d1, 32'h40d9df8a},
  {32'hc4c38c47, 32'hc20713a6, 32'hc1d0f7b3},
  {32'h44541e6a, 32'h42e7d6bd, 32'hc10de5b8},
  {32'hc4d475e6, 32'h43fec8e3, 32'h4169a8cc},
  {32'h450aa2f9, 32'h4405f8b7, 32'h3efa271a},
  {32'hc4f6dbda, 32'hc2adabce, 32'hc2861338},
  {32'h4405ec54, 32'h4382421a, 32'hc0aac1a6},
  {32'hc395614c, 32'hc3630eda, 32'hc1d0e522},
  {32'h446af56a, 32'hc34f0999, 32'hc2bcd364},
  {32'hc3bddb34, 32'h42b4207c, 32'h4267e34c},
  {32'h42718390, 32'hc30c5f31, 32'hc16acdc4},
  {32'hc4f50093, 32'h41fc76dd, 32'h43fa0b3c},
  {32'h43a0fbdf, 32'hc32d763f, 32'hc328072a},
  {32'hc430b6dc, 32'h43836fa6, 32'hc1db1365},
  {32'h44a00616, 32'hc198ffce, 32'h433a9c23},
  {32'hc445995c, 32'h438f5844, 32'hc232dd41},
  {32'h44b7842c, 32'h42a3a652, 32'hc2165748},
  {32'hc4d4906d, 32'hc37805f1, 32'h43ca13fd},
  {32'h44cb29b4, 32'hc32f4ab1, 32'hc39bcfe5},
  {32'hc4df75f4, 32'hc176004c, 32'h435f756e},
  {32'h44032bf0, 32'hc1be5230, 32'h423f822f},
  {32'hc45f4d46, 32'h428c969a, 32'h435108b3},
  {32'h44eb7ae9, 32'hc1e32774, 32'hc323604f},
  {32'hc3bd3ee2, 32'h434cbcd1, 32'h4399efdc},
  {32'h44c73683, 32'hc32cd1c2, 32'hc3dc317e},
  {32'hc4390458, 32'hc1835267, 32'h427d42f1},
  {32'h43f13408, 32'hc3883141, 32'hc34a0ef3},
  {32'h445ace20, 32'hc3d99b68, 32'hc35fdd24},
  {32'hc4b1cc5c, 32'h430fbb77, 32'hc32d2e5b},
  {32'h44fa6b88, 32'h4343697e, 32'h430dcaad},
  {32'hc4f789f8, 32'h40bf940d, 32'h42ae5bde},
  {32'h44b92134, 32'hc4051fbb, 32'hc3bf740c},
  {32'hc4871682, 32'h43620119, 32'h42c9f2e7},
  {32'h41ef8cc0, 32'h41affd24, 32'hc3f2042c},
  {32'hc4d46949, 32'h4314987b, 32'hc13006f9},
  {32'h440a49e2, 32'h4357ddef, 32'hc219dd0a},
  {32'hc4ced447, 32'hc38607db, 32'h40c61a51},
  {32'h4396ad30, 32'hc2af1133, 32'hc3218342},
  {32'hc51183b3, 32'hc3068fe6, 32'hc30f6c3d},
  {32'h450cf51d, 32'h435dc1ff, 32'h42ed5499},
  {32'hc3a80566, 32'h42a73330, 32'hc1f79fc3},
  {32'h44962412, 32'h43bf8fca, 32'h4356572a},
  {32'hc4e781a8, 32'hc24157c8, 32'h43824864},
  {32'h450940c0, 32'hc34d12cb, 32'h42eb202d},
  {32'hc4bb6570, 32'hc395d481, 32'h43314f21},
  {32'h440c150d, 32'hc3873ea6, 32'hc2fe46a9},
  {32'hc4042b60, 32'hc2045fa2, 32'h43541feb},
  {32'h449d3753, 32'h435d8023, 32'h43da81ac},
  {32'hc503facd, 32'hc38d1d92, 32'h421256de},
  {32'h42e65860, 32'h4380bb2d, 32'hc41d14fc},
  {32'hc484d4be, 32'hc302a790, 32'h438e77b8},
  {32'h44a5c245, 32'h42a40491, 32'hbf266840},
  {32'hc3e9d8b4, 32'h431b419b, 32'h3f77b380},
  {32'h451b9883, 32'hc3af45fc, 32'h4402178d},
  {32'hc51525f4, 32'hc2e5a300, 32'h43b65257},
  {32'h44191ede, 32'h43dfa9e3, 32'hc2922e98},
  {32'hc510bb19, 32'h4296c2be, 32'hc2fbfd2e},
  {32'h44236128, 32'hc3b33a81, 32'h42d9c9dc},
  {32'hc4b4673b, 32'hc398c825, 32'hc34d2ebf},
  {32'h44bd6716, 32'hc30b89bb, 32'hc2264b5b},
  {32'hc4d52df6, 32'hc1a094f2, 32'h42e02103},
  {32'h45055e88, 32'h43518a8d, 32'hc3057fab},
  {32'hc4ed8b6a, 32'h4245844e, 32'h41c00040},
  {32'h4433e670, 32'h433918fc, 32'hc2a9300f},
  {32'hc48aaf03, 32'h43c5c7c7, 32'h41b05f86},
  {32'h4405c59b, 32'h431caa16, 32'h430e5ffe},
  {32'hc465da8a, 32'hc2e81ee7, 32'h43601a1d},
  {32'h44b72eb2, 32'hc0033fca, 32'hc345ccb5},
  {32'hc41d557e, 32'h437ae2df, 32'h43cc044e},
  {32'h45109a50, 32'hc23cc672, 32'h43b01a94},
  {32'hc50a8d2c, 32'hc220ce2e, 32'hc29ee6c6},
  {32'h442a929e, 32'hc2f3225b, 32'h430e7866},
  {32'hc3ec7ad0, 32'hc26e78d0, 32'h42bbe94e},
  {32'h448d2c15, 32'hc2e03dc0, 32'h434c1136},
  {32'hc49598c6, 32'h4322d57a, 32'hc3bdc53d},
  {32'h4403d60c, 32'hc27a21e4, 32'h43b89857},
  {32'hc50043b3, 32'hc3cdf5e4, 32'h43f4cfeb},
  {32'h43678ba0, 32'hc3433713, 32'hc2ff8f0a},
  {32'hc499c29e, 32'h43c3ef12, 32'hc3ae49ed},
  {32'h44a6b71c, 32'hc2ab4823, 32'hc3584032},
  {32'hc48bb410, 32'hc3af5012, 32'hc3e4a98e},
  {32'h4353c1f4, 32'hc2299ee9, 32'hc33459f4},
  {32'hc4a1fa8e, 32'h42d0e10c, 32'hc39841f1},
  {32'h4503fe92, 32'hc29290f4, 32'hc29c7e8d},
  {32'hc4ae79bf, 32'hc33a494e, 32'h4270ef5d},
  {32'h44c01294, 32'h431522e0, 32'h43c23cd5},
  {32'hc4d4d18d, 32'h43bda7b2, 32'hc3bb8d30},
  {32'h451cd687, 32'hc255d7cf, 32'hc3b42ba6},
  {32'hc3e18bfb, 32'h405b2c01, 32'hc3749ac9},
  {32'h44a03143, 32'hc3dc4cdb, 32'hc30ea2d4},
  {32'hc47f53a4, 32'hbfed59a4, 32'hc23ae020},
  {32'h44b21143, 32'h4319b212, 32'h41dc06a8},
  {32'hc510ce29, 32'h4372523e, 32'h43438d49},
  {32'h44bccde2, 32'hc36bb4ce, 32'h425638f2},
  {32'hc5081e99, 32'hc2e4e32e, 32'hc0eba931},
  {32'h4506535d, 32'hc359b426, 32'hc32ab49b},
  {32'hc2fe7390, 32'h42d3f09a, 32'h4293c6d1},
  {32'h44779e72, 32'h42c1215e, 32'h438192ba},
  {32'hc4244bea, 32'hc371a4a0, 32'h431af847},
  {32'h44909dc9, 32'h43938c39, 32'h4325a6d8},
  {32'hc5003549, 32'hc1a442d4, 32'h42c62be7},
  {32'h4468009d, 32'h4365256c, 32'h43dde08c},
  {32'hc3b0179f, 32'h43aed937, 32'hc30c0329},
  {32'h43ecded0, 32'h42da2a15, 32'hc07aa3a5},
  {32'hc4e3b8ca, 32'h43a057aa, 32'h4385e82e},
  {32'h43abab20, 32'hc38406b6, 32'h4224c0ce},
  {32'hc4a25da9, 32'h43485bd0, 32'h42b62262},
  {32'h44c7b47f, 32'hc26e4b8b, 32'h437953c8},
  {32'hc4aa5550, 32'hc0beb4da, 32'hc2c2317b},
  {32'h440aeea9, 32'h42ff83e2, 32'hc261c1fb},
  {32'hc3d2498c, 32'hc2c794cd, 32'h42bb8f0b},
  {32'h44dc3c8d, 32'hc3106138, 32'hc3377fc2},
  {32'hc4d3f35e, 32'hc2d18c9a, 32'h43996078},
  {32'h4416ebf2, 32'hc1b83d0b, 32'hc3322527},
  {32'hc48add36, 32'hc12fc8b7, 32'h430cd551},
  {32'h441faad1, 32'hc3488703, 32'h43f46d62},
  {32'hc4885c72, 32'hc389d627, 32'hc321020f},
  {32'h44ebdf0d, 32'hc3451aad, 32'hc3252b55},
  {32'hc3ab4620, 32'hc313af43, 32'h4107001c},
  {32'h4503e225, 32'hc325e49a, 32'hc3bbc4a4},
  {32'hc4bbb354, 32'h437d6cad, 32'hc30ff8fb},
  {32'h44c45004, 32'hc287c2ed, 32'h43971b46},
  {32'hc4ce55c9, 32'hc2af1602, 32'h43a8b53b},
  {32'h44d49dbb, 32'hc2875d21, 32'h42cd0b85},
  {32'hc35e6d00, 32'hc2b4ba79, 32'h42b7c1ca},
  {32'h4388113c, 32'hc23e4497, 32'h4376afc2},
  {32'hc4b11706, 32'hc13d3e48, 32'hc17e623f},
  {32'h4477af8c, 32'h43832593, 32'h423e34b7},
  {32'hc4238d00, 32'h4236f906, 32'h43feb2c3},
  {32'h4502da5c, 32'h4312901f, 32'h435c995a},
  {32'hc3dc15c6, 32'hc2b76ffc, 32'h4397238d},
  {32'h4484a898, 32'hc1144003, 32'h4334ba37},
  {32'hc4ea2d07, 32'h438a1281, 32'h42e54aae},
  {32'h4421a2da, 32'hc1992b51, 32'hc2811b44},
  {32'hc3963a08, 32'hc3d537c8, 32'hc2b53468},
  {32'h4461d08c, 32'hc28d6037, 32'h4314e4e3},
  {32'hc4c895d1, 32'hc37296b5, 32'h4331e1af},
  {32'h443fa801, 32'hc403d624, 32'hc32c34cd},
  {32'hc4dfd05e, 32'h42f6c957, 32'h42bf800a},
  {32'h44ded553, 32'h41f3d93d, 32'hc366a9d4},
  {32'hc49defbd, 32'h42b4df26, 32'h434f3089},
  {32'h44cab334, 32'h424310ea, 32'hc06a9f7a},
  {32'hc489170e, 32'h4224480e, 32'hc34523aa},
  {32'h44862592, 32'hc3202034, 32'h43371867},
  {32'hc32b4e5c, 32'h434c04c3, 32'hc2b53e93},
  {32'h44b5dd7d, 32'hc2bd88d6, 32'h4239ff98},
  {32'hc5018973, 32'h433b86e4, 32'hc3960131},
  {32'h44069987, 32'hc42c86ad, 32'h41f4a044},
  {32'hc511fbab, 32'hc3655986, 32'hc313f327},
  {32'h4473403e, 32'h4301ad9a, 32'h4225c792},
  {32'hc4d08081, 32'hc3a5cfe8, 32'h42d94a8d},
  {32'h4408cdf3, 32'h432107f6, 32'hc3697eae},
  {32'h42fd87a0, 32'h41f7e066, 32'hc229f774},
  {32'h43bc692a, 32'hc305a0f9, 32'h42d95d34},
  {32'hc3e01d20, 32'h43b6e9f8, 32'hc2decd9d},
  {32'h451ac7c4, 32'h43976a0b, 32'h42bbcd7a},
  {32'hc4843985, 32'h4389caa3, 32'h436ec7f6},
  {32'h4514ab6a, 32'hc419e960, 32'h43fbf538},
  {32'hc5085ddb, 32'h4474c947, 32'hc0b7176a},
  {32'h44986cd0, 32'hc363e521, 32'h421b2cd9},
  {32'hc4567a98, 32'hc2fa3e43, 32'hc32d667b},
  {32'h43724e90, 32'h435e48f5, 32'h42e2d3e9},
  {32'hc4bc92cf, 32'hc30a5746, 32'h43178efe},
  {32'h44654fb2, 32'h43da1a91, 32'hc1103b58},
  {32'hc5038433, 32'h4349d125, 32'h436bfc3b},
  {32'h44d947a5, 32'hc3cb50f7, 32'h4330ad35},
  {32'hc2babb20, 32'h418119b8, 32'hc21ac356},
  {32'h438578e6, 32'h42e129d6, 32'hc295e89e},
  {32'hc5023650, 32'h42a647b2, 32'h43d9b4c6},
  {32'h43cb0ef7, 32'h43b132fc, 32'h43b0eea4},
  {32'hc36ae870, 32'hc3c90cc2, 32'hc32d0a27},
  {32'h42fba6c0, 32'h43cddec7, 32'hc3211b64},
  {32'hc4b9eef9, 32'h42703be2, 32'hc35c183f},
  {32'h44eb4edd, 32'h42d2b507, 32'hc3b33db5},
  {32'hc439ca87, 32'h427d452c, 32'h43c5f0b3},
  {32'h44c55350, 32'h423d18f0, 32'hc30ea863},
  {32'hc48245ca, 32'h42bf4581, 32'h4362713e},
  {32'h44af123e, 32'hbfc36478, 32'h435d61ce},
  {32'hc492eef0, 32'h42e05586, 32'h411d2c8c},
  {32'h445edb20, 32'h43355b7d, 32'hc201e3aa},
  {32'hc2a3ab49, 32'hc2daaba5, 32'h4208d174},
  {32'h44fbb537, 32'h4280636d, 32'h429f80fa},
  {32'hc4255d86, 32'hc2825711, 32'h42e2778b},
  {32'h43ee8f58, 32'hc305c6de, 32'h42e94c43},
  {32'hc43d3c2d, 32'hc3238f2e, 32'hc3b19679},
  {32'h43aca4cf, 32'hc1d514c3, 32'hc31ed298},
  {32'hc5077737, 32'h44110c99, 32'h4309c9a7},
  {32'h44faccce, 32'h4314764a, 32'hc254d887},
  {32'hc4270ad2, 32'hc1a1ceb2, 32'h42c1967d},
  {32'h447feff8, 32'hc1e61647, 32'h42f0ac46},
  {32'hc4bc2558, 32'hc3c28a5c, 32'hc2eecccc},
  {32'h445a0726, 32'h41985425, 32'hc329a0d5},
  {32'hc3a337b8, 32'h42af4ef2, 32'h4390766f},
  {32'h443a39c4, 32'h43e49438, 32'hc32c3b4f},
  {32'hc4b609a7, 32'hc337abf2, 32'hc333f1f4},
  {32'h43746a0c, 32'hc3b2e2d8, 32'h43de78d4},
  {32'hc4c66a22, 32'hc41fd624, 32'h43fcddc3},
  {32'h444c7664, 32'h432ec1ac, 32'h4376588d},
  {32'hc3ff58b8, 32'hc375731b, 32'h42e529c4},
  {32'h44c15f07, 32'h4337eaec, 32'hc23e1e71},
  {32'hc3395c35, 32'h43074fc5, 32'hc2e21561},
  {32'h44db368c, 32'hc26d5c73, 32'hc2d39726},
  {32'hc4ff8f48, 32'hc25c7d3f, 32'hc100f855},
  {32'h448757df, 32'h4339408f, 32'hc1ddb6de},
  {32'hc3c5d2c4, 32'h432b722e, 32'h4138dcea},
  {32'h44f1ee0d, 32'h42adbd91, 32'hc3a34a33},
  {32'hc3aaf389, 32'hc35e02c9, 32'hc30fbd81},
  {32'h450a8e68, 32'h418ebe66, 32'hc407dedf},
  {32'h42408e80, 32'h43061b65, 32'hc2687f3b},
  {32'h445c1800, 32'hc370afcd, 32'h423de2e2},
  {32'hc455eed0, 32'h4380a388, 32'h4377777c},
  {32'h448e8903, 32'hc22c81a8, 32'hc1a8e15d},
  {32'hc48be2b2, 32'h41d69ed7, 32'h43217982},
  {32'h44847645, 32'h43fbaf5d, 32'hc316b456},
  {32'hc49d7fa9, 32'h42e30ce6, 32'h43df8ff0},
  {32'h442f7a02, 32'hc348d273, 32'h439ada08},
  {32'hc47c302e, 32'hc381169f, 32'hc3c5078d},
  {32'h450225d5, 32'h4351d84a, 32'h4205403a},
  {32'hc4fdd887, 32'h3fce0454, 32'h42aea250},
  {32'h4519a5f5, 32'h4367b970, 32'h43047941},
  {32'hc4cbfae5, 32'hc1dc740a, 32'h41171882},
  {32'h44a8ba62, 32'hc3116a95, 32'h4315b0b1},
  {32'h409c72b8, 32'hc38cd1b0, 32'h43263639},
  {32'h44b7f7be, 32'h4371feb8, 32'hc39df3c1},
  {32'hc502cc9d, 32'h42b6236e, 32'h42b15bd1},
  {32'h4489d7d4, 32'hc35b4e02, 32'h43a55154},
  {32'hc4b0695e, 32'hc3017712, 32'h432c4123},
  {32'h449772f2, 32'h42948f35, 32'hc2b31c64},
  {32'hc49b8edc, 32'hc2803cad, 32'h4209dba7},
  {32'h4420a6cc, 32'h432480f3, 32'hc18a43db},
  {32'h432c93a4, 32'hc28cffb7, 32'hc347c868},
  {32'h44ef2e1c, 32'hc266c1c4, 32'h440805af},
  {32'hc4d7550a, 32'hc326aef9, 32'hc3a0b61f},
  {32'h44add72a, 32'h4255d739, 32'hc3d98b4e},
  {32'hc5033753, 32'hc30679c7, 32'hc397d4bd},
  {32'h4492121b, 32'hc20194b5, 32'h43b48d91},
  {32'hc46242db, 32'hc35db662, 32'h43e3ee53},
  {32'h450fb658, 32'hc0c2f963, 32'hc43d2714},
  {32'hc4e9fe94, 32'hc338232e, 32'hc295fbf4},
  {32'h4388a75a, 32'h41b236e1, 32'h42e35cc9},
  {32'hc4b8a9f6, 32'h4380de41, 32'h4309c363},
  {32'h44127fd0, 32'h423da1d5, 32'h42eedca2},
  {32'hc3fd0e20, 32'hc25ebf2c, 32'h431aad41},
  {32'h44d98549, 32'h424b35f0, 32'hc3bab2d0},
  {32'hc51821fa, 32'h42e617db, 32'h43a440f4},
  {32'h44305638, 32'hc3d6db9e, 32'h431607fe},
  {32'hc400e1a2, 32'hc33fbe0c, 32'hc390cfd1},
  {32'h435d7c50, 32'h434ce0f7, 32'h4281c502},
  {32'hc44ebcf2, 32'h42ca5a40, 32'h429efff7},
  {32'h4481f828, 32'hc2201efc, 32'hc2266674},
  {32'hc4db742b, 32'hc2af1ab8, 32'hc38bc99a},
  {32'h44f39440, 32'hc2b4fdc8, 32'h41be218a},
  {32'hc485de8e, 32'hc3a90bb4, 32'hc2d7ee0d},
  {32'h44b44718, 32'hc303c572, 32'h439ffa62},
  {32'hc4c62386, 32'h43932f6a, 32'hc318bd80},
  {32'h450afb9a, 32'h43885937, 32'hc2bd252c},
  {32'hc409cce6, 32'h4381ef53, 32'hbf936ec1},
  {32'h45159cc9, 32'hc0c958da, 32'hc36b741f},
  {32'hc44b2ca0, 32'hc2f8c7a6, 32'hc2109f2e},
  {32'h43ab8f88, 32'hc28c7f59, 32'hc381c231},
  {32'hc41c551c, 32'h42f9dc0b, 32'h43001c8c},
  {32'h4406fb48, 32'hc2283f40, 32'hc3c1fe41},
  {32'hc4d1aec1, 32'hc1971c7b, 32'hc40ab0b4},
  {32'h424422c4, 32'h43485674, 32'h4360734b},
  {32'hc4d5cf65, 32'hc3755735, 32'h42b0e318},
  {32'h448365c0, 32'h43938c81, 32'hc3e950ba},
  {32'hc498080f, 32'h4305a1a6, 32'h43ce6676},
  {32'h4508f5a0, 32'hc2f23ae7, 32'h43802b81},
  {32'hc4b803e0, 32'h42e7e1c0, 32'hc395c4ff},
  {32'h4420fa60, 32'h429a9df9, 32'hc2b7d919},
  {32'hc513fa70, 32'hc2913618, 32'h427cd3d3},
  {32'h44ff4a86, 32'hc2ba7c00, 32'h41d6db8f},
  {32'hc4b204a5, 32'hc1a7e973, 32'hc38808f7},
  {32'h442f6c87, 32'h422780a7, 32'hc38e7a4a},
  {32'hc2e7bc78, 32'hc2a3ce4a, 32'h43a005ff},
  {32'h447be719, 32'h43d7312e, 32'hc22446e7},
  {32'hc4c0f3ee, 32'h4357b361, 32'h435f2e80},
  {32'h44dc9fdb, 32'h4338af4c, 32'h43bada37},
  {32'hc4c0bc7b, 32'hc3802796, 32'h432b889f},
  {32'h448a67d3, 32'h43fb7958, 32'hc3e76b24},
  {32'hc4a87e8a, 32'hc1f80ca7, 32'hc29673bd},
  {32'h43ded300, 32'hc372ce65, 32'h42ecca20},
  {32'hc3c183aa, 32'hc3b1adcc, 32'hc38e6b77},
  {32'h44ecce86, 32'hc3700742, 32'hc2887a67},
  {32'hc505d529, 32'h4311596e, 32'h42c78e1d},
  {32'h449bf12f, 32'hc2ece9e4, 32'hc4029f02},
  {32'hc411e959, 32'h4314a259, 32'h436a5db6},
  {32'h44035dc9, 32'hc3df8127, 32'h42f50b74},
  {32'hc3f6a0dc, 32'hc37c8d4d, 32'h4109c2b6},
  {32'h450f7916, 32'h44095a19, 32'h43be07ef},
  {32'h422e8fe0, 32'h43039b60, 32'h3efe9450},
  {32'h440594fc, 32'hc4468434, 32'h43150624},
  {32'hc37c0f45, 32'hc30946e4, 32'hc383c37d},
  {32'h45168e95, 32'h439a9890, 32'hc3918e83},
  {32'hc4c7339f, 32'h43160732, 32'h4285ff97},
  {32'h445737d7, 32'h429d0ddf, 32'hc34428b6},
  {32'hc4ea446b, 32'hc08eeeac, 32'hc3c20243},
  {32'h451c8c99, 32'hc38bb87d, 32'h42e40d5c},
  {32'hc503069a, 32'hc29f6e8c, 32'h437e3dc2},
  {32'h44da1775, 32'h41899579, 32'hc2ae2b73},
  {32'hc3df5c24, 32'h431de68a, 32'hc35c1680},
  {32'h45227bdb, 32'hc322b362, 32'hc2e366b5},
  {32'hc4f794b6, 32'h4367071f, 32'hc3187ea6},
  {32'h450b8bd7, 32'h437518c3, 32'hc35eb702},
  {32'hc4cc5983, 32'h4195dbbe, 32'hc30c6cac},
  {32'h431d2428, 32'hc30c9315, 32'h42a4b48a},
  {32'hc4974902, 32'h43037cf5, 32'hc3aeb02e},
  {32'h43bfec84, 32'h41bd3a65, 32'h434faa4d},
  {32'hc509a96b, 32'hc0588ee0, 32'h419db7e0},
  {32'h44b6533e, 32'h437e1b63, 32'h43a75e53},
  {32'hc447e747, 32'hc2befe77, 32'h420ac983},
  {32'h44e60156, 32'h4219a7b5, 32'hc34209e1},
  {32'hc4a856a4, 32'hc21378d3, 32'hc28d384e},
  {32'h451d43c5, 32'hc1e05566, 32'hc28449ca},
  {32'hc510e9d7, 32'h4313e6d7, 32'hc2820c3a},
  {32'h44efeccd, 32'h43c8f982, 32'h43bf2681},
  {32'hc1ce5140, 32'h430ecead, 32'hc3aad70d},
  {32'h44a1ef92, 32'h435b0d10, 32'hc3b50b6a},
  {32'hc50f6274, 32'h432e56f0, 32'h436855a8},
  {32'h44b0d4b8, 32'hc1d0d4f4, 32'h42b56b97},
  {32'hc5126dda, 32'h438fbb72, 32'h436a4281},
  {32'h4353544a, 32'h43152ed5, 32'hc3bdb3d1},
  {32'hc50bddd6, 32'h43b8a280, 32'hc2f74200},
  {32'h44e3fc2b, 32'h4135cc8b, 32'hc2f758ea},
  {32'hc42a6c5b, 32'hc1983d2e, 32'hc2662498},
  {32'hc3ca6bb5, 32'hc30d78b1, 32'h4354394c},
  {32'hc216f380, 32'hc31d1433, 32'hc382f09b},
  {32'h44ebe8ae, 32'hc224da5e, 32'hc3390ba0},
  {32'hc4b848ac, 32'h43bdce6c, 32'hc30d6321},
  {32'h4520e80a, 32'h43650e54, 32'hc31c414d},
  {32'hc4b809da, 32'hc27b71d0, 32'hc3c3acf3},
  {32'h4426431a, 32'h43800663, 32'hc3a27412},
  {32'hc482396e, 32'hc1d28c85, 32'h43a67960},
  {32'h440ade58, 32'h43e1be37, 32'hc2d2147e},
  {32'h42f433e0, 32'h440e1cc7, 32'hc312cb37},
  {32'h4475857e, 32'hc39b5fea, 32'h43a3eea5},
  {32'hc4de2849, 32'hc2d26822, 32'h43ea8163},
  {32'h4518b3bc, 32'hc2c2977a, 32'hc2f62f28},
  {32'hc4b40db4, 32'hc22804bb, 32'h421b4d70},
  {32'h4487b723, 32'h4169e852, 32'h436c9d4e},
  {32'hc51802ec, 32'hc3165730, 32'h42be7635},
  {32'h4512418f, 32'hc343fd34, 32'h42d3f367},
  {32'hc4f36021, 32'hc2705bd9, 32'h4335e62c},
  {32'h441b3124, 32'h43280999, 32'hc28c1678},
  {32'hc4cf2f20, 32'hc2cc151c, 32'h43e1822e},
  {32'h44c9c2d0, 32'hc2ee700e, 32'hc3808479},
  {32'hc4f0905c, 32'h4383ffb7, 32'hc3b1f53b},
  {32'h44d6564d, 32'h4313422f, 32'h4394f402},
  {32'hc47a2592, 32'hc2e508c6, 32'h43b3ce30},
  {32'h44bf44a6, 32'h41dd2996, 32'h43600c19},
  {32'hc4c36e59, 32'h41c8ba32, 32'hc376f50f},
  {32'h44d517ff, 32'h42f81f25, 32'hc1cec9c9},
  {32'hc4ac45c6, 32'h42a5ca1e, 32'hc3b7d57b},
  {32'h45013e3f, 32'hc334cf2d, 32'h43275397},
  {32'hc4788757, 32'h41f51de0, 32'hc304e97b},
  {32'h44cef54b, 32'h43345874, 32'h43987774},
  {32'hc5118f22, 32'hc3361981, 32'hc3c3a953},
  {32'h44f108f6, 32'h43274cd3, 32'h432c19c5},
  {32'hc49b4724, 32'hc2dfd048, 32'h43a6f860},
  {32'h4510f736, 32'h42e47e73, 32'hc370f9dd},
  {32'hc39fe4de, 32'hc37e8bee, 32'hc3e5d6bf},
  {32'h44d17ada, 32'h42d02966, 32'hc38b8045},
  {32'hc40772e4, 32'hc11e573e, 32'hc302854a},
  {32'h450d1edb, 32'hc1c39311, 32'hc2866c25},
  {32'hc4a91827, 32'h430fad12, 32'hc34c9675},
  {32'h4452ce01, 32'hc2c5c90f, 32'h428a0862},
  {32'hc4cd7bbf, 32'hc4082050, 32'hc3134d36},
  {32'h44dc09df, 32'h43c70a5a, 32'hc1d50d6b},
  {32'hc4a0d8ea, 32'hc3bad4df, 32'hc3390681},
  {32'h448b413c, 32'h43bd90c0, 32'h4314b5d7},
  {32'hc4f61371, 32'h425c9bb9, 32'hc304fcd5},
  {32'h4488eb99, 32'h42531de0, 32'hc3c496bb},
  {32'hc4014d7c, 32'hc2809b5c, 32'h41b35420},
  {32'h449d18a2, 32'hc431a216, 32'hc3586680},
  {32'hc493fde2, 32'h438aa79a, 32'h4314840a},
  {32'h4462d688, 32'hc29c5122, 32'hc390c58f},
  {32'hc4c7974c, 32'h438ae6bf, 32'hc2cf2040},
  {32'h43982f68, 32'h4354766e, 32'h435d2e1c},
  {32'hc4c8a78e, 32'h429a613b, 32'h422d658e},
  {32'h4497fe3b, 32'h4312236f, 32'hc336908a},
  {32'hc4fe8e55, 32'hc2f86cc1, 32'h40d6f62a},
  {32'h4510b56b, 32'h431d8189, 32'h430328df},
  {32'hc4512d5e, 32'h437873b8, 32'hc2883cb4},
  {32'h43c9b87b, 32'hc3840908, 32'h438d70b4},
  {32'hc41f4037, 32'hc42872ad, 32'h3fd031ad},
  {32'h44cb24ec, 32'h42c1dc8c, 32'hc27fc3e6},
  {32'hc494c303, 32'h433a5179, 32'h4320fe45},
  {32'h434b8e60, 32'h430ca14d, 32'h42954b81},
  {32'hc500cff7, 32'h3f11adbc, 32'h41c2bbe3},
  {32'h44d116bf, 32'hc2dac010, 32'hc290a9e6},
  {32'hc499f655, 32'hc2a36700, 32'h439afec4},
  {32'h44df505a, 32'hc34303fe, 32'h42a3ddf8},
  {32'hc5022a3e, 32'hc384591c, 32'hc3068e38},
  {32'h4446e650, 32'hc0dc5c1a, 32'hc3300949},
  {32'hc2d88b78, 32'h437a7ff9, 32'h431c9058},
  {32'hc2797fe0, 32'h435b9cfc, 32'hc3a2068f},
  {32'hc50fc012, 32'h43d3f1e6, 32'h433f58b9},
  {32'h44302c30, 32'h43308668, 32'h420bec0d},
  {32'hc3c5460c, 32'hc3d918b5, 32'h42d45050},
  {32'h449054b8, 32'hc390cfe6, 32'hc4119549},
  {32'hc4910ab6, 32'h42123d90, 32'hc2afd9a0},
  {32'h44899873, 32'h433780fe, 32'hc0e345d4},
  {32'hc4ef039f, 32'hc30327c4, 32'hc26741bd},
  {32'h3fabf100, 32'hc2dd27bb, 32'hc35fbc26},
  {32'hc48b445f, 32'hc3938f10, 32'hc3b4d420},
  {32'h4422d000, 32'h41972906, 32'h429429c6},
  {32'hc510ee8a, 32'hc3234eb6, 32'hc387073b},
  {32'h44d3345f, 32'hc33d19f1, 32'hc0ed8383},
  {32'hc4685a2c, 32'hc22bed09, 32'hc1d16ae8},
  {32'h44e4f5ca, 32'hc3486b9e, 32'hc3563b9f},
  {32'hc5001dff, 32'hc32cc155, 32'hc247bb76},
  {32'h44727aea, 32'hc2466ce1, 32'h4203c685},
  {32'hc40fb044, 32'hc32797e9, 32'hc1413460},
  {32'h44f67994, 32'hc30dc189, 32'h42996f6d},
  {32'hc4e67ed3, 32'h43cb84a5, 32'hc23fa97a},
  {32'h44392fb9, 32'h40609893, 32'h42dbbe83},
  {32'hc4cc70ef, 32'hc3c1e098, 32'hc332fedd},
  {32'h4433b512, 32'hc363c131, 32'hc3808943},
  {32'hc34bae08, 32'hc3198588, 32'hc13d3334},
  {32'h43883678, 32'h4200d4ec, 32'hc24ea888},
  {32'hc48c1762, 32'hc3681e38, 32'h43a30e04},
  {32'h45014600, 32'hc2c752da, 32'hc2dba747},
  {32'hc4d1161e, 32'hc32b6cd4, 32'hc416f618},
  {32'h44eb1e22, 32'hc329ee21, 32'h42cc3b40},
  {32'hc3a97484, 32'h42da2aa6, 32'h43835436},
  {32'h444b9c26, 32'h43853550, 32'h437a86e0},
  {32'hc4917a94, 32'hc28f5d32, 32'hc2e878d9},
  {32'h44c1c317, 32'hc3c14c93, 32'h43662624},
  {32'hc4a70df7, 32'h431473e3, 32'hc41a0b8d},
  {32'h44eab000, 32'hc2bb582f, 32'h442469bf},
  {32'hc40480eb, 32'h3fd33ac0, 32'h4335838e},
  {32'h44202c9a, 32'hc373460d, 32'h4393e6e7},
  {32'hc357e9be, 32'hc32cf96c, 32'h421ca292},
  {32'h448c6a76, 32'h4201a4d4, 32'hc20eb2ff},
  {32'hc46b213d, 32'hc305bbc1, 32'hc37daa0c},
  {32'h449b8d21, 32'h43af85dc, 32'h43828be8},
  {32'hc503577c, 32'h43496813, 32'h41db86dc},
  {32'h44edbe07, 32'h4345a2f1, 32'h42f39c12},
  {32'hc4a02c0a, 32'hc220cbd4, 32'h417708e4},
  {32'h44eccbd5, 32'hc28d75f6, 32'hc1c60645},
  {32'hc4652715, 32'hc38dbd04, 32'hc2ad50a1},
  {32'h43e74e3c, 32'h40cf750d, 32'h42edb3e8},
  {32'hc4ba5dd5, 32'hc2dc500b, 32'h415f4fb5},
  {32'h43edd4ac, 32'hc3324339, 32'h42dbbd0e},
  {32'hc4eae664, 32'h422a281a, 32'hc1848c47},
  {32'h44aed384, 32'hc40e8770, 32'h4393c5fe},
  {32'hc439e8e6, 32'hc3bc0c5e, 32'h43533cd7},
  {32'h44c25b02, 32'hc2b3d591, 32'h42ed0dd7},
  {32'hc4f63726, 32'h42a8c9ec, 32'hc40934b5},
  {32'h4485555f, 32'hc187673f, 32'h43ff8d70},
  {32'hc38ed500, 32'h43212bb9, 32'hc295f2fc},
  {32'h4419252b, 32'hc218b61f, 32'h43468a69},
  {32'hc46e4e93, 32'hc2ee6f29, 32'hc322ca43},
  {32'h43f97ca8, 32'h430c1a7c, 32'h42733dd7},
  {32'hc4c1c95e, 32'h42d26ae0, 32'h4251a686},
  {32'h448ab286, 32'hc2f38bbc, 32'h43a5878d},
  {32'hc4ed00ea, 32'h42a9366b, 32'h4055bda8},
  {32'h44ad5476, 32'h41df4ab8, 32'h42c3b275},
  {32'hc45be975, 32'hc392c243, 32'hc289116e},
  {32'hc49c03c3, 32'hc35aaccb, 32'h431aa354},
  {32'h437b5c80, 32'hc3442aac, 32'h438606f4},
  {32'hc45a066e, 32'hc419b41b, 32'hc30870aa},
  {32'h44ac6eca, 32'hc308a85f, 32'h431d1db7},
  {32'hc46da57e, 32'hc3d883a7, 32'h410cfe6b},
  {32'h43e4a8b6, 32'h43941291, 32'hc332207a},
  {32'hc517e230, 32'h41635dc0, 32'hc30c8b86},
  {32'h446b5c1f, 32'h41c7cd0b, 32'hc2107716},
  {32'hc4c32ab9, 32'hc04580ce, 32'hc3017b1d},
  {32'h439a9730, 32'hc3e3490d, 32'hc2e46ea6},
  {32'hc3086d20, 32'hc376916e, 32'hc354d8a6},
  {32'h44a969f7, 32'h42e998d6, 32'hc32c8431},
  {32'hc4938187, 32'hc203d5f0, 32'h435fb219},
  {32'h44f29402, 32'h42097230, 32'h4270cfa2},
  {32'hc40d6199, 32'h42480147, 32'hc26ee9e3},
  {32'h43a05e0b, 32'h42c57121, 32'h42a45ff4},
  {32'hc4913916, 32'hc07652dc, 32'hc34df39f},
  {32'h44c537ed, 32'h433fa98d, 32'hc20c8a94},
  {32'hc42420de, 32'h43a1202c, 32'h4358e696},
  {32'h431efa68, 32'hc2aaf645, 32'h42cdf165},
  {32'hc32c45d8, 32'hc3d96e2c, 32'hc3d9b1cd},
  {32'h44f84adb, 32'h437254e9, 32'h440ed7d7},
  {32'hc515934a, 32'h429fcd06, 32'h438c77b6},
  {32'h448b826a, 32'hc32be60f, 32'h435ce6e0},
  {32'hc4843e68, 32'hc3b9b183, 32'hc381a4a6},
  {32'h4487b367, 32'hc2a5d76c, 32'hc2dffb4a},
  {32'hc38a7748, 32'hc2b52e93, 32'hc36b2021},
  {32'h4489afa0, 32'hc3939515, 32'hc2bfcbf3},
  {32'hc49ee26b, 32'h4336f430, 32'hc3f85022},
  {32'h443dd319, 32'hc3824562, 32'hc291eba3},
  {32'hc4111438, 32'h431458e0, 32'h42bbf12a},
  {32'h43dab1fc, 32'hc3bb567f, 32'hc1d4852e},
  {32'hc4fd4d5d, 32'hc3223520, 32'hc2b760a6},
  {32'h4502fe0e, 32'h43c1d451, 32'h429aaf2b},
  {32'h434e9d4e, 32'hc3f9f82b, 32'h41a46a1b},
  {32'h4473590e, 32'hc1fb87f7, 32'hc303d9eb},
  {32'hc319c290, 32'hc3578159, 32'hc3a7d028},
  {32'h44cca9ca, 32'h434f40e2, 32'h428bf0ea},
  {32'hc383fbb8, 32'hc2fd03cd, 32'h430ec397},
  {32'h44c9a39e, 32'h434645e7, 32'h4375bde9},
  {32'h4107caa6, 32'hc40fc983, 32'h43001c17},
  {32'h443883d5, 32'hc28df285, 32'h430ff1d1},
  {32'hc4a02b05, 32'hc238fdc6, 32'h437db410},
  {32'h44bdc9c0, 32'hc2b7dc71, 32'hc3c302ea},
  {32'hc44f70e8, 32'hc1a469ca, 32'hc2aa7ed4},
  {32'h44ac974c, 32'h43ceaaf4, 32'h41b13e51},
  {32'hc4cf1871, 32'hc3ce072f, 32'h435b74b8},
  {32'h4285a9d9, 32'h4083b883, 32'hc36fba84},
  {32'hc4cf2080, 32'h42edc302, 32'h4341382d},
  {32'h435133d0, 32'hc33323e6, 32'h4199cfc0},
  {32'hc4f2888c, 32'h435da5ed, 32'hc073d669},
  {32'h449f987a, 32'h42a63137, 32'hc2792d0b},
  {32'h4413de7a, 32'h4244f5d2, 32'hc22580c3},
  {32'h44119eea, 32'h42bfa58f, 32'h42eb8b55},
  {32'hc47fed62, 32'h43093b37, 32'hc1870aaa},
  {32'h446bb8e0, 32'h430254fd, 32'h4354c5b9},
  {32'hc4d6aa04, 32'hc3b15d81, 32'hc23e6366},
  {32'h44fddc8e, 32'hc3c63d9a, 32'hc37c3193},
  {32'hc4e9785a, 32'h438a02b4, 32'hc378b250},
  {32'h44bf9fd7, 32'hc30b2906, 32'hc1b0c21b},
  {32'hc4e09111, 32'hc3afb42c, 32'hc3036b57},
  {32'h449cfcd1, 32'hc2db0e3c, 32'h4371eb78},
  {32'hc4ac9d7f, 32'h4237214a, 32'hc38d7d6f},
  {32'h441e5ad6, 32'hc38fba43, 32'h421c7d1d},
  {32'hc3f689e4, 32'h4369e66b, 32'h428bffbd},
  {32'h433583d3, 32'hc3bdd2bd, 32'h42f45673},
  {32'hc3b226e8, 32'h42d487e7, 32'hc317c274},
  {32'h44f252a7, 32'hc29926ae, 32'hc318a77e},
  {32'hc3f7f3d0, 32'h43061acc, 32'hc3a50eaa},
  {32'h444d94dc, 32'h42d7fb6e, 32'h440deb33},
  {32'hc47d1a2e, 32'hc34b0a6e, 32'h433457cf},
  {32'h44b9f1f6, 32'hc333415e, 32'h42b74e31},
  {32'hc4fcc0dd, 32'hc232472a, 32'hc1e0b0dc},
  {32'h446b5eec, 32'h4387c93a, 32'hc1bb2a29},
  {32'hc50ca24c, 32'h436400f6, 32'hc316628b},
  {32'h44bdff31, 32'h43a3f8e8, 32'hc31e69d3},
  {32'hc4c00174, 32'h42a1cc72, 32'h41118584},
  {32'h44c80fac, 32'h4326c2cb, 32'h42a3b458},
  {32'hc482bca3, 32'hc3970264, 32'hc37506d5},
  {32'h435afbca, 32'hc2affca2, 32'h40e46a9a},
  {32'hc4aa031d, 32'hc3522a8a, 32'h432ac71c},
  {32'h44a14526, 32'hc3728150, 32'h4408903f},
  {32'hc4b847de, 32'h43e23e49, 32'h435cd4cc},
  {32'h448c492a, 32'h434ad8ea, 32'hc2f9953a},
  {32'hc4a84883, 32'h42e7fa23, 32'h437a3a99},
  {32'h44eeb19e, 32'hc3b8bbbe, 32'hc334935a},
  {32'h4410d3b1, 32'hc3a95a4d, 32'hc38604eb},
  {32'h441581de, 32'hc38d039c, 32'hc376dfe4},
  {32'hc5064787, 32'h43873c23, 32'h4180feba},
  {32'h4502ab1d, 32'hc2c9daed, 32'h42f9dd17},
  {32'hc4b6c431, 32'hc1cc3118, 32'h430403af},
  {32'h443602f4, 32'h432ab8d7, 32'hc2372d5f},
  {32'hc3c802fc, 32'hc34c7b9f, 32'h436ba3a3},
  {32'h450ba9fd, 32'h4271e1f0, 32'h435e95ae},
  {32'hc4b0755c, 32'h42a88e79, 32'hc4086466},
  {32'h44f60965, 32'h432cd9e9, 32'hc3c2f458},
  {32'hc2072900, 32'hc111cc0c, 32'h43141924},
  {32'h44135fc5, 32'h42a64acf, 32'h43400977},
  {32'hc4edbefe, 32'hc393d18c, 32'hc377938f},
  {32'h442a71f0, 32'h41f2b541, 32'h42ac6876},
  {32'hc289ba78, 32'h43251e78, 32'hc3122f19},
  {32'h44ef21ea, 32'hc3a4b9b8, 32'h42125963},
  {32'hc4b6d2ee, 32'hc28379a8, 32'h41a73fb2},
  {32'h44d29316, 32'h440b33b5, 32'hc2b3ec0c},
  {32'hc49d07df, 32'hc33b0515, 32'h44019469},
  {32'h448fb957, 32'h42b7323c, 32'h432fee5f},
  {32'hc48d90f9, 32'h4244597e, 32'h427e5b1f},
  {32'h44e538b1, 32'hc3857eca, 32'hc307dcaa},
  {32'hc4683e5d, 32'hc29ad78b, 32'hc1244c19},
  {32'h444b58d6, 32'hc29930dd, 32'hc329dd1d},
  {32'hc4903038, 32'hc2e65f45, 32'h4346834c},
  {32'h448b3230, 32'h435b175e, 32'hc3091716},
  {32'hc2415ab0, 32'hc3d37d6d, 32'h4385937f},
  {32'h438b5588, 32'h4384890e, 32'h4350f31f},
  {32'hc4c67b61, 32'h42e65252, 32'hc365af8d},
  {32'h44ce95a4, 32'hc3660155, 32'h43bbe7c0},
  {32'h41925f00, 32'hc3060966, 32'h43ab3be5},
  {32'h441ad3ac, 32'h42cf5e4a, 32'h44230466},
  {32'hc1c28580, 32'hc2ba951b, 32'hc344a07c},
  {32'h44df3597, 32'h434b8634, 32'h43b4e05e},
  {32'hc4cbed80, 32'h413ee184, 32'h42d5dc5b},
  {32'h44efa3d8, 32'hc348428f, 32'hc3714146},
  {32'hc48e8011, 32'h43484f34, 32'h43af47cb},
  {32'h450a43ab, 32'hc40f1c4b, 32'h42e92518},
  {32'hc4e28d21, 32'h43ca338a, 32'h430daafb},
  {32'h44d45e08, 32'h431da149, 32'hc3071498},
  {32'hc27c69f0, 32'h439a88a6, 32'h428a9fa7},
  {32'h4460b63e, 32'hc3e0a727, 32'h432bf889},
  {32'hc4d158f7, 32'hc238b411, 32'h42312906},
  {32'h44eca704, 32'h439fe319, 32'hc3822846},
  {32'h43dd9ff0, 32'hc305c7ad, 32'h43b621aa},
  {32'h43577270, 32'hc3000e40, 32'h43ec6c19},
  {32'hc5087a9a, 32'h41902d96, 32'h43b1b875},
  {32'h433ea3e0, 32'h435e378a, 32'h4319c81e},
  {32'hc4c77654, 32'hc33a6a78, 32'h44324155},
  {32'h443d95ce, 32'h42a1dda9, 32'h4245c240},
  {32'hc49764d8, 32'hc199c5cc, 32'h428e5ad6},
  {32'h44d3aefb, 32'h4384f739, 32'hc112ed6a},
  {32'hc4fbad46, 32'hc2b6c1bc, 32'h426f69b2},
  {32'h44eb76c6, 32'h4299d97b, 32'h42a064a8},
  {32'hc38e7cb0, 32'h425a3ed3, 32'h42a1e0a5},
  {32'h45156dee, 32'h42d4fe08, 32'hc3433fce},
  {32'hc44a3372, 32'hc32a4753, 32'h4308e711},
  {32'h44983cbb, 32'hc3e549da, 32'h4303ffe6},
  {32'hc4f3bf69, 32'hc38009e9, 32'hc1e93a62},
  {32'h45049781, 32'hc256b348, 32'h4314ad04},
  {32'hc4fbee77, 32'hc40aad0a, 32'h4386b3bf},
  {32'h445ca1ab, 32'hc30cbe7f, 32'hc31a2809},
  {32'hc452470c, 32'h42d9805f, 32'h43740db6},
  {32'h44910cfc, 32'h41e036a9, 32'hc25145f9},
  {32'hc423c80a, 32'hc33235aa, 32'hc32a3a43},
  {32'h43fe677c, 32'h4304f64a, 32'h4382ce68},
  {32'hc40f23e8, 32'hc1f37100, 32'hc3743cb1},
  {32'h4332b18f, 32'h4347fa58, 32'h434f0ea2},
  {32'hc4a47e46, 32'h426725d3, 32'hc339de44},
  {32'h44f11c51, 32'h41dafac0, 32'hc3629d7b},
  {32'hc4c37f62, 32'hc144698b, 32'hc3bc2c54},
  {32'hc3571e60, 32'hc291de31, 32'hc41c064a},
  {32'hc49c87a6, 32'hc3a77c2c, 32'hc3872c0b},
  {32'h438f683c, 32'h422f062a, 32'h439618e7},
  {32'hc4b6ac24, 32'hc1581aa0, 32'hc2f580e6},
  {32'h4484415c, 32'h432b9635, 32'hc37b4017},
  {32'hc453a6d6, 32'hc29ee7e7, 32'hc1678748},
  {32'h44a49610, 32'h42621a90, 32'hc27fe78e},
  {32'hc4293922, 32'hc3b038cc, 32'h43f517f2},
  {32'h450fe327, 32'hc2c7dd9d, 32'hc3e5e0cd},
  {32'hc48122d8, 32'h3f6a5220, 32'hc2aa4eaa},
  {32'h43d89710, 32'hc377b3de, 32'hc2ae593b},
  {32'hc4cc70dc, 32'h42f045e4, 32'h422a0691},
  {32'h44bee32b, 32'hc2df213e, 32'hc3382465},
  {32'hc50495cf, 32'h4397c968, 32'h43c245c5},
  {32'h446a959a, 32'h4203a9cf, 32'hc2e6e85f},
  {32'hc41b954f, 32'h40ec77e0, 32'hc1345dd1},
  {32'h4443da89, 32'h426f10da, 32'hc3d27360},
  {32'hc4e9d5fb, 32'hc1b79f8a, 32'hc3bb1ec2},
  {32'h428081a0, 32'h428e7b07, 32'h43481444},
  {32'hc4beef18, 32'h438fc3e9, 32'hc41aaa76},
  {32'h44da0aba, 32'hc1bcb3ce, 32'h42b63bbc},
  {32'hc3bbd09a, 32'h431b6fc0, 32'hc3ad4266},
  {32'h44576b96, 32'hc2f5634d, 32'h43f55fcc},
  {32'hc4b3357a, 32'hc237f576, 32'hc121ed88},
  {32'h45186c1d, 32'hc384c9ec, 32'hc31b7889},
  {32'hc325c15e, 32'hc342cb51, 32'hc3df9df3},
  {32'h44ffc182, 32'hc10f3b1b, 32'hc20e6e56},
  {32'hc4f0c427, 32'hc356115d, 32'h42443566},
  {32'h450207e7, 32'hc3af85d7, 32'hc26b4805},
  {32'hc46a5553, 32'hc3055cfa, 32'hc2ef6bdd},
  {32'h449d4f06, 32'h43de08a5, 32'h436570f2},
  {32'hc4f6af8e, 32'h43bf4b75, 32'h418e94e4},
  {32'h4417b7dc, 32'hc2d91e49, 32'hc383eb62},
  {32'hc4caa02c, 32'hc33d0c55, 32'hc3129efc},
  {32'h4499aaf1, 32'hc298a9b3, 32'h414696ea},
  {32'hc5054bb1, 32'hc39f7a9d, 32'h415f095c},
  {32'h45180432, 32'h4335d01b, 32'hc385c664},
  {32'hc4954a50, 32'h4338c85d, 32'h42ee88e0},
  {32'h43594c5a, 32'h42eb7d04, 32'h4214b402},
  {32'hc431fde3, 32'h42cabb2e, 32'h40fbcfb7},
  {32'h44ef03e0, 32'h43c623ab, 32'h43b0d1f2},
  {32'hc518cc82, 32'hc39093fa, 32'h437fe596},
  {32'h4461b0aa, 32'hc32984ea, 32'hc2be159a},
  {32'hc3deed10, 32'h42ebb36c, 32'h435e02e6},
  {32'h44e31466, 32'h41cc3845, 32'h4301b8ad},
  {32'hc3f7a766, 32'hc3cac0c1, 32'h43542d53},
  {32'h44fa34e8, 32'h43420876, 32'hc2071b76},
  {32'hc48e33d3, 32'hc2eeb4ef, 32'h43737d87},
  {32'h44e335d9, 32'h42d7b409, 32'h42b8b64a},
  {32'hc47a0f2e, 32'h43dab05b, 32'h430209f9},
  {32'h4480ba34, 32'hc3c40d7e, 32'h42dcdb3a},
  {32'hc38bef68, 32'hc35aba9a, 32'hc2aa313a},
  {32'h4484f4f3, 32'hc3cd9a91, 32'hc2a7fe0a},
  {32'hc4e03b0a, 32'hc3040be8, 32'h42ae9527},
  {32'h440a37e3, 32'h42eb5dc3, 32'h42b09f89},
  {32'hc4bf990e, 32'h42138357, 32'h43ab522d},
  {32'h4451671c, 32'hc3a81178, 32'h42c7f5a2},
  {32'hc37289ac, 32'h42db73ef, 32'h421ce807},
  {32'h44d6b625, 32'hc32f34d9, 32'h43032e80},
  {32'hc506abbc, 32'hc3414399, 32'hc3860541},
  {32'h43d61778, 32'hc2d9e9f5, 32'hc2d8fc91},
  {32'hc3ceb980, 32'hc21d2331, 32'h432ff4f6},
  {32'h43b20d2c, 32'hc33d066f, 32'h43c5cd83},
  {32'hc3fae735, 32'hc29b4526, 32'h41b8d684},
  {32'h441714ea, 32'h4304e58e, 32'h43b6fc49},
  {32'hc4e45297, 32'h439cfe7e, 32'hc336ef76},
  {32'h43828d92, 32'h43bf33ab, 32'h42d7d464},
  {32'hc4880395, 32'h43883803, 32'h421ef284},
  {32'h433c0a68, 32'h43b55642, 32'hc222cd19},
  {32'hc4a5da0e, 32'hc245942d, 32'h41539c5e},
  {32'hc3d38514, 32'hc27858af, 32'hc3a6a02c},
  {32'hc4adb60c, 32'hc3049e1b, 32'h4383b942},
  {32'h441f841a, 32'h429fd5c3, 32'hc3aaa61c},
  {32'hc4139a64, 32'h42adc9b6, 32'hc2e7c4e3},
  {32'h440f5766, 32'hc3889e18, 32'h42f92893},
  {32'hc514c6f7, 32'hc2afb68f, 32'h42b74f37},
  {32'h4431228c, 32'h3fe3b6a0, 32'h415c4a78},
  {32'hc442a653, 32'hc2a4d5a7, 32'hc2882fd3},
  {32'h4509e6f4, 32'h432c60c8, 32'hc2a45107},
  {32'hc5079922, 32'hc35f6c9d, 32'hc3e6d5d2},
  {32'h44790476, 32'h4343e807, 32'hc285af91},
  {32'hc386e79c, 32'hc2c8cd22, 32'hc239a0cc},
  {32'h44808b1d, 32'h44138622, 32'h43fcc344},
  {32'hc502ac4b, 32'h4407322b, 32'hc2a04ab0},
  {32'h44c33b1e, 32'hc3fbde4d, 32'hc39b1eff},
  {32'hc281a6e0, 32'hc1ad6df6, 32'h438e96aa},
  {32'h44696904, 32'hc39646ef, 32'h432026f0},
  {32'hc4d21ac7, 32'hc306c3fe, 32'hc3496bf1},
  {32'h451069bd, 32'h418f5bd4, 32'hc2b44a17},
  {32'hc4d6ce28, 32'h43669480, 32'hc2b90bf0},
  {32'h44ea8940, 32'hc394bd71, 32'hc0bc2d70},
  {32'hc4ec2871, 32'h43574a6d, 32'hc3fa6a9e},
  {32'h4384d360, 32'hc3e6a447, 32'hc41eb9ff},
  {32'hc47a6e16, 32'hc1ab1f74, 32'h431dd356},
  {32'h44e1a489, 32'h437b2d88, 32'hbfcfd540},
  {32'hc3a52ee4, 32'hc3dbe955, 32'h439f1b66},
  {32'h44e9b471, 32'hc340827f, 32'hc19bb715},
  {32'hc4dac5c0, 32'hc36a078c, 32'h43166e1b},
  {32'h4424a27c, 32'h43e0cc3e, 32'h434b9b17},
  {32'hc4045222, 32'hc393c63e, 32'h41fb40f2},
  {32'h4402ae5d, 32'h43c12fcc, 32'h43da5f00},
  {32'hc504f3e8, 32'h429aa8d1, 32'hc38bdf1b},
  {32'h4382ddf7, 32'h4312e775, 32'h438837d1},
  {32'hc46ff3b2, 32'h423f9272, 32'hc31e39b9},
  {32'h43d20801, 32'h4397e611, 32'hc2e89433},
  {32'hc4f5c79c, 32'h434ea9cb, 32'h43325b23},
  {32'h43bac4b4, 32'hc334bf8f, 32'h431f82e0},
  {32'hc492b238, 32'hc233d3df, 32'hc0a60bf6},
  {32'h44c85658, 32'h43b4464c, 32'h436bf226},
  {32'hc4e07d76, 32'h435b6b69, 32'h421f1ef6},
  {32'h450d652b, 32'hc2f86c0e, 32'hc3320aaa},
  {32'hc3cf91f7, 32'h434241ba, 32'h42b1e981},
  {32'h44f9b490, 32'hc359a40f, 32'h42193792},
  {32'hc458af68, 32'hc1e10248, 32'h440aa541},
  {32'h45007023, 32'h4361a5fe, 32'hc234c65b},
  {32'hc417debc, 32'h43baa7cc, 32'h4339adb7},
  {32'hc1a99208, 32'hc328073c, 32'h42fc0a17},
  {32'hc0b75b80, 32'hc3476001, 32'hc382c850},
  {32'h44cd7f14, 32'h40ed9873, 32'hc33c9b1d},
  {32'hc4e191d0, 32'hc3dab8ff, 32'h43528def},
  {32'h44fe53b8, 32'h4220d326, 32'h433907a0},
  {32'hc48c881b, 32'h42a7fbab, 32'hc30d5d81},
  {32'h44187dcc, 32'h4316511d, 32'hc268497e},
  {32'hc4952ad7, 32'h441de075, 32'hc2e43cbe},
  {32'h413b7300, 32'hc39c70eb, 32'hc36d2a4d},
  {32'hc4270380, 32'hc219ef4c, 32'hc391b1f1},
  {32'h45163536, 32'h412fbd29, 32'h40c0a3c8},
  {32'hc48d336a, 32'hc2b45992, 32'hc32fa352},
  {32'h44da5035, 32'h43121fd2, 32'h4361dcc1},
  {32'hc46a18aa, 32'h43368019, 32'hc26e8eea},
  {32'h4453b022, 32'hc29fc4bd, 32'hc2c8a4e2},
  {32'hc38a82a6, 32'hc3c107df, 32'hc255fc7e},
  {32'h44a86a64, 32'h42a8b164, 32'h4384b241},
  {32'hc444afac, 32'h4236f472, 32'hc35d1dea},
  {32'h4362702f, 32'h435eada8, 32'h41229b2f},
  {32'hc3a58019, 32'hc28f9ae4, 32'hc07f97ff},
  {32'h449c6826, 32'hc38967f1, 32'h4222f83b},
  {32'hc4296a7c, 32'hc3744fd7, 32'hc27316c6},
  {32'h43858727, 32'hc390259d, 32'h42ad3a78},
  {32'hc4535710, 32'h425dbb00, 32'hc27f6f09},
  {32'h448ea425, 32'hc082a8d1, 32'h438517c9},
  {32'hc48e3cf4, 32'h4398fe03, 32'h4377b152},
  {32'h44c4cee8, 32'h42e46b2f, 32'hc361e64e},
  {32'hc502fabf, 32'hc24ce6d1, 32'hc358cda0},
  {32'h44aaaf2c, 32'hc1f7d071, 32'hc3c7b0bf},
  {32'hc51e0ea2, 32'hc31b226e, 32'h41c92aa8},
  {32'h450c222c, 32'hc398aa51, 32'h427b589c},
  {32'hc51aa065, 32'h43588c67, 32'h434ccf38},
  {32'h448e9291, 32'h42039702, 32'hc2344670},
  {32'hc50f950f, 32'hc38d90f3, 32'h42b56cb6},
  {32'h451776b2, 32'hc2dac4a0, 32'hc2d8f3b1},
  {32'hc3ad43ec, 32'hc39ca135, 32'h4339d502},
  {32'h45103591, 32'h43cbc964, 32'h43cfff95},
  {32'h41fd914a, 32'hc370dc45, 32'hc04a038c},
  {32'h446ca600, 32'hc3030fe4, 32'h42ed6067},
  {32'hc51ad15a, 32'hc2b90d14, 32'hc2d983be},
  {32'h43b3d860, 32'h42e7801e, 32'h43962957},
  {32'hc4e6810a, 32'hc1e27892, 32'hc2e7241b},
  {32'h43e03784, 32'h428e85a8, 32'h43a1bd61},
  {32'hc3a1112c, 32'h439720d4, 32'hc3205408},
  {32'h44ec9eba, 32'hc3269c20, 32'hc2bcd319},
  {32'hc45677ea, 32'hc346599c, 32'hc2bcb4cb},
  {32'h45354da2, 32'h427e3629, 32'h4281056b},
  {32'hc47ebcac, 32'h42255f1e, 32'hc312de96},
  {32'h45075b90, 32'hc34201f3, 32'h425af72f},
  {32'hc4dc6bc8, 32'h42ff4260, 32'hc36ef915},
  {32'h4366960d, 32'h433d0da2, 32'h43c11c6f},
  {32'hc49fd2dc, 32'hc2fcc574, 32'h428cf9a4},
  {32'h444d40da, 32'h43969019, 32'hc2936913},
  {32'hc45dce90, 32'hc4077feb, 32'hc40aa277},
  {32'h4471f7fd, 32'hc1c27834, 32'h432a4119},
  {32'hc503ff2c, 32'hc1086fdb, 32'h41f93e5f},
  {32'h4485eb6a, 32'h42639ed2, 32'h421b66ba},
  {32'hc39bf528, 32'hc387ec40, 32'h42bf43f7},
  {32'h44db4b85, 32'hc376c1f1, 32'h4397ad9a},
  {32'hc4e13308, 32'h43e8e1b2, 32'hc3590a29},
  {32'h450ebb22, 32'hc31b9dcf, 32'h423a0834},
  {32'hc4030404, 32'h4360fd5c, 32'hc1c72f56},
  {32'h44b40ba9, 32'h42549d91, 32'h42ec99d1},
  {32'hc48e91f8, 32'hc237f20b, 32'h4380e1e7},
  {32'h45127c04, 32'h4282a5fa, 32'h42348202},
  {32'hc4fd4661, 32'hc3f0d19e, 32'h435eab4c},
  {32'h45274093, 32'h42e2c56a, 32'h42e3cd73},
  {32'hc4b59dbd, 32'hc1b5d6d2, 32'hc3300e06},
  {32'h44cac5d8, 32'hc0a2b120, 32'hc3bd3f62},
  {32'hc4b4e884, 32'h439300a8, 32'h42e486b1},
  {32'h4471e32f, 32'hc2e83c15, 32'h43332c03},
  {32'hc42f340e, 32'hc28cd0e8, 32'hc30f46a5},
  {32'h44a74433, 32'h42fa7570, 32'h426e74c8},
  {32'h421b455c, 32'h4319d8e5, 32'hc1eb8de9},
  {32'h44c4308f, 32'hc2639b69, 32'hc2fbb1b4},
  {32'hc506f9e8, 32'hc251312d, 32'hc0bbb9e7},
  {32'h44bc867c, 32'hc3c03baa, 32'hc3848092},
  {32'hc498c5f2, 32'hc2af4dd0, 32'h43ca99b1},
  {32'h4391a885, 32'hc40307fc, 32'h435ce600},
  {32'hc4f2c8c0, 32'hc2ad0061, 32'h440ac7c6},
  {32'h438ace30, 32'hc3f4bffa, 32'hc23d17a6},
  {32'hc4793d56, 32'h3f8523c5, 32'hc21132fe},
  {32'h452bbdc7, 32'hc3746a0c, 32'hc3b354e7},
  {32'hc510a7a8, 32'h435de8e3, 32'hc396ef67},
  {32'h44cded65, 32'hc2a839e4, 32'hc2939fb5},
  {32'hc42d33a0, 32'h42a34d0b, 32'hc3e691e0},
  {32'h4512ed20, 32'hc3489d15, 32'h43857b08},
  {32'hc394637c, 32'hc314c79c, 32'h425ce533},
  {32'h4493b1ad, 32'h4340cac7, 32'hc315efb9},
  {32'hc3b5c342, 32'hc11a5d52, 32'hc35daf1b},
  {32'h44dc82b9, 32'h435982aa, 32'h43910ace},
  {32'hc47511b1, 32'hc28f0501, 32'h41c5debe},
  {32'h4509dc54, 32'h4287b72a, 32'h4207caa1},
  {32'hc4b08254, 32'h429b57d7, 32'h40aa63ea},
  {32'h450946fd, 32'hc26f6783, 32'hc288d016},
  {32'hc2978b10, 32'h430e2692, 32'h4355d407},
  {32'h44e18b01, 32'h4265301f, 32'h43a4ab49},
  {32'hc512e0f3, 32'h4373189c, 32'hc2ae136b},
  {32'h44897828, 32'hc291fcff, 32'hc3cdae64},
  {32'hc4d79209, 32'hc34d2c1e, 32'hc3212631},
  {32'h44a12a81, 32'hc3abad26, 32'hc1390e12},
  {32'hc4dbfd96, 32'hc252e3ec, 32'h4316f6fe},
  {32'h452e50a1, 32'h441d3e85, 32'h4314ea70},
  {32'hc4eb5326, 32'h43645a7a, 32'h43a95bcd},
  {32'h440a00c6, 32'hc31d409a, 32'h44189b18},
  {32'hc41728f2, 32'h43afc35b, 32'hc2582fbd},
  {32'h450eac8b, 32'h43525f90, 32'h43fb3bb4},
  {32'hc4aa53d4, 32'h42fb4079, 32'hc22258b8},
  {32'h44bccf1d, 32'h439fb7e5, 32'hc33f8661},
  {32'hc47edaa3, 32'hc3ce0b58, 32'h42f8b6ef},
  {32'h44b949ee, 32'hc282bb12, 32'hc328d923},
  {32'hc3cf9c30, 32'h42cb9fce, 32'h40a69fd0},
  {32'h4446a2f7, 32'hc34c0d11, 32'hc36c4ca2},
  {32'hc4378986, 32'hc2aa27fc, 32'hc24fc289},
  {32'h43cfd338, 32'hc3665752, 32'h439b768f},
  {32'hc42e0e7a, 32'hc3b3529b, 32'hc33e68e9},
  {32'h450e1e28, 32'h43cea33a, 32'hc14217fd},
  {32'hc4d9e9b2, 32'h42571f6c, 32'hc21a4aa6},
  {32'h4518d532, 32'hc38dac6d, 32'hc2e2faec},
  {32'hc4d3e3b9, 32'h43457e4a, 32'h435086f6},
  {32'h438b2ddc, 32'h43b4868b, 32'h426538fa},
  {32'h431f12c8, 32'hc1241136, 32'hc24b724d},
  {32'h441030e4, 32'h43155c56, 32'hc3d8d698},
  {32'hc4bc9d51, 32'h3ecd4b02, 32'hc32a7737},
  {32'h450c463a, 32'h42ff541a, 32'hc3020168},
  {32'hc43d875f, 32'hc38bb8a4, 32'h434203cf},
  {32'h44e84821, 32'hc30e4b34, 32'hc1c16545},
  {32'hc4a299ae, 32'h4229eac7, 32'h40ccd592},
  {32'h450d9053, 32'h439840be, 32'hc3b5c6b2},
  {32'hc460dd0e, 32'hc1cfc59b, 32'h435b4968},
  {32'h450486cd, 32'h425567f2, 32'h43173c3a},
  {32'hc4b78434, 32'hc28ce2d2, 32'h431d8a48},
  {32'h44b7689d, 32'h41eebf98, 32'h3ea1f9a7},
  {32'hc49fd071, 32'hc353b19e, 32'h42fc5320},
  {32'h44c142a9, 32'h4318773c, 32'hc3d3be82},
  {32'hc3a5b29a, 32'h429c95e0, 32'h438ed062},
  {32'h43c9eabb, 32'h4029b635, 32'hc3c1d9b4},
  {32'hc46dae8a, 32'h42de2a66, 32'h41e4cfe0},
  {32'h44c9c5d5, 32'h43516428, 32'hc3c7204d},
  {32'hc4844a39, 32'hc2da721d, 32'hc2ac43ea},
  {32'h44e356cc, 32'h4371f86f, 32'h4300eeec},
  {32'hc4cdba0c, 32'hc33b774e, 32'h430431b5},
  {32'h44a3e4de, 32'h433e1c5e, 32'hc3431ab4},
  {32'hc5047e36, 32'h41f02ffc, 32'h43aab57f},
  {32'h44d72f38, 32'h42e0d0f2, 32'hc193d692},
  {32'hc4fc0043, 32'hc3152ced, 32'hc2a329c6},
  {32'h4382ec5c, 32'h43e5dce1, 32'hc391e077},
  {32'hc36fd260, 32'hc3035f30, 32'h43afdd93},
  {32'h4445e856, 32'h4195b69b, 32'h42fa96b5},
  {32'h41b1d41e, 32'h41aa1e80, 32'h43a239a4},
  {32'h44de4e77, 32'hc3681156, 32'hc1a0dc30},
  {32'hc47dc132, 32'h42c05674, 32'h430be9a4},
  {32'h44c0edfe, 32'h42e82742, 32'hc37e1480},
  {32'hc4a89220, 32'hc41463eb, 32'hc31e4b11},
  {32'h44d7bd13, 32'h42d91a05, 32'hc26b3742},
  {32'hc4f9b25f, 32'h436f828e, 32'h439c2a6f},
  {32'h44abf60d, 32'hc3bbdd6a, 32'hc42366df},
  {32'hc4af9fdb, 32'hc29bc942, 32'hc2e53330},
  {32'h444bc8e0, 32'h43d09af8, 32'hc34ee75f},
  {32'h446d9c7c, 32'hc3326502, 32'hc2b03c44},
  {32'hc4549596, 32'h43c9257d, 32'hc2ff85dd},
  {32'h43dfe8e2, 32'hc338f517, 32'h42b968ea},
  {32'hc4d880fa, 32'hc3377621, 32'hc365bb03},
  {32'h43ef79c4, 32'h434b5ec9, 32'hc39017e9},
  {32'hc4affc72, 32'h43606241, 32'hc20e37c7},
  {32'h44cd327b, 32'hc264812c, 32'hc27d40a2},
  {32'hc4fe8b20, 32'hc423c8f6, 32'h439e98df},
  {32'h44bb1832, 32'hc3298d6a, 32'hc2ae079c},
  {32'hc3902322, 32'h438355cc, 32'h4325ce97},
  {32'h44fe3ec4, 32'hc3838e41, 32'h432a4aef},
  {32'hc3718628, 32'hc404d347, 32'hc40fbafa},
  {32'h45089bf6, 32'h43d1e137, 32'hc204b888},
  {32'hc30baba0, 32'hc35c9269, 32'hc2adb8a0},
  {32'h447cce96, 32'hc32e97e4, 32'h42b932a4},
  {32'hc50e2849, 32'h41283bf2, 32'hc231697f},
  {32'h4487b05d, 32'h43d6dc47, 32'hc2cbbc84},
  {32'hc50a0bf4, 32'h440f8cd5, 32'hc226165e},
  {32'h445938ac, 32'h43a4650e, 32'hc204e4bf},
  {32'hc515a261, 32'h439a7035, 32'hc32aa7f6},
  {32'h44ce32ce, 32'h43026c18, 32'hc212e8c0},
  {32'hc45fce41, 32'h42cbaa8d, 32'h42d5dba5},
  {32'h450288ce, 32'hc37848c7, 32'h42fb248b},
  {32'hc196fda0, 32'h4358605d, 32'hc08f3027},
  {32'h44fc9763, 32'hc370c8c8, 32'h427cc6fa},
  {32'hc430de48, 32'h43eab72d, 32'h434c9be0},
  {32'h44d5cead, 32'hc29a9753, 32'h42e63250},
  {32'hc3ffff37, 32'hc34264e1, 32'h43bdcb26},
  {32'h435476bc, 32'h43bb2692, 32'hc22aa348},
  {32'hc4c90e97, 32'h42915143, 32'h43c60095},
  {32'h445b234c, 32'h41d920fb, 32'hc3e05440},
  {32'hc47d6694, 32'hc3e9e49c, 32'h43e9636b},
  {32'h449de859, 32'h42b67d0f, 32'hc3177e06},
  {32'hc48145bb, 32'hc2af7d32, 32'hc382a173},
  {32'h44ee04bd, 32'h430ab714, 32'hc18ca6c2},
  {32'hc4ef20fe, 32'hc3c1964d, 32'h42ab7625},
  {32'h4508704e, 32'hc3680683, 32'h43146149},
  {32'hc4ae3094, 32'h43330d72, 32'h43b94521},
  {32'h44d7b67e, 32'hc39cee22, 32'hc3006ef3},
  {32'hc48c8001, 32'h438fb824, 32'h43ab6816},
  {32'h4514709b, 32'hc38c34da, 32'h417be59c},
  {32'hc492ced6, 32'hc2bec681, 32'h406cbd24},
  {32'h44077c1a, 32'hc3d082bd, 32'h41bb9929},
  {32'h4290f660, 32'hc3627ed1, 32'hc304aedd},
  {32'h451b317c, 32'hc2a3dd7e, 32'h430904e8},
  {32'hc39128d2, 32'h43ae8eab, 32'h42c9e22a},
  {32'h44d8445f, 32'h4333da93, 32'hc20e27a0},
  {32'hc4c0a8a7, 32'hc3b4c091, 32'h4229a436},
  {32'h44fe5942, 32'h409fb65b, 32'h42ac3c80},
  {32'hc4faea10, 32'hc100c5f8, 32'h41e92e51},
  {32'h4496e09e, 32'h43c8a868, 32'hc3eb2b39},
  {32'hc49d70fe, 32'hc386c257, 32'hc35eb2bb},
  {32'h44675d32, 32'h42a16928, 32'hc275f10f},
  {32'hc38c95a4, 32'h432dd3c7, 32'hc1dbc717},
  {32'h448f3a18, 32'hc2a44975, 32'hc2b190bf},
  {32'hc506fb19, 32'hc320947c, 32'hc3268010},
  {32'h44d4873c, 32'hc37d34a0, 32'hc23ed003},
  {32'hc5096171, 32'hc206ea27, 32'hc3570dad},
  {32'h441dfd0f, 32'h43b83f67, 32'hc12280ec},
  {32'hc154a800, 32'hc302a39e, 32'hc2d4591c},
  {32'h44c3f480, 32'hc3a97050, 32'h4311d425},
  {32'hc4b3fcef, 32'h439deff0, 32'h435e0900},
  {32'h43e6e23e, 32'hc3a4c8e7, 32'hbfc4cbae},
  {32'h42a7b8c0, 32'h42ed202d, 32'h427d17dd},
  {32'h430aa188, 32'hc2c8421b, 32'h4367c3f5},
  {32'hc50c4b7b, 32'hc3013420, 32'h429b3f48},
  {32'h450a618b, 32'h42972c2d, 32'hc3147d79},
  {32'hc4da15db, 32'hc33812ae, 32'h436d4403},
  {32'h450f2454, 32'h4363040d, 32'h43991acb},
  {32'hc5053c87, 32'hc3b239ea, 32'hc2ab3f4e},
  {32'h45021389, 32'h4386e898, 32'hbfe2ca10},
  {32'hc40ab438, 32'hc3bf6b6f, 32'h43e9899b},
  {32'h44c80661, 32'hc29bd8b6, 32'h43469c71},
  {32'hc4c42814, 32'h43899325, 32'h42c10722},
  {32'h44fac622, 32'hc3508591, 32'h430bec92},
  {32'hc5033348, 32'h43b8fdd6, 32'hc37a8e20},
  {32'h43f7d46c, 32'h4114cd35, 32'h4305b044},
  {32'hc3a7ab10, 32'hc333aa3e, 32'h42b03db0},
  {32'h45171d4a, 32'h433faad3, 32'h4303d219},
  {32'hc515ded3, 32'hbfcb9630, 32'hc2fc4e2d},
  {32'h4191bac0, 32'hbed8ef40, 32'h43e79597},
  {32'hc4eb60d8, 32'h43eb4c33, 32'h42bc9395},
  {32'h449618ba, 32'hc325148e, 32'h43b79a23},
  {32'h430099b0, 32'h437f68ca, 32'h437e8ec7},
  {32'h44842657, 32'h42abc4b5, 32'h42df3c09},
  {32'h406c7c00, 32'h425ee112, 32'h42523d38},
  {32'h444edf94, 32'h4403ade4, 32'h41a18650},
  {32'hc4cae200, 32'hc2d50fe3, 32'hc2740672},
  {32'h45010d36, 32'hc199542c, 32'hc3868246},
  {32'hc4fdca07, 32'hc3aca827, 32'hc380faae},
  {32'h451a5c4b, 32'h430fecee, 32'hc1bc78fc},
  {32'hc4ef5f86, 32'hc3610b95, 32'h4323ef52},
  {32'h4503b95b, 32'h429a2068, 32'h43db064e},
  {32'hc4b2592b, 32'hc2273df2, 32'hc2da22f1},
  {32'h43d9178e, 32'h43964770, 32'h437d1d82},
  {32'hc3c12000, 32'hc3094d74, 32'h42d21031},
  {32'h44c22d31, 32'h430196d3, 32'h428aab05},
  {32'hc4f8d3bc, 32'hc2aa5de6, 32'h42e9a91a},
  {32'h42f97a88, 32'h437b4acc, 32'hc387608e},
  {32'hc4ab9c15, 32'hc3a0c154, 32'h43278382},
  {32'h450a4f5f, 32'hc39a691e, 32'h41c0a77e},
  {32'hc489524a, 32'h434b2b05, 32'hc34933d2},
  {32'h440e67e0, 32'hc3e7f4cf, 32'hc25051f2},
  {32'hc4f97226, 32'hc24d557a, 32'h439cb3d1},
  {32'h448cc2e7, 32'h43d76fae, 32'h42bc54e5},
  {32'hc4a5de84, 32'hc35d5bef, 32'hc1ff2db2},
  {32'h43f930a8, 32'hc34f7f81, 32'hc2a74d1a},
  {32'hc42000f8, 32'hc390e9f1, 32'hc22ff8ad},
  {32'h4436d9dc, 32'hc2d8c7c2, 32'hc3682182},
  {32'hc4556816, 32'h42283d86, 32'h435c0c25},
  {32'h43921baf, 32'hc3debaf2, 32'hc38c0a9a},
  {32'hc39f27b0, 32'h43864be5, 32'hc23d1537},
  {32'h43c8cd82, 32'h423bfeca, 32'hc2ea8cff},
  {32'hc51536aa, 32'hc2d3bb48, 32'hc333c1d3},
  {32'h44e14938, 32'hc2c7adfa, 32'h43157c75},
  {32'hc502ae38, 32'hc342ee51, 32'h438c9175},
  {32'h43c07524, 32'hc3975dca, 32'h4375878e},
  {32'hc4c33838, 32'hc3e87966, 32'hc334683c},
  {32'h43808390, 32'h436cda39, 32'h43e7a6a0},
  {32'hc3101e50, 32'hc28f0e44, 32'hc2d01874},
  {32'h44dc4bdf, 32'h43e83eae, 32'hc34c54fc},
  {32'hc475c566, 32'hc21252fd, 32'h428c4521},
  {32'h430814a8, 32'hc1b1a8d8, 32'h43708660},
  {32'hc4208975, 32'h434f4b1f, 32'hc2e6862c},
  {32'h44f3a061, 32'h412ed372, 32'hc3e7e6ec},
  {32'hc4f1bdc3, 32'hc321c329, 32'h42d30316},
  {32'h44d2870c, 32'hc229431e, 32'h430aa564},
  {32'hc5155e8e, 32'h440aee92, 32'h41efc017},
  {32'h4482d4fb, 32'hc3362702, 32'h43e11877},
  {32'hc4b085d8, 32'h40d9ccda, 32'h438e4ae2},
  {32'h448d0370, 32'h43534a53, 32'h435b7440},
  {32'hc4fddf02, 32'h42905dd4, 32'h43a05665},
  {32'h43ce2598, 32'hc228a3a9, 32'h43c83eec},
  {32'hc4a6fbfd, 32'h437dcc3a, 32'h434d35ca},
  {32'h4420e68e, 32'hc21a9c20, 32'hc1e14813},
  {32'hc4fb5667, 32'hc38191b6, 32'h41c75dd5},
  {32'h44d44ae3, 32'hc2a0ad83, 32'hc2c74d7d},
  {32'hc3cc4f94, 32'hc24372d4, 32'h4307fa29},
  {32'h44f26bc2, 32'hc3b3ecd5, 32'hc1761584},
  {32'hc4f398e8, 32'h43333757, 32'hc3873f1e},
  {32'h44c6c818, 32'hc3b08333, 32'hc31e983a},
  {32'hc4a708a1, 32'hc1b05276, 32'hc39c4bec},
  {32'hc304b518, 32'hc2b9f67c, 32'h4323789a},
  {32'hc4cb9d08, 32'hc38350d1, 32'hc2b2e571},
  {32'h44fc87c1, 32'hc3052062, 32'h42e53668},
  {32'hc4bcea10, 32'h42bcdf41, 32'h417cec71},
  {32'h4347bce0, 32'hc3d459f2, 32'h43921b1b},
  {32'hc29a9722, 32'h432780a5, 32'hc30410a6},
  {32'hc010d800, 32'hc1bdb5bc, 32'h41817700},
  {32'hc3d2c7fc, 32'h43d0b757, 32'hc2752836},
  {32'h43d73e60, 32'hc306aa38, 32'h41bb1034},
  {32'hc4893636, 32'hc21871ea, 32'h42475028},
  {32'h450f3072, 32'h43b40a61, 32'h42380321},
  {32'hc4d4272b, 32'h4206a334, 32'hc38946bc},
  {32'h44adcbf2, 32'h43421520, 32'hc2a168c5},
  {32'hc4991280, 32'h42186e8f, 32'h4185bc20},
  {32'hc2091290, 32'hc2c2a4f3, 32'h43060b71},
  {32'hc44a9df5, 32'h4357984a, 32'h4105c5fa},
  {32'h4487fbb0, 32'hc2996b00, 32'hc3f92cf0},
  {32'hc3f71452, 32'hc3511157, 32'h42a71dd8},
  {32'h45089620, 32'h42b447d7, 32'h432f3d5a},
  {32'hc4f21c8e, 32'hc1d5d600, 32'hc3119a73},
  {32'h4502096a, 32'hc319bd00, 32'h41bb674a},
  {32'hc480f910, 32'h435b9980, 32'hc2236bf2},
  {32'h450bb559, 32'h430a6276, 32'h4299c820},
  {32'hc49a11e0, 32'hc1ce53f2, 32'hc3339674},
  {32'h442446b5, 32'h410285d8, 32'h42e8d293},
  {32'hc458b62e, 32'hc1f44710, 32'hc32f08c1},
  {32'h44639576, 32'h4393b486, 32'hc260dcfa},
  {32'hc5091bd1, 32'h42fca0a2, 32'hc32ef6cb},
  {32'h44f4f06c, 32'h4321be7a, 32'hc36835c7},
  {32'hc4624cc7, 32'h41713c77, 32'hc3812014},
  {32'h4506786f, 32'h43ab2c7a, 32'hc21394c0},
  {32'hc47fd58e, 32'hc2819e81, 32'hc3851fc1},
  {32'h44358014, 32'hc3085af7, 32'h436ffbcc},
  {32'hc4b752c4, 32'hc16f1b9f, 32'h434db67a},
  {32'h44e1a5ff, 32'h4246f5a5, 32'h4284df43},
  {32'hc4911bc0, 32'h431cddd5, 32'hc19d6dba},
  {32'h44ef9a36, 32'hc35db0b1, 32'h42f930c1},
  {32'hc4fff211, 32'hc3c1525b, 32'hc361cc34},
  {32'h4488f20c, 32'h4331f1e3, 32'hc3ec6f7a},
  {32'hc495e9fa, 32'hc33a73ad, 32'hc2e1e1ac},
  {32'h44d7c61e, 32'hc19771c2, 32'h43decd54},
  {32'hc4dd67f0, 32'hc3b93cd7, 32'h438d5752},
  {32'h4486be5f, 32'hc370d05c, 32'hc3b204f9},
  {32'hc4adcc76, 32'h4337c11a, 32'h42cf9fd1},
  {32'h43c08c98, 32'hc190f71d, 32'hc343a4ea},
  {32'hc4ec3a74, 32'hc1d2ad3d, 32'hc29b6ace},
  {32'h43f948c8, 32'h419aa888, 32'hc0846b62},
  {32'hc4ca3e49, 32'h4394e968, 32'h43303269},
  {32'h448f3b2d, 32'h4321df83, 32'hc28c3584},
  {32'hc4b336dd, 32'h41806d21, 32'hc30bdca1},
  {32'h44b3333f, 32'h4331a1ce, 32'h43c97a15},
  {32'hc48255df, 32'hc32827d4, 32'h4363fb25},
  {32'h446a975c, 32'hc2c2aa20, 32'h4395232c},
  {32'hc429abe6, 32'hc242d7ed, 32'h41e2e4c6},
  {32'h4413ba1b, 32'hc1dbba7c, 32'hc2a88ded},
  {32'hc41febe7, 32'hc415573e, 32'hc2a9eeae},
  {32'h44ad4c48, 32'h4295c4d7, 32'h431352be},
  {32'hc4cc8232, 32'hc36158b1, 32'h43c2dea7},
  {32'h44ed6825, 32'h430024f8, 32'h43f842ca},
  {32'hc49738d2, 32'h4369b808, 32'hc1e38d90},
  {32'h4485cb2b, 32'hc354119b, 32'hc321b34c},
  {32'hc4a1deda, 32'hc38ece0d, 32'hc31868c1},
  {32'h44ad15f3, 32'hc3936332, 32'h4313c5e6},
  {32'hc3ba2458, 32'h43a4bfbd, 32'h433140ab},
  {32'h44d90b6e, 32'hc3be9cc3, 32'h43d8744c},
  {32'hc43c557e, 32'hc38a1d46, 32'hc40e9dd2},
  {32'h44dc6840, 32'hc3b78cdf, 32'h43a45093},
  {32'hc4d647df, 32'hc3214fe0, 32'h43854cca},
  {32'h4364c810, 32'hc3227217, 32'h43a277c3},
  {32'hc496672e, 32'h43151fea, 32'h43bab1d9},
  {32'h423abba0, 32'h43b83e09, 32'hc3cce33a},
  {32'hc4823a02, 32'hc065407b, 32'h439f1c82},
  {32'h439dc380, 32'hc26e6830, 32'hc2ca733e},
  {32'h439c4450, 32'hc3c1f493, 32'h4385112d},
  {32'h4411c24f, 32'hc3383d5e, 32'hc318f933},
  {32'hc488370d, 32'h4388bf31, 32'h43f6c7a2},
  {32'h440b0a80, 32'hc2bd6a29, 32'hc2d1a0ab},
  {32'hc47ed1bd, 32'h43a04768, 32'h43793c5f},
  {32'h44263546, 32'hc2fb84d9, 32'h43771dad},
  {32'hc4f5b116, 32'hc3177d30, 32'h4322eaea},
  {32'h43c81df0, 32'hc38dfb67, 32'hc2b58af3},
  {32'hc4a5136a, 32'hc238f5c2, 32'h429bcbf9},
  {32'h44f098f4, 32'hc43860a0, 32'h437f9ff0},
  {32'hc454facb, 32'hc3ff6848, 32'hc2f84767},
  {32'h450bc017, 32'h430bf8f2, 32'hc27764ea},
  {32'hc4bab830, 32'hc28c3f7a, 32'hc22bb5ac},
  {32'h437373a8, 32'hc01cea56, 32'h43432d53},
  {32'hc4ae863d, 32'h42c3de11, 32'h43086556},
  {32'h44f0931a, 32'h4386ce49, 32'hc37805e2},
  {32'hc436b9f0, 32'hc316fb63, 32'hc21b80da},
  {32'h44afd10a, 32'hc42a1dd1, 32'h42d78bd3},
  {32'h416f9500, 32'hc324a81d, 32'hc2f33d29},
  {32'h44d1228e, 32'h4339a002, 32'hc24e9121},
  {32'hc4b48db0, 32'hc2f9fc3f, 32'hc3032fec},
  {32'h450e21ae, 32'h43a30183, 32'hc33190e6},
  {32'hc4165310, 32'hc2944e96, 32'h42be7440},
  {32'h44bba66d, 32'hc2aa4e53, 32'h4395c5fd},
  {32'hc4c4bc9c, 32'hc38ff644, 32'hc38be05d},
  {32'h44e9cfad, 32'hc22ef227, 32'hc302ba3e},
  {32'hc36f32b4, 32'hc411d536, 32'hc3a70d9b},
  {32'h44ec992d, 32'hc2223764, 32'hc3be4b48},
  {32'hc49bbbb9, 32'h4384f777, 32'h438ca36b},
  {32'h450a5d4f, 32'h43213d3d, 32'h4322850d},
  {32'hc4bb1f76, 32'hc1fb2120, 32'h4214809c},
  {32'h44b5b1e0, 32'h429e056b, 32'hc3aaf819},
  {32'hc3c81312, 32'h42926236, 32'h413c8f44},
  {32'h44f13a84, 32'hc2009a72, 32'hc3a6cbd3},
  {32'hc402705b, 32'h438844c1, 32'hc2d9fbab},
  {32'hc2f09ea0, 32'hc2887a7c, 32'h435dc31f},
  {32'hc4a99191, 32'hc2d56b44, 32'h425a5c68},
  {32'h451beba5, 32'hc3302613, 32'h438f8885},
  {32'hc4502662, 32'h41bb6854, 32'h4324b804},
  {32'h43a5973c, 32'h43066bff, 32'hc30c482f},
  {32'hc4da3661, 32'h42a0a857, 32'hc2f71807},
  {32'h44ab17f4, 32'hc327f0ae, 32'hc300bd5b},
  {32'hc4ccab7d, 32'hc31b06cd, 32'hc2d584b8},
  {32'h43313f90, 32'hc39a1e7e, 32'hc0023ffc},
  {32'hc31ce4b8, 32'h4391a099, 32'h438c6c59},
  {32'h44aed4c2, 32'hc14bc1f0, 32'hc2f02459},
  {32'hc42cd6c3, 32'h433e8cce, 32'hc1edf1c6},
  {32'h450c1169, 32'h42a4dffa, 32'h43a6d256},
  {32'hc48bc6ef, 32'hc1a0f540, 32'hc1c82d1c},
  {32'h451fcde8, 32'hc3eb9dbe, 32'h43e33959},
  {32'hc3922da0, 32'h43cd1e5e, 32'hc387b744},
  {32'h4406cd3e, 32'hc3b4db74, 32'h4320ce10},
  {32'hc3aac798, 32'h43cdeefe, 32'h43302085},
  {32'h4380c8b1, 32'h43c329d2, 32'h43af7ad4},
  {32'hc2f6135e, 32'h40a4f9c0, 32'hc361524e},
  {32'h44d01411, 32'h44018ac3, 32'hc18a5156},
  {32'hc43ec578, 32'h4390ca56, 32'h4334d122},
  {32'h43f08638, 32'h42d9b6b6, 32'hc1b7e59e},
  {32'hc507a140, 32'h41e79572, 32'hc3b59605},
  {32'h44773dd2, 32'hc365272c, 32'h418fe726},
  {32'hc506a908, 32'hc344b8fe, 32'h42d4fa81},
  {32'h444f2bba, 32'hc39902f6, 32'hc332b4a1},
  {32'hc4029802, 32'h4239ad4f, 32'h41d9c7c0},
  {32'h4410e75c, 32'h438375e8, 32'hc21a4ddc},
  {32'hc48582d2, 32'hc37928be, 32'hc2e2e3f3},
  {32'h450e42e2, 32'h41450200, 32'h43bd1ec5},
  {32'hc4877bff, 32'hc2bddc23, 32'hc2cda728},
  {32'h44e97c3c, 32'hc1c8286c, 32'h42b73f78},
  {32'hc48d5f6e, 32'h43630a24, 32'hc39d282d},
  {32'h443598b8, 32'h42e13650, 32'hc299534b},
  {32'hc4bf271c, 32'hc233cdbb, 32'hc2c65cdc},
  {32'h44cdb4d6, 32'h4383592e, 32'hc30095b5},
  {32'hc4a55e6a, 32'h43aaf9dd, 32'h43c21f21},
  {32'h44bb3793, 32'hc11ea728, 32'h42c4efc9},
  {32'hc4d4995c, 32'h4336cf6d, 32'hc3431ee4},
  {32'h44d24100, 32'hc396029e, 32'hc29ed185},
  {32'hc41f8b6c, 32'h43a9deb9, 32'hc35f3c5b},
  {32'h44ecc161, 32'hc3002c75, 32'hc2270648},
  {32'hc39b968d, 32'hc2a4411c, 32'h4288dd67},
  {32'h44855fce, 32'hc3728c5d, 32'h4387558a},
  {32'hc50a9d35, 32'h43124824, 32'h430592c2},
  {32'h43f28845, 32'h437248a2, 32'h42f9f0a3},
  {32'h41ea7700, 32'h431a07d1, 32'hc33c5bd5},
  {32'h445a36e2, 32'h43cf4591, 32'hc22bfa24},
  {32'hc3b409f8, 32'hc282d779, 32'hc334d3de},
  {32'h44b782da, 32'hc2b4747c, 32'hc31aff61},
  {32'hc4aa2687, 32'h438ce408, 32'hc2a2a86e},
  {32'h451af63e, 32'hc282a8ac, 32'h429f9460},
  {32'h424bddfe, 32'h42887775, 32'h4316cddc},
  {32'h44388e23, 32'h42c3b484, 32'hc3e255f0},
  {32'hc4b1c6ec, 32'hc2ce1ac1, 32'hc331c7d7},
  {32'h44c65f4f, 32'h43fa2353, 32'hc30f1f65},
  {32'hc37b29e8, 32'hc2b25c55, 32'h427b4687},
  {32'h44f99d3e, 32'h417fa0e3, 32'hc24f9e79},
  {32'hc2bd2714, 32'h432ca1f5, 32'hc3e9925f},
  {32'h4500a128, 32'h4388c7f4, 32'hc3e3e0cc},
  {32'hc4950fa2, 32'hc313d4a8, 32'hc38bd73b},
  {32'h44dcf23a, 32'h42bf98e2, 32'h4363eacf},
  {32'hc482ea54, 32'hc2c25ab4, 32'h433fcb63},
  {32'h44590a82, 32'h42210ff7, 32'hc3247327},
  {32'hc4412ecc, 32'h41f8cc52, 32'hc370bbc2},
  {32'h45094361, 32'h4181d030, 32'h421bde95},
  {32'hc5110c9f, 32'h4180890c, 32'h4393f718},
  {32'h450e5e7e, 32'hc2df6fdb, 32'hc2f0e4ad},
  {32'hc4561f9d, 32'h42541afb, 32'hc333e99d},
  {32'h44c8aa8c, 32'h42e7b3ed, 32'hc2eaadb2},
  {32'hc4467284, 32'h439eba4f, 32'hc2a0eb95},
  {32'h44220a0b, 32'hc342b321, 32'h42a875f3},
  {32'hc5031c40, 32'hc3b2a976, 32'hc2fe090f},
  {32'h44053b52, 32'hc35b8d84, 32'hc2405375},
  {32'hc48b5156, 32'h43333f89, 32'hc33d054a},
  {32'h44b61f46, 32'h4306c87c, 32'hc2de046e},
  {32'hc3a41788, 32'h433e9c4a, 32'h430407bc},
  {32'h446a38aa, 32'h422efbdd, 32'h4346f56c},
  {32'hc3c001a8, 32'h42177352, 32'hc3911f2d},
  {32'h44700920, 32'h4166acbc, 32'hc208a16d},
  {32'hc46b0867, 32'h43143897, 32'hc2b516e0},
  {32'h434e4110, 32'hc38a5ff2, 32'hc2827078},
  {32'hc312a3ec, 32'h43c3db86, 32'h431d7f0e},
  {32'hc23261f0, 32'hc32853d5, 32'hc2bb3b93},
  {32'hc4e634bc, 32'hc20c79e1, 32'h42f9a52f},
  {32'h45140c76, 32'hc367767f, 32'h427739b8},
  {32'hc4ef1f78, 32'hc35bceef, 32'h432c7a2f},
  {32'h4420bb8c, 32'h4257ba90, 32'h43700ead},
  {32'hc3b9d919, 32'h42f26451, 32'h420a982b},
  {32'h44d28388, 32'h42e82a14, 32'hc32daa97},
  {32'hc396e198, 32'h433d3251, 32'hc34557f0},
  {32'h4514654c, 32'h43229030, 32'hc29b23e6},
  {32'hc4c5e419, 32'hc2d7fd3a, 32'hc2c06724},
  {32'h442a56e8, 32'hc20d55be, 32'hc2f83a5c},
  {32'hc5105237, 32'hc2cbea39, 32'h43406008},
  {32'h451b91c6, 32'h43803a1a, 32'hc225df46},
  {32'hc48aa40e, 32'hc3481039, 32'h438f01ba},
  {32'h4535f60b, 32'h419182a4, 32'h41afae14},
  {32'hc505f0fb, 32'hc36bcddf, 32'hc22f0ca2},
  {32'h446eecae, 32'hc38f492d, 32'h43189ca4},
  {32'hc4d7c160, 32'hc28670b2, 32'h41c0adae},
  {32'h44df67c0, 32'hc33de4ea, 32'h4388c2e3},
  {32'hc4862966, 32'hc2081f6e, 32'h43810871},
  {32'h44b144e4, 32'hc36d62ed, 32'hc3b5c1b9},
  {32'hc4cecc9d, 32'h433b4722, 32'hc245d871},
  {32'h44b0acc8, 32'h43096a12, 32'hc2cf539b},
  {32'hc2bf4100, 32'hc38f4ee4, 32'hc2489223},
  {32'h43c69174, 32'hc324a199, 32'h41623425},
  {32'hc49032f5, 32'hc35836fc, 32'h43498566},
  {32'h45008356, 32'hc31cdfef, 32'hc32140de},
  {32'hc4e566e7, 32'h436ca803, 32'hc1e566d0},
  {32'h44a423ab, 32'h42ada60c, 32'hc37db942},
  {32'hc4a5b4fd, 32'h42c2a8e6, 32'h42146cb8},
  {32'h45186faf, 32'hc2d2f9da, 32'h432df04a},
  {32'hc4b50307, 32'h43b9429a, 32'hc3b3a5e6},
  {32'h4493c647, 32'hc30eb1b0, 32'h43877f4f},
  {32'hc4b05f04, 32'h440f716e, 32'h42eaff6d},
  {32'h44aea7ee, 32'h437a9c81, 32'hc34783a6},
  {32'hc49e127b, 32'h409dd37d, 32'h433b2fb2},
  {32'h4506beca, 32'h438b2acd, 32'hc3f3c096},
  {32'hc4829142, 32'hc1fbf8e8, 32'hc33dc47e},
  {32'h44884e62, 32'hc325da73, 32'hc35b1332},
  {32'hc50e2c9a, 32'hc205bffc, 32'h43700a14},
  {32'h440716de, 32'hc30c963d, 32'hc3ebae4e},
  {32'hc3c27990, 32'h43202daf, 32'h42266e1c},
  {32'h44911150, 32'hc2bbac9e, 32'hc300407f},
  {32'hc45a07d0, 32'h42b92c53, 32'h43765dd6},
  {32'h43e41914, 32'hc1ae0b7e, 32'hc1a10502},
  {32'hc5062961, 32'h42ab4a22, 32'hc397b88b},
  {32'h45065e9f, 32'h4216efbf, 32'h426f220f},
  {32'hc4518105, 32'h43ad7f0f, 32'hc24ecfa8},
  {32'h44ef6db8, 32'hc3981d3f, 32'hc20130f6},
  {32'hc4e79a4a, 32'hc2c86b74, 32'h438c93d4},
  {32'h4457f078, 32'hc379c45b, 32'h439a02a5},
  {32'hc4a49679, 32'hc1911960, 32'hc21860e0},
  {32'h44492450, 32'h4383c4d0, 32'h42aaf50c},
  {32'hc4ee46b9, 32'hc0cfc4f8, 32'h4363e238},
  {32'h449a8ebe, 32'hc1f560a1, 32'h4281f1e2},
  {32'hc508a3b9, 32'h429798eb, 32'hc27db4d2},
  {32'h450a12b8, 32'h42c6ae6c, 32'h438f83d1},
  {32'hc5045c2d, 32'hc3ad6f0e, 32'h429e9454},
  {32'h42d8d768, 32'hc38b735a, 32'hc30592fc},
  {32'hc404acac, 32'h42992ba5, 32'h4300596b},
  {32'h4518144f, 32'hc2a17c0f, 32'h426fd446},
  {32'hc4e3e8f7, 32'hc270704e, 32'hc34516dd},
  {32'h448bf70c, 32'hc336bdc1, 32'h42a5a1e6},
  {32'hc49d009f, 32'h437fb6c9, 32'h434c44a2},
  {32'hc1e1aa80, 32'hc3e7fd25, 32'hc33a0ee1},
  {32'hc3d42376, 32'h43b2681c, 32'hc32eb3cb},
  {32'h444c4e89, 32'hc21b8d89, 32'h42df2edc},
  {32'hc4b860b5, 32'h4342add3, 32'hc407bf19},
  {32'h4459202e, 32'hc224cc82, 32'h3f426207},
  {32'hc4867076, 32'h4326d1af, 32'hc266f776},
  {32'h45039b0a, 32'h43212ad8, 32'h42df38e0},
  {32'hc503d235, 32'h43638c10, 32'hc367fa4a},
  {32'h43c4133a, 32'hc1c31046, 32'h42b7188c},
  {32'hc5008382, 32'h42ea8c8f, 32'hc2832e4d},
  {32'h4514c7b8, 32'hc3837ac7, 32'h432193c3},
  {32'hc50326c5, 32'hc3991e89, 32'hc15fc545},
  {32'h42186b40, 32'h434c52dc, 32'h43428570},
  {32'hc470dd10, 32'h43c7b0d7, 32'h41c47f4f},
  {32'h44ff31f6, 32'hc39fb373, 32'hbf32ab40},
  {32'hc495216d, 32'hc1e22d80, 32'h4283d5b8},
  {32'h44cc9dc4, 32'h43203a3f, 32'hc2113e71},
  {32'hc47b8701, 32'hc19d7368, 32'hc399d9f2},
  {32'hc297ffe0, 32'hc3ba1871, 32'h4401cffd},
  {32'hc4b2b697, 32'h422b12bb, 32'hc2b821f4},
  {32'h421ba62f, 32'hc3ea0566, 32'h41e26243},
  {32'hc50414ef, 32'h4334779f, 32'hc39a31dc},
  {32'h43ac9a5e, 32'h42400e32, 32'hc2a13faf},
  {32'hc4b4f54a, 32'h42dc32c1, 32'hc252f98c},
  {32'h43423b20, 32'hc34c8169, 32'hc2e31674},
  {32'hc4b47eca, 32'h4300b873, 32'h4200686e},
  {32'h43933796, 32'hc1745363, 32'h42ff688d},
  {32'hc42794d8, 32'h40922176, 32'hc0989bdb},
  {32'h43344370, 32'h43030105, 32'h430b0467},
  {32'hc3a401c3, 32'h42502f1e, 32'hc3292fdd},
  {32'h4373dd80, 32'hc35de133, 32'h421b2b3f},
  {32'hc4d87ecc, 32'h43148cc9, 32'hc3c9185f},
  {32'h4489a0c2, 32'hc402e5b2, 32'h43b9589d},
  {32'hc40761f1, 32'hc33198b7, 32'hc2a72e01},
  {32'hc4fcf0ac, 32'h4301a91a, 32'h42bc292c},
  {32'h43a6a0d2, 32'hc37cd77c, 32'h430fbd00},
  {32'h432f3dac, 32'h44008310, 32'hc32a2065},
  {32'h44ac8deb, 32'hc2cb6589, 32'hc1e506bf},
  {32'hc4d75c3e, 32'hc31b21be, 32'hc2b76332},
  {32'h4311b43c, 32'hc3186e0b, 32'h43b42528},
  {32'hc4c52847, 32'hc3243bc0, 32'hc39c36a3},
  {32'h43ab3330, 32'h436c1644, 32'hc38209df},
  {32'hc4eaff0e, 32'hc2e58737, 32'hc24a8342},
  {32'h441cb14f, 32'h435113e7, 32'h43a492f4},
  {32'hc40a7774, 32'h4347b6e4, 32'h420da30e},
  {32'h4476d5b2, 32'h42ef96b6, 32'h43210aee},
  {32'hc46fe2f0, 32'hc37174f3, 32'hc3884e72},
  {32'h4407c175, 32'hc28ab3a7, 32'hc31e2615},
  {32'h429bfa05, 32'h43c9dbe6, 32'h416d98da},
  {32'h43c95c50, 32'hc397ec16, 32'hc42c7a8e},
  {32'hc488aafa, 32'h42bdd81c, 32'h4223d1ce},
  {32'h45052c3e, 32'hc369feb7, 32'hc049db13},
  {32'hc4a973bf, 32'h42b7df01, 32'hc22c0ec7},
  {32'h4507cf0a, 32'hc28cb8d0, 32'h42bd9154},
  {32'hc419a8c4, 32'h4327a8c3, 32'hc23aee39},
  {32'h44855046, 32'hc381c508, 32'h42bc0d5e},
  {32'hc4f8fee8, 32'hc394f448, 32'h43217106},
  {32'h449add14, 32'h43a21ba5, 32'h4376066b},
  {32'hc5041799, 32'hc2ac2c1b, 32'hc3af6576},
  {32'h432e6ad1, 32'h436531d2, 32'h4384117f},
  {32'hc4f2245f, 32'h423e067a, 32'h430b1163},
  {32'h44e25019, 32'hc3ac1cd7, 32'hc33b1726},
  {32'hc50db495, 32'hc29dfbdb, 32'hc378afdb},
  {32'h4505b22d, 32'h43155975, 32'hc394c2b5},
  {32'hc3740504, 32'hc2c5fa0c, 32'hc255d008},
  {32'h44054c52, 32'h437d5bd4, 32'h434086e6},
  {32'hc4cadbed, 32'hc3be3300, 32'hc3b6c4cb},
  {32'h44ccbd76, 32'hc367f334, 32'h42ac2740},
  {32'hc4fc49db, 32'h43d5b2cb, 32'h43292027},
  {32'h44cbf714, 32'hc2e85254, 32'h40cb5790},
  {32'hc4719210, 32'hc2169782, 32'hbfc94850},
  {32'h4391852e, 32'hc2600348, 32'hc307f378},
  {32'hc49457cf, 32'h40f45f53, 32'h437514c6},
  {32'h441896c6, 32'hc240f52d, 32'hc2b04f4f},
  {32'hc428f9d0, 32'h43257107, 32'hc23b760f},
  {32'h43ad8f4c, 32'h3f349069, 32'h438335fb},
  {32'h42a3421e, 32'hc3eb733e, 32'h43a8daca},
  {32'h43480030, 32'h42f1d6f0, 32'h433fee17},
  {32'hc481fa5d, 32'hc40851ca, 32'h41fef594},
  {32'h43c08218, 32'hc30bc508, 32'hc2dd827f},
  {32'hc4ebf1fc, 32'hc307ef67, 32'hc29e850e},
  {32'h443cb7c8, 32'hc33480ac, 32'hc385c6ec},
  {32'hc4f0c7b6, 32'hc39ed06b, 32'hc26d14ba},
  {32'h444223d6, 32'hc3a3b1bf, 32'hc2070262},
  {32'hc447e5b8, 32'hc28ad626, 32'hc2950678},
  {32'h44a895d1, 32'h440b6ed8, 32'h433cfe24},
  {32'hc4c3e430, 32'h43068a89, 32'hc23f8f92},
  {32'h44ed7a67, 32'h43a4d1ff, 32'hc37502b6},
  {32'hc444760c, 32'h428d7147, 32'hc29a9f24},
  {32'h43d8eed5, 32'hc3bb8337, 32'hc37cb975},
  {32'hc3e028f3, 32'hc2f8baff, 32'h42f9f007},
  {32'h4452efc4, 32'h42f8e8b4, 32'hc2fea071},
  {32'hc1094000, 32'h4228f208, 32'hc3ad2eb2},
  {32'h444c4e52, 32'hc29da485, 32'hc31019f8},
  {32'hc4fd4fec, 32'h431e7f53, 32'h41c425ac},
  {32'h446a2a9a, 32'hc3d0f356, 32'h437cd6fb},
  {32'hc4e21642, 32'hc26d859e, 32'h43216ed9},
  {32'h45148fb3, 32'hc3f8d910, 32'hc0c11a4c},
  {32'hc4360622, 32'h439b3e07, 32'h439a95b5},
  {32'h450641fc, 32'h438f77c5, 32'h4332549d},
  {32'hc5139238, 32'h43257f6b, 32'hc2b41559},
  {32'h443f4cdf, 32'h42cb96dc, 32'hc3224bc5},
  {32'hc493705e, 32'h41f22f38, 32'h4363b376},
  {32'h44a7f505, 32'hc328cee6, 32'h42a4a404},
  {32'hc50768f3, 32'h43ac00af, 32'hbfa724f4},
  {32'h440bf8ff, 32'hc38a84a2, 32'hc32f911f},
  {32'hc49a6c09, 32'hc360278e, 32'h43692e9a},
  {32'h44bc7b6d, 32'h4353e8d1, 32'h4269a59c},
  {32'hc4f0a2ad, 32'hc2e98edd, 32'hc4070411},
  {32'h44e703a6, 32'hc3281ddf, 32'h42686626},
  {32'hc48fda5b, 32'h41fe731a, 32'hc3298e9e},
  {32'h446915bd, 32'h4207f8fc, 32'hc39f37ae},
  {32'hc4c43e25, 32'hc3242619, 32'hc29f5c33},
  {32'h43c06874, 32'hc43e1bce, 32'h43412d13},
  {32'hc506ce2c, 32'h43345f78, 32'hc34be3cc},
  {32'h450a38b3, 32'hc3a9d00a, 32'hc29b1f4d},
  {32'hc4818983, 32'hc3191795, 32'hc3cb24c6},
  {32'h44493a80, 32'h43965f4a, 32'hc3dc328f},
  {32'hc3bc0c44, 32'h43e9e5c0, 32'h43783b88},
  {32'h4500e3fc, 32'hc38c4029, 32'h433a85ee},
  {32'hc4cead50, 32'h41fdc5fb, 32'hc1badaa1},
  {32'h44b4a50c, 32'h43f9a4bc, 32'hc3345048},
  {32'hc4e5eb5a, 32'hc33993c8, 32'h4224d6df},
  {32'h44915a2d, 32'hc3256daf, 32'hc26b1635},
  {32'hc4a3519b, 32'h418ac125, 32'hc3b03f6e},
  {32'h44f2c02e, 32'h41ff4c77, 32'hc312ede6},
  {32'hc419a484, 32'h41bc8e13, 32'hc35ac366},
  {32'h43000330, 32'hc1eb1d7f, 32'h43a7270e},
  {32'hc48c042a, 32'hc3d21c8f, 32'hc3a0f220},
  {32'h445cbdd0, 32'hc327da05, 32'h41247f38},
  {32'hc502146f, 32'hc2d13631, 32'hc3088b6d},
  {32'h44fd80fb, 32'h4386fa6b, 32'hc328cef6},
  {32'hc304246c, 32'hc308b148, 32'h431459bd},
  {32'h440cc84e, 32'hc2a03f3c, 32'hc3629fdd},
  {32'hc47c6d36, 32'h4250c0fb, 32'h42ec1cb8},
  {32'h43ada20c, 32'h43031b8a, 32'hc368145d},
  {32'hc502d2c3, 32'hc3061c55, 32'h4328f4c0},
  {32'h442079ea, 32'hc1c98724, 32'hc20f3ceb},
  {32'hc440dfcc, 32'h439d8abd, 32'hc21bbe79},
  {32'hc2970474, 32'h43235aa9, 32'hc3074f19},
  {32'hc3ccb46b, 32'h43e091c0, 32'hc2e16cbf},
  {32'h43de51a0, 32'hc3420f03, 32'hc2f14423},
  {32'hc1be7a17, 32'h4336cc60, 32'hc34989b4},
  {32'h451aaf7b, 32'h418a378d, 32'hc38354cb},
  {32'hc48ce587, 32'hc2e9a235, 32'h435f0558},
  {32'h44aa83c6, 32'h43884479, 32'h439d3247},
  {32'hc4ecdffc, 32'h42c52087, 32'h43234d47},
  {32'h44b488a3, 32'h43231cc2, 32'h42dd25d9},
  {32'hc499f06e, 32'h439f9927, 32'hc3034fb4},
  {32'h4456f44e, 32'hc25981f6, 32'hc38e539a},
  {32'hc4bbfbe8, 32'hc24835c8, 32'h439158e1},
  {32'h445c6b37, 32'h434e72ed, 32'h434a3467},
  {32'hc4e7a000, 32'h43d582f3, 32'h4288cbf6},
  {32'h449ce2c8, 32'hc3576e3a, 32'h426c10cb},
  {32'hc4f639c6, 32'h43e42023, 32'hc20c086b},
  {32'h44ca2241, 32'hc2121490, 32'h427b9152},
  {32'hc422b42b, 32'hc3989431, 32'h42a08bba},
  {32'h44f9fee6, 32'h4389072a, 32'h434185c9},
  {32'hc3a1fc8c, 32'h42569723, 32'hc3d29661},
  {32'h4481e2d4, 32'hc287ab3b, 32'hc2fb362b},
  {32'hc4a638c6, 32'h43310518, 32'h43ab1121},
  {32'h43dc4667, 32'h42af5d8f, 32'h43880737},
  {32'hc2900040, 32'h42246084, 32'h43c912ef},
  {32'h44cf3c32, 32'h435e0060, 32'hc382ccfc},
  {32'hc4b05d10, 32'h43e78eaa, 32'h436cb8b6},
  {32'h450bf5dd, 32'hc3e1ab39, 32'h440974a3},
  {32'hc4fcaffb, 32'h42e3fc11, 32'h42fbab6d},
  {32'h44b6e900, 32'h42e6fde4, 32'hc2b986d6},
  {32'hc4e3dc67, 32'hc3ac339a, 32'h43a047a0},
  {32'h451372a8, 32'h42b57e25, 32'hc35298f0},
  {32'hc4f5d41c, 32'hc3440eb0, 32'hc29508b2},
  {32'h44dd71e6, 32'h43c344bc, 32'hc3da4557},
  {32'hc4be0b97, 32'h4323c96b, 32'h431df34f},
  {32'h44635dd8, 32'hc38463ea, 32'hc11f292b},
  {32'hc46600af, 32'hc1f2089e, 32'hc2646396},
  {32'h44fa375a, 32'hc35b8424, 32'hc38cae1d},
  {32'hc4c75d0c, 32'h430467dd, 32'h4361c30c},
  {32'h43f84f30, 32'hc393e8c0, 32'hc28492ca},
  {32'hc4f99c4a, 32'h42a8c9dc, 32'hc34f3251},
  {32'h448856ee, 32'h42b5b6e9, 32'h43410d7e},
  {32'hc48aea0b, 32'h42d33923, 32'h4357a101},
  {32'hc004bdc0, 32'h432b52fe, 32'hc34be9d7},
  {32'hc487f2f4, 32'hc4396ba3, 32'h440293bb},
  {32'h4458235a, 32'hc2d73fd1, 32'h438298eb},
  {32'hc4bd3a64, 32'h42a43c7c, 32'hc3466cd3},
  {32'h44b948d7, 32'h42f532d1, 32'h4351a5b4},
  {32'hc4a6f81c, 32'hc34606ef, 32'hc37a025c},
  {32'h444cd6f2, 32'h433fe569, 32'h43f313d3},
  {32'h4165ec00, 32'h426a6b30, 32'hc204256b},
  {32'h44e73531, 32'h4395e287, 32'hc31aa949},
  {32'hc49c9630, 32'hc3266d22, 32'hc2b4bbad},
  {32'h43932b8d, 32'hc28cc5d1, 32'hc2fc50fd},
  {32'h3fa70b40, 32'h4016dcf7, 32'hc3225930},
  {32'h440547d1, 32'h42929895, 32'h42540cfa},
  {32'hc40a7f37, 32'hc35d2059, 32'hc22d4e48},
  {32'h442c81a8, 32'h439df5d1, 32'h43215a89},
  {32'hc47540f0, 32'hc2e39254, 32'h41a0d7e9},
  {32'h43f6e732, 32'h4356dd87, 32'hc337e900},
  {32'hc4350f34, 32'hc364d3ab, 32'h3f3b0768},
  {32'h441bf68f, 32'hc38f90cd, 32'h428da6c9},
  {32'hc4af9f55, 32'h430c1461, 32'hc40113b5},
  {32'h44d79b38, 32'h43952177, 32'hc38f8d87},
  {32'hc1d9ffa0, 32'hc3e9c182, 32'h42c029a9},
  {32'h43a92650, 32'hc4007cda, 32'h4399950b},
  {32'hc4f9b45a, 32'hc383fe85, 32'h438d2ada},
  {32'h448b8f60, 32'h43ea9463, 32'h43699580},
  {32'h41cf73c0, 32'hc364f4c3, 32'hc407cfff},
  {32'h4481c4f7, 32'h431fa247, 32'hc361706f},
  {32'hc5022299, 32'hc398be61, 32'h402fbf72},
  {32'h450d11fa, 32'hc1b0596d, 32'h429b429e},
  {32'hc3f2e22f, 32'h427f3814, 32'h4263bf33},
  {32'h43b9d1e8, 32'hc38e0bfa, 32'h42b4491b},
  {32'hc3b22da6, 32'hc3885ee3, 32'h43306b1f},
  {32'h4305c30e, 32'h4288c9c3, 32'h422ae108},
  {32'hc4539594, 32'h434d2846, 32'h4041d4ac},
  {32'h447c5130, 32'h430be859, 32'hc3c420a4},
  {32'hc48f3160, 32'hc30553f3, 32'hc30fe521},
  {32'h43616ed0, 32'h42b07f12, 32'hc3256fa5},
  {32'hc436d276, 32'hc20c898d, 32'hc1cf3dc9},
  {32'h442825aa, 32'hbf1ac4ec, 32'h43ebdd96},
  {32'hc4d76a34, 32'h437166dd, 32'h428556ab},
  {32'h44cfa84c, 32'hc29617a7, 32'h40b1c927},
  {32'hc50ae2b2, 32'hc3b0c1b1, 32'h42151117},
  {32'h45190d54, 32'h42e10eeb, 32'h41ea9161},
  {32'hc4b79b1e, 32'h438f192e, 32'hc2f7ce80},
  {32'h45009bbd, 32'hc333a786, 32'hc1893343},
  {32'hc4fd8098, 32'hc2770cca, 32'h42e33af0},
  {32'h43326912, 32'h433b1b47, 32'h42d20449},
  {32'hc4f4d7de, 32'h425c7ea3, 32'hc2bc213a},
  {32'h44218ba5, 32'hc3d934ca, 32'hc20cf6e6},
  {32'hc4e4298b, 32'h43a974d7, 32'h42875d22},
  {32'h448d7b9d, 32'hc3106e9e, 32'h4242e344},
  {32'hc390206d, 32'h4267f598, 32'h412512a3},
  {32'h448d90c8, 32'hc2999386, 32'h41e289e8},
  {32'hc4f59ca6, 32'hc3d014a7, 32'hc324fc94},
  {32'h44710acc, 32'h42bccdab, 32'hc28f6361},
  {32'hc48079d1, 32'h4369db30, 32'hc3bf043a},
  {32'h44370798, 32'h41deeafe, 32'hc3226752},
  {32'hc50ebfdf, 32'h4388c7e4, 32'hc208563d},
  {32'h4493471c, 32'hc2c4d5c3, 32'hc2a47036},
  {32'hc4f5e031, 32'hc369fb86, 32'h433ad9d4},
  {32'h43fb7078, 32'hc1a96c44, 32'hc223a29a},
  {32'hc4d7bdea, 32'hc2d19511, 32'hc4329a8a},
  {32'h447a1e31, 32'h43e40610, 32'h43257ffd},
  {32'h43279f86, 32'h416cc251, 32'h43832a37},
  {32'h439e84c2, 32'hc34e3dba, 32'hc06e2c90},
  {32'hc4e2fdf3, 32'h42e5990f, 32'h4338f63f},
  {32'hc2b69fb0, 32'h414ae0c0, 32'h4305c9e7},
  {32'hc315eaa2, 32'h438c4539, 32'h4403ab58},
  {32'h44e88b98, 32'hc29771f2, 32'hc3b96795},
  {32'hc493a0bb, 32'h4387080a, 32'hc3b090bf},
  {32'h432e7b98, 32'h42122202, 32'h42880f15},
  {32'hc4745917, 32'hc350e6cb, 32'h417e4cb8},
  {32'h44f42754, 32'hc3435f01, 32'hc39f034d},
  {32'hc501de32, 32'hc35f4b33, 32'hc0f7671d},
  {32'h44edcbd6, 32'hc32bd0fd, 32'h42d7a0ba},
  {32'hc4b06162, 32'h43be4f36, 32'h429bec05},
  {32'h44e4af1b, 32'hc236f8db, 32'hc3b1bb21},
  {32'hc4280e8b, 32'hc3386cd1, 32'hc2397c18},
  {32'h4451991a, 32'h4305bc3f, 32'hc3e28772},
  {32'hc4d2596a, 32'h424163dc, 32'h43a54c15},
  {32'h43c1fcbc, 32'h420077ac, 32'h43190e18},
  {32'hc503bec2, 32'hc3abe94f, 32'h42cd395f},
  {32'h44c832a3, 32'hc2f979e0, 32'hc353104d},
  {32'hc4a0d33a, 32'h439bd7b4, 32'h43598ac8},
  {32'h443f8fc8, 32'h428a8dc6, 32'h439e831a},
  {32'hc4305c97, 32'h437395e3, 32'hc33383aa},
  {32'h44d6969c, 32'hc3036290, 32'hc27d7ee8},
  {32'h431a2cd6, 32'hc30dbd2b, 32'hc3581226},
  {32'h443f4fa3, 32'h42dae3a6, 32'h4239bae2},
  {32'hc4843bc4, 32'hc39906cf, 32'hc0e59fa8},
  {32'h4483bcd6, 32'hc24018ee, 32'h432b651c},
  {32'hc51570df, 32'hc405f762, 32'hc2cae3b5},
  {32'h43fc5efc, 32'hc28b97ba, 32'hc2e2271a},
  {32'hc3e49a66, 32'hc227f6e2, 32'h43ec524f},
  {32'h44f87144, 32'h4362950f, 32'h43120bb4},
  {32'hc502a424, 32'hc3134cb2, 32'h43e3f1af},
  {32'h44591988, 32'hc3475be2, 32'hc217bb54},
  {32'hc47a646d, 32'h42fb8731, 32'hc1196dbb},
  {32'h44d90597, 32'hc33a322c, 32'h43c7564e},
  {32'h42030450, 32'h4287dfe7, 32'hc3d7caac},
  {32'h445067cc, 32'hc386f287, 32'h437efcf1},
  {32'hc480fe3b, 32'h42a08e9c, 32'hc389cd72},
  {32'h44d649d5, 32'hc358ba98, 32'h4335e91c},
  {32'hc4e090db, 32'h429ae273, 32'hc3115afc},
  {32'h44c78eb1, 32'hc35ca8d6, 32'h423370c9},
  {32'h432a92a0, 32'hc2b56886, 32'hc3588a79},
  {32'h4433f05c, 32'hc3ba8007, 32'hc36b6fc1},
  {32'hc4d58085, 32'hc343d1e2, 32'h42e3cb5f},
  {32'h449ac8d2, 32'hc3fcf3a6, 32'h43a1401d},
  {32'hc4f1d5bc, 32'h429052ba, 32'hc3535428},
  {32'h43956a84, 32'hc2bf0116, 32'h429d28b8},
  {32'hc4ce5224, 32'h42b81f40, 32'hc3412438},
  {32'h443d6f6e, 32'hc2a2fcd3, 32'hc234ab49},
  {32'hc4866fc5, 32'h430310c9, 32'h4266f09b},
  {32'h44df8b04, 32'hc26ee2d7, 32'h430618d7},
  {32'hc454eb44, 32'h442bac64, 32'h437dfe5f},
  {32'h441a95cf, 32'h42ec7bc7, 32'hc3d63bf1},
  {32'hc42cca9c, 32'h41212c38, 32'hc233d9c4},
  {32'h4303d63c, 32'h437ef194, 32'hc31cb833},
  {32'hc502fc47, 32'h424e3116, 32'h430273c2},
  {32'h4423957d, 32'h43bba364, 32'h434a61fb},
  {32'hc286c260, 32'h430b1321, 32'h4198c97b},
  {32'h43f13930, 32'h419ddc46, 32'h4354f80d},
  {32'hc3a596ef, 32'hc16984c7, 32'h421e8d5c},
  {32'h43ad0020, 32'hc38cdb24, 32'hc30ff2ae},
  {32'hc4c363da, 32'h4370253b, 32'hc2ea848a},
  {32'h44dee0ec, 32'h4392050a, 32'hc2fc9576},
  {32'hc4e79259, 32'hc3919248, 32'hc2b13317},
  {32'h44775298, 32'hc41365bf, 32'hc3764fb2},
  {32'hc415ea3c, 32'hc252c28c, 32'hc2e780f6},
  {32'h451939c8, 32'hc2d10c78, 32'h40befc2a},
  {32'hc5141fbb, 32'hc0df9ad4, 32'hc39a1b20},
  {32'h44090a82, 32'hc36d9b98, 32'h43966acd},
  {32'hc498d3af, 32'hc207621a, 32'hc2e43367},
  {32'h44ff742d, 32'h42e34d80, 32'hc3dd438a},
  {32'hc427bc31, 32'h4392f13b, 32'h435ae956},
  {32'h413fef80, 32'hc2cdfaab, 32'hc3908ed4},
  {32'hc4a98b8a, 32'h437431c9, 32'hc3379908},
  {32'h45102d13, 32'hc28ba50b, 32'hc1a12e70},
  {32'hc487c368, 32'hc34eefce, 32'h43791bc9},
  {32'h45164d28, 32'hc389a6eb, 32'h3f9dc76c},
  {32'hc5076af8, 32'hc290c968, 32'hc261c482},
  {32'h448a84ac, 32'h4337a795, 32'hc247a18d},
  {32'hc3a2c880, 32'hc3df62dc, 32'h4376c5a6},
  {32'h42bdadb8, 32'hc2616890, 32'h43284551},
  {32'hc50c3dfa, 32'hc233f192, 32'h419b096e},
  {32'h44917ff3, 32'hc38c9dc8, 32'h42c80a5c},
  {32'hc4c25dc5, 32'hc3956c43, 32'hc33015c6},
  {32'h451ad4a7, 32'h435a637e, 32'h432a2052},
  {32'hc50df364, 32'h40e74340, 32'hc385b1bf},
  {32'h450048eb, 32'h432abaa6, 32'h43d19a8d},
  {32'hc417f46a, 32'h44117443, 32'h43ad4d59},
  {32'h44b95a4a, 32'hc2a1f06a, 32'hc3076ef8},
  {32'hc4e04c9c, 32'h435a37ac, 32'hc30a8ebb},
  {32'h42050a6c, 32'h431638b6, 32'hc35af343},
  {32'hc51d7eb8, 32'h43834ce7, 32'h43ba4046},
  {32'h44cf0ecb, 32'h429ff75b, 32'hc380362a},
  {32'hc4a18f76, 32'hc3402271, 32'h43b92d75},
  {32'h4491ae80, 32'h4376a5c2, 32'hc302eb70},
  {32'hc19e6040, 32'h43046edb, 32'hc381e9c0},
  {32'h450824ac, 32'hc346f340, 32'hbfaca014},
  {32'hc15d321b, 32'h42eca120, 32'h4334ee06},
  {32'h44343482, 32'hc3901d0e, 32'h4315205b},
  {32'hc4187b3b, 32'hc3c8734b, 32'h4356394f},
  {32'h452a04c8, 32'h42bf383d, 32'hc33c843f},
  {32'hc4dcaf0c, 32'h4303b000, 32'h42343407},
  {32'h44b9f1bc, 32'h42f08ccb, 32'h43115131},
  {32'hc515ae6e, 32'h42348ade, 32'hc3fe09d5},
  {32'h4530cff4, 32'h440c6972, 32'h432a384c},
  {32'hc4b94c6a, 32'h423bc188, 32'hc37e42a2},
  {32'h445d88f0, 32'hc3220f3d, 32'hc2ce6303},
  {32'h42d7d420, 32'h42df9659, 32'h42e44797},
  {32'h42d3a234, 32'h4373fddc, 32'hc2fbc048},
  {32'hc493eb74, 32'hc3112265, 32'hc3ed84ca},
  {32'h43f443b4, 32'hc3bbe7ee, 32'h43647656},
  {32'hc4b8c000, 32'hc2b20d3c, 32'hc43ffa44},
  {32'h44a7b488, 32'hc2c1c026, 32'h43836acf},
  {32'hc38deb80, 32'hc3be5091, 32'hc2eb8e98},
  {32'h447563d6, 32'h42c36b4e, 32'h42c3aacd},
  {32'hc4fb13ce, 32'h420f36e2, 32'hc38558f2},
  {32'h449d909f, 32'h434122e3, 32'h42f3036b},
  {32'hc500dcfd, 32'hc2b81149, 32'hc2ab4442},
  {32'h446d4148, 32'hc1d2dab9, 32'hc326272a},
  {32'hc509ab87, 32'hc3875202, 32'h420c682e},
  {32'h44dd4b72, 32'hc3042281, 32'hc2f02061},
  {32'hc41f21c3, 32'h438e17b2, 32'h43058830},
  {32'h44a99d67, 32'hc22247c8, 32'hc3f135a7},
  {32'hc51b105a, 32'h43825115, 32'h43510fd2},
  {32'h450b0cee, 32'h4341c080, 32'hc39a691f},
  {32'hc4b829ed, 32'hc296f50a, 32'h42116fd0},
  {32'h441b29cd, 32'h430a2b11, 32'hc34b6bc2},
  {32'hc4917a12, 32'h43a942ee, 32'h4389f505},
  {32'h44fc1a8a, 32'h436ac948, 32'h42202c77},
  {32'hc4f8fa8e, 32'h42889ca5, 32'hc30ce12b},
  {32'h43c8dbee, 32'hc2dc8279, 32'hc33721ac},
  {32'hc3a9b610, 32'h42c4f881, 32'h42d926aa},
  {32'h44c5010e, 32'h43b9ac31, 32'hc37cc3cf},
  {32'hc5037ae4, 32'h42a27f4a, 32'h434edbb9},
  {32'h43d723be, 32'h423ddfe0, 32'hc2c5150a},
  {32'hc4d857f9, 32'h4199e47f, 32'h41dccb04},
  {32'h449a0dca, 32'hc1590cc4, 32'h429d93c7},
  {32'hc4f99e6b, 32'hc1c2ba8a, 32'hc08df92c},
  {32'h44ebfd0b, 32'hc1d8a220, 32'hc3580a58},
  {32'hc49b2ae4, 32'hc3fedcd8, 32'hc1b7e30e},
  {32'h44139e96, 32'hc2330f34, 32'h435ff43f},
  {32'hc480c74a, 32'hc351e2c8, 32'h4423c8fd},
  {32'h4481d368, 32'h429d690e, 32'h4384196d},
  {32'hc4de6600, 32'h433f227c, 32'hc342b072},
  {32'h448208d6, 32'hc3d657ff, 32'h42c126eb},
  {32'hc50806d0, 32'hc2c2e51c, 32'hc2de71ed},
  {32'h450e2995, 32'h43722727, 32'h42ff96f1},
  {32'hc44a6a04, 32'hc2d1481e, 32'hc34c117f},
  {32'h44fc180e, 32'hc1f359ec, 32'h42d7dc19},
  {32'hc50253cc, 32'hbfcc976c, 32'hc3cfe3fa},
  {32'h4438c4af, 32'hc3be3385, 32'h43dcdbab},
  {32'hc3d7e132, 32'h43b08e83, 32'h429d69ae},
  {32'h4401231b, 32'h43897d34, 32'hc314c991},
  {32'hc500cd55, 32'hc359d20c, 32'h4368ac3a},
  {32'h44f5fd38, 32'hc365ed3a, 32'h42aa9f4c},
  {32'hc416ea5c, 32'h42bf8102, 32'h43b14159},
  {32'h43e9d212, 32'hc299737c, 32'hc38dd073},
  {32'hc45f819f, 32'h4302365c, 32'hc4099650},
  {32'h44b14710, 32'hc39619e1, 32'h43017cee},
  {32'hc4da0021, 32'hc292d13f, 32'hc2f2c7dc},
  {32'h44b64843, 32'hc428b86f, 32'hc2504558},
  {32'hc51b6aa2, 32'h4235d87b, 32'h4269380e},
  {32'h451fa95a, 32'h42414e09, 32'h425a6d1e},
  {32'hc40c9888, 32'h432b5cee, 32'hc3ea78e8},
  {32'h44f4f9f2, 32'hc363f8fb, 32'h43008d12},
  {32'hc3abca28, 32'h420cf54e, 32'hc3b75830},
  {32'h44d1b533, 32'h43a15139, 32'h4285f72f},
  {32'hc3ea01aa, 32'hc3b55715, 32'hc343e2f8},
  {32'h4510b252, 32'hc38b9fe2, 32'hc377f5ec},
  {32'h41a8bfc0, 32'hc2928ee3, 32'h43560c21},
  {32'h444fc582, 32'h42beb7cf, 32'h41e22245},
  {32'hc511d334, 32'hc2b6c339, 32'h4319edd7},
  {32'h44eae9c9, 32'hc3516b07, 32'hc2f1051c},
  {32'hc515c1b6, 32'hc36e62e6, 32'h43149306},
  {32'h44bcbeb6, 32'hc403924f, 32'h43022fda},
  {32'hc4972844, 32'h43ef2adb, 32'hc2218e2a},
  {32'h4506ef16, 32'h41dabd2e, 32'hc40d992e},
  {32'hc509c7ec, 32'h43fdc869, 32'hc3897898},
  {32'h4514f48a, 32'hc30a1d55, 32'hc20a51e5},
  {32'hc500ff4f, 32'h4349b850, 32'hc391cdd1},
  {32'h43df72f2, 32'hc342b220, 32'hc1e01f00},
  {32'hc32ca249, 32'h43a3aaf2, 32'hc2a8edf8},
  {32'h44cc4b3c, 32'hc3ebbcdf, 32'hc2f86d8a},
  {32'hc4a5a961, 32'h434819a2, 32'h43db05a5},
  {32'h44c48e78, 32'h42461244, 32'hc2f66252},
  {32'hc4453066, 32'hc2b5ad51, 32'h43b316b9},
  {32'h45031493, 32'hc37b7d42, 32'hc29efa09},
  {32'hc3b30b5a, 32'h4287ed66, 32'h438876fb},
  {32'h432f7bae, 32'hc2cf767b, 32'hc40d7b60},
  {32'hc4892b3e, 32'h43b63ca4, 32'h4304ea1e},
  {32'h450498d7, 32'hc2f53175, 32'hc395a01e},
  {32'hc4cc9eea, 32'hc21dc4fe, 32'hc380c3ab},
  {32'h439a5a60, 32'h43815208, 32'hc36b4d8a},
  {32'hc48bc547, 32'h426a23ba, 32'h424db4a7},
  {32'h445726d3, 32'hc396c273, 32'h423e96bf},
  {32'hc3e25308, 32'h4338f683, 32'hc329d7e5},
  {32'h448122a0, 32'hc2e4fa7a, 32'hc36ac236},
  {32'hc428f63c, 32'h432ac4c7, 32'h42dd414e},
  {32'h44c8e534, 32'h439c30a3, 32'hc1d8794e},
  {32'hc50ac257, 32'hc2cb432e, 32'h43d50f94},
  {32'h450f53b8, 32'hc3c45a7b, 32'h43347f47},
  {32'hc4cede1c, 32'h41aa0612, 32'h43b38b63},
  {32'h45056324, 32'hc2b614e5, 32'hc08fe4dc},
  {32'hc40d6664, 32'hc30ac389, 32'h434087b5},
  {32'h43d87474, 32'h43233231, 32'hc2225742},
  {32'hc5063a42, 32'h43028a93, 32'h438c84c6},
  {32'h44d9aa62, 32'hc19d14e6, 32'hc30a129a},
  {32'hc48f1978, 32'hc3df2d1f, 32'h42e8c842},
  {32'h450628f3, 32'h415ee628, 32'hc2c0548d},
  {32'hc442e6ba, 32'hc2ccc4c6, 32'h43065fb0},
  {32'h44d44b69, 32'h426b37a9, 32'hc2b6075c},
  {32'hc488d11b, 32'h4200ddbe, 32'hc2abf6ed},
  {32'h44f670a9, 32'hc359fb1b, 32'h422f6441},
  {32'h41164600, 32'h43e5033d, 32'h43a360c0},
  {32'h43a61efa, 32'hc2b63d19, 32'h437b6c93},
  {32'hc5020882, 32'h4295b136, 32'hc381803f},
  {32'h44a1831c, 32'hc28197e7, 32'hc32ffd58},
  {32'hc4f8241d, 32'hc4036021, 32'h43181911},
  {32'h44278635, 32'hc38aeb0c, 32'h4312abc8},
  {32'hc4dc69e6, 32'hc329a604, 32'h435c9e30},
  {32'h4500ae2f, 32'hc3755a90, 32'h438a2e8d},
  {32'h448f4924, 32'hc1d2ac50, 32'h430831c7},
  {32'hc3457ca8, 32'hc3bb8c40, 32'h43a2a4c6},
  {32'h43c450b0, 32'hc3e66368, 32'hc2c9cc81},
  {32'hc3bc0792, 32'h422b9066, 32'h42f9540a},
  {32'h44ff3d33, 32'hc337b4d0, 32'hc3d9e95e},
  {32'hc51a8a47, 32'hc18a4dff, 32'h42b97886},
  {32'h4506bf1c, 32'hc39d24c6, 32'hc33167b1},
  {32'hc4665180, 32'h42f868c8, 32'hc368f3da},
  {32'hc2064340, 32'h43a27a0b, 32'hc3805126},
  {32'h420ebe20, 32'h42ff764e, 32'hc2d802c1},
  {32'h441e7a76, 32'hc311aa0e, 32'hc348a65d},
  {32'hc4241a5a, 32'hc1da962e, 32'hc29cf8ae},
  {32'h44da280e, 32'hc2833c57, 32'h4293b877},
  {32'hc4aa5498, 32'hc24d8972, 32'hc3755211},
  {32'h4482acf9, 32'hc2976667, 32'h43907af8},
  {32'hc4fdc322, 32'hc247e418, 32'hc3136440},
  {32'h443925ec, 32'hc2f010a3, 32'hc3669a2c},
  {32'hc4f655c1, 32'h439bf813, 32'h43e44d6b},
  {32'h4421ad75, 32'hc216370d, 32'h43f11bcb},
  {32'hc4d72018, 32'hc23d69a9, 32'h43b119b6},
  {32'h4478568f, 32'hc2066ac5, 32'h43128bde},
  {32'hc4a3a533, 32'hc33350c4, 32'hbf41d877},
  {32'h4457a36f, 32'h423417ad, 32'hbff2344f},
  {32'hc508bb28, 32'hc183fb8c, 32'h426d4579},
  {32'h45093887, 32'hc3a03e9f, 32'hc309b6ff},
  {32'hc500a9b4, 32'hc3c30e44, 32'h436edab4},
  {32'h44a93831, 32'h42c0d957, 32'hc2ab55f2},
  {32'hc38dbc75, 32'h429f116d, 32'h42736f7b},
  {32'h45095076, 32'h4383275d, 32'hc3172e9f},
  {32'hc502ef7f, 32'hc221b2e1, 32'h434bc20b},
  {32'h44ac07dc, 32'h4392f287, 32'hc308910f},
  {32'hc438577e, 32'hc3c31d92, 32'hc310ca75},
  {32'h44be0cf1, 32'h43118cfc, 32'h435df1a5},
  {32'hc4bbd47f, 32'h42b14aba, 32'hc37a24f3},
  {32'h44498d93, 32'h429f9459, 32'hc2e1ad1d},
  {32'hc48f51d7, 32'h40d6f16b, 32'hc1cf2ffe},
  {32'hc2af67e0, 32'h41da60c4, 32'h42290a52},
  {32'hc4444d70, 32'hc2d00b38, 32'h4324ec42},
  {32'h45155411, 32'hc3bcc0d0, 32'hc29b2b31},
  {32'hc4ab466b, 32'h43842bfb, 32'hc309f54b},
  {32'h448d490e, 32'hc2612aae, 32'h43806f43},
  {32'hc4e16686, 32'hc2ab13d8, 32'hc37a859b},
  {32'h44b05748, 32'h4307ee3b, 32'h438aa6b1},
  {32'hc5146eae, 32'hc3597e62, 32'hc3542758},
  {32'h43b73d36, 32'h42588d36, 32'h426f1e89},
  {32'hc4f98360, 32'h4386211d, 32'h4384e965},
  {32'h44a0be42, 32'hbf6296c4, 32'h42a02b4c},
  {32'hc357f350, 32'h42d0f29a, 32'hc2adf206},
  {32'h45087fae, 32'h4330b12c, 32'h42c15142},
  {32'hc4e45acc, 32'h437d7196, 32'hc29ce112},
  {32'h44929522, 32'h4311525a, 32'h434554df},
  {32'hc4951c60, 32'h43a0be1f, 32'hc37d6493},
  {32'h451a91a9, 32'hc2cf16e7, 32'h434fad1c},
  {32'hc3fc3090, 32'h430acbdc, 32'h42322f84},
  {32'h44a69a47, 32'h42ebb5e1, 32'h4325bbef},
  {32'hc415a9a0, 32'h432a58d9, 32'hc3c6eb77},
  {32'h44666930, 32'hc12e3a56, 32'hc33b3806},
  {32'hc478c595, 32'hc3a0ec35, 32'hc21e056f},
  {32'h42447a84, 32'h43c8ca95, 32'h406711f3},
  {32'hc4017e31, 32'h43401886, 32'hc39365b9},
  {32'h451907f2, 32'hc3b0e8d4, 32'h42ae8439},
  {32'hc3645160, 32'hc338855d, 32'hc3ce9cc0},
  {32'h45078723, 32'h4360b4ff, 32'hc2e6c3a0},
  {32'hc4637931, 32'h429d910d, 32'hc235d42a},
  {32'h446fcaa0, 32'h3f3b3408, 32'hc3ab7954},
  {32'hc50c307c, 32'hc38469e9, 32'hc273f55d},
  {32'h44acfa37, 32'hc291fa99, 32'hc2873830},
  {32'hc440dc19, 32'h43224df8, 32'hc3337547},
  {32'h4503a217, 32'h42b7f028, 32'h4300e980},
  {32'hc4f155b8, 32'hc31f1b92, 32'hc2799a2e},
  {32'h43a989ff, 32'h43bc3cf0, 32'hc1fa45e5},
  {32'hc35712b4, 32'hc2d6bc03, 32'h420860f1},
  {32'h449eb07e, 32'h427ab166, 32'h42f96a38},
  {32'hc4e1dfaf, 32'hc345bae6, 32'hc2f1de4f},
  {32'h44055aca, 32'hc200986a, 32'h431ad1d5},
  {32'hc448480e, 32'hc29d854a, 32'h43a83134},
  {32'h44509273, 32'hc32eb8b6, 32'hc315b372},
  {32'hc4f03677, 32'h4202d990, 32'hc2f7b02e},
  {32'h44d62b5c, 32'hc36f8cdc, 32'h4383cbb0},
  {32'hc4184bd2, 32'hc310b351, 32'h424d8a44},
  {32'h44de69a8, 32'hc20afd53, 32'h43f7b7a5},
  {32'hc507001f, 32'hc0fb0c3a, 32'hc39fa0b7},
  {32'h44ecb663, 32'h431021e4, 32'hc1a92a10},
  {32'hc45c1c73, 32'h441eabbb, 32'hc39f5a8d},
  {32'h440fbce5, 32'hc3bcf0ed, 32'hc298f41d},
  {32'hc3a26a80, 32'h42f0e38e, 32'h42ce54c0},
  {32'h4376aa4c, 32'hc2853ecf, 32'h43401143},
  {32'hc515db50, 32'hc2160366, 32'hc39b933c},
  {32'h44cf47f7, 32'hc310fd71, 32'h41ee7cbb},
  {32'hc51b4028, 32'hc14744f1, 32'hc347f7cd},
  {32'h44913500, 32'hc3750e99, 32'h43c066c3},
  {32'hc4ce5076, 32'h4235249a, 32'h431216c2},
  {32'h447a99ed, 32'h4373ac6d, 32'hc35362b4},
  {32'hc4f31b09, 32'h44478082, 32'h4347cb9c},
  {32'h444651bd, 32'hc36be3c2, 32'h4370bae6},
  {32'hc38479f0, 32'h41bc8207, 32'h4132882c},
  {32'h449c1b4d, 32'h422151e2, 32'h4371a345},
  {32'hc391c3fe, 32'h41906afd, 32'hc1afa667},
  {32'h44fdbdc7, 32'hc3e07297, 32'hc301e94d},
  {32'hc457929a, 32'hc33cc5be, 32'h43089f18},
  {32'h4390f540, 32'h432dcdc3, 32'hc2185dfe},
  {32'hc5044e11, 32'hc30ed3c9, 32'hc36b0ea2},
  {32'h445759b8, 32'h43c5221a, 32'h439941fe},
  {32'hc474441a, 32'hc3ef0025, 32'h438b839d},
  {32'h446491e6, 32'hc23ca79b, 32'h42241d48},
  {32'hc3536eb0, 32'hc3a2cd5f, 32'h43834e0b},
  {32'hc2876690, 32'hc3095f5f, 32'h41e591f4},
  {32'hc5052b2a, 32'hc2fcce92, 32'h42eea3fe},
  {32'h43da2290, 32'hc3236cfc, 32'hc225b7a5},
  {32'h42bd2880, 32'hc32033de, 32'h435c9c67},
  {32'h44f8b3ec, 32'h41870326, 32'h43c51f82},
  {32'hc4e64843, 32'h428c112d, 32'h429d7955},
  {32'h44f6323b, 32'h4323b8db, 32'hc1d34a6d},
  {32'hc50e9148, 32'h43152a75, 32'h41b4837a},
  {32'h44ed643c, 32'hc305e345, 32'h43a121cc},
  {32'hc3ed5b68, 32'h422417be, 32'hc2c20721},
  {32'h44c67213, 32'hc20c6188, 32'hc3018beb},
  {32'hc3bc67dc, 32'hc2e57e03, 32'hc2af3730},
  {32'h44c31969, 32'hc1a29bd7, 32'h42318c1f},
  {32'hc4a3324f, 32'hc3845c37, 32'h436d19dc},
  {32'h4478f5bf, 32'hc30b9adc, 32'h42b893bd},
  {32'hc4a1acb6, 32'hc38545be, 32'hc303ac4e},
  {32'h43ccf2f4, 32'h4347b2af, 32'hc23d416c},
  {32'hc39a495c, 32'h42bc3292, 32'hc249bc32},
  {32'h44b582dc, 32'hc21ea781, 32'h42fafa32},
  {32'hc4926b14, 32'h43137628, 32'h437b04a3},
  {32'h45111408, 32'hc324d31c, 32'hc2568f80},
  {32'hc499a1d6, 32'h428f6ab4, 32'h434122db},
  {32'h44ab523f, 32'h41b57e58, 32'h41cd5ad0},
  {32'hc4dae25c, 32'h43a89509, 32'h4328c291},
  {32'h450f270c, 32'hc269bd29, 32'h43187534},
  {32'hc48598dc, 32'h4289b8e2, 32'h3ff85aba},
  {32'h4479a06d, 32'hc3390242, 32'hc2b19ac1},
  {32'hc4a0038a, 32'h42dfe816, 32'h43f543a0},
  {32'h44712f88, 32'hc33c67f2, 32'hc30cd26b},
  {32'hc30d5350, 32'h3ef4c700, 32'hc38c67ed},
  {32'h44cff73b, 32'hc28210b1, 32'hc37f7db8},
  {32'hc3fdccd8, 32'hc3b766fc, 32'hc4115096},
  {32'h44aa8880, 32'h43013791, 32'hc3b492cf},
  {32'hc4b4a81e, 32'h42fb7506, 32'h435c1c2a},
  {32'h44ea629c, 32'h43c33bf4, 32'h43498c93},
  {32'hc316a8d8, 32'hc3214c51, 32'h4290f115},
  {32'h44940574, 32'h42d0d662, 32'h42a2cb1f},
  {32'hc4e07f73, 32'hc32a3207, 32'h42f9d01c},
  {32'h44833b86, 32'h43851707, 32'h42fa1b2b},
  {32'h433114d4, 32'hc38ff828, 32'hc2ab7d55},
  {32'h44727e33, 32'h41889113, 32'hc33712a6},
  {32'hc4d912ff, 32'h4298deff, 32'hc387ff1d},
  {32'h4500242e, 32'hc2a9b18c, 32'hc2d9794a},
  {32'hc3147e72, 32'h434e2f95, 32'h410991de},
  {32'h43e626d0, 32'h43b9eed3, 32'h41964468},
  {32'hc4d754f3, 32'h42d0e635, 32'h430e439b},
  {32'h4420be84, 32'h4204985a, 32'h413e2b88},
  {32'hc486e498, 32'hc34177ee, 32'hc232f855},
  {32'h44a0ba19, 32'hc37f43f3, 32'h42c97c48},
  {32'hc36bf240, 32'h4279c771, 32'h431ae46e},
  {32'h44e5bae9, 32'h431d9dd2, 32'h4212eb3d},
  {32'hc4b13abb, 32'h438c8461, 32'hc2833793},
  {32'h44264b3e, 32'hc200426b, 32'hc3144aea},
  {32'hc48615e7, 32'h41ba490c, 32'hc3929fc4},
  {32'h43e4a968, 32'h428d96f6, 32'h43b2158a},
  {32'hc473b7b6, 32'h4216a831, 32'h434fb7c6},
  {32'h4464207c, 32'hc34e58a3, 32'hc38cbd7b},
  {32'hc503bdea, 32'h43a3bc40, 32'hc3a478f0},
  {32'h44bb31f6, 32'hc2c37f40, 32'h435bd8e0},
  {32'hc505b3e7, 32'h432394d1, 32'h438e0732},
  {32'h441a8798, 32'hc2e2a5a9, 32'h422251f8},
  {32'hc3cfb5f8, 32'hc19ed7b9, 32'h42db1747},
  {32'h43f0a9ef, 32'hc2f66f34, 32'h43141c9b},
  {32'hc4cfe015, 32'hc3eb1bcc, 32'hc15e8b0d},
  {32'h445fee4d, 32'hc2b2b4a6, 32'h3eea9d2e},
  {32'hc509fac1, 32'hc3cc1b75, 32'h43a6409a},
  {32'h449e3986, 32'hc3a49876, 32'h431c89e7},
  {32'hc4ffd2b3, 32'h42b6cb46, 32'hc372fc11},
  {32'h44c4af68, 32'h43842afc, 32'h432003c0},
  {32'hc488e1a9, 32'hc2806815, 32'h42b6e088},
  {32'h44d46e54, 32'hc3651faa, 32'hc2e0bfb6},
  {32'hc4af7608, 32'hc3289ea9, 32'hc38be053},
  {32'h450210b9, 32'hc300de47, 32'h437e6352},
  {32'hc3f9a1ec, 32'hc2c1159a, 32'h4387126c},
  {32'h450ae62f, 32'h4394d4d5, 32'hc397d8bd},
  {32'hc4b1def7, 32'h436890d3, 32'hc3acc527},
  {32'h447126e2, 32'h42908f87, 32'h438c8b5f},
  {32'hc4b4dd5f, 32'h434a029a, 32'h4296a864},
  {32'h439c36b8, 32'hc33e07ff, 32'h421b49e1},
  {32'hc4fe136f, 32'h42b91788, 32'h409bf2d2},
  {32'h44c50e2b, 32'hc3a067ce, 32'hc23e4726},
  {32'hc3893d80, 32'h43298b6c, 32'h4336d986},
  {32'h44f14df5, 32'hc327623d, 32'hc248e548},
  {32'hc4921919, 32'h43b2f47d, 32'h43300b6d},
  {32'h44fe1a10, 32'h422fc501, 32'hc2b64da6},
  {32'hc3dcd4f6, 32'hc2bcb921, 32'h42ea11d9},
  {32'h44f34712, 32'hc22e3d08, 32'hc332faf5},
  {32'hc4953bcc, 32'h422d99da, 32'hc2e3143b},
  {32'h443ff395, 32'hc130b7f7, 32'hc2500c35},
  {32'hc482a9b3, 32'hc3177a50, 32'h43f882c0},
  {32'h437b46a8, 32'h438b97a4, 32'h43038aca},
  {32'hc4cf75ca, 32'h42e1d578, 32'hc1b37189},
  {32'h44838324, 32'hc1bb72d6, 32'h43cec27c},
  {32'hc3cba3b5, 32'hc25a296e, 32'h4393b96b},
  {32'h44a1ff6b, 32'h44199df9, 32'h415d3bec},
  {32'hc4255c18, 32'h417adf42, 32'h40a92630},
  {32'h44457fa2, 32'h429cf1f8, 32'hc39b4854},
  {32'hc4b9e2cd, 32'h4354209e, 32'hc3446f0f},
  {32'h448f0049, 32'hc34ab098, 32'h4293f1e2},
  {32'hc4bbeac3, 32'hc380d06b, 32'h43668035},
  {32'h44bf3c33, 32'hc35de62a, 32'h4255601e},
  {32'hc4c9ec1d, 32'h43c0f923, 32'hc30a6d6f},
  {32'h45018108, 32'hc2100c32, 32'hc10c0616},
  {32'hc2ba3520, 32'h41a6b5e4, 32'hc247f8c0},
  {32'h446200b6, 32'h432e495c, 32'h4314dd76},
  {32'hc3c2f545, 32'hc26927b9, 32'h42e34d83},
  {32'h43f478d4, 32'hc2ffea9d, 32'hc38c8b25},
  {32'hc4fb5a10, 32'h42fb9fad, 32'h4323c549},
  {32'h4473e946, 32'h43375864, 32'hc2fa9e04},
  {32'hc4962387, 32'hc3289738, 32'hc3635895},
  {32'h4284a208, 32'h438dfd29, 32'h433fcaa2},
  {32'hc4daf21b, 32'hc3c70732, 32'h433cb024},
  {32'h44c6a59d, 32'hc3e0e34f, 32'hc2806066},
  {32'hc505d3fb, 32'hc33960f3, 32'h4169fd9b},
  {32'h448af0e2, 32'h43d484f2, 32'h43a93d03},
  {32'hc463e960, 32'h42033982, 32'h438d2ed8},
  {32'h4328a8d0, 32'hc1e709f1, 32'hc2e1ca1b},
  {32'hc4af6a34, 32'hc3b2609a, 32'hc3b45636},
  {32'h4455de52, 32'hc36d78be, 32'hc3d5103f},
  {32'hc4f5f42d, 32'hc33c19b7, 32'hc3bcca75},
  {32'h44bedf54, 32'hc337e49e, 32'hc21b2a5d},
  {32'h41905500, 32'h4306c434, 32'hc335670f},
  {32'h44d1183d, 32'hc33a8cc8, 32'h432246bc},
  {32'hc421eb66, 32'h43f7bcac, 32'h42941e37},
  {32'h44dabdbe, 32'hc2d1e29a, 32'h41c336d7},
  {32'hc3327d10, 32'hc1f1214c, 32'hc3919ca6},
  {32'h448beaa1, 32'h43028f1d, 32'h43fa43d6},
  {32'hc50ac918, 32'hc2128f08, 32'h42a81bb8},
  {32'h450d3ffa, 32'hc330d658, 32'h40af01d8},
  {32'hc5019b39, 32'hc3b0f52d, 32'h4323d80c},
  {32'h440875d8, 32'h43937fdc, 32'hc25e4c2a},
  {32'hc481f854, 32'hc345cb53, 32'h4334a6b9},
  {32'h4426727c, 32'hc3fdd8e4, 32'hc3f41235},
  {32'hc44b6f1a, 32'hc2df1d9c, 32'hc2b18ece},
  {32'h44a8f1cb, 32'h402e02f4, 32'hc1db4c31},
  {32'hc5024dca, 32'h42a45ae1, 32'h4387ff65},
  {32'h44576a28, 32'h43346e32, 32'hc35bc62b},
  {32'hc4273327, 32'h43648930, 32'h436fcbad},
  {32'h44580f4b, 32'hc3c41071, 32'hc1c3427c},
  {32'hc3e6f6f6, 32'hc318dae3, 32'h41b0d9be},
  {32'h44f49916, 32'hc33a3d83, 32'hc0570ee9},
  {32'hc3ac1942, 32'hc361c62b, 32'h42d947bd},
  {32'h4459c724, 32'hc303b49d, 32'h4286c5ff},
  {32'hc443eed5, 32'hc36b57f8, 32'h4380b518},
  {32'h442ffdfd, 32'hc2b24099, 32'hc2f6f34a},
  {32'hc4abe984, 32'h41f4fbba, 32'h439f326d},
  {32'h44640e1c, 32'h4412a2f9, 32'h428bb760},
  {32'h4385d84c, 32'hc343a20b, 32'hc2af141d},
  {32'h44b0d1df, 32'hc38051ef, 32'hc3a52d9a},
  {32'hc502a057, 32'h42d4ef70, 32'hc22b0bd3},
  {32'h44d8df20, 32'hc2f47aba, 32'hc35317ad},
  {32'hc48c16b0, 32'hc37754d4, 32'h4347d59e},
  {32'h43d77da4, 32'hc22a00a4, 32'h436159ed},
  {32'hc507bc42, 32'hc3a7ece4, 32'h43888a76},
  {32'h44c4df76, 32'h41866bd0, 32'h439960af},
  {32'hc4ba67f8, 32'hc24c0083, 32'h435e4259},
  {32'h44ef2121, 32'h41f45187, 32'hc3b391b7},
  {32'hc43f2723, 32'h43d37e27, 32'h429b76e1},
  {32'h4507d994, 32'h428e4c0e, 32'hc2cffb6f},
  {32'hc4eae7c0, 32'h438a8a31, 32'h43a3d46a},
  {32'h4339f3a0, 32'hc1a1d3f0, 32'hc33d7a9f},
  {32'hc4f31230, 32'hc2a48d00, 32'h43805c55},
  {32'h4483b047, 32'h43cbb5cc, 32'h43971ce7},
  {32'hc4be2cf3, 32'hc3223e27, 32'h42e2f951},
  {32'h44aa7aee, 32'h4282a05d, 32'hc3043878},
  {32'hc483eacf, 32'h431798bc, 32'h441d9b3d},
  {32'h44511d10, 32'hc31281a8, 32'hc40e06e2},
  {32'hc43eac62, 32'hc309fc08, 32'h43a111f2},
  {32'h45063178, 32'h430058e0, 32'hc3c8922a},
  {32'hc364d348, 32'hc3b781e7, 32'h42c7efae},
  {32'h44a9c5ef, 32'h439280be, 32'hc33d2740},
  {32'h41a19380, 32'hc231ebe2, 32'hc1f25957},
  {32'h44523df2, 32'hc32a7dc3, 32'h431472a7},
  {32'hc498df0a, 32'hc327913c, 32'h426c81ca},
  {32'h439e1764, 32'h43129aea, 32'h4384a611},
  {32'hc4195461, 32'hc1b6aac6, 32'hc394f9ba},
  {32'h44b0327c, 32'hc36c0302, 32'h4379f893},
  {32'hc4e3712d, 32'h429840f9, 32'h43fab78b},
  {32'h4486f57f, 32'hc253b1b2, 32'hc2143cd0},
  {32'hc4ccfd27, 32'h42a61da8, 32'h42adf121},
  {32'h45048b2c, 32'h42255031, 32'h43d05a55},
  {32'hc44cb0e2, 32'hc2dd43e1, 32'hc3a3b9b0},
  {32'h439f83d6, 32'hc2ed4abd, 32'hc3b030e2},
  {32'hc4f43fac, 32'h430a02c6, 32'h4246f7d6},
  {32'h44b52f7b, 32'h41831510, 32'h43768ba1},
  {32'hc5119aa4, 32'h43a9f5f2, 32'h43ceed71},
  {32'h438a7321, 32'hc310d091, 32'h4319e682},
  {32'hc47d0342, 32'hc1df241c, 32'hc351f11a},
  {32'h450bde88, 32'h439aedfe, 32'hc21e26c1},
  {32'hc4fee4aa, 32'h4388f8ad, 32'hc3024bea},
  {32'h44d2558c, 32'hc2b978f2, 32'hc24295e4},
  {32'hc4dca158, 32'h405d8d20, 32'h4434d4c3},
  {32'h43fa0297, 32'hc356bd2d, 32'h43c1686e},
  {32'hc4e33d3a, 32'h435e1cb3, 32'hc41b5bca},
  {32'h4508d9e3, 32'hc31a8384, 32'hc38ff187},
  {32'h43b17404, 32'hc39dea9c, 32'hc30e387b},
  {32'h45224782, 32'hc2f0d918, 32'hc38da772},
  {32'hc4623af2, 32'hc3c8742b, 32'hc30c7639},
  {32'h4511b77b, 32'h428ad942, 32'h421e22d1},
  {32'hc45ec94c, 32'hc2f5ccf1, 32'hc272ded8},
  {32'h44f6fdfc, 32'h43204eae, 32'h43374baa},
  {32'hc4ebe7b0, 32'hc3e11885, 32'h423ceaaa},
  {32'h44b4a9d6, 32'hc1a6a665, 32'h43aaa680},
  {32'hc49b5bcd, 32'hc3a9fc29, 32'h4343b675},
  {32'h440af7ee, 32'h432331ae, 32'hc2778183},
  {32'hc4dde89e, 32'h4370745a, 32'h43df3e57},
  {32'h4459bf1f, 32'h42d42056, 32'hc2b88b77},
  {32'hc3be4e4d, 32'h42da6b48, 32'h43152c32},
  {32'h451f10d0, 32'hc34f727d, 32'hc24158f3},
  {32'hc4171448, 32'hc31991f7, 32'h3ea0cfd7},
  {32'h4493f45f, 32'h3ff51e40, 32'hc34a6eaa},
  {32'hc4e59e40, 32'h43d237bc, 32'hc2cc7dab},
  {32'h44179716, 32'hc2f505ac, 32'hc305df6c},
  {32'hc490caf7, 32'h42635a41, 32'hc34cad86},
  {32'h44721364, 32'hc3b0c72d, 32'hc34ca1d2},
  {32'hc40b123e, 32'hc3d7ef56, 32'hc27b35aa},
  {32'h44a98dd5, 32'hc0ea915a, 32'hc20c3652},
  {32'hc4c5b827, 32'hc3bca989, 32'hc31e92c5},
  {32'h448d8a57, 32'h43af0c16, 32'hc27a5032},
  {32'hc47613e4, 32'h4372047d, 32'hc1d389f2},
  {32'h44cf59b4, 32'hc0c249a9, 32'hc3665503},
  {32'hc4f82e02, 32'hc307ebdd, 32'hc2b7b9b3},
  {32'h4416cad3, 32'hc2a7071e, 32'hc33fb042},
  {32'hc3bda924, 32'h4328e9d6, 32'h4394eb0b},
  {32'h450983d7, 32'hc2c7247d, 32'h3ef60890},
  {32'hc50b52a8, 32'h4339a79e, 32'h400975c2},
  {32'h44c970af, 32'h437e0423, 32'hc39eb442},
  {32'hc49cf78c, 32'h437cefb4, 32'hc2dfe20d},
  {32'h44a3e77c, 32'hc234ca07, 32'hc12b646c},
  {32'hc3e60470, 32'hc1076c25, 32'h43f4a0bd},
  {32'h44829c88, 32'h4200f6f1, 32'hc38d68e2},
  {32'hc4f45986, 32'hc35878a5, 32'hc2174dd4},
  {32'h44ed4e8a, 32'h433e8065, 32'h42702f93},
  {32'h42c61438, 32'hc2bc287d, 32'hc2f6d6c4},
  {32'h43f4ec72, 32'h43a6545f, 32'h43394469},
  {32'hc4d7c5d2, 32'h43243d43, 32'hc42c3f70},
  {32'hc25dcca0, 32'h424f0d00, 32'h43a0a5a9},
  {32'hc390fdb0, 32'h438a978e, 32'hc345bfb5},
  {32'h43d6cc30, 32'h4339b477, 32'hc179ca75},
  {32'hc3c9ea44, 32'hc0256b87, 32'hc18d6505},
  {32'h42eac920, 32'hc421c7b3, 32'hc356d3c8},
  {32'hc36d4710, 32'hc33e9d5f, 32'h41b7f83a},
  {32'h44eed943, 32'hbf0438b0, 32'hc301b3d3},
  {32'hc4dbf557, 32'hc33f300e, 32'hc2e615c3},
  {32'h447cf35d, 32'h420f21dd, 32'h44274633},
  {32'hc48159e1, 32'h4309fdc0, 32'h431ee4d6},
  {32'h450a5e12, 32'hc25678f8, 32'hc3032fca},
  {32'hc3ec2f79, 32'hc40a16a4, 32'hc1bd2ae9},
  {32'h445a842b, 32'h42955849, 32'h43f5eedc},
  {32'hc505829a, 32'hc3cef8bc, 32'h42b75be2},
  {32'h441072a6, 32'h435d95a1, 32'h438b98cf},
  {32'hc4da52ae, 32'hc3853d55, 32'h42cc0176},
  {32'h44e2f24a, 32'h434c54fc, 32'h4355a130},
  {32'hc42bc3de, 32'hc367325d, 32'h40a5bc44},
  {32'h44bab727, 32'hc39aa0df, 32'h42ca4f25},
  {32'hc3b7d27c, 32'h436962e3, 32'hc297d963},
  {32'h44e778f1, 32'hc369b4f3, 32'hc3364388},
  {32'hc3064970, 32'h423ab933, 32'hc1712fe4},
  {32'h44ce870a, 32'hc2e6e4c3, 32'hc3e8c031},
  {32'hc4ed73f7, 32'hc26b056f, 32'hc3a572c5},
  {32'h44dfd10d, 32'h4381befc, 32'hc3b82f71},
  {32'hc40c9778, 32'hc31cd9d6, 32'h436d3d72},
  {32'h441bd573, 32'h432b1b11, 32'hc31bf63c},
  {32'hc4c1ee88, 32'hc3af55cb, 32'h436bc47f},
  {32'h450c39bf, 32'h42ae8040, 32'hc0a8a490},
  {32'hc46e4234, 32'hc41d585c, 32'h418b64f0},
  {32'h450af4f9, 32'hc39ddc87, 32'h43efd8cf},
  {32'hc49d73a6, 32'h41df14b7, 32'h43d322e7},
  {32'h43b73e7e, 32'hc3de9e70, 32'h412ef100},
  {32'hc4cbf160, 32'h42cb72bb, 32'h42e70bbb},
  {32'h44ae4a95, 32'h42db80fe, 32'hc3541d69},
  {32'hc4f14af4, 32'h4222e12d, 32'hc2fbbcd1},
  {32'h43ff5bf8, 32'h42379760, 32'h42b36bbc},
  {32'hc42084af, 32'h437591a5, 32'h4357130f},
  {32'h43f90ce4, 32'h4380e0b7, 32'hc36df958},
  {32'hc524d1df, 32'hc3c07243, 32'h42eb52f5},
  {32'h44fca6e7, 32'hc3b8cb32, 32'h427d4a18},
  {32'hc28f37c0, 32'hc3755595, 32'hc3c6e932},
  {32'h441771b2, 32'h434b5196, 32'h43c243e6},
  {32'hc473befc, 32'hc32d155b, 32'hc2aaf56f},
  {32'h43c603c8, 32'hc359822a, 32'hc2fdcf0c},
  {32'hc4aebb1b, 32'h433b5ca9, 32'h4412170c},
  {32'h44e08e2e, 32'h42cabda5, 32'hc2e79718},
  {32'hc508db6f, 32'h42491c70, 32'h43276755},
  {32'h4476274f, 32'h42f90921, 32'hc4267268},
  {32'h43043218, 32'hc3a3a134, 32'h4375aef7},
  {32'h4488ed33, 32'h439f6ca9, 32'hc3b2a216},
  {32'hc31ed346, 32'h43241ac8, 32'hc3209ebc},
  {32'h4482ab63, 32'h42398f4f, 32'hc38c50b1},
  {32'hc4ebc1a5, 32'hc2f34256, 32'hc3bf4119},
  {32'h44a1246b, 32'hc2c76b65, 32'h41e89e60},
  {32'hc4c7f5e8, 32'h4393a477, 32'hc3302ccc},
  {32'h44a98518, 32'hc3452cde, 32'hc2cc1ba2},
  {32'hc41c4980, 32'hc2c48c68, 32'hc339a93a},
  {32'h44cb7999, 32'hc309999a, 32'hc324c4f0},
  {32'hc4e7a17f, 32'hc3dbdf73, 32'hc3731233},
  {32'hc286bdb8, 32'hc216dd49, 32'h435cfbc0},
  {32'hc47c97e4, 32'hc355ed75, 32'hc3b3e6e2},
  {32'h438eadd0, 32'hc3a3b5b5, 32'h43d437f3},
  {32'hc500c9df, 32'h4201ca92, 32'hc347da0b},
  {32'h44978fdc, 32'h422af481, 32'h438e42ff},
  {32'hc4234a78, 32'hc354dda9, 32'hc3b584af},
  {32'h444ef731, 32'h43354c7d, 32'h43a7a4cc},
  {32'hc3bbf730, 32'hc2e4f0fc, 32'hc303cb62},
  {32'h439b4654, 32'hc36c501a, 32'h43382697},
  {32'hc4a49bd5, 32'h4399797c, 32'h404eebbc},
  {32'h43e479e0, 32'hc32f99be, 32'h435ffe25},
  {32'hc4c5fc4f, 32'hc28e7ba8, 32'h43923dd2},
  {32'h4503339e, 32'h42bc7b4a, 32'h42897156},
  {32'hc3f0324f, 32'hc4009a62, 32'hc29739f1},
  {32'h44bfd75e, 32'hc1930be4, 32'h43a382a0},
  {32'hc3229e00, 32'h43012a23, 32'hc35c4cf8},
  {32'h43cee390, 32'hc3747a68, 32'h439e1e2a},
  {32'hc4a575ba, 32'h42c7fc48, 32'hc39a01a1},
  {32'h45130455, 32'h431c98f0, 32'h431dbfd6},
  {32'hc38ce758, 32'hc3258661, 32'hc4342274},
  {32'h4414009a, 32'h4229c718, 32'h43511e43},
  {32'hc4890336, 32'h41d29c06, 32'hc3309d1b},
  {32'h4440bb88, 32'hc2bde73b, 32'h4252cb10},
  {32'hc4f06c98, 32'hc30a6dd9, 32'hc3979ab0},
  {32'h44c591ce, 32'hc335b2ac, 32'hc2436ec7},
  {32'hc440f6b6, 32'hc3bbf794, 32'hc25e927b},
  {32'h4383770c, 32'h43df880f, 32'hc29823ab},
  {32'hc4c83b45, 32'hc392744f, 32'h40c6452c},
  {32'h44dd6c6c, 32'hc2f4392e, 32'h42981867},
  {32'hc451c02f, 32'hc332e213, 32'h4286d3e3},
  {32'hc4d8299b, 32'h4104f9ca, 32'h429e6817},
  {32'h44da1a5e, 32'hc354497c, 32'h43e90cf2},
  {32'hc4beadf7, 32'hc3624378, 32'h4304de54},
  {32'h44d50c96, 32'hc380b0e4, 32'h423fa3b5},
  {32'hc4d602cc, 32'hc28b9ca4, 32'h409f43e6},
  {32'h448bb104, 32'h42adbc8b, 32'h4442c4fa},
  {32'hc4bb6be3, 32'hc33091a8, 32'hc312fc44},
  {32'h449f3a4f, 32'hc2d6f5c7, 32'hc3876fd1},
  {32'hc51ae8ff, 32'h4279a7ae, 32'hc38dffac},
  {32'h45003c48, 32'h43ae5fe9, 32'hc320356d},
  {32'hc44e76d6, 32'h427ab648, 32'hc2d26d68},
  {32'h444aef78, 32'hc29124e0, 32'h4387d0f8},
  {32'hc4d2ba04, 32'h42218247, 32'hc2ba70bb},
  {32'h451514fc, 32'hc3e84ded, 32'h43dbbcb7},
  {32'hc4b1391e, 32'hc05787e4, 32'hc2880d9c},
  {32'h42acc904, 32'h4305932c, 32'h42f52a4d},
  {32'hc3e6cdd8, 32'h42c5453d, 32'hc389a177},
  {32'h44057414, 32'h426928f6, 32'h43b250b6},
  {32'hc4ca1d49, 32'h4405c39d, 32'h42438cf0},
  {32'h43f9a95c, 32'hc3792168, 32'h43aa3b7f},
  {32'hc2c150f0, 32'h4311db16, 32'hc36ba8ee},
  {32'h438956f3, 32'h43ea930a, 32'hc19d9585},
  {32'hc2cfab40, 32'hc3697380, 32'hc22b6348},
  {32'h449c901f, 32'h43318851, 32'h43411a96},
  {32'hc4c0b0be, 32'hc3814a46, 32'hc36dfeb4},
  {32'h44ca646b, 32'h422d2abc, 32'h42fe84bd},
  {32'hc4c99ea2, 32'hc3ab3b00, 32'hc3496a1d},
  {32'h4505bec9, 32'h430c11a2, 32'h41e0c0df},
  {32'hc3866537, 32'h431d66ee, 32'h42d4206d},
  {32'h44568a7e, 32'hc293be59, 32'hc34c466c},
  {32'hc4c631de, 32'hc38b11bc, 32'h43334b99},
  {32'h44fd33ef, 32'hc31b9a67, 32'h42ece0c7},
  {32'hc4cbf0b0, 32'hc21998da, 32'hc33e4738},
  {32'h44d14a6f, 32'h4280c969, 32'h43be5eb1},
  {32'hc4166d30, 32'h42feb9f4, 32'hc3b816bf},
  {32'h450d2b74, 32'hc1a9b5f5, 32'hc2b9e784},
  {32'hc4540b30, 32'h426e65cc, 32'h42fba01a},
  {32'h43583928, 32'hc31a2731, 32'hc2c961a6},
  {32'hc4c0dd65, 32'hc3a5e1bb, 32'h4318e19f},
  {32'h430a8b08, 32'h42cc4acf, 32'h43a62d0f},
  {32'hc46519d8, 32'hc351b38d, 32'h41c0b415},
  {32'h433d482e, 32'h413aa15b, 32'h433bdfb0},
  {32'h43e87d90, 32'h429a724b, 32'h4212b54e},
  {32'hc2af1c60, 32'hc3f4a4ee, 32'h4303d481},
  {32'hc4c3254d, 32'h4386dd22, 32'h436b89ff},
  {32'h450000e0, 32'hc3580ebf, 32'h42d9dcd6},
  {32'hc514cf24, 32'hc3112406, 32'h41837474},
  {32'h44f65d00, 32'hc3cf037e, 32'h440083da},
  {32'hc4345668, 32'hc2717dc2, 32'hc0b74998},
  {32'h446fee7e, 32'h42ac03c1, 32'h4276783e},
  {32'h42e17139, 32'h42f906b9, 32'hc3e0b03d},
  {32'h44d41569, 32'h425e1c7a, 32'h4360a88c},
  {32'hc38e1378, 32'hc2dbe3fa, 32'h427e1eb0},
  {32'h44e2ded5, 32'hc373d7b2, 32'h41f22dbc},
  {32'hc36547e8, 32'h4332e15a, 32'h41543eb2},
  {32'h446476f4, 32'h41cabd3f, 32'h4203eedf},
  {32'hc4216a10, 32'h43448633, 32'h4322aa01},
  {32'hc2ed4d90, 32'hc336d435, 32'hc26fb823},
  {32'hc3ece8a8, 32'h4330a2d0, 32'hc36a5740},
  {32'h450a840c, 32'h43bb5ab5, 32'h42e3f62f},
  {32'hc370e998, 32'hc411aec5, 32'hc312efba},
  {32'h42c395d0, 32'h42bf857e, 32'hc2e1c463},
  {32'hc42c8f58, 32'h41c39510, 32'h429a68d4},
  {32'h44c892df, 32'hc2d554c2, 32'h41d90e4a},
  {32'hc38a9860, 32'h4294d23c, 32'hc32f34da},
  {32'h43d26c40, 32'h420a64a3, 32'hc325dd0b},
  {32'hc500c555, 32'hc316f587, 32'h4314aee0},
  {32'h4339c72b, 32'hc2114f14, 32'hc312767a},
  {32'hc4c41083, 32'h410a8b92, 32'hc2c25505},
  {32'h41432c00, 32'hc190b4fd, 32'h433f44f8},
  {32'hc4048f4e, 32'h43bd5c69, 32'h43c0a404},
  {32'h4255af10, 32'hc3dffa6a, 32'hc2b2e44a},
  {32'hc41b5938, 32'h43a5c7a6, 32'hc3ff80aa},
  {32'h44ba02f7, 32'h43382b01, 32'hc396ee28},
  {32'hc49a8c86, 32'hc39d660c, 32'h431a51b6},
  {32'h42acc500, 32'hc198d3ba, 32'h436ac7e8},
  {32'hc4872dd0, 32'hc2a045cc, 32'hc3ab9f25},
  {32'h42cecf40, 32'h42aecfb6, 32'h431e60f5},
  {32'hc4f665ae, 32'hc2fd8cb3, 32'h43657875},
  {32'h44bcbf2c, 32'h421d5f86, 32'hc1b31b3c},
  {32'hc4fe6576, 32'h434c1729, 32'h42e3a56e},
  {32'hc35ec5cc, 32'h422315f9, 32'h438f4e3d},
  {32'hc3f5c368, 32'hc3c4b78b, 32'h4398d6a3},
  {32'h42804a00, 32'h4317a910, 32'hc324b859},
  {32'hc46a69af, 32'h42ffb520, 32'hc28be751},
  {32'h446759ce, 32'h42ae5068, 32'hc26a5beb},
  {32'hc4906089, 32'h43893cd1, 32'hc3bd20d6},
  {32'h44e5f4d4, 32'h43646895, 32'hc3639992},
  {32'hc4bbbd00, 32'hc3ed42fe, 32'h43a27be2},
  {32'h443a2e7f, 32'h42d85b68, 32'h43b03341},
  {32'hc4da9290, 32'hc38061e6, 32'h42bdd34b},
  {32'h41f03908, 32'hc30204a9, 32'h434199b8},
  {32'hc49c9751, 32'hc3548e2e, 32'h43c10a07},
  {32'h44859452, 32'hc3ac31a6, 32'hc1e6b261},
  {32'hc404c98e, 32'hc24b0011, 32'hc21d27f8},
  {32'h43ce82c8, 32'h42a4a6d1, 32'h42ba809b},
  {32'hc48de501, 32'hc2d84405, 32'h421ac175},
  {32'h44909d1d, 32'hc3121394, 32'hc311c17c},
  {32'hc2f3b9d0, 32'hc38d4ab4, 32'h42513cdd},
  {32'h44e70fd4, 32'h43199fa8, 32'h441bfe27},
  {32'hc4fb2b7c, 32'h4344fdbc, 32'h4415065f},
  {32'h43340920, 32'h43a6d043, 32'hc223c775},
  {32'hc4b40e34, 32'hc31be183, 32'hc3288888},
  {32'h4483946a, 32'hc2b5700e, 32'hc3349ea2},
  {32'hc4be2899, 32'hc24677eb, 32'h42c36e80},
  {32'h44b3b40d, 32'hc1860452, 32'hc310fa0a},
  {32'hc4811dd5, 32'hc214923e, 32'h43dad067},
  {32'h44de9fd3, 32'hc34e9dbc, 32'hc1dee8d4},
  {32'hc50653ef, 32'hc36edd39, 32'h426eb5b2},
  {32'h44f247ec, 32'h4381edd0, 32'hc3c299dc},
  {32'hc483da03, 32'hc239ca1d, 32'h436b14af},
  {32'h44b7f4ec, 32'h43bc563e, 32'h42ac14f8},
  {32'hc4fdb5c6, 32'hc406e3ac, 32'h42978f8e},
  {32'hc298e71c, 32'hc3d0b4b3, 32'h435cf997},
  {32'hc4d2c67e, 32'h43c31c8e, 32'h4352e561},
  {32'h451742af, 32'h42ffd72e, 32'hc3bf6c41},
  {32'hc3e73f5c, 32'h4315f5b6, 32'h43c0d26c},
  {32'h451102f2, 32'hc39ed0b3, 32'h42d14a31},
  {32'hc514de8d, 32'h43c7da7c, 32'hc2561eda},
  {32'h45069efc, 32'hc2e17d93, 32'h43546abf},
  {32'hc502778e, 32'h4332cc74, 32'h431e51ec},
  {32'h43938da5, 32'h42b3d80b, 32'h43c3e063},
  {32'hc50199f2, 32'hc2a4f6f8, 32'h4380c404},
  {32'h44870dd0, 32'h40f4585a, 32'h43a155a4},
  {32'hc485189d, 32'hc35f6867, 32'h43b639a4},
  {32'hc0c7ca80, 32'h439f3739, 32'hc34ecf33},
  {32'hc4004378, 32'h415a5a88, 32'h431d8868},
  {32'h44414492, 32'h43053b27, 32'hc2d4e6da},
  {32'hc49d8183, 32'h43a0ea0d, 32'h43a28162},
  {32'h4427b4b0, 32'h430cb452, 32'h42f84553},
  {32'hc4cd221e, 32'hc3203d1c, 32'h42c08d96},
  {32'h43cfc5f8, 32'h43111563, 32'hc36d8ecc},
  {32'hc42076c8, 32'h40d42400, 32'h42e74943},
  {32'h44316062, 32'hc34e84eb, 32'h438ebee5},
  {32'h43317090, 32'h431b0aff, 32'h42ffb434},
  {32'h43aadcaf, 32'h43161c53, 32'hbf1f6f84},
  {32'hc3cae888, 32'h438deed4, 32'h43c525d1},
  {32'h448de9c9, 32'hc36384b9, 32'hc3c367e8},
  {32'hc494559c, 32'h4376a261, 32'h42c8504b},
  {32'h44e842c1, 32'h43d3611a, 32'hc1b4cd6f},
  {32'hc3789e90, 32'hc284f148, 32'h4347a0bf},
  {32'h44e76caf, 32'h43482a5a, 32'h4380744a},
  {32'hc479f054, 32'hc33298a7, 32'h41ecf6d9},
  {32'h44ac3906, 32'h4314d369, 32'hc25c450a},
  {32'hc387bfc8, 32'h428aacaf, 32'hc29b5be4},
  {32'h44e3cafa, 32'h418de951, 32'h42460468},
  {32'hc4fd8c69, 32'hc3a19a40, 32'hc231cb03},
  {32'h44075bbc, 32'hc151ed54, 32'h432635ff},
  {32'hc3de6d8e, 32'h41a8ad67, 32'h438da0dc},
  {32'hc2d11f5a, 32'h43a8a827, 32'hc39747b4},
  {32'hc50195fa, 32'hc2d8c627, 32'hc35ae55c},
  {32'h442d7a16, 32'h436e295c, 32'hc3496665},
  {32'hc4e1ee72, 32'hc399d656, 32'h435ecdbb},
  {32'h44543742, 32'hc1ba0dbc, 32'h4302b844},
  {32'hc5080f67, 32'hc34d9323, 32'h42a12b16},
  {32'h44e9ee2e, 32'hc34d989f, 32'h418a9c57},
  {32'hc4b46a89, 32'hc313d6e8, 32'hc3027855},
  {32'h4517bdc0, 32'hc1980d61, 32'hc3dca49a},
  {32'hc4ca368e, 32'h4373ab4b, 32'hc09514ca},
  {32'h44d8cef6, 32'hc1677082, 32'h41632666},
  {32'hc3e9b360, 32'h42c7055b, 32'h43bb7e2b},
  {32'h42c6efc0, 32'hc35a1239, 32'hc2f6cae1},
  {32'hc445f730, 32'hc3972185, 32'hc20fe0f9},
  {32'h446f80d2, 32'hc3b2e513, 32'h428caabf},
  {32'hc474efb4, 32'h43abce61, 32'hc407fd50},
  {32'h43a4e308, 32'h4393ff76, 32'hc3b8551b},
  {32'hc3a5e0ac, 32'h42c28679, 32'h438c3662},
  {32'h45019c22, 32'hc1ee4eaa, 32'h3ea89808},
  {32'hc5014035, 32'h431e6ce1, 32'hc2f3e87f},
  {32'h433be471, 32'h4385f740, 32'h4320a390},
  {32'hc3957510, 32'h4329e1fb, 32'hc3821b38},
  {32'h44ff51a5, 32'hc2969c53, 32'hc38418d6},
  {32'hc4c0154e, 32'hc22b080c, 32'h438fcee4},
  {32'h446721ac, 32'h43adcb47, 32'h41a90e8a},
  {32'hc4b95535, 32'h42936b10, 32'h427dcf96},
  {32'h44a87cc0, 32'hc3238ca7, 32'hc247a8d7},
  {32'hc3f75062, 32'h43a1c008, 32'h43b9459e},
  {32'h451133a8, 32'hc25c988c, 32'h43896c9d},
  {32'hc504e624, 32'h434b6a38, 32'h4191c16b},
  {32'h4463f370, 32'hc1d50464, 32'hc40ac1f4},
  {32'hc50065ca, 32'hc27c7273, 32'hc2846a3e},
  {32'h4473c5ee, 32'hc3c7e47d, 32'hc34d144d},
  {32'hc4dceedf, 32'h4378eb52, 32'h41b275ab},
  {32'h44879785, 32'h42ac9b1b, 32'h4335e54c},
  {32'hc4d1dc0a, 32'h413c91d2, 32'h42a4597b},
  {32'h43a22d78, 32'h417a5784, 32'hc24d40fa},
  {32'hc478678b, 32'h42063b23, 32'h421ff139},
  {32'h440d1eb2, 32'h43b6a01e, 32'h41dcc925},
  {32'hc420ffba, 32'h42d975ab, 32'hc2c7d36d},
  {32'h4462d818, 32'hc39362be, 32'h42bcff89},
  {32'hc3422430, 32'h42956eff, 32'h4292c71f},
  {32'h4412a422, 32'hc1c3eec3, 32'hc37d9351},
  {32'hc36cfe40, 32'hc3ad6813, 32'h4290da11},
  {32'h41ac2880, 32'h434b5534, 32'hc0584ea7},
  {32'hc4e2263b, 32'hc11a81a1, 32'h43503aec},
  {32'h449c81e8, 32'h42007348, 32'h4404adb9},
  {32'hc393ce98, 32'hc311b581, 32'h427c1dda},
  {32'hc29018d0, 32'h4171c672, 32'h42b8beca},
  {32'hc3e43934, 32'hc3c12fab, 32'hc3f7962b},
  {32'h450c7bd3, 32'hc3732751, 32'hc21b4cc2},
  {32'hc4a9752f, 32'h436ea79e, 32'hc3c98c3c},
  {32'h44871de0, 32'h4370a285, 32'h431b880c},
  {32'hc4eba89e, 32'hc3161012, 32'hc1ba1468},
  {32'h439a4a50, 32'h42f2749c, 32'hc3805c00},
  {32'hc2e12ae0, 32'h42929a1e, 32'hc29194e7},
  {32'h43b10da4, 32'h43295f61, 32'h4288fee2},
  {32'hc4bf9e61, 32'h43aa9f14, 32'hc3628f14},
  {32'h43bad969, 32'h425b861e, 32'hc2ccedb0},
  {32'hc502ee32, 32'hc311b73c, 32'hc3abe8ca},
  {32'h4493a42e, 32'hc2960c5d, 32'hc33fb322},
  {32'hc3b55838, 32'h43cab661, 32'hc304e010},
  {32'h4514888c, 32'h434e20c1, 32'hc3892e62},
  {32'h42d3234a, 32'hc25f44a4, 32'hc3258a57},
  {32'h45154b9d, 32'h44020632, 32'hc2c80265},
  {32'h43a6f09f, 32'h429efc4f, 32'h42987ae3},
  {32'h449f67de, 32'hc32418ca, 32'h4158096e},
  {32'hc40ddafc, 32'hc2703193, 32'hc2badf2e},
  {32'h43b0d79c, 32'h41fe844f, 32'h43b3de90},
  {32'hc26042a0, 32'hc1722bd5, 32'h42429e45},
  {32'h44b2c302, 32'hc2cd79b4, 32'h42b15f96},
  {32'hc49d7a19, 32'hc38d791a, 32'hc2ba4117},
  {32'h441f3eb4, 32'h4325e617, 32'hc31e99d0},
  {32'hc400d4af, 32'hc414ddab, 32'hc1b0ca97},
  {32'h4427beb0, 32'hc324b59c, 32'hc19d8864},
  {32'hc484a3f9, 32'h43963075, 32'h426f72a1},
  {32'h44c8f528, 32'h435e450d, 32'hc34cfe3c},
  {32'hc24018b8, 32'h437454a6, 32'h41a52697},
  {32'h44315808, 32'h43767dac, 32'hc36a9b85},
  {32'hc40e5d0b, 32'hc36f02e3, 32'h427ee523},
  {32'h44bcbc32, 32'h420120ad, 32'hc1fefb10},
  {32'hc3a7ef0c, 32'h42a17a92, 32'h42f8057f},
  {32'h44bd81ab, 32'hc302c08e, 32'hc36ce9f1},
  {32'hc425abab, 32'h41c3eb3b, 32'h432cde44},
  {32'h44735480, 32'hc18538cf, 32'hc2ed1cd4},
  {32'hc5134c21, 32'h41c9e589, 32'h434aaf7d},
  {32'h448b494c, 32'h42f51809, 32'h41cbdcc4},
  {32'hc44fd3c3, 32'h41e84204, 32'hc35e7d7b},
  {32'h449ce6cb, 32'h42eb295c, 32'h41910267},
  {32'hc506b991, 32'hc3310401, 32'h40a0f08d},
  {32'h4423a673, 32'hc399868d, 32'hc288b3ae},
  {32'hc4ab4564, 32'h4363a2a7, 32'h437bf88a},
  {32'h44a37c23, 32'hc2b42532, 32'hc3302b9c},
  {32'hc41f74e8, 32'hc2efd3a8, 32'hc3845e57},
  {32'h44c472d2, 32'h4327a325, 32'h431dd418},
  {32'hc3d51db6, 32'h438ac487, 32'hc2e1ed69},
  {32'h44cfaf9d, 32'hc2a3f28c, 32'hc39f65fd},
  {32'hc4f97ad4, 32'hc2a98744, 32'h43aa7905},
  {32'h44a78424, 32'hc30c2087, 32'h41942014},
  {32'hc47e109c, 32'h429108c7, 32'hc2c90d8c},
  {32'h449a81f1, 32'h4231d862, 32'hc39fdea1},
  {32'hc514b963, 32'hc3842437, 32'hc24ecea7},
  {32'h4265bd00, 32'hc35d68e5, 32'hc2c87a9a},
  {32'hc3f435c8, 32'hc333c856, 32'hc367bdb6},
  {32'h451e6e39, 32'hc30b2a34, 32'h43294212},
  {32'hc506c014, 32'h439ead49, 32'hc2cf390b},
  {32'h441eff2b, 32'hc1e82cc0, 32'hc0b7dd79},
  {32'hc4b975da, 32'hc338b95b, 32'hc3222fbb},
  {32'h444e7afe, 32'h4317ae2e, 32'hc1b5ff78},
  {32'hc48aa6cb, 32'hc0738da2, 32'h42763fb0},
  {32'h44bde58c, 32'h4304e7e5, 32'hc2c24b5e},
  {32'hc51d7500, 32'h428720fe, 32'hc3a94d6c},
  {32'h450df726, 32'h4308daf7, 32'h42afec49},
  {32'hc50a7a5b, 32'h42a2d455, 32'h434448bd},
  {32'h446600a6, 32'hc3823928, 32'h43a7f4ab},
  {32'hc4f7c374, 32'hc33dbae8, 32'hc38267d9},
  {32'h44edbab3, 32'h43565691, 32'h42dbc6ea},
  {32'hc4e97990, 32'hc3754660, 32'hc2d46eb3},
  {32'h44d88a20, 32'hc35ba0b7, 32'h41902b0f},
  {32'hc4c70988, 32'hc21ddb07, 32'hc36719b1},
  {32'h4520e3b8, 32'h42928dc9, 32'h4365dc3c},
  {32'hc4b58e5d, 32'h42f35cd3, 32'h43ad1b07},
  {32'h446c27b2, 32'h432c4755, 32'h42819275},
  {32'hc4c488b8, 32'h42407190, 32'h43911b2f},
  {32'h44c92f78, 32'hc20d1c31, 32'hc341a8fb},
  {32'hc42587da, 32'hc42d0271, 32'hc3bb3394},
  {32'h449dcf7d, 32'hc240607b, 32'hc340df55},
  {32'hc29f0600, 32'h433d2f3a, 32'h41bcf1f7},
  {32'h443ddf9a, 32'h42cb1800, 32'hc1c1732c},
  {32'h4229fd20, 32'h41b62a5b, 32'hc3ded945},
  {32'h42e80e77, 32'h43870bee, 32'h43f8ec4a},
  {32'hc4d6d745, 32'h43c4597e, 32'hc3b4977a},
  {32'h444ddf54, 32'hc0cbfd2a, 32'hc263d7ea},
  {32'h41d5c580, 32'h42ba4cf3, 32'hc3e13aa4},
  {32'h44323284, 32'hc3a5962a, 32'hc30b2114},
  {32'hc3d42870, 32'h43431e96, 32'h3fb46898},
  {32'h43a80a60, 32'hc2a08d6f, 32'h4363741e},
  {32'hc48731d6, 32'h43a5fb73, 32'h432eed2c},
  {32'h44f63519, 32'h42ceaf02, 32'h40de1590},
  {32'hc4fd8115, 32'hc2b0e13b, 32'h42c42937},
  {32'h4491d1d0, 32'h439e5fcc, 32'h43005ce5},
  {32'hc3a634d8, 32'h43406247, 32'hc31c13b6},
  {32'h4508440d, 32'hc318871f, 32'hc27cf93d},
  {32'hc5050119, 32'hc2d5c18a, 32'hc2dc9069},
  {32'h448e1ef7, 32'h43df0cce, 32'h4350ab80},
  {32'h42f8387c, 32'hc17aca35, 32'h419771cb},
  {32'h4470a9f2, 32'h41b73e9a, 32'hc2099dcc},
  {32'hc4fc5a3a, 32'hc29cc32d, 32'hc2bca04a},
  {32'h448cdfb1, 32'h42bb8aed, 32'h412d6496},
  {32'hc4dbefcb, 32'h42b2cedd, 32'hc1afd6b5},
  {32'h44e28388, 32'hc31ec8b6, 32'h43989137},
  {32'hc509d563, 32'hc108e740, 32'hc3a01f1e},
  {32'h450f43d1, 32'hc2a23e12, 32'hc3df217c},
  {32'hc1b21900, 32'hc3afa09b, 32'hc24ef7e5},
  {32'h448f7a74, 32'hc3196b14, 32'hc2a6ab2d},
  {32'hc386d42e, 32'hc26635f2, 32'h423d692f},
  {32'h44ecaec0, 32'h4353f63b, 32'hc2cad7e7},
  {32'hc47bef9c, 32'h427f61ec, 32'hc316ee1b},
  {32'h4413501e, 32'hc1b1cdb9, 32'hc389f626},
  {32'hc4718229, 32'hc30471d1, 32'h440a052e},
  {32'h44a74807, 32'hc2b4ee5e, 32'h42007e36},
  {32'hc49cf399, 32'hc2e19faf, 32'hc35c2cd4},
  {32'h44c42aa9, 32'h43232ece, 32'h42b15d2b},
  {32'hc4462cb0, 32'hc341add1, 32'hc19f9e06},
  {32'h44958e64, 32'hc2ba0dc2, 32'h4330f654},
  {32'hc4226644, 32'hc35f40a0, 32'h3f88f080},
  {32'h44f9a795, 32'h42f40fa1, 32'h3fea80f4},
  {32'hc4745444, 32'h43190568, 32'h42caf4bb},
  {32'h44fc664c, 32'hc354ce0f, 32'h4347cf99},
  {32'hc501f2a4, 32'h438ca9a2, 32'hc3754db1},
  {32'h44b169ec, 32'h42e319ec, 32'h4320d418},
  {32'hc47d4269, 32'h43290fea, 32'hc38a7f32},
  {32'h44e83641, 32'h43f0a93e, 32'hc2e743c5},
  {32'hc408d1d4, 32'h4384fbda, 32'hc2955b45},
  {32'h44deba71, 32'hc3f25ca5, 32'hc2d5578f},
  {32'hc43613b4, 32'hc3a1730d, 32'hc30f725e},
  {32'h44135010, 32'h429f322e, 32'h43fdf1e0},
  {32'hc4c88305, 32'hc4121f0e, 32'h4290457e},
  {32'h445a4b10, 32'hc2391a0e, 32'h42b22f7c},
  {32'hc3297001, 32'h41f5cef0, 32'h43d38558},
  {32'h44d472e0, 32'hc0addbcb, 32'hc28d355b},
  {32'hc42bc1f8, 32'hc3979e55, 32'hc338da54},
  {32'h450eac66, 32'hc32cbfca, 32'hc3bf970b},
  {32'hc5015829, 32'h435367aa, 32'h430240c7},
  {32'h45132344, 32'h41d34c7c, 32'hc394fce0},
  {32'hc41b6014, 32'h42ed8e30, 32'hc37a5647},
  {32'h42b534a0, 32'h43a5b905, 32'hc39c0464},
  {32'hc524b62e, 32'h433246e5, 32'h4323e59a},
  {32'h448146b8, 32'hc1f94ffd, 32'h42d9b9ed},
  {32'hc46a55d2, 32'hc3224ce7, 32'h42b06ce0},
  {32'h44a98b23, 32'h43bdcee4, 32'h4370f654},
  {32'hc45f99d1, 32'h4347dc22, 32'hc37b657d},
  {32'h44c71ed0, 32'h4355e6ed, 32'hc39eeb08},
  {32'hc4bd6c05, 32'h42ccf774, 32'h4130d334},
  {32'hc20c01c4, 32'h4221f16f, 32'hc2b3e329},
  {32'h41475080, 32'h427dc621, 32'h42751baf},
  {32'h44d28c26, 32'hc2f08fde, 32'hc30942b6},
  {32'hc3cbb177, 32'hc351eccf, 32'h42d4104a},
  {32'h435599b8, 32'h4347a7da, 32'hc33f9bc8},
  {32'hc49c302e, 32'hc39c8522, 32'hc08388de},
  {32'h44eddff6, 32'h43478880, 32'hc2700d0b},
  {32'hc5128c54, 32'hc3bc0b09, 32'h43d540e0},
  {32'h446d9a08, 32'hc2d0be50, 32'hc2a63325},
  {32'hc4c21780, 32'hc3da580e, 32'hc217204e},
  {32'h43cd6f78, 32'h437141e3, 32'hc223591c},
  {32'hc4930d56, 32'hc3a4b0fc, 32'hc363fa5a},
  {32'h45161967, 32'hc3e9c17f, 32'h4347c02c},
  {32'hc48b5cf2, 32'h4327fd62, 32'h42ab1e63},
  {32'h43f7d966, 32'h4402bd67, 32'hc39ea3cf},
  {32'hc4e91d3b, 32'h43b2ba85, 32'hc30f8de7},
  {32'h43140d88, 32'h4232ebbe, 32'h43bfad32},
  {32'hc3da9650, 32'hc35fb5d3, 32'hc3706670},
  {32'hc2c8de10, 32'h427b03a6, 32'hc279e8f3},
  {32'hc4ad8fdd, 32'hc37962b2, 32'h420763f8},
  {32'h42906cc0, 32'h42924441, 32'hc299178e},
  {32'hc3e2020e, 32'h436ae9e8, 32'h429cc089},
  {32'h45013daa, 32'hc135c854, 32'h42552eaa},
  {32'hc40297c2, 32'h435ff2d6, 32'h438b4afc},
  {32'h44d1756e, 32'h433398ee, 32'h435596f8},
  {32'hc410df3c, 32'h43909ba8, 32'h43c0aae9},
  {32'h45030b9f, 32'h42598e86, 32'h4274fe38},
  {32'hc389c4d0, 32'hc34b8aa8, 32'hc3a2fded},
  {32'h44ffe81c, 32'hc2615cc5, 32'h4338790e},
  {32'hc3c722b1, 32'h428a9312, 32'hc2f404d6},
  {32'h44486725, 32'hc368aa61, 32'hc3aa5939},
  {32'hc51a0721, 32'h43a3bf10, 32'hc293c8ad},
  {32'h453090b8, 32'h43af1307, 32'hc2356790},
  {32'hc4a4615e, 32'h41ec4b14, 32'h435e16f3},
  {32'h4447488d, 32'h41d8f1b5, 32'hc20e1178},
  {32'hc4245dc2, 32'hc38a8bb7, 32'hc2baa7d5},
  {32'h44ec9be4, 32'h43439c94, 32'h43801d4a},
  {32'hc2dc7880, 32'h43253550, 32'hc3f30cc5},
  {32'h449279e6, 32'h429a5351, 32'hc219add7},
  {32'h422ef81e, 32'hc4146538, 32'hc2dccafe},
  {32'h44e104aa, 32'hc2ac5b71, 32'hc30824f9},
  {32'hc5189389, 32'hc35f8de0, 32'hc376ca8a},
  {32'h452e34ed, 32'hc30a9400, 32'h43d8136c},
  {32'hc5074ec4, 32'hc3c3d828, 32'h41e6efb0},
  {32'h44c822aa, 32'h42010a72, 32'hc21a9d08},
  {32'hc437cb7f, 32'hc3905a0e, 32'h43bfe55d},
  {32'h4296a450, 32'h438f9486, 32'hc36c7206},
  {32'hc4a9ce19, 32'hc355ffcf, 32'hc3009d06},
  {32'h449edc2b, 32'h4378b99f, 32'hc3cc1af5},
  {32'hc4c424ee, 32'hc30570b5, 32'h43b25368},
  {32'h44d3b033, 32'h436a6e08, 32'h425c1d6c},
  {32'hc485ff3d, 32'h42942895, 32'hc2c32d29},
  {32'h43d85e44, 32'hc31d8403, 32'h420ad2b5},
  {32'hc4921780, 32'hc31e4aec, 32'hc0c2eeb9},
  {32'h442c47ec, 32'hbf052b26, 32'hc38caa0b},
  {32'hc4aa2b23, 32'h42d104b4, 32'h42b379fe},
  {32'h44240e30, 32'hc2f97477, 32'hc2e893a1},
  {32'hc4470ae3, 32'h42302902, 32'hc221b72e},
  {32'hc2b75b10, 32'h42860c34, 32'hc378386d},
  {32'hc5037870, 32'hc2a5a952, 32'hc36bd484},
  {32'hc14c0200, 32'h43a02b3b, 32'hc289033e},
  {32'hc4bf887d, 32'h435cd1e1, 32'h43e9a79c},
  {32'h45086cc9, 32'h43aa1fcf, 32'hc2581c3d},
  {32'hc4353342, 32'h428fb632, 32'h420237f6},
  {32'h43ed06b0, 32'hc380e606, 32'hc398a595},
  {32'hc4360ef7, 32'hc0592314, 32'h43d4d3f7},
  {32'h44044c2a, 32'h4304d90b, 32'hc25c2f4a},
  {32'hc3fdb4f0, 32'h41dc08cc, 32'h41d1dfc7},
  {32'h42230010, 32'hc2287c20, 32'hc3c59b31},
  {32'hc5051076, 32'hc402bb7c, 32'hc388be1f},
  {32'h44b3b53d, 32'h428c2d12, 32'hc3666fda},
  {32'hc4d9bdec, 32'h43c1fb5b, 32'h43455a15},
  {32'h4489a0b2, 32'h438147dc, 32'h4243d944},
  {32'hc4cee63a, 32'hc21f65f6, 32'h434116c8},
  {32'h45138eba, 32'h42def2e4, 32'hc3ebd603},
  {32'hc4f43e53, 32'h438c0c20, 32'h4229881a},
  {32'h4429cc9c, 32'hc2c48638, 32'hc3dcee55},
  {32'hc42c8920, 32'hc330589a, 32'h4304b1af},
  {32'h438639f8, 32'hc2d0ab45, 32'hc2f64a1d},
  {32'hc5094c13, 32'h43850ab7, 32'h438e19d4},
  {32'h44cf093d, 32'h425158d5, 32'hc357a7d1},
  {32'hc50c5c52, 32'hc245abaa, 32'h429877d3},
  {32'h4508eaf2, 32'h438ac077, 32'hc2e8bec9},
  {32'hc4f1b953, 32'hc25f0609, 32'hc3081d04},
  {32'h444becd6, 32'h439af572, 32'hc28bd4f3},
  {32'hc39219d0, 32'hc2ccc590, 32'h432a1fa8},
  {32'h44c282d7, 32'hc3467016, 32'h43389dbe},
  {32'hc46960f6, 32'h42bb4046, 32'h43b155d7},
  {32'h44dfbda6, 32'hc30c0ca7, 32'hc32d7bd8},
  {32'h44fb4c0e, 32'h4339828f, 32'hc2ac050a},
  {32'hc4bf001a, 32'h43afcce7, 32'hc1f68e6d},
  {32'h44ccbaa4, 32'h42db11ee, 32'hc356eaaa},
  {32'hc4a0660b, 32'hc28f2c0e, 32'h42cb3cf6},
  {32'h44399bda, 32'hc387703b, 32'hc2383318},
  {32'hc4938d28, 32'h4399d321, 32'hc2b7bed1},
  {32'h43c72028, 32'hc364d2f9, 32'h4391bb07},
  {32'hc4cef2d4, 32'hc2efe04e, 32'h424b8b20},
  {32'h450e23c0, 32'h433503f9, 32'hc2bd7c18},
  {32'hc4ad0d82, 32'hc3308fb7, 32'h438fec84},
  {32'h449458ca, 32'hc3399b97, 32'hc346fe7f},
  {32'hc4aded9c, 32'hc305c5b8, 32'hc3748fcf},
  {32'h43eecd60, 32'hc229d2af, 32'h43d990cf},
  {32'hc4b8f2e3, 32'hc18405b6, 32'hc3d89dcb},
  {32'h44502526, 32'hc37adbb2, 32'hc3c666b2},
  {32'hc32e07a4, 32'hc23e75d6, 32'hc1eaf6c7},
  {32'h45018e3d, 32'h4376cd10, 32'hc1abddcb},
  {32'hc40855c0, 32'hc29c4201, 32'h4395a119},
  {32'h4405c68c, 32'hc30c0a8f, 32'hc2053813},
  {32'hc4f3ea7d, 32'h42858c12, 32'hc2ac02dd},
  {32'h4502face, 32'h438e919c, 32'h41e0782a},
  {32'hc4af83e8, 32'h41b82247, 32'h422b8226},
  {32'h42b8b8c4, 32'hc2877251, 32'h42913f5b},
  {32'hc4faa9fe, 32'hc217c130, 32'hc30cd176},
  {32'h45160700, 32'h43bda010, 32'h434fb0a7},
  {32'hc4cb464c, 32'h43b4452f, 32'hbfdb9970},
  {32'hc2fd6b4e, 32'h435a975c, 32'h42adcdcf},
  {32'hc4bac174, 32'hc2b9da87, 32'h42a65738},
  {32'h441a0218, 32'hc2fceaf4, 32'hc3b8c7e8},
  {32'hc4403be0, 32'hc393995c, 32'hc37eb90f},
  {32'h44d7cff5, 32'hc305f89f, 32'hc3620f76},
  {32'hc42526b0, 32'hc20d929c, 32'hc28745e9},
  {32'h43ec899e, 32'hc2cd3f3d, 32'h426507d4},
  {32'hc4dd6a6e, 32'h43147dc7, 32'hc340df4e},
  {32'hc2f8e718, 32'h41b77472, 32'hc3450592},
  {32'hc4876996, 32'hc2dc7b45, 32'hc21264f6},
  {32'h41614780, 32'hc3a57814, 32'hc3e594d5},
  {32'hc4bc40ee, 32'h42aa9ccc, 32'h435f6002},
  {32'h44e6f2a3, 32'hc3550476, 32'h4368fc2c},
  {32'hc4e66583, 32'h437fa228, 32'hc39ad783},
  {32'h4458d4c6, 32'hc3b02a73, 32'hc3809567},
  {32'hc3bd2c80, 32'hc26b7332, 32'hc20fbb23},
  {32'h443e5f14, 32'h41e1dcd4, 32'h433292a3},
  {32'hc40b4e40, 32'hc385bc8d, 32'h43881e89},
  {32'h450f8dcb, 32'hc23cf6e7, 32'hc24f62a9},
  {32'hc433a1dd, 32'hc3827a95, 32'hc3e50856},
  {32'h4511957e, 32'hc33eb4a0, 32'h42422b7b},
  {32'hc3467b3e, 32'h43d0f290, 32'h4357ef33},
  {32'h44c70779, 32'h4259bd7c, 32'hc3848b8d},
  {32'hc3ee18c8, 32'hc2d3191f, 32'h434a2e32},
  {32'h441f8082, 32'hc2ca257b, 32'h42b4a5a2},
  {32'hc4a32928, 32'hc34ad53a, 32'h437639e9},
  {32'h44fb415e, 32'hc378127b, 32'h43addb3b},
  {32'hc4bec153, 32'h430d6966, 32'h414fa75c},
  {32'h451a4f83, 32'h4181b7a1, 32'hc3d7069e},
  {32'hc41281b7, 32'hc3bb4be8, 32'hc399e6b1},
  {32'h441f65c0, 32'h42ae8ef6, 32'hc20a7e66},
  {32'hc507928e, 32'h42ab808a, 32'hc3b7256c},
  {32'h44ef42b3, 32'hc42f170b, 32'hc3961f48},
  {32'hc501be42, 32'hc30b89e0, 32'hc3124770},
  {32'h44d00fc5, 32'hc2e234b4, 32'hc38608c0},
  {32'hc42dc66a, 32'h44061bfa, 32'h438bab89},
  {32'h4409338a, 32'h41d730fc, 32'hc2e2f44c},
  {32'hc41d5e1e, 32'hc3a40d64, 32'hc24b70e8},
  {32'h45058e95, 32'hc39b8474, 32'hc32a3dc0},
  {32'hc519647f, 32'hc35c8c06, 32'hc1d00864},
  {32'h447557af, 32'h41fdfa44, 32'hc371ee90},
  {32'hc4eceadf, 32'hc232efeb, 32'hc401eb94},
  {32'h44554199, 32'h42907a1e, 32'h3f8ea4b8},
  {32'hc4f8af98, 32'hc36af9f0, 32'h433c85f5},
  {32'h451ae456, 32'hc313f20c, 32'h437c75fc},
  {32'hc3f57ba5, 32'h42a0422b, 32'hc30708de},
  {32'h43f98cbd, 32'hc3da978c, 32'hc09f5b21},
  {32'hc49c7f71, 32'h414146e8, 32'h43a38620},
  {32'h45210894, 32'hc329e298, 32'h43473b2a},
  {32'hc4b9fad4, 32'h41f5ce87, 32'h436d6121},
  {32'h43aa29c4, 32'hc407bb85, 32'hc32fac5b},
  {32'hc41eaece, 32'hc2d45bb2, 32'hc29cb705},
  {32'h44ad1214, 32'hc36afe53, 32'h430db44e},
  {32'hc4886226, 32'hc325eb7a, 32'hc24119ba},
  {32'h44b35566, 32'hc3db218a, 32'h43822c8e},
  {32'hc437b4ec, 32'hc2c6e810, 32'h43bacd06},
  {32'h450ad9a1, 32'h42d6509a, 32'hc24acb34},
  {32'hc3fdb7d0, 32'h42ab79fe, 32'h42ad7630},
  {32'h44fde952, 32'hc3bc4c85, 32'h43fffeab},
  {32'hc28f2a70, 32'hc31ad067, 32'h4181f7b4},
  {32'h44f6ba17, 32'h4301aa8f, 32'hc352f58a},
  {32'hc4a7f874, 32'hc386b3fc, 32'h4283694d},
  {32'h449f9339, 32'hc3185cd6, 32'h41c0df6f},
  {32'hc4b703c6, 32'hc377ceb5, 32'h431a0f6e},
  {32'h451807d5, 32'h4148759b, 32'hc3a2ad34},
  {32'hc4c4b8ef, 32'h44036c4e, 32'h43504cc7},
  {32'h444db5d0, 32'h43d7078a, 32'h40c853bc},
  {32'hc39ca2ce, 32'hc2b4d57c, 32'hc3b4cc3c},
  {32'h442ed1ec, 32'h437f1d3b, 32'hc32314a2},
  {32'hc4501375, 32'hc3ace46e, 32'h4294fc2b},
  {32'h4509d2b1, 32'h42119fcc, 32'hc25efc3a},
  {32'hc4dda802, 32'hc2fab10c, 32'h40ff1b20},
  {32'h45065558, 32'hc1e21bcd, 32'hc2b608a5},
  {32'h425619c0, 32'hc2ade8c0, 32'h43df84fa},
  {32'h451a029b, 32'h440be71f, 32'h42f39e60},
  {32'hc501610f, 32'hc394e51e, 32'h439103b1},
  {32'h4483c92a, 32'hc314cf46, 32'h4380fe80},
  {32'hc487714a, 32'hc3425d7f, 32'h430222d6},
  {32'h4480ec5e, 32'h43b37a80, 32'h4326f409},
  {32'hc2e3f762, 32'h42914935, 32'hc2234868},
  {32'h44ba7b3a, 32'hc2014c25, 32'hc219c1c5},
  {32'hc4dd8dd6, 32'h4314218d, 32'h41939a9a},
  {32'h4446f1de, 32'h42c78941, 32'hc348b8ac},
  {32'hc500dbb6, 32'h436e70d5, 32'hc33a238d},
  {32'h43faed98, 32'hc383a73c, 32'hc3edf545},
  {32'hc4b5b884, 32'hc309837d, 32'hc337d148},
  {32'h4384b65a, 32'hc4239785, 32'h429eafc9},
  {32'hc491b0ae, 32'hc33a8bd4, 32'h4342752c},
  {32'h447d5c3e, 32'hc300170d, 32'h4400448d},
  {32'hc4846634, 32'h422f446a, 32'hc1da7e72},
  {32'h45191191, 32'hc3b28662, 32'h42e3064f},
  {32'hc4f4b616, 32'hc3bbff35, 32'h431f07fd},
  {32'h44a2f81c, 32'h42d1d1e9, 32'h421265c4},
  {32'hc4bee527, 32'hc3510e2b, 32'h43c42fd7},
  {32'h429413a8, 32'hc144aa73, 32'h4378a673},
  {32'hc51f5bf2, 32'h432763b9, 32'h4287b3d2},
  {32'h44869846, 32'hc2ceb541, 32'h43721632},
  {32'hc4a3a0b2, 32'hc408a410, 32'h421b9ddf},
  {32'h4409fdd1, 32'hc2f60b15, 32'h4365aff4},
  {32'hc4bc84dd, 32'hc283c38a, 32'hc1983255},
  {32'h437c3d00, 32'h42f7a53c, 32'h42891f65},
  {32'hc50c2bbc, 32'hc3244dd7, 32'h4331bade},
  {32'h4493d0d6, 32'hc3111a0a, 32'h4284cad4},
  {32'hc466ae16, 32'h436a7379, 32'h4331ba06},
  {32'h44f0b415, 32'h437f3695, 32'h43c58363},
  {32'hc5067761, 32'hc3ab9db8, 32'hc3215b54},
  {32'h43177824, 32'h43ad23be, 32'h436e17df},
  {32'hc3910e2a, 32'h434d2d49, 32'hc2cf7fb9},
  {32'h4491fbc1, 32'hc30bfa92, 32'hc2d040cb},
  {32'hc5019d4a, 32'h41c15bab, 32'hc2d54557},
  {32'h441c2811, 32'h437e59d3, 32'h438c021e},
  {32'hc3d82b48, 32'hc3c12956, 32'h4287ff26},
  {32'h44f58427, 32'hc2e272cb, 32'hc35e53ba},
  {32'hc406e3fa, 32'h42069ba8, 32'h42bc9f1a},
  {32'h445df640, 32'h42e916d2, 32'h42d07348},
  {32'hc4da8ba6, 32'hc3cd5601, 32'hc33ae24a},
  {32'h44d1b56b, 32'hc40abee4, 32'h434a0308},
  {32'hc3a89e40, 32'h43940ce5, 32'hc3103052},
  {32'h43c02a24, 32'hc2b81674, 32'h43411256},
  {32'hc4186073, 32'h42445351, 32'h431b5ba2},
  {32'h45003cc0, 32'hc3339fc0, 32'h43cbb8bf},
  {32'hc38e647e, 32'h42b1c77a, 32'h43a009d4},
  {32'h44d8f4e2, 32'h436ba18e, 32'hc12d9e0a},
  {32'hc0af3000, 32'hc34fce79, 32'hc3a656e7},
  {32'h44b6b304, 32'h43dd57ac, 32'h4391e928},
  {32'hc5042470, 32'hc33fe16a, 32'hc3a66bd1},
  {32'h44ce1332, 32'hc3f95fac, 32'hc2a18872},
  {32'hc5021425, 32'hc206fe3c, 32'hc3de7aaa},
  {32'h44f3435d, 32'h4283e50a, 32'h42fecd19},
  {32'hc3c6b729, 32'h431d40e5, 32'hc359b1d4},
  {32'h450bf040, 32'hc2d27701, 32'hc02ece6d},
  {32'h431b0498, 32'hc359bb7a, 32'hc362cc58},
  {32'h4411b59a, 32'h42834656, 32'hc29ead61},
  {32'hc41a3867, 32'hc38c1567, 32'h43ac9fd9},
  {32'h44cda9c4, 32'hc38893f4, 32'h436efa1f},
  {32'hc4a242b2, 32'hc2eac90f, 32'hc19939e8},
  {32'hc355daa8, 32'hc33634a5, 32'hc32215bd},
  {32'hc5148206, 32'hc3ab37fa, 32'h42942cdd},
  {32'h43cca504, 32'hc3c241bd, 32'hc4179ae8},
  {32'hc30b4738, 32'hc304a228, 32'h42f346b6},
  {32'h44ec86a9, 32'hc1f52c68, 32'hc2423308},
  {32'hc3de1290, 32'hc3c1017c, 32'hc260588d},
  {32'h4422135e, 32'h43cded74, 32'h431a9363},
  {32'hc407aa1a, 32'h43047264, 32'h438dddad},
  {32'h44e6db58, 32'h42e878ee, 32'hc2fbccd3},
  {32'hc4a546e3, 32'h43a22f23, 32'hc30fa379},
  {32'h44e60322, 32'hc357e8e7, 32'h416cd6ca},
  {32'hc4f1ea77, 32'hc2f521b2, 32'hc386f423},
  {32'h44ba8b14, 32'h433c1647, 32'hc2bd20a2},
  {32'hc4643e8f, 32'hc2849063, 32'h4389eed7},
  {32'h43e3e012, 32'h42842260, 32'h42e8f340},
  {32'hc4cf9a85, 32'hc19ba128, 32'h43bcb2c0},
  {32'hc3205b32, 32'hc3169f85, 32'h436e2074},
  {32'hc4e5eea6, 32'h4318d8ee, 32'hc2e1c79b},
  {32'h415d955c, 32'hc38dcdaf, 32'h426c774c},
  {32'hc5046451, 32'h4258c284, 32'hc326b3e8},
  {32'h44fe5cd7, 32'hc2f97024, 32'hc332cc08},
  {32'hc4dfbb68, 32'h43a3a8a7, 32'hc3ac3d50},
  {32'h446d4b56, 32'hc3395b70, 32'h42833998},
  {32'hc49bde63, 32'h42f94ee1, 32'h439602ee},
  {32'h44790e0a, 32'h42a29903, 32'hc365b302},
  {32'hc4bb6234, 32'h42b98383, 32'hc3e184bc},
  {32'h4486526c, 32'h435bc6d9, 32'hc26d348a},
  {32'hc4fccb4f, 32'h43334140, 32'hc1ff9e77},
  {32'h4428c79d, 32'h4377d064, 32'h437f77ba},
  {32'hc4d927fc, 32'h433b518e, 32'hc391ec14},
  {32'h44ef9d1e, 32'h42cf9e3f, 32'hc315c778},
  {32'hc3f65c06, 32'hc334b02c, 32'hc2da37d4},
  {32'h448a70a4, 32'hc3115661, 32'h438e354e},
  {32'hc3a03fb0, 32'h418c7315, 32'h42edfe2b},
  {32'h44663418, 32'hc32800d2, 32'hc331d988},
  {32'h40946d94, 32'h42ffc285, 32'hc276d050},
  {32'h44be7034, 32'h42ad1690, 32'h42b01f99},
  {32'hc264d800, 32'hc379ae87, 32'hc36503df},
  {32'h44331032, 32'h42370e7c, 32'h42c97ec7},
  {32'hc4b180d6, 32'hc333fd1f, 32'h43039d6c},
  {32'h43cf51f0, 32'hc31899d1, 32'hc2d3ba2c},
  {32'h42cbbbbf, 32'hc3618e60, 32'hc38334ee},
  {32'h44849c14, 32'h4347ad50, 32'hc31cb1ab},
  {32'hc483fb5c, 32'hc268db11, 32'hc2adc461},
  {32'h44de89bb, 32'hc400523a, 32'hc2beb63c},
  {32'hc4aca88b, 32'hc33c848b, 32'hc3abce63},
  {32'h450c84ee, 32'hc399c343, 32'h42c37c72},
  {32'hc4002a52, 32'hc3822c34, 32'hc29f122a},
  {32'h44e1eca6, 32'h423521e8, 32'h434413ad},
  {32'hc4be41b4, 32'h41548774, 32'hc139311a},
  {32'h443b4249, 32'h43573e49, 32'hc367beee},
  {32'hc34f5370, 32'hc3e70bc3, 32'hc36b770b},
  {32'h4511c3a4, 32'h43b26442, 32'hc3c10365},
  {32'hc4ff4f0f, 32'h40208a17, 32'h436d9e1d},
  {32'h44568a93, 32'hc32745d3, 32'hc138ee76},
  {32'hc40250fc, 32'hc1099592, 32'h43586c78},
  {32'h448e3de1, 32'hc153a5be, 32'h429a7f2d},
  {32'hc4ee8fb8, 32'h41e124ca, 32'hc348619d},
  {32'h450a3593, 32'hc2fd7b4e, 32'h41259435},
  {32'hc3d4835b, 32'h4089d9c8, 32'h438e9849},
  {32'h44142c93, 32'hc31cd769, 32'hc1ab15ab},
  {32'hc4c23ac0, 32'hc27b7413, 32'h4343b7c2},
  {32'h445961d2, 32'hc27eebd7, 32'hc3374ab0},
  {32'hc4af2c70, 32'hc291c0d7, 32'hc352ac63},
  {32'h4456ec43, 32'h439e97ed, 32'hc342002d},
  {32'hc40d1b84, 32'hc38a525e, 32'h42910af2},
  {32'h44855892, 32'hc2e491ce, 32'h435cebb5},
  {32'hc2e18c50, 32'h426bdeb8, 32'h42f232f0},
  {32'h44a4d768, 32'h43e45d31, 32'h426423fa},
  {32'h43026de4, 32'hc2e7385c, 32'hc2c500aa},
  {32'h451c254d, 32'h4322c9f4, 32'h4351fabc},
  {32'hc49793fc, 32'hc349ed32, 32'h43273ba9},
  {32'h44e25617, 32'h436aeb98, 32'h435985f5},
  {32'hc4645642, 32'h42df6e4e, 32'hc29b9ea8},
  {32'h44449540, 32'hc2416672, 32'h43c20cf8},
  {32'hc4d4c184, 32'h4192c719, 32'hc323bec3},
  {32'hc1b78920, 32'hc34b5da1, 32'hc368a16b},
  {32'hc4cfd977, 32'h43b716b4, 32'h42a49fdf},
  {32'h44f45bc4, 32'hc2ce1b87, 32'hc29229fc},
  {32'hc4a494a6, 32'hc30ff669, 32'h4209349a},
  {32'h4447af1c, 32'hc4297be7, 32'h42fe5414},
  {32'hc505047d, 32'h43bedc94, 32'hc3841cf2},
  {32'h443b2474, 32'h43515250, 32'hc1308570},
  {32'hc4e38857, 32'h4284af5f, 32'hc28bcfd4},
  {32'h44bab22e, 32'hc06a2918, 32'h42c177da},
  {32'hc4143f7d, 32'hc2eb0b84, 32'hc374744a},
  {32'h437157f8, 32'h43510f4d, 32'h428131b0},
  {32'hc3249a40, 32'h432a6433, 32'hc2deece1},
  {32'h450d2981, 32'h4369f868, 32'h42df1949},
  {32'hc313dd8c, 32'hc30b19cd, 32'h4387cf32},
  {32'h4454b028, 32'hc3053914, 32'h430751f2},
  {32'hc485dd1e, 32'hc29eae92, 32'hc2db1542},
  {32'h44898446, 32'hc1fb801f, 32'h43634310},
  {32'hc24fff00, 32'h440d7ffc, 32'h42c21bab},
  {32'h44e95f2f, 32'h432ac1fa, 32'hc2e1bbe7},
  {32'hc4f1b32e, 32'h4069891c, 32'h4384e818},
  {32'h443f95d8, 32'hc38004f9, 32'hc385c33b},
  {32'hc47b842d, 32'hc1c47f24, 32'hc138f0c0},
  {32'h444695f0, 32'h4401cb3b, 32'h434e77a2},
  {32'hc4de4f61, 32'h43c0c504, 32'h42d6dae7},
  {32'hc28a0904, 32'h43497dc7, 32'h4361e428},
  {32'hc48fba22, 32'hc3b42810, 32'h4319e5f4},
  {32'h44067856, 32'h4425c1a6, 32'hc45c8dbb},
  {32'hc40c77e3, 32'h43750787, 32'h43dc5b5c},
  {32'h44578e00, 32'h4392dee4, 32'hc39d62e7},
  {32'hc48efa37, 32'h4339e901, 32'hc32c50eb},
  {32'h430756e0, 32'hc31b540d, 32'h42724c08},
  {32'hc4fc5ee9, 32'hc32af96d, 32'hc348faa1},
  {32'h4444267c, 32'h44007623, 32'h423d51e4},
  {32'h3fad1800, 32'h43bbc6d4, 32'hc1c0eed8},
  {32'h43b285df, 32'hc218afd4, 32'hc39327c4},
  {32'hc50a221f, 32'h42c0e931, 32'hc2ae2260},
  {32'h44e637f5, 32'hc2b1fad5, 32'hc36a08b3},
  {32'hc449cfb0, 32'h433c7812, 32'hc30bac29},
  {32'h44bebe23, 32'h428d90f7, 32'h42346f89},
  {32'hc5108330, 32'hc2f86d40, 32'hc330b347},
  {32'h443b2ae8, 32'hc1e0d7f1, 32'h43ab96a7},
  {32'hc2f5be22, 32'hc25e67e7, 32'h43813fb8},
  {32'h43739b40, 32'h4393a0eb, 32'h432428d4},
  {32'hc3802d27, 32'h42c76271, 32'hc3137494},
  {32'h4426dd14, 32'hc3cac6be, 32'hc25eaaf8},
  {32'hc3fdef56, 32'h43b419f6, 32'hc336ac0a},
  {32'h44aeeacc, 32'h431c9c0e, 32'hc19d643e},
  {32'hc4a6439b, 32'hc365f291, 32'hc326e11f},
  {32'h44849f60, 32'hc05954da, 32'hc2d86882},
  {32'hc4670e44, 32'hc2d15150, 32'hc3964d1a},
  {32'h42e72350, 32'hc3d0b56d, 32'h4354da4c},
  {32'hc43caa00, 32'h43e341a7, 32'hc340e7d3},
  {32'h4491a45b, 32'h41b52f72, 32'hc1722969},
  {32'hc36ff6f0, 32'h427e1c48, 32'h43ff31e0},
  {32'h4500bd67, 32'hc39c2cc8, 32'h4317d369},
  {32'hc4ebf3f3, 32'hc1d09b39, 32'hc1f32792},
  {32'h44c51445, 32'hc372982e, 32'hc27e2b39},
  {32'hc4bc5cc8, 32'hc2b8bb58, 32'h42cfd015},
  {32'h449e6c26, 32'hc2219535, 32'h433c8661},
  {32'hc5002044, 32'h42e1d1e2, 32'h426564f8},
  {32'h43981aa8, 32'hc373ea92, 32'h418f0964},
  {32'hc50972ec, 32'hc3b788f5, 32'h4347efc6},
  {32'h44821070, 32'h434512f8, 32'h4190987e},
  {32'hc2e2aed0, 32'h43dde093, 32'hc3e3a8a7},
  {32'h4515b124, 32'h43252f04, 32'hc3bbca5e},
  {32'hc46939ae, 32'h42b0f833, 32'h412a780e},
  {32'h43777f8c, 32'hc36fdd55, 32'hc366896f},
  {32'hc4f40f88, 32'h41827c32, 32'h431e80dd},
  {32'h44a3be22, 32'h4407a684, 32'h415c519b},
  {32'hc444bcc8, 32'h4346242e, 32'h434bc960},
  {32'h4438a3b8, 32'h439219d3, 32'hc39c22b8},
  {32'hc4b8b265, 32'h41734c17, 32'hc2bd4591},
  {32'h445a2c0a, 32'hc36cba3b, 32'hc34879a0},
  {32'hc4f70d9b, 32'hc0b29190, 32'h433e7238},
  {32'h448d4e3b, 32'hc375d847, 32'hc36e2a3d},
  {32'hc3ca68ae, 32'hc31feccd, 32'h4316a70a},
  {32'h43b7b006, 32'hc3227382, 32'hc1af6de9},
  {32'hc485f7b6, 32'h437c95b5, 32'h42e2eae5},
  {32'h426a8f80, 32'hc302830a, 32'h42f6e929},
  {32'hc32bbb52, 32'hc2d0085c, 32'h438cefcd},
  {32'h450f4c77, 32'h42b55079, 32'hc281f245},
  {32'h416777a2, 32'hc3fa5856, 32'h4342a034},
  {32'h450807f2, 32'h428dcee2, 32'hc42a2d59},
  {32'hc468dcd2, 32'h43fc3a43, 32'hc2992124},
  {32'h450d9c82, 32'h426f8e5b, 32'h43b4da96},
  {32'hc461500e, 32'hc3972ae5, 32'h42812b2f},
  {32'h4415e757, 32'h43654baa, 32'h41af5b4d},
  {32'hc22b76a0, 32'h42064ca8, 32'hc35c5a22},
  {32'h43855581, 32'hc35d80b9, 32'h426721de},
  {32'hc4e0a5de, 32'h43176910, 32'h434556be},
  {32'h450f5083, 32'hc3a0874a, 32'hc2f96225},
  {32'hc5017cb2, 32'h4221dfa9, 32'hc222aadf},
  {32'h44b863d4, 32'hc36ee684, 32'hc3904738},
  {32'h43099d30, 32'hc3117721, 32'hc2301ca2},
  {32'h44d46c0a, 32'hc20a3b72, 32'hc2c2d3da},
  {32'hc519a2ad, 32'hc1d54900, 32'hc2f77cba},
  {32'h4497f402, 32'hc24a0cb2, 32'h43613105},
  {32'hc3cb3f06, 32'hc3c0d6b6, 32'h439eca75},
  {32'h44c5ac26, 32'hc3805d40, 32'hc3125242},
  {32'hc4dec27f, 32'h431dddd5, 32'hc30832c4},
  {32'h45114abd, 32'h42fe0060, 32'h421da82f},
  {32'hc4359e47, 32'hc2dff3fa, 32'h4354dea3},
  {32'h44a112ed, 32'h41905398, 32'h4117c348},
  {32'hc4e4ef37, 32'h432d3161, 32'h4241b944},
  {32'h450e4606, 32'h442f5a47, 32'hc3425164},
  {32'hc48dc5bc, 32'hc290b0ca, 32'hc39d20ae},
  {32'h45072a52, 32'h43866bc8, 32'hc414e049},
  {32'hc490de51, 32'h43807001, 32'h421435f5},
  {32'h44758cd9, 32'h435eeec9, 32'hc320476a},
  {32'hc48844d3, 32'hc2f80963, 32'h4386f652},
  {32'h44e5d83a, 32'hc2cf1ba4, 32'hc38e6775},
  {32'hc50057d2, 32'hc36d0c59, 32'h43054411},
  {32'hc0ade100, 32'hc3926093, 32'h418e78fe},
  {32'hc4d573eb, 32'hc3196d20, 32'hc19b0cfa},
  {32'h435afb9a, 32'h41b7923c, 32'h431a0bdf},
  {32'hc4c7a966, 32'hc3858d79, 32'hc322bf3c},
  {32'h446219df, 32'hc4069a24, 32'h432c0573},
  {32'hc4f3a278, 32'hc2727d87, 32'hc329908b},
  {32'h442372ee, 32'h43297b9f, 32'h42ae1064},
  {32'hc237d2f0, 32'hc0c1ce64, 32'h42ddfbd1},
  {32'h44b88414, 32'hc2d1b76f, 32'hc3874b6a},
  {32'hc4e683b4, 32'h43477a40, 32'h433dedaf},
  {32'h44f95f69, 32'hbfb8ebd0, 32'h44058a18},
  {32'hc4bcd98b, 32'h425778ad, 32'hc21b90b0},
  {32'h44c1a658, 32'hc36497ad, 32'h43f0e297},
  {32'hc1384a00, 32'h42618490, 32'hc3d81104},
  {32'h44497ca5, 32'hc352b62a, 32'h3e8ddb23},
  {32'hc3367a90, 32'h42e7bc70, 32'h438a1540},
  {32'h446202f6, 32'hc296cf4d, 32'hc37d60ba},
  {32'hc49b5b20, 32'h43248814, 32'hc289a27a},
  {32'h449ea435, 32'h432c2306, 32'h438c994e},
  {32'hc4a18c8a, 32'h43a2d9de, 32'h4229b059},
  {32'h44807c32, 32'h4354fab2, 32'hc3691733},
  {32'hc407ae06, 32'hc20df009, 32'h428cf112},
  {32'h4508d74b, 32'hc2f86f72, 32'hc2a41091},
  {32'hc34d8eb0, 32'h432a9911, 32'h4362dab6},
  {32'h4474897a, 32'h42baffb2, 32'hc2af9cac},
  {32'hc5063f55, 32'hc05282b8, 32'hc2d9268c},
  {32'h44187299, 32'h43c552a4, 32'h42e4f725},
  {32'hc424a200, 32'hc3e6c86e, 32'hc2aab5b3},
  {32'h4391d3a0, 32'h414caa28, 32'h4412292a},
  {32'hc2d66a48, 32'h42ae19a1, 32'hc292ffa2},
  {32'h44c48485, 32'h43975cf0, 32'h430ad2ad},
  {32'hc5234e5a, 32'hc35f77be, 32'h4385a5de},
  {32'h43b660ac, 32'hc3116c30, 32'hc2ea1b8f},
  {32'hc48f4afc, 32'hc2727dd9, 32'hc321860a},
  {32'h44aef14d, 32'hc1feec39, 32'hc31b2f71},
  {32'hc4ddaed5, 32'hc215962a, 32'hc3683af5},
  {32'h448b6c0b, 32'h42a5ad96, 32'h42a442df},
  {32'hc45959bd, 32'hc380f476, 32'h437efb09},
  {32'h437619c8, 32'hc288ba92, 32'hc2ddcbbf},
  {32'hc523d89d, 32'hc3584f7c, 32'h429132e9},
  {32'h44e0e0d6, 32'h43e8add7, 32'hc1911dde},
  {32'hc4e8eaf1, 32'h438d39c1, 32'h4321a36c},
  {32'h44091051, 32'hc33e61f1, 32'hc28d4ee4},
  {32'hc2c704f0, 32'h429404f9, 32'hc09c8ab0},
  {32'h44caf549, 32'h4373ab35, 32'h433421d6},
  {32'hc41902a4, 32'h4402baec, 32'h4381830f},
  {32'h44fc4354, 32'hc4012921, 32'hc1b21906},
  {32'hc4e8eb1f, 32'h436e1ec2, 32'h4217cb6e},
  {32'h43c4ab50, 32'hc3a4de5e, 32'h43abf931},
  {32'hc4195f62, 32'hc3a8e2b2, 32'hc3a32054},
  {32'h439c8d08, 32'hc22d73f8, 32'hc248ada9},
  {32'hc4afe54d, 32'h4389fa45, 32'h423be732},
  {32'h43a2d7e8, 32'hc38cfe0c, 32'hc309db43},
  {32'hc4f4b9ce, 32'hc32bd1c0, 32'hc3ae0705},
  {32'h450a5391, 32'hc36f63e1, 32'h42bfb453},
  {32'hc4ef5de0, 32'h42e22859, 32'hc31e73a2},
  {32'h4499e7a2, 32'h4403d683, 32'hc2ed2f61},
  {32'h43554950, 32'h431b19f6, 32'hc39c44b7},
  {32'h44b5f5e4, 32'hc2ddf38b, 32'h4376e6ab},
  {32'hc4ff9908, 32'hc30b774a, 32'hc1abdb71},
  {32'h44838bcb, 32'hc2af8a1d, 32'h422b1d56},
  {32'hc4b5225c, 32'h438c533c, 32'h4256c289},
  {32'h44271b51, 32'h42bf39d8, 32'h43858e55},
  {32'hc433ae50, 32'h438024d7, 32'hc2b4dcee},
  {32'h43fa952d, 32'h438fd4d6, 32'h433b3553},
  {32'hc46385dd, 32'hc3be9aac, 32'hc300baa2},
  {32'h42c017b0, 32'h4293e5f6, 32'h43b25bbd},
  {32'hc4dbffd8, 32'hc313b495, 32'hc2b2d3cc},
  {32'h438839cf, 32'h43613f29, 32'h429f0eb0},
  {32'hc4925ff4, 32'hc18e96f3, 32'h41c5089d},
  {32'h443e8640, 32'h42638c21, 32'h43832822},
  {32'hc2ec38f6, 32'hc2e482a5, 32'h40fd1ab3},
  {32'h44a134f1, 32'hc3b88a3f, 32'hc27d2901},
  {32'hc51a88bd, 32'h40d6ce20, 32'h420e32c6},
  {32'h44b06275, 32'h431fdea3, 32'hc3270c19},
  {32'hc344d670, 32'h4326ea62, 32'h43b7b171},
  {32'hbf4c9800, 32'h44162efe, 32'hc4054449},
  {32'hc4453aae, 32'h42113afa, 32'hc2aef302},
  {32'h44f0e38d, 32'h42198231, 32'h404fc6e8},
  {32'hc4d934aa, 32'h41a510bf, 32'h4358ea01},
  {32'h43d72553, 32'hc20bc6dc, 32'h436f09c5},
  {32'hc3654560, 32'h433e69e1, 32'hc37cc718},
  {32'hc4ad1548, 32'hc3c9c023, 32'hc3586a51},
  {32'h441e22da, 32'hc2dd6c8a, 32'hc2076bba},
  {32'hc4e3095f, 32'h42b7012e, 32'h434ac8ea},
  {32'h4444df0c, 32'h433cfbc9, 32'hc1481d18},
  {32'hc44c6178, 32'h428e9fa8, 32'h42bf2163},
  {32'h445b1054, 32'hc31d185f, 32'hc2adbd54},
  {32'hc346ba38, 32'hc3544c65, 32'hc3df39aa},
  {32'h4482c832, 32'hc30a368e, 32'hc2b334bc},
  {32'hc39a5be0, 32'h43939340, 32'h421b0fa7},
  {32'h43b7e282, 32'hc11aa27a, 32'hc38aeb2e},
  {32'h41e578e6, 32'hc346884e, 32'hc37b49a8},
  {32'h43f6d0b0, 32'h423c99db, 32'h436216ab},
  {32'hc4896606, 32'hc2461f9b, 32'hc3b9a329},
  {32'h447b2fe5, 32'h43d3c362, 32'hc31a6767},
  {32'hc45a2e5c, 32'h42b280be, 32'h4377a7dd},
  {32'h44c135c8, 32'h4290b70a, 32'hc192f780},
  {32'hc44f2229, 32'hc372a732, 32'h4344654c},
  {32'h44d7812a, 32'hc38f49a9, 32'h43c652ed},
  {32'hc4c78b4b, 32'hc2823616, 32'h42236d8b},
  {32'h447fdad7, 32'hc21d3278, 32'hc30dc1cc},
  {32'hc4ea6898, 32'h42d7026b, 32'hc2d1f355},
  {32'h44841d21, 32'h42b67fdb, 32'hc347d6ac},
  {32'hc480217c, 32'hc2012e1f, 32'hc3a8ab34},
  {32'h44ff3246, 32'h41ccc86c, 32'h42649f9a},
  {32'hc486ef23, 32'hc20ce193, 32'hc385823d},
  {32'h443c8f20, 32'h428b7ad8, 32'h40b10045},
  {32'hc30d6c60, 32'hc38feb4b, 32'hc20dc07b},
  {32'h4391f288, 32'hc3b5f7f8, 32'h432d5cdd},
  {32'hc4b3d7f1, 32'h4387b69d, 32'hc3bdbe53},
  {32'h44c06917, 32'h43b087c2, 32'hc1d2666b},
  {32'hc4d183dd, 32'hc1d00cbd, 32'hc3564172},
  {32'h440ef4a9, 32'hc3aa1a2d, 32'h422bc7a9},
  {32'hc4ed2fb7, 32'hc3a26290, 32'hc316a94f},
  {32'h4430dfae, 32'hc348531c, 32'h43b5c421},
  {32'hc4806405, 32'hc25373ca, 32'hc39ff272},
  {32'h44d04f2a, 32'hc34552dd, 32'h434467e6},
  {32'hc49cffad, 32'hc26ac9e2, 32'hc309b886},
  {32'h4430a62c, 32'hc2ae8b45, 32'h43f54c4d},
  {32'hc4af73c3, 32'h40f4266d, 32'h42dfe79a},
  {32'h440d4aea, 32'hc30ccf94, 32'hc3ac69ed},
  {32'hc39724d0, 32'hc2c3095c, 32'hc35d4ea6},
  {32'h43f460ec, 32'h43e8e764, 32'hc0e6d9c7},
  {32'hc4ebc09a, 32'h43403add, 32'h4395fe98},
  {32'h448dd568, 32'h422276c7, 32'h4377720f},
  {32'hc4f68bde, 32'hc1d23609, 32'hc3123c0e},
  {32'h44c5e1de, 32'h42a19dec, 32'h42e4568a},
  {32'hc4c896be, 32'hc3362305, 32'hc3321a6a},
  {32'h451d68ae, 32'hc309069e, 32'hc3104209},
  {32'hc4297e22, 32'h4180aadf, 32'hc2d2652a},
  {32'h447641e4, 32'hc3102e0c, 32'hc3a7b705},
  {32'hc4f49640, 32'hc3693d45, 32'hc3a8f79c},
  {32'h44a1e45f, 32'hc3092604, 32'hc2b0e644},
  {32'hc44e1492, 32'h437df669, 32'hc3e6678d},
  {32'h44d566af, 32'hc375bc45, 32'h4296b48c},
  {32'hc4fc0391, 32'h43651265, 32'h3f51d700},
  {32'h4503f57c, 32'hc24fdf17, 32'hc38b97f6},
  {32'hc472c8d5, 32'h43af0059, 32'h413a3b79},
  {32'h44f861f3, 32'h43d4f846, 32'hc3b1e3c6},
  {32'hc437a67a, 32'hc3a5e66c, 32'hc307efa4},
  {32'h445a9400, 32'hc190fd13, 32'h43013298},
  {32'hc4808385, 32'h42750432, 32'h415cacb9},
  {32'h44c975da, 32'hc3389951, 32'h43496e3c},
  {32'hc4d1333a, 32'hc324cad0, 32'hc36c44d6},
  {32'h45139272, 32'hc296fe50, 32'h4334db99},
  {32'hc43ce649, 32'h428f8f01, 32'h42b65f8d},
  {32'h44c6146d, 32'h43ef1f52, 32'hc324a960},
  {32'hc4350358, 32'hc28f2b20, 32'h43e9bd29},
  {32'h44627966, 32'hc34f4221, 32'hc418b316},
  {32'hc48853ff, 32'h43721f99, 32'h44029765},
  {32'h44f35ffd, 32'hc36a43a3, 32'hc3894b06},
  {32'hc3f5dbac, 32'h44129328, 32'h439eec72},
  {32'h4482255e, 32'hc3352403, 32'hc362d117},
  {32'hc4f2cd1f, 32'h42f69dbf, 32'h42839e28},
  {32'h44cc8d5a, 32'h43232bb4, 32'h412c8f37},
  {32'hc489c47d, 32'h43645baa, 32'hc400f3c4},
  {32'h43dc5940, 32'hc2264304, 32'h434e4ed7},
  {32'hc4fe4768, 32'h43d9b617, 32'hc302b13d},
  {32'h448d7b99, 32'hc177c0f6, 32'h42ec9a74},
  {32'hc4b71ac7, 32'h42dc84ad, 32'h4311d56d},
  {32'h45057ae6, 32'h431e7882, 32'h43d5f2e4},
  {32'hc490dc1e, 32'h4294a3c5, 32'h431aeba3},
  {32'h444df6d7, 32'h42e6b4cc, 32'h436520c4},
  {32'hc4ad7294, 32'h434308ee, 32'hc3f3ade1},
  {32'h44c9613d, 32'h42c407d5, 32'h43a28d31},
  {32'hc5193947, 32'hc209534a, 32'hc350e8da},
  {32'h440a729a, 32'h415edf33, 32'hc18de088},
  {32'hc4cc3b5e, 32'hc300c622, 32'h413db21b},
  {32'h44c0f5b0, 32'h428ebf18, 32'hc2b1ce74},
  {32'hc4ba94ac, 32'h431d1fc0, 32'h438dfad2},
  {32'h43bfa0f8, 32'hc32e2eda, 32'h4298cfbe},
  {32'hc3d68c22, 32'hc3c74074, 32'h435dab71},
  {32'h440cbc55, 32'hc37777d8, 32'hc2f8b361},
  {32'hc392db00, 32'h43a80c84, 32'h431728d9},
  {32'h44f7da9b, 32'h43315346, 32'h41a1955e},
  {32'hc4fb88e4, 32'h43a27bb4, 32'h43b5d5d1},
  {32'hc296307c, 32'h42976fcb, 32'h42841dd6},
  {32'hc4989532, 32'hc2c6bbf7, 32'h422c5536},
  {32'h450b4c79, 32'h43641ff2, 32'h430245fc},
  {32'hc398b828, 32'h42d2ebd0, 32'h43eaccc4},
  {32'hc3a8ac74, 32'hc280437c, 32'h42b54082},
  {32'hc3b40ef8, 32'hc3693ff4, 32'hc3ae8c1e},
  {32'h44b3fc92, 32'h41c0de9e, 32'hc34fe861},
  {32'hc391f5a4, 32'hc38996a0, 32'hc3accdad},
  {32'h450e3984, 32'hc320d354, 32'h43ce6145},
  {32'hc4f672e0, 32'h433574bc, 32'h43a59132},
  {32'h44d890c2, 32'hc1017c96, 32'hc30bd6a0},
  {32'hc4ce2110, 32'h43135ce2, 32'hc354aaf1},
  {32'h446c5ad4, 32'hc2bb106c, 32'h434459a4},
  {32'hc3e011e4, 32'h410a46a8, 32'h42a23e07},
  {32'hc2d3be60, 32'h42f95e8c, 32'hc3c30ebc},
  {32'hc4add0f7, 32'h44131db4, 32'h42318a90},
  {32'h43a500e8, 32'hc2b8da3b, 32'h420f21bd},
  {32'hc2af4920, 32'h42d55212, 32'h428b840c},
  {32'h44aa7b48, 32'h43896624, 32'hc2ed12ac},
  {32'hc413e7a4, 32'h425412c1, 32'hc3c6b45d},
  {32'h44d1fdf2, 32'hc2eb8cd0, 32'h4320464c},
  {32'hc40a4b0a, 32'h43b1b25a, 32'h41600d9b},
  {32'h430bf590, 32'h426a23bf, 32'hc2a37856},
  {32'hc434c0c8, 32'h435aed93, 32'h42ec8f66},
  {32'h44893d97, 32'h4359b97a, 32'h434d4164},
  {32'hc4acb5c9, 32'h42f11889, 32'h4387872a},
  {32'hc3379408, 32'h4334c6af, 32'h421a1660},
  {32'hc4f1501e, 32'h4215e8e9, 32'hc2b17409},
  {32'h44ba1f3e, 32'hc3011b8f, 32'hc288876c},
  {32'hc32a4758, 32'h432729e3, 32'h416a645f},
  {32'h44de67c6, 32'h41a93e92, 32'h4361e0c7},
  {32'hc4654305, 32'hc23d0c8d, 32'h432b5aa0},
  {32'h43cc8f92, 32'hc347ea85, 32'h431acbad},
  {32'hc3fe9ba8, 32'h4311938e, 32'h42525eab},
  {32'hc1e7ad20, 32'hc22edbe8, 32'hc3c351c4},
  {32'hc3c95f68, 32'hc3aeea20, 32'h42fa4385},
  {32'h440a5bef, 32'h434299cc, 32'h41ec69c7},
  {32'hc4fbcc9c, 32'hc290730e, 32'hc35482d4},
  {32'h44ff44fe, 32'hc080b1d8, 32'hc2ad7f68},
  {32'hc4af7596, 32'h42a0bf8d, 32'hc276dc2a},
  {32'h44ca887c, 32'hc3033cde, 32'hc20efa5d},
  {32'hc49be152, 32'h43017f6d, 32'h4341bd9e},
  {32'h43e156a0, 32'h420206ce, 32'hc3d3ee09},
  {32'h4375c321, 32'h43b3d327, 32'h43166d4c},
  {32'h45069c5e, 32'hc4335068, 32'h42a172bb},
  {32'hc4589666, 32'h423bf556, 32'h43adef38},
  {32'h4467612d, 32'hc39288fa, 32'hc2ca3d43},
  {32'hc4dac3a6, 32'h421418f1, 32'hc2745d87},
  {32'h451448ae, 32'h42940c6d, 32'hc2259c72},
  {32'hc50656ca, 32'hc209a550, 32'hc2aa26a3},
  {32'h4416ee7e, 32'h43784b97, 32'hc2c3ce9d},
  {32'hc4eaae57, 32'h42e836e6, 32'hc2261bf4},
  {32'h44eed1d6, 32'h42d99ebc, 32'hc36921e8},
  {32'hc3da1fd0, 32'h4429f5c0, 32'hc28831b8},
  {32'h4508cd82, 32'h42d7c2aa, 32'hc35d924a},
  {32'hc3b55061, 32'h438a1dd0, 32'h418b3d16},
  {32'h44dca60d, 32'hc2a75112, 32'h436e800f},
  {32'hc5031034, 32'hc3a0b325, 32'h43a1766e},
  {32'h44eda526, 32'h438499a3, 32'h42cc874c},
  {32'hc4c94018, 32'hc2b2bed0, 32'h42703187},
  {32'h450873f9, 32'h433a2611, 32'h43f9d52d},
  {32'hc48db4f4, 32'hc2122e2e, 32'h43181cde},
  {32'h4513f704, 32'hc4188824, 32'h437849a6},
  {32'hc442b06a, 32'hc363ec6a, 32'hc3273a6e},
  {32'h4507ca6f, 32'h430641d6, 32'hc332920c},
  {32'hc4ea7e1c, 32'hc3838f85, 32'hc374172c},
  {32'h4498535f, 32'hc3ad2ba5, 32'hc28d0f02},
  {32'hc4d7e367, 32'hc2c4bb7b, 32'hc369440d},
  {32'h432978e8, 32'h43207622, 32'hc3ddfd33},
  {32'hc42adb5c, 32'hc0b41e70, 32'h43b900b8},
  {32'h431b9110, 32'hc3a150e6, 32'h42d3b816},
  {32'hc3df34f4, 32'h418b07fb, 32'hc2fedc85},
  {32'h4411c221, 32'h43610a85, 32'hc3e64291},
  {32'hc40fe5c1, 32'hc383f2b4, 32'h435c281e},
  {32'h44a34c4a, 32'h437bfb8e, 32'h43ee3010},
  {32'h418ab980, 32'h4384b3f8, 32'h432997ca},
  {32'h44ce980a, 32'h438d6042, 32'hc35f9aa5},
  {32'hc4b98da4, 32'hc3f4e044, 32'h435ff048},
  {32'h448c473f, 32'hc30e78aa, 32'h438b3fdd},
  {32'hc4948ada, 32'h42afe224, 32'hc2b3edf9},
  {32'h44d76f79, 32'h43651ebe, 32'h434d57ff},
  {32'hc4e67716, 32'h43246c42, 32'hc3f08337},
  {32'h45165c05, 32'hc397cf30, 32'h43475053},
  {32'hc38b3b2a, 32'hc284cf82, 32'h438278ad},
  {32'h449a2b8d, 32'hc16253a2, 32'hc17a7e4b},
  {32'hc49dd443, 32'hc34fd992, 32'h423a0816},
  {32'h44be6400, 32'h43f22983, 32'h4367840e},
  {32'hc4db4655, 32'h428d663d, 32'h41cc56d7},
  {32'h44e064ba, 32'h4293083b, 32'hc28c27b7},
  {32'hc509155a, 32'hc288d5f9, 32'hc317bd41},
  {32'hc31c122c, 32'h430cb779, 32'h429d39aa},
  {32'hc514f9eb, 32'hc3248f76, 32'h428188b6},
  {32'h44c59b08, 32'h4230341f, 32'h41505749},
  {32'hc4619222, 32'hc2d89af0, 32'h4418ddbb},
  {32'h450cc34e, 32'hc3140f10, 32'h438906b3},
  {32'hc4185d28, 32'h43947805, 32'hc263bf2d},
  {32'h44c60574, 32'h43718681, 32'hc3a8add0},
  {32'hc482f49c, 32'h430d91f1, 32'hc31ab442},
  {32'h448a6fca, 32'h43c40bc4, 32'h434c6023},
  {32'hc41c5ea0, 32'hc2d7f788, 32'hc3987cee},
  {32'h449ffc22, 32'hc362ad8a, 32'hc3a666de},
  {32'hc2a14055, 32'h430fc909, 32'h438e073d},
  {32'h445414d8, 32'hc3394bc5, 32'h420823b9},
  {32'hc35bf950, 32'h42ef23ae, 32'h40a87850},
  {32'h440bf6c4, 32'h440007a4, 32'h41a017a7},
  {32'hc44b687d, 32'h42e3d7af, 32'hc3582cc3},
  {32'h44f0e85d, 32'h42e792e2, 32'h41737edb},
  {32'hc47063e4, 32'hc2dd8c25, 32'hc1490ff5},
  {32'h44bc8305, 32'h43765be4, 32'h43931da7},
  {32'hc4fad52a, 32'h43aa33ed, 32'h42c83eb9},
  {32'h4462cb53, 32'h43b53732, 32'hc31eb2d2},
  {32'hc45805b0, 32'h409bceb0, 32'h4344a29a},
  {32'h44c115bf, 32'h438d7c62, 32'h43e635fe},
  {32'hc2e268e0, 32'hc2b0b8ec, 32'hc3740041},
  {32'h450b821a, 32'hc1d85fd0, 32'hc0bff86a},
  {32'hc4ec43f0, 32'h4393cfed, 32'hc23def24},
  {32'h45118797, 32'hc3b6738e, 32'h43224da0},
  {32'hc4dc45d1, 32'hc26c800e, 32'hc2800de6},
  {32'h448b6320, 32'hc425a84a, 32'h43297329},
  {32'hc3171738, 32'h42d332b6, 32'h43ddc5f4},
  {32'h44aa4cea, 32'hc318d794, 32'hc2bc7932},
  {32'hc36eef18, 32'h428d7995, 32'h42af1990},
  {32'h44f52585, 32'h43658da9, 32'hc2c68929},
  {32'hc3e7f8d8, 32'h42e436d9, 32'h43952736},
  {32'h44b0ae24, 32'h420abd94, 32'hc2bab3f0},
  {32'hc435d30c, 32'h41b0975b, 32'hc1ddd16e},
  {32'h4487d35e, 32'hc42ce63c, 32'hc3a6c4d2},
  {32'hc3ce4e84, 32'h43b36fd7, 32'h428754a6},
  {32'h42691529, 32'h4349bc55, 32'h422157ce},
  {32'hc4d13bd8, 32'hc2783e61, 32'h42b52212},
  {32'h44cac793, 32'h43f862d5, 32'h417404a4},
  {32'hc424b1b5, 32'hc2ce459d, 32'h43c00411},
  {32'h44e89fa2, 32'h4337fd07, 32'hc2374e9b},
  {32'hc4b9c5b0, 32'h438837c8, 32'hc23f77cc},
  {32'h45110e68, 32'hc2d02fae, 32'h4317bca8},
  {32'hc4d521ec, 32'h43468941, 32'h43705916},
  {32'h450a2453, 32'h43ffa781, 32'hc20aede1},
  {32'hc36735e0, 32'h43cf7b1f, 32'h43a8db65},
  {32'h4494b672, 32'hc295633a, 32'h42749a91},
  {32'hc43bcc11, 32'hc182c56f, 32'hc3f03445},
  {32'h45072876, 32'hc3f73cdc, 32'h43b4d912},
  {32'hc4c6a59e, 32'h40d577f4, 32'hbda04c90},
  {32'h450fe174, 32'h43282a52, 32'hc2f931b4},
  {32'hc50095eb, 32'h438a14a7, 32'h3f62ebb8},
  {32'hc2d06dd0, 32'hc37c0774, 32'h43684b4d},
  {32'hc3e6e6b8, 32'h42695c41, 32'h42290280},
  {32'h44cb8728, 32'h42f815c4, 32'h42f33831},
  {32'hc4ed0fc8, 32'h4332f7f3, 32'hc260093b},
  {32'h44c4afdf, 32'hc2d9b840, 32'hc3120cd1},
  {32'hc465e530, 32'h427d1c86, 32'hc1f98a0b},
  {32'h43c8ce73, 32'hc34ed14d, 32'hc344a0f3},
  {32'hc4af24af, 32'h42427ba3, 32'h4089ffbd},
  {32'h4333f13c, 32'hc35ae951, 32'hc26de6ef},
  {32'hc50609c2, 32'h420cc1b5, 32'h430ba2a0},
  {32'h44e7bacf, 32'hc3d36bb3, 32'hc165b3a2},
  {32'hc4c03624, 32'h438c4c50, 32'hc34e1d26},
  {32'h44bdb148, 32'hc28c8e05, 32'hc202ff7b},
  {32'hc3b52870, 32'hc43f3f61, 32'h428b57c2},
  {32'h3ec10000, 32'h42b264b4, 32'h438d67e6},
  {32'hc45a28e8, 32'hc161b2c7, 32'hc369c2fb},
  {32'h43accd92, 32'h430fef7a, 32'hc2292db0},
  {32'hc3ddb234, 32'h43bfb6d8, 32'h43021360},
  {32'h44e67926, 32'hc2cfefd7, 32'h43101ec6},
  {32'hc4e5fcd6, 32'hc2b4c429, 32'hc3940280},
  {32'h44e85044, 32'h43909edb, 32'h43b7ea12},
  {32'hc4a62abb, 32'h43476c68, 32'h438a7197},
  {32'h44aaed6b, 32'hc301793e, 32'h43b3473b},
  {32'hc508ddcc, 32'h43544a57, 32'hc339caf9},
  {32'h44b479b7, 32'h42bd24ee, 32'h42864a0c},
  {32'hc4a14ad1, 32'hc33529fd, 32'h43dfe7a9},
  {32'h4506c0e6, 32'h4391add2, 32'hc3ef4f3f},
  {32'hc2601140, 32'hc3770c6d, 32'hc35362db},
  {32'h45166c72, 32'hc3565ad2, 32'h428fb101},
  {32'hc50a675e, 32'h425fb880, 32'hc3b36e43},
  {32'h4498cad9, 32'h42c67ee3, 32'hc37e8a18},
  {32'hc3fa6958, 32'hc07ba613, 32'h433dcb24},
  {32'h44fd278c, 32'hc3e3bcf4, 32'h43788ff7},
  {32'hc4073094, 32'hc2cfca45, 32'hc4263380},
  {32'h44952edb, 32'h433b613f, 32'hc31c8e69},
  {32'hc4d36dca, 32'h43bcff0a, 32'h42b46fa2},
  {32'h450d6ef2, 32'h4326d1f0, 32'h4171bfd4},
  {32'hc504648a, 32'hc32a4756, 32'h4388f039},
  {32'h446b5c34, 32'h42485282, 32'hc2c41896},
  {32'h42534930, 32'hc31afdde, 32'hc33c892d},
  {32'h4513af34, 32'hc301503f, 32'h42f61ccf},
  {32'hc4c6b3d0, 32'hc1bf1f63, 32'hc1d4a783},
  {32'h4504d75c, 32'hc3159e17, 32'hc20b7be0},
  {32'hc496e134, 32'h417a1501, 32'hc34211a2},
  {32'h44b57d90, 32'hc2f9c800, 32'h43865078},
  {32'hc3ab2a54, 32'h42f64239, 32'h42f7dc37},
  {32'h44dcc3a2, 32'h426f30fc, 32'h43c627b0},
  {32'hc3acf15c, 32'h4357564d, 32'h4394ad3c},
  {32'h449b9b4c, 32'hc399ec02, 32'hc26dd372},
  {32'hc4eab2bb, 32'h43062202, 32'hc30bb045},
  {32'h44b80910, 32'h440e3d82, 32'h42a2eb08},
  {32'hc4255404, 32'hc3b91aa6, 32'hc1c744d8},
  {32'h4481a9f7, 32'hc19caab3, 32'hc30d61f0},
  {32'hc4e93cfe, 32'hc2a75faf, 32'hc25785c5},
  {32'hc2d21a60, 32'h44183e99, 32'hc35b1b63},
  {32'hc4a1e3a4, 32'h43e99017, 32'hc28409ba},
  {32'h4491fca0, 32'h42a85b5b, 32'hc3cf721c},
  {32'hc514bd7c, 32'h4353ee8b, 32'h424f3b59},
  {32'h445a08a4, 32'h439c5b8c, 32'h420cd187},
  {32'hc4ffb670, 32'h431593d9, 32'h4408fd41},
  {32'h44fc510c, 32'hc201e753, 32'h416c8cbe},
  {32'hc397b329, 32'h428d3278, 32'hc2ee6b06},
  {32'h44976ad3, 32'hc3699f67, 32'hc348151c},
  {32'hc4c276c2, 32'hc1140655, 32'hc3fcd760},
  {32'h44cf943f, 32'h438ef5ef, 32'hc388d341},
  {32'hc50849e7, 32'hc3853fd3, 32'hc2cc8465},
  {32'h44619db8, 32'hc2b7007c, 32'h42a267ec},
  {32'hc44ade38, 32'hc331e787, 32'hc3975f19},
  {32'hc1166910, 32'h431dc1ea, 32'h43591c34},
  {32'hc507d1da, 32'hc31d3bcf, 32'h43d57c19},
  {32'h4429f002, 32'h4017af34, 32'hc2f17a3a},
  {32'hc417b6da, 32'hc38b0284, 32'h417030e4},
  {32'h43afda18, 32'h423d665d, 32'h41a40fd0},
  {32'hc4b5329d, 32'hc339f44a, 32'h430e25e2},
  {32'h43e7ebc4, 32'hc37f01fe, 32'h438f2baf},
  {32'hc50d0c55, 32'hc2845ad7, 32'h4322cd9b},
  {32'h43f98f40, 32'h43db11a0, 32'h43303d46},
  {32'hc468a051, 32'h422e8749, 32'hc24e97e8},
  {32'h43cab2b0, 32'h43676f1b, 32'hc31467ae},
  {32'hc3be9c20, 32'h4390cc02, 32'hc378f209},
  {32'h447044c9, 32'hc3386e18, 32'hc33f0929},
  {32'hc4d45de3, 32'h41cdfa9a, 32'hc331424e},
  {32'h445c2708, 32'hc3eac8c7, 32'h43bbb0cc},
  {32'hc51ed65c, 32'hc2a20977, 32'hc35b8fec},
  {32'h44165744, 32'hc2d632a9, 32'h42e37d81},
  {32'hc419e736, 32'hc29bf2de, 32'hc3b5271b},
  {32'h448abeb3, 32'h43ca32d9, 32'hc305d74f},
  {32'hc2bc8f90, 32'h414a0f20, 32'h4211e3df},
  {32'h451e2ec7, 32'h4315df3f, 32'h431e973e},
  {32'hc4d1cf4e, 32'h4049909f, 32'h42d86668},
  {32'h440fe56c, 32'h430493c2, 32'h42274053},
  {32'hc451e2b2, 32'hc362ce21, 32'h432adf2f},
  {32'h43d1a1e7, 32'hc28b9318, 32'h42467abe},
  {32'hc4db8c72, 32'h43279c52, 32'h433dac9a},
  {32'h449bd7c2, 32'hc391bc2a, 32'hc32a8cb4},
  {32'hc4951785, 32'hc350c273, 32'hc3890381},
  {32'h430bca00, 32'h40282980, 32'h44029966},
  {32'hc4967911, 32'h43f64b54, 32'hc40493cd},
  {32'h44c65826, 32'hc2ed5eac, 32'hc3148634},
  {32'hc3633e78, 32'hc2930f92, 32'h4351d938},
  {32'h440960a4, 32'h43279b02, 32'h43290453},
  {32'hc4ef81e7, 32'hc3404366, 32'hc2f89827},
  {32'h439069c6, 32'hc3a72085, 32'hc31d01fb},
  {32'h41f5bd80, 32'h4246a1de, 32'h412e8ad2},
  {32'h44be7aaa, 32'hc0e321c0, 32'hc235c2c6},
  {32'hc4f9a7c4, 32'h43be9478, 32'h41552c79},
  {32'h450595db, 32'h43a0d490, 32'hc304f5ca},
  {32'hc50f6e4a, 32'h4277757c, 32'hc2fb48bf},
  {32'h44f16c73, 32'hc3a8cbea, 32'hc327691b},
  {32'hc4335bd8, 32'hc2aaa225, 32'hc39b67e9},
  {32'h4489616b, 32'h42ad90e1, 32'h4324aab2},
  {32'hc4134d23, 32'hc282a5f3, 32'h419aa440},
  {32'h422ab870, 32'hc345144d, 32'hc33219e2},
  {32'hc40a2730, 32'hc34ff209, 32'h4310f77b},
  {32'h44efc0a4, 32'hc2799f3d, 32'hc1d50bd2},
  {32'hc3f1b900, 32'h43ba42aa, 32'hc3ffd080},
  {32'h442a9b60, 32'h42851546, 32'h432f5449},
  {32'hc2596300, 32'h43402158, 32'h431aec32},
  {32'h44c4bf1c, 32'hc2c243d1, 32'hc39c9216},
  {32'hc21cd248, 32'h4399f38b, 32'h42f6f96c},
  {32'h43e18748, 32'h4281e285, 32'h43832d27},
  {32'hc4be7940, 32'hc30eccbb, 32'hc34bf411},
  {32'h44ca1afd, 32'h41fa6836, 32'h43d8166c},
  {32'hc4c7cfff, 32'h4305134c, 32'h40b587a0},
  {32'h44a44c7c, 32'hc32f4e50, 32'hc283162e},
  {32'hc2e11fd2, 32'hc377f8e4, 32'h4254e8c9},
  {32'h44d510d8, 32'h42b5dfe0, 32'h42adf0c1},
  {32'hc4e72424, 32'hc1946f97, 32'hc2f5aa18},
  {32'h448c5159, 32'h4132e2e3, 32'h419affac},
  {32'hc3917ae0, 32'h430b920f, 32'h440d400a},
  {32'h434bd4e8, 32'hc29f1bb3, 32'h4392c899},
  {32'hc3ca6b8d, 32'h4386f6b5, 32'hc2c8975c},
  {32'h4408f09c, 32'hc3ba9b4f, 32'hc2b10c39},
  {32'hc4eedd22, 32'h435cab2b, 32'hc2575856},
  {32'h43f855e0, 32'hc2d61d44, 32'hc2b96294},
  {32'hc37c40e7, 32'hc3854bd1, 32'hc2591dba},
  {32'h441ac306, 32'hc192ae61, 32'hc3656092},
  {32'hc4f27481, 32'h43cd1a8d, 32'hc3797cfd},
  {32'h436f968a, 32'h4336fef4, 32'hc2f681e2},
  {32'hc4e0ce22, 32'h43466de5, 32'hc31bab67},
  {32'h44e91f0f, 32'h43836aa6, 32'h4377f51b},
  {32'hc50a6fac, 32'hbe1c0646, 32'h439367ee},
  {32'h44d42d83, 32'hc3331c8e, 32'h4364c499},
  {32'hc4dccd70, 32'hc1a2e181, 32'h432b13ac},
  {32'h44a3e93c, 32'hc2fdcfc2, 32'h415c1b34},
  {32'hc5128657, 32'h40b20e8d, 32'h429c2479},
  {32'h44ea37c6, 32'h439c6aaf, 32'h43444a0f},
  {32'hc4e7f7b1, 32'hc3493a1d, 32'h428e2bd8},
  {32'h44de2e8e, 32'hc403a5ba, 32'h420aa20d},
  {32'hc4dbbd03, 32'h437b86c0, 32'hc382c4c2},
  {32'h439d48bc, 32'hc190cb70, 32'hc2d7d127},
  {32'hc4f22fa7, 32'h429d6ee0, 32'h42c0f983},
  {32'h450eec10, 32'h417de096, 32'h43f0cd57},
  {32'hc47aed40, 32'h4319d96a, 32'hc2953e52},
  {32'h44c657c4, 32'h42e2703a, 32'hc33075ca},
  {32'hc47c39f2, 32'h4332ec8a, 32'h43441903},
  {32'h4466c6aa, 32'h436f2e14, 32'h42dea114},
  {32'hc48f3209, 32'h41b977fa, 32'h438a86d1},
  {32'h444fd230, 32'hc37c1c0c, 32'hc44e91e4},
  {32'hc44e19c3, 32'h424900fc, 32'h411423ec},
  {32'h44f569ea, 32'h41d48d04, 32'hc326c45d},
  {32'hc3fd8578, 32'h4280e568, 32'hc31b192b},
  {32'h44ce61c1, 32'hc3cb7d41, 32'hc432b6f3},
  {32'hc4f6d864, 32'hc295b1be, 32'h42c8442d},
  {32'h44ebcd7e, 32'h4343ee49, 32'hc311bf72},
  {32'hc48a4a3a, 32'h42102728, 32'hc35642e7},
  {32'h43ff8d64, 32'hc29c49c6, 32'hc3228e6b},
  {32'hc4799dff, 32'hc20e3962, 32'h43501d12},
  {32'h44aef35d, 32'hc32371f9, 32'h3f172739},
  {32'hc3c0e77c, 32'hc11665ea, 32'h43cd7620},
  {32'h44eee096, 32'h411f8c88, 32'h42e41a2d},
  {32'hc4f8cb37, 32'hc2d74014, 32'h43b39099},
  {32'h444d4380, 32'h429519c7, 32'h4346b745},
  {32'hc3ad193b, 32'hc2fac2ac, 32'h42ae9655},
  {32'h44e77072, 32'h432f49c8, 32'hc32c9321},
  {32'hc5063c14, 32'hc311b717, 32'hc360668d},
  {32'h442b4e10, 32'hc3bd1717, 32'hc316b9f4},
  {32'h436650e5, 32'hc241f66e, 32'h436cd6ee},
  {32'h448f6759, 32'h42ad9ab6, 32'hc2846a0b},
  {32'hc50687d3, 32'hc2d21e0c, 32'h4278899c},
  {32'h44ba9b5a, 32'hc32bb507, 32'hc319f0cc},
  {32'hc4c456c4, 32'h42c01b81, 32'h43880fdd},
  {32'h44a6540d, 32'hc20aa1b6, 32'hc23e85e9},
  {32'hc4ec0d94, 32'h423de9d7, 32'h430dd3f2},
  {32'h4431bc64, 32'h43032974, 32'h432d1cb8},
  {32'hc200b0b0, 32'h43694349, 32'h42bfb961},
  {32'h4494e28a, 32'h42f92af0, 32'h42913a81},
  {32'hc424b8fe, 32'h42bb259d, 32'hc3087ed3},
  {32'h448981fa, 32'hc31e1478, 32'hc36d7b42},
  {32'hc4eab053, 32'hc37020f6, 32'hc2e22687},
  {32'h4359e8dc, 32'hc366665d, 32'hc309d80e},
  {32'hc41e45ec, 32'h42e94de8, 32'h4118e9b5},
  {32'h44cd296e, 32'hc30ce21c, 32'h4455a64b},
  {32'h446c9782, 32'hc3803675, 32'h43855d0b},
  {32'hc4ca4846, 32'h43d51585, 32'h41057348},
  {32'h45007c68, 32'h4332f651, 32'hc0d7b375},
  {32'hc46fb4ea, 32'hc3195d89, 32'h431b5a85},
  {32'h43bd7192, 32'hc3aa4029, 32'hc335cc76},
  {32'h42bc2140, 32'hc3125155, 32'hc3adc5fb},
  {32'h44517e2d, 32'h43792e10, 32'hc3bb764d},
  {32'hc39a3ece, 32'hc3ae4dd3, 32'hc2a13a26},
  {32'h44b6c837, 32'hc2877268, 32'hc2cc0c6a},
  {32'hc4f6dae8, 32'h4324f585, 32'hc34ce0d6},
  {32'h44dc6069, 32'h4210f596, 32'hc2d04e21},
  {32'hc4d3c89b, 32'hc3e2db00, 32'hc152ee05},
  {32'h44eb2825, 32'hc255b134, 32'h42eb6623},
  {32'hc50a6e9d, 32'h438d21c3, 32'hc32eb1e2},
  {32'hc3063878, 32'h40fda391, 32'h43b699c4},
  {32'hc4a86fe1, 32'h43e54238, 32'h42103b74},
  {32'h4510f63e, 32'hc305c4ac, 32'h439abddb},
  {32'hc4c8991a, 32'h43774d68, 32'hc39f9ea8},
  {32'h44db2d6d, 32'hc28c2ea9, 32'h4401895f},
  {32'hc4237f40, 32'hc15c22d6, 32'hc32ce61f},
  {32'h4485bae4, 32'h42cfd5ce, 32'hc295238d},
  {32'hc483cbd2, 32'hc385ba7e, 32'hc31bfd95},
  {32'h4471f325, 32'hc3086dc6, 32'hc419555c},
  {32'hc465ef9e, 32'hc324b914, 32'h4261a5b7},
  {32'h4504dbba, 32'h42a8fb15, 32'h438703fb},
  {32'hc5125d04, 32'hc24574ee, 32'h4329766d},
  {32'h44a7e5eb, 32'hc38baa4d, 32'h41f51484},
  {32'hc494a150, 32'hc2d3cbdf, 32'h43c91a38},
  {32'h44cdd569, 32'h431cce9f, 32'hc3b5e8ff},
  {32'hc421dfae, 32'hc38e1421, 32'hc348a821},
  {32'h44123cf4, 32'h41943e3d, 32'h43118292},
  {32'hc3bc2370, 32'hc3756b16, 32'h4395297b},
  {32'h44bc2ef4, 32'hc280c9a6, 32'h43632bea},
  {32'hc4f5c4cb, 32'hc3a8a0e1, 32'hc2f661d6},
  {32'h43e171d8, 32'h437598ba, 32'hc326aace},
  {32'hc0907000, 32'hc2f224ca, 32'h4368bbbc},
  {32'h44f4f8c2, 32'hc256d219, 32'hc2b74a88},
  {32'hc50bb40f, 32'h43ff5099, 32'hc12262e9},
  {32'h446f88cc, 32'h424fc363, 32'h412acae3},
  {32'hc42242f9, 32'h43ce6818, 32'hc35a48a8},
  {32'h4435b217, 32'h4204acd2, 32'hc06570db},
  {32'hc38c86a4, 32'hc251b1a0, 32'h43dd5e8b},
  {32'h44b30b85, 32'hc39e4626, 32'h43a86a98},
  {32'hc3caf935, 32'hc38dbedb, 32'hc3bd1293},
  {32'h44df7ccd, 32'hc2bf357e, 32'h41e438c7},
  {32'hc4867463, 32'h42748bc3, 32'hc2a3a5d0},
  {32'h442fb30e, 32'h43576986, 32'h42e36b21},
  {32'hc373bc5b, 32'h43377dbc, 32'h4302877d},
  {32'h45184107, 32'h4312c5a9, 32'hc40687ce},
  {32'hc515aa8b, 32'hc1a2123e, 32'hc2e2f334},
  {32'h44c9eecd, 32'h438a8b6a, 32'hc17acc12},
  {32'hc4fa2b12, 32'h431716dd, 32'hc30be321},
  {32'h4302fb11, 32'h40f3ff8a, 32'hc355d0bd},
  {32'hc317b22f, 32'h436dddd1, 32'h440538fc},
  {32'h4509bd4d, 32'h43b0ec58, 32'hc2b95d96},
  {32'hc4e274af, 32'h43bc3216, 32'hc0137b28},
  {32'h442228f2, 32'h4346ed25, 32'h4390c3e8},
  {32'hc46baf37, 32'hc3077821, 32'hc34ac579},
  {32'h44a812c3, 32'h4220682f, 32'h43114bb5},
  {32'hc48ff1c2, 32'hc2ccebdc, 32'hc3af1516},
  {32'h44da77e8, 32'hc30e8793, 32'h41600ad0},
  {32'hc4b081e2, 32'hc3e45fd5, 32'hc32deae1},
  {32'h4418e665, 32'hc38281ea, 32'hc2d7e33d},
  {32'hc4ebf954, 32'h42b07c74, 32'h420edb70},
  {32'h44f0e08d, 32'h441c96a5, 32'hc33d3c9f},
  {32'hc3e01552, 32'h4317f97c, 32'h4233a175},
  {32'h4375a7ce, 32'h430f88aa, 32'hbecba6f3},
  {32'hc42b839c, 32'h4342223c, 32'hc39938c8},
  {32'h43403f78, 32'h4376f144, 32'h43104c3a},
  {32'hc49cc6e2, 32'hc322d23b, 32'hc2eedc4e},
  {32'h440fafdd, 32'hc307950e, 32'h43a9e26b},
  {32'hc42befe8, 32'h41fab350, 32'hc3cfc09b},
  {32'h4455be44, 32'h40e2f907, 32'h43d7cedf},
  {32'hc3f0e13b, 32'h43bc5d46, 32'hc3765ddf},
  {32'h44e268a5, 32'h43a0f4df, 32'h41f1fc1e},
  {32'hc4bc49a4, 32'hc3326dd6, 32'h43c0fb2b},
  {32'h448b30fc, 32'hc340f6de, 32'hc3a6ca9a},
  {32'hc3ab47ee, 32'h44114b0d, 32'hc2763e46},
  {32'h44cd7ba0, 32'hc3a58003, 32'h43a9cc7a},
  {32'hc415fc99, 32'h436453b7, 32'h42fdcc15},
  {32'h45062107, 32'hc2b67372, 32'h4258d04d},
  {32'hc4a09e9c, 32'hc300d13e, 32'hc39d888e},
  {32'h42aeba4e, 32'h430d9084, 32'h430512d3},
  {32'hc50e68e8, 32'h42e3f395, 32'hc34750c4},
  {32'h434deaf0, 32'hc32e17ed, 32'hc31fe99e},
  {32'hc481248e, 32'hc43ef1f1, 32'h42e4e434},
  {32'h44f886cb, 32'h42ed5ee1, 32'hc3d68021},
  {32'hc3de1724, 32'h4318400f, 32'hc328eb38},
  {32'h4425bc30, 32'h428f253c, 32'h4383293e},
  {32'hc4f6753c, 32'hc34caab2, 32'h42118620},
  {32'h43eb9fc0, 32'h420c4af4, 32'hc300a17f},
  {32'hc50e2af9, 32'hc229c022, 32'hc3d3523a},
  {32'h44b26e01, 32'h43a6d922, 32'h434ba59e},
  {32'hc4ab630c, 32'h42216a44, 32'h440e7a61},
  {32'h4417c2a7, 32'hc305697d, 32'h428e1bda},
  {32'hc4c88995, 32'hc0fc1259, 32'h43eb1532},
  {32'h435d785b, 32'hc27fb79d, 32'h43e9c770},
  {32'hc4f50bd7, 32'hc3233d26, 32'h4323c749},
  {32'h44deee43, 32'hc318279d, 32'h425c6f2f},
  {32'hc3bf5c45, 32'hc200f0b2, 32'hc1cd0752},
  {32'h44fcb82e, 32'h43b22e5b, 32'h4314f42b},
  {32'hc481a58f, 32'hc3723c2e, 32'hc28fe53f},
  {32'h44028948, 32'h423adb07, 32'h42acbae0},
  {32'hc3ad08c4, 32'h42a25fd6, 32'h42cb57c2},
  {32'h41f9d390, 32'h4177b586, 32'h4267a0e0},
  {32'hc50ffc32, 32'h430d91a8, 32'h428cc31d},
  {32'h44f35394, 32'h40616080, 32'hc3b3b6d3},
  {32'hc4929b79, 32'hc4025576, 32'hc2258ff3},
  {32'h446ae674, 32'h4201315e, 32'h4331808e},
  {32'hc41af2e6, 32'h42c09fc6, 32'h43abad94},
  {32'h44145544, 32'h42a4d6ce, 32'hc387418e},
  {32'hc492f03c, 32'h4342b8dd, 32'h4325e08b},
  {32'h4497d2f6, 32'hc3acfbde, 32'h43947ad3},
  {32'hc4f09167, 32'hbfb35121, 32'h40b99dfc},
  {32'h448c21ac, 32'h42295a0d, 32'hc259ed19},
  {32'hc4420c6a, 32'hc06aadc0, 32'h42c76211},
  {32'h4487e062, 32'h423ba57b, 32'hc30e2d34},
  {32'hc421a3b7, 32'hc2befe45, 32'hc3900205},
  {32'h44ceab2b, 32'hc3c02247, 32'hc15545fb},
  {32'hc35018fa, 32'h439e280c, 32'h4345e099},
  {32'h44b91768, 32'hc32237b4, 32'hc39c49d6},
  {32'hc506d857, 32'hc3a47f3d, 32'h43e06a35},
  {32'h44326745, 32'h4308e796, 32'h42a02514},
  {32'hc5039f7f, 32'h434d917b, 32'h44277725},
  {32'h44e3382a, 32'h42827324, 32'h427fe39f},
  {32'hc4bd1be8, 32'h42c99d03, 32'hc3070e37},
  {32'h44634a0e, 32'h4324e7f8, 32'hc2f13f67},
  {32'hc36bca50, 32'h43d681ec, 32'h41969c38},
  {32'h44ca9352, 32'hc201b6fc, 32'hc02f5ebf},
  {32'hc4afd7d4, 32'h43c67671, 32'h43535704},
  {32'h450bbee2, 32'h41ed8c4f, 32'h433e9ccc},
  {32'hc2f313c0, 32'h4382848d, 32'h438abc68},
  {32'h439d3bc4, 32'hc341c921, 32'hc357cd2f},
  {32'hc36897b2, 32'hc3d60ecd, 32'hc36f1072},
  {32'h44ab6f7b, 32'h42b8375e, 32'hc37e94b9},
  {32'hc4d60d6a, 32'hc3b49a58, 32'hc1b33bbc},
  {32'h4442099c, 32'hc2f555ed, 32'h4306beb5},
  {32'hc5001d79, 32'h43101524, 32'h4373c427},
  {32'h44b348de, 32'h43adfbe9, 32'h42bb32a1},
  {32'hc4b6509e, 32'hc3c9b720, 32'h41bf40f8},
  {32'h450e67fc, 32'hc243d04e, 32'h4244b42c},
  {32'hc3ef2dcc, 32'hc3ad814d, 32'hc275e93a},
  {32'h4441f44a, 32'h406fb41c, 32'h4358c0de},
  {32'hc4c8af12, 32'hc3e1e2be, 32'h422ec39a},
  {32'h43f67838, 32'hc321d448, 32'h4120875f},
  {32'hc4bb431f, 32'hc2c8dee2, 32'hc30dd255},
  {32'h421ca320, 32'hc34d7c32, 32'hc2e08424},
  {32'hc4829df9, 32'h428c9d98, 32'hc32d0c90},
  {32'h450223d6, 32'hc35e6030, 32'hc3bf6dfb},
  {32'hc5015737, 32'hc2d538c2, 32'h4316bfe7},
  {32'h44b2750d, 32'hc3954f7e, 32'h42e37c28},
  {32'hc506b67c, 32'hc3cae79a, 32'hc2bc99f1},
  {32'h44dd0857, 32'hc2eb220b, 32'hc3b1d511},
  {32'hc40b5bb2, 32'h43087eec, 32'hc38b314b},
  {32'h44bcff96, 32'hc2e485e3, 32'hc40c2192},
  {32'hc4a8ab9c, 32'hc3b8db97, 32'h43530288},
  {32'h4494ba5f, 32'hc32c14e6, 32'hc334b59c},
  {32'h434944d0, 32'h439a678a, 32'h422e95ee},
  {32'h44f6a62a, 32'h41cda6f2, 32'hc367e24a},
  {32'hc32dc7e0, 32'h437147a4, 32'hc2ffdfda},
  {32'h439f07e0, 32'h42fd668d, 32'h43a5a1b5},
  {32'hc4caf3f9, 32'h42fe5dd4, 32'hc28d8a6c},
  {32'h44dc9681, 32'h41b8cb9a, 32'h41861af0},
  {32'hc42c085b, 32'hc3ea32b7, 32'hc33e9372},
  {32'h42b1cd00, 32'hc2a031a8, 32'hc3a243f7},
  {32'hc4d5a3c0, 32'h42e668c4, 32'hc27f89ce},
  {32'h43d59664, 32'h4332c858, 32'h41f0bba9},
  {32'hc4eacbcb, 32'h43b97487, 32'h431ac226},
  {32'h45055047, 32'hc23a09cf, 32'h43d4f32c},
  {32'hc4426f9b, 32'hc2a6e131, 32'h4255fdb0},
  {32'h443b4d62, 32'h4393383e, 32'hc3bc62a2},
  {32'hc5061788, 32'hc36dbcd1, 32'hc2f74b74},
  {32'h4296f5c0, 32'h42ac8f82, 32'hc23c186d},
  {32'hc4d42084, 32'hc31c1b28, 32'hc3320a73},
  {32'h449ba514, 32'hc34ce74f, 32'hc3410cd0},
  {32'hc33d1bb0, 32'hc3db1084, 32'hc3a6266f},
  {32'h4517c9c2, 32'hc383d2a2, 32'h4343d0ef},
  {32'hc3d777f4, 32'hc3ced469, 32'h433b37ce},
  {32'h44199719, 32'h42a501ce, 32'h42a41624},
  {32'hc339bc48, 32'hc2f4815e, 32'h428cb521},
  {32'h4504c086, 32'h42d7dc90, 32'h42a3564e},
  {32'hc4347bac, 32'hc347dfbb, 32'hc395dafa},
  {32'h450a5665, 32'h439daf41, 32'hc396aece},
  {32'hc3573a0c, 32'hc3612506, 32'h43035100},
  {32'h4339771d, 32'hc3aa63de, 32'h4248914b},
  {32'hc43683a6, 32'h4388c4c2, 32'hc38d69fa},
  {32'h441835e6, 32'h425db088, 32'h4113221c},
  {32'hc511297d, 32'hc16be7e4, 32'hc405ce5d},
  {32'h44e5a9dd, 32'hc2db4f84, 32'hc34c5ab1},
  {32'hc50908e3, 32'hc2158554, 32'h426859d6},
  {32'h44a9b716, 32'hc2d9cc1b, 32'h437d418a},
  {32'hc4fef1e3, 32'hc2067d85, 32'h43b65b8d},
  {32'h4463dd04, 32'hc3273e62, 32'hc2d5dd5e},
  {32'hc4227e38, 32'h42532807, 32'h436d010b},
  {32'h440f8c2e, 32'hc32169a7, 32'h43a81b23},
  {32'hc462a1c8, 32'h41eb4245, 32'hc37a1b27},
  {32'h43c220a6, 32'h43cc6039, 32'h43d77d42},
  {32'hc4c49dcf, 32'hc1403d5e, 32'hc2a5eb14},
  {32'h42de1823, 32'h4389f321, 32'h43a0bbc6},
  {32'hc44c4ed7, 32'h4350a84a, 32'h434e77a8},
  {32'h44b97728, 32'h43d31624, 32'hc2ee2c3e},
  {32'hc4167eb0, 32'h42810e12, 32'hc3cd4e18},
  {32'h44a90300, 32'h420b3a2c, 32'h431f4006},
  {32'hc2aaaf7c, 32'hc1063ef2, 32'hc357710b},
  {32'h4515f950, 32'hc39a9a1b, 32'hc252be54},
  {32'hc39b3b04, 32'hc28af5a8, 32'hc11515fc},
  {32'h443a68e7, 32'hc392bdc1, 32'h418d6f88},
  {32'hc485687a, 32'h43eed478, 32'h418a57d6},
  {32'hc2a06f90, 32'h41e36986, 32'h42a87b9b},
  {32'hc3388328, 32'hc2e0bbfa, 32'h432b2552},
  {32'h4508f61b, 32'h42b64545, 32'hc343e343},
  {32'hc4ac37e3, 32'h42779b7d, 32'hc35aadbe},
  {32'h44c5bfcb, 32'hc25f9460, 32'h4330e162},
  {32'hc44e6460, 32'h43434732, 32'h42e79073},
  {32'h43960360, 32'h43202f61, 32'h42676183},
  {32'hc4b2ce7c, 32'hc343cb54, 32'hc2a566e3},
  {32'h44d7ad1c, 32'hc35d5149, 32'hc357be6c},
  {32'hc51106c7, 32'hc3688c02, 32'h43592408},
  {32'h44edf16e, 32'h4379f873, 32'hc3434896},
  {32'hc2b7c3c8, 32'hc2cb992b, 32'h4165a24e},
  {32'h44d1d97c, 32'h426812f3, 32'h424477be},
  {32'hc48825cf, 32'hc3f8b9ce, 32'h437defac},
  {32'hc0f5a3c0, 32'h439b80e2, 32'hc23e7eea},
  {32'hc44b3d26, 32'hc40b7405, 32'hc3802a0d},
  {32'h43eab1b0, 32'hc2fe9f59, 32'hc3cf6ae2},
  {32'hc424aeee, 32'h42962437, 32'h43814cca},
  {32'h44e7c8c0, 32'h43116ea6, 32'hc36244a9},
  {32'hc5144f75, 32'h42a371de, 32'h4360a0fd},
  {32'h44a0e891, 32'hc34b42bd, 32'hc0cd6eee},
  {32'hc4a55b52, 32'hc27e2626, 32'hc37468d8},
  {32'h442e9e84, 32'hc222a022, 32'h42e997a0},
  {32'hc5007125, 32'hc2c045b3, 32'h43a99b64},
  {32'h4482e9ec, 32'hc36129e4, 32'h41d51fe7},
  {32'hc416e9ad, 32'h41dd8fd6, 32'h43508ce1},
  {32'h44f9c6fa, 32'hc2aa5410, 32'h419fafa8},
  {32'hc4b9c4f6, 32'h4357ae6a, 32'h43b91058},
  {32'h445a78b9, 32'hc28899b3, 32'h4214c6be},
  {32'hc49767c2, 32'hc302cffa, 32'h4156df5d},
  {32'h4449d6aa, 32'hc3d7588e, 32'hc3aa3a1e},
  {32'h42a71920, 32'hc3fa370a, 32'hc2e6130c},
  {32'h44d73425, 32'h44075351, 32'hc38e0c43},
  {32'hc430f0d8, 32'h438938e6, 32'hc330d5d7},
  {32'h44cd96d0, 32'hc32ac88a, 32'h43663afe},
  {32'hc4bb4849, 32'h43079b1f, 32'hc3563305},
  {32'h42ccba30, 32'hc2b5f907, 32'hc34c12b1},
  {32'hc41aca44, 32'hc38d9719, 32'h43d5143a},
  {32'hc3ad5568, 32'h4386d20a, 32'h430de43a},
  {32'hc4ea116c, 32'h411919d7, 32'hc3876328},
  {32'h44cb7a2d, 32'h43a1fe94, 32'hc2f265b6},
  {32'hc47878a2, 32'hc2aaa955, 32'h42f87e73},
  {32'h43bf8db4, 32'h423eb5b8, 32'hc310abfe},
  {32'hc41d5a2d, 32'hc3400953, 32'h430b0077},
  {32'h439a23e0, 32'hc23b4bff, 32'hc3171627},
  {32'hc2300588, 32'h436e61f4, 32'hc33acf13},
  {32'h44c3476e, 32'hc40d5777, 32'h437f4e7a},
  {32'hc4feb50f, 32'hc387d5f1, 32'hc358ecbc},
  {32'h43d099fc, 32'h412fc181, 32'hc3824000},
  {32'hc4075c8d, 32'h42cb658a, 32'hc2595bad},
  {32'h438ec8b4, 32'h438fa186, 32'hc2b9b1d8},
  {32'hc32e1daa, 32'h42db9d1a, 32'hc38c861b},
  {32'h43fa2b2f, 32'hc25b2dec, 32'h438d713a},
  {32'hc30a717c, 32'hc3ba9193, 32'hc225e332},
  {32'h451e5a17, 32'h42db13d5, 32'hc3758847},
  {32'hc4a5c118, 32'h43beb9d2, 32'h420303bd},
  {32'h446a495c, 32'hc3c5ac7b, 32'hc3931257},
  {32'hc4751064, 32'hc257f104, 32'h3fa5e9ba},
  {32'h44e0cc09, 32'h4325d8a5, 32'hc3756d9b},
  {32'hc43303e7, 32'hc3362c24, 32'h442ddbc2},
  {32'h449e4600, 32'h41d23d71, 32'hc1d2e48a},
  {32'hc4ead62c, 32'h42851eb1, 32'hc35a9d22},
  {32'h44f13ab2, 32'hc26bde3e, 32'hc2a089c1},
  {32'hc4dde9b0, 32'hc4407b86, 32'h436dfd9a},
  {32'h43b13901, 32'hc3787ae4, 32'hc394010d},
  {32'hc38037fc, 32'hc355f960, 32'h42636e1e},
  {32'h4516aa3a, 32'hc12c29e3, 32'hc2e27d1f},
  {32'hc49128be, 32'hc33db872, 32'h426c1d2d},
  {32'h4520cbfb, 32'h42887086, 32'hc3c83d3c},
  {32'hc5085df1, 32'hc1a1bdf0, 32'hc108b53f},
  {32'h44da5a8d, 32'hc2d2c0f6, 32'hc2877426},
  {32'hc4e91985, 32'hc398b9ae, 32'hc34dce46},
  {32'h450bed8e, 32'h42f14418, 32'hc3a74c45},
  {32'hc491f0a3, 32'hc31a7671, 32'hc28cae82},
  {32'h4468b772, 32'h410c7b3d, 32'hc097deb8},
  {32'hc4d2c8ee, 32'hc343a55d, 32'h43876d9b},
  {32'h45307324, 32'hc14ea16e, 32'h439019f7},
  {32'hc2d80420, 32'hc3801634, 32'hc1d1128e},
  {32'h447cbfa4, 32'h4382ff7c, 32'h433ca7fe},
  {32'hc40b2976, 32'hc266e969, 32'h42cdd455},
  {32'h4402370e, 32'h43cb6821, 32'h4334b6f9},
  {32'hc18eca56, 32'h43c91a84, 32'h438768e0},
  {32'h4511cf93, 32'h43343b5d, 32'h421b29c3},
  {32'hc5082b44, 32'hc347ea0e, 32'hc418d74d},
  {32'h44f04a88, 32'h429fb6fd, 32'h43114637},
  {32'hc4829882, 32'h42201531, 32'h4308fdd4},
  {32'h44729ce6, 32'h4340ce49, 32'h42ec367b},
  {32'hc4342875, 32'hc39ce2c5, 32'hc35cd6ff},
  {32'h4417591c, 32'h427e4368, 32'hc19e08b1},
  {32'h43107ea0, 32'h43569095, 32'hc271df34},
  {32'h449fe1ed, 32'hc2e298aa, 32'hc24c3d11},
  {32'hc45921ff, 32'h43451896, 32'h4355b6b8},
  {32'h43e396f0, 32'h41916bdc, 32'h440a5627},
  {32'hc4d4d359, 32'h42b4c8f0, 32'hc1f86d82},
  {32'h44edde68, 32'h42e21cc9, 32'hc3ae2f05},
  {32'hc51e954b, 32'hc3200a50, 32'hc159fa20},
  {32'h44e2b481, 32'hc3bd67c4, 32'hc32254fd},
  {32'hc4bd20dc, 32'hc2aa5f05, 32'h420218e4},
  {32'h4505106c, 32'hc3266b97, 32'h42fe77db},
  {32'hc5007b26, 32'hc3ad311e, 32'h442a44ad},
  {32'h4510c96b, 32'h42d8b8ef, 32'h43e8681c},
  {32'hc3609d10, 32'h4357431a, 32'h417f348a},
  {32'h4399ac32, 32'h4286666f, 32'hc338b02a},
  {32'hc4bde023, 32'h42296b2a, 32'h43393ee4},
  {32'h43b27e5e, 32'hc32a352a, 32'h429b9a1c},
  {32'hc4cb36b7, 32'hc2c93868, 32'hc3598904},
  {32'h44b6438e, 32'h4318c6e9, 32'hc3e26f19},
  {32'hc45542ee, 32'h43735d25, 32'hc370caf5},
  {32'h45118156, 32'h436faa34, 32'h428e5973},
  {32'hc4780ef8, 32'h3f055ab7, 32'h434c31a7},
  {32'h44e2a866, 32'h43c34681, 32'hc30ccf8c},
  {32'hc4d22400, 32'hc3aff2da, 32'hc31d4a8a},
  {32'h4512a78a, 32'hc37ae17c, 32'h433b0ab5},
  {32'hc3a22292, 32'hc40a5472, 32'hc1d63cf2},
  {32'h43fa0a54, 32'hc09e558d, 32'hc31fa648},
  {32'hc40218d8, 32'hc33efcab, 32'hc2a4a3a9},
  {32'h43d0ce20, 32'h42b2f491, 32'hc31152aa},
  {32'hc462323f, 32'h43c50016, 32'hc21c59d2},
  {32'h4488942a, 32'hc1592882, 32'hc3964085},
  {32'hc348f4f4, 32'hc28f8fd6, 32'h42dda300},
  {32'h4514ceb8, 32'h42243ced, 32'hc31c0b15},
  {32'h437c14e0, 32'hc186b61c, 32'h42365e66},
  {32'h4523d8c0, 32'h42dd9d08, 32'hc225b7c8},
  {32'hc4c009fe, 32'h43807aa1, 32'hc207b8e4},
  {32'hc1e37f00, 32'hc329b4a2, 32'h433cead1},
  {32'hc4368544, 32'h43e37fb4, 32'hc3d1078f},
  {32'h44b5d2c6, 32'hc338f50c, 32'h42b1f353},
  {32'hc50a1ca9, 32'hc35189d8, 32'h42f2c4f7},
  {32'h45107fbe, 32'hc3e09a3b, 32'hc3aa80f8},
  {32'hc2cb4140, 32'h4176f108, 32'hc303f91b},
  {32'h4387e940, 32'hc32ad738, 32'h43b1f830},
  {32'hc3ee5802, 32'hc35aa6f2, 32'hc2861dcd},
  {32'h438e509a, 32'h431b7edc, 32'h436df3c7},
  {32'hc491f930, 32'hc382d1b5, 32'hc3a35a91},
  {32'h45099db6, 32'hc3857272, 32'hc3db2353},
  {32'hc4c29734, 32'hc274f7ea, 32'h436dcecf},
  {32'h45112e21, 32'h4385c53c, 32'h42ee3d44},
  {32'hc4daac1d, 32'hc308924e, 32'hc2dc93f9},
  {32'h4509b55e, 32'hc33796ad, 32'hc2116256},
  {32'hc48f4c00, 32'h43a3bc8b, 32'hc2a8702e},
  {32'h44b36fd5, 32'h429f3fe7, 32'hc2f70979},
  {32'hc495db32, 32'h4206b463, 32'hc2fc069f},
  {32'h44e61385, 32'h41c1e105, 32'hc2906f0f},
  {32'hc50147e1, 32'h43862a01, 32'hc1cf60f7},
  {32'h44af7dba, 32'hc33c5628, 32'hc38f5c0f},
  {32'hc48dd06b, 32'hc2a2618e, 32'hc1e68bc2},
  {32'h4512a49a, 32'h42109b05, 32'h435703f5},
  {32'hc4f99822, 32'hc194a712, 32'h43a765cc},
  {32'h44a4fb86, 32'hc22caff8, 32'hc2cdcad9},
  {32'hc421d998, 32'hc385f04d, 32'h4358772c},
  {32'h446016aa, 32'h438af8f4, 32'h405a6ccb},
  {32'hc4948a40, 32'hc1d7636c, 32'hc1258dea},
  {32'h44d43a8d, 32'h421e5cc0, 32'h439c3e55},
  {32'hc4c2854c, 32'hc29cb67a, 32'hc31646b2},
  {32'h424940e0, 32'hc2ee08d0, 32'h4330ad63},
  {32'hc4b8ac61, 32'h437c52c3, 32'h42d52bcc},
  {32'h444f4835, 32'hc37a468d, 32'h4327bcb5},
  {32'hc4b3468b, 32'hc2dcdfe3, 32'hc218d3bc},
  {32'h450b96d6, 32'h4303b1e0, 32'hc2914fc2},
  {32'hc42a2685, 32'hc26e6948, 32'h440ac28f},
  {32'h450c74d0, 32'h43bdc6fe, 32'h4307fd9a},
  {32'hc492e5f9, 32'hc39f36b2, 32'h4258f2e5},
  {32'h445913dc, 32'hc34f77f6, 32'h4292edb5},
  {32'hc4de3be4, 32'hc322d7fc, 32'hc3283f6b},
  {32'h43e4ffce, 32'h43480a12, 32'h429cf456},
  {32'h42a54598, 32'hc330dcc1, 32'hc19e0e22},
  {32'h443a6236, 32'hc2f61db5, 32'hc2738017},
  {32'hc4801af5, 32'hc33d2ec9, 32'h43846ed9},
  {32'h441f61a4, 32'h430be911, 32'hc3c1d22b},
  {32'hc3079e65, 32'hc39c9f38, 32'h431a45cf},
  {32'h4506c5a5, 32'h438cc332, 32'h42e204aa},
  {32'hc4ecbacf, 32'hc335c076, 32'h43a58bf3},
  {32'h44a15fe0, 32'h430852ab, 32'h43811735},
  {32'hc466fa92, 32'hc28a7a07, 32'h43adb976},
  {32'h446c1d0a, 32'hc304994a, 32'h41b3d4df},
  {32'hc42f7960, 32'h420906ff, 32'hc2fddc52},
  {32'h44a8f30c, 32'h42ba6745, 32'h4304ba44},
  {32'hc4f6a7d3, 32'hc22c5ea2, 32'h435fc96c},
  {32'h448d7efc, 32'hc2a89963, 32'h426d7907},
  {32'hc451d1bc, 32'hc313032d, 32'hc1eed0be},
  {32'h4508d0b6, 32'h43a620be, 32'h43967b8f},
  {32'hc4932dca, 32'hc3da983d, 32'hc39322e7},
  {32'h4503671f, 32'hc3599b7d, 32'hc2b88d64},
  {32'hc4e3db97, 32'h438fa0ec, 32'h441778f1},
  {32'h45075ac0, 32'hc292d6be, 32'h439406b4},
  {32'hc448de87, 32'hc27d9f56, 32'hc353032c},
  {32'h4505b108, 32'h4148a9a8, 32'hbfb63660},
  {32'hc4520984, 32'h43057c56, 32'hc3b76fab},
  {32'h44bc813d, 32'hc2c42755, 32'hc217f244},
  {32'hc3bb0b08, 32'hc397766a, 32'hc3874f73},
  {32'h44a92590, 32'h43e61b72, 32'hc344937d},
  {32'hc503fd40, 32'hc265b2a4, 32'hc332475e},
  {32'h437b124e, 32'h43d9ae8b, 32'h431b8e4e},
  {32'hc50df4c0, 32'hc3991272, 32'h43018f3d},
  {32'h449305a8, 32'hc33a5236, 32'h438ee7ce},
  {32'hc40d760c, 32'h42fc8fd0, 32'hc3fef186},
  {32'h450e88a3, 32'hc35ba86b, 32'hc184eed9},
  {32'hc4b7579d, 32'hc3705e52, 32'h42013556},
  {32'h450d872b, 32'hc379b219, 32'h4219b2bb},
  {32'hc3c3cc10, 32'h41f6373e, 32'hc3a1b332},
  {32'h4438eba2, 32'hc2553670, 32'h42b363a7},
  {32'hc4c34566, 32'h426f4ce6, 32'hc19aba91},
  {32'h44524a54, 32'hc22e71dc, 32'h43c2e4c1},
  {32'hc508a4d3, 32'hc1f2c7b2, 32'hc3c469bf},
  {32'h440078d2, 32'hc29f5f67, 32'hbfd74670},
  {32'hc4aa1ce4, 32'hc2d124af, 32'h43989135},
  {32'h44d7dcfc, 32'hc27396ed, 32'h420b2ca3},
  {32'hc4603866, 32'hc2d710a6, 32'hc36de473},
  {32'h44d764c6, 32'h4324abfd, 32'h43156796},
  {32'hc5099a59, 32'h42a137e8, 32'h428f19fa},
  {32'h44e96340, 32'hc17f64f6, 32'h42ccd1ff},
  {32'hc4730670, 32'hc288b87c, 32'h42040fa4},
  {32'h4446580f, 32'hc22700c6, 32'hc2b231af},
  {32'hc3b357e8, 32'hc2e6a940, 32'h4385ea32},
  {32'h45071941, 32'h411c741e, 32'h43872917},
  {32'hc3ed9bea, 32'h438cedf8, 32'hc3347894},
  {32'h44d6fce3, 32'hc2b1c550, 32'hc1e27a2d},
  {32'hc4f3d472, 32'hc2a21af1, 32'hc30de9db},
  {32'h44a0d3e9, 32'hc1acebdb, 32'hc2bdcdb4},
  {32'hc4eacc99, 32'hc333388d, 32'h438cf716},
  {32'h44e08fd5, 32'hc341243a, 32'h43249008},
  {32'hc4564bcf, 32'hc38ad4e2, 32'hc147e100},
  {32'h452622d3, 32'hc3a7fef3, 32'hc32a73c6},
  {32'hc2ce6dd8, 32'hc2bad790, 32'hc2535020},
  {32'hc093c7e0, 32'hc369b511, 32'hc2f6b134},
  {32'h44f73d2a, 32'hc40961b3, 32'hc307687b},
  {32'hc4805552, 32'hc3cd987b, 32'h43e9d8ef},
  {32'h44cf910a, 32'h43e32bd0, 32'hc24e30e6},
  {32'hc49fbe56, 32'h3feda6c8, 32'hc3a02385},
  {32'h448f54f7, 32'h42cbbf3d, 32'h4428998a},
  {32'hc4c3de76, 32'hc3cd2ba0, 32'h430b59b8},
  {32'h44b78585, 32'h42a05fcb, 32'h43e82dcf},
  {32'hc4896c03, 32'h43b399d8, 32'hc3563cda},
  {32'h449d6872, 32'h43aef4f6, 32'hc38c6375},
  {32'hc4eb214b, 32'hc38bf35a, 32'hc329da4c},
  {32'h4506ac46, 32'h4403cd28, 32'hc274d384},
  {32'hc4588434, 32'hc28e9d24, 32'h42f91292},
  {32'h449279d7, 32'h43bc22a0, 32'hc1e16f06},
  {32'hc456c418, 32'h4311e801, 32'hc2984a42},
  {32'h44a20fe4, 32'hc20e8a33, 32'h43abcf3f},
  {32'hc4ec14c2, 32'h4280f03a, 32'h42d16e41},
  {32'h43fd10cc, 32'hc3403b73, 32'h42b55cbf},
  {32'hc35cdeac, 32'hc0e399d6, 32'hc255bdd3},
  {32'h44572b54, 32'h4248b0ae, 32'h42f7dfa3},
  {32'hc50a4000, 32'hc33d5555, 32'hc3b0abf9},
  {32'h44b34ac3, 32'h4363fe50, 32'h4301b6e5},
  {32'hc49ac4b0, 32'h42a10c92, 32'h43212f7e},
  {32'h443b8876, 32'h42c28450, 32'h4355cdb6},
  {32'hc48d40d2, 32'hc325193e, 32'h421f954f},
  {32'h451f6b20, 32'hc3598205, 32'hc27f22b7},
  {32'hc4b92b55, 32'hc31d8e1d, 32'h426c23b2},
  {32'h44185610, 32'h41d31bd8, 32'h4315b7c6},
  {32'hc44e5d3e, 32'hc3304637, 32'hc376a515},
  {32'h43ed85f0, 32'h42bddc59, 32'h4363716a},
  {32'hc4616337, 32'h438a3179, 32'hc2b7db26},
  {32'h43fa9a18, 32'hc2d8d30a, 32'h42c270d1},
  {32'hc4ea917a, 32'hc3810f03, 32'h428322c6},
  {32'h44715b0f, 32'h43a8c064, 32'h42b69286},
  {32'hc413850a, 32'hc2bf0e06, 32'hc381d072},
  {32'h4417a5f1, 32'h4309526c, 32'hc32501a9},
  {32'hc4495027, 32'hc38ddb8f, 32'h432d99ee},
  {32'h44b21db1, 32'hc2277421, 32'h42772d10},
  {32'h4369ff66, 32'hc2acf8de, 32'h4369df54},
  {32'h45016a74, 32'hc38130ea, 32'h43a03321},
  {32'hc4c38f50, 32'h438248e9, 32'h430e0994},
  {32'h441d9e5c, 32'hc1aa6e76, 32'hc2ddc3f0},
  {32'hc50f2655, 32'h4340539d, 32'h41e612ec},
  {32'h45063e8a, 32'hc425b9e4, 32'h43993ebf},
  {32'hc4d101e8, 32'hc393a9a9, 32'h43ea4130},
  {32'h44eb3e0a, 32'h41555de4, 32'h440044b5},
  {32'hc4a6deef, 32'hc2d09870, 32'hc2a2114f},
  {32'h4462c9d6, 32'h42d7eb32, 32'h43c83e0f},
  {32'hc488a5bf, 32'h433a63ad, 32'h42a6b976},
  {32'h44b3bf56, 32'hc27b592c, 32'hc373181f},
  {32'hc5212e42, 32'hc1d3ff88, 32'h43a4b632},
  {32'h44caca5e, 32'hc38a4002, 32'h434e23ff},
  {32'h43a2d899, 32'hc3350ea4, 32'h432d2406},
  {32'h44a1b472, 32'hc22dd88a, 32'h43a64eb6},
  {32'hc38171e2, 32'hc3a7ce8b, 32'h42b5e7ae},
  {32'h44e1bb12, 32'hc150e554, 32'hc41ada7f},
  {32'hc4f3bec3, 32'hc3442203, 32'h431d726a},
  {32'h45025e39, 32'hc30548a8, 32'hc347bf52},
  {32'hc3c50666, 32'hc1bfe853, 32'hc3b8da39},
  {32'h4499f162, 32'hc1ca4968, 32'hc28b07d1},
  {32'hc45d3950, 32'hc2ba58e5, 32'hc345fc11},
  {32'h435113e2, 32'hc398478a, 32'h42ba8fa9},
  {32'hc40e4a14, 32'hc3924a61, 32'hc2d466fa},
  {32'h443aded9, 32'h4302425d, 32'h42456301},
  {32'hc456a493, 32'h430ca3f8, 32'hc2121e9d},
  {32'h43d33f20, 32'h43ba4dd0, 32'h43ddd3c5},
  {32'hc447d070, 32'h419410f6, 32'hc391abdf},
  {32'h445e67f4, 32'h4251c006, 32'hc365e7c8},
  {32'hc501ac72, 32'h4365e0f8, 32'hc32212fb},
  {32'h450224e5, 32'h437b68a8, 32'hc3850205},
  {32'hc4d0d490, 32'h4359b057, 32'hc2a9f162},
  {32'h448e99c1, 32'h43133d1e, 32'h43c1c39b},
  {32'hc41a8560, 32'hc379ce3a, 32'h43b9587a},
  {32'h448c5f26, 32'h4352b61b, 32'h430c083e},
  {32'hc4a0a108, 32'hc35b8b0c, 32'h433976aa},
  {32'h42a6d430, 32'hc303503d, 32'hc3b5f860},
  {32'hc36687a0, 32'hc2b5cc3a, 32'h434b2e2c},
  {32'h44eac973, 32'hc2d1d113, 32'hc33c4db0},
  {32'hc367e040, 32'hc1584c24, 32'hc2c06334},
  {32'h44bdf2bc, 32'h41078e6d, 32'hc3648c94},
  {32'hc5134356, 32'h429ead89, 32'hc38b8c9e},
  {32'h443c4dd4, 32'h409b7aef, 32'hbec676b2},
  {32'hc4eb7bac, 32'hc361d045, 32'hc328004e},
  {32'h451ed234, 32'hc209dd1e, 32'h4283966c},
  {32'hc44582ca, 32'h4382ad50, 32'h438e3068},
  {32'h4413625c, 32'hc323ec42, 32'hc3618452},
  {32'hc4e517be, 32'h42ff25b3, 32'hc323a595},
  {32'h4507d420, 32'hc3583c9f, 32'hc383a336},
  {32'hc40ed224, 32'hc3fe0706, 32'h41e7f58c},
  {32'h43074134, 32'hc2d060ed, 32'h43157bcf},
  {32'hc3b58c2e, 32'hc2aa6e52, 32'hc2a23b3e},
  {32'h44d95189, 32'hc35e3f6c, 32'h42e09fc2},
  {32'hc423b8f2, 32'hc397a511, 32'h438d5594},
  {32'h44c0c711, 32'hc38154dc, 32'hc36bf49d},
  {32'hc464963e, 32'hc14e3e0c, 32'h438f0aca},
  {32'h44a1d575, 32'h4014ce54, 32'hc3044713},
  {32'hc4a0b308, 32'h434d49fb, 32'h43ea4004},
  {32'h450c2848, 32'h43b51729, 32'hc3b5d475},
  {32'hc4690d86, 32'h425e82bd, 32'h426b5ce7},
  {32'h44d28bfb, 32'hc30de1a4, 32'h430d3e37},
  {32'h42cb827a, 32'h43a954d3, 32'h43169638},
  {32'h4485ef98, 32'h436f020a, 32'hc2ec7ab4},
  {32'hc50fa6ad, 32'h43359318, 32'hc24296de},
  {32'h44b61919, 32'h43e7c89d, 32'h439d3011},
  {32'hc3ef78fc, 32'hc3a72cf7, 32'h43db6b83},
  {32'h44a2a519, 32'hc2724681, 32'hc2c44aea},
  {32'hc19eae00, 32'hc29d1b45, 32'h4324eeb4},
  {32'h42c96310, 32'hc3373c2c, 32'h438a6dc7},
  {32'hc4950f7a, 32'hc384b703, 32'h42ba1502},
  {32'h44cb85f9, 32'h4272367a, 32'hc350b251},
  {32'hc5017286, 32'hc30f9bbe, 32'h42072f73},
  {32'h44cd16ea, 32'h42f4bf40, 32'h4313eeaf},
  {32'hc40ad3ba, 32'hc3a90c3c, 32'h3f77ed02},
  {32'h44e86f72, 32'hc370e20e, 32'h418d3e8a},
  {32'hc36e4126, 32'hc1cdb0dc, 32'h430d0c00},
  {32'h44dbe7b5, 32'h43962b48, 32'hc3cab93a},
  {32'hc4bb9fe6, 32'h42e27a63, 32'h442b146a},
  {32'h448539fc, 32'hc3eb60ba, 32'hc36ea94e},
  {32'hc4021354, 32'hc294c0cd, 32'hc359c178},
  {32'h43ce7f50, 32'hc3285da7, 32'hc3599e26},
  {32'hc494fc7e, 32'hc3202839, 32'h4344166d},
  {32'h445ae6d6, 32'hc3b03e1e, 32'hc2e27e25},
  {32'hc2b4fe6d, 32'h43ab96ca, 32'h43569a45},
  {32'h44f87532, 32'h430859a2, 32'h43d6bfe8},
  {32'hc41a61b8, 32'hc35e2062, 32'h437c7a31},
  {32'h4482f3ed, 32'h41a2cf5d, 32'hc2990bb7},
  {32'hc4dc3291, 32'h435a7fae, 32'hc268c52d},
  {32'h44f2e28b, 32'hc2716e2e, 32'h420ecb2a},
  {32'hc4001aab, 32'h42683140, 32'h41ba2edf},
  {32'h44bcc661, 32'h42bf01b0, 32'hc3070fea},
  {32'hc4eb573f, 32'h43349be9, 32'hc2d07718},
  {32'h43d0e9a0, 32'hc3484fdf, 32'h43503e78},
  {32'hc49c7580, 32'h43885472, 32'h43c21bdd},
  {32'h452f9fdc, 32'h43687340, 32'hc240741c},
  {32'hc439bcd1, 32'h439101b6, 32'hc3c7fe82},
  {32'h43410d90, 32'hc32f35bc, 32'hc409d131},
  {32'hc36e9938, 32'h43a2343b, 32'h4325b25d},
  {32'h450388a4, 32'h433fdf92, 32'hc2a76ef3},
  {32'hc4608308, 32'hc2ee7abc, 32'h42afd19f},
  {32'h449c97c0, 32'h43b2839b, 32'h437e658e},
  {32'hc5015b3c, 32'hc334dd60, 32'h4385275c},
  {32'h447ad790, 32'hc20e88a2, 32'h429da732},
  {32'hc48284d3, 32'hc3e45671, 32'h44465377},
  {32'h445dadb7, 32'h42c28f4a, 32'hc3d849b0},
  {32'hc48d6a48, 32'hc39e712f, 32'h42f65b90},
  {32'h43c4fadc, 32'h426c1632, 32'h430fd104},
  {32'hc4c93a87, 32'hc36d44e8, 32'h43544c87},
  {32'h449f6280, 32'h41809c39, 32'hc1c31736},
  {32'hc423e144, 32'h41d94270, 32'h435b67f5},
  {32'h44ff273b, 32'hc34021f9, 32'hc24ad7ca},
  {32'hc4c4cf35, 32'h428ffe9a, 32'hc2232529},
  {32'h441403da, 32'h42419388, 32'h432b46f4},
  {32'hc4244943, 32'hc239542c, 32'h432134f5},
  {32'h44936a67, 32'hc3dcb8b7, 32'hc3d5aa03},
  {32'hc49c9868, 32'h432db040, 32'hc390ea7b},
  {32'h44ff3ba6, 32'h432f5419, 32'hc22cd17f},
  {32'hc4168abe, 32'h43559c90, 32'h424ea343},
  {32'h428fe558, 32'h41791d93, 32'h43b62c4d},
  {32'hc41b80a4, 32'h4362c302, 32'hc419772c},
  {32'h44fb1046, 32'h43223c44, 32'hc39395a6},
  {32'hc43ee395, 32'hc1f47f53, 32'hc36d36ea},
  {32'h442bd950, 32'h3e8b1b00, 32'hc3865337},
  {32'hc492501a, 32'h434a5c06, 32'h43223a19},
  {32'h44e8cf8c, 32'hc3c3c7ea, 32'hc2785cf4},
  {32'hc4e068c2, 32'hc03625e1, 32'h434360f7},
  {32'h4514d888, 32'h431f54d7, 32'h433ed815},
  {32'hc4101a64, 32'hc31c59e7, 32'hc390539e},
  {32'h44f590a2, 32'hc361a279, 32'hc2e468e7},
  {32'hc48814b0, 32'h43809b27, 32'hc30280cb},
  {32'h4411010e, 32'h438be5b6, 32'hc2061ee8},
  {32'hc2af87f0, 32'h435d4536, 32'h4380c3fa},
  {32'h44a62623, 32'hc2638a4e, 32'h43cc44f1},
  {32'hc4e191bc, 32'h43c50fe4, 32'h4386babf},
  {32'h44be0dad, 32'hc31d10cf, 32'hc400d224},
  {32'hc5070f79, 32'hc350c749, 32'h43201265},
  {32'h44f25288, 32'h41e25738, 32'h4259e16e},
  {32'hc47d55fe, 32'hc2d5f265, 32'h43b7aa9f},
  {32'h4503d309, 32'h42df48d6, 32'hc1c95c91},
  {32'hc41830ee, 32'hc2c7e26e, 32'hc38b4865},
  {32'h450e8f26, 32'h42accd38, 32'h423adb8f},
  {32'hc4b2e59a, 32'h430d7800, 32'h42a4d224},
  {32'h44d9c4ba, 32'hc385b006, 32'h424da5d6},
  {32'hc443d6b5, 32'hc38fe2ae, 32'hc26c1722},
  {32'h44c5f309, 32'hc27160b9, 32'h43601643},
  {32'hc3948874, 32'h40de14e8, 32'h4258a343},
  {32'h447bf737, 32'h43a8f284, 32'h4290870a},
  {32'hc4546fca, 32'hc3048df6, 32'hc2b28fd7},
  {32'h451f5509, 32'h437ce797, 32'h4124362e},
  {32'hc506cb36, 32'hc2aff49b, 32'h4239330d},
  {32'h4480a5bb, 32'hc1d15c79, 32'hc2ad3ee8},
  {32'hc51161d6, 32'h43042043, 32'hc21547e1},
  {32'h43372418, 32'h431a2bb1, 32'h4372b8e3},
  {32'hc4a4561f, 32'hc38a73f6, 32'h43226eb5},
  {32'h445e26f5, 32'h4369b85b, 32'h428a69cb},
  {32'hc50306b5, 32'hc29900a7, 32'hc2abc159},
  {32'h45055e30, 32'h429b2c23, 32'hc3bc168f},
  {32'hc4f1faf4, 32'h4380a8e4, 32'h42a772ae},
  {32'h4518b77b, 32'h43b91339, 32'h440aa829},
  {32'hc4482586, 32'hc35abc71, 32'hc39d7f29},
  {32'h4456701e, 32'hc062cb1e, 32'h420b90b2},
  {32'hc506ba94, 32'h435a5582, 32'h438ffb0b},
  {32'h45220962, 32'h430b78a6, 32'h43df52ef},
  {32'hc49f3677, 32'hc3c537a3, 32'hc1ebaa9a},
  {32'h4458d341, 32'hc3766d5a, 32'hc31ddfa8},
  {32'hc482df64, 32'hc3c1957e, 32'hc296005a},
  {32'h4324b4f8, 32'h43650fa2, 32'hc353fb5e},
  {32'hc330cb00, 32'h43ad766c, 32'hc2fbdfe5},
  {32'h4454ff78, 32'hc3b1af3d, 32'h433ec6ca},
  {32'hc48f5a0e, 32'hc25ead29, 32'hc269b4e6},
  {32'h43f93e84, 32'hc37b5c37, 32'hc3cf7743},
  {32'hc49c0a0e, 32'hc38d0d96, 32'h4221ad15},
  {32'h43bc5a2c, 32'hc2d8c848, 32'hc2ff6888},
  {32'hc2e28f10, 32'h43026032, 32'hc33da194},
  {32'h44edb469, 32'h43662855, 32'hc08f6d00},
  {32'hc4d19ff0, 32'h438101c1, 32'h43724372},
  {32'h44381e72, 32'hc35b12cd, 32'h42afbed7},
  {32'hc4749152, 32'hc15627fc, 32'hc393aec2},
  {32'h448f4035, 32'h428e0381, 32'h43195978},
  {32'hc40912e0, 32'hc2bf4782, 32'hc0ab0c90},
  {32'h44e01be7, 32'hc2a400da, 32'hc2934218},
  {32'hc50e85ce, 32'hc3c49022, 32'h41558cd7},
  {32'h44ffde6c, 32'h43714cf0, 32'hc1f278a8},
  {32'hc4105fcb, 32'h435ca7df, 32'h43836c7f},
  {32'h449cab83, 32'hc2a01216, 32'hc37fd536},
  {32'hc4e19aa6, 32'hc3b7cee3, 32'hc0d21760},
  {32'h4488309e, 32'h42c5480c, 32'hc301b3d9},
  {32'hc47001d6, 32'hc2b31391, 32'hc3bdc54b},
  {32'h44e3aea9, 32'h43805937, 32'h42e8ea87},
  {32'hc37b9981, 32'hc3a22a76, 32'h42658b4f},
  {32'h44ee4d6a, 32'hc1bb3b52, 32'hc2eda426},
  {32'hc50896da, 32'hc30c86ee, 32'hc18ecdc2},
  {32'h43863790, 32'hc2f562df, 32'hc21a1792},
  {32'h42cdb3d6, 32'hc233ca3e, 32'h42a7e1fe},
  {32'h4493df1c, 32'hc16e8615, 32'h43a3dc12},
  {32'hc496899e, 32'h4252cb9c, 32'h3e129e78},
  {32'h44270d1c, 32'h428349c6, 32'hc2803983},
  {32'hc4108d54, 32'h431c4ef1, 32'hc309875e},
  {32'h450413b8, 32'hc2d23759, 32'h43e2647f},
  {32'hc4ef5505, 32'hc32aa5b2, 32'hc2149417},
  {32'h444eb47a, 32'hc31fa8b9, 32'h42a5653a},
  {32'hc48674d3, 32'h43795048, 32'hc203084f},
  {32'h4442cbd4, 32'hc171fe44, 32'hc2decda5},
  {32'hc4f89e34, 32'hc1b0b7ca, 32'h42e71218},
  {32'h4463037c, 32'h43074646, 32'h430dc569},
  {32'hc4ceee11, 32'hc31ad3e8, 32'h43873acb},
  {32'h44bf85a4, 32'hbd4f0400, 32'hc2982c5f},
  {32'hc4cc8c96, 32'h4368d42e, 32'hc33f7fb7},
  {32'h417998c0, 32'h43a0d4b0, 32'hc37e81e5},
  {32'h439a1d98, 32'h41c6ce00, 32'hc3207d67},
  {32'h42608251, 32'h4380b949, 32'hc2f79273},
  {32'hc4a8c830, 32'hc3bfb1a5, 32'h430ad2f7},
  {32'h44dd864e, 32'h43433468, 32'h43bac8ab},
  {32'hc4f7cd7a, 32'hc1d72f27, 32'h4288ab43},
  {32'h43a9f8d6, 32'hc220ff85, 32'h42c9b0bf},
  {32'hc4338f10, 32'hc39c445c, 32'hc33f2a9f},
  {32'h44c5082f, 32'h43d9e692, 32'hc3864446},
  {32'hc48ab497, 32'hc2789a02, 32'hc29ed078},
  {32'h44ac875e, 32'h42de5e06, 32'h413296e1},
  {32'hc41d8950, 32'h44127ffc, 32'h432a7155},
  {32'h449cf93b, 32'hc28043a5, 32'h4369de1f},
  {32'hc3bf459b, 32'hc3683d9d, 32'h421b2d15},
  {32'h4511ace3, 32'hc33020cd, 32'h43447d14},
  {32'hc4c3c9d7, 32'hc39191d6, 32'hc35c0aba},
  {32'h44b71855, 32'h432b55ad, 32'h42c1a7c5},
  {32'hc450a85a, 32'hc21f3c49, 32'h4266aa2a},
  {32'h44b3a555, 32'h43901b3f, 32'h42a08f45},
  {32'hc48841de, 32'h432099aa, 32'hc3d65de1},
  {32'h4426f8b4, 32'h431a6f01, 32'h432f05d3},
  {32'hc483b614, 32'hc2ba20d3, 32'h43dca3fb},
  {32'h4487a4f4, 32'h4338784c, 32'hc1a97564},
  {32'hc4dad6a3, 32'hc3b1966b, 32'hc3439f82},
  {32'h41198880, 32'h42aae290, 32'hc22df96c},
  {32'hc4d93b03, 32'h434e6e97, 32'h4292e6c9},
  {32'hc2715ca0, 32'h4370ce08, 32'hc31acf49},
  {32'hc42c2418, 32'hc36d3410, 32'hc2dfa591},
  {32'h44a612a2, 32'hc260fddd, 32'h43a65e54},
  {32'hc4e193da, 32'h432c27f9, 32'h440f51a9},
  {32'h44efb4d1, 32'h425ce8a3, 32'h42f63cc3},
  {32'hc51e2ea2, 32'hc35f33ba, 32'hc3a9b962},
  {32'h44bd6dae, 32'h434aa239, 32'hc2b6dc29},
  {32'hc4b8faa0, 32'h41445b80, 32'h4366bccd},
  {32'h42d4e300, 32'hc35e14ce, 32'h43160c66},
  {32'hc482ba60, 32'hc2e17ae1, 32'hc283409c},
  {32'h44e7b40c, 32'h4393efed, 32'hc391389d},
  {32'hc4fc0d48, 32'hc3e06e73, 32'h41c8a095},
  {32'h447c7d2e, 32'hc3291cfa, 32'h431f5cbe},
  {32'hc4c5c388, 32'hbf1bf810, 32'h428578c1},
  {32'h450a3982, 32'hc3948a05, 32'hc321ea45},
  {32'hc4fbcf42, 32'hc29620cb, 32'hc2dc762e},
  {32'h450aadbe, 32'hc2c5a3c5, 32'hc331d9b6},
  {32'hc43c6bc8, 32'hc3a8c8ea, 32'hc28f2b5a},
  {32'h43ea8708, 32'h437bb3df, 32'h4395f12b},
  {32'hc494d79e, 32'h42cc1b1f, 32'h4276f662},
  {32'h441a1fe1, 32'h42cbd2c2, 32'h43218dbc},
  {32'hc384a040, 32'h43672d77, 32'hc3447490},
  {32'h4509cd90, 32'h42a4a1af, 32'h43d077b1},
  {32'hc4026060, 32'h4395ebc6, 32'h4339b80f},
  {32'h4523afc7, 32'hc3572b28, 32'hc242977e},
  {32'hc4c56cec, 32'hc3e30bc9, 32'h43a3e833},
  {32'h450038b2, 32'hc2fdd9ff, 32'hc3138ed5},
  {32'hc3cfa89b, 32'h43979bcf, 32'hc353d286},
  {32'h4481d65c, 32'h43a47a4f, 32'h43aba1dd},
  {32'hc503dc4f, 32'hc38bcc37, 32'h434cef26},
  {32'h44de6bcb, 32'h420fea8f, 32'hc151075c},
  {32'hc4b8de2a, 32'h4385627f, 32'h432d38ca},
  {32'h44ba6c9e, 32'hc341cf8d, 32'h434c0a35},
  {32'hc502f35d, 32'h4231f24d, 32'h4238f863},
  {32'h44deea84, 32'h416462d0, 32'hc0e1b7a5},
  {32'hc2af56c0, 32'h426b0d5a, 32'h43366b13},
  {32'h44686e6e, 32'h433e71b1, 32'h4272fb24},
  {32'hc2cc8bbd, 32'hc312cd15, 32'hc3356548},
  {32'h45020fe3, 32'hc3bb8ff4, 32'h413daffe},
  {32'hc43e4e97, 32'h43c36ef8, 32'hc2a864b1},
  {32'hc32f8928, 32'hc2a2348a, 32'h4269cf5e},
  {32'hc4f97fd5, 32'h4389a0ac, 32'hc1f3f4cb},
  {32'h4389c59f, 32'hc20a2169, 32'h423eec04},
  {32'hc502f5fd, 32'h42016f5b, 32'h43f48647},
  {32'h44b1506e, 32'hc081aaff, 32'hc2724a3f},
  {32'h41aaaf40, 32'h43b5d6d2, 32'h437eb8e4},
  {32'h44d469cc, 32'h4333d003, 32'hc1f9f210},
  {32'hc4fc443b, 32'h434ae4ad, 32'h4357ecd9},
  {32'h4507f578, 32'hc36cf26c, 32'h4306cb80},
  {32'hc4e2a5b5, 32'h432b8bdf, 32'hc335eaca},
  {32'h451c76a2, 32'h4229999b, 32'h437a3670},
  {32'hc42ba3b8, 32'h430a5968, 32'h41ccc2f8},
  {32'h445d3620, 32'h410e4f3b, 32'h430f1d13},
  {32'hc4ea6814, 32'hc3bd9cc5, 32'hc1e38411},
  {32'h44c8a51b, 32'h43b15cf2, 32'h439047be},
  {32'hc506d24a, 32'hc2970cd1, 32'hc271ed8a},
  {32'h434840d0, 32'hc1853c06, 32'h42f94a28},
  {32'hc516c9fe, 32'h430b1705, 32'hc310a254},
  {32'h449e7010, 32'h440f9cd7, 32'hc287f765},
  {32'hc45395ef, 32'hc2c1e75d, 32'h438749cd},
  {32'h439b596c, 32'hc3878ab4, 32'hc24cb0c2},
  {32'hc51aec3c, 32'hc344d73e, 32'h42e3b131},
  {32'h43d9a7d5, 32'hc3a3e57a, 32'hc396993d},
  {32'hc515d362, 32'h42f2a7ae, 32'hc2761a96},
  {32'h4462f33e, 32'h43c1cd8f, 32'h43a56a85},
  {32'hc498e7fd, 32'hc19317e0, 32'hc2a3b8cb},
  {32'h4527276e, 32'hc28498c6, 32'h425e18bd},
  {32'hc4235210, 32'h42477159, 32'hc244621c},
  {32'h44d64ffa, 32'h42ea6caf, 32'hc2d29d76},
  {32'hc48bc11b, 32'h439ab48b, 32'hc29c5ab9},
  {32'h4388dc80, 32'hc1e02b2b, 32'h4343ba12},
  {32'hc4acfdb2, 32'hc302cd7f, 32'hc3f99f16},
  {32'h43a5a20c, 32'h44010efd, 32'h432fa745},
  {32'hc5153472, 32'h4379a0ba, 32'h43124d06},
  {32'h44d8daf6, 32'h412ebd64, 32'hc2bd14da},
  {32'hc4fd4a52, 32'hc371e9b4, 32'hc373acf8},
  {32'h4492c707, 32'hc3b7220c, 32'hc2af83bf},
  {32'hc5201399, 32'hc3019344, 32'hc388f044},
  {32'h44fa1c5f, 32'hc3a09f4c, 32'h43138f9e},
  {32'hc51b5067, 32'h433f522d, 32'h430a5709},
  {32'h450bcfa4, 32'h43b385ed, 32'h4398655b},
  {32'hc38468f8, 32'h43782e1a, 32'hc3a94a49},
  {32'h449bc5d2, 32'hc1fe0abc, 32'hc2befdf7},
  {32'hc4f4a908, 32'hc217f2a7, 32'hc3bfa6e0},
  {32'h4473679c, 32'hc3463729, 32'hc2bce437},
  {32'hc339eb6e, 32'h4372ee95, 32'hc3de8cbe},
  {32'h4502897e, 32'hc329f381, 32'h42f9b038},
  {32'hc3561c20, 32'hc2c2fff6, 32'hc387e1ba},
  {32'h45167cf1, 32'hc3d87ea6, 32'h427df11d},
  {32'h43297179, 32'hc367a6bb, 32'h42b2da75},
  {32'h43fbe9b0, 32'h43817824, 32'h42567504},
  {32'hc450bc5c, 32'h42fdb80a, 32'hc250314c},
  {32'h43c161c0, 32'hc2d47798, 32'hc0d53442},
  {32'hc32783d0, 32'h4294ac2e, 32'h43b30826},
  {32'h450a4878, 32'hc204d95b, 32'hc23628a4},
  {32'hc5068c2a, 32'h42f5a4bb, 32'h43a02915},
  {32'h4517ceea, 32'hc340985f, 32'h4398cc15},
  {32'hc41ec633, 32'hc399db0f, 32'hc2e7d2a6},
  {32'h44f9ff11, 32'hc23e760d, 32'h43ab6080},
  {32'hc3d4c14c, 32'hc30dfcc8, 32'h42845da6},
  {32'h450dff84, 32'hc2f8468c, 32'h414d5bd2},
  {32'hc48e1df2, 32'h42a0ac3a, 32'hc3230fbf},
  {32'h4303091c, 32'hc36d2183, 32'hc23278af},
  {32'hc4ef8af3, 32'hc355b5da, 32'h43167c7e},
  {32'h4445c758, 32'h433474fc, 32'hc391d6ab},
  {32'hc3fc6c72, 32'hc38d5ca5, 32'h435e5a21},
  {32'h42e1d6f4, 32'h43972f9f, 32'h42a60432},
  {32'hc1372800, 32'h42946a1e, 32'hc3a328b1},
  {32'h4486971f, 32'h436fe200, 32'hc374c20e},
  {32'hc4d4838b, 32'hc3820721, 32'h4207a7c5},
  {32'h4493d1c3, 32'hc352fede, 32'h432c5c7c},
  {32'hc5010720, 32'h43afedd9, 32'h43adb140},
  {32'h448bc158, 32'h4317168b, 32'hc42a8979},
  {32'hc46d3568, 32'hc3eccdc7, 32'hc398e73a},
  {32'h4472db60, 32'h41269a42, 32'hc11e201d},
  {32'hc50538d0, 32'hc14cf39b, 32'hc3085555},
  {32'h4349f55c, 32'h428433ed, 32'hc3c6c6ed},
  {32'hc41af410, 32'hc2a31767, 32'h411c4aa4},
  {32'h449cfba4, 32'h422775c6, 32'h42ffd2c4},
  {32'hc4df4f59, 32'hc316aa06, 32'h435b4cdc},
  {32'h435445fc, 32'h437ade25, 32'hc38eb3ab},
  {32'hc4e258a8, 32'hc2800176, 32'h439fe76f},
  {32'h4518f224, 32'hc3889399, 32'h431ab7f2},
  {32'hc48b1f70, 32'h43556d06, 32'h42a6a97c},
  {32'hc2df8d49, 32'h43a627b6, 32'hc2600ab4},
  {32'hc48ce62f, 32'hc395c53f, 32'h409424fe},
  {32'h45063420, 32'hc139b993, 32'hc2c83e2e},
  {32'hc41e1dda, 32'hc2c7b378, 32'h42e30e8b},
  {32'h44abac32, 32'h42b888e6, 32'hc17e3cc6},
  {32'hc44740c7, 32'hc2ccb880, 32'h421bf567},
  {32'h4490c28a, 32'h43844c99, 32'hc3d0965a},
  {32'hc4c20baf, 32'hc3c69822, 32'h43a4457b},
  {32'h450ba35d, 32'hc3862ed5, 32'h42fd8112},
  {32'hc5023252, 32'hc2cc5b80, 32'hc3266795},
  {32'h4511b3e2, 32'h42214e9f, 32'hc36f3b58},
  {32'hc3d504ec, 32'h42f27be2, 32'h4341a988},
  {32'h43bd6c3d, 32'hc3c80794, 32'hc19c741d},
  {32'hc4fb2846, 32'h42cad66f, 32'hc1d488c3},
  {32'h451e800c, 32'h436f1ff7, 32'h43b25132},
  {32'hc46fa6c4, 32'hc4096efb, 32'hc372e20f},
  {32'h448a1b46, 32'h42b2a932, 32'hc3e88eba},
  {32'hc4bf0712, 32'h429c4cc2, 32'h43a8a065},
  {32'h438974e4, 32'h4232c58c, 32'hc28f632d},
  {32'hc43dc11f, 32'hc30b4303, 32'h43867456},
  {32'h438170ad, 32'hc337c674, 32'hc309c871},
  {32'hc466d365, 32'h43a8a772, 32'h43a8d757},
  {32'h44b981f7, 32'h42a7750e, 32'hc351c4bf},
  {32'hc49041e0, 32'h432d86ee, 32'hc30598fc},
  {32'h4438144e, 32'h42d80351, 32'hc30b21b0},
  {32'hc3921e19, 32'h432d3b65, 32'hc2ae2cb0},
  {32'h44cc3ad2, 32'h42f1bb4a, 32'hc325ec14},
  {32'hc484f728, 32'h431e8c93, 32'h43f6d3b4},
  {32'h43fc8090, 32'h4315c650, 32'hc446123c},
  {32'hc40e632b, 32'hc3c7f833, 32'h4330cecf},
  {32'h42a24530, 32'hc31c3874, 32'h42bd9fcb},
  {32'hc51262f9, 32'h410b84cd, 32'h434eca5e},
  {32'h450aa494, 32'hc3a5c516, 32'hc39edb76},
  {32'hc44d9f59, 32'hc28d2d11, 32'h438c6788},
  {32'h45050773, 32'h41a97ea6, 32'h4352b3e5},
  {32'h42da34e0, 32'hc1d8f643, 32'h41c6a3e6},
  {32'hc4e0483f, 32'h4333fda7, 32'hc404f983},
  {32'h43cbd54a, 32'hc3a45f82, 32'h439be3d9},
  {32'hc4925e53, 32'hc2dbe3c1, 32'h435c82c9},
  {32'h43215398, 32'hc391cf51, 32'hc278165f},
  {32'hc49d7b83, 32'h42fc8e13, 32'h42b1125a},
  {32'h446bebec, 32'hc304e662, 32'hc3bf51fe},
  {32'hc4f3d71d, 32'hc3094780, 32'h438869a1},
  {32'h443489a6, 32'hc08d1273, 32'hc32e6895},
  {32'hc3b4c588, 32'hc14201d6, 32'hc40bf3ae},
  {32'h44f672ce, 32'h43a356cd, 32'hc2d3c37d},
  {32'hc3e08674, 32'hc3a9f0b7, 32'h42336458},
  {32'h44b4bce2, 32'hc38ac454, 32'hc3baef0d},
  {32'hc4d59c93, 32'hc2289cd8, 32'h42c608e8},
  {32'h4505b3c8, 32'hc13ac7c2, 32'h430746ae},
  {32'hc2d59ad0, 32'hc324ef3e, 32'hc2bbb17a},
  {32'h450ae4f9, 32'h439064f8, 32'hc3ba8d64},
  {32'hc417e06d, 32'hc1d00dae, 32'h43296123},
  {32'h44e3c7ac, 32'hc2119cf9, 32'h42d1652d},
  {32'hc3aebf07, 32'h438961aa, 32'hc299b9ab},
  {32'h4405c3c0, 32'h43052cf6, 32'h42855564},
  {32'hc41c8ed0, 32'h4381f401, 32'hc296ed49},
  {32'h43c89a19, 32'hc33960c0, 32'hc3827eee},
  {32'hc4095a59, 32'h4306bb63, 32'h42f115a3},
  {32'h45055804, 32'h4289f1ee, 32'hc336763b},
  {32'hc4d1c12a, 32'hc1028440, 32'h435f8778},
  {32'h44d0938f, 32'h436771bc, 32'hc2968c54},
  {32'hc3b9a572, 32'h440489db, 32'h42df4c38},
  {32'h44315356, 32'h43baa5f0, 32'h4332052e},
  {32'hc5026c95, 32'hc347dec2, 32'hc340c5ca},
  {32'h44e5ea89, 32'h42ea3189, 32'hc28433d8},
  {32'hc4ab0141, 32'h4318a708, 32'hc2adc20c},
  {32'h43b555e8, 32'h431d9027, 32'hc2f6e9b7},
  {32'hc43810ba, 32'hc33b7264, 32'h41cc2e7a},
  {32'h433b9120, 32'hc31fefa9, 32'hc32f3e67},
  {32'hc498bf79, 32'hc1ebb2aa, 32'hc1c8f98d},
  {32'h445a403e, 32'hc3902390, 32'hc2df11cf},
  {32'hc3a6c590, 32'hc2ac63d6, 32'h429aadca},
  {32'h436d5910, 32'h4217ab26, 32'h425be5cb},
  {32'hc417e398, 32'hc374ffda, 32'hc3dac7e0},
  {32'h44dddb94, 32'hc441c587, 32'hc2c130bd},
  {32'hc3a41e80, 32'hc34bb5c7, 32'h4342cb86},
  {32'h445f345a, 32'h430fb9bc, 32'hc08f09f0},
  {32'hc491cbf9, 32'hc3ab185f, 32'hc2e0aca0},
  {32'h44461e6a, 32'hc30c03e3, 32'h423bd096},
  {32'h430e022e, 32'hc3999cbb, 32'hc14370a5},
  {32'h450bf76a, 32'h4333718c, 32'hbe575a30},
  {32'hc3d08a1c, 32'h42f67b67, 32'hc376024a},
  {32'h43fd6c2d, 32'h4432bde1, 32'hc212fae5},
  {32'hc4cc1d32, 32'h41573ee8, 32'hc374191b},
  {32'h44f3eda2, 32'hc30e06ac, 32'hc2aa4c47},
  {32'hc4f63a4b, 32'hc3809980, 32'hc22957ab},
  {32'h44df5499, 32'hc3096fa1, 32'h4223e164},
  {32'hc41a3878, 32'h41999eea, 32'hc2b46fd2},
  {32'h44d01f9b, 32'hc3680f0c, 32'hc3d7c208},
  {32'hc36a2655, 32'hc2da41c4, 32'hc2ea4c0a},
  {32'h44e2fbe7, 32'hc379506e, 32'hc396f535},
  {32'hc3a18c14, 32'hc2c8711f, 32'hc30a16b1},
  {32'h44848a56, 32'hc3cd15be, 32'h4217e246},
  {32'hc4d6b21e, 32'hc16f6d36, 32'hc33258c6},
  {32'h44f45940, 32'hc3e89b0c, 32'h42d1eaac},
  {32'hc385259b, 32'hc3700334, 32'hc302e6e1},
  {32'h44eebc68, 32'h43b01f05, 32'hc342f847},
  {32'hc512be16, 32'hc21f12dc, 32'hc2bd003c},
  {32'h431ad990, 32'hc2d08526, 32'h41c9d089},
  {32'hc417d442, 32'hc30d50a7, 32'h4432903b},
  {32'h441d2138, 32'h433992c5, 32'hc406a44d},
  {32'hc4f5737d, 32'hc3cfd247, 32'h4254a9bf},
  {32'h44a2e898, 32'h42b2d522, 32'h43c467b8},
  {32'h430f8a48, 32'hc2c8b7f4, 32'h4312881e},
  {32'h44cb8c0f, 32'hc3bacfe2, 32'h42f67a0b},
  {32'hc48ee8c3, 32'h4282e820, 32'hc12f176e},
  {32'h44394737, 32'hc4174c50, 32'h4338de60},
  {32'hc4e4fba4, 32'h43a2dc0d, 32'h426f3a32},
  {32'h44e7b2fa, 32'hc1f5871a, 32'hc36c6de2},
  {32'hc45100e6, 32'h41f7ca02, 32'h43233c3d},
  {32'h44b8a7e4, 32'h41c67366, 32'hc2a0f81f},
  {32'hc3afd620, 32'h4384a314, 32'hc40a0515},
  {32'h4481636a, 32'hc26663c8, 32'h43e815f3},
  {32'hc4e9605e, 32'hc259d196, 32'hc1f528b0},
  {32'h424f54a8, 32'hc36faf44, 32'h43820e8c},
  {32'hc35c8430, 32'hc23b2329, 32'h438dd37a},
  {32'h44956b49, 32'h41796bee, 32'h43351e75},
  {32'hc424cf84, 32'hc2286f01, 32'h435ecef2},
  {32'h451ee152, 32'h431a48ee, 32'h431716a6},
  {32'hc51236e7, 32'hc3066ed7, 32'hc32331ea},
  {32'h445a013c, 32'hc20a2e30, 32'hc32520b9},
  {32'hc45013b5, 32'hc311b917, 32'h41b2f3c9},
  {32'h44570156, 32'hc306deb4, 32'h43153917},
  {32'hc48a7868, 32'hc38e1d15, 32'hc36ec661},
  {32'h4413c974, 32'hc36a1bb7, 32'hc382b4d8},
  {32'hc486ab29, 32'hc383735a, 32'hc1905a7a},
  {32'h441f11c0, 32'hc2f86d0e, 32'h4325ac2d},
  {32'hc50667e8, 32'hc32933fb, 32'hc3b1d56b},
  {32'h45064a1c, 32'hc3a80757, 32'h43815cbd},
  {32'hc2dc4364, 32'h42418dfb, 32'h4327f9ca},
  {32'h4492e911, 32'hc3623328, 32'hbf77437b},
  {32'hc390bae8, 32'h42b3e2e3, 32'h43452d56},
  {32'h44801889, 32'hc33d05a2, 32'hc316dc32},
  {32'hc3e3861e, 32'h42c06088, 32'hc302a31a},
  {32'h44a2e0fb, 32'hc1d69ea6, 32'hc214a119},
  {32'hc4a66596, 32'h437481c5, 32'hc2295dea},
  {32'h43649450, 32'h432d5f43, 32'h4388997a},
  {32'hc4eec445, 32'hc24b5d68, 32'h434d8218},
  {32'h43f601f8, 32'hc304be6a, 32'h437aa004},
  {32'hc484a9ac, 32'h428364dc, 32'h42e89a0d},
  {32'h44a873a3, 32'hbef63773, 32'h42b7d831},
  {32'hc5068574, 32'hc2980f90, 32'hc3877dcd},
  {32'h44d85d6c, 32'hc374ba9a, 32'hc27bbb32},
  {32'hc44bea84, 32'h43f33a9a, 32'h43642a23},
  {32'h44f39416, 32'h43959157, 32'h3c20a000},
  {32'hc2f1c0d0, 32'h41d0da38, 32'h431a9ed1},
  {32'h4502a3f6, 32'hc2908ef5, 32'h42e154e5},
  {32'hc4c0e2dc, 32'hc2b29630, 32'h43a3b6f4},
  {32'h437c2430, 32'h431ad0db, 32'h427333aa},
  {32'hc3c6d088, 32'h432ef372, 32'hc394ce90},
  {32'h439271a8, 32'h4399a10c, 32'h41a1d42a},
  {32'hc350d664, 32'h43c28e84, 32'hc3bdc1f5},
  {32'h448b2e6b, 32'hc29eefa6, 32'h4208a210},
  {32'hc394b8e7, 32'hc392b36f, 32'h41278d6a},
  {32'h4492972e, 32'hc2c596d2, 32'h428ac3e8},
  {32'hc44c93d1, 32'hc1772f7f, 32'hc3bb0e27},
  {32'h4448a841, 32'hc10f4fee, 32'h43381793},
  {32'hc4bc57f0, 32'hc2d64b5f, 32'hc2ef653f},
  {32'h45051176, 32'h43c3ff3d, 32'hc23cc529},
  {32'hc4642149, 32'h43f4c443, 32'hc2e3f4a9},
  {32'h44ee0fd8, 32'hc27cb8d0, 32'hc323dab5},
  {32'hc4c831c0, 32'h42ca28ac, 32'hc2bf1e5f},
  {32'h44f7d52f, 32'hc35c21e7, 32'h414799b2},
  {32'hc444ad3a, 32'h432da5c6, 32'h43e181c8},
  {32'h43a5d878, 32'hc32385a8, 32'h4379b2e5},
  {32'hc46e5243, 32'hc38b07f2, 32'h432345f7},
  {32'h44cbd7ce, 32'h43be9adb, 32'hc1ad7466},
  {32'hc4f9cada, 32'h439cf674, 32'h4310b7be},
  {32'h43df828a, 32'hc2480d4d, 32'h431098b8},
  {32'hc37c7b20, 32'hc343024d, 32'hc17de35d},
  {32'h44b2f8e0, 32'h4331acf8, 32'h43502d58},
  {32'hc473ce00, 32'hc2901732, 32'hc2bc7c66},
  {32'h449d1bfa, 32'h43b06739, 32'hc2a69f03},
  {32'hc28a3100, 32'h4324654e, 32'hc3954900},
  {32'h44b42e0b, 32'hc382dc77, 32'hc39ed935},
  {32'hc48fe7b8, 32'hc21d4c7a, 32'hc385a95b},
  {32'h4512b389, 32'hc3890de3, 32'h42ed9811},
  {32'hc3746ec4, 32'h43cd7599, 32'hc2169868},
  {32'h44d30871, 32'h42edc38f, 32'h41f92cf3},
  {32'hc4f2a385, 32'hc2790060, 32'h42a8b068},
  {32'h44d68891, 32'h43696f44, 32'h428792eb},
  {32'hc4e985e2, 32'h4313033d, 32'h43846570},
  {32'h446e9ec3, 32'h43044f7a, 32'hc392498e},
  {32'hc5057881, 32'h429e8288, 32'h43958ac8},
  {32'h44e93a49, 32'h42d0509e, 32'h42b1df5e},
  {32'hc3f105b6, 32'hc384facc, 32'h42d80b01},
  {32'h43361c3b, 32'h4052540d, 32'hc2c841aa},
  {32'hc41bbbec, 32'h43295aaf, 32'hc38836dc},
  {32'h4510dbaa, 32'h42a1111c, 32'hc35ce7c3},
  {32'hc3858a70, 32'h4323e7e0, 32'h43ffcdca},
  {32'h45102d8a, 32'hc16e2dfc, 32'hc4008e99},
  {32'hc516a501, 32'h435bd06a, 32'hc34a9fd0},
  {32'hc15d46c0, 32'hc20c1f07, 32'hc37ae9ca},
  {32'hc4ea8bed, 32'hc28b4461, 32'h439c0dca},
  {32'h4519a9e2, 32'h439a36e5, 32'h4313ed92},
  {32'hc4af10aa, 32'hc2ee8b42, 32'h43aae70e},
  {32'h443c236f, 32'h42899195, 32'h40f620dd},
  {32'hc501d00c, 32'h4231bf91, 32'hc2100d3d},
  {32'h44a1b461, 32'hc2307ddc, 32'hc38c8b09},
  {32'hc4e779e2, 32'hc3778cc6, 32'h434ae331},
  {32'h4494112e, 32'h43452f7e, 32'hc36f777b},
  {32'hc3da6fa0, 32'hc388db12, 32'h42dfb3fe},
  {32'h44c7ca2b, 32'h42637edb, 32'hc3aba0e9},
  {32'hc4a88d96, 32'h437df06c, 32'hc2b2ee49},
  {32'h439c9860, 32'hc3641b80, 32'h4387d78a},
  {32'hc3ef3488, 32'hc3126bb5, 32'h440dbb20},
  {32'h44bf8e60, 32'hc3efdd19, 32'hc3975e9e},
  {32'hc454c735, 32'hc3902817, 32'hc23b0623},
  {32'h43f76812, 32'h433607d3, 32'h4171199a},
  {32'hc50d0ef5, 32'hc2b4eef6, 32'hc34a0949},
  {32'h45088ce4, 32'hc31764f4, 32'hc36b022d},
  {32'hc195ea80, 32'hc354c767, 32'h436571de},
  {32'h43954ae6, 32'h40c2e405, 32'hc31682e2},
  {32'hc49eb16e, 32'hc3f96228, 32'hc37ca441},
  {32'h4411db9c, 32'hc3af083a, 32'hc20caf25},
  {32'h42649b40, 32'hc2ddde18, 32'hc1b63324},
  {32'h447fcaae, 32'h4322cee1, 32'h43459089},
  {32'hc49015be, 32'h43001aa4, 32'h411ae2d3},
  {32'h44d7cc38, 32'hc2659198, 32'hc26c9e5b},
  {32'hc4ae2548, 32'h4398aea1, 32'h42a96578},
  {32'h44224d3c, 32'h427cc191, 32'hc3c363d7},
  {32'hc5156dca, 32'h41adc272, 32'hc3a8b87a},
  {32'h43454db9, 32'h42fab490, 32'hc35063c9},
  {32'hc49a7fe4, 32'h42571646, 32'hc359e72c},
  {32'h44a73332, 32'h428a2bf2, 32'hc3647270},
  {32'hc4f3b13f, 32'h437818e4, 32'h43232365},
  {32'h4515f5e4, 32'hc3252577, 32'hc3b51a7d},
  {32'hc4fbebb4, 32'h425b1924, 32'hc049483a},
  {32'h45072581, 32'h43557e40, 32'h438e1351},
  {32'hc4a0eb9a, 32'h4215649e, 32'h4282c417},
  {32'h4511b013, 32'h432a6c0c, 32'h441ea00f},
  {32'hc4a83d26, 32'h43864b94, 32'h42f1f7fb},
  {32'h43d004ba, 32'h43ae8211, 32'hc3aac660},
  {32'hc40bc1da, 32'hc396d813, 32'h43926c42},
  {32'h4345a288, 32'h425c93ca, 32'h428476d0},
  {32'hc4ed8236, 32'h42c887ba, 32'hc2c97485},
  {32'h44afb98c, 32'hc420ca25, 32'h4323da71},
  {32'hc3ce0956, 32'hc2d8020b, 32'h43bd3d7b},
  {32'h43fd823a, 32'hc38ffcbf, 32'hc2902d09},
  {32'hc4c9b1b9, 32'h42359f38, 32'hc188e2cd},
  {32'h440ebd99, 32'h43a59bba, 32'h416497ef},
  {32'h41308500, 32'h41d93be1, 32'hc34c5d60},
  {32'h44a62491, 32'hc27f602b, 32'h4329f346},
  {32'hc41f6e48, 32'h439d6a5b, 32'h4365ae19},
  {32'h4516f617, 32'hc34dcfc8, 32'hc36077fa},
  {32'hc41df380, 32'hc3534da0, 32'h433379c7},
  {32'h44676cf3, 32'h429a38c8, 32'h42793e17},
  {32'hc4b47437, 32'hbeda5842, 32'h43f3f8b6},
  {32'h44f9b571, 32'h43465b59, 32'hc302e7aa},
  {32'h40ae1365, 32'h4307848c, 32'h42ab1f74},
  {32'h44a6ea09, 32'h4354fb68, 32'hc2c6405d},
  {32'hc4256ffa, 32'hc28fbd11, 32'hc2b9b532},
  {32'h449cc0c1, 32'hc35c6196, 32'hc28c2874},
  {32'h42e23dc8, 32'h43cf2732, 32'h438db5dd},
  {32'h4418d72e, 32'h4350afe2, 32'h42f84e1d},
  {32'hc4c48133, 32'h4398a4f7, 32'hc2937af2},
  {32'h45020fcf, 32'h43ad757d, 32'h42e8bc91},
  {32'hc4e78ee3, 32'hc252e6da, 32'h43012c64},
  {32'h442ae4a6, 32'h42de2e7f, 32'hc344400b},
  {32'hc424b9b3, 32'hc3f11e32, 32'hc3a3c4d6},
  {32'h450fad5b, 32'h435558aa, 32'h42f7218a},
  {32'hc4d2a535, 32'h42a12253, 32'hc2e1de1e},
  {32'h44aae836, 32'h42c87d54, 32'hc319b6ab},
  {32'hc4e81b00, 32'h4194627f, 32'hc398cc9b},
  {32'h450d43db, 32'h431039ac, 32'hc31bdc9b},
  {32'hc3eb0892, 32'h423e9c18, 32'hc3389f2e},
  {32'h43b8881c, 32'h42af695d, 32'h42c3a371},
  {32'hc4e0fd52, 32'hc2409188, 32'h438dc8b8},
  {32'h43939143, 32'h436b08a7, 32'h43651228},
  {32'hc419836b, 32'hc2f02493, 32'hc3a72339},
  {32'h44eacd07, 32'hc349ef55, 32'h438d0328},
  {32'hc4f8c903, 32'h4264b118, 32'h43754389},
  {32'h43171e20, 32'hc2ae52a5, 32'hc33c6b4a},
  {32'hc4a1cd48, 32'hc14a5cae, 32'hc3a587e7},
  {32'h44e395ee, 32'h42193ab0, 32'h41f9a65a},
  {32'hc4a406e5, 32'hc34bacb0, 32'h429d8294},
  {32'h44cb351e, 32'hc209222b, 32'h43584e24},
  {32'hc4b8bb76, 32'hc20adea8, 32'h43831f85},
  {32'h450448d6, 32'h42c573df, 32'hc28e31d6},
  {32'hc4610ace, 32'hbf6fc634, 32'hc1d54eed},
  {32'h43eb2a8f, 32'hc34b566c, 32'hc11746c4},
  {32'hc42ea438, 32'h4232d698, 32'h43c162ec},
  {32'h43bb72f8, 32'h439adba3, 32'hc0942a47},
  {32'hc491f5b3, 32'hc3280885, 32'hc2cfce40},
  {32'h44f9fae4, 32'h428fed09, 32'h402c9ab0},
  {32'hc4752a34, 32'h439e52c6, 32'hc2041662},
  {32'h43b3931c, 32'hc3dae66c, 32'hc34854d8},
  {32'hc4a9efd2, 32'hc2f97c3a, 32'hc2287268},
  {32'h44f5e9d0, 32'h4358d3b0, 32'hc36977cd},
  {32'hc41422be, 32'h434b09c1, 32'h431b1cd4},
  {32'h447986d8, 32'h43a301fb, 32'h4383b875},
  {32'hc412476e, 32'h435c2310, 32'h435817d2},
  {32'h43d06b70, 32'hc3f47387, 32'h43863100},
  {32'hc2937823, 32'hc384fa66, 32'h43334bba},
  {32'h44c5ee43, 32'hc2f46091, 32'h412d784d},
  {32'hc5004dac, 32'h42c62ed6, 32'hc3b18aba},
  {32'h4519adf0, 32'h430479d4, 32'h43ee3d6e},
  {32'hc4fb4ed7, 32'hc24d9790, 32'hc2998dae},
  {32'h4320bea7, 32'h43f3e956, 32'hc3f7e4f0},
  {32'hc4b34eae, 32'h43a14a13, 32'h42cb8f57},
  {32'h440861cc, 32'hc37b9974, 32'hc2bf3f29},
  {32'hc38b19fc, 32'h431cf2a3, 32'h43ac841d},
  {32'h44984d9c, 32'h43981692, 32'hc415b4a1},
  {32'hc4aefe56, 32'hc1adbdec, 32'hc26f7fe7},
  {32'h450e3094, 32'h42af209f, 32'hc2172ef2},
  {32'hc41db66c, 32'h428c05fd, 32'h4244e778},
  {32'h446c65b0, 32'h4345a040, 32'hc1d84397},
  {32'hc3ebd794, 32'hc3a7b28d, 32'hc26fc6c5},
  {32'h44a33a11, 32'hc3aeb67b, 32'h434fcc4a},
  {32'hc503f10c, 32'h432c65b7, 32'h42fbd754},
  {32'h44f617b3, 32'h431cecf0, 32'hc3c4c841},
  {32'hc4bc7654, 32'hc16246e8, 32'h411e763e},
  {32'h44b6db1b, 32'hc2c10fc8, 32'h426dfa5d},
  {32'hc47ec31a, 32'h43d46e8d, 32'h42e02094},
  {32'h44f5955b, 32'h43cceadf, 32'h40b5c402},
  {32'hc50c1889, 32'hc3734c62, 32'hc358e544},
  {32'h448c63af, 32'h438e443f, 32'h42e98507},
  {32'hc3c42400, 32'hc3443cfd, 32'h437e7ad0},
  {32'h424996e8, 32'h43477809, 32'hc259c4e9},
  {32'hc441c3c6, 32'h439f8658, 32'h4332ddfa},
  {32'h43decdfc, 32'hc2d8b91b, 32'h42a8a55b},
  {32'hc4086106, 32'h423829b6, 32'h40845e4a},
  {32'h442b875b, 32'hc3246df8, 32'hc36a8e3f},
  {32'hc4fb8443, 32'hc2b87b52, 32'hc39088fa},
  {32'h43d400c2, 32'hc35b2e2b, 32'hc3ca5251},
  {32'hc4bc662b, 32'hc399ae53, 32'hc1c56514},
  {32'h43b346b5, 32'h42145b35, 32'hc37670ac},
  {32'hc48b7515, 32'h42640465, 32'hc0eb43ed},
  {32'h44e1c75b, 32'h42d5f7cf, 32'hc308dbb2},
  {32'hc4e2da48, 32'h43099ec4, 32'hc24e640c},
  {32'h451723ce, 32'hc329fb9c, 32'h439de6f4},
  {32'hc283d7e0, 32'h42f61436, 32'h43527478},
  {32'h446e80ee, 32'hc10fa61c, 32'h43545fd0},
  {32'hc4e41b3c, 32'h42ae7ac7, 32'h41f15cc1},
  {32'h444c8e77, 32'h4293fea0, 32'hc3fd544d},
  {32'hc4f94cea, 32'hc369f162, 32'h4357fb24},
  {32'h44ad712f, 32'h42cc8125, 32'h42a0f542},
  {32'hc3d6c9dc, 32'h41c6d7aa, 32'h4391e1a5},
  {32'h450d067e, 32'h40e36cac, 32'hc3080418},
  {32'hc52155ca, 32'hc38a289c, 32'h430717ad},
  {32'h412a9f80, 32'h43abc4a1, 32'h42b5df3a},
  {32'hc4ffe71c, 32'h431e11a1, 32'h43762e38},
  {32'h44d1c709, 32'hc368d8d6, 32'h4310327b},
  {32'hc4781834, 32'h42b62c90, 32'h4280f852},
  {32'h4432331d, 32'hc32fe869, 32'h43cdf856},
  {32'hc1a69020, 32'h427edff1, 32'hc29054e2},
  {32'h43faeade, 32'h4281a51c, 32'h435b2010},
  {32'hc506d6ec, 32'hbfbde540, 32'h43441e92},
  {32'h4420c518, 32'h42b534c0, 32'hc2d31c68},
  {32'hc42102b8, 32'hc3b00cf3, 32'h43412156},
  {32'h43acbc0c, 32'h4218552a, 32'hc35c9614},
  {32'hc50a0af0, 32'hc2c32af8, 32'h4302f7ab},
  {32'h440d93c4, 32'hc2e62240, 32'h436e0981},
  {32'hc4c02fa4, 32'h42b9f565, 32'h4341abfc},
  {32'h45072ca6, 32'hc2ab60bd, 32'hc36b02c8},
  {32'hc4b70f92, 32'h43d5d90d, 32'h43b5c1f4},
  {32'h44a313ef, 32'h43c4f997, 32'h4302b0c6},
  {32'hc38a31aa, 32'hc2b81ffd, 32'hc2a9fb78},
  {32'h44d9b21e, 32'h435e2985, 32'h4326e710},
  {32'hc47836c8, 32'hc2422dc2, 32'hc31903de},
  {32'h44c85521, 32'hc3a9324c, 32'h42630abe},
  {32'hc509fe52, 32'hc395f20d, 32'h433870a1},
  {32'h441c4a2a, 32'hc3ce9cb9, 32'hc185eb5c},
  {32'hc4cdb1ce, 32'h4340fe3a, 32'h4319dd67},
  {32'hc26d78c0, 32'h40b72fc8, 32'hc395825c},
  {32'hc510ce45, 32'hc2dfec99, 32'hc3aa073b},
  {32'h44f55e50, 32'h4257fd1e, 32'hc36e76b6},
  {32'hc457abb4, 32'h430c601f, 32'h433b5463},
  {32'h44c25c66, 32'h43b63482, 32'h42712633},
  {32'hc490644b, 32'hc25c2267, 32'hc39252d7},
  {32'h44356712, 32'hc2a07641, 32'hc323e3de},
  {32'hc3b234ec, 32'hc3506966, 32'hc3be4e04},
  {32'h450bef56, 32'h41388008, 32'h42ae2cad},
  {32'hc4aae658, 32'h43081b86, 32'hc0145420},
  {32'h445252b2, 32'h428e35c1, 32'hc30f130b},
  {32'hc49d3313, 32'h438e3b01, 32'hc1baf50d},
  {32'h44dc0598, 32'h439aac59, 32'h42bf9ab5},
  {32'hc4498b4a, 32'hc3040e1b, 32'hc32a98c6},
  {32'h44d01d80, 32'h430e1bca, 32'hc2d3e830},
  {32'hc147f700, 32'h4304010b, 32'h41bec0d4},
  {32'h450295f1, 32'h4342c946, 32'hc36d7bd3},
  {32'hc4ffdb9e, 32'hc272a76d, 32'hc2e39c66},
  {32'h42140a38, 32'hc281634f, 32'hc1a1a584},
  {32'hc48cb2e5, 32'hc2423297, 32'h4384b0d1},
  {32'h44c26a97, 32'hc2928e9b, 32'h431acb0b},
  {32'hc4b415e0, 32'hc2b6123a, 32'hc184c357},
  {32'hc1c44120, 32'hc23e0363, 32'h42e1e543},
  {32'hc2c58b40, 32'h43d29f6f, 32'h44031374},
  {32'h44ee5590, 32'hc406ea79, 32'hc3d401d7},
  {32'hc485a032, 32'h42e28228, 32'h42c0b673},
  {32'h45097a36, 32'h43390bc1, 32'h439244bd},
  {32'hc4a40da4, 32'h42dffb81, 32'hc3728919},
  {32'h44b76a37, 32'h433c75e1, 32'h42d706b9},
  {32'hc4f1f3c8, 32'hc30b5681, 32'hc33c39a2},
  {32'h44b6ace5, 32'h42699dbe, 32'h42c44843},
  {32'hc4e72b84, 32'hc397e7ad, 32'hc24a24a8},
  {32'h4516cd2d, 32'h43712959, 32'h439d90db},
  {32'hc49f3b5a, 32'h435874e0, 32'h43f711c7},
  {32'h436d10e8, 32'h42b9fba4, 32'hc3943566},
  {32'hc4ebdb89, 32'h42b80ef6, 32'h42a71136},
  {32'h44f3843a, 32'hc20635ee, 32'h434f7bf4},
  {32'hc4c593e8, 32'h4364d124, 32'h4253663d},
  {32'h451599d3, 32'h43939819, 32'h43bb287a},
  {32'hc4aef493, 32'hc191b48a, 32'h427422be},
  {32'h45029eff, 32'h3fb697dc, 32'hc35ef028},
  {32'hc4a5554e, 32'hc33a9c28, 32'hc3101b9f},
  {32'h44d8737e, 32'hc3cbbd16, 32'h42b9c48c},
  {32'hc381bc28, 32'hc0223ba6, 32'hc1bc291f},
  {32'h4391c4c0, 32'h432d6da9, 32'hc1e5d44e},
  {32'hc4127afe, 32'h438ac14d, 32'hc2ee2bd0},
  {32'h446d54d8, 32'hc2f272e8, 32'hc2ad7daf},
  {32'hc504f7a4, 32'hc23333d0, 32'hc3246ca3},
  {32'hc212fbc0, 32'h417094b3, 32'h42c28366},
  {32'hc3b61d76, 32'h43de67e2, 32'h42f7c9d7},
  {32'h4514ea92, 32'h43cb49cb, 32'h4397e354},
  {32'hc4e4f722, 32'h43c9890a, 32'hc3a2e74b},
  {32'h44338c4e, 32'hc29247cd, 32'hc261f2f5},
  {32'hc5051276, 32'h43b9c739, 32'h43dd6c5f},
  {32'h44b30504, 32'hc2d58a70, 32'hc270a615},
  {32'hc484160e, 32'hc21c4626, 32'hc3abc1d4},
  {32'h43ea53b8, 32'hc20f3d08, 32'hc1d3c5bb},
  {32'hc5074135, 32'hc3680aab, 32'h43806c5f},
  {32'h44a6473e, 32'h424e50cd, 32'hc39608af},
  {32'hc4cb53d4, 32'h42cde399, 32'hc3098588},
  {32'h4515beb0, 32'hc229a46e, 32'h4365598e},
  {32'hc503d171, 32'h41845c21, 32'hc2975140},
  {32'h4275af40, 32'h426b9e04, 32'hc37a3e8c},
  {32'hc45001a1, 32'hc3e0ec85, 32'h4408404a},
  {32'h4410afa4, 32'h414eeb1e, 32'hc31ab1c3},
  {32'hc3e35dd1, 32'hc3ab1cf0, 32'hc21eebf5},
  {32'h44ce88a6, 32'hc32689cf, 32'h4339fe6d},
  {32'hc5261d2d, 32'h42e6fbc4, 32'h439cf50e},
  {32'h44ed5372, 32'hc346dc94, 32'h42468b7e},
  {32'hc4ef9f94, 32'hc2d96b25, 32'hc3906b00},
  {32'h4496feef, 32'hc306739a, 32'h437f9eb3},
  {32'h420ebbc0, 32'h42651c74, 32'hc28dbf5c},
  {32'h445a6a74, 32'h41cd5acb, 32'hc40fd8d2},
  {32'hc4c5da38, 32'h4216e2be, 32'h4226541a},
  {32'h448ace22, 32'hc2c8a5c6, 32'hc21257c0},
  {32'h4381adc5, 32'h43a36d44, 32'hc399ab78},
  {32'h45221b7a, 32'h4398e1d2, 32'h431a9a87},
  {32'hc4f0e74a, 32'hc33ca29e, 32'hc368f26e},
  {32'h43f37c4f, 32'h4331a1b9, 32'h43bad8cf},
  {32'hc39ee520, 32'h43ba8daa, 32'hc2ce4b90},
  {32'h44f8f56a, 32'h430ea8aa, 32'hc382c481},
  {32'h4391ad30, 32'h42f485a3, 32'hc2e2b36d},
  {32'h44a4ae4d, 32'h4308bc0e, 32'hc37dd7cc},
  {32'h43a43a48, 32'hc3afb174, 32'hc399f533},
  {32'h445aeccf, 32'h43b7a4a7, 32'h43e61b7b},
  {32'hc45ab970, 32'h4350c0ac, 32'h43754302},
  {32'h4413845a, 32'hc3b2f570, 32'h43a4058e},
  {32'hc4b03fa5, 32'h42f1ef94, 32'h429fd861},
  {32'h4513209d, 32'hc2a70514, 32'hc3bbce69},
  {32'hc4be3187, 32'hc1f34cdb, 32'hc292a4e7},
  {32'h44fd4ddd, 32'h43561440, 32'h429659aa},
  {32'hc3ee9aac, 32'h43d3004d, 32'hc398ddd3},
  {32'h4489d654, 32'hc32d0163, 32'hc2a00034},
  {32'hc3bde74c, 32'h428d9dde, 32'hc3853c0f},
  {32'h44fd7098, 32'h43650993, 32'hc184d6de},
  {32'hc4ba87ca, 32'hc2926690, 32'h41d07f52},
  {32'h4328d6f0, 32'h43790192, 32'hc395186d},
  {32'hc3cdd2da, 32'hc29aa10f, 32'h4382203e},
  {32'h44857493, 32'hc1d5ea02, 32'h42d005ea},
  {32'hc4b7984b, 32'hc2faeaec, 32'h42dd46f6},
  {32'h44fa355b, 32'h422392c9, 32'h435480a2},
  {32'hc477780c, 32'hc2e1d88c, 32'h43b9b91a},
  {32'hc5076636, 32'hc36f15ab, 32'hc2e7f9e1},
  {32'h450c1267, 32'h435ce79a, 32'h432ee56d},
  {32'hc4f4d7a7, 32'h430d23c1, 32'hc26a08ac},
  {32'h44198db2, 32'h42981fa0, 32'h437e1da8},
  {32'hc4f4be33, 32'h43b545f9, 32'hc2acd177},
  {32'h4494144a, 32'h42a0063e, 32'h43621d20},
  {32'hc51455fd, 32'hc3407d69, 32'hc35c769f},
  {32'h44dcd23e, 32'h42de91b2, 32'h435114ac},
  {32'hc5073bb8, 32'h437d0602, 32'hc326f3e0},
  {32'h4510546c, 32'hc372b159, 32'hc2a6c1ac},
  {32'hc4cf9a69, 32'h433085a7, 32'hc3cd539c},
  {32'h450b611a, 32'hc3341fd4, 32'h43d2878f},
  {32'hc5175f56, 32'h424644ea, 32'h433ba5cd},
  {32'h444d6ef8, 32'hc31cf932, 32'h43d1d3e3},
  {32'hc44c1b37, 32'hc4022562, 32'hc27eda3a},
  {32'h44f2bf8e, 32'hc2d6cd58, 32'h42686cc8},
  {32'hc4d6e06c, 32'h43836c19, 32'h42533e49},
  {32'h44165336, 32'hc30f7223, 32'h432858af},
  {32'hc504bba2, 32'h435bcaea, 32'h41ee8e04},
  {32'h44157fe4, 32'hc295d868, 32'hc2d1fb6c},
  {32'hc3f213e8, 32'hc22d0b3e, 32'hc39a3c64},
  {32'h444544b2, 32'hc34ae9f1, 32'h420a0a66},
  {32'hc5028210, 32'hc22c3c92, 32'hc3e0a209},
  {32'h44aeb43e, 32'h43f616d1, 32'h43336e91},
  {32'hc494f7fe, 32'hc3a05f6d, 32'hc3a76a15},
  {32'h44c6d8a6, 32'h427d436e, 32'h439387c6},
  {32'hc3baf5be, 32'h43aed708, 32'h42abec3a},
  {32'h44a669da, 32'hc2dffd0a, 32'h4367483b},
  {32'hc4c88df7, 32'hc2057f55, 32'hc41b7a57},
  {32'h43b86b5a, 32'h42b12d98, 32'h424e252a},
  {32'hc4d3503f, 32'h439fcd44, 32'h43d2a64f},
  {32'h4411caf4, 32'h405e16cc, 32'hc0e22d7a},
  {32'hc34d0850, 32'h433ba083, 32'h4371ef94},
  {32'h4458af36, 32'h426bef9f, 32'h432f684d},
  {32'hc35e0ee0, 32'hc159f516, 32'hc329c7b6},
  {32'h4311e990, 32'hc26e3720, 32'h427fe21a},
  {32'hc3578690, 32'h41cf0c3a, 32'hc31de6b0},
  {32'h44925fac, 32'hc3dc315b, 32'h43924cff},
  {32'hc3c01caa, 32'h43d12d04, 32'h437ac8e2},
  {32'h449a1d16, 32'h4240c95c, 32'h434c810b},
  {32'hc4d78db8, 32'h430ccce5, 32'h432ffb91},
  {32'h4468ca67, 32'hc040dabb, 32'hc40bfc76},
  {32'hc3836965, 32'h4338feca, 32'h431951d4},
  {32'h44e0091f, 32'hc31d2bc1, 32'h43c10f40},
  {32'hc42f8848, 32'hc3916af5, 32'h4216ee3f},
  {32'h44994016, 32'h420a21a5, 32'h42e4785a},
  {32'hc4c9096c, 32'h42fbefc0, 32'hc29ca0ac},
  {32'h4515142a, 32'hc07bcb62, 32'h43e333ab},
  {32'hc4ce9896, 32'h4329ff7b, 32'hc2fcd0d4},
  {32'h43342660, 32'h4247d7b2, 32'h42b05459},
  {32'h42b93d5d, 32'hc2b46f84, 32'h4154e426},
  {32'h4427cc40, 32'h43184152, 32'h429bac95},
  {32'hc4f4c916, 32'hc2eae4a0, 32'hc3178136},
  {32'h4482ec25, 32'hc38bf030, 32'h42a08000},
  {32'hc4a33604, 32'h42f045ea, 32'h4269b94b},
  {32'h448b1a50, 32'h438de451, 32'h41ed85ea},
  {32'hc49133a4, 32'h42cd9513, 32'hc3d2dead},
  {32'h449e60cb, 32'hc29acdf2, 32'hc3afc8ee},
  {32'h428c6620, 32'hc413888a, 32'hc3b6687e},
  {32'h435a097c, 32'h434eed34, 32'hc3ba9de6},
  {32'hc484f0b6, 32'h438a45f0, 32'h433463ab},
  {32'h451ffc32, 32'hc3835252, 32'h43d4137d},
  {32'hc4d11d33, 32'hc1c63b4a, 32'hc187faa7},
  {32'h43aaceba, 32'hc1eeecbc, 32'h438f4cf5},
  {32'hc4176dc7, 32'hc2d02fdb, 32'h43c8ec40},
  {32'h45150ae3, 32'h43f04369, 32'h43d5abbc},
  {32'hc45bef6e, 32'hc372019c, 32'h4316b216},
  {32'h43a61613, 32'h43b49175, 32'h4359bae3},
  {32'hc30ead18, 32'h44034ec2, 32'h420fd638},
  {32'h445947c9, 32'hc37f7c85, 32'h41e4d043},
  {32'hc496bccf, 32'hc21f15f4, 32'h4308c72c},
  {32'h437252b0, 32'h431aca94, 32'h4378cb79},
  {32'hc4b14d3c, 32'hc29f0d0a, 32'hc2c4908c},
  {32'h44b33b65, 32'h43120cd7, 32'hc2e63971},
  {32'hc50734fc, 32'hc260c169, 32'hc3692622},
  {32'hc0867900, 32'h42a508d4, 32'h40a78655},
  {32'hc467fe76, 32'hc2a6162e, 32'h4396e649},
  {32'h446f9eac, 32'hc31aaaad, 32'hc41fa858},
  {32'hc4cbcebd, 32'h3f967ba0, 32'hc3005bd7},
  {32'h449f4bec, 32'h431bd262, 32'h43194c05},
  {32'hc36bdce0, 32'hc3e4f19a, 32'hbfaff3ac},
  {32'h43a0d8a8, 32'h416b8190, 32'hc2f075f2},
  {32'hc1fd3642, 32'hc2b3b9f3, 32'hc392eb77},
  {32'hc38e6b59, 32'hc1da227b, 32'hc335a6e4},
  {32'hc4c09531, 32'hc213cbac, 32'h4264395a},
  {32'h448dee6c, 32'h43854920, 32'h43911d5f},
  {32'h432735c0, 32'hc1f57ac8, 32'hc15ec5c2},
  {32'h44ed68c5, 32'h4307e179, 32'hc2315bd1},
  {32'hc50e1888, 32'hc3584b3b, 32'hc40ecdb8},
  {32'h44c4f4f2, 32'h424e6300, 32'h42b50cba},
  {32'hc4bf784f, 32'h41e9fdd6, 32'h4396743b},
  {32'h449a60af, 32'h430c4d24, 32'hc2cbaf3c},
  {32'hc4836117, 32'h4417621c, 32'hc35605c3},
  {32'h44bd5296, 32'h434b28e0, 32'h43bc644c},
  {32'hc4bf9327, 32'hbf1d6d6c, 32'h437cd088},
  {32'h43aedf56, 32'hc3c7fc86, 32'h4310292b},
  {32'hc4d33297, 32'h4362ff76, 32'h421cc2b8},
  {32'h44057cc6, 32'h4317fb9a, 32'hc2c5bdc4},
  {32'hc4acb8ce, 32'hc3e1d3ba, 32'h44011a7a},
  {32'h44aa3a50, 32'h438a7ded, 32'h414ad6c9},
  {32'hc4a2bcac, 32'h42aa8791, 32'h42b4b484},
  {32'h431a0df0, 32'h42a8bb9c, 32'h41d0fdbd},
  {32'hc4966bc1, 32'h43a0e1ec, 32'h41a6fc84},
  {32'h448b47d8, 32'h42895fef, 32'hc365b056},
  {32'h420e0d4e, 32'h4168831f, 32'h41cfcda8},
  {32'h43c58cee, 32'hc3a04a7a, 32'hc391fbbb},
  {32'hc4e10589, 32'hc34961fa, 32'h433ff791},
  {32'h45119680, 32'hc37384db, 32'hc31d327c},
  {32'hc39b4704, 32'hc35cb96c, 32'h419f28d8},
  {32'h44a6f970, 32'h42068710, 32'h4329ea16},
  {32'hc4d94180, 32'hc294ef36, 32'hc1a42106},
  {32'hc2639ba0, 32'hc1e0595e, 32'hc273bae8},
  {32'hc40c9b37, 32'h436a7e6b, 32'hc3da4dba},
  {32'h44989495, 32'hc2b320ca, 32'hc20b036c},
  {32'hc3d08fe0, 32'hc306329a, 32'h43852790},
  {32'h43bf5bcf, 32'hc2d03e0e, 32'hc3036bb8},
  {32'hc478a2de, 32'hc2f12f73, 32'hc3c09302},
  {32'h44adb102, 32'h3f1edcc0, 32'hc32c1997},
  {32'hc2abe088, 32'hc230c358, 32'h4166bdec},
  {32'h43ea9ea0, 32'hc243ea3e, 32'h436c5454},
  {32'hc5007eaf, 32'h42d26470, 32'hc327c524},
  {32'h4480a156, 32'h422ff128, 32'hc2999398},
  {32'hc504c7ef, 32'hc38650c7, 32'h42f835cb},
  {32'h44ce5a02, 32'hc348f7ea, 32'hc32c2fc6},
  {32'hc4136ba8, 32'h42b84984, 32'hc22bf869},
  {32'hc2fc5bf0, 32'h43f79dc3, 32'h42dcec3b},
  {32'hc4d7cf62, 32'hc32eb31a, 32'h43707f69},
  {32'h4313def8, 32'h43169349, 32'h43b9fba6},
  {32'hc490f320, 32'hc388d749, 32'hc3159d94},
  {32'h43dad2ba, 32'hc27e75b3, 32'hc1f99f84},
  {32'hc4682246, 32'h420f2dcf, 32'hc299a7bf},
  {32'h4400430e, 32'h42231ee4, 32'hc29089a6},
  {32'hc481dbc2, 32'hc25e8a8a, 32'h42bc2525},
  {32'h44aebf32, 32'hc36b757b, 32'h432aa821},
  {32'hc503b690, 32'h430544d9, 32'hc2d3c173},
  {32'h44f8e29d, 32'hc2c0033e, 32'hc39390bf},
  {32'hc3b4f2f4, 32'h42a5d20b, 32'hc2221f1f},
  {32'h447ca0d0, 32'h43c984a0, 32'h432faa5f},
  {32'hc4b233b7, 32'h43180ad6, 32'hc1ad235d},
  {32'h4418227e, 32'hc3257b37, 32'hc363f372},
  {32'hc3d1f596, 32'h43a3c222, 32'h432706f5},
  {32'h44f40c30, 32'hc37c2133, 32'hc27691ad},
  {32'hc4babce7, 32'h42555990, 32'hc3ae7cbc},
  {32'h4495412e, 32'hc2130670, 32'hc0d8abb5},
  {32'h43064235, 32'h43fd6db3, 32'hc31f4fba},
  {32'hc29f9780, 32'hc30fe855, 32'hc309fb82},
  {32'hc4cdb838, 32'h4397731e, 32'h43000c19},
  {32'h444113be, 32'h430f6e10, 32'hc3f8ef05},
  {32'hc50146d1, 32'hc3803952, 32'h433eb613},
  {32'h43e08850, 32'h43b49d97, 32'hc37c63cd},
  {32'hc50a9b5a, 32'hc2fb0148, 32'h43fc0224},
  {32'h451ad556, 32'h43871994, 32'h41b4d374},
  {32'hc1cb8080, 32'hc385c22d, 32'hc3a3b223},
  {32'h44e26075, 32'hc3bdf469, 32'h433b9ab9},
  {32'hc4d085a4, 32'h43d34b30, 32'h438a602d},
  {32'h44339f81, 32'hc312ae43, 32'h42f82bb6},
  {32'hc50dbc6b, 32'h421bbf76, 32'hc31e48ba},
  {32'h449e0336, 32'hc2fa75f9, 32'hc30c87bf},
  {32'hc3fe90eb, 32'h423e9e00, 32'h4248a9c2},
  {32'h44f9726f, 32'h424b9880, 32'h42c499e6},
  {32'hc506baa7, 32'hc39c9489, 32'hc2834571},
  {32'h4406a21e, 32'hc3691c9a, 32'hc336cb1a},
  {32'hc23049d2, 32'hc333a7f1, 32'h431fe823},
  {32'h44fed2dc, 32'hc2ebd193, 32'h42d9b0f2},
  {32'hc4feb9a0, 32'h4332c40e, 32'h43464b6d},
  {32'h440dd8d1, 32'hc303f1f3, 32'h41eee056},
  {32'hc3e2bc74, 32'h42ed273b, 32'h4408e581},
  {32'h447cf338, 32'hc30cab53, 32'hc30682ba},
  {32'hc3f154f0, 32'hc3b23f51, 32'hc348fc57},
  {32'h449235a4, 32'hc3f4d29e, 32'hc23370d2},
  {32'hc4fdda14, 32'h42f03ee5, 32'hc3aa0e87},
  {32'h44964a4e, 32'h439a5f93, 32'h437c5a67},
  {32'hc5043561, 32'h43593f0a, 32'hc3315f69},
  {32'h4437390c, 32'h42b66f93, 32'h421414cf},
  {32'hc48edbda, 32'hc2f704fc, 32'h43037e11},
  {32'h444b50a2, 32'hc33d7240, 32'hc2e0cd01},
  {32'hc35a6390, 32'h4283238f, 32'h42898270},
  {32'h442be43e, 32'hc291d369, 32'hc310db85},
  {32'hc4e48e88, 32'h42b9227b, 32'hc33bb7b1},
  {32'h44c3c709, 32'hc2cc1669, 32'hc3a57f74},
  {32'hc27a9c20, 32'h4376fd46, 32'hc39406bd},
  {32'h4518caed, 32'h43c99ce3, 32'hc3c537a6},
  {32'hc2c8f6a7, 32'hc3a4d479, 32'h4349bcc8},
  {32'h44cd8a6b, 32'hc38b40e3, 32'hc23cacda},
  {32'hc504f1f2, 32'h42938a1c, 32'h43a24ba0},
  {32'h44bcb9ca, 32'hc2dde174, 32'hc373e0c4},
  {32'hc50bdcf9, 32'hc3379600, 32'hc3bec770},
  {32'h44254832, 32'h43383b47, 32'hc39149cc},
  {32'hc49b0cf7, 32'hc3a048aa, 32'h4369d2f6},
  {32'h41850540, 32'h42b5931a, 32'h40454450},
  {32'hc455bd58, 32'h430194c5, 32'hc38f2252},
  {32'h44d01087, 32'h425d77f8, 32'hc362885c},
  {32'hc3cc9850, 32'hc11af286, 32'hc3961dda},
  {32'h44899252, 32'h4319b11b, 32'hc1bb9752},
  {32'hc45e7135, 32'hc3ad71e6, 32'h427f0d41},
  {32'h414f4fb0, 32'hc3a6e728, 32'hc2ec675e},
  {32'hc4e9a85c, 32'h430f334c, 32'h436af6c6},
  {32'h44cb322a, 32'h430c7a77, 32'hc2f054c7},
  {32'hc4d27e99, 32'hc3a62b7b, 32'hc3972821},
  {32'h43d0fd45, 32'hc3c78bb0, 32'h43074662},
  {32'hc4ea12d9, 32'hc34da5d8, 32'h4206883e},
  {32'h45095033, 32'hc34fa6f6, 32'hc30325b5},
  {32'hc3a21360, 32'h429e9122, 32'hc3d3d1a9},
  {32'h44c606a2, 32'h43643d4f, 32'hc2159993},
  {32'h4311bef0, 32'h436b46c8, 32'hc356f5f9},
  {32'h44604cbd, 32'h420ca876, 32'hc303784b},
  {32'hc5055284, 32'hc3e9a276, 32'h42eabfd7},
  {32'h450c5b66, 32'hc2b1a57a, 32'h4387b847},
  {32'hc50a1770, 32'hc397066e, 32'h4240996a},
  {32'h44c2bc38, 32'hc2021d39, 32'hc30f35e9},
  {32'hc4e8310f, 32'hc3c86b95, 32'h4206d4dd},
  {32'h44e724ce, 32'hc319672e, 32'hc4340014},
  {32'hc4c561e3, 32'h42d9114f, 32'h432e9113},
  {32'h449eb5b7, 32'hc0a25bd0, 32'h43f1fef1},
  {32'hc482cec6, 32'h432d4ab1, 32'h43de39c5},
  {32'h43d48526, 32'hc2a3cc19, 32'h43b936ef},
  {32'hc4d7fcac, 32'h42af2738, 32'h42a09451},
  {32'h4484718b, 32'h430a95bc, 32'h4405adfc},
  {32'hc4e0e445, 32'h41045a90, 32'h43734d9d},
  {32'h4476af35, 32'h434c64e3, 32'hc3f1768e},
  {32'hc299b5e0, 32'h4280014c, 32'h439ab896},
  {32'h4505ecd5, 32'hc3aec4df, 32'h433a43a3},
  {32'hc426d880, 32'hc14e8cd8, 32'h439dca57},
  {32'h44830454, 32'hc3ab52cf, 32'hc30d5ef1},
  {32'hc40806e1, 32'h42d7f6fb, 32'h429046c7},
  {32'h441c14cc, 32'h4210ea11, 32'h41986482},
  {32'hc4a3ff41, 32'hc224edc0, 32'hc3884448},
  {32'h44b608ef, 32'hc18454c5, 32'h42f1ac1d},
  {32'hc4957d51, 32'hc324f154, 32'h431532b4},
  {32'h4457f552, 32'h43b938bc, 32'h4198785b},
  {32'hc432ec22, 32'h4272a098, 32'h42eb8d56},
  {32'h44f026f0, 32'h4283265a, 32'h430dd931},
  {32'hc3ab56f2, 32'hc1999094, 32'hc3c3eeff},
  {32'h44c2065a, 32'hc453e7d5, 32'h42e11248},
  {32'h4298759e, 32'hc2cfed8f, 32'hc36c9101},
  {32'h43d9ede7, 32'hc32cfe8b, 32'hc260509d},
  {32'hc48c2e4a, 32'h42103c9b, 32'h41af9028},
  {32'h4433286e, 32'h422718bc, 32'hc243fbc5},
  {32'hc4c148c9, 32'hc24f5396, 32'hc2f7d0a3},
  {32'h43d1ee1c, 32'hc30e661b, 32'h43ddadc3},
  {32'hc3d8d6ec, 32'hc3a21c82, 32'h41f5dc68},
  {32'h4428ca0c, 32'hc31e6817, 32'hc12e3ef9},
  {32'hc44b5a6c, 32'hc2b23ba4, 32'h43cd26c4},
  {32'h44bdb0b6, 32'hc23378b5, 32'hc3c6fe6b},
  {32'hc28b039c, 32'h4301a62c, 32'h404e882e},
  {32'h448ef47a, 32'hc3505195, 32'h42f2c56d},
  {32'hc3e240e9, 32'h43bd16ae, 32'hc339c86b},
  {32'h4486363c, 32'h435dbac4, 32'h40c403da},
  {32'h42d36840, 32'h43c7e8e2, 32'h430d950f},
  {32'h44eebe19, 32'h42da039f, 32'hc2af2149},
  {32'hc4ee1f5c, 32'h4352071b, 32'hc35fa006},
  {32'h446cc41a, 32'hc3accb62, 32'h424714df},
  {32'hc50e1b77, 32'hc014b070, 32'h438c98be},
  {32'h44a547ce, 32'hc2787ed3, 32'hc2a52359},
  {32'hc357b238, 32'hc3099f57, 32'hc3cfb439},
  {32'h43ae6b3b, 32'hc3538362, 32'h429f99ae},
  {32'hc321fdc0, 32'h43b757ec, 32'h421e485e},
  {32'h44d51d3a, 32'hc3137b8c, 32'h413aa3cc},
  {32'hc418b2b2, 32'hc20bd88d, 32'h43c364d4},
  {32'h43c5e9dc, 32'hc1d110bc, 32'h43d6235d},
  {32'hc502e6bb, 32'h44010f54, 32'hc2987808},
  {32'h44b48b26, 32'hc314b905, 32'h430aea36},
  {32'hc3b84ab0, 32'h4345447d, 32'h43b3d5b2},
  {32'h450e8533, 32'h43b95abe, 32'hc369f928},
  {32'hc4e9b622, 32'hc2f0f1f6, 32'h4214c2c5},
  {32'h44c0a4fb, 32'h43098a88, 32'h41b13277},
  {32'hc493deb2, 32'hc4015eba, 32'h42ec976c},
  {32'h43a764d0, 32'hc34f91ed, 32'hc38a69dc},
  {32'hc3aeafec, 32'h42d6358b, 32'hc3d946a1},
  {32'h441073ed, 32'h437f94fc, 32'hc2c5cce7},
  {32'hc42816a4, 32'hc3993800, 32'hc1bdada7},
  {32'h44c4cf0f, 32'hc403d5d0, 32'hc3dcbe86},
  {32'hc50f5cb0, 32'hc3905923, 32'hc281b8ed},
  {32'hc3a62e50, 32'hc2ca5739, 32'hc15d7789},
  {32'hc44d71cc, 32'hc399301b, 32'hc2d03cf9},
  {32'h428f2016, 32'hc3976535, 32'h43a72dc5},
  {32'hc436a7d2, 32'hc302e3cd, 32'hc2ebabf0},
  {32'h42ff3977, 32'h434d0482, 32'h42eabfe1},
  {32'hc4fed314, 32'h436ede0f, 32'h438ffbb5},
  {32'h449d677b, 32'hc420b3bb, 32'hc2a7cdfa},
  {32'hc48dedc9, 32'hc2622a07, 32'h43e07692},
  {32'h4486ad8f, 32'h434a6e91, 32'hc3544683},
  {32'hc492c576, 32'h439e49d9, 32'h4209b2d8},
  {32'h4415da84, 32'h42292d2a, 32'hc2c78d40},
  {32'hc4ecfff9, 32'h43404de9, 32'h433f0c3b},
  {32'h4408f795, 32'hc31dde37, 32'h43ee93db},
  {32'hc3eb36d6, 32'h436eb686, 32'h42b9c985},
  {32'h447aa418, 32'hc07a8728, 32'hc2ac8570},
  {32'hc4918d5d, 32'hc3cb4772, 32'h435aa1b9},
  {32'h441406cc, 32'h439797bc, 32'h428fa34e},
  {32'hc4eecc8a, 32'hc33a046b, 32'h4240770c},
  {32'h44033178, 32'hc3e98bb1, 32'h43d9fe1b},
  {32'hc3c4d786, 32'h4327a2b1, 32'h4277f5ad},
  {32'h448f6214, 32'hc274f0d8, 32'hc2bcc0de},
  {32'hc4bd0b22, 32'hc1ccb779, 32'hc33bc677},
  {32'h44f7a472, 32'hc3c64b41, 32'h43f1eae9},
  {32'hc46bc0b4, 32'hc1db33d4, 32'hc24e40c5},
  {32'h45130d92, 32'hc24b7230, 32'h43d97f06},
  {32'hc21ea900, 32'h4421f92a, 32'h412d07f0},
  {32'h437fc474, 32'hc2ff7d4c, 32'hc13d37c6},
  {32'hc502e67f, 32'h4262f9d7, 32'h40d11a60},
  {32'h44601a4f, 32'hc344443c, 32'h431e464f},
  {32'hc40117a8, 32'h44188ea4, 32'hc36624d3},
  {32'h44ddbc6c, 32'h434a2d0b, 32'hc32e67f9},
  {32'hc51d5d06, 32'hc3488115, 32'h43e5309c},
  {32'h41a5a400, 32'hc33a77ef, 32'hc313a109},
  {32'hc526c916, 32'h42bd6301, 32'hc3b6276a},
  {32'h44e05dde, 32'hc2de54aa, 32'h430cf0e0},
  {32'h4318a548, 32'hc246ee81, 32'h43bb6de7},
  {32'h444d9c7c, 32'h42ccb07e, 32'h4216a6d6},
  {32'hc4eb143e, 32'hc3129ee8, 32'h435588f7},
  {32'h44de086d, 32'h43ad502a, 32'hc0d3e501},
  {32'hc5006566, 32'h43abd280, 32'h430b32ef},
  {32'h43ae0733, 32'h433b898e, 32'hc3a30d23},
  {32'hc45f606d, 32'h43766b51, 32'hc3d8f973},
  {32'h44d71c38, 32'h4127435c, 32'hc344f851},
  {32'hc421fb73, 32'h43082669, 32'hc3e9d798},
  {32'h44d4e256, 32'hc2a0bd7a, 32'h42b45047},
  {32'hc4dbeaf8, 32'hc24c9ef1, 32'hc3007e2e},
  {32'h442b5c30, 32'hc3913d25, 32'hc38e8332},
  {32'hc4af00c1, 32'hc312fc22, 32'hc3464203},
  {32'h4501ec80, 32'h4348f008, 32'hc34b7da1},
  {32'hc51458ed, 32'h42c78a8f, 32'hc3cfb34c},
  {32'h43ca83b8, 32'hc417221d, 32'hc3061982},
  {32'hc47b8d2c, 32'hc1719341, 32'h42ad5930},
  {32'h44f0bb32, 32'hc318b30a, 32'h43c652f1},
  {32'hc3f9a0e8, 32'h43a0cc69, 32'h42e3c358},
  {32'h45149e54, 32'h41c35ba1, 32'h426c0d1c},
  {32'hc4a5a4c9, 32'hc32be6ef, 32'hc3342e15},
  {32'h44034060, 32'h43a6ae67, 32'hc3499052},
  {32'hc49a8e46, 32'hc40b662e, 32'hc1ce8066},
  {32'h447f7c4a, 32'hc2fd1a53, 32'hc291091e},
  {32'hc50101aa, 32'hc24d9152, 32'h428880e6},
  {32'h44d26ad2, 32'hc2db2682, 32'hc3db983f},
  {32'hc487ed70, 32'hc36dd7e1, 32'hc2d175b7},
  {32'h447ea1d0, 32'h4215e582, 32'hc3b28705},
  {32'hc49c2e98, 32'h439ff9f9, 32'h43f48211},
  {32'h44deaee0, 32'h435cde9a, 32'h4406652d},
  {32'hc36e2d10, 32'hc2e6cd84, 32'h42a2bca2},
  {32'h43abeb44, 32'h41ce9e1e, 32'hc23f9913},
  {32'hc2bece54, 32'hc3ceaa13, 32'hc32ae3d5},
  {32'h44ae0340, 32'hc205de80, 32'hc1f3d625},
  {32'hc52f23d0, 32'h4336bbd1, 32'h405561af},
  {32'h42502be0, 32'h414a87d3, 32'hc25919ac},
  {32'hc4566294, 32'hc3b2c3d6, 32'h40da6fcc},
  {32'h44e6f61d, 32'h42952d58, 32'hc1bf5829},
  {32'hc3d5b6b8, 32'h427e29ca, 32'h4348dd54},
  {32'h44f6ba5e, 32'hc38a4029, 32'hc30ae0aa},
  {32'hc4c57e5c, 32'h42d546d9, 32'hc3b1b00c},
  {32'h438be3f3, 32'hc3a5c766, 32'h425f0efc},
  {32'hc50f54dc, 32'hc2b8f013, 32'hc0911f0f},
  {32'h45142f8b, 32'hc35835d7, 32'hc38cde77},
  {32'hc41d43da, 32'h43046413, 32'h42c93700},
  {32'h43f728a2, 32'hc16c0510, 32'hc30e7b10},
  {32'hc4437836, 32'h43730e6b, 32'h43cb8a9a},
  {32'h443700fb, 32'h423f7cac, 32'h42b11f8f},
  {32'hc2c34160, 32'hc408f52f, 32'hc10b58e2},
  {32'h44d13ef6, 32'hc20cea93, 32'hc30b68e8},
  {32'hc4fa3701, 32'h40af363f, 32'hc34d0f36},
  {32'h4484c23c, 32'hc3ab8389, 32'h430889d2},
  {32'hc3953746, 32'hc34c39b7, 32'hc3a06586},
  {32'h445351e6, 32'h43416d97, 32'hc3987bbd},
  {32'hc4b1450d, 32'hc09ca223, 32'hc3443143},
  {32'h44c790e0, 32'hc23a1bc2, 32'h431debb7},
  {32'hc3ff3f4c, 32'hc342d03b, 32'h42e736fd},
  {32'h441762d0, 32'h43784572, 32'hc04fa990},
  {32'hc4836c6a, 32'h4301bd70, 32'hc2a4d787},
  {32'h44ab37bb, 32'hc265678e, 32'hc33523c2},
  {32'hc49eeb65, 32'h42cca79f, 32'hc117201f},
  {32'h44c047a2, 32'h41a064aa, 32'h43db3d75},
  {32'hc49d679c, 32'h4235fb4c, 32'hc1a92a12},
  {32'h448cb6b8, 32'hc20c14f0, 32'hc35ba3b6},
  {32'hc4ea40fc, 32'h415c7244, 32'h423ae564},
  {32'h44db3b24, 32'hc1a3e383, 32'hc32dff7d},
  {32'hc402ca9c, 32'h42738ca4, 32'hc40ffe24},
  {32'h450da5e5, 32'hc3ae25fa, 32'h428bcb11},
  {32'hc46a7d3a, 32'hc2ae9933, 32'h43a33747},
  {32'h44f69893, 32'hc2bf7f02, 32'h4385e7eb},
  {32'hc50184b9, 32'hc0ea4040, 32'hc376972c},
  {32'h44c6d900, 32'hc3321fcf, 32'h43221e68},
  {32'hc38c1508, 32'h4305ca87, 32'hc22c9b16},
  {32'h4408a70c, 32'h4348072c, 32'h3fd19f64},
  {32'hc4d14fb5, 32'h4312b70b, 32'hc236d6c7},
  {32'h449faa71, 32'hc2dc50b9, 32'hc25f6f6d},
  {32'hc4982412, 32'h436d14d9, 32'h435271c9},
  {32'h44929bd6, 32'hc4178596, 32'h4342d3d4},
  {32'hc4f9e926, 32'h4320c141, 32'h43aed8c9},
  {32'h44d6a068, 32'hc35786ee, 32'hc3430347},
  {32'hc50a3279, 32'h43af54ec, 32'h43b16b8c},
  {32'h43e1d3b8, 32'h426d3683, 32'hc35b5ada},
  {32'hc46b203a, 32'h433887a7, 32'h429a7f27},
  {32'h45103d12, 32'hc32965ce, 32'hc38a77af},
  {32'hc4271ef0, 32'h4359d0ed, 32'h42e2ee78},
  {32'h45089c9f, 32'h438e7f16, 32'h4334c7af},
  {32'hc483073c, 32'hc2832c99, 32'hc1df852c},
  {32'h43e2ed7e, 32'hc382af77, 32'hc27d9f7a},
  {32'hc436cdd8, 32'hc2612f14, 32'h41d4c9f5},
  {32'h450bc6bf, 32'h42338e1b, 32'hc3004764},
  {32'hc4216e85, 32'h42920b8a, 32'h4314492a},
  {32'h44b9dfe1, 32'h43b7339d, 32'hc354f236},
  {32'hc3d714a1, 32'hc1542e1f, 32'h42caf187},
  {32'h44b81d27, 32'hc2cd73de, 32'hc3862520},
  {32'hc4e90555, 32'h42290943, 32'h43548aba},
  {32'h44b410cd, 32'h428781c1, 32'hc37fea89},
  {32'hc4dec086, 32'hc2fb2f0e, 32'h430ddc18},
  {32'h44d08d02, 32'hc1541ac8, 32'h432b9e37},
  {32'hc489f374, 32'h4308b998, 32'hc30e1cce},
  {32'h44c84b03, 32'hc1a2f3ad, 32'hc386ac04},
  {32'hc4a13005, 32'h43843f0f, 32'h437c7b0e},
  {32'h447e2e35, 32'h426703d3, 32'h4357ad16},
  {32'hc4cd4999, 32'hc2836604, 32'h437c091f},
  {32'h44da7b0c, 32'hc2c21c06, 32'hc22aced1},
  {32'hc50af19f, 32'hc307c8a1, 32'h4286751b},
  {32'h45116538, 32'hc30f480e, 32'h4382932c},
  {32'hc49ec7b7, 32'hc36ed7e7, 32'h43a06630},
  {32'h44b5f4f8, 32'hc38fbc68, 32'hc2a85633},
  {32'hc4f3ee55, 32'h4362281f, 32'hc1a0d0d9},
  {32'h44c2c7fe, 32'hc212d40f, 32'hc3c914b8},
  {32'hc512738e, 32'h432c2143, 32'h43bf357f},
  {32'h44dc09d6, 32'h41a0306e, 32'h43a4a516},
  {32'hc02b5c00, 32'h4386f53d, 32'hc2e70ef3},
  {32'h44b61476, 32'h4300129a, 32'hc1f883f2},
  {32'hc413e55c, 32'hc3af69b4, 32'h4330b4ab},
  {32'h44a91c60, 32'h4325d036, 32'h4293eb3a},
  {32'hc4df408d, 32'hc2ea9a12, 32'h42be4e9c},
  {32'h44f355c2, 32'h41e1b2de, 32'hc117c8ed},
  {32'hc4fdeae1, 32'h430543d3, 32'h42450c7e},
  {32'h43cd2978, 32'hc23c7d12, 32'hc30f59cb},
  {32'hc4d79746, 32'hc31c1be9, 32'h42a2f82e},
  {32'h44cfcdc2, 32'h4358d0dd, 32'h423ea31e},
  {32'h4396b45f, 32'h42bf61bb, 32'hc2cbdbfe},
  {32'h43ad77da, 32'hc2779a3f, 32'h42ae47de},
  {32'h444e106e, 32'hc3433d3b, 32'h422aada4},
  {32'hc44a5291, 32'hc2bc11f5, 32'h412e4809},
  {32'h449efc1b, 32'h438cd528, 32'hc14dd06b},
  {32'hc4964bf7, 32'h4381268f, 32'h434f1ff8},
  {32'h44e3571c, 32'hc34f6943, 32'h43102e6c},
  {32'hc4bda9fc, 32'hc1ec7c06, 32'h40f5e5a6},
  {32'hc2dc7a60, 32'h430970ad, 32'hc2dcea4c},
  {32'hc410b72a, 32'h436dd1dc, 32'hc2e3422d},
  {32'h44ec1dd4, 32'hc0ea1330, 32'hc358a83b},
  {32'hc43d7988, 32'h4280913c, 32'h425740d2},
  {32'h45209269, 32'hc2ed211a, 32'hc334387e},
  {32'hc41e6b1a, 32'h42e89ba8, 32'h4398f6bf},
  {32'h44edc1a0, 32'h42aef138, 32'h433059c3},
  {32'hc420430b, 32'hc3050d36, 32'hc39ce759},
  {32'h450f123c, 32'hc399f8c0, 32'h42dc7199},
  {32'hc511aa3e, 32'h4230fd3f, 32'hc2673cd7},
  {32'h44828236, 32'h438d319a, 32'hc391e53a},
  {32'hc4f78c77, 32'hc2c40640, 32'h43bbc0cb},
  {32'h44a02f0d, 32'hc0201528, 32'h4345f075},
  {32'hc337b688, 32'h4233587e, 32'hc34b9fa6},
  {32'h44cb4a23, 32'h40199d2e, 32'h42a338b6},
  {32'hc3175b00, 32'h4369d6f4, 32'hc3b5167d},
  {32'h4493c544, 32'h43268b03, 32'hc3878ff5},
  {32'hc4d6d93e, 32'h429d1217, 32'h432de5ce},
  {32'h45164c7b, 32'hc116dc64, 32'hc334d2af},
  {32'hc4ff2f74, 32'hc380d06a, 32'hc38af628},
  {32'h442bd887, 32'h423782a3, 32'h4280db6c},
  {32'hc4822c0b, 32'h429085ad, 32'hc32e6701},
  {32'h44a3c8c1, 32'h431f87ed, 32'hc3641687},
  {32'hc4dbe417, 32'h43362e8e, 32'hc308764d},
  {32'h43ef7450, 32'hc09a4a1e, 32'hc392745d},
  {32'hc4aec85e, 32'h431ad500, 32'hc32a1957},
  {32'h44f086e4, 32'hc2bb3469, 32'h40862365},
  {32'hc5023544, 32'h433153a9, 32'hc2d5b116},
  {32'h44e7c8be, 32'h437adb9e, 32'hc2de2003},
  {32'hc4ad50a5, 32'hc2633171, 32'h4385c417},
  {32'h4503f282, 32'h41ca2697, 32'hc381870f},
  {32'hc4e145a2, 32'hc3a9ab60, 32'h43b7f654},
  {32'h4512dd7e, 32'hc42a257d, 32'h428e9aea},
  {32'hc27f61a8, 32'hc3a10d8f, 32'h4383c833},
  {32'hc2877cb0, 32'h43548d1a, 32'h4315a55a},
  {32'hc4ba457a, 32'hc352373c, 32'hc2d76f38},
  {32'h43be68d0, 32'h43c38f3b, 32'hc1ae4ffa},
  {32'hc5132d30, 32'h438757ef, 32'h428e9e91},
  {32'h45184651, 32'hc20c08d8, 32'h43a09387},
  {32'hc4fd1b61, 32'h4317f27c, 32'h42d7c5e6},
  {32'h450d0c00, 32'h4208b41b, 32'hc1eba905},
  {32'hc5166005, 32'h437f36cd, 32'hbfcda0e4},
  {32'h448e5013, 32'hc2d1f71b, 32'h439f8f97},
  {32'hc4a42f67, 32'hc258367e, 32'hc2299f9e},
  {32'h453125ed, 32'h41a3a414, 32'h42cce7eb},
  {32'hc5026df0, 32'h42fee6e1, 32'h423b1d12},
  {32'hc1040000, 32'h432723cd, 32'hc37a7191},
  {32'h42572a00, 32'hc221caa7, 32'h4336b95b},
  {32'h44e91820, 32'h4383cb53, 32'hc2a7bbc9},
  {32'hc4f6477a, 32'h431407d0, 32'hc2f60607},
  {32'h44061176, 32'h42b9d46f, 32'h42f85d2d},
  {32'hc3864c08, 32'hc31120e0, 32'hc3d5fc9f},
  {32'h43ec609c, 32'hc3fcff71, 32'hc398724c},
  {32'h4097c700, 32'h4194613d, 32'hc3ac7f74},
  {32'h4508c8dc, 32'hc20bb5b1, 32'h42ab59ed},
  {32'hc5058bfe, 32'hc4016e27, 32'hc34e8c2b},
  {32'h44e7f60e, 32'h43870b66, 32'hc179d958},
  {32'hc4327964, 32'hc2308a75, 32'h43562832},
  {32'h44f5238a, 32'h43c746df, 32'h43a177c5},
  {32'hc453352c, 32'h43a5d4ce, 32'h43b44083},
  {32'h44ed9ce9, 32'h43210a5c, 32'hc3e76816},
  {32'hc4ffbb79, 32'h4356cf89, 32'hc0fbf569},
  {32'h449c7f82, 32'h4280b767, 32'h431aa53c},
  {32'hc3c2e504, 32'hc32cd037, 32'hc39cbcce},
  {32'h44a36de1, 32'h41fe5439, 32'h4376c4a6},
  {32'hc5015166, 32'h42d0c0e7, 32'h42f843cf},
  {32'h4509b9c2, 32'hc36aad2f, 32'h43bca5e2},
  {32'hc4c03e8d, 32'h419681af, 32'hc1b8d04f},
  {32'h446f1301, 32'h4332c86e, 32'h43936d45},
  {32'hc4520fa2, 32'h43d7b036, 32'hc393ea0c},
  {32'h450ca75b, 32'h43596454, 32'hc29be0c3},
  {32'hc4c9982f, 32'h43f04934, 32'h42cd1358},
  {32'h45094d16, 32'hc19d053a, 32'h43211c9a},
  {32'hc4ee10ea, 32'hc3ae5a43, 32'hc3d77e55},
  {32'h4460e48a, 32'h438d4454, 32'h422991dd},
  {32'hc4bd3539, 32'h42caf390, 32'h420b0cee},
  {32'h44ba5322, 32'h430b0399, 32'h42f61fe1},
  {32'hc486bcdd, 32'h426cd4ce, 32'hc31827b1},
  {32'h44a6ebfa, 32'hc368973b, 32'h429b9c62},
  {32'hc282df90, 32'hc225ea1c, 32'h4233b6dd},
  {32'h4375bcd0, 32'h429128b1, 32'hc33f76b2},
  {32'hc4d10166, 32'h43128f07, 32'h4233ea0a},
  {32'h450e72ba, 32'hc3c3c66d, 32'h41bf50d4},
  {32'hc50061ff, 32'h40bf5229, 32'hc350a095},
  {32'h45116cd3, 32'hc186bb17, 32'hc331fa26},
  {32'hc511b698, 32'hc2ef214b, 32'hc0803906},
  {32'h44ae0e71, 32'h4351fc7d, 32'h4292a6c3},
  {32'hc22aaac0, 32'hc195ff57, 32'hc2c77d5a},
  {32'h449cae68, 32'h42ba26e4, 32'hc2066cba},
  {32'hc419ef5c, 32'h429f22e7, 32'h426ee02d},
  {32'h452ac7d7, 32'hc294ed3f, 32'h4296b582},
  {32'hc503db08, 32'hc37f8793, 32'h432f25e0},
  {32'h451434e2, 32'h42ba02d7, 32'h434c05d2},
  {32'hc40cb579, 32'hc268fb48, 32'hc3e080d4},
  {32'h43f7f540, 32'hc3ec69ad, 32'hc25c951d},
  {32'hc32ac7c4, 32'h42b1e89f, 32'hc28f03a3},
  {32'h451d4dcd, 32'h42212e52, 32'hc4005806},
  {32'hc42cf27e, 32'hc2db167e, 32'h429825f7},
  {32'h44fd3e88, 32'hc187ffc7, 32'hc2701006},
  {32'hc4ce5cc6, 32'hc3ce0e3e, 32'h439547d8},
  {32'h44069428, 32'h43e1aa15, 32'hc2e0787e},
  {32'hc4fc9407, 32'hc2799e17, 32'hc39b9262},
  {32'h450080ba, 32'hc39118d9, 32'hc243daa3},
  {32'hc364a870, 32'h43d6da82, 32'h42dc36ea},
  {32'h444e97bd, 32'hc3104a19, 32'hc39a979f},
  {32'hc2844fa0, 32'h4352c755, 32'h43caa4c4},
  {32'h43bbff00, 32'h431236d5, 32'h41ef1266},
  {32'hc4bbb05f, 32'h4358e052, 32'h43283dcd},
  {32'h42ba3bb4, 32'h3ff23d62, 32'h4275b207},
  {32'hc48e2051, 32'h43836f74, 32'hc2abc65b},
  {32'h44d36a60, 32'h41c82868, 32'h4313b5b4},
  {32'h435d81f0, 32'h431921e7, 32'hc329c5d0},
  {32'h44d7509a, 32'hc2799bae, 32'hc22bddcf},
  {32'hc38dd9b4, 32'h41b8ec16, 32'h426cbdb2},
  {32'h441e7ed9, 32'h41d18213, 32'hc3487281},
  {32'hc379aca8, 32'hc181cfc4, 32'h4377d1db},
  {32'h44c868bc, 32'hc131ba86, 32'hc267dc78},
  {32'hc48238f8, 32'h428b83ef, 32'h43b70fb4},
  {32'h44885b97, 32'hc27c7af4, 32'h40c4fae5},
  {32'hc50c0a2e, 32'h42c7d6c8, 32'h42993d8f},
  {32'h44ece620, 32'hc2ade32b, 32'h4379e8f0},
  {32'hc39217a2, 32'hc3657473, 32'h41c47daa},
  {32'h42e43510, 32'hc34af361, 32'hc358de76},
  {32'hc4f4233a, 32'h43e45f18, 32'h420b1a15},
  {32'h44e04fc8, 32'hc3cc0e35, 32'h42827f4a},
  {32'hc4c00378, 32'hc37799a6, 32'hc29cca5c},
  {32'h43989268, 32'hc3afd463, 32'h424c245f},
  {32'hc4ca3621, 32'hc3a255c5, 32'hc3fdad47},
  {32'h44f3b3c0, 32'h43a04b6b, 32'hc13ed19e},
  {32'hc3ba3104, 32'hc3a1e745, 32'h420cabc6},
  {32'h44dfc4e5, 32'h42b31e81, 32'hc34ec60f},
  {32'hc48ef205, 32'h435ce3be, 32'h43905969},
  {32'h44430616, 32'h4288d78c, 32'hc396b93a},
  {32'hc31b1825, 32'hc3b0f01c, 32'hc3acc555},
  {32'hc30d0418, 32'hc34748e2, 32'hc1d8ac94},
  {32'hc4349ec8, 32'hc317a3c9, 32'hc3a96822},
  {32'h44ca0c55, 32'h43d25896, 32'h43669b4e},
  {32'hc468c72b, 32'hc31d31c3, 32'hc33c63e6},
  {32'h44ebeb1f, 32'h41e8a1be, 32'h4286b75a},
  {32'hc48eafd7, 32'hc20022f7, 32'hc2bcfacf},
  {32'h44a85544, 32'h4181a0d1, 32'hc2083c02},
  {32'h4208a9c8, 32'h432e9cf2, 32'h43ae107a},
  {32'h451e7cb4, 32'h42bd27ec, 32'hc376a9bb},
  {32'hc49c3a2f, 32'hc1549669, 32'h42c40bf7},
  {32'h44f2df65, 32'h43152a95, 32'hc37f96ac},
  {32'hc41dab56, 32'hc3900970, 32'hc2d98283},
  {32'h445d6d28, 32'h43b95027, 32'hc3de90ad},
  {32'hc4bfa230, 32'h429f13c2, 32'h4309ba9f},
  {32'h44567dea, 32'h43baf7b6, 32'hc2b1b170},
  {32'h42447790, 32'hc14e94a6, 32'h413cd80c},
  {32'h44bcddba, 32'hc2938e77, 32'hc38725fe},
  {32'hc4ab38e7, 32'hc1a5e370, 32'hc39d43df},
  {32'h4454ec0f, 32'h422ff0b0, 32'hc36562b7},
  {32'hc44c734b, 32'hc2d5a056, 32'hc0727e06},
  {32'h4414f1ca, 32'h42dd013d, 32'hc348a6d6},
  {32'hc440ab4e, 32'h4365dffa, 32'hc3377f65},
  {32'h439a1c22, 32'h40471ca5, 32'h43114411},
  {32'hc4ac31c7, 32'h42db4e13, 32'hc3093c64},
  {32'h435fb2e0, 32'hc28123dc, 32'h42934dda},
  {32'hc500c996, 32'hc2ff5b21, 32'hc2ca3bf2},
  {32'h4509e302, 32'hc391d216, 32'h42dafdbf},
  {32'hc42bbeb6, 32'h43225af1, 32'hc277ccbc},
  {32'h44934ce8, 32'hc2d0565d, 32'hc2b16da3},
  {32'hc4c24c13, 32'hbff345bf, 32'h432adda4},
  {32'h43e28c2d, 32'hc20bca8d, 32'h42fd3121},
  {32'h43ad11c8, 32'hc3c0c1ee, 32'h42e963b5},
  {32'h4503f6ee, 32'h439499bb, 32'h438ff1b8},
  {32'hc4b57584, 32'h434c5c8a, 32'h430d854b},
  {32'h44a46f0d, 32'h42486ecc, 32'h4351fb3e},
  {32'hc4916ef8, 32'h42505f9a, 32'hc377071a},
  {32'h44f1014a, 32'hc3a93ec4, 32'hc3381a4e},
  {32'hc4c647d4, 32'hc0b4c89c, 32'h41eb65b6},
  {32'h437f04c8, 32'h43bf4456, 32'h436ca97d},
  {32'hc50ae077, 32'hc2dc0a55, 32'h42247a14},
  {32'h44f972e6, 32'h43b9d40e, 32'hc2d68f6e},
  {32'hc4a3b113, 32'hc376fffa, 32'h430f3eff},
  {32'h448cdb2d, 32'hc3dbf9af, 32'h42ac6034},
  {32'hc4c7236b, 32'hc3645de4, 32'h427fcfc9},
  {32'h442592a4, 32'hc3687971, 32'hc2964413},
  {32'hc491f616, 32'h43d7af0d, 32'h4298b010},
  {32'h43f0da30, 32'h43c835f2, 32'h42bb53cf},
  {32'hc4def654, 32'hc360b691, 32'h439e0eda},
  {32'h44b39dc8, 32'hc049afc0, 32'hc243ba26},
  {32'hc46ee454, 32'h437f8a43, 32'h42173fec},
  {32'h44fa418d, 32'hc2b9b148, 32'h43a1c959},
  {32'hc4293156, 32'h433fe2db, 32'hc36cc445},
  {32'h43d7d823, 32'hc1bf43e8, 32'hc3be83a8},
  {32'hc4702f61, 32'h43618303, 32'h4323e36b},
  {32'h44bba55d, 32'hc3a5c320, 32'h42dae283},
  {32'hc45c5f53, 32'h41474f49, 32'hc38228fb},
  {32'h44c6fb1e, 32'h42c97ccd, 32'hc31646a6},
  {32'hc4e1e4e8, 32'h439d7e0c, 32'hc0a3b418},
  {32'h44a27b13, 32'h434a050a, 32'h42afef78},
  {32'hc401a4dc, 32'h42271102, 32'hc295577d},
  {32'h4426cf18, 32'hc312fcd0, 32'h439eaa45},
  {32'hc401995c, 32'h437c5735, 32'h43eccbfe},
  {32'h44e1fb14, 32'h4166d602, 32'h43446cd0},
  {32'hc450b2fa, 32'h43296f1b, 32'hc3605523},
  {32'h42c95df4, 32'h43a4c7b5, 32'hc2a7089c},
  {32'hc42975dd, 32'h437efcb8, 32'hc377bd18},
  {32'h4488d71a, 32'h438fff0d, 32'h437351bd},
  {32'h43003804, 32'hc2b8ac63, 32'hc2c5d2ed},
  {32'h441c4d26, 32'hc23d1b96, 32'h416a05a6},
  {32'hc4a2af33, 32'hc2cc67f5, 32'hc2e4ba29},
  {32'h44ac8540, 32'hc36ebb77, 32'hc232d41d},
  {32'hc4c0ccdf, 32'hc28a6bf1, 32'h4348af3a},
  {32'h441c4932, 32'h41627abd, 32'h426b3cac},
  {32'hc3023aa0, 32'hc3df100b, 32'h43b0d960},
  {32'h43a33ad0, 32'h43823b9e, 32'h43057df7},
  {32'hc3ca9970, 32'hc313cbd9, 32'hc3229e1c},
  {32'h44eb27a0, 32'hc2705bfb, 32'hc3347b0a},
  {32'hc46a83c2, 32'hc2cf04e1, 32'h431aafd2},
  {32'h445c4227, 32'h43167cb0, 32'hc3461594},
  {32'hc4d6f5bc, 32'h42bef08b, 32'hc25b5a78},
  {32'h426c0ac0, 32'hc33cf404, 32'h43cdbc6e},
  {32'hc3e8fe58, 32'h42ec1d2c, 32'hc2914a40},
  {32'h44ea0d86, 32'h41eb4ce2, 32'h4116d1e6},
  {32'hc4454fd3, 32'h43099443, 32'h434513f2},
  {32'h450720f6, 32'hc3c99590, 32'h430cb065},
  {32'hc4580eb8, 32'h43373db0, 32'h42aa5bcc},
  {32'h43929ab8, 32'h43930577, 32'hc31d2632},
  {32'hc3f0cbf8, 32'h42c96080, 32'hc2d9f291},
  {32'h44820290, 32'hc1bd1ff4, 32'hc21c5631},
  {32'hc4fe16de, 32'h42f09209, 32'h4357a75a},
  {32'h44d31df1, 32'h4327e036, 32'h43620a96},
  {32'hc397b1fc, 32'hc26fffe1, 32'hc2f2d832},
  {32'h44a2a3bc, 32'h423d01be, 32'hc2319b1a},
  {32'hc1cdbf18, 32'h42d31b59, 32'h431838d0},
  {32'h44ee8ea0, 32'hc2ef9aa6, 32'h42999f32},
  {32'hc4544396, 32'hc2c70027, 32'h416b433b},
  {32'h446789d1, 32'hc2b69de7, 32'hc2f3dcf4},
  {32'hc4bf8659, 32'h43500a15, 32'h42550833},
  {32'h44ccb456, 32'hc435cd7d, 32'h4369669b},
  {32'hc32946e0, 32'hc345f644, 32'hc24e3453},
  {32'h44da97f3, 32'h4354e243, 32'hc3ecd9d6},
  {32'hc4777d68, 32'h431fb1ef, 32'h42d8eed7},
  {32'h450aaebd, 32'h42a33d48, 32'hc3e49ad5},
  {32'hc4955ca0, 32'h419e2e4a, 32'h43d131b3},
  {32'h44bdeccf, 32'hc326698a, 32'hc37ebb2e},
  {32'hc38773e5, 32'h42c572a1, 32'hc31ce9af},
  {32'h44c09cbf, 32'h43026a2c, 32'h42c8c303},
  {32'hc47bad02, 32'hc34ee0b3, 32'hc35fd477},
  {32'h44d155e6, 32'h404e38a7, 32'hc249ab4b},
  {32'hc4b38286, 32'hc290e86e, 32'h40da0738},
  {32'h44a3986f, 32'hc36ae14d, 32'h43271e93},
  {32'hc4d45bc5, 32'h41764d7e, 32'h430410d3},
  {32'h4367ccf2, 32'hc02a7e49, 32'h439b498b},
  {32'hc504c0b8, 32'h43300164, 32'hc2de3752},
  {32'h43967ee6, 32'hc41da9d8, 32'hc3a9db1d},
  {32'hc4eb763e, 32'h438d67c2, 32'hc099c3dc},
  {32'h44846053, 32'h42f0b2e8, 32'hc3c30eba},
  {32'hc4427d06, 32'h43e25d2b, 32'hc31ecdf6},
  {32'h44af92a3, 32'hc2235497, 32'hc2accbd5},
  {32'hc4913fa0, 32'hc23eebca, 32'h43087670},
  {32'h45103ca4, 32'hc420b8a1, 32'hc1c57faf},
  {32'hc32bedc8, 32'hc394b1ef, 32'h4103ed57},
  {32'h44f04f1c, 32'h43ca68f4, 32'hc34d8474},
  {32'hc3f20618, 32'h43b94b52, 32'h43553bb3},
  {32'h4492c379, 32'hc1c5de69, 32'hc2df4efc},
  {32'hc3e3c3f0, 32'hc353f7b6, 32'h4349e44c},
  {32'h42aacc30, 32'hc2c74aa4, 32'h431cdc42},
  {32'hc340d8f8, 32'hc37671e8, 32'hc1bbcc4e},
  {32'h44f1d611, 32'hc1709271, 32'h41c9e4a0},
  {32'hc4a12652, 32'hc306dbad, 32'hc15fb9e9},
  {32'h449f8513, 32'hc34faa36, 32'h430956cb},
  {32'hc4b6873f, 32'h43e7befb, 32'h428a71c6},
  {32'h447912fb, 32'hc301ffa1, 32'hc3a86c2e},
  {32'hc4cbb81e, 32'hc3866e07, 32'h42920fb2},
  {32'h438ac6dc, 32'hc30f7ea7, 32'h43390f74},
  {32'hc43a3560, 32'h43002a90, 32'hc3d63824},
  {32'h448cf700, 32'hc3bc697c, 32'hc35ad2bc},
  {32'hc4842ba0, 32'h42797b45, 32'hc3822f34},
  {32'h45045eab, 32'hc354d6cc, 32'hc23dfb30},
  {32'hc4dacf79, 32'hc0eeb2a8, 32'hc2923b7d},
  {32'h44a5cc9c, 32'h42f215b3, 32'hc15241ec},
  {32'hc4b21cd0, 32'hc338ee62, 32'hc216c763},
  {32'h44f9bebd, 32'hc2e0dc52, 32'h4245ae1a},
  {32'hc494156a, 32'hc2c1d492, 32'h41edd80b},
  {32'h441a4107, 32'h41e394d1, 32'hc21148ee},
  {32'hc4e44651, 32'h430bfd24, 32'h434ff06d},
  {32'h42ce5a60, 32'h40c8954c, 32'h42fd7c2e},
  {32'hc4f5994f, 32'hc2ba164c, 32'hc2957540},
  {32'h44c30f17, 32'h4328c092, 32'h43a3c4aa},
  {32'hc49dde82, 32'h43805a94, 32'h43b6550f},
  {32'hc2e132c0, 32'hbfcddbb0, 32'h434c2fb1},
  {32'hc4f82631, 32'hc388a17d, 32'h438268cf},
  {32'h44eea92e, 32'h42ce617e, 32'hc304dc83},
  {32'hc4d73ac6, 32'h42b60367, 32'hc134d8bd},
  {32'h450a61a0, 32'h43b572ea, 32'h420558e3},
  {32'hc3f846ac, 32'h4276137f, 32'h43118224},
  {32'h447a2a45, 32'h41ff32c5, 32'h43cf709a},
  {32'hc4cc4c97, 32'hc2fdac32, 32'h4347c56d},
  {32'h4510ae07, 32'h4287072f, 32'h43492282},
  {32'hc4a6b637, 32'hc17bb4c7, 32'hc32ddd8b},
  {32'h4399d2e0, 32'hc2f9414f, 32'hc3b5256e},
  {32'hc4b0a636, 32'hc3c6f367, 32'h439042b1},
  {32'h44c8b094, 32'h433016f9, 32'hc31ed8f1},
  {32'hc4fe2d90, 32'hc2eccfc2, 32'hc39756f8},
  {32'h43ba15cc, 32'hc2f5aaa3, 32'hc2b426cc},
  {32'hc50ec49d, 32'h41cb8ea5, 32'h438034ab},
  {32'h44864251, 32'hc32a267c, 32'hc37f1310},
  {32'hc49474c7, 32'hc33a017f, 32'h435e394e},
  {32'h43fd9bd2, 32'h4330afc0, 32'h4395b073},
  {32'hc50c5d15, 32'hc30f2791, 32'h4428e34c},
  {32'h44c8d24a, 32'h42aa7756, 32'h430b464b},
  {32'hc4206222, 32'hc1c8a1b8, 32'h432dfc26},
  {32'h43f05f9b, 32'hc3212ff6, 32'h44001248},
  {32'hc502c54d, 32'h42832515, 32'hc2fb89bf},
  {32'h44d7c524, 32'h42968a85, 32'hc1c49b41},
  {32'hc4a886ee, 32'hc36327da, 32'hc34a101c},
  {32'h44ee0910, 32'h430f685a, 32'h4366f7d9},
  {32'hc4df63f5, 32'h431527c0, 32'h4386cc43},
  {32'h44ec1e79, 32'h42aff0c1, 32'hc39a33a2},
  {32'hc38d0fff, 32'hc3632549, 32'hc444ecba},
  {32'h448758bb, 32'hc38134e1, 32'hc28a04a8},
  {32'hc48623fc, 32'hc3354519, 32'hc29b9223},
  {32'h4506e9d5, 32'h439e7d3f, 32'h42d132fc},
  {32'hc45f4478, 32'hc356a475, 32'hc300785e},
  {32'h4161c9f0, 32'h40d32f22, 32'h4340a006},
  {32'hc49d5b9e, 32'hc2d402d2, 32'hc3992a69},
  {32'h43282eb0, 32'h4373e60c, 32'hc2dee03a},
  {32'hc4e8a232, 32'h42e752ed, 32'hc16085bd},
  {32'h45171f8f, 32'hc3a45d58, 32'h439a42cb},
  {32'hc44cb358, 32'h434cf412, 32'hc071b2f8},
  {32'h43809c10, 32'h43042300, 32'hc304c358},
  {32'hc509260a, 32'hc324bedc, 32'hc36f10d5},
  {32'h448d20d0, 32'h43bf8aef, 32'hc3b73b4b},
  {32'hc4bcfd28, 32'h403f9806, 32'h43038273},
  {32'h43601f7a, 32'h42dbaf1d, 32'hc3ce5919},
  {32'hc388753b, 32'h42aeb4df, 32'hc39074d6},
  {32'h43a6236d, 32'h41ab5c8f, 32'hc31c42b6},
  {32'hc432581c, 32'h43895a70, 32'h42488816},
  {32'h442b7c9c, 32'hc2764a38, 32'hc249ce94},
  {32'hc49a08cb, 32'hc3203e78, 32'h41fc8cb8},
  {32'h44179de6, 32'h43249010, 32'hc2c88bc8},
  {32'hc52911b9, 32'h4375a2a3, 32'hc2f81480},
  {32'h43ada484, 32'hc3c96f96, 32'h434f6962},
  {32'hc4de2c20, 32'hc2ebe18e, 32'hc3b85cee},
  {32'h441cca2b, 32'hc0615dac, 32'hc3da26e7},
  {32'hc4474740, 32'hc361be00, 32'h413f72e2},
  {32'hc27c8080, 32'hc3df5217, 32'h43369810},
  {32'hc48b5b40, 32'h43133a40, 32'h438d8bdd},
  {32'h440aa6fc, 32'hc3c80b3a, 32'h42849576},
  {32'hc4d1fe26, 32'hc38ae631, 32'hc1f583eb},
  {32'h4409c3ba, 32'h4160c92e, 32'hc1fb73b4},
  {32'hc38a5c2a, 32'hc39830c1, 32'h431dfb4a},
  {32'h44d68133, 32'hc2da74ac, 32'h42a67b51},
  {32'hc3563090, 32'h4299b9b9, 32'h43ce1030},
  {32'h440814bc, 32'hc142b9c1, 32'h4337dc18},
  {32'hc49ed82f, 32'h431030a0, 32'h430b6a75},
  {32'h4488a61a, 32'h42fc4c12, 32'hc38244fa},
  {32'hc46a4b00, 32'hc34d7869, 32'hc31506eb},
  {32'h4476975f, 32'hbfc4a239, 32'h40262558},
  {32'hc4f7226c, 32'hc31a0342, 32'h43158726},
  {32'h44344246, 32'hc33e4704, 32'hc2804d6a},
  {32'hc50b3555, 32'hc1fcaf6e, 32'hc32f4494},
  {32'h441a6338, 32'h4352e4ad, 32'hc38e24dc},
  {32'hc46a6032, 32'hc3acb13b, 32'h43352f8d},
  {32'h44f3786b, 32'h431e9704, 32'h411cea6b},
  {32'hc3900a50, 32'h42736001, 32'hc352d8c0},
  {32'h45135bdf, 32'hc0e3eae8, 32'hc2877112},
  {32'hc4e35532, 32'hc3abbb39, 32'h42a2f97f},
  {32'h44bff077, 32'hc34e9fa5, 32'h42935e6f},
  {32'hc509794e, 32'hc3c6dfae, 32'hc3a733b5},
  {32'h448fddfd, 32'hc2f6927e, 32'hc3ef9e2c},
  {32'hc4b8e02a, 32'hc2d79cdc, 32'hc2704002},
  {32'h4418f103, 32'h42091c2b, 32'hc3c91450},
  {32'hc4e6674d, 32'h42cd783f, 32'h43a65c39},
  {32'h44884eb5, 32'hc1d35487, 32'hc38e62f3},
  {32'hc48bebed, 32'hc34533f0, 32'h43b58f93},
  {32'h451b2385, 32'h432b4930, 32'h429fa9a8},
  {32'hc50f6dbe, 32'hc32a6138, 32'hc3ae50ac},
  {32'h44b35593, 32'hc168b164, 32'hc2fceb52},
  {32'hc4d02a19, 32'hc3758a2d, 32'h426a1d8d},
  {32'h452f855d, 32'hc280ceba, 32'hc199b38b},
  {32'h4269a960, 32'h42ac5e54, 32'hc34cf8d6},
  {32'h44d76ff6, 32'hc2eab84c, 32'h432e86bf},
  {32'hc4af9502, 32'hc2950c41, 32'hc24e1884},
  {32'h44a72176, 32'h42ecdc71, 32'h437a8c14},
  {32'hc4034440, 32'hc32dd67a, 32'hc3c5f2cb},
  {32'h442818a6, 32'hc3e29e1c, 32'h428fa201},
  {32'hc4c09def, 32'hc28e2b32, 32'h43b3ce0e},
  {32'h44da8fa8, 32'h4353b265, 32'hc3be1139},
  {32'hc3a1b363, 32'hc2f672d1, 32'h423de65f},
  {32'h44dd56f8, 32'hc27f02b4, 32'hc2df7249},
  {32'hc3ae85ba, 32'hc3dea0f3, 32'hc2829726},
  {32'h43158058, 32'h43971211, 32'h436f71be},
  {32'hc407a7a4, 32'hc261c688, 32'h424a9b9c},
  {32'h44828aa7, 32'h42fa5ebb, 32'h4263690b},
  {32'hc51b1a3d, 32'hc08bd7c8, 32'hc3acee34},
  {32'h44aea726, 32'h427f8081, 32'hc1a3bf01},
  {32'hc3f49684, 32'hc2dee612, 32'h420155e3},
  {32'h450c0666, 32'h420b0818, 32'hc31a6ed0},
  {32'hc4390306, 32'h432d7978, 32'hc37c9cf5},
  {32'h44847cce, 32'hc380d5e4, 32'hc3df861e},
  {32'hc333a4f8, 32'h43759492, 32'h42a82eba},
  {32'h4382a718, 32'h43b559f8, 32'hc3d3bf7f},
  {32'h43278d18, 32'hc303a8de, 32'hc3a53816},
  {32'h44f98ff4, 32'hc30f32aa, 32'h430e4c36},
  {32'hc1034b00, 32'hc3deed1c, 32'hc399bfdf},
  {32'h44f508f6, 32'hc37c6deb, 32'hc3b27bcf},
  {32'hc4f050a4, 32'h4282ffe1, 32'hc3891ba5},
  {32'h4522d308, 32'h440bcb9d, 32'h4301e6ad},
  {32'hc512e2a5, 32'h4334b529, 32'h4323c580},
  {32'h4416c37c, 32'h42702991, 32'h42b01a42},
  {32'hc46cd8a3, 32'hc2ecea5c, 32'hc2de8f57},
  {32'h443c6c10, 32'hc35d2af4, 32'hc2ec45f8},
  {32'hc2e7adc0, 32'h3faf9c30, 32'hc399e013},
  {32'h4503d9a4, 32'hc3439744, 32'hc393bd08},
  {32'hc38c8dc0, 32'hc3a0662f, 32'hc3c74e38},
  {32'h43d860d2, 32'h42ecfb7c, 32'h435fbe88},
  {32'hc423dc5d, 32'h42933e58, 32'hc397da7e},
  {32'h447b50c1, 32'hc36d275f, 32'h43b20220},
  {32'hc49abcc6, 32'hc1a936f9, 32'hc3d3b915},
  {32'h43e869f8, 32'h433beddc, 32'h42e94c4d},
  {32'hc4d938f4, 32'hc009bb80, 32'hc3108172},
  {32'h44b71a2f, 32'hc3607a83, 32'h42bfe531},
  {32'hc493af44, 32'hc3884c27, 32'h42f387c8},
  {32'h448f149e, 32'h4360a7b4, 32'h4313b8cf},
  {32'hc4f3a2e7, 32'hc383d318, 32'hc30f12ea},
  {32'h44d5e056, 32'h4205a9de, 32'hc30c41ae},
  {32'hc3c429ea, 32'hc3b0acdf, 32'h4297a606},
  {32'h43eb9839, 32'h436f800c, 32'hc0d7590f},
  {32'hc3dd2623, 32'hc32984fc, 32'hc1a9fff1},
  {32'h43ba9908, 32'h43c39cb4, 32'h435d36d2},
  {32'hc2f25430, 32'hc3899ede, 32'hc2211a80},
  {32'hc4091058, 32'hc350c8c2, 32'h4340f952},
  {32'hc28c8f8c, 32'hc2a35a82, 32'h42bc9a1f},
  {32'hc47a3441, 32'hc38e1c43, 32'hc138baf4},
  {32'h44ac26b8, 32'hc2ea1093, 32'h435b4c79},
  {32'hc5075830, 32'h4273a828, 32'hc38227c8},
  {32'h4426dd82, 32'h429d5279, 32'h4332c2ed},
  {32'hc475d09a, 32'h433cac80, 32'hc20b73d6},
  {32'h44eceae3, 32'h43f0c48a, 32'hc2f6f728},
  {32'hc4b8dbfe, 32'h430a4327, 32'hc3bc84fc},
  {32'h44d134bb, 32'hc3aea789, 32'h436e2cc1},
  {32'hc3b6d5ce, 32'h43564727, 32'hc1e558c9},
  {32'h44db27de, 32'h43b94a0f, 32'hc3888bb8},
  {32'hc2528f70, 32'hc2bb0190, 32'h431592e0},
  {32'h44614a66, 32'hc25430ef, 32'h431df599},
  {32'hc4f5b15c, 32'h42cf5ca0, 32'h4305f8ac},
  {32'h44184805, 32'h41a58557, 32'hbfc92810},
  {32'hc4b8ca52, 32'h433d5c74, 32'hc2a5f370},
  {32'h4474ae9e, 32'h43739b91, 32'h43689919},
  {32'hc489dc4c, 32'hc31da240, 32'h409a581e},
  {32'h44ac2028, 32'hc3841a7a, 32'h43869c93},
  {32'hc4126bc4, 32'hc39304c8, 32'hc35d9548},
  {32'h43f7ee60, 32'hc3bcb6c1, 32'hc3169f73},
  {32'hc3a2b480, 32'hc304b68d, 32'h4330bbad},
  {32'h431c4d3b, 32'h42787b0f, 32'h4352a569},
  {32'hc4d28519, 32'hc24f18e7, 32'hc38dd7da},
  {32'h450a2288, 32'h4030fcf8, 32'h435fa278},
  {32'hc4c4a758, 32'hc39d242f, 32'hc29db656},
  {32'h44f2bf9a, 32'h40dcc6e1, 32'h431f8d5d},
  {32'hc4f0c7f1, 32'hc2826720, 32'hc3af871b},
  {32'h44743520, 32'h432befbb, 32'hc1f8e932},
  {32'hc49e31c5, 32'h428ba609, 32'hc30ba990},
  {32'h44966c8c, 32'h420b9d00, 32'hc1cda534},
  {32'hc46953f2, 32'hc3855850, 32'hc30dad75},
  {32'h450537be, 32'h428b0b5d, 32'h434096ba},
  {32'hc516599d, 32'h4349650e, 32'hc36bc739},
  {32'h4500960c, 32'h42a6bb08, 32'hc0f9425c},
  {32'hc507dd0b, 32'h4293df88, 32'hc23f307a},
  {32'h438c1bd0, 32'h4335f01c, 32'h437cda9c},
  {32'hc43666f9, 32'hc3876577, 32'h42d27d47},
  {32'h44858d7d, 32'hc36bc625, 32'hc12e2f0c},
  {32'hc4310f73, 32'hc3546f84, 32'hc3122a42},
  {32'h45048fc4, 32'h43348312, 32'h439aa9d4},
  {32'hc45ae0a0, 32'h43194db9, 32'h428e6a92},
  {32'h4518ee8c, 32'h43184624, 32'h4338122b},
  {32'hc4fc4461, 32'h43a52573, 32'h43c4d042},
  {32'hc0f31880, 32'h425acc41, 32'h43a4fccf},
  {32'hc4a602c8, 32'h42bc6b5e, 32'h4232afdd},
  {32'h4505e924, 32'h42bf09c4, 32'hc3c2aaf9},
  {32'hc3d8c950, 32'hc207d198, 32'h43af185a},
  {32'h449ff31e, 32'hc2792392, 32'h42f5d755},
  {32'hc4ca750e, 32'h443edd64, 32'hc207daa4},
  {32'h45165524, 32'h436748dd, 32'hc326fdd3},
  {32'hc40b0a44, 32'hc3b794e8, 32'h42c7754b},
  {32'h4321f058, 32'hc3c16a67, 32'h43433db2},
  {32'hc4ac7b53, 32'hc228852d, 32'hc3a48ef7},
  {32'h445d0491, 32'hc3027b82, 32'hc41e2998},
  {32'hc34a4dc8, 32'hc332defb, 32'hc38a5326},
  {32'h450656af, 32'hc2547324, 32'hc3be598c},
  {32'hc49450d9, 32'hc31cb9ba, 32'hc349defa},
  {32'h44900992, 32'hc2498cdc, 32'h43133a7c},
  {32'hc5053ca5, 32'hc309921e, 32'h42b5c3c5},
  {32'h423be5e4, 32'h4381ec27, 32'h439e8e0b},
  {32'hc398b638, 32'h42d75083, 32'h43446623},
  {32'h44df3c11, 32'h42439812, 32'h421c7269},
  {32'hc3a8fed8, 32'h42148b9e, 32'h432ac146},
  {32'h43235c50, 32'hc444234c, 32'hc225c14e},
  {32'hc1fece80, 32'hc1851fdb, 32'hc3b0cb06},
  {32'h449b1f87, 32'h43ad56b3, 32'hc38c0283},
  {32'h4280ea0e, 32'hc365cbe4, 32'hc3acac0a},
  {32'h4436f3ce, 32'hc2880958, 32'h438381f6},
  {32'hc51b8cb8, 32'h4358981f, 32'h432bc3c1},
  {32'h44e8122c, 32'hc3fab786, 32'h41cd66b2},
  {32'hc4f08394, 32'hc19191a7, 32'hc217db77},
  {32'h44c2fa8a, 32'h41c1728d, 32'h4332432c},
  {32'hc41c919c, 32'hc30eda7e, 32'hc2abb806},
  {32'h447f992a, 32'h411e2fa0, 32'h427f9af2},
  {32'hc3c6de50, 32'hc1350ebc, 32'hc12b4e80},
  {32'h44dc9e5a, 32'h42d80e3d, 32'h42b0d788},
  {32'hc389709c, 32'hc1dccfcd, 32'h4378f677},
  {32'h448fdf52, 32'hc17e09f5, 32'h438ac80d},
  {32'hc3927c6c, 32'h430629b5, 32'h427759e4},
  {32'h44e491d6, 32'hc3a63946, 32'hc2fab162},
  {32'hc1c29048, 32'hc32d1863, 32'hc3642dc7},
  {32'h44b34aca, 32'h433371fc, 32'hc2bbc4a6},
  {32'hc5206502, 32'hc39528a7, 32'h409a84ea},
  {32'h44540f00, 32'hc2e5eec7, 32'h40842a66},
  {32'hc39bd24f, 32'h43cae3c7, 32'hc352bb0a},
  {32'h44e5852f, 32'hc3527bf5, 32'hc328962a},
  {32'hc4efd7e7, 32'hc3e99038, 32'h439faf5e},
  {32'h44a386e5, 32'h418d48f8, 32'h42852924},
  {32'hc44b22ab, 32'hc36f089a, 32'hc1aaacd1},
  {32'h44e38fe0, 32'hc1eae4ae, 32'hc1f3a428},
  {32'hc42f70bc, 32'h43bf9a79, 32'h4381d802},
  {32'hc2231794, 32'h4208753d, 32'h43807d3c},
  {32'hc49dfe54, 32'h432bb9e0, 32'h42500532},
  {32'h4462948c, 32'hc34f0085, 32'hc38adb46},
  {32'hc43a0b56, 32'h440f08ff, 32'h43338f47},
  {32'h448f1c97, 32'hc2f8dbea, 32'h430544c2},
  {32'hc5087907, 32'h43395a21, 32'hc22d617c},
  {32'h44a927a3, 32'h439880f9, 32'h440eb13d},
  {32'hc50ba339, 32'h439267b5, 32'h437a7670},
  {32'h44e0c2b2, 32'h42b30d61, 32'h418e5d83},
  {32'hc42ebf58, 32'hc299c27e, 32'h430687ad},
  {32'h44884339, 32'h43e61c0a, 32'h43b3a0dc},
  {32'hc47c685c, 32'hc3a0e11a, 32'h436870f5},
  {32'h44073406, 32'hc36c7fdf, 32'hc35e5b45},
  {32'hc4cfd235, 32'hc36cb3a6, 32'h41c88697},
  {32'h4514c0df, 32'hc373f610, 32'h434c38a0},
  {32'h40c91960, 32'h43cc940c, 32'hc3e1e561},
  {32'h4461ebfc, 32'h432aaed7, 32'hc35a3e0b},
  {32'h42a7f800, 32'hc186fec8, 32'h42f6ad33},
  {32'h450c77cc, 32'h4301f81b, 32'hc31111d4},
  {32'hc4e1aafa, 32'h43aa90d7, 32'hc387bfa4},
  {32'hc29177d8, 32'hc3733a42, 32'h43aaa874},
  {32'hc52b3ba2, 32'hc38ef164, 32'hc1d61a5a},
  {32'h44ba8d3f, 32'hc3d416ad, 32'hc38330a1},
  {32'hc3cd9377, 32'hc3a1bdcb, 32'hc1907425},
  {32'h44b93c07, 32'h4289ca83, 32'hc290c4ae},
  {32'hc4e75fd9, 32'hc388e6fb, 32'h43b06a76},
  {32'h44ab2b0a, 32'h4300bbba, 32'h429523b6},
  {32'hc4ff0473, 32'hc2781b40, 32'h4282f9ea},
  {32'h450c8902, 32'h42ef8fc1, 32'hc319b27e},
  {32'hc5099114, 32'h436531a6, 32'h43a65188},
  {32'h4425ce76, 32'hc2ce07a7, 32'h430fe9a8},
  {32'hc4dc8c74, 32'h42811b42, 32'hc30c7b15},
  {32'h450581e4, 32'h42c4a2d1, 32'hc3d3aeb2},
  {32'hc5037940, 32'hc393c504, 32'h42172635},
  {32'h4415e28a, 32'h43e507dc, 32'hc31a1cd7},
  {32'hc4b38a0b, 32'hc367df09, 32'hc388beee},
  {32'h451e87a4, 32'hc26f2b1a, 32'h424c2e57},
  {32'hc4ecce3d, 32'hc4048873, 32'h434305f4},
  {32'h4410e0c3, 32'h42024a05, 32'hc2c8a813},
  {32'hc4af26a0, 32'h439b3c18, 32'hc4001b00},
  {32'h44953208, 32'hc2d91508, 32'hc1cbb513},
  {32'hc5115c45, 32'hc3c2710c, 32'h438109fe},
  {32'h4354a452, 32'h42517b44, 32'hc35dac0a},
  {32'hc45a0e23, 32'hc37fa89a, 32'h42bdc83b},
  {32'h44fb8148, 32'h431e227a, 32'hc2904af4},
  {32'h4293c8a0, 32'hc33beb8a, 32'hc30b3cd6},
  {32'h44e69282, 32'h424465b5, 32'hc28c74c5},
  {32'h4368ab24, 32'h421812e1, 32'h43587d30},
  {32'h44fd9098, 32'hc3349b65, 32'h42390f8f},
  {32'hc3fd2860, 32'hc3af4321, 32'hc2a96d8c},
  {32'h45013371, 32'hc2799d15, 32'hc381c071},
  {32'hc5016bef, 32'hc3460173, 32'hc1e1e036},
  {32'h43bf6478, 32'hc1baf609, 32'h438f91cb},
  {32'hc51664d7, 32'hc403416c, 32'h431b7776},
  {32'h441e1fa7, 32'h437115ce, 32'h421206fb},
  {32'hc4f1fffa, 32'hc0dba747, 32'h43938b8c},
  {32'h44b14d96, 32'h4374b7e8, 32'hc3657574},
  {32'hc50f8cb4, 32'h438d39c6, 32'hc2437a1f},
  {32'h44b99d92, 32'hc3a9e1ec, 32'h4388c8a0},
  {32'hc4d5513b, 32'hc192f754, 32'hc2ba57a8},
  {32'h42f32180, 32'hc0fef294, 32'h43923935},
  {32'hc4f9ab06, 32'h3f1a74b8, 32'hc3811f2d},
  {32'h45007662, 32'h438be6cc, 32'h43118d16},
  {32'hc4f176b6, 32'hc299951f, 32'hc37def95},
  {32'h44feee6d, 32'h437e5bd8, 32'hc3d151dc},
  {32'hc4d0b06e, 32'h431d4a22, 32'hc11e6ab0},
  {32'h448224ee, 32'hc2ed9706, 32'hc2b17f92},
  {32'hc3dd06e8, 32'hc3052c8b, 32'hc3bbc47b},
  {32'h45112f76, 32'h42e5f054, 32'h415ef248},
  {32'hc48750a4, 32'hc3362165, 32'hc386a384},
  {32'h440bcc51, 32'hc2bc3272, 32'hc2be2b67},
  {32'hc44cbd11, 32'hc40ab695, 32'hc345f07d},
  {32'h44f5a4b1, 32'h41fcf17d, 32'hc3936ea9},
  {32'hc4c18606, 32'h4317900b, 32'h41e4fd4d},
  {32'h44a388be, 32'h43caa5a1, 32'h43392e1d},
  {32'hc273c678, 32'h42451a96, 32'h4345b17b},
  {32'h44fd3f86, 32'hc2c44ed2, 32'hc241997e},
  {32'hc4982b8a, 32'h41798519, 32'hc3970f3a},
  {32'h44a85408, 32'h42d93599, 32'hc328c040},
  {32'hc3f785aa, 32'h42c68fa9, 32'h42d03072},
  {32'h44e23326, 32'hc3582524, 32'h432527d5},
  {32'hc49c43f5, 32'hc39b15d2, 32'hc313c7ba},
  {32'h44bb6feb, 32'h43ba7b76, 32'h440a6a54},
  {32'hc46f6256, 32'hc27bfba9, 32'hc33a844a},
  {32'h44d5ea25, 32'hc2135ef8, 32'hc389d908},
  {32'hc4c8ee4e, 32'hc332f380, 32'hc41123df},
  {32'h4384e728, 32'hc229ee58, 32'h422cd82e},
  {32'hc402d166, 32'hc3adfc01, 32'h438256ad},
  {32'h441ce773, 32'h41b7caa8, 32'hc19f0644},
  {32'hc41b6e61, 32'hc385e458, 32'h4285b1ca},
  {32'h44b073d9, 32'h41c58942, 32'hc3568165},
  {32'hc4d714e7, 32'hc38d14f2, 32'h42e66db0},
  {32'h4475c1a8, 32'h4306f00c, 32'h42b5d3ed},
  {32'hc4345d19, 32'h4223df96, 32'hc241d5f5},
  {32'h4473bad0, 32'h43a6934b, 32'h4302002f},
  {32'hc4990544, 32'hc30d9413, 32'h43816574},
  {32'h44e8decc, 32'hc31eeb88, 32'h437ce9f1},
  {32'hc4dbd962, 32'hc3a94f38, 32'h41ede600},
  {32'h43a27c14, 32'h43b5c4b6, 32'hc0bbd3f4},
  {32'hc48bdae8, 32'h421f2440, 32'h4229c099},
  {32'h4384c934, 32'h4106a119, 32'h421887a6},
  {32'hc40fac97, 32'hc2e7fccc, 32'hc2b21cee},
  {32'h450f720e, 32'h4176babc, 32'h432cb674},
  {32'hc3adf315, 32'hc2d8d599, 32'hc0595f97},
  {32'h44fc41e5, 32'hc178342b, 32'h436d0e5f},
  {32'hc3ecd05e, 32'hc2d8eb51, 32'hc36df854},
  {32'h438c4e4a, 32'hc30fb92e, 32'h43b5d7e1},
  {32'hc50ca0a5, 32'hc34ed648, 32'h438072bb},
  {32'h44e90f29, 32'hc210d868, 32'hc1bb630a},
  {32'hc3a129d0, 32'hc31786c5, 32'h43dcd52b},
  {32'h44926d23, 32'h430a4310, 32'hc385615f},
  {32'hc4914208, 32'hc34e20ee, 32'h42f6b0ee},
  {32'h450dc2c2, 32'h42e2d9fb, 32'hc2bf0f4f},
  {32'h43b5e008, 32'h4364b608, 32'h4341254d},
  {32'h4323ee7e, 32'hc32625f4, 32'hc33fab60},
  {32'hc5021601, 32'h42c6600b, 32'hc1dc1a49},
  {32'h44eebd12, 32'hc28834d8, 32'h422628ee},
  {32'hc44475aa, 32'h40710251, 32'hc3166487},
  {32'hc2d34130, 32'h439b8dc2, 32'hc1042652},
  {32'hc44be144, 32'h42158901, 32'hc1f06629},
  {32'h4505005e, 32'h422ceb2c, 32'h42b18eb8},
  {32'hc489062f, 32'hc2ed0d92, 32'hc29ec75a},
  {32'h43d82b9b, 32'h43456cd0, 32'h436defdc},
  {32'hc4e463c1, 32'h43370c10, 32'h43731600},
  {32'h44fae290, 32'h435cd404, 32'hc38c3c21},
  {32'hc4d9df42, 32'h42746ed4, 32'hc2cb9b1c},
  {32'h4478ade7, 32'hc1ae0337, 32'h43ad6337},
  {32'hc43e8606, 32'h41ac7f82, 32'h409bb368},
  {32'h446dc504, 32'h4299d457, 32'h4224dae2},
  {32'hc4bf0146, 32'h43a1e9ec, 32'h41b6247e},
  {32'h4504bb7c, 32'h4325bc5d, 32'hc1f60837},
  {32'hc50cf98c, 32'hc243da95, 32'h430029f5},
  {32'h4493140e, 32'hc09c563c, 32'hc3322610},
  {32'hc4fe86df, 32'h4360d2e8, 32'hc43a2e7e},
  {32'h44db2f56, 32'h438c87ec, 32'hc32e1452},
  {32'hc5225546, 32'h4391729f, 32'h43917434},
  {32'h449d5e5a, 32'hc19253aa, 32'hc30196a0},
  {32'hc497796a, 32'h434458ff, 32'h427c0167},
  {32'h43dc2504, 32'h423d8da2, 32'hc3944ec7},
  {32'hc3479cd0, 32'h42b7d61b, 32'h422e3648},
  {32'h45035437, 32'h43466860, 32'h43a3d675},
  {32'hc4e7524b, 32'h42fe2b3b, 32'h4287914e},
  {32'h43ac3c12, 32'h4313422e, 32'h4346c54a},
  {32'hc4b7cfbf, 32'hc320cf13, 32'hc2fe2fde},
  {32'hc29e6e6c, 32'hc384f142, 32'hc38b7524},
  {32'hc45f4466, 32'h4271be1a, 32'h43d32362},
  {32'h43edf458, 32'h43a31b4b, 32'h42d320ba},
  {32'hc5162b7b, 32'h41b6ad44, 32'h423f0c0c},
  {32'h4459cd8f, 32'hc2eb8993, 32'hc24c7d60},
  {32'hc4ddce24, 32'h428200f6, 32'h418609e6},
  {32'h446cf8b2, 32'h43669226, 32'h42de1b79},
  {32'hc34c143c, 32'hc00ec504, 32'h438b8a88},
  {32'h44910b3b, 32'hc1db9035, 32'h43d0de6b},
  {32'hc4ed2dce, 32'h43a23b86, 32'h42ad46d9},
  {32'h447feddb, 32'hc38faf57, 32'hc3719c04},
  {32'hc50d1a62, 32'h435133ed, 32'h42d93411},
  {32'h44f7a885, 32'h43d86eed, 32'hc3fd5637},
  {32'hc461e6b2, 32'h42e9811b, 32'h43442476},
  {32'h44fc075e, 32'hc2b489dc, 32'h43884bb6},
  {32'hc45e20a9, 32'hc37e9514, 32'h426a3926},
  {32'h4468f53c, 32'h41c69204, 32'h42e1c9cc},
  {32'hc4c783ec, 32'hc2a3667f, 32'h42d5fdb8},
  {32'h435e0717, 32'hc3989fbf, 32'hc2df7c3c},
  {32'hc4a74584, 32'hc3371010, 32'hc3461d7a},
  {32'h45123785, 32'hc2c40bb4, 32'hc1e1bab3},
  {32'hc4a12874, 32'h430269b4, 32'hc39a1649},
  {32'h45188b45, 32'hc1552788, 32'hc342fe68},
  {32'hc4ce759f, 32'hc2a3f7eb, 32'h4318dbc7},
  {32'h44edabfe, 32'h42d60d6d, 32'hc2a1b776},
  {32'hc38d9bb4, 32'h427dbb70, 32'hc2c6b0fc},
  {32'h44db97a4, 32'h42c59afc, 32'hc3066683},
  {32'hc4ce3408, 32'h42c2cac8, 32'hc3717c74},
  {32'h44e811b8, 32'hc31d4b53, 32'h4422c156},
  {32'hc4f7414c, 32'hc3943105, 32'h434f26f0},
  {32'h448be566, 32'hc37fc689, 32'hc333e2ed},
  {32'hc4c28ae5, 32'h4206f695, 32'h43b997b3},
  {32'h44e8241f, 32'hc32d7d13, 32'h43200c15},
  {32'hc431df13, 32'h430640ef, 32'hc24e9b0f},
  {32'h44218763, 32'h433991b2, 32'hc2a3f2b0},
  {32'hc3bce73c, 32'h4430e0ad, 32'hc33864d7},
  {32'h44fbd3f8, 32'hc227d13c, 32'hc2b91765},
  {32'hc4e38c67, 32'hc2aa946c, 32'hc2920a8a},
  {32'h4304a8a6, 32'h428ccf80, 32'h42c8e641},
  {32'hc4c19912, 32'h43c8c688, 32'hc26600ea},
  {32'h44a83a47, 32'hc220494f, 32'h4291e064},
  {32'hc4b700a8, 32'h4225c004, 32'hc2de735c},
  {32'h449a6684, 32'h42c6dace, 32'hc2711122},
  {32'hc45d9984, 32'h42d45a98, 32'hc383fd7c},
  {32'h44ef43d6, 32'hc3341866, 32'hc329677f},
  {32'hc4c7bd2a, 32'h433f6d34, 32'hc27ab3f9},
  {32'h44e75b84, 32'hc2babea9, 32'h43fa47e4},
  {32'hc4db5c8a, 32'h42a29472, 32'hbf47bba0},
  {32'h44ad9635, 32'h43c1feec, 32'h42565950},
  {32'hc4aa19b7, 32'h438afcc8, 32'h431edde9},
  {32'h450f4a7c, 32'hc314a873, 32'hc36ca648},
  {32'hc49f4e31, 32'hc3ce92b3, 32'hc3186b86},
  {32'h44154b38, 32'h431d0439, 32'hc3bb92c0},
  {32'hc50f380f, 32'h423b5ccf, 32'h43dfba29},
  {32'h448c3189, 32'hc3c72167, 32'hc362d5b0},
  {32'hc44bd70c, 32'hc2b7b799, 32'hc38e108e},
  {32'h4497e169, 32'h439270e2, 32'h43116cfe},
  {32'hc4b09af9, 32'hc3965107, 32'h42be67cb},
  {32'h440013e2, 32'h424b9f84, 32'h426ec2f0},
  {32'hc48dfe27, 32'hc36a7567, 32'hc39eb491},
  {32'h450b8b62, 32'h42a98b80, 32'h43a7ec6f},
  {32'hc424228c, 32'hc30104f8, 32'hc317ce1d},
  {32'h45184fee, 32'h4378f75e, 32'hc37014a3},
  {32'hc48e3aa8, 32'hc26808dd, 32'hc2e7d6d0},
  {32'h44e69f04, 32'h43894ade, 32'hc3557ab4},
  {32'hc47d7698, 32'hc3c9201b, 32'h42613eb8},
  {32'h43c205a8, 32'h43820e54, 32'hc29f168a},
  {32'hc5114069, 32'hc389debb, 32'h422d0c46},
  {32'h44a2c7f6, 32'h428b3ba1, 32'h4349d562},
  {32'hc2e14360, 32'h427179c0, 32'hc20696ae},
  {32'h4397f868, 32'hc2cabde6, 32'h419a1a5a},
  {32'hc3da3438, 32'hc374f9e2, 32'h4229e5e7},
  {32'h43800476, 32'h4329da87, 32'h437404c1},
  {32'hc4b0e491, 32'h4384f645, 32'hc31ed0f7},
  {32'h4496171a, 32'h4320e0c3, 32'h428676ca},
  {32'hc4818399, 32'h42f83ba7, 32'hc3858d22},
  {32'h444a2331, 32'hc3238698, 32'h43233ae2},
  {32'hc4deff23, 32'h42980946, 32'hc319fab1},
  {32'h442f2c9d, 32'h430d36b6, 32'hc33de560},
  {32'hc47b8c9a, 32'h441a3381, 32'h431e38bc},
  {32'h44d82c82, 32'hc338dbef, 32'h43fde83e},
  {32'hc47ea234, 32'hc352c34f, 32'h42be517c},
  {32'h44b53df2, 32'hc36d4af1, 32'h420b0010},
  {32'hc41ea9a4, 32'hc37bdb18, 32'hc2919105},
  {32'h43fe7be0, 32'hc32324ea, 32'h43a056f5},
  {32'hc2aec8d0, 32'h421df6c0, 32'h4368dd51},
  {32'h45220426, 32'h43dfd15f, 32'hc30ff773},
  {32'hc3cdbace, 32'hc2b19fba, 32'hc3b5ae47},
  {32'h44805fe0, 32'h43b5a8a3, 32'h437ff452},
  {32'hc4db913a, 32'hc3d98cac, 32'hc3e7d97c},
  {32'h43f6ab5c, 32'h42837f2e, 32'hc2191c11},
  {32'hc4845253, 32'h4341c6ac, 32'hc31f4abe},
  {32'h445b99fa, 32'hc2dab479, 32'h4388d7a2},
  {32'hc4366ffb, 32'h42983eb2, 32'hc344cb8b},
  {32'h443118e8, 32'h42fdc91a, 32'h43a077f1},
  {32'hc50ad56f, 32'h4386d51f, 32'h3fcf678c},
  {32'h44ab91f5, 32'h42f20a73, 32'hc389e9eb},
  {32'hc405582c, 32'h4351cde5, 32'hc1a82dfd},
  {32'h43a29c8b, 32'hc137ce4c, 32'hc3f93859},
  {32'hc4c42ca4, 32'hc27187e3, 32'h43669a73},
  {32'h432e37d0, 32'hc32a52f9, 32'h430b92be},
  {32'hc3987948, 32'h422cb586, 32'h409a5570},
  {32'h450f368b, 32'h43a095ed, 32'hc33b9aa7},
  {32'hc50f9baa, 32'hc322e281, 32'h4266fb10},
  {32'h449b2b1b, 32'h4230062a, 32'h42bda408},
  {32'hc4e4f0a8, 32'hc246d689, 32'h4210b1da},
  {32'h45114b6a, 32'h4289f92a, 32'h42f53712},
  {32'hc4c251f1, 32'h430798b1, 32'hc3386128},
  {32'h44b89249, 32'hc3b1dc4f, 32'h421b695f},
  {32'hc4dc50d1, 32'h437dee88, 32'h43c409e7},
  {32'h449953f8, 32'hc2f23d28, 32'hc18c50ca},
  {32'hc482da2e, 32'h41a363cd, 32'hc39446cf},
  {32'h446675e6, 32'hc2d71743, 32'h42b7e08c},
  {32'hc4423bf4, 32'hc3ea3a8e, 32'h43591518},
  {32'h43e5fea2, 32'hc31ec8cb, 32'h4203f496},
  {32'hc45c80ea, 32'h4207bf3d, 32'hc270f9fb},
  {32'h4528ebf2, 32'hc2f85142, 32'hc3db06b3},
  {32'hc440aa82, 32'hc332eb86, 32'hc326a583},
  {32'h45021ea7, 32'hc27ea62c, 32'hc1164a02},
  {32'hc4bdf75f, 32'h4228ea68, 32'h421bd90a},
  {32'h4470165c, 32'hc3815e53, 32'hc3cd8bde},
  {32'hc446b6ac, 32'h43a54e69, 32'h436c72fb},
  {32'h42bfa170, 32'hc2fbe98d, 32'hc066f41a},
  {32'hc48bfed9, 32'hc3caef8f, 32'hc39aa1a0},
  {32'h45043d58, 32'hc3b0ce92, 32'h42e88750},
  {32'hc4ba4255, 32'hc2c56ff7, 32'h420e23f0},
  {32'h44770658, 32'hc2f5f8d0, 32'hc35c0d44},
  {32'hc34165f0, 32'h4209bb42, 32'h43000cbe},
  {32'h435b21af, 32'h41f2c587, 32'h432bf884},
  {32'hc4149450, 32'h427d4213, 32'h428f0db8},
  {32'h44aa6273, 32'h43c45744, 32'hc3606ab6},
  {32'hc4e297c8, 32'h43cd7824, 32'hc3ab82a4},
  {32'h442ef997, 32'hc3087cfc, 32'hc2b878ed},
  {32'hc4bf85f5, 32'h43959bc9, 32'hc1d88dd1},
  {32'h448261f8, 32'h42f99081, 32'h4209d27e},
  {32'hc3b6d554, 32'hc1f02bde, 32'hc1a63a98},
  {32'h439445bf, 32'h407ac112, 32'hc3ab3dbc},
  {32'hc3c47c10, 32'hc2150ff3, 32'hc31a8f2e},
  {32'h4491c152, 32'hc35e3209, 32'h429421b9},
  {32'hc4a0c835, 32'h42b47cfd, 32'h43ea317d},
  {32'h442f06dc, 32'hc3a48bb7, 32'h42d200a6},
  {32'hc50fe192, 32'hc28acb8e, 32'h42c4cc74},
  {32'h436d8193, 32'hc3506213, 32'hc0813564},
  {32'hc488bd5f, 32'h43823c84, 32'hc2dcb411},
  {32'h448597c1, 32'h42fc9e90, 32'h41515f8e},
  {32'hc2317e64, 32'h424054f4, 32'hc3274dbf},
  {32'h44ec96da, 32'hc29a2c39, 32'h43a539dc},
  {32'hc506e946, 32'h4390ec77, 32'h4389d722},
  {32'h444e734f, 32'h4386d0b2, 32'hc3a5dff0},
  {32'hc3aa4b33, 32'h42507573, 32'h422d8898},
  {32'h4515677b, 32'hc3baa2d3, 32'h421b1cd2},
  {32'hc5184178, 32'hc28edba6, 32'h43a7c3db},
  {32'h44870ec8, 32'h43b19898, 32'hc109c5fa},
  {32'hc293eae0, 32'h4398f1c8, 32'h438f62a7},
  {32'h44643d00, 32'h3d69c400, 32'hc0d6faac},
  {32'hc504649c, 32'hc3875aaf, 32'h43971eb7},
  {32'h44e43596, 32'h42910970, 32'hc386be2e},
  {32'hc4f7eca4, 32'hc3f19994, 32'hc089f67d},
  {32'h44ad7610, 32'hc2f20078, 32'hc2916a9f},
  {32'hc4f43f7c, 32'hc2b36cab, 32'h427be99a},
  {32'h44ac40f6, 32'h4350757c, 32'hc3aa8bba},
  {32'hc3965480, 32'hc2a0a3ef, 32'hc2e4ddc1},
  {32'h41f6f900, 32'hc217c0aa, 32'hc2127f62},
  {32'hc39de5ec, 32'hc3418088, 32'h43a079f6},
  {32'h44c15c50, 32'h4360a22a, 32'hc2be2722},
  {32'hc48452d8, 32'hc003b178, 32'hc1c22f04},
  {32'h443d93cc, 32'hc387d3bb, 32'h437e55e5},
  {32'hc48b4b96, 32'hc302148c, 32'h42ea4536},
  {32'h44b20ec6, 32'h43ca8df2, 32'hc3818dd8},
  {32'hc44d3cea, 32'h439e5499, 32'h43855af7},
  {32'h44c11637, 32'hc21b61ff, 32'h4278507a},
  {32'hc49cb792, 32'hc38f3d61, 32'h43b43ad7},
  {32'h43240b23, 32'h430f503c, 32'hc380a03a},
  {32'hc438ff46, 32'hc304e375, 32'h431739d5},
  {32'h44863447, 32'hc2be65d4, 32'h4186609d},
  {32'hc4d45d27, 32'hc2dd96eb, 32'hc37ac394},
  {32'h444428f6, 32'h437aee28, 32'hc2e812e4},
  {32'hc4304748, 32'h419342b2, 32'h43d6ae9b},
  {32'h438b5408, 32'h4233cb92, 32'h4262463b},
  {32'hc514e216, 32'hc2ab3170, 32'h4301b48d},
  {32'h44fa30d7, 32'h44287f78, 32'h433fa1cb},
  {32'hc488b31a, 32'hc3054ed1, 32'h43b6e9a7},
  {32'h44d1c690, 32'hc3826650, 32'hc32c9e94},
  {32'hc5042be4, 32'h43b6a9d4, 32'h43a7ec3c},
  {32'h43cd6670, 32'hc24d7154, 32'h4106fcff},
  {32'hc3e6f58e, 32'hc2c995c1, 32'h42a1f1c9},
  {32'h44ba23c3, 32'h41b1ca84, 32'hc15964ac},
  {32'hc4bcf892, 32'hc3004ffc, 32'hc1e0b7ac},
  {32'h44b516bc, 32'hc2000123, 32'hc3e75c63},
  {32'hc4dce90f, 32'hc3a49971, 32'hc3213b36},
  {32'h44f87b2a, 32'hc03f80b8, 32'h42f85b60},
  {32'hc41338c3, 32'h430607c6, 32'h4295d256},
  {32'h44e615e8, 32'hc3c4fad2, 32'hc3b06358},
  {32'hc4abc170, 32'h43b0958f, 32'hc372d7e9},
  {32'h448fcfab, 32'h438a5917, 32'h4344f892},
  {32'h44d862ea, 32'h43021894, 32'h436f008f},
  {32'hc4d08605, 32'h4389f69b, 32'h432ce372},
  {32'h4462a950, 32'hc33f1e21, 32'hc34d899f},
  {32'hc363445c, 32'h42a7cc93, 32'h43b0f9da},
  {32'h447a1474, 32'hc3adf28a, 32'hc2cb5abc},
  {32'hc4a14977, 32'h43a0865a, 32'hc130895b},
  {32'h44b9b9ec, 32'h425468ae, 32'hc2c32c22},
  {32'hc31411c1, 32'h4112f22b, 32'h4359c1c1},
  {32'h447a7d34, 32'hc32aecf9, 32'hc3805c4e},
  {32'hc50b0d29, 32'h433e6c01, 32'hc31f75c3},
  {32'h448ac344, 32'h43460a4a, 32'h429fb1d5},
  {32'hc26ff336, 32'hc436601f, 32'h438f1f58},
  {32'h44850c0e, 32'h436f4598, 32'h426566ad},
  {32'hc4e914c7, 32'hc330ae43, 32'hc1f7b6e3},
  {32'h44cc4ce0, 32'hc23aadee, 32'h431d4cdc},
  {32'hc445e290, 32'hc34a763b, 32'hbfde8969},
  {32'h43dba7c6, 32'hc381bc38, 32'hc1fbf815},
  {32'hc489b1fe, 32'h434aa4e5, 32'hc37c17f9},
  {32'h44e1f3c7, 32'h43bdbb86, 32'hc1e95e88},
  {32'hc48f8fcf, 32'h43d10a62, 32'h431ecaab},
  {32'h445eb8f7, 32'h422b3249, 32'h42a932d0},
  {32'hc4f80927, 32'h431dad83, 32'h4197be77},
  {32'h44393870, 32'h42b09a12, 32'h425553ce},
  {32'hc4eaa602, 32'h435a5acd, 32'h4374be92},
  {32'h43eea7d1, 32'hc26c1780, 32'h42325e1e},
  {32'hc4c471ea, 32'hc27208e6, 32'h43932ebb},
  {32'h44db67dd, 32'hc307728f, 32'hc1d927fd},
  {32'hc4be8300, 32'h438c1982, 32'hc2afc6f0},
  {32'h448a3ea7, 32'hc3002390, 32'hc3bb3742},
  {32'hc32a8528, 32'hc32e2765, 32'hc3213c43},
  {32'h449006ae, 32'hc232f8ca, 32'hc33afdf9},
  {32'hc4658010, 32'hc31f5ec6, 32'hc38b4612},
  {32'h433fa3a9, 32'h41a2eeb0, 32'h430767e6},
  {32'hc469ea31, 32'hc28e7b35, 32'h438ecccb},
  {32'h450f9437, 32'hc32b1475, 32'h4353fd9a},
  {32'hc3badfab, 32'hc30f4628, 32'hc3ac79de},
  {32'h442bc980, 32'hc40ff5fc, 32'hc31677e6},
  {32'hc4bed8a8, 32'h42d3c4b7, 32'h42064ec5},
  {32'h443dfd36, 32'hc35abe22, 32'hc26fe850},
  {32'hc47e657d, 32'hc074a7d4, 32'hc3dd5057},
  {32'h44ef33fc, 32'hc3215f61, 32'h411b5f76},
  {32'hc3b11e0c, 32'h427e65d8, 32'h4228a2a8},
  {32'h44655778, 32'hc33dffba, 32'h43b71187},
  {32'hc4b1ea39, 32'hc3b3fdd4, 32'h43bfe2d2},
  {32'h440b994c, 32'hc271a4e4, 32'hc24c434e},
  {32'hc50e200e, 32'h437c910f, 32'h4343558f},
  {32'h44a36938, 32'h42cab67a, 32'hc27c3186},
  {32'hc40bf8d0, 32'h4351d038, 32'h42f2d0f9},
  {32'h44b08079, 32'h428f4698, 32'h42073174},
  {32'hc4b32fb8, 32'hc31b9881, 32'h42c003ba},
  {32'h44679289, 32'h43ba4a3f, 32'hc386b71a},
  {32'hc4a1be95, 32'hc3c9267a, 32'h4249c3a2},
  {32'h44254c63, 32'hc25172e8, 32'hc35b6d0c},
  {32'hc45c86f7, 32'hc3c6eca4, 32'h42eee2b7},
  {32'h44f06ecf, 32'h41a704fe, 32'hc36fefa4},
  {32'hc4f024c5, 32'h42623e3c, 32'h42454968},
  {32'h449cca01, 32'h428da6e8, 32'hc191b751},
  {32'hc42551ea, 32'h437c5112, 32'hc401cd5e},
  {32'h4419bbe2, 32'hc2dd3c6a, 32'hc3b1b545},
  {32'hc494c0de, 32'h42b38dd9, 32'hc3123b64},
  {32'h43db1e18, 32'hc4023526, 32'hc224023f},
  {32'hc4921c56, 32'h4306bab7, 32'hc30276dd},
  {32'h442fa946, 32'h4200d2b6, 32'hc2bf9fc3},
  {32'hc4feeca6, 32'h403818b8, 32'hc2cc89c8},
  {32'h445bd540, 32'hc27b02b6, 32'h43559bfa},
  {32'hc390d4e0, 32'hc3ad4285, 32'hc22614c7},
  {32'h44fd73c2, 32'hc3185ec0, 32'hc23d672c},
  {32'hc48a2d82, 32'hc2a55d05, 32'hc1eb8911},
  {32'h44de014a, 32'h438f5603, 32'h422281e3},
  {32'hc517f722, 32'hc3a96747, 32'hc30fde56},
  {32'h443daf6b, 32'h42ae6789, 32'hc307648a},
  {32'hc4be6f90, 32'hc35f0341, 32'hc2c8f431},
  {32'h4495d850, 32'h4373bbbe, 32'h4369004d},
  {32'hc4b1c1b1, 32'h42a0a43f, 32'h440baebe},
  {32'h44f6f86c, 32'hc2694a8a, 32'h42ec2eca},
  {32'hc3f3afef, 32'hc2059075, 32'hc378cfe5},
  {32'h44e0e480, 32'h43ca99e3, 32'hc191097c},
  {32'hc4e93d3c, 32'hc37801a8, 32'hc3686655},
  {32'h45080f3e, 32'h428df51c, 32'hc2d88a26},
  {32'hc4943d3a, 32'hc2a599b3, 32'hc1fe6757},
  {32'h441d397e, 32'hc185423d, 32'hc28c75a9},
  {32'hc4c060e0, 32'h4399f2df, 32'hc26c1a9f},
  {32'h44a288ad, 32'hc317fed1, 32'h42bfb321},
  {32'hc4a7ddda, 32'h4217add3, 32'hc2f53a22},
  {32'h4404aa32, 32'h42f5b601, 32'h43546bb7},
  {32'hc48c4214, 32'h42e16654, 32'h42245cab},
  {32'h44d38d38, 32'h431f4ac9, 32'h422631f6},
  {32'hc4a3d678, 32'hc2f9ec02, 32'h4310c351},
  {32'h443e11ee, 32'hc348578c, 32'h4170215a},
  {32'hc507f0ed, 32'h42b6f70a, 32'h42c32e08},
  {32'h450df817, 32'h430e9853, 32'h436a37fe},
  {32'hc50dc164, 32'hc30575fe, 32'hc40c0fcc},
  {32'h44b3569b, 32'hc3ec34a1, 32'h4225ea9b},
  {32'hc44ac406, 32'hc2472638, 32'hc3a49a1e},
  {32'h44f3290e, 32'hc34539c0, 32'hc29673ef},
  {32'hc50c7229, 32'hc3c6b274, 32'hc32f5ae9},
  {32'h450c80a8, 32'h439feed9, 32'hc3979599},
  {32'hc4b71a69, 32'hc2b0906e, 32'h42eb55a8},
  {32'h44d804b6, 32'hc2e7703f, 32'hc2381ac6},
  {32'hc4f76059, 32'h436682ad, 32'hc37963f9},
  {32'h44b29f11, 32'h440ba0c7, 32'h43dff5f7},
  {32'hc503d9f3, 32'h43f176c2, 32'hc39defca},
  {32'h4442ec50, 32'hc3192b45, 32'h430ffc80},
  {32'hc3dd2dc6, 32'h42c8d9c5, 32'h43f09152},
  {32'h44cd79d0, 32'h42a8d95a, 32'h43859598},
  {32'hc3fe398c, 32'hc28deaf9, 32'h4185d39a},
  {32'h451b9a38, 32'h4353b4ec, 32'h3fadb120},
  {32'hc46d7354, 32'hc2f58e41, 32'h42d582bf},
  {32'h45072886, 32'hc34f4b53, 32'hc23e4ff9},
  {32'hc4ab9ab6, 32'h4287c61c, 32'h4214da22},
  {32'h4409e9d8, 32'h431f5510, 32'h4384d22c},
  {32'hc4628cb6, 32'h428e6073, 32'hc3446a23},
  {32'h44839e57, 32'hc3d61af2, 32'h428d30aa},
  {32'hc4e08d7f, 32'h429def4d, 32'h439a601c},
  {32'h44ca2a82, 32'h4340a869, 32'hc2ac3927},
  {32'hc46f8628, 32'hc1173e45, 32'h4323a852},
  {32'h44c57ff8, 32'h42118bc4, 32'h43b728cd},
  {32'hc4022803, 32'hc2314fb0, 32'h43817b74},
  {32'h450da0ae, 32'hc32ec9de, 32'hc10a830b},
  {32'hc489ec42, 32'hc39082bd, 32'h4290fa49},
  {32'h441a1032, 32'hc17ae052, 32'h4353af31},
  {32'hc3133722, 32'h435affe1, 32'h43762a17},
  {32'h45053bd8, 32'hc3ab4580, 32'h43211782},
  {32'hc4bfe7f6, 32'hc309e456, 32'h431d0a50},
  {32'h44c582ed, 32'h439b6e46, 32'h42a52ebc},
  {32'hc4f2e5cd, 32'hc360a0ea, 32'h43017614},
  {32'h4402d380, 32'h42f40557, 32'h42ae5fb3},
  {32'hc4972556, 32'hc39f4bdd, 32'h42852a77},
  {32'h4415e85e, 32'hc3128b00, 32'hc19a50b7},
  {32'hc3d2e286, 32'hc278278a, 32'h4320242a},
  {32'h449e336d, 32'h4368877d, 32'h43622aa7},
  {32'hc4fe7bab, 32'hc3c959a3, 32'h4393e3f5},
  {32'h43f92f5c, 32'hc285dad3, 32'h420e41b2},
  {32'hc3dde197, 32'h42eb1418, 32'h42cebe87},
  {32'h45209b49, 32'hc3a05628, 32'hc38e955d},
  {32'hc4ca55be, 32'hc2a3fc93, 32'hc2d97827},
  {32'h44ed8b62, 32'h432458b2, 32'h40efd382},
  {32'hc4b7bc49, 32'h42988b40, 32'h41e3211d},
  {32'h44c1c727, 32'hc33e91cd, 32'hc33983fe},
  {32'hc43c9c23, 32'h431f162c, 32'hc09308b3},
  {32'h44d26404, 32'h4341f796, 32'hc37f66e7},
  {32'hc37f6d70, 32'h43ae6b78, 32'hc2670c9e},
  {32'h44c927a2, 32'h42cc4afd, 32'hc3228fb5},
  {32'hc48f61a7, 32'h41cff8f6, 32'hc10051f4},
  {32'h4404832c, 32'hc2940a1c, 32'h436b2707},
  {32'hc48ccf32, 32'hc36d00ce, 32'hc2c4c86f},
  {32'h441b1ed8, 32'h4344fb08, 32'h42089e75},
  {32'hc42e235e, 32'h4357753f, 32'h4368ebcb},
  {32'h441ebd79, 32'hc38af9cb, 32'h42dbce57},
  {32'hc4290782, 32'hc34088fc, 32'hc376d437},
  {32'h4515559e, 32'hc30a261f, 32'hc24d043b},
  {32'hc503a6a1, 32'h43dfd3b7, 32'h43660c1b},
  {32'h4513da69, 32'hc3bea168, 32'hc2e9a0bd},
  {32'hc5027aca, 32'hc30299fc, 32'hc216cffb},
  {32'h44d114f3, 32'h43385554, 32'hc39d0f91},
  {32'hc4a38804, 32'h43077cb7, 32'h439ac8b0},
  {32'h440b22d0, 32'hc2ec7ebc, 32'hc08962c6},
  {32'hc37c9c20, 32'hc3f04bb2, 32'h42b3bfcf},
  {32'h447c9223, 32'h435a221f, 32'hc36918fb},
  {32'hc39cbf06, 32'h41d17ade, 32'h431b77d3},
  {32'h4456c1f2, 32'hc3b21658, 32'h430baf42},
  {32'hc461c4af, 32'hc286fc82, 32'h4236c65d},
  {32'h43094de4, 32'hc25d6816, 32'h43cd74e0},
  {32'hc5022f68, 32'h41424f77, 32'hc2918759},
  {32'h43925d2f, 32'hc2770925, 32'hc25b4b38},
  {32'hc4f55599, 32'hc3a81649, 32'hc31c3564},
  {32'h44246c4a, 32'h44078efc, 32'hc2dba31c},
  {32'hc3b29b9d, 32'hc344f168, 32'hc0e3aefc},
  {32'h4367b770, 32'h42f57178, 32'hc294ce21},
  {32'hc4dc0e3a, 32'hc285d93d, 32'hc2b66283},
  {32'h44f55dfc, 32'h429c2938, 32'hc320d186},
  {32'hc3f0ec04, 32'hc38d3648, 32'h43d04c50},
  {32'h44b9cd3e, 32'h407bf356, 32'h4066766e},
  {32'hc402d438, 32'hc39057bc, 32'h42d193d1},
  {32'h44e36d2d, 32'h43a2c3ab, 32'hc293ecab},
  {32'hc3fa5688, 32'h41cc6dbc, 32'h42bade3e},
  {32'h443cb118, 32'hc2434538, 32'h43121945},
  {32'hc4a70148, 32'h41b747b6, 32'h43586e84},
  {32'h44e24b56, 32'hc21a1d07, 32'h40b110f0},
  {32'hc4a5f469, 32'hc235ae06, 32'h42b0852d},
  {32'h4454741b, 32'hc1e196b9, 32'hc2ab636b},
  {32'hc31f718b, 32'hc295745d, 32'hc3e86587},
  {32'h44f7b72a, 32'h4134e506, 32'h4400e23d},
  {32'hc3d57fc0, 32'hc32decae, 32'hc2e7d69c},
  {32'h43efcb9f, 32'hc34c4814, 32'h434fb093},
  {32'hc4f67d95, 32'hc1dc1582, 32'h41a1d541},
  {32'h4500b902, 32'h43b0caa3, 32'h42909098},
  {32'hc4c0f11a, 32'h42aeb9c1, 32'h43093ece},
  {32'h44b82d6a, 32'hc364c7e2, 32'hc36836fd},
  {32'hc496e2b0, 32'hc3a794d4, 32'h43626ad3},
  {32'hc112d510, 32'hc28ea4b8, 32'h43fa389e},
  {32'hc50a9849, 32'hc298f89a, 32'hc226452c},
  {32'h44b41326, 32'h4176ff4a, 32'hc35a35c2},
  {32'hc4893c5c, 32'hc17f2c42, 32'h426ae0bf},
  {32'h44586330, 32'hc31a1740, 32'hc27956dc},
  {32'hc460af5f, 32'hc30efbbb, 32'h421b30ef},
  {32'h446aff68, 32'hc3795d57, 32'hc279bb05},
  {32'hc3d69940, 32'h4208d599, 32'hc2608439},
  {32'h442dab34, 32'hc3a979d3, 32'hc322f925},
  {32'hc4e945ff, 32'hc31f33e0, 32'h43a99234},
  {32'h445b9f24, 32'h43e82aa2, 32'hc24ecdf6},
  {32'hc486ef8b, 32'hc3808c11, 32'h43658cbf},
  {32'h44385930, 32'h42aa6dae, 32'hc3129f79},
  {32'hc4714454, 32'h42cdadf2, 32'h4318ce99},
  {32'h4407ee84, 32'h4348bad8, 32'h42db978c},
  {32'hc412fa51, 32'h4404d09b, 32'hc3817ac0},
  {32'h44e1e634, 32'hc213ab8c, 32'hc20b05f3},
  {32'hc44b104f, 32'h41c4ac7f, 32'hc3942c7c},
  {32'h449d5b54, 32'hc3a0f5bc, 32'h43ce034e},
  {32'hc4a364e4, 32'hc3c5e8ac, 32'h43086e4f},
  {32'h44a27b93, 32'hc2e3f2f2, 32'hc339ad10},
  {32'hc438aa46, 32'h435cd5fa, 32'h439f3a2b},
  {32'h44910fca, 32'h43238e82, 32'hc28a2a3a},
  {32'hc3bdb120, 32'h442d619d, 32'hc1fd3a38},
  {32'h440a8fc0, 32'hc1211a5f, 32'hc29ddae9},
  {32'hc4962421, 32'h43c0251e, 32'h4302aeb9},
  {32'h43946bd0, 32'hc3717eec, 32'hc2c27822},
  {32'hc4138611, 32'hc2248a80, 32'hc2e268c4},
  {32'h445e187a, 32'hc1b191ce, 32'h422531cb},
  {32'hc3964538, 32'hc1811600, 32'hc29bb72a},
  {32'h45031ef8, 32'hc3241aaa, 32'hc3b406f6},
  {32'hc4db5504, 32'h4326a59b, 32'h4333af5a},
  {32'h431b9cea, 32'h433058aa, 32'h4330eb68},
  {32'hc4b7e86f, 32'h40a76bd4, 32'hc223ba30},
  {32'h4425cd32, 32'h42ea3b6f, 32'hc352f636},
  {32'hc485daed, 32'h43849c59, 32'hc3fb49ba},
  {32'h44355f93, 32'hc39464e9, 32'h41a63404},
  {32'hc4ac7fc3, 32'hc2c863f9, 32'h4238b115},
  {32'h44635c84, 32'hc3bd49ac, 32'h41ae427c},
  {32'hc3f3a954, 32'h435cae58, 32'hc328f49e},
  {32'h4406df76, 32'h430d07e1, 32'h43bf0e91},
  {32'hc507d4ac, 32'h415affca, 32'h41cb0de3},
  {32'h43784c5c, 32'hc2196fd4, 32'h4308249a},
  {32'hc4db1564, 32'h41df8cae, 32'h42c02798},
  {32'h44b2ae9c, 32'h432fa773, 32'hc3368598},
  {32'hc3ebf6a0, 32'h436d9289, 32'hc351c866},
  {32'h44dbae67, 32'h4122afd8, 32'hc3450b40},
  {32'hc48babb1, 32'hc348aced, 32'h422fcf53},
  {32'h44206071, 32'hc35c1745, 32'hc35d552a},
  {32'hc4a010b8, 32'h421acf17, 32'hc14e53a5},
  {32'h4492a8b8, 32'h429e6641, 32'hc408f495},
  {32'hc448a5f9, 32'h42be9fb6, 32'hc2c575d0},
  {32'h447394e7, 32'hc2dd90f1, 32'h4240f8a0},
  {32'hc491eb9b, 32'hc1efb8c4, 32'h43b508b4},
  {32'h4483aff5, 32'h434a3a08, 32'h42f15ee9},
  {32'hc50a4a72, 32'h42049cc9, 32'h42f915fd},
  {32'h44b2db57, 32'hc360db17, 32'h4235ca51},
  {32'h4382ab1d, 32'h43a47278, 32'h42ba928e},
  {32'h44a4b13c, 32'h43cc5af5, 32'h43893109},
  {32'hc5038ef3, 32'hc39aeb6d, 32'hc366d66e},
  {32'h4481d413, 32'hc0dc58f8, 32'h43c67778},
  {32'hc505756f, 32'h42eff098, 32'hc3274edb},
  {32'h44f0b2a3, 32'h41a0e74e, 32'h436bc26b},
  {32'hc4a8cc91, 32'h42b1a3a6, 32'h42c5d3cd},
  {32'h44be983c, 32'hc2b8116c, 32'h417f13e6},
  {32'hc437e2a2, 32'h422b80a4, 32'hc38cdf80},
  {32'h44133e80, 32'hc3b26e07, 32'h40d1735f},
  {32'hc4325758, 32'h42650c66, 32'h43400e49},
  {32'h44b4c216, 32'hc2d4f2ee, 32'h43d04dd6},
  {32'h433888f0, 32'hc3a28998, 32'hc25abcce},
  {32'hc39b0c26, 32'h42fece65, 32'hc346e63e},
  {32'h427e388c, 32'h437f2aca, 32'h4218b1e6},
  {32'h44f6b406, 32'h4396443c, 32'h433973a8},
  {32'hc4f431a2, 32'hc2892d3b, 32'h42c30030},
  {32'h4503b325, 32'hc261e130, 32'hc190b2c7},
  {32'hc4c2b535, 32'hc22fa157, 32'h434492e7},
  {32'h44c392be, 32'h42f6036c, 32'hc3700b72},
  {32'hc46ecd50, 32'h4355cccc, 32'h42fa9c8e},
  {32'h44661133, 32'h43e27084, 32'h43678fba},
  {32'hc4f97a2c, 32'hc35ecc8e, 32'hc271b0c8},
  {32'h441c1180, 32'h42e96604, 32'h43b05e60},
  {32'hc4c7845e, 32'h417381ff, 32'h43603bb0},
  {32'h45087649, 32'hc38fcd4b, 32'hc3512e79},
  {32'hc3a7cd34, 32'h4321ebb7, 32'h4216de95},
  {32'h449392b4, 32'hc30c9cb0, 32'hc3968ac5},
  {32'hc513aaed, 32'h43b58353, 32'h416f6926},
  {32'h43dcf795, 32'hc33d4833, 32'hc3c0205c},
  {32'hc49b17e3, 32'hc298d784, 32'h42ee29a8},
  {32'h44eb12d1, 32'hc3a0a095, 32'hc346066a},
  {32'hc4bd3860, 32'h428b7e0b, 32'h43485886},
  {32'h44cac08d, 32'h442081b2, 32'h431f9c24},
  {32'hc45aaed9, 32'hbecf0460, 32'hc39d9a9b},
  {32'h446af038, 32'hc26a5b57, 32'hc2bcb7c2},
  {32'hc4ce7730, 32'hc28bff5c, 32'h41fc5bc6},
  {32'h44f6a78e, 32'hc09c5543, 32'hc28c96c9},
  {32'hc4bb5485, 32'hc106b84e, 32'h42cddf73},
  {32'h4500673f, 32'hc27b8705, 32'h4321216f},
  {32'hc4decfa8, 32'hc340bf84, 32'hc31eb4ca},
  {32'h44eea74b, 32'hc3492a3f, 32'hc337c243},
  {32'hc4c58a74, 32'h430b92b7, 32'hc236a783},
  {32'h45004ac7, 32'hc3249466, 32'hc343c8a8},
  {32'hc4f6b026, 32'hc3099f56, 32'h40864538},
  {32'h44eaf523, 32'hc3264ec4, 32'h43ac27c0},
  {32'hc48f1a5f, 32'hc3b49ec3, 32'h42b19823},
  {32'h450288ef, 32'h42ce3fc8, 32'hc38c72a4},
  {32'hc426756e, 32'hc2e3448c, 32'hc2a1c09f},
  {32'h44ea479c, 32'hc3863565, 32'h430339a3},
  {32'hc41307b6, 32'h43857a87, 32'h429bb1d9},
  {32'h44c86448, 32'h43460311, 32'h43cc6e4d},
  {32'h42fefba0, 32'hc363b23f, 32'hc36d478f},
  {32'h4486665b, 32'h4304ea1c, 32'hc34d82fa},
  {32'hc51117f0, 32'h43975b90, 32'h430b89d0},
  {32'h43a66628, 32'h410c55e0, 32'hc317033f},
  {32'hc4ed90c3, 32'h43c8b601, 32'h43321278},
  {32'h4485315e, 32'h4281a128, 32'hc30f7e90},
  {32'hc41b9ab7, 32'hc1ce4b01, 32'hc309f8f1},
  {32'h44707e70, 32'hc1d019e6, 32'hc3fa603a},
  {32'hc50d3c78, 32'h4336038b, 32'hc2231b3c},
  {32'h448d18c5, 32'hc29cee93, 32'h43c586b0},
  {32'hc50c7a51, 32'hc3e40ce3, 32'h4203e5be},
  {32'h44117ddc, 32'hc3ffe098, 32'hc3008ee2},
  {32'hc4b64cfa, 32'h43d69b1b, 32'hc2d13c98},
  {32'h450d39a9, 32'h435e080b, 32'hc2f51f1e},
  {32'hc4b3bd00, 32'hc1fe169c, 32'hc1d4c240},
  {32'h4449b933, 32'h43201776, 32'hc394f07a},
  {32'hc3647cd0, 32'hc332ce3e, 32'h42fcfe8a},
  {32'h443c4592, 32'h4323a298, 32'hc0d915d3},
  {32'h4250c180, 32'hc2af665c, 32'h3e3e3550},
  {32'h44949180, 32'hc2a4497f, 32'h4327bbf3},
  {32'hc49db993, 32'hc32305d8, 32'hc393f948},
  {32'h444bef7f, 32'h42f8d66d, 32'h43902f13},
  {32'hc486fa95, 32'h436c02bc, 32'hc2a05a53},
  {32'h44e83382, 32'h436ee167, 32'hc259d9a2},
  {32'hc4ec85f5, 32'h415660a3, 32'hc29a48d4},
  {32'h44e3e61e, 32'h43b5ce2e, 32'h434315f8},
  {32'hc5035e24, 32'hc2b84a3a, 32'h42f65b2f},
  {32'hc1cab920, 32'hc34925dc, 32'h4341a399},
  {32'hc45c9e4a, 32'h440327b0, 32'h439e9e2f},
  {32'h44d8f731, 32'hc26c2bb5, 32'hc24b328d},
  {32'hc4b94087, 32'h43b0262e, 32'h439a461b},
  {32'h447c0bd3, 32'hc32593ce, 32'hc2d78e36},
  {32'hc2e28fa0, 32'hc1be275c, 32'hc2827383},
  {32'h450db6f5, 32'hc01fa6fe, 32'hc255654d},
  {32'hc39634da, 32'h43202eec, 32'hc360fe63},
  {32'h44fd4729, 32'h422cc3ef, 32'h43782e98},
  {32'hc40b1765, 32'hc35abc01, 32'hc3adcf82},
  {32'h43a09f0c, 32'h433265d1, 32'h42b5f4c5},
  {32'hc4cc3716, 32'hc3abe4bd, 32'h42faed19},
  {32'h43d0e9fc, 32'hc2aa7946, 32'hc38b7bdb},
  {32'h4391f4cc, 32'h426b291c, 32'h43344ed6},
  {32'h4442cd6c, 32'hc2dfddc3, 32'hc3ab75c7},
  {32'hc4482f00, 32'h42b21e7e, 32'hbfb71d40},
  {32'h450df3d4, 32'hc2face07, 32'h43ad12dd},
  {32'hc4c9a812, 32'h433f8c92, 32'h432fc8f8},
  {32'h44eb7c71, 32'h42e439cf, 32'hc2180b90},
  {32'hc4c025a6, 32'h431c782f, 32'hc0cd6968},
  {32'h439b76e8, 32'h4176d3d4, 32'h43a8bd5d},
  {32'hc3e65a1e, 32'h433b95a2, 32'h442576b5},
  {32'hc1d84860, 32'hc304164f, 32'hc29f0f72},
  {32'hc40d862c, 32'hc1d64e84, 32'hc2f7a995},
  {32'h44cf1f68, 32'h41a2e402, 32'h437eecfd},
  {32'hc47b8f0e, 32'hc10633b5, 32'hc286feb9},
  {32'h44a8a7d4, 32'h43679bbb, 32'hc3065cf1},
  {32'hc4f37024, 32'hc31d2bee, 32'hc3b4c44d},
  {32'h4498e815, 32'hc40fc2f5, 32'hc3086bf0},
  {32'hc502c79f, 32'h43d610ba, 32'hc31ec2ab},
  {32'h44a65c9c, 32'h43002cae, 32'h43088487},
  {32'hc3e26698, 32'h42bfb160, 32'h42960bf4},
  {32'h4512bf72, 32'hc28aa09f, 32'hc35bd15b},
  {32'hc3ac70f4, 32'hc34250ad, 32'h431097eb},
  {32'h44a1b17d, 32'hc2c95791, 32'h3f3cbd5a},
  {32'hc48bceae, 32'h4359a7fc, 32'hc314f9ff},
  {32'h43bc9bcc, 32'h42a8e91d, 32'h41b54f55},
  {32'hc4990637, 32'h4319fb8c, 32'hc321b508},
  {32'h45068e3e, 32'hc2ae4d17, 32'hc3805a3d},
  {32'hc43c35d3, 32'h434a73e5, 32'h42f92420},
  {32'h44ce807a, 32'hc23e5f32, 32'h43a0ae57},
  {32'hc3fc0580, 32'h401f9f18, 32'hc30384a3},
  {32'h450ef11d, 32'h4293547c, 32'h430b1b46},
  {32'hc4fa3b07, 32'hc3a42eed, 32'h43e76e43},
  {32'h45481d77, 32'h4394588a, 32'hc343a004},
  {32'hc4be8fd0, 32'hc3ff4e8e, 32'hc32b9b89},
  {32'h44eeb856, 32'hc2ae7c80, 32'hc32906f4},
  {32'hc410b610, 32'hc329ff7d, 32'hc3901186},
  {32'h448e46e5, 32'hc39e37a5, 32'h434bc4d1},
  {32'hc402d63c, 32'h40543438, 32'hc2cb275d},
  {32'h45092b3c, 32'hc36ed49f, 32'h42109f6a},
  {32'hc499766c, 32'hc2bdfe88, 32'h42d1ddc6},
  {32'h43d8b390, 32'h407a602a, 32'hc2efdc2e},
  {32'hc4a3e587, 32'h415ada0d, 32'h436e3c9e},
  {32'h442d38e6, 32'hc2829044, 32'hc28569c2},
  {32'hc4248fca, 32'h4376aba2, 32'hc3838cc8},
  {32'h4461ea64, 32'hc3379349, 32'hc3b4f175},
  {32'hc46d5674, 32'h42978c5d, 32'hc2d0e49a},
  {32'h451ac5b2, 32'hc29a7573, 32'h42d4f909},
  {32'hc45ddf5a, 32'h440374a0, 32'hc2db8a80},
  {32'h4530fdf8, 32'h421c5ac4, 32'h42b6f264},
  {32'hc36934b8, 32'hc2c39008, 32'hc3b4d10c},
  {32'h4456b670, 32'hc33c5578, 32'hc19426a2},
  {32'hc32b831d, 32'h43ae5457, 32'hc3c0590b},
  {32'h4506187e, 32'h431586ed, 32'h42d0aa8f},
  {32'hc4b320f2, 32'hc21c0c86, 32'hc385bcc3},
  {32'h4510e633, 32'h436ede58, 32'h42fe7aa5},
  {32'hc4e01a2c, 32'hc2e8d389, 32'h430cf169},
  {32'h43daddd8, 32'h42770b22, 32'h42f26ebe},
  {32'hc2aaf75e, 32'h421be8ee, 32'hc34a1865},
  {32'h42eba970, 32'h4282b587, 32'h4225c5fb},
  {32'hc4c79b7f, 32'h43132707, 32'h432ce2aa},
  {32'h44e5b339, 32'hc2d55a8a, 32'hc17ba9cd},
  {32'hc4b5f119, 32'hc10504e6, 32'hc3f0d013},
  {32'h44ffd6c5, 32'h432f7e3a, 32'hc2101c32},
  {32'hc507e86e, 32'h43d492b5, 32'hc3eef7a0},
  {32'h44b30af2, 32'h42be03ff, 32'h425b0a6d},
  {32'hc466ae40, 32'hc2a1a4e6, 32'hc1db366d},
  {32'h446410e2, 32'h430e931f, 32'h438e0aa6},
  {32'hc489bee2, 32'h43376dd2, 32'hc3427a6c},
  {32'h449df601, 32'hc181a0be, 32'h43a28c20},
  {32'hc4f29498, 32'hc38a6427, 32'hc370b48e},
  {32'h44ec3656, 32'hc30ff0f6, 32'hc282b73c},
  {32'hc4e1a427, 32'h412cf72f, 32'h41d5e019},
  {32'h429607ec, 32'h4325151b, 32'h433d1b16},
  {32'hc39bc114, 32'hc25a1f18, 32'hc2bfe3db},
  {32'h439530f2, 32'h43a0fa00, 32'h4317e154},
  {32'hc48faffe, 32'h4322ad0f, 32'h42e76c5c},
  {32'h4430c440, 32'h42c45c68, 32'h4396eead},
  {32'hc2eecfd0, 32'h43840897, 32'hc30afe24},
  {32'h41fe13a0, 32'hc2e93944, 32'h43991507},
  {32'hc40519eb, 32'hc321fca4, 32'hc29abd8b},
  {32'h43c6e3f0, 32'h437c661b, 32'h43040996},
  {32'hc4b7b33e, 32'h440d9b92, 32'hc3dac22d},
  {32'h4383d5ff, 32'hc23c29cc, 32'h4319cab1},
  {32'hc42197ba, 32'h4349f58b, 32'hc392ab99},
  {32'h449c1850, 32'hc1914126, 32'hc20d8252},
  {32'hc40e3547, 32'hc3d63408, 32'h4319fd7c},
  {32'h424caa30, 32'h418d03d0, 32'h43858b2f},
  {32'hc3a91718, 32'h4320bc9c, 32'hc356daac},
  {32'h45000ffd, 32'h43a94933, 32'h4263bd96},
  {32'hc4d66c94, 32'h42964300, 32'hc2c49e3f},
  {32'h448bc9f8, 32'hc2e10089, 32'hc303e78a},
  {32'h431461c7, 32'hc409fa93, 32'hc3602af1},
  {32'h451c8f0e, 32'h438a5104, 32'hc2764e40},
  {32'hc49900b5, 32'hc2feaede, 32'hc3d86a26},
  {32'hc3c58fc4, 32'hc309f6f3, 32'h42a3552d},
  {32'h441e82be, 32'h433b131f, 32'hc1fc56ea},
  {32'hc4e8c08e, 32'h4415af1f, 32'h4326c902},
  {32'h44e2ba24, 32'hc3002236, 32'h41d227a5},
  {32'hc4972362, 32'hc30992a2, 32'hc320d2c6},
  {32'h44b4313d, 32'h4347c9fa, 32'hc2f6cccf},
  {32'hc48223fc, 32'hc267eda1, 32'hc398712a},
  {32'h44577a9a, 32'h428e5403, 32'h432003f1},
  {32'hc4935eca, 32'hc215027c, 32'hc2f2ed4f},
  {32'h44c68eb9, 32'h430fac64, 32'h427d634c},
  {32'hc3703484, 32'h431cadae, 32'hc341035c},
  {32'h43f06dc4, 32'hc3bd2fce, 32'hc25eb25c},
  {32'hc4e64449, 32'hc2fe6efc, 32'hc3192227},
  {32'h447ff4fb, 32'h43b01db8, 32'h434a3fac},
  {32'hc4f3d62a, 32'h428f08d6, 32'hc310c01e},
  {32'h44203627, 32'h4350ca7a, 32'hc433abbf},
  {32'hc4ac3159, 32'hc323bbbb, 32'hc2ca5baa},
  {32'h44697c37, 32'h41fa58df, 32'h425a0109},
  {32'h42f48018, 32'h431575c6, 32'h43374194},
  {32'h43190544, 32'h4377120a, 32'h432471e8},
  {32'hc49c7133, 32'h4396274c, 32'h434fe059},
  {32'h44604330, 32'h42ecd1e9, 32'h419867f2},
  {32'hc465d78c, 32'h432ecb0b, 32'hc294e966},
  {32'h450fd49d, 32'h4326833b, 32'h433c31ee},
  {32'hc48d9fce, 32'h439a61d3, 32'hc3f16724},
  {32'h44c5747a, 32'h415de6c1, 32'h433133e9},
  {32'hc46cdb0e, 32'hc0409fae, 32'hc380a2d6},
  {32'h44947fb3, 32'hc28cb0d3, 32'h4108cf77},
  {32'h426ac900, 32'h4368c9a6, 32'hc3117c47},
  {32'h45114398, 32'h43de9bb2, 32'h42de1109},
  {32'hc46f6a18, 32'h431bd91b, 32'hc3a4c945},
  {32'h4502b843, 32'hc2dab19f, 32'h43d955a6},
  {32'hc403f24a, 32'h43003ed3, 32'hc339d8e8},
  {32'h44ab7d08, 32'h43140bfe, 32'h4361300f},
  {32'hc3c54b10, 32'h436663a9, 32'hc327c09d},
  {32'h442cb6da, 32'hc207b393, 32'hc3a04b33},
  {32'hc48503b0, 32'hc34ce1f1, 32'hc41858c5},
  {32'h44989516, 32'h438bc8fe, 32'h419266e8},
  {32'hc3cfb2f0, 32'h42b317a1, 32'h4389edb3},
  {32'h43e6c3a8, 32'h41ed805b, 32'h4363bdd0},
  {32'hc413380d, 32'hc25b32de, 32'hc183e47a},
  {32'h43b1e5c4, 32'h424b7cf9, 32'hc38630c9},
  {32'hc50fd81d, 32'hc31119c1, 32'hc0fecc23},
  {32'h451602a3, 32'h4325c0bd, 32'h43338970},
  {32'hc4e39a3a, 32'hc3780343, 32'h432eaf9e},
  {32'h44c43480, 32'hc28379df, 32'hc1d11344},
  {32'hc386faf5, 32'hc1c26c7a, 32'hc20a620d},
  {32'h451bb89b, 32'h437c1c87, 32'h43284fe5},
  {32'hc4674f7c, 32'h42aec36c, 32'h42b56408},
  {32'h44963dfb, 32'h43ce5b7a, 32'hc2b1dd19},
  {32'hc4e81498, 32'h433ba9c1, 32'hc30c1491},
  {32'h4504ab5b, 32'h42bd382e, 32'h4358ee59},
  {32'hc46f79e8, 32'h4322e0c7, 32'hc3ced086},
  {32'h426db570, 32'h43a96666, 32'h424d4df1},
  {32'hc4dfd46a, 32'h43252f84, 32'hc33cad2b},
  {32'h43752e04, 32'h41a6f641, 32'h41ac317e},
  {32'h418fb3c0, 32'h4343b8ef, 32'hc3b77688},
  {32'h43cc7f5c, 32'hc36f6d5f, 32'h438feec1},
  {32'hc4c10862, 32'h43257e0e, 32'hc300b724},
  {32'h4430598c, 32'h433625a6, 32'h426d637c},
  {32'hc487fd5d, 32'h435c2be0, 32'hc381e6ba},
  {32'h4465544a, 32'hc2a71f51, 32'h42bd7fbd},
  {32'hc3cbcdc0, 32'h401d412d, 32'hc3289b54},
  {32'h42281630, 32'hc38ce97f, 32'hc2792441},
  {32'hc45c58eb, 32'h41bc8b80, 32'h4419a2e0},
  {32'hc3750864, 32'h4386b225, 32'h43f36561},
  {32'hc2596bc0, 32'hc2274f8b, 32'h43174ad4},
  {32'h450e8b48, 32'h431d66c4, 32'hc3100734},
  {32'h432b9bbf, 32'h439187c8, 32'h42c6e434},
  {32'h43bd6ce8, 32'hc34c00fc, 32'hc3bdaad4},
  {32'h4333793d, 32'h4353232f, 32'hc2bc67e0},
  {32'h44c117df, 32'hc24f42a1, 32'hc286242f},
  {32'hc313a5a0, 32'h3f00f026, 32'h43bda3d0},
  {32'h44f1060f, 32'h43948ceb, 32'hc31ae2a4},
  {32'hc419ff74, 32'hc2fefec6, 32'h435ad9b6},
  {32'h3f0f2800, 32'h435525d3, 32'hc340721c},
  {32'hc4f6d047, 32'hc3a1fbaa, 32'hc226cf63},
  {32'hc19708c0, 32'h43e265e5, 32'h438d1c30},
  {32'hc482f25f, 32'h435c5d70, 32'h425ec22a},
  {32'h44e612f6, 32'hc337af7b, 32'h444420ef},
  {32'hc4d8c6c8, 32'hc3233880, 32'h435953cc},
  {32'h44ba3c76, 32'hbf1e5da8, 32'h42e337cb},
  {32'hc3bb1ba4, 32'h431922e4, 32'hc31c0005},
  {32'h44ea1d03, 32'h428d1d01, 32'h42cf6afa},
  {32'hc3ec5200, 32'hc296dda5, 32'hc3615d8a},
  {32'h441e1547, 32'h4318f0e7, 32'h429a4aad},
  {32'hc4c01d42, 32'hc338e4d1, 32'h4144a8ff},
  {32'h433a76c0, 32'h43d1a0f4, 32'hc3228f44},
  {32'hc371a291, 32'h435a1163, 32'h431b93f3},
  {32'h42f1889f, 32'h436c8985, 32'h42a5452f},
  {32'hc3b2ed70, 32'hc2823785, 32'h42aab174},
  {32'h44b031e8, 32'hc1aeefcf, 32'h438797b2},
  {32'hc4a65856, 32'hc2a71934, 32'h42fc0471},
  {32'h44e8eb55, 32'hc326936f, 32'h442f918d},
  {32'hc51ccad8, 32'h4390084b, 32'hc1a2c192},
  {32'h42f1bca0, 32'hc24d288b, 32'hc20819ce},
  {32'hc2a30b70, 32'hc2fcb370, 32'h4403dd47},
  {32'h451557ba, 32'h41c0abb7, 32'hc379ffaf},
  {32'hc49e3736, 32'h41d16b53, 32'h42a23cda},
  {32'h44861bea, 32'hc2f262e2, 32'hc2d3417c},
  {32'hc4e72416, 32'h41a9d0e6, 32'hc1c56182},
  {32'h44fdb450, 32'h43805f90, 32'hc3134b9e},
  {32'hc4f52b03, 32'hc13125cb, 32'hc29441bc},
  {32'h448b5961, 32'hc34aae90, 32'h42d54625},
  {32'hc416b40a, 32'h43e80a38, 32'h43b54e3c},
  {32'h44f191eb, 32'h40ee43cc, 32'h42743a42},
  {32'hc42ad63a, 32'h42330c14, 32'hc2750a86},
  {32'h45006480, 32'hc31cd59d, 32'h43083990},
  {32'hc4fa0db8, 32'h429b165c, 32'h4279fde6},
  {32'h45007ef6, 32'h42c8b3ca, 32'h440e3b28},
  {32'hc3a0b268, 32'h425dfc6f, 32'h430139cf},
  {32'h44cda564, 32'h42238e7f, 32'hc2e4c5c2},
  {32'hc47fda32, 32'h4403d2ca, 32'h431d1ffd},
  {32'h41c66570, 32'h43ee1628, 32'h42b4396c},
  {32'hc47a4eb7, 32'h42aac3a1, 32'h437e6a6d},
  {32'hc30b08fc, 32'hc3253904, 32'h422ca61f},
  {32'hc4b66a7d, 32'hc38c85a9, 32'h42f62dbc},
  {32'h43f4103c, 32'hc1c24680, 32'hc3368f0b},
  {32'hc3f0cb94, 32'h41c6a180, 32'h4400bd7c},
  {32'h44918deb, 32'h43662a63, 32'h433261c6},
  {32'h4313b530, 32'hc23182f6, 32'h4308fd6a},
  {32'hc2f07780, 32'hc27a99d6, 32'h43a90d61},
  {32'hc39eef7c, 32'hc320566a, 32'h42b0654d},
  {32'h4445414b, 32'hc30998de, 32'h41d9f762},
  {32'hc4cc5525, 32'hc2fcfed5, 32'h437587c7},
  {32'h4501b9a7, 32'hc2998fe0, 32'hc2c1bb7f},
  {32'hc4f1ce26, 32'h43aa9ef7, 32'hc333a730},
  {32'h443c35ba, 32'hc35bb984, 32'hc33c0514},
  {32'hc509f0be, 32'h42cbb0e7, 32'hc3b04c13},
  {32'h44bf9199, 32'h43c1df42, 32'hc2a9739c},
  {32'hc4b27974, 32'hc393d8de, 32'h437cde35},
  {32'h42a8bf8a, 32'h43bbff15, 32'h40374cc8},
  {32'hc37e1e88, 32'hc2c20d75, 32'h4136bcbb},
  {32'h44aeff3b, 32'hc114a531, 32'hc35b55c9},
  {32'h42a498a8, 32'hc07fb3d4, 32'h42f3c4f6},
  {32'h449b001b, 32'h428e78dd, 32'hc34908be},
  {32'hc4c336c3, 32'hc3d7b200, 32'hc3ae3e9e},
  {32'h448f76a7, 32'h43c32393, 32'hc39eea92},
  {32'hc4004768, 32'h42c00e8f, 32'hc29dee30},
  {32'h450a583f, 32'h4355778f, 32'h42c83f14},
  {32'hc487c83e, 32'h43334ed9, 32'h4268e7af},
  {32'h44a5afef, 32'hc2a1e536, 32'hc2eb41f0},
  {32'hc4c02034, 32'h42cebc0f, 32'h435181ce},
  {32'h44d90610, 32'hc233763a, 32'hc39c54af},
  {32'hc4aeb456, 32'hc23e2f68, 32'h42f0be95},
  {32'h44f709b4, 32'hc15edcf6, 32'hc2b496e4},
  {32'hc4927464, 32'h441ea2ef, 32'h435c31cb},
  {32'h448002e0, 32'h424bc85a, 32'h43cac991},
  {32'hc4cc0500, 32'h430f7148, 32'h43eb5ada},
  {32'h44dda5ce, 32'h438b3782, 32'hc335a929},
  {32'h411a224c, 32'hc41a4688, 32'hc1c64970},
  {32'h44e911c0, 32'h43a827f6, 32'hc252ca1f},
  {32'hc5022bf4, 32'hc18cef34, 32'h427343f6},
  {32'h43759540, 32'h42b90529, 32'h43953e29},
  {32'hc4e75fc4, 32'hc328d57e, 32'hc3240c9c},
  {32'h44d0ec9a, 32'hc2fc799e, 32'hc3348710},
  {32'hc50161d9, 32'hc29acecd, 32'h436a9c40},
  {32'h44a03170, 32'hc2e5c8c7, 32'hc321ca60},
  {32'hc50740f8, 32'hc1402df4, 32'hc25c9196},
  {32'h44f21d96, 32'hc40bf826, 32'hc2e486c1},
  {32'hc324026a, 32'h41ff80ce, 32'h4347c4ec},
  {32'h441ec8e4, 32'h43706a91, 32'h43828afc},
  {32'hc48656c7, 32'hc21025bf, 32'hc24cbc87},
  {32'h44c99dce, 32'h433de19b, 32'hc3357c79},
  {32'hc4f7a8c0, 32'hc22fe567, 32'hc2fd941b},
  {32'h44e824a2, 32'h4385bf2e, 32'h42f75f34},
  {32'hc3ddf762, 32'hc255209c, 32'hc3dfb481},
  {32'h43952540, 32'h43851c46, 32'h43f8437a},
  {32'hc4965070, 32'hc2183ec5, 32'hc342c368},
  {32'h451b9d84, 32'hc3111106, 32'h437a3345},
  {32'hc30971cc, 32'h434cf204, 32'hc2368394},
  {32'h44c28583, 32'hc3705305, 32'hc3af4f1a},
  {32'hc4987809, 32'h43b0051a, 32'hc1e2cead},
  {32'h44f62be0, 32'hc300f816, 32'h430efb00},
  {32'hc486b3fd, 32'hc2897a26, 32'hc3143f37},
  {32'h441010da, 32'hc43b1536, 32'h430160e5},
  {32'hc402b7a7, 32'hc2ece4c0, 32'hc315ddc3},
  {32'h4420e650, 32'hc3e69d49, 32'hc2e0f269},
  {32'hc4917226, 32'hc3cf0144, 32'hc380fbc9},
  {32'h44b71898, 32'h42f03555, 32'h439f2319},
  {32'hc4e60032, 32'hc314e60a, 32'hc3889257},
  {32'h4422c562, 32'hc0a6d74f, 32'h42501efb},
  {32'hc4a50564, 32'hc39c14ff, 32'hc217961f},
  {32'h44d5f21a, 32'h43e807c6, 32'h4306ceaa},
  {32'hc3df8560, 32'hc33569d3, 32'h438e1c52},
  {32'h445ca4c4, 32'hc1fd65e2, 32'h412e4ff0},
  {32'hc50c2114, 32'hc30e7423, 32'hc32d3e2a},
  {32'h4474b902, 32'hc307fb94, 32'hc14de928},
  {32'hc4091a88, 32'hc2fc2e3c, 32'h43112b66},
  {32'h450725a9, 32'h43f831c5, 32'hc1ad5217},
  {32'hc47e4e14, 32'h43b16522, 32'h42fa3097},
  {32'h44ebee94, 32'hc27a9fc2, 32'h4268c46b},
  {32'hc4a2de15, 32'h43164095, 32'h41f31372},
  {32'h4432d488, 32'h43761942, 32'h42417ac7},
  {32'hc49e8a5a, 32'hc229dd90, 32'h432a7815},
  {32'h44e9a311, 32'h438bd326, 32'h428259ba},
  {32'hc4dc0291, 32'hc3eb8a34, 32'h439736b6},
  {32'h43e151b0, 32'hc2e7b341, 32'h43e8cd1b},
  {32'hc4c4a27a, 32'h431ccb4a, 32'h432df52b},
  {32'h4362c418, 32'h42fec142, 32'h4223e328},
  {32'hc50c39c0, 32'hc39f71ea, 32'h42ddedf7},
  {32'h4440fee2, 32'h438e4426, 32'h4384728d},
  {32'hc44b17e9, 32'hc2e1d26a, 32'h43310ed5},
  {32'hc29d5cbc, 32'h43a46a53, 32'hc3bf820f},
  {32'hc452dd08, 32'h402c0420, 32'h4367cf47},
  {32'h445ef43c, 32'hc390d505, 32'hc2c5ab39},
  {32'hc4d389ca, 32'hc30b1a20, 32'hc2cdb8ff},
  {32'h43cf5960, 32'h41a07a1d, 32'hc35672e1},
  {32'hc4bbe27e, 32'h42ea2521, 32'hc30187d3},
  {32'h43193f43, 32'h423485d9, 32'hc3f45bce},
  {32'h43a4e70e, 32'hc1082bfa, 32'h43f76dea},
  {32'h43e1cd97, 32'hc39d6059, 32'h41d2910d},
  {32'hc3d21dc0, 32'h4365b265, 32'hc3951975},
  {32'h43cd9bb0, 32'h42436909, 32'h431dca98},
  {32'hc4d8c10a, 32'h42fad38d, 32'h43bf36ab},
  {32'h44d6e12b, 32'hc18c812e, 32'hc25ef3e7},
  {32'hc3ca03ec, 32'h43a71e59, 32'h427fdeb4},
  {32'h44c5bfca, 32'h438410dc, 32'h41e66530},
  {32'hc48fef2e, 32'hc315c947, 32'h439b1679},
  {32'h44fcbd6e, 32'hc358de68, 32'h42953b08},
  {32'hc4c7538e, 32'hc39c36e7, 32'hc35af138},
  {32'h43d8594a, 32'hc31d83b0, 32'h435c9be2},
  {32'hc48fc49a, 32'h42edbf47, 32'h43aa8832},
  {32'h444bda20, 32'h422f4397, 32'hc36d0d94},
  {32'hc2950980, 32'hc3cb1776, 32'hc0c2cc40},
  {32'h443a3236, 32'hc3010808, 32'hc329b3c5},
  {32'hc3a8cc78, 32'hc3867393, 32'hc3c71e73},
  {32'h43bb23d5, 32'h4334d2f9, 32'hc396deef},
  {32'hc4627650, 32'hc2826a2e, 32'hc36ac994},
  {32'h45047221, 32'hc30bbe0c, 32'h4328c02c},
  {32'hc4aaab11, 32'hc3318973, 32'h42a90cf3},
  {32'h43eb65f8, 32'h435ee343, 32'hc3f96de9},
  {32'hc44c12ce, 32'h41f40875, 32'h4309b36d},
  {32'h4477685b, 32'hc3b5fe6f, 32'h430ac9c0},
  {32'hc2d2d8e8, 32'hc2d81941, 32'hc3817504},
  {32'h44969ecb, 32'hc26efb12, 32'hc38d6231},
  {32'hc3a05bd6, 32'hc39a47de, 32'h436cf36c},
  {32'h44f1e659, 32'hc3838b34, 32'hc352762e},
  {32'hc4dd1501, 32'hc2917f70, 32'hc2c4492c},
  {32'h42c1bf79, 32'hc3b5d4e0, 32'hc248e2ee},
  {32'hc4adf69a, 32'hc182d33e, 32'hc336afdd},
  {32'h44246dd8, 32'h42c8f388, 32'hc4368834},
  {32'hc4ab1b1b, 32'h4356e866, 32'h436b1cb8},
  {32'h4412076d, 32'h443ba00e, 32'hc3a32694},
  {32'hc3129d30, 32'h4387b2fc, 32'h42a6b7ef},
  {32'h45008712, 32'hc3185e59, 32'h42f928aa},
  {32'hc4ba5085, 32'hc30cca27, 32'hc2b6ffe6},
  {32'h44138ee0, 32'hc324e19a, 32'h441bd848},
  {32'hc2c6eaa0, 32'h43c0fb38, 32'h42c43918},
  {32'h44398bd2, 32'h4213eb47, 32'h43919925},
  {32'hc5028653, 32'h42ce8874, 32'h425f873b},
  {32'h45058fb0, 32'h4306a5e1, 32'h43a0d86c},
  {32'h42a6fdd0, 32'h413efc70, 32'h426e14c4},
  {32'h44e3d56a, 32'h42fd2d69, 32'hc31f956c},
  {32'hc4694b84, 32'hc3a2024e, 32'hc3bf591d},
  {32'h450973b2, 32'hc3a52804, 32'h42fd2ca6},
  {32'hc4ede90c, 32'hc2c6aea9, 32'h42bc4d97},
  {32'h44fb70b2, 32'h4346a5b2, 32'h41bb9d0a},
  {32'hc4cfe652, 32'h431ad56f, 32'h42b49086},
  {32'h442e072e, 32'h43f7ddad, 32'h42d3fe7a},
  {32'hc391087a, 32'h4092f9f4, 32'hc257bf0e},
  {32'h43aa5c5c, 32'hc34d0e98, 32'h42dbbb0d},
  {32'hc438e8e7, 32'h423abe2a, 32'hc2d5c595},
  {32'h4433d401, 32'hc20e27df, 32'hc2609560},
  {32'hc3ae55f8, 32'hc271a98c, 32'h435a780c},
  {32'h45038499, 32'h433479c6, 32'h431cf035},
  {32'hc4d2a753, 32'h4415e17a, 32'h43a84e32},
  {32'h4510ee36, 32'h41acaf4b, 32'h425277de},
  {32'hc4faa85b, 32'h434b27f6, 32'hc28f83a2},
  {32'h44067929, 32'hc30966ef, 32'hc1b030ae},
  {32'hc3e40b56, 32'h4301e903, 32'h428023a9},
  {32'h44f0663d, 32'hc3dffa44, 32'hc35927ad},
  {32'hc4c2176a, 32'hc2c00ae3, 32'hc3c917d4},
  {32'h440e15f8, 32'h4385a9e2, 32'hc2d28684},
  {32'hc4beb26c, 32'hbfc0fe30, 32'hc1e118f4},
  {32'h4432ca37, 32'hc30fddca, 32'hc37d2eeb},
  {32'hc4d7d5d0, 32'hc3fe3f27, 32'h432baa07},
  {32'h4472687e, 32'hc320715f, 32'h4342293c},
  {32'hc3b728b0, 32'h439cb537, 32'h41c0102d},
  {32'h4326a554, 32'hc2da5cb4, 32'hc34ec134},
  {32'hc4bdfd40, 32'hc1f70688, 32'hc09e47ea},
  {32'h448ee2cd, 32'hc2c7f602, 32'hc272706a},
  {32'hc4328dd5, 32'h438356df, 32'h4434360a},
  {32'h445c82f9, 32'h42cc4a13, 32'hc2f23c9a},
  {32'hc4dec624, 32'hc311d21a, 32'h4218c62d},
  {32'h45212fc1, 32'hc28973f0, 32'h433530c7},
  {32'hc49bdf66, 32'h4333c243, 32'h42c495af},
  {32'h44e4a7e7, 32'h42c39222, 32'h41efe602},
  {32'hc5197f80, 32'h431c5df3, 32'h42b509b6},
  {32'h435240dc, 32'h4387eca1, 32'h43b98a8c},
  {32'hc4987096, 32'hc3655874, 32'hc291de4c},
  {32'h44f49214, 32'h433ad214, 32'h41dfb3d4},
  {32'hc5117e68, 32'h4351f4e2, 32'hc3bc38aa},
  {32'h44f2d42b, 32'hc3211cdd, 32'h4246a352},
  {32'hc2b69370, 32'hc387dbe7, 32'hc3b72bdc},
  {32'h443691cf, 32'hc3aecb1b, 32'hc3dcd821},
  {32'hc4d545d0, 32'h43114069, 32'h41a37453},
  {32'h4455a7e4, 32'h43623253, 32'h3ff86f40},
  {32'hc496a7bb, 32'hc38fff31, 32'h4378e3aa},
  {32'h4410be25, 32'h40510105, 32'h435406f2},
  {32'hc35a5a58, 32'hc31c32bd, 32'hc355293c},
  {32'h44970c1b, 32'h427224fb, 32'hc2ef871c},
  {32'hc49ba5c0, 32'h42a79851, 32'hc3d62d8a},
  {32'h43860631, 32'hc341264d, 32'hc3a51968},
  {32'hc51cc3fa, 32'hc3e666b0, 32'hc2a03084},
  {32'h4501e5fa, 32'hc3ae98b0, 32'hc300cac2},
  {32'hc44bdd08, 32'h43dcf918, 32'hc392621b},
  {32'h4357cd72, 32'hc3a4407c, 32'h44379a41},
  {32'hc4462aab, 32'h42676e88, 32'h4098f4f9},
  {32'hc159cf80, 32'hc398ae2a, 32'h43972d2a},
  {32'hc467bf5c, 32'hc36c3315, 32'h439a48cd},
  {32'h450eee00, 32'h43875e8f, 32'h4379152b},
  {32'hc4cab20c, 32'h43648a2f, 32'hc187617e},
  {32'h44e488f4, 32'h4307fa87, 32'h43ec5557},
  {32'hc4525f40, 32'hc325b0a9, 32'hc40f7cb6},
  {32'h43e37ac8, 32'hc3b96c9e, 32'hc2eaf7e0},
  {32'hc5002566, 32'hc1e514dd, 32'hc3b53bb4},
  {32'h44d01658, 32'hc33bd631, 32'h431f9211},
  {32'hc51234ee, 32'hc181e01d, 32'h423d1439},
  {32'h4498402d, 32'hc352143e, 32'hc3211aaa},
  {32'hc3d590a8, 32'h43e969b3, 32'h4321d934},
  {32'h445cb7c8, 32'hc3ebda44, 32'hc35829a1},
  {32'h42db1210, 32'h4298423e, 32'hc39f7d74},
  {32'h45140eca, 32'hc37f1172, 32'hc31d0b98},
  {32'hc4ea47f1, 32'hc1a52ac2, 32'h420ccd50},
  {32'h44acf661, 32'hc3130bdc, 32'hc3948ff1},
  {32'hc3a4430f, 32'h42c01d56, 32'h41dcb0b5},
  {32'h44b42cbc, 32'h439c1e55, 32'h4239611b},
  {32'hc4603214, 32'hc4098636, 32'h432b455a},
  {32'h44848401, 32'hc3153c3c, 32'h4220c3b2},
  {32'hc4bfc592, 32'hc3d4ffe3, 32'hc3017b28},
  {32'h44fe5457, 32'h42f67487, 32'h4398f2aa},
  {32'hc2e1ce20, 32'h434a98a2, 32'hc3ac81c1},
  {32'h4394b918, 32'hc3715e90, 32'h4343a28c},
  {32'hc49d916b, 32'h430d16bf, 32'hc22484e6},
  {32'h44c79a4c, 32'hc20adcc8, 32'hc382085f},
  {32'hc50285f3, 32'hc29e62b0, 32'h43b6a505},
  {32'h44d733f2, 32'hc28d7762, 32'h42bf66c0},
  {32'hc5195945, 32'h432cafe7, 32'hc371937b},
  {32'h44bf8d1e, 32'h43d6dc54, 32'h436cc7ec},
  {32'hc4a43269, 32'hc22c93ec, 32'h4367a92e},
  {32'h436fe6c0, 32'h400b8382, 32'hc2bcc591},
  {32'hc450c9c8, 32'h43155386, 32'h42d35eac},
  {32'h44d18240, 32'h43e7181a, 32'hc3d02bd7},
  {32'hc3af41c9, 32'hc21dc406, 32'h42d70d40},
  {32'h41fcfcc0, 32'h4341d0f3, 32'h429d71b6},
  {32'hc4010f78, 32'h42802924, 32'h42e95eb6},
  {32'h449997b8, 32'h423bae0f, 32'hc294e913},
  {32'hc516854e, 32'h42ddbfe6, 32'h429784e2},
  {32'h443d2fb0, 32'hc0aad16a, 32'h4352b023},
  {32'hc515218c, 32'h439f32de, 32'hc2902aa1},
  {32'h451c4ec6, 32'hc3a8e7d2, 32'hc2f84324},
  {32'hc4a44dd4, 32'hc314067f, 32'hc3c91f5f},
  {32'h44b058b0, 32'h431ffed6, 32'h4389b284},
  {32'hc4ef592a, 32'hc366be8c, 32'hc212df6c},
  {32'h4487ee22, 32'hc3160e21, 32'hc2b7eaa1},
  {32'hc4a77f54, 32'hc2a9ba0a, 32'hc23a4695},
  {32'h44e3fe60, 32'hc2518d7b, 32'h4283c26e},
  {32'hc4fb886e, 32'hc3a934c5, 32'h438f3571},
  {32'h450013bc, 32'hc2521d67, 32'hc175eb48},
  {32'hc50fa39f, 32'hc33ec10b, 32'h43264ae4},
  {32'hc18df800, 32'h441b1c3c, 32'hc30dfe99},
  {32'hc43307e8, 32'h4331f01c, 32'hc2a66286},
  {32'h4452cf10, 32'hc3da5d9f, 32'hc1efb720},
  {32'hc4428a12, 32'hc3d65511, 32'h43cac921},
  {32'h449ecbda, 32'h43949c35, 32'h43616522},
  {32'hc50ec89f, 32'hc284e6cd, 32'hc3ad85e7},
  {32'h45024360, 32'hc1720188, 32'hc33b0410},
  {32'hc40c2aca, 32'h425970fc, 32'h437fe5d9},
  {32'h42881abe, 32'hc3898eed, 32'h43be9a4f},
  {32'h433bd3ef, 32'h4306f3e2, 32'h4369c139},
  {32'h44dc2998, 32'hc2c0a774, 32'h42c8ae3c},
  {32'hc4a72835, 32'h42c0bd0f, 32'h432a98d7},
  {32'h45119378, 32'hc304791e, 32'h43c0f9a0},
  {32'hc413348e, 32'hc26481af, 32'h4330fd44},
  {32'h44b3a0e1, 32'h4362e61f, 32'h42c43a94},
  {32'hc508255a, 32'hc3b5d101, 32'h439d0ddf},
  {32'h449b1596, 32'h43cd1a7d, 32'hc3960b40},
  {32'hc4b8ec9e, 32'hc3fd526c, 32'h42da7cb8},
  {32'h44ca7448, 32'h436d76d8, 32'hc2e63c7d},
  {32'hc47e00e5, 32'h42ba9cba, 32'hc2812c69},
  {32'h44bb163b, 32'hc2be64d0, 32'hc2679004},
  {32'hc4b9b99b, 32'hc2588858, 32'h407d66f0},
  {32'h441c607c, 32'hc3990d26, 32'h42a2791e},
  {32'h43649c1f, 32'hc2e0f3ab, 32'h429bd506},
  {32'h4488a3bd, 32'h4280b94e, 32'hc384b92b},
  {32'hc3016ae0, 32'h424c7aa4, 32'h4214fc8e},
  {32'h44ddc906, 32'hc254fcb3, 32'hc30b1124},
  {32'hc4abff12, 32'h42daa241, 32'h41101d2c},
  {32'h452d5930, 32'hc1af1b6a, 32'hc3720e18},
  {32'hc3c0647c, 32'hc29eaa96, 32'hc375b69a},
  {32'h440e02cd, 32'hc361bfe6, 32'h4386b419},
  {32'hc4d9cbfb, 32'h43ae2897, 32'h4393b64a},
  {32'h448cbe07, 32'hc2032ff0, 32'h4327c1ad},
  {32'hc3c77aa6, 32'hc3841316, 32'h4266e50f},
  {32'h44116ccf, 32'hc391ed9a, 32'h42c36efd},
  {32'hc3a6402e, 32'hc2c1aeb9, 32'h4327838d},
  {32'h4412ca67, 32'hc3aaa1d2, 32'h436fed79},
  {32'hc52ec77e, 32'h43c8202e, 32'h42ba6c20},
  {32'h440beb7d, 32'h4386e601, 32'hbfb06c5e},
  {32'hc4ff3004, 32'hc2c80208, 32'h43a80b67},
  {32'h43f18784, 32'h42c8dea8, 32'hc314003b},
  {32'hc401962c, 32'hc3570783, 32'h43fce894},
  {32'h43911206, 32'hc409e1e9, 32'hc321ae5e},
  {32'hc4982f10, 32'hc2fd5ed2, 32'h43e171c5},
  {32'h441fa818, 32'hc3029402, 32'hc2e029d2},
  {32'hc4306de6, 32'h435ca7c3, 32'hc35bdbb0},
  {32'h449fb48f, 32'h431c4c13, 32'hc26bbea9},
  {32'hc4a72990, 32'h42c8efe1, 32'h42cf0efa},
  {32'h44c53176, 32'h4327d55d, 32'h4230fef3},
  {32'hc5063b79, 32'h4378bc4a, 32'h41e1c4cd},
  {32'h441947f8, 32'hc33d70a4, 32'h42e2caec},
  {32'hc4ae4087, 32'hc2cf80f1, 32'h430e6d5a},
  {32'h44343401, 32'h4201f8b7, 32'hc33b38c2},
  {32'hc50c0f93, 32'hc291db67, 32'hc29eed16},
  {32'hc338a0e8, 32'hc1569600, 32'hc2b00ddf},
  {32'hc42c2d98, 32'h439e6f42, 32'h43480d98},
  {32'h448338ed, 32'hc329f187, 32'hc2c68b1c},
  {32'hc499695d, 32'h42cc2112, 32'h42f04720},
  {32'h44c448c6, 32'hc292b082, 32'hc3796bbf},
  {32'hc3d351a0, 32'hc31280ba, 32'h428c5ee1},
  {32'h4435ca59, 32'h4333d893, 32'h439dede3},
  {32'hc48fc55c, 32'hc3024080, 32'h43998382},
  {32'h419135c0, 32'hc3916b64, 32'hc2eb5cde},
  {32'hc4208e45, 32'h432f1485, 32'h4439d83d},
  {32'h4355f88c, 32'hc353a9e4, 32'hc384f97d},
  {32'hc1240818, 32'hc37cde34, 32'hc2da1fd3},
  {32'h44b969de, 32'h42b19e7d, 32'hc2a9b416},
  {32'hc48eb887, 32'h4293787f, 32'h424d27e5},
  {32'h45003c5c, 32'hc1155c61, 32'hc3a97373},
  {32'hc4f79522, 32'hc3b7dcea, 32'hc2ca30e4},
  {32'h44836c89, 32'hc3d49baf, 32'h43434ba7},
  {32'h43a728d0, 32'h42293bd2, 32'h420c09ab},
  {32'hc46675d2, 32'h4380564f, 32'hc38d8f03},
  {32'h435fa5f8, 32'hc3c3296e, 32'hc30f6b9c},
  {32'hc403e4a4, 32'hc16b89c0, 32'h43ccf429},
  {32'h44190c3c, 32'h42aa70a1, 32'h432925ab},
  {32'hc43e3ddc, 32'h423a89c6, 32'h41d016d6},
  {32'h4513344d, 32'hc302a6d7, 32'hc3ee12ae},
  {32'hc4fc2c98, 32'h42ee6fc6, 32'hc3e42b7d},
  {32'h44e8878b, 32'hc32ea8c0, 32'hc30da5aa},
  {32'hc4ca32c7, 32'h42e82bb3, 32'h42f3ced0},
  {32'h44c9b9f0, 32'h40f93c46, 32'h4308b786},
  {32'hc4584857, 32'hc2691a46, 32'h42d8f74e},
  {32'h441d4b81, 32'h43681db4, 32'hc383c089},
  {32'hc5020dd8, 32'h43903852, 32'hc3e1017e},
  {32'h44354db1, 32'h437ba554, 32'hc2c502dc},
  {32'hc507cf8d, 32'h43a083bc, 32'h430d42e0},
  {32'h444d9e99, 32'h42786223, 32'hc00c1ec1},
  {32'hc500969e, 32'hc3a2c82d, 32'hc1fbe334},
  {32'h44ef7a28, 32'hc3baf42d, 32'hc2a98020},
  {32'hc4fb8ee3, 32'hc17ff93a, 32'hc35d38ee},
  {32'h4519c807, 32'h4315332b, 32'h4327d70f},
  {32'hc32f47d2, 32'hc38b0ce5, 32'h438d9566},
  {32'h4500ec00, 32'h435efef0, 32'hc1fa81ff},
  {32'hc489139b, 32'hc22855bf, 32'h4308203f},
  {32'h44c416fd, 32'h42a00b7f, 32'hc3790334},
  {32'hc480c8be, 32'hc3ce1bec, 32'h4332d7ad},
  {32'h44865d4e, 32'h43053d30, 32'hc333673f},
  {32'hc4f16919, 32'hc283aceb, 32'h42e75717},
  {32'h444315a8, 32'h43408dbd, 32'h423bd2b7},
  {32'hc4ce25b6, 32'hc3462fb3, 32'h434b3430},
  {32'h44758390, 32'hc2f03b38, 32'hc21a760f},
  {32'hc3ef4e4e, 32'hc37cdb86, 32'h438ecc94},
  {32'h44ee63b2, 32'h425b0364, 32'h436abfba},
  {32'hc4d5f1a1, 32'h416aa00c, 32'h4170bb4e},
  {32'h440e9382, 32'h43a54645, 32'hc3be802a},
  {32'hc4e870b8, 32'h42977e04, 32'h4358560c},
  {32'h43c04cdc, 32'hc34f596b, 32'hc299e75c},
  {32'hc4cc74e6, 32'h43d819fd, 32'hc38df02f},
  {32'h430babb0, 32'hc39e013e, 32'h4290f9d2},
  {32'hc4d29008, 32'h43ab481c, 32'h40b10e58},
  {32'h444f48ee, 32'h42107c84, 32'h423c4762},
  {32'hc445ea60, 32'h433b7b52, 32'hc2ebefbc},
  {32'h4416a40e, 32'hc36d7028, 32'h43910d5a},
  {32'hc4ba10ee, 32'h42e986d9, 32'h4215ee96},
  {32'h450c5d0d, 32'hc31db431, 32'h43575dd4},
  {32'hc49a2921, 32'hc35c0fc8, 32'hc29ceae2},
  {32'h452339b2, 32'h430102c4, 32'h41a1b90b},
  {32'hc5083c69, 32'h43388f79, 32'hc3857343},
  {32'h439c434a, 32'h4377abeb, 32'h42a488df},
  {32'hc3d0b069, 32'hc34ed90a, 32'hc242b458},
  {32'h450b6d28, 32'h43cd6d6b, 32'h4254a909},
  {32'hc48c6f35, 32'h41843d97, 32'hc1ea74f6},
  {32'h44e9b672, 32'hc39422f1, 32'h428b8e52},
  {32'hc40cab8c, 32'h41aa6afb, 32'hc2b7d15c},
  {32'h447a4634, 32'h42ef6550, 32'hc1f58544},
  {32'hc4de7c70, 32'h426e117e, 32'hc2fc1ef1},
  {32'h443d451d, 32'hc3238bbb, 32'hc09f7f3f},
  {32'hc46c6368, 32'h43155f50, 32'hc300beac},
  {32'h44113344, 32'hc3583b52, 32'hc31ca22c},
  {32'hc4d83563, 32'h43ce063e, 32'hc24099c8},
  {32'h44a41cda, 32'h439fb3e1, 32'hc2afe87c},
  {32'hc495c765, 32'hc2e44231, 32'hc3aaaadc},
  {32'h43a4247c, 32'h428f8c38, 32'h437e3a9d},
  {32'hc48eeb6b, 32'hc3075ebd, 32'h43964304},
  {32'h44df8c97, 32'h443b4dfe, 32'hc31a87ba},
  {32'hc4fce5f2, 32'h4316d7c0, 32'h43a47002},
  {32'h44c53e96, 32'h42e572b4, 32'h433029a4},
  {32'hc4bf4cf7, 32'h428f20a8, 32'hc2ce5bc3},
  {32'h4425db4c, 32'h42fb6dac, 32'hc299a62e},
  {32'hc4653cf2, 32'hc3e4a120, 32'hc3cc6e7b},
  {32'h44988c9e, 32'h43e6281f, 32'h41cae606},
  {32'hc470ceda, 32'h410d9dfc, 32'hc2da4dc7},
  {32'h44d9faf6, 32'h41a2c701, 32'h43e66883},
  {32'hc48e6cf5, 32'h42d1d997, 32'h40b5e0de},
  {32'h44193a02, 32'h43f36bf7, 32'h43584457},
  {32'hc45c4989, 32'h438b4c0e, 32'hc38cd5aa},
  {32'h4408e796, 32'h41b16368, 32'hc12002a6},
  {32'hc1ac5f80, 32'hc399cbe2, 32'h43dd1e02},
  {32'h4463ea81, 32'h4309a11f, 32'h43a0c950},
  {32'hc510e1be, 32'hc393d149, 32'hc2aa5199},
  {32'h4473bca2, 32'hc070bf93, 32'h433a0677},
  {32'hc488f343, 32'h432265c9, 32'hc2539e45},
  {32'h450b95ea, 32'h42c6ef54, 32'h430e3dba},
  {32'hc3f83640, 32'h427e1675, 32'hc357e586},
  {32'h44f1f810, 32'hc3086b00, 32'hc35a5f9a},
  {32'hc4967ed2, 32'hc1cfce9a, 32'hc232adeb},
  {32'h4423e5ac, 32'hc30eb59a, 32'hc445a198},
  {32'hc363d358, 32'h416e3b51, 32'h437f588c},
  {32'h44099668, 32'hc213fec0, 32'hc32d58cf},
  {32'hc4737f6f, 32'hc1946e4e, 32'hc275c9ac},
  {32'h44cbb6e4, 32'h42644545, 32'hc36226c3},
  {32'hc4d95ecf, 32'hc0c2e504, 32'h42f3fc5c},
  {32'h44fbcd71, 32'h4360258e, 32'h42bfea4a},
  {32'hc4aadc60, 32'h44233e13, 32'h42e8d79a},
  {32'h42a1bab2, 32'hc1ed51a6, 32'h42862568},
  {32'hc4e69aaa, 32'hc3d0e334, 32'h43f77885},
  {32'h44895ec6, 32'hc33b7e8e, 32'hc358fd36},
  {32'hc4bf1f2a, 32'h42c5592b, 32'hc3a9d099},
  {32'h443f1182, 32'hc0227418, 32'h431c67cf},
  {32'hc4d44a3e, 32'hc2355c74, 32'h428fc1c8},
  {32'h44d89f21, 32'h4341b5c4, 32'h4315f532},
  {32'h4375c8af, 32'h4350a6ed, 32'h431c6f0b},
  {32'h44aac7bc, 32'h43bbc883, 32'h43e95351},
  {32'hc49391ec, 32'h430b1e8a, 32'h43130ebf},
  {32'h4463d517, 32'h430c5265, 32'hc377cd73},
  {32'hc3c61710, 32'hc4358773, 32'h43215e40},
  {32'h441a6ae8, 32'hc0f9da95, 32'hc364502a},
  {32'hc4d8c865, 32'hc3a40891, 32'hc3b6a22a},
  {32'h450f6f07, 32'h433e3ee6, 32'h428bb61e},
  {32'hc4e34cb2, 32'hc20e0b90, 32'hc3255bb7},
  {32'h43805216, 32'hc31a4ad4, 32'h43702b01},
  {32'hc4a06a77, 32'hc167b346, 32'h43eb78b1},
  {32'h44db4786, 32'h436585f6, 32'h43580567},
  {32'hc3ee9ef0, 32'hc1ae109f, 32'hc215b337},
  {32'h445dee32, 32'hc251a270, 32'h42b4e3e8},
  {32'hc4ab9ae6, 32'h43958d31, 32'h431fffad},
  {32'h44f2c436, 32'hc3724472, 32'h42a78700},
  {32'hc503a1eb, 32'hc344d540, 32'h433eba5d},
  {32'h44e0191b, 32'h438d3abc, 32'h4245df15},
  {32'hc3191000, 32'h4331dd81, 32'h4417cad2},
  {32'h43e6daf2, 32'h419dd929, 32'h426edaff},
  {32'hc4b05c1f, 32'hc3ac41b5, 32'h41b8285c},
  {32'h443324f8, 32'hc35f4723, 32'h411b8553},
  {32'hc492d6d1, 32'hc30f5d5a, 32'hc16094f4},
  {32'h446bd7db, 32'h43aaa0f5, 32'h43ec51ae},
  {32'hc4b60508, 32'h42023cfe, 32'h43758c11},
  {32'h449fd8ec, 32'hc27921c4, 32'h4141e87f},
  {32'hc4feb36e, 32'hc387ffb2, 32'h43b1527d},
  {32'h4403a07e, 32'h42e48f33, 32'hc327af2b},
  {32'hc47430f0, 32'h4353f98b, 32'h42e4599e},
  {32'h4409331d, 32'h4402ea28, 32'h43edfbec},
  {32'h411cfdb0, 32'h43ad4d58, 32'h43193316},
  {32'h43b481e4, 32'h43911d92, 32'h430a0d94},
  {32'hc48dce50, 32'hc31a2308, 32'hc303bc96},
  {32'h44f483ad, 32'hc366e7da, 32'h43a6b293},
  {32'hc4deaca6, 32'hc40672da, 32'hc3160c1d},
  {32'h44f758ca, 32'h431c441d, 32'h40833dea},
  {32'hc4121c84, 32'hc3340015, 32'h432dd335},
  {32'h450b7e99, 32'h41d280be, 32'h43148245},
  {32'hc4523a62, 32'h431e0d9a, 32'hc24412cc},
  {32'h4483dfee, 32'h4332df2f, 32'h4260cbf3},
  {32'hc492cdc9, 32'hc0459476, 32'h42a37f4f},
  {32'h44f351b1, 32'h430f8ecc, 32'h43889ea6},
  {32'hc4e0e9b2, 32'hc2e9cd6e, 32'hc2dd065a},
  {32'h44aedda3, 32'h42b7bdde, 32'h42b7b170},
  {32'hc49c0f3e, 32'h41fc4a7a, 32'h4285d19a},
  {32'h45105576, 32'h436b9dcf, 32'h441210df},
  {32'hc4a896b5, 32'h433d776a, 32'h435d6829},
  {32'h4457f0af, 32'hc2d1b7b3, 32'h418c02c0},
  {32'hc38909de, 32'h43200ae8, 32'h43045f95},
  {32'h44da5a7d, 32'h42dcbfe7, 32'hc32195e1},
  {32'hc4c3fdac, 32'hc212ec62, 32'hc214003c},
  {32'h45083a82, 32'hc2c404d2, 32'h42159726},
  {32'hc4f62e87, 32'hc237f557, 32'h43a16762},
  {32'h44bf622d, 32'h41cb4f50, 32'hc1e19810},
  {32'hc4d34137, 32'h43058741, 32'h42cecf94},
  {32'hc0df3100, 32'h43adcb8f, 32'h42e40ecc},
  {32'hc4d75cc0, 32'hc39489f7, 32'hc34c2e7e},
  {32'hc294f29c, 32'hc2448761, 32'hc331da89},
  {32'hc4c04243, 32'h4417e179, 32'hc3d82270},
  {32'h43cc7d26, 32'h435225f9, 32'h430f2813},
  {32'hc4836005, 32'h4121fbba, 32'hc4175d33},
  {32'h44972019, 32'h420a5b83, 32'h431a19cc},
  {32'hc4b4efc4, 32'hc3d72efc, 32'hc29d0c1a},
  {32'h44608588, 32'hc14b8b7f, 32'hc33ff91e},
  {32'hc3890760, 32'hc34a480d, 32'h440ff160},
  {32'h44f34c44, 32'h423bbc82, 32'h40d23127},
  {32'hc4a211fe, 32'h4286273d, 32'hc38000af},
  {32'h446c67be, 32'h424e0bfd, 32'h439e7fb0},
  {32'hc4447cea, 32'h43bc4e7c, 32'h426022b0},
  {32'h44e1a357, 32'hc394f1e5, 32'h42d250d0},
  {32'hc489c59d, 32'hc410b839, 32'h425e7340},
  {32'h44ce8d64, 32'hc24553ce, 32'h433e4990},
  {32'hc2210558, 32'h419cdf65, 32'hc33495f3},
  {32'h444d525f, 32'hc387d671, 32'hc2c43511},
  {32'hc508135e, 32'h418da499, 32'h4115e8cb},
  {32'h449416b4, 32'hc3151d9e, 32'h436d15a7},
  {32'hc424a17c, 32'h42e99ada, 32'h42ca83f2},
  {32'h432b5b30, 32'h4226e70a, 32'hc3717737},
  {32'hc4ef14d5, 32'hc38f0a68, 32'hc3a12e36},
  {32'h424d37a0, 32'h42137014, 32'h42dd9af6},
  {32'hc50cf8b4, 32'hc42655e2, 32'h43277274},
  {32'h448c47e3, 32'h42885350, 32'hc307d258},
  {32'hc443b236, 32'hc309cae2, 32'h3fbdc224},
  {32'h4351f5a0, 32'h42450312, 32'hc2304e4c},
  {32'h4313d9e4, 32'h43022ea8, 32'hc35ca64b},
  {32'h4397eb38, 32'h431b3a84, 32'h43d06b20},
  {32'hc403f392, 32'hc28c40f5, 32'hc38c6273},
  {32'h44cdce72, 32'hc3922f63, 32'hc3768238},
  {32'hc4651723, 32'hc3ae9125, 32'hc2e87749},
  {32'h44b86e18, 32'hc363af1b, 32'h432a9688},
  {32'hc421e305, 32'h43a13142, 32'h43697cc9},
  {32'h446081fb, 32'hc307c5a0, 32'hc33f50e2},
  {32'hc4fb0afb, 32'h4353e8dd, 32'hc38ef5e0},
  {32'h448b8e01, 32'h424b2ea7, 32'h431ebda8},
  {32'hc3fd0ca8, 32'hc3056fac, 32'h43e3dce8},
  {32'h44efeedc, 32'hc3f71584, 32'hc1d25a4b},
  {32'hc4fb6a44, 32'hc2ccf023, 32'h410f30c0},
  {32'h4509bd8e, 32'h4362cbf6, 32'hc2977db7},
  {32'hc499eeb8, 32'hc40554a0, 32'h42d97579},
  {32'h4502babc, 32'h421b0bf9, 32'h4335d7b9},
  {32'hc4ab381a, 32'hc1434ac4, 32'hc37ad0b8},
  {32'h45028cc0, 32'h43863da1, 32'hc387ca67},
  {32'hc424216a, 32'h4121c22f, 32'hc2a82cc3},
  {32'h44871ea0, 32'h42d5aafd, 32'h43882ed2},
  {32'hc40d9628, 32'hc3f407ae, 32'h43baf19f},
  {32'h44291a42, 32'h4241d2cd, 32'hc28a5fe5},
  {32'hc50ab8db, 32'hc3012694, 32'hc3c1ffec},
  {32'h43fb7c81, 32'hc30003d6, 32'h4303b86a},
  {32'hc4b80f8c, 32'hc24293dc, 32'hc3743ac6},
  {32'h440d23cc, 32'h4394ed38, 32'h434eaff1},
  {32'hc441a5b9, 32'h4275ee3a, 32'h430dfa68},
  {32'h449b0456, 32'hc308e9c6, 32'hc3076a24},
  {32'hc4be65d3, 32'h426f0d44, 32'h43c31991},
  {32'h43b67968, 32'hc101fa87, 32'h4244c404},
  {32'hc4e7352a, 32'hc3fcad3b, 32'hc38a299f},
  {32'h44f6f905, 32'h434fe2c1, 32'h431518e6},
  {32'hc4e71411, 32'hc36091c6, 32'h432a34ce},
  {32'h439cd6a1, 32'hc39fe3f0, 32'h436ee2ae},
  {32'hc4f19e6a, 32'hc2f93429, 32'h43844ed1},
  {32'h4430c223, 32'hc3cbc32f, 32'hc10cb17b},
  {32'hc416eb20, 32'hc0e4d910, 32'hc2f7ffcd},
  {32'h433cc176, 32'h430c13da, 32'hc2c1ddf9},
  {32'hc492bc9a, 32'hc2afa973, 32'h43bc9589},
  {32'h450d4c27, 32'hc3058658, 32'hc3b80d67},
  {32'hc3cc4eee, 32'h438bfc77, 32'h430cb3a4},
  {32'h44babd44, 32'hc2e4a2c6, 32'h43646c5f},
  {32'hc488f2ec, 32'h439b28cc, 32'hc16dc62f},
  {32'h444961d8, 32'h43174ff4, 32'h43391bf4},
  {32'hc4d8b3b0, 32'hc3b52ea1, 32'h43b029ef},
  {32'h4480e9a0, 32'hc0cf1d21, 32'h429ec1ac},
  {32'h42a01200, 32'hc2960188, 32'h420f0832},
  {32'h449b7b7f, 32'hc2041514, 32'h430751f9},
  {32'hc4441b77, 32'h436549a6, 32'h4323d3e1},
  {32'h44cd858c, 32'h438c23ca, 32'hc32e69a4},
  {32'hc4a6d51e, 32'hc28702ba, 32'hc33a069e},
  {32'h4502c46e, 32'hc30a2ae9, 32'hc2f7124d},
  {32'hc4e63ccc, 32'h43559e58, 32'hc3940dc6},
  {32'h450bbdd5, 32'hc25affb6, 32'hc16591a7},
  {32'hc44ed30c, 32'h42a5c078, 32'h435a072a},
  {32'h440fc27a, 32'h431ffcf8, 32'h421e725b},
  {32'hc493b0f3, 32'h4346035b, 32'hc21031a7},
  {32'h450f0d9e, 32'h434ee2b8, 32'h4167fb30},
  {32'hc4b25bce, 32'h4371beca, 32'hc1cbb1f3},
  {32'h44cf2c42, 32'hc32fb442, 32'h42b0041f},
  {32'hc49bf947, 32'h4256e379, 32'h435e92f4},
  {32'h4407950e, 32'h43bc44d4, 32'hc3293729},
  {32'hc4897c28, 32'h424f0d2b, 32'hc27c5a45},
  {32'h44548658, 32'hc3a0e346, 32'hc2712762},
  {32'hc4a07a58, 32'hc22bc3fa, 32'hc1361e46},
  {32'h44d759a0, 32'h4359ccfb, 32'h421817e0},
  {32'hc44597a8, 32'hc3af3396, 32'h439581d2},
  {32'h450534e9, 32'h4400ea3d, 32'hc3c231f5},
  {32'h43122d7f, 32'h41be41c8, 32'h3f2f430f},
  {32'h44da0822, 32'hc2033573, 32'hc33c10c5},
  {32'hc4e10dd3, 32'h43501492, 32'hc402251c},
  {32'h44ec9242, 32'hc37fecda, 32'h428e63e9},
  {32'hc50d635c, 32'h3f51cfbf, 32'hc338cc7d},
  {32'h445368dd, 32'hc333d73d, 32'h42185946},
  {32'hc502b2b4, 32'h43665002, 32'hc1b2bb64},
  {32'h4416fc78, 32'h430d5676, 32'h431e3003},
  {32'hc4b1b482, 32'h43af6b6b, 32'h4308a4fc},
  {32'h43584d40, 32'hc2ead241, 32'h42c98ff8},
  {32'h41a63408, 32'hc152d7ae, 32'hc216c759},
  {32'h430e70ac, 32'hc4413adf, 32'h42b7a30d},
  {32'hc4a49516, 32'h42e88ffe, 32'h43b1a366},
  {32'h44980fec, 32'h42d24996, 32'hc3b22f88},
  {32'hc4f4d929, 32'hc2994a6b, 32'hc1221c4a},
  {32'h44861062, 32'h432ff816, 32'h431dc855},
  {32'hc4f3db2a, 32'h42aa5248, 32'hc19a055a},
  {32'h442e6bbd, 32'hc337b721, 32'h428d069b},
  {32'hc5268034, 32'hc384901b, 32'h43b50af1},
  {32'h44ae4557, 32'h41fadd50, 32'hc3170dce},
  {32'hc4ebf067, 32'hc319615a, 32'h411b373c},
  {32'h442bf77a, 32'hc2a09f12, 32'hc2a57b06},
  {32'hc4c72f17, 32'hc37197a0, 32'hc385e567},
  {32'h445cf376, 32'h41441471, 32'h42648a9a},
  {32'hc5010b98, 32'h434d7fc6, 32'hc291d845},
  {32'h448ba692, 32'hc1a15c60, 32'h43d835b9},
  {32'hc5055c77, 32'h435a2f3f, 32'hc319e7db},
  {32'h4445d94e, 32'hc315ce51, 32'hc320e4d4},
  {32'h43943d60, 32'h43435f4a, 32'hc2ab2542},
  {32'h428c9240, 32'hc324d16d, 32'hc32a71bf},
  {32'hc4a3d471, 32'h431aaa14, 32'h42b93572},
  {32'h44ea464c, 32'h42a66eab, 32'hc2ebe56c},
  {32'hc4e00aba, 32'hc35bd407, 32'h40c1ba42},
  {32'h450abc8d, 32'h42f44e1d, 32'h430393b1},
  {32'hc42fbda3, 32'h42b7108f, 32'h44050a4d},
  {32'h43430a6e, 32'h437adb7a, 32'h42d3545f},
  {32'hc4ccfe4a, 32'h40ca141c, 32'hc2a57582},
  {32'h449cda51, 32'h428a2a87, 32'h40cb02e1},
  {32'hc4f11bd2, 32'h411fc258, 32'hc300b8bf},
  {32'h44d016c3, 32'h41ba97ff, 32'hc328f10b},
  {32'hc5168c0e, 32'hc24d88ea, 32'h4285947c},
  {32'h449a0bc1, 32'h41701dbf, 32'hc374ae45},
  {32'hc3f66ec0, 32'h40f9666e, 32'h423d6287},
  {32'h449fb21f, 32'hbf2076e9, 32'h4372edc3},
  {32'hc49ffb71, 32'hc34c5bab, 32'h420330de},
  {32'h44c60eba, 32'h438a113f, 32'hc1a79eea},
  {32'hc32f4d60, 32'hc2e277d8, 32'hc39e2038},
  {32'h44285429, 32'hc2742788, 32'h42c88b25},
  {32'hc484b35c, 32'h4317dde9, 32'h429e4ce0},
  {32'h443ce0e8, 32'h43bbdebe, 32'h4386dedd},
  {32'hc367c7f0, 32'h423f41f2, 32'h42b52cf5},
  {32'h44c958f2, 32'h434b8a61, 32'h428037ca},
  {32'hc3f951ea, 32'hc3c77bb8, 32'h4405a427},
  {32'h445cd08a, 32'hc2847a3b, 32'hc38ec609},
  {32'hc4e2dff3, 32'hc29f18e4, 32'h41f509cb},
  {32'h4503e332, 32'hc22443c9, 32'h4411124a},
  {32'hc4245846, 32'hc39e5038, 32'h43ca076f},
  {32'h44822fea, 32'h40ac3aca, 32'h438728d4},
  {32'hc4a4ecdc, 32'hc3d2c819, 32'hc31cfa90},
  {32'h440f5c26, 32'h434449fc, 32'h41cc0336},
  {32'hc49618b6, 32'h42a900af, 32'hc2e6591a},
  {32'h450c6598, 32'hc2c9e126, 32'hc3aaeecd},
  {32'hc45d3ed2, 32'hc2e40920, 32'hc252dae6},
  {32'h45059ae7, 32'hc2839bea, 32'hc2dc56d0},
  {32'hc3de9600, 32'h431cc6a1, 32'h43a6f168},
  {32'h43bfb628, 32'h43ab2237, 32'hc39a1961},
  {32'h42d90c40, 32'hc326e96f, 32'h428b4d4a},
  {32'h451dfa8f, 32'h430579b4, 32'hc38c9e88},
  {32'hc4888e5d, 32'hc113c4e9, 32'hc3a32174},
  {32'h43bbf390, 32'hc33d053b, 32'hc3649488},
  {32'hc46f2d52, 32'h42091687, 32'h41d2cb14},
  {32'h44f519e3, 32'h4399be8d, 32'hc1c93c40},
  {32'hc49611d6, 32'hc34d7f63, 32'hc31c6875},
  {32'h44ba7fc4, 32'h43bb0358, 32'h41e63624},
  {32'hc3e3c1ae, 32'hc39e7569, 32'h438b29c7},
  {32'h448fd2f2, 32'hc3816c3a, 32'hc31d1a71},
  {32'h424b06c0, 32'h4305df0d, 32'h40fbe2a8},
  {32'h44011468, 32'h4271d1fc, 32'h4303370a},
  {32'hc49f4bdc, 32'hc3643e40, 32'h432b1941},
  {32'h44e45ee9, 32'hc2c393cd, 32'hc3ab38ba},
  {32'hc4d64cf4, 32'hc2ffb552, 32'hc3fba95f},
  {32'h43987790, 32'h439f8c1c, 32'hc35b1ebb},
  {32'hc4c73a58, 32'hc35f9c26, 32'hc201916c},
  {32'h433b1230, 32'h43d26478, 32'hc2594334},
  {32'hc43d1e41, 32'h433d9910, 32'hc3a0d809},
  {32'h45100396, 32'h429e880a, 32'hc35f3a48},
  {32'hc4ff6108, 32'h435b7239, 32'h436764eb},
  {32'h44fbfc60, 32'h42e18352, 32'hc31e3a80},
  {32'hc4fe4920, 32'hc35bdac0, 32'hc34b634c},
  {32'h43f7bc40, 32'h42f8be80, 32'h42e0773d},
  {32'hc4a4adeb, 32'h431d5c3f, 32'hc33232e6},
  {32'h439ec7fe, 32'h436d5800, 32'hc336d58d},
  {32'hc4f02e66, 32'h421f0138, 32'hc28d64d9},
  {32'h44aeaba4, 32'hc1fc56e8, 32'hc2d0be02},
  {32'hc4c533c3, 32'hc3232fb9, 32'hc37aecc2},
  {32'h45001273, 32'hc3a384d5, 32'hc35655a2},
  {32'hc39d1736, 32'hc2265526, 32'h43930e21},
  {32'h449220dd, 32'h4293a769, 32'hc2a9fe11},
  {32'hc3808c38, 32'hc3dedc3a, 32'h43d5209f},
  {32'h4319ab9c, 32'h4415bebb, 32'hc3c78ec3},
  {32'hc50809a1, 32'h43e189c3, 32'hc36753c6},
  {32'h44b8014c, 32'hc30ee400, 32'hc395702f},
  {32'hc4810401, 32'hc2ce5bf6, 32'hc3190dae},
  {32'h4508445a, 32'hc363cccf, 32'h42d5f761},
  {32'hc4a6bc12, 32'hc3b747c7, 32'hc195c8d0},
  {32'h446d5bb5, 32'h43407734, 32'h42d622ae},
  {32'hc32e0930, 32'hc2632af2, 32'h42c64891},
  {32'h44089086, 32'hc20b5877, 32'h3f5ca020},
  {32'hc4f8682f, 32'hc34b1f38, 32'h421603ae},
  {32'h4428226c, 32'hc345648f, 32'hc3351f8f},
  {32'hc402063a, 32'hc2c98e21, 32'h42a2a9d4},
  {32'h4492bbf4, 32'hc29c0638, 32'hc3cd305a},
  {32'hc415f3c2, 32'h436bbe61, 32'hc36f87e0},
  {32'h44ac4898, 32'h43506e03, 32'hc386026b},
  {32'hc3e3b084, 32'h41d63b9b, 32'hc2d834c5},
  {32'h45068b17, 32'hc350d741, 32'h43cef98b},
  {32'hc31265f2, 32'hc33001ef, 32'h42aeff83},
  {32'h44fd9073, 32'h41e81e4d, 32'hc2ebb74b},
  {32'hc50fd88c, 32'hc384fafc, 32'hc2ed2377},
  {32'h450ea4c5, 32'h42757251, 32'hc3189788},
  {32'hc4751462, 32'h4234801c, 32'hc3fe6241},
  {32'h44251692, 32'hc30f12b6, 32'hc2397cf8},
  {32'hc4ad61d6, 32'h43a61359, 32'hc30d493c},
  {32'h444273e2, 32'h414056c2, 32'hc342569d},
  {32'hc4792415, 32'h43a28e3e, 32'hc1bd6ddf},
  {32'h4260c9a0, 32'hc35045fc, 32'h42becbe0},
  {32'hc3fa1885, 32'hc2628160, 32'hc2be1b22},
  {32'h44ec754c, 32'hc307d50f, 32'hc2602bf5},
  {32'hc3a72b80, 32'h4266d876, 32'hc3130662},
  {32'h449a6470, 32'h4258f71b, 32'hc31af635},
  {32'hc4dd9b5d, 32'h4286f669, 32'h41bd5f56},
  {32'h42fa0300, 32'hc18a05a7, 32'h43a01d80},
  {32'hc5068037, 32'hc30869b3, 32'h433d582d},
  {32'h45137875, 32'hc174c800, 32'h4129ac64},
  {32'hc4934f8c, 32'hc26dc4b2, 32'h43558cad},
  {32'h4404524a, 32'h42d5c58b, 32'h4304c90b},
  {32'hc45469e0, 32'h433c36e9, 32'h433afb6c},
  {32'h43b0007c, 32'h42480645, 32'h438ec2a5},
  {32'hc4a71891, 32'hc38da044, 32'h42ce26f1},
  {32'hc3b18aaf, 32'h439d61bf, 32'hc39ca320},
  {32'hc4b5d497, 32'hc1b1fa5f, 32'hc3a7d663},
  {32'h4483b211, 32'h43785adc, 32'h43106fd4},
  {32'hc4f3d940, 32'h432b084f, 32'h4399d40d},
  {32'h4495f38c, 32'hc32c47cb, 32'hc2dfab94},
  {32'hc4db5bd5, 32'h431ad059, 32'h43cf611a},
  {32'h45166d95, 32'hc29a2875, 32'hc2f3bcb0},
  {32'hc4fb5eb3, 32'hc36d82cb, 32'hc39497a2},
  {32'hc35c4134, 32'hc30ada60, 32'h439e3787},
  {32'hc50c621f, 32'h4271cb69, 32'hc352c042},
  {32'hc41e68aa, 32'hc319ec14, 32'hc2b67ab1},
  {32'hc4ad04c3, 32'h419fdfbb, 32'hc0977e37},
  {32'h447625f6, 32'hc3de275e, 32'h43056949},
  {32'hc43a8dba, 32'hc40d7ab4, 32'hc3220ec8},
  {32'h44d0569f, 32'h42c6ed36, 32'hc2b5724a},
  {32'hc407a682, 32'hc3260291, 32'h3f549a60},
  {32'hc3108068, 32'hc32cc927, 32'h400cb9ae},
  {32'hc2d96a1c, 32'hc2dc84e9, 32'h42bf38e5},
  {32'h44db67ac, 32'hc28d97ca, 32'hc384246b},
  {32'hc4e35b2d, 32'hc3374ecb, 32'hc352d5b9},
  {32'h44e12eea, 32'h42a6a225, 32'hc3b80c66},
  {32'hc4f022af, 32'h43eff385, 32'h43a14688},
  {32'h445bfa10, 32'hc3397bff, 32'h43f7655b},
  {32'hc41e1c7a, 32'hc2ba518c, 32'hc323077c},
  {32'h43fd3c98, 32'hc393bef9, 32'h434bf8a6},
  {32'hc507c0c5, 32'hc32af038, 32'hc244e7d5},
  {32'h4453bfe2, 32'hc277caed, 32'h43c14f70},
  {32'hc4f825a1, 32'hc3c7ad16, 32'hc2a52152},
  {32'h44a66070, 32'h42aeaa60, 32'h4347a633},
  {32'hc3db28ea, 32'h4275bcfb, 32'hc239587c},
  {32'h44b7d182, 32'hc33575c8, 32'h4351d401},
  {32'hc4bed443, 32'h42eb57e6, 32'h43c8422e},
  {32'h43c98f44, 32'h43a9ac86, 32'h43b31446},
  {32'hc4a19fc6, 32'hc36a57c8, 32'hc14b3507},
  {32'h44a830d1, 32'h42b51f66, 32'hc30eaa19},
  {32'hc5066731, 32'hc3b93edd, 32'hc38324f1},
  {32'h436e0c18, 32'h42fed802, 32'h43c0db47},
  {32'hc4c11d9a, 32'hc3bef115, 32'hc3351206},
  {32'h4458cf7e, 32'h43a1ccdb, 32'hc291fdff},
  {32'hc4ae1576, 32'h429529fc, 32'hc3087f92},
  {32'hc0e67600, 32'h43033b4c, 32'h432d3058},
  {32'h44004e24, 32'h4305d6c8, 32'h438532ec},
  {32'hc4e6c63a, 32'hc3687822, 32'hc29f074a},
  {32'h43fa77c8, 32'h43c360e5, 32'hc1fddb29},
  {32'h43b4d19f, 32'h42d33697, 32'h3f096034},
  {32'h448da4b4, 32'hc23e5e18, 32'hc367af3f},
  {32'hc4de20b6, 32'h4391ac54, 32'h43872815},
  {32'h43d7a26c, 32'hc2a0b3d9, 32'h43e3fc9c},
  {32'hc4e82902, 32'hc2685ae4, 32'hc2a48415},
  {32'h44caec3b, 32'h42b6c921, 32'hc33281ba},
  {32'hc42953a1, 32'hc38925d0, 32'hc4119b21},
  {32'h42953458, 32'h43bb2d71, 32'h431802c1},
  {32'hc441c108, 32'h438c372c, 32'hc2ce7234},
  {32'h43bad2d8, 32'hc39dbfb2, 32'h42a3097c},
  {32'hc48f724c, 32'h434c5964, 32'h42139916},
  {32'h4510cd8d, 32'h4394c4c2, 32'h4341308f},
  {32'hc4eca82c, 32'h436f1af1, 32'hc318c54c},
  {32'h450a79d2, 32'h4409ad18, 32'hc4052c4d},
  {32'hc457f3a6, 32'h43ad71c3, 32'h42271068},
  {32'h44a88854, 32'h4258dfa6, 32'h43913acf},
  {32'hc488866a, 32'hc31d98ff, 32'hc404070f},
  {32'h439d04b8, 32'hc1dba070, 32'h42d17a3f},
  {32'hc4b97dc9, 32'h4280899a, 32'hc2d3f950},
  {32'h44998ee4, 32'hc3763b9a, 32'h4347e167},
  {32'hc287940e, 32'hc3432547, 32'hc3d84e7b},
  {32'h43cb1aa2, 32'hc1f440d7, 32'hc2a63b51},
  {32'hc4696a40, 32'hc3a42e04, 32'h4394bcd8},
  {32'h440dd153, 32'hc384f185, 32'hc347183e},
  {32'hc4f3fc38, 32'hc1a472a4, 32'hc3278495},
  {32'h44827469, 32'hc2a9f4d9, 32'h43801124},
  {32'hc4244c0c, 32'h42bc9da6, 32'hc3f5e223},
  {32'h44a92c78, 32'h42e0aeb0, 32'h436ee165},
  {32'hc4d575cc, 32'hc354887e, 32'h42e774dd},
  {32'h44b70f82, 32'h422ef6c1, 32'hc327c78d},
  {32'hc50201e1, 32'hc2c9ed35, 32'hc3d9c174},
  {32'h4443c340, 32'hc394504e, 32'hc2fc845c},
  {32'hc4841deb, 32'hc312738a, 32'hc406bf09},
  {32'h44f26d40, 32'h43497f8c, 32'h41fa41e2},
  {32'hc38a44ea, 32'h4295cfc8, 32'h4351b758},
  {32'h450f9fd2, 32'hc25c33d9, 32'hc388f51b},
  {32'hc50fbb8a, 32'h439d1f43, 32'h43291f58},
  {32'h45030be4, 32'h4415d2e3, 32'hc1ae3045},
  {32'hc509c353, 32'hc2b498ae, 32'h433d6184},
  {32'h447c4bb4, 32'hc24c06cb, 32'h4339494c},
  {32'hc492208c, 32'h43b4402a, 32'hc2c5a5e7},
  {32'h44eec8e7, 32'hc39d79b2, 32'hc2f5c9a1},
  {32'hc4c0a14f, 32'h43c08c5f, 32'hc2935606},
  {32'h44167da6, 32'h4408eb36, 32'hc3d40687},
  {32'hc429295c, 32'hc25f6913, 32'hc39113d2},
  {32'h44ee04ce, 32'hc289a8a1, 32'h4278523e},
  {32'hc4d93eda, 32'hc319a501, 32'h4308c819},
  {32'h448d0479, 32'hc345e586, 32'hc10d15f0},
  {32'hc456c0c8, 32'hc393d667, 32'h438f1486},
  {32'h43865e90, 32'hc4032f16, 32'h43240187},
  {32'hc4f0aea9, 32'h439d353f, 32'h4313a405},
  {32'h43d3594c, 32'hc33073d3, 32'hc38ee0c1},
  {32'hc4ecf44d, 32'hc30fbf68, 32'h4422eeba},
  {32'h4414731a, 32'hc2211023, 32'hc418ab5a},
  {32'hc4c07c19, 32'hc305e487, 32'h4383f689},
  {32'h448fddf9, 32'h433bc840, 32'h43c58cb6},
  {32'hc4c1e68a, 32'hc2621b40, 32'h41e27bcd},
  {32'h437fc87b, 32'h426be528, 32'hc35f7b85},
  {32'hc43171f9, 32'hc3c76b8b, 32'hc3c77e5a},
  {32'h43e52d87, 32'h431a9aea, 32'h42b579f0},
  {32'hc50a4164, 32'h43321209, 32'hc2dd1fe0},
  {32'hc2bcc440, 32'hc354fd58, 32'h44465199},
  {32'h430e33c9, 32'h41b99687, 32'h41bfc532},
  {32'h44f16391, 32'h432098cd, 32'hc29f03c8},
  {32'hc431cb43, 32'hc34ce55e, 32'hc35fd123},
  {32'h44f9911e, 32'h434dfb84, 32'h4347e260},
  {32'hc4b9560d, 32'hc3025e5c, 32'hc1de200b},
  {32'h44bd4b0d, 32'hc2d09901, 32'h436e27b7},
  {32'hc496ac79, 32'h430579b2, 32'hc32202c8},
  {32'h445ca24a, 32'h43063e07, 32'hc38a2964},
  {32'hc4ee4dce, 32'hc3ba97d4, 32'h43c075fa},
  {32'h40fc8b00, 32'h436ffa01, 32'hc3995e68},
  {32'hc43912da, 32'h430cabfe, 32'hc34fe0fc},
  {32'h43ee78ec, 32'h439f9aef, 32'hc2cb6446},
  {32'hc3bc1871, 32'hc35222ce, 32'h42fdcc4a},
  {32'h4508cf40, 32'h43bcbac3, 32'h43bca977},
  {32'hc43a73df, 32'hc1e36188, 32'hc3024599},
  {32'h45202bc7, 32'hc3b85d18, 32'hc21c691b},
  {32'hc37060d0, 32'hc3e56823, 32'hc37c3177},
  {32'h445f803c, 32'hc14b3fb3, 32'hc343a9c4},
  {32'hc30f84d9, 32'h43c251ea, 32'h437d06e2},
  {32'h44be1db2, 32'h43649113, 32'h43bc7b1f},
  {32'hc5060abe, 32'h4349c9fc, 32'h4341bd59},
  {32'h437b1718, 32'h43523564, 32'hc3994845},
  {32'hc5031a13, 32'hc2dc0288, 32'hc3078001},
  {32'h440f49c2, 32'h4264d256, 32'hc338c324},
  {32'hc5083938, 32'hc33d8813, 32'hc0ad3df1},
  {32'h44110fc8, 32'h4201d0c8, 32'hc2f69be0},
  {32'hc46a4851, 32'hc325de83, 32'hc36dd451},
  {32'h44fedd10, 32'h438631ce, 32'hc28980b6},
  {32'hc5106963, 32'hc32d0c01, 32'hc3d17be5},
  {32'h44804837, 32'hc257536b, 32'hc38636d0},
  {32'hc509ca63, 32'h436f1ce1, 32'hc2bb0da5},
  {32'h4383cb48, 32'hc213faec, 32'hc290587a},
  {32'hc48b6c3a, 32'hc2ac02f9, 32'hc281352e},
  {32'h44a43786, 32'h433a51c5, 32'h43267d80},
  {32'hc48f9e6c, 32'h438b1bf9, 32'h4302422d},
  {32'h44ed980a, 32'h42fc91f2, 32'h435daaa1},
  {32'hc4ac25d6, 32'hc368833d, 32'hc34dd44c},
  {32'h44504bf6, 32'h4383debc, 32'hc341e967},
  {32'hc3257408, 32'hc3436370, 32'h43ba745d},
  {32'h44d09fba, 32'h4289ae4c, 32'hc2c04617},
  {32'hc4c489bc, 32'hc18670bc, 32'hc374eabf},
  {32'h43e4d1ba, 32'hc3dcd194, 32'hc3982868},
  {32'h426afe40, 32'hc0a326fc, 32'h41d404e3},
  {32'h44add3ed, 32'hc36777f2, 32'hc31e1d45},
  {32'hc5087d94, 32'hc388e47d, 32'hc0d233a6},
  {32'hc341cc28, 32'h43596e24, 32'hc3db8a60},
  {32'hc502b30b, 32'hc0b83fb0, 32'hc236d730},
  {32'h44d5772e, 32'h4344d5f1, 32'hc1133cd4},
  {32'hc4870400, 32'hc40d1ef6, 32'h433786c6},
  {32'h45141cec, 32'hc402ad53, 32'hc3280751},
  {32'hc3d279cc, 32'hc3602b89, 32'h43b57a0d},
  {32'h449ee122, 32'hc351e218, 32'hc3b14064},
  {32'hc4891c1e, 32'hc2a6ce2e, 32'hc2b4f8d9},
  {32'h4508da65, 32'hc39b297f, 32'hc3d674d5},
  {32'hc4780abd, 32'hc25e93d7, 32'h4384bcb5},
  {32'h439d317c, 32'hc3bacde8, 32'hc35f191f},
  {32'hc1c654c0, 32'hc306ef06, 32'h43bdd728},
  {32'h44a28132, 32'h42daa9c1, 32'hc33227f9},
  {32'hc4568182, 32'h4408981b, 32'hc1bb8709},
  {32'h44dbb8d8, 32'hc3c54a36, 32'hc343e7d1},
  {32'hc526b02a, 32'h4288d930, 32'hc148dd10},
  {32'h44eaaa55, 32'h42d94dc0, 32'h42ec7915},
  {32'hc4f71475, 32'h4395c50d, 32'h43d30093},
  {32'h450111d6, 32'h4315d8e5, 32'hc0ae2498},
  {32'hc4a88c3e, 32'hc2de2802, 32'h43beb646},
  {32'h44e74008, 32'h43020201, 32'h43055273},
  {32'hc50083ee, 32'h4305dc78, 32'h41a01629},
  {32'h44929f44, 32'h430d7d9e, 32'hc2985d8f},
  {32'hc4b67bcb, 32'hc0a6b828, 32'hc10e291c},
  {32'h45157d39, 32'hc14898cc, 32'hc3f2b9ea},
  {32'hc5121cbb, 32'h41f5268e, 32'hc3c3b144},
  {32'h451a6837, 32'h43be0d52, 32'hc0c8c298},
  {32'hc492d79d, 32'hc3bb24f0, 32'h438a3676},
  {32'h445c07aa, 32'h4343d3f6, 32'h43a28878},
  {32'hc34f000d, 32'h41f5dd62, 32'h4335174a},
  {32'h44723578, 32'h41b414e6, 32'h42e2eac3},
  {32'hc4db3fbe, 32'hc2585471, 32'hc18ac7e7},
  {32'h43784e3e, 32'hc36b2b04, 32'h420352e0},
  {32'hc37cc330, 32'h41902810, 32'h4308864a},
  {32'h449202dd, 32'hc0e23761, 32'h42cf48ca},
  {32'hc4e677b0, 32'hc309dcbe, 32'h422df3f3},
  {32'h42ea3d40, 32'hc348ea52, 32'h431b2016},
  {32'hc3b1ce80, 32'hc2eeb497, 32'h42e78e2e},
  {32'h44a2df22, 32'hc38a3cf8, 32'h431aca85},
  {32'hc2dfd200, 32'h409bf02e, 32'hc31186c7},
  {32'h4506fb81, 32'h4354b406, 32'hc321bfa8},
  {32'hc5004eb4, 32'h4426d0ad, 32'hc392582f},
  {32'h445b36c6, 32'hc3487e6d, 32'hc28c9e6b},
  {32'hc21a25c2, 32'h4126b003, 32'hc3afe7de},
  {32'h426488c0, 32'h4388607f, 32'hc3e53814},
  {32'hc46d2c28, 32'h43136806, 32'hc108d804},
  {32'h446a1462, 32'hc243c6a6, 32'hc3809ee2},
  {32'hc4f1910d, 32'h42ca4a1c, 32'hc351dc8f},
  {32'h44ae877a, 32'h42eb0f30, 32'h4323a664},
  {32'hc5105ec2, 32'h42c6e1f1, 32'h4318fa28},
  {32'h4488c2a4, 32'hc38e7541, 32'h42b90df7},
  {32'hc35e2883, 32'hc1f6177a, 32'h429551ae},
  {32'h44c4c2c0, 32'h43857f27, 32'hc1a202a8},
  {32'hc44fec81, 32'h40f96772, 32'hc2504b6e},
  {32'h43ed4e26, 32'hc22d742c, 32'hc21b5e35},
  {32'hc4908aee, 32'h42cbb1a6, 32'hc33399ba},
  {32'h44a520b0, 32'hc3ae7485, 32'h40d49ace},
  {32'hc4dad48a, 32'h41bd3937, 32'hc1e3d56e},
  {32'h44228be4, 32'hc2d77b4e, 32'h42b3f389},
  {32'hc4b1deff, 32'hc2a4c798, 32'hc316977c},
  {32'h43fd80ba, 32'hc22faeec, 32'h41e0fc06},
  {32'hc452feb6, 32'hc29edf12, 32'hc2a6d6a9},
  {32'h43970758, 32'hc30d65f1, 32'h43611ea7},
  {32'hc48af268, 32'h41f162d0, 32'hc3c920b2},
  {32'h43bb0640, 32'hc26a8260, 32'h4316760c},
  {32'hc41fc26b, 32'h42ca8603, 32'hc32cad04},
  {32'h44261a7c, 32'h418a7498, 32'hc397ab44},
  {32'hc4988ab5, 32'h42aae581, 32'h4309f96e},
  {32'h44bc2a2a, 32'h4326f288, 32'hc3d2b247},
  {32'hc4a9d01b, 32'hc201a358, 32'hc3b5eac3},
  {32'h449a8540, 32'hc31d5f99, 32'hc26a9503},
  {32'hc354529c, 32'hc353a45f, 32'h431e8990},
  {32'h44cdeda5, 32'h421766c4, 32'h4255084d},
  {32'hc4e8973e, 32'hc3724934, 32'hc2ebd5fe},
  {32'h4462e962, 32'h42b7374a, 32'h412c8b04},
  {32'hc4be7852, 32'hc34e257f, 32'h4302af1d},
  {32'h44aaaf7e, 32'h43c31ea2, 32'hc1a3f9ed},
  {32'hc4818910, 32'h42781fe2, 32'hc2b74c45},
  {32'h44c5e3ee, 32'hc3455d26, 32'hc280ee54},
  {32'hc4810be4, 32'h434eb461, 32'hc357aec0},
  {32'h44837701, 32'h4404d534, 32'h436e6c12},
  {32'h434f4080, 32'hc3c84b36, 32'hc2a9c173},
  {32'h44b563fe, 32'hc32c6ff9, 32'hc38047b7},
  {32'hc46e2952, 32'h43d920d2, 32'h42e41369},
  {32'h4420cf8e, 32'h42d950f2, 32'hc29627ad},
  {32'hc42db74d, 32'hc2966852, 32'h4345a909},
  {32'h44918ae4, 32'hc372201d, 32'h413937dc},
  {32'hc4f07264, 32'hc31498f9, 32'h4193fe78},
  {32'h44f39482, 32'hc380af4a, 32'h42bf94b2},
  {32'hc4ccc7ea, 32'hc3897ee3, 32'h43c43b8a},
  {32'h440b0b0c, 32'hc35dc4d8, 32'h431d3696},
  {32'hc3add486, 32'hc3b66849, 32'hc2a824d6},
  {32'h4354a050, 32'hc19de764, 32'hc2080631},
  {32'hc4f2d0a7, 32'hc30f62fb, 32'h42f97c3d},
  {32'h450eb0ae, 32'hc3183036, 32'h431c5311},
  {32'hc4ee1a26, 32'h44316bac, 32'hc374ef09},
  {32'h44bda141, 32'hc2760d4e, 32'h42856c33},
  {32'hc45a376d, 32'h429e9877, 32'hc3427d80},
  {32'h43c2104c, 32'hc32a7318, 32'hc393d8b3},
  {32'hc4aef0ba, 32'h43b2fa33, 32'h4381ce90},
  {32'h4502e58c, 32'h436e679b, 32'hc36f33a9},
  {32'hc4f60f56, 32'hc1cbe2d2, 32'h40ed0776},
  {32'h44b664c6, 32'hc1a4fa5a, 32'h43802c64},
  {32'hc4b289dd, 32'hc3e2658d, 32'hc334a592},
  {32'h4487811a, 32'hc30805ea, 32'h436b9f6b},
  {32'hc405b8f0, 32'hc2c06d81, 32'hc34d8c58},
  {32'h44966f8c, 32'h41eb570b, 32'h4305ce87},
  {32'hc43f29f2, 32'h42b88cb4, 32'h433bb2c0},
  {32'h448b9ff6, 32'h4252dc28, 32'h4398903d},
  {32'hc46f3acc, 32'hc2b8063f, 32'h431bf746},
  {32'h45032336, 32'h435bd96d, 32'hc3862d51},
  {32'hc4cf36cc, 32'h43ac362c, 32'h430049c0},
  {32'h444aadf5, 32'h418bd1b8, 32'hc3cb1179},
  {32'hc40b53a6, 32'h4222a182, 32'hc33d10be},
  {32'h45059f13, 32'hc3dd9d69, 32'h43ef5c2b},
  {32'hc4381d4a, 32'h439a19cf, 32'hc2b1ab7b},
  {32'h44998610, 32'h433446c2, 32'hc34d5867},
  {32'hc4fbe652, 32'hc37d0970, 32'h42d29cad},
  {32'h440677c6, 32'h4336bfcb, 32'h42a5223f},
  {32'hc4d8ced8, 32'h4185a2e8, 32'hc36146c7},
  {32'h42b40688, 32'hc206f003, 32'h40e1fe80},
  {32'hc3c4b0d8, 32'hc391528c, 32'hc1a45eca},
  {32'h44fb5efe, 32'hc2906599, 32'h43b8d77b},
  {32'hc502de66, 32'h41bcf81a, 32'hc33167ad},
  {32'h44f33321, 32'hc343ed6d, 32'hc262c0be},
  {32'hc4d61874, 32'h4288c3d4, 32'h418b2aff},
  {32'h449f4046, 32'hc2ea1772, 32'h43ad552f},
  {32'hc3106f91, 32'hc2c2631f, 32'hc409634a},
  {32'h4501b340, 32'h43e431da, 32'h43c5c71a},
  {32'hc50ac3f4, 32'h430005ae, 32'h42b0f8a3},
  {32'h44ec73fa, 32'hc2889a86, 32'hc3967aa0},
  {32'hc4b5328b, 32'hc2a63e7c, 32'h434e415d},
  {32'h44566110, 32'hc2be01e4, 32'h4278201c},
  {32'hc38d4b22, 32'h42b528a1, 32'hc377c337},
  {32'h44d1af38, 32'h43daf970, 32'hc31434ed},
  {32'hc4381fb7, 32'h427d4d5f, 32'h431b425c},
  {32'h428d2ef0, 32'h43cfda03, 32'hc3199268},
  {32'hc5168f21, 32'hc393ca59, 32'h434a0838},
  {32'h44d47b9b, 32'h43db5f82, 32'h422a8f6c},
  {32'hc4375714, 32'hc3c54141, 32'h430414ae},
  {32'h450ef4e3, 32'hc352053d, 32'h42a7a964},
  {32'hc40231e4, 32'hc31ea722, 32'h3ea7989c},
  {32'h44a79306, 32'hc2083226, 32'h4286c8d5},
  {32'hc4f87c00, 32'h4145a734, 32'hc2d3c7dc},
  {32'h44a9adb4, 32'h43c22037, 32'h42b65074},
  {32'hc48dde0d, 32'hc28e7765, 32'hc380db96},
  {32'h449d28e9, 32'h436a1f0e, 32'hc1c45922},
  {32'h41c8cfc0, 32'h42da4878, 32'h4294d8df},
  {32'h4508305a, 32'hc3319678, 32'hc32a6f23},
  {32'hc4a930a8, 32'h436ed667, 32'hc387ce6b},
  {32'h443d7510, 32'h438a292a, 32'h4368ab71},
  {32'hc40dc578, 32'h42976c67, 32'hc306c3b1},
  {32'h4406dca7, 32'hc37f05ed, 32'hc2c0d565},
  {32'hc4d54698, 32'h4120763f, 32'h42e7591d},
  {32'h43acbe69, 32'h42c596ce, 32'hc2fc4474},
  {32'hc485b43c, 32'hc37847c8, 32'h416531aa},
  {32'hc2348e28, 32'hc30ee7a9, 32'hc3c37ff4},
  {32'hc4550ed8, 32'hc2c62507, 32'h42c18d99},
  {32'h43b5f506, 32'h42bd5dec, 32'h4288edde},
  {32'hc3d1c310, 32'hc36d1d0c, 32'hc254e052},
  {32'h449ec4b2, 32'hc013d334, 32'h42b338d6},
  {32'hc4c8d2c9, 32'hc30854c1, 32'hc39401ec},
  {32'h44f5cc8a, 32'hc2b6f0c6, 32'h43441e81},
  {32'hc43cc4bc, 32'hc329aa69, 32'h43122444},
  {32'h44af6524, 32'h42cef0f7, 32'hc339719f},
  {32'hc4748b8d, 32'h42bd1f54, 32'h43799c27},
  {32'h44d316c1, 32'h43961d2a, 32'hc2bce134},
  {32'hc462931e, 32'hc26e14a1, 32'h433394b6},
  {32'h4518e93f, 32'hc33c183c, 32'h43c5f7e7},
  {32'hc49e9318, 32'hc15f98db, 32'hc3ac71f1},
  {32'h450fddf7, 32'hc2fb93e2, 32'hc1e6bd9c},
  {32'hc4128e94, 32'h40a7d174, 32'h436f062c},
  {32'h43f765c8, 32'h4222e71a, 32'hc0dc3bbe},
  {32'hc2ebd6e0, 32'h42d32718, 32'hc39b4270},
  {32'h44a94a7e, 32'hc230bac8, 32'h43bc44cf},
  {32'hc4992cb2, 32'h421caba3, 32'h4246de13},
  {32'h4435f722, 32'h42f64ae3, 32'hc2faab7c},
  {32'hc47fef7a, 32'hc0afdfe6, 32'hc379c99c},
  {32'h44bd7646, 32'hc3a51813, 32'hc2dd6a2d},
  {32'hc2bb9960, 32'h43425294, 32'hc376adaa},
  {32'h44373de6, 32'h4303a946, 32'hc3a36214},
  {32'hc4ff5e37, 32'hc2235bd3, 32'hc30c6379},
  {32'h43400488, 32'hc32bf17d, 32'h4286d629},
  {32'hc505b98e, 32'hc21a0e9c, 32'h42c46b0b},
  {32'h44e184f4, 32'h438c4ba1, 32'h4389d340},
  {32'hc218c147, 32'hc3644eec, 32'hc37814b2},
  {32'h451a11af, 32'h42de2be6, 32'hc2d95283},
  {32'hc4ab32e7, 32'hc235307a, 32'hc2f9a49d},
  {32'h4429fa8c, 32'hc40b5e97, 32'hc1646f78},
  {32'hc462b3ee, 32'hc36bf24a, 32'hc380c18c},
  {32'h450a945a, 32'h43801910, 32'hc3f97014},
  {32'hc4a55a22, 32'h43247d2a, 32'h42fc625e},
  {32'h4494c91c, 32'hc34f57e2, 32'hbe8273c0},
  {32'hc516e3d3, 32'hc37e31fc, 32'hc2f5abd7},
  {32'h44147070, 32'h42ec7c03, 32'h428cfea7},
  {32'hc4030e17, 32'hc281b5e6, 32'h4400c44e},
  {32'h4518cf5f, 32'h43484643, 32'hc38e2b4b},
  {32'hc441cfa6, 32'hc183a485, 32'h4401994a},
  {32'h44eeb229, 32'hc3006c99, 32'hc2410a7f},
  {32'hc483a53f, 32'hc2aa0c47, 32'hc27f11ac},
  {32'h450cf500, 32'h43c5bdb2, 32'h42e3bd26},
  {32'hc3e54ba1, 32'h4297dfc6, 32'h4386dd97},
  {32'h450e4784, 32'hc34adada, 32'hc2e2f0c2},
  {32'hc48f6cfe, 32'h43ac1cdc, 32'h4353ed54},
  {32'h43d748fa, 32'h43488389, 32'hc23d4f00},
  {32'hc418e160, 32'h4344dc91, 32'hc34078f0},
  {32'h44bd9041, 32'hc2f4d498, 32'h437b4f0f},
  {32'hc4097068, 32'h428a6060, 32'h423df827},
  {32'h43d1ad48, 32'h41fbc2c9, 32'h420fdc0b},
  {32'hc4a8ebce, 32'h44030823, 32'hc2abb00f},
  {32'h43e2e02c, 32'h4372ea4f, 32'hc35a16ec},
  {32'hc5039bab, 32'h43b21ea2, 32'h425c9eec},
  {32'h44d8d90a, 32'h440bf5bd, 32'h439b068f},
  {32'hc3dc0084, 32'h428991f0, 32'hc2972d27},
  {32'h4399240c, 32'h42f65f86, 32'h4216110c},
  {32'h4347e860, 32'hc322f84b, 32'h4231878c},
  {32'h44a5fe42, 32'h43bb981d, 32'h42c02433},
  {32'hc5069ae9, 32'hc368d36a, 32'h435a1bb0},
  {32'h4497b61d, 32'hc136b466, 32'h430c8402},
  {32'hc4403ef4, 32'hc3f45923, 32'h42e0e6ac},
  {32'h4440591b, 32'hc1f61259, 32'h43ac3383},
  {32'hc510c82a, 32'hc30e80cd, 32'h43b0c19e},
  {32'h4461d1aa, 32'hc2b7de8a, 32'hc395b868},
  {32'hc46f1bfb, 32'h435952ed, 32'hc2568b95},
  {32'h44e7b2a8, 32'hc319155f, 32'hc310f9c2},
  {32'hc4e971c4, 32'hc3504975, 32'h42feff13},
  {32'h450d8f5f, 32'h426c367b, 32'hc352246f},
  {32'hc5046a86, 32'hc3330f2d, 32'hc3c8e0e1},
  {32'h44832b46, 32'hc1f42125, 32'hc3bf55b7},
  {32'hc50b33e6, 32'h40ea42cc, 32'h42296d4e},
  {32'h450275f0, 32'h42cbdf44, 32'hc394f197},
  {32'h436424cd, 32'h4181e3a2, 32'h42aced72},
  {32'h44ca7282, 32'h42c56745, 32'hc2e1d61d},
  {32'hc4ad9186, 32'hc3425fcd, 32'hc40fbf05},
  {32'h440d20d3, 32'h43a05f66, 32'hc3c8aa6b},
  {32'hc504b14e, 32'h42a31aa4, 32'hc2f43f3f},
  {32'h44a16d39, 32'hc3518865, 32'h434cb1c7},
  {32'hc4e5ac64, 32'hc3c9067e, 32'h430211b1},
  {32'h45027381, 32'hc2b735a2, 32'hc3d6cf32},
  {32'hc4ce2e6a, 32'hc37d284c, 32'h432e7c0b},
  {32'h440f4d1a, 32'hc175dd61, 32'hc2551821},
  {32'hc4947c26, 32'h43007bb6, 32'h4319cd34},
  {32'h432673d0, 32'h4308fd58, 32'h43b3e79f},
  {32'hc499c97d, 32'h42ceb889, 32'h40894da9},
  {32'h451f81cc, 32'hc34399c2, 32'hc31f5aa7},
  {32'hc3d99885, 32'hc1223885, 32'hc2e3468c},
  {32'h44ebf654, 32'h3f0dbbaa, 32'hc3b7e36a},
  {32'hc32dbd50, 32'h43984442, 32'hc2bb1820},
  {32'h450b371e, 32'hc06737c9, 32'h43a0f861},
  {32'hc396017c, 32'hc31108a6, 32'h431224ed},
  {32'h442ae6a0, 32'hc344c6c9, 32'h4275fa0b},
  {32'hc36b6280, 32'hc2b07e6e, 32'hc2ba5fda},
  {32'h44b0c092, 32'h43dafa0b, 32'h431760da},
  {32'hc3b7470c, 32'h41ebfb83, 32'h43a0654c},
  {32'h43eb2c1c, 32'h42e1ee64, 32'hbfe8b540},
  {32'hc4e25f7a, 32'h40547d32, 32'h43a9a7e1},
  {32'h45130c92, 32'hc1b0287f, 32'hc32c63a3},
  {32'hc50c3204, 32'hc364cb43, 32'h426bf5b5},
  {32'h4494fa58, 32'h42f638f8, 32'h42d4bc93},
  {32'h42e36b60, 32'hc402bc21, 32'hc385e249},
  {32'h4386e388, 32'h42620da7, 32'h42a950db},
  {32'hc49388d6, 32'hc2630ecb, 32'hc34d4405},
  {32'h44ec38a6, 32'hc2077310, 32'h4279e79b},
  {32'h43c5a019, 32'h43366a7b, 32'hc35fa37f},
  {32'h44b0fb4c, 32'h436b4318, 32'hc384f457},
  {32'hc462250c, 32'hc2dba872, 32'h43b1b672},
  {32'hc3027af8, 32'hc3534bfc, 32'h43272e9a},
  {32'hc3b40360, 32'h42b3b7b9, 32'hc36b61ec},
  {32'h450fa060, 32'h43c3b02d, 32'h4372cdd1},
  {32'hc5171c1d, 32'hc2f2effb, 32'h43fa21bf},
  {32'h444e9368, 32'h42445202, 32'hc30a3b3e},
  {32'hc2161048, 32'h42b81ef6, 32'h433ef075},
  {32'h450e1f64, 32'hc29a4c4c, 32'h42ab3748},
  {32'hc47d5318, 32'h422c94ea, 32'h43237af7},
  {32'h451616d2, 32'hc2b4dc33, 32'h4306c582},
  {32'hc4810b27, 32'h41535a0f, 32'h4280fec9},
  {32'h44935ce0, 32'h41e24b22, 32'h41a5d3fa},
  {32'hc50ced48, 32'h4331522d, 32'h42352b59},
  {32'h4407f132, 32'h441bb387, 32'h42fd39f1},
  {32'hc508a795, 32'hc24bdd02, 32'hc2a2aa88},
  {32'h44164d85, 32'hc3a2e2c3, 32'h42fa5e77},
  {32'hc39de009, 32'h42a533c8, 32'h418db494},
  {32'h45026887, 32'h43b5eea2, 32'h43249f8d},
  {32'hc3bec36b, 32'hc2b88897, 32'h438c6607},
  {32'h45108393, 32'hc217ce91, 32'hc3ad9856},
  {32'hc4f51068, 32'h43dc852b, 32'hc24ab0ed},
  {32'h44ce5051, 32'hc2a8b42c, 32'hc2a2fb1c},
  {32'hc428f13d, 32'hc32f6554, 32'hc1c96ed0},
  {32'h447ac858, 32'h432f66f0, 32'hc2c38fdc},
  {32'hc4d10a4a, 32'hc237e51d, 32'h42fe054a},
  {32'h43febf98, 32'h43b3d301, 32'h429b4e60},
  {32'hc2e22ab8, 32'h41cff5ad, 32'h43a1870f},
  {32'h44c157b4, 32'hc309593d, 32'hc354e7a1},
  {32'hc4357c00, 32'h4286e329, 32'hc238de9e},
  {32'h436b0b28, 32'h43058d89, 32'hc2033e8e},
  {32'hc4b69a61, 32'hc332b958, 32'hc31a18a2},
  {32'h44e28194, 32'h4384b7d2, 32'hc397238f},
  {32'hc49626de, 32'h43825ff2, 32'h43707468},
  {32'h4510aaac, 32'h43a75659, 32'h43dba668},
  {32'hc4d744dd, 32'h41a825c1, 32'h4212b75a},
  {32'h44fd705f, 32'hc3261010, 32'hc2296171},
  {32'hc4dd49c5, 32'h42b7e7d4, 32'h42b56eb5},
  {32'h439e0230, 32'h429b82c7, 32'hc3629051},
  {32'hc415bb74, 32'h433220b6, 32'h43184bda},
  {32'h43e27ac0, 32'hc3211a6f, 32'h41ab2ec4},
  {32'hc4c7c156, 32'hc3eb6628, 32'h433d8bf9},
  {32'h4494c785, 32'h42fadb71, 32'h431e51df},
  {32'hc4ee3f2c, 32'hc3be3d85, 32'h42a1089b},
  {32'h44b3bcac, 32'h43440b10, 32'hc36ac7db},
  {32'h4281f7f4, 32'hc2a2e93d, 32'h433c061c},
  {32'h44aa110f, 32'hc3bd6062, 32'h43a1fd12},
  {32'hc420e0d2, 32'hc18573c5, 32'h43a3139c},
  {32'h44aa3e87, 32'hc2d39b12, 32'hc31d3005},
  {32'hc2f98d1e, 32'h4329d77e, 32'h43bc577a},
  {32'h44f4c69c, 32'hc26c6f2a, 32'hc33a82e3},
  {32'hc4d3f010, 32'hc3491256, 32'hc29e59e3},
  {32'h445d7952, 32'h4334f80e, 32'hc1c63d7e},
  {32'hc51b4dc3, 32'h43a56060, 32'hc3033713},
  {32'h44474dce, 32'hc3930419, 32'hc37a286a},
  {32'hc4e38437, 32'h42f96f3e, 32'h40a5e51b},
  {32'h450ea0fc, 32'hc30c7cbc, 32'hc363216f},
  {32'h44a2c3b6, 32'hc2837b63, 32'h43041a31},
  {32'hc4b88968, 32'hc2de9938, 32'hc3237689},
  {32'h43098320, 32'hc40b83d8, 32'h42279b04},
  {32'hc4940efe, 32'hc30526ac, 32'hc37343d6},
  {32'h44b32b97, 32'hc295d9db, 32'h43108c15},
  {32'h41817500, 32'hc2bf269a, 32'h4290b486},
  {32'hc2cf8160, 32'hc27073d3, 32'hc35a85b9},
  {32'hc49fcd44, 32'hbf9f5d60, 32'hc22d8568},
  {32'h44f9aabd, 32'h436ad613, 32'h43592cd1},
  {32'hc4a588da, 32'h4391068e, 32'hc21f21b7},
  {32'h44ffcdf2, 32'h43a91176, 32'hc38e6686},
  {32'hc498e0a2, 32'hc34eb5fb, 32'h43286e6e},
  {32'h437fd2b0, 32'h435161c2, 32'hc3fdeb84},
  {32'hc4ced3e7, 32'hc2c3a9d6, 32'h42df5994},
  {32'h439c6e88, 32'hc382a910, 32'hc13c272a},
  {32'hc40c55ee, 32'hc267cded, 32'h4402ae64},
  {32'h44df4659, 32'h435956c6, 32'hc3af5b3d},
  {32'hc4964ba0, 32'h4249d44d, 32'h41caa449},
  {32'hc2f83610, 32'h43a0b9f4, 32'h42aa8e09},
  {32'hc4e7a9d9, 32'hc2e6aa3f, 32'hc38e99b0},
  {32'h447cccb8, 32'h43354954, 32'h424c1896},
  {32'hc40d9924, 32'hc3134a38, 32'h43d60111},
  {32'h44976b4f, 32'h42a6bf50, 32'hc26794bc},
  {32'hc4ca7168, 32'h43833d40, 32'hc3193e3f},
  {32'h44b8dd02, 32'h4394022f, 32'hc2a06d70},
  {32'hc4f7ffcb, 32'h4251174f, 32'hc2c7da27},
  {32'h44eb68ff, 32'h429ec262, 32'h422f3533},
  {32'hc4fe4c6a, 32'hc348d449, 32'hc32545c8},
  {32'h44958346, 32'hc35e27ce, 32'hc307a990},
  {32'hc4d10bea, 32'hc336e193, 32'h412b53e8},
  {32'h44c7615f, 32'hc2251838, 32'h433ca7f3},
  {32'hc501d6b7, 32'hc331d026, 32'h43912494},
  {32'h44cbee4a, 32'h42b39303, 32'hc2c8fff5},
  {32'hc40a5a36, 32'hc365122c, 32'hc3bc2a5d},
  {32'h446b4a41, 32'hc14829d0, 32'hc32b5e34},
  {32'hc186f500, 32'hc2436c90, 32'hc281b8c7},
  {32'h4365fa16, 32'hc3a9a43d, 32'hc3f2401d},
  {32'hc4db5e3f, 32'h43a2ed96, 32'hc31bccf0},
  {32'h44c1b30d, 32'hc284dba3, 32'hc35914dc},
  {32'hc40ba5bc, 32'hc182c3b0, 32'h439b627d},
  {32'h4383e560, 32'hc348517f, 32'hc389831f},
  {32'hc4c2420f, 32'h42d41398, 32'hc28c4d65},
  {32'h44f02d3f, 32'hc381fa4d, 32'h437b08c7},
  {32'hc3b7b136, 32'hc34c594a, 32'h42948469},
  {32'h45104fe5, 32'hc311e0bc, 32'h43fde14c},
  {32'h436d668a, 32'hc37f011b, 32'hc35f016d},
  {32'h451cdf1f, 32'h4135481a, 32'h4317a823},
  {32'hc4ddc439, 32'hc2821f95, 32'hc3ae899d},
  {32'h4500cc7e, 32'h44243921, 32'hc3b185ab},
  {32'hc41d57c0, 32'h42b077ad, 32'hc3672f1e},
  {32'h451358ca, 32'h430a0da5, 32'h43860fd3},
  {32'hc4198a0e, 32'hc3e1807f, 32'h4346a908},
  {32'h432b74f0, 32'h431f45d7, 32'h432da8f3},
  {32'hc4f175ed, 32'hc24e86a3, 32'h41990756},
  {32'h44f82908, 32'h423ff33d, 32'hc3e70439},
  {32'hc4bcf017, 32'hc26cf188, 32'hc2a3a5a9},
  {32'h4501e8d2, 32'hc2b60aa3, 32'h42130530},
  {32'hc454eb46, 32'h4256151e, 32'h4313c6f3},
  {32'h4398b753, 32'hc376bf88, 32'h43486831},
  {32'hc3e3e1b1, 32'hc3502ba7, 32'h43ca62d1},
  {32'h4356233a, 32'hc2ae9aa7, 32'h43a0ebc1},
  {32'hc4babea9, 32'hc1b24557, 32'hc3bbb5d9},
  {32'h44944e5e, 32'h42a4998c, 32'h40941b34},
  {32'hc4a409ec, 32'h4349d602, 32'h42c6f557},
  {32'h4512809a, 32'hc31211cc, 32'h42fc08ed},
  {32'hc3aa9e80, 32'hc4206bf0, 32'h4392fa75},
  {32'h44ec7024, 32'h43ad2ba2, 32'h4381e60b},
  {32'hc4fa5f6a, 32'hc36755e4, 32'hc3742224},
  {32'h44fe59d0, 32'h43eb979c, 32'h42c4bc08},
  {32'hc4ccf0ce, 32'h4354a75f, 32'hc071d610},
  {32'h4382f3a2, 32'hc362b172, 32'h4153be4c},
  {32'hc4f53e49, 32'hc3185eb5, 32'h431963d6},
  {32'h44d66373, 32'h43155ee2, 32'hc3724322},
  {32'hc43da91b, 32'hc26c4a9a, 32'h433908a4},
  {32'hc356535a, 32'hc28a376d, 32'hc210eca8},
  {32'hc4d8d99a, 32'hc3890a32, 32'hc1150fff},
  {32'h442aa41e, 32'hc39cac31, 32'hc40c06e1},
  {32'hc4ecd080, 32'hc2ea6d1f, 32'h42e53ad0},
  {32'h44b4dad4, 32'h43ac5fe8, 32'hc3c9fd9a},
  {32'hc4ad4c4b, 32'hc3738615, 32'h4275d484},
  {32'h449037a6, 32'hc3bd74ba, 32'h432a4568},
  {32'hc30b4268, 32'h42d2e07e, 32'h4348999a},
  {32'h44b21dd3, 32'h429f4b90, 32'h4181b82d},
  {32'hc503b9c0, 32'hc2fcff1b, 32'h4315b8f4},
  {32'h42536120, 32'h429c59db, 32'h43f2d12b},
  {32'hc4b8cef0, 32'h43a7989d, 32'hc330af8d},
  {32'h44b39bf0, 32'hc2dc6b87, 32'hc28419ee},
  {32'hc48ebbc4, 32'h4252a66f, 32'hc39b81b6},
  {32'h448067e6, 32'h42d95cb8, 32'hc281cae1},
  {32'hc496fa72, 32'hc3a010f8, 32'hc3b241d5},
  {32'h45033af2, 32'h42957506, 32'hc3c9c247},
  {32'h4158c630, 32'hc39dc712, 32'h41fb1419},
  {32'h448e3b47, 32'hc3a0c7ad, 32'hc2f83ed9},
  {32'hc4a14466, 32'h423beef2, 32'hc32d3522},
  {32'h44bc0226, 32'h42eb90e5, 32'hc32f48e9},
  {32'hc1e1e800, 32'hc2cb978f, 32'h41b95f22},
  {32'h44c23277, 32'hc286f491, 32'hc3390173},
  {32'hc326ccb7, 32'h440e113a, 32'hc2ba88a6},
  {32'h4424435e, 32'h42b2287b, 32'h4309f9ca},
  {32'hc494779d, 32'h42d0c454, 32'hc247b428},
  {32'h44706cc4, 32'h43318e0a, 32'h43dffd53},
  {32'hc5087cf8, 32'hc36ec666, 32'hc335bb3c},
  {32'h448f0dec, 32'h433b82ae, 32'h436b997a},
  {32'hc3760a12, 32'h43462b7b, 32'hc241b4ab},
  {32'h44b76916, 32'h440568d3, 32'hc1c849e4},
  {32'hc5197796, 32'h418ebb0e, 32'hc2d5ccd0},
  {32'h44de53e0, 32'hc3862b38, 32'hc202de97},
  {32'hc483f3a0, 32'h41a425da, 32'h42945881},
  {32'h44bc5530, 32'hc31c02f9, 32'h423b1558},
  {32'hc48705a1, 32'hc2597c53, 32'hc2ddfa87},
  {32'h44c3379f, 32'hc1cb3905, 32'h4080f068},
  {32'hc4f6c90d, 32'h4382b0bf, 32'h437842d4},
  {32'h4430e6bb, 32'h42e4ea14, 32'h440000bb},
  {32'hc451d030, 32'hc2fd7983, 32'h43853b57},
  {32'h43aa480a, 32'hc3c2a368, 32'hc2fd2395},
  {32'hc49194e6, 32'h42a215ae, 32'h42b87a81},
  {32'h44eefdd6, 32'h431d8602, 32'hc3915746},
  {32'hc3a1b3ba, 32'h43d89f1a, 32'h41b5ff4a},
  {32'h440cb650, 32'h426afb9d, 32'h435a3aa9},
  {32'hc30e8a01, 32'h41448ae0, 32'h42cfbe10},
  {32'h44c6b03f, 32'h43e3c206, 32'hc3c0a92f},
  {32'hc3ee78b8, 32'h43bb4c0a, 32'h42fe6548},
  {32'h4423a4c0, 32'h431eb24c, 32'hc20588fb},
  {32'hc4e86a18, 32'h43b4822c, 32'h41b1208e},
  {32'h43da90c8, 32'hc3622c39, 32'h43203641},
  {32'hc3f64b78, 32'h4310c13c, 32'hc1a6029d},
  {32'h449dc089, 32'hc2a956bd, 32'hc35ae681},
  {32'hc4430a74, 32'hc18e1062, 32'h433e00eb},
  {32'h44acbc1e, 32'hc203328c, 32'h432d766b},
  {32'hc4f0be84, 32'hc4085ba2, 32'h4407ff70},
  {32'hc304ff44, 32'h438d0d27, 32'hc215ee31},
  {32'hc512d812, 32'hc1b14539, 32'hc2d02a02},
  {32'h4481332e, 32'h4428c8a9, 32'hc018aace},
  {32'hc463bdb7, 32'h42763444, 32'h428304de},
  {32'hc3416d70, 32'h4393d6cc, 32'h42d220d4},
  {32'hc46f63cc, 32'hc33d4d07, 32'hc3375884},
  {32'h45018d8c, 32'h420cbac5, 32'hc2da1bc4},
  {32'hc49a1fe1, 32'h42467686, 32'hc292b782},
  {32'h44a1e652, 32'h426cf432, 32'h43781c42},
  {32'hc50ce712, 32'hc2ab57b0, 32'h42a08c4c},
  {32'h44af5f5a, 32'hc08fe4f7, 32'hc313c980},
  {32'hc4a0cd4a, 32'h43185d6a, 32'h4306123e},
  {32'h4502ca4d, 32'hc21939e4, 32'hc3a1c559},
  {32'hc11f6c00, 32'h43e3ca59, 32'hc2d9e9fe},
  {32'h445f7f7a, 32'hc3408937, 32'h42c9e361},
  {32'hc29ecf40, 32'h43445373, 32'hc2402766},
  {32'h44684595, 32'h433d61cd, 32'h43d70c1f},
  {32'hc4fe5f84, 32'hc25756a9, 32'h4325f7f1},
  {32'h44ca0a2b, 32'h43691c8b, 32'h438ff9f4},
  {32'hc45bab62, 32'h4218d005, 32'h42623c73},
  {32'h44e890c5, 32'h4163abd5, 32'hc2fef5f4},
  {32'hc504e85d, 32'h43bbd3f4, 32'h43090819},
  {32'h4483c2f0, 32'hc2a7351e, 32'hc2d244f9},
  {32'hc4b6094b, 32'hc330440d, 32'hc241decf},
  {32'h43a0638e, 32'h42f64597, 32'hc31d0c77},
  {32'hc45129cc, 32'h43398660, 32'hc330f4d6},
  {32'h44e915b4, 32'h4055b7f7, 32'h41134379},
  {32'hc503d3cf, 32'hc341d431, 32'hc421c17f},
  {32'h448b93ac, 32'h42897f85, 32'h42ecfab4},
  {32'hc4d893bb, 32'h43ede692, 32'h43801768},
  {32'h44afc1da, 32'hc2b6e756, 32'h438e3531},
  {32'hc38956e4, 32'h42741434, 32'h43b739f3},
  {32'h44e67e87, 32'hc3889fe5, 32'hc24c1651},
  {32'hc42ffa11, 32'hc36352be, 32'hc3371116},
  {32'h43b1ff08, 32'h3fc30d60, 32'hc38c8e50},
  {32'hc4c6f0f1, 32'hc35b0719, 32'hc310c8fc},
  {32'h44f8dadb, 32'h441aecaa, 32'hc12f57bc},
  {32'hc4409e8c, 32'h437e7a9e, 32'hc3208db7},
  {32'h4482c7ac, 32'h4383f166, 32'hc38aa667},
  {32'hc465bb58, 32'h434e72c2, 32'h41cb649e},
  {32'h44f58b39, 32'h42aa27f2, 32'hc2cfc2e4},
  {32'hc4f52622, 32'hc2ce07ea, 32'h43908684},
  {32'h44fb4692, 32'hc0f85b2c, 32'hc2e100c4},
  {32'hc4ed1ab2, 32'h439ec587, 32'hc35f45f5},
  {32'h44aecead, 32'h43609fde, 32'h432f4776},
  {32'hc40790da, 32'h42200295, 32'h44184d59},
  {32'h438f1250, 32'h4210f532, 32'hc3b00eb6},
  {32'hc4a559a6, 32'hc37bbdae, 32'hc302e64d},
  {32'h450a3a03, 32'h4197b11e, 32'h426ed27e},
  {32'hc3cdb68c, 32'hc2e769db, 32'hc2e52a3c},
  {32'h443c9f41, 32'hc392800e, 32'hc33e76da},
  {32'hc503e0a8, 32'hc39fe96a, 32'hc38698a5},
  {32'h44eb3044, 32'hc0c43477, 32'h41341b20},
  {32'hc4d55edc, 32'h43afb2dd, 32'h433efcf8},
  {32'h44845066, 32'h421d931c, 32'hc315e517},
  {32'hc3eb49e8, 32'hc2bb7578, 32'hc367a532},
  {32'h44b6065e, 32'hc19f375d, 32'h414685aa},
  {32'hc4318d4a, 32'h42dd5d5b, 32'hc3b0e82a},
  {32'h4495bfd4, 32'hc2a03fbd, 32'h43643f8d},
  {32'hc4825d48, 32'hc30b38ac, 32'h428717d3},
  {32'h44c00ff4, 32'h4317f018, 32'h4330a3de},
  {32'hc46bc598, 32'h43b33dea, 32'h42fdeaec},
  {32'h44bf1875, 32'h438fdd26, 32'h435e2347},
  {32'hc4263032, 32'h432acb7f, 32'h42c284dd},
  {32'h449bf7e6, 32'h42d036c8, 32'hc1c57c84},
  {32'hc41002c4, 32'h4380cf84, 32'h43156bc6},
  {32'h442bd3cc, 32'hc237713a, 32'h42f3dc56},
  {32'hc2fac5a4, 32'h4275812e, 32'h436f2be4},
  {32'h44127d8c, 32'h43c38e5b, 32'hc3278344},
  {32'hc50ee5cb, 32'hc3c0c170, 32'h437cb95e},
  {32'h448c4d65, 32'h41cfe3a2, 32'h43cfe57b},
  {32'hc48177d5, 32'hc37b07f4, 32'h42111311},
  {32'h4377e280, 32'hc3d38a52, 32'h430c8fa6},
  {32'hc473921c, 32'h431fb63a, 32'h440f4658},
  {32'h4518efb2, 32'hc2c4bd35, 32'hc37e6314},
  {32'hc4860669, 32'hc262db68, 32'hc3f58326},
  {32'h44a15d58, 32'hc30ba0d3, 32'hc21d2708},
  {32'hc4f0c549, 32'h4340fce4, 32'hc33a900d},
  {32'h4504275f, 32'hc39c370d, 32'h43c2b6a3},
  {32'hc5050b26, 32'h42dffa73, 32'hc2b0fbf3},
  {32'h4501e0eb, 32'hc317304a, 32'hc2d8d191},
  {32'hc4914cb2, 32'hc17ea164, 32'h431a00d2},
  {32'h442f098f, 32'h4325be5f, 32'h432a25c4},
  {32'hc47abc83, 32'h43954ced, 32'hc3f80c88},
  {32'h44920132, 32'h4341aab3, 32'h43945890},
  {32'hc4f3b9d4, 32'hc2ca8998, 32'hc2f1a30a},
  {32'h4483a1c1, 32'hc314c5b1, 32'hc3044e06},
  {32'hc49b33f5, 32'hc29d47b5, 32'hc3a9a00b},
  {32'h44ca2ae5, 32'hc34880d7, 32'h42444dfa},
  {32'hc4be8ad9, 32'h435d993e, 32'h43843d9a},
  {32'h43e2f213, 32'hc29dda82, 32'h42e079fe},
  {32'hc436acf0, 32'h433d27a7, 32'h43700c60},
  {32'h42957f87, 32'h405e180f, 32'hc306f95a},
  {32'hc409cac0, 32'h4397808a, 32'hc2969c23},
  {32'h43fd2074, 32'hc2cf81de, 32'hc2d313cb},
  {32'hc4da9af9, 32'hc30b7336, 32'hc1a4a8f0},
  {32'h44adfd4a, 32'hc3f26189, 32'h4400b770},
  {32'hc4b300dd, 32'h420e03ef, 32'h433fa848},
  {32'h441d7c5c, 32'hc307d94e, 32'h437c90ac},
  {32'hc49a670e, 32'hc27da14e, 32'hc327a3a2},
  {32'h436f88c0, 32'hc284b20e, 32'h43a3efbf},
  {32'hc4a94081, 32'hc1820777, 32'h4310a87a},
  {32'h44be6fd2, 32'hc395c945, 32'h4360e940},
  {32'hc3e75b38, 32'hc2f5c993, 32'h42a1d5a4},
  {32'h450ceeb1, 32'h4238167f, 32'hc361d04b},
  {32'hc4e603ba, 32'hc3362128, 32'hc20f947a},
  {32'h44e1bc66, 32'h43babbb5, 32'hc39211bc},
  {32'hc4897079, 32'hc0ef7b76, 32'h442bb204},
  {32'h4504bf17, 32'hc28250b1, 32'hc3353aae},
  {32'hc4fe13f3, 32'hc29bd6e5, 32'h427505f4},
  {32'h44c18a1b, 32'hc25d892d, 32'hc382c4cb},
  {32'hc33dd3c2, 32'hc2494399, 32'h409a66c9},
  {32'h449ef171, 32'hc1a0f06e, 32'h41fa880f},
  {32'hc5027c6f, 32'h4303be95, 32'h44067d50},
  {32'h44a551a7, 32'h424eedb2, 32'h42458b88},
  {32'hc49f0952, 32'hc2e5446e, 32'h428d58e2},
  {32'h435154e4, 32'h42f31ec8, 32'hc34901b3},
  {32'hc4ccaaa1, 32'h43600022, 32'h4355610a},
  {32'h449e4bcb, 32'h4327eea0, 32'hc350e632},
  {32'hc4842c37, 32'h42334b23, 32'hc45f727b},
  {32'h449be5f0, 32'hc29136d6, 32'h4232a92b},
  {32'hc4fa2e68, 32'h42dda2ac, 32'h43807a0e},
  {32'h44c2eb98, 32'h3f90a4f8, 32'h42a63da0},
  {32'hc4afd262, 32'h42b35d25, 32'h4395a49e},
  {32'h448b2e24, 32'hc39bb501, 32'hc3681f09},
  {32'hc4e76f9e, 32'hc38b999a, 32'hc417adc9},
  {32'h44552f8e, 32'h43e08d11, 32'hc1ed6f55},
  {32'hc4e1a0ab, 32'hc2c6a53a, 32'hc2634736},
  {32'h44d9260c, 32'h4290490c, 32'hc3e74bd9},
  {32'hc3851dcc, 32'hc3be8fe2, 32'h432de09c},
  {32'h450cd1ea, 32'hc1f46dd2, 32'h4343d7d3},
  {32'hc5242f29, 32'h42dcfaea, 32'hc24a07b6},
  {32'h44a8bb02, 32'h41ab84c9, 32'h430d6446},
  {32'hc4829ec4, 32'hc2890350, 32'h435e28f6},
  {32'h45187495, 32'h4307f464, 32'h420b53c5},
  {32'hc4f26b52, 32'hc2d68c2b, 32'hc2c21835},
  {32'h4487b110, 32'h436f450d, 32'h4016342c},
  {32'hc4ad8c98, 32'h43e0bd40, 32'hc22041e1},
  {32'h447e3dec, 32'hc3d50e60, 32'h43275300},
  {32'hc30a34e0, 32'h425183d6, 32'hc32cd0cd},
  {32'h45108574, 32'hc3137065, 32'hc31936ac},
  {32'hc5008593, 32'hc311569b, 32'h41d72dc0},
  {32'h45090ff0, 32'hc30a5266, 32'h430cf401},
  {32'hc49ed957, 32'h43bbdebe, 32'hc3134125},
  {32'h43a6a7fd, 32'hc402f6d5, 32'hc3063053},
  {32'hc49cb052, 32'hc32b322f, 32'h43091da6},
  {32'h42fc8808, 32'h41bc73b0, 32'h4225889c},
  {32'hc50c91ee, 32'hc13957f7, 32'hc3b150b0},
  {32'h44cbd809, 32'h4401d146, 32'h43cedbec},
  {32'hc3a3c6d5, 32'h41b47463, 32'hc2c2ed30},
  {32'h44746384, 32'hc18fd050, 32'h42cf8b1d},
  {32'hc338f13b, 32'h43ad7d23, 32'hc1821b33},
  {32'h448f032d, 32'hc2b9c930, 32'h42b65707},
  {32'hc4726e8c, 32'h42812991, 32'h428be356},
  {32'h45012101, 32'h422391bb, 32'h432d87af},
  {32'hc4cf852e, 32'hc3217996, 32'h4347852e},
  {32'h450dfbe8, 32'h4172f07e, 32'hc38a1751},
  {32'hc44850d9, 32'hc3222213, 32'hc2e6e2f4},
  {32'h44ac0d6d, 32'hc3055b92, 32'h4355b625},
  {32'hc40bbb34, 32'h42ee22ca, 32'hc3dea887},
  {32'h450d8202, 32'hc3442175, 32'hc31b4cb4},
  {32'hc3120259, 32'h43abbd41, 32'hc39603d7},
  {32'h440ea2fe, 32'h43afa9ac, 32'h41f6fb18},
  {32'hc3dc1f14, 32'hc2986a44, 32'hc2c7fb8d},
  {32'h44f41c23, 32'h436f6451, 32'h3fcaf928},
  {32'hc34a0396, 32'h43a905d3, 32'hc23f34c9},
  {32'h444278fa, 32'h42942bd5, 32'h416bb82c},
  {32'hc4afeb09, 32'h4358bbaf, 32'hc28d4a65},
  {32'h44a9f54d, 32'h433fa3fa, 32'h430ad824},
  {32'hc4d995ed, 32'hc3605d74, 32'hc2cbff17},
  {32'h43761d80, 32'hc17dc938, 32'hc2bfa7c4},
  {32'hc4290716, 32'h430cb03d, 32'hc2e5d7ac},
  {32'h44c0ab41, 32'hc3a47279, 32'hc1a31081},
  {32'hc432c0c4, 32'hc08ee0ac, 32'h42cf06f6},
  {32'h44c11a86, 32'hc398ccab, 32'hc38c3f87},
  {32'hc49c0ca8, 32'hc337e578, 32'hc33255bd},
  {32'h446b8a58, 32'h44091532, 32'h40a472dc},
  {32'hc511782c, 32'h42ac9687, 32'h439c4b97},
  {32'h43971cd4, 32'hc2e940a6, 32'h4231f84e},
  {32'hc4e06969, 32'h430ff2fa, 32'h43c16c57},
  {32'h44ec3950, 32'hc387d18b, 32'h441ec9d2},
  {32'hc45a304c, 32'hc3a36634, 32'h422b1790},
  {32'hc34c7504, 32'h42a3ef43, 32'h4349cc9b},
  {32'hc50192fc, 32'h41b47387, 32'hc33df4f1},
  {32'h44a11d87, 32'hc3864f3b, 32'h43f9d65c},
  {32'hc43d3f38, 32'hc236e4fd, 32'hc3f3cb24},
  {32'h45113da5, 32'h4288a3b2, 32'hc36a6aa3},
  {32'hc515f624, 32'hc20ebbb6, 32'h4386660d},
  {32'h44a33f51, 32'hc2118636, 32'h41dff712},
  {32'hc35da5e8, 32'hc1ddd3bd, 32'hc25ce2a3},
  {32'h43331478, 32'hc325347e, 32'hc36b30d4},
  {32'hc4f53ffe, 32'h43ea9ce6, 32'hc2b779ae},
  {32'h444715e6, 32'h4384487a, 32'hc36de53a},
  {32'hc38231d3, 32'h4385adb1, 32'h433b51a5},
  {32'h44c3c47b, 32'h43050ba4, 32'hc36d7bdf},
  {32'hc4a7e0d4, 32'h40d19022, 32'h43b51665},
  {32'h44eab8b7, 32'h41f63d15, 32'hc2a54909},
  {32'hc416f390, 32'hc2aede22, 32'hc3880c5f},
  {32'h44011546, 32'hc31796ef, 32'h438a634c},
  {32'hc4f766f8, 32'h43aea8b1, 32'h4307b130},
  {32'h44527c68, 32'h425d6dc1, 32'h41f408d5},
  {32'hc4009f4c, 32'h4310addf, 32'hc1835e54},
  {32'h44062aa0, 32'hc394cbd0, 32'hc3279b8e},
  {32'hc4b36442, 32'h4376d45a, 32'h427330e0},
  {32'h44b234f7, 32'h42364129, 32'hc2ca6e31},
  {32'hc3aa8cd8, 32'h42be4861, 32'h43a1313d},
  {32'h43c69cd8, 32'h436d850b, 32'hc39cb051},
  {32'hc3f02ba8, 32'hc2be90f5, 32'hc1b4aca8},
  {32'h44e55f89, 32'h4233289a, 32'h41179881},
  {32'h43766cb2, 32'h429cfb3d, 32'hc2100ca1},
  {32'h448b53e2, 32'hc24c93a4, 32'h431bb231},
  {32'hc4dbba1b, 32'h4211d83e, 32'hc3e863aa},
  {32'h4495786b, 32'h40e75b50, 32'hc2464e62},
  {32'hc3921898, 32'h43272f25, 32'hc391465f},
  {32'h442ac760, 32'h4315490b, 32'h425d2510},
  {32'hc485a1e7, 32'h43092bfb, 32'h4114fddd},
  {32'h44804392, 32'hc3027978, 32'h43c67807},
  {32'h43842038, 32'h42a76009, 32'h440f99bc},
  {32'h4514bdb6, 32'hc403006b, 32'h43020542},
  {32'hc47881fe, 32'h41e29c20, 32'h41f20b17},
  {32'h4510d309, 32'hc3062c66, 32'h4236d177},
  {32'hc3899ae7, 32'hc2cc2960, 32'hc190252b},
  {32'h44d3cd02, 32'hc2bb0e3f, 32'hc3affbdf},
  {32'hc51768de, 32'hc2cde0f2, 32'h41eb875c},
  {32'h4414e182, 32'hc2a0805c, 32'hc356064c},
  {32'hc4414710, 32'hc0865d48, 32'hc0c804f5},
  {32'h43f13964, 32'h43a5cd92, 32'hc1ea79d2},
  {32'hc367e0a4, 32'hc315177d, 32'hc2d35c19},
  {32'h45294386, 32'h42eb15dd, 32'h42b2a5a1},
  {32'hc5054f37, 32'hc307a406, 32'h436636b9},
  {32'h444a73a3, 32'hc0bf9ea1, 32'hc240dc85},
  {32'hc48e930a, 32'h42b7cbf7, 32'h4293a874},
  {32'h44bc12ee, 32'h43802990, 32'h40a8461f},
  {32'hc424c4b2, 32'h42800079, 32'hc3a0f38f},
  {32'h450a0e43, 32'h429017e0, 32'hc22a42ce},
  {32'hc503c5cc, 32'h430f1b55, 32'hc316bfac},
  {32'h446a92db, 32'hc3129735, 32'h43ef39ac},
  {32'hc35fe984, 32'h43292f2b, 32'hc3a5cb4f},
  {32'h446d576c, 32'hc34dac61, 32'h44165b0a},
  {32'hc49eb0b4, 32'hc1d20d00, 32'h424ebfaf},
  {32'h434253b8, 32'hc3dfe69a, 32'h4370eb1a},
  {32'hc50c394f, 32'hc374547f, 32'h41975848},
  {32'h445c2a3a, 32'h42c3c40a, 32'hc3964c3f},
  {32'hc23052a0, 32'hc39cf75f, 32'h43534aaa},
  {32'h42ee7a21, 32'h42e73130, 32'hc1b6a68d},
  {32'hc4d8155a, 32'hc394f23f, 32'h432a44f6},
  {32'h44ad67cd, 32'h43869aa4, 32'h4301b067},
  {32'hc4c31a37, 32'hc3404ca7, 32'hc32ef386},
  {32'h450fc377, 32'h4388a7c0, 32'h43eb6d9a},
  {32'hc51261bf, 32'h431a43f5, 32'h42e9d4ef},
  {32'h44dc0248, 32'h42b68e9f, 32'h3f9232ad},
  {32'hc4a555dc, 32'h42d46a88, 32'hc2c3f559},
  {32'h44a3866e, 32'hc2219829, 32'h429c4d1f},
  {32'hc4fb93c7, 32'hc299e82e, 32'h43c9c7ab},
  {32'hc363f27c, 32'h43cc203f, 32'h4303b9c5},
  {32'hc4bc8503, 32'hc36f0a43, 32'hc310fa1b},
  {32'h450e8dbf, 32'h41dc05b6, 32'hc289867a},
  {32'hc505c2e2, 32'hc1f07ebe, 32'h43018285},
  {32'h450c8835, 32'h43130bfb, 32'h42d813ce},
  {32'hc2b6daf8, 32'hc32b5d75, 32'hc3161ebb},
  {32'h44f62058, 32'h42ba26b8, 32'h42a4a77d},
  {32'hc4acf290, 32'h430c1dab, 32'h42bf8c2b},
  {32'h4336bd40, 32'hc313e277, 32'h4247754a},
  {32'hc3c6e761, 32'hc3334c32, 32'hc326e3a3},
  {32'h45129b6c, 32'hc2af1cf7, 32'hc0a3d3eb},
  {32'hc4defad2, 32'h438e9eba, 32'hc3271f5c},
  {32'h44d488ba, 32'hc2e272e3, 32'h42adcdef},
  {32'hc0b74100, 32'h43c25cb4, 32'h43464196},
  {32'h43915641, 32'h4396e51c, 32'hc383ae38},
  {32'hc4859595, 32'h43ca3c0f, 32'hc2d84866},
  {32'h44e1afbe, 32'hc32c4804, 32'h437d712d},
  {32'hc50bf10a, 32'h43cca15e, 32'hc2b21896},
  {32'h43cd3732, 32'h43923f83, 32'h428e67de},
  {32'hc50a2b1b, 32'hc397f52e, 32'h42f2e9d4},
  {32'hc1bb02a0, 32'hc2693527, 32'h421b159d},
  {32'hc3421a98, 32'h427adc3c, 32'hc3a2d0eb},
  {32'h44a9656d, 32'hc30db1a2, 32'h41edf900},
  {32'hc4369784, 32'hc39987d6, 32'hc325fdd0},
  {32'h43ae28f8, 32'hc2b644ce, 32'h434c5906},
  {32'hc45775c3, 32'h43cb1ef8, 32'hc1017a18},
  {32'h44d76131, 32'h441cba70, 32'h42eb1b27},
  {32'hc4c7d0ce, 32'h4311e085, 32'h41a30f28},
  {32'h44e865a0, 32'hc2f97d5d, 32'hc399865d},
  {32'hc49f51a8, 32'h4082b109, 32'h43d18c3e},
  {32'h44bd5cdb, 32'h434bf2c6, 32'hc33e3b8f},
  {32'hc48e5964, 32'hc294b9dc, 32'h43375fe7},
  {32'h45083316, 32'h422bbd90, 32'h43b44b5f},
  {32'hc50d1219, 32'h431a09ef, 32'hc223f327},
  {32'h450260ee, 32'h43e266c3, 32'h43519e80},
  {32'hc28d7be0, 32'h4295328f, 32'hc2ffe546},
  {32'hc2cd78e0, 32'hc35ccb53, 32'h4362b976},
  {32'hc392d9e0, 32'h42f4fd9e, 32'h4119343c},
  {32'h44fa72ea, 32'hc210dc2c, 32'h42880244},
  {32'hc4adec64, 32'hc35fef2b, 32'hc418d786},
  {32'h4507249d, 32'h41ee7381, 32'hc31cc594},
  {32'hc4dbaa00, 32'h43838aab, 32'hc294c7b3},
  {32'h44d2b033, 32'hc3114c0f, 32'hc19c4ae7},
  {32'hc48ad376, 32'h434aa560, 32'hc285b0a1},
  {32'h4285e5c0, 32'hc392ad5c, 32'h423d56c2},
  {32'hc4997dee, 32'hc36a9036, 32'h42fc33ec},
  {32'h44aca40b, 32'h43066621, 32'h43424560},
  {32'hc50a2d67, 32'h415a3f5e, 32'h435c6897},
  {32'hc493fb71, 32'hc3a6fd93, 32'h43000c88},
  {32'h411ec17c, 32'hc3269e7d, 32'h41d32a8a},
  {32'hc447b5d4, 32'h42e54b83, 32'hc411c881},
  {32'h44f0d301, 32'h4140873c, 32'h43907da7},
  {32'hc438c466, 32'hc242f78c, 32'h427b7266},
  {32'h449338c8, 32'hc3a92291, 32'h43713929},
  {32'hc4ae6d3d, 32'h4270cb6c, 32'hc2fbd84a},
  {32'h445c49e6, 32'h428f4e0f, 32'hc2c763f7},
  {32'hc2946d60, 32'h42555e06, 32'hc3ab2837},
  {32'h448c3c1c, 32'hc3a4f7c8, 32'hc387b4e2},
  {32'hc4258154, 32'hc1a5db4f, 32'hc2279765},
  {32'h448742ce, 32'hc22c0cf6, 32'h43c9e81e},
  {32'hc2f92800, 32'hc229c6de, 32'hc2d6288a},
  {32'h44c47422, 32'h41e1042f, 32'h42f193fb},
  {32'hc42b3f10, 32'h43955941, 32'hc3e05c21},
  {32'h442d5396, 32'h43b80deb, 32'h4264878c},
  {32'hc4613198, 32'h427d6d9e, 32'hc33ff874},
  {32'h44cfe815, 32'hc38308f2, 32'h4376bc15},
  {32'hc2be3210, 32'h424fe35c, 32'h42bca426},
  {32'h432f6c6e, 32'hc39979cd, 32'h4321b06b},
  {32'hc4faf86f, 32'h4288b55c, 32'hc0e9e5d6},
  {32'h44d03c56, 32'hc236da64, 32'hc2a6a1df},
  {32'hc4f53d13, 32'hc1be6b3a, 32'h43219b85},
  {32'h44b56832, 32'h42bbf83f, 32'h42f79f2f},
  {32'hc4a2ff54, 32'hc2d3ef65, 32'hc39adb4f},
  {32'h44d3fbb2, 32'h43d29ca8, 32'h41c4a1fd},
  {32'hc416df79, 32'hc259f5f4, 32'h4329e8a9},
  {32'h449dfc53, 32'h41af7318, 32'h43b86a88},
  {32'hc510429b, 32'hc2f66c2f, 32'h43175140},
  {32'h44d9e91d, 32'h4233a1d1, 32'h431af1b8},
  {32'hc4dae916, 32'h437d62e1, 32'hc42117d6},
  {32'h43a1c158, 32'h40f5660c, 32'h438032ea},
  {32'hc3893ea0, 32'h4206fa96, 32'hc39473d9},
  {32'h45034154, 32'hc387e104, 32'h43adfabc},
  {32'hc4df9a5e, 32'h439745d5, 32'hc364ab30},
  {32'h4421ee2e, 32'hc3ae1161, 32'h437d58c9},
  {32'hc501bb1c, 32'hc2e81a91, 32'hc3f6485e},
  {32'h45025846, 32'h42f4fad8, 32'h432b0064},
  {32'hc496f351, 32'h4345277d, 32'hc2c1f50d},
  {32'h440f164f, 32'hc2bcf996, 32'hc19e1c11},
  {32'hc4c02f35, 32'hc273170e, 32'h43602609},
  {32'h4434350f, 32'h42df9c54, 32'hc39314e0},
  {32'hc4fa5586, 32'hc3a97164, 32'hc397b963},
  {32'h43f7f997, 32'h421740e0, 32'hc3de386f},
  {32'hc5093db4, 32'hc300a7d8, 32'h41d8b702},
  {32'h45119016, 32'hc1b11868, 32'hc373a05c},
  {32'hc4a1fb3c, 32'h419c806c, 32'hc1862b3a},
  {32'h4484d95c, 32'hc322a696, 32'hc3549656},
  {32'hc489b5f7, 32'h425c67c5, 32'hc0b992dc},
  {32'hc15a3400, 32'hc34959ec, 32'h4056a060},
  {32'hc4d78f33, 32'hc25d04fb, 32'hc2a42bc8},
  {32'h45173c20, 32'h42638073, 32'hc3165c25},
  {32'hc4f5f685, 32'h4382dbf7, 32'hc381956f},
  {32'h4491a1f0, 32'h4268fd32, 32'hc2402e02},
  {32'hc45bc779, 32'h4389210e, 32'hc3afb495},
  {32'h45048a0e, 32'h41ee589c, 32'hc320cb51},
  {32'hc2549a80, 32'h433132c0, 32'h42007da2},
  {32'h450612fa, 32'hc20dc503, 32'h425a1ebd},
  {32'hc5082c93, 32'hc3931e08, 32'h4380236e},
  {32'h44f333a8, 32'h42cd741c, 32'h439b02df},
  {32'hc4fe41e8, 32'h423edad0, 32'h4347fe81},
  {32'h43503020, 32'hc3ca480f, 32'hc39b0c51},
  {32'hc4ad80af, 32'h4321387d, 32'hc28e5197},
  {32'h44c9842e, 32'hc3a947ac, 32'hc2154abf},
  {32'hc48826c0, 32'h43391bbc, 32'h4401d562},
  {32'h4505afc5, 32'h43b25e33, 32'hc2f37bf7},
  {32'hc4b2c1cc, 32'h431cd632, 32'h435222ef},
  {32'h44b7ee31, 32'hc3a82e9e, 32'hc32b9c04},
  {32'hc4862b93, 32'h431e109a, 32'hc2c71244},
  {32'h44d260a0, 32'hc31674ce, 32'h41da2445},
  {32'hc1f752c0, 32'hc3101bc5, 32'h4366a543},
  {32'h44b4bf50, 32'hc3f29770, 32'h432ab25a},
  {32'hc3ccc380, 32'h43d661ac, 32'h435aee71},
  {32'h4497db22, 32'h4373637a, 32'h4077cb09},
  {32'hc415f13c, 32'hc0a81248, 32'h43a7c5df},
  {32'h44804d02, 32'h42beb08c, 32'hc3c2ec10},
  {32'h429f5660, 32'h426c132d, 32'h41b21a3f},
  {32'h4469c62c, 32'hc30281ac, 32'h42f809d3},
  {32'h42f51720, 32'h3e3db800, 32'hc00bb9d0},
  {32'h44da0752, 32'hc3c88796, 32'h44081a69},
  {32'hc478ed89, 32'h42b39ddd, 32'h4270e58b},
  {32'hc377b030, 32'hc23af7f8, 32'hc23cc7fb},
  {32'hc1f4c2f2, 32'h440c58e2, 32'hc3d25b73},
  {32'h451c56d0, 32'hc246547a, 32'hc318f294},
  {32'hc4d58cbf, 32'h43b4181e, 32'h43a08668},
  {32'h44e2b93c, 32'h42fd8263, 32'hc20ace62},
  {32'hc40d765c, 32'h41f8b3a9, 32'h42825312},
  {32'h4441e9ac, 32'h44011f2b, 32'hc39a63d8},
  {32'hc45a0ee7, 32'h42b82d73, 32'h4387d1bd},
  {32'h44b52620, 32'h433fdadf, 32'h4262602d},
  {32'hc4abb8ef, 32'h43a88900, 32'hc3ac6575},
  {32'h44dbf4d5, 32'h421a2535, 32'hc30a8f7d},
  {32'hc4e566ce, 32'h432e7c7c, 32'hc006ab26},
  {32'h442b3a27, 32'h43403629, 32'hc2ab329c},
  {32'hc49ea927, 32'h4409504f, 32'h424f97c9},
  {32'h451306db, 32'h41c681c5, 32'hc3d8bcc3},
  {32'hc4e2c5d5, 32'hc3031754, 32'h423f396d},
  {32'h44772644, 32'h42d0c778, 32'hc3228f27},
  {32'hc4f4b5f7, 32'h433224d2, 32'h42f6a47b},
  {32'h44ce5e69, 32'hc314dd85, 32'h43455a1c},
  {32'hc512e8cc, 32'h425bf5a4, 32'h414fa59e},
  {32'h44990950, 32'h42869aa5, 32'h43cfc117},
  {32'hc4150e4a, 32'h42612fdb, 32'h41f8c0d1},
  {32'h4413d1d0, 32'h44005f18, 32'h440f76e3},
  {32'hc1896240, 32'h421901fb, 32'h40920602},
  {32'h449382e6, 32'hc3845a3b, 32'hc329d785},
  {32'hc4d19696, 32'h42d680db, 32'h430abc00},
  {32'h4510da98, 32'h42877ce8, 32'hc34bf792},
  {32'hc46e08b9, 32'h42a32c4b, 32'hc30f79ce},
  {32'h44ae0ad7, 32'h43890829, 32'h42e991d5},
  {32'hc5096d61, 32'hc2cbb0fb, 32'hc2bd6a6a},
  {32'h44f70853, 32'h432a7e8d, 32'hc3bfaa6d},
  {32'hc2dd1997, 32'h439b0720, 32'h42da7447},
  {32'h43a25938, 32'hc2f26ed2, 32'h4330c642},
  {32'hc3adb612, 32'h42b31f9a, 32'h4199c329},
  {32'h44c6fd1e, 32'h43c1cc0f, 32'hc40b377e},
  {32'hc410621c, 32'h43974b6a, 32'h42e1c23a},
  {32'h44c6e23b, 32'hc397f427, 32'hc3593cd7},
  {32'hc48ca1a7, 32'hc3029aec, 32'h43201d11},
  {32'h4435b154, 32'hc217986c, 32'h43660e5b},
  {32'hc456e85c, 32'h41eb2156, 32'hc31cedc4},
  {32'h433d37e0, 32'hc205ec48, 32'hc30f5764},
  {32'hc442545c, 32'hc34eb480, 32'h4318d1b7},
  {32'h43f024a8, 32'h42a4103e, 32'hc1dea5f7},
  {32'hc45b966a, 32'hc31c05f5, 32'h4340e388},
  {32'h4440253e, 32'hc3b7c351, 32'hc19f9960},
  {32'hc4ddf4ca, 32'h43a77ed2, 32'h42a55d7e},
  {32'h44cc32e8, 32'hc2b26e9e, 32'h42dc9636},
  {32'hc4002e0e, 32'h409e7194, 32'hc37cad21},
  {32'h44d44229, 32'hc39fc5cf, 32'hc3dfc1de},
  {32'hc4413ec7, 32'hc35657d4, 32'hc2d57afe},
  {32'h446ff3ae, 32'hc34d5f95, 32'h433d0c5a},
  {32'hc39f3006, 32'hc2c80566, 32'h431a0349},
  {32'h432be3ed, 32'h43710053, 32'hc379f8ed},
  {32'hc2d0e8f8, 32'hc37cdc8b, 32'hc2253ad3},
  {32'h42ee2a38, 32'hc3041a3a, 32'hc386442f},
  {32'hc4019645, 32'h42724619, 32'hc3ca1b9e},
  {32'h43824bbe, 32'h4368fcd9, 32'hc30c4516},
  {32'hc5086995, 32'hc0a452ef, 32'h43cce399},
  {32'h44a74d5c, 32'hc3b39373, 32'h42798328},
  {32'hc465fb6c, 32'hc0a1d03f, 32'h436fe848},
  {32'h443b8584, 32'hc33da88c, 32'h4372820d},
  {32'hc4cafae1, 32'h43a61a15, 32'h4302606a},
  {32'h44ddfec9, 32'hc3863d2f, 32'hc2f4be39},
  {32'hc3f112fe, 32'h439a41fa, 32'hc39e2d9e},
  {32'h430a9404, 32'hc2688b45, 32'hc3b872f4},
  {32'hc4e6cecc, 32'h4131875c, 32'h430e30e5},
  {32'h4516370e, 32'h43057ec1, 32'hc28840ad},
  {32'hc4aa93b0, 32'hc39160cb, 32'h42f68185},
  {32'h449672e8, 32'h43a68bec, 32'hc2842444},
  {32'hc4f04ca0, 32'h430cc4d7, 32'hc2d01c16},
  {32'h4385b6ed, 32'h42bee4c1, 32'h4220e74a},
  {32'hc3fba47e, 32'h43c2beec, 32'h43b9143b},
  {32'h432adc60, 32'h41aa818b, 32'h3d061200},
  {32'h4236ffa8, 32'h4353bc5f, 32'hc3cb9c2b},
  {32'h44ee1f14, 32'h43027698, 32'h420825ed},
  {32'hc44fa1c4, 32'hc345c7d2, 32'h43d45231},
  {32'h442529e2, 32'h4315bb6c, 32'hc3b5e17d},
  {32'hc49a05b0, 32'h41f67c91, 32'hc34aefe1},
  {32'h44b2ed6a, 32'hc32eea3c, 32'h43981496},
  {32'hc23bd740, 32'hc1248fbe, 32'hc2fead56},
  {32'h44bb24bf, 32'hc2aa78d9, 32'hc342db05},
  {32'hc5062f76, 32'h40ba0be2, 32'hc2bc7dfa},
  {32'h44ab4198, 32'hc22314cd, 32'hc35946ee},
  {32'hc4b8a7ad, 32'hc38d47b9, 32'h42095fec},
  {32'h448800dd, 32'h42dad472, 32'h427a9290},
  {32'hc4e098ee, 32'hc30f2902, 32'hc4110e6e},
  {32'h44cc17b4, 32'hc338fd96, 32'hc3c08827},
  {32'hc4f18577, 32'hc2543453, 32'hc3aee314},
  {32'h44fafea0, 32'hc3ae9c48, 32'h43c27562},
  {32'hc39e9959, 32'h42b25768, 32'hc2d7f134},
  {32'h44d85cef, 32'hc1cb0d48, 32'hc2793775},
  {32'hc4e71a62, 32'h432c24e6, 32'hc3a2bbec},
  {32'h4508496b, 32'h4373afd7, 32'hc3a85f14},
  {32'hc4f3c956, 32'hc2085db5, 32'hc2b7e3c4},
  {32'h44e2c4b6, 32'hc38bfec5, 32'h422265e7},
  {32'hc4758f5e, 32'h4283717c, 32'hc2d1205b},
  {32'h444c1520, 32'hc32be50d, 32'h42f7c7db},
  {32'hc438a5f3, 32'h430baca8, 32'hc3958cd9},
  {32'h449ed225, 32'h42b5ae97, 32'h431c1745},
  {32'hc4b80046, 32'h430bcc1d, 32'h411eaad0},
  {32'h429a10c0, 32'h42025638, 32'hc382a8fd},
  {32'hc41cb50c, 32'hc30c9aaf, 32'hc308bf16},
  {32'h451501fe, 32'h428cec66, 32'hc3942e00},
  {32'hc46d4462, 32'hc3173e13, 32'h425f5841},
  {32'h44bd4cfb, 32'h429e91c3, 32'h438a80f0},
  {32'hc481cda9, 32'hc2188960, 32'h4285a456},
  {32'h44f9e8c8, 32'h42cec655, 32'h415f784c},
  {32'hc4ff2760, 32'h423d5b61, 32'hc38eaad1},
  {32'h449a2e7a, 32'h430ada90, 32'h4296dea8},
  {32'hc4d824c1, 32'hc3011501, 32'hc2128b9a},
  {32'h44a8594c, 32'h4397cbbe, 32'h431bb911},
  {32'hc4ae21bf, 32'hc25e1613, 32'hc06380cf},
  {32'h44015c18, 32'hc39bd7ae, 32'h439334be},
  {32'hc3ac1120, 32'h42b75976, 32'hc3b322cf},
  {32'hc1b62400, 32'hc3b02bf0, 32'hc2804b6e},
  {32'hc4e46004, 32'h4355a4da, 32'hc2bf0e75},
  {32'hc2e87ea8, 32'hc17350e1, 32'h43d82d0c},
  {32'hc47b252e, 32'hc3510123, 32'hc37fb833},
  {32'h44d3a5ed, 32'h43dff97c, 32'hc2229d53},
  {32'hc41e7f84, 32'h430e99d8, 32'h4150a05d},
  {32'h450c6fae, 32'h43885169, 32'h43c0f6ca},
  {32'hc42e9a3c, 32'hc39d5a38, 32'hc31f8331},
  {32'h43b7b6de, 32'hc16cd740, 32'h431594f1},
  {32'hc46b3da0, 32'hc38877f0, 32'h43387b42},
  {32'h44a63b1c, 32'hc3a4b2ee, 32'h41c49d27},
  {32'hc4ae933a, 32'h431acb64, 32'h43938f5a},
  {32'h4511856e, 32'hc3975cce, 32'hc2361c97},
  {32'hc354ccc8, 32'h424d0db0, 32'hc215f613},
  {32'h411c6ac0, 32'h427d08ea, 32'hc35c6512},
  {32'hc3f587bc, 32'hc334384d, 32'h43cac69d},
  {32'h44ef2de4, 32'hc404b1e6, 32'h42eb6b79},
  {32'hc43e5f81, 32'h41440a61, 32'h41266e15},
  {32'h44361acc, 32'h42a36305, 32'hc13f1185},
  {32'hc3aa9d36, 32'hc299efb5, 32'h43892dc6},
  {32'h43cd41bd, 32'hc358e900, 32'h435c924c},
  {32'hc4d51c47, 32'hc07b7f24, 32'hc3db7d0b},
  {32'h44fa3dba, 32'h42fa9b89, 32'hc400e35c},
  {32'hc3d028c8, 32'hc343f922, 32'hc24638e1},
  {32'h44f9bdb4, 32'hc3291cca, 32'h4311bd70},
  {32'hc4bafe6f, 32'hc3e25ace, 32'h438355b5},
  {32'h44b5a64e, 32'hc357565e, 32'h43e9aef9},
  {32'hc3418a88, 32'h43a02f8e, 32'hc3966880},
  {32'h4456c427, 32'hc217d62b, 32'h431eb07f},
  {32'hc41aaf72, 32'hc38d688c, 32'hc4087efc},
  {32'h4483c63a, 32'h438dc521, 32'hc194c333},
  {32'hc404b6ad, 32'h43b80fc9, 32'h42c43c5e},
  {32'h44723108, 32'hc14ac041, 32'hc38f836d},
  {32'hc45f4dc2, 32'hc2f5b927, 32'h425e9f00},
  {32'h44e2a331, 32'hc2b653e1, 32'hc2147512},
  {32'hc500ce38, 32'h434e6429, 32'hc3bff347},
  {32'h40488200, 32'hc324a230, 32'h41e290cb},
  {32'h4222db00, 32'h4323bc38, 32'h4296e1a0},
  {32'h4423eb31, 32'h4316da3d, 32'hc2cc20bc},
  {32'hc4dd92a2, 32'hc23e571a, 32'h4206dd81},
  {32'h442c1dcf, 32'hc3d34648, 32'h436ea895},
  {32'hc4f7b87c, 32'h42f9b052, 32'h4327b2a9},
  {32'h44cdffa3, 32'hc3b3a5e9, 32'hc3c66d9f},
  {32'hc4d355f1, 32'hc2ebb155, 32'h42c59df2},
  {32'h44776b8b, 32'h435ac49c, 32'h41d1d14e},
  {32'hc4c27a88, 32'hc257e9fb, 32'hc3ba3c0e},
  {32'h44c50602, 32'h43a2eb92, 32'hc3bdede5},
  {32'h42926902, 32'hc3881795, 32'h43249109},
  {32'h44a13372, 32'hc3850db8, 32'h4328666c},
  {32'hc4928464, 32'hc34b820a, 32'h43b9289a},
  {32'h44cc2539, 32'hc35eef7a, 32'h43272369},
  {32'hc461f648, 32'h4341bcf6, 32'hc36b7dfd},
  {32'h44a9fb8e, 32'hc1231d7c, 32'h4240551f},
  {32'hc48467ec, 32'hc30d8ceb, 32'hc3c77ba9},
  {32'h4441fca4, 32'hc39124de, 32'hc39814e4},
  {32'hc44deb7a, 32'h432d0ac0, 32'hc235aa0d},
  {32'h43e08290, 32'hc1963293, 32'hc1b87bb8},
  {32'hc4869123, 32'h419834f1, 32'hbec3a678},
  {32'h43c5e7aa, 32'hc408ae85, 32'hc20dbf92},
  {32'hc504d7af, 32'h436a4013, 32'hc39cf02a},
  {32'h44b82f72, 32'hc28913e0, 32'hc3408587},
  {32'hc48dc291, 32'hc3031782, 32'hc31e56a4},
  {32'h448b7e7f, 32'h43b922ff, 32'h426e853f},
  {32'hc442bdbe, 32'h43956860, 32'hc2f71411},
  {32'h44939604, 32'hc2ee8f66, 32'hc3b683da},
  {32'hc44d0c3e, 32'hc10e0f02, 32'hc2b1dc31},
  {32'h43b07de9, 32'hc2a7bcca, 32'h43272bb7},
  {32'hc4b9b39e, 32'h43d47e02, 32'hc3b71db2},
  {32'h44e2819c, 32'hc3c5986a, 32'hc1a6ab5c},
  {32'hc4f8b386, 32'hc2ba3ac9, 32'h3f050de7},
  {32'h452b9a91, 32'h408c3507, 32'h433fa9d0},
  {32'hc4fbef63, 32'h4389e813, 32'h421a68c3},
  {32'h44d07d09, 32'hc384c066, 32'hc2b41c34},
  {32'hc3a53a46, 32'h42033d9d, 32'h431cafa9},
  {32'h43a359b8, 32'hc2bace46, 32'h43963f9c},
  {32'hc512b33f, 32'hc3923057, 32'hc3d16cbf},
  {32'hc21eb990, 32'hc36665f5, 32'hc2ed079f},
  {32'hc470ed18, 32'hc36bec0d, 32'hc3dec664},
  {32'h442e8570, 32'hc2d673f9, 32'hc34d79a5},
  {32'hc3fa530e, 32'h43e9b959, 32'hc3977b0e},
  {32'h450b7f13, 32'hc2ab210a, 32'hc22c7625},
  {32'hc3b46c0e, 32'h40c5e258, 32'hc2d7ea9e},
  {32'h42100ebc, 32'hc26cc091, 32'h425b5e09},
  {32'hc3bd7368, 32'hc27a79be, 32'hc3158028},
  {32'hc215d4c8, 32'hbf9ee51b, 32'hc27f9bd0},
  {32'hc45fcfd1, 32'h43a5f2f0, 32'hc30a35fc},
  {32'h4505740d, 32'hc2f0b918, 32'hc294ddef},
  {32'hc4bce795, 32'hc38b4c91, 32'hc2a75ea9},
  {32'h4419626e, 32'hc352681c, 32'h4280181a},
  {32'hc4f2e2df, 32'h430f9401, 32'h430dcc36},
  {32'h44ca62d5, 32'hc39d100e, 32'hc31c3c3e},
  {32'hc2db11f0, 32'h41b7fa00, 32'h432f9ef2},
  {32'h4515f53d, 32'h432a0851, 32'h4391cdf3},
  {32'hc4d2d7da, 32'hc324bde6, 32'hc329fbf0},
  {32'h445cdce4, 32'h42d55c56, 32'h427604b4},
  {32'hc46cb242, 32'hc3992197, 32'h427962c7},
  {32'h44a63cc1, 32'hc337b82a, 32'h436304f1},
  {32'hc5205804, 32'h431fa87b, 32'hc101505d},
  {32'h4488e753, 32'h431b6f42, 32'hc3afb9d9},
  {32'hc33229f0, 32'hc370016e, 32'hc3a3d0b5},
  {32'h44d538e5, 32'h40cf8f7a, 32'h439b3054},
  {32'hc4bae9b1, 32'hc1b2e59a, 32'h41dfba77},
  {32'h44b2adc0, 32'h431a1333, 32'h4294cd77},
  {32'h42f79d40, 32'h42b853d6, 32'hc35bf290},
  {32'h44b1555f, 32'h4089947e, 32'h43d9c02a},
  {32'hc382ad90, 32'hc28dec4b, 32'h41a3a122},
  {32'h444b5ab4, 32'hc3265d42, 32'hc30175b2},
  {32'hc50b1748, 32'h4330a792, 32'h40028500},
  {32'h44d379db, 32'h4386faa1, 32'h431bdcff},
  {32'hc3c6cc04, 32'hc2d6d69b, 32'h4327b7fc},
  {32'h450e2fd8, 32'hc3430a02, 32'hc2af1f74},
  {32'hc3efbf31, 32'h42b042e2, 32'h42f8b1b9},
  {32'h439655b8, 32'hc3c171c2, 32'hc3a17ce6},
  {32'hc48e03f9, 32'h42503129, 32'h4314f33e},
  {32'h44476de6, 32'h428dc7a4, 32'h43143db5},
  {32'hc456fa58, 32'h42f19b73, 32'hc2aa4fb3},
  {32'h44a8cf11, 32'hc127e8f0, 32'h42b6a916},
  {32'hc51005af, 32'hc3a7ecc7, 32'h42c2ced2},
  {32'h445cbe0e, 32'h436ca5e2, 32'h435f301e},
  {32'hc5071768, 32'hc2fdf43e, 32'h42d8204f},
  {32'h44bb0efa, 32'h42a418d9, 32'hc33c1234},
  {32'hc4c770e3, 32'h42e0a965, 32'hc399b779},
  {32'h421807a0, 32'hc29fe721, 32'h42fa5531},
  {32'hc441c04c, 32'h43d93831, 32'h4244e115},
  {32'h4368ae0c, 32'hc3d0d03e, 32'hc3921e0a},
  {32'hc50a941c, 32'h4389df57, 32'hc2c3a777},
  {32'h451948ab, 32'hc413eea8, 32'hc3ad792f},
  {32'hc448fec1, 32'hc304f95b, 32'hc3bd4cbc},
  {32'h44d140c4, 32'hc1d1c1f1, 32'h43167f7f},
  {32'hc5144260, 32'hc27f1e46, 32'hc2f97aa3},
  {32'h45080019, 32'h4361037a, 32'hc3890caf},
  {32'hc5082164, 32'h4342b824, 32'h42ee989f},
  {32'h44ce1d1b, 32'h438e88a0, 32'h4346a74b},
  {32'hc4c30677, 32'h43238e2e, 32'h41164cd8},
  {32'h44fa2c2d, 32'hc393dd70, 32'h438e533b},
  {32'h435466b0, 32'hc1e16c9f, 32'h439377fa},
  {32'h437922a8, 32'hc286bdbd, 32'h42782384},
  {32'hc5056cdd, 32'h42281579, 32'hc31cea7a},
  {32'h45149786, 32'hc34e6876, 32'hc3518fe3},
  {32'hc4461f62, 32'hc3bf12a2, 32'h43bc65f8},
  {32'h44cb6a53, 32'hc205d5b2, 32'hc23d95a2},
  {32'hc3c98660, 32'h419c7a25, 32'h42c22154},
  {32'h44bade40, 32'hc21af675, 32'h4240959d},
  {32'hc49ae4f7, 32'h4312b3c3, 32'h4200dcac},
  {32'h43e0ecb0, 32'h4325c1b4, 32'h43711e1d},
  {32'hc4e88854, 32'h419a1331, 32'h427fe4b9},
  {32'h4511d4ce, 32'hc3aaf931, 32'hc21d3973},
  {32'hc4c8973f, 32'h43f567d5, 32'h43ce1271},
  {32'h44d716c4, 32'h435b4de4, 32'hc3e6c4ff},
  {32'h429e0150, 32'hc212f87f, 32'hc23ee62d},
  {32'h44cc9f1e, 32'h423c5946, 32'hc323356a},
  {32'hc4d52f4e, 32'hc3b831c6, 32'hc2b78ca1},
  {32'h44fd671e, 32'hc35365d0, 32'hc3d7169e},
  {32'hc5106a92, 32'h43082d7a, 32'hc338723e},
  {32'h450619a1, 32'hc11b6a08, 32'hc2fd3ae7},
  {32'hc4497169, 32'hc2b59516, 32'hc256ddcd},
  {32'h44e08dce, 32'hc3cc4544, 32'hc3a291f1},
  {32'h4332552b, 32'h41fa7742, 32'hc36b7565},
  {32'h450afe00, 32'h4359996c, 32'h42d99f6f},
  {32'hc41f798a, 32'h43a1b66a, 32'h43e085a4},
  {32'h443b2797, 32'hc3a36714, 32'h4312f8cc},
  {32'hc4fa5c30, 32'hc39d7486, 32'h41beb214},
  {32'h450c2960, 32'hc2746d3d, 32'hc35c71d4},
  {32'hc3a79900, 32'hc13ba51a, 32'h43307ee0},
  {32'h44f1e13a, 32'h43b0ca77, 32'hc2c7c9f0},
  {32'hc50f4bb2, 32'h43918c7d, 32'h43202b16},
  {32'h432690d0, 32'h42d122bc, 32'h4417972c},
  {32'h4333192f, 32'hc3193a67, 32'hbde3d5a8},
  {32'h450b241c, 32'h4147ab33, 32'hc1a86726},
  {32'hc4c1bec8, 32'hc32220e3, 32'h439a87e0},
  {32'h44aeca68, 32'hc4016ffc, 32'h4335d4ee},
  {32'hc32ec670, 32'h42ba1e2a, 32'h4205c11e},
  {32'h4489f1c2, 32'hc1fdf841, 32'h431ff849},
  {32'hc4a3f088, 32'h431538ba, 32'hc37c0ff4},
  {32'h43a6064c, 32'hc3d3c9bc, 32'h438d0d98},
  {32'hc381818e, 32'h4323ec06, 32'h42a64a46},
  {32'h44e87fa0, 32'hc2bd21f1, 32'h4207a140},
  {32'hc507399c, 32'hc38e2fd7, 32'hc359517c},
  {32'h446c753b, 32'hc2e4be09, 32'h42f75c9f},
  {32'hc5047e1d, 32'h41e5f4f8, 32'h42fa4e12},
  {32'h442fc3f0, 32'h42085825, 32'hc2975dbb},
  {32'hc4802dbd, 32'h43584aa8, 32'hc2c8dca8},
  {32'h44544efc, 32'h405c61f6, 32'hc2c52107},
  {32'h41fd6600, 32'hc3a09cde, 32'hc3e4c694},
  {32'h44cb3d4a, 32'h42c84de6, 32'h43ab5f86},
  {32'hc482c35a, 32'h43d2f16e, 32'h40cbeba5},
  {32'h450b0ad1, 32'hc3484cd5, 32'h413311ff},
  {32'hc4386c19, 32'h4225d9c5, 32'h4362082a},
  {32'h45135850, 32'h40ad6150, 32'hc225e7f2},
  {32'h429d6703, 32'h4356c796, 32'h4114fc18},
  {32'h44435d26, 32'hc340f676, 32'h43356a93},
  {32'hc4ed764d, 32'hc2a1079d, 32'hc32f6c2e},
  {32'h44ceba16, 32'hc370201e, 32'hc343a9dd},
  {32'hc50e446d, 32'h4296d783, 32'h428f536c},
  {32'hc1c7817c, 32'hc3870f02, 32'h4081e91d},
  {32'hc4880efe, 32'hc317bc4c, 32'hc2904560},
  {32'h450068e0, 32'hc36b341b, 32'h42adbe51},
  {32'hc4c09dfe, 32'h3fbdfdc0, 32'h3f104240},
  {32'h4471617f, 32'hc1e3ac6c, 32'h42c10d18},
  {32'hc50a0513, 32'h438756df, 32'h430c64a4},
  {32'h442284f4, 32'hc36c3984, 32'hc3a5947f},
  {32'hc34b2611, 32'hc2dd5689, 32'h424c332a},
  {32'h44c867ea, 32'hc3a448b2, 32'hc3084e86},
  {32'hc4e46387, 32'h435c9ebb, 32'hc2b9130a},
  {32'h44e5006a, 32'h434b4790, 32'hc325da66},
  {32'hc4771655, 32'hc1ca1daa, 32'h439899ba},
  {32'h44074d84, 32'h42e8671e, 32'hc2c11120},
  {32'hc3dd37b0, 32'hc2d39ae2, 32'h4353e4e8},
  {32'h44d1657d, 32'hc35630b3, 32'hc2f18e0f},
  {32'hc507b4a0, 32'h438a1ea7, 32'hc31c5242},
  {32'h4474b44e, 32'h41896e21, 32'hc211e799},
  {32'hc4eca4b8, 32'hc391e0c7, 32'h431d98c3},
  {32'h4371c060, 32'hc2a9f1a7, 32'hc3488e9d},
  {32'hc4cff57b, 32'h430123d8, 32'h3fa69300},
  {32'h44a9d404, 32'hc2ecbe63, 32'hc3a93fc4},
  {32'hc4105f3c, 32'hc28b8e6b, 32'h42479f08},
  {32'h4498e876, 32'h42c40678, 32'h43002706},
  {32'hc44b0510, 32'h42311196, 32'h434da097},
  {32'h437e781c, 32'hc2d599f9, 32'h410c677f},
  {32'hc480e04c, 32'h42d465cc, 32'h43bdf2cd},
  {32'h448c0c57, 32'hc3c5c692, 32'hc2f082bd},
  {32'hc48a76c2, 32'h419b65e4, 32'h43ad8895},
  {32'h44dad912, 32'hc38ba6a2, 32'hc1aad0e9},
  {32'hc4c64265, 32'h417ea769, 32'h432fd186},
  {32'h44ed925d, 32'hc2980456, 32'hc3686c02},
  {32'hc443c278, 32'hc1978ab1, 32'h42dbd3e6},
  {32'h44e5021f, 32'h43216a5e, 32'hc2ce222f},
  {32'hc3e8e864, 32'h43fd9f1f, 32'h43ac93b8},
  {32'h44ba7a4c, 32'h43c22e99, 32'hc2938061},
  {32'hc457fe7a, 32'hc2aec436, 32'h42226e0e},
  {32'h446d330c, 32'hc307c7ab, 32'hc3736307},
  {32'hc4a9a945, 32'h42be3410, 32'hc11980e5},
  {32'h449309f1, 32'h4282bbf5, 32'hc38ec56a},
  {32'hc4a15018, 32'hc320076f, 32'h427e576b},
  {32'h43bb0b98, 32'h41854cc8, 32'h430f2396},
  {32'hc46bf5fa, 32'h434b3d58, 32'h422cc93e},
  {32'h4337ecd9, 32'hc3616ec0, 32'hc1d7fe32},
  {32'h44e27f11, 32'hc2b80043, 32'hc25c652a},
  {32'hc4fafb60, 32'h43b5419b, 32'hc0cb06dd},
  {32'h44682b70, 32'h42eafab9, 32'hc2c35cb3},
  {32'hc5234414, 32'h41ef2f1c, 32'hc1ec80a7},
  {32'h4491c398, 32'hc32c408a, 32'hc3c6dc7e},
  {32'hc48d9b78, 32'h43c6a123, 32'h43b91f96},
  {32'h44ef2919, 32'h43e576a4, 32'hc3c2eee1},
  {32'hc42bd036, 32'h427fe0ad, 32'hc2ccfd24},
  {32'h45089725, 32'h41a0b048, 32'h429d3fe5},
  {32'hc4dbc993, 32'hc19228b5, 32'hc35fa354},
  {32'h449b82d8, 32'hc38fef6b, 32'hc3a2163f},
  {32'hc4df615a, 32'hc34fa043, 32'h42a1e72a},
  {32'h43d14f68, 32'hc3527dbc, 32'hc2f28d72},
  {32'hc4c2ef9c, 32'hc3b2c807, 32'hc33254f3},
  {32'h438cc82d, 32'hc30a4e0d, 32'hc31f168f},
  {32'hc44fee48, 32'h4397d309, 32'hc3b6d3c4},
  {32'h450717ef, 32'hc39281e5, 32'hc389f145},
  {32'hc4b5ef56, 32'hc25c2724, 32'hc114e080},
  {32'h442b8961, 32'hc25819a1, 32'hc3378ccf},
  {32'hc4de9859, 32'h3fe8d620, 32'hc2d19527},
  {32'h422fc590, 32'h42846e27, 32'hc2ebbb1e},
  {32'hc47b3fa5, 32'h41e98e1a, 32'hc37123d8},
  {32'h4504579f, 32'h42dfab53, 32'h424c4df9},
  {32'hc4ac2057, 32'h436ad167, 32'hc30391d2},
  {32'h4517fb35, 32'h429a5dc8, 32'h4277482d},
  {32'hc34d41c8, 32'hc25a12d5, 32'h434ab708},
  {32'h44d8f5f4, 32'hc431f99d, 32'hc3eeeacf},
  {32'hc417959e, 32'hc16d83ff, 32'hc3cb2a0d},
  {32'h450c0889, 32'h43fbcd83, 32'h428ea6e0},
  {32'hc4587d98, 32'h43165bb8, 32'h4317fc8b},
  {32'h44d2e7d5, 32'hc0a14f1a, 32'h43228e05},
  {32'hc48dc409, 32'h425f01ea, 32'hc1d660ea},
  {32'h44a564c9, 32'h42533456, 32'h436bd020},
  {32'hc4543f72, 32'h4317b3de, 32'hc3365bf6},
  {32'h43b5a5ac, 32'h43572ab1, 32'h42ca4c37},
  {32'hc4dabf8c, 32'hc2a5a13d, 32'h43680aba},
  {32'h44dddebb, 32'h40b9e550, 32'h435d291d},
  {32'hc3113540, 32'h439fa05c, 32'h43b3b67b},
  {32'h4504521b, 32'hc353c5d9, 32'h4240cd3a},
  {32'hc388c938, 32'h434a068b, 32'hc3470bc9},
  {32'h43fea37f, 32'hc02b3b35, 32'hc1d1b131},
  {32'hc4c5778a, 32'h41470d40, 32'hc30ccbb8},
  {32'h443213f4, 32'hc38f5e16, 32'hc359f1d7},
  {32'hc4d62929, 32'hc3027c3f, 32'hc368df9c},
  {32'h44fdde30, 32'h42d061d2, 32'h4312ef4d},
  {32'hc4cb1ed4, 32'h4327d785, 32'h432b6e5e},
  {32'h43ecf6e4, 32'h4321d60e, 32'hc22c51cc},
  {32'hc42b99ba, 32'h43595ee7, 32'h43443b26},
  {32'h441d32e9, 32'h43897668, 32'h42f19cb0},
  {32'hc4949d26, 32'hc3a9e7af, 32'h438f2ac7},
  {32'h44ebde55, 32'hc379b67b, 32'hc3dc7332},
  {32'hc48f7982, 32'h421ead32, 32'hc2355eae},
  {32'h4499fdf4, 32'hc391e91b, 32'hc3aa7bda},
  {32'hc4ceae2b, 32'h41a19354, 32'h42bd7000},
  {32'h44b5bc32, 32'h436e7d26, 32'hc358a461},
  {32'hc1c02580, 32'h435de225, 32'hc348f8b1},
  {32'h44c274e8, 32'hc230bc34, 32'hc38fd714},
  {32'hc5036bd1, 32'hc38fd737, 32'h42acaea9},
  {32'h44e38bfb, 32'h43a2632d, 32'h3d603110},
  {32'hc50010e5, 32'h422aaeac, 32'hc4157ea4},
  {32'h42f996c0, 32'h438aca96, 32'h4396ac09},
  {32'hc4cf25ec, 32'hc32d8f44, 32'hc3852c66},
  {32'h4513662b, 32'h4134b0af, 32'hc3291701},
  {32'hc510b27e, 32'hc32b9592, 32'hc253098d},
  {32'h450c4960, 32'h442984cc, 32'hc30c4ee6},
  {32'hc3b78de4, 32'hc3316718, 32'h430926c4},
  {32'h450df2d7, 32'h4297b42a, 32'h41b2b2a0},
  {32'hc48b9ee2, 32'hc3cff1aa, 32'hc3df29c3},
  {32'h44ad0a34, 32'hc1bcc365, 32'hc21136f4},
  {32'hc4dd4027, 32'hc2d2a2ee, 32'hc1944dc0},
  {32'h44fab942, 32'hc30ddd94, 32'h42d030e8},
  {32'hc4ffdaab, 32'hc2a958d8, 32'hc30dbd98},
  {32'h449819c2, 32'h429c2ea0, 32'h43040570},
  {32'hc352b2c2, 32'h43a972f0, 32'hc2d93c6a},
  {32'h45000e3c, 32'h43573634, 32'h43737afd},
  {32'hc4fcd63d, 32'h43497248, 32'hc38c4488},
  {32'h45136abe, 32'h437fbf7e, 32'h435279c7},
  {32'hc510ab94, 32'h4345ebae, 32'h43707c51},
  {32'h445c20b0, 32'hc384667f, 32'h4350bb2d},
  {32'hc4b1ed8a, 32'h43001a5b, 32'hc35bbe5a},
  {32'h44392300, 32'hc3c27780, 32'h4346cd3b},
  {32'hc4e5a8be, 32'hc2ac93e8, 32'h43945b72},
  {32'h45188718, 32'hc3602b56, 32'hc32e257a},
  {32'hc48a688d, 32'hc36aa143, 32'hc317ad48},
  {32'h443ad300, 32'h43b51c7e, 32'h42583593},
  {32'hc445e15a, 32'hc3880133, 32'hc2edb11e},
  {32'h451094f3, 32'h43da18cc, 32'hc37ce002},
  {32'hc4da1531, 32'hc34c0b3d, 32'h432e7c07},
  {32'h450f5a42, 32'hc31c7e66, 32'hc04129c4},
  {32'hc3ef9dec, 32'hc2ac62ea, 32'hc15253bf},
  {32'h45050eed, 32'hc2a87b72, 32'h4384fafa},
  {32'hc4b67689, 32'h427e7999, 32'hc271319d},
  {32'h450d8340, 32'h42c2acd0, 32'h41de0734},
  {32'hc37407fa, 32'h43c56f39, 32'hc307a6cb},
  {32'h44d474ba, 32'h430557c5, 32'h42ac9402},
  {32'hc4fd2b9f, 32'hc28248fd, 32'h435b0fe2},
  {32'h43a1fe6b, 32'h42d01f39, 32'h43ce7aa7},
  {32'hc4be8e84, 32'h4265a25b, 32'h427b691e},
  {32'h44be936b, 32'h43409318, 32'h43fde5d0},
  {32'hc48a56bb, 32'hc34233d8, 32'h43b3179c},
  {32'h4515f210, 32'h43a69dea, 32'hc3805de0},
  {32'hc4fc5f4b, 32'hbffb1b1e, 32'hc3e1ec99},
  {32'h44067f94, 32'hc380bab0, 32'hc1fea6b3},
  {32'hc39c758c, 32'hc36f436e, 32'h43055d33},
  {32'h451b7332, 32'h41a7d5ac, 32'h4308bb91},
  {32'hc47fbb68, 32'h4148bdd5, 32'h42c0c590},
  {32'h44db05fd, 32'h43c55ebb, 32'hc39b1c38},
  {32'hc4675f06, 32'hc3504dab, 32'h42697002},
  {32'h434c0289, 32'hc2b083fe, 32'hc2fbb2ec},
  {32'hc5008967, 32'hc3281524, 32'hc3798822},
  {32'h43e27d86, 32'h4213ff72, 32'hc1b8ec44},
  {32'hc4c34b7e, 32'h4313f795, 32'h430d4a97},
  {32'h44c1a635, 32'h4368f11d, 32'hc303d118},
  {32'hc4426a66, 32'h4357f8f0, 32'h42cc8f7a},
  {32'h44f5fc63, 32'h431ed37e, 32'hc3250729},
  {32'hc5011f01, 32'h4350429c, 32'hc2099e61},
  {32'h450b2a65, 32'h4120a010, 32'hc1d0a008},
  {32'hc4c413d8, 32'hc1b4cc02, 32'hc399789d},
  {32'h44e748bd, 32'hc3e2e4ec, 32'hc29b7a7b},
  {32'hc4396ee7, 32'h42182954, 32'h40c1e850},
  {32'h4507b68c, 32'h42212007, 32'hc34aa2c9},
  {32'hc4d867d1, 32'hc26b0c94, 32'h42b12b76},
  {32'h44a740b4, 32'h436e81e0, 32'h43a0a049},
  {32'hc4b5ae82, 32'hc1ce2382, 32'h42a97611},
  {32'h44cc6f79, 32'h42849086, 32'hc33b5cb8},
  {32'hc2fb4280, 32'hc40f2f57, 32'h42b9b273},
  {32'h425fde80, 32'hc2c65418, 32'h43cb06cc},
  {32'hc48d431d, 32'hc3552b0a, 32'hc308c4ae},
  {32'h441d7f0f, 32'h42c0e0e2, 32'hc16cd55f},
  {32'hc4585f46, 32'hc29ca5a8, 32'hc313f3f3},
  {32'h43d30619, 32'hc2ca16f6, 32'h424fe8e5},
  {32'hc4e8ca06, 32'h43400438, 32'hc2c78d5e},
  {32'h44f1b694, 32'h4343735e, 32'h42d4203b},
  {32'hc4faa044, 32'hc09285e2, 32'h4352354e},
  {32'h44f3d90a, 32'h418fb413, 32'h42eee042},
  {32'hc4a453a7, 32'hc35737dc, 32'hc3aee240},
  {32'h44646e02, 32'h41b4a93e, 32'h422b6743},
  {32'hc50508b4, 32'hc37d43d9, 32'hc364deb4},
  {32'h446f9fa5, 32'hc30d5902, 32'h419260de},
  {32'hc4cfec63, 32'h440a9155, 32'h434f377c},
  {32'h4501df83, 32'h42183ad3, 32'hc3be9055},
  {32'hc4e30072, 32'hc38b8e6a, 32'hc31eabf6},
  {32'h44bb2de4, 32'h4337f710, 32'hc37d5183},
  {32'hc4e685ad, 32'h42016b37, 32'hc232de1c},
  {32'h448d9dbb, 32'h438a8cc4, 32'h42bed376},
  {32'hc3550a80, 32'h4280b00e, 32'hc29391d9},
  {32'h44a96464, 32'hc339e13e, 32'hc1c89fd1},
  {32'hc48b5ebd, 32'h42a92878, 32'hc3b1a303},
  {32'h451b9ecf, 32'h43e24200, 32'h41ff96cd},
  {32'hc4fe2ae7, 32'h42ce3085, 32'hc338c6a1},
  {32'h451182eb, 32'h4256b751, 32'hc2268d54},
  {32'hc41128a8, 32'hc3b7774a, 32'h41dfcb14},
  {32'h45000686, 32'hc1d2816d, 32'hc3ef57b4},
  {32'hc48ee12e, 32'hc2d73def, 32'h436066dd},
  {32'h44634208, 32'h42808fc8, 32'hc317082d},
  {32'hc4b90a22, 32'hc1d8649a, 32'hc3325a86},
  {32'h431441c6, 32'hc3b0eb55, 32'hc1b7ceff},
  {32'hc4fe838f, 32'hc3e2fc70, 32'hc397665a},
  {32'h4506bde8, 32'h435bc662, 32'hc3ef5188},
  {32'hc21e0741, 32'hc392250a, 32'h428f321c},
  {32'h44f19a38, 32'h43dcbfb2, 32'h42e68d8c},
  {32'hc4c04870, 32'hc2f5e3e6, 32'hc33483a6},
  {32'h43ad3155, 32'h42e6a694, 32'hc20e686a},
  {32'h42ee00d0, 32'h434eb24e, 32'hc432307c},
  {32'h44924ed0, 32'h43a0b16f, 32'h425ef50c},
  {32'hc4aa7ffb, 32'h4347c41e, 32'hbfe1b902},
  {32'h44beaf1d, 32'h429e9997, 32'h4402e35b},
  {32'hc4cdc5b4, 32'h433b7415, 32'h42436c73},
  {32'h44fde82b, 32'hc37f05f8, 32'h4347bbef},
  {32'hc49e1341, 32'h424e063a, 32'h416a675f},
  {32'h4500b9c0, 32'h4310011d, 32'h42f8bf5b},
  {32'hc4ea38ea, 32'h41bff8d8, 32'hc1c050cd},
  {32'h44bc9538, 32'hc1895abb, 32'hc2a92604},
  {32'hc4329cf8, 32'h43192194, 32'hc2efdc54},
  {32'h444a3619, 32'h43419f88, 32'hc381b22c},
  {32'hc4fbef8b, 32'h430c4f58, 32'hc2c4028a},
  {32'h44cc60b3, 32'h40ba1e33, 32'hc36cd0f2},
  {32'hc44202cc, 32'hc3c3485d, 32'h43f3026d},
  {32'h44a2fdbc, 32'hc25ad333, 32'h4368a558},
  {32'hc4e1ab78, 32'hc38638c5, 32'h431e4a09},
  {32'h4315c564, 32'h4327c515, 32'h42ec85b2},
  {32'hc4821072, 32'h4376c055, 32'h42954e2a},
  {32'h4470b637, 32'hc2730e6b, 32'hc2e4da60},
  {32'hc3f14028, 32'hc11294c4, 32'hc2e07966},
  {32'h43e99321, 32'h43167001, 32'h42e9bcaf},
  {32'hc3585e00, 32'h439a7a3b, 32'hc36e576a},
  {32'h44de0853, 32'hc37adf01, 32'h4039ad90},
  {32'hc416433e, 32'h42f6fdeb, 32'h41c6526e},
  {32'hc241e440, 32'hc29c88bb, 32'h42f11506},
  {32'hc505cb77, 32'hc110f7dd, 32'hbffa7dea},
  {32'h44de85a8, 32'h4202ccd3, 32'h43d32a09},
  {32'hc473f3b6, 32'hc3b44146, 32'h43839d18},
  {32'h44dfa0b7, 32'hc2b70164, 32'hc2e024ae},
  {32'hc49139f5, 32'hc17ef301, 32'h42e39347},
  {32'h43cdeb9c, 32'h429875bc, 32'h43185012},
  {32'hc4d16fc4, 32'h4239c38a, 32'h42761ea4},
  {32'h44d356f7, 32'h4410b208, 32'h3f3f4b00},
  {32'hc498be2e, 32'hc33f0d14, 32'h41d56f4c},
  {32'h4466dadc, 32'h42812ef3, 32'hc2c4ea9c},
  {32'hc36a5a78, 32'h4236d131, 32'h435226e3},
  {32'hc299fc28, 32'h43965c0f, 32'hc27aba70},
  {32'hc4a67bac, 32'h42b067e5, 32'hc33b7ce6},
  {32'h43b82541, 32'h43aefda1, 32'hc315d53b},
  {32'hc4ccc681, 32'h4323e2d5, 32'hc1afb09f},
  {32'h44a6bbdd, 32'hc3541254, 32'h42cb9b54},
  {32'hc5065cc6, 32'hc26cec37, 32'hc23a498c},
  {32'h436daa90, 32'h431eab4e, 32'hc3568f0a},
  {32'hc4da8e55, 32'h440ddacb, 32'h42c60e88},
  {32'h43d69c2c, 32'hc287e5f1, 32'hc0a493ca},
  {32'hc4d72e4c, 32'h431a815f, 32'h4396e6cb},
  {32'h446f466c, 32'h4310664b, 32'h4317f1f7},
  {32'hc4015e59, 32'hc23c7624, 32'h41233fc7},
  {32'hc2d88188, 32'hc2ba54fe, 32'hc345e4c0},
  {32'hc45400ab, 32'h411d565c, 32'h43840cd1},
  {32'h44b8de34, 32'h42655aa9, 32'h42a1acf4},
  {32'hc4df4b2e, 32'hc20304a7, 32'h436d6065},
  {32'h4451b4d0, 32'hc1375dca, 32'hc3171e26},
  {32'hc4ad17e5, 32'h43e01e39, 32'h438c6fab},
  {32'h44efc540, 32'hc367497f, 32'h42e8b788},
  {32'hc4976a49, 32'hc35bb2a2, 32'hc262d0b4},
  {32'h438122a8, 32'hc3903b97, 32'h42f81c73},
  {32'hc4b3c4f8, 32'h43482463, 32'hc28f2fb4},
  {32'h44b83f4a, 32'h433403fd, 32'hc32f304c},
  {32'hc46c1f90, 32'hc38f3639, 32'hc3282aac},
  {32'h44f83e94, 32'hc35d584c, 32'h41856be9},
  {32'hc4f20efe, 32'hc0d35659, 32'hc284b2c7},
  {32'h445bd52e, 32'h438aac42, 32'h42e67acf},
  {32'hc36830c0, 32'hc2f018df, 32'hc3cc1118},
  {32'h43821ed2, 32'hc388e68b, 32'hc36af4ff},
  {32'h406b2800, 32'hc372b5fe, 32'h427b0d0d},
  {32'h4485b83c, 32'hc202f8da, 32'h424770d2},
  {32'hc4f71e93, 32'h4301e136, 32'hc20a13a5},
  {32'h4437e7cd, 32'h43a2488f, 32'hc34da0e4},
  {32'h4203e33c, 32'hc1e7c80c, 32'h43bfe671},
  {32'h440c8ff0, 32'h4396eada, 32'hc3f8195f},
  {32'hc401210a, 32'hc305fbc1, 32'hc3a8abe6},
  {32'h44a2d672, 32'hc353e069, 32'hc307ad96},
  {32'hc4b36209, 32'hc2ed249e, 32'h4311b98e},
  {32'h45003e02, 32'hc3b02f80, 32'hc36fdc43},
  {32'hc4ff054d, 32'hc343cdca, 32'h423f6d63},
  {32'h44d66bea, 32'hc2be6809, 32'hc2e45f3e},
  {32'hc50392bd, 32'hc2ed8715, 32'h43ac079a},
  {32'h44f39794, 32'hc3a7e53f, 32'h438bb6ca},
  {32'hc36f70eb, 32'h43c5fb36, 32'hc400ebb5},
  {32'h45292a9f, 32'hc3964c89, 32'h424f2904},
  {32'hc494994d, 32'hc3792b7e, 32'hc3860ad5},
  {32'h43f5557c, 32'h43b80239, 32'h41775b81},
  {32'hc444c23e, 32'hc30c2981, 32'h4338efd2},
  {32'h442d124f, 32'h435c952b, 32'hc37f3c40},
  {32'hc38e15e9, 32'hc386fe43, 32'h42bc602b},
  {32'h44e5f46c, 32'h4308fed4, 32'hc3b2c2b9},
  {32'hc4d11418, 32'hc114943b, 32'h430cc0ff},
  {32'h431cac90, 32'h420ce269, 32'hc3ec206d},
  {32'hc4063562, 32'hc3a55079, 32'hc3858475},
  {32'h4427f857, 32'hc413a12f, 32'h436e6e48},
  {32'hc4f2bdd2, 32'h42e911b4, 32'hc37470fc},
  {32'h4498a214, 32'hc3976163, 32'hc36e0d0a},
  {32'hc4ffcd18, 32'hc2b4617e, 32'h41c8dae5},
  {32'h4503b89c, 32'h429a843f, 32'h433188a8},
  {32'h427c7380, 32'hc13ef302, 32'h43b97327},
  {32'h439baafb, 32'h42059d2a, 32'h41a2c91a},
  {32'hc48f7738, 32'hc3361a68, 32'h4367b9de},
  {32'h4387253c, 32'h428eb9e3, 32'hc39b5983},
  {32'hc4f46958, 32'hc2666c37, 32'hc1237160},
  {32'h43b6ea48, 32'hc2282b84, 32'h43541029},
  {32'hc501c442, 32'hc3854a1e, 32'hc34fbe2b},
  {32'h4335e34a, 32'hc2bcac91, 32'h42390b18},
  {32'hc4921107, 32'hc3b84d65, 32'hc347f89a},
  {32'h45207c1a, 32'hc30e2fe7, 32'hc2b20c0b},
  {32'hc4e6c690, 32'h434d2eb6, 32'hc387aba6},
  {32'h44b09b4a, 32'h421dcbde, 32'h43214ca4},
  {32'hc481bd7e, 32'hc3c5b4f1, 32'hc3add062},
  {32'h43c66770, 32'hc3f32182, 32'hc33103ea},
  {32'hc4bc956b, 32'hc332ddd4, 32'h41e6f228},
  {32'h44939eb2, 32'h43e4e1df, 32'hc3748207},
  {32'hc50923f9, 32'hc213f1c6, 32'h429e5c34},
  {32'h44d472e3, 32'h438b7b2b, 32'hc3a976ec},
  {32'hc3da3a5c, 32'h42b285d2, 32'hc3058bb1},
  {32'h445b3fe9, 32'hc2d7fb98, 32'hc34497ac},
  {32'hc5047855, 32'hc1d4708b, 32'h4284b582},
  {32'h44f7b2b0, 32'hc3454bf6, 32'h412f2ef4},
  {32'hc38cbd4c, 32'hc30a41ca, 32'hc2041588},
  {32'h430313d0, 32'h439c637b, 32'h435099c5},
  {32'hc4893e20, 32'hc2d94ff2, 32'h43f7f4d7},
  {32'h448992ce, 32'hbf701e30, 32'hc33c89aa},
  {32'hc4e2e8f8, 32'h431a639c, 32'hc28ead45},
  {32'h44a32089, 32'h4131b725, 32'h40f2a818},
  {32'hc4c47790, 32'h42f4415f, 32'h3fcb622c},
  {32'h413b8c80, 32'hc30e06af, 32'h43334aa2},
  {32'hc50d35b5, 32'hc3112693, 32'h42c60f6c},
  {32'h445bd5ee, 32'hc2b90f29, 32'hc372a74e},
  {32'hc4c47036, 32'h4180f8cf, 32'h43d8e4bc},
  {32'h432befe0, 32'hc3a579cf, 32'h43ecc825},
  {32'hc34c8b77, 32'h433d4d48, 32'hc2429a85},
  {32'h44e89946, 32'h437e6486, 32'h43826584},
  {32'hc2072680, 32'hc39577ad, 32'hc2d0af32},
  {32'h45022087, 32'h42236186, 32'h43bb275a},
  {32'hc4a75e05, 32'h43b739db, 32'h430750f5},
  {32'h4516df4c, 32'hc38a7d21, 32'h42cc76dc},
  {32'hc4c36578, 32'hc2912be8, 32'hc2c93124},
  {32'hc2876d90, 32'h43e32449, 32'hc3f00a38},
  {32'hc514b998, 32'hc2274ca6, 32'h438d1427},
  {32'h4401f08a, 32'hc3238c11, 32'hc327a6fb},
  {32'hc428791c, 32'hc2bf528d, 32'h42871fb7},
  {32'h446336bb, 32'hc368330e, 32'h43b32de9},
  {32'hc3ec7270, 32'h435d5d19, 32'h428fc7ec},
  {32'h44cfaea9, 32'hc261de43, 32'hc33a8c3a},
  {32'hc49b6692, 32'hc23cf420, 32'h43b19114},
  {32'h450e931e, 32'hc3a23d89, 32'h43a55ba2},
  {32'hc4be95ba, 32'hc3d44d4a, 32'h421448f0},
  {32'h44117d53, 32'hc134c43d, 32'h42ca239b},
  {32'hc4b3447c, 32'h4183edae, 32'h42ef84da},
  {32'h448a2453, 32'h439c7370, 32'h43af30f0},
  {32'hc4a4fa15, 32'h42431a9c, 32'h4363f29c},
  {32'h42b26890, 32'h43b9e333, 32'hc283bb73},
  {32'hc402674c, 32'hc32bfa9a, 32'h440d266b},
  {32'h44961945, 32'hc3182528, 32'hc354ec71},
  {32'hc4e86d0b, 32'h43936e34, 32'h428f2ce8},
  {32'h4461d12a, 32'h431a3f70, 32'hc3964780},
  {32'hc3e82d7c, 32'h42f08259, 32'h420ee191},
  {32'h44fd701c, 32'hc1b5ab8f, 32'h43076788},
  {32'hc472d9de, 32'hc36055b2, 32'h41542966},
  {32'h451488f2, 32'h4379d15e, 32'hc3304612},
  {32'hc3e3bcfe, 32'hc3d1162e, 32'hc213d4bd},
  {32'h44550180, 32'hc28c3bab, 32'h42f0efc0},
  {32'hc3a708be, 32'hc1e80ec6, 32'h4295575b},
  {32'h442bc0d0, 32'h42f0466e, 32'h41e0cfc9},
  {32'hc496924a, 32'h424627e1, 32'h429fbece},
  {32'h44f9bb1c, 32'h43c989e4, 32'hc384783c},
  {32'hc4a9c3dd, 32'h4277d5e3, 32'hc2c46084},
  {32'h44ff882c, 32'h435b394d, 32'h4304cc0e},
  {32'hc3c1d449, 32'hc2f45332, 32'h432f7c62},
  {32'h44fd984d, 32'h43213bee, 32'hc354a336},
  {32'hc5037deb, 32'hc3a8028e, 32'h43a7c9c1},
  {32'h449e45bc, 32'hc262a158, 32'h438ae59a},
  {32'hc4bbde18, 32'h42c94b82, 32'h4233e717},
  {32'h450dcb0e, 32'hc400f09a, 32'hc38dadab},
  {32'hc32f5188, 32'hc32b0a47, 32'h428215be},
  {32'hc249dd40, 32'hc268591c, 32'h43a679d5},
  {32'hc4a09e24, 32'h41b68b77, 32'hc448effe},
  {32'h44927ef2, 32'hc30d2b9d, 32'h42db1547},
  {32'hc4a4cdce, 32'h439adaf2, 32'h4142b4e9},
  {32'h44db30ab, 32'h43db123e, 32'h43b81615},
  {32'hc4a3045b, 32'hc1cae4d7, 32'h41f12e6a},
  {32'h44b3a6d3, 32'h43aa6815, 32'hc33210d7},
  {32'hc3b04b4a, 32'hc37dcb65, 32'hc38f689f},
  {32'h44dbd975, 32'hc20566a7, 32'hc32ef0f2},
  {32'hc51b02ce, 32'h43c4ff60, 32'h440073f8},
  {32'h440041cf, 32'h4125afe8, 32'h424f01fc},
  {32'hc3c68060, 32'hc24c60a0, 32'h41cf5e96},
  {32'h44d208e7, 32'h420a41ba, 32'h43290932},
  {32'hc4fcfc0b, 32'h43485308, 32'hc0bd890c},
  {32'h447b652a, 32'hc2e4c332, 32'h410edfe0},
  {32'hc505927f, 32'h423653cf, 32'hc29fa8f4},
  {32'h451fd4f4, 32'h4396921f, 32'hc37941c8},
  {32'hc3bc9046, 32'hc32a9779, 32'hc32b7937},
  {32'h450aceb8, 32'h410c913d, 32'hc174c011},
  {32'hc4242c74, 32'hc3d3fe91, 32'hc2eb0013},
  {32'h42cad878, 32'h438cc2b2, 32'h430d58f9},
  {32'hc38320b7, 32'hc17108d7, 32'hc1eccd0a},
  {32'h44c6ed14, 32'hc1fa5e67, 32'hc393636c},
  {32'hc4bdf6a3, 32'h437c689f, 32'h433e24e1},
  {32'h451b0970, 32'hc337f847, 32'hc343a54d},
  {32'hc454fc7e, 32'hc2fa7fe9, 32'h432fdf48},
  {32'h4448f68a, 32'hc390649c, 32'h42aaee24},
  {32'h4312b6b0, 32'h4315be16, 32'hc38df8ae},
  {32'h42a79900, 32'hc306329e, 32'h43594bc8},
  {32'hc2965da0, 32'h42f318a3, 32'h421e6f7d},
  {32'h4408bb9b, 32'hc2c65a2d, 32'h42ea1043},
  {32'hc513cc26, 32'h435a56ea, 32'h43ad6aad},
  {32'h448cc667, 32'h43a32e6f, 32'hc2d12a02},
  {32'h42c71e57, 32'hc376cb02, 32'hc31afb97},
  {32'h44ddcd6f, 32'h43bacfe2, 32'h428a9eac},
  {32'hc50b7d80, 32'h4300c6a6, 32'hc26aa012},
  {32'h445a2844, 32'hc2fe299e, 32'h4354efec},
  {32'hc5057131, 32'hc3a91dff, 32'hc30ee853},
  {32'h44f8eef6, 32'h435c6832, 32'hc2f7908c},
  {32'hc4302f69, 32'h426d273a, 32'hc2b5cb01},
  {32'h44bb49b8, 32'h4347d962, 32'h43b45b01},
  {32'hc4a1a3aa, 32'h435878d3, 32'hc285f3c1},
  {32'h44ed89ac, 32'hc2335a6e, 32'hc2b69276},
  {32'hc4ddf400, 32'h422e3b46, 32'h437df1dd},
  {32'h451006a7, 32'h41bc196e, 32'h43262886},
  {32'hc4bf11aa, 32'h433b8f32, 32'hc42de3e4},
  {32'h4483bb6f, 32'hc20be653, 32'hc2b6b1d9},
  {32'hc3b02e12, 32'hc2ffc150, 32'hc2123043},
  {32'h449f2635, 32'hc2fdad69, 32'hc2ee2a9f},
  {32'hc3125c10, 32'hc2cdd16a, 32'h4328b1d7},
  {32'h44a548f5, 32'h439c42ae, 32'hc2bb1c56},
  {32'hc5131dbd, 32'h3fc555de, 32'h4267385a},
  {32'hc2974bdc, 32'h4312cf0b, 32'hc3085837},
  {32'h438ce921, 32'hc423e32c, 32'hc302d2b5},
  {32'h448d7e75, 32'h435682cd, 32'hc1199a5c},
  {32'hc4d1cf81, 32'h43733fc8, 32'h432380cb},
  {32'h44313100, 32'hc2faed23, 32'hc3306c43},
  {32'hc449968e, 32'hc38e21dc, 32'hc36985a3},
  {32'h445ee6e0, 32'hc1c89384, 32'h4348548c},
  {32'hc377fcf6, 32'h43b6ee16, 32'hc3a65a6f},
  {32'h43a121e4, 32'h430f34ac, 32'hc23a04f3},
  {32'hc4378218, 32'h432aa7fd, 32'h42033748},
  {32'h45205be7, 32'hc3546588, 32'hc344e70f},
  {32'hc4028a28, 32'h42d8f0e9, 32'hc30e5a7a},
  {32'h43c9e500, 32'hc1ad42e6, 32'h41849298},
  {32'hc4eacab2, 32'hc20dd671, 32'hc35b91c8},
  {32'h436c64fc, 32'hc369c110, 32'h43a90220},
  {32'hc49cb278, 32'h432f08eb, 32'hc35f16bf},
  {32'h44a700e6, 32'h41800381, 32'hc28b7ad9},
  {32'h41ac3a00, 32'h4314a24e, 32'h43200850},
  {32'h4509d456, 32'h4380d157, 32'h42fc3002},
  {32'hc431133e, 32'hc2a6ad94, 32'h433de0c6},
  {32'h44cb1a9b, 32'hc33a6513, 32'h438017b7},
  {32'h43d6c44c, 32'hc3b67854, 32'hc23afc90},
  {32'h4478b85c, 32'hc39914b8, 32'h42c7823b},
  {32'hc45c95ef, 32'hc3c152a8, 32'h4388a4fd},
  {32'h43b72830, 32'hc321cac0, 32'hc25bab32},
  {32'hc514466a, 32'h43211dcd, 32'h43ba0f5f},
  {32'h44cc9e57, 32'h41d0bcfa, 32'h435cf750},
  {32'hc45bc1ee, 32'h43730316, 32'hc29980b3},
  {32'h447fac94, 32'hc2e09f42, 32'h430e8061},
  {32'hc48bd4e2, 32'h424fc195, 32'hc15637e4},
  {32'h43daf477, 32'h4344f6ab, 32'h428c7637},
  {32'hc4e1b6bb, 32'h4293e504, 32'hc3bdac3d},
  {32'h44a59af7, 32'h432cef28, 32'hc315fdaf},
  {32'hc41343c8, 32'h43c4fd1e, 32'hc3a781b5},
  {32'h44836dc2, 32'hbe851526, 32'h435a860a},
  {32'hc4f05b12, 32'h43c4e3b8, 32'hc3b66d7b},
  {32'h44a4fdb1, 32'h42f4a600, 32'hc216888b},
  {32'hc496423c, 32'h42a85c6a, 32'h42f77eea},
  {32'h438ba77c, 32'h42a6d0e8, 32'h43368156},
  {32'hc4cf072c, 32'hc34de1cc, 32'hc23fc207},
  {32'h44fa034d, 32'hc26186d1, 32'h429e8b18},
  {32'hc48a524b, 32'hc399ac00, 32'hc39963c1},
  {32'hc47d2782, 32'hc2d23b4d, 32'h432db9f8},
  {32'h43c11fbc, 32'hc391df13, 32'hc0d5bfa4},
  {32'hc5096050, 32'h432ed2f9, 32'hc3f99577},
  {32'h44da5030, 32'hc10beef2, 32'hc3c21fb1},
  {32'hc3e90c1b, 32'hc3b10112, 32'hc338c893},
  {32'h44f2affa, 32'hc29001fc, 32'h43c342f8},
  {32'hc440fd92, 32'h43266208, 32'hc34e4da5},
  {32'h44cb2b89, 32'h439b4152, 32'hc3bc72fa},
  {32'hc5128b76, 32'hc23fe388, 32'hc3042a31},
  {32'h44f184db, 32'h43428abe, 32'h436bca78},
  {32'hc504fd18, 32'hc3575106, 32'h4147f878},
  {32'h44d46649, 32'h41c86fe0, 32'hc188b7a6},
  {32'hc4c939d4, 32'h43060846, 32'hc35d9357},
  {32'h450f7d57, 32'h3f913456, 32'h4170c48b},
  {32'hc499b497, 32'h43944b25, 32'hc372e6f9},
  {32'h44c6094c, 32'hc2db9bf6, 32'hc37ebac2},
  {32'hc4a01e26, 32'h41ed95e4, 32'hc2a45472},
  {32'h44dcce6d, 32'hc3027922, 32'h431121a8},
  {32'hc4a7ee14, 32'h43457608, 32'hc29686a8},
  {32'hc274e750, 32'h429f2a20, 32'h4343c9d7},
  {32'hc4c50422, 32'h4305ec58, 32'hc31612a7},
  {32'hc2778340, 32'hc2e420ee, 32'hc25f6034},
  {32'hc4f49601, 32'hc387cf06, 32'hc31b4c6d},
  {32'h4389d5fa, 32'hc2cbc517, 32'h42238f57},
  {32'hc3f0bd55, 32'hc32f829b, 32'h42a63ed3},
  {32'h44e30644, 32'hc3d18186, 32'hc32395ae},
  {32'hc4f7f098, 32'h4377af02, 32'h42b14d32},
  {32'hc3608f3e, 32'h425de431, 32'h4304544f},
  {32'hc4cd0c30, 32'h42aec541, 32'hc33ea189},
  {32'h44fbf64d, 32'hc2c12674, 32'hc2c2181c},
  {32'hc4127951, 32'h4320d2d8, 32'hc3615eeb},
  {32'h44f0f28c, 32'h42f94e84, 32'h443584c8},
  {32'hc442dec8, 32'hc35d75a5, 32'h4306e668},
  {32'h44faf92f, 32'h4344a653, 32'h431fcf1f},
  {32'hc4c4b637, 32'hc40296cb, 32'hc332e209},
  {32'h44e08d08, 32'h422e5124, 32'hc346116c},
  {32'h42a35c14, 32'hc3054330, 32'hc0d9ef7a},
  {32'h4422f1a8, 32'h4354a74d, 32'h43824b0a},
  {32'hc2a295c0, 32'hc408e0f8, 32'h432f6768},
  {32'h449df86a, 32'h4081fff8, 32'hc208b99f},
  {32'hc4a35434, 32'hc30f0e35, 32'h438f5488},
  {32'h44fd5b34, 32'hc177aa40, 32'hc388d2c1},
  {32'hc4c35e67, 32'h42723190, 32'h435a1dbc},
  {32'h44c75394, 32'hc3b16f68, 32'h4397413d},
  {32'hc50a4704, 32'h43c13bc7, 32'hc2facea3},
  {32'h449b5d8a, 32'h41fe5260, 32'h4384a45b},
  {32'hc3a22a8a, 32'h41f1759b, 32'h3f960bd2},
  {32'h449dd298, 32'h4277f428, 32'hc3e84714},
  {32'hc4ff8f93, 32'h4357d878, 32'h422e57d4},
  {32'h450f489b, 32'hc2061148, 32'hc29c9d5a},
  {32'hc49cb308, 32'h43c14206, 32'h43455730},
  {32'h44cd8a26, 32'h4336ca44, 32'h4396224b},
  {32'hc5071958, 32'hc3ca2d3d, 32'hc33f9a8f},
  {32'h451612c2, 32'hc2ea0332, 32'h438f3ff6},
  {32'hc458a3bc, 32'hc2d3b939, 32'h42def222},
  {32'h44937b75, 32'hc3944f07, 32'hc32ea22c},
  {32'h41cdaff0, 32'h4348add4, 32'h43519547},
  {32'h44154ce6, 32'hc3bba028, 32'hc352ee32},
  {32'hc4096127, 32'hc3c117a3, 32'h43057461},
  {32'h449c0e8c, 32'h438a01e5, 32'hc31d08e6},
  {32'hc4b7e1b2, 32'h40aed16e, 32'h43513ecb},
  {32'h44e4166c, 32'hc2a07c7f, 32'hc30d62c5},
  {32'hc39a2eb5, 32'hc38bbe8d, 32'h41fc14f8},
  {32'h449c9719, 32'hc33e160d, 32'h436915e9},
  {32'hc453bb26, 32'h4166b80c, 32'h42f882cd},
  {32'h437db2b1, 32'hc3a4d517, 32'h438d1773},
  {32'hc35bdf40, 32'h4311dd83, 32'h43750e07},
  {32'h44e2fe95, 32'hc2a18628, 32'hc30d0f21},
  {32'hc45aeea2, 32'hc2a6aad8, 32'hc2120656},
  {32'h44409f44, 32'hc2811d5e, 32'h43696bb3},
  {32'hc4761c42, 32'h43d085e6, 32'hc2aeb5d1},
  {32'h44ab8fbe, 32'h422ebdd5, 32'h42e964ec},
  {32'h43176654, 32'hc305f955, 32'hc40b7ef4},
  {32'h44517c54, 32'hc2d6bc21, 32'h42f165db},
  {32'hc4fb0d96, 32'hc2dbd6c2, 32'h436faf6b},
  {32'h4493bd00, 32'hc1a45ef3, 32'h43537107},
  {32'hc48eb02d, 32'hc39928c3, 32'hc2ed761b},
  {32'h4478b4d6, 32'h41aabc21, 32'hc321290f},
  {32'hc4483210, 32'hc344435e, 32'h422f5daf},
  {32'h44c4ec0e, 32'hc2fcf349, 32'hc3efc7dc},
  {32'hc52af0c0, 32'hc3d4f5bb, 32'hc3835bb1},
  {32'h44a97d8a, 32'hc2d8c30a, 32'hc2b2b0df},
  {32'h43780796, 32'hc3d9c42b, 32'h43b19502},
  {32'h43fdd420, 32'h4341e1c0, 32'hc2b74c39},
  {32'hc4b9ccc8, 32'hc39d1abb, 32'hc389d0a3},
  {32'h44108f94, 32'hc3986f04, 32'hc2a483de},
  {32'hc43500dc, 32'h43f7e7f9, 32'h43e41b37},
  {32'hc1abda80, 32'hc3924fe4, 32'h4315b742},
  {32'hc512192a, 32'hc3856a0c, 32'hc2a7de0a},
  {32'h4385cf88, 32'h42920ff1, 32'hc328b0a5},
  {32'hc518c3a1, 32'h4263c9bc, 32'hc1f45583},
  {32'h45058b18, 32'h41cbb17f, 32'hc3474b64},
  {32'hc4be50fa, 32'hc3c2567a, 32'hc3870a1e},
  {32'h450c1260, 32'h4369efc6, 32'h43961aa6},
  {32'hc4fe70a8, 32'hc22c0d49, 32'hc38e7906},
  {32'h43b92296, 32'h4349d626, 32'h4284d80a},
  {32'hc4d5dd25, 32'hc21bd17f, 32'hc2a2a229},
  {32'h44362f10, 32'hc3428406, 32'h4020d940},
  {32'hc4f5456d, 32'hc37a1dea, 32'h42202f42},
  {32'h443c747a, 32'h43ad6489, 32'hc21920b9},
  {32'hc50e5187, 32'hc23fb804, 32'h4399d311},
  {32'h44b66530, 32'h42b12acd, 32'h43db5e22},
  {32'hc2ae2a58, 32'h42ec65d8, 32'h437e2bf0},
  {32'h44a8f6c2, 32'hc1f306cb, 32'hc3a270f2},
  {32'hc50b24b6, 32'h41bb9f90, 32'h43b419fb},
  {32'h44d5ad0a, 32'h4339db5a, 32'hc29c85f0},
  {32'hc4b322f2, 32'hc30288b9, 32'hc2068add},
  {32'h4513e8d0, 32'hc23391b5, 32'hc2b9f03e},
  {32'hc49fab73, 32'h418811c7, 32'h435b11a0},
  {32'h440b8916, 32'h43951cf3, 32'h42e0c1f5},
  {32'hc50e641c, 32'hc40cbf1b, 32'hc3983081},
  {32'h4465e964, 32'h43df2d52, 32'h43c4ff87},
  {32'hc391fd38, 32'hc308be0e, 32'hc2ce4a30},
  {32'h44c699a0, 32'h43cb01a4, 32'h436cef2e},
  {32'hc4568c4e, 32'hc378e844, 32'h44123b0a},
  {32'h44490d34, 32'hc2b0f980, 32'hc2dcb634},
  {32'hc3d28126, 32'hc3a287fb, 32'h3fc3549f},
  {32'h45003022, 32'h4253556f, 32'hc38d1535},
  {32'hc4e30523, 32'hc28947fc, 32'hc2c4bc36},
  {32'h451afc90, 32'hc390d39c, 32'hc3b43295},
  {32'hc42a4850, 32'h4315eac0, 32'hc0374cdc},
  {32'h44e18fb4, 32'hc2b815f9, 32'h422f929e},
  {32'hc4c0c910, 32'hc206683d, 32'h4311b3b9},
  {32'h4408849c, 32'hc1e7140b, 32'hc314905c},
  {32'hc49c4932, 32'h42605d0a, 32'h40c9fa13},
  {32'h43181034, 32'hbf46edc4, 32'h436f2905},
  {32'hc3dbc15c, 32'h436e9821, 32'h432cf15b},
  {32'h415e0a0a, 32'hc315b32e, 32'h4307ca32},
  {32'hc3f0fcc9, 32'hc388ef75, 32'hc271fe60},
  {32'h45255883, 32'h429558c6, 32'hc2ed7bfc},
  {32'hc4a2861b, 32'hc2f577fc, 32'h438e366b},
  {32'h44918ae6, 32'hc3d17590, 32'h43bef16a},
  {32'hc4d2e18c, 32'hc21aec3f, 32'h43414011},
  {32'h44c9fd17, 32'h42f931f9, 32'hc297d4e1},
  {32'hc38bf8c9, 32'h43b46358, 32'hc3868a27},
  {32'h45276fae, 32'h43645fa6, 32'hc195e911},
  {32'hc40eabcc, 32'hc2fcb26e, 32'h43172f7a},
  {32'h44f98f1e, 32'hc3634df4, 32'hc3abf048},
  {32'hc0e7ae00, 32'hc35cfe60, 32'hc397db3e},
  {32'h44655a90, 32'h43ac6a05, 32'h42f080c8},
  {32'hc48e2fc5, 32'h43acec4f, 32'h4304a6ec},
  {32'h44a08528, 32'h43cbbdcc, 32'hc381ad51},
  {32'hc4d2fe50, 32'hc3d893db, 32'h43a04070},
  {32'h44f9f104, 32'hc350ee2b, 32'hc0011cce},
  {32'hc475fbcc, 32'h41fd1594, 32'h437dc9dd},
  {32'h44efb291, 32'h41577c00, 32'h4354df3c},
  {32'hc4cc7154, 32'hc3051a85, 32'hc3016360},
  {32'h447f036e, 32'hc29e7dd4, 32'hc2d46ba8},
  {32'hc4945b90, 32'hc2c22056, 32'h435edf15},
  {32'h44f7267c, 32'hc266e4de, 32'h431b7608},
  {32'h42aa6e90, 32'h436ef653, 32'hc344b48b},
  {32'h449ea02e, 32'h43aac5e0, 32'hc3132ef4},
  {32'hc3dab7a6, 32'h41391d28, 32'hc34df790},
  {32'h4505b631, 32'hc395c07b, 32'hc3935b5d},
  {32'h43100e98, 32'hc2ebcbc0, 32'hc2dda662},
  {32'h4504860e, 32'hc2765cf4, 32'h430aec3f},
  {32'hc435ccde, 32'hc3c4bb4b, 32'h42c7955e},
  {32'h4499352e, 32'h429e6c06, 32'hc4069eb7},
  {32'hc49593a9, 32'h43000f1b, 32'hc2686426},
  {32'h44badadf, 32'hc35b518e, 32'h42e9bf79},
  {32'hc4d7b271, 32'h433f187a, 32'hc33d27b2},
  {32'h44f4ae98, 32'hc1edaabf, 32'hc32b273e},
  {32'hc50fe142, 32'hc3625585, 32'h42d24da8},
  {32'h44bd7689, 32'hc2ade755, 32'h419315ae},
  {32'hc5031784, 32'hc31ce831, 32'hc33f46d0},
  {32'h44758f7c, 32'hc342791e, 32'h42b06b52},
  {32'hc4cee1f3, 32'hc346979e, 32'hc1d3a15e},
  {32'h44d1b9df, 32'h42cca80a, 32'h428d4b59},
  {32'hc4d6290c, 32'hc15cc016, 32'hc190ff2e},
  {32'h4510155d, 32'hc2901bd3, 32'h42cfdbf6},
  {32'hc503be0c, 32'h43ad513a, 32'h428201dc},
  {32'h4504377c, 32'hc3205865, 32'hc32f4152},
  {32'hc4e8fff2, 32'h4358c945, 32'h43496139},
  {32'h450e044a, 32'h42a02459, 32'hc1f84cfa},
  {32'hc47a85ec, 32'h4253ca3a, 32'h42cf9c19},
  {32'h433cf438, 32'h420ba3e5, 32'h42488294},
  {32'hc4e66d4e, 32'h4396306d, 32'hc250dfd2},
  {32'h450deb56, 32'h422717e9, 32'h4345ee4d},
  {32'hc4b2c1a1, 32'h4386d972, 32'hc2bb40b8},
  {32'h44ebd5ea, 32'h416eb4e0, 32'hc2d7da26},
  {32'hc4882547, 32'hc303492a, 32'hc3a727e5},
  {32'h440ad668, 32'h42ae20eb, 32'h4187791a},
  {32'hc4e4fda0, 32'hc3f1cb9e, 32'hc3bb6b2f},
  {32'h44c25dd0, 32'hc27a71c8, 32'h431c7984},
  {32'hc3dd52cc, 32'hc1a43d77, 32'hc18ef5d0},
  {32'h44e35a40, 32'h42bed82d, 32'hc3b07477},
  {32'hc3ecc57c, 32'hc375bcf8, 32'hc36f03fd},
  {32'h45041288, 32'h4394c46f, 32'h42dd87dc},
  {32'hc4f83597, 32'h4304ae1f, 32'hc30d2dd1},
  {32'h4511e8f4, 32'hc391295e, 32'hc2be77ea},
  {32'hc481029b, 32'h42997d7d, 32'h428cb128},
  {32'h44f954b1, 32'h42612550, 32'h4399023c},
  {32'hc4418030, 32'hc0c65dec, 32'hbf02d6c0},
  {32'h45185564, 32'hc2de2336, 32'hc322c598},
  {32'hc3b072d0, 32'hc2ed1f76, 32'h4335e585},
  {32'h45203eac, 32'h437ce507, 32'h43d0409c},
  {32'hc4f57c10, 32'h4393849a, 32'hc2da1004},
  {32'h44a4c035, 32'h41ac2f3c, 32'hc3903013},
  {32'hc4c4079a, 32'hc32e4e57, 32'hc2dd85f6},
  {32'h44221eb2, 32'hc34148b1, 32'hc202cf05},
  {32'hc35502ec, 32'h42ec8306, 32'h426b2c06},
  {32'h450ab3ff, 32'h434800af, 32'h4328103f},
  {32'hc5086985, 32'hc3324d1d, 32'hc2204d1f},
  {32'h44a3a570, 32'h43c855ef, 32'h42a745d8},
  {32'hc3e96308, 32'h4105ae6e, 32'h4291c492},
  {32'h440124d6, 32'hc35568f2, 32'h434cd30c},
  {32'hc4d65206, 32'h42c4e415, 32'hc3461484},
  {32'h44ca2052, 32'hc3462bc8, 32'h43035cab},
  {32'hc16b4180, 32'hc3201516, 32'h432d420b},
  {32'hc35c41e8, 32'hc3b0dcf5, 32'h41cbb128},
  {32'hc51010e9, 32'hc2ad1c5e, 32'hc3855d28},
  {32'h4506cfaa, 32'h42e92103, 32'h438801d3},
  {32'hc4d6be7a, 32'h437162f0, 32'h42cc6393},
  {32'h419cbd00, 32'hc404b493, 32'h42db5344},
  {32'hc4e0b932, 32'hc34ba884, 32'h43ae9f71},
  {32'h42c20aa0, 32'hc35332f5, 32'h43b2693d},
  {32'hc3697be0, 32'hc3ad348b, 32'hc2e812a9},
  {32'h44ad6682, 32'hc3188361, 32'h42d90555},
  {32'hc50661a0, 32'h42ab81b5, 32'hc2c5b1cd},
  {32'h44889bcf, 32'hc2ac5038, 32'h41585188},
  {32'hc5009523, 32'hc1e70494, 32'h4292fdfc},
  {32'h43e52050, 32'h4289fb44, 32'hc36160c5},
  {32'hc4c5f5f1, 32'h4322f661, 32'h427322ea},
  {32'h4439b840, 32'hc3756430, 32'hc3e58d9f},
  {32'hc42779d4, 32'hc31ceff3, 32'h4329896e},
  {32'h44f748fe, 32'hc38cda46, 32'h434dfa42},
  {32'hc4fd36c7, 32'h43597dcd, 32'h430d9baf},
  {32'h441ad3f6, 32'h439e25d6, 32'h43bb25bb},
  {32'hc4844783, 32'h42f014d3, 32'h436c283b},
  {32'h451fc6f0, 32'h42b462ce, 32'hc318aae7},
  {32'hc40ef148, 32'hc2dcd15d, 32'h424aeb5c},
  {32'h44945c00, 32'h429241f1, 32'h42d5a31b},
  {32'hc4d302ae, 32'hc32d343d, 32'h430b2a3f},
  {32'h44fb8781, 32'h439c5f8a, 32'h42e91789},
  {32'hc42a290a, 32'hc2f40dad, 32'hc28b353f},
  {32'h4498e0b0, 32'hc3ac0b91, 32'h4336aa96},
  {32'hc50cbfe5, 32'hc3e7bf79, 32'hc2d95499},
  {32'h44d30d28, 32'h43aaf326, 32'h43bd39e1},
  {32'hc4fdbb81, 32'hc37e834c, 32'hc3886e65},
  {32'h449a5c47, 32'h435d980d, 32'hc18a8878},
  {32'h439e89e9, 32'h4281129e, 32'hc3b5d898},
  {32'h44a842b0, 32'hc315c824, 32'hc2b8207a},
  {32'hc4bcf1e9, 32'h431098d0, 32'hc2abbd78},
  {32'h451d59dd, 32'h4304641b, 32'h43324203},
  {32'hc4a088bd, 32'h42fec5ee, 32'hc3013869},
  {32'h4504dbbe, 32'hc1d6364e, 32'h431b77d5},
  {32'hc50a83bf, 32'h436a9034, 32'hc1e93f31},
  {32'h44d715a4, 32'hc22b8f40, 32'hc38a20d8},
  {32'hc4b9f429, 32'hc2310803, 32'hc06b62dc},
  {32'h44fed670, 32'h43c8740f, 32'hc17d9cec},
  {32'hc39e8188, 32'hc3203b5f, 32'h4382450e},
  {32'h44333dc7, 32'hc30953c5, 32'hc385887a},
  {32'hc299332b, 32'hc2e54bb0, 32'hc31034f8},
  {32'h4494694e, 32'hc2ab0a43, 32'h423c5900},
  {32'hc4c55632, 32'hc3ce57b0, 32'h421b91af},
  {32'h45074e43, 32'hc1b675be, 32'hbfbb1810},
  {32'hc448577a, 32'hc2de17be, 32'h436dae0d},
  {32'h4446bd6a, 32'h430ce589, 32'h439da461},
  {32'hc516d4f8, 32'hc2e5791b, 32'h4315e695},
  {32'h446fdc7f, 32'h43b73063, 32'h433ff90e},
  {32'hc356bbf0, 32'hc1903deb, 32'hc3a4bf2e},
  {32'h449f99f9, 32'h42b69f95, 32'h428c633a},
  {32'hc529b2f2, 32'h421c30e9, 32'h42475840},
  {32'h4411a480, 32'h41f1d8f5, 32'h4372225a},
  {32'hc44f4e3c, 32'hc2f4239a, 32'h4093ee0a},
  {32'h4514428f, 32'hc2ce38e5, 32'h43b71ea7},
  {32'hc4bacf86, 32'h439103ea, 32'h43a4ebe4},
  {32'h450b853c, 32'h43d49cf0, 32'hc37baba2},
  {32'hc512dded, 32'hc311aa34, 32'h43202c90},
  {32'h429c7af0, 32'hc303349b, 32'hc23a7220},
  {32'hc4ec7a61, 32'hc378859c, 32'hc2f3f1e6},
  {32'h450dec5a, 32'hc20b2888, 32'h42fe2fd6},
  {32'hc3ae7980, 32'hc3be359e, 32'hc3839b48},
  {32'h44f44604, 32'h43274e5d, 32'hc2e3b1ce},
  {32'hc500c2ae, 32'hc401a337, 32'hc2ba4b04},
  {32'h44ef9ad0, 32'h430a81f2, 32'h43126430},
  {32'hc33de143, 32'hc395428c, 32'hc2180c17},
  {32'h44512b66, 32'hbf463d82, 32'h434b9362},
  {32'hc510c989, 32'h4306dfc4, 32'hc381527a},
  {32'h4508bf13, 32'h434f2109, 32'hc2b9d251},
  {32'hc5036946, 32'h42dbdb42, 32'hc380b736},
  {32'h44748b84, 32'h423e7cd7, 32'h42a1ffbf},
  {32'hc500369a, 32'hc219cb9f, 32'h401236b2},
  {32'h44970194, 32'hc2e6d589, 32'h43195356},
  {32'hc4aea136, 32'h437366ae, 32'h418461ee},
  {32'h45249289, 32'h416af636, 32'h431cf5f3},
  {32'hc492feac, 32'hc1328707, 32'hc38882b2},
  {32'h4240d680, 32'h4283425a, 32'hc38112cc},
  {32'hc3d3fc7c, 32'hc3c5ec7d, 32'hc2df21d5},
  {32'h44fcf797, 32'h42ac74ba, 32'hc313e0ed},
  {32'hc3501080, 32'h4305cbc8, 32'hc3921a8c},
  {32'h44e1bddc, 32'h435ef0e7, 32'h43682884},
  {32'hc4fff616, 32'hc32e2814, 32'h40886052},
  {32'h4482d852, 32'h41523868, 32'hc3426a94},
  {32'hc4816cfe, 32'hc309275e, 32'h438457d5},
  {32'h44d192e5, 32'hc349be8f, 32'hc2f05684},
  {32'hc50311b3, 32'h42b8fba2, 32'hc26bb9b0},
  {32'h451a9b69, 32'h42b95854, 32'hc1c7455c},
  {32'h4205a0f2, 32'hc24a6e23, 32'hc3d8f2f4},
  {32'h449e9432, 32'hc369a210, 32'hc28d3240},
  {32'hc4a2ac8c, 32'h441430a5, 32'hc29a99ba},
  {32'h446f76ab, 32'h4325eb02, 32'hc37129e9},
  {32'hc1c6bba4, 32'hc32ba0ca, 32'h423a2013},
  {32'h4501fc85, 32'hc180a266, 32'hc3269e76},
  {32'hc4ffe25e, 32'hc3a2ffa7, 32'hc3a67f00},
  {32'h452ea4d3, 32'h435b6112, 32'h440350e0},
  {32'hc4af07c4, 32'hc33c2a3b, 32'hc2fc2007},
  {32'h45176baa, 32'h40110cf8, 32'hc38ac144},
  {32'hc50e7d9a, 32'h401adc35, 32'h41fce508},
  {32'h451647ea, 32'h439713c0, 32'h42e81a4a},
  {32'hc32c11c4, 32'hc391fd0f, 32'h424d94ec},
  {32'hc13c5880, 32'hc3944e01, 32'hc23af2ca},
  {32'hc5102731, 32'h438989a4, 32'h436bf4bc},
  {32'h45155bdb, 32'h4338b548, 32'h435e81f0},
  {32'hc32b9ed0, 32'hbf145610, 32'hc30c86e0},
  {32'h45088820, 32'hc02aac50, 32'hc1976f14},
  {32'hc3d0076a, 32'hc3a24bce, 32'hc3d0bc02},
  {32'h437bbbd0, 32'hc34d44d0, 32'h42c489f0},
  {32'hc3d2a3af, 32'hc3161e76, 32'hc40d8fac},
  {32'h450cd2e0, 32'hc3a5ff73, 32'h43c27aac},
  {32'hc4df3e02, 32'h4413915d, 32'h411fdcb2},
  {32'hc22fd440, 32'hc3a326c0, 32'hc283a0ee},
  {32'hc49596ac, 32'h43acd552, 32'hc33b8473},
  {32'h448fff3a, 32'h43022f1e, 32'h4301a4d8},
  {32'hc4ce0be0, 32'h430ccaee, 32'h42e8cb21},
  {32'hc2fd6060, 32'hc37e7c41, 32'h43c57c3a},
  {32'hc3b1c69d, 32'hc3efeb44, 32'h42cc7381},
  {32'h45061fe3, 32'h4206771e, 32'h438801f5},
  {32'hc3084bc0, 32'hc2571744, 32'h42db4f3c},
  {32'h4227ead0, 32'h43f1baed, 32'hc2cd781c},
  {32'hc4980d98, 32'hc39c482a, 32'h42a5f98b},
  {32'h45279e23, 32'h43446e1e, 32'h435720b4},
  {32'hc4b675c5, 32'hc2b33660, 32'h43988e3d},
  {32'h447048e5, 32'h438e2664, 32'hc2aa6363},
  {32'hc4c92513, 32'h415ced34, 32'hc3b17a6c},
  {32'h4491c218, 32'hc3a8ae53, 32'hc1486d1f},
  {32'hc50ee853, 32'h438cd8bb, 32'hc2c9db00},
  {32'h442b74a0, 32'hc308c9a7, 32'h4315e320},
  {32'hc4f4f492, 32'hc29f3780, 32'hc315382c},
  {32'h44b4cf22, 32'hc2fb8c4c, 32'h43c917c9},
  {32'hc4664b65, 32'hc337726c, 32'hc37e7592},
  {32'h44d212b6, 32'h43d591b6, 32'hc2117fc8},
  {32'hc436396c, 32'hc3ad76d1, 32'hc383cd3e},
  {32'h449f9878, 32'hc3209a0e, 32'h43ebd688},
  {32'hc50d5d48, 32'h42b4f213, 32'hc36ef6e2},
  {32'h44f1b948, 32'hc199807c, 32'hc3b1b8b2},
  {32'hc4dc0e12, 32'h412cfb36, 32'h4299196c},
  {32'h4443d5d3, 32'h43632dee, 32'hc2a3e96c},
  {32'hc4a7d97d, 32'h43859469, 32'hc3718595},
  {32'h4488e40b, 32'h429c2621, 32'hc31e8e5a},
  {32'hc41dd498, 32'hc37216e4, 32'hc3182e82},
  {32'h450dc3e6, 32'hc21ee2f3, 32'hc324b136},
  {32'hc329abf6, 32'hc1437e1a, 32'h43210589},
  {32'h451625c0, 32'hc2f9584f, 32'h43d062a6},
  {32'hc509cd13, 32'h43103aa2, 32'h415d387d},
  {32'h4503962b, 32'hc312440d, 32'h425145e8},
  {32'hc4f1fb66, 32'h422ce4a2, 32'h418882e1},
  {32'h44c1ba7c, 32'hc383bdf0, 32'hc3236446},
  {32'hc41d1f4c, 32'h42daa4da, 32'h419b5eb8},
  {32'h446db756, 32'hc3bf763d, 32'h4399b741},
  {32'hc3d75a4c, 32'hc20f81b4, 32'h4203da23},
  {32'h44fed067, 32'hc353267f, 32'h43293cae},
  {32'hc391d2cc, 32'hc33e3349, 32'hc38c104d},
  {32'h44c50029, 32'hc3d3def5, 32'h42be0fb8},
  {32'hc3981ad8, 32'hc3be1c38, 32'h43cd0a87},
  {32'h448439d4, 32'h43a84001, 32'h4367bb34},
  {32'hc346ea60, 32'hc2e738aa, 32'h435d4a99},
  {32'h450f4682, 32'h43ab6f24, 32'h43c75107},
  {32'hc5000e6a, 32'h4298786f, 32'h438596f7},
  {32'h4517a589, 32'hc33bbf10, 32'h43546e34},
  {32'hc4345f54, 32'h4301ff51, 32'h43be1c5a},
  {32'h44fa665e, 32'hc26e3211, 32'h43b03c79},
  {32'hc479459e, 32'hc363e3a0, 32'h41cbba1b},
  {32'h44fcb746, 32'hc2cebdbd, 32'hc2e381a5},
  {32'hc4a2f921, 32'h421d2e4c, 32'hc3a221f3},
  {32'h43f18674, 32'hc2c508ca, 32'hc2519082},
  {32'hc4e57438, 32'h433ad5ad, 32'hc2204104},
  {32'h448f1b8c, 32'hbf1268fa, 32'h4373a137},
  {32'hc3838190, 32'h42c79037, 32'h4402b031},
  {32'h447228b0, 32'h43541948, 32'hc3ead7c6},
  {32'hc38b1930, 32'hc35a5ed8, 32'h437bb95f},
  {32'h451f52ac, 32'h4365d2a0, 32'hc39fe198},
  {32'hc517a4a4, 32'h43f031c9, 32'hc3727d71},
  {32'h44866ef2, 32'h423a57e0, 32'hc1f70ca6},
  {32'hc4a65764, 32'hc2bd6751, 32'h42d43f2e},
  {32'h450977bf, 32'h42a45764, 32'h42a99ef7},
  {32'hc4130eb4, 32'hc3efae3b, 32'hc2bde8fe},
  {32'h45122d3c, 32'h42fd5765, 32'hc38e4a93},
  {32'hc4f11159, 32'hc2a0b788, 32'hc38e3dc5},
  {32'h44f04add, 32'hc3384ff7, 32'hc1efcd2a},
  {32'hc5046ac7, 32'hc23294e2, 32'hc28b319a},
  {32'h44832baf, 32'h420ae85a, 32'hc3b055a7},
  {32'hc292e2ba, 32'h43460dd4, 32'h435cbf72},
  {32'h44e2b666, 32'h424f86d8, 32'hc3111003},
  {32'hc2e716ca, 32'h43cebc07, 32'h43854cf6},
  {32'h44584bcc, 32'hc2c6d9c8, 32'hc0d0d418},
  {32'hc44d1f8e, 32'hc3a1d988, 32'hc314aa48},
  {32'h44aaafd4, 32'h444dfe88, 32'hc3277203},
  {32'hc3f61d84, 32'hc30eccd8, 32'hc1f19cec},
  {32'h43bd68a4, 32'h4323e2ca, 32'h42cf6c1d},
  {32'hc50bcdc5, 32'h4359c154, 32'hc3744937},
  {32'hc28b72bc, 32'h42c1c9fc, 32'hc406094a},
  {32'hc4a47914, 32'hc1d8a1a0, 32'hc28e2e49},
  {32'h42f2fefc, 32'hc2d39429, 32'h424e0d1b},
  {32'hc5047ed8, 32'hc3a3845a, 32'h43f4219b},
  {32'h44e2512f, 32'hc31bf050, 32'hc3c510a4},
  {32'hc49ffd41, 32'h4371fb41, 32'hbf5214d8},
  {32'h452e123f, 32'h4305bdeb, 32'hc3b8c38c},
  {32'h433d21c6, 32'h432ed4bb, 32'hc36babd1},
  {32'h445145cf, 32'h3f77dfe3, 32'h437c1e51},
  {32'hc466837c, 32'h42d4528b, 32'h43e30ce1},
  {32'h449312eb, 32'h4170aff5, 32'hc2e75202},
  {32'hc4bdc286, 32'hc2ca9b0e, 32'hc300b302},
  {32'h449dc6bb, 32'h41330caf, 32'h4340ba50},
  {32'hc42b029c, 32'h43909b0d, 32'h43a677d7},
  {32'h450dc59a, 32'hc2a7139e, 32'hc2d7a9fe},
  {32'hc39e1100, 32'h4362ff44, 32'h43069c7d},
  {32'h44f6789b, 32'h438f6ab2, 32'hc3c2c08d},
  {32'hc4a061eb, 32'hc3139816, 32'hc2bce776},
  {32'h448de845, 32'h4397f71e, 32'hc3386fb4},
  {32'hc4fc5e60, 32'h41c8342c, 32'h4161be09},
  {32'h4437e402, 32'h42bdb33b, 32'hc3296766},
  {32'hc4df1df8, 32'h4312d791, 32'hc2558eb1},
  {32'h45082247, 32'hc3629752, 32'hc3c4a2b1},
  {32'hc435c038, 32'hc385466e, 32'h4418a314},
  {32'h44ad9fa1, 32'h43a8ce04, 32'hc328cc22},
  {32'hc4eafd42, 32'hc38d9177, 32'hc1a9dab4},
  {32'h444dbf9e, 32'hc38ef4a2, 32'hc2a6852a},
  {32'hc4cae90a, 32'hc31fcc36, 32'h42e45510},
  {32'h4428e79c, 32'hc3491ed1, 32'h425393dd},
  {32'hc4c9ec51, 32'hc315f7dc, 32'h433d9955},
  {32'h449a1802, 32'h42eb77b2, 32'h42d60372},
  {32'h440ebaa8, 32'hc324d84c, 32'h4238ac6a},
  {32'hc3963ca0, 32'h41c64bd7, 32'h4292a4bb},
  {32'h43d54b02, 32'hc40c51ae, 32'hc0222790},
  {32'hc4464e92, 32'hc2af9d5f, 32'h4248dc13},
  {32'h44b9ab40, 32'hc30f42c9, 32'hc3817c0c},
  {32'hc43341ca, 32'h433ddac8, 32'h428eb5f2},
  {32'hc38752b8, 32'h41a0a126, 32'hc29fef86},
  {32'hc4e6466e, 32'hc3c5491d, 32'hc2483356},
  {32'h439596f0, 32'h4125dfbe, 32'hc316c662},
  {32'hc4edd07c, 32'h42248347, 32'hc3ba4531},
  {32'h448733a1, 32'hc22eddaa, 32'h41267d2e},
  {32'hc50c2ad1, 32'h42454e14, 32'h41106260},
  {32'h44dbaad9, 32'h43497082, 32'hc2a3c710},
  {32'hc44be95c, 32'h42eaaa39, 32'h423d50f8},
  {32'h44eae816, 32'hc3865511, 32'h421ce092},
  {32'hc4f798da, 32'h41677888, 32'h42a398c0},
  {32'h44cd8169, 32'hc34134bd, 32'h3fd86860},
  {32'hc4c475fe, 32'h43515548, 32'h434e4079},
  {32'h441614cf, 32'hc218ea5e, 32'h4389298c},
  {32'hc3e39b98, 32'h43c02bef, 32'h433518a0},
  {32'h44e2a89c, 32'h43ccf3f6, 32'h4337a9b8},
  {32'hc4d180fc, 32'h42f85c72, 32'h431eade5},
  {32'h4414175b, 32'hc34bef27, 32'hc349917b},
  {32'hc4908b9e, 32'hc35c44bc, 32'h42027554},
  {32'h44d2a854, 32'h42ac0384, 32'hc2b22abe},
  {32'hc4745208, 32'hc3807a8e, 32'h43b100f0},
  {32'h449a21fe, 32'h43854187, 32'hc2f1961c},
  {32'hc47bda33, 32'h431dee22, 32'hc32f9350},
  {32'h44f65ada, 32'hc210544b, 32'hc3a1bd03},
  {32'hc4f9a4b1, 32'h4332721e, 32'h4337c7b9},
  {32'h4493f469, 32'hc2fa5708, 32'h4320ff66},
  {32'hc4f688f7, 32'h439ddb73, 32'hc2a5ea83},
  {32'h43044464, 32'h432d799f, 32'hc3a367c0},
  {32'hc5055eb6, 32'h43281905, 32'h42a5ad6c},
  {32'h43c3907b, 32'hc36394e2, 32'hc3abc2a8},
  {32'hc39644ae, 32'hc2fb8e5f, 32'h4291057b},
  {32'h44de55e9, 32'h4313a6e9, 32'h437eb77a},
  {32'hc4897301, 32'h43729f48, 32'hc35f1556},
  {32'h4497a4ea, 32'hc3b5b3f0, 32'h43bb6b0e},
  {32'hc4d468ea, 32'h43084feb, 32'hc3465b11},
  {32'h440b70c0, 32'hc398bd28, 32'h43071184},
  {32'hc4d80ffa, 32'h4235df44, 32'hc352fe7c},
  {32'h45149c96, 32'h420824ea, 32'h42b67ccb},
  {32'hc503a7fa, 32'h4168c4a9, 32'h43b02345},
  {32'h44a619af, 32'hc190544d, 32'h42984d74},
  {32'hc498759e, 32'hc30608f7, 32'h4262e696},
  {32'h443260f0, 32'hc2598fd0, 32'hc3257e7d},
  {32'hc4989290, 32'hc302fd7d, 32'hc2719d47},
  {32'h44d3e36d, 32'h439b1eb4, 32'hc2d1bde6},
  {32'hc4a1ffc9, 32'h42ac136b, 32'hc38120a0},
  {32'h44b064f5, 32'h43641971, 32'hc2c905d7},
  {32'hc4feb458, 32'hc302ab2a, 32'h429a5af5},
  {32'h45083b5c, 32'h427b83bf, 32'h4305dd37},
  {32'hc286f9ac, 32'hc338c17a, 32'h43488709},
  {32'h450a971c, 32'h4330dfd2, 32'hc3a19104},
  {32'hc48cbcc3, 32'hc3c5e13d, 32'hc3a205dc},
  {32'h452b8929, 32'hc2300792, 32'hc32e4ddd},
  {32'hc4ce2f65, 32'hc2310d3d, 32'hc33ff360},
  {32'h44be973e, 32'hc3fdb0f3, 32'hc227a6a1},
  {32'hc5051831, 32'hc3d57098, 32'hc3a55c54},
  {32'hc3ff389a, 32'hc3b31e56, 32'hc38b22d0},
  {32'hc392f49d, 32'h429a6133, 32'hc38e31a1},
  {32'h438cb852, 32'hc2bae7cb, 32'hc0286b2f},
  {32'hc483f1f4, 32'hc1638dd7, 32'h431bc777},
  {32'h44fae6e2, 32'hc340c404, 32'h42e0977e},
  {32'hc347334e, 32'hc2af4289, 32'h43590805},
  {32'h4503ba5a, 32'h433f9ab7, 32'hc3d65513},
  {32'h41fecee8, 32'hc353d1df, 32'hc2b92008},
  {32'h445e9deb, 32'hc32074fc, 32'hc272755c},
  {32'hc4c4272f, 32'h41216a63, 32'hc31770aa},
  {32'h44d55c0e, 32'h430103bc, 32'h43cdcbe2},
  {32'hc4d5e709, 32'h42d199eb, 32'h42dc278f},
  {32'h442b1055, 32'hc33e695c, 32'hc30224a5},
  {32'hc4ef6698, 32'h434d9fa1, 32'h431b1fb8},
  {32'h4371fee8, 32'h4177978f, 32'h410d3e60},
  {32'hc4d71586, 32'hc3592f3f, 32'hc2ea9d98},
  {32'h44c35813, 32'hc385692e, 32'h42e6b7a0},
  {32'hc4f5b343, 32'h43945859, 32'hc210cd3c},
  {32'h450ad155, 32'h435c533e, 32'h428e5e20},
  {32'hc3cc45f2, 32'h4383da91, 32'h433d1aed},
  {32'h441428b2, 32'hc3b24b44, 32'h4386e740},
  {32'hc4fc59e5, 32'h438b3e43, 32'h42bc57ab},
  {32'h448fa5d3, 32'h421569cd, 32'h432bd85d},
  {32'hc47e9fb2, 32'hc291aedf, 32'h43032d45},
  {32'h44bfe66c, 32'hc214f9a6, 32'h436587e2},
  {32'hc416e457, 32'h431d9b7f, 32'h42b01332},
  {32'h44efa529, 32'hc396a135, 32'h428cb6ed},
  {32'hc36f98bd, 32'h40813155, 32'hc3723fda},
  {32'h44b2a56d, 32'hc2a145ec, 32'h432f766c},
  {32'hc505faec, 32'hc305182d, 32'h43229660},
  {32'h4428f010, 32'h4303b26e, 32'h42dc6df5},
  {32'hc42d4998, 32'h4352c2c5, 32'hc2bb4db9},
  {32'h450ee268, 32'hc33985cc, 32'hc321123b},
  {32'hc4f77d1f, 32'h4354a2c9, 32'hc386cd30},
  {32'h44d95c62, 32'h442a7c3c, 32'h43318e56},
  {32'hc4bbb3db, 32'h43422b8a, 32'h43a950f5},
  {32'h44dd4d70, 32'h41585d4b, 32'h430ba382},
  {32'hc50701f8, 32'hc380038d, 32'hc2e276d8},
  {32'h4496b144, 32'h432c1f1a, 32'h42a123ab},
  {32'hc50d086d, 32'h430403ac, 32'h4395f259},
  {32'h4514a8e4, 32'h43453661, 32'h420bd639},
  {32'hc444d992, 32'h431d58ab, 32'h434d7920},
  {32'h45219627, 32'h41ed67ff, 32'hc2a6248c},
  {32'hc48d2ab6, 32'h42e50e08, 32'h42fed8a7},
  {32'h44138c05, 32'hc3e2f7cd, 32'h42a55218},
  {32'hc4013691, 32'hc2a002a2, 32'hc2936577},
  {32'h44ca5a5e, 32'hc3d44b39, 32'hc3e44e22},
  {32'hc50901f5, 32'hc216b75f, 32'h4310dde2},
  {32'h435badd2, 32'hc3dbbbf7, 32'hc29f7456},
  {32'hc4514ba0, 32'h42972fb3, 32'h41d27d80},
  {32'h449d00b3, 32'hc3e489be, 32'hc3013b2e},
  {32'hc50708f7, 32'h439df64b, 32'hc2969f9b},
  {32'h4474c0e3, 32'h42bbfa61, 32'h434668e9},
  {32'hc4e8eeb8, 32'h43a096da, 32'hc0130088},
  {32'h43c61ce0, 32'hc2ac87ba, 32'h432c2c55},
  {32'hc4fe9916, 32'h42517380, 32'h432b89b8},
  {32'h44c95edc, 32'h41ed6a35, 32'h42fce162},
  {32'hc49f0143, 32'h4297bfb1, 32'h43d9945d},
  {32'h450e5d51, 32'h43c4041f, 32'h42328a95},
  {32'hc505751b, 32'h42ea2d73, 32'hc34f39b0},
  {32'h4437ca4e, 32'h435ab28e, 32'h439d5d01},
  {32'hc4aa16a2, 32'h42dad602, 32'hc2d9395b},
  {32'h44b2e246, 32'h431c00ce, 32'hc0f4eb60},
  {32'hc391eda8, 32'hc2c2f083, 32'hc2a78485},
  {32'h43c4d7e6, 32'hc226d937, 32'hc2ba6d6d},
  {32'hc5123708, 32'hc2266dfc, 32'h417b1223},
  {32'h44d66720, 32'h429e838e, 32'h43560a5d},
  {32'hc48f7d6e, 32'h433f5844, 32'h43174288},
  {32'h449bf804, 32'hc230815e, 32'h43a985ba},
  {32'hc4633364, 32'hc255c1ce, 32'h43803356},
  {32'h449aaf0e, 32'h43c02e52, 32'hc360d9d1},
  {32'hc4d53d42, 32'h418edee6, 32'hc0489150},
  {32'h4503494c, 32'h42ad3720, 32'h42c9ea76},
  {32'hc42e9182, 32'hc2677ea6, 32'h42d48491},
  {32'h44d5372a, 32'hc37ab239, 32'h42ec397e},
  {32'hc4421fcc, 32'hc37763da, 32'hc3ad671f},
  {32'h42f22aa4, 32'hc28e183c, 32'hc3388aca},
  {32'hc4cf6100, 32'hc2e8d9f0, 32'h440bd1e0},
  {32'h4440bc02, 32'hc381afda, 32'hc39e8389},
  {32'hc495ff54, 32'hc2e8c47a, 32'hc2384ead},
  {32'h45244204, 32'h432af24b, 32'h439bce87},
  {32'hc4f96c76, 32'h42cf4bb9, 32'h43873a73},
  {32'h443f0685, 32'hc421918f, 32'hc234bd56},
  {32'hc501da74, 32'hc2acc609, 32'h42148b5e},
  {32'h44908eaa, 32'hc311feb7, 32'h41eac031},
  {32'hc40ff666, 32'h4192946f, 32'hc3c9bbab},
  {32'h449416ce, 32'h431492a3, 32'hc2454e22},
  {32'hc4c60bd3, 32'hc2597038, 32'hc2825ba7},
  {32'h44ec4d6b, 32'hc341ca1b, 32'hc3cf0ab7},
  {32'hc2add43a, 32'h43b8e872, 32'hc318b7f4},
  {32'h443aedfe, 32'hc302df2e, 32'hc2d253c3},
  {32'hc4dc0d19, 32'hc213a241, 32'hc185255b},
  {32'h44d93812, 32'hc0aa0b70, 32'hc35ea7ff},
  {32'hc414a6b8, 32'h42e30852, 32'hc34b4b0a},
  {32'h4508a8d4, 32'h4381b7e3, 32'hc1b010e6},
  {32'hc515e335, 32'h4304e9f3, 32'h433c53ce},
  {32'h4424b65c, 32'hc3882405, 32'hc339de60},
  {32'hc505450e, 32'h4299f5dd, 32'hc3104b17},
  {32'h43969b90, 32'h42f5ad5f, 32'hc31a3ba9},
  {32'hc4797c07, 32'hc2a9ea0f, 32'h438d66cc},
  {32'h44b73b25, 32'h42a6b390, 32'h43c2008f},
  {32'h4300a570, 32'hc388105d, 32'hc3141fa1},
  {32'hc10da680, 32'hc3afa541, 32'hc2769081},
  {32'hc2815f20, 32'hc34e6154, 32'h434a60f4},
  {32'h444e6c12, 32'h432e19fa, 32'hc3bf3dbd},
  {32'hc50015f2, 32'hc31965b2, 32'hc38faad1},
  {32'h44cb85d9, 32'h4338fd70, 32'hc360cfb5},
  {32'hc3890394, 32'hc2fb1d21, 32'hc3600275},
  {32'h4459464e, 32'hc38d6378, 32'hc36a0550},
  {32'hc498a58e, 32'hc0b62690, 32'hc24f4f52},
  {32'h431c8914, 32'h42396d1b, 32'h421cf676},
  {32'hc3d278a0, 32'h444d6c0d, 32'h43e0e828},
  {32'h44c0e202, 32'hc3d20eea, 32'hc3965c7a},
  {32'hc4ec40a8, 32'h42026e8b, 32'h42beb287},
  {32'h4504ba71, 32'hc2d04d3b, 32'h423398e9},
  {32'hc4bec825, 32'h42a9381d, 32'hc347ca3b},
  {32'h43bc2665, 32'h42547d96, 32'h4379d4d1},
  {32'hc4bde3c0, 32'hc404e318, 32'h43cc806f},
  {32'h438e18f0, 32'hc2dae14c, 32'h4203e6df},
  {32'hc2fb1000, 32'hc218b5da, 32'hc370a9a1},
  {32'h44beb59a, 32'h40d77da4, 32'hc385699c},
  {32'hc4e138ce, 32'hc13ead07, 32'hc3b261a7},
  {32'h44c3fc0a, 32'h435d49b6, 32'h432f4244},
  {32'hc432abf9, 32'h423381ad, 32'h418cd703},
  {32'h44ce8df0, 32'hc3a39558, 32'h4354968e},
  {32'h41fb1b80, 32'hc2f3eb9f, 32'h41f1fc6a},
  {32'h43a95db2, 32'h421c0811, 32'hc2264b94},
  {32'hc4063274, 32'h4328115b, 32'h41dce706},
  {32'h425ddbc0, 32'h4217305e, 32'hc3960884},
  {32'hc44510b2, 32'h427b7981, 32'h42ace2be},
  {32'h44bcbe42, 32'h4287fb77, 32'h42c8a33c},
  {32'hc3109185, 32'hc266ea6a, 32'h43a6adac},
  {32'h450c3d46, 32'h430aec18, 32'h442a4104},
  {32'hc3018738, 32'h42943124, 32'h42e1aa99},
  {32'h444d1a61, 32'hc25082fe, 32'hc3086b1a},
  {32'hc491ede5, 32'h438a7098, 32'h4197f2d2},
  {32'h43cfbeb8, 32'hc2e8bdd0, 32'hc2caf02a},
  {32'hc5031f98, 32'h42cd203c, 32'hc27b3e3f},
  {32'h44d9e7b1, 32'hc28b35ed, 32'hc3705a41},
  {32'hc50704d8, 32'h43755b1b, 32'h42687ef2},
  {32'h450f065b, 32'hc341e81a, 32'hc2dcbba4},
  {32'hc4cc9fd9, 32'hc3477a44, 32'h435440d5},
  {32'h43e6c658, 32'hc3d625ae, 32'hc0c1ef3c},
  {32'hc50a9bc9, 32'h42b6122c, 32'hc1073836},
  {32'h4501eb20, 32'hc38683c6, 32'h40a97d60},
  {32'hc4de2cb5, 32'hc3087176, 32'h42c34670},
  {32'h448009a9, 32'hc35cfe06, 32'hc220a6c1},
  {32'hc40f31c0, 32'h443dd6d8, 32'h42004f31},
  {32'h44df7333, 32'hc3fba503, 32'h434f76ea},
  {32'hc4af91a2, 32'h43178bfc, 32'hc3266306},
  {32'h44f5d0c2, 32'hc2c0145e, 32'hc281e423},
  {32'hc4ec1386, 32'h42912f32, 32'hc312ba0a},
  {32'h445cafa4, 32'hc314d347, 32'hc2aa4b49},
  {32'hc4df9e70, 32'h4426dc13, 32'hc2fd3cd8},
  {32'h43c4ba79, 32'hc2d7c6a6, 32'h419c3266},
  {32'h43008990, 32'h42195fe7, 32'hc3a36aa9},
  {32'h450f6dc4, 32'hc3b31e65, 32'hc22631c1},
  {32'hc4105e3a, 32'hc33550a3, 32'h436e466f},
  {32'h44f270ac, 32'h43786760, 32'h42e0a2f9},
  {32'hc40bd378, 32'h43e0d240, 32'h437bb61b},
  {32'h44746326, 32'hc3841ddc, 32'hc298a923},
  {32'hc3d0fb98, 32'h43c03d6e, 32'h43a86627},
  {32'h45023d1e, 32'h43b8c158, 32'h4263fe64},
  {32'hc4511542, 32'h41ed850c, 32'h43ff920b},
  {32'h44bd4f6a, 32'h433f4b52, 32'hc32315d0},
  {32'hc3db5784, 32'h42c7d795, 32'h436cbdbd},
  {32'h44efa130, 32'h42d73ab6, 32'h433c17d0},
  {32'hc38d1cfc, 32'h428160c1, 32'h43043bf6},
  {32'h450c4244, 32'hc28dda3e, 32'hc3e1fe3c},
  {32'hc4d75a70, 32'h43c5a236, 32'h422f7cea},
  {32'h44ecb4ab, 32'h43305e64, 32'hc30224c2},
  {32'hc4cc5687, 32'hc37d1a7b, 32'hc32085bf},
  {32'h43e31347, 32'hc33936f8, 32'h433df820},
  {32'hc33a00f0, 32'h41fe902a, 32'h43ab65c2},
  {32'h444d56c2, 32'h4117030c, 32'hc24eec98},
  {32'hc487e48c, 32'hc20abb81, 32'hc30ab4a6},
  {32'h44d7ad4c, 32'h429b5eae, 32'h43010f60},
  {32'hc2125d00, 32'hc263f871, 32'h4224fddf},
  {32'h4478a296, 32'h4218604a, 32'hc3115da2},
  {32'hc4fcdbec, 32'h439b28e1, 32'h41c431e1},
  {32'h43ff8980, 32'h42aeb110, 32'h434cb39e},
  {32'hc489cfc4, 32'hc250ef9b, 32'h43062b88},
  {32'h441615e2, 32'hc3b5db04, 32'h42b47a32},
  {32'hc45149d4, 32'hc36cfbda, 32'h4312d98d},
  {32'h4443935f, 32'h42b0459c, 32'hc358f848},
  {32'hc4a999e0, 32'h42b23e45, 32'h416a9db2},
  {32'h44e89fb4, 32'hc2fabd8b, 32'hc2db7fca},
  {32'hc4fa5e82, 32'hc39df7e1, 32'h4397b41f},
  {32'h45087eed, 32'h4367e44f, 32'hc2b92646},
  {32'hc422e163, 32'hc3769e09, 32'hc36d584e},
  {32'h44fd3cb4, 32'hc09003e8, 32'hc2930943},
  {32'hc465e006, 32'hc3822424, 32'h4408274f},
  {32'h43f0dd78, 32'hc404ea3c, 32'h42e1c754},
  {32'hc46c7212, 32'h43abd5ab, 32'hc3834889},
  {32'h448fc436, 32'hc078bb12, 32'hc3280769},
  {32'hc4223909, 32'h43d203ea, 32'hc399b5a1},
  {32'h44fda352, 32'hc3cecff1, 32'h4323feb4},
  {32'hc4d9e955, 32'hc28ef18e, 32'h439ec7ba},
  {32'h43ec0358, 32'hc3817ba3, 32'h42fdfcb8},
  {32'hc482d6a2, 32'h42128d6c, 32'h430b12f2},
  {32'h45166da4, 32'hc0768640, 32'hc403a412},
  {32'hc4dee569, 32'hc3cb3c20, 32'h4204a336},
  {32'h44e67a60, 32'h4325bbee, 32'hc3a3d0f4},
  {32'hc3ecb42c, 32'hc3a71e33, 32'h435ddee0},
  {32'h441209ce, 32'hc1e5bef4, 32'hc31b2fdd},
  {32'hc4c43af8, 32'hc3bfff4e, 32'h4356a404},
  {32'h44cce0ea, 32'hc3279e7c, 32'hc2a0cf34},
  {32'hc43c6070, 32'h437949b7, 32'h439fd2db},
  {32'h4495e8ec, 32'hc392471a, 32'h402b6ed9},
  {32'h42298840, 32'h4352df86, 32'hc34398ab},
  {32'h4501e560, 32'h43d10371, 32'hc23fab1f},
  {32'hc4d54a34, 32'hc2b131d8, 32'h421bec39},
  {32'h450182a9, 32'hc33cbf4c, 32'hc38209fd},
  {32'hc4920c35, 32'h438273d3, 32'h435a2061},
  {32'h442265c9, 32'hc31e4acb, 32'hc3b56ba9},
  {32'hc42c8a80, 32'h43a2c32e, 32'h429071de},
  {32'h444d2a21, 32'h430f37a3, 32'hc113dd8f},
  {32'hc4df3fd4, 32'h42c0c661, 32'h42860548},
  {32'h44563a6e, 32'h412fc66b, 32'hc33b5760},
  {32'hc3cf7268, 32'h438811af, 32'h4375b781},
  {32'h44f55a84, 32'hc314b5d4, 32'h43e65cea},
  {32'hc40e8096, 32'h438c55b9, 32'hc30d11d5},
  {32'h44e80f13, 32'h4354f9c3, 32'h420089a9},
  {32'hc480a90e, 32'hc1f916fc, 32'h42e3490c},
  {32'h447c1687, 32'hc32292a5, 32'h4287fe60},
  {32'hc5021506, 32'h438cee62, 32'hc3380b1d},
  {32'h44ed2be7, 32'hc07d012c, 32'hc2dd2e88},
  {32'hc4d56368, 32'hc2edf224, 32'hc18a72a9},
  {32'h44da6723, 32'hc39b1ce5, 32'hc2caffbe},
  {32'hc3a27255, 32'h433cc730, 32'hc3ac6838},
  {32'h44fa4c6e, 32'hc2dceb71, 32'hc351fb66},
  {32'hc4cd2b9e, 32'h43df1b23, 32'h43b20155},
  {32'h450122c4, 32'hc3ad5932, 32'hc3b4fec7},
  {32'hc5097530, 32'hc38338fa, 32'hc2fd4505},
  {32'h441d8bba, 32'h433c80b1, 32'hc3051bc8},
  {32'hc4d9705d, 32'hc3b90eec, 32'h428adc5a},
  {32'h44fd64e2, 32'hc21e2878, 32'h4389445d},
  {32'hc3fbbec6, 32'h41f5b1e9, 32'h4364cc00},
  {32'h44b13020, 32'hc29edef8, 32'hc3216339},
  {32'hc50132de, 32'h42c36ccc, 32'h433c07dd},
  {32'h44eb9d71, 32'h4454d206, 32'h4209cb34},
  {32'hc4f1d847, 32'h43734529, 32'hc231cd7e},
  {32'h44b738b6, 32'hc28b1af4, 32'hc199ef16},
  {32'hc515c544, 32'h42515aa8, 32'hc1f36654},
  {32'h43f725f8, 32'hc3104c41, 32'hc25fe281},
  {32'hc40463e2, 32'hc305bef8, 32'h42f92f60},
  {32'h45155f99, 32'hc2d529e4, 32'hc2fe0376},
  {32'hc47a79b1, 32'hc1842580, 32'h43de0806},
  {32'h44820778, 32'h426b7e7d, 32'hc36c6c73},
  {32'hc3b00790, 32'h434da934, 32'hc27c608c},
  {32'h441a76f8, 32'hc390700e, 32'hc3656bc7},
  {32'h43a02280, 32'hc302b92f, 32'h40bf3230},
  {32'h44057b4a, 32'hc3534ac9, 32'hc1afdd8f},
  {32'hc5017697, 32'hc112ad80, 32'hc36aebbd},
  {32'h4521c74f, 32'hc2065cb5, 32'hc2a0e757},
  {32'hc4d4c158, 32'h42d13fd2, 32'h43a354c6},
  {32'h44cd994a, 32'hc245f647, 32'hc33b3094},
  {32'hc4114d9c, 32'hc2dd6f34, 32'h43436c56},
  {32'h446823fc, 32'hc3d76fb1, 32'h41de02a8},
  {32'hc4b01a06, 32'h42517990, 32'h433b54a5},
  {32'h4368b508, 32'hc1952f2b, 32'h42e7824e},
  {32'hc3c84cb8, 32'h430e7f7f, 32'h42d724ef},
  {32'h44079d36, 32'h4391e83d, 32'hc312bfce},
  {32'hc49986f8, 32'h42215696, 32'h41d9b9c6},
  {32'h451462ad, 32'h4386459a, 32'hc389529e},
  {32'hc4e98212, 32'hc3865845, 32'hc0de9a4d},
  {32'h432c6ca8, 32'h4221c45e, 32'h43a4045c},
  {32'hc44df47a, 32'h43463f71, 32'h43115dda},
  {32'h4478f7f8, 32'hc3abd12e, 32'hc1f3f952},
  {32'hc4b14564, 32'h43a8e914, 32'h41e95896},
  {32'h4509da92, 32'h430b486a, 32'h43823b91},
  {32'hc4184658, 32'h4336ba42, 32'h43cd1dde},
  {32'h44f0a18d, 32'hc2fc25d4, 32'hc3f5a602},
  {32'hc50a6d4b, 32'h43c66a84, 32'h42de7de9},
  {32'h44832fe4, 32'h43563bbc, 32'h4193bf38},
  {32'hc391d290, 32'h43482f32, 32'h43a48240},
  {32'h45103abc, 32'hc31efa8c, 32'hc3848f2e},
  {32'hc47e7988, 32'h42fb1188, 32'h4384ef2c},
  {32'h4478a708, 32'hc2fe19ce, 32'hc2c314df},
  {32'hc477c3e7, 32'h438b72da, 32'hc3e54712},
  {32'h44bc00d3, 32'hc3759192, 32'h438cbb5b},
  {32'hc40b23e0, 32'hc1c99d7f, 32'hc3b2c487},
  {32'h433debd0, 32'h42d83358, 32'hc39afe3f},
  {32'hc5094054, 32'hc375e240, 32'hc3b8abd0},
  {32'h43642786, 32'hc295b350, 32'hc2f42bca},
  {32'hc41a8139, 32'h430fce82, 32'h433b32f4},
  {32'h4508e147, 32'h439d1d59, 32'hc18e744b},
  {32'hc4047975, 32'hc1d04a89, 32'hc2be2f3d},
  {32'h4406cf8a, 32'hc3297653, 32'h42a08d6e},
  {32'hc4c50eef, 32'hc3c6e8a9, 32'h43abb98d},
  {32'h4506b334, 32'hc25e8172, 32'hc36b8b31},
  {32'hc473f495, 32'hc2c610e1, 32'h42ebe681},
  {32'h45016ffa, 32'h436f4b2b, 32'hc37bf596},
  {32'hc4cf220f, 32'hc39dd9f5, 32'hc3a77586},
  {32'h450dfa19, 32'h42ef0708, 32'h420f32a8},
  {32'hc489538b, 32'hc319602c, 32'h43715b65},
  {32'h44612176, 32'h430de96c, 32'h428c26ad},
  {32'hc4de1653, 32'h441bc1f1, 32'h43ea49aa},
  {32'h441f8468, 32'hc399a45b, 32'hc33decc6},
  {32'hc3d67de8, 32'hc2001dbb, 32'h42e1a38e},
  {32'h44e4c954, 32'h4349afb2, 32'hc37e81a1},
  {32'hc454c0d8, 32'h430e18fd, 32'hc2f2ffdc},
  {32'h4426b3d6, 32'hc2045fbb, 32'h42abfb59},
  {32'hc4965119, 32'h436870d6, 32'hc24d2075},
  {32'h4401de3c, 32'h4395a233, 32'hc296ff52},
  {32'hc5131bb0, 32'h4115a49c, 32'hc1bd15e9},
  {32'h44e04b76, 32'h41b66486, 32'h416fcf36},
  {32'hc516eed4, 32'hc315775e, 32'h42920b52},
  {32'h425b2618, 32'hc2f15280, 32'h43443e11},
  {32'hc3a9ffb3, 32'h43c9cc88, 32'h422867b1},
  {32'h44cbcc41, 32'h424bbdab, 32'h4226ee94},
  {32'hc4bb0dca, 32'hc2f74bc8, 32'h43e3f721},
  {32'h4507649a, 32'hc38feb30, 32'h4387c9be},
  {32'hc50b91aa, 32'h4331c341, 32'hc3a6b1c0},
  {32'h44546032, 32'hc37998fd, 32'h4380c062},
  {32'hc4cda939, 32'h424ed29a, 32'h4328433d},
  {32'h4471aa81, 32'hc324689d, 32'hc38cfb35},
  {32'hc3ce32a1, 32'hc1fe079f, 32'h4345b91c},
  {32'h446d12d0, 32'h42ed2fa7, 32'h432fce0e},
  {32'hc415b19d, 32'hc2cc5ef4, 32'h42b71d44},
  {32'h45068650, 32'h43831ebd, 32'hc2a8b452},
  {32'hc51322c6, 32'hc2a93884, 32'hc2aad152},
  {32'h449402b7, 32'hc2285fda, 32'h440439b9},
  {32'hc49887d2, 32'h419dfcb9, 32'hc27f76c1},
  {32'h45292cdf, 32'hc338808d, 32'h43affa89},
  {32'hc4e969ff, 32'hc394f376, 32'hc3a0369b},
  {32'h44e819d5, 32'h4379a64a, 32'h42edcdf0},
  {32'hc306c868, 32'hc245493d, 32'hc35a0a06},
  {32'h447b7530, 32'h42748e8b, 32'hc1f3d2e3},
  {32'hc4178b2c, 32'h41b2c9a1, 32'hc38120b6},
  {32'h4480b6a4, 32'h43a4110c, 32'hc2fb89b6},
  {32'hc4b76a78, 32'h40555e68, 32'h42b341f5},
  {32'h452a5b2b, 32'h4240816d, 32'h4367c1e2},
  {32'hc3cdc3bc, 32'hc296a24a, 32'h423dc1e8},
  {32'h44c25caa, 32'hc380bcd7, 32'h42de243c},
  {32'hc446e97f, 32'hc28515be, 32'hc301d5b5},
  {32'h44e706b9, 32'hc39b7179, 32'h4234ca1a},
  {32'hc492b4a3, 32'h435a7128, 32'hc252c97e},
  {32'h44104678, 32'hc31cf67f, 32'hc2b6d32e},
  {32'hc4950b53, 32'h43392297, 32'hc32a4eb6},
  {32'h44b94065, 32'hc2588b09, 32'h42d54f21},
  {32'hc283bde8, 32'h42a6d61f, 32'hc280adec},
  {32'h43e44c83, 32'hc311ff12, 32'h438438aa},
  {32'hc4bea84f, 32'hc31e0a1a, 32'hc32b5e95},
  {32'h4506a587, 32'hc3a35e4e, 32'hc2b46fda},
  {32'hc50dc573, 32'h42861d98, 32'hc1856927},
  {32'h43b4edb0, 32'h43aadc4a, 32'hc2a594fa},
  {32'h41ee6119, 32'h42f7c597, 32'hc3a04ac9},
  {32'h4421dd99, 32'h434783e8, 32'h4375a96a},
  {32'hc5175784, 32'hc364dd1e, 32'h422ae8f1},
  {32'h443a755e, 32'hc30f5fdb, 32'h4378b755},
  {32'hc3b48140, 32'hc1f90a26, 32'hc29601fa},
  {32'h4387fc97, 32'h4372a674, 32'h42bc72a0},
  {32'hc46f3a60, 32'hc2b10505, 32'hc303c0bb},
  {32'h44f522fa, 32'h43676707, 32'h4297de0f},
  {32'hc48c2c33, 32'hc3bd337c, 32'hc35918af},
  {32'h4391f302, 32'hc2ac88b4, 32'h43c43ddd},
  {32'hc400ca14, 32'hc1e116e9, 32'h43d94bf0},
  {32'h450b4b56, 32'h4241b0fe, 32'hc21e2adb},
  {32'hc4bf589a, 32'h42797c6f, 32'hc4022a49},
  {32'h4424b02d, 32'hc3941591, 32'h436c5bf3},
  {32'hc4b669c6, 32'h43aa7d35, 32'h435f7315},
  {32'h45120c0a, 32'hc38514c6, 32'hc2a9ed64},
  {32'hc4f58cdc, 32'hc3274f80, 32'hc1c88fb8},
  {32'h44aa3897, 32'h43288748, 32'h42a10805},
  {32'h4296a052, 32'h432fc36b, 32'hc3582260},
  {32'h4386d788, 32'hc2a9cf10, 32'h435d58df},
  {32'hc47221ac, 32'hc1cfbefe, 32'h410b2118},
  {32'h45095f3a, 32'hc2e6ce88, 32'hc383a325},
  {32'hc34fbbee, 32'h42ba1f9d, 32'hc2abbe76},
  {32'h4492606c, 32'h42dbdffa, 32'hc168c952},
  {32'hc4c5d88d, 32'hc33bdb16, 32'hc34b5bc5},
  {32'hc4264417, 32'hc3bfff9d, 32'hc2ec9ff0},
  {32'h44f39f30, 32'h42cbb462, 32'h42413967},
  {32'hc4974f0a, 32'hc3117176, 32'hc3e4b874},
  {32'h448fe5f7, 32'hc348896e, 32'hc2d16d83},
  {32'hc283af60, 32'h42ef912d, 32'h42b7e22e},
  {32'h44f43707, 32'hc28c3ab1, 32'hc313ff69},
  {32'hc4ef629e, 32'h42a7c1c6, 32'hc302d6f7},
  {32'h44b8a4c0, 32'hc0c59ec6, 32'hc38066f2},
  {32'hc4dfb373, 32'h4229090c, 32'hc2826e29},
  {32'h44966f19, 32'hc3397076, 32'h42ae07e0},
  {32'hc4ec7b7b, 32'h41faacbe, 32'h414e28f8},
  {32'h4373609e, 32'h428f9243, 32'h41f0b396},
  {32'hc4947045, 32'h439d59d0, 32'h436318ba},
  {32'h436d9040, 32'h42cf8a02, 32'hc305ff08},
  {32'hc3f751e0, 32'h42598523, 32'hc40ddb02},
  {32'h4507787a, 32'h42ed0543, 32'h434adaef},
  {32'hc51451df, 32'h41a83cf3, 32'h42e1eac3},
  {32'h44db5b71, 32'hc15e15c6, 32'h42b8b79b},
  {32'hc4b7b2b0, 32'hc38f4a33, 32'hc308b2ce},
  {32'h4502d0a3, 32'h42057b15, 32'h4190a3e2},
  {32'h42662dcc, 32'h440467c5, 32'h405622ed},
  {32'h44bdbbfe, 32'h4200948b, 32'h4363b42a},
  {32'hc4b2cf89, 32'hc3257e3e, 32'hc33575bc},
  {32'h42739060, 32'hc3dea32d, 32'h4391f30c},
  {32'hc52079f3, 32'hc336ecc9, 32'h4319dbd1},
  {32'h4464f58c, 32'h4383739d, 32'h436fef94},
  {32'hc431bb92, 32'h419afba6, 32'h43817b36},
  {32'h44b53de1, 32'hc3422a9a, 32'h42d32e35},
  {32'hc514fdc0, 32'hc3be59f0, 32'hc3829e31},
  {32'h44e34edb, 32'h43b94a0d, 32'h4282689d},
  {32'hc4beff9e, 32'hc1c5d7e4, 32'hc3827855},
  {32'h4513b31e, 32'h4315b408, 32'h439ad415},
  {32'hc483f0a8, 32'hc330182e, 32'hc2ade6b2},
  {32'h440cec57, 32'hc360efd4, 32'h432ada94},
  {32'hc4255636, 32'hc29b092b, 32'hc334240d},
  {32'h43dd09ea, 32'hc12c500a, 32'hc26cff5b},
  {32'hc5131fdc, 32'hc2ee224b, 32'hc37cab28},
  {32'h449716fb, 32'h425f2158, 32'h43cc7be5},
  {32'hc4d41ccd, 32'h434593cb, 32'h42ff0c78},
  {32'h445f5223, 32'hc1926a64, 32'h431fb01a},
  {32'hc297ad20, 32'hc351e699, 32'h42900f7b},
  {32'h43ec4418, 32'hc3ca4f86, 32'h444312b8},
  {32'hc41db8bc, 32'h41dc7c9f, 32'hc398bd45},
  {32'h44dca88d, 32'h433a82b6, 32'hc339897d},
  {32'hc3de7c48, 32'h432c4d44, 32'h41681b14},
  {32'h44b85c01, 32'h41bd50b4, 32'hc1759b15},
  {32'hc45061fa, 32'hc1e9e5b3, 32'h412ce4f2},
  {32'h4484a918, 32'hc1822fb8, 32'hc40ab94b},
  {32'hc337fa8c, 32'h43108242, 32'h430d5d7a},
  {32'h44d15144, 32'h4314be58, 32'h43056ef7},
  {32'hc47631a8, 32'hc3c83597, 32'hc38b6b75},
  {32'h436c6270, 32'hc205c653, 32'h4279199c},
  {32'hc255c240, 32'h43a2c749, 32'hc28b9281},
  {32'h44942918, 32'h431e6728, 32'hc36cbb95},
  {32'hc4c12ab8, 32'h428c7b98, 32'h4315651e},
  {32'h43c45610, 32'hc35af105, 32'hc3c17c65},
  {32'hc4d6cfb7, 32'h41a47a92, 32'hc33705f0},
  {32'h43595020, 32'hc273e583, 32'hc243cf2e},
  {32'hc5036b20, 32'h42b1b844, 32'hc3a38e8d},
  {32'h44308177, 32'hc2f2d499, 32'h4370919e},
  {32'hc4ec8ab6, 32'hc32d7c34, 32'h431c5612},
  {32'h44b6a9d0, 32'hc38b8d36, 32'hc33e0016},
  {32'hc4fbf437, 32'hc352388f, 32'hc2c10852},
  {32'h44474d42, 32'hc33cad7b, 32'hc3214b72},
  {32'hc507db55, 32'h43a09423, 32'h433dda93},
  {32'h449af80c, 32'h4349330b, 32'hc37ae1ca},
  {32'hc4de8659, 32'h434abcb8, 32'h41b3663d},
  {32'h44dc8384, 32'h42be8f55, 32'hc3957bb1},
  {32'hc331f290, 32'h4248a16a, 32'hc2091bb2},
  {32'h44f4a88c, 32'hc2eb2687, 32'h43dca1a5},
  {32'hc49e71bc, 32'hc2e10d24, 32'h431739c4},
  {32'h448b69cb, 32'hc38747bf, 32'h43ad3319},
  {32'h42907c50, 32'h43142994, 32'h4298f5a6},
  {32'h44e50d2d, 32'hc3625b18, 32'h43127966},
  {32'hc32b62ea, 32'h43362188, 32'hc1544fba},
  {32'h44ded175, 32'h439110ef, 32'hc20f4169},
  {32'hc4018266, 32'h41dfb0da, 32'h4379043e},
  {32'h4392b8fe, 32'h43bcac3f, 32'hc1901b7c},
  {32'hc4dc961d, 32'h4306a7a1, 32'h431c633a},
  {32'h41d07800, 32'h424b93a8, 32'h433d7ca1},
  {32'hc4fddc75, 32'hc381aa16, 32'hc28ef065},
  {32'hc3559068, 32'h42cbc264, 32'hc408b702},
  {32'hc417eb40, 32'h433324af, 32'h4333fb1a},
  {32'hc301a488, 32'h41bf3e33, 32'hc1a38a1b},
  {32'hc449f01e, 32'hc2027648, 32'hc1fa3be1},
  {32'h43919598, 32'hc36cc572, 32'h41c09640},
  {32'hc3b37120, 32'hc31a81af, 32'h437890b5},
  {32'h44ecd7f6, 32'h4314efac, 32'hc31b98e5},
  {32'hc31c15e8, 32'h428b712c, 32'h42e3161d},
  {32'h450dd1d4, 32'h43030fd4, 32'hc26f4c8f},
  {32'hc419ea64, 32'h42a3f948, 32'h432ff16e},
  {32'h44747c0e, 32'hc359d9ce, 32'hc31177d3},
  {32'hc3e86eac, 32'hc3c93853, 32'h425d17f7},
  {32'h44b166dc, 32'h4383b937, 32'hc3689dd1},
  {32'hc4a5a6fa, 32'h428b47bc, 32'hc3d42872},
  {32'h44a7b0a0, 32'hc373e4ba, 32'hc0fbab54},
  {32'hc4ee1581, 32'hc33cbee7, 32'hc351afce},
  {32'h42b23062, 32'hc2b768b2, 32'hc32f230f},
  {32'hc441900e, 32'h43552adb, 32'h42d1a622},
  {32'h44c85474, 32'hc4343ce6, 32'h439fbf6e},
  {32'hc40b608d, 32'h4301c8ca, 32'hc3c6827f},
  {32'h42f852f0, 32'h42e7c67e, 32'h4386f15f},
  {32'hc4b9db61, 32'h4324359a, 32'hc32a1735},
  {32'h450c9353, 32'h428656ad, 32'h430c2798},
  {32'hc40521f2, 32'h4313c556, 32'h431afdf2},
  {32'h44a4df4e, 32'hc3023f56, 32'h42f7a990},
  {32'hc4d88a03, 32'h433f42b5, 32'hc3067de3},
  {32'h4441e8bc, 32'h4303254c, 32'hc3901bf2},
  {32'hc4385f7e, 32'hc2a3fadb, 32'hc33ae7d7},
  {32'h44c59f1d, 32'h430fc220, 32'h43e52635},
  {32'hc3dca12c, 32'h4278146e, 32'h41602309},
  {32'h43be4778, 32'h43b9f8bd, 32'h4348d379},
  {32'hc4bd1231, 32'hc384147b, 32'h43857e9e},
  {32'h44a5c0c3, 32'h428e43ba, 32'h43ac9a3a},
  {32'hc4854b6d, 32'h4321ea65, 32'hc33280f5},
  {32'h442fb4f7, 32'h43954eba, 32'hc3ccd37f},
  {32'hc451e9c6, 32'hc34a3dae, 32'h42f57e19},
  {32'h44c933b3, 32'hc2d4a7ae, 32'hc27db033},
  {32'hc43243d0, 32'h4380e93a, 32'h437dfbbb},
  {32'h43e59570, 32'h437e2b42, 32'h43f5d4a7},
  {32'hc466986a, 32'hc21caf25, 32'h4281628d},
  {32'h4452c790, 32'h42f9e7e4, 32'h43b77d77},
  {32'hc42bf7f2, 32'hc2ef0497, 32'hc2b44ec5},
  {32'h44f19888, 32'h4383bff4, 32'h438290d5},
  {32'hc4fb1cd1, 32'h42cf72b5, 32'h435817ed},
  {32'h44a0a46d, 32'h428a4369, 32'h42f786b4},
  {32'hc31580ae, 32'h4351a088, 32'h42d6b9b9},
  {32'h4333600a, 32'h43614253, 32'h432ac8ab},
  {32'hc4362148, 32'hc3d8bca3, 32'hc180ccfe},
  {32'h44fcdaa2, 32'hc238afcf, 32'hc36c9b57},
  {32'hc3d63a68, 32'hc22efe1c, 32'hc313d3dd},
  {32'h44b748be, 32'hc103d601, 32'hc329ff58},
  {32'hc38b412e, 32'hc39bab30, 32'hc2f98093},
  {32'h44339cfe, 32'h427f9346, 32'hc2c0dadd},
  {32'hc41a37c1, 32'hc3445620, 32'h42a76836},
  {32'h4445fed6, 32'h4391090f, 32'h425c3b44},
  {32'hc48bc655, 32'h431ac0e3, 32'h435d73ed},
  {32'h42db2f80, 32'hbee31760, 32'hc3d4e238},
  {32'h43c33309, 32'h438c8f76, 32'hc1be4a54},
  {32'h44be2160, 32'h420dbd74, 32'hc38fe7b5},
  {32'h43882808, 32'hc39b8ee7, 32'h43c8a50c},
  {32'h45204447, 32'hc20e7789, 32'hc2daf221},
  {32'hc345f0c8, 32'h43857c41, 32'hc2881b5a},
  {32'h450c0a0f, 32'hc3377742, 32'h4305e8d4},
  {32'hc48f0502, 32'hc3928508, 32'h4284ce0a},
  {32'h443231dc, 32'hc2990b06, 32'hc3a222b9},
  {32'hc417f5b0, 32'hc0696678, 32'h43159e8c},
  {32'h4435f730, 32'h438be190, 32'hc247a6c2},
  {32'hc30af074, 32'h431f1b7a, 32'h4386272a},
  {32'h44f762af, 32'hc2f17d91, 32'hc3808e6b},
  {32'hc4c14224, 32'hc341c5d4, 32'h4392bf51},
  {32'h44556966, 32'h4289ba17, 32'h438213a5},
  {32'hc4fd3696, 32'hc2a7968e, 32'h43043f46},
  {32'h4483ce43, 32'hc2173d3a, 32'h43c55356},
  {32'hc4f16df3, 32'h429afeac, 32'h424bafe6},
  {32'h43e00ef4, 32'hc3560bce, 32'hc39869a6},
  {32'hc3641b58, 32'h439fcdac, 32'h43556598},
  {32'h4493880b, 32'hc3cb0676, 32'hc392550c},
  {32'hc506b2d4, 32'hc3a86dab, 32'hc371c23c},
  {32'h45070d51, 32'hc2284be6, 32'h42f258fa},
  {32'hc4d7973c, 32'h42fe5765, 32'hc2e4f43a},
  {32'h44a84c37, 32'h426372f4, 32'h42e1bae5},
  {32'hc3856bb8, 32'h42d26282, 32'h42668d4e},
  {32'h43e21b38, 32'h43a7df44, 32'hc3848dd5},
  {32'hc40548de, 32'hc21e9424, 32'h43a92664},
  {32'h450bb851, 32'hc2c8cb15, 32'h4341524b},
  {32'hc4a19f9c, 32'h439dd3e1, 32'h426be225},
  {32'h448cc1e3, 32'h4286cba9, 32'hc2c90f0c},
  {32'h421b3980, 32'hc2840cdd, 32'hc35380cd},
  {32'h44b4cb5d, 32'hc3b2f993, 32'h4413b7fe},
  {32'hc4b5fb86, 32'hc2e1339a, 32'hc2524df6},
  {32'h44e2abfc, 32'h434ffdf8, 32'h4401fa86},
  {32'hc4b936dd, 32'h4377ff5a, 32'hc2fd9137},
  {32'h44828eb3, 32'hc3613ecb, 32'hc401dcf3},
  {32'hc3afc07e, 32'hc1a1060c, 32'hc210d002},
  {32'h44ba4400, 32'hc3727c72, 32'h429967f4},
  {32'hc5028b2a, 32'hc28a9f28, 32'hc310d7a7},
  {32'h450883c1, 32'hc3199ee1, 32'h432fc8bc},
  {32'hc4be9732, 32'h428b3dfe, 32'hc3c1e05e},
  {32'h44b67c27, 32'hc307d96a, 32'h433c0bd0},
  {32'hc483d7f6, 32'hc2bd26de, 32'h43717c34},
  {32'h44424250, 32'h417ae6b2, 32'h4306014c},
  {32'hc3c62af0, 32'hc211eb45, 32'hc11fce9b},
  {32'h44c24fa2, 32'hc243a5a6, 32'h42757c82},
  {32'hc49e24cb, 32'h429fb427, 32'hc37ba516},
  {32'h450685c2, 32'h426b3dda, 32'h43420046},
  {32'hc436f032, 32'h435b4676, 32'h41d51e7e},
  {32'h45193c83, 32'hc36b0a05, 32'hc28ab354},
  {32'h429ff220, 32'h43014f97, 32'hc284e3fc},
  {32'h442cb508, 32'h43d36266, 32'hc18d3a05},
  {32'hc4e26fe6, 32'hc214e841, 32'hc28bc37a},
  {32'h450cacd4, 32'h43312451, 32'h42bd1451},
  {32'hc4acf18c, 32'h43145f2a, 32'h42d2ae60},
  {32'h44bef582, 32'h432de0f3, 32'h42bd7ccd},
  {32'hc3b1f874, 32'h42e48f1d, 32'hc0db0a3b},
  {32'h45163ad3, 32'hc3745b4f, 32'h424d22fd},
  {32'hc4ad895e, 32'hc32f6c5f, 32'h436436b5},
  {32'h43bbec50, 32'hc20b4a28, 32'hc30df887},
  {32'hc3c3e930, 32'hc3e3b9a8, 32'h4374edb3},
  {32'h4346eacc, 32'hc3c05a9b, 32'h439ef803},
  {32'hc3da11c8, 32'hc30f52d6, 32'h4141e538},
  {32'h4435a5a4, 32'h43b6378b, 32'h43d53efc},
  {32'hc4f26960, 32'hc1a9218a, 32'hc29ee9d0},
  {32'h42774a08, 32'hc29b0970, 32'h437c97f5},
  {32'hc5192ca2, 32'h42f374da, 32'h41e657a5},
  {32'h42e59400, 32'hc35aec7c, 32'h43bbc7cb},
  {32'hc45e9174, 32'hc3d9fb6a, 32'h4391999c},
  {32'h43ad8318, 32'hc2150900, 32'h4300ff20},
  {32'hc4b0c9a4, 32'hc3360431, 32'h4337a94b},
  {32'h443af806, 32'h42433143, 32'hc3498bb2},
  {32'hc4c5663e, 32'h4325b24b, 32'hc31d0871},
  {32'h428ef752, 32'hc439ef2a, 32'hc3777810},
  {32'hc3cc2ff8, 32'hc381c395, 32'hc28310e9},
  {32'h439a0440, 32'hc3070042, 32'hc387a52a},
  {32'hc4e62602, 32'h42e01a08, 32'h4407f211},
  {32'h44a6efda, 32'h431e79ac, 32'h436feb3d},
  {32'hc4f87b5c, 32'hc35c9cb9, 32'h42e9e71a},
  {32'h44fd509d, 32'hc2661e67, 32'h424e156d},
  {32'hc411ce0a, 32'hc27334b3, 32'hc314059f},
  {32'h4420b0d8, 32'h42ea68f3, 32'h432d5b90},
  {32'hc4c3d573, 32'hc24470f4, 32'h42f957c1},
  {32'h44da00e6, 32'hc38e6d45, 32'hc2dfc69d},
  {32'hc4f0e615, 32'h433e9af2, 32'h439cd392},
  {32'h44adbf93, 32'h423be498, 32'hc2e2f33c},
  {32'hc429f750, 32'h43b6c29e, 32'h43103af0},
  {32'h4431a5ac, 32'h437a0f92, 32'hc2a322c8},
  {32'hc506c5c8, 32'h42949a2e, 32'hc329215d},
  {32'h445e1a53, 32'h428b7a37, 32'h433c9173},
  {32'hc4fed882, 32'hc232cfda, 32'hc2937b48},
  {32'h429471a0, 32'hc1149330, 32'h43cbb314},
  {32'hc4f2d4f5, 32'h42a86a3d, 32'hc39a30d0},
  {32'h44d2b6b2, 32'hc31a03d3, 32'h4365bf17},
  {32'hc3e75676, 32'h4277faaf, 32'hc3b94630},
  {32'h44660648, 32'h42a3bfc6, 32'hc321d221},
  {32'h42821ae0, 32'h410d6828, 32'h4329388a},
  {32'h441df2fc, 32'hc37c7e60, 32'h44113e90},
  {32'hc4e44e96, 32'h419fcd04, 32'hc387391f},
  {32'h44e45a7b, 32'h3fbeffc1, 32'hc2e8f8b1},
  {32'hc508f8ce, 32'h4234d610, 32'h422a75aa},
  {32'h44799f3a, 32'hc3310793, 32'hc2b3be67},
  {32'hc486c78f, 32'hc3802c19, 32'hc38b22eb},
  {32'h4502145a, 32'h42c6fad2, 32'h431d60ed},
  {32'hc4de7d1a, 32'hc28e5849, 32'hc383e70c},
  {32'h44deea2f, 32'h42a85ee7, 32'hc3c57bff},
  {32'hc43e4307, 32'h434effff, 32'h43bc6c63},
  {32'h45185140, 32'hc343cb20, 32'h43bdd83c},
  {32'hc493b2f4, 32'hc1e71486, 32'hc304c9b8},
  {32'h448e221b, 32'hc43c6e0a, 32'h4300765d},
  {32'hc436a516, 32'h40f410cb, 32'hc1f2f7e3},
  {32'h44233201, 32'hc28b6396, 32'hc39db817},
  {32'hc4dc509a, 32'h42543ccc, 32'h4226e0e8},
  {32'h44ede99d, 32'h43c94fa7, 32'h4333ddcf},
  {32'hc3bd8a32, 32'hc315d370, 32'h4317c915},
  {32'h449bf66a, 32'hc1119ac8, 32'h4315587b},
  {32'hc4eda584, 32'hc2f3dacd, 32'hc3586fd2},
  {32'h4360939a, 32'hc2e55d25, 32'h42690ca8},
  {32'hc4a0dda6, 32'hc2abe3e5, 32'h42e601e4},
  {32'h4482cffd, 32'hc0b8d9a4, 32'h428fc69e},
  {32'hc4c7e6ac, 32'h43a5071e, 32'hc3bb0778},
  {32'h450a90bc, 32'hc2ae5919, 32'h43cdc94b},
  {32'hc4e688e8, 32'hc3b7b2c0, 32'hc2d01e88},
  {32'h44cfb797, 32'hc39b1e90, 32'h42a33997},
  {32'hc3cd8d93, 32'hc38d7967, 32'h43872974},
  {32'h4440dc20, 32'hc382d544, 32'h4365d231},
  {32'hc4d6ceb0, 32'hc2ec115e, 32'h433e9668},
  {32'h4522e70e, 32'hc382c478, 32'h432e2c09},
  {32'hc4c2340d, 32'h42396013, 32'h43e4befb},
  {32'h44d6f487, 32'hc3a2d2d9, 32'hc1660c8d},
  {32'hc44af077, 32'h42aa6c36, 32'hc3aa93a8},
  {32'h448878a3, 32'h43611300, 32'h42591710},
  {32'hc5158d36, 32'hc394fe3f, 32'hc149380f},
  {32'h4494074d, 32'hc38c129c, 32'h41a3f750},
  {32'hc4fa0ec5, 32'hc2e75168, 32'h4299dd8b},
  {32'h431d8d3a, 32'hc3358472, 32'hc33052e8},
  {32'hc47915c8, 32'hc1c4042a, 32'h4286e7df},
  {32'h444c6310, 32'hc281dddb, 32'hc342bd08},
  {32'hc4e79418, 32'h428472a8, 32'h440a6cfb},
  {32'h44ceeaaa, 32'h418a326d, 32'hc2b3caf7},
  {32'hc4d0381e, 32'h4393b77a, 32'hc418193d},
  {32'h449636b8, 32'hc352b9de, 32'h43e038bb},
  {32'hc456711f, 32'hc2f7ef85, 32'hc2d67449},
  {32'h44e25080, 32'hc2ec6d56, 32'hc2ae40d5},
  {32'hc4dde176, 32'h42d7c689, 32'hc0a769cd},
  {32'h44f11afc, 32'hc25648fd, 32'h41566851},
  {32'hc3bc4708, 32'hc2052e03, 32'h436a6efe},
  {32'h43cbad84, 32'h42bf276a, 32'h43727f9c},
  {32'hc497cc9d, 32'h42263f01, 32'hc31b1a28},
  {32'h44f8edec, 32'h431c5970, 32'hc3281f38},
  {32'hc2f12fe0, 32'h42ce5b6f, 32'h43460923},
  {32'h44203db9, 32'hc2932175, 32'hc2f793dd},
  {32'hc4f33d9a, 32'h41d2e6cc, 32'h4229b310},
  {32'h44566e93, 32'hc34e9b93, 32'hc2eca2d8},
  {32'hc50220a4, 32'h434a857b, 32'h42f25708},
  {32'h44fd8915, 32'hc34b8ba0, 32'hc3437564},
  {32'hc45fd3b1, 32'hc2670f76, 32'hc362a33a},
  {32'h4453a56c, 32'h42b5e0b6, 32'h431dcdd3},
  {32'hc51e6aa4, 32'hc2bde228, 32'h42256f7f},
  {32'h43799245, 32'hc1983837, 32'hc26e4619},
  {32'hc40b1640, 32'hc3facdc6, 32'hc29c7265},
  {32'h445f9df8, 32'h436dee9b, 32'h41b5aaf8},
  {32'hc2f79a00, 32'h41a3e5b8, 32'hc35fe257},
  {32'h427cc858, 32'h429effdd, 32'h43d17ca2},
  {32'hc41b3f58, 32'hc18068ba, 32'h42fa68b4},
  {32'h44c8056b, 32'hc37e164b, 32'hc2e275a7},
  {32'hc4af38fe, 32'h4136395a, 32'hc2dde7b6},
  {32'h44b3c9ce, 32'hc361a57a, 32'h420ae54c},
  {32'hc50c19ee, 32'hc39f3a00, 32'h42c95388},
  {32'h450c954a, 32'hc36fa7b9, 32'h431ad47d},
  {32'hc418c03c, 32'hc2be999d, 32'h43438b70},
  {32'h44bf5b9e, 32'h421ac8da, 32'hc3237062},
  {32'hc4abe9a7, 32'hc309e045, 32'h43c22f24},
  {32'h44b829e5, 32'h429c1c88, 32'h43976b5e},
  {32'hc4f9993e, 32'h4385e16a, 32'hc40c31bf},
  {32'h44911cc4, 32'hc2d7d82c, 32'h439a5715},
  {32'hc49437d6, 32'hc2e67cb0, 32'h3f2e95f2},
  {32'h447ea1bc, 32'h42d31028, 32'hc1e1982f},
  {32'hc4de07aa, 32'hc1c0892e, 32'hc3efd5f1},
  {32'h43eaa45c, 32'hc3199221, 32'hc3bc6b9a},
  {32'hc14c175b, 32'h438c549f, 32'h43ccbf88},
  {32'h42ba59ec, 32'h4319cc79, 32'hc222e529},
  {32'hc31a82a0, 32'hc26884be, 32'hc42f0212},
  {32'h43d1a988, 32'h43029b2d, 32'h430fb17c},
  {32'hc50108cc, 32'hc3e65cfa, 32'hc328f86a},
  {32'h437a3b90, 32'hc146a85e, 32'hc3daf832},
  {32'hc50d4f94, 32'hc2ab00e7, 32'h43aabc65},
  {32'h44ed9dba, 32'h42927811, 32'h437a5e4c},
  {32'hc39ebb06, 32'h43837531, 32'hc1b9b479},
  {32'h433fe218, 32'h41fa9d33, 32'h4280e10a},
  {32'hc3d3d970, 32'h42ce075e, 32'hc37b486f},
  {32'h44fae672, 32'hc38e1039, 32'h422d6740},
  {32'hc2447b20, 32'hc30b3445, 32'h43d8bd8d},
  {32'h452b5a98, 32'h4421f640, 32'h4264ce23},
  {32'hc3aa69d8, 32'hc2257cf0, 32'h42106170},
  {32'h44890726, 32'hc32b22fe, 32'hc18d5cca},
  {32'hc4e4cd3e, 32'h42987a16, 32'hc2b46b50},
  {32'h44330ae8, 32'h439c02a5, 32'hc36fd538},
  {32'hc2e44c00, 32'h43327f6a, 32'hc12b817c},
  {32'h44fe2d38, 32'hc2d63462, 32'h42699980},
  {32'hc4ba74c9, 32'hc1b5aafa, 32'h43bc544c},
  {32'h44931a3e, 32'hc2c03132, 32'h4391a154},
  {32'hc2c0f4da, 32'hc363adcf, 32'h41106f93},
  {32'h448357da, 32'h424d2f80, 32'hc3857898},
  {32'hc4f5b613, 32'h430c80ef, 32'hc0189d88},
  {32'h44a612f2, 32'h432ce7ca, 32'h42ea13a1},
  {32'hc3d41770, 32'h43e6e40b, 32'hc10323c3},
  {32'h44be123a, 32'hc261b8f4, 32'hc3e37b36},
  {32'hc5038c1e, 32'hc27d1623, 32'hc305f6be},
  {32'h4450f59c, 32'h431f1702, 32'h422e9aa6},
  {32'hc4dedf1f, 32'hc305bb8a, 32'h4351462f},
  {32'h43a416f8, 32'h4305bd2b, 32'hc335845c},
  {32'hc41e1923, 32'hc26727cb, 32'h438ef739},
  {32'h43bc48a8, 32'hc33cce97, 32'h42bf1c42},
  {32'hc3950b58, 32'h430a1150, 32'h430f53cf},
  {32'h444d242c, 32'h41cbe2e6, 32'h4115abe8},
  {32'hc3906410, 32'h434332bf, 32'h42399af4},
  {32'h4442925d, 32'hc38ad2a6, 32'h425062c9},
  {32'hc4e77814, 32'h4288b464, 32'hc337b672},
  {32'h443ac1c0, 32'hc32191b4, 32'h43222b5e},
  {32'hc4a4f3e4, 32'h42bbf45f, 32'hc193afe1},
  {32'h442d15cc, 32'hc312d4fd, 32'hc3e89f05},
  {32'hc40036ba, 32'hc2feb52b, 32'hc28fc5f1},
  {32'h44cb02dc, 32'h43947611, 32'hc294eaaa},
  {32'hc4f92baa, 32'hc3220c64, 32'h43a02875},
  {32'h44345700, 32'h431385b8, 32'h445534aa},
  {32'hc44461e9, 32'hc31ac420, 32'hc3fce92f},
  {32'h4402ea17, 32'h41e1d387, 32'hc30cf3e4},
  {32'hc4ade2d2, 32'hc3cd41eb, 32'hc2923423},
  {32'h451adf70, 32'hc3a7cfa6, 32'h4198d34c},
  {32'hc510d08e, 32'h42089ff0, 32'h4392866e},
  {32'h44d456ae, 32'hc2845c5c, 32'h419caa04},
  {32'hc50ae987, 32'h42947246, 32'h43d3cfd0},
  {32'h44a5d350, 32'h429c7654, 32'hc2f3e915},
  {32'hc4e00e50, 32'hc324aefe, 32'hc3479098},
  {32'h43fdf310, 32'h433227de, 32'hc36e24ce},
  {32'hc2cc0830, 32'hc38d9cb8, 32'h42d6a30a},
  {32'h4484332e, 32'h4244cad1, 32'hc22c2faa},
  {32'hc4746b7e, 32'h438a0ae4, 32'h43304fcd},
  {32'h4416c3fc, 32'h4339b7e6, 32'hc3b31e5d},
  {32'hc4e63985, 32'hc2186833, 32'h42e6b834},
  {32'h4359fb69, 32'h4310bc53, 32'hc32ee964},
  {32'hc4eb7b06, 32'hc25a7119, 32'h4385780f},
  {32'h4482d0ba, 32'h42873e2d, 32'hc29a0f0b},
  {32'hc4095a6a, 32'hc1814f87, 32'hc4047b53},
  {32'h44f16b46, 32'hc3c9f7e6, 32'h424e5a3e},
  {32'hc2440c40, 32'h42fbf5ac, 32'h428bc8fc},
  {32'h44a02554, 32'h421ac98c, 32'hc33fe986},
  {32'hc4e9eabd, 32'hc327d9fc, 32'h41b92ec8},
  {32'h449d8a52, 32'hc2e91859, 32'hc34049b5},
  {32'hc3cad138, 32'h435602a5, 32'h4411166a},
  {32'h44b972f0, 32'hc19dee88, 32'hc40d5195},
  {32'hc5056db3, 32'h4139f15e, 32'h423ca7d0},
  {32'h44bd8704, 32'hc3b853ad, 32'hc3312e12},
  {32'hc4936bd3, 32'hc242ef0a, 32'h4265e4b9},
  {32'h45127f37, 32'hc4259b4f, 32'h429e195f},
  {32'hc3abd958, 32'h4152968c, 32'hc3275b11},
  {32'h44330b80, 32'h430d5cbd, 32'hc307f2b0},
  {32'hc434e6dc, 32'hc297491c, 32'hc185fbde},
  {32'h44376600, 32'h428b642b, 32'h434359c8},
  {32'hc398a5f0, 32'h42e997ce, 32'h43935890},
  {32'h44898ace, 32'hc36df4e6, 32'hc2fdc092},
  {32'hc48b4564, 32'hc3747e3e, 32'h432bb19a},
  {32'h44f0dd05, 32'h4347a3e2, 32'h418d31e0},
  {32'hc3b44ed0, 32'hc2343848, 32'h42366722},
  {32'h44e74f08, 32'h4382e5b2, 32'hc3b36b82},
  {32'hc475c34a, 32'h4272160e, 32'hc29e759a},
  {32'h4508e1b6, 32'h41de5db8, 32'h43cad26b},
  {32'hc48d2a9c, 32'h43b0c712, 32'hc2388d0a},
  {32'h449f7c41, 32'h425e43ca, 32'hc34df4f9},
  {32'hc3df4a6e, 32'hc27e77f9, 32'h441429c8},
  {32'h4464147c, 32'hc31ce27f, 32'hc31fbc9b},
  {32'hc486c78b, 32'h4336d6d8, 32'h43758c61},
  {32'h449113f7, 32'hc28ed5aa, 32'h42951951},
  {32'hc38c992f, 32'h439064a6, 32'hc317f26c},
  {32'h439ddf02, 32'h424a6fc4, 32'hc30e4ade},
  {32'hc5093511, 32'hc31d57b0, 32'h4310e2fb},
  {32'h43bce4fc, 32'h4271a6ee, 32'h4244804a},
  {32'hc483d1c3, 32'h4350d8c2, 32'h44035a31},
  {32'h44833a67, 32'h42fc4472, 32'hc1beaeda},
  {32'hc519806b, 32'hc2fd47fe, 32'h43808b82},
  {32'h4443cec2, 32'hc4116fbc, 32'hc4157023},
  {32'hc4843c2d, 32'hc3525a52, 32'h4352c901},
  {32'h44f9cd96, 32'hc31117f6, 32'h437e7be4},
  {32'hc503822b, 32'hc3f0c74f, 32'h439b3451},
  {32'h450ba429, 32'h42b14681, 32'h42d73738},
  {32'hc2f42e00, 32'hc1fd2099, 32'h43eeadd3},
  {32'h45002728, 32'hc0830a49, 32'hc2f95b7a},
  {32'hc441f63c, 32'hc32321fa, 32'h43330b1e},
  {32'h450bd1ad, 32'h42f98bc7, 32'hc22e9b16},
  {32'hc4e960c7, 32'hc3196246, 32'h42c014c7},
  {32'h44968295, 32'hc35f7d64, 32'h416d9cc9},
  {32'hc4d5d26e, 32'h428e1723, 32'hc31fc938},
  {32'h4506b64c, 32'hc4026325, 32'hc39346ab},
  {32'h448cd01b, 32'h43833f6d, 32'hc3194b4c},
  {32'hc43024ce, 32'hc415cc10, 32'hc0f05abc},
  {32'h43ef4c40, 32'h43b7f2bb, 32'hc40feaaf},
  {32'hc31df676, 32'hc39962d1, 32'h4301e8eb},
  {32'h44e08aa8, 32'hc4139552, 32'h4309e927},
  {32'hc44295b9, 32'h43323888, 32'hc351cd20},
  {32'h44d5ed0e, 32'h429ee413, 32'hc34d2010},
  {32'hc4aa519c, 32'h4291c263, 32'h42c1dcc6},
  {32'h42cec1d0, 32'h4331de75, 32'hc386c0b6},
  {32'hc4069e00, 32'hc2505442, 32'hc2bbbfb6},
  {32'h44bea724, 32'h43b5ceb4, 32'hc34a6946},
  {32'hc396523c, 32'hc29b1c04, 32'h40c19914},
  {32'h44882962, 32'hc3ad6c14, 32'h42b8906c},
  {32'hc4fd03a3, 32'h43e0a363, 32'hc39272f4},
  {32'h4463519c, 32'h438f4b97, 32'h4187f957},
  {32'hc51a5347, 32'h40f5d0fa, 32'hc3199d0d},
  {32'h43a88c70, 32'h438c13c2, 32'h43a476da},
  {32'hc199bbc0, 32'h42be148d, 32'h42ffcee1},
  {32'h43fc2e6e, 32'hc2e2a17e, 32'hc2c2d307},
  {32'hc506627c, 32'hc1b72f51, 32'h42ac9100},
  {32'h44fc5235, 32'hc2ecb21b, 32'hc34fbd88},
  {32'hc3ca4000, 32'hc31450a2, 32'hc3411692},
  {32'h440bc665, 32'h42f7a7e8, 32'hc30988bf},
  {32'hc4206d14, 32'h4190e4fc, 32'h42a3c088},
  {32'h43f4d6c6, 32'h430d22c1, 32'hc3b05c36},
  {32'hc4c7c425, 32'h43364aae, 32'h435dde89},
  {32'h44942b8f, 32'hc39ad1bf, 32'h41715c22},
  {32'h43929e58, 32'h43402e7b, 32'h43627edb},
  {32'h437ff011, 32'h42d3ffae, 32'hc39292bc},
  {32'hc50167a5, 32'h4367061d, 32'h4339b983},
  {32'h44b75441, 32'h425ec4ad, 32'hc176f2f6},
  {32'hc330b320, 32'hc32ed13e, 32'h42f593b4},
  {32'h44c6d62d, 32'h42c5a5ff, 32'hc3e5acb2},
  {32'hc2877815, 32'hc1e58a04, 32'h430e2b4e},
  {32'h44def5af, 32'h43d86ca0, 32'hc37cd986},
  {32'hc43581d4, 32'hc3838e1a, 32'h42d5cdd3},
  {32'h45165428, 32'hc1e7b85c, 32'h41cb65cc},
  {32'hc3bf64a0, 32'hc2e16c42, 32'h4400e22a},
  {32'h44f5e014, 32'hc403465f, 32'h438d709f},
  {32'hc4fbe775, 32'hc190e017, 32'h43375540},
  {32'h44e8e234, 32'hc06f13a0, 32'h43a21ef4},
  {32'hc3c541a0, 32'h42e34896, 32'hc38d61ba},
  {32'h44ac08c5, 32'hc280a066, 32'h43d3f93d},
  {32'hc4b418ae, 32'hc2dff9b6, 32'hc20d7058},
  {32'hc1386b00, 32'h41ef57b3, 32'h44055b84},
  {32'hc206ee80, 32'h429b23f2, 32'h43b0dd27},
  {32'h44be9b4d, 32'h43c39758, 32'h42bcf31d},
  {32'hc4400254, 32'h434de7cb, 32'h432cb97c},
  {32'h4448154a, 32'h43857146, 32'h425cdf0b},
  {32'hc42634e6, 32'h41da92d8, 32'h431a6170},
  {32'h448a9a4d, 32'hc2aed2c9, 32'h4257bdc4},
  {32'hc4b20fd5, 32'hc29844b3, 32'h43100c92},
  {32'h44c08429, 32'hc2a1d883, 32'hc314f29c},
  {32'hc46e0621, 32'h41abcb31, 32'h3fbb67d3},
  {32'h4423ba94, 32'hc36bae68, 32'h42882c0d},
  {32'hc3259020, 32'hc3040b6e, 32'hc39435a8},
  {32'h44d2ff2b, 32'hc2a43613, 32'hc0d2a564},
  {32'hc504abad, 32'hc35427d0, 32'hc3886df0},
  {32'h448b2a99, 32'hc226f46a, 32'h4255f726},
  {32'hc366dac1, 32'hc4090cdf, 32'h42877f3b},
  {32'h4485b321, 32'hc40493bc, 32'hc221de7d},
  {32'hc398f9c2, 32'hc32a9b4f, 32'hc378e62e},
  {32'h438986c8, 32'h43003d11, 32'h434034ec},
  {32'hc50510f9, 32'hc36854ee, 32'h42181a7b},
  {32'h442be2dc, 32'hc344e660, 32'hc2362384},
  {32'hc501b56e, 32'hc2d72ced, 32'h42e6e02b},
  {32'h44a0c910, 32'hc353bc8e, 32'hc37dc6c5},
  {32'hc4a83b0b, 32'hc2e1dff6, 32'h4042fd6a},
  {32'h44a5e838, 32'h42ce99cf, 32'h43892e65},
  {32'hc4844abf, 32'hc3bc4277, 32'hc3a1e201},
  {32'h451bc07c, 32'h42d603a0, 32'h43ca8810},
  {32'hc41336b4, 32'hc0e7b6a8, 32'hc29e5688},
  {32'h44738501, 32'hc38b3f6e, 32'hc27186e6},
  {32'hc5120ba4, 32'hc355b9ec, 32'h42c226ae},
  {32'h43aef6b4, 32'h4383432e, 32'hc3091f76},
  {32'hc4c13f3c, 32'h42ab7af2, 32'h4212d866},
  {32'h43a7d43c, 32'hc24395d6, 32'hc1140f1a},
  {32'hc45a7102, 32'h4326f641, 32'h4347d195},
  {32'h43acf418, 32'h429c38e9, 32'h40b2ddf8},
  {32'hc31bec10, 32'hc339b97f, 32'h4348941c},
  {32'h451ca38f, 32'hc2f823bc, 32'h430247bb},
  {32'hc5049f08, 32'hc3247c44, 32'hc0bcf999},
  {32'h44149eb9, 32'h41dbaf36, 32'hbe42c380},
  {32'hc51abcc9, 32'h4354fc17, 32'hc3218655},
  {32'h449cc0fa, 32'h43400771, 32'h4257d3de},
  {32'hc43c83ce, 32'hc1198260, 32'hc36eb4f3},
  {32'h44f47e7c, 32'h42978fd2, 32'hc3a4e37a},
  {32'hc4a7a8fd, 32'hc2f030c2, 32'hc38135e7},
  {32'h451fd35c, 32'hc36743be, 32'hc28d6f50},
  {32'hc511950e, 32'h435e95e3, 32'hc3816303},
  {32'h440d894b, 32'hc36947a1, 32'h4394f311},
  {32'hc45a02dc, 32'hc1e8a83c, 32'h434f5c57},
  {32'h45158922, 32'h4302ba35, 32'h430946ed},
  {32'hc51297e9, 32'hc28ea95d, 32'hc1e0018e},
  {32'h4494fe40, 32'hc0520d86, 32'hc08a876c},
  {32'hc4363177, 32'hc2079292, 32'h43e38167},
  {32'h43e9e420, 32'h42976a93, 32'h43e996d7},
  {32'hc5045c3e, 32'hc369c1c3, 32'hc365bf2d},
  {32'h44a984d2, 32'h428e2d9e, 32'h43083045},
  {32'hc4f84dfd, 32'h434888e6, 32'hc3693946},
  {32'h43b92264, 32'hc3159801, 32'hc3aea972},
  {32'h438b8549, 32'hc203743f, 32'hc1a768f3},
  {32'h4469dca0, 32'h43adf9d7, 32'h435c9a9b},
  {32'hc477247a, 32'hc3275848, 32'hc1b5d9af},
  {32'h44661478, 32'hc227d866, 32'h432799eb},
  {32'hc497441e, 32'h43107dfc, 32'hc306f7f3},
  {32'h44df3a82, 32'h417e2fca, 32'hc363fcf3},
  {32'hc4915287, 32'hc27d1387, 32'h43afd15a},
  {32'h44c8b8f8, 32'hc1a48a6e, 32'hc28c651c},
  {32'hc4965c89, 32'hc2d26902, 32'hc34712b0},
  {32'h443298be, 32'hc31e16da, 32'h42354001},
  {32'hc4a6643f, 32'h4379e73f, 32'h437ae31d},
  {32'h443aff40, 32'hc35ef44c, 32'hc2a20462},
  {32'hc401f072, 32'h438e5d71, 32'hc365ad5d},
  {32'h44d534a1, 32'hc2eb4fc6, 32'h43de6ea1},
  {32'hc4918899, 32'h415038aa, 32'h419ce728},
  {32'h44bbd397, 32'hc3a653fa, 32'h430f7029},
  {32'hc43686c5, 32'h43446001, 32'h4346b517},
  {32'h45137ba4, 32'hc410b5c3, 32'h4318c2bb},
  {32'hc4b70855, 32'hc3596912, 32'hc23405f0},
  {32'h449e1001, 32'hc20f1b13, 32'h42d3a274},
  {32'hc492c8b0, 32'hc3664ec2, 32'h43ca495c},
  {32'h44c15111, 32'h42a8c14f, 32'h43626f5c},
  {32'hc2d0b6b0, 32'hc31168de, 32'h422bc9f4},
  {32'h43e1a7ec, 32'h436d8f52, 32'h43c5c3d2},
  {32'hc4b211fa, 32'h41fb7a84, 32'h4301bb7e},
  {32'h44c412da, 32'h40984014, 32'hc1fcbd26},
  {32'hc4ce5b5b, 32'hc385298e, 32'h41f9972e},
  {32'h4504373d, 32'hc2a3212c, 32'hc2ed6deb},
  {32'hc4d47ceb, 32'h43706cd5, 32'h43800d71},
  {32'h44cce9a6, 32'hc38cbba8, 32'h440b5519},
  {32'hc4993c04, 32'h43e2deff, 32'h42b9eb8a},
  {32'h44919c72, 32'h42f1b9d7, 32'h4333b380},
  {32'hc41cd574, 32'hc3203692, 32'hc3bb649b},
  {32'h450906ac, 32'hc2f71f40, 32'hc33724e9},
  {32'hc5183f54, 32'hc3460e6f, 32'h427c0e3c},
  {32'h44a48172, 32'h43929616, 32'h4327043e},
  {32'hc2d4bd80, 32'h42a3e57b, 32'h43cc35ab},
  {32'h44b41dc7, 32'h42df492d, 32'hc295d19c},
  {32'hc4d31510, 32'h413fa915, 32'h43115d5a},
  {32'h44624b31, 32'h4304b1a3, 32'hc342b1d8},
  {32'hc4837676, 32'h4327af44, 32'hc35729cf},
  {32'h44fa95ac, 32'h432b9b8d, 32'h42307b95},
  {32'hc40a53a0, 32'hc39799ca, 32'hc1e1ef86},
  {32'h44dd1052, 32'h4372fcaf, 32'hc2ea6e64},
  {32'hc4deab62, 32'h3fd88962, 32'hc1cf81a6},
  {32'h444fc093, 32'h42af2c53, 32'hc36f9019},
  {32'hc49f2e9a, 32'hc2707f8e, 32'hc2f2ff4d},
  {32'h44e5e3d2, 32'hc28b6165, 32'h41032330},
  {32'hc425d421, 32'hc26a3147, 32'h43667838},
  {32'h44e20428, 32'h4254d750, 32'hc3ce2826},
  {32'hc43b6cbb, 32'h43561e07, 32'hc2b2d6de},
  {32'h448b333e, 32'hc3653aa1, 32'h428dc271},
  {32'hc3258f90, 32'h425097d4, 32'h428ac70e},
  {32'h4500a9bc, 32'h43690a60, 32'hc1404562},
  {32'h41eab108, 32'hc1aa4e44, 32'h4317af48},
  {32'h45155866, 32'hc2c6f365, 32'hc33a94da},
  {32'hc50225f7, 32'hc2964092, 32'h41e8ba27},
  {32'h45024f60, 32'h43784c79, 32'hc367e6c1},
  {32'hc5114f06, 32'h43a51933, 32'hc303ea98},
  {32'h4492f710, 32'hc12ac218, 32'h43ab0f6b},
  {32'hc4e493d9, 32'h436b10f5, 32'hc27d4f0b},
  {32'h44b72c37, 32'hc3423009, 32'h4140e912},
  {32'hc4fe4d3a, 32'hc3c55896, 32'h425f8403},
  {32'h449eac94, 32'hc281242e, 32'hc31e26b3},
  {32'hc4675a2a, 32'hc3b9571e, 32'h41ff7923},
  {32'h42921622, 32'hc38409be, 32'h42e89ac7},
  {32'hc48a1a55, 32'h43f4534b, 32'hc3255137},
  {32'h44a84a1e, 32'h410defa3, 32'h4357e2b8},
  {32'hc50e5266, 32'h426b8550, 32'hc2145764},
  {32'h44b9dabf, 32'hc1af2532, 32'h431500a7},
  {32'hc4faa519, 32'h42db7f9f, 32'h40a1b6b7},
  {32'h44404284, 32'hc2c752c9, 32'hc29fda91},
  {32'hc400928c, 32'hc3738576, 32'hc2e2596b},
  {32'h449f8732, 32'hc32ef78c, 32'hc309fca3},
  {32'hc4eb0658, 32'h43361049, 32'hc3e67c3c},
  {32'h432039f0, 32'hc1f6f815, 32'h4313aca8},
  {32'hc39282a8, 32'hc1a447a0, 32'hc328f336},
  {32'h441a47f4, 32'h43acb121, 32'hc310840d},
  {32'hc41e5313, 32'hc3f4a6c7, 32'h42fec6aa},
  {32'h44ccddaf, 32'h4326cab3, 32'h42b169f6},
  {32'hc438313d, 32'hc39da678, 32'h4261740d},
  {32'h44b8b93e, 32'h432e557b, 32'hc33eb168},
  {32'hc4a10981, 32'hc29acb00, 32'hc2910863},
  {32'h4514d3d8, 32'h43024d6f, 32'hc2a44fc1},
  {32'hc43ec0e1, 32'h423ab6f4, 32'h43153d2b},
  {32'h43a6e2b8, 32'h43408fd8, 32'hc3e8f428},
  {32'hc502663d, 32'h435ceb5b, 32'hc2be5e0c},
  {32'h44b9c144, 32'h43b18fbe, 32'hc2955096},
  {32'hc443900a, 32'hc1823c25, 32'h43f38fa9},
  {32'h43e94398, 32'h42756374, 32'hc30aea4c},
  {32'hc393a1a2, 32'hc307e710, 32'hc3fc07f6},
  {32'h4433d5d8, 32'h42195394, 32'hc108f013},
  {32'hc4c1c31a, 32'hc2d02863, 32'h42ad3de9},
  {32'h44fcdebf, 32'hc301938a, 32'h431dd57c},
  {32'hc48c000d, 32'hc0af5a28, 32'h43c27449},
  {32'h448af5a1, 32'h4183dfc0, 32'hc31f7ac1},
  {32'hc496c4b0, 32'h43113bfa, 32'h426eee6f},
  {32'h43901f33, 32'hc29bdd6f, 32'h42a6e7b2},
  {32'hc41bf306, 32'h438f5b91, 32'h438fef54},
  {32'h44b464c2, 32'hc2f92ac1, 32'h42b4351a},
  {32'hc5043ee7, 32'hc117d056, 32'h43e206cf},
  {32'h449f4cdd, 32'h4346ddcd, 32'hc296fe99},
  {32'hc40fc164, 32'h43842f76, 32'hbfe60a20},
  {32'h44da4356, 32'h439c4cd1, 32'hc1444fb1},
  {32'hc31f7448, 32'hc301f5bb, 32'h434ae820},
  {32'h43230614, 32'h41f71f89, 32'h42d51a77},
  {32'hc4c0f3ee, 32'hc35f846e, 32'hc3d86be4},
  {32'h450e175f, 32'h439d989b, 32'h419814b2},
  {32'hc38406c8, 32'h4187fc28, 32'h432a8157},
  {32'h437f3c70, 32'h43e2b24c, 32'hc31f2ba2},
  {32'hc256e1a0, 32'hc3150995, 32'hc38ae999},
  {32'h4368fc30, 32'h43b0b95f, 32'h43868df0},
  {32'hc5120294, 32'hc2f6f5d8, 32'hc353bc86},
  {32'h44bb13ce, 32'h42a44124, 32'h43013fa0},
  {32'hc4178a3b, 32'hc3f920c3, 32'hc2ac4dae},
  {32'h43f6a7cb, 32'hc39b35b7, 32'h42a3a3cc},
  {32'hc4921ed8, 32'h43723631, 32'hc283be76},
  {32'h44aea233, 32'hc0c88614, 32'h42e5f41c},
  {32'hc3f3740e, 32'h40d4b502, 32'h432dc570},
  {32'h44e9b42c, 32'hc33e037b, 32'hc2856fde},
  {32'hc4a2d4f0, 32'h43a5f7c9, 32'h425095f4},
  {32'h43e0b826, 32'h43098435, 32'hc2c8f264},
  {32'hc4d995bf, 32'hc2fa24d6, 32'h4318870e},
  {32'h449e8d3b, 32'hc38e452c, 32'hc4058ae4},
  {32'hc484904b, 32'h435ea3fa, 32'hc2d35121},
  {32'h44d768e4, 32'hc304fd31, 32'hc128d78a},
  {32'hc475777b, 32'h42eb6002, 32'h429684c9},
  {32'h4496508f, 32'hc2b93818, 32'hc321a91d},
  {32'hc4819472, 32'hc322d807, 32'hc385f959},
  {32'h43c281ae, 32'hc26e8e7f, 32'h42f8e52d},
  {32'hc5110987, 32'h43961b45, 32'hc316aeb8},
  {32'h43effe08, 32'h4370ace8, 32'hc21b24de},
  {32'hc3d220bc, 32'hc2c3678a, 32'hc18b434d},
  {32'h444120f8, 32'h4295450b, 32'hc3c84427},
  {32'hc3b9c53b, 32'h423de18c, 32'hc3a290f7},
  {32'h45148470, 32'hc2e4118f, 32'hc304f6ee},
  {32'hc403c33e, 32'hc1f8d441, 32'h43580e98},
  {32'h450dc7d2, 32'hc396b5e8, 32'h43494b91},
  {32'hc4274e2d, 32'h4275b231, 32'h42624cba},
  {32'h450a28a6, 32'h43e3ebd1, 32'hc36ced23},
  {32'hc497e031, 32'h42eeb199, 32'h43b8b692},
  {32'h43af2a88, 32'h43913912, 32'hc326d2a1},
  {32'hc38f66bc, 32'hc293b83d, 32'h43020f2e},
  {32'h44d4c3ce, 32'hc35a4c11, 32'h434a4f2c},
  {32'hc4fd7fcd, 32'hc2eb86f5, 32'h4378d9c1},
  {32'h44ddb02e, 32'h42bc058a, 32'h432b5d0a},
  {32'hc4095e05, 32'h4196e45a, 32'h42697437},
  {32'h4514dbc9, 32'hc325dcb5, 32'h43583a4d},
  {32'hc3722a38, 32'hc3eed3f5, 32'h4240daf7},
  {32'h44d89fb6, 32'hc2b9efa5, 32'h436e0b58},
  {32'hc430bb5c, 32'hc2e56c0a, 32'h4395958c},
  {32'h45161ecd, 32'h41e187e7, 32'h42ffb7ca},
  {32'hc480fb5a, 32'h41a1e2a4, 32'h4219bf3c},
  {32'h44160624, 32'h432104a1, 32'hc303e92a},
  {32'hc4ab503c, 32'h41ce2885, 32'hc347feb6},
  {32'h4511d492, 32'hc3a34390, 32'hc2a20a9c},
  {32'hc487f15a, 32'hc21a546d, 32'h4397bcda},
  {32'h444548b6, 32'h439cff22, 32'hc2ba9f2f},
  {32'hc4fe0925, 32'hc2440069, 32'h42df758d},
  {32'hc1564340, 32'h439f9847, 32'hc2442714},
  {32'hc425e546, 32'hc2598eed, 32'h426f2093},
  {32'h44034f57, 32'h43090232, 32'h41e75ded},
  {32'hc50108d2, 32'hc202af57, 32'h41ed930d},
  {32'h4441d2a8, 32'hc13e9556, 32'h4318c59d},
  {32'hc513246a, 32'hc2bc3ab6, 32'h43901ab4},
  {32'h44787592, 32'h431790e4, 32'hc397dd8c},
  {32'h424965b6, 32'h41d0b05d, 32'hc12071e4},
  {32'h4505836c, 32'hc344638b, 32'hc34dce38},
  {32'hc469f669, 32'h42b9ebd1, 32'h43a69ced},
  {32'h4488ad2a, 32'hc164f0ce, 32'hc29f55a1},
  {32'hc430ade8, 32'h43a43000, 32'h429721ae},
  {32'h4492f10e, 32'hc20e40c8, 32'hc2ef43c7},
  {32'hc2c687ea, 32'h43daaab6, 32'h43a0cb47},
  {32'h43ef0c96, 32'hc1ab6f60, 32'hc3aaf3e6},
  {32'hc4435534, 32'hc3c00727, 32'hc1f8cb6e},
  {32'h44444c47, 32'hc2a7e19f, 32'hc2bd9a22},
  {32'hc4a6ea57, 32'hc25e0d9f, 32'h4331a78c},
  {32'h43c323f8, 32'hc26b5c89, 32'h435db4ac},
  {32'h4347e128, 32'hc3b291f0, 32'h43981e5b},
  {32'h44f84ac3, 32'hc3a3210b, 32'hc3981393},
  {32'hc49e302c, 32'hc14405ee, 32'hc12fdc7e},
  {32'h44d3c59a, 32'h42efc2d3, 32'h4355ebba},
  {32'hc395105e, 32'h4310d112, 32'hc27fe986},
  {32'h449b8a3f, 32'hc349d424, 32'h42de7ce8},
  {32'hc35079e8, 32'h432066ee, 32'h43b9e3b2},
  {32'h44646c14, 32'hc37d4344, 32'hc316b619},
  {32'hc42bf5e9, 32'hc368ca4b, 32'hc2de9318},
  {32'h44f86933, 32'h431ce05c, 32'h4329c42c},
  {32'hc49eabf5, 32'hc2ff7ca2, 32'hc34d343c},
  {32'h44a50df2, 32'h42e00c71, 32'h43870e33},
  {32'hc3c12f3f, 32'hc35fe71e, 32'hc165ea10},
  {32'h44a35d1f, 32'hc31c9f76, 32'h438317fd},
  {32'hc4f16d96, 32'h428fa529, 32'hc2ca5044},
  {32'h449a2760, 32'h43758a39, 32'h418f357a},
  {32'hc4bc3633, 32'h41974f6e, 32'h434e5f7b},
  {32'h4511820e, 32'h42892d6f, 32'h43ee841e},
  {32'hc41fbb34, 32'h42196351, 32'hc33c2442},
  {32'h44e0c053, 32'h419d518f, 32'h422c938e},
  {32'hc4eaae99, 32'h42976406, 32'h438fb7a3},
  {32'h44993d1a, 32'hc3e7b870, 32'hc1033629},
  {32'hc4b3dd66, 32'hc39692bc, 32'h43937772},
  {32'h44a82cc0, 32'h428486b8, 32'h43c532b3},
  {32'hc4f2fa1f, 32'hc2f4e184, 32'hc305e2c0},
  {32'h44a22555, 32'hc3485367, 32'hc380f9d4},
  {32'hc4fb80e5, 32'hc35fba1e, 32'h43a09f1c},
  {32'h44c3d5ef, 32'hc34bd6b7, 32'h419089f1},
  {32'hc5139344, 32'h42290efb, 32'hc335b944},
  {32'h44b5423a, 32'hc3516932, 32'h4396250a},
  {32'hc4806cdf, 32'hc2f99b41, 32'h41e18f7c},
  {32'h44da8276, 32'hc394b8b4, 32'hc20da587},
  {32'hc42fcbba, 32'h42b7597a, 32'h42201c1e},
  {32'h4504edf0, 32'h430c2923, 32'h43636c95},
  {32'hc49b24f1, 32'hc2948783, 32'hc1efe3e6},
  {32'h4515655c, 32'hc39bd6f6, 32'h431890b6},
  {32'hc44510de, 32'hc2af77f9, 32'h4366bee4},
  {32'h44b0aef8, 32'hc36ba053, 32'hc14a2fe3},
  {32'hc496f8e4, 32'h439461f6, 32'h430f8f3e},
  {32'h44fff16f, 32'hc24a99c6, 32'hc2b47393},
  {32'hc48d4965, 32'hc3295ae5, 32'hc31e7db2},
  {32'h44ccf7c5, 32'hc24df40c, 32'h41fa2e1f},
  {32'hc4a0f066, 32'hc32cc94d, 32'hc310668c},
  {32'h44875489, 32'h40e3de16, 32'hc2fa8166},
  {32'h41221d6a, 32'hc3ff927a, 32'hc3399781},
  {32'h450cba02, 32'hc2c19a1f, 32'hc37dc55f},
  {32'hc50b8161, 32'h438680b7, 32'hc39dd620},
  {32'h44edc8fe, 32'h439fdeae, 32'hc2c97fe3},
  {32'hc4224f8f, 32'hc1814018, 32'h43164d94},
  {32'h44ed3f6c, 32'h4342f18b, 32'h436148cd},
  {32'hc50829c4, 32'hc10695f8, 32'hc1abab92},
  {32'h451586fe, 32'h431b8f5d, 32'h4372598d},
  {32'hc42373ed, 32'h43b5b094, 32'h43586864},
  {32'h446d7062, 32'hc1368c2d, 32'hc343b221},
  {32'hc4d98eac, 32'hc32f0b6d, 32'hc39ef734},
  {32'h44c329d6, 32'hc2c73141, 32'hc2b6f092},
  {32'hc49ff316, 32'h42c0678f, 32'hc2b3e411},
  {32'h43502ab0, 32'h43d40cb8, 32'hc2c44b04},
  {32'hc1067f00, 32'h430133d6, 32'hc3925e9a},
  {32'h44f4443e, 32'h42fbbba9, 32'h42d0c62d},
  {32'h43974951, 32'hc31d2df0, 32'hc0ab9dcc},
  {32'h450e6598, 32'hc1504593, 32'hc287d3f6},
  {32'hc4aef414, 32'h43b78d1c, 32'hc3f277b9},
  {32'h420c6b30, 32'hc3cab5ba, 32'h43a6af1c},
  {32'hc39a9868, 32'h436b164c, 32'hc15deef5},
  {32'h44afee2e, 32'h42e40182, 32'h41b6c88d},
  {32'hc50832e0, 32'hc3a3371f, 32'hc3207889},
  {32'h446ea108, 32'hc30734b6, 32'h438793c8},
  {32'hc4d34ece, 32'h43d35bf6, 32'h43a7f37d},
  {32'h44f16fcb, 32'h43a31182, 32'hc386d8b9},
  {32'hc4a3fbda, 32'hc33a1eaa, 32'hc38a49d1},
  {32'h44b0e254, 32'h42dbe758, 32'h43dcfdf4},
  {32'hc4e74226, 32'h4317f2be, 32'hc28383d1},
  {32'h450129ca, 32'hc3475248, 32'h430f26f2},
  {32'hc402b9c8, 32'h4367c4c9, 32'h41f662cb},
  {32'h4444664a, 32'h408b2981, 32'hc3a746fa},
  {32'hc40e95b2, 32'hc298c1c2, 32'hc2041dd8},
  {32'h44b3431a, 32'hc383875e, 32'hc1be87c7},
  {32'hc4a05bd8, 32'h41ed8791, 32'h44050f1c},
  {32'h44fc1204, 32'h433a3db3, 32'h43c588af},
  {32'hc4db828e, 32'h4073a2d8, 32'h42562e95},
  {32'h44965da8, 32'h42f71dc5, 32'h42e9254e},
  {32'hc3e6f7a7, 32'hc3346e24, 32'hc37a3b34},
  {32'h44c06caa, 32'hc39062bb, 32'hc33ac6ff},
  {32'hc4d64bfc, 32'hc30828f8, 32'h43db4e08},
  {32'h4519f17f, 32'h43b1740e, 32'h4366daad},
  {32'hc3a864fc, 32'h4185b6a3, 32'hc3120a66},
  {32'h4522a605, 32'hc2a1877d, 32'hc05f9a48},
  {32'hc43b603b, 32'h437d81e2, 32'h43388d24},
  {32'h45216b81, 32'hc323a2a3, 32'hc3933bf1},
  {32'hc4e16502, 32'hc35bf047, 32'hc2509dba},
  {32'h43a44fc0, 32'h40ab7722, 32'hc2df74a8},
  {32'hc50acc5d, 32'hc33cc274, 32'h423fa818},
  {32'h44a5423e, 32'h431c679c, 32'h4369f50b},
  {32'hc3f7c5d4, 32'hc2eb03e6, 32'h428c5a6e},
  {32'h44923d83, 32'hc2dfd42c, 32'h43430fee},
  {32'hc356c0d8, 32'hc3b9326d, 32'hc2f4efb8},
  {32'h44800527, 32'hc27caa19, 32'h4351da09},
  {32'hc3780374, 32'h42c04e14, 32'hc2c79b4b},
  {32'h450a75c5, 32'h4281d5d7, 32'h43af1702},
  {32'hc46ba085, 32'hc0ef43b5, 32'h42770627},
  {32'h44b49960, 32'h4396a09f, 32'h42e1fb38},
  {32'hc328c8ee, 32'h438dfdb2, 32'hc33eae37},
  {32'h45137d0c, 32'hc26b13fa, 32'h434aea9c},
  {32'hc448a05a, 32'h4264c691, 32'hc3660b97},
  {32'h4457e6b6, 32'h43b4082c, 32'hc1d61dd3},
  {32'hc45a936a, 32'hc3a64440, 32'h43efae4c},
  {32'h44f8ea7c, 32'h4298e354, 32'hc2a7126c},
  {32'hc4918c2e, 32'hc1c0a03a, 32'h42a26d04},
  {32'h4469b778, 32'hc36d8e60, 32'h4142fae0},
  {32'hc493cd74, 32'h436c5a57, 32'hc339a5cb},
  {32'h42099c28, 32'h43691dd9, 32'hc2fe1cee},
  {32'hc49f8eea, 32'hc3aa722e, 32'hc3392312},
  {32'h449a39bb, 32'hc21742c7, 32'hc306d4fb},
  {32'hc4e7533f, 32'h40a1cdda, 32'h439c91f0},
  {32'h4501287b, 32'h4314bd50, 32'h439b1dd8},
  {32'hc50cc34a, 32'h4118b4b7, 32'h4379cebc},
  {32'hc38e5a5b, 32'h4283f8bc, 32'hc2d060c2},
  {32'hc505ad1e, 32'hc1c93fb7, 32'hc31ddb5a},
  {32'h4507107f, 32'h3f3b8e4a, 32'hc31eb4e4},
  {32'hc44b4be8, 32'hc2bb3a57, 32'hc327c3ad},
  {32'h43061d02, 32'hc393a012, 32'h43ac437d},
  {32'hc4b4ccf8, 32'h42c92f73, 32'hc3be6690},
  {32'h41e6e480, 32'hc3978068, 32'h4431d742},
  {32'hc4d26b07, 32'h41726d78, 32'hc3c4907f},
  {32'h45203c76, 32'h42c7295f, 32'h42a036e6},
  {32'hc501837e, 32'h422754b4, 32'hc310a865},
  {32'h43719328, 32'h439a92f0, 32'hc35406b9},
  {32'hc4b2b4ea, 32'h42aaf6f6, 32'h4232f75c},
  {32'h4501bce1, 32'h43512d0d, 32'hbf9f39ce},
  {32'hc50c89a1, 32'hc386c499, 32'hc3109611},
  {32'h44a98f9a, 32'hc2c6046b, 32'h432bbea6},
  {32'hc3e08d00, 32'hc25d47d6, 32'h43636e63},
  {32'h44588777, 32'hc3a6cd88, 32'h437a80e3},
  {32'h4112f300, 32'hc32a03d0, 32'hc16cece4},
  {32'h44504b8e, 32'hc1bc75f7, 32'h41c1ee68},
  {32'hc4e91d5a, 32'h42dd1227, 32'hc339cfa4},
  {32'h43f9ad3c, 32'h437f7473, 32'h421e2fab},
  {32'hc28e0fdd, 32'hc029924b, 32'h436dc307},
  {32'h44e33908, 32'h41814361, 32'hc38d71ed},
  {32'hc43d613b, 32'hc3eb52fc, 32'hc2cc04bf},
  {32'h44f83b3f, 32'hc31ce34e, 32'h423d3fb1},
  {32'hc4f895b6, 32'h42f3b6e7, 32'hc22962f2},
  {32'h448f57b5, 32'h406115d3, 32'h419f2941},
  {32'hc4038a10, 32'hc1f862dc, 32'hc3917115},
  {32'h45061659, 32'h42aa61cf, 32'h43244de0},
  {32'hc50f8afc, 32'h41c55676, 32'h43bb9f98},
  {32'h3fb4d400, 32'hc231a1c5, 32'h4409bc1d},
  {32'hc4c53201, 32'h42b92c1c, 32'hc33f8f6a},
  {32'h4403014a, 32'hc39346f4, 32'h43a8cd7c},
  {32'hc383f488, 32'h438f7e15, 32'hc2d565e9},
  {32'h449cd96f, 32'h4153c139, 32'h4320cf09},
  {32'hc4d1bc9d, 32'hc23251e7, 32'hc1dd2f74},
  {32'hc460098e, 32'h423d2b5b, 32'hc391fb98},
  {32'h44cff286, 32'h426ae258, 32'h41b4900b},
  {32'hc4e71cfc, 32'hc077c85b, 32'hc26da397},
  {32'h43c54b6c, 32'hc345da01, 32'hc35847dc},
  {32'hc40d9a04, 32'hc22b4e31, 32'hc31f78b4},
  {32'h44cb5a28, 32'h426799ed, 32'hc353329c},
  {32'hc4f2c405, 32'h4413111f, 32'hc279dc3a},
  {32'h44bca0d3, 32'hc20395d5, 32'h43523fea},
  {32'hc4334c44, 32'h41ea8ee9, 32'hc2dc0620},
  {32'h43fb26de, 32'hc3a3a1bc, 32'h42494439},
  {32'hc4a0b4d0, 32'hc3a9ee9e, 32'hc41822b3},
  {32'h4510f5d1, 32'hc2b03c18, 32'hc29e02ca},
  {32'hc31a9900, 32'hc291e386, 32'hc384c1e8},
  {32'h43e6a593, 32'h428d79cf, 32'hc3c8e296},
  {32'hc504a13e, 32'hc3c0e669, 32'hc2842b30},
  {32'h45050bbc, 32'h43dff0f7, 32'hc37168b6},
  {32'hc4b56e30, 32'hc2027e73, 32'hc15e1e4e},
  {32'h449e8ef4, 32'h42c70bde, 32'h431ef11f},
  {32'hc4d6c890, 32'hc2965422, 32'h42981036},
  {32'h42278090, 32'h43a17fcf, 32'hc213b6a9},
  {32'hc3aa6f00, 32'hc342c3bb, 32'hc3c9fac5},
  {32'h4373677f, 32'hc3260e79, 32'hc2f23d97},
  {32'hc45cbee8, 32'hc3911794, 32'hc16eeafc},
  {32'h43c1fbe0, 32'hc3937930, 32'h42f53b33},
  {32'hc500a2f3, 32'h4318e1e8, 32'hc3793da2},
  {32'h44a1db30, 32'hc3db0b5f, 32'h41fd9e4e},
  {32'hc47a86c3, 32'hc253673c, 32'hc396e94e},
  {32'h4492d634, 32'h435af77a, 32'h43b424fb},
  {32'hc50725b6, 32'hc259545e, 32'hc3938d73},
  {32'h44f18ff8, 32'hc0a0a7a0, 32'hc31d4cb7},
  {32'hc40d4452, 32'h43297d26, 32'hc2e506c0},
  {32'h44e79b5e, 32'hc3b6cb31, 32'hc3c7c329},
  {32'hc49c8642, 32'hc3343f2e, 32'h43886282},
  {32'h44e04ba4, 32'h433c5b30, 32'h438286a9},
  {32'hc5088681, 32'h4029c982, 32'hc39fc7ed},
  {32'h44dce48a, 32'hc36e2426, 32'hbe3150a0},
  {32'hc4b20516, 32'hc352ca5f, 32'hc3e15b2e},
  {32'h44e7ff93, 32'hc187f19f, 32'hc0f8fcdf},
  {32'hc4c05f23, 32'hc37a734e, 32'h43852c5a},
  {32'h45131687, 32'h41d26eac, 32'h4402fc51},
  {32'hc486a8b0, 32'hc232afc5, 32'hc2673057},
  {32'h4460b911, 32'h43534cda, 32'h43765f4c},
  {32'hc3e89550, 32'hc3330c1f, 32'hc2a372ee},
  {32'h44c33b36, 32'hc41df810, 32'h43ad230f},
  {32'hc488ea06, 32'h440bb4fa, 32'h40a02de1},
  {32'h426ac740, 32'h43252d06, 32'hc3486db4},
  {32'hc4fb39c4, 32'h422a5078, 32'hc0294d08},
  {32'h43f021e9, 32'h437d321c, 32'h43640fae},
  {32'hc3cdef34, 32'h437e2ebd, 32'hc2c235b9},
  {32'h44e26f6f, 32'hc34c12d6, 32'hc09800c8},
  {32'hc417f86e, 32'h43f320d2, 32'h43c1e06a},
  {32'h43c1c458, 32'hc29a2736, 32'hc2cdf926},
  {32'hc4995509, 32'hc32b7ca4, 32'hc2b623cc},
  {32'hc3ae46dc, 32'hc3b0b1cb, 32'h43665934},
  {32'hc2ac9a97, 32'hc3832cc5, 32'hc3b2cf2c},
  {32'h431fd660, 32'hc394df07, 32'hc42fe1e0},
  {32'hc3ec8fdf, 32'hc1c807a8, 32'h42d74b88},
  {32'h44c7170a, 32'hc288e675, 32'h42c777d5},
  {32'hc4554a0a, 32'h42a7f1b0, 32'hc3bd19ab},
  {32'h4317b19e, 32'hc38ac055, 32'hc33d19de},
  {32'hc2b485e0, 32'hc3a20f71, 32'hc38ae070},
  {32'h4498d514, 32'hc2b278bb, 32'hc3721aa0},
  {32'hc48b8674, 32'h42f76aa4, 32'h3f0a073e},
  {32'h44010146, 32'h4325656d, 32'h431dae9d},
  {32'hc44b6a92, 32'hc325115b, 32'h439b2d89},
  {32'h447a2d36, 32'hc11a2592, 32'hc1c468be},
  {32'hc50cc23c, 32'hc1a22ea2, 32'hc14901d3},
  {32'h438556cc, 32'h43a28dc3, 32'h42fd968e},
  {32'hc4d91006, 32'hc3207efc, 32'hc3b4c363},
  {32'h439ba05c, 32'h43362a47, 32'hc3d811bc},
  {32'hc5065fc4, 32'hc3781a1d, 32'h438ed02a},
  {32'hc3477530, 32'hc33f4420, 32'h439179ad},
  {32'hc50873fe, 32'hc3d09cb0, 32'h438ab84b},
  {32'h45115f0c, 32'hc3978b4d, 32'hc38af8b7},
  {32'hc49a9e59, 32'hc2d37504, 32'h42e2d284},
  {32'h45122d74, 32'h43435b6d, 32'hc04da11c},
  {32'hc4cf7d4f, 32'hc2c94f10, 32'hc322470d},
  {32'h44bf489a, 32'hc3038195, 32'hc2cc72a1},
  {32'hc443234a, 32'h43b702fa, 32'h433b7ae7},
  {32'h4447e2cc, 32'hc3ababfa, 32'hc3a0951b},
  {32'hc503b04a, 32'h43187e52, 32'hc34cc8a8},
  {32'h443961db, 32'h4309c807, 32'hc409d263},
  {32'hc482caac, 32'h43105c44, 32'h43322cfb},
  {32'h450397ae, 32'h4296326f, 32'hc35c52a8},
  {32'hc3a40be0, 32'hc191b85a, 32'hc2d98238},
  {32'h44acef32, 32'hc395789e, 32'h439033f9},
  {32'h4414f927, 32'h43c7f910, 32'hc3c7b997},
  {32'h44949762, 32'hc18d5eec, 32'hc308fb0c},
  {32'hc341bb70, 32'h432ff33b, 32'h42ca8275},
  {32'h41c05b78, 32'h4345f9ef, 32'hc2ed66f8},
  {32'hc4d6cd30, 32'h42b3ab61, 32'hc34e7bda},
  {32'h41a1e480, 32'hc3848024, 32'h43481334},
  {32'hc3cdc4da, 32'hc2bba1ae, 32'hc33896a0},
  {32'h44255538, 32'hc3b9cc43, 32'hc182003b},
  {32'hc4bb7bb3, 32'h420578de, 32'hc284a8a4},
  {32'h45067421, 32'h4363a626, 32'hc2c2e92f},
  {32'hc507a538, 32'hc1c35db6, 32'hc2eca85f},
  {32'h44ee1c20, 32'hc32c733c, 32'h43428332},
  {32'hc4469441, 32'hc3f35c49, 32'h43afc1fb},
  {32'h4535136a, 32'h4282b7f1, 32'h42e23886},
  {32'hc3cd5792, 32'h434c5593, 32'hc0f98046},
  {32'h43ab942a, 32'h41d1ce45, 32'h42a1c2aa},
  {32'hc4d9f241, 32'hc3a1e3d0, 32'h42c0b507},
  {32'h44973355, 32'hc26253a3, 32'hc3468580},
  {32'hc0576b20, 32'h4314eb6a, 32'h44016af3},
  {32'h44cbbdcf, 32'h439d540e, 32'hc3200ed4},
  {32'hc40610bd, 32'hc2892a6d, 32'hc37d6909},
  {32'hc20265f0, 32'hc37ee7c8, 32'h42907cb8},
  {32'hc4802d18, 32'hc14e1c45, 32'hc2a1e224},
  {32'h43a56243, 32'h43918b04, 32'h4331299a},
  {32'hc455d24b, 32'hc4082b02, 32'h43aeb6d8},
  {32'h42b555f4, 32'h4257f6d7, 32'hc3b66d28},
  {32'hc49a0dba, 32'hc0d86f0e, 32'h43ebd0c5},
  {32'h42ce28cb, 32'h42c7d5ae, 32'h4285ff13},
  {32'hc4ba83da, 32'hc2f11c6b, 32'h43cfb468},
  {32'hc32e1120, 32'h432624b0, 32'hbfea48c8},
  {32'hc509748c, 32'hc317f9c2, 32'h42fbd6d4},
  {32'h450ade82, 32'h4198642e, 32'hc30cb726},
  {32'hc5130136, 32'h438f5b0e, 32'hc28d7f5f},
  {32'h44860ee0, 32'h422c0ebe, 32'hc2bd7e93},
  {32'hc408ca44, 32'hc3a0331e, 32'h4372c0e4},
  {32'h45106fb0, 32'h42955616, 32'hc284486b},
  {32'hc490c224, 32'h43cc912a, 32'h424f08a1},
  {32'h44688178, 32'hc3a72e04, 32'hc31bf9e5},
  {32'hc4e6a4fe, 32'hc136f43f, 32'hbf7719b4},
  {32'h44b63fec, 32'hc33b6805, 32'h43753b22},
  {32'hc51da389, 32'hc3089446, 32'hc308b09a},
  {32'h43d4cc5d, 32'hc3c8fe4f, 32'h4286efeb},
  {32'hc4fc9bc3, 32'hc2dc9454, 32'hc27a8b60},
  {32'hc3876584, 32'h43b91244, 32'h43b36b97},
  {32'hc4715bf5, 32'h431a8395, 32'h438b0bc8},
  {32'h44f7be40, 32'hc37823c4, 32'h433105b2},
  {32'hc3f076a2, 32'h3f05632d, 32'h43055a17},
  {32'h44ea3d03, 32'h430039c0, 32'h42b5c428},
  {32'hc4816739, 32'h43f2085b, 32'h430b5eef},
  {32'h44fe0793, 32'hc1b737d7, 32'hc3743810},
  {32'hc50a3200, 32'h43b9b025, 32'hc28fc929},
  {32'h449ae6ed, 32'hc37f7acf, 32'hc3c327f9},
  {32'hc48fd540, 32'hc38a48f3, 32'h429e156c},
  {32'h44aadf84, 32'h439593ed, 32'hc375ace6},
  {32'hc4d48f1a, 32'h430caa22, 32'hc3773f8b},
  {32'h443cad60, 32'hc2d42b2a, 32'hc37df144},
  {32'hc4d27e14, 32'hc2213d8a, 32'hc1a8226b},
  {32'h44c1a8b0, 32'hc3d5bb90, 32'h42683f1f},
  {32'hc4f4b16c, 32'hc20fda68, 32'hc2ec569f},
  {32'h448ea986, 32'hc338d78b, 32'hc3fc66e0},
  {32'hc359e4f0, 32'hc23836a3, 32'h41b0ef3f},
  {32'h4508b632, 32'h417807aa, 32'hc356c649},
  {32'hc3fa80f4, 32'hc3c38763, 32'hc1cb2530},
  {32'h42726d90, 32'hc363d94c, 32'hc33fe7b2},
  {32'hc445016e, 32'h4359fb14, 32'hc238eba8},
  {32'h446c2841, 32'hc386a727, 32'h43cbd9c7},
  {32'hc46f4672, 32'hc102e4e1, 32'hc3a39b9e},
  {32'h43f9060a, 32'hc294020f, 32'h43b29d61},
  {32'hc4b645f6, 32'h42feaaf4, 32'h4326c8b0},
  {32'h4491dac3, 32'hc124c1a0, 32'hc27e29ca},
  {32'hc4c8f036, 32'hc34c0e68, 32'hc212fd1a},
  {32'h4274a8a0, 32'hc34f4d3d, 32'h439bed8b},
  {32'hc09e0d00, 32'h430beb39, 32'hc3407464},
  {32'h43d2f3d2, 32'hc2e03ac3, 32'h439a254b},
  {32'hc2996320, 32'h42316b91, 32'h43d52bc7},
  {32'h450b82de, 32'h42e3ff04, 32'h42ca5073},
  {32'hc2e8c3a0, 32'h43d5c174, 32'h43768722},
  {32'h44fd9c68, 32'h4373b99c, 32'hc1c8438a},
  {32'hc442ec3e, 32'hc3baf71d, 32'hc345172b},
  {32'h4480b454, 32'hc33cfbf2, 32'hc1a9e984},
  {32'hc4c18105, 32'h43478c4b, 32'h43845240},
  {32'h44e2d432, 32'hc30af0f1, 32'hc353d529},
  {32'hc43e8d7c, 32'h42eee34f, 32'h4327b24c},
  {32'h4461b978, 32'h4365f9da, 32'h4408e33b},
  {32'hc3325a6e, 32'hc2d79c9c, 32'h4341f542},
  {32'h448ac496, 32'h43af612d, 32'hc2b754be},
  {32'hc48ca344, 32'h432558cd, 32'h3fff1882},
  {32'h4435002c, 32'hc2bdbd5f, 32'h43a86ddb},
  {32'hc44a0990, 32'hc2ac15f2, 32'hc233904a},
  {32'h431fb6ae, 32'h43cb7cf2, 32'hc38ea5c6},
  {32'hc4ca346a, 32'h43710780, 32'hc30bd473},
  {32'h446508a6, 32'hc1c209c5, 32'hc328d075},
  {32'h43fdf2d6, 32'hc3c70ad9, 32'hc3f2e962},
  {32'h44f651da, 32'hc2c82dec, 32'hc28a5c70},
  {32'hc4f2cbd8, 32'h42d97afa, 32'hc35ea1a2},
  {32'h44ddaf78, 32'hc3985fbb, 32'hc342c447},
  {32'hc3792cf8, 32'hc2efea7e, 32'h43a64476},
  {32'h44cce658, 32'h431e3678, 32'hc310b702},
  {32'hc3e08f4c, 32'hc318290a, 32'hc119c2a8},
  {32'h44e5757a, 32'h40e8b012, 32'h43a4d21c},
  {32'hc4e65a8c, 32'h438998fd, 32'hc3390684},
  {32'h4518b6ab, 32'h43f8ea7e, 32'hc2721e5a},
  {32'hc4fe5dd9, 32'hc25bcf24, 32'hc3477ec4},
  {32'h44d68d87, 32'h42ade802, 32'hc39efc29},
  {32'hc4eabc2a, 32'hc3e67abf, 32'hc2dc6b7a},
  {32'h44f734ed, 32'h41c1a0e8, 32'h4386eb45},
  {32'hc385955a, 32'hc3a96fc1, 32'h41f68f92},
  {32'h4502213c, 32'hc3033cb3, 32'h433fe182},
  {32'hc48f8222, 32'hc2f906b1, 32'hc31f45e8},
  {32'h447f2d77, 32'h42d4e372, 32'hc3e7475f},
  {32'hc4f1dddc, 32'h441ce74c, 32'h42d2142c},
  {32'h4478063c, 32'h43360cb9, 32'h42db07ca},
  {32'hc50146bb, 32'hc3630de6, 32'hc277c352},
  {32'h44bff1b0, 32'h41a26d92, 32'h42c4f567},
  {32'hc4e3292a, 32'hc3a57b54, 32'hc317b932},
  {32'h44a0cc3d, 32'hc1fe67ef, 32'h4241c0b1},
  {32'hc3c3f9bf, 32'hc2eb343f, 32'hc2dee7c4},
  {32'h434a0640, 32'hc28bbc4f, 32'h42e3665e},
  {32'hc4f0f032, 32'hc1a08a3e, 32'h43243949},
  {32'h4498e43d, 32'h41d4fee6, 32'h42d676e8},
  {32'hc4847ba1, 32'hc2b1322a, 32'hc2b2e384},
  {32'h43eb83c2, 32'hc3caacbd, 32'h434d7530},
  {32'hc49c83b1, 32'h42954b2f, 32'hc337195e},
  {32'h427dce80, 32'h4263f44f, 32'hc38a8a57},
  {32'hc4b4aabd, 32'hc3f94bd3, 32'hc2880ad4},
  {32'h44987828, 32'h432c5b87, 32'hc3a5083c},
  {32'hc4a06a1e, 32'h43c174d1, 32'h43acff00},
  {32'h4480e9b3, 32'hc340678b, 32'h3f7684c0},
  {32'hc4b3ad0d, 32'hc2334d3c, 32'hc2d19612},
  {32'h440265e8, 32'h42935d54, 32'h43c2b51d},
  {32'hc4fcafe7, 32'hc34136da, 32'hc34a2ca6},
  {32'h43d6f38b, 32'h440ddf57, 32'hc29257bb},
  {32'hc4dd191b, 32'h43333c1c, 32'h421b5cc3},
  {32'h44bbb028, 32'hc43c69c7, 32'h4388e30c},
  {32'hc4e1d64d, 32'h422cfb53, 32'h439335fa},
  {32'h4501cf31, 32'h43a356a0, 32'h43980c58},
  {32'hc437b680, 32'h4389b60e, 32'hc3a3feaa},
  {32'h4487451c, 32'h4304aba1, 32'hc372d043},
  {32'hc473041c, 32'h437dcc48, 32'hc3486c04},
  {32'h4442c205, 32'hc38a8f33, 32'h429d32df},
  {32'hc5047b6a, 32'hc3a76c5f, 32'h42a2dd30},
  {32'h4490925c, 32'h43305e2e, 32'h42f52104},
  {32'hc3c08ebb, 32'hc369956e, 32'hc3100e08},
  {32'h440a251a, 32'h43fa382c, 32'hc1fc448d},
  {32'hc502ab11, 32'hc3c7b027, 32'hc2f269fa},
  {32'h44aba0a4, 32'hc31ff266, 32'h430cae80},
  {32'hc3f73236, 32'h42b2473a, 32'hc38955c6},
  {32'h44f21463, 32'h43a1ce4e, 32'hc3777861},
  {32'hc4e35e3f, 32'hc38006ee, 32'hc291108f},
  {32'h44baeab3, 32'hc148b88c, 32'hc31687d6},
  {32'hc339c9a0, 32'hc3aa5468, 32'hc2b0f35b},
  {32'h44d57640, 32'h439f22e3, 32'h4310b724},
  {32'hc49c0078, 32'hc2eb192a, 32'hc30139ed},
  {32'h44095ffc, 32'hc3da56cf, 32'h43e7b858},
  {32'hc3d94390, 32'h43c73192, 32'hc30b19d5},
  {32'h450286e6, 32'h4384b36f, 32'hc2cf9ff5},
  {32'hc48c47dd, 32'hc34a6f99, 32'hc22cd8d7},
  {32'h44be4fda, 32'h42faca9c, 32'hc2e1356d},
  {32'hc477e71e, 32'hc2c4f407, 32'hc36e1740},
  {32'h450f993b, 32'hc3261d19, 32'hc2be6890},
  {32'hc435b338, 32'h40811ac8, 32'hc39be61a},
  {32'h42e36390, 32'hc3027dc2, 32'h44004486},
  {32'hc406bbf0, 32'h434e1dec, 32'h43325ff9},
  {32'h44e9e50e, 32'h43848d4d, 32'hc3c9eff7},
  {32'hc4d15aea, 32'hc34a7dda, 32'h43b29de7},
  {32'h4412a472, 32'h4370e9f7, 32'hc3993662},
  {32'hc3eb0dec, 32'h431e905a, 32'h42a5c30c},
  {32'h44a76ce1, 32'hc31c222e, 32'h438a082b},
  {32'hc501f31b, 32'hc3f8fe6c, 32'h438f5b7b},
  {32'h44c7decc, 32'h426af7e2, 32'hc202cb3f},
  {32'hc45b8200, 32'hc388969b, 32'h430f8bab},
  {32'h44f0fb1e, 32'hc2af3938, 32'h429d95c4},
  {32'hc3a00f74, 32'h4343b964, 32'hc341f0df},
  {32'h44c1ce8a, 32'h42dd9d52, 32'hc30c57dc},
  {32'hc4ed6a4c, 32'hc33dd2ad, 32'h4367c9d4},
  {32'h430a3db0, 32'hc2804ca3, 32'hc3273faa},
  {32'hc3d84888, 32'hc1077190, 32'hc1199641},
  {32'h451293c5, 32'hc3039c28, 32'h420f543b},
  {32'hc3c2cfd2, 32'hc319adb9, 32'hc0bdd472},
  {32'h44e65dcc, 32'hc30ab1b2, 32'h42fb29e9},
  {32'hc4f08a2d, 32'h431e466b, 32'h435c1699},
  {32'h4506f904, 32'h407d565d, 32'h429650a4},
  {32'hc4c9609d, 32'hc3031f71, 32'hc3814d2b},
  {32'h447aa125, 32'h42d87b49, 32'hc2662caf},
  {32'hc4ed18d1, 32'hc1119818, 32'h436f9caf},
  {32'h44daf7fc, 32'hc2bf1d07, 32'h43e0c1b1},
  {32'hc47ffb36, 32'hc2c5029e, 32'hc26837b9},
  {32'h447b7448, 32'h43772428, 32'hc33d2b1b},
  {32'hc4c7baba, 32'hc3a9407c, 32'hc3f20534},
  {32'h450c2020, 32'h4285acb0, 32'hc1d16c72},
  {32'hc4a27d14, 32'h43918d5c, 32'hc38843f4},
  {32'h444ab529, 32'h433d1756, 32'h3f00f875},
  {32'hc36593e5, 32'h429fc433, 32'h4388847b},
  {32'h434730a8, 32'h42c84703, 32'hc2618333},
  {32'hc484a18f, 32'h4313c6ca, 32'hc3af2307},
  {32'h44cfc1ab, 32'h434f7e8d, 32'hc381dd88},
  {32'hc3d29ef2, 32'hc31a4163, 32'hc362f711},
  {32'h44d55fad, 32'hc31869a6, 32'h424c3648},
  {32'hc49b53ff, 32'h43ef70fa, 32'h4320c23c},
  {32'h4501af34, 32'hc27c8e18, 32'h437e43fe},
  {32'hc3eecfa0, 32'h42849ca7, 32'h42f0038c},
  {32'h44e889e4, 32'h43141cfd, 32'hc2dad254},
  {32'hc4ed820f, 32'hc1a1c61d, 32'hc32f7ef0},
  {32'h449c19b4, 32'hc2c69685, 32'hc3164a06},
  {32'hc4385fb8, 32'h4374ceb0, 32'hc3f041f7},
  {32'h446d65d4, 32'h43ea270b, 32'h3f43e661},
  {32'hc48411c0, 32'hc3668ff6, 32'hc3a19afe},
  {32'h44c5553f, 32'hc2a45122, 32'h43697b02},
  {32'hc3e236a0, 32'hc388edae, 32'hc2c95453},
  {32'hc2f2e030, 32'h439fa6d3, 32'hc2a88fa7},
  {32'hc47d8fe0, 32'h438fd4ef, 32'h43902030},
  {32'h44a1b8e3, 32'h43c65d10, 32'h43b0a05c},
  {32'hc4d27ce8, 32'h432d9423, 32'h43846396},
  {32'h43e06fb8, 32'hc2fa84c1, 32'h42a9f8b2},
  {32'hc4f85922, 32'h43668f92, 32'hc3445359},
  {32'h43968c44, 32'h4300682a, 32'hc2a151b6},
  {32'hc5154e35, 32'hc339956d, 32'hc3292ec8},
  {32'h44327e68, 32'h4394ee80, 32'hc2b79127},
  {32'hc4cf0a06, 32'h4343ad42, 32'h4171b946},
  {32'h4511c60c, 32'h43cd2a73, 32'hc25a0eef},
  {32'hc4a18ad3, 32'h42c1c982, 32'h42d34d5c},
  {32'h445a5038, 32'h438c4556, 32'h40ccb4f0},
  {32'hc4d0e629, 32'hc3916472, 32'hc3477001},
  {32'h43d9befe, 32'h42a494cc, 32'h42d319f5},
  {32'hc50c6feb, 32'h43eec143, 32'hc33669bb},
  {32'h4044b400, 32'hc35f1459, 32'hc28e34ec},
  {32'hc4cc4da9, 32'h434cc2a2, 32'hc34ec622},
  {32'h44c93483, 32'hc2472539, 32'hc1c21972},
  {32'hc4feb30a, 32'h424ce394, 32'hc27cebee},
  {32'h43e4af6c, 32'hc3813581, 32'hc2868fed},
  {32'hc5006947, 32'h43845473, 32'h42ef8100},
  {32'h44b2095d, 32'hc1b4ffbd, 32'h4373558d},
  {32'hc512a038, 32'hc2a6910f, 32'h422b4139},
  {32'h449c0608, 32'h435c0fd0, 32'h42c12dfc},
  {32'hc3a40758, 32'h42c069f1, 32'h43d23414},
  {32'h445306b0, 32'hc369ac7e, 32'h440216f0},
  {32'hc50cd64e, 32'h43d52016, 32'h4202e1f6},
  {32'h4268ae30, 32'hc29d2e88, 32'h409f2590},
  {32'hc3bd72f8, 32'hc41199a3, 32'hc32dfbbc},
  {32'h4444a444, 32'hc383f5d2, 32'h42baf2df},
  {32'hc4969b7e, 32'hc3f3dc29, 32'h43d564ab},
  {32'h4514395e, 32'h437ed4cf, 32'h440585fa},
  {32'hc49b3da1, 32'hc3748482, 32'h437a2350},
  {32'h450b5ee0, 32'hc313a98c, 32'hc39b7ce4},
  {32'hc4cccb36, 32'h4388a0dd, 32'hc2f85279},
  {32'h4489becd, 32'hc2aff284, 32'h43f7d89d},
  {32'hc3b82749, 32'hc2207643, 32'h43a43598},
  {32'h4385f935, 32'h43896411, 32'h405be70d},
  {32'hc50c342c, 32'hc244724b, 32'hc37b82c8},
  {32'h450dd488, 32'h40e7cfdc, 32'h43c1e48f},
  {32'hc4942205, 32'h439501de, 32'hc3202668},
  {32'h44aaa591, 32'hc394ef9c, 32'hc38b5277},
  {32'hc4ad15ea, 32'hc353b974, 32'h43894edb},
  {32'h441287a0, 32'hc38ccf84, 32'h435f1e20},
  {32'hc344a810, 32'h42720286, 32'hc3ea2171},
  {32'h451f7b92, 32'h43962ea7, 32'h431ac2bc},
  {32'hc490b678, 32'hc2f5b642, 32'h43d577ac},
  {32'h4370e340, 32'hc2149e03, 32'hc31ebee4},
  {32'hc4d7f0de, 32'h43207dd9, 32'h42f6a979},
  {32'h44f6b0e0, 32'h43b35daf, 32'hc3debe38},
  {32'hc445cd9f, 32'hc3b2ef3d, 32'h43c7adf3},
  {32'h44fa1f71, 32'hc1dc0a71, 32'h4224b7a3},
  {32'hc4e9026a, 32'hc2e526a7, 32'hc291b70e},
  {32'h43b15ef0, 32'hc2b41b4e, 32'h431b65bc},
  {32'hc3ef8190, 32'h416a4041, 32'hc35ceb79},
  {32'h430c74e0, 32'h42aa9a16, 32'h437704ae},
  {32'hc4612da9, 32'hc2817a12, 32'h42a1a487},
  {32'h45239f69, 32'hc1a8c03f, 32'hc36d8a60},
  {32'hc4bb5764, 32'hc2d6fd2f, 32'hc350ae30},
  {32'h45136d99, 32'h432f27d8, 32'hc3626d44},
  {32'hc473657d, 32'hc282c15f, 32'h410eb44a},
  {32'h451070f3, 32'h416a484a, 32'h42b822b7},
  {32'hc4c23ff6, 32'h418092c6, 32'h43429023},
  {32'h44c003ae, 32'hc3830c54, 32'h42a68394},
  {32'hc4b110a5, 32'hc28fb16a, 32'hc3828d73},
  {32'h44c27303, 32'hc39652ed, 32'h41ee95c7},
  {32'hc47b6ed6, 32'hc32a3949, 32'h42503635},
  {32'h44047c9c, 32'h4306c9e0, 32'h42efdfee},
  {32'hc4d29e4e, 32'h431ae3ea, 32'h42d7739f},
  {32'h44e596d0, 32'h428133db, 32'hc14d7b00},
  {32'hc34e05f6, 32'hc3b805e7, 32'hc3834ae3},
  {32'h44e71274, 32'hc2e57e18, 32'h413d58ab},
  {32'hc491cb16, 32'h42a7e436, 32'hc2d9d051},
  {32'h450d3e72, 32'hc334923c, 32'h425179bc},
  {32'hc4c70fe3, 32'h42f922de, 32'hc2d8391a},
  {32'h444f4176, 32'hc2bad277, 32'hc3f06640},
  {32'hc525aec0, 32'h43b76a9e, 32'hc228ee3e},
  {32'h450533e8, 32'hc2ebf1f8, 32'h428d23f4},
  {32'hc4ee8cd0, 32'h426c6886, 32'hc34cb518},
  {32'h44cb6934, 32'h42d0bc4a, 32'h436c9246},
  {32'hc2a60b36, 32'h431f22b6, 32'h43718933},
  {32'h434d6fb8, 32'hc3999eac, 32'hc234da63},
  {32'hc471a154, 32'hc0501a28, 32'hc360f9ed},
  {32'h44bdecb6, 32'hc3582f08, 32'h4419a7db},
  {32'hc33065a0, 32'hc1e9a024, 32'hc0b19834},
  {32'h44bb77c9, 32'h4306c271, 32'hc305a65c},
  {32'hc5073471, 32'h425c14d2, 32'hc30b0b26},
  {32'h44550453, 32'hc324b36e, 32'hc2bacb1a},
  {32'hc47ff7ae, 32'hc3ca94fe, 32'h431bd25a},
  {32'h44f22d52, 32'h43516138, 32'h4218f235},
  {32'hc443d00c, 32'h4203ee2e, 32'hc3027adc},
  {32'h448073aa, 32'h42187e52, 32'hc35f1648},
  {32'hc48c1dbe, 32'hc389f2f0, 32'h426641e0},
  {32'h44dc7eca, 32'hc32caf17, 32'h42624fb6},
  {32'hc505bcb3, 32'h4209ccec, 32'h42805817},
  {32'h45055d13, 32'h4313025b, 32'h43c6e09e},
  {32'hc301b1eb, 32'h4312b81b, 32'h42d65c6a},
  {32'h438f5f68, 32'h42a8f36c, 32'h416b95ee},
  {32'hc407de89, 32'h4278a99e, 32'hc1adf047},
  {32'h449ff015, 32'hc2d90a49, 32'hc2f7da8e},
  {32'hc4451274, 32'h42a75dd4, 32'h44024dab},
  {32'h4480c1c6, 32'h425c2f8c, 32'h427dd273},
  {32'hc3befc6c, 32'h430373af, 32'h433cab2d},
  {32'h43719a6e, 32'h418de7ce, 32'hc3cb36f5},
  {32'hc2a8cad8, 32'hc35dfe72, 32'hc361dc95},
  {32'h43d6d500, 32'h4305b437, 32'hc4108dc1},
  {32'hc4db6043, 32'h41f1a031, 32'hc2fc78ba},
  {32'h45291840, 32'h438d0a22, 32'hc3ca5fd8},
  {32'hc4039156, 32'h43a393dc, 32'hc3b18a61},
  {32'h44422056, 32'h431fb04b, 32'hc014ba30},
  {32'hc43e03a2, 32'hc2b44e72, 32'hc200c9bb},
  {32'h44ae2806, 32'h4011f696, 32'hc2d54e9b},
  {32'hc4e17119, 32'h438741cb, 32'h4219eb8f},
  {32'h4508b016, 32'hc335362d, 32'h43ba33af},
  {32'hc4aa52b7, 32'hc1b1d559, 32'h42fdf938},
  {32'h44b5d302, 32'hc3104525, 32'hc3aa3197},
  {32'hc2cb3a98, 32'h424a6aa1, 32'hc3354a03},
  {32'h44c27a1a, 32'hc32c9320, 32'h435c9875},
  {32'hc4cfb20b, 32'h436bd02f, 32'h43f21bdc},
  {32'h44de07c2, 32'hc235a3fa, 32'hc2c0f2b6},
  {32'hc4f470b8, 32'h429fc9cb, 32'h433f2a7d},
  {32'h448eb826, 32'h41dd06e0, 32'h41a078cd},
  {32'hc464250a, 32'h42df4b0c, 32'hc273292c},
  {32'h44fdbed0, 32'hc33a5374, 32'hc343fef7},
  {32'hc4c0397e, 32'hc3b2b18c, 32'hc33213d5},
  {32'h446abdd2, 32'h424ece63, 32'hc33ef082},
  {32'hc40068c4, 32'hc3530de6, 32'h439b931b},
  {32'h451d65e3, 32'hc3055a4f, 32'h42195235},
  {32'hc4f1ba73, 32'h433bef91, 32'h42a97c30},
  {32'h43b4bafa, 32'h4341f345, 32'hc36e7647},
  {32'hc412ed3b, 32'hc2a81a3a, 32'h4357ad1c},
  {32'h44200527, 32'h4394f3e3, 32'hc2d825de},
  {32'hc4902348, 32'hc33a34b6, 32'hc2826740},
  {32'h44f28a1c, 32'hbf9a8338, 32'h4253fbe0},
  {32'hc4ee08f0, 32'h438d8f6c, 32'hc1d9bba0},
  {32'h42f31bcd, 32'h40e0d849, 32'h439224fc},
  {32'h44e835ba, 32'h43b86738, 32'hc3be0fae},
  {32'hc330e740, 32'h42ce2fa5, 32'hc2eab44e},
  {32'h4505094f, 32'h429f6c31, 32'h41b046b3},
  {32'hc4172e36, 32'h430ba814, 32'h434e8f75},
  {32'h43edb259, 32'h4305b1c4, 32'h4315d09c},
  {32'hc4ae3841, 32'h4384e98f, 32'h43905452},
  {32'h4443f62c, 32'h4315efb8, 32'h43ff548f},
  {32'hc3be11fc, 32'hc239d93e, 32'h420c66e3},
  {32'h449c2e66, 32'h42b4a472, 32'h42733689},
  {32'hc4b3667f, 32'h43baabc2, 32'hc1acfb16},
  {32'h4424ad40, 32'h43aa3baa, 32'h42e82983},
  {32'hc4e24215, 32'h42a52922, 32'hc273d0a2},
  {32'h44b36267, 32'hc293e403, 32'hc305b002},
  {32'hc5158d66, 32'hc312e239, 32'h42e8c8bc},
  {32'h44e95760, 32'h439ecf3f, 32'hc21b5cda},
  {32'hc31ae350, 32'hc33ae2e8, 32'h433d3b67},
  {32'h43901592, 32'h42d956ed, 32'hbf5d6e80},
  {32'hc378c74c, 32'hc3d776e7, 32'hc2e4219b},
  {32'h4459a380, 32'h439ca9de, 32'h42fa93f2},
  {32'hc29ebb60, 32'hc1a3d1b3, 32'h42421a69},
  {32'h452139b1, 32'h43d56899, 32'h43541a51},
  {32'hc4b614a4, 32'h420d9c3a, 32'h43318c89},
  {32'h44a5ccba, 32'h429f69c8, 32'hc3b1f8a3},
  {32'hc4ae895e, 32'h411c1314, 32'h42a9500b},
  {32'h44cab03d, 32'h4399920c, 32'hc3a9b01b},
  {32'hc3b38eb2, 32'h43970783, 32'h41c51ab4},
  {32'h44fe9aa3, 32'h434d8462, 32'h4297390b},
  {32'hc4103024, 32'h43384123, 32'hc38d7ed7},
  {32'h44b8fe94, 32'h434568ad, 32'hc37d8972},
  {32'hc4acf029, 32'h42032d00, 32'hc19a0fbf},
  {32'h44d9bcf1, 32'h4170ea28, 32'hc2cd3cd5},
  {32'hc498049e, 32'hc2883e5c, 32'hc2d25974},
  {32'h44ec4faf, 32'h4213ad7b, 32'hc2c0da2b},
  {32'hc3b8495c, 32'hc3e0bd59, 32'h42e68638},
  {32'h44e4550c, 32'hc30cc9cc, 32'hc31f6fbc},
  {32'hc4c237d8, 32'hc2d50c8b, 32'h43902cf6},
  {32'h44fc00f6, 32'h43046da1, 32'h429ed6ac},
  {32'hc3d588f8, 32'h443ba448, 32'h43bd43fd},
  {32'h4401d352, 32'hc25db3be, 32'hc2e1d986},
  {32'hc4a4b814, 32'h431de152, 32'hc3782374},
  {32'h44f92afc, 32'hc3907e99, 32'h3dc45780},
  {32'hc4ab23ad, 32'h43159d32, 32'hc2ad0c93},
  {32'h44b29ec1, 32'hc3200fd1, 32'h4394336a},
  {32'hc4c34a0b, 32'h436aa654, 32'h4239ea84},
  {32'h451580c2, 32'hc2e42fd8, 32'h4091372c},
  {32'hc4085610, 32'h43005502, 32'hc2bca11e},
  {32'h44565680, 32'h434b4fd0, 32'h43229e12},
  {32'hc500b07c, 32'h439414db, 32'h41895fdd},
  {32'h44f0b054, 32'h4311df4a, 32'hc3572ac6},
  {32'hc4fda2a0, 32'hc32a2f3a, 32'h42c6775e},
  {32'h44935073, 32'h41c98b51, 32'hc22f916c},
  {32'hc41c25f0, 32'hc32365fb, 32'hc3d597a0},
  {32'h450c2468, 32'h41ac692b, 32'h43c1f9e3},
  {32'hc5087097, 32'hc2d58738, 32'h42b69c2d},
  {32'h4487ebd0, 32'hc32cba69, 32'hc1f8cdb6},
  {32'hc3b63720, 32'h43ca22a1, 32'hc415d793},
  {32'h4499a50a, 32'h4003fe58, 32'hc3414b2b},
  {32'hc394e1c0, 32'hc37fb6d6, 32'hc316d7ba},
  {32'h43a6b802, 32'h433be829, 32'hc34cb3c6},
  {32'hc4200f42, 32'hc3c154a8, 32'hc326d968},
  {32'h43a9c015, 32'hc3db5e05, 32'hc4158187},
  {32'hc3b2ebf0, 32'h443354f0, 32'hc3ce90fb},
  {32'h40040700, 32'h413b4702, 32'hc27f1180},
  {32'hc4e7ecc8, 32'h438ed2f5, 32'h4289c8d0},
  {32'h450f9db5, 32'h413d363c, 32'h43bcadf8},
  {32'hc4bed431, 32'h4405f630, 32'hc44d9f98},
  {32'h440c53d8, 32'h43f9a2bc, 32'hc3bb16c9},
  {32'h42b964c4, 32'hc355ce5e, 32'hc2d2645b},
  {32'h44a6dcbc, 32'hc31915b0, 32'h429173fa},
  {32'hc50a7b46, 32'h431a0306, 32'hc28cd512},
  {32'h4493b65c, 32'hc316abc0, 32'h438b5449},
  {32'hc44e0d7e, 32'h42bf0c4e, 32'h42f967d4},
  {32'h44b5ebca, 32'hc4095766, 32'h431d304e},
  {32'hc4459613, 32'h4387ab76, 32'hc25bdbf9},
  {32'h44cfe0e7, 32'hc34f1851, 32'h43700ab6},
  {32'hc4780d14, 32'h4353006e, 32'hc374625d},
  {32'h451ec5bb, 32'h4230e95f, 32'hc2a716d3},
  {32'h4237d140, 32'h425d3f14, 32'hc3db785d},
  {32'h450a1193, 32'h42bbcfe0, 32'hc3973fba},
  {32'hc50b1508, 32'hc35faa91, 32'hc2ac7494},
  {32'h44fdfeb2, 32'hc3b4c97b, 32'h432b6545},
  {32'hc423154e, 32'h435f619d, 32'h43acd209},
  {32'h441bc740, 32'h43d9daff, 32'h43ae4e6d},
  {32'hc42f93e9, 32'h430660e3, 32'hc3820369},
  {32'h4234aac0, 32'h415f1a5a, 32'h423a831e},
  {32'hc480c054, 32'hc1fe67ce, 32'hc2eb29bd},
  {32'h4389aaee, 32'h43558d30, 32'h42dfba92},
  {32'hc4f1ccc1, 32'h436b96fc, 32'hc2528451},
  {32'h4495b300, 32'hc3e24b2a, 32'h44194bfb},
  {32'hc487eb1e, 32'hc3603d07, 32'h42bb975f},
  {32'h43f851da, 32'h43a69e5b, 32'hc296fee0},
  {32'hc48b1044, 32'h43caa9bc, 32'hc2ac5f99},
  {32'h44448ce0, 32'hc3b4427f, 32'h432de24d},
  {32'hc32a9c60, 32'h422b6236, 32'hc36f1fe8},
  {32'h431e9534, 32'h4381949e, 32'hc1a05bbd},
  {32'hc4ed2ba2, 32'hc39789bf, 32'h439803b3},
  {32'h4506ab68, 32'h420cdbe9, 32'hc3cedac3},
  {32'hc48c8251, 32'h43e53235, 32'h42d0b768},
  {32'h44bf4c86, 32'hc34afdc0, 32'hc36d9045},
  {32'hc500f9a1, 32'hc29a872f, 32'h43a21eda},
  {32'h45015f35, 32'h41e2a24e, 32'h435dfa2f},
  {32'hc4bd2e81, 32'hc345db31, 32'h4354d8bf},
  {32'h44e3b5c9, 32'hc1566db0, 32'h436fd885},
  {32'hc35c2de0, 32'h43076ad9, 32'h43b6387e},
  {32'h434bf188, 32'h437ca530, 32'h4397081b},
  {32'hc4a1bf66, 32'h43723731, 32'hc398c573},
  {32'h44994bb1, 32'hc2100d37, 32'hc288fef8},
  {32'hc4be815b, 32'hc3c7f110, 32'h42807876},
  {32'h45021498, 32'h431ca5ed, 32'hc35701e8},
  {32'hc3939b50, 32'h43cd414d, 32'h433aefe7},
  {32'h442d15e0, 32'hc38d783c, 32'hc3c5b6bc},
  {32'hc4e9c29b, 32'hc36830a5, 32'hc30f1c91},
  {32'h4423ac7c, 32'hc39d4823, 32'h4348abaf},
  {32'hc4a1fa34, 32'hc0784c3b, 32'h43a095a3},
  {32'h44681102, 32'h4320d449, 32'h432034de},
  {32'hc46ff27e, 32'h4265211c, 32'hc353b294},
  {32'h43c1be41, 32'h43078a66, 32'hc2d45141},
  {32'hc4fc8c30, 32'h43ad08bd, 32'hc26edef9},
  {32'h43ffd1f0, 32'h42a5e85c, 32'hc25b9e64},
  {32'hc4ee376f, 32'h43a60acb, 32'h413cc910},
  {32'h43c8b2af, 32'hc3d19b2a, 32'h43f24498},
  {32'hc4feeb34, 32'hc20903c5, 32'h4368bec4},
  {32'h439258a0, 32'hc2526e1b, 32'h42c44e9e},
  {32'hc4195976, 32'h4222ea16, 32'hc32acfc0},
  {32'h4429ff5d, 32'hc3085e6d, 32'h42196cec},
  {32'hc481041a, 32'h4383582f, 32'hc350501e},
  {32'h450dbc2d, 32'hc2375d6a, 32'h4387391a},
  {32'hc4beccf2, 32'h439f04b4, 32'h429e4e79},
  {32'h44f51b03, 32'hc301d188, 32'hc395a3e8},
  {32'hc4a895c3, 32'hc330fd94, 32'h43d10e83},
  {32'h43aeaa98, 32'hc1ba79c9, 32'h433cb531},
  {32'hc4775d53, 32'h422cf631, 32'h4270179a},
  {32'h4485dbc1, 32'h42bc2806, 32'h420efc75},
  {32'hc3df31da, 32'h4289dae9, 32'h431e61a9},
  {32'h43e5a560, 32'hc37a7382, 32'h436ed51c},
  {32'hc493dae4, 32'h421fd3af, 32'hc2a6f19c},
  {32'h446780a9, 32'h437f12fe, 32'h42cc3086},
  {32'hc515efc0, 32'hc0cf7658, 32'h43c83f32},
  {32'h43de5b1a, 32'hc3b64b88, 32'h432fe457},
  {32'hc4bf65fd, 32'h441259b9, 32'hc3124a8c},
  {32'h44aa62a4, 32'h42ea9e22, 32'h437b6913},
  {32'hc448f8c6, 32'hc2f475be, 32'hc19b149c},
  {32'h4484a805, 32'hc38d290c, 32'h40d59c4f},
  {32'hc4a23cb6, 32'h43fbc076, 32'h43146968},
  {32'h44b9488e, 32'hc3393460, 32'hc148feec},
  {32'hc3a5b910, 32'h42eee6b3, 32'hc2dfffe3},
  {32'h44de2f95, 32'h41d3011f, 32'hc3121974},
  {32'hc0f4eb12, 32'hc391b161, 32'hc3b47fd3},
  {32'h4465653a, 32'hc3a96fca, 32'hc2dcadbe},
  {32'hc3079370, 32'h4341a02d, 32'h434fbf7e},
  {32'h43d13378, 32'h4363608b, 32'h42b1cc36},
  {32'hc334ec18, 32'hc31afaab, 32'hc35f29d9},
  {32'h44fc598e, 32'h43f8b4e1, 32'h42d39479},
  {32'hc400828a, 32'h438d1502, 32'hc3cb23f2},
  {32'h4495e5dc, 32'h42adc4b3, 32'hc3552126},
  {32'hc51ce286, 32'h431a2954, 32'h4247c93a},
  {32'h443289b2, 32'hc3773652, 32'h43bb29e1},
  {32'h438470c8, 32'hc27b07e0, 32'h4208246d},
  {32'h451420ff, 32'h42a42365, 32'hc39d2bab},
  {32'hc2a53b60, 32'hc2cd2ada, 32'h4297c598},
  {32'h44fc0503, 32'h428c6e7d, 32'hc310bc5d},
  {32'hc3338ce0, 32'h42281ab4, 32'h42ca7cd0},
  {32'h440bb4ab, 32'hc2ffee01, 32'hc3371301},
  {32'hc4bdf7e4, 32'h4300f430, 32'hc2554774},
  {32'h441c0d14, 32'hc3ad1d80, 32'h411d992f},
  {32'hc42cb2f8, 32'hc3a4a4a8, 32'hc1e58e96},
  {32'h452232fd, 32'hc106526e, 32'h421a7e10},
  {32'hc4ccfb15, 32'h422b8e37, 32'hc1e0a13b},
  {32'h4486e5a1, 32'h42d70a84, 32'h42bd215c},
  {32'hc4e4a2e6, 32'h43a5cc4a, 32'hc27f33cf},
  {32'h43b05232, 32'hc1f1cba7, 32'h42ad7a3d},
  {32'h420f4120, 32'h435f9056, 32'hc09b6006},
  {32'h444385e8, 32'hc32d90ff, 32'hc2ec608a},
  {32'hc489cf3d, 32'h41f750b0, 32'h4399741e},
  {32'h44fa4e55, 32'h43d7b67b, 32'h430905e2},
  {32'hc43dd9b4, 32'hc3436ba1, 32'hc3404ed4},
  {32'h44758f4e, 32'h4280386b, 32'h4349e501},
  {32'hc4b1af9f, 32'h430deb4b, 32'hc2e0faff},
  {32'h445ce5b0, 32'hc109c1b0, 32'hc2fc2fb6},
  {32'hc5076722, 32'h431907d6, 32'hc3ef73b8},
  {32'h44872bf1, 32'hc3ac19a1, 32'h428ed3d9},
  {32'hc489c368, 32'h428114f2, 32'h436655f8},
  {32'h441b354e, 32'hc3ab2510, 32'hc2529d46},
  {32'hc4927587, 32'h439d6698, 32'hc2d0d5d8},
  {32'h43b6741c, 32'hc31569bf, 32'hc2fb26b0},
  {32'hc4c2de16, 32'hc2f6db42, 32'h4255a475},
  {32'h44b4df61, 32'hc2eb11de, 32'hc3434e36},
  {32'hc4b230be, 32'h43b3a147, 32'h42d27acb},
  {32'h44e64ff5, 32'hc301c91d, 32'hc3b3c6d6},
  {32'hc5077456, 32'hc379fe39, 32'hc2e16517},
  {32'h43a5cfb8, 32'h42c94f70, 32'h43851709},
  {32'hc5115250, 32'h4400e18f, 32'h437e99bd},
  {32'h450b12fd, 32'h436b0738, 32'hc2ce734e},
  {32'hc503e4aa, 32'hc226ca6d, 32'hc3fd4cb7},
  {32'h4480886e, 32'hc1522a6b, 32'h4083dc3e},
  {32'hc38e842e, 32'h410af72a, 32'h43ae5e89},
  {32'h45118df0, 32'h43809d96, 32'h430b4f74},
  {32'h437197e2, 32'h432ba57d, 32'h4220565a},
  {32'h440a8322, 32'hc3602b25, 32'hc22a9b10},
  {32'hc499ad33, 32'h42c706b7, 32'hc209d1fa},
  {32'h44d4d164, 32'h43b37d6d, 32'h4363d6e3},
  {32'hc412a96a, 32'hc3ed9f0c, 32'h427f126b},
  {32'h44b57a35, 32'h43516d11, 32'hc3c96a8b},
  {32'hc4abaaa4, 32'hc27aad3b, 32'h43233dbc},
  {32'h4516db29, 32'hc402386d, 32'h435dc548},
  {32'hc4d6ef66, 32'hc1928d21, 32'h4285d54d},
  {32'h44df7ac4, 32'h4386428e, 32'hc16caaab},
  {32'hc4e4dfe0, 32'hc3ac4fce, 32'hc35b8c78},
  {32'h44116d98, 32'hc2ad60d5, 32'h42c469cf},
  {32'hc36e0100, 32'h4322b8f7, 32'h43128242},
  {32'h4494dbb0, 32'hc16ddf18, 32'h42022bac},
  {32'hc482a2dc, 32'hc3192b0f, 32'h424930d3},
  {32'h4459f9d2, 32'h438d92f1, 32'hc3c452e6},
  {32'hc4ab80ae, 32'hc3301de1, 32'h442b96de},
  {32'h44a8a510, 32'h43814ac3, 32'h4379acb2},
  {32'hc43b0dd4, 32'h43872947, 32'h42ea1882},
  {32'h451923b2, 32'hc2bd319e, 32'hc33e25fc},
  {32'hc122c7c0, 32'h42675d63, 32'h42d098bb},
  {32'hc3965240, 32'hc2ef15d1, 32'h431eeca8},
  {32'hc41c8886, 32'h43969bbe, 32'hc2240777},
  {32'h44f7b746, 32'h4326f892, 32'h42e674fc},
  {32'hc4d39198, 32'h434a70dd, 32'hc345a1f0},
  {32'h44eed189, 32'hc30e7366, 32'hc334505d},
  {32'hc50dce0b, 32'hc34c392a, 32'hc3adc15c},
  {32'h44f41d8e, 32'h420c9216, 32'hc38c805d},
  {32'hc4816a93, 32'hc398140b, 32'hc3867479},
  {32'h44dc3614, 32'hc31013b6, 32'h42ec3168},
  {32'hc4b3680b, 32'hc3259474, 32'h42b351c7},
  {32'h44f483b4, 32'hc12a2a10, 32'hc37cbc30},
  {32'hc49ca10f, 32'hc2c6c7aa, 32'hc36de511},
  {32'h43069dd0, 32'h43a99118, 32'hc377af7a},
  {32'hc43e759c, 32'h4291fbe4, 32'hc34a107d},
  {32'h43c77bac, 32'hc38b54a1, 32'hc3db34ab},
  {32'hc431b2f5, 32'hc367174f, 32'hc28030b2},
  {32'h4490e0f4, 32'h430f96a1, 32'hc3985db8},
  {32'hc36f42d8, 32'h42baeef0, 32'hc264e690},
  {32'h44528198, 32'hc32cc5d4, 32'h428c2890},
  {32'hc4ca2954, 32'hc39b0510, 32'hc3993b15},
  {32'h44d70c6e, 32'h42f2b942, 32'h42fd06e9},
  {32'hc3eef108, 32'hc3953667, 32'h439428da},
  {32'h44edf85e, 32'hc200faae, 32'hc2bb8fd0},
  {32'hc46b8e17, 32'h42fef2cd, 32'hc177b366},
  {32'h44fb3567, 32'h422f8c44, 32'h41928f72},
  {32'hc4d38a93, 32'h4242861a, 32'h4292be45},
  {32'h4467bc78, 32'hbfbd3b76, 32'h432f7c34},
  {32'hc4d944a4, 32'hc390d306, 32'h43816284},
  {32'h4493bdae, 32'hc3a4b973, 32'h4309b922},
  {32'hc4c2096f, 32'h42d35a88, 32'hc2175f61},
  {32'h43b5826c, 32'hc31d7fca, 32'hc31fe632},
  {32'hc4029a78, 32'hc30a9728, 32'hc3b5490a},
  {32'h4401f768, 32'hc33a935a, 32'hc26e2805},
  {32'hc38bd190, 32'hc344438b, 32'h432a83f1},
  {32'h440bb02e, 32'hc2a3334f, 32'hc2e35840},
  {32'hc5024fd1, 32'h4300cdf4, 32'hc214055d},
  {32'h44cc1db3, 32'hc301f581, 32'h4387a9ee},
  {32'hc49c3dea, 32'h4309b504, 32'hc3f9fd1e},
  {32'h44f407d0, 32'hc30545ac, 32'hc2d23abf},
  {32'hc4b5d50b, 32'hc2b36a8b, 32'h43a0f13e},
  {32'h43f04168, 32'h43878d80, 32'h43926ca0},
  {32'hc3e6f290, 32'hc34792c6, 32'h4213c4c5},
  {32'h449f56d1, 32'h4342783e, 32'hc382e735},
  {32'hc3bba27a, 32'h4412d5d9, 32'hc1315e10},
  {32'h44a91e54, 32'hc2ebb6c5, 32'hc3f48a6b},
  {32'hc443e202, 32'hc3889717, 32'hc22ef5b6},
  {32'h44354608, 32'h440b20c5, 32'h43572697},
  {32'hc3e13334, 32'h43197602, 32'h43b8f09e},
  {32'h44803cf4, 32'h4378e5fc, 32'h4415c36e},
  {32'hc4e81f80, 32'h435932c9, 32'h42fbd098},
  {32'h45029c80, 32'h42a9f48f, 32'hc2abb965},
  {32'h42c0d320, 32'h424fe177, 32'hc3be3bd8},
  {32'h4514af7d, 32'h415cb317, 32'h4313c863},
  {32'hc4bb33ad, 32'hc2a3442a, 32'hc2b5f61c},
  {32'h4496b7ee, 32'hc3089f47, 32'hc2ea8f27},
  {32'hc51d8d00, 32'hc351f322, 32'h43832b33},
  {32'h44fd9b58, 32'hc0f4d9bf, 32'h424f9786},
  {32'hc508fe7a, 32'h4320af1a, 32'hc252ca80},
  {32'h44acb406, 32'hc3139c17, 32'hc343709d},
  {32'hc4eabe64, 32'hc33641d0, 32'h42812d92},
  {32'h44a1c5b3, 32'hc1fd9fdb, 32'hc34546f2},
  {32'hc4808f52, 32'h432f96c8, 32'h43a2a656},
  {32'h44f93443, 32'h42cacb25, 32'hc1ab9ea6},
  {32'hc45867a2, 32'hc2e89ba3, 32'h42ed7275},
  {32'h4508c097, 32'h4291ee28, 32'h42978b02},
  {32'hc4bb62ee, 32'h433849d9, 32'h42f2de14},
  {32'h44fb4ba2, 32'h43ba32f4, 32'hc1d5c695},
  {32'hc4685d8e, 32'hc2359941, 32'hc221449d},
  {32'h43fec158, 32'h42f23520, 32'h43b75080},
  {32'hc3aecfb2, 32'h430e676b, 32'hc31ce8b0},
  {32'h448c43ac, 32'hc3681fdd, 32'hc32d9be2},
  {32'hc464a054, 32'hc1b309ef, 32'hc3f77c42},
  {32'h44d82add, 32'hc2ba95ce, 32'h43a1252a},
  {32'hc4ad656f, 32'hc29e4a0d, 32'hc3b078b6},
  {32'h44388404, 32'hc38559b4, 32'hc281fe67},
  {32'hc4cfd928, 32'hc3983f58, 32'h42dff6e4},
  {32'h44803d70, 32'hc2866276, 32'hc35bd4a1},
  {32'hc1a6ea00, 32'h42c9f27a, 32'hc36ffcf6},
  {32'h452ada90, 32'hc2f44403, 32'hc2e32073},
  {32'hc4eb338c, 32'h43d4bac6, 32'hc30048bd},
  {32'h44588090, 32'hc2d7d2ef, 32'h43a57f8a},
  {32'hc4c8c4ca, 32'hc31e1ba4, 32'h43861961},
  {32'h45061eb2, 32'h442cb972, 32'hc3780cf6},
  {32'hc4efc3da, 32'h42147ce9, 32'h434d2585},
  {32'h44c04580, 32'h3c4f64c0, 32'h4327369a},
  {32'hc4ed3651, 32'h427c1cc0, 32'hc16acc23},
  {32'h44cfaf56, 32'hc10b960b, 32'hc3b4d68a},
  {32'hc506e394, 32'h436501a5, 32'h41bb298b},
  {32'h45262967, 32'h43a252af, 32'hc3fd1829},
  {32'hc4aba299, 32'h42e9d14d, 32'h42bcf693},
  {32'h44f995d3, 32'hc324834a, 32'h43949d37},
  {32'hc44b7e6e, 32'h43448d1f, 32'hc26198df},
  {32'h4452a927, 32'h42e701cf, 32'h4198bac1},
  {32'hc4d0f4ea, 32'hc1f08ddb, 32'hc3ad764c},
  {32'h4452105c, 32'h437a6ff4, 32'h43894f97},
  {32'hc4950dda, 32'hc39c5130, 32'h432b4a90},
  {32'h43bf89c2, 32'hc3304e50, 32'h3ffcdcb0},
  {32'hc46255b8, 32'h41f9e4d4, 32'hc332c6ab},
  {32'h4500e8aa, 32'h42119006, 32'h421d7e17},
  {32'hc4bc350a, 32'hc34d9b41, 32'h441f40cc},
  {32'h441674d8, 32'h4419c3f6, 32'hc3138e82},
  {32'hc455cf19, 32'hc053a91b, 32'hc3ac68aa},
  {32'h44a25f50, 32'hc04317a5, 32'h43a5e005},
  {32'hc4a5c037, 32'h414d39ad, 32'hc3b638e3},
  {32'h44aef73a, 32'h430f0e3e, 32'hc0ef3f38},
  {32'hc4733034, 32'h42571764, 32'h4284cad5},
  {32'h4491ab06, 32'h43a737de, 32'h43b7463c},
  {32'hc50286b9, 32'hc31d45a5, 32'h421714e3},
  {32'h42e9f338, 32'hc3aa8af1, 32'h43b84e29},
  {32'hc50d937f, 32'hc12ed1c9, 32'hc1f60850},
  {32'h44dd3d86, 32'hc21d42bc, 32'hc31cef70},
  {32'hc488f422, 32'hc269ce6e, 32'h438e66bd},
  {32'h44c0f718, 32'hc2372e18, 32'h434493b6},
  {32'hc32a2b67, 32'hc2b6237a, 32'h4343b17f},
  {32'h44e7f0b4, 32'h434af857, 32'hc3285f81},
  {32'hc432235a, 32'h43926d5b, 32'h421dca06},
  {32'h44bd7508, 32'hc389820d, 32'hc3135b1f},
  {32'hc4d39de5, 32'hc387b5b6, 32'hc35a6949},
  {32'h451295bb, 32'hc3f017ac, 32'hc341d214},
  {32'hc4d5ee81, 32'h437daac1, 32'hc39e31ba},
  {32'h450eff70, 32'h4095f6b4, 32'hc178dbd3},
  {32'hc4d04689, 32'hc40acae9, 32'h42ed5b10},
  {32'h44ed5f8a, 32'hc32c2ee7, 32'h433f76bc},
  {32'hc4c72284, 32'h430ed9ff, 32'hc3b29728},
  {32'h450594c7, 32'h4220d7ff, 32'hc3585ddd},
  {32'hc4cf9251, 32'hc28824c2, 32'hc4078b7a},
  {32'h44a1d592, 32'hc1de63e4, 32'hc385ffe6},
  {32'hc3775354, 32'h43804012, 32'hc3092a3d},
  {32'h44d472c8, 32'h427226d8, 32'hc1df4e34},
  {32'hc4c27bb2, 32'hc10c63f1, 32'h42c0b9d6},
  {32'h414b8780, 32'h42f404c5, 32'hc23e1f66},
  {32'hc43755e6, 32'hc26866ee, 32'h4255108e},
  {32'h44e510b1, 32'h42e6552c, 32'hc209cd9b},
  {32'hc362bbb0, 32'hc2df4945, 32'h426e21fb},
  {32'h446e9245, 32'hc2ddbcf9, 32'h4301cbf6},
  {32'hc4f25454, 32'hc39d8462, 32'hc3dec1b6},
  {32'h4349fc38, 32'h4312c2c4, 32'hc251fcbe},
  {32'hc3cae93c, 32'hc1d59438, 32'h4317ccbd},
  {32'h445aac18, 32'h43b5bd07, 32'h4151afe1},
  {32'hc492df99, 32'h436b49d7, 32'hc221c363},
  {32'h451c45d7, 32'hc1911798, 32'h4364b774},
  {32'hc49a7d80, 32'hc2866a0a, 32'h42ab3262},
  {32'h44f425ef, 32'hc225ff96, 32'hc329c7cc},
  {32'hc4f1f84c, 32'hc2ccb06c, 32'h43b0b8e5},
  {32'h44cec103, 32'hc34321f0, 32'hc2ba1f73},
  {32'hc4de028e, 32'h42da5f08, 32'h42b5abb6},
  {32'h4512cb22, 32'hc30d2057, 32'hc2b76da2},
  {32'hc424e4a0, 32'h439ebd68, 32'h42f14f59},
  {32'h4512d77d, 32'h4335aed3, 32'h4315124e},
  {32'hc4934bed, 32'hc335deb5, 32'h4394d94d},
  {32'h434787e0, 32'hc2a37514, 32'hc249aa32},
  {32'hc4dfd90e, 32'h43b32512, 32'hc3b5bcbb},
  {32'h45187fe8, 32'h43832b82, 32'hc34e013c},
  {32'hc4fc60a1, 32'hc32835c8, 32'hc31c652d},
  {32'h44b23d57, 32'hc2ca68da, 32'hc3870191},
  {32'hc2e30d20, 32'h4336fa5f, 32'hc34d40a8},
  {32'h451c5bfb, 32'hc394c58e, 32'hc2b8ac20},
  {32'hc480e917, 32'h41d1d60d, 32'hc2897c34},
  {32'h45070efc, 32'h41ce17a8, 32'hc3b1267a},
  {32'hc4174873, 32'hc30d5071, 32'h42d75d2e},
  {32'h445b2182, 32'h4315e93f, 32'h43c053a8},
  {32'hc5059d1b, 32'hc3798d9f, 32'hc09e0161},
  {32'h442123c8, 32'h43cff680, 32'hc1cfd757},
  {32'hc4d860cb, 32'hc1b0b7fd, 32'hc34ebf88},
  {32'h4497414d, 32'hc359a834, 32'h43c918fa},
  {32'hc32afe40, 32'h43ce1c82, 32'hc15f7304},
  {32'h43df435a, 32'h431979b1, 32'h42c94992},
  {32'hc4392372, 32'h42ded444, 32'h42859ed8},
  {32'h44b5b19b, 32'hc32080fd, 32'hc09544f9},
  {32'hc4bd2f78, 32'hc38234c4, 32'h43a304fb},
  {32'h44ca9df7, 32'h42f46578, 32'h43a2d02c},
  {32'hc3187150, 32'h440edf1e, 32'hc2ea6c42},
  {32'h44cf6cd8, 32'h4389c3d1, 32'h429b7f71},
  {32'hc40cfc92, 32'h43103c29, 32'hc35b71a7},
  {32'h44c27dc9, 32'h43854784, 32'hc3130fcc},
  {32'hc4e3da2c, 32'h432a36f7, 32'hc333bdba},
  {32'h44368d2c, 32'h43d2af37, 32'h43996862},
  {32'hc3842154, 32'h43a20147, 32'hc35e7f06},
  {32'h4425bb20, 32'hc3097fe8, 32'h439ffad8},
  {32'hc41de342, 32'h42b2c17f, 32'hbfa5a003},
  {32'h44fe695a, 32'h4317e1ef, 32'hc321626d},
  {32'hc3e03f35, 32'h43a058f8, 32'hc32faa8b},
  {32'h43b50dc6, 32'hc377c727, 32'h439ec263},
  {32'hc3f8bc10, 32'hc33bd992, 32'hc311bc45},
  {32'h4511fd93, 32'hc2c844fa, 32'h4399782f},
  {32'hc3bf55c0, 32'h4395e771, 32'h4286d713},
  {32'h44db71e5, 32'h432d9b24, 32'hc37cd471},
  {32'h42502d80, 32'h43cd7569, 32'hc27cdd2b},
  {32'h44645c84, 32'h431f700b, 32'h4344df2b},
  {32'hc4aa3eb1, 32'hc28b16b2, 32'hc393a7c6},
  {32'h44e34f5d, 32'h433b0a50, 32'h437920dc},
  {32'hc31611d0, 32'hc2f52f51, 32'hc3772013},
  {32'h449dfa50, 32'hc3995243, 32'h42326576},
  {32'hc464f924, 32'h42fe5c5e, 32'h4163c320},
  {32'h448293b3, 32'h437d41ad, 32'h431aa7d6},
  {32'hc39bcb30, 32'h4310329d, 32'hc379384f},
  {32'h4501b3ad, 32'h436f8d20, 32'h4346bd4e},
  {32'h42af6444, 32'h4304741c, 32'hc2f80b3f},
  {32'h44d64b90, 32'h40d6b060, 32'h436c5e1e},
  {32'hc4072a03, 32'h42243ca6, 32'h438c3985},
  {32'h450538fb, 32'h4035b0ba, 32'hc3c4ea75},
  {32'hc43aab2c, 32'h439ce0b0, 32'hc346c030},
  {32'hc2693868, 32'h429d5b57, 32'h435b2def},
  {32'hc5088faa, 32'h420c98c1, 32'h42cbe507},
  {32'h4392a868, 32'hc195d5be, 32'hc286f1ea},
  {32'hc4db5fbf, 32'hc3410070, 32'hc3a9d4fc},
  {32'h44400212, 32'h412004d8, 32'h43989668},
  {32'hc4851636, 32'h4224c948, 32'hc3d3a429},
  {32'h4452cc86, 32'hc38b9718, 32'h4330f313},
  {32'hc50b57ad, 32'h4337bef5, 32'hc195cb31},
  {32'h448100b5, 32'hc39a8d7e, 32'h43b45147},
  {32'hc52dd3d6, 32'h43a90aec, 32'h42b62463},
  {32'h44586ece, 32'hc25bc9e6, 32'h43d9926b},
  {32'hc4d0d124, 32'h42adbf66, 32'hc2ce6d29},
  {32'hc50e6e26, 32'hc31d1ff3, 32'hc2b1325e},
  {32'h4227d878, 32'h421ce86a, 32'h423437ae},
  {32'hc48063d4, 32'h41a45ef0, 32'hc3a56906},
  {32'h44d183a5, 32'hc2df0bae, 32'h41e92766},
  {32'hc46f9b28, 32'h429a079a, 32'hc3bd8cf2},
  {32'h42829610, 32'h44194994, 32'hc0821a27},
  {32'hc50232aa, 32'h4341e36e, 32'hc38a4ab5},
  {32'h44b15fd3, 32'h4293b60d, 32'hc36e2592},
  {32'hc3ada89c, 32'hc3bb975d, 32'hc0de20d0},
  {32'h449214dd, 32'hc1ffee4a, 32'hc29e6444},
  {32'hc4b2c3f9, 32'hc2ec2e90, 32'hc3aae3c0},
  {32'h44d1bfdd, 32'hc12e3f22, 32'h43180839},
  {32'hc45f7aa0, 32'h423960d6, 32'h4355f20e},
  {32'h44925939, 32'hc146964c, 32'h438488fd},
  {32'hc4042b51, 32'h42eac1a9, 32'h416be25b},
  {32'h44d244ff, 32'hc30231cd, 32'h40f22fae},
  {32'hc3f8d041, 32'h41ac24c1, 32'h4374a370},
  {32'h44ee0347, 32'h4385db7b, 32'hc314c8c9},
  {32'hc484fa4c, 32'hc37b5cca, 32'hc309cb1f},
  {32'h4525d2b5, 32'h4171992f, 32'h437c12d8},
  {32'hc4dc5d9a, 32'h40e1c3da, 32'hc2e0a084},
  {32'h44efbd8b, 32'h43ad1aef, 32'h4397eb9c},
  {32'hc404166e, 32'hc3305d66, 32'h43c1b146},
  {32'h45067bd2, 32'h42ff7e93, 32'hc2459d7a},
  {32'hc4b5c4b1, 32'hc3a95a97, 32'hc3a81197},
  {32'h44bfa4e1, 32'h43592c7e, 32'hc384fcd1},
  {32'hc47746bc, 32'hc360945f, 32'hc21513ed},
  {32'h449c5bfa, 32'hc417316c, 32'hc381660d},
  {32'hc45ba2c6, 32'h428cae9a, 32'hc4257199},
  {32'h442858b9, 32'h4325fe6f, 32'h41977760},
  {32'h41462100, 32'hc3135e3f, 32'hc36f7db4},
  {32'h4401a893, 32'hc3c72b4d, 32'hc3ba5a91},
  {32'hc470870d, 32'hc3f69f2f, 32'hc30ed917},
  {32'h445abecc, 32'hc3087762, 32'h40d7072d},
  {32'hc47fde33, 32'h43ffe343, 32'hc3843c7b},
  {32'h44c955b9, 32'h429a9571, 32'h438056f1},
  {32'hc5003e97, 32'h437e34d7, 32'h4318eb1a},
  {32'h450211c7, 32'hc35c0a02, 32'h43d13f14},
  {32'hc507151a, 32'h42bcef6c, 32'hc19afa6c},
  {32'h451446ea, 32'hc3e73066, 32'h43ac19ec},
  {32'hc418b30c, 32'h43796897, 32'h43530340},
  {32'h451127ba, 32'h426a33f4, 32'hc3a6e5ab},
  {32'hc44dca7a, 32'h43ab6929, 32'h41c153a9},
  {32'h42c1afd0, 32'h42c05740, 32'h44091038},
  {32'hc3b233c4, 32'h42aa4f5d, 32'hc114d437},
  {32'h4526112a, 32'hc272148a, 32'hc2c986bc},
  {32'hc4fed006, 32'h43db3efe, 32'hc393b636},
  {32'h4440a32e, 32'hc38a33c4, 32'h42dea4e9},
  {32'hc503bbe7, 32'hc24cc49f, 32'hc3af661e},
  {32'h450be57b, 32'h43c35634, 32'h43a6140e},
  {32'hc40aa670, 32'hc3b58832, 32'hc1add0a1},
  {32'h442679f8, 32'h43270414, 32'hc2ba8246},
  {32'hc495f401, 32'h431857b7, 32'hc3e6af81},
  {32'h44127aca, 32'h43bdfc42, 32'h426bfc3d},
  {32'hc49cea28, 32'hc3938908, 32'hc1fb1d55},
  {32'h4503bbb5, 32'h4384e970, 32'hc2467b7b},
  {32'hc4a7232b, 32'h4359049a, 32'h433676be},
  {32'h4412c689, 32'hc21442a7, 32'hc2e7a732},
  {32'hc3e24e70, 32'h42025096, 32'hc3916dbe},
  {32'h443b0e9c, 32'h43e111a2, 32'hc29d18ee},
  {32'hc36d3efe, 32'h439580d8, 32'h434699b6},
  {32'h44aac235, 32'hc13fb426, 32'h417bbcef},
  {32'hc41cb7e2, 32'hc3b6f78e, 32'hc25f8c16},
  {32'h42dd29df, 32'h42a250bb, 32'hc387702d},
  {32'hc4c69dec, 32'h41c6118a, 32'h42f0b6f8},
  {32'h439acc9c, 32'h42a179bd, 32'h43b8bd93},
  {32'hc4d8a42c, 32'hc38a1844, 32'hc2e06312},
  {32'h45234d38, 32'hc205b91a, 32'hc30480b6},
  {32'hc487f412, 32'hc3280eaa, 32'h4425e07c},
  {32'h443c514e, 32'hc301ba5e, 32'hc13a3b6d},
  {32'hc35609ee, 32'hc38f8865, 32'h42dd8836},
  {32'h44ac17ef, 32'hc387a0c6, 32'hc32b291c},
  {32'hc48b54e2, 32'h441fd663, 32'hc3cbc996},
  {32'h441ac68c, 32'hc3149ddf, 32'h413d2e90},
  {32'hc4a2148f, 32'h4316947e, 32'h43b42ce5},
  {32'h44d17e18, 32'h42eb8bd1, 32'h43d8fe10},
  {32'hc51f10d7, 32'h440c6285, 32'hc3bad9ab},
  {32'h43fee2f8, 32'h430c49d8, 32'h4219fa76},
  {32'hc4e520de, 32'hc247642d, 32'hc2b7c117},
  {32'h415f18b8, 32'h415e3e24, 32'h437be8f8},
  {32'hc4d224b8, 32'hc39708eb, 32'hc29b4c78},
  {32'h45009677, 32'h432ec1cf, 32'hc358625b},
  {32'hc507104f, 32'h41f436ce, 32'hc32d8421},
  {32'h44c3498f, 32'hc2a7b082, 32'hc412fcd3},
  {32'hc446f82e, 32'hc3f2dbe7, 32'h420f3338},
  {32'hc301f13d, 32'h425c5939, 32'h433a9d48},
  {32'hc4356ef7, 32'hc37c8823, 32'hc350dcc6},
  {32'h44b05d75, 32'hc295dfa5, 32'hc24ec142},
  {32'hc4fc5ffe, 32'h41893482, 32'hc08f7ff1},
  {32'h444e6fde, 32'hc2077a9d, 32'hc28cba36},
  {32'hc4b83841, 32'h43215bf8, 32'h430673df},
  {32'h4472d56e, 32'h42756c17, 32'hc33147e4},
  {32'hc41442c2, 32'hc1d46862, 32'h43c435a5},
  {32'h443db96a, 32'h4360618c, 32'h43c89bdd},
  {32'hc5138625, 32'hc39a5565, 32'hc37833dc},
  {32'h448f13c8, 32'h42d01045, 32'h43363c6f},
  {32'hc4f000ca, 32'hc3066673, 32'hc340017f},
  {32'h44418970, 32'hc3c2d8d9, 32'hc2a77172},
  {32'hc4d22195, 32'hc33aaf8e, 32'hc40ff748},
  {32'h4491e646, 32'hc3bdb35a, 32'h4391a497},
  {32'hc5072936, 32'h4330f6a0, 32'hc2bef45b},
  {32'h446b16ab, 32'hc3906ccc, 32'hc3a25e54},
  {32'hc413e23c, 32'hc2174763, 32'h42bffa4d},
  {32'h44de8796, 32'hc18e296f, 32'h43aec73f},
  {32'hc4483313, 32'h43622678, 32'hc336403f},
  {32'h4504840e, 32'hc29494a6, 32'h436cfc4d},
  {32'hc4b113ec, 32'h434d6bfb, 32'hc253b281},
  {32'h446503ef, 32'h3f381f50, 32'hc397917e},
  {32'hc4e1e022, 32'h430dce4f, 32'h4387448a},
  {32'h445b4f94, 32'h438cf23f, 32'hc3030461},
  {32'hc4ecbdc8, 32'hc24366b0, 32'h433b8770},
  {32'h43ac0c98, 32'h432cb98a, 32'h43936fbb},
  {32'hc51dee63, 32'hc2dd23be, 32'h42947d49},
  {32'h44ffbe76, 32'h43638b69, 32'h43074cae},
  {32'hc502dbba, 32'h4210bf7a, 32'h4297f13e},
  {32'h44c1e75d, 32'hc27034fc, 32'hc364f5db},
  {32'hc4aa0426, 32'hc403684d, 32'h431d9e78},
  {32'h4519a2df, 32'h4335495f, 32'h436284ff},
  {32'hc4d3ee3a, 32'h42430377, 32'hc289a2a3},
  {32'h43a91bbe, 32'hc2878f52, 32'h439300e6},
  {32'h42bbcdc0, 32'hc355412d, 32'h434ffeee},
  {32'h4505b558, 32'h41eb3c2c, 32'hc3ada866},
  {32'hc4f39200, 32'h428d46b0, 32'hc2ce8dbe},
  {32'h444b2b6e, 32'h42f38f70, 32'hc2abd7e8},
  {32'h42e83ae0, 32'h43815422, 32'hc2936ba1},
  {32'h44a2f450, 32'h43943f91, 32'hc2802164},
  {32'hc40f04b8, 32'hc314c6ba, 32'hc363945d},
  {32'h44c2cccc, 32'h42e961f4, 32'hc28a5cd2},
  {32'hc4b8465e, 32'h4272af14, 32'h434a4829},
  {32'h4455f4b0, 32'hc005fb18, 32'hc1b29edc},
  {32'hc4eb3ac0, 32'h425d1515, 32'hc39398d0},
  {32'h44ce56d9, 32'hc28a4759, 32'h432042a2},
  {32'hc5016f1d, 32'h439f5562, 32'h43811278},
  {32'h445ac543, 32'h42b2bc6d, 32'hc2be1d74},
  {32'hc518d39f, 32'h431a28a8, 32'hc317909e},
  {32'h43813720, 32'hc35bbef7, 32'hc3af9d55},
  {32'hc48385a4, 32'hc33ddc77, 32'h43369a30},
  {32'h44f52a61, 32'hc3a5db52, 32'hc1b428d5},
  {32'hc4277282, 32'h4370b63a, 32'hc2a95f6e},
  {32'h449ba6ca, 32'hc31b3d2c, 32'h432ba7b8},
  {32'hc465b688, 32'h432b4e2e, 32'h4329b38a},
  {32'h449483b0, 32'hc128c0d2, 32'hc23a7d1e},
  {32'hc505f23c, 32'h42f65ad5, 32'h41885cea},
  {32'h4222d722, 32'hc3b41a25, 32'hc17a21ef},
  {32'hc437c278, 32'h42a00c38, 32'hc2ba4a02},
  {32'h450ad6ab, 32'h42091777, 32'h43109597},
  {32'hc4103b5a, 32'h42a23a0b, 32'h4229cd22},
  {32'h44e69bb0, 32'h42a30762, 32'h43b3f91a},
  {32'h433ba124, 32'h43f1ce86, 32'h4371a0de},
  {32'h44bb1d6a, 32'h4332e7e3, 32'hc37c09ef},
  {32'hc4367f34, 32'hc39485f3, 32'h42b1c1ce},
  {32'h43d9df46, 32'hc33a19ab, 32'hc3c24b41},
  {32'hc4184734, 32'hc27f420e, 32'hc296a6b0},
  {32'h42ca69d0, 32'h3f9dd813, 32'h42a01652},
  {32'hc379b014, 32'h43241914, 32'h43340fc9},
  {32'h439fd50c, 32'h42530e90, 32'h4309b368},
  {32'hc4745bd8, 32'hc39b3f4b, 32'hc2f7278a},
  {32'h446266b4, 32'h422fca83, 32'h42f2aacf},
  {32'hc48b56bf, 32'hc23459a8, 32'h4337f6ed},
  {32'h44e423f8, 32'h42eb353e, 32'hc3da8024},
  {32'hc4f05555, 32'hc308d016, 32'hc33a2994},
  {32'h4500a760, 32'hc3809163, 32'h42bcea00},
  {32'hc5073946, 32'h42e36424, 32'hc3810cbc},
  {32'h44fb803a, 32'h42bfd87f, 32'hc3162e43},
  {32'hc4a10caf, 32'hc36c188d, 32'hc2dc842f},
  {32'h4320ca48, 32'h42244d92, 32'h42942d7d},
  {32'hc4325ffc, 32'h43ecbf62, 32'h4286e299},
  {32'h448cf6b4, 32'h433ae204, 32'h42973d7c},
  {32'hc3638dbc, 32'hc215a4ee, 32'h43809120},
  {32'h44edfa8c, 32'hc22e0c0d, 32'h43033aa5},
  {32'hc49ac4b8, 32'hc1a6f877, 32'hc2ca2d4b},
  {32'h4503fbbb, 32'hc315b793, 32'hc3c47e03},
  {32'hc333d2ae, 32'h433df2a0, 32'h429f378d},
  {32'h439c4050, 32'h441855fb, 32'hc2f3fffb},
  {32'hc4061691, 32'h4399f1c4, 32'h42c66dee},
  {32'h4508ed6e, 32'hc3cb849a, 32'h433483ed},
  {32'hc5024053, 32'hc2dbff10, 32'hc4174648},
  {32'h440f68c4, 32'hc2a3b975, 32'hc1d0d5ad},
  {32'hc4e2791b, 32'hc36f3aac, 32'h43385ac0},
  {32'h44df3dca, 32'hc30890e3, 32'hc3a4a34a},
  {32'hc5067e75, 32'h42f4b035, 32'h416c0302},
  {32'h447c27e3, 32'hc3392afa, 32'hc3b4d39d},
  {32'hc50ae784, 32'hc427def2, 32'h434d8055},
  {32'h4500baf4, 32'h435dbef1, 32'hbfb07620},
  {32'hc4aeccaf, 32'hc413b072, 32'hc29c4116},
  {32'h45039663, 32'h43198a7e, 32'hc30260bd},
  {32'hc4c5819c, 32'h42a71032, 32'h43ffca6e},
  {32'h44c3362f, 32'hc2bfdd00, 32'h439399cf},
  {32'hc46483e3, 32'hc306c953, 32'hc23ef00b},
  {32'h44b6d400, 32'h42c82383, 32'hc311893b},
  {32'hc4b188a8, 32'hc39a3e1a, 32'h42eecaf3},
  {32'h4525db56, 32'h42a78276, 32'hc2a46303},
  {32'hc4af15e5, 32'h43145f34, 32'hc37e4877},
  {32'h449720dd, 32'hc39f7dd5, 32'h42bd17ac},
  {32'h4373dd31, 32'hc33a83c3, 32'h421cb579},
  {32'h450144f4, 32'h43237ab2, 32'h4225834c},
  {32'hc4f9e963, 32'h424e7e8e, 32'hc31a48d2},
  {32'h44f0183a, 32'h42d47228, 32'hc2bb5ad6},
  {32'hc4977bd1, 32'h4319933e, 32'hc3430d4f},
  {32'h44aeb97d, 32'hc355f2a9, 32'hc2c3ad7a},
  {32'hc4bdf960, 32'hc117a6fe, 32'hc31202c0},
  {32'h43f234bc, 32'hc2e8551c, 32'hc22e3e9c},
  {32'hc4acdb7c, 32'h43c5d4c3, 32'hc356ed7e},
  {32'h44ff0414, 32'h43428edb, 32'h437075a1},
  {32'hc34e54e0, 32'hc3acfee2, 32'hc1eafe9d},
  {32'h44fc5ecf, 32'hc30f9f2d, 32'hc3219d0b},
  {32'hc4e5f259, 32'h427bc6ab, 32'h432fae66},
  {32'h4500ff2e, 32'h43966f2f, 32'h439e6212},
  {32'hc4da6cc5, 32'hc355b9d7, 32'h4304e961},
  {32'h43e8116c, 32'h432f30b6, 32'h4349c2bf},
  {32'hc478b756, 32'h439f306c, 32'h4387b43c},
  {32'h44c81f73, 32'hc3e289f6, 32'hc424e09c},
  {32'hc4e6f191, 32'hc3810844, 32'hc20f6088},
  {32'h449665e2, 32'hc3ca4d09, 32'h42f94313},
  {32'hc4850bc0, 32'h438eddfb, 32'h43a5067b},
  {32'h44de062d, 32'h41449dfb, 32'h42a631fc},
  {32'hc444c456, 32'hc301a2e9, 32'hc39545f0},
  {32'h4402b1c5, 32'hc34fe488, 32'hc38d93d3},
  {32'hc44d722f, 32'hc3509dc8, 32'hc1c5ba07},
  {32'h451ae469, 32'hc24a4a03, 32'hc3993513},
  {32'hc46b8532, 32'hc25223a4, 32'h43a91839},
  {32'hc2485165, 32'h438fc44c, 32'h43845b3c},
  {32'hc4ba7ae6, 32'h42c28693, 32'hc387f43b},
  {32'h446f9578, 32'h42acf88f, 32'hc380f8bc},
  {32'hc48dae97, 32'hc1aaf803, 32'hc28320c4},
  {32'h444b145a, 32'h431cc971, 32'h430af873},
  {32'hc45a80f3, 32'h44390c6c, 32'h4387ccec},
  {32'h45232937, 32'h4059d268, 32'h423765ac},
  {32'hc488b544, 32'h428d13fb, 32'h43cb3ed2},
  {32'h44183617, 32'h414c676c, 32'hc2d3430c},
  {32'hc4eb2e59, 32'hc358085d, 32'hc2a05de1},
  {32'h44aaaac0, 32'h43abfe10, 32'hc3910647},
  {32'hc4c610d8, 32'hc2aec997, 32'h423ad4ba},
  {32'h4488b246, 32'hc39c0f19, 32'h43a26e0e},
  {32'hc415227c, 32'h4133e6f2, 32'hc320409e},
  {32'h44ce3e5a, 32'h42c135e9, 32'hc377afd3},
  {32'hc508560a, 32'h42da4c8e, 32'h43ac1363},
  {32'h44716cd1, 32'h42f513ed, 32'hc34e37e6},
  {32'hc30ccccc, 32'hc1b58c07, 32'hc3de7b73},
  {32'h44e6a1ee, 32'hc304e99a, 32'h432f58ab},
  {32'hc4a1dc04, 32'hc3e50f57, 32'hc23485fa},
  {32'h44e27d8a, 32'hbe75c6ef, 32'hc3526405},
  {32'hc4ded888, 32'h43271c60, 32'hc2d516b1},
  {32'h451f3168, 32'hc369dc0f, 32'hc31b89c1},
  {32'hc4ab334b, 32'hc149eec1, 32'hc2a1c151},
  {32'h4441054a, 32'hc234dc0e, 32'h4347b102},
  {32'hc4617229, 32'h440f2b4d, 32'hc34103a6},
  {32'h44f4677e, 32'hc2579b4c, 32'h425d6e6b},
  {32'hc4c017e2, 32'hc27b36da, 32'hc3af7010},
  {32'h434a635a, 32'hc41115c3, 32'hc3168def},
  {32'hc4f38804, 32'h4313fe78, 32'hc3160653},
  {32'h434729ad, 32'hc1b54c3d, 32'h438265ea},
  {32'hc50ef22e, 32'hc29fc174, 32'hc25a7b00},
  {32'h449bb0f8, 32'h42faa6ff, 32'h41a8372f},
  {32'hc514e887, 32'hc14a4347, 32'h43f06f5f},
  {32'h4500fc0b, 32'hc3317ed7, 32'h42b76c35},
  {32'hc4440834, 32'hc3239f04, 32'hc3bbfda8},
  {32'h44040d78, 32'hc2f4aeaf, 32'h4187cab3},
  {32'hc4af25b3, 32'h42cb0cf4, 32'h429327ef},
  {32'h44e639be, 32'h430eb527, 32'h432f917e},
  {32'hc449a470, 32'h4132f4ff, 32'h42815bce},
  {32'h44e076a8, 32'h4239f638, 32'h42803280},
  {32'hc50757b8, 32'h43ecb973, 32'h429c9fa9},
  {32'h4509d85c, 32'h4310ffec, 32'h43faf55a},
  {32'hc4af2a7c, 32'hc359bba2, 32'h4356199a},
  {32'h43678f28, 32'h40b18757, 32'h42203008},
  {32'hc4bfdaf8, 32'h41bdee47, 32'hc314ad3d},
  {32'h4505ec02, 32'h43d9ea87, 32'hc33a3fc9},
  {32'hc4f44528, 32'h43cf151b, 32'hc3a3162f},
  {32'h430b6330, 32'h43a6a4c0, 32'hc2165f14},
  {32'hc3e53d51, 32'hc38110e2, 32'hc18022ef},
  {32'h44f6cfd2, 32'h42ac691a, 32'hc34a1d91},
  {32'hc4ce64f4, 32'hc2997778, 32'hc29006dc},
  {32'h450013ae, 32'hc14f1c09, 32'hc21e0ca6},
  {32'hc4159502, 32'hc2f2edb7, 32'h4398dd52},
  {32'h44af9721, 32'hc20338a6, 32'hc3800b17},
  {32'hc506d0c8, 32'hc3b8665f, 32'h429bfc3c},
  {32'h44be6d6e, 32'h4332632f, 32'hc246a605},
  {32'hc4cb5d86, 32'h432fc00d, 32'hc316265d},
  {32'h4461847c, 32'hc30fbad7, 32'hbfc78ea5},
  {32'hc4428cec, 32'hc28a0000, 32'hc31efb49},
  {32'h441a3874, 32'hc36470f3, 32'h432f79cb},
  {32'hc48d5cc9, 32'h4328d38b, 32'h4388eb28},
  {32'h44805b10, 32'hc355361b, 32'h43973338},
  {32'h4231f962, 32'h42998b6f, 32'hc307ed72},
  {32'h4490e6b9, 32'hc347cef9, 32'h43ebf0e2},
  {32'hc4d5e65f, 32'h42149227, 32'h43df20ca},
  {32'h441ed738, 32'hc37544ac, 32'hc2b9fda0},
  {32'hc4f1ab57, 32'h4390654d, 32'h43912284},
  {32'h43eb9244, 32'h4396d04a, 32'hc322db47},
  {32'hc301f500, 32'hc3992842, 32'hc21defc5},
  {32'h449cb1f0, 32'hc206578b, 32'hc3144b9d},
  {32'hc456271c, 32'h430b9d82, 32'h44235720},
  {32'h43d3977a, 32'hc34fb9eb, 32'hc40e00dc},
  {32'hc4993a90, 32'h41f766fd, 32'h4114b5c8},
  {32'h4444e380, 32'hc38b6a10, 32'hc30d8ae0},
  {32'hc4d1ba63, 32'hc2b42083, 32'hc2ce3739},
  {32'h448ed838, 32'hc37b93df, 32'h41e580d6},
  {32'hc3ccd750, 32'hc3d80548, 32'hc33bbc42},
  {32'h448a4f92, 32'h4137f55c, 32'h42a7e042},
  {32'hc49413dc, 32'h4345d398, 32'h417f4d5d},
  {32'h44433218, 32'h42df9da4, 32'hc31c3d93},
  {32'hc4b84090, 32'h42e53c7a, 32'hc383b565},
  {32'h44452609, 32'hc3a9e21d, 32'hc3da7072},
  {32'hc426608c, 32'h43399a7d, 32'hc1b0b534},
  {32'h44f13d97, 32'hc3afda62, 32'hc3985a15},
  {32'hc42c4998, 32'h4211d095, 32'h4225f02d},
  {32'h447bd9cc, 32'h41f8c32b, 32'hc317e4ca},
  {32'hc48555fa, 32'h428be4f8, 32'h43a117e3},
  {32'h441a36a3, 32'hc2f344a9, 32'h438d6442},
  {32'hc4ab4b5a, 32'hc0112c88, 32'h41e08564},
  {32'h44400e9c, 32'h4331dff1, 32'hc1ad8119},
  {32'hc4089a44, 32'h419e238f, 32'hc314dcfb},
  {32'h4484f8f7, 32'hc2d69fee, 32'hc21d4953},
  {32'hc4b0e0e5, 32'h41f563fb, 32'h41be20a6},
  {32'h45111bdb, 32'hc3510867, 32'h4363ba84},
  {32'hc3ec1fd0, 32'h438f8ce1, 32'hc40126a9},
  {32'hc26f58a0, 32'h42340a2e, 32'h4341a062},
  {32'hc4d5193c, 32'hc3242b3e, 32'hc30a96ec},
  {32'h415ad600, 32'h42c3b0ff, 32'hc280eda4},
  {32'hc386eb58, 32'h43383ece, 32'hc424cd9a},
  {32'h4433be83, 32'hc3d368c5, 32'h43083274},
  {32'h436b6d00, 32'hc3b32aa6, 32'hc305ea66},
  {32'h441a6c98, 32'hc3cff074, 32'h43d96b70},
  {32'hc4713f9d, 32'hc2ad2a7f, 32'h42faa1f6},
  {32'h43ee56ca, 32'h42ef751e, 32'h41cbdaca},
  {32'hc5149986, 32'hc212a019, 32'hc38ff061},
  {32'h43d3a02c, 32'h43b7b79d, 32'hc293221a},
  {32'hc409a3ab, 32'h42ff501e, 32'hc39ec241},
  {32'h44ca4241, 32'hc2cd9240, 32'hc355895b},
  {32'hc4b3932c, 32'h4432d459, 32'h434fff87},
  {32'h43a2e850, 32'hc37881cb, 32'hc3166e2e},
  {32'hc4d01c81, 32'h42e7c058, 32'hc318a0b1},
  {32'h451d462b, 32'hc3e32cbf, 32'h41b36e8d},
  {32'hc39f0533, 32'h434f4663, 32'hc4089746},
  {32'h451af9b9, 32'hc33b135f, 32'hc331c1de},
  {32'hc4cf4397, 32'hc2461176, 32'hc452ae02},
  {32'h450807ab, 32'hc27a807d, 32'hc342647a},
  {32'hc484397c, 32'hbf9301f0, 32'h42ebddda},
  {32'h446fb1d4, 32'hc3436bc7, 32'h42a7e9d9},
  {32'hc4ed7c29, 32'h43603830, 32'h43c6b908},
  {32'h44a1b672, 32'h43080b12, 32'hc3731df1},
  {32'hc3027b28, 32'hc2a7a74f, 32'h431dd6ca},
  {32'h44c433d7, 32'h437b776e, 32'hc3bb55bc},
  {32'hc5019950, 32'hc366167c, 32'hc2c357da},
  {32'h448c0454, 32'h4327e502, 32'hc39df4ef},
  {32'hc50f82a3, 32'h43200d67, 32'h42a4e127},
  {32'h440cc1a7, 32'h414ffed8, 32'h4380478b},
  {32'hc5191213, 32'hc2abcea1, 32'hc2d4f060},
  {32'h44fae7f8, 32'h427e3bc0, 32'hc378c4fe},
  {32'hc4ab0e78, 32'hc391db4d, 32'h42098efb},
  {32'h446729c0, 32'hc3c59466, 32'h4162370a},
  {32'hc41a4040, 32'h4424e0f7, 32'h430ace24},
  {32'h44fb2468, 32'hc3748403, 32'hc2302334},
  {32'hc3718850, 32'h434537e3, 32'hc3775b25},
  {32'h44dc1399, 32'h43124229, 32'h43223da1},
  {32'hc4070347, 32'hc0070ba4, 32'h4322cd01},
  {32'h4400c698, 32'hc3b2c92e, 32'h434f84a6},
  {32'hc4a6e14c, 32'h429b8c91, 32'h41d659af},
  {32'h443ffda6, 32'hc3a8359c, 32'h430b9d55},
  {32'hc4730cf6, 32'hc36dff8c, 32'hc3b46d32},
  {32'h44fd92a0, 32'h4341f780, 32'h42d5e2ba},
  {32'hc2f29aa0, 32'hc33dcd67, 32'h433b76fc},
  {32'h43e2f928, 32'hc2b3dadd, 32'h430cf05c},
  {32'hc515c57e, 32'hc3417832, 32'h4385cb70},
  {32'h4409c63c, 32'h433162dc, 32'hc25e9b74},
  {32'h40387a00, 32'h42b3da03, 32'hc3ca9e95},
  {32'h44bdbe8e, 32'hc31c9de3, 32'hc34e5e66},
  {32'hc49190fd, 32'h43240b26, 32'hc36b8cda},
  {32'h4500ce90, 32'h423a96ee, 32'hc3099fa6},
  {32'hc4ad137d, 32'hc3842284, 32'h4305a83d},
  {32'h452560d6, 32'h42d3f14d, 32'hc30eed51},
  {32'hc436b8c8, 32'h3f88071b, 32'hc292bf29},
  {32'h43e05bff, 32'hc39273f2, 32'hc2e905b4},
  {32'hc4fe6e7a, 32'h421ef42b, 32'hc2bfcc15},
  {32'h4516f97c, 32'hc3f4cc32, 32'h43507521},
  {32'hc4050c84, 32'h439f674b, 32'hc2c336e2},
  {32'h44e5a11b, 32'h3f901605, 32'h438930d0},
  {32'h4200eec0, 32'h421f6270, 32'h4289dec6},
  {32'h44eb428f, 32'hc1eb6785, 32'hc08d8eda},
  {32'hc350ecc2, 32'hc3538a93, 32'hc1547dd9},
  {32'h44f10867, 32'h437b450f, 32'h43ec0846},
  {32'hc4d5c2c5, 32'hc36862d5, 32'h43b127d7},
  {32'h45107938, 32'hc37a19fd, 32'h42060f52},
  {32'hc51277e3, 32'h429966de, 32'hc326d783},
  {32'h448dbfc5, 32'hc07afab5, 32'hc393a283},
  {32'hc21c32b0, 32'hc34f06ce, 32'h4315dd73},
  {32'h437b28f0, 32'hc2a04d58, 32'h42d3215c},
  {32'h4343bda8, 32'h410c80c6, 32'h438049be},
  {32'h4509a31d, 32'h427f28fb, 32'h41e08769},
  {32'hc4f4f3b2, 32'h41444935, 32'h43997160},
  {32'h44ea7ec8, 32'hc3002e14, 32'h43549d8b},
  {32'hc3f4f8b8, 32'hc3eef518, 32'h435ebca1},
  {32'h44907519, 32'hc3a459b1, 32'h41f7f24a},
  {32'hc517675b, 32'h43ad58ed, 32'hc32962bc},
  {32'h44a58322, 32'h435cae29, 32'hc31577b8},
  {32'hc4956c8c, 32'hc2933bf8, 32'h424cf232},
  {32'h4509c4f2, 32'hc2cd4fde, 32'hc358bbd7},
  {32'hc498277e, 32'hc3354c06, 32'h4337777c},
  {32'h4429ae18, 32'h4290dc58, 32'hc44b5f55},
  {32'hc4c1db91, 32'hc1c637e8, 32'hc2d21386},
  {32'h44466650, 32'h42a6ebd2, 32'hc34837a9},
  {32'hc4b432d2, 32'hc3f92031, 32'h439a38a4},
  {32'h434a554e, 32'hc3d67ddd, 32'h43c4a3ef},
  {32'hc5031809, 32'hc3c0ef86, 32'h433efa1b},
  {32'h446092d2, 32'h42e62f42, 32'h42b3af1b},
  {32'hc4063668, 32'hc2999a6a, 32'hc0b282e4},
  {32'h44ee88d4, 32'hc329b016, 32'hc3c82298},
  {32'hc3d66b14, 32'h4387276a, 32'h41fefc1a},
  {32'h444a9747, 32'h440e3869, 32'h430a4399},
  {32'hc4879108, 32'h4333ad2e, 32'h42f5c8e1},
  {32'h4498faad, 32'h42e27229, 32'h437d5abd},
  {32'hc5122074, 32'h437e97b3, 32'h43246867},
  {32'h440e1124, 32'hc33c53b2, 32'hc23ab5c6},
  {32'hc47784a1, 32'h42c359a0, 32'h434abcca},
  {32'h44323821, 32'hc31c2d91, 32'h4258c0a4},
  {32'hc51ef205, 32'h4348f53f, 32'h430c8140},
  {32'h444df2b6, 32'h424c58ac, 32'hc31d8b01},
  {32'hc4885a37, 32'hc34c219a, 32'h43d41d22},
  {32'h44f7c577, 32'h435fe7ad, 32'hc33f579a},
  {32'hc4857dd7, 32'h43bb6ea9, 32'hc3da801a},
  {32'h43b0e130, 32'h42e3d83a, 32'hc32e2580},
  {32'hc34334f0, 32'h43903cca, 32'h43836bf4},
  {32'hc23b8b6e, 32'h43ad57d4, 32'hc4310269},
  {32'hc45c3387, 32'hc28c5651, 32'h439d01ad},
  {32'h4514fc99, 32'hc3053f62, 32'h42ee1254},
  {32'hc444b195, 32'h43097109, 32'h43375047},
  {32'hc20efe68, 32'hc266f03d, 32'h4391b57b},
  {32'hc4de81d0, 32'h41fb0042, 32'h41784ca6},
  {32'h438590ec, 32'hc3c003f5, 32'hc33f1342},
  {32'hc4c0f934, 32'hc1725f88, 32'hc22ca70a},
  {32'h443ae242, 32'hc369ba60, 32'h43b3aed0},
  {32'h433c8f08, 32'hc39af969, 32'h436ef0d8},
  {32'hc411b030, 32'h42d4def8, 32'h43382c7c},
  {32'h4260cca0, 32'hc2ea67c0, 32'h440ac032},
  {32'hc5021da0, 32'h42fd9f44, 32'hc1e24cfa},
  {32'h44e58f01, 32'hc37d794a, 32'h43363a80},
  {32'hc4c84ae2, 32'h41ef2d28, 32'h43b1aaff},
  {32'h451e4e69, 32'hc3fbb21b, 32'hc362bff3},
  {32'hc4f06d0d, 32'hc2de6bbf, 32'hc336a014},
  {32'h44da1754, 32'hc337e867, 32'hc36c742e},
  {32'hc4c229cb, 32'h42fad97f, 32'hc37e3c4f},
  {32'h446836ec, 32'hc3456bf3, 32'hc30b88bf},
  {32'hc496d093, 32'hc2f62557, 32'h4313f728},
  {32'h447a94dc, 32'h4379b830, 32'h412adb5b},
  {32'hc49d88e8, 32'h434f37e0, 32'hc37a2b1f},
  {32'h44a4f081, 32'hc3633b44, 32'hc3574f85},
  {32'hc3a86f40, 32'h4100e2e8, 32'h438b15ea},
  {32'h45050244, 32'hc3ad58ad, 32'h4308c9a8},
  {32'hc50b737b, 32'h423277ec, 32'h4303f136},
  {32'h44d10f4e, 32'hc317a7f6, 32'h432b7197},
  {32'hc4abd291, 32'h43f494e3, 32'h43ab67a5},
  {32'h443b2886, 32'hc2e5de37, 32'h42f51bb4},
  {32'hc4e95410, 32'hc32c2e97, 32'h437ca473},
  {32'h44134c22, 32'hc3488ad8, 32'hc3601f21},
  {32'h427a03e4, 32'h428dff1f, 32'h4317f394},
  {32'h44ddd24e, 32'h433404b0, 32'hc1e907b0},
  {32'hc38492c5, 32'hc2f17192, 32'h41a46163},
  {32'h4441f665, 32'hc300069e, 32'hc3912b50},
  {32'hc50cbce5, 32'hc32e758e, 32'hc3269d39},
  {32'h444ff37a, 32'h43664079, 32'h428bc0a1},
  {32'hc4e8f82a, 32'h435fae28, 32'hc37c5588},
  {32'h44edee59, 32'hc2595ccc, 32'hc383ef4e},
  {32'hc4fd8458, 32'hc3c57969, 32'h426360f8},
  {32'h44dbd5ec, 32'hc26d0c79, 32'hc245e706},
  {32'hc47da37b, 32'hc369dfe8, 32'hc27d0da0},
  {32'h44e3ffa2, 32'h42521241, 32'hbdf22780},
  {32'hc470e5e0, 32'h432b9d1d, 32'h42eafa5c},
  {32'h44ac3c48, 32'hc393d677, 32'hc299f02e},
  {32'hc4696b24, 32'h43eccf12, 32'h412987db},
  {32'h42be5540, 32'hc291e0b3, 32'hc36b357c},
  {32'hc493c803, 32'h43bf97a2, 32'hc336d32d},
  {32'h450ce487, 32'h4385d4f7, 32'hc385aa26},
  {32'hc4e7c7a2, 32'hc29988c9, 32'h4386e464},
  {32'h44eefaa9, 32'h421d4a3e, 32'h42f3b283},
  {32'hc4fa8c30, 32'h4314dc21, 32'h43885957},
  {32'h4504ed07, 32'hc3634ef5, 32'h4359c39e},
  {32'hc4ed0cb2, 32'h435f1322, 32'hc3932e7f},
  {32'h4501dd74, 32'h43cc346d, 32'hc3c40e2a},
  {32'hc4cf6fad, 32'h419e8b4e, 32'h42b240f7},
  {32'h44465052, 32'hc38a2581, 32'h439af994},
  {32'hc4a6ffba, 32'h43729e6a, 32'h42b93bf6},
  {32'h441356dd, 32'hc30ddd84, 32'h43b1cedf},
  {32'h4147c730, 32'h428640fb, 32'hc3653637},
  {32'h44ea8a7c, 32'hc3e64d1c, 32'h43808bd7},
  {32'hc4c3f575, 32'hc337bd17, 32'h43471d40},
  {32'h450d683f, 32'h42fde0d7, 32'hc2b56ac5},
  {32'hc4e6e246, 32'h41bfcf1c, 32'h426415d6},
  {32'h44b9481e, 32'h42979a27, 32'h431416d5},
  {32'hc4508640, 32'hc357c1aa, 32'h4323fdcd},
  {32'h4514b9b3, 32'h42b69a46, 32'h4232ecc4},
  {32'hc50b7a1a, 32'h430caef8, 32'hc2c63077},
  {32'h44df7971, 32'h42b8cd95, 32'h4199b010},
  {32'hc453671d, 32'hc2696617, 32'hc339e2d3},
  {32'h443fa6ca, 32'h42b54cc9, 32'hc3809286},
  {32'hc502e97c, 32'hc22f1d46, 32'hc3ac71b7},
  {32'h444bd40b, 32'hc2a6b069, 32'h43813e4b},
  {32'hc35a8aa0, 32'hc2cb34cc, 32'h42b49a94},
  {32'h43a9822f, 32'h421ac84e, 32'h43354e5b},
  {32'hc4f7fb10, 32'hc321d365, 32'h42b44b4e},
  {32'h443dd321, 32'h41a75ca6, 32'h4337b69b},
  {32'hc4d062a1, 32'hc25d4acc, 32'hc384d86a},
  {32'h44adf083, 32'h431819b9, 32'hc22c5791},
  {32'hc49b35ee, 32'hc341cfc5, 32'hc34b2f8f},
  {32'h44add002, 32'h421468fa, 32'h42ca0530},
  {32'hc32c0304, 32'h43010ea9, 32'hc401e457},
  {32'h4518e8ad, 32'h4213bca9, 32'hc285eb55},
  {32'hc5156fcc, 32'h436a8418, 32'hc392205a},
  {32'h4508d0ad, 32'hc09414cc, 32'hc22468b8},
  {32'hc30e3167, 32'h43eaa393, 32'h438d996e},
  {32'h44018d76, 32'h4181ac8e, 32'h42aae9f1},
  {32'hc424c9c0, 32'h43a852bd, 32'h428a5ea3},
  {32'h442039e2, 32'hc2c38485, 32'h41d625f5},
  {32'hc446cda0, 32'h4302925d, 32'h43897d51},
  {32'h44d14130, 32'hc33d42bc, 32'h4343065a},
  {32'hc49de2b8, 32'h42b9c3e4, 32'hc3c9a2c0},
  {32'h451516f2, 32'h40dcd833, 32'hc3363915},
  {32'hc4f26ad5, 32'hc3df9ebb, 32'hc2e13029},
  {32'h445bf53c, 32'hc28a764b, 32'hc2e2bec4},
  {32'hc4adda08, 32'hc39a2549, 32'hc22f93d8},
  {32'h44773002, 32'hc39f28a3, 32'hc198f83c},
  {32'hc419176e, 32'h430697f1, 32'hc33091c4},
  {32'h44601532, 32'hc21fc57f, 32'hc3ed37e0},
  {32'hc31a31de, 32'h41e1e69a, 32'hc2a3429f},
  {32'h44a13ce1, 32'hc354904a, 32'h4325b24a},
  {32'hc50ff7b7, 32'h439214d4, 32'h41e5e78b},
  {32'h44a4fafd, 32'hc37ad176, 32'hc31c05eb},
  {32'hc4143294, 32'h42eb27a1, 32'h431e469f},
  {32'h43e1f88f, 32'hc2c7864a, 32'h435740d0},
  {32'hc414911a, 32'hc3901d77, 32'hc293afbd},
  {32'h44cfa4d2, 32'hc314b611, 32'hc295d6a2},
  {32'hc118d000, 32'hc2cef04e, 32'h43292728},
  {32'h450c571c, 32'h43563221, 32'h3f8d9ec8},
  {32'hc4634814, 32'h410b39fb, 32'hc3552e2a},
  {32'h44ebf9b8, 32'h4282b7d1, 32'h4386e398},
  {32'hc359ef50, 32'hc328c374, 32'hc2a0dd1e},
  {32'h4506c4ba, 32'h401ce55a, 32'h42da3dcd},
  {32'hc4efda2c, 32'h438ef03f, 32'h42751b5b},
  {32'h450713f0, 32'hc184e229, 32'h42a768cd},
  {32'hc4b7b8dc, 32'hc3567755, 32'hc36e1be0},
  {32'h44389e10, 32'h438f2a48, 32'hc24a33f6},
  {32'hc49aecb0, 32'hc3057baa, 32'hc334ad20},
  {32'h43b3f258, 32'h438b5154, 32'hc26d8174},
  {32'hc48733cf, 32'hc1f33a49, 32'hbf950afe},
  {32'h449b367c, 32'h43a35ada, 32'h42238466},
  {32'hc5045f6e, 32'hc3687212, 32'hc2a70b7c},
  {32'h44b374fd, 32'hc3715220, 32'h43710a57},
  {32'hc5150ccc, 32'h434568a7, 32'h43a0dca8},
  {32'h43284830, 32'hc2ec1b0b, 32'hc3931cfa},
  {32'hc48e0d4e, 32'hc27f3167, 32'hc2f19a38},
  {32'h44e8b77e, 32'h424d9877, 32'h42c96846},
  {32'hc40f83ef, 32'hc2a0e232, 32'h42fbf965},
  {32'h44a89db0, 32'hc310b9de, 32'h4384fcbc},
  {32'hc4b884db, 32'hc36cae50, 32'hc3047edb},
  {32'h43b6d5d4, 32'h436b2705, 32'h4408727c},
  {32'hc48bfe07, 32'h4321f97f, 32'h436756d5},
  {32'h44c01dc6, 32'h436b6b65, 32'h4383a1b6},
  {32'hc4557bf8, 32'h40cdca28, 32'hc3420100},
  {32'h43a9f0d7, 32'h43626405, 32'hc2e94731},
  {32'hc4457af9, 32'hc22120df, 32'h42dedaae},
  {32'h442d40a2, 32'h4224a296, 32'h421c2942},
  {32'hc4ebe2b6, 32'h430902ef, 32'hc2d90a33},
  {32'h44b4e791, 32'hc10320a8, 32'h428e4e6d},
  {32'hc5185126, 32'h440d4fc7, 32'h439ebc3a},
  {32'h44a36f3a, 32'hc34ef854, 32'hc3407e60},
  {32'hc4d829f0, 32'h4321ad54, 32'h4213625d},
  {32'h445a803c, 32'h43c07fcb, 32'hc1ec7130},
  {32'hc508cf00, 32'hc3523f03, 32'h4387c28a},
  {32'h4276a3c0, 32'h42c238ac, 32'hc3ad8e46},
  {32'hc4ae184f, 32'h4258645b, 32'hc19e0e5a},
  {32'h45073fb1, 32'h4312746c, 32'hc38a9943},
  {32'hc31a6570, 32'hc2a640b0, 32'hbff4bda0},
  {32'h4457bf24, 32'h44088456, 32'hc2e84316},
  {32'hc3d12fda, 32'h4224a132, 32'h42ecec43},
  {32'h447e4a3e, 32'h440ec896, 32'h4347db39},
  {32'h41acb140, 32'hc33f8bc6, 32'hc2cebcc6},
  {32'h448c92d0, 32'h42c9f7e2, 32'h437ee9d5},
  {32'hc4fb1d42, 32'h435c15e6, 32'hc35fe0ae},
  {32'h44e7c9c3, 32'hc2d4c61a, 32'hc25edff8},
  {32'hc3d6cc38, 32'h43543593, 32'hc3538cb4},
  {32'h431dab8a, 32'h43a97046, 32'hc1915ac8},
  {32'hc3ce3ea9, 32'h43d2109f, 32'h4345f24d},
  {32'h43c041a0, 32'h43c8bcba, 32'h4336c747},
  {32'hc325f55f, 32'h436dad6e, 32'hc1a8393f},
  {32'h44862c9f, 32'hc37cc634, 32'hc300b3e9},
  {32'hc409e1b1, 32'h438bea4a, 32'hc374e08c},
  {32'h44a6990e, 32'h43edf92d, 32'hc301d82c},
  {32'hc5172dd2, 32'h4273299c, 32'h43a20a3d},
  {32'h44505265, 32'hc335566d, 32'h43030623},
  {32'hc48ff299, 32'h42973353, 32'hc2ce905b},
  {32'h44773b99, 32'hc2e3b58a, 32'hc280996e},
  {32'hc4ebfcf5, 32'hc2a11549, 32'h4199c6b5},
  {32'h450fd0ce, 32'h42a21c51, 32'hc3a2f90f},
  {32'hc45a5f92, 32'h42e274a8, 32'hc1e85962},
  {32'h4423e190, 32'hc1a7879a, 32'h43bfa077},
  {32'hc48203f2, 32'hc3813812, 32'h44203732},
  {32'h44a510aa, 32'hc0bb03d0, 32'h4052c520},
  {32'hc4ffc09b, 32'hc36eaf9b, 32'h43975f60},
  {32'h44c857e3, 32'hc3a41872, 32'hc2bef3f3},
  {32'hc4585660, 32'h43b9c308, 32'h42766451},
  {32'h44fa18dc, 32'hbfa58750, 32'h439a0b7c},
  {32'hc4f5f3d7, 32'hc334c680, 32'h43a56a11},
  {32'h43f40e65, 32'hc3648a46, 32'hc2390e0f},
  {32'hc4e76472, 32'h4368b9e0, 32'hc17666dc},
  {32'h43c5565e, 32'h4316d706, 32'hc39266da},
  {32'h431fb620, 32'h4292f793, 32'hc350fc48},
  {32'h44bae8dc, 32'h42918aba, 32'h420f4b4b},
  {32'hc4ae7650, 32'h43dc63ae, 32'hc1e8b9b2},
  {32'h44bdecaa, 32'h41e9d2ff, 32'hc2b283fd},
  {32'hc3df5f08, 32'hc315f6b5, 32'hc13fdac8},
  {32'h44d3353f, 32'h42a76024, 32'hc1ede737},
  {32'hc4a5dde5, 32'hc40dae31, 32'hc3126fe8},
  {32'h44f29de6, 32'h42e311e2, 32'hc36456e3},
  {32'hc50bad6a, 32'h422f5de0, 32'h414b80b0},
  {32'h4430cc7c, 32'h429c5f9f, 32'hc384c71f},
  {32'h42e232a0, 32'h436b2b39, 32'h436e9d0e},
  {32'h44d59e73, 32'h42268e19, 32'hc25d396b},
  {32'hc4d33898, 32'hc371535e, 32'hc312d0b1},
  {32'h429881e0, 32'h432696fd, 32'h41dbdcfd},
  {32'hc4b6547a, 32'hc258f6a3, 32'h42df63c1},
  {32'h449315c5, 32'h42fd4d53, 32'h42478d8d},
  {32'hc50cf354, 32'h439f0a3f, 32'hc0866e1c},
  {32'h451a26cc, 32'h432ead40, 32'hc2c238ec},
  {32'hc4d7764b, 32'h41962bfb, 32'h427946bb},
  {32'h44ee52bd, 32'h414b6990, 32'h43a2b881},
  {32'hc4c1fcb6, 32'h428af4a7, 32'hc3a10645},
  {32'h4436a414, 32'hc221e0b2, 32'hc38b1cf4},
  {32'hc4fba53c, 32'hc40fd65e, 32'hc18b71a7},
  {32'h445e962e, 32'hc24045fd, 32'hc13f8e6c},
  {32'hc432360e, 32'h43154058, 32'h429b28bf},
  {32'h4426ce0e, 32'hc22cf645, 32'h43a58f0d},
  {32'hc5074bc3, 32'hc3c3c6f3, 32'h42ccbd66},
  {32'h44e3b00e, 32'h428c4544, 32'h41f2a1ca},
  {32'hc3b0f8a0, 32'hc39a076c, 32'hc3ae7e84},
  {32'h44d5b6d3, 32'hc37692c5, 32'hc3b85f78},
  {32'hc4b48325, 32'h4380398f, 32'hc3535338},
  {32'h440b5f4e, 32'h436879f1, 32'hc3357a49},
  {32'hc342e850, 32'h439f5daf, 32'hc33bd0b4},
  {32'h44fcb878, 32'h43b2f192, 32'h43528178},
  {32'hc4f47b00, 32'hc24c6a3e, 32'hc288ca33},
  {32'h4515133b, 32'h43010c66, 32'h43332415},
  {32'hc3ed5b3c, 32'hc3172ce6, 32'h42cf4ee6},
  {32'h44e417bc, 32'h429d3838, 32'h42a38300},
  {32'hc437c8d6, 32'h43689b36, 32'h43051fae},
  {32'h43491f6c, 32'h4309b9a0, 32'hc2e7631f},
  {32'hc4add43d, 32'hc34b4610, 32'h42465d30},
  {32'h44ad28e7, 32'hc33cd6a0, 32'hc2c1a5cc},
  {32'hc2d992dc, 32'hc3899c47, 32'h43b17e99},
  {32'h43f9373d, 32'h4371d182, 32'hc3517f4c},
  {32'hc436a946, 32'hc32e9d16, 32'h43d92b05},
  {32'h451e892d, 32'hc39b8205, 32'hc1ccd57f},
  {32'hc505cfa6, 32'h424c6a22, 32'h422d07d9},
  {32'h44f38df0, 32'hc318a01c, 32'hc390140f},
  {32'hc3f501d0, 32'h4407a6d4, 32'hc0888f04},
  {32'h44f0f589, 32'h432e402f, 32'hc229a20e},
  {32'hc5088c76, 32'h42f993d9, 32'hc15cd8ce},
  {32'h442f63c4, 32'hc30eba71, 32'h43ba2c9e},
  {32'hc4226b5e, 32'hc2bc5feb, 32'h4214848f},
  {32'h44ed13ac, 32'h419210e1, 32'h4383a974},
  {32'hc113f300, 32'h43f6424c, 32'hc3649b82},
  {32'h45035cca, 32'hc354b8fb, 32'hc36f7566},
  {32'hc4321b38, 32'h42e58d8c, 32'h4037bb7b},
  {32'h44a59952, 32'hc11cf291, 32'h42832769},
  {32'hc4d81815, 32'hc20ff7d0, 32'h43cb5bf8},
  {32'h43bbfef8, 32'h43ee70b3, 32'h4361bfcd},
  {32'hc4ec2c97, 32'h43040f79, 32'h4384eb96},
  {32'h44a51009, 32'h42aae0f0, 32'hc378d063},
  {32'hc50e03cb, 32'hc31baa0f, 32'hc212f3b5},
  {32'h442f6f5a, 32'h42577b96, 32'hc386bd8f},
  {32'h428a5906, 32'h429e69a6, 32'h43a0b943},
  {32'h43a03bb0, 32'hc34948e9, 32'h43945dcd},
  {32'hc4e568bd, 32'hc33c7db5, 32'hc384a415},
  {32'h44e9e004, 32'h42821a60, 32'hc35c12b2},
  {32'hc46a9bd5, 32'h430ec280, 32'hc349348e},
  {32'h43fc37b2, 32'h4386c7cb, 32'hc36304ca},
  {32'hc46e2c52, 32'h42fa81b8, 32'hc2239cb7},
  {32'h445aaccd, 32'h4118ff32, 32'h437977ec},
  {32'hc3aa23b8, 32'h432128de, 32'h42ea20ff},
  {32'hc17d3700, 32'h42a1706c, 32'h43967933},
  {32'h41924f00, 32'hc37fb6ea, 32'h42c5acd8},
  {32'h42e6d9c8, 32'h43a1665d, 32'h43aa3afa},
  {32'hc44dbd20, 32'hc2f8e352, 32'hc326e341},
  {32'h44351f99, 32'h41fd2425, 32'h43669e04},
  {32'hc4f8d98c, 32'h432c1cfd, 32'hc2adb5d2},
  {32'h44709d2c, 32'hc39954e4, 32'hc3c3fb51},
  {32'hc431fe9f, 32'hc1e698f0, 32'hc35ebfed},
  {32'h44a5845d, 32'hc2d74451, 32'hc382bf58},
  {32'hc506298b, 32'h42adf1ab, 32'hc3731030},
  {32'h44bd6202, 32'hc3019633, 32'hc343691e},
  {32'hc49e08d0, 32'h4318e71d, 32'hc24c0860},
  {32'h45059b30, 32'hc2ddd5b3, 32'hc38a254a},
  {32'hc3d171a4, 32'hc38e59b4, 32'hc3b65fe4},
  {32'h44a662da, 32'h42aaf20a, 32'hc37a4aa7},
  {32'hc4cdd962, 32'hc2b2a4dc, 32'hc2abb4fa},
  {32'h44ca0c36, 32'h43b1a4f7, 32'h4318c214},
  {32'hc3e858a8, 32'h43f15f62, 32'h42235f16},
  {32'h43e2c689, 32'hc321162a, 32'h43964893},
  {32'hc30d9980, 32'hc3032447, 32'h43434758},
  {32'h448e4db5, 32'h424443c8, 32'h43041688},
  {32'hc47c58e3, 32'hc3ae71b0, 32'h44346635},
  {32'h450bc1fb, 32'hc348e74f, 32'hc2bf9d6e},
  {32'hc42bb1fa, 32'h41d39aa4, 32'h42c208f9},
  {32'h44e8d889, 32'hc3b312c7, 32'hc23a5bec},
  {32'hc4f4e860, 32'hc3816498, 32'hc3702afc},
  {32'h44ec522a, 32'h42ce9c11, 32'hc4147e95},
  {32'hc4820876, 32'h3f6edf74, 32'hc39a2e6e},
  {32'h441489ef, 32'h42217468, 32'hc330a5f6},
  {32'hc4fadea4, 32'h42be60c4, 32'h4397a2ca},
  {32'h431cab20, 32'h3fbaf7c0, 32'hc3e7df5b},
  {32'hc2dd2398, 32'h42c2b083, 32'hc2e0fd41},
  {32'h439140fa, 32'hc32eb94c, 32'h43863091},
  {32'hc40fd353, 32'hc2f845df, 32'hc30774c4},
  {32'h446b6d0b, 32'h438e2f5b, 32'hc3194b2d},
  {32'hc50290c2, 32'hc1e10e68, 32'h4262df35},
  {32'h44818ac9, 32'h43135969, 32'h431ddec7},
  {32'hc47e729b, 32'hc3c29bd0, 32'h433dcdd2},
  {32'h450b45c9, 32'h43533b6a, 32'hc1d72047},
  {32'hc47fe1a2, 32'hc36e2633, 32'hc2911d3a},
  {32'h45042402, 32'hc36b34e2, 32'hc33ff33e},
  {32'hc48cdcd2, 32'hc3988df2, 32'h42a7f0b7},
  {32'h43c2c439, 32'hc3028c39, 32'h435b7d6b},
  {32'hc4bf7235, 32'h41a1f466, 32'h43695b0c},
  {32'h44e02dd4, 32'h43d06856, 32'hc4031096},
  {32'hc4adbe25, 32'h4314ae78, 32'h42890f64},
  {32'h44fbf414, 32'hc265a1dc, 32'hc32690c6},
  {32'hc4cd1e26, 32'hc369c339, 32'hc2cb6b8d},
  {32'h4506f667, 32'hc33bf5b5, 32'hc204d0eb},
  {32'hc4f59af8, 32'hc307719f, 32'h429fd1fb},
  {32'h4454db72, 32'hc2bba9b4, 32'h434d25c0},
  {32'hc3422096, 32'h4272be50, 32'h431bdcc7},
  {32'h4386fca4, 32'hc36d40ba, 32'h439bff64},
  {32'hc4a2bd88, 32'hc2285745, 32'h40ced3cc},
  {32'h446998f4, 32'hc3714fdc, 32'hc3753902},
  {32'hc4116e53, 32'hc18f90a7, 32'hc1caedc9},
  {32'h43fdbc4d, 32'hc30803bf, 32'hc1b55c92},
  {32'hc4b46759, 32'hc400a21e, 32'hc37a2e24},
  {32'h4468b666, 32'h439ab10b, 32'h420f034c},
  {32'hc3d66d33, 32'hc40a5fff, 32'hc34ac6e6},
  {32'h44f2b21a, 32'hc3aaee7a, 32'hc2e90df3},
  {32'hc4c85990, 32'h43a83b73, 32'h40ef107f},
  {32'h44822def, 32'h42f5f097, 32'hc32b4c1e},
  {32'hc42df550, 32'hc385aa74, 32'h435ff32b},
  {32'h44f7a55b, 32'h423dab50, 32'h431845fb},
  {32'hc4c2d573, 32'hc38e93b6, 32'hc30473b2},
  {32'h44f39c9a, 32'hc2b8b406, 32'h4339f9e5},
  {32'hc4540d92, 32'h4374382c, 32'hc1ec2052},
  {32'h451fd2c9, 32'hc414a023, 32'hc30db134},
  {32'hc4a498d3, 32'h435a0fdc, 32'hc383de09},
  {32'h451afdcd, 32'hc2e2dd55, 32'h43ab7dbd},
  {32'hc5053d20, 32'h42cced96, 32'hc3152f90},
  {32'h445f07b3, 32'h431e1f76, 32'hc178be7a},
  {32'hc4b459f1, 32'hc3c3b02f, 32'hc21c0f40},
  {32'hc3142168, 32'h42cbeb90, 32'hc3c3993b},
  {32'hc48a0224, 32'hc38f4bec, 32'hc28d5ed5},
  {32'h449a3efc, 32'h415d2376, 32'hc270c048},
  {32'hc50c9bfe, 32'hc2de6001, 32'h41cd8ee8},
  {32'h449481f6, 32'h405f7fd2, 32'h43783d9e},
  {32'hc47f1858, 32'hc33b3d8b, 32'h4297d079},
  {32'h43458210, 32'h425a172e, 32'h4324e312},
  {32'hc02c7000, 32'hc303f60c, 32'h43947404},
  {32'h45227ab4, 32'h42bb0734, 32'hc26d4f56},
  {32'hc491e5a8, 32'h41de883c, 32'hc317d69c},
  {32'h44c027f3, 32'h41a14222, 32'h41ae5fed},
  {32'hc4d6191d, 32'hc1e52b77, 32'h4136f702},
  {32'h4495ed66, 32'h4384f824, 32'hc232f7fe},
  {32'hc3bbd7f0, 32'h4417bafa, 32'hc365f42c},
  {32'h44948813, 32'hc1a9d050, 32'hc2b4e2d5},
  {32'hc4d11f8e, 32'hc2402d8c, 32'hc1b15595},
  {32'h44c2b8a4, 32'hc2c0fba9, 32'hc3b51624},
  {32'hc4d53744, 32'h4097f2ac, 32'hc3ad8081},
  {32'h44c7df2c, 32'hc29831c4, 32'hc0120b4c},
  {32'hc3eb88dc, 32'h431e822e, 32'hc3326d3d},
  {32'h44ad3d5e, 32'h43f22ceb, 32'hc2e95c36},
  {32'hc45d2ce4, 32'h42410e52, 32'hc3d1f43e},
  {32'h448e83b9, 32'hc3a3e276, 32'hc0b4f670},
  {32'hc4e50a48, 32'hc3ba843b, 32'hc244897e},
  {32'h442c5a78, 32'h4392298b, 32'hc3d39bc8},
  {32'hc494864e, 32'h43538ca4, 32'h416b8cff},
  {32'h45257497, 32'h4245fc60, 32'hc3675d27},
  {32'hc52094f0, 32'hc2a46398, 32'hc390ee20},
  {32'h44e02d93, 32'hc3446b12, 32'hc2f602f1},
  {32'hc51fdc07, 32'h436656ac, 32'h43bf660c},
  {32'h43d6b6f2, 32'h43283fa1, 32'h43912446},
  {32'hc4b0d155, 32'h4124aa32, 32'hc153ebf9},
  {32'h450c8bcc, 32'h424eda76, 32'hc3868ae8},
  {32'hc51d3e1f, 32'hc2511930, 32'h42f23e98},
  {32'h449d84d9, 32'h431d5210, 32'h4298d63d},
  {32'hc4946c57, 32'hc30e3e26, 32'hc126e045},
  {32'h4492de21, 32'h439f3cc0, 32'h415d3fc6},
  {32'hc5120fa4, 32'hc3650ebe, 32'h441a1579},
  {32'h44c0053d, 32'h43211084, 32'hc2886413},
  {32'hc4140630, 32'hc1cdd087, 32'h430fe92c},
  {32'h44892d6d, 32'h427909be, 32'h422f93bb},
  {32'hc485b58e, 32'h41a0cc76, 32'h43844977},
  {32'h4400648a, 32'hc3d5827c, 32'hc3aee632},
  {32'hc508de28, 32'hc37dd1b8, 32'h438f4c1e},
  {32'h440194b6, 32'hc1bcebdc, 32'hc22a00f4},
  {32'hc4152768, 32'h437c0aa1, 32'h43260584},
  {32'h445584b6, 32'h4204fcd3, 32'hc3aa725f},
  {32'hc391288e, 32'hc1b04575, 32'hc3ac43f9},
  {32'h451e474e, 32'hc38126aa, 32'hc1726b90},
  {32'hc4fa83cb, 32'hc246f541, 32'hc370261e},
  {32'h448ffa09, 32'h42c39716, 32'h4307f424},
  {32'hc4db0750, 32'hc2e42fb3, 32'h434a678b},
  {32'h4427be10, 32'hc25a82d6, 32'hc35b810c},
  {32'hc27e2480, 32'hc3ae5050, 32'hc23acd45},
  {32'h44fa6d42, 32'hc39288e0, 32'h43102ce6},
  {32'hc40b8ab4, 32'h428a2597, 32'hc33bb7e1},
  {32'h4429bcdc, 32'h43c4be5b, 32'hc28f686e},
  {32'hc44708ba, 32'hc24d040b, 32'h43052933},
  {32'h449a2f5e, 32'h422bfae1, 32'hc2951ad2},
  {32'hc3c46a20, 32'hc21094cc, 32'h4383d1b6},
  {32'h4356a38a, 32'hc26fbcec, 32'h43042567},
  {32'hc463344e, 32'hc16991ef, 32'hc3048516},
  {32'h43dea248, 32'hc2729605, 32'h430dd942},
  {32'hc4d31ad0, 32'hc2176eb3, 32'h42c75db8},
  {32'h4308c9d1, 32'hc3b607c8, 32'h42da0e59},
  {32'hc387be52, 32'hc3902e63, 32'hc30d765f},
  {32'h43888344, 32'h430c677c, 32'hc2983b54},
  {32'hc4038a43, 32'h427909b9, 32'h434ea58e},
  {32'h4516ca83, 32'hc3afed1e, 32'h439d074c},
  {32'hc41f2953, 32'hc3987fc7, 32'h4384006a},
  {32'h44f06359, 32'hc33a2a21, 32'h42d52162},
  {32'hc3b1a142, 32'hc2b853d1, 32'hc316bd01},
  {32'h44895e5c, 32'h43bca7c6, 32'hc350618d},
  {32'hc501a186, 32'hc312d920, 32'hc33e287f},
  {32'h44ab6e32, 32'hc3594e80, 32'hc32a2399},
  {32'hc4850522, 32'h430ef2c1, 32'h429a4e9c},
  {32'h4500dd5a, 32'h431f191b, 32'hc3077aa2},
  {32'hc4056e46, 32'hc248bb6e, 32'hc3129763},
  {32'h434946a8, 32'hc32bac7a, 32'h424387aa},
  {32'hc4e53560, 32'hc3af92b7, 32'hc3a7c9e0},
  {32'hc2c47ca8, 32'hc270c6f4, 32'h43158843},
  {32'hc4badde9, 32'h43c2c39d, 32'hc3b588d4},
  {32'h45004392, 32'hbe5c8f00, 32'h43e727d0},
  {32'hc4ee0450, 32'hc404a95b, 32'hc24dbf44},
  {32'h43dcbe72, 32'h438d1066, 32'h42419284},
  {32'hc4c71e53, 32'hc3d70885, 32'hc2e9009c},
  {32'h449a92bd, 32'hc2db4b15, 32'h432f0ca5},
  {32'hc30ed141, 32'hc2794ca9, 32'hc3ba968e},
  {32'h44198562, 32'h43c98be6, 32'h431dcb0f},
  {32'hc4979c7a, 32'h42594fce, 32'hc35dd655},
  {32'h44ddd7c2, 32'hc38155fd, 32'h43321a84},
  {32'hc46f0ccb, 32'hc382fa08, 32'h433ad2e9},
  {32'hc1393480, 32'h4137c904, 32'hc148ef00},
  {32'hc4645180, 32'hc31749f9, 32'h43494c93},
  {32'h44d0bef4, 32'hc2c737f8, 32'hc1c6a0b4},
  {32'hc4955945, 32'hc3ba89a5, 32'hc3a0d85f},
  {32'h44672106, 32'h42fbe28a, 32'h3f9cf9aa},
  {32'hc4a9e59b, 32'h4252d36c, 32'hc3e378ef},
  {32'h44d05343, 32'hc303ac98, 32'hc2aa5c30},
  {32'hc40cfe9a, 32'hc3d11710, 32'hc30647e4},
  {32'h440bf5e0, 32'h42abee44, 32'h4376343b},
  {32'hc4f6b426, 32'hc3d4d2e2, 32'h42cc1ac6},
  {32'h43f72190, 32'h42f80e45, 32'h4327664c},
  {32'hc4c1de55, 32'hc338b4a4, 32'hc2676104},
  {32'h42f936f4, 32'hc33955fc, 32'h43a492c5},
  {32'hc1e325c0, 32'hc30c0950, 32'hc37aa527},
  {32'h44fd4d82, 32'hc352b704, 32'h424b1a45},
  {32'hc4a66884, 32'hc40e2bc6, 32'hc3919432},
  {32'h44d3fed2, 32'hc35f5ce9, 32'h41d33993},
  {32'hc483e23d, 32'hc30fed31, 32'hc37eaac5},
  {32'h4481181e, 32'hc365c604, 32'hc37d1d82},
  {32'hc485bb57, 32'hc292a69e, 32'hc3814355},
  {32'h43389610, 32'hc39e85c8, 32'hc4003581},
  {32'h44f19b42, 32'h43555945, 32'hbfd71043},
  {32'hc40d4a14, 32'hc3aed735, 32'h4384a4f4},
  {32'h45197622, 32'h43323dbe, 32'h43ce7320},
  {32'hc4cd22bc, 32'h43e538bf, 32'hc331109a},
  {32'h44bfeda6, 32'h4245f0c4, 32'h4405a020},
  {32'hc274d03c, 32'hc3ac9f1c, 32'hc425b5a2},
  {32'h4379a648, 32'hc2bb7e4f, 32'h428b344f},
  {32'hc40c770e, 32'h42f7489f, 32'hc284734f},
  {32'h44858f2c, 32'h43075e23, 32'hc399cc5d},
  {32'hc4f7b8c0, 32'h42c2bfb8, 32'hc3ee53df},
  {32'h44b5ee4c, 32'h431f7783, 32'h4379b1e6},
  {32'hc50208f4, 32'hc21012e3, 32'hc33c7483},
  {32'h44fb2686, 32'h43a9c88b, 32'h4380df09},
  {32'hc3c364b4, 32'h422e17d0, 32'h42159f05},
  {32'h44afdeb4, 32'hc3276512, 32'h428be908},
  {32'hc4accc7b, 32'hc27bed26, 32'hc32b9cbe},
  {32'h438afdb1, 32'hc3100154, 32'h439579d4},
  {32'hc47b9f30, 32'h42c45b89, 32'hc3cc82ca},
  {32'h4357bf0c, 32'h42b843fa, 32'hc2bbde3e},
  {32'hc4252448, 32'hc32ffa01, 32'hc2727a55},
  {32'h44aa51b6, 32'hc14854de, 32'h4335647e},
  {32'hc2aa54ce, 32'h420e80ec, 32'hc2d9d1ee},
  {32'h435661a1, 32'h41db8190, 32'hc1ae82da},
  {32'hc482f1be, 32'h433b9e19, 32'h42e029ba},
  {32'h44c033e4, 32'hc24ae4ac, 32'hc1f75789},
  {32'hc392faf8, 32'hc2f6fc79, 32'h42186e9c},
  {32'h43d29e88, 32'hc1fe9250, 32'h4371b906},
  {32'hc4cc40c9, 32'h409522ca, 32'h427dfd6f},
  {32'h444c912a, 32'hc161891b, 32'h438d8268},
  {32'hc4c4db32, 32'h431248e7, 32'h42ae9d49},
  {32'h4314b650, 32'h434a4b53, 32'h43bc3189},
  {32'hc4a1b4fe, 32'h42da4128, 32'hc3a5906a},
  {32'h430edc14, 32'h4324136c, 32'h424584e9},
  {32'hc4fb74be, 32'h436e8fde, 32'hc3800fbc},
  {32'h450fe796, 32'h439092d8, 32'h43627171},
  {32'hc4c0081d, 32'hc2a267b6, 32'hc298b26a},
  {32'h45020f4c, 32'hc2068293, 32'hc229c7ec},
  {32'hc414bc70, 32'hc29d5f96, 32'h42f29e2f},
  {32'h44eec9fe, 32'hc336d777, 32'h42fc4797},
  {32'h41ba8780, 32'hc33a3ba8, 32'hc331f765},
  {32'h44b5c8e1, 32'hc2bd589b, 32'hc13d700b},
  {32'hc4fe9051, 32'hc1c332d4, 32'h43515cf4},
  {32'h450df816, 32'hc30a2f6b, 32'hc28266f2},
  {32'hc3f6042c, 32'hc330fe5c, 32'h4144334c},
  {32'h448cf0c1, 32'h4365ec87, 32'h43193c30},
  {32'hc48ad596, 32'hc2ad1d59, 32'hc3782011},
  {32'h4508aff8, 32'hc2c999d6, 32'h41e3438e},
  {32'hc49bae7e, 32'h438aa8b2, 32'h411dba4e},
  {32'h43d169db, 32'hc2102714, 32'h420209d2},
  {32'hc406019e, 32'h43da79a0, 32'hc367ee7c},
  {32'h43792300, 32'h42338475, 32'hc382cd2d},
  {32'hc4aaa5e9, 32'hc15ea8b6, 32'hc3261fd5},
  {32'h42aae8dd, 32'hc388d853, 32'hc3a36d77},
  {32'hc31db844, 32'hc1cce616, 32'hc243ab51},
  {32'h43facab0, 32'hc3aad417, 32'hc2c73aa9},
  {32'hc4f70662, 32'hc2830752, 32'hc3c12463},
  {32'h4483513a, 32'h4246645c, 32'hc187b60d},
  {32'hc4951821, 32'h43d20c57, 32'hc3b6e38e},
  {32'h43713794, 32'hc4026bc0, 32'h43faf2b2},
  {32'h42fa2420, 32'hc3281399, 32'hc3920efa},
  {32'h44dd4f36, 32'hc28db0cb, 32'hc37b35d7},
  {32'hc4bbeea7, 32'hc250b648, 32'hc41e0c6c},
  {32'h44fbfc8d, 32'hc2d81d5f, 32'h43af114f},
  {32'hc4e24750, 32'h41bedb6f, 32'h43aaf711},
  {32'h44b005ac, 32'hc43b9bf5, 32'h42a23232},
  {32'hc4cefe65, 32'hc26e941f, 32'h42bcc636},
  {32'h443b0cf3, 32'h40a49524, 32'h431c9439},
  {32'hc50f3022, 32'h41707eb5, 32'hc3840a69},
  {32'h43c351bc, 32'hc370b8ca, 32'h443cdf93},
  {32'hc41deb86, 32'hc32986ac, 32'h41ca64e6},
  {32'h44c0bde2, 32'hc29405b2, 32'h43460947},
  {32'hc4cc0653, 32'hc3cbec68, 32'hc2d1fc22},
  {32'h442271c0, 32'hc2bbecb0, 32'h432d92c2},
  {32'hc51c8efc, 32'hc31e77f4, 32'hc2f6528e},
  {32'h43c34f06, 32'h43890839, 32'h43eb5a50},
  {32'hc5004ac7, 32'h4347cf45, 32'hc39036a0},
  {32'h45158f57, 32'hc12b18f8, 32'hc3d30878},
  {32'hc4f2b466, 32'hc36843d9, 32'hbfa303c8},
  {32'h4514c57a, 32'h43eb981b, 32'h43bfa967},
  {32'hc513eace, 32'h432f3f39, 32'hc2b7ad96},
  {32'h450b006e, 32'hc3b0b89a, 32'h43cc7887},
  {32'hc34f127c, 32'h434a502c, 32'h436477bc},
  {32'h44d1f323, 32'h415cb9a6, 32'hc3b0eacf},
  {32'hc4072598, 32'hc3caa259, 32'h439d3c0e},
  {32'h437436b8, 32'h40e7f16d, 32'h41293be5},
  {32'hc44bea52, 32'h436677d6, 32'hc2e13c24},
  {32'h450e14ee, 32'h420b8eca, 32'hc3753488},
  {32'hc30e8b8c, 32'hc2e223d3, 32'h43fe1973},
  {32'h43dd954b, 32'hc2caef82, 32'h42c592cc},
  {32'hc4287dc6, 32'hc3b4e580, 32'hc298cf2e},
  {32'h430102e6, 32'h43081de5, 32'hc2904518},
  {32'hc4ee3480, 32'hc2bc07be, 32'hc3ca77e6},
  {32'h44c24aed, 32'hc0a79b18, 32'h43eb8d3e},
  {32'hc493bd29, 32'hc201c79c, 32'hc3becdd5},
  {32'h449d8086, 32'hc37031dc, 32'hc29da7e3},
  {32'hc4d96d0c, 32'hc2ad1044, 32'hc3018016},
  {32'h4433fcbc, 32'h4344a446, 32'hc3286c2f},
  {32'hc4bd6a30, 32'hc37b887b, 32'hc397ef15},
  {32'h4505f72f, 32'hc2b79703, 32'hc2d03b82},
  {32'hc26e5823, 32'hc1f6b5b0, 32'h42baa87f},
  {32'h44c54389, 32'hc27fa957, 32'hc2d050f2},
  {32'hc4251710, 32'hc35071d4, 32'h430a5b53},
  {32'h4502c193, 32'h431deb39, 32'h4398a1a0},
  {32'hc431cd50, 32'hc13fe442, 32'hc302f81e},
  {32'h4494f9f2, 32'hc3546cb7, 32'h41c16cef},
  {32'h43672a5c, 32'hc287e3d6, 32'hc2d86747},
  {32'h449dbda9, 32'hc2a78a30, 32'h418e1906},
  {32'hc48050d7, 32'hc26208a5, 32'h430e9c5a},
  {32'h45195134, 32'h42fdcf66, 32'hc3f00742},
  {32'h4355ab0a, 32'hc31cb5c5, 32'hc3e0b915},
  {32'h44584130, 32'hc289209c, 32'h431229ca},
  {32'hc4d636fb, 32'h437f4322, 32'hc391b778},
  {32'h4507b0cd, 32'hc391fc09, 32'h4300ddfb},
  {32'hc2428300, 32'hc2fc3f92, 32'h435be48b},
  {32'h451cd6dc, 32'h43c50f58, 32'hc243b517},
  {32'hc48c6caa, 32'hc19abe20, 32'hc2e8de21},
  {32'h439a0240, 32'h41ae99d4, 32'h41f53ba0},
  {32'hc4f3f616, 32'h43737f55, 32'h438e7b6e},
  {32'h451e4984, 32'hc41f9512, 32'h4208177c},
  {32'hc4d8a908, 32'hc2b74bbb, 32'h43ebbba2},
  {32'h450b3dc0, 32'h4319579d, 32'hc3e495a2},
  {32'hc22cbb10, 32'hc37af3c6, 32'hc2183f48},
  {32'h43f37948, 32'hc30d8a25, 32'hc2d4a977},
  {32'hc4cc3114, 32'h4408a03b, 32'hc271e384},
  {32'h450b5a5c, 32'hc2cc1c30, 32'h438b273c},
  {32'hc4634920, 32'hc2cf325f, 32'h438b4b3a},
  {32'h447ca58d, 32'hc385e1cd, 32'h43082c28},
  {32'hc4f43294, 32'hc2a696a3, 32'h421f20aa},
  {32'h44df35e8, 32'hc336821d, 32'hc3607ab6},
  {32'h432e3630, 32'h43cbf4a6, 32'hc2a8449a},
  {32'h42aa15e0, 32'hc27028e6, 32'h4336fd2b},
  {32'hc28e0c27, 32'h43e73f74, 32'h4389dd5e},
  {32'h44516f69, 32'hc2579c36, 32'hc301b751},
  {32'hc4e55ada, 32'h44169477, 32'h4359232d},
  {32'h453ed515, 32'h43e1e63e, 32'hc29d8572},
  {32'hc4955e24, 32'h422dd430, 32'h43809906},
  {32'h4506bb70, 32'hc313c0b4, 32'h43348107},
  {32'hc4ffd5b2, 32'hc31aee44, 32'h43873dbb},
  {32'h44df7dc7, 32'h43bc1d7a, 32'hc34c0760},
  {32'hc436cbc4, 32'hc36e1bf7, 32'h419c4503},
  {32'h446c8f9e, 32'hc30115d5, 32'hc39ad820},
  {32'hc51f8337, 32'hc1dab371, 32'hc2855ea0},
  {32'h441d51c4, 32'h43aaa1f3, 32'hc29c2fb7},
  {32'hc480cce4, 32'h434a9154, 32'h43d4b3d6},
  {32'h448d5fd4, 32'h429035f3, 32'h4245ff43},
  {32'hc44fc4c8, 32'hc401ca9c, 32'hc2190fd9},
  {32'h44511250, 32'h42b15247, 32'hc21e85f8},
  {32'hc272dc20, 32'h42066074, 32'h42a06924},
  {32'h44a57016, 32'hc1950524, 32'h421ff789},
  {32'hc48e7559, 32'hc38b8021, 32'h42d7045a},
  {32'h43c05804, 32'hc388330d, 32'hc391ede2},
  {32'hc4f0e778, 32'h43260c25, 32'hc0e74dc4},
  {32'h44d02896, 32'hc25ee279, 32'hc38a12a2},
  {32'hc4251c26, 32'h438a0cc6, 32'hc364c5e8},
  {32'h43cf78d6, 32'h43449a6e, 32'h43612c10},
  {32'hc45c58e4, 32'h43967bdc, 32'hc3b21572},
  {32'h44ca1a5a, 32'hc3538e52, 32'h4315eb92},
  {32'h4374f37f, 32'h42eb0d54, 32'h42fc5a56},
  {32'h42733800, 32'h438c4028, 32'hc3e51df1},
  {32'hc4cb0e84, 32'h4218ca6f, 32'h437dbae8},
  {32'h44eb49ce, 32'hc1b511ab, 32'hc08e63e0},
  {32'hc3ff86bc, 32'hc3766dbc, 32'hc33c1607},
  {32'h44974daa, 32'hc3bf5d2a, 32'h429a0963},
  {32'hc422d7d4, 32'hc2a8394e, 32'h43478615},
  {32'h44c9859a, 32'hc34895c2, 32'hc0827914},
  {32'hc3a88f20, 32'hc29fe2f5, 32'hc1b52a04},
  {32'h4470c810, 32'h4317019e, 32'hc36d5f14},
  {32'hc3a92f6e, 32'hc308eaec, 32'h425467bb},
  {32'hbfabb500, 32'hc367efb5, 32'h4326baa3},
  {32'hc41af30a, 32'hc2bb095f, 32'h42bf441f},
  {32'h44678393, 32'hc39f819e, 32'hc2fcff92},
  {32'hc4cf33c2, 32'hc36aa517, 32'hc291a609},
  {32'h448a6d52, 32'h439efd5d, 32'hc31e890e},
  {32'hc4d3ce10, 32'hc3bc48cf, 32'hc3156fb4},
  {32'h446844d4, 32'hc3675918, 32'hc3890c04},
  {32'hc4cfa84f, 32'h439c32ec, 32'h43ee70dd},
  {32'h43ca0760, 32'hc32b933f, 32'h42a5d717},
  {32'hc4b8b9cf, 32'h4366fdba, 32'hc3cdfad5},
  {32'h4502df89, 32'hc3474eb3, 32'hc21327d9},
  {32'hc40d903d, 32'hc3699c08, 32'h42ed04e7},
  {32'h438d11d0, 32'hc29386b4, 32'hc2a6f5f5},
  {32'hc450847a, 32'hc3041f1a, 32'h44121837},
  {32'h44a5beb0, 32'h43891fc8, 32'hc14e30e8},
  {32'hc4f47ea2, 32'hc30c6ef4, 32'hc3022030},
  {32'h44198276, 32'hc30dd646, 32'h438135ea},
  {32'hc49bd219, 32'hc31e7e6a, 32'h430d7d32},
  {32'h429e43f7, 32'h43d9302c, 32'hc20a3e7a},
  {32'h4309c1ae, 32'hc2a1bde7, 32'h4394a922},
  {32'h4517fc99, 32'hc35d6cd0, 32'hc3113d7a},
  {32'hc3322d10, 32'h42a9cec0, 32'h43a159e4},
  {32'h43db2a38, 32'hc22ac64f, 32'h4373d7ae},
  {32'hc47efbb6, 32'hc31ad16a, 32'h43bfb9e2},
  {32'h44fcb0fc, 32'hc27a87d5, 32'h4313b818},
  {32'hc4d35858, 32'h4318e7b7, 32'hc39665cb},
  {32'h44b82b06, 32'h42e7e088, 32'h4389c325},
  {32'hc496c275, 32'h432d81a2, 32'hc360b850},
  {32'h450df7ad, 32'h43a6a569, 32'h42cef070},
  {32'hc342fdca, 32'h43ac57d0, 32'hc282e8cb},
  {32'h43fe9e0a, 32'hc310f1e1, 32'hc31e7353},
  {32'hc186f850, 32'h413d5edd, 32'h43717369},
  {32'h44135d40, 32'hc2e0954f, 32'h415d3f60},
  {32'hc47a43b0, 32'hc236905f, 32'hc286e91a},
  {32'h44bbebde, 32'h42b7e6b6, 32'h42c1439a},
  {32'hc41caab0, 32'hc31ccd86, 32'h43df25ce},
  {32'h4349c888, 32'h43930906, 32'h438376b6},
  {32'h4043dc00, 32'h440d3154, 32'h42b593b8},
  {32'h451281aa, 32'h42af9c7c, 32'hc22a635c},
  {32'hc4c1f433, 32'h4332031d, 32'hc39c85b4},
  {32'h445bce66, 32'hc34d7c3e, 32'h4359fca7},
  {32'hc3827ef0, 32'hc2c5e8f8, 32'h43baa875},
  {32'h44650976, 32'h4386fdaa, 32'h4246e443},
  {32'hc4b2d6a4, 32'hc259f91a, 32'h431798c9},
  {32'h42fac778, 32'hc3ff55bc, 32'hc26e4acd},
  {32'hc4fcbb7d, 32'hc1c43436, 32'hc0bf7808},
  {32'h44e1571c, 32'hc390d7da, 32'hc3c134f3},
  {32'hc28e07c4, 32'hc3851b78, 32'hc3842cbe},
  {32'h44ebefa3, 32'hc32f665f, 32'hc3ae84b8},
  {32'hc4b6b144, 32'hc35a81f8, 32'h42a9df2b},
  {32'h44b9e050, 32'hc0dda4c1, 32'h43830935},
  {32'hc3b23528, 32'hc3b9c2f1, 32'h41ff3b0f},
  {32'h44dd051a, 32'h42346844, 32'hc2d8fcfd},
  {32'hc50fd229, 32'hc182a639, 32'h43b5374f},
  {32'h43e1f7c0, 32'h43621fe6, 32'h42b2b1d4},
  {32'hc44068d8, 32'h433a02cc, 32'hc2f29864},
  {32'h435b38d2, 32'h435d1567, 32'hc37c860c},
  {32'hc4d114ad, 32'hc2c25ad6, 32'hc36db698},
  {32'h44bb8caf, 32'h442d8cba, 32'hc32a1def},
  {32'hc4a800b6, 32'hc43f56ac, 32'h43c1204b},
  {32'h452801bc, 32'h430cdcd4, 32'hc2ea20ac},
  {32'hc46304a3, 32'hc2af25ce, 32'h44092c47},
  {32'h450eecfc, 32'h437f46c9, 32'h437f4155},
  {32'hc50cec5d, 32'h402d2fad, 32'hc19f10d8},
  {32'h44cfcd3e, 32'hc317b3a4, 32'h432843be},
  {32'hc50673cd, 32'h41e4ff13, 32'h43360c99},
  {32'h44d55b46, 32'h43de1a56, 32'h4386c133},
  {32'hc4c4ed16, 32'h418a9ab0, 32'hc2c90dc0},
  {32'h42fecfd0, 32'hc28756d8, 32'h436c2b2f},
  {32'hc4b05712, 32'hc347ecc6, 32'h42870a4a},
  {32'h44af5b75, 32'h420a67eb, 32'hc34a8f03},
  {32'hc3ac5e76, 32'hc2b509a6, 32'h4345b7e4},
  {32'h4430db75, 32'h424a3062, 32'hc2c96c68},
  {32'hc4affc3a, 32'h429b9a3f, 32'h431e7fc9},
  {32'h443a4014, 32'h431b229f, 32'h40642029},
  {32'hc419e7bc, 32'h43c61329, 32'h4363058d},
  {32'h441a2bb5, 32'h439a4a69, 32'h43cad873},
  {32'hc4969fe3, 32'h42495155, 32'h42814094},
  {32'h44d4ce9e, 32'hc31887e2, 32'h4329c9c3},
  {32'hc4f5f596, 32'hc314ff03, 32'h435555fb},
  {32'h4445bcf4, 32'h435c01cf, 32'hc307fbd8},
  {32'hc444e222, 32'hc38e945a, 32'h434e856a},
  {32'h448f956f, 32'h430ca0a7, 32'h425ae4dc},
  {32'hc32f3890, 32'h4319ad12, 32'hc211d5c8},
  {32'h45154785, 32'h43501b2a, 32'hc2c891f5},
  {32'hc40d15e4, 32'hc388a3fe, 32'hc1110852},
  {32'h4486a296, 32'h4383653a, 32'hc3a75309},
  {32'hc2c489f0, 32'hc3d24b56, 32'h435cb220},
  {32'h44360f0f, 32'h43c17e8b, 32'hc2dca219},
  {32'hc4ff336e, 32'h427263a8, 32'hc15523de},
  {32'h43aa9fc6, 32'h42654380, 32'h41b8e419},
  {32'hc48464bc, 32'hc2484e8a, 32'hc20eb132},
  {32'h44a89f62, 32'h4357668a, 32'hc34e4b49},
  {32'hc505fbd4, 32'h41e89610, 32'hc15d5837},
  {32'h45024ea7, 32'h4307bc72, 32'hc25ec052},
  {32'hc4996fad, 32'hc2de42f7, 32'hc3505dcd},
  {32'h44f2109c, 32'hc3927da5, 32'h4382c248},
  {32'hc4844646, 32'hc2809099, 32'hc382ab88},
  {32'h44b9c6d8, 32'h436ca66d, 32'hc34c87ef},
  {32'hc49bdd92, 32'hc31d358a, 32'hc3940dff},
  {32'h4510bf0d, 32'hc332429c, 32'hc42c9012},
  {32'hc4d65e62, 32'h42bb62fe, 32'hc2b24f64},
  {32'h446c5e76, 32'h430d56bd, 32'hc31748e6},
  {32'h42314392, 32'h42f20bc3, 32'h433dff5f},
  {32'h44665e00, 32'h4348b739, 32'h43692ec3},
  {32'hc19fd02c, 32'hc40837c3, 32'hc3df5a7f},
  {32'h445e542e, 32'h4269e6ec, 32'hc0dfc9c9},
  {32'hc46ea550, 32'h41df37b5, 32'h4376c01e},
  {32'hc2b475d0, 32'hc2b4f0d6, 32'h43a02247},
  {32'h42690340, 32'h438d0603, 32'h42858f63},
  {32'hc327aafc, 32'h43034396, 32'h4310fc45},
  {32'hc39d07a0, 32'h437bdc57, 32'h43ab67ec},
  {32'h451873aa, 32'h43957de2, 32'hc3a51abd},
  {32'hc44e2652, 32'hc2f712a0, 32'h42270836},
  {32'h4119bb00, 32'hc2c282e7, 32'hc2d6bec8},
  {32'hc504b152, 32'h42aa6f9f, 32'h43876b6e},
  {32'h448d5620, 32'h42b8bf8e, 32'hc374afc8},
  {32'hc44fb520, 32'h43d10cbf, 32'h40e07b66},
  {32'h450c0ff6, 32'h43c1afe3, 32'hc3072b8a},
  {32'hc414fab8, 32'h42830016, 32'h4032f005},
  {32'h44e56780, 32'h43509fbb, 32'hc3895106},
  {32'hc495b361, 32'hc235382c, 32'h418c7100},
  {32'hc1332b80, 32'h440f486a, 32'h41c724df},
  {32'hc4e10edb, 32'h43189af6, 32'hc372116a},
  {32'h441d39e8, 32'h428f76ae, 32'hc22403c5},
  {32'hc42a0d18, 32'hc1d2b9bb, 32'hc32d121f},
  {32'h44e253e8, 32'hc1908d97, 32'h430a318b},
  {32'hc4bfba4a, 32'hc08285c8, 32'hc31e5ef0},
  {32'hc17f8800, 32'h439bcbea, 32'h430ec06e},
  {32'hc510bae8, 32'h42be04e7, 32'h415241a5},
  {32'h44a0f730, 32'hc3493934, 32'h43732f75},
  {32'hc500b0d5, 32'hc3c1a9cd, 32'hc0b86c50},
  {32'h44aeaa7d, 32'hc2d16e75, 32'hc3b5e5e6},
  {32'hc4465002, 32'hc3791b29, 32'h434371a8},
  {32'h43cea818, 32'h42843c8c, 32'h4287c698},
  {32'hc4971f33, 32'h436074ee, 32'hc3df46ff},
  {32'h44d00d37, 32'h4303b035, 32'hc1414f88},
  {32'hc496698b, 32'h423ab376, 32'hc3526a73},
  {32'h448966e3, 32'h41c332f5, 32'hc399b47e},
  {32'hc481ff26, 32'h42bf52cf, 32'hc298c67e},
  {32'h44e939df, 32'hc2a89685, 32'h432aa6ae},
  {32'hc3a02106, 32'hc3f7207b, 32'h4362e74e},
  {32'h438beaec, 32'h4202ef6c, 32'h42e602da},
  {32'hc3ce96f8, 32'h432595e4, 32'hc2271f35},
  {32'h4500fd05, 32'hc27bafe2, 32'h42a991c3},
  {32'hc45cda24, 32'h43c8992f, 32'h4398c2fb},
  {32'h44de8b68, 32'h43a25637, 32'hc1faa04e},
  {32'hc3e859d2, 32'h436b3bad, 32'h439fb396},
  {32'hc3417167, 32'hc356df8d, 32'h425fb772},
  {32'hc4e079da, 32'h41d9d674, 32'hc25ce0a6},
  {32'h44542af2, 32'hc3b4f680, 32'h4386b39b},
  {32'hc4c909ad, 32'h43c84a1c, 32'hc35be37e},
  {32'h44ea0d57, 32'hc3b99d17, 32'h438c0a73},
  {32'hc399f5a0, 32'h42b5357a, 32'hc0bacb1a},
  {32'h4433e990, 32'h43d18be5, 32'h43d4117e},
  {32'hc4a4ba5b, 32'h434d73e1, 32'hc31cbbc2},
  {32'h43d46a3a, 32'h42c939ab, 32'h43d0e970},
  {32'hc3641912, 32'hc3efbf83, 32'h43da6246},
  {32'h44d8a1be, 32'h43b00df3, 32'hc2c84f52},
  {32'hc2c32570, 32'hc376e687, 32'hc1e6e9d7},
  {32'h44645c40, 32'h432d586a, 32'hc3667dae},
  {32'hc45fac2c, 32'hc395e2c8, 32'h42b1cc3d},
  {32'h451b7418, 32'h43616cf9, 32'h4273963f},
  {32'hc45c8182, 32'h436d6ba0, 32'h42995820},
  {32'h44289601, 32'h42c35dff, 32'hc220f3a8},
  {32'hc4ebcb4a, 32'h432e3ffe, 32'hc2f23ec1},
  {32'h44a20bb8, 32'hc2f8baec, 32'h404b75b7},
  {32'hc4c50f2e, 32'h43c15000, 32'h42dbdc77},
  {32'h44fb66ba, 32'hc217ea0c, 32'hc319b7ff},
  {32'hc44af90f, 32'hc3c5ed17, 32'hc3c3f06a},
  {32'h451a550c, 32'h43d3b508, 32'hc288cba0},
  {32'hc43a44a2, 32'h42f0cd0e, 32'h411035b8},
  {32'h44ee7f02, 32'hc2b7f359, 32'hc29eb282},
  {32'hc3a973d5, 32'hc3369443, 32'h438c6101},
  {32'h44f9e146, 32'h42a4ed10, 32'hc3188c22},
  {32'hc4dca9d5, 32'h42a393e1, 32'hc21cb9a9},
  {32'h4501f6c7, 32'h4398da45, 32'h438b9fc7},
  {32'hc46443ce, 32'hc2f9dd27, 32'hc2d426ea},
  {32'h450ffc13, 32'hc0cb8b3b, 32'hc32d3f69},
  {32'hc48722dc, 32'hc19e199b, 32'hc3dfbc6e},
  {32'h45005eae, 32'h42d5108d, 32'h409fb45e},
  {32'hc32d325b, 32'hc3b50364, 32'h439e4dda},
  {32'h44b3fcab, 32'h438ecc8b, 32'hc1bc294b},
  {32'hc518a52b, 32'hc2b4deae, 32'hc415718c},
  {32'h451298fa, 32'h4302c628, 32'hc286030c},
  {32'hc5141608, 32'h41b3ca8a, 32'hc3846583},
  {32'h448c4549, 32'hc23b8bec, 32'hc2f72926},
  {32'hc4cad475, 32'h43cc7f79, 32'h424a6748},
  {32'h43818b80, 32'hc35c17f7, 32'hc3170d4e},
  {32'hc4e651be, 32'h43d1fba8, 32'hc25d43fd},
  {32'h45157f10, 32'h43086162, 32'h41e521ea},
  {32'hc504fa84, 32'hc38a0944, 32'h4195f0e3},
  {32'h44b4fa6d, 32'hc33133da, 32'h43559cec},
  {32'hc4168c08, 32'hc27f2791, 32'hc24058b5},
  {32'h44b8e5e9, 32'h43014025, 32'hc3917064},
  {32'hc501b4ad, 32'h42af3588, 32'h4374c406},
  {32'h426c1818, 32'h4385768e, 32'hbea550b1},
  {32'hc27da420, 32'h42d2ac94, 32'h44091011},
  {32'h4433d761, 32'hc27f272b, 32'hc2f3744e},
  {32'hc5294460, 32'h43453ae6, 32'hc3346880},
  {32'h44cba5dc, 32'hc0cef0ea, 32'h43339111},
  {32'hc4bd7eec, 32'h43ecca42, 32'h4372d24f},
  {32'h434aa800, 32'h421d7e9b, 32'hc36db15a},
  {32'hc4326761, 32'h42fd5d41, 32'h428dd8a0},
  {32'h44ef3ca7, 32'h439ce6dc, 32'h415cab04},
  {32'hc444f47a, 32'h43846a2c, 32'hc2b581ea},
  {32'h450fc3f4, 32'h4343b2ef, 32'h43c6ffad},
  {32'hc499cfd7, 32'hc1d250e4, 32'h439cb7bb},
  {32'h44f385ed, 32'h42bae5d1, 32'hc2918163},
  {32'hc37e1f3b, 32'hc373f843, 32'h434024ef},
  {32'h44e90939, 32'hc253e4aa, 32'hc34a2979},
  {32'hc454738e, 32'h4385d617, 32'hc381a3e3},
  {32'h45236907, 32'h43a47804, 32'h42969bec},
  {32'hc4a57dda, 32'hc2e6455d, 32'hc328f4cc},
  {32'h44a6b517, 32'hc297d159, 32'h43042b33},
  {32'hc4f18132, 32'hc2bedff2, 32'h43985135},
  {32'h44399414, 32'hc39b18be, 32'hc317df1e},
  {32'hc45699a4, 32'h42ea7731, 32'hc341e91d},
  {32'h44b30320, 32'h43d719af, 32'hc3b200d8},
  {32'hc4d586dc, 32'h4082132e, 32'h4433241b},
  {32'h43cd5d0c, 32'h43309058, 32'hc2f59cd2},
  {32'hc3ac941c, 32'hc2dec7b5, 32'h420dbf8a},
  {32'h44cf684c, 32'hc21a0d2c, 32'hc3a086da},
  {32'hc3e3a080, 32'h430d00c0, 32'hc3994dcd},
  {32'h450deb9e, 32'hc370bd5f, 32'hc2302d3b},
  {32'hc4f242ed, 32'h434fc677, 32'h4313ea5e},
  {32'h44728a86, 32'hc381f584, 32'hc07ccf00},
  {32'hc179a600, 32'hc3571ff0, 32'h410dd7cd},
  {32'hc2e8fdd3, 32'hc374e848, 32'hc29ff615},
  {32'hc4ac75f6, 32'h432bea5e, 32'h43561407},
  {32'h444461a2, 32'h414e3992, 32'hc28c4c08},
  {32'hc475eb78, 32'hc1713ff3, 32'hc314d086},
  {32'hc239bae0, 32'hbfa7ff50, 32'hc32eb233},
  {32'hc4c5b55b, 32'h42bbbb58, 32'hc32401bf},
  {32'hc2240550, 32'h4371a243, 32'hc3a49015},
  {32'hc489d97f, 32'hc286218b, 32'h439f864b},
  {32'h43efc7b0, 32'hc3947032, 32'hc3c431fb},
  {32'hc3dc97d0, 32'h43f68441, 32'h42dd01cd},
  {32'h452d81ee, 32'h4363936d, 32'hc30c8245},
  {32'hc3f20f3f, 32'h43cbcbf9, 32'h43412404},
  {32'h449e97e7, 32'h426c8dec, 32'hc2fdec63},
  {32'hc48d5fde, 32'hc1f32382, 32'h441a170a},
  {32'h44e6a12f, 32'hc187a11b, 32'hc1fc569f},
  {32'hc4bf93f2, 32'h43faa0d2, 32'h42687367},
  {32'h445ec778, 32'hc32c9b47, 32'hc39e7129},
  {32'hc4d05ab6, 32'h43a4fdaa, 32'hc2bfaa04},
  {32'h44064b73, 32'h439283e0, 32'h41bab812},
  {32'hc40fcd7d, 32'hc35b8a0e, 32'h4410f862},
  {32'h44f32fca, 32'h431ed86b, 32'hc1a1113b},
  {32'hc4cb7b2d, 32'h43f9320b, 32'h41782bae},
  {32'h4474b8c6, 32'h42a23ea6, 32'hc38b5a4f},
  {32'hc4bf4e9f, 32'hc2148902, 32'hc35c746a},
  {32'h43f0716c, 32'h41f19a6a, 32'hc35ed352},
  {32'hc4c37ab1, 32'h43191e52, 32'h439b54c7},
  {32'h44af195e, 32'hc332b916, 32'h4214f4b7},
  {32'hc4bedb24, 32'hc1cca3f3, 32'h42b1026b},
  {32'h44e59eab, 32'h4338469e, 32'hbfbda957},
  {32'hc4d24b42, 32'h40ca9547, 32'h4277ea97},
  {32'h437b9d43, 32'hc2b9bdf5, 32'hc1cc1de5},
  {32'hc464fb20, 32'hc30407c0, 32'h43e55b44},
  {32'h44ee51f7, 32'hc26f3fcf, 32'hc3d21cb4},
  {32'hc50362aa, 32'h420b5e55, 32'hc3862728},
  {32'h4499c663, 32'h43a3d7f3, 32'h43396b00},
  {32'h44d32e96, 32'h43bc83d4, 32'hc3d0fadb},
  {32'hc49d3968, 32'h43b31060, 32'hc2b7bd64},
  {32'h44de3ee7, 32'hc2e95838, 32'hc31d8464},
  {32'hc4669816, 32'hc396be63, 32'h4411d91b},
  {32'h43670280, 32'hc3307f39, 32'hc369830a},
  {32'h4276eec0, 32'h43bb197a, 32'hc38cedaf},
  {32'h41e6e080, 32'hc36348c5, 32'hc3cedd11},
  {32'hc48a6deb, 32'h43712661, 32'h42ccf7d5},
  {32'h446c7926, 32'hc1c57be3, 32'hc32b869d},
  {32'hc3d5d360, 32'hc29bbec3, 32'h432d87cf},
  {32'h44badd3c, 32'h42a3c6a8, 32'hc2cc7083},
  {32'hc4a47591, 32'hc236c7e4, 32'h4217a7b4},
  {32'h44ad5374, 32'hc3832e29, 32'hc253e858},
  {32'hc4e1c59c, 32'h4197aebc, 32'hc3360189},
  {32'h4314009e, 32'hc2d2644a, 32'h43350f60},
  {32'hc4c45e5c, 32'h43974842, 32'h416d308f},
  {32'h450b1e5e, 32'h42bf3f95, 32'h423eb100},
  {32'h3ec57000, 32'hc3f36c77, 32'h41fdcf70},
  {32'h450fb1b0, 32'h43894168, 32'h43bfd9a6},
  {32'hc50f4cf0, 32'hc200e05e, 32'hc38931d8},
  {32'h44dce22f, 32'h43fc8b81, 32'hc277f19c},
  {32'hc4d2db2e, 32'h42efe51d, 32'h43686db5},
  {32'h45127a38, 32'hc2518297, 32'hc3148919},
  {32'hc32f34c6, 32'hc343f068, 32'h40f95556},
  {32'h4503a59b, 32'hc2a23eda, 32'h41c6c920},
  {32'hc4917a4e, 32'h43025f6c, 32'h42ba8427},
  {32'h43b37c20, 32'h437475e6, 32'h43584302},
  {32'hc491cc2d, 32'hc3b5cfdc, 32'hc327beca},
  {32'h44c80e96, 32'hc2adf082, 32'h4336b939},
  {32'hc4c4e059, 32'hc36aae07, 32'hc3436a82},
  {32'h43f888d8, 32'h42e1d582, 32'hc0d9c4fa},
  {32'hc4a63203, 32'hc2af9488, 32'h42fbb79b},
  {32'h44975d68, 32'h4404cda2, 32'h43de38e1},
  {32'h438f87e4, 32'hc291fa96, 32'h43930329},
  {32'h4516d46c, 32'hbfde7a5c, 32'hc21ec9d3},
  {32'hc495e79b, 32'hc3e1b8b2, 32'h423d714a},
  {32'h44b9374c, 32'hc166e74c, 32'h42609825},
  {32'hc4ea848e, 32'h4378557a, 32'h43a57060},
  {32'h4436396d, 32'hc08f08dc, 32'h4390f635},
  {32'hc4b93bb2, 32'hc2c40e79, 32'hc33e21a8},
  {32'h44986e85, 32'hc210259b, 32'hc314e178},
  {32'hc468ab50, 32'hc2f9048c, 32'h43141767},
  {32'h4471823e, 32'h417b67da, 32'h43acbda0},
  {32'hc4cf9f53, 32'hbf97599c, 32'hc2e13132},
  {32'h44cc5165, 32'h4107734a, 32'hc376b545},
  {32'hc4efc530, 32'hc3d5aa98, 32'h42b992c2},
  {32'h4323fb24, 32'h42b97235, 32'h43ac7060},
  {32'hc49d26e4, 32'h430dda47, 32'hc3cc400e},
  {32'h442edffc, 32'h43d80197, 32'hc2e92140},
  {32'hc4d63c0b, 32'h427bdcd6, 32'hc2d5aa7f},
  {32'h43a15f5c, 32'h43268447, 32'h43349824},
  {32'hc507ccf2, 32'hc41ba4ce, 32'hc372e6e7},
  {32'h44ad6df2, 32'h4424d4e6, 32'hc3ad87a9},
  {32'hc4ba31d0, 32'hc157ac6d, 32'h43afdb85},
  {32'h44da7052, 32'hc3f24340, 32'hc2eaa33b},
  {32'hc43311a0, 32'hc359ab1b, 32'h42c8f555},
  {32'h43a7e304, 32'h43d6a9e3, 32'hc2d52feb},
  {32'hc4c5b0e2, 32'hc248e692, 32'hc0c4b312},
  {32'h433c1630, 32'hc2aa154c, 32'hc3f29a6d},
  {32'hc4c6111f, 32'hc389727d, 32'hc2f913fc},
  {32'h4482b7aa, 32'hc3d1c79e, 32'h40f99868},
  {32'hc4f1a5d7, 32'h436ec516, 32'hc2b769f7},
  {32'h44d4075d, 32'hc33f5aa8, 32'hc3624051},
  {32'hc4b34fb2, 32'hc302dc32, 32'h42919ca0},
  {32'h44dd7459, 32'hc3041d3c, 32'hc1bee7bc},
  {32'hc4d4af5e, 32'hc396219b, 32'hc3c67707},
  {32'h450d960c, 32'h43843ac6, 32'hc3f0b984},
  {32'hc2f4cfa0, 32'hc39de307, 32'hc3f8be94},
  {32'h44201903, 32'hc20322c9, 32'hc2984222},
  {32'hc3dec808, 32'h4362a6b4, 32'h43e001a2},
  {32'h44ae377c, 32'hc2dde631, 32'h426aafe0},
  {32'hc4793cc2, 32'h4057e0c8, 32'h4363afce},
  {32'h43960625, 32'hc3079ac9, 32'hc31bb6be},
  {32'hc335df86, 32'h3f81ad61, 32'h433d4e1c},
  {32'h445f41a7, 32'hc030c1ec, 32'h42ac5794},
  {32'hc3a22c78, 32'h43971059, 32'h435aab93},
  {32'h44f8e439, 32'h4293ec37, 32'hc3faac27},
  {32'hc3056887, 32'h437972a9, 32'h4236b5e2},
  {32'h432bf970, 32'h42baf364, 32'hc3597070},
  {32'hc4e8b22f, 32'h4382a9b9, 32'h42875b15},
  {32'h4453b9dc, 32'hc2646548, 32'h439f8e5b},
  {32'hc504466d, 32'hc25f7803, 32'hc3278daa},
  {32'h44bc9a12, 32'h42c49d91, 32'h43ccd9a4},
  {32'hc505cd64, 32'h42d392a4, 32'h43171e22},
  {32'h4485955e, 32'h438f2db2, 32'h424971ad},
  {32'hc49f26b6, 32'h433a4242, 32'h42a8479c},
  {32'h44760c94, 32'h43b05422, 32'hc3283259},
  {32'hc51b4df0, 32'hc32dd318, 32'hc3a2b1fb},
  {32'h4500d57f, 32'h4298855f, 32'hc2ba4022},
  {32'hc3702190, 32'hc215bdfd, 32'hc22f8632},
  {32'h4503bb0d, 32'hc1b91a9e, 32'hc297d2be},
  {32'hc509e4b9, 32'h4289b775, 32'hc37109a0},
  {32'h4445e826, 32'h43d4b8ec, 32'hc3df6cc1},
  {32'hc4f03196, 32'hc3210b08, 32'hc33311d8},
  {32'h44ef32a6, 32'h42e65bcf, 32'h437eae94},
  {32'hc465dd0c, 32'hc36409b5, 32'h42e16f5b},
  {32'h44e38fdd, 32'h436df4e4, 32'h427370a0},
  {32'hc4352ae8, 32'hc3a2ad73, 32'hc307334a},
  {32'h44b01395, 32'hc33126fc, 32'hc2f9ffbd},
  {32'hc4b73e1f, 32'hc231de16, 32'h4223fbea},
  {32'h44b5be9d, 32'hc3451c5b, 32'hc36b13e8},
  {32'hc42680f2, 32'h43245d76, 32'h42ee69b4},
  {32'h44e6e4a1, 32'h42b889b8, 32'h43a24937},
  {32'hc5050c4c, 32'h4204af32, 32'h433dba6a},
  {32'h44f7d522, 32'h4336aace, 32'h4332ccc6},
  {32'hc4065255, 32'h4233b903, 32'h41d9eea4},
  {32'h4506ded1, 32'hbf8fef2c, 32'h3f05aa88},
  {32'hc4bdccb0, 32'hc22b0342, 32'hc31d9ca9},
  {32'h4458a79b, 32'hc2df242e, 32'hc2181b53},
  {32'hc39964e5, 32'h41021ab9, 32'hc336c577},
  {32'h44fccd33, 32'h437e1296, 32'hc3205b4f},
  {32'hc49dff9c, 32'h43e45958, 32'h43466f5e},
  {32'h44d5efab, 32'h4321af30, 32'hc24e0a83},
  {32'hc414a1d5, 32'hc2909633, 32'h42a54573},
  {32'h44d6c158, 32'hc288a714, 32'hc19ace1c},
  {32'hc4736b30, 32'hc3318574, 32'h426bde4a},
  {32'h44c6bd4e, 32'hc39c9512, 32'hc3599acf},
  {32'hc4f65789, 32'h43162a7b, 32'h432b3faf},
  {32'h45261682, 32'hc3de2a63, 32'h41bc2291},
  {32'hc46562c0, 32'h42ad880a, 32'h437d354d},
  {32'h44dff1c2, 32'hc2c942c9, 32'h4272b1c1},
  {32'hc42abf0a, 32'h42af18a5, 32'hc32a5471},
  {32'h44c3215a, 32'hc3aaa865, 32'hc19505b0},
  {32'hc4a2581a, 32'hc21ab52a, 32'h4367431e},
  {32'h451c3c5c, 32'h4348a6a0, 32'hc2f217fa},
  {32'hc4f1f3b1, 32'hc3aecc96, 32'hc2e8608c},
  {32'h44c5e5ef, 32'h437afe3e, 32'h4300af57},
  {32'hc5008bf8, 32'hc309beb6, 32'hc312206c},
  {32'h4515e21d, 32'h4346e523, 32'h41c372e8},
  {32'hc2e0aff0, 32'h436dc643, 32'h433215d5},
  {32'h451601c4, 32'hc33383e7, 32'h43cba127},
  {32'hc3f288a4, 32'hc3695e1c, 32'hc2919389},
  {32'h4484628e, 32'h43dda160, 32'h432be1d0},
  {32'hc4a59dcb, 32'h43a1d448, 32'h43248bab},
  {32'h43e74d5a, 32'h41f9ae6c, 32'h416de088},
  {32'hc4e5d04c, 32'h4284b646, 32'hc320ba50},
  {32'h44922ff9, 32'h41ea07c2, 32'h43225c89},
  {32'hc4f372cb, 32'hc380554f, 32'h43a01bbe},
  {32'h44dc25c4, 32'hc3071bfb, 32'hc2f1a88d},
  {32'hc4c5a190, 32'h435fb2fc, 32'hc329128f},
  {32'h44b00b7f, 32'hc35596c9, 32'hc2b3d871},
  {32'hc48f805a, 32'h43597ce7, 32'hc2c119c4},
  {32'h43e526e0, 32'hc40318e6, 32'hc31fcc53},
  {32'hc36a6a10, 32'h432ee1ae, 32'hc2cb755c},
  {32'h449856dc, 32'hc108c03d, 32'h4359f909},
  {32'hc4998558, 32'h43d1c27c, 32'hc0027bf0},
  {32'h4504d95b, 32'h44610203, 32'hc166040b},
  {32'hc467cfdc, 32'h4168abfa, 32'h4276d154},
  {32'h44a7a7a3, 32'hc2ff523f, 32'h4387a612},
  {32'hc4f43dbf, 32'h438b9f1b, 32'h424379b7},
  {32'h43ba7eae, 32'h40d3718d, 32'h434410ed},
  {32'hc3f79d04, 32'h42ebbf98, 32'h41c63f4f},
  {32'h437b0ab8, 32'hc265f84f, 32'hc33897ff},
  {32'hc3918254, 32'hc34eed15, 32'h434f872f},
  {32'h44c39a1a, 32'hc302de8e, 32'hc3aa196f},
  {32'h4374fb9c, 32'hc246798d, 32'hc2492043},
  {32'h450d83a3, 32'h420f43b6, 32'hc3b27366},
  {32'hc510fc6c, 32'h4323a21f, 32'h3f90e430},
  {32'h4425c1b6, 32'h43b52b01, 32'hc34d4b62},
  {32'hc3963c8d, 32'hc25a3f85, 32'h43b09a17},
  {32'h44e5b612, 32'h43590733, 32'hc1b645b5},
  {32'hc3ce5029, 32'hc3c20b9c, 32'hc37e4650},
  {32'h449ce590, 32'hc0c1fb00, 32'hc2d007dc},
  {32'hc4e7d504, 32'h43b9943b, 32'h42c82927},
  {32'h44be462c, 32'hc1702d92, 32'hc2b4eb75},
  {32'hc4b1ff0e, 32'h432ed3b5, 32'h42208264},
  {32'h4413e9fd, 32'hc257d875, 32'h42fb96e1},
  {32'hc4588667, 32'hc385b6dd, 32'h43820aea},
  {32'h44bcab90, 32'h404a123c, 32'hc322caca},
  {32'hc4a5b23b, 32'hc2d6439e, 32'hc38b4a1c},
  {32'h44ce733c, 32'hc2179759, 32'h4338a2b5},
  {32'hc4ba682a, 32'hc2ffbe5e, 32'h431771e8},
  {32'h4416f2e1, 32'hc3a34b78, 32'hc3b11340},
  {32'hc509a1ce, 32'hc2c4af04, 32'h4204024a},
  {32'h4464f143, 32'hc380e894, 32'h4307a49c},
  {32'hc524554f, 32'hc2bc4e87, 32'hc26a3e37},
  {32'h44b41546, 32'hc2f36d7d, 32'hc359d81d},
  {32'hc4f84543, 32'h422a6c00, 32'h429d3068},
  {32'h44b3e0b9, 32'h43a92ad3, 32'hc3754908},
  {32'hc4420966, 32'hc3aa1d1c, 32'hc407f4bb},
  {32'h44bb30fb, 32'hc3bbaae1, 32'h4289e5b7},
  {32'hc2d75100, 32'hc311c1de, 32'hc307c805},
  {32'h42c92da0, 32'hc3562db8, 32'h4236a79b},
  {32'hc4995a63, 32'h41e008c2, 32'h4268b38e},
  {32'h4453ffac, 32'hc3a1e949, 32'h43847ade},
  {32'hc4de5842, 32'h43843cea, 32'hc20861b0},
  {32'h4519dc90, 32'h43e5b879, 32'hc3964c63},
  {32'hc3cfcbba, 32'h43ef764f, 32'hc3700783},
  {32'hc4019b97, 32'h40a6c894, 32'hc20fe52c},
  {32'hc50353f6, 32'h428d931d, 32'hc36c04a2},
  {32'h446ca053, 32'hc2b1093c, 32'hc30acbaf},
  {32'hc4e06101, 32'h3dc14e00, 32'h43802e54},
  {32'h450dece3, 32'hc2897665, 32'h43067858},
  {32'hc32180d7, 32'hc274f198, 32'h43972017},
  {32'h4510ccd5, 32'h4304c392, 32'h438b3200},
  {32'hc4ebe787, 32'h4393570c, 32'hc3484e72},
  {32'h44922e43, 32'hc2606696, 32'hc2c736ff},
  {32'hc4e5038e, 32'hc397091d, 32'hc29e398e},
  {32'h440b478b, 32'h4243d3d8, 32'h4324d4e3},
  {32'hc503f9cb, 32'h43c512dd, 32'h4318772f},
  {32'h4466a28c, 32'h434cf620, 32'h430b4c8e},
  {32'hc33969ee, 32'hc1dc6813, 32'h43310a71},
  {32'h45054780, 32'h429b492b, 32'h4281d4bf},
  {32'hc45794b6, 32'h432665dc, 32'h40310050},
  {32'h440828d9, 32'h3fb7eead, 32'h4373941f},
  {32'h4323e018, 32'h4309efc0, 32'h41a8c3e4},
  {32'h449e980c, 32'hc38df0f1, 32'hc2d8b7a9},
  {32'hc4288169, 32'h43a40ae3, 32'hc41a4b24},
  {32'h4480a360, 32'hc3bf4198, 32'hc190ec76},
  {32'hc47b26c0, 32'h43080934, 32'hc3e7bb8c},
  {32'h445a88b8, 32'hc330323b, 32'hc304a6c9},
  {32'hc3118239, 32'hc3b5ac5c, 32'h428d3b9a},
  {32'h44ad0630, 32'h4306aad1, 32'hc3728c7c},
  {32'hc490c08a, 32'h4431998d, 32'h43b667b2},
  {32'h44abf856, 32'h4336de08, 32'hc296dadd},
  {32'hc3236f2a, 32'h423c47cf, 32'hc1ff0134},
  {32'h44fd81ad, 32'hc3316bcc, 32'hc383e81a},
  {32'hc4f65b7e, 32'hc2a8a607, 32'hc3bd6fbc},
  {32'h437c61c0, 32'hc391f685, 32'hc134276e},
  {32'hc48311c8, 32'hc2a246b1, 32'h4327416b},
  {32'h44b6808e, 32'hc379d990, 32'hc2302625},
  {32'hc4f7611b, 32'h43602bc8, 32'hc3735a6c},
  {32'h44b6094f, 32'hc11032d3, 32'h4308615a},
  {32'hc498723f, 32'hc3c99b08, 32'h438afed7},
  {32'h44ee8566, 32'h423c8c9a, 32'h4286f795},
  {32'hc50c439f, 32'h434e37ac, 32'hc3633641},
  {32'h44b16618, 32'h43846c8a, 32'hc3302214},
  {32'hc4943ff8, 32'hc3be7bb5, 32'hc295484e},
  {32'h4350d6e0, 32'h425b36dd, 32'h3f877bd0},
  {32'hc50bf53a, 32'hc33a0496, 32'h436d4f68},
  {32'h44dfb2da, 32'h429406fb, 32'hc3798784},
  {32'hc47dc872, 32'h430494dd, 32'h42978434},
  {32'h43a7df62, 32'hc2b5cfcd, 32'hc359d1cc},
  {32'hc5045b1c, 32'hc34a53de, 32'h41536b65},
  {32'h4492647d, 32'h43ac5550, 32'hc380b768},
  {32'hc465fd2b, 32'hc261c22f, 32'hc3256553},
  {32'h44dfaf52, 32'h43542cec, 32'h42764f38},
  {32'hc492c268, 32'h42ef7880, 32'hc34f002e},
  {32'h44031560, 32'hc28d63a0, 32'h42d71b53},
  {32'hc4e124b2, 32'hc19fc01d, 32'h41b10fea},
  {32'h44f56766, 32'hc30d022b, 32'hc38760e7},
  {32'hc4a0b512, 32'hc22a9f34, 32'h4238be1d},
  {32'h44b23a1a, 32'hc337be32, 32'hc2ebc0a5},
  {32'hc476d5f5, 32'hc2cc790c, 32'hc20e3418},
  {32'h4400cf10, 32'h433929be, 32'h421468e4},
  {32'hc4430147, 32'h42915804, 32'h42b325e0},
  {32'h44926972, 32'hc2c3c0a0, 32'h4213a087},
  {32'hc505c8d1, 32'h43653ba3, 32'hc2129826},
  {32'h45141998, 32'h440ad590, 32'hc34edb47},
  {32'hc3a5da30, 32'hc3c2aea7, 32'h43825af0},
  {32'h44c108ba, 32'h42ebf114, 32'hc38a48b2},
  {32'hc4669e5e, 32'hc35872e6, 32'h426a4ac1},
  {32'h443f73ff, 32'h418f4178, 32'h42ec396d},
  {32'hc4fa989c, 32'hc2d0b011, 32'h42dd2fe4},
  {32'h436532c8, 32'h42e48c14, 32'hc364e1f2},
  {32'hc4badc94, 32'hc3941017, 32'h434b0fef},
  {32'h440f2441, 32'hc20ebdeb, 32'h42bf1343},
  {32'hc4992aea, 32'h42a881f9, 32'h42b1a53f},
  {32'h44db777d, 32'h43c88f26, 32'hc29568c0},
  {32'hc4ab6b30, 32'hc347fac5, 32'h43241089},
  {32'h43607fc0, 32'h42ead9d4, 32'hc41c0714},
  {32'hc4d88be4, 32'h4323733f, 32'hc25d0f47},
  {32'h442e53da, 32'hc2a4b176, 32'hc39e4c9c},
  {32'hc4d43ad6, 32'h4243528a, 32'h42a57df4},
  {32'h44eaa9af, 32'h434b9555, 32'hc3d3d841},
  {32'hc41dfb0e, 32'hc24443ac, 32'h43de8a24},
  {32'h44d16a47, 32'hc399f410, 32'hc3b51cd9},
  {32'hc3b732d8, 32'h42e9af9a, 32'h435b5ae2},
  {32'h44e94b0f, 32'hc37432f8, 32'h41b2cf53},
  {32'hc4bc1acf, 32'hc306b8a7, 32'hc341293e},
  {32'h4424dd86, 32'h42aa737f, 32'hc36f1f31},
  {32'hc48e1683, 32'h43b50b5e, 32'h44365ca0},
  {32'h44d25282, 32'h4308ef0d, 32'hc2e34dfb},
  {32'hc4d792d0, 32'h41297f96, 32'hc311a669},
  {32'h422988a4, 32'hc3840289, 32'h43147c0e},
  {32'hc3e3e180, 32'hc3c16b5b, 32'h4337ebee},
  {32'h442e0bf9, 32'hc30b5321, 32'hc380fcd4},
  {32'hc4a4dbda, 32'hc18a9e6a, 32'h435ef5d9},
  {32'h450a5d68, 32'hc327d5fb, 32'h430f5f69},
  {32'hc519f6f9, 32'h431b5342, 32'hc36b0c5f},
  {32'h441513b5, 32'h43db33d2, 32'h42a0a150},
  {32'hc4b0ac58, 32'hc364b365, 32'hc406140f},
  {32'h44f7ba79, 32'hc360b29b, 32'h43a76c5c},
  {32'hc512349f, 32'hc1d7f71a, 32'hc1c404d0},
  {32'h44534a00, 32'hc3b1f8ff, 32'hc239a76a},
  {32'hc28708f2, 32'h43582e74, 32'hc309929b},
  {32'h4456258a, 32'hc2d040ec, 32'h439987ce},
  {32'hc4406493, 32'hc31d468f, 32'hc211fb98},
  {32'h429af384, 32'hc3ae77c1, 32'h418f0ea4},
  {32'hc44cfe6a, 32'h4381e002, 32'hc2ecb67d},
  {32'h43689504, 32'hc335c92c, 32'h42decea3},
  {32'hc4eb3761, 32'h42c61b4d, 32'h4386b0e0},
  {32'h4437ae93, 32'h4285d641, 32'hc3a17b58},
  {32'hc494a2d8, 32'h43de384f, 32'hc1fbac36},
  {32'h4204c3c0, 32'hc370e9dc, 32'hc28f7b98},
  {32'hc4c4983c, 32'hc3901577, 32'h41de167d},
  {32'h44bec192, 32'h428824a8, 32'h43521199},
  {32'hc46fdf5e, 32'h433649aa, 32'h436b5345},
  {32'h451ba5b7, 32'h40d2e214, 32'h43828435},
  {32'hc3ceddae, 32'hc3ab0f9e, 32'h43c9fb81},
  {32'h449aa8f9, 32'h417a740b, 32'hc348200b},
  {32'hc4e3a8aa, 32'h4307819a, 32'hc380d407},
  {32'h4508a019, 32'hc2e5f3ee, 32'hc064fc72},
  {32'hc47b193c, 32'h434cf0d2, 32'hc32b4b2d},
  {32'h44a3e1bd, 32'h42ab4025, 32'hc33cd5f3},
  {32'hc4bc7c49, 32'hc3ed8893, 32'h42a6d250},
  {32'h449e0810, 32'h434dad44, 32'hc40f47a6},
  {32'hc502a032, 32'h4155abad, 32'hc2860d60},
  {32'h4482939e, 32'h43937692, 32'hc34bc1c4},
  {32'hc4eb54cd, 32'h4277d088, 32'h4256e9aa},
  {32'h4528c3fa, 32'hc3c304d3, 32'hc222be61},
  {32'hc513ecc7, 32'hc3193471, 32'hc2e5df9e},
  {32'h43fc1eae, 32'h42187790, 32'hc29922a8},
  {32'hc4f47acd, 32'hc1fe2930, 32'h3f24b134},
  {32'h450a7ab6, 32'h4292431e, 32'hc2c9aae9},
  {32'hc3f4dd60, 32'h41c1ce34, 32'h440493b7},
  {32'h4519f96b, 32'hc260dae5, 32'hc19e06c2},
  {32'hc31187f0, 32'hc3c9534a, 32'h43a846d9},
  {32'h4485fe88, 32'hc3610909, 32'hc40f2e70},
  {32'hc4456e27, 32'h435ef043, 32'hc29e0a0d},
  {32'h450040c3, 32'hc2ffacc7, 32'hc3ce7070},
  {32'hc4a73146, 32'h43acb54a, 32'hc3686270},
  {32'h4445f45a, 32'hc29e6e5c, 32'h4314ef04},
  {32'hc4899854, 32'hc3410509, 32'hc2d57549},
  {32'h442837be, 32'hc323e594, 32'hc23f57af},
  {32'hc4ba7452, 32'h429b3183, 32'hc25b0651},
  {32'h44b5ace4, 32'hc19309d6, 32'h4311ed75},
  {32'hc5017f3a, 32'h43bb889e, 32'h43b14110},
  {32'h44ba43ac, 32'hc2bc6b88, 32'h435b1011},
  {32'hc3504870, 32'hc1138fac, 32'hc32539b9},
  {32'h44a89dc0, 32'hc16fd168, 32'h42df6c6d},
  {32'hc51a542a, 32'h43669327, 32'h43433f1b},
  {32'h449ee5c4, 32'hc3a3761c, 32'hc3035346},
  {32'hc3ec53e3, 32'hc26a57d2, 32'hc36e779b},
  {32'h45015dd2, 32'h429ac2b4, 32'h429fc350},
  {32'hc45c6abe, 32'h439769a2, 32'hc3acef72},
  {32'h44cbba46, 32'hc0bed4a4, 32'hc2d04d77},
  {32'hc44c0d7f, 32'hc20e1f1f, 32'h4313e0f8},
  {32'h4493bf83, 32'h4307344a, 32'hc212b22c},
  {32'hc4ed34ad, 32'hc189058e, 32'hc4038229},
  {32'h44e7a9a2, 32'h4243609e, 32'h42a2e0ed},
  {32'hc3b2ebbc, 32'h42dd40de, 32'h4293973d},
  {32'h441cc1de, 32'h431f3485, 32'h42f3e96c},
  {32'hc4dd5eab, 32'hc3f19670, 32'hc05e9ad0},
  {32'h44dd31de, 32'h436a396f, 32'hc3afd7d3},
  {32'hc4cd4927, 32'h42cbcd11, 32'h415de700},
  {32'h42d54d6c, 32'h42d01805, 32'hc296b569},
  {32'hc3d5eeba, 32'h4402d71b, 32'hc394e384},
  {32'h45105f51, 32'h41fb7937, 32'hc36ae97a},
  {32'hc4ea3cf2, 32'hc2417b0d, 32'h432fa681},
  {32'h445103ea, 32'h4324eea9, 32'h433a00e2},
  {32'hc4cdf691, 32'hc34d9e70, 32'hc0917628},
  {32'h45186746, 32'hc2a6c803, 32'hc3ae047e},
  {32'hc402810d, 32'hbfb6a649, 32'hc30f5a87},
  {32'h4486b7ff, 32'hc3e7abc4, 32'hc36e8e35},
  {32'hc48d5c56, 32'hc1771ffd, 32'hc2574e5c},
  {32'h44bb9569, 32'h4270bfbf, 32'hc0f60e3c},
  {32'hc4d65ab6, 32'hc305917b, 32'h42893f83},
  {32'h4366ccc8, 32'h43fa5fb8, 32'h42600e16},
  {32'hc451ccd3, 32'hc2ba369b, 32'hc31cdded},
  {32'h44a1dad1, 32'h437cbaba, 32'h43b7f570},
  {32'hc4de5408, 32'h4313992d, 32'hc2473e8e},
  {32'h441e6eb8, 32'hc3b4f31a, 32'h42f3f04a},
  {32'hc4b50f50, 32'h41aa7590, 32'hc2388079},
  {32'h443d6324, 32'hc3e2be77, 32'hc1f07119},
  {32'hc50a6aaf, 32'h43a28d8e, 32'hc38305cb},
  {32'h43fa1728, 32'hc2dc78f9, 32'hc2c30086},
  {32'hc5034734, 32'h438edb3f, 32'h43ae0958},
  {32'h437bcfe0, 32'h434e3795, 32'h42de31b0},
  {32'hc3142f1c, 32'h439691bd, 32'h42407977},
  {32'h435583d0, 32'h4356e0a7, 32'hc3ad1ce0},
  {32'hc47094e0, 32'hc3a22fa9, 32'h42b36d1e},
  {32'h451dc248, 32'hc321aa92, 32'hc2aaf31d},
  {32'hc3b5d71c, 32'hc2be9529, 32'hc3d68999},
  {32'h44cde537, 32'h42ff0dac, 32'h43942961},
  {32'hc46c8312, 32'h430bafef, 32'h416f557f},
  {32'h43c809f8, 32'h40f4f603, 32'hc18c5190},
  {32'hc514358c, 32'h437b98f0, 32'hc26727d9},
  {32'h43a199a8, 32'h43872eb7, 32'h4392bf7c},
  {32'hc42def01, 32'h439c26f8, 32'hc1c22f46},
  {32'h43f485df, 32'h43b25b62, 32'hc28663dc},
  {32'hc3b5bb6d, 32'h437c372d, 32'hc1983adf},
  {32'h4291b920, 32'h42fe2291, 32'h42a6bf92},
  {32'hc41993d6, 32'h43836247, 32'hc31428be},
  {32'h4522f1d4, 32'hc37b0355, 32'h440bee91},
  {32'hc4d813d6, 32'hc3861716, 32'h42b3932f},
  {32'h441cc42d, 32'hc38c4767, 32'h43636bce},
  {32'hc4e2fc00, 32'h41eb09a6, 32'h4338b103},
  {32'h44ffd6d5, 32'h41f6eb10, 32'h43788e77},
  {32'hc4e6ae78, 32'hc3d526d6, 32'hc3600cd9},
  {32'h44f3030a, 32'hc38ad24b, 32'h428af2d7},
  {32'hc2e274fe, 32'h433a0939, 32'h42a39135},
  {32'h44b8c24a, 32'hc31745d5, 32'hc20b2340},
  {32'hc4c16876, 32'hc3a6f519, 32'hc34010bf},
  {32'h45036b74, 32'h41e3eaf6, 32'hc36d22be},
  {32'hc4e16ffd, 32'hc283137a, 32'hc3a247b6},
  {32'h433500c8, 32'hc2bf1ae3, 32'h4373855f},
  {32'hc420dcf4, 32'h42db2932, 32'hc2fe8681},
  {32'h450916a8, 32'h42ced371, 32'hc39695f6},
  {32'hc38d20de, 32'h414f477c, 32'hc33ec187},
  {32'h44849383, 32'h430e99ce, 32'h439947cb},
  {32'hc4ccf4fa, 32'h42c98075, 32'hc3ebfe3e},
  {32'h43241980, 32'hc32a3a2e, 32'h42b7a94d},
  {32'hc350a930, 32'h4349513a, 32'h420e99ce},
  {32'h4501d251, 32'hc22cd5a8, 32'h435ea2e2},
  {32'hc43bfa40, 32'h43c4718a, 32'h42dc5d54},
  {32'h44fd7e99, 32'h438f4cf1, 32'h4307e276},
  {32'hc4ccf229, 32'hc33747e5, 32'hc3ad19ae},
  {32'h44929ea0, 32'h435ca2ed, 32'h43a0c0bb},
  {32'hc4f76662, 32'h430e2e34, 32'h420e2c56},
  {32'h430669e0, 32'h4246957a, 32'h40a636fc},
  {32'hc4a3e52a, 32'hc30335d7, 32'hc32329b7},
  {32'h450c6c3a, 32'h437f74e3, 32'hc4196a58},
  {32'hc4fd027c, 32'hc2fee8c4, 32'h42cd6ded},
  {32'h44c77e1e, 32'h42814196, 32'h439ae3af},
  {32'hc4b86402, 32'h42bf3f6f, 32'h4398325b},
  {32'h44d36329, 32'hc10f9e44, 32'h442620a7},
  {32'hc326fea2, 32'hc1e4fabd, 32'hc3660fba},
  {32'h44e86434, 32'h407f8ac7, 32'hc31c0398},
  {32'h433c5670, 32'h43f16344, 32'hc2d2da5e},
  {32'h4403b0b4, 32'hc359e399, 32'h42cd31bd},
  {32'hc4b2c5fb, 32'h43e042c7, 32'h434471a5},
  {32'h43204990, 32'hc38d7f58, 32'hc23636ec},
  {32'hc42e0b0c, 32'h4406f3c9, 32'hc39686a0},
  {32'h44363a80, 32'h421c6489, 32'h43a66e9d},
  {32'hc4cd4e30, 32'h436a55c1, 32'hc2c7228a},
  {32'h44b9c89e, 32'hc2c8cee8, 32'hc18360d9},
  {32'hc4f1b84f, 32'hc13e6e8f, 32'hc1722e0a},
  {32'h44d155a5, 32'hc382b472, 32'h4326f317},
  {32'hc51c717e, 32'h43141f8f, 32'hc32cff13},
  {32'h44f06f53, 32'hc3632d6b, 32'h432721bd},
  {32'hc472d4d5, 32'hc3ed4703, 32'hc3fdeab7},
  {32'hc4c7d696, 32'hc32f0ff8, 32'h436b5f22},
  {32'h4508a256, 32'h437eba1b, 32'h43973949},
  {32'hc347b2c5, 32'h4391cec1, 32'hc2cf3e31},
  {32'h43bcd1a4, 32'hc2cf349b, 32'h430184fb},
  {32'hc4c161a8, 32'hc3bf3616, 32'hc282b23c},
  {32'h44fabdc7, 32'hc41453ab, 32'h41a74241},
  {32'hc4b62b80, 32'h42b17fbc, 32'hc3c11208},
  {32'h443d2801, 32'h43413320, 32'h420cf423},
  {32'hc4fa73dd, 32'h40f6a80b, 32'hc11e006a},
  {32'h4457fbcc, 32'hc3113b9e, 32'h42a4618c},
  {32'hc4965694, 32'h425c3048, 32'hc3af8474},
  {32'h443a2eec, 32'h429bf344, 32'hc2b35c8a},
  {32'hc41b9f14, 32'h4367ed6d, 32'hc3827d30},
  {32'h4495c005, 32'h43e2d7a3, 32'h43b71482},
  {32'hc4fd3fa6, 32'hc356c16f, 32'h42e84e08},
  {32'h4506656d, 32'h433dc326, 32'h4268b256},
  {32'hc4fecd28, 32'hc31407c0, 32'hc3327d92},
  {32'h440028a9, 32'hc13e59e3, 32'hc18d7d0e},
  {32'hc39ae3c8, 32'h434ea338, 32'hc3404ec6},
  {32'h44987e21, 32'h43870236, 32'h429bd48f},
  {32'hc50a458e, 32'h4377b496, 32'hc34516e2},
  {32'h44f41738, 32'hc251bd66, 32'hc2a18b5e},
  {32'hc398ea74, 32'h43429bdc, 32'hc3a5b8fa},
  {32'h44a8ce56, 32'h4314954e, 32'h43186f8d},
  {32'hc41b8d40, 32'h423a950c, 32'hc364863f},
  {32'h445491e0, 32'h43b8b2f7, 32'h435f97ce},
  {32'hc513f7a4, 32'hc3137546, 32'h437ce404},
  {32'h429f105f, 32'hc31745c2, 32'hc399d1f0},
  {32'hc4b33dfa, 32'hc319b920, 32'hc3b4b70d},
  {32'h44641624, 32'h438d1a03, 32'h4261477b},
  {32'hc49499ce, 32'h42e9e586, 32'h43205415},
  {32'h428e5c70, 32'hc0e0ebad, 32'h43e43d34},
  {32'hc46c244a, 32'h4258a240, 32'hc34b5ca2},
  {32'h4475ae6c, 32'hc3318448, 32'h438a1a72},
  {32'hc3fdaff1, 32'h434b841a, 32'hc322eec9},
  {32'h42a5aba8, 32'hc35522b9, 32'hc2c745fe},
  {32'hc4fc7e54, 32'hc1aaabed, 32'h42c95638},
  {32'hc0874900, 32'hc30d0115, 32'hc2aef7b8},
  {32'hc4d00ce7, 32'hc1de2aac, 32'h416fa3f1},
  {32'h4405d06b, 32'hc3079085, 32'h41dee455},
  {32'hc4ab1a64, 32'hc31014a9, 32'h4273f422},
  {32'h448bcd59, 32'h434c5e52, 32'hc3080c1f},
  {32'hc4c52209, 32'hc230fce4, 32'h419f21a2},
  {32'h44a8f90d, 32'h429d4b69, 32'h440e2688},
  {32'hc46842a8, 32'h42e63c7d, 32'h420b0765},
  {32'h4510b174, 32'h435b7d83, 32'h43c6d928},
  {32'hc3a266b0, 32'h42e85525, 32'hc335f94c},
  {32'h44360080, 32'hc35badf8, 32'h437e275a},
  {32'hc4228232, 32'hc386af76, 32'hc2b6096a},
  {32'h43eba594, 32'hc373b837, 32'h42ef8eeb},
  {32'hc41e04b6, 32'hc3b91128, 32'hc3612100},
  {32'h43b21a18, 32'h4318425f, 32'h42873fa9},
  {32'hc4daafd6, 32'h42f6982c, 32'hc3d89cdf},
  {32'h44a295e0, 32'hc2fd0f7d, 32'h42ab4694},
  {32'hc4eb22c4, 32'h43402910, 32'h4366c12e},
  {32'h43ffd579, 32'h41fbdcc8, 32'h42caca74},
  {32'hc486b75a, 32'h42dbcc18, 32'hc3147961},
  {32'h44cf3b10, 32'h429297b1, 32'hc342298d},
  {32'hc4506149, 32'h42a0b0b0, 32'h431e8bf9},
  {32'h44ebe584, 32'hc28a778a, 32'h43b12f21},
  {32'hc35b487c, 32'h433e35e0, 32'hc2f0588f},
  {32'h45249269, 32'hc3f30cdf, 32'h43b4974f},
  {32'hc46a2456, 32'hc2e63012, 32'hc3a5e04f},
  {32'h44e718f2, 32'hc39b6f13, 32'hc3b72887},
  {32'hc420d4c8, 32'hc3acd9d2, 32'hc29c6725},
  {32'h452317f1, 32'h436c87aa, 32'h437250af},
  {32'hc4387f90, 32'h42ded34c, 32'hc1ad2e8d},
  {32'h441d7239, 32'h40f236bd, 32'hc33df7d9},
  {32'hc3ed23d8, 32'h437e23b1, 32'hc1cf9e6e},
  {32'h44f9951e, 32'hc38d6290, 32'hc3a7f34c},
  {32'hc4aa8de8, 32'h42846793, 32'h41f22641},
  {32'h44bf83cb, 32'hc3cc021e, 32'h43e74050},
  {32'h4412b274, 32'h44326153, 32'h430d177e},
  {32'h44b4206c, 32'h42d1158e, 32'h430f05e3},
  {32'hc50d69ef, 32'hc213610c, 32'h43731912},
  {32'h4460ba18, 32'h42db1814, 32'hc353b8bf},
  {32'hc5175da9, 32'hc2ddff9c, 32'h41e84aa3},
  {32'h447948de, 32'hc2ae4de0, 32'hc4057c88},
  {32'hc50f5fda, 32'h42fa2a36, 32'hc193de9a},
  {32'h450051a0, 32'hc388ba2a, 32'h4416e591},
  {32'hc3d1835a, 32'hc32c3982, 32'hc31a70c4},
  {32'h450a76b4, 32'hc3be1913, 32'hc2a64ab4},
  {32'hc4d2919b, 32'h437317c1, 32'hc3916b73},
  {32'h44f74732, 32'h43c9a4e0, 32'h42542724},
  {32'hc4fc5110, 32'h437c8b08, 32'h43b41247},
  {32'h446084eb, 32'h42a9b852, 32'hc2d2f6cd},
  {32'hc4c12baa, 32'hc2062125, 32'h43778320},
  {32'h44ae810e, 32'hc37624a8, 32'hc3682c4b},
  {32'h43dde3fb, 32'hc271621c, 32'h43dd76f1},
  {32'h448e5df0, 32'hc386d3dc, 32'h42ff03f6},
  {32'hc5120c95, 32'h42c0bcee, 32'h4242a7f4},
  {32'hc2656ea0, 32'hc3633a24, 32'hc35cf747},
  {32'hc4b3f666, 32'h439b7768, 32'hc27263d5},
  {32'h44297da9, 32'hc2df3da8, 32'h421472f9},
  {32'hc4c56abc, 32'hc3d0ed20, 32'hc3a81954},
  {32'h44f35b0d, 32'hc1f538f0, 32'hc379af08},
  {32'hc4261388, 32'hc39af26e, 32'h43166416},
  {32'h4507ffa9, 32'h41f0dc97, 32'hc2240251},
  {32'hc477dd04, 32'h438d9047, 32'hc391003d},
  {32'h43dbf4d0, 32'hc34e1788, 32'hc269b0ae},
  {32'hc4286a6e, 32'h436ba6f6, 32'hc2b41daf},
  {32'hc2eeea02, 32'h413248c2, 32'hc385523e},
  {32'hc4f208f4, 32'hc22d0e46, 32'hc2ddb2bd},
  {32'h44cd6fa4, 32'hc335fbfb, 32'h43c837fb},
  {32'hc50ae636, 32'h41b252a3, 32'h4312e6a3},
  {32'h44cd59ea, 32'hc2064888, 32'hc36e49c4},
  {32'hc1db8580, 32'h4338c717, 32'h3f601f10},
  {32'h44f65699, 32'hc2c40966, 32'hc3b4a803},
  {32'hc3c19e88, 32'hc23c2b8b, 32'hc316f8a1},
  {32'h44b44e81, 32'h442c39d8, 32'hc380b552},
  {32'hc512ab67, 32'hc28dd093, 32'hc32108ce},
  {32'h44cb532c, 32'h4363b370, 32'hc38605b0},
  {32'hc4db74f8, 32'h41fc5ab7, 32'hc2abc129},
  {32'h435ab8a0, 32'h4125aac8, 32'h43ed1eef},
  {32'hc3cf8185, 32'hc3da7d28, 32'hc2427a55},
  {32'h44eee4dd, 32'h43a5cb51, 32'hc3a99fa5},
  {32'hc4747098, 32'hc2cadb1a, 32'h419566e9},
  {32'h44e81728, 32'h43d5b0e3, 32'h43e6126e},
  {32'hc4941adc, 32'hc2f1b789, 32'h4331b689},
  {32'h4505637c, 32'hc252bc08, 32'h430f63a4},
  {32'hc48ee155, 32'h427c9457, 32'h43478ace},
  {32'h450560f0, 32'hc282e175, 32'h42174380},
  {32'hc4dfa220, 32'h42add88b, 32'h431e00db},
  {32'h44290fde, 32'hc29a7258, 32'hc1827073},
  {32'hc4ad5c99, 32'hc2b65818, 32'hc0e9a3b5},
  {32'h44fd18be, 32'hc1853c3f, 32'hc2a63404},
  {32'hc4013726, 32'h4358e419, 32'h4227fbc4},
  {32'h44fc4a30, 32'hc1544ba4, 32'hc2d281b3},
  {32'hc4b798cc, 32'hc1c97f38, 32'h4346a09c},
  {32'hc34b9da0, 32'hc3f40dff, 32'hc339e02e},
  {32'hc493abf8, 32'hc2a0f072, 32'hc320464c},
  {32'h41b2ce80, 32'hc33b8122, 32'h41a0be72},
  {32'hc41672c5, 32'hc2dc1436, 32'h4338dc12},
  {32'h44e7ca96, 32'hc3473c69, 32'hc2e2b87a},
  {32'hc4b6bede, 32'h43351677, 32'h4293bb94},
  {32'h4504b10d, 32'hc2e693f7, 32'hc3ac9492},
  {32'hc4533141, 32'h4303fe98, 32'hc3ac2919},
  {32'h418b2c00, 32'h4242db4d, 32'hc3ce0da9},
  {32'hc4142ec0, 32'hc2a08ae9, 32'h435af468},
  {32'h44367c38, 32'h43989885, 32'h41cbf3df},
  {32'hc4e4c40e, 32'h43cc34bf, 32'h433df486},
  {32'h44b71e3b, 32'hc3287bc4, 32'hc202eeb1},
  {32'hc4188d96, 32'h43ae6b34, 32'h41a72d0b},
  {32'h44b44478, 32'hc3892241, 32'h43904820},
  {32'hc5000bf4, 32'h435c6f63, 32'h43124c44},
  {32'h44f3077a, 32'hc32451ec, 32'hc39073b6},
  {32'hc477cc3c, 32'h42addf8b, 32'h429e0c05},
  {32'h451450eb, 32'h430fc6ee, 32'hc275b58e},
  {32'hc485b839, 32'h43d47bd6, 32'h4317263f},
  {32'h44214bb4, 32'hc287ee58, 32'hc335c43a},
  {32'hc4f25a87, 32'h42ce911b, 32'h428d44e4},
  {32'h43fe76ac, 32'h43ddb539, 32'hc26ca9ad},
  {32'hc4fcc2b0, 32'h4361d351, 32'h42db2c56},
  {32'h43bf1e18, 32'hc376cefc, 32'hc389d69b},
  {32'hc481b590, 32'h42507bfc, 32'h421efa99},
  {32'h4515ddc2, 32'h43aa064e, 32'h43a226e4},
  {32'hc3675af8, 32'h42bf34f0, 32'hc0d2ae9b},
  {32'h4506e234, 32'h41f2bbf2, 32'h4360e730},
  {32'hc4df10ba, 32'hc2c261c2, 32'h43a0b1a1},
  {32'h44d118a8, 32'h421085a0, 32'h40bbee88},
  {32'hc4f96ef6, 32'h3e29fd80, 32'hc23ea6fa},
  {32'h44c54d2e, 32'h424e001a, 32'hc3ab1e81},
  {32'hc4d1cabc, 32'h437d9dd4, 32'hc31bbdfd},
  {32'h44b523c7, 32'h43083072, 32'h43809c02},
  {32'hc44f2257, 32'h4175557e, 32'h43353c21},
  {32'h446d98d7, 32'h41bd6d27, 32'hc31cb125},
  {32'hc359f03f, 32'hc307ae36, 32'h435511ed},
  {32'h44798728, 32'hc3cb6902, 32'h43886896},
  {32'hc45090b0, 32'hc3c6e823, 32'h43547cdd},
  {32'h443a35ab, 32'hc39839dc, 32'h43a1a95d},
  {32'hc46931a8, 32'h43ab6805, 32'hc19eddb2},
  {32'h44ffb6b0, 32'h4321cfa5, 32'hc389b286},
  {32'hc5119161, 32'h41b65722, 32'h42b764a5},
  {32'h44fd6d10, 32'h4327796f, 32'h4381af07},
  {32'hc4730454, 32'h435fa10f, 32'h4311f504},
  {32'h44058c3e, 32'hc3614486, 32'h4223f0ed},
  {32'hc4ed1643, 32'h42e181da, 32'h43ab7d44},
  {32'h44aee328, 32'h3fcac33a, 32'hc3a7870a},
  {32'hc3fab288, 32'hc3e34dcb, 32'hc3842d6c},
  {32'h45012956, 32'h42eb14e6, 32'hc383656c},
  {32'hc4bf1f65, 32'h435c3140, 32'h42c38703},
  {32'h44a1a0da, 32'hc2ed6fc1, 32'hc41a8588},
  {32'hc48905ea, 32'h43745817, 32'hc3ed573f},
  {32'h43f022ce, 32'h440209cb, 32'h41f64de1},
  {32'hc4d0d380, 32'hc33dc2f5, 32'h42d49754},
  {32'h43d9b99c, 32'h4262271a, 32'hc34f2ab4},
  {32'hc38e80cc, 32'h432c1df6, 32'hc32d27d8},
  {32'h44934c6b, 32'h3f33947f, 32'h42e6c6ec},
  {32'hc4f8923b, 32'hc318483b, 32'hc38d2914},
  {32'h4501fb3f, 32'h43b735ba, 32'hc397fff8},
  {32'hc39f790e, 32'h43bca23d, 32'h4326e568},
  {32'h44ba96b2, 32'hc2c5671e, 32'hc375b654},
  {32'hc5068104, 32'hc358b895, 32'h4379fbb1},
  {32'h445db35e, 32'hc28aa0e9, 32'h430fdbd7},
  {32'hc4697cb0, 32'h3f8c5014, 32'hc19cfb19},
  {32'h44999728, 32'hc36c9665, 32'hc388e966},
  {32'hc48412e4, 32'h42e23868, 32'h42a30207},
  {32'hc352d238, 32'hc0bfbc71, 32'h431c528f},
  {32'hc42f0bb4, 32'h4179af42, 32'h436c3a63},
  {32'h43cdae54, 32'hc23bbb70, 32'h4281bdf8},
  {32'hc48f4cde, 32'h438887bb, 32'h43892c31},
  {32'h440901fc, 32'h434107ca, 32'h42a0430e},
  {32'hc4d88613, 32'hc178e2de, 32'hc28d3830},
  {32'h44af89e1, 32'h43a0bf60, 32'hc36a3c8a},
  {32'hc487069d, 32'h439f50e9, 32'hc1a6e242},
  {32'h445c5eb9, 32'hc3664979, 32'h43b557aa},
  {32'hc51373af, 32'hc3493d48, 32'h42e74617},
  {32'h440102f9, 32'hc35ae5fc, 32'h4055fadc},
  {32'hc4aa7674, 32'h440b1053, 32'hc0d6ba0c},
  {32'h451b6c6a, 32'hc24c79bd, 32'hc395bda8},
  {32'hc3ea0394, 32'h4350fb60, 32'h439b2582},
  {32'h44a3a50e, 32'h44100233, 32'hc1974c4e},
  {32'hc4c5e2a0, 32'hc38a6a97, 32'h42a12feb},
  {32'h4424bf2b, 32'hc344008e, 32'hc2a15bb4},
  {32'hc410ae0a, 32'h43ad7dac, 32'h43a0cd01},
  {32'h43a85940, 32'hc2f51d83, 32'h42e2f6b1},
  {32'hc3c55124, 32'hc1791498, 32'hc3814fc5},
  {32'h44ec008b, 32'hc181794a, 32'h42d6187a},
  {32'hc4becaf5, 32'hc1822f9e, 32'hc30bb7cf},
  {32'hc2302988, 32'hc2a594f3, 32'hc2eaf07e},
  {32'hc3b1e0c0, 32'hc3982f41, 32'hc3136b86},
  {32'h445c8fc5, 32'hc36f0c29, 32'hc2b99f80},
  {32'hc3da8769, 32'h437463a4, 32'h42c4bfb5},
  {32'h448ec7aa, 32'hc232dd53, 32'hc33396e1},
  {32'hc2f6ee80, 32'hc2f5fb16, 32'hc0b253ae},
  {32'h44097dd8, 32'h4382e7d3, 32'h4387e6d5},
  {32'hc4edb754, 32'h42c61990, 32'hc3980331},
  {32'h44813204, 32'h43912d58, 32'h435e711b},
  {32'hc4f14543, 32'h435806a9, 32'h439b8a1a},
  {32'h44c184c4, 32'hc1c0ecde, 32'hc2a43305},
  {32'hc49d641b, 32'h42d8b4cb, 32'hc344378c},
  {32'h44d30c3e, 32'h43c10aeb, 32'hc2c640dd},
  {32'hc4d39a42, 32'hc2974650, 32'h4376c85f},
  {32'h449763cc, 32'hc29b0c28, 32'h43b11954},
  {32'hc4a69295, 32'hc2a748d2, 32'h43d97a93},
  {32'h4416a31c, 32'h429a5164, 32'h430c282f},
  {32'hc4ca9c23, 32'hbec2de2e, 32'hc182cb20},
  {32'h44f29a60, 32'hc3b7ca0f, 32'hc3abf103},
  {32'hc3d37cd3, 32'hc2166908, 32'hc3bf85e2},
  {32'h44bc7bec, 32'h43298f63, 32'h43c0244f},
  {32'hc4edc3c6, 32'h4312f540, 32'hc3b39eb2},
  {32'h441a3c32, 32'h430be1a5, 32'hc302d5c0},
  {32'hc50e59b4, 32'h4393cf14, 32'h42d95350},
  {32'h44f27b06, 32'hc39bf28a, 32'hc2bc7064},
  {32'h4256c680, 32'h4398d3d0, 32'hc21c8bf5},
  {32'h4444bd08, 32'h42b19cf5, 32'h438ddfa6},
  {32'hc4cdcf97, 32'h432bcfff, 32'h43affabd},
  {32'h43a39303, 32'hc37147bd, 32'h4388800f},
  {32'hc400456a, 32'h43dc63a6, 32'h4308413d},
  {32'h44157dad, 32'hc429b8c0, 32'h4375a95d},
  {32'hc4d7f711, 32'h41930d12, 32'h434cbe52},
  {32'h4501ffca, 32'h42fdfc20, 32'h43a33acb},
  {32'hc48b74de, 32'hc2cba031, 32'h438058a6},
  {32'h447cde82, 32'h435f2d63, 32'hc3dde85e},
  {32'h430b295b, 32'hc39ef320, 32'hc3bb8a49},
  {32'h44dafa6f, 32'hc3a24546, 32'hc23cc793},
  {32'hc503e7be, 32'hc208ba76, 32'hc3c9f435},
  {32'h4455e64a, 32'h43780321, 32'h41f95df0},
  {32'hc4b665b0, 32'h43ed35b1, 32'h436aaf45},
  {32'h4495cd6c, 32'hc3327f79, 32'hc39a7cd3},
  {32'hc38886f9, 32'hc32f0459, 32'hc2d58641},
  {32'h4503b4e8, 32'hc36b1fec, 32'h42d411a6},
  {32'hc4908731, 32'h427ff7f1, 32'hc3d091e3},
  {32'h450fbdfc, 32'h426a52a7, 32'h4383979e},
  {32'hc41987a8, 32'hc32078d0, 32'hc39e2866},
  {32'h450d3036, 32'h43038ce5, 32'hc2cd29a8},
  {32'hc4faaf15, 32'h44409462, 32'h4320d704},
  {32'h44629734, 32'hc2226feb, 32'h43bbe2ba},
  {32'hc3557ace, 32'h43a6be8a, 32'hc38757ae},
  {32'h44a4f2a2, 32'hc3867c39, 32'h4215e63d},
  {32'hc4e3e5c0, 32'h434f3b22, 32'hc367e829},
  {32'h451fa06d, 32'hc3d25777, 32'h42e46065},
  {32'hc2c94be0, 32'h42db46e5, 32'hc36bc9c4},
  {32'h43e3876c, 32'hc383d6a6, 32'h41bbe1cc},
  {32'hc500b6aa, 32'h4373b641, 32'hc34c7d15},
  {32'h44c207f5, 32'h424cbbbe, 32'h423c8327},
  {32'hc2308297, 32'hc3815611, 32'h413be0a0},
  {32'h440254c6, 32'hc2026f95, 32'hc3003698},
  {32'hc49aeaca, 32'hc315b4f4, 32'h4361624e},
  {32'h446340e8, 32'h42a0c7a8, 32'hc233d3a9},
  {32'hc2d0b6d0, 32'hc2ee3413, 32'h43a1dff7},
  {32'h44d07888, 32'hc297b4d4, 32'hc3f38444},
  {32'hc49207bd, 32'h43fc21ac, 32'h437af780},
  {32'h430a362a, 32'hc3a7776b, 32'hc39d1007},
  {32'hc397b190, 32'hc09f0c4a, 32'hc38b1654},
  {32'h44f243ca, 32'hc3dafb81, 32'h43205951},
  {32'hc4bb0aca, 32'hc22b6180, 32'h42960a43},
  {32'h443398aa, 32'h434674bd, 32'h4226fe23},
  {32'hc500bcf8, 32'hc362425e, 32'hc33732c1},
  {32'h42ad67a0, 32'h43e6f78e, 32'hc36e2302},
  {32'hc4ea891f, 32'hc388b593, 32'h432d201f},
  {32'h45235a24, 32'hc2549b16, 32'hc34c22f3},
  {32'hc42eb628, 32'h43270f67, 32'hc2a8235b},
  {32'h44ca7c45, 32'hc2c99592, 32'hc28f8042},
  {32'hc511fbd7, 32'h423fe84b, 32'hc3b3c4ae},
  {32'h44696f17, 32'h433879c0, 32'hc20a830d},
  {32'hc4c1fad4, 32'h43c26fb4, 32'hc2a40ef6},
  {32'h44ec323e, 32'hc25d7c7e, 32'h43c30d03},
  {32'hc38a505c, 32'h430e5e09, 32'h4326448c},
  {32'h44e0afba, 32'hc2845dc2, 32'h418b7d6b},
  {32'hc51e6800, 32'h43072df9, 32'h438c1c51},
  {32'h44d310ef, 32'hc38245fa, 32'hc359cd4b},
  {32'hc5124cf4, 32'h430c55e3, 32'h42d9a27a},
  {32'h4434ee17, 32'hc111f251, 32'h425612eb},
  {32'hc50dfa9b, 32'hc3c6327e, 32'hc218d718},
  {32'h451b37c6, 32'hc3687841, 32'hc26abd0f},
  {32'hc483d4d0, 32'h4342cf32, 32'h42047dfc},
  {32'h45134210, 32'hc3696ee2, 32'hc154082b},
  {32'hc4767975, 32'hc38a9162, 32'h42bc8f39},
  {32'h44bf343a, 32'h440273c2, 32'hc29141d3},
  {32'hc4d5e0cc, 32'hc2b9db67, 32'h43578f31},
  {32'h44b415e2, 32'hc2dd369f, 32'h43275d71},
  {32'h430c37fb, 32'h42104151, 32'hc1493bed},
  {32'h44ebfa9e, 32'h42a87b5f, 32'h4319dd64},
  {32'hc4a6a19a, 32'h41f51243, 32'h423af7f4},
  {32'h42e4d790, 32'hc36ec8b4, 32'hc36a9fd0},
  {32'hc3851d8a, 32'hc33641fc, 32'hc3116b49},
  {32'h446ccba2, 32'hc3881e2b, 32'hc2b5c955},
  {32'hc4ce776d, 32'h43bcdfb5, 32'hc41ad967},
  {32'h450c0572, 32'hc39548c4, 32'hc37a2aae},
  {32'hc4de1656, 32'h4226ecf7, 32'hc39522d3},
  {32'h4487bdb6, 32'h43bf87e9, 32'hc35762b6},
  {32'hc49702ca, 32'hc325285b, 32'hc385a08b},
  {32'h450ed10a, 32'h43b8b2d0, 32'hc1e2fa7c},
  {32'hc3691dfc, 32'h431d6c31, 32'h42a67fc8},
  {32'h4355f9a8, 32'h44013cbd, 32'hc28a7413},
  {32'hc403be36, 32'hc2d43993, 32'h42b861c4},
  {32'h42db1a90, 32'h439e7663, 32'hc21846cf},
  {32'hc42ff9d6, 32'hc30add51, 32'hc32c422b},
  {32'h44c27b5c, 32'hc3084c46, 32'h4304675c},
  {32'hc4ff94f2, 32'hc2ed29fd, 32'hc3048721},
  {32'h44da1614, 32'h439e3048, 32'h43e7cde6},
  {32'hc3d108f8, 32'h4390f69c, 32'hc33d2fed},
  {32'h448d7c78, 32'hc38abb53, 32'hc3bef4f2},
  {32'hc4b71776, 32'hc29a0094, 32'hc318c60a},
  {32'h440333b5, 32'hc1d588ef, 32'hc3315cc4},
  {32'hc4a7befe, 32'h42a7cc28, 32'hc377f216},
  {32'h4511c8c9, 32'hc271a976, 32'h42145e39},
  {32'hc3244db8, 32'h43b083f8, 32'h43ce8f47},
  {32'h44779950, 32'hc304f1bd, 32'hc387a95e},
  {32'hc4958668, 32'hc3d55137, 32'h41a121a7},
  {32'h439ff13c, 32'hc31e09e3, 32'hc408ac4b},
  {32'hc44eaf98, 32'h41c972f7, 32'h43a40cad},
  {32'h4410a886, 32'hc20ac290, 32'h42ae5228},
  {32'hc4969311, 32'hc2d2a300, 32'h42add76a},
  {32'h43ebe308, 32'h42821168, 32'hc3552862},
  {32'hc4ca311a, 32'hc3327f52, 32'h4222350a},
  {32'h448fb085, 32'hc1465e19, 32'hc384eabd},
  {32'hc2d81780, 32'hc1b8cabc, 32'hc3864a7e},
  {32'h44012030, 32'hc18b6ca5, 32'h434e3586},
  {32'hc50e8540, 32'hc336838d, 32'h42b48d9d},
  {32'h4348e838, 32'hc1f51b57, 32'hc2a2dfcb},
  {32'hc50a4891, 32'h43a99771, 32'hc2b0a844},
  {32'h445264cc, 32'h4354e70d, 32'h43d89a4f},
  {32'hc4c76b23, 32'h43bb7712, 32'h436566ca},
  {32'h44fce585, 32'hc3113565, 32'h430299c0},
  {32'hc49b4fd7, 32'h4390c287, 32'h4382eff4},
  {32'hc1721800, 32'hc40764f7, 32'hc38d80dd},
  {32'hc3c82048, 32'hc2adca1a, 32'hc16e165d},
  {32'h4404a438, 32'hc39eb9c5, 32'hc1d579c6},
  {32'hc4e1f2fa, 32'h43a07efb, 32'hc2c2a05c},
  {32'h44ad8db6, 32'h43b70f55, 32'h434ec0f0},
  {32'hc5001fde, 32'h3fb9a4d2, 32'hc3b9c278},
  {32'h450cce67, 32'hc3c353c6, 32'hc2ac1fad},
  {32'hc41b2075, 32'hc3111d97, 32'h421a7f2d},
  {32'h44d857bb, 32'h42c270f0, 32'hc39b96d4},
  {32'hc46210ac, 32'h42c19dfe, 32'hc3ba10f0},
  {32'h43ab6ce4, 32'h41715050, 32'hc28c5e34},
  {32'hc3cc50b8, 32'hc3dd2d3d, 32'hc1b9a0fa},
  {32'h45102022, 32'hc26bd1f7, 32'hc3241595},
  {32'hc4ec347e, 32'h43028af6, 32'hc3702475},
  {32'h4410377e, 32'hc27fe66a, 32'hc292fb31},
  {32'hc458b1a4, 32'h438bd9ea, 32'h432c9222},
  {32'h449b2378, 32'hc38ae520, 32'hc37f1f4d},
  {32'hc3d40f37, 32'hc2637e49, 32'hc3bdf0d3},
  {32'h43f7ddcd, 32'hc4064700, 32'hc3560c0a},
  {32'hc4a79bd4, 32'hc3be0fe8, 32'h41ddb7f0},
  {32'h44878270, 32'h437257bf, 32'hc39a0d38},
  {32'hc4b26105, 32'h431e2883, 32'hc340cfaf},
  {32'h4443a8b3, 32'hc3a6a5cc, 32'hc2918634},
  {32'hc40f5728, 32'hc307b759, 32'hc2afbbdc},
  {32'h45130aec, 32'hc3cb1f04, 32'h42ebe22d},
  {32'hc4e230b6, 32'hc3c40bcd, 32'h421c1f1a},
  {32'h44225b4c, 32'hc3c6f797, 32'hc3886450},
  {32'hc4e3e3fa, 32'h4281ce14, 32'h3f92a660},
  {32'h449b4012, 32'hc2eb313f, 32'hc23495c4},
  {32'hc49701aa, 32'hc3e0b623, 32'hc2fd384d},
  {32'h449fc4a4, 32'hc404fe83, 32'hc3a10044},
  {32'hc32071e1, 32'h4110641c, 32'h40e86e58},
  {32'h4358c710, 32'h43cd5272, 32'hc24d21d2},
  {32'hc4a815fc, 32'h42c1b262, 32'hc1aa9682},
  {32'h449bb07c, 32'h40a16172, 32'hc2e2d169},
  {32'hc4feefb6, 32'h42db644c, 32'h43a23535},
  {32'h44c1ab78, 32'hc292b7be, 32'hc3d81807},
  {32'hc4f3b64e, 32'hc39b2814, 32'hc37144e4},
  {32'h44375434, 32'h428f1eda, 32'hc33ed76b},
  {32'hc502f1e3, 32'hc253e528, 32'hc2032b11},
  {32'h44de9b63, 32'hc281f3c9, 32'h424b0789},
  {32'hc4c191e1, 32'h43935a32, 32'h43bd6c36},
  {32'h451e1d9d, 32'hc303386f, 32'hc3b8c5af},
  {32'hc49bd6f5, 32'hc2f225d1, 32'hc3ae9412},
  {32'h4421db50, 32'hc3e6c9fe, 32'hc360ff98},
  {32'hc4150f20, 32'hc34c5daa, 32'h4261e8a9},
  {32'h44046b9c, 32'h4220a55e, 32'hc40429fa},
  {32'h42ef5bce, 32'hc232ca8c, 32'h4371ca69},
  {32'h450ec84e, 32'hc2a078e8, 32'h439497ae},
  {32'hc2a6b3e4, 32'h42f44b06, 32'hc0fe47ac},
  {32'h45191d56, 32'hc345f022, 32'hc3350d85},
  {32'hc41588e9, 32'h43cbb448, 32'h429b41f8},
  {32'h44ad3b74, 32'hc3608eab, 32'h420835c5},
  {32'hc3d20584, 32'h4356e4a1, 32'h43c52886},
  {32'h445fbd7a, 32'hc2b5a8c0, 32'h43c64fcd},
  {32'hc3c67f6d, 32'hc3122caf, 32'h4104ce05},
  {32'h44d1b35c, 32'hc39d41ed, 32'hc3dfd80c},
  {32'hc4c4c577, 32'h43efa102, 32'h4298286f},
  {32'h44b190dc, 32'hc3896dcd, 32'hc2cad18b},
  {32'hc4c86916, 32'h43616272, 32'h43ff289b},
  {32'h44eaba50, 32'h43a7d561, 32'hc2af7ab9},
  {32'hc3bd5083, 32'hc3abc86e, 32'h438e7087},
  {32'h450d4974, 32'h4364cdd2, 32'h4293238c},
  {32'hc405266e, 32'h428d9cd8, 32'h433fc4dd},
  {32'h44db98e8, 32'hc2a5fb57, 32'h42f2e0c5},
  {32'hc4d7160a, 32'hc36803db, 32'h43a4b032},
  {32'h44aeec80, 32'h438ed7ee, 32'hc28f210c},
  {32'hc4f3384a, 32'hc39fabcd, 32'hc25d7140},
  {32'h44f27dde, 32'h40b16380, 32'h42886a76},
  {32'hc411ab5c, 32'h43357680, 32'h42e2d3c8},
  {32'h44bd77af, 32'h42bd589b, 32'hc39778d6},
  {32'hc2dc9620, 32'h4223eb5c, 32'h437c6bca},
  {32'h4397696a, 32'hc40c7f52, 32'h4376f1b4},
  {32'hc4d32e76, 32'h42ed5fc4, 32'h435560bd},
  {32'h44a00944, 32'hc366781e, 32'hc3e39d9b},
  {32'h44f4dd96, 32'h41dc9064, 32'h43705e9e},
  {32'hc26ccb50, 32'h43624a12, 32'h4361cfb8},
  {32'h44cdbb27, 32'hbf912354, 32'h4325633d},
  {32'hc3c47c8a, 32'hc34a4adb, 32'h42c235d6},
  {32'h44c38063, 32'hc34abb42, 32'h43423b6c},
  {32'hc416a7c0, 32'h42a62db6, 32'hc364c482},
  {32'h451db53c, 32'hc3d3d3a3, 32'hc031c3e9},
  {32'hc3c83563, 32'h42e7dfa3, 32'hc38e1e78},
  {32'h44719182, 32'hc367682c, 32'hc25d11ff},
  {32'hc4624f9c, 32'h43818ddc, 32'h43582f56},
  {32'h44f6b9f3, 32'hc3a111f7, 32'hc3391ba4},
  {32'hc4099d21, 32'hc3598d47, 32'h44146e9a},
  {32'h447ea15c, 32'hc35316a2, 32'hc24f66d0},
  {32'hc49543c0, 32'hc30c2458, 32'hc3153ed9},
  {32'hc2d26548, 32'hc30310d6, 32'h43b3b861},
  {32'hc503920c, 32'hc3948ee3, 32'h41c4df0e},
  {32'h449b404c, 32'hc2e4f124, 32'hc3b51e78},
  {32'hc3589088, 32'h419c9f49, 32'h42c1a690},
  {32'h440a3d7b, 32'hc36587a9, 32'h43a4afbf},
  {32'hc3fd8e62, 32'hc38b4839, 32'h42b0c50d},
  {32'h440b78ab, 32'hc113c71e, 32'h430193de},
  {32'hc48b00e8, 32'hc3a9214a, 32'h428d89bd},
  {32'h44b2119b, 32'h4365c8d3, 32'hc36f9409},
  {32'h421e33c0, 32'h414fa5ad, 32'h43b6e98e},
  {32'h44c62313, 32'hc234750c, 32'hc39e9b90},
  {32'hc0d9da88, 32'h428c68ca, 32'hc327374c},
  {32'h446819bd, 32'h429bd974, 32'hc3c366ce},
  {32'hc473a8ce, 32'hc347992a, 32'hc2ef240c},
  {32'h4426f140, 32'h43020198, 32'hc3ab8a22},
  {32'hc36d215a, 32'h43802f71, 32'hc31153ee},
  {32'h44983561, 32'h428f7c63, 32'hc21efa49},
  {32'hc49e63df, 32'hc1c37fc1, 32'h43c3aaf9},
  {32'h449c7a77, 32'h42ff7027, 32'h4364e2e9},
  {32'hc3459737, 32'hc26d4f6d, 32'hc3532bc5},
  {32'h44e42d73, 32'hc35e8a63, 32'hc377aafe},
  {32'hc435897b, 32'h43200a31, 32'h4212606a},
  {32'h4386cc10, 32'h42e5e1ac, 32'hc27d7557},
  {32'h439ac638, 32'h43007cba, 32'h43b26f57},
  {32'h43c2beec, 32'h436a79aa, 32'h43108294},
  {32'hc4a75033, 32'h431e98ca, 32'hc3a99013},
  {32'h44cabeae, 32'hc3028d41, 32'h43a06dc9},
  {32'hc3994522, 32'hbeaea9b5, 32'hc2ebbd75},
  {32'h43dc6cb0, 32'h436ef1a6, 32'h42351f4b},
  {32'hc4be3328, 32'hc1c2cc21, 32'hc29f6a91},
  {32'h438bac30, 32'h423a6230, 32'h43d78638},
  {32'hc3987820, 32'h438da4e7, 32'h419e9dd6},
  {32'h447a2d18, 32'h433c7777, 32'h433fcce2},
  {32'hc4899f51, 32'h43bc10ff, 32'hc381b500},
  {32'h450296c3, 32'h439473f0, 32'h41a7a972},
  {32'hc4d8547b, 32'hc2b0ee22, 32'hc280048d},
  {32'h4503957c, 32'hc1cfe87a, 32'hbfe77140},
  {32'hc42b30d4, 32'hc28127ec, 32'hc38b5774},
  {32'h44213ca0, 32'hc2ecf640, 32'hc36e59c6},
  {32'hc50d7b78, 32'hc36b8562, 32'h4356e670},
  {32'h45068bd4, 32'hc281838b, 32'h4172ff5e},
  {32'hc42a2154, 32'h429c250e, 32'h421ad617},
  {32'h4512e3d3, 32'h4387bae2, 32'hc36bbf19},
  {32'hc2fd87e5, 32'hc3833adf, 32'h4365a589},
  {32'h4506ba40, 32'h441a7a2d, 32'h43fcdd5b},
  {32'hc4078fc8, 32'h4391ba14, 32'hc47a35e8},
  {32'h44d05b4a, 32'hc2d17a9a, 32'h43417e08},
  {32'hc49b4bd2, 32'hc3664c24, 32'hc366bfaf},
  {32'h44ed9e97, 32'hc39c6262, 32'h42cd8a80},
  {32'hc4be9e6c, 32'h42bb6399, 32'h42ee5df6},
  {32'h44168806, 32'h43e92c0d, 32'hc3512d7b},
  {32'hc4f509c9, 32'h42c86a3a, 32'hc2318417},
  {32'h4418fdd4, 32'h438516f5, 32'h42517378},
  {32'hc4852b72, 32'hc2f77272, 32'hc27781fb},
  {32'h44de1c55, 32'hc344e822, 32'hc2675db3},
  {32'hc26a66b8, 32'hc26dddac, 32'h40808176},
  {32'h44bf97b6, 32'hc23ce097, 32'h42d86eda},
  {32'hc344a820, 32'h42452a73, 32'h41d6f60b},
  {32'h44ce8e9d, 32'h439997e1, 32'hc304ec45},
  {32'hc4fea7c8, 32'hc1b951e8, 32'hc3d06454},
  {32'h45216cc6, 32'h433e60d6, 32'h435253d4},
  {32'hc4e377b1, 32'h42c1e302, 32'hc36c9d28},
  {32'h448406b5, 32'hc2f67109, 32'h42133348},
  {32'hc4056aaa, 32'h43e9a060, 32'h438471df},
  {32'h43e92986, 32'h42bd6704, 32'hc258cb1f},
  {32'hc4c14105, 32'h439482a7, 32'hc23f554e},
  {32'h449352a7, 32'hc2a5191a, 32'h4336188d},
  {32'hc40c66fe, 32'h42ebae88, 32'hc35dd08b},
  {32'h439f8204, 32'h43acbf98, 32'h42c48b48},
  {32'hc4035a0e, 32'h43597d34, 32'hc3ff00e8},
  {32'h44d7419f, 32'h4296b6b3, 32'h42cf6997},
  {32'hc50e508e, 32'hc39ddc9c, 32'hc35055d4},
  {32'h445d8ee0, 32'h4308b97a, 32'hc32284cc},
  {32'hc4dddec4, 32'h43257223, 32'hc2e4a1aa},
  {32'h44b4b422, 32'hc337c757, 32'h43025aff},
  {32'hc4751474, 32'h436c3984, 32'h41dee667},
  {32'h4439cc78, 32'hc33d5042, 32'h42e888ee},
  {32'h421a5ff8, 32'hc2ddbd42, 32'h431730cb},
  {32'h451cd108, 32'h418a1eac, 32'h42b1ee7b},
  {32'hc4c7d422, 32'h43972c53, 32'hc3bddfef},
  {32'h44ddc4cd, 32'hc3687b49, 32'h42a4f77f},
  {32'hc4c949b6, 32'hc330979f, 32'h43a00c2d},
  {32'h450e8ce2, 32'hc2b8cdb1, 32'h42b5c3d8},
  {32'hc4f90b06, 32'h43c8aa02, 32'h42abe2f6},
  {32'h451647a8, 32'hc3bfe174, 32'h42c7f443},
  {32'hc51340d0, 32'hc3906fbe, 32'h43b06014},
  {32'h443aee13, 32'h436cb662, 32'h43a76d46},
  {32'hc4f3fcf0, 32'hc2ecad0f, 32'hc1f8595d},
  {32'h44e383b6, 32'h43e60fe0, 32'h44284d52},
  {32'hc420277d, 32'h43665988, 32'hc10f930c},
  {32'h449a7c6f, 32'h430ecf1f, 32'h4345dcf8},
  {32'hc40150d8, 32'hc38c2ffb, 32'h44024da9},
  {32'h442b239a, 32'h4308977e, 32'hc2b03821},
  {32'hc4628429, 32'hc39b5fd5, 32'hc3ddce37},
  {32'h44a1d9a0, 32'hc3e73648, 32'hc3cfce12},
  {32'hc4598ffe, 32'h43db3b69, 32'h41827a24},
  {32'h44a79757, 32'h4384bcff, 32'hc0b6b398},
  {32'hc3ea8e80, 32'h43603b1a, 32'h434bdc8a},
  {32'h448b12c8, 32'h42b9fe64, 32'h4322d4f6},
  {32'hc437f7e2, 32'hc1aad8ff, 32'hc2dcc7e0},
  {32'h44c688c1, 32'h42b05273, 32'h436f9e3a},
  {32'hc4a8c502, 32'hc38cb03e, 32'h4398a75a},
  {32'h44ce5200, 32'hc39ab4a4, 32'h437ca2a0},
  {32'hc4c8f927, 32'h4391b566, 32'hc2809bc5},
  {32'h4409694f, 32'h43831d13, 32'hc247750c},
  {32'hc4b01c63, 32'hc404d9f2, 32'h43a2dc9e},
  {32'h44a938a3, 32'hc38a7937, 32'h4374e8c7},
  {32'hc396b578, 32'hc3885318, 32'hc38c70de},
  {32'h44e9a59d, 32'h43e18e2c, 32'h43ddf730},
  {32'hc48b8018, 32'h427cdffe, 32'h43415764},
  {32'h44f659fc, 32'h42025026, 32'h4301ba49},
  {32'hc4df5575, 32'h4381c994, 32'h4316c7a5},
  {32'h450feefd, 32'h4193c5b6, 32'hc39887c0},
  {32'hc4c0ed28, 32'h42e1b208, 32'h43f35be6},
  {32'h4532d11f, 32'h43239393, 32'hc360aa27},
  {32'hc35cc120, 32'h43fbe713, 32'h4318f71c},
  {32'h44163ee4, 32'hc390cc20, 32'h4419d63e},
  {32'hc4c5be64, 32'h44330afd, 32'hc37bf3ab},
  {32'h42b2d098, 32'hc2b7b706, 32'hc32237cd},
  {32'hc48f5e7c, 32'hc383308f, 32'hc24dde99},
  {32'h4510a7dc, 32'hc303ac4e, 32'hc2e43910},
  {32'hc463aad0, 32'hc31d0510, 32'hc3021ad3},
  {32'h44e012ba, 32'h4394fd4f, 32'h4213b6f0},
  {32'h42d2b200, 32'hc37bdeec, 32'hc3e5e1c6},
  {32'h44073f48, 32'h42234e9c, 32'hc3294a4c},
  {32'hc4aa1aad, 32'h434cd6a6, 32'h439bbe7b},
  {32'h44efa3cf, 32'h4328deac, 32'h41cc56af},
  {32'hc428fec2, 32'hc3257d99, 32'hc2b7f7cc},
  {32'h449e9f84, 32'h44045553, 32'h431ebd1d},
  {32'hc425c374, 32'hc3adf389, 32'h427ead44},
  {32'h447cb631, 32'hc368c809, 32'h4207c930},
  {32'hc4a7340e, 32'h4322c626, 32'h4111000e},
  {32'h44bb3f7b, 32'h4387b41e, 32'h418a2b6d},
  {32'hc40c6030, 32'hc3617113, 32'h43017421},
  {32'h44db0854, 32'h420f19ee, 32'hc2f5d725},
  {32'hc46d821e, 32'h43690265, 32'h438eb063},
  {32'h44c426f5, 32'h431253c2, 32'hc35c6d1e},
  {32'hc4454b1d, 32'h433410b2, 32'h42327352},
  {32'h42de07e4, 32'hc28e4255, 32'h43ae4127},
  {32'hc4bd6f0a, 32'hc23f1f5c, 32'h4355eb44},
  {32'h44326ec4, 32'h43570835, 32'hc398bb2d},
  {32'hc44de030, 32'hc2138a7a, 32'h42c11b4a},
  {32'h44a44168, 32'hc2db958e, 32'h416844a5},
  {32'hc4b14232, 32'h430e8039, 32'h4341d9e6},
  {32'h44f5edf5, 32'h40f06099, 32'hc2fb9fa1},
  {32'hc4d6ca0a, 32'hc2c05dc5, 32'h409ba21e},
  {32'h449492a1, 32'h418f832f, 32'h431a8756},
  {32'hc5111881, 32'h438c6dc2, 32'hc386e7ab},
  {32'h43c399fa, 32'hc3ad0de0, 32'hc15d3919},
  {32'hc5089aa4, 32'hc3bcefb1, 32'hc295e330},
  {32'h4512907d, 32'hc293f091, 32'h4391fcea},
  {32'hc28e6ea0, 32'hc229bbbc, 32'h41253e95},
  {32'h446368cc, 32'h437e9245, 32'hc20938e2},
  {32'hc485f4f8, 32'hc2fa5b53, 32'h42f0c4ef},
  {32'h4452e470, 32'hc18f512f, 32'hc2973614},
  {32'hc3bf23ed, 32'hc3e95a51, 32'h4350b978},
  {32'h444f62b2, 32'h42c1612e, 32'hc299ce8c},
  {32'hc5074bdd, 32'h43aeb0ef, 32'hc28e2c44},
  {32'h44e972b3, 32'hc2873cae, 32'hc349a54f},
  {32'hc407406c, 32'hc31fffca, 32'hc2a09bb6},
  {32'h45059bb8, 32'h3f8fa34a, 32'hc1f54ad1},
  {32'hc39a3b4f, 32'hc31cb79f, 32'hc1c8510c},
  {32'h44127f78, 32'h436a6921, 32'hc18c0210},
  {32'hc50414c1, 32'hc292fb0c, 32'hc20ff291},
  {32'h44b56550, 32'h43814de9, 32'hc1d78e47},
  {32'hc4808f6a, 32'hc39e3236, 32'h43044c46},
  {32'h44ef20c2, 32'hc285ea42, 32'hc31100e7},
  {32'hc285a37f, 32'h43930217, 32'h4360eefd},
  {32'h448db2d1, 32'hc2d74f22, 32'h3fafe060},
  {32'hc3f1e6f3, 32'h43acd123, 32'hc38e829e},
  {32'h43f327c4, 32'h43725e75, 32'hc2953063},
  {32'h40f2f600, 32'h420acdb2, 32'h43c8558c},
  {32'h44819b69, 32'h43178174, 32'hc398a15c},
  {32'hc48c4425, 32'hc3589259, 32'h431d5505},
  {32'h41d77a80, 32'hc38aea27, 32'hc1d503ce},
  {32'hc38935a7, 32'h43d170f1, 32'h4319108c},
  {32'h449d75de, 32'hc224f1bc, 32'h440e2fdb},
  {32'hc4ad27ee, 32'h43106641, 32'hc326e281},
  {32'h436967c0, 32'h434502a8, 32'hc0d076e8},
  {32'hc3fd619a, 32'h42e6010b, 32'hc217b2c5},
  {32'h44e327cb, 32'h42c6cbc0, 32'h435a8883},
  {32'hc3bcad05, 32'h4362fa70, 32'h43c1200d},
  {32'h450e6ddf, 32'hc3a0061c, 32'h42b9ef4c},
  {32'hc4020022, 32'hc287eb4d, 32'h438bcb44},
  {32'h44803b51, 32'h4342fd62, 32'h437f17a7},
  {32'hc41abef6, 32'h4374c994, 32'h43c8b6c5},
  {32'h45146935, 32'h4393df15, 32'h43a9993a},
  {32'hc4ca3a1e, 32'h421e774e, 32'hc32dfbdc},
  {32'h42cd2692, 32'hc376e279, 32'hc2d4a4fe},
  {32'hc4ff1dd5, 32'h4398ec01, 32'h429807a8},
  {32'h4497f126, 32'h43a76d03, 32'h430a6136},
  {32'hc44aa988, 32'hc2d061da, 32'hc35790f8},
  {32'h446b64c3, 32'hc393ea1a, 32'h4277ec52},
  {32'hc473aa93, 32'h42db1cee, 32'hc2dca254},
  {32'h4297fe78, 32'hc2bfecec, 32'hc36aa48c},
  {32'h3f9f5800, 32'h42d4e3a5, 32'h3f9acca0},
  {32'h4420a7fa, 32'h43e5e58e, 32'h42e46ad1},
  {32'hc485b33a, 32'h42c6e5b6, 32'hc1f6c210},
  {32'hc2d3d040, 32'hc17dbf25, 32'h42e5003a},
  {32'hc4c4ae2c, 32'hc3c050c4, 32'hc3023643},
  {32'h4509b8dc, 32'h42ef4907, 32'hc393b25c},
  {32'h42ec8428, 32'hc3879b27, 32'h432331d1},
  {32'h4497d090, 32'h43d2aa54, 32'hc332ec9f},
  {32'hc5186bcb, 32'h4325f8ab, 32'h42a5f447},
  {32'h44ba900d, 32'hc3cd6290, 32'h431222dc},
  {32'hc49767ac, 32'hc0f48272, 32'h42a2f98e},
  {32'h449fff6f, 32'h4345f1e6, 32'h4302df1a},
  {32'hc4afc5b5, 32'h420d195e, 32'h42cb9b4b},
  {32'h4499ab5c, 32'h4383ac21, 32'hc33a4eee},
  {32'hc4dbf4d5, 32'hc350ba0c, 32'h431ccdec},
  {32'h44dfa074, 32'hc350d46a, 32'h4359400d},
  {32'hc4a079c7, 32'h43680d52, 32'h41b1fcf2},
  {32'h43f1e1db, 32'hc2900c3b, 32'hc2f98609},
  {32'hc3edbaea, 32'h4418a584, 32'h429593ad},
  {32'h4496e6a8, 32'hc1c4866b, 32'h41319130},
  {32'hc48ada31, 32'h4337ac01, 32'hc303da38},
  {32'hc224b000, 32'hc37806f9, 32'h42e4414f},
  {32'hc440cadd, 32'h42433f2f, 32'hc2eff0e2},
  {32'h44dc4b4c, 32'h430cc6a6, 32'h440daa2b},
  {32'hc463c614, 32'h42ed0ffa, 32'h432893b7},
  {32'h44b65de2, 32'h42d401d5, 32'hc2e30cf9},
  {32'hc460a546, 32'hc2ed1c7f, 32'h438e5dc0},
  {32'h44f3e23f, 32'hc2cd9be5, 32'h43203d07},
  {32'hc441b732, 32'hc37931b6, 32'h42abae63},
  {32'h4456be1c, 32'h434f3a97, 32'h43d321a7},
  {32'hc44ea8ce, 32'h4301eaa6, 32'h43557052},
  {32'h4442f8b2, 32'h437f2705, 32'hc3186ec9},
  {32'hc3aa2f3e, 32'h433aa363, 32'h435d9b6e},
  {32'h43a8fe24, 32'hc3988136, 32'h43c3afba},
  {32'hc50f4511, 32'hc1821e51, 32'h4421395e},
  {32'h4436dd1e, 32'hc2291b1a, 32'h428b5130},
  {32'hc503e20a, 32'hc3390c56, 32'hc41c7366},
  {32'h4443f1b4, 32'h43df197d, 32'hc32957f8},
  {32'hc510b40d, 32'hc2e3523b, 32'hc380b69c},
  {32'h4458ea48, 32'h4426c3c8, 32'h4336edfe},
  {32'hc4903132, 32'h4359d99a, 32'h438dd086},
  {32'h44360685, 32'hc33d97d8, 32'h4341c2ae},
  {32'hc494ad77, 32'h418cad2d, 32'h43f98974},
  {32'h450b3ffd, 32'h410ff89c, 32'h434ce4d1},
  {32'hc4f69dbb, 32'hc0c768d6, 32'h43654fac},
  {32'h444f57bc, 32'hc3127846, 32'hc4028e08},
  {32'hc4b513c9, 32'hc39cf692, 32'h432aa6b0},
  {32'h450127ad, 32'hc1bfb57f, 32'h42bc2e5a},
  {32'hc4c70dcb, 32'h433f5d3f, 32'hc0e424e4},
  {32'h44a684f4, 32'h423df34d, 32'hc366dda7},
  {32'hc44a592f, 32'h43a8fc5d, 32'h433598c3},
  {32'h44e65396, 32'hc31d837c, 32'hc3468c2e},
  {32'hc4061b32, 32'hc3290c91, 32'hc1c349f9},
  {32'h4431a68c, 32'hc353cb13, 32'hc312ff14},
  {32'hc47444d5, 32'h438b7e6e, 32'hc308c59b},
  {32'h45126ede, 32'hc29d85b0, 32'hc236da7f},
  {32'hc4a8fb95, 32'hc3007b3d, 32'h438ce4fc},
  {32'h4505ea0d, 32'h43dc30d7, 32'hc318fc7b},
  {32'hc50a21e4, 32'h425f2fcc, 32'h42edc494},
  {32'h4480371f, 32'h42f10b3d, 32'hc34fa940},
  {32'hc4b303ce, 32'hc22ce4b9, 32'h41dcfa74},
  {32'h43de6409, 32'h435e81a5, 32'hc33fa880},
  {32'hc3f621b0, 32'hc3114ec0, 32'h4282785e},
  {32'h4343b6f0, 32'hc353df3c, 32'hc3688629},
  {32'hc4b98c88, 32'hc37b39f8, 32'hc295e72a},
  {32'h451913ea, 32'hc3d3f871, 32'h426f655d},
  {32'hc41e2d8f, 32'h43c8ef7e, 32'hc2dec3ed},
  {32'h43bc3c0a, 32'h42eb1292, 32'h425aa23c},
  {32'hc4607b80, 32'hc3c6f030, 32'h406ae9a4},
  {32'h44c2603f, 32'hc2d04295, 32'hc37c51a0},
  {32'hc3b0b79d, 32'hc0a79efc, 32'h43a658fa},
  {32'h44b4cf16, 32'hc1d69bb6, 32'h42cba1da},
  {32'hc46a0a97, 32'hc30be0d2, 32'hc2dde045},
  {32'h436c9410, 32'h4267705c, 32'h4383df3a},
  {32'hc2c1cf60, 32'h43456b95, 32'hc3985378},
  {32'h44e0c794, 32'hc2f747c8, 32'hc35075f2},
  {32'hc2e1ab38, 32'hc2c971ff, 32'h43c0df9f},
  {32'h43803d6a, 32'hc1922d3b, 32'hc31c0439},
  {32'h43dbed20, 32'hc30da265, 32'hc18f86d5},
  {32'h44aebb44, 32'hc354f555, 32'h436bfb08},
  {32'hc2843923, 32'h43b45e42, 32'hc39645c8},
  {32'h448421ca, 32'hc356beb9, 32'hc3ca963f},
  {32'hc3c25395, 32'hc2113478, 32'h43d068cc},
  {32'h44d71d32, 32'h4080fc06, 32'h43419081},
  {32'h42870260, 32'h4308cb86, 32'h43a8b3d0},
  {32'h44ebdd6c, 32'h429a708c, 32'hc3acb13d},
  {32'hc4ed94ae, 32'h423ade10, 32'h4238bcd6},
  {32'h4506edef, 32'h4124be71, 32'h437b5ae3},
  {32'hc5128368, 32'hc22b7ba4, 32'h436720d5},
  {32'h449de2fb, 32'hc3527700, 32'h42263572},
  {32'hc4ad03c6, 32'h42b9b32c, 32'hc2e5ea82},
  {32'h44c133a4, 32'hc3ae7204, 32'hc3eec434},
  {32'hc4b3d076, 32'h4370096b, 32'h417de52c},
  {32'h43ba68d0, 32'h43b17245, 32'h43293c15},
  {32'hc4a8e449, 32'h43259520, 32'h3f56e164},
  {32'h448c9e68, 32'hc1e9b6f5, 32'h41ffbe73},
  {32'hc4b2673b, 32'hc2208ceb, 32'h431cb57c},
  {32'h445c18a1, 32'hc28325b0, 32'h4268bc74},
  {32'hc4643c26, 32'hc19aff5a, 32'h430efd67},
  {32'h44330d6c, 32'h438e7145, 32'hc1ece2df},
  {32'hc4f9902e, 32'hc2fdfd40, 32'h43b4327d},
  {32'h43f5841c, 32'h4253555d, 32'h43062fa0},
  {32'hc5106434, 32'h43350c69, 32'hbec91018},
  {32'h44968c97, 32'h438ef173, 32'h43c39a4c},
  {32'hc50b2d69, 32'hc335fa4f, 32'h4258a71c},
  {32'h4416f9ed, 32'h4374b0f8, 32'hc2cd1c09},
  {32'hc4d64e10, 32'hc20c8cc3, 32'hc3bd9f79},
  {32'h438a5c34, 32'hc236e94c, 32'hc257b36c},
  {32'h428cfc7c, 32'h42a6b649, 32'h4127a160},
  {32'h43e37cbe, 32'hc33c4811, 32'hc3fab8a7},
  {32'hc4d61f54, 32'h41a4dc1c, 32'hc3700831},
  {32'h44ebd86d, 32'hc2f472e3, 32'hc396e4e3},
  {32'hc4a86304, 32'hc381f24f, 32'h43599824},
  {32'h449eeb12, 32'h429fb5e4, 32'hc357cb15},
  {32'h42ef5ae0, 32'hc1559aea, 32'h424612f1},
  {32'h446f5289, 32'h423d898d, 32'h431d2b83},
  {32'hc341d273, 32'h438a65d4, 32'hc2deb4be},
  {32'h448c7f18, 32'hc2c4cf10, 32'hc3605125},
  {32'hc4ecff4e, 32'h4349d719, 32'h439e5038},
  {32'h44dc5764, 32'h43398eda, 32'hc3a4479e},
  {32'hc4c17396, 32'hc2d3387a, 32'h43960024},
  {32'h4465bb79, 32'hc25011c5, 32'h42a28af2},
  {32'h429482b8, 32'hc2e4d39e, 32'hc19bf99e},
  {32'h44e48798, 32'hc346e77c, 32'hc3af38d2},
  {32'hc4f3ef50, 32'hc2e509c7, 32'hbf004727},
  {32'h44e43ba8, 32'h42d9cea5, 32'h42f0d251},
  {32'hc48867c2, 32'hc2b98672, 32'hc2e7d6ab},
  {32'h44c66bc4, 32'hc39ab4d0, 32'hc3b2a654},
  {32'hc3ee1eb8, 32'hc351da3d, 32'hc38646dd},
  {32'h44a7320a, 32'hbf271bac, 32'hc341095f},
  {32'hc452b4e5, 32'hc2349ad4, 32'hc3145c8e},
  {32'h4454b17a, 32'hc3c8f66b, 32'h43a304a8},
  {32'hc36d574c, 32'h438446b6, 32'hc3f43452},
  {32'h4400f5c8, 32'h4326f93f, 32'h4358da4f},
  {32'hc476b4b4, 32'h4229868c, 32'hc31d5cbe},
  {32'h44d560dc, 32'hc380e83c, 32'h42f63e17},
  {32'hc4eefc98, 32'hc2dac1ba, 32'hc2c4bb70},
  {32'h44f77be1, 32'hc39d47fa, 32'hc34f6b76},
  {32'hc5178763, 32'h43c290e6, 32'h4292beb5},
  {32'hc2063d90, 32'h437386e3, 32'hc0bc1076},
  {32'hc4b804b7, 32'hc40136b2, 32'h4236f05e},
  {32'h426ffab0, 32'h4366bd4d, 32'h42c39acd},
  {32'hc4c4705a, 32'hc3cd9ca3, 32'h43929bc0},
  {32'h4447f30e, 32'h41988aba, 32'hc3184d54},
  {32'hc45afe92, 32'h424b2057, 32'hc13d1150},
  {32'h44808312, 32'hc2cf5758, 32'hc3d02198},
  {32'hc4e3765c, 32'hc34bf12d, 32'hc14af2ea},
  {32'h44e77193, 32'h40ad67b4, 32'h433d9702},
  {32'hc50ad42a, 32'h41663e2a, 32'hc2494d97},
  {32'h44bd2d7d, 32'h423dd9ea, 32'hc38c5eee},
  {32'hc496619e, 32'hc394a45b, 32'h423dd73c},
  {32'h424d7190, 32'h42e54648, 32'h4286755a},
  {32'hc4876743, 32'hc329ac2b, 32'h4373253f},
  {32'h44571096, 32'hc206a430, 32'h43a4381e},
  {32'hc42d4b09, 32'hc26718f2, 32'h433d01df},
  {32'h44afd056, 32'hc37ac194, 32'hc38b732e},
  {32'hc4c4b5ec, 32'h43574aa2, 32'hc29a2a88},
  {32'h43dcf904, 32'hc3bf4c04, 32'h43215bea},
  {32'hc414420e, 32'h429b3c32, 32'h43d60adf},
  {32'h41c78c80, 32'h419fb150, 32'h42bcb1fa},
  {32'hc4585c48, 32'hc39aef8a, 32'h418d7fc7},
  {32'h43dfec10, 32'hc36adf3b, 32'h4193c0e6},
  {32'hc3d96b84, 32'h4342dbd8, 32'h41b740b0},
  {32'h44e2a1a5, 32'h4311ba31, 32'h43d7666a},
  {32'hc5021af8, 32'h432dda84, 32'h42f32530},
  {32'h44db760f, 32'hc364669d, 32'h434e2334},
  {32'hc5157512, 32'hc209404f, 32'hc357c01d},
  {32'hc2eaba50, 32'hc23d7690, 32'h42d9f925},
  {32'hc4f3386c, 32'hc2b0b511, 32'hc3ca17ff},
  {32'h44bf5b26, 32'h436f0c21, 32'h4333de30},
  {32'hc5057b36, 32'h431c5ef6, 32'hc2383b02},
  {32'h450c16a4, 32'hc3d63ff4, 32'h43867585},
  {32'hc4738456, 32'h43f89a69, 32'h4279df0b},
  {32'h450cd8e3, 32'hc2e0528b, 32'hc39ba5c8},
  {32'hc4a3bcb6, 32'hc3f2a297, 32'h41293ca2},
  {32'h450f3699, 32'h420aae3a, 32'h42ee0b09},
  {32'hc4da3b62, 32'hc321a672, 32'hc3c5ee0b},
  {32'h447df194, 32'h43476efc, 32'hc09f7360},
  {32'h41fe3262, 32'hc3158837, 32'h4350857f},
  {32'h44d1538b, 32'h438ca0fa, 32'h4363fbfa},
  {32'hc4923e5a, 32'h43320695, 32'h437f613e},
  {32'h446ee7d2, 32'hc414845e, 32'hc1163fdc},
  {32'hc446476e, 32'hc2a2e610, 32'hc393227d},
  {32'h438252ac, 32'h43392cf4, 32'h438cd90b},
  {32'hc4d468b7, 32'h44045bcf, 32'hc3b08efb},
  {32'h43d9dcc8, 32'h422e3638, 32'hc3828cfd},
  {32'hc4e7be8c, 32'hc2951438, 32'hc2929a1e},
  {32'h431fd2ec, 32'h437366f5, 32'h432f1a9f},
  {32'hc522a6f8, 32'h439b88cf, 32'hc31448a8},
  {32'h44f24c52, 32'h42651e33, 32'hc38deb37},
  {32'hc4efe653, 32'hc334e74a, 32'h4250d011},
  {32'h44acbd63, 32'h43a73b11, 32'hc35fc8f3},
  {32'hc50f192d, 32'hc314f547, 32'hc3c1aa63},
  {32'h4514e623, 32'h4321ec3d, 32'h418ebe84},
  {32'hc4b7cb33, 32'hc1449c2d, 32'h41a2b2be},
  {32'h44721158, 32'hc2f361a9, 32'h4324f937},
  {32'h41cddc80, 32'hc3763e2b, 32'h428c5a67},
  {32'h43ab8a71, 32'hc3ae0596, 32'hc303752b},
  {32'hc47258a6, 32'hc14ec888, 32'hc3c744fd},
  {32'h44ca6381, 32'hc33ce57c, 32'h43937db2},
  {32'hc509bf79, 32'h3fb50c00, 32'hc34d9e42},
  {32'h44cf8194, 32'h431bb5ca, 32'h430df4a1},
  {32'hc5010e00, 32'hc37d8130, 32'h4211efd0},
  {32'h44338ed4, 32'h4313e976, 32'hc1b3adde},
  {32'hc431aa70, 32'h41abca42, 32'hc3ae7c38},
  {32'h44e3c6b3, 32'hc3dd8a61, 32'h428d0267},
  {32'hc50bb88d, 32'hc3679c42, 32'h43384ec3},
  {32'h448851e4, 32'h42af0ddc, 32'h4364eb6e},
  {32'hc52061ab, 32'h42df4274, 32'h41bdf484},
  {32'h420d86d8, 32'hc390c9e0, 32'hc1e20ab7},
  {32'hc4c02664, 32'h433c3419, 32'h40c3ce14},
  {32'h442b105a, 32'h43b5d08d, 32'hc2c4f3d3},
  {32'hc49fe3ec, 32'hc33dc919, 32'h424adba4},
  {32'h446af0d0, 32'hc3b6c8b7, 32'h42bacf4c},
  {32'hc26315da, 32'h424e8e20, 32'hc389d211},
  {32'h450df51e, 32'h427a2a6a, 32'h40b94140},
  {32'hc4cff78c, 32'hc39e912e, 32'hc30ae0e5},
  {32'h4486b753, 32'h43c315d3, 32'h4159ade6},
  {32'hc50b00eb, 32'hc399df3c, 32'hc36e61c3},
  {32'h44c34bef, 32'h43535186, 32'h443c94bd},
  {32'hc4e3c9d5, 32'hc2b01ede, 32'h43716e35},
  {32'h44567c25, 32'hc20de698, 32'hc314e01b},
  {32'hc4b7f46a, 32'hc1e0a168, 32'h41336724},
  {32'hc4c40f8e, 32'hc21bddbb, 32'h40521e6d},
  {32'h44b14b10, 32'h426e88ee, 32'h438f5c2d},
  {32'hc3d6d0a8, 32'hc3c2a281, 32'hc3754317},
  {32'h44597a34, 32'h42e0a2d4, 32'h43a3df50},
  {32'hc4e4915e, 32'hc3865ae5, 32'hc31c934d},
  {32'h44b32af0, 32'h400fb979, 32'hc3293ee2},
  {32'hc4c695aa, 32'h421816d4, 32'h41c0cf95},
  {32'h44f93a9c, 32'hc2db96cd, 32'hc282a92b},
  {32'hc4bcf306, 32'h43cd10ca, 32'h43e2e78c},
  {32'h45057b37, 32'hc2b9e893, 32'h433d5827},
  {32'h43024230, 32'hc262ca67, 32'hc3d7906f},
  {32'h440b0ffa, 32'h4329f3ba, 32'h42288282},
  {32'hc4d65b62, 32'h42bce1ec, 32'hc32d2dec},
  {32'h445077fa, 32'h4197a4b1, 32'h4234cfe5},
  {32'hc4201b36, 32'h430b51f7, 32'hc0f41f48},
  {32'h444734cc, 32'hc292e8c2, 32'h43e43803},
  {32'hc4e88786, 32'hc282c674, 32'h4386085b},
  {32'h44d884e7, 32'h42f74db3, 32'hc36fd3fb},
  {32'hc4048427, 32'hc3779f99, 32'h4280b172},
  {32'h45138a16, 32'hc35c1c84, 32'h432f2214},
  {32'hc4622102, 32'h42b2a989, 32'hc3c755ac},
  {32'h43ba4ff0, 32'h40b41ac6, 32'h429ebada},
  {32'hc4c537bb, 32'hc28d04d7, 32'hc0622dc0},
  {32'h4492e8b2, 32'h42199915, 32'h40cf8f0e},
  {32'hc4c34865, 32'hc3770499, 32'h42f4830d},
  {32'h44af0281, 32'hc3ff10d5, 32'h42db28f0},
  {32'hc4c2b51e, 32'h42917626, 32'h43939df0},
  {32'h44d1157c, 32'hc359d946, 32'h436a6155},
  {32'hc3bf9058, 32'hc2606368, 32'hc3a44da8},
  {32'h44be122d, 32'hc3505b68, 32'hc12aa303},
  {32'hc494eda1, 32'hc3921b7f, 32'hc31e98c4},
  {32'h43d05b78, 32'hc3dbc70a, 32'hc352e878},
  {32'hc4fad085, 32'h40446f45, 32'hc435b9b0},
  {32'h446c155a, 32'hc21dc5ec, 32'h43964a0e},
  {32'hc490632e, 32'hc2749c90, 32'hc3611a7c},
  {32'h44bf7c6f, 32'h415d1188, 32'hc34e4ddb},
  {32'hc4d8bf4c, 32'h4305397d, 32'h42aaf54f},
  {32'h43c125c8, 32'hc2e3622c, 32'hc23b10aa},
  {32'h43d232db, 32'hc323c466, 32'hc2b23722},
  {32'h438e4e46, 32'h42d9df10, 32'hc35fb5f0},
  {32'hc1010970, 32'hc323528f, 32'hbee54d12},
  {32'h4412353e, 32'h43152c7e, 32'h3ecfa1b4},
  {32'hc3fa84c8, 32'hc3536f3c, 32'hc295b508},
  {32'hc2877820, 32'hc391b9b7, 32'h42b3aae9},
  {32'hc4463c5c, 32'h41ccc2f1, 32'hc3b1b29c},
  {32'h44552fa0, 32'h437293f2, 32'h427367f4},
  {32'hc517e9de, 32'hc3be668f, 32'hc2112387},
  {32'h44e317d4, 32'h435dd374, 32'hc2ec8b24},
  {32'hc50734b5, 32'h42e8d6e3, 32'h40f332c1},
  {32'h44fb947d, 32'hc304f7d8, 32'hc37d2eec},
  {32'hc50929b0, 32'hc28a5dc3, 32'hc40981cc},
  {32'h450ba214, 32'h42b9c98c, 32'h43d314ad},
  {32'hc46db566, 32'hc3b3127f, 32'h4367773c},
  {32'h44e40719, 32'hc30f0c35, 32'h425dc29d},
  {32'h43349c60, 32'hc2f6d448, 32'hc308c1c2},
  {32'h450cb172, 32'h4373ea0d, 32'hc351de15},
  {32'hc4871de5, 32'h40d5dc1b, 32'h4310badf},
  {32'h438b48cd, 32'hc33dc62f, 32'hc32c647c},
  {32'hc502387c, 32'h43640fb2, 32'h4407ed99},
  {32'h443dfb4a, 32'hc3412db7, 32'hc2f0d394},
  {32'hc4c4416e, 32'hc40530ef, 32'hc30c2b34},
  {32'h44c18c78, 32'hc2bada6f, 32'h41fd04f5},
  {32'hc5158d50, 32'hc3ab6a86, 32'hc4108dc3},
  {32'h44f17d3d, 32'h43a7d194, 32'hc38ddbda},
  {32'hc430363f, 32'hc41e69f3, 32'h429dce95},
  {32'h4500dc1d, 32'h42a6e042, 32'hc2adcd23},
  {32'h43036550, 32'h4315eed6, 32'hc2a4268c},
  {32'h43081ea0, 32'h43cb925b, 32'hc1ff9ad0},
  {32'hc4ace502, 32'hc364f6d5, 32'hc31262f0},
  {32'h446e7959, 32'h426df83c, 32'h428c52c7},
  {32'hc40563ac, 32'hc19926de, 32'hc1b62f05},
  {32'h4452c886, 32'hc3ae6a34, 32'h434acb0c},
  {32'h43d5bea0, 32'hc399134f, 32'hc3654a51},
  {32'h442d20b0, 32'h41e0235f, 32'hc399399b},
  {32'h42a2aca8, 32'hc1bd35dc, 32'hc2a9f653},
  {32'h43ed47b8, 32'h4307d783, 32'h438392c2},
  {32'hc36f1080, 32'h42550a9c, 32'hc30cc788},
  {32'h44ea9558, 32'h428478c6, 32'hc39c5f93},
  {32'hc4f8c499, 32'hc2c23913, 32'hc3567a26},
  {32'h43c12ddb, 32'h439234e5, 32'h43c4d38d},
  {32'hc511b60d, 32'h43dddb62, 32'hc3bd96de},
  {32'h4466874c, 32'h43b8227e, 32'hc420ac5f},
  {32'hc47a6e02, 32'hc30b7eb1, 32'h439bd077},
  {32'h4506b4a0, 32'h43775f1e, 32'hc3a9226b},
  {32'hc480fb0f, 32'hc240222a, 32'h43808714},
  {32'h450a3bee, 32'h42622a76, 32'hc27da016},
  {32'hc483552d, 32'h435de17a, 32'h4315e2fa},
  {32'h44fa16b8, 32'hbedb4998, 32'hc32f3c5e},
  {32'hc480c642, 32'h4387a419, 32'hc3ecb8bd},
  {32'hc381c960, 32'h436aec2f, 32'hc380c551},
  {32'hc497f32e, 32'hc35b442b, 32'hc3422fb6},
  {32'h44d43f87, 32'hc3303272, 32'h41b11ff9},
  {32'hc5141e66, 32'h42592f68, 32'h4272134c},
  {32'h44cd222e, 32'hc324cfdb, 32'h43839a01},
  {32'hc38fac90, 32'h40f54b3f, 32'hc2966b5c},
  {32'h4317bc3c, 32'h4296e122, 32'hc262676c},
  {32'hc498c4cb, 32'h4386613d, 32'hc24613aa},
  {32'h44c0d376, 32'h42069959, 32'h4205f60d},
  {32'hc474f08c, 32'h4323a66f, 32'h43b995de},
  {32'h450e334c, 32'hc38a6fe5, 32'h4392299a},
  {32'hc395150c, 32'h43408538, 32'h422d1d9c},
  {32'h4505c7fe, 32'h43eca104, 32'h437c0903},
  {32'h42904ed9, 32'hc3929c2e, 32'hc195cdd6},
  {32'h4457531d, 32'h42ad6788, 32'hc2362e5d},
  {32'h43a0e532, 32'h437170d5, 32'hc236b2a2},
  {32'h42425ee0, 32'hc23cd2f0, 32'h424aff76},
  {32'hc508cf1a, 32'hc18bc2df, 32'hc255e101},
  {32'h4512daab, 32'hc1d3defb, 32'h42c69526},
  {32'hc36626c0, 32'h429841f8, 32'hc371b713},
  {32'h44dbcfdc, 32'hc3829ee2, 32'hc10ec129},
  {32'hc3d9fc06, 32'hc22d3dc7, 32'hc39e9075},
  {32'h442b7bf8, 32'hc28d0830, 32'hc31e7693},
  {32'hc4edc76a, 32'hc345f034, 32'h435eefb8},
  {32'h4289f748, 32'hc2ef0b62, 32'h4286f1ac},
  {32'hc475e178, 32'h4311d864, 32'h44109e5c},
  {32'h4430d317, 32'hc2d6f8d4, 32'hc3a59e05},
  {32'hc3b28774, 32'h42847870, 32'h43ef4984},
  {32'h438b54fc, 32'hc3267d82, 32'hc275f117},
  {32'hc401ecae, 32'hc32da0d0, 32'h439bf889},
  {32'h450cdf01, 32'hc399c894, 32'h4359064c},
  {32'hc3c0fabe, 32'h414e9b16, 32'hc385203e},
  {32'h43b6edb4, 32'h4385b608, 32'h41809306},
  {32'hc50fe808, 32'h42dc76c3, 32'h439521b3},
  {32'h442a1aa7, 32'hc3387a91, 32'hc37cdea8},
  {32'hc4d5e7a4, 32'h42f42096, 32'h4392850a},
  {32'h4522f3bd, 32'h429b0dee, 32'hc4175cc6},
  {32'hc41fe6fc, 32'hc31aa39b, 32'hc3059cca},
  {32'hc2584280, 32'hc40d2371, 32'h43d04289},
  {32'hc490b7aa, 32'hc26412ad, 32'hc29bd56b},
  {32'h44878a73, 32'hc3b134f9, 32'hc328117b},
  {32'hc4976e88, 32'hc3d2bbe8, 32'h435fdbfb},
  {32'h44b13f14, 32'h41057174, 32'h43bd2964},
  {32'hc508b79b, 32'hc2e8e3f9, 32'h4324ce50},
  {32'h44b1038c, 32'hc3926be7, 32'h4306a65e},
  {32'hc434b9ea, 32'h439af2d0, 32'h434b74f1},
  {32'h451533b2, 32'h4353ee07, 32'hc3dd3570},
  {32'hc4130b26, 32'h41cb5da2, 32'h430baf1a},
  {32'h44c51b06, 32'hc2b8c76e, 32'h43d9e90e},
  {32'hc3f8de2b, 32'hc337d125, 32'hc28ddd91},
  {32'h45000d82, 32'h43ad0c27, 32'hc300f60c},
  {32'hc4ba4270, 32'h43b7dce0, 32'h43883f1a},
  {32'h44c6e649, 32'h412a7c55, 32'hc3c5a210},
  {32'hc42d86e0, 32'hc39330a3, 32'hc321bfa3},
  {32'h43e36200, 32'h4306817b, 32'h431b5df2},
  {32'hc49a90f1, 32'hc2083fbe, 32'h4347f23c},
  {32'h44cb993b, 32'h434e00cf, 32'h43533c24},
  {32'hc4cad708, 32'hc3e12d03, 32'h439e21cc},
  {32'h42f06aba, 32'h431905a5, 32'hc3022fb0},
  {32'hc4f68273, 32'h428f990a, 32'h43b8b71a},
  {32'h44279e30, 32'hc250f7a8, 32'h42abf144},
  {32'hc3a9ea72, 32'hc08af46d, 32'h42dd6da9},
  {32'h44ed2956, 32'hc2ffbf43, 32'hc1d876b0},
  {32'hc35508e8, 32'hc2d12572, 32'hc3c1d15c},
  {32'h451b66a7, 32'h420d707e, 32'hc32a12c6},
  {32'hc4d679a4, 32'hc2110f93, 32'hc2169d55},
  {32'h450dc6a2, 32'h4300c431, 32'h42b26f76},
  {32'h422cf6f0, 32'h43564eba, 32'hc2e839a0},
  {32'h447d929b, 32'hc3a1e41f, 32'h4319f659},
  {32'hc3411dc0, 32'hc0e94524, 32'h42a5f503},
  {32'h4507b62a, 32'h43a3323a, 32'hc20549b9},
  {32'hc358e7e6, 32'hc38f7861, 32'hc38f6d1d},
  {32'h447cbe48, 32'hc31a26ec, 32'h435bd544},
  {32'hc4a6a2e8, 32'h42d4d77c, 32'h43c76338},
  {32'h4380bf34, 32'hc2bf6128, 32'h4376fdb4},
  {32'hc32cb1e7, 32'h4397d19d, 32'h42ede24b},
  {32'h44a29989, 32'h40c338ec, 32'hc28ead69},
  {32'hc4eb8712, 32'hc36b40ca, 32'h437899f5},
  {32'h44da2ea7, 32'hc33d8ca6, 32'hc35d085b},
  {32'hc4bc86f7, 32'h42907a74, 32'hc2c4433b},
  {32'h43933b54, 32'h436f0247, 32'hc140a5f6},
  {32'hc40c2ff3, 32'h43b36569, 32'hc12a2a5c},
  {32'h44778374, 32'hc38d2459, 32'h429411ed},
  {32'hc436d36d, 32'hc2ba95aa, 32'h432b56fc},
  {32'h44b02a32, 32'hc256e5d7, 32'hc3ce0b45},
  {32'hc3d6aae0, 32'h4286665a, 32'h4389a13f},
  {32'h44fdc4dc, 32'h4323c6fc, 32'h42d8ae02},
  {32'hc50dfde2, 32'hc350d899, 32'hc3704511},
  {32'h45078248, 32'h4153c158, 32'hc154abc5},
  {32'hc4eb24b1, 32'hc1eb558f, 32'h4302a4e2},
  {32'h4493d05c, 32'hc28d4683, 32'hc2086971},
  {32'hc4878ec0, 32'hc385a5e9, 32'hc3a9f5db},
  {32'h44e342de, 32'h4142a049, 32'hc3307bf2},
  {32'hc40c66fd, 32'h438cacc1, 32'h433c803f},
  {32'h44aa4c95, 32'hc326ad33, 32'h4345a6da},
  {32'hc43faa94, 32'hc3767ad6, 32'h41bde22a},
  {32'h44e34142, 32'hc22e5363, 32'h43ef2065},
  {32'hc5018e73, 32'h42cbab71, 32'h438000d7},
  {32'h4388f8a4, 32'h437791f8, 32'hc3103957},
  {32'hc41a7724, 32'h427faeda, 32'hc118eebe},
  {32'h43cbb72a, 32'hc1f49f11, 32'hc29c916c},
  {32'hc373738e, 32'h41a58208, 32'hc30d63df},
  {32'h45009f5c, 32'h43100383, 32'h43f0ac75},
  {32'hc30fe40a, 32'hc317ba4b, 32'hc29f93ba},
  {32'h438c5e6c, 32'hc2d9d320, 32'h419b2995},
  {32'h4367ecaa, 32'hbf134b14, 32'h435e447d},
  {32'h44db628a, 32'hc1989789, 32'h433bff6b},
  {32'hc446437c, 32'hc28717cd, 32'hc24d6cf1},
  {32'h445c197c, 32'h42b59785, 32'h43333284},
  {32'hc34c70ac, 32'hc2566bec, 32'h4327d576},
  {32'h44cffcd7, 32'hc39a2549, 32'h4302fb76},
  {32'hc50f36d4, 32'h4406b8d8, 32'h433205a2},
  {32'h45194669, 32'h4337763a, 32'h42dfba71},
  {32'hc4f65b2c, 32'h419f0cfe, 32'h43a312fa},
  {32'h44e4b418, 32'hc33f447e, 32'h42c34ca6},
  {32'hc4c6da72, 32'h42925129, 32'hc314fc8b},
  {32'h4482ab09, 32'h42c184ca, 32'h41178a93},
  {32'hc493fb07, 32'h43c18745, 32'h43844f36},
  {32'h44c9bd8f, 32'hc3007fa0, 32'h421258a2},
  {32'hc401614f, 32'h42a7227a, 32'hc3985726},
  {32'h4406c114, 32'hc2ff9e8f, 32'h4319ce22},
  {32'hc5079f34, 32'h40e0bf85, 32'hc3f1f1bd},
  {32'h450f3843, 32'h42f5c631, 32'hc3b93666},
  {32'hc41a9a93, 32'h43ae3189, 32'hc2963a39},
  {32'h44a57817, 32'h42aec0ba, 32'h4160d59c},
  {32'hc4421970, 32'hc2ac9c88, 32'hc34f1b66},
  {32'h4498ab4e, 32'h42e898c5, 32'h424e9f55},
  {32'hc4267744, 32'hc2da560b, 32'h438a988f},
  {32'h4515a677, 32'hc35e8ad9, 32'hc2883f90},
  {32'hc4a1719c, 32'hc3aca246, 32'h42f95146},
  {32'h44019482, 32'h434d1702, 32'h4380267e},
  {32'hc506295d, 32'hc3f1a690, 32'hc395a69e},
  {32'h44c11060, 32'h439524f1, 32'hc39cf782},
  {32'hc49ddb73, 32'h431ca294, 32'hc39647ab},
  {32'h441b430a, 32'h429e4f31, 32'hc245f8e4},
  {32'hc4c24124, 32'hc29f20d9, 32'h41abeffe},
  {32'h44f6ba0f, 32'hc2304cab, 32'h4390890e},
  {32'hc2a6f168, 32'h43918f9c, 32'hc2de53f2},
  {32'h44a7d382, 32'h437c63a4, 32'h43b4d3fd},
  {32'hc48aa111, 32'hc303982e, 32'h427542bd},
  {32'h44c0b908, 32'h429767ed, 32'hc30352c5},
  {32'hc49fb3e5, 32'hc074da46, 32'h401ca040},
  {32'h44a0d844, 32'hc268886c, 32'hc353d912},
  {32'hc4fd4031, 32'hc293edd1, 32'hc31e1c80},
  {32'h448beb1e, 32'hc31777ec, 32'h432a8577},
  {32'hc3e72078, 32'hc1c81221, 32'hc20735a8},
  {32'h449b5e04, 32'h433ec8c2, 32'h42811ee2},
  {32'hc3fcd140, 32'hc2853d80, 32'h4175fb6a},
  {32'h45016d56, 32'hc3821c5d, 32'hc3697d12},
  {32'hc50cf336, 32'h430a784d, 32'hc3737813},
  {32'h44f2c4f6, 32'h436cb81a, 32'h436ee7ad},
  {32'hc47e3174, 32'hc2eea1dc, 32'h43872963},
  {32'h4455e7b4, 32'h42c8ef5e, 32'hc3fee9b8},
  {32'hc4bf8d52, 32'hc21c66f4, 32'h43639330},
  {32'hc372fd31, 32'hc3316391, 32'h437530e0},
  {32'h433ebf00, 32'h431ea874, 32'hc30ba936},
  {32'h448236ed, 32'hc1c75f9d, 32'hc1aac608},
  {32'hc43a67fc, 32'h42f43b17, 32'hc2b537bd},
  {32'h4468de62, 32'h4396debf, 32'hc3327b63},
  {32'hc2ba6348, 32'h40bad004, 32'h4304470d},
  {32'h44015b12, 32'h42f8f53e, 32'hc2b4aa52},
  {32'hc50c7e36, 32'h42376952, 32'hc2a92f96},
  {32'h44c57e35, 32'h43dd1363, 32'h41d9ddd0},
  {32'hc2aa0240, 32'hc38236ce, 32'h428f7f79},
  {32'h43d94f63, 32'hc3b63638, 32'h432b344f},
  {32'hc4f69b7c, 32'hc2ca2265, 32'hc3083bb3},
  {32'h448c9fa0, 32'h42796778, 32'h434b1374},
  {32'hc4b23648, 32'hc3abea81, 32'hc34d5610},
  {32'h44c87184, 32'h42f1878b, 32'hc2704c0a},
  {32'hc490cf3a, 32'h43104372, 32'h40c95dbe},
  {32'h442cd2aa, 32'h435a6bc6, 32'h43821be9},
  {32'hc458f21a, 32'hc3947aaf, 32'h43b0fef4},
  {32'h44b711ba, 32'h4370f0b8, 32'h42794fc6},
  {32'hc4c36f18, 32'hc3c083d8, 32'h435f388f},
  {32'h444281ad, 32'hc35462ee, 32'h4346073c},
  {32'hc4d0f801, 32'h43e858cb, 32'hc28ba652},
  {32'h44ea9559, 32'h43428d62, 32'h426bb043},
  {32'hc4eeb4ff, 32'h43c2ff6c, 32'hc2a2c023},
  {32'h444b5ae6, 32'h42b1865a, 32'hc3444505},
  {32'hc4262eb3, 32'hc3250204, 32'h432ce4c0},
  {32'h451c2c5e, 32'h43f0cb5a, 32'h42ae6690},
  {32'hc5161687, 32'h42ff23df, 32'hc2c52939},
  {32'h440f3e34, 32'h438f306b, 32'h431486f7},
  {32'hc499d4f2, 32'h43987817, 32'hc3a57dba},
  {32'h447e800a, 32'h417d43ac, 32'h42858293},
  {32'hc47c0cb6, 32'hc3647054, 32'hc3b1824c},
  {32'h44d671a0, 32'h43ca4185, 32'hc31893f3},
  {32'hc518b799, 32'hc20f2942, 32'hc3c919dd},
  {32'h44e0762e, 32'hc3ae006f, 32'h4326219a},
  {32'hc50659ca, 32'h435f845f, 32'hc2d716e2},
  {32'h448bf6e4, 32'h430eb34f, 32'h413dc94d},
  {32'hc424fb13, 32'hc34012c9, 32'h43df8e66},
  {32'h44b36b6a, 32'hc2a216b0, 32'h427b7761},
  {32'hc4dd0a22, 32'h436fc68a, 32'h418f9e6d},
  {32'h448d38ea, 32'h428a5566, 32'h42abe5b7},
  {32'hc4a90114, 32'hc2167710, 32'h4047ba4a},
  {32'h448be48f, 32'hc2d589a1, 32'hc1c851f5},
  {32'hc400f390, 32'h43186dad, 32'hc38a3db7},
  {32'h44dea9a2, 32'h426a985f, 32'h4323e760},
  {32'hc4adda4d, 32'hc20f9ff4, 32'h430c07bb},
  {32'h44fb889b, 32'hc3575af4, 32'hc31373b6},
  {32'h4266a304, 32'h4337096d, 32'hc38a1649},
  {32'h44820361, 32'hc2074c24, 32'hc370cb73},
  {32'hc4d575c2, 32'hc328e803, 32'h432cf8c3},
  {32'h4506586d, 32'hc35e5196, 32'h43b5b068},
  {32'hc4f9e3ac, 32'h431cf9c7, 32'h410bd12c},
  {32'h441f6414, 32'hc2251652, 32'hc33d55e7},
  {32'hc4d13233, 32'h43611087, 32'hc3d85b15},
  {32'h4395114c, 32'h412048f2, 32'h436c5d67},
  {32'hc4aae6ab, 32'h436c7cde, 32'h40ed613d},
  {32'h451c837b, 32'h42429b26, 32'h43841162},
  {32'hc4c52289, 32'hc35e415a, 32'hc3f971e7},
  {32'h451180a6, 32'h4388dfc0, 32'hc335026e},
  {32'hc45db2be, 32'hc3a45694, 32'hc28cf905},
  {32'h451a1775, 32'h43912da3, 32'h43fc398d},
  {32'hc51b2f49, 32'h425b0d84, 32'h42572b44},
  {32'h43f86174, 32'hc09f613e, 32'hc30e0b8a},
  {32'hc3f679f0, 32'hc202feb6, 32'hc39914c3},
  {32'h440b11b6, 32'hc41608df, 32'hc31fc38f},
  {32'hc4e3b702, 32'hc3423152, 32'h42a5c301},
  {32'h4505dc6c, 32'h4281ce5e, 32'h4389fcef},
  {32'hc4f933a2, 32'h4296e7ce, 32'h43002e3b},
  {32'h447c034e, 32'hc125575a, 32'hc31ee8a1},
  {32'hc500bf4e, 32'hc2d127a1, 32'hc3372080},
  {32'h44c604c4, 32'h42b9204c, 32'h435c63e7},
  {32'hc405eca1, 32'hc39bbd09, 32'h420b73d9},
  {32'h44809d47, 32'hc2551f00, 32'h43ab209d},
  {32'hc4cea14b, 32'h4104ef51, 32'hc3d92f88},
  {32'h44911d9f, 32'hc226fcc4, 32'h433bfb80},
  {32'hc4521b9a, 32'h430a3de8, 32'h42839772},
  {32'h4503d419, 32'h4287cccc, 32'h4295aefc},
  {32'hc3b08b34, 32'hc2861fe2, 32'h43570e8c},
  {32'h4500d38a, 32'hc3387854, 32'hc4559730},
  {32'hc50d9081, 32'h4388e614, 32'h42ce9814},
  {32'h44b5dd9e, 32'h438bccef, 32'h43b28e74},
  {32'hc50f8311, 32'hc326aca9, 32'h42c6960e},
  {32'h4511a797, 32'hc2a5e651, 32'hc10b89e6},
  {32'hc4943718, 32'hc40dd6b9, 32'hbf7b7020},
  {32'h4416c473, 32'hc3656484, 32'hc27f2b0f},
  {32'hc516d348, 32'hc18e2b2e, 32'h4405288f},
  {32'h448770ec, 32'h43a8c9ff, 32'h434c8c48},
  {32'hc5133bec, 32'h4172084d, 32'hc3238a20},
  {32'h44e44d51, 32'hc2ae981a, 32'hc3a13856},
  {32'hc4ff04e5, 32'h439b8274, 32'h4256ac08},
  {32'h44554e72, 32'h43b12c89, 32'h4298ebcd},
  {32'hc272e48f, 32'h426ca7c4, 32'hc2f09f0f},
  {32'h4314bc78, 32'hc3d43c28, 32'h42f2cbec},
  {32'hc4ce953a, 32'h437827be, 32'h426fbe29},
  {32'h442668be, 32'hc19d7607, 32'hc3495b10},
  {32'hc482ae04, 32'hc311495c, 32'h429713d5},
  {32'h444ce295, 32'h44131834, 32'h42e0da89},
  {32'hc4e46c9b, 32'hbfce885c, 32'h4144c650},
  {32'h40c2a0f8, 32'hc34998e6, 32'h42ca7e61},
  {32'hc399a750, 32'h42c97950, 32'hc1a587d0},
  {32'h42075308, 32'hc3b19319, 32'h4327ea58},
  {32'hc3cb9796, 32'h43692db2, 32'hc323d7c3},
  {32'h41e7d740, 32'h42888941, 32'hc28bbe0d},
  {32'hc4a3503b, 32'hc2c9a2c8, 32'h438b5f52},
  {32'h4462fd35, 32'h43eac954, 32'h43567233},
  {32'hc4ab2014, 32'h432d7498, 32'h3fcc173b},
  {32'h4412904c, 32'hc363d9e7, 32'hc3170e44},
  {32'hc40d4715, 32'hc2758efe, 32'h42b27a85},
  {32'h450d9120, 32'h431f0d28, 32'hc2b42b88},
  {32'hc4da32ab, 32'h4281b5d1, 32'hc3f64282},
  {32'h446ecf20, 32'hc355f73e, 32'hc20409e2},
  {32'hc4f6ea9c, 32'h4369085e, 32'hc2f3597b},
  {32'h4502e584, 32'h41494c38, 32'h43d06df5},
  {32'hc49ecd16, 32'h43830d41, 32'h41a31bc5},
  {32'h44e90aa0, 32'hc305b36c, 32'hc294ee48},
  {32'hc4a27784, 32'h43008da0, 32'h4201a5f0},
  {32'h439f1248, 32'h42bba4cc, 32'h4307ea88},
  {32'hc41d80b2, 32'hc3a708c0, 32'hc2c918a2},
  {32'h43a72f70, 32'h43de207f, 32'hc3b06542},
  {32'hc4fe2aa3, 32'h420af3b3, 32'h4233f90a},
  {32'h44eb8193, 32'h433aa1d8, 32'h43f04ab6},
  {32'hc3b6f1e0, 32'h40206e10, 32'hc3c071d1},
  {32'h4464cd51, 32'hc257a0d5, 32'h432f3a6a},
  {32'hc4f8f117, 32'hc312ee31, 32'hc1b02fd0},
  {32'h448691a5, 32'hc1f60eae, 32'hc284d450},
  {32'hc5187a4c, 32'h432b2758, 32'h43e01598},
  {32'h44c00b61, 32'hc306a9a2, 32'h43d2a65b},
  {32'hc4c32538, 32'h42adfd9f, 32'h435346a2},
  {32'h450d13b3, 32'h42ac26b2, 32'h41198da4},
  {32'hc4186b18, 32'h4194467c, 32'hc29d5f69},
  {32'h44dd43cf, 32'hc20760a6, 32'hc30a4223},
  {32'hc501c722, 32'h41f469d4, 32'h441491b3},
  {32'h4478a21a, 32'h3f252d70, 32'hc2a03f00},
  {32'hc44502e6, 32'h41472ac8, 32'h42e225ad},
  {32'h4504f5ba, 32'hc3700440, 32'h43311900},
  {32'hc50ab076, 32'h439887c9, 32'h4292468b},
  {32'h44b1b03e, 32'h4394f3e4, 32'h43a6bf94},
  {32'hc4beeab6, 32'hc3c67727, 32'hc3da2c66},
  {32'h44d9463e, 32'hc274e5db, 32'hc3887ab3},
  {32'hc4848c96, 32'hc411276c, 32'hc3ebb90b},
  {32'h4517bdac, 32'h42269fd8, 32'h42ce077f},
  {32'hc5053fc1, 32'hc0689f98, 32'h43a7fd5e},
  {32'h4509cb1c, 32'hc31600f8, 32'h436b29e7},
  {32'hc4e15943, 32'hc2e3af11, 32'hc1ce7b7b},
  {32'h43d021e2, 32'hc399038e, 32'h4254e235},
  {32'hc5077c76, 32'hc3a624fd, 32'h43683718},
  {32'h44bb58f7, 32'h417eff0f, 32'hc42d0050},
  {32'hc3dce820, 32'h43bf272a, 32'h434d498b},
  {32'h44a8e3eb, 32'h4341e818, 32'h438c8b7e},
  {32'hc4a13b50, 32'h42df2ab5, 32'hc2b80fa9},
  {32'h450a0a44, 32'h42fc5916, 32'h435663a3},
  {32'hc4198bf6, 32'h43e74c13, 32'h434497f4},
  {32'h43dc00c0, 32'h42d1e29f, 32'h4322849d},
  {32'hc42c906a, 32'h41205ff7, 32'hc2ffb162},
  {32'h44983c7c, 32'hc26bf85a, 32'hc2d2776f},
  {32'hc413b0ec, 32'hc38e8944, 32'hc2d28acc},
  {32'h4398e69c, 32'h43e47ed0, 32'hc3618f2a},
  {32'hc49ce161, 32'h418a69bb, 32'h42a1ed87},
  {32'h4501b59e, 32'h438eb041, 32'h423670e0},
  {32'hc39ca8a5, 32'hc1f882a2, 32'h43977056},
  {32'h432ad718, 32'h43301a13, 32'h43cb142b},
  {32'hc2d7ec4d, 32'h435f6dd7, 32'hc1ee8fb8},
  {32'h44e96ff4, 32'hc369c596, 32'h40437af5},
  {32'hc4980e78, 32'h43e7a7aa, 32'h42ce0e6c},
  {32'h433c43be, 32'h43513596, 32'hc33b0f30},
  {32'hc35ab349, 32'h428bdf4d, 32'h43d390b6},
  {32'h440a6651, 32'hc2379a5a, 32'hc3ee94ca},
  {32'hc3f39578, 32'h4303aeb2, 32'hc1642f0c},
  {32'h44dd06be, 32'hc24f58d0, 32'h42b26610},
  {32'hc3d533a4, 32'hc328b305, 32'hc2fc1536},
  {32'h4505690b, 32'h4371b203, 32'hc3a93783},
  {32'hc3e5c1d0, 32'hbbda4000, 32'hc3297309},
  {32'h445bd3ce, 32'h41e1c818, 32'h406543a8},
  {32'h43aa1869, 32'h43a76653, 32'hc2af345d},
  {32'h452164cb, 32'h4365479b, 32'hc37bf0c9},
  {32'hc500f5db, 32'h42332a87, 32'h439203fd},
  {32'h4504d52a, 32'hc2bfc212, 32'hc38792b9},
  {32'hc467964e, 32'h42d42907, 32'h42985aab},
  {32'h43485b28, 32'h41023f09, 32'h43175f28},
  {32'hc31315c0, 32'hc3179000, 32'hc31c7e9e},
  {32'h43079894, 32'hc393ec8b, 32'hc404a50a},
  {32'hc3e5be10, 32'h42a5d62a, 32'h410c575f},
  {32'h43b80c59, 32'h42cc6076, 32'hc32a0605},
  {32'hc4e86cd6, 32'h418e865f, 32'hc337f471},
  {32'h44d72dcb, 32'hc3406bcd, 32'hc2895433},
  {32'hc4db56a9, 32'h42c1cd96, 32'h435bfadd},
  {32'h43e96cc8, 32'hc3fc0815, 32'hc420cbd6},
  {32'hc510bbac, 32'h435018be, 32'hc350c9ab},
  {32'h43f17cf0, 32'hc3479990, 32'hc399e976},
  {32'h44cd219c, 32'h41402731, 32'hc2831775},
  {32'hc43cf6eb, 32'h412af552, 32'hc28799ae},
  {32'h44397cfa, 32'hc390ce8a, 32'hc372892d},
  {32'hc4b82218, 32'h434171c2, 32'h428e6cf3},
  {32'h44eb7d89, 32'h4219b5a8, 32'h43067c5c},
  {32'hc40b5d14, 32'hc35a74f3, 32'h43b4c5e6},
  {32'h44922d2b, 32'hc296f666, 32'h42f1d5c1},
  {32'hc4e67fc8, 32'h43a0217b, 32'hc416153b},
  {32'h44aac00c, 32'hc2bf3e52, 32'hc2fb5baf},
  {32'hc417fedc, 32'h4388768a, 32'hc3ae6f34},
  {32'h43349470, 32'hc31071f9, 32'hc3429171},
  {32'hc4d662c8, 32'hc218440f, 32'h43a8011a},
  {32'h44e4ebf8, 32'hc3e3d6d0, 32'hc34f6884},
  {32'hc49ddc1c, 32'hc3201472, 32'hc2d9de9f},
  {32'h440f67a2, 32'h41d6f769, 32'h425969cc},
  {32'hc4fac3c2, 32'h438eab4f, 32'h436f7fe7},
  {32'h44630d42, 32'hc1e33915, 32'hc3ba916a},
  {32'hc4c5b796, 32'h44086f58, 32'h4334256e},
  {32'h440cc042, 32'h43739a87, 32'hc30d88c9},
  {32'hc4123599, 32'h43371546, 32'hc21042e7},
  {32'h433b4400, 32'hc31059f5, 32'hc3e64bdc},
  {32'hc5191828, 32'h4392c097, 32'hc3670c36},
  {32'h44c654a1, 32'h433352f9, 32'hc1fb1a41},
  {32'hc506646e, 32'hc2dad878, 32'hc1e56c8c},
  {32'h44b5f7fd, 32'hc35ac006, 32'hc276ef0c},
  {32'hc2a09100, 32'hc33d8450, 32'hc29fd33f},
  {32'h44d45604, 32'h430066ce, 32'h430223dd},
  {32'hc4c8707e, 32'h42f9c4ee, 32'hc4093580},
  {32'h44df094b, 32'hc323baa0, 32'h43234c35},
  {32'hc3ca0178, 32'hc2e9093a, 32'hc30552a9},
  {32'h436129b8, 32'h42335b96, 32'hc3ab5097},
  {32'hc439ee0d, 32'hc33f6828, 32'h423a410a},
  {32'h44eb8dc9, 32'hc2ef1061, 32'h42d08985},
  {32'hc50d1760, 32'hc3d39df7, 32'hc253c4d3},
  {32'h4510e9f0, 32'h4355b0c0, 32'hc2db8ee1},
  {32'hc4b23147, 32'h430e1e80, 32'h4338b641},
  {32'h450e82bb, 32'h4337c2a6, 32'h42be00f0},
  {32'hc3d48d2a, 32'hc141f8e8, 32'hc31dde7d},
  {32'h445b9c8c, 32'hc3462f90, 32'h430bf75f},
  {32'hc3fa749e, 32'h4357e029, 32'hc3722ef1},
  {32'h3f846780, 32'h414acc6b, 32'h428183f8},
  {32'hc4aceddd, 32'h42f02a2d, 32'h4386412b},
  {32'h4440cdff, 32'h42a87a33, 32'h4399e3f6},
  {32'hc502a42c, 32'h4335e6ed, 32'h42bcccd0},
  {32'h45032169, 32'hc28cc631, 32'h4332f9a1},
  {32'hc4f73217, 32'h43abc4ef, 32'h4384c5ea},
  {32'h451546e1, 32'h42e37a64, 32'h440392ca},
  {32'hc432bcf8, 32'h439d136f, 32'h41b8e278},
  {32'h43c14bc8, 32'hc2406fb3, 32'hc3296d5a},
  {32'hc505898d, 32'h43151075, 32'h431dcab0},
  {32'h44f8e29e, 32'h42a7a84b, 32'h43c2b19e},
  {32'hc4cffc63, 32'hc34ac260, 32'hc27ab013},
  {32'h44fd30a6, 32'h420a3a44, 32'h438ac0b6},
  {32'hc4ad18e5, 32'hc33193db, 32'h43210635},
  {32'h44149bfa, 32'h43528f49, 32'h4259cc72},
  {32'hc3ad02e0, 32'hc3492f0c, 32'hc3686fca},
  {32'h4495ec6f, 32'hc352a80b, 32'hc345567c},
  {32'hc50a4ff8, 32'hc360df7d, 32'hc3a34eec},
  {32'h451f4b29, 32'hc10cbd5a, 32'hc2bb930e},
  {32'h4137bd80, 32'hc3133ee3, 32'hc30a2a23},
  {32'h44d93af8, 32'hc1af1afb, 32'h43313325},
  {32'hc4e64b6f, 32'h43d34857, 32'h42927c44},
  {32'h450c4ac2, 32'hc2fefa22, 32'hc3a9ea81},
  {32'hc492628e, 32'h41007e3c, 32'h430b194d},
  {32'h447ef38d, 32'h421409c0, 32'h43ab9cb2},
  {32'hc4261f22, 32'hc29a409a, 32'h41d6767d},
  {32'h4460ecb0, 32'h44065d48, 32'hc3c2960e},
  {32'hc4e2a87a, 32'hc386c084, 32'hc3b0e1f5},
  {32'h43f98285, 32'h4376296f, 32'h42cee622},
  {32'hc4d109f5, 32'hc2f78b92, 32'h430bdbe8},
  {32'h4441fd6c, 32'h430af6b6, 32'h435205ef},
  {32'hc483b2f6, 32'hc1a50849, 32'hc1c561a9},
  {32'h449ec812, 32'h427f3f75, 32'h4316a742},
  {32'hc484ca16, 32'hc322addd, 32'h4392e22f},
  {32'h43d2abcc, 32'hc30e5764, 32'hc3a80ab9},
  {32'hc41a93f2, 32'hc337374a, 32'h44009d5d},
  {32'h44c8f6aa, 32'hc3ae6f4f, 32'h4365b765},
  {32'hc4f9dbb7, 32'h4280f0f2, 32'hc40b2521},
  {32'h44c86c21, 32'hc388bb5a, 32'h42e2183c},
  {32'hc5096c79, 32'hc323cbca, 32'hc23b67f9},
  {32'h44e23953, 32'hc3c77b9d, 32'h4328a84e},
  {32'hc4af0dee, 32'hc31f6aec, 32'hc0ea5178},
  {32'h44fc0af7, 32'h42c8b3fd, 32'h428850b6},
  {32'hc4b5d960, 32'h421b006c, 32'h425961f5},
  {32'h44d46bc2, 32'h42c1e322, 32'h43557d09},
  {32'hc3528082, 32'h42f71f7b, 32'h43269f94},
  {32'h451aa8c4, 32'h4286f2d6, 32'hc314b1eb},
  {32'hc50be60a, 32'hc3827707, 32'h43d47a09},
  {32'h44981c15, 32'hc39d3305, 32'hc2dafeae},
  {32'hc4591924, 32'hc38f24a6, 32'h43861586},
  {32'h44d5e4a6, 32'h4270cbe4, 32'h429c1b3b},
  {32'hc4fd352a, 32'hc397b935, 32'h4344f8d3},
  {32'h44785961, 32'hc3197d01, 32'h43b5e557},
  {32'hc4e8e9a6, 32'hc29d5a19, 32'hc3b631fe},
  {32'h450e38d5, 32'hc2996b74, 32'h435d68eb},
  {32'hc3909f13, 32'hc2a69102, 32'hc2ce2c5e},
  {32'h438e93ca, 32'hc3af6418, 32'hc3ba14bb},
  {32'hc42b385b, 32'hc2a6c5db, 32'hc2bd4064},
  {32'h4502c9c7, 32'h42a56387, 32'hc3b45e79},
  {32'hc2fdeb90, 32'hc2ad2df3, 32'h43188587},
  {32'h44f0e0c5, 32'h43f8e35e, 32'h43681795},
  {32'hc32eb8b0, 32'h4350e887, 32'h434afc3e},
  {32'h444572f6, 32'h431755a7, 32'h43817b3c},
  {32'hc4048ad7, 32'h41948786, 32'h4356058b},
  {32'h44cea130, 32'hc3d628bb, 32'h439f0c30},
  {32'hc4db3d7c, 32'hc38a4c94, 32'hc32835f6},
  {32'h43d15a10, 32'h42db3655, 32'h418c27bd},
  {32'hc43bbd48, 32'h40cabad0, 32'h437e0132},
  {32'h441007e4, 32'h42d6ac93, 32'h434ff347},
  {32'hc49524b1, 32'h42b2cc99, 32'h41a3a2f5},
  {32'h44d120f1, 32'hc2d8cc28, 32'hc3b803c7},
  {32'hc4897595, 32'h41cfb040, 32'h4203ff04},
  {32'h4508c3f9, 32'hc21c8a57, 32'hc2e3f806},
  {32'hc413ca0a, 32'h434a0b67, 32'h4387e24a},
  {32'h44c96a9e, 32'h413b55f0, 32'h43b2cd07},
  {32'hc43ba03c, 32'hc31e6bf9, 32'hc2ddd47e},
  {32'h448481eb, 32'h438650a5, 32'hc3507ae6},
  {32'hc4b71e33, 32'hc3a47f4d, 32'h43bb1046},
  {32'h44c51e02, 32'h43c366fc, 32'hc2a4845c},
  {32'hc4b141cc, 32'hc35f0ade, 32'h433c9edc},
  {32'h4517b2b3, 32'h4317bdcf, 32'h4311f362},
  {32'hc4d9f163, 32'h43e858ba, 32'h439056ae},
  {32'h44c49ab4, 32'hc2f4f9c2, 32'h439dccd8},
  {32'hc4dfd9b1, 32'h43108bde, 32'hc2badf2f},
  {32'h44bc3356, 32'hc35bc254, 32'hc2bfe07a},
  {32'hc5101e92, 32'hc28fe7ba, 32'hc2876ffa},
  {32'h43e1f6c0, 32'h43e6597c, 32'h4352d02e},
  {32'h43b7c4a8, 32'h42db290c, 32'hc322ace3},
  {32'h450977b0, 32'hc3932201, 32'hc1e4c4a4},
  {32'hc2b04af2, 32'hc29dae5d, 32'h43ed0be2},
  {32'h44fa7310, 32'hc21d5f5c, 32'hc2873e69},
  {32'hc41760eb, 32'h42c136f0, 32'h43145d46},
  {32'h450c789e, 32'hc20fa4e1, 32'hc37128cc},
  {32'hc492326a, 32'hc2a29fa4, 32'hc3855526},
  {32'h445705a4, 32'hc2be39c8, 32'hc317101f},
  {32'hc49a83b2, 32'hc2d26d18, 32'h42dbd908},
  {32'h4505a5ef, 32'hc3c0add3, 32'h432e12ed},
  {32'hc4246a36, 32'hc3e41cb0, 32'hc2f15981},
  {32'h43c0d1dc, 32'hc30c946c, 32'h43809d14},
  {32'hc3c32964, 32'h43b2d3e6, 32'hc048e748},
  {32'h450c028c, 32'hc1ad8148, 32'h43b14177},
  {32'hc4b9b1b2, 32'h430da5e2, 32'hc2075b68},
  {32'h42720ab0, 32'hc3aa12e5, 32'h432e9551},
  {32'hc5126548, 32'h421c5f98, 32'hc28198a3},
  {32'h4485491a, 32'hc29d49b6, 32'h436338f8},
  {32'hc46c0783, 32'h42811b4a, 32'hc285b820},
  {32'h4422056c, 32'h439315ee, 32'h41a95ee7},
  {32'hc4fab578, 32'hc11ae660, 32'h435d5d3d},
  {32'h440be7aa, 32'h437e516b, 32'h43390ec4},
  {32'hc42b5587, 32'hc1135697, 32'h43810d19},
  {32'h4388e0b2, 32'hc2d10618, 32'h436e447b},
  {32'hc43a398c, 32'hc3b7ad82, 32'hc3ce2dab},
  {32'h4517f33b, 32'hc39b7cb7, 32'h425d2524},
  {32'hc2f57b80, 32'hc375d526, 32'h42377260},
  {32'h44576e54, 32'hc214795e, 32'hc1ffe0c7},
  {32'hc3ec605b, 32'h43968d64, 32'h42803e4b},
  {32'h44821522, 32'h42291d0d, 32'h4315ad04},
  {32'hc4bcb730, 32'h441391e9, 32'h43031447},
  {32'h448e07bc, 32'hc1c0d7cc, 32'hc166f80b},
  {32'hc4aa8f6e, 32'h411ee4f0, 32'h435d5de9},
  {32'h451688b7, 32'h4281b64a, 32'hc37a9e04},
  {32'hc505c170, 32'hc2e9a67f, 32'hc2edf53f},
  {32'h44eaa222, 32'h42d00e57, 32'hc1daa548},
  {32'hc4f15e88, 32'h42b6a80b, 32'h4273f422},
  {32'h45169d00, 32'h4187cd8d, 32'hc3f6c736},
  {32'hc438d264, 32'h43031edf, 32'hc28b215d},
  {32'h451033dd, 32'hc32d2864, 32'hc36333c6},
  {32'hc4e8377a, 32'h4102df84, 32'hc397ad2d},
  {32'h446dc0f4, 32'h434d895e, 32'hc2d6a850},
  {32'hc4302932, 32'h41aa5524, 32'hc2542e36},
  {32'h43c7c911, 32'hc269f415, 32'h43cb01c7},
  {32'hc4f11fa0, 32'h43d703de, 32'h42cc2725},
  {32'h4279a690, 32'h3fea45a5, 32'h42562ea4},
  {32'hc3796b04, 32'hc2fc174f, 32'h41ccd7ce},
  {32'h44100878, 32'h40919f4d, 32'h433ab7eb},
  {32'hc4ee51f5, 32'h42e58952, 32'h43bf6027},
  {32'h44a2f8d1, 32'hc292e1ef, 32'hc35bf590},
  {32'hc44acecf, 32'hc424de0d, 32'hc34d71fb},
  {32'h44ac6393, 32'hc3b86c0e, 32'h428fcbe0},
  {32'hc4eef730, 32'h4311ce19, 32'hc30acc34},
  {32'h44726866, 32'hc2cf3e74, 32'h43eca8a7},
  {32'hc511a28e, 32'h40cf5b1d, 32'h43137973},
  {32'h43b93c44, 32'h42dfd6fa, 32'hc2e8b5c9},
  {32'hc444e8e6, 32'hc3e613da, 32'h42375407},
  {32'h450ca574, 32'hc33660af, 32'h4392d758},
  {32'hc4eb94a7, 32'hc1e368b5, 32'h43238fca},
  {32'h41f32720, 32'hc35e5796, 32'hc2cc6800},
  {32'hc4a6702c, 32'hc23bd272, 32'h41735272},
  {32'h45095b92, 32'hc30107bb, 32'hc390209e},
  {32'h4325c9a8, 32'h42c75674, 32'h42c9fd64},
  {32'h4334171c, 32'hc395cdbb, 32'h435ce271},
  {32'hc49391ac, 32'h43cc92ae, 32'h437b26ed},
  {32'h44c63da1, 32'hc3a1f229, 32'hc3220db9},
  {32'hc3b777f8, 32'h432b46d4, 32'h425b8c6c},
  {32'h4518caa0, 32'hc1d86c58, 32'h4379720c},
  {32'hc4b07f8a, 32'hc2abb346, 32'hc2aa36a2},
  {32'h44f90eea, 32'h433c51a4, 32'h4373ce9e},
  {32'hc4e99200, 32'hc2608337, 32'h42ee60c2},
  {32'h420781e0, 32'hc36a2678, 32'h420b1d5d},
  {32'hc4d8607f, 32'hc38a3c2b, 32'hc0eb723a},
  {32'h451956c1, 32'h436737c1, 32'h41b81caf},
  {32'hc4eaa3b1, 32'h42f1e7f8, 32'hc3206b3f},
  {32'h446aae3e, 32'h3faf9375, 32'hc29c7877},
  {32'hc3eda73c, 32'hc3673302, 32'h433e4b3c},
  {32'h450d8032, 32'hc3e5786e, 32'h41305664},
  {32'hc5043dd9, 32'h438ae966, 32'h41c5f091},
  {32'h44320733, 32'hc2f5cad4, 32'h4335ce83},
  {32'hc34296b8, 32'h43729f04, 32'hc3cef9b8},
  {32'h45024519, 32'hc3478280, 32'h432b5a56},
  {32'hc4c06c10, 32'h42a1c373, 32'hc2e15f85},
  {32'h44c662d9, 32'hc326fbb0, 32'h4320baf6},
  {32'hc47f4466, 32'hc3db9f42, 32'h43201174},
  {32'h44b74d21, 32'hc095e661, 32'hc30cee8d},
  {32'hc4793016, 32'h42aa6634, 32'h43289ac9},
  {32'h446335c5, 32'h4391fea7, 32'h43098972},
  {32'hc4193dd0, 32'hc23d22ff, 32'hc2fb4b85},
  {32'h450432cb, 32'hc30cbccf, 32'hc36c9466},
  {32'hc3c7ae6c, 32'hc319dba7, 32'h4311b932},
  {32'h44f8127e, 32'h43a81882, 32'hc2f7f5b3},
  {32'hc4191e89, 32'hc3c3acc2, 32'h43899d08},
  {32'h4468427a, 32'h42d41c03, 32'h43980ea0},
  {32'hc4b2c498, 32'h43453a72, 32'h42dc3a33},
  {32'h44ccae91, 32'hc38e5f4f, 32'hc2609d39},
  {32'hc47f845c, 32'hc2a51561, 32'hc31e237f},
  {32'h43e0e560, 32'h436c57fa, 32'h4352a45a},
  {32'hc4607d72, 32'h4194d560, 32'hc311d942},
  {32'h43629c4e, 32'h43bc3e94, 32'h4389aa7f},
  {32'hc4aa5afe, 32'hc28b741f, 32'h419fa470},
  {32'h441aeb0c, 32'hc180656a, 32'h41b120e0},
  {32'hc4bd1114, 32'h4241339b, 32'hc2ee9afe},
  {32'h449eec8e, 32'h433d1314, 32'hc361854b},
  {32'h42af5a00, 32'h42862bdf, 32'hc2305726},
  {32'h443ae6b8, 32'hc2b3121d, 32'h430f8099},
  {32'hc44a729e, 32'hc311965c, 32'h42b38716},
  {32'h44d15c62, 32'hc300a4fa, 32'hc269741c},
  {32'hc507997c, 32'hc39dfb97, 32'h429eb9a8},
  {32'hc2274fc0, 32'h4398de8e, 32'hc2b81757},
  {32'hc460d596, 32'h430811b7, 32'h4283b5f8},
  {32'h441b106e, 32'hc343f7e1, 32'h426ed1ca},
  {32'hc433c535, 32'hc3c7bdcd, 32'hc369e75d},
  {32'h4418b276, 32'h42480a54, 32'hc214ec3e},
  {32'hc4b29c6d, 32'h421bd058, 32'hc35656b6},
  {32'h44d7fc47, 32'hc3090663, 32'h43b8db91},
  {32'hc4749ded, 32'h41b5cd47, 32'h424234bd},
  {32'h44059e34, 32'h41e4bd2e, 32'hc268ad19},
  {32'hc47a11c8, 32'h43055fd6, 32'hc2ac8d9a},
  {32'h44ddca06, 32'hc3648cbc, 32'h43c0afb8},
  {32'hc3096cd8, 32'h43aa6104, 32'h43026907},
  {32'h4485e128, 32'h439bacd6, 32'h426a6e5d},
  {32'hc45873e0, 32'h42a6e1cf, 32'hc407eb7a},
  {32'h43a7b992, 32'hc293cb73, 32'h4266b75d},
  {32'h42de6c94, 32'h428878c2, 32'h438eddbc},
  {32'h44ce4469, 32'h432f77f9, 32'hc28cb66e},
  {32'hc42110b2, 32'h41e60c37, 32'h42b54a64},
  {32'h445f8875, 32'h4290bc04, 32'h431859b8},
  {32'hc412d4a0, 32'hc3cbd1b7, 32'h432ae69c},
  {32'h4413f362, 32'h440446a2, 32'hc1eecf7b},
  {32'hc50019af, 32'h4300f74b, 32'h41f492bc},
  {32'h44f93d40, 32'h423bd778, 32'hc3636f0a},
  {32'hc4a587c5, 32'hc396450f, 32'hc373ab2c},
  {32'h431d8ee0, 32'hc16b75a8, 32'hc266ea3f},
  {32'hc38cd52e, 32'h419df28c, 32'hc3982f7e},
  {32'h435c1ee0, 32'h41895d08, 32'hc3317a46},
  {32'hc4d6be84, 32'hc366df33, 32'hc31bee98},
  {32'h44e0890e, 32'h4295a03e, 32'hc329590a},
  {32'hc505b4e0, 32'h4414193e, 32'h435ecc29},
  {32'h440148fa, 32'hc2a8c3d9, 32'hc100ba4a},
  {32'hc4c79167, 32'hc25fa86d, 32'h43b7d7e0},
  {32'h44d05c68, 32'h43536456, 32'hc381ad4a},
  {32'hc4126cb7, 32'hc1f335e8, 32'hc41a5fb5},
  {32'h44eddc60, 32'h43b1a7d5, 32'hc290904d},
  {32'hc4be7924, 32'hc12350eb, 32'h42ac542d},
  {32'h44656682, 32'hc38c6e70, 32'hc2b33c47},
  {32'hc4d289a3, 32'hc355bef6, 32'hc36da760},
  {32'h44bbb59a, 32'hc3e2d61b, 32'h431fca89},
  {32'hc1fe93c0, 32'hc19129f4, 32'h42ab02b4},
  {32'h449f7b7f, 32'h430a2442, 32'h43b95430},
  {32'hc50ea4b1, 32'h40a81109, 32'h420e2a6e},
  {32'h44fe6ef2, 32'h4366be9f, 32'h438fff5c},
  {32'hc4673ba3, 32'hc3abf2d0, 32'hc302f18d},
  {32'h44b49af8, 32'h42e61b20, 32'h424e9c14},
  {32'hc4bf1a49, 32'hc389af30, 32'hc3460cca},
  {32'h44afa556, 32'h4385370a, 32'h41f07e66},
  {32'hc5128668, 32'hc143a5c1, 32'h40cd4574},
  {32'h4460115c, 32'hc2db16ca, 32'hc30e4a03},
  {32'hc4bb0508, 32'h438a8a0d, 32'hc2bc3b92},
  {32'h44e4bf31, 32'hc2ea1feb, 32'h42b25ef9},
  {32'hc50345dd, 32'h4160aaa2, 32'h439439a1},
  {32'h44e69462, 32'hc3002cfd, 32'h41e9d1a3},
  {32'hc4c60b03, 32'hc315e314, 32'hc3187c8c},
  {32'h4345c750, 32'hc140ee2c, 32'h4314f1eb},
  {32'hc3bf5154, 32'hc18f7a0c, 32'h430b9eb3},
  {32'h4462e656, 32'hc2900a64, 32'h439ac94a},
  {32'hc1e38500, 32'h43b3a472, 32'hc2633450},
  {32'h44e45614, 32'h43500580, 32'hc2b725ec},
  {32'hc51c7b3b, 32'hc3a3a7cd, 32'hc1486b29},
  {32'h4503cbb1, 32'hc3647c5a, 32'h4298b73b},
  {32'hc2a9e250, 32'h4211e7f2, 32'h41de2783},
  {32'h444cc411, 32'hc3c0d978, 32'h3ff9c63e},
  {32'hc4d6b4bd, 32'hc28d2722, 32'hc2309ff2},
  {32'h45079cfa, 32'h42ab9a5a, 32'h43470bca},
  {32'hc34c07b8, 32'h430cd435, 32'h4282b2b8},
  {32'h439cc518, 32'h42e6e3b1, 32'h4193a782},
  {32'hc432cd5e, 32'hc10b8b65, 32'h4300d3f7},
  {32'h440516b5, 32'h42be0c13, 32'h4308260f},
  {32'hc51e988e, 32'hc2e07220, 32'hc38c971a},
  {32'h44d0f1ea, 32'h42cab5d5, 32'h4322f0c9},
  {32'h43ddec9b, 32'hc3b2248e, 32'hc3219aef},
  {32'h4461471d, 32'h43737f64, 32'hc32279a7},
  {32'hc50cfa75, 32'h440b7e59, 32'h43a70f70},
  {32'h44bb29b2, 32'h4403aa2d, 32'hc3023069},
  {32'hc4cea429, 32'h419376d0, 32'h4304ad73},
  {32'h44626a76, 32'hc3a6f6ad, 32'h438f8fb8},
  {32'h417ea900, 32'h428b7e4a, 32'h429939e3},
  {32'h445e766c, 32'hc3d3f4c2, 32'h435cde5b},
  {32'hc4a59e4b, 32'hc297ea79, 32'h434f49c9},
  {32'h44fb57f1, 32'h41baa42c, 32'hc381fc12},
  {32'hc4c075dc, 32'hc2dae224, 32'h4406f9eb},
  {32'h449b1cf2, 32'h4349fb77, 32'hc2e3d690},
  {32'h42c751f0, 32'hc31d0088, 32'hc310880c},
  {32'h44ab0a96, 32'hc23670a9, 32'h4301eeef},
  {32'hc4ae798a, 32'h43e8d13b, 32'h432f39f6},
  {32'h44e53848, 32'h43b6a887, 32'hc332a9da},
  {32'hc48501e6, 32'hc30ce0f0, 32'h439ddf81},
  {32'h441a2fb4, 32'h430a79a3, 32'hc287f493},
  {32'hc39b8610, 32'h438c0403, 32'hc2c1719d},
  {32'h430a0408, 32'hc378282d, 32'h433a8df0},
  {32'hc44b6c94, 32'h432e2da1, 32'h42851ff1},
  {32'h41f67820, 32'h43cf88fe, 32'hc357f137},
  {32'hc44d638a, 32'hc1b79de2, 32'h439a0936},
  {32'h452a675d, 32'hc329991b, 32'h41619544},
  {32'hc2903900, 32'h43a0633a, 32'h432676a7},
  {32'h445bf514, 32'hc297b604, 32'h42d0e8e4},
  {32'hc47e6842, 32'h426807c2, 32'hc400f259},
  {32'h446a2cc6, 32'hc39da285, 32'h4220dc56},
  {32'hc50ac0fe, 32'hc2e2f08f, 32'hc084436e},
  {32'h44b52b2a, 32'hc2d66ed0, 32'hc4029c44},
  {32'hc49b92b2, 32'h400ea2ab, 32'hc32871cc},
  {32'h4452ec13, 32'h41c9f427, 32'hc2c36345},
  {32'hc2b28c30, 32'hc2220da2, 32'hc39459d0},
  {32'h43471050, 32'h42af9bc9, 32'hc22df730},
  {32'hc3f22280, 32'hc317e552, 32'hc32fb4a7},
  {32'h4453931c, 32'hc394b627, 32'hc3262f6c},
  {32'h43aabc7f, 32'hc2241c42, 32'hc257a2a7},
  {32'h430621ac, 32'hc2e3f7d8, 32'hc36b177e},
  {32'hc4d1d928, 32'hc296887e, 32'hc25ede2e},
  {32'h4519cb82, 32'h4357664d, 32'h431c26aa},
  {32'hc4e701e2, 32'hc2181ec8, 32'h42085110},
  {32'h4514998e, 32'hc3fe3b50, 32'h439e9d14},
  {32'hc51c51ec, 32'h432d304d, 32'hc2eb1e23},
  {32'h44b64338, 32'hc2968b22, 32'hc2967132},
  {32'hc4be67ff, 32'hc3d90f83, 32'h42b3fd4f},
  {32'h440a3e0a, 32'h42b3667c, 32'hc2c9c83e},
  {32'hc4c39731, 32'hc30e66cc, 32'hc1a55a7d},
  {32'h44f6f74d, 32'hc31ba7b4, 32'h438824a0},
  {32'hc4f4a28a, 32'hc2c7e8d5, 32'hc31cd166},
  {32'h44edda32, 32'hc2bf902b, 32'h420a44ea},
  {32'hc4b6fe27, 32'h43b4d860, 32'hc3828ba6},
  {32'h44b04e68, 32'hc29bd485, 32'hc30d3549},
  {32'hc3c93fe8, 32'h4268829d, 32'h438746b2},
  {32'h4207ad88, 32'hc33d56ea, 32'hc329e8fd},
  {32'hc5029d1a, 32'h42074958, 32'hc390aac5},
  {32'h44cc1ad4, 32'h4316f1ee, 32'h421d862d},
  {32'hc4cd032a, 32'hc2b140c7, 32'h43eb454e},
  {32'h44d7733e, 32'hc3abd3e0, 32'h41eb514b},
  {32'hc418b006, 32'h4316b08f, 32'hc1281a1a},
  {32'h451c5fe2, 32'hc2507293, 32'hc3146728},
  {32'h430054d0, 32'h439be5cc, 32'hc3c794dc},
  {32'h43f6e4d8, 32'h42d0ad6a, 32'h439c1dc2},
  {32'hc387cd10, 32'hc3941066, 32'hc1324254},
  {32'h44adecdb, 32'hc33fa934, 32'h438a8862},
  {32'hc38f74bc, 32'h425c61b8, 32'hc36a618a},
  {32'h44e455f9, 32'hc10a5444, 32'hc3802882},
  {32'hc5077d1c, 32'h41ea052e, 32'hc31c8582},
  {32'h43e58430, 32'hc360097d, 32'h430286a8},
  {32'hc4644a2a, 32'hc36b81cf, 32'hc36a4c60},
  {32'h450ba5be, 32'hc34cae26, 32'h43bfeeaf},
  {32'hc3eae1af, 32'hc36e9272, 32'hc3a4563b},
  {32'h441c83e8, 32'h43866377, 32'h421e9f8a},
  {32'hc4cfd008, 32'hc3c3ad99, 32'h4241c6c7},
  {32'h4434fd71, 32'h42dbf80e, 32'h42c1ba32},
  {32'hc486c001, 32'h441984d8, 32'hc2973636},
  {32'h452176bb, 32'hc2811482, 32'hc3c5da8a},
  {32'hc488c24c, 32'hc32252b4, 32'h43105b99},
  {32'h44d5ce56, 32'hc35a0c49, 32'hc2962920},
  {32'hc4560558, 32'h422c348b, 32'h435d5317},
  {32'h451073b6, 32'hc29944bf, 32'hbfc53670},
  {32'hc4f0a228, 32'hc0836c99, 32'h4312bf40},
  {32'h44dc69fe, 32'hc1e86ead, 32'h425daa3a},
  {32'hc4313b36, 32'hc34b13ba, 32'hc220f19f},
  {32'h4450cfec, 32'h429be13f, 32'h43c67392},
  {32'hc4689c31, 32'hc315688a, 32'hc1218216},
  {32'h44d29eb0, 32'hc2f7da62, 32'h42b06238},
  {32'hc4e701be, 32'hc2fc08ae, 32'h4359f2da},
  {32'h44f14105, 32'h436c377b, 32'hc2f36194},
  {32'hc3c34e16, 32'hc2a230c7, 32'hc3f61930},
  {32'h44169a68, 32'h42d0e684, 32'h42a2c0b8},
  {32'hc45b639c, 32'h43a847e5, 32'h432c7133},
  {32'h45063634, 32'h4229a0e6, 32'hc2ef83f8},
  {32'hc406432c, 32'h43298104, 32'hc2c69150},
  {32'h44f3935b, 32'h43b1b5d2, 32'h43311e8e},
  {32'hc4624bac, 32'h43d3031b, 32'hc341a558},
  {32'h44b94170, 32'hc2e42523, 32'h42fc6f96},
  {32'hc4e634da, 32'hc3064540, 32'hc307205b},
  {32'h44d4a473, 32'hc26a5bf8, 32'h430e0f77},
  {32'hc45668c2, 32'h43b34ee1, 32'h4230ef5f},
  {32'h447f62c4, 32'h4296b2fa, 32'h42c21903},
  {32'hc3c63470, 32'h424f1a8e, 32'hc34cc89f},
  {32'h44d7039b, 32'hc214f3a8, 32'h434c3153},
  {32'hc4b614f0, 32'h432e5e27, 32'hc283de39},
  {32'h4474dd56, 32'h4278530c, 32'hc32d11ba},
  {32'hc35e3af0, 32'hc241214e, 32'hc237dc05},
  {32'h444682fb, 32'h43a0135f, 32'hc354a44c},
  {32'hc502ba83, 32'h436cf2f3, 32'hc27ab62a},
  {32'h44a7f8a0, 32'hc208cf12, 32'h43c7ca88},
  {32'hc325314c, 32'h43162738, 32'hc346fc7c},
  {32'h443950cd, 32'hc31eb1af, 32'h441cd40a},
  {32'hc500ff7a, 32'h41df28de, 32'h435d012e},
  {32'h44627d9e, 32'h433cd52f, 32'h42f1bdc8},
  {32'hc280c408, 32'h43401dfe, 32'hc3912727},
  {32'h4434ec6d, 32'hc395c101, 32'hc2219c05},
  {32'hc5153039, 32'h434a34ae, 32'h433d79a8},
  {32'h44f07c55, 32'h418fff12, 32'h438a8b01},
  {32'hc3c05780, 32'hc3ccbcbe, 32'hc3f94a8a},
  {32'h445f516c, 32'h43327b4e, 32'h4296e14a},
  {32'hc4dabd55, 32'hc195e054, 32'hc28ffc75},
  {32'h44f396bb, 32'hc2dbb429, 32'hc39525d4},
  {32'hc4342b06, 32'h43084c82, 32'h4357b5cd},
  {32'h44410104, 32'hc38ec286, 32'hc25903cc},
  {32'hc4cca1a4, 32'hc2a61ae4, 32'hc402d391},
  {32'h434ffe94, 32'hc37eff19, 32'h43aec293},
  {32'hc4b7f080, 32'hc37f7470, 32'hc04a8d46},
  {32'hc4d8fd7a, 32'hc11914dc, 32'h42a6fee2},
  {32'hc2239c10, 32'h4028ba86, 32'h42ce4561},
  {32'hc5094f52, 32'hc2f57159, 32'hc3384c6e},
  {32'h43f3a2ba, 32'hc35b3a23, 32'h43999dca},
  {32'hc4fb9f39, 32'h4199edda, 32'h42ead50f},
  {32'h443a6b59, 32'hc22e9cef, 32'hc30f267b},
  {32'hc39ef6a8, 32'hc3b89a57, 32'hc32bc4b0},
  {32'h44a9c9fa, 32'h43185641, 32'h43804c71},
  {32'hc49d306b, 32'h431a7976, 32'h424505a6},
  {32'h43c88610, 32'hc406127f, 32'hc2511f78},
  {32'hc4fc8446, 32'h42bd6d4d, 32'hc2177ffe},
  {32'h44e91559, 32'hc30a0ef0, 32'h4295703c},
  {32'hc4f772b1, 32'h42ca2fba, 32'h43e06a2d},
  {32'h45041c32, 32'h438ef191, 32'h42b3cb05},
  {32'hc49d0721, 32'h42ec2719, 32'hc3114bfa},
  {32'h44c767ff, 32'h41e92606, 32'h42e9bedc},
  {32'hc4aab9c3, 32'hc1861893, 32'h430ea243},
  {32'h450bfded, 32'hc3784bf8, 32'h43a900c2},
  {32'hc5008b02, 32'hc205dbcc, 32'hc3285c17},
  {32'h4442e67e, 32'h41bd95d5, 32'h43557107},
  {32'hc46a7a93, 32'h4307f5be, 32'hc3033e0c},
  {32'h44b5eb31, 32'hc1e1eb81, 32'hc0c7c213},
  {32'hc4894390, 32'hc31191a9, 32'hc3dbee58},
  {32'h4303ef30, 32'hc2ab0f3a, 32'h433d40ce},
  {32'hc3b298ea, 32'h418c9dfa, 32'hc1ab043a},
  {32'h44f5b85c, 32'h4314241e, 32'hc2e5f5ba},
  {32'hc4b7efa0, 32'h430661c0, 32'h42fbdd92},
  {32'h44e3737a, 32'hc32f23d7, 32'h430a969a},
  {32'hc42d35da, 32'hc204156c, 32'hc3949814},
  {32'h448181d7, 32'h431dbc4d, 32'h41dd6f4f},
  {32'hc50268a3, 32'hc332da60, 32'h42adba5f},
  {32'h436c3d40, 32'hc326ed1f, 32'h417bef63},
  {32'hc491f90a, 32'hc2454b5e, 32'hc275c423},
  {32'h440e85ee, 32'h434783fd, 32'hc30ef968},
  {32'hc50558be, 32'hc32477e4, 32'h4367b077},
  {32'h447458b2, 32'hc301287b, 32'hc38ae671},
  {32'hc4b3d8d0, 32'hc2fa782f, 32'hc3b1012a},
  {32'h44c0ab3a, 32'hc264e284, 32'hc19b65f6},
  {32'hc2f04080, 32'h43313796, 32'h43205fa6},
  {32'h44f88ba3, 32'h43aaf45f, 32'h438040a3},
  {32'hc511a26d, 32'h4236f922, 32'h4390b5e6},
  {32'h443d10d2, 32'hc293353e, 32'h43850372},
  {32'hc2ff9bb0, 32'h43949cf9, 32'h434845c0},
  {32'h41822dc0, 32'hc3a79c30, 32'h43ba2130},
  {32'hc45ef584, 32'hc327d565, 32'h42ea01ea},
  {32'h442860ce, 32'hc2942589, 32'h431e8780},
  {32'hc4c0116c, 32'h42c1cf6b, 32'h438c34ab},
  {32'h44448dbc, 32'hc384ae20, 32'hc1c120d6},
  {32'hc40d6818, 32'h432a2e75, 32'hc244424b},
  {32'h448ea3d7, 32'h42d2e3e2, 32'h435b8092},
  {32'hc4c185fb, 32'hc375b6ce, 32'hc258fae7},
  {32'h44341f6c, 32'hc309f9ae, 32'h4378d211},
  {32'hc506d058, 32'h42d30b7a, 32'h42ad4b23},
  {32'h44fe5ebf, 32'hc399ff3e, 32'hc25dcf90},
  {32'hc4812db4, 32'h43886bfa, 32'h42a3b1d6},
  {32'h447fd4ae, 32'h42c25d35, 32'hc332e4fa},
  {32'hc42ca9bc, 32'h4367e0ab, 32'h430e3414},
  {32'h44eaca68, 32'h43d3e638, 32'hc2c8f0d7},
  {32'hc4bec48c, 32'hc00d62da, 32'h437f147e},
  {32'h44d19190, 32'h436cdf17, 32'h43bb689e},
  {32'hc3f89808, 32'h42250ae4, 32'hc223cebe},
  {32'h448bbe37, 32'hc2182c6d, 32'hc07a8520},
  {32'hc4d919d1, 32'hc3d48b95, 32'hc29800b5},
  {32'h446cb766, 32'h41ecccd4, 32'hc2c84711},
  {32'hc47d37c4, 32'hc35cfec1, 32'h438b98ba},
  {32'h450b7b6e, 32'h441cabda, 32'hc2e08400},
  {32'hc47e9e34, 32'h43220cec, 32'h4296c13f},
  {32'h441b6024, 32'hc3214ba6, 32'hc30d3884},
  {32'h4201b540, 32'h4381b8ed, 32'h42a370ca},
  {32'h4405d7ac, 32'hc2bcd394, 32'hc221b1f3},
  {32'hc38c6240, 32'h4371e696, 32'h41390b58},
  {32'h42e32fc4, 32'hc30a912f, 32'h4330308c},
  {32'hc5029c8a, 32'hc33188d9, 32'h439e459a},
  {32'h439e7f99, 32'hc255d4bd, 32'h4292e211},
  {32'hc2a98aa0, 32'hc35633b4, 32'h4339e836},
  {32'h44e5659f, 32'h4335ff92, 32'hc30d4dba},
  {32'hc4f7972d, 32'h4340fe61, 32'h42ec0527},
  {32'h433fe0ce, 32'h4357fed6, 32'hc3e6d294},
  {32'hc4d877cb, 32'h433e3322, 32'h43172266},
  {32'h448685ae, 32'h43a7d6fe, 32'h439b82d3},
  {32'hc5039daa, 32'hc3b4412d, 32'hc3b771c6},
  {32'h44365591, 32'hc25167c9, 32'hc3af3d1a},
  {32'hc35b9d4b, 32'h43ff20ae, 32'h437b9d5f},
  {32'h45091dbe, 32'h42ca1351, 32'h40bef6cf},
  {32'h42f9c3e6, 32'hc3476829, 32'hc3909fbc},
  {32'h4516e55e, 32'h436ebe5f, 32'h4311a91b},
  {32'hc4291e0c, 32'h41ff6607, 32'h4023add3},
  {32'h44f7810f, 32'h436eb827, 32'hc3939e67},
  {32'hc43375a4, 32'h41e3c443, 32'hc25817f0},
  {32'h44d27131, 32'hc350009a, 32'h422383a6},
  {32'hc4028644, 32'h423700f0, 32'hc2d2047c},
  {32'h4507e986, 32'h411188d8, 32'hc336935b},
  {32'hc4e3b2a0, 32'hc2b335d2, 32'hc33263bc},
  {32'h4356ef18, 32'h42a1d430, 32'hc3751899},
  {32'hc4fd4ec5, 32'h43f2f086, 32'h4336a045},
  {32'h44dee41e, 32'hc368275d, 32'hc31c574d},
  {32'hc437eb72, 32'h4377eb1b, 32'h4371a28b},
  {32'h44702f3b, 32'h4363b5f6, 32'h426cd642},
  {32'hc4ec975f, 32'h435fa2b9, 32'hc3899380},
  {32'h443442e0, 32'hc33254d2, 32'h43c2583b},
  {32'hc4be3976, 32'hc3611892, 32'h42842c0a},
  {32'h4399ee7c, 32'hc3a4d0fd, 32'h42576ba5},
  {32'hc45dce36, 32'hc3ea874c, 32'h43c358b7},
  {32'h447d76b0, 32'hc3bd81d4, 32'h424dea8a},
  {32'hc4c7bd54, 32'h42f2af3b, 32'h433155dc},
  {32'h43e03bae, 32'hc2a66939, 32'hc3b5c93a},
  {32'hc3b7defe, 32'h42538593, 32'hc2c724a2},
  {32'h43ef7bc4, 32'hc42c29b0, 32'hc3b70ea5},
  {32'hc490dec6, 32'hc24b37ce, 32'hc140978a},
  {32'h44c95596, 32'hc16eae8c, 32'hc266bf9e},
  {32'hc4cc821d, 32'h4384d8cf, 32'h434cc218},
  {32'h43e62104, 32'hc1dcc69c, 32'h43e85276},
  {32'hc4371e92, 32'hc293f7e5, 32'hc298a1cf},
  {32'h4469141f, 32'h426a1124, 32'hc2b519a7},
  {32'hc4e0bfea, 32'h43bcd4ec, 32'h4398a354},
  {32'h424d11a0, 32'h418638a9, 32'hc3bc2c95},
  {32'hc4a46d5c, 32'h439900d7, 32'hc19f9ffe},
  {32'h4432473e, 32'hc39c0e69, 32'hc397b06f},
  {32'h4250cb60, 32'h43a94d08, 32'h430f2fbe},
  {32'h45049797, 32'h431319c8, 32'h4282b886},
  {32'hc406bb9a, 32'h438b0da8, 32'hc336391a},
  {32'h45164d52, 32'hc31c4861, 32'hc2f1fa44},
  {32'hc427ecf9, 32'hc1754ce2, 32'h4332417d},
  {32'h44d095e4, 32'h42db2ab1, 32'hc33a20d8},
  {32'hc4e0c9b5, 32'hc3a2d5f7, 32'h42777539},
  {32'h44bdb601, 32'h41e37df1, 32'hc1fbad0c},
  {32'h42cc1f06, 32'hc2803024, 32'hc2f770d3},
  {32'h44ef31bf, 32'h42fd09da, 32'h43a57bf5},
  {32'hc49b83b0, 32'h430b4b98, 32'hc297e314},
  {32'h4086f1c0, 32'h436d73c3, 32'h40c42248},
  {32'hc4dc624c, 32'h4401567f, 32'hc29fc83a},
  {32'h44ff4164, 32'hc382d921, 32'h430b7624},
  {32'hc4fe4bfe, 32'hc2879b76, 32'h43b68476},
  {32'h439f9094, 32'hbed13180, 32'h4334c99d},
  {32'hc4b8d86c, 32'hc3420c57, 32'h4224fd7f},
  {32'h44c17e4c, 32'hc3783e1b, 32'h41eb0458},
  {32'hc42a4a98, 32'h4161415f, 32'h43ef8bf4},
  {32'h449df1f4, 32'h43c71d87, 32'hc2bf91c5},
  {32'hc504b232, 32'hc39c3a54, 32'h439a1df9},
  {32'h4404cbf4, 32'hc3d48a8a, 32'h438d3f9a},
  {32'h42f96df0, 32'h436f37b9, 32'h4396cc29},
  {32'h44b83181, 32'h4244c272, 32'hc332a8f1},
  {32'hc43c384e, 32'h42e6e831, 32'h43707557},
  {32'h44fe2cf2, 32'hc301918b, 32'h431cb75e},
  {32'hc38040a8, 32'hc3b6b20b, 32'h43430971},
  {32'h44b2af05, 32'h439a8f6a, 32'hc40cd324},
  {32'hc42bd1f7, 32'h441751df, 32'h438e94cd},
  {32'h447506dc, 32'hc38123be, 32'h43258123},
  {32'hc3c711a8, 32'hc29014f0, 32'h44059544},
  {32'h446fca6f, 32'h4371a9b6, 32'hc39de282},
  {32'hc4734cdc, 32'h4184cc8e, 32'hc30ea224},
  {32'h448d1945, 32'h43c61d04, 32'h42f56c80},
  {32'hc3b9f7a0, 32'hc3830829, 32'hc37cf8d6},
  {32'h4449b1b9, 32'h4321026f, 32'hc2cae161},
  {32'hc3da5a07, 32'h436f2578, 32'h42b1b358},
  {32'h450b76a4, 32'hc28e6b63, 32'h42f8a6b3},
  {32'hc4fc7a69, 32'h437b1b48, 32'h4246403c},
  {32'h43113c52, 32'hc35793b3, 32'h43ad6e5a},
  {32'hc49ef072, 32'hc380c204, 32'h42bc5904},
  {32'h42f5ee50, 32'h4279188a, 32'hc28c9326},
  {32'hc4a46f88, 32'h42bda648, 32'h421fc605},
  {32'h44fade52, 32'h43a64006, 32'h4204e8b1},
  {32'hc4d87824, 32'hc254b6e5, 32'hc2a69bb5},
  {32'h440d460c, 32'h43602933, 32'hc2f38d41},
  {32'hc27ca0c0, 32'hc336d146, 32'h43cb750a},
  {32'h44717d3c, 32'h4343d2e4, 32'h43aa5a17},
  {32'hc40f0e64, 32'h43a1ab7c, 32'hc3968d87},
  {32'hc34eec39, 32'h440a26e5, 32'hc38a4105},
  {32'hc44ad3b0, 32'h42903050, 32'hc38cd035},
  {32'h437d20e0, 32'hc39bfb8d, 32'h435f4bd7},
  {32'hc47e3496, 32'h4213a2e8, 32'hc3283b2a},
  {32'h44b9d142, 32'h41c495dd, 32'hc38f90db},
  {32'hc4a34a8f, 32'hc3c957dd, 32'h43a93bb9},
  {32'h4438fd3d, 32'hc3358b5e, 32'hc4142583},
  {32'hc4a407d3, 32'h4329f691, 32'h428a8505},
  {32'h433785da, 32'h42c4b0a2, 32'h4206f3d0},
  {32'hc3c282eb, 32'h4301ea5f, 32'hc32359eb},
  {32'h43f1a0cc, 32'hc31e1464, 32'hc2fdd570},
  {32'hc46b9869, 32'h42855147, 32'hc3ae39d4},
  {32'h405d6400, 32'hc34190f3, 32'h4242a164},
  {32'hc502e51c, 32'hc34352bd, 32'h419232b4},
  {32'h4480208c, 32'h43e5e80b, 32'h4339050f},
  {32'hc4d13d17, 32'hc38a4e2e, 32'h439bc6f2},
  {32'h44d50f93, 32'hc3052c8c, 32'hc30120ca},
  {32'hc3b83328, 32'h436d69fd, 32'hc38d1918},
  {32'h43bdfd3a, 32'h42adec7a, 32'h439ae7a3},
  {32'hc4d3d833, 32'h429f0acb, 32'h43383dcb},
  {32'h449d30a9, 32'hc39e68a4, 32'hc2b43e7d},
  {32'hc40ed714, 32'h42a960bd, 32'h421e41b4},
  {32'hc31b99d5, 32'hc0e7c252, 32'h422970da},
  {32'hc5056867, 32'h42cdf7b2, 32'hc34255a7},
  {32'h43c17ac8, 32'h43925e50, 32'h4349fb18},
  {32'hc4a031e8, 32'h4319622d, 32'hc298a79e},
  {32'hc2551cc0, 32'hc32da3e1, 32'h4198a99b},
  {32'hc4fd8bb0, 32'hc2eab0ec, 32'hc30b6306},
  {32'h451be3c6, 32'h4304d7bf, 32'h437a6806},
  {32'hc4fd2f04, 32'h42e3a921, 32'h40b9d9bb},
  {32'h43a2e179, 32'hc2916a1a, 32'h42014f9c},
  {32'hc4b01030, 32'hc2af9436, 32'h441ab4f3},
  {32'h43e16d70, 32'h42285a35, 32'h435566c1},
  {32'hc2ac1880, 32'hc2fc9ce9, 32'h4263ec99},
  {32'h43d676cc, 32'h4345e1e0, 32'h43e3aeb6},
  {32'hc378e6d4, 32'h43c7d360, 32'h42a65be7},
  {32'hc3388150, 32'h43ae7a34, 32'h42ef1ac6},
  {32'h41625200, 32'h431dfd5e, 32'h433f9c2e},
  {32'h44db2dd6, 32'h4340fb4a, 32'h42fee276},
  {32'hc4cf4118, 32'hc3a467ed, 32'h4391811a},
  {32'hc32db788, 32'h4308e8ce, 32'hc33c1460},
  {32'h4348a5a8, 32'h40b40e7c, 32'h4387b281},
  {32'h4506f877, 32'h4228b0ed, 32'hc377e5d9},
  {32'hc4ae5689, 32'hc2376435, 32'h41e06ec2},
  {32'h45077b9e, 32'hc2910562, 32'hc4245663},
  {32'hc428cfde, 32'h4388a1b4, 32'h4327fc91},
  {32'h4497ee2d, 32'h42642a06, 32'h4311e7e0},
  {32'hc4a0e280, 32'h43f5455d, 32'h438c6102},
  {32'h44cbb658, 32'hc316e849, 32'hc357a4d0},
  {32'hc4fbb0dc, 32'hc3a3def4, 32'hc38f4806},
  {32'h44758aa2, 32'h4333008d, 32'h4282ee42},
  {32'hc458c206, 32'hc2141497, 32'h43fa9c95},
  {32'h442f0167, 32'h43a0caf9, 32'hc38692fe},
  {32'hc28b9f76, 32'h430553ab, 32'h4121536a},
  {32'h442d5ba4, 32'h43654fe1, 32'h43afcb93},
  {32'hc43cb91a, 32'h436f2f79, 32'h4383a2c0},
  {32'h43b828a8, 32'hc200c58f, 32'hc39a9f5e},
  {32'hc4f5fca2, 32'hc2e090ef, 32'hc16b64da},
  {32'h450573ea, 32'hc1f6c77f, 32'h42660747},
  {32'hc4b70333, 32'h43fb451d, 32'h44022444},
  {32'h44eca259, 32'hc32a7c7f, 32'h43812c80},
  {32'hc44c802a, 32'hc3b6d541, 32'h431f058b},
  {32'h4502beba, 32'hc397301f, 32'hc31f7274},
  {32'hc4264e20, 32'hc35e3f7d, 32'hc0dd1e68},
  {32'h443552f8, 32'hc312f4b3, 32'hc3bbb92d},
  {32'hc49d4771, 32'hc186938d, 32'h4373d576},
  {32'h44b77609, 32'hc39c11d3, 32'hc2ef7dd8},
  {32'hc455b244, 32'hc34a81aa, 32'hc3c48283},
  {32'h4502091b, 32'hc3c2af6e, 32'h428081c5},
  {32'hc418dee0, 32'hc41790ed, 32'h42a94bff},
  {32'h44c0907a, 32'hc3b67d0d, 32'hc3b4068d},
  {32'hc437f96f, 32'h40bd98bc, 32'hc38ea1a4},
  {32'h4451e3e9, 32'hc33b8836, 32'hc20f5e78},
  {32'hc3ab55a0, 32'hc38a6cfe, 32'hc2d09152},
  {32'h44ddbc38, 32'h4293d931, 32'hc27cdda1},
  {32'hc3efea8c, 32'hc3da35e6, 32'hc3e72ae3},
  {32'h44d2b979, 32'hc3d7a98a, 32'hc2f37ac9},
  {32'hc3b70c52, 32'hc2bf02ba, 32'h42512de3},
  {32'h45277733, 32'hc38c516e, 32'h42e61670},
  {32'hc41da3a7, 32'h423bde09, 32'h4310d5a5},
  {32'h4408366f, 32'hc34f11f4, 32'h4319be7b},
  {32'hc4fd0750, 32'hc29f7df0, 32'hc3c6a801},
  {32'h45019cdb, 32'hc3b0c480, 32'h438ab288},
  {32'hc3c8e577, 32'h43aaf0e0, 32'h430c5f75},
  {32'h44152b51, 32'hc326c695, 32'hc366b501},
  {32'hc4bd03e1, 32'hc3188ae0, 32'hc1f9cdb8},
  {32'h44b13cb0, 32'h41213b93, 32'hc35d93b7},
  {32'hc4550bd2, 32'hc2064dd1, 32'h422068eb},
  {32'h45048f2f, 32'h436b2dd2, 32'hc3494459},
  {32'hc4805f5e, 32'hc1ee17b3, 32'hc2c97bbe},
  {32'h44e371ed, 32'h43692035, 32'h42f794a7},
  {32'hc4dceb6f, 32'h43ad831f, 32'h41ab9f01},
  {32'h44a6caa9, 32'hc306659e, 32'hc3b8f5f2},
  {32'hc3d9ce25, 32'h42c8a042, 32'h43ca9bb8},
  {32'h4485ec96, 32'hc343ca33, 32'h43192e57},
  {32'hc484b09b, 32'h4318ac50, 32'h429eb1fe},
  {32'h448bf7da, 32'h418b45f8, 32'hc3b9c836},
  {32'hc4ae69c6, 32'hc3ff3438, 32'hc220b2a3},
  {32'h44bf58c2, 32'hc273c379, 32'h4352081a},
  {32'hc50950c6, 32'h4342ab16, 32'hc3cc90e0},
  {32'h43c4b77c, 32'h416ddd3c, 32'h4343afae},
  {32'hc506919d, 32'hc33ec7fa, 32'h425c8cd6},
  {32'h43b66686, 32'hc2bcbb1e, 32'h438f1df9},
  {32'hc4953d7e, 32'hc1904f8a, 32'h43b768d5},
  {32'h450ab6c5, 32'hc3ae2313, 32'h42aa550c},
  {32'h42524869, 32'hc3e2d659, 32'hc1195ef6},
  {32'h44ea323e, 32'hc13938f6, 32'hc2b10070},
  {32'hc38f61be, 32'h43346907, 32'hc2f68b4a},
  {32'h4249b220, 32'h438f41da, 32'h42eeaadc},
  {32'hc5196718, 32'h435e83cc, 32'h437ee06e},
  {32'h44204dca, 32'h43ebab0d, 32'hc2465c0d},
  {32'hc48b5a7c, 32'h41db13bd, 32'hc37e4f7e},
  {32'h42b9fa38, 32'h4309dbe7, 32'hc34a20ca},
  {32'hc50abd48, 32'hc2bcd738, 32'h4399051e},
  {32'h43fff824, 32'h429d1017, 32'hc3a9aeff},
  {32'hc36759b8, 32'h4270b982, 32'h4358bf5d},
  {32'h44e0d937, 32'h429f8a15, 32'h43ab26aa},
  {32'hc4170a8b, 32'hc33cf04e, 32'h43807df0},
  {32'h4456925c, 32'hc38ea6e1, 32'h436057ac},
  {32'hc465fbb5, 32'h413601e3, 32'h3f33ca38},
  {32'h44d820d5, 32'h418f23e1, 32'h433babdf},
  {32'hc4b232fc, 32'hc38ff7c3, 32'h42e9857f},
  {32'h430332b0, 32'hc290b8ea, 32'h43949e8b},
  {32'hc51ebbcf, 32'h42b56da8, 32'hc391277f},
  {32'h43d9e01c, 32'hc2455bd4, 32'h41dd8c7f},
  {32'hc4311c02, 32'h431878fe, 32'hc3511e55},
  {32'h4404a2f9, 32'h440ba404, 32'h41063db4},
  {32'hc50c8292, 32'hc33eec6b, 32'hc39d6322},
  {32'h4389c60c, 32'hc365a942, 32'h42d07587},
  {32'hc4caa8e0, 32'h41f1a390, 32'hc29194c8},
  {32'h448a0c92, 32'hc28bc884, 32'h438dab7e},
  {32'h43477399, 32'hc30ea4e6, 32'h430ac91a},
  {32'h44b47808, 32'h422b4c50, 32'hc2879061},
  {32'hc4f4d132, 32'h43eaba5e, 32'h4321fc72},
  {32'h435bfdc4, 32'h43a0412c, 32'hc391b83a},
  {32'hc50f80f1, 32'hc328f91c, 32'h43a9ec2c},
  {32'h45200566, 32'h40a58118, 32'hc33ae97f},
  {32'hc4cd8cff, 32'h41b96c20, 32'h42665cbe},
  {32'h44aa52b5, 32'hc41953c4, 32'h430e488e},
  {32'hc49d7614, 32'h4202c096, 32'hc36e057d},
  {32'h444cabec, 32'h4326e4d8, 32'h4247c74d},
  {32'hc4ecae16, 32'h415907f5, 32'h4286d235},
  {32'h43c53462, 32'h42432ab8, 32'hc2f49844},
  {32'hc321dcf0, 32'h433354cc, 32'hc2c5c472},
  {32'h4485b6f0, 32'hc2cb5a3e, 32'hc336d14e},
  {32'hc514d1d4, 32'hc1616d15, 32'h3faac09a},
  {32'h4437089a, 32'h42b8d177, 32'hc334037f},
  {32'hc5099560, 32'h41e4a79a, 32'hc3ffed27},
  {32'h4499362e, 32'hc32c81c2, 32'h4009c18c},
  {32'h43699b3d, 32'h4252b9d0, 32'h437470b3},
  {32'h446a5290, 32'hc30871a0, 32'hc2d53e62},
  {32'hc42aec36, 32'h43e9c301, 32'hc315b9de},
  {32'h44f14727, 32'hc0d14305, 32'h43345bce},
  {32'hc3e43318, 32'hc38dc018, 32'hc389c69c},
  {32'h44a0163a, 32'hc3bca0b5, 32'hc3455ab2},
  {32'hc33abde8, 32'h432d5289, 32'hc2e45bd8},
  {32'h449e1f84, 32'hc2960c3f, 32'h432a0bbb},
  {32'hc4bac19c, 32'h42ac984c, 32'hc34c4742},
  {32'h43cbc395, 32'hc2fa5085, 32'h42453fc7},
  {32'hc4c92840, 32'hc39f32c1, 32'h438f5b86},
  {32'h44d3109c, 32'hc3033d81, 32'hbf6b2dbe},
  {32'hc50ef7a0, 32'hc34e7892, 32'h439847fd},
  {32'h44df2b57, 32'h42c99784, 32'h4332a8ea},
  {32'hc3f42f40, 32'hc387b34d, 32'hc390a6c6},
  {32'h44d5c0a7, 32'hc307c734, 32'h434ffa51},
  {32'hc38f00d8, 32'h42db6763, 32'hc1ee8126},
  {32'h444b2d72, 32'hc2b08330, 32'h41fc74ed},
  {32'hc5006748, 32'hc316b225, 32'hc1d0cdad},
  {32'h43e8e2e8, 32'hc27ac549, 32'hc29dd2ed},
  {32'hc520564e, 32'h43206741, 32'h432ab56e},
  {32'h42f81e70, 32'h438d2191, 32'hc3d966dd},
  {32'hc4fa0cd0, 32'hc321c6cb, 32'h426c0865},
  {32'h44d59c5a, 32'h42bce068, 32'h43971626},
  {32'hc484318e, 32'h4246ac7a, 32'hc166955e},
  {32'h45100984, 32'h438e51b4, 32'hc3640aa9},
  {32'h439480cd, 32'hc23ac4e4, 32'h4288aa10},
  {32'h44bb4208, 32'hc23bd1d4, 32'h42c2607a},
  {32'hc3b6dfb5, 32'h42813772, 32'hc31da02f},
  {32'h43b6db67, 32'h4313e36e, 32'hc39decb3},
  {32'hc500de07, 32'hc3365559, 32'hc27d2131},
  {32'h44ee0966, 32'hc2f5b0fa, 32'hc38ca1c5},
  {32'hc4c34632, 32'hc20326d6, 32'h429df661},
  {32'h43378ed8, 32'hc2c01a5d, 32'h42bcd257},
  {32'hc4ff33d0, 32'h4283f6bc, 32'h42043a44},
  {32'h438b15a8, 32'hc3477755, 32'hc2804df8},
  {32'hc4969030, 32'hc1c780ba, 32'h4398dc47},
  {32'h44c507a5, 32'hc3628e13, 32'h43167713},
  {32'hc4e96c1e, 32'h4004f5ee, 32'h40936260},
  {32'h451af50e, 32'h425a5366, 32'hc388c79f},
  {32'hc3d98508, 32'hc1d7c7cd, 32'h4393a52e},
  {32'h448ac7aa, 32'h42e75ca5, 32'h439a6642},
  {32'hc4c63ea6, 32'hc20d3b07, 32'hc23e03a6},
  {32'h4449e9ae, 32'hc10c545d, 32'hc3230f24},
  {32'hc508d8d6, 32'hbf926212, 32'hc3151dbe},
  {32'h4483569d, 32'hc2556958, 32'hc3751fdf},
  {32'hc42f0b70, 32'hc1fe802b, 32'hc3e6321b},
  {32'h44fa4d6e, 32'h434d85f8, 32'h420369a9},
  {32'hc28fe3ba, 32'hc32c2639, 32'hc35987d2},
  {32'h4395d528, 32'hc37cacbd, 32'hc3644532},
  {32'hc506567e, 32'hc2d31240, 32'hc3ba1856},
  {32'h45051026, 32'h43443f96, 32'hbfca9ed0},
  {32'hc4cc8871, 32'h41acc0e6, 32'hc32cc959},
  {32'h448607d8, 32'hc24a4438, 32'hc40a3231},
  {32'hc4df94f8, 32'hc3ac3827, 32'h43917e1a},
  {32'h446c3b80, 32'h42845848, 32'hc1818d61},
  {32'hc5016562, 32'h42e34c4e, 32'h42559ffb},
  {32'h4484ef7a, 32'hc2caccba, 32'hc32069c8},
  {32'hc484284d, 32'hc3b6b72e, 32'hc2b39976},
  {32'h44fb3e18, 32'hc2ba44b3, 32'h42a62707},
  {32'hc51fd286, 32'hc2d995b6, 32'hc2d26b21},
  {32'h451169e6, 32'h439f468f, 32'hc30426e3},
  {32'hc4ba216e, 32'h42b2c108, 32'hc2c4f63e},
  {32'h44c2baa9, 32'hc1ded4bb, 32'hc3308f29},
  {32'hc49b0ab7, 32'h41cda697, 32'h43287a32},
  {32'h44fa2689, 32'h4326fb7f, 32'h43b56de3},
  {32'hc2363c4c, 32'h4291bd23, 32'h435fa50a},
  {32'h4419ca68, 32'hc2332965, 32'h43227116},
  {32'hc3ef0f91, 32'h43979fdf, 32'hc2c419f8},
  {32'h4507e917, 32'hc209e71b, 32'hc2e5e2f8},
  {32'hc36c0a4f, 32'h436c8a87, 32'h438a3b6b},
  {32'h45151949, 32'hc3127358, 32'h42ded9b0},
  {32'hc3d87dc8, 32'h430de4e1, 32'hc2f062a4},
  {32'h4506eecc, 32'hc1a5f35c, 32'h42378ae4},
  {32'hc1cc0580, 32'hc30ba195, 32'h43a840cc},
  {32'h4333f5e0, 32'hc3884e35, 32'hc3b19410},
  {32'hc4a6b8ad, 32'hc2cda3f7, 32'hc3744a37},
  {32'h43e44920, 32'h418494e7, 32'h42a8f52e},
  {32'hc4518e7c, 32'h43580e90, 32'hc3b9abea},
  {32'h44f1805c, 32'hc2a56e04, 32'h420058ab},
  {32'hc4373250, 32'h402a63d8, 32'h4207dd02},
  {32'h44248535, 32'hc3935b82, 32'hc2d7789d},
  {32'hc4a84e30, 32'h42b9694e, 32'h4282fc69},
  {32'h44ec012e, 32'h4391387e, 32'hc396c137},
  {32'hc4afca22, 32'h43858018, 32'hc386459a},
  {32'h44f53308, 32'h426f2d42, 32'h41c78412},
  {32'hc50924f4, 32'hc2f11738, 32'h429639a7},
  {32'h44ca0322, 32'hc38f467d, 32'h430f367c},
  {32'hc3d50500, 32'hc2a26bac, 32'h43c45a3a},
  {32'h451e64c4, 32'hc0d56ddd, 32'h3f9bf758},
  {32'hc344fc80, 32'h438f7dd9, 32'h43c52602},
  {32'h4425b93c, 32'hc28970eb, 32'hc3aaad1e},
  {32'hc4aee724, 32'h43942d68, 32'h43e9558e},
  {32'h4505a65c, 32'h41dc04f2, 32'hc3102c1b},
  {32'hc50582c5, 32'h43916a94, 32'hc2fed116},
  {32'h44b213d9, 32'hc32fc41f, 32'h43423f1a},
  {32'hc4ce09c3, 32'hc1a12025, 32'h4358aa05},
  {32'h443269d0, 32'hc3bcd07f, 32'hc272510a},
  {32'hc3394ac4, 32'hc282e97b, 32'hc369bcb7},
  {32'h44a08045, 32'hc2e2b00d, 32'hc1bbad4e},
  {32'hc422d1d0, 32'hc30b23cc, 32'h43f0fd87},
  {32'h44ea5900, 32'h413ca8af, 32'hc2cf9965},
  {32'hc44de7d0, 32'hc36c5130, 32'h439d37e3},
  {32'h443ed16d, 32'hc3cdb640, 32'hc44a28d4},
  {32'hc4365ebd, 32'hc380f3e0, 32'h42d53c62},
  {32'h44316f53, 32'h416e1678, 32'hc2bb5ca2},
  {32'hc4c7ff6c, 32'h4304f75a, 32'hc378c4d6},
  {32'h447b0517, 32'h438c303c, 32'h43968502},
  {32'hc502a32f, 32'h42c4f783, 32'hc238f3aa},
  {32'h44886f8d, 32'h42943612, 32'hc356672e},
  {32'hc4f137c5, 32'h41ffcfb8, 32'h43bb9565},
  {32'h4488f9be, 32'h42eb33d6, 32'hc30cb8a4},
  {32'hc4696502, 32'h436ddcfe, 32'hc35d1662},
  {32'h40e8c900, 32'hc3b1dbaa, 32'h40bd7a35},
  {32'hc4373fe3, 32'h423d3ba0, 32'h437d2b4e},
  {32'h4484d0b1, 32'hc3a33b52, 32'h425fa0cc},
  {32'h4329eb20, 32'hc3c1a68a, 32'hc3986cbf},
  {32'hc47245c9, 32'h41fc5066, 32'h436ef73c},
  {32'h44ba030d, 32'h42899cb8, 32'hc21fcbb9},
  {32'hc3907db0, 32'hc29bb6fa, 32'h43a18982},
  {32'h44741c02, 32'hc34bbfa6, 32'hc188d194},
  {32'hc49c0fb8, 32'hc3051147, 32'h427cf185},
  {32'h45044354, 32'h436945dd, 32'hc21f502c},
  {32'hc4816fdf, 32'h437a00f7, 32'h42c06b95},
  {32'h44bb87f8, 32'h43101b35, 32'hc324262d},
  {32'hc4e4adbc, 32'h432ffbe1, 32'h433a850c},
  {32'h44c9b520, 32'h4291d50e, 32'h42529f02},
  {32'hc4135b25, 32'h436dfad3, 32'h435a4c6c},
  {32'h44fc8fa8, 32'h438abf0e, 32'h43ae2ad5},
  {32'hc480cd3a, 32'h438a2305, 32'h413d04ee},
  {32'h45156765, 32'h436135a9, 32'hc390b9f3},
  {32'hc4aa73c2, 32'hc0be26c4, 32'hc32cdf4c},
  {32'h43f7377e, 32'hc385846a, 32'hc28c1822},
  {32'hc429c87c, 32'hc2b8f63e, 32'h4309d722},
  {32'h43e64794, 32'hc3025233, 32'hc3abc658},
  {32'hc4fae388, 32'h43c04fa2, 32'h42ec3931},
  {32'h44bfc6b6, 32'hc0ab0696, 32'hc3a43019},
  {32'hc2c4f300, 32'h43407198, 32'hc3bcc156},
  {32'h44b35ad2, 32'h42850318, 32'hc4005168},
  {32'hc4a94fcd, 32'h4264305d, 32'hc2b56d6e},
  {32'h44ea0f8f, 32'h42c92ec4, 32'h427f8835},
  {32'hc3394eb8, 32'h42df12e6, 32'h43a0946f},
  {32'h4516875c, 32'h419c4b8a, 32'hc3576d61},
  {32'hc3d09464, 32'h43998c9e, 32'hc3067518},
  {32'h44ef77d3, 32'hc3c003e7, 32'hc34854fb},
  {32'h41beb680, 32'h42a79ed4, 32'hc330cb19},
  {32'h4508218d, 32'h42e97490, 32'h425c3a7b},
  {32'hc4f29051, 32'h41b36dc1, 32'hc2ac20ab},
  {32'h4456cf28, 32'hc2dcba78, 32'h4308fd6f},
  {32'hc4ba9754, 32'h43695e62, 32'hc2fd9243},
  {32'h442dfd3e, 32'h432ada05, 32'hc3c80c3a},
  {32'hc4a38950, 32'hc33bed8d, 32'hc30f17aa},
  {32'h44421686, 32'hc0063288, 32'hc25abd08},
  {32'hc406816b, 32'h42db1a28, 32'h42fef1ab},
  {32'h44910f6d, 32'hc2fc1c7e, 32'h42976f01},
  {32'hc4481639, 32'h42cab9d9, 32'hc3ede91d},
  {32'h44a242a9, 32'h433dafdc, 32'hc370e5ef},
  {32'hc4f3161e, 32'h416b71f9, 32'hc37a4946},
  {32'h437914a0, 32'hc4130cf7, 32'h437713b3},
  {32'hc4625015, 32'hc24a898a, 32'h43df3c81},
  {32'h44af4895, 32'hc37e9652, 32'h42c04cde},
  {32'hc3065116, 32'h428e8126, 32'h4356079d},
  {32'h44fe426f, 32'hc2b23a1d, 32'h42f588dd},
  {32'hc50fc9ea, 32'hc2c8a750, 32'h4399b4c1},
  {32'h44c8c220, 32'h4326a15e, 32'h429a187e},
  {32'hc4827351, 32'h4339e755, 32'h43877980},
  {32'h448267af, 32'hc24e33c0, 32'h426d9c1b},
  {32'hc5127b5c, 32'hc334066e, 32'hc1f59370},
  {32'h4472eb30, 32'hc2975c4a, 32'hc331cc0c},
  {32'hc4b82684, 32'h42cfbb94, 32'h42db2d0d},
  {32'h45089ab8, 32'h43a244a4, 32'hc0c2759f},
  {32'hc4e4a3d2, 32'h43b84cb0, 32'hc38559e8},
  {32'h44da1bd2, 32'h42dd2e85, 32'hc2a85010},
  {32'h43004e10, 32'h42054f08, 32'hc3859e34},
  {32'h44d3686a, 32'hc3062c7f, 32'h41b59b76},
  {32'hc435e7c8, 32'h43b06ca8, 32'h42c4dc14},
  {32'h40372400, 32'h42bdcd20, 32'hc3af74fb},
  {32'hc4fc7f19, 32'hc3a744ff, 32'hc34cae28},
  {32'h43bffb50, 32'hc017c5a4, 32'h43b0b79f},
  {32'hc43e6938, 32'h4352a369, 32'h437bbd7f},
  {32'h449a9681, 32'h439cf4e5, 32'hc275e93b},
  {32'hc4ace0b1, 32'hc3972ffb, 32'h439c0f85},
  {32'h450f9158, 32'h4262a04d, 32'hc3c5eddd},
  {32'hc3a0e379, 32'h41ac360e, 32'hc2ed9af8},
  {32'h436effa4, 32'h4371896d, 32'hc32f1d35},
  {32'hc4af44b2, 32'h430de55c, 32'hc3049801},
  {32'h44d10891, 32'h423789be, 32'hc1f6062f},
  {32'hc488d6f1, 32'hc394a8f3, 32'h42977c8e},
  {32'h4442fd9c, 32'h43dae6c8, 32'h4386e2f6},
  {32'hc487885b, 32'h42c86deb, 32'hc2ea54a7},
  {32'h446548a2, 32'h43691275, 32'h41eb9014},
  {32'hc4c7ef76, 32'h439c3c59, 32'hc1dad968},
  {32'h451a091b, 32'hc119b065, 32'hc2aa204c},
  {32'hc48daf9c, 32'h42cf11bb, 32'hc35843e5},
  {32'h451ce271, 32'hc062a8b8, 32'h42043f01},
  {32'hc40c6806, 32'hc24b5d2a, 32'h4364949b},
  {32'h4510413e, 32'h4112e899, 32'hc2c5c189},
  {32'hc4c9e8dc, 32'h4387ddc2, 32'hc2e9b284},
  {32'h441cade6, 32'hc29b202c, 32'hc2120e8a},
  {32'hc4eaf0ec, 32'h42d4347c, 32'hc3914604},
  {32'h4444dac0, 32'h42132033, 32'h429a49b7},
  {32'hc42c38c4, 32'hc2d4a50e, 32'h4296008e},
  {32'h44d3521b, 32'hc1c5e796, 32'hc39920f3},
  {32'hc492c8cf, 32'hc19a3041, 32'hc3917346},
  {32'h44cc6a94, 32'hc0932190, 32'h42700260},
  {32'hc491f0a0, 32'h4368f337, 32'hc1ea830c},
  {32'h440300c5, 32'h42c0022f, 32'hc2ef65cf},
  {32'hc4e3a72a, 32'hc29510b8, 32'h4386cf85},
  {32'h450bab77, 32'h4256fc70, 32'h43936785},
  {32'hc47d31fc, 32'h4357f871, 32'hc357ae50},
  {32'h45137d81, 32'hc3ab4566, 32'h41e1061c},
  {32'hc4bf3bdc, 32'hc361d146, 32'h43c010b0},
  {32'h4502e438, 32'h4167d332, 32'h3e87e9c7},
  {32'hc45cd14f, 32'hc29bd6af, 32'hc1f47668},
  {32'h4476c4fb, 32'h43929a9b, 32'h419b77ea},
  {32'hc4824218, 32'hc29e35bf, 32'hc2f9e841},
  {32'h446d8bda, 32'hc308a6c0, 32'h419461ac},
  {32'hc4e71781, 32'hc3879eae, 32'h4266590f},
  {32'h44b3ba59, 32'hc12fde7a, 32'hc380e043},
  {32'hc4a48d04, 32'h43a86a33, 32'h4388638b},
  {32'h4434c74c, 32'h43230074, 32'h43dc1dee},
  {32'hc48236c8, 32'h42ba0300, 32'h43926284},
  {32'h44e753fc, 32'h4361fa70, 32'hc342eb93},
  {32'hc4e59c1a, 32'h4259d581, 32'hc28c28f3},
  {32'h43d6889e, 32'hc3c9ef08, 32'hc38fd1e5},
  {32'hc4f44cf4, 32'h4290c331, 32'hc2e78a87},
  {32'h448c4cb6, 32'h434047d1, 32'h42f8beb8},
  {32'hc49cebaf, 32'h4208077c, 32'h43022d10},
  {32'h43a33802, 32'h43db26bb, 32'hc2b395af},
  {32'hc416b17d, 32'h42c9ea38, 32'h435dfe07},
  {32'h440a1b1e, 32'hc2eaf2fb, 32'h438289da},
  {32'hc4c77810, 32'h438d293f, 32'h43248b64},
  {32'h43bb013a, 32'hc2875b44, 32'h43e2d38f},
  {32'hc4728f0a, 32'h428ca7e0, 32'hc3f081be},
  {32'h44b602eb, 32'h4361a43e, 32'hc30cd7a2},
  {32'hc4f6271b, 32'h4365c3c3, 32'h437e8430},
  {32'h44f53078, 32'hc2bd0b7a, 32'h42b4404f},
  {32'h41b6bea0, 32'hc1aa3445, 32'h440cc01a},
  {32'h44f369fb, 32'hc32470db, 32'h41ee3cdf},
  {32'hc4ecbb22, 32'h434b68d6, 32'h43aa251b},
  {32'h44f8162d, 32'h43fc60c1, 32'hc254d068},
  {32'hc500ef7b, 32'hc175064d, 32'hc2227546},
  {32'h44942f74, 32'hc2e543b1, 32'h42131c24},
  {32'hc4ae3ec9, 32'h42ebc026, 32'hc3ee512a},
  {32'h44ba1b49, 32'hc2dfe0b3, 32'hc38402d7},
  {32'hc4d6b0e4, 32'h432bc3e1, 32'hc3293009},
  {32'h446f635d, 32'hc3ef0009, 32'h43d7d3c0},
  {32'hc427d634, 32'h441eed9b, 32'h429e088b},
  {32'h44d6da24, 32'h3f4b83d0, 32'h42d95d61},
  {32'hc3ec810e, 32'h422d49a4, 32'hc1e4841b},
  {32'h449b18be, 32'h42ca3f12, 32'hc35e0697},
  {32'hc49fb45d, 32'hc3bff328, 32'hc375427f},
  {32'h4395f9b2, 32'h42682b8a, 32'hc31ae667},
  {32'hc49b5da5, 32'hc392d93c, 32'hc1e8ef2c},
  {32'h44f893bf, 32'hc3b28fe9, 32'h436cd94a},
  {32'hc45c5a45, 32'h43b15b3c, 32'h43a513b7},
  {32'h4417798e, 32'h431cb222, 32'h42f228bc},
  {32'hc208a3c0, 32'hc381bd97, 32'hc3a6df50},
  {32'h428936a0, 32'h4391ff5c, 32'hc3104ba9},
  {32'hc4da1c8c, 32'hc2a79353, 32'hc1a5c371},
  {32'h44c7c2ea, 32'h43922fd4, 32'h42385872},
  {32'h42b02730, 32'hc24f15c9, 32'hc18b5554},
  {32'h44c77c98, 32'hc0a595bc, 32'hc207762b},
  {32'hc499a8ad, 32'h43221982, 32'hc38e89ac},
  {32'h43e66671, 32'hc34e1958, 32'h42830bac},
  {32'hc45f1ba4, 32'h41da456b, 32'hc2f22682},
  {32'h44687891, 32'h43c208b3, 32'h4225b8a8},
  {32'hc47a5f39, 32'h429640dc, 32'h4310bce1},
  {32'h44fd77ec, 32'hc2f85f14, 32'hc1b657ac},
  {32'hc4bb7210, 32'h428fe008, 32'hc2adff19},
  {32'h438745ac, 32'h439aa5ef, 32'h429c1593},
  {32'hc3f85374, 32'hc35bce68, 32'h42e1a813},
  {32'h45119c1e, 32'hc3063062, 32'hc20c9a03},
  {32'hc4a12dc4, 32'hc382d2c4, 32'h409ce8c0},
  {32'h44b0d61a, 32'hc20cf39e, 32'h43236afe},
  {32'hc48c767a, 32'h437731e3, 32'h43852a39},
  {32'h44f9e331, 32'h42915b54, 32'h434b9d3f},
  {32'hc365cdfc, 32'h4311d4e8, 32'h43649aee},
  {32'h44624819, 32'hc307983d, 32'h42c3e3c4},
  {32'hc4709b64, 32'h425832a6, 32'hc306ce5c},
  {32'h438f3b49, 32'hc2b4133c, 32'hc2250464},
  {32'hc4a16b78, 32'hc1c06524, 32'hc33b44e7},
  {32'h45140a16, 32'hc38c0aec, 32'hc2de451c},
  {32'hc45dce4e, 32'h436ba76a, 32'h431399f2},
  {32'h44d95c7f, 32'hc2d44ecd, 32'hc2eaf644},
  {32'hc4c6a287, 32'h437000f5, 32'h440a368f},
  {32'h44a3db58, 32'h43635f09, 32'hc39ee206},
  {32'hc30e743f, 32'h431bf29a, 32'h43c540da},
  {32'h442c9c98, 32'h4216540b, 32'hc261db0b},
  {32'hc4eb4207, 32'h43e6e962, 32'hc3337621},
  {32'h43de0fa5, 32'hc3b8514f, 32'hc4115acf},
  {32'hc4c54112, 32'h408c5854, 32'h433ff6c3},
  {32'hc32925fd, 32'h430842c6, 32'h4390805e},
  {32'hc4cd3aa5, 32'h43157e39, 32'hc23c24da},
  {32'h448c28f4, 32'h42e66875, 32'hc1f447a7},
  {32'hc4b42074, 32'h4312267c, 32'h42efd113},
  {32'h4426c018, 32'h4355741e, 32'hc342aba3},
  {32'hc4d44416, 32'hc334d20e, 32'hc11d07bf},
  {32'h447a33fe, 32'h42226bdb, 32'h4141b639},
  {32'hc40de40c, 32'h41f1663a, 32'hc1d0a8a1},
  {32'h44585951, 32'hc2f5c3d7, 32'hc2a53995},
  {32'hc4ad2fc8, 32'hc3450e58, 32'hc2414f37},
  {32'h44e25ff9, 32'hc2c4ebd8, 32'h43ce44c7},
  {32'hc3c67a74, 32'h3f30c02e, 32'hc3f2360c},
  {32'h43c53062, 32'hc33e9a36, 32'h43e371c0},
  {32'hc4c5dcc6, 32'hc2dffd3f, 32'hc39c4624},
  {32'h44323510, 32'h41d2a79c, 32'h439cbf90},
  {32'hc4ccb5f2, 32'hc4284584, 32'hc2c24141},
  {32'h44f1fda2, 32'hc21970b2, 32'hc2944145},
  {32'hc5099e6f, 32'h42b86da5, 32'hc3c46cda},
  {32'h429c5c82, 32'h42660184, 32'hc387990d},
  {32'h42700e80, 32'hc3ecc64a, 32'h42bbed7c},
  {32'h44ce5376, 32'h430f58e6, 32'hc331d973},
  {32'hc4359907, 32'hc25bfeb5, 32'h4259d7ef},
  {32'h44c7895d, 32'h43200b00, 32'h43bb6fff},
  {32'hc4942076, 32'h42504c68, 32'hc16eb978},
  {32'h447ece29, 32'h4321017f, 32'hc3f4a86e},
  {32'hc4a2b590, 32'h418c26ea, 32'h4252608d},
  {32'h45003cf0, 32'h436b423c, 32'hc3b2015b},
  {32'hc5014953, 32'hc2870f33, 32'hc25b0bac},
  {32'h44e97c73, 32'hc2e8546f, 32'hc3a634d3},
  {32'hc51510e6, 32'hc3e8e8f3, 32'h42a4ca1a},
  {32'h44f78c84, 32'hc2049c8c, 32'hc00f6514},
  {32'hc469fdf9, 32'hc3beb844, 32'hc21fc166},
  {32'hc397fa12, 32'hc32871d5, 32'hc22c4b59},
  {32'hc5086a59, 32'h43004c72, 32'h4340654d},
  {32'h44e879f6, 32'hc24e3f13, 32'hc39fb4b2},
  {32'hc44ba5f4, 32'hc383b45a, 32'hc2eee095},
  {32'h44c5a41f, 32'hc3864ac6, 32'h440bd02b},
  {32'hc4e7e2d4, 32'hc37bc7c7, 32'hc4058488},
  {32'h440eedd7, 32'h432110e5, 32'h43902e3c},
  {32'hc4da9098, 32'hc33ae43b, 32'h43d33392},
  {32'h4488dfbe, 32'h438630a0, 32'hc3567cc2},
  {32'hc4ff8e14, 32'h42cb3d27, 32'h433fd03b},
  {32'h4457c310, 32'hc26ac833, 32'h43ad8e71},
  {32'hc506ffe0, 32'hc26f7dd0, 32'h42a646ae},
  {32'h452345d0, 32'h43602750, 32'h431c9514},
  {32'hc5015300, 32'hc26c7d70, 32'h41ce03a6},
  {32'h450ae44c, 32'h4027f0c6, 32'hc405a2ef},
  {32'hc364359d, 32'h4361573e, 32'hc3e137e2},
  {32'h44d02891, 32'h435cc2c7, 32'hc3bc9eef},
  {32'hc41853ab, 32'h433cf846, 32'h43a0f2dd},
  {32'h44fca0ea, 32'h3f344b50, 32'h421de862},
  {32'hc4c8ab80, 32'h42d05a63, 32'hc35beaba},
  {32'h44c3aa10, 32'hc38a18bb, 32'h42394e39},
  {32'hc4b2e027, 32'h439fbf8c, 32'hc2acf177},
  {32'h44912037, 32'hc30d9f38, 32'hc31f623d},
  {32'hc2a73660, 32'h4351dfd4, 32'h433ceaca},
  {32'h450974f3, 32'hc3dc1ec6, 32'hc08b5fd8},
  {32'hc4cc165a, 32'hc33cb80d, 32'h431499cc},
  {32'h445030f2, 32'h435b3756, 32'hc335903d},
  {32'hc508f07b, 32'h4370eea1, 32'hc2945aa1},
  {32'h442329ee, 32'hc39933da, 32'hc1742faa},
  {32'hc4b0cae8, 32'hc2415a15, 32'hc28d0502},
  {32'h451019a3, 32'hc4193c39, 32'hc3b6ec2a},
  {32'hc5059402, 32'h4207f7f8, 32'h438c4c05},
  {32'h44fbbca7, 32'h431e7c0d, 32'hc3c924ac},
  {32'hc4f19a2e, 32'h43b006d6, 32'hc2b30e1f},
  {32'h4458d513, 32'h41c82589, 32'h4343e8e0},
  {32'hc4ce41a3, 32'h420e7586, 32'h4425a505},
  {32'h44dc4004, 32'hc2a38050, 32'h4338ded7},
  {32'hc236ade2, 32'h43039dd2, 32'h433c4c1e},
  {32'h442fd6c4, 32'h43cb52db, 32'hc2185d08},
  {32'hc49eddb9, 32'hc41deb3e, 32'h4309f5c0},
  {32'h45002e5c, 32'h435276f7, 32'hc389d5d9},
  {32'hc488d21a, 32'h430bfe7b, 32'hc32462c3},
  {32'h44597d0f, 32'h41a0ad38, 32'h428be78e},
  {32'hc46b4b44, 32'h4206e7cd, 32'h42976ab9},
  {32'h44fb34ea, 32'h440d6f84, 32'h42fde986},
  {32'hc2a35a3f, 32'hc21c2f82, 32'h43659223},
  {32'h45001b50, 32'hc3616001, 32'hc385d88a},
  {32'hc3a4931f, 32'hc329397d, 32'hc38d69c2},
  {32'h447e38f1, 32'hc382a064, 32'hc287cba3},
  {32'hc3d18588, 32'h407e7723, 32'hc0b58b7e},
  {32'h44ceccd0, 32'hc38c4a00, 32'hc23272ce},
  {32'hc4c07703, 32'h42dc55d8, 32'hc20d5cd6},
  {32'h44f1b766, 32'h42eef356, 32'h43a3bd9e},
  {32'hc4bfea1e, 32'hc344acd6, 32'hc29ccc3a},
  {32'h450238b2, 32'h43488775, 32'h4297d5ac},
  {32'hc4442ad9, 32'h43fc4059, 32'hc21b18fe},
  {32'h444f5962, 32'hc3b45a6d, 32'h43adf1a1},
  {32'hc507c634, 32'h44358461, 32'h41067482},
  {32'h445ee518, 32'hc369dd5d, 32'hc2dd9198},
  {32'hc3d49911, 32'hc32d1823, 32'h43c84d16},
  {32'h44becb12, 32'hc38742cd, 32'hc296463b},
  {32'hc1a69180, 32'h42c05864, 32'h42c75d5a},
  {32'hc28f7470, 32'h42ceb24a, 32'hc3c80f3e},
  {32'hc44ef267, 32'hc2dd8ebd, 32'h43ca03c4},
  {32'h4464b4a6, 32'hc30a04dc, 32'hc38c2f5b},
  {32'hc4ad76bd, 32'h4277e372, 32'h434081ac},
  {32'h444ec970, 32'hc368d308, 32'hc1343518},
  {32'hc3e25915, 32'hc3fd5a8e, 32'h4392ad10},
  {32'h44d2bbe2, 32'h435cf82b, 32'h3e2c7f80},
  {32'hc414af4f, 32'hc381df21, 32'h43bec799},
  {32'h451b5d4d, 32'hc3611108, 32'h43871d0d},
  {32'hc43d7702, 32'hc2b759f5, 32'h4236848b},
  {32'h44948abb, 32'hc2dab2f6, 32'hc35fe3a3},
  {32'hc4bb481a, 32'h42f13620, 32'hc237f240},
  {32'h446d5eaa, 32'h43db72d5, 32'h431dab71},
  {32'hc496e2cc, 32'h440624a4, 32'hc160401e},
  {32'h44f1b21e, 32'hc2aa1b67, 32'h4215ffd1},
  {32'hc41b7626, 32'hc38b2e4d, 32'hc1e26e23},
  {32'h440e00e1, 32'hc2f81c27, 32'h439fb06c},
  {32'h430a6158, 32'hc3866d3c, 32'hc25b902b},
  {32'h4440756a, 32'h41b9d7c2, 32'h438b126e},
  {32'hc42bd1b6, 32'hc1cbd778, 32'hc34dcaee},
  {32'h446b3df1, 32'hc3b13fd5, 32'hc390a1c2},
  {32'hc3e03836, 32'h43a0be8d, 32'h431a820d},
  {32'h44c9265a, 32'hc2975afd, 32'hc27aecfe},
  {32'hc492f687, 32'h4389b168, 32'hc36ee04c},
  {32'h4491d218, 32'h426f3e7b, 32'hc390d12e},
  {32'hc486ad26, 32'h42fed092, 32'hc2246d40},
  {32'h441672ac, 32'h4292aa7b, 32'hc20eec00},
  {32'h4202e6f6, 32'hc3582c18, 32'h4313a4ce},
  {32'hc07c3e00, 32'h430874be, 32'h436fea2d},
  {32'hc25a6fc0, 32'hc314cba8, 32'h437f607c},
  {32'h44b66f90, 32'h42b801bf, 32'hc3aa92e2},
  {32'hc40d632c, 32'hc4050900, 32'h415b0614},
  {32'h44e0a183, 32'hc1c814b9, 32'hc1fb6459},
  {32'hc4ace362, 32'hc208e7a8, 32'hc32d9069},
  {32'h44e27e9d, 32'hc207f6db, 32'hc393141f},
  {32'hc4c90eba, 32'hc38978f5, 32'h42dbda05},
  {32'h4505ac26, 32'hc019c099, 32'hc3b299dc},
  {32'hc513cb67, 32'hc37708a6, 32'hc438fe6d},
  {32'h43ce0858, 32'hc37a6282, 32'h43344551},
  {32'hc4e5b53e, 32'hc35a87ba, 32'h42ec350c},
  {32'h44d7d2e0, 32'h42bf505e, 32'h4127f692},
  {32'hc48012a8, 32'h41b46d2b, 32'h430ac822},
  {32'h445a5199, 32'h43085594, 32'h4390f649},
  {32'hc3539d80, 32'hc32caf12, 32'h435f4c9d},
  {32'h44a4fad0, 32'h43020087, 32'hc2286ded},
  {32'hc4d35cdb, 32'h42b0db94, 32'hc2c492f0},
  {32'h44ab6f53, 32'hc2a296af, 32'hc25eeadf},
  {32'hc3df68f8, 32'h410822e6, 32'hc247eee2},
  {32'h44b69712, 32'h422be18b, 32'hc2dd0eda},
  {32'hc449f900, 32'hc35858f0, 32'hc200f87c},
  {32'h44b440fa, 32'hc356ffda, 32'hc33882a3},
  {32'h423c7781, 32'hc2fa2cf6, 32'hc3d6330f},
  {32'h44ea2225, 32'hc33d252c, 32'h4308c561},
  {32'hc481e4e4, 32'hc3ae0276, 32'hc3e186c2},
  {32'h44d4c505, 32'hc33b3031, 32'h431d8ef0},
  {32'hc4fd080c, 32'h4379e4f8, 32'h4277ea63},
  {32'h44fed4c0, 32'h433a6de1, 32'h42df37ef},
  {32'hc4ab2ca3, 32'hc307ebdb, 32'h4259f31c},
  {32'h440e0402, 32'hc2cc9530, 32'hc380d52c},
  {32'hc4a253bb, 32'h438c5c7a, 32'hc31a649e},
  {32'h44839267, 32'hc3af8027, 32'hc2972ef6},
  {32'hc510e3b4, 32'h435717ec, 32'h3f955897},
  {32'h440df766, 32'h428c6a68, 32'hc3e2b840},
  {32'hc29c9cd8, 32'hc3d5b0ac, 32'h4308d2ad},
  {32'hc3df4c0e, 32'hc3188bf7, 32'hc4277ad8},
  {32'hc4fe9337, 32'h41e87596, 32'hc2901e81},
  {32'h4499e3fb, 32'hc396b82a, 32'hc331a5b5},
  {32'hc4fd3c86, 32'h420e6fa9, 32'hc35547df},
  {32'h44bb20f4, 32'h43366eec, 32'hc36db8ff},
  {32'hc3f2ca54, 32'h42d0cbc0, 32'hc3b85626},
  {32'h44d5db62, 32'hc3473712, 32'h4377e328},
  {32'hc3f025b4, 32'hc1a57030, 32'hc4113a6b},
  {32'h44eea050, 32'hc3461b28, 32'h43bc98ae},
  {32'hc4f66614, 32'h426ac2e7, 32'hc2a4a798},
  {32'h448085fc, 32'h43b00cda, 32'hc3b1b6e4},
  {32'hc3307684, 32'h43d4b875, 32'h430615ca},
  {32'h450f7504, 32'hc331c6bb, 32'h434ef49a},
  {32'hc3daebe8, 32'h437dcd79, 32'h42b9a2e5},
  {32'h44815f6a, 32'hc3660ca0, 32'hc36cadab},
  {32'hc39cc4b0, 32'hc31d139f, 32'h43234c23},
  {32'h43ff887e, 32'h4352eb2a, 32'hc20e9315},
  {32'hc300dd80, 32'hc3d6cdd0, 32'h4317753d},
  {32'h45184560, 32'h41c6d6f2, 32'hc1f08644},
  {32'hc4208008, 32'h43457ec0, 32'hc3716a89},
  {32'h443a237d, 32'hc38491fb, 32'h4260d8b0},
  {32'h41a88605, 32'hc3314add, 32'hc234c8f9},
  {32'h449bb4cb, 32'hc2ae2df2, 32'h434c1cd6},
  {32'h435419a0, 32'hc2fb2947, 32'h425df181},
  {32'h44c9ac7c, 32'h432915e0, 32'h42a9f8ef},
  {32'hc4af740f, 32'hc2b368ac, 32'h419a272f},
  {32'h44d77fd5, 32'h4307c6c0, 32'h420b4c35},
  {32'hc3f2aa48, 32'h438abfde, 32'hc02e20e0},
  {32'h44eb7457, 32'hc1af8a7e, 32'h4388a245},
  {32'hc49194ec, 32'h42fbe0cd, 32'h42e7479d},
  {32'h43b4aa65, 32'h43b4cb0c, 32'h3f5f4dd8},
  {32'hc3ad2c14, 32'h43319d52, 32'hc373a5fa},
  {32'h44bce9a8, 32'h4397ff60, 32'hc3aba5bc},
  {32'hc510fc96, 32'hc35673df, 32'h4281f028},
  {32'h451e441f, 32'hc271b4d3, 32'h432bf191},
  {32'hc4d65336, 32'hc2b05608, 32'h43b87a36},
  {32'h4510778a, 32'h4249cc9e, 32'h42d2324c},
  {32'hc481f32c, 32'h434af3a4, 32'h431cc39d},
  {32'h441ba340, 32'hc2be4757, 32'h4312c2c1},
  {32'hc4b767d1, 32'h426ed162, 32'h43620804},
  {32'h44c1f556, 32'hc3f9a141, 32'h43374f7c},
  {32'hc2f45d20, 32'hc334246c, 32'h432e0807},
  {32'h4444a638, 32'hc1829264, 32'h424dfb9d},
  {32'hc4c9f79c, 32'hc34bd175, 32'hc31bc2e8},
  {32'h449d9344, 32'hc15b0802, 32'h43925104},
  {32'hc50e8907, 32'hc39e14d6, 32'hc30fc055},
  {32'h448d6f81, 32'h42f5535a, 32'h43a8f5bf},
  {32'hc4d88cdc, 32'h43c6f1d6, 32'hc36b33e1},
  {32'h44baad85, 32'h42b75732, 32'hc40f252c},
  {32'h439236b0, 32'h42d15a8d, 32'h437f0584},
  {32'h43c98b54, 32'h4389e6e0, 32'h42ce088a},
  {32'hc5097d0a, 32'h432e5d9f, 32'h41c6eb06},
  {32'h450b4d66, 32'hc2ff7412, 32'hc3199336},
  {32'hc456305c, 32'hc3579f46, 32'h43349a28},
  {32'h4512d216, 32'h432f3bb0, 32'hc3565ab2},
  {32'hc4a6c620, 32'h430999d7, 32'hc381939d},
  {32'h44c62551, 32'hc3ba2dac, 32'hc375f1e6},
  {32'hc50eb9e0, 32'hc32ec2a0, 32'h43ec4a2e},
  {32'h4404d775, 32'h433d136d, 32'hc3a99af2},
  {32'hc4699607, 32'hc3540f4a, 32'h4365bef3},
  {32'h43a97ccf, 32'hc2e02acf, 32'hc2ed52b8},
  {32'hc3d925c8, 32'hc370e587, 32'hc22f1e6f},
  {32'h43a77194, 32'hc3ae8403, 32'h431fe51e},
  {32'hc4448eac, 32'h43203d54, 32'h4307fab5},
  {32'h43c6e1d4, 32'h4237d8ab, 32'hc2ce912e},
  {32'hc3b223c8, 32'h4345035e, 32'hc33adc3f},
  {32'h4411ce32, 32'hc2ab1838, 32'h42cf4596},
  {32'hc3c2dd47, 32'hc2e8a89d, 32'hc353e74d},
  {32'h448f0311, 32'hc3af60b6, 32'h43f9ebdf},
  {32'hc4669f5a, 32'hc3238e91, 32'h43002918},
  {32'h4449fbd4, 32'h4369467f, 32'h4387c4d6},
  {32'hc3ce571a, 32'hc3c96f9a, 32'hc2d72fb6},
  {32'h434e515a, 32'h429d1340, 32'h437abd5a},
  {32'hc42e9874, 32'hc22b1825, 32'h43835f01},
  {32'h44a1baae, 32'h42313605, 32'h43887933},
  {32'hc4b90059, 32'h4385873c, 32'hc32a094c},
  {32'h45007207, 32'hc37ed637, 32'h439bac15},
  {32'hc4912c8a, 32'h41d11bf7, 32'hc39127c8},
  {32'h44b988e9, 32'hc2d71767, 32'hc2128821},
  {32'hc3576640, 32'hc30ffc9f, 32'hc1a8f39e},
  {32'h43db8964, 32'hc2327a9b, 32'h434fadab},
  {32'hc50a1cb9, 32'hc2d9f8ce, 32'h40372a10},
  {32'hc1db3600, 32'h42603f9e, 32'h434c58aa},
  {32'hc486592f, 32'h431efe67, 32'h42426c4a},
  {32'h4504d323, 32'hc3713141, 32'h439e7a14},
  {32'hc4136870, 32'hc3e63ccf, 32'h4289f885},
  {32'h44b28f41, 32'h43ff3a43, 32'h425132a8},
  {32'hc2e2847e, 32'hc2017743, 32'hc2e7fb0e},
  {32'h44932776, 32'hc3da5fb7, 32'h427ba39e},
  {32'hc50a5ba0, 32'h429915fc, 32'hc2b2c8c7},
  {32'h4445fe76, 32'h42a34740, 32'h4162ae02},
  {32'hc467cc46, 32'h42d40110, 32'hc38c25d4},
  {32'h444c3d7c, 32'hc315f1dc, 32'h43633621},
  {32'hc3d2f7c7, 32'hc32e1545, 32'hc3047840},
  {32'h44c9490a, 32'hc3122d97, 32'h42361876},
  {32'hc4c21150, 32'h4330c8cb, 32'h43d9e069},
  {32'h43ea306e, 32'h43de4eff, 32'h431c1bb9},
  {32'hc4e57326, 32'hc35d2f3e, 32'hc322938c},
  {32'hc479b0ca, 32'hc2ec0983, 32'hc33759a6},
  {32'h44c43534, 32'h43d4ebc0, 32'h42e0dddc},
  {32'hc4bcb204, 32'hc213cfdc, 32'hc43d6c20},
  {32'h44e9896f, 32'hc3a25f02, 32'h438553eb},
  {32'hc40fa38e, 32'hc324182b, 32'hc362c1d2},
  {32'h44c7330c, 32'h41122e08, 32'hc390901d},
  {32'hc453faf7, 32'h4399785d, 32'hc396fa13},
  {32'h4483cf7e, 32'h4316cdd9, 32'hc2aa3aef},
  {32'hc4c91d88, 32'h42513c0a, 32'hc2e284f1},
  {32'h44d9a28e, 32'h43123d9b, 32'hc3ba4225},
  {32'hc4e9675e, 32'h4262dc6e, 32'hc290e50f},
  {32'h4481c089, 32'hc1a43462, 32'hc2967f10},
  {32'hc45c1388, 32'h43fb5fa7, 32'hbfd529e0},
  {32'h452369d5, 32'hc295c66f, 32'hc26b0e7a},
  {32'hc4adc437, 32'hc2bcd822, 32'hc319cfcd},
  {32'hc28fc245, 32'hbf921bf3, 32'h4311cf53},
  {32'hc4f479eb, 32'hc28237bc, 32'hc36d8939},
  {32'h4421beec, 32'h43214083, 32'h42a76713},
  {32'hc5106e76, 32'h42f53eb1, 32'hc28c0620},
  {32'h45076a8c, 32'h43c1601a, 32'h425f4dd0},
  {32'hc4dff372, 32'hc31ff8fc, 32'h428b403d},
  {32'h44845c88, 32'h423a2fb7, 32'hc1d51b66},
  {32'hc50b10af, 32'hc2925e8e, 32'hc2beb622},
  {32'h45071b2e, 32'hc3ba589b, 32'hc3368a11},
  {32'hc4cecdc4, 32'hc2d504ca, 32'h42e1fa30},
  {32'h43f45c47, 32'hc3cf5c74, 32'h437a504a},
  {32'hc500f577, 32'h416fe476, 32'hc31e38aa},
  {32'h442f38ac, 32'h4299aa91, 32'h43588968},
  {32'h3ffc8362, 32'h4383c884, 32'hc3c2d85a},
  {32'h4487c58d, 32'h43ae0be0, 32'hc283adeb},
  {32'hc4d381cd, 32'h430b4198, 32'h43af96ac},
  {32'h4409b86b, 32'hc34e998e, 32'h4322e942},
  {32'hc4cacaa6, 32'h428dfbbc, 32'hc3af44d8},
  {32'hc2aacdf0, 32'hc3fd614d, 32'hc241c622},
  {32'hc4120ef4, 32'hc3e8e414, 32'hc38016d7},
  {32'h42020160, 32'hc3509cca, 32'hc32028e2},
  {32'hc41466e0, 32'hc35a806d, 32'h43b78c6f},
  {32'h441eff54, 32'h438dfd6c, 32'hc38469dd},
  {32'hc49a6e1e, 32'hc21a9b5b, 32'h43476460},
  {32'h43389296, 32'h4297538a, 32'hc308ba57},
  {32'hc4f44e48, 32'h426e31a1, 32'h42c5eec9},
  {32'h44c75631, 32'hc2444812, 32'hc2b487d0},
  {32'hc4ab7236, 32'h4309e07a, 32'hc3ac6d99},
  {32'hc1802760, 32'hc1d8a955, 32'h4366bb23},
  {32'hc40ba336, 32'hc2aebc0a, 32'h420f47ac},
  {32'h44f1576c, 32'hc26dbadc, 32'h43129f05},
  {32'hc45429ac, 32'hc38dc179, 32'hc2fbe960},
  {32'h450f3d87, 32'h414a1735, 32'hc289a01f},
  {32'hc4adbe60, 32'h43a9ad81, 32'h4219ed7d},
  {32'h450be72a, 32'hc2a9a4f1, 32'h433c540c},
  {32'hc4569b34, 32'h42ee73d6, 32'hc401bbd3},
  {32'h43d8c4b8, 32'hc3ceda44, 32'h43960059},
  {32'hc3846188, 32'h427ffc87, 32'hc34091d4},
  {32'h44f93826, 32'hc34609e7, 32'h43b246b3},
  {32'hc44664ca, 32'h42826fcc, 32'hc2810701},
  {32'h44e0a798, 32'h4236119e, 32'hc3205c4e},
  {32'hc4b1376c, 32'hc3b99079, 32'hbfd09b9d},
  {32'h44ffd2f6, 32'h4358cf80, 32'hc3941929},
  {32'hc4d091ea, 32'h43f8cc6f, 32'hc1c76566},
  {32'h440d56a5, 32'hc3a6aba9, 32'h41eef4f9},
  {32'hc2707d00, 32'hc3a07808, 32'hc3581b7f},
  {32'h4405b6c0, 32'h431a6ea0, 32'h429c0d37},
  {32'hc46748b8, 32'h41252c05, 32'hbfaa4797},
  {32'h443ab07e, 32'h431a4c50, 32'h42b73a40},
  {32'h42057748, 32'hc21105b9, 32'h43a79628},
  {32'h448a157b, 32'hc3971161, 32'h42ec9746},
  {32'hc484d9c0, 32'hc28127f2, 32'hc2b351f8},
  {32'h44a8838c, 32'h432c9cbb, 32'h4293e3e9},
  {32'hc51250a1, 32'hc34222d6, 32'h43229f8f},
  {32'h439f9fec, 32'hc3f079db, 32'h43df2233},
  {32'hc47c3f68, 32'hc3391d86, 32'hc1e545a8},
  {32'h4477ca5e, 32'hc308fbaf, 32'h43948953},
  {32'hc4f4bd39, 32'hc36051aa, 32'h42ab58a9},
  {32'h44ec8a24, 32'hc2970db9, 32'h42e36406},
  {32'hc4279403, 32'h411e5b49, 32'hc318120f},
  {32'h440964b1, 32'h436c7900, 32'hc09f0479},
  {32'hc460aa52, 32'h4331582c, 32'hc3869c52},
  {32'h43bc61e4, 32'h427057b6, 32'hc385b8c6},
  {32'hc41af2ac, 32'h4398dfff, 32'h42ae1a85},
  {32'h44a6e751, 32'hc322717c, 32'h43449b16},
  {32'hc43fa2a6, 32'hc3b1285d, 32'h43643929},
  {32'h43985842, 32'hc20a03cb, 32'h43d8497b},
  {32'hc39c6a60, 32'hc3cb9b28, 32'h43a41a64},
  {32'h44ddcf3f, 32'h43e7daf3, 32'hc3a042a7},
  {32'hc4b64c45, 32'h43977fbb, 32'hc2df6d7b},
  {32'h4489a3b5, 32'h4325d376, 32'h42b71596},
  {32'hc492d0cc, 32'h435d8822, 32'hc32cdc78},
  {32'h44244616, 32'hc32a8be9, 32'hc2da13d5},
  {32'hc4d12705, 32'h43770df9, 32'hc3a30af1},
  {32'h44e50a00, 32'h43045344, 32'h43abaac7},
  {32'hc4b127ac, 32'hc3d0e789, 32'hc389f808},
  {32'h43f6384c, 32'hc3a10964, 32'hc31b6a85},
  {32'hc46e0728, 32'h437c8cbe, 32'h4386fc72},
  {32'h43fe3523, 32'hc228e84c, 32'h42581e76},
  {32'hc4ed0998, 32'h434dca7c, 32'hc12e5c1a},
  {32'h44e27abc, 32'hc24b6680, 32'hc27a3bac},
  {32'hc479d332, 32'h40099917, 32'h43f33535},
  {32'h450c19a7, 32'h431c4133, 32'hc2f826ba},
  {32'hc5075190, 32'hc1ead49f, 32'hc38457b5},
  {32'h43aee46a, 32'hc3f7fa5d, 32'h42949471},
  {32'hc483672a, 32'h438201ab, 32'h4286ec90},
  {32'h44d60da6, 32'hc1536bff, 32'h4383832a},
  {32'hc2be2248, 32'h43159f5d, 32'h43aa57e7},
  {32'h44197c9c, 32'hc38ad409, 32'h4413ed26},
  {32'hc3818f98, 32'h42af413e, 32'h4395b88c},
  {32'h44196a8c, 32'h41acaf73, 32'hc36a72d3},
  {32'hc51b1c84, 32'h438579f0, 32'hc35e3a18},
  {32'h43b97c4c, 32'hc2192d46, 32'hc3430940},
  {32'hc5088514, 32'hc39e61fa, 32'h436ad59e},
  {32'hc1605380, 32'h4361fec0, 32'h43a2b21e},
  {32'hc263e297, 32'hc39be6e7, 32'hc3847261},
  {32'h44c5ef0f, 32'h43a93025, 32'h42a44477},
  {32'hc411e6e2, 32'h432b2f78, 32'h42d01945},
  {32'h44e945d0, 32'h415458b2, 32'hc3a6733c},
  {32'hc3a1edb4, 32'h4305e15a, 32'h4349e8f6},
  {32'h449ea2b6, 32'h42e17bc6, 32'hc3e93682},
  {32'hc4fdebe5, 32'h411c2d94, 32'h44246828},
  {32'h435fb220, 32'hc39ba075, 32'hc3701611},
  {32'hc40c5962, 32'h428fb9a8, 32'hc32de49a},
  {32'h4460d5d2, 32'hc19bab98, 32'hc37d5f43},
  {32'hc2baea40, 32'hc320a798, 32'hc1940f5c},
  {32'h44a0f8e7, 32'h42fd32bf, 32'hc3d5b9d9},
  {32'h4317f570, 32'h439b700a, 32'h412ce288},
  {32'h4504369e, 32'h432ac4c6, 32'hc25c7f2a},
  {32'hc41278b6, 32'h43e52f88, 32'h42579668},
  {32'h449baf1a, 32'hc1b14c6b, 32'h435cc6e0},
  {32'hc41706e1, 32'h43872420, 32'hc295c7a5},
  {32'h44338b43, 32'hc2287ffc, 32'hc339aa4e},
  {32'hc4cba8d8, 32'h427d68e0, 32'h439aa656},
  {32'h44824a9b, 32'h43d81494, 32'h43e79359},
  {32'hc3b921fc, 32'hc395e78f, 32'h437b17e5},
  {32'h44d53375, 32'hc2e4fff3, 32'h43650ee3},
  {32'hc508372a, 32'hc3c28614, 32'h42eb0e2b},
  {32'h43fcb6c8, 32'hc33b24e2, 32'hc18c9170},
  {32'hc4889075, 32'h4360a4a7, 32'hc3970ad6},
  {32'h448db646, 32'hc3b42d3e, 32'hc37b22d3},
  {32'hc500c55e, 32'hc365768c, 32'hc27f6aee},
  {32'h44c18409, 32'h4288e5ab, 32'h431beefd},
  {32'hc437d209, 32'hc3279d26, 32'h426e17fb},
  {32'h4444fb6a, 32'h43cf24c3, 32'h422acdf6},
  {32'hc48c4838, 32'hc29ebbd8, 32'hc379dbef},
  {32'h44873761, 32'h414db1bf, 32'h43dda117},
  {32'hc4ee08d7, 32'h43365ca5, 32'h4352e9e0},
  {32'h41ac8bc0, 32'hc34f3597, 32'h42c61866},
  {32'hc2629fc0, 32'h4317ff27, 32'h422c8fd5},
  {32'h44a5b261, 32'hc33e08e5, 32'hc32e8b29},
  {32'hc445d880, 32'hc3ee3f35, 32'hc40cf3ac},
  {32'h44a8da26, 32'hc3295f59, 32'hc313db61},
  {32'hc4ff1c96, 32'h4221ffb5, 32'h438506bc},
  {32'h44b8190c, 32'hc3c1d37d, 32'h440765e9},
  {32'hc49c3d66, 32'h42603cc0, 32'hc3c53372},
  {32'h4481e7a9, 32'h4300e0d9, 32'hc3bd7f5d},
  {32'hc45ee6e7, 32'h42d03561, 32'h41908fcb},
  {32'h44d780fa, 32'h425e1903, 32'hc30293da},
  {32'hc4d183ad, 32'hc28b626d, 32'h430fbeaa},
  {32'h450b14a2, 32'h41eade05, 32'hc3bdf1a5},
  {32'hc45bb2cb, 32'hc3da21b6, 32'hc24663f5},
  {32'h431094e0, 32'hc1dbc4b3, 32'hc401009e},
  {32'hc40c8cdb, 32'hc347c3d5, 32'hc3577302},
  {32'h44aa1fd3, 32'h42cf5364, 32'h41e0bf96},
  {32'hc3db446e, 32'hc31aaa83, 32'hc3b320fe},
  {32'h4363da30, 32'hc35d865a, 32'h435d6449},
  {32'hc4fc255b, 32'h41a3697e, 32'hc2037088},
  {32'h441ce18c, 32'h42b7ba94, 32'h42f7a4a7},
  {32'hc4d59f03, 32'h433a47ba, 32'hc3b98360},
  {32'h44953818, 32'hc28f18f2, 32'hc329e482},
  {32'hc428ff88, 32'h439d9e32, 32'hc28b2dcc},
  {32'h436cc45c, 32'hc35030b6, 32'h42c7525d},
  {32'hc491f3aa, 32'h4399a595, 32'hc327186a},
  {32'h447b1f60, 32'h43876cb5, 32'hc2995f77},
  {32'hc4136996, 32'hc165214c, 32'hc3579c48},
  {32'h44a42f3c, 32'hc36dcc53, 32'hc1a8b8fb},
  {32'hc4c93cd0, 32'hc388647a, 32'hc23a266a},
  {32'h44776524, 32'hc3792ade, 32'h40ab770a},
  {32'hc4b3faa0, 32'hc34030a3, 32'hc26d58a4},
  {32'h448b9e2a, 32'h434183ca, 32'h4175e5e2},
  {32'hc48fe951, 32'h424a2c54, 32'hbee571b0},
  {32'h450eb1e8, 32'h414e6e2a, 32'hc301b197},
  {32'hc4f20c0c, 32'h42f47ae8, 32'h41df879d},
  {32'h43ba16cc, 32'hc3288977, 32'hc329a9e9},
  {32'hc34ba3e8, 32'hc1af8b4f, 32'h43f23c80},
  {32'h4383d854, 32'h43c2fddc, 32'hc2d12e5b},
  {32'hc4a8bafa, 32'hc3cdccdc, 32'hc301480f},
  {32'h4453c6b0, 32'hc367261f, 32'h435620cc},
  {32'hc46a9ac9, 32'hc3dd3d02, 32'h4356834d},
  {32'h44e5c80a, 32'hc2767531, 32'h42f6dde3},
  {32'hc49a5597, 32'hc341ed99, 32'h433f8711},
  {32'h44bc3684, 32'h42e857be, 32'h430d365d},
  {32'hc4549a22, 32'h43e47032, 32'hc0f88214},
  {32'h4503e1e3, 32'hc3574f1e, 32'hc36f22f8},
  {32'hc4dbe581, 32'h431b16be, 32'hc2df1754},
  {32'h44f97887, 32'hc20af9ef, 32'h435e4387},
  {32'hc41180ba, 32'h4302cf3c, 32'hc3868c2b},
  {32'h450a4b40, 32'hc3347265, 32'h43877b6d},
  {32'hc4a697ca, 32'hc24731a0, 32'hc2f4be28},
  {32'h4502f4ff, 32'h431aa2c3, 32'hc303dec5},
  {32'hc24079c0, 32'hc323b8d8, 32'hc131fb8a},
  {32'h4506b639, 32'h43299069, 32'h43e65e12},
  {32'hc49019cb, 32'hc396977d, 32'hc27002b6},
  {32'h44624676, 32'h42319e58, 32'h41b3b61e},
  {32'hc46c3412, 32'h415e2ed1, 32'h4389da69},
  {32'h42a9cbd4, 32'hc2c6beb7, 32'h432e3a44},
  {32'hc4167b24, 32'hc37c3158, 32'h430b8600},
  {32'hc3640612, 32'hc31e90f9, 32'h439c0081},
  {32'hc36e79d8, 32'h4300c0d9, 32'h43a82896},
  {32'h44081854, 32'h43748ba9, 32'h43040139},
  {32'hc5038609, 32'h43d4cfb9, 32'hc34096b2},
  {32'h4394b42c, 32'hc10cda79, 32'hc31c1986},
  {32'hc40f3718, 32'hc33c5564, 32'h434726f7},
  {32'h4507eead, 32'hc37495c0, 32'hc34bdde0},
  {32'hc3fb82cc, 32'hc2895710, 32'h42d1a90b},
  {32'h44f7bdee, 32'hc2ec8cf4, 32'hc3e04197},
  {32'hc3329c00, 32'h43833fb6, 32'h424d2c49},
  {32'h44c9fd74, 32'h433baf6a, 32'h43188b6f},
  {32'hc4fa319e, 32'h420fb678, 32'h420199ff},
  {32'h4413a98a, 32'h42118ae1, 32'h4100e8e0},
  {32'hc487a5db, 32'h428e12c9, 32'hc0a31cfa},
  {32'h44c0697a, 32'h43722cbc, 32'hc2e0331e},
  {32'hc4342a13, 32'h4285b2e8, 32'hc2fc2deb},
  {32'h443abdce, 32'h43991566, 32'hc38e4417},
  {32'hc414a8e8, 32'h410fb339, 32'h434ecd86},
  {32'h4434a260, 32'h43342b31, 32'hc220dd66},
  {32'hc467a4af, 32'hc2ae626a, 32'h42347430},
  {32'h449a6c64, 32'h430b6e8f, 32'hc366101c},
  {32'hc4b17e23, 32'hc13a4be4, 32'hc2b39012},
  {32'h442a1a08, 32'hc43065fd, 32'h4337a580},
  {32'hc45b061e, 32'hc3577207, 32'hc27cafa3},
  {32'h44f72337, 32'h431130ad, 32'h41ec877f},
  {32'hc4ad2d81, 32'hc30047bc, 32'h441e7fac},
  {32'h44e63db3, 32'hc30334b5, 32'hc3ad2397},
  {32'hc4e0af4d, 32'hc35758bf, 32'h431b359f},
  {32'h44cf010d, 32'h425dd9fd, 32'h42504418},
  {32'hc41a2aab, 32'h436b933d, 32'hc195f4b0},
  {32'h431146be, 32'hc308eb9e, 32'hc313ddfb},
  {32'hc4ead357, 32'h43190275, 32'hc2fff923},
  {32'h44da2a4f, 32'h441f9ac2, 32'h432055ed},
  {32'hc4e7f62e, 32'hc2d0e2a2, 32'h430d6a9c},
  {32'h4444ffba, 32'hc2e36909, 32'hc2291026},
  {32'hc367e348, 32'hc25ed6dd, 32'h412cee8c},
  {32'h44865aa6, 32'h4386485a, 32'h42149e2a},
  {32'hc5288060, 32'hc2f20484, 32'hc3649188},
  {32'h44bf037a, 32'hc23755d8, 32'h439cbecd},
  {32'hc2d7c8c8, 32'hc35d4d58, 32'h432cdf7b},
  {32'h44f57f01, 32'hc28b3443, 32'hc344c109},
  {32'hc4dce40b, 32'h440839da, 32'hc30d4c02},
  {32'h44a18830, 32'h41a1ac87, 32'h4372eb07},
  {32'hc4732ae2, 32'hc33bb4a4, 32'hc32eb8d6},
  {32'h4292d020, 32'h43082dee, 32'hc292fc5b},
  {32'hc462cc2c, 32'hc23391be, 32'hc3885288},
  {32'h44424afe, 32'h43230899, 32'h43c41a0b},
  {32'hc4b7cb14, 32'hc2fe571c, 32'h42d4db86},
  {32'h44353dc6, 32'h437b8627, 32'hc2c068c9},
  {32'hc46b1044, 32'hc2d4fce9, 32'hc2fe7a15},
  {32'h4420f2ea, 32'h4330f6db, 32'h431fd207},
  {32'hc468b9d8, 32'hc32bbc61, 32'hc33ae9dc},
  {32'h438300be, 32'h43e6f332, 32'hc315c9f3},
  {32'h41b94280, 32'hc30f7a96, 32'hc272e2c3},
  {32'h44fc343e, 32'hc3a27126, 32'h43a07e5f},
  {32'hc39fc7c0, 32'h43966ced, 32'hc2acd94d},
  {32'h448105a9, 32'h4227a60d, 32'h42a750fa},
  {32'hc4e8943f, 32'h4291cdd2, 32'h436ec535},
  {32'h44eae5cf, 32'hc2d4bd66, 32'hc332e692},
  {32'hc4fadce8, 32'h430e7c27, 32'hc254a7d3},
  {32'h44969cc8, 32'hc2075148, 32'h4316e029},
  {32'hc43cb446, 32'h42245424, 32'hc3818a8b},
  {32'h4457f1c4, 32'h439cbd02, 32'h438f3016},
  {32'hc5101e2a, 32'hc240fb24, 32'h433cc92c},
  {32'h4516d5c4, 32'h44087e08, 32'hc30adb54},
  {32'hc4095556, 32'h43d652cf, 32'hc1fba997},
  {32'h43fbda18, 32'hc228d9d6, 32'hc29b15b2},
  {32'hc3b0382a, 32'h43a52451, 32'h42ace611},
  {32'h4523d289, 32'h4237f94c, 32'h4316ec36},
  {32'hc4a4207e, 32'h43bd98d8, 32'h4302dfd7},
  {32'h438d0110, 32'hc283caa3, 32'hc3d1a8a1},
  {32'hc503b3de, 32'h42199dcf, 32'hc280009a},
  {32'h4408bc70, 32'hc247468f, 32'h42fd876d},
  {32'hc39a8ff7, 32'h43121f0f, 32'h4310dc47},
  {32'h433d3654, 32'h43008cd3, 32'h42ce1051},
  {32'hc5001f88, 32'hc289c69d, 32'hc29412df},
  {32'h4440c9e0, 32'h416b9e54, 32'h43e633ea},
  {32'hc50e07eb, 32'h44163801, 32'hc3576900},
  {32'h44033bad, 32'hc239ccc8, 32'h422df9bd},
  {32'hc488d2b8, 32'h419639f7, 32'hc361db4c},
  {32'h43f5ed01, 32'hc310ffcd, 32'hc234df51},
  {32'hc4ea29c5, 32'hc1c6b5ed, 32'h4398b70a},
  {32'h4513fd63, 32'hc3659bce, 32'h422c0f31},
  {32'hc3d5f520, 32'h43a64ab1, 32'h430e6fdc},
  {32'h450e30ef, 32'h434856c8, 32'h438aa275},
  {32'hc4af8f6e, 32'h436159e1, 32'hc236d5cf},
  {32'h44c9f138, 32'h4230e84d, 32'hc3288712},
  {32'hc3ba7b0c, 32'h41573b67, 32'hc3d030b6},
  {32'h44c8273c, 32'h43944864, 32'hc2bdeb35},
  {32'hc495e04c, 32'hc3c77b1a, 32'hc3902faa},
  {32'h4399b050, 32'h4387f50f, 32'h4330747c},
  {32'hc480f67b, 32'h43c5f92c, 32'hc2fcfb4d},
  {32'h451bbab8, 32'hc3236dda, 32'hc389ce73},
  {32'hc2eec240, 32'hc2af9b1e, 32'h4285a7c8},
  {32'h43ae223a, 32'h421bb575, 32'h4382760d},
  {32'hc407b557, 32'hc2d5a585, 32'hc384a732},
  {32'h4500e03e, 32'h4211803c, 32'h42865649},
  {32'hc490e48f, 32'h43723f88, 32'hc370daa9},
  {32'h45059838, 32'h419b9934, 32'h42425af3},
  {32'hc2a96036, 32'h43b4fe0a, 32'hc12a0ead},
  {32'h44f346d2, 32'h42a8c0d7, 32'hc16f014a},
  {32'hc4583463, 32'hc2057b1e, 32'hc302529e},
  {32'h44b6dd52, 32'hc2f9b758, 32'hc38a2079},
  {32'hc4a468fe, 32'h4336acbe, 32'h433a6622},
  {32'h4412db76, 32'h43928306, 32'hc3834d12},
  {32'hc44b4614, 32'hc3568d1d, 32'h437567b7},
  {32'h44caba68, 32'hc27f9d5b, 32'h4402b010},
  {32'hc50700eb, 32'hc2eca411, 32'h41fd8919},
  {32'h4506da2e, 32'hc271e4d2, 32'hc368c18c},
  {32'hc50b948e, 32'h42af0914, 32'hc32809ea},
  {32'h43cc0080, 32'h42f29c40, 32'h43dd36c3},
  {32'hc43d9072, 32'hc29b92fe, 32'hc3c0a0f0},
  {32'h442dff67, 32'hc3412b79, 32'h4175c798},
  {32'hc49ea0a0, 32'hc3e67c1f, 32'hc3c1e7d4},
  {32'h44e8df87, 32'hc3395431, 32'h42c8e7a8},
  {32'hc4a899f8, 32'h428f0657, 32'h43ce5f0a},
  {32'h432477c0, 32'h433fb0ea, 32'h40bc6552},
  {32'hc507bb91, 32'h43ab5fae, 32'hc3c3659c},
  {32'h44a3b045, 32'hc4131aa3, 32'h4432c7c1},
  {32'hc4d8636a, 32'h43730787, 32'h4232b757},
  {32'h448d43b4, 32'h43857380, 32'h439dbfdb},
  {32'h435941e8, 32'hc0a8b3a5, 32'h438d61a3},
  {32'h44cc967b, 32'hc35ada41, 32'hc08c9bd8},
  {32'hc489cbd8, 32'hc3b75abf, 32'h4338bb14},
  {32'h45078852, 32'h4279ebbe, 32'hc33ff57d},
  {32'hc4437022, 32'hc2b8ac88, 32'h425f77ca},
  {32'h44b1879e, 32'hc3457dda, 32'hc19bd9e7},
  {32'hc35ba0cf, 32'hc251cc0b, 32'hc4008de6},
  {32'h44870b57, 32'hc3828894, 32'h42852e15},
  {32'hc4dc5072, 32'hc3642105, 32'h4294c08d},
  {32'h4331c298, 32'hc33a1a97, 32'h4309dafe},
  {32'hc4729bfb, 32'h426b5863, 32'h4306f02c},
  {32'h44fa32f4, 32'hc318dd6c, 32'hc3269fdb},
  {32'hc40e6a87, 32'h4383e90b, 32'hc2ae265e},
  {32'h44b52272, 32'hc2cd2702, 32'hc33c4d13},
  {32'hc5130e6a, 32'hc3416354, 32'hc2e7491c},
  {32'h45165dea, 32'hc397cc20, 32'hc326713a},
  {32'hc321f08e, 32'hc30e864d, 32'h43473070},
  {32'h45118759, 32'hc385a040, 32'hc22bb6c8},
  {32'hc29a2ec0, 32'hc39b558a, 32'h419f3d30},
  {32'h44894c7f, 32'h41c3216c, 32'hc30abb26},
  {32'hc4b451d0, 32'hc401dbb9, 32'hc40be874},
  {32'h44b9ff96, 32'h4446a7e2, 32'h42e118c7},
  {32'hc3df9aa2, 32'hc3862b67, 32'h43a24bbe},
  {32'h43a4da18, 32'h418ea4b7, 32'hc3e64e07},
  {32'hc508262f, 32'h432dd615, 32'h439aac27},
  {32'h44cc3671, 32'hc328027e, 32'hc3880215},
  {32'hc512256c, 32'h435a321c, 32'hc2b9515a},
  {32'h4511ae8a, 32'h419a63ef, 32'hc2a35c4d},
  {32'hc44a75a0, 32'h43a855ef, 32'h4000e602},
  {32'h45066993, 32'h41f029bf, 32'hc3b5fbc1},
  {32'hc504c164, 32'h4326b55d, 32'h426ee926},
  {32'h44b3a8ef, 32'hc31f01a5, 32'hc21ff787},
  {32'hc1c86d80, 32'hc390c5d6, 32'h415aea82},
  {32'hc2ded830, 32'h4411f667, 32'h421aad6e},
  {32'hc4e81ec6, 32'hc3162133, 32'h4331696e},
  {32'h446339f9, 32'h4256331d, 32'hc2223e38},
  {32'hc4cef113, 32'h41146443, 32'hc1188bfe},
  {32'h44ef53f6, 32'hc313f7d9, 32'hc13e8d30},
  {32'hc507d9ca, 32'hc3233e37, 32'hc12bdb3d},
  {32'h441d542e, 32'h42fdf385, 32'h43928ffc},
  {32'hc4a86f0a, 32'hc1051334, 32'h432dfa98},
  {32'h443ce0da, 32'h42b91bb2, 32'hc33294ba},
  {32'hc35a62fc, 32'hc3d309e7, 32'hc30d0f5d},
  {32'h441cc6ae, 32'h42d8d785, 32'hc323d1a5},
  {32'hc4088410, 32'h4200e629, 32'h42ec25c4},
  {32'h451bb674, 32'h4146899b, 32'hc23d5683},
  {32'hc1a89100, 32'hc3b1a239, 32'h43f64246},
  {32'h44c7777a, 32'h42c89549, 32'hc2134b41},
  {32'hc4d849c7, 32'h43dcef84, 32'h42479eaf},
  {32'h449de9a7, 32'hc2f6dacc, 32'h4111f354},
  {32'h43507e89, 32'hc2a9948e, 32'hc3b1f072},
  {32'h44e63bbb, 32'h42b4a204, 32'hc34da69a},
  {32'hc3bd10b0, 32'hc2c3a25d, 32'h43f5d2ba},
  {32'h44f05e02, 32'hc377bf95, 32'hc2ee309c},
  {32'hc5057016, 32'h42ea3435, 32'h41ec113f},
  {32'h44bff45e, 32'h4403102d, 32'h4347aac4},
  {32'hc4c1e91b, 32'h42e41027, 32'h432f8c30},
  {32'h448e013a, 32'hc254d4cb, 32'h4381273f},
  {32'hc4fc0224, 32'hc4054b0b, 32'hc2364f7b},
  {32'h44adb192, 32'hc35490c9, 32'hc203d294},
  {32'hc32edc80, 32'h430f6b69, 32'h435c5e8a},
  {32'h448ff828, 32'hc389d805, 32'hc31e77a0},
  {32'hc489b0d8, 32'h42f3923c, 32'hc262c0e9},
  {32'h44f39cd7, 32'h42b505c7, 32'hc2fe8084},
  {32'hc4594390, 32'hc208a8c3, 32'h43ec89f6},
  {32'h4502a3b5, 32'hc2d580b0, 32'hc42e514b},
  {32'hc4994124, 32'h43d92330, 32'hc28bbf37},
  {32'h44e64fc7, 32'h4145320f, 32'hc18de3cc},
  {32'hc3d4fca0, 32'h4298c49c, 32'h412a410e},
  {32'h4465d7b8, 32'hc2a3a8fe, 32'hc3422e23},
  {32'hc4d9c650, 32'hc38c1173, 32'h434c820a},
  {32'h44f734b2, 32'hc30910a4, 32'h42a3f0a0},
  {32'hc44d56f7, 32'h42fa6c47, 32'hc27c45ad},
  {32'h446e8435, 32'hc0be0c43, 32'hc36b24b9},
  {32'hc498f46e, 32'hc2be2d77, 32'h4320f05a},
  {32'h438e399c, 32'h432940fa, 32'hc3a2ca3c},
  {32'hc47667eb, 32'hc3452191, 32'h4397d105},
  {32'h4496241a, 32'h4311ad25, 32'hc3a8af1e},
  {32'hc4919212, 32'hc33e6a24, 32'hc3121d04},
  {32'h43c461bc, 32'h42278a70, 32'hc21fc4f0},
  {32'hc4002e69, 32'hc3ac7b35, 32'h43542019},
  {32'h449a833c, 32'hc22526df, 32'hc3fa9607},
  {32'hc4e63024, 32'h43bb3702, 32'h43bbd1de},
  {32'h44ba7a3c, 32'h42b034cd, 32'hc383d192},
  {32'hc4bbe604, 32'h42dc3044, 32'h43b69ded},
  {32'h44c57aeb, 32'h4393b96a, 32'h42d4e595},
  {32'hc4152bf8, 32'hc18aa662, 32'h431ec14b},
  {32'h44ed0b2e, 32'h440087e6, 32'hc3a6361a},
  {32'hc50891df, 32'hc2800859, 32'hc306e72d},
  {32'h44159ef5, 32'hc25f7ffc, 32'hc3149086},
  {32'hc4de0f06, 32'hc2e1aecc, 32'h421abfa4},
  {32'h451a327c, 32'hc2e5fe16, 32'hc3c6f52a},
  {32'hc4c12e10, 32'h41dc838d, 32'h42628dff},
  {32'h448d1bf8, 32'hbf473fd4, 32'hc2489a73},
  {32'hc493d73f, 32'hc314e23a, 32'hc3332eb5},
  {32'h433cb9b0, 32'h43a6ca8e, 32'hc297d772},
  {32'h4296019e, 32'h429d69fa, 32'h43c3f0dd},
  {32'h450c3256, 32'hc0872039, 32'h427dc2b8},
  {32'hc4b065ba, 32'hc25d7b14, 32'h440e716f},
  {32'h449f8218, 32'h406e240d, 32'hc3a4df42},
  {32'hc2b42050, 32'h42b38486, 32'h435445b2},
  {32'h45034ecc, 32'hbf881bb2, 32'h43929823},
  {32'hc4a869a7, 32'hc391fda4, 32'hc20f3ef0},
  {32'h43958193, 32'hc13cee96, 32'h3f9d38de},
  {32'hc5002c68, 32'h42c573dc, 32'h42c44ef9},
  {32'h445b976a, 32'hc40c34a5, 32'hc3cbc65b},
  {32'hc370e440, 32'hc39884dc, 32'hc32a3881},
  {32'h429348c0, 32'hc29e69dc, 32'hc37830cb},
  {32'h44b390a2, 32'h42b62aaa, 32'h42382342},
  {32'hc4444c66, 32'h43778c5f, 32'h42791c75},
  {32'h43460638, 32'hc2f42c23, 32'h42022862},
  {32'hc4a7f1af, 32'hc2a3f59c, 32'hc36fb458},
  {32'h44cec742, 32'hc2966a30, 32'hc336e069},
  {32'hc4fab8b3, 32'h40d22996, 32'hc2be5425},
  {32'h44d059e3, 32'h431f76e1, 32'hc2c24ac7},
  {32'hc389e36c, 32'hc2abc5cc, 32'h42fed60e},
  {32'h4449b968, 32'hc395f42a, 32'h4281e1bf},
  {32'hc4ea3752, 32'hc295e3c8, 32'hc3d60d28},
  {32'h44f28ef6, 32'hc2ec3176, 32'h43a9ae1f},
  {32'hc323dc1a, 32'hc1f93e6f, 32'hc41c2449},
  {32'h448b45ff, 32'hc2b4ab72, 32'hc34647a7},
  {32'hc3c689e4, 32'hc3f46180, 32'h42d20ce1},
  {32'h43f61dfa, 32'h428d2b15, 32'hc293f6ef},
  {32'hc506931b, 32'h43f2af54, 32'hc38bb22f},
  {32'h44a3b6c2, 32'h439f42f3, 32'h43b55308},
  {32'hc1bec700, 32'hc40c11d7, 32'h421903cf},
  {32'h450706b8, 32'h4381fde0, 32'h42a99fb3},
  {32'hc3db8f22, 32'h4407ee1a, 32'hc19405f2},
  {32'h44ae97f5, 32'hc399bf10, 32'hc390c3f6},
  {32'hc3b6a500, 32'h4291099e, 32'h42e50210},
  {32'h44f32f30, 32'h42da862f, 32'hc30bf285},
  {32'hc4d58de4, 32'h4209f2f2, 32'h424a76ae},
  {32'h44d315e8, 32'hc31f83ab, 32'hc377e02d},
  {32'hc4bfc12d, 32'h42b87837, 32'h43b51a10},
  {32'h44f89733, 32'hc288fe4d, 32'hc2a955ef},
  {32'hc4efd7c0, 32'h42246797, 32'hc2a7f4d7},
  {32'h440a6640, 32'h4303151a, 32'hc38d1f1a},
  {32'hc3f72078, 32'h4286684b, 32'hc3da73ab},
  {32'h44d49519, 32'hc364a217, 32'h431102f0},
  {32'hc3e3a472, 32'hc31ee026, 32'h42d9837c},
  {32'h452053e9, 32'h4334e13b, 32'hc2ac8417},
  {32'hbfbb0500, 32'hc2a06fdd, 32'h423c3103},
  {32'h44975625, 32'hc396101f, 32'hc38785e1},
  {32'hc4ac387e, 32'hc3b97152, 32'h4398655e},
  {32'h44bb0901, 32'hc365902a, 32'h432e5335},
  {32'h439e3f50, 32'hc330e8b8, 32'hc3f34232},
  {32'h44cc6c9e, 32'hc378529d, 32'h41e8f8f2},
  {32'hc2e8e078, 32'hc3ad254d, 32'hc30732a2},
  {32'h44f6d8ab, 32'h430b9c4a, 32'h42c5daa3},
  {32'hc491a224, 32'h428d1392, 32'hc37e3281},
  {32'h450672f7, 32'hc3bab08b, 32'h43f3ed62},
  {32'hc4824d40, 32'h43c4006b, 32'h432e9592},
  {32'h4440f01c, 32'h4371ea76, 32'hc23d86a2},
  {32'hc50dc415, 32'hc3eee042, 32'hc3ac48b6},
  {32'h44fdbd56, 32'h42829176, 32'h4339d595},
  {32'hc4e51d0b, 32'h43599afe, 32'h43c28f39},
  {32'h4514fcd2, 32'h42839f90, 32'h41b17b94},
  {32'hc5097c1a, 32'h436276aa, 32'hc316a470},
  {32'h43c22f2c, 32'h43523ec2, 32'hc360fdb5},
  {32'hc42365d4, 32'h43418348, 32'h43aa988d},
  {32'h43d4381a, 32'h4287c489, 32'h4390f3a7},
  {32'hc4b11b74, 32'h4357befd, 32'h41b906b7},
  {32'h450f9e0e, 32'hc3a36e02, 32'hc343b250},
  {32'hc4dda42a, 32'hc20b72ce, 32'h4135cf0b},
  {32'h440ce1b4, 32'hc340967a, 32'hc3e57f76},
  {32'hc51092c1, 32'h44020d14, 32'hc40c7183},
  {32'h45157baf, 32'hc2983a85, 32'hc2bc525c},
  {32'hc4ecf4c1, 32'h430bd3f6, 32'hc270c739},
  {32'h44659872, 32'hc34b964b, 32'h43108388},
  {32'hc50fb12d, 32'h42863d80, 32'hc3829ded},
  {32'h449183c9, 32'hc3bfedaa, 32'h425ee0c5},
  {32'hc41f9a50, 32'h4297fe7f, 32'hc2a33fd0},
  {32'h44bd8994, 32'h43784ee5, 32'hc1e81a76},
  {32'hc50c9c50, 32'h43b895b8, 32'h4315319f},
  {32'h43c36950, 32'h42cd93ab, 32'hc3aca465},
  {32'hc48867b4, 32'h4302d9e1, 32'h42910e9e},
  {32'h44c7538b, 32'h42e76942, 32'h44154ba6},
  {32'hc40611da, 32'hc38840f7, 32'h43c1aaf2},
  {32'h4500d9eb, 32'hc387d51d, 32'h43254b86},
  {32'hc4f75bd2, 32'hc30a09ae, 32'h420843b1},
  {32'h442e9ed8, 32'h42d2ceaf, 32'hc2a8b7af},
  {32'hc496a3e2, 32'hc2a64750, 32'h426e2026},
  {32'h44b78973, 32'hc2ebc35b, 32'hc31ae4e8},
  {32'hc40555ec, 32'hc1bd74b2, 32'h4335d5e7},
  {32'h44f5cbe9, 32'h428519b8, 32'hc36b049e},
  {32'hc460fa03, 32'hc2019bbf, 32'h424efe4e},
  {32'h44a0f297, 32'h41bc170b, 32'h416d3868},
  {32'hc495b060, 32'h3ea51c7c, 32'hc3423e45},
  {32'h449ae518, 32'h42b1987d, 32'hc2bdc7ab},
  {32'hc4a1b580, 32'hc3d2069f, 32'h41cbe950},
  {32'h44f4e157, 32'hc2bf14b1, 32'hc3e3ed01},
  {32'hc4f44ff8, 32'hc34bda8e, 32'hc3a7f402},
  {32'h44ac3085, 32'hc355c051, 32'hc2dcc8eb},
  {32'hc4fe60f1, 32'h439b40a6, 32'hbf548b20},
  {32'h44f0ea66, 32'hc29d7e71, 32'hc2beb579},
  {32'hc12e6c6a, 32'hc2ba7ce0, 32'hc28fc7c8},
  {32'h448800b0, 32'h431f9061, 32'h41c4a6ff},
  {32'hc4fd672b, 32'h4317ba25, 32'hc393dd5a},
  {32'h45037269, 32'hc29ad0a4, 32'h41888104},
  {32'hc36377ac, 32'h42a1aa52, 32'hc2067a55},
  {32'h44ee6703, 32'h43c3f069, 32'hc3aa11fd},
  {32'hc29e6ab0, 32'hc3455137, 32'hc3f7c039},
  {32'h44ab54c5, 32'h44082d05, 32'h434e3ee6},
  {32'hc35df7bc, 32'hc228eb40, 32'hc3622576},
  {32'h44365f05, 32'hc40de28d, 32'h4400c7e4},
  {32'hc438a61b, 32'hc292d068, 32'hc39fa23c},
  {32'h441178ed, 32'hc42cc80f, 32'hc289e683},
  {32'hc460f718, 32'h43855320, 32'h418bee7f},
  {32'h44830d30, 32'hc2de9963, 32'h429927e9},
  {32'hc3c4ecc0, 32'h428026d1, 32'hc331ef45},
  {32'h44ce95c6, 32'h42b1a71e, 32'h43a0ed1c},
  {32'hc340fe58, 32'hc22460e6, 32'h40baa390},
  {32'h447f62bb, 32'hc2fd1c94, 32'hc2dda250},
  {32'hc5146a32, 32'hc29f989d, 32'hc2556666},
  {32'h44bde651, 32'hc28a9671, 32'hc3b416a1},
  {32'hc4d209cc, 32'hc241a4dc, 32'hc343962c},
  {32'h444fe8a4, 32'hc3200517, 32'h4341cf24},
  {32'hc4fcd18b, 32'h4350b6c3, 32'h414117fa},
  {32'h44e96540, 32'h434671bf, 32'hc38179dd},
  {32'hc4e67c49, 32'hc31a59a8, 32'hc35dc90c},
  {32'h442f2529, 32'hc3baf964, 32'h43bab5d3},
  {32'hc4f80111, 32'h417d9cd5, 32'h439d9993},
  {32'h451fb482, 32'h434d227b, 32'hc2260a30},
  {32'hc3f6eea4, 32'hc322b896, 32'hc3a57d11},
  {32'h44d00ab7, 32'hc2e89dff, 32'h42a51c11},
  {32'hc32dcbd8, 32'hc3734a8f, 32'h43b27e0e},
  {32'h44fbc0bc, 32'hc27bdd31, 32'hc0c929df},
  {32'hc4a70830, 32'hc3047322, 32'hc3b68fb0},
  {32'h435fa7e0, 32'hc36c47e8, 32'h4385a9dc},
  {32'hc365b2ae, 32'hc38376b5, 32'h429ed3d9},
  {32'h44a0810c, 32'hc3355f74, 32'h43dc03a0},
  {32'hc4d13748, 32'hc2e96129, 32'h42c21990},
  {32'h4501687c, 32'hc1e77ce6, 32'h4381990a},
  {32'hc4da6d54, 32'h435b80de, 32'h42b4275b},
  {32'h43c81b84, 32'hc33c416f, 32'hc3fea256},
  {32'hc4e50f0e, 32'hc391b40c, 32'hbfc9dec2},
  {32'h44af22b0, 32'h43ca3f32, 32'hc27cc15b},
  {32'hc4ecd700, 32'hc37f6738, 32'h43acfb74},
  {32'h451dbdae, 32'h4322ffc4, 32'h42c501d6},
  {32'hc4cbc4e0, 32'hc37bd935, 32'hc3156f21},
  {32'h42d224c0, 32'h428d7886, 32'h43060b5d},
  {32'hc3c90586, 32'h43401f41, 32'h4344e246},
  {32'h447d3a29, 32'h432edcf7, 32'hc3ca5826},
  {32'hc4a4c08b, 32'h4167e4ca, 32'hc2b391a1},
  {32'h44e85995, 32'h429f4073, 32'h41e24f71},
  {32'hc5170a1c, 32'hc30c4536, 32'h428a5a0c},
  {32'h444be004, 32'hc3c886cf, 32'hc3333e97},
  {32'hc3b87b06, 32'hc31f3f07, 32'hc289d033},
  {32'h447d0339, 32'h4299baf8, 32'hc34a67b3},
  {32'hc512cd4e, 32'hc34692ca, 32'h4312a450},
  {32'h44651a5b, 32'hc30890d4, 32'hc3225386},
  {32'hc2c0b260, 32'h41509a44, 32'h407a6f58},
  {32'h451bc0b1, 32'h428c48ee, 32'h42d2ab7d},
  {32'hc3d3ae20, 32'hc3bb41f8, 32'h43a6ea33},
  {32'hc36afcb8, 32'hc3898a30, 32'h436722dc},
  {32'hc49240b9, 32'h433ccec4, 32'h43966e82},
  {32'h42f6d090, 32'hc3258c2f, 32'h43b57361},
  {32'hc4aef5f9, 32'hc36a6089, 32'hc352a94a},
  {32'h44ae646e, 32'h439c7f10, 32'hc29fd0f1},
  {32'hc4abeca9, 32'hc17b2c2c, 32'h42191a72},
  {32'h43d8007b, 32'h43928af2, 32'hbf897e53},
  {32'h42c11b79, 32'hc277f733, 32'h4268d78f},
  {32'h438de608, 32'hc354c75b, 32'h4255a1e1},
  {32'hc38519b0, 32'hc21e35a3, 32'h411e72fa},
  {32'h449152e8, 32'h43b536b6, 32'hc30cfed2},
  {32'hc42860a6, 32'h4353b51d, 32'h43a1720a},
  {32'h44ff0d54, 32'h434d4f57, 32'hc40224cd},
  {32'hc4a7db78, 32'h41853df2, 32'hbebecb88},
  {32'h44cfff23, 32'h42ec9c2d, 32'h4390811b},
  {32'hc349b834, 32'hc3d153c4, 32'hc2003c14},
  {32'h44b211eb, 32'h43cb9e46, 32'hc36691eb},
  {32'hc4dd13bc, 32'hc2169ffb, 32'h440746a5},
  {32'h438a86ec, 32'h430b00dd, 32'h4373c821},
  {32'hc3c808c4, 32'h42e0b42a, 32'hc3413125},
  {32'h44a663eb, 32'hc2cfbd9e, 32'hc1a9edd8},
  {32'hc4e43191, 32'hc33ef1c6, 32'hc3adbf20},
  {32'h4509fee8, 32'hc2ae1719, 32'hc2f9bb28},
  {32'hc2b93c40, 32'hc3866ce8, 32'h4294568d},
  {32'h450b36bd, 32'hc2525758, 32'hc348e274},
  {32'hc508cd53, 32'hc3e69a6d, 32'h42ef16fe},
  {32'h44486f66, 32'h438d33a2, 32'h431477cc},
  {32'hc4cf2577, 32'h4316748f, 32'hc3639cd4},
  {32'h44ee8e1a, 32'h434c2145, 32'hc21f0612},
  {32'hc4f5ddf6, 32'h43e2bd23, 32'h42b1caf7},
  {32'h437f8989, 32'h41de0745, 32'h4399257d},
  {32'hc4d42b86, 32'hc3c1192e, 32'hc31384fc},
  {32'h436e3c60, 32'hc34bba72, 32'h437d77e4},
  {32'hc4fd18d9, 32'hc38dd7ad, 32'h439119f8},
  {32'h43f67d17, 32'h41e18fb5, 32'h43b425fc},
  {32'hc4f7d157, 32'hc38c9aa0, 32'hc3c0f3a5},
  {32'h4472aa36, 32'h4128c19a, 32'hc36b1fa2},
  {32'hc410be82, 32'hc3903a27, 32'hc362c17d},
  {32'h442046dc, 32'h43082859, 32'hc320b9c3},
  {32'hc49dca63, 32'hc096db9a, 32'hc254fc6c},
  {32'h44d78e35, 32'h43338efc, 32'hc3391970},
  {32'hc37d24fe, 32'h42539ed4, 32'hc2c29b32},
  {32'h448ab9c4, 32'hc39d3295, 32'hc22611a4},
  {32'hc3f299df, 32'hc1453a13, 32'h43310e88},
  {32'h44957bdc, 32'h425734f0, 32'h4371adde},
  {32'hc4b31a98, 32'h437ff4ed, 32'h43bbe23e},
  {32'h44451bf3, 32'h43012ca2, 32'h43078be3},
  {32'hc504fd94, 32'hc3603972, 32'hc219187b},
  {32'h450a9bdb, 32'h43daa942, 32'h432faab2},
  {32'hc487ab40, 32'h420d6d6d, 32'h43212d23},
  {32'h44bc4692, 32'h4393f2c6, 32'hc3847b3e},
  {32'hc4fecd51, 32'hc308a1c7, 32'h43591f7f},
  {32'h441b44a4, 32'h4298dea5, 32'h43ae3e6c},
  {32'hc4466d02, 32'h43413fcd, 32'h41aaef86},
  {32'h4403c818, 32'hc41d2675, 32'h43149141},
  {32'hc38b9cd0, 32'hc3209be4, 32'hc2ff8e94},
  {32'h44ff6a24, 32'hc3926591, 32'hc3afdf7a},
  {32'hc4cd7a5e, 32'hc29a8934, 32'h4168c001},
  {32'h44bbf15b, 32'hc42e2bf9, 32'h43b49aa4},
  {32'hc50f1441, 32'h43c506d2, 32'hc2e1b5e4},
  {32'h4508bf33, 32'hc344d47a, 32'hc3bc3464},
  {32'hc47e2796, 32'h44152f18, 32'hc365b976},
  {32'h440baae4, 32'h43a9565d, 32'hc301f53f},
  {32'hc50bd143, 32'h42f062cf, 32'h4369b43c},
  {32'h446d8e58, 32'h42adbe6c, 32'hc1bc8524},
  {32'hc40f6f74, 32'hc36eb11a, 32'h4271d27e},
  {32'h44c295ad, 32'h43df0bc7, 32'h43aff273},
  {32'h42bd4f20, 32'h4336aac5, 32'h43c22c41},
  {32'h44568838, 32'h430176d5, 32'h43bcb1a9},
  {32'hc4f5bf5a, 32'hc2e83194, 32'hc2e865b5},
  {32'h44d82ac3, 32'hc3876bec, 32'hc3cb1e7f},
  {32'h430daa7c, 32'hc3468481, 32'h43c1fd05},
  {32'h44a2f1de, 32'h420eee6d, 32'hc35e80fe},
  {32'h43357acc, 32'h43d98737, 32'hc2042017},
  {32'h44a986b7, 32'hc32f322b, 32'h424d46f4},
  {32'hc4e49dcf, 32'h42da5b8a, 32'h4382710a},
  {32'h44fa116e, 32'h4387a2d1, 32'h429e34c4},
  {32'hc50cde4a, 32'hc35296e5, 32'hc23b1a11},
  {32'h450f6167, 32'hc43be5f1, 32'hc2bc0fdd},
  {32'hc4b1b706, 32'h4211b4f4, 32'h42ba07e2},
  {32'h4394d221, 32'h42332a55, 32'hc2413aee},
  {32'hc4cbf5a8, 32'hc180950c, 32'hc30f672d},
  {32'h450031e2, 32'h43840e90, 32'h4395e3ce},
  {32'hc487bf5f, 32'hc1f7b762, 32'hc2a13f04},
  {32'h44961c4f, 32'h434f3016, 32'h42a6ff45},
  {32'hc3de9a44, 32'h42d925fc, 32'hc3320af5},
  {32'h450b19d6, 32'hc32b09f3, 32'h4399a4bd},
  {32'hc4144ef0, 32'hc3186d0b, 32'hc3491da0},
  {32'h4515be59, 32'hc28531eb, 32'h436f319f},
  {32'hc4e0e779, 32'h42a26e10, 32'h42401345},
  {32'h44d54627, 32'hc317a39b, 32'hc2aa8195},
  {32'hc4e0a285, 32'hc4004800, 32'hc3ef3262},
  {32'h445351b2, 32'hc305615b, 32'h4327166e},
  {32'hc515c7b8, 32'hc21568f9, 32'h435936a5},
  {32'h4407deb6, 32'h436f884e, 32'hc3d8b25c},
  {32'hc3446810, 32'hc1f53290, 32'hc1332784},
  {32'h441ed954, 32'hc3904162, 32'h438458c0},
  {32'hc4ee1bd6, 32'h42ed9f0d, 32'hc23c4659},
  {32'h45070c82, 32'hc353bd10, 32'hc4117da1},
  {32'hc4870f0e, 32'h42cd6758, 32'hc350f0d8},
  {32'h442710e8, 32'hc35aec18, 32'h4377a9cc},
  {32'hc47938f7, 32'h4381f331, 32'hc320f39a},
  {32'h44a9ac1a, 32'h43b4d2ea, 32'hc30cf405},
  {32'hc4da567a, 32'h41272efd, 32'hc344cdf4},
  {32'h442de612, 32'hc2668660, 32'hc35e874f},
  {32'hc4d1fcd9, 32'h43951935, 32'hc2a762fe},
  {32'h444b0971, 32'hc3450561, 32'h4335024f},
  {32'hc4f298b2, 32'hc3cc82f2, 32'h4358b66e},
  {32'h44ce655e, 32'h43621c93, 32'hc38b2970},
  {32'hc365d01d, 32'hc3211034, 32'hc410da55},
  {32'h450d273d, 32'h435c40e8, 32'h43ab705b},
  {32'hc3e54d72, 32'hc239c552, 32'hc341f322},
  {32'h449932e2, 32'hc1a5565a, 32'h435d8af5},
  {32'hc4a1d0dd, 32'hc38e3983, 32'hc3e16074},
  {32'h45167c7d, 32'hc0c8c596, 32'hc184b29c},
  {32'h430029b0, 32'h439e0b02, 32'hc205d9ef},
  {32'h444d5435, 32'hc3a06f75, 32'hc33c644b},
  {32'hc45968d0, 32'hc38f2db1, 32'hc292fafd},
  {32'h451626d4, 32'h4118af16, 32'h42e8f6e3},
  {32'h432b1220, 32'hc1d08137, 32'h43b8bc44},
  {32'h44ed4252, 32'h4381690c, 32'hc2919ca8},
  {32'hc4a71bb7, 32'h4340f607, 32'h43a14d8e},
  {32'h44236de8, 32'hc315f724, 32'hc29c2bb4},
  {32'hc41fec40, 32'hc2adff90, 32'hc259f834},
  {32'h448ed0cc, 32'h43835ee9, 32'hc278716c},
  {32'hc508f822, 32'h438d0604, 32'h43db549a},
  {32'h431fa160, 32'h4222c1b4, 32'h418a589e},
  {32'hc4012188, 32'h42814daa, 32'hc2de2ff8},
  {32'h44e90c28, 32'hc2d81c98, 32'hc2b7a019},
  {32'hc4b2597e, 32'hc393d032, 32'h4343f7bd},
  {32'h44e2c68b, 32'h42ee584d, 32'hc21968e0},
  {32'hc46da3a3, 32'hc3a2ecc9, 32'h438db774},
  {32'h434de9f3, 32'h43ebcd5b, 32'hc32bb7d3},
  {32'hc50be72e, 32'h43db7b43, 32'hc23bf306},
  {32'h44cfa095, 32'h43a8fe2e, 32'hc3054256},
  {32'hc505932f, 32'hc39073bc, 32'h43590f72},
  {32'h44376348, 32'h42fe3c72, 32'h42eb88df},
  {32'hc35158c8, 32'h4347b6ad, 32'hc2cfe921},
  {32'h43eeac9e, 32'h4288de5c, 32'h42440471},
  {32'hc4f9e808, 32'hc333d38a, 32'hc3122371},
  {32'h44d9f755, 32'h429daf02, 32'h4313b7cf},
  {32'hc3889978, 32'hc2ba625a, 32'hc315d4ad},
  {32'h4441a356, 32'hc33f6dab, 32'hc38c2356},
  {32'hc50b15bb, 32'hc34b4727, 32'h43bee310},
  {32'h44cb3477, 32'hc3329b83, 32'h4341b4f4},
  {32'hc45944c8, 32'h4390b075, 32'hc3e7b723},
  {32'h44fb33f7, 32'hc0b92fe3, 32'hc295c705},
  {32'hc4597a72, 32'h435e640d, 32'h42b71d44},
  {32'hc24d4a80, 32'hc3fce8c9, 32'hc2d3e618},
  {32'hc4690d81, 32'hbf26792e, 32'hc2efb3ae},
  {32'h44dd2497, 32'h41792452, 32'h43f2f990},
  {32'hc51b8d8c, 32'hc25a4279, 32'h4367df99},
  {32'h42d39750, 32'hc30d15fd, 32'hc2f5764e},
  {32'hc332e480, 32'h43ecf116, 32'hc353c80a},
  {32'h4521b31c, 32'h43c088e8, 32'hc3c98262},
  {32'hc300f075, 32'hc20550f9, 32'h434c77d3},
  {32'h4516289f, 32'hc386d68d, 32'hc38678e2},
  {32'hc2ce3810, 32'h43282b6d, 32'hc2d1a0e1},
  {32'h451459c6, 32'hc2dc35ba, 32'hc3e0e576},
  {32'hc48f395e, 32'h424dccdb, 32'hc2f72e76},
  {32'h44bcd0e8, 32'hc3c094e8, 32'hc26713bd},
  {32'hc4bea1a3, 32'h42f5925a, 32'hc26dfc89},
  {32'h44fe53e8, 32'hc2cb09af, 32'hc3a70d99},
  {32'hc4da9043, 32'h433e1803, 32'h42d14886},
  {32'h43f264a0, 32'h434d7f77, 32'hc2473d51},
  {32'hc4ccf934, 32'h4384ed9d, 32'hc2bf323c},
  {32'h451610d2, 32'h42445e63, 32'h433e417e},
  {32'hc48105f0, 32'h4397a9c1, 32'hc321472d},
  {32'h450c07de, 32'h4375aec8, 32'hc316b466},
  {32'hc4af3372, 32'hc14c79f1, 32'h4415e768},
  {32'h447e7a0e, 32'hc399f34a, 32'hc33f85d7},
  {32'hc5049de5, 32'hc39f92be, 32'h432cb9a4},
  {32'h44fd6234, 32'hc29c56d2, 32'hc209eb11},
  {32'hc45a34be, 32'h42c2ae6d, 32'h434d9109},
  {32'h44e96f32, 32'hc2931ce1, 32'hc3ee02f5},
  {32'hc4620bc6, 32'h43bf6e5b, 32'h431fdd1d},
  {32'h4498bf4c, 32'h426e0d9b, 32'hc19c89de},
  {32'hc4c34c56, 32'hc323fe7f, 32'hc35c4ef8},
  {32'h44e6c319, 32'h41b7e8e2, 32'h41c22f52},
  {32'hc4cce1bd, 32'hc196233f, 32'hc1ba290e},
  {32'h4441bdac, 32'hc28e5f44, 32'hc24e4200},
  {32'hc4f119a1, 32'hc291b7bf, 32'hc37d3dc0},
  {32'h44edd244, 32'hc3c81da4, 32'hc3b6fc50},
  {32'h43a1fa64, 32'h436bf2de, 32'hc2533c7f},
  {32'h44f27b9a, 32'hc2f755fb, 32'hc3307ef5},
  {32'hc4c66336, 32'hc15e2158, 32'hc2e860f0},
  {32'h44ca974c, 32'h4076a2d0, 32'hc349abd7},
  {32'hc3a412c5, 32'h4380869b, 32'h42fe6210},
  {32'h4359e109, 32'hc2e92e70, 32'hc360f3f0},
  {32'hc443caf4, 32'hc2f0e09e, 32'h425e73ed},
  {32'h43b7c612, 32'h431e5799, 32'h43c9ce36},
  {32'hc4dd740b, 32'hc4180cd1, 32'hc25d9f83},
  {32'h4501406d, 32'hc141a9d3, 32'hc30e3c15},
  {32'hc3bb4008, 32'hc177efec, 32'hc41d426e},
  {32'h44944437, 32'hc31dfde7, 32'h402278f8},
  {32'hc477af2d, 32'hc3501e21, 32'hc1b1a9c7},
  {32'h4424ea05, 32'hc1901a9c, 32'h43b8fd5c},
  {32'hc4bfe325, 32'h44005d9b, 32'hc2d17db9},
  {32'h44fa407c, 32'h435a55c8, 32'hc2e949ef},
  {32'hc449879d, 32'h435d58b5, 32'h436dc1e9},
  {32'h44ff3a7e, 32'hc38c97c5, 32'hc274b39e},
  {32'hc47b964c, 32'h430e668d, 32'h42a554ee},
  {32'h443c6cb1, 32'h42b5efc1, 32'hc22840b4},
  {32'hc4be9654, 32'hc3c0ce33, 32'hc2923989},
  {32'h44acf9e8, 32'hc32681c5, 32'h4334beda},
  {32'hc4afaa58, 32'hc24a553e, 32'h435f2495},
  {32'h436776ff, 32'hc2ae5630, 32'hc326921d},
  {32'hc50eed15, 32'h4198f9d6, 32'h414346be},
  {32'h43a1d97a, 32'hc10862c6, 32'hc2d8bc43},
  {32'hc500e965, 32'h43a4c37c, 32'h43c54111},
  {32'h450df33c, 32'h436788a2, 32'hc262d4c9},
  {32'hc5118304, 32'hc1c5f988, 32'h420bdc24},
  {32'h441e891d, 32'h43f25b72, 32'h42b65b52},
  {32'hc4db384a, 32'hc36ae0fa, 32'hc387ea60},
  {32'h43ba505c, 32'h41bb0102, 32'h438957b7},
  {32'hc4e74c67, 32'hc3040d1d, 32'hc3743115},
  {32'h40c97a00, 32'hc3523783, 32'hc37c9af5},
  {32'hc485db70, 32'h4058db68, 32'hc3377fee},
  {32'h43b706f6, 32'h42cedbf8, 32'hc38c7c8b},
  {32'hc4a66f4c, 32'h438e55a9, 32'hc2d8fefc},
  {32'h45249252, 32'hc36bf2a5, 32'hc2009555},
  {32'hc41fa437, 32'h438c220c, 32'hc34874f1},
  {32'h44decf2b, 32'hc38eca9f, 32'hbfa30b73},
  {32'hc49fbc2d, 32'h421851a6, 32'h43780d22},
  {32'h44dc1740, 32'h42a6fda7, 32'hc28d7642},
  {32'hc4b449e4, 32'hc315f631, 32'hc34648be},
  {32'h451ea44d, 32'hc338c3c2, 32'hc3a5a827},
  {32'hc48741db, 32'h438cb529, 32'hc1fefee6},
  {32'h4514a3f4, 32'h43e221ae, 32'hc32a4fdf},
  {32'hc30656e0, 32'h433e34ba, 32'h4317cf2b},
  {32'h45164c7c, 32'hc19fc7ef, 32'h41dfcafc},
  {32'hc472c45a, 32'hc3bed939, 32'h431f3004},
  {32'h451edae1, 32'h437adf2e, 32'h43c68671},
  {32'hc488362e, 32'hbff352c0, 32'h4373f661},
  {32'h445939e3, 32'h43791849, 32'hc2821cf6},
  {32'hc518c849, 32'h439c8f03, 32'hc209b627},
  {32'h43b0f081, 32'hc33c2416, 32'h439a32dc},
  {32'hc2857da0, 32'h4381f479, 32'h432b88d2},
  {32'h44878dd3, 32'h43a53137, 32'h427b65c3},
  {32'hc48fc9cc, 32'h42a2d39c, 32'h43199c8a},
  {32'h4514e552, 32'hc37d157d, 32'h429e4fb3},
  {32'hc4e11aeb, 32'h42d67bf2, 32'h439d06b9},
  {32'h44474648, 32'hc2232132, 32'hc327f9cb},
  {32'hc3dec2d8, 32'hc2a987ca, 32'hc3ab8398},
  {32'h448694b7, 32'hc3663238, 32'h41e82d5f},
  {32'hc41a2117, 32'hc35c8f32, 32'hc37368a2},
  {32'h4482e638, 32'h42cb2c62, 32'hc34ae472},
  {32'hc4a62461, 32'hc360446d, 32'hc2f3acde},
  {32'h44f1ae03, 32'h42726166, 32'hc3a2551f},
  {32'hc4ccf7be, 32'hc3c3ead7, 32'hc29a37e4},
  {32'h449b7261, 32'hc272a488, 32'h42f07530},
  {32'hc4dbcdcc, 32'h429e0d63, 32'hc2511f76},
  {32'h4413d3d4, 32'h4315b8d2, 32'hc3a16f15},
  {32'hc50934d3, 32'h43b25487, 32'h42ab4f91},
  {32'h43efec2b, 32'hc291fa2f, 32'h418ec899},
  {32'hc4ba1615, 32'h40b7a26f, 32'h40faaa53},
  {32'h44678a56, 32'hc2b2af71, 32'h427652cb},
  {32'hc4e558c3, 32'h43d97a27, 32'h43857204},
  {32'h44977579, 32'h4218a5a9, 32'h43935488},
  {32'hc4efd32a, 32'hc220a260, 32'h42b66a13},
  {32'h44e74c2f, 32'hc2a676c5, 32'hc2fb7d8c},
  {32'hc34298fc, 32'hc3448ca9, 32'hc2ee67c0},
  {32'h44ce0c8e, 32'h427bbccd, 32'h43f0fd82},
  {32'h41c85e80, 32'h43705bbe, 32'hc39dca93},
  {32'h448fd50b, 32'h44089033, 32'hc387d857},
  {32'hc5153aa6, 32'hc2f183f5, 32'hc39b7726},
  {32'h45180caa, 32'hc267a77c, 32'hc27a99b7},
  {32'hc3498000, 32'h4342dcdb, 32'hc2c49082},
  {32'h44f5a972, 32'h42d2ada8, 32'h426f8f58},
  {32'hc3b8bb7c, 32'h442d4a45, 32'hc3e6ef0f},
  {32'h447a9e8c, 32'hc32d2af9, 32'h41c8dd38},
  {32'hc49865a4, 32'h43453e5f, 32'h432efc3b},
  {32'h4398d09a, 32'h434c6893, 32'h42278c82},
  {32'hc4538776, 32'hc2b59975, 32'hc2edb0d4},
  {32'h444b09fa, 32'hc3be9510, 32'h43c082e3},
  {32'hc4601a84, 32'h430c4320, 32'hc3c085b8},
  {32'h44e69ae2, 32'h43e9315f, 32'h42a4ec9b},
  {32'hc42ff20f, 32'hc30f522e, 32'h41de8a89},
  {32'h45022801, 32'h432220aa, 32'h430f8aab},
  {32'hc4f7c9fb, 32'h42f4365e, 32'h42d7a343},
  {32'h44da23cc, 32'h4250711e, 32'h427efd5e},
  {32'hc369183a, 32'hc2009483, 32'hc2eaaf3c},
  {32'h44d123b6, 32'h43996c5d, 32'h431fed76},
  {32'hc3d0393a, 32'hc3b85cd3, 32'hc3ba1e5f},
  {32'h4486c62e, 32'hc405b63c, 32'hc3900e8e},
  {32'hc5036138, 32'hc380d391, 32'hc253120a},
  {32'hc3d1c808, 32'hc25f5a9c, 32'hc2bd6358},
  {32'h44f9b190, 32'h41b2afbf, 32'hc3839c30},
  {32'hc4aecd03, 32'hc1f6b8e6, 32'hc38370ce},
  {32'h44c8f3ca, 32'h42e3439b, 32'h43d039bc},
  {32'hc4d97922, 32'hc2aa788c, 32'hc2bdaae9},
  {32'h44f8486a, 32'h414a264c, 32'h42b3dcbe},
  {32'hc4fea94f, 32'hc130563d, 32'h4314b180},
  {32'h4481c22a, 32'hc2d05d7d, 32'h4340f99c},
  {32'hc36d7f98, 32'h411a7e9c, 32'hc3b098e3},
  {32'h44869f1a, 32'hc3b24766, 32'hc1dd6055},
  {32'hc3d17f14, 32'h4394b696, 32'hc2bc9184},
  {32'h45124e8c, 32'h427ea6ea, 32'hc2f131c3},
  {32'hc3cbccec, 32'hc32111b1, 32'h43674ea4},
  {32'h43e055d7, 32'h43a4f503, 32'h43397057},
  {32'hc2ff9f40, 32'h41f1d453, 32'hc161ed64},
  {32'h447a2f6e, 32'h43477cf5, 32'h4347371e},
  {32'hc47ade26, 32'h43cb2f06, 32'hc3e9d497},
  {32'h44949ee0, 32'hc1f0bb72, 32'h433a4289},
  {32'hc4d562db, 32'h4158c492, 32'hc171c37b},
  {32'h44ef8266, 32'h433f8a57, 32'h426b4a6b},
  {32'hc4840e20, 32'h424c30b1, 32'hc38b606e},
  {32'h42bedd6c, 32'hc21c8c79, 32'h42b31241},
  {32'hc4de3baf, 32'hc2a4b669, 32'hc37c79a2},
  {32'h44174de6, 32'h43c7201e, 32'h42c015c8},
  {32'hc49acbbb, 32'h42a5773f, 32'hc1ea6a22},
  {32'h44e9fb40, 32'h42d72fae, 32'hc2e57eb6},
  {32'hc43493c6, 32'h436c130c, 32'h42a0a9b2},
  {32'h44cff374, 32'hc3d92bce, 32'h43071b00},
  {32'hc500bd6f, 32'hc200c238, 32'hc39ca5f4},
  {32'h433be5e0, 32'h435d300c, 32'hc30b5527},
  {32'hc512a48a, 32'hc3ba4add, 32'h4386bb2d},
  {32'h44d5ed4e, 32'h42b5c6dc, 32'hbea11370},
  {32'hc2dd39b0, 32'h4356759f, 32'h42380312},
  {32'h44fe05b8, 32'hc3a1ca93, 32'h43c934c2},
  {32'hc4cae70a, 32'hc38e3bdd, 32'hc3b35738},
  {32'h44a27f0a, 32'h4344fcc1, 32'hc34377e1},
  {32'hc50a1bb8, 32'h3fe94003, 32'hc407e4ab},
  {32'h447b6e5c, 32'h432fd3ef, 32'h43d2932b},
  {32'hc4b7266d, 32'h41057881, 32'h435f1887},
  {32'h45087b3d, 32'h4350a2d9, 32'h4356dda4},
  {32'hc35f851f, 32'hc2eb996e, 32'hc38e5426},
  {32'h4525a422, 32'h43b21755, 32'hc3b67020},
  {32'hc5179508, 32'h430faed8, 32'hc28d4f8a},
  {32'h444a58b2, 32'h42362e64, 32'h438d68af},
  {32'hc50fa192, 32'h4386d163, 32'hc31910ec},
  {32'h44b4fc82, 32'h434311f1, 32'hc136efbf},
  {32'hc49fdd5b, 32'h402c9384, 32'h4222635d},
  {32'h44c751f3, 32'h420edb22, 32'hc3550cf9},
  {32'hc5042b1b, 32'hc321ae4f, 32'hc25ae9f6},
  {32'h440e5022, 32'h433154c4, 32'h44138cd6},
  {32'hc5014da3, 32'h425d7413, 32'h43a6a8a6},
  {32'h44946102, 32'h431aeed1, 32'h4229c655},
  {32'hc50f4261, 32'h43603357, 32'h420659e5},
  {32'h44a3aa79, 32'h43b74cdc, 32'h42a69bc2},
  {32'hc4f655db, 32'hc341e778, 32'hc3798e81},
  {32'h4504325c, 32'h4224b210, 32'hc3af5351},
  {32'h42e2aba2, 32'hc33f3e45, 32'hc130ad27},
  {32'h440c690b, 32'h42e1445b, 32'hc27d593f},
  {32'hc51d0b89, 32'hc16ec570, 32'hc24cbf56},
  {32'h44a5a753, 32'hc2d45383, 32'h43330f7d},
  {32'hc4add8c9, 32'hc21aa85f, 32'hc2397ed8},
  {32'h43ada7f8, 32'h42898a57, 32'hc39d4a40},
  {32'hc3515408, 32'hc201df1e, 32'hc32cb95d},
  {32'h4521048e, 32'h434de82a, 32'h42e1e9e3},
  {32'h427172ec, 32'h431d9fbb, 32'hc2a3155e},
  {32'h4424de50, 32'h435ca264, 32'h428e972a},
  {32'hc383f270, 32'h43107389, 32'hc2fe661b},
  {32'h44fb4bb9, 32'hc37b40b4, 32'h432279f4},
  {32'hc4ff9955, 32'hc2b05b14, 32'hc20b5350},
  {32'h43e91faa, 32'hc01ee255, 32'h42b2c52e},
  {32'hc4beaebd, 32'hc341c94c, 32'h435e8c35},
  {32'h44a9f136, 32'hc3344dc5, 32'h426f1767},
  {32'hc4c5214f, 32'h43a643a7, 32'hc3545157},
  {32'h4500ef5a, 32'h4349b698, 32'hc35947ab},
  {32'hc51a9372, 32'h42d2f8de, 32'hc3b43e5a},
  {32'h4481d0f5, 32'h438c56ac, 32'h43127b61},
  {32'hc4bc74db, 32'h4383e939, 32'hc29dd807},
  {32'h44287b1a, 32'hc259cba4, 32'h426fa5dc},
  {32'hc4d83065, 32'h408fc006, 32'h43286cfd},
  {32'h44fe5496, 32'hc222d48d, 32'h43c61b54},
  {32'hc4e1cbdc, 32'hc32934e2, 32'hc397e2b5},
  {32'h4381c934, 32'hc2da173f, 32'h4316be15},
  {32'hc4b51f84, 32'h4382c8a7, 32'hc307c4a5},
  {32'h44b84a5e, 32'h4408356a, 32'hc40a8624},
  {32'hc3b43d28, 32'hc33860a3, 32'hc353ff3f},
  {32'h44a6e0e0, 32'h4301f9b0, 32'h4222bd93},
  {32'hc4b6fa7f, 32'h42473fb2, 32'h429b806d},
  {32'h44c1840f, 32'h43deaedd, 32'hc396aabc},
  {32'hc4f8d11e, 32'hc308b237, 32'h43ae9267},
  {32'h44013c04, 32'h41a88642, 32'hc38e9ef7},
  {32'hc39aa92f, 32'h42057b1f, 32'h43a4fc74},
  {32'h44cfd852, 32'h42121a20, 32'h4333245e},
  {32'hc4b08486, 32'hc265113b, 32'h4223f754},
  {32'h44895a9d, 32'hc2660184, 32'h43e673b0},
  {32'hc465eef2, 32'h43b51ed5, 32'h44096001},
  {32'h44ac608f, 32'hc3250f33, 32'h43a9bcca},
  {32'hc45d6db4, 32'hc32b6640, 32'h438d4959},
  {32'h450040ae, 32'h4395c8b0, 32'hc2914659},
  {32'hc4fa2877, 32'h43a5d8ab, 32'hc139b83d},
  {32'h447bc402, 32'hc394b748, 32'hc1598dc7},
  {32'hc3c05699, 32'hc3c82b5e, 32'h43aa6575},
  {32'h441eec7c, 32'h43d8a905, 32'h41e9027e},
  {32'hc5073a2f, 32'h40c170dc, 32'hc33facd6},
  {32'h43c4bd78, 32'hc2c18eae, 32'h41b75857},
  {32'hc496779f, 32'h42e63ab4, 32'hc1ae28fe},
  {32'h44e8663e, 32'hc3a5ad88, 32'h438b1504},
  {32'hc360a196, 32'h40abae77, 32'hc3928f49},
  {32'h44421ff7, 32'hc40de575, 32'hc2a8c042},
  {32'hc4886419, 32'h42b4ed1b, 32'h42701a44},
  {32'h44ed5d8d, 32'h43d0ea4d, 32'h42a4ab49},
  {32'hc3fe1d98, 32'h42b788bf, 32'h432e68f7},
  {32'h448b6db9, 32'hc3017b6a, 32'hc3c767cc},
  {32'hc4cb36ae, 32'h42510466, 32'h431dad9f},
  {32'h4421e4b8, 32'hc31ae484, 32'h439f72c2},
  {32'hc4d7e57a, 32'h43c70739, 32'h43851e67},
  {32'h44a5131f, 32'hc3115ff0, 32'hc3816ec4},
  {32'hc503ae62, 32'h42a60b8d, 32'h42de2719},
  {32'h44169b7a, 32'hc03a4726, 32'h42a7b9e4},
  {32'h42b0d8f0, 32'hc300c144, 32'h440344ae},
  {32'h44d3455c, 32'h431beffd, 32'h430685e6},
  {32'hc5126b86, 32'hc2986765, 32'h41a45022},
  {32'h440356c0, 32'h43c90ff0, 32'h43db6aed},
  {32'hc3c48ed0, 32'hc3298e64, 32'h439df4c2},
  {32'h44e422a0, 32'hc2ee41b3, 32'h4320dab5},
  {32'hc4551d20, 32'h42f01499, 32'h4314c366},
  {32'h44cf130f, 32'h42cb6010, 32'hc1e3a529},
  {32'hc45ccd00, 32'h4341a9e8, 32'hc33047ec},
  {32'h44c7a8d8, 32'h42a8cfca, 32'hc2ed1381},
  {32'hc43129e7, 32'h432bac2c, 32'hc304bcc2},
  {32'h44771aee, 32'h430b3d48, 32'hc31fdc5b},
  {32'hc32cd308, 32'hc2101c18, 32'h43171a11},
  {32'h447aff60, 32'h41ef37d2, 32'h43daab3f},
  {32'hc4aac38e, 32'h43055d21, 32'hc34dcfaa},
  {32'h45027e3c, 32'hc34f2779, 32'h436887d9},
  {32'h43420ca0, 32'hc2304141, 32'hc320fa70},
  {32'h42c566c0, 32'h430f2ed0, 32'h42e01d33},
  {32'hc50c5228, 32'hc2188202, 32'h42662abb},
  {32'hc234f148, 32'h4310a931, 32'hc36312d6},
  {32'hc46d90aa, 32'h432fa488, 32'hc10ee811},
  {32'h44e2a21d, 32'hc422c917, 32'hc17fb158},
  {32'hc3e532c8, 32'hc24b9f68, 32'hc2898368},
  {32'h450191de, 32'hc34cd9e4, 32'hc1db7a31},
  {32'hc435d9ac, 32'h42f55489, 32'h4375416d},
  {32'h4453d034, 32'hc33caaa1, 32'hc3d56af3},
  {32'hc4751880, 32'hc26c1166, 32'h4383e975},
  {32'h44ec1801, 32'hc13eb100, 32'hc2919648},
  {32'hc4a7433a, 32'hc22bb7c9, 32'h432823b7},
  {32'h444a6ea0, 32'h42420a81, 32'hc300ef1b},
  {32'hc4f95e83, 32'hc345ff06, 32'h43593f79},
  {32'h43a89a3c, 32'h43a5e343, 32'hc33b3b3a},
  {32'hc333a481, 32'hc244f81a, 32'h436ccfd4},
  {32'h45090cc0, 32'h42c2c48b, 32'hc2ef4b76},
  {32'hc4f6fe44, 32'h43d86f2d, 32'hc14cb72e},
  {32'h45171882, 32'h41bfb8d4, 32'hc30841e1},
  {32'hc494052b, 32'h41bae0c3, 32'hc30df53d},
  {32'h44b3d3a8, 32'h430ef251, 32'h43d210cc},
  {32'hc4b95355, 32'hc20ff4e4, 32'h42c47655},
  {32'h44212704, 32'hc35c3b45, 32'h43f29f27},
  {32'hc42439a6, 32'h432bf59c, 32'h4219ee36},
  {32'h442334b7, 32'h4365fad7, 32'h43f3ff51},
  {32'hc44744c4, 32'h42650d3c, 32'h431dc2bf},
  {32'h4482671e, 32'h43b7cee5, 32'hc3cc545f},
  {32'hc4bfe3a0, 32'h4109a9b6, 32'hc3696f56},
  {32'h4451af03, 32'h431ebdb2, 32'hc2485182},
  {32'hc49d6e1b, 32'hc2ad8789, 32'hc3a3c14a},
  {32'h44dcebf2, 32'h4369ad95, 32'h43421126},
  {32'hc4b41147, 32'h4394ab8a, 32'hc311e400},
  {32'h4509356c, 32'hc3a7a819, 32'hc2fc73b4},
  {32'hc505e962, 32'h435c185e, 32'hc3bf0d3c},
  {32'h4389f754, 32'hc395e893, 32'h429a0fe5},
  {32'hc4a1d360, 32'h439f4597, 32'hc33c6b2a},
  {32'h44c7b3de, 32'h42e7036d, 32'h40f1d610},
  {32'hc50b5f12, 32'h41e91b4c, 32'h435ecaa4},
  {32'h4498f430, 32'hc20ec560, 32'hc383f8d3},
  {32'hc4a9d7f5, 32'h43118622, 32'hc38f1198},
  {32'h426836a0, 32'h420afce8, 32'hc1850a24},
  {32'hc4ec0dbc, 32'hc3ca71ab, 32'hc3c0b9d3},
  {32'h44f2ba89, 32'hc3678686, 32'hc2cad670},
  {32'hc4a21f66, 32'h431ce996, 32'hc354e9fb},
  {32'h4481d874, 32'h437b3b7a, 32'h433b69e1},
  {32'hc3aa4460, 32'h43716ac8, 32'hc22d567c},
  {32'h44bcff4e, 32'hc2a56895, 32'h42bdad11},
  {32'hc3f3f282, 32'h42c42a2e, 32'hc37dfbf2},
  {32'h44abf126, 32'h42af1239, 32'hc26f0f46},
  {32'hc238da60, 32'hc1e24db6, 32'h430950d0},
  {32'h442a8a75, 32'hc30e48be, 32'hc3b01ccf},
  {32'hc47c389a, 32'h43e0a1bb, 32'hc3283912},
  {32'h44f6336e, 32'hc34fb05c, 32'hc2b3450b},
  {32'hc4ea788b, 32'hc34ec38d, 32'hc340043b},
  {32'h443fe04d, 32'hc187db68, 32'hc40c3dc9},
  {32'hc4313908, 32'h436a7a68, 32'h432a3148},
  {32'h44db772c, 32'hc3810056, 32'h427e2dd4},
  {32'hc4bc4fe6, 32'h43053780, 32'h42caf4b6},
  {32'h44bcc3e2, 32'h41a0996c, 32'h4299eb84},
  {32'hc4579528, 32'h43b649a9, 32'hc292daa5},
  {32'h43fab0d4, 32'hc3552b1b, 32'h40639da9},
  {32'hc31ae17e, 32'h43343932, 32'h420ec874},
  {32'h450ca77d, 32'hc3bde4b6, 32'h4392f937},
  {32'hc4578366, 32'h438de758, 32'h4306b08a},
  {32'h44699dda, 32'h43d20641, 32'h438563d6},
  {32'hc429c700, 32'hc4138c22, 32'h418108be},
  {32'h44a22676, 32'h41cc1083, 32'hc2b6e749},
  {32'hc45ea6e1, 32'h436ca0ba, 32'hc38643d0},
  {32'h441c07a6, 32'hc288fee8, 32'hc3fb7f76},
  {32'hc50f2cd6, 32'hc377c4e4, 32'hc33a7fd4},
  {32'h438fd200, 32'hc2915893, 32'hc307d2bf},
  {32'hc3e5b445, 32'h42cf74be, 32'h429c8260},
  {32'h44db9c4f, 32'h43278351, 32'hc3696d7d},
  {32'hc316fbdf, 32'h42fb427a, 32'hc2968d87},
  {32'h451a9258, 32'hc08516ac, 32'hc3d209d0},
  {32'hc50c7d42, 32'h424c6223, 32'h4346570e},
  {32'h4485e762, 32'hc40da36e, 32'hc4808434},
  {32'hc3594a48, 32'hc33c3119, 32'hc363a9b3},
  {32'h44a3a7c6, 32'hc3db95ff, 32'h42e15446},
  {32'h433c41f7, 32'h4230c661, 32'h42347715},
  {32'h44b56350, 32'h42e59fe0, 32'h43b3b153},
  {32'hc4cac110, 32'h431b712e, 32'h42b8e4d6},
  {32'h44ce64ec, 32'h4304b5ce, 32'h43819009},
  {32'hc41ff7f6, 32'hc2830ea0, 32'hc2636d7a},
  {32'h44781d62, 32'h43809c98, 32'hc33380c8},
  {32'hc4fce432, 32'hc2d6e588, 32'h421c37ee},
  {32'h451951ba, 32'h42c8f8e2, 32'hc2c3d5f9},
  {32'hc50581df, 32'hc2bd96f2, 32'h436450b8},
  {32'h43be1e34, 32'h4226254b, 32'hc1a5f5fe},
  {32'hc48c658e, 32'hc073c8e8, 32'hc2887cb8},
  {32'h44c5ebcc, 32'h43031eb7, 32'h430444b5},
  {32'hc4841252, 32'h4318998c, 32'h420db1ea},
  {32'h447a9bea, 32'h42fcbdf1, 32'hc395d2a2},
  {32'h43255084, 32'hc0ee1ea7, 32'hc382c633},
  {32'h44c8b37f, 32'hc3b2831c, 32'h42de962a},
  {32'hc4b4c223, 32'h4216783e, 32'hc25bee7a},
  {32'h44f3359c, 32'hbff684dd, 32'hc3c67efb},
  {32'hc4be0813, 32'h438b20f1, 32'hc3748d8c},
  {32'h450845c1, 32'hc36ecd80, 32'h43c21ab3},
  {32'hc2c856a0, 32'h438b84bf, 32'h432a6165},
  {32'h44b5b7d8, 32'hc21fe4f2, 32'hc3266402},
  {32'hc4d6cfc0, 32'h43694c49, 32'h421957c8},
  {32'h449210a9, 32'hc38aa6b2, 32'hc393d1d7},
  {32'hc47f20b9, 32'hc31e70d7, 32'hc341edd7},
  {32'h445cf3c3, 32'hc287696a, 32'hc329ad01},
  {32'hc4d47cc0, 32'hc18bb20d, 32'hc3b1a204},
  {32'h4493ef61, 32'h436e3232, 32'hc3ff70bf},
  {32'hc49240b2, 32'h418bec88, 32'h42e9ec60},
  {32'h44faf4cd, 32'hc3052273, 32'h41aae895},
  {32'hc50482f0, 32'h431b18f6, 32'hc2abbd9c},
  {32'h44f5065a, 32'h42b7d4a7, 32'h42225a87},
  {32'hc5055c41, 32'hc344e47f, 32'h431db181},
  {32'h44e3ad96, 32'hc2a7a39d, 32'h4183549b},
  {32'hc45cb432, 32'hc3768224, 32'h4370d30b},
  {32'h443fedaa, 32'hc3c86931, 32'hc287b07e},
  {32'hc40f99a4, 32'h434cb918, 32'hc22a2afb},
  {32'h44c7f880, 32'hc0bf142c, 32'h430552d9},
  {32'hc3a71dac, 32'h43828e3c, 32'h417bfcae},
  {32'h44bd0463, 32'h43503590, 32'hc299c9dd},
  {32'hc49975d9, 32'hc341f75a, 32'hc2ce4eed},
  {32'h44a1dcc9, 32'h41f90f35, 32'hc33e92d6},
  {32'hc3bc6e20, 32'h405a6920, 32'h439d57d7},
  {32'h45032203, 32'hc3511d5d, 32'hc352c939},
  {32'hc471439c, 32'hc2209c65, 32'hc3c9cafb},
  {32'h4504fef2, 32'h43f71117, 32'hc2b7d936},
  {32'hc3dfcb68, 32'hc330d70e, 32'h43464f84},
  {32'h43a30adc, 32'hc3d46ef0, 32'h43697112},
  {32'hc502fbad, 32'h43b88506, 32'hc342beaf},
  {32'h43f9d4d0, 32'hc29c2070, 32'hc32c39ad},
  {32'hc45ac7a8, 32'hc2fbf466, 32'h42cfd8b5},
  {32'h44017226, 32'h420d622c, 32'hc371b79e},
  {32'hc50c3710, 32'hc373d469, 32'hc04f7cea},
  {32'h44ce210a, 32'h434acf63, 32'h41f66d3c},
  {32'hc41758cc, 32'h4330047b, 32'hc14b614c},
  {32'h44592e4e, 32'hc2dccba1, 32'hc2e6dec3},
  {32'hc4ec62dc, 32'hc3085903, 32'h42df9dbe},
  {32'h44fe5c23, 32'h41c92fe6, 32'hc344228a},
  {32'hc3a07474, 32'hc2cfc496, 32'hc3a796bc},
  {32'h4434ff6a, 32'hc2e4ba81, 32'h41cf3600},
  {32'hc3e677ec, 32'h43a644dd, 32'hc3ae8de8},
  {32'h442866db, 32'hc199a7d4, 32'h4382ad7a},
  {32'hc3c48618, 32'h42eb86b3, 32'hc3e696c4},
  {32'h42ed8270, 32'h426895f0, 32'h429a80ba},
  {32'hc506ea5f, 32'hc37dc021, 32'h435812e3},
  {32'h451989a0, 32'h42208f68, 32'h436bb11c},
  {32'hc4f40f02, 32'h43cf7afb, 32'hc2dfc502},
  {32'h44ebef98, 32'hc2e27c68, 32'hc1fd9d62},
  {32'hc484f324, 32'hc29df00f, 32'hc0f834fc},
  {32'h442ce306, 32'hc323dde8, 32'hc25f9f87},
  {32'hc3d062f0, 32'h43bfae27, 32'hc402a2f2},
  {32'h44c8dd21, 32'hc39c54a8, 32'h428fefbe},
  {32'hc39cc844, 32'h40e3049d, 32'hc3974700},
  {32'h44305790, 32'hc3b954c0, 32'hc2e1b15f},
  {32'hc432347e, 32'hc31e1e59, 32'h42b81b99},
  {32'h449b4d46, 32'h43137f18, 32'h439d5ce8},
  {32'hc5151fb4, 32'hc2029a7d, 32'h4249c4e1},
  {32'h4475ee62, 32'h4183b29c, 32'hc2db0b28},
  {32'hc4ab941d, 32'h432bbed4, 32'h438fe5f7},
  {32'h450eb692, 32'hc3b787b3, 32'h43bf158f},
  {32'hc457dc65, 32'hc36c60c2, 32'hc3320181},
  {32'h44cc71c0, 32'hc379e123, 32'h42d47734},
  {32'hc407e4bc, 32'h42666a5c, 32'hc31761e6},
  {32'h45163d0e, 32'hc3040296, 32'h439d5e17},
  {32'hc50e1746, 32'h404ed819, 32'h4332a099},
  {32'h4454c7b4, 32'h425d7ad3, 32'hc2d053db},
  {32'h4333edf0, 32'hbfb47418, 32'hc31b7dbd},
  {32'h44c2fc84, 32'hc0c6c3ac, 32'h43565c1a},
  {32'hc2c695a0, 32'h431de2ae, 32'h43f26273},
  {32'h43ecf30c, 32'hc3499a2a, 32'hc26d1eb1},
  {32'hc3d77668, 32'hc4131504, 32'h4391c91c},
  {32'h43af2070, 32'h43f7359a, 32'h431f4937},
  {32'hc50c7fda, 32'hc2b621ae, 32'hc0a1fde2},
  {32'h439b0cd8, 32'h4360159e, 32'hc35b436a},
  {32'hc3a5f312, 32'hc358ab3d, 32'h433dcabc},
  {32'h450b1830, 32'h40bfdd70, 32'h43b2f456},
  {32'h4349a7bf, 32'h43b3e8f6, 32'h439d321f},
  {32'h44cdb5c3, 32'h42836281, 32'hc22f1f04},
  {32'h40ef6c00, 32'hc1b2042f, 32'h43c34311},
  {32'h442cef88, 32'h43963bd4, 32'h43614de9},
  {32'hc4336898, 32'h432ce42b, 32'hc3a82e9d},
  {32'h44863b8b, 32'hc2a0c1a8, 32'hc2385799},
  {32'hc4d275b4, 32'h42aa1b4a, 32'hc3f8438a},
  {32'h438e90ba, 32'h44023e76, 32'h439fc33a},
  {32'hc4a73f87, 32'hc367b8b4, 32'hc3216da0},
  {32'h445618fa, 32'hc272e921, 32'h40bd5c2c},
  {32'hc43e2308, 32'hc396854a, 32'hc403e905},
  {32'h438e086f, 32'hc3983285, 32'hc1cb47cf},
  {32'hc3923730, 32'hc3ca2e76, 32'hc3216471},
  {32'h42caa0e4, 32'hc40cdfc8, 32'h4282ef27},
  {32'hc4aedc71, 32'h434fac34, 32'hc3a5f739},
  {32'h447b3ec4, 32'hc3360b82, 32'hc3df48d6},
  {32'hc4725066, 32'hc36da534, 32'h430b88a9},
  {32'h4421530e, 32'h43326d5a, 32'h430a8807},
  {32'h428c32b3, 32'h439c4218, 32'h41824389},
  {32'h44408364, 32'h433884c6, 32'h43a02cb3},
  {32'hc3a0255f, 32'h41b3b0f3, 32'hc335f07a},
  {32'h438de41e, 32'h429dc5ae, 32'h42e125fc},
  {32'hc46a1154, 32'hc2d9a099, 32'h422d28b2},
  {32'h44eca15a, 32'hc36c8a23, 32'hc37a47b2},
  {32'hc3f2b806, 32'h41a4dc8d, 32'hc26d04f4},
  {32'h45079262, 32'h43bdfc44, 32'hc31949a6},
  {32'hc42edf16, 32'h434df17a, 32'hc410dbcf},
  {32'h449e0bf0, 32'h42ba54b3, 32'h429d35aa},
  {32'hc439441e, 32'h4387fd2e, 32'h42d0bc59},
  {32'h4487e009, 32'h439cc875, 32'h4337b501},
  {32'hc4f80cd5, 32'h431c87f6, 32'h43c63083},
  {32'h44afda01, 32'hc27418e7, 32'hc28acefc},
  {32'hc1f9e6fe, 32'h434afff0, 32'hc28e1f84},
  {32'hc250efa0, 32'hc2caca17, 32'hc2fbe37a},
  {32'hc4d8e28b, 32'h42d6444c, 32'h40a8dda0},
  {32'h4436b988, 32'h4387d76d, 32'h4325c580},
  {32'hc3b9b421, 32'hc3b78b09, 32'h433d8737},
  {32'h4326a22c, 32'hc16f224d, 32'hc28072f1},
  {32'h418ee6bc, 32'hc3134dcb, 32'hc3932e46},
  {32'h44234b32, 32'h42e32194, 32'hc27161fa},
  {32'hc4d384c2, 32'h438e69e4, 32'hc13e4819},
  {32'h45259757, 32'hc3546184, 32'h422a94c8},
  {32'hc5217d2d, 32'h43a2a9fb, 32'h41cd6357},
  {32'h436c1528, 32'h42880354, 32'h41acbd41},
  {32'hc32249a8, 32'h43b78f03, 32'hc1731546},
  {32'h44f7b148, 32'hc21b1342, 32'h43b23daa},
  {32'hc4987446, 32'h41a17b56, 32'hc30f272a},
  {32'h44ae1352, 32'hc30c0a3e, 32'hc29b1107},
  {32'h4260de10, 32'h405e0ab8, 32'h41b7b414},
  {32'hc329b608, 32'hc385727a, 32'h42808cad},
  {32'hc4a73728, 32'h437a8947, 32'h4271294b},
  {32'h450307ea, 32'h42d0c74e, 32'h433aa3e3},
  {32'hc4e9dd62, 32'h41400ee3, 32'hc2a34615},
  {32'h44d01461, 32'hc2978690, 32'hc2b0cd36},
  {32'hc5004e9a, 32'hc380a707, 32'h43d71eac},
  {32'h448ae0cb, 32'h436a9cbf, 32'hc36812fc},
  {32'hc4e1254c, 32'hc2275198, 32'hc26a1a99},
  {32'h4388585e, 32'h433f65f9, 32'hc3ade25c},
  {32'hc4d6cf1e, 32'hc2323e86, 32'h43822043},
  {32'h4494ec5e, 32'h413f08bd, 32'hc229d406},
  {32'hc435b040, 32'hc13007e8, 32'h435eadad},
  {32'h44fcc3cb, 32'hc350db2e, 32'h43004ae8},
  {32'hc4f9017d, 32'h42733b69, 32'hc2270875},
  {32'h43d0ab78, 32'hc1975c6a, 32'h42a00a92},
  {32'hc4dddf86, 32'hc3b3abbd, 32'h43404d0a},
  {32'h44c4b75c, 32'hc37ff285, 32'h4219b911},
  {32'hc3f4a751, 32'hc23da648, 32'h423bbbd2},
  {32'h44fd138a, 32'hc37948b8, 32'hc2aae59d},
  {32'hc4e5f0de, 32'h43819f96, 32'hc33f3862},
  {32'hc270d744, 32'h4388cc00, 32'hc2f1935f},
  {32'hc452889d, 32'hc1d744c4, 32'hc392dfc8},
  {32'h434bae74, 32'h41ed769f, 32'h4299c48c},
  {32'hc4d522c0, 32'h42bf2927, 32'h41934fab},
  {32'h43a41399, 32'h434d1173, 32'h402424e5},
  {32'hc4804237, 32'h433d12f6, 32'h43b03a54},
  {32'h445efaa2, 32'h41704194, 32'h42c335cb},
  {32'hc438ec82, 32'hc2cb3f37, 32'h419811b8},
  {32'h44aefead, 32'hc2e3beba, 32'h43a0c856},
  {32'hc4dc5b9a, 32'h442e22f7, 32'h44062485},
  {32'h44c4cd36, 32'hc0f1d9f2, 32'hc32037da},
  {32'hc486286f, 32'h3f2cc900, 32'h42b8c9fa},
  {32'h44be9cf8, 32'hc0dc88d5, 32'h431a8ced},
  {32'hc3d1b8f0, 32'hc39aced2, 32'hc2afc45c},
  {32'h44b72c6f, 32'h42eb5af8, 32'hc360f463},
  {32'hc500488e, 32'hc2a996e8, 32'h43675384},
  {32'h43927096, 32'hc3415713, 32'hc32004a2},
  {32'hc4af0cde, 32'hc2724394, 32'hc348aea5},
  {32'h43c1b180, 32'hc3c7e43b, 32'hc303ba3c},
  {32'hc4613e3a, 32'h43880b82, 32'h43582205},
  {32'h44ea1830, 32'hc2cf9295, 32'hc39cb6cb},
  {32'h428b2e40, 32'hc2752ee6, 32'hc393778c},
  {32'h440438dc, 32'hc35b554e, 32'hc35c761a},
  {32'hc3eb2878, 32'h41db7d9a, 32'h428f88ed},
  {32'h44ffe2ff, 32'hc319bcf1, 32'hc30d021e},
  {32'hc49cfa99, 32'h43345b65, 32'h433ef51a},
  {32'h44d6e63c, 32'hc1ac8f64, 32'hc374b029},
  {32'hc4f828fe, 32'h43427264, 32'h42256cd6},
  {32'h4417da25, 32'hc3007daf, 32'hc34c5a36},
  {32'hc4b8985f, 32'h439b182b, 32'h437fc2e7},
  {32'h4501b251, 32'hc2a56d76, 32'hc293c472},
  {32'hc4c9a945, 32'hc275b6e0, 32'hc3a98b3e},
  {32'h4504ae6c, 32'hc3706994, 32'h416f89ba},
  {32'hc4594fa8, 32'hc32770eb, 32'h42743d24},
  {32'h44aed46d, 32'hc38b6f7e, 32'hc1b7513e},
  {32'hc4bc86a0, 32'hc15ba36c, 32'h4347e92a},
  {32'h44974a8e, 32'h424f8346, 32'hc1d4aa09},
  {32'hc4e2ceb6, 32'hc370827b, 32'h4385c4a5},
  {32'h4457a236, 32'hc2bfe272, 32'h428c4b32},
  {32'hc3a9dffc, 32'h41de6fb8, 32'h41cab0ae},
  {32'h44575f0f, 32'hc2898e6a, 32'hc2eda351},
  {32'hc4afc6d2, 32'hc2cc8ca9, 32'hc32a6952},
  {32'h44615b74, 32'h431f408f, 32'hc2d377ec},
  {32'hc4a2a749, 32'hc29dc791, 32'h43b52c05},
  {32'h44b47c2d, 32'h43754863, 32'hc2421c48},
  {32'hc4d62932, 32'h41e67398, 32'hc248fcdb},
  {32'h450017d5, 32'h436df0cc, 32'hc3a87a11},
  {32'hc4ec493d, 32'h4330644f, 32'h430e0594},
  {32'h44f95f56, 32'hc29cfdc1, 32'h42826560},
  {32'hc3d158b0, 32'h435782e4, 32'h435da0fc},
  {32'h442636ca, 32'hc3ec3013, 32'h4348064f},
  {32'hc38c37fe, 32'h4323209c, 32'h439d6ce7},
  {32'h43df95d0, 32'hc39991eb, 32'h436ca806},
  {32'h4407fb20, 32'h43044642, 32'hc3816d55},
  {32'hc48dd63d, 32'h43509b76, 32'h438af2a4},
  {32'h44bcb526, 32'h4398f2b4, 32'hc2d137fe},
  {32'hc4d190ef, 32'hc25d1214, 32'h429a3d94},
  {32'h44ae427b, 32'hc3ad7c56, 32'hbff9ea8f},
  {32'hc494f042, 32'h42eed305, 32'h42bdaaf6},
  {32'hc20a3c40, 32'h440c5a9d, 32'hc39745e6},
  {32'h43871730, 32'hc32bc448, 32'h4360f612},
  {32'h44ccab46, 32'hc359c386, 32'hc2b21972},
  {32'hc4c43105, 32'hc3b487a2, 32'h42e82880},
  {32'h44a6e965, 32'hc3b9d19f, 32'hc332a74e},
  {32'hc48579f9, 32'h41497c32, 32'h436fbba6},
  {32'h43d5e133, 32'hc123c45e, 32'h42e5483c},
  {32'hc42c58ab, 32'h42eaf904, 32'hc32bf036},
  {32'h4485af99, 32'h43407c8c, 32'h43813d70},
  {32'hc48c33eb, 32'h43d32487, 32'h434373d2},
  {32'h44f7517c, 32'h43a09266, 32'hc320964c},
  {32'hc427b6db, 32'h42de2d4d, 32'h439ece53},
  {32'h4507c072, 32'hc2c856f5, 32'h429bc9f8},
  {32'hc4dc7717, 32'hc34102c2, 32'h400538ce},
  {32'hc27fbea3, 32'h41217268, 32'h3faf02b2},
  {32'hc419a5d0, 32'h4349d659, 32'hc303fbd5},
  {32'h44e0d668, 32'hc2d06a8a, 32'h425004c3},
  {32'hc36a25e0, 32'hc330c432, 32'h43747949},
  {32'h447b70a6, 32'h4307efa5, 32'hc3913fcd},
  {32'hc483d4aa, 32'hc36149c5, 32'h420bc4a1},
  {32'h44c2a37f, 32'hc3aadbd2, 32'hc3bfa227},
  {32'hc3c163b0, 32'hc10aa89b, 32'hc3ff6aeb},
  {32'h4501649a, 32'h435cda7b, 32'hc242bf3d},
  {32'hc2168680, 32'hc061bfec, 32'hc28e3f56},
  {32'h44772a53, 32'hc34937c8, 32'hc25269fd},
  {32'hc3faddda, 32'hc33136f0, 32'hc3e2032c},
  {32'h44be51be, 32'hc33069f3, 32'h4424fe8d},
  {32'hc44ee75e, 32'hc2d01067, 32'hc2fff28e},
  {32'h447ef7fc, 32'h438d354d, 32'hc30952a7},
  {32'hc4239dbf, 32'hc2fefa53, 32'h4421ea25},
  {32'h44ca2ee0, 32'hc1c616a0, 32'h426c4870},
  {32'hc4b4f582, 32'hc394c6fb, 32'h43caecbd},
  {32'h4510dc7f, 32'h439d8757, 32'hc36b5ed9},
  {32'hc50d0ecb, 32'h43cbb184, 32'hc3988e36},
  {32'h44b2e3c9, 32'h42f09945, 32'h43e4035b},
  {32'hc2fff01a, 32'h439d4d8b, 32'hc35e85d9},
  {32'h450a47e9, 32'hc2fd0e1c, 32'h42e46abb},
  {32'hc4524d7d, 32'h4350a76e, 32'h4387e783},
  {32'h4387f34c, 32'h433f2aa8, 32'h41fa507c},
  {32'hc4da5ede, 32'hc1b8730f, 32'h43105fa1},
  {32'h44902e73, 32'h3f535ae0, 32'h43a7eb01},
  {32'hc4137400, 32'hc34920bf, 32'hc21de794},
  {32'h448b4a88, 32'h42c7927a, 32'h426744e2},
  {32'hc4254b5c, 32'hc39b0393, 32'hc205021e},
  {32'h42c8beca, 32'hc23dd528, 32'hc0ff7bbd},
  {32'hc4b4a1f0, 32'h428d69cb, 32'hc29cc728},
  {32'h4516cc0a, 32'hc37e9839, 32'hc2ac4528},
  {32'hc4985fd7, 32'h4303743f, 32'hc34744fc},
  {32'h41ab28d0, 32'h436bdef8, 32'hc371f1ca},
  {32'hc4426dff, 32'h434bd817, 32'h419bb345},
  {32'h43f97b24, 32'hc2c4ea4a, 32'h430ee66b},
  {32'hc50a12ad, 32'h426602ae, 32'hc2ee8b92},
  {32'h446ff65c, 32'h432a4b66, 32'hc0c27880},
  {32'hc4c885e8, 32'hc361722a, 32'hc3c2af1a},
  {32'h42aac170, 32'h42d28881, 32'h433fc22a},
  {32'hc507386d, 32'hc1f37654, 32'h43b70e21},
  {32'h44d29a07, 32'hc3433270, 32'h42c44379},
  {32'hc4a05c1b, 32'h42902345, 32'h42a1aab4},
  {32'h440bae55, 32'h42f6496a, 32'h43a32ffc},
  {32'hc4af0fa1, 32'hc38e063f, 32'hc2fac261},
  {32'h44522f50, 32'hc1568912, 32'h43193f46},
  {32'hc50b11ec, 32'h40bdc21c, 32'hc39b655d},
  {32'h442d364c, 32'h43a8a799, 32'h4250387e},
  {32'hc2b67dd0, 32'h409a0418, 32'hc3ccfbd3},
  {32'h44444b4a, 32'h43a4468c, 32'hc2e76736},
  {32'hc5018f22, 32'hc34f5370, 32'h42846846},
  {32'h4500e668, 32'hc29b97e4, 32'h421a2eaf},
  {32'hc5006c50, 32'h43b5cc05, 32'h43861068},
  {32'h44a06490, 32'h42f5b5d6, 32'hc21f2b41},
  {32'hc4930f5e, 32'h43f8d4ca, 32'hc398c68f},
  {32'h4502df38, 32'h42a724da, 32'hc3edf3a4},
  {32'hc4bc16ce, 32'h42e0b31a, 32'h42fb236e},
  {32'h44f1c7bf, 32'hc3775dbd, 32'hc3a345e9},
  {32'hc50dd2c5, 32'h42953e0d, 32'h43382270},
  {32'h448ff529, 32'hc1e2d5eb, 32'h420bb65d},
  {32'hc3acc774, 32'hc087cdb0, 32'hc39ca06c},
  {32'h44bac108, 32'hc2a275df, 32'hc3237384},
  {32'hc4b8b98a, 32'h4435041d, 32'hc27259b6},
  {32'h44c6a2ed, 32'hc352e8b1, 32'h428b5bf3},
  {32'hc3132a90, 32'hc2e55790, 32'h42aec7fa},
  {32'h44c2f503, 32'hc2353e50, 32'h430a0b56},
  {32'hc4897ee1, 32'hc3095fb1, 32'hc3864e2f},
  {32'h445c3181, 32'hc1c474e1, 32'hc24a6d71},
  {32'hbf365000, 32'hc2baff77, 32'h43b08909},
  {32'h45086fde, 32'hc27c577c, 32'hc324349d},
  {32'hc4df2b7d, 32'h4186cd3e, 32'hc233069c},
  {32'h438968a2, 32'h4342c18f, 32'h42f3382b},
  {32'hc34cb0ad, 32'h4325256e, 32'h430e01c8},
  {32'h4460ae5d, 32'hc36d058a, 32'hc0abf0ca},
  {32'hc505926f, 32'h438c155d, 32'h43543575},
  {32'h450804b0, 32'h43ce3590, 32'hc3665128},
  {32'hc40e432e, 32'hc36a3ffe, 32'hc281f8df},
  {32'h44313fc7, 32'h44013af8, 32'hc35092a8},
  {32'hc4d1859d, 32'h42de6c67, 32'h4305349f},
  {32'h44d6c581, 32'h42ce8666, 32'h438f9720},
  {32'hc30f1431, 32'h404a1760, 32'hc3285465},
  {32'h44aa066e, 32'h43120ba2, 32'h43252516},
  {32'hc3fd4d40, 32'h427e90ce, 32'h43a3d142},
  {32'h4408af9a, 32'h42863109, 32'hc36d66c3},
  {32'h4362e777, 32'hc387ea84, 32'hc2914ee2},
  {32'h448c5454, 32'h42e17634, 32'hc3ebacce},
  {32'hc4f77b72, 32'hc392b926, 32'hc31eeeb0},
  {32'h44a6b0c8, 32'hc35ebdbe, 32'hc2cb27ab},
  {32'hc4fe8c31, 32'hc3069632, 32'hc24b300f},
  {32'h44f1d49d, 32'h436a021c, 32'hc35630e0},
  {32'hc44e8aaa, 32'h42deae97, 32'h430945db},
  {32'h4482458f, 32'h420079da, 32'h430471ec},
  {32'hc43f6dca, 32'hc1e8b6e0, 32'h436889cd},
  {32'h448e5a08, 32'hc2ac8272, 32'hc304550c},
  {32'hc49ea093, 32'hc2a7f367, 32'hc1812904},
  {32'h444a9dde, 32'hc1ee2117, 32'hc359d862},
  {32'hc4eab0aa, 32'h43852a53, 32'hc2ede123},
  {32'h450a3240, 32'h424357eb, 32'hc3d8a84b},
  {32'hc41f3c98, 32'h4338bde6, 32'h43c57979},
  {32'h44ab44fd, 32'hc36f4b84, 32'h4214b24e},
  {32'hc45a5860, 32'hc2fe58da, 32'h4318ea03},
  {32'h44a2eb86, 32'h43a8f8ea, 32'hc1a64e34},
  {32'hc4ad200c, 32'hc1b8fb0a, 32'h43866e54},
  {32'h416a6300, 32'hc1c7124c, 32'hc3752d57},
  {32'hc4a322b0, 32'h4328bd17, 32'hc1478680},
  {32'h44d33066, 32'hc3c7aabc, 32'hc2fb4476},
  {32'hc468e8b1, 32'h43c86246, 32'h429dd896},
  {32'h4489cbbe, 32'hc309d839, 32'hc39f9fc4},
  {32'hc51fd8f0, 32'h42e7e65d, 32'h42c00e2c},
  {32'h44042c23, 32'h436aaaec, 32'h43bfc832},
  {32'hc369e3ec, 32'hc2ea6307, 32'hc3983d53},
  {32'h450373ce, 32'h42c99223, 32'hc363d628},
  {32'hc486b68a, 32'hc39983d0, 32'h42601458},
  {32'h443fc918, 32'h439a70ef, 32'hc090e222},
  {32'hc4a3b59c, 32'hc33430d6, 32'hc358d92c},
  {32'h44b97e6e, 32'h43b20d43, 32'hc2196dc9},
  {32'hc45945fc, 32'hc3b7dc48, 32'hc38a8c93},
  {32'h444ed985, 32'h40867b42, 32'hc3c7828f},
  {32'hc42ae04a, 32'h436398cd, 32'hc39e6541},
  {32'h42308620, 32'h4340fed2, 32'h42d30e73},
  {32'hc4e83fb0, 32'h4383b884, 32'h42683436},
  {32'h44659cb2, 32'hc09a6dbe, 32'h43676dcd},
  {32'hc446ae3c, 32'hc3183e04, 32'h424ea672},
  {32'h450dfa71, 32'h42893fc4, 32'h4360d691},
  {32'hc4ada580, 32'h4264ed64, 32'hc408c0ac},
  {32'h4428605c, 32'hc32b0668, 32'hc21bcaeb},
  {32'hc4a35d99, 32'hc2878e22, 32'hc3021c47},
  {32'h44cee7fa, 32'hc321aac2, 32'h42eb1ec4},
  {32'hc4f63518, 32'h4205ed73, 32'h422f0435},
  {32'h44f501be, 32'h41deb561, 32'hc32976bd},
  {32'hc4a9af1a, 32'hc313da07, 32'hc205162b},
  {32'h44f1e0b7, 32'h439d2fb2, 32'h409777d3},
  {32'hc4bea99f, 32'hc2d12884, 32'h43675d4a},
  {32'h44c5fdbc, 32'hc353ae45, 32'hc3065883},
  {32'hc4c3caae, 32'h42e5890d, 32'h42eafd08},
  {32'h43f7c168, 32'hc151d2a6, 32'h4284bc09},
  {32'hc4ec8340, 32'hc3c720ca, 32'hc3ff7564},
  {32'h4509feea, 32'hc21793f1, 32'hc3e8c85d},
  {32'hc4fdb586, 32'h43a64e93, 32'hc414f591},
  {32'h44337bd6, 32'hc2fa5edf, 32'hc1f134ef},
  {32'hc4864946, 32'hc3215efc, 32'h4353f88c},
  {32'hc2f31c4c, 32'hc24d1df9, 32'h43463fe8},
  {32'hc35cb73c, 32'h43d2cf2e, 32'hc39341c3},
  {32'h43eee348, 32'hc38d2e65, 32'h433fdbbe},
  {32'hc4b68ea4, 32'h430119f0, 32'h42da8590},
  {32'h43730cf8, 32'hc2e374f8, 32'hc2ec4939},
  {32'hc524ab34, 32'hc11e2ca2, 32'h435969b3},
  {32'h44ed9e78, 32'hc31b6390, 32'h436bc6cf},
  {32'hc4ef649c, 32'h430f5f1b, 32'hc28f2322},
  {32'h4522ff20, 32'h438275b0, 32'h43969adf},
  {32'hc4687b54, 32'hc3f67378, 32'h433c0055},
  {32'h442ea00a, 32'h439adfb1, 32'hc394aabc},
  {32'hc48e4e02, 32'h43288e40, 32'hc3e1ab8e},
  {32'h4187c2f0, 32'h42e47cef, 32'h42d8f0da},
  {32'hc4cbbc8c, 32'hc317da75, 32'hc3276a27},
  {32'h44c80672, 32'hc0e8b2fa, 32'hc27e6f87},
  {32'hc4937ed0, 32'hc31d7565, 32'h416dd681},
  {32'h44d8e077, 32'hc2f2c554, 32'h438ba0b3},
  {32'hc4092260, 32'hc36e2b9a, 32'h433b0bcc},
  {32'h44881aca, 32'h42ed5ebd, 32'hc222d0c3},
  {32'hc4e89f7b, 32'h4211d88d, 32'hc238bd94},
  {32'h44d8410a, 32'h43138a46, 32'hc3f4e3df},
  {32'hc4ccbec1, 32'hc2cd38c0, 32'hc325f840},
  {32'h4472dd72, 32'h439c2895, 32'h42da5356},
  {32'hc5090b17, 32'hbfc441c8, 32'hc220964d},
  {32'h44e74cb5, 32'hc364d89e, 32'hc354f417},
  {32'hc34597bc, 32'hc36c3a9c, 32'h4206c58f},
  {32'h43eb503e, 32'hc2ff4bc4, 32'hc309475d},
  {32'hc506f6c1, 32'h439fd036, 32'hc1a4f099},
  {32'h42a15af8, 32'h432a2907, 32'hc2f348eb},
  {32'hc4eec815, 32'hc24ea458, 32'hc31be658},
  {32'h4524e467, 32'hc3d1f95b, 32'h4284d3ee},
  {32'hc4ee1a45, 32'h435d1fd6, 32'h438d454c},
  {32'h44fb9168, 32'hc2962b7a, 32'h43e15b82},
  {32'hc4b8a427, 32'hc33bb72a, 32'h43cc25c3},
  {32'h452b7f8c, 32'hc391c779, 32'h43684236},
  {32'hc49142f6, 32'h424ec56c, 32'h43889f1d},
  {32'h44eb2962, 32'hc1a91aec, 32'hc11a0ef8},
  {32'hc4fc0f7a, 32'hc39e7606, 32'hc218cd49},
  {32'h43e56e9a, 32'h41617f47, 32'h429b82ac},
  {32'hc3f99230, 32'h42ea52fb, 32'h3fa296e0},
  {32'h44efc165, 32'h43e83aba, 32'h4261bc9b},
  {32'hc4de3af2, 32'h42bd4560, 32'hc3826490},
  {32'h44b0154c, 32'hc2c893f5, 32'h41da7039},
  {32'hc42f29a2, 32'hc193281c, 32'hc243ac28},
  {32'h43c74bc0, 32'hc32ffe95, 32'hc1f7cd58},
  {32'hc4983ddb, 32'hc34da396, 32'hc4055f5f},
  {32'h41f84380, 32'h42dda730, 32'hc24b1bf3},
  {32'hc42f2ffc, 32'hc39bdd0f, 32'hc2c37d5e},
  {32'h44b88b44, 32'h43888a5d, 32'hc26599ca},
  {32'hc4835703, 32'hc2ccf3af, 32'h437a0ea7},
  {32'h44c4331c, 32'h4319ba80, 32'hc3845ce9},
  {32'hc4494ba9, 32'h42564a6f, 32'h4207ef2e},
  {32'h44e18121, 32'hc2054123, 32'hc3240cfa},
  {32'hc4d9d4d8, 32'hc2dd86d4, 32'hc2f41344},
  {32'h44e3aece, 32'hc04efd63, 32'h4329d3f0},
  {32'hc3d3806c, 32'h43e713ec, 32'hc3008f54},
  {32'h44cc6118, 32'hc28cd10e, 32'h4373bc6e},
  {32'hc4c3d72c, 32'h428614d0, 32'h42eda2ab},
  {32'h44aaccd4, 32'h42a22e95, 32'h43808a96},
  {32'hc4c373b0, 32'hc304879a, 32'h43125aa5},
  {32'h445dd7f0, 32'h430f4401, 32'h435458c9},
  {32'hc376e778, 32'h431dceca, 32'hc401716b},
  {32'h4480276f, 32'h43b59c1e, 32'h43a20f78},
  {32'hc32788fd, 32'hc329eab9, 32'hc37013a8},
  {32'h44bd6320, 32'h4351d192, 32'hc385669e},
  {32'hc4628fe8, 32'h43d1edf8, 32'h42d762e3},
  {32'h44f87f31, 32'h4330656a, 32'hc407054e},
  {32'hc42050db, 32'hc277f421, 32'hc31a22bc},
  {32'h43ce157c, 32'hc373e70b, 32'h431983c3},
  {32'hc4a6e1fa, 32'h42c03632, 32'hc156179a},
  {32'h450eae94, 32'h430561f8, 32'h435ade1b},
  {32'hc4a7ea3a, 32'hc28719fe, 32'hc32dbc8d},
  {32'h44de681f, 32'h434e81e7, 32'hc36b75c0},
  {32'hc4f41930, 32'h41b428fe, 32'hc3395d97},
  {32'h44c2a1bf, 32'h42a459a8, 32'hc39dca7c},
  {32'hc4eda00a, 32'hc3cbfdd2, 32'h436a7bd6},
  {32'h44ebd3a0, 32'h432f9f10, 32'h43ae62c4},
  {32'hc374c860, 32'h419ac8a7, 32'hc2c74eb4},
  {32'h449fbb64, 32'h4389e8b2, 32'h43c1a54f},
  {32'hc50371c6, 32'h439bed53, 32'h43947712},
  {32'h44b75ce3, 32'hc28fe003, 32'h42e59d3e},
  {32'hc4a31fd9, 32'hc311514f, 32'h4308793a},
  {32'h446fe3ac, 32'hc33695b9, 32'h437d1dfe},
  {32'hc48c3127, 32'h41af7ccf, 32'hc263445e},
  {32'h44d0647a, 32'h43b546c1, 32'hc356e564},
  {32'hc3c600b0, 32'hc3ba13ff, 32'h41da52a9},
  {32'h44e382f3, 32'hc292f21e, 32'h4313a42b},
  {32'hbf30aa00, 32'hc3effc99, 32'hc00dd5e3},
  {32'h44fc1e3d, 32'h42ed20de, 32'hc225e62a},
  {32'hc4f8e89a, 32'h423aa576, 32'h428aaecd},
  {32'h4456d2b8, 32'h4388725a, 32'hc35102d6},
  {32'hc48b2cb2, 32'h439e74ba, 32'h42cd9a0c},
  {32'h4517a520, 32'hc38d8d35, 32'h435de967},
  {32'hc42b6fd7, 32'hc28fac95, 32'hc362cb76},
  {32'h4432a9be, 32'hc3155131, 32'hc1311057},
  {32'hc50c8aa7, 32'h42c9a036, 32'h424322a5},
  {32'h4499b7b7, 32'hc116e4e5, 32'hc225da5f},
  {32'hc4e2d75a, 32'hc30aa284, 32'h43806301},
  {32'h44fed594, 32'hc2d0bf0d, 32'h43448e83},
  {32'hc4b48268, 32'hc09f4546, 32'hc302e7aa},
  {32'h436a3e30, 32'h4398080e, 32'hc114297c},
  {32'h42dacf10, 32'h43e2c29f, 32'hc356722a},
  {32'h44ff1dad, 32'h4328f94c, 32'hc3ab2f16},
  {32'hc4dbc7ad, 32'hc20d5f34, 32'h432a7415},
  {32'h43107b18, 32'hc22526a3, 32'hc3c5d469},
  {32'hc4696a8a, 32'hc332aec4, 32'hc0599a54},
  {32'h445fef72, 32'h42e90d9c, 32'hc226c2c2},
  {32'hc4f5763f, 32'h427d430f, 32'hbfdf2a65},
  {32'h44c1700e, 32'hc31e9fbb, 32'hc14c70cf},
  {32'hc40698dc, 32'hc3cc55a9, 32'h41ec5032},
  {32'h43aa6fac, 32'h435a8398, 32'hc32465c3},
  {32'hc50f160d, 32'hc3b7d5ee, 32'hc399d275},
  {32'h44494b16, 32'h42098383, 32'hc3ab46cc},
  {32'hc50b7d8f, 32'h4404bd1e, 32'hc366f08b},
  {32'h45034ad4, 32'h4349e9c3, 32'hc3ce7459},
  {32'hc42434cf, 32'h43356cdd, 32'h43278594},
  {32'h44cbb415, 32'h42cded6f, 32'h4327cd7a},
  {32'hc4b9a535, 32'hc29b4af8, 32'hc37606c2},
  {32'h44c3a93d, 32'hc3ca5d8f, 32'h434f15ea},
  {32'hc49128bd, 32'h43c71dd0, 32'hc312aa52},
  {32'h445ca881, 32'h42aabed6, 32'h42ec541a},
  {32'hc39dfc50, 32'hc2060de6, 32'h43a3f0c9},
  {32'h448b73af, 32'h436bc266, 32'hc2f118c1},
  {32'hc4ed80d6, 32'hc2788c16, 32'hc2468592},
  {32'h442f0222, 32'hc22c95cd, 32'h4341bfbe},
  {32'hc49893d4, 32'hc28ae6a6, 32'h42b6cbfe},
  {32'h42dfa980, 32'h437777c3, 32'h436e798c},
  {32'hc3ada76e, 32'h423acb81, 32'h43732a72},
  {32'h440fc9ae, 32'h43c1ae65, 32'hc2a4ab66},
  {32'hc504140c, 32'hc290d916, 32'hc2f62faf},
  {32'h4517bf52, 32'h4060070f, 32'hc319cd0f},
  {32'hc49af088, 32'h4396d1b4, 32'hc28bdbdc},
  {32'h44119ee0, 32'h3eb3d080, 32'hc237b562},
  {32'hc493e941, 32'hc285a594, 32'hc316ea11},
  {32'h44cfd8d2, 32'hc36bbf73, 32'h42fe6523},
  {32'hc42e9be7, 32'hc2e93634, 32'h435b4253},
  {32'h44a49d36, 32'hc2ef864d, 32'hc25259a0},
  {32'hc48aac8d, 32'h429a1f04, 32'hc325211c},
  {32'h4471b841, 32'hc3656828, 32'hc30cfb62},
  {32'hc3790ed0, 32'hc3764175, 32'h42f9586d},
  {32'h423863b0, 32'h4403acf3, 32'hc2155e2e},
  {32'hc3bb0c85, 32'hc34da38f, 32'hc4088852},
  {32'hc2f32240, 32'hc2ee2059, 32'hc3d66753},
  {32'hc4c87008, 32'hc3624b3c, 32'hc3079f3b},
  {32'h43e597e0, 32'hc1bd7511, 32'hc3c5e4dc},
  {32'hc2dff5d6, 32'h43b9e453, 32'hc3207015},
  {32'h448d862a, 32'h43d9d231, 32'hc37ddbf1},
  {32'hc4d190ca, 32'hc2e430c1, 32'hc2c862ab},
  {32'h450afb4b, 32'h433ef5e1, 32'h42906f65},
  {32'hc4f48523, 32'hc30476e4, 32'hc38421eb},
  {32'h444aef68, 32'h433893ca, 32'h4314d3b6},
  {32'hc4f3b300, 32'h42df7731, 32'hc2c3f706},
  {32'h444c38d2, 32'h431652f8, 32'hc3b41f72},
  {32'hc31f78f0, 32'hc38d22e9, 32'h433360ba},
  {32'h4410c4ee, 32'h4315c083, 32'hc2a87d6c},
  {32'hc40b93d1, 32'h42ac00bb, 32'h433951e3},
  {32'h43964888, 32'hc1e41e4c, 32'hc36fd400},
  {32'hc4868d71, 32'hc3d59ee6, 32'hc39616fe},
  {32'h43d2482f, 32'hc3075094, 32'hc2f026b5},
  {32'h407c6800, 32'h4375666f, 32'hc31745d0},
  {32'h4431456d, 32'h43dddcb1, 32'h4250b7f8},
  {32'hc4eeedba, 32'hc2c100aa, 32'hc38b1ebc},
  {32'h44b21167, 32'h42188786, 32'hc3dff044},
  {32'hc43935a4, 32'h43a8284d, 32'h42969eb9},
  {32'h4438f46a, 32'h4209036e, 32'h43b527d1},
  {32'hc4bfbaf2, 32'h42926c90, 32'h43031c56},
  {32'h45056082, 32'h433836d4, 32'hc2a3a2c8},
  {32'hc3e2b5a2, 32'h431bbefa, 32'h42d01164},
  {32'h417bfd80, 32'hc33e576b, 32'h437edd48},
  {32'hc46cc714, 32'h42c05fe9, 32'h423ad314},
  {32'h449644c4, 32'hc30aa4bb, 32'hc33f920c},
  {32'hc3b82253, 32'h43cf35ed, 32'hc3bb2132},
  {32'h44f9fa68, 32'h4300ab6a, 32'hc2e41775},
  {32'hc4f2be07, 32'h423584d6, 32'h42ff4316},
  {32'h429dd960, 32'h40602cff, 32'h422f72c6},
  {32'hc4f9213b, 32'hc358bc39, 32'h426fdb3c},
  {32'h438798a4, 32'hc2982499, 32'h438f5195},
  {32'hc48f4b7a, 32'hc33a1e60, 32'hc1f231f5},
  {32'h44987c6d, 32'hc1a6cde7, 32'h4072efe6},
  {32'hc47b8ac4, 32'h43075da3, 32'h41edefa0},
  {32'h449c1950, 32'h428683a7, 32'hc3a6e509},
  {32'hc51908f3, 32'hc2e48729, 32'h4262f837},
  {32'h452129e1, 32'h425099a9, 32'h40d09fc1},
  {32'hc4917516, 32'hc35cb5e0, 32'hbfbd09fa},
  {32'h448f4f31, 32'h43dc8d9e, 32'h443ad4c9},
  {32'hc48c9198, 32'h438ad6dd, 32'hc244b4f5},
  {32'h44ef9663, 32'h435596d4, 32'hbf133a15},
  {32'hc35c99d8, 32'h428aebea, 32'hc2f9bd89},
  {32'h44c6ea6a, 32'h41f5a59d, 32'h437cd45e},
  {32'hc0a97c00, 32'hc3486fa4, 32'h4271a670},
  {32'h44cdc8d0, 32'hc12ad258, 32'hc2c90591},
  {32'hc415386f, 32'h438693ce, 32'h4185702d},
  {32'h44afa5b8, 32'hc2c2f5fe, 32'h42a5e293},
  {32'hc4b70a13, 32'hc3ce54be, 32'hc2d2d6ed},
  {32'h444973e0, 32'hc20b47a3, 32'h4334b7eb},
  {32'hc4c828d6, 32'hc388903c, 32'h42971558},
  {32'h44fa0ef6, 32'h43c2a3d9, 32'hc34d45bd},
  {32'hc4c76dad, 32'hc341a2f9, 32'hc376a23f},
  {32'h449c8ff5, 32'h43ba6357, 32'hc224d4f0},
  {32'hc50048dc, 32'h432fbdb7, 32'hc35c54d7},
  {32'h44c6d87a, 32'h429d6c5b, 32'h42c7a826},
  {32'hc4796362, 32'hc1ec1ad6, 32'h421d9d8a},
  {32'h44f42b42, 32'hc37ad124, 32'h43f7f772},
  {32'hc51087fe, 32'h429926a1, 32'hc35acfea},
  {32'h44fe490b, 32'h4305d0a8, 32'h42a356cf},
  {32'hc4bba90d, 32'hc39b2fa7, 32'hc27f3d13},
  {32'h44ecdc9a, 32'h42fc5ca9, 32'hc304ae5e},
  {32'hc3ec9a1a, 32'h42a92937, 32'h43332079},
  {32'h434a521e, 32'hc32bbd55, 32'h4381b448},
  {32'h42f362b4, 32'hc261132f, 32'hc1f66a02},
  {32'h44e9c54e, 32'h4302b9db, 32'hc301b3f3},
  {32'hc50b92ec, 32'hc1f660cd, 32'hc33aee51},
  {32'h44a877a2, 32'hc3ca6578, 32'h434c3576},
  {32'hc520c276, 32'hc368244d, 32'h4274107f},
  {32'h4506e95e, 32'h432a719c, 32'hc3339f57},
  {32'hc4d84cf9, 32'hc0fcd247, 32'hc2ae60c1},
  {32'h441b2be7, 32'hc1e49dae, 32'hc195e60c},
  {32'hc29341c0, 32'h424fbf1f, 32'h42954c1d},
  {32'hc2236000, 32'h43911ad8, 32'h40ca4090},
  {32'hc4a0eec3, 32'hc2dc0bac, 32'h43b4d74f},
  {32'h4513d448, 32'hc231ebec, 32'hc2f45696},
  {32'hc4d74c2b, 32'hbf4e9af6, 32'h437edfa2},
  {32'h44153df0, 32'h43334abd, 32'hc32954f7},
  {32'hc4829a88, 32'h4304b938, 32'hc3f30d3c},
  {32'h44c09734, 32'hc1b16503, 32'hc35c1d5f},
  {32'hc2f01918, 32'hc111d036, 32'hc41f30e6},
  {32'h4504e690, 32'h434a4af4, 32'h435a425e},
  {32'hc4139340, 32'h4447c6b0, 32'hc3db7701},
  {32'h450ae619, 32'hc2aad910, 32'hc330c0f0},
  {32'hc492c7e5, 32'hc39c7955, 32'h42a37584},
  {32'h44751961, 32'hc1e6f3ad, 32'hc40f700d},
  {32'hc42b4f24, 32'hc393c114, 32'h41acb0c4},
  {32'h44c95095, 32'h3f058be8, 32'hc0813440},
  {32'hc40b69a3, 32'hc364e59b, 32'hc3406646},
  {32'h43d69774, 32'hc2e09bf0, 32'hc1c08eda},
  {32'hc41b26f1, 32'hc2d0cea7, 32'hc3259383},
  {32'h43f27de6, 32'h4332c947, 32'h435af1ec},
  {32'hc4e268ff, 32'hc17488ae, 32'hc39a0616},
  {32'h449fb02c, 32'hc300d620, 32'hc2786b18},
  {32'hc4affdde, 32'h4348ba73, 32'hc32ac67c},
  {32'h43d7aafa, 32'hc3f2bfbb, 32'h427ab18f},
  {32'hc4384966, 32'h43f57df2, 32'hc24f0a89},
  {32'h44a524e6, 32'h43618f01, 32'h42e78ce9},
  {32'hc1e56380, 32'h43809cf9, 32'hc399c966},
  {32'h44fdeff9, 32'h42cf060d, 32'hc2ee1291},
  {32'hc4f41b8d, 32'hc388ac4b, 32'hc0d1142a},
  {32'h43898391, 32'hc2b0cc97, 32'h4222c39f},
  {32'hc49a0e9d, 32'h4287679e, 32'h4287eb3c},
  {32'h44afc2eb, 32'h4202a3d3, 32'h3f859594},
  {32'hc469ce9e, 32'hc2e5927b, 32'h42d2af05},
  {32'h44de8612, 32'h434a371e, 32'hc21eab91},
  {32'hc38c9345, 32'hc3905fcf, 32'hc33da848},
  {32'h446b40ee, 32'hc4036864, 32'hc18fd081},
  {32'hc48ed44a, 32'hc40b5980, 32'hc3911642},
  {32'h44866f96, 32'hc3117734, 32'hc20b917e},
  {32'hc2231878, 32'hc21aeccf, 32'h43052809},
  {32'h4512f339, 32'h42e26d36, 32'hc3018cb9},
  {32'hc39d056c, 32'h42545c84, 32'h428d3ee0},
  {32'h4507dd19, 32'h42402fa3, 32'h433dd26d},
  {32'hc4fb81f1, 32'hc3c0ef09, 32'h42ceec08},
  {32'h43e60cec, 32'hc38949d4, 32'h43287566},
  {32'hc4f17785, 32'hc3467a63, 32'hc371ca36},
  {32'h44ecc086, 32'h43831a51, 32'h433b6ad4},
  {32'hc3acd394, 32'hc364b558, 32'h40ef6ab3},
  {32'h4491633a, 32'hc37452ab, 32'h437a826a},
  {32'hc46011f4, 32'hc3834951, 32'h431651ee},
  {32'h4501455c, 32'h42df1e6e, 32'h4298ad4a},
  {32'hc44ca958, 32'hc2256322, 32'hc2f0b6cb},
  {32'h441414ca, 32'hc2d0b601, 32'h43820c91},
  {32'hc4e1cac1, 32'hc2815a74, 32'hc3803345},
  {32'hc465ee24, 32'h42e9aed0, 32'hc28e2dcd},
  {32'h4503d656, 32'hc2905b01, 32'hc389189e},
  {32'h439a5b04, 32'hc3ccb005, 32'h4389626e},
  {32'h44d44064, 32'h429f8142, 32'hc2852da0},
  {32'hc50c6166, 32'hc360701e, 32'hc34534d4},
  {32'h450ae4fc, 32'hc2a5e421, 32'hc32e35f1},
  {32'hc3ea78c0, 32'h42f158b8, 32'hc3d8bf74},
  {32'h44d6c10e, 32'hc2c323b9, 32'h43f3b8a3},
  {32'hc4e13070, 32'h4328454f, 32'hc3a7fa68},
  {32'h441499d2, 32'h43281378, 32'hc38b1cb9},
  {32'hc3c35b28, 32'h428d5c56, 32'hc3b783b5},
  {32'h44f89b18, 32'h43232f33, 32'h430bcc0c},
  {32'hc48ee16c, 32'hc39e96c1, 32'hc3d6e291},
  {32'h44c24a59, 32'hc198e060, 32'h432f6ae2},
  {32'hc4e27e0d, 32'h40b9c1d2, 32'h41f98d8c},
  {32'h45079fdb, 32'h40db8ff0, 32'hc304ccf2},
  {32'hc4c5deb7, 32'h434e9ffe, 32'h42c99512},
  {32'h45028068, 32'h4397f755, 32'h4212aedb},
  {32'hc4a9cf26, 32'h422f90c5, 32'hc368e683},
  {32'h451322fb, 32'hc18afe56, 32'h4345b31e},
  {32'hc506abb8, 32'h431b892a, 32'hc3c0a39c},
  {32'h4478b994, 32'hc261ce58, 32'h4300414a},
  {32'hc4d24bd2, 32'h4411f169, 32'hc2546064},
  {32'h44edc9af, 32'hc3175d88, 32'h41d30a95},
  {32'hc50ae2d2, 32'hc332e1d3, 32'hc2d432d7},
  {32'h44ce3650, 32'h4104c116, 32'h4320f34b},
  {32'hc4fa2b08, 32'hc38663b8, 32'h4359224f},
  {32'h44c1c75f, 32'hc33f308d, 32'hc3226e64},
  {32'hc4d9ef4a, 32'h436cfcca, 32'hc3d0ff25},
  {32'h448b146c, 32'h402d2048, 32'h43b06508},
  {32'hc4b6e10c, 32'hc207d076, 32'hc3597dc2},
  {32'h4468798f, 32'hc38faf8c, 32'h42bcf3e3},
  {32'hc3f8a840, 32'hc27fe120, 32'hc2000879},
  {32'h43746059, 32'h42ca0f52, 32'hc261097a},
  {32'hc511224d, 32'hc34b4618, 32'hc2c4a074},
  {32'hc2204c80, 32'hc20ed76c, 32'h43a22a3d},
  {32'hc4f3ea32, 32'h42e8c3aa, 32'hc179c739},
  {32'h44ac8a80, 32'h43505782, 32'hc2a6140b},
  {32'hc4ef6f71, 32'hc24a2a56, 32'hc31df17d},
  {32'h446b116e, 32'h432c0ff9, 32'hc2972b38},
  {32'hc4eecf99, 32'hc33866ba, 32'h42d5e346},
  {32'h421b7080, 32'h437b0993, 32'hc28ff843},
  {32'hc3402168, 32'h435ec320, 32'hc2bc7f08},
  {32'h44460e2a, 32'h4358ee71, 32'hc3cfb25e},
  {32'hc4238aa8, 32'hc3d3038c, 32'hc06949a6},
  {32'h44f5fe8a, 32'hc37cbdbb, 32'h4338633b},
  {32'hc3c9bd48, 32'h437ae00c, 32'hc141f56b},
  {32'h44770138, 32'h43cf2a98, 32'h43dc3b7c},
  {32'hc396c3b0, 32'h42d81061, 32'h43537f40},
  {32'h44c06c77, 32'h4382fa9f, 32'h43404a8d},
  {32'hc504b67c, 32'h42c22787, 32'hc2a2e6e3},
  {32'h44e18411, 32'hc2e419a3, 32'h42862e8e},
  {32'hc4aa62e5, 32'h42262c1f, 32'hc2e1b22a},
  {32'h441e5458, 32'h43d45da2, 32'h42b8882c},
  {32'hc3ca7642, 32'hc3866e3c, 32'h420963ef},
  {32'h4511b853, 32'hc31a7815, 32'hc38c6481},
  {32'hc3be8e90, 32'hc29c64ca, 32'hc2b8916f},
  {32'h44a17852, 32'hc35fb2de, 32'h42869da4},
  {32'hc3ee802f, 32'hc2225cd8, 32'h41c1d6c6},
  {32'h4403ae70, 32'hbfeeac40, 32'hc2524f26},
  {32'h42b5063a, 32'hc37d79e1, 32'hc3c2d08b},
  {32'h44fbe17a, 32'hc2c9e418, 32'h4287528d},
  {32'hc4f01611, 32'h4287abac, 32'hc3f84457},
  {32'h44eedc94, 32'hc361aa5d, 32'hc1ff7cb1},
  {32'h42acb33a, 32'hc2a19f29, 32'h4380e09a},
  {32'h450e7268, 32'hc18f650a, 32'hc35e1db6},
  {32'hc2dacf00, 32'h4397abc0, 32'hc37187de},
  {32'h4381a940, 32'h42f9b7e9, 32'hc3f6efef},
  {32'h43173100, 32'hc32c6e2f, 32'hc39c9bc0},
  {32'h4415ece2, 32'hc33462a1, 32'hc315e122},
  {32'hc43c2940, 32'hc3af57aa, 32'h42988ca3},
  {32'hc2c4b0b8, 32'hc2ce5882, 32'hc34d7551},
  {32'hc22bf7c0, 32'h43aae8f3, 32'h431dc40b},
  {32'hc34556e7, 32'h4306795b, 32'hc25da134},
  {32'hc382b6a9, 32'hc321cc23, 32'h4299c807},
  {32'h44746ace, 32'h42bbbf14, 32'hc295fa8b},
  {32'hc38b005c, 32'h436215e1, 32'hc1e565b6},
  {32'h41cb9c90, 32'hc32871a5, 32'hc2acb44e},
  {32'hc407b1ee, 32'hc346389f, 32'hc0fe3702},
  {32'hc35c70b6, 32'hc3d5f227, 32'h3f3c7e9c},
  {32'hc497e8b4, 32'hc3c23258, 32'hc26b6782},
  {32'h44924d97, 32'hc3df3c20, 32'h43f797ea},
  {32'hc50a90d1, 32'hc38414ac, 32'h432fd293},
  {32'h45296c72, 32'h4291247e, 32'hc1a9c4d6},
  {32'hc3a9ee00, 32'h43415e7d, 32'h43e47a94},
  {32'h443d8fba, 32'hc29987c2, 32'h42716108},
  {32'hc43cc334, 32'h42b3da98, 32'hc2bdb5c9},
  {32'h450abf10, 32'h3fcb4e5f, 32'hc30e812f},
  {32'hc4f61f3e, 32'hc10fa5de, 32'h42f4000d},
  {32'h45034d7c, 32'hc3871de3, 32'h42686a71},
  {32'hc50b464f, 32'hc38c23a1, 32'hc1ae9982},
  {32'h44c49cff, 32'h4342a908, 32'h42fbfa3a},
  {32'hc300c916, 32'h43bd4adb, 32'hc31b087a},
  {32'hc2c98a60, 32'hc338eeb9, 32'h430aaf27},
  {32'hc412e686, 32'hc38213c9, 32'h43a9d7ed},
  {32'h4402807a, 32'h42a1d898, 32'hc2125dd5},
  {32'hc4bc74c6, 32'hc21a93e2, 32'h4300c204},
  {32'h43bf6a12, 32'h415703da, 32'hc405a62c},
  {32'hc1211e84, 32'h43b381fd, 32'h4308a416},
  {32'h4352ed88, 32'h434e0008, 32'h439ecfa2},
  {32'hc3c7830f, 32'h42bb19c1, 32'hc216b05e},
  {32'h445fd5cc, 32'h4395828b, 32'hc3020270},
  {32'hc44c3a28, 32'hc3d10238, 32'h4287a700},
  {32'h44e35c72, 32'hc3bceb6a, 32'hc31c9003},
  {32'hc4be56f5, 32'hc3d8261f, 32'h42605d80},
  {32'h44e666ca, 32'hc28c86f0, 32'hc2a0d445},
  {32'hc3c07ff9, 32'hc1e1503f, 32'h4347fa8f},
  {32'h44fd1f94, 32'hc2242a06, 32'h4291c6e4},
  {32'hc4c12655, 32'hc3378890, 32'h423aa7b0},
  {32'h43a13730, 32'h4409aa02, 32'hc1ad08d9},
  {32'hc4a45105, 32'hc3d9b6c7, 32'h428ba5a0},
  {32'h43f4870b, 32'h43a3d73d, 32'hc3a13d39},
  {32'hc3482ce8, 32'hc32d32a8, 32'hc22dab21},
  {32'h44b12574, 32'hc1edbf09, 32'hc3f52dcb},
  {32'h42b968d1, 32'hc2d5feaa, 32'h43e63432},
  {32'h451c62da, 32'h429d1505, 32'hc3063a12},
  {32'hc4f70256, 32'h41e5815c, 32'hc215aefd},
  {32'h44c3be50, 32'hc35f21c1, 32'h42a58c98},
  {32'hc4730c89, 32'hc166c5f5, 32'h4398da3b},
  {32'h44bb7cf2, 32'hc289c074, 32'hc36ed6b9},
  {32'hc0a37a00, 32'h431a8c90, 32'h431b381c},
  {32'h4327f0d8, 32'h44093eb5, 32'h437d83d6},
  {32'hc3678b3e, 32'hc1a9251d, 32'h43adc7be},
  {32'h44caefce, 32'hc34257cb, 32'h440cadf4},
  {32'hc4cde14d, 32'hc35e84ea, 32'hc1c4a5c3},
  {32'h44d3f264, 32'h42ce94df, 32'hc30af8f1},
  {32'hc50a57d6, 32'hc3ddfb66, 32'hc2db5c2a},
  {32'h44a5cb65, 32'h4358da4f, 32'hc3089909},
  {32'hc314ca88, 32'hc374ffcb, 32'hc27d10bc},
  {32'h44cc7ada, 32'h4353cc38, 32'hc32d79ba},
  {32'hc4176eb2, 32'hc323eb58, 32'hc35f2f47},
  {32'h432e24c0, 32'hbfad7150, 32'hc2befdf1},
  {32'hc4022828, 32'h43a0a167, 32'hc3c0d569},
  {32'h44986ed8, 32'hc2d71469, 32'h42d6d099},
  {32'hc4e651d2, 32'h42ece7ee, 32'hc378ff67},
  {32'h44e1b2e6, 32'hc3796aaf, 32'hc3612243},
  {32'hc4ac6725, 32'h43239565, 32'hc1ad8198},
  {32'h44fc07b4, 32'h431ad24d, 32'hc30ed891},
  {32'hc42a22e8, 32'hc0bb9686, 32'hc38e9cdd},
  {32'h439813e5, 32'h41e8f434, 32'h42eecd01},
  {32'hc4d6820e, 32'h4342ffba, 32'hc2b635b8},
  {32'h433217f4, 32'hc241e2cf, 32'h42791c31},
  {32'hc42a3ade, 32'hc37afb1e, 32'h4392dc4f},
  {32'h44c243fc, 32'h41c7787a, 32'hc3608066},
  {32'hc501a967, 32'h428776f4, 32'hc3361ff9},
  {32'h446b6c45, 32'hc2a08391, 32'hc3f704f1},
  {32'hc51a4960, 32'hc3d78301, 32'h40e99e54},
  {32'h4466dcb6, 32'h442fe0a3, 32'hc398c656},
  {32'h42bcba15, 32'hc32e7c82, 32'hc365a000},
  {32'h443cb460, 32'h411c4e1a, 32'h43a110f1},
  {32'hc3379598, 32'h43754718, 32'hc2824734},
  {32'h44ed9494, 32'h43cd7b73, 32'h43361449},
  {32'h423a9180, 32'hc389c316, 32'h43b83c72},
  {32'h44b38fa9, 32'hc3765912, 32'hc2d4969c},
  {32'hc4f0af79, 32'h4147d29d, 32'hc280d635},
  {32'h433bad0a, 32'h4370729c, 32'hc2e88241},
  {32'hc33a11ea, 32'hc2a27c58, 32'h43a979f3},
  {32'h44c55c2b, 32'h43811229, 32'h4288cc46},
  {32'hc4908dca, 32'h43a0ccce, 32'h42d52839},
  {32'h44c27aaa, 32'h419b9ea3, 32'hc1d174ca},
  {32'hc3dcb1e8, 32'hc389ce89, 32'h42afa62f},
  {32'h448b4158, 32'hc2b8040f, 32'h41fd9dc0},
  {32'hc405c2ec, 32'h4388ffa9, 32'h4330b591},
  {32'h44f5074f, 32'h4308f787, 32'hc234c5d7},
  {32'hc481d836, 32'hc208fca0, 32'h431d7aee},
  {32'h444d0e91, 32'h431c2844, 32'hc10c7252},
  {32'h42a6d04c, 32'hc283dfa5, 32'h4389edcb},
  {32'h44917c49, 32'hc277642a, 32'hc2d4de00},
  {32'hc389cbb0, 32'h4216d126, 32'hc33becde},
  {32'h44b49952, 32'h42086140, 32'h4254fa38},
  {32'hc40983e2, 32'h42e632a1, 32'hc2b3ab40},
  {32'h44b5d7ed, 32'hc2480907, 32'hc34cf2ff},
  {32'hc4fc39e2, 32'h43263ba3, 32'hc3652412},
  {32'h444aec2c, 32'h419f151a, 32'hc29dbed6},
  {32'hc439093d, 32'hc2ad9aad, 32'h43112120},
  {32'h4503b226, 32'hc28be833, 32'h420030eb},
  {32'h4290c4e0, 32'h4281d46e, 32'h42c133ad},
  {32'h43d6e18f, 32'hc28a1cb5, 32'hc24c8728},
  {32'hc5049f3e, 32'h431136f9, 32'hc381e756},
  {32'h45045702, 32'hc3887ae8, 32'hc2237b18},
  {32'hc41e2d7e, 32'h4284c5b7, 32'h432e48bc},
  {32'h44f3eaf2, 32'h438566c5, 32'hc14caa17},
  {32'hc417c09e, 32'h437f0bb8, 32'hc2aee8d1},
  {32'h44850774, 32'h42efa0ad, 32'h42c6ded4},
  {32'hc4b1efd6, 32'hc3150d4e, 32'h4302e57c},
  {32'h435b1f06, 32'h42ee3509, 32'hc356693d},
  {32'hc1aec14f, 32'hc2b95aaa, 32'h42a3ab99},
  {32'h4298eaf8, 32'h4404b31a, 32'hc232ead4},
  {32'hc431685c, 32'hc311be96, 32'h424655f5},
  {32'h44d24b48, 32'h4303ae27, 32'h43307c52},
  {32'hc42a979e, 32'h41b65517, 32'hc3460ef4},
  {32'h44fb8cd3, 32'hc296e7b2, 32'hc1a40f38},
  {32'hc3058140, 32'hc33035b4, 32'h4303991d},
  {32'h44d918e1, 32'h42fdc5c6, 32'hc24c1b42},
  {32'hc48d6022, 32'h43b129bd, 32'hc39771b9},
  {32'h450625d4, 32'h42cb3c06, 32'hc3e21775},
  {32'hc510853d, 32'hc387851e, 32'hc1db6b95},
  {32'h426ce300, 32'h4383f146, 32'hc15e8898},
  {32'hc4edb67f, 32'h40d6fac8, 32'h435f35b9},
  {32'h44413c9e, 32'h42fca99e, 32'h431215ff},
  {32'hc4c39787, 32'h434e0b99, 32'h4304761f},
  {32'h4500be7f, 32'hc34177a0, 32'h42ff65c6},
  {32'hc4284a18, 32'hc3667fb2, 32'hc3964471},
  {32'h42e588b6, 32'hc356f26d, 32'h431c983f},
  {32'hc4c7739c, 32'hc39fee0f, 32'hc25612b6},
  {32'h44c10cf4, 32'hbe3c7d52, 32'hc1b2ac8e},
  {32'hc4bd78d0, 32'hc31ffdb0, 32'h431e3bb9},
  {32'h4507ca4a, 32'hc34198b2, 32'hc1f201d4},
  {32'hc5138534, 32'hc2339d14, 32'hc3845c52},
  {32'h448c5feb, 32'hc41a827f, 32'h42f03c44},
  {32'hc4e9a49c, 32'hc3cb9954, 32'h424a7092},
  {32'h44ed1707, 32'hc3b381aa, 32'hc3d30f4d},
  {32'hc49870ec, 32'h4352ec2e, 32'h42c6622d},
  {32'h44d3aa46, 32'h41ad5a12, 32'hc380258d},
  {32'hc291ce76, 32'hc30e89ac, 32'h41cc848a},
  {32'h451204ca, 32'h43b029fd, 32'hc35e3d7c},
  {32'hc50b0464, 32'hc380a1be, 32'h41941a12},
  {32'h4500408d, 32'hc2cb5020, 32'hc3920818},
  {32'hc3fb8718, 32'hc359a781, 32'hc3a3e8b2},
  {32'h45014440, 32'h43747614, 32'h4218122d},
  {32'hc4ee0397, 32'h4261c41c, 32'h436dacf8},
  {32'h4418adb8, 32'h430b0edb, 32'h4389dea0},
  {32'hc48db12e, 32'hc290d09b, 32'hc3110256},
  {32'h44f03783, 32'h43cbdebf, 32'hc317b6b7},
  {32'hc4eb7a35, 32'h4153651c, 32'h435cfa42},
  {32'hc30b8380, 32'h434e0416, 32'h43140c13},
  {32'hc35b6f80, 32'h42b28c70, 32'h434f1284},
  {32'h43312528, 32'hc31fd77e, 32'h42260fca},
  {32'h41826b1f, 32'hc299f1c5, 32'h40040281},
  {32'h44c5cbb6, 32'hc3e7cdaa, 32'hc3555b90},
  {32'hc4a6554e, 32'h434fea45, 32'h440d3036},
  {32'h44aba860, 32'hc2e95b62, 32'hc31b39ad},
  {32'hc4bf0c36, 32'hc39db143, 32'h4286bb87},
  {32'h44c83008, 32'h4406d419, 32'hc3124680},
  {32'hc4432558, 32'h42c04273, 32'hc34a24de},
  {32'h44bf7834, 32'hc1e6019e, 32'h41c4634a},
  {32'hc4d5204d, 32'h42fc88d2, 32'hc28236fa},
  {32'h43120361, 32'h44205dfd, 32'hc31185c5},
  {32'hc37a3b8f, 32'hc3301ef2, 32'h426a7e4f},
  {32'h44a02c28, 32'h428c14d7, 32'h411a8de8},
  {32'hc4fe421c, 32'hc363e207, 32'h420a9a46},
  {32'h44fe6182, 32'hc37363b8, 32'hc40e5ffc},
  {32'hc49db25f, 32'h417295ce, 32'h43f49c59},
  {32'h445e385a, 32'h43a8e9c3, 32'hc2f1e433},
  {32'hc42bcba4, 32'h42ac90eb, 32'hc3324739},
  {32'h4502a1ee, 32'hc27353e2, 32'h438cd7f2},
  {32'hc38def8f, 32'hc37ef451, 32'hc2f04a25},
  {32'h44f1e70e, 32'h41ffe4ac, 32'h4368ea10},
  {32'hc45f5b7d, 32'hc3923b97, 32'hc244a13e},
  {32'hc26b9450, 32'hc2925478, 32'hc3519ecd},
  {32'hc44e3656, 32'hc3602962, 32'hc2ac2d15},
  {32'h44fcd854, 32'h439cd39a, 32'h43f3c5ea},
  {32'hc4bcd06e, 32'hc1b5b73d, 32'h40d48d7d},
  {32'h44fc1b47, 32'hc250bbd8, 32'h42652b77},
  {32'hc4d4e17e, 32'hc04cce3f, 32'hc3209a26},
  {32'h4416ad2a, 32'h43064764, 32'h425b9d35},
  {32'hc49c54dc, 32'hc23c8ae3, 32'hc3acb9e0},
  {32'h449fa2e1, 32'hbf3eebc0, 32'h424f7b30},
  {32'hc4c2e14a, 32'h434354fa, 32'hc329d690},
  {32'h44f753e1, 32'h40529053, 32'h43fbf49a},
  {32'hc4e2bf5c, 32'h43757acb, 32'h435222dd},
  {32'h451144d8, 32'hc109f0dc, 32'h43c8ddd3},
  {32'hc4ca031f, 32'h4348d125, 32'hc21d5073},
  {32'h43f61300, 32'hc380d224, 32'h418ce5c6},
  {32'hc429f868, 32'hc37bde35, 32'hc295d714},
  {32'h45183fa9, 32'h42cd510f, 32'h42e44975},
  {32'hc4abe86a, 32'hc3a8f315, 32'hc3f1cc7c},
  {32'h442f8eec, 32'h42db6298, 32'h4396d40f},
  {32'hc4641b00, 32'h421a7c3a, 32'hc1c89dcc},
  {32'h450ba0a6, 32'h42be03e2, 32'hc2300dc8},
  {32'hc33aaa90, 32'h4340c091, 32'h4398c7c8},
  {32'h44e0ef2c, 32'h43594099, 32'hc384abc0},
  {32'hc4d62a29, 32'hc243d098, 32'h43a72fcd},
  {32'h44cc467c, 32'hc22371f3, 32'hc306f035},
  {32'hc4549f02, 32'h42116001, 32'hc2c4451e},
  {32'h44221d34, 32'hc3311b5b, 32'hc2ce6f78},
  {32'hc516a5d7, 32'hc1b5d50e, 32'h439524e4},
  {32'h451a671d, 32'hc20b6267, 32'hc3066607},
  {32'hc44a16fd, 32'hc2e3ae66, 32'hc2f1cfe8},
  {32'h4429c3f8, 32'h43016358, 32'hc3434a0e},
  {32'hc4606d16, 32'hc275212e, 32'h437115f7},
  {32'h44a5dc14, 32'hc3b12c38, 32'hc1221e9c},
  {32'hc49ef6d2, 32'h42ae31c4, 32'h4340271c},
  {32'h44843e88, 32'h439fd373, 32'hc2a3d6df},
  {32'hc48426e1, 32'h42946b23, 32'hc2dcb3a6},
  {32'h44fa72fc, 32'hc2dfc5e0, 32'h434de624},
  {32'hc4a19c79, 32'hc3c6a754, 32'h4341a2eb},
  {32'h449bf327, 32'h438437ae, 32'h42e0e0bc},
  {32'hc3b94249, 32'hc3cbf0f1, 32'hc36fecf0},
  {32'h44b8f29c, 32'hc39bf6cd, 32'hc4069268},
  {32'hc49b6845, 32'hc27b0f38, 32'h42343a26},
  {32'h44da3f63, 32'hc37c56bd, 32'h430d5034},
  {32'hc3479230, 32'h43372920, 32'h424e2155},
  {32'h444a9ca4, 32'h440c57d8, 32'h430dc885},
  {32'hc4d08bc1, 32'h433cd1f0, 32'h42025bd2},
  {32'h441d9668, 32'h4085d0a8, 32'h42edaf73},
  {32'hc4f3b820, 32'h42f67f5a, 32'h438069c4},
  {32'h4424f08a, 32'h43b7a5f4, 32'h4383aaf7},
  {32'hc4375be6, 32'hc20ce5b2, 32'hc3967656},
  {32'h44b5f8f0, 32'h438a130c, 32'h42b114bc},
  {32'hc4a55cb7, 32'hc2fcf8d9, 32'hc2b94ed2},
  {32'h44a428ea, 32'h430a1feb, 32'hc21a2acf},
  {32'hc49e049a, 32'hc2692452, 32'hc202177b},
  {32'h45009d2e, 32'h438e9337, 32'hc2c60b58},
  {32'hc42f3ffb, 32'h42bbec0a, 32'hc31a5b94},
  {32'h44666e36, 32'h4334cb05, 32'h43385742},
  {32'hc4dd29a6, 32'hc3b40e32, 32'hc3e4ecaa},
  {32'h45092fd0, 32'h43fbe4e5, 32'hc225ec7a},
  {32'hc4f0f028, 32'h427a1f07, 32'h4145a6aa},
  {32'h43ff9ee4, 32'h4336d50d, 32'h4314272d},
  {32'hc4eac4a7, 32'h433513f7, 32'h42e2f8b9},
  {32'h44ffa940, 32'hc193f20a, 32'h42b4ea0f},
  {32'hc4cb2b42, 32'h436bc407, 32'hc2043b31},
  {32'h4504ca61, 32'hc2cb21a6, 32'h43486fb7},
  {32'hc3b5142f, 32'h43b9d83d, 32'hc33872f9},
  {32'h449304e0, 32'h433d5966, 32'hc2cb8b81},
  {32'hc4b5bb4e, 32'hc23f7987, 32'hc321179e},
  {32'h45097272, 32'h42e58f7f, 32'h418aa2fb},
  {32'hc504941a, 32'hc28fe99d, 32'h42380b17},
  {32'h448801ec, 32'hc22e29ca, 32'h436683bd},
  {32'hc50b4df3, 32'h430791d5, 32'hc2e6aa11},
  {32'h44013e28, 32'hc204948c, 32'h42e17767},
  {32'hc4fc851c, 32'h43466078, 32'hc3232d76},
  {32'h42aad100, 32'h43bedccb, 32'h4321814f},
  {32'hc50590f3, 32'h42911e40, 32'h42ab6434},
  {32'h44f26a72, 32'h433c2a97, 32'h43735f3f},
  {32'hc43eb2f4, 32'hc1c78273, 32'h4384d58b},
  {32'h44ebed4d, 32'hc3902e8a, 32'hc38c521f},
  {32'hc3f935c8, 32'hc3a84d8b, 32'h4156776a},
  {32'hc19af040, 32'h41eb01c1, 32'hc3ee5d1f},
  {32'hc4e60aba, 32'hc2d5248a, 32'hc2360d2b},
  {32'h43b3f1a3, 32'hc3653a6e, 32'hc2640188},
  {32'hc49176a8, 32'hc32fe9c9, 32'hc34589ee},
  {32'h45186a14, 32'hc28294d9, 32'hc3b422e0},
  {32'hc486dc0e, 32'h42d4b444, 32'hc41acb0a},
  {32'h44863c9a, 32'hc18aa9f6, 32'hc379085f},
  {32'hc50992be, 32'h42d9515e, 32'hc28e08f6},
  {32'h446e26a5, 32'hc24eeeb4, 32'hc38c1b64},
  {32'hc48ef9bc, 32'hc39dcefe, 32'hc204d6ed},
  {32'h44eb1250, 32'h4281557e, 32'h43ad7486},
  {32'hc503112c, 32'hc38d3f4d, 32'hc3a412b9},
  {32'h448fac40, 32'h43c73c54, 32'hc2e654a2},
  {32'hc5141877, 32'h42045bdb, 32'hc2d1666d},
  {32'h44ab6ffd, 32'h42abfefc, 32'h427e22f4},
  {32'hc50625d2, 32'h4276d026, 32'hc25e8027},
  {32'h44e45ac3, 32'hc28d1453, 32'hc3812c9c},
  {32'hc4906f78, 32'hc270ee36, 32'hc3848574},
  {32'h43877058, 32'hbf88e82a, 32'h42b5c664},
  {32'hc487b336, 32'h4360edbf, 32'hc34fd12e},
  {32'h44d18333, 32'hc3dddf75, 32'hc31319c2},
  {32'hc5086886, 32'h434480e5, 32'h41855e1a},
  {32'h43cd0721, 32'hc23ccf2c, 32'h42f5f818},
  {32'hc502e565, 32'h4303f0e9, 32'hc40b25ef},
  {32'h44b15e10, 32'h42aa50b7, 32'hc217be7c},
  {32'hc49fba1b, 32'hc1393da8, 32'hc2ed2278},
  {32'hc287c970, 32'hc3d9c435, 32'h438d9cae},
  {32'hc506b963, 32'hc3975e0b, 32'h419b8e5b},
  {32'h44e122f6, 32'hc215c4a2, 32'hc3bf21a3},
  {32'hc50a9165, 32'hc33d66c5, 32'h42a8cb52},
  {32'h4296f2b0, 32'hc4050726, 32'hc199885d},
  {32'h43d85468, 32'hc336ccd9, 32'hc38e03e5},
  {32'h44d20c0b, 32'hc2ffd2f4, 32'h43210b9f},
  {32'hc4f3d774, 32'hc304b888, 32'hc3ae0f11},
  {32'h45139b08, 32'h4397d0dc, 32'hc21f42fe},
  {32'hc3f1a7c8, 32'h42f1df1e, 32'hc28c85b1},
  {32'h444c726f, 32'hc0908ec4, 32'h431c2bda},
  {32'hc50f3190, 32'hc32bd8b2, 32'h4330d26f},
  {32'h44f1f6aa, 32'hc31faa2b, 32'hc20b2028},
  {32'hc51a21e2, 32'h41a95b36, 32'hc22355b6},
  {32'h43b7bdff, 32'h427fdb35, 32'hc2940883},
  {32'hc4e26884, 32'h42c29c88, 32'h43d2d2a7},
  {32'h432629a2, 32'h42a2d437, 32'h437fbde5},
  {32'hc4835b3e, 32'h432781dd, 32'hc3db77f9},
  {32'h43b2201c, 32'hc3aacef2, 32'hc3a35b62},
  {32'hc476b740, 32'h432c46ca, 32'h42df7166},
  {32'h44dc9cdf, 32'h438f7c5e, 32'hc18ac3fa},
  {32'hc452eb0e, 32'hc2d96e73, 32'h43844f17},
  {32'h44c0041b, 32'h434bcaf3, 32'h425df182},
  {32'hc46789a2, 32'hc287a7ff, 32'h42db1078},
  {32'h44812c5d, 32'hc3b85dc7, 32'hc3b55035},
  {32'hc4bef81a, 32'h3e734c00, 32'h429f70fe},
  {32'h44c178ef, 32'h4362dd77, 32'hc3550dc4},
  {32'hc4f0f49e, 32'hc304b37f, 32'hc3e3bea4},
  {32'h43c00b10, 32'h43b434af, 32'h42e010f0},
  {32'hc5006860, 32'h423374ff, 32'h41356c4a},
  {32'h44b6931a, 32'h428d50f0, 32'h41d7d7cb},
  {32'hc2bd4dd8, 32'hc2f9b327, 32'h4327e111},
  {32'h43b53fac, 32'hc3aa345d, 32'h42eda87d},
  {32'hc3a8c341, 32'hc3822a1a, 32'h42c459f3},
  {32'h4488108e, 32'h4307c596, 32'hc3606f2b},
  {32'hc41141c2, 32'hc0d17682, 32'h43d5dfec},
  {32'h44eda6d0, 32'h435bc108, 32'hc3bc089c},
  {32'hc51ce174, 32'hc3a7ec2e, 32'h43f2a0b4},
  {32'h44971e1e, 32'hc38a8c16, 32'hc26ea71a},
  {32'hc4846b14, 32'hc38c76c4, 32'h43939e98},
  {32'h450d0aee, 32'hc3a33d74, 32'h429e3203},
  {32'hc4e9c584, 32'h436f6658, 32'hc3d37cbe},
  {32'hc35c4988, 32'h42c77f59, 32'h4305b66c},
  {32'hc44833ca, 32'hc308a937, 32'h42804e2e},
  {32'h44a724e5, 32'h43be9454, 32'hc2d29efe},
  {32'h424e64db, 32'hc2dfe4a6, 32'h423764f9},
  {32'h440f1af3, 32'h432f195e, 32'hc3305ff5},
  {32'hc3a16c78, 32'h401c63d8, 32'h41608782},
  {32'h44b57ba8, 32'h433abd87, 32'hc3c05142},
  {32'hc512989c, 32'hc299a016, 32'h43618aca},
  {32'h4412b238, 32'h4398cfad, 32'h4383c0ed},
  {32'hc517085a, 32'h43a1e28a, 32'h4264a509},
  {32'h450dff76, 32'hc2dffbe3, 32'h434090ae},
  {32'hc3506540, 32'hc245a884, 32'hc23c6121},
  {32'h43cd33a2, 32'hc28fbefe, 32'h42d6cf01},
  {32'hc4c8a939, 32'hc193fe23, 32'hc2a7e6da},
  {32'h447903e4, 32'h43076dd2, 32'hc30017b5},
  {32'hc4a7a131, 32'hc31daba3, 32'hc3c47ec6},
  {32'h445f95fd, 32'hc25f339d, 32'h4307a0da},
  {32'hc4eeedd9, 32'hc2d3c4e8, 32'h42b39da7},
  {32'h43e1fcfc, 32'hc32a1f86, 32'hc337256b},
  {32'hc5144596, 32'h43c85abf, 32'h43c1bc90},
  {32'h44bf1817, 32'h425044fc, 32'hc33b2d81},
  {32'hc4db0eae, 32'hc2eb2dd7, 32'h43d10d3d},
  {32'h44d0bb97, 32'h4362b263, 32'h41a17a58},
  {32'hc3a3e0db, 32'h43ec5a61, 32'hc2f9f77a},
  {32'h449fd350, 32'h401078d2, 32'h436853a7},
  {32'hc44b9dd1, 32'h4182f4c8, 32'h427a15f3},
  {32'h4414ae56, 32'h4273cefc, 32'hc3178fb5},
  {32'hc435de30, 32'hc2097c31, 32'h43f37ff1},
  {32'h43562dd7, 32'h42fac1f4, 32'hc391538c},
  {32'hc388b1eb, 32'h41a5fbfa, 32'h40f7a34f},
  {32'h42ed4e20, 32'hc2e9910d, 32'hc351143b},
  {32'hc4adbda1, 32'hc344c470, 32'h43516ab7},
  {32'h44efefa3, 32'h42849ccf, 32'hc0507481},
  {32'hc42e7404, 32'hc35c2661, 32'hc164359b},
  {32'h444b1663, 32'hc358bc48, 32'h4208bd65},
  {32'h44597f3c, 32'hc2eeb818, 32'hc351a834},
  {32'hc4dad492, 32'h42d4038f, 32'hc2b52542},
  {32'h44b4cc8c, 32'hc3ba1d1b, 32'h429da4c2},
  {32'h4304c120, 32'h43bd66d8, 32'h425c5fba},
  {32'h445ce3a7, 32'hc3772be0, 32'hc3b54dd3},
  {32'hc47fa7c4, 32'h4422542a, 32'hc3609ebf},
  {32'h4497ec88, 32'h4384882c, 32'hc35b3380},
  {32'hc50956e7, 32'h4298c602, 32'hc23367dc},
  {32'h44604c8a, 32'hc3959c1a, 32'h43328d6a},
  {32'hc4acd009, 32'h43cdbdea, 32'hc286516b},
  {32'h4490733b, 32'h427d667c, 32'hc3778928},
  {32'hc440a126, 32'hc39c6a46, 32'h42921ed5},
  {32'h4513bd2f, 32'h43e0e2b2, 32'h40536fea},
  {32'hc4de1e25, 32'hc23f63d4, 32'hc2c43e9e},
  {32'h451151ba, 32'h430f1a4f, 32'h432932a8},
  {32'hc49f67e4, 32'hc37fda0a, 32'h432db42a},
  {32'h44b05afc, 32'h437d0421, 32'h42b03ae6},
  {32'h42d3e893, 32'h4309be05, 32'h42c6db1e},
  {32'h44a41839, 32'h43c27a0d, 32'hc32b8344},
  {32'hc4ca8426, 32'h437ac9fd, 32'hc352ff1c},
  {32'h43077b64, 32'hc12fe2c1, 32'hc1aec22e},
  {32'hc4f521da, 32'hc2612186, 32'hc2b22619},
  {32'h44ad9929, 32'h43a95af7, 32'hc3427279},
  {32'h41a837f0, 32'h43a6827a, 32'hc3124675},
  {32'h44b05aae, 32'hc3c57a8e, 32'h43055e47},
  {32'hc4f2a1c7, 32'h436aeb0e, 32'h43901060},
  {32'h44aa35f4, 32'h42990132, 32'hc2bc8fa4},
  {32'hc488915e, 32'h43b06b00, 32'hc26ae573},
  {32'h44a5a830, 32'h43b4a511, 32'hc01fa230},
  {32'hc4e30084, 32'h437248f2, 32'hbf990ef2},
  {32'h43cb99a0, 32'hc2544ccf, 32'h4236edf8},
  {32'hc429b149, 32'h4397dafe, 32'h42f0614e},
  {32'h44973e08, 32'h436163d8, 32'h433fecb5},
  {32'hc4e18d98, 32'hc362be52, 32'h43cb0e4b},
  {32'h442d669e, 32'hc3b046f3, 32'h42f1563d},
  {32'hc3c0f157, 32'hc342efd6, 32'hc2dabc76},
  {32'h448e448c, 32'hc32d8406, 32'hc20b994c},
  {32'hc4ae5ffc, 32'h42690d0d, 32'hc38fa05c},
  {32'h451ce3b5, 32'h43158d3b, 32'hc38998a6},
  {32'hc4999463, 32'h4270569a, 32'h4291edb4},
  {32'h44fa0968, 32'h40b8b868, 32'h4310cedb},
  {32'hc4958bf8, 32'hc35df086, 32'h43727e3f},
  {32'h451ccf0c, 32'hc3a49aaa, 32'h43381f56},
  {32'hc43e0bac, 32'hc29572b6, 32'h42a9497a},
  {32'h44db8f5e, 32'h420e04cc, 32'hc26e0a28},
  {32'hc47ad489, 32'h423a7323, 32'h42c01a2b},
  {32'h44a39960, 32'hc344fc81, 32'h43493134},
  {32'hc49ba496, 32'h43988472, 32'h43efa34c},
  {32'h4500d054, 32'h43a1f797, 32'h432ff538},
  {32'hc468e6ea, 32'hc01a435c, 32'h42f5612a},
  {32'h44c267e4, 32'h431048f8, 32'h423328da},
  {32'hc50b6090, 32'h4287006e, 32'h41798613},
  {32'h44e1869c, 32'hc282f02c, 32'h42722273},
  {32'hc513a2e8, 32'hc327ced3, 32'h431bc9d6},
  {32'h44adf131, 32'h43a494c0, 32'hc3d992df},
  {32'hc3916850, 32'h42d83d66, 32'hc43711a4},
  {32'h44d8681d, 32'h40d809bc, 32'h43beb107},
  {32'hc5022b60, 32'hc249cbc3, 32'h4354fe38},
  {32'h4523946d, 32'hc37b8f68, 32'h437da90c},
  {32'h422daa04, 32'h4383d6b0, 32'h4380290d},
  {32'h44a61cba, 32'h42bdc682, 32'h42dd71f4},
  {32'hc43957fe, 32'hc055aa9a, 32'hc301d054},
  {32'h43b3b5d0, 32'h430e0e80, 32'h4216979b},
  {32'hc50db16f, 32'hc1e7e27b, 32'hc2f668d4},
  {32'h45181cc8, 32'h42982718, 32'hc284a12b},
  {32'hc4fe7d27, 32'hc2c409dd, 32'h4399b837},
  {32'h44efb37e, 32'h42f50d32, 32'hc366478f},
  {32'hc43625d5, 32'hc416a674, 32'hc3b31357},
  {32'h44bffb23, 32'h43fcce42, 32'h41319f40},
  {32'hc35ab47c, 32'h4297334a, 32'h41a64da0},
  {32'h448dcb65, 32'hc248c3b2, 32'hc280c651},
  {32'hc42e211c, 32'hc36dd11e, 32'h43b0a1b1},
  {32'h44ce4986, 32'h427898a0, 32'hc327845c},
  {32'hc4b7246c, 32'h430ce810, 32'hc35997ea},
  {32'hc33e1588, 32'hc38bb43e, 32'h42798dee},
  {32'hc434b30f, 32'h42924f48, 32'hc3cd0265},
  {32'h4403d6e2, 32'h43a57942, 32'h4362716a},
  {32'hc4938b2a, 32'hc1b8b6ae, 32'h430e0da4},
  {32'h44d7a5d7, 32'hc3818b00, 32'h433feabf},
  {32'hc43b553d, 32'hc3adaf8d, 32'hc374019e},
  {32'h44c2b239, 32'hc3a3de10, 32'hc195e6b4},
  {32'hc457aecc, 32'h4315bcc8, 32'hc34af9ba},
  {32'h438e7bcc, 32'h43a11a40, 32'hc3543154},
  {32'hc4f554d0, 32'hc2df2aed, 32'h41a06460},
  {32'h44a380bc, 32'h4260f285, 32'h437c311a},
  {32'hc50ca49c, 32'h433923a6, 32'h42418b87},
  {32'h444102c8, 32'hc1d4254b, 32'hc40a8e05},
  {32'hc47597a4, 32'hc391b760, 32'hc1da47c2},
  {32'h447d0334, 32'hc2c7af1a, 32'h436b1eb0},
  {32'hc4a4ed2d, 32'hc3c8952f, 32'hc16e3b9f},
  {32'h44a21ad2, 32'h42267298, 32'h43143bd7},
  {32'hc4dd2e46, 32'hc3590e31, 32'h43c9a20f},
  {32'h44d45c20, 32'h434140be, 32'hc1927a6d},
  {32'hc5019d19, 32'h43f540a1, 32'h41770cc2},
  {32'h44cf7233, 32'h42c2598b, 32'hc2acfb29},
  {32'hc4021664, 32'hc3b88440, 32'h43480d14},
  {32'h44dc505c, 32'hc2ff1974, 32'hc3e3bace},
  {32'hc50a24fa, 32'hc24ff244, 32'hc3cf850a},
  {32'h44822a7a, 32'hc2d94f75, 32'hc2eca576},
  {32'hc428578c, 32'h436bc747, 32'h4393b488},
  {32'h448c3771, 32'h439e1802, 32'hc1a6c568},
  {32'hc40f7c94, 32'h43a7fa68, 32'hc31bc45d},
  {32'h44a528eb, 32'hc1442526, 32'h4412c348},
  {32'hc50db21b, 32'hc31fbdad, 32'h42acd09d},
  {32'h44d521e1, 32'h43bd0ec5, 32'h42865707},
  {32'hc4faed39, 32'hc32197dd, 32'hbe4460ad},
  {32'h4351448c, 32'hc2df7229, 32'h434b883c},
  {32'hc3ad42da, 32'h42a19c3e, 32'h427f87a1},
  {32'h43aa85de, 32'hc2938501, 32'hc3066a45},
  {32'hc47e1fdc, 32'h43333c78, 32'hc084fa7c},
  {32'h43952ec9, 32'hc365e806, 32'hc38be9ca},
  {32'hc4d8b5b8, 32'hc401d5db, 32'hc3b7bcfe},
  {32'h44c9e170, 32'hc3a6a9dc, 32'h4222db15},
  {32'hc4be6ce1, 32'hc30c6062, 32'h4322832b},
  {32'h43e542f7, 32'h43a1ee22, 32'h4366e89e},
  {32'hc4187c84, 32'hc1890d95, 32'h42c6b1b2},
  {32'h450dbdea, 32'hc38083e6, 32'h4369d952},
  {32'hc4fdf290, 32'hc3841d3f, 32'h4385db68},
  {32'h449eb872, 32'h417da0c0, 32'h41f8417a},
  {32'hc474420e, 32'h438ffeb7, 32'h418a968c},
  {32'h44fc3997, 32'hc3b415f0, 32'h4232e92c},
  {32'hc4f33b55, 32'h4287c9fc, 32'h44129158},
  {32'h44f0b7cc, 32'hc3a7d41a, 32'h4263d200},
  {32'hc5013d35, 32'hc36b89df, 32'h41a415b0},
  {32'h4485e352, 32'h433ce681, 32'hc31060eb},
  {32'h43be4da8, 32'h42e7d8c2, 32'hc3a1530b},
  {32'h450b3add, 32'hc394cc52, 32'h4246da61},
  {32'hc4d84365, 32'hc2b7de8e, 32'h439f27fd},
  {32'h43d9cb44, 32'hc38f5955, 32'h4266461c},
  {32'hc3de4ecc, 32'hc2e202ab, 32'h432e7b83},
  {32'h43b621f5, 32'h42616dff, 32'h43579e0c},
  {32'hc4c1a984, 32'hc3c2c37d, 32'h433f0933},
  {32'h44aabb46, 32'h4400628e, 32'hc27209ed},
  {32'hc3cfc584, 32'hc2863fa6, 32'hc33939f0},
  {32'h44e5f0f8, 32'h42dac901, 32'hc2ce689c},
  {32'hc500999f, 32'hc2be19a2, 32'hc316a22a},
  {32'h44ec9f90, 32'h435ced50, 32'h4332db54},
  {32'hc4bbfa32, 32'hc35599b5, 32'h415ebf79},
  {32'h44c2aed8, 32'hc30d1528, 32'h428f80b2},
  {32'hc48a1556, 32'h439b95af, 32'hc36043d6},
  {32'h450e1ff7, 32'h421c857f, 32'hc2189490},
  {32'hc4380df6, 32'h42c47f93, 32'hc2cc4753},
  {32'h44c7e3ab, 32'hc3a94017, 32'hc2bf69d0},
  {32'hc392bc18, 32'hc3baa110, 32'h440a144c},
  {32'h4506146a, 32'hc3d47c37, 32'h4385fdc1},
  {32'hc4f7e494, 32'hc31cf199, 32'h43641bdf},
  {32'h43f67294, 32'hc21901de, 32'hc0d0dab0},
  {32'hc4c4043a, 32'h43105197, 32'h42308058},
  {32'h44af267e, 32'hc310a926, 32'h434ec25a},
  {32'hc51e3756, 32'hc2d7d21d, 32'hc3a63e87},
  {32'h43d301e0, 32'hc38409b1, 32'hc25226d1},
  {32'hc4398232, 32'h4315c654, 32'hc38e3efc},
  {32'h433823d4, 32'hc30831d7, 32'hc3084879},
  {32'h429d92c0, 32'hc2bac856, 32'hc2b8aada},
  {32'h44d55527, 32'h431dcced, 32'hc170385d},
  {32'hc4c8e491, 32'h438ba9c0, 32'h40a8fc70},
  {32'h4199c140, 32'h425b727a, 32'h41111bfb},
  {32'hc4f3e8a9, 32'h43965101, 32'hc1846d4c},
  {32'h447e418d, 32'hc31b9cfa, 32'h43121a1b},
  {32'hc4c64861, 32'h410f9652, 32'h42baa88e},
  {32'h44ae3bb0, 32'h432995bc, 32'h4082a820},
  {32'hc430ff5e, 32'hc33eafaf, 32'hc2547f9d},
  {32'h4418752c, 32'hc339374d, 32'hc3cf9c56},
  {32'hc4d7cd3c, 32'h4348e846, 32'h4312094e},
  {32'h448599f4, 32'h4343a3d1, 32'h42d936d0},
  {32'hc3d9b7b4, 32'hc2a97961, 32'h432732e8},
  {32'h44a1a75c, 32'h4245e494, 32'h4408b162},
  {32'hc4bff58a, 32'hc356c46b, 32'h44087326},
  {32'h432cbe50, 32'h44296135, 32'hc2a63cf2},
  {32'hc48db68a, 32'h4383fcc2, 32'h433a4bb5},
  {32'h443a4e42, 32'h431e8fdc, 32'h437ad498},
  {32'hc5010717, 32'h43ef794f, 32'h42dc1d72},
  {32'h44fe8c96, 32'hc35594e7, 32'h42bced2c},
  {32'hc4c9b544, 32'h42dfd7a3, 32'hc3450383},
  {32'h450b0791, 32'h426c894b, 32'h41d2e47c},
  {32'hc44863d2, 32'h42e59448, 32'h437c348b},
  {32'h44dcbc75, 32'h421f4943, 32'hc3058979},
  {32'hc5265bba, 32'h42eaaf5c, 32'h4272b085},
  {32'h443f97bc, 32'hc433a13a, 32'hc2d0a2bf},
  {32'hc4a37469, 32'hc2a4040e, 32'h425b3d76},
  {32'h4418624a, 32'hc3ad0606, 32'h4369e2b7},
  {32'hc4adc8b8, 32'h43cb6d4d, 32'h424b56d2},
  {32'h44a7f886, 32'hc375d1f3, 32'hc2dc9ffe},
  {32'hc4fe7903, 32'hc40a2432, 32'h435c6033},
  {32'h44c5022d, 32'hc38067ac, 32'hc27b70e9},
  {32'hc49b6b57, 32'h43cb2480, 32'hc2695085},
  {32'h44f1b053, 32'h43f074bd, 32'hc1ecb011},
  {32'hc40a0b3b, 32'h439291ac, 32'hc353441a},
  {32'h45049083, 32'hc1f19b84, 32'hc30a96d1},
  {32'h42d2ff80, 32'hc3b6134f, 32'hc2b63428},
  {32'h44d19173, 32'hc0ef5a80, 32'h42d62ea4},
  {32'hc50c0091, 32'h42bbe68d, 32'hc30f6920},
  {32'h44cf8e78, 32'hc1d27a4e, 32'h439b8606},
  {32'hc44b1c5a, 32'hc2d4a84f, 32'h40ed39d7},
  {32'h43d484e0, 32'h43a83ee5, 32'hc2e036c3},
  {32'hc4c81148, 32'hc215e30a, 32'hc1ff8eb0},
  {32'h450eeb4c, 32'hc250e168, 32'h4390ce08},
  {32'hc4b42d90, 32'hc227aed8, 32'hc177e200},
  {32'h43cf24e0, 32'h43dc1a69, 32'h4204f4f9},
  {32'hc50ff1d6, 32'h424235fc, 32'hc20089e0},
  {32'h451bc941, 32'h439ec258, 32'h42fe98df},
  {32'hc4dccb1e, 32'hc38ab395, 32'h41baf99a},
  {32'h44d2a814, 32'hc19cca7c, 32'hc310666f},
  {32'hc4c033ce, 32'h4168263b, 32'h42e2551b},
  {32'h43ae011d, 32'hc3949e57, 32'h43a255cd},
  {32'hc4ec57e1, 32'h432c47de, 32'hc3b1f991},
  {32'h44fe4f24, 32'hc3c07efd, 32'h43fc3863},
  {32'hc4e56bb4, 32'h427c713f, 32'hc3d4e4a3},
  {32'hc383d41e, 32'h42d19d13, 32'h432da37d},
  {32'hc50b0c4a, 32'hc376b86a, 32'h43444c4f},
  {32'h44275ad3, 32'h438258bf, 32'h43281cb9},
  {32'hc4ffde0b, 32'h42ff7b17, 32'h43a89583},
  {32'h42e0cf30, 32'h42e0c084, 32'hc3b74cf8},
  {32'hc4e51a32, 32'h4245f3e6, 32'h43c3f134},
  {32'h444385c0, 32'h42f34834, 32'h435a2ba2},
  {32'hc4323eee, 32'hc2cbdc98, 32'hc221a7fd},
  {32'h4380f67c, 32'hc317528b, 32'h42c6bcd2},
  {32'hc4993d6a, 32'h4357c61b, 32'hc4177141},
  {32'h43e8ce00, 32'hc3a9a00e, 32'h4311983b},
  {32'hc4b976e4, 32'hc2843fb0, 32'h42cddf42},
  {32'h44fe6dec, 32'hc2a09aec, 32'hc22ea186},
  {32'hc431cb64, 32'h43660af1, 32'h43357de6},
  {32'h450ba163, 32'h43a95f7e, 32'h40b1fe63},
  {32'h41a1cb00, 32'hc18d5450, 32'hc307f3a0},
  {32'h440c510d, 32'h40823517, 32'hc1821895},
  {32'hc2cc5060, 32'h42dde494, 32'hc32927b8},
  {32'h4488e855, 32'h43874cf7, 32'hc38bba1c},
  {32'hc4085c20, 32'hc2a85fc9, 32'hc31ae0cd},
  {32'h444913e6, 32'hc28a775b, 32'h436e087f},
  {32'hc4f89a84, 32'h42a75535, 32'h42c8b25b},
  {32'h44939430, 32'h432603cc, 32'hc406cf5d},
  {32'hc3dd5a57, 32'hc28aa766, 32'h437ef51d},
  {32'h44205742, 32'hc3112abf, 32'hc2ab56be},
  {32'hc50f3778, 32'h41ef2049, 32'h426b87dc},
  {32'h44fa45f0, 32'h42d0d588, 32'hc2f0a27b},
  {32'hc4f917bf, 32'h4299cd66, 32'hc24c49a3},
  {32'h44b4d375, 32'hc26f7b81, 32'h42aed57b},
  {32'hc3f543f2, 32'h428861b1, 32'h431dfbea},
  {32'h44cd1f04, 32'hc1497f96, 32'h428e4a1d},
  {32'hc5195240, 32'hc2a19f51, 32'hc316da04},
  {32'h44ba5006, 32'hc37e2c0c, 32'hc0bfeaca},
  {32'hc4db455f, 32'h423b5f5c, 32'hc2a6a55e},
  {32'h41dc4140, 32'hc37a1b1d, 32'hc3978d22},
  {32'hc411ccb0, 32'hc348d894, 32'hc342deef},
  {32'h44c84d7a, 32'h42d17b76, 32'h42526487},
  {32'hc40269b5, 32'h42f24618, 32'h439ae70c},
  {32'h45022b1e, 32'hc3d1a51e, 32'hc29ee152},
  {32'hc506bcaa, 32'h437052f8, 32'h42bce86b},
  {32'h4510ab44, 32'h43399b6d, 32'h43c543b1},
  {32'hc50db560, 32'hc3d86b16, 32'h438d05d5},
  {32'h44f48125, 32'h4385a2ef, 32'h4313c92f},
  {32'hc4dcb8fc, 32'h436f8b1e, 32'h42d5f899},
  {32'h44f5e500, 32'hc31c4b3b, 32'h42e3d61f},
  {32'hc2eb4d00, 32'h42c56c52, 32'h438c7346},
  {32'h4502ef02, 32'hc375e65c, 32'hc3b9505e},
  {32'hc43eeb8c, 32'h43e62a76, 32'hc331ed04},
  {32'h44c6f49f, 32'h414de62e, 32'h42df51a8},
  {32'hc3d255a8, 32'h4403f2e4, 32'h43106f25},
  {32'h44fbffcf, 32'hc23b756b, 32'hc2cb8901},
  {32'hc505643f, 32'hc3acc646, 32'h431bbfd3},
  {32'h4352d920, 32'h416cc40e, 32'h42f70f00},
  {32'hc3ca97fe, 32'h42bf5c22, 32'hc36e51e2},
  {32'h440e9426, 32'h431669e7, 32'hc30055f4},
  {32'hc48714aa, 32'hc29f9000, 32'h42c7f9a5},
  {32'h4401191f, 32'hc39bfea3, 32'h4305d6c3},
  {32'hc4b555ab, 32'h4324f02a, 32'h43b699a1},
  {32'h448c1e05, 32'hc38a33bf, 32'h42959714},
  {32'hc4be625c, 32'h424852f1, 32'h430806fa},
  {32'h44c9c44c, 32'h4309b908, 32'hc3e1a763},
  {32'hc2cdc740, 32'h42b2ce1a, 32'hc3efec3f},
  {32'h44151102, 32'h4237c0f9, 32'hc3446757},
  {32'hc4919723, 32'h439bcfe0, 32'h43ad9850},
  {32'h4514dd68, 32'hc38b71e9, 32'hc3562617},
  {32'hc4526f7f, 32'hc29b6824, 32'hc2ec30e8},
  {32'h43c01d70, 32'hc2a01ddb, 32'hc36c8829},
  {32'hc4cf0aed, 32'h43009ad6, 32'hc293bcb9},
  {32'h44c04c98, 32'hc29fb665, 32'h4350d72c},
  {32'hc4e1e58a, 32'h42890794, 32'h43be2b4e},
  {32'h447116bc, 32'hc3951d41, 32'hc32a94f9},
  {32'hc45fddd1, 32'hc3a8a58b, 32'hbfd6c5f4},
  {32'h44e18053, 32'h41e7760a, 32'h40c19b9b},
  {32'hc5092c81, 32'hc3c26b36, 32'hc306510a},
  {32'h441636b2, 32'hc32c68a0, 32'hc36621e9},
  {32'hc36d3b64, 32'hc2f6e4aa, 32'h4299c7be},
  {32'h45213bfd, 32'hc2019b13, 32'h431cd02b},
  {32'hc4843b48, 32'h436e5ba9, 32'h438fe643},
  {32'h45087f1e, 32'hc30b560a, 32'h422d325e},
  {32'hc40bc842, 32'h42d039b1, 32'h4275045a},
  {32'h44fddaf6, 32'h42b9deb2, 32'hc31fd097},
  {32'hc5068b13, 32'hc39e2327, 32'h439040c6},
  {32'h44bb6991, 32'hc3e031cf, 32'hc259d964},
  {32'hc393f01a, 32'h42900e7f, 32'h42a16c7f},
  {32'h44c4bed2, 32'h4283417f, 32'hc1cee361},
  {32'hc4de93cd, 32'h4354766c, 32'hc36b384e},
  {32'h443093f1, 32'hc3dcb535, 32'h4294c9af},
  {32'hc507666c, 32'hc3e0c0a8, 32'hc2afbb8a},
  {32'h44d03b3d, 32'h42a144c4, 32'hc34acf98},
  {32'hc4e349f9, 32'h429ea956, 32'h43a8eb45},
  {32'h44d1cd29, 32'h430a3cf5, 32'hc3c1b770},
  {32'hc436bf3f, 32'h412ed141, 32'h429a8c67},
  {32'h4426c748, 32'h40425aa0, 32'h4204eceb},
  {32'hc4a9d5f0, 32'hc3236435, 32'h4244e611},
  {32'h449e20d2, 32'hc21f3123, 32'hc33eba7d},
  {32'hc498f7b4, 32'h43862b12, 32'hc396166f},
  {32'hc2634390, 32'h43a000cd, 32'h42583463},
  {32'hc46505a8, 32'h427d631c, 32'h42b617df},
  {32'h44f30829, 32'h432c1194, 32'hc293b63d},
  {32'hc5110945, 32'h43551d31, 32'h424b92e7},
  {32'h4426e934, 32'h433d0427, 32'h4395ea9d},
  {32'hc4630116, 32'h4371232b, 32'h435eae6a},
  {32'h44a6a665, 32'h42247865, 32'hc3a87f4e},
  {32'hc4a21c71, 32'hc39a2266, 32'hc307b76f},
  {32'h45141fd5, 32'h42ab30d1, 32'h42220224},
  {32'hc3fef0b3, 32'h41d6799e, 32'h430dba15},
  {32'h4490da98, 32'hc20421ff, 32'h42b8c938},
  {32'hc50a9682, 32'hc21bef7d, 32'hc32aece9},
  {32'h449f7259, 32'hc388c652, 32'hc2ead631},
  {32'hc454744d, 32'hc35e4cf4, 32'h42218391},
  {32'h43923a80, 32'h43d9c664, 32'h432997e6},
  {32'hc4d5c16e, 32'hc2026db7, 32'hc36e6cbc},
  {32'h4506975b, 32'h434cd052, 32'h441e91af},
  {32'hc4a87aac, 32'hc318cd24, 32'hc280a5f3},
  {32'h4504fd7d, 32'h41c751fd, 32'h4348251c},
  {32'hc4ef65b6, 32'h43a9f3e1, 32'hc2a983dd},
  {32'h42ffcff0, 32'h417714e2, 32'hc2a3f08d},
  {32'hc380be4a, 32'h414c2dac, 32'h43ec9d17},
  {32'h4474ed7c, 32'hc30a8c9a, 32'hc3700f84},
  {32'hc480cb09, 32'h43601d9e, 32'h40d32c46},
  {32'h44da1302, 32'hc289c5f2, 32'h42f3d02f},
  {32'hc41d702c, 32'h42fa5b4e, 32'hc3c1db9f},
  {32'h438bc580, 32'hc266fd70, 32'hc0a34764},
  {32'hc4080190, 32'hc2ad65d4, 32'h42be248a},
  {32'h44aa4cb1, 32'hc35615e2, 32'hc34407fa},
  {32'hc1582300, 32'h43b487a1, 32'h4264177b},
  {32'h439508ea, 32'h431649fd, 32'hc23a7db9},
  {32'hc49f1e88, 32'hc23db299, 32'h434c9a29},
  {32'h440a6834, 32'h4361a56d, 32'hc36bb134},
  {32'hc34255e7, 32'h41922324, 32'h434e305d},
  {32'h4509f798, 32'hc2f884d3, 32'h427d402d},
  {32'hc4010a40, 32'h41444713, 32'hc24c97bb},
  {32'h45100a56, 32'hc2304b19, 32'h42f9096e},
  {32'hc43a6cdc, 32'h43982875, 32'hc28e42df},
  {32'h449fb04a, 32'hc36d7f9d, 32'hc33332e2},
  {32'hc4105bb7, 32'hc3063c61, 32'hc372a5de},
  {32'h446bb448, 32'hc1cc861d, 32'hc308d115},
  {32'hc510c9de, 32'h4253ed48, 32'h437a2488},
  {32'h43f76bf2, 32'h4276aafb, 32'h435a4abd},
  {32'hc43ac773, 32'h43b52d04, 32'hc1715e85},
  {32'h44e085c1, 32'h430d5f2c, 32'h4403ab26},
  {32'hc48a8fbf, 32'hc2bb8e02, 32'hc27edaaf},
  {32'h44e1703c, 32'hc28f9ee8, 32'h420b6b49},
  {32'hc3de3574, 32'hc36d5ecf, 32'h42f3caa1},
  {32'h44f804c0, 32'hc13c848c, 32'hc32ae970},
  {32'hc508f989, 32'h4250eb43, 32'h431d9b0a},
  {32'h443b153c, 32'h43ac8010, 32'h43217a87},
  {32'hc4b55312, 32'h4336c061, 32'hc32f0375},
  {32'h44cd1eb5, 32'h43bb9360, 32'hc2f1df02},
  {32'hc4a8d9a3, 32'hc42218f4, 32'h42cf0898},
  {32'h450dac65, 32'hc1bd8597, 32'h4353087f},
  {32'hc34b0140, 32'hc30adf86, 32'h42dae868},
  {32'h44802ab9, 32'hc30971dc, 32'hc3c3a418},
  {32'hc4bc4ad0, 32'h4371d76e, 32'hc2b14311},
  {32'h450f6ae9, 32'h43860ebf, 32'h43395eec},
  {32'hc307ae70, 32'h4336789e, 32'h42bb1616},
  {32'h44e3d18f, 32'hc323c450, 32'hc3011f1f},
  {32'h4324b954, 32'h43471ddd, 32'h43964f61},
  {32'h44d968ba, 32'h42fca4bc, 32'hc37cfc73},
  {32'hc4a3491e, 32'hc351ec0e, 32'h4315e931},
  {32'h44914863, 32'h42f7de90, 32'h41b39ed6},
  {32'hc50ac558, 32'h4332f72e, 32'h43e5c83c},
  {32'h43e804d4, 32'h43d512ee, 32'hc2166a3a},
  {32'hc49096a6, 32'hc2a35eb8, 32'hc31bb176},
  {32'h44890f42, 32'h438f784f, 32'hc375ab7b},
  {32'hc4ab69a4, 32'hc378e442, 32'h43d1c54a},
  {32'h42f14ea8, 32'h422699c5, 32'hc31ff0e7},
  {32'hc4c9d9a3, 32'h429fb963, 32'h4286d326},
  {32'h44f9c63b, 32'h43919b90, 32'h4225010f},
  {32'hc5014841, 32'h42ee34d5, 32'h4361f088},
  {32'h44d6e9ac, 32'hc01460c0, 32'h43970c84},
  {32'hc460f202, 32'hc2a39360, 32'h4284143d},
  {32'h4518cef0, 32'h41dffb22, 32'hc28720df},
  {32'hc478e976, 32'hc18c271d, 32'h42e76c4c},
  {32'h44835424, 32'hc202d6dc, 32'h42354272},
  {32'hc4a40e5b, 32'h43edf823, 32'h41ef23de},
  {32'h443875de, 32'hc3a066ba, 32'h42976e2c},
  {32'hc3903c9f, 32'h4321a174, 32'h438841b7},
  {32'h44d87e33, 32'h43b0c20d, 32'hc37124f9},
  {32'hc4073690, 32'hc1c06518, 32'h43c5472e},
  {32'h450590eb, 32'h43806e72, 32'h42da7701},
  {32'hc4ec4c2d, 32'h42e59a20, 32'h428b1d8b},
  {32'h448adb64, 32'h4302dfc4, 32'hc28da8ce},
  {32'hc3a224a0, 32'h41452ee9, 32'hc2c47f4a},
  {32'h44f105c7, 32'h436f8bfd, 32'h4268f1e1},
  {32'hc44c7d6a, 32'hc3c8ec90, 32'hc2cdb8a7},
  {32'h44979700, 32'hc181cebe, 32'h41a72e5e},
  {32'hc510c358, 32'h433fa5a0, 32'h42be4864},
  {32'h44cb97f2, 32'hc14f5dc0, 32'hc324dc7f},
  {32'hc3b87ee7, 32'hc2e9aa95, 32'hc205414b},
  {32'h446bd32f, 32'h420f238e, 32'h40d1f349},
  {32'hc3ddb77e, 32'h43755626, 32'hc317fefa},
  {32'h44ee5c29, 32'h426e9232, 32'h43b2a35a},
  {32'hc4abed0a, 32'h430d02d2, 32'hc294e413},
  {32'h44d058a7, 32'hc218ce6e, 32'h42db5e96},
  {32'hc4f3438e, 32'hc33597c5, 32'hc29cfcde},
  {32'h45069e5a, 32'hc213dc60, 32'h4387ad81},
  {32'hc473207a, 32'h4339358a, 32'hc29944b9},
  {32'h450dd913, 32'h4329c637, 32'hc324a219},
  {32'hc50b7ac3, 32'h430ceb25, 32'hc2fb325f},
  {32'h438ae030, 32'hc23346ca, 32'hc372e41e},
  {32'hc4a3fdc4, 32'h425fe8ea, 32'hc2a0a780},
  {32'h435fea70, 32'h430840d4, 32'h435563a7},
  {32'hc3887a08, 32'hc1ea4d07, 32'h42bfd23f},
  {32'h45027431, 32'hc37052b2, 32'h43251a63},
  {32'hc4e58224, 32'h437ba785, 32'h43f5bb6e},
  {32'h448e9a79, 32'h4295352c, 32'h43c82f42},
  {32'hc4b2260c, 32'hc3a39d0e, 32'h43b3a940},
  {32'h44f34dcb, 32'hc2e6ccf2, 32'h42c0983e},
  {32'hc41381ee, 32'h42af619c, 32'hc241cc74},
  {32'hc38e5bce, 32'hc3345453, 32'hc39cd8b7},
  {32'hc4ec7ee0, 32'h43977832, 32'h42a86f40},
  {32'h4488be72, 32'hc30c4b99, 32'h42d0c2a3},
  {32'hc33492c8, 32'h4265ff34, 32'hc1801afa},
  {32'h4427bc68, 32'h41953a74, 32'hc0d95e12},
  {32'hc40cb51c, 32'hc3a2c151, 32'hc40fea2d},
  {32'h45064de5, 32'h43873349, 32'hc312166d},
  {32'hc4014edb, 32'hc2a11feb, 32'hc2fa74e7},
  {32'h44a748c6, 32'h43183a76, 32'hc34f3366},
  {32'hc4f44640, 32'h4111a9d8, 32'hc191f993},
  {32'h44ee657c, 32'hc2569756, 32'h4363dd4f},
  {32'hc4299247, 32'hc2e9102e, 32'hc304b0f0},
  {32'h43b6712f, 32'hc3a0bb4d, 32'h4334cb29},
  {32'hc4dde116, 32'hc3963310, 32'hc24a1f9d},
  {32'hc3dc5c3f, 32'hc341628d, 32'h42f4dbc1},
  {32'h44bb91b3, 32'hc325ddc0, 32'h436d2f96},
  {32'hc511e7c6, 32'h4373dd41, 32'hc3e5a6be},
  {32'h4493d0e1, 32'h421ba527, 32'h4276a317},
  {32'h43222ca4, 32'h431de76f, 32'hc304bd78},
  {32'h44ec3630, 32'hc33342f7, 32'h42051aaf},
  {32'hc4180175, 32'hc19dc63b, 32'hc232df55},
  {32'h4500913a, 32'hc3b204bd, 32'hc2b4f3c2},
  {32'hc30e6d30, 32'hc357d62e, 32'hc2b9a8cd},
  {32'h45021336, 32'hc32a1651, 32'hc2ca798e},
  {32'hc470a4fe, 32'hc0b311a4, 32'h433bb782},
  {32'h43c12090, 32'h424ec0eb, 32'h43c92c8f},
  {32'hc4c56e61, 32'hc2b09785, 32'hc3237c7d},
  {32'h44e0d0cf, 32'h43c810b5, 32'h4396f3dd},
  {32'hc3b68340, 32'h4331e70f, 32'hc3689205},
  {32'h43604671, 32'hc379fbce, 32'hc2f60a5f},
  {32'hc4edddda, 32'h42aea6b3, 32'hc310ebf2},
  {32'h43ba4520, 32'h4283a167, 32'h41e30b66},
  {32'hc45466b0, 32'hc2d44953, 32'hc253e030},
  {32'h44c8e68d, 32'h43250cc6, 32'hc06d09eb},
  {32'hc4e9520c, 32'h42233764, 32'h428d5361},
  {32'h4282a6f0, 32'hc3442885, 32'h4256b452},
  {32'hc4cd3df4, 32'hc3b55666, 32'hc361fb9a},
  {32'h447b3af2, 32'h42579743, 32'h43955dd6},
  {32'h4236aacb, 32'h43a2ade5, 32'hc3a68acf},
  {32'h44f5b2b4, 32'hc346d23e, 32'hc1eda2d5},
  {32'hc2656a56, 32'h42ef2050, 32'h4322eb5a},
  {32'h44ebb584, 32'hc243e823, 32'hc1643311},
  {32'h430804de, 32'h43a249ce, 32'hc408d2a8},
  {32'h4334d8e0, 32'h432fbf6a, 32'hc249f411},
  {32'hc45c72c2, 32'h430f68bb, 32'hc38cdc96},
  {32'h44ab565c, 32'h42842473, 32'hc3019340},
  {32'hc4cd1b07, 32'h3e7cc8b0, 32'hc2c0ab30},
  {32'h44dd698b, 32'h410a62b8, 32'hc3043713},
  {32'hc34f40a0, 32'h440c4ea6, 32'hc205e10e},
  {32'h44e40f9c, 32'h424793ca, 32'hc289d5b0},
  {32'hc3f26106, 32'h42394574, 32'hc29e2d1d},
  {32'h44ea37bf, 32'hc20ee94a, 32'h434b28d6},
  {32'hc2f0d308, 32'h433cc3ec, 32'hc37805e4},
  {32'h450b3696, 32'h4250becd, 32'hc2253b2d},
  {32'h42162639, 32'hc3194cd6, 32'h422781ff},
  {32'h44f06cda, 32'h43f2f9f3, 32'h42becc8d},
  {32'hc4ee2e03, 32'h4103d9e8, 32'h43028626},
  {32'h44fd9693, 32'hc3e999f1, 32'h42e9443c},
  {32'hc4a985ae, 32'hc383dd85, 32'hc11338a5},
  {32'h44a4cf86, 32'hc2bacddf, 32'hc349fa4d},
  {32'hc4eb50c2, 32'h438fabd9, 32'h42bc6eda},
  {32'h44b484f2, 32'hc19936f9, 32'h4387dcfb},
  {32'hc4b052c3, 32'hc2cd51be, 32'hc27cbd16},
  {32'h4435e15b, 32'h41712704, 32'h4393f86f},
  {32'hc364e48e, 32'hc3f341fd, 32'h42fe274b},
  {32'h44596ca4, 32'hc2a09641, 32'hc39a4dba},
  {32'hc2b69320, 32'h424e5d8e, 32'hc247cc4a},
  {32'h44e7d017, 32'h421ffd2c, 32'h42c81c92},
  {32'hc4bd4d44, 32'h433de4f9, 32'h3f0049e0},
  {32'h43ce36f5, 32'h4385c8ed, 32'hc2987d86},
  {32'hc4eba2b6, 32'h42823ba0, 32'hc292350f},
  {32'h44c4986f, 32'hc2a03320, 32'hc2ce5274},
  {32'hc2a5a580, 32'h42a8cc47, 32'h42895efa},
  {32'h451aba5b, 32'h43d293c9, 32'hc2badecd},
  {32'hc4e86bf3, 32'hc2fafbac, 32'h42fbc28e},
  {32'h44fd1b8e, 32'hc3e8b7b0, 32'h439ca68f},
  {32'hc4ab3cdc, 32'hc245bffd, 32'hc3abc858},
  {32'h4421123d, 32'hc3b7b537, 32'h42cb761a},
  {32'hc4cff64a, 32'h430bb812, 32'h43ea2b10},
  {32'h4442de3f, 32'h43acb43a, 32'h4289b4b8},
  {32'h427e9df8, 32'h4241df2d, 32'h434593f1},
  {32'h4411c987, 32'hc294a0e7, 32'hc2e0427a},
  {32'hc4436b03, 32'h436c51d4, 32'h4244f272},
  {32'h449e9672, 32'hc30c878a, 32'hc2924e97},
  {32'h43947844, 32'h440b9973, 32'h42df413d},
  {32'h446d24f9, 32'h42ae841c, 32'h438199da},
  {32'hc4a4cc6a, 32'h43bb35b7, 32'hc35cfee4},
  {32'h44b3256a, 32'h42311108, 32'h4384a102},
  {32'hc3031af0, 32'hc1901fbd, 32'h4330e974},
  {32'h44c82f9b, 32'h4367991d, 32'h43b262c8},
  {32'hc4a2cb8b, 32'h43c0968b, 32'hc408736d},
  {32'h450e370b, 32'hc2b38714, 32'h432fabea},
  {32'hc38498e0, 32'hc1fe98ec, 32'h436147f6},
  {32'h450c26e8, 32'hc3d84da8, 32'h43eea36f},
  {32'hc503fa7d, 32'h426b00ae, 32'h42abcf94},
  {32'h450efefc, 32'h4264f7ad, 32'h416eed07},
  {32'hc40919b6, 32'h437474c9, 32'hc40c5e0b},
  {32'h448980c0, 32'h418fe8e4, 32'h42c92119},
  {32'hc49acdc4, 32'h42538ce8, 32'hc376c77e},
  {32'h4179fc40, 32'hc3180fb8, 32'h439cc21f},
  {32'hc459829e, 32'hc29c62a3, 32'hc1875db8},
  {32'h438d23b4, 32'h43644fe8, 32'hc35708e2},
  {32'hc46ffd2a, 32'h437abab0, 32'h42803c71},
  {32'h448968ab, 32'hc2c1efd9, 32'h422290cf},
  {32'hc4ee19fe, 32'h428d9765, 32'hc2eaac6c},
  {32'h4441f8ca, 32'h42038746, 32'hc3215722},
  {32'hc4c7ccfb, 32'hc387a37d, 32'h43a3b774},
  {32'h4512653f, 32'h43bf70b5, 32'h426625b2},
  {32'hc3415e12, 32'h43311788, 32'h43c1d5af},
  {32'h44f1d555, 32'h4209c024, 32'hc3e4c48e},
  {32'h42dd57e0, 32'h4315dea3, 32'h42b42428},
  {32'h450ab789, 32'hc362f660, 32'h42f840e4},
  {32'hc50c85f2, 32'h43fb6b5b, 32'hc234fed5},
  {32'h450d98de, 32'hc3b8a38f, 32'h424d341a},
  {32'hc21ff440, 32'hc2d5c637, 32'h437f5796},
  {32'h4421fa60, 32'h43a70d53, 32'hc3428495},
  {32'hc3315a80, 32'hc3e49d5d, 32'h43ce51f2},
  {32'h444f22bf, 32'hc1540e1b, 32'hc1c30c96},
  {32'hc4a6473b, 32'h429865f0, 32'h4349c493},
  {32'h444d4038, 32'h42dcd978, 32'h418b8d26},
  {32'hc480257a, 32'h439bae16, 32'h42bd36b8},
  {32'h44cce5d0, 32'hc3daff0e, 32'hc39c99cb},
  {32'hc39b3770, 32'hc358f817, 32'h42c5957c},
  {32'h44f11e27, 32'h41086042, 32'h3ff555e4},
  {32'hc32ffcd0, 32'h423ac4ef, 32'hc270b6a0},
  {32'h442c9f22, 32'h43d4f0d6, 32'hc38ec85b},
  {32'hc43c3009, 32'h43bd267b, 32'hc21bd1be},
  {32'h44823b32, 32'h422d53da, 32'h437c7f8f},
  {32'hc41b1ea8, 32'h43b8a11f, 32'h42acd032},
  {32'h44257e34, 32'hc104d7a7, 32'hc3a15794},
  {32'hc50490da, 32'h4305de0d, 32'h41a86c84},
  {32'hc34dd8c4, 32'hc2fc2937, 32'h42b9733f},
  {32'hc4dee09f, 32'h43824e46, 32'h42d54d89},
  {32'h44070180, 32'hc3ac751e, 32'h4350bc51},
  {32'hc4882534, 32'h42353815, 32'h435b8575},
  {32'h44f7439a, 32'hc35af4a4, 32'h433cdafa},
  {32'hc4e9b0df, 32'h43934d00, 32'h42a2263d},
  {32'h44af4962, 32'hc3147233, 32'h4335d6ae},
  {32'hc2d28ed0, 32'hc315a3b5, 32'hc2e5fcfa},
  {32'h44228c17, 32'h42fef03e, 32'h439c95af},
  {32'hc49542e0, 32'h43a4924b, 32'h435a9e8b},
  {32'h448fcee7, 32'h42fa6282, 32'h415df1d0},
  {32'hc50324b3, 32'hc34d87ea, 32'h439d7779},
  {32'hc1f1b680, 32'h4330450b, 32'hc1a7bca8},
  {32'hc4972ee9, 32'hc38cb2e4, 32'hc202d313},
  {32'h43de0cc0, 32'hc259938d, 32'hc2234ac5},
  {32'hc5079c32, 32'h438f8d0c, 32'hc20cc62a},
  {32'h44aabaa9, 32'hc28e5609, 32'h423222e8},
  {32'hc50ee92f, 32'h41e726e3, 32'hc271c1a7},
  {32'h430d6a2d, 32'hc2cdcfc7, 32'hc2f5d99e},
  {32'hc3c06d2c, 32'hc27b3d75, 32'h43e13e0c},
  {32'h44fdad8a, 32'hc33186c1, 32'hc340e412},
  {32'hc4bf94a2, 32'h42a38a79, 32'hc3320732},
  {32'h44895ae9, 32'hc2ceb69c, 32'h435d1af5},
  {32'hc3377330, 32'h43932c1d, 32'h43f59672},
  {32'h4461dd96, 32'hc3b9e520, 32'h429567b5},
  {32'hc3ef1710, 32'h411ade43, 32'h435e9229},
  {32'h450f13fe, 32'hbfbade01, 32'hc3b14d1e},
  {32'hc3d8f5b6, 32'hc1f28cb6, 32'h42bce519},
  {32'h42f80150, 32'h4286cd64, 32'hc3ef1033},
  {32'hc40ba298, 32'h43178c03, 32'h42b4d2c1},
  {32'h44300e68, 32'h43c38d9f, 32'hc302af8c},
  {32'hc49fbf3d, 32'h43854738, 32'h4384e92c},
  {32'h43003ec6, 32'h420a66f1, 32'hc36c1dd2},
  {32'hc5097e39, 32'h42584656, 32'h43298252},
  {32'h4525f511, 32'hc3441693, 32'h4254f573},
  {32'hc4a31394, 32'hc2588dc6, 32'h432df6b0},
  {32'h44cdda3a, 32'h4382ad88, 32'h42046db2},
  {32'hc43eafe6, 32'h43850a19, 32'h42d096ce},
  {32'h44fb25ec, 32'hc325e707, 32'hc3495259},
  {32'hc486d79a, 32'h43917946, 32'h42a1f6de},
  {32'h451f20b8, 32'hc416ffd5, 32'h42a90676},
  {32'hc2f6259a, 32'h42a3059c, 32'hc34ff906},
  {32'h44921e08, 32'h434591ad, 32'h4384af89},
  {32'hc502644e, 32'hc307af47, 32'h42870955},
  {32'h44f6b908, 32'hc3a67f25, 32'h43b752c5},
  {32'hc380d01c, 32'hc1ebaea8, 32'hc3bee25a},
  {32'h45029384, 32'hc2861158, 32'h4315d864},
  {32'hc5045f16, 32'hc2ffb751, 32'hc27451da},
  {32'h44bc2458, 32'h42bc99d9, 32'hc3aad85d},
  {32'hc4f6e3ca, 32'h4401084a, 32'h43d93d5b},
  {32'h44a7c3b8, 32'hc3599566, 32'hc2d6c24a},
  {32'hc4ccbe42, 32'hc2c4b968, 32'h4306091e},
  {32'h4442317f, 32'hc38e6c7b, 32'h42a28e44},
  {32'hc50dd44f, 32'hc33f73f0, 32'h4329aa84},
  {32'h44ff902e, 32'h430f403a, 32'hc1d98b5c},
  {32'hc3a0a400, 32'hc227b950, 32'hc35434aa},
  {32'h44ebd4be, 32'hc318933e, 32'h41fcbf90},
  {32'hc4e3f4db, 32'h4304b57d, 32'hc389bfbc},
  {32'h448dfe39, 32'hc2e888ed, 32'hc2b66bd5},
  {32'hc42a6ac9, 32'h4140531c, 32'hc2c5df85},
  {32'h44762a6a, 32'h423a0feb, 32'hc2cd2f4f},
  {32'hc4a6f308, 32'h43e7cd0a, 32'h42ff2fda},
  {32'h446367cc, 32'hc2bf71d4, 32'hc3976ebe},
  {32'hc417aa46, 32'h43b0e9ea, 32'h40f3d0e3},
  {32'h45157998, 32'h43885c1e, 32'hc1527c6d},
  {32'hc4b899e0, 32'h4313d507, 32'hc20ebe01},
  {32'h45033dcc, 32'h41c7cb70, 32'hc3b420f0},
  {32'hc4877915, 32'hc314b39a, 32'hc2cac751},
  {32'h44bed735, 32'h431472f6, 32'h43c6ac0a},
  {32'hc3a72bce, 32'h43836236, 32'h431aacdd},
  {32'h44f72ad0, 32'h43820331, 32'hc28c441c},
  {32'hc42edfc6, 32'h42c5dc18, 32'hc2e6cb18},
  {32'h4474fda2, 32'h436576de, 32'hc26810d7},
  {32'hc47c68ec, 32'h433b1064, 32'h433db73d},
  {32'h43845cce, 32'h4319e265, 32'hc386aeb3},
  {32'hc374b310, 32'hc33f48f8, 32'hc2770161},
  {32'h44cf64e9, 32'h42df36fc, 32'h429f030e},
  {32'hc48aab79, 32'h41d12e5e, 32'hc2a0813e},
  {32'h448a1f81, 32'h430426bd, 32'h417ea53c},
  {32'h427b5f1d, 32'h4019a27f, 32'h42e21dc0},
  {32'h44e99bd6, 32'hc330e727, 32'hc282428b},
  {32'hc4b76f86, 32'h438da5d7, 32'h43da5ef8},
  {32'h449a1952, 32'h434cdf35, 32'h42841996},
  {32'hc2b51690, 32'hc3933455, 32'h42f86895},
  {32'hc27ca670, 32'h421e76ce, 32'h432572ec},
  {32'hc4f95f23, 32'h43be493a, 32'hc3339336},
  {32'h4459b6dd, 32'hc2e56404, 32'hc2e8dfb8},
  {32'hc41e2f9e, 32'hc2808e41, 32'hc3b1c9a4},
  {32'h429643f8, 32'h431fd22b, 32'hc39e1927},
  {32'hc4b1999c, 32'hc398186e, 32'h4320a2e7},
  {32'h44fcac24, 32'hbfa726c8, 32'h4309288b},
  {32'hc36b60e1, 32'hc331c804, 32'h401f47a0},
  {32'h43f7e312, 32'h413feb26, 32'h43bf5d58},
  {32'hc484a04a, 32'h42fd96a3, 32'h41360f8f},
  {32'h440828ca, 32'hc3f38bc3, 32'hc42e611a},
  {32'hc4eac35e, 32'hc3251c8f, 32'h431d214c},
  {32'h4287b580, 32'hc34cbfa6, 32'h430bc6ff},
  {32'hc4c5c30e, 32'h43821395, 32'hc28163e2},
  {32'h44f0e280, 32'hc2d87986, 32'hc2ee25f6},
  {32'hc505e465, 32'hc2d2400d, 32'hc34ad1e4},
  {32'h44e90ab4, 32'hc3014467, 32'hc2b45fa8},
  {32'hc5020465, 32'h4337a85e, 32'h43a22292},
  {32'h44877e2f, 32'hc2c71342, 32'h427acc44},
  {32'hc4e69a0a, 32'hc2bee769, 32'h4323d1a7},
  {32'h4496a8da, 32'h438d773c, 32'hc31d359b},
  {32'hc3803910, 32'h43508f75, 32'h43255868},
  {32'h44656900, 32'hc327d428, 32'hc372353e},
  {32'hc4a5c5df, 32'hc2f30d3d, 32'h439b5bcc},
  {32'h450015a9, 32'h432ebc0c, 32'hc3f62592},
  {32'hc4f8dd3c, 32'h43913934, 32'h42e02b84},
  {32'h44e6da38, 32'h41eedc63, 32'h418cd2f0},
  {32'hc40fce4c, 32'h439f088a, 32'hc29e7a73},
  {32'h44792edd, 32'h411851ea, 32'hc30e5e4a},
  {32'hc424122c, 32'hc3744c11, 32'h421b9be1},
  {32'h448c2e4a, 32'hc396779f, 32'hc29da0af},
  {32'hc4ef8049, 32'h43956b9b, 32'h42d4a659},
  {32'h450fbb78, 32'hc40f6bd9, 32'h43917304},
  {32'hc44fda7b, 32'h439098a4, 32'hc30c146c},
  {32'h4377e9fe, 32'h41928cbc, 32'h43c836e7},
  {32'hc4345f2a, 32'hc2b212db, 32'h42e37dd0},
  {32'h42ca07f0, 32'hc3ab75b9, 32'h42a1dd4a},
  {32'hc4bedaa5, 32'hc337ac84, 32'h4386bfea},
  {32'h4493939e, 32'hc33d03d8, 32'h435bdc32},
  {32'hc4eb442c, 32'h42da3ff4, 32'hc3988ef4},
  {32'hc289a490, 32'h4073045a, 32'hc33bea81},
  {32'h434c1a0b, 32'h434488ae, 32'h43d90ea9},
  {32'h452695ee, 32'h43ccc1b8, 32'h431c8d06},
  {32'hc4ff801f, 32'h441707de, 32'h430998c2},
  {32'h447c3c94, 32'h427fcfe1, 32'h42e16b5b},
  {32'hc4101d52, 32'hc241d6d6, 32'hc3b1a362},
  {32'h45025778, 32'h423a5228, 32'hc31386fc},
  {32'hc4e683de, 32'h438e1a07, 32'h42f0a706},
  {32'h44f2be4a, 32'hc26f7874, 32'hc388fc42},
  {32'hc2f1965e, 32'h428f687f, 32'h4312bea7},
  {32'h43c46b16, 32'hc3b31ca5, 32'hc351aaaa},
  {32'hc4849694, 32'hc18294c4, 32'h43bd9c2a},
  {32'h44c456fa, 32'h42cb41f4, 32'hc35013e5},
  {32'hc4ec9f15, 32'hc0c95baa, 32'h432dff85},
  {32'h43c42958, 32'h4351497c, 32'hc1db11ec},
  {32'hc4daf741, 32'hc35c73c8, 32'hc227bf86},
  {32'h4487a8e4, 32'hc2e846fa, 32'hc390d3c4},
  {32'hc4ea1900, 32'h42723912, 32'h41e0062a},
  {32'h449f2696, 32'hc39fdd38, 32'hc37c3142},
  {32'hc4209ea0, 32'h43804149, 32'h431c6ee3},
  {32'h43cbae86, 32'hc315215a, 32'hc1a52db2},
  {32'hc51794aa, 32'h43cfff23, 32'hc3b1d14e},
  {32'h450afe52, 32'hc31698d9, 32'h43c9530d},
  {32'hc3e5b164, 32'hc35b9c08, 32'h40d02e56},
  {32'h44696253, 32'hc3a0104c, 32'h43863fbe},
  {32'hc3e0baab, 32'hc2b83417, 32'hc3ea339f},
  {32'h4510e7a7, 32'h434362ca, 32'hc2e8c093},
  {32'hc508bce7, 32'hc366d616, 32'hc2974c8f},
  {32'h433e4c26, 32'h41c1eb3c, 32'h41bf3abb},
  {32'h42550b00, 32'h421fcb4a, 32'h429ad276},
  {32'h44d28e58, 32'h42d36be1, 32'h41cf742d},
  {32'hc485e2d2, 32'h4361a698, 32'hc38ca134},
  {32'h44e8c870, 32'h431dcb7e, 32'hc306999c},
  {32'hc4cf8f4c, 32'h43a60790, 32'hc32c7711},
  {32'h440d36e1, 32'h43126b70, 32'h437c7a8e},
  {32'hc5002c33, 32'h42a49167, 32'hc311e631},
  {32'h442da14c, 32'hc3049761, 32'hc2e3f479},
  {32'hc44ce3d7, 32'h4262faa2, 32'h439db8e2},
  {32'h42f9abd4, 32'hc2f67f5a, 32'h42aa691a},
  {32'hc48ebf40, 32'h41aa8c56, 32'hc31e4806},
  {32'h443027cc, 32'hc36d8c87, 32'hc380148c},
  {32'hc3c72ef8, 32'h41e1e1a9, 32'h436e7941},
  {32'h44f82322, 32'hc3cda253, 32'hc24d70e9},
  {32'hc4839857, 32'h4363f2f1, 32'hc1c37cbd},
  {32'h444e69ed, 32'h435ed65b, 32'h432ee7b3},
  {32'hc51225aa, 32'h41c301bd, 32'h4283eaa6},
  {32'h43d88c74, 32'hc389070a, 32'h42542050},
  {32'hc41d23d4, 32'hc06d0a10, 32'hc287bc8d},
  {32'h44fd8f59, 32'h42e1b73a, 32'h44020100},
  {32'hc41e321c, 32'hc3d63d7a, 32'h431fe121},
  {32'h44802702, 32'hc2a23762, 32'h427136e5},
  {32'hc391fd88, 32'h434ae344, 32'hc1bb2706},
  {32'h43e882e8, 32'h43f1455b, 32'hc2039cfe},
  {32'hc505da7e, 32'h4187088c, 32'h4366d733},
  {32'h44920810, 32'hc3383708, 32'h41a685e6},
  {32'hc5092e81, 32'hc3033f7f, 32'hc31963d3},
  {32'h44490fe9, 32'hc33259c0, 32'h439ddcbc},
  {32'hc41d6489, 32'h433a5ef1, 32'h430dfb5e},
  {32'h4412fa8c, 32'hc2cf9e3d, 32'h42cee695},
  {32'hc43bf960, 32'hc316a9e1, 32'h4092f41c},
  {32'h44ffff9a, 32'hc32cb55b, 32'hc363c30a},
  {32'hc3fe3b94, 32'h43acc57b, 32'hc2b7c8c4},
  {32'h43d47bc8, 32'h423dba82, 32'hc3c2692d},
  {32'hc4937a42, 32'hc3fd6159, 32'h436ff082},
  {32'h45134f52, 32'hc2f9baa0, 32'h439dbcdf},
  {32'hc35177d8, 32'hc2d43a8a, 32'hc3736a9a},
  {32'h44c7ed0f, 32'hc36ede1d, 32'h43037621},
  {32'hc487e616, 32'h431a83e7, 32'hc3d2379e},
  {32'h44e44d7d, 32'hc09e496d, 32'h43e91806},
  {32'hc428a03a, 32'h4385a1f7, 32'h41c0876a},
  {32'h447f2dbe, 32'h437b6c3e, 32'h438e8e47},
  {32'hc25586c0, 32'hc31a9db4, 32'h42e3d56a},
  {32'h42319e08, 32'h42b6de8f, 32'h43cb2c11},
  {32'hc45544ee, 32'hc38b2ae6, 32'hc36b078c},
  {32'h44e2b413, 32'hc33c064f, 32'h420bca36},
  {32'hc41966a2, 32'h42c96b71, 32'hc3d5da75},
  {32'h45212665, 32'hc2e59317, 32'h43a62c62},
  {32'hc44b30f4, 32'h43ef1f74, 32'hc407ba24},
  {32'h4498b4ce, 32'hc3b48e08, 32'hc1e103d7},
  {32'hc4e345f7, 32'h43092343, 32'hc34f4266},
  {32'h44aa9b4a, 32'h42683144, 32'hc3c26d43},
  {32'hc4960459, 32'hc37af01b, 32'hc40569a0},
  {32'h4408a0a8, 32'h42ca529e, 32'h43013594},
  {32'hc338b090, 32'h43ca5bc7, 32'hc3d815bf},
  {32'h45181c38, 32'h431f9097, 32'hc289859a},
  {32'hc502a930, 32'h43342dcc, 32'hc21ce553},
  {32'h44a9b642, 32'hc34912a4, 32'hc3dac450},
  {32'hc4c28d0e, 32'h43fab9e9, 32'h43089822},
  {32'h438b10ac, 32'h43c0912b, 32'h41964267},
  {32'hc1ea2800, 32'hc29da112, 32'hc3a02365},
  {32'h4496c5e7, 32'h43ec0722, 32'h43b10064},
  {32'hc47b3634, 32'h4307a6e2, 32'hc3c54862},
  {32'h4486ed4f, 32'h41c93350, 32'h434eece8},
  {32'hc4665a3e, 32'hc1f0cab6, 32'h4343245d},
  {32'h44ecac23, 32'hc3072ea0, 32'hc1f1c2dc},
  {32'hc4b9517a, 32'hc015138e, 32'hc20c9ecd},
  {32'h44dd46bd, 32'h4305d7cd, 32'h4226156b},
  {32'hc4ecd770, 32'hc355fd7c, 32'hc2b91143},
  {32'h43ea9288, 32'h4275566d, 32'h430e9bdb},
  {32'hc40cb991, 32'h4226417a, 32'h43bc85c1},
  {32'h4394084c, 32'h42d97975, 32'hc33aa4cd},
  {32'hc46b6d12, 32'h43f8592f, 32'h432e20d4},
  {32'h450582e8, 32'hc2a6e834, 32'hc3ee84c1},
  {32'hc48a43dd, 32'hc2a6ed92, 32'hc3f0301d},
  {32'h44476b84, 32'hc2799ab1, 32'h42cd672a},
  {32'hc4b49c50, 32'hc2919bea, 32'hc181d4fa},
  {32'h44faaefe, 32'hc397d924, 32'h434b21aa},
  {32'hc49c823c, 32'hc2aae102, 32'hc3d94cf9},
  {32'h4478f8a8, 32'h4299611a, 32'hc2a8941c},
  {32'hc4c350c6, 32'hc3a37258, 32'h431ed442},
  {32'h431a27b0, 32'hc39595b1, 32'hc30d728e},
  {32'hc5120a26, 32'hc20d6657, 32'hc379f586},
  {32'h451b207c, 32'h42e2c8fb, 32'hc32cb89a},
  {32'hc413e64b, 32'h43b03e5f, 32'hc08f4104},
  {32'h44d14c28, 32'hc2fb8a07, 32'h42b19ab2},
  {32'hc40e7e6d, 32'h439cfcc7, 32'hc3179be8},
  {32'h44f679c2, 32'hc3ab9720, 32'hc3d610e4},
  {32'hc474a15c, 32'hc2361cfa, 32'h42d19c57},
  {32'h449b41cf, 32'hc25f4473, 32'hc329f9a1},
  {32'hc3e0044c, 32'h43844602, 32'h41c3db1f},
  {32'h44c51472, 32'hc26146e1, 32'h422879cb},
  {32'hc4aa772d, 32'hc3229bb8, 32'h4384e01a},
  {32'h446ffbb5, 32'hc31cd9d0, 32'h414dee9f},
  {32'hc4fc8cfa, 32'h428711ae, 32'hc40d4aa0},
  {32'h4432a037, 32'hc4093f1c, 32'hc29f81da},
  {32'hc47a194d, 32'hc38999cc, 32'h430c7a4c},
  {32'h4469e864, 32'hc370b16c, 32'hc3affb7a},
  {32'hc41b4a09, 32'h434cefe5, 32'h4343de27},
  {32'h440c12a2, 32'hc38b7370, 32'hc3fd9821},
  {32'hc5114319, 32'hc242c5cb, 32'h4326d9bc},
  {32'h451be44f, 32'h4355b78a, 32'h427b0652},
  {32'hc424eb4a, 32'h43205ccf, 32'hbff01258},
  {32'h45117bc2, 32'hc3774841, 32'h43ce7587},
  {32'hc2fb7150, 32'h42831efc, 32'h41e3e6a4},
  {32'h43dcc158, 32'h429a06c0, 32'hc3b9eea7},
  {32'hc4dd4937, 32'h43a903e3, 32'h4352c66a},
  {32'h44728240, 32'h4338093e, 32'hc29a9dae},
  {32'hc4ced5d2, 32'hc108fe19, 32'hc24b8f0d},
  {32'h43e08750, 32'h43a7d55d, 32'h431dc8f2},
  {32'hc50f2145, 32'hc26402fd, 32'hc3713ef1},
  {32'h44d959ea, 32'h40dd05e7, 32'h42446269},
  {32'hc4acf4eb, 32'hc188098b, 32'hc38597a6},
  {32'h4429c621, 32'h423dfc90, 32'hc39f83fc},
  {32'hc502c283, 32'hc38b3f49, 32'h41f5cf02},
  {32'h44151298, 32'hc35ac80d, 32'hc1874eb0},
  {32'hc4d53567, 32'hc3b23796, 32'hc3c6df23},
  {32'h440988c7, 32'hc349c41c, 32'h42640627},
  {32'hc483afb1, 32'h439ccd1d, 32'h44056897},
  {32'h45071d05, 32'hc3be6a15, 32'hc0edb3aa},
  {32'hc35e52f0, 32'hc36277dc, 32'hc3777d9b},
  {32'h4494530c, 32'hc12bc6cc, 32'hc37b8dea},
  {32'hc4eb3664, 32'hc3ba4892, 32'h4105778d},
  {32'h44a3f34c, 32'h42d3342e, 32'hc3f0174e},
  {32'hc39897aa, 32'h43312013, 32'h427c311a},
  {32'h4302e604, 32'hc3ed45a8, 32'h439ac623},
  {32'hc4066c2b, 32'hc1d2e47b, 32'h436b7836},
  {32'h43e94e60, 32'hc2b6e84a, 32'h430bc888},
  {32'hc3d73c38, 32'h4330be2e, 32'h429bd431},
  {32'h4508d7fb, 32'h4301092a, 32'hc3f0b3b3},
  {32'hc4a9beba, 32'hc2b60cf4, 32'hc336cc52},
  {32'h43eb05e2, 32'hc2844979, 32'hc43247e0},
  {32'hc45731b1, 32'h4338291d, 32'h4356fa0a},
  {32'h44bc7f32, 32'h4313cff9, 32'h4359c5ce},
  {32'hc46e04ae, 32'h437098a4, 32'h434f7e73},
  {32'h44bbb960, 32'hc1ae58e5, 32'hc2b3b3ab},
  {32'hc4a0203d, 32'hc2dabc81, 32'hc388f0a9},
  {32'h43acf708, 32'hc31c051b, 32'hc297a63f},
  {32'hc455ea11, 32'h43820f2b, 32'h4336f837},
  {32'h4441f754, 32'hc30d3e53, 32'hc345477c},
  {32'hc497553e, 32'h420fd0d3, 32'h42d61859},
  {32'h4488b3b8, 32'h434f6f7e, 32'h43971124},
  {32'hc421ad4e, 32'hc29babaa, 32'h43b4e699},
  {32'h451372ca, 32'hc346a8a6, 32'hc386764f},
  {32'hc41aa51a, 32'hc1633a2b, 32'h43247321},
  {32'h44170715, 32'hc3bebd2f, 32'hc3b14761},
  {32'hc481a35d, 32'h43883474, 32'h438e53b2},
  {32'h43ed34c4, 32'hc33d20f2, 32'hbfc4a962},
  {32'hc51e7176, 32'hc38c3378, 32'h4362ac9a},
  {32'h44b4fba8, 32'hc295c0da, 32'hc38c67d5},
  {32'hc484a5bf, 32'h42db7cb9, 32'h42c58984},
  {32'h44dea8b8, 32'hc2d654f0, 32'hc24a1c8c},
  {32'hc4378cc4, 32'hc3b7d043, 32'h43863677},
  {32'h4494d4e3, 32'h43a3b8e4, 32'hc399e170},
  {32'h42302408, 32'hc3108ea5, 32'h43ebc374},
  {32'h4428d03c, 32'h43247882, 32'hc2b6f9fe},
  {32'h428f9ec0, 32'h435bf5d1, 32'h4367945f},
  {32'h447d01b2, 32'hc2e4bcd8, 32'h438f5017},
  {32'hc4aa9271, 32'h41c1af88, 32'hc35c4976},
  {32'h426e6620, 32'hc3a91191, 32'hc2aa889f},
  {32'hc478cf8a, 32'hc1ff7304, 32'h431ffd84},
  {32'h448a0928, 32'h4315472c, 32'hc3675aa8},
  {32'h4492bf28, 32'h4356b33f, 32'hc3891eff},
  {32'hc50a2cca, 32'h4306ccda, 32'h42296869},
  {32'h45090ea5, 32'h42b1d0a9, 32'h437ca7bf},
  {32'hc4c3ac9a, 32'h4408e3bb, 32'h42873079},
  {32'h43bfb85c, 32'hc382785e, 32'h4168e720},
  {32'hc5008ff1, 32'hc3a5ee24, 32'h4256bc2e},
  {32'h4508564b, 32'h43dca17d, 32'hc2f2cfef},
  {32'h43a695ac, 32'h430eb1d3, 32'hc3c9d39a},
  {32'h43a0fc3b, 32'h42674b94, 32'hc2fa98ae},
  {32'hc502fa1e, 32'h412be476, 32'hc3adc2ca},
  {32'h4442e58c, 32'h40468dd0, 32'h42dcc0b1},
  {32'hc3e37a90, 32'h42f350bb, 32'hc31e6ac4},
  {32'h44ab3e60, 32'hc31f8208, 32'h42d35bf5},
  {32'hc46c0c54, 32'hc2cc69ca, 32'hc359546b},
  {32'h438ca450, 32'h42daa327, 32'h434a114f},
  {32'hc4b17de7, 32'hc2dbc556, 32'hc32a158d},
  {32'h44991e13, 32'hc2c11bdf, 32'hc3299c34},
  {32'hc501ec75, 32'h42ff25f1, 32'h431297ff},
  {32'h443eaa2a, 32'h4320ca5f, 32'h43a63352},
  {32'hc418a196, 32'hc2c76d27, 32'h42c03ca5},
  {32'h43e12995, 32'h43247b70, 32'hbea6edb3},
  {32'hc3c2160a, 32'hc376587d, 32'h434fb990},
  {32'h43bf931e, 32'h435bb4c9, 32'h41f7f0c3},
  {32'hc4fb2d91, 32'hc1a593a4, 32'h429b025f},
  {32'h4461023c, 32'h43090cc8, 32'hc3b519d0},
  {32'hc49011ce, 32'hc209ba96, 32'h437ddcf9},
  {32'h441768e5, 32'hc3cac758, 32'hc319bfff},
  {32'hc3f29bbf, 32'h428d10e0, 32'hc3f45a77},
  {32'h4206cc50, 32'hc296207d, 32'hc39f7359},
  {32'hc4bea18e, 32'hc2a75ad1, 32'h43df9b96},
  {32'h4382f916, 32'hc2331162, 32'hc2d9c57d},
  {32'hc4dd7ee3, 32'hc3b194a4, 32'h43b1aad1},
  {32'h4511d2a6, 32'hc1115398, 32'h44458718},
  {32'hc3c70ef7, 32'h4346e8e2, 32'h438546bd},
  {32'h44a29809, 32'h4123a74c, 32'hc35c8932},
  {32'hc4af6279, 32'hc32aad30, 32'h43e8bc02},
  {32'h44ca5758, 32'h429ad83e, 32'h435becb1},
  {32'hc4ca8c52, 32'h428cc3e5, 32'hc2a39a80},
  {32'h44ce2bc8, 32'hc2ab5bfd, 32'hc3d4f9d4},
  {32'hc4d10f30, 32'hc363ae23, 32'hc286f7be},
  {32'h44267300, 32'hc3d8b614, 32'hc022f204},
  {32'hc49ac77e, 32'hc2b7da29, 32'hc32326f6},
  {32'h43cad502, 32'hc099acca, 32'h43b9befc},
  {32'hc50e0907, 32'hc308dc3d, 32'h43475317},
  {32'h44f5a3ba, 32'h429a0b21, 32'hc2957a1b},
  {32'hc4110e7a, 32'h4306249f, 32'hc34a252b},
  {32'h450fa1c6, 32'h43ac401b, 32'h42597527},
  {32'hc4e9c2b9, 32'h425d096b, 32'h42ce310f},
  {32'h44c92932, 32'h4252c995, 32'h41acfad1},
  {32'hc3960bfe, 32'hc28a7582, 32'hc2b6630e},
  {32'h44735480, 32'hc34462a5, 32'h427f4a44},
  {32'hc4b69e41, 32'h43b96cad, 32'hc3bd76b8},
  {32'h450c34e9, 32'hc2fa4453, 32'hc2ccb28e},
  {32'hc4ad55b5, 32'hc2d8ae6e, 32'hc30f9e1b},
  {32'h44802bc2, 32'hc3912164, 32'hc2c45ead},
  {32'hc427f8ee, 32'h42105285, 32'hc3a65caa},
  {32'h450736f1, 32'hc2f7cf6f, 32'hc30b0cbe},
  {32'hc4e6b785, 32'hc2ab23bc, 32'h41d1eca3},
  {32'h4434a43e, 32'h438cdef8, 32'hc2cefee6},
  {32'hc4f0bf8a, 32'h43581ea5, 32'hc2c88568},
  {32'h43dbfb1c, 32'hc389381c, 32'hc3cc8f88},
  {32'hc405c440, 32'hc3197ce2, 32'h4320a906},
  {32'h4476fb6e, 32'hc26ed8de, 32'h42e9360a},
  {32'hc4873a6f, 32'hc2c871c0, 32'h42c9d76f},
  {32'h43aa77a0, 32'hc19a8fba, 32'h42cce432},
  {32'hc400e636, 32'h43cc494b, 32'h43bfbdd5},
  {32'h44233496, 32'h413ac4dc, 32'h3ebbe664},
  {32'hc5025aba, 32'hc3a8bd85, 32'hc3e29a21},
  {32'h44f00660, 32'hc4183952, 32'h42be43db},
  {32'hc4de7123, 32'hc2bd430d, 32'hc2a0ef42},
  {32'h4430d43e, 32'h43534798, 32'h43fb917f},
  {32'hc4de0a5c, 32'hc36a05a1, 32'hc34900df},
  {32'h44c71c9a, 32'h43e501e0, 32'hc37cc66e},
  {32'hc4fef5b9, 32'hc3af8029, 32'h433b2640},
  {32'h451eee7b, 32'h43603623, 32'h43bec17c},
  {32'hc4d4d974, 32'h4418ca95, 32'hc4228c74},
  {32'h4480210a, 32'h4389e35b, 32'h42649dba},
  {32'hc4a75243, 32'h426290ac, 32'h435238d5},
  {32'h44913fe0, 32'hc4023bd5, 32'h437d52c9},
  {32'hc4f7e437, 32'h41b1094e, 32'hc30215c7},
  {32'h43c6aa71, 32'h41ef4b1e, 32'h428bcb7f},
  {32'hc5137f9f, 32'h433e75d6, 32'hc3a95789},
  {32'h44d9a89f, 32'h442cd30c, 32'hc30daa82},
  {32'hc36ac932, 32'hc2b96c52, 32'hc381e5e4},
  {32'h44e9602f, 32'hc3b8680a, 32'hc39ce82d},
  {32'hc44aecd1, 32'hc39198ac, 32'h42b7f930},
  {32'h44cd62de, 32'hc21d704a, 32'hc3b9d7b9},
  {32'hc4d9ec84, 32'hc34c09a5, 32'h43017389},
  {32'h44cb3b41, 32'hc3a2b86d, 32'h429d6c76},
  {32'hc3d1c6a5, 32'hc2d190c7, 32'h43224de8},
  {32'h43b1e6e4, 32'hc344f442, 32'hc36dc17a},
  {32'hc4ce0494, 32'hc29553d1, 32'h42bd1e96},
  {32'h4491bb03, 32'h433c0399, 32'hc381390a},
  {32'hc50dd259, 32'h420a2fae, 32'hc2852f4c},
  {32'h443b0ff9, 32'hc3afd05f, 32'h43b5705f},
  {32'hc46c3198, 32'hc2d2fef9, 32'hc2fada8e},
  {32'h44a40b53, 32'hc2d788c2, 32'h43c21fe8},
  {32'hc4ca73df, 32'h436d90bc, 32'hc3b45b04},
  {32'h43f7a188, 32'h42a3a026, 32'hc38cc0a4},
  {32'hc41655fb, 32'h4261292a, 32'h4384d83a},
  {32'h44d9d7af, 32'h42bfd4f1, 32'hc2da33e8},
  {32'hc4a125b7, 32'hc39d3756, 32'hbf151634},
  {32'h44c50234, 32'h4318b1b6, 32'h41e06ba5},
  {32'hc4cae4d2, 32'hbfb2cb31, 32'hc1790de5},
  {32'h442adebe, 32'h40489f20, 32'hc23c836d},
  {32'hc49936fa, 32'hc2ab99ce, 32'h435258e7},
  {32'h44a289a4, 32'hc3945434, 32'hc2dbdeaa},
  {32'hc428028c, 32'h4316e5a3, 32'h42ac841b},
  {32'h44922232, 32'hc2c2cf13, 32'hc1a91d49},
  {32'hc3e635d1, 32'h41fff793, 32'hc390c892},
  {32'h44d72614, 32'hc31233bd, 32'hc20d023e},
  {32'hc4574b1c, 32'h436c81e7, 32'h42cca4bf},
  {32'h4463473f, 32'hc31da78a, 32'h43e3964b},
  {32'hc48e1b29, 32'h431b47c3, 32'hc2a9e085},
  {32'h445e48ee, 32'hc2c549f2, 32'h439f5523},
  {32'hc42ecf1c, 32'h42a061e0, 32'h3f98abec},
  {32'h44239b69, 32'hc1418b5d, 32'h42dd6d24},
  {32'hc4503b94, 32'h42e55340, 32'hc1a92eef},
  {32'h440e5ce8, 32'hc0684b9a, 32'h43a4d425},
  {32'hc3f705a8, 32'hc25ba698, 32'h435bc3da},
  {32'h43712c00, 32'hc3536135, 32'hc1e389d0},
  {32'hc41f2a38, 32'hc3b444ea, 32'hc344b095},
  {32'h450b3b1d, 32'h439fd85b, 32'h439664bc},
  {32'hc3c2faa8, 32'hc2f5e3ff, 32'h43984146},
  {32'h44ac1ed2, 32'h430f9e71, 32'hc2f0a131},
  {32'hc5015a7a, 32'h42ab35f2, 32'hc313b00c},
  {32'h44203d26, 32'hc24738b0, 32'hc25e03a3},
  {32'hc4821164, 32'h41a37e51, 32'hc344fadc},
  {32'h44aecdd4, 32'hc3209a66, 32'hc3308626},
  {32'hc42aaba8, 32'h43435898, 32'hc3542394},
  {32'h449e40fc, 32'h419bcb64, 32'h433817cb},
  {32'hc4b5a75d, 32'h4061e304, 32'hc184cf7e},
  {32'h44a41c08, 32'hc36743fa, 32'hc357de89},
  {32'hc4e6fa4a, 32'hc3ec93ad, 32'hc3025bd7},
  {32'h44fc4b76, 32'h43a20685, 32'h42a1f253},
  {32'hc499e863, 32'hc345c0b6, 32'h40865f21},
  {32'h44f1fb54, 32'hc3c834be, 32'h436632fb},
  {32'hc4ec37b6, 32'h42bbd505, 32'h433dd478},
  {32'h45115bbc, 32'hc2d8e470, 32'hc3143650},
  {32'hc41dbd28, 32'h42715a8d, 32'h4448d7b0},
  {32'h446e2111, 32'h430c855a, 32'hc34b9306},
  {32'hc4b2905a, 32'h4125ea96, 32'hc3d3b4bd},
  {32'hc2388490, 32'hc2b3378d, 32'h4359ed59},
  {32'hc4afd00c, 32'hc37d81af, 32'hc2229350},
  {32'h443bccbc, 32'hc2ceaff7, 32'hc29f54fe},
  {32'hc3fcb6e9, 32'hc2d63c82, 32'hc341d2fe},
  {32'h44d850bd, 32'h439f5d88, 32'hc324d6a3},
  {32'hc4e4b1bd, 32'hc3427814, 32'h4352b836},
  {32'h4427bf82, 32'h43625960, 32'h432fd4ee},
  {32'hc410a49b, 32'hc2c7cdc3, 32'h42493afd},
  {32'h44627c5f, 32'hc2943d58, 32'hc31e6ae3},
  {32'h41810980, 32'hc39687cb, 32'h430730d7},
  {32'h43b51d40, 32'hc1f57bb1, 32'hc383cf0e},
  {32'hc41057f0, 32'h4267d35d, 32'hc2ae7705},
  {32'h447e845e, 32'h43bce62c, 32'h425f6022},
  {32'hc42254ee, 32'hc3889f83, 32'h42b27851},
  {32'h42fc2da0, 32'hc2a31d5c, 32'h43bb7375},
  {32'hc4dfc0dd, 32'hc2322d43, 32'h43a64f00},
  {32'h44845135, 32'h428a2b3e, 32'hc3a43780},
  {32'hc4ab1bd5, 32'hc38d861e, 32'h436a20da},
  {32'h44db363f, 32'hc205791a, 32'hc381fa6b},
  {32'h42f54840, 32'h42f2a578, 32'hbd281200},
  {32'h4481236f, 32'hc2a69362, 32'hc3193353},
  {32'hc3f83d0c, 32'hc303a2ca, 32'h422d1b2e},
  {32'h44ca736c, 32'h43a4c2c3, 32'hc285b769},
  {32'hc4ed5401, 32'hc30b2ca2, 32'hc31c2886},
  {32'h44a0305f, 32'h43a21eb9, 32'h43332601},
  {32'hc4fe846e, 32'h42627eeb, 32'h43a4b923},
  {32'h439149ec, 32'h43588d26, 32'h431000c0},
  {32'hc4a26918, 32'h4277a3f8, 32'h42f554d4},
  {32'h45125926, 32'h41c9ac07, 32'h43ac80cc},
  {32'hc3a656c0, 32'h43b9fab6, 32'h439ad6b9},
  {32'h447abd64, 32'hc3058d4b, 32'hc1d60a16},
  {32'hc50c656a, 32'hc2b6b32c, 32'hc248cd55},
  {32'h4492db14, 32'hc2b22e90, 32'hc3898284},
  {32'hc4bceea2, 32'h43f8b7ef, 32'h40b5fa5c},
  {32'h4407856e, 32'h422960e1, 32'h438e64c2},
  {32'hc3db7ba4, 32'hc35b6791, 32'hc21e7a2c},
  {32'h42d00718, 32'h43148f51, 32'h4328cec6},
  {32'hc4aae763, 32'hc3f1d32a, 32'h439fba27},
  {32'h4475f4ba, 32'h434b3e30, 32'hc24e6bac},
  {32'hc2393dc8, 32'h4311971c, 32'hc0eb69ca},
  {32'h44cad277, 32'h426f4012, 32'hc319d361},
  {32'h432b34e0, 32'h4374f883, 32'hc364255e},
  {32'h44a5adbc, 32'hc39e08ed, 32'hc359f6a7},
  {32'hc4b1299c, 32'hc2e923b2, 32'hc2ff1e53},
  {32'h44b78418, 32'hc3dcf24a, 32'hc2f7e757},
  {32'hc5027892, 32'hc388138a, 32'h4397ca1e},
  {32'h44d7bfb4, 32'hc2b7c366, 32'hc362421b},
  {32'hc4b0b77e, 32'h43132631, 32'h42b18dd5},
  {32'h44c32302, 32'hc2f9ae8b, 32'h430c2198},
  {32'hc50326a7, 32'hc2c868b6, 32'h4286613b},
  {32'h44ffc8ed, 32'hc2fe4b61, 32'h432c4a34},
  {32'hc48eaf46, 32'h42d7ee5f, 32'hc34db80f},
  {32'h450c85b0, 32'h42d3287d, 32'h43806f94},
  {32'hc415ddf8, 32'hc3946167, 32'hc305c95b},
  {32'h444295fd, 32'h42bc0f81, 32'hc321029a},
  {32'hc50bf1ac, 32'hc0258218, 32'hc3065f17},
  {32'h44e9fa2d, 32'h4393b412, 32'hc1b1c60c},
  {32'hc4f730da, 32'hc36fdb00, 32'h4353f5d4},
  {32'h4406b2ed, 32'hc275d27f, 32'hc2d1594e},
  {32'hc4a27368, 32'hc39b6714, 32'hc28dcb8b},
  {32'h4504df2e, 32'h42a7cf09, 32'hc3863063},
  {32'hc52f3dda, 32'h43717817, 32'h437676d2},
  {32'h424de480, 32'hc0e7918e, 32'h431bd694},
  {32'hc3ad34e8, 32'hc1948f17, 32'h428243d9},
  {32'h449fa1b9, 32'hc3dd8834, 32'hc34948ae},
  {32'hc4950084, 32'h4353de3e, 32'hc316f387},
  {32'h444e1b4e, 32'hc31d789b, 32'h42eb8b78},
  {32'hc503cbbf, 32'h43104390, 32'h40596ac1},
  {32'h439b9663, 32'h43e480ee, 32'h43c9944f},
  {32'hc4f3ec9f, 32'hc3556727, 32'h43640542},
  {32'h447f251e, 32'hc2ae0936, 32'h43861edf},
  {32'hc4a42e46, 32'hc12ec45f, 32'h405efd93},
  {32'h4500ae91, 32'hc2aacd10, 32'hc2dd1bbf},
  {32'h4309dfad, 32'h42b66604, 32'hc3190e61},
  {32'h4409db1e, 32'hc34ce190, 32'hc332a398},
  {32'hc4f3491e, 32'hc34c776b, 32'h439ae322},
  {32'h43894594, 32'h432c1744, 32'hc35626a2},
  {32'hc4eabbff, 32'hc374a2b2, 32'hc2170244},
  {32'h4502f562, 32'h432c8e15, 32'h43960614},
  {32'hc4820ed0, 32'hc33cb4dc, 32'hc21b9b97},
  {32'h44e92924, 32'hc29900ec, 32'h42d482cc},
  {32'hc3f55c36, 32'hc2e4408e, 32'h42c2fbe5},
  {32'h4478731b, 32'h43671593, 32'hc3d670ff},
  {32'hc2aa04d0, 32'h416d5924, 32'h430b66f0},
  {32'h439fbe80, 32'hc2040c47, 32'hc35c42b1},
  {32'hc48827ba, 32'hc1e912fe, 32'h435d4e86},
  {32'h44b786f8, 32'hc2614f3d, 32'h430bff40},
  {32'hc3786bfe, 32'hc2a6d074, 32'h430e4425},
  {32'h450babf3, 32'h439b2ecc, 32'hc2ec6373},
  {32'hc4af4aaa, 32'h42e01e07, 32'hc379099e},
  {32'h44dc6852, 32'hc382e48d, 32'h42b69b5f},
  {32'hc4b75a30, 32'h42d00c80, 32'h43b59153},
  {32'h44b07152, 32'hc32ae960, 32'hc292167b},
  {32'hc4dd01d5, 32'hc24c62dc, 32'h42c433f2},
  {32'h4423a853, 32'hc3bfe9cf, 32'h4358de2b},
  {32'hc4fa76a2, 32'hc3992a60, 32'hc313e4d4},
  {32'h45161b68, 32'hc3bac7d7, 32'hc3e9b0e6},
  {32'hc51193a2, 32'h436e3cca, 32'h43d2d172},
  {32'h43ac28ee, 32'hc340d05a, 32'hc32bb1ce},
  {32'hc48da3e1, 32'h4339eb23, 32'hc3c6db36},
  {32'h44c76cc5, 32'hc210a1af, 32'h43809f6a},
  {32'hc4f690ff, 32'h436ae465, 32'hc29ee9a8},
  {32'h44f0f654, 32'hc2e59110, 32'h4303de88},
  {32'hc504a972, 32'h431870c2, 32'h436e1b9e},
  {32'h44a533a3, 32'h42d1652c, 32'hc2402c38},
  {32'hc47cc8a9, 32'hc3b9ec1a, 32'h434b472e},
  {32'h44128bf8, 32'h418704ee, 32'h42874c35},
  {32'hc39d1246, 32'hc1b4d638, 32'h40a61d19},
  {32'h45048213, 32'h41b501fa, 32'h426fa07b},
  {32'hc48f1054, 32'hc3b86fa4, 32'h42cd1e05},
  {32'hc2f4f434, 32'hc290a2d1, 32'h43080465},
  {32'hc4a6a722, 32'h435109bd, 32'h42a87d6c},
  {32'h44354fd2, 32'hc40f2d2e, 32'hc1d13ef6},
  {32'hc4041a5e, 32'h42ec3dda, 32'h43209d7e},
  {32'h44c7e514, 32'hc3c835cc, 32'hc2467a96},
  {32'hc327d9b5, 32'h42e4cb77, 32'h42f61468},
  {32'h450f89ec, 32'hc34a7505, 32'h42112a55},
  {32'hc1cd4800, 32'hc31ac748, 32'hc3e9fb65},
  {32'h442d2747, 32'h43dd5953, 32'hc167b211},
  {32'hc4995582, 32'h43973192, 32'h43c2e008},
  {32'h45279d4f, 32'h4183e642, 32'h4322e89e},
  {32'hc45b988a, 32'hc3253149, 32'hc30894b4},
  {32'h448102f6, 32'hc42bd522, 32'hc2a0542e},
  {32'hc482f1c4, 32'h428a48c9, 32'hc1f06e8e},
  {32'h44fc99ae, 32'hc2039758, 32'h42e01b15},
  {32'hc36de2a0, 32'h41169a1a, 32'h43f37941},
  {32'h441cd615, 32'h42a6ad00, 32'h41aadbe4},
  {32'hc3a7efee, 32'h427e47b0, 32'hc385aab5},
  {32'h44495eef, 32'hc1f489a8, 32'h42ceefcb},
  {32'hc407d76b, 32'hc2ab5036, 32'h4135613e},
  {32'h4467aed3, 32'h4330b4bf, 32'h4317768a},
  {32'hc4bc75c6, 32'h430ce148, 32'hc205c616},
  {32'h44e2650e, 32'hc4195213, 32'hc40ca90d},
  {32'hc4339638, 32'hc4058ffb, 32'hc38d5a55},
  {32'h44bf8941, 32'h4386afe7, 32'hc3a06a9b},
  {32'h4280c8c8, 32'hc32201c6, 32'h42fe9f44},
  {32'h43c4eb1d, 32'h4187948c, 32'h4324db9a},
  {32'hc466b232, 32'h4375151f, 32'h44037167},
  {32'h44a4a492, 32'hc263f32f, 32'hc36a9db2},
  {32'hc3958010, 32'hc229d957, 32'h423a1a92},
  {32'h43264240, 32'hc36d9efa, 32'h43f8358d},
  {32'hc449384a, 32'h3ff74916, 32'hc31672a7},
  {32'h43b128b8, 32'h43b436f3, 32'h421bd3e0},
  {32'hc4014dd4, 32'hc3a32709, 32'h43007ff4},
  {32'h42db79b0, 32'hc38f3e89, 32'h429ca456},
  {32'hc2e57063, 32'hc308a9f7, 32'h42c06e6a},
  {32'h4452e957, 32'h43cb9b53, 32'h437a3ff9},
  {32'hc50ee3c8, 32'hc31d1f8a, 32'h43331acf},
  {32'h44c040ab, 32'h433d033b, 32'hc28eb412},
  {32'hc3ee017c, 32'h4201e997, 32'h414e012c},
  {32'h438df070, 32'hc2498b5d, 32'hc292a44a},
  {32'hc3afcdd4, 32'hc316f1d1, 32'hc35a554b},
  {32'h44fbb782, 32'h43a154bf, 32'hc2bde7bc},
  {32'hc3689006, 32'h42a91d98, 32'h431fade7},
  {32'h43a04b08, 32'h42187959, 32'h436ef245},
  {32'hc51de3bb, 32'h434c9e08, 32'h4355c66e},
  {32'h448f2dc6, 32'h42e8ecee, 32'hc22dd196},
  {32'hc461ba19, 32'hc30fb5fd, 32'hc2c67f36},
  {32'h44fad812, 32'hc2f60596, 32'h4361cd8e},
  {32'hc4db7538, 32'h43410168, 32'h4297c241},
  {32'h44c1af41, 32'h429325ed, 32'h42fb412b},
  {32'hc5222471, 32'hc3366399, 32'h42fddf4f},
  {32'h45103690, 32'hc3c06c09, 32'h43cc9956},
  {32'hc445b824, 32'h430aa42b, 32'h43f5982a},
  {32'h44239810, 32'hc225544b, 32'h43691c2c},
  {32'hc4976885, 32'hc1286016, 32'hc2d5c35c},
  {32'h4445e9bc, 32'hc376bf64, 32'h43871093},
  {32'hc4fc25c7, 32'hc07c26ae, 32'hc2eee4c3},
  {32'h4390aa1e, 32'hc2b5875d, 32'h434977b7},
  {32'hc522ae2d, 32'hc1019114, 32'hc316a2c4},
  {32'h4508e31a, 32'h43839835, 32'h43c490a2},
  {32'hc4eeb6b7, 32'hc192bdb7, 32'h41a3a762},
  {32'h44e54a12, 32'h431a8447, 32'h42d96d5d},
  {32'hc4cc5cab, 32'h4026e8d8, 32'hc352a446},
  {32'h438e4180, 32'hc3340375, 32'hc34a3e34},
  {32'hc4be5c16, 32'hc23dc313, 32'h4308a95d},
  {32'hc22b6280, 32'h435a3cd4, 32'hc2e2c211},
  {32'hc4cda394, 32'hc24d69ce, 32'hc405cc2b},
  {32'h435854e0, 32'h43866b3a, 32'hc2fbb5f0},
  {32'hc4f3990a, 32'hc289b6ce, 32'hc3ada30d},
  {32'h44106638, 32'h4419c45c, 32'h41ce7936},
  {32'h433922a0, 32'hc39877b8, 32'h43238890},
  {32'h449d0fd0, 32'h42c3b35d, 32'hc39c2be2},
  {32'hc506e232, 32'hc3934c7c, 32'h43c442ed},
  {32'h450a59f4, 32'h432a47a3, 32'hc2eeebfe},
  {32'hc501471a, 32'h43931f4b, 32'h42c77028},
  {32'h44947147, 32'hc3a78572, 32'hc1676cb0},
  {32'hc4f46ab6, 32'hc36d86d9, 32'h424c9fdc},
  {32'h44ce1dfc, 32'h43940bd8, 32'h43c6d3bc},
  {32'hc5102384, 32'hc306d6b2, 32'h415719b4},
  {32'h44982f22, 32'hc34e3f8b, 32'hc3607147},
  {32'hc3383688, 32'h4338331a, 32'hc1bcd183},
  {32'h43d610f2, 32'h42e29821, 32'hc262922f},
  {32'hc3ecb549, 32'hc2b73887, 32'hc3894140},
  {32'h4526d2a6, 32'hc20e25a1, 32'h42bdb4a7},
  {32'hc4e3b9cb, 32'hc25bdbbf, 32'hc2665740},
  {32'h4511d385, 32'h4304fc1d, 32'h41a33dec},
  {32'hc502742d, 32'hc0e5d073, 32'hc249ca70},
  {32'h442f9060, 32'h4357defb, 32'hc31c3b60},
  {32'hc3153cfc, 32'h439510fc, 32'hc4083a5c},
  {32'h43d2d070, 32'hc28607bc, 32'h438ac94e},
  {32'hc4b9c797, 32'h4232ede5, 32'hc291f89e},
  {32'h4513b13b, 32'hc27a3bda, 32'h4288190f},
  {32'hc3afc440, 32'h3fe7073c, 32'hc34a3d13},
  {32'h4503fc7e, 32'hc3242afc, 32'hc2a825c5},
  {32'hc4b13490, 32'h4310652f, 32'hc2bc1ced},
  {32'h44b9c857, 32'h424609ea, 32'hc42155f7},
  {32'hc516d203, 32'hc36a8909, 32'hc1cf2e88},
  {32'h43c750a6, 32'h41928fe7, 32'hc29f874d},
  {32'hc387c228, 32'hc3213ce0, 32'h42d56a13},
  {32'h4389964a, 32'hc334bd9b, 32'hbfb5b6f2},
  {32'hc3c469f0, 32'hc3b846c9, 32'hc3094964},
  {32'h43d89528, 32'h41e863c6, 32'h42ba3f08},
  {32'hc416dc3c, 32'hc3871334, 32'h4319a900},
  {32'h448fbec3, 32'hc3756059, 32'h43816cbb},
  {32'hc4accb74, 32'hc2ab6ba3, 32'h43ba180b},
  {32'h4503b83b, 32'h436a3ed8, 32'hc15229c4},
  {32'hc43e3407, 32'hc18ff8d1, 32'h43a478ed},
  {32'h451e97bd, 32'hc3a319ff, 32'hc36dc5f0},
  {32'hc4e4097a, 32'hc371eaa4, 32'h432e4b87},
  {32'h44f60c7c, 32'h435d135e, 32'h43c4f429},
  {32'hc4caf92a, 32'h43ba8661, 32'hc1e4fb86},
  {32'h43082f40, 32'h42939400, 32'h431f7606},
  {32'hc3b42418, 32'h43a8a91d, 32'hc31f7893},
  {32'h44786b0e, 32'hc2989e40, 32'hc38562cc},
  {32'hc43e04a6, 32'h438cba12, 32'h42b0fcdd},
  {32'h45079a6b, 32'hc252f050, 32'h438f4797},
  {32'hc4aa0153, 32'hc2c9b0b2, 32'h437bf388},
  {32'h44d11118, 32'h439875c9, 32'hc3551d48},
  {32'hc509fe41, 32'hc1c6ac53, 32'hc2f5c223},
  {32'h45184cc4, 32'hc4085289, 32'hc392a746},
  {32'hc4a51274, 32'h42de7f49, 32'h4318dbaf},
  {32'h445ff4d4, 32'hc3fadb96, 32'h403f8f78},
  {32'hc3c90820, 32'hc3a409cd, 32'h428a7dfe},
  {32'h451d152f, 32'h43816d61, 32'hc3368e5a},
  {32'hc2c50d34, 32'hc255d26c, 32'hc2842131},
  {32'h43fd7f38, 32'h42d6e686, 32'h419c1083},
  {32'hc4ae5320, 32'hc2109ee4, 32'h435124e5},
  {32'h44f71648, 32'h437ecce6, 32'h4358674c},
  {32'hc5118c5f, 32'hc28c026b, 32'hc189bfcf},
  {32'h43bc75ac, 32'hc2aaa435, 32'h43163c75},
  {32'hc4e88490, 32'h4265886c, 32'hc3a162b0},
  {32'h442cf288, 32'h415a929e, 32'h43c9293d},
  {32'hc5205ffc, 32'hc2245be8, 32'hc2625934},
  {32'h4495c651, 32'hc370882e, 32'hc38e3672},
  {32'h4382166c, 32'hc3cf8183, 32'hc3b3b904},
  {32'h451ba7ee, 32'h438e525e, 32'h420a19e8},
  {32'hc3534490, 32'hc3088112, 32'h43bdce81},
  {32'h434e27d6, 32'hc1d50929, 32'h4275a2c1},
  {32'hc467c872, 32'hc3829de5, 32'h42f36acd},
  {32'h44f641f3, 32'hc3504b7a, 32'hc39356b4},
  {32'hc2f29e06, 32'hc30f2c2f, 32'h42d3718d},
  {32'h44df8dcb, 32'h4331100c, 32'h428c0f6c},
  {32'hc28a5400, 32'h435df657, 32'h42a279f8},
  {32'h44f6c022, 32'hc3de7272, 32'h42d7ce21},
  {32'hc4df6cb5, 32'h43b55822, 32'hc3102630},
  {32'h44d6bcfd, 32'h4363a20f, 32'hc2fc00fd},
  {32'hc495da7a, 32'h424dd3a5, 32'hc392189f},
  {32'h44c02f67, 32'hc304a22c, 32'h42805c81},
  {32'hc4a30d5e, 32'h42e2dd9b, 32'hc41d2c5e},
  {32'h4507baa6, 32'h42ec7836, 32'h432ee7f2},
  {32'hc4316a72, 32'hc39bc2c7, 32'hc3d19dca},
  {32'h444403a6, 32'hc375777e, 32'h41a8e3e7},
  {32'hc5075304, 32'hc141411c, 32'hc30afa21},
  {32'h44e82ebf, 32'h42c210d8, 32'h42d69402},
  {32'hc31c3100, 32'hc36c1c6c, 32'hc3bdea24},
  {32'h442932cc, 32'hc23a5998, 32'h43c39ec3},
  {32'hc4e4a169, 32'hc2d9be7e, 32'hc377b97e},
  {32'h4459680b, 32'h43390c02, 32'h43d296cd},
  {32'hc3a6019b, 32'hc3f8fa93, 32'hc30660d5},
  {32'h4498789a, 32'hc25f4317, 32'hc2582f40},
  {32'hc4de8f86, 32'h42df851f, 32'h43dbae23},
  {32'h449f1030, 32'h4227ebae, 32'h439416eb},
  {32'hc4834693, 32'hc2fe9871, 32'hc1a02daf},
  {32'hc26a1e68, 32'h43931e97, 32'h42700d5a},
  {32'hc4b9cc62, 32'h4333c9cc, 32'hc251135f},
  {32'h42f242a0, 32'h421c8319, 32'h42e03727},
  {32'hc4fda9fd, 32'hc3d95afc, 32'hc0dc7c91},
  {32'h44355540, 32'h4353467f, 32'h4317c3f5},
  {32'hc4339aea, 32'hc22225c0, 32'hc2c15a80},
  {32'h440a77c9, 32'hc1e603f1, 32'h4378b827},
  {32'hc4fb444e, 32'h43c57d4a, 32'hc36d94d6},
  {32'h43b995e4, 32'h4381f92b, 32'hc1aaa88d},
  {32'hc44ac46a, 32'h437994e4, 32'hc3a1f5c0},
  {32'h441ee94b, 32'h425725ad, 32'h43929aa3},
  {32'hc3dac2bd, 32'hc323f0f0, 32'hc1fc84ea},
  {32'h451c9c2b, 32'h4300f5d6, 32'hc1ee4ed2},
  {32'hc4e2744f, 32'h42c76b42, 32'h428153e5},
  {32'h448209bf, 32'h4331d2d6, 32'h3ff31390},
  {32'hc3bea1f8, 32'hc3326635, 32'hc3d17c9b},
  {32'hc46a23b1, 32'h42a4ab2f, 32'h4350b916},
  {32'h44ba95a1, 32'hc2ac37ea, 32'hc1fceaf2},
  {32'hc4838475, 32'hc2961b5d, 32'hc386a039},
  {32'hc3787dc8, 32'h42167660, 32'h429e5e9f},
  {32'hc4c0f891, 32'h4344b9a1, 32'hc3bafa71},
  {32'h44e6bfaa, 32'h438ad52a, 32'hc3b23f40},
  {32'hc466d5e6, 32'h434f2f11, 32'hc37cd2ef},
  {32'h442438ca, 32'hc237db90, 32'h43ea685b},
  {32'hc31af930, 32'hc2ddb91c, 32'h42586031},
  {32'hc30c9838, 32'h42021dc0, 32'hc3a4a43f},
  {32'hc488d37e, 32'h433a6fc9, 32'h42d6fec0},
  {32'h43d2f598, 32'h43bac2e9, 32'h43b91ca3},
  {32'hc386e0e0, 32'h434bd2e4, 32'h41cbb052},
  {32'h432e4f00, 32'h435a3879, 32'h43ba331f},
  {32'hc4c354f3, 32'h42961bcd, 32'hc26226d1},
  {32'h42fe7f80, 32'hc22bb199, 32'h4189021b},
  {32'hc4f74bbf, 32'h42e16e7d, 32'h42e5a038},
  {32'h4255f4a0, 32'hc0a51e48, 32'h43ca32c1},
  {32'hc485b16a, 32'h43222a44, 32'hc38582f3},
  {32'h4459fce3, 32'hc3a5e4ec, 32'h412f5ac0},
  {32'hc491a44b, 32'hc34c7c98, 32'hc3a34b3e},
  {32'h44db2a77, 32'hc1e38112, 32'h43ae1ba4},
  {32'hc505f2a2, 32'h42d16655, 32'hc3754a6c},
  {32'h44dc9172, 32'hc2d47e0d, 32'hc3422aa0},
  {32'hc4f56cd9, 32'h43222c3b, 32'h42de9ea1},
  {32'h451c8d03, 32'hc3336afa, 32'h43082d83},
  {32'hc4918aaa, 32'hc31eb3fd, 32'hc2a45ca0},
  {32'h44ef5c27, 32'h4303a42a, 32'h42929f65},
  {32'hc485f29e, 32'hc3c305ff, 32'hc1ad34e6},
  {32'h43145270, 32'hc238b70c, 32'hc370aaee},
  {32'hc4b220f3, 32'h432bcf94, 32'h42b5baf8},
  {32'h44822176, 32'hc3dcb930, 32'hc3011165},
  {32'hc4bec188, 32'hc294d148, 32'h43431310},
  {32'h43254fb0, 32'h43245f85, 32'hc32bcf67},
  {32'hc50f5cc7, 32'hc2a3f49b, 32'hc31f5e51},
  {32'h43efce0e, 32'h418d1a1b, 32'hc30e80ef},
  {32'hc493e5c0, 32'hc3902e1f, 32'hc235e646},
  {32'h435385bb, 32'h422a5b41, 32'hc36e2652},
  {32'hc4d40e70, 32'hc347d658, 32'h42fe139d},
  {32'h4487b8a9, 32'hc3a24b97, 32'hc3640008},
  {32'hc4cdfd96, 32'hc3836eff, 32'hc277eeb8},
  {32'h44b1fb48, 32'h42a8db20, 32'h42c18c1f},
  {32'hc405e1b9, 32'hc3c6151c, 32'hc202923b},
  {32'h448fa85f, 32'hc37d6943, 32'h433f6116},
  {32'hc4ef01f4, 32'h43eb8863, 32'h42f21123},
  {32'h445732c2, 32'h42cf6e8d, 32'hc25f855f},
  {32'hc447f6e4, 32'h42b5f0a6, 32'hc32cb2b0},
  {32'h441566c4, 32'hc22dab50, 32'hc37fff7c},
  {32'hc4973e07, 32'h42d1ba3f, 32'h41c3c138},
  {32'h3e9dfc80, 32'hc30d90c1, 32'hc3ee0e78},
  {32'hc388a018, 32'h43238cf5, 32'h42ece9d1},
  {32'h44955720, 32'h43833214, 32'h42d2e669},
  {32'hc4f25510, 32'hc3b4a7d1, 32'hc3562a67},
  {32'h4384ed32, 32'hc302ea09, 32'h43579bc8},
  {32'h4339e468, 32'hc3df2494, 32'h42f200b3},
  {32'h450b9f04, 32'hc3722f7a, 32'hc2394321},
  {32'hc47378e4, 32'h4315e6d7, 32'hc12c8d02},
  {32'h44a6b478, 32'hc3ab4bbe, 32'hc35164bb},
  {32'hc4346ba6, 32'hc3c15556, 32'hc3436578},
  {32'h44717dd4, 32'hc2030a8b, 32'h43ee6ff5},
  {32'hc3ce1028, 32'hc3b53034, 32'hbfcd0878},
  {32'h440ab2da, 32'hc2e4b1ac, 32'hc363aea3},
  {32'hc40c1294, 32'hc2e95ff7, 32'h4263048a},
  {32'h44cbe3f4, 32'h42d1e304, 32'h433a6fda},
  {32'hc50b9a28, 32'h43a1bd66, 32'hc3abd78d},
  {32'h449a52d9, 32'h40994fab, 32'h439f399e},
  {32'hc42c2e00, 32'hc302192e, 32'hc233b522},
  {32'h448d4da0, 32'h431da5dd, 32'hc3671efc},
  {32'hc5145c94, 32'hc37f34d8, 32'hc3e8a636},
  {32'h4483bb01, 32'h4163b315, 32'h42f843fa},
  {32'hc49a6585, 32'h42b930e8, 32'hc1cc2470},
  {32'h43404334, 32'hc3509e92, 32'h43bc1ea0},
  {32'hc416e5cd, 32'h41dc7283, 32'h43573d9e},
  {32'h44c19534, 32'h43174fec, 32'hc3a1c64b},
  {32'hc3a4564e, 32'hc33dbca7, 32'h42f1f5e4},
  {32'h443e59b3, 32'h433a4427, 32'hc2ed3304},
  {32'hc2b9481f, 32'hc38d5856, 32'hc31c3b14},
  {32'h41bc6f70, 32'h437be457, 32'hc2ac8ded},
  {32'hc4a6b7a7, 32'hc35db0f4, 32'h4290a93d},
  {32'h44f52676, 32'h42c15bc8, 32'h431dd481},
  {32'hc34d31f0, 32'h4220c6fe, 32'hc33beceb},
  {32'h44d70877, 32'hc402d7b9, 32'h43936199},
  {32'hc4046b04, 32'hc312c73a, 32'h43abb0a9},
  {32'h44e7ed89, 32'h43bbb32a, 32'h429520c0},
  {32'h43872f7a, 32'hc194dd81, 32'h43596928},
  {32'hc2e32fb0, 32'hc3eeee32, 32'hc2b6b724},
  {32'hc45ed9b8, 32'h43146d0f, 32'h431047c1},
  {32'h44bbc5e0, 32'hc3c5e23e, 32'hc22b13d8},
  {32'hc5151d8f, 32'h42e67d3c, 32'hc3911393},
  {32'h450fc095, 32'hc314b8f6, 32'hc2b0078b},
  {32'hc43d06d1, 32'hc332e496, 32'h438e8953},
  {32'h4481f21f, 32'hc3154c6c, 32'hc2ed48fc},
  {32'hc4e72d8a, 32'hc38d6833, 32'h42ae3801},
  {32'h4503977f, 32'h427281cf, 32'h412e6f9c},
  {32'hc4967a66, 32'h413adf14, 32'hc24bae37},
  {32'h4436833a, 32'h433a02b4, 32'hc3006d27},
  {32'hc2ea2cd9, 32'hc3d90472, 32'h42aac1b4},
  {32'h45001fb6, 32'h430d608a, 32'hc3e29bc0},
  {32'hc5041cf0, 32'hbeea7dd0, 32'h42681e5f},
  {32'h44bedca6, 32'h425e071d, 32'hc39745e9},
  {32'hc4b69557, 32'h439cc07d, 32'h431a5553},
  {32'h442d6e58, 32'h4389b5ae, 32'hc2b5b230},
  {32'hc3a79762, 32'h41a75680, 32'hc2f58182},
  {32'h448f3e89, 32'h4399b288, 32'hc28379e4},
  {32'hc2802370, 32'hc40da7f6, 32'hc315b86e},
  {32'h4472ea14, 32'hc380e675, 32'h43289bb6},
  {32'hc510a738, 32'h421e3e22, 32'h4282b7e1},
  {32'h440bf066, 32'hc398cf65, 32'h4378fc68},
  {32'hc5012462, 32'hc3946418, 32'h43d80848},
  {32'h4488f05b, 32'h438f6767, 32'h42f1fcc5},
  {32'hc4a5a448, 32'hc41d4590, 32'h4381e954},
  {32'h44accf08, 32'h432e87e1, 32'hc3559c38},
  {32'hc506704d, 32'hc3c49aae, 32'hc3078f00},
  {32'h44116170, 32'hc40a1742, 32'hc3a271b9},
  {32'hc49137d2, 32'h430f1865, 32'h4393f57d},
  {32'h4428f2e4, 32'h42483878, 32'hc352074a},
  {32'hc5118714, 32'hc4214a7f, 32'h42f2829e},
  {32'h43c21cac, 32'hc23703f6, 32'hc3275ad1},
  {32'hc47dc644, 32'hc365fec3, 32'h43158c06},
  {32'h43dc2ee9, 32'h423e78f0, 32'hc3a74d16},
  {32'hc494b598, 32'hc2fee59a, 32'h4303788d},
  {32'h4495f5fa, 32'hc270bbc0, 32'hc389bd94},
  {32'hc45279a4, 32'h433718d0, 32'h43d39475},
  {32'h44f77f41, 32'h434b5498, 32'h433f2c6b},
  {32'hc4493aff, 32'hc1ef9460, 32'hc2a67f7a},
  {32'h442313b2, 32'h431ede17, 32'hc366c100},
  {32'hc486db64, 32'h42e94918, 32'hc3100da4},
  {32'h4450ee3c, 32'hc23e7e76, 32'h43681733},
  {32'hc48ad5b5, 32'hc3d51027, 32'hc25ce015},
  {32'h4503d22e, 32'h432132c8, 32'h42ec473a},
  {32'hc4342d62, 32'hc330a413, 32'h4361e0ac},
  {32'h44de8f50, 32'hc3a54823, 32'h43789da0},
  {32'hc42a0723, 32'h42c6fc8c, 32'hc3820b19},
  {32'h44a3ebd2, 32'h43d63be5, 32'hc1aa44ae},
  {32'hc4e2100b, 32'h43458c36, 32'h4387d74f},
  {32'h42848550, 32'hc3ace81f, 32'hc3e0cb76},
  {32'hc4e35dd6, 32'h43842002, 32'h4327cac3},
  {32'h44cb8048, 32'hc2c1ca2b, 32'h43011f8b},
  {32'hc486dbec, 32'hc30fa62d, 32'h439966cb},
  {32'h44e01c1f, 32'h43c1160c, 32'hc3846a92},
  {32'hc4d4069e, 32'hc35efca2, 32'hc155530f},
  {32'h44ea2c0c, 32'h43917fb1, 32'h43807516},
  {32'hc4cc318f, 32'hc2b80985, 32'h43748eae},
  {32'hc3a9e72c, 32'hc2db9ff8, 32'hc2a0297e},
  {32'hc4a4b793, 32'hc38f3657, 32'h42971460},
  {32'h44a5e574, 32'hc2dd74fd, 32'h4378644d},
  {32'hc4b90b6d, 32'h434b47ca, 32'hc11adc4c},
  {32'h44d1f5ee, 32'h42f3b5a1, 32'h4282b877},
  {32'hc31adba8, 32'h4232a994, 32'h422c4aa2},
  {32'h444285ab, 32'h4354023a, 32'h4293d990},
  {32'hc3f7a99d, 32'hc1f13086, 32'h43034b5d},
  {32'hc2b6ebac, 32'h42bb6091, 32'hc3835969},
  {32'hc508e4b8, 32'hc2c00d00, 32'hc2bdad3a},
  {32'h44f6c515, 32'hc22b8d9a, 32'hc3840eba},
  {32'hc3d1011c, 32'hc325aa9b, 32'hc3ce601e},
  {32'h444ad734, 32'hc19a19f2, 32'h40bc6e98},
  {32'hc4facbad, 32'h42ab3a1f, 32'h431133b7},
  {32'h44f90d1a, 32'h431e75bb, 32'h4373de33},
  {32'hc273ed80, 32'h43d42d3a, 32'hc28e81fc},
  {32'h443216d2, 32'hc2eb3fa6, 32'h42c37bdd},
  {32'hc43adb16, 32'hc30608c6, 32'h437e198f},
  {32'h4517c6c8, 32'hc2ebb60a, 32'h43627633},
  {32'hc4bb4e1e, 32'h431abab7, 32'h41aba2b3},
  {32'h44340d31, 32'hc3b89b2c, 32'hc32ccf7a},
  {32'hc4044c80, 32'h43972b28, 32'h440debad},
  {32'h448cd781, 32'hc25b2694, 32'hc31ae6d6},
  {32'hc438efaa, 32'hc3917d4b, 32'h437bb32e},
  {32'h449e7eef, 32'h4356b0ce, 32'hc2cef573},
  {32'hc4da4f4f, 32'h434c9c57, 32'hc32b30bf},
  {32'h4428f0c4, 32'hc36498bc, 32'hc4010327},
  {32'hc5099c52, 32'hc191998a, 32'hc2884219},
  {32'h439043e0, 32'hc2f922a6, 32'h429a82b9},
  {32'hc4a830cd, 32'h431937e4, 32'h4392f943},
  {32'h43d494af, 32'hc2e6059c, 32'hc2dcf005},
  {32'hc4af68da, 32'h41f7d4cb, 32'h4377d57e},
  {32'h42bd40dc, 32'h4368d207, 32'hc17b68da},
  {32'hc4fa9f68, 32'hc3d5f3a1, 32'hc389d972},
  {32'h44886cf4, 32'h4344e988, 32'h437027ba},
  {32'hc4cf6c67, 32'hc2f8ce1e, 32'hc362dd02},
  {32'h445723f6, 32'hc3260689, 32'hc19db4a7},
  {32'hc3ea6cb0, 32'hc34119cd, 32'hc3d44e98},
  {32'h44cf4159, 32'hc41a118a, 32'h4182a80f},
  {32'hc4d5d071, 32'hc231b529, 32'hc33a49e6},
  {32'h43eab590, 32'h438db1bc, 32'hc330be86},
  {32'hc4eeb8ce, 32'hc369e8eb, 32'hc142ec8a},
  {32'h42e104a4, 32'h4309c99f, 32'h42a97fc9},
  {32'hc4c4bd5d, 32'h4308e749, 32'hc1878e39},
  {32'h44903ff1, 32'hc2b1dbf1, 32'h42e02150},
  {32'hc4e45058, 32'hc0250fbd, 32'h41d29c50},
  {32'hc1e917ce, 32'hc3038040, 32'hc2750b6c},
  {32'hc4d652f4, 32'hc2bb4802, 32'hc306e39a},
  {32'h44445702, 32'h437a784e, 32'hc3a2bd83},
  {32'hc41367d7, 32'h425cfcb6, 32'hc3cb8e4d},
  {32'h43c6bade, 32'hc31b1a47, 32'h4386f8cb},
  {32'hc4a71c9d, 32'hc3039106, 32'hc3b1f9ec},
  {32'h445354b1, 32'hc32f93b2, 32'h43270c7b},
  {32'hc4e4bc3f, 32'hc1fc8c06, 32'hc2b90f10},
  {32'h44a72ad4, 32'hc3285c62, 32'hc269a23c},
  {32'hc4af263e, 32'hc3059762, 32'h43995038},
  {32'h44822868, 32'hc39453af, 32'h43976354},
  {32'hc2da21e0, 32'h4340bafc, 32'h43068973},
  {32'h44808974, 32'h415ea984, 32'h4350d207},
  {32'hc49fd181, 32'hc20fa7eb, 32'hc1f40fd7},
  {32'h43036438, 32'hc395f1c2, 32'h43384be0},
  {32'hc4f8de15, 32'h42c523ae, 32'h42f4058f},
  {32'h444e5a60, 32'h42db81f8, 32'hc313c005},
  {32'hc422f142, 32'h4369e18a, 32'h43afbb68},
  {32'h44af87fa, 32'hc2961750, 32'hc312962f},
  {32'hc5070eae, 32'h434e0a9b, 32'hc2d9f02b},
  {32'h43af8d60, 32'hc254c352, 32'h402171b0},
  {32'hc51d4ca8, 32'hc315865d, 32'h436e58ed},
  {32'hc2a51d35, 32'h41b714f4, 32'h4302b1e6},
  {32'hc4d6c45a, 32'h43af7db1, 32'h43420113},
  {32'h45053705, 32'h43bf1d7a, 32'h41f8f50e},
  {32'hc483f63f, 32'hc0c15fdc, 32'h42535a7f},
  {32'h44e5220d, 32'h437abf0f, 32'hc25a8644},
  {32'hc4aa6d54, 32'hc3f3dfb6, 32'hc2d54de8},
  {32'h441d2af5, 32'h3f2f8c5c, 32'h4400e94a},
  {32'hc2d6442c, 32'hc3879a78, 32'hc3d35ec1},
  {32'h4485bb45, 32'h440586ad, 32'h440a828b},
  {32'hc33a26d8, 32'h43820594, 32'hc3a03671},
  {32'h4488fb2d, 32'h418c64ce, 32'hc3018eb7},
  {32'hc4b17a38, 32'hc246046e, 32'h42a06809},
  {32'h45039db7, 32'h434aadc3, 32'hc337079e},
  {32'h4365a38c, 32'h420b7c50, 32'h424f314f},
  {32'h450d02e2, 32'hc3b31cc6, 32'h435adf6c},
  {32'hc50e3ab3, 32'h435dd703, 32'h42757762},
  {32'h4500a92c, 32'h432b89cc, 32'h4321a81d},
  {32'hc4ecebcc, 32'hc346fc95, 32'hc1a6af68},
  {32'h450de51b, 32'hc32e603b, 32'h437a3250},
  {32'hc4525038, 32'hc28a18e0, 32'h41bf9da4},
  {32'h445e69bf, 32'hc3942263, 32'hc3592e8c},
  {32'hc408638f, 32'hc3a0e9b6, 32'h430e1430},
  {32'h4397c8c2, 32'hc37f98d5, 32'h436c46aa},
  {32'h42b82460, 32'h42d0543f, 32'hc3906f5a},
  {32'h43849418, 32'hc21cb936, 32'hc38038a7},
  {32'hc4862c6e, 32'hc2feac78, 32'hc354bf64},
  {32'h44aadfaa, 32'h42e251ff, 32'h42d3a2da},
  {32'hc4a5e32a, 32'hc335f349, 32'h42b2ef85},
  {32'h45052243, 32'h42ec7e71, 32'h42d6da45},
  {32'hc405a787, 32'hc2fd730f, 32'hc39e38f2},
  {32'h4405ebe6, 32'hc118dc89, 32'h423c6e6e},
  {32'hc4d4c99a, 32'h42f12f61, 32'hc264a29c},
  {32'h42ccba82, 32'h43363cb2, 32'hc3866643},
  {32'hc4b3f920, 32'h43246a13, 32'hc26fd4ea},
  {32'h44ad3bf2, 32'hc39187a3, 32'h429a5664},
  {32'hc49a76be, 32'h42366960, 32'hc392a12a},
  {32'h447a03d4, 32'hc376e003, 32'hc239075a},
  {32'hc3e65800, 32'hc38175d0, 32'h422e7e97},
  {32'h4432bb83, 32'h431f6ee7, 32'h420d2972},
  {32'hc4bf5a58, 32'h43736345, 32'h43a33c78},
  {32'h44761511, 32'h41013106, 32'h43697aa7},
  {32'hc49747e2, 32'hc3acc544, 32'h432315ec},
  {32'h44177598, 32'h43869ba7, 32'hc2f18e07},
  {32'hc3dc96d9, 32'hc395a8b3, 32'hc3172c67},
  {32'h43fe4e2c, 32'h43a74da8, 32'h433f1196},
  {32'hc2eb5446, 32'h428b2e48, 32'h438122a0},
  {32'h4503b177, 32'h43445fc0, 32'hc2e55ac3},
  {32'hc50a1ca9, 32'h431891d3, 32'hc35ffb06},
  {32'h44b94afc, 32'hc350408e, 32'h43937f03},
  {32'hc40713fe, 32'h438b8de5, 32'hc3d9e4fe},
  {32'h44ebb46e, 32'h42b73a79, 32'hc34f8d28},
  {32'hc43a4f48, 32'h431951b6, 32'h43672b52},
  {32'h4467f0ea, 32'hc376a491, 32'hc1a8bd8c},
  {32'hc502deae, 32'hc29560eb, 32'hc367e027},
  {32'h449ca2ec, 32'h434ad2af, 32'hc1ad4cb0},
  {32'hc42a9c32, 32'hc380b1ac, 32'hc2dd9860},
  {32'h44078484, 32'h437a64dd, 32'h4339b3a1},
  {32'hc4c44ecc, 32'hc22f9ccd, 32'h42e2539b},
  {32'h4420e332, 32'h42a1f758, 32'hc29d4cca},
  {32'hc3f61328, 32'h438d88d4, 32'hc0db34ce},
  {32'h45046c92, 32'h429f1eee, 32'hc3864834},
  {32'hc4429488, 32'hc18999b8, 32'hc2df1caf},
  {32'h450358b1, 32'hc2556787, 32'h42db4815},
  {32'hc4c84b36, 32'hc3a31980, 32'hc33a8d20},
  {32'h44a105be, 32'h420fba27, 32'h43c04d65},
  {32'hc4825639, 32'h43245187, 32'h43688831},
  {32'h44e900d3, 32'hc2160fd8, 32'h43191d1f},
  {32'hc47b9510, 32'hc1be45db, 32'h3f7cf405},
  {32'h451294d7, 32'hc1bdfadb, 32'hc29ad4a0},
  {32'hc382d754, 32'h437a05b7, 32'h439def26},
  {32'h45126a86, 32'h4408ccc8, 32'hc1c1a1f4},
  {32'hc4c00518, 32'h420d9aad, 32'h426f3454},
  {32'h44ef4625, 32'hc18eb6c6, 32'hc39b8003},
  {32'hc3720500, 32'h433e225e, 32'h4383a462},
  {32'h44ed098e, 32'hc37b323c, 32'hc25da19d},
  {32'hc4b621a2, 32'h438e15d3, 32'hc244ea3d},
  {32'h446781e4, 32'hc37c92c5, 32'hc39536db},
  {32'hc3f7cf24, 32'h42a891eb, 32'h42e782e9},
  {32'h43c6fff0, 32'h4318927b, 32'hc3afb25f},
  {32'hc4fa0346, 32'hc2e0114d, 32'h43f09278},
  {32'h43fbb72d, 32'h43c79aeb, 32'hc38c6b17},
  {32'hc4563668, 32'h437ac6f6, 32'hc2ad675e},
  {32'h44bae3ae, 32'hc28825de, 32'h42c63268},
  {32'hc4578119, 32'h43bd4fc9, 32'hc2d69fa2},
  {32'h44def294, 32'hc22db4e6, 32'hc1cdee73},
  {32'h4395fa20, 32'h43a919c6, 32'hc29f9fe2},
  {32'h44c4b124, 32'hc31c7910, 32'hc26435ee},
  {32'hc415445c, 32'h42add087, 32'h431b1b53},
  {32'h44585770, 32'hc32130aa, 32'h432b0779},
  {32'hc4a57239, 32'h4226ff55, 32'hc2840d55},
  {32'h44252cc0, 32'h43dfa622, 32'hc28ee6bc},
  {32'hc39776ec, 32'hc351d0bb, 32'hc2745020},
  {32'h4464f0bc, 32'h4359e909, 32'hc2bf7830},
  {32'hc522254f, 32'h41be3b6a, 32'hc401b16c},
  {32'h447f325b, 32'h4343e008, 32'h4203cdef},
  {32'hc315b3c0, 32'h418190ca, 32'h429e0c4c},
  {32'h45179a36, 32'h42b4a695, 32'hc3872f91},
  {32'hc3583644, 32'h43b617e3, 32'hc289b858},
  {32'h440a675c, 32'h43345e81, 32'h44010684},
  {32'hc3cc33b0, 32'hc25d6147, 32'hc39476a4},
  {32'h44057315, 32'h4109ca24, 32'hc2adebef},
  {32'hc4cf4692, 32'h43b9f60c, 32'h41efdbbd},
  {32'h4406062c, 32'hc394f24e, 32'hc1f22e3a},
  {32'hc3f2fd60, 32'hc3ad0674, 32'h421e4634},
  {32'hc3954ae0, 32'h435a2076, 32'h41ac5b38},
  {32'hc4c17554, 32'hc2a8ce76, 32'h42dabc78},
  {32'h447676e6, 32'h43303546, 32'h43c81495},
  {32'hc4d36d8c, 32'h4318bc27, 32'h4340cf2f},
  {32'h44ff5b86, 32'h434d73e7, 32'h42dcc542},
  {32'hc42bdb0e, 32'h4418a584, 32'hc0b4ff08},
  {32'h43a5ad14, 32'h42eb2fb2, 32'hc1589506},
  {32'hc5164a04, 32'h431c7a3f, 32'h42f7b156},
  {32'h43f859ec, 32'h43b9dcdb, 32'h42551028},
  {32'hc4cd5f98, 32'hc222484a, 32'h4045d5f8},
  {32'h450bcbba, 32'h43db4d34, 32'h42dd60a4},
  {32'hc408c640, 32'h4322a073, 32'h43a0f298},
  {32'h43e29c14, 32'h4344b6e4, 32'h43b86c14},
  {32'hc507be0e, 32'h435b8612, 32'hc2db2580},
  {32'h44ce926d, 32'h430ab228, 32'h435dcb20},
  {32'hc47c27a7, 32'hc37db94e, 32'hc2b87c87},
  {32'h440cf2ea, 32'h43fa493b, 32'h42834367},
  {32'hc4f125b0, 32'hc3c07ef6, 32'h439f7cb8},
  {32'h44120a98, 32'hc29ac30e, 32'h42b7c7ea},
  {32'hc4e68f08, 32'h4330b7dd, 32'hc28974ce},
  {32'h440b8ad8, 32'h41686f72, 32'hc300387c},
  {32'hc358def0, 32'h42aa3b92, 32'hc295d2f7},
  {32'h43bdb740, 32'h42b3b008, 32'h431f26d6},
  {32'hc4914d11, 32'hc3d407cd, 32'hc10c43ed},
  {32'h44e6e3ee, 32'h4394c4ba, 32'hc30aee4e},
  {32'hc3fbafb5, 32'h43c2ff39, 32'hc341fe30},
  {32'h443bb9be, 32'h4136197a, 32'hc32c18ee},
  {32'hc4982145, 32'hc32884d9, 32'hc2b9a7f5},
  {32'h44ffebc4, 32'h4276e6fe, 32'h4303f06d},
  {32'hc511f326, 32'hc19d7921, 32'hc3d23b30},
  {32'h4500ebdb, 32'h4409315f, 32'hc3856ae8},
  {32'hc505f742, 32'h43734e1b, 32'hc2a58180},
  {32'h450c5823, 32'hc38cbe09, 32'hbe08937b},
  {32'hc3bc9fca, 32'hc2c84d1a, 32'hbebb5718},
  {32'h443764b5, 32'hc31481cd, 32'h423e0c3e},
  {32'hc47871b3, 32'h432b2cbf, 32'h43f88aab},
  {32'h44a26eb3, 32'hc2927d90, 32'hc35b50e2},
  {32'hc4246519, 32'h41a9ed11, 32'h42d487b7},
  {32'h44892c2e, 32'h42b66daf, 32'h41bad539},
  {32'hc1124220, 32'hc27a413c, 32'h43b2aa46},
  {32'h4379c1b0, 32'hc2582e31, 32'hc1b92d20},
  {32'hc3e1f820, 32'h427ad141, 32'hc37839e6},
  {32'h449b5d90, 32'hc3a517a5, 32'h41593220},
  {32'hc4627338, 32'h434c043c, 32'hc2bf207f},
  {32'h44e22ca7, 32'hc23138ce, 32'h43cb5463},
  {32'hc4df871b, 32'hc21380fc, 32'hc3415eae},
  {32'h44531052, 32'hbf8bcf98, 32'hc269eacf},
  {32'hc4a94b73, 32'hc359f1b3, 32'hc3a56bfa},
  {32'h4511914b, 32'h4339b23b, 32'h3fc5fb30},
  {32'hc454bf4e, 32'hc33104dd, 32'h429a9d80},
  {32'h4511d18d, 32'h41b9eeeb, 32'hc311183b},
  {32'hc4be077e, 32'hc3c936f0, 32'hc24354fc},
  {32'h44970c75, 32'h435aaf57, 32'hc2e9e7b8},
  {32'hc4eaf968, 32'hc31ca122, 32'h42fbf01a},
  {32'h44350f80, 32'h436c8c27, 32'h43ce9037},
  {32'hc401798d, 32'h4243925f, 32'hc3a166d4},
  {32'h44345d3a, 32'h44000b83, 32'h43de6dad},
  {32'hc4d740dd, 32'hc2acc091, 32'hc36936d1},
  {32'h4481cbf7, 32'hc390dea3, 32'h4220e750},
  {32'hc483dbeb, 32'h4130e369, 32'h433b33f2},
  {32'h43dacb00, 32'hc2a76c21, 32'h432649b2},
  {32'hc3d058a0, 32'h42987460, 32'h43e7a236},
  {32'h448eacf4, 32'h4372be2d, 32'hc3a1d0fd},
  {32'hc4d4ad7b, 32'hc36411ed, 32'h438af124},
  {32'h4422963c, 32'h428d5582, 32'hc355c5a2},
  {32'hc4b2b7d6, 32'hc2f4d9e0, 32'hc32b400e},
  {32'h4436d148, 32'h43699bee, 32'h41cff33f},
  {32'hc4e68fd1, 32'h42f879a4, 32'h43a06e9a},
  {32'h44e9432f, 32'hc3b4e92d, 32'h43183419},
  {32'hc49b381b, 32'h420d1622, 32'hc28e4c30},
  {32'h441ac124, 32'hc317e86e, 32'hc364f38c},
  {32'hc45c103e, 32'hc2d8a37b, 32'h3f741df7},
  {32'h44740618, 32'hc1d1719a, 32'h43831fa1},
  {32'h41bea280, 32'hc0ede368, 32'h438be83f},
  {32'h44e12131, 32'hc2a195b8, 32'h418b9fd6},
  {32'h42e75f20, 32'hc16408a8, 32'h419fc80c},
  {32'h436bc090, 32'h42d9ce48, 32'hc3883e54},
  {32'hc509082a, 32'hc313edc9, 32'hc2916a4b},
  {32'h448bc659, 32'h43780d33, 32'hc362ba4a},
  {32'hc4d98c2c, 32'h4308a6a1, 32'hc32bf6af},
  {32'h4515d451, 32'h42400026, 32'h438ef861},
  {32'hc4f022be, 32'h438c015c, 32'h42be67ba},
  {32'h43d3f2d5, 32'h430332a6, 32'h43563d7b},
  {32'hc49d89ec, 32'hc3a07d94, 32'h43c111ab},
  {32'h4481d352, 32'h43ec3481, 32'hc33022b1},
  {32'hc50b3672, 32'h42f402be, 32'h42a27d7d},
  {32'h44b9505a, 32'h438d6c6e, 32'hc315cb0e},
  {32'hc3023ed9, 32'hc2630231, 32'h4383e1d5},
  {32'h449ed8d0, 32'h424d8137, 32'hc382b08d},
  {32'hc5151bea, 32'h42a7bfc7, 32'h41717165},
  {32'h43e71a04, 32'hc2049c12, 32'hc37a9fb5},
  {32'hc47d6a9c, 32'hc2465f43, 32'h42e6fa9d},
  {32'h442aacba, 32'hc299082c, 32'hc0937481},
  {32'hc4806070, 32'hc33dfb7e, 32'h438e6a23},
  {32'h445776b3, 32'h432835e4, 32'hc3dde0a0},
  {32'hc4bcd3d8, 32'h4254f703, 32'hc31aa5de},
  {32'h44db90ca, 32'hc3047239, 32'h42ecfcbc},
  {32'hc450a3e6, 32'hc2d4d528, 32'hc38e62b9},
  {32'h44eccca8, 32'hc3385d4e, 32'h42fdc2d2},
  {32'hc2d16590, 32'h43871835, 32'hc1b9bb4d},
  {32'h443098a8, 32'h42039b80, 32'h41e10910},
  {32'hc4f76bd6, 32'h43823795, 32'hc243a14c},
  {32'h43e3f468, 32'hc2f64985, 32'hc2ef14fb},
  {32'h4310cb96, 32'h42cf0de5, 32'h4403d746},
  {32'h448e8407, 32'h4376aafa, 32'hc36e5173},
  {32'hc38a730d, 32'hc31a912f, 32'h418610f4},
  {32'h44965fe2, 32'h4329f0d3, 32'h42e8cef9},
  {32'hc4ce2d7c, 32'hc32cc62a, 32'h43dbf374},
  {32'h44bced2b, 32'hc418ee60, 32'hc37c6b16},
  {32'hc4a2f1dc, 32'hc35ec8c8, 32'h43f6f0fc},
  {32'h4470c368, 32'h4347a243, 32'hc3d669b5},
  {32'hc4fc9534, 32'hc2355c04, 32'h431c7535},
  {32'hc1522600, 32'h4305f846, 32'h42b1aead},
  {32'hc41ee2ef, 32'h42c52733, 32'hc2899d66},
  {32'h44bf533c, 32'hc412a786, 32'hc3c764a4},
  {32'hc338b378, 32'h4350277c, 32'h43977a79},
  {32'h44b3a4f3, 32'hc29a4262, 32'h4305dc50},
  {32'hc272b890, 32'hc33cd97a, 32'hc36043f5},
  {32'hc38bf379, 32'h42fce6c5, 32'h42d35e6f},
  {32'h4470220e, 32'h435ce6bb, 32'h43955475},
  {32'hc4859085, 32'h43ad3ccb, 32'hc03662ff},
  {32'h44c2f881, 32'hc37da43e, 32'h42e924a8},
  {32'hc4d2deed, 32'hc282494d, 32'h43283ca6},
  {32'h429d1d88, 32'hc3bc5d2c, 32'hc38feedb},
  {32'hc4bd8b7b, 32'hc2b5281a, 32'hc3bb8bc3},
  {32'h44f021f8, 32'h4319e570, 32'hc2bb42ae},
  {32'hc4b45ac5, 32'h43c9ca8b, 32'h42a13838},
  {32'h440cbe86, 32'h42cc6361, 32'hc285b441},
  {32'hc50bb922, 32'h41ecc126, 32'h41ebdfde},
  {32'h450f3fe9, 32'hc34a3e89, 32'hc2c930f1},
  {32'hc20b5760, 32'h4379b983, 32'h430f7d48},
  {32'h447d6aa5, 32'hc1cece63, 32'hc362e326},
  {32'hc4ea1526, 32'hc2bb8cce, 32'h4411d86e},
  {32'h429d9e24, 32'hc2f8f67f, 32'hc3107f34},
  {32'h43747ab0, 32'h426ae608, 32'hc2653a42},
  {32'h44da3efa, 32'h43633998, 32'hc2e960d3},
  {32'hc4e2d204, 32'hc243b57f, 32'h4372d001},
  {32'h44ab376d, 32'h430460a4, 32'hc38b3d3e},
  {32'hc4d2143c, 32'hc1fd284c, 32'h4006a2f0},
  {32'h444d26ae, 32'h4236765f, 32'hc3b2c2ee},
  {32'hc4f825b8, 32'h4191cb36, 32'h431611fa},
  {32'hc0895080, 32'hc3bddfab, 32'hc3203e98},
  {32'hc503bfc0, 32'h43ac1e62, 32'h429d26fd},
  {32'h44550d8a, 32'hc343156d, 32'hc12ddc62},
  {32'hc22bc000, 32'hc2ef72c0, 32'hc2cb19b8},
  {32'h44c34735, 32'h43087bb1, 32'hc32b3f6d},
  {32'hc4abc37a, 32'h427610cc, 32'h439f048b},
  {32'h446130cc, 32'h439c4fc0, 32'hc399d1df},
  {32'hc313cad0, 32'hc390f55b, 32'h4284ba58},
  {32'h44153aa8, 32'h43e48ea3, 32'h42ee66df},
  {32'hc502a55e, 32'h40f54a38, 32'hc34ba900},
  {32'h44f2fe77, 32'h42d40d2b, 32'hc39b7426},
  {32'hc471a9a4, 32'h43845fd0, 32'h435cfafc},
  {32'h448eaaa1, 32'hc35f6f59, 32'hc3760bcb},
  {32'hc3904b3b, 32'h42c2204e, 32'h42c63205},
  {32'h44a4c0ca, 32'hc20badaf, 32'h43b4a7e7},
  {32'hc32b3c9e, 32'hc34c2bdf, 32'hc41d104d},
  {32'h44b7edd2, 32'h42aeebeb, 32'h438a30b5},
  {32'hc510af94, 32'h429a367e, 32'hc3321c5a},
  {32'h4370c040, 32'hc38249fd, 32'h42330c54},
  {32'hc4665093, 32'hc3cf29e7, 32'h40a65bf6},
  {32'h44df8892, 32'hc3456c3f, 32'h429aec8f},
  {32'hc532eb5f, 32'hc3a725bf, 32'h4286d0fe},
  {32'h44c5e1e3, 32'hc3bf328e, 32'h4383bd3e},
  {32'hc3a7c5d2, 32'h42bed0c7, 32'h43c3f6c2},
  {32'h44a49708, 32'h438e39ba, 32'h434d9fd4},
  {32'hc4e178b9, 32'hc32c34a0, 32'h42d7e390},
  {32'h440ced18, 32'h429a2686, 32'h4343d7a8},
  {32'hc4ca3a7d, 32'hc3ca5be7, 32'h41426e18},
  {32'h450f4843, 32'hc2c71cc3, 32'h433b7f60},
  {32'hc430d984, 32'hc362ccfc, 32'h4364ef72},
  {32'h4384527d, 32'h41e61492, 32'hc245fefb},
  {32'hc47f9169, 32'h438d8ad2, 32'hc33cda83},
  {32'h44a06497, 32'h4342956a, 32'h42800d31},
  {32'hc503c201, 32'hc3814e2b, 32'hc41619c7},
  {32'h44837546, 32'hc3918480, 32'hc3465fb1},
  {32'hc48128ea, 32'h4287292b, 32'h43a11c66},
  {32'h4428ec48, 32'hc3634146, 32'hc30abdde},
  {32'hc378eeb0, 32'hc24c4ef8, 32'h4347cd55},
  {32'h44b63828, 32'h4263b370, 32'h43199c41},
  {32'hc508e8f2, 32'h4342b616, 32'hc2f0c0c2},
  {32'h42aa66c4, 32'h418d36e2, 32'h436b36bd},
  {32'hc390b385, 32'h430c073e, 32'h43249bd1},
  {32'h44841b15, 32'h43453f1f, 32'hc3e19a10},
  {32'hc4acd217, 32'hc212f07e, 32'h42fd8736},
  {32'h445312af, 32'hc33af72a, 32'hc3379a42},
  {32'hc50473a8, 32'hc301b2de, 32'h43b2b9ff},
  {32'h450f329c, 32'h41f96665, 32'h4069cdc1},
  {32'hc4474010, 32'hc3604eec, 32'h42b29ebc},
  {32'h445cc336, 32'hc4041f17, 32'hc3a13898},
  {32'hc434900f, 32'h42084819, 32'hc2b90fa5},
  {32'h4515a065, 32'h4353b98f, 32'hc2243e32},
  {32'hc3c2a198, 32'h439184e2, 32'hc30dbf0d},
  {32'h443728a8, 32'h42d49f5b, 32'h435add1c},
  {32'hc4c03374, 32'hc28df45e, 32'hc364ee8e},
  {32'h4436eab7, 32'hc39f350d, 32'hc1b4fbf7},
  {32'hc4cdcac5, 32'hc33b3bba, 32'h42ee4ce8},
  {32'h449f997e, 32'hc38daaf8, 32'h4390fa4d},
  {32'hc22aeec0, 32'h43cbfa5a, 32'hc38a229c},
  {32'h43e59b83, 32'h430f54ed, 32'hc1c51598},
  {32'hc4ede363, 32'hc2a9759a, 32'h436fb1e8},
  {32'h438c05c0, 32'hc287c12b, 32'h4402620e},
  {32'hc4ce6842, 32'hc2910068, 32'h427aa760},
  {32'h44644d32, 32'h432233b0, 32'h417324fc},
  {32'hc5185c1b, 32'hc284818b, 32'h424ce2de},
  {32'h4490a384, 32'h42872b90, 32'h4395de00},
  {32'hc4a29a4a, 32'hc3d0e8f6, 32'h43623284},
  {32'h44e3eeba, 32'hc3025cce, 32'hc0e75f20},
  {32'hc3520e78, 32'h435f6015, 32'h43094c98},
  {32'h44e82dfd, 32'h43a96a81, 32'h438383c1},
  {32'hc4ae41d9, 32'hc30d679a, 32'hc2d5aecc},
  {32'h4502aa7f, 32'h425c3feb, 32'hc3214144},
  {32'hc3ffe298, 32'hc385ac6a, 32'hc1cbb4eb},
  {32'h440a8688, 32'h4388ed1c, 32'h435e4455},
  {32'hc26e5640, 32'h43a84d55, 32'hc22e0516},
  {32'h42ae6a40, 32'hc34af859, 32'hc31ae357},
  {32'hc4967ab4, 32'hc29d4813, 32'h43718520},
  {32'h4434a5ca, 32'h43a5fc70, 32'hc2a2ffdf},
  {32'hc4994e94, 32'h43750462, 32'hc2bdc4ae},
  {32'h4426ffdc, 32'hc1ef7819, 32'h437313de},
  {32'hc4957716, 32'hc3908d3e, 32'hc3efbd55},
  {32'h4505ae49, 32'h420466c6, 32'h41513049},
  {32'hc5107cbb, 32'h42b64768, 32'hc10541eb},
  {32'h44328cf6, 32'hc3007d90, 32'hc3f45152},
  {32'hc3f79230, 32'hc2082caa, 32'hc28157cf},
  {32'h44a7a84d, 32'hc20cb3c3, 32'hc2d65ff0},
  {32'hc4d00de8, 32'hc2f1987d, 32'hc280b066},
  {32'h4495a2e1, 32'hc31951c5, 32'h42926d70},
  {32'hc4f11f11, 32'hc3c2bc45, 32'hc1c08c64},
  {32'h4485edd0, 32'hc3b65b71, 32'hc2bbf3a6},
  {32'hc49f0b69, 32'hc2be1668, 32'h43872d8f},
  {32'h44929291, 32'h42a08722, 32'h43ca8bcb},
  {32'hc49b82b3, 32'h43720672, 32'hc15f7e8c},
  {32'h4499cf64, 32'h43b7f308, 32'h42d5eb2a},
  {32'hc4d5b70d, 32'h43fab5de, 32'h435bad28},
  {32'h45062038, 32'hc14dfc9b, 32'h41e30d68},
  {32'hc437db68, 32'hc3c90687, 32'hc2b693bc},
  {32'h4514dadb, 32'hc2b0d960, 32'hc3ae5b6d},
  {32'hc4851435, 32'h422a1365, 32'h43e666e1},
  {32'h45076b03, 32'hc3ba31dd, 32'h418f85d4},
  {32'hc4c923da, 32'hc34cb7a6, 32'hc343e658},
  {32'h4418db42, 32'hc341034f, 32'h435b87d3},
  {32'hc389c982, 32'h434e62d2, 32'hc34dde34},
  {32'h44275104, 32'hc0df896b, 32'h43556b56},
  {32'hc36ae72c, 32'h42b443a5, 32'hc2d225ce},
  {32'h45111bbf, 32'h428ff20a, 32'hc2907cf0},
  {32'hc48c6d31, 32'hc2dd4869, 32'h4399e558},
  {32'h450b70b4, 32'h437eb51a, 32'hc17f236a},
  {32'hc43668d1, 32'hc3ab0a22, 32'h41a6d73c},
  {32'h44821aa7, 32'h43db396d, 32'hc3842393},
  {32'hc4d8d053, 32'h4392fbdf, 32'h432fdfed},
  {32'h44d8f8d6, 32'h43563964, 32'h4339e2f3},
  {32'hc3e610f8, 32'hc25f09f2, 32'hc290906a},
  {32'h444186c3, 32'h42c5e41e, 32'hc2a6cca9},
  {32'hc37007f0, 32'h43e53306, 32'hc375a2da},
  {32'h44d8842f, 32'hc3b5ffaa, 32'h426173c6},
  {32'hc44323fb, 32'hc302a120, 32'hc3aef691},
  {32'h44f1c35e, 32'hc2277927, 32'h4109793e},
  {32'hc5031751, 32'h426b294d, 32'hc36abdbc},
  {32'h44e6c1bf, 32'hc363faa4, 32'hc382f81f},
  {32'hc4d1cdd7, 32'h43c3b151, 32'h42721bae},
  {32'h4309fc62, 32'hc3970669, 32'h44114718},
  {32'hc4169fd8, 32'h42e8dd9d, 32'h4374fc00},
  {32'h44e0aca1, 32'hc39ab859, 32'hc338d774},
  {32'hc4f10c09, 32'h40aecd98, 32'h43193a39},
  {32'h450b7490, 32'hc39756d4, 32'h43abcb4c},
  {32'hc457f4e9, 32'hc35861f8, 32'hc323f897},
  {32'h4501397b, 32'hc304da74, 32'h421e011b},
  {32'hc36346d0, 32'h42d28780, 32'h434d0cd0},
  {32'h43b38ed7, 32'hc23107b0, 32'hc3370904},
  {32'hc3931858, 32'h4371c333, 32'h4335164a},
  {32'h4489282f, 32'h43bae111, 32'hc3aa68e7},
  {32'hc48b78b6, 32'h43625dfe, 32'h433ce567},
  {32'h44051846, 32'hc30707b1, 32'hc38ef75b},
  {32'hc4821cae, 32'hc33f5120, 32'hc354348d},
  {32'h44e9d9a2, 32'hc2afa2b2, 32'hc3b2a822},
  {32'hc4700a64, 32'hc403c6a5, 32'h43dbb3a0},
  {32'h44d6a98c, 32'h41ce93c4, 32'h4303dd2b},
  {32'hc4fb6ee9, 32'hc301a9c4, 32'h42eca851},
  {32'h44a8f16e, 32'hc2312df1, 32'hc270e03c},
  {32'hc5186c12, 32'hc2178b14, 32'h42b18ac6},
  {32'h43cca24c, 32'hc314d536, 32'hc39f7b6a},
  {32'hc506f2c8, 32'hc3378e52, 32'h43a4fdba},
  {32'h4510c6f2, 32'hc1aee938, 32'h4288088e},
  {32'hc4d8b176, 32'hc3a53ad6, 32'h4350c0b3},
  {32'h443db867, 32'h43e838df, 32'hc3cf80f5},
  {32'hc4b1600e, 32'hc332acbd, 32'hc35d69a0},
  {32'h442fe2e8, 32'h433aca42, 32'hc33c5028},
  {32'hc4e3ced2, 32'hc3793a98, 32'hc3484783},
  {32'h43f3fa04, 32'h418e7c5a, 32'h42d354de},
  {32'hc397785c, 32'hc3095bca, 32'hc16f7910},
  {32'h44b09598, 32'hc2bca074, 32'hc128d0f2},
  {32'hc4ef98a8, 32'hc306d025, 32'hc386cded},
  {32'h4507347d, 32'h43a60bee, 32'hc1fd2073},
  {32'hc4f8932e, 32'h4353b06f, 32'h43076b8e},
  {32'h441d540d, 32'h4293de9c, 32'h42f2194e},
  {32'hc2dbcdc0, 32'h43b0eb64, 32'hc3aa98ea},
  {32'h435fb589, 32'hc3baf439, 32'h428dec5b},
  {32'hc4cd4e5d, 32'hc325e021, 32'hc23d4323},
  {32'h44b58e15, 32'h4395e6ba, 32'h43885560},
  {32'h4314fcd0, 32'hc2b7b7b6, 32'h4175df38},
  {32'h446e1cb2, 32'hc397cf85, 32'h43289218},
  {32'hc5186fbc, 32'hc1ff13fa, 32'h41b5376f},
  {32'h44ca790b, 32'h4333d4f9, 32'hc3ac5eef},
  {32'hc2c01820, 32'h4368c598, 32'h431109ab},
  {32'h44556410, 32'hc2e58da6, 32'hc2e1144c},
  {32'hc5173a35, 32'hc3a212fd, 32'h43721f1a},
  {32'h450de77d, 32'h43756468, 32'h438fcaf0},
  {32'hc404df2e, 32'hc3dc69e3, 32'h4222be0f},
  {32'h44d67542, 32'h43626a2e, 32'h429987d6},
  {32'hc4d67a3b, 32'h430ad63b, 32'hc314dd79},
  {32'h44c93464, 32'h43bf9a47, 32'h4228af65},
  {32'hc45abc96, 32'h43a6fb13, 32'h42d1218b},
  {32'h44b40200, 32'hc287537a, 32'hc182cfae},
  {32'hc33cb6f9, 32'hc3968301, 32'h418c5c73},
  {32'h440fcbbd, 32'hc2facc5d, 32'h42324a69},
  {32'hc5038b38, 32'hc31a4772, 32'hc2c52aee},
  {32'h4476a909, 32'h4200b3c3, 32'h4383f57c},
  {32'hc49ae866, 32'hc3a496af, 32'h4330149f},
  {32'h44cec58a, 32'hc2d32085, 32'h4336ba17},
  {32'hc512619a, 32'h43071010, 32'h429dae8a},
  {32'h44e16acd, 32'h43d20f25, 32'h42e95700},
  {32'hc4a29a17, 32'h43e89a1b, 32'h42e0544f},
  {32'h44bab995, 32'hc2d4d7fe, 32'h438e1598},
  {32'hc4e395f4, 32'h4382239b, 32'hc24b3902},
  {32'h4485662f, 32'hc387e0c1, 32'hc3704a53},
  {32'hc4cd5c60, 32'h420b3a74, 32'hc3e16a86},
  {32'h44282ad4, 32'hc152d4ba, 32'h438b1264},
  {32'hc439d85e, 32'h42de2d98, 32'hc2b2cd06},
  {32'h42ec9d20, 32'h438ad339, 32'hc3d9a5ea},
  {32'hc392a6ba, 32'hc3a23e58, 32'hc2c0c3aa},
  {32'h44ccbec9, 32'h4395c02e, 32'hc28fff2b},
  {32'hc4a5592a, 32'h42845af8, 32'hc2d166a4},
  {32'h4483a06d, 32'hc2ff095a, 32'hc1fdd43b},
  {32'hc4238a56, 32'h438e55e2, 32'h41ffe14c},
  {32'h44e67a30, 32'hc2f42618, 32'h42de41d4},
  {32'hc48b03e0, 32'hc3511d4b, 32'h43c2cb15},
  {32'h44a56b3e, 32'hc3757189, 32'hc343eff5},
  {32'hc42cbb9e, 32'h4327dcfe, 32'h427b35d2},
  {32'h44b480ec, 32'h42cd409d, 32'hc3c83182},
  {32'hc38801ba, 32'h42ed027b, 32'hc202ba0b},
  {32'h44bf8bd8, 32'h43262821, 32'h42cf9f87},
  {32'hc4abba70, 32'h4331f7d3, 32'hc286f1eb},
  {32'h44c073dd, 32'h432b7260, 32'h43c5b2f3},
  {32'hc50bd175, 32'hc1828b0f, 32'h41b356da},
  {32'h45032a04, 32'hc349b10a, 32'hc3a4a760},
  {32'hc4ec4fc6, 32'hc1027338, 32'h42200c12},
  {32'h44e2d9f0, 32'h43673b6f, 32'hc39190c0},
  {32'hc334af70, 32'h43811640, 32'hc20312dc},
  {32'h44c52a52, 32'h43a44bfe, 32'hc2d0ab2e},
  {32'hc4e3715a, 32'hc32647da, 32'h42e58f22},
  {32'h44075948, 32'h424471ee, 32'hc39b86b7},
  {32'hc4824a8e, 32'hc26c3aeb, 32'h43b9b59e},
  {32'h4414949a, 32'h429dee16, 32'hc3b3b482},
  {32'hc4c8f518, 32'hc3568180, 32'h43e06eca},
  {32'h44ac0a0c, 32'hc30d8948, 32'hc1092bc6},
  {32'hc3fc7bb7, 32'hc36e7d23, 32'h43bc8a2e},
  {32'h44682196, 32'hc29cb076, 32'hc38cc510},
  {32'hc42f8c04, 32'hc2ed0db7, 32'hc20cd8f5},
  {32'h44e090d6, 32'hc41a1a36, 32'hc35386d9},
  {32'hc4d734b7, 32'hc35be79e, 32'h432c5726},
  {32'h44cac1ae, 32'hc2d4af75, 32'h436af278},
  {32'hc50c7fa8, 32'hc150003c, 32'h435dea96},
  {32'h41282700, 32'h42a8bbf3, 32'hc3ca367c},
  {32'hc515ce90, 32'hc3a20da5, 32'h43441109},
  {32'h45139201, 32'h43b9dcbb, 32'hc3c29268},
  {32'hc46e4e10, 32'h427b68dc, 32'hc1a5ce99},
  {32'h4425df84, 32'h43007701, 32'hc2ca0f30},
  {32'hc468b677, 32'h439788e4, 32'hc20d8c2c},
  {32'h44695c00, 32'hc2735e74, 32'hc2b80cae},
  {32'hc4bb409a, 32'h4357b503, 32'h4269d794},
  {32'h44ca5adb, 32'h43f31d9d, 32'hc3546c0c},
  {32'hc48d019e, 32'hc35f9f9c, 32'hc216b167},
  {32'h442ba290, 32'hc3a7a797, 32'hc291599f},
  {32'hc507bf60, 32'hc28afb2b, 32'h430f65b4},
  {32'h44b7a8fe, 32'h43052d9e, 32'hc31260b8},
  {32'h4339b9cd, 32'h422f6dc5, 32'hc2a05ac9},
  {32'h4401d1d8, 32'h435e0602, 32'hc25fbb11},
  {32'hc4a7131a, 32'hc33a42d6, 32'h42ac4c39},
  {32'h44b7f0dc, 32'h429d5018, 32'h431cdca6},
  {32'hc4f3bc94, 32'hc3c6395a, 32'hc2abd834},
  {32'h44a9ca8c, 32'h42189f72, 32'hc2284d75},
  {32'hc500dcb8, 32'h42a57b0d, 32'h438b417c},
  {32'h44a0f594, 32'h42ba3c45, 32'hc29ef0d6},
  {32'hc4e78e5b, 32'hc18a2f79, 32'h429af494},
  {32'h44f965d0, 32'hc269e642, 32'h430665da},
  {32'hc4f9d22e, 32'hc33df507, 32'hc23cb15e},
  {32'h43f58b82, 32'h4388ae4e, 32'h432b16cd},
  {32'hc42da4ce, 32'h42c30570, 32'h429091d0},
  {32'h44fd33e1, 32'hc3c84072, 32'hc3eb1c5b},
  {32'hc5111af6, 32'hc39f3baf, 32'h42c08105},
  {32'h447f77f4, 32'hc30e1857, 32'hc41e9d97},
  {32'hc3e465e4, 32'hc3cee063, 32'hc2ac1607},
  {32'h44fc3930, 32'hc2d47e43, 32'hc112c3b7},
  {32'hc4d09b96, 32'h43449b81, 32'hc2c80f6a},
  {32'h44d9bbcb, 32'h4381451d, 32'hc30c89cb},
  {32'hc4f2d3bf, 32'h425bdb02, 32'h420f90f8},
  {32'h444eeec9, 32'h41a4cb1a, 32'h4256ae6e},
  {32'hc3d75eee, 32'h41ed1c8d, 32'h4212299b},
  {32'h44e0ba95, 32'hc301b932, 32'hc2473c33},
  {32'hc4b21dae, 32'h4314a139, 32'hc2c774bf},
  {32'h45011a4f, 32'hc30a3bcb, 32'h42c93971},
  {32'hc4dd1d60, 32'h4378b563, 32'h43b11316},
  {32'h447726e1, 32'hc310ad1a, 32'h4389b0b8},
  {32'hc4fcea44, 32'h42ac5050, 32'hc2d69f9e},
  {32'h4506c374, 32'h42acead2, 32'hc33ae3cf},
  {32'hc440856b, 32'h431613d2, 32'h4291a65e},
  {32'h4471d3d9, 32'hc395e917, 32'hc391c428},
  {32'h428e7dc0, 32'h4165c3dc, 32'h43f63cce},
  {32'h437f7500, 32'h42f3417a, 32'h4256c0ba},
  {32'hc31bafb0, 32'hc246ab8c, 32'hbfc3fee0},
  {32'h44e199f9, 32'h428abba2, 32'hc21bbac4},
  {32'hc4ebb92d, 32'hc402bef6, 32'h42fb52e7},
  {32'h448aeef2, 32'h43ced95d, 32'h423450eb},
  {32'hc4e683ad, 32'h431936dc, 32'h43b4d1c4},
  {32'h4457b08a, 32'h423b489b, 32'h437dbd0c},
  {32'hc4a96734, 32'hc33f21ec, 32'hc2eb9dd0},
  {32'h451e191b, 32'hc312f550, 32'hc2c94309},
  {32'hc41e0178, 32'h42f7ba9e, 32'h426c2144},
  {32'h44bce988, 32'h41da2039, 32'h4355b703},
  {32'hc45c51c6, 32'h42bc9690, 32'hc2b1106e},
  {32'h45090d18, 32'hc387dbb4, 32'hc399a659},
  {32'hc3bf6038, 32'hc30811e2, 32'hc2b9de9d},
  {32'h44b954fa, 32'h42bd84f9, 32'hc25fbb33},
  {32'hc48b5c80, 32'hc18b9bda, 32'hc2fec01a},
  {32'h4500f0ed, 32'h431daf18, 32'hc29969c0},
  {32'hc35c0710, 32'h410806e6, 32'hc233b372},
  {32'h441847e4, 32'hc343365d, 32'h42c1aada},
  {32'hc342e5a0, 32'h432ca512, 32'h42807904},
  {32'h44772904, 32'hc32b3800, 32'h433203cf},
  {32'hc502468f, 32'hc217a611, 32'hc3341ec5},
  {32'h446a3bd2, 32'h4252519a, 32'hc313cd8b},
  {32'hc3ca377b, 32'hc31ac4db, 32'h432e28cf},
  {32'h4484ec31, 32'hc39f8d52, 32'hc226dc55},
  {32'hc407a684, 32'hc22a7d91, 32'h4396fc82},
  {32'h442fc922, 32'h431419a1, 32'hc407bfa4},
  {32'hc491c5ad, 32'h42418f70, 32'hc2319cbb},
  {32'h44d1ccba, 32'h4348dbb3, 32'h4380adad},
  {32'hc510e350, 32'h434a8f98, 32'h41fa5038},
  {32'h44792298, 32'hc2c09645, 32'h428274c7},
  {32'hc42ddfcc, 32'h438c91b6, 32'h439b68fc},
  {32'h4105b400, 32'hc3491eab, 32'hc2f2c34f},
  {32'hc4a84879, 32'h4336953e, 32'h4298cc2a},
  {32'h450463a7, 32'hc38aa7dc, 32'hc34edacf},
  {32'hc503d847, 32'h428fa172, 32'h42c4c5c1},
  {32'h43278e08, 32'hc35804f8, 32'hc34594b5},
  {32'hc351aa66, 32'h421add55, 32'h435421db},
  {32'h451125fb, 32'h440a9bcd, 32'h43c4bf3b},
  {32'hc4093576, 32'h43b63258, 32'hc325d5f8},
  {32'h431d0fb0, 32'hc420eb56, 32'hc3183ae2},
  {32'hc50504f7, 32'h41bc9bcd, 32'hc3e57f79},
  {32'h44ab2f66, 32'hc39a38a3, 32'h4343185c},
  {32'hc47bd727, 32'hc2fbff86, 32'hc3153ead},
  {32'h443a420e, 32'h3fe76ee5, 32'hc2f9a4f7},
  {32'hc2af5cc0, 32'hc30b1c35, 32'h43945464},
  {32'h44bae2dc, 32'h42f36172, 32'hc31b82ab},
  {32'hc3a44910, 32'hc3b18b08, 32'hc386c122},
  {32'h438ae960, 32'hc28f365e, 32'h43dc06eb},
  {32'hc51445de, 32'h43406579, 32'h42937dad},
  {32'h4437633a, 32'h4394233c, 32'h42db693c},
  {32'hc4b7867f, 32'hc18aa9b7, 32'h4190a91a},
  {32'h4519216f, 32'h436f1b40, 32'hc3b7aa64},
  {32'hc4ae7823, 32'h435c173f, 32'hc34a9d1d},
  {32'h4483d64b, 32'hc2a9464c, 32'hc25a12b5},
  {32'hc4b2d13d, 32'h433f2b47, 32'h420924f6},
  {32'h44d0ebfc, 32'hc1cf8e6c, 32'hc38d82ae},
  {32'hc3e7adf8, 32'hc380044e, 32'h438d9809},
  {32'h42ef57c8, 32'hc3c77182, 32'hc30528b6},
  {32'hc50249d9, 32'hc3738272, 32'h439b7e45},
  {32'h43a37c00, 32'hc1ebbc79, 32'hc38f348f},
  {32'hc442b96c, 32'hc2454361, 32'h42eaa7e2},
  {32'h4523374e, 32'hc43cf018, 32'h425e88b0},
  {32'hc3ced02a, 32'hc3330f67, 32'h41c8138c},
  {32'h44d87fdf, 32'hc3b58d23, 32'h423bd860},
  {32'hc2f7345c, 32'hc39a4663, 32'h43830d5a},
  {32'h44f6ce26, 32'hc30a6db0, 32'hc2fdae72},
  {32'hc4edb318, 32'h43a499a4, 32'hc37d9e56},
  {32'h450cb197, 32'h435f7a2f, 32'h438b789c},
  {32'hc48aa938, 32'hc2fa7a35, 32'h4119207a},
  {32'h44b463fb, 32'h43918125, 32'h4290010e},
  {32'hc4dc684c, 32'h436d1a56, 32'hc263d5ce},
  {32'h44d17651, 32'hc350ce60, 32'hc2de8614},
  {32'hc4e5549e, 32'h430b4f12, 32'hc21ffce3},
  {32'h44902286, 32'h43a4a9ba, 32'h43106074},
  {32'hc51a0716, 32'h435a70c3, 32'hc3875441},
  {32'h44853d23, 32'hc1afbd41, 32'h411b4633},
  {32'hc4c3ca7c, 32'hc28513c6, 32'h43887a63},
  {32'h43f8cd25, 32'h4386b612, 32'hc383d436},
  {32'hc4c18f06, 32'hc2ff463e, 32'h41914898},
  {32'h447378fe, 32'h3f25f1b0, 32'hc0de8ee8},
  {32'hc430c6a6, 32'h4257c368, 32'h43f66174},
  {32'h450729b4, 32'h4341cd30, 32'h439ddada},
  {32'hc44ae640, 32'h40dda464, 32'hc3329f3a},
  {32'h44c0cc34, 32'hc2ffa9ed, 32'hc37d8900},
  {32'hc4434304, 32'hc29e731d, 32'h43d054f1},
  {32'h44f135f9, 32'h43937291, 32'h4306d772},
  {32'hc4dbcfb1, 32'hc24a58e5, 32'hc322175c},
  {32'h44f08da3, 32'h43dc25ae, 32'h42063a1a},
  {32'hc3a9e7a0, 32'hc35e4483, 32'hc332d5e7},
  {32'h44cf0496, 32'h42ea8269, 32'hc12549f0},
  {32'hc3a0245a, 32'h4350142e, 32'hc11f75a7},
  {32'h446a64d9, 32'hc31dd9fb, 32'h41ad9c28},
  {32'hc3821592, 32'h43b05a06, 32'hc3e1c8f5},
  {32'h44c1bae7, 32'hc2603e90, 32'hc2364f9b},
  {32'hc4160f85, 32'h41c7c1be, 32'hc3af0609},
  {32'h45053b3c, 32'hc3217097, 32'hc392b46e},
  {32'hc3aa0834, 32'hc35878f5, 32'hc29763f0},
  {32'h44261d38, 32'h43be996b, 32'h42e6e523},
  {32'hc4fb9513, 32'h42261c13, 32'h4358c8e3},
  {32'h44b53834, 32'h42a5028c, 32'hc2f93549},
  {32'hc505eb89, 32'hc339ce9a, 32'h4342e9d8},
  {32'h42c779e0, 32'h42e2efb0, 32'hc2cbfa10},
  {32'hc3a84fe6, 32'hc387b99c, 32'hc22be14d},
  {32'h44a4634c, 32'h4271bc72, 32'h429595b4},
  {32'hc44f7c1c, 32'h4360d875, 32'hc274bacf},
  {32'h4504c64c, 32'hc2a43b50, 32'hc3aeda1f},
  {32'hc4c28443, 32'hc2bdc4e8, 32'h42867cb8},
  {32'h44b2e193, 32'hc360117b, 32'h43b47986},
  {32'hc4e3e564, 32'h43d44270, 32'hc401c130},
  {32'h450548a4, 32'h43f82d85, 32'hc2b1013f},
  {32'hc4e8f5b1, 32'hc2dab919, 32'h441a78cd},
  {32'h450600c0, 32'h41a2964f, 32'hc383b6b8},
  {32'hc429f382, 32'h429be662, 32'hc3c39c34},
  {32'h4483a066, 32'h43a9745f, 32'hc2eabcce},
  {32'hc3ce9578, 32'hc3c59e6c, 32'h4135bf06},
  {32'h43c4e418, 32'hc30e79de, 32'h42b6adc4},
  {32'hc456a603, 32'hc314ffea, 32'hc2ba854e},
  {32'h44fab6b2, 32'h425b62b7, 32'hc39ea470},
  {32'hc4b9ca67, 32'hc204defe, 32'hc33cd3c8},
  {32'h4452a3d1, 32'h4377b830, 32'hc0beaad8},
  {32'h420a4b02, 32'h437b30c9, 32'hc240cb0a},
  {32'h42f44cd0, 32'h436416b3, 32'h4200a78d},
  {32'hc3445fb2, 32'h43713126, 32'hc3875d26},
  {32'h44b9f6d5, 32'hc2bc520d, 32'h4411d173},
  {32'hc334d32c, 32'h435a1d40, 32'h4174c5ec},
  {32'h44f2662a, 32'h439a728a, 32'hc36eb876},
  {32'hc4f86e63, 32'hc2367ea3, 32'hc3560249},
  {32'h450be65b, 32'hc2e78bc5, 32'hc336e267},
  {32'hc4d644c4, 32'h413c9d3a, 32'h41d4c8fc},
  {32'h444616fa, 32'hc1eee97d, 32'hc1dd0360},
  {32'hc4460eec, 32'hc18e44f6, 32'hc40698cb},
  {32'h45034268, 32'hc3087986, 32'hc25812ef},
  {32'hc4481d6f, 32'h42aa1a77, 32'h406f6e0b},
  {32'h4474c838, 32'hc304944f, 32'h4402a36e},
  {32'hc3feb50b, 32'hc3c078b9, 32'hc3ed3850},
  {32'h45172622, 32'h41cbe14d, 32'hc32da402},
  {32'hc4317993, 32'hc38ca08b, 32'hc3f83e4a},
  {32'h4496aefc, 32'h43a5b0e4, 32'h44293f0b},
  {32'hc4b76936, 32'hc32ea098, 32'h42f1c607},
  {32'hc4ab15f9, 32'hc303635c, 32'h4310e952},
  {32'h4492809d, 32'h431858db, 32'hc2b24755},
  {32'hc4ca718f, 32'h42560304, 32'hc426d830},
  {32'h43b1d2fd, 32'hc323dd52, 32'h43f2a2d7},
  {32'hc49c1ec2, 32'hc32e2681, 32'hc114f6a8},
  {32'h451090d9, 32'h43804012, 32'hc36f454f},
  {32'hc34baa18, 32'h42de49be, 32'hc34a8744},
  {32'h44a0ad81, 32'hc354e27b, 32'h422186c8},
  {32'hc4a2b8f7, 32'h434b74dd, 32'hc30a11d6},
  {32'h43d3fe60, 32'hc2c2204c, 32'hc3694ea7},
  {32'hc4c0c82e, 32'h429a4193, 32'h420b058e},
  {32'h43e97226, 32'hc3cab56d, 32'h43f38cda},
  {32'hc3665880, 32'h43e7b0c5, 32'hc1d6238c},
  {32'h451718db, 32'h43495e1c, 32'h43a95b9c},
  {32'hc1c78810, 32'h4235e10a, 32'h426d23c9},
  {32'h44956196, 32'hc22c36f0, 32'h428928b7},
  {32'hc504d928, 32'hc274bb29, 32'h41000307},
  {32'h431d85d2, 32'h439e8eec, 32'hc28fa5d8},
  {32'hc147a800, 32'hc3bae181, 32'hc37abc06},
  {32'h446ad42c, 32'hc157b297, 32'hc135fd4d},
  {32'hc3cbc37a, 32'h431a10b9, 32'hc3fc1a8f},
  {32'h4436f43c, 32'h43909468, 32'hc3940aca},
  {32'hc4146659, 32'hc3e48295, 32'hc3772179},
  {32'h431fc94e, 32'hc2bea32b, 32'h430876ad},
  {32'hc4527288, 32'h435412a7, 32'hc3486426},
  {32'h450b4379, 32'h42d3893a, 32'hc2df1ea1},
  {32'hc40d8bac, 32'hc33f11ff, 32'hc33f5d59},
  {32'h44cdf4ee, 32'h42a4ea83, 32'h4207cf30},
  {32'hc48fac22, 32'h435a6443, 32'hc45750bf},
  {32'h44a201f4, 32'hc2493fc7, 32'h4394e094},
  {32'hc3a5a888, 32'hc2bc9c91, 32'hc38a4752},
  {32'h44d05248, 32'hc387d9ff, 32'hc17d9da4},
  {32'hc4bc3996, 32'hc3a41074, 32'h43cba9b7},
  {32'h44f4f9c3, 32'hc311d28d, 32'h4293f773},
  {32'hc4e6b7bc, 32'h41e995f3, 32'hc3713024},
  {32'h44decd76, 32'h42a3a510, 32'h4353babe},
  {32'hc503c8d2, 32'hc3647ec2, 32'hc38077f4},
  {32'h44e81c04, 32'h42d32930, 32'h434bc24e},
  {32'hc4a816c4, 32'h40a9e4fa, 32'h43dc75e7},
  {32'h4487d0d3, 32'h43979d63, 32'hc147b1af},
  {32'hc44d7acc, 32'h41dab0ee, 32'hc2c36f45},
  {32'h44783cf5, 32'h439e3099, 32'h42823c09},
  {32'hc4b8382e, 32'h424aa669, 32'hc2da7768},
  {32'hc2634ad0, 32'hc2c4f2ce, 32'h42efe3ae},
  {32'hc48e83fd, 32'hc312a805, 32'h426c0a06},
  {32'h4426abb8, 32'hc385c79a, 32'hc3a8ba11},
  {32'hc4f03b4e, 32'h43ec8266, 32'hc3d9a427},
  {32'h4521c07d, 32'h438c8d00, 32'hc2d83e5c},
  {32'hc4d484eb, 32'hc0760ed5, 32'h429ea75c},
  {32'hc334e2ac, 32'h4215484c, 32'h433a34a0},
  {32'hc4931e7d, 32'h41db27b7, 32'h439e7184},
  {32'h44dfd358, 32'h413b0d4c, 32'hc34b18af},
  {32'hc41bd8ca, 32'h3ec8fe60, 32'hc3c4b6b0},
  {32'h43f66eac, 32'h4335a7ec, 32'h43c35185},
  {32'hc50b4705, 32'h434b9726, 32'hc1790109},
  {32'h44d4ded3, 32'h4380e808, 32'hc36865da},
  {32'h4320baba, 32'h42cc4150, 32'h423cf719},
  {32'h441ec326, 32'hc253b4ce, 32'hc24daa92},
  {32'hc498875d, 32'hc32e0c69, 32'h42a350c2},
  {32'h44cd58fe, 32'h43f4b481, 32'hc2753d4c},
  {32'hc443f4b8, 32'hc316ec9a, 32'h423434c4},
  {32'h451e91fc, 32'hc20de090, 32'h432f13f5},
  {32'hc443e556, 32'h411768b8, 32'hc369f29b},
  {32'h447640c0, 32'hc22baa60, 32'h436d231d},
  {32'hc4dc6f10, 32'h42419f0c, 32'h4227ea4f},
  {32'h43c3be1a, 32'h42aa9026, 32'h4397b4b8},
  {32'hc44b911e, 32'h42b99dff, 32'hc2f4ce86},
  {32'h45000008, 32'h41deab96, 32'hc30d6f2f},
  {32'hc4993b55, 32'h41d6a528, 32'hc30ae70c},
  {32'h44a1dd78, 32'h42fbbc42, 32'hc3afa259},
  {32'hc43706d3, 32'h42dbc809, 32'h4368f1b2},
  {32'h44991e77, 32'hc2b3afed, 32'h43c7dca6},
  {32'h434529cd, 32'hc3dbca17, 32'h443998ea},
  {32'h439d10d6, 32'h4300639c, 32'h436cb9ba},
  {32'hc3fb28ce, 32'h41423d8d, 32'h43802279},
  {32'h44dc8011, 32'h42dca751, 32'hc2e0f8af},
  {32'hc4f10606, 32'h4303a06d, 32'h416fcd58},
  {32'h449bd728, 32'h43f8185e, 32'hc1f008ba},
  {32'hc4f054b8, 32'h43708214, 32'h42c1a9b6},
  {32'h4509ef37, 32'hc355a2b8, 32'h4435972a},
  {32'h43e384c8, 32'hc3d23fdd, 32'hc37dcb5b},
  {32'h44514df4, 32'h438405f1, 32'hc35c647f},
  {32'hc4974532, 32'h4281adc7, 32'hc3705db2},
  {32'hc22028e0, 32'h4174c060, 32'hc355b0ac},
  {32'hc501bf32, 32'hc3aeb2f8, 32'h43cd7d2e},
  {32'h4463cb3e, 32'hc18fb9ea, 32'h43915417},
  {32'hc4fab08a, 32'h430d6116, 32'h43df6c41},
  {32'h44d3b988, 32'hc26b91cc, 32'hc36ee4f3},
  {32'h436082c0, 32'h42dee1b5, 32'h42f09518},
  {32'h445f9a4e, 32'hc280e63b, 32'hc3dc3bc0},
  {32'hc48f69be, 32'h4320900a, 32'hc2bc2f8b},
  {32'h4500ae6c, 32'h3e6be880, 32'hc35eec96},
  {32'hc516af3f, 32'h43282036, 32'h43720271},
  {32'h44373f5e, 32'h43b6391d, 32'hc3027af8},
  {32'hc456cc2e, 32'h4403aa07, 32'h428bfeb2},
  {32'h44b40ebe, 32'hc3537022, 32'h41e73362},
  {32'hc2fa0040, 32'hc2b69357, 32'h43a08d30},
  {32'h42973f20, 32'h43201c88, 32'hc38828b3},
  {32'hc518ccfc, 32'hc2d09ce8, 32'hc2df935d},
  {32'h431f6f70, 32'hc0dd5407, 32'hc1014668},
  {32'hc3133808, 32'hc3a1215d, 32'hc28efb2f},
  {32'hc2cb225a, 32'h43632477, 32'hc2bf3cc5},
  {32'hc49541b8, 32'h420ee7a8, 32'hc2f925d5},
  {32'hc3cc8a54, 32'h437eec33, 32'h43cddb5b},
  {32'hc444e9a8, 32'hc274676b, 32'h4402ee67},
  {32'h44a3e954, 32'hc37befdc, 32'hc34ada36},
  {32'hc5047111, 32'h42c3d151, 32'hc0593037},
  {32'hc35b5018, 32'hc3ea8ff2, 32'h43425509},
  {32'hc4dcaaec, 32'h438752c2, 32'h43452f30},
  {32'h44f96b26, 32'hc12cf255, 32'hc3cf0c65},
  {32'hc4c7bf5d, 32'hc2d677f7, 32'hc39c7314},
  {32'h451cd328, 32'hc37c5dcb, 32'hc3e62bbb},
  {32'hc423121e, 32'hc3bcf2ea, 32'hc389048d},
  {32'h443f6d54, 32'h4338e792, 32'hc236550e},
  {32'hc330bd90, 32'h43c694d6, 32'h42e03ace},
  {32'hc401f3ad, 32'h4316713f, 32'hc2f27b9e},
  {32'hc4d5a0d0, 32'h43828d54, 32'h430d4503},
  {32'h44c84a8e, 32'hc37d95d1, 32'h426ef813},
  {32'hc46f0df9, 32'h40eea37e, 32'h43ac6453},
  {32'h44a9daa8, 32'h426da5a2, 32'h438f3905},
  {32'hc40371ba, 32'hc31f23f3, 32'hc38b388d},
  {32'h44d24d84, 32'hc38396bd, 32'hc3a19434},
  {32'hc51268fb, 32'h42a0f9a8, 32'h410fe05a},
  {32'h44956392, 32'h430aaeff, 32'hc39466d5},
  {32'hc28610b8, 32'h43dc99ca, 32'h434c8529},
  {32'h43e7a810, 32'hc334843f, 32'h41e9cc72},
  {32'hc4498624, 32'hc2e72fbd, 32'h433d130f},
  {32'h445a8bc1, 32'h43e756b8, 32'hc314e481},
  {32'hc3cf7af0, 32'hc317faf0, 32'hc338ad1b},
  {32'h4445fd75, 32'h436066f6, 32'hc2cc4b8e},
  {32'hc502ad24, 32'h439da5c7, 32'h43943670},
  {32'h44ff8d83, 32'h4353ae49, 32'h4351d8a8},
  {32'hc4aaa41e, 32'hc39553e4, 32'hc30e8ead},
  {32'h439079a2, 32'hc3c186bb, 32'hc3064206},
  {32'hc368da54, 32'hc2daca13, 32'hc3addfe6},
  {32'hc2e55948, 32'hc1734996, 32'hc22dff0a},
  {32'hc500cb5a, 32'hc2a0f5ee, 32'h42a5f8be},
  {32'h4488c827, 32'h4327a212, 32'h4375dc09},
  {32'hc48e9eec, 32'hc21c76b4, 32'h429085ba},
  {32'hc190bbf0, 32'hc31d7977, 32'hc26e453b},
  {32'hc4d52bd8, 32'h430d6bb3, 32'h439ba414},
  {32'h44472789, 32'hc32adb59, 32'h4309a6a0},
  {32'hc50b4172, 32'h439905b8, 32'h43a64aef},
  {32'h43f29784, 32'hc3dee690, 32'hc31e2ee9},
  {32'hc4f10d80, 32'h4109cbd4, 32'h4322bc8c},
  {32'h449d0d25, 32'h4410f09e, 32'hc374ba15},
  {32'h436bdf00, 32'h44037d8b, 32'hc38999d5},
  {32'h4500074a, 32'h43ba1e33, 32'hc38b2e6f},
  {32'hc431101d, 32'hc4198d20, 32'hc1bb29fa},
  {32'h4489d600, 32'hc282b2db, 32'hc19fc45c},
  {32'hc41c15fa, 32'h43fbac3a, 32'hc2aa441c},
  {32'h44ae1e24, 32'h43bda3fb, 32'h43c98300},
  {32'h431422f0, 32'hc2d53603, 32'h42352543},
  {32'h44779a48, 32'hc292800f, 32'h44004465},
  {32'hc40c85ea, 32'h42e6979c, 32'hc3576a12},
  {32'h44bc7f5a, 32'h4288f556, 32'h433acf0a},
  {32'hc47252b4, 32'hc333667e, 32'h42520aa1},
  {32'h439c62a2, 32'hc3f4d183, 32'hc3967d72},
  {32'hc4eb4f44, 32'hc2a983f8, 32'hc3182f2c},
  {32'h443af0dc, 32'hc1f90966, 32'h42a1242e},
  {32'hc4a938e4, 32'hc0acb0b6, 32'hc3885f4c},
  {32'h448e027c, 32'h43e664d5, 32'h41907580},
  {32'hc44fbc90, 32'h436466fe, 32'hc31f2c0c},
  {32'h4451b083, 32'h435a6bcf, 32'h408a4c10},
  {32'hc4fec9af, 32'hbfc209e0, 32'hc3652a25},
  {32'h44e49cfa, 32'h42f7f7f4, 32'h42f176aa},
  {32'hc4b88c12, 32'hc3cf989c, 32'hc4452fed},
  {32'h44c45768, 32'h436baade, 32'h42c870a9},
  {32'hc4a3e92c, 32'h4280efda, 32'hc18abab6},
  {32'h44a96286, 32'hc417b1c7, 32'h4372b123},
  {32'hc449bf50, 32'hc3bb4777, 32'h422ec56c},
  {32'h44fd0d97, 32'h426dad30, 32'hc2e905cf},
  {32'hc5087537, 32'h43755fd3, 32'hc13716f2},
  {32'h44ebccb5, 32'hc3dfb56e, 32'hc30e8a67},
  {32'hc4f67bdd, 32'h42bd7c9b, 32'hc24ecb1b},
  {32'h44187684, 32'hc357f1d5, 32'hc2b1d2d5},
  {32'hc4b7aa56, 32'hc1989c46, 32'hc3cff4ce},
  {32'h44548c6a, 32'hc1f50c3c, 32'h40f38ac6},
  {32'hc4f4408e, 32'hc17d2581, 32'h427c3b1c},
  {32'h44de93dd, 32'h43564ede, 32'h430bf1c8},
  {32'hc50b0be4, 32'h43f829f0, 32'hc36b5d88},
  {32'h4503439d, 32'h438a7724, 32'h43a4c55d},
  {32'hc3893c9f, 32'hc32313e4, 32'hc3bfe285},
  {32'hc3d27424, 32'hc2813c6e, 32'h43bd624b},
  {32'hc4d8869e, 32'hc32ef9ea, 32'h43218620},
  {32'h4507846a, 32'hc33bfde1, 32'h425e3003},
  {32'hc47a920c, 32'h42d559e3, 32'hc1d02f47},
  {32'h43f8c017, 32'hc330f831, 32'hc2a462ba},
  {32'hc428f2a2, 32'hc3eb447b, 32'hc319b5a0},
  {32'h44a46bf4, 32'hc34e3fc2, 32'hc2efeea5},
  {32'hc3493070, 32'h430d301d, 32'hc31f93a4},
  {32'h448538fb, 32'hc2521243, 32'h43086514},
  {32'hc3e08ddd, 32'hc0bc2b17, 32'h4285ae7e},
  {32'h441a9099, 32'h43739d8d, 32'hc317dd12},
  {32'hc29be4e0, 32'h43986b1e, 32'h4324fe7a},
  {32'h4453f6d3, 32'hc1af521f, 32'hc3213237},
  {32'hc50a556e, 32'hc39867c6, 32'h43a4cd69},
  {32'h43881e6c, 32'h4393c358, 32'h434ce3c9},
  {32'hc4fc508a, 32'hc294fb9b, 32'hc278c5bf},
  {32'h44c6ed08, 32'hc3418de7, 32'h43afd47c},
  {32'hc4b2aa16, 32'hc2d9a444, 32'h42005da5},
  {32'h4484674e, 32'h438e0f73, 32'hc2cd2405},
  {32'hc48e8655, 32'hc38feaff, 32'h431fe7cf},
  {32'h4500dfb1, 32'h43081710, 32'hc3ae7651},
  {32'hc4d4b66b, 32'h4303fad7, 32'h430fbbd3},
  {32'h43ffdc88, 32'h43aaae64, 32'hc357e288},
  {32'hc4733338, 32'hc1ba68c2, 32'hc384ba9c},
  {32'h44b7e486, 32'hc3e9dcad, 32'h411b739b},
  {32'hc5074059, 32'h42b30078, 32'hc266a6a5},
  {32'h44d3ae2b, 32'h43ea6b8d, 32'hbf910428},
  {32'hc424ccf6, 32'h438d386c, 32'hc1cd9e69},
  {32'hc3822040, 32'hc250e1fa, 32'hc2b17a83},
  {32'hc46054fc, 32'hc2352f06, 32'h4314a212},
  {32'h44388340, 32'hbfbc87ac, 32'hc2cba1ed},
  {32'hc4b1c443, 32'h43813f4b, 32'h43fe242b},
  {32'h44117d84, 32'hc26ee32a, 32'h434bd8c3},
  {32'hc4e89c86, 32'hc2ea9f3c, 32'h43bf9451},
  {32'h44be64b0, 32'h43012d02, 32'hc2c66dba},
  {32'hc4cb1673, 32'h42b33bfd, 32'hc2bc624a},
  {32'h45078244, 32'h430211ba, 32'h431f04df},
  {32'hc435e861, 32'hc08e5f71, 32'hc2e4866b},
  {32'h45021451, 32'hc2d89688, 32'hc1c21c30},
  {32'hc3e1eaa0, 32'h434e970e, 32'hc205f24a},
  {32'h4492bc3e, 32'h40d88b3c, 32'h43051f57},
  {32'hc3b02d2e, 32'hc1ebccc4, 32'hc392c8c5},
  {32'h446bdb88, 32'h43ac6e33, 32'h4186989f},
  {32'hc413de74, 32'hc39aad8c, 32'h42d850c8},
  {32'h44f49e8a, 32'h3e6892e0, 32'hc1f83647},
  {32'hc4cb4fac, 32'hc20fef66, 32'h42a0b62f},
  {32'h44e54fd2, 32'h43ee477a, 32'hc3c01ae5},
  {32'hc4cab7b2, 32'h42e39461, 32'h4445606e},
  {32'h44d9dba1, 32'hc3a200f4, 32'hc3116850},
  {32'hc4b5bd29, 32'hc3239adf, 32'hc32e83d4},
  {32'h444b05bc, 32'hc3bffc0b, 32'h42e38b7e},
  {32'hc473b761, 32'h42ea2b9a, 32'h43b754e7},
  {32'h4483d1a3, 32'hc4521db8, 32'h43473c73},
  {32'hc4b14c9a, 32'hc2fe4f36, 32'h422b4db5},
  {32'h44798c7e, 32'h406f6316, 32'h43143b26},
  {32'hc498f473, 32'hc3ce1c98, 32'hc2971e52},
  {32'h44f49100, 32'h4282fb6a, 32'hc35efb08},
  {32'hc3c45b80, 32'hc30827a0, 32'hc277ad87},
  {32'h44a53dc7, 32'h42870c32, 32'hc3640cbd},
  {32'hc49b7749, 32'h42c81c5c, 32'h432192ea},
  {32'h44b4cd7d, 32'h4204caeb, 32'h42d0eb20},
  {32'hc4d2e0d5, 32'h438b6071, 32'hc30d3e9e},
  {32'h433de921, 32'hc32a30c0, 32'h41d8b518},
  {32'hc50319fd, 32'hc312ce2f, 32'h43006d6c},
  {32'h448ae81e, 32'h419d2334, 32'hc322a1ba},
  {32'hc1a4cf40, 32'h427a7d8a, 32'h41062346},
  {32'h44435692, 32'hc2c2f5c2, 32'hc2b7a902},
  {32'hc498d174, 32'h428dcac4, 32'hc21ce26b},
  {32'h44586061, 32'h4391df0b, 32'hc2124341},
  {32'hc505537e, 32'hc32b569a, 32'hc1d1317b},
  {32'h445bd7ac, 32'h437f0581, 32'h42b6e74c},
  {32'hc4c6a288, 32'hc3b85381, 32'h4315cea6},
  {32'h447e7e82, 32'h43b9cb41, 32'h42d91805},
  {32'hc4940b27, 32'h42ed1fb5, 32'h42c051b9},
  {32'h45085495, 32'hc1f976eb, 32'hc3154575},
  {32'hc50a5b0a, 32'h4363d492, 32'hc2d63f0e},
  {32'h4478a6f0, 32'hc2864c92, 32'h44110ee6},
  {32'hc4ab69e0, 32'hc1c4b17a, 32'h4253b0e4},
  {32'h450f4e3d, 32'hc3618c88, 32'hc3b55764},
  {32'hc3e82882, 32'hc38ce68f, 32'h4184d9f8},
  {32'h44843bc8, 32'h43a873a3, 32'h433eab9f},
  {32'hc4cbaec7, 32'hc20cd586, 32'hc24bae73},
  {32'h44b0706e, 32'h4320fb71, 32'h438edfe1},
  {32'hc48ebdca, 32'hc3143ae0, 32'hc3723f88},
  {32'h450be652, 32'h42e3514b, 32'h43b5b713},
  {32'hc4a4cfc2, 32'hbf90fc78, 32'h42f77285},
  {32'h4509b0da, 32'h4301f002, 32'hc40d328d},
  {32'hc4e1fccf, 32'h4239f7b3, 32'h439835bb},
  {32'hc239d540, 32'hc2ea3914, 32'h433bb13a},
  {32'hc4a8806a, 32'h4169687d, 32'hc1d703f6},
  {32'h44d6c548, 32'hc3753604, 32'h3fcdaf60},
  {32'hc484e6dd, 32'h42bb35cf, 32'hc262d985},
  {32'h44c17510, 32'hc3981625, 32'hc3c74f3e},
  {32'hc4835171, 32'h404e4569, 32'hc3cff123},
  {32'h44bca29c, 32'h438d4811, 32'h43f957ac},
  {32'hc4ff83ad, 32'h43ef79c6, 32'hc3205928},
  {32'h43852acc, 32'hc3b9e84a, 32'hc1981744},
  {32'hc498b0ca, 32'hc231ab58, 32'h43b404ee},
  {32'h44dbe540, 32'hc2448a78, 32'h42b89485},
  {32'hc39f2365, 32'h43b54cb4, 32'h4370e0a1},
  {32'h43c4ee28, 32'h4346771d, 32'h41c99b24},
  {32'hc47ef2a6, 32'hc2fcae1d, 32'h424ce8fc},
  {32'h44fb390f, 32'h421bcbe4, 32'hc15edaf3},
  {32'hc48f73d4, 32'h43bb87bc, 32'hc1544153},
  {32'h44b9e302, 32'hc3a6e183, 32'hc16794ac},
  {32'hc459cb5a, 32'hc3112eca, 32'h43d3b545},
  {32'h44f3e73a, 32'h433e0f55, 32'h43791054},
  {32'hc48359b9, 32'h425b36a6, 32'h4166745c},
  {32'h43dd82f0, 32'hc283be6e, 32'h434d3c87},
  {32'hc3284cf0, 32'h41dfe156, 32'hc2eb95bd},
  {32'h44d0967a, 32'h436ec4bc, 32'hc304aa77},
  {32'hc4c5c6c0, 32'hc347eea3, 32'hc290ee9d},
  {32'h449af8c0, 32'hc30bd082, 32'hc3887fc6},
  {32'hc472da9a, 32'hc3e66eb5, 32'hc21352f2},
  {32'h4504433c, 32'hc3d60d1a, 32'h440653ea},
  {32'hc46dbb1a, 32'h42e14e54, 32'h43055771},
  {32'h44db5356, 32'hc36a64b9, 32'h434befb1},
  {32'hc5169740, 32'h438f2f26, 32'h4302c446},
  {32'h43f30e30, 32'hc33ef2e2, 32'hc2921707},
  {32'hc4f6680c, 32'h43962902, 32'hc3611952},
  {32'h44b41432, 32'h43a377ec, 32'hc22c6dba},
  {32'hc46375d4, 32'hc3f772af, 32'hc1a4be58},
  {32'h4456aedc, 32'hc34a92ba, 32'hc2d52d76},
  {32'hc4949382, 32'h42de0618, 32'h4385c52f},
  {32'h44bcb5d5, 32'hc3b650ec, 32'h41dfe4d2},
  {32'hc396ceb8, 32'hc33101cd, 32'h43238564},
  {32'h440d8864, 32'h43cb70c6, 32'hc0755e70},
  {32'hc3562d58, 32'h432d8824, 32'h430f9238},
  {32'h423b7040, 32'h439ad1c4, 32'h41c4eafa},
  {32'hc45b2d55, 32'hc3c7bac8, 32'hc2210249},
  {32'h432ecf2a, 32'h432793f3, 32'hc2bb63eb},
  {32'hc50b026b, 32'hc3962ccb, 32'h427dc246},
  {32'h44392f08, 32'h42f65dc1, 32'hc2e6b81b},
  {32'hc48faa52, 32'hc0837f89, 32'hc3d084fb},
  {32'h4508cd4e, 32'h42a81eca, 32'hc2bde0af},
  {32'hc39fdce0, 32'h44024308, 32'hc3d0d070},
  {32'h44754cd6, 32'hc3215948, 32'hc3c8db94},
  {32'hc4a1ff70, 32'h43652424, 32'hc42722ed},
  {32'h448ccf4a, 32'hc290b49b, 32'h42b7187e},
  {32'hc3801728, 32'h437a5892, 32'h428dc864},
  {32'h44ddc016, 32'h43311863, 32'h434ce34b},
  {32'hc4c65e6b, 32'hc2f98e2f, 32'h43a546a6},
  {32'h448793c0, 32'h43dcb258, 32'hc320ee19},
  {32'hc4b43cf7, 32'hc1aa9d34, 32'h430c6fb8},
  {32'h43d521a0, 32'hc223b370, 32'h43925bd4},
  {32'hc479529e, 32'h4379b269, 32'hc3a33f62},
  {32'h44cc2852, 32'h437ea646, 32'h426547b6},
  {32'hc50deec1, 32'hc1af5691, 32'hc2b58b63},
  {32'h43a34a8c, 32'h438f430f, 32'hc2f94241},
  {32'hc3e9fb20, 32'h4417dc3e, 32'h4214aa20},
  {32'h44b13112, 32'hc175e79e, 32'h43075a9c},
  {32'hc4a9d290, 32'h42700082, 32'hc37ba909},
  {32'h4281c82c, 32'hc186ace8, 32'hc32a6197},
  {32'hc5198112, 32'hc305c66c, 32'hc3cf7af1},
  {32'h451be9a4, 32'hc3765688, 32'hc25a4d13},
  {32'hc4b38900, 32'hc349171f, 32'h4034d238},
  {32'h44a0cfd2, 32'h43876439, 32'h41829dc4},
  {32'hc4007c91, 32'h42d6fe56, 32'h433600d6},
  {32'h450dd284, 32'h41b5475f, 32'h42d94b52},
  {32'hc4c62cb5, 32'h43680ade, 32'h428bc833},
  {32'h4508cce1, 32'h4290dc6a, 32'h422fc814},
  {32'hc42869b1, 32'hc300f296, 32'h42dd1365},
  {32'h452364d0, 32'hc30c09b4, 32'h42a02a78},
  {32'hc488b402, 32'hc38c5118, 32'hc2c26c9a},
  {32'h45047a9a, 32'h43ce5380, 32'h4336cced},
  {32'hc484368c, 32'h434f706a, 32'hc3aafe27},
  {32'h44b36767, 32'h436d2f62, 32'h421904df},
  {32'hc2594140, 32'h4295378e, 32'h43a2327a},
  {32'h437b8a00, 32'h4395555c, 32'h4316cbea},
  {32'hc4992219, 32'h43f046bc, 32'h41891809},
  {32'h451ed384, 32'hc28dcbdc, 32'h428828d8},
  {32'hc508cd9e, 32'hc3131091, 32'h42a575b6},
  {32'h449259bd, 32'hc3b8ccb3, 32'hc2c06faa},
  {32'hc4e92cb4, 32'h4301fb3f, 32'hc3277216},
  {32'h4442dec4, 32'hc32ff4da, 32'hc29dd536},
  {32'hc4ab69b0, 32'hc30a711d, 32'h42f46e85},
  {32'h42475804, 32'hc1e6cfae, 32'h434941b0},
  {32'hc4c0a0dd, 32'hc3acfca3, 32'hc38fc276},
  {32'h447f36d2, 32'hc39808a3, 32'h4336ab81},
  {32'hc48049d2, 32'hc30655d3, 32'h430b7528},
  {32'h44758060, 32'h4368f396, 32'h41fdcf64},
  {32'hc4f5b48a, 32'hc334b4ca, 32'hc33fe761},
  {32'h4521080c, 32'hc36898ed, 32'h435368d0},
  {32'hc3d2d6b0, 32'hc2e37b80, 32'hc32b3336},
  {32'h4520f47a, 32'hc2d1c7f8, 32'h4321388e},
  {32'hc409082e, 32'hc208aeec, 32'h41fc327a},
  {32'h44c5a9ec, 32'h422f5694, 32'h4307b6f0},
  {32'hc506f1ba, 32'h4395bf54, 32'h4348e065},
  {32'h44d38496, 32'hc216eee4, 32'hc2109046},
  {32'hc4ef76ff, 32'hc2a0d953, 32'h43835367},
  {32'h43d5a250, 32'h40ccc196, 32'h42c5145f},
  {32'hc4b8396b, 32'hc311b330, 32'hc2cec903},
  {32'h44f156b6, 32'hc2601e13, 32'h42b7fb8f},
  {32'hc485bba3, 32'h4392f4e1, 32'h43720694},
  {32'h44479601, 32'hc1ae5460, 32'hc3830b39},
  {32'hc44f82e0, 32'hc0dfc329, 32'h437c51b1},
  {32'h44fc9bac, 32'h4231c06c, 32'h430c3b95},
  {32'hc354273b, 32'hc2b90586, 32'h413ceba6},
  {32'h44e0fddd, 32'h43c7de32, 32'h43c9eaea},
  {32'hc3d30364, 32'h430de007, 32'h4275c85b},
  {32'h44c5e384, 32'h42e7a7fc, 32'hc13ee6b4},
  {32'hc4729d4d, 32'h43dc1889, 32'h42d600f9},
  {32'h440c86b6, 32'hc2fa833b, 32'h4299409a},
  {32'hc48f3702, 32'hc3004fae, 32'hc2ba6a4d},
  {32'h450d00fe, 32'hc23ddb80, 32'h4381440a},
  {32'hc4085164, 32'h4419745d, 32'hc34d2f57},
  {32'h44972941, 32'h4056bbbc, 32'hc3b70f2a},
  {32'hc3ce37fe, 32'h43437778, 32'h4284f078},
  {32'h44aa2fb0, 32'h4384ddf0, 32'h43001cce},
  {32'hc4a2f8f8, 32'hc2d73658, 32'h42bcad6a},
  {32'h44300316, 32'hc2343426, 32'hc39db454},
  {32'hc4b24094, 32'hc2f5bb3c, 32'h424c1b69},
  {32'hc3104040, 32'hc35b52b7, 32'hc37ff37d},
  {32'hc4147470, 32'h42ce636f, 32'h4189e922},
  {32'h44c73484, 32'h43b3d413, 32'hc3b66850},
  {32'hc46ed088, 32'h4229b985, 32'h434969ec},
  {32'h448aa2f8, 32'hc1eb55f6, 32'hc2bb68ee},
  {32'hc3ea8e9c, 32'hc1d9ac25, 32'hc3909c31},
  {32'h448c4f0a, 32'h4358751f, 32'hc32a049b},
  {32'hc3b5042c, 32'hc18006f8, 32'h430cb4eb},
  {32'h44991281, 32'hc24e9432, 32'hc2cee5c0},
  {32'hc50cab3c, 32'hc38ecefa, 32'hc018aa20},
  {32'h44af32ce, 32'h4217fd82, 32'hc3673b16},
  {32'hc51d295a, 32'hc1814e9a, 32'h43111272},
  {32'h44fe9548, 32'hc2d5a9ce, 32'hbf685870},
  {32'hc36aa55a, 32'hc2466a7d, 32'h439e3a08},
  {32'h43d3ecea, 32'hc3872641, 32'h42bfebfb},
  {32'hc4c6d7db, 32'hc2086a77, 32'h42877c7e},
  {32'h4505d1f0, 32'hc3050da6, 32'h43614379},
  {32'hc4f630ba, 32'h42f78dc8, 32'hc1494e05},
  {32'h4485a3bd, 32'hc31f0939, 32'h434ddc6f},
  {32'hc4621cd0, 32'hc0b74d81, 32'h42a12cf4},
  {32'h44d749d7, 32'hc148cf06, 32'hc3518e5c},
  {32'hc4142c85, 32'hc3353279, 32'hc1a64d18},
  {32'h44855d29, 32'hc2ddcb66, 32'hc145feae},
  {32'hc30444ad, 32'hc3a6554b, 32'h434b6fba},
  {32'h44fe35a1, 32'hc38657cb, 32'h42be1ee9},
  {32'hc3a40310, 32'h42931880, 32'h4213708c},
  {32'h446d7054, 32'hc35e4279, 32'hc2c1e808},
  {32'hc411c5f0, 32'hc3f51572, 32'h417d8b84},
  {32'h44ddbeab, 32'hc24391e3, 32'hc3ab6766},
  {32'hc49e08eb, 32'hc2cd01e3, 32'h43bce5a0},
  {32'h44eeb921, 32'hc294f561, 32'hc3299b73},
  {32'hc40fb683, 32'h436fa2af, 32'hc3510cb9},
  {32'h44837e65, 32'hc3f17097, 32'h437c5624},
  {32'hc405ca04, 32'h42e4da5e, 32'h434490fc},
  {32'h44fa226d, 32'h43ce61c6, 32'hc346800d},
  {32'hc483e5aa, 32'h42f2484d, 32'h42e22d3d},
  {32'h44c8ebc0, 32'hc3da7ac7, 32'hc2fd21cb},
  {32'h44540742, 32'hc3c7ae7d, 32'h432619cd},
  {32'hc35fd2ec, 32'h415d0f95, 32'h42c41908},
  {32'h45085ba6, 32'h432b623b, 32'h4356d54c},
  {32'hc48bcdd4, 32'h42efcc1d, 32'hc3081a58},
  {32'h4470f26f, 32'hc33128fb, 32'h431a8c0b},
  {32'hc3592130, 32'h438e45d4, 32'h43a5950b},
  {32'h44a0aa2c, 32'hc2c3dddf, 32'hc3e9cbde},
  {32'hc431f91c, 32'h437c83d6, 32'hc308dd67},
  {32'h43986120, 32'h4371cf80, 32'hc2df3b7e},
  {32'hc484ff63, 32'hc34a9876, 32'hc3debc4b},
  {32'h43117170, 32'hc3651e49, 32'hc321e3fb},
  {32'hc35f326c, 32'hc323a639, 32'h440546f2},
  {32'h44c79229, 32'h43fa72d2, 32'hc325d66c},
  {32'hc501851b, 32'hc35c6945, 32'h43798bb1},
  {32'h450774c5, 32'hc2e384da, 32'h42b1e3b7},
  {32'hc49808f8, 32'h433e97ec, 32'hc3a49670},
  {32'h448dfbef, 32'h42bed457, 32'hc409dec0},
  {32'hc3542560, 32'hc2337576, 32'h430d611e},
  {32'h4476abc6, 32'hc2897a58, 32'hc3e80791},
  {32'hc373e1f8, 32'hc2f1ae15, 32'hc356df1c},
  {32'h449018ad, 32'h42c29aba, 32'hc37b078c},
  {32'hc498252b, 32'h42b443df, 32'h437bd0dd},
  {32'h4410b530, 32'h436b0c78, 32'hc1a33194},
  {32'hc4eb0678, 32'h42168368, 32'h426aa1eb},
  {32'h43d7b128, 32'h431acd8c, 32'hc2f599e6},
  {32'hc4abf51b, 32'h41d556fe, 32'h4388e9c2},
  {32'h4405202d, 32'hc2675567, 32'hc2951a3f},
  {32'hc226ecc0, 32'hc38186dd, 32'h42241ce0},
  {32'h44dc9940, 32'h42218fe2, 32'h42a3ad77},
  {32'hc3f0e02c, 32'h437bb23c, 32'hc23461e6},
  {32'h442583b9, 32'h42bf1888, 32'h42df5898},
  {32'hc50d2f06, 32'hc3fa1449, 32'h4399df30},
  {32'h44d479ae, 32'h4329b6ac, 32'hc312115d},
  {32'hc2ae0065, 32'hc2b22470, 32'hc385f488},
  {32'h444cb82f, 32'h4358e2a1, 32'hc3120761},
  {32'hc49eb0b1, 32'hc34f75d6, 32'hc1bb548a},
  {32'h43499708, 32'hc2009187, 32'h43c5f3e3},
  {32'hc48bd3ba, 32'h4400816a, 32'hc3ee71b0},
  {32'h4413ca15, 32'h42bf97cf, 32'h432297dc},
  {32'h430650a8, 32'h4342f666, 32'hc3aaded9},
  {32'h44daeb93, 32'hc236f872, 32'hc013eefa},
  {32'hc41e6567, 32'h42b310cd, 32'h43a6a94c},
  {32'h449d71d6, 32'h43cfb56e, 32'hc385ce37},
  {32'hc495104b, 32'h4271a690, 32'hc2b8d63c},
  {32'h4453834d, 32'h438d283a, 32'hc3f0a4b2},
  {32'hc25a1a52, 32'h43ac1c46, 32'h4349ca8c},
  {32'h448fc2ec, 32'hc32e2d86, 32'h430c55ba},
  {32'hc3c4d156, 32'hc37388c3, 32'hc26e29a7},
  {32'h4423444a, 32'h4381842a, 32'hc122137a},
  {32'hc511e462, 32'h4324a15c, 32'hc333f9a0},
  {32'h433177a0, 32'hc36336e2, 32'hc3210f2f},
  {32'hc4f4540f, 32'h432d880e, 32'h43303562},
  {32'h438ee550, 32'h418593e4, 32'h41f18e92},
  {32'hc3d36d17, 32'hc3bc2cd4, 32'hc37c4e61},
  {32'h44b69815, 32'hc3769e61, 32'hc34004d9},
  {32'hc3e9ca90, 32'hc1f13a2f, 32'hc3804b17},
  {32'h44acef36, 32'hc30f56b2, 32'hc2f3eb70},
  {32'hc40e17d0, 32'hc287a8d1, 32'h438d1131},
  {32'h450c73ac, 32'h44566a78, 32'hc2948fa7},
  {32'hc5120459, 32'h4300b152, 32'hc39996c7},
  {32'h44efce23, 32'hc411c619, 32'h422a8912},
  {32'hc3d12d63, 32'hc379f8be, 32'hc3021765},
  {32'h4344d836, 32'h436ac4c9, 32'hc337082a},
  {32'hc40bb264, 32'h4382c257, 32'h433a6f89},
  {32'h443a5dbf, 32'h43c7567c, 32'h430449e2},
  {32'hc4c9fc41, 32'h4423ae9e, 32'hc2e701f7},
  {32'h45071cad, 32'hc20f8e54, 32'hc3bb9199},
  {32'hc4c77e3f, 32'hc3416af9, 32'hc34ffee8},
  {32'h44f73fed, 32'hc30da5db, 32'hc352a84d},
  {32'hc299a41a, 32'h41fe5a96, 32'h42aa0988},
  {32'h4404b452, 32'h429e9b9e, 32'hc2d8555c},
  {32'hc4f1800d, 32'hc381932b, 32'h429e3057},
  {32'h450507c5, 32'hc3ec66a2, 32'hc37b2fcc},
  {32'hc51813ee, 32'h413831e4, 32'hc3e60510},
  {32'h44f84968, 32'h42244a8e, 32'h433232ba},
  {32'hc4f49abf, 32'hc2c664f4, 32'h419d6f91},
  {32'h451374d6, 32'h430bd75e, 32'hc272b242},
  {32'hc48911c9, 32'hc392faff, 32'h4234579f},
  {32'h44f4b7b0, 32'hc28b8b56, 32'h436df763},
  {32'hc4c9c817, 32'hc3329762, 32'hc21d481b},
  {32'h44efe9d0, 32'h42723b27, 32'h4309b705},
  {32'hc3cf0200, 32'h40db4a26, 32'h4308f863},
  {32'h44908197, 32'h435a7229, 32'hc1c32f5e},
  {32'hc395f344, 32'hc2666192, 32'hc36109b6},
  {32'h4416f4c1, 32'hc333d84f, 32'hc24405a1},
  {32'hc494776b, 32'hc3b21600, 32'hc2ab41f4},
  {32'h4406b78b, 32'hc2e22129, 32'hc329cb3d},
  {32'hc4bd1e05, 32'hc22da935, 32'hc3ba4c78},
  {32'h4518e95f, 32'h439a879b, 32'h4172b6d5},
  {32'hc4a9e3de, 32'h4297e00f, 32'hc346b2cf},
  {32'h447df407, 32'h43155739, 32'h41b09e50},
  {32'hc387ff10, 32'h439458c9, 32'h434bcc98},
  {32'h4465d454, 32'h433b4386, 32'hc208dfa2},
  {32'hc49bc63f, 32'hc1c95a5b, 32'hc24a533a},
  {32'h44c30570, 32'h429c9361, 32'hc22daff4},
  {32'hc4c48d16, 32'hc3896df6, 32'h42efd33d},
  {32'hc1b6a380, 32'h438f994b, 32'h436b2497},
  {32'hc39ea326, 32'hc11f9dd6, 32'h42a39793},
  {32'h448bf4f8, 32'h43b193b1, 32'h40a5614e},
  {32'hc50ea4e6, 32'hc390101e, 32'hc3858517},
  {32'h43e8142f, 32'h436adbaa, 32'h423d048b},
  {32'h43a078c8, 32'hbe38d000, 32'h41937abe},
  {32'h44db8a3c, 32'h4343879d, 32'hc34fb217},
  {32'hc4bb1ba8, 32'h43bb191f, 32'h4390db46},
  {32'h43838b00, 32'h433d4910, 32'hc380c88c},
  {32'hc504c525, 32'hbfe56400, 32'h42b7a9e0},
  {32'h44fb8e86, 32'h420cc27e, 32'hc3b5b86b},
  {32'hc4ae079e, 32'hc39bdc6c, 32'hc292578e},
  {32'h4457bd48, 32'hc291da9f, 32'h41189f9a},
  {32'hc51f4727, 32'hc1076446, 32'hc300f2af},
  {32'h4526d016, 32'h43183e14, 32'hc3272fb1},
  {32'hc51855d6, 32'hc2edf617, 32'h427e1164},
  {32'h44ba0820, 32'h42f5392c, 32'hc0bc19d6},
  {32'hc388f8d8, 32'h439652c6, 32'h41d11a2e},
  {32'h451f593e, 32'h42afb932, 32'hc350f747},
  {32'hc50580cc, 32'hc2838003, 32'hc1dbca6e},
  {32'h448a6c9f, 32'hc24fe3a0, 32'hc38d4932},
  {32'hc2babbc0, 32'h430563d0, 32'hc29f4aed},
  {32'h45173a99, 32'hc39228ee, 32'h4382b932},
  {32'hc4eec65e, 32'hc22c2de4, 32'h435c3059},
  {32'h4416168d, 32'h430ce409, 32'h433c7839},
  {32'hc4a9cc24, 32'hc2c5bbc4, 32'hc0338bc0},
  {32'h42f8eca0, 32'hc3ace27b, 32'h43018744},
  {32'hc4e6f2cc, 32'hc3acc568, 32'h430640b8},
  {32'h44e0006f, 32'hc2bcc50f, 32'h43e674ac},
  {32'hc498fb9d, 32'hc3c19717, 32'hc2d3197a},
  {32'h4503d8c8, 32'h43fecfba, 32'h4395b15e},
  {32'hc4f4dc98, 32'h42962f1c, 32'hc267a5bc},
  {32'h44981c99, 32'h42c004dd, 32'h436d83b1},
  {32'hc4f517d8, 32'h4379ea84, 32'h440c9634},
  {32'h4446d65a, 32'hc38cf37e, 32'h43d7ef51},
  {32'hc4cb22d8, 32'h43fe9d97, 32'hc252461d},
  {32'h44cebde4, 32'h424b2029, 32'hc390bf0a},
  {32'hc4e1e1e3, 32'hc3ac54d3, 32'h43e3b696},
  {32'h44efe2ac, 32'hc35a943c, 32'hc31608d5},
  {32'hc1ce7e80, 32'h41fb417f, 32'h42b5f0eb},
  {32'h443e124a, 32'h4360b88c, 32'h43be6d21},
  {32'hc51ba7f0, 32'hc227c383, 32'h43822c9a},
  {32'h44df3d2c, 32'hc2e2845d, 32'h43a3b156},
  {32'hc49cee8c, 32'hc3c8dd14, 32'h43adeddb},
  {32'h445b3002, 32'hc07bdfa4, 32'hc30d4acc},
  {32'hc3934a68, 32'h42e14624, 32'hc25def66},
  {32'h44f76c39, 32'h420f1767, 32'h42237f95},
  {32'hc3c377c0, 32'hc397e6ed, 32'h42b1ed79},
  {32'h443b9bfa, 32'hc3bbc952, 32'h4341e09f},
  {32'hc4e84c8e, 32'hc300e828, 32'h42e443f8},
  {32'h450e516b, 32'h42883516, 32'hc39b330a},
  {32'h4360fb80, 32'h43ac5a78, 32'h43828b3c},
  {32'h45195903, 32'h42b75874, 32'h439443c7},
  {32'hc4972538, 32'h4296cb79, 32'hc3aae6d0},
  {32'h4480fd00, 32'h43106ffc, 32'hc28bb950},
  {32'hc4c13122, 32'hc3056702, 32'h4359db01},
  {32'h44e1ff50, 32'h4388d440, 32'h423bf1a5},
  {32'hc4f3ae2c, 32'hc132efe3, 32'h42bb5f47},
  {32'h4371dc33, 32'h42e52f77, 32'h42ebd3cc},
  {32'hc4fbca64, 32'hc3051d89, 32'hc223afc6},
  {32'h451317a3, 32'hc404208b, 32'hc321c265},
  {32'hc38463e0, 32'h428bdf28, 32'hc3131241},
  {32'h43ea3f2b, 32'hc03e6bc0, 32'h41e53ea9},
  {32'hc4eda88a, 32'h4395917f, 32'h42884302},
  {32'h44c06b03, 32'h42c8dcaa, 32'h4357bee5},
  {32'hc42951a7, 32'hc3bf3f12, 32'h429d47be},
  {32'h4502235f, 32'h42f2cf77, 32'hc33e5983},
  {32'hc488828b, 32'h431c33e2, 32'h438d6982},
  {32'h449c1eff, 32'h43700c0c, 32'h434692c7},
  {32'h42830760, 32'h435184c4, 32'h43910675},
  {32'h44d86a98, 32'hc33c6faa, 32'hc294c2b1},
  {32'hc3fcc6e4, 32'h4365d4a1, 32'hc3a0d460},
  {32'h445d8673, 32'h426af08c, 32'h437c9b8b},
  {32'hc46fc948, 32'hc3b7fb35, 32'hc281df93},
  {32'h44918d44, 32'h43e9ea75, 32'h42c20e2e},
  {32'hc2c64480, 32'hc29696bb, 32'hc34fe586},
  {32'h44d30fa0, 32'h4408a05e, 32'h43296380},
  {32'hc50b31f5, 32'h435d8384, 32'hc3a6514b},
  {32'h440bdd20, 32'hc2a1c377, 32'h4347240f},
  {32'hc4148440, 32'h423d4429, 32'hc282da71},
  {32'h448f27de, 32'h428b7f6e, 32'hc2a242ba},
  {32'hc4a29408, 32'hbf7509bc, 32'h42ac4637},
  {32'h43e7800c, 32'h4389d349, 32'h41b4e21c},
  {32'hc4f9ae6a, 32'hc3ce0bfe, 32'hc38995e0},
  {32'h4519a8fe, 32'h43300dfb, 32'h4296d019},
  {32'h434c71f0, 32'hc1296770, 32'hc2391413},
  {32'h44ebd0ff, 32'h428f1318, 32'h42c2ca35},
  {32'hc49ab941, 32'hc281c756, 32'hc14ad006},
  {32'h44a7b9fc, 32'hc2d60234, 32'h423a50ee},
  {32'h4236cbc0, 32'h42a77c3b, 32'hc3436853},
  {32'h45127ec1, 32'hc3687f94, 32'hc315a28f},
  {32'hc38e1e24, 32'h412a48c2, 32'h41d26386},
  {32'h44942128, 32'hc1131e65, 32'h4323adff},
  {32'hc46d0363, 32'h432c9581, 32'h430877e6},
  {32'h436df260, 32'hc350b579, 32'h43938d43},
  {32'hc3c078a4, 32'hc25e0983, 32'hc3997771},
  {32'h450adadd, 32'hc306aded, 32'hc33bc85a},
  {32'hc321204e, 32'hc1dca3fb, 32'h4372fbda},
  {32'h447d4345, 32'h439724bb, 32'h431b5eee},
  {32'hc4b109f0, 32'h432322e4, 32'h42bf3aac},
  {32'h437dd21a, 32'h43ea3984, 32'h43bbc311},
  {32'hc4e9914a, 32'hc3166d32, 32'h4299dd17},
  {32'h433d3200, 32'h41f4cebf, 32'h432a78e6},
  {32'hc4d938c9, 32'h4357cbe2, 32'hc2adab65},
  {32'h45082b3b, 32'h423a0af4, 32'hc302a745},
  {32'hc43511cd, 32'h4328a779, 32'h436c5fed},
  {32'h44e469b8, 32'h439f22d7, 32'hc40397ab},
  {32'hc50ba78c, 32'hc3de976c, 32'h43d43a18},
  {32'h442482d4, 32'h4381e5e4, 32'h412fdccc},
  {32'hc497e359, 32'h4340bda5, 32'h4359e113},
  {32'h45084f70, 32'hc3524c19, 32'hc21ee1de},
  {32'hc4ec500b, 32'h43d6020f, 32'hc384eacc},
  {32'h4485c912, 32'h42ff5cef, 32'h42009490},
  {32'hc48d3347, 32'hc3c490cf, 32'h439c7a6e},
  {32'h44221f1a, 32'h43bb5444, 32'h431d9667},
  {32'hc4fca7d5, 32'h430be1d0, 32'hc1fc7393},
  {32'h440ca1f0, 32'hc23c9847, 32'hc306eb76},
  {32'hc3a52224, 32'hc3c27acb, 32'h408dfdc2},
  {32'h4498cfc4, 32'hc2964b70, 32'h4283518f},
  {32'hc40abf0c, 32'hc3a4753b, 32'hc358dfa0},
  {32'h44df4ca0, 32'h42aaa8ed, 32'hc2cba44b},
  {32'hc4cde06e, 32'hc1e8ad49, 32'h42191440},
  {32'h4400b394, 32'hc295cd2c, 32'hc35e38b8},
  {32'hc2afaace, 32'hc38ab88e, 32'hc22a8a3b},
  {32'h439f4175, 32'h416c9f1a, 32'h40c23077},
  {32'hc40aa500, 32'hc3175f6f, 32'h432ff51c},
  {32'h44fd0639, 32'hc1201aa7, 32'h4279b52b},
  {32'hc4c19deb, 32'h435ce55b, 32'hc38b83c1},
  {32'h435aec00, 32'hc1233ffc, 32'hc2c90baa},
  {32'hc4ca2887, 32'h4322e5dc, 32'hc2b40039},
  {32'h4431e9f2, 32'h43fe69da, 32'h42dc7e02},
  {32'hc37fae96, 32'h43ba1493, 32'hc2fa81aa},
  {32'h436aee90, 32'hc319a17c, 32'h430151cb},
  {32'hc35cc956, 32'h42f1d8e9, 32'hc42c90c4},
  {32'h44d55a6d, 32'hc33ce45a, 32'h4224a03f},
  {32'hc518583a, 32'h4310f358, 32'hc38521d7},
  {32'h449039f1, 32'hc1afcd32, 32'hc33b6cd5},
  {32'hc4021a34, 32'h421ee46f, 32'h427cd524},
  {32'h4491177b, 32'hc028e070, 32'hc29635a9},
  {32'hc352f630, 32'hc2bdc74f, 32'hc33ae743},
  {32'h4425dea6, 32'h430d32e9, 32'h43735242},
  {32'hc4e6519e, 32'hc3a2dc36, 32'hc360e29f},
  {32'h42694050, 32'hc45372aa, 32'h43290b7c},
  {32'hc3871d48, 32'hc22fca58, 32'h430ca860},
  {32'h44a4267b, 32'hc39287b0, 32'hc39b6e24},
  {32'hc4e63425, 32'h41a38c55, 32'hc299d621},
  {32'h44ddb42d, 32'h43c0e8bc, 32'h42dd963a},
  {32'hc4940450, 32'h421b687f, 32'h43a8edff},
  {32'h4442cb98, 32'hc1897b98, 32'hc34b5f80},
  {32'hc4dbf66b, 32'h4390c662, 32'hc3fca7c7},
  {32'h44f1af90, 32'hc32d63f0, 32'hc1796c11},
  {32'hc4706ce8, 32'hc37c0ac8, 32'hc2553476},
  {32'h450146d6, 32'h4329231f, 32'h43053b3b},
  {32'hc430316a, 32'hc37698aa, 32'h4385ea4d},
  {32'h44816581, 32'h4341deb6, 32'hc32c8f94},
  {32'hc2873594, 32'hc20a0441, 32'hc1bc66bc},
  {32'h44e59775, 32'hc3d432bf, 32'h43d858a2},
  {32'hc475bc58, 32'hc34f7072, 32'hc363dd3c},
  {32'h44c79036, 32'hc2b0b089, 32'hc2c3665c},
  {32'h42b21cc0, 32'hc3889f1e, 32'hc2de5904},
  {32'h44b3d3f4, 32'hc289f45e, 32'hc3519bc8},
  {32'hc47dea24, 32'hc27f6fee, 32'hbfe0feb0},
  {32'h447910e8, 32'h428e32f8, 32'h4232ad72},
  {32'hc4ee741e, 32'hc3c5bfb2, 32'h43656655},
  {32'h44f93bfe, 32'hc3a0f6f5, 32'hc2ad5bd0},
  {32'hc4963d34, 32'hc3aa76ef, 32'hc2c3bc43},
  {32'h452090a4, 32'hc15f1ee8, 32'h41e3730a},
  {32'hc3fd22a1, 32'hc381e4d6, 32'hc2a56704},
  {32'h44c0236f, 32'h42d8f0c1, 32'hc176e62a},
  {32'hc4ebe2b0, 32'hc3022eb0, 32'hc30b1870},
  {32'h44dfded3, 32'h424abc6b, 32'h418b07d4},
  {32'hc4df1ce5, 32'h43246e7d, 32'h43118ad1},
  {32'h44bbb646, 32'hc19aeda2, 32'h4093c4c7},
  {32'hc4fe9ee7, 32'hc1837c4b, 32'hc38eb32f},
  {32'h4333a22c, 32'hc3a64cd8, 32'h41d668d6},
  {32'hc3bfbe20, 32'h428fb4d5, 32'h43c21b18},
  {32'h44c5ace2, 32'h4317b348, 32'hc412362c},
  {32'hc51b736a, 32'hc286717e, 32'h42e43053},
  {32'h45051e73, 32'hc33f8156, 32'hc3fff7f4},
  {32'hc4266a1a, 32'hc327042c, 32'h43b934a0},
  {32'h440713b2, 32'hc3a1605c, 32'h426d8c9c},
  {32'hc42a3afc, 32'hc2c38eb5, 32'h4303fa3a},
  {32'h44bc5e65, 32'hc09a5ea2, 32'h43a9d58c},
  {32'hc50b067d, 32'h440d0b4d, 32'hc34c3758},
  {32'h44021828, 32'hc3ce9fa9, 32'hc36c0c52},
  {32'hc47eaa16, 32'h4301d569, 32'hc4071a37},
  {32'h44b16e11, 32'h42eb12a7, 32'h43007760},
  {32'hc4e065bc, 32'hc3b62e11, 32'h4271359c},
  {32'h45248c12, 32'hc29943c7, 32'h4363d998},
  {32'hc4b3b93d, 32'hc3b4a689, 32'hc1d1f5e8},
  {32'h42ea0670, 32'h438b6f7f, 32'hc38e1c12},
  {32'hc4ceefde, 32'h41ee9fdc, 32'hc23180c7},
  {32'h44d949bc, 32'hc3283947, 32'h4319448c},
  {32'hc5072be4, 32'h42f46c45, 32'hc3c06018},
  {32'h44134728, 32'hc41a8e3d, 32'h43ac443d},
  {32'hc4ef5b92, 32'h435464e8, 32'h439394b7},
  {32'h447c0e60, 32'h43034ed1, 32'h432aef47},
  {32'hc50a3f22, 32'h4372e80a, 32'h435bfa3f},
  {32'h44945ee3, 32'h3fb05dc4, 32'hc2e78ad8},
  {32'hc436ad77, 32'hc383e9d4, 32'h42411532},
  {32'h44c89c5a, 32'h43899789, 32'h43125678},
  {32'hc508afae, 32'h42f11847, 32'h4400a6f6},
  {32'h4473fe17, 32'h43e6957e, 32'h421ef361},
  {32'hc4d2c36d, 32'h4366b112, 32'h435cad90},
  {32'h4481b75f, 32'hc3b19405, 32'hc3313ce5},
  {32'hc48d523b, 32'hc05c0024, 32'h43c5230c},
  {32'h4495272e, 32'h414dbac9, 32'hc29055a4},
  {32'hc459a17d, 32'hc1bdc4b1, 32'h42c785de},
  {32'h44a0d768, 32'hc3050633, 32'h41832a56},
  {32'hc4419ea6, 32'h4354578a, 32'h440f1db5},
  {32'h45257035, 32'h40d2029e, 32'h42be1aa8},
  {32'hc4cf50af, 32'hc13eae9e, 32'hc2e31bc7},
  {32'h4502e744, 32'h4309ac46, 32'h434c268f},
  {32'hc44a11b5, 32'h407d43be, 32'h4397bc4c},
  {32'h436127a0, 32'h4396b890, 32'h41144516},
  {32'hc4e0fb14, 32'hc3007e6d, 32'hc330164f},
  {32'h44a23043, 32'h43bd1068, 32'h43846f02},
  {32'hc41d148a, 32'hc31c50b6, 32'h41c120d8},
  {32'h4467bc7e, 32'h40ee65b6, 32'hc32706b6},
  {32'hc40864e6, 32'hc383e2da, 32'hc413da61},
  {32'h44fc154a, 32'h438f1d55, 32'h43565019},
  {32'hc3a5dcb8, 32'h438fcdd3, 32'hc29ac5f2},
  {32'h44f0f6bc, 32'h438facb8, 32'hc27f22d3},
  {32'hc4e5a162, 32'hc3efe6df, 32'hc3f87413},
  {32'h440d66a8, 32'hc39457a0, 32'hc30d7939},
  {32'hc4adb9d7, 32'hc3825e5b, 32'hc2ca5a56},
  {32'h44d003f3, 32'h43c426e6, 32'h434e57ad},
  {32'hc4b61c4f, 32'hc3269c3f, 32'hc3131762},
  {32'h44578ca4, 32'hc2b2ebd4, 32'h4388da1f},
  {32'hc50d5ec8, 32'h42e41254, 32'hc3a5410b},
  {32'h450d4e3e, 32'h4335e064, 32'hc30426e4},
  {32'hc49a037a, 32'hc3168371, 32'hc2c647d4},
  {32'h4424eee4, 32'hc1b67d28, 32'hc391448b},
  {32'hc48e4644, 32'h432eb118, 32'h4401ca31},
  {32'h444855ed, 32'hc290deb4, 32'hc1daa3e8},
  {32'hc4f6fce7, 32'h431f1e6c, 32'hc3494e07},
  {32'h44130a10, 32'hc3146041, 32'hc2bf2b5c},
  {32'hc42b4724, 32'hc2a53db2, 32'h42d31674},
  {32'h43493b74, 32'h4308bd3a, 32'h424b1b31},
  {32'hc507cbdd, 32'hc2c18417, 32'hc2d0e04c},
  {32'h45159227, 32'hc212dddf, 32'h425ce9da},
  {32'hc363ec04, 32'hc37a8d79, 32'hc39cf4e6},
  {32'h44eb318f, 32'h420d895d, 32'hbfe80666},
  {32'hc4649bda, 32'hc397fe94, 32'h435eca38},
  {32'h43344f80, 32'hc11637d3, 32'hc37d0a43},
  {32'hc488e372, 32'h43a17ac6, 32'hc236f427},
  {32'h442bf570, 32'hc356062a, 32'h42e8066c},
  {32'hc4808132, 32'hc1c3c67d, 32'h42ec22b1},
  {32'h450635d4, 32'hc2415c62, 32'hc3ce8197},
  {32'hc3c4c608, 32'h42e2c207, 32'hc3164374},
  {32'h44689a8e, 32'h426f6326, 32'hc39e1da9},
  {32'hc4efab48, 32'h43641936, 32'hc3ca7a0f},
  {32'h45062000, 32'h438392bf, 32'hc3f22899},
  {32'hc4bf25d0, 32'hc22d87e8, 32'h433a81e2},
  {32'h43eb9124, 32'hc0098711, 32'h43c23032},
  {32'hc3b919c5, 32'h43943a6e, 32'h4119224a},
  {32'h4455c4fe, 32'h42c4e9f1, 32'hc38ae2f2},
  {32'hc4e475bc, 32'h43926bb8, 32'hc36fe2a3},
  {32'h444e8602, 32'h43b7299f, 32'hc389c0dc},
  {32'hc4d61e08, 32'h42e37f1e, 32'hc21bf605},
  {32'h44e8a524, 32'hc2b7a6df, 32'hc29d6f4d},
  {32'hc4e81d5b, 32'hc28c402a, 32'hc0bbe058},
  {32'h443b8e5e, 32'h4361c1d0, 32'hc203b693},
  {32'hc4b3e456, 32'h42ee3996, 32'h43743e17},
  {32'h44819514, 32'h42bcae23, 32'h43687f7c},
  {32'h43617ea8, 32'hc3a7d318, 32'hc3b537b4},
  {32'h44c4d166, 32'hc32f763d, 32'hc2cec187},
  {32'hc4d86f8e, 32'h435e62a1, 32'hc32825ed},
  {32'h444fe3db, 32'hc38cca32, 32'h42f8f25a},
  {32'hc4d69e85, 32'hc2e294af, 32'hc38ed5eb},
  {32'h44a19db2, 32'h416a3b88, 32'hc1baf3c8},
  {32'hc4f8d6cd, 32'hc0d35bbe, 32'hc3026967},
  {32'h450acdd1, 32'hc2ba48f4, 32'h42414137},
  {32'hc363c6c0, 32'hc39da91a, 32'h43927deb},
  {32'h44549529, 32'h42489bdb, 32'h42519b96},
  {32'hc3771130, 32'h42a27379, 32'hc307e5fe},
  {32'h4382d600, 32'h42898914, 32'hc268590a},
  {32'hc408f160, 32'h42e2de4b, 32'hc1af8857},
  {32'h43ed5200, 32'hc1083a0e, 32'h42458b4e},
  {32'hc49d474e, 32'h42a3dd78, 32'h42a4f280},
  {32'h4519ab04, 32'h4282ca33, 32'h43197664},
  {32'hc3c3a2f1, 32'h439b6314, 32'hc2b33580},
  {32'h44149501, 32'hc2882ebc, 32'h436c41de},
  {32'hc312661b, 32'hc30f3b33, 32'h42eb21ba},
  {32'h4488ac40, 32'hc3522980, 32'h42d0120f},
  {32'hc4f4062a, 32'hc33d29ee, 32'h43eee60a},
  {32'h44039b62, 32'h422459a0, 32'hc3340ef0},
  {32'hc50212ca, 32'h43f10103, 32'h42c189ac},
  {32'h43920302, 32'hc335dcc6, 32'hc30ef8f9},
  {32'hc35b9728, 32'hc39cbf7e, 32'h43a27d4d},
  {32'h44c7c372, 32'hc3e00737, 32'hc19c8df5},
  {32'hc497747c, 32'h43ab9830, 32'hc3838105},
  {32'h4424561c, 32'h43fb8f32, 32'h430270ec},
  {32'hc358a710, 32'hc08f4d98, 32'h4381ccdc},
  {32'h448e8465, 32'h4364adac, 32'hc31c551a},
  {32'h42020f00, 32'hc2d496ba, 32'hc2b9f383},
  {32'h44aec2b7, 32'h434c9d75, 32'hc3f4bab5},
  {32'h4129fecc, 32'hc40efca7, 32'hc32a565b},
  {32'h44eb5128, 32'h43809622, 32'hc37a3c2c},
  {32'hc4c54501, 32'hc20eee1a, 32'hc20f3e20},
  {32'h439fe488, 32'h4128dab0, 32'hc29f8790},
  {32'hc4908299, 32'h429218b3, 32'hc2f077b6},
  {32'h44f156ea, 32'h41a87cbf, 32'h4350a962},
  {32'hc4ff36a6, 32'h4312d459, 32'h4380fb52},
  {32'hc3e3c36e, 32'hc442e2f0, 32'hc2239322},
  {32'hc45a6d72, 32'h4262044a, 32'hc32492bb},
  {32'hc2bd7740, 32'h4392afdc, 32'h43ea1082},
  {32'hc3dd760c, 32'h42547464, 32'hc280dee4},
  {32'h449077d5, 32'h42b5a251, 32'h419f9fb2},
  {32'h41d21780, 32'hc2f4673a, 32'h428c4bdf},
  {32'h44c06ece, 32'h43bfbbae, 32'hc09ce422},
  {32'hc43cce66, 32'hc2fc7684, 32'hc3eb2ccf},
  {32'h44f3f2dd, 32'h43603dfb, 32'h43993705},
  {32'hc3f917bf, 32'h4295c92e, 32'h421052f4},
  {32'h4490ccc4, 32'h43b250a5, 32'h42930f77},
  {32'hc4d79c0f, 32'h4261c022, 32'hc2794670},
  {32'h4458b331, 32'h433cfee5, 32'hc2ecbc14},
  {32'hc4d8b1d1, 32'hc1b56588, 32'hc195195a},
  {32'h44b6fe7d, 32'h409aee6c, 32'h4294a8fa},
  {32'hc44d2f61, 32'h41c4a0b1, 32'hc25392f6},
  {32'h44937310, 32'hc2e5a313, 32'h43891dad},
  {32'hc501dbc7, 32'h43ddf33e, 32'h433fa7e3},
  {32'h44dd6fb1, 32'hc3fe9009, 32'h43032811},
  {32'hc4d8b4c8, 32'h420e2006, 32'hc307b147},
  {32'h432f60b0, 32'h429bd836, 32'h4284fadf},
  {32'hc42e08a3, 32'hc3e94fff, 32'hc3d880c0},
  {32'h4520d5f3, 32'hc2115fac, 32'h41bdec73},
  {32'hc49b46bb, 32'h428507a5, 32'hc3b70627},
  {32'h4502c80f, 32'h42200d3a, 32'hc303f0d7},
  {32'hc46262a3, 32'h429df45d, 32'hc2ced62f},
  {32'h44e861e1, 32'h42b25e32, 32'hc4152fcf},
  {32'hc4d5af64, 32'hc41ddf57, 32'hc37987db},
  {32'h4491f6c0, 32'h43e7f5fa, 32'h42cba99f},
  {32'hc4860487, 32'hc30bcdba, 32'hc3214908},
  {32'h44fc6f81, 32'h421f6b9c, 32'h42c11af8},
  {32'hc4a821ab, 32'hc3e964d2, 32'h434eacc5},
  {32'hc4bf9401, 32'h4219b6ef, 32'hc3106c5a},
  {32'h448252be, 32'h40b00950, 32'h42808a68},
  {32'hc32dc3c4, 32'hc3ad8e33, 32'h43d70b3a},
  {32'h44852c22, 32'h4349428a, 32'hc2dcf798},
  {32'hc4bb7d3d, 32'hc2e5d5de, 32'hc33e3202},
  {32'h4412fe0e, 32'h4392d560, 32'hc350e656},
  {32'hc46fe6e3, 32'hc0f8d2fd, 32'hc2e5361d},
  {32'h44ca6ca0, 32'hc3d28335, 32'h423f25e9},
  {32'hc516e767, 32'h4396aca1, 32'hc394151f},
  {32'h42f94f38, 32'h43198b01, 32'h42d03ed9},
  {32'hc4401eb2, 32'h42ac2f54, 32'hc37bbe14},
  {32'h445a9894, 32'h43ce9cd4, 32'h4347db68},
  {32'hc4837056, 32'h43ee4a04, 32'h412fb80b},
  {32'h44f49150, 32'h43294ec7, 32'h43a01edd},
  {32'hc4299490, 32'h43cc0a77, 32'h40c59dc5},
  {32'h449421ef, 32'h431f6a3b, 32'h431ba5e9},
  {32'hc495cdb6, 32'h42c8882e, 32'h4131b207},
  {32'h44d1618d, 32'hc2b5a4a5, 32'h42ac6c1b},
  {32'hc3cbf768, 32'h43abd266, 32'h430ab497},
  {32'h44db1f77, 32'hc359dfd4, 32'hc3278da2},
  {32'hc4a03e8e, 32'hc20c0530, 32'hc2fb94e6},
  {32'h44e0ff99, 32'hc395f6f3, 32'h43110011},
  {32'hc411d2a8, 32'hc3b33597, 32'hc385352d},
  {32'h4505da5a, 32'h433e63d5, 32'h42510fbf},
  {32'hc39f3208, 32'hc3c8cb7a, 32'h4290269b},
  {32'h44381527, 32'hc37c8a25, 32'h43749e48},
  {32'hc4fb9b50, 32'hc2e362bb, 32'h43b61ebc},
  {32'h42dbfeb8, 32'hc34315e4, 32'h43521157},
  {32'h404e0d32, 32'hc1fe2c68, 32'hc3c8e76f},
  {32'h436b1344, 32'h42b9cbd8, 32'hc30acf4d},
  {32'hc50bd2e2, 32'hc36e6608, 32'hc0cbf571},
  {32'h440c5b12, 32'hc32fa4a0, 32'hc2a02df5},
  {32'hc4fd4bc6, 32'h42657517, 32'h43c0e6b5},
  {32'h450153d8, 32'hc31eb034, 32'hc1a7967b},
  {32'h42fc41a8, 32'hc2859028, 32'hc2e6753a},
  {32'h4493b2d2, 32'h435eef15, 32'hbf8faab5},
  {32'hc46b9dc2, 32'h43816a25, 32'hc449cd81},
  {32'h44cb9760, 32'h42b21615, 32'h43710148},
  {32'hc47a9aa0, 32'hc10aa8e6, 32'h432af3bb},
  {32'h44965f90, 32'h42c12c96, 32'hc208215d},
  {32'h42be2670, 32'hc3400940, 32'hc2704a84},
  {32'h44e40aa3, 32'h3f5a6bd8, 32'h43740165},
  {32'hc16e4040, 32'hc21c4e51, 32'hc2a36b5d},
  {32'h44013d28, 32'hc3d93d9a, 32'hc2fa8343},
  {32'hc50c5f36, 32'hc315fc4a, 32'hc390f8fc},
  {32'h44320652, 32'h43a9728c, 32'hc2a61fe2},
  {32'hc5047c71, 32'h42a551f1, 32'hc37ba1e5},
  {32'h43efac40, 32'h43ab1c8c, 32'h440f0a8c},
  {32'hc49b432a, 32'h433e45a5, 32'hc2a29fea},
  {32'h44b9ce1d, 32'h42c5d25c, 32'h42de9966},
  {32'hc4524ade, 32'hc20f59a0, 32'h40ea6f2b},
  {32'h4415173c, 32'hc3514448, 32'hc2a85854},
  {32'hc45a2c14, 32'h4336f1f7, 32'hc315edf4},
  {32'h44b50718, 32'h41cd8680, 32'hc385e432},
  {32'hc3a77c64, 32'hc30ed988, 32'h4250ea64},
  {32'hc0e8a300, 32'hc37ac1c7, 32'hc407d3b6},
  {32'hc47c3b60, 32'hc35a7c40, 32'h42cf5a2b},
  {32'h45004f78, 32'hc2495550, 32'h42a3fa19},
  {32'hc4d20b88, 32'hc2cb8f98, 32'h42ba7231},
  {32'h438cae75, 32'hc2e23993, 32'hc2471e6b},
  {32'hc3feea60, 32'hc3d18d89, 32'hc232884c},
  {32'h450bc488, 32'h42e44a37, 32'h42864292},
  {32'hc4525327, 32'h43a62ef5, 32'hc26ae13a},
  {32'h44e88d8a, 32'hc3ca1b90, 32'h43042c84},
  {32'hc4adbff0, 32'hc32831b5, 32'hc37a493d},
  {32'h44e8231e, 32'hc3437e90, 32'h428ab1de},
  {32'hc4da7fce, 32'hc286c989, 32'h431f6310},
  {32'h450f172a, 32'hc338166a, 32'h43789919},
  {32'hc46e79c4, 32'hc2f42e9a, 32'hc2adb1a9},
  {32'h44ef87ec, 32'h438178a4, 32'h440ad2d7},
  {32'hc263fea2, 32'h4376105b, 32'hc2513df2},
  {32'h43fa26ff, 32'hc39bbab8, 32'h43a3503c},
  {32'hc4f6c4b0, 32'h4368dc6a, 32'hc3adca4f},
  {32'h45046b2d, 32'h42cb3684, 32'hc32ef7eb},
  {32'hc5088392, 32'hc3afb314, 32'h42776692},
  {32'h44f3e88c, 32'h42882bb4, 32'hc385bced},
  {32'hc4387d5c, 32'hc3a3103f, 32'hc3543e22},
  {32'h4494c35a, 32'h439952e4, 32'hc39aa134},
  {32'hc38c3fe0, 32'h4308b169, 32'hc364a301},
  {32'h449f6054, 32'hc33db8eb, 32'h4367633c},
  {32'hc4ce2710, 32'h432bdb1d, 32'hc3b3d100},
  {32'h4432fb34, 32'hc25d3292, 32'h42f56dd6},
  {32'hc4d83f2d, 32'h434812c2, 32'h43e73cba},
  {32'h43da5388, 32'hc37b8ac7, 32'h432a2b7d},
  {32'hc4cf1432, 32'hc374fa1a, 32'hc3b29b8f},
  {32'h44cde4e2, 32'hc3943059, 32'h418a6a78},
  {32'hc4148d4e, 32'hc2392293, 32'hc2ec1987},
  {32'hc3142810, 32'hc383278d, 32'h429e9ca2},
  {32'hc3dcfc34, 32'hc3b775fd, 32'h4269af09},
  {32'h444ca01a, 32'h4348e7a0, 32'hc3402d3a},
  {32'hc4da86f8, 32'hc380a7c1, 32'hc1067e66},
  {32'h450429ad, 32'h43652a70, 32'h4220e11f},
  {32'hc4e248fe, 32'h41d0bc6b, 32'hc2fa89ce},
  {32'h44519d22, 32'hc349380c, 32'h4166aefc},
  {32'hc402a80a, 32'h41b1d153, 32'h4290bca2},
  {32'h450bfbf4, 32'hbf40116b, 32'hc36df221},
  {32'hc4a2bce1, 32'h42cc36c2, 32'hc3a790ed},
  {32'h4411ce21, 32'hc2d70683, 32'h42900327},
  {32'hc4c32246, 32'hc3b7df5e, 32'h40c612cb},
  {32'h44994700, 32'h42a84662, 32'hc2d4ce3f},
  {32'hc4a3ae44, 32'hc3f61d1f, 32'h42800149},
  {32'h44e943b2, 32'h435665c4, 32'hc325a323},
  {32'hc45a7f4e, 32'h4322c92c, 32'hc355479d},
  {32'h451ba02d, 32'hc3211c86, 32'h4311e159},
  {32'hc4d4f732, 32'hc3ad29bd, 32'h431e33e2},
  {32'h43cbb192, 32'hc3abc9a0, 32'h42d685de},
  {32'hc4ef2f40, 32'hc3336c4b, 32'hc337266c},
  {32'h43bc04c8, 32'hc39faaba, 32'h42262f7a},
  {32'hc4c7b6d9, 32'h43168c09, 32'hc24f8026},
  {32'h440edb9e, 32'h4261a851, 32'hc3547dae},
  {32'hc4788ce4, 32'hc31a2d7a, 32'h412df058},
  {32'h44a35539, 32'h43b06a04, 32'h421e81f8},
  {32'hc4c83377, 32'hc379b9ba, 32'h43227ec9},
  {32'h437194d5, 32'hc214582c, 32'hc35cad5a},
  {32'hc3670950, 32'hc2a1666a, 32'h434e54ce},
  {32'h444697d5, 32'hc3c96d3b, 32'hc35e34b5},
  {32'h43f84810, 32'hc29e31f5, 32'h4303635d},
  {32'hc30f7030, 32'h43998cb5, 32'hc13c3aa9},
  {32'h44f6f5cf, 32'hc3262729, 32'hc212a978},
  {32'hc3fb0d54, 32'h429a7451, 32'h42970974},
  {32'h43ab81a8, 32'h43e734d0, 32'hc32df1bf},
  {32'hc493ee2c, 32'h43947d58, 32'h43330139},
  {32'h44bc6b0a, 32'h439546cd, 32'h42eacd79},
  {32'hc46f7bd9, 32'hc20ddbf7, 32'h4358cb6b},
  {32'h4493a603, 32'h438dc8a7, 32'hc354c744},
  {32'hc3f16640, 32'hc2b5c21e, 32'h43747043},
  {32'h43b3d858, 32'h42736fba, 32'hc2ed8d43},
  {32'hc4b8efab, 32'hc40472e1, 32'h430b1550},
  {32'h43367c44, 32'hc28a9e3a, 32'hc30145bd},
  {32'hc3c2ee60, 32'hc14d4e9b, 32'hc25405b6},
  {32'h44df73d6, 32'hc3aab973, 32'h439abac7},
  {32'hc44fb83c, 32'h429c2236, 32'hc3aea5b6},
  {32'h4490409e, 32'hc2ec6b82, 32'h42d04f58},
  {32'hc338b6b7, 32'h42b5c6a7, 32'hc3a703f7},
  {32'h450040d6, 32'hc2f046be, 32'h431064f5},
  {32'hc4f6bd08, 32'h438f149a, 32'h42a1388b},
  {32'h44ecdc52, 32'h422b4cad, 32'hc24e83a4},
  {32'h420bc48a, 32'hc3c800f1, 32'h430e47d8},
  {32'h43b40b6c, 32'h43607007, 32'hc3412d8e},
  {32'h42350740, 32'h41dbadb0, 32'h4309b1eb},
  {32'h44d6d90c, 32'h41b37e7e, 32'hc3bdfdcc},
  {32'hc455ecc8, 32'h433ba459, 32'h442e2d78},
  {32'h4461da15, 32'h4375191c, 32'hc385be4c},
  {32'hc488a1b4, 32'h42194d62, 32'hc40e00ba},
  {32'h4461cb36, 32'h42e7d0d3, 32'h437703ac},
  {32'hc4cbe0cf, 32'hc24b257f, 32'hc0875b37},
  {32'h450c832a, 32'h42ddc54c, 32'hc0109e8e},
  {32'hc4ffc7a5, 32'hbfdbb450, 32'h4329f783},
  {32'h44d1cf18, 32'h42957268, 32'hc30d70e6},
  {32'hc3b7a2ea, 32'hc3099c76, 32'hc34d0f7f},
  {32'h44d134f7, 32'h438736a5, 32'hc2485792},
  {32'hc519630c, 32'h424cbdd4, 32'h41301e63},
  {32'h45152b04, 32'hc32925b5, 32'hc30ef2db},
  {32'hc4902f93, 32'h430dde99, 32'hc2915d4c},
  {32'h450c1044, 32'h42f0c67d, 32'hc2e7de47},
  {32'hc427da6c, 32'hc2b2e949, 32'hc337e266},
  {32'h451ed275, 32'hc25ff78f, 32'hc3ef7123},
  {32'hc4f917db, 32'h43864c41, 32'hc2b22005},
  {32'h4383a440, 32'hc2e8db7e, 32'hc30ada58},
  {32'hc2a3ce44, 32'hc27f9e6d, 32'hc18956cd},
  {32'h44241d78, 32'hc34cee53, 32'h41d655bc},
  {32'hc48595c6, 32'h4183ff92, 32'h436d2015},
  {32'h44cb8c89, 32'hc3472dd4, 32'hc232caa2},
  {32'hc4b9752b, 32'hc36b0b2e, 32'hc3b3471e},
  {32'h43c141b2, 32'h43925c0f, 32'hc36a594d},
  {32'hc4f4c25b, 32'h4240d9d2, 32'hc1d0be58},
  {32'h4389dcf0, 32'hc2fd7d6c, 32'h430bb193},
  {32'hc39cbc78, 32'hc28dbf7a, 32'h42c990cf},
  {32'h43c44149, 32'h43cc629d, 32'hc3375a8d},
  {32'hc430aae7, 32'h42a1de15, 32'h43de067e},
  {32'h44ce5b40, 32'h42af9dee, 32'hc3aaa3ff},
  {32'hc4f9fdb8, 32'hc30a6eee, 32'hc31a19d1},
  {32'h43bc717a, 32'h41e22a67, 32'h43c6d492},
  {32'hc4f15d2a, 32'hc33eaad5, 32'h43284e06},
  {32'h44f4688c, 32'h43ab0356, 32'h422fcaf1},
  {32'hc432a954, 32'h43e08946, 32'h42f03d74},
  {32'h447aa2d6, 32'hc34d409b, 32'hc3bd01c8},
  {32'hc4a5de04, 32'h42cfcdc2, 32'h404237e0},
  {32'h44b94452, 32'hc2a25393, 32'hc1e95aa8},
  {32'hc4af60d9, 32'hc221292f, 32'hc3a223e6},
  {32'h4406256f, 32'hc33ecdc1, 32'hc2abc6ec},
  {32'hc4191a98, 32'h43cd2669, 32'hc32196f2},
  {32'h44a0af9e, 32'h433c9134, 32'h43639084},
  {32'hc4bba7ee, 32'h4187091b, 32'hc26012c3},
  {32'h43ba4704, 32'h4391210c, 32'h43c4cbf3},
  {32'hc46177ff, 32'hc296ca92, 32'hc2a99658},
  {32'h4506ceca, 32'hc218908d, 32'hc37638b4},
  {32'hc435b05a, 32'h43c744ea, 32'h433e4bd2},
  {32'h44dad68c, 32'hc3244e7e, 32'h42de9fb5},
  {32'hc4c79424, 32'h43107a3e, 32'hc31ff8d8},
  {32'h44de23e9, 32'h4341562f, 32'h43b45207},
  {32'hc12c6d4c, 32'hc2a1861e, 32'h42bb43c1},
  {32'h438e0c3d, 32'h42224b73, 32'h436e8c5a},
  {32'hc495f3fc, 32'hc3110e5c, 32'hc3bd3103},
  {32'h44b5b690, 32'hc3872af6, 32'hc25b92a0},
  {32'hc4999c61, 32'h43961e50, 32'hc3655b24},
  {32'h44b8b877, 32'h40c25b2d, 32'hc25a8930},
  {32'hc325f2d6, 32'hc308d5f1, 32'hc1a1f4dd},
  {32'h446c0f14, 32'hc354a67f, 32'h432511d0},
  {32'hc2a0d736, 32'hc2efa085, 32'h4283edf5},
  {32'h445019e0, 32'hc3f7a0d8, 32'h43c347cd},
  {32'hc45929e0, 32'hc31751bd, 32'h4316dea2},
  {32'h45069778, 32'hc38639a4, 32'hc3772cb0},
  {32'hc4ae4913, 32'hc2bc90f1, 32'hc127a38a},
  {32'h44ca9e3c, 32'hc3965871, 32'h4341f536},
  {32'hc4ef80ef, 32'h443543e3, 32'hc3607c28},
  {32'h4508ef08, 32'hc3c5b074, 32'h4326d16f},
  {32'h423e29c0, 32'hc3731d0b, 32'hc399ed94},
  {32'h446b80b2, 32'h42b120c4, 32'h43a43fee},
  {32'hc490f6cf, 32'hc245fe7c, 32'h43816193},
  {32'hc394bfa8, 32'hc3a7d546, 32'h4247038e},
  {32'hc4d13ae8, 32'h4382c897, 32'h42665f22},
  {32'h4454b310, 32'h4302b9d8, 32'hc2c1774e},
  {32'hc4c824af, 32'hc2e387d3, 32'hc231dade},
  {32'h43ab8fd0, 32'h4306b39f, 32'h43c86956},
  {32'hc4ed4dd6, 32'h435ace7a, 32'h4340d34d},
  {32'h44d30a4b, 32'h4211fb42, 32'hc2c05bc5},
  {32'hc452f358, 32'hc3714293, 32'hc34df074},
  {32'h448003cb, 32'hc3139eb5, 32'h42b12a05},
  {32'hc50ce130, 32'hc2be34b0, 32'hc2543ec0},
  {32'h449347c5, 32'h42897e7e, 32'hc301a67f},
  {32'hc50c66e2, 32'hc17eefbd, 32'h42a465b3},
  {32'h45002a8a, 32'h437bc226, 32'hc308a4c1},
  {32'hc514d818, 32'hc29b6532, 32'h429b1fd6},
  {32'h446e95d6, 32'h4193c0a9, 32'hc300c2d7},
  {32'hc36bff7e, 32'h43ef293a, 32'h43b09448},
  {32'h44bb819c, 32'h42dfa9aa, 32'hc34f59d6},
  {32'hc4a82c9e, 32'hc4200e1e, 32'h43a8d190},
  {32'h449928fa, 32'h43e88d7d, 32'hc25015bf},
  {32'hc4aabbe4, 32'h43b991e8, 32'h43e0daed},
  {32'h449374a4, 32'hc32b2ff2, 32'hc223edc2},
  {32'hc2273dc3, 32'h42ff7462, 32'hc3f49077},
  {32'h44c3d28e, 32'h42bb5251, 32'hc2a6cb1c},
  {32'hc3d08a3c, 32'h432e2cf4, 32'hc25a98f2},
  {32'h436a7270, 32'hc303a3a9, 32'h439292ec},
  {32'hc40de20c, 32'hc293d9b6, 32'hc2809203},
  {32'h4502a99e, 32'h437637de, 32'h43932a72},
  {32'hc4c2d1a2, 32'hc146be0c, 32'hc386e67b},
  {32'h44849b31, 32'h436b8e07, 32'hc14c4909},
  {32'hc4bcd859, 32'hc292180b, 32'h43f1c056},
  {32'h4491c62c, 32'hc2e632f6, 32'hc3a5a34b},
  {32'hc4923e75, 32'h4277870c, 32'h43ba99aa},
  {32'h44ccfd6f, 32'h42b7d12a, 32'h43950e7d},
  {32'hc4d46160, 32'hbf82aec5, 32'hc2de30ba},
  {32'h43b936b4, 32'h43ac9769, 32'h43452146},
  {32'hc4e2f367, 32'h4387def1, 32'h4303b1ea},
  {32'h44ef472a, 32'hc36f9409, 32'h428ca2f6},
  {32'hc50f3b07, 32'hc3571b30, 32'h433a6188},
  {32'h43e18676, 32'h4391ccaa, 32'hc2257c05},
  {32'hc4650722, 32'hc31d69ef, 32'hc288296d},
  {32'h44e9bba2, 32'h434f7b59, 32'hc36232af},
  {32'hc35cc7c0, 32'hc3eb5cfa, 32'h43780829},
  {32'h44b87700, 32'h43782b46, 32'hc2ce4a1b},
  {32'hc4853ac2, 32'hc3bf9656, 32'h428246e7},
  {32'h4403fade, 32'hc3795053, 32'h436f4733},
  {32'hc4eee996, 32'hc3b5cdaf, 32'hc3195cba},
  {32'h448b7460, 32'h43b489ca, 32'h4240f5d3},
  {32'hc322421b, 32'h439ac343, 32'hc32620d0},
  {32'h432b208c, 32'hc37ab647, 32'h4354867d},
  {32'hc5022e71, 32'hc29902d4, 32'h43545e3e},
  {32'h4504717a, 32'h4330e0ba, 32'h42097873},
  {32'hc341ede0, 32'h4242d2e8, 32'hc157805a},
  {32'h44585ad2, 32'hc2217af7, 32'h41ef85c0},
  {32'hc4bf02d8, 32'h42025c3d, 32'hc34abed1},
  {32'h44bf3fef, 32'h433a5611, 32'h431f2a48},
  {32'hc43126f0, 32'hc39df841, 32'hc2c00878},
  {32'h45026879, 32'h43729cbf, 32'hc382a437},
  {32'hc44a4016, 32'h43006cc4, 32'hc39366e8},
  {32'h450aea96, 32'h43578bc1, 32'h41b51015},
  {32'hc4ac2ea6, 32'h429e8a8f, 32'h4336b61a},
  {32'h44bfa78e, 32'h43258191, 32'h425e4917},
  {32'hc4e1cc8d, 32'h427e6ce2, 32'hc2f19175},
  {32'h4473859c, 32'h434bf4e1, 32'h42184b45},
  {32'h436e8893, 32'hc3b27d98, 32'hc41ca417},
  {32'h44ddb36e, 32'h42d5d2db, 32'hc1febc1c},
  {32'hc4ed3616, 32'h4309bf16, 32'hc37d098c},
  {32'h43a8f754, 32'hc32b6715, 32'hc391f63e},
  {32'hc4af71f4, 32'h4324179a, 32'hc394cf37},
  {32'h45025158, 32'h44338af0, 32'h4286ef02},
  {32'hc48e2195, 32'h431fe909, 32'hc21647e5},
  {32'h430aaf83, 32'h433bc114, 32'h43b5613d},
  {32'hc4360306, 32'hc2debd4e, 32'hc2aa712a},
  {32'h44cfd597, 32'hc2f3fa18, 32'hc3854fb6},
  {32'hc51b9e80, 32'h4162d955, 32'hc305d553},
  {32'h4498b4be, 32'h42691e78, 32'h43fe843e},
  {32'hc46c1c2e, 32'h43e7d62b, 32'h42e95601},
  {32'h4396c9f8, 32'hc2340cbb, 32'hc37658d6},
  {32'hc475c072, 32'h429f6781, 32'h4296fe7b},
  {32'h440ed637, 32'hc3072607, 32'h42111686},
  {32'hc4839d3c, 32'hc3d10bd6, 32'hc3d48c26},
  {32'h441fe102, 32'hc2a04049, 32'hc339adfb},
  {32'hc4c143fa, 32'h42d227d4, 32'h42f59a4d},
  {32'h44df4657, 32'hc2345f67, 32'h434f58f7},
  {32'h436b01b0, 32'h438d5dd2, 32'h3f426320},
  {32'h449d8df9, 32'h43221be9, 32'h42598814},
  {32'h4208a900, 32'h439f34b3, 32'h43bfbc1c},
  {32'h44f1b19b, 32'hc3153a76, 32'hc20926dc},
  {32'hc5202e7a, 32'h42a15918, 32'h43fd1904},
  {32'h4486701c, 32'h426b7f1a, 32'h43769359},
  {32'hc3822e38, 32'h41d0a2e8, 32'h41642184},
  {32'h44fbda84, 32'h43c2b103, 32'hc3505919},
  {32'hc514654c, 32'hc2bc26d9, 32'hc3bb80f2},
  {32'h43184960, 32'h3fd37af6, 32'hc338a3e1},
  {32'hc4398d33, 32'h42e39e89, 32'hc3241c3b},
  {32'h430e26f0, 32'h41f9f29a, 32'hc34af593},
  {32'hc3665612, 32'h43630291, 32'h42deca8f},
  {32'h448effbb, 32'h42732d62, 32'hc3896292},
  {32'hc3bcce84, 32'h4358cd9b, 32'h41fb2c0e},
  {32'h440caabc, 32'h43293bc3, 32'h438a8bb2},
  {32'hc5039a7e, 32'hc1455bb4, 32'h43688ab7},
  {32'h4499bbf2, 32'hc2a9aa39, 32'h43031f71},
  {32'hc496d4cf, 32'h41ff781b, 32'h42ef4042},
  {32'h44d97948, 32'hc39587b2, 32'h43920d06},
  {32'hc2826220, 32'hc37619ce, 32'hc29d33b4},
  {32'h44acf952, 32'h431b42b6, 32'h43c0a5c5},
  {32'hc23cdd90, 32'h43ca1931, 32'h43cf45ff},
  {32'h44675aba, 32'h42ef24ed, 32'h41c31418},
  {32'hc4aabd70, 32'hc1c30a42, 32'h40d7b9c0},
  {32'h44e55e69, 32'hc1d8fd24, 32'h42bcc70d},
  {32'hc43b6c92, 32'h42f7be92, 32'hc2ecac85},
  {32'h440b31f8, 32'hc3aa9e2b, 32'h43c99532},
  {32'hc500f2ca, 32'h43d0221a, 32'hc33af0cd},
  {32'h4504481a, 32'h42fafb87, 32'hc2ce59b0},
  {32'h436e447a, 32'hc3190eb9, 32'h429171fa},
  {32'h443788f2, 32'h3f876118, 32'h4174ca80},
  {32'hc4a02354, 32'hc337a32c, 32'h424ff80e},
  {32'h44fe1c66, 32'hc3520a61, 32'hc2e25d22},
  {32'hc505c311, 32'hc36f5a12, 32'h4317726e},
  {32'h44cce57a, 32'h431353ae, 32'h42e13a85},
  {32'hc3d9b84e, 32'h430359b5, 32'hc3b9aa88},
  {32'h45311fdc, 32'h43a8252d, 32'h409e2432},
  {32'hc4565471, 32'hc2a5d762, 32'hc29ccf3a},
  {32'h447f482e, 32'hc285117f, 32'hc21572fa},
  {32'hc4809497, 32'h431f2913, 32'hc37edbd7},
  {32'h451b3cf6, 32'h4274edcf, 32'hc2d6d52c},
  {32'hc525baf1, 32'h437d37d6, 32'h438390c1},
  {32'h444f34a4, 32'hc3a8bc66, 32'hc19675db},
  {32'hc5065ee9, 32'h4286ec81, 32'h43afc642},
  {32'h44dfe1ac, 32'hc3f61f61, 32'h42c86878},
  {32'hc5026281, 32'hc3a613ff, 32'hc39dbeb8},
  {32'h444c42f0, 32'hc3ccde40, 32'hc37b4a11},
  {32'hc4591c91, 32'h43476457, 32'hc2b98e28},
  {32'h441eff56, 32'h42bdac12, 32'hc2dcf67b},
  {32'hc5055e58, 32'hc2a80602, 32'h43335774},
  {32'h44b95cb5, 32'hc290df29, 32'hc2d89a65},
  {32'hc4322203, 32'hc3844cf9, 32'hc3800c9f},
  {32'h4520004c, 32'h4368645a, 32'hc3cba1d3},
  {32'hc500bf18, 32'hc0c95f96, 32'hc2e1d225},
  {32'h4479d37e, 32'hc3ac1b25, 32'hc136751b},
  {32'hc48618ca, 32'hc300324d, 32'h43fc78de},
  {32'h44d87c5c, 32'h42a91bca, 32'h41cf4534},
  {32'hc3281b18, 32'h435e7b31, 32'h4389c777},
  {32'hc25d2a74, 32'hc3b9e690, 32'h418d49ab},
  {32'hc40c741d, 32'hc165cb8f, 32'hc3a80a1d},
  {32'h447d75f2, 32'hc31ccfea, 32'h421826f9},
  {32'hc50427fa, 32'h434f60a4, 32'h43a8f4a4},
  {32'hc29c0190, 32'hc34636f0, 32'hc26e0dea},
  {32'hc51751d5, 32'h420be28b, 32'hc1c70683},
  {32'h44f725e8, 32'h420bf04d, 32'h432a1cff},
  {32'hc5027c22, 32'hc31b7ad6, 32'hc327ef5b},
  {32'h44fd7ab4, 32'h4254f156, 32'h4263b9c1},
  {32'hc3f04dee, 32'hc1a5e7ce, 32'hc34d52c1},
  {32'h442a6806, 32'hc0c68fe1, 32'h42b90eea},
  {32'hc46b5041, 32'h430426c6, 32'hc322a2cd},
  {32'h435227ac, 32'h4288cd09, 32'hc213c03d},
  {32'hc513ee13, 32'hc3468406, 32'hc0f3a67b},
  {32'h441a711b, 32'h434df489, 32'hc2e55cc7},
  {32'hc4cd3c66, 32'hc3b7e77f, 32'hc30b5b2d},
  {32'h45147be8, 32'hc2c0b482, 32'h4318ce91},
  {32'hc2b15a64, 32'hc36f1591, 32'h43cd2767},
  {32'h44d79b03, 32'hc3886df8, 32'h4307b964},
  {32'hc3d957d0, 32'h3f68687c, 32'hc38c0a80},
  {32'h450d7aff, 32'h42cac1e9, 32'hc1d21cb9},
  {32'hc3cf33d4, 32'h42803841, 32'h41bf3fbd},
  {32'h4509fce4, 32'h43907439, 32'h432d4683},
  {32'hc4c45089, 32'h41ae33c3, 32'h43031b83},
  {32'h44a40608, 32'h4302ae58, 32'hc230c72b},
  {32'hc50a9be0, 32'hc3a1fc2b, 32'h42d91d78},
  {32'h44c72da5, 32'h419dd4db, 32'h44031982},
  {32'hc4ad27f2, 32'h4284d156, 32'hc3249724},
  {32'h45096378, 32'hc31a726e, 32'hc3c2f300},
  {32'hc5052547, 32'hc338f7ed, 32'h431d33cf},
  {32'h44415a8c, 32'h4340c980, 32'hc29580f3},
  {32'hc4017422, 32'hc3450fbb, 32'hc3b2c59f},
  {32'h44609598, 32'hc35419f6, 32'hc2827c9d},
  {32'hc4e72743, 32'h4208f4ea, 32'hc34bc1ed},
  {32'h450463e4, 32'h43c71d69, 32'hc2849226},
  {32'hc48e3e27, 32'hc2baf156, 32'h4400e6d6},
  {32'h44afe7ad, 32'hc30e7bfd, 32'hc3a8187f},
  {32'hc32a59a8, 32'hc28fa464, 32'hc29f5242},
  {32'h4493a83a, 32'h435822ae, 32'hc379ff7c},
  {32'hc422b9da, 32'h438ecbc2, 32'hc2cdf1d4},
  {32'h450d1152, 32'h436ad5f4, 32'hc1833527},
  {32'hc4914a6c, 32'h43398e9c, 32'hc329dc75},
  {32'h445f6c7c, 32'hc3507027, 32'hc2ee03e4},
  {32'hc4c45184, 32'hc1c38cc8, 32'hc32833a0},
  {32'h43a05334, 32'hc2acd4c4, 32'hc2df505a},
  {32'hc4493c06, 32'hc2aaa301, 32'hc086e450},
  {32'h44f7b0ad, 32'hc305c661, 32'hc3930691},
  {32'hc2cf23f0, 32'hc35bd5a2, 32'h436d0247},
  {32'h44a26d3f, 32'h4318a8b2, 32'hc381ea79},
  {32'hc1d429e4, 32'hc2bf2e28, 32'h4388e00f},
  {32'h44cc0bf1, 32'h433f728e, 32'h430ecd1b},
  {32'hc48b46e0, 32'h421f165a, 32'h438a1653},
  {32'h42ab6760, 32'h43486a50, 32'hc3344dc2},
  {32'hc4a7d370, 32'h43d2d802, 32'hc269bdb0},
  {32'h44d45355, 32'hc1c2644b, 32'hc398e887},
  {32'hc4ea4c52, 32'h432a6584, 32'h438bd5c4},
  {32'h4513cb8f, 32'hc1f2b536, 32'hc31bc0e3},
  {32'hc0f0f600, 32'h43328418, 32'h41adb888},
  {32'h4451a3df, 32'h439d90e2, 32'hc393e8ea},
  {32'hc5098c55, 32'hc405e4ea, 32'hc38dfa98},
  {32'h438dad08, 32'hc32ed05a, 32'hc38f3878},
  {32'hc4f0f987, 32'h428c1e48, 32'h430caa39},
  {32'h442bdea2, 32'hc1cf43e2, 32'hc1851c9c},
  {32'h43583da0, 32'h43f1f7f1, 32'hc307cc07},
  {32'h4492453e, 32'h4388d977, 32'h430dc553},
  {32'hc4cbe97a, 32'h42c2ce79, 32'h42fbf5b1},
  {32'h44b81a76, 32'h4345a9cf, 32'hc36195a8},
  {32'hc4136d75, 32'h4364bdb4, 32'h41c077a5},
  {32'h44638f88, 32'h406ecabf, 32'hc3629ee8},
  {32'hc4b7a8d9, 32'h4214f8ee, 32'h43a9ab04},
  {32'h44879c53, 32'hc2a55fce, 32'hc3e32bda},
  {32'hc50c0a14, 32'h4336e608, 32'h4389babf},
  {32'h442412d4, 32'h43400e1d, 32'hc1b068fc},
  {32'hc4e1efec, 32'hc2ceac39, 32'h42d60852},
  {32'h44b06e0d, 32'h42a56014, 32'hc1cf19ee},
  {32'hc4d1e2e0, 32'h43a53a8b, 32'hc2c4ecad},
  {32'h448c7fb1, 32'hc3f246c6, 32'hc41db530},
  {32'hc4cc5a46, 32'hc24fbd8c, 32'h438ea5ef},
  {32'h44bcd522, 32'h43047b3b, 32'hc3050eff},
  {32'h44c631c3, 32'h43568224, 32'hc2a8a1f3},
  {32'hc3d68429, 32'hc2d27cf2, 32'h434c0d47},
  {32'h44dd3eac, 32'hc3c407a6, 32'h43bdaf42},
  {32'hc408bbd6, 32'h42643e8b, 32'hc29ab553},
  {32'h448d87ca, 32'hc2bb4d52, 32'hc31ff7ce},
  {32'hc4ade09d, 32'h42efb1dd, 32'hc27cd24a},
  {32'h44f96c9c, 32'hc2f9de01, 32'hc2c91119},
  {32'hc4417eb6, 32'hc2f16003, 32'h4165e6ca},
  {32'h44ee80b2, 32'hc1ebb078, 32'h41cfcb79},
  {32'hc355f080, 32'hc2ea19a4, 32'h41e690ac},
  {32'h44af03a7, 32'h434cab57, 32'hc2f58a18},
  {32'hc44df432, 32'h41d59c4e, 32'h43a0fa2b},
  {32'h44925563, 32'hc3089f8a, 32'hc2a93a9f},
  {32'hc484f6c5, 32'h437d1ebb, 32'hc277fd59},
  {32'h43c2d614, 32'hc397e1cc, 32'hc2b9fec0},
  {32'h40d0bc00, 32'hc37acdbf, 32'h440f82ca},
  {32'h44bab7a3, 32'h42b88ab0, 32'hc226a196},
  {32'hc46fa5df, 32'hc38cdbb3, 32'h43771f69},
  {32'h44aca8b5, 32'h43dc70a3, 32'hc380b66e},
  {32'hc518b2d3, 32'h432fe903, 32'hc3946927},
  {32'h44dfc016, 32'hc349e205, 32'h42bb6feb},
  {32'hc5221b95, 32'h439e88e5, 32'h42bdb437},
  {32'h43b2753a, 32'h407b0e13, 32'hc3868da8},
  {32'hc49bf3a5, 32'hc154434e, 32'hc2826c0a},
  {32'h44fb3072, 32'h42746f48, 32'hc34f17b6},
  {32'hc4b17d74, 32'h43034c40, 32'h4341d252},
  {32'h44b59fd7, 32'h439d5b22, 32'hc3284e6c},
  {32'hc3aad377, 32'h4230e3ae, 32'h41f887ee},
  {32'h445997ef, 32'h43529c3b, 32'h431cda88},
  {32'hc324a8e0, 32'hc3445a96, 32'hc24cea06},
  {32'h43e4ade1, 32'hc29cdc4e, 32'hc2a51528},
  {32'hc47ac2ae, 32'hbf8a6bfa, 32'hc2edc47d},
  {32'h44ef3dfa, 32'h42f67999, 32'h43b1382c},
  {32'hc4cd2171, 32'h4181bb7e, 32'hc35a8f14},
  {32'h44de73a8, 32'hc1e418ff, 32'hc2c13211},
  {32'hc512bfab, 32'hc2b825f2, 32'h4306e1ea},
  {32'h44b46fbb, 32'h42c39f94, 32'hc405f026},
  {32'hc3ca9548, 32'hc3839a73, 32'h41f6d170},
  {32'h4433d8b4, 32'hc3dabb56, 32'h41b10f75},
  {32'hc4e047f2, 32'h4344e326, 32'hc38e4d35},
  {32'h44cccb10, 32'hc29da49f, 32'h43885930},
  {32'hc4ebf978, 32'h4276ee79, 32'h42639109},
  {32'h439f1028, 32'hc401f4f0, 32'h42cbd5dd},
  {32'hc4a41689, 32'hc3695570, 32'h4346f5a2},
  {32'h447f9036, 32'h429e810c, 32'h437c982a},
  {32'hc4e44788, 32'h42197af6, 32'hbfa08750},
  {32'h45138327, 32'h42873d99, 32'h43206e9c},
  {32'hc4c6685d, 32'h43c86a9c, 32'hc3be9fd5},
  {32'h446d5c5a, 32'h442b2255, 32'hc38f7cb6},
  {32'hc4a5950c, 32'h43267b2c, 32'hc2858e8d},
  {32'h453156d6, 32'hc31f2fc7, 32'h4311bf09},
  {32'hc4d66867, 32'hc27c698d, 32'hc35b3285},
  {32'h44e74ce2, 32'hc2a053b6, 32'hc27d1a66},
  {32'hc50037a7, 32'h4292628a, 32'h42964532},
  {32'h43f6c080, 32'hc35123e5, 32'hc2fe1e9a},
  {32'hc3b094fe, 32'h4353e91f, 32'hc400afb7},
  {32'h44a120af, 32'h41dac96d, 32'hc3589fe9},
  {32'hc5098760, 32'h4407d01c, 32'hc4345d1d},
  {32'h44d864af, 32'hc32249e7, 32'h434140a9},
  {32'hc3851c06, 32'hc384f862, 32'hc1894797},
  {32'h450a0631, 32'hc3531315, 32'h44098749},
  {32'hc41bf732, 32'h43730185, 32'h42c945b8},
  {32'h44ff203b, 32'hc38c799e, 32'hc22718e2},
  {32'hc51d7e61, 32'h42853201, 32'h431884e5},
  {32'h42f7b020, 32'h42723426, 32'h43820380},
  {32'hc4c247c6, 32'h43d34233, 32'hc2cabc35},
  {32'h443985ac, 32'h43784783, 32'hc384e8ca},
  {32'hc4bad055, 32'hc39fddc8, 32'hc2a8f8d6},
  {32'h4502726a, 32'h43ac3d8d, 32'hc20ac0fb},
  {32'hc4ccbe48, 32'h42af8642, 32'h4189a71f},
  {32'h452233d9, 32'hc034b656, 32'h43272265},
  {32'hc4897cca, 32'h41754859, 32'h404b8a80},
  {32'h44f90c8d, 32'h4302b491, 32'h430a7407},
  {32'hc41ee0a0, 32'hc2145271, 32'hc350759b},
  {32'h45030f5c, 32'hc40dd050, 32'hc38bf4ae},
  {32'hc38b81fd, 32'h426af204, 32'h434a9808},
  {32'h4433e072, 32'hc35d63bd, 32'hc38c4e14},
  {32'hc4e03d43, 32'h4313c071, 32'h4232717d},
  {32'h44a7fbe9, 32'hc239c213, 32'h426c6c82},
  {32'hc4ebe0f1, 32'h430cd295, 32'hc19faa10},
  {32'h43b5f0e0, 32'hc32accb3, 32'hc2a36efb},
  {32'hc3f6d87c, 32'h41f2eb8e, 32'h42a37315},
  {32'h446b4a74, 32'h427bb1a1, 32'h43851e6d},
  {32'hc4e01087, 32'hc395b03a, 32'hc17dbbda},
  {32'h44c687c8, 32'hc0285820, 32'h43683482},
  {32'hc510a2a9, 32'h405f5a90, 32'hc30443e9},
  {32'h438040d4, 32'h43e6ef95, 32'h42ebd234},
  {32'hc39b8020, 32'hc3be61f9, 32'h43efcfba},
  {32'h43d0e678, 32'hc36e6769, 32'h43ac919c},
  {32'hc39f8349, 32'h4350843d, 32'hc38a6e3c},
  {32'h438f3b64, 32'h430fbbe1, 32'h4262ba90},
  {32'hc44d6f31, 32'h4350b9f8, 32'h43171ed5},
  {32'h45163c0d, 32'hc201529a, 32'h438e3cb5},
  {32'hc49711ab, 32'h41f900e6, 32'hc3604722},
  {32'h4503b7f2, 32'h43fb24e1, 32'hc31312a7},
  {32'hc479e105, 32'h41d27bf9, 32'hc32a0b54},
  {32'h44fd5fcd, 32'h4323d39d, 32'hc36305c8},
  {32'hc470f2d1, 32'hc306b2c8, 32'hc3412513},
  {32'h44860034, 32'hc3b6ef8d, 32'h413deef9},
  {32'hc48f0cc2, 32'hc38d12df, 32'h435041c9},
  {32'h45124ad1, 32'h430c9409, 32'h43471869},
  {32'hc3d679f7, 32'h43c749e8, 32'hc2b6e26f},
  {32'h43c6cfd6, 32'h430c32eb, 32'h43ce4e57},
  {32'hc409cbed, 32'h4383d323, 32'h43e8672f},
  {32'h4406d178, 32'hc37999dd, 32'hc22b04e0},
  {32'hc4af4025, 32'h43399c30, 32'hc3018f7b},
  {32'h451ba990, 32'h43c69970, 32'hc22c09d7},
  {32'hc4b96d20, 32'hc2ce613f, 32'hc194f1da},
  {32'h44391686, 32'hc303c55b, 32'hc2fef36d},
  {32'hc31e19e7, 32'hc39d2c4f, 32'h43a3d586},
  {32'h44f4ef55, 32'hc30bee10, 32'h428c5f78},
  {32'hc3c76c47, 32'hc2a6694e, 32'h43044160},
  {32'h4401a3d6, 32'hc340cd3c, 32'hc31aee40},
  {32'hc4da5516, 32'hc3027f36, 32'h42914665},
  {32'h44832d2c, 32'h431d677a, 32'h4387221a},
  {32'hc42d1886, 32'h434452ca, 32'hc32e3114},
  {32'h45160e35, 32'hc335db8c, 32'h421e2040},
  {32'hc4d06dd3, 32'h4381a3c7, 32'h42847fba},
  {32'h44380521, 32'hc1d07f56, 32'h425803e3},
  {32'hc4098700, 32'h4297a503, 32'h42c43f1a},
  {32'h44dc317a, 32'h43ba8603, 32'hc357177e},
  {32'hc50c546a, 32'hc331f88e, 32'h430cf41a},
  {32'hc3251d70, 32'h424281e1, 32'h4246491a},
  {32'hc49ff4e8, 32'hc2b1ac64, 32'h42be4ac3},
  {32'h447748e4, 32'hc34ec536, 32'hc393f266},
  {32'hc4c557bc, 32'h422d91df, 32'hc308b6b3},
  {32'h41f46580, 32'hc331efbb, 32'hc3b85da4},
  {32'hc5045995, 32'h422cea90, 32'h4340d2b5},
  {32'h44ef447c, 32'hc238f0b8, 32'h4291cf9e},
  {32'hc4f70c58, 32'hc38571e0, 32'h43863cea},
  {32'h448c5f7f, 32'h4295f65b, 32'h4315c7ac},
  {32'hc4399018, 32'hc371f14f, 32'h43009702},
  {32'h44617660, 32'h43e61a6b, 32'hc1dedaef},
  {32'hc3cfb242, 32'h437172ec, 32'hc2d43e70},
  {32'h43c99d2a, 32'hc2b92d8d, 32'hc2c3637b},
  {32'hc4f2be35, 32'h422d6f56, 32'h415c3ec2},
  {32'h44e90732, 32'h42de101e, 32'h43a10c37},
  {32'hc5006232, 32'h42086102, 32'h43d4f15f},
  {32'h4386f615, 32'hc3502603, 32'hc29b46e3},
  {32'hc4cb6e67, 32'hc37f8933, 32'hc3637dfe},
  {32'h44c1252d, 32'h432d94f7, 32'hc3a020ca},
  {32'hc2556d80, 32'hc3d33b28, 32'h4387546f},
  {32'h450c9ded, 32'hc29f2f1c, 32'hc3e6c79a},
  {32'hc3f8dcd6, 32'hc2662757, 32'h43f42585},
  {32'h43b69270, 32'h42aa2fb0, 32'h43d6e452},
  {32'hc3eba130, 32'h41ddf02f, 32'hc30953ae},
  {32'h438f43fc, 32'hc378343f, 32'hc397d82f},
  {32'hc4937423, 32'h431d473b, 32'h431c910a},
  {32'h44f7ea4c, 32'h40c7c802, 32'h41815d54},
  {32'hc40cc541, 32'h439feba6, 32'hc2a11312},
  {32'h448856e8, 32'h43904e7d, 32'hc3a91cd3},
  {32'hc48892c9, 32'hc34df9b7, 32'hc21aee63},
  {32'h43f13af4, 32'h43003285, 32'hc357bfe3},
  {32'hc4cf4fef, 32'h41885f8a, 32'hc3f1bc79},
  {32'h4504d435, 32'h4332446b, 32'hc258da6d},
  {32'hc51248c6, 32'h43a5e29d, 32'h4283dc75},
  {32'h45016467, 32'hc4244f57, 32'hc36001ea},
  {32'hc293f872, 32'hc3abe103, 32'h4351c1bb},
  {32'h441a19bf, 32'h4301b9fe, 32'hc2035087},
  {32'hc4540532, 32'hc3a838ed, 32'h4385dc83},
  {32'h44461f23, 32'hc35ee6ec, 32'h42e8c793},
  {32'hc5043bb2, 32'hc36cc4cc, 32'h42335b33},
  {32'h439f4c72, 32'hc2e0df8d, 32'h435935a7},
  {32'hc46d67e2, 32'hc293a052, 32'h434ac375},
  {32'h44aa1a2c, 32'hc375a553, 32'hc2010afb},
  {32'h42e32590, 32'hc13dff8f, 32'hc3bd6898},
  {32'h44803963, 32'hc358ff45, 32'h439131eb},
  {32'hc4d13fe9, 32'hc20cb1de, 32'hc32ca987},
  {32'h44beb2f0, 32'hc3e38651, 32'h427dc048},
  {32'hc4bfb083, 32'hc30220bf, 32'hc289cc5e},
  {32'h44f63282, 32'hc17935b0, 32'hc2f46fbb},
  {32'hc49fc572, 32'hc2f0742f, 32'h432af6ce},
  {32'h44f9dc5c, 32'hc3e6d04c, 32'h4366323c},
  {32'hc41257ea, 32'h42beaa2f, 32'hc3072d64},
  {32'h4505546b, 32'h43fe6af0, 32'h42eefe03},
  {32'hc4bd084e, 32'hc2edbf2b, 32'hc32190fa},
  {32'hc2304060, 32'h42c55038, 32'h43003216},
  {32'hc4bc6159, 32'h432cef88, 32'h435bdab1},
  {32'h45134a4c, 32'hc35bf817, 32'hc31b5927},
  {32'h41f73100, 32'h43b0e100, 32'hc321e055},
  {32'h44097c75, 32'h42b80c1c, 32'hc3d31f0c},
  {32'hc4f106a6, 32'hc38eadd3, 32'hc3f09b82},
  {32'h450688ef, 32'hc366c8de, 32'hbe900d80},
  {32'hc30befe0, 32'hc31a85ff, 32'hc2f77044},
  {32'h44df5d68, 32'hc39fff4d, 32'h438f1386},
  {32'hc4d28b70, 32'h435e8029, 32'h42b42f4c},
  {32'h43ee77c4, 32'h4288cfe0, 32'h43173efe},
  {32'hc48b7d53, 32'h4356e861, 32'hc39a41ba},
  {32'h44fbf3b9, 32'hc3ba6ed3, 32'h42873605},
  {32'h42ca9e62, 32'hc376dd91, 32'h4314cbac},
  {32'h44ff9221, 32'h4139329c, 32'h42bef9ba},
  {32'hc45b8c1c, 32'h4384b94a, 32'hc29d74b5},
  {32'h43c521bc, 32'hc3947887, 32'hc401eab9},
  {32'h413d9c00, 32'hc2c0b00e, 32'hc18ef864},
  {32'h444c58d0, 32'h426bd5b2, 32'h4326865f},
  {32'hc4d8cf83, 32'hc20b14cf, 32'h41e48b12},
  {32'h452ab924, 32'hc402acb3, 32'h432221cd},
  {32'hc4b8bbc6, 32'h4323f6f0, 32'hc08902e5},
  {32'h44fec025, 32'h42662edc, 32'hc32c8932},
  {32'hc4810ab8, 32'h42aa9ebf, 32'hc2f4b383},
  {32'h44e414a4, 32'h4398b9c7, 32'hc3254670},
  {32'hc4d0eea7, 32'hc31bf77b, 32'h430732e2},
  {32'h450b4dfc, 32'hc3b51f53, 32'hc38b7db2},
  {32'hc5124de0, 32'h422c3ce2, 32'hbfa4f38a},
  {32'h44e496fd, 32'hc3ea5247, 32'h42f65337},
  {32'hc4e4b166, 32'h43f229cd, 32'h410d45ca},
  {32'h44d70cf7, 32'hc3cf7c60, 32'h4417939c},
  {32'hc4b5b5d5, 32'h43b9e9c2, 32'h43421099},
  {32'h42280f30, 32'hc15f260b, 32'hc331105a},
  {32'hc4c77f7b, 32'hc36501a7, 32'h43aa34b1},
  {32'h4312d520, 32'h42a6dadd, 32'h43c97d6f},
  {32'hc3d03c3b, 32'hc367c496, 32'h421e8edf},
  {32'h44be4f64, 32'h43ba97b6, 32'h43a6bf7e},
  {32'hc38c2022, 32'hc3ddcae3, 32'h431476b0},
  {32'h449f253f, 32'h431d154b, 32'h432e919f},
  {32'h42cd28d7, 32'h4387968d, 32'h435783cd},
  {32'h4486bc3a, 32'h43975112, 32'hc2c0362e},
  {32'hc4b65fc8, 32'h43255e57, 32'hc3624e92},
  {32'h440b6694, 32'hc30b4192, 32'h43b67964},
  {32'hc2a09f60, 32'hc1a3546c, 32'hc2bb19a0},
  {32'h43fc102f, 32'h43aa7d1d, 32'h43a0acbd},
  {32'hc438f504, 32'hc2590c1d, 32'h43d056eb},
  {32'h43f81518, 32'hc301adb7, 32'h436ec4e1},
  {32'hc51a4fcc, 32'h43a6670f, 32'h43986122},
  {32'h44c310a9, 32'h430f9e17, 32'h42b8d513},
  {32'hc44eb528, 32'h4348c520, 32'hc333c7d3},
  {32'h43a608e8, 32'h43b60500, 32'hc32ee674},
  {32'hc4c5afbc, 32'h416d289c, 32'hc31807e9},
  {32'h437dd593, 32'hc403f8cc, 32'hc196bc3c},
  {32'hc4407429, 32'h427772fe, 32'hc38722f2},
  {32'h447b587f, 32'h436a7323, 32'h432db9d0},
  {32'hc4b84308, 32'hc348bf8b, 32'hc361cdc5},
  {32'h44d09b23, 32'hc3bcb6c8, 32'hc223c9ee},
  {32'hc4e5df65, 32'hc2b2fd2e, 32'h4242bb41},
  {32'h44b891e3, 32'h43fd7ed5, 32'hc3bb4364},
  {32'hc4e003be, 32'hc29d5627, 32'hc327ced9},
  {32'h451383f5, 32'h42839b1d, 32'hc2285425},
  {32'hc509bbed, 32'hc33326fe, 32'hc3954b8b},
  {32'h44ba5370, 32'h42ac15f5, 32'h4378d2cb},
  {32'hc4dc1a2a, 32'hc16c0208, 32'hc3d40299},
  {32'h44ef2bcb, 32'hc2b088fd, 32'h43c81bf8},
  {32'hc45b3562, 32'h42ce3ab3, 32'hc2f241d9},
  {32'h446c8500, 32'hc30bf7a6, 32'hc2a97ceb},
  {32'hc4a74d81, 32'h41cddd64, 32'h43d85420},
  {32'h44bde900, 32'hc32e8cfb, 32'h41ff9723},
  {32'hc4be7f92, 32'hc2250e42, 32'h42955dc0},
  {32'h43bc5f02, 32'h439bcc11, 32'h420ca0c0},
  {32'hc4d37716, 32'hc3cb1403, 32'h421ca1a9},
  {32'h450391b5, 32'h42826f88, 32'h433231c4},
  {32'hc37d6f7c, 32'hc212035d, 32'hc3fb07b0},
  {32'h439057ed, 32'hc2ec779f, 32'hc1204d61},
  {32'hc4d49f62, 32'h4360a711, 32'hc30b924f},
  {32'h44a54fd6, 32'hc37c7aeb, 32'hc3875664},
  {32'hc453c850, 32'hc30eafcb, 32'hbe8a0c24},
  {32'h44832701, 32'h42f193c2, 32'h433d9a3d},
  {32'hc501a03d, 32'hc3a6237d, 32'hc3adcc08},
  {32'h4500d8a8, 32'h43a6d431, 32'hc295e8b5},
  {32'hc4c9f22b, 32'hc28b2c83, 32'h43918925},
  {32'h4458bb72, 32'h42cda8f3, 32'h41cbfc5a},
  {32'hc4c6ed8a, 32'h42ae683e, 32'hc1d0c4a6},
  {32'h44b82911, 32'h41e816bf, 32'hc355ce3e},
  {32'hc506e308, 32'hc4060fd2, 32'h43031466},
  {32'h449e423a, 32'h438add8e, 32'h3f9fc76e},
  {32'hc51ffbf2, 32'h422e8c88, 32'hc2a1aeaf},
  {32'h44073d14, 32'h440e7758, 32'hc42879b3},
  {32'hc4c7bc65, 32'hc2dcabef, 32'h43b28273},
  {32'h4489e58c, 32'hc2697b81, 32'hc404730b},
  {32'hc51cc39a, 32'h4327c92b, 32'hc32276e9},
  {32'h44921522, 32'h432d7c75, 32'hc369fc69},
  {32'hc2ffb3e0, 32'hc3105a95, 32'hc298de40},
  {32'h44ed0c85, 32'h42d14811, 32'hc2e4a973},
  {32'hc4e85a55, 32'hc36e8c08, 32'h433c44bd},
  {32'h44abdbc2, 32'hc36b7288, 32'hc2394c81},
  {32'hc507f20c, 32'hc31ca7ef, 32'hc3e33aea},
  {32'h451e1670, 32'h43619ec7, 32'hc2ce8c45},
  {32'hc500810c, 32'hc3707df6, 32'h436d2da2},
  {32'h44d96300, 32'h43870b34, 32'hc1fa8771},
  {32'hc4b0fd8e, 32'h4083d52d, 32'hc1af2a0c},
  {32'h45145bbf, 32'hc34ac915, 32'hc300ca72},
  {32'hc51992e9, 32'h438fe803, 32'hc34436a8},
  {32'h42f17400, 32'h43e64662, 32'h42ab87bc},
  {32'hc361c510, 32'hc013b490, 32'h3e092c78},
  {32'h44cc222e, 32'h438cbc0b, 32'h42fe85f4},
  {32'hc40ad4a6, 32'hc329261d, 32'h42380193},
  {32'h437f58d1, 32'hc1780314, 32'h409bbe16},
  {32'hc48f352f, 32'h438461c5, 32'h4210f3d4},
  {32'h44ea981f, 32'hc245b746, 32'h4356b3bf},
  {32'hc4c5135e, 32'hc392472c, 32'h435cd1d8},
  {32'h44caaa24, 32'h4134cbab, 32'h42b43fc5},
  {32'hc4f1ece4, 32'hc346116e, 32'hc3f1f61b},
  {32'h45091346, 32'hc37f0b4c, 32'hc3ba7878},
  {32'hc4bd6b3a, 32'h43af9574, 32'hc2bdfe5f},
  {32'h4438541f, 32'h438b18d3, 32'h425dc5fc},
  {32'hc269cab2, 32'hc386615c, 32'hc1b05b4b},
  {32'hc30b289c, 32'hc3ef0220, 32'hc1d90d4e},
  {32'hc48a2773, 32'hc2c81118, 32'h43ad0f39},
  {32'h451196f0, 32'hc300de20, 32'h43d1c864},
  {32'hc405a031, 32'h438f36b1, 32'h433c498c},
  {32'h44ef19e5, 32'h438bee03, 32'h43f2c9b6},
  {32'hc490ed99, 32'hc3695456, 32'hc2a80bb9},
  {32'h4490eb81, 32'hc1b5f16e, 32'hc37e1a60},
  {32'hc4014ff2, 32'h43a92ccc, 32'hc3a8db4f},
  {32'h44d91173, 32'hc3b7a0a6, 32'h401a06f8},
  {32'hc46e397e, 32'h438365f5, 32'hc35df1e4},
  {32'h44007a64, 32'hc2aeacdd, 32'hc2fbf5e5},
  {32'hc512be0f, 32'hc28f4e10, 32'h43886c52},
  {32'h45129b93, 32'h43e92e93, 32'h41cd2bb8},
  {32'hc508d7f8, 32'hc319aa28, 32'h429e1d44},
  {32'hc29c203c, 32'h439e2e9c, 32'h42ee530e},
  {32'hc4d3eb60, 32'h43b24db6, 32'hc39b8beb},
  {32'h44c7b6cc, 32'hc281cba9, 32'hc340f032},
  {32'hc512e7af, 32'h41a88709, 32'hc2ac0254},
  {32'h449b26bc, 32'h4308485d, 32'h44364d09},
  {32'hc50fe6f3, 32'h42576f44, 32'h42fd1954},
  {32'h448ee917, 32'hc3be9ca2, 32'h4375164f},
  {32'hc485030d, 32'hc2648ff2, 32'h41d52072},
  {32'h4511be4b, 32'h422fc12e, 32'h42a66961},
  {32'hc3d67338, 32'hc39a12dd, 32'h435b461c},
  {32'h44bc0631, 32'h435ccda2, 32'hc38ff0f1},
  {32'hc4866274, 32'hc18308df, 32'h4222485b},
  {32'h45052f53, 32'h4300ac98, 32'h43b744dd},
  {32'hc4927d3a, 32'h4375b1ce, 32'h4382d2f7},
  {32'h43731c68, 32'hc321c474, 32'h413c6a22},
  {32'hc50ee5da, 32'hc34cc6a3, 32'h4226d0f4},
  {32'h449abc9f, 32'h434def9f, 32'hc3273d0b},
  {32'h41267480, 32'hc31bde8a, 32'h439b2684},
  {32'h44e53f14, 32'hc2bb5471, 32'h430c8fc3},
  {32'h404bb000, 32'h42915d0d, 32'h43447fba},
  {32'h4485bbc4, 32'hc38e28e7, 32'hc33d9bc3},
  {32'hc5005af5, 32'hc3469124, 32'h42b3e5ab},
  {32'h4509a22f, 32'h4429723f, 32'h439ff8ff},
  {32'hc511c7b6, 32'hc34eec06, 32'hc325b7da},
  {32'h450a7c13, 32'h4103d5eb, 32'hc3796b53},
  {32'hc49ed99e, 32'h424f9742, 32'h43106af3},
  {32'h44f72636, 32'hc3b695ea, 32'h43e043be},
  {32'hc4576094, 32'hc38e6b6f, 32'h42dc0a53},
  {32'h44975946, 32'h42ba2f67, 32'hc3e8b5c4},
  {32'hc4e5a14b, 32'hc3bade86, 32'hc326d5e0},
  {32'h43204100, 32'h42fc37f2, 32'hc25354fd},
  {32'hc4b5b3b2, 32'hc2262e69, 32'h435115ab},
  {32'h43081c0c, 32'h405d4d92, 32'h43afe179},
  {32'hc4a8017c, 32'hc3616e7c, 32'hc3525c04},
  {32'h4512f522, 32'h42129e42, 32'hc3415e68},
  {32'hc45352ef, 32'h4148633c, 32'hc281f4f5},
  {32'h4514f78c, 32'h424fc5b7, 32'hc3a1743a},
  {32'hc38f9398, 32'h4350ffd3, 32'hc1eb5c91},
  {32'h451dc5a1, 32'hc258d3d9, 32'h42cbe923},
  {32'hc4c1ae63, 32'hc2a44e44, 32'h4382ea13},
  {32'h443ae138, 32'h430fbb1c, 32'hc2e6669f},
  {32'hc51c8016, 32'h4300f9d2, 32'h4329dab8},
  {32'h450a2008, 32'hc278bf94, 32'h433dc4cc},
  {32'hc4698f8f, 32'hc316ca1a, 32'h435a3578},
  {32'h42ec5ef4, 32'hc2a82b9a, 32'h438f8252},
  {32'hc40c9bd0, 32'hc2f0fbab, 32'h43793a99},
  {32'h4472c37c, 32'hc3edafaf, 32'hc34adfe4},
  {32'hc4c530ed, 32'h4240f63a, 32'hc24adc5a},
  {32'h44125fcd, 32'hc27606fa, 32'hc2da0e03},
  {32'hc3059be0, 32'hc3362b98, 32'h437ae4df},
  {32'h44b26c3a, 32'h42f3309a, 32'h438bbd94},
  {32'hc49d5ea0, 32'h41bcfc2f, 32'h43937f8e},
  {32'h44a347cd, 32'hc2840099, 32'h42b77313},
  {32'h40adccc8, 32'h43e8cbdc, 32'hc3871185},
  {32'h44f4b820, 32'hc0d3cdfc, 32'h439e4fa1},
  {32'hc4af7fd3, 32'h421cd839, 32'h435c0ca2},
  {32'h450b6e98, 32'hc32122db, 32'hc1c65dfb},
  {32'hc48f436c, 32'h43cbf0b1, 32'hc38d0671},
  {32'h44776ae0, 32'h43ae5f6d, 32'hc2bde72a},
  {32'hc384026c, 32'hc1290d19, 32'hc318fe00},
  {32'h4464ebbc, 32'h42afa747, 32'h441a5aaa},
  {32'hc4f88b0b, 32'h43a5fcbb, 32'h43b4570c},
  {32'h4387d850, 32'h43320b8f, 32'h4390094d},
  {32'hc46d878f, 32'hc2b550d7, 32'hc3329b79},
  {32'h44ff6683, 32'hc1db875c, 32'h43485da2},
  {32'hc494250a, 32'hc3351ddc, 32'hc24f14f0},
  {32'h44749c24, 32'hc176a725, 32'hc3aed78c},
  {32'hc4fe8a85, 32'h4313ca4c, 32'hc3c2b2f4},
  {32'h450f0031, 32'hc368294b, 32'h43da443e},
  {32'hc48caceb, 32'hc1e2d84c, 32'hc323a9eb},
  {32'h440af776, 32'h43b43fba, 32'h4301107d},
  {32'hc4103bd2, 32'h435e2bcd, 32'h435c2890},
  {32'h4536ea27, 32'h4135d58f, 32'h432df7c8},
  {32'hc2041fc0, 32'h43c1d710, 32'h43b48383},
  {32'h45163569, 32'hc28cf717, 32'hc3b1f347},
  {32'hc3e6b212, 32'h43cc784f, 32'h434b7634},
  {32'h43ef0afb, 32'hc310675e, 32'hc1fb3672},
  {32'hc4ca9e9a, 32'hc32bed00, 32'h426deceb},
  {32'h44e05dbd, 32'h4327fd87, 32'hc2238472},
  {32'hc4c3da97, 32'hc3c37240, 32'h4289ac3e},
  {32'h44955764, 32'hc1a46073, 32'hc35cf989},
  {32'hc40c1408, 32'h4327652a, 32'hc3641864},
  {32'h4515e4bf, 32'h4329d15e, 32'h42725fe4},
  {32'hc4eafb07, 32'hc1e5b17e, 32'hc2b5ffab},
  {32'h447ad552, 32'h437e33f4, 32'hc2aad63b},
  {32'hc4a7ff3c, 32'h42c5b699, 32'hc2dd89e4},
  {32'h452566ce, 32'hc296537c, 32'hc28d9068},
  {32'hc51390a4, 32'hbea1e3d4, 32'hc2072492},
  {32'h41a68f10, 32'hc357353f, 32'h4370ac01},
  {32'hc46e6f3c, 32'hc23c63c2, 32'hc38b4219},
  {32'h443d2582, 32'hc2e7497c, 32'hc2c8c8d7},
  {32'hc439f146, 32'h43319d4f, 32'h42a413b0},
  {32'h43fb59e8, 32'hc30e6520, 32'h424ba1d9},
  {32'h4181bec0, 32'h436a373e, 32'hc434c522},
  {32'h4499455b, 32'h44044efd, 32'hc311c71d},
  {32'hc2b115c4, 32'hc00ced10, 32'h420d6cdd},
  {32'h450b9e29, 32'hc33b911d, 32'hc33bdac8},
  {32'hc47a4b90, 32'h438178d9, 32'hc1b85662},
  {32'h44ce55b1, 32'h4263ee81, 32'h43c44964},
  {32'hc388a630, 32'hc37e0104, 32'h42d519f2},
  {32'h448487b7, 32'h436f9c4c, 32'h43c7f03d},
  {32'hc4758a0a, 32'h43523264, 32'hc2676104},
  {32'h44ef22ff, 32'hc05e3028, 32'hc3c5f7e9},
  {32'hc3243617, 32'h430eb488, 32'hc112ac71},
  {32'h449f1c0a, 32'h439f719a, 32'h43c6c4de},
  {32'h415ac7a0, 32'hc2fb3c87, 32'h42ef2155},
  {32'h44360923, 32'h435ee1d7, 32'h42fbf478},
  {32'hc2a11140, 32'hc341fcc9, 32'h438a69e2},
  {32'h44b59352, 32'hc28bc060, 32'h43d1849e},
  {32'hc4e57867, 32'h438325f8, 32'hc23d702f},
  {32'h44fc212e, 32'h42db257c, 32'hc31b0a8f},
  {32'hc4c5f2a1, 32'h43afde82, 32'hc2f94ad0},
  {32'h449c59e6, 32'h40b546ee, 32'hc29ebe26},
  {32'hc48d631c, 32'h434041a8, 32'hc16d4655},
  {32'h445d24f2, 32'h4319a77a, 32'hc255cba6},
  {32'hc4a1df88, 32'hc2c650a8, 32'hc3ae46fb},
  {32'h44facb36, 32'h4108bd90, 32'hc301ed65},
  {32'hc4f4a8ec, 32'hc19c2af8, 32'hc25e86a7},
  {32'h44fb2891, 32'hc3427266, 32'hc33e6d23},
  {32'hc45908a7, 32'hbf0f89e0, 32'h42e98eca},
  {32'h446a1033, 32'hc3b06e18, 32'h42a4f466},
  {32'hc52c8869, 32'h43564278, 32'h4354fc2c},
  {32'h440ca025, 32'h3f20d4cf, 32'h431b11a1},
  {32'hc4d9a209, 32'hc3142645, 32'h4258c236},
  {32'hc3fa8658, 32'hc39414a2, 32'hc317d43e},
  {32'h44dbbba3, 32'hc27bf308, 32'hc2d815bd},
  {32'hc50d24f7, 32'h4188dc0c, 32'hc1f68472},
  {32'h44d466df, 32'hbf8cacb7, 32'h432e9273},
  {32'hc4da56ba, 32'hc31fd360, 32'hc20405a8},
  {32'h445db41f, 32'hc341ce28, 32'h43bcf888},
  {32'hc4de669f, 32'hc3dbb66d, 32'hc39608c6},
  {32'h44f407c8, 32'hc288b112, 32'h438c167b},
  {32'hc4a85580, 32'hc33447c8, 32'h417b29fc},
  {32'h42e5aa20, 32'h425a365c, 32'hc30c4588},
  {32'hc4d0276b, 32'h43956ab7, 32'hc32bc1f7},
  {32'h44e4d10e, 32'hc254c633, 32'hc35a13c3},
  {32'hc48d120e, 32'hc1bbe176, 32'hc33b30ef},
  {32'h450efda8, 32'h4272e7ca, 32'hc331bfb8},
  {32'hc4fb2b40, 32'h42f95079, 32'h430f0f52},
  {32'h444647c8, 32'hc06895a0, 32'h4248c8bd},
  {32'hc4a4cb44, 32'hc289b95c, 32'h42f61594},
  {32'h44d30ab2, 32'h43189ff7, 32'h41b76c88},
  {32'hc4bcc9ee, 32'hc33ccff3, 32'hc3c24fda},
  {32'h44006ea1, 32'h40353150, 32'hc2c8949d},
  {32'hc505ef26, 32'h43062933, 32'h4246a415},
  {32'h44c4bf54, 32'h41cfd942, 32'h42661fbc},
  {32'hc5042f5a, 32'hc31481f0, 32'hc28b0f21},
  {32'h44549d46, 32'h43879fdc, 32'hc2fdb370},
  {32'hc4b30b86, 32'hc332c1a3, 32'hc35e24c5},
  {32'h44dfdfb4, 32'hc15173f1, 32'hc2e92997},
  {32'hc44ca68d, 32'hc2058a18, 32'h4396dbd9},
  {32'h4446db22, 32'hc359fde0, 32'hc32cbd12},
  {32'hc4bde4ad, 32'hc301a704, 32'hc3986a2d},
  {32'h44587040, 32'h4305ec74, 32'hc24cef99},
  {32'h41fbc8a8, 32'h43e3697e, 32'hc2c94820},
  {32'hc390ecd8, 32'hc2998ded, 32'h44057ab1},
  {32'hc50d4e22, 32'hc2e9331f, 32'h41d0a6e7},
  {32'h44b7897b, 32'hc1aa1599, 32'hc2017cd4},
  {32'hc5209cd5, 32'hc334fbf5, 32'h436d4e06},
  {32'h43f70fda, 32'hc314d605, 32'hc3884e9c},
  {32'hc4ab7a47, 32'hc36986bd, 32'hc37c25d5},
  {32'h44a2464c, 32'h440b97b2, 32'hc2cfae82},
  {32'hc292c14a, 32'hc2af9d76, 32'hc3878709},
  {32'h418d6000, 32'h42aae41c, 32'hc3a927bd},
  {32'hc3df05c8, 32'hc25fe0fe, 32'hc33f6e78},
  {32'h445799fe, 32'hc2c170b8, 32'hc3c4aead},
  {32'hc463776d, 32'h438f6358, 32'h4389bbc3},
  {32'h4481d01c, 32'h433fa62d, 32'h43305272},
  {32'hc509d4d9, 32'h4386441c, 32'h432aa9f3},
  {32'h44b43fc4, 32'hc3955aec, 32'hc34e34d8},
  {32'hc3a37c74, 32'hc2ff280f, 32'h43c4c325},
  {32'h44f50980, 32'hc2b92882, 32'h438f757e},
  {32'hc4ba20cb, 32'hc2f1de48, 32'hc33ca5fd},
  {32'h4491477b, 32'hc2a1123c, 32'hc13f0cde},
  {32'hc4b7223b, 32'hc381778a, 32'h42159893},
  {32'h446659ec, 32'h43c50574, 32'h43709cae},
  {32'hc506a0bf, 32'hc313d392, 32'hc3303ecd},
  {32'h448e6047, 32'h42ad3899, 32'hc1f3b251},
  {32'h42ef7cae, 32'hc35d9638, 32'hc19835bd},
  {32'h44af9d2d, 32'hc3797fe5, 32'hc31bb7a9},
  {32'hc46f66ac, 32'h43c4c546, 32'hc242eedf},
  {32'h447b0dcc, 32'h42a4874a, 32'hc3a9d92a},
  {32'hc4801e79, 32'hc324c186, 32'h4281199f},
  {32'h4226a236, 32'hc3b24e81, 32'h44225c80},
  {32'hc50e3ecc, 32'hc39fa40e, 32'h42f00750},
  {32'h44ad6de4, 32'hc2ad944d, 32'h42046d91},
  {32'hc50c0a8d, 32'hc2bb8f72, 32'hc3d63f41},
  {32'h449c1ffd, 32'h43bd1a96, 32'h431d10c6},
  {32'hc4b40785, 32'h435e2df5, 32'h43d7eedc},
  {32'h4388b220, 32'h431aeb92, 32'h43db43e0},
  {32'hc4ed34e5, 32'hc29c06ca, 32'hc2a16af8},
  {32'h4482b5bb, 32'hc3c7a639, 32'hc3704bcc},
  {32'hc38ce182, 32'h43163584, 32'hc2e6d09f},
  {32'h4471c440, 32'hc3bf512c, 32'hc3c88410},
  {32'hc50273f2, 32'h437f80f1, 32'h42d66eb6},
  {32'h44f92cea, 32'hc319affa, 32'h43652722},
  {32'hc5056752, 32'hc1a4bd42, 32'hc35569f4},
  {32'h44ad881c, 32'h43110556, 32'h43c494ea},
  {32'h4397355c, 32'h41d22c9d, 32'h437b3011},
  {32'h43b41ec0, 32'h42e0a4ca, 32'h43c0331d},
  {32'hc426db80, 32'h42049321, 32'h42c27ace},
  {32'h45019750, 32'h42ab56f7, 32'hc37a0887},
  {32'hc4c7f5f2, 32'h4306287b, 32'h41c00d60},
  {32'h448c08c2, 32'hc2fafb39, 32'h43e63c83},
  {32'hc519bc96, 32'hc33f26ab, 32'hc2d57232},
  {32'h442a322a, 32'hc3a28029, 32'h4339ea40},
  {32'hc436fa87, 32'h42a114b4, 32'hc30aec1a},
  {32'h44cd2367, 32'hc33d515f, 32'h44226115},
  {32'hc4c284b0, 32'hc0cb1f28, 32'h42450018},
  {32'h44c951c3, 32'hc36ac351, 32'hc2b5f013},
  {32'h41885580, 32'h42f6b438, 32'hc383cad7},
  {32'h4302cbbb, 32'h430d81ec, 32'h437c2dde},
  {32'hc4e8598b, 32'h4309549d, 32'hc30df896},
  {32'h44fb3aee, 32'hc3322bb2, 32'h42efcf73},
  {32'hc3e0d220, 32'hc2e489d4, 32'h410e6094},
  {32'h44a5764b, 32'h42865a17, 32'h42859c16},
  {32'hc3b764c2, 32'hc2eacb2e, 32'h3f2fc36c},
  {32'h4491f266, 32'h438dce49, 32'h431536be},
  {32'hc50e3b6c, 32'hc2f0302d, 32'hc34fe09a},
  {32'h45068ef2, 32'h4336a7db, 32'hc397a6f0},
  {32'hc2d55020, 32'h412807ab, 32'h43d37056},
  {32'h44af2049, 32'h42be5d37, 32'h42ae124d},
  {32'hc4d7a52c, 32'hc39bb65a, 32'h4397d220},
  {32'h440bdc66, 32'hc391f26a, 32'h4402f2d4},
  {32'hc1455754, 32'h41acc738, 32'hc372c194},
  {32'h44e43000, 32'hc3101013, 32'h41963943},
  {32'hc4b7279a, 32'hc2b0b18a, 32'h42c6e4d6},
  {32'h44005515, 32'hc153d0eb, 32'h43f1a3dc},
  {32'hc4400645, 32'h43915b1d, 32'h438aabf8},
  {32'h44d3b1c1, 32'hc1e44191, 32'h41d839d0},
  {32'hc48e06d1, 32'h431bed2c, 32'h43157e10},
  {32'h4508c81b, 32'hc1c4d79e, 32'h404da758},
  {32'hc4234164, 32'h41df66a2, 32'hc1696a12},
  {32'h44ebfc4d, 32'h4341286b, 32'h433d7e5a},
  {32'hc4d78f1c, 32'hc37465da, 32'hc3c32906},
  {32'h43c6da58, 32'h4383c1cc, 32'hc2d80adf},
  {32'hc505114a, 32'h4321f2ed, 32'hc31675b8},
  {32'h445e2e2c, 32'h427dd39d, 32'hc324e73e},
  {32'hc413ce6c, 32'hc330629a, 32'hc31e5d31},
  {32'hc4057d4a, 32'h4285c18e, 32'hc282c490},
  {32'hc4055e92, 32'hc2c03f7b, 32'h43469a22},
  {32'h44e4243f, 32'hc2e7d147, 32'h4372dad9},
  {32'hc4e8d49a, 32'h4373a068, 32'h42abd099},
  {32'h4527a30e, 32'h434e626a, 32'hc40310ee},
  {32'hc41bc6cc, 32'hc2e50ed8, 32'h42c31d8f},
  {32'h43e73960, 32'h429eba88, 32'h43e050c4},
  {32'hc4da9aae, 32'hc3a341fe, 32'hc2c0990b},
  {32'h4494c334, 32'hc28d2896, 32'hc2a1ba70},
  {32'hc4b155ef, 32'hc3258306, 32'h436a35b8},
  {32'h44958bc0, 32'h435cc481, 32'h4302ff93},
  {32'hc3973cd2, 32'hc292839f, 32'h432b7689},
  {32'h4493f753, 32'hc39d8ffd, 32'hc26bb789},
  {32'hc42b1e06, 32'h436740b3, 32'hc366cf53},
  {32'h44e5d7d4, 32'hc2a4b86d, 32'hc341ae88},
  {32'hc4086f19, 32'hc3a49414, 32'h432376f9},
  {32'h44fc75e1, 32'hc3ece23e, 32'h4438d24b},
  {32'hc3136d50, 32'hc388678e, 32'h420b60ed},
  {32'h4457eb5f, 32'hc2850572, 32'hc200bb30},
  {32'h42f863ca, 32'hc2f3a8e7, 32'hc33c14cb},
  {32'h44f78e04, 32'hc354b846, 32'hc32ba56f},
  {32'hc48c7b5f, 32'hc1b9757c, 32'hc30af91f},
  {32'h451003dc, 32'hc2887158, 32'hc25bc013},
  {32'hc387dfa6, 32'h41b54bb6, 32'hc3942ce1},
  {32'h450a1fa2, 32'h439a2e11, 32'h438c3a3a},
  {32'hc4b9f743, 32'h4389e3bc, 32'h435bd2c2},
  {32'h43a536f6, 32'hc37a004b, 32'hc2b9cd66},
  {32'hc308f05c, 32'h437638f5, 32'h435f7e77},
  {32'h440e7c56, 32'hc38069cd, 32'hc3ca69da},
  {32'hc488e504, 32'h429a3d37, 32'h432e5d41},
  {32'h44fed74d, 32'h425e9586, 32'hc3ae07b1},
  {32'hc4690c36, 32'h4326a61c, 32'h429f0e8b},
  {32'h45133d0c, 32'hc2c89422, 32'h427a3565},
  {32'hc43764a1, 32'hc4142557, 32'h43b7c93d},
  {32'h44499358, 32'h40e16b46, 32'hc3fc6543},
  {32'hc3753188, 32'h43544eea, 32'hc2f7e0ef},
  {32'h41eb4000, 32'h421fbe3b, 32'h4247a454},
  {32'hc4e37c80, 32'h423c7fee, 32'h428a96db},
  {32'h42992a20, 32'hc1c42784, 32'h43c78aea},
  {32'hc4ad77a3, 32'hc3aa8414, 32'hc3145c34},
  {32'h44d67c2e, 32'hc3ac9b27, 32'hc36b507b},
  {32'hc34fdc88, 32'hc32057c9, 32'h430fed28},
  {32'h4407d8b0, 32'hc33abb12, 32'h438f504f},
  {32'hc489d598, 32'hc321b92f, 32'hc28a4d5a},
  {32'hc1625380, 32'h43682821, 32'h41a122b6},
  {32'hc50f555a, 32'h404e6c61, 32'h42c6e0ef},
  {32'h4403e440, 32'h4354ca9a, 32'h43959eb0},
  {32'hc3eea79a, 32'hc1e0b172, 32'h4316c092},
  {32'h4464e264, 32'hc29a012b, 32'h42931e2e},
  {32'hc3d13046, 32'hc31f80df, 32'h433c0832},
  {32'h43d31430, 32'hc32536b8, 32'h416723b4},
  {32'hc492dd48, 32'hc373b9c6, 32'hc47a70d7},
  {32'h44cea5bc, 32'h432fd9c3, 32'h43d44d3f},
  {32'hc16ba500, 32'hc3118432, 32'hc3120458},
  {32'h44b65e12, 32'hc3ea4dea, 32'h43e708b0},
  {32'hc4101894, 32'h43a1ffbc, 32'hc1d041ca},
  {32'h43fa98f0, 32'h4024ca40, 32'hc28fd036},
  {32'hc4c9363e, 32'hc37e68a7, 32'h4375596b},
  {32'h450195be, 32'hc2cc113c, 32'hc2eec770},
  {32'hc4a9c89a, 32'h43204f26, 32'h434f89cd},
  {32'h45069864, 32'hc3c646d6, 32'h439c5d96},
  {32'hc46b4b30, 32'h430586c7, 32'hc27adf54},
  {32'h44f6d7e0, 32'hc32763da, 32'hc328e2c4},
  {32'hc4af243b, 32'hc369d5eb, 32'hc360842c},
  {32'h451ae05a, 32'h42ce8197, 32'hc32f7080},
  {32'hc50861a0, 32'h43934f9f, 32'hc36bcdc5},
  {32'h444c5380, 32'h43fd0867, 32'h434fa9b6},
  {32'hc463c95e, 32'h41609ff1, 32'hc3ded692},
  {32'h442e3dac, 32'h43db5840, 32'hc308bcb1},
  {32'hc40ec520, 32'hc2c4c67c, 32'h437179eb},
  {32'h43a99fc0, 32'h4301199a, 32'h429a1ed7},
  {32'hc4d33b9b, 32'h43287a88, 32'h42fc30c9},
  {32'h441674d0, 32'hc1987f38, 32'h42fc8e57},
  {32'hc513bf4f, 32'h41d3dc03, 32'h432b5e08},
  {32'h4398607e, 32'h43c67108, 32'h434034fc},
  {32'hc42eda9d, 32'h41b07c10, 32'hc2d387ed},
  {32'h42cb8260, 32'hc269a52b, 32'hc2fd857a},
  {32'hc38b1c50, 32'hc381418b, 32'hc31c7af2},
  {32'h4492a3b2, 32'hc3db6891, 32'h427647e0},
  {32'hc4a6141e, 32'h4392e4f2, 32'hc2d2a59e},
  {32'h451191e2, 32'hc2fb7d45, 32'h43558451},
  {32'hc50ee4f0, 32'hc2f9a451, 32'h436b11dc},
  {32'h44c5137e, 32'hbfff8194, 32'hc2547a13},
  {32'h427c66a4, 32'hc3516b67, 32'h42ff6c84},
  {32'h42f4df1e, 32'hc3ba7e80, 32'h4390389b},
  {32'hc4a88aad, 32'hc34377e8, 32'h43698d70},
  {32'h44482e5a, 32'h42de39ac, 32'h42628bbe},
  {32'hc4a5a3b5, 32'hc3729c23, 32'h429a7de4},
  {32'h450cda4d, 32'h433497b3, 32'h42b8fe2f},
  {32'hc44e9600, 32'h431a6a46, 32'hc2d00cdc},
  {32'h42e54b70, 32'hc3249aa1, 32'h430613e2},
  {32'hc4955348, 32'hc26fc012, 32'h43bbde2d},
  {32'h44e6f700, 32'h4370cb4c, 32'hc0b4a85d},
  {32'hc401670c, 32'h426ad344, 32'hc313b8e8},
  {32'h450e391b, 32'hc2340321, 32'hc2be424a},
  {32'hc4a569ae, 32'h43251569, 32'h43233cdc},
  {32'h44add57d, 32'h42d8e24a, 32'hc2658704},
  {32'hc4caa31b, 32'h43ce0a4c, 32'h434169dd},
  {32'h43fe9244, 32'hc3fe8c03, 32'hc241c58b},
  {32'hc4efd05e, 32'h42efcf75, 32'h42f8ed90},
  {32'h450fea9b, 32'hc3184c59, 32'h430cb7cf},
  {32'hc4f09ee3, 32'h42d2142b, 32'hc343104d},
  {32'h450097a8, 32'hc32b2eba, 32'hc2f95e74},
  {32'hc4b81712, 32'h43a3dfa9, 32'hc28b93d6},
  {32'h44f0da6b, 32'hc395572f, 32'hc26db41a},
  {32'hc3fe04c0, 32'hc3a43278, 32'h411a1d06},
  {32'h44949b61, 32'hc413fe3c, 32'hc34c90ea},
  {32'hc458ede2, 32'h43d284b2, 32'hc372c192},
  {32'h44aec294, 32'h42899db1, 32'hc2cf05de},
  {32'hc4bdbb58, 32'h4213ca29, 32'h4304704d},
  {32'h4508fdcd, 32'h43921246, 32'h4332ccf5},
  {32'hc4f19bc6, 32'h43a64724, 32'hc387479d},
  {32'h4387a470, 32'hc2ff1bb8, 32'hc37a1915},
  {32'hc4f75782, 32'h4212610b, 32'h4325d265},
  {32'h448c5268, 32'h43700f6e, 32'hc1de1062},
  {32'hc4444d73, 32'h429ee722, 32'hc361f005},
  {32'h441a0428, 32'h41e814d8, 32'hc290fa9d},
  {32'hc505ac9e, 32'h4320c9f4, 32'hc25b329a},
  {32'h44f029f6, 32'hc3811219, 32'h42221314},
  {32'hc487b4a8, 32'hc3803921, 32'hc1b27ff4},
  {32'h4469aebe, 32'hc3e3679d, 32'hc23aced0},
  {32'hc4de7105, 32'h43453622, 32'h41765bf1},
  {32'h434c28d0, 32'hc32619c8, 32'hc353b05c},
  {32'hc50ed408, 32'hc2678da3, 32'hc257abe7},
  {32'h44dca18a, 32'hc31f7181, 32'h4382c5ad},
  {32'hc4ed20e5, 32'h438b1297, 32'hc391f34e},
  {32'h44fe3e0b, 32'h428eb690, 32'h438c7eec},
  {32'hc3a05808, 32'h42d7a9ab, 32'hc2c65e38},
  {32'h44dbac10, 32'hc2582453, 32'h43243dc9},
  {32'h42490640, 32'h42dcb52f, 32'hc2c95ee0},
  {32'h449f2ba4, 32'h43b10dd4, 32'h43435081},
  {32'hc5036288, 32'hc2db3c56, 32'h4386771a},
  {32'h44a59708, 32'hc23d5b98, 32'h43a49ce2},
  {32'hc44150f6, 32'hc3b91ece, 32'hc38df05d},
  {32'h4494b7ec, 32'hc33738aa, 32'h41e8e24f},
  {32'hc3d88324, 32'h435544d8, 32'h43b48f3b},
  {32'h44e8e40b, 32'hc27b5682, 32'hc3a73331},
  {32'hc42145f0, 32'hc40615ef, 32'h43759a24},
  {32'h442226d3, 32'h413488f8, 32'hc3bde558},
  {32'hc4849b2d, 32'hc3fbab77, 32'hc2ee91ce},
  {32'h4468fdc4, 32'h439b7864, 32'h429967a4},
  {32'h41c01984, 32'h43debb3e, 32'h427f0112},
  {32'h439a1518, 32'h41dc4e4d, 32'hc3885780},
  {32'hc4e9fd1a, 32'h43393a76, 32'hc3aa81b7},
  {32'h448e043e, 32'h43484156, 32'hc23b2dd4},
  {32'hc48119f3, 32'hc2a0d740, 32'hc3797021},
  {32'h44b2e232, 32'hc3a18114, 32'hc1e118b8},
  {32'hc420c882, 32'hc11ed903, 32'h43a713d2},
  {32'h43c2cba6, 32'h438ea994, 32'h43a5533d},
  {32'hc4d0f4ed, 32'hc320a1c2, 32'hc3376142},
  {32'h4441fcbc, 32'h435c6e3c, 32'h42f62b07},
  {32'hc241ed70, 32'hc1859fc3, 32'h41e24296},
  {32'h43bd253c, 32'hc18d947c, 32'h4232c2ae},
  {32'hc4a0c27f, 32'h41062893, 32'h42dad6a4},
  {32'h44a46231, 32'hc30d5112, 32'h42cd604d},
  {32'hc4f567d0, 32'h435408b4, 32'h433acc80},
  {32'h4504e135, 32'hc364ba4e, 32'hc31712d2},
  {32'hc26038c0, 32'h42ea642f, 32'hc347ba96},
  {32'h45044b8e, 32'h42730540, 32'hc259da54},
  {32'hc4309cb4, 32'h42e4e058, 32'hc2bd3bb1},
  {32'h44d5d999, 32'hc3516a45, 32'hc3474a81},
  {32'hc408e71d, 32'hc32389af, 32'h439cd8cf},
  {32'h42061bb0, 32'h42ee0e8d, 32'h4226da9c},
  {32'hc3ef8351, 32'hc3938e28, 32'hc1bf8901},
  {32'h44e67d35, 32'hc24cce3a, 32'h431de900},
  {32'hc490a676, 32'hc2e42be3, 32'h431c5b6e},
  {32'h43927af0, 32'hc32d4d82, 32'h4244910d},
  {32'hc348db14, 32'h43a18315, 32'h439ea5dc},
  {32'h44b8a506, 32'h410f4bc6, 32'h439836f3},
  {32'hc499573e, 32'h42e40ee9, 32'hc170f6ac},
  {32'h450d4411, 32'hc355236a, 32'h419e0515},
  {32'hc510dc2a, 32'h43a82f0a, 32'h42c057e7},
  {32'h44f8692c, 32'h43430efe, 32'h43381722},
  {32'hc2d35820, 32'h4218cd3a, 32'h4315d3fb},
  {32'h4475472d, 32'hc19c08f8, 32'h432c4568},
  {32'hc4f25eec, 32'hc32ac797, 32'h4327af4f},
  {32'h45142491, 32'h4375f011, 32'h43806bdc},
  {32'hc32fc440, 32'h43635d03, 32'h432fdbc8},
  {32'h45073c82, 32'h4354ddde, 32'hc32072c6},
  {32'hc4e0605a, 32'hc28298f2, 32'hc33f1507},
  {32'h44944aaa, 32'hc3af9fa8, 32'hc416b357},
  {32'hc48fc894, 32'h4319d176, 32'h43a690c9},
  {32'h4513b9b7, 32'hc2d8b9c0, 32'h43673094},
  {32'hc3f0cd14, 32'hc1050d93, 32'h4376dc40},
  {32'h442f8156, 32'hc3889902, 32'hc26d6ebc},
  {32'hc3094148, 32'h433c6ee4, 32'hc3be1589},
  {32'h44aed226, 32'hc347c95e, 32'hc39f3bba},
  {32'hc4a15f8c, 32'h442e3f01, 32'hc30d04af},
  {32'h44141604, 32'h41e98855, 32'hc2f5e97c},
  {32'hc4818383, 32'hc42b8dc7, 32'h435cf162},
  {32'h44dfc07d, 32'hc1b6f7c8, 32'h427fbd85},
  {32'hc4a905bd, 32'h42981133, 32'hc2e2568b},
  {32'h442d5268, 32'hc3e12697, 32'hc1fc2765},
  {32'hc498a70d, 32'hc36d76cf, 32'h4322ec9c},
  {32'h44ed70f2, 32'h4419bc1a, 32'hc2d6691b},
  {32'hc4326984, 32'hc383c65c, 32'hc2bb023b},
  {32'h44ee3d41, 32'h4127cd33, 32'h43188faf},
  {32'hc16fd000, 32'hc36bc048, 32'h420731c7},
  {32'h443bdf0d, 32'h43e070f5, 32'h42e6faa7},
  {32'hc2c8fd80, 32'h43db6bc1, 32'hc3061335},
  {32'h441dbedd, 32'hc362495f, 32'hc313bc64},
  {32'hc4fc4c9b, 32'h4346a76a, 32'hc30ebb9c},
  {32'h44806773, 32'h42ffe1a0, 32'hc21f56c2},
  {32'hc4961b57, 32'h43c1ff19, 32'hc30edf69},
  {32'h44ecfbf4, 32'h423dfa84, 32'h432ace98},
  {32'hc4618bfa, 32'hc40bd9df, 32'hc2eff293},
  {32'h4485b9dc, 32'hc3633d9a, 32'hc346d136},
  {32'hc4c04497, 32'h422849fd, 32'hc4357bd3},
  {32'h43e951f0, 32'hc385bb93, 32'h42dbc263},
  {32'hc2eff648, 32'h435ca026, 32'hc0bda425},
  {32'h44dece78, 32'hc1aca048, 32'h42b428ca},
  {32'hc0f67100, 32'h43b1e572, 32'h435f9423},
  {32'h4507dc18, 32'h43d61cca, 32'h423f207c},
  {32'hc4b94b0f, 32'h437b62d6, 32'h430abc0c},
  {32'h4513381b, 32'h433c7e3e, 32'hc3f09895},
  {32'hc4a5c131, 32'hc306681c, 32'hc2a213ef},
  {32'h4515a911, 32'h42d3c856, 32'h433c659d},
  {32'hc5049bc3, 32'h419dcb67, 32'hc30d1c4c},
  {32'h450404a7, 32'h42f277b3, 32'hc2f67952},
  {32'hc504003d, 32'hc2b052e0, 32'hc1cbdef0},
  {32'h44dad2d1, 32'h4264c622, 32'hc31759b2},
  {32'hc45ae9de, 32'h440d18c8, 32'hc3b278cb},
  {32'h44abaf4c, 32'h430914ca, 32'hc307c415},
  {32'hc4fb7c66, 32'hc238507c, 32'hc3577d5d},
  {32'h4444adb2, 32'h4316a2ea, 32'h42d16dbf},
  {32'hc1d4e600, 32'hc3f19586, 32'h41e05314},
  {32'h44e4dfe6, 32'hc32e8a40, 32'hc3168902},
  {32'hc44b96d5, 32'h4321878e, 32'h432d9587},
  {32'h44ead4ca, 32'hc07d0fb4, 32'hc0a814a8},
  {32'hc5257ffb, 32'hc2a9ef26, 32'hc2e557a3},
  {32'h45074940, 32'h437855da, 32'hc358799d},
  {32'hc4a87d56, 32'h43233c16, 32'h42da3fe1},
  {32'h44dac1da, 32'h432a4dd2, 32'hc11238c8},
  {32'hc4c6ff13, 32'h4302a9d4, 32'hc1afcc8f},
  {32'h450bedb9, 32'h43292446, 32'hc3a31383},
  {32'hc30cd401, 32'hc3a2446d, 32'h43bd7e1e},
  {32'h450da5e0, 32'hc3365bdf, 32'hc39e700a},
  {32'hc5101cf2, 32'h42d81ce1, 32'hc21389f7},
  {32'h4434df3e, 32'hc400137b, 32'h43498190},
  {32'hc50b167d, 32'hc3944252, 32'hc3afbb80},
  {32'h448e46ac, 32'hc376bea7, 32'h43bbe5a7},
  {32'hc48893e9, 32'hc380b80e, 32'hc307e0ec},
  {32'h43a9f343, 32'hc383fadc, 32'h4372309b},
  {32'hc47d148c, 32'hc21ed5b1, 32'hc2594440},
  {32'h44e331d4, 32'hc2dcb08d, 32'h421c5e94},
  {32'hc51344ba, 32'h42c55e6a, 32'hc1b98539},
  {32'h449c77fa, 32'h3e0d4c80, 32'h43805cea},
  {32'hc4e1c02f, 32'h43ca4ea8, 32'hc080c1cd},
  {32'h43f89063, 32'hc26e91c3, 32'h4391165f},
  {32'hc4fad0f4, 32'hc3a2a7c0, 32'h4309f7f2},
  {32'h4457014f, 32'hc2f2a53c, 32'hc32f7200},
  {32'hc4bab47e, 32'hc350cdb6, 32'hc36f4376},
  {32'h44f11269, 32'h430fb852, 32'hc37d10d3},
  {32'hc4c7b91e, 32'h43c49549, 32'h42d0c668},
  {32'h44fba896, 32'h41dae6f8, 32'hc0234370},
  {32'h43215bda, 32'h4313df49, 32'h437cd656},
  {32'h44e430d3, 32'hc14cdd07, 32'hc2471484},
  {32'h435b1a78, 32'h429b1544, 32'hc30ae82b},
  {32'h43e51902, 32'hc2b9140d, 32'h428f654c},
  {32'hc4180df8, 32'h439cc55b, 32'hc4199b15},
  {32'h44870d24, 32'hc32000b8, 32'h40af5d7a},
  {32'hc449417c, 32'hc1e28c88, 32'h41747243},
  {32'h451f39f3, 32'hc25c2ac7, 32'hc345c419},
  {32'hc36c01e8, 32'hc21ace3d, 32'hc3173ddd},
  {32'h4407d2ec, 32'h4230475f, 32'h428e0b1b},
  {32'hc4410862, 32'h43507318, 32'hc312147d},
  {32'h4492eb0a, 32'hc32e816a, 32'h42d006ce},
  {32'hc41bbc16, 32'hc2f3faa0, 32'h43a4913b},
  {32'h44993c4e, 32'hc2ee77f7, 32'h42c73583},
  {32'hc4a524e3, 32'hc30ac0a6, 32'h43617e64},
  {32'h446e3704, 32'h42450303, 32'h436ca953},
  {32'hc43e4812, 32'hc33cbc17, 32'h41d4c081},
  {32'h4312a040, 32'hc41139f3, 32'hc3228b41},
  {32'hc51027dd, 32'h4409b2b2, 32'hc10ad210},
  {32'h44e0905b, 32'hc344cc64, 32'hc3133f2e},
  {32'hc4e4b398, 32'h42cfb9cb, 32'h43718232},
  {32'h43267390, 32'hc3c54134, 32'h42d24b9b},
  {32'hc4a2a7d7, 32'h43298b1f, 32'hc2ac5518},
  {32'h450b2d1a, 32'hc3aec50b, 32'hbf2e33a8},
  {32'hc3af669c, 32'hc302b251, 32'h42de7a05},
  {32'h44943d51, 32'hc3b63886, 32'h4210e488},
  {32'hc516a58f, 32'h4103ccf3, 32'hc36af77c},
  {32'h431a2ec2, 32'hc38aaa4b, 32'hc34b1f4b},
  {32'hc4cb9602, 32'h41a8ed08, 32'h43e77158},
  {32'h438c8300, 32'hc230d618, 32'hc3bd3ffa},
  {32'hc50745ca, 32'h437fd471, 32'h425785b9},
  {32'h44442e48, 32'hc3b4ad54, 32'hc395b00f},
  {32'hc3766eb0, 32'hc333de7f, 32'hc24e23f6},
  {32'h44e48d54, 32'hc3b33d24, 32'hc3138ed7},
  {32'hc4b4fdd4, 32'h43053be9, 32'h43283ea5},
  {32'h447ca385, 32'h42adc43c, 32'h43f1ae26},
  {32'hc4b2c863, 32'hc27729aa, 32'hc2dcf656},
  {32'h44b8d62a, 32'hc3ad007b, 32'hc304176f},
  {32'hc4e6cebe, 32'h43db2841, 32'h41a97906},
  {32'h427bbca0, 32'h43571101, 32'h432255e7},
  {32'hc4708e21, 32'h43b9c974, 32'h43fff0fb},
  {32'h4461b2ab, 32'h43b29c67, 32'h4322545f},
  {32'h41b58380, 32'hbf014594, 32'h429681ff},
  {32'h45154a95, 32'h43650c52, 32'hc18f96d4},
  {32'hc3fbcd08, 32'h40157693, 32'h43b9b557},
  {32'h449d19b4, 32'hc3b6b491, 32'hc2e39622},
  {32'hc3edb375, 32'h4342823e, 32'h434b8abe},
  {32'h44eb0614, 32'hc2073f93, 32'hc352260b},
  {32'hc4b7f515, 32'h42e03426, 32'h4361b3c1},
  {32'h432f1ce8, 32'hc1cb0e16, 32'hc3370a90},
  {32'hc4940fca, 32'h42136bca, 32'hc32db583},
  {32'h44ae3a2f, 32'hc196a4c4, 32'hc2a4bb11},
  {32'hc50cfcd6, 32'hc32b9d87, 32'h43366d34},
  {32'h4512f2cf, 32'hc271a188, 32'hc32c46ef},
  {32'hc46afc5a, 32'hc1b3eea1, 32'h438d8c4a},
  {32'h444d28ac, 32'hc328d48c, 32'h42f7219c},
  {32'hc49bb83a, 32'h432fd122, 32'h43030191},
  {32'h44071960, 32'hc22aa8dc, 32'hc3fe71b7},
  {32'hc3df6960, 32'h42b1f602, 32'h44013707},
  {32'h44be2f78, 32'hc3423c5b, 32'hc1c8bc9b},
  {32'hc4fc4c7c, 32'hc2f701ba, 32'hc10ade65},
  {32'h444cacac, 32'h43130bcc, 32'hc32cf699},
  {32'h4446201b, 32'hc350e5f9, 32'h4367b3bb},
  {32'hc4f6d715, 32'h437ff120, 32'hc3853425},
  {32'h44c48324, 32'h42d4ba38, 32'h4284b1b0},
  {32'hc2ffefa6, 32'hc345aede, 32'h4344356a},
  {32'h44c1cef8, 32'hc3a44efe, 32'h41d29f72},
  {32'hc41f5870, 32'hc2ba1eb9, 32'hc30fc09d},
  {32'h440dc051, 32'h4353bb89, 32'hc3b17db6},
  {32'hc4ee1d49, 32'hc34d59a4, 32'hc35744ea},
  {32'h4454e5ed, 32'h43a5bc22, 32'hc396de2c},
  {32'hc4f5f1c8, 32'hc32f1412, 32'h428ef3ef},
  {32'h44cd6d3a, 32'h423c6d10, 32'hc2a060eb},
  {32'hc517da0f, 32'hc1a2a72b, 32'h418bbca9},
  {32'h441d07b6, 32'h43881e30, 32'hc339736b},
  {32'hc50900f0, 32'hc2fa9393, 32'h429ff85d},
  {32'h44c8eb0e, 32'hc3183881, 32'hc3a5cff0},
  {32'hc38056e1, 32'hc3ad0c96, 32'h42c67c65},
  {32'h44769f8e, 32'h42fc3d52, 32'hc3c31fc2},
  {32'hc3ceb7b7, 32'hc3cf8ca5, 32'hc2b04ee5},
  {32'h44def178, 32'h41d5dc8a, 32'h43780e47},
  {32'hc4c0e073, 32'hc38c4fe4, 32'h437bcb17},
  {32'h44ede99b, 32'hc285e3d7, 32'h43766056},
  {32'hc41d0a1a, 32'hc39dedc6, 32'h42a3dad3},
  {32'h4452356d, 32'hc28eb925, 32'hc3da8ac2},
  {32'hc3b61630, 32'hc3e77af1, 32'h43fc8f86},
  {32'h43c63600, 32'h4339a0d6, 32'hc2c232e4},
  {32'hc47ed954, 32'hc2e41344, 32'h42f69ae5},
  {32'h44290954, 32'hc35a958e, 32'hc34d2c30},
  {32'hc394a3e0, 32'hc2101112, 32'hc3d87e4c},
  {32'h44e78996, 32'h418a9302, 32'h43b0ba1b},
  {32'hc4b9040c, 32'h43727ac0, 32'h433b0c0a},
  {32'h4468a9d6, 32'hc2ed0402, 32'hc2833a1d},
  {32'hc4e81ef3, 32'hc22dd54d, 32'hc1dd755b},
  {32'h44b5146e, 32'h3f0172a0, 32'hc31e88c3},
  {32'hc502df99, 32'hc3a7f8ff, 32'hc2e79732},
  {32'h44cb35e8, 32'hc2f64ec3, 32'hc360bec0},
  {32'hc48db5b7, 32'hc28546ca, 32'h43c68fd8},
  {32'h45012d96, 32'h43729357, 32'hc2cc2538},
  {32'hc519c2b5, 32'h436e84d4, 32'hc30f68ce},
  {32'h44b8b334, 32'hc245248c, 32'hc2a649f0},
  {32'hc528a0b6, 32'h429c3ac7, 32'hc3a63814},
  {32'h43fc4f0e, 32'hc31df1ee, 32'hc38977fe},
  {32'hc495439a, 32'hc28fd536, 32'hc3c3c1a8},
  {32'h44364eae, 32'h42785101, 32'h4309fb9d},
  {32'hc4bc31a6, 32'hc36d47dc, 32'hc39936e4},
  {32'h44f3297a, 32'h42ebad08, 32'h43242b70},
  {32'hc3b43114, 32'h434e5062, 32'hc36c153f},
  {32'h45043afd, 32'hc1d61410, 32'h4185f084},
  {32'hc4884be3, 32'hc2e21edd, 32'hc23037c2},
  {32'h441579f6, 32'hc36bd9c6, 32'h43a5de18},
  {32'hc475912e, 32'h42f0f2de, 32'h42f14969},
  {32'h4435b4d0, 32'h41aa0fac, 32'hc3910729},
  {32'hc24fd4c0, 32'hc1efeaf4, 32'hc262cb8c},
  {32'h451e4699, 32'hc35987f6, 32'hc2b1292a},
  {32'hc45c7914, 32'h42c69ef9, 32'hc3ba785e},
  {32'h3f79ac00, 32'h424e1f60, 32'hc35c9c74},
  {32'hc4b3b3be, 32'hc10b42b2, 32'hc41e7c4e},
  {32'h438cc9e4, 32'h431e46fb, 32'h43827658},
  {32'hc3d60a74, 32'h40cde35c, 32'h4012463c},
  {32'h45197522, 32'hc2b2393b, 32'h43251987},
  {32'hc4bbd2db, 32'h438992cd, 32'hc3519367},
  {32'h4512bf29, 32'h431bf762, 32'hc3d9d515},
  {32'hc447e4fa, 32'h43867d5f, 32'h418382e7},
  {32'h442763dd, 32'h430b6044, 32'h44052558},
  {32'hc50789f4, 32'hc37bf297, 32'hc264af66},
  {32'h44633c0a, 32'h425fb15d, 32'hc38fe03e},
  {32'hc448b686, 32'h43a07c49, 32'h4413a3ae},
  {32'h4514cfdc, 32'h430cce85, 32'hc3a3be1f},
  {32'hc49d8e37, 32'hc383f115, 32'hc382be3c},
  {32'h44e5f53e, 32'hc3916513, 32'h42761bd0},
  {32'hc4aecf5a, 32'hc27e56a2, 32'hc3340ec0},
  {32'h44abc197, 32'h438965b0, 32'h42e791b1},
  {32'hc488808f, 32'hc3b1ca94, 32'h43207525},
  {32'h44060b6e, 32'h42d44c89, 32'hc295c8e3},
  {32'hc32aa168, 32'h419f5021, 32'h418c24be},
  {32'h45052610, 32'h432c5c28, 32'h431f426a},
  {32'hc452415b, 32'h43df2410, 32'hc266601b},
  {32'h43f0cd4c, 32'h4294d6ea, 32'hc33d03bc},
  {32'hc4f2edfd, 32'h43a36ce4, 32'h432058a7},
  {32'h45000f34, 32'h42080919, 32'hc29b0b4a},
  {32'hc509afee, 32'h4203a346, 32'h432a8be6},
  {32'h431870d4, 32'h4393644d, 32'h43495b87},
  {32'hc5264424, 32'h41c0ece1, 32'hc2bf5784},
  {32'h4409ae9c, 32'h42b96ab9, 32'h43a21fe5},
  {32'hc50b31d2, 32'hc2fc569e, 32'hc342c578},
  {32'h44ce308a, 32'h42be95b4, 32'hc3877734},
  {32'hc4e3ba0d, 32'hc33d5dbd, 32'h40077f1c},
  {32'h44042014, 32'hc3049173, 32'hc2e455e9},
  {32'hc4b6079e, 32'hc2aa866a, 32'hc330f516},
  {32'h44b48aec, 32'h41bef38d, 32'h42aaf302},
  {32'hc44a94ae, 32'h42ce9686, 32'h41c75942},
  {32'h4439ec82, 32'h43d82a74, 32'h407de9a4},
  {32'hc306f3e5, 32'hc3c58ab3, 32'h42a40466},
  {32'h43c91917, 32'h4345b2c2, 32'hc2bf5b85},
  {32'hc3fce1c8, 32'hc268136a, 32'h423969bd},
  {32'h44ffc5f7, 32'h4352acac, 32'hc3673a70},
  {32'hc49b1028, 32'hc3261c1e, 32'h438ba99a},
  {32'h4486efad, 32'hc3406b97, 32'h43b674f0},
  {32'hc4c7c5f2, 32'h42bae3ff, 32'h40c2565c},
  {32'h44f4ae22, 32'hc3654edc, 32'h42748f8c},
  {32'hc429a883, 32'hc358ae73, 32'h432440e7},
  {32'h44d143d8, 32'h437bf056, 32'hc337c5e5},
  {32'hc443349a, 32'hc2db06f1, 32'h413424b2},
  {32'h43b2a1a8, 32'h4378ef89, 32'hc3c0f956},
  {32'hc4c85098, 32'h42c9fca2, 32'h42b05b52},
  {32'h44eedfd4, 32'hc409dbd8, 32'hc1d77518},
  {32'hc4351a21, 32'h418aa086, 32'h4321dd29},
  {32'h4508b62a, 32'hc264e17c, 32'hc3285071},
  {32'hc48d1184, 32'hc3bfd879, 32'h4314d38f},
  {32'h43690450, 32'hc283614e, 32'hc0f5df70},
  {32'hc53ddcd8, 32'hc2fd9b2e, 32'hc385ab78},
  {32'h43527da0, 32'hc2ddd1ff, 32'h41a7fd6c},
  {32'hc4d16b0e, 32'h428d58dc, 32'h436ab6f6},
  {32'h45104dd6, 32'h43716808, 32'h428d6f8b},
  {32'hc5099f6b, 32'hc3055a75, 32'hc19996a5},
  {32'h451e54f4, 32'h411f8670, 32'hc223529e},
  {32'hc3f42c00, 32'h40003090, 32'hc21cf89e},
  {32'hc2e7e3d0, 32'h4082c6c7, 32'h43693926},
  {32'hc3c41948, 32'hc3209466, 32'hc1dc93c5},
  {32'h4368a738, 32'hc2e84d02, 32'hc1cfec07},
  {32'hc498d3d1, 32'hc24b2762, 32'h43a6c059},
  {32'h450df240, 32'hc2ea57bd, 32'h438b887c},
  {32'hc46ac9f6, 32'hc2705951, 32'hc247c2a9},
  {32'h44f84681, 32'hc32120f6, 32'h43932c3b},
  {32'hc49f50ea, 32'hc2dc1644, 32'h4376da14},
  {32'h440299b7, 32'h431ed321, 32'hc2817e05},
  {32'hc4e5ca6e, 32'hc29eb230, 32'hc2ea2a44},
  {32'h43b18ea8, 32'h43acd052, 32'h42f813d5},
  {32'hc4b3280f, 32'h42f34aee, 32'hc3fdafb4},
  {32'h43e5fb94, 32'h42f48e4b, 32'hc1a58d82},
  {32'hc4ebfc6b, 32'h43c2d0a4, 32'h435e9dc1},
  {32'h44f87188, 32'hc2e41834, 32'h43442b88},
  {32'hc47a72ae, 32'h41a73daa, 32'hc36e613c},
  {32'h4508f7b5, 32'hc30e6468, 32'hc307f112},
  {32'hc4c189e8, 32'hc2eb0de4, 32'hc30c24d4},
  {32'h449eea09, 32'h441d4efe, 32'h42ad52b3},
  {32'hc45159bb, 32'hc346c790, 32'hc359a104},
  {32'h44f6c3d1, 32'hc3abe2ff, 32'h427afc2d},
  {32'hc49e7b51, 32'hc1a223f0, 32'h4275d996},
  {32'h4492a766, 32'hc3a44d42, 32'hc1eccd2c},
  {32'hc4d7a4ed, 32'h43d389c3, 32'h4282ab4e},
  {32'h4475979c, 32'hc32fac51, 32'hc30a22ad},
  {32'hc420abb0, 32'hc3922a79, 32'hc2deedde},
  {32'h44f46970, 32'hc1bb5bb4, 32'h41f38b9e},
  {32'hc4bdc23c, 32'hc3ab064e, 32'h4247a754},
  {32'h44b52c1d, 32'h43a670df, 32'hc2873bb0},
  {32'h42988852, 32'hc31c1051, 32'hc402a10c},
  {32'h43f8ded6, 32'hc3e46944, 32'h41d7f1cc},
  {32'hc50bea1a, 32'h431f650a, 32'h42a990a1},
  {32'h44bcc201, 32'hc2a1a05b, 32'h42b69c1f},
  {32'hc48801e9, 32'h436d51be, 32'h430e7243},
  {32'h4500322a, 32'h434a4b4e, 32'h4287606e},
  {32'hc4efbf1c, 32'hc370524a, 32'h433e2416},
  {32'h44e1633f, 32'hc313e760, 32'hc36b786c},
  {32'hc4c9af09, 32'hc305a856, 32'h43c2335f},
  {32'hc2bb4888, 32'h41a05cb4, 32'h41b9d3db},
  {32'h43119200, 32'h427381a8, 32'h432c9c63},
  {32'h44e57a49, 32'hc337012a, 32'h43133149},
  {32'hc3bfce36, 32'h42da25df, 32'h41e908ed},
  {32'h44d1af16, 32'hc127c2d6, 32'h42a33a07},
  {32'hc4afdcaa, 32'hc391cbad, 32'hc299dcb8},
  {32'h448e2e82, 32'h42c426ae, 32'hc218e7f9},
  {32'hc3261710, 32'h42ca8e8e, 32'hc3ce9e44},
  {32'h431ce4a0, 32'h435e5130, 32'hc3106324},
  {32'hc3c175a2, 32'h4395aa6e, 32'h42ae0d30},
  {32'h4508695e, 32'h43c4368f, 32'h43f1cf7c},
  {32'hc4dcde66, 32'h4340c155, 32'hc27e5600},
  {32'h44ef87fa, 32'hc2fdc27d, 32'hc3469c03},
  {32'hc4455b7a, 32'h41eb862a, 32'h434b6098},
  {32'h44fa03e1, 32'hc34ad1c9, 32'h42985e04},
  {32'hc4fe5c28, 32'hc3247d4a, 32'h437ce415},
  {32'h446f24bf, 32'h42593541, 32'hc2c1d728},
  {32'hc3ff9330, 32'h43806ca9, 32'hc318ebe2},
  {32'h44ccf8c5, 32'hc3bdfca0, 32'hc3078f70},
  {32'hc507ab67, 32'h432e7eda, 32'hc38cb5c4},
  {32'h45162f2e, 32'hc18a4c8c, 32'h419065a0},
  {32'hc4a9c25f, 32'h4389e412, 32'hc3869c14},
  {32'h44f5c434, 32'h419c5d59, 32'h3fabbb68},
  {32'hc4273518, 32'hc3c3ee1f, 32'h42cde91d},
  {32'h437f36f0, 32'hc319cb2b, 32'h441607e3},
  {32'hc50fd7f4, 32'h42ca09a4, 32'hc3377166},
  {32'h448cdc3e, 32'hc2f66c27, 32'hc309b8b3},
  {32'hc1cd87c0, 32'hc2bb1161, 32'hc34820b8},
  {32'h44fc5603, 32'h420a69a6, 32'h43017689},
  {32'hc416ab28, 32'h428871b7, 32'h437fbdd2},
  {32'h43da8071, 32'hc25ac05f, 32'hc2f60ef9},
  {32'hc5027d28, 32'hc2812f14, 32'hc2b54172},
  {32'h44c2ea1a, 32'hc3e3a26f, 32'hc31352ef},
  {32'h43051868, 32'hc324347c, 32'hc2f2849a},
  {32'h44c6c1c0, 32'hc18f3f2b, 32'hc33a6339},
  {32'hc4adde2a, 32'h4319987c, 32'hc2c1e10f},
  {32'hc33b44f8, 32'h43612b2d, 32'h435df157},
  {32'hc3edcf30, 32'hc02fc14c, 32'h420d40c6},
  {32'h43a1cff0, 32'hc2c8fafe, 32'hc2d1685a},
  {32'hc48b0179, 32'hc398b319, 32'hc358b1ac},
  {32'h450428b4, 32'hc30df943, 32'hc262b55c},
  {32'hc4c66959, 32'h420412f7, 32'h43db2807},
  {32'h4507a04b, 32'h4377735e, 32'h41ee7ae2},
  {32'hc4c4048c, 32'hc3288ea2, 32'hc2d5fdb4},
  {32'h44b79f30, 32'hc33f7fde, 32'h43c75d75},
  {32'hc38f913a, 32'h4382d4f6, 32'h437a61be},
  {32'h44778620, 32'h42e24fea, 32'h42f5ae6c},
  {32'hc4f14bb8, 32'hc316f474, 32'h4306dbea},
  {32'h446d4f7f, 32'h42524299, 32'h42d06bcb},
  {32'hc50ede51, 32'h4231a085, 32'h41a8fc63},
  {32'h44173396, 32'h4304aa36, 32'hc2c86b8d},
  {32'h42ebb6e0, 32'hc2118194, 32'h43e35c0d},
  {32'h44ea209a, 32'hc124d8ac, 32'h41ca7d0d},
  {32'hc4d8afc8, 32'hc343cd75, 32'hc383e5a9},
  {32'h451fa12d, 32'hc10e26f8, 32'hc34dc512},
  {32'hc3b18c3e, 32'hc37a1122, 32'h439f5c9b},
  {32'h4422e9fc, 32'h43628a8f, 32'hc172adbc},
  {32'hc493ca46, 32'hc34b0f8f, 32'h4368338a},
  {32'h44c0227c, 32'hc2df6065, 32'hc00bd03b},
  {32'hc29a1627, 32'hc38d7dce, 32'hc3066ae2},
  {32'h43d6b478, 32'h43a551ca, 32'hc29e750c},
  {32'hc4eb7670, 32'hc3ced7c9, 32'hc29dafb5},
  {32'h44b1ed1a, 32'hc28acaa6, 32'hc415f533},
  {32'hc493873d, 32'hc28d3db1, 32'h4286040e},
  {32'h44f1a863, 32'hc2548791, 32'h41122ced},
  {32'hc4191fc9, 32'hc21ab2dc, 32'h4301dc08},
  {32'h4486a971, 32'hc3cf4d0d, 32'h4318e627},
  {32'hc48035ec, 32'h43aaaeaf, 32'h4224ca36},
  {32'h44fd0ff8, 32'hc39f2cde, 32'hc1af3056},
  {32'hc4caec14, 32'h424847b5, 32'hc32af843},
  {32'h4505b058, 32'h42da5f56, 32'h43eb9acf},
  {32'hc31c397e, 32'h4385e280, 32'h42b45302},
  {32'h44d97f7d, 32'h4286bb00, 32'h43252762},
  {32'hc4b70df9, 32'hc34d8aa9, 32'hc3a69a4a},
  {32'h44b19881, 32'hc343c321, 32'h437160e4},
  {32'hc480d652, 32'hc2bdeeb5, 32'hc3326bd1},
  {32'h44f0b1f3, 32'h436db015, 32'h4283968d},
  {32'hc4f78d99, 32'h42c974ba, 32'hc3055a6e},
  {32'h4435633a, 32'h4388d753, 32'hc34381f7},
  {32'hc4eb187a, 32'hbff10890, 32'hc1fbe73d},
  {32'h4514bf0c, 32'hc386ae84, 32'hc28327d0},
  {32'hc4069f08, 32'hc29e76ca, 32'h42e26d33},
  {32'h44a89fc7, 32'hc32221a6, 32'hc34e45a0},
  {32'hc43a3b80, 32'hc36a2286, 32'hbfacb1e4},
  {32'h44a5aebc, 32'hc39c0aad, 32'hc31e8cd0},
  {32'hc3a96278, 32'h43875920, 32'h434803e0},
  {32'h44a0515a, 32'h42b551f0, 32'h42d83204},
  {32'hc4f72537, 32'h4332ca26, 32'h428e38b4},
  {32'h448a46e1, 32'h43891c35, 32'hc2e8403f},
  {32'hc4845a40, 32'h43234de7, 32'h4185a4b9},
  {32'h446ff348, 32'hc3011def, 32'h4322210d},
  {32'hc4e8ba33, 32'h4284cdb0, 32'hc3d84a79},
  {32'h448a22a1, 32'h43cfd533, 32'h413b56b6},
  {32'hc489b494, 32'hc385adee, 32'h43142787},
  {32'h44a8b6ec, 32'h43b21b89, 32'hc3c3b0fc},
  {32'hc43004fb, 32'h4183df5d, 32'hc1979850},
  {32'h413e1a00, 32'h420a45b9, 32'hc1dc46bc},
  {32'hc4bef5d6, 32'h421c46c3, 32'h426167cd},
  {32'h4504e663, 32'h438b1bac, 32'hc3cf5836},
  {32'hc379beb5, 32'h43913372, 32'hc2ea6416},
  {32'h4467cf59, 32'hc313d4ff, 32'h43083b52},
  {32'hc4f57b41, 32'hc272fe24, 32'hc33ae466},
  {32'h449f01aa, 32'h40cbdb4e, 32'hc3906652},
  {32'hc4b1a4ac, 32'hc277ef52, 32'hc2b034d2},
  {32'h44d8b99d, 32'hc39493f7, 32'hc30b2d29},
  {32'hc4c96abd, 32'hc34cd0db, 32'hc1d918ff},
  {32'h43f65244, 32'hc4162b21, 32'h42c9e6aa},
  {32'hc46ff317, 32'h43a44680, 32'h43b8b469},
  {32'h4483027e, 32'hc32d7adf, 32'hc3b39274},
  {32'hc50231dc, 32'h425adb72, 32'h436b44b8},
  {32'h4443b5dc, 32'hc307c71d, 32'h43569c29},
  {32'hc4c6be8e, 32'hc35daaa5, 32'h42e374d5},
  {32'h449e415f, 32'hc1dd9b95, 32'hc3e85c10},
  {32'hc5160a7d, 32'hc1dfb11a, 32'h429cd0e0},
  {32'h44634f27, 32'h43cb61d6, 32'h42c019a0},
  {32'hc4c4b737, 32'h432a3926, 32'hc1baf219},
  {32'h44f851a0, 32'hc3456c0c, 32'h42d87098},
  {32'hc3585200, 32'hc3518979, 32'hc2b7a35f},
  {32'h448cc96e, 32'h40f914ea, 32'hc2411a00},
  {32'hc4fe2c46, 32'hc3aeea90, 32'h410eb397},
  {32'h44101a87, 32'hc1b0fde9, 32'hc3eebeb1},
  {32'hc4739efc, 32'hc40a4424, 32'hc37b0456},
  {32'h44b914e5, 32'hc28ccf52, 32'hc31ab4ce},
  {32'hc4a3ea41, 32'hc376f293, 32'hc125436c},
  {32'h44917e7f, 32'h42a8aad7, 32'hc2ee061d},
  {32'hc432e7e8, 32'hc21074d7, 32'hc1940b8f},
  {32'h44f31688, 32'hc3021333, 32'hc32fc530},
  {32'hc45ded0b, 32'hc350bef4, 32'h434826b5},
  {32'h441f446a, 32'hc3495e47, 32'h438a247b},
  {32'hc4b8c13a, 32'h438ff4c1, 32'hc194fc32},
  {32'h42550f70, 32'h4304e991, 32'hc2d58744},
  {32'hc3e00f04, 32'hc35084c3, 32'h4363d832},
  {32'h442a0fa5, 32'hc13d23d6, 32'hc206dff5},
  {32'hc5106fad, 32'hc2d03d3b, 32'h428d25d1},
  {32'h448e1ffb, 32'hc35d06d0, 32'h42a44a8e},
  {32'hc418941d, 32'h4321bdae, 32'h4396a639},
  {32'h44e796ea, 32'h42e3b23b, 32'hc3d95527},
  {32'hc48ca4ff, 32'h43115117, 32'h444aa78f},
  {32'h44c2e740, 32'hc125623c, 32'h418812d8},
  {32'hc51a5c42, 32'hc22bbf3e, 32'h42a7ce08},
  {32'h4508865d, 32'h4392c30a, 32'hc31f9087},
  {32'hc43f0926, 32'hc31d729c, 32'hc3ad27fa},
  {32'h449a2ef4, 32'hc31404a1, 32'h4272aef2},
  {32'hc50c61fa, 32'h4331a1bc, 32'h4384628d},
  {32'h44e65413, 32'hc0aa0a44, 32'hc34a17b0},
  {32'hc4c01499, 32'h430d8f0b, 32'h438edf21},
  {32'h44043082, 32'hc3997979, 32'hc3b8e664},
  {32'hc4b11746, 32'hc3808419, 32'h43b9e3f8},
  {32'h44aede0e, 32'h430744c9, 32'hc287269c},
  {32'hc3bf288c, 32'hc34f4fde, 32'hc3f8569e},
  {32'h43c2cd60, 32'hc1b8b244, 32'h436e39be},
  {32'hc34e3afc, 32'h4364608d, 32'h43a5d0ec},
  {32'h44dd22fe, 32'hc147581b, 32'h42990258},
  {32'hc4f1ff20, 32'hc34599fb, 32'h44232fd2},
  {32'h43c93a78, 32'h43a99644, 32'hc280a746},
  {32'hc4f17d5a, 32'hc33f17a6, 32'h43fe76c1},
  {32'h44d64ce9, 32'hc24796da, 32'h42e68078},
  {32'hc505717e, 32'h4382425d, 32'h43dcc89b},
  {32'h44fbddc2, 32'h43354173, 32'h433a48e2},
  {32'hc50dfcdb, 32'hc2599814, 32'h43027699},
  {32'h44f3fdd1, 32'hc2c7068a, 32'h423367e7},
  {32'hc4c9ae88, 32'hc390b703, 32'h43496a3c},
  {32'h43db04dc, 32'h43094804, 32'h427e5de0},
  {32'hc4302efa, 32'h42f78def, 32'h433d390f},
  {32'h43818064, 32'h431003c8, 32'hc31b7112},
  {32'hc46b9687, 32'hc3c56224, 32'hc365fb7e},
  {32'h4509872f, 32'hc36674cf, 32'h42b0419a},
  {32'hc48e55d6, 32'hc3ac66e8, 32'hc33bc7fa},
  {32'h44f29c86, 32'hc193d9e6, 32'h426d5a45},
  {32'hc507e860, 32'hc2dbdb8e, 32'hc316b471},
  {32'h44f89fb3, 32'h421fad7b, 32'hc30b57d1},
  {32'hc508c62e, 32'h442edd0f, 32'hc40457d0},
  {32'h44db6519, 32'h42b1ef18, 32'hc3507e78},
  {32'hc4b09516, 32'h41a2a18e, 32'h430df783},
  {32'h4453738e, 32'h4282c6b0, 32'hc32b997d},
  {32'hc45a29ec, 32'hc3044716, 32'h434bd5b3},
  {32'h4457a4cd, 32'hc3619dd4, 32'h436c05be},
  {32'hc257bd40, 32'h4341d508, 32'h3f8e69c8},
  {32'h44500aac, 32'h436d0518, 32'hc37929d6},
  {32'hc4a68f65, 32'hc1a61c75, 32'hc33bd03c},
  {32'h45066181, 32'h43541948, 32'h4387417a},
  {32'hc4bedd75, 32'hc3575364, 32'hc33ae44d},
  {32'h43c1d1b2, 32'h420f3cf6, 32'h409335a4},
  {32'hc3b7226a, 32'hc33e2a62, 32'hc1fe9cce},
  {32'h44ed3d7e, 32'h4321c403, 32'hc061fe74},
  {32'hc410cd0d, 32'h42974666, 32'h41704418},
  {32'h451447df, 32'h424efa4b, 32'hc31e193e},
  {32'hc2286900, 32'h43921878, 32'hc3df25e8},
  {32'h42dd26ac, 32'hc2373cbc, 32'h42d04ca9},
  {32'hc3aa52a4, 32'hc348047c, 32'h42d47d34},
  {32'h444ed290, 32'h43aa6c13, 32'hc3fd661a},
  {32'hc50d6802, 32'hc3832a40, 32'hc1965a71},
  {32'h4506b070, 32'hc2c92743, 32'hc3526c95},
  {32'hc51bb136, 32'h43d0befa, 32'h4317430a},
  {32'h450a3a04, 32'h43b96278, 32'hc3b20f46},
  {32'hc4a09640, 32'h42aedef3, 32'h42d6d93d},
  {32'h42de6730, 32'hc2ff332c, 32'h41c207bc},
  {32'hc4d80166, 32'h438d8419, 32'hc2327e9d},
  {32'h451a5fb1, 32'h4235a1e6, 32'hbff78932},
  {32'hc4be4f50, 32'hc2d7c794, 32'hc37838d3},
  {32'h432d7c62, 32'h4416bd2f, 32'hc0304ecf},
  {32'hc409f466, 32'hc2fb3d98, 32'hc304e5ad},
  {32'h442beb44, 32'hc34fd986, 32'h411f5104},
  {32'hc504bb67, 32'h40f1e9c6, 32'h43465ad1},
  {32'h44d802a1, 32'h43617cca, 32'h43b3d48a},
  {32'hc504b8fe, 32'hc33ebd89, 32'h43bde17a},
  {32'h440f7880, 32'hc32033c5, 32'h431ea486},
  {32'hc50e552a, 32'hc3b57b22, 32'hc0feb0f7},
  {32'h4482ab10, 32'h42446735, 32'h4268b868},
  {32'hc409777a, 32'hc2d487c2, 32'h4396ecec},
  {32'h44513deb, 32'hc421061e, 32'h436e409f},
  {32'hc504e831, 32'h422fcf64, 32'hc2d48d3f},
  {32'h450aba10, 32'hc207cba1, 32'h426267fc},
  {32'hc5131216, 32'hc38c3255, 32'h42866183},
  {32'h443c6830, 32'hc29f5429, 32'h4363b7fa},
  {32'hc503ed23, 32'hc39d810e, 32'hc3571149},
  {32'hc37c2bce, 32'hc2905c0d, 32'h43218afe},
  {32'hc421db2c, 32'h42b5c062, 32'hc1f52f4e},
  {32'h43efd5c0, 32'hc03f6060, 32'hc4102b88},
  {32'hc4523e9a, 32'hc0d35338, 32'h43cc72b8},
  {32'h44e39fa0, 32'hc39a09a8, 32'h4337dc60},
  {32'h4211c620, 32'hc36f832d, 32'h423049cc},
  {32'h441d1110, 32'h432a2f19, 32'hc3378247},
  {32'hc4b15aff, 32'h43d64df9, 32'hc3aa9f24},
  {32'h44078034, 32'h42ab508b, 32'h433d878d},
  {32'hc457df90, 32'h4209ff67, 32'h41161190},
  {32'h4510719a, 32'hc2e28606, 32'hc3084aba},
  {32'hc502ce70, 32'hc32a7454, 32'h42f073d4},
  {32'h445d0a4d, 32'h42c3698c, 32'h42a1fedc},
  {32'hc42d0f64, 32'hc3c48373, 32'hc37fcb64},
  {32'h43413b10, 32'h43270670, 32'h434b738c},
  {32'hc4f02754, 32'hc307d736, 32'hc19087c0},
  {32'h450cd811, 32'hc2ed1265, 32'h41a65e80},
  {32'hc423e117, 32'hc3c58887, 32'h433b4b95},
  {32'h4480c17c, 32'h4376e41a, 32'h40fe836d},
  {32'hc4da4338, 32'hc28d2bf4, 32'hc34d31fe},
  {32'h44fd83fa, 32'hc2f67294, 32'h4260e1d0},
  {32'hc38c5094, 32'hc3c2b22e, 32'hc30a7e97},
  {32'h4468f0b2, 32'h441b8aba, 32'hc34aeffb},
  {32'hc501a5ba, 32'h435e01de, 32'hc3374f59},
  {32'h43cebd1a, 32'h43423287, 32'hc28df300},
  {32'hc46c5dba, 32'hc2428e15, 32'hc392167f},
  {32'h44afa01e, 32'hc10a0ad9, 32'hc332705a},
  {32'hc3aba8f0, 32'h42b793b2, 32'h4341b3aa},
  {32'h44eeb3b6, 32'h426f0d3a, 32'hc340e685},
  {32'hc3428f4a, 32'hc310acf2, 32'hc3d22ebe},
  {32'h44e54b7b, 32'hc31d1993, 32'h43984e8c},
  {32'hc50bd220, 32'h4291d7ca, 32'hc34dd24e},
  {32'h44b041c2, 32'h4325d359, 32'hc3930972},
  {32'hc313caf0, 32'h43967ba8, 32'hc2d1f75e},
  {32'h4488cfdc, 32'h436dad21, 32'h4317392c},
  {32'hc4a1ad24, 32'hc3831a4e, 32'hc282db53},
  {32'h44844346, 32'hc42f67da, 32'hc2b5fa51},
  {32'hc4653107, 32'h4318f06c, 32'hc32b36f9},
  {32'h45039d9f, 32'hc307dd11, 32'h426b875b},
  {32'hc420f983, 32'h437a0520, 32'hc3a1419e},
  {32'h44d5045e, 32'hc3e201dc, 32'hc2204d84},
  {32'hc48c7a94, 32'hc345f85a, 32'h4193286e},
  {32'h44a0edc8, 32'h430b1b7a, 32'hc298bcad},
  {32'hc258d947, 32'hc2cdf419, 32'h43ca636e},
  {32'h43d2df74, 32'hc348844b, 32'h43dc1046},
  {32'hc4defbb3, 32'hc38875c9, 32'h41b79119},
  {32'h441e18bc, 32'hc2364af5, 32'h428146e1},
  {32'hc5052e5f, 32'h4383894a, 32'hc327ba91},
  {32'h450af6ce, 32'hc3c6079a, 32'h43901c1a},
  {32'hc4b59a2f, 32'hc3221c4e, 32'hc35947f1},
  {32'h43843cd4, 32'hc2158baf, 32'hc2106f11},
  {32'h43cef6d4, 32'h41b4a8d8, 32'hc38c31c0},
  {32'h44e48ec5, 32'h431caffe, 32'hc2e29476},
  {32'hc41a17ce, 32'hc35f86f9, 32'hc3a27b57},
  {32'h42e0d0e0, 32'hc321fe09, 32'h43d8a52e},
  {32'hc4167e02, 32'hc18f5bf2, 32'hc3c2d114},
  {32'h439f8888, 32'hc226c48f, 32'hc35e01a4},
  {32'hc4aeb13e, 32'hc3bafbc9, 32'h41e46013},
  {32'h44effdc7, 32'h43403479, 32'h41b208fe},
  {32'hc363fd12, 32'hc3894e11, 32'h424a30fe},
  {32'h4468002d, 32'h43070206, 32'hc3326cb9},
  {32'hc4c17ffe, 32'hc3acc5c8, 32'hc2a90442},
  {32'hc3ee4980, 32'hc2a5291c, 32'hc2c323e9},
  {32'h44217b4a, 32'hc23e5fc4, 32'h431dce6e},
  {32'hc45b6b32, 32'h42f54939, 32'hc3a9c247},
  {32'h44af6546, 32'h426832bd, 32'h41d7dfae},
  {32'hc4be361b, 32'hc28dfe8d, 32'hc2ae6a1f},
  {32'h441d32ef, 32'h439a97c4, 32'hc305ec78},
  {32'hc439fbfc, 32'hc33f6761, 32'h43e34db7},
  {32'h44788d54, 32'h437bd777, 32'h4355aa00},
  {32'hc4897767, 32'h43569e1b, 32'h422a9a04},
  {32'h44ef354e, 32'hc39d837b, 32'h431ab865},
  {32'hc503c5e5, 32'hc25790c6, 32'hc2d98380},
  {32'h44ca2b64, 32'h42237e4f, 32'hc209a5c4},
  {32'hc47f59e0, 32'h43c4293a, 32'hc21732f7},
  {32'h4514a796, 32'h421c1437, 32'h437254da},
  {32'hc49bbf77, 32'hc3ea4150, 32'h42a40709},
  {32'h44e230b2, 32'h42cbe655, 32'hc36bf649},
  {32'hc35af3c0, 32'h439d346d, 32'hc33bf3e9},
  {32'h451c02c7, 32'h43c0b707, 32'hc32f28bd},
  {32'hc3a0f190, 32'h43af240a, 32'hc3f2c90b},
  {32'h449111d2, 32'h41729c90, 32'h44048e49},
  {32'hc4633cf9, 32'h439adca1, 32'hc3a34825},
  {32'h43a96fca, 32'hc28b17cd, 32'hc3527424},
  {32'hc34f5618, 32'hc30f8779, 32'hc283cdf1},
  {32'h45118b7f, 32'hc24482c8, 32'hc2c62dba},
  {32'hc3d36b44, 32'hc3061b38, 32'hc0211e28},
  {32'h43cf25d8, 32'hc2ee08f8, 32'h4333b41a},
  {32'hc3ec78c3, 32'h42eccfaf, 32'hc28c4f37},
  {32'h4506e303, 32'h432612a4, 32'h42be9cbf},
  {32'hc50c7475, 32'h43170ee2, 32'hc394d551},
  {32'h44e8967e, 32'hc30c38fd, 32'h42d1c875},
  {32'hc37893d3, 32'h4295c0d6, 32'hc37ddc4e},
  {32'h44f83054, 32'h4210273f, 32'h44073606},
  {32'hc50645c8, 32'h41ddf4c0, 32'h4385efbd},
  {32'h4428fa23, 32'h43661f5d, 32'hc2fb7162},
  {32'hc380bb10, 32'hc35fa9bb, 32'hc371b2b0},
  {32'h44ce7f7c, 32'h438cc683, 32'hc2631179},
  {32'hc412598a, 32'h42f9587f, 32'hc414046a},
  {32'h44e5494b, 32'h435872dc, 32'h432bf7d9},
  {32'h42dd1c00, 32'hc33fd55f, 32'hc3078253},
  {32'h449a7c61, 32'h4335e807, 32'hc3870966},
  {32'hc3552852, 32'hc29df7b8, 32'h41ac0c5c},
  {32'h451d3158, 32'h43252b3f, 32'hc2a24bdf},
  {32'hc43a7918, 32'hc0f7a781, 32'hc3c2da3f},
  {32'h44e03b36, 32'hc29a54f0, 32'h42c0905b},
  {32'hc4821b3d, 32'h42cff22e, 32'h41faf002},
  {32'h444b24c2, 32'h422116de, 32'h42c0ed0e},
  {32'hc508bbf3, 32'h42873414, 32'h437aed10},
  {32'h44cf3170, 32'hc1b3604a, 32'h43fb3242},
  {32'hc4870922, 32'h43d99fbe, 32'hc2c307ab},
  {32'h44d9eaa5, 32'hc3a9626f, 32'h42dd04d4},
  {32'h434bf4c7, 32'h432dcaea, 32'hc3a15cb4},
  {32'h437b5988, 32'h41bb27c1, 32'hc351abb4},
  {32'hc4a300fc, 32'hc2772f2e, 32'hc38bd347},
  {32'h44c14156, 32'hc211a9d5, 32'h42bf1d97},
  {32'hc41c9eae, 32'hc2a99562, 32'h427dbbe4},
  {32'h42c83774, 32'hc34896c4, 32'hc40f7f72},
  {32'hc4cf4873, 32'hc383ee25, 32'hc1f05d1f},
  {32'h44dd920e, 32'hc1fd3929, 32'hc4097dde},
  {32'hc3c4e098, 32'h4309b6ae, 32'hc3b46eee},
  {32'h43806db8, 32'hc30815de, 32'h43cf0dd2},
  {32'hc4b70c70, 32'h431d366a, 32'h42fe0048},
  {32'h44d63518, 32'hc305d7a6, 32'h43ef9771},
  {32'hc4e1e086, 32'h433546f6, 32'hc357709b},
  {32'h4449ba64, 32'h40d996aa, 32'h41e7ca18},
  {32'hc4f6aad0, 32'hc3a08720, 32'h4280701e},
  {32'h447885d6, 32'hc3a22373, 32'h41e347f5},
  {32'hc4be5bb7, 32'h41b69c88, 32'h4361c744},
  {32'h451d6352, 32'h43034bcd, 32'hc1806e96},
  {32'hc50e823e, 32'hc2328abc, 32'hc32dc273},
  {32'h44792da4, 32'hbdced000, 32'h42f27f5e},
  {32'hc4dadaa3, 32'hc39d70a7, 32'h4379da5c},
  {32'h44874862, 32'h4202493b, 32'h43c7f1de},
  {32'hc380d6ec, 32'h42e5ab40, 32'hc440150e},
  {32'h44ee987a, 32'hc0387432, 32'h4285be8d},
  {32'hc4ec57d2, 32'h437beadd, 32'h4203d5d2},
  {32'hc35b7700, 32'h42317992, 32'hc3a72d87},
  {32'hc3766760, 32'hc3188d5a, 32'h43dac2ae},
  {32'h44dec34f, 32'hc311a8f2, 32'hc2544d14},
  {32'hc50c928e, 32'hc2a65565, 32'h4301dcdd},
  {32'h451cc88a, 32'h44229f0f, 32'h42e0ac72},
  {32'hc4fc1a39, 32'h43534186, 32'hc3603fef},
  {32'h448a3ce7, 32'h3ea806a2, 32'hc3117a8c},
  {32'h434d10b8, 32'hc354444b, 32'h43afa26e},
  {32'h450a4920, 32'h43b6ceb2, 32'h43576877},
  {32'hc513c054, 32'hc204d2aa, 32'hc2d17550},
  {32'h450e3e0c, 32'hc3b04d42, 32'h43d51f32},
  {32'hc4e1ba17, 32'h4321ae7f, 32'hc2e4ac9b},
  {32'h4451eaf4, 32'hc3b629e6, 32'h433b7597},
  {32'hc4df5902, 32'hc32baf42, 32'hc26ed31e},
  {32'h446f0d91, 32'hc3e94fa8, 32'hc3372994},
  {32'h436b860d, 32'hc2e29cff, 32'hc2b8ea5c},
  {32'h450973bc, 32'hc25b87e5, 32'hc30144b5},
  {32'hc4e478c8, 32'hc324705a, 32'h435fee0c},
  {32'h441c5a52, 32'hc360ca6f, 32'h43b1e92f},
  {32'hc390aee8, 32'hc07af856, 32'h42998f16},
  {32'h44114492, 32'hc37eab99, 32'h423aa645},
  {32'hc4b1178f, 32'hc380c2a4, 32'hc2beebf9},
  {32'h4506a401, 32'h431d11e3, 32'hc362d47f},
  {32'hc3343800, 32'hc345179b, 32'h4380e23c},
  {32'h44c2dde3, 32'h42ba4454, 32'h43c622b2},
  {32'hc483252f, 32'hc2dbb08d, 32'hc2a6f6cc},
  {32'h44e343d7, 32'hc3b58c97, 32'hc332041f},
  {32'hc4926b68, 32'h4389c70e, 32'h42d43b8b},
  {32'h439b7739, 32'h43810b75, 32'h437bd2f6},
  {32'h43a482b1, 32'hc3579960, 32'hc3143b74},
  {32'h44618b3b, 32'hc340ae32, 32'h41595310},
  {32'hc4528291, 32'hc3850715, 32'hc34961bf},
  {32'h44f4b36c, 32'h4343e0e6, 32'h4390cb6e},
  {32'hc4bd3416, 32'hc36b3e12, 32'h439147d1},
  {32'h451a971d, 32'h42bdbf87, 32'hc3f4708d},
  {32'hc082a700, 32'hc2971eb8, 32'hc28f027a},
  {32'h423f7f50, 32'h42ccc59d, 32'hc2297662},
  {32'hc50e437f, 32'h42fc638d, 32'h434ae361},
  {32'h44890d1e, 32'hc335c9cb, 32'hc319a40d},
  {32'hc5099ce4, 32'h434c16d5, 32'h41e91997},
  {32'h43e94c48, 32'hc3e712c3, 32'hc3cf5592},
  {32'h44831580, 32'h4243339a, 32'hc2f5e169},
  {32'hc46a77e0, 32'h435a7ea6, 32'hc29acf74},
  {32'h44e0ac96, 32'h42f1336d, 32'hc24ed228},
  {32'hc414c155, 32'h434d0aef, 32'hc1c27ab2},
  {32'h44af360f, 32'hc25149a4, 32'hc091599a},
  {32'hc511adbe, 32'hc2571a5f, 32'h4395caf5},
  {32'h450ddd40, 32'hc2c80028, 32'h42c50ec2},
  {32'hc4c2e3b7, 32'h43cd170f, 32'hc2a6b9cc},
  {32'h439eb847, 32'h43f029ec, 32'h41ddfad6},
  {32'hc4b6283d, 32'hc353cda1, 32'hc37423ac},
  {32'h44c2f4c8, 32'hc1ac880f, 32'h42ab8b81},
  {32'hc47c9a4b, 32'hc3a7a90e, 32'h435d9245},
  {32'h4503b11d, 32'h43786951, 32'hc3624a5d},
  {32'hc4bb459a, 32'h422879e3, 32'h433e003f},
  {32'h44b62e18, 32'h43113cff, 32'h43c14d56},
  {32'hc46c8535, 32'h42ee37b1, 32'h43d0a48f},
  {32'h44f416b2, 32'h42e1dcde, 32'hc1e1b144},
  {32'hc451a764, 32'hc1e598a1, 32'h43d3d2f3},
  {32'h44bfc25e, 32'hc3d37981, 32'hc37e6b16},
  {32'hc35e9b94, 32'h421bb25a, 32'h42ee8de3},
  {32'h44a82508, 32'h4347db22, 32'hc2670675},
  {32'hc4c72d23, 32'h434f5c90, 32'hc05497c0},
  {32'h450e6834, 32'h42b0d132, 32'h42939c35},
  {32'hc4f0cb58, 32'h43039e3e, 32'h4122316b},
  {32'h43ba8670, 32'hc2c6f0ec, 32'h43462f8d},
  {32'hc50de8ca, 32'hc33fc8ab, 32'h43c2a576},
  {32'h44001c20, 32'h438c2622, 32'h431654bb},
  {32'hc41365f0, 32'h431dea36, 32'h439f6bf2},
  {32'h440858c6, 32'hc2e6a2e2, 32'hc31e7778},
  {32'hc49f06f2, 32'h43476598, 32'hc39f4397},
  {32'h44673fe0, 32'h4332f4da, 32'hc22ee664},
  {32'hc487f668, 32'hc2b03e2b, 32'h42e2c5d8},
  {32'h44ec86ca, 32'h43929fc6, 32'hc30ed4bf},
  {32'hc42f9b00, 32'hc380cb96, 32'hc35004a2},
  {32'h450c061b, 32'h437bea30, 32'hc314d612},
  {32'hc488f780, 32'h431580ea, 32'hc3325452},
  {32'h44411e34, 32'hc29a6aea, 32'h4293ed95},
  {32'hc3c7b7a4, 32'hc2c49fb3, 32'hc2ad068d},
  {32'h444b0d80, 32'h43e8e0a0, 32'h432d3200},
  {32'hc46bc55a, 32'h42d57e92, 32'hc3434b98},
  {32'h44ad7909, 32'h429fd804, 32'h4377977c},
  {32'hc4243bcd, 32'h42ca0fdc, 32'hc3b74ff0},
  {32'h44f3bd42, 32'h4227bc6a, 32'hc3522da9},
  {32'hc387951c, 32'hc3b87eeb, 32'hc33e6919},
  {32'h4502f1eb, 32'h432a14a9, 32'hc31d1ee9},
  {32'hc32a7d70, 32'hc2e9e716, 32'hc31b8f71},
  {32'h4477924c, 32'h42fca937, 32'hbfea39e0},
  {32'h42527b82, 32'hc264d0a3, 32'hc31626ba},
  {32'h44ab5db0, 32'h425f24a0, 32'hc1729164},
  {32'hc4872d2c, 32'h42d6fb5a, 32'h42418884},
  {32'h43922fe4, 32'h43a861bf, 32'h42b19e46},
  {32'hc490ff26, 32'hc26a7199, 32'hc2e8c064},
  {32'h448eb45e, 32'hc2d414f9, 32'h42e53b72},
  {32'hc3c2fb38, 32'h4400eb28, 32'h43717f74},
  {32'h4386c994, 32'h43bfe3b3, 32'h422d5a31},
  {32'hc4add72c, 32'h42baa026, 32'h430fa717},
  {32'h42b93d40, 32'h42340f65, 32'h42ccaa67},
  {32'hc4fbc76a, 32'hc301251d, 32'hc2d68ff9},
  {32'h43afbfc8, 32'h4402bc5a, 32'h43e38f2c},
  {32'hc4451b76, 32'h4330981a, 32'h41a02d04},
  {32'h450496fa, 32'h435b2ce6, 32'h438d1cfc},
  {32'hc4781316, 32'h4323cfe1, 32'hc3d780dc},
  {32'h44b6e64e, 32'h41ee2c48, 32'hc3bd3bb3},
  {32'hc4b28ce5, 32'h418f005b, 32'h429b5d7a},
  {32'h44a4cfb4, 32'h429ae308, 32'hc41cc6fc},
  {32'hc34e4a00, 32'h42032742, 32'h43c4f2f5},
  {32'h44970b1b, 32'h43981aac, 32'h43360266},
  {32'hc4b194a5, 32'h42e8ac4d, 32'h4274871c},
  {32'h442dc718, 32'h4341febe, 32'hc228f4d2},
  {32'hc50b6d04, 32'hc2c87732, 32'hc334a0e3},
  {32'hc2b74b58, 32'hc367772b, 32'hc3895999},
  {32'hc3b63b52, 32'h431aa9ee, 32'h43418f3c},
  {32'h447da1fc, 32'h438f9109, 32'hc2e0a1c1},
  {32'hc460936b, 32'hc30633f1, 32'hc335ac40},
  {32'h44c7c1a2, 32'h43a9cf05, 32'h439db463},
  {32'hc4b6e973, 32'hc2e02405, 32'h43b330ac},
  {32'h44fdd8fc, 32'h436bdf9f, 32'h42652508},
  {32'hc2d97d70, 32'hc1f7c4b3, 32'h438f2667},
  {32'h44d46f18, 32'h439cffab, 32'hc31f5b8b},
  {32'hc4cf5054, 32'h4324e92c, 32'hc3274de1},
  {32'h43cc2280, 32'hc36e74e5, 32'hc2a88f78},
  {32'hc50adc98, 32'h43091d99, 32'hc306e1b5},
  {32'h44a9d40e, 32'hc33c609a, 32'h436a3fc8},
  {32'hc4b3169e, 32'hc25389f4, 32'hc2dcfc94},
  {32'h44646e00, 32'hc19963cf, 32'h43a0bb56},
  {32'hc3ec0519, 32'hc3bf7e13, 32'hc303bff1},
  {32'h4494babe, 32'h43a00437, 32'h430687b1},
  {32'hc46a1618, 32'h3e92e480, 32'h434731d4},
  {32'h44ed740d, 32'h40775412, 32'h42633074},
  {32'hc4ddecde, 32'h43c5a484, 32'hc37d8318},
  {32'h4426ba21, 32'h42ae9115, 32'h43069c9a},
  {32'hc2a9d500, 32'hbfc97146, 32'hc34a30a8},
  {32'h44a8742a, 32'hc308151a, 32'hc3e54b5e},
  {32'hc3b78278, 32'hc3e42a92, 32'hc1a8741f},
  {32'h43dd6082, 32'h4396c206, 32'hc3e675b7},
  {32'hc4159d58, 32'hc24c7b79, 32'hc3a89d2e},
  {32'h44461a64, 32'h4396deef, 32'hc32d0f9c},
  {32'hc4819678, 32'hc35cf353, 32'h42981353},
  {32'h449eb514, 32'h40c769d8, 32'h439a54c1},
  {32'hc505990a, 32'h433911b6, 32'hc2aeb462},
  {32'h448d3d43, 32'hc2fb668d, 32'h42690308},
  {32'hc50e4fa5, 32'hc28952aa, 32'h43a5d9f9},
  {32'h44638e64, 32'hc18fb25c, 32'h440d6b47},
  {32'hc4688e8c, 32'hc2d76616, 32'h436d4791},
  {32'h44c5faaf, 32'h435ef9bf, 32'hc333402a},
  {32'hc474d799, 32'h410ca89d, 32'hc2b96ef0},
  {32'h44efa070, 32'h434f26a7, 32'h422f3f9a},
  {32'hc302b670, 32'h437304a1, 32'hc3498ad5},
  {32'h42a9ce40, 32'h42788481, 32'h4295c137},
  {32'hc465b557, 32'h431454d9, 32'h42e1e942},
  {32'h43eab428, 32'hc30d068e, 32'hc382fb89},
  {32'hc4875495, 32'hc3acccff, 32'h43d72705},
  {32'h44784f74, 32'hc2a9b4e1, 32'hc3a6806e},
  {32'h435a1575, 32'h42c7d94a, 32'hc39a45e7},
  {32'h4465b43b, 32'h420fd907, 32'hc383dc87},
  {32'hc4aec456, 32'hc2ba0389, 32'hc23481c8},
  {32'h4505c032, 32'h42887037, 32'hc39d79f7},
  {32'hc507536c, 32'hc33aa1bd, 32'hc1b860ff},
  {32'h43eb7221, 32'h42c8589e, 32'h4383f066},
  {32'hc4d505dd, 32'hc283f170, 32'h40f4deae},
  {32'h44ea6cdb, 32'h42e17930, 32'h412b8b1b},
  {32'hc4dacd05, 32'hc3c0b8e9, 32'h42c126d3},
  {32'h449a491e, 32'h428acd51, 32'hc20e3ae4},
  {32'hc3b68e4c, 32'h406ae170, 32'hc28d14f6},
  {32'h449f8921, 32'h4230a5a0, 32'hc29ac077},
  {32'hc44277a4, 32'h42a9d6a0, 32'h4294ed14},
  {32'h42e9fa20, 32'h424a423e, 32'hc32287bf},
  {32'hc4a0871d, 32'h439abafc, 32'hc3cad42f},
  {32'h43c0d3e4, 32'h435fff43, 32'hc150dc52},
  {32'hc505d30d, 32'h4311697d, 32'h4330a867},
  {32'h44373918, 32'hc3100a6f, 32'hc183464c},
  {32'hc45bcb4c, 32'h4364871f, 32'hc22a673e},
  {32'h4465dc60, 32'h43ba451e, 32'hc466a500},
  {32'hc47d8ac8, 32'hc3445a7b, 32'h426cd168},
  {32'h445de4ee, 32'h4391b721, 32'h42cc7c34},
  {32'hc4c019b4, 32'hc37bc19a, 32'h42ebed97},
  {32'h444da01a, 32'h410a2f46, 32'hc2cbebf4},
  {32'hc475e998, 32'hc362e51c, 32'hc1b6880f},
  {32'h44283ca8, 32'hc38b9c43, 32'hc207b6b4},
  {32'hc41ca454, 32'hc35aadcb, 32'hc0dcc54f},
  {32'h44f0ff99, 32'h4284f307, 32'h43545bcb},
  {32'hc4b5a4f1, 32'h43b4fe4d, 32'hc2258cad},
  {32'h44f7be18, 32'h43371bc3, 32'hc38a3e48},
  {32'hc465f214, 32'hc1c56892, 32'hc33264db},
  {32'h43bede7c, 32'hc39e4029, 32'hc2c7cc3f},
  {32'h42084370, 32'h41301b5c, 32'h42c74da8},
  {32'h44a319d5, 32'h430b9f63, 32'hc1e01147},
  {32'hc4c6ea64, 32'hc345627e, 32'hc368af8c},
  {32'h44e6c570, 32'hc374ced2, 32'h435d5073},
  {32'hc45bed3a, 32'h43ada352, 32'hc3eba9bd},
  {32'h43faa614, 32'h4382abc1, 32'h4324fa76},
  {32'hc395cc00, 32'hc2beefaf, 32'h41a0f45d},
  {32'h44808ccc, 32'h43da034b, 32'h412f2adb},
  {32'hc494aa0e, 32'h41c4d397, 32'hc39504b1},
  {32'h450c1164, 32'h42824b34, 32'hc3aa5f3e},
  {32'hc4ba1dec, 32'hc206ab2c, 32'h4375cca8},
  {32'h4419eeea, 32'h4394e3d5, 32'hc3dd6a26},
  {32'hc4ee8bb2, 32'h432a6db7, 32'h4151f5da},
  {32'h44e45240, 32'hc3bedea9, 32'hc2df8e20},
  {32'hc491205f, 32'hc2215ee7, 32'h4382902d},
  {32'h4470668a, 32'hc310726c, 32'h42eec416},
  {32'hc48dcf53, 32'h43b043b8, 32'hc1d395b6},
  {32'h44ce4500, 32'h3ef230dd, 32'hc2cd172a},
  {32'hc364d1bb, 32'h42f8c915, 32'hc0b3dcb0},
  {32'h44bbb128, 32'hc2a0b313, 32'h438d05a6},
  {32'h424a9ac0, 32'h423dc6e6, 32'hc1a9ef3c},
  {32'h4487d8fd, 32'hc2c7bd88, 32'hc3ccc663},
  {32'hc503eb9e, 32'hc26f9fc3, 32'hc30fbdaa},
  {32'h450f0f45, 32'hc08b6fd0, 32'h424f4a37},
  {32'hc4286332, 32'hc2d8b69e, 32'hc2a7c2c2},
  {32'h44d7f7f2, 32'h43b61be9, 32'hc1b7c2b0},
  {32'hc41e6c5e, 32'hc305c917, 32'h42c064bf},
  {32'h448f5f59, 32'hc392c1a4, 32'h42f862be},
  {32'hc3c4bdc7, 32'hc1bdf7d0, 32'hc3a6adb4},
  {32'h440ceab8, 32'hc352abe1, 32'h41028640},
  {32'hc45e47a2, 32'h433ee936, 32'h427e17aa},
  {32'h44c427b6, 32'hc3c49a05, 32'h43954c03},
  {32'hc48b1c86, 32'hc3725ebc, 32'hc39eea47},
  {32'h44061d78, 32'h4331a53c, 32'hc2880753},
  {32'hc40bf8c0, 32'h435584a6, 32'h4406bc24},
  {32'h44251210, 32'h43f517dc, 32'hc18ed73c},
  {32'hc5024c81, 32'hc31ef0fd, 32'h438a5de6},
  {32'h447ea7c4, 32'hc2beb653, 32'hc1013546},
  {32'hc41d5406, 32'h43d5934f, 32'hc39cfb67},
  {32'h4511c185, 32'hc210a340, 32'h4167fa2a},
  {32'hc47015f8, 32'hc38cb7ca, 32'h43c1aeb6},
  {32'h44dbf7d3, 32'h432f60e9, 32'hc34fc709},
  {32'hc3a574ac, 32'h42f6ce8a, 32'hc30d47c4},
  {32'h44b80fd6, 32'h43016555, 32'h42c53a90},
  {32'hc45990c0, 32'h4041f874, 32'h4281ce74},
  {32'h4522febc, 32'h439821b9, 32'hc33eee25},
  {32'hc4cef830, 32'h43535fa0, 32'h4309834e},
  {32'h43ace084, 32'h43882d35, 32'h4397da61},
  {32'hc45248a4, 32'hc2fd9799, 32'h43839c67},
  {32'h44ed7c50, 32'h43a0d9f6, 32'h43a4b567},
  {32'hc35ab265, 32'h41a26353, 32'h432f8c5f},
  {32'h45318dd0, 32'hc2445222, 32'h43615eaa},
  {32'h426bfd40, 32'h42f0b1d2, 32'hc3b673d6},
  {32'h44885268, 32'hc0d93647, 32'h4303f841},
  {32'hc3f96169, 32'h4364b633, 32'h43c15974},
  {32'h4495cddb, 32'hc308d7f2, 32'h43bc7875},
  {32'hc3daecc2, 32'hc380112d, 32'h41dffe99},
  {32'h44941a1e, 32'hc305e6f1, 32'h3f344220},
  {32'hc40f5990, 32'h435df501, 32'hc39e6cda},
  {32'h4424df7b, 32'hc3554a73, 32'h4357c4c8},
  {32'hc502d93e, 32'h42e2ca5b, 32'hc323bb57},
  {32'h443a6bf2, 32'h43f84d44, 32'h4391cedc},
  {32'hc4e18e62, 32'h4100127b, 32'h4261a469},
  {32'h44a39e13, 32'hc40cc686, 32'h4406e5f1},
  {32'hc47d6a06, 32'h42283f33, 32'h4408056e},
  {32'h44855b60, 32'hc3435119, 32'h4397121f},
  {32'hc42433cc, 32'hc3f4e0d5, 32'h41e754b4},
  {32'h44d173c0, 32'h4190754a, 32'hc31bd3fd},
  {32'hc4f968c7, 32'hc380c444, 32'hc37419c6},
  {32'h44211a14, 32'hc309d16f, 32'hc343bc18},
  {32'hc5100c21, 32'h424bd15b, 32'hc1841575},
  {32'h450c4cde, 32'hc2104937, 32'hc33e366b},
  {32'hc5032bea, 32'hc30b8a91, 32'hc1a67300},
  {32'h44967418, 32'hc2330a70, 32'hc35ce4e2},
  {32'hc3d75f65, 32'h4338492b, 32'h41899b83},
  {32'h440c90e8, 32'h4274a9c0, 32'hc1cd80e0},
  {32'hc502b2f2, 32'h41a6da9a, 32'hc3dd0728},
  {32'h45063bf6, 32'hc32f67b2, 32'hc2c5ae82},
  {32'hc4ab8119, 32'hc308f0fa, 32'h4230e1c3},
  {32'h43c56360, 32'hc1b59dbe, 32'hc33870d4},
  {32'hc4a70b2a, 32'h43390d4b, 32'hc206708b},
  {32'h4377eccc, 32'hc335d381, 32'hc1ddeef5},
  {32'hc3239dc0, 32'h431bbf5a, 32'hc223ed0e},
  {32'h450553e6, 32'h436b7c3b, 32'h43c91de0},
  {32'hc4f06535, 32'h42562015, 32'hc382fbee},
  {32'h44bea3c4, 32'hc3002750, 32'h4306a2c7},
  {32'hc40207df, 32'h43adadb3, 32'h41ac74ba},
  {32'h44c0bd62, 32'h41e5461d, 32'hc3620425},
  {32'h43061c56, 32'hc2b73e2e, 32'hc3ace6f5},
  {32'h45018be7, 32'h4343232d, 32'h42ea4581},
  {32'hc34a859c, 32'hc310460c, 32'hc23d868e},
  {32'hc215a390, 32'h431eb6c7, 32'hc25439f0},
  {32'hc3edd218, 32'hc34f2f23, 32'h421bfaff},
  {32'h44f7c994, 32'hc4286127, 32'h42a73ef1},
  {32'hc4a37005, 32'h439bacf7, 32'hc24887af},
  {32'hc362507d, 32'h42ae68ce, 32'hc34e1852},
  {32'hc501908a, 32'hc2f886f1, 32'h426e2f9d},
  {32'h448723d2, 32'hc3100c09, 32'hc3f0b3f6},
  {32'hc4c147c8, 32'h43a68787, 32'hc2ff1c3b},
  {32'h44bc4564, 32'hc3be3316, 32'h42c4a75c},
  {32'hc33f6fc0, 32'h41e1ffa1, 32'hc2716d74},
  {32'h43046bb0, 32'h416eb44c, 32'h43180625},
  {32'hc4fe5c63, 32'h43b93f32, 32'h43955616},
  {32'h44f20000, 32'hc3582aac, 32'h4357f8c9},
  {32'h43a9b0d4, 32'hc31e920d, 32'h423898b0},
  {32'h45000b82, 32'h428b2b15, 32'hc38a8f31},
  {32'hc5189198, 32'h43987124, 32'h425ddff6},
  {32'h42c4dd1c, 32'h43851139, 32'h43a7b856},
  {32'hc497639a, 32'h425d53da, 32'h43a5c0c4},
  {32'h44ad9fe6, 32'h41996fe6, 32'hc2e97429},
  {32'hc48ca32d, 32'h4384391d, 32'hc3b1e252},
  {32'h45077dab, 32'hc3404566, 32'h4241119f},
  {32'hc5062e38, 32'hc39e1899, 32'hc3cc96c1},
  {32'h439cc841, 32'h4285172e, 32'hc315edc1},
  {32'hc4574030, 32'hc22c58ab, 32'h408272ec},
  {32'h43604030, 32'hc2a39ab5, 32'h42778f92},
  {32'hc31454c0, 32'hc2c381cd, 32'h43a89fc5},
  {32'h4479881c, 32'hc3a0cf7e, 32'hc2c48ce4},
  {32'hc48c33d0, 32'hc34156cf, 32'hc269544b},
  {32'h43e9149c, 32'h43922d8c, 32'hc1aec676},
  {32'hc342aef0, 32'hc4006a76, 32'h4363f9bc},
  {32'h4511c51a, 32'h43238012, 32'hc2c9cbc3},
  {32'hc513889b, 32'hc2b5419b, 32'h42c7314c},
  {32'h45034f79, 32'hc3e4f542, 32'h4342e0be},
  {32'hc4c0e6e6, 32'hc4430de1, 32'hc2542789},
  {32'h44f07e2e, 32'hc309d213, 32'hc21b488c},
  {32'hc4d7c8ea, 32'hc2900eab, 32'hc2d10884},
  {32'h445cacd0, 32'hc3743933, 32'hc2d667ee},
  {32'hc3ee7e6e, 32'h4321b544, 32'h428711eb},
  {32'h42b1eb48, 32'hc2f9a5a5, 32'h438e7b5e},
  {32'hc466e4bc, 32'h42cf0a39, 32'h4179c50f},
  {32'h4462706c, 32'hc29668d6, 32'hc35fc19e},
  {32'hc51134cc, 32'hc3acec9b, 32'hc0d7d20d},
  {32'h4469fe30, 32'hc1cf86da, 32'hc33d8ae2},
  {32'hc45a8c28, 32'h435f802a, 32'h43e56345},
  {32'h44de001b, 32'h43f2eddb, 32'hc2b54538},
  {32'hc520a7a9, 32'hc2d7f3b7, 32'h43597130},
  {32'h44af2087, 32'hc0f0a6c6, 32'hc2c56533},
  {32'hc4a61f1c, 32'h429e8146, 32'hc29c4954},
  {32'h44eeb0fa, 32'hc18086ce, 32'h42f13500},
  {32'hc3862270, 32'hc3755e5e, 32'h437bf25a},
  {32'h44724a1a, 32'h435fecb2, 32'hc24afe5b},
  {32'hc5079ac9, 32'h42734cc7, 32'h43886be6},
  {32'h44a53cf8, 32'h417449ac, 32'hc19a5798},
  {32'hc504cfac, 32'hc33c08e7, 32'h43120f53},
  {32'h45053d89, 32'h42c174bd, 32'hc3059552},
  {32'hc3ed6384, 32'hc269a927, 32'h43741b94},
  {32'h451a78a4, 32'h42eb427d, 32'h437eb6b0},
  {32'hc3ce9058, 32'h4384a788, 32'h43fd3dc5},
  {32'h44710862, 32'hc2a7970c, 32'hc2dbef05},
  {32'hc3f93285, 32'h42e934cc, 32'h4404a04b},
  {32'h444f5792, 32'hc2f03c52, 32'hc283aac1},
  {32'hc497d6f1, 32'h437691d6, 32'h42b67b99},
  {32'h44851991, 32'h4329179e, 32'hc394a6a9},
  {32'hc40c5b35, 32'hc2745d2d, 32'h4380fd0c},
  {32'h43baa7e0, 32'h43e04f26, 32'h438f5575},
  {32'hc49eec24, 32'hc2c0d15c, 32'h433b6c98},
  {32'h44bd147d, 32'h435bd01c, 32'hc1d3aae6},
  {32'hc4e32916, 32'h435b2c5b, 32'hc30be313},
  {32'h43f0066c, 32'h431afbde, 32'hc356952d},
  {32'hc43ceb88, 32'hc3b84b2c, 32'hc198f570},
  {32'h42d5a820, 32'hc2c6be91, 32'hc4079699},
  {32'hc4d38c84, 32'h42807a4f, 32'h4387eaab},
  {32'h43f61e7c, 32'hc233a5eb, 32'hc291ae43},
  {32'hc4ff028d, 32'h42c91894, 32'h4393342c},
  {32'h4497bc03, 32'h432fdf6d, 32'h43119242},
  {32'hc28bd63d, 32'h43a22555, 32'h439a63ea},
  {32'h44fcc8bc, 32'hc3b993cc, 32'h41630b5c},
  {32'hc3389404, 32'h4304813d, 32'h430c8ec5},
  {32'h449c38ea, 32'h43799c76, 32'h43743683},
  {32'h43cd5460, 32'hc28c6bfb, 32'hc3e5766a},
  {32'hc463b531, 32'h431e7fe6, 32'h43069d86},
  {32'h43b1f7f0, 32'hc417fa75, 32'hc2dabcb1},
  {32'hc335adb1, 32'h43732b97, 32'h43d796b1},
  {32'h44f08448, 32'hc3716f10, 32'h43e0d9f2},
  {32'hc464aafd, 32'hc101bed4, 32'hc320eb69},
  {32'h41e7f9c0, 32'h432567d5, 32'hc33a9474},
  {32'hc343a2c8, 32'hc34aa4f3, 32'h42cd246d},
  {32'hc2e4a2e0, 32'hc33c04cf, 32'h431a80d9},
  {32'hc4da5950, 32'h431c198b, 32'hc2e86291},
  {32'h44907970, 32'h40888589, 32'h42a70c80},
  {32'hc3f2b06c, 32'hc32af3f1, 32'hc37c0f71},
  {32'h44cc2cde, 32'h438a35da, 32'hc3894dc5},
  {32'hc4acbfd4, 32'hc2b26463, 32'hc39be022},
  {32'h44f77ffc, 32'h43adaa3d, 32'hc344647f},
  {32'hc4d3dacc, 32'hc2a679b2, 32'h43922d91},
  {32'h448b860c, 32'h434fed15, 32'hc2a1efc4},
  {32'hc3d2b0a0, 32'hc28e45b2, 32'h430d07bb},
  {32'h44a57d0a, 32'hc293481a, 32'h41d522ce},
  {32'hc50215b6, 32'h42532fc6, 32'hc27c4e34},
  {32'h44f499d3, 32'hc39ea5fd, 32'h430b2df2},
  {32'hc48c0b8c, 32'hc310d994, 32'hc2a09c94},
  {32'h43c0c02e, 32'hc3955073, 32'hc37f87a5},
  {32'hc4149980, 32'h43a93a00, 32'h42f9f6dc},
  {32'h43ed3ec0, 32'hc03de1f7, 32'hc36aef8f},
  {32'hc49cad8d, 32'hc3833bc6, 32'hc2c843f2},
  {32'h43e0baf8, 32'h4271f6dd, 32'hc374c870},
  {32'hc470feee, 32'hc38ee07d, 32'h42866cfa},
  {32'h4500a64b, 32'hc1ef022d, 32'hc2a17a85},
  {32'hc48aaa45, 32'hc2b5f80a, 32'h43219217},
  {32'h450008cd, 32'h42681580, 32'h42b1d8d9},
  {32'hc3acd22a, 32'h43d85808, 32'hc31a0c48},
  {32'h449bd9d8, 32'h43f61718, 32'h425b077f},
  {32'hc4b8173d, 32'h43f81b3c, 32'hc39ef158},
  {32'h44124628, 32'h431c96a7, 32'hc3ba9d8d},
  {32'hc4210653, 32'h42d738c5, 32'hc320ec62},
  {32'h44b4ebd4, 32'hc35fe050, 32'h41cd9902},
  {32'hc43e6afd, 32'h435d4e29, 32'h4317d748},
  {32'h4430032a, 32'hc2ef9c7c, 32'hc1917c59},
  {32'hc43cb71c, 32'h43315c97, 32'hc3d71679},
  {32'h44900fe7, 32'hc39c8167, 32'hc1532283},
  {32'hc437c958, 32'h43a5a7af, 32'hc34a0fb4},
  {32'h45242730, 32'h428708e9, 32'h42e675d5},
  {32'hc4d25ae5, 32'h419877f8, 32'hc305ce70},
  {32'h44c3e94f, 32'hc3270067, 32'hc2e01bb2},
  {32'hc500fa6a, 32'h4241f96f, 32'h436f9497},
  {32'h4514ea1e, 32'hc1b7d15b, 32'hc2d605a2},
  {32'hc4dda10f, 32'h43abb929, 32'hc3187692},
  {32'h4502f3d2, 32'h43bbbee0, 32'h4152ba79},
  {32'hc3ab8de8, 32'hc2f206e0, 32'h42a2b5f9},
  {32'h4493f84b, 32'h43ebb5db, 32'hc3620c71},
  {32'h42d07de0, 32'hc33ab5c5, 32'h436d8967},
  {32'h44546306, 32'h43eba41b, 32'h43d15a23},
  {32'hc4c5c7d2, 32'h418f4477, 32'hc3596664},
  {32'h447f28d0, 32'hc3c4781e, 32'hc3597f72},
  {32'hc4099a0f, 32'h4352b72c, 32'hc36c7acf},
  {32'h441a53bc, 32'hc2e4661e, 32'h42d6fb2a},
  {32'hc44fb6ca, 32'h41aa2a34, 32'hc27b85a5},
  {32'h44369433, 32'h4352441a, 32'hc33edaa5},
  {32'hc406b404, 32'h423f56c2, 32'hc2f67064},
  {32'h4477eace, 32'hc3b88078, 32'hc410cdd2},
  {32'hc446ec7e, 32'hc2f6ab80, 32'hc36dccdd},
  {32'h44658082, 32'hc3bb036b, 32'h410c7a59},
  {32'hc4fedd7e, 32'hc38a236c, 32'h433fe80a},
  {32'h441be66e, 32'hc31c4009, 32'hc312e9c4},
  {32'hc3aabfed, 32'hc3561a85, 32'h42b6e3a4},
  {32'h4507568a, 32'h42eaa66d, 32'h41cd2698},
  {32'hc4f09b7a, 32'h42cdd764, 32'hc36b4331},
  {32'h44cf2e14, 32'h43bad6e4, 32'hc2f6b7e0},
  {32'hc4c6da3c, 32'hc34b8241, 32'h423de4fb},
  {32'h45055663, 32'hc3824867, 32'h4283caae},
  {32'hc4568401, 32'hc3107563, 32'h42b10872},
  {32'h44fc1cec, 32'hc20220c9, 32'hc1085fd6},
  {32'hc4f181e2, 32'h438bd52e, 32'hc30732c0},
  {32'h43c75104, 32'hc393141d, 32'hc2c29f37},
  {32'hc07a2400, 32'h437b9add, 32'h437eb663},
  {32'h44f7e384, 32'hc37000ee, 32'h42003bd1},
  {32'hc3d05e6d, 32'h43c86466, 32'h41751763},
  {32'h44c5a8af, 32'h4375da34, 32'hc3d6da46},
  {32'hc4b42b4f, 32'h3f52bb08, 32'hc203a695},
  {32'h4498c334, 32'hc3e2e49f, 32'h43a66b12},
  {32'hc45ab0fb, 32'hc379065a, 32'h43bdc588},
  {32'h44fe7448, 32'h432db14e, 32'hc25ee210},
  {32'hc4f0e49e, 32'h41cfffd8, 32'hc25fbb9a},
  {32'h437164c0, 32'h42549447, 32'h42723f0c},
  {32'hc4aeeae2, 32'h42889e1d, 32'h43e194fc},
  {32'h44c38d2b, 32'hc14d483d, 32'h427fea2b},
  {32'hc4c4c388, 32'hc1c4fac1, 32'hc3e78bae},
  {32'h4433947b, 32'hc383d5ca, 32'h436005d4},
  {32'hc50ffd4b, 32'h430013ca, 32'hc3a35647},
  {32'h44dbaba4, 32'h42f4227d, 32'h4378c178},
  {32'h429dcf20, 32'h430a4923, 32'h4140aeb0},
  {32'h447db034, 32'h43c9bf9b, 32'h42f7200e},
  {32'hc3b925f7, 32'hc2be01dd, 32'hc3acd076},
  {32'h45178a8d, 32'h424acb92, 32'hc371a972},
  {32'hc38f0882, 32'hc3826fcc, 32'hc2994673},
  {32'h44629588, 32'hc33ce484, 32'h41c37334},
  {32'h41891000, 32'h42805e4c, 32'hc1c424e1},
  {32'h44f6e646, 32'h434c8ca7, 32'h42f32908},
  {32'hc4b13e57, 32'hc382d0a2, 32'h43148968},
  {32'h44cdcea8, 32'h4293ca20, 32'h43247900},
  {32'hc50ffa3e, 32'h42af060b, 32'hc098fbf0},
  {32'h4511b858, 32'h43726a49, 32'h43efb26b},
  {32'hc48e0686, 32'h42cd337f, 32'hc2d359a3},
  {32'h44d2fde1, 32'h4313e096, 32'hc2bf5448},
  {32'hc40144c8, 32'h42319caf, 32'hc384569e},
  {32'h44b2c402, 32'hc3e2ce05, 32'hc35f59be},
  {32'hc490d768, 32'h434d5623, 32'h42a8383c},
  {32'h43ec1a38, 32'hc3a0d0bf, 32'hc2d88c73},
  {32'h435152e8, 32'h439e7e39, 32'hc3c76f50},
  {32'h4429d157, 32'hc2a4e518, 32'h4331f7d6},
  {32'hc480a66f, 32'h41d65e5e, 32'hc343d958},
  {32'h44adffb0, 32'h4339365b, 32'hc35176cb},
  {32'hc50060e4, 32'hc28eb7be, 32'h43acce4b},
  {32'h43604c20, 32'hc3031700, 32'h4409a070},
  {32'hc4f2e43c, 32'hc0082d41, 32'h42efccc7},
  {32'h420889e0, 32'h43cfaca8, 32'h4210c9c2},
  {32'hc40c0d96, 32'h4343ca8d, 32'hc415f390},
  {32'h43191cee, 32'hc3060b33, 32'hc3eacdb9},
  {32'hc50a57a6, 32'hc304eb94, 32'h438deb92},
  {32'h44cb5113, 32'hc3c24d9f, 32'h42329d87},
  {32'hc4d14154, 32'hc30805cb, 32'h4382c360},
  {32'h44442a5d, 32'h433933ee, 32'h43967f06},
  {32'hc4f257e3, 32'hc2af8ac5, 32'hc30778b4},
  {32'h44e7aad0, 32'hc26f69ce, 32'hc35dbd0c},
  {32'hc450c5c0, 32'h43a7b647, 32'h435d9f46},
  {32'h44f258c6, 32'h429a3645, 32'h42f5f62a},
  {32'hc47d103e, 32'hc305bb60, 32'hc2b5e9c8},
  {32'h4501bb22, 32'hc3c3941d, 32'h43c7aea0},
  {32'hc3fee064, 32'h4153676c, 32'h437db506},
  {32'h4422da48, 32'hc2272f63, 32'hc28d72be},
  {32'hc4a27f71, 32'hc3373a94, 32'h429b3d0d},
  {32'h4452ad5e, 32'h426c0e95, 32'h43408f0d},
  {32'hc50a375e, 32'h42b5e446, 32'hc38d925b},
  {32'h43cdb277, 32'h42dea404, 32'h434df04b},
  {32'hc4a01185, 32'h41852faf, 32'hc35c95c0},
  {32'h4460bd68, 32'h4409f25e, 32'h4350dce9},
  {32'hc481f745, 32'hc21fd44b, 32'h4306bbbd},
  {32'h447a7b24, 32'hc23753ea, 32'hc3743d17},
  {32'hc41f6330, 32'hc391756c, 32'h43a328b4},
  {32'h43de0306, 32'hc343da04, 32'h42fa2ae3},
  {32'hc396b0e4, 32'h432fc697, 32'hc365c041},
  {32'h45079f8a, 32'h422c706b, 32'hc2ab450c},
  {32'hc504e563, 32'h436560ba, 32'hc26acf63},
  {32'h4500fc2f, 32'h432ccc21, 32'h432400b1},
  {32'hc2a347fc, 32'hc2d60cf8, 32'hc3c00b58},
  {32'h44d4ae8f, 32'h43838cbe, 32'h429859ba},
  {32'h434119d8, 32'h42dbe6c2, 32'hc342d6a2},
  {32'h447ae20c, 32'hc3247edd, 32'hc0bd92bc},
  {32'hc465a2cb, 32'hc37a5cf5, 32'hc230f78c},
  {32'h4510c982, 32'h42fce58a, 32'h4336e6ee},
  {32'hc4f4812c, 32'hc318f491, 32'h4243efcb},
  {32'h443c4f84, 32'hc32be1d3, 32'hc2c20fa6},
  {32'h420baf28, 32'hc3addf9a, 32'h42bf4b2d},
  {32'h44ba7a8e, 32'h42605e99, 32'hc34301d4},
  {32'hc4759545, 32'h4384ec1e, 32'h43464139},
  {32'h445e21ac, 32'hc24ca9d9, 32'hc2a46590},
  {32'hc4a62f64, 32'hc283ee84, 32'hc34c16e3},
  {32'h44d8e012, 32'h431fd54b, 32'h42007c58},
  {32'hc4332f60, 32'h431a62ef, 32'h43635261},
  {32'h43f980e0, 32'hc39a8757, 32'hc280f258},
  {32'hc4cf12a0, 32'hc2d4ac19, 32'h42b28332},
  {32'h44ef4c9f, 32'hc29db1e0, 32'h4311670d},
  {32'hc3b5e2e8, 32'hc27d56be, 32'hc318f27a},
  {32'h44c09a88, 32'h4215cc78, 32'hc372d49d},
  {32'h432bed30, 32'hc0a06757, 32'hc394be67},
  {32'h43e5d1d0, 32'hc148287d, 32'hc34f07f6},
  {32'hc487fb48, 32'hc3479345, 32'h4364d83b},
  {32'h443461bc, 32'hc2129353, 32'h42eccc7a},
  {32'hc4d1b6e6, 32'h41582729, 32'h43112e33},
  {32'h43bfb2e4, 32'hc290dbda, 32'hc37824f0},
  {32'hc4c2c886, 32'h4414da25, 32'h438dbfc3},
  {32'h44909926, 32'hc3ba1770, 32'hc3801623},
  {32'hc48e2f44, 32'h428497f8, 32'h41314cec},
  {32'h45031d96, 32'h428f519d, 32'h431afbcd},
  {32'hc3049d23, 32'hc2b67aaa, 32'h437b7b23},
  {32'h43a52fc2, 32'h4208ef85, 32'hc185a776},
  {32'h429337f0, 32'hc3015d80, 32'hc3195ff0},
  {32'h4433f557, 32'hc3982687, 32'hc244a489},
  {32'hc4a913ba, 32'hc34edde6, 32'hc28b5cfd},
  {32'h44896578, 32'h4333e47d, 32'h430df314},
  {32'hc3450550, 32'hc2720770, 32'hc3881205},
  {32'h44e59c17, 32'h4210c2c9, 32'h43a3a418},
  {32'hc47ee489, 32'hc2dd9b8e, 32'h4286ec8a},
  {32'h438a9df0, 32'hc3e5ec52, 32'h42622f23},
  {32'hc4e4038e, 32'h43670dcd, 32'h41a7fb2c},
  {32'h44042b24, 32'h4312cbee, 32'hc30898af},
  {32'hc386da26, 32'h43467e1e, 32'hc35ec982},
  {32'h43fe6942, 32'h429fa8bd, 32'h43d2780f},
  {32'hc4b3c796, 32'h416fca9a, 32'hc3131d39},
  {32'h450aaeb0, 32'h426991df, 32'h432b6b5d},
  {32'hc3c77f64, 32'h4351ebf4, 32'h429e63cc},
  {32'h44c9a813, 32'h42163448, 32'h43304c9d},
  {32'hc4ed3da0, 32'h41d4bec8, 32'hc30c7819},
  {32'h44e72030, 32'h42f2e714, 32'hc24b4605},
  {32'hc50411a4, 32'hc387a3f6, 32'h41521af0},
  {32'h439eda84, 32'h43e6b1a0, 32'h429644ff},
  {32'hc415ff98, 32'hc3b76324, 32'h439a76ee},
  {32'h45075406, 32'hc39d844b, 32'h4303fda4},
  {32'hc4dc8b7e, 32'h434f9186, 32'hc2b82464},
  {32'h44ae2a4a, 32'hc351ef6e, 32'hc2fb9602},
  {32'hc2fb2b86, 32'h42704e13, 32'h43af37c2},
  {32'h447a39e3, 32'hc339a23e, 32'hc26ccc0b},
  {32'hc4f02274, 32'hc2fe26b5, 32'h42ad5c19},
  {32'h44c3bb11, 32'hc40a346b, 32'h4410d9e9},
  {32'hc3628375, 32'hc217dcb1, 32'hc20e7ad0},
  {32'h44384796, 32'hc3a1c02f, 32'hc2928adc},
  {32'hc4f8bb7e, 32'hc27df177, 32'hc3d9dacd},
  {32'h45012956, 32'hc3ef37d9, 32'hc102e4ee},
  {32'hc40a2930, 32'hc2e4d463, 32'hc3357202},
  {32'h44ebf235, 32'hc3c71a72, 32'h418fa5dc},
  {32'hc48afac0, 32'hc30405c6, 32'h437a7e5b},
  {32'h446d90ea, 32'h42dec8c7, 32'h43c9ef3b},
  {32'hc48060be, 32'hc3878646, 32'h438b1d7c},
  {32'h445b2a34, 32'hc25d425c, 32'h4228a1bf},
  {32'hc4a70084, 32'h4328da76, 32'h437b9bf8},
  {32'h44c42dcc, 32'h43b90b7f, 32'h425db5d5},
  {32'hc4b78e87, 32'h432f03be, 32'hc3a914b3},
  {32'h44574859, 32'hc1e88d53, 32'hc1b61c39},
  {32'hc26b9b40, 32'h4336df9a, 32'h43aec10b},
  {32'h44b20b9a, 32'hc31e1d7f, 32'hc3955fd5},
  {32'hc4303edf, 32'h41df7193, 32'h43aa409c},
  {32'h41a41ff8, 32'h43571a72, 32'hc1c0a38b},
  {32'hc3cb0418, 32'h434689e8, 32'h43e44763},
  {32'h44185496, 32'hc3cd5d18, 32'hc3c45ddc},
  {32'hc419d72a, 32'hc2a8871a, 32'h421783a8},
  {32'h44cb9932, 32'h436713af, 32'h41bddef2},
  {32'hc47d24d4, 32'hc23c1965, 32'hc387b17b},
  {32'h44fe45db, 32'h435035ae, 32'h4182e971},
  {32'hc38b5cae, 32'hc232fdbd, 32'hc2f32bc7},
  {32'h44e38ab7, 32'hc1bb9b84, 32'h42849c1a},
  {32'hc4a054c1, 32'h4379c470, 32'hc334e49b},
  {32'h45138af2, 32'hc2e01296, 32'h437b0cfe},
  {32'hc4ba82e4, 32'hc39ca1e2, 32'h4374bd29},
  {32'h444a62d0, 32'h428cd8ee, 32'h431fac86},
  {32'hc4d2cf2c, 32'hc3364d1c, 32'h4268a9bb},
  {32'h44b54f9a, 32'h4391b4f4, 32'hc2c69298},
  {32'hc50f788c, 32'hc2843840, 32'hc379ff9a},
  {32'h44286012, 32'hc384fb34, 32'h43b2cca8},
  {32'hc49d4495, 32'hc2696270, 32'hc3195bee},
  {32'h44e41ed1, 32'hc38c4f41, 32'hc37fdd96},
  {32'hc3e10ba0, 32'hc2b22776, 32'h427dc1cd},
  {32'h44ea7ffa, 32'hc3b6643d, 32'hc3c53095},
  {32'hc50c9020, 32'h4404d7be, 32'h4026a7ac},
  {32'h45014d88, 32'h438a3cbb, 32'hc414b9b7},
  {32'hc4d5cfa7, 32'h43514ad1, 32'h431e48c5},
  {32'h4417249b, 32'h429b2a2a, 32'hc3bdf946},
  {32'hc5031d5b, 32'hc326ad3d, 32'h42b43743},
  {32'h43aa7dac, 32'hc2d590a6, 32'h43499240},
  {32'hc3f28c72, 32'hc3a632cd, 32'h4313cf18},
  {32'h4507f455, 32'h438677dd, 32'hc36ad43f},
  {32'hc4d30054, 32'hc302fd80, 32'h42d8277f},
  {32'h4311652f, 32'hc357a8dc, 32'h429bafc1},
  {32'hc4b20bde, 32'hc064a868, 32'h437993d3},
  {32'h4510d999, 32'hc31d2122, 32'hc349f448},
  {32'hc384f1ce, 32'h432552b8, 32'hc32fcb2c},
  {32'h43e9dc4c, 32'hc33ac06c, 32'h43a6510e},
  {32'h41ff0e00, 32'h437a072d, 32'hc2168084},
  {32'h42fadc40, 32'h44036735, 32'h4315c0bb},
  {32'hc3849a54, 32'hc38a41d4, 32'h4064b908},
  {32'h4454f1fa, 32'hc2c41f00, 32'h429fa495},
  {32'hc458af08, 32'h417d4792, 32'hc265feac},
  {32'h44374a7d, 32'h42e41dbc, 32'hc2afbea8},
  {32'hc4ec88ea, 32'h42470286, 32'h42a07662},
  {32'h42ff9920, 32'hc2ab5cbb, 32'hc3b38d1a},
  {32'hc42abe55, 32'h4333f140, 32'h41f1a86b},
  {32'h4501f1ee, 32'h43d95eae, 32'h42281e6c},
  {32'hc4fe1f41, 32'h437ba698, 32'hc266a6c8},
  {32'h43c92536, 32'hc38daec5, 32'h43406bf5},
  {32'hc42a6948, 32'hc29034be, 32'hc255ac14},
  {32'h444309b0, 32'h43f1c4be, 32'h4359585a},
  {32'hc38bfcc2, 32'h42928795, 32'hc2a31d4d},
  {32'h43de9aa8, 32'h435ef849, 32'hc334372a},
  {32'hc32cdbe6, 32'h43881fe2, 32'h41db1fa5},
  {32'h44138032, 32'hc3e1dbf1, 32'h42de6a10},
  {32'hc4b454a9, 32'hc2fa3e7e, 32'h434d4942},
  {32'h44b43665, 32'hc301deb5, 32'hc3a38a88},
  {32'hc513d0a6, 32'h41b5248c, 32'h42ae6027},
  {32'h4511836c, 32'hc2c6530d, 32'hc2aceafc},
  {32'hc4c86a55, 32'hc35b58b1, 32'h438857f6},
  {32'h44bdea86, 32'hc24917b2, 32'hc32fc5e7},
  {32'hc4b40a1a, 32'h427972a6, 32'h439c71a8},
  {32'h449834e8, 32'hc34e7efa, 32'hc2bebee6},
  {32'hc4f18ebd, 32'h426397a3, 32'h42fbdaa5},
  {32'h44b28314, 32'hc0496ce0, 32'h421f1fe5},
  {32'hc4a835a1, 32'h43999feb, 32'hc3473af0},
  {32'h449dc636, 32'h42a5d4de, 32'h42f6e4fe},
  {32'hc4f97252, 32'hc21e6ebe, 32'h4207a5ae},
  {32'h440f7f56, 32'hc0b08551, 32'h43b3efb3},
  {32'h430b72b8, 32'hc2750fe7, 32'hc3d16072},
  {32'h44fe940f, 32'hc35d287e, 32'h43855944},
  {32'hc4f050fc, 32'h42a00258, 32'hc2b93164},
  {32'h44d62fea, 32'hc1213e74, 32'hc1ebc6f9},
  {32'hc396a420, 32'hc299fc44, 32'h425f6834},
  {32'h449bf8b6, 32'hc3808ef8, 32'hc3a24a3c},
  {32'hc458a78c, 32'h42f9ec5c, 32'h42e7225e},
  {32'h44b43db9, 32'h4066d111, 32'h42d8e274},
  {32'hc4f6dcab, 32'h43c1f956, 32'h43954f1f},
  {32'h4510e6fb, 32'h437031a8, 32'hc282414f},
  {32'hc510e5e1, 32'hc2700553, 32'h43957e33},
  {32'h44c467ab, 32'h43aaef86, 32'hc2faa832},
  {32'hc507f947, 32'hc3a714df, 32'hc1a1389c},
  {32'h450ebd3d, 32'h41cb9f22, 32'h42862c26},
  {32'hc4925f10, 32'h43649db1, 32'h438f64ed},
  {32'h446a8aee, 32'hc2007e18, 32'hc357bf61},
  {32'hc4ebfe72, 32'h43e21b71, 32'h43cd0f09},
  {32'h45034161, 32'h4367ecaa, 32'hc38330fa},
  {32'hc4a247be, 32'h4310a2ca, 32'hc360df1c},
  {32'h444ace86, 32'h43f6f60d, 32'h41270de8},
  {32'hc5202547, 32'h4337ec0f, 32'h43f3d103},
  {32'h42854d3e, 32'h42cbebde, 32'hc17ffaf1},
  {32'hc3ce3ad5, 32'h3feffb4a, 32'hc35e5b52},
  {32'h4287c850, 32'hc33dc821, 32'h433e1a03},
  {32'hc518617d, 32'hc2d89ed3, 32'h42236e06},
  {32'h44f301a1, 32'hc361e014, 32'h42fe9ba2},
  {32'hc508b4a5, 32'h43e3c12d, 32'hc312c0b2},
  {32'h43097694, 32'hc31dc298, 32'hc3c2369f},
  {32'hc4b80815, 32'h425d73e8, 32'h43e45217},
  {32'h44c87910, 32'h433a49e3, 32'hc2b1a7a4},
  {32'hc2c6c84c, 32'h42ca74b6, 32'hc127eff1},
  {32'h4432b15e, 32'hc2ac8748, 32'hc2a19d8f},
  {32'hc3b92240, 32'h42a1ddd4, 32'hc21d5b27},
  {32'h438f5b80, 32'h420a0ef7, 32'hc2842bfc},
  {32'hc5034abc, 32'h438b55bd, 32'hc0e0a0eb},
  {32'h44e08348, 32'h4354615e, 32'h42cfa58f},
  {32'hc48db090, 32'hc2a004be, 32'h43976c75},
  {32'h43ba19b4, 32'hc3d32b8e, 32'h4336e722},
  {32'hc4d05ae6, 32'hc355d8ec, 32'h42210d8d},
  {32'h440ec576, 32'hc3beeca1, 32'hc36e19f3},
  {32'hc302f8a0, 32'h4388ae86, 32'hc335a42d},
  {32'h445fea74, 32'hc31210a4, 32'hc2f05433},
  {32'hc50f0fc6, 32'hc2338668, 32'h43a4e8d2},
  {32'h44a02941, 32'h43593847, 32'hc39b0212},
  {32'hc493591f, 32'h40641b38, 32'hc3141743},
  {32'h44222c7b, 32'hc215bf96, 32'hc11c34bd},
  {32'hc4e62fcb, 32'hc3be1a4d, 32'h4306439a},
  {32'h43ad5468, 32'h434ca59d, 32'hc1f1560d},
  {32'hc3c2ae34, 32'h43116c5c, 32'h43a357da},
  {32'h43e6b384, 32'h42211868, 32'hc34814e0},
  {32'hc49de526, 32'hc32339c0, 32'hc3924dac},
  {32'h42a0369c, 32'hc0038b14, 32'h436f9b00},
  {32'hc4ed456d, 32'hc2b0060e, 32'hc33c3117},
  {32'h44de9efc, 32'hc1d68526, 32'h43b7335b},
  {32'hc507ed79, 32'hc346785c, 32'hc2a33441},
  {32'h44a340fa, 32'h42437252, 32'hc3e87927},
  {32'hc3f3c67e, 32'h4296ae37, 32'hc20c2a02},
  {32'h4510b2d0, 32'hc37714ba, 32'hc1ff3342},
  {32'hc445fd12, 32'h43cee5ba, 32'h432c6564},
  {32'h44993e5a, 32'h43c22fb9, 32'hc3c0b8e7},
  {32'hc500c4a4, 32'hc3741023, 32'h43ff840c},
  {32'h44be3b8b, 32'h4257e100, 32'h430a4328},
  {32'hc4c0ed70, 32'hc2c2a99f, 32'hc2627e71},
  {32'h4429f4b6, 32'h437724f4, 32'h4393d597},
  {32'hc415c29a, 32'hc12bdb29, 32'hc3a448e0},
  {32'h451c23da, 32'hc4002d64, 32'h4308f02d},
  {32'hc4083058, 32'h43172125, 32'h4379be82},
  {32'h44aba934, 32'hc34f901b, 32'hc326bda1},
  {32'hc3ee3837, 32'hc309f596, 32'h40a6c300},
  {32'h44be7c0a, 32'h42cdcf8c, 32'hc2c280a3},
  {32'h438889f0, 32'h4361a618, 32'h43b5be36},
  {32'h450d28ad, 32'hc3cfaed9, 32'h42f29edb},
  {32'hc51bfe08, 32'hc2f6ef28, 32'h43130d94},
  {32'h439d5398, 32'hc3b62994, 32'hc30debbb},
  {32'hc4f52082, 32'hc2344b92, 32'h43a14bfd},
  {32'h4480cad6, 32'h41a58735, 32'hc3d3753a},
  {32'hc4a0ee2b, 32'h43437976, 32'h435609d0},
  {32'h4481cff2, 32'hc399966b, 32'h41b4002b},
  {32'hc46960d7, 32'h43850a31, 32'h4335095c},
  {32'h4412c68a, 32'h430c395f, 32'h43fae274},
  {32'hc40e8410, 32'h421b7754, 32'hc266274f},
  {32'h4524ad3c, 32'h43d05cbc, 32'hc2a85d32},
  {32'hc4f4f2bf, 32'h40ffcba0, 32'hc3503a30},
  {32'h445b08aa, 32'hc2a386b9, 32'h439a13ea},
  {32'hc50a4397, 32'h43058008, 32'h422b0749},
  {32'h432bbeb1, 32'h43d9ee59, 32'h42e7e3c4},
  {32'hc4f61532, 32'h43c5f026, 32'h4372e47b},
  {32'h4244a128, 32'hc30aaa17, 32'hc175df48},
  {32'hc40a96f1, 32'hc3024b8b, 32'hc3857671},
  {32'h44a7608d, 32'h429022c0, 32'h43d15ed0},
  {32'hc51ffed6, 32'hc2bec99c, 32'hc30b12e7},
  {32'h45136ce9, 32'h42c06916, 32'h42cefe3c},
  {32'hc4f4a5cd, 32'h42a35360, 32'h4382552d},
  {32'h449971c3, 32'hc38264b5, 32'h42ec3673},
  {32'hc2f77ba6, 32'hc37cda98, 32'h421f3c70},
  {32'h43bb8fac, 32'h43556276, 32'h42cb5a25},
  {32'hc49b1469, 32'hc276dd22, 32'hc3be2f50},
  {32'h44c2dc20, 32'hc31bdac0, 32'h43b2a0e4},
  {32'hc4bfdb27, 32'h42a1bd8a, 32'hc30947d1},
  {32'h45133bf9, 32'hc314c078, 32'h433a93e7},
  {32'hc4374f32, 32'h42b0ed87, 32'hc2155974},
  {32'h447985c5, 32'hc23ab112, 32'h43071edc},
  {32'hc4e188b0, 32'h41d285e2, 32'hc2b23b26},
  {32'h4484d7f8, 32'hc29b4660, 32'hc212bde7},
  {32'hc464ce86, 32'hc3b9f00b, 32'hc25f81cf},
  {32'h44af8047, 32'hc350b892, 32'hc30b4455},
  {32'hc504a67d, 32'hc28ec426, 32'hc320bcfd},
  {32'h4478919d, 32'h418a38a9, 32'hc35e87d7},
  {32'hc4d81f7c, 32'hc23d3ae8, 32'h429e327d},
  {32'h442c5f49, 32'hc36f0202, 32'hc305a0dd},
  {32'hc450f2af, 32'hc2dbbb93, 32'h438f69d5},
  {32'h44956b33, 32'h42a8193a, 32'h435c10dc},
  {32'hc41c1c7c, 32'h439a6c72, 32'hc3afb92d},
  {32'h44d86ad3, 32'hc34e5d27, 32'hc2c054a8},
  {32'hc2d964d2, 32'hc1b5d9bc, 32'h428b8ba0},
  {32'h4493a91e, 32'hc2f517cf, 32'h438ac437},
  {32'hc4b2ca9d, 32'h42f90efc, 32'hc39f40f0},
  {32'h4525ff8d, 32'h4290b377, 32'h43312fa7},
  {32'hc50cca4e, 32'hc316f0c4, 32'hc2a1bc39},
  {32'h441957ca, 32'h434cf6c8, 32'h43a57468},
  {32'hc50004a1, 32'h434211d8, 32'h42f20804},
  {32'h451526da, 32'hc326407d, 32'h430371f3},
  {32'hc4f60641, 32'hc30f5703, 32'hc27d7bbe},
  {32'hc2f981c2, 32'h431616c0, 32'hc2cfc778},
  {32'hc4a04148, 32'h43420373, 32'h43730323},
  {32'h448269fa, 32'hc1e2adb9, 32'h430c5c9a},
  {32'hc2289ffc, 32'hc2734a44, 32'h431fea55},
  {32'h4503a136, 32'h4221ae8c, 32'h415ef5f8},
  {32'hc4fb84b3, 32'h431ef137, 32'h42201d56},
  {32'h444899a5, 32'h404d4a00, 32'h436330d5},
  {32'hc49870b0, 32'h433b6f03, 32'hc3876499},
  {32'h44edbfa0, 32'h423ec109, 32'h43067889},
  {32'hc4a0e9ff, 32'h434d71d6, 32'hc31442a9},
  {32'h43ec1885, 32'hc335b0df, 32'hc03d7738},
  {32'hc47d6722, 32'hc249a7c8, 32'hc3a292ca},
  {32'h447a5c1b, 32'hc3100ffe, 32'h4328af91},
  {32'hc493386a, 32'h439f648a, 32'hc3aff7a3},
  {32'h4471b2f2, 32'h430e235e, 32'h4026e344},
  {32'hc4dad6d8, 32'hc24e8739, 32'hc28020dc},
  {32'h444aea3a, 32'hc39b7d9d, 32'h4342be56},
  {32'hc50cd535, 32'h430cb994, 32'hc2ae7f82},
  {32'h451a67b3, 32'h41b7d379, 32'h43aa3b26},
  {32'hc4e5cb9b, 32'hc26f9212, 32'h43be10d4},
  {32'hc3b8b00a, 32'h428ec0ac, 32'hc39df348},
  {32'h44071fd2, 32'hc3af25ed, 32'h438338a2},
  {32'hc3e2f082, 32'h440a2e2d, 32'h41db8af6},
  {32'h44673584, 32'hc20c8fb2, 32'h4378ff08},
  {32'hc414b600, 32'h4362b530, 32'hc3d8813f},
  {32'h44958917, 32'hc263806a, 32'h431d0b64},
  {32'hc4af9c2e, 32'hc2a9b029, 32'hc37fc3b9},
  {32'h448068e8, 32'h439102a4, 32'hc34f6e5e},
  {32'hc3b780d9, 32'hc36261eb, 32'hc321d2ef},
  {32'h432a7659, 32'hc3257828, 32'h420d07f0},
  {32'hc439ceb4, 32'hc39d5de3, 32'hc3e3589d},
  {32'h44596a16, 32'h4264acd2, 32'h4342c58f},
  {32'hc414a683, 32'hc3d12357, 32'hc35c9420},
  {32'h404b3800, 32'h43620b04, 32'h436916d1},
  {32'hc4f90803, 32'hc3801faf, 32'h437f9659},
  {32'h431f6f2c, 32'hc348970e, 32'hc3d37dd0},
  {32'hc4e0e2e2, 32'h4395ca22, 32'hc385be1b},
  {32'h43b945e8, 32'hc3457f23, 32'hc0e025fc},
  {32'hc41b6a3d, 32'h43d1fd44, 32'hc3466c28},
  {32'h43f26be0, 32'hc2d180bc, 32'hc3100c18},
  {32'hc48a0b79, 32'h43967892, 32'hc384b1d0},
  {32'h44edc084, 32'h4212f816, 32'h43c5f8b5},
  {32'hc446d71b, 32'hc3c44591, 32'hc254bf5a},
  {32'h442a59f6, 32'h436dd480, 32'hc32e7046},
  {32'hc5052115, 32'h43195bd7, 32'h42aa84e7},
  {32'h4399adb0, 32'hbd6bf89c, 32'h42b86984},
  {32'h43cf9160, 32'hc36e4204, 32'hc2a025f8},
  {32'h44922305, 32'h4307b157, 32'h42351ffd},
  {32'h4290446c, 32'h42addb35, 32'hc385446f},
  {32'h44aa524e, 32'hc3082ee0, 32'h41726065},
  {32'hc3f2189c, 32'h438e7f0a, 32'hc37c6cd8},
  {32'h44a33cc3, 32'hc3c975ce, 32'h4393a343},
  {32'hc4a7d56f, 32'hc29cba43, 32'hc2980ced},
  {32'h44a1c150, 32'hc302411d, 32'h4262d819},
  {32'hc4857f6c, 32'hc38c3558, 32'hc39b9ff8},
  {32'h44b38910, 32'hc28b0e4d, 32'h42e4a954},
  {32'hc487f247, 32'h42e31ba9, 32'hc3242eb3},
  {32'h43c2fddc, 32'hc326474e, 32'h43d1cf71},
  {32'hc468fe84, 32'h42ced3bb, 32'hc3937547},
  {32'h4504c329, 32'h439615f8, 32'h431f347e},
  {32'hc513dc22, 32'hc3903535, 32'h41d1d6cd},
  {32'h449f2ecd, 32'h42cb0654, 32'h44117bac},
  {32'hc4393788, 32'hc3b62572, 32'hc321eb36},
  {32'h44027475, 32'h4266d0d2, 32'hc303a11e},
  {32'hc306ee00, 32'hc2e3a200, 32'hc333b8bb},
  {32'h450d7030, 32'hc319891a, 32'h439ccdc5},
  {32'hc339a378, 32'h43937e42, 32'hc2096698},
  {32'h451b36df, 32'h435670cd, 32'hc37c8871},
  {32'hc4d97b7d, 32'h43630330, 32'hc334fe9e},
  {32'h43a6eeaf, 32'hc35d45f6, 32'hc34a2462},
  {32'hc464c4f0, 32'hc3a9f833, 32'h43216f48},
  {32'h44e1dd3e, 32'hc34788ab, 32'hc2ad474c},
  {32'hc29be8d8, 32'hc3129bf3, 32'h42a18b75},
  {32'hbfd83400, 32'h439c0f8d, 32'hc33a58e1},
  {32'hc50d66da, 32'hc2b5124e, 32'hc3a7c883},
  {32'h444efbdd, 32'hc3178146, 32'hc32f2591},
  {32'hc508a0a5, 32'h437f0364, 32'h42b2703b},
  {32'h44d4f9aa, 32'h4339a744, 32'hc3b52305},
  {32'hc4ba2a7e, 32'hc3abbdfb, 32'h4114d0ff},
  {32'h40c50d00, 32'h42615140, 32'hc1ec8610},
  {32'hc4ee62f2, 32'hc2c7516e, 32'h415e868c},
  {32'h43b5ed62, 32'hc3580905, 32'hc2e8c6bb},
  {32'hc4f448c7, 32'hc2c7adf3, 32'hc3fb6604},
  {32'h44dd252f, 32'h43a9911f, 32'h43b3af4d},
  {32'hc5067713, 32'h41c3b461, 32'h43ef2384},
  {32'hc25bfc48, 32'h43b3c7d0, 32'h4410f4b9},
  {32'hc4acc5f7, 32'hc2898244, 32'h41aed4f5},
  {32'h438ee1ea, 32'hc2d3fc52, 32'hc0157435},
  {32'hc4ce48a4, 32'hc338c8e2, 32'hc3c4f4fa},
  {32'h4501c2b4, 32'hc2ae0fdc, 32'hc23c73a5},
  {32'hc1a0e85a, 32'h42dadd2a, 32'hc320fa45},
  {32'h43ad102c, 32'hc38f6488, 32'h4382852f},
  {32'hc2847760, 32'h43735df3, 32'h443e447c},
  {32'h44f7944e, 32'hc3a90302, 32'hc2ccdcd9},
  {32'hc4801268, 32'h42d1f177, 32'hc3acf47d},
  {32'h449a98e2, 32'h42c3930c, 32'hc38d9741},
  {32'hc44c262a, 32'hc3064b96, 32'hc0f45111},
  {32'h44f02269, 32'h43823018, 32'h42e23fce},
  {32'h4131f200, 32'h43aa1797, 32'h42eba4c2},
  {32'hc3840d23, 32'hc31e3456, 32'h439bab48},
  {32'hc2cffbf0, 32'h423339af, 32'hc2c0036d},
  {32'h44237250, 32'h439c9d8b, 32'h42521d52},
  {32'hc4eaadac, 32'hc39ca4c6, 32'hc381d484},
  {32'h447b755e, 32'hc2b59409, 32'hc3573cf7},
  {32'hc4dd5da9, 32'h438aaf3b, 32'h431eb225},
  {32'h45104141, 32'h43912303, 32'hc08d5a1e},
  {32'hc4bf922a, 32'h4313e6d9, 32'h436eefd8},
  {32'h44fdef0c, 32'h42a531b7, 32'hc2acd04a},
  {32'hc3f51121, 32'h42ba5419, 32'h42f1c022},
  {32'h44c5fe3a, 32'hc326d12b, 32'h42c9b4ab},
  {32'hc505df6b, 32'h4356f7fe, 32'hc36634cd},
  {32'h44d31c56, 32'h428504c0, 32'hc31a34ea},
  {32'h43158479, 32'h438d2572, 32'hc36890ad},
  {32'h450345a1, 32'h42d9d117, 32'h433e299a},
  {32'hc4de75e6, 32'hc3a6a2cf, 32'hc24ab71a},
  {32'h43419320, 32'h42339b72, 32'hc3e6046a},
  {32'hc4a4e6b0, 32'hc2e23f53, 32'hc109561a},
  {32'h41ac9170, 32'hc2eb6773, 32'hc3011bfc},
  {32'hc4868240, 32'hc20e8b65, 32'h433a46f8},
  {32'h449adb06, 32'h43d5cd11, 32'hc3545aac},
  {32'hc4abde68, 32'hc37b5289, 32'h430a4b74},
  {32'h44ae1bc8, 32'h3eadada1, 32'hc2da5516},
  {32'hc45c2162, 32'h433d35bc, 32'hc28aaf66},
  {32'h4371bad0, 32'hc31fa2e0, 32'h42baea47},
  {32'hc4855cdf, 32'h439f0abf, 32'h43310717},
  {32'h44b3a776, 32'hc38759e6, 32'hc1ea4ed0},
  {32'hc509c494, 32'h42b81dda, 32'h43442e73},
  {32'h43a1b710, 32'h43782d62, 32'hc349c18d},
  {32'hc4175634, 32'h42b27cf4, 32'h43a66ac4},
  {32'h44411260, 32'hc3360964, 32'hc18da952},
  {32'hc3417fb0, 32'hc180afa0, 32'h431a95a3},
  {32'h445e5de4, 32'hc2bbd2fb, 32'hc34168dd},
  {32'hc494fd16, 32'hc3d6c9cc, 32'h4249fc34},
  {32'h44fe4447, 32'h434f2447, 32'h438261c5},
  {32'h430e66f0, 32'hc2a4be1a, 32'h429914a6},
  {32'h44c24742, 32'hc2355fcb, 32'hc3c7f7cc},
  {32'hc3601390, 32'hc31a38fe, 32'hc2e5b1c7},
  {32'hc31f0db8, 32'h423fc356, 32'h439e9d9d},
  {32'hc4fca0f5, 32'h42084efe, 32'h439127df},
  {32'h444ef781, 32'h43d0c5c4, 32'hc22992f1},
  {32'hc463ecf6, 32'h42918b35, 32'h43526029},
  {32'h449db49c, 32'hc3780e63, 32'h42939fe6},
  {32'hc481cb23, 32'hc2afea69, 32'h43a6c6e2},
  {32'h4436a0e3, 32'hc2f05186, 32'h4369789c},
  {32'hc42f5fda, 32'hc24fcbd7, 32'hc1597446},
  {32'h450109c5, 32'hc131cbe7, 32'hc1e2d737},
  {32'hc3fc6fe4, 32'hc346e263, 32'hc39d5392},
  {32'h44bfda28, 32'hc330e53c, 32'h42f365d2},
  {32'hc44f8c14, 32'h42833ed6, 32'h428cec40},
  {32'h44efb5f2, 32'h435ffeaf, 32'hc3bb8dff},
  {32'hc20ae328, 32'hc3b05b4f, 32'hc399578e},
  {32'h4416c321, 32'hc3109eb2, 32'hc31cef33},
  {32'hc491f5fa, 32'hc3538e24, 32'hc19dfd1d},
  {32'h442e05b7, 32'hc0875b37, 32'hc1a61e86},
  {32'hc44e39d3, 32'h42b5ef0e, 32'h42c6d658},
  {32'h448f2779, 32'hc2837627, 32'hc3bfe296},
  {32'hc5013556, 32'h425fedb1, 32'h41a9d82f},
  {32'h4502041c, 32'h419c69a2, 32'hc40116ef},
  {32'hc4b0d5ae, 32'h4325d474, 32'h433f8e8d},
  {32'h44ed7c10, 32'h428d43e8, 32'h440d27ab},
  {32'hc417d660, 32'h42be8236, 32'hc31b8e56},
  {32'h447607b6, 32'hc27100c8, 32'h40920646},
  {32'hc4eda27d, 32'h401e6d70, 32'h4350ba50},
  {32'h44f11377, 32'h430f50a5, 32'hc249ce57},
  {32'hc403b378, 32'h40948e6b, 32'h421f0090},
  {32'h441a8f1e, 32'h42e2108c, 32'hc328e25b},
  {32'hc2915c00, 32'hc307566d, 32'h44190c9f},
  {32'h44980186, 32'h432a1b12, 32'h43a6082d},
  {32'hc4a3208b, 32'hc39ba7c5, 32'h4385acd8},
  {32'h45193af3, 32'h43622acd, 32'hc2b27374},
  {32'hc4d7268e, 32'h43103f53, 32'hc2936abb},
  {32'h44da4700, 32'h43f9929d, 32'h43ed963c},
  {32'hc3bafb43, 32'hc2f6389c, 32'hc3aac202},
  {32'h44a1c920, 32'hc2cce567, 32'h41995e59},
  {32'hc4d7bb60, 32'h42bc8fa8, 32'h417357e4},
  {32'h44168964, 32'h4276284c, 32'hc32e6153},
  {32'hc508ebb5, 32'h42670904, 32'hc385b1cb},
  {32'h449b1a46, 32'hc32d898f, 32'h43acaf9e},
  {32'hc4c40838, 32'h43c9e309, 32'hc368c9b0},
  {32'hc38aa721, 32'hc2042828, 32'h43e8a8b2},
  {32'hc38e3318, 32'hc084c230, 32'hc34052d6},
  {32'h44e47c2a, 32'h42ff3236, 32'hc38310a8},
  {32'hc3c6e8ac, 32'hc326a4ed, 32'h42f3940c},
  {32'h44288bd3, 32'h43846447, 32'hc3317fa2},
  {32'hc4dc8d19, 32'hc0e33f80, 32'hc2cf913b},
  {32'h44ed72e4, 32'h41a1e2ac, 32'hc30b6555},
  {32'hc2e3f6dc, 32'hc36880a1, 32'h432005b8},
  {32'h43261b56, 32'h43303414, 32'h42db5991},
  {32'hc43cc9d3, 32'hc2aeafd0, 32'hc20ae6ae},
  {32'h443a32b7, 32'hc3d50212, 32'hc067503c},
  {32'h42e463d9, 32'hc16978a9, 32'hc2d3e08c},
  {32'h44902d8e, 32'hc3bc63dd, 32'hc2d1f39f},
  {32'hc4b8caf1, 32'hc414fe0c, 32'h4179f8b8},
  {32'h4479e3b4, 32'h430c9efd, 32'hc3207e63},
  {32'hc506528a, 32'hc29fd71d, 32'hc3224b99},
  {32'h44bd6d2a, 32'h43e71e4b, 32'h44027b02},
  {32'hc5058567, 32'h420fa68a, 32'h4339090e},
  {32'h43d63738, 32'hc2c6091a, 32'h42b5b462},
  {32'hc48b66ca, 32'h43b9785a, 32'hc2cc2902},
  {32'h44d1bb6c, 32'hc2f4dec4, 32'hc3607ae7},
  {32'hc5113e57, 32'h421c85f3, 32'hc2e52030},
  {32'h447fc0a0, 32'hc30a5a06, 32'h429aad14},
  {32'hc4025d2c, 32'hc2220288, 32'hc3c827b9},
  {32'h448826cf, 32'h4081c086, 32'h3fc268c2},
  {32'hc4109d02, 32'hc39a1830, 32'hc32a05b7},
  {32'hc23b4ed0, 32'h4324fb9b, 32'hc31b9bcd},
  {32'hc4c313e3, 32'h4304779d, 32'h434580ad},
  {32'h451678e7, 32'h3f641818, 32'hc38f80d3},
  {32'hc3ef0bc4, 32'h42951d39, 32'hc20a0df1},
  {32'h428223f2, 32'hc2fc2f6d, 32'h425c704c},
  {32'hc5022cdb, 32'h43e512ab, 32'h42c47a8c},
  {32'h444ce198, 32'h40b5c692, 32'h43eee326},
  {32'hc4320b38, 32'hc3be40f0, 32'hc2d0cf88},
  {32'h45147adf, 32'h41a19091, 32'h42d3b322},
  {32'hc49f99f4, 32'h43405c14, 32'h436a029b},
  {32'h44f4c2dc, 32'hc24f9feb, 32'h439aead5},
  {32'hc4b1c906, 32'h43dde040, 32'hc2926b86},
  {32'h44b09797, 32'hc304f5eb, 32'h43878bb9},
  {32'hc3c5bd59, 32'hc3cd05ac, 32'h431b3be2},
  {32'h44e3184d, 32'h43b8d84c, 32'h4284dbdc},
  {32'hc4e7a70e, 32'hc400b10c, 32'h431ee6e6},
  {32'h440c4644, 32'h42732aa0, 32'hc3716193},
  {32'hc49db8f4, 32'hc3469a9a, 32'h41f44bf4},
  {32'h450b62f1, 32'h42c73ecc, 32'hc3d4085c},
  {32'hc49d9373, 32'h43c62ff0, 32'h43ed9a1d},
  {32'h44833b5a, 32'hc38923d4, 32'h438e12ef},
  {32'hc44d2916, 32'hc3955a78, 32'h432cc5f4},
  {32'h44b31259, 32'hc38653f3, 32'hc247ce0a},
  {32'hc510a787, 32'h432baacc, 32'hc2803441},
  {32'h448106c7, 32'hc239c513, 32'hc2719711},
  {32'hc4a65172, 32'h4337b5b8, 32'h432496bf},
  {32'h44bf943c, 32'hc38db02d, 32'hc4064fcc},
  {32'hc3462c8c, 32'hc12a4d16, 32'hc34749ca},
  {32'h45016b42, 32'hc35d7f58, 32'h43a9e9e4},
  {32'hc3b905c4, 32'h43a4a853, 32'h43d0da5e},
  {32'h44aeb577, 32'hc3d12bab, 32'hc28b7615},
  {32'hc4aa8155, 32'hc34d37fd, 32'hc1b4cb07},
  {32'h436d2e76, 32'h44029223, 32'h441e0555},
  {32'hc5004f2b, 32'hc38995d3, 32'hc337b373},
  {32'h43b53534, 32'h435106de, 32'hc24c82b3},
  {32'hc4a18c2c, 32'hc3d7f332, 32'hc331f2d6},
  {32'h44cbd06e, 32'h437f0140, 32'hc2adc45a},
  {32'hc4f83627, 32'hc31f66a6, 32'hc1af7d56},
  {32'h44bd5ea2, 32'h424ebe32, 32'hc2fff06d},
  {32'h42cc8833, 32'hc2d4958b, 32'hc36631bc},
  {32'h4516f2cf, 32'h42eb2c42, 32'hc33c4e32},
  {32'hc489935a, 32'hc367a87d, 32'hc260c97c},
  {32'h45088381, 32'hc3af0de6, 32'hc2d98203},
  {32'hc406dec5, 32'hc30aa604, 32'h42c12a11},
  {32'h4291ea80, 32'hc3af7a49, 32'h421f5e6f},
  {32'hc4df7610, 32'h41bb56f1, 32'h42d45b82},
  {32'h4383d1b8, 32'h434ae77b, 32'hc3195672},
  {32'hc4e012b6, 32'hc3427c1d, 32'hc3a91554},
  {32'h4498c2a5, 32'hc25116d6, 32'hc364d980},
  {32'hc494b76f, 32'hc2cb56f2, 32'hc24c54da},
  {32'h448c1993, 32'hc339f3c6, 32'hc39a53e9},
  {32'hc3b024d8, 32'hc20f494d, 32'h4383736d},
  {32'h44cb4142, 32'h42aca4eb, 32'hc3baf627},
  {32'hc4f2115c, 32'h41a11b2f, 32'h43a22866},
  {32'h44919eab, 32'h4280e3ca, 32'h434216c1},
  {32'hc4125efe, 32'hc33920e0, 32'hc391fbad},
  {32'h440fcf60, 32'hc2e42b99, 32'h42a6e643},
  {32'hc4b63f6b, 32'h43331eaa, 32'hc38639a4},
  {32'h43c8b85c, 32'h426c2302, 32'h4328d2f7},
  {32'hc50c5f60, 32'h43a9957e, 32'h437b3081},
  {32'h451d7a3c, 32'hc44b3a65, 32'h42747f23},
  {32'h4290afc2, 32'h4335076b, 32'hc37923c1},
  {32'h44e14a11, 32'hc36ed6c9, 32'hc24d82bc},
  {32'hc490e1c7, 32'h4371594f, 32'h43acd7ed},
  {32'h44f42451, 32'hc21064de, 32'h410a000a},
  {32'hc42c1e2e, 32'h435c30fe, 32'hc313b26f},
  {32'h444b7692, 32'hc2f38066, 32'h43a53032},
  {32'hc41e6b2c, 32'hc30638fb, 32'hc3570bbb},
  {32'h44cfd755, 32'h433cf21a, 32'h430c63b6},
  {32'hc4943ed5, 32'h41e1f83a, 32'h42e04642},
  {32'h43a68f46, 32'hc3814d02, 32'hc2320694},
  {32'hc4a0686e, 32'hc36f0f5b, 32'hc333d698},
  {32'h440bedd8, 32'h439557d7, 32'h43bb4495},
  {32'hc3f01303, 32'hc3586952, 32'h438a4054},
  {32'h450270c2, 32'h43cd41bb, 32'hc11c47b5},
  {32'hc45b4346, 32'h42be7bf6, 32'hc29226dd},
  {32'h451c5249, 32'hc40ce01f, 32'h4330dcc4},
  {32'hc5052573, 32'h4362b6e3, 32'hc110aa37},
  {32'h44ecb4f3, 32'h43adb948, 32'h42c266c6},
  {32'hc47976e4, 32'hc38e09fc, 32'hc34e27ed},
  {32'h4452df34, 32'h438f7cbb, 32'h434f6016},
  {32'hc4fa7316, 32'h42a6cd47, 32'h41900b08},
  {32'h44d057ba, 32'hc392d4d6, 32'h43ccd03c},
  {32'hc45dc3db, 32'hc3a3014a, 32'hc36dcff1},
  {32'h441f5f5a, 32'hc27182fe, 32'h42a70286},
  {32'hc468d29c, 32'h432ff09c, 32'h43156d50},
  {32'hc20916e0, 32'hc35cc764, 32'h42f54cac},
  {32'hc501120f, 32'hc001533e, 32'hc12304d4},
  {32'h44e2d076, 32'hc2813eb5, 32'h42cda6e3},
  {32'hc40d8a48, 32'h42d43669, 32'hc30c47d1},
  {32'h44c4a7fc, 32'h4363677a, 32'hc37b6cc3},
  {32'hc4fee4d2, 32'h433e6c57, 32'hc329de77},
  {32'h44a593b0, 32'h434a39d2, 32'h43376c57},
  {32'hc48d11a9, 32'hc2643610, 32'hc3b5d6aa},
  {32'h450d8da8, 32'hc3792f1b, 32'h41960ba2},
  {32'hc5014328, 32'h433a74a5, 32'h43fe28fe},
  {32'hc2440ad0, 32'h422f33b4, 32'h418b2242},
  {32'hc4ffb134, 32'h42a141ac, 32'hc1b970d3},
  {32'h44866e3a, 32'hc32587f0, 32'h438d60de},
  {32'hc49d8354, 32'h42cf058a, 32'h4382b182},
  {32'h444d7300, 32'h433415c6, 32'h430ef43c},
  {32'hc4353d51, 32'hc2e1b960, 32'h42a92ccb},
  {32'h44314984, 32'hc398cd3a, 32'hc2c0bb5a},
  {32'hc4c1c534, 32'hc1bfc1d2, 32'h42d707d4},
  {32'h44fd4cf6, 32'h4372c67a, 32'h43c204e0},
  {32'hc4a6b900, 32'hc32752f2, 32'hc1a253c9},
  {32'h41dfcfa0, 32'h4382717a, 32'hc3038fc5},
  {32'hc4506066, 32'hc3d70820, 32'h43432edd},
  {32'h4507608e, 32'hc3428fba, 32'hc30cb2f3},
  {32'hc409dc6a, 32'hc384910c, 32'hc3687057},
  {32'h44a5c536, 32'h42aafefb, 32'hc3aa6b80},
  {32'hc2328800, 32'hc2b47f65, 32'h404e2054},
  {32'h4367a340, 32'h4343ff28, 32'h42bca486},
  {32'hc390a1b0, 32'hc2784964, 32'hc33c7bad},
  {32'h4487a1aa, 32'hc283bdbf, 32'hc26c461c},
  {32'h42b26130, 32'hc39aa94f, 32'h42887762},
  {32'h4444dd50, 32'hc0e924a0, 32'hc32cc690},
  {32'hc49e0bfc, 32'h433f2cbc, 32'h4401052b},
  {32'h446ac01c, 32'hc28f2e06, 32'hc37de624},
  {32'h41617c70, 32'hc0f83e1a, 32'h41839b4d},
  {32'h44a34bb6, 32'h43135a42, 32'hc2ef7c42},
  {32'hc43aa34c, 32'h41f094bf, 32'hc4081d0f},
  {32'h450c32f4, 32'h41eb5e3e, 32'h4371be53},
  {32'hc4a6dce0, 32'hc32c6b0b, 32'hc3257e82},
  {32'h45068197, 32'h42052e93, 32'h434915f3},
  {32'hc481079f, 32'h433b505c, 32'h407a8c80},
  {32'h44e9e589, 32'hc2ea8b81, 32'hc2011458},
  {32'hc4d8d4e3, 32'hc39abeb2, 32'h4353d222},
  {32'h44ca46b3, 32'h41b53f75, 32'h42e8bf7e},
  {32'hc5065228, 32'hc302e01a, 32'h42e32b66},
  {32'h446c1ff9, 32'h42f77197, 32'hc389a643},
  {32'hc4abe53b, 32'h43bc7572, 32'hc3907284},
  {32'h4451c78c, 32'hc2906246, 32'hc404f810},
  {32'hc43c86cc, 32'hc2500eea, 32'h40ea745e},
  {32'h44b2e166, 32'hc39edfc5, 32'hc322714a},
  {32'hc4160162, 32'hc2d2f3c6, 32'hc1fe2fe9},
  {32'h44820aea, 32'h43324688, 32'h42a91752},
  {32'hc480abd4, 32'h439c55c1, 32'hc120f3d1},
  {32'h440b34f8, 32'h41c6ee9d, 32'h42bdaed2},
  {32'hc3a79038, 32'hc2e66efa, 32'h420cf925},
  {32'h44a6d109, 32'h4316c93b, 32'h42520560},
  {32'hc503e506, 32'h439c584e, 32'h4287b450},
  {32'h43fc9578, 32'h42748641, 32'hc0940385},
  {32'hc49a76a7, 32'h42377049, 32'hc2cf42a6},
  {32'h44589c98, 32'h4353ebd7, 32'hc2e1377a},
  {32'hc5043fa6, 32'hc37cb962, 32'h43b85fa5},
  {32'h442787f8, 32'hc36d8ac7, 32'h43728964},
  {32'h41867600, 32'h42980874, 32'hc41250aa},
  {32'h44e7c575, 32'h43036aee, 32'hc3e9de9c},
  {32'hc489633e, 32'hc28430dd, 32'h437660e8},
  {32'h441e078e, 32'h41ff1626, 32'h432c0c48},
  {32'hc3c13a3c, 32'hc359836f, 32'h42c963f1},
  {32'h430b5ce8, 32'h432f5b53, 32'hc3efecad},
  {32'hc33446f0, 32'hc33c8450, 32'hc1a3a1b0},
  {32'h44e0c5ad, 32'hc3a3feac, 32'h438e9756},
  {32'hc4afa8f1, 32'h422149c2, 32'h427a3f25},
  {32'h4392b65a, 32'h4379e7aa, 32'hc400e135},
  {32'hc400dfe8, 32'h42de0a6c, 32'h434a6257},
  {32'h4388ba8c, 32'h43820f76, 32'hc37a6b95},
  {32'hc516c930, 32'hc37d88c8, 32'hc38c2467},
  {32'h44fb2d95, 32'h42ae50a6, 32'hc15aefa5},
  {32'hc366634f, 32'hc05f2627, 32'hc397085f},
  {32'h44d94506, 32'h42536d81, 32'hc38972af},
  {32'hc4491a84, 32'hc2140dfd, 32'hc31149ea},
  {32'h43f41138, 32'h42c5065f, 32'h43011c66},
  {32'h4313f19c, 32'hc232286f, 32'h43956593},
  {32'h43a70c56, 32'hc31f41a3, 32'h4322dcea},
  {32'hc452a068, 32'hc1caae2a, 32'h43a20fc2},
  {32'h44eb48a8, 32'hc3a3e615, 32'h437b4330},
  {32'hc3952744, 32'h43c4d3c3, 32'hc2bb77d4},
  {32'h44f1efbc, 32'hc34772d5, 32'h42bc6bd1},
  {32'hc4af1ec1, 32'h4405a77b, 32'h42de51e5},
  {32'h441d2658, 32'hc30ca3cc, 32'hc36f913d},
  {32'hc32eb498, 32'h4303f874, 32'h4336592c},
  {32'h447c1cb0, 32'hc3dbf306, 32'h436ee295},
  {32'hc50ce549, 32'h43fa86b2, 32'h425b9f3d},
  {32'h44537d70, 32'h43ba2d02, 32'hc32740c2},
  {32'hc4de54d8, 32'hc269a8f6, 32'hc2b996a7},
  {32'h44e6cff4, 32'hc3a1e51a, 32'h433a216b},
  {32'hc4f7d164, 32'hc3b2b1e1, 32'h43765080},
  {32'h444b4c88, 32'h43128541, 32'hc3786291},
  {32'hc36e1e88, 32'hc31ba3e3, 32'hc3bf9fc9},
  {32'h4516ca91, 32'h4306d7c8, 32'hc1e9c3bc},
  {32'hc4e39f1e, 32'h419b9761, 32'h43284ac7},
  {32'h44d50a81, 32'hc32e4ee4, 32'h42eb0cd5},
  {32'hc47160d5, 32'hc258d2d2, 32'h439b1e4b},
  {32'h44535bae, 32'h43954516, 32'hc2a02cd8},
  {32'hc402b000, 32'h418b98b5, 32'h420f1eb0},
  {32'h44dd9734, 32'hc335d553, 32'h439b92b9},
  {32'hc5019119, 32'hc22fd981, 32'h400a2454},
  {32'h43882570, 32'h4315380b, 32'h4223a419},
  {32'hc502eb60, 32'hc3cd67e3, 32'hc2812f6b},
  {32'h4507a9d0, 32'h4389490d, 32'hc257b32c},
  {32'hc46bd6ca, 32'h439a2de0, 32'h42c5daf2},
  {32'h4511a62c, 32'h4206a9c2, 32'h42cd36b1},
  {32'hc421967c, 32'h4404a562, 32'h40d5ddfc},
  {32'h4525333e, 32'hc36d598b, 32'hc2582016},
  {32'hc4591692, 32'hc36420c3, 32'h435d760a},
  {32'h43414280, 32'h425230e2, 32'hc388bedc},
  {32'hc450e354, 32'hc2e3f278, 32'h436c624c},
  {32'h439f1c3e, 32'h43024e77, 32'hc31a0c86},
  {32'hc395ffb2, 32'h41f0a683, 32'hc3b0ab9c},
  {32'h4473ab64, 32'hc3ff6e40, 32'hc1fdc777},
  {32'hc4e5733c, 32'hc2c88881, 32'h439414e0},
  {32'h449ddb4c, 32'h4395be44, 32'hc38115f5},
  {32'hc3d5b461, 32'hc3a63e0e, 32'hc2c3ab49},
  {32'h44457e28, 32'h42f29ef8, 32'h43dfef71},
  {32'h4287bb60, 32'h42b8e234, 32'hc398412e},
  {32'h44ad174a, 32'hc09b1142, 32'hc10d5850},
  {32'hc40533c3, 32'h4346f227, 32'h42298997},
  {32'h44974f7e, 32'hc3015cb5, 32'h4251ffa7},
  {32'hc50b048a, 32'h432212aa, 32'hc3aa8a01},
  {32'h449d1653, 32'hc219df1f, 32'hc1cd68cc},
  {32'hc4beabe1, 32'h42b9e010, 32'h428942f4},
  {32'h451bc5f9, 32'hc27052a7, 32'hc375bc57},
  {32'hc4fc9501, 32'hc361133a, 32'hc288114f},
  {32'h45079faa, 32'h40fe696a, 32'h41711688},
  {32'hc3f313b8, 32'h420de917, 32'hc33eaa75},
  {32'h44dd43bf, 32'hc28903a2, 32'hc3b10c9e},
  {32'hc4fdda2c, 32'h4122474e, 32'h42503ef3},
  {32'h440d22e5, 32'hc3ae913b, 32'h43a8a669},
  {32'h4271213a, 32'hc3d319ca, 32'hc0c96f63},
  {32'h44f1fa06, 32'hc2e83eac, 32'h428c5c9b},
  {32'hc505ec60, 32'h4293c105, 32'h432c1d2d},
  {32'h44c43ec5, 32'h43b20264, 32'h40b75898},
  {32'hc497d79c, 32'h42b89fdc, 32'hc232b28a},
  {32'h435fcb80, 32'hc240074d, 32'hc2dbb366},
  {32'hc5049eec, 32'hc31da152, 32'hc32af44f},
  {32'h4508de8c, 32'h438dd95a, 32'hc27ce62b},
  {32'hc4b278cd, 32'hc32722aa, 32'h440fc763},
  {32'h44dd5f04, 32'h42be8c8c, 32'h42243b33},
  {32'hc50c769b, 32'h4291d598, 32'h43538335},
  {32'h44f86af2, 32'hc0a38f08, 32'h42bbdc07},
  {32'hc5102aa9, 32'hc24b26cf, 32'h43ecaad1},
  {32'h4511e326, 32'h42d408e2, 32'hc32edf9f},
  {32'hc4f21cc8, 32'hc3711380, 32'hc3872a12},
  {32'h449b3070, 32'hc2661319, 32'hc20ddc9c},
  {32'hc2477064, 32'hc1c85182, 32'hc397d5ec},
  {32'h44c72175, 32'h43396557, 32'hc2aefb83},
  {32'hc38a590c, 32'hc286d78a, 32'h43df4cf2},
  {32'h4344b1c4, 32'h433762cd, 32'h432f5734},
  {32'hc1d9c860, 32'h425ce7a2, 32'h439d0475},
  {32'h444788f5, 32'hc34a0ff3, 32'hc2991dad},
  {32'hc33491cb, 32'h4380d728, 32'hc2e45656},
  {32'h4420d6b6, 32'hc30e686f, 32'hc36a0a04},
  {32'hc50eda55, 32'h42e6f6f3, 32'hc1a45b6b},
  {32'h44ba9851, 32'hc3e52e48, 32'hc341f7ff},
  {32'h44ffdad4, 32'hc2232a36, 32'h431f6c48},
  {32'hc48b16a8, 32'h4284e1ad, 32'h41e75fa6},
  {32'h4462fbd6, 32'h3fb105d6, 32'h43ab12d4},
  {32'hc4bbae74, 32'h42ac589a, 32'h42c04cbe},
  {32'h44dff58b, 32'hc29f1306, 32'hc23f1d12},
  {32'hc478dcc7, 32'h4316cb93, 32'hc3ce1d12},
  {32'h43ab1388, 32'hc1848bd2, 32'hc3c5de4f},
  {32'hc0af0000, 32'hc2e8a901, 32'h438ec361},
  {32'h45012070, 32'hc2e89c6e, 32'hc389c675},
  {32'hc3f7022c, 32'h4393b8b2, 32'h4316d22c},
  {32'h44d01df5, 32'hc364ed34, 32'h40d1e6c9},
  {32'hc4b1d146, 32'h43b2adcd, 32'h43e34881},
  {32'h43d5e0a1, 32'h412ab273, 32'h433beada},
  {32'hc5182711, 32'hc1389a9a, 32'h424cc1b4},
  {32'h4417e2a7, 32'hc313d6f6, 32'h4395a855},
  {32'hc3d719ce, 32'h42ad5715, 32'hc149dcd5},
  {32'h44b42e3c, 32'hc108b10a, 32'hc3081d83},
  {32'hc48da8ba, 32'h429e8a65, 32'h42fc841a},
  {32'h452d5f41, 32'hc3397257, 32'h43ff9061},
  {32'hc45f513e, 32'hc260b84e, 32'h42a39d0c},
  {32'h44a89cdb, 32'hc3303868, 32'h42e7ad4c},
  {32'hc49ea655, 32'h433bb3ec, 32'h432f770d},
  {32'h44041b93, 32'h43840126, 32'hc2af47c8},
  {32'hc4c35ab3, 32'hc22e2200, 32'h42c1a576},
  {32'h4449836a, 32'hc2bcc936, 32'hbf47e77a},
  {32'hc43710bf, 32'h43944e7e, 32'h43bac122},
  {32'h449df09c, 32'h40806e9a, 32'h407a1660},
  {32'hc49ad104, 32'h438e68b4, 32'h43688032},
  {32'h4496122c, 32'h43419a8c, 32'hc4048337},
  {32'hc4d3f83e, 32'h43e79eef, 32'hc311abf9},
  {32'h448f28da, 32'h42913272, 32'h43a0bc35},
  {32'hc4b14fc6, 32'hc3ae285e, 32'h42918eb5},
  {32'h4442fcd4, 32'h431ffae5, 32'h4301accd},
  {32'hc4486964, 32'hc312de92, 32'h439194e3},
  {32'h44e90159, 32'h42edb0ca, 32'h429c98b1},
  {32'hc4ea47c7, 32'hc228e1af, 32'h42d165b8},
  {32'h44c402c6, 32'hc2b246b1, 32'h43538467},
  {32'hc5173e10, 32'h440a57c8, 32'hc222a1e8},
  {32'h44d7ab12, 32'hc387d527, 32'h428e1a24},
  {32'hc491cabe, 32'h42cbb322, 32'hc30cdd55},
  {32'h45047b9b, 32'h421b9a58, 32'h434b497d},
  {32'hc514db12, 32'hc34af919, 32'hc34decd5},
  {32'h44fa663d, 32'h43c10bd4, 32'h43aa46b1},
  {32'hc4d35984, 32'hc37750c8, 32'hc3b25074},
  {32'h4457ed86, 32'hc1b9a9c2, 32'hc36f589d},
  {32'hc2382e80, 32'hc21a36d6, 32'h4356f5d2},
  {32'hc1e6a1c0, 32'hc196671e, 32'h433c4844},
  {32'hc4988886, 32'hc3158aad, 32'h42620515},
  {32'h43618c50, 32'hc2303862, 32'h42b7f71e},
  {32'hc507bfbf, 32'hc3131f3f, 32'hc1b53771},
  {32'h443e8a02, 32'h4388e5df, 32'h431c91f5},
  {32'hc4f5e2e4, 32'h435d6d8f, 32'hc415e3b1},
  {32'h45045c79, 32'h42972c7d, 32'hc293e622},
  {32'hc505e557, 32'h41d0b8f8, 32'hc0907fe8},
  {32'h43b95f86, 32'h435434c4, 32'hc309ac23},
  {32'hc50a1c26, 32'h4366b915, 32'hc2976cbc},
  {32'h450a91d0, 32'hc2d9f035, 32'hc36e57bd},
  {32'hc49c4712, 32'hc3745b45, 32'hc2e944e7},
  {32'h450db8f4, 32'h434a5b9a, 32'h4382df41},
  {32'hc4ccbef2, 32'hc346eafe, 32'hc37bb4a1},
  {32'h4406689d, 32'hc2dbf67a, 32'hc3bc5365},
  {32'hc3cd4102, 32'hc155d554, 32'hc36a59ac},
  {32'h44f7fe0f, 32'hc18a3d52, 32'h43bdbf55},
  {32'hc3e8dce5, 32'hc1376056, 32'h440f9634},
  {32'h43f22d1d, 32'hc30a97d4, 32'hc35bef64},
  {32'hc46805e0, 32'hc1b246b2, 32'hc2062cc5},
  {32'h450ff2eb, 32'hc2840f62, 32'h423e076f},
  {32'hc4149847, 32'hc24d92d3, 32'hc31da80a},
  {32'h44a0ec7a, 32'h435cce87, 32'h43298331},
  {32'hc2becd20, 32'h42f7b252, 32'h43b6e566},
  {32'h44fe5c83, 32'hc3012894, 32'hc1b31850},
  {32'hc4c21ff1, 32'hc3a68e85, 32'h4313e2d5},
  {32'h43877cbc, 32'hc3b0b43d, 32'hc3b20a9d},
  {32'hc488e052, 32'hc306b17d, 32'h42d252b7},
  {32'h44e4c2f9, 32'h43d8f83d, 32'h42bb0137},
  {32'hc4c27436, 32'h42bc1920, 32'hc3a92717},
  {32'h43efa11c, 32'hc2b62627, 32'hc365741d},
  {32'hc3e06cf8, 32'hc1aa1a84, 32'hc3010c26},
  {32'h4505378a, 32'hc307e010, 32'hc1b2889e},
  {32'hc4928ec5, 32'hc2bae816, 32'h40e46644},
  {32'h45149447, 32'h42f39d31, 32'h43bc879a},
  {32'hc4d57a70, 32'h43cdc53d, 32'hc3b44436},
  {32'h44429d3a, 32'hc391c45a, 32'h43687c8d},
  {32'hc4234f5c, 32'h4282940d, 32'hc39f4a5a},
  {32'h450132ed, 32'h421f7ca0, 32'hc32f7eb9},
  {32'hc4f5fff4, 32'hc3208e07, 32'hc2f98b73},
  {32'h442e3965, 32'hc29b9cbf, 32'hc3817c2c},
  {32'hc3c56e38, 32'h435d1f39, 32'hc3058b95},
  {32'h44e292ef, 32'hc3cf7cb9, 32'h43427e91},
  {32'hc3882260, 32'hc35adb2c, 32'h42939dd4},
  {32'h448727c5, 32'hc417712b, 32'hc2bf174b},
  {32'hc48b48c7, 32'h435e4fc5, 32'h42f05fc1},
  {32'h429c702c, 32'h433d95b1, 32'h428ada7b},
  {32'hc41e58fd, 32'hc3597fe4, 32'h438ddff9},
  {32'h43bfc02b, 32'h4306aff2, 32'hc317f455},
  {32'hc41c5090, 32'h43230af0, 32'hc12ddd24},
  {32'h44b64792, 32'hc36e8803, 32'h424dfc39},
  {32'hc4a99a3b, 32'hc3f14ed5, 32'hc3b0d08e},
  {32'h444b4d01, 32'h43832b7b, 32'h432c4076},
  {32'hc4dd94e1, 32'hc3c334c0, 32'hc33f57b1},
  {32'h44e13d7d, 32'hc29e5ad1, 32'hc04b01a6},
  {32'hc3fb203c, 32'hc2a73a40, 32'h42b579c7},
  {32'h443038d0, 32'h44123cdd, 32'hc32c24ff},
  {32'hc4908274, 32'h43b40429, 32'h43198fd8},
  {32'h44e7d1e1, 32'h42e7e547, 32'hc396b07d},
  {32'hc4af5943, 32'hc32a3beb, 32'h436abca4},
  {32'h44687f64, 32'h434f43d5, 32'hc370fcfa},
  {32'hc3b7322e, 32'hc40ab53d, 32'h433b377d},
  {32'h44ac54bf, 32'hc255c3d3, 32'hc29a223c},
  {32'hc45d5148, 32'hc37bfbf8, 32'hc32062d8},
  {32'h43e6e748, 32'hc34c1a50, 32'hc316abe4},
  {32'hc48412e8, 32'h434d634d, 32'h44029772},
  {32'h44b81cc7, 32'hc2cb8a95, 32'h4369b047},
  {32'hc486d7fa, 32'h41f083ec, 32'hc3306e69},
  {32'h44d28b8e, 32'h3f501a30, 32'h430f3616},
  {32'hc4fe8646, 32'h42df7ac3, 32'hc1bd4d71},
  {32'h447245cb, 32'h43861576, 32'h42cc6f31},
  {32'hc38a318e, 32'hc300f6dd, 32'hc3ada8ec},
  {32'h448d3ab9, 32'h42fb42f2, 32'hc308c42a},
  {32'hc4ef5195, 32'h4262c0ef, 32'hc20ea6ed},
  {32'h448c01d5, 32'hc215e79d, 32'hc28706c5},
  {32'hc46e8a5c, 32'hc3d1796b, 32'h44271f9e},
  {32'h44634acf, 32'hc1d2868d, 32'h42d3e975},
  {32'hc48fa542, 32'hc3dc43da, 32'hc2740411},
  {32'h44efb17d, 32'h422c0d2f, 32'hc38369c5},
  {32'hc4ad9db9, 32'h4312673a, 32'h42d751d3},
  {32'h4401b11c, 32'h418d3a74, 32'h43937a66},
  {32'h42b1b920, 32'hc383e0ff, 32'h43406d8f},
  {32'h43974934, 32'h436a9fa7, 32'hc347cc8e},
  {32'hc3aab98a, 32'h434b9059, 32'h430bbaf1},
  {32'h44fdf061, 32'hc2fd4c5f, 32'h44132fb2},
  {32'hc40dc3d9, 32'hc36d38bf, 32'hbf6ebcc2},
  {32'h43c80d6b, 32'hc30f73e7, 32'hc39a39e0},
  {32'hc502ad5c, 32'hc2881492, 32'hc350fc6f},
  {32'h42fbb0a0, 32'hc2645c5f, 32'h42cbf5ba},
  {32'hc40200f0, 32'h429a7b06, 32'hc2eb92b6},
  {32'h42dcd290, 32'h42f1a01a, 32'hc3c44581},
  {32'hc43c036e, 32'hc2da7e9a, 32'h419f281b},
  {32'h43c3f496, 32'h438d2cb9, 32'hc2edba9b},
  {32'hc2aaad08, 32'h432592cc, 32'hc29fd720},
  {32'h43c60ea4, 32'h43865984, 32'h436696cf},
  {32'hc4c94a4d, 32'hbf54267c, 32'h4319451f},
  {32'hc33c04d6, 32'h435a4f5b, 32'hc2eae886},
  {32'hc4d72df0, 32'h4330804a, 32'h434ce891},
  {32'h43cc78a0, 32'h42916da6, 32'h436b9184},
  {32'hc4bd4b83, 32'hc1774251, 32'hc3c8482f},
  {32'h44fc0c14, 32'h43d411d8, 32'h43471f46},
  {32'hc4fce514, 32'hc3160297, 32'hc28ad955},
  {32'h44b4e3b0, 32'hc246c057, 32'hc25074b6},
  {32'hc4bb3288, 32'hc2a64b75, 32'hc3df369f},
  {32'h4471aeca, 32'h431d029b, 32'h4382da13},
  {32'hc4eb6fb3, 32'h4388df5b, 32'hc250b894},
  {32'h430fb308, 32'hbec38880, 32'h42210b05},
  {32'hc4b20d7c, 32'h433c8c6b, 32'hc318a52b},
  {32'h4505d505, 32'hc3200e40, 32'h4197864e},
  {32'hc4133cbf, 32'hc22ffd50, 32'h41fdff8f},
  {32'h448bb276, 32'hc34f6096, 32'hc399295d},
  {32'hc4fcd74f, 32'h41a4b6b3, 32'hc384c00b},
  {32'h44799bc6, 32'h42d2e3de, 32'hc2f15eb8},
  {32'hc4501374, 32'h43d82cea, 32'hc3084494},
  {32'h450628c1, 32'h4394d2d0, 32'h40bca7a3},
  {32'hc3ec51d6, 32'hc131bba0, 32'hc29b426a},
  {32'hc33a84f0, 32'h4354c81a, 32'h435b6613},
  {32'hc3edb5a4, 32'h439f1219, 32'hc27d8e4c},
  {32'h448643fc, 32'hc3051ad8, 32'hc2bf509d},
  {32'h41071180, 32'hc3876e3c, 32'h43d965f1},
  {32'h44808518, 32'hc3818374, 32'hc13a18e2},
  {32'hc490a122, 32'h439dab3b, 32'hc31027ff},
  {32'h439b14e3, 32'hc3a02466, 32'hc28d6e60},
  {32'hc44165fd, 32'hc3958c91, 32'h4212b05f},
  {32'h448701f7, 32'hc11e6c30, 32'h429c8996},
  {32'h42bd0600, 32'h42f0531a, 32'hc2fb285e},
  {32'h426150ec, 32'hc2ed05dd, 32'hc3e59ac0},
  {32'hc50f6e73, 32'h41cfed8e, 32'h429a84f7},
  {32'h4332bef8, 32'h42ad1c8b, 32'h424e7176},
  {32'hc4c5003e, 32'h43a34ba1, 32'h426a1bec},
  {32'h45008f52, 32'hc27cd57e, 32'hc3e77aec},
  {32'hc4c49289, 32'hc2c13721, 32'hc1da57d7},
  {32'h44a8fcff, 32'hc283c7fd, 32'h43726dfc},
  {32'hc4e83d03, 32'hc291e801, 32'h4332739e},
  {32'h44912078, 32'h42d18d12, 32'hc364c136},
  {32'hc3a46ba6, 32'hc3411d36, 32'hc3b4414d},
  {32'h45089bc0, 32'hc302453a, 32'h420e7fcc},
  {32'h42e4d060, 32'h43f4beed, 32'h42fc6764},
  {32'h4494b0d9, 32'h425934be, 32'h42d49beb},
  {32'hc40cbb1f, 32'h431606a0, 32'h42c2f684},
  {32'h4517052a, 32'hc376901c, 32'hc259113a},
  {32'hc41d90dc, 32'hc3740955, 32'hc2571fd5},
  {32'h452881b8, 32'h42e49d63, 32'hc2a6020c},
  {32'hc3f2e89c, 32'hc2c881ee, 32'hc352692c},
  {32'h42f6c524, 32'hc3239c7a, 32'hc3875f33},
  {32'hc3956d8b, 32'hc329c7f4, 32'h429e48c1},
  {32'h445da510, 32'hc39f6a24, 32'h42f1184a},
  {32'hc4afdbb9, 32'h420058be, 32'hc38cead5},
  {32'h447ce846, 32'hc38b311f, 32'h439f7cc7},
  {32'hc40ad04c, 32'hc27a14c0, 32'hc2ef2943},
  {32'h44fac298, 32'h436d5f9c, 32'hc2ac863b},
  {32'hc31aad50, 32'hc31471dc, 32'h41f8f5a7},
  {32'h44b2ad4e, 32'h42966f7b, 32'h436bcd6b},
  {32'hc4872f36, 32'h4156c7dc, 32'hc35e2d90},
  {32'h45041b49, 32'h42d920a5, 32'h41b6579b},
  {32'hc4e17660, 32'hc0e386aa, 32'h4389f749},
  {32'h450602b0, 32'hc34e834e, 32'hc1c0ba5d},
  {32'hc516c6d8, 32'h4341abb5, 32'h42bc1875},
  {32'h43cc17e4, 32'hc3bdda45, 32'hc34f4262},
  {32'hc3ac9d2f, 32'hc38ea76c, 32'h442273c8},
  {32'hc1818630, 32'hc3097576, 32'hc327078a},
  {32'hc32f4ec0, 32'h432c2da9, 32'hc32e11aa},
  {32'h44f39040, 32'h42c74072, 32'h435fa749},
  {32'hc4de2803, 32'h4246496a, 32'hc36f4371},
  {32'h43351758, 32'h43d3b19c, 32'h423c8828},
  {32'hc48a58b2, 32'hc3c59274, 32'h4395a122},
  {32'h448caaf0, 32'h43188856, 32'hc2632d99},
  {32'hc4ff8033, 32'hc1edbde9, 32'h42b70148},
  {32'h44684bd5, 32'h43030971, 32'h426a1da3},
  {32'hc43c56af, 32'hc4010080, 32'hc31aacb1},
  {32'h4302fb90, 32'hc27503b7, 32'hc2958516},
  {32'hc4fe248c, 32'h406b7a88, 32'hc2241342},
  {32'h44998a75, 32'hc35c643c, 32'h42d35f93},
  {32'hc342c47c, 32'h423fbb5a, 32'hc1792151},
  {32'h445c526d, 32'h42fd83e8, 32'h434ca41c},
  {32'hc1bb21b3, 32'hc2a1c5dc, 32'h42945082},
  {32'h43eadec4, 32'h43d67184, 32'hc246b4c6},
  {32'hc3a024a0, 32'hc35e6a40, 32'h425d5b64},
  {32'h43fa3a0c, 32'hc349981a, 32'hc2de5895},
  {32'hc4f5172d, 32'h43526474, 32'h43282281},
  {32'h44c150a2, 32'h427e94e6, 32'hc2e7dd83},
  {32'hc4dccb18, 32'h43e81ed8, 32'h4331ef7e},
  {32'h44282370, 32'h429517c0, 32'h42e680d0},
  {32'hc3512000, 32'hc34c41bb, 32'h42cef2d8},
  {32'h44cf1b11, 32'h4383be3d, 32'hc283dc7a},
  {32'hc3add9a6, 32'hc35c1452, 32'h42b5dffd},
  {32'h450e0896, 32'hc33fe332, 32'h43c2c6fa},
  {32'hc4a52ec6, 32'h431aaef1, 32'h436a2fd5},
  {32'h44330b37, 32'h427ccad4, 32'hc28fc58e},
  {32'h408de000, 32'hc2414d64, 32'hc21e147c},
  {32'h448db312, 32'hc2f646eb, 32'hc3597376},
  {32'hc50748f8, 32'hc2db40fd, 32'hc31eaabd},
  {32'h4427c6a4, 32'hc41a702e, 32'h43ea643a},
  {32'hc4cf54f9, 32'h429a9608, 32'h43dda33f},
  {32'h43ca82b0, 32'hc3481da2, 32'h429730c2},
  {32'hc4cb66a9, 32'h43336f4c, 32'h42f6ea1a},
  {32'h449f94ed, 32'hc2bb3da9, 32'hc33ef16e},
  {32'hc4fbe2a5, 32'h43ef2ef0, 32'h43c850fc},
  {32'hc26156b0, 32'hc240e4fc, 32'h4372dd5d},
  {32'hc2687694, 32'hc3c774fe, 32'hc2acdb20},
  {32'h444dfd7d, 32'hc25e28bc, 32'h3f3b469c},
  {32'hc4248826, 32'h430f47c7, 32'h43b99bf3},
  {32'h44cc5b08, 32'hc30dd480, 32'hc175bbda},
  {32'hc3708104, 32'hc28f4fe7, 32'h42cf136f},
  {32'h44f330cf, 32'hc2c3d5a3, 32'hc0b27709},
  {32'hc506885f, 32'hc217b941, 32'hc3b610a8},
  {32'h44fc8457, 32'h43a42e29, 32'hc33d3436},
  {32'hc4e04a27, 32'hc33f02ab, 32'hc291ff21},
  {32'h446c090f, 32'hc3ffa799, 32'h4201952c},
  {32'h4283f724, 32'hc392a8bc, 32'h42eff92d},
  {32'h439f8fc4, 32'h40a9df0a, 32'hc1adf097},
  {32'hc2d010d8, 32'hc10228b5, 32'h41886007},
  {32'h450ff130, 32'hc3097a73, 32'hc320902c},
  {32'hc4e4db8d, 32'h439c2772, 32'hc324475a},
  {32'h43c86919, 32'h432e845b, 32'hc352bab3},
  {32'hc4307601, 32'hc37eb339, 32'hc2706cd9},
  {32'h44dfea0f, 32'hc2b3c440, 32'h42dda80a},
  {32'hc4ca7434, 32'h43a4bca9, 32'h439184a2},
  {32'h44c2b4a4, 32'hc1cc520d, 32'hc15b1a5d},
  {32'hc3a753b4, 32'h41e7b716, 32'h437f7b3b},
  {32'h44f96354, 32'hc26e3f63, 32'hc31c1dee},
  {32'hc5072174, 32'hc261fb0b, 32'h435d8dd9},
  {32'h43a109e4, 32'h437407b3, 32'hc39f7441},
  {32'hc4ea1d49, 32'h42a78c10, 32'h43166ce2},
  {32'h44a4b3bd, 32'hc25c42c0, 32'hc2165c09},
  {32'hc3d02e56, 32'h42bb2dc5, 32'h4382df94},
  {32'h4501bca3, 32'h432e8f18, 32'hc38c1feb},
  {32'hc5037bad, 32'hc365403b, 32'hc34a8c47},
  {32'h450d0598, 32'hc3db4150, 32'hc4039ea1},
  {32'hc49cec88, 32'h438d1a65, 32'hc3313221},
  {32'h43ad9b0b, 32'hc37b2330, 32'hc2a78234},
  {32'hc501f5ae, 32'hc24b1782, 32'h4318d9ab},
  {32'h450f5426, 32'h42844b67, 32'hc26a1c5f},
  {32'hc50d5ebb, 32'h430b8bb3, 32'hc16e1060},
  {32'h4400fa83, 32'hc31bf75b, 32'hc1f6695a},
  {32'hc4488342, 32'h43cb68ec, 32'hc0ff0d6e},
  {32'h440f776c, 32'h4322063c, 32'hc337b68e},
  {32'hc3ca68e6, 32'h438abd39, 32'hc2f4b564},
  {32'h44b2a58c, 32'hc30dffa5, 32'h4316cd2a},
  {32'hc4b16d8c, 32'h430ea92c, 32'h43d97280},
  {32'h44b79a72, 32'h438a92ea, 32'h4362207b},
  {32'hc5057a69, 32'h4313a8aa, 32'h41969736},
  {32'h450e8705, 32'hc32a0d74, 32'hc3d44658},
  {32'hc5010f0e, 32'hc2a31d55, 32'hc3cb261b},
  {32'h4497c53c, 32'h4149eade, 32'hc3660d2f},
  {32'hc4132b45, 32'hc308a2db, 32'h43566f9a},
  {32'h43b925fa, 32'hc302aa77, 32'hc1d8201a},
  {32'hc41e1fae, 32'hc2b6d298, 32'hc19eecff},
  {32'h44e4bf35, 32'h431ff956, 32'h428d6a1f},
  {32'hc4eed4af, 32'hc2be6c7d, 32'hc2ab60b1},
  {32'h4512c591, 32'h42db0ed8, 32'h42fdb1c5},
  {32'hc45ec123, 32'hc4092f97, 32'h43903876},
  {32'h42d4fe10, 32'h430a3bb0, 32'h415627ce},
  {32'hc5132bff, 32'h42f334b4, 32'hc3824e9d},
  {32'h4316eb68, 32'hc20e979a, 32'h43c232d7},
  {32'hc376904b, 32'hc2714ac0, 32'h43a52d4f},
  {32'h446d722e, 32'h426fb0ff, 32'hc03f9bc8},
  {32'hc527bf66, 32'hc13e5283, 32'hc360fccc},
  {32'h443084cc, 32'hc295c65d, 32'h437097cb},
  {32'hc3e68778, 32'h43d236d6, 32'h43ffcf79},
  {32'h44e2813f, 32'hc209beed, 32'hc35f015a},
  {32'hc5077aaa, 32'hc2b1ee49, 32'h444d321c},
  {32'h40164000, 32'h42524b14, 32'hc1ac749e},
  {32'hc4c3780a, 32'hc23cfa6a, 32'hc26ed422},
  {32'h442cc4ac, 32'h429154f4, 32'h433ea0eb},
  {32'hc4f1b7c4, 32'hc24d7cac, 32'hc2ed809c},
  {32'h444750b7, 32'h438ff5b7, 32'h425bad2c},
  {32'hc48002ac, 32'hc1d4857a, 32'h439960f1},
  {32'h451870fa, 32'hc227e474, 32'h43caa250},
  {32'hc4916474, 32'hc3152034, 32'hc315cc48},
  {32'h450a3add, 32'h432be7e7, 32'hc3a14391},
  {32'hc48497bf, 32'h438c5998, 32'h430c074b},
  {32'h4461af5a, 32'h43cdf69b, 32'hc29c0174},
  {32'hc3dfd63a, 32'hc36fe9b8, 32'hc3b8bccb},
  {32'h443efc3a, 32'hc3838bb5, 32'hc321c137},
  {32'hc50a789e, 32'hc344bcbe, 32'hc213749f},
  {32'h43a06878, 32'h4380e2b9, 32'hc3c4ed67},
  {32'hc4a88d50, 32'h43048321, 32'hc3a9f157},
  {32'h42434b40, 32'hc391b451, 32'hc395d7ec},
  {32'hc4c915a7, 32'h4314aedf, 32'hc2dc54b0},
  {32'hc2b39fee, 32'h42cb7c76, 32'hc17bf6ae},
  {32'hc50e1434, 32'hc2982f53, 32'hc24fdc9c},
  {32'h45089ca0, 32'h4386cba4, 32'hc287d655},
  {32'hc4b22a79, 32'hc28ad094, 32'hc27281bc},
  {32'h44688c98, 32'hc344b262, 32'h43b6ecc8},
  {32'hc3e06708, 32'hc3403f94, 32'hc26cc827},
  {32'h44351c11, 32'h4368ec45, 32'hc400a59e},
  {32'hc4e34d04, 32'h42995e79, 32'h4398143c},
  {32'h44a12855, 32'h429e762c, 32'hc229148d},
  {32'hc4cea74a, 32'h43215394, 32'h402ed38f},
  {32'h450230fa, 32'hc2b3515c, 32'hc37a9660},
  {32'hc505fe7b, 32'h41c7f15f, 32'hc32186e2},
  {32'h4504124b, 32'h4386bcd1, 32'hc38e76b8},
  {32'hc4a9cd69, 32'hc0b6b2d0, 32'h42ee2f77},
  {32'h43283fd8, 32'hc38b3ae7, 32'h431363ff},
  {32'hc47949c4, 32'hc2498be7, 32'hc34c5b5a},
  {32'h44fe6f45, 32'hc2593622, 32'hc2eed124},
  {32'hc38b9a88, 32'h4393efef, 32'hc302f9bd},
  {32'h44a347b6, 32'hc38c34aa, 32'h425f8af9},
  {32'hc40c9718, 32'hc3579126, 32'hc204bf53},
  {32'h4438d60f, 32'h42ca6ee2, 32'hc3711cec},
  {32'h41282840, 32'h43c25683, 32'h437dfc53},
  {32'h44d03ff6, 32'h43353324, 32'h41de4774},
  {32'hc3c46916, 32'hc2a9b168, 32'h42b8ab8a},
  {32'h4482c005, 32'hc2e2ade4, 32'h43908530},
  {32'hc4a01f37, 32'hc3d789c4, 32'h4397b7b8},
  {32'h44943858, 32'hc306a850, 32'h4111f1d4},
  {32'hc35e56b8, 32'hc2e51c0d, 32'h438e8d10},
  {32'h44a907f1, 32'h43739145, 32'h43a45342},
  {32'hc4aa9383, 32'h4105f9f2, 32'hc2a51c0a},
  {32'h44358f9e, 32'h4384bb75, 32'hc2f34fa2},
  {32'hc5038857, 32'hc35e80af, 32'hc36e0ef2},
  {32'h44eda184, 32'hc324fdf7, 32'h41ab89c2},
  {32'hc32560ec, 32'hc32ceebc, 32'h41b4d714},
  {32'h440045d4, 32'h4318049c, 32'h43f55d1e},
  {32'hc426daef, 32'h420bb500, 32'hc32ca787},
  {32'h4506eb54, 32'hc310f54a, 32'h42fca866},
  {32'hc4b02caa, 32'h42a2e4ce, 32'hc33821da},
  {32'h450b0fbe, 32'hc2333b2a, 32'h44002387},
  {32'hc507b5ca, 32'hc21b849b, 32'h4335bd7f},
  {32'h44696687, 32'h42d437db, 32'hc2fd96b0},
  {32'hc501d6d5, 32'hc3332e0a, 32'hc08ed98f},
  {32'h4522266a, 32'h43323a0d, 32'h437e24e0},
  {32'hc4ac91a4, 32'hc2a5e3d9, 32'hc373e521},
  {32'h434d724e, 32'h42963d21, 32'h43f899bf},
  {32'hc4be4fda, 32'hc32e3686, 32'hc35a08a3},
  {32'h4492a2de, 32'h3e7c87b0, 32'hc3049c6f},
  {32'hc4d91f38, 32'h4096963f, 32'h436708f1},
  {32'h44dc6887, 32'hc2e5c1ae, 32'hc2c506a8},
  {32'hc4ec2417, 32'hc2e5471a, 32'h433e1362},
  {32'h4391123a, 32'hc3065bf5, 32'hc329399b},
  {32'hc389abcc, 32'hc377da97, 32'hc30e4e1d},
  {32'h4501aeb5, 32'hc32edc84, 32'hc2abdb18},
  {32'hc45a9d5c, 32'hc3a31b77, 32'h43228f75},
  {32'h450d33ee, 32'hc2da7b56, 32'hc2bdf9e1},
  {32'hc4b2228c, 32'h42d139ba, 32'hc38babe9},
  {32'h446ae9ba, 32'hc348f6e0, 32'hc1b6a39e},
  {32'hc4fd745e, 32'hc2cc4b00, 32'h43ab072f},
  {32'h442dc524, 32'h42b878f6, 32'h42f39e4f},
  {32'h430081aa, 32'hc324dfb2, 32'hc2b92e60},
  {32'h44a15f76, 32'hc3987328, 32'h429bb6a8},
  {32'hc4f47d28, 32'h43683dfe, 32'h435a4790},
  {32'h450668cf, 32'h42c94b01, 32'hc1bed99d},
  {32'hc50d8f43, 32'h42b6cb73, 32'h436cf59f},
  {32'h44470b82, 32'h43596a95, 32'h431b8b8e},
  {32'hc445eb3a, 32'h429f246e, 32'h4350a8e7},
  {32'h448127ba, 32'hc202e840, 32'hc34f821b},
  {32'hc45636b3, 32'hc2e5e875, 32'hc32a11e9},
  {32'h44ed7cef, 32'h43cf99a5, 32'hc3811d03},
  {32'hc43636f7, 32'h4209efe5, 32'hc3b55455},
  {32'h44f24648, 32'hc35c1824, 32'hc1e80cf7},
  {32'hc4cf2793, 32'h432705d4, 32'hc30471c2},
  {32'h4381f684, 32'h4398e2a0, 32'h430f8399},
  {32'h4334fb30, 32'hc3095072, 32'hc1936896},
  {32'h450e03e1, 32'h41ca986f, 32'hc294a4ca},
  {32'hc50c271d, 32'hc3aca22c, 32'hc34dd688},
  {32'h4500e0bd, 32'hc26cd34e, 32'h4352b22a},
  {32'hc51e2502, 32'hc3ee1379, 32'hc1e7875e},
  {32'h45082f5b, 32'h42dcb2aa, 32'h43ec9efa},
  {32'hc4b4ec34, 32'hc2e3a0de, 32'hc22a09d5},
  {32'h44bb7a41, 32'hc2e613ab, 32'h436689a5},
  {32'hc4daf6ea, 32'hc390ea30, 32'hc1ea353d},
  {32'h44aec379, 32'h4166e226, 32'h43482b07},
  {32'hc3980165, 32'hc32605b6, 32'hc2aecb35},
  {32'h432a8ed0, 32'hc3f65829, 32'h43aaff11},
  {32'hc4c7e764, 32'hc3cb6f2e, 32'h419b10cd},
  {32'h44aa41a4, 32'hc309d601, 32'hc1b7c904},
  {32'hc491fa04, 32'h439c4ea5, 32'hc25cc9bd},
  {32'h4410ec96, 32'hc389ea50, 32'h438878cb},
  {32'hc4a9bced, 32'hc37230ea, 32'hc3a19020},
  {32'h4495a9fa, 32'h439e05a1, 32'h4394eaa1},
  {32'hc4917f06, 32'hc22d3a9f, 32'hc213a524},
  {32'h44650e22, 32'hc353f142, 32'hc21398e6},
  {32'hc4a65502, 32'hc392ed66, 32'h42a15411},
  {32'h449e5cc7, 32'h4305e002, 32'h4393fbe4},
  {32'hc28f2d30, 32'h43716007, 32'hc2c39cf2},
  {32'h43c33754, 32'hc2d3fbdd, 32'h43101c43},
  {32'hc40b05c8, 32'hc3078a73, 32'hc3741e52},
  {32'h43534060, 32'h4217018e, 32'hc2b1af31},
  {32'hc46638cd, 32'hc1771fa1, 32'hc220572f},
  {32'h43699ac0, 32'hc300446f, 32'h4021a4b7},
  {32'hc3ad371c, 32'hc1f437be, 32'hc38ea4c8},
  {32'h4458ecb4, 32'h43ad3b0b, 32'h43921465},
  {32'hc498a235, 32'hc2a378f2, 32'h43578865},
  {32'h4436ae5a, 32'h42934cee, 32'hc2b81aeb},
  {32'hc49fad4b, 32'hc32c71e9, 32'h40d3facc},
  {32'hc4b9b42b, 32'hc2a798d7, 32'h4343e003},
  {32'h44ddce96, 32'h43ad7149, 32'h40efc8dd},
  {32'hc4eb63c8, 32'h41dfb3cb, 32'hc3abca2d},
  {32'h43d458dc, 32'h42572481, 32'h436c1940},
  {32'hc4102025, 32'hc2c1b09f, 32'hc3f48200},
  {32'h4419b5c6, 32'hc37d9187, 32'h43bab214},
  {32'hc424a041, 32'hc2da8977, 32'h4340b0bc},
  {32'h449390f2, 32'h40db507c, 32'h4291d468},
  {32'hc40212c4, 32'hc2cb7bb2, 32'h414fe8d6},
  {32'h43cc07bc, 32'hc218d364, 32'h42aae6a3},
  {32'hc4bd281c, 32'h43b52752, 32'hc3193b1f},
  {32'h44bd5052, 32'hc2041695, 32'hc30d9df6},
  {32'hc47a5dc2, 32'h44072c31, 32'hc2458d75},
  {32'h4439dd0d, 32'hc2bcef8c, 32'h411b75bf},
  {32'hc504c08f, 32'hc38630fe, 32'hc32f9f4e},
  {32'h450c03f1, 32'h431dc0f1, 32'h4232de0b},
  {32'h42f851fe, 32'h439a7169, 32'hc398d7ec},
  {32'h43b0cbf4, 32'hc30dff0a, 32'h43a527dc},
  {32'hc4e18b8e, 32'h426e3139, 32'h43044304},
  {32'h449075a4, 32'hc140f875, 32'h43b18b94},
  {32'hc50dfb21, 32'hc35e720c, 32'hc21c1b8d},
  {32'h44e88012, 32'hc22db760, 32'hc2c1ff08},
  {32'hc4d7f0d9, 32'h439a0f81, 32'hc4073448},
  {32'h44fee44a, 32'h4140470b, 32'hc357f9e4},
  {32'hc4f04f36, 32'h42fe17e3, 32'hc2fdc024},
  {32'h43426e66, 32'hc41fa5eb, 32'h430ca62b},
  {32'hc47a2aae, 32'h429d61e5, 32'h43ab094e},
  {32'h449478f7, 32'h4229f03a, 32'h41fa553a},
  {32'hc456fd12, 32'h433b1ddd, 32'hc37afc12},
  {32'h44b857d4, 32'hc3a8c487, 32'h41c0be99},
  {32'hc5007136, 32'hc34b1d72, 32'hc31a8391},
  {32'h44cb7c1c, 32'hc3a82e63, 32'h4285f49d},
  {32'hc477246d, 32'h424269d6, 32'h4324ee8a},
  {32'h44aa970f, 32'h43a72129, 32'h428634a5},
  {32'hc4543e26, 32'hc3e77260, 32'hc3cc04b7},
  {32'h43b2fa68, 32'hc3cd5c13, 32'h4259ba0a},
  {32'hc4c6cb43, 32'hc3609f3a, 32'hc2dff254},
  {32'hc1df7a00, 32'h43945804, 32'h433808c0},
  {32'hc43a4246, 32'hc200741a, 32'hc3362edb},
  {32'h43825e42, 32'h43a0040b, 32'hc34dbca8},
  {32'hc4499fae, 32'hc1b92d36, 32'h42fb5dc1},
  {32'h440f1664, 32'h42093ba2, 32'h43bd6290},
  {32'hc4c52188, 32'hc2721e7c, 32'hc39310b0},
  {32'h4517a2de, 32'h42bd50a6, 32'hc36b352f},
  {32'hc410b4aa, 32'h41688636, 32'hc368cd1a},
  {32'h44ddcbf4, 32'h4391e8a6, 32'hc3233f06},
  {32'hc51d5eb8, 32'h43ae30ba, 32'h412c85e3},
  {32'h42c04660, 32'h429036ff, 32'hbe790960},
  {32'hc41f6e02, 32'hc1c4097b, 32'h42933705},
  {32'hc1ff0f80, 32'h43031f16, 32'h42cca13f},
  {32'hc50ec42a, 32'h43d04626, 32'hc3acdca4},
  {32'h44fad05c, 32'h42a4d0c3, 32'hc331bc7b},
  {32'hc4dc397e, 32'hc34969fd, 32'hc36dd905},
  {32'h4503a862, 32'hc305a3c0, 32'h43120934},
  {32'hc41adfbe, 32'hc290aa7c, 32'hc37226fb},
  {32'h448e3ede, 32'hc2bb28a4, 32'hc339ccf5},
  {32'hc5159bbc, 32'h42cdab84, 32'hc385a3e0},
  {32'h44f5289e, 32'h4318d024, 32'h429bbf6d},
  {32'hc518021c, 32'h438764fd, 32'hc3753ddb},
  {32'h450eccd3, 32'hc347df17, 32'h434bc311},
  {32'hc4d48120, 32'hc3ebf297, 32'hc395ce72},
  {32'h44dba36c, 32'hc30471c4, 32'h41c80ebb},
  {32'hc4fe0893, 32'h441a7e95, 32'hc309e216},
  {32'h44af26ac, 32'hc33beab0, 32'hc3246d37},
  {32'hc41cb4e1, 32'hc288bea6, 32'h42fc40bb},
  {32'h4487f32a, 32'hc3894b90, 32'h427f1ec2},
  {32'hc50a8159, 32'hc2d665ce, 32'hc252811b},
  {32'h4490f7ae, 32'h4272a9b1, 32'h4372ddd3},
  {32'hc41a96ea, 32'hc34c3c08, 32'hc31c9de8},
  {32'h448d74da, 32'h43a19ed9, 32'h4384bb89},
  {32'hc4c25675, 32'hc2d3ced4, 32'hc2030a75},
  {32'h44a13b2e, 32'hc24137b4, 32'h439b3d90},
  {32'hc46aced4, 32'hc193a80c, 32'h42ee2267},
  {32'h44d27016, 32'hc24e9504, 32'h4203837f},
  {32'hc4c2a9c8, 32'hc31f1fd8, 32'hc327c877},
  {32'h44f8c1e8, 32'h439cd111, 32'h40d8e050},
  {32'hc45edc53, 32'hc3e5fab5, 32'h42c3087d},
  {32'h451abfc8, 32'hc1f6d57e, 32'hc2dd7e76},
  {32'hc4653c5e, 32'hc3926d8e, 32'h427783f1},
  {32'h44e34120, 32'h4242b7e6, 32'h439e37bb},
  {32'hc49bf454, 32'hc3b68e39, 32'h42b17ea5},
  {32'h44c517b2, 32'hc3d5e3a8, 32'h43e0a074},
  {32'hc4ae6c1b, 32'hc242d66a, 32'hc329a57d},
  {32'h45038b6a, 32'hc3fa0750, 32'hc326d926},
  {32'hc50becb9, 32'h43493df0, 32'h42faf8c6},
  {32'h44ff0c7a, 32'h4388e76a, 32'h43a838c4},
  {32'hc4938327, 32'h43a2a836, 32'hc2d5c7d5},
  {32'h44dec15d, 32'hc34eb1a1, 32'hc36226fa},
  {32'hc47c914a, 32'h42e8c5b9, 32'h4316b7c3},
  {32'h4487c381, 32'h430f9083, 32'hc261d046},
  {32'h43278ee8, 32'h42172f0b, 32'h42a4de4c},
  {32'h440a7c48, 32'hc267f948, 32'hc22e4a70},
  {32'hc3977b84, 32'hc3753f7e, 32'h42db635d},
  {32'h44933802, 32'h4257f931, 32'h43bc4cee},
  {32'hc3daf4e4, 32'hc24c4bb3, 32'hc2d98af5},
  {32'h4380f560, 32'hc395adca, 32'hc2a9a880},
  {32'h4321f80d, 32'h43c6f56a, 32'hc30920ab},
  {32'h442527f2, 32'h43a87fa2, 32'h4284a60e},
  {32'hc3790e00, 32'h43eebb3c, 32'hc26f7748},
  {32'h45190b79, 32'h42c1cc35, 32'h44013165},
  {32'hc4b3f2cb, 32'h4255130d, 32'h43cc7c87},
  {32'h45068bd8, 32'hc2d27fef, 32'hc229f7c8},
  {32'hc32e3ba0, 32'hc0fdad04, 32'h4341af42},
  {32'h44f12afc, 32'h430090be, 32'h43ecd828},
  {32'hc4c8ab4e, 32'hc2ab274b, 32'h439177e0},
  {32'h449e83c0, 32'h43768afd, 32'hc2062d34},
  {32'hc234ad12, 32'hc29ecf27, 32'hc3b79066},
  {32'h43b0e478, 32'hc2718e32, 32'h435bc6e7},
  {32'hc4f871d8, 32'h43ce8452, 32'hc237366a},
  {32'h44964f65, 32'h431ff2b0, 32'h418c6015},
  {32'hc40a7ec3, 32'hc2991914, 32'h432800b8},
  {32'h447ef271, 32'h42e3543d, 32'h434d4640},
  {32'hc4f4d990, 32'hc378da6e, 32'h43cd11a0},
  {32'h442c5d9e, 32'h432f674a, 32'hc2bd7d60},
  {32'hc508795c, 32'hc3b8becd, 32'h441c1909},
  {32'h4518b6f3, 32'h42afd8a4, 32'hc398b22d},
  {32'h438ac145, 32'hc34be812, 32'hc1f4b69e},
  {32'hc350ef8b, 32'h41eb39a4, 32'h42f3a2cf},
  {32'h450163ee, 32'hc06d3024, 32'hc305862c},
  {32'hc26decc0, 32'h42f65961, 32'h43133a43},
  {32'h446fffea, 32'hc40e7bfe, 32'h4321e51b},
  {32'h42e1b978, 32'h43128b99, 32'h4341896a},
  {32'h43b260f0, 32'h43d24e92, 32'h42b2225a},
  {32'hc4b9fc38, 32'h439c0f38, 32'hc2f77ab0},
  {32'h4467912c, 32'h43540318, 32'h42fcfc57},
  {32'hc49eed91, 32'h426e8fe1, 32'h4230dfac},
  {32'h44847f06, 32'h42ef7356, 32'hc39cde51},
  {32'hc4e23b6f, 32'hc2bd8152, 32'h43a53fc0},
  {32'h44347936, 32'h42c1f808, 32'h435ca324},
  {32'hc45b625c, 32'hc327ef12, 32'h43c11dcc},
  {32'h43ca21b0, 32'hc2ba5afc, 32'h43090731},
  {32'hc44d5bbc, 32'h43a645bb, 32'h425265ae},
  {32'h4393e478, 32'h42c2eeac, 32'hc1c3989e},
  {32'h437763f8, 32'h4343c45a, 32'h436e93c4},
  {32'hc325a860, 32'hc301e16f, 32'hc2f3c332},
  {32'hc40d1632, 32'h43e4c79b, 32'h439086f8},
  {32'h42a18630, 32'hc2775881, 32'h42cd45cb},
  {32'hc419114d, 32'hc2fd71f2, 32'hc31d4900},
  {32'h44dd34f2, 32'h43b3861a, 32'hc3472592},
  {32'hc4e8ccb6, 32'h4386fe2a, 32'h42b77ccd},
  {32'h44a3d9f8, 32'hc32d5d1c, 32'hc31922fd},
  {32'hc4cae989, 32'hc2db3050, 32'h4358c02d},
  {32'h43312240, 32'hbf859ae9, 32'hc37265ec},
  {32'hc414642a, 32'hc1dd3272, 32'hc2d0138b},
  {32'h43f0ba35, 32'hc2b608d8, 32'hc3230258},
  {32'hc4924f58, 32'hc2adf818, 32'h431e82fa},
  {32'h44bb8bc0, 32'hc30d11da, 32'hc379657b},
  {32'hc2e63c60, 32'hc2b792da, 32'h43806dee},
  {32'h44e033d3, 32'hc2f8ec95, 32'hc2bcd472},
  {32'hc46208de, 32'h42f7d986, 32'hc384ca44},
  {32'h4398624a, 32'hc4181a03, 32'hc31c1c3d},
  {32'hc48bcbb2, 32'hc2008ff2, 32'hc301e4de},
  {32'h44b6e8de, 32'hc31699c2, 32'h432970e5},
  {32'hc47a8c03, 32'h43a0e5c4, 32'h425cce8f},
  {32'h43a36440, 32'hc2d1846c, 32'hc2b8eee5},
  {32'hc49bf9f4, 32'h43433631, 32'hc3967dde},
  {32'h45037cd8, 32'h43a5f556, 32'h4308d23e},
  {32'hc501f92c, 32'h43a14382, 32'hc13435bf},
  {32'h44ca0b97, 32'hc38ab850, 32'hc1789cf0},
  {32'hc43963a1, 32'hc314217d, 32'hc322af07},
  {32'h44f9841e, 32'hc1fab56d, 32'hc2521d58},
  {32'hc38c4a8c, 32'hc2a2dc72, 32'hc24b950a},
  {32'h44bdb2fa, 32'hc28dc738, 32'hc2e7c9c2},
  {32'hc4296a0e, 32'h432f4162, 32'h431a6768},
  {32'h4452be90, 32'hc2121e3c, 32'hc28e0868},
  {32'hc43a99be, 32'h42b0133f, 32'hc3841316},
  {32'h43e49e20, 32'hc3d25b6e, 32'hc31528ea},
  {32'hc50bb71f, 32'h43515435, 32'hc3527866},
  {32'h43b4914e, 32'h422ecdfd, 32'hc381ca4f},
  {32'hc4409cc2, 32'h42f849fa, 32'hc3a1054f},
  {32'h43a2a4f8, 32'hc2c3fcbd, 32'hc327beca},
  {32'hc2380880, 32'hc33057f8, 32'hc211f5bc},
  {32'h434efa78, 32'hc315b290, 32'hc30dedc3},
  {32'hc4de38a0, 32'hc38d4c94, 32'hc3d22c78},
  {32'h44b7f303, 32'h43d5f55b, 32'h43a05048},
  {32'hc4659941, 32'h4320a797, 32'hc2402ed6},
  {32'h449568c9, 32'h426ebc60, 32'h42463d2c},
  {32'hc4ec3ee6, 32'hc1feb548, 32'hc30f6da4},
  {32'h446496f2, 32'hc302b2cb, 32'h437242ea},
  {32'hc4c79e8a, 32'hc2b4b125, 32'h42e9c3c3},
  {32'h43f6ff68, 32'h42dead10, 32'hc2e410c1},
  {32'hc41cd596, 32'hc341e8f3, 32'hc2b6db4b},
  {32'h44a7565d, 32'h43ae904b, 32'h437e4da7},
  {32'hc4cea229, 32'hc2b33033, 32'h432a6d9b},
  {32'h44342ed4, 32'h43162e64, 32'hc26e2b5a},
  {32'hc4bbe3b8, 32'h42685a58, 32'h43328623},
  {32'h43e1dbad, 32'h42d8310e, 32'h42657617},
  {32'hc4544fba, 32'hc3bf3bab, 32'hc38e78a8},
  {32'h44cc9485, 32'h42c3b3ae, 32'hc34e0243},
  {32'hc4c9417b, 32'hc30f7d93, 32'h428c2401},
  {32'h44a23d73, 32'hc335663a, 32'hc1bd7afe},
  {32'hc3ab60ac, 32'hc36677e3, 32'hc280e397},
  {32'h44404cb7, 32'hc2032250, 32'h430a4f03},
  {32'hc4cd2756, 32'h42f3c935, 32'hc18b18d2},
  {32'h44bff826, 32'h434e8ba0, 32'hc3d91dda},
  {32'hc501fd2d, 32'hc31bd9fe, 32'hc39d94ef},
  {32'h43bec3b0, 32'h42a60936, 32'h42c08482},
  {32'hc40f6de8, 32'h42bd5ad9, 32'h43c50d89},
  {32'h44afeb37, 32'hc0505ab2, 32'h42a6dafe},
  {32'hc407cdd2, 32'h430a4c9d, 32'h429bfa2f},
  {32'h441268e5, 32'h40911545, 32'hc29a0790},
  {32'hc4c92ca4, 32'hc11af72b, 32'h42d2b165},
  {32'h44e8ec60, 32'h4214acbd, 32'hc2dd1b92},
  {32'hc4391493, 32'hc30eaf25, 32'h43c0fe48},
  {32'h450eadad, 32'hc365b16e, 32'hc1d99958},
  {32'hc4cf30b0, 32'h43834507, 32'hc2d1751f},
  {32'h450c3a90, 32'hc213a40a, 32'h42d97437},
  {32'hc4b33da0, 32'hc387fed6, 32'h4363f78f},
  {32'h446e5e8c, 32'hc1f185f5, 32'hc173cf5c},
  {32'hc4bf321c, 32'hc3422fda, 32'hc2dd29d7},
  {32'h44a4abc0, 32'h42343548, 32'hc20b5c66},
  {32'hc4305227, 32'h4356a010, 32'hc2f5568c},
  {32'h44bbef3a, 32'h42cfe451, 32'hc2169e41},
  {32'hc511448e, 32'hc14bb7d1, 32'h416196aa},
  {32'h4517a283, 32'hc33605d3, 32'hc33a3971},
  {32'hc4f83454, 32'hc3991d11, 32'hc37dc265},
  {32'h43d9b060, 32'hc3ae4280, 32'h43e8d5aa},
  {32'hc2a0da08, 32'hc325b681, 32'hc32d071e},
  {32'h448eb094, 32'h4303dcdb, 32'h439bd407},
  {32'hc43021ec, 32'hc3833794, 32'h43314efb},
  {32'h44e2c082, 32'h43c0c164, 32'hc32e76c3},
  {32'hc42c8c2b, 32'h4259ecab, 32'hc394b403},
  {32'h44f929ef, 32'h43171709, 32'h417c29f9},
  {32'hc487b80a, 32'hc3856466, 32'hc3a35bff},
  {32'h44229304, 32'hc34d7f1c, 32'hc20e61fc},
  {32'hc448ce06, 32'hc385b97c, 32'hc393bf31},
  {32'h448a4a34, 32'hc01f46a0, 32'hc3804991},
  {32'hc503c241, 32'hc3acb5fe, 32'h42c8f7fc},
  {32'h44c10e39, 32'hc381ebaa, 32'hc24c801d},
  {32'hc4a6ffdc, 32'h43f05963, 32'h437e361a},
  {32'h44c0be14, 32'hc1f35cd3, 32'hc3e6b0d1},
  {32'hc4cce99e, 32'hc296abff, 32'h41debec0},
  {32'h445c480e, 32'hc157ae8a, 32'hc3699714},
  {32'hc4057839, 32'h42836ffb, 32'hc2c1521d},
  {32'h44a356d6, 32'hc3ccdd4f, 32'h430bd9cf},
  {32'hc3b06ac0, 32'h43954d89, 32'hc20f3104},
  {32'h448ba42a, 32'h42ce53a1, 32'hc294be90},
  {32'hc4f61c88, 32'hc270734b, 32'hc2fd72d7},
  {32'h449797f0, 32'h4295403c, 32'h433363fe},
  {32'hc4786aee, 32'h42d9f7c5, 32'hc300cf49},
  {32'h4435b082, 32'hc36a3e6e, 32'h423b9235},
  {32'hc4e0d5be, 32'hc2b02087, 32'h43661db0},
  {32'h41c5a060, 32'h42e54311, 32'hbec330b7},
  {32'hc4ead405, 32'h42ad90ce, 32'h4332c5e2},
  {32'h442a9ac2, 32'h43530266, 32'hc0c2135e},
  {32'hc2e8bd20, 32'h41806a26, 32'hc3858b76},
  {32'h450efca2, 32'hc400c0c2, 32'hc3c8d520},
  {32'hc4049cc5, 32'h42e4cfd9, 32'h42a4ba9d},
  {32'h44a66889, 32'h4397aef9, 32'h41480199},
  {32'hc4c1289e, 32'h43b80af5, 32'hc2094f56},
  {32'h443b9d18, 32'h43a3402e, 32'hc3b257e7},
  {32'hc4a916d4, 32'hc3860cc4, 32'hc30b53ad},
  {32'h450bf1a0, 32'hc26e6e52, 32'hc3d732c2},
  {32'hc485eb54, 32'hc2b70c42, 32'h428206a7},
  {32'h441af64c, 32'h43b80802, 32'h430fe3a7},
  {32'hc4c7cd5f, 32'hc3d7aed7, 32'hc37ef696},
  {32'h44bc9b26, 32'h431fa39a, 32'h40d2ba69},
  {32'hc4b535ca, 32'h435eedb9, 32'hc2e3bfc4},
  {32'h44a28930, 32'h43978ede, 32'h424838d8},
  {32'hc39b2580, 32'hc3596ade, 32'hc34995ed},
  {32'h44bbfef9, 32'h432fc3af, 32'hc2f68d72},
  {32'hc4be3e6a, 32'h42ed659b, 32'hc2fa6786},
  {32'h43c82e3a, 32'h43d00757, 32'h437ae961},
  {32'h412a1940, 32'hc32e952a, 32'hc1d76530},
  {32'h440b0253, 32'h433b8972, 32'h4137b378},
  {32'hc4b0c373, 32'hc31de6b0, 32'h43203bbc},
  {32'h42b45490, 32'h42b9ee31, 32'h427e2217},
  {32'hc496456a, 32'h43434253, 32'hc180fcfd},
  {32'h4315f7d0, 32'h43444583, 32'hc349e0a2},
  {32'hc4a275d1, 32'h418aec50, 32'h43c4b91a},
  {32'h44f1f2c4, 32'hc2a8348c, 32'h431946ba},
  {32'hc503154b, 32'h42b5fe2f, 32'h430a659e},
  {32'h44f304ee, 32'hc336049d, 32'hc147cd92},
  {32'hc50f9bb3, 32'hc10949cb, 32'h42e457c6},
  {32'h43f70f42, 32'hc130a14a, 32'h43207bbf},
  {32'hc4849d42, 32'h4098206a, 32'h421df9fd},
  {32'h44eb4e00, 32'h42234666, 32'hc33508c8},
  {32'hc51fbc2f, 32'hc30da850, 32'hc395deca},
  {32'h4527340e, 32'h42449ab2, 32'h43b2e5a4},
  {32'hc3d6e00c, 32'h4417500a, 32'h41137aca},
  {32'h448ca7cf, 32'h40a0d744, 32'hc31667ba},
  {32'hc4853154, 32'h42c88671, 32'hc2f1918a},
  {32'h4462a9d0, 32'hc305e9c4, 32'h42e307d4},
  {32'hc3b4e8aa, 32'hc2deba54, 32'h43caffd4},
  {32'h44edcd4a, 32'hc29926d1, 32'h4391fa96},
  {32'hc4372214, 32'h43a3e733, 32'h43432164},
  {32'h4440bbee, 32'h4372d896, 32'hc1ba0ec5},
  {32'hc3a07ae0, 32'hc36361e2, 32'h434639f6},
  {32'h4511466f, 32'hc2ee6b09, 32'h424f16e9},
  {32'hc4b18230, 32'hc2f7ca05, 32'hc310068b},
  {32'h44aac29f, 32'hc226f65e, 32'h42862a88},
  {32'hc39f9d6b, 32'h42f0d93b, 32'h42a6b9cb},
  {32'h4498dfb5, 32'hc34ccd40, 32'h43649941},
  {32'hc46a1c08, 32'h412364f7, 32'h438ded96},
  {32'h450ecdf0, 32'hc3858d24, 32'hc3013c22},
  {32'hc3830fe8, 32'h432c3ce2, 32'hc2f933df},
  {32'h44c1a129, 32'h411976da, 32'h433a304d},
  {32'hc4aa6d0b, 32'h439129fc, 32'hc12a5cf2},
  {32'h450627b8, 32'h4331da63, 32'h43d1274c},
  {32'hc4b4f5a0, 32'h44167e8a, 32'hc25f098a},
  {32'h43ae2000, 32'h4143ff1e, 32'hc2af3f7a},
  {32'hc5076938, 32'hc111d25e, 32'hc3578f4e},
  {32'h43da1a28, 32'hc308a2f9, 32'h438107d7},
  {32'hc4594f7f, 32'hc20cf4bf, 32'hc353ea84},
  {32'h449fe9a2, 32'h43850bea, 32'hc239ac16},
  {32'hc4a366c4, 32'h432cbc3d, 32'h42580552},
  {32'h4387b804, 32'hc38479b5, 32'hc34dad21},
  {32'hc49dbcc4, 32'h430781e6, 32'hbe896e74},
  {32'h44e0b567, 32'h440ef2d4, 32'hc310f4e9},
  {32'hc46c786c, 32'hc322930b, 32'hc2effa14},
  {32'h44f6ea26, 32'hc196234d, 32'h430e6363},
  {32'hc5065f6b, 32'hc27475f6, 32'hc2945c06},
  {32'h446c7182, 32'h439b263a, 32'h43ddaf04},
  {32'hc469805e, 32'hc2783e5b, 32'hc30b9896},
  {32'h44eb7be3, 32'h42ea7e49, 32'h4321af11},
  {32'hc475f924, 32'h43c7ae09, 32'hc19c04c5},
  {32'h450c00bd, 32'hc2b8507c, 32'hc33919bb},
  {32'hc511011f, 32'h432967eb, 32'hc224146d},
  {32'h44e00294, 32'hc334bd1d, 32'h42b0c623},
  {32'hc494b21b, 32'h4223fb10, 32'hc33b8838},
  {32'h441a9864, 32'h41ab2ce7, 32'h42037cc2},
  {32'hc453a3aa, 32'h43b3a5a8, 32'hc29c0c79},
  {32'h43d322a7, 32'h43a0176f, 32'h43b5ba20},
  {32'hc3b02ff0, 32'hc38477bd, 32'hc2c55a48},
  {32'h43ae7e5d, 32'hc00fa350, 32'h435312ef},
  {32'hc4fa2e6e, 32'hc39925ff, 32'hc1689e9e},
  {32'h43eadfd4, 32'hc25f0bb4, 32'h4323b3fe},
  {32'hc4389b10, 32'hc2d362c6, 32'hc27d1952},
  {32'h44aac052, 32'hc30c575a, 32'h41241c62},
  {32'hc3de8a30, 32'hc376bf2a, 32'h42d2bc60},
  {32'h44ec3126, 32'h43812b2c, 32'hc1d24388},
  {32'hc50ac155, 32'h43b37811, 32'hc257e092},
  {32'h4509c488, 32'hc32695aa, 32'hc2b59ef6},
  {32'hc485d197, 32'hc33752ac, 32'hc3502507},
  {32'h44e5fbaa, 32'hc3883f50, 32'hc39e461d},
  {32'hc4ec84f0, 32'hc082ba39, 32'hc0450345},
  {32'h44c6dfbe, 32'h43d615e0, 32'h426d87ad},
  {32'hc4bcbfde, 32'hc3bd3ad7, 32'h419fca32},
  {32'h4496155f, 32'h43a96651, 32'h41c017d3},
  {32'hc4b2359e, 32'h42f791cb, 32'hc24ea882},
  {32'hc3018cb0, 32'hc0b24adc, 32'hc38b45b0},
  {32'hc34a5c70, 32'hc2bd4762, 32'h430590f6},
  {32'h44da1b1c, 32'h42ba2fc3, 32'hc2203f17},
  {32'hc4037850, 32'hc2d527c3, 32'h43060ebe},
  {32'h4462f206, 32'h4267eedc, 32'hc3983b45},
  {32'hc481eaae, 32'hc2d6bab0, 32'h438ef926},
  {32'h4486dfc4, 32'hc1d58a02, 32'h42a42955},
  {32'hc26bbba2, 32'h42b3f265, 32'hc37dc776},
  {32'h448f33f7, 32'hc318a351, 32'hc395dff1},
  {32'hc4168f53, 32'hc3c58092, 32'h422b666e},
  {32'h45255ccd, 32'h4384ded4, 32'h40686f28},
  {32'hc45acd3d, 32'hc37488ee, 32'h42187f87},
  {32'h450faaac, 32'h43045fbc, 32'hc164f2e7},
  {32'hc4be742e, 32'h4350c1b9, 32'hc0869a25},
  {32'h451c20fc, 32'hc263d00e, 32'h42c86e30},
  {32'hc41d8cef, 32'h412e74be, 32'hc3735bc6},
  {32'h45136332, 32'h43c1537e, 32'hc3897c9b},
  {32'hc4a703d9, 32'h431661c1, 32'hc2a2407c},
  {32'h44ec7e9e, 32'hc334ca5d, 32'hc37f0de0},
  {32'hc34be740, 32'hc3232eef, 32'h42735346},
  {32'h450f98e9, 32'h43594589, 32'h438427b8},
  {32'hc3c672aa, 32'hc28d797b, 32'hc350eb92},
  {32'h43e01ec0, 32'h4374f3c4, 32'h423a90cd},
  {32'hc4e35df2, 32'h43925069, 32'h403b812b},
  {32'h44196f0c, 32'h4409641b, 32'h434a2df0},
  {32'h41afda00, 32'h415ab780, 32'h42f7b6e8},
  {32'h4416fe22, 32'hc1e3c766, 32'hc3deff98},
  {32'hc525f0cb, 32'h4310def8, 32'hc3a8234c},
  {32'h44b859be, 32'h432ded4b, 32'h43d98a39},
  {32'hc4f1855a, 32'h43eb5bc5, 32'hc2f6b8df},
  {32'hc2c88300, 32'hc3574fc2, 32'h41f413ae},
  {32'hc4f93a0b, 32'h425b2b91, 32'hc31c8942},
  {32'h44997083, 32'hc3aac29a, 32'hc0fe6520},
  {32'hc306baa0, 32'h43b346ba, 32'hc371b65f},
  {32'h447096c4, 32'h433ba6f6, 32'hc3288996},
  {32'hc40f0611, 32'hc37412a7, 32'hc2cb7f66},
  {32'h42d37930, 32'hc3801255, 32'h43034814},
  {32'hc4583854, 32'hc300c2d4, 32'h432ea67b},
  {32'h451ae7ef, 32'h43621c20, 32'h42c6b26b},
  {32'hc32d12ae, 32'hc1452ad1, 32'hc41d0ed3},
  {32'h44c46c0e, 32'h42b44193, 32'hc2998c6d},
  {32'hc4566d14, 32'h4324d9f1, 32'h422f6874},
  {32'h44e8c4bc, 32'hc2fe8f27, 32'h439a1005},
  {32'h4277c440, 32'h4321fdf2, 32'hc25277b0},
  {32'h444ed2cc, 32'h4300034e, 32'hc3a6db71},
  {32'hc476635a, 32'hc3a1226e, 32'h42673b81},
  {32'h43696c24, 32'hc30f0497, 32'hc2f484c8},
  {32'hc47b31d4, 32'h4335b4fb, 32'h4321e70f},
  {32'h4412fc74, 32'h420accfb, 32'hc3178ade},
  {32'hc3187270, 32'hc2b633a3, 32'hc31ea8c1},
  {32'h448dba33, 32'h435a49a2, 32'h42ebf4dd},
  {32'hc4234790, 32'h4123617d, 32'hc1df28d7},
  {32'h44cda561, 32'h439b61b7, 32'hc1ec5355},
  {32'hc4f97286, 32'hc3f6eba5, 32'hc1ec5534},
  {32'h432772bc, 32'hc3890561, 32'h41a4b93f},
  {32'hc4b341d7, 32'h4294b673, 32'h422e559b},
  {32'h450ac03d, 32'h425ac4f1, 32'hc291e65e},
  {32'hc477e8a8, 32'hc27967d8, 32'h4246356e},
  {32'h449c5f33, 32'h42569736, 32'hc396e250},
  {32'hc49636f5, 32'hc30b8359, 32'hc35c5db9},
  {32'h4481ecd4, 32'hc38c592f, 32'hc2b9a57f},
  {32'hc3dd23bc, 32'hc334dc8f, 32'h4324f652},
  {32'h449e32c6, 32'h435feb78, 32'hc3a871a7},
  {32'hc4f64ae9, 32'h43132233, 32'h4356b75c},
  {32'h44c57a77, 32'hc17f24d8, 32'h4301fa5a},
  {32'hc4f6b81e, 32'h4396121e, 32'h441443fa},
  {32'h44b48b92, 32'hc314352b, 32'hc41d394a},
  {32'hc50b23af, 32'hc275e7a5, 32'h4239f4dc},
  {32'h4450c95c, 32'h428537de, 32'hc3fcefd2},
  {32'hc4c2fa01, 32'hc32dbcb9, 32'h4389323a},
  {32'h44b20948, 32'h43829fd6, 32'hc375aafd},
  {32'hc4c0a3b8, 32'hc23eeedf, 32'hc2be8b88},
  {32'h4438e845, 32'hc2c4cf74, 32'hc23df2b0},
  {32'hc3dbd9d0, 32'h42ee9290, 32'hc34ab4ad},
  {32'h450465e6, 32'h42e1db26, 32'h42b4ed9a},
  {32'hc453ce88, 32'hc3da9152, 32'h429dc538},
  {32'h4397145f, 32'h433a95cc, 32'h42fd783c},
  {32'hc449a37a, 32'h43480fd6, 32'h43a022be},
  {32'h44998d4e, 32'hc2fbe839, 32'hc3e785f6},
  {32'hc4cad280, 32'h42e9fde3, 32'hc24e43e5},
  {32'h4525a54a, 32'hc14ba1d8, 32'hc2fabab7},
  {32'hc4f6de14, 32'h41a83ba2, 32'h437029e7},
  {32'h450cd7eb, 32'hc1e0f425, 32'h42e4c8a1},
  {32'hc4cc2733, 32'h4312932d, 32'h4323d937},
  {32'h44600c95, 32'h433b3681, 32'hc3b76827},
  {32'hc4dbb2ac, 32'h42c8404e, 32'hc2384702},
  {32'h4383e988, 32'h4316f73f, 32'hc2a81ca2},
  {32'hc428c5b0, 32'hc241381d, 32'h4186396d},
  {32'h44b4a282, 32'hc22516c8, 32'hc38643f6},
  {32'hc4dcbc6d, 32'hc3270418, 32'h42c7193f},
  {32'h443ce0cc, 32'h42c9549a, 32'hc2f762d8},
  {32'h433691b0, 32'hc0ebed32, 32'h4367500d},
  {32'hc4a08c3a, 32'hc0f3073c, 32'hc1155cc0},
  {32'h442d90dd, 32'hc3671eb0, 32'h42b1bda6},
  {32'hc4855bc7, 32'hc25a7570, 32'h42862d3d},
  {32'h43805d36, 32'h4455145f, 32'h414c5593},
  {32'hc3c4c288, 32'h44089499, 32'h431d9f84},
  {32'h44ea7223, 32'hc33bdd78, 32'h429f5758},
  {32'hc18073c0, 32'hc38960a0, 32'h42dd656e},
  {32'h449ec9c5, 32'hc18e77c7, 32'hc34d6cf3},
  {32'hc3d48378, 32'h4284964b, 32'hc2bf9d07},
  {32'h448a096a, 32'h437e6ce8, 32'hc38cba16},
  {32'hc4ae9b24, 32'hc1b8e285, 32'h42968a19},
  {32'h443b6b33, 32'h40b51d10, 32'hc2fe671f},
  {32'hc457bc84, 32'h431eb3f6, 32'hc38ab44a},
  {32'h44d46863, 32'hc39efefe, 32'hc2860388},
  {32'hc4dfdf97, 32'h42f4b718, 32'hc38462b3},
  {32'h44ad26a4, 32'h4372f389, 32'hc356b7db},
  {32'hc2107240, 32'h439b0663, 32'h4324044e},
  {32'h4509e504, 32'hc384aafb, 32'hc36f5736},
  {32'hc497423d, 32'hc32014f5, 32'hc36e14fc},
  {32'h44317dee, 32'h41db89cf, 32'h41d67b1e},
  {32'hc500c543, 32'h4304dbb0, 32'hc2e49b46},
  {32'h43d986f6, 32'hc38c02da, 32'hc3ea5412},
  {32'hc3889ecc, 32'hc2230e35, 32'h423de826},
  {32'h44f09f58, 32'hc281e765, 32'h41635a84},
  {32'hc4a3499e, 32'hc247a594, 32'h4357100c},
  {32'h432539f2, 32'h437aa792, 32'h41840809},
  {32'hc468935c, 32'h42e12c77, 32'h41c0c098},
  {32'h44ce4fea, 32'h4323b600, 32'hc304662a},
  {32'hc4052070, 32'h426b7692, 32'hc3b74e43},
  {32'h44ee36d0, 32'h423087e5, 32'h43ab53b7},
  {32'hc480ffa6, 32'hc3a5e58f, 32'h41fef1a5},
  {32'hc24613d0, 32'hc2281159, 32'hc1d5c174},
  {32'hc46be6ac, 32'h43d4b814, 32'h40663a14},
  {32'h444ef8f5, 32'h4271b2a1, 32'hc34a64a3},
  {32'hc3fd60c0, 32'hc388419d, 32'hc2cad67d},
  {32'h4303749e, 32'hc36a6980, 32'hc31bc6d3},
  {32'hc4970d64, 32'h4367a2b3, 32'hc39380b4},
  {32'h442c4f68, 32'h425af40f, 32'hc3088824},
  {32'hc3fa8544, 32'hc222c1db, 32'hc40510de},
  {32'h43e8eae4, 32'hc3a116aa, 32'hc34b229f},
  {32'hc4460da2, 32'hc197a9da, 32'h438c8a7f},
  {32'h44112090, 32'hc3159ef6, 32'h4301c70f},
  {32'hc473460e, 32'h432d5b45, 32'h43aa0700},
  {32'hc2c348c0, 32'h4085db48, 32'h4229c889},
  {32'hc4303b0a, 32'hc298b3c2, 32'hc37d8c30},
  {32'h45080427, 32'h4324300f, 32'hc32d0f4e},
  {32'hc50253bd, 32'hc343d45c, 32'hc2ae6b66},
  {32'h44017b90, 32'h440fd774, 32'hc248a1a7},
  {32'hc5000d99, 32'hc3056ac8, 32'hc245e6ed},
  {32'h4471ba14, 32'hc310960d, 32'h434f915e},
  {32'hc4c7a582, 32'h42b441e5, 32'h41adb8b1},
  {32'h44e31ad2, 32'hc35e04ae, 32'h42b7cf5a},
  {32'hc49fdccc, 32'h4098321c, 32'h432547c6},
  {32'h4426229c, 32'hc277735a, 32'hc2602e86},
  {32'hc4343ffc, 32'hc36f6fab, 32'hc39c3ebf},
  {32'h450bb496, 32'hc3758fbc, 32'hc38d493c},
  {32'hc4edfc59, 32'hc3710664, 32'hc3288f71},
  {32'h4434d2fe, 32'hc2923283, 32'hc366e312},
  {32'hc4e600bb, 32'h42c9772a, 32'h42bacae8},
  {32'h43a23810, 32'h431c0682, 32'hc345cd42},
  {32'hc3b74d24, 32'h425a627f, 32'h436b85e0},
  {32'h4439f97c, 32'hc3c4450f, 32'hc38fcdcf},
  {32'hc4873a6e, 32'h41891ed2, 32'h43119846},
  {32'h44cf43a2, 32'hc1f1e5cc, 32'h4244de28},
  {32'h437d8370, 32'hc3712bb2, 32'h4377981a},
  {32'h45358dc2, 32'hc10ea69d, 32'hc346c944},
  {32'hc48db2f5, 32'hc35c78be, 32'hc3163a03},
  {32'h44868437, 32'h4354f79a, 32'h42f1cf49},
  {32'hc36700fc, 32'h4298bb59, 32'h43d5c92f},
  {32'h450faeaf, 32'hc30eae38, 32'h4302ca45},
  {32'hc429ebcf, 32'h4277d255, 32'h4302d41b},
  {32'h445a4abb, 32'hc35b830f, 32'h43d7b72f},
  {32'hc4aef123, 32'h4113614b, 32'h4313e040},
  {32'h44f5216f, 32'hc2a04cad, 32'hc0bf03a6},
  {32'hc42481f4, 32'hc323fdfa, 32'h437dd83d},
  {32'h44caf4ad, 32'hc2835964, 32'hc30759f1},
  {32'hc4e63edd, 32'h421b7498, 32'hc2f8689a},
  {32'h45109866, 32'hc3014bee, 32'hc371b2c0},
  {32'hc4d38dd3, 32'hc39f1858, 32'h432c3584},
  {32'h43e927dc, 32'h4296bf35, 32'hc19149bb},
  {32'hc4ec6e4b, 32'h42fe67b6, 32'h43ac5dd7},
  {32'h438df1b8, 32'hc3b39f32, 32'h434ba524},
  {32'hc4eef75e, 32'hc36813ed, 32'h40bc8d19},
  {32'h432135b8, 32'h42c840d2, 32'h43b95149},
  {32'hc51d2da2, 32'hc31605d7, 32'h42a50c16},
  {32'h425df7c0, 32'h4392ab09, 32'h42918420},
  {32'hc4bb20fc, 32'hc2e0e2c7, 32'h435124ec},
  {32'h44a0a6f2, 32'h42251260, 32'hc13471c6},
  {32'hc3ef1c98, 32'h430eb202, 32'h408098e8},
  {32'h44d6ed30, 32'h4285487b, 32'hc422b1b1},
  {32'hc52e4caa, 32'hc26f6c15, 32'h439ba665},
  {32'h44f32468, 32'hc35e4d36, 32'hc2bdf7e7},
  {32'hc4871a56, 32'hc20afc24, 32'h4192f41f},
  {32'h444d39ca, 32'h43b632ea, 32'h43bcea93},
  {32'hc4e2bcea, 32'hc2beeda3, 32'h43ab8107},
  {32'h449d3d78, 32'hc261fe35, 32'h42fc954e},
  {32'hc4f41370, 32'h423f1ddb, 32'hc30adde0},
  {32'h436ca750, 32'hc410703d, 32'h428b701f},
  {32'hc4a73503, 32'h433c0c24, 32'h42764932},
  {32'h4508f4cd, 32'hc2159a75, 32'h437b7df6},
  {32'hc4e13df4, 32'hc093a42c, 32'hc2efc51d},
  {32'h44c41b2f, 32'h432c9b57, 32'h42a00bb5},
  {32'hc4f7ca1b, 32'hc392949d, 32'h430b8343},
  {32'h44091e4e, 32'hc2f6f287, 32'h43aefd96},
  {32'hc4cc61bc, 32'hc220636a, 32'hc35c90d0},
  {32'h44bf44d0, 32'hc31d2df8, 32'hc1c78d33},
  {32'hc4891958, 32'h43a9ef54, 32'hc1c1d614},
  {32'h44a337d1, 32'hc2cadd35, 32'hc35226ab},
  {32'hc3ecd4c3, 32'h43cfcc9a, 32'h429af816},
  {32'h440d42fc, 32'hc322fe30, 32'hc34f4227},
  {32'hc4f97cee, 32'h43989bde, 32'h4386a9f4},
  {32'h449cd77c, 32'hc307ab76, 32'hc16c65be},
  {32'hc51bf110, 32'h42cbd0cf, 32'hc330356b},
  {32'h43a967bf, 32'hc2c46785, 32'h43a6c4e2},
  {32'hc50be95d, 32'hc252c208, 32'hc205813d},
  {32'h44bdf220, 32'h4390bae1, 32'hc2376906},
  {32'hc4ef6de4, 32'h435b5414, 32'h43b75340},
  {32'h446dc39f, 32'hc39267e0, 32'hc19afbcd},
  {32'hc4691812, 32'hc39e4640, 32'h41ab5ed8},
  {32'hc2a59c98, 32'h41ea2969, 32'h42c9932a},
  {32'hc4ac7f8e, 32'h423f8376, 32'h43e1c21e},
  {32'h42f60f30, 32'h41efeb5e, 32'hc3159b02},
  {32'hc4a09996, 32'hc39b6572, 32'h42548750},
  {32'h45008f2e, 32'h4301a718, 32'h42462a66},
  {32'hc4f12c2f, 32'hc2612b0b, 32'hc2b92c53},
  {32'h443fa547, 32'h43817562, 32'h42b6c81e},
  {32'hc4347e64, 32'h4230cd6d, 32'h4401e3bc},
  {32'h44e5235e, 32'hc35ca430, 32'h43eacb61},
  {32'hc4d38d37, 32'hc291d8c0, 32'hc302c771},
  {32'h44e2f180, 32'hc3327e62, 32'h43c57fbf},
  {32'hc4d69a08, 32'hc1cf3474, 32'hc2adb361},
  {32'h4491d244, 32'h43bffac8, 32'hc311f8ca},
  {32'hc4c98569, 32'h43803d98, 32'hc33aef00},
  {32'h44c6c870, 32'hc03c60f8, 32'hc218f5c5},
  {32'hc4c311a4, 32'h42a3300c, 32'hc2870f74},
  {32'h44326b84, 32'h43bb73cb, 32'h43538874},
  {32'hc487e6b0, 32'hc3fc81e0, 32'hc2ba05fe},
  {32'h44cee14e, 32'hc31c6046, 32'hc3af3732},
  {32'hc4f1b6c4, 32'h424757f5, 32'hc3ba38b2},
  {32'h4467a691, 32'hc3621fc2, 32'hc2869a0a},
  {32'hc494dd6b, 32'h43be554e, 32'h412bc9e6},
  {32'h44c7ecbc, 32'h42aeb116, 32'hc3278400},
  {32'hc4972748, 32'hc4040299, 32'hc30cf059},
  {32'h437a35ac, 32'h4345ed04, 32'h42b4af67},
  {32'hc4fe1c5f, 32'hc3120c04, 32'hc2d3b064},
  {32'h446cd225, 32'h4332c2a2, 32'h40df331c},
  {32'hc41e1855, 32'h43206861, 32'h43294e3f},
  {32'h4463a62f, 32'hc2f152ec, 32'hc30f0a9c},
  {32'hc3d13d08, 32'hc3127dd7, 32'h429fa47f},
  {32'h447434d8, 32'hc1f598f3, 32'hc32ce1e3},
  {32'hc4f62593, 32'h42002d52, 32'h43130ffe},
  {32'h45150007, 32'hc2423f8f, 32'h43409b1a},
  {32'hc509ba36, 32'hc3c31b13, 32'hc1f39e7e},
  {32'h4503aa68, 32'h423876c6, 32'hc38319b0},
  {32'hc4e18877, 32'hc352b2b5, 32'h434768ed},
  {32'hc350b9a8, 32'hc287fdbc, 32'h43d93c62},
  {32'hc5033cd2, 32'h43df339e, 32'hc322ea09},
  {32'h43c35548, 32'h429e3386, 32'hc36909f2},
  {32'hc4a4259e, 32'hc27ca489, 32'h42b432df},
  {32'hc318dd7a, 32'hc414ccb5, 32'hc39bd761},
  {32'hc48fa673, 32'hc3b4c240, 32'h42aa8196},
  {32'h44e3c374, 32'hc2144a9c, 32'hc268e79c},
  {32'hc4bd942b, 32'hc3621062, 32'h43b9dcbc},
  {32'h43e90794, 32'hc1c4740d, 32'h4299e8d4},
  {32'hc4bb0840, 32'hc413b847, 32'h4205347d},
  {32'h44cd3fa3, 32'h435e3ee9, 32'hc39858f6},
  {32'hc501f1d6, 32'h42dd7767, 32'hc239870b},
  {32'h449409a2, 32'hc3507c41, 32'hc346e9d5},
  {32'hc4bb19ca, 32'hc30f1c56, 32'hc2c7f1cc},
  {32'h44e237e3, 32'hc1b1205e, 32'h42a67485},
  {32'hc4b02cd5, 32'h43d25e44, 32'h41743ad2},
  {32'h43280b0c, 32'hc1c7df61, 32'h43215132},
  {32'hc40487d2, 32'hc3963cde, 32'h43457585},
  {32'h4521c8be, 32'hc2a1510c, 32'h433897c7},
  {32'hc4833be3, 32'hc27ec870, 32'hc27808c8},
  {32'h44829f7e, 32'h42de0868, 32'h42c86c9f},
  {32'hc49244b2, 32'h42bae11d, 32'h42075d6d},
  {32'h44bd0b63, 32'hc33dd79d, 32'h4304de54},
  {32'hc4bf9285, 32'hc2f246ee, 32'h407ba448},
  {32'h450162b6, 32'hc30a49d3, 32'hc253bcdd},
  {32'hc360eb21, 32'hc2c8a6e0, 32'hc380e054},
  {32'h44fe262d, 32'hc1c97d30, 32'hc0b2f7a5},
  {32'hc47b0788, 32'h4363d59a, 32'hc1cc63f9},
  {32'h44d57828, 32'hc39cc9ce, 32'h42df701c},
  {32'hc3b9e826, 32'hc1cc09d8, 32'hc2f2fc90},
  {32'h4507099c, 32'hc33528c3, 32'h426e88f0},
  {32'hc3d3cbb4, 32'h42e99d2c, 32'hc3c07cc4},
  {32'h44ccd12d, 32'hc281bcdf, 32'hc38e4fcd},
  {32'hc503b986, 32'h42f1c127, 32'hc3265ce3},
  {32'h43991e08, 32'hc26183c5, 32'h42a87991},
  {32'hc398b9a2, 32'hc3af6cbb, 32'hc12c9909},
  {32'h4464e8dc, 32'h432f8dff, 32'h422d385d},
  {32'hc5028fd2, 32'h4279e1ee, 32'hc2e95db6},
  {32'h44637ada, 32'hc364489c, 32'hc2f7bb25},
  {32'hc4657318, 32'hc3a2d874, 32'h43af3699},
  {32'h44969470, 32'h43b51448, 32'h43daa351},
  {32'hc510f2c1, 32'hc2d692eb, 32'h427576e5},
  {32'h44ead953, 32'hc2a0f8c4, 32'hc3793ef1},
  {32'hc4a34772, 32'hc2b4fa60, 32'h436d8a02},
  {32'h44a3a7b2, 32'hc2a3b63f, 32'h4355a918},
  {32'hc4c25bc5, 32'hc3077b4f, 32'h4357c012},
  {32'h45026d6b, 32'hc07417e4, 32'h4210dedd},
  {32'hc44f263c, 32'h427a167f, 32'h43b3a46f},
  {32'h44e0931c, 32'hc413ff06, 32'h43da573a},
  {32'hc4f27cd2, 32'h41085092, 32'h4214596d},
  {32'h439e3f5a, 32'h43562959, 32'h433f0661},
  {32'hc5118bec, 32'h4255c38d, 32'hc3d59d59},
  {32'h4491ecd4, 32'hc3a171c3, 32'h4368fd6e},
  {32'hc40cdf66, 32'hc1549eb8, 32'h42f65c93},
  {32'h4515a863, 32'hc32fa20b, 32'hc1658f81},
  {32'hc50d5b28, 32'hc3518d92, 32'h4405c8d4},
  {32'h44ad206a, 32'h42578fce, 32'hc34ed645},
  {32'hc448ec16, 32'hc393ddc5, 32'h43c7f261},
  {32'h4461d1f0, 32'h43b5ba26, 32'h429a57c6},
  {32'hc4cb9d18, 32'h42e8bd58, 32'h43b6023a},
  {32'h44e8a070, 32'hc37eda63, 32'hc3c6d635},
  {32'hc4516096, 32'h431f3b32, 32'h423f5c0a},
  {32'h44dbc414, 32'hc24d5bf8, 32'h42a80d25},
  {32'hc498af7d, 32'hc35eb772, 32'hc3807805},
  {32'h44c76164, 32'h43977556, 32'hc28197e1},
  {32'hc4af1b75, 32'h417e8b6e, 32'h43732212},
  {32'h43979cda, 32'h41e6070d, 32'h438a4710},
  {32'hc485ea40, 32'hc3a6feb4, 32'h42bc1fb7},
  {32'h441e64da, 32'h43982bbe, 32'hc382097a},
  {32'hc43e22f6, 32'hc3b58e16, 32'hc30fdc11},
  {32'hc21954f8, 32'h43995d6a, 32'h43546dbb},
  {32'hc4847e8b, 32'h41ddaed9, 32'hc2d783e3},
  {32'h44490eaf, 32'h42e95c20, 32'h43139f20},
  {32'hc4f219b1, 32'h41893a43, 32'h41e0a343},
  {32'h4493ff22, 32'h426f8f92, 32'hc356a416},
  {32'hc4a470d4, 32'h4335aaa8, 32'hc212a4d2},
  {32'h44cd9acc, 32'hc33b0721, 32'hc26b3fbc},
  {32'hc4d31f60, 32'hc32cb363, 32'h432afdd3},
  {32'h44ef01c1, 32'h4385182d, 32'h42b73029},
  {32'hc50c5266, 32'hc3b787ed, 32'h428d8501},
  {32'h45081b20, 32'h430b9e9f, 32'h418b9d06},
  {32'hc4c7f7e2, 32'hc3c0423d, 32'h42acc8a9},
  {32'h44a76df8, 32'h42621e24, 32'hc2c41f38},
  {32'hc2128968, 32'hc34d814a, 32'h44179689},
  {32'h44db4f3b, 32'hc36de97c, 32'hc340d50e},
  {32'hc4edf33e, 32'hc2a5150f, 32'h42091bb9},
  {32'hc2c0cc54, 32'hc36b5ce0, 32'hc3aeb298},
  {32'hc47f905c, 32'h42b3fc51, 32'h425c77fd},
  {32'h44edb0c6, 32'hc3017788, 32'hc2c80daa},
  {32'hc50e0e2c, 32'hc29ce3b5, 32'h4398ba57},
  {32'h44e3c74b, 32'h43f65419, 32'hc396f1f1},
  {32'hc20931e5, 32'h4393b150, 32'hc1d10948},
  {32'h4469b47a, 32'hc253048f, 32'hc3a2fe91},
  {32'hc4eada43, 32'hc362fa72, 32'hc28c9e48},
  {32'h44b65b77, 32'h435055b3, 32'h4287d377},
  {32'hc45e35a5, 32'h43763a9b, 32'hc3a22a54},
  {32'h44b23b33, 32'hc3eb71c1, 32'h40afbef1},
  {32'hc48b2846, 32'h43811f5a, 32'hc2c144c8},
  {32'h4489a41c, 32'hc380387f, 32'hc3253138},
  {32'hc4cc1bbe, 32'h4384ea87, 32'hc35d9022},
  {32'h4498df78, 32'hc362d514, 32'hc373b044},
  {32'hc4f74d76, 32'hc2a74fe4, 32'h433e09d8},
  {32'h42946aa0, 32'hc29038a3, 32'h41ac013c},
  {32'hc445b526, 32'h439e194b, 32'h4265ab97},
  {32'h43a94ca8, 32'hc2b2348b, 32'h43e3c0f8},
  {32'hc49c6533, 32'hc28fec34, 32'h43508ea9},
  {32'h44349cc4, 32'h417b45bc, 32'hc210f7bc},
  {32'hc45958e3, 32'h42a2e9c3, 32'h434d29d9},
  {32'hc2856100, 32'h4320eec6, 32'h43bf0f1e},
  {32'hc48f8912, 32'h4109de56, 32'h42bda3c7},
  {32'h44d90998, 32'h41a52c3f, 32'hc2c2f97b},
  {32'hc41f3118, 32'h43016928, 32'h429fc2a6},
  {32'h44813112, 32'h43fe139b, 32'h43241aad},
  {32'hc2e66f90, 32'h427f61a7, 32'hc436bc9f},
  {32'h4512ac23, 32'hc278eeca, 32'hc1fe90e4},
  {32'hc4651d0e, 32'h428bc582, 32'h43a18bc5},
  {32'h44b5b231, 32'hc2a14089, 32'h4245899f},
  {32'hc4cdd200, 32'hc1f5294a, 32'h425f94b0},
  {32'h44db0824, 32'hc3835d5a, 32'h4183be74},
  {32'hc446e1c6, 32'h430f4735, 32'hc143c740},
  {32'h44d5e471, 32'hc2e45d8e, 32'h42386a4c},
  {32'hc4d54586, 32'h42ea2379, 32'h4383fad3},
  {32'h4505529f, 32'h430cea70, 32'hc30686ce},
  {32'hc4814b47, 32'hc32dc84a, 32'h436f29d7},
  {32'h4347c860, 32'h43b1db73, 32'h4297c4ca},
  {32'hc3a167b0, 32'hc31899f3, 32'h421379d3},
  {32'h44c0a210, 32'hc319e514, 32'hc22b2da9},
  {32'hc4e03e87, 32'hc2eac4c1, 32'hc2988dfe},
  {32'h450311d2, 32'h4394567d, 32'h4243234f},
  {32'hc4171ade, 32'hc20796ed, 32'h4353cc60},
  {32'h44b2a59b, 32'h42ffe91f, 32'h4395d798},
  {32'hc5102227, 32'hc1744a2e, 32'h4338f5e3},
  {32'h43ef744c, 32'hc222c4c8, 32'hc29bbf45},
  {32'hc3c3ccba, 32'h43a4b244, 32'hc2dc4046},
  {32'h42930318, 32'hc30ca934, 32'hc3e725c5},
  {32'hc3f603bc, 32'hc2f6c836, 32'hc3b4c815},
  {32'h44cb4523, 32'hc2d19075, 32'hc1aec214},
  {32'hc4016c2e, 32'h43d480d6, 32'h43418439},
  {32'h44f088d9, 32'hc158aa09, 32'hc3cfdcdc},
  {32'hc4d72c85, 32'hc3f2db46, 32'h41ca366e},
  {32'h43ec740a, 32'h43534873, 32'h43dea6b6},
  {32'hc41607bd, 32'h414383eb, 32'hc2beaf9b},
  {32'h44e232de, 32'h42f5902a, 32'hc3254c6e},
  {32'hc4ff74bc, 32'hc2d83656, 32'hc27808e6},
  {32'h442ff712, 32'h429a7a40, 32'hc2c11322},
  {32'hc3c6f5e0, 32'hc2d3198a, 32'h427b5b99},
  {32'h44b2ac48, 32'h43844170, 32'h43751aad},
  {32'hc4d5e860, 32'h436c78bd, 32'h43724fa7},
  {32'h4371f75a, 32'hc39cf368, 32'h42cc1c66},
  {32'hc4d7c299, 32'hc3036e55, 32'h42c06262},
  {32'h448c53b4, 32'h4218c3f2, 32'hc33f382f},
  {32'hc3203988, 32'hc24d962f, 32'h41a5ad52},
  {32'h45104061, 32'hc1d105f5, 32'h43dbd73f},
  {32'hc50fc803, 32'h4455c07f, 32'h42cb8e82},
  {32'h4454942b, 32'hc3824178, 32'h41f71c82},
  {32'hc50c2bf5, 32'hc14d5334, 32'h4358efc6},
  {32'h451a1784, 32'hc1ba2265, 32'hc1d84ef9},
  {32'hc4f8334a, 32'hc3668172, 32'h422c5c27},
  {32'h44ec4899, 32'hc1e82892, 32'hc2ba4c2a},
  {32'hc4304086, 32'h42808bb9, 32'h438474d3},
  {32'h44f9854f, 32'hc34b0c76, 32'h4245eed7},
  {32'hc4bec662, 32'h438dc4e3, 32'hc20f4924},
  {32'h4483e59a, 32'hc41cfeb7, 32'h4311565e},
  {32'hc50c2d6b, 32'h427ccbfc, 32'hc3f2c294},
  {32'h4508bfc1, 32'h429502d4, 32'h43a0d2e3},
  {32'hc497e54d, 32'h43c9cd97, 32'h41e945ff},
  {32'h44ac29d1, 32'h43ae980c, 32'h43293561},
  {32'hc4c860f3, 32'h42e63592, 32'h43c19a7b},
  {32'h440e35ef, 32'hc2d67889, 32'h433db786},
  {32'hc4fa32e6, 32'hc29427f0, 32'hc24ec37c},
  {32'h434bea3c, 32'hc3c617b8, 32'hc26f8a98},
  {32'hc4835f85, 32'h42b4b98a, 32'h40a7d1a2},
  {32'h442e12be, 32'hc30fd5e3, 32'h424a9bcc},
  {32'hc311ff80, 32'h41f7fbb2, 32'hc3e13ae5},
  {32'h450b90aa, 32'hc3396d43, 32'h422ee7d5},
  {32'hc4bc6d74, 32'hc172f823, 32'hc3e5abec},
  {32'h43c5f08a, 32'hc3b81dfd, 32'hc3819b3a},
  {32'hc473201c, 32'h43760dea, 32'h420f6e6b},
  {32'h4475ca80, 32'h437ef8b8, 32'hc367784f},
  {32'hc4ba7030, 32'h427861b1, 32'h4125763b},
  {32'h44c83c52, 32'h43658dc3, 32'hc3709280},
  {32'hc47890ed, 32'hc1db3f1b, 32'h438f820a},
  {32'h44c999a7, 32'hc360bb49, 32'h42f7e5c8},
  {32'hc50535c5, 32'h43908894, 32'hc3e52c32},
  {32'h4440d195, 32'h42e6e40b, 32'hc29baa44},
  {32'hc461d29e, 32'h43d2d184, 32'hc3984c9b},
  {32'h45158758, 32'h44249535, 32'hc34cd3b2},
  {32'hc4eb562f, 32'hc313da35, 32'hc26069b5},
  {32'h43b0a8e0, 32'h432a7f1e, 32'h3ff776a0},
  {32'hc50bcdc4, 32'h430b3f59, 32'h436f6fdb},
  {32'h43be79b0, 32'h431b9ab5, 32'h43a5fc70},
  {32'hc4dcd578, 32'hc2ba97d2, 32'hc2b9fa61},
  {32'h44ae8104, 32'h42fb6c8a, 32'h43501816},
  {32'hc50c76f3, 32'hc35c9153, 32'h43e40138},
  {32'h44e51ea7, 32'hc4060c9b, 32'hc337a79d},
  {32'hc4908e22, 32'hc287df88, 32'hc279d278},
  {32'h44af0edc, 32'h428076c4, 32'hc21087b5},
  {32'hc517b36c, 32'hc2ad9cb6, 32'h438b261a},
  {32'h445a8158, 32'h432cc7cf, 32'h429d91ce},
  {32'hc5020fc0, 32'h42e9669a, 32'hc2cc9a6c},
  {32'hc0fc1f40, 32'h421d5b27, 32'h431f10c3},
  {32'hc4e12bc4, 32'h43e0405e, 32'h43c78ada},
  {32'h447f2109, 32'h4394c162, 32'hc125587a},
  {32'hc4aa24e0, 32'hc330e61d, 32'h43835e10},
  {32'h4486f2f5, 32'hc32ace95, 32'hc3b9e6ce},
  {32'hc470105b, 32'hc358a5d1, 32'h43732dbb},
  {32'h452108ae, 32'h43a83829, 32'h433bb915},
  {32'hc4e86b11, 32'h43d312f6, 32'hc31e6b60},
  {32'h42a43d80, 32'hc39e38e3, 32'h40e6f7cb},
  {32'hc3d99f88, 32'h4397e36e, 32'hc3944556},
  {32'h43dd99f8, 32'h41e1d068, 32'hc2a929fd},
  {32'hc483fe3e, 32'h434c8af0, 32'h4246988c},
  {32'h4363fdee, 32'h4257d6d3, 32'h43871135},
  {32'hc4fc6250, 32'hc3af1d09, 32'h43feb7f2},
  {32'h43cf4794, 32'hc30d9de3, 32'h43cbc569},
  {32'hc2de5760, 32'h42ef2a93, 32'h42ed5a6f},
  {32'h44c7dc53, 32'hc3c5ceb3, 32'h42b4821e},
  {32'hc388cbb4, 32'h431759db, 32'hc3b75d7d},
  {32'h44878062, 32'h4372947e, 32'h435b6e50},
  {32'hc46b9bb4, 32'hc30bc50c, 32'h432d7a63},
  {32'h42235fe8, 32'hc355eb58, 32'hc2234335},
  {32'hc4a66af8, 32'hc380202c, 32'hc1f76633},
  {32'h443b5e06, 32'h4411b4ab, 32'h4367422a},
  {32'hc512a97a, 32'h42328c5e, 32'hc31b49be},
  {32'h44c66482, 32'hc0d7088d, 32'h42caf290},
  {32'hc33de75b, 32'h42932d77, 32'hc2219573},
  {32'h4506d6da, 32'hc2be4226, 32'hc400fae6},
  {32'hc4e18acb, 32'h421fd59d, 32'h428219d0},
  {32'h43908f90, 32'hc29b792d, 32'hc22101c9},
  {32'hc4290682, 32'h43c25009, 32'h42bb77d0},
  {32'hc3136992, 32'hc20e3910, 32'h41ead74a},
  {32'hc4513ffc, 32'hc3985e5f, 32'h429b557d},
  {32'h43b8605f, 32'h42ecd34e, 32'h4203bce2},
  {32'hc2aaa560, 32'h44316f5a, 32'hc3bd0411},
  {32'h4425f73a, 32'h42e51686, 32'h43f8f8af},
  {32'hc50899f5, 32'h431865e0, 32'h44003805},
  {32'h44f2d3d0, 32'h43c1ad8a, 32'hc2222d2a},
  {32'hc4b05ccc, 32'h434b9082, 32'h42818320},
  {32'h4459c57a, 32'hc304c4b3, 32'h4309742e},
  {32'hc487aca4, 32'hc2da3a40, 32'h4308c71d},
  {32'h4412b500, 32'h4252c13d, 32'hc3698de3},
  {32'hc3ec9b8c, 32'h43351fdc, 32'hc30488a3},
  {32'h43695360, 32'hc3f0f6d6, 32'hc2c7bd1d},
  {32'hc2ee5dbc, 32'hc2f04ce0, 32'hc38aaa1f},
  {32'h43a5b846, 32'hc3a011d3, 32'h4361b3f4},
  {32'h4312df0b, 32'h43046b21, 32'h4225c912},
  {32'h4503ca32, 32'hc2b853f3, 32'h42d2b88d},
  {32'hc4eb1a20, 32'hc3519ad9, 32'h442c35e8},
  {32'h451504a3, 32'h4332d916, 32'hc3333d54},
  {32'h439b8300, 32'h432a5239, 32'hc3b13026},
  {32'h438c1dcc, 32'h42f2653a, 32'h43159b0b},
  {32'hc4ac4bc7, 32'hc38e6c41, 32'hc3aa67c4},
  {32'h4502f0b1, 32'hc35ef3f1, 32'h41f56c9c},
  {32'hc5166714, 32'h43c6d555, 32'h4319b936},
  {32'h44ec7c3c, 32'h4356e1d7, 32'h4239874a},
  {32'hc39f9004, 32'h41128e7a, 32'hc13abfd4},
  {32'hc2afde78, 32'h432fc6e6, 32'h41bb13ea},
  {32'hc504b14c, 32'h43938288, 32'h430df1dc},
  {32'h4477445c, 32'h42ed8ace, 32'h43900682},
  {32'h43159062, 32'hc2978ed4, 32'h44018eeb},
  {32'h44decd1a, 32'h42ec99ea, 32'h4361a593},
  {32'hc1c7869e, 32'hc3bbbd86, 32'h4360dde8},
  {32'h4456c4a6, 32'hc27fe619, 32'h424f5f5b},
  {32'hc4b69fe1, 32'h440328ff, 32'hc349f9db},
  {32'h4493fff2, 32'hc33566a8, 32'h4416461c},
  {32'hc4bf248e, 32'h432b5251, 32'hc323a1a2},
  {32'h448238f7, 32'h4316c867, 32'h4328a00c},
  {32'hc4357348, 32'h428219a7, 32'hc2f336fb},
  {32'h44ae9e35, 32'h430eb0b6, 32'h42692860},
  {32'hc48239cd, 32'h43c0e70b, 32'hc3d1568f},
  {32'h439253ab, 32'h4365d29f, 32'hc30a97f1},
  {32'hc3b680b8, 32'h40b9f632, 32'h437e0314},
  {32'h43b3392e, 32'h430b16d3, 32'h432bf058},
  {32'hc4c79b0a, 32'hc35c6ec6, 32'hc39127f5},
  {32'h4452a342, 32'hc3b60814, 32'hc335a15e},
  {32'hc4b25336, 32'hc2a6ae2a, 32'h41af6ba6},
  {32'hc3331d6c, 32'h431f767c, 32'hc3301279},
  {32'h44e184f3, 32'h438932e8, 32'h41189534},
  {32'hc50827ee, 32'h42a59d6c, 32'hc21ccff8},
  {32'h44d22427, 32'h412f8e68, 32'h42d497c7},
  {32'hc514f633, 32'hc2abac28, 32'hc281029d},
  {32'h447fac31, 32'hc3825c32, 32'hc25998c7},
  {32'hc430377e, 32'hc40a699d, 32'hc410746c},
  {32'h444cbdfc, 32'hc1ee5979, 32'hc38119ea},
  {32'hc4d4b68d, 32'hc1971d36, 32'hc3360f2f},
  {32'h450cc509, 32'hc2d92841, 32'hc36426d4},
  {32'hc4d3f88c, 32'hc2a893e2, 32'h420019f7},
  {32'h44b86421, 32'hc32a3ec8, 32'h41d7aaed},
  {32'hc4f390bd, 32'h42b17643, 32'h42a77ec9},
  {32'h4508b1f4, 32'h43f085c9, 32'h43b18141},
  {32'hc4149929, 32'h4133f21e, 32'h43c72cfd},
  {32'h4362f130, 32'h433ff8bc, 32'hc383d998},
  {32'hc1fe9c20, 32'hc23b6cbe, 32'hc35838c0},
  {32'h438341aa, 32'h42a48968, 32'hc3513db9},
  {32'hc439b541, 32'hc303f4db, 32'hc3039a1e},
  {32'h441f4ea7, 32'h41a8c85c, 32'hc2b3c192},
  {32'hc50de664, 32'h428b0806, 32'hc0eff9a0},
  {32'h44e59f3e, 32'h42466426, 32'h42d564ad},
  {32'hc50cce71, 32'h41b5109f, 32'hc3176950},
  {32'h4482af43, 32'h438a170f, 32'h43314102},
  {32'hc4e66253, 32'hc3407531, 32'hc223e1e7},
  {32'h44c6a19c, 32'hc225c044, 32'h42164f4e},
  {32'hc5070ceb, 32'h42578967, 32'h42ffb8c4},
  {32'h44c19a6f, 32'hc3a00839, 32'h41a179ac},
  {32'hc454b2e0, 32'h4388ffb3, 32'hc4055ee8},
  {32'h44e4591a, 32'h4342fb62, 32'hc1e390ac},
  {32'hc2ebcf20, 32'hc3a55ad6, 32'hc381d362},
  {32'h440748dc, 32'h425d8094, 32'h4431b635},
  {32'hc4c84593, 32'hc391edba, 32'hc35392ee},
  {32'h4480f5ba, 32'hc315389d, 32'h423e513a},
  {32'hc3de3d64, 32'hc3b2b2ee, 32'hc352ae0c},
  {32'h44afb438, 32'hc2e3c96a, 32'h4316b922},
  {32'hc3bce938, 32'hc39630a0, 32'hc32cf999},
  {32'h439b302c, 32'hc1b512f8, 32'h439cafb3},
  {32'hc494816b, 32'hc2f6c7ef, 32'h40d2e398},
  {32'h43f9abc0, 32'hc1ab25d2, 32'h43591941},
  {32'hc2a72d98, 32'hc2e0b906, 32'hc3839f98},
  {32'h44f4ec76, 32'h43f80584, 32'h438b05fe},
  {32'hc3b75dcc, 32'hc23e9d13, 32'h43d1e948},
  {32'h451e1344, 32'h432d87f4, 32'h42dbf392},
  {32'hc34ccd99, 32'hc3797a12, 32'hc2d737a0},
  {32'h44150d68, 32'h429aa2a8, 32'h43200c88},
  {32'hc4d1d2e3, 32'h43706511, 32'hc3134972},
  {32'h45284a86, 32'h4426bec6, 32'h42aae802},
  {32'hc5035554, 32'hc2057da6, 32'hc31b64b5},
  {32'h4416751a, 32'hc215b76c, 32'h42d64a4a},
  {32'hc3b20b7a, 32'hc3650c29, 32'hc29c8d00},
  {32'h431c4c34, 32'h43c000bc, 32'h410f8df0},
  {32'hc50e561f, 32'h440c5da4, 32'hc4098ad8},
  {32'h44d21a2a, 32'hc2a71a3c, 32'h42d5ae2e},
  {32'hc45665ac, 32'h43cc743b, 32'hc3d52e31},
  {32'h446361fb, 32'h42bfdcfc, 32'hc2aa70f6},
  {32'hc46fd94e, 32'h4365c8d2, 32'hc2b79807},
  {32'h4399a424, 32'hc0347aa0, 32'hc2fcafa0},
  {32'hc418a593, 32'h4381260a, 32'h424fc7ac},
  {32'h437a7e7c, 32'h426a01f9, 32'hc3394ac0},
  {32'hc513514d, 32'h428dfee8, 32'h43820118},
  {32'h4525ef45, 32'hc3acc68c, 32'h43cec3e3},
  {32'hc457306b, 32'h43b9996d, 32'hc38545fc},
  {32'h44fd3506, 32'hc392fcca, 32'h42a9f26a},
  {32'hc4f435c3, 32'h42126d19, 32'h428d6f1e},
  {32'h450ee7dc, 32'h4398bcb7, 32'h419d54c6},
  {32'hc48413da, 32'h42b80694, 32'h42dff9c6},
  {32'h44d79a9f, 32'h400e9edc, 32'hc38db6d7},
  {32'hc42970a9, 32'h4381a2a0, 32'h426c1ca3},
  {32'h440b16d6, 32'h40cc07da, 32'hc2f7d008},
  {32'hc42ceada, 32'h44136020, 32'h42a06101},
  {32'h448d9d8f, 32'hc37ede94, 32'hc385d409},
  {32'hc2256270, 32'h435ea084, 32'hc28e28b5},
  {32'h4460c10c, 32'hc3b11dde, 32'h43751dcc},
  {32'hc4b2e41f, 32'hc361657d, 32'h434d0436},
  {32'h44b70e16, 32'h439be440, 32'h4346f066},
  {32'hc2810c50, 32'hc224b4b8, 32'hc2c691eb},
  {32'h44f01b57, 32'hc387fad9, 32'hc3cb999f},
  {32'hc3a00e3c, 32'hc2e096fd, 32'hc2f109a5},
  {32'h4508e6fe, 32'hc39aa0f7, 32'h440b13f1},
  {32'hc49aeedc, 32'hc4177bdf, 32'hc37b7425},
  {32'h443989f2, 32'hc2d16f3a, 32'hc23e0f0e},
  {32'hc4baa386, 32'h43b66683, 32'hc3cc2efb},
  {32'h445f6fc0, 32'h424902e6, 32'hc100d5fe},
  {32'hc3c4004e, 32'h43ff370f, 32'h42fa8c1b},
  {32'h442d6f52, 32'h432e27de, 32'h41c16fcd},
  {32'hc4c5c8f2, 32'h42f7f77f, 32'hc36337d3},
  {32'h43f5b548, 32'h43c5614b, 32'hc3997187},
  {32'hc48a9fc4, 32'h4287217b, 32'h42772045},
  {32'h4484c48d, 32'h42ee2e22, 32'hc37acd8d},
  {32'h42f09144, 32'hc2824a0e, 32'hc300a1ca},
  {32'h44c267d6, 32'h4188f676, 32'hc30c3d21},
  {32'hc4f829a6, 32'h42ee327f, 32'hc2f1ceae},
  {32'h43f4adfc, 32'h439ba95e, 32'hc3647336},
  {32'hc3967c2d, 32'h435850df, 32'h43b8ed3e},
  {32'hc314d2b2, 32'h42ee657e, 32'h423b0be8},
  {32'hc4f1a4a7, 32'hc3888803, 32'hc316ec2d},
  {32'h44365d41, 32'hc30a27e5, 32'hc23ec424},
  {32'hc50a611b, 32'h437aaf27, 32'hc20c14fc},
  {32'h445dfaa0, 32'hc2cd5d4e, 32'hc2887bd6},
  {32'h426503c0, 32'hc3113d3a, 32'h42c4f852},
  {32'h43f8a7f2, 32'h439980ca, 32'h4393dcfa},
  {32'hc472789e, 32'hc39448f5, 32'hc3f3acbf},
  {32'h450ce3de, 32'hc384b73a, 32'h436e9b78},
  {32'hc39b54ea, 32'h43247002, 32'hc21f640e},
  {32'h449719f6, 32'h415fc300, 32'h43d0a2f6},
  {32'hc4cc2805, 32'h43604c92, 32'hc3c0a63f},
  {32'h44d662ea, 32'hc3424249, 32'hc37a25af},
  {32'hc48ab641, 32'h42f9241d, 32'h42f78525},
  {32'h4518a5b7, 32'h41959bfb, 32'hc0ed10b8},
  {32'hc240da00, 32'h435e8b60, 32'hc28b0fc8},
  {32'h43c2e39f, 32'hc21c6fdd, 32'hc29921fe},
  {32'hc3b3ec3e, 32'h43ae4ca9, 32'hc37e3ca7},
  {32'h44cca269, 32'h43babc0a, 32'hc3480930},
  {32'hc4bf6889, 32'h43031e0a, 32'h43d5031f},
  {32'h44b34d7c, 32'h42cdb789, 32'hc3f112b4},
  {32'hc440ed04, 32'hc33144c6, 32'h43923ad8},
  {32'h45161a71, 32'hc3960729, 32'h42998a92},
  {32'hc3d1700d, 32'hc33f9ff1, 32'hc31c6143},
  {32'h450819dc, 32'h42998496, 32'h42281cc0},
  {32'hc4234880, 32'hc2aa6696, 32'h42bc4307},
  {32'h4320a418, 32'hc238fede, 32'h43e3f694},
  {32'hc4d5f4b8, 32'h437a77e4, 32'h43867ff3},
  {32'h449ccd5e, 32'h41554bb4, 32'hc3afea1e},
  {32'hc405e65a, 32'h43a03123, 32'h4389068f},
  {32'h43b6b89e, 32'hc1ed95d3, 32'h43733df9},
  {32'hc50a2210, 32'h41aefb3f, 32'h43a64676},
  {32'h450a3334, 32'h4317ad32, 32'h43b5a1b4},
  {32'hc4fde2de, 32'hc38181de, 32'h4221ec27},
  {32'hc35188b8, 32'h42816c2e, 32'hc20ab0a9},
  {32'hc4f604b6, 32'h43418a52, 32'hc39596a4},
  {32'h44aee917, 32'h4220948b, 32'h42bf97c2},
  {32'hc4a063fb, 32'h42d194dd, 32'h43d1415e},
  {32'h44cff878, 32'hc358db3e, 32'hc2535f33},
  {32'hc4efbb4d, 32'hbe7cb280, 32'hc32cd66c},
  {32'h439d5066, 32'hc209d9a4, 32'h42cfdd0c},
  {32'hc32816db, 32'h42fcc0e5, 32'hc2fdd770},
  {32'h448f6983, 32'hc3d6d9de, 32'hc371770b},
  {32'hc1bc2680, 32'hc31d1dd3, 32'h4069a228},
  {32'h44017b24, 32'hc385850e, 32'h438c893f},
  {32'hc438d7cc, 32'h42e0a744, 32'h41c4c3b7},
  {32'h43324580, 32'h41edea20, 32'hc2113387},
  {32'hc4f75b61, 32'h435f427f, 32'h43102c36},
  {32'h446f254f, 32'h42de3101, 32'h439bee81},
  {32'hc43f3f7c, 32'hc258ebf2, 32'h438313c8},
  {32'h44c959dc, 32'h42c4fd07, 32'hc452f025},
  {32'hc4deacff, 32'h431bd324, 32'h434d569c},
  {32'h44e9d044, 32'h42b94964, 32'hc3874cd8},
  {32'hc3be260e, 32'h41c8ebee, 32'hc282d68d},
  {32'h443095e2, 32'hc339d045, 32'hc3be6021},
  {32'hc4e8b20e, 32'h427201b5, 32'hc2ae7d3c},
  {32'h44addad9, 32'h43a0c014, 32'h43617a96},
  {32'hc274ba65, 32'h41300a32, 32'h41574331},
  {32'h4503c8a4, 32'hc2cd7cca, 32'hc2d770c4},
  {32'hc354140c, 32'hc33b832a, 32'hc293166a},
  {32'h42472a68, 32'hc3702316, 32'h4253fda0},
  {32'hc4b76204, 32'hc2c2e79d, 32'h425f0e94},
  {32'h44d14b15, 32'hc285ad70, 32'h3f584163},
  {32'hc46009bc, 32'hc2a2bc70, 32'hc35883d6},
  {32'h44d829fe, 32'hc30af59b, 32'h43d03fb6},
  {32'hc4a95ab4, 32'h428ae6dc, 32'hc1b80e03},
  {32'h44f8c104, 32'h4281dc8e, 32'hc1249736},
  {32'hc3031c29, 32'hc1a9bbb4, 32'h41df8ef4},
  {32'h445595aa, 32'h43a10c63, 32'hc34ff9a4},
  {32'hc4b43d9b, 32'hc39753b7, 32'h4167375a},
  {32'h42a1e58c, 32'hc1cb237c, 32'hc24eddaf},
  {32'hc46a3c57, 32'hc27abda8, 32'h432e065c},
  {32'h43296ae6, 32'h43a878d4, 32'hc1e2300b},
  {32'hc4f4a32b, 32'h42d15144, 32'hc2867253},
  {32'h44760888, 32'hc407072b, 32'h412c8d02},
  {32'hc50595fc, 32'hc3c7e3ce, 32'h420e5fe8},
  {32'h448d2fd9, 32'h42ef59e3, 32'hc39d2565},
  {32'hc5105fec, 32'hc1eb7e75, 32'h432b1b79},
  {32'h44f2f0c6, 32'h4219f895, 32'hc31e51ba},
  {32'hc3e29259, 32'h42cf4239, 32'hc2c9a9e3},
  {32'h43c496a4, 32'h43732706, 32'hc1c3ebf0},
  {32'hc4916910, 32'h42eb3cb0, 32'hc3824e20},
  {32'h45027d9d, 32'hc31d2141, 32'hc24e82b3},
  {32'hc4d447a8, 32'h422c20ee, 32'h4204efcc},
  {32'h44bfa859, 32'h42c8b7b8, 32'h43ae8df5},
  {32'hc4bb5c89, 32'hc3901a8e, 32'h40a9fcd2},
  {32'h4490175c, 32'hc31ad4b3, 32'h4317e107},
  {32'hc28eae12, 32'h41fd30e1, 32'hc3b643dc},
  {32'h44235c73, 32'h4364093b, 32'h43ad6ec0},
  {32'hc497eef2, 32'h43868d9a, 32'h4305a241},
  {32'h45008e0f, 32'hc34ce8d9, 32'h43841d3a},
  {32'hc47695d6, 32'h43cf154a, 32'hc27e1e6f},
  {32'h449588ff, 32'h42c4b2d4, 32'hbfcb4050},
  {32'hc439f3e1, 32'hc38733e5, 32'h433da7e6},
  {32'h44d610a4, 32'hc388989c, 32'hc37d5fec},
  {32'hc4a9016e, 32'h4312af62, 32'hc3328131},
  {32'h44b2d849, 32'hc31a6efe, 32'h42d84561},
  {32'hc50427e4, 32'h437fe780, 32'h4331855d},
  {32'h44c884a6, 32'h431b0575, 32'h430f55a9},
  {32'hc4ac6baa, 32'h42404046, 32'hc25aa0b9},
  {32'h44eeaf38, 32'h402a12c8, 32'hc2c187f4},
  {32'hc4b4c82e, 32'h437094d7, 32'h43957a9b},
  {32'h44dc704a, 32'hc2d6b2d4, 32'hc35dbfc5},
  {32'hc508e0f6, 32'h42da18e7, 32'h429b0c85},
  {32'hc1f49ad0, 32'h4370c13a, 32'hc34ce8d2},
  {32'hc4f6deff, 32'h426d2bab, 32'hc39ac498},
  {32'h4503d63c, 32'h43b28709, 32'h42426f05},
  {32'hc4ed8b28, 32'h432cc07d, 32'hc3c07555},
  {32'h44c86684, 32'h43133ec6, 32'h436ec575},
  {32'hc4938d58, 32'h43c8638d, 32'h4400e8c1},
  {32'h450170c7, 32'hc1998c7d, 32'hc2e02cb9},
  {32'h42cdd160, 32'hc3b64bba, 32'h424c8c9b},
  {32'h440d8d48, 32'hc3171983, 32'hc3029ea1},
  {32'hc3bcb527, 32'hc2bcdabf, 32'hc34e44d8},
  {32'h451bbb30, 32'hc358adcd, 32'hc3a15599},
  {32'hc506412b, 32'h42adf2de, 32'h4321d566},
  {32'h445b465d, 32'hc402fc5c, 32'hc3920112},
  {32'hc5079032, 32'hc3c0066b, 32'hc324db44},
  {32'h44ae20a1, 32'h41cb9997, 32'h410d6128},
  {32'hc4f768f7, 32'h42fdddcf, 32'h41911673},
  {32'h44ca1eba, 32'hc38df919, 32'hc3264fde},
  {32'hc4b0e718, 32'hc28d04d4, 32'hc419d9bb},
  {32'hc39346c0, 32'h41d06479, 32'h42d26f8d},
  {32'hc3fa4b7c, 32'h429acf00, 32'hc28b7db6},
  {32'h43d006a0, 32'h43c09f71, 32'hc299ec62},
  {32'hc4f441d5, 32'h42d09574, 32'hc38651d2},
  {32'h44f46f52, 32'hc2b21e4d, 32'hc24e8412},
  {32'hc45be1de, 32'h42c87f66, 32'h43abbe7f},
  {32'h4505d19b, 32'hc2563b06, 32'hbe781e80},
  {32'hc4b9ebe1, 32'hc250a4c2, 32'h420112a7},
  {32'h4506bd9f, 32'hc3574649, 32'hc2a0d2c5},
  {32'hc47ef210, 32'h4363b8fe, 32'hc276993e},
  {32'h43cc44fe, 32'h42e60653, 32'hc27a214f},
  {32'hc494c830, 32'hc37a5a41, 32'h43900e1d},
  {32'h422f4270, 32'hc383fe38, 32'hc3419427},
  {32'hc42b2f54, 32'h436a3443, 32'hc370a3b4},
  {32'h44c9b8f8, 32'h41c8c995, 32'hc264909e},
  {32'hc424c098, 32'h43e56bb3, 32'h43d6c240},
  {32'h4500516a, 32'hc3848980, 32'h43b33229},
  {32'h4389ca33, 32'h43975907, 32'h42d4ecc8},
  {32'h44d2a489, 32'hc2b52d87, 32'hbff4059a},
  {32'hc50e51e6, 32'hc3e2d2fc, 32'hc2432854},
  {32'h44669d2a, 32'hc3ae931c, 32'hc38081e3},
  {32'hc509970b, 32'h431d81ec, 32'hc2781f41},
  {32'h44824aca, 32'hc146cf14, 32'h4358e058},
  {32'hc42b2195, 32'hc36404ee, 32'hc2f224dc},
  {32'h44042cb8, 32'h41249f16, 32'hc1ccf0e3},
  {32'hc51230fe, 32'h432e3a53, 32'hc1062c46},
  {32'h44b7976d, 32'hc2e28521, 32'hc35a62ac},
  {32'hc432d6a7, 32'h42f45e04, 32'h43134529},
  {32'h44c63808, 32'h42e863d3, 32'h42f46d68},
  {32'hc43a0594, 32'h438ef718, 32'hc1dd64e7},
  {32'h44c6f3b4, 32'h42b52956, 32'hc2204386},
  {32'hc4f540b6, 32'h422782ef, 32'hc27c08f6},
  {32'h4500d494, 32'hc19893fc, 32'hc38f9bc6},
  {32'hc4c4f6e1, 32'h43cea7eb, 32'hc27258b8},
  {32'h43a0976e, 32'hc3a31262, 32'hc3944a1c},
  {32'hc429af30, 32'hc3e07d9e, 32'h434d4724},
  {32'h44509d40, 32'hc28bfb70, 32'hc3b942d7},
  {32'hc4df101b, 32'hc2cc772e, 32'hc3da21b3},
  {32'h44b526d2, 32'h42e01143, 32'h431003aa},
  {32'hc4f7075a, 32'h4290044d, 32'hc3b69b14},
  {32'h42cb94d0, 32'h438351e8, 32'h431ed98d},
  {32'hc4ba5464, 32'h43a355c0, 32'h435f5436},
  {32'h435a13dc, 32'h4239820f, 32'h42da1e8f},
  {32'hc468d464, 32'hc22370e4, 32'hc26af313},
  {32'h44e8c7fc, 32'hc401d1ee, 32'h43871d4c},
  {32'hc418431c, 32'h439c9d77, 32'h43c8356c},
  {32'h44755ca1, 32'hc2233163, 32'hc2a7508d},
  {32'hc49dc138, 32'h43164852, 32'hc39ba03f},
  {32'h4394b8a2, 32'hc2aba3de, 32'hc2b42044},
  {32'hc4833a8d, 32'hc29dc28c, 32'hc3228a30},
  {32'h450a9df6, 32'h4229bdc9, 32'h422e2e01},
  {32'hc5139183, 32'h4380f806, 32'hc389897d},
  {32'h45112f55, 32'hc353ceb0, 32'h4328c5b9},
  {32'hc4a0ea17, 32'hc348bff7, 32'hc06a722c},
  {32'h450b8d33, 32'hc379bc3c, 32'h41d341dc},
  {32'hc50d532a, 32'hc33c0df1, 32'hc318b08a},
  {32'h445dbf6c, 32'h438c952d, 32'h421eda6f},
  {32'hc4fda102, 32'hc10c9651, 32'h41c5ba69},
  {32'h443a07fe, 32'hc39f320d, 32'h420fc8c9},
  {32'hc38ba0a0, 32'h421976e8, 32'hc334cb03},
  {32'h4468b3b0, 32'h43612fc5, 32'hc36f7f7e},
  {32'hc4c05e4e, 32'h433d1728, 32'hc40c74f6},
  {32'h44dc959d, 32'h41e8dcce, 32'h41b446aa},
  {32'hc4f55b7b, 32'h43629f90, 32'h43c7bdf9},
  {32'h44fe15d3, 32'h42ccf0d2, 32'hc38cddf1},
  {32'hc4349723, 32'h42f10b8f, 32'h435c78bb},
  {32'h43ac335f, 32'hc3d568d1, 32'hc2ad306c},
  {32'hc4891b22, 32'h4337aef9, 32'hc32c47a0},
  {32'h44180b58, 32'hc2a7e94c, 32'h4400e07d},
  {32'hc4f77ceb, 32'hc2d27f08, 32'h43c636aa},
  {32'h44cfcc2a, 32'hc19a0b68, 32'h43379f82},
  {32'hc49f677c, 32'h42a7520d, 32'h42309949},
  {32'h445f9f6d, 32'h42f89a65, 32'hc2654052},
  {32'hc33a5d4e, 32'hc3530021, 32'h421230da},
  {32'h44029604, 32'h42bf3476, 32'h4182bc22},
  {32'hc4a27e14, 32'hc3185f76, 32'h42a751c4},
  {32'h45144f48, 32'hc3b27750, 32'h43990bd5},
  {32'hc4d8b731, 32'hc28dbb9e, 32'h4332a622},
  {32'h4468484b, 32'hc3ee8562, 32'hc3bd86e1},
  {32'hc519ef87, 32'h43c7dd50, 32'hc22dd2ee},
  {32'h44fb110d, 32'h4286b9ef, 32'hc345e518},
  {32'hc5078208, 32'hc295204e, 32'hc23fd485},
  {32'h44eee3fb, 32'hc399a579, 32'h44015da1},
  {32'hc2bb819f, 32'h430879ab, 32'hc2ea86e2},
  {32'h447927ba, 32'hc35b0041, 32'hc2a40582},
  {32'hc4d69c12, 32'h43a5a478, 32'h438f0e8e},
  {32'h44ad9b70, 32'h41aaa5c0, 32'hc35a8c73},
  {32'hc5293880, 32'hc38da636, 32'hc289d8f5},
  {32'h44e1e86a, 32'hc3b74875, 32'h42a1f8de},
  {32'hc43e6ad1, 32'hc30352ae, 32'hc395cee6},
  {32'h44a3831f, 32'hc31417c0, 32'h4304bf50},
  {32'hc4f0bb6a, 32'h4277ec0e, 32'h43342779},
  {32'h44f4abd0, 32'h418138e4, 32'h4316da1b},
  {32'hc407c320, 32'hc3c3167e, 32'h43a509d3},
  {32'h4453371c, 32'h427a993e, 32'hc2989341},
  {32'hc3b446f4, 32'h42c2857b, 32'h43a44969},
  {32'h44ce2906, 32'h4363795c, 32'hc1e0e8f3},
  {32'hc23c6546, 32'hc30c69bc, 32'hc3bc5006},
  {32'h44bf47f0, 32'h430051c9, 32'h43161856},
  {32'hc50e58ce, 32'hc395296b, 32'hc3348ea8},
  {32'h432a85a6, 32'hc33021d3, 32'hc2b5c47b},
  {32'hc3f9ced8, 32'h43aae8de, 32'hc3b59ba2},
  {32'h44ff9458, 32'h42406011, 32'hc33d2a9c},
  {32'hc4a2e47d, 32'h42447171, 32'hc3277b50},
  {32'h449153d4, 32'h43dba3b4, 32'h43434f74},
  {32'hc49adb36, 32'hc227c3ab, 32'hc2ea9e59},
  {32'h45021929, 32'hc0eba400, 32'h411177bc},
  {32'hc3180de0, 32'h436003be, 32'h4312b3e9},
  {32'h44f29cfb, 32'h42de6a47, 32'h43b57771},
  {32'hc37f637a, 32'h43747841, 32'hc204d647},
  {32'h450a3eb8, 32'hc2993127, 32'hc33550a2},
  {32'hc508d614, 32'h42b1dd49, 32'hc267a1ec},
  {32'h447b3907, 32'h4323bf4c, 32'h431f4b2d},
  {32'hc41b7efa, 32'hc3029feb, 32'hc34273c0},
  {32'h433ff710, 32'hc31a6e9e, 32'h4344f6ef},
  {32'hc4940c5a, 32'h441b6a5b, 32'h429ef6b0},
  {32'h42ad7c8c, 32'h43d77f9e, 32'hc4051e95},
  {32'hc44ad968, 32'h41b6dc72, 32'hc43dd661},
  {32'h432c5d79, 32'hc3836609, 32'h4197500a},
  {32'hc50635a1, 32'hc2ddf8a7, 32'hc41ac4cf},
  {32'h43f302c0, 32'hc3355a13, 32'hc36ade03},
  {32'hc50ac1ef, 32'hc326c771, 32'h43004419},
  {32'h44bb9c19, 32'h43bac7f0, 32'h4332063e},
  {32'hc33cb2e0, 32'h4301471f, 32'hc3cd8f07},
  {32'h448f666f, 32'hc38c5461, 32'hc18e9975},
  {32'hc4236e2c, 32'h421b94c3, 32'h4295afa7},
  {32'h44d9a58c, 32'h4321ab1a, 32'hc38a133a},
  {32'hc388eafa, 32'hc324be96, 32'h42a00b05},
  {32'h451a04b8, 32'hc2e63218, 32'hc3ce1177},
  {32'hc3f056d8, 32'hc3d0f882, 32'h41962f7a},
  {32'h44d510d6, 32'hc3a06c5c, 32'hc38987d7},
  {32'hc4645bcf, 32'hc13b5378, 32'hc2e80552},
  {32'h44f5d728, 32'hc29e1d53, 32'hc2dc7980},
  {32'h42027a62, 32'h434405e6, 32'h43d18539},
  {32'h42d0d3ee, 32'h4216cdfd, 32'hc2a24c21},
  {32'hc5126992, 32'h43a9f9bf, 32'hc284f6e0},
  {32'h4466f556, 32'h41c9f61b, 32'h43d3d09a},
  {32'hc38569f2, 32'h42d986fe, 32'h44502675},
  {32'h44301245, 32'hc35ed345, 32'hc1f33fe5},
  {32'hc4f3049a, 32'h42f334da, 32'hc384cd00},
  {32'h43d07951, 32'hc2f51d13, 32'hc36ae16c},
  {32'hc3b408c5, 32'h42c8934b, 32'h4334284d},
  {32'h44a310f0, 32'hc384a2de, 32'h4382ac77},
  {32'hc5015955, 32'h430ffc17, 32'h42f43b06},
  {32'h44c7e90b, 32'h437f7833, 32'hc29b6c9a},
  {32'hc4e92de2, 32'h435c270c, 32'h40e7ecfb},
  {32'h4447ae20, 32'h410697dc, 32'h441bb8ec},
  {32'hc45b6749, 32'hc38109d6, 32'h42aa8ae9},
  {32'h44a51363, 32'h41983443, 32'hc32f2be4},
  {32'h4254989d, 32'hc300d389, 32'hc4043568},
  {32'h4478e825, 32'hc128ef1a, 32'hc3fd7f3e},
  {32'hc430f321, 32'hc34edf48, 32'h43409d5f},
  {32'h44d5d950, 32'hc1a27ec1, 32'h42c9f787},
  {32'hc4863b74, 32'h430d1a19, 32'h42fe9b42},
  {32'h44e92bf7, 32'h42eab32c, 32'h4307d4f9},
  {32'hc4fa2753, 32'hc2c60365, 32'hc3d8cd68},
  {32'h444ba1db, 32'hc294bfbe, 32'hc0b0804f},
  {32'hc3875be0, 32'h42999ef6, 32'hc315b58d},
  {32'h45279c96, 32'h43909c91, 32'hc3475098},
  {32'hc3b030c0, 32'hc28c5570, 32'hc33d9df5},
  {32'h44278c78, 32'h43ee66fc, 32'hc3027737},
  {32'hc5041422, 32'h42519b97, 32'hc324bc78},
  {32'hc32afb38, 32'h43f83c21, 32'hc3433f69},
  {32'hc44ed97c, 32'h413b979e, 32'h41c67efe},
  {32'h44fa3560, 32'hc2044052, 32'hc305f194},
  {32'hc506397f, 32'hc2d7db14, 32'h42059bbb},
  {32'h4488af5d, 32'hc30e3c06, 32'hc22981fe},
  {32'hc46a2fba, 32'h42f9ac74, 32'hc3449cfd},
  {32'h44b84e42, 32'hc413ae2b, 32'h43df2b0f},
  {32'hc4d3390b, 32'h43e5ffa0, 32'hc1d33c2c},
  {32'h4390c97c, 32'hc3651af9, 32'hc206b3ac},
  {32'hc4f61946, 32'h440f27f4, 32'hc3a30796},
  {32'h446339e8, 32'h4230d7ed, 32'h43439f31},
  {32'hc3d1e138, 32'h422d5de6, 32'h40787400},
  {32'h4482707f, 32'hc25b3f11, 32'h41639a0b},
  {32'hc3d97b78, 32'hc227b4cf, 32'h42909dfb},
  {32'h44454fb8, 32'hc14cf47a, 32'hc351dcf4},
  {32'hc4d29922, 32'h427e7adf, 32'h417ad9b8},
  {32'h44a5b5de, 32'h4373502b, 32'h43326b7a},
  {32'hc295cea0, 32'hc29f4125, 32'hc2b952a8},
  {32'h44c8d2be, 32'h43ad9ec4, 32'hc3a4734c},
  {32'hc3d2632c, 32'h42ae6a84, 32'h439d31f0},
  {32'h44c06132, 32'h437297bf, 32'hc366aea7},
  {32'hc49f9780, 32'h4320edea, 32'h4286108d},
  {32'h44b7a947, 32'hc2a49f04, 32'hc38830a7},
  {32'hc3194530, 32'hc2f3860e, 32'h442217d2},
  {32'h44c17ec4, 32'h3fce8e1c, 32'hc21d42e6},
  {32'hc4cc568a, 32'h41865d3a, 32'hc279b588},
  {32'h448e6602, 32'hc2de0a55, 32'hc239e216},
  {32'hc4c25144, 32'h436a1afb, 32'hc3a3e606},
  {32'h44423f6a, 32'hc32e169f, 32'hc2b0f066},
  {32'hc48c9ccc, 32'h43245d51, 32'h435a7443},
  {32'h44b92750, 32'h43511a8f, 32'hc30aa9cf},
  {32'hc43546fa, 32'h4291152a, 32'h4308219a},
  {32'h447145c0, 32'hc10be1c8, 32'h4405dc26},
  {32'hc4f4651e, 32'hc2d0f9fa, 32'hc27cf00c},
  {32'h450e67b3, 32'hc2e49f73, 32'hc2891870},
  {32'hc513859c, 32'hc384c62f, 32'hc34619b5},
  {32'h43703970, 32'h4319020c, 32'h4312b36c},
  {32'hc40d9304, 32'hc36d9245, 32'h43c1526c},
  {32'h44839ac4, 32'hc350eff4, 32'h41c04b6e},
  {32'hc3072a50, 32'hc3493718, 32'h425eb349},
  {32'h44dc65b9, 32'hc2f89149, 32'hc2b6997e},
  {32'hc38c0ba6, 32'h432d4562, 32'h430fcf43},
  {32'h4452ff5c, 32'h43045b5f, 32'h41446dc1},
  {32'hc4c03078, 32'hc39adf4e, 32'h438b8d68},
  {32'h44a6e719, 32'h436669fc, 32'hc3265938},
  {32'hc43776d0, 32'h4305ddf7, 32'h42f21d3c},
  {32'h44ff1f50, 32'hc33dd635, 32'hc375c551},
  {32'hc3c2edae, 32'h435f755e, 32'h422f20f0},
  {32'h4379d4bb, 32'h42248e0b, 32'hc31b6635},
  {32'hc5007e68, 32'hc347559e, 32'h4321648a},
  {32'h43e2f0c4, 32'hc32d2b94, 32'hc2383d50},
  {32'hc4d6f541, 32'hc3269cde, 32'hc3194b8a},
  {32'h447ffdde, 32'hc3356b1e, 32'hc3190a87},
  {32'h44f39abf, 32'h41788a5e, 32'hbe976285},
  {32'hc4284498, 32'hc409e12c, 32'h421b6089},
  {32'h4449539c, 32'h43f2e37e, 32'hc35f70c5},
  {32'hc4fd3938, 32'h428e559f, 32'h4409a158},
  {32'h4424528d, 32'hc3361be7, 32'hc30b0781},
  {32'hc4f498f1, 32'h427dc558, 32'h437fde7d},
  {32'h441b9abe, 32'hc2cc0549, 32'h417bb8d8},
  {32'hc4d823b9, 32'hc2ef1fab, 32'hc2adedd7},
  {32'h4431381c, 32'hc145a86e, 32'hc2aa267e},
  {32'hc519a96c, 32'h436dc212, 32'h43a41a49},
  {32'h444d16d4, 32'hc3a97901, 32'hc2b40055},
  {32'hc435e2b1, 32'hc24f2c3a, 32'h43336c73},
  {32'h450d2ac3, 32'h43478522, 32'h43af52de},
  {32'hc4427dd9, 32'hc37a640f, 32'hc3908dcc},
  {32'h442809d0, 32'h43869a43, 32'hc188b266},
  {32'hc518d62c, 32'h421724cf, 32'h4332a8ce},
  {32'hbfedf880, 32'hc218098e, 32'hc19050d4},
  {32'hc4b8a4f4, 32'hc3ac2400, 32'hc203cb10},
  {32'h43a3d5d5, 32'h4259dd30, 32'hc34854e2},
  {32'hc4106d8c, 32'h43a27ff2, 32'h43d5c7c8},
  {32'h45021234, 32'h41f2ebd9, 32'hc3585252},
  {32'hc4c90555, 32'h4133c166, 32'h43c03ea8},
  {32'h44762e4c, 32'hc20f38ec, 32'hc2bbf0e1},
  {32'hc39704dd, 32'hc3f43c13, 32'h42d3854b},
  {32'h433e18d0, 32'hc2c5ba2a, 32'hc3b50181},
  {32'hc500ab4c, 32'h433b97e7, 32'h4283fba9},
  {32'h45022fb0, 32'hc3d2aa23, 32'hc413ed3f},
  {32'hc518fdbe, 32'hc3ee0df3, 32'hc33e7316},
  {32'h451af0cd, 32'h440c6c86, 32'h42c2f71b},
  {32'hc4c51b9a, 32'hc2db2c7f, 32'h438918e0},
  {32'h43c0540e, 32'hc2ff246b, 32'hc22717dd},
  {32'hc4d4128a, 32'h42b3006b, 32'hc2adda44},
  {32'h44daabfe, 32'hc2e17296, 32'h44121b7e},
  {32'hc4a111ea, 32'hc27e46ea, 32'hc1c7b0ae},
  {32'h443b3692, 32'h42879a3d, 32'hc29e4d97},
  {32'hc51215d9, 32'hc1cd79bb, 32'h42e3b350},
  {32'h44f1211c, 32'hc27cec46, 32'h4318d690},
  {32'hc4b20a8c, 32'hc3925fe5, 32'h434428ea},
  {32'h44ff074c, 32'h42d738da, 32'h42aaad7b},
  {32'h43ee8673, 32'h42fd508e, 32'h43ae04bf},
  {32'h44f01888, 32'h42b222cd, 32'h43353677},
  {32'hc4c484c8, 32'h433bc0a4, 32'hc3c6eddc},
  {32'h431f4778, 32'h439d2574, 32'h43110b9c},
  {32'hc47347a5, 32'h42da4a55, 32'hc31f1b3b},
  {32'h4525dd89, 32'hc201235a, 32'hc0ced753},
  {32'hc4b1403e, 32'hc27adc77, 32'h41c1e9c8},
  {32'h450fc0a0, 32'h4284f7df, 32'h427bd8a0},
  {32'hc516cd22, 32'hc279650e, 32'hc2e63f32},
  {32'h442d38c0, 32'hc0af19fc, 32'h4376e853},
  {32'hc43b2bef, 32'h423b6d03, 32'h42e3c313},
  {32'h4418109a, 32'hc3d0ff12, 32'h4316cd05},
  {32'hc48d3f86, 32'h441745f0, 32'hc3d19e2c},
  {32'h450ef406, 32'hc32b8b2c, 32'h3ff38b40},
  {32'hc4be9a1a, 32'hc308fcd3, 32'h43170ae6},
  {32'h44a34a4f, 32'hc26065c2, 32'hc2e26362},
  {32'hc4b43d15, 32'h4300e50e, 32'hc388b42d},
  {32'h44556a36, 32'h42b8c9dc, 32'h43c71d44},
  {32'hc4ccb910, 32'hc2f08afd, 32'hc24ee792},
  {32'h4481fa2d, 32'h43ae1ce4, 32'hc27208d2},
  {32'hc423120e, 32'h4178f354, 32'hc2803ea9},
  {32'h44e409ce, 32'h42ed00ec, 32'h42e390be},
  {32'hc336daea, 32'hc3ad03ef, 32'hc2a4c089},
  {32'h44f8235c, 32'h41918aa9, 32'hc303a71f},
  {32'hc3d8d40e, 32'hc32f3fee, 32'h42dbc545},
  {32'h451058bf, 32'h4346a16f, 32'h42c4f0a1},
  {32'hc474c47a, 32'hc2c54f91, 32'hc28dbc38},
  {32'h44347e4c, 32'h4327a608, 32'hc3b76f12},
  {32'hc38e780e, 32'hc3bba773, 32'hc334fbb3},
  {32'h44f1bbb6, 32'hc41f1999, 32'hc23a890f},
  {32'hc4cc8d78, 32'hc3ee9568, 32'hc38a7b36},
  {32'h45052c8e, 32'hc332c805, 32'hc31ec0df},
  {32'hc4197451, 32'hc36dda27, 32'hc210439a},
  {32'h444c6b4b, 32'h43c7d636, 32'h43b28b72},
  {32'hc4902997, 32'h4386a624, 32'h43b84888},
  {32'h445aac98, 32'hc2684fee, 32'h43576d27},
  {32'hc4a92c1d, 32'h4381747d, 32'hc3a5a121},
  {32'h4520b9e9, 32'h42cf105c, 32'hc40522c6},
  {32'hc4e15f62, 32'hc2ce8ff1, 32'hc390fc45},
  {32'h431bf9a8, 32'hc3998405, 32'h43514983},
  {32'hc51365f4, 32'hc397dd67, 32'h4285fe4b},
  {32'h45030a5e, 32'hc2a9ef2c, 32'h42cd423f},
  {32'hc50e868b, 32'h434ebb41, 32'hc34597ee},
  {32'h43dcd0bb, 32'h434069ea, 32'hc35cd562},
  {32'hc449b12b, 32'hc2b65d81, 32'hc3aa3e55},
  {32'h44cfb324, 32'hc3464a58, 32'hc2a6db4d},
  {32'hc333c1a9, 32'hc1d47c8d, 32'h4298cd66},
  {32'h44e4a25c, 32'h43285dbc, 32'hc429859d},
  {32'hc50a3fba, 32'hc1b9065d, 32'hc3d6e30e},
  {32'hc1f02020, 32'hc1e2f077, 32'hc2d3eddf},
  {32'hc4bc2bf5, 32'hc35aeadb, 32'h43298d1e},
  {32'h44baed91, 32'h43a640d8, 32'hc33b02a0},
  {32'hc4b94558, 32'h431ba18c, 32'h4304f9a8},
  {32'h4431dc28, 32'h43bc0615, 32'hc2be7388},
  {32'hc4238fe6, 32'h435f413f, 32'hc1ac67a2},
  {32'h44fd63cd, 32'h4315c8c7, 32'hc38f8ad2},
  {32'hc4c2a7a5, 32'hc31f5640, 32'h43bbf5c9},
  {32'h44f2d0da, 32'hc351a287, 32'h429f88d8},
  {32'hc4392faf, 32'h432a6e7f, 32'h4334e363},
  {32'h44e66d02, 32'hc428944f, 32'hc26d3da1},
  {32'hc3a44ef0, 32'hc2ebb310, 32'h4334a2c3},
  {32'h43a6d408, 32'h4306097f, 32'hc1fff741},
  {32'hc43e6aa8, 32'h42f34662, 32'h44260450},
  {32'h447f21da, 32'h432431b4, 32'hc263b046},
  {32'hc4c94ee7, 32'hc365b486, 32'h420cacd8},
  {32'h4411cad2, 32'h4324a5ee, 32'h41b44ad1},
  {32'hc4199544, 32'hc24ce43a, 32'h4202e6e6},
  {32'h44555c0e, 32'h43280acc, 32'hc397e02f},
  {32'hc496a750, 32'h42a77105, 32'h42c2e30a},
  {32'h43c4d898, 32'h437a91c8, 32'hc29060a1},
  {32'hc4b82006, 32'hc2ccd5db, 32'h432b2ad8},
  {32'h438b00c9, 32'h423efc1a, 32'h426d23f4},
  {32'hc24b0345, 32'h43a9c118, 32'h43516d3a},
  {32'h44e32062, 32'h42ae8d53, 32'h42b80cf2},
  {32'hc4ddc6b5, 32'h42dcc885, 32'h433d0ffe},
  {32'h44b9b3ba, 32'hc397019a, 32'h42bcd51e},
  {32'hc4abfa60, 32'hc3143312, 32'h433cbbe9},
  {32'h44f31c06, 32'hc3859782, 32'hc3807aaa},
  {32'hc4771425, 32'hc24c4d1e, 32'h409dbe64},
  {32'h44cce6c2, 32'h438b0d48, 32'hc3a84877},
  {32'hc4cdb8df, 32'h4248f6bc, 32'h43122555},
  {32'h443eb6cf, 32'hc240b205, 32'h428cb76d},
  {32'hc48f1461, 32'hc3dbc7a1, 32'h42f0df37},
  {32'h44aad75c, 32'h435d2115, 32'h4320817b},
  {32'hc4b06c10, 32'hc3ca6ebd, 32'hc2c4c157},
  {32'h44df23f2, 32'hc152db61, 32'hc39acf08},
  {32'hc3a1b440, 32'hc37dc6b8, 32'hc38240c2},
  {32'h4474a3bb, 32'h420a928c, 32'h42aa3db0},
  {32'hc476670a, 32'h431c3456, 32'hc32ac8ba},
  {32'h446d10f5, 32'h432a2afd, 32'hc3daa9f5},
  {32'hc40085b8, 32'h43b950f0, 32'h432cda37},
  {32'h443d2723, 32'h43e211dd, 32'h43ffb99d},
  {32'hc33875bc, 32'h42cf1715, 32'h43a97b62},
  {32'h44812001, 32'hc2e83994, 32'h43dd1793},
  {32'hc44480d3, 32'hc2f4e2c5, 32'hc30a554e},
  {32'h44fb0a2d, 32'hc27cd14e, 32'hc2d0d6d4},
  {32'hc5086222, 32'hc3839e6d, 32'h42f5d426},
  {32'h4421115d, 32'h43716eee, 32'h431dacf8},
  {32'hc3b3c848, 32'hc355733d, 32'hc2c89a8f},
  {32'h446d4e5e, 32'h4400caac, 32'hc2732e09},
  {32'hc4691e4d, 32'h42d51cca, 32'h43b70603},
  {32'h43be2926, 32'hc29b4ff5, 32'hc317b808},
  {32'hc313cc00, 32'h43343599, 32'hc32259b5},
  {32'h43088aa0, 32'h4335ddc6, 32'h43c1a8a1},
  {32'hc4944415, 32'hc35cbb53, 32'hc3128ca7},
  {32'h441f87ee, 32'h43a9d50f, 32'h427747c1},
  {32'hc4b10ebf, 32'h4326ec7e, 32'hc1e9814e},
  {32'h44eb53dc, 32'h43425c97, 32'hc3a72aa1},
  {32'hc46119cc, 32'h42ceac65, 32'hc2644d59},
  {32'h431821f0, 32'hc1fc548e, 32'h4007f782},
  {32'hc437b223, 32'h4324cab8, 32'h437428cc},
  {32'h44a196b5, 32'hc29362a2, 32'h435c5852},
  {32'hc474c75f, 32'hc1a71e2c, 32'hc08bac72},
  {32'h4487e6ab, 32'h43408028, 32'hc3f89bea},
  {32'hc4f23adf, 32'hc3087874, 32'hc2c534a3},
  {32'h44d0a1fa, 32'hc31c9573, 32'h422de2f2},
  {32'hc4a01c8e, 32'h42930624, 32'hc21e505b},
  {32'hc347f926, 32'hc32a726d, 32'hc30846cf},
  {32'hc42aa40a, 32'h42c9387d, 32'hc33e4f53},
  {32'h44a96013, 32'h430fe371, 32'hc36f1550},
  {32'hc4e5dfde, 32'h42298610, 32'hc2df0d70},
  {32'h449226f0, 32'hc2acba01, 32'h4287b6b3},
  {32'hc4570a72, 32'hc1ad0cd4, 32'hc38161ac},
  {32'h44c0de12, 32'h431a39fa, 32'hc38c39ef},
  {32'hc3e3feec, 32'h433b3fee, 32'hc3a8dd1d},
  {32'h44a62cc2, 32'h4307d0e7, 32'hc36e8ea5},
  {32'h430fdf90, 32'h43137364, 32'h42c83734},
  {32'h450d4849, 32'hc3b57456, 32'hc2a38416},
  {32'hc50df2e2, 32'hc23beef3, 32'h4301ba6a},
  {32'h43e63873, 32'hc2f44b55, 32'h42c222bf},
  {32'hc454898c, 32'hc3089ae9, 32'h430a946b},
  {32'h4449ef38, 32'h435f4e44, 32'hc39232b1},
  {32'hc4a8aafe, 32'h43a69f3e, 32'h440d3b27},
  {32'h440250a2, 32'h42e1c92c, 32'hc256ebd0},
  {32'hc4d8c890, 32'hc28fbec1, 32'h426e1d2e},
  {32'h446e1d2a, 32'hc39eea91, 32'h42964ce1},
  {32'hc4d12cc6, 32'h43036ce6, 32'hc2dc6425},
  {32'hc23cc960, 32'h430db66a, 32'h420f1c3d},
  {32'hc496db1c, 32'h42af221d, 32'hc26d27d0},
  {32'h44ecf6a0, 32'hc30d9032, 32'h4371dbad},
  {32'hc40670c0, 32'hc317549c, 32'h42389f3f},
  {32'h4410d86d, 32'h41ff6d3a, 32'h423a6e96},
  {32'hc4b9604c, 32'hc2dc8034, 32'h432e4d3e},
  {32'h4507ce42, 32'h437f1887, 32'h4305ddde},
  {32'hc423e0ba, 32'h40fc35fe, 32'hc296d5e0},
  {32'hc2ef9270, 32'hc3d88566, 32'hc409c971},
  {32'hc505b06d, 32'h42a3d85a, 32'hc239528c},
  {32'h44ae3292, 32'h421ef38f, 32'hc3360d1e},
  {32'hc481c16e, 32'h425febce, 32'hc37c78a3},
  {32'h44aa33e2, 32'h4389e89c, 32'hc30120af},
  {32'hc50ec11d, 32'h436b5ffb, 32'h4222e235},
  {32'h450352c6, 32'h410c9c9c, 32'h43d9fc41},
  {32'hc3ddc5ec, 32'hc238821c, 32'hc33a8796},
  {32'h45146e0a, 32'h41e851f9, 32'h428811e3},
  {32'hc4998192, 32'h43ba6dcd, 32'h4369bbc6},
  {32'h451342c0, 32'h4216df36, 32'h43bc62bd},
  {32'hc447e186, 32'h42e9fead, 32'hc27aa552},
  {32'h448199ac, 32'h4218a5d0, 32'hc312af2d},
  {32'hc4f0cb9d, 32'h42283a82, 32'h43cd2efe},
  {32'h438698e6, 32'hc334debf, 32'h4305c2db},
  {32'hc4cd955f, 32'hc37c7012, 32'h4356a416},
  {32'h4506d1c1, 32'h430d8942, 32'h4284ee80},
  {32'hc501cef4, 32'hbe4eb900, 32'hc3989b51},
  {32'h435fda6c, 32'h430358a4, 32'hc3df8992},
  {32'hc4cbfc0c, 32'h41a31658, 32'hc2365124},
  {32'h44f39778, 32'h4302b5a5, 32'h4297fcfa},
  {32'hc44fd088, 32'h43124a7f, 32'h438d56ce},
  {32'h44e4954a, 32'h440a7018, 32'h439abfff},
  {32'hc4619f28, 32'hc2a18d10, 32'hc3a8f6ec},
  {32'h44d2305f, 32'hc3e58e84, 32'hc3a16039},
  {32'hc4d8b9e5, 32'hc2eb68f7, 32'hc3896706},
  {32'h450b8b79, 32'h43969feb, 32'hc414c6f8},
  {32'hc4c9d018, 32'h42a17e3f, 32'hc3783941},
  {32'h44b7b7a6, 32'h4248096f, 32'hc3613b83},
  {32'hc4e751a3, 32'h42d46b91, 32'h431943bc},
  {32'h448c23c3, 32'h426b9cf2, 32'h41a25aa6},
  {32'h4348c47b, 32'hc3a05b5a, 32'h42cd05e2},
  {32'h43ab2fda, 32'hc104e599, 32'hc2a36f03},
  {32'hc3584f54, 32'h44056a75, 32'hc28ae283},
  {32'h43ceac64, 32'hc3954d59, 32'h4347979e},
  {32'hc4048898, 32'hc173026c, 32'hc329ca37},
  {32'h44793955, 32'hc3253db0, 32'hc380d42f},
  {32'hc49d17a0, 32'h4334599c, 32'h42e01d11},
  {32'h44abf9ca, 32'hc2868faa, 32'h4320ce9d},
  {32'hc4c0e188, 32'hc32fc521, 32'hc28fffb0},
  {32'h44225537, 32'hc39605a9, 32'hc397d925},
  {32'hc4389df2, 32'hc3989659, 32'hc397a2c8},
  {32'h44d07cc8, 32'hc17594f0, 32'hc2638198},
  {32'hc4d696f9, 32'h43a45f9c, 32'h43292e90},
  {32'h43a6f868, 32'hc1c53b57, 32'hc2ba47a8},
  {32'hc46afcf5, 32'h425f675b, 32'hc22b95ab},
  {32'h450d01eb, 32'hc3a2afac, 32'hc1c777d4},
  {32'hc4a94d47, 32'hc2baa742, 32'h43762cf8},
  {32'h44fd219a, 32'h43592561, 32'h42ab7a21},
  {32'hc436e066, 32'h41abf275, 32'h4349f610},
  {32'h44c306d9, 32'h42c7d645, 32'h420e08b0},
  {32'hc3a3c600, 32'h434ac715, 32'h438838b4},
  {32'h450ac724, 32'h42ca55e8, 32'h4328e376},
  {32'hc4d07702, 32'h42bdf6ba, 32'h439931cc},
  {32'h44fdcd15, 32'h430ab4c9, 32'h41046978},
  {32'hc39171e4, 32'hc3e43ae9, 32'hc320c2a1},
  {32'h44d10d18, 32'hc2a63b63, 32'hc3213edb},
  {32'hc4a77b44, 32'hc06a5600, 32'hc357ef6b},
  {32'h44aad098, 32'hc2618f09, 32'hc261cad5},
  {32'hc49ead36, 32'hc34e82f6, 32'h4384b9db},
  {32'h44494384, 32'h42a87510, 32'hc3692697},
  {32'hc4efee57, 32'h4202ad3f, 32'hc3820159},
  {32'h442c5276, 32'h43bd222e, 32'h41924ef2},
  {32'hc3a26802, 32'h4288c550, 32'h42774014},
  {32'h44401316, 32'hc39aea34, 32'hc2caeb62},
  {32'hc4da562c, 32'h432271aa, 32'hc32abff0},
  {32'h44f7e2cc, 32'hc33578db, 32'h4342117e},
  {32'hc43177b4, 32'hc1f39e40, 32'h43f88528},
  {32'h441d3172, 32'hc30f9924, 32'hc11ce7e2},
  {32'hc2d4c168, 32'h43b0cdba, 32'hc33c6d10},
  {32'h44f067e1, 32'hc3bbe75c, 32'h438477c5},
  {32'hc4a7aadc, 32'h41a31801, 32'hc30a157e},
  {32'h44ca7206, 32'hc28a4a47, 32'hc3224f14},
  {32'hc4e742d9, 32'h430431ea, 32'h424e89d5},
  {32'h434c93c0, 32'h4380dae2, 32'h428be1ae},
  {32'hc4469c3a, 32'h429b83cc, 32'h42fb196c},
  {32'h437c875a, 32'h4364f547, 32'hc1893ae1},
  {32'hc49586cf, 32'hc38f8e13, 32'hc216e6c2},
  {32'h45049596, 32'h439ed0aa, 32'h430a6c60},
  {32'hc45a9b8c, 32'h43bd629a, 32'hc20e8aa3},
  {32'h44ebd854, 32'hc204a34c, 32'h42e63714},
  {32'hc4d81833, 32'h430bb3d0, 32'h4336cd83},
  {32'h43ab1920, 32'hc31af4af, 32'hc3a1c733},
  {32'hc5025f1c, 32'h42b325ac, 32'h43105bc4},
  {32'h44ba7ea5, 32'h418fea1e, 32'hc1fddece},
  {32'hc4b21d3d, 32'h42a1653f, 32'hc3a7077e},
  {32'h44af2f74, 32'hc380bffa, 32'hc221ca64},
  {32'hc4ebe839, 32'hc34dee90, 32'hc382c970},
  {32'h440a003a, 32'h43712bce, 32'hc2439aec},
  {32'hc511e0f8, 32'hc2922b41, 32'h425cd1f2},
  {32'h4502f8ae, 32'hc307cfc2, 32'hc3bced87},
  {32'hc4d7c5d3, 32'h437dc3fb, 32'h43498cba},
  {32'h440c7230, 32'hc2b6f770, 32'h433646e0},
  {32'hc4160408, 32'h432c295d, 32'hc19b77a7},
  {32'h43c0f5f3, 32'h42f81f45, 32'hc38c61a3},
  {32'hc4f49a6b, 32'hc361251c, 32'hc2eff4f3},
  {32'h43a5b5a0, 32'hc413e9d9, 32'hc29302c6},
  {32'hc47e6cb1, 32'hc294166b, 32'hc33b6f44},
  {32'h44f23670, 32'hc30111de, 32'hc2c73044},
  {32'hc37a4c08, 32'hc33521d4, 32'h435ce58f},
  {32'h44f6ca74, 32'h409aa4c6, 32'hc326de0d},
  {32'hc479103c, 32'h42b4e29a, 32'h441285ef},
  {32'h42002b1c, 32'h43107c56, 32'hc280b63d},
  {32'hc418eff0, 32'h43ce6d2e, 32'h43b2fbad},
  {32'h449b7eb8, 32'hc3508b55, 32'h43636efa},
  {32'hc48c63c7, 32'h43d1646c, 32'h429bd546},
  {32'h448a5278, 32'h41b2db9f, 32'h421959e9},
  {32'hc47bb3f8, 32'h427cc635, 32'hc2d4f137},
  {32'h44e4d0cf, 32'hc31321cb, 32'h42b219d9},
  {32'hc4495658, 32'h439281e4, 32'hc36f6118},
  {32'h44685813, 32'h426cee83, 32'hc3ca0196},
  {32'hc41bc01a, 32'h4313b24a, 32'h43bbe74e},
  {32'h45046a99, 32'h42745c0d, 32'h437b649c},
  {32'hc4b7336e, 32'hc32767ee, 32'h4410f7b6},
  {32'h4266d0d0, 32'h42893ad9, 32'h4260c04e},
  {32'hc4d204dc, 32'h40799aaa, 32'hc25f4b68},
  {32'h4475ad7c, 32'hc3503176, 32'hc3934677},
  {32'hc473ee18, 32'h43131ad0, 32'hc240d436},
  {32'h44dff710, 32'h4375de82, 32'hc2364d56},
  {32'hc50f2cf4, 32'hc3423025, 32'h4327cb4c},
  {32'h43d9b30c, 32'h435a72ce, 32'h43364fd5},
  {32'hc509740d, 32'hc3418670, 32'h41076251},
  {32'h44258866, 32'hc210f8a9, 32'h434a9667},
  {32'hc4f49265, 32'hc25b722e, 32'hc2bab2f3},
  {32'h45156410, 32'hc2b1d5cf, 32'h42bc81c7},
  {32'hc50411aa, 32'h4319db6b, 32'h42bbd997},
  {32'h442b1d0a, 32'h43644501, 32'hc32d39de},
  {32'hc4611860, 32'hc3ee1fe6, 32'hc284f816},
  {32'h43e48a92, 32'hc392f185, 32'h4294245c},
  {32'hc4d04511, 32'h42d10c39, 32'h42b80f68},
  {32'h44279966, 32'h4348203b, 32'hc3034b89},
  {32'hc4bcf0d6, 32'hc2a8ddc7, 32'h4281f976},
  {32'h44dfca51, 32'hc27c479d, 32'h438ae910},
  {32'hc4455522, 32'hc227f9e9, 32'hc224555a},
  {32'h44ecfdec, 32'h4309547f, 32'hc4301193},
  {32'hc3d50745, 32'hc227caae, 32'hc1dab036},
  {32'h44ce7206, 32'hc38996bd, 32'hc38bd2da},
  {32'hc4253a2d, 32'hc3652512, 32'hc3bff9c6},
  {32'h440ea1db, 32'hc341622e, 32'hc31ec05d},
  {32'hc4cbd348, 32'hc39c7b0e, 32'hc3034f23},
  {32'h44aadce5, 32'hc22eff9d, 32'hc3951ecc},
  {32'hc4a61be7, 32'h43196c50, 32'hc33885ef},
  {32'h44b23ce0, 32'h43735c8c, 32'hc3689295},
  {32'hc47da563, 32'h4323d9cd, 32'hc379cc87},
  {32'h44d318ef, 32'hc1881075, 32'hc2826516},
  {32'hc4f69adc, 32'hc343177f, 32'h433774f3},
  {32'h4512082a, 32'h431ce2fe, 32'h426c75dd},
  {32'hc4f8a1a0, 32'hc324431d, 32'h4328a61d},
  {32'h44c280e8, 32'h439ae958, 32'hc23fc2ba},
  {32'hc4d4220f, 32'h425bf572, 32'h43744c90},
  {32'h44b98ddc, 32'hc32dfc64, 32'h42fb6d73},
  {32'hc50aa1d8, 32'hc1991120, 32'hc24696a8},
  {32'h43b22e42, 32'hc2b40b74, 32'h4237c96a},
  {32'h430fb718, 32'hc3053862, 32'hc386fd46},
  {32'h44f09494, 32'h433c37e6, 32'hc3837ccf},
  {32'hc4a63188, 32'h42c99b52, 32'hc1d08d76},
  {32'h44dda9e2, 32'h43ce5d4d, 32'hc110c596},
  {32'hc4125c44, 32'h430dfec2, 32'h433f9d65},
  {32'h44132eb4, 32'h43373706, 32'h43246a78},
  {32'hc512c07b, 32'hc22015c4, 32'hbf62b564},
  {32'h450b1805, 32'hc16e32d8, 32'hc31fa367},
  {32'hc484aa3c, 32'hc1834ce2, 32'hc3306904},
  {32'h44cd1237, 32'hc352f23e, 32'h43f8b15c},
  {32'hc51c4330, 32'h43918aca, 32'hc23c6549},
  {32'h44942538, 32'hc2f2b9c1, 32'hc3a61dec},
  {32'hc51320fd, 32'hc380fab3, 32'h42c95fb9},
  {32'h4515c128, 32'h4339a6dc, 32'hc2401195},
  {32'h4200ea40, 32'hc4242aa4, 32'h4345ab57},
  {32'h45275b32, 32'h4389aa37, 32'h42a66a60},
  {32'hc34cd90c, 32'h425be106, 32'h429d09dc},
  {32'h4501c166, 32'hc297447a, 32'hc2e8c541},
  {32'hc4d17245, 32'h41d78a05, 32'h4053e42b},
  {32'h44a47b64, 32'hc2a29f99, 32'h43c12727},
  {32'hc508e635, 32'h428501e1, 32'h428d7a53},
  {32'hc26224d0, 32'h4356e1d1, 32'h4379c146},
  {32'hc4d08c60, 32'hc3036ef2, 32'hc2fd3661},
  {32'h447a83d4, 32'h43c37bff, 32'h4234b045},
  {32'hc5035b5d, 32'h420f4f59, 32'hc34968ee},
  {32'h44e72db3, 32'hc34ea267, 32'hc375382a},
  {32'hc484edc6, 32'hc34d2085, 32'hc2ce2f2d},
  {32'h43ad82e4, 32'hc2f5d9c6, 32'h432ca7b3},
  {32'hc33f91f1, 32'h42484fa1, 32'hc38bac10},
  {32'h44f9975e, 32'h42584bad, 32'hc34b6ef2},
  {32'hc424f297, 32'h4188845a, 32'hc36879f3},
  {32'h450f902b, 32'hc335bbe0, 32'h43c90146},
  {32'hc490f52a, 32'hc303c644, 32'h432b92f6},
  {32'h43c033e0, 32'hc3d96a4b, 32'h42434921},
  {32'h428a8b20, 32'h42433350, 32'h42d1fae7},
  {32'h441aa86a, 32'hc37378f4, 32'h42ac106b},
  {32'hc450c932, 32'h3fdd5068, 32'h43c832b6},
  {32'h45145549, 32'hc3c4e817, 32'hc3ef093d},
  {32'hc3d468c8, 32'hc3994f3f, 32'hc324d64e},
  {32'h40aa4c00, 32'h42c7e174, 32'hc31b059f},
  {32'hc4a497d3, 32'h435e7f13, 32'hc1dd491c},
  {32'h4517e0a1, 32'hc28c6584, 32'h429bb5dd},
  {32'hc4e2c4f2, 32'hc33aeb9d, 32'h4232b229},
  {32'h4516eb52, 32'h43703661, 32'h439e35b5},
  {32'hc481360a, 32'hc1967471, 32'h4305303d},
  {32'h450f127d, 32'h418370ae, 32'h42cc9b8f},
  {32'hc0eecc40, 32'h428ab82d, 32'hc387be8d},
  {32'h44453232, 32'h42927526, 32'h430f0a40},
  {32'h421a8522, 32'h430a3715, 32'hc3b83ada},
  {32'h43dcc7a0, 32'h4380d32f, 32'h42a0a496},
  {32'hc4a99339, 32'h43bff40c, 32'h43b3bdd5},
  {32'h44878ab0, 32'hc2bd7509, 32'hc3454a8e},
  {32'hc428d832, 32'h438d4df1, 32'h420407be},
  {32'h43e37708, 32'hc3ec7672, 32'hc3300c64},
  {32'hc4b7010a, 32'h4027a2cc, 32'h438491ec},
  {32'h44c1158f, 32'hc3041ba6, 32'hc3273c37},
  {32'hc42288db, 32'hc39e4d9d, 32'hbea07a20},
  {32'h446b919e, 32'h4380b892, 32'h41e6f1a4},
  {32'hc498f020, 32'h4290aa70, 32'hc33b4781},
  {32'h43f2c300, 32'hc3d4f421, 32'h42267da2},
  {32'hc4b241a8, 32'h4344c2bb, 32'h43d93f6d},
  {32'h44589ca0, 32'h42c5f90b, 32'h41a5eea2},
  {32'hc3e27892, 32'h425c1a69, 32'hc39dd142},
  {32'h44c2cece, 32'hc18165b2, 32'hc22cdc75},
  {32'hc3cf94f1, 32'hc3e3f99a, 32'h42b444c7},
  {32'h450e5457, 32'hc2fcada9, 32'h43916a51},
  {32'hc4da4c3b, 32'hc32e9f41, 32'h4357e0a9},
  {32'h4502f5c7, 32'hc26923a5, 32'h4186451a},
  {32'h43bb2df1, 32'hc39b7909, 32'h43367035},
  {32'h44d5ad49, 32'h4307267a, 32'h41a623ee},
  {32'hc4835fd1, 32'hc32d210e, 32'hc41420b3},
  {32'h4503880b, 32'h434c4958, 32'h440865d3},
  {32'hc4daa900, 32'h4340299f, 32'hc2c246bb},
  {32'h43fb98af, 32'h42b1dfb3, 32'hc2bb367f},
  {32'h44017918, 32'hc30bc026, 32'h420152d8},
  {32'h4418c4ac, 32'hc2aa5468, 32'h4248c338},
  {32'hc4f7b40f, 32'h433c3db3, 32'h43446422},
  {32'h44900f04, 32'h42003538, 32'h4293eb38},
  {32'hc43e5c29, 32'hc3510080, 32'hc3056eb5},
  {32'h442a87f4, 32'h43747bb9, 32'h42271b1e},
  {32'hc476be35, 32'h40f47af2, 32'hc3db1743},
  {32'h43559f4e, 32'hc1c9fe14, 32'h43a4e45b},
  {32'hc4259c72, 32'hc3cef230, 32'hc20dc117},
  {32'h44da38fd, 32'hc1e26060, 32'h43818aa0},
  {32'hc4d7a866, 32'hc156749c, 32'hc3abb5bb},
  {32'h42d3dbe0, 32'hc3e0fa6d, 32'h431c2a07},
  {32'hc4e45f4f, 32'h43a5faa9, 32'hc30eecb3},
  {32'h44eb22ac, 32'h439f869e, 32'h430d9ef8},
  {32'hc4a5a260, 32'h4299777c, 32'hc33a6acf},
  {32'h442cd950, 32'hc37a7fff, 32'h4394dd1d},
  {32'hc50c2457, 32'hc3a27bc6, 32'hc33a2331},
  {32'hc24c9e48, 32'h43976ae8, 32'hc2d0c182},
  {32'hc30f8586, 32'h4279915b, 32'hc1d4f826},
  {32'h4383837a, 32'h43e332f3, 32'h436be3fd},
  {32'hc3e4dd76, 32'hc30f2975, 32'hc3613d4a},
  {32'hc47ba16b, 32'h42ed076e, 32'h43770f68},
  {32'h41371a00, 32'hc2117212, 32'h4325d0f6},
  {32'hc4bd891a, 32'h4237a022, 32'h422dea7a},
  {32'h44fbb183, 32'h43b067a4, 32'h431f6571},
  {32'hc45b1eb6, 32'hc2f4fea5, 32'hc2bad44b},
  {32'h4420fbba, 32'hc3bd07d6, 32'h43ef25a7},
  {32'hc50c796a, 32'h432f1cc0, 32'hc357f58e},
  {32'h44724108, 32'hc25a0d00, 32'h42949839},
  {32'hc44bcfcb, 32'h43b5ff96, 32'h4118f919},
  {32'h44cccc90, 32'h4242109a, 32'hc315a4b8},
  {32'hc4bf76de, 32'h42766335, 32'hc3cceecb},
  {32'h44da5349, 32'h43d8d16b, 32'hc3bf2d45},
  {32'hc4825db1, 32'h439c08b8, 32'hc2dfbacb},
  {32'h44e9cad6, 32'h42f6a5a0, 32'h433a313d},
  {32'hc415e952, 32'h440222ba, 32'hc333ba7e},
  {32'h45009692, 32'h435036d7, 32'hc2f72bd2},
  {32'hc48cc7d7, 32'h432f32bc, 32'hc28a077c},
  {32'h4507d901, 32'h43437de1, 32'h433af724},
  {32'hc4331b66, 32'h43ce7265, 32'hc30c3adc},
  {32'h434ed970, 32'h4347323f, 32'hc112cdd2},
  {32'hc3e92d70, 32'h43001771, 32'hc3efd546},
  {32'h450292c8, 32'h4349d141, 32'h4324dc52},
  {32'hc462ca3a, 32'h42c3d7b6, 32'h42ce9549},
  {32'h448e9be1, 32'hc281a11a, 32'h43c246a5},
  {32'hc410499a, 32'h43947b7c, 32'hc311d248},
  {32'h4502e455, 32'hc1322a72, 32'h41d96c46},
  {32'hc4e76174, 32'hc3dd5ebb, 32'h436e1c29},
  {32'hc2d9efc9, 32'hc29e3540, 32'hc1ade0df},
  {32'hc4fb6930, 32'hc16a3aea, 32'hc336c839},
  {32'h4485ab20, 32'hc2a1e7b3, 32'hc3056d80},
  {32'h42fe0f94, 32'h41031aca, 32'hc2e56dc7},
  {32'h4500f5ff, 32'hc1ae01d4, 32'h43d531b1},
  {32'hc494791e, 32'h429dee83, 32'hc3761e19},
  {32'h44db0640, 32'h42a245d0, 32'h431196b8},
  {32'hc5110ec3, 32'hc31d90a1, 32'hc28608b6},
  {32'h44a1b7c8, 32'hc35836bd, 32'h41f6d268},
  {32'hc3f2600a, 32'hc37336c4, 32'hc38e3337},
  {32'h44fb395c, 32'hc3a5c2b4, 32'hc2ac0305},
  {32'hc44220d0, 32'hc3ac3607, 32'h43213266},
  {32'h443ccce6, 32'h43c77c5c, 32'h434e0160},
  {32'h4384a3c7, 32'h429e350c, 32'hc3a3e8d4},
  {32'h43ee4708, 32'h4273db03, 32'hc2fca914},
  {32'hc502c447, 32'h42a0da25, 32'h43537bab},
  {32'h44b98bc6, 32'h42b80159, 32'hc3688506},
  {32'hc3fcaada, 32'hc24ce9e5, 32'hc39a0745},
  {32'h44d72b14, 32'hc0e9a270, 32'h437d4cd4},
  {32'hc480b1dc, 32'h4352868a, 32'hc389e53d},
  {32'h451fc740, 32'h4301ec08, 32'h42975f0d},
  {32'hc4eb56ec, 32'h42da710b, 32'hc18c721b},
  {32'h44f2fbac, 32'h43540abc, 32'hc2f4b81a},
  {32'hc40b47d4, 32'h43b9d399, 32'hc344c2e5},
  {32'h44a49203, 32'hc2b742c8, 32'h43208060},
  {32'hc3fc1d8e, 32'hc36ae6cf, 32'h43ab8ac1},
  {32'h44f812f2, 32'h41cff077, 32'hc23750be},
  {32'hc4ef48be, 32'h438269d0, 32'h4254a15a},
  {32'h43eeaac5, 32'h42b8a1e6, 32'hc36dfa6c},
  {32'hc4a6e51e, 32'hc2a13597, 32'hc380a26d},
  {32'h44741bb9, 32'hc394e3e5, 32'hc4165a67},
  {32'hc502f602, 32'hc242fb59, 32'hc2bfc00e},
  {32'h4407405b, 32'hc36be326, 32'hc2e8b6a7},
  {32'hc5145c98, 32'hc2b3380f, 32'h42bfa750},
  {32'hc29cc2d0, 32'h4408719c, 32'hc38fa6b3},
  {32'hc4cd062f, 32'hc1d79bb6, 32'hc386f08d},
  {32'h445aa568, 32'hc2f6876f, 32'h421fb574},
  {32'hc49f5965, 32'h4314ccda, 32'h4192b8cb},
  {32'h43460920, 32'h41f62692, 32'hc3e23a53},
  {32'hc44ccec0, 32'hc2246222, 32'h4380e7c3},
  {32'h44190f35, 32'hc3bae4e8, 32'hc2d8cf7a},
  {32'hc4d7d8b4, 32'hc207379c, 32'hc30d26d3},
  {32'h43aebfbc, 32'hc370810a, 32'h41002f4a},
  {32'h43b45810, 32'h42a34b01, 32'hc32b97d4},
  {32'h43965aa8, 32'hc2bd8c27, 32'h436d6064},
  {32'hc44f4db3, 32'h42a894e5, 32'hc2434de3},
  {32'h40be4a00, 32'h43393775, 32'hc361a36e},
  {32'hc495911a, 32'hc36f54bf, 32'h43c87b11},
  {32'h42c4aab8, 32'h42ba3658, 32'h43b2f73a},
  {32'hc3129117, 32'hc3adc4b9, 32'hc332026d},
  {32'h4510e73a, 32'h43c8cd03, 32'h42b10e0a},
  {32'hc47eb76a, 32'hc32c06cb, 32'h41f84044},
  {32'h44d51e4b, 32'hc301714a, 32'hc2e5441b},
  {32'hc4e4a602, 32'h42877d36, 32'h42c27b78},
  {32'h43e85570, 32'h42a68620, 32'hc2821c47},
  {32'hc3aebd8c, 32'h434e1514, 32'hc17bc6aa},
  {32'h44a26b62, 32'hc26b1c45, 32'h42e817b4},
  {32'hc4321d98, 32'h435f7741, 32'h432bbd4d},
  {32'h431ce060, 32'h429226c4, 32'hc341ef37},
  {32'hc4ca9fc8, 32'h3f09073c, 32'hc0757acb},
  {32'h44e48776, 32'h4393f963, 32'hc369c010},
  {32'hc4eaff14, 32'h433a625c, 32'h4222d5f4},
  {32'h44841200, 32'hc38fc534, 32'hc407c5f9},
  {32'hc47cdbc0, 32'hc3a9c68b, 32'h43cd55f5},
  {32'h44a30952, 32'hc317d3ca, 32'hc2835d2a},
  {32'hc354d970, 32'h4139d302, 32'h431b08d5},
  {32'h44f9b61a, 32'hc38c2dc9, 32'hc39ec61e},
  {32'hc304c4a8, 32'h427e9559, 32'h431495c3},
  {32'h4444bc7c, 32'h4314fa68, 32'hc2dd234a},
  {32'hc49e2ee1, 32'h42d499fa, 32'h42a707ee},
  {32'h43838fbe, 32'hc39950cf, 32'hc3a44dde},
  {32'hc4a3f762, 32'hc2cd180b, 32'hc33a3a2e},
  {32'h44c1bcd0, 32'hc28d6881, 32'hc39375a4},
  {32'hc510b0a2, 32'h430f7e00, 32'hc2ae7c6c},
  {32'h44d5dfb4, 32'h3fca27ff, 32'h43711db2},
  {32'hc4d86014, 32'hc32e6db7, 32'hc35bf4e4},
  {32'h44d1c1f6, 32'h41a2c521, 32'h4357c096},
  {32'h427e993d, 32'h42c6fb84, 32'h43e31773},
  {32'h446c6540, 32'hc2e01c2d, 32'hc28ad3c9},
  {32'hc5016479, 32'hc2cf2c6d, 32'h42a4121b},
  {32'h4506d86e, 32'hc31e715a, 32'hc3a50d73},
  {32'hc444e666, 32'h4301b1a7, 32'hc332bb1a},
  {32'hc2955b50, 32'h431e38b8, 32'hc3875a64},
  {32'hc4f156f8, 32'hc333b461, 32'h4341ba30},
  {32'h4491dea1, 32'hc2ddf5ed, 32'h4336e005},
  {32'hc28eece8, 32'hc40bbc7d, 32'h43a68c23},
  {32'h43c3dd18, 32'hc3d423a1, 32'h43ebde2e},
  {32'hc510e162, 32'hc2884cff, 32'h439f1456},
  {32'h43d7fbf8, 32'h4403168f, 32'h42cecd92},
  {32'h43d71da0, 32'h43016358, 32'hc2dceb3f},
  {32'hc460eb9a, 32'hc2802aa4, 32'h42da53db},
  {32'h43b1f06e, 32'h43d23ac7, 32'h432fb3e2},
  {32'hc4ef6c79, 32'hc0f5c615, 32'hc2bf058a},
  {32'h450c865c, 32'hc3eb089d, 32'h4399dfc4},
  {32'hc48ba42b, 32'h40a7d035, 32'hc36c7bd4},
  {32'h444338e6, 32'h412e1740, 32'hc2c546f8},
  {32'hc4207354, 32'h420fac86, 32'h41b78a10},
  {32'h43ea8c68, 32'hc1782444, 32'h4284f9cc},
  {32'hc501bfed, 32'hc3a66ddd, 32'hc352b417},
  {32'h4508db37, 32'hc3b0720c, 32'hbe705800},
  {32'hc50339c4, 32'hc38d6d25, 32'hc369451a},
  {32'h450c51a1, 32'hc3059050, 32'hc2f49542},
  {32'hc2c5b244, 32'hc406be4b, 32'hc23101cc},
  {32'h44b19cd6, 32'h428aa5b7, 32'h42d44205},
  {32'hc48d1f5a, 32'h43274539, 32'h41efd416},
  {32'h440717ec, 32'h429c805e, 32'hc322e611},
  {32'hc48876d3, 32'hc3385377, 32'hc28f4222},
  {32'h451780f2, 32'hc3ac2df1, 32'hc31cedf3},
  {32'hc3351bf8, 32'h43097e8c, 32'h4271366b},
  {32'h448dfa28, 32'hc3b83aa7, 32'hc2ba8d62},
  {32'hc43cf760, 32'hc397aa47, 32'h42010e4c},
  {32'h438159a0, 32'h434c3f24, 32'hc240a482},
  {32'hc3743948, 32'h432bf4aa, 32'h432577fc},
  {32'h4444e34e, 32'hc391f8a7, 32'hc2b7f0e9},
  {32'hc44998e2, 32'hc365f6f7, 32'h42b71d9f},
  {32'h4423c852, 32'h429bfb51, 32'h43860a98},
  {32'hc4f4b223, 32'h432cac37, 32'h4302452f},
  {32'h44789924, 32'hc2dc8c3b, 32'h438b4ce7},
  {32'hc383d099, 32'hc40b3ac0, 32'h43aa7475},
  {32'h44e8d5a2, 32'hc3083a6e, 32'hc3887b72},
  {32'hc4de53b9, 32'h41dd5016, 32'hc34ad278},
  {32'h4371748e, 32'h43589dd6, 32'h430b173f},
  {32'hc4c1c77a, 32'hc3057a8d, 32'hc330ab47},
  {32'h44ad5cb2, 32'h433b5886, 32'hc3878692},
  {32'hc4da0c06, 32'h43669e68, 32'h43535d66},
  {32'h44bc908f, 32'h4362e670, 32'h418e070c},
  {32'hc4284bde, 32'hc2dbc326, 32'h429f7967},
  {32'h44b89b04, 32'h43750064, 32'hc3814281},
  {32'hc3e3edd0, 32'hc3a3e7d0, 32'h4085d978},
  {32'h44618660, 32'hc398f740, 32'hc0f6a2d4},
  {32'hc4d815ba, 32'h408653c2, 32'hc3b344e9},
  {32'h44a24540, 32'hc2cce562, 32'h4294db77},
  {32'hc33f8364, 32'h41e9898d, 32'h4239f367},
  {32'h43b85124, 32'h42ed87fb, 32'hc16aa80c},
  {32'hc3bf8780, 32'hc25df32a, 32'h43031ddb},
  {32'h44dfc0f2, 32'hc36e8dd6, 32'hc356473e},
  {32'hc3e28798, 32'hc3dd1f5d, 32'h4323ab24},
  {32'h44f1dc1d, 32'h41b7fe82, 32'hc207cf8a},
  {32'hc13a977c, 32'hc2d5c8ac, 32'hc207eef0},
  {32'h449d8487, 32'hc29d229a, 32'hc395b0b9},
  {32'hc5054ad1, 32'h43b306ae, 32'hc32a0e58},
  {32'h43c55a48, 32'h434771e5, 32'hc3499493},
  {32'hc5090d33, 32'h42fd6542, 32'hc2f45a6a},
  {32'h44827497, 32'hc36c7e41, 32'h426c3f53},
  {32'hc3762440, 32'h434eaba5, 32'hc3809284},
  {32'h45016832, 32'h400ea270, 32'h43cd212f},
  {32'hc4d46faa, 32'hc3607be7, 32'h42173688},
  {32'hc3917a50, 32'h43e8e7b4, 32'hc1842780},
  {32'hc467c48d, 32'h43a17a6c, 32'h421c48a9},
  {32'h448d4d9c, 32'hc33354a6, 32'hc388a1c9},
  {32'hc4f4be71, 32'hc354a9f4, 32'hc3017644},
  {32'h449569b7, 32'h42b85e66, 32'h43a0e431},
  {32'hc4de1c02, 32'h42d4baa0, 32'hc314ea27},
  {32'h440a1804, 32'h4382f9eb, 32'hc38f648e},
  {32'hc464d6df, 32'h411906eb, 32'h4299f8cb},
  {32'h446f66b0, 32'h43555d6d, 32'hc35f6577},
  {32'hc3e0257a, 32'hc307a2ee, 32'h4306faae},
  {32'h414db100, 32'h41d5e910, 32'hc16c73a0},
  {32'hc1a93980, 32'h42e05250, 32'hc3160448},
  {32'h4508dbb8, 32'h43062383, 32'hc3979a98},
  {32'hc507f3ae, 32'h43adcec6, 32'hc3bd6c36},
  {32'h45048678, 32'hc3925ded, 32'hc2b3aebc},
  {32'hc49c98e9, 32'hc2a163fe, 32'hc3a7bd09},
  {32'h42b627f0, 32'hc34e085d, 32'hc2269915},
  {32'hc3c7108c, 32'hc2cfdbd8, 32'hc2898d2b},
  {32'h44ab18ec, 32'h42eba8db, 32'h43345cce},
  {32'hc50ae335, 32'h41af643e, 32'hc38948bc},
  {32'h4364c24e, 32'h4401b7f6, 32'h430b53d0},
  {32'hc43e6a04, 32'hc222b0cd, 32'h42d1e5d8},
  {32'h448dc269, 32'hc35c5526, 32'hc337089e},
  {32'hc38fcc50, 32'h43b446e1, 32'hc2d8e47b},
  {32'h4491962d, 32'h4205f7d6, 32'h4289ac29},
  {32'hc4ba6aa2, 32'h4357b62a, 32'h4370bab1},
  {32'h442b78f2, 32'hc34f34aa, 32'h433570c7},
  {32'hc500c62c, 32'hc33f600c, 32'hc2a95760},
  {32'h44b36142, 32'h42147ca7, 32'hc31f8f3d},
  {32'hc18a8e00, 32'hc20dc297, 32'h43fb9b1f},
  {32'h44f7376a, 32'h43d7137f, 32'hc15deb76},
  {32'hc4130e1e, 32'h43db9b6d, 32'hc19282fd},
  {32'h44ca159e, 32'h436b34c1, 32'h43768e39},
  {32'hc483ceee, 32'h43a7532a, 32'hc31603cc},
  {32'h44700806, 32'hc3daa079, 32'h43000f3a},
  {32'hc41bcd43, 32'hc3ad26e7, 32'hc0aa3433},
  {32'h4421c760, 32'hc2f76964, 32'h436ff0b9},
  {32'hc3f269fc, 32'hc14dbdad, 32'h432be23f},
  {32'h44989116, 32'hc2b6daed, 32'h4332aa0d},
  {32'hc477eab3, 32'h425bfe64, 32'h4268daa7},
  {32'h45097eec, 32'h438e4569, 32'hc3e806fb},
  {32'hc4543d0a, 32'hc2a57065, 32'hc3186145},
  {32'h44aebaf6, 32'hc30779f4, 32'hc2ad75fb},
  {32'hc48bb264, 32'hc17716a1, 32'hc091bb6a},
  {32'h448f00f9, 32'h4484dc23, 32'h4343513e},
  {32'hc3a74f2c, 32'h41d6f8d1, 32'h4263e687},
  {32'h43cd1d35, 32'h42925f3e, 32'h435b9168},
  {32'hc4986b96, 32'hc3c0ec9e, 32'hc3dbd139},
  {32'h4401515c, 32'h3edd5c0b, 32'hc36d69c7},
  {32'hc4d7d8c3, 32'hc38d3016, 32'h42c67239},
  {32'h4423c92a, 32'hc31cf990, 32'hc3d49dec},
  {32'hc43fce2c, 32'hc41e9212, 32'hc343f090},
  {32'h44fea374, 32'hc32a7463, 32'hc305b617},
  {32'hc412d753, 32'hc376adda, 32'h428fd3c6},
  {32'h43a9ba54, 32'h429acfcb, 32'h429f26ee},
  {32'hc2455b20, 32'h433c54c2, 32'hc2c646f0},
  {32'h4526ad12, 32'h43a0bf88, 32'hc3a3aa8c},
  {32'hc42dfdbf, 32'hc3113676, 32'hc32d3338},
  {32'h44b74d8b, 32'h43c825cc, 32'hc395d97c},
  {32'hc4bcb5ac, 32'hc3c2ea92, 32'hc2165e45},
  {32'h43110e60, 32'hc3246cd5, 32'h43e13b01},
  {32'hc2c2b120, 32'h42b6c008, 32'h42fd2273},
  {32'h44b29f66, 32'h4383de5b, 32'hc3229e0d},
  {32'hc32fdd22, 32'hc2120979, 32'h42681c03},
  {32'hc21ab430, 32'h43307d56, 32'hc11fb984},
  {32'hc4d2945e, 32'hc32361f0, 32'hc3549e7a},
  {32'h4474140b, 32'hc2c6e2f6, 32'h42ef1856},
  {32'hc4a12b56, 32'h42a77da7, 32'hc1a9bed5},
  {32'h44f14d83, 32'h42a94b40, 32'h438bde63},
  {32'hc471b81c, 32'h43b490ef, 32'h42ff3487},
  {32'h44ff37cb, 32'hc32abc63, 32'h4387057b},
  {32'hc4fe86e2, 32'hc364bbad, 32'hc3bdacbf},
  {32'h447864de, 32'hc2e9fc67, 32'hc379fe89},
  {32'hc2f179f0, 32'h42c25554, 32'hc2fc85f6},
  {32'h44eee931, 32'h43dfad34, 32'hc3b0f002},
  {32'hc4e3525e, 32'hc3bd0fe0, 32'hc36f28f4},
  {32'h45062ee6, 32'h4347ee35, 32'h43dddd1d},
  {32'hc26f8b40, 32'hc1901561, 32'h4314983e},
  {32'h44950657, 32'h43964931, 32'hc2827cba},
  {32'hc414c342, 32'hc2f6ba7e, 32'hc2b951db},
  {32'h44655352, 32'h42d8537d, 32'hc32fd97a},
  {32'hc4cf8e1c, 32'hc3ff3a16, 32'hc41218d0},
  {32'h449e8862, 32'h43232279, 32'h42af4a84},
  {32'hc39ca4f0, 32'hbf686200, 32'hc35b13b8},
  {32'h44a8907b, 32'hc2b30860, 32'hc1cbb3c8},
  {32'hc4ac19b8, 32'hc3852fa9, 32'h439cf1b0},
  {32'h44b3baa6, 32'h4388248d, 32'h4284f3e5},
  {32'hc342b400, 32'hc2220b05, 32'h433fc44c},
  {32'h45059ad2, 32'h4381edfe, 32'hc38c8199},
  {32'hc4b73f22, 32'hc1015440, 32'hc29d7d44},
  {32'h4404d823, 32'h4366cdd8, 32'h437020c1},
  {32'hc4779b8f, 32'hc27edba1, 32'hc2588840},
  {32'h450d96ca, 32'h4394cb50, 32'h42ee4341},
  {32'hc3ee73a0, 32'h433e7869, 32'h431cacad},
  {32'h44f21ee1, 32'hc314bbcc, 32'hc3a4ad83},
  {32'hc4b3a953, 32'hc385c2a7, 32'hc33b30d0},
  {32'h4490a5da, 32'h438af3a1, 32'hc28272cc},
  {32'hc41d1a5c, 32'hc3a71858, 32'hc31086d5},
  {32'h4253a1e0, 32'h42febbed, 32'hc2e29558},
  {32'hc383ba3e, 32'hc3e9325d, 32'hc3da86fa},
  {32'h44a7662a, 32'h4312d443, 32'h438c05d8},
  {32'hc4255fc7, 32'hc2d13214, 32'hc26c322d},
  {32'h43cfb454, 32'hc2d56d3c, 32'h42c91f62},
  {32'hc4f4c7fe, 32'h4248fdb5, 32'h432bb6eb},
  {32'h4469fb4e, 32'hc29d6427, 32'h43473b83},
  {32'hc4af9bd6, 32'h43a1ffb5, 32'h42a667ec},
  {32'h435c93bc, 32'h42357878, 32'hc3c1cd4b},
  {32'hc4006170, 32'h4387c084, 32'h434bdfba},
  {32'h4507c824, 32'hc38f069b, 32'h42ec135d},
  {32'hc4809064, 32'h42e2d810, 32'h42f20a72},
  {32'h44b60293, 32'hc2eceead, 32'h42687345},
  {32'hc501f918, 32'hc3343372, 32'hc369b396},
  {32'h44b640eb, 32'hc2a54078, 32'hc3b2d4d5},
  {32'hc4ba4d94, 32'hc2b30c89, 32'h4316db27},
  {32'h450a9b19, 32'hc2acad3c, 32'h42967f46},
  {32'hc4d8447d, 32'h427933cd, 32'hc34cb894},
  {32'h45095595, 32'hc3cfe9cc, 32'hc1b102cb},
  {32'hc5048591, 32'hc406afbb, 32'h4386cdd4},
  {32'h4499c6e6, 32'h4428543e, 32'h4378e9b7},
  {32'hc4bad451, 32'h44044890, 32'hc3132093},
  {32'h44ad2709, 32'hc2e51633, 32'hc34856ec},
  {32'hc4181cc4, 32'h439a8a06, 32'h410e9e38},
  {32'h44db30c5, 32'hc3a3bf76, 32'h433cf2a8},
  {32'hc4de3d4a, 32'h43b79765, 32'h439dc545},
  {32'h452251e4, 32'hc31acf66, 32'hc2c64e6c},
  {32'hc514af22, 32'hc32e041c, 32'hc364c9d7},
  {32'h4461a9e3, 32'h43788aa6, 32'hc1a8fbc8},
  {32'hc3923e8a, 32'h40843758, 32'hc32303f5},
  {32'h443962bc, 32'hc2f15e9f, 32'hc3d36d93},
  {32'hc4b3eaa1, 32'h431c39af, 32'hc3e4dbdb},
  {32'h45025dcf, 32'h42a277bd, 32'h439dc151},
  {32'hc483ec54, 32'hc3b7a81d, 32'hc3c27715},
  {32'h43b7eece, 32'hc29eb61a, 32'h42f42fba},
  {32'hc4ab32a0, 32'hc2c3c1c6, 32'h427b8dfc},
  {32'h449047fe, 32'h434847f4, 32'hc25420c5},
  {32'hc49bd85d, 32'hc2187937, 32'h438b47cc},
  {32'h43a0d988, 32'h42094617, 32'h43a6f076},
  {32'hc470bca7, 32'hc33a1a24, 32'hc2439b2f},
  {32'h449f7516, 32'hc26b9481, 32'hc22b2b7e},
  {32'hc34383fa, 32'hc3ab3d46, 32'hc31a05c2},
  {32'h448cde68, 32'h43a1237f, 32'hc380155a},
  {32'hc34f87c7, 32'hc247af0b, 32'h4238a20d},
  {32'h43d4c78c, 32'hc3adb1d2, 32'h43b58c36},
  {32'hc2ec3aa8, 32'hc28dc352, 32'h4382f995},
  {32'h44e8518e, 32'hc325aad1, 32'hc0fe471f},
  {32'hc4c12d13, 32'h4291a674, 32'hc3bd7000},
  {32'h4501d722, 32'hc382c927, 32'h4319404d},
  {32'hc444153a, 32'h42bb9b13, 32'hc3aa8c25},
  {32'h44d8f012, 32'h430638bf, 32'h4338336f},
  {32'hc33e8dfa, 32'hc1d93451, 32'h42d49476},
  {32'h44e30ef2, 32'hc2967a5e, 32'h431c0b1f},
  {32'h41fbdbc0, 32'hc338bc9a, 32'h43d20405},
  {32'h44478720, 32'h438bfa60, 32'h434f67f4},
  {32'hc4c12bac, 32'h42ce739e, 32'hc304bfc4},
  {32'h4390c699, 32'h43b9ad78, 32'hc0fdb46a},
  {32'hc331c274, 32'h431bf9cc, 32'hc2abc93c},
  {32'h44b3c957, 32'h4203bc10, 32'hc31c3786},
  {32'hc46f8095, 32'hc36db4a5, 32'hc34fdf83},
  {32'h4342f6b0, 32'h43012e24, 32'h42fc4de9},
  {32'hc4c60687, 32'h4338d46e, 32'hc2bc0a83},
  {32'h444e5873, 32'hc3f1027d, 32'hc0b47ecb},
  {32'hc3e62d05, 32'hc2877872, 32'h4384dee1},
  {32'h440a21d6, 32'hc1c3aef1, 32'hc2dec79a},
  {32'hc4c5f30c, 32'hc41ddb13, 32'h421eb3bf},
  {32'h44b6f388, 32'hc39234f4, 32'h438dcb98},
  {32'hc20215ba, 32'h43b3ef2c, 32'hc35b3261},
  {32'hc2af31c4, 32'h428d9326, 32'hc33d0eed},
  {32'hc505030d, 32'hc3457079, 32'hc3035111},
  {32'h44520052, 32'hc32bd260, 32'h439923c4},
  {32'hc4754414, 32'h4294c347, 32'h427ac349},
  {32'h4500b402, 32'hc308b14f, 32'h4329a623},
  {32'hc4ccf1fc, 32'h42d08b52, 32'h412ef153},
  {32'h4463685c, 32'hc2fa87e8, 32'h43396159},
  {32'hc4465f8d, 32'hc216d9a7, 32'h428da988},
  {32'h45125248, 32'h41a75aca, 32'hc18b7c08},
  {32'hc4c9d536, 32'hc2bcc351, 32'h43e492c8},
  {32'h44b9c8ef, 32'hc2210cf0, 32'h43cb1b46},
  {32'hc40d87c0, 32'h4286a9d2, 32'hc30ad9c4},
  {32'h4484ea1e, 32'h425d2d3f, 32'hc3323921},
  {32'hc3c5fe02, 32'hc2ddec04, 32'hc21562e5},
  {32'h440fd0f6, 32'h3e966980, 32'h43626083},
  {32'hc4a3d8d8, 32'hc213cb52, 32'hc2fe0d13},
  {32'h4425f890, 32'h43f771e1, 32'hc30e0f0f},
  {32'hc4934418, 32'hbf8a3712, 32'hc318a9e7},
  {32'h45107c0c, 32'hc19fbcf8, 32'hc150af28},
  {32'hc4200539, 32'hc37ee204, 32'hc3993dac},
  {32'h44966830, 32'hc2e216b5, 32'h427c8d63},
  {32'hc45b6918, 32'h4294b940, 32'hc2a744d6},
  {32'h4489710e, 32'h4315b5e4, 32'h43a8fbef},
  {32'hc2f94900, 32'hc2a0d853, 32'hc36e35fc},
  {32'h44380551, 32'hc381819b, 32'h4394be59},
  {32'hc47ee234, 32'hc35efa9e, 32'hc34e1a13},
  {32'h448ea752, 32'h431f5e0b, 32'hc22e0940},
  {32'hc4c0ec6e, 32'h43150019, 32'h435540c3},
  {32'h44a6407a, 32'h41dd97f1, 32'h404936a0},
  {32'hc3eb5a66, 32'h43096243, 32'h44040f6a},
  {32'h44e22f25, 32'h438f3deb, 32'h43a940f2},
  {32'hc4db865d, 32'hc387ee06, 32'hc2010930},
  {32'h44519562, 32'hc289224d, 32'h438e6374},
  {32'hc45a7eef, 32'hc2042912, 32'h414599ae},
  {32'h4508a8f2, 32'h4387a1b2, 32'h432be370},
  {32'hc4a4bbd5, 32'h4285adfe, 32'h4246acfe},
  {32'h449313f6, 32'hc3e57a11, 32'hc387808d},
  {32'hc50e39bd, 32'hc274930b, 32'h43b38d2f},
  {32'h43379c90, 32'h409ce7dc, 32'hc29bb1e4},
  {32'hc513cc93, 32'h435f83d0, 32'h435cdbd2},
  {32'h443a8624, 32'h435d1bac, 32'h43a396b9},
  {32'hc50aff8c, 32'h42843bc2, 32'hbfe4bf6f},
  {32'h4487df6c, 32'h433e525b, 32'hc2cfce17},
  {32'hc4e9c5b0, 32'h42b9b62b, 32'hc3800493},
  {32'h44a556b4, 32'hc2fedf6f, 32'hc24074be},
  {32'hc2ef4d40, 32'hc1a1b2c9, 32'hc14a379a},
  {32'h4322c6f1, 32'h4163ce15, 32'hc3d6118c},
  {32'hc4bb1c62, 32'hc386a83a, 32'h43a8eead},
  {32'h448e9981, 32'h41f7e903, 32'hc388a804},
  {32'hc50d07cc, 32'hc2004dde, 32'hc2f24686},
  {32'h45123562, 32'h42dbff2c, 32'h4359a883},
  {32'hc50e4b1c, 32'hc3054dcc, 32'h425266b1},
  {32'h44ccf3e9, 32'hc332e430, 32'h42f4cf13},
  {32'hc4b30f65, 32'hc13812f3, 32'hc34bb2bf},
  {32'h452f92f2, 32'hc2c964f4, 32'h42569bb7},
  {32'hc4f53b1a, 32'h43290a0d, 32'hc2dba6a9},
  {32'h44f4a5f3, 32'hc2dcd164, 32'hc2fa3520},
  {32'hc4b4299f, 32'hc3a3cd68, 32'h43251bf2},
  {32'h4304802e, 32'h43edaacb, 32'h41e3c490},
  {32'hc450e982, 32'h433e5467, 32'hc2627095},
  {32'h449cbce0, 32'hc1131cc2, 32'h432dea93},
  {32'hc4f2b164, 32'h42b5d07f, 32'hc37e9459},
  {32'h44697040, 32'h43fd4f36, 32'h4326b2a1},
  {32'hc48535b0, 32'hc2d87a46, 32'h4376070e},
  {32'h449b8f4e, 32'h42167041, 32'h42734ac9},
  {32'hc518f90a, 32'hc24e46a1, 32'h43528200},
  {32'h44d071d2, 32'hc2023159, 32'h42c24213},
  {32'hc46c8c48, 32'hc3a137d6, 32'h42430db5},
  {32'h44dd8d7a, 32'hc3965cd1, 32'hc3e9ada2},
  {32'hc5168489, 32'hc3425d5e, 32'h4114583a},
  {32'h450aa6e4, 32'hc2f25fa4, 32'hc25d2b88},
  {32'hc3c9a34c, 32'hc231f860, 32'h42b0a1f4},
  {32'h4439d6d1, 32'h40092a4b, 32'hc28fe9bc},
  {32'hc444927c, 32'h43540ff7, 32'h432b662a},
  {32'h451f4912, 32'h438e24f6, 32'hc23654a8},
  {32'hc3eb45ce, 32'hc393c82c, 32'h42855424},
  {32'h4363f13d, 32'hc1dd9efd, 32'hc314f5ce},
  {32'hc3ae6bc5, 32'hc2209498, 32'hc34f4913},
  {32'h43a15ba4, 32'hc36de275, 32'hc40ef9a8},
  {32'hc47a9f30, 32'hc1e78521, 32'h432eada5},
  {32'h44e4401f, 32'hc34042ba, 32'hc353a721},
  {32'hc49a5685, 32'h42e80260, 32'hc22b9bd0},
  {32'h444580b4, 32'h42ba681d, 32'hc399312e},
  {32'hc503a236, 32'hc389333f, 32'hc1a9f307},
  {32'h44ce4f2a, 32'h432937f6, 32'hc306efe0},
  {32'hc4836098, 32'hc26024b6, 32'h438d8244},
  {32'h44afc817, 32'hc30c5816, 32'h422cacd5},
  {32'hc49b4406, 32'h439dcec4, 32'hc2e482f2},
  {32'hc261b740, 32'hc30b230a, 32'h42bea0b2},
  {32'hc4068e30, 32'h42995c16, 32'h43358561},
  {32'h44853b4f, 32'h42d69652, 32'hc15fa240},
  {32'h44c2e0fb, 32'hc375c00d, 32'hc33f36f7},
  {32'hc48636d6, 32'h43609e6f, 32'hc32f24c7},
  {32'h449f5852, 32'h41d2b0d1, 32'h42ec78c0},
  {32'hc4f54741, 32'hc22764f8, 32'hc37ea194},
  {32'h44fd1888, 32'h42254168, 32'hc32c131f},
  {32'hc2abb656, 32'h41d8526f, 32'h431aea2a},
  {32'h44ecb611, 32'hc3a0eee4, 32'h432bbca1},
  {32'hc483016d, 32'h4318444d, 32'hc3835019},
  {32'h4487f68c, 32'h41d2eb1a, 32'hc38351f6},
  {32'hc4e6cce6, 32'hc30448f5, 32'hc300d7f4},
  {32'h44295aa4, 32'h43a8a1b2, 32'hc32e3151},
  {32'hc49f1159, 32'hc38f77af, 32'h429936cc},
  {32'h44d80348, 32'hc273ccf8, 32'hc3ebbcb7},
  {32'hc5116cee, 32'hc366ff38, 32'hc377e37d},
  {32'h44fd7eae, 32'h440c19a6, 32'hc33a6628},
  {32'h42c27ab0, 32'hc30847a5, 32'h43f3ea6f},
  {32'h444b7432, 32'h4322cd0b, 32'hc3873cf8},
  {32'hc4f9c035, 32'hc26fac37, 32'hc2fa43bb},
  {32'h44eaa0c4, 32'h434d5b5f, 32'hc2019244},
  {32'hc460fbfc, 32'h42aac39a, 32'h4391e8e8},
  {32'h44616fcc, 32'hc380f9f4, 32'hc3c350a3},
  {32'hc507654a, 32'h4387fa94, 32'h427ebd64},
  {32'h43dcb8a8, 32'h42d5fb22, 32'hc3632a7b},
  {32'hc435a088, 32'h435bb306, 32'hc36969f8},
  {32'h44a5b132, 32'h42d747b4, 32'hc3bc2909},
  {32'hc44ac9a4, 32'h4303b356, 32'h41ef7dbc},
  {32'h44f80b20, 32'h422990d5, 32'hc193f565},
  {32'hc43d433f, 32'hc243e920, 32'hc28799d4},
  {32'h44c3cd93, 32'h431fcf97, 32'hc389803b},
  {32'hc4fda568, 32'hc2c7c1cb, 32'h43854aa5},
  {32'h44f3c2d0, 32'hc38e0d3a, 32'h435d3ff1},
  {32'hc50284d4, 32'hc385c1fd, 32'h42d713bc},
  {32'h45088b5b, 32'h42027b25, 32'h43e85bb3},
  {32'hc4ae9059, 32'h43d64fcb, 32'h42e9c5ca},
  {32'h44a31c9d, 32'hc3eac495, 32'h41086ac6},
  {32'hc3dfc9b0, 32'hc39bf112, 32'hc2040c89},
  {32'h4430d316, 32'hc21bfe2b, 32'h422953ab},
  {32'hc4e3a71a, 32'hc324185d, 32'h4312f3af},
  {32'h45057af5, 32'hc27db6ae, 32'h427f9ce6},
  {32'hc4d34146, 32'hc337ee47, 32'h4168c185},
  {32'h44d9ac1c, 32'h4347391c, 32'h430a6764},
  {32'hc40bcabc, 32'hc236e3b8, 32'h43833dfb},
  {32'h44cd03a3, 32'hc35b8872, 32'h430b2a2d},
  {32'hc3c9f6fc, 32'h41527cfe, 32'h43944cc6},
  {32'h445729c0, 32'h4333ddca, 32'h4391cf37},
  {32'hc4ee8252, 32'hc3a408ea, 32'hc3759654},
  {32'hc1acbc80, 32'hc31de631, 32'hc2cbdb41},
  {32'hc3fd2504, 32'h43c73196, 32'h438e90a8},
  {32'h42353860, 32'h42aa5b94, 32'hc33119ef},
  {32'hc4be664f, 32'hc3b2f023, 32'h42c4a048},
  {32'h4511ee70, 32'hc2f233ef, 32'hc247080b},
  {32'hc4e4fbb2, 32'h434686b9, 32'h41891062},
  {32'h4506f192, 32'hc2bae9b1, 32'h42ce15c2},
  {32'hc4cf4120, 32'hc31ae866, 32'h43083789},
  {32'h43dc75a0, 32'h42b26745, 32'hc37ea80e},
  {32'hc4aa698b, 32'h43888037, 32'hc38ced38},
  {32'h43dd0340, 32'h42ca808d, 32'h437a5281},
  {32'hc3cb0d98, 32'hc3b7ea1c, 32'hc2da6976},
  {32'hc0ad6e00, 32'hc3a519cf, 32'hc1bc7335},
  {32'hc4407ac9, 32'hc43ab57e, 32'h41a56e45},
  {32'h4481ecca, 32'hc3e5483d, 32'hc33349b3},
  {32'hc4cebb7e, 32'h4310a8c9, 32'hc305df06},
  {32'h44c9f037, 32'h43213453, 32'h439e01db},
  {32'hc38667d8, 32'hc204344b, 32'h432af3b3},
  {32'h44a354fb, 32'hc298af94, 32'h42c2b4fb},
  {32'hc44cd0a0, 32'hc2b094f2, 32'h4386e6c2},
  {32'h44bb785a, 32'hc1692d39, 32'hc39f8e4b},
  {32'h43cc5820, 32'hc346f179, 32'h41197e04},
  {32'h44056b4a, 32'hc2d892a2, 32'hc3387728},
  {32'hc3c60ff4, 32'hc333f10b, 32'hc33813ae},
  {32'h445765ae, 32'h42d3690a, 32'h42810900},
  {32'hc50c9427, 32'hc3985924, 32'h4283a80e},
  {32'h44999cf9, 32'hc335a0d1, 32'h441c303d},
  {32'hc47a97b9, 32'h423c1d88, 32'hc19fc3b9},
  {32'h441c58c5, 32'hc3efaab0, 32'hc15366e9},
  {32'hc45b930d, 32'hc24cdecf, 32'h43489c35},
  {32'h4480cd7f, 32'hc1310882, 32'h433749f8},
  {32'hc503679c, 32'hc2ca235c, 32'hc1834345},
  {32'h4466a27a, 32'hc2e285fc, 32'h437c110d},
  {32'hc4f565c2, 32'hc2620563, 32'h42d0fe83},
  {32'h42e6626c, 32'hc277f4f6, 32'h435dcff0},
  {32'hc3c85488, 32'h435fde7a, 32'hc2b4f805},
  {32'h4507f4be, 32'h431b5da5, 32'h4387670a},
  {32'hc503a8c1, 32'h422fea78, 32'h43807172},
  {32'h450a0a3a, 32'hc0a74d6e, 32'h4400bcbd},
  {32'hc376bca8, 32'hc3459b43, 32'h4235bc8e},
  {32'h44fd1df0, 32'hc334782e, 32'hc3a27c7c},
  {32'hc3fd0db0, 32'hc3384fad, 32'hc2cd4213},
  {32'h44ddcbc4, 32'hc3943c90, 32'h430acda8},
  {32'hc4c88607, 32'h42eb07c4, 32'hc36cc561},
  {32'h430b5c30, 32'hc36cd9bc, 32'h429c0234},
  {32'hc5197e7a, 32'h43933765, 32'h4300fcc3},
  {32'h44bc4fc9, 32'hc2bc79d9, 32'h434b9854},
  {32'hc48c685e, 32'hc1d4ebd0, 32'hc33ec9b8},
  {32'h44b685b5, 32'h4391c7b6, 32'h42be9b72},
  {32'hc3cfec63, 32'hc3848161, 32'h42b58831},
  {32'h446985ed, 32'h43a5117c, 32'hc3ae50e4},
  {32'hc5138669, 32'h42e4cca2, 32'hc3951233},
  {32'h44088ee2, 32'hc329289c, 32'h4102444c},
  {32'hc509cf20, 32'h41d32096, 32'h43ce6b4e},
  {32'h4513fde0, 32'h42ad495b, 32'hc3d2aef3},
  {32'hc4d61f07, 32'h42b681cf, 32'hc28ef02f},
  {32'h450390af, 32'h40a20f26, 32'h433f387c},
  {32'hc43c33cf, 32'h431dd07a, 32'h432ddd49},
  {32'h44484de9, 32'hc2ed9fcd, 32'hc3833220},
  {32'hc1155500, 32'h423b1ab0, 32'hc30666fd},
  {32'h45143721, 32'hc3a0ef83, 32'h438348f2},
  {32'hc454adc4, 32'hc180e221, 32'h42869151},
  {32'h4514e7fe, 32'h4321d162, 32'hc3632084},
  {32'hc3ac785c, 32'h42817834, 32'hc1981466},
  {32'h4503dcfc, 32'hc1d1808c, 32'hc1e17c1e},
  {32'hc410ceaf, 32'h44140fae, 32'hc3890756},
  {32'h44aa98ff, 32'hc3949f1e, 32'h42a7e4f0},
  {32'hc4d9dbbb, 32'hc32536c9, 32'hc3ad7f64},
  {32'h43f67422, 32'h42e9b90a, 32'h41fea7dc},
  {32'hc50900c2, 32'hc21914fa, 32'h42414215},
  {32'h44650ce0, 32'h3f0a1580, 32'h42bb9054},
  {32'hc413fb1e, 32'hc3a13a68, 32'h43b655a8},
  {32'h4510cbd2, 32'hc3256d6b, 32'h420a4616},
  {32'hc5120877, 32'hc385cbeb, 32'h438f3de4},
  {32'h44da921b, 32'h440562d6, 32'hc3801192},
  {32'hc49575c1, 32'h4366f8cc, 32'h43acc8c5},
  {32'h44c3b0b3, 32'h41157fd1, 32'hc2b1818c},
  {32'hc450cc34, 32'hc2762567, 32'hc24d2f1b},
  {32'h4502fc6c, 32'h426ab3b8, 32'hc31bd82f},
  {32'hc1c84760, 32'hc3631b5e, 32'h43925182},
  {32'h44c77cd7, 32'hc3828e7d, 32'hc27b7564},
  {32'hc3ad2084, 32'h43966bac, 32'h434c1049},
  {32'h4513e193, 32'hc34121e6, 32'hc35c7f08},
  {32'hc4e2ed25, 32'hc30ed832, 32'h437a8189},
  {32'h45050ebc, 32'h4389ec16, 32'h42f83a42},
  {32'hc4028d9a, 32'hc2e6831e, 32'hc24788ad},
  {32'hc2f520a0, 32'hc33cc7ee, 32'h43c2bc0b},
  {32'hc505b256, 32'h43d7742a, 32'h42f2a3ac},
  {32'h4431c0c2, 32'h42fd93a8, 32'h43d96688},
  {32'hc364bfc8, 32'h40da852c, 32'h4289a4ac},
  {32'h44a1bcf6, 32'hc3079ae6, 32'hc2416e0c},
  {32'hc4ec0a61, 32'hc382c39b, 32'hc36d346b},
  {32'h450e5a90, 32'hc2e8b1ce, 32'h4110b998},
  {32'h4274a6c0, 32'h4324b24d, 32'hc379cf01},
  {32'h44f899cf, 32'h42ee9eea, 32'hc2b3b739},
  {32'hc2dc77e9, 32'hc3b3c004, 32'h431ad4b5},
  {32'h44ef1390, 32'hc3883b38, 32'h41d2ac0a},
  {32'hc4cfe163, 32'hc38aecc1, 32'h4370c011},
  {32'h4501fcc3, 32'hc34f19ea, 32'h4394d89c},
  {32'hc4fb9ff6, 32'hc2f39b71, 32'hc367e617},
  {32'h43ad8feb, 32'hc3ba1a06, 32'hc3001fe5},
  {32'hc4c7bd40, 32'hc3450084, 32'h4360674c},
  {32'h450430db, 32'h42f5b530, 32'h42318a79},
  {32'hc4de59ee, 32'h4358cf68, 32'h4359a928},
  {32'h44e01919, 32'hc344ecee, 32'hc16b76b4},
  {32'hc48844bc, 32'hc390c890, 32'h424b0f6d},
  {32'h44fd99de, 32'h432f4f18, 32'h440f5aea},
  {32'hc4e1039b, 32'h4352d382, 32'hc246fafb},
  {32'h444b83df, 32'hc38f6ba4, 32'hc380c147},
  {32'hc4e29f6f, 32'h438aea77, 32'h42eb90bb},
  {32'h446af42c, 32'hc340949e, 32'h41517cbe},
  {32'hc4b281db, 32'h43847808, 32'h41b98b73},
  {32'h4476aa02, 32'h4254cb83, 32'hc38632ee},
  {32'hc4d5ac1d, 32'h43046504, 32'h437a82d3},
  {32'h4500fe8b, 32'h43639704, 32'h43c5db09},
  {32'hc4187bd2, 32'hc38d2a83, 32'h41523bbb},
  {32'h44cb60f1, 32'hc30660f9, 32'hc2a362ff},
  {32'h3f96fc00, 32'h42b15cc9, 32'hc385f79d},
  {32'h4425e0aa, 32'hc211e071, 32'hc380db5f},
  {32'hc48abe2a, 32'hc1ddf472, 32'h42c71b54},
  {32'h44f9fa79, 32'h43324d17, 32'hc38fcd7e},
  {32'hc4b725ce, 32'h43847939, 32'hc3533a2a},
  {32'h44de7254, 32'h43ad3152, 32'h42a7090b},
  {32'h4267a3c7, 32'h432a27c1, 32'h42e5bf09},
  {32'h4437ed25, 32'h42796e0a, 32'hc2d36ef8},
  {32'h437deeb0, 32'hc1f0a8f6, 32'h442a614b},
  {32'h4431f5dc, 32'hc360d4e7, 32'h42dbca33},
  {32'hc40bac48, 32'hc2f0ba01, 32'h43859c71},
  {32'h44b77857, 32'hc25e2632, 32'h422cf688},
  {32'hc481aec8, 32'hc2b56ed6, 32'hc33cbed3},
  {32'h43e7bd70, 32'hc16aa969, 32'hc22eefab},
  {32'hc473be78, 32'hc34c5956, 32'hc291d62a},
  {32'h4424a770, 32'hc3984efe, 32'h42c06a09},
  {32'hc4412db8, 32'h4240347a, 32'hc3a0da9b},
  {32'h44b30f24, 32'hc2c1fcbe, 32'hc1fc1651},
  {32'hc488eeee, 32'h419ea88a, 32'hc381fa3d},
  {32'h44a2b26f, 32'h402d01c6, 32'h445f4450},
  {32'hc3cc3360, 32'h43c44f86, 32'h42df128f},
  {32'h449bc170, 32'hc3970060, 32'hc300900f},
  {32'hc4c849d0, 32'h431285e1, 32'h42b37b40},
  {32'h450435d2, 32'hc30ba094, 32'hc330560f},
  {32'hc4031d3d, 32'h43c54eeb, 32'h430b5daf},
  {32'h44f0f88a, 32'hc3db2752, 32'h427b75bc},
  {32'hc4d02797, 32'hc2a86048, 32'h4354ef16},
  {32'h440b03e2, 32'h4116c9d1, 32'hc376a9b0},
  {32'hc42443e8, 32'h4395dd72, 32'h42ed41cd},
  {32'h445beb53, 32'hc312d35d, 32'h4204c760},
  {32'hc4068419, 32'h42fb083d, 32'h42b6c5b3},
  {32'h44ca25a9, 32'hc2c24e5c, 32'h429b7e41},
  {32'hc485be24, 32'h42cf70f1, 32'h42c32bf0},
  {32'h45190297, 32'hc3a22e1c, 32'h430133ee},
  {32'hc4f709ae, 32'hc213d2de, 32'h42d1864f},
  {32'h44aaf4ca, 32'hc3017290, 32'h42a3144b},
  {32'hc4a0cc3e, 32'hc39d06d0, 32'h42eeed6b},
  {32'h44c79ba2, 32'hc38e7d6e, 32'h4371b114},
  {32'h42cce510, 32'h42930774, 32'h42e64b60},
  {32'h4482a5e8, 32'hc345b06f, 32'hc23868c7},
  {32'hc4e2c07c, 32'hc03d0d4a, 32'h439d750a},
  {32'h43ab022c, 32'h4390bcf0, 32'hc1133253},
  {32'hc4cf2be6, 32'h431c378c, 32'h4407d85e},
  {32'h443fc0c4, 32'h438cd2e6, 32'h43a016d0},
  {32'hc4911bb2, 32'hc30a8423, 32'hc41bb988},
  {32'h4447576c, 32'hc3b85df1, 32'h41245cc3},
  {32'hc505759a, 32'hc3238fc8, 32'h3fe16fbe},
  {32'h44d159a3, 32'hc228ddbe, 32'hc316ef50},
  {32'hc42fa6d7, 32'hc2fe11e5, 32'h43547f34},
  {32'h44a3006e, 32'h439a9794, 32'hc2b709da},
  {32'hc514e170, 32'h41cd6fd2, 32'hc3952700},
  {32'h451039c1, 32'h41eb41a1, 32'h42836a90},
  {32'h42843c40, 32'hc36bba1f, 32'h434417ca},
  {32'h4473f43a, 32'h432acfc6, 32'hc1e90a5c},
  {32'hc4c37636, 32'h43400f4c, 32'h42fe3d8e},
  {32'h4429a64c, 32'hc20e8055, 32'h42d91685},
  {32'hc4747b02, 32'h430bde66, 32'hc28e8d81},
  {32'h441aa62c, 32'hc206bf26, 32'hc2c4c43d},
  {32'hc4fc600b, 32'h41828a6a, 32'hc370cb51},
  {32'h445131d0, 32'h43377890, 32'hc2af0548},
  {32'hc4649356, 32'h43266244, 32'hc2a64c12},
  {32'hc2268d50, 32'h42935111, 32'hc2c04962},
  {32'hc5193284, 32'hc2d79dd7, 32'h42873d16},
  {32'h45123552, 32'h43e82c2b, 32'h432425ea},
  {32'hc46b12fd, 32'hc2be11f3, 32'hc304ab7b},
  {32'h44b48287, 32'h439ed14a, 32'hc234ee72},
  {32'hc4b9f25d, 32'hc1f9be24, 32'h411cddc6},
  {32'h449b847e, 32'h42d83d5f, 32'h4288d917},
  {32'hc3855fd6, 32'h42436119, 32'h42b6623d},
  {32'h44c77249, 32'hc2cf7414, 32'h4326e343},
  {32'hc35c95e0, 32'hc2ab6682, 32'hc2e87b13},
  {32'h43e0ab98, 32'hbf9a66b0, 32'hc2f11e51},
  {32'h42089940, 32'hc39f56e7, 32'h41fd482e},
  {32'hc2310600, 32'h431d98e1, 32'h435188c7},
  {32'hc43cc0a8, 32'h435c638e, 32'h4123106d},
  {32'h43f1ffaf, 32'hc2a3486d, 32'hc3193ee5},
  {32'h429e5a40, 32'hc30e9a84, 32'hc30e4533},
  {32'h448ce6c9, 32'hc387cb2b, 32'hc2f00d63},
  {32'hc5013e1e, 32'h435dd70d, 32'hc3081291},
  {32'h44113b68, 32'hc28f4b9c, 32'h434fa29f},
  {32'hc4062819, 32'h42d907b8, 32'hc2b0daf1},
  {32'h449fac3b, 32'h43c2a014, 32'h434d447c},
  {32'hc496612b, 32'hc306cbec, 32'h437b2610},
  {32'h448da9d8, 32'hc38007fc, 32'hc20d07f1},
  {32'hc4e7329f, 32'hc36a9429, 32'h432ec7b9},
  {32'h44b00824, 32'h43bc90ab, 32'h43f1c2be},
  {32'hc4f5e833, 32'hc2d72b48, 32'hc3027c48},
  {32'h447b7b50, 32'h43aee482, 32'h42d2ef76},
  {32'hc49dbea9, 32'h430fe05a, 32'hc3ceaa78},
  {32'h44f59971, 32'hc3d26925, 32'h4304ae74},
  {32'hc4c3047b, 32'hc36d2993, 32'h427a61d0},
  {32'h44d39970, 32'hbd772900, 32'hc3cac02f},
  {32'hc42ee970, 32'hc3c4ca22, 32'h43d628e8},
  {32'h43689cb2, 32'hc40c254e, 32'h42a0036a},
  {32'hc46875a3, 32'hc3ac5f86, 32'hc36ca732},
  {32'h450b9232, 32'hc2aa2a00, 32'hc37def0e},
  {32'hc3a366db, 32'hc2aa604c, 32'h43c7422f},
  {32'h4346f1ac, 32'h439a2a59, 32'h43000b9e},
  {32'hc4887695, 32'h423b3565, 32'hc28aa614},
  {32'h44a79c41, 32'h42746f69, 32'hc35ac759},
  {32'hc4b92ba8, 32'h42b042fe, 32'hc30eb040},
  {32'h44e04f2b, 32'h418dca18, 32'hc12d6b17},
  {32'hc4b20883, 32'h43a20eda, 32'hc3b37b40},
  {32'h43dc66e8, 32'h439dd0d5, 32'hc2b96317},
  {32'hc39974d2, 32'h440710ae, 32'hc2264b96},
  {32'h42da5460, 32'h433a3a14, 32'h43804a47},
  {32'hc4a8df7a, 32'hc3dbac48, 32'hc31c2b75},
  {32'h43a99100, 32'hc1938562, 32'hc2b9779e},
  {32'hc3c71178, 32'hc13ed6ae, 32'hc2826b32},
  {32'h447ed4ac, 32'h42a7fb7a, 32'hc3558380},
  {32'hc4a9218e, 32'hc367f34c, 32'hc0db5e26},
  {32'h43ff2dfc, 32'hc3b87858, 32'hc2e9b1e8},
  {32'h4240fb00, 32'hc3530492, 32'h431eaedf},
  {32'h44d73946, 32'h42d56bed, 32'h43862390},
  {32'hc49f1c8d, 32'h417e4582, 32'h43d9746d},
  {32'h4495e191, 32'h4373867a, 32'h41dd8ed2},
  {32'hc3add824, 32'hc3b826d8, 32'hc365bf19},
  {32'h448010e4, 32'hc35e0ad0, 32'hc2d901fa},
  {32'hc4495974, 32'h43116f92, 32'h4266186c},
  {32'h43f0ab60, 32'hc20e2c63, 32'hc38d28d8},
  {32'hc3b6a2d6, 32'h41ae7d5f, 32'h42dcff27},
  {32'h450dd250, 32'h43dff45e, 32'h4222cc2e},
  {32'hc45732c8, 32'h41eed3b0, 32'h42a798d0},
  {32'h43848dd0, 32'hc24a028b, 32'h42e46287},
  {32'hc4a07494, 32'hc1fc364e, 32'h435b1aca},
  {32'h449df142, 32'hc2be9395, 32'hc2cc45fe},
  {32'hc4d8d403, 32'h43864bc4, 32'hc3a8b702},
  {32'h44fa3b3f, 32'hc3f48aa3, 32'hc3b9f0d9},
  {32'hc4d8b0c4, 32'h42efe110, 32'h42ab6f14},
  {32'h44bcccae, 32'hc27b3878, 32'h41d2e9cd},
  {32'hc48b9142, 32'h4309f335, 32'hc294e7dc},
  {32'hc259c0e0, 32'hc3d368b9, 32'h437975b9},
  {32'hc3cba70c, 32'h3fe67754, 32'h41d0efee},
  {32'h45008da9, 32'h3f1cabbb, 32'h432ccd4f},
  {32'hc49bc512, 32'h4399dde8, 32'h42d8bc54},
  {32'h44842074, 32'h43e38ad3, 32'h43a0c1c8},
  {32'hc4bfa898, 32'hc397e356, 32'hc39479a6},
  {32'h43369868, 32'h43bfea15, 32'hc3bec0fe},
  {32'hc49896b2, 32'hc3b95890, 32'h416787d6},
  {32'h44d855b2, 32'hc2aa13fd, 32'hc2a2bdca},
  {32'hc4a54db9, 32'h43159fe0, 32'h4037c759},
  {32'h44af6e85, 32'hc31e6dfa, 32'hc3803703},
  {32'hc4050267, 32'hc2369a4a, 32'h429d10f4},
  {32'h4507fcfc, 32'h43b57c02, 32'hc18e3b54},
  {32'hc49aeb40, 32'h42d56994, 32'h40f39d9b},
  {32'h45127c14, 32'h432d1f32, 32'hc26bae9a},
  {32'hc4a54b1a, 32'h43164b12, 32'h43bccb09},
  {32'h4493d2ce, 32'hc3be2015, 32'h432f45b2},
  {32'hc4032530, 32'h42e97316, 32'h434c75c3},
  {32'h44122100, 32'h420b698b, 32'hc211ee40},
  {32'hc50daa78, 32'hc28bd08d, 32'hc3471cf2},
  {32'h44bbdd5d, 32'h4324c234, 32'hc3337498},
  {32'hc46334e8, 32'hc1caae5e, 32'hc3b0f8b3},
  {32'h441198c8, 32'h42aee880, 32'hc2ddfa2d},
  {32'hc4fe9474, 32'h435c242c, 32'h442af31c},
  {32'h448d141e, 32'h43e87503, 32'hc3fe7c66},
  {32'hc464ccb4, 32'hc282d22f, 32'h4323105a},
  {32'h44a81f0a, 32'h43794e30, 32'hc100645c},
  {32'hc4b6cc27, 32'h43739c57, 32'hc2103f5b},
  {32'h440aa6d4, 32'h439aac04, 32'hc32fb658},
  {32'hc48a417c, 32'h43ca4171, 32'h44072f46},
  {32'h446091ec, 32'hc1559def, 32'h433acdc8},
  {32'h42852780, 32'h437a3136, 32'h437c2ae4},
  {32'h44fb6fa2, 32'hc31b88e3, 32'hc3352d08},
  {32'hc4052dee, 32'h436a062d, 32'h43786ee7},
  {32'h44ae55c8, 32'hc302e59a, 32'h420c1b2a},
  {32'hc5070d80, 32'hc33c43f3, 32'h42ca4031},
  {32'h43e2e021, 32'h42f313eb, 32'hc28fa393},
  {32'hc4bb9a2c, 32'h4379c3c2, 32'h43a213b4},
  {32'h445eb00a, 32'hc343d1a2, 32'hc43b4e81},
  {32'hc4c4024a, 32'h438a51d4, 32'hc2ec1361},
  {32'h451d0302, 32'hc22d6726, 32'h43bcce86},
  {32'h42435f00, 32'hc2f5b9ae, 32'hc2d6187e},
  {32'h44dc1229, 32'hc3969b7e, 32'hc3875b59},
  {32'hc504076e, 32'hc263018e, 32'hc3d3ffdc},
  {32'h4406dc7a, 32'h42836c6c, 32'hc348a2ac},
  {32'hc4cc5e2c, 32'h43ada36e, 32'h43545816},
  {32'h4492cedb, 32'h437f7e1a, 32'hc09c60ea},
  {32'hc47c5b00, 32'h441766c2, 32'hc3bc9a88},
  {32'h450c93bc, 32'h43860f8c, 32'h4350a426},
  {32'hc42c54e4, 32'hc2273e63, 32'hc322ced0},
  {32'h43e3474c, 32'h43c28174, 32'hc31c5d25},
  {32'hc518f56a, 32'h42c9b282, 32'h43b3f8f9},
  {32'h4506e2b9, 32'h42b11cc8, 32'h426f679a},
  {32'hc4a21b06, 32'hc273d62d, 32'h43f7ecfd},
  {32'h44bcc389, 32'hc2cfbe47, 32'h40fe03c2},
  {32'hc4d4670e, 32'hc1afd410, 32'hc28c1465},
  {32'h44ed92c3, 32'hc3502abf, 32'h419a0cc5},
  {32'hc49beb2e, 32'hc3092d94, 32'hc3bdae14},
  {32'h44878e2e, 32'hc37c5d52, 32'h42ad874f},
  {32'hc437d254, 32'hc3ca762b, 32'h4227b5be},
  {32'h452c748c, 32'hc4046cc7, 32'hc254c258},
  {32'hc50e1232, 32'h42b995fe, 32'hc36fdd2e},
  {32'h45135399, 32'hc3aea735, 32'hc117034d},
  {32'hc5173ce8, 32'h42fb138c, 32'hc0429b4d},
  {32'h44b226ee, 32'h4364e433, 32'hc19c63b7},
  {32'hc492ef40, 32'hc4107294, 32'hc3324705},
  {32'h44059aa0, 32'hc318cd3b, 32'hc2e0ef28},
  {32'hc3d92385, 32'h436d32db, 32'hc242137a},
  {32'h423d2680, 32'h42a435c3, 32'h433e27a7},
  {32'hc4b58bd6, 32'h434b04a8, 32'h4295c108},
  {32'h448c85e8, 32'hc3b6d2b7, 32'hc318cd11},
  {32'hc4b0289d, 32'h42d6a5b9, 32'h4263fd34},
  {32'h432d8800, 32'h438e21c1, 32'hc2a74186},
  {32'hc4dd53a0, 32'h4334870c, 32'hc29681e5},
  {32'h44010780, 32'h430c90a2, 32'h438f4db0},
  {32'hc4de431a, 32'h4388dd65, 32'hc2d08296},
  {32'h44cc82f8, 32'h42bbb650, 32'hc380d64a},
  {32'hc45ed310, 32'h42eafb58, 32'h418c5663},
  {32'h43a42f66, 32'h42b1ac54, 32'hc38355fb},
  {32'hc51de0e7, 32'h433b121b, 32'hc2a4ac43},
  {32'h44ee1cb8, 32'h439d8980, 32'hc1dd1454},
  {32'hc378864c, 32'hc27a8ebb, 32'hc3299015},
  {32'h4513e4bc, 32'hc392bada, 32'h42a0f609},
  {32'hc50d8194, 32'h43880776, 32'h43649114},
  {32'h42b930c0, 32'hc3b42d1e, 32'hc26bf0a9},
  {32'hc4bc35eb, 32'hbecc2c00, 32'h43832b16},
  {32'h4505a4e3, 32'h43df5e3a, 32'h430251ff},
  {32'hc31ec61e, 32'h42c9a880, 32'hc2b1e3dc},
  {32'h44fe810b, 32'h422dfa42, 32'hc344bd89},
  {32'hc37ce0b4, 32'hc373448b, 32'hc36980b7},
  {32'h44f1d59e, 32'hc2fcd774, 32'h4316e849},
  {32'h42a18977, 32'h42b4cb66, 32'h433a0955},
  {32'hc259afbc, 32'h42e963c5, 32'h4322d88f},
  {32'hc364ee5d, 32'hc4043649, 32'h42e3806d},
  {32'h441324a1, 32'hc264b44e, 32'h41e35062},
  {32'hc3a1b49b, 32'hc3cabb90, 32'hc34b17e7},
  {32'h450f0c0a, 32'h433746be, 32'hc377b386},
  {32'hc3a008f0, 32'hc3aa008d, 32'hc1f515cd},
  {32'h447a9888, 32'h43b3cc2b, 32'hc2b48e93},
  {32'hc50aa5fa, 32'hc1f32d08, 32'hc391a677},
  {32'h451fd22b, 32'hc21eec00, 32'hc2af32ef},
  {32'hc3a9e920, 32'hc38ae612, 32'hc3abeb3d},
  {32'h438f2910, 32'hc28e02b0, 32'h4317361a},
  {32'hc49c1a60, 32'h43e32711, 32'h4373353f},
  {32'h4488b98b, 32'hc3f473ca, 32'h42f69c49},
  {32'hc4c46ad7, 32'h43ad278e, 32'h4284b289},
  {32'h43f6df28, 32'h42542449, 32'h43794201},
  {32'hc4100993, 32'h432602e4, 32'hc341b591},
  {32'h440713c0, 32'h4294a08e, 32'h433e3a6a},
  {32'hc4c1ea37, 32'hc3193792, 32'hc2f0b81b},
  {32'h44809ba2, 32'hc2762124, 32'h41fa7a2a},
  {32'hc4eb99f0, 32'h41a63e7f, 32'hc3550b35},
  {32'hc2e317a0, 32'h44034574, 32'hc39dd98b},
  {32'hc4a8ca95, 32'hc3606404, 32'hc3bc924e},
  {32'h44b9a7cc, 32'h4379acaa, 32'h43da4784},
  {32'hc4898844, 32'hc33d0dbc, 32'hc38c6a61},
  {32'h44c1af8b, 32'h43d9f021, 32'h432c6915},
  {32'hc43654e0, 32'h425a2af8, 32'hc2ec82aa},
  {32'h44cdc706, 32'h43dfdd24, 32'hc3e75388},
  {32'hc2885b80, 32'hc3b01882, 32'hc31735f2},
  {32'h4508fc50, 32'hc273d7d1, 32'hc2390c2e},
  {32'hc4d77000, 32'hc31cf641, 32'h40d0d9b4},
  {32'h44bfa27d, 32'hc2d1c81a, 32'h4360d2c5},
  {32'hc44e35c8, 32'hc0f8d166, 32'hc3ba0d7f},
  {32'h4496ee16, 32'h42d2d673, 32'hc213011c},
  {32'hc3838350, 32'h42aed890, 32'hc34f6572},
  {32'h4499252c, 32'hc32f3e0f, 32'h4414ee5a},
  {32'hc31db2a8, 32'h43770a17, 32'hc36091d2},
  {32'h4523b164, 32'hc3a10e31, 32'h4279703f},
  {32'h4368b830, 32'hc306cd2a, 32'h43a175b5},
  {32'h43ba0fa6, 32'h4238a46a, 32'h43ca09ff},
  {32'hc4f379cc, 32'h428160e7, 32'hc31475d9},
  {32'h44c9540e, 32'h43cf51ab, 32'h425cfc53},
  {32'hc42014d9, 32'h416b7dde, 32'h423a3094},
  {32'h4502d10f, 32'hc3e6c7b5, 32'hc32fb5d1},
  {32'hc464a5c0, 32'hc372e95a, 32'hc3987fad},
  {32'h4460b7e4, 32'h43d921cc, 32'h43aa1d96},
  {32'hc4541ce5, 32'h4281cf4e, 32'h42cfa058},
  {32'hc50bfbfa, 32'hc2f006f6, 32'h4358742f},
  {32'h43ef6577, 32'hc3dfe0e7, 32'h42f6047f},
  {32'hc50d557f, 32'hc387a1ed, 32'hc34a1b92},
  {32'h4503123c, 32'h42c68597, 32'h42c9125e},
  {32'h42ab671a, 32'hc3b4e942, 32'h42d2d2b1},
  {32'h43c26790, 32'h42eea43b, 32'h4317352d},
  {32'hc206cf60, 32'hc3b4ab2c, 32'hc3b43460},
  {32'h44fe3ecb, 32'hc3288b5c, 32'h4390ae97},
  {32'hc5020699, 32'h433ff4c7, 32'h42e5ca28},
  {32'h44fb2eea, 32'hc32c2b9d, 32'hc1564035},
  {32'hc4cf205d, 32'hc31bf5d5, 32'h4293426d},
  {32'h43d90aba, 32'hc217eeab, 32'h436351a2},
  {32'hc4ce3a24, 32'h4304cc40, 32'h4354ac79},
  {32'h44075ac2, 32'hc2452d8b, 32'hc34d5eb5},
  {32'hc4945efd, 32'hc3815f3a, 32'hc4081d28},
  {32'h4514b47d, 32'h43fa305e, 32'hc10f8451},
  {32'hc4f26a6a, 32'h42f59d3e, 32'h439995a8},
  {32'h44bb2772, 32'hc3387f8c, 32'h4372d5a6},
  {32'h42652272, 32'h430545a2, 32'h4273fec5},
  {32'h44b7df53, 32'h42213480, 32'h43e6a621},
  {32'hc415c0da, 32'h43515bba, 32'hc2b2c058},
  {32'h44b1dd50, 32'hc3121aa2, 32'h437929de},
  {32'hc47edf68, 32'hc2b7dc49, 32'hc39189aa},
  {32'h44915ae7, 32'h4261daf4, 32'h437a74e9},
  {32'hc3e0dca8, 32'h43a55d53, 32'hc182926c},
  {32'h44f2ab41, 32'hc2c03aea, 32'hc387a5b7},
  {32'hc4c12a7b, 32'h43130224, 32'h43902a75},
  {32'h43af439c, 32'h435b6adc, 32'h418522a2},
  {32'h43ab3910, 32'hc381af06, 32'hc3a6f968},
  {32'h432ddfd8, 32'h42973848, 32'h42ab2ada},
  {32'hc42546bd, 32'h414db90c, 32'hc38f667c},
  {32'h449b7962, 32'hc29bd639, 32'h4308cc7b},
  {32'hc43fc2a8, 32'hc2753bf8, 32'hc3704f5d},
  {32'h44ebbe59, 32'h42aa45a1, 32'h42806071},
  {32'hc399da50, 32'h438af3ca, 32'hc31fe7c6},
  {32'h441101d0, 32'h422f02b4, 32'h4200920b},
  {32'hc4d73c44, 32'h419e3e9f, 32'h4361ba75},
  {32'h4480cb6e, 32'h40f0ec22, 32'h44198f84},
  {32'hc40de370, 32'hc2cbc02c, 32'h42a8caf8},
  {32'h445c083e, 32'hc38c6e8a, 32'h4240b431},
  {32'hc38b2998, 32'h436256dc, 32'h4374995a},
  {32'h44aba137, 32'hc344e0ff, 32'hc2eeaae3},
  {32'hc4900575, 32'hc262a145, 32'h43691fd6},
  {32'h44ff25fd, 32'h43648cf5, 32'h42946b88},
  {32'hc500c5ff, 32'hc3ad11ce, 32'hc32bd78a},
  {32'h44829e99, 32'h422073d0, 32'h437c1595},
  {32'hc41b55c2, 32'h435a5b54, 32'hc3349f16},
  {32'h432b482a, 32'h414894de, 32'hc3869871},
  {32'hc4e4e7ad, 32'hc301f6d1, 32'hc253be46},
  {32'h451187b2, 32'h420e67ca, 32'h423fcea4},
  {32'hc4d79bc0, 32'h42e178f2, 32'h3f77e3a0},
  {32'h4507087d, 32'h423fccf9, 32'hc224acf4},
  {32'hc4d62b87, 32'h4238aba4, 32'h42d19768},
  {32'h450956d6, 32'h43bcc74e, 32'hc256d3d6},
  {32'hc509d53f, 32'hc38bcf01, 32'h42f0ab34},
  {32'h43d542ab, 32'hc2dec0c4, 32'hc2e1cacf},
  {32'hc4d578ba, 32'h4355efea, 32'hc390153d},
  {32'h4511aaac, 32'h436c80e2, 32'h4270b8d0},
  {32'hc340e4f0, 32'h4298b4fc, 32'h42f22d6d},
  {32'h450910ff, 32'h433889f0, 32'h428d3e3e},
  {32'hc4711568, 32'h420f148f, 32'h4252919c},
  {32'h44a97de9, 32'hc219d000, 32'h43835fa9},
  {32'hc4df65d5, 32'h4281ba3b, 32'hc2fd1ca8},
  {32'hc2c1b250, 32'hc2402e68, 32'h43976668},
  {32'hc4a19933, 32'h42bf7dcf, 32'h4406f366},
  {32'h45153163, 32'hc38cda5c, 32'hc22c634d},
  {32'hc50dea37, 32'h422da572, 32'hc294bb3c},
  {32'h447f8d5a, 32'hc30c995f, 32'hc3155944},
  {32'hc4bc4db7, 32'h43664a64, 32'hc20a1428},
  {32'h44d5f8c7, 32'hc358caee, 32'hc2f07915},
  {32'hc439a858, 32'h438c1ae6, 32'hc379ec37},
  {32'h443ffe84, 32'hc2f0426c, 32'h4396e613},
  {32'hc4854377, 32'h4371ea22, 32'h4402a8f7},
  {32'h44050df8, 32'h423aa5e2, 32'hc340e025},
  {32'hc4305838, 32'h417bd37c, 32'h433aec73},
  {32'hc2ab3cc0, 32'h43faed77, 32'h4298c0ed},
  {32'hc39a5cec, 32'hc2b8aa31, 32'hc30e4496},
  {32'h446e9cbc, 32'h437551e6, 32'hc39f5a54},
  {32'h430cac00, 32'h43a17ae4, 32'h43aa57ec},
  {32'h44c38bb6, 32'h42ed3693, 32'h43ad21b8},
  {32'hc51485cf, 32'h425bcfae, 32'h42f3b886},
  {32'h44b83de3, 32'h435a1376, 32'hc3007b55},
  {32'hc50ac235, 32'h430e3243, 32'hc38d8059},
  {32'h4492da4f, 32'hc40c9d4b, 32'hc38222d1},
  {32'hc41c1ff8, 32'hc3a77729, 32'hc31c5fed},
  {32'h44f917fb, 32'hc2941009, 32'hc367e25e},
  {32'h422373d0, 32'hc3623431, 32'hc111ec70},
  {32'h44c99d4c, 32'h436ab893, 32'hc2008ed0},
  {32'hc33ab880, 32'h4325f93d, 32'h4308bb1e},
  {32'h45061794, 32'h43384d0f, 32'h42ce74a2},
  {32'hc3d70762, 32'hc3e6669a, 32'hc2439d9a},
  {32'h435aaf48, 32'hbedc32a0, 32'h438b7099},
  {32'hc4c9c5a3, 32'hc3a345e4, 32'hc2a83133},
  {32'h44470fa6, 32'h433416dd, 32'hc2824e61},
  {32'h417f6238, 32'hc306df63, 32'h438d2e78},
  {32'h444d46ae, 32'hc2bd4248, 32'hc38b84e8},
  {32'hc4819964, 32'h4317caff, 32'h43adb350},
  {32'h44c88008, 32'hc3af9fbc, 32'hc31f19fb},
  {32'hc48635d4, 32'h443613a4, 32'hc095d56e},
  {32'h441911cc, 32'hc3a5a830, 32'h437d0587},
  {32'hc4fbf782, 32'hc1480509, 32'h433298f3},
  {32'h43f90396, 32'h43929852, 32'h435a003b},
  {32'h43403ac6, 32'h4311055a, 32'h43299ea7},
  {32'h450305a7, 32'hc1cfaf2b, 32'h429f3bd6},
  {32'hc4a0f70f, 32'h43f8b84b, 32'hc2e796ca},
  {32'h44d52b0c, 32'hc2c44d42, 32'h43316df6},
  {32'hc3f95519, 32'hc3973fea, 32'hc34dd631},
  {32'h44bac36d, 32'hc19f7c52, 32'hc317ffa1},
  {32'hc49cc13a, 32'hc2dadd9e, 32'h43041fb4},
  {32'h451399fd, 32'h435de9aa, 32'h43f74a01},
  {32'hc43bb2f4, 32'h434eb706, 32'h4261e0ca},
  {32'h4486eefc, 32'h430a72e9, 32'h438074e4},
  {32'hc451f032, 32'h43751ad8, 32'h44115e87},
  {32'h4388c560, 32'h427ed9a4, 32'h4342648f},
  {32'hc4f370d7, 32'h43a5b9c8, 32'h43ff3ab1},
  {32'h445d3424, 32'hc3111a26, 32'hc3c6e140},
  {32'hc3f6bceb, 32'h429cd2e7, 32'h42cf83b3},
  {32'hc31f58a4, 32'hc2d363c2, 32'hc2f00f04},
  {32'hc5014463, 32'hc1a1d296, 32'h433ce2c7},
  {32'h44493d8c, 32'hc21dd8a6, 32'hc31e9778},
  {32'hc49a5b97, 32'h43a98200, 32'hc29d24c2},
  {32'h44dc7b61, 32'hc33c8e0f, 32'hc38f475b},
  {32'hc4f61e35, 32'hc3bfd963, 32'hc1221d67},
  {32'h442901d8, 32'hc33f383c, 32'h43014542},
  {32'hc441b798, 32'hbf735740, 32'h43c57fdb},
  {32'h44ffcd2f, 32'h40ca65fd, 32'h42252740},
  {32'hc5043d60, 32'hc168fa09, 32'h42f6ec8d},
  {32'h43f59818, 32'h43b29a9b, 32'hc3167946},
  {32'hc3f07c30, 32'h43b96457, 32'hc3b77cb8},
  {32'h45073da3, 32'h432940cb, 32'hc34291b9},
  {32'hc450c11e, 32'h435624ab, 32'hc3bdc645},
  {32'h44a0547c, 32'h4203f57c, 32'h43a6db2b},
  {32'hc390d6a1, 32'h4286d53d, 32'h42d6a5f1},
  {32'h44b6bd4d, 32'hc3082a52, 32'h42f1067f},
  {32'hc465885b, 32'h42c8ab43, 32'h4369d198},
  {32'h444360ec, 32'h42aea698, 32'hc3bdb005},
  {32'hc42869cd, 32'h43a12851, 32'h4366217e},
  {32'h43ca35e0, 32'hc33641df, 32'h439cfdae},
  {32'hc3075190, 32'h43d02ef9, 32'hc388b47a},
  {32'h44b51c6c, 32'hc3ba110b, 32'h4363aa7b},
  {32'hc404e669, 32'h431bfe83, 32'hc158ca5b},
  {32'h43a129c6, 32'h43120e20, 32'hc29cb060},
  {32'hc3fcef3d, 32'h439dcefd, 32'h43767f48},
  {32'h4470abfc, 32'hc3c715ce, 32'h422fdb0a},
  {32'hc40ab808, 32'h431a4ee2, 32'hc28c4cb7},
  {32'h443ed1a4, 32'hc3aec3e6, 32'hc39ec912},
  {32'h440b6c13, 32'h434f50c9, 32'hc2d3d9fe},
  {32'h44138d7a, 32'h40a1d29c, 32'h427cb256},
  {32'hc4ae1a92, 32'hc4147fa7, 32'h43cbaef5},
  {32'h445e294a, 32'h429fb67e, 32'hc348c52c},
  {32'hc4dea5e6, 32'hc20c7369, 32'h438330a1},
  {32'h4340d278, 32'h4408737a, 32'h43771443},
  {32'hc4cc4812, 32'h41f82435, 32'hc335beec},
  {32'h44e41bcb, 32'hc3808965, 32'hc2cc7b96},
  {32'hc4b3607c, 32'hc1834275, 32'hc29e3bf5},
  {32'h44d2b445, 32'h43dbb6d8, 32'h4191d4aa},
  {32'hc4de0ebe, 32'hc11b3fea, 32'h4345f164},
  {32'h44f1a952, 32'hc3609bfa, 32'hc2f22ff0},
  {32'hc373447e, 32'hc0f77f75, 32'hc22819e4},
  {32'h43d41a45, 32'hc2bd0b20, 32'h43fd2802},
  {32'hc3b0e46a, 32'h43341d59, 32'h4350537d},
  {32'hc227b0a8, 32'hc4056322, 32'hc3450355},
  {32'hc48c828c, 32'h417907f3, 32'hc159e2de},
  {32'h44b7b3c7, 32'h437ae22d, 32'hc3898ee1},
  {32'hc4af01fc, 32'hc2e3f49e, 32'h43288898},
  {32'h447f5c71, 32'hc2a8e23a, 32'hc3309497},
  {32'hc4ea7523, 32'h3fb231b9, 32'h42934880},
  {32'h4433d691, 32'h43865cbd, 32'h43c62f6d},
  {32'hc3d7ebc7, 32'hc3e3c6e6, 32'hc405fdc9},
  {32'h43e59dbb, 32'h43b4e599, 32'h43048976},
  {32'hc4db472a, 32'hc30d9bca, 32'hc278f0fa},
  {32'h44961ea2, 32'hc404a13c, 32'h42012a86},
  {32'hc4ee574f, 32'h42887f37, 32'h43403da0},
  {32'h44e1dd40, 32'hc2c00687, 32'hc3bce6ff},
  {32'hc40a6b8f, 32'hc2ffc4d7, 32'hc2695844},
  {32'h4444a080, 32'hc2ecf588, 32'hc309470a},
  {32'hc50046dc, 32'h436d82f3, 32'h43174d3d},
  {32'h4316314c, 32'h4281e2d5, 32'hc217f1c0},
  {32'hc505f1d4, 32'h43414618, 32'hc1dd57c4},
  {32'h44051d19, 32'h428bcbe9, 32'h40d9aa1c},
  {32'hc5054c50, 32'hc305070b, 32'hc331b118},
  {32'h4476edfe, 32'h431953c2, 32'hc393db0d},
  {32'hc49eaacb, 32'h415e75bc, 32'hc2d9957c},
  {32'h43c7f008, 32'h42f1d289, 32'h43420947},
  {32'hc4d8f64a, 32'h438cde3b, 32'h430e6d80},
  {32'h43905a26, 32'hc085df84, 32'h439016d0},
  {32'hc4b13a85, 32'h439b37e8, 32'h42fb2878},
  {32'h44ee7e02, 32'hc27188bf, 32'h42d92a81},
  {32'hc513a277, 32'hc38a0d17, 32'h4384924f},
  {32'h43ef1362, 32'h404d1d82, 32'hc3397fcd},
  {32'hc4d95e88, 32'h436d2519, 32'hc344102e},
  {32'h44fd9c34, 32'h42aa2215, 32'h431d5113},
  {32'hc44a35ff, 32'hc34a2afa, 32'h42c67f68},
  {32'h44ad4479, 32'h426e043a, 32'h4349ff5e},
  {32'hc4b6bb80, 32'h430976eb, 32'hc283f1ba},
  {32'h4503276c, 32'hc3713711, 32'h40f7cef8},
  {32'hc4daab62, 32'h433e84e2, 32'h432e174f},
  {32'h44cffe57, 32'hbf7dbb80, 32'hc2b54a4b},
  {32'hc3d43b96, 32'hc1203575, 32'h428d2cac},
  {32'h44032320, 32'h42de3206, 32'h420b188b},
  {32'hc4f0908b, 32'hc3987efe, 32'h427fa1c1},
  {32'h448194fc, 32'hc2f0349b, 32'h4324c1e1},
  {32'hc4e66378, 32'hc2f7343c, 32'hc0b3f95d},
  {32'h44673cdc, 32'hc1ced436, 32'hc26056b4},
  {32'hc466ad2e, 32'hc21902fa, 32'h425d8e13},
  {32'h42b7b305, 32'hc33c7d2b, 32'hc374f549},
  {32'hc4ec6f7b, 32'hc2f56f84, 32'h437dd717},
  {32'h447e5790, 32'h4166fddd, 32'h439c4f10},
  {32'hc460d10c, 32'hc35675a4, 32'hc2a595f7},
  {32'h44043749, 32'hc30aabba, 32'hc30695e6},
  {32'hc48d910c, 32'h4386f62d, 32'h4222499e},
  {32'h43788d2c, 32'hc3099fab, 32'h418f2962},
  {32'hc4b0712e, 32'h427a188e, 32'hc2a1d4d4},
  {32'h44c9b049, 32'hc2821fc0, 32'h43188acf},
  {32'hc4c8e79e, 32'h43691a85, 32'hc120f832},
  {32'h44a74631, 32'hc2864bcd, 32'hc33dd1f9},
  {32'hc33a06a0, 32'h42a1652f, 32'hc1f95088},
  {32'h44065816, 32'h42bbfcea, 32'h427f76d3},
  {32'hc2a09bf8, 32'hc3a05c9f, 32'h43238560},
  {32'h451a406e, 32'h431b6086, 32'h4307f431},
  {32'hc4d0fbb9, 32'h421ce702, 32'hc38961fa},
  {32'h4523bcc4, 32'h4337beb2, 32'h41e2a77c},
  {32'hc4cc4976, 32'h4313d4c4, 32'hc3dc1ffa},
  {32'h446018c0, 32'hc2e6aad8, 32'h41d146eb},
  {32'hc46ca1bb, 32'h42f9c929, 32'hc31a4778},
  {32'h44cedfa4, 32'hc1ec4cd6, 32'h42d070b8},
  {32'hc4187472, 32'hc37b3d32, 32'hc32085b5},
  {32'h43c378e4, 32'hc2c9145e, 32'h3ff31db0},
  {32'hc3a76738, 32'hc35db39f, 32'hc31cf2a7},
  {32'h446adc3a, 32'h43716874, 32'hc2c076aa},
  {32'hc4b0652c, 32'hc2c17e64, 32'h4311f4b1},
  {32'h4337c5f4, 32'hc3dc0291, 32'h43784380},
  {32'hc4a652fc, 32'h42997f47, 32'h427aae89},
  {32'h43a25eb8, 32'h41eead60, 32'hc30dc839},
  {32'hc4b718fe, 32'hc38c8e41, 32'h4304f691},
  {32'h44b43198, 32'h41064f08, 32'h43b04eb7},
  {32'hc2c47ae8, 32'hc3d0ac5b, 32'h42d97ab1},
  {32'h44e0b8d2, 32'h4362babe, 32'hc2fdf8f2},
  {32'hc4d85fa0, 32'hc3861bf1, 32'hc35cce33},
  {32'h44c0361d, 32'hc2572231, 32'h423b1ee4},
  {32'hc492defa, 32'h43277a4b, 32'hc20336a8},
  {32'h443ecf88, 32'hc38fff90, 32'hc39eb7d2},
  {32'hc4fbaa97, 32'h432da337, 32'h436393ce},
  {32'h44a9a920, 32'h41ae66d8, 32'hc3384557},
  {32'hc4c51f9b, 32'h42b4767d, 32'h43904276},
  {32'h44df2553, 32'hc3ae0d40, 32'hc3915db4},
  {32'hc2cd4aa3, 32'h4355e371, 32'hc3b81dc7},
  {32'h426a2000, 32'hc33fa48a, 32'h43812b43},
  {32'hc4e2a26a, 32'hc3af3d5e, 32'hc16fc25b},
  {32'h445a9398, 32'h438d5702, 32'hc3a90d42},
  {32'h429360a4, 32'h4385d9a7, 32'hc2953cbd},
  {32'h442ee3bc, 32'hc3fc1862, 32'hc3020fa7},
  {32'hc504c4e0, 32'hc2af3e68, 32'h436c7ae0},
  {32'h44d25df0, 32'hc3037663, 32'h42f97487},
  {32'hc4f7c3d2, 32'hc1a0007f, 32'hc440978a},
  {32'h44fa0252, 32'hc2f0b4a1, 32'h429f19c7},
  {32'hc4eca7d4, 32'h42279003, 32'hc2f1f05d},
  {32'h44d269a3, 32'h436fc42b, 32'h43a38ca8},
  {32'hc12ac0c0, 32'h4343ca9a, 32'h43d986fa},
  {32'h445f8038, 32'hc300f004, 32'h4381581b},
  {32'hc3f8a7b8, 32'h429d5b02, 32'hc37c0b04},
  {32'h44b601ec, 32'hc384f0df, 32'hc367c8e1},
  {32'hc4b1989b, 32'h43a61edc, 32'hc399d64b},
  {32'h441fa410, 32'hc34fffcb, 32'hc4007c01},
  {32'hc5078edc, 32'h4289ca4d, 32'hc2c51f97},
  {32'h431d8594, 32'h42946260, 32'hc3133e75},
  {32'hc4a5bda4, 32'hc1f8c92e, 32'hc3578c20},
  {32'h44907ab4, 32'hc33e77aa, 32'h42d7221e},
  {32'hc3996f78, 32'h40e07c0e, 32'h41d9093f},
  {32'h445aa818, 32'hc132b9df, 32'h43e26517},
  {32'hc50b3bba, 32'h42ae2e28, 32'h42d7141f},
  {32'h44680488, 32'hc2dec908, 32'h43157da7},
  {32'hc3dd3138, 32'hc3ab7a3e, 32'hc3d1f045},
  {32'h44530156, 32'h4091c96a, 32'hc2e9e9de},
  {32'h42b39bc0, 32'h438a7943, 32'hc29f7391},
  {32'hc282b05f, 32'h42edcd4e, 32'h43a571b4},
  {32'hc50c0dc2, 32'hc30fc245, 32'hc365b086},
  {32'h4026b400, 32'h43961e49, 32'hc2a97a29},
  {32'hc4d816ae, 32'hc0ec5f7a, 32'hc3337d5b},
  {32'h44f867c1, 32'hc2d9c592, 32'h4364be1f},
  {32'hc4ec686e, 32'hc36120a0, 32'h418d0caa},
  {32'h44831cca, 32'hc30e0776, 32'h425af1c9},
  {32'hc439fef4, 32'h437041e4, 32'hc2e89b6f},
  {32'h44d4dc82, 32'h428ebb58, 32'h43839e89},
  {32'hc3e711e4, 32'h4399c0df, 32'h422c1e76},
  {32'h44c8116e, 32'h43994d7b, 32'hc31bbacb},
  {32'hc503e790, 32'h410a9144, 32'h431b6460},
  {32'h439085e5, 32'hc3a99d67, 32'h4324081e},
  {32'hc448fb84, 32'h42081cdd, 32'hc2a93fcd},
  {32'h442a6b76, 32'h43532af2, 32'h4333ff8c},
  {32'hc4e0e4cc, 32'hc32d7213, 32'h432ceec8},
  {32'h448328a0, 32'h433a65bb, 32'hc2e333c1},
  {32'hc40c159a, 32'h42fb68e0, 32'h436adef1},
  {32'h43e348bd, 32'h436ce447, 32'h436ab516},
  {32'hc5006046, 32'h429269bf, 32'hc1b49817},
  {32'h44bfaa2b, 32'hc34388cd, 32'hc45edbc5},
  {32'hc4f7a8ba, 32'hc303a739, 32'h420bfca9},
  {32'h447a4345, 32'h436607d8, 32'h4267f9db},
  {32'hc51ade66, 32'h40e00d77, 32'h42967302},
  {32'h44e10d34, 32'hc3281523, 32'h44096b38},
  {32'hc49f903b, 32'h428cacd8, 32'hc3722f88},
  {32'h45109d97, 32'hc2b80085, 32'hc2e7653e},
  {32'hc513251d, 32'hc311678e, 32'h43c29417},
  {32'h4524e1ca, 32'h4285d093, 32'hc38819ed},
  {32'hc46334f2, 32'hc348e1b0, 32'h41a665bb},
  {32'h443cdf64, 32'hc0eadcb7, 32'h43eb1153},
  {32'hc48bd8e0, 32'h43a41f9c, 32'hc31c3de0},
  {32'h44ea924d, 32'h43aea8e0, 32'hc343bc6f},
  {32'hc37a9530, 32'h43779d05, 32'hc325932d},
  {32'h4432baf0, 32'hc411a49e, 32'h433bfa4b},
  {32'hc3df3372, 32'h42e5142d, 32'hc3778af4},
  {32'h44e9b0d2, 32'hc2eb0f12, 32'h4351a024},
  {32'hc4ff9580, 32'hc3792fb5, 32'hc293a9f1},
  {32'h424d6f60, 32'hc3bb1819, 32'hc37b1fd0},
  {32'hc505cf17, 32'h43c02362, 32'hc38417ec},
  {32'h449b2fd4, 32'hc3ab8485, 32'h4309ea55},
  {32'hc47de2fc, 32'h43862ad7, 32'hc353c869},
  {32'hc307d7d0, 32'h4328a5d6, 32'hc30171dd},
  {32'hc4c58013, 32'hc2a2a4db, 32'hc3a09b14},
  {32'h44c299f6, 32'hc30cb1b7, 32'hc33b2fd0},
  {32'hc4f7cae4, 32'hc365c931, 32'hc326219d},
  {32'h4503175d, 32'hc3dcd2f6, 32'h43f06470},
  {32'hc4debde9, 32'hc3051cc7, 32'h4061a216},
  {32'h44af8e41, 32'hc2e72187, 32'h439ec915},
  {32'hc50350d2, 32'h41c36ef4, 32'h42d283d2},
  {32'h43203f70, 32'h43ff2053, 32'hc257619e},
  {32'hc5012eed, 32'hc3a71041, 32'hc3b0aea0},
  {32'h438e9708, 32'hc30b2269, 32'h4202e340},
  {32'hc4d47ddf, 32'h43c537d8, 32'h435bdb3f},
  {32'h450bacf1, 32'hc199aacf, 32'hc2339628},
  {32'hc3b4f40c, 32'hc254c910, 32'hc3179ab0},
  {32'h44c00b0e, 32'h439403f2, 32'h439e9dab},
  {32'hc509f43f, 32'h43208082, 32'hc308e75c},
  {32'h450f2f39, 32'hc28afe09, 32'hc3c0560b},
  {32'hc5143f36, 32'h43dd9073, 32'h429417c0},
  {32'h439bb85e, 32'h43692a28, 32'hc3ef15bf},
  {32'hc4ff209e, 32'hc3a02b16, 32'hc24827c2},
  {32'h451053f2, 32'hc3afb1f2, 32'hc285316d},
  {32'hc4b1c105, 32'h43485ddd, 32'hc3890744},
  {32'h44cb526c, 32'hc3c2a479, 32'h43861b1b},
  {32'hc2e58030, 32'hc40cfbf4, 32'h41a1a0f0},
  {32'h446add90, 32'hc39101b6, 32'hc2afc520},
  {32'hc48f7acd, 32'h420cb900, 32'h4322c96a},
  {32'h448ff165, 32'h42a69a99, 32'h429028b6},
  {32'hc517b8ec, 32'hc316c3be, 32'h430b77a2},
  {32'h4514eac3, 32'h4357dc93, 32'h409b3301},
  {32'hc40dba84, 32'h40cc3fc2, 32'hbf750b3a},
  {32'h43f2e838, 32'h432f7b7e, 32'h42cd9922},
  {32'h43446cc8, 32'hc1f865b0, 32'hc3d207e5},
  {32'h4492a302, 32'hc258d0eb, 32'hc2d7b5ad},
  {32'hc4f35ddc, 32'h4392f9fd, 32'h40930321},
  {32'h44d88200, 32'hc3a481bf, 32'h408ec868},
  {32'hc4033c8f, 32'hc2a89a3d, 32'hc28bbdfc},
  {32'h44dca2da, 32'h4317ccd0, 32'h43a30942},
  {32'hc4828e89, 32'h4268a298, 32'hc1b36c1f},
  {32'h442cbe39, 32'hc373fd49, 32'h4331147f},
  {32'hc4d4a698, 32'h4376c6ba, 32'h41a82630},
  {32'h438cfd82, 32'hc3aaf055, 32'h431bf36d},
  {32'hc2855d80, 32'hc2c4a8a9, 32'hc2660cd5},
  {32'h4478e9a6, 32'hc15085e6, 32'h429674c6},
  {32'hc43f8f65, 32'h4356ddcd, 32'hc3ab5caa},
  {32'h43ff4c34, 32'hc352e639, 32'hc3224d2a},
  {32'hc469a4b8, 32'hc30358fc, 32'h440c0a34},
  {32'h44b6255d, 32'h436005b4, 32'hc30dee8e},
  {32'hc4bc4a7a, 32'hc3d1da5d, 32'hc336ed00},
  {32'h451f5f0c, 32'hc30a7345, 32'h41ba7568},
  {32'hc50643c8, 32'hc369f99b, 32'hc13653f3},
  {32'h44f927af, 32'h43202c6b, 32'hc237bf26},
  {32'hc2bc78d1, 32'hc312d0cc, 32'h44031d53},
  {32'h4485e99e, 32'hc315d7ff, 32'hc38c68a0},
  {32'hc4b260f8, 32'h411b5072, 32'h4280a387},
  {32'h44ea94f5, 32'h431837e8, 32'hc28ef444},
  {32'hc47b9cc8, 32'hc2ba1f15, 32'hc30f366c},
  {32'h450e55de, 32'hc330d356, 32'h4166ba29},
  {32'hc4c826a4, 32'h42b8a6f4, 32'h42f3a08f},
  {32'h448654dc, 32'hc30ac9bc, 32'hc3042895},
  {32'hc48c2b54, 32'h43c7b020, 32'h42276d32},
  {32'h4434e972, 32'h4385edb1, 32'hc38481f9},
  {32'hc415f5ef, 32'h431d10ca, 32'h423b34b9},
  {32'h44665e07, 32'h4242a854, 32'h420378e0},
  {32'hc34b7700, 32'hc3774d93, 32'h42fdc254},
  {32'h4326b0b4, 32'h43219859, 32'hc224bbe7},
  {32'hc49a039b, 32'hc31fc2be, 32'h4192e55b},
  {32'h44ba1154, 32'h4334b49a, 32'hc304d005},
  {32'hc505382a, 32'h421b6d0f, 32'h43a25473},
  {32'h44b9647a, 32'h4253b15e, 32'hc3086d1c},
  {32'hc4128d44, 32'hc33c61fc, 32'hc1bef1af},
  {32'h4521528e, 32'hc35aa769, 32'hc26c3a03},
  {32'hc4a2fab6, 32'h42f3ce81, 32'h43e859e7},
  {32'h43ef4710, 32'h438738e7, 32'hc36a14e3},
  {32'hc4bb7a78, 32'h4284383d, 32'hc2db9186},
  {32'h43f38cdb, 32'hc2b6bd4c, 32'h42e09e04},
  {32'hc39ab888, 32'hc3208212, 32'h41859a4d},
  {32'h44f64303, 32'hc279ec36, 32'h43cb5779},
  {32'hc4e35972, 32'hc3cc3b8d, 32'hc2da1f71},
  {32'h44ee1e55, 32'hc30c0edc, 32'hc2ce11e9},
  {32'hc4f57984, 32'hc32bdeff, 32'hc36b5cee},
  {32'h4314c33c, 32'h439129bd, 32'hc27aad17},
  {32'hc50a1c1a, 32'h4353c63a, 32'h410b3009},
  {32'h45127ac3, 32'h42aa5beb, 32'hc37e1b0f},
  {32'hc42dde31, 32'h4348fc73, 32'h43c4b76c},
  {32'h44be22d8, 32'hc380e598, 32'h41867764},
  {32'hc4da7874, 32'h4232d6a5, 32'h42b36b00},
  {32'h44cdd793, 32'h437638ae, 32'hc3915af6},
  {32'hc4be4bcd, 32'h439a8e8e, 32'hc303e3c9},
  {32'h44d5e8d0, 32'hc2cec9f8, 32'h437eaec2},
  {32'hc4f4c45c, 32'h432e0214, 32'hc2183a23},
  {32'h43be8e44, 32'hc342399e, 32'hc3e01714},
  {32'hc48bee78, 32'h42f5ad20, 32'h433c460d},
  {32'h435bd6f0, 32'h42f2b414, 32'h426b6834},
  {32'hc51dd19d, 32'h434dd434, 32'hc3c1e286},
  {32'h44d2e39a, 32'hc28e9973, 32'hc3b3a71a},
  {32'hc4d9974e, 32'h43006d67, 32'hc302ec56},
  {32'h451bb706, 32'h42c35d7a, 32'hc30c66fa},
  {32'hc4b98165, 32'hc30896e6, 32'hc3022720},
  {32'h44fd395a, 32'h42097948, 32'hc1bd26cf},
  {32'hc48b2e9e, 32'h42f273c5, 32'h422df637},
  {32'h44b0cf0b, 32'hc35ed369, 32'h40b969ab},
  {32'hc48c7dec, 32'hc29c2176, 32'hc2cbaf9f},
  {32'h447c28c2, 32'hc35162e1, 32'hc28cbc64},
  {32'hc4f500bc, 32'hc38b7dad, 32'h438de6c9},
  {32'h44cfc793, 32'hc31a0810, 32'h42a3fd0f},
  {32'hc3bd399c, 32'h437dabbb, 32'h43a85767},
  {32'h44f84b82, 32'h42a589b8, 32'hc2b6c739},
  {32'hc3b9d290, 32'h41fb9c51, 32'h43961850},
  {32'h44845942, 32'hc3a6e8bd, 32'hc30fae41},
  {32'hc452eb2c, 32'h42ac2138, 32'hc383ad87},
  {32'h450ac29f, 32'hc0184d4a, 32'hc2b2adcd},
  {32'hc41d6868, 32'hc30227ef, 32'h43cf5c84},
  {32'h440022ae, 32'hc34df048, 32'hc29d4c5f},
  {32'hc4eb58e8, 32'hc182ea9f, 32'hbfc2e97c},
  {32'h452ff588, 32'h419e9f37, 32'h4384ddf1},
  {32'h44569542, 32'hc3602427, 32'hc2c01245},
  {32'hc4c3eee3, 32'hc2a1a657, 32'hc2ded231},
  {32'h445cc78c, 32'h4324b777, 32'hc2166f41},
  {32'hc43d0020, 32'hc34ebccc, 32'h438db053},
  {32'h4482284b, 32'h437b05d0, 32'hc2ecdda0},
  {32'hc49d6803, 32'h43614903, 32'hc3021e1c},
  {32'h43fd6027, 32'h4312d5c0, 32'hbfdd0018},
  {32'hc4cb3465, 32'h431d8574, 32'h41abef25},
  {32'h446d34bd, 32'h438ee298, 32'hc37f99e7},
  {32'hc2a44600, 32'h43ea804a, 32'hc330bf0f},
  {32'h4488a587, 32'hc204df5e, 32'hc31d85a6},
  {32'hc413340b, 32'h43ac49d0, 32'h4296f1ef},
  {32'h43977704, 32'h417037de, 32'hc376fe37},
  {32'hc22bb630, 32'h43984f9f, 32'hc1e74b05},
  {32'h44c1aac8, 32'hc22ae0ad, 32'h4301353b},
  {32'hc4dcf5c4, 32'hc22e3a6b, 32'h43b85e83},
  {32'h4504fd0b, 32'hc31305a2, 32'hc28334fa},
  {32'hc427239d, 32'hc33effed, 32'h4309342b},
  {32'h4519e17e, 32'hc29d02e0, 32'hc3154f45},
  {32'hc4c06c8c, 32'h43158cef, 32'h435fb484},
  {32'h430943df, 32'hc38b695a, 32'hc3359bfa},
  {32'hc4f3b1da, 32'h434e5738, 32'hc33fb494},
  {32'h44bde5de, 32'hc2b7ad31, 32'hc38f594d},
  {32'hc4855107, 32'hc31b5cbe, 32'h40d4dd5c},
  {32'hc1ec4640, 32'h43cd44cc, 32'hc317ee79},
  {32'hc4fbe797, 32'h43f55295, 32'h436dba5b},
  {32'h44b12412, 32'hc405e862, 32'hc2dd0893},
  {32'hc4e605c8, 32'hc37932ca, 32'h4112cc98},
  {32'h44f3d450, 32'h432db95c, 32'hc30c8df5},
  {32'hc383ae8c, 32'h433f3dae, 32'hc22bf85b},
  {32'h43a24112, 32'h44082c6f, 32'h4314f608},
  {32'hc3f63c7d, 32'hc30669d9, 32'h42947479},
  {32'h426182e0, 32'hc2855a6f, 32'h42cfce2c},
  {32'hc460539b, 32'hc2c2923b, 32'h42a1464a},
  {32'h44852675, 32'hc2467cce, 32'hc219f2cb},
  {32'hc4ac94d9, 32'hc24ce924, 32'h439c8532},
  {32'h450cf196, 32'h4331c780, 32'h43a25fca},
  {32'hc42d2110, 32'h43287f7c, 32'hc2546552},
  {32'h450b4fed, 32'h4391c79a, 32'hc369ab6c},
  {32'hc3403380, 32'h43b581cb, 32'hc3ca9407},
  {32'h444b38dc, 32'h428ae55f, 32'h41b8f976},
  {32'hc3e12e70, 32'h419ff7f6, 32'h43387206},
  {32'h443776de, 32'hc3585017, 32'hc28bf0ac},
  {32'hc4f131f9, 32'h43358972, 32'h43bb2e38},
  {32'h435a1d9e, 32'h40b8bf5c, 32'hc3925a34},
  {32'hc4ff3350, 32'hc28068c7, 32'hc33023ec},
  {32'h439ad468, 32'h43b40217, 32'h42aee3cb},
  {32'hc448218c, 32'hc28814e6, 32'hc2a4e56b},
  {32'h44559032, 32'h4348597a, 32'h42d9270f},
  {32'hc4995482, 32'hc0f056c7, 32'h436ad167},
  {32'h444d2e07, 32'h42cc2bba, 32'h428232ff},
  {32'hc507ba89, 32'h42ff8cc8, 32'h43223163},
  {32'h44d09635, 32'h429aeffb, 32'hc2d523f2},
  {32'hc4803dce, 32'h4381b765, 32'hc28684c2},
  {32'h448abf61, 32'h43319d2f, 32'h435e9422},
  {32'hc4b2b617, 32'h4381d132, 32'hc3a25ac2},
  {32'h44a46bbf, 32'h43806091, 32'h41e59f8d},
  {32'hc44caa26, 32'hc12d56aa, 32'hc2f47140},
  {32'h44ef3b45, 32'h435a8c00, 32'hc35fe715},
  {32'hc4bc3b4a, 32'h426e7532, 32'h41ebf8cf},
  {32'h449e5fe5, 32'hc3788109, 32'h42e346d6},
  {32'hc4751600, 32'hc392b518, 32'h42b2661a},
  {32'h43442313, 32'hc300a491, 32'hc2cdba42},
  {32'hc44f09e1, 32'h431649eb, 32'hc2ca3976},
  {32'h440da16c, 32'h43978d43, 32'h4386f6fe},
  {32'hc48580c1, 32'hc38429ae, 32'hc17ad81d},
  {32'h439d59ae, 32'h43f681eb, 32'h43da67a5},
  {32'hc41a5696, 32'hc117dca0, 32'hc21fe8f9},
  {32'h44d188d7, 32'hc40aa560, 32'h4295089a},
  {32'hc490b020, 32'h4321155e, 32'h438f0fd2},
  {32'h449152df, 32'hbf6636d0, 32'hc3817509},
  {32'hc5084104, 32'hc31cfd89, 32'h4339e51e},
  {32'h44d4c637, 32'h424c0526, 32'hc3a18032},
  {32'hc42927e0, 32'h4385b6bb, 32'h43b201db},
  {32'h451411c3, 32'h437e13fa, 32'h432ad420},
  {32'hc452a901, 32'h4373b809, 32'hc2a2b90e},
  {32'h4507f1e0, 32'h42e989c0, 32'hc365eb54},
  {32'hc2ca14c0, 32'h437d6319, 32'hc339f587},
  {32'h4253e0e0, 32'hc2bd733e, 32'hc3231fee},
  {32'hc432c290, 32'hc2aebf94, 32'hc386cf2b},
  {32'h4482a3b2, 32'hc3151e19, 32'h43614a4b},
  {32'hc49c7aaa, 32'h42f6e0dd, 32'hc319bec9},
  {32'h44234b00, 32'h435856c0, 32'h435eadbb},
  {32'hc4f7f4db, 32'h436c1cc1, 32'hc3710f74},
  {32'h43b1aba8, 32'hc216a0b3, 32'h43480bf4},
  {32'hc4a038ea, 32'hc2e738e4, 32'h42f1d5ef},
  {32'h44c456bf, 32'hc23ba057, 32'hc39f6bc4},
  {32'hc41a262d, 32'h42941c6b, 32'hc4087e5f},
  {32'h44c0edc2, 32'hc3babdbe, 32'hc29e045e},
  {32'hc508e770, 32'h41ef4eba, 32'h42e53455},
  {32'h44e6319f, 32'h41bdc8ac, 32'hc2d3aee2},
  {32'hc4640d78, 32'hc388e896, 32'hc33fcc3b},
  {32'h4449de84, 32'h4295ff94, 32'hc383bdcd},
  {32'hc4d0942c, 32'hc31e0b47, 32'h41841e62},
  {32'h44adcc65, 32'hc32098a9, 32'hc2787aa8},
  {32'hc44fbc56, 32'h42a204f8, 32'h43d8f749},
  {32'h44877120, 32'hc3acd441, 32'h4394ef19},
  {32'hc49cde58, 32'hc39d2f65, 32'hc10fc4fd},
  {32'h45135689, 32'h43184155, 32'h42e77fb3},
  {32'hc4ac2f41, 32'hc33032f7, 32'hc2935265},
  {32'h449a0591, 32'h420967f0, 32'h42b2c7f0},
  {32'hc5083e5b, 32'hc3616003, 32'hc324bea5},
  {32'h44ff9024, 32'hc38b984c, 32'h43eeb5df},
  {32'hc4ca274f, 32'h425ab608, 32'h42dae875},
  {32'h44be0c2c, 32'hc107d344, 32'hc158a606},
  {32'hc45589a5, 32'h42380b91, 32'h439ef15d},
  {32'h4478f8b8, 32'hc168cfa2, 32'hc19945df},
  {32'hc3bd7468, 32'hc2b6b451, 32'hc18cf741},
  {32'h43bee194, 32'h439b981a, 32'hc2022adf},
  {32'hc3be1b79, 32'h4403bb4e, 32'hc2035413},
  {32'h45177643, 32'hc3321feb, 32'h43958874},
  {32'hc4f33ace, 32'h421972ec, 32'h439ed5b4},
  {32'h447abd42, 32'h43badca8, 32'hc1ac6579},
  {32'hc4cf5bbe, 32'h43823e83, 32'h438c1cbf},
  {32'h449cde6a, 32'h42849498, 32'h43842d9d},
  {32'hc44129ef, 32'h424d255c, 32'hc30e17aa},
  {32'h439ad998, 32'hc2931dd6, 32'hc26cc320},
  {32'hc4d2128f, 32'h424dbef7, 32'hc14a80ad},
  {32'h447be1a6, 32'hc2834ae4, 32'hc34149a6},
  {32'hc5009e2c, 32'h42c0d399, 32'h43327ac5},
  {32'h44f22929, 32'hc348ef99, 32'hc0f7c097},
  {32'hc4a413ca, 32'hbfe15364, 32'h4347e63e},
  {32'h44e2c49f, 32'hc31d1a70, 32'h4365a9a8},
  {32'hc42d1dec, 32'h42a516cd, 32'hc2bebd6c},
  {32'h4478267a, 32'h41c3176d, 32'h42bac970},
  {32'hc480b7d3, 32'hc3bd6fb3, 32'hc221775d},
  {32'h450db0bf, 32'hc28ea49e, 32'hc2465f02},
  {32'hc371d538, 32'h4383abdc, 32'hc2fa9f7e},
  {32'h448050ad, 32'h42c71676, 32'h4364578f},
  {32'hc45bd73d, 32'hc38048e6, 32'hc39b00ca},
  {32'h44a9a368, 32'hc272af75, 32'h4303bec6},
  {32'hc4d6f6e5, 32'h43b59fbf, 32'hc4135234},
  {32'h441d0b9c, 32'hc217b7bb, 32'h416d2911},
  {32'hc471d0cd, 32'hc3dc4bc6, 32'hc32bb80a},
  {32'h44c9631b, 32'h4315c01a, 32'hc3673ead},
  {32'hc42d8ea6, 32'hc328050c, 32'hc3e24a2c},
  {32'h43d6d610, 32'h4329074f, 32'h4291855f},
  {32'hc49e1f2c, 32'h421997ba, 32'h40807953},
  {32'h448c8c55, 32'h42e909ac, 32'hc3891b42},
  {32'hc4a73297, 32'hc31dcc18, 32'h4384996a},
  {32'h44558710, 32'h43320a06, 32'h419ebc2c},
  {32'hc4e0b09a, 32'h41524ca5, 32'hc3078a4c},
  {32'h44fa1d76, 32'hc219a78b, 32'h4301c6c9},
  {32'hc2e721e0, 32'hc35e61e9, 32'h41ac248c},
  {32'h43d10d84, 32'h43a0d708, 32'h432e64c1},
  {32'hc47c23f2, 32'hc0e3ce3d, 32'hc3319dec},
  {32'h4363bbd8, 32'h42494517, 32'h41910826},
  {32'hc405ae09, 32'hc2c7a73c, 32'h433e3225},
  {32'h45155810, 32'hc3592f4b, 32'h413fd7be},
  {32'hc4bcfba0, 32'h43c2ee76, 32'h43ddfef7},
  {32'h44339370, 32'hc3586fde, 32'h432a1abf},
  {32'hc4b3de5a, 32'hc31ea9ac, 32'h439e8dfb},
  {32'h4509060f, 32'hc2e70eca, 32'h42ef3f6e},
  {32'hc4584c99, 32'hc29b5a69, 32'h42239b72},
  {32'h44d208de, 32'hc2426e1e, 32'h421286fe},
  {32'hc50991d4, 32'hc191451a, 32'h434ac3e0},
  {32'h44e8a5b4, 32'hc35aac64, 32'h43041393},
  {32'h42e641d9, 32'hc30c2865, 32'hc09b5347},
  {32'h441244c0, 32'h430cb224, 32'hc39ebe0b},
  {32'hc494561e, 32'hc2ab9983, 32'hc3a44df0},
  {32'h44b7f220, 32'hc24d4220, 32'h437f36b6},
  {32'h43b34208, 32'hc407dc07, 32'hc3d46054},
  {32'h4498c67f, 32'h43b88b7e, 32'hc305947f},
  {32'hc4092ef9, 32'h4335d22d, 32'hc3b79f66},
  {32'h451080bb, 32'h4355eda5, 32'h4395268e},
  {32'hc3a3886c, 32'h4369d46f, 32'hc38b37a6},
  {32'h44fa9b81, 32'hc1a8097e, 32'h4323430b},
  {32'hc4ddc2fb, 32'h42e1f0bf, 32'h438cd298},
  {32'h44c9c59e, 32'hc3e7a26a, 32'hbe9c47dd},
  {32'hc4a6d55e, 32'h43a083ba, 32'h43a6eec0},
  {32'h44c0d663, 32'hc2b5f5aa, 32'hc2a77313},
  {32'h42819e3e, 32'hc3dc77b9, 32'h4383a270},
  {32'h450b36b6, 32'hc0d4bb4a, 32'hc3939645},
  {32'hc49cc45e, 32'hc38c1851, 32'h42e7c1e5},
  {32'h449cd861, 32'hc3e38484, 32'hc27d8683},
  {32'hc3eef4b1, 32'h4286cbdf, 32'hc3189670},
  {32'h4506a9ac, 32'h42659b38, 32'h4298d8da},
  {32'hc43434c2, 32'hc40b5878, 32'h43ec0041},
  {32'h428ebd68, 32'hc349c84e, 32'h43ace8d8},
  {32'hc4c22711, 32'hc307a537, 32'hc30188d5},
  {32'h43ff2d54, 32'h407c7e48, 32'hc0c43311},
  {32'hc5009eb8, 32'hc303748d, 32'hc325bd05},
  {32'h4507e179, 32'h4222475e, 32'h42daf9a5},
  {32'hc4d2b388, 32'hc3aaae4d, 32'hc2b77ae6},
  {32'h448c1068, 32'hc20e57b3, 32'h428ded1c},
  {32'hc4e73000, 32'hc1654a10, 32'h432a763d},
  {32'h44178938, 32'h424644d2, 32'hc2ed8773},
  {32'h4264d580, 32'h43b7952c, 32'h43442849},
  {32'h44cfc384, 32'h42e7a2d7, 32'hc301979a},
  {32'hc4b239ce, 32'h42f02574, 32'h42bf57de},
  {32'h449cf0bc, 32'hc2e08cda, 32'h4408a5a6},
  {32'hc513547b, 32'h43513ad9, 32'hc2af66ee},
  {32'h43f776c7, 32'hc1c1a628, 32'h4304c34f},
  {32'hc472e808, 32'h428fbc26, 32'hc03c7ec5},
  {32'h43aea803, 32'h439af907, 32'hc1a3a1bd},
  {32'hc50b80dc, 32'hc114df5a, 32'h43a7b006},
  {32'h44da68fb, 32'hc2a17b6a, 32'hc24b3fa7},
  {32'hc41ac694, 32'hc31caadb, 32'h4197b5f6},
  {32'h44f3251e, 32'h435e9735, 32'hc293fbe5},
  {32'hc4830c15, 32'hc3a8fa0b, 32'hc2c4748c},
  {32'h448e8b1d, 32'h4400df7f, 32'h43feeae6},
  {32'hc50541a8, 32'h43133153, 32'hc312ed1d},
  {32'h449f1792, 32'h43259c0c, 32'hc3e922ad},
  {32'hc4038e55, 32'hc3454565, 32'hc1c9ba88},
  {32'h43bb5297, 32'hc30d0ac4, 32'hc34d0537},
  {32'hc4780f4a, 32'hc322d59e, 32'hc359afa7},
  {32'hc3b62e8e, 32'h4324c3bd, 32'h44075062},
  {32'hc48841dc, 32'hc361c5f9, 32'hc38aecd0},
  {32'h44861b88, 32'h42987fdb, 32'h43e3edcd},
  {32'hc483e5ae, 32'hc20ee66d, 32'h43ad6c88},
  {32'h4496d86d, 32'h4390ec94, 32'h43627745},
  {32'hc4b29798, 32'h41cce22f, 32'h430ae764},
  {32'h44c68c74, 32'hc21b3930, 32'h42908752},
  {32'hc4c8bb32, 32'h42b9c9c3, 32'h43992e84},
  {32'h44d84ef8, 32'h42af2e8f, 32'hc214afe3},
  {32'hc3bb2ebb, 32'hc3192eaa, 32'h433389cd},
  {32'hc2fff620, 32'hc1c48eeb, 32'h4307f23b},
  {32'hc41314a2, 32'h4316c40a, 32'h44014f2f},
  {32'h441bfdf0, 32'hc3928e9a, 32'hc1d25774},
  {32'hc49f9086, 32'h42939c33, 32'h430c1e98},
  {32'h4504c988, 32'h425e1219, 32'hc185051d},
  {32'hc468b5ad, 32'hc25b008b, 32'h41d1cde0},
  {32'h44c6be82, 32'hc2bd4f1d, 32'hc3114961},
  {32'hc4834220, 32'hc26ccda8, 32'h42ce5581},
  {32'h44dd51cb, 32'hc2dcd420, 32'hc325cddf},
  {32'hc49fdad3, 32'h435c29d0, 32'h41f3d163},
  {32'h449c4ac1, 32'hc3db0766, 32'h42cbb553},
  {32'hc3f285c9, 32'h43d06355, 32'h43692249},
  {32'h44f79f1f, 32'h42ca1b8c, 32'hc419d2d8},
  {32'hc509babd, 32'h42a6634e, 32'hc34d1013},
  {32'h44536f5a, 32'hc3715f2f, 32'h418e64ae},
  {32'hc4e297ec, 32'h43000aea, 32'hc32f542e},
  {32'h450215d7, 32'h4383ef87, 32'h42bdeec0},
  {32'hc50bc398, 32'hc159b2d5, 32'h42b5425e},
  {32'h446a19e8, 32'hc2f79852, 32'hc299a8c6},
  {32'hc4bea0a9, 32'hc2c66ef5, 32'hc3bd4d90},
  {32'h44db52c1, 32'hbe17ef78, 32'hc35a9474},
  {32'hc4654940, 32'hc2943a36, 32'h441209bd},
  {32'h42376ac8, 32'hc1f3970a, 32'h440ab51a},
  {32'hc34a23fe, 32'hc34532ee, 32'h40c480ea},
  {32'h44e9df66, 32'hc25610c6, 32'h43144a01},
  {32'hc43d8b41, 32'h430e80e7, 32'hc2bdec3b},
  {32'h44fc1cf6, 32'hc34e141c, 32'hc30789a8},
  {32'hc3bac098, 32'h4365f47f, 32'h43839fa8},
  {32'h44d0aff0, 32'hc37ab4fe, 32'hc38d2c45},
  {32'hc4808e6a, 32'h42f8e96c, 32'h4278db04},
  {32'h44a9b28e, 32'hc0e823de, 32'h42e06c38},
  {32'hc33ecd24, 32'hc29e5545, 32'h438fc1ad},
  {32'h44434ec2, 32'h437025e4, 32'h433817ea},
  {32'hc4d27cc6, 32'h436b9746, 32'hc3246db2},
  {32'h449542c8, 32'hc2225dc4, 32'hc35c9932},
  {32'hc464abe3, 32'h43140176, 32'hc3a24647},
  {32'h44e3ce24, 32'hc144fcc6, 32'hc36ded34},
  {32'hc449e20e, 32'h436f563f, 32'hc2b7cd70},
  {32'h451e601e, 32'hc261fce3, 32'hc2855be7},
  {32'hc4c93c41, 32'h42043327, 32'hc3a32c08},
  {32'h44592a4c, 32'h433eb171, 32'hc3cc830b},
  {32'hc2ad003c, 32'h42a9ff94, 32'hc30e7f64},
  {32'h445575b1, 32'hc2abc5f5, 32'hc2ab231c},
  {32'hc41216b6, 32'h42fd6b45, 32'h43a4254f},
  {32'h4502db6f, 32'hc1302832, 32'hc31a43aa},
  {32'hc4875e05, 32'hc3918adc, 32'h4293021c},
  {32'h44d08f1a, 32'hc2b01b8f, 32'hc360ee35},
  {32'hc4f8a23a, 32'hc399850a, 32'hc3c88c8f},
  {32'h44b3e452, 32'h4185608f, 32'hc1963c8a},
  {32'hc505eba0, 32'h41213bdb, 32'h435f54ea},
  {32'h44b8856d, 32'h434c3609, 32'h42530c34},
  {32'hc4fc4c8d, 32'h42249b8b, 32'hc2c7f706},
  {32'h41007bc0, 32'h432fc430, 32'hc1beca06},
  {32'hc3fc48c4, 32'h43527daa, 32'h43923347},
  {32'h4500e0c6, 32'hc3bd67ed, 32'hc2683f13},
  {32'hc3a44bda, 32'hc38b21c1, 32'hc35faeeb},
  {32'h44b357e1, 32'h4366ba74, 32'hc320e13a},
  {32'hc4dcfb64, 32'h430e961d, 32'hc18db029},
  {32'h44b9f4b2, 32'h42b76230, 32'hc332cdfd},
  {32'hc3301d80, 32'hc32ced0b, 32'h430ace7b},
  {32'h44c91825, 32'hc3099952, 32'hc356a498},
  {32'hc502eb9f, 32'h42451b4c, 32'hc2ea89d1},
  {32'h44959736, 32'hc2b6c361, 32'h438d7b4f},
  {32'hc504a9de, 32'hc39131c5, 32'hc05c0992},
  {32'h44bb7d5f, 32'hc2902cf8, 32'hc335034a},
  {32'hc400e23e, 32'h42f130ed, 32'hc3b23058},
  {32'h44a0b2ed, 32'h42bc2c3f, 32'hc161d423},
  {32'hc4ba0f4a, 32'hc3ef2a62, 32'h4329b79c},
  {32'h43a8b788, 32'h43105a1b, 32'h4238111b},
  {32'hc4312c7e, 32'hc1ec35b1, 32'hc31223b9},
  {32'h45101d08, 32'hc3d83766, 32'hc2e6acf0},
  {32'hc513ca2c, 32'hc312a785, 32'h430c212d},
  {32'h44a385bf, 32'h437b2410, 32'h436f936e},
  {32'h429887d0, 32'h4208222f, 32'hc2923fef},
  {32'h4425d335, 32'hbfd9a751, 32'h4257b421},
  {32'hc34f97ec, 32'hc33b9b33, 32'hc3739758},
  {32'h43eb6230, 32'hc2bb8184, 32'h439b1c53},
  {32'hc501c8e0, 32'h43a7f5f6, 32'hc31f09bf},
  {32'h450241c6, 32'hc31151ef, 32'hc3788250},
  {32'hc4104de8, 32'h3f09daf0, 32'h432fbec6},
  {32'h44866c80, 32'hc0b5edab, 32'h43a99cdd},
  {32'hc39895b8, 32'h41b58122, 32'h433c6deb},
  {32'h43dc0a46, 32'hc2ab3f1d, 32'h4218c9e2},
  {32'h43459280, 32'h431871c7, 32'hc2934a60},
  {32'h4501e0f9, 32'hc30d4739, 32'hc3cb4ae1},
  {32'hc425209a, 32'hc380cd41, 32'hc29fef69},
  {32'h44878f37, 32'h43630b21, 32'hc2d6a956},
  {32'hc38ac348, 32'hc29e7b18, 32'hc437ca7f},
  {32'h4452330c, 32'hc3bfea11, 32'h4312180b},
  {32'hc4e9371a, 32'h43208896, 32'h43908479},
  {32'h44b4d905, 32'hc3e1031a, 32'hc206dbdc},
  {32'hc4c06c84, 32'hc29ad9c4, 32'h42e1bdce},
  {32'h446a0fb4, 32'hc383c024, 32'h43fd2a42},
  {32'hc49efdfc, 32'h42f4e652, 32'hc3084292},
  {32'h4455c789, 32'hc09cc563, 32'hc3462b6a},
  {32'hc4929d28, 32'hc26ecc71, 32'h418e8d4b},
  {32'h44c9d0ca, 32'h43b1e8f5, 32'h43455a2a},
  {32'hc4e7dc41, 32'hc03d4eb8, 32'h4328c8c5},
  {32'h450b6c87, 32'h4390c0af, 32'hc3d92a3f},
  {32'hc3576320, 32'hc36bfdf9, 32'hc3af55d5},
  {32'h44a54a8f, 32'hc2b31206, 32'hc3386d8f},
  {32'hc4961338, 32'h43790b18, 32'h43abffb1},
  {32'h4503c742, 32'hc37e8b14, 32'h420ea369},
  {32'h43593800, 32'h4315b927, 32'hc309b016},
  {32'h443ff31e, 32'hc2ae1851, 32'hc222160f},
  {32'hc34b6fae, 32'hc2e33d5c, 32'h4404f2a7},
  {32'h45070ddd, 32'hc3813a71, 32'hc2cbeb2d},
  {32'hc504def1, 32'h42fac3da, 32'hc30904fa},
  {32'h43fb0734, 32'hc35ebd97, 32'hc30471fd},
  {32'hc4e56fab, 32'h433a9a33, 32'hc3304a70},
  {32'h44a0bbcc, 32'h423eecc2, 32'hc162c16d},
  {32'hc48c89a8, 32'hc378385a, 32'h42a0890f},
  {32'h44642fb6, 32'h405349f0, 32'hc305c217},
  {32'hc4f4075c, 32'h429c14d1, 32'h42faa722},
  {32'h43d3bbf4, 32'hc306743b, 32'h43986f53},
  {32'hc4b21133, 32'hc2382bb4, 32'h42c49841},
  {32'h44a88af0, 32'h40889ea8, 32'h430cabfe},
  {32'hc45ed464, 32'h43e6c660, 32'hc3a4199d},
  {32'h442e12ee, 32'hc266588b, 32'h43995e5e},
  {32'hc4f157bf, 32'hc36556ad, 32'hc31cddfc},
  {32'h447b58b0, 32'hc341f8eb, 32'h439c0a74},
  {32'hc4a6e3c7, 32'h43ead34e, 32'h4192522e},
  {32'h441db046, 32'h43960630, 32'h4396ea79},
  {32'hc4f2d3b4, 32'hc2352d7a, 32'hc2979841},
  {32'h45214abd, 32'hc3ac8e82, 32'h444754da},
  {32'hc50c883d, 32'h438a2f78, 32'hc3d6e1a8},
  {32'h44dd4458, 32'h42ac2e84, 32'h4201a76f},
  {32'hc4aff0de, 32'hc2a80ffd, 32'hc2c83eb4},
  {32'h42255720, 32'hc30050d9, 32'h42ef81a9},
  {32'hc4d36b86, 32'h428ac3c6, 32'hc15037bb},
  {32'h444f064a, 32'h41c53bea, 32'hc3361b97},
  {32'hc3b59404, 32'hc1856475, 32'h41fa1c1f},
  {32'h4407e0dc, 32'hc303dc2b, 32'hc3804426},
  {32'hc51e1628, 32'h43810507, 32'h4330afef},
  {32'h43e8f694, 32'h4321381d, 32'h42ca9322},
  {32'hc297c8e0, 32'h42d5eae6, 32'hc1f69cea},
  {32'h4521cf6f, 32'hc31241c1, 32'h42eb363c},
  {32'hc4a968ef, 32'h43a04a0c, 32'h41550ebb},
  {32'h44a80096, 32'hc312d3b8, 32'h427189bb},
  {32'hc4911c20, 32'hc3291bb1, 32'hc136159a},
  {32'h4485d27e, 32'h438ee38f, 32'h4217d674},
  {32'hc4bcab0c, 32'h43900ffe, 32'hc376af2a},
  {32'h449ad299, 32'h4390276d, 32'hc146530d},
  {32'hc33d2cc0, 32'hc359ed54, 32'h439f2889},
  {32'h44b3eb63, 32'hbffa2514, 32'h42763140},
  {32'hc3c74dee, 32'hc35b005b, 32'h4408a52c},
  {32'h442e695c, 32'hc224f792, 32'hc2580f73},
  {32'hc486518b, 32'hc1b22c86, 32'hc2946565},
  {32'h44aa783a, 32'hc37a9bc8, 32'h43b5ce64},
  {32'hc4df45e9, 32'hc1c6cb86, 32'h419b09da},
  {32'h450151c8, 32'h42e9523b, 32'hc32443b3},
  {32'hc515fdde, 32'hc2460171, 32'hc3444bbe},
  {32'h44b4cafc, 32'hc3a01868, 32'hc30d9ec5},
  {32'hc416f08e, 32'hc3fa21fa, 32'h433d63cf},
  {32'h44f99b0a, 32'hc1888d85, 32'h43a6ec17},
  {32'hc4ba76d8, 32'hc35dce57, 32'h4309c35b},
  {32'h44534d7e, 32'h4306e2c9, 32'hc3019cca},
  {32'hc4ea0ae2, 32'hc12f14ea, 32'hc3e34c07},
  {32'h44bebdca, 32'hc39b0ca9, 32'h4305fcb0},
  {32'hc464d8f6, 32'h43b03177, 32'hc30cbfad},
  {32'h44f18833, 32'hc19ca2cb, 32'hc3ac362b},
  {32'hc4f709db, 32'h4253cff0, 32'hc35a2d80},
  {32'h44b7b607, 32'h43887abc, 32'h43aa35b4},
  {32'hc4ed76a1, 32'hc391ab30, 32'hc368dd81},
  {32'h44b2506b, 32'h43148618, 32'hc25b2aa2},
  {32'hc4d7d010, 32'hc0682af0, 32'hc382921e},
  {32'h44b52a21, 32'hc25c9b4b, 32'hc2b3d862},
  {32'hc43f5c1c, 32'h428a4d7c, 32'hc2c6b57e},
  {32'h44cff682, 32'h4382d70c, 32'h4220ed5d},
  {32'hc5004c99, 32'h435d4bde, 32'hc336edf6},
  {32'h44d7464f, 32'h425864f9, 32'hc365c3fc},
  {32'hc4c17134, 32'hc29f8eb1, 32'hc1e612b4},
  {32'h439ac71c, 32'hc39eb46b, 32'h43183191},
  {32'hc43a96b8, 32'h428ae35f, 32'hc1e95929},
  {32'h4365e21e, 32'h433ddb96, 32'hc260b017},
  {32'hc3a01120, 32'hc42d0d47, 32'h4324a59d},
  {32'h45149545, 32'h430fd9e6, 32'hc1c9a321},
  {32'hc30d68be, 32'h41d6aa77, 32'hc3664337},
  {32'h42f0f600, 32'hc2bcd626, 32'h42c6c92b},
  {32'h427fe5c0, 32'hc389e6fc, 32'hc37d1757},
  {32'h43678530, 32'hc3c9b5a4, 32'hc0181c88},
  {32'hc4b2c6ed, 32'h418d2ac9, 32'h418b89a2},
  {32'h446c9996, 32'hc28f67ad, 32'h4249b500},
  {32'hc466d429, 32'hc33cf940, 32'hc33884dc},
  {32'h451413dd, 32'hc355a055, 32'h437d84c2},
  {32'h3fc50800, 32'h42f1acad, 32'hc400996e},
  {32'h422cace6, 32'h42cb10fb, 32'h43dbb337},
  {32'hc4c6c6e8, 32'h4265d07a, 32'hc2b55382},
  {32'h44fd998b, 32'h418272ac, 32'hc208cd83},
  {32'hc488313c, 32'hc2f9f1eb, 32'h438aa6a5},
  {32'h42cf45e8, 32'h42a7fea8, 32'h43b1dc9b},
  {32'h41aab0dc, 32'h4248dc46, 32'hc1d2ddb1},
  {32'h44b8c59b, 32'h43853ec0, 32'h4389f00d},
  {32'hc397a3d4, 32'hc3c674d9, 32'hc351136a},
  {32'h450d71b0, 32'hc355599a, 32'hc38de655},
  {32'hc4a16f97, 32'hc304b071, 32'h42a62f99},
  {32'h4502ea6c, 32'hc3b71b67, 32'h4351c893},
  {32'hc3947430, 32'h42c578d0, 32'hc28eb789},
  {32'h4500ab8b, 32'hc2c5f5c9, 32'h43ce7349},
  {32'hc3cbad7d, 32'hc3dede0e, 32'hc2b9401c},
  {32'h450ea94d, 32'h432f72b5, 32'hc3cbc0bd},
  {32'hc4aa214a, 32'hc3ab1fbc, 32'hc2bc6398},
  {32'h449d0a50, 32'hc3033a49, 32'h42f6a668},
  {32'hc2cc3168, 32'hc2e930ef, 32'hc3063629},
  {32'h443b1040, 32'h4348c922, 32'hc2bbd0ad},
  {32'hc42c9550, 32'hc15d7b92, 32'hc4293690},
  {32'h4509461b, 32'h42da06a9, 32'h438bd4d8},
  {32'hc29c14e0, 32'h42f69ac5, 32'h4358f950},
  {32'h44bf41c0, 32'hc2cec2d5, 32'h425999a8},
  {32'hc3a6feb8, 32'h40794620, 32'hc3d96c4f},
  {32'h44ecd244, 32'hc33097eb, 32'hc280da60},
  {32'hc4e94470, 32'hc33e029c, 32'hc3066e84},
  {32'h450ba5e6, 32'h43337b61, 32'h42a774e8},
  {32'hc47072fc, 32'hc3526733, 32'hc20236bd},
  {32'h44eb2524, 32'hc38998b6, 32'h43828ae1},
  {32'hc36e6bb0, 32'hc33e55d6, 32'hc37e356a},
  {32'hc46dcb95, 32'h42104347, 32'hc37d674f},
  {32'h43a6ebb0, 32'h43ac91bd, 32'h4341e0a8},
  {32'hc384fe6e, 32'hc0dff242, 32'hc3bc5a71},
  {32'h445101d4, 32'h4342f88c, 32'hc0121c34},
  {32'hc45cb876, 32'h43122304, 32'hc37657dd},
  {32'h44557e0e, 32'h42c4a04d, 32'h43c48099},
  {32'hc51293b5, 32'h41e2d18c, 32'h432434fb},
  {32'h4297e5b2, 32'h442cb91a, 32'hc219a560},
  {32'hc4cc2f3a, 32'h42dc957b, 32'h42b2de21},
  {32'h4493913a, 32'h3e653480, 32'hc36b4e5a},
  {32'hc4f3a2cb, 32'h435186e0, 32'h4255c55c},
  {32'h443ff50c, 32'h42d5dc48, 32'h43b235ee},
  {32'hc48c947d, 32'h43a1f410, 32'hc318ce77},
  {32'h44b2dc89, 32'h428bc874, 32'h435068ac},
  {32'h42dc7460, 32'h435b733c, 32'hc29e8891},
  {32'h440a6857, 32'h437dba5a, 32'h43929e83},
  {32'hc41a4558, 32'hc2b0fc17, 32'hc0b0038c},
  {32'h4473ef27, 32'h41f7c955, 32'h43668296},
  {32'hc4a7f5de, 32'h41806870, 32'h4326e7d8},
  {32'h44424be3, 32'h428e971f, 32'hc2859a2e},
  {32'hc47ebbc8, 32'h436c1fca, 32'hc3802d1a},
  {32'h443c0f61, 32'h429f5482, 32'h42aa6fba},
  {32'hc2bc6d90, 32'h425f6287, 32'hc35d8bc9},
  {32'h447f439a, 32'hc3055942, 32'hc3164bf9},
  {32'hc400cac4, 32'hc38774c3, 32'h4365a19b},
  {32'h425904e0, 32'h4313532e, 32'h42b693eb},
  {32'hc481f537, 32'hc35a8eac, 32'h42a4fa1f},
  {32'h43dea1fc, 32'hc355d1ea, 32'h43a4d791},
  {32'hc4e4da10, 32'h416da778, 32'hc386d046},
  {32'h44f170f2, 32'hc337af70, 32'hc261118d},
  {32'hc4856d89, 32'hc3225124, 32'hc2bc394a},
  {32'hc39a4453, 32'hc1bff69d, 32'h4360b30b},
  {32'hc4b68cda, 32'hc363f531, 32'hc2b6c309},
  {32'h44042fc9, 32'hc1a7bc9a, 32'h429fdeb3},
  {32'hc4c0cd54, 32'hc3bdc3b8, 32'h43304eed},
  {32'h4447e19c, 32'hc3065952, 32'h409b9692},
  {32'hc4085312, 32'hc22727cd, 32'hc41be817},
  {32'h444e2e51, 32'h436e8933, 32'hc36c43f9},
  {32'hc4694289, 32'hc38ad877, 32'h4300cbcb},
  {32'h4454b964, 32'h435af610, 32'h42a803a7},
  {32'hc4cacfad, 32'h430b2547, 32'h43a56411},
  {32'h440c11ca, 32'h43c87444, 32'hc201bc60},
  {32'hc4e779d9, 32'hc38fbeb2, 32'h42cfb61c},
  {32'h44e93688, 32'hc441c5c5, 32'h42ca17f0},
  {32'h4197cfd8, 32'hc378442b, 32'hc2a1da9a},
  {32'h430f0b40, 32'h430cb181, 32'hc2a0ab17},
  {32'hc4afa2bd, 32'h42ed1952, 32'hc2e446ab},
  {32'h43ab0f38, 32'h4433c8d9, 32'h43a75719},
  {32'hc409a422, 32'h4419af22, 32'hc3148fed},
  {32'h44687aeb, 32'hc3055113, 32'h431e0a71},
  {32'hc4f04946, 32'h440850e2, 32'h43203a79},
  {32'h43b6f7c0, 32'h42e919da, 32'h42bfc182},
  {32'hc44d0fb4, 32'h40be4688, 32'hc3be203a},
  {32'h440d2f34, 32'hc386218c, 32'hc092edb2},
  {32'h42a17e20, 32'hc2e1a45a, 32'h42343fd0},
  {32'h4484e394, 32'h42bedcaf, 32'hc3ae2bc7},
  {32'hc4b305d9, 32'hc29f3311, 32'h432ae278},
  {32'h443cdd67, 32'h43030641, 32'h434ec739},
  {32'hc514dcc8, 32'hc1e0865b, 32'hc40686bd},
  {32'h450ff330, 32'hc3acef79, 32'hc38dccd6},
  {32'hc483adff, 32'hc35ca388, 32'hc38aa85b},
  {32'h44a26331, 32'h42870913, 32'hc20e39cf},
  {32'hc4610230, 32'hc28ac703, 32'hc2bdb8c9},
  {32'h448176df, 32'h43504075, 32'h431ca986},
  {32'hc5029844, 32'hc431ac71, 32'h42ab6865},
  {32'h435d4bcc, 32'hc13e1aaa, 32'h434971c2},
  {32'hc4c9788a, 32'h426ea94b, 32'hc1699599},
  {32'h44f328d6, 32'h43a338b4, 32'hc3826550},
  {32'hc4945436, 32'hc31144ca, 32'hc3baac11},
  {32'h44cef5db, 32'h4329baee, 32'h441a3d01},
  {32'hc4cece5f, 32'h42d3c4f4, 32'h433f2f5a},
  {32'h43ccb0c2, 32'hc2d85f18, 32'h42b0f1f2},
  {32'hc44ffecf, 32'h42bb9745, 32'h432e2430},
  {32'h44f94dcf, 32'hc2de9614, 32'h4318d373},
  {32'hc4fdac4c, 32'hc21793c4, 32'h4394b24a},
  {32'h448ca06c, 32'hc237c7f7, 32'h4348fc9c},
  {32'hc4d870cc, 32'hc2c0c0f4, 32'hc3fbba78},
  {32'h43e6199c, 32'h43a6843c, 32'hc342b6b4},
  {32'hc4056000, 32'h439d88b5, 32'h431d3bcc},
  {32'hc31193a4, 32'hc3e978ca, 32'h43f7e8f0},
  {32'hc4dc21a8, 32'h427903e9, 32'h437a3060},
  {32'h43b56648, 32'hc37ae974, 32'h43a41cf0},
  {32'hc4ddf826, 32'hc355d765, 32'h42730ab2},
  {32'h4503e272, 32'h43a65eaa, 32'hc2125db7},
  {32'hc37bb530, 32'h42b1749c, 32'h442a9277},
  {32'h43f1b330, 32'hc2225670, 32'h432c34a6},
  {32'hc4a91299, 32'h42ec9c2e, 32'h43d4555b},
  {32'hc2971d20, 32'hc366616e, 32'h41df5ef7},
  {32'hc46d67b0, 32'h42bbb419, 32'h434411b1},
  {32'h448fe335, 32'hc3b8456c, 32'hc381d0cb},
  {32'h438b4710, 32'hc35d7c73, 32'hc1187401},
  {32'h44052676, 32'hc28a8ae5, 32'h4250f4e2},
  {32'hc4f52677, 32'hc30bfb80, 32'hc1ac80a6},
  {32'h44ac2a47, 32'hc2b84a76, 32'h43a54a42},
  {32'hc4ff5aaa, 32'h43e13ef4, 32'h42571a29},
  {32'h44e2ccda, 32'h42224814, 32'hc3346fb2},
  {32'hc5024b8a, 32'hc300bb10, 32'h42224ec8},
  {32'h44c4a405, 32'h43533b46, 32'hc30e29e8},
  {32'hc505fe62, 32'hc1dd4542, 32'h43ac6937},
  {32'h44bee4ff, 32'h42b56832, 32'h43499831},
  {32'hc4c651d3, 32'h429c0b36, 32'h42f1c1f6},
  {32'h44e47eb4, 32'h439cfb3b, 32'hc1f7926c},
  {32'hc4b0f66e, 32'hc38f76c0, 32'h436921ae},
  {32'h4354fa50, 32'h4319f3fc, 32'hc309a7f0},
  {32'hc3fa4d80, 32'hc3dd987c, 32'hc2d2642a},
  {32'h43c823b2, 32'hc1ab5287, 32'hc39b89d7},
  {32'hc4c52452, 32'hc35d18fc, 32'hc2db8d41},
  {32'h4511351a, 32'hc34fc37f, 32'hc384e4e9},
  {32'hc3d13d0b, 32'hc40caa9a, 32'hc0f115a2},
  {32'h45178262, 32'h43ceb587, 32'hc317e86e},
  {32'hc400fbc8, 32'hc342c021, 32'h433f051c},
  {32'h4482ea0e, 32'h435f429a, 32'hc28f1d8c},
  {32'hc0e6be00, 32'hc405aeef, 32'h43c7f81b},
  {32'h450544c1, 32'hc38f8f20, 32'hc2b20dfb},
  {32'hc4edcaa3, 32'hc3c656e1, 32'h430437cf},
  {32'h439522ea, 32'hc361dea0, 32'hc3779ad2},
  {32'hc1c23f00, 32'hc03ec920, 32'h428c1012},
  {32'hc4a3ee82, 32'h43858497, 32'hc28a310d},
  {32'h44be0adc, 32'hc3244dab, 32'h423ce7e3},
  {32'hc364e296, 32'hc10d4969, 32'hc3ecfbd0},
  {32'h43153ba8, 32'h4392ca53, 32'h4314adff},
  {32'h435d3e9e, 32'h4397fe8f, 32'hc0d711f4},
  {32'h448afcd5, 32'hc276a798, 32'hc3b45191},
  {32'hc4c0a94f, 32'h440000b3, 32'hc3318bac},
  {32'h44fec16b, 32'hc2cd10a3, 32'h430149e9},
  {32'hc52ac1b4, 32'hc33e6611, 32'h431974f1},
  {32'h4416df62, 32'hc39ad18e, 32'h4315e7ff},
  {32'hc30061b0, 32'hc36dcd86, 32'hc3065889},
  {32'hc141006e, 32'h4365cae4, 32'hc37a7ce0},
  {32'h42b75060, 32'h4358fe10, 32'hc35f1fc4},
  {32'h4412cb6b, 32'hc409a504, 32'h432c70d3},
  {32'hc413537a, 32'h42b67740, 32'h41dadf6e},
  {32'h440a0686, 32'h42675951, 32'hc1609e2c},
  {32'hc10cb800, 32'hc25e1535, 32'hc2747bdc},
  {32'h4503bfbc, 32'hc378500b, 32'hc34e9b55},
  {32'hc49998b6, 32'hc363fc92, 32'h4309ce12},
  {32'h44efc32a, 32'h43c0e7a3, 32'hc31233a6},
  {32'hc4964704, 32'h42a596e2, 32'h42307f94},
  {32'hc2c8fa78, 32'h431980e2, 32'h4187b4b9},
  {32'hc4b4a857, 32'h41e4480d, 32'h43113f7f},
  {32'h44d22394, 32'hc31551fd, 32'hc28599c3},
  {32'h420acac0, 32'hc36f0d68, 32'hbf464d20},
  {32'hc3958160, 32'h419d54a2, 32'h42225f6d},
  {32'hc2e1aec0, 32'hc32b2eab, 32'h43d5667a},
  {32'h44aa855f, 32'hc2b6b2b2, 32'hc3b910cb},
  {32'h42d67ee0, 32'hc2b42671, 32'h43886398},
  {32'h442dd5fe, 32'hc208231e, 32'h42bf2a0e},
  {32'hc3fa16ba, 32'hc38be03a, 32'hc3ebeb69},
  {32'h44bcd988, 32'hc34d3a6c, 32'h42b92eea},
  {32'hc40116b0, 32'hc1fe19c1, 32'h423050cf},
  {32'h4400740e, 32'h424ac21a, 32'h436abe18},
  {32'hc3c5d9c6, 32'hc3862fee, 32'h4318ca67},
  {32'h43e037b4, 32'h4362c398, 32'h4343ecb9},
  {32'hc2b07590, 32'hc31178ef, 32'hc369e481},
  {32'h450b6c91, 32'h42f581cc, 32'hc3803c32},
  {32'hc4a9472e, 32'hc3a7673e, 32'h430df133},
  {32'h450c9374, 32'hc3c57b17, 32'hc1ef6d3c},
  {32'hc4f423be, 32'h41f15988, 32'h43024f0a},
  {32'h41e68b2e, 32'hc2a7957b, 32'h4390936a},
  {32'hc4c98d0c, 32'hc37b2e0c, 32'h43ad72c6},
  {32'h4402b9c0, 32'hc345a223, 32'hc37c7783},
  {32'hc39871a8, 32'h4158affc, 32'h42dcf86f},
  {32'h44cf2112, 32'h43340074, 32'h40a35364},
  {32'hc4f44323, 32'hc0f3f6c4, 32'h438a9f09},
  {32'h44477778, 32'h4345c851, 32'hc2dfbf62},
  {32'hc4b0e2fc, 32'h43ac5e73, 32'hc3630312},
  {32'h450402b7, 32'h43771e08, 32'hc3c14e2d},
  {32'hc50944ce, 32'h43ad469d, 32'hc35f9e6d},
  {32'hc16105c0, 32'hc38a97e9, 32'h43229a68},
  {32'hc4fd19ea, 32'h42c089a7, 32'hbfeb830b},
  {32'h449f2fee, 32'hc29a30e8, 32'h435b435a},
  {32'hc45e92b4, 32'hc3933351, 32'h412f9d72},
  {32'h44fed480, 32'hc28b20ca, 32'hc3bdfbdd},
  {32'hc3ba58f4, 32'h406f19ae, 32'hc28695bb},
  {32'h44c14666, 32'h43a97f25, 32'h4400bde6},
  {32'hc41b989c, 32'h431cc99f, 32'hc2242f13},
  {32'h4482e84c, 32'hc12010f4, 32'h436a149c},
  {32'hc449041c, 32'hc3d9111b, 32'h4385533e},
  {32'h444db148, 32'hc27dc542, 32'hc3a2b25f},
  {32'hc36c82c4, 32'hc319deb8, 32'hc20a17c6},
  {32'h45035c9c, 32'hc3091ab0, 32'hc380082c},
  {32'hc44b7d0a, 32'h42a8e903, 32'h4314f501},
  {32'h43ac622c, 32'hc31913c7, 32'hc12e1584},
  {32'hc4f36778, 32'h42ca6cb3, 32'h42a28e98},
  {32'h44e36667, 32'h41627bf0, 32'h428caa67},
  {32'hc4fd76a1, 32'hc2336dde, 32'h43184163},
  {32'h44dfa08d, 32'h439fc425, 32'hc30542a6},
  {32'hc3d0cd28, 32'h42c393a4, 32'h42bdcbcc},
  {32'h435bbea0, 32'h434d46e4, 32'hc1f351fd},
  {32'hc3be1290, 32'hc42e0579, 32'h42d795d3},
  {32'h428d6232, 32'h440525a2, 32'h43d25f10},
  {32'hc4acb07f, 32'hc3581212, 32'h4291ffcc},
  {32'h44f06960, 32'hc3be8526, 32'h43c37c2b},
  {32'hc50e7d56, 32'hc3c761b0, 32'h414b7b1e},
  {32'h441df004, 32'h4221d950, 32'h42e0355b},
  {32'hc510e8b2, 32'h430e236a, 32'h43910d71},
  {32'h45044f9e, 32'h439c4f7a, 32'h43532314},
  {32'hc48de609, 32'hc3d62c1f, 32'h439b4e4e},
  {32'h4398768d, 32'h42d97366, 32'h43152f54},
  {32'hc50f7f87, 32'h432f18af, 32'h44118da6},
  {32'h439cc390, 32'hc32cc3e5, 32'h433e2b5c},
  {32'hc50a042d, 32'hc28fdc8b, 32'h4286d1b4},
  {32'h43723a78, 32'hc38100fe, 32'h43b40c40},
  {32'hc4dd7af6, 32'h42c224ae, 32'hc1a3d378},
  {32'h44677b1e, 32'h42badee8, 32'hc23bb48d},
  {32'hc3e865b3, 32'hc1a8aa7a, 32'h431caae8},
  {32'h441a03e0, 32'hc38c68fe, 32'h437d7692},
  {32'hc4bebce1, 32'h4325046a, 32'hc2b2e3c4},
  {32'hc332eed8, 32'hc3957008, 32'hc27ace57},
  {32'hc49fe42a, 32'hc278dd3a, 32'hc34d36d0},
  {32'h42782560, 32'hc3315dcd, 32'h422c4cc3},
  {32'hc3ce8ae2, 32'h401e4778, 32'hc36391f2},
  {32'h448c00de, 32'hc2be389c, 32'h43929991},
  {32'hc3e72c30, 32'hc25cb842, 32'hc0cb4108},
  {32'h450d2f67, 32'h4383ff16, 32'h425149c0},
  {32'hc4da6bd9, 32'hc3da1ecb, 32'hc353df1f},
  {32'h43e9bcb0, 32'hc24ecb98, 32'h43297e5a},
  {32'hc43b2d98, 32'h4147595e, 32'hc319fdc4},
  {32'h44b24028, 32'hc355374a, 32'h43360520},
  {32'hc3cf2352, 32'h4347785b, 32'hc3714d6a},
  {32'h44ded51c, 32'h434b9d58, 32'hc3797606},
  {32'hc3c9444c, 32'hc1b811b2, 32'hc2daf573},
  {32'h44933cc3, 32'hc2251068, 32'hc3896370},
  {32'hc43b7c52, 32'h4341b9dc, 32'hc2f16c48},
  {32'h44c04522, 32'hc321bc0b, 32'h4348b23a},
  {32'hc4af328e, 32'h42839ff1, 32'h43b0aafb},
  {32'h448f0596, 32'h434b5d2c, 32'h42aced2c},
  {32'hc4f2fe2a, 32'hc31d63d3, 32'h4376bf5f},
  {32'h44880427, 32'hc3834089, 32'hc2cd3c01},
  {32'hc48e5b06, 32'hc2dce828, 32'h440cbcca},
  {32'h44e5e488, 32'h42a889fe, 32'h42d89bed},
  {32'hc30b37f8, 32'hc318676c, 32'h425da0be},
  {32'h44c987c6, 32'h442f30fb, 32'hc37dab52},
  {32'hc3e06674, 32'hc287dcb7, 32'hc300eacd},
  {32'h44b062dc, 32'h41378cac, 32'h41d0a12e},
  {32'hc49da19c, 32'h42c8db3a, 32'h431b1f11},
  {32'h44a9739a, 32'h426514a4, 32'h42a0d01d},
  {32'hc3c65fa2, 32'h421b68ee, 32'hc25e8e0e},
  {32'h44ebde90, 32'h43841cbd, 32'h42cc79bc},
  {32'hc474265e, 32'hc2fac15b, 32'h426a25f4},
  {32'h44850ec2, 32'h42ba5eb2, 32'hc31a697a},
  {32'hc4e0caf7, 32'hc314b716, 32'h43a228cc},
  {32'h43a84f18, 32'hc3452cae, 32'h41c48840},
  {32'hc5030673, 32'hc293fdf0, 32'h4367af4a},
  {32'h441b13b0, 32'h43b8eec7, 32'h43831d19},
  {32'hc460a138, 32'h428d3ece, 32'hc3aca560},
  {32'h44d038a8, 32'hc383ba5c, 32'h4352ce4c},
  {32'hc51897e8, 32'h4315e76f, 32'hc3bd309a},
  {32'h4440fcf0, 32'h43479e0a, 32'hc354c98a},
  {32'hc4478d38, 32'hc399d596, 32'h433e9ef5},
  {32'h44d818db, 32'h4339986a, 32'h415ca6de},
  {32'hc3d9aa8a, 32'hc40468a1, 32'h41d7b736},
  {32'h44b48c17, 32'h4391fea0, 32'hc1fba836},
  {32'hc4986e62, 32'hc38434af, 32'hc2b9049e},
  {32'h441919d6, 32'h436475fc, 32'h42f10b13},
  {32'h42465280, 32'hc3186158, 32'hc30c6a11},
  {32'h44c7a421, 32'hc3792b52, 32'hc2d70351},
  {32'hc4c413c2, 32'h43c74e2d, 32'hc38fe68d},
  {32'h44252366, 32'h42e0164e, 32'h43186a7c},
  {32'hc409668a, 32'h42ef5892, 32'hc3af205a},
  {32'h4502f8c4, 32'hc178f1b4, 32'h436d5240},
  {32'hc4ab7460, 32'hc3b24307, 32'h42a59e75},
  {32'h445a5da2, 32'hc351a958, 32'hc210f680},
  {32'hc4d05715, 32'h430b9dba, 32'hc2d815b5},
  {32'h44fcacf2, 32'hc385ec61, 32'h43a4186b},
  {32'hc5012129, 32'h42b41d67, 32'hc35f50b9},
  {32'h4402c04e, 32'h430f92c0, 32'h42c0f445},
  {32'hc3d0d630, 32'hc1b144e6, 32'hc26e109c},
  {32'h450a7f10, 32'h42b32867, 32'h42dee143},
  {32'h42fbf720, 32'hc3d77bcb, 32'h429e4076},
  {32'h43afb531, 32'hc31cf00c, 32'hc19737d1},
  {32'hc36199ab, 32'hc25a997c, 32'hc3c5f368},
  {32'h4481103a, 32'h43340f29, 32'hc284b2bb},
  {32'hc466c4fa, 32'hc2a7864b, 32'h433db35a},
  {32'hc30a0600, 32'h432ce06b, 32'hc2fa9fe8},
  {32'hc4e02d2a, 32'hc38c4297, 32'h425fe8e7},
  {32'h4470bfb5, 32'h431abe9f, 32'hc3aa0452},
  {32'hc4e27f00, 32'hc1ffbddf, 32'h42f9e807},
  {32'h443d0249, 32'hc3538fa5, 32'hc31b30a6},
  {32'hc3a0d65d, 32'h425f1cc5, 32'h43472905},
  {32'h45142e7a, 32'h430403c3, 32'hc1ec44c6},
  {32'hc50101e3, 32'h42921ff1, 32'hc337d8bc},
  {32'h449086fc, 32'h42beaa67, 32'hc3ea2c9c},
  {32'hc4ebb4e7, 32'h434776d4, 32'h42f4de66},
  {32'h443ead20, 32'hc24230f0, 32'h42245dfd},
  {32'hc41376e8, 32'h41bd09c6, 32'hc32fd6b4},
  {32'h4440bee7, 32'h42a4cb9f, 32'h43542283},
  {32'hc4eb6679, 32'hc3695ed5, 32'hc2b26566},
  {32'h44d99440, 32'hc3477e74, 32'hc3d446f7},
  {32'h4179d980, 32'hc150b384, 32'hc3043c4a},
  {32'h438d712e, 32'hc28e99d6, 32'h42078936},
  {32'hc3e8c640, 32'hc2bfe56f, 32'hc37f1bb0},
  {32'h44b4f826, 32'hc2dfc5bb, 32'h427eed30},
  {32'hc4b88f28, 32'hc30f1c4c, 32'hc392ad62},
  {32'h42775614, 32'hc2a5eb27, 32'h428f3446},
  {32'hc4c94a0d, 32'h4347f92c, 32'hc3855f67},
  {32'h43bec285, 32'h42a23a4f, 32'h43565ed2},
  {32'hc48b6312, 32'h431285e0, 32'h4326fe86},
  {32'h4514ddac, 32'hc2b69288, 32'h438e0410},
  {32'hc4d90968, 32'h437ff425, 32'hc324d2ff},
  {32'h44d47df8, 32'hc1e8581e, 32'h409c00a3},
  {32'hc4e45fa2, 32'h42887643, 32'h42d20cdd},
  {32'h443731a5, 32'hc31fcd16, 32'hc3b76502},
  {32'hc3bba39e, 32'hc2e76df1, 32'hc26af2e4},
  {32'h450f5601, 32'h43a46226, 32'hc312b5aa},
  {32'hc4bc5ae9, 32'hc1ba8af1, 32'hc384b4ee},
  {32'h442c5443, 32'hc3a0c4f0, 32'hc2d4138b},
  {32'hc4fa7654, 32'hc31a5ca3, 32'h42ce921d},
  {32'h4502cdc2, 32'h42d00ed0, 32'hc3947059},
  {32'hc1e1df80, 32'hc33abfbe, 32'hc3282002},
  {32'h4508a554, 32'h423f3f62, 32'h42e35d37},
  {32'hc3d3b934, 32'hc2824720, 32'h430fbf00},
  {32'h44accb5f, 32'hc1a79fc9, 32'h43828a47},
  {32'hc526054a, 32'hc3e6cfd8, 32'h43213304},
  {32'h44c2c899, 32'h43886d34, 32'hc1dde360},
  {32'hc49e5c32, 32'h43ea7f55, 32'hc3311d22},
  {32'h448e0816, 32'hc276911a, 32'h43107bb9},
  {32'hc4484c1e, 32'h420b43b0, 32'hc1f4f77e},
  {32'h449e61ed, 32'h4351f747, 32'h439fe87d},
  {32'hc41b94ee, 32'hc3706fc8, 32'hc36376dc},
  {32'h44211062, 32'hc26828a1, 32'h42ca4997},
  {32'hc456c4bd, 32'hc2500654, 32'hc3454d17},
  {32'h450a6724, 32'h43b96509, 32'h43cb9774},
  {32'hc3a155a4, 32'hc3ada934, 32'hc3832806},
  {32'h43ceb55c, 32'h438a0254, 32'h42104d02},
  {32'hc4a8d91a, 32'h41124eaf, 32'h43f91270},
  {32'h44f995d5, 32'hc1f21e3e, 32'h424b8f2b},
  {32'hc48ce9f1, 32'h42f6371e, 32'hc3401d20},
  {32'h43d11d38, 32'h43a5335c, 32'hc375290b},
  {32'hc4817a9c, 32'hc3a6fdd5, 32'h42127872},
  {32'hc0691400, 32'hc3905e15, 32'h429fce9c},
  {32'hc3bfbb2e, 32'h4068e938, 32'hc36efb72},
  {32'h4480514a, 32'h4272816d, 32'hc3d645d4},
  {32'hc4992d8f, 32'hc2fcfbf9, 32'hc3e5823b},
  {32'h44bfda35, 32'h428ef0ef, 32'hc2f0d9ed},
  {32'hc3901842, 32'hbf13a030, 32'h4302310c},
  {32'h4203bb40, 32'hc3526701, 32'hc2212721},
  {32'hc5174067, 32'hc3229218, 32'hc383f302},
  {32'h44c4f6e8, 32'hc27a3849, 32'h428d8e3c},
  {32'hc318d470, 32'h42686d04, 32'h439aeb4a},
  {32'h44ea43ae, 32'hc3a3c8cd, 32'hc2630a81},
  {32'hc35c43d0, 32'hc390211b, 32'hc33b8ab3},
  {32'h41044e80, 32'hc3909d5a, 32'h42f13242},
  {32'hc498fde4, 32'hc30161fb, 32'hc4031c04},
  {32'h438bbb54, 32'h42a9c95c, 32'h42b4fb4c},
  {32'hc4b0316c, 32'hc2c82cff, 32'hc1f6488e},
  {32'h45086329, 32'hc39b58ec, 32'hc23c0337},
  {32'hc4563927, 32'h438c655c, 32'h41c6b3b5},
  {32'h44fa0730, 32'h4200631d, 32'hc29671e8},
  {32'hc50e5298, 32'h3fd4bbf0, 32'hc33c8dec},
  {32'h4313f4b8, 32'h43174043, 32'hc3201b13},
  {32'hc4ee1527, 32'hc0c6b998, 32'h43945214},
  {32'h44879f1e, 32'hc1827abe, 32'hc28ba44b},
  {32'hc4e07c12, 32'h41e1df14, 32'hc39adb3c},
  {32'h45234b16, 32'h42db18cc, 32'h4372c214},
  {32'h43553a50, 32'hc2d0036b, 32'h4397fe0f},
  {32'h450fc949, 32'h42f7cdf7, 32'hc3cdf9a2},
  {32'hc50d54a5, 32'h42bba09a, 32'h410505c2},
  {32'h451ca52c, 32'hc27171c8, 32'hc39b9e97},
  {32'hc4f1d2b4, 32'hc3c7b9e2, 32'h41edc239},
  {32'h450cd020, 32'hc39c038c, 32'h41ae5873},
  {32'hc3241ab0, 32'h426c5754, 32'hc3baada3},
  {32'h44b6f9ed, 32'h43e3d5ae, 32'hc2840e94},
  {32'hc49ed669, 32'h3d9cb7a2, 32'h42f8a7ee},
  {32'h44b885f9, 32'hc2ffd728, 32'h4354ab9f},
  {32'hc4cbd2b4, 32'hc0962c20, 32'hc0428698},
  {32'h449ba6a6, 32'h438b2187, 32'hc29d1465},
  {32'hc4a4bf37, 32'hc1b1ddfa, 32'hc3582433},
  {32'h44caae86, 32'h438b6724, 32'h4318ac84},
  {32'h42b82e2b, 32'hc3e2a99b, 32'h4232daed},
  {32'h43fe2eb4, 32'h43ba3952, 32'h4347a5e3},
  {32'hc2e09d20, 32'hc32c04ef, 32'h435178ad},
  {32'h44d4d890, 32'h43291b6e, 32'hc2f0cb58},
  {32'hc4a1fbe9, 32'hc2cd196c, 32'h426c5f01},
  {32'h452d5a42, 32'h42ecef97, 32'hc3c233d2},
  {32'hc49958f2, 32'hc31a8019, 32'hc2f8c1c6},
  {32'h44d43a2c, 32'h420efe57, 32'hc24c7bc6},
  {32'hc50faf12, 32'hc345d81c, 32'hc214668a},
  {32'h44ecd857, 32'h43d200e2, 32'h42a6a469},
  {32'hc48eb655, 32'h43ae67f5, 32'hc3702834},
  {32'h4474e872, 32'h434d0a58, 32'hc2d1a4d9},
  {32'hc3c727b6, 32'h423111fa, 32'h4231e330},
  {32'h44bd6d2b, 32'h415afd68, 32'h40b8c5a9},
  {32'hc50b9ce5, 32'h42b96a6c, 32'h4399fbf0},
  {32'h4479427d, 32'h42d789ee, 32'hc396d7f9},
  {32'hc4e27522, 32'hc4007b58, 32'h432ce894},
  {32'h44a8eb7c, 32'hc082fc78, 32'hc31da5e0},
  {32'hc50bd7ba, 32'hc3201b05, 32'hc3d6892c},
  {32'h4474b5c4, 32'hc369a040, 32'hc2fa1de8},
  {32'hc4e492a4, 32'h42df8137, 32'hc22ff98e},
  {32'h42685a80, 32'h43653b92, 32'hc2b7f11b},
  {32'hc3853134, 32'h42db3645, 32'h42eaf20c},
  {32'h43d414b5, 32'h42e94c34, 32'h434fe694},
  {32'hc5065022, 32'hc381c81d, 32'h4327fa2a},
  {32'h452388c0, 32'h438bc849, 32'hc388625d},
  {32'hc12dd3b8, 32'hc324da83, 32'h431b1f1d},
  {32'h445fbd82, 32'h428bacdf, 32'hc362fd2e},
  {32'hc481e512, 32'hc3727b4f, 32'h4266e4b7},
  {32'h44abbbfc, 32'h438d8389, 32'hc396e633},
  {32'hc3de91b4, 32'hc3a9354d, 32'h4345b7f2},
  {32'h445a3baa, 32'hc2b6182d, 32'h4340f7fa},
  {32'hc483828f, 32'h435e368f, 32'hc0941a60},
  {32'h43c5add7, 32'hc3958c41, 32'hc2744760},
  {32'hc48494d1, 32'h405fdc2c, 32'h42fc1432},
  {32'h44e3a393, 32'hc283db20, 32'hc2a363c6},
  {32'hc4357696, 32'hc265f23f, 32'hc160d64e},
  {32'hc26c7b20, 32'hc2c9440b, 32'hc2d8eb06},
  {32'h425aede8, 32'h42e48ad6, 32'hc331d55d},
  {32'h4409af66, 32'hc3bf5421, 32'hc2a6a9f5},
  {32'hc4b26ae2, 32'h4304f38d, 32'h42e1ab30},
  {32'h4500adf6, 32'hc1d5ec8c, 32'hc316c211},
  {32'h433915c4, 32'h4249fca9, 32'hc3175f03},
  {32'h44496097, 32'hc3d4f731, 32'hc388a7e4},
  {32'hc372d268, 32'h43a113c8, 32'h437f981f},
  {32'h428347b2, 32'h424ffb38, 32'h43500d05},
  {32'hc484cc9e, 32'h437a8900, 32'h43b36d5a},
  {32'h44f2ef42, 32'hc0d4dc47, 32'hbf206c22},
  {32'hc4ab6ade, 32'hc28b118a, 32'h43445ea6},
  {32'h4346ea68, 32'h43d6b546, 32'hc3b3b94f},
  {32'hc39be2d0, 32'hc33fccc3, 32'h434924b2},
  {32'h444aa596, 32'h43167274, 32'hc30edd49},
  {32'hc4b2886e, 32'hc21fd9b6, 32'hc2b5bd76},
  {32'h44e34128, 32'hc393425e, 32'hc0584ce2},
  {32'hc3bef5be, 32'h42cd7c0a, 32'h431daf76},
  {32'h44449610, 32'h420d51ae, 32'hc3809ebc},
  {32'hc47b3de6, 32'hc17e06a1, 32'hc3330315},
  {32'h4513d26c, 32'hc2cbf724, 32'hc379e37e},
  {32'hc4afc7c2, 32'hc33a2989, 32'h439d64e9},
  {32'h44b1991e, 32'h431beb8a, 32'hc2aa281b},
  {32'hc48fe2e8, 32'hc25b833a, 32'h43a55793},
  {32'h445afd83, 32'h438dded5, 32'hc2d7f470},
  {32'h43a2ff43, 32'hc31d0989, 32'hc3f2845b},
  {32'hc4bae12a, 32'h43088be0, 32'hc4264eac},
  {32'h44ded4c1, 32'hc38a2b12, 32'h4380b55d},
  {32'hc473dffc, 32'hc3620944, 32'hc3349ce6},
  {32'h45017aec, 32'hc26c7df3, 32'hc3854728},
  {32'hc4e0b85b, 32'h43187e82, 32'hc1a3c4a9},
  {32'h44954122, 32'hc367a3c9, 32'hc306cb2f},
  {32'hc4d3ca4a, 32'h430122ba, 32'hc3aaaf1c},
  {32'h44835d65, 32'hc2ef985e, 32'hc2e7018e},
  {32'hc4aa2667, 32'h43be49a4, 32'hc294aeee},
  {32'h4420b85b, 32'h424dd1f0, 32'hc301e9a9},
  {32'hc4e19e3d, 32'hc2c50b02, 32'h4225ba05},
  {32'h44b2dd6f, 32'hc38caf05, 32'hc3ccc512},
  {32'hc4d6d478, 32'h4346a654, 32'h4215898a},
  {32'h43f14e7c, 32'hc2c0581d, 32'hc1858351},
  {32'hc51bdfa9, 32'h439a85c4, 32'h438fbd1b},
  {32'h449a4972, 32'hc3739464, 32'hc3240335},
  {32'hc50a688d, 32'h431e90c3, 32'hc35f3923},
  {32'h44c38cfe, 32'h4321fa95, 32'hc29fb426},
  {32'hc501f627, 32'hc25e38a2, 32'hc2fd1077},
  {32'h44d228e0, 32'h43b68aca, 32'h438e2a1d},
  {32'hc517ea91, 32'h440a2248, 32'h426ec0fc},
  {32'h43e8068e, 32'hc20def91, 32'hc3443baf},
  {32'hc3f0e5d2, 32'hc386edfa, 32'h431d3c05},
  {32'h44b70660, 32'hc366dad8, 32'hc382fa54},
  {32'hc41c4a0a, 32'hc31fabd4, 32'h437a064a},
  {32'h441367f1, 32'h42e67384, 32'h41fa13fc},
  {32'hc46d778c, 32'h43a0c025, 32'hc3d38229},
  {32'h4457fc17, 32'hc2888de0, 32'h41e6aeb2},
  {32'hc4fde8d2, 32'h436d5f75, 32'h43c84b5a},
  {32'h4494bdc0, 32'hc1c6fe39, 32'h437e3df8},
  {32'hc4e82d99, 32'hc392d814, 32'h429573b9},
  {32'hc2a6ba1c, 32'h42a0ba80, 32'hc384d8d5},
  {32'hc3a5671c, 32'h42b8d06e, 32'h41d5e5e0},
  {32'h44d71f79, 32'h42bc930e, 32'hc38372b1},
  {32'hc4d19125, 32'h438145eb, 32'h431a654e},
  {32'h44ed0501, 32'hc339e88a, 32'hc29d7cd6},
  {32'hc4dad633, 32'h42fb93d4, 32'h429a44eb},
  {32'h449619c5, 32'hc2d141fb, 32'h435cad2a},
  {32'hc4ae3c3e, 32'h430131c7, 32'hc3cfb282},
  {32'h44d44743, 32'hc334c187, 32'h401bfcba},
  {32'hc3cb7877, 32'h43811d59, 32'hc32ee094},
  {32'h43f3302e, 32'hc38b7a92, 32'h43015541},
  {32'hc5185f31, 32'hc33a30af, 32'h430bbb9c},
  {32'h4517a09b, 32'h43546063, 32'hc18fd78a},
  {32'hc4fb84d1, 32'h436dbba8, 32'h4388af0b},
  {32'h4489b75d, 32'h431a0833, 32'h43453195},
  {32'hc5164e9e, 32'h42f37828, 32'hc26caf40},
  {32'h44d75649, 32'h43963426, 32'hc338c134},
  {32'hc29cb31a, 32'h40e214f0, 32'h43933c00},
  {32'h4419bfb0, 32'hc3328e4a, 32'h4279b83a},
  {32'hc49c5cef, 32'hc2bc4e56, 32'h43a7d58b},
  {32'h4457e9b0, 32'h429e68dd, 32'h434538ea},
  {32'hc4565af5, 32'hc2c71853, 32'h41f24b7e},
  {32'h444da341, 32'hc1003e5e, 32'hc37920d2},
  {32'hc488f266, 32'hc329f266, 32'hc3f1572b},
  {32'h4456f9cb, 32'h440dfc64, 32'h42934640},
  {32'hc48476ca, 32'hc33e8caa, 32'hc3a2bb96},
  {32'h452e7747, 32'hc34f5aea, 32'hc3519b6f},
  {32'hc4d86444, 32'hc2b3b375, 32'hc2cd70f5},
  {32'h443fddb4, 32'hc3ed28d8, 32'hc24afdb0},
  {32'hc4c640bc, 32'h4383520e, 32'hc2d54bc3},
  {32'h44f60a62, 32'hc3b6bdbe, 32'hc2ddf7fc},
  {32'hc48cb6ab, 32'h438c862b, 32'hc212db88},
  {32'h4336b612, 32'hc1f183de, 32'h438f7dbd},
  {32'hc4ddb33a, 32'h44079621, 32'hc4054ade},
  {32'h43a4c250, 32'hbd740200, 32'h421d8fc7},
  {32'hc45cac02, 32'hc3edbec7, 32'h43aac312},
  {32'h44ec0f3e, 32'h43e55d6f, 32'h4213c688},
  {32'hc506b993, 32'h412d2ce4, 32'h437f5987},
  {32'h45172c5c, 32'h437c58d7, 32'hc38ad07e},
  {32'hc442281e, 32'hc366159e, 32'h4386de13},
  {32'h44b1dfa0, 32'h438ebf2e, 32'hc2870c6c},
  {32'hc50edba8, 32'hc11943d5, 32'hc20b5d9e},
  {32'h4470e8c9, 32'hc326b5c8, 32'h42fffb95},
  {32'hc4e4117f, 32'hc2e3572c, 32'hc2f79063},
  {32'h4511e7f1, 32'h42f7654a, 32'h436a3481},
  {32'hc4ef51e3, 32'h428745d4, 32'hc40946d7},
  {32'h43eb1242, 32'hc2f6f9b4, 32'hc123b4c8},
  {32'hc4f3c9ff, 32'hc2523f58, 32'hc21d6756},
  {32'h44f8d107, 32'hc353a032, 32'h43e000eb},
  {32'hc500f234, 32'h43dd613d, 32'h42b75500},
  {32'h4412d135, 32'h43c47dcb, 32'h42927562},
  {32'hc499f01e, 32'hc1fb0932, 32'hc31a1a70},
  {32'h44a6eb74, 32'h4302663d, 32'h429ef054},
  {32'hc26352af, 32'hc22f0f45, 32'hc0173506},
  {32'h446bd57b, 32'hc306aa75, 32'hc296e058},
  {32'hc4cfbe64, 32'hc33dd45d, 32'hc23914b5},
  {32'h4404b3f6, 32'h43158680, 32'hc32c5d2a},
  {32'hc3b5fd48, 32'h43b36448, 32'hc35d596d},
  {32'h449d1208, 32'h43c46b6a, 32'h43840fb4},
  {32'hc3729e10, 32'hc3b2cb70, 32'h42af27d4},
  {32'h43fd9f1a, 32'hc3725e0f, 32'hc34fe623},
  {32'hc4d3ef8a, 32'hc257d24e, 32'hc3a4e6d4},
  {32'h4496ff5d, 32'h42fb7983, 32'hc3aa4bcf},
  {32'hc3041f60, 32'hc35f0bb8, 32'hc3291199},
  {32'h4477cdc8, 32'h42a5cd43, 32'h43906b45},
  {32'hc253cb80, 32'h4418b9dc, 32'hc2b699a3},
  {32'h4528926c, 32'hc32c8b7e, 32'hc2160791},
  {32'hc44e7f1b, 32'h43590505, 32'h431c8d59},
  {32'h44c1ac33, 32'h43e09bab, 32'h4392bce7},
  {32'hc4bfa8f5, 32'h41e73706, 32'h43744b02},
  {32'h44bca01d, 32'h42ac0a3e, 32'h43e1dad8},
  {32'hc393434f, 32'h43472d58, 32'h431ebe96},
  {32'h4485758b, 32'hc315c21e, 32'hc2a6cd9c},
  {32'hc4c40651, 32'hc18c4ce7, 32'h439a0d4a},
  {32'h4516e629, 32'h437f287e, 32'hc3597e81},
  {32'hc435fa48, 32'hc333eb21, 32'h42feb117},
  {32'h441bf129, 32'h42e18eab, 32'hc2cbb8ce},
  {32'hc326bfc8, 32'hc2ac478e, 32'h42369525},
  {32'h441549d6, 32'hc2ae864e, 32'hc2bfbd7b},
  {32'hc4eb5d5e, 32'hc3b9e1ea, 32'hc173209e},
  {32'h44fe4c92, 32'hc31d050b, 32'hc1cb9b24},
  {32'hc51b6a1a, 32'hc2e91485, 32'h42375a3e},
  {32'h43f0714b, 32'h43f8df04, 32'h42ea329d},
  {32'hc41573b4, 32'hc3393ec7, 32'hc21b027b},
  {32'h44b34cc0, 32'h4271f771, 32'h43483a0f},
  {32'hc3b726af, 32'hc32bcf6a, 32'hc3871eb2},
  {32'h44a76c93, 32'hc1020f0b, 32'h42bf7951},
  {32'hc4945892, 32'h42c24a8c, 32'h43163292},
  {32'h4515dfe6, 32'h42afb28d, 32'hc2e8baca},
  {32'hc44c30c8, 32'h43a50771, 32'h43162210},
  {32'h4507ebb5, 32'hc3d9e8d5, 32'h4349ad48},
  {32'hc49774b8, 32'h43cc71f0, 32'h4314312b},
  {32'h44c5e792, 32'h42acf166, 32'hc332d56d},
  {32'hc3af72de, 32'h43f8ec27, 32'hc2b533be},
  {32'h4506a838, 32'hc383ac47, 32'hc3428b55},
  {32'hc4b34182, 32'h42e4a351, 32'h41936279},
  {32'h438c7196, 32'hc3cae43c, 32'hc1c70397},
  {32'hc51ab650, 32'hc1ce7832, 32'h434d18ad},
  {32'h45089580, 32'h425af147, 32'h42c78248},
  {32'hc41be49e, 32'hc254a78a, 32'h42d28dba},
  {32'h43e9d798, 32'h435c501f, 32'h4341f4da},
  {32'hc3be0a22, 32'hc1b1069a, 32'h43080a56},
  {32'h4493f10d, 32'hc22012d7, 32'h42ef1b5d},
  {32'hc4a8ee68, 32'hbfb61ed0, 32'hc3029fc3},
  {32'h44c349d0, 32'h43a04e2e, 32'h42c2b3da},
  {32'hc4ed9fcf, 32'h43c3ec1b, 32'h433bfaf8},
  {32'h447b411b, 32'h4265a848, 32'h43aa0634},
  {32'hc47b9934, 32'h4201e632, 32'h40cb7f1e},
  {32'h42cd5be8, 32'hc3e7e719, 32'hc1aa1632},
  {32'hc500c658, 32'h41dc67ec, 32'h43bd4e51},
  {32'h4393c6d8, 32'hc39b2caa, 32'h42c76fe4},
  {32'hc2b38e00, 32'h43d1b508, 32'hc3581112},
  {32'h44b56849, 32'h432d3589, 32'h43672a86},
  {32'hc3b659c8, 32'hc2eab7e2, 32'hc32115e3},
  {32'h44115032, 32'h4211cd8e, 32'h439d5d9b},
  {32'hc4a9d73c, 32'h42e33b51, 32'h43879639},
  {32'h44e0ceb3, 32'h42b1978a, 32'h427841b8},
  {32'hc405a8db, 32'hc346c75b, 32'hc3705371},
  {32'h446b14fa, 32'hc2f44db7, 32'hc17a8b99},
  {32'hc46c3c80, 32'hc344e05f, 32'hc293e886},
  {32'h44ebb351, 32'h43b3b1a8, 32'h42ed7c30},
  {32'hc504cc58, 32'hc3d6ab8e, 32'hc33a6d53},
  {32'h44b4a951, 32'h43d4ed31, 32'h4397e42b},
  {32'hc4fc6123, 32'h4264336e, 32'hc2298906},
  {32'h45069000, 32'hc23f6e89, 32'hc3a2acba},
  {32'hc4f356f3, 32'hc3a25489, 32'hc36f9997},
  {32'h445e0398, 32'h42b03f67, 32'h428228ce},
  {32'hc4a48a46, 32'h43d523c9, 32'h4243e1ea},
  {32'h44f80031, 32'h431bf802, 32'h4259a3a3},
  {32'hc4704f0b, 32'h424be75b, 32'hc2ed8860},
  {32'hc3672f48, 32'h43781c2c, 32'h434766ca},
  {32'hc5188aa2, 32'h42ca3fa7, 32'h43151ea8},
  {32'h450c51db, 32'h42a14bc6, 32'h42c60235},
  {32'hc4f4b262, 32'hc05cdcf5, 32'h423182d8},
  {32'h44bc953d, 32'h43857449, 32'hc36b1c25},
  {32'hc4ade228, 32'hc35307b9, 32'h43a779cb},
  {32'h45196510, 32'h4370d10b, 32'hc29682e4},
  {32'hc40283c6, 32'hc31f33de, 32'h41dc81bd},
  {32'h44c686cc, 32'h431922ea, 32'h43321598},
  {32'hc494d3fa, 32'h42f76199, 32'hc35ac64a},
  {32'h44ae1100, 32'hc2b57718, 32'hc33eaec2},
  {32'hc4df2089, 32'hc3880db7, 32'h42b4413d},
  {32'h450144ba, 32'hc10f2ae6, 32'h433789b2},
  {32'hc4b38aa9, 32'hc1dab2dc, 32'hc306b1c3},
  {32'h448059ff, 32'h42aefaad, 32'h42ec068c},
  {32'h43822438, 32'hc2b279a8, 32'h43b57861},
  {32'h44164944, 32'hc3953723, 32'hc2722605},
  {32'hc39c28a0, 32'hc358368d, 32'h431aa3a1},
  {32'h44bcadf5, 32'h41b8d488, 32'hc3c6b5dd},
  {32'hc19da468, 32'h42f4cf16, 32'hc3298f56},
  {32'h44efad47, 32'hc1d0ad49, 32'h42bf5129},
  {32'hc4d9097c, 32'h428217ba, 32'hc2f9e478},
  {32'h44d3f9c4, 32'hc1b4d3a2, 32'h43118492},
  {32'hc4e44baf, 32'h4321d8ec, 32'h4319eac6},
  {32'h449d1217, 32'hc263779e, 32'hc385d5d3},
  {32'hc2941658, 32'h43c78d12, 32'hc23b0ec2},
  {32'h443d1722, 32'h42abb287, 32'h43974cdc},
  {32'hc504a2b0, 32'h433bd76f, 32'h42fe5345},
  {32'h4510d67f, 32'hbf13d50a, 32'h42d91326},
  {32'hc4420cba, 32'h43019937, 32'hc2edf72e},
  {32'hc3144c50, 32'h42a8d793, 32'hc384f31c},
  {32'hc511d514, 32'hc39c0818, 32'hc3483fe6},
  {32'h448814e6, 32'hc2514976, 32'hc27048b5},
  {32'hc3daf8ef, 32'h43cfd9f8, 32'hc2b152ab},
  {32'h44a909d8, 32'h43207d24, 32'h43051ce4},
  {32'hc4bc67a6, 32'h42365b5a, 32'h42b96308},
  {32'h43eb06c2, 32'hc36f98fe, 32'hc233f8b1},
  {32'hc4833850, 32'h425ea0c8, 32'hc2dafc14},
  {32'h446c3626, 32'h433a77c9, 32'h43bc708e},
  {32'hc4877ec9, 32'hc3249a10, 32'h4288e59d},
  {32'h44c21971, 32'hc32805c8, 32'hc3035514},
  {32'hc48cb8f0, 32'hc3210800, 32'h4283fce5},
  {32'h447589a6, 32'hc40f2dda, 32'h43ba77f0},
  {32'hc4c23482, 32'h43029bdf, 32'hc02c3534},
  {32'h44e4f8fe, 32'h4319c498, 32'hc2afbe44},
  {32'hc500a854, 32'h4221aede, 32'hc3bf7aa2},
  {32'h44deb95a, 32'hc34d810d, 32'h42b524cc},
  {32'hc516e7c5, 32'hc32c5408, 32'h438f3bac},
  {32'h44d9b4f9, 32'hc3b8f604, 32'hc32effd0},
  {32'hc44136e4, 32'h41cfca36, 32'h43930781},
  {32'h44529f94, 32'h41bbea42, 32'hc3a637c0},
  {32'hc4e84246, 32'h428aed5c, 32'h439b3354},
  {32'h4454ff03, 32'h43589757, 32'h42dc1414},
  {32'hc4f30093, 32'hc293d89a, 32'hc36fac68},
  {32'h44be5c88, 32'hc2e4e002, 32'hc3b157e4},
  {32'hc396a600, 32'hc2c10a10, 32'hc2eccc92},
  {32'h449d77f0, 32'hc313fd7d, 32'hc18b90cc},
  {32'hc501e0dc, 32'h437812fb, 32'h43c9d8a8},
  {32'h44dd5aac, 32'hc2fa3d69, 32'hc302fd13},
  {32'hc2328d46, 32'h434696b1, 32'h43a9a851},
  {32'h440bad70, 32'hc30829fd, 32'h413b8b39},
  {32'hc3819a88, 32'h41349477, 32'h42a4bb69},
  {32'h44871425, 32'h43337c27, 32'hc3285036},
  {32'hc5029243, 32'h430e3b0c, 32'hc33fbfb2},
  {32'h4449179e, 32'h43b99969, 32'hc3e1cbba},
  {32'hc42e0c4f, 32'hc37246ea, 32'hc39ddaa7},
  {32'h43bc8dbc, 32'hc2048cdc, 32'h4217f164},
  {32'hc2775df8, 32'hc3163aa7, 32'h4265ab17},
  {32'h448b3092, 32'h43a5849d, 32'hc3438859},
  {32'hc48f91ec, 32'h43221b84, 32'hc30995f7},
  {32'h44cb75d8, 32'hc2e4b99d, 32'hc3a73218},
  {32'hc4852864, 32'hc2618dc2, 32'h40cb1f60},
  {32'hc377d696, 32'h42975c04, 32'h42eb1fb0},
  {32'hc3ed1788, 32'hc1b851d9, 32'hc2ca65a1},
  {32'h44b70327, 32'h434b27ce, 32'h43033755},
  {32'hc417d958, 32'h4334599c, 32'hc2482163},
  {32'h44e43f1a, 32'h42f7acc9, 32'h43895629},
  {32'hc5030e27, 32'hc2d05e2b, 32'hc32508ce},
  {32'h4508f690, 32'h43c1eb1d, 32'hc419c68c},
  {32'hc4897c82, 32'hc31d4312, 32'h42cb51c2},
  {32'h44c6ad9f, 32'hc2e0882a, 32'h428fa01e},
  {32'hc48a3c9c, 32'hc26e2512, 32'h4308e69b},
  {32'h44fde759, 32'h4383174b, 32'h429b2869},
  {32'hc4fbffe8, 32'hc3141d20, 32'hc205a143},
  {32'h44f4a885, 32'hc1bc2236, 32'hc3c05ac2},
  {32'hc507a42b, 32'hc20c60c6, 32'h43b1c9b3},
  {32'h448af5b9, 32'hc20451a2, 32'h42f8e9af},
  {32'hc3dd0f4b, 32'hc3a11ec9, 32'h434b6939},
  {32'h4508365b, 32'h4338ea74, 32'h43708a3b},
  {32'hc4df563b, 32'h42d64c6f, 32'hc0e0b5f1},
  {32'h44b565f8, 32'hc235caa9, 32'h43e82c85},
  {32'hc4b0a85d, 32'hc3195e28, 32'hc2b8f82e},
  {32'h44f56e51, 32'h435d5b28, 32'h428ae3b0},
  {32'hc4e5b193, 32'hc2315301, 32'hc3bc346e},
  {32'h449dc081, 32'hc30b125c, 32'hc28b5af6},
  {32'hc40b7a60, 32'h434724d1, 32'h42827fb7},
  {32'h448478bd, 32'h42c3fee4, 32'h4220f346},
  {32'hc505b854, 32'h403d6d68, 32'hc141dc3d},
  {32'h451a460f, 32'h42b5ed3d, 32'hc1a5a139},
  {32'hc262d6c0, 32'h43907327, 32'hc0d8efb5},
  {32'h44c64cef, 32'hc2839521, 32'hc300f765},
  {32'hc4668a66, 32'hc3900679, 32'h44027c8b},
  {32'h4482fcaf, 32'hc24259fb, 32'h401c8f31},
  {32'hc5003f06, 32'hc3634b83, 32'h41c5d720},
  {32'h444b5268, 32'h41b3298c, 32'hc32f6ddf},
  {32'hc432bf8a, 32'h4404b1d2, 32'h42d0fd3f},
  {32'h44b630e0, 32'hc2be0402, 32'hc2b648f4},
  {32'hc4a2169c, 32'hc3c068ba, 32'hc31a12cc},
  {32'h43995600, 32'hc2c7ac33, 32'hc2ed8479},
  {32'hc4189255, 32'h42a1b58f, 32'h43091a60},
  {32'h44cbb0ec, 32'hc2f7de36, 32'hc3d0761e},
  {32'hc394d304, 32'hc300c693, 32'hc3518e71},
  {32'h4344c1c8, 32'hc4041ab7, 32'hc35c3e9d},
  {32'hc5065a8b, 32'h43e9441f, 32'hc1f9c651},
  {32'h4437fcc7, 32'h42cfdd47, 32'hc14c1bf0},
  {32'hc4e9a0dd, 32'hc30c2aaa, 32'h425b7127},
  {32'h438ae108, 32'h43c4cd78, 32'hc3d7bb69},
  {32'hc4ac1dde, 32'h43189cdb, 32'h41ce2986},
  {32'h448dd5b9, 32'h43a70281, 32'hc2642ca7},
  {32'hc4810d82, 32'hc3948cf5, 32'h429939b5},
  {32'h4310d450, 32'hc03957f9, 32'hc26ac794},
  {32'hc3a6d1f0, 32'hc3682d82, 32'h42ac5058},
  {32'h4485ffbc, 32'hc382b2b7, 32'hc2961592},
  {32'h42575b80, 32'hc015e308, 32'h428f6496},
  {32'h44265e11, 32'hc2bfb1f6, 32'h439473bb},
  {32'hc492049e, 32'h439c86c5, 32'hc25b7e5e},
  {32'h436857f0, 32'hc3bc0904, 32'hc12c7150},
  {32'hc4691a1a, 32'h43814c2a, 32'hc1721647},
  {32'h432c384c, 32'hc27e0e81, 32'hc29d0db8},
  {32'hc4b3510a, 32'h4372ace6, 32'hc2cc625b},
  {32'h44c69e3b, 32'h42296f13, 32'hc2bbdd9a},
  {32'hc4bcd2a8, 32'hc3d7b5f2, 32'h42640a5c},
  {32'h43dcdd48, 32'hc33c50c7, 32'hc37f7b8f},
  {32'hc4db4fec, 32'hc2b5facd, 32'h432ffb75},
  {32'h44f20faa, 32'h42c2e157, 32'hc1fe23e8},
  {32'hc2f1b50a, 32'h4334b90f, 32'h439a95ba},
  {32'h44bd5d92, 32'h43b55154, 32'hc33fc2c4},
  {32'hc487e9a8, 32'hc2b17b09, 32'h429d35a6},
  {32'h45096bb2, 32'h43a52a5c, 32'hc37ca1e8},
  {32'hc4e9eff5, 32'hc267b161, 32'hc3e2d9b3},
  {32'h44ffee84, 32'h421ba5fc, 32'hc0f7cfb1},
  {32'hc4c019f4, 32'h42f75034, 32'h4136572c},
  {32'h44095690, 32'h42817b9c, 32'hc38b871e},
  {32'hc4284b60, 32'hc33db816, 32'h43657723},
  {32'h451b3e68, 32'h438e08e4, 32'hc40a9bb9},
  {32'hc485b2f2, 32'hc2d916b2, 32'hc27dafad},
  {32'h44ade330, 32'h437aa6ff, 32'h42e2cae2},
  {32'hc4f90e09, 32'h40cf3f34, 32'h43739a66},
  {32'h4363689d, 32'hc39c85d9, 32'hc31a1d8d},
  {32'hc4906da6, 32'h438762da, 32'h4217a569},
  {32'h450579b5, 32'h429299ee, 32'h4197fe48},
  {32'hc4e1a97f, 32'hc31f41c8, 32'h4392d3ad},
  {32'h44f98b52, 32'h4401632c, 32'h42937d4c},
  {32'hc4ab732a, 32'h4370cb33, 32'h43a21b57},
  {32'hc2d9c788, 32'hc2de2e4c, 32'hc36e788d},
  {32'hc4eda6f4, 32'hc30a12d6, 32'hbf3ed874},
  {32'h441532fc, 32'h42b916ec, 32'h40b1add4},
  {32'hc4f38358, 32'h431d06e8, 32'hc39f9aa6},
  {32'h4494d5d2, 32'h434cdaca, 32'h4384dabb},
  {32'hc4e3780a, 32'h43802efb, 32'hc38ef95c},
  {32'h4405a267, 32'hc31a6f75, 32'h435e864e},
  {32'hc50fdc2d, 32'hc2a8459d, 32'h4318119c},
  {32'h4475a14f, 32'hc3a3495a, 32'hc34ed302},
  {32'h4362aa3b, 32'h4310730e, 32'h43875067},
  {32'h449a42c6, 32'hc3acd388, 32'h42e84fee},
  {32'hc4e39cc2, 32'h43340336, 32'h42cf386d},
  {32'h4399e288, 32'hc38e61ff, 32'hc3736a6e},
  {32'hc329a0d0, 32'h41fb43c5, 32'hc32f4734},
  {32'h450c7bf2, 32'h435d5e47, 32'h43da8a17},
  {32'hc4b50f02, 32'hc2788ede, 32'hc21e7ca4},
  {32'h4420df74, 32'h4305364f, 32'hc36b78d5},
  {32'hc41c72e1, 32'h412ceb01, 32'hc3a4109f},
  {32'h45034eb4, 32'h42eb5f08, 32'hc1eb577b},
  {32'hc5048a57, 32'hc3be2bb6, 32'hc381db21},
  {32'h440328a4, 32'h4331b8c2, 32'h4378fad1},
  {32'hc4cfd966, 32'h429aa813, 32'hc2f2bc03},
  {32'h44d82d40, 32'h42f202aa, 32'hc158f07b},
  {32'hc3546438, 32'h42f4d994, 32'hc394cb7a},
  {32'h4328b660, 32'h43514c24, 32'hc2fbf29e},
  {32'hc4c8b61f, 32'h41ea237b, 32'hc39d7bd5},
  {32'hc0df9bc0, 32'h433543d2, 32'hc38c9013},
  {32'hc3c81788, 32'hc282e68c, 32'hc2350479},
  {32'h4416a3e0, 32'h4293f13e, 32'hc1f01908},
  {32'hc35c5f60, 32'hc3339575, 32'hc3656368},
  {32'h439a11d0, 32'hc2e6d9a8, 32'h417f5f41},
  {32'hc4269d1e, 32'hc28b60b7, 32'h43a26f7f},
  {32'h43315544, 32'hc2cc809d, 32'hc31d0fc6},
  {32'hc4d71a3f, 32'hc3b4e5b5, 32'h43248207},
  {32'h44e1e6ca, 32'hc1c9d8b0, 32'h43576693},
  {32'hc50e811b, 32'hc320ec47, 32'h436376ab},
  {32'h44e2e66b, 32'h42d92535, 32'hc38c6bfc},
  {32'hc41533e4, 32'hc2519808, 32'hc393de2f},
  {32'h453a3abc, 32'hc4235646, 32'h432bcd45},
  {32'hc4584190, 32'hc36615c6, 32'h42d7629d},
  {32'h44566342, 32'h434f76bc, 32'hc2caf414},
  {32'hc4e5f50a, 32'h41da7b52, 32'hc37f695e},
  {32'h44ce5bb1, 32'h434793bd, 32'h430ae8ea},
  {32'hc51b3f36, 32'hc36625d0, 32'hc09fa1d4},
  {32'h44d3b318, 32'h42f9a997, 32'h43a6d6b3},
  {32'hc424e204, 32'h42b0a22e, 32'hc286e150},
  {32'h438810c0, 32'hc3a123e8, 32'hc412c204},
  {32'hc433cc59, 32'h41906ade, 32'h430221e0},
  {32'h44723748, 32'hc39137c2, 32'hc354126e},
  {32'hc3ce0bf0, 32'h43d572cb, 32'hc33c4576},
  {32'h4457c2f6, 32'hc4123998, 32'hc2ebf7aa},
  {32'hc50540b6, 32'h43d58f9c, 32'hc131da9d},
  {32'h44a393af, 32'h415dd5b6, 32'hc387d359},
  {32'hc502b391, 32'hc2aff946, 32'h42cb137e},
  {32'h452248ff, 32'h43802dbd, 32'hc26cc0f8},
  {32'h42d6a008, 32'h429c235b, 32'hc3685458},
  {32'h4429f304, 32'h418724ea, 32'hc2d7fcc7},
  {32'hc5072112, 32'hc344efb0, 32'hc2809b83},
  {32'hc316c820, 32'h438aadab, 32'h42ec9fb0},
  {32'hc4e157b6, 32'hc142fa1c, 32'hc26762ee},
  {32'h44acd9d2, 32'h432fe857, 32'hc2a3c1a4},
  {32'hc4cdf02f, 32'hc2eefaf8, 32'h405526a1},
  {32'h451513cf, 32'h43567ba7, 32'h436ef89b},
  {32'hc4a73f10, 32'hc38c8e34, 32'hc32d955b},
  {32'hc26d5be0, 32'hc25c57df, 32'hc36bdd01},
  {32'hc4c795d0, 32'hc35f386f, 32'hc2634a81},
  {32'h45021a1f, 32'hc3945a81, 32'h4370bc5d},
  {32'hc513d4d1, 32'hc292dc30, 32'h43f07dfd},
  {32'h4481ac9e, 32'h41534f80, 32'h436b6ef8},
  {32'hc4b257b2, 32'hc2cc5c42, 32'hc2fa3cc3},
  {32'h4514c589, 32'hc2a132aa, 32'hc303e074},
  {32'hc34ebb60, 32'hc40fe929, 32'h42aa67ce},
  {32'h4415cd5b, 32'h43213126, 32'hc305adbb},
  {32'hc4c1d85e, 32'h438a4ebe, 32'h43aab8e2},
  {32'h4321e8f8, 32'h43288ecd, 32'hc393519c},
  {32'hc5115f54, 32'hc18f664a, 32'h434642ac},
  {32'h443cd9e1, 32'h431a0612, 32'hc2cbdc65},
  {32'hc49cccee, 32'hc3b735dc, 32'hc2d15bac},
  {32'h43590df0, 32'h43e23e83, 32'h438ac1b3},
  {32'hc4faa596, 32'hc28bb652, 32'hc34815bc},
  {32'h435f0000, 32'hc2077326, 32'h43f4c2cb},
  {32'hc39ac21b, 32'hc0bc31e1, 32'h4365e275},
  {32'h4509ffec, 32'h4338c80a, 32'hc39e72dc},
  {32'hc380807b, 32'h43c75889, 32'hc2d8d2d3},
  {32'h4334cbe8, 32'h42bc9be5, 32'h42970445},
  {32'hc3333d27, 32'h438cf92b, 32'hc2f58b3e},
  {32'h44ec4ad0, 32'h405a8d24, 32'h4285c181},
  {32'hc4c6674f, 32'hc278946a, 32'hc3d78c15},
  {32'h44fc897d, 32'h42375e05, 32'h434f1bd8},
  {32'hc4f8cdbe, 32'h42f74321, 32'hc1befa1c},
  {32'h44a3245c, 32'h43cf2e73, 32'hc33ed959},
  {32'hc4c83390, 32'hc3c037f5, 32'h40e99b89},
  {32'h44edaef1, 32'h41f89f84, 32'hc2172bd8},
  {32'hc50569b8, 32'h42a99ff0, 32'hc3cb7433},
  {32'h43aeb6d8, 32'h428795b3, 32'h43102136},
  {32'hc49d6c7c, 32'hc235bf8c, 32'hc24a94ff},
  {32'h44a5d651, 32'h43b37ba6, 32'hc40ca16a},
  {32'hc381c3b0, 32'hc323eda8, 32'hc3586f15},
  {32'h4395e7ba, 32'h42da3d7b, 32'h416223ef},
  {32'h4279ffb8, 32'hc3350c32, 32'hc330607d},
  {32'h450be297, 32'hc34b74cf, 32'h434ca8bc},
  {32'hc401c17a, 32'h433b3517, 32'h43747651},
  {32'h4482083c, 32'h438d6d7f, 32'h40110032},
  {32'hc4a4b318, 32'h42013f4d, 32'hc2069c87},
  {32'h44fd6504, 32'hc2f96d9e, 32'h42e2028e},
  {32'hc42951ba, 32'h432268fa, 32'h420918e0},
  {32'h4500da78, 32'hc1f24179, 32'hc2f89116},
  {32'hc4a1a538, 32'h42b9cc85, 32'hc3d9c8ba},
  {32'h450170af, 32'hc339b2ca, 32'h425d6f94},
  {32'hc4909947, 32'hc29f9084, 32'hc389b8f2},
  {32'h44a9a2de, 32'h4357e354, 32'hc3c654bd},
  {32'hc44b36e2, 32'h42ec5e6f, 32'hc28c612b},
  {32'h43883d80, 32'h43c21775, 32'h4337c1f8},
  {32'hc4bfbdf7, 32'h41a7f0be, 32'hc40db3f1},
  {32'h446920a1, 32'h438946c2, 32'h42609ff6},
  {32'hc4ab5c52, 32'hc310761e, 32'h43c939e8},
  {32'hc4d4b859, 32'hc3e18256, 32'h435188d9},
  {32'h44da87a6, 32'h432734f9, 32'hc188a413},
  {32'hc50ad635, 32'h43e75868, 32'hc32f0ac1},
  {32'h4505fd63, 32'h4396e5d4, 32'h43033716},
  {32'hc4ed5467, 32'h42c256be, 32'hc131e2a4},
  {32'h4452bf4c, 32'hc227cef1, 32'hc3649d8c},
  {32'hc396d084, 32'h430010a7, 32'hc3af1b08},
  {32'h448337fe, 32'h43aae47e, 32'h40fe5f50},
  {32'hc48bcd63, 32'h42a4ec9e, 32'hc11ae7ab},
  {32'h4446768c, 32'h42a9bc94, 32'hc313c277},
  {32'hc4bfeeae, 32'h41aef5f9, 32'hc3fb4a61},
  {32'h450c83ae, 32'hc38c6b22, 32'h422c8ab1},
  {32'hc3fcb58c, 32'hc3d8cc70, 32'h42872e4d},
  {32'h431ffd4c, 32'hc2adeba0, 32'h42f324e6},
  {32'hc40b7656, 32'hc1fecc8e, 32'h4322016a},
  {32'h4366b7d8, 32'hc351eaaa, 32'h42aaea96},
  {32'hc478d067, 32'h43d0d042, 32'hc3a8ac1f},
  {32'h43aa21ba, 32'hc3638632, 32'h43015410},
  {32'hc4c78c7a, 32'h432a43ce, 32'hc3008633},
  {32'h44e6c15b, 32'h43278a4a, 32'h41b78795},
  {32'hc2df03a0, 32'h42fad030, 32'h422dc0d1},
  {32'h4438615e, 32'hc20c2f37, 32'h428c62b9},
  {32'hc5043210, 32'hc3035bac, 32'h41d8923e},
  {32'h4423296a, 32'h423d06d4, 32'h43bf894e},
  {32'hc38b0635, 32'h4246da71, 32'hc33017f1},
  {32'h4505e8aa, 32'h43762e5f, 32'h43462718},
  {32'hc423deac, 32'h4391faeb, 32'hc2d646fc},
  {32'h435d9fe0, 32'hc40d4833, 32'hc3ec9682},
  {32'hc4c54cf6, 32'hc29e0a24, 32'h427f11a6},
  {32'h4511de92, 32'h43c98039, 32'h4282fe2e},
  {32'hc40f11aa, 32'h43176636, 32'hc3686706},
  {32'h43689160, 32'h43396267, 32'h42913b26},
  {32'h42067c00, 32'h43a9a446, 32'h42dd0506},
  {32'h44ec9036, 32'h42adca15, 32'h42dab30d},
  {32'hc4748b64, 32'hc3229e77, 32'hc3bd7d1e},
  {32'h43324820, 32'h43528569, 32'h42cc8ce5},
  {32'hc3f87d38, 32'hc15e1a3c, 32'hc3976703},
  {32'h44a5c0a6, 32'hc223fe0e, 32'hc38a352a},
  {32'hc469addc, 32'h436633e3, 32'h423ea0c2},
  {32'h43dbac6c, 32'hc38e6aa0, 32'h4206c0d1},
  {32'h4357ac02, 32'h42ae5273, 32'hc14093de},
  {32'h4506f7ab, 32'hc3825bb9, 32'hc353fbc4},
  {32'h41bd9c80, 32'hc3b22e04, 32'h43896970},
  {32'h446eea12, 32'h4232f893, 32'h43848e83},
  {32'hc3935588, 32'h43160cb6, 32'h42ef0b7e},
  {32'h4505b0ec, 32'h41e22a28, 32'h4351914f},
  {32'hc4576ffd, 32'h4291a66e, 32'hc11a5069},
  {32'h45158a1f, 32'h43917e64, 32'hc3ce4e01},
  {32'hc4fe3e8e, 32'hc397accf, 32'h410617c0},
  {32'h4486e1af, 32'h41b2634d, 32'h42520c3f},
  {32'hc3871156, 32'hc3178c40, 32'h418744a5},
  {32'h450e1038, 32'h422835dd, 32'h432e6e75},
  {32'hc5056914, 32'hc29ffd62, 32'h432af83c},
  {32'h4384a2d2, 32'hc16488cd, 32'h439e5619},
  {32'hc4d9f739, 32'h434d78a2, 32'hc255de9e},
  {32'h43874109, 32'h41aa24f3, 32'hc31c97ad},
  {32'hc507b9b2, 32'h434fc149, 32'h41b44704},
  {32'h44bd09e5, 32'h43dc8f40, 32'h42b425c6},
  {32'hc48c1455, 32'hc3a5ffbe, 32'hc390e9c3},
  {32'h4515886e, 32'h42a37be1, 32'h42528ab1},
  {32'hc503d975, 32'h43894c50, 32'h42b1b9bd},
  {32'h45033502, 32'h412fcb3d, 32'h427a7ddc},
  {32'hc4a0e1c4, 32'h4167d53b, 32'h41a95fab},
  {32'h450987ad, 32'hc16ae451, 32'h4374b4ae},
  {32'h4380f149, 32'hc325eacd, 32'hc302a1e7},
  {32'h43ea7cb1, 32'h42906584, 32'h439d79f1},
  {32'hc46df9b8, 32'h43c58da1, 32'h42bfa352},
  {32'h449a5abd, 32'hc3060022, 32'hc2d1a4e7},
  {32'hc49a8673, 32'h4295ff3c, 32'hc2ded23d},
  {32'h450e95a2, 32'hc38f3005, 32'hc324777b},
  {32'hc4c9c9bd, 32'h40e79684, 32'h429f986b},
  {32'h44d855c9, 32'hc359961c, 32'hc360b60d},
  {32'hc41323e6, 32'h439c6675, 32'h43752eb8},
  {32'hc20d21e0, 32'h42ef283a, 32'hc22f9674},
  {32'hc501178e, 32'hc2fa3683, 32'h434cfc9d},
  {32'h45122af8, 32'hc34f27c5, 32'h43d5e67c},
  {32'hc46cadef, 32'h42a13f84, 32'h43590ffd},
  {32'h4503a0ae, 32'hc37bdeb1, 32'h4254aa9d},
  {32'hc51f5cfd, 32'h42d0284b, 32'hc295a7cb},
  {32'h449bbb73, 32'hc36d4af3, 32'h4395d1a4},
  {32'h414f4600, 32'hc372604a, 32'hc14fc020},
  {32'h45013fe5, 32'hc35e2eff, 32'hc2a1fd8b},
  {32'hc3935f72, 32'hc3d8fee9, 32'hc3bbdf20},
  {32'h44b9301f, 32'hc3086aff, 32'h4329aeb1},
  {32'hc49cc08a, 32'h43ac0862, 32'h42b2c053},
  {32'h44666320, 32'hc22c1ec6, 32'h4397d468},
  {32'h42101d80, 32'hc1b164f4, 32'h436f225b},
  {32'h44cf5f31, 32'hc1bfbd23, 32'hc336c638},
  {32'hc4aeb2ef, 32'h42f1496e, 32'hc1a9ffd5},
  {32'h44ae95cb, 32'h428411cb, 32'hc3c28ef7},
  {32'hc4da788e, 32'h433f360b, 32'h414b9e0a},
  {32'hc3145c44, 32'h4107836f, 32'h433bb948},
  {32'hc45473a1, 32'h4374bdd8, 32'h41d7b1a1},
  {32'h44cc76a4, 32'h4304ac0c, 32'h43530508},
  {32'hc5097984, 32'hc3e45aa9, 32'hc39b2c57},
  {32'h44326293, 32'hc36f7e03, 32'h42d77cef},
  {32'hc48e1e03, 32'h42945bd9, 32'h433bd935},
  {32'hc0b4ba40, 32'hc1b46e35, 32'hc212182d},
  {32'hc50dd7ca, 32'h43f0456a, 32'hc1c6d08b},
  {32'h44fa94f5, 32'h3fe28054, 32'hc2dad892},
  {32'hc506158b, 32'h42ea18b2, 32'hc2d72a70},
  {32'h44bfa55b, 32'h435399ec, 32'h42d609a3},
  {32'hc4200f8e, 32'hc2eb0f62, 32'h43963247},
  {32'h444f0a97, 32'h42a10134, 32'h42ccd66e},
  {32'hc4d98af0, 32'h430980c4, 32'hc20e3beb},
  {32'h43bb124c, 32'hc398a0ca, 32'hc360b465},
  {32'h42b236cc, 32'h42976979, 32'hc29d9d17},
  {32'h448cef78, 32'h42f777eb, 32'hc3a46e9c},
  {32'hc4f6b95c, 32'h42b1a897, 32'h43021318},
  {32'h44e5d48c, 32'h42495889, 32'hc2f5bba9},
  {32'hc5013770, 32'h41e5f0ea, 32'h434fc510},
  {32'h4468b3ff, 32'h43b2094c, 32'hc31e26b1},
  {32'hc4e60036, 32'h43a010f7, 32'h43e16ae8},
  {32'h432ec922, 32'h43e4e5f7, 32'h4103c766},
  {32'hc347ab94, 32'h4082c1c8, 32'h43a3a921},
  {32'h44e659bd, 32'hc334c52b, 32'hc40d947d},
  {32'hc4ddb4f2, 32'h439bff96, 32'h432bd93f},
  {32'h4505223b, 32'hc384b1ef, 32'h4298feae},
  {32'hc3f0eed4, 32'h4345d56d, 32'h43d2f696},
  {32'h4504661a, 32'hc1c7ba7f, 32'h428ca482},
  {32'hc4bf579a, 32'h41ccdea6, 32'h42561cc4},
  {32'h442c3e40, 32'h41d2730d, 32'h4307a54d},
  {32'hc5072e22, 32'h40e19c4b, 32'h43adc488},
  {32'h44ac2e20, 32'hc1c1b5d0, 32'h41848691},
  {32'hc5044d20, 32'hc3ebc9b9, 32'h4315ea6c},
  {32'h44a5887a, 32'h42c35370, 32'h41a49572},
  {32'hc344b150, 32'hc14328e6, 32'hc2883ba8},
  {32'h44b10e9e, 32'h4367f5b5, 32'h41f2b1ea},
  {32'hc4a3e4c8, 32'h41f3b444, 32'hc2c52f24},
  {32'h44f80e32, 32'hc1ad543c, 32'hc3296767},
  {32'hc4f19086, 32'h4204c8f1, 32'hc292ca45},
  {32'h4484a005, 32'h430511bb, 32'h432534bb},
  {32'hc27e07e8, 32'hc3521d35, 32'hc2ac967a},
  {32'h444dfa7a, 32'hc329ebe7, 32'hc2c64186},
  {32'hc4956b94, 32'hc30e63b9, 32'h42f384bd},
  {32'h45154f05, 32'h4392b6ea, 32'hc3bf44c5},
  {32'hc3a7d5c4, 32'h438100f8, 32'h439e2ab8},
  {32'h44cfe8d2, 32'hc355dcef, 32'hc34ccb5e},
  {32'hc4fa81d6, 32'hc3367f9c, 32'hc2b9a797},
  {32'h448b03b0, 32'hc3f1b8cf, 32'hc2baa52e},
  {32'hc393998c, 32'h430d2037, 32'h41998138},
  {32'h44212ef7, 32'hc364e71e, 32'h43195a9d},
  {32'hc4aa8a35, 32'h41ae131f, 32'hc1c3d2d7},
  {32'h44b3a591, 32'hc38e1c36, 32'h4388fdbf},
  {32'hc41c83e4, 32'h440b386a, 32'hc39cb742},
  {32'h44cbc3b2, 32'hc3adfbf1, 32'hc2d13cd4},
  {32'hc4d3e01c, 32'hc1f2aca3, 32'h43805d8f},
  {32'h432b42a0, 32'hc1ede655, 32'h42effe3c},
  {32'hc3cdd5a0, 32'hc304f67b, 32'h42e969ac},
  {32'h44e7a6e4, 32'h424c8822, 32'hc3213f23},
  {32'hc4dcf397, 32'h4312d767, 32'h43792fd7},
  {32'h44af6cde, 32'h42b22c67, 32'h42e05c78},
  {32'hc406e6ee, 32'h42f56324, 32'hc2415f55},
  {32'h451fcedd, 32'h41e65538, 32'hc3805c5d},
  {32'hc4cd0f30, 32'h431289ec, 32'h41b966ed},
  {32'h4507975c, 32'hc0a313c6, 32'h415f4b99},
  {32'hc513a86d, 32'hc38d5994, 32'h43b223e8},
  {32'h44eb97a0, 32'h439c3092, 32'h431e5cbd},
  {32'hc4afaeb7, 32'h42d6fd88, 32'hc2a85f1e},
  {32'h440b0644, 32'h42651d7c, 32'h43515e0a},
  {32'hc4a48e14, 32'h425a246d, 32'hc351a207},
  {32'hc32b7890, 32'hc314695d, 32'hc3af53a7},
  {32'hc4ac419d, 32'h437c6d77, 32'h432fff8b},
  {32'h4407aa7c, 32'h435ba89f, 32'hc3ace27c},
  {32'hc49c90c3, 32'hc2700097, 32'h43284fb0},
  {32'h4414f4a7, 32'hc3690fe8, 32'h41a026d4},
  {32'hc468d4c4, 32'hc283a549, 32'h4353bb70},
  {32'h4383ada8, 32'h42c200e3, 32'h43a4c121},
  {32'hc438817c, 32'hc406d836, 32'hc30b626e},
  {32'h449ef6aa, 32'h43347995, 32'hc2bd52b8},
  {32'hc522a418, 32'hc3c25459, 32'hc3129c67},
  {32'h448af3a7, 32'hc3df731c, 32'hc1e09380},
  {32'hc4c6497c, 32'h434ebd13, 32'hc285a177},
  {32'h446d808f, 32'h4303a677, 32'hc29f423e},
  {32'hc4d8c482, 32'h41d5dd16, 32'hc2812908},
  {32'h44ae8c71, 32'hc2c5b47f, 32'h417319e2},
  {32'hc4e8b5fa, 32'h42631f84, 32'hc407056b},
  {32'h44af8300, 32'hc374657b, 32'hc32c9948},
  {32'hc1a2b280, 32'hc3e2a6b9, 32'h4419825f},
  {32'h4487544b, 32'hc28da9ae, 32'hc2128c2a},
  {32'hc294e410, 32'h4345ffbc, 32'hc2cee657},
  {32'h4405bcf0, 32'h42a59b79, 32'hc2e62e81},
  {32'hc49e9aca, 32'h42949cf6, 32'h42ba1176},
  {32'h43cb7e70, 32'h43d4fad4, 32'h42836ae9},
  {32'hc4b47d79, 32'h4362978a, 32'hc323983d},
  {32'h43dc3b2b, 32'h421b7f90, 32'h41871144},
  {32'hc50f26d3, 32'hc287e6bc, 32'hc1c0ea3b},
  {32'h42cabd10, 32'h4333a67a, 32'h43602a2b},
  {32'hc3c9ed90, 32'hc390f6a2, 32'hc2495538},
  {32'h432b9f94, 32'hc39b9e6c, 32'hc2b4ab55},
  {32'hc3165924, 32'h42c5a8e0, 32'hc223f659},
  {32'h4500aea0, 32'h43423884, 32'hc385b1fb},
  {32'hc3960f3a, 32'hc2b096ab, 32'hc31dd1cc},
  {32'h43013e18, 32'h4347108f, 32'h430c88b6},
  {32'hc437316a, 32'h4332f943, 32'hc352db3d},
  {32'h44645416, 32'hc3f0ab9a, 32'h43164f2f},
  {32'hc505ee6a, 32'hc39cdb25, 32'h43466646},
  {32'h3fe00000, 32'h40c054f6, 32'h42844f4c},
  {32'hc44c490a, 32'h42250f3e, 32'hc24fb506},
  {32'h44126dba, 32'h41123898, 32'h43c06af7},
  {32'hc373c2a0, 32'h4309f605, 32'h4268c9fd},
  {32'h44c8b013, 32'h43769b2d, 32'h431beee1},
  {32'hc4f83105, 32'h439067a8, 32'h438da8df},
  {32'h42f7eaa0, 32'h42963ae1, 32'h432a1452},
  {32'hc28f5120, 32'h418339ee, 32'h42e23e1d},
  {32'h448c3d4a, 32'hc35b7b06, 32'h4315d5ad},
  {32'hc4a84a5a, 32'hc3a98b6f, 32'h432a421d},
  {32'h44f84e98, 32'h43d51178, 32'h40f353e0},
  {32'hc351442a, 32'hc1863105, 32'h42287cf1},
  {32'h44bede28, 32'hc2699c56, 32'hc2edba30},
  {32'hc5005593, 32'hc385bead, 32'hc25e96d0},
  {32'h45149ddb, 32'h3e34efb6, 32'hc40d84cb},
  {32'hc4d13977, 32'h434b074f, 32'h413f6258},
  {32'h4417f0bc, 32'h43218e3b, 32'hc12184df},
  {32'hc4893d0d, 32'h425a4e0a, 32'h42ca9f66},
  {32'h43efcf78, 32'hc3a8778e, 32'hc22be5e4},
  {32'hc3deecb8, 32'h43075dee, 32'hc2af9b2f},
  {32'h44d0b80a, 32'hc278e102, 32'hc3369735},
  {32'hc4fc6cdc, 32'h42fd80b0, 32'h43d9ae27},
  {32'h448da254, 32'hc2f6d5f7, 32'h427eed18},
  {32'hc4cfe043, 32'hc31f4675, 32'h42eaef0d},
  {32'h445b6046, 32'hc3864055, 32'h41988930},
  {32'hc4dd1f85, 32'h42c69d76, 32'h410d1d1c},
  {32'h441ad29e, 32'hc34b6c3c, 32'hc2ebe7e2},
  {32'hc426d67f, 32'hc2b0ac5a, 32'hc3093351},
  {32'h44c7c7e7, 32'h43eabad6, 32'hc226e2a2},
  {32'hc41aa1a2, 32'h44033098, 32'hc333103c},
  {32'h447a646e, 32'h41aa95df, 32'hc36ff1e6},
  {32'hc4e5a1a9, 32'hc29f63e4, 32'hc251fe7b},
  {32'h448c2485, 32'hc3dcae18, 32'hc304b4af},
  {32'hc4dcb36c, 32'hc2b623af, 32'h43c598fb},
  {32'h44d808b9, 32'hc348fabd, 32'h429f4680},
  {32'hc40014a4, 32'h42d6080f, 32'hc39da34c},
  {32'h4429d140, 32'hc4118bb0, 32'h42bcfae1},
  {32'hc4229120, 32'hc32175d0, 32'h42cd8df7},
  {32'h425985f0, 32'hc2865025, 32'h4407457e},
  {32'hc3f99d08, 32'hc4219369, 32'h4249bc3b},
  {32'h44d0abf4, 32'hc2fd4daf, 32'hc3a77b73},
  {32'h43262790, 32'h42f03c44, 32'hc32801e2},
  {32'h448f8bc1, 32'h41f65919, 32'hc1be4a59},
  {32'hc44542e2, 32'hc34c913c, 32'hc3143a4f},
  {32'h44990315, 32'h4401add8, 32'hc3e08c04},
  {32'hc4f3edec, 32'h42a68d57, 32'h424f5e29},
  {32'h43566978, 32'hc293dc1b, 32'hc319b1bc},
  {32'hc4b395f2, 32'hc2e997bc, 32'h43197a67},
  {32'h450a992f, 32'hc2f19512, 32'h43c397c5},
  {32'hc4cf2e5f, 32'h43651bf6, 32'hc261a9f6},
  {32'h44c1c508, 32'hc3bac60f, 32'h42fc065f},
  {32'hc4655cee, 32'h4302098c, 32'hc34175f0},
  {32'h44927b64, 32'hc39f1111, 32'hc2dc4835},
  {32'hc4c03963, 32'h43af400f, 32'hc3b18d4d},
  {32'h4431a128, 32'hc3f542f1, 32'hc308d4c9},
  {32'hc51a51ab, 32'hc34ef80b, 32'h434e87c5},
  {32'h439d7f90, 32'hc39204df, 32'hc3303639},
  {32'hc47cfc54, 32'hc3af24c9, 32'hc3bdb407},
  {32'h4502df7e, 32'hc30bb435, 32'h42da7b65},
  {32'hc40adee4, 32'h429ea61c, 32'hc2810e60},
  {32'h45104c14, 32'h435171ba, 32'hc2d5c1d3},
  {32'hc4b5c5e6, 32'hc2ddf4ec, 32'hc3d3e3ea},
  {32'h44bd79f4, 32'h4414c3b8, 32'h438a9f7b},
  {32'hc41dd148, 32'h436f419e, 32'h42b99bf4},
  {32'h449deaf6, 32'hc339ca2f, 32'h42e9fabe},
  {32'hc4b1de86, 32'h43b9bc9a, 32'h42d5c450},
  {32'h44148eac, 32'hc21199e9, 32'hc30a406b},
  {32'hc4bd3da6, 32'hc36de868, 32'h4374263f},
  {32'h43a450d0, 32'h42b1bd8a, 32'h42d847c3},
  {32'hc2fd556c, 32'h40ab3956, 32'hc2b9b56b},
  {32'h438f1124, 32'hc3236931, 32'hc1821220},
  {32'hc47a8b9b, 32'h430c23f3, 32'hc249f2da},
  {32'h4476f06b, 32'hc32f081a, 32'h43fde2ac},
  {32'hc409afd4, 32'hc27a3bea, 32'hc30427fb},
  {32'h43ffbfc1, 32'hc3bfe2df, 32'h4217adba},
  {32'hc413c09b, 32'hc38511c8, 32'hc39cb230},
  {32'h44c5a4f4, 32'hc2fd63a4, 32'h41f0c0e3},
  {32'hc4ba2d4a, 32'hc3a8962e, 32'h439ba251},
  {32'h4404ea1c, 32'hc366ba58, 32'hc31ee20f},
  {32'hc3f1abae, 32'h43cb6473, 32'hc10cdb9c},
  {32'h441ffe66, 32'h42dc1038, 32'h41f9d94b},
  {32'hc43ccb1a, 32'hc28676b9, 32'hc3971231},
  {32'h430e3b28, 32'h41c3a587, 32'hc10a7c47},
  {32'hc4fbe446, 32'hc2d06716, 32'h43577f70},
  {32'h44c38814, 32'h436c0048, 32'hc3896650},
  {32'hc46a258b, 32'hc0deec46, 32'h42b9a850},
  {32'h44ee0bd3, 32'hc0921642, 32'h43864d88},
  {32'hc4231daa, 32'hc263df83, 32'h43598243},
  {32'h445802ee, 32'h420f6f15, 32'h4183db36},
  {32'hc416d67d, 32'h42972dfb, 32'hc36b5a88},
  {32'h44857eda, 32'h42081f0d, 32'hc2926e19},
  {32'hc4ba204f, 32'h437966f0, 32'h43f48020},
  {32'h43eed921, 32'h441030ed, 32'h439b6d9d},
  {32'hc2329180, 32'hc3a95737, 32'hc2eca419},
  {32'h444bdec9, 32'h431188a5, 32'hc2d5a506},
  {32'hc50a54df, 32'hc2f2d961, 32'h432dfead},
  {32'h44ea7849, 32'h416d5656, 32'hc234a38b},
  {32'hc4fe8c4c, 32'h4290baf2, 32'hc24e82be},
  {32'h44ef726c, 32'hc2fbd393, 32'hc2b5d791},
  {32'hc5099c37, 32'hc38f9a5f, 32'h42546c33},
  {32'h4500b129, 32'hc2d59346, 32'hc17b0216},
  {32'hc3cbb1be, 32'h43ed61a2, 32'h42c1ee0c},
  {32'h44e12d13, 32'hc207ebc6, 32'hc28763f6},
  {32'hc498e704, 32'h43b84cc4, 32'hc20dd075},
  {32'h44a34443, 32'h4323ea2c, 32'h427fe36b},
  {32'hc4983951, 32'h41e21be6, 32'h4323b5df},
  {32'h44e71ffb, 32'hc19d6738, 32'hc374e2c8},
  {32'hc3fd5aa4, 32'hc39e6beb, 32'h432ad4ec},
  {32'h44dc8734, 32'hc39d1084, 32'hc396e4b7},
  {32'hc4a258cb, 32'hc128d832, 32'hc40f579e},
  {32'h43f9bb90, 32'h42466211, 32'hc32f1ad5},
  {32'h43da5155, 32'h41bf8c87, 32'h436e77e9},
  {32'h44a4989e, 32'hc3b1b72c, 32'h4353750b},
  {32'hc4e9cbb0, 32'hc303b33c, 32'h4343e4a8},
  {32'h449d5410, 32'h433a0208, 32'h438aa88e},
  {32'hc3fda334, 32'hc37ffa5e, 32'h42b1ad14},
  {32'h45054430, 32'hc3a107ae, 32'h43c86e9c},
  {32'hc2c9e6a0, 32'h43b1d62d, 32'hc3cfbeca},
  {32'h451370fb, 32'h42f8d33d, 32'h422e15f1},
  {32'hc4ba6e98, 32'h4289ae42, 32'hc3e063c9},
  {32'h44919bbc, 32'hc3066d00, 32'hc2ae0ea4},
  {32'hc4a24c96, 32'hc39597c1, 32'hc38286fc},
  {32'h4483b441, 32'hc32a6d18, 32'h423f6a84},
  {32'hc46dfa83, 32'hc2ee138b, 32'hc2f7f5ec},
  {32'h44e166b7, 32'hc282824b, 32'hc2bf5c16},
  {32'hc424f690, 32'hc33b4f3e, 32'h42b33e48},
  {32'h44291340, 32'h4308094a, 32'h4314102c},
  {32'hc40f98fc, 32'hc392f1eb, 32'hc37d97ee},
  {32'h431f0afc, 32'hc12fc75f, 32'h4253e4ca},
  {32'hc3c70e98, 32'h4373fe11, 32'hc289f790},
  {32'h43bd0fb0, 32'h436e766e, 32'hc298aa78},
  {32'hc4bbcd10, 32'h411ae27c, 32'hc3af06ac},
  {32'h44cbf801, 32'h4369561f, 32'h4225f910},
  {32'hc4ba6d7f, 32'hc154e6e5, 32'h43496864},
  {32'h4410a2f0, 32'h439db5ed, 32'h43322ba6},
  {32'hc51088fa, 32'h42fb0fdd, 32'hc2d87052},
  {32'hc21d0c20, 32'h43868b01, 32'hc3d36de6},
  {32'hc47f5e87, 32'h43ace0a9, 32'hc3bbaa97},
  {32'h44602192, 32'hc3520260, 32'hc300550f},
  {32'hc3a1733f, 32'h431daa64, 32'hc3469ce1},
  {32'h4471791b, 32'h4313d1f7, 32'hc35a80c3},
  {32'hc491fe0d, 32'h430c0899, 32'h435d904f},
  {32'h43d1544e, 32'h41457fba, 32'h4316c65c},
  {32'hc4b80c74, 32'hc31eeeef, 32'hc286f29d},
  {32'h45082da7, 32'hc2cda205, 32'hc1dc1f52},
  {32'hc5107149, 32'h42b12eee, 32'h41d0f282},
  {32'h448dea2e, 32'h436e15e4, 32'h421acf3c},
  {32'hc4db73bc, 32'hc2c92743, 32'hc30974ea},
  {32'h44c7f814, 32'hc30a9cd9, 32'h43c8d416},
  {32'hc4d3b512, 32'hc27bf40e, 32'hc1937c5a},
  {32'h43d6c412, 32'h42fbd16d, 32'hc3a5d7e2},
  {32'hc47631f2, 32'hc3528e13, 32'hc292d025},
  {32'h43cfa18e, 32'hc1b8628c, 32'h42afe3f1},
  {32'hc480b420, 32'hc3a05a82, 32'h42f52506},
  {32'h44a38308, 32'hc2340ef2, 32'hc38bf2ee},
  {32'hc4343ee4, 32'hc2ae6804, 32'h42a44804},
  {32'h452679cf, 32'hc1cd2f3d, 32'hc38bfa23},
  {32'hc3f00ecc, 32'h4402cda7, 32'hc2109d14},
  {32'h4309f040, 32'hc38b7550, 32'h439915d0},
  {32'h43a122e8, 32'h43cfbd0f, 32'hc2c758b0},
  {32'h42eb84f0, 32'hc3cad864, 32'hc28dfb81},
  {32'h42fa17ca, 32'hc228e809, 32'h43a82140},
  {32'h44af53dd, 32'hc3e353c9, 32'h4311cbce},
  {32'hc40de832, 32'h42207531, 32'h43ebd74a},
  {32'h44869ee5, 32'hc3eccf33, 32'hc3305810},
  {32'hc4d1041d, 32'hc329832f, 32'h425c954c},
  {32'h447151a8, 32'hc2d301c5, 32'hc3472336},
  {32'hc524b3f9, 32'h4384202b, 32'hc4034e2d},
  {32'h45180d19, 32'hc178d685, 32'hc280f286},
  {32'hc50db312, 32'hc2b1bea5, 32'hc360faf8},
  {32'h4505b27d, 32'h42163bab, 32'hc1403c9e},
  {32'hc514c4fe, 32'hc31d253d, 32'hc33e6dfb},
  {32'h44a05fe6, 32'hc35eabd9, 32'hc336e0ac},
  {32'hc4831960, 32'h418d0271, 32'h434e1845},
  {32'h44963540, 32'hc2969151, 32'hc3a4e2be},
  {32'hc4b5156e, 32'hc34e3a84, 32'h439389ad},
  {32'h44b97d05, 32'hc36483fc, 32'hc1133208},
  {32'hc40aa044, 32'h437e6a7c, 32'hc3dfe634},
  {32'h44aa68ab, 32'h421a4d52, 32'hc3236a7e},
  {32'hc4790601, 32'h438aa4b4, 32'hc33cc2b8},
  {32'h44a18aff, 32'hc3d7e3d0, 32'hc31e705e},
  {32'hc31692c0, 32'hc259367d, 32'h433647a5},
  {32'h42ea6cc6, 32'h41acda2d, 32'hc2e8e838},
  {32'hc498fff8, 32'h429b87ee, 32'hc31f6100},
  {32'h45042f7f, 32'h42ec96df, 32'hc39574d8},
  {32'hc4e81452, 32'h4252688a, 32'h423be418},
  {32'h44a4b7b0, 32'hc29ed6bf, 32'h43857219},
  {32'hc4614098, 32'h4327c281, 32'h425586e0},
  {32'h44c56936, 32'h4012fe32, 32'hc34f1054},
  {32'hc508b43b, 32'hc31b6ba7, 32'h4324283f},
  {32'h451261a2, 32'hc3897e24, 32'h43359823},
  {32'h4213cf00, 32'hc2c022cb, 32'h43a7044e},
  {32'h4427ea3b, 32'h43321b0e, 32'hc3af7c13},
  {32'hc482d6ae, 32'hc194f03d, 32'h420a0636},
  {32'h4383b357, 32'hc35cc4ce, 32'hc25d35bb},
  {32'hc480046a, 32'hc2dfd53e, 32'hc2e7a1f2},
  {32'h437e6d20, 32'hc323279e, 32'h415bdba4},
  {32'hc4cd1090, 32'hc1e73aa0, 32'h40fef69c},
  {32'h4495a018, 32'h4210bb31, 32'hc31966cf},
  {32'hc501404c, 32'hc138ef68, 32'h3fd42379},
  {32'h4526eeb0, 32'hc182afc4, 32'hc35f382c},
  {32'hc4eca307, 32'hc19b2c5e, 32'hc33438ee},
  {32'h45141c4d, 32'h424a8c6c, 32'hc2d23105},
  {32'hc44b3652, 32'h439793e1, 32'h43815c46},
  {32'h44a23f7c, 32'hc3f1f18e, 32'hc3df02f7},
  {32'hc42e6948, 32'hc2c69827, 32'h43ba31cf},
  {32'h4479a7c8, 32'hc31f80b2, 32'hc2d04a17},
  {32'hc498d553, 32'h43c58899, 32'hc30da6f2},
  {32'h44fb9bfc, 32'h417c851c, 32'h4289bcdf},
  {32'hc478de41, 32'h420216a5, 32'hc34cabea},
  {32'h4485e3f4, 32'h43254d1b, 32'hc33b40ea},
  {32'hc498761c, 32'h42dc1810, 32'hc2061848},
  {32'h4451dfee, 32'hc20c5432, 32'hc35e19b6},
  {32'hc4b7b610, 32'hc2c0763b, 32'h4404b240},
  {32'h446bf7bb, 32'hc40385b6, 32'hc38f5def},
  {32'hc49a6954, 32'h42c21625, 32'h41d521d5},
  {32'h44235f60, 32'h42aeb8dc, 32'hc327eefb},
  {32'hc3f51998, 32'hc31da2d9, 32'h42ec7902},
  {32'h43de8c4a, 32'h4312ac40, 32'hc1812fb9},
  {32'hc3ec8780, 32'hc32885e3, 32'hc342029b},
  {32'h445dd064, 32'hc265f956, 32'h42939697},
  {32'hc3fdb85f, 32'h431880ea, 32'h42856cd3},
  {32'h4479bd42, 32'hc34e1b4e, 32'hc39b22e0},
  {32'hc33e5bec, 32'hc29b1ab0, 32'hc2bb53ca},
  {32'h442e33a4, 32'h43a5690e, 32'h430febc0},
  {32'hc4edc87d, 32'hbe9d4a8c, 32'hc23166a3},
  {32'h44d067d5, 32'hc334a93c, 32'hc3c39dd0},
  {32'hc319826b, 32'h431f21f6, 32'hc2cfaf1d},
  {32'h447d3d28, 32'h43c2d19e, 32'h42ddd744},
  {32'hc50ad413, 32'h42c9019c, 32'hbfa8f24d},
  {32'h44d52111, 32'hc22e349e, 32'hc34da1b1},
  {32'hc4091c36, 32'h4329664d, 32'h43857a4c},
  {32'h450ac460, 32'h425a1194, 32'hc30e7774},
  {32'h42f9a170, 32'h43c3ed1e, 32'hc212d01c},
  {32'h43783ff0, 32'hc32703d8, 32'hc223bc0a},
  {32'h44e010b4, 32'h43acfea7, 32'hc3bef2f5},
  {32'hc39bc382, 32'h422d9eb9, 32'h4111891a},
  {32'h44159840, 32'h43298706, 32'h4234bc09},
  {32'hc5349474, 32'h438e3b7a, 32'hc29ef983},
  {32'h43e24ca6, 32'hc2bb66d7, 32'hc373b79c},
  {32'hc475a8e0, 32'h4308d087, 32'h41f53b9a},
  {32'h44bfdb2a, 32'hc3a52c22, 32'hc30b0a61},
  {32'hc504fd9e, 32'hc2b8a4af, 32'h428cdfc2},
  {32'h44d5136f, 32'hc2b45b97, 32'hc2da0509},
  {32'hc3734e68, 32'hc389db23, 32'hc2f62ddf},
  {32'h44b3a397, 32'hc3792416, 32'hc380db48},
  {32'hc2e13146, 32'hc31216b8, 32'h43c18324},
  {32'h44ab977d, 32'h430b4566, 32'hc377b356},
  {32'hc444f9c0, 32'hc304c68a, 32'hc34b8877},
  {32'h45107b9d, 32'h438fce5a, 32'h4146f76c},
  {32'hc4e7f9dc, 32'hc305486f, 32'hc32a1965},
  {32'h41b2e3a0, 32'hc30c75b7, 32'h43a4c963},
  {32'hc4cef813, 32'h434b7fb0, 32'h43289984},
  {32'h44f8f4b7, 32'hc312e790, 32'hc1248b0a},
  {32'hc4ee5acd, 32'h428167f8, 32'h435b87a7},
  {32'h41a20900, 32'h4354117c, 32'hc20535b6},
  {32'hc4bfe5e0, 32'h41ebfa44, 32'h438caf30},
  {32'h44ca37bd, 32'h43244016, 32'hc3236812},
  {32'hc5116307, 32'h411b7148, 32'h42dbc858},
  {32'h44f73a40, 32'h4323e049, 32'hc149d348},
  {32'hc449f530, 32'h4365ff07, 32'h438c0c73},
  {32'h434bc408, 32'h42628b6b, 32'h426ae680},
  {32'hc4bb86e8, 32'hc2830140, 32'hc38acafd},
  {32'h447d8173, 32'h4288288a, 32'hc3bb4a27},
  {32'hc4a9c3d3, 32'hc3581bb4, 32'hc352f817},
  {32'h4405338a, 32'hc2f08207, 32'h43356732},
  {32'hc4fa574f, 32'hc3af63e7, 32'hc3f6898c},
  {32'h44c3e4b8, 32'h42abd15b, 32'hc3a4e81b},
  {32'hc2808900, 32'hc2c46fac, 32'hc224bdcd},
  {32'h44eb352e, 32'h428746cc, 32'hc3a83f26},
  {32'hc4a0c06a, 32'hc19e86d3, 32'h43567089},
  {32'h4498bea1, 32'hc1ed99a0, 32'hc32291eb},
  {32'hc5030367, 32'h441d93de, 32'hc3871639},
  {32'h4507f236, 32'hc42a5cb9, 32'h4241bdaf},
  {32'hc37bbcc0, 32'hc2fee83b, 32'hc283fc3c},
  {32'h450eee80, 32'h434ba007, 32'h42bc76b8},
  {32'hc40841ce, 32'h4287930a, 32'hc372e556},
  {32'h44ce5560, 32'h4310d0d1, 32'h4371b0a8},
  {32'hc3003606, 32'h42326ff2, 32'h438b8b98},
  {32'h44c4b443, 32'hc34c337d, 32'h42bdb8cd},
  {32'hc4ddcd83, 32'h43576f15, 32'h433c2dd1},
  {32'h45100f65, 32'h4460c971, 32'hc39e6a99},
  {32'hc4774432, 32'h432922ba, 32'h42d97401},
  {32'h43daee4d, 32'h432274b9, 32'h430f95ac},
  {32'hc46aab0a, 32'h4396eeb9, 32'h4386a50f},
  {32'h43f1af86, 32'hc328aa0f, 32'h43520262},
  {32'hc4333a21, 32'h438c0538, 32'h4303326d},
  {32'h44a7896d, 32'h426c9c3e, 32'hc3d01729},
  {32'hc3afc54c, 32'hc28ee5e4, 32'hc26a0119},
  {32'h450766d1, 32'hc2bf084f, 32'hc2986ac9},
  {32'hc44106f2, 32'hc22e8225, 32'hc2b25eca},
  {32'h450a441e, 32'hc239345c, 32'h42f20b3f},
  {32'hc405054c, 32'h432c879c, 32'hc339028a},
  {32'h44ac3835, 32'hc33681f2, 32'h42ef8dc2},
  {32'hc39cf980, 32'h425ebc23, 32'hc4108730},
  {32'h44b455e1, 32'hc4067ff2, 32'hc3be0e07},
  {32'hc243b340, 32'hc3563112, 32'hc354bf19},
  {32'h43e11dbc, 32'h42cd046a, 32'hc1cf37a0},
  {32'hc43c82d2, 32'hc30cc37d, 32'h4340be83},
  {32'h445b2dba, 32'h438d2df3, 32'hc3a99558},
  {32'hc4ac7ee3, 32'h4372ac04, 32'h42c46d0a},
  {32'h45130dbe, 32'h434f5ff7, 32'hc3c16ce1},
  {32'hc492e486, 32'h42c271eb, 32'h434807fb},
  {32'h44edc5e8, 32'h420fc3c0, 32'hc38a824c},
  {32'hc4600c72, 32'hc334574b, 32'h4250301d},
  {32'h4516995d, 32'hc2c0643f, 32'h42776df0},
  {32'hc49f5e83, 32'hc30dcd7a, 32'hc28e3238},
  {32'h44c8c7fc, 32'hc33c5dbd, 32'hc175203e},
  {32'hc48ea755, 32'h43477f77, 32'hc37c9860},
  {32'h45183051, 32'h43b9542e, 32'h43591ddc},
  {32'hc3ef7465, 32'h4377897c, 32'hc341d01d},
  {32'h4502a5b3, 32'hc2893bfa, 32'hc37dd0a5},
  {32'hc505a84d, 32'h435d8712, 32'hc032d880},
  {32'h44e63c29, 32'hc4090d6b, 32'h440bb62e},
  {32'hc4dc6ecc, 32'hc232559d, 32'hc323bf83},
  {32'h44cc2fb9, 32'hc317c440, 32'h429ad071},
  {32'hc33fc43a, 32'h437a2988, 32'hc30b8361},
  {32'h4501e600, 32'h41a221d6, 32'h4312749e},
  {32'hc3eee58e, 32'h436e5167, 32'hc3bf5d16},
  {32'h4448b5d0, 32'h42e0e32f, 32'hc2226921},
  {32'hc42e460b, 32'hc363c605, 32'hc2fd2d62},
  {32'h43a2195c, 32'h43039449, 32'hc35c807f},
  {32'hc3932578, 32'hc2b2fe82, 32'hc3b19ea3},
  {32'h44ccd972, 32'hc38da91a, 32'h403412e1},
  {32'hc3b6338e, 32'hc2579cdc, 32'hc25e57e8},
  {32'hc0f0a200, 32'hc3b8c084, 32'hc3284bf8},
  {32'hc20518c0, 32'hc38517a8, 32'hc35da862},
  {32'h44e42e12, 32'h41c5b520, 32'hc29c57a9},
  {32'hc5067fdd, 32'h4363a42f, 32'hc33e9547},
  {32'h443f1e56, 32'hc296337c, 32'hc0b2eec9},
  {32'hc3a7d1ec, 32'h4300a1d9, 32'h438ec899},
  {32'h450a974a, 32'hc2702ad6, 32'hc27ee822},
  {32'hc3d017f0, 32'hc251459c, 32'h428406d1},
  {32'h4413a410, 32'h42a080fd, 32'hc36d672a},
  {32'hc3decbb8, 32'h42df0991, 32'hc36ca355},
  {32'h449fe6fb, 32'h42052db5, 32'h421d1b5f},
  {32'hc4e5d452, 32'hc38a8390, 32'hc2ad0eb5},
  {32'h43a9c3b8, 32'h44020e8a, 32'hc2f835f9},
  {32'hc4bf6b97, 32'h42c0ade2, 32'h431cb75a},
  {32'h44c67c0f, 32'hc2b69175, 32'h41c36291},
  {32'hc45abaa4, 32'hc385114b, 32'h42c6fca7},
  {32'h45020272, 32'h4346a56d, 32'hc38a9593},
  {32'hc4de1585, 32'hc37df5ac, 32'hc375fc3d},
  {32'h441fb68b, 32'hc3a99f7f, 32'hc2cdffd8},
  {32'hc44402cc, 32'h431f20ed, 32'hc3485f4d},
  {32'h43e93250, 32'hc30dc293, 32'h4286970d},
  {32'hc4e07a02, 32'hc3330153, 32'h434a4c29},
  {32'h443dc578, 32'hc3169e52, 32'h43148d75},
  {32'hc4997174, 32'h4333a28a, 32'h42cb0626},
  {32'h4505d4c3, 32'hc286b9e2, 32'h428068c3},
  {32'hc50554d8, 32'h43594f0f, 32'hc2593162},
  {32'h44a92e89, 32'hc364392b, 32'hc2700dae},
  {32'hc49a058a, 32'h431cefb6, 32'h43364484},
  {32'h4422bbaa, 32'hc38cdc70, 32'h4355d804},
  {32'hc50a407a, 32'h423a5109, 32'hc2b7e272},
  {32'h44e870aa, 32'hc3291e59, 32'h42badc2a},
  {32'hc483bae8, 32'h42a89a4b, 32'h43eda8c1},
  {32'h44f66759, 32'h43ce14d0, 32'h4376d7e9},
  {32'hc4127001, 32'hc26721be, 32'h4398bd1c},
  {32'h43cecac9, 32'h439a8478, 32'hc2cd807c},
  {32'hc5084882, 32'h42e3ebe1, 32'h4311b884},
  {32'h445f44c2, 32'h432f3453, 32'hc38e0530},
  {32'hc481b4fa, 32'h4319c322, 32'h42147bff},
  {32'h44ed92a6, 32'h434a24fa, 32'hc1d7cdc9},
  {32'hc4ffaa95, 32'h438a18b0, 32'h429b024a},
  {32'h43dcc708, 32'hc32c7152, 32'hc327be9c},
  {32'hc38ddc5a, 32'hc3a2bab4, 32'hc30d3e84},
  {32'h43bfd17f, 32'h421ff347, 32'hc27b629c},
  {32'hc3c7e776, 32'hc2e5a9e4, 32'h41a90008},
  {32'h451672c0, 32'h432a6c70, 32'h42827a93},
  {32'hc3d2d81c, 32'hc390b17a, 32'hc3ba844d},
  {32'h44e3803e, 32'h428061d3, 32'hc3255533},
  {32'hc512bef0, 32'hc3ebb43e, 32'h4328836b},
  {32'h442c0540, 32'h4323a565, 32'hc359dcfe},
  {32'hc4adc119, 32'h4334a7b7, 32'h439a2e1b},
  {32'h45083395, 32'h41bf7579, 32'hc2d8e744},
  {32'h427d8720, 32'h42870c04, 32'h426d3a92},
  {32'h45054953, 32'hc144817a, 32'h43c63cea},
  {32'hc4196150, 32'hc2f205ad, 32'hc2af1f43},
  {32'h44df6fe7, 32'h42347331, 32'hc2bc190b},
  {32'hc4daef9c, 32'h42185aff, 32'hc3d1c1ca},
  {32'h432fb060, 32'hc332b9f4, 32'hc32e3155},
  {32'hc4ea7f62, 32'h415b92f4, 32'h42280462},
  {32'h44c6ac9e, 32'hc2c5da29, 32'h41867ee7},
  {32'hc4c2b700, 32'hc2f8147d, 32'hc302f5ba},
  {32'h44e9a3c7, 32'h41e58973, 32'hc3bc1ace},
  {32'hc3185292, 32'hc39d2437, 32'h42e117ce},
  {32'h450d25ba, 32'h43a63437, 32'hc3d41178},
  {32'hc3936634, 32'h43a2e33a, 32'hc369193e},
  {32'h44c250f8, 32'h431315f2, 32'hc253f697},
  {32'hc3746310, 32'hc32b898e, 32'h4239509e},
  {32'h44cf0916, 32'hc3d0b002, 32'hc3dc877d},
  {32'hc48f7c64, 32'h438ee3e5, 32'hc2b1191a},
  {32'h440142b8, 32'hc31b171a, 32'hc307f372},
  {32'hc3fde20a, 32'h4415313c, 32'hc2a6558d},
  {32'h44fd14d8, 32'h4105fff4, 32'hbf26f74a},
  {32'hc490f078, 32'h43254c29, 32'hc2ff5eca},
  {32'h44638004, 32'h42f3e7e4, 32'h43108ba3},
  {32'hc4ada228, 32'h42098d07, 32'hc367d6f4},
  {32'h450c6055, 32'h432410e9, 32'h428bcbcb},
  {32'hc2958bd0, 32'h43a448df, 32'h423c2dfc},
  {32'h44ffeb48, 32'h435e2c94, 32'h432ae450},
  {32'hc51dd0fb, 32'h4387b1cd, 32'h4355d6f9},
  {32'h44302a7f, 32'h434ab157, 32'h43c41a9f},
  {32'hc4d336e6, 32'h42f7fe98, 32'h432084d1},
  {32'h448e26bc, 32'hc2677616, 32'h409612c0},
  {32'hc43d6534, 32'hc3835bea, 32'h42e4ca7b},
  {32'h45046efc, 32'hc2ab472b, 32'hc24ddf91},
  {32'hc35746c4, 32'hc3677c05, 32'hc38addab},
  {32'h43acfcc0, 32'hc380b14e, 32'h40ab0338},
  {32'hc474171c, 32'h42905b99, 32'hc104748e},
  {32'h44012816, 32'hc1cf7904, 32'hc25dbdc1},
  {32'hc31c3518, 32'hc3153ddc, 32'hc3303af6},
  {32'h4500c1eb, 32'h4379384d, 32'hc3a6e815},
  {32'hc4b0b359, 32'hc3b96ba7, 32'hc1dd0bcf},
  {32'h4500ac13, 32'h43ede7d8, 32'hc3386979},
  {32'hc4bcd899, 32'hc22a3b8d, 32'hc2a769b3},
  {32'h443e9f3d, 32'hc3bed329, 32'h4321db93},
  {32'hc488f4f1, 32'hc3336552, 32'hc3efda5c},
  {32'h441f6c5c, 32'hc29e89f0, 32'hc27e37fc},
  {32'hc457924f, 32'h41cba236, 32'h428f1c34},
  {32'h44b60881, 32'h439d2e57, 32'hc31d9979},
  {32'hc490f255, 32'hc39475b6, 32'h41437297},
  {32'h4474ecd0, 32'h4289de08, 32'h42ebf8e7},
  {32'hc4ed201d, 32'hc2f51d52, 32'hc30cd38a},
  {32'h44fa5543, 32'h42da459b, 32'h4310ced5},
  {32'hc4d2a436, 32'hc2ab0cb4, 32'hc3773693},
  {32'h44ee3faf, 32'hc381df3d, 32'hc3139a90},
  {32'hc487d1b4, 32'hc29ae892, 32'h43840c33},
  {32'h44844ef7, 32'h4191c112, 32'hc31836bc},
  {32'hc4c4c7e9, 32'h4171e46b, 32'h438dc86e},
  {32'h4469583f, 32'hc108498d, 32'hc1332986},
  {32'hc4e2c0fd, 32'h431205b8, 32'h420b2648},
  {32'hc0f0e760, 32'h426f6d02, 32'h434abaf4},
  {32'hc4c05be3, 32'hc3bb4e09, 32'hc2be0bdd},
  {32'h44a461d3, 32'h43821fd2, 32'h423c8d5c},
  {32'hc426ef7e, 32'hc3211994, 32'hc37b9843},
  {32'h449d0e40, 32'h435cb995, 32'hc3621d9c},
  {32'hc40cf992, 32'h43f0c9be, 32'hc39f7c81},
  {32'h44aebef0, 32'hc2b07621, 32'h418de138},
  {32'hc4c75efa, 32'h4239678e, 32'hc3155713},
  {32'h41799980, 32'h42d6760a, 32'h438603c8},
  {32'hc4b92210, 32'hc28dcdca, 32'hc3cf97c9},
  {32'h43877ba0, 32'hc30d6c07, 32'h42e127a6},
  {32'hc507ee0a, 32'h41494312, 32'h42454946},
  {32'h45142170, 32'h425803a2, 32'hc32ac365},
  {32'hc4b181ad, 32'h42f9e2cd, 32'hc3eb9243},
  {32'h43a4009f, 32'hc32c7a6a, 32'hc33e9584},
  {32'hc3c970ae, 32'hc325b456, 32'h437b575e},
  {32'h44ed0fa2, 32'hc31c5ad1, 32'hc00ce9de},
  {32'hc4622eb6, 32'hc1317386, 32'h42701e87},
  {32'h44cdd558, 32'h43b90a26, 32'h4216b632},
  {32'hc33eed6e, 32'h4391817a, 32'h42845ad5},
  {32'h44da5420, 32'hc392ffe3, 32'h40be30d5},
  {32'hc4246eac, 32'hc3a5eb92, 32'hc2e1b24e},
  {32'h44608b5a, 32'hc004bd60, 32'hc1882bba},
  {32'hc521ace2, 32'h43115b36, 32'hc2e9a202},
  {32'h44886aa2, 32'h434c0276, 32'hc3001bf4},
  {32'hc4c5c781, 32'hc3aeca31, 32'hc31f7fe6},
  {32'h43a4ccb0, 32'hc3503a2c, 32'hc39a80be},
  {32'hc4b4d05b, 32'h42c525bc, 32'h41efc1d4},
  {32'h43a1882a, 32'h430c8cb7, 32'hc33afcde},
  {32'hc4deab5e, 32'h42f3280a, 32'hc24871a3},
  {32'h450d4505, 32'hc2153552, 32'hc2b90dff},
  {32'hc4eb4b70, 32'h43d7f5cd, 32'hc3418b2c},
  {32'h44cfafdc, 32'hc354430a, 32'hc297bfb6},
  {32'hc0cb2cc0, 32'h4392117e, 32'hc30acbc2},
  {32'h446fd818, 32'h4131596f, 32'hc33746e1},
  {32'hc47e5a20, 32'hc30951bd, 32'hc3973847},
  {32'h450ce1e7, 32'hc328548a, 32'hc3637e0c},
  {32'hc45669e2, 32'h43463eae, 32'hc3130334},
  {32'h43e6610a, 32'hc3e28e59, 32'h4352aa63},
  {32'hc4ea7d86, 32'hc3353eb3, 32'h43484aeb},
  {32'h449ef19c, 32'hc3889fb4, 32'h430de155},
  {32'hc459eab0, 32'hc2ce8838, 32'h42bde3c5},
  {32'h44900b82, 32'h438c3de6, 32'h42bd9fed},
  {32'hc37849f0, 32'h4333efd6, 32'hc210e7cc},
  {32'h4443731c, 32'hc240aa8b, 32'hbfefc908},
  {32'h4203bb80, 32'h439d1851, 32'hc437e17d},
  {32'h4503daec, 32'hc1ee677e, 32'h42124fc4},
  {32'h4218a2f0, 32'hc37308ef, 32'h4318ef7d},
  {32'h44862d7c, 32'h42308eac, 32'hc3985de0},
  {32'hc40b02a8, 32'hc36cf3f0, 32'h434a9c42},
  {32'h440113cd, 32'h4382006e, 32'hc28f663e},
  {32'hc4b394b0, 32'h428cb7ba, 32'hc2fb9fa6},
  {32'h4402822c, 32'hc3185f3d, 32'h42c8aa3d},
  {32'hc3e1d768, 32'hc3a8c4e4, 32'hc3fd1967},
  {32'h4511bc97, 32'h43e9894b, 32'hc11ccdd3},
  {32'h4234a820, 32'h41634bc6, 32'h43b8009d},
  {32'h44f40714, 32'hc3476843, 32'hc32dab65},
  {32'hc43d740e, 32'hc35a27e1, 32'h421f197e},
  {32'h44afb4b8, 32'h432ebf0a, 32'hc365d05e},
  {32'hc44c5852, 32'h43b7721f, 32'hc3355cb7},
  {32'h4305f140, 32'hc3de8f07, 32'hc3d24bfe},
  {32'hc3846e8c, 32'h4285448f, 32'hc3a599f9},
  {32'h44f0d314, 32'hc3dd4cba, 32'hc35ee2c4},
  {32'hc4a898ea, 32'hc2e6470d, 32'h43375fa5},
  {32'h4518f799, 32'h43533d56, 32'hbf4e342e},
  {32'hc4adad70, 32'h436c87b7, 32'hc39b4a3a},
  {32'h43e0bebc, 32'hc288dc77, 32'h43ccfb9a},
  {32'hc49c9bd2, 32'hc2b68006, 32'h4328439a},
  {32'h44a1768f, 32'h437ebe06, 32'h42b4b765},
  {32'hc4558bf6, 32'hc30de072, 32'h438d6d08},
  {32'h439f62e1, 32'h42e041d9, 32'hc3f34176},
  {32'hc49fc2aa, 32'hc280beb7, 32'hc288bb25},
  {32'h450fbde1, 32'hc324b09d, 32'h43227580},
  {32'hc50145f6, 32'hc31bff32, 32'h4414a7d1},
  {32'h4427fb2a, 32'h4395a182, 32'h42272631},
  {32'hc483a8c2, 32'hc1c093c9, 32'hc3886d70},
  {32'h443b3a9d, 32'hc2320f3e, 32'hc32270bd},
  {32'hc472d7be, 32'h4378f0cd, 32'h43cbd01f},
  {32'h44a73561, 32'hc2f2a688, 32'hc3996268},
  {32'hc429cb5b, 32'hc3840ea9, 32'h42cfa217},
  {32'h447cfd86, 32'h40634acd, 32'h42948ea6},
  {32'hc46cb735, 32'h414fe6de, 32'hc38ccb31},
  {32'h4491885c, 32'hc31b7afa, 32'hc28a9e7f},
  {32'hc441baa8, 32'hc220d121, 32'hc3e52663},
  {32'h4490de69, 32'hc3d57610, 32'h440260b6},
  {32'hc4f8306a, 32'hc21e02f2, 32'h42c9299a},
  {32'h434c2a48, 32'h4303b80c, 32'hc3115bb3},
  {32'hc3f95870, 32'hc2f2a845, 32'h42cbfb78},
  {32'h42c30118, 32'hc23edd3a, 32'hc34e6a97},
  {32'h43bf1828, 32'hc3595578, 32'hc280445c},
  {32'h45255c50, 32'h43c3cc6b, 32'h4421aa3c},
  {32'hc4abcabd, 32'h433814ae, 32'hc1b8db6c},
  {32'h44b302bf, 32'h43eac6d7, 32'hc3489e87},
  {32'hc4b26aa2, 32'h43b9543a, 32'hc26aaf3f},
  {32'h443a2052, 32'hc1b0dbd0, 32'h43728239},
  {32'hc445bd27, 32'h42560cfe, 32'h42610778},
  {32'h449a82b8, 32'h42ed893c, 32'hc32c3d01},
  {32'hc4665326, 32'hc2236518, 32'h42577ba0},
  {32'h44224a74, 32'hc2f6f0fa, 32'hc31b0196},
  {32'hc510176b, 32'hc23510a1, 32'h431fbd32},
  {32'h44fcbd66, 32'hc34b9b13, 32'hc19acfda},
  {32'hc511c4ed, 32'h42c5823e, 32'hc3e71bdb},
  {32'h437991e0, 32'hc38affe6, 32'hc338daf1},
  {32'hc44064ce, 32'h431f5833, 32'hc1e7913c},
  {32'h4509f576, 32'h42ce2186, 32'hc388c9f7},
  {32'hc3e43f1c, 32'hc3cb9667, 32'hc33115bc},
  {32'h4468708a, 32'hc31d2308, 32'h43d0e16e},
  {32'hc400e80c, 32'h429b9b40, 32'h43973134},
  {32'h43f4991a, 32'hc3051df3, 32'h42eb3267},
  {32'hc42d58b6, 32'h42d08318, 32'h43a23d20},
  {32'h44e4fa1c, 32'h43284b95, 32'h439b1eea},
  {32'hc4efce54, 32'hc3828d00, 32'h43ea4cac},
  {32'h44743289, 32'hc2f07314, 32'h42ec563c},
  {32'hc442e8f9, 32'hc1c7f6d5, 32'h4250a4f9},
  {32'h441671c8, 32'h4346b072, 32'h434b009d},
  {32'hc516b38e, 32'hc34bc434, 32'hc3395594},
  {32'h4515bed4, 32'h42231365, 32'hc354f936},
  {32'hc41f651c, 32'h4269b237, 32'h42ecd3ca},
  {32'h44f3e68f, 32'h436c78a0, 32'h42a27022},
  {32'hc519214e, 32'hc38f2bb2, 32'h43147efd},
  {32'h44a7b21e, 32'hc270a1a8, 32'h41304483},
  {32'hc3a933a8, 32'h437f4ee4, 32'hc2179466},
  {32'h45243e0c, 32'hc30ab74b, 32'h435cae36},
  {32'hc49e6371, 32'hc38a011d, 32'hc2e1a66f},
  {32'h4452b074, 32'h435d8d9a, 32'h43161267},
  {32'hc5045407, 32'h4168b4e6, 32'hc3554140},
  {32'hc3414ba9, 32'hc3629a5e, 32'hc3d5bfe6},
  {32'hc44a564a, 32'hc25b4f43, 32'hc11cb3ef},
  {32'h44c94522, 32'h42d94253, 32'h41587a96},
  {32'hc41f6a6b, 32'hc237109d, 32'hc34be606},
  {32'h4509b27a, 32'h430dac3d, 32'h42ee6866},
  {32'hc3c6c8fe, 32'h43bdb8ee, 32'h43b8f344},
  {32'h4500b66f, 32'hc296f116, 32'h42644eca},
  {32'hc4fa0d0e, 32'hc3352c74, 32'h43261fb3},
  {32'h44ef022b, 32'h42b1d6b1, 32'h427447b7},
  {32'hc2939e90, 32'hc251ee28, 32'h40d30454},
  {32'h4500b342, 32'hc2a0a897, 32'hc1a2361c},
  {32'hc32bd3d1, 32'h429e6c26, 32'h42aa1931},
  {32'h45032ab6, 32'hc3c72d11, 32'h42588980},
  {32'hc49e756a, 32'h4268466b, 32'hc3e83d8e},
  {32'h451e3e5d, 32'h432e61be, 32'hc2f47e8e},
  {32'hc3a9eca0, 32'hc2a43a47, 32'hc395f4f6},
  {32'h4494f3ca, 32'h4321203b, 32'h43146118},
  {32'h41849e80, 32'hc2719575, 32'hc3e48998},
  {32'h4521b6a0, 32'h4331f92f, 32'h428721b3},
  {32'hc465a820, 32'h421b85ba, 32'hc31bac95},
  {32'h45101139, 32'h42835034, 32'h424103c6},
  {32'hc4fe6d00, 32'h41bf110f, 32'hc390aba6},
  {32'h44bf6684, 32'hc22cf95c, 32'hc3605ba5},
  {32'hc4bb1239, 32'h426486eb, 32'hc37151b5},
  {32'h448533fe, 32'h42c5ff97, 32'h42fbcbfb},
  {32'hc502d25f, 32'h42da2269, 32'hc280ac44},
  {32'h448ee813, 32'hc3e0c1a3, 32'hc324cfe0},
  {32'hc506eebc, 32'hc0da426f, 32'hc285516a},
  {32'h44d27e75, 32'hc32429e6, 32'hc33602db},
  {32'hc501747b, 32'h41236bb9, 32'h423fe6ab},
  {32'h4492cb06, 32'hc2fdb015, 32'h43871b2a},
  {32'hc333852c, 32'h42008e74, 32'hc2c380a4},
  {32'h44477046, 32'h43a49aa9, 32'h42c2aff4},
  {32'hc420e98e, 32'hc3a2105e, 32'h43880d9a},
  {32'h45044a95, 32'h43808f1e, 32'h43685d29},
  {32'hc4d99d92, 32'hc302d226, 32'hc3503f9d},
  {32'h4310bf0c, 32'hc377059d, 32'h433b6635},
  {32'hc4d715e0, 32'h415ce2da, 32'h428e6bfb},
  {32'h450fd003, 32'hc3affd13, 32'h431e75b9},
  {32'hc3d1ce81, 32'h4285b1ab, 32'h4207ae6f},
  {32'hc127bfe0, 32'hc27b3044, 32'hc287b8af},
  {32'hc51659d6, 32'hc23f93b6, 32'hc2d9cf10},
  {32'h44fdeb3d, 32'hc2248d68, 32'h428c2da4},
  {32'hc522b16a, 32'h420c6f0e, 32'hc25801f2},
  {32'h43c0f442, 32'h438dcff2, 32'hc38b6e97},
  {32'hc47ca78a, 32'hc2eab9fa, 32'h42466d0d},
  {32'h45071455, 32'hc284339e, 32'h42b70a44},
  {32'hc4210ccf, 32'hc359b0c2, 32'h4312f0ba},
  {32'h452d8897, 32'h43b74718, 32'h42fb6098},
  {32'hc5119074, 32'h42b8e5fe, 32'h40ac95b4},
  {32'h441cbc77, 32'h421e1e9b, 32'h4280ccd1},
  {32'hc41a222c, 32'h42c697fc, 32'h416adb08},
  {32'h45142cc8, 32'h4201c61f, 32'h42cea246},
  {32'hc513c7af, 32'hc29f7caa, 32'hc32c889b},
  {32'h450c752a, 32'h44055291, 32'hc3014a7e},
  {32'hc5032cea, 32'hc1d5ed0e, 32'hc2187494},
  {32'h44a01192, 32'h433c4cf6, 32'h4395d704},
  {32'hc2c6f250, 32'hc3012225, 32'hc36e6d40},
  {32'h451570f0, 32'hc36bda75, 32'h43245216},
  {32'hc4ec8946, 32'h43041ed3, 32'hc327b21e},
  {32'h43e3ffbc, 32'h43903912, 32'h433ed29b},
  {32'hc5092775, 32'hc2d4f59d, 32'h426250f3},
  {32'h435e4e8f, 32'h4295612d, 32'hc33c8228},
  {32'hc37f7c88, 32'hc3180349, 32'hc3a44af5},
  {32'h44e1e9d1, 32'h43158533, 32'h437a4110},
  {32'hc42e9b3c, 32'h438aaf23, 32'hc2715298},
  {32'h433b6390, 32'h43bf0232, 32'hc36b4efe},
  {32'hc4a6be51, 32'hc39c6499, 32'h41f4a785},
  {32'h44fd62e1, 32'h41be0467, 32'hc41358b4},
  {32'hc4df9a44, 32'hc31dd3ea, 32'h41ac9550},
  {32'h44f38660, 32'h43885d6b, 32'hc3554f18},
  {32'hc42b1f1d, 32'hc30a6a79, 32'hc3c5c6f7},
  {32'h44cb2c94, 32'hc3be8689, 32'h43939a81},
  {32'hc4eef170, 32'h433367a0, 32'h42811bc1},
  {32'h449aed7f, 32'h43571811, 32'h432a26e6},
  {32'hc35d74c8, 32'hc262c108, 32'hc363b09f},
  {32'hc3440580, 32'hc3958802, 32'hc2cdb806},
  {32'hc2a17e00, 32'hc19cf7d6, 32'hc3c83194},
  {32'h450dd507, 32'h438c9923, 32'h43da5dac},
  {32'hc38434d4, 32'hc2e44c4b, 32'hc3eb2cfa},
  {32'h45076684, 32'h4338a411, 32'h43e8cd7a},
  {32'hc516fef5, 32'h4301b8c0, 32'hc394c104},
  {32'h44890352, 32'h434d1b4e, 32'hc2805ba0},
  {32'hc35a8204, 32'hc2b1f2ff, 32'hc395e542},
  {32'h43a74780, 32'h435d750c, 32'hc19bcb09},
  {32'hc3abec37, 32'hc21c927d, 32'hc3644e3a},
  {32'h441b84de, 32'hc13a9604, 32'h439477fa},
  {32'hc4fad0b0, 32'hc360c040, 32'hc2408d2f},
  {32'h428430f8, 32'hc3655399, 32'hc284d1bb},
  {32'hc4ad94f9, 32'h43127f19, 32'h43ca53b3},
  {32'h45003cda, 32'h42bc87e0, 32'hc30d26ef},
  {32'hc49612b9, 32'hc3991693, 32'hc34d4dea},
  {32'h43ece258, 32'h43726400, 32'h42bb9090},
  {32'hc5078e33, 32'h43427df6, 32'h42a99d76},
  {32'h413d3e50, 32'hc306a867, 32'hc2b2f57d},
  {32'hc457de06, 32'hc3ce7f4d, 32'h427e5354},
  {32'h448aff27, 32'h43a4e4ab, 32'hc2690eb5},
  {32'hc3b1900a, 32'hc2c46f49, 32'h4237f4eb},
  {32'h44a7349b, 32'hc2592191, 32'h43f6325c},
  {32'h41cd5b00, 32'hc0de09d8, 32'hc3b68631},
  {32'h4451818e, 32'h42e1f4a5, 32'hc2566750},
  {32'hc48cf9fa, 32'h4217e377, 32'hc2f61824},
  {32'h44e1e98f, 32'hc158058e, 32'hc3f59ed2},
  {32'hc4cdf4be, 32'hc35ef13b, 32'hc2f364a7},
  {32'hc333c948, 32'hc3701cdf, 32'h434591c7},
  {32'hc30fa388, 32'hc26a5c80, 32'hc2aad971},
  {32'h4501b9cf, 32'h426acd39, 32'h4255853d},
  {32'hc4c6e7db, 32'hc2c4626e, 32'hc30f0387},
  {32'hc21de070, 32'hc30cf11d, 32'hc3907cbf},
  {32'h4512c35f, 32'hc3950cd2, 32'h427c9e34},
  {32'hc4df1928, 32'h43237eed, 32'hc1ea00ec},
  {32'h44f90a12, 32'h438a0e62, 32'hc2f10ed0},
  {32'h41a95f6d, 32'hc403e505, 32'h4280bfb2},
  {32'h446b3df8, 32'hc37c172b, 32'h43aa332f},
  {32'hc5083d92, 32'h43c8a073, 32'hc286f772},
  {32'h4455a0a2, 32'h43269122, 32'h4310439e},
  {32'hc4672543, 32'h42f9a954, 32'h428e621a},
  {32'h44ebfa01, 32'hc28fa333, 32'h41a45736},
  {32'hc4c9e1de, 32'h438186d5, 32'hc362d1f4},
  {32'h4495c09e, 32'hc3b2dc93, 32'hc2eac04c},
  {32'hc483a10c, 32'h438dbf30, 32'h428c853e},
  {32'h44bad555, 32'hc36e343e, 32'hc2990834},
  {32'hc47455ba, 32'h434907de, 32'hc2c328dc},
  {32'h450b5940, 32'h432513d4, 32'h4347e86c},
  {32'hc4f4fcf1, 32'h42486575, 32'h42976d53},
  {32'h4518fb1f, 32'hc32bb44b, 32'h4273eef2},
  {32'hc43f5e3c, 32'h436ddfb0, 32'h41758f4c},
  {32'h445a11f4, 32'h42fcd98f, 32'h43c66736},
  {32'hc42f854c, 32'hc33516de, 32'hc2fa6f5e},
  {32'h44e60731, 32'hc24a9e8c, 32'h43065885},
  {32'hc44f9a64, 32'hc2b1d3f6, 32'hc345dfc8},
  {32'h4441a173, 32'h4267b18a, 32'h43358e4e},
  {32'hc49da1ce, 32'hc3ee5f94, 32'h4306971b},
  {32'h43c24650, 32'h438894e0, 32'hc2fb522d},
  {32'hc48bfb64, 32'hc25e717c, 32'hc3a0d7eb},
  {32'h4516a70f, 32'hc3d30768, 32'h4208b6aa},
  {32'hc4e12879, 32'hc389e264, 32'hc3ef3228},
  {32'h450efca2, 32'hc3898587, 32'h427a2e0c},
  {32'hc3223258, 32'hc017308b, 32'hc38043de},
  {32'hc3cfbe50, 32'hc37000dd, 32'h42e068a5},
  {32'hc42d3cc4, 32'hc38c5b1a, 32'h42a15283},
  {32'h4494ddac, 32'hc2ff9994, 32'hc226b8fa},
  {32'h431775c3, 32'hc2a09f0a, 32'hc22f8bf9},
  {32'h450617a4, 32'hc34c017b, 32'h437b616e},
  {32'hc43c2d6f, 32'hc307ccb2, 32'h42afbdb1},
  {32'h4429fa74, 32'h43490877, 32'hc2ba409a},
  {32'hc45730e4, 32'hc380a81c, 32'h4300f147},
  {32'h44ad76d8, 32'hc1a46546, 32'hc1972a2a},
  {32'hc3e805dc, 32'hc38fb057, 32'h439a2e82},
  {32'h44e9324d, 32'hc300b9b8, 32'h426fd5a4},
  {32'hc44f6382, 32'hc286c5f1, 32'h423753f1},
  {32'h44c2d147, 32'hc41b39a0, 32'h438c7ff7},
  {32'hc4a6f480, 32'h434168a2, 32'h42aaf57e},
  {32'h44c059d6, 32'h4251db28, 32'hc3452d33},
  {32'hc3b48758, 32'hc2071ec4, 32'h427ab870},
  {32'h436338b1, 32'h4427ee55, 32'h431318b9},
  {32'hc48b79f6, 32'hbefe3640, 32'hc2fe560a},
  {32'h448faf0c, 32'h41c35a91, 32'h41635c4d},
  {32'hc45a4c0a, 32'h439e39ab, 32'hc25d6060},
  {32'h4357b8f0, 32'hc2300edf, 32'h428f9b92},
  {32'hc47781fd, 32'hc1139c52, 32'h4319a5f5},
  {32'h44caf48a, 32'hc33c8ed1, 32'h436af1eb},
  {32'hc493446c, 32'hc3d70cea, 32'hc391d7a9},
  {32'h433c2f3a, 32'hc35ab4c6, 32'hc3dfbce5},
  {32'hc27c7167, 32'hc395d4b5, 32'h4348fdd7},
  {32'h450e9202, 32'hc3939297, 32'hc3c49e9d},
  {32'hc3fd9c13, 32'hc343c0ca, 32'h433e841f},
  {32'h448ade0c, 32'hc3844828, 32'h433ccd1b},
  {32'hc4cf23a4, 32'hc2c1f7ed, 32'hc241e0ea},
  {32'h43e6dd65, 32'hc2ad43ab, 32'hc37ad504},
  {32'hc5092ae1, 32'hc3a2b255, 32'hc3793027},
  {32'h4406d34e, 32'hbf37b1b0, 32'h42ab6b63},
  {32'h42c8cd60, 32'hc33446ac, 32'h43946f67},
  {32'h448c9798, 32'hc35d193a, 32'h430b2385},
  {32'hc51092b8, 32'hc3082e59, 32'hc29a30d2},
  {32'h426ebe60, 32'h4370220c, 32'hc31d976c},
  {32'hc4b9440b, 32'hc3216422, 32'hc34b8e07},
  {32'h43b2d820, 32'hc3465904, 32'h43e66c09},
  {32'hc5030773, 32'hc34e2470, 32'h421eddd2},
  {32'h44882a1a, 32'hc304bf4b, 32'h433bf6c3},
  {32'hc4d20a96, 32'hc2b28202, 32'h42dd0b14},
  {32'h444d9190, 32'h43086be8, 32'hc2e2bc57},
  {32'hc50140b1, 32'hc313474f, 32'h42f12b10},
  {32'h42fa9f04, 32'hc181313a, 32'hc3284357},
  {32'hc50a9141, 32'h43c20668, 32'hc209c7b7},
  {32'h44a19268, 32'hc2084dff, 32'hc38c2f26},
  {32'hc287e8c0, 32'hc25d11b8, 32'hc38d24f1},
  {32'h44e01c13, 32'h42c91c3a, 32'h434922a8},
  {32'hc4b36eb6, 32'h43a2fc81, 32'hc392f85c},
  {32'h4436eaa8, 32'hc26423c7, 32'hc22c4c73},
  {32'hc4e4a29a, 32'hc2957a7a, 32'h43643d39},
  {32'h4502579b, 32'h439256b6, 32'h43a30dd6},
  {32'hc28da460, 32'hc143b5c6, 32'h418f3b2d},
  {32'h430149a4, 32'hc1d34bf6, 32'hc1adce24},
  {32'hc4826e7b, 32'h436b9530, 32'h432ece4b},
  {32'h44e324b2, 32'hc23196de, 32'hc3032005},
  {32'h433d05a8, 32'h42800ccf, 32'h431c246c},
  {32'hc0fca100, 32'hc2da5743, 32'hc35bf194},
  {32'hc2fa76f4, 32'hc3bef5da, 32'hc2d6340d},
  {32'h41913880, 32'hc28f8024, 32'hc22b458a},
  {32'hc5005935, 32'hc35900f3, 32'hc28af923},
  {32'h43810fe0, 32'hc3486442, 32'hc3f568ae},
  {32'hc4c34847, 32'hc2df6f95, 32'hc30a4605},
  {32'h450549e8, 32'hc19a0bbc, 32'h42233471},
  {32'hc4e3e9fd, 32'h411994c8, 32'hc2d9b7c9},
  {32'h4475f22e, 32'hc31a992f, 32'hc352cce6},
  {32'hc43066e9, 32'h44039f7c, 32'h414cee71},
  {32'h448e7423, 32'hc3b97d22, 32'h431dc6b6},
  {32'hc45050f7, 32'h439a1fce, 32'h4179dded},
  {32'h44bf86da, 32'h428848e7, 32'h421d1809},
  {32'hc422a97a, 32'h4332989c, 32'hc3a598d2},
  {32'h43fac254, 32'hc35737ab, 32'h442b9eee},
  {32'hc4e9dda8, 32'hc3ebc7fc, 32'hc3338e56},
  {32'h439b63f8, 32'hc1bb1b32, 32'hc290ab25},
  {32'hc37f2ea0, 32'hc3e6cab2, 32'hc302c4b1},
  {32'h42465d88, 32'h40cc35b6, 32'hc398de5b},
  {32'hc508b299, 32'hc3d58af7, 32'h43505b69},
  {32'h44cc78e6, 32'h42d849dc, 32'h42a1eeb5},
  {32'hc5116af3, 32'hc3c5fda7, 32'hc33b3fce},
  {32'h44a185c2, 32'h43944aef, 32'h43271709},
  {32'hc351cd50, 32'hc3b174b0, 32'h42f360c2},
  {32'h44be7d2e, 32'h4345733f, 32'hc301f211},
  {32'hc40cae1e, 32'hc3acd72f, 32'h42d919ab},
  {32'h42814fd4, 32'hc437f1d5, 32'hc3669c6c},
  {32'h44e1eb4e, 32'hc30a9927, 32'hc31e3532},
  {32'hc4d38e46, 32'h439b1e52, 32'hc3c2aa46},
  {32'h4421f0a4, 32'hc16a326f, 32'hc2b86588},
  {32'hc343f16c, 32'h437d966a, 32'h42cdb806},
  {32'h4506a457, 32'h430c8d22, 32'h43eb3cea},
  {32'hc48297cd, 32'h4372300a, 32'hc2c89eb6},
  {32'h44574a38, 32'hc1c42043, 32'hc29d7fad},
  {32'hc4596b40, 32'h428a48d1, 32'h438135ae},
  {32'h44651bf4, 32'hc186ec42, 32'h42fab44e},
  {32'hc4a599c6, 32'hc0ff7e0f, 32'h420d1203},
  {32'h450c06e1, 32'hc2ff63db, 32'h4336c8e3},
  {32'hc38ba9dc, 32'hc3410fd8, 32'hc2a9dfda},
  {32'h445f7822, 32'hc213e7e7, 32'hc208fcc4},
  {32'hc4d8e708, 32'hc3ab4003, 32'h4385d450},
  {32'h44873dd3, 32'hc39c5c8e, 32'h42f5d5d4},
  {32'hc4915307, 32'hc343e4a4, 32'h43878a3b},
  {32'h44d2ca71, 32'hc329832c, 32'h437903ae},
  {32'hc28f33e0, 32'hc11b8f82, 32'hc397f416},
  {32'h440694ec, 32'hc3027dd0, 32'hc362ae2a},
  {32'hc4c8bee5, 32'hc23e9e2d, 32'hc2925ed3},
  {32'h442160b0, 32'hc2c0aa27, 32'h42cbf658},
  {32'h43260462, 32'hc3b7f94e, 32'hc0eb345d},
  {32'h44de6de4, 32'h438f8ff2, 32'hc32c243b},
  {32'hc44b8671, 32'h43a1f7c6, 32'hc3249808},
  {32'h4429590d, 32'hc38fb2ea, 32'hc2216521},
  {32'hc481ffc6, 32'hc3713844, 32'hc2a78eec},
  {32'h447190f0, 32'hc2360dc3, 32'hc20d48f0},
  {32'hc4f58784, 32'h43ae78e8, 32'h4398a02c},
  {32'h44e52647, 32'h42934d2f, 32'h4364e210},
  {32'hc4e1451c, 32'hc3012707, 32'hc101af19},
  {32'h44f2505a, 32'hc309553d, 32'hc267bca3},
  {32'hc48485e0, 32'hc395c6e8, 32'hc33fe657},
  {32'h442cbfde, 32'h42063378, 32'hc397c543},
  {32'hc50b10d2, 32'h42c3b57a, 32'hc3845a4c},
  {32'h4415e112, 32'h42a8285f, 32'h41e95036},
  {32'hc4305f3f, 32'hc36dedd6, 32'h428a0ffa},
  {32'h44a66c9f, 32'hc246ed7f, 32'h40cfb020},
  {32'hc3687d2f, 32'hc2d8e02a, 32'hc276794f},
  {32'h44eb613a, 32'hc3131d1a, 32'h423ce28e},
  {32'hc3e9bddc, 32'h437f7e64, 32'hc310b00a},
  {32'hc2d6f390, 32'hc2658e3c, 32'hc415303f},
  {32'hc4ce9cc3, 32'h439c6346, 32'hc2e872dd},
  {32'h438f47c3, 32'hc389c749, 32'h4329dac2},
  {32'hc510c697, 32'h43224027, 32'h428901d4},
  {32'h44b486e0, 32'hc33419d9, 32'h428247ea},
  {32'hc4e327a3, 32'hc3c6094d, 32'hc38b42b4},
  {32'h449cd1b2, 32'hc1a12905, 32'h434b2156},
  {32'hc497816c, 32'hc3696977, 32'hc3405675},
  {32'h42b90ba8, 32'h42174b6c, 32'hc35c71cb},
  {32'hc48203b6, 32'h4398907a, 32'h422d5c16},
  {32'h43247989, 32'hc41fa1fa, 32'h42c5d1fe},
  {32'hc4cd0e90, 32'h430d4026, 32'h43063da8},
  {32'h45020db4, 32'hc301f1a4, 32'h42f30d75},
  {32'hc4d4a2bc, 32'h429608f7, 32'hc12dd34b},
  {32'h449c1fd1, 32'hbf4077c0, 32'h41efb8fc},
  {32'hc499290e, 32'hc2bc4d89, 32'hc35e302d},
  {32'h4444623c, 32'h42707270, 32'h43a413ae},
  {32'hc42f1ea0, 32'h4320934e, 32'h3e241600},
  {32'h44e52e63, 32'h43c5e1b9, 32'hc1845459},
  {32'hc4cb48f6, 32'hc204648d, 32'h434af71e},
  {32'h4513d4c4, 32'h40bbc8ed, 32'h432f49b6},
  {32'hc4dd4cef, 32'hc338dfed, 32'h4187de7d},
  {32'h441f033e, 32'h41b25ed9, 32'hc3660cbe},
  {32'hc46cea22, 32'h432f4fff, 32'h42976b82},
  {32'h44b79f0f, 32'h433383ff, 32'hc190f8f7},
  {32'hc45889e6, 32'h43c1a54c, 32'hc2b4e0fd},
  {32'h43970405, 32'h43e36deb, 32'hc374e48c},
  {32'hc5077893, 32'hc316ebb2, 32'hc1fb4122},
  {32'h4471d6e3, 32'h43e9e69f, 32'h43b5d5f5},
  {32'hc503949c, 32'hc392d4d4, 32'hc22801b2},
  {32'h4342e334, 32'h43a41b99, 32'h4031c8af},
  {32'hc427cfdd, 32'hc29f31c4, 32'h439128b4},
  {32'h3d8bc800, 32'hc182a3fd, 32'hc2e8ae5d},
  {32'hc4f66b7a, 32'hc296d848, 32'hc2f1a6de},
  {32'h449855b9, 32'h4355bde3, 32'hc239d990},
  {32'hc4c15d65, 32'h4214951c, 32'h438d5558},
  {32'h4516070b, 32'h428e2a70, 32'h4373df79},
  {32'hc4d78f5f, 32'h4089a91b, 32'hc38ab953},
  {32'h442adc3a, 32'h4331aaea, 32'hc37baae3},
  {32'hc3fa3728, 32'hc3769f25, 32'h42b24347},
  {32'h44b09930, 32'h43bb9917, 32'h43b566a3},
  {32'hc4addf44, 32'hc4256ff4, 32'hc1b2b8ac},
  {32'h44e5fd67, 32'h4390c4f3, 32'h42b8515a},
  {32'hc42070f6, 32'hc2858a24, 32'hc37331a8},
  {32'h44fb5b5c, 32'h437f4200, 32'hc30ab4e4},
  {32'hc5003cd0, 32'hc3b2f281, 32'h42b90867},
  {32'h45097b82, 32'hc26fb5c8, 32'h43257d07},
  {32'hc4956d71, 32'h4115a5b5, 32'h430a188d},
  {32'h44f9c8aa, 32'hc20495b3, 32'hc3191490},
  {32'hc3961628, 32'h428ea00d, 32'hc118ec72},
  {32'h450a0702, 32'hc1b9726c, 32'h43aded09},
  {32'hc4df97b4, 32'h41ec5d3d, 32'hc3b03114},
  {32'h447bfbec, 32'hc36fd28b, 32'hbe5b14a8},
  {32'hc4b45d9d, 32'hc32fa4e1, 32'h4403f76b},
  {32'hc2f6efd0, 32'h43778ea6, 32'h43dbd635},
  {32'hc495c416, 32'h4395ab66, 32'h430d29fc},
  {32'h44e56557, 32'hc2871186, 32'h439425ff},
  {32'hc4623720, 32'h42e99a68, 32'hc34ebaf3},
  {32'h44e43b54, 32'h42add011, 32'h433afb1c},
  {32'hc4b3546e, 32'hc1b815d9, 32'h436d9900},
  {32'h44c5068f, 32'hc3026af9, 32'hc3495562},
  {32'hc42bf080, 32'hc31f01e3, 32'hc196d3de},
  {32'h43e70fd8, 32'hc18d4b9c, 32'h43cbaa94},
  {32'hc39a2e10, 32'hc3dfb65f, 32'h42f24ff8},
  {32'h44c66840, 32'hc288f825, 32'h42c69000},
  {32'hc4bea18d, 32'hc33efd52, 32'h43af42f9},
  {32'h44acfd84, 32'h4313d143, 32'hc3624661},
  {32'hc4eed4dd, 32'hc377ed5b, 32'hc2fa9aa0},
  {32'h4437bbfb, 32'h42ce4465, 32'h43f04ca9},
  {32'hc50c0309, 32'h42d2ee87, 32'h43c854cb},
  {32'h440edb56, 32'hc30ad0d9, 32'hc3cd82a4},
  {32'hc3c88700, 32'h430c2513, 32'h4116aa00},
  {32'h44db0e54, 32'h4399599a, 32'hc305ceac},
  {32'hc4f5f0c6, 32'hc2fdad55, 32'hc314224b},
  {32'h44eec175, 32'h428cd4a2, 32'hc3a73ca8},
  {32'hc4c34069, 32'hc31d6f1e, 32'hc33051dd},
  {32'h44a80811, 32'h43229e54, 32'hc1f7dc30},
  {32'hc3d64600, 32'h3d845900, 32'hc33f94b5},
  {32'h44bb4435, 32'hc35c1126, 32'h420f69b9},
  {32'hc4a82423, 32'h4195e709, 32'h419744b6},
  {32'h43ef747e, 32'h43a9961a, 32'h431a5a62},
  {32'hc4d87a05, 32'h4293727e, 32'hc3367ca6},
  {32'h44e0bd1c, 32'h4165d259, 32'h437631e6},
  {32'hc334c8f8, 32'h4278d274, 32'h41e6c835},
  {32'h44f0c7e6, 32'h43ca2488, 32'h4261b24f},
  {32'hc460a750, 32'h429777e2, 32'hc235d0e9},
  {32'h42f97518, 32'h4338f37f, 32'h41beae07},
  {32'hc2792e20, 32'h43bfe542, 32'h42b3267d},
  {32'h4502de21, 32'h4322604d, 32'h401bfe95},
  {32'hc318ac30, 32'hc25b735e, 32'h43364180},
  {32'h44a36359, 32'hc36aa0dc, 32'h4309f291},
  {32'hc4ba0fce, 32'hc311e9ce, 32'h42c44bd2},
  {32'h44f11e0e, 32'hc224cacc, 32'hc3860c12},
  {32'hc4a9b243, 32'h4322f8af, 32'hc3217c59},
  {32'h43b40403, 32'hc2518a26, 32'h436d8a95},
  {32'hc18eeeb5, 32'hc37a6e1a, 32'h42ab49b7},
  {32'h44bec9dc, 32'h4357f80c, 32'h423cefd1},
  {32'hc46207ac, 32'h4369018c, 32'h4392b678},
  {32'h450466ef, 32'h42fdf435, 32'hc18b2678},
  {32'hc4bfa221, 32'hc2afbad8, 32'h4329cfdd},
  {32'h44db3ad4, 32'h435dfba6, 32'h435ecc07},
  {32'h43d20238, 32'h4209eeb6, 32'h43b33053},
  {32'h4485f492, 32'hc2f1d738, 32'h43634747},
  {32'hc43af47e, 32'h4262ab96, 32'h42a6bb06},
  {32'h446e8e84, 32'hc2e501b2, 32'h43652996},
  {32'hc4f1bbef, 32'hc2acf540, 32'h42e2629b},
  {32'h44b72497, 32'h436b6371, 32'hc31a72db},
  {32'hc36b7180, 32'h41f629c2, 32'hc35ac302},
  {32'h448af1e6, 32'hc35eb8e3, 32'h439c3134},
  {32'hc427710e, 32'hc2564046, 32'hc30fe32e},
  {32'h44994b90, 32'hc32ff269, 32'h410e160b},
  {32'hc40afbb4, 32'hc28db755, 32'hc384f654},
  {32'h44485010, 32'hc2ea2f9f, 32'hc24ff271},
  {32'hc2988382, 32'hc246bd55, 32'hc20b49dd},
  {32'h451f8ef8, 32'h418a6ba2, 32'h438b3272},
  {32'hc4a8cdeb, 32'h42edefc3, 32'hc23cf8af},
  {32'hc28f98f2, 32'hc23c7004, 32'hc36889ae},
  {32'hc3fb3aab, 32'hc3167a57, 32'hc3168f2c},
  {32'h442546a6, 32'hc3456582, 32'h4380d659},
  {32'h418c02d7, 32'h41d23c31, 32'h42a4e488},
  {32'h44948c08, 32'h4278b1ca, 32'h431f9e7e},
  {32'hc4d0c2d6, 32'h430c1ac6, 32'h413c3082},
  {32'h44e77b33, 32'h438e6d4b, 32'h438811d8},
  {32'hc3d58ed4, 32'h43b537cd, 32'h4227434e},
  {32'h4487d1ff, 32'h41fb315c, 32'hc3c6a222},
  {32'hc47d3ab0, 32'h4330453f, 32'hc303149c},
  {32'h44689e0d, 32'hc30b5d72, 32'h43212d0a},
  {32'hc51a0c27, 32'hc2f5704a, 32'h43a02caf},
  {32'h440ba992, 32'h42a06617, 32'h43a2a769},
  {32'hc47e0387, 32'hc2f93b6a, 32'h41d0de31},
  {32'h43cfd06c, 32'h42c70998, 32'h431952b5},
  {32'hc4acd78a, 32'hc2ead53f, 32'hc29faed9},
  {32'h449f431c, 32'h433bfb42, 32'h430568a3},
  {32'hc4e41091, 32'hc307dc81, 32'hc36af09a},
  {32'h44dfa3e8, 32'h432ae1a6, 32'hc3b95db2},
  {32'hc4234a82, 32'hc36a0b07, 32'h418d93de},
  {32'h44b567ad, 32'h43f0fc7a, 32'h43239e7d},
  {32'hc4e8a436, 32'hc3831677, 32'hc3899f35},
  {32'h443283b2, 32'h4299fb5a, 32'h41f63b2e},
  {32'h42cdaae4, 32'h43b79f06, 32'hc281042b},
  {32'h44d40657, 32'h43aaaa29, 32'hc2fc22f9},
  {32'hc5024a14, 32'h415bf2b7, 32'h440bb8f4},
  {32'h42aa1010, 32'hc375f8a3, 32'h43e17041},
  {32'hc49582a3, 32'h4304c9b2, 32'hc35fad90},
  {32'h448f3c00, 32'h4400192b, 32'hc3907e3d},
  {32'hc4e1c5c2, 32'hc3c45951, 32'hc1759a5c},
  {32'h4420d446, 32'hc314777f, 32'h43866033},
  {32'hc2cee646, 32'h42e2e344, 32'h43ab6bfc},
  {32'hc3876023, 32'h41fc35e0, 32'h409dd21e},
  {32'hc4166b98, 32'h43403b76, 32'hc3917c2a},
  {32'h4493ccdf, 32'h42b57b2e, 32'hc329aaca},
  {32'hc3959bc8, 32'hc396d3f7, 32'h4362ffc4},
  {32'h451fe342, 32'hc3129b5c, 32'h4381bc3e},
  {32'hc3812b5e, 32'hc37c7b18, 32'h428b378d},
  {32'h4497d52d, 32'h42fed4ef, 32'h421bfa46},
  {32'hc3b045c6, 32'hc26a8322, 32'h43ac5b7e},
  {32'h44288cf8, 32'hc38954dc, 32'h4334b030},
  {32'hc521a69d, 32'h43390ce0, 32'hc337f12c},
  {32'h4496521a, 32'hc266511a, 32'h43bce156},
  {32'hc4b1de64, 32'hc31ca1bf, 32'hc3c05518},
  {32'h451776e8, 32'hc2ea0df2, 32'hc38dcab3},
  {32'h42fa3898, 32'h41815070, 32'hc18230ff},
  {32'h44b9c849, 32'h43c95ce2, 32'h43ccd83d},
  {32'hc49d74ba, 32'h440ed10d, 32'h43a05bfc},
  {32'h44df3ae0, 32'hc411cd06, 32'h4303207c},
  {32'hc4606b86, 32'h43eb5b02, 32'hc31b04f5},
  {32'h450f0ac9, 32'h43f01f77, 32'hc2fd628a},
  {32'hc46db4d0, 32'hc2a2a138, 32'hc2ad713b},
  {32'h44d4e874, 32'hc36558b3, 32'h43c869ec},
  {32'hc41caaa8, 32'h42159884, 32'hc3c0bf67},
  {32'h45146354, 32'hc026f956, 32'hc330002b},
  {32'hc4397a62, 32'h430d9b70, 32'h41925e80},
  {32'h43abfe3b, 32'h42041991, 32'h4302d502},
  {32'hc48a4db4, 32'hc2e509a5, 32'hc3623143},
  {32'h43b690a0, 32'h4387c90f, 32'hc3165f9b},
  {32'hc50d242e, 32'hc30bd330, 32'hc2e5fde3},
  {32'h44b5a2db, 32'hc35d2d11, 32'h423aedad},
  {32'hc466087a, 32'hc2de7201, 32'hc307ec56},
  {32'h4436c079, 32'hc354c418, 32'h43294ba4},
  {32'hc4a4333b, 32'h4046ef78, 32'hc3115571},
  {32'h450ce02b, 32'h43e9c288, 32'h4322b854},
  {32'hc4fe56ef, 32'hc2592bb2, 32'h434dadfd},
  {32'h451bf809, 32'hc2c4ea10, 32'h437c2534},
  {32'hc503006b, 32'hc3650d9f, 32'hc385f6ae},
  {32'h4423ff74, 32'hc3ac2433, 32'hc2d6a69a},
  {32'hc4e5f7db, 32'h4068ada8, 32'h42006609},
  {32'h44d18f45, 32'hc32c477c, 32'h428b9c34},
  {32'h431e99bf, 32'h4356238e, 32'hc38ac9eb},
  {32'h43dd93f4, 32'h413c06e2, 32'h43777651},
  {32'hc518b9df, 32'h41b7d6f7, 32'h4312b6d8},
  {32'h4428792c, 32'hc304d9a4, 32'h43088b4d},
  {32'hc3ba1f0b, 32'hc3270bc0, 32'hc33e65d0},
  {32'h448ab898, 32'hc3289fb2, 32'h42fab82b},
  {32'hc37f4dc0, 32'hc362ab84, 32'h43fa2028},
  {32'h4499018f, 32'hc310eed9, 32'h428dde51},
  {32'hc4f6c9b2, 32'hc4185167, 32'hc4001018},
  {32'h443ed3a8, 32'hc388c707, 32'hc1d37b12},
  {32'hc5172932, 32'hc0ad4f54, 32'h43176b12},
  {32'h449813a8, 32'hc2cca2c5, 32'hc2f404b8},
  {32'hc3e581ec, 32'h435b745d, 32'hc2cfc5b0},
  {32'h442f8866, 32'hc332e760, 32'hc371860d},
  {32'hc507ea9c, 32'hc1654238, 32'hc3601f8a},
  {32'h44345c4b, 32'hc2f836eb, 32'h43568856},
  {32'hc4fe6658, 32'hc3e8286b, 32'hc31cfa91},
  {32'hc28fb3f0, 32'hc32ae8e5, 32'hc3c66c1a},
  {32'hc4dc8459, 32'hc388068b, 32'hc3de0b2d},
  {32'h44f34218, 32'h430fef18, 32'hc308cf64},
  {32'hc414a120, 32'hc2009b84, 32'hc38000c9},
  {32'h447a7eb5, 32'h43700795, 32'hbeffc310},
  {32'hc48a1cd7, 32'hc382700f, 32'h43963a7a},
  {32'h4328c6c2, 32'hc32d5236, 32'hc370a659},
  {32'hbf1a5000, 32'h43bb4aa6, 32'h43e34847},
  {32'h449d2968, 32'h43bd45e8, 32'h433e35f6},
  {32'hc4a638f3, 32'hc21a3fc9, 32'hc2b24457},
  {32'h448b3df1, 32'h437ec885, 32'hc3231f3c},
  {32'hc4b28156, 32'h4319afe0, 32'hc358337e},
  {32'h448df90a, 32'h43a9b02d, 32'h41a8f00f},
  {32'hc450b7c7, 32'h43ca4131, 32'hc28159ad},
  {32'h4486eba3, 32'hc33a0264, 32'hc2f4b523},
  {32'hc38a2490, 32'h43a77ef3, 32'h421f4952},
  {32'h43ca0508, 32'h43c24aac, 32'hc130a284},
  {32'hc4f1597b, 32'hc25953d7, 32'h42aee1a3},
  {32'h41439670, 32'h426f1cb4, 32'h43411ffa},
  {32'hc474d84d, 32'h428a6003, 32'h4401ccff},
  {32'h44f69048, 32'h41915231, 32'h42c31c16},
  {32'hc4c2c6f5, 32'h41c7f43d, 32'h43355b0f},
  {32'h44108338, 32'h439b1fc0, 32'hc22e88c2},
  {32'hc39cfd24, 32'hc30bc632, 32'hc3021953},
  {32'h44bb5513, 32'hc351e5e7, 32'h436a398c},
  {32'hc508a7e3, 32'h4330d3ff, 32'hc2b17f78},
  {32'h43b8da8c, 32'hc2f6ee85, 32'h421abb52},
  {32'hc4910a78, 32'hc3a90586, 32'hc30152e3},
  {32'h443a0655, 32'h42aaf170, 32'hc2326896},
  {32'hc4b63940, 32'hc2cb5c81, 32'h41d0bd9e},
  {32'h44889ed4, 32'hc352dce7, 32'h4209ebfa},
  {32'hc4484080, 32'h4389126e, 32'h409e958c},
  {32'h43ddbf07, 32'hc39032df, 32'hc3b2a866},
  {32'hc396ae14, 32'h435091d6, 32'h419873fc},
  {32'h4423794e, 32'hc2449a78, 32'hc2f02787},
  {32'hc4e955be, 32'h42d5671d, 32'hc3f0f2d2},
  {32'h44437de4, 32'hc25d2f1f, 32'hc19d05ae},
  {32'hc5126e59, 32'h4296b979, 32'h43772934},
  {32'h444421d8, 32'hc28b1d5e, 32'hc3aa1626},
  {32'hc4ec8aa2, 32'h42d267f0, 32'hc361cbc1},
  {32'h44a8c028, 32'hc26e8f27, 32'hc3c1f21e},
  {32'hc465be6a, 32'hc211927d, 32'h4134d1b2},
  {32'h44289a60, 32'h43aaeafe, 32'hc3971428},
  {32'hc4aef372, 32'hc2f7a680, 32'h42e82eef},
  {32'h44ed06c4, 32'h430f58ce, 32'h435e3bb9},
  {32'hc3dbdc78, 32'hc14620db, 32'hc14183c0},
  {32'h44c732a1, 32'h40187c8c, 32'hc409f57e},
  {32'hc3974e43, 32'h430ed978, 32'h4369caf2},
  {32'h44f3afea, 32'h40b11311, 32'hc41a7454},
  {32'hc3330986, 32'h433516a7, 32'h438e24fd},
  {32'h44ee0d3c, 32'hc3075925, 32'hc3fd26eb},
  {32'hc3e9c5f0, 32'hc3f5eb2d, 32'h42ef9af8},
  {32'h441e1bbb, 32'hc29865f2, 32'hc3876548},
  {32'hc3448c08, 32'h44118652, 32'h43a2b696},
  {32'h42ab7200, 32'hc01c0e78, 32'h43991d48},
  {32'hc4a33598, 32'h41d9e1b0, 32'hc2c6af60},
  {32'h442b9476, 32'h43754ad7, 32'h4372b918},
  {32'hc4d7ec0b, 32'h43adc928, 32'hc350a08b},
  {32'h440671bc, 32'hc21e4fad, 32'hc2eb137c},
  {32'hc457e7a2, 32'h3fc9f9ce, 32'h428d4d0e},
  {32'h451c09f2, 32'hc2033c34, 32'h437c93e8},
  {32'hc3e49e2c, 32'hc30ed20f, 32'h43c66a1c},
  {32'h44851f9b, 32'hc3b9be7f, 32'hc3018947},
  {32'hc4e74c88, 32'hc30b7e59, 32'h43406d1d},
  {32'h448613c6, 32'h439051bd, 32'h43c96d0e},
  {32'hc42403ca, 32'hc3e0b817, 32'h4323839b},
  {32'h449e84ec, 32'hc2ac8ee6, 32'hc413fe49},
  {32'hc4f5c06c, 32'h42c7d584, 32'h43cc1755},
  {32'h44961a3e, 32'hc3088fb3, 32'h3fa49e20},
  {32'hc349c3f4, 32'hc264d7b0, 32'h42eb0a86},
  {32'h444bb70c, 32'hc14cac33, 32'hc39e4597},
  {32'h4372b9d0, 32'hc29fbc78, 32'hc3bc5fc7},
  {32'hc483b6a7, 32'h428b1815, 32'h432af1a7},
  {32'h44e478fe, 32'hc2149e70, 32'h4329e862},
  {32'hc4c0500d, 32'hc233a736, 32'hc1c3a1d4},
  {32'h44d1572a, 32'hc2f3e8da, 32'hc3907903},
  {32'hc4ca77d5, 32'h433f4277, 32'h43600f9c},
  {32'h43f824e5, 32'hc35fcd2b, 32'h4218f9ff},
  {32'hc482d99f, 32'hc321fee8, 32'hc2c914d9},
  {32'h436f7220, 32'hc3a68080, 32'hc1b14768},
  {32'h42d5f731, 32'h4333bb22, 32'hc42c9412},
  {32'h44864c5c, 32'h435b6df8, 32'hc37b748c},
  {32'hc3389e56, 32'h43495fb6, 32'h4397da81},
  {32'h439dcc0a, 32'h429f5e1e, 32'h434a84cc},
  {32'hc45ee106, 32'hc3834620, 32'hc39c5225},
  {32'h4492cc39, 32'hc376b379, 32'hc2170fda},
  {32'hc4c689b2, 32'hc38c8413, 32'hc1165568},
  {32'h449fef71, 32'hc3358603, 32'hc3daf2b2},
  {32'hc38fee38, 32'h413245ac, 32'hc29e31bb},
  {32'h4507878b, 32'hc2cb4e78, 32'hc330ce7d},
  {32'hc1424080, 32'h4397cc12, 32'hc123fdc6},
  {32'h44e23ee6, 32'h42308220, 32'h42253984},
  {32'hc3f077d0, 32'h4329948e, 32'h42dd14ab},
  {32'h44c24fc4, 32'hc3526117, 32'hc228b62f},
  {32'hc49058f2, 32'hc2d2bdf0, 32'h4304921e},
  {32'h4405320a, 32'hc3d99f9d, 32'hc34c9c12},
  {32'hc3bf986e, 32'hc30dd62b, 32'hc125b77c},
  {32'h441342e7, 32'h43071c81, 32'h4398a57d},
  {32'hc459dc7b, 32'h43e5390a, 32'hc317f0a5},
  {32'h44cb0184, 32'hc28a041e, 32'h43156888},
  {32'hc47f9daa, 32'h40d0048c, 32'h4311ff09},
  {32'h447e5904, 32'h418a9e28, 32'h430044f7},
  {32'hc4f2b75e, 32'hc2c1ab26, 32'hc3dfe885},
  {32'h449305de, 32'hc3f8379f, 32'hc24aa723},
  {32'hc455f620, 32'hc2d5e56d, 32'h42bd0f76},
  {32'h42bfbee2, 32'hc4005f24, 32'hc2e96747},
  {32'hc50d7d8e, 32'hc30d16e1, 32'h42d25275},
  {32'h446a0ad7, 32'hc38b5a6b, 32'hc2ecd18b},
  {32'hc4da661b, 32'hc2de90fe, 32'hc319e83c},
  {32'h43984b64, 32'hc2ab9710, 32'hc15be358},
  {32'hc4a7373a, 32'h42ab5038, 32'hc3d8ee59},
  {32'h4487c541, 32'h43969782, 32'hc2836c5a},
  {32'hc45f5982, 32'h436d3478, 32'hc2ae9da1},
  {32'h45142bc6, 32'hc391c744, 32'hc2d85560},
  {32'hc4f79aaa, 32'hc3886c5a, 32'h42ec5008},
  {32'h44a2b1db, 32'h43c315ca, 32'h4287c962},
  {32'hc4cc113c, 32'hc402a23e, 32'hc304cd94},
  {32'h44925a6b, 32'hc3920e66, 32'hc3813eec},
  {32'hc4dc455e, 32'hc2af3a64, 32'hc27ee1e8},
  {32'h4325a524, 32'hc2251ab3, 32'h438aba6e},
  {32'hc4e84990, 32'hc3687f28, 32'h417d4cfa},
  {32'h45022e81, 32'hc26875ad, 32'h4260ba33},
  {32'hc4a54cfd, 32'hc387df4d, 32'hc31f8763},
  {32'h4508d62d, 32'hc31882de, 32'h43b186ed},
  {32'hc301ee38, 32'hc3b5fd92, 32'hc289a895},
  {32'h44b39aa4, 32'h43b56ef5, 32'hc332d864},
  {32'hc4be7890, 32'hc297af08, 32'hc21e95b2},
  {32'h45000904, 32'hc0094724, 32'hc2e83050},
  {32'hc4b051ec, 32'h434802ab, 32'hc3905568},
  {32'h44b27c60, 32'hc13e86c2, 32'hc36d5711},
  {32'hc4b322a7, 32'hc376427d, 32'hc34403e7},
  {32'h451031f5, 32'hc2ac0c21, 32'h41aa4315},
  {32'hc445769c, 32'h43ae9651, 32'h419f6804},
  {32'h44dda964, 32'h4388d32c, 32'h4283d92f},
  {32'hc4f5e73a, 32'h42fc9853, 32'hc319dc50},
  {32'h43e07af4, 32'h4165aecb, 32'h43894633},
  {32'hc46cbadb, 32'h43bacce6, 32'hc34644d4},
  {32'h43968fa0, 32'h43c572d1, 32'h43158a1c},
  {32'hc50287ea, 32'hc39d607e, 32'hc227f197},
  {32'h450a4053, 32'h43743c9c, 32'h439c1eda},
  {32'hc4f3cc4f, 32'h42ccb593, 32'hc273d3a4},
  {32'h443392c5, 32'h3edbeb6f, 32'h4302288f},
  {32'hc3faab58, 32'h426887ae, 32'h43859899},
  {32'h44032af0, 32'hc386365c, 32'h43c0e91e},
  {32'hc5094c21, 32'hc2a8339f, 32'h4329b9c2},
  {32'h43f73ea8, 32'hc3b6c6d2, 32'h43b6ef33},
  {32'hc4728acd, 32'hc35adcc4, 32'h430c021e},
  {32'h44da398e, 32'h429d5cb3, 32'h43a3d4f5},
  {32'hc4400965, 32'hc316e078, 32'hc34e07d7},
  {32'h449dd8df, 32'h42b9c12d, 32'h4300916a},
  {32'hc4d09b98, 32'hc26fe174, 32'hc299c712},
  {32'h445787fd, 32'hc35e4f63, 32'h4350b906},
  {32'hc5010c6e, 32'hc35e617b, 32'h4318947d},
  {32'h4354ac84, 32'h4375d14e, 32'hc28abefd},
  {32'hc4eaf1e7, 32'hc3bb2430, 32'h42f38672},
  {32'h44a3b382, 32'h430d49c3, 32'h43443d93},
  {32'hc4612214, 32'h43ab5d17, 32'h43405619},
  {32'h43e307a7, 32'h40b89263, 32'h4356ac29},
  {32'hc50498da, 32'h42baa4f2, 32'hc3f27dd9},
  {32'h441b1357, 32'hc14405d1, 32'h43b155a6},
  {32'hc5170c44, 32'hc3d1dffd, 32'h4364b0e7},
  {32'h42bc2270, 32'hc2130b44, 32'h435ece0d},
  {32'hc50d7d5e, 32'hc32978d6, 32'hc32a631f},
  {32'h44018680, 32'h4349ddaf, 32'h4348dc85},
  {32'hc3d4702c, 32'h422533d5, 32'h4245add0},
  {32'h451f3dd8, 32'hc13262c4, 32'hc15cd236},
  {32'hc4ff85cb, 32'hc2e81025, 32'hc35a55a7},
  {32'h4513002a, 32'h4248f75e, 32'h42428790},
  {32'hc4ee1961, 32'h432d51d7, 32'hc3cc5d26},
  {32'h44afeff8, 32'hc18e4191, 32'hc2de380f},
  {32'hc4463eb3, 32'hc387d6dc, 32'h43a9c0c5},
  {32'h44924879, 32'hc37bae64, 32'hc32ba7f9},
  {32'hc4aff65a, 32'h4334e2a7, 32'hc3b2d896},
  {32'h44b5e12a, 32'h439145c0, 32'h41841e6e},
  {32'hc48f0caa, 32'h43052757, 32'hc2841551},
  {32'h44becd9e, 32'h4320ae0c, 32'h4310ff31},
  {32'h432f658b, 32'hc3803c38, 32'h4215f439},
  {32'h44d56dbe, 32'h420a9bb1, 32'hc2a16c86},
  {32'hc323bfd0, 32'h408a1388, 32'hc2af13d3},
  {32'h450623cd, 32'hc37007aa, 32'hc26efd2d},
  {32'hc5022deb, 32'h424caf8c, 32'h42a3f75f},
  {32'h443d7f54, 32'hc224fb92, 32'hc3b21087},
  {32'hc4e8bfc0, 32'hc2408902, 32'h429dff8f},
  {32'h43a96a88, 32'h42ea5ecd, 32'h4218c8e8},
  {32'hc4f4465e, 32'h4180641c, 32'hc3172054},
  {32'h4503a11c, 32'hc28e8a47, 32'hc0f828a0},
  {32'hc28ea970, 32'hc2a48fb0, 32'hc2b97b9e},
  {32'h4513c793, 32'h43660f70, 32'hc2d5d158},
  {32'hc336fd30, 32'hc362972c, 32'hc39c67d6},
  {32'h4444f67e, 32'h434e0236, 32'h4334c643},
  {32'hc420744f, 32'hc316a3eb, 32'hc2e10e03},
  {32'h445721a0, 32'hc3dd6deb, 32'hc3ce8545},
  {32'hc4ac75cf, 32'h40e59b25, 32'h430604ce},
  {32'h43a656c4, 32'hc2faa86e, 32'hc101f690},
  {32'hc4e7a9f4, 32'h43d1268f, 32'hbf313b22},
  {32'h4225aef0, 32'hc1be48e6, 32'hc3d8ee44},
  {32'hc4cd5736, 32'h426807ba, 32'hc3189a3c},
  {32'h439ca40a, 32'hc1375129, 32'hc2b82ce3},
  {32'hc4f457e5, 32'h435ac499, 32'h4284e7ca},
  {32'h43f26a1a, 32'hc3d0e1b0, 32'hc38ef9c6},
  {32'h431127b8, 32'hc29b2802, 32'h4398a74b},
  {32'h44ecaef3, 32'hc3c4d74b, 32'h43bc56c9},
  {32'hc42290d9, 32'hbf1b3abc, 32'hc1d792eb},
  {32'h40677e00, 32'h44129f00, 32'hc38a3ba0},
  {32'hc4e918fb, 32'h440ce50a, 32'hc2284e1c},
  {32'h44c66062, 32'hc21f3df6, 32'h43b23740},
  {32'hc4ced415, 32'hc35cbb4c, 32'hc2824994},
  {32'h44d3b824, 32'h424d8f6a, 32'h43ca17e5},
  {32'hc44dbc32, 32'hc3b1f17c, 32'h43acb357},
  {32'h4495d5a9, 32'hc346247f, 32'hc2f6f3fc},
  {32'hc42a3e6a, 32'h43e7c0c4, 32'hc2902888},
  {32'h45046297, 32'h43b0742d, 32'hc3029a46},
  {32'hc4507900, 32'hc34f80c0, 32'h428a82cb},
  {32'h4471a195, 32'hc2e0bd05, 32'hc2a1bb1c},
  {32'hc4b68659, 32'h43c2102d, 32'hc20abf8e},
  {32'h44906788, 32'h42b9a325, 32'h42ef1686},
  {32'hc4eadb25, 32'hc21a3e89, 32'h4034303c},
  {32'h4502f920, 32'h431318b6, 32'hc29f066a},
  {32'hc4c3b3ba, 32'h43aa4a97, 32'h43a22eee},
  {32'h42b226a0, 32'h43be2888, 32'hc337a2a3},
  {32'hc52d5f35, 32'h43064b62, 32'h436872e5},
  {32'h44ad3ed7, 32'h43883913, 32'h43b28628},
  {32'hc4c15d46, 32'hc398cc1a, 32'h43a018b0},
  {32'h4499a3ae, 32'h429848b0, 32'hc2f7d9dd},
  {32'hc4c1f1cf, 32'hc2d31133, 32'hc39a8079},
  {32'hc37b730c, 32'h4286149e, 32'h43f296ce},
  {32'hc4a2ea3b, 32'h43351426, 32'hc3b8bf91},
  {32'h44f47e95, 32'hc37e4792, 32'hc2cd7f44},
  {32'hc4fd1b47, 32'hc29126ca, 32'hc31b6fb4},
  {32'h43a51943, 32'h42a50519, 32'hc303dba1},
  {32'hc4e8ccd5, 32'hc3a1cfec, 32'h43a1040c},
  {32'h43e5d04e, 32'h41febf02, 32'hc2cdd10f},
  {32'hc455415c, 32'h4373d44d, 32'hc32664d2},
  {32'h44532044, 32'hc217c35f, 32'h434c7ebe},
  {32'hc441b66c, 32'h4319b3e7, 32'hc24c80e3},
  {32'h44af3efe, 32'h432125e7, 32'hc30a0a7a},
  {32'hc4f7864c, 32'h4360d855, 32'hc3b78010},
  {32'h44b18fd5, 32'hc39e7bad, 32'h4400f178},
  {32'hc4c31caf, 32'hc25e40cf, 32'hc34d9b0e},
  {32'h44da883d, 32'hc2e6b55b, 32'h4275c97a},
  {32'hc4a563fd, 32'h4323b1ca, 32'hc3a631f6},
  {32'h44a2cb72, 32'hc273e0d4, 32'hc34d6e3f},
  {32'hc339d286, 32'h43910a3d, 32'h44130ea1},
  {32'h44cc6043, 32'hc3a38979, 32'h42e81d1b},
  {32'hc42c54de, 32'hc2d4ad19, 32'hc2c691b6},
  {32'h446cb1ae, 32'hc1873ea2, 32'hc22dc6a3},
  {32'hc4ab9a80, 32'h429c7091, 32'h43a58423},
  {32'h44917b7e, 32'h42f110f8, 32'hc293b1f2},
  {32'hc50ce1f2, 32'hc366fcac, 32'hc389c1b4},
  {32'h44bb8fd2, 32'hc38d91f9, 32'hc12a47e9},
  {32'hc3b2fc00, 32'hc41a7a0c, 32'hc3d12158},
  {32'h44c51996, 32'hc2fd88a8, 32'h4384ec0b},
  {32'hc3bfb4a5, 32'h43793144, 32'h421b73f2},
  {32'h45050806, 32'hc39a273c, 32'hc11decb3},
  {32'hc4ef3c81, 32'hc418d8dc, 32'hc31e5a35},
  {32'h44ff9f74, 32'hc372eb19, 32'h423d28fb},
  {32'hc4196e38, 32'h42e9e21c, 32'h430a96bc},
  {32'h44ba0ff1, 32'h42d5c43e, 32'hc31225a5},
  {32'hc463d063, 32'h4391e2ba, 32'h43147024},
  {32'h44d25511, 32'h425e1e76, 32'h41c6e84c},
  {32'hc4805eeb, 32'hc35e8ca9, 32'h40863208},
  {32'h44ff3fcb, 32'h4219c783, 32'h413dbfa4},
  {32'hc4fb1eb2, 32'h438d15ed, 32'h42888cee},
  {32'h441161ae, 32'h432afad9, 32'h43506d75},
  {32'hc4a4f167, 32'h42cb3a54, 32'hc3310f36},
  {32'h44dfaad6, 32'hc39d9abf, 32'h42c62428},
  {32'hc4f12c09, 32'hc2f127cc, 32'hc3da7b2a},
  {32'hc2e0cec0, 32'h43c84fc1, 32'h437386ab},
  {32'hc3938234, 32'hc1d3aa50, 32'h43704063},
  {32'h44eb1a36, 32'h42064966, 32'hc3b871d2},
  {32'hc3c5fcbd, 32'h4291653f, 32'h42e580ae},
  {32'h4307e380, 32'hc38ff669, 32'h432430ab},
  {32'hc5098e5d, 32'hc314c4a8, 32'h43a04df1},
  {32'h43ceaa2c, 32'hc3be7d88, 32'hc30369f6},
  {32'hc4ba49aa, 32'hc1aeab48, 32'h432321d4},
  {32'h451d6247, 32'h43848b3d, 32'hc2ad7622},
  {32'hc4f0fa9e, 32'h4363a142, 32'hc2ad73ea},
  {32'h451395b1, 32'h432694a3, 32'hc230895c},
  {32'hc4e95591, 32'h4380f469, 32'hc3d16dd9},
  {32'h44eceadf, 32'hc387b13f, 32'hc3f31e5a},
  {32'hc4dec22c, 32'hc354accb, 32'h4250bf2f},
  {32'h44a61bd2, 32'hc2512712, 32'h43d6ed99},
  {32'hc37938c8, 32'hc2ccac6a, 32'hc1c0dcd2},
  {32'hc25c77f0, 32'hc191ca87, 32'h43aa3440},
  {32'hc31c8cbe, 32'hc3a322c9, 32'h42f91b72},
  {32'h45025076, 32'h43c7fa80, 32'h430bbf28},
  {32'hc4f5fb5f, 32'h421fd4dc, 32'hc320bfa3},
  {32'h4501766a, 32'hc326a78e, 32'hc18340fc},
  {32'hc3a130d8, 32'h423e371f, 32'h437d7f8a},
  {32'h44f2fc9a, 32'h4215c120, 32'h423a8851},
  {32'hc456a199, 32'hc33ba813, 32'h435de20b},
  {32'h431b8a54, 32'hc3a96dc5, 32'h42ef64a4},
  {32'hc42b5a42, 32'hc2c6d39f, 32'h4398826d},
  {32'h44ab21b0, 32'h433781de, 32'h42ffcdc9},
  {32'hc425a638, 32'hc38c006d, 32'h432dbec5},
  {32'h44d68ee3, 32'h43ba5786, 32'hc3881ab4},
  {32'hc3d133c0, 32'hc2ebd9bf, 32'hc3ca650e},
  {32'h44f77712, 32'hbfa07098, 32'hc31d7b54},
  {32'hc45bbd34, 32'hc2977eb3, 32'h4266dc08},
  {32'h45083037, 32'hc396487d, 32'h43b3de3d},
  {32'hc2d26598, 32'hc32e915e, 32'hc2fe8484},
  {32'h44dbc747, 32'h428bf9b6, 32'hc3a6b0cd},
  {32'hc4beace7, 32'hc2b525d4, 32'hc2a817e8},
  {32'h44cca0ec, 32'h4381b3d2, 32'hc1c9c1b2},
  {32'hc288cbeb, 32'h42af4987, 32'h437fd3db},
  {32'h44f427e9, 32'hc2e6d71b, 32'h42df9a33},
  {32'hc4ffd52e, 32'h436b1a03, 32'hc36abe18},
  {32'h445499f9, 32'h43389f62, 32'h4328a290},
  {32'hc45633d2, 32'h4265532d, 32'hc326fad0},
  {32'h449a563e, 32'hc32a4822, 32'h434a9780},
  {32'hc3e2d7e6, 32'h41f6d6c8, 32'h4320f837},
  {32'h4460482a, 32'hc10daf3e, 32'hc2dd0ccc},
  {32'hc48127a6, 32'hbf9f0e82, 32'hc32bc150},
  {32'h451459a4, 32'h4377d4c6, 32'hc29ff6e7},
  {32'hc502c666, 32'h43841de9, 32'hc1a5e8f0},
  {32'h431d61ae, 32'h43c19580, 32'h437ed2b6},
  {32'hc4a8ed0c, 32'hc3ae3184, 32'h4307e970},
  {32'h4497ab38, 32'h417723d5, 32'hc369c8d3},
  {32'hc4b23402, 32'h431e19d1, 32'hc3230243},
  {32'h44f95168, 32'hc22103fa, 32'hc23ab6cc},
  {32'hc5075298, 32'hc2cb201e, 32'hc30751b6},
  {32'h4380d327, 32'hc176a23b, 32'hc2b89c2d},
  {32'hc38f10b8, 32'h4326182b, 32'hc2b44019},
  {32'h45012ec0, 32'hc309997e, 32'h42995861},
  {32'hc3f75127, 32'hc378ecbe, 32'h42c58424},
  {32'h438ea4fc, 32'hc37de10c, 32'hc3334e45},
  {32'hc4c396c3, 32'hc38cbac7, 32'hc3565269},
  {32'h44bebf82, 32'h425dd4d4, 32'hbfebc13c},
  {32'hc3bf8cd8, 32'h43a1b239, 32'hc2439058},
  {32'h43714a68, 32'h431c1bc2, 32'hc390499f},
  {32'hc1eea030, 32'hc2117e58, 32'hc2842860},
  {32'h44097149, 32'hc1e35d1f, 32'h431244c2},
  {32'hc4377470, 32'hc2c37982, 32'hc29f40e1},
  {32'h44fdc6fb, 32'h43a712db, 32'hc3ba2a71},
  {32'hc39fc2d0, 32'hc3693d90, 32'hc19a5c1a},
  {32'h449c9808, 32'h4268c2e8, 32'h42e088cb},
  {32'hc39d1468, 32'hc3407eb9, 32'hc32734f4},
  {32'h4471b3a7, 32'hc19e0171, 32'hc40f931f},
  {32'hc35d3ae0, 32'h44059905, 32'hc3059516},
  {32'h43f446db, 32'h43c3b17b, 32'hc3ead986},
  {32'hc4d5ef5c, 32'hc12054b4, 32'hc21b5675},
  {32'h450f9e52, 32'hc2c8809e, 32'hc38319a2},
  {32'hc38e4d3a, 32'h4390128a, 32'hc23834b6},
  {32'h443e60e8, 32'h431a68ea, 32'hc2c141a3},
  {32'hc42faa50, 32'hc30592e9, 32'hc3a22c3a},
  {32'h451a4e3a, 32'h42647bf6, 32'h4257b45b},
  {32'hc4aa0468, 32'h43309686, 32'hc2fadc9b},
  {32'h44ee9590, 32'h4390db04, 32'h43b32848},
  {32'hc502c3dd, 32'h4235acda, 32'h42d38d93},
  {32'h4512754c, 32'h43cfceda, 32'hc2065964},
  {32'hc4fd00eb, 32'h43bb0f1e, 32'h4196ebb8},
  {32'h432e40f4, 32'h43b34141, 32'h435c6885},
  {32'hc507f897, 32'hc18616f7, 32'h4319a712},
  {32'h43e84f20, 32'h428aabcc, 32'h432720cd},
  {32'hc4b3a872, 32'hc30c399d, 32'h4323eb46},
  {32'h44ac7478, 32'h41788626, 32'h4332ff47},
  {32'hc4311610, 32'hc385a0cc, 32'h42f53549},
  {32'h44e6ef2f, 32'h42dc6641, 32'hc3ed8111},
  {32'hc4f59dae, 32'hc33ab5f2, 32'h428d2aae},
  {32'h444539e4, 32'hc4000f17, 32'h43c4665d},
  {32'hc45b71ad, 32'h42106178, 32'hc34ce45a},
  {32'h44d2a357, 32'h431d708f, 32'hc3712de4},
  {32'hc46dbfaf, 32'h42163f67, 32'h42f3ab07},
  {32'h435b7276, 32'hc397e682, 32'hc3b4a140},
  {32'hc4ca7f41, 32'hc3f1391a, 32'hc372c1c9},
  {32'h4516748e, 32'hc1a22792, 32'h416e3054},
  {32'hc4c5e8de, 32'h41efdf1d, 32'hc2963961},
  {32'h4402fefe, 32'h4356f865, 32'h43db24c5},
  {32'hc31f4d94, 32'h435a4c4f, 32'hc3424694},
  {32'h44b6b550, 32'hc343b282, 32'h430a2c3c},
  {32'hc4846831, 32'h413a1b7a, 32'h4385e1e5},
  {32'h44b09b48, 32'h439be28b, 32'hc2f77dbc},
  {32'hc4d434c6, 32'h40febda0, 32'h4335ae73},
  {32'h4438f450, 32'h42ac09b7, 32'h432e05ba},
  {32'hc4ed572b, 32'h436b594c, 32'h42d80640},
  {32'h4384ed24, 32'hc31d8ec9, 32'hc29f43a3},
  {32'hc4a49a07, 32'hc30554c4, 32'h434642a0},
  {32'h44e1b484, 32'hc327c7e6, 32'hc350e7d7},
  {32'hc42dc695, 32'hc2a274ce, 32'hc237050b},
  {32'h45083f6f, 32'hc2427f10, 32'h441acd6f},
  {32'hc41b99c2, 32'hc20d26f6, 32'h4229cd0e},
  {32'h447e1e0a, 32'hc28104a6, 32'hc2998a09},
  {32'hc47b17b8, 32'h418461fd, 32'hc2ad1001},
  {32'h44be3fd3, 32'h4371f684, 32'hc21936a8},
  {32'hc34eb142, 32'h439687e9, 32'h4283937b},
  {32'h42b0ffcb, 32'hc32250c4, 32'h4306982c},
  {32'hc4dfd29f, 32'h4296b724, 32'hc38d7d58},
  {32'h449281e5, 32'hc3729fd2, 32'hc3d8deda},
  {32'hc4f601da, 32'hc36b03f0, 32'hc2acf95a},
  {32'h4510869c, 32'hc3a282df, 32'h42b68319},
  {32'hc49f01e6, 32'hc1af990f, 32'hc3d73ec7},
  {32'h44e6da8c, 32'h4269368f, 32'h41df2559},
  {32'hc4893407, 32'hc289f151, 32'hc2db07de},
  {32'h449bf7b2, 32'h41d1b2d5, 32'hc2210fa6},
  {32'hc4d6d537, 32'hc20aabd6, 32'hc16503ec},
  {32'h44aafa3a, 32'hc3b849cd, 32'h43d9bd35},
  {32'hc4ce0e5b, 32'hc2a6a3c2, 32'h4213d44b},
  {32'h44e45135, 32'hc2973f58, 32'hc2e6b490},
  {32'hc4906f42, 32'h43aea9cb, 32'h437d04bf},
  {32'h42c0b380, 32'hc29c6337, 32'h425b4600},
  {32'hc47d77ca, 32'h43a2bfe6, 32'h42a0815c},
  {32'h44cd2532, 32'hc2ec8622, 32'h4346a777},
  {32'hc44c1e6b, 32'h42cf4f0f, 32'h42fe7cd8},
  {32'h44f34b46, 32'h41581242, 32'hc392ee6e},
  {32'hc51ba68c, 32'h41dbac09, 32'h439447b3},
  {32'h43d1c1d9, 32'h42730180, 32'h43789c7b},
  {32'hc4edfe71, 32'hc3c849bb, 32'hc3a3363f},
  {32'h42a2f240, 32'hc2afeb21, 32'hc3154c0e},
  {32'hc4811947, 32'h43b6afd3, 32'hc34093e6},
  {32'h4514eafd, 32'h40684594, 32'h42632355},
  {32'hc4456822, 32'h4379ac1e, 32'hc368bf3c},
  {32'h4516ed19, 32'h423d138e, 32'hc261830a},
  {32'hc3a58f0e, 32'hc305e668, 32'hc3a99aa4},
  {32'h4409f2a6, 32'h42953b9b, 32'hc382a701},
  {32'hc49f88b5, 32'hc3093cda, 32'h41bfe58c},
  {32'h447ca524, 32'hc287fd1d, 32'hc2b28532},
  {32'hc5125026, 32'h4411d004, 32'hc3b21bf7},
  {32'h448a1df4, 32'h420d77c1, 32'h43a3dce0},
  {32'hc5188018, 32'hc12ef7e7, 32'h4229fb97},
  {32'h44679853, 32'hc1648875, 32'hc220957e},
  {32'hc5149462, 32'hc281947e, 32'h43fdd6d3},
  {32'h4346b9da, 32'hc1b12bad, 32'h42859db7},
  {32'hc5007aae, 32'hc391fb6a, 32'h438c0121},
  {32'h4509e776, 32'hc2af921b, 32'h4302aa96},
  {32'hc4940a2e, 32'hc25eb77c, 32'h438a9d6b},
  {32'h44e5d119, 32'hc2457b1b, 32'hc1fc6e2d},
  {32'hc51371fa, 32'h432faf2c, 32'hc1324f40},
  {32'h44b62e74, 32'hc27039c1, 32'hc3845c42},
  {32'hc4851d69, 32'h41a844a8, 32'h41b7f564},
  {32'h4512643e, 32'h42bd49c2, 32'hc345ae22},
  {32'hc518fab7, 32'hc32e68a2, 32'h43794bbf},
  {32'h44f62b0d, 32'hc3e5e895, 32'hc3988c99},
  {32'hc4e7a495, 32'hc2523f7d, 32'h42e34d39},
  {32'h4504d09c, 32'h4342e076, 32'h42680526},
  {32'hc3c7f828, 32'h4351c38c, 32'h42eb7418},
  {32'h44cce22b, 32'hc36d4dca, 32'h41a63667},
  {32'hc4ee3f1f, 32'h43852c7d, 32'hc2b08099},
  {32'h44400ff0, 32'h43186d7a, 32'hc2ae42c4},
  {32'hc31666c0, 32'h41912716, 32'hc3e8c8bc},
  {32'h44975c68, 32'hc1a38d04, 32'h43616f8f},
  {32'hc375dfa8, 32'hc27d96b8, 32'h41f1fdd0},
  {32'h451a69c5, 32'h4358e8b5, 32'hc3ede044},
  {32'hc36f7f10, 32'h435deafe, 32'h4390085d},
  {32'h440a6420, 32'h41038518, 32'h434415d0},
  {32'hc3e895fa, 32'hc2dd5a26, 32'h421ffbb9},
  {32'h44679e99, 32'h4343d370, 32'hc2ee94d6},
  {32'hc50c60c8, 32'hc3a54e53, 32'h43d1cf9f},
  {32'h4499de7e, 32'h436ac631, 32'h41f58d93},
  {32'hc47374ac, 32'h4333b780, 32'h41e10055},
  {32'h440a9134, 32'h43597e41, 32'h4391a897},
  {32'hc50c805e, 32'hc3823082, 32'hc2dd4ce3},
  {32'h45155403, 32'hc32bd676, 32'hc1e89857},
  {32'hc4d877b0, 32'hc2c03325, 32'h4216af3b},
  {32'h441c7544, 32'hc3c66b57, 32'h41d126d3},
  {32'hc42f161c, 32'h43435564, 32'h43977c01},
  {32'h435bf10c, 32'hc2081ec6, 32'h4389e8b1},
  {32'hc42abe66, 32'hc2250a74, 32'hc35aeb6b},
  {32'h44b9503b, 32'hc341f5b2, 32'hc283b258},
  {32'hc49e7386, 32'hc3b28fc6, 32'h42d40c80},
  {32'h44eab7a2, 32'h42406510, 32'hc364b01f},
  {32'hc4972e25, 32'hc2b09726, 32'h421c6f97},
  {32'h4507f734, 32'h433cc809, 32'hc292f56f},
  {32'hc4c0488c, 32'h42063e61, 32'h43481b0d},
  {32'h43f6febc, 32'h42684248, 32'hc288a22c},
  {32'hc4c3fd6d, 32'hc3ae9510, 32'h43ad18fc},
  {32'h44eb39e3, 32'h42ac0cb1, 32'hc2d230fb},
  {32'hc5199ce0, 32'hc333766e, 32'hc3dc8008},
  {32'h442c0552, 32'hc202a804, 32'hc336d501},
  {32'hc3e38547, 32'hc30c2538, 32'hc34b6d79},
  {32'h43943328, 32'hc380952d, 32'hc34cda97},
  {32'hc400cfd0, 32'h42886206, 32'h4293405f},
  {32'h446e861b, 32'hc211a150, 32'h4254b6d8},
  {32'hc4430da6, 32'h43811e6a, 32'hc3a0d227},
  {32'h44fedfda, 32'h43ecd352, 32'h42792b57},
  {32'hc49a0c09, 32'h43b6dca6, 32'hc3878d34},
  {32'h44b974ba, 32'hc34b7cbf, 32'hc349ccbc},
  {32'hc3eb083c, 32'hc32e7239, 32'hc36ad609},
  {32'h450ff471, 32'hc3100612, 32'h43712d64},
  {32'hc3a331d8, 32'hc36c3bd0, 32'hc2b9e70f},
  {32'h441c2348, 32'h40aa0f78, 32'h43d0c3c9},
  {32'hc403fac8, 32'h42915cbb, 32'h42548d8a},
  {32'h44400830, 32'h439a6b51, 32'h43b6e94e},
  {32'hc4d7df28, 32'hc228052d, 32'h4311a178},
  {32'h44f10b25, 32'hc33f709f, 32'h436cf244},
  {32'hc4ddc261, 32'h42a451d5, 32'h42cdcbf2},
  {32'h448c37f4, 32'h426eb886, 32'h42994ba7},
  {32'hc46c8b9a, 32'h4291a575, 32'hc2c76083},
  {32'h44dc90f1, 32'h43374f69, 32'h436e3f35},
  {32'hc493bb96, 32'h4196a798, 32'h42bd0aec},
  {32'h44861db8, 32'h4374fe8e, 32'h43cf8bd7},
  {32'hc484b5b5, 32'hc3377893, 32'hc41575ca},
  {32'h450859d5, 32'hc39e315d, 32'h40b3b400},
  {32'hc170f7b0, 32'h431baf41, 32'hc20c5902},
  {32'h44317612, 32'h43902d07, 32'h42119e48},
  {32'hc50fc81e, 32'hc0ed949f, 32'hc2cd2fbe},
  {32'h44e2bbf4, 32'h42743fae, 32'h43f5f95f},
  {32'hc4a4f2c0, 32'hc20b288c, 32'hc38f4bf4},
  {32'h44873705, 32'hc3292d96, 32'h439fee10},
  {32'hc4818fc9, 32'h42ea7f8a, 32'h416c3ee1},
  {32'h44679172, 32'h4387800d, 32'hc386792f},
  {32'h41b856e0, 32'hc3d226e3, 32'hc3093c83},
  {32'h4512469f, 32'h42a8fd54, 32'hc3600b70},
  {32'hc3fc5b3c, 32'h42e14551, 32'hc206587f},
  {32'hc50ef182, 32'hc1e9009c, 32'h4341cfbc},
  {32'h441f1c16, 32'hc21148a8, 32'hc33ea9ee},
  {32'hc4caa436, 32'h431a0123, 32'hc32488c0},
  {32'h44d06859, 32'hc41d0b93, 32'h43bafef1},
  {32'h4314f278, 32'h438b0b6e, 32'hc1ea2b76},
  {32'h444c1ac2, 32'hc3877f7c, 32'hc29aecc1},
  {32'hc3a41f98, 32'h430fe1fa, 32'hc3ba0ecf},
  {32'h423d4ac0, 32'h43c77380, 32'hc38c3cb3},
  {32'hc4844bee, 32'h43a895ac, 32'hc300b9d4},
  {32'h43815eb6, 32'h43b331cd, 32'h41949bce},
  {32'hc3418740, 32'h432eba65, 32'hc391307c},
  {32'h444c923c, 32'hc216198c, 32'h43a63b90},
  {32'h42c10ad4, 32'h43eccb29, 32'h42f7f1b8},
  {32'h44a12a85, 32'h4307ca58, 32'hc39fea3e},
  {32'hc2bf3e10, 32'hc3526337, 32'hc402ca0e},
  {32'h4421b9a8, 32'hc29c5c0a, 32'h431ebf2f},
  {32'hc4b305c8, 32'h431ffefd, 32'h425021d2},
  {32'h44b1c81b, 32'h4295f877, 32'h42e0a9bb},
  {32'hc4622976, 32'hc3db4d52, 32'hc3a7d9ad},
  {32'h4450354d, 32'h4347cc0a, 32'h43ddc76c},
  {32'hc4c142da, 32'h4389236c, 32'hc3a06bbd},
  {32'h4508c4f3, 32'h428e6d31, 32'hc2bad442},
  {32'hc39ac3a8, 32'h4210c79e, 32'h42053657},
  {32'h44928d98, 32'h4288baa9, 32'h42649cde},
  {32'hc4b96106, 32'hc286cf32, 32'h43297758},
  {32'h447d8f12, 32'h4366c932, 32'h43664416},
  {32'hc51437fe, 32'h4205b418, 32'h4347a17e},
  {32'h451d379c, 32'hc39f6410, 32'hc2a44215},
  {32'hc3afde44, 32'h43aee58d, 32'hc3c30626},
  {32'h450a5daf, 32'hc3632e03, 32'hc1ab7a2b},
  {32'hc4475382, 32'hc264fe58, 32'h42ee6757},
  {32'h44d984f8, 32'hc3270932, 32'h43246847},
  {32'hc4df96b3, 32'hc2d66633, 32'h435b4c24},
  {32'h4475f86a, 32'hc249016f, 32'hc24a2063},
  {32'hc4a9e1dc, 32'h43ffd3e8, 32'h4285baa3},
  {32'h44dfa9bd, 32'hc30b0891, 32'h4214f80d},
  {32'hc45b3562, 32'h433fde1a, 32'hc32b8431},
  {32'h447e000b, 32'hc2603b81, 32'h433ab853},
  {32'hc3ead98c, 32'hc2837c08, 32'hc2c86b2e},
  {32'h42fcef2c, 32'h4322177c, 32'hc301da0f},
  {32'hc22ddd30, 32'h418b62ef, 32'h428ae0c4},
  {32'h4508d349, 32'hc398539a, 32'hc320024d},
  {32'hc4759df4, 32'h4380e049, 32'h43412c2c},
  {32'h45033279, 32'hc3cdee07, 32'hc36ffa4a},
  {32'hc3b82744, 32'hc10f5f3c, 32'h437c8114},
  {32'h443c82b8, 32'hc26fa82b, 32'hc381d6dd},
  {32'hc412b24c, 32'hc2bc79f7, 32'h42df8bbc},
  {32'h43e19938, 32'h41706ba2, 32'h42ffde97},
  {32'h42bd1dfd, 32'h4318e254, 32'h427712d9},
  {32'h450ca934, 32'h437f3e01, 32'h4309e22b},
  {32'hc4df830c, 32'hc2f1b826, 32'hc19cfe67},
  {32'h442b9d12, 32'hc19d4192, 32'h4351f702},
  {32'hc418fcf8, 32'h43ca6102, 32'hc30f3742},
  {32'h44e25ed9, 32'hc32d41a2, 32'h434dd176},
  {32'h406ccc00, 32'hc2f8bec3, 32'hc31ddc1b},
  {32'h4379de38, 32'hc34c8add, 32'h42219cc4},
  {32'hc43dea36, 32'h42686acc, 32'hc322d79a},
  {32'h43c2775c, 32'h43a23a68, 32'h42bc356c},
  {32'hc4e7e2d3, 32'h428cd53a, 32'hc355820e},
  {32'h44c35a65, 32'h4333f3cc, 32'hc35a40f6},
  {32'hc46e42fe, 32'h43820216, 32'hc2eaef56},
  {32'h449b6f86, 32'h41ffd890, 32'h435a5f9a},
  {32'hc50f2020, 32'hc38dd0ac, 32'hc356e100},
  {32'h4494133e, 32'hc383a29a, 32'h437fbd78},
  {32'hc4b5ee72, 32'hc30ef426, 32'hc37d0286},
  {32'h449e1d16, 32'h43560af8, 32'h4427b0d3},
  {32'hc29100e0, 32'hc304890f, 32'hc315f5e6},
  {32'hc2ae7eaa, 32'hc10497a3, 32'hc3a7dddc},
  {32'h438b51ed, 32'h43fbdb92, 32'h423505d8},
  {32'h44dae2aa, 32'hc1c43ec8, 32'h42b01226},
  {32'hc506292a, 32'h433c3f4a, 32'h423d2a11},
  {32'h42ef4490, 32'hc39b2667, 32'h43121a85},
  {32'hc4f514eb, 32'h4338abf1, 32'hc3f78328},
  {32'h445a78aa, 32'h42f2bc1e, 32'h4213fc89},
  {32'hc441e1f0, 32'hc317c416, 32'hc241d6cc},
  {32'h44fba60a, 32'h43c8324a, 32'h41ed9e0b},
  {32'hc3b92008, 32'hc380dfaa, 32'hc30bdd66},
  {32'hc2db0cd0, 32'hc2f199b0, 32'h421400f5},
  {32'h4382c567, 32'h4391525c, 32'h430afbc6},
  {32'h44d45c9b, 32'hc37693e2, 32'h4407e92a},
  {32'hc50e72bb, 32'h40ac353a, 32'h42d8d69a},
  {32'h44b48c39, 32'h4140e473, 32'hc327ba80},
  {32'hc4f589af, 32'h43240fd4, 32'hc35bbca3},
  {32'h4481e4b1, 32'hc2ad310f, 32'hc41037c3},
  {32'hc4c00803, 32'h43831125, 32'h421a22e8},
  {32'h44b104be, 32'h42b995ad, 32'hc262713e},
  {32'hc4a60ac3, 32'h429d8f37, 32'h425b48d4},
  {32'h4396cff0, 32'h4384febf, 32'h42da7b9c},
  {32'hc4607c4c, 32'hc2a2a284, 32'hc321e87d},
  {32'h45098e18, 32'h4394ec91, 32'hc3e32f45},
  {32'hc4e439f5, 32'h434cd887, 32'h428f23ce},
  {32'h44b6f396, 32'h40fa35ce, 32'hc3164516},
  {32'hc2ed694a, 32'hc3b32b5f, 32'hc328633e},
  {32'h44e8e38a, 32'h431c7516, 32'h43aaca94},
  {32'hc4e3c028, 32'h415fe5d3, 32'h433c8131},
  {32'h44d81bb3, 32'hc29189d6, 32'hc2cc5a1e},
  {32'hc50a5210, 32'h436e13c9, 32'hc281d700},
  {32'h4514c3a6, 32'h42fdff49, 32'hc26075db},
  {32'hc3a9dd5e, 32'hc2fbd4b2, 32'hc2703102},
  {32'h44dd3cc1, 32'hc379b626, 32'hc261f22e},
  {32'h42e59c26, 32'hc3277e2a, 32'h4361cc7d},
  {32'h4466a522, 32'h43d9f070, 32'hc340e5d0},
  {32'hc4d746ae, 32'hc287ff37, 32'h42fb2303},
  {32'h44f270e4, 32'hc38d6807, 32'h43820116},
  {32'h43286ab4, 32'h4404a4da, 32'h4289d4af},
  {32'h45089f08, 32'h438ed002, 32'h42f2104f},
  {32'hc4e66ad8, 32'h430df8ff, 32'hc3aac6d5},
  {32'h4441ca32, 32'hc4072aa9, 32'hc288ebc4},
  {32'hc50341a0, 32'h41516ed2, 32'h43ac534e},
  {32'h44d6f8dd, 32'h43e08e7c, 32'hc38c579f},
  {32'hc4dc7502, 32'h43d9055c, 32'h420f4afa},
  {32'h451ccfe2, 32'h43bfe773, 32'h4250afdb},
  {32'hc4a647fb, 32'hc285f19e, 32'hc2976b68},
  {32'hc1525bc0, 32'h42c6cdea, 32'hc2994e3c},
  {32'hc504ada5, 32'h438d2673, 32'h4293b10c},
  {32'h451308a5, 32'hc291a9f2, 32'hc3c7f747},
  {32'hc4ff005e, 32'h4336edca, 32'h43973c39},
  {32'h44a6f915, 32'h43159d7a, 32'hc31473ab},
  {32'hc3d9188a, 32'hc2f91696, 32'hc2962f0d},
  {32'h44df7eb8, 32'h430b8466, 32'hc195fc98},
  {32'hc3a8e20c, 32'hc30ed096, 32'h42d8824c},
  {32'h44cf9dcb, 32'h431f0aa5, 32'hc38e086d},
  {32'hc4fb432f, 32'h41a4d646, 32'h42973885},
  {32'h44b69d45, 32'hc2e4b4cc, 32'hc2f0d1a7},
  {32'hc403c8aa, 32'hc30f10cc, 32'h43473bc1},
  {32'h4387934c, 32'hc346b74b, 32'h43a92b09},
  {32'hc3e747ab, 32'h43816da2, 32'h42b0860a},
  {32'h43a0af70, 32'hc35de903, 32'h42e18f51},
  {32'hc4a24603, 32'hc3af9fe1, 32'hc25ee6b6},
  {32'h44bf8140, 32'h432cf885, 32'hc1a653cc},
  {32'hc43b60bb, 32'hc30af5e1, 32'hc34add41},
  {32'h42b83ed0, 32'hc1d63759, 32'h43d6f48d},
  {32'hc3f0e916, 32'hc2f72fce, 32'h4278e531},
  {32'h44b38c02, 32'hc3542849, 32'h43a5792c},
  {32'hc41bb2c6, 32'h4295853e, 32'h3f0861b8},
  {32'h44df1bb4, 32'h43bc5d8e, 32'h42e5e395},
  {32'hc4a70a0a, 32'hc32c0536, 32'h434d98da},
  {32'h44864fa8, 32'h43734c5c, 32'h4290211f},
  {32'hc450368c, 32'h436b1964, 32'hc30bdb9b},
  {32'h45037556, 32'hc38ae129, 32'hc386d9ea},
  {32'hc48770ee, 32'h434ffd13, 32'h424ccbc8},
  {32'h44fb010e, 32'h423662c9, 32'hc3c68900},
  {32'hc4ddac6c, 32'h425c7b03, 32'h441c83ea},
  {32'h442d2d5d, 32'hc319e622, 32'hc24f554d},
  {32'h408181e0, 32'h43981f1c, 32'h43b8e924},
  {32'h44e349ea, 32'h43ad96dd, 32'hc400950a},
  {32'hc397b0f5, 32'hc3003f00, 32'h42e2ea36},
  {32'h45073ad3, 32'h43a7301e, 32'hc3777812},
  {32'hc45f3e0c, 32'h43bc8225, 32'hc388c4b7},
  {32'h44bc2486, 32'h43e72bf4, 32'hc36e8092},
  {32'hc46acf92, 32'h4314ae39, 32'hbfe246f8},
  {32'h45060f56, 32'hc336f527, 32'hc3c2878b},
  {32'hc495210a, 32'hc2f292ec, 32'hc265b07a},
  {32'h440603cc, 32'hc338d00a, 32'hc27ffb0b},
  {32'hc4bb17ff, 32'h42bc6981, 32'h42d0d1d8},
  {32'h448905e4, 32'hc2f85eeb, 32'hc18f29c4},
  {32'hc4e5ec61, 32'hc29f05b8, 32'h4316fa53},
  {32'h44bb2973, 32'h4259132d, 32'h4327e4ab},
  {32'hc506da24, 32'h431162ae, 32'hc33cf1eb},
  {32'h447badbe, 32'hc38b7ed0, 32'h43aeb9fd},
  {32'hc4b36a60, 32'h43641358, 32'h41c2de7d},
  {32'h4406814c, 32'h4171f27c, 32'h4197c67b},
  {32'hc5144f7d, 32'hc279369e, 32'hc2e10f5d},
  {32'h4494ca3e, 32'h434528fa, 32'h438311e3},
  {32'hc37126f0, 32'h41aedf66, 32'h42e2ed41},
  {32'h43378fe0, 32'h4348f802, 32'hc3141cbe},
  {32'hc4cb19dc, 32'hc30ddbf7, 32'h433eba7e},
  {32'h42d2dc84, 32'h42cf7a88, 32'hc33a7b9f},
  {32'hc2bc62e2, 32'h437d63ae, 32'hc1fe6a5e},
  {32'h449d4af0, 32'hc326af7c, 32'h438ea902},
  {32'hc4285717, 32'h4344996a, 32'h42ea9782},
  {32'h44597962, 32'hc209bb80, 32'hc33294b4},
  {32'hc4fee734, 32'h42b7cf24, 32'hc265040a},
  {32'h44c831b2, 32'h428cb9d1, 32'hc366e60c},
  {32'hc4f2b555, 32'h40d1b8b0, 32'hc25c2245},
  {32'h44fbfae7, 32'hc2adb545, 32'h42b0a782},
  {32'hc49d97a9, 32'hc24ca5c6, 32'hc3dde834},
  {32'h44c25de2, 32'h41410042, 32'hc22855f2},
  {32'hc4edd3c1, 32'hc3275c95, 32'hc33bea95},
  {32'h4473a101, 32'hc393d907, 32'h4364e67f},
  {32'hc502acb0, 32'h438816a9, 32'h42f32310},
  {32'h445c5b2f, 32'hc3524469, 32'hc2a073b1},
  {32'hc507f632, 32'hc328cc3d, 32'hc21dd256},
  {32'h44a9c6ce, 32'h4373eca8, 32'hc34aff0e},
  {32'hc50ab468, 32'hc3853935, 32'hc30d0894},
  {32'h446a5905, 32'h42a45e86, 32'h44050ab7},
  {32'hc42c9a86, 32'hc1c5fb3f, 32'h42a0e7e7},
  {32'h441392ac, 32'h43061a9e, 32'h4340cbbd},
  {32'hc503ae18, 32'hc25d2532, 32'hc1adff80},
  {32'h44ba1878, 32'h438461bb, 32'hc308e00d},
  {32'hc45849ce, 32'hc25ce41b, 32'h41535219},
  {32'h451c276c, 32'hc2658170, 32'h40aea81c},
  {32'hc4ba80e8, 32'h423f97a9, 32'h436de2cd},
  {32'h44ae9230, 32'hc2876c6a, 32'h42f59197},
  {32'hc29a3ee0, 32'h439989fe, 32'hc29e6a51},
  {32'h43bca630, 32'hc2edb0bc, 32'hc24e999e},
  {32'hc356a360, 32'h4212a702, 32'h4365303d},
  {32'h416a0580, 32'hc386c6d6, 32'hc2e98a23},
  {32'hc44e6558, 32'hc1946582, 32'h420f09c1},
  {32'h44d8778e, 32'hc25c71f5, 32'h42b283b6},
  {32'hc50ca6d9, 32'h42b8a2b3, 32'hc3926a2a},
  {32'h44bd6e78, 32'h41201fcc, 32'h439e88ee},
  {32'hc4bb8c66, 32'hc39edd46, 32'h43202242},
  {32'h44d958a3, 32'h422e7448, 32'hc117b345},
  {32'hc4bf9301, 32'hc38a2b77, 32'hc331cdab},
  {32'h44ccdc4e, 32'h4387f058, 32'h4315cf52},
  {32'hc432d276, 32'hc31289f3, 32'h42c404ab},
  {32'h448091c3, 32'h430211db, 32'hc36fb43a},
  {32'hc435ce50, 32'h436bbf9c, 32'hc3a6b7f4},
  {32'h43c91dc2, 32'hc1e9c4ea, 32'h426b0e1a},
  {32'hc4143c52, 32'h43d1de2a, 32'h43c21b8f},
  {32'h450ee7e1, 32'hc2f5636b, 32'hc39935cb},
  {32'hc4ab580b, 32'hc186483e, 32'h42893f92},
  {32'h44981544, 32'hc41b5d8b, 32'h41bc2d92},
  {32'hc4fdfa0e, 32'hc3084eaa, 32'h42d829fb},
  {32'h43f2a9b2, 32'hc3b7f552, 32'h41b89bde},
  {32'hc39c0205, 32'hc3ce5469, 32'h4259033c},
  {32'h44bcd567, 32'hbf01c989, 32'h43c79252},
  {32'hc4abd0f2, 32'h41275814, 32'hc3ab1b74},
  {32'h44ae7073, 32'h431df31c, 32'h4245949d},
  {32'hc43b615d, 32'h428857c8, 32'hc36b80aa},
  {32'h44807cb6, 32'hc0297f35, 32'h434b5088},
  {32'hc485baac, 32'hc233bb74, 32'hc3b2c253},
  {32'h45014404, 32'h42df9746, 32'hc35f475b},
  {32'hc4cbb023, 32'hc154a494, 32'hc16684f4},
  {32'h416f7e00, 32'h4262a62a, 32'h437888be},
  {32'hc4c7992b, 32'h4381bf17, 32'hc2e748bf},
  {32'h44e5e592, 32'hc2cea3c6, 32'h40354f1c},
  {32'hc4d1c3fd, 32'h43928e13, 32'h431e9c3d},
  {32'h440fae18, 32'h42fdd8a2, 32'hc1ffaaf4},
  {32'hc4dead2e, 32'h43739a8d, 32'h4293f3fc},
  {32'h44c86c11, 32'hc26bd7ee, 32'h42257a37},
  {32'hc4564af1, 32'hc26fb5dc, 32'h43c3dfc6},
  {32'h43a6e168, 32'hc30aec3b, 32'hc0cfa992},
  {32'hc4eb072a, 32'hc349ad47, 32'hc3a0cb6a},
  {32'h45134cc1, 32'hc37a1838, 32'h42c58974},
  {32'hc46d2c34, 32'hc3a630cb, 32'h431ad30f},
  {32'h43aeb200, 32'hc298e22a, 32'h43312bf2},
  {32'hc4f3da68, 32'hc417b398, 32'hc3b35abc},
  {32'h4434de27, 32'hc374a089, 32'hc1350300},
  {32'hc38d5a80, 32'h43f03ca5, 32'hc2fbe89d},
  {32'h44816666, 32'h43aaf973, 32'hc33945ca},
  {32'hc380e320, 32'h42e97912, 32'hc39326c5},
  {32'h4514aaef, 32'h42a8b29c, 32'hc38047d4},
  {32'hc4d34dbd, 32'h43544b63, 32'h44299e94},
  {32'h442719a9, 32'h42bd3655, 32'hc2a438c9},
  {32'hc47434d8, 32'h436a7d8f, 32'hc20d860a},
  {32'h43a775f8, 32'hc3b64abf, 32'h43204dce},
  {32'hc3750c19, 32'hc2e23c7e, 32'hc3dd7101},
  {32'h44f0e602, 32'hc26518e2, 32'hc3a392f3},
  {32'hc3a25ce4, 32'hc2c948cd, 32'hc370e043},
  {32'h44f45ffa, 32'hc28217ee, 32'h4299e11c},
  {32'hc4270961, 32'hc27096f9, 32'h433ea2e5},
  {32'h441dc90e, 32'hc0fe0ae0, 32'hc3a0ab72},
  {32'hc4d754b6, 32'h433582b0, 32'hc306649a},
  {32'h4488aefe, 32'hc2b538bc, 32'hc390aac5},
  {32'hc4fbc3a7, 32'h4311db8e, 32'h42de9463},
  {32'h4500dae4, 32'h4223d4df, 32'hc2c649ae},
  {32'hc21e6ca0, 32'h43ae4773, 32'h42eee19d},
  {32'h44d3f104, 32'h424f49a6, 32'h441cd24c},
  {32'h431581d8, 32'hc217cb5a, 32'hc32a580e},
  {32'h44b6d244, 32'hc389daf0, 32'hc2e3d139},
  {32'hc41ddec0, 32'h41e62a81, 32'h42943346},
  {32'h44d2d69e, 32'h43945d49, 32'hc38073f6},
  {32'hc4c15d02, 32'hc1d1f322, 32'h42156546},
  {32'h442bc888, 32'hc15b84b6, 32'h439543b4},
  {32'hc409e97b, 32'hc1a896cc, 32'hc3677d27},
  {32'h4511acdc, 32'h430cd738, 32'hc339cc1e},
  {32'hc47ef07b, 32'h43e357f4, 32'hc3cd62c1},
  {32'h450ed691, 32'hc3abace1, 32'hc37f013b},
  {32'hc36f5804, 32'hc3385565, 32'h4304e033},
  {32'h44c3c8d2, 32'hc3203486, 32'h435253e9},
  {32'hc4d26e92, 32'hc3a8462b, 32'h431683b1},
  {32'h4415dbe2, 32'h4307efb0, 32'h429dcf2b},
  {32'hc47bef16, 32'hc332aa14, 32'h4308c04d},
  {32'h451e9879, 32'hc325f58d, 32'hc325ef22},
  {32'hc51604b1, 32'h430111ff, 32'h43a5598f},
  {32'h44bcaa6a, 32'h4304b488, 32'h4365d5f7},
  {32'hc513a21b, 32'h4384bf8d, 32'h4250ebb0},
  {32'h4500c0f2, 32'hc3572fdd, 32'h40d2af69},
  {32'hc4ce4be8, 32'h42be5b4c, 32'h43cc8fdd},
  {32'h44e84a64, 32'h427bd3ff, 32'h433a3fb2},
  {32'hc39350d8, 32'h421005c8, 32'h4349c897},
  {32'h4416219e, 32'hc2552688, 32'h428f0828},
  {32'hc488ba01, 32'h41072cce, 32'h429d2fc2},
  {32'h43e8f398, 32'hc3510f72, 32'h43c01181},
  {32'hc5020797, 32'h42925f79, 32'h435e1454},
  {32'h45168896, 32'hc329a826, 32'h41761994},
  {32'hc4f5f352, 32'hc3677b7f, 32'h41003a38},
  {32'h44017b4c, 32'h4400b1cf, 32'h4310026e},
  {32'hc48de4e0, 32'hc298a8e5, 32'hc3c52292},
  {32'h45032a20, 32'hc3287ac7, 32'h43859b4a},
  {32'hc4c2ce54, 32'hc2d36c29, 32'h42d6b092},
  {32'h4501293d, 32'hc28eaa38, 32'hc27f9b16},
  {32'hc506f621, 32'hc31d0c7b, 32'hc2cae0db},
  {32'h4494c4be, 32'hc20a4376, 32'hc3bf16c3},
  {32'h41af2aea, 32'h42ce167f, 32'h4383f164},
  {32'h44891cf8, 32'hc2c6ec0c, 32'hc2a12277},
  {32'hc4b27258, 32'h43a18100, 32'h436d4a4a},
  {32'h44e47576, 32'h42502aca, 32'h43a3cfa2},
  {32'h430f1ba0, 32'hc33505fa, 32'hc384bfac},
  {32'h4480a284, 32'hc34d4945, 32'hc2ac04bd},
  {32'hc493f19b, 32'h4439cf75, 32'h4379b920},
  {32'h45189768, 32'h439f33c3, 32'hc1e9af56},
  {32'hc37d4408, 32'hc18af26e, 32'h436a5f5a},
  {32'h44a2e684, 32'h42e2b956, 32'h412a0722},
  {32'hc4441b42, 32'hc3410b97, 32'hc2b61cb3},
  {32'hc2b2eaa0, 32'hc3a8d6be, 32'h43d0c0df},
  {32'hc4cddc10, 32'h4310c276, 32'h43955ac6},
  {32'h44a40e56, 32'hc1ecd937, 32'h43b0813b},
  {32'hc4b50960, 32'h41f7dc78, 32'hc12bdb42},
  {32'h448bd526, 32'hc2be1a40, 32'h422da338},
  {32'hc4af0c4a, 32'hc395e30d, 32'hc13279ae},
  {32'h438ae385, 32'h42e3ef3a, 32'h43cffdd5},
  {32'hc0eb655d, 32'h43a55a2b, 32'hc3cbe359},
  {32'h433aaea0, 32'h418a79c6, 32'hc3c49732},
  {32'h434e3358, 32'h42eec4f1, 32'hc3753a94},
  {32'h44158b4e, 32'h43a2676c, 32'h42c1c36a},
  {32'hc4d80f24, 32'hc122fe6d, 32'hc0d9a01e},
  {32'h4482d984, 32'hc2cb0f6b, 32'h4317dfa1},
  {32'hc4c8fee8, 32'h439bd245, 32'hc386518c},
  {32'h4460238c, 32'hc34e6dd4, 32'h4373adfd},
  {32'hc4d97fae, 32'h4228733b, 32'hc403a24b},
  {32'h42e198e0, 32'hc356b6d0, 32'h43ad28d2},
  {32'hc3908cdc, 32'h4281a324, 32'hc3ba8c89},
  {32'h44f57165, 32'hc36dd92d, 32'h41bf152c},
  {32'hc404a9ac, 32'hc1aeb39e, 32'h41adeb01},
  {32'h43d2d420, 32'h40a6d840, 32'h437672f4},
  {32'hc435698a, 32'hc3b38864, 32'hc32bbb3e},
  {32'h42ad0ff8, 32'h4271f4f2, 32'h43631d63},
  {32'hc4b5fe5f, 32'hc2285cb7, 32'h42b58678},
  {32'h4483b54f, 32'h41a0d106, 32'h42710568},
  {32'hc4a88bdd, 32'h43dfe9fc, 32'h435c5e20},
  {32'hc22d2d0b, 32'h43f8b5b9, 32'hc3e8dc7f},
  {32'hc4832bd1, 32'hc1b22f0c, 32'hc334eec1},
  {32'hc2832ae0, 32'hc3b1547d, 32'hc0e38188},
  {32'hc3ddde34, 32'h43531c18, 32'hc3b0b936},
  {32'h449e6f3d, 32'h42c6ca1a, 32'hc2bc5991},
  {32'hc4b80aef, 32'h43251ee4, 32'hc2b99a6b},
  {32'h449edef9, 32'h43aaf911, 32'h423b4842},
  {32'hc48bea3a, 32'hc23b463b, 32'h4214f8d6},
  {32'h449d64d2, 32'hc2915bb4, 32'h413415bb},
  {32'hc421b138, 32'hc28d5110, 32'hc33ba2cf},
  {32'h43e6d390, 32'h43082c5d, 32'hc349f90f},
  {32'hc4bb5640, 32'hc24c8ca2, 32'h42ec3a98},
  {32'h44be2034, 32'h431cc297, 32'h41b9fd3a},
  {32'hc4a9dc18, 32'hc3fa7dbd, 32'hc230455e},
  {32'h4476a42a, 32'h413d66fb, 32'hc3a42b1e},
  {32'hc501568b, 32'h42d7ac16, 32'hc31e4104},
  {32'h4306e990, 32'hc15d19aa, 32'hc3aab5c9},
  {32'hc4903b4d, 32'hc3a37833, 32'hc3484264},
  {32'h442d1030, 32'h4372ed92, 32'hc2c4427e},
  {32'hc5162459, 32'h44073837, 32'h411cbb6a},
  {32'h45024497, 32'h415746b0, 32'h43293c4c},
  {32'h42d08d9d, 32'h43a9da5c, 32'hc30c2ec4},
  {32'h4449cbc5, 32'hc2637b46, 32'hc1e1a938},
  {32'hc45a2b20, 32'hc334d5ca, 32'h431888fe},
  {32'h441837ca, 32'hc3d8b020, 32'hc1b4608e},
  {32'hc426179a, 32'hc2d7634c, 32'hc29c1e17},
  {32'h4500ba6d, 32'h423f85d4, 32'hc23872b2},
  {32'hc41b6c96, 32'hc1ec2113, 32'h4404bdf9},
  {32'h449ba27c, 32'hc2abfd46, 32'h42213bd2},
  {32'hc3b99e6a, 32'hc30fd985, 32'hc3a33497},
  {32'h450c4eae, 32'h4045f888, 32'h4393113a},
  {32'hc4be6347, 32'hc3c73684, 32'h4348eda9},
  {32'h4492953e, 32'hc0bcd448, 32'hc352669e},
  {32'h4373f4bc, 32'h4324e862, 32'hc410a9c8},
  {32'h447390f4, 32'h434f3718, 32'h43111422},
  {32'hc46067b1, 32'hc3662288, 32'h43439f29},
  {32'h445502d4, 32'h42e979ca, 32'hc2e3ceff},
  {32'hc350f151, 32'hc31f0dbb, 32'h435ac467},
  {32'h44aea109, 32'hc385dd52, 32'h441667d0},
  {32'hc473b8af, 32'h413425b6, 32'h433d7143},
  {32'h44d8a7c5, 32'h435e7f5e, 32'hc37382cb},
  {32'hc4ac5f80, 32'h4176f1c0, 32'h43d2be5f},
  {32'h44abd790, 32'hc333cd07, 32'hc3a455bb},
  {32'hc50928e9, 32'hc33cf697, 32'h43b7d804},
  {32'h44f499e5, 32'h43d1b71c, 32'hc2f0d9d4},
  {32'hc4084fea, 32'h42194490, 32'hc28def65},
  {32'h44c334de, 32'h423570e5, 32'h43bb49fd},
  {32'hc5044bfc, 32'h43b16c3a, 32'hc3265390},
  {32'h4509140a, 32'hc30c6b36, 32'h439e0426},
  {32'hc501fd0a, 32'hc3bd7781, 32'h418e1384},
  {32'hc319b2ec, 32'hc38bf2a4, 32'hc3826d5a},
  {32'hc50fe4b1, 32'hc318ca7c, 32'h43a08412},
  {32'h44a34a92, 32'hc32a9e6b, 32'h427e0a3b},
  {32'hc51ff99a, 32'h4240adf4, 32'h4354151f},
  {32'h44c0c48a, 32'hc3aa8719, 32'hc2ec2f62},
  {32'hc3003023, 32'hc39a7740, 32'h43c43f0b},
  {32'h43fae4be, 32'hc3894535, 32'hc3c0cdcf},
  {32'hc4fc2e62, 32'h439ac8b5, 32'h42571653},
  {32'h44efa7cc, 32'hc10b0c50, 32'hc24f7843},
  {32'hc4d8ad74, 32'hc23887f0, 32'hc34e310b},
  {32'h44099416, 32'hc3c9dc3c, 32'h43a0d4f2},
  {32'hc4166e3e, 32'hc1d00292, 32'hc24829b3},
  {32'h45182434, 32'h430d8afe, 32'h42a363c0},
  {32'hc421ea50, 32'hc3a7c5e8, 32'h43acbb51},
  {32'h4418141e, 32'h40f1f509, 32'hc3027fd1},
  {32'hc49f1a8c, 32'h436a6d5f, 32'hc36b6129},
  {32'h42c7be42, 32'hc10ffc33, 32'hc4136552},
  {32'h43309d67, 32'h43179969, 32'h43034df1},
  {32'h44bb247c, 32'hc28ac261, 32'hc44f8af0},
  {32'hc4f41229, 32'hc26830df, 32'h43079689},
  {32'h44a34f7d, 32'hc342522a, 32'hc2ade9da},
  {32'hc39750f0, 32'h430aa21a, 32'h4304abb0},
  {32'h44a8c8a3, 32'h433216d1, 32'hc1f09f9b},
  {32'hc4f333a0, 32'h42504968, 32'h4139577e},
  {32'h44c8c93b, 32'hc37d5f66, 32'hc352f5d8},
  {32'hc45c97d8, 32'h4246d56f, 32'h42c8483f},
  {32'h4293e000, 32'h43011fc5, 32'h43a902b6},
  {32'hc4057a38, 32'hc22efd35, 32'h43531773},
  {32'h4517e4a4, 32'h439f1c2c, 32'h40cf7c40},
  {32'hc3dd2878, 32'h4143ec8c, 32'hc33e40ea},
  {32'h44e6eb4f, 32'hc3b2dffa, 32'h431c3dbc},
  {32'hc511cb26, 32'hc350f6b5, 32'h43faeac7},
  {32'h451412e2, 32'h428e8bcd, 32'h439d0900},
  {32'hc4f8225a, 32'h4299979c, 32'hc1c94c61},
  {32'h44c95282, 32'hc2bbd270, 32'hc2edd014},
  {32'hc2e56de8, 32'hc28e4abc, 32'h435c3fe5},
  {32'h44b50f64, 32'hc2e86c48, 32'hc36b54a4},
  {32'hc40d00a2, 32'h433272d4, 32'hc319112d},
  {32'h434a3cf0, 32'h41a8ccda, 32'hc3436a55},
  {32'hc46ebb10, 32'hc2995896, 32'hc3428439},
  {32'h44d2b287, 32'h43cbf4af, 32'h40bffb95},
  {32'hc4e19b8b, 32'hc344aabe, 32'h4388096e},
  {32'h450dba43, 32'h431ac7d9, 32'hc30d4b99},
  {32'hc4fa157a, 32'hc13346e1, 32'hc227fe98},
  {32'h44d566b3, 32'h42a31d28, 32'hc39c55b5},
  {32'hc46c3402, 32'hc3785740, 32'h425246bf},
  {32'h43b7869e, 32'h43afa6f0, 32'hc26579cc},
  {32'hc475f95b, 32'h40cdcccc, 32'h4214c897},
  {32'h44e91793, 32'h43d8f1b1, 32'hc3a71912},
  {32'h45163587, 32'h432251c5, 32'h43eb5f35},
  {32'hc3c07f66, 32'h416c4a69, 32'hc2283c84},
  {32'h44c9aa32, 32'h4344faff, 32'h439285cc},
  {32'hc4cad4bb, 32'h422f8e1f, 32'hc20b1af6},
  {32'h44df5f7e, 32'hc2ffbd30, 32'hc2f495fb},
  {32'hc5049d07, 32'hc180661b, 32'h431c8d2c},
  {32'h44e0ad3c, 32'h420735de, 32'hc2897879},
  {32'hc49c5992, 32'h42f1911a, 32'h42b07c3c},
  {32'h44589c8c, 32'h431779a0, 32'hc385342c},
  {32'hc500d4ca, 32'hc3a420ca, 32'hc3d080be},
  {32'h43be7497, 32'h4338ebe7, 32'hc3073907},
  {32'hc44a03f3, 32'hc3cae641, 32'h438d350f},
  {32'h45093e92, 32'h4306a31f, 32'h43ec666a},
  {32'hc3beb8ab, 32'hc32b3869, 32'hc30cd8c4},
  {32'hc1f2771c, 32'hc3255c8b, 32'hc3c04d7c},
  {32'hc4db1221, 32'h43a1950d, 32'hc30c575f},
  {32'h44186187, 32'hc3f296ea, 32'hc391f903},
  {32'hc405687b, 32'hc38280a2, 32'h41ed0239},
  {32'h450fe4e5, 32'h43ab6409, 32'hc1bbbdfe},
  {32'hc479ffe8, 32'hc2f8772e, 32'h43bc9290},
  {32'h4505dc64, 32'h4338416f, 32'hc33246b8},
  {32'hc47d8d9e, 32'hc1dd3182, 32'h43b8f092},
  {32'h45147ce7, 32'h4304421a, 32'hc20f95c6},
  {32'hc4e20026, 32'hc3379754, 32'hc36f4587},
  {32'h44b81607, 32'hc1ce96bd, 32'hc318c9b2},
  {32'hc4fe4e9f, 32'hc34e4823, 32'h42ca3a1d},
  {32'h44b08dba, 32'hc3e175cf, 32'h411ec24c},
  {32'hc361bc68, 32'h4310848e, 32'h42c059f5},
  {32'h449aaf6d, 32'h40f09624, 32'h433a8acd},
  {32'hc4cac9df, 32'h43ae4dc2, 32'h4316fd26},
  {32'h42867cd4, 32'h43f83964, 32'hc2a16ed5},
  {32'hc3adc2aa, 32'hc31bef45, 32'hc2f31b6e},
  {32'h450255b2, 32'h41968290, 32'h42d34534},
  {32'hc32ff34c, 32'hc3042d09, 32'h432d382f},
  {32'h4507ed98, 32'h4166251c, 32'hc36c7795},
  {32'hc31d563e, 32'hc3a403e8, 32'h438d401e},
  {32'h44ccadff, 32'hc2f67374, 32'hc020e2ee},
  {32'hc377eac8, 32'h433cc477, 32'h413fd965},
  {32'h440b39be, 32'h40d2f4e3, 32'hc32cdf77},
  {32'hc487f330, 32'hc3a5f38f, 32'hc40da512},
  {32'h450ec7b4, 32'hc3397c6c, 32'hc3822cc0},
  {32'hc49b2daa, 32'hc2855cf4, 32'hc3e000c7},
  {32'h45188f7b, 32'h4225f666, 32'h438ebf5f},
  {32'hc4c709d8, 32'hc3072ff9, 32'hc2c662ab},
  {32'h4474673d, 32'hc3c881f7, 32'h42901f9c},
  {32'hc48d552d, 32'hc10ba21f, 32'h43bad5bc},
  {32'h438d5fca, 32'h4180d7b7, 32'hc31901dd},
  {32'hc36b3810, 32'hc2db9bae, 32'hc315cc43},
  {32'h4470bbe4, 32'h43b0e404, 32'h438da164},
  {32'hc50c7f5e, 32'h431de6ae, 32'h42395bad},
  {32'h4432398f, 32'h435bcde1, 32'hc2838c14},
  {32'hc49ea91a, 32'hc3222db3, 32'hc2c7940c},
  {32'h44acd2e5, 32'hbe6ff900, 32'h43a8bb06},
  {32'hc5100a50, 32'hc37090c9, 32'h43049438},
  {32'h43da9b08, 32'h42b7941c, 32'hc375db15},
  {32'hc4b61422, 32'hc306498b, 32'hc3859360},
  {32'h442c4b2e, 32'h42af1156, 32'h4314e282},
  {32'hc4a984f4, 32'h42cb213d, 32'hc3338922},
  {32'h450c8935, 32'hc2acba9c, 32'h424c2ff6},
  {32'hc2e5d2e0, 32'hc3ea4e81, 32'h44566f3e},
  {32'h44d93586, 32'hc361fd1d, 32'hc42919ea},
  {32'hc43aab6b, 32'h42955cca, 32'h424a8519},
  {32'h448b9e96, 32'h4316c33a, 32'h43a56aba},
  {32'hc46fbc7b, 32'h4395f139, 32'hc35049e9},
  {32'h450e96a3, 32'h4408621e, 32'h4392f728},
  {32'hc34800b0, 32'h43043652, 32'hc1fddb12},
  {32'h447ae460, 32'h42cd9d31, 32'hc3016f26},
  {32'hc480ba01, 32'h438cec5f, 32'h4307dde2},
  {32'h45002942, 32'hc1ca67cd, 32'hc2895b6f},
  {32'hc4a094d6, 32'h434f0d99, 32'hc351d1c8},
  {32'h448cc6a1, 32'hc2cf738d, 32'h4343e306},
  {32'hc4b65db9, 32'hc402b6ac, 32'hc2dafae3},
  {32'h44c04ac5, 32'h43382a8c, 32'h439d7a08},
  {32'hc512738a, 32'hc19abec8, 32'h440c08ed},
  {32'h43cc1e67, 32'h43594211, 32'h434cea38},
  {32'hc46b206f, 32'hc2b4b7a8, 32'h4165a252},
  {32'h4514e326, 32'hc35eb918, 32'hc3d0e981},
  {32'hc4b91507, 32'h43aa4d10, 32'h43962b81},
  {32'h44c14147, 32'h4345e5ea, 32'h43b41cd3},
  {32'hc4130d18, 32'h42c65538, 32'hc397e480},
  {32'h44d8a711, 32'h437c5482, 32'hc23aaa54},
  {32'hc4e0ac72, 32'h41b98e63, 32'hc2ff7bcb},
  {32'h449550dd, 32'h434c46fa, 32'h42d668b0},
  {32'hc4ee57cf, 32'h43d77c18, 32'h41140f7b},
  {32'h45080886, 32'hc2ce1170, 32'h42e7b2ca},
  {32'hc4083304, 32'hc2179b3a, 32'hc18ed445},
  {32'h44be9163, 32'hc3526d11, 32'h42405bf7},
  {32'hc456e193, 32'hc3803d1c, 32'h42831a06},
  {32'h4463c4f2, 32'hc3babd76, 32'h436a1491},
  {32'hc4e881a6, 32'h4322ed4a, 32'h41a047d8},
  {32'h45110036, 32'h435a9d98, 32'h41b0a6b4},
  {32'hc470a432, 32'h4309ff69, 32'h4384c05d},
  {32'h44690a00, 32'hc38ce33b, 32'hc306247f},
  {32'hc3ac1c3a, 32'h43ba4315, 32'hc3196cd0},
  {32'h43e574f7, 32'hc340adfb, 32'h4336d672},
  {32'hc16f810c, 32'h430d37f0, 32'hc36bafd9},
  {32'h448c68e8, 32'h4307675d, 32'h43a420f0},
  {32'hc50b4dc6, 32'hc20b226d, 32'hc3e0d678},
  {32'h44d11ada, 32'hc33708b7, 32'hc3b3916b},
  {32'hc4150a45, 32'h428ebde5, 32'hc228ec36},
  {32'h44bdcd78, 32'h43114a79, 32'hc2977a5a},
  {32'hc4d1d962, 32'hc1d8f0d0, 32'hc03c8c28},
  {32'h44959d9e, 32'h430a9797, 32'h42aee210},
  {32'hc4e2f643, 32'h429ddb4a, 32'h438779a2},
  {32'h44d1cf61, 32'h43934ce2, 32'h42ddabb7},
  {32'hc4c83655, 32'hc36d680a, 32'h42860dc9},
  {32'h43b7c15d, 32'h43337b39, 32'hc3663497},
  {32'hc4dcae94, 32'h43831918, 32'hc1b99977},
  {32'h4482c3b5, 32'hc3c8a9e0, 32'h43854d1d},
  {32'hc4159a04, 32'hc311e34e, 32'hc2c6bd32},
  {32'h44e7662c, 32'h43a53070, 32'h4387336e},
  {32'hc4d2965a, 32'h42ad2a25, 32'h43532c4c},
  {32'h42f4a908, 32'h43308726, 32'hc2039204},
  {32'hc492c0e6, 32'h432067cc, 32'h42c49418},
  {32'h44e61b48, 32'h4295ebd9, 32'hc32e20a0},
  {32'hc42f840f, 32'hc19b4d7e, 32'hc3100687},
  {32'h44f3287d, 32'h4335da3e, 32'hc06de9a1},
  {32'hc50fb22a, 32'h4367a478, 32'h4176152a},
  {32'h439d085a, 32'hc337d34e, 32'hc2a8389a},
  {32'hc4b06908, 32'h41b0c7db, 32'hc2e6ab3c},
  {32'h4505fbe5, 32'hc2f8c097, 32'h4380247b},
  {32'hc291f6a0, 32'h4045c450, 32'h4359c4a2},
  {32'h44f476f4, 32'h430363a6, 32'h415950e6},
  {32'hc4dbe648, 32'hc13289fa, 32'h436e673c},
  {32'h443e3191, 32'hc386b1d5, 32'hc3f96891},
  {32'h41d77090, 32'h432c36dc, 32'hc2dc9359},
  {32'h44a421ef, 32'hc29f4005, 32'h43ed9faa},
  {32'hc48de7bf, 32'h430284aa, 32'hc2921b19},
  {32'h44b74de5, 32'h42d44e95, 32'hc36dc676},
  {32'hc4b352a2, 32'h43949276, 32'h42df1508},
  {32'h44da83c5, 32'hc35e0562, 32'h43ae4bf0},
  {32'hc4ea23dd, 32'h435d9af8, 32'hc2ee7343},
  {32'h440f4200, 32'hc38da125, 32'hc38c96fa},
  {32'hc30a3c00, 32'hc3636838, 32'hc29e520a},
  {32'h449418a0, 32'h43e6ada0, 32'hc137403a},
  {32'hc4e7c50a, 32'hc2ebb33c, 32'hc3044aa5},
  {32'h44f04a24, 32'hc1d03dda, 32'hc287a553},
  {32'hc4af1654, 32'h42acde63, 32'h43b564aa},
  {32'h44a781e2, 32'h42afe452, 32'hc20c86aa},
  {32'h41cad8e0, 32'hc4564b49, 32'h430598d6},
  {32'h44c6dc3f, 32'hc35e222e, 32'hc29fde3f},
  {32'hc42a15cc, 32'hc32a038c, 32'hc3a9e8cc},
  {32'h441e7ecf, 32'h4312af76, 32'h42f035b6},
  {32'hc4defdbe, 32'hc0f34206, 32'h42fc8db7},
  {32'h442df5e8, 32'hc3977653, 32'h43adc47f},
  {32'hc3f75ac6, 32'hc01eb413, 32'hc3a71b11},
  {32'h441563d7, 32'h438e4a36, 32'hc327b21f},
  {32'hc469c714, 32'hc3307ded, 32'hc25adf67},
  {32'h4338328e, 32'h421d3c8b, 32'hc27e665f},
  {32'hc4b578ac, 32'hc2c04312, 32'h425942a3},
  {32'h44b6b267, 32'hc300bc3f, 32'h428469a2},
  {32'hc4f3fb9c, 32'h421a05a7, 32'h43182499},
  {32'h44b92cc4, 32'hc3a968eb, 32'hc34aee70},
  {32'hc2f979f0, 32'hc1f9fdce, 32'h437121b3},
  {32'h4426f1a6, 32'h42f53b4b, 32'hc37f4767},
  {32'hc407f938, 32'hc14607ea, 32'h43074453},
  {32'h44e25496, 32'hc3b7539c, 32'hc37560e0},
  {32'hc51e13f2, 32'hc37a2ca2, 32'hc36dcc08},
  {32'h44b40c49, 32'h4386a402, 32'hc3c98a9b},
  {32'hc41e8ee0, 32'hc1aa28d8, 32'hc0d177c1},
  {32'h44f07775, 32'hc2ea4133, 32'hc375c468},
  {32'h42738a40, 32'h4323ec89, 32'h43aae7a5},
  {32'h44002f69, 32'h42e88f8e, 32'hc3adc577},
  {32'hc4eb9a69, 32'hc0f0d330, 32'hc3383695},
  {32'h450a3246, 32'h42f94af6, 32'h42dbd69e},
  {32'hc3e37d13, 32'h420dc3ff, 32'hc39cc1f2},
  {32'h450e6d34, 32'hc38bde35, 32'hc34087a9},
  {32'hc49afe7d, 32'hc30fc306, 32'h4350e17c},
  {32'h446a3bc2, 32'hc282494e, 32'hc1010b24},
  {32'hc4f212d0, 32'h42b7f2d0, 32'hc0dc2f85},
  {32'h44bb0586, 32'hc33ac293, 32'hc2012e0e},
  {32'hc48d4c35, 32'hc2351e8d, 32'hc289c4bc},
  {32'h44a5079d, 32'hc3c53e40, 32'hc400dc8d},
  {32'hc45e5527, 32'hc2f03aa7, 32'hc37fd4a7},
  {32'h442b428e, 32'hc2ed9ee8, 32'h436adeb4},
  {32'hc494daa4, 32'h4285fa08, 32'h42c531b7},
  {32'h450afef1, 32'hc3fd9397, 32'hc368cf21},
  {32'hc3f051a8, 32'h4352e5b2, 32'hc299462f},
  {32'h446591ab, 32'h4271c6dc, 32'hc33cdb18},
  {32'hc43b2000, 32'hc29ce095, 32'h42d4b672},
  {32'h4476ea76, 32'h42858128, 32'hc2fc0794},
  {32'hc47bad93, 32'hc22f0de4, 32'h43b0e309},
  {32'h44d076c5, 32'h3f7ec797, 32'h41c38988},
  {32'hc447b07b, 32'hc2aa1141, 32'h433507fa},
  {32'h43e70288, 32'h4322c6f4, 32'h41f765fc},
  {32'hc318a340, 32'hc2ba4f37, 32'h43853b2c},
  {32'h44e7e27f, 32'h43625302, 32'hc382a7bc},
  {32'hc4f455e9, 32'h410eaf8b, 32'h439fa72a},
  {32'h45212012, 32'h4303a394, 32'hc3602a19},
  {32'hc4f48daa, 32'h43f3b37d, 32'hc2e21a0c},
  {32'h441ab8d8, 32'hc375d839, 32'h44128230},
  {32'hc4d0a6e3, 32'hc1eabb18, 32'hc4311752},
  {32'h447a4764, 32'hc2999fcc, 32'hc402a97a},
  {32'hc380e8f8, 32'h4352fd2c, 32'h438db260},
  {32'h44955cc3, 32'h41dccbb7, 32'hc257ae32},
  {32'hc493ee4d, 32'hc262453d, 32'hc2a55270},
  {32'h44616d10, 32'hc36de2a0, 32'hc21c094b},
  {32'hc4aa5b25, 32'h420a92a4, 32'hc1a89986},
  {32'h44cf15e1, 32'h43ad534b, 32'h43552e69},
  {32'hc43f492c, 32'hc31e830e, 32'h420b3428},
  {32'h450b71dd, 32'h42712749, 32'h43ad6a06},
  {32'hc4d23af5, 32'h4303c161, 32'h42f24de2},
  {32'h44a30f7d, 32'hc1f9a1dc, 32'h42049bf8},
  {32'hc473c2b1, 32'hc30a1d4c, 32'h4305a804},
  {32'h4442891e, 32'h434ddcce, 32'hc1cc7106},
  {32'hc469eb09, 32'h43656345, 32'hc18f7e5c},
  {32'h42b2efe4, 32'hc2ae34cb, 32'hc224ba2b},
  {32'hc5007c9f, 32'h42f61e6b, 32'h43ddfd42},
  {32'h450cb008, 32'h42a66f15, 32'h4118e751},
  {32'hc4d81286, 32'h4392105e, 32'hc33c1bf1},
  {32'h43de42b9, 32'h43c4b264, 32'hc2467fe1},
  {32'hc402a24a, 32'h422d539e, 32'hc3f295c1},
  {32'h4462616e, 32'hc304f586, 32'h43b90ab9},
  {32'hc374fbe0, 32'hc3bbb4b5, 32'h4344ba68},
  {32'h44ce9765, 32'hc2a50434, 32'h43dcd927},
  {32'hc3cb2625, 32'hc32eb421, 32'hc37e7cbc},
  {32'h445a3eda, 32'h431e368d, 32'hc288664d},
  {32'h430718f0, 32'h422e5936, 32'h42830975},
  {32'h44343ce6, 32'h425f7109, 32'h433af964},
  {32'hc4bd7b68, 32'hc394f8e3, 32'h40949acf},
  {32'h4409e6f4, 32'h431bb8e1, 32'hc21daf8b},
  {32'hc2e70540, 32'h42d30676, 32'h43cb6d31},
  {32'h44833cc8, 32'h4303ad29, 32'hc2956083},
  {32'hc498cdbf, 32'hc386541b, 32'hc3972740},
  {32'h4412eda0, 32'h435b24e3, 32'h439a244f},
  {32'hc48cde24, 32'h42e0b579, 32'hc311fbf1},
  {32'h44f6749e, 32'hc2f18274, 32'hc3251f86},
  {32'hc503d1ff, 32'h438ff0bf, 32'hc2ed1992},
  {32'h433956f0, 32'hc321d664, 32'hc34dc42a},
  {32'hc505d21a, 32'h424f1a4e, 32'hc11df436},
  {32'h443929be, 32'h433b88b4, 32'hc30cce76},
  {32'hc416d498, 32'h43150806, 32'hc35a44fc},
  {32'h44367b27, 32'h424f41d8, 32'hc31ac132},
  {32'hc4e335ea, 32'h4295c46a, 32'h4219611a},
  {32'h44075d84, 32'hc297cbd8, 32'hc34a41fa},
  {32'hc482822e, 32'h43693f54, 32'hc37f49eb},
  {32'h44ec2f00, 32'hc24b7113, 32'hc2b64929},
  {32'hc309e5f0, 32'h431d68bb, 32'h413189ac},
  {32'h446d6a08, 32'h4310eafc, 32'h42a23994},
  {32'hc4898a5a, 32'h439a27bd, 32'h42ea71de},
  {32'h4501ea2d, 32'hc1d7c59b, 32'h42be0682},
  {32'hc505b271, 32'h427dbcaa, 32'hc33db8f4},
  {32'h43a65050, 32'hc23c9f8e, 32'h425f7a4e},
  {32'hc4259700, 32'h42a9f745, 32'h42bd845a},
  {32'h439fd837, 32'hc38622f0, 32'hc3408532},
  {32'hc2ce88e0, 32'h4378d89a, 32'hc24e7662},
  {32'h44776c47, 32'h43641331, 32'hc3508e14},
  {32'hc4dd71c6, 32'hc3cf88dd, 32'h423782d1},
  {32'h44c56d9a, 32'hc21e9be2, 32'hc2fbde2f},
  {32'hc42f717e, 32'hc4047ff7, 32'h438c94cf},
  {32'h44794b4a, 32'h4280cb32, 32'hc1de5795},
  {32'h438f2d76, 32'hc37b615c, 32'hc34b8212},
  {32'h4482c363, 32'h43de478b, 32'hc11ee486},
  {32'hc4172268, 32'hc3529a07, 32'h432afade},
  {32'h44db8309, 32'hc3ce2f08, 32'h431210c7},
  {32'hc4c999c2, 32'h43583dbb, 32'hc40933ee},
  {32'h43e0f6ac, 32'hc288ab8e, 32'h42ed7c37},
  {32'hc40e0dc8, 32'hc242b4e0, 32'h433808e3},
  {32'h451c68c9, 32'hc342d34c, 32'h4396f7dc},
  {32'hc49662ec, 32'h42d10b5f, 32'h436d778c},
  {32'h440ca39c, 32'hc403f4d6, 32'h42c273a0},
  {32'hc50ee5d4, 32'hc34d7dba, 32'h434b2ecd},
  {32'h444aaa86, 32'hc2d98213, 32'h423701d9},
  {32'hc3457b43, 32'hc08fd299, 32'h43403325},
  {32'h44aed21b, 32'hc2d25898, 32'hc2cb36ce},
  {32'hc48e2928, 32'hc2db216c, 32'h4381b78f},
  {32'h430c98ae, 32'hc3a61863, 32'h42740756},
  {32'hc42a9ef9, 32'h42f848c7, 32'h423653e1},
  {32'h4414b33c, 32'h429fc439, 32'hc3cfdf80},
  {32'hc4a6ef5f, 32'hc22f3092, 32'h42d079b6},
  {32'h4434976c, 32'hc3888a17, 32'hc3bd97b3},
  {32'hc388e072, 32'h426b06d5, 32'h43394223},
  {32'h44aed198, 32'hc2310829, 32'hc3a7a5f2},
  {32'hc474273e, 32'h4363000a, 32'hc2721e23},
  {32'h43cb0a71, 32'h42041a60, 32'hc351dfc5},
  {32'hc4f58e83, 32'h430fa5e5, 32'hc2a26171},
  {32'h45072cf4, 32'hc1bb75f9, 32'hc0d46fa3},
  {32'hc48ac258, 32'hc2126812, 32'hc1a260ae},
  {32'h443317a5, 32'hc3246b33, 32'hc2ca5eb0},
  {32'hc4261615, 32'hc3a662e6, 32'hc32cb35a},
  {32'h4490490d, 32'hc38c915e, 32'hc27aecfc},
  {32'hc4c150ec, 32'h42d13c91, 32'hc2b05b91},
  {32'h441c168e, 32'h4332421e, 32'h42cf10b8},
  {32'hc4dfd945, 32'h42041a48, 32'h42fc06ba},
  {32'h446a2b61, 32'h438ce8cc, 32'hc38bb9a1},
  {32'hc4daf532, 32'hc328504e, 32'hc35dc205},
  {32'h43b7e5d7, 32'hc341ffe3, 32'h4307896f},
  {32'hc3bd05c1, 32'h44052d77, 32'h43ce3f24},
  {32'h43bf3c13, 32'h42b52f2e, 32'h416dee6b},
  {32'hc4e91ea1, 32'hc1dc0e4f, 32'hc2c7b1c6},
  {32'h44a7a262, 32'hc352902d, 32'hc38e1580},
  {32'hc44069da, 32'hc379dc54, 32'h43c3700d},
  {32'h44d429e4, 32'h42ec907a, 32'h42be28e4},
  {32'hc446bcec, 32'hc22e7914, 32'h4341b7a1},
  {32'h43086d00, 32'h439c65ee, 32'hc35db5d5},
  {32'hc33f5173, 32'hc302462a, 32'hc308a57e},
  {32'h4468e914, 32'h4239e5b3, 32'h438c7ab6},
  {32'hc4c9f031, 32'hc389d0f5, 32'hc2d65cd3},
  {32'h44ae88e4, 32'hc3065599, 32'hc311a979},
  {32'hc428edb4, 32'hc0e4e27e, 32'h3fd66966},
  {32'h44962388, 32'hc3e00a55, 32'hc180f6e2},
  {32'h42f5e9e0, 32'hc3964a1b, 32'hc34b60b4},
  {32'h44cce9b9, 32'h4230ced5, 32'hc3281e8f},
  {32'hc4fadade, 32'hc403add8, 32'h4277fab4},
  {32'h4489dc40, 32'hc318a133, 32'hc16a0e1e},
  {32'hc4c9c9a1, 32'h3ea80370, 32'h43634256},
  {32'h44dd9f2a, 32'h43bff8ac, 32'h4002ae9c},
  {32'h42ce4100, 32'hc3a99ffc, 32'h43b36bf2},
  {32'h44b6dc52, 32'h420fcf12, 32'h44417bbc},
  {32'hc4fec8ae, 32'h438828b1, 32'hc39f9fe2},
  {32'h4460f8da, 32'h432ef879, 32'h43456c32},
  {32'hc4e1d01c, 32'hc288e1ea, 32'hc2a293cc},
  {32'h44e2b446, 32'hc29ae7e2, 32'h42940a39},
  {32'hc4c598d4, 32'hc16d0c1e, 32'h42b17928},
  {32'h452126b5, 32'hc3ac6715, 32'hc3a3c648},
  {32'hc4ce2da2, 32'hc322e084, 32'h42c539ac},
  {32'hc0e0c2c0, 32'h430b9883, 32'hc2bda3e7},
  {32'hc41ad5a0, 32'h439c33e7, 32'h438b3e63},
  {32'h439c611b, 32'hc354fe35, 32'h42a870bd},
  {32'hc42b3f8e, 32'hc30e8b90, 32'h422cad37},
  {32'h450b0543, 32'hc336765f, 32'h434b33f0},
  {32'hc4eb27fe, 32'hc3fda582, 32'hc2b6f7d9},
  {32'h43d57751, 32'hc3a7fb5b, 32'hc371740c},
  {32'hc422a014, 32'hc31d9226, 32'h4284e45c},
  {32'h447dbbda, 32'h430b8ec3, 32'h43535c34},
  {32'hc463944e, 32'hc2e7f714, 32'hc30c4fe3},
  {32'h444a0533, 32'h432fcc09, 32'h42c02196},
  {32'hc516bfcb, 32'hc3a981df, 32'h4366f0c7},
  {32'h44f38a1d, 32'hc28d5104, 32'h426754c2},
  {32'hc4249948, 32'hc312617c, 32'h416f103d},
  {32'h44dcb770, 32'hc30120cd, 32'h42a2cdcf},
  {32'hc4c84f8c, 32'h43722c2e, 32'hc39ee992},
  {32'h4499201d, 32'h439b6b03, 32'hc354a7ee},
  {32'hc48090a3, 32'hc34b02d0, 32'h4394d8e6},
  {32'h44cd7a8e, 32'h428e1214, 32'hc3ad70b7},
  {32'hc4f103c8, 32'hc31c5708, 32'hc2718617},
  {32'h444f9753, 32'hc3247da5, 32'h41daaf1b},
  {32'hc3e5e6ac, 32'hc2397b00, 32'hc2a8230a},
  {32'h44c80061, 32'h430ca04d, 32'hc2bd2a4d},
  {32'hc3d16968, 32'hc3248dd7, 32'h42f5f610},
  {32'h44dd1963, 32'h4395faf7, 32'h42e10519},
  {32'hc3b849ce, 32'hc2cbd2c4, 32'hc3be5c89},
  {32'h44a01415, 32'h42e72f7e, 32'h43b3bbe6},
  {32'hc4f3f097, 32'h416d0497, 32'hc29e8834},
  {32'h43349d50, 32'hc313e199, 32'h433191c3},
  {32'hc414fcaa, 32'h4385da56, 32'hc3185069},
  {32'h45094d1a, 32'hc34c7c5a, 32'hc34095c1},
  {32'hc47017f2, 32'h433f3977, 32'h40c62cda},
  {32'h43371018, 32'hc395ed6e, 32'h4256f24b},
  {32'hc4c97d35, 32'hc328d66a, 32'hc365c901},
  {32'h450283b2, 32'hc3442e08, 32'h433f2fba},
  {32'hc4842ca4, 32'h434c943e, 32'h4293232e},
  {32'h441cdad1, 32'h4386b219, 32'hc3cf159b},
  {32'hc51b4dac, 32'h438786c5, 32'h42d2ba16},
  {32'h450c28fb, 32'hc35aaa98, 32'hc31edc3b},
  {32'hc30eca0c, 32'h42a61af8, 32'h41bf6d6f},
  {32'h44b34afd, 32'hbfcb01e8, 32'h43d970e7},
  {32'hc4cbf6ba, 32'hc354e3e1, 32'h4243cf31},
  {32'h44fd1ff5, 32'hc3758deb, 32'hc1a959aa},
  {32'hc480b0a2, 32'hc31851f2, 32'h43b49fde},
  {32'h4522df62, 32'hc3d1b32d, 32'hc38d47d7},
  {32'hc4b4baaa, 32'h438f45bd, 32'hc254b83c},
  {32'h4515d376, 32'hc3126834, 32'h4383a855},
  {32'hc51c3e33, 32'h43923a08, 32'hc3b19b87},
  {32'h450a02ea, 32'hc36f0151, 32'h43c4621c},
  {32'hc4e76cab, 32'hc3b4759a, 32'hc397901b},
  {32'h449ff500, 32'h42c305f4, 32'hc37017bc},
  {32'hc4f5a1fa, 32'hc19e3830, 32'hc244f0a0},
  {32'h44bb4310, 32'h4225d205, 32'hc250ff8f},
  {32'hc49ac09c, 32'hc3f5d1fa, 32'hc11d762e},
  {32'h44ddaef0, 32'hc3834a43, 32'hc333e2ca},
  {32'hc419f2c2, 32'hc2d7fa87, 32'h4054ffed},
  {32'h44dcd93e, 32'h43b47a93, 32'h422a1032},
  {32'hc477d86b, 32'hc1d4ebac, 32'hc27430c2},
  {32'h4509b0b0, 32'hc2b84123, 32'hc2b21c95},
  {32'hc42af418, 32'h42fa3c31, 32'h420e74a7},
  {32'h45009347, 32'h4405d9a9, 32'h41bf22f0},
  {32'hc49ed2e5, 32'hc1dd0cd4, 32'hc241fd86},
  {32'h445b1e48, 32'hc17775d8, 32'h43742458},
  {32'hc3b9b390, 32'hc2e1fd30, 32'h43824ca0},
  {32'h430d1230, 32'hc2e5e3cb, 32'hc392a602},
  {32'hc4369e01, 32'h439184d6, 32'hc2a7d676},
  {32'h439e59f7, 32'hc2994c93, 32'h4331a754},
  {32'hc51cd9df, 32'hc18c077c, 32'hc3e71df1},
  {32'h4509f070, 32'hc2d49cbd, 32'hc3218983},
  {32'h43155cd0, 32'h43009af7, 32'hc404e72c},
  {32'h4445cd68, 32'hc342b7f1, 32'h4298a1b4},
  {32'hc4ee1c55, 32'h433fa943, 32'h429489c3},
  {32'h445a0645, 32'hc35be448, 32'h43ca189f},
  {32'hc47ceacb, 32'h43dc9d3e, 32'hc31febd4},
  {32'h43cd5368, 32'hc3da23f0, 32'hc256af8b},
  {32'hc40b2252, 32'hc3b1c3c7, 32'h43777a5c},
  {32'h44dff26d, 32'h4013525b, 32'hc318c5bd},
  {32'hc522a48a, 32'h44178426, 32'hc3cfbe27},
  {32'h449668b0, 32'h43a55fda, 32'hc29d1ef4},
  {32'hc4af13da, 32'hc38c90dc, 32'hc2bd1523},
  {32'hc1ab0170, 32'h42e14171, 32'h406a757c},
  {32'hc4b18b1b, 32'h439db641, 32'h4380c2a9},
  {32'hc19db480, 32'h4345e197, 32'h4395f5f0},
  {32'h42588ec0, 32'hc38814db, 32'hc2a475a0},
  {32'h43d434d1, 32'hc3ee50dd, 32'hc357f1c3},
  {32'hc28f9a3c, 32'h43b24080, 32'hc29ef2b0},
  {32'h44ac93e0, 32'h44094536, 32'h439531a6},
  {32'hc48e405e, 32'hc35bfde6, 32'hc304c890},
  {32'h44a01da7, 32'hc2744ff9, 32'h43a344c4},
  {32'hc3ebc9a0, 32'hc3f23d67, 32'hc2cf86cc},
  {32'h44348b9c, 32'hc3a4e287, 32'h416f3bc0},
  {32'hc4c334ea, 32'h4293b5fb, 32'hc2e16d89},
  {32'h42cd5cc0, 32'h4384ef89, 32'h4367f79a},
  {32'hc4a5f48e, 32'hc1a0d3a6, 32'h42ac3615},
  {32'h440fa6d4, 32'h43f75419, 32'h41cb5c44},
  {32'hc4f5b1c1, 32'hc2aadf5c, 32'h413dc5c6},
  {32'h44bfab61, 32'hc34ebb46, 32'h43f8508d},
  {32'hc4b8cde4, 32'hc37a7527, 32'h43180de8},
  {32'h44ea9e55, 32'hc1c0630f, 32'h4343fa78},
  {32'hc4117984, 32'hc3841e66, 32'h435a88dd},
  {32'h450547b7, 32'h433619f1, 32'h42ba567d},
  {32'hc3fe96aa, 32'h421a7f6a, 32'hc17d8da8},
  {32'h44edd660, 32'hc38e24ff, 32'h42b48f75},
  {32'hc38cffa8, 32'h41a0ba6a, 32'hc05f8480},
  {32'h43cb4f34, 32'hc26903a2, 32'hc2b1b9f0},
  {32'hc5096912, 32'h431e2e56, 32'h43557b39},
  {32'h44ad9729, 32'h42665c09, 32'h431e60c8},
  {32'hc4be48f7, 32'h42c70151, 32'hc1f69a9b},
  {32'h444db7be, 32'h431c9aef, 32'hc1efab30},
  {32'hc49bcd3a, 32'h4326a949, 32'hc38ee9a7},
  {32'h44b44699, 32'h42f03f12, 32'h4245354b},
  {32'hc490917e, 32'h42f0bc9f, 32'hc29865b5},
  {32'h44ab8a13, 32'hc243982d, 32'h429151ff},
  {32'hc390cb40, 32'hc26379df, 32'h4325161e},
  {32'h449ec9f7, 32'hc33fa2c2, 32'hc2b7cecd},
  {32'hc4bc17bf, 32'h42c7eb4f, 32'hc364f182},
  {32'hc47ac34a, 32'h4367e50b, 32'hc2cfc7a1},
  {32'h440375ce, 32'h42e163fd, 32'hc2f3416c},
  {32'hc41aa2b0, 32'hc3acd34a, 32'hc433d0bb},
  {32'h44b3cf85, 32'h434f986c, 32'h42cbbb96},
  {32'hc4c998f0, 32'hc3bb28e9, 32'hc372dfe0},
  {32'h4481044c, 32'hc2ee749b, 32'h43e34482},
  {32'hc303d260, 32'h42ea5880, 32'hc31d9aa2},
  {32'h44006062, 32'h41f800c3, 32'h431899d6},
  {32'hc515254f, 32'hc39ffd81, 32'hc358594d},
  {32'h44ffd950, 32'h42e3fc7a, 32'h433e4e2c},
  {32'h4406a7f9, 32'h42840038, 32'hc31952b4},
  {32'h44b86352, 32'h43a673f0, 32'h423c272a},
  {32'hc4e93d81, 32'h43ad0d13, 32'h42fc22c4},
  {32'h44ee5175, 32'hc39046e5, 32'h434b576a},
  {32'hc333bc78, 32'h43ae62ef, 32'hc1f68390},
  {32'h439b36d2, 32'hc2e83590, 32'hc23ef062},
  {32'hc2d95e60, 32'h438f9596, 32'h42e3908e},
  {32'h443dbc2b, 32'hc1ed6bf2, 32'h437590ee},
  {32'hc38a86b2, 32'hc29fa6f2, 32'h41d7a556},
  {32'h4432e94c, 32'hc2a2667f, 32'h434180b1},
  {32'hc49ac375, 32'hc2974ae6, 32'hc39884e8},
  {32'h445ce96e, 32'h43268be6, 32'h4221c3b3},
  {32'hc470dc89, 32'hc29f9c2c, 32'hc3961722},
  {32'h4440401a, 32'h41b5fa73, 32'h43992262},
  {32'hc43a2e88, 32'hc426fa09, 32'hc3498f5e},
  {32'h450cff86, 32'hc2035e90, 32'h430555ee},
  {32'hc40e7550, 32'hc1b4b480, 32'hc39a0a91},
  {32'h45036551, 32'hc35ef935, 32'h429e490c},
  {32'hc5118b4e, 32'hc380fba6, 32'hc3dd510f},
  {32'h439756b4, 32'hc3608abd, 32'h43391659},
  {32'hc3ee3147, 32'hc2c6b927, 32'hc3149309},
  {32'h44608884, 32'h429e22e9, 32'h43764833},
  {32'hc41ac1bc, 32'hc27a9c3c, 32'hc2d54386},
  {32'h448916d4, 32'h42115921, 32'hc3c4bc64},
  {32'hc4842c1d, 32'hc320e8cc, 32'hc25e1dee},
  {32'h446f5aa8, 32'hc33e4f7a, 32'hc2840040},
  {32'hc48548d6, 32'hc1d4d10d, 32'h40edefa8},
  {32'h45013ac2, 32'h3e177ad8, 32'hc1c7683e},
  {32'hc460d2ca, 32'hc3880f52, 32'h433de537},
  {32'h44f84e25, 32'hc309f618, 32'h44173c2f},
  {32'hc3aa2fb7, 32'hc34dd5ac, 32'h42857de8},
  {32'h42f12790, 32'h43335cb5, 32'h4349b722},
  {32'hc4bfa1f4, 32'h41f38920, 32'hc1a86e48},
  {32'h432abadf, 32'h41857ca2, 32'h43c94f19},
  {32'hc50e123e, 32'hc2364d0b, 32'hc3f523c8},
  {32'h450a4851, 32'hc316088c, 32'h425bbf39},
  {32'hc4c0fda2, 32'hc3138b1d, 32'h429fc45f},
  {32'h451cc48e, 32'hc32983c0, 32'h43033791},
  {32'hc4e0994a, 32'h428ee373, 32'h429c7c1e},
  {32'hc3a95788, 32'h4380696f, 32'hc3cb488b},
  {32'hc2d4b4e0, 32'hc1cf594a, 32'hc35403bc},
  {32'h4520789e, 32'hc103ffaa, 32'h43d9ed36},
  {32'h43eaefa2, 32'hc3a5c848, 32'h431993b9},
  {32'h437af0a6, 32'hc15f4bdd, 32'h427395bf},
  {32'hc4d3708a, 32'hc34b09a4, 32'h422d5f96},
  {32'h4486db63, 32'hc2d3fce2, 32'hc2e1b87e},
  {32'hc2b78fef, 32'hc3a5396b, 32'h435e7268},
  {32'h449c3c5c, 32'hc4004f44, 32'hc38f7102},
  {32'hc469df7c, 32'h4369521b, 32'hc3cd2f3b},
  {32'h4383290c, 32'hc3b63290, 32'hc3554d70},
  {32'hc511d2c0, 32'hc3086f11, 32'h42cd1c43},
  {32'h442b219a, 32'h441a37aa, 32'hc3e626e1},
  {32'hc4b5b2b9, 32'h43997d00, 32'hc3abd2ab},
  {32'h4514b0f1, 32'hc3ec4039, 32'h42057572},
  {32'hc40d5574, 32'h436a023d, 32'h437a6424},
  {32'h450502f6, 32'hc3a1639c, 32'hc346823f},
  {32'h433113e0, 32'h4302b8d3, 32'hc35c75ac},
  {32'h44a2c782, 32'h42fbe27c, 32'hc25e03c1},
  {32'hc405a010, 32'hc2c483fa, 32'hc2e92308},
  {32'h44d6c017, 32'h43b1d312, 32'hc32e7267},
  {32'hc4e8ca84, 32'hc353ff43, 32'h43398783},
  {32'h44fdce36, 32'hc31a588f, 32'h4207101c},
  {32'hc3ce3d27, 32'h43b053d3, 32'hc3b38b13},
  {32'h428ab72c, 32'h4383791b, 32'hc35861db},
  {32'hc4aa66a4, 32'hc3ba40dd, 32'hc26bdcdd},
  {32'h443d4d34, 32'h42a32276, 32'h424c3899},
  {32'h42dd7054, 32'hc3911a93, 32'hc38a4b6a},
  {32'h44a916c7, 32'h43a9825a, 32'hc2e669f9},
  {32'h43025f90, 32'hc3be8b47, 32'h43540856},
  {32'h45058698, 32'h434b34b2, 32'h42c20d9f},
  {32'h428f026a, 32'hc3210158, 32'hc2cf5d86},
  {32'h45070f76, 32'hc30be628, 32'hc31f2a02},
  {32'hc4957f16, 32'hc25d2c09, 32'h43a00438},
  {32'h44b9d236, 32'hc029a568, 32'hc36548f9},
  {32'hc2fdc180, 32'hc376ca77, 32'h43125738},
  {32'h43193c24, 32'h42e2f68f, 32'hc3dbd2d4},
  {32'h432f0ee0, 32'h43028604, 32'hc2d37b02},
  {32'h44089a56, 32'h431ae256, 32'hc3249cdb},
  {32'hc36f95c9, 32'hc3a9591c, 32'h43bfc5d6},
  {32'h4457a37b, 32'h421f3325, 32'hc3e83b8f},
  {32'hc49f3edf, 32'h43166755, 32'h4262013f},
  {32'h44b61715, 32'hc26ae014, 32'h42a0f37e},
  {32'hc51f2cd9, 32'hc306b5b6, 32'h405e1548},
  {32'h442a56e3, 32'hc377ab86, 32'h3fdc924c},
  {32'hc4f22a49, 32'hc237af8c, 32'hc381c9fa},
  {32'h44e43af4, 32'h4200a992, 32'hc33892f1},
  {32'hc289b740, 32'hc38c61ba, 32'h43ca0af2},
  {32'h44cf65b3, 32'hc27393fb, 32'hc21538b0},
  {32'hc33edba0, 32'h42bc6c8a, 32'h43436920},
  {32'h41ccfe00, 32'hc166ba3b, 32'hc325a062},
  {32'hc4cce031, 32'hc22242e1, 32'h439ec8fc},
  {32'h45021bde, 32'h419e576d, 32'h40ae6a1e},
  {32'hc50659cb, 32'h42615cb6, 32'h436e7cb7},
  {32'h43e6d1be, 32'hc3274151, 32'h42824f13},
  {32'hc502e92c, 32'hc3d53c3a, 32'hc307aa1d},
  {32'h4499f0a6, 32'hc1ea148d, 32'hc3e82d6a},
  {32'hc4d06d5a, 32'h4275f9c0, 32'hc3319652},
  {32'h45011d09, 32'hc34e822b, 32'hc3c43d83},
  {32'hc2fe1498, 32'h42c234fb, 32'hc312f956},
  {32'h4504b65d, 32'hc1a65d46, 32'hc3fac9d1},
  {32'hc4bff22a, 32'hc2c7f104, 32'hc24fd8fc},
  {32'h44a9d408, 32'h420ba78b, 32'h4267782a},
  {32'hc4a5402f, 32'h439f994d, 32'hc34c587b},
  {32'h44435038, 32'hc3ad2896, 32'h43b4832d},
  {32'hc3e47dc0, 32'hc190968f, 32'h437812c1},
  {32'h436a0e9c, 32'hc3767f19, 32'hc3284c5f},
  {32'h43833a10, 32'hc2f8ae1d, 32'hc34e3f7c},
  {32'hc51036bb, 32'h424c327d, 32'h42d9c7fa},
  {32'h447d44e4, 32'h42aa8be0, 32'hc395f8b0},
  {32'hc3b9b12c, 32'h4336719d, 32'h42221381},
  {32'h43a3bd94, 32'h43b6cdd7, 32'h4326fb8a},
  {32'hc39453a2, 32'h43065617, 32'h4313f6ee},
  {32'h44d28255, 32'h4320f716, 32'hc307bd59},
  {32'hc480f970, 32'h4300692f, 32'h42f41012},
  {32'h45015d34, 32'h42a34d76, 32'hc1ec7134},
  {32'hc4ad7f30, 32'hc331385b, 32'hc2efebba},
  {32'h450154c0, 32'hc2b70a5a, 32'hc2994aae},
  {32'hc5013ab0, 32'hc372b8c8, 32'h438c45fc},
  {32'h4444a3e6, 32'h43ef1251, 32'h44149155},
  {32'hc315dfd0, 32'hc40fcca8, 32'h427269c5},
  {32'h43a8f19c, 32'hc3aa5695, 32'hc3549816},
  {32'hc32f5d00, 32'h436f7669, 32'h42aa37dc},
  {32'h450be5b8, 32'h42f91e82, 32'h43388aab},
  {32'hc508e1fc, 32'h4215bb6c, 32'h43aaac62},
  {32'h451a4a8a, 32'hc2ac0409, 32'hc3015520},
  {32'hc18efed0, 32'h43898e23, 32'hc369f373},
  {32'h44dce1be, 32'hc382b057, 32'h428472f0},
  {32'hc4f08954, 32'hc1b47baa, 32'h43a1f52f},
  {32'h44f8dfb4, 32'h42fc679e, 32'hc3895ca9},
  {32'hc4905dd6, 32'h42c3cfe7, 32'hc12e9310},
  {32'h450e5a24, 32'h4287739f, 32'hc38efa65},
  {32'hc4990866, 32'hc38ce98b, 32'hc26cb13f},
  {32'h44caa0a9, 32'hc3812b00, 32'h42bb15bf},
  {32'hc490d6f3, 32'h421686db, 32'h4299f1a4},
  {32'h441fa1fa, 32'hc3450b82, 32'h433e8a22},
  {32'hc51e09af, 32'hc412179a, 32'h42614d76},
  {32'h450c78a8, 32'h4429489c, 32'h43afbf15},
  {32'hc4e679ba, 32'h4157e259, 32'h4397de02},
  {32'h42396610, 32'hc3812292, 32'hc32b4b2f},
  {32'hc1dda2da, 32'hc26102f3, 32'hc37c6128},
  {32'h449d4787, 32'h4338315f, 32'hc3691fe7},
  {32'hc50d456e, 32'hc3a3c0fe, 32'h4338f2e9},
  {32'h44f2d52d, 32'h431c2e77, 32'h438a480d},
  {32'hc34496a8, 32'hc3019739, 32'h43071003},
  {32'h44ebf8a7, 32'h4285179b, 32'hc0b8f673},
  {32'hc4d78133, 32'hc02cfad4, 32'hc10ab7f3},
  {32'hc1a2b4c0, 32'hc23ee8c9, 32'hc2da82df},
  {32'hc3b2e2ca, 32'h4372bf89, 32'hc3deb581},
  {32'hc2734500, 32'hc2748cec, 32'hc3a08791},
  {32'hc344bc58, 32'hc28858be, 32'hc395a720},
  {32'h44b71ccc, 32'h42248e0b, 32'hc21b1baa},
  {32'hc38cbb82, 32'h435cf499, 32'h431d069d},
  {32'h44e12748, 32'hc24a60e2, 32'hc2ba0b96},
  {32'hc4b1b88d, 32'h41442bf6, 32'hc2013736},
  {32'h44fd86dd, 32'hc3e07902, 32'hc33d3f03},
  {32'hc440e77e, 32'hc28aa1ca, 32'hc345b854},
  {32'h43719b86, 32'hc402edf3, 32'h432d7a0b},
  {32'hc500a334, 32'h438172fc, 32'h422447d0},
  {32'h4516c8c9, 32'hc26d438e, 32'h42529ec8},
  {32'hc3e289f0, 32'h4203a83d, 32'h42b8b822},
  {32'h45099a8d, 32'h43636b3a, 32'h436b4cff},
  {32'hc4b50586, 32'h436bdaae, 32'hc2464978},
  {32'h44859232, 32'hc29f4672, 32'hc345ee7c},
  {32'hc4f2ddd7, 32'h420956ae, 32'hc2e2028f},
  {32'h44c1c75c, 32'h430cf4eb, 32'h429779b3},
  {32'hc3c12a8b, 32'hc30dde82, 32'hc3663e54},
  {32'hc0c40e80, 32'hc2565282, 32'hc201a3b0},
  {32'hc45f93d6, 32'hc2b1c67f, 32'h41b2b513},
  {32'h4417357a, 32'h42a41aea, 32'hc3bdabaf},
  {32'hc49ca062, 32'hc31a3283, 32'h4229d44a},
  {32'h4400aac8, 32'h43cf4d01, 32'hc3a4d226},
  {32'hc4cbd1e1, 32'h4249e41e, 32'hc30881c4},
  {32'h441db8f0, 32'h41586a14, 32'h43896ae6},
  {32'hc50679e2, 32'hc00a253c, 32'h42ea435c},
  {32'h44875584, 32'h42d9e116, 32'h438cb3b8},
  {32'hc4f13418, 32'h4360cbec, 32'h4308583e},
  {32'h4506029d, 32'h4399aa31, 32'hc314446d},
  {32'hc487bc49, 32'h42f4b024, 32'hc38ba612},
  {32'h44d9da4e, 32'h433f67f0, 32'hc3e00895},
  {32'hc4a1be46, 32'hc2b5d5f3, 32'h43ccd8ab},
  {32'h44e54854, 32'h41796346, 32'h4363d9f1},
  {32'hc390f5a5, 32'hc3209e0c, 32'h4365cacc},
  {32'h449c0660, 32'h42d5c226, 32'h430289f6},
  {32'hc3668c88, 32'h41dc09bb, 32'hc3b02fc1},
  {32'h4524c417, 32'h435159b2, 32'h4409ffbf},
  {32'hc3f1943d, 32'hc2cf08b0, 32'h4355e256},
  {32'h44d5a5ce, 32'h43b929d7, 32'h436406a9},
  {32'hc4e8f1ba, 32'hc351ed22, 32'hc339fe08},
  {32'h44eb16a4, 32'h43054275, 32'h439ac851},
  {32'hc4f56ee8, 32'hc40acedc, 32'h422f6122},
  {32'h43deed56, 32'h437b6067, 32'h431ca2e5},
  {32'hc3cdbd3e, 32'h42b57738, 32'h41ade8aa},
  {32'h44ea2369, 32'hc12dd862, 32'h435337a8},
  {32'hc3258359, 32'h421016ab, 32'h43d8889b},
  {32'h44105085, 32'h438c9a1d, 32'h4348ea11},
  {32'hc51050b8, 32'h4309e9b5, 32'hc3917e09},
  {32'h44996aba, 32'h4294e622, 32'h403ffa98},
  {32'hc517a08a, 32'h40a9acee, 32'hc3dcf83c},
  {32'h4462592e, 32'hc3b66d56, 32'h40d6acca},
  {32'hc5174322, 32'hc16a72d7, 32'h43c5ba6e},
  {32'h444d4985, 32'h439f2a8f, 32'h424cacd5},
  {32'hc4ecc0dd, 32'hc38a51bd, 32'hc35be36a},
  {32'h44cc7ed2, 32'hc3ac7e40, 32'hc385ed0f},
  {32'h41904300, 32'hc3814632, 32'hc30239a7},
  {32'h4518864c, 32'hc2830c12, 32'hc3eb664b},
  {32'hc2f6e720, 32'h40c68e74, 32'hc39e2512},
  {32'h44e17501, 32'hc21720cc, 32'h41845f0d},
  {32'hc474b4a7, 32'hc2ab0066, 32'h4296210b},
  {32'h44958025, 32'h43edea10, 32'h43bb36bc},
  {32'hc50ed34f, 32'hc32e231d, 32'hc13772c4},
  {32'h44995dbb, 32'h4382cb15, 32'hc122e783},
  {32'hc4d4ec81, 32'h43ce798c, 32'hc377810f},
  {32'h4186cdcc, 32'h439dcba3, 32'h434cebf8},
  {32'hc5258cac, 32'h42694805, 32'hc331b08a},
  {32'h4504b757, 32'hc3e382c1, 32'h43baf6c9},
  {32'hc40033f0, 32'hbe4ac720, 32'h42b07e7e},
  {32'h442c318d, 32'h42a4720a, 32'hc3447853},
  {32'hc4ad542d, 32'hc395c406, 32'hc0a017d5},
  {32'h43c8a490, 32'hc3312cb4, 32'hc3f95418},
  {32'hc4307cdd, 32'hc306e881, 32'h429f4624},
  {32'h45052247, 32'hc00bb0e0, 32'h422333b7},
  {32'hc41a1244, 32'h42d4877d, 32'h42df0a7e},
  {32'h44aa5881, 32'h43a81ed8, 32'hc36d2df8},
  {32'hc4ecd343, 32'hc390861d, 32'hc3680f47},
  {32'h44b451ae, 32'h43c44ada, 32'h439ffea0},
  {32'hc4036866, 32'h430861a0, 32'h428294ca},
  {32'h45018edc, 32'hc3a1656e, 32'h438bebd4},
  {32'hc5100748, 32'h412f0d6b, 32'hc32f29da},
  {32'h4429a6f0, 32'hc3290a6b, 32'h4397ae7e},
  {32'h43b0f247, 32'hc3614232, 32'hc2048866},
  {32'h44b421fd, 32'h4221ab74, 32'hc3887620},
  {32'hc4c31435, 32'h425ce2c3, 32'h43449736},
  {32'hc2e1bb40, 32'h40bea976, 32'h438efe36},
  {32'h4285e509, 32'h43383e1a, 32'h41c61669},
  {32'h435b1dcf, 32'h42ad74e1, 32'hc26097ec},
  {32'hc3c9be18, 32'hc2fa8f8a, 32'h42b3b649},
  {32'h44db38ff, 32'hc1fb29b6, 32'hc29b03e9},
  {32'hc4f54c0b, 32'hc227d627, 32'hc2a49ba3},
  {32'h450da748, 32'hc22c7731, 32'h435288b5},
  {32'hc499f058, 32'hc23c4efd, 32'h439202ee},
  {32'h44ea1639, 32'h43216e7a, 32'h4428a8e8},
  {32'hc3248610, 32'hc31e1a2e, 32'h42198e26},
  {32'h43b2a43c, 32'h439f9598, 32'h42418b64},
  {32'hc4161533, 32'h43cdd0b8, 32'h424613a2},
  {32'h4519291a, 32'hc332993e, 32'hc3728ea8},
  {32'hc39e117c, 32'hc38abb1c, 32'h42c636ba},
  {32'h43a1de20, 32'hc1ca5f18, 32'h42bed050},
  {32'hc49683a8, 32'h420e1e07, 32'hc2a88db5},
  {32'h44f54f0c, 32'h42f026a9, 32'h43665ddb},
  {32'hc4ff61bb, 32'hc306a3c6, 32'hc3bf350a},
  {32'h43adc066, 32'h4138d573, 32'hc38675ae},
  {32'hc39f3d4c, 32'hc313ec4f, 32'h437772cd},
  {32'h44c92224, 32'hc3bd2f34, 32'h43a8313b},
  {32'hc44b7a4a, 32'hc39354d2, 32'hc379e031},
  {32'h44404664, 32'h4242b8b0, 32'h42a73b11},
  {32'hc46d9504, 32'h438b906d, 32'hc3b83888},
  {32'h44e64a5f, 32'h42f79ea9, 32'h40570ba3},
  {32'hc4663de6, 32'h43c6c5c7, 32'h42c37080},
  {32'h4499ad8f, 32'h440512a0, 32'hc237eea3},
  {32'h43865a5b, 32'hc363768d, 32'hc2e645c1},
  {32'h44170c1a, 32'h43312c04, 32'hc28015bc},
  {32'hc4ca8812, 32'hc3327093, 32'hc30b35e9},
  {32'h4453411c, 32'h42a40f84, 32'hc34457d6},
  {32'hc4271456, 32'hc3c0c0b9, 32'hc3a26a66},
  {32'h44f86a54, 32'h427bbc20, 32'h43bb207f},
  {32'hc4d470f8, 32'h43744a22, 32'h440b6e19},
  {32'h43ac3fdc, 32'h423e22be, 32'h4370b3e7},
  {32'h438cef58, 32'h43335c46, 32'hc359d0fc},
  {32'h4408d692, 32'h426e8bfc, 32'h40c6930a},
  {32'hc3b49ee0, 32'h439425ac, 32'h43b21d1f},
  {32'h4432477c, 32'h4335140f, 32'h435ca11b},
  {32'hc383dff6, 32'h434f7772, 32'h438523a2},
  {32'h442c01f9, 32'hc2d2cd77, 32'hc32d96ae},
  {32'hc4bea44e, 32'hc1d9cb42, 32'h43115515},
  {32'h43dce18c, 32'hc179dfef, 32'h43548c5f},
  {32'hc4bb49f5, 32'hc3433200, 32'h43218166},
  {32'h45090276, 32'h438b03fc, 32'hc3a2219c},
  {32'hc4b7996f, 32'hc3162802, 32'h41c07170},
  {32'h450f5548, 32'hc2b0732a, 32'h402bc10e},
  {32'hc4b7610a, 32'hc3379b9a, 32'hc1fc32e4},
  {32'h44bb93ea, 32'hc2099582, 32'hc1a5375f},
  {32'hc4c5590c, 32'hc24dbe74, 32'hc2c307e9},
  {32'h448d2664, 32'h44034380, 32'h42b7e142},
  {32'hc4c3ceb8, 32'h4412c773, 32'hc3061e3f},
  {32'h44edea90, 32'h438043e1, 32'h43b25dfb},
  {32'hc4cffaea, 32'hc3385f1b, 32'hc339a598},
  {32'h450489ef, 32'hc142e008, 32'h432b8319},
  {32'hc46f7bdc, 32'h426f6466, 32'h422a2023},
  {32'h43a93078, 32'hc3bd3dc4, 32'h4277739c},
  {32'hc36462b6, 32'hc185a832, 32'hc2fbb94b},
  {32'h44b4f7c6, 32'hc3b8e4de, 32'h4133b44c},
  {32'hc4ef1b5a, 32'hc35021ef, 32'hc2aa69c6},
  {32'h449412ec, 32'hc2222822, 32'hc1c913e6},
  {32'hc490b76f, 32'h431b5a11, 32'hc35b914a},
  {32'h44fd2015, 32'h4056286d, 32'h4335e557},
  {32'hc4d139e0, 32'hc3a46ed6, 32'hc4229427},
  {32'h450aff6c, 32'h4400548e, 32'h41b245f9},
  {32'hc48d9ec3, 32'h40fe7737, 32'hc2420d70},
  {32'h452736d6, 32'hc32cf553, 32'h43acd49a},
  {32'hc36e52d8, 32'hc3b7e29c, 32'hc2162a1d},
  {32'h4333e8f0, 32'h42bde0a1, 32'hc2ba071e},
  {32'hc4113df7, 32'h42996997, 32'h4392c70a},
  {32'h4476636c, 32'hc397f3d9, 32'hc2994697},
  {32'hc47de00f, 32'h41b1436f, 32'h42a7a585},
  {32'h44c52065, 32'h417fd8e2, 32'h432bb8c9},
  {32'hc401a0e5, 32'hc3b0aadf, 32'hc35dd616},
  {32'h4362091d, 32'h429876a3, 32'h4283f254},
  {32'hc4e4552f, 32'h3fcac239, 32'hc3849f6f},
  {32'h44a424b2, 32'hc2c45b9d, 32'hc0e09de2},
  {32'hc4c87411, 32'h417da309, 32'h42b146a0},
  {32'h44f65aea, 32'hc3e32922, 32'h41d3b5a9},
  {32'hc4399e10, 32'h4348f362, 32'hc3b14e5a},
  {32'h450d4a2f, 32'h4412edaa, 32'h43167c2e},
  {32'hc4da0a97, 32'hc35a26c3, 32'h42abb0c8},
  {32'h44a262f4, 32'h42d787d9, 32'h426c2542},
  {32'hc471d95e, 32'hc39a5829, 32'h439bf8f1},
  {32'h4509f436, 32'h42c50b41, 32'h4372f39d},
  {32'hc44c81ab, 32'hc31d0c5f, 32'hc1982ad1},
  {32'h44d55c5e, 32'hc1936fa1, 32'h43b61b94},
  {32'hc511a5d0, 32'hc266c553, 32'hc1e56d7a},
  {32'h4483166f, 32'hc30974d4, 32'h43a3c287},
  {32'hc4c702f8, 32'hc217f842, 32'h425f4e11},
  {32'h4207e312, 32'h4250fb46, 32'h4016cb0d},
  {32'hc477906c, 32'hc3178d54, 32'h4113eb5e},
  {32'h449b375a, 32'hc2f6b0f2, 32'hc39b54e3},
  {32'hc4a1d282, 32'hc315273c, 32'h42df6fee},
  {32'h44fcfd06, 32'hc27f381f, 32'hc0babe2f},
  {32'hc4fe8a2d, 32'hc3e87161, 32'h40fe51dd},
  {32'h444504fa, 32'h42894edc, 32'hc30fa0a9},
  {32'hc4ab0ef0, 32'hc34de428, 32'hc164eeca},
  {32'h43b46af1, 32'h4247d1c3, 32'h4333a9e9},
  {32'hc44f2d90, 32'hc30875ac, 32'h43c89879},
  {32'h43fe35ec, 32'h42f12baf, 32'hc392f8e2},
  {32'hc419e9db, 32'hc29e606f, 32'h42dc5db3},
  {32'h44d618c9, 32'hc31754c9, 32'h4181757f},
  {32'hc499afed, 32'hc33f63eb, 32'h43c12fe1},
  {32'h44486f00, 32'h4384b5ca, 32'h420616ed},
  {32'hc395037d, 32'hc31f420e, 32'hc2adad04},
  {32'h443443d0, 32'hc3606112, 32'h431d6274},
  {32'hc42e47e2, 32'hc30fe4db, 32'hc30fa4a8},
  {32'h45148001, 32'h425e9a7f, 32'hc2ac9ff9},
  {32'hc4561c42, 32'h439c8418, 32'h43237578},
  {32'h41732280, 32'hc2ea5146, 32'hc31edbe6},
  {32'hc3eb1544, 32'h439e2db2, 32'hc3524db0},
  {32'h4507029f, 32'hc33e8da0, 32'hc2c6c375},
  {32'hc395a514, 32'h4250e9c5, 32'hc2dcdf44},
  {32'h4510aa0a, 32'h42f47db4, 32'hc316ed8a},
  {32'hc4315964, 32'h432c144e, 32'h43cdb9e0},
  {32'h4458df2c, 32'hc2fda393, 32'h43466456},
  {32'hc502684e, 32'hc32cf27e, 32'hc432d921},
  {32'h44ae7960, 32'hc39f5b96, 32'h4320c0a8},
  {32'hc313fb00, 32'hc2d7b511, 32'h43b718b8},
  {32'h451cb0d0, 32'hc188fb30, 32'hc39c629a},
  {32'hc4808d10, 32'h41763f65, 32'hc2b3fa79},
  {32'h43212200, 32'h43ce6f80, 32'h4390bc3b},
  {32'h40c12c40, 32'hc2f78e1f, 32'hc34165c6},
  {32'h4401db04, 32'h42d0a474, 32'hc31b3d6e},
  {32'hc2c7a488, 32'hc2fe05c9, 32'h43428688},
  {32'h44e8b692, 32'hc14c2e51, 32'h4367679a},
  {32'hc4ef1106, 32'hc18f131d, 32'hc396339b},
  {32'h4305f7a1, 32'hc1027a51, 32'h4182eb74},
  {32'hc47ff3c8, 32'h431a3b19, 32'hc2f171c4},
  {32'h42382a20, 32'hc392202a, 32'hc39ff536},
  {32'hc5074224, 32'h434527af, 32'h43eb826e},
  {32'h4525cf98, 32'h43d54dc9, 32'h430a8be8},
  {32'hc4665f17, 32'h42e259a5, 32'h43dbf8db},
  {32'h451573ae, 32'hc235d3ff, 32'h43c6cbb4},
  {32'hc47d41a9, 32'h43783cf2, 32'h429a3357},
  {32'h439353e4, 32'hc38c43f9, 32'h42b856e4},
  {32'hc4e02add, 32'hc33a23cd, 32'h4224e6c1},
  {32'h4429dce2, 32'h43789bc6, 32'hc2a43f18},
  {32'hc4bf35c6, 32'h44433635, 32'h419ff487},
  {32'h43941b88, 32'h42bc18b5, 32'hc429ca8c},
  {32'hc4a4ad36, 32'hc24555f1, 32'hc297f079},
  {32'h43c98111, 32'h43547a51, 32'hc2bcf348},
  {32'hc4bff915, 32'h42f4245b, 32'h439dc425},
  {32'h437354ad, 32'hc2c8be57, 32'h42f92be4},
  {32'hc458085e, 32'hc380b9b1, 32'hc33f1abb},
  {32'h44d0adfd, 32'h43a56621, 32'hc29bb8e0},
  {32'hc430e1c6, 32'hc1affc5c, 32'h43ce3ccc},
  {32'h44d4d5a0, 32'h43b11260, 32'hc25535ec},
  {32'hc3e08fa9, 32'hc298fdb9, 32'h4359718f},
  {32'h439a5741, 32'hc376121b, 32'hc3609dec},
  {32'hc4c3a9fc, 32'h42de7f3a, 32'hc2967706},
  {32'h44eb33aa, 32'hc39c0e83, 32'hc21ed614},
  {32'hc4e83f6c, 32'hc36b4791, 32'h43f574bd},
  {32'h44421dc6, 32'hc28d9c9d, 32'hc337f3d2},
  {32'hc4cc3336, 32'hc3936f24, 32'h42bb46bb},
  {32'h4500be5d, 32'hc34d43b5, 32'h43137db2},
  {32'hc4c8bacc, 32'hc311fd1d, 32'hc225dc83},
  {32'h44caf7b7, 32'hc231979d, 32'hc425836a},
  {32'hc3bf7cb0, 32'h422bc9ea, 32'hc1e8e016},
  {32'h450205b7, 32'h4281f8dd, 32'h4370a4ed},
  {32'hc4fc8f00, 32'hc35b8f02, 32'h43bd19ab},
  {32'h44fecae0, 32'h430d5504, 32'h41c10734},
  {32'hc485ed62, 32'h433ddbf6, 32'h435614b0},
  {32'h442392ba, 32'h420a43dd, 32'hc285dd24},
  {32'hc18ac908, 32'h435fc054, 32'h430e3267},
  {32'h44f90c16, 32'hc3c34a32, 32'hc1d6bc9f},
  {32'hc488f55e, 32'h43bf44be, 32'h429bb1f4},
  {32'h45009732, 32'h4340181f, 32'h430ab448},
  {32'hc4eec870, 32'hc2abc87f, 32'hc390c530},
  {32'h44d8c854, 32'h436196fa, 32'hc269d639},
  {32'hc3aaefaf, 32'h42983624, 32'h43be4488},
  {32'h4474c0a0, 32'h42ed1d9c, 32'hc2c2e22a},
  {32'hc3f18344, 32'h44097dd4, 32'h43c006d0},
  {32'h44bcc740, 32'h42abee0c, 32'h43103769},
  {32'hc515328b, 32'h427126ae, 32'hc22282f3},
  {32'h44d01af7, 32'h42f68bc4, 32'h42b5cf3a},
  {32'hc4714e00, 32'hc1a124f9, 32'hc147e20a},
  {32'h445634e8, 32'hc3813a63, 32'hc368486d},
  {32'hc4c33132, 32'h43b2f956, 32'h4283f60c},
  {32'h44d0b7c4, 32'hc35d5043, 32'hc30707a9},
  {32'hc4d6cffa, 32'hc28a38f4, 32'h4298d237},
  {32'h44e2037a, 32'h431b70dd, 32'hc3851898},
  {32'hc42cf694, 32'hc371d162, 32'h438c98ad},
  {32'h442a679e, 32'h432a0b31, 32'h40d492a0},
  {32'hc50fed40, 32'h418a9cd7, 32'h43593876},
  {32'h448c5b0c, 32'hc415d42d, 32'hc3f97eea},
  {32'h42ea9b60, 32'hc2d9fe1c, 32'h41ac4b3a},
  {32'h4496a733, 32'hc2b1b3b7, 32'hc2869e09},
  {32'h44cd600d, 32'h42b8fdfa, 32'hc033a1e6},
  {32'hc50b6c7a, 32'h413c0f6c, 32'h429ba924},
  {32'h43a11524, 32'hc426bee8, 32'hc2c78c28},
  {32'hc4e74789, 32'hc307aa8c, 32'hc318097d},
  {32'h43855c25, 32'h43e8793c, 32'h43261647},
  {32'h42c698c2, 32'hc31a5bf3, 32'h42c71c93},
  {32'h442d0f28, 32'hc26bf982, 32'hc3de2af7},
  {32'hc3d30144, 32'h434f440d, 32'h43080697},
  {32'h4480abc0, 32'h431c2f31, 32'h418d2041},
  {32'hc3c1928c, 32'hc397e165, 32'h4387997b},
  {32'h44b72877, 32'h43017dfc, 32'hc1cbf48a},
  {32'hc4e65a78, 32'hc3149c4f, 32'h430ed5ea},
  {32'h440e4d98, 32'h430059e5, 32'h41935820},
  {32'hc4dcd81d, 32'h43ed97df, 32'hbfac8ff0},
  {32'h44a80b1a, 32'hc335f151, 32'hc0af8288},
  {32'hc31b9950, 32'h3f1dc9c8, 32'h431a0bf3},
  {32'h44bfd37e, 32'h438bd8d8, 32'hc3fae7b7},
  {32'hc47a17a4, 32'h42b33a69, 32'h4304e020},
  {32'h4512f45b, 32'hc39bc77e, 32'hc389fe1d},
  {32'hc3a5d957, 32'h42c8319f, 32'h41a13275},
  {32'h44e9c290, 32'h435f2c58, 32'h4251043a},
  {32'hc4d304d4, 32'hc274e0fb, 32'hc293a76a},
  {32'h44ef3df7, 32'h43447303, 32'hc321ecc9},
  {32'hc3210d10, 32'h4224e756, 32'hc0739c08},
  {32'h4496c6c0, 32'h420a5032, 32'hc3a1f0d3},
  {32'hc4bedf15, 32'hc28f1b85, 32'h42b218f4},
  {32'h442a8028, 32'h41f80649, 32'h42d1e93d},
  {32'hc3845a80, 32'hc34fd888, 32'hc2e9f996},
  {32'h44dab7a3, 32'hc2048152, 32'hc324d7fa},
  {32'hc4c8ca5a, 32'hc2e6efe4, 32'hc281125d},
  {32'h44a147f2, 32'hc296fc47, 32'hc35cea61},
  {32'hc3e6ebd8, 32'h4264ee4c, 32'h4281d4c7},
  {32'h42775df0, 32'hc353f566, 32'hc2e2045a},
  {32'hc312b58a, 32'hc36d72f9, 32'hc22b6442},
  {32'h44a1fb7e, 32'h4318e720, 32'hc329c386},
  {32'hc4dec55b, 32'h429ae3e9, 32'h4294614b},
  {32'h44b3c0c3, 32'hc2578d2a, 32'hc3818453},
  {32'hc50196ed, 32'hc31aaf57, 32'h43ba45e7},
  {32'h44a4a86a, 32'hc33ad41e, 32'h43b8765b},
  {32'hc4c3a86c, 32'hc3ab9b77, 32'h40c16e71},
  {32'h448c7298, 32'hc3624e35, 32'hc322d4ce},
  {32'hc4334b4e, 32'h43b30fb9, 32'h438a377c},
  {32'h450c290c, 32'h42f9c418, 32'hc3715b4d},
  {32'hc4fc0077, 32'h4220fb8c, 32'hc222428e},
  {32'h4519cde2, 32'h43094fe0, 32'h423be75b},
  {32'hc4d74fa0, 32'h430867a3, 32'h4300f872},
  {32'h4520ad72, 32'hc2364ab4, 32'hc15efce1},
  {32'hc4a70cc7, 32'h4361a4ae, 32'h43ec5b7f},
  {32'h44dceb9f, 32'h4390967e, 32'hc3a59d7b},
  {32'hc4453918, 32'h4295af79, 32'hc35b2382},
  {32'h4512e2d7, 32'hc39c3bb4, 32'h42d42c29},
  {32'hc4bd3475, 32'hc3d0576f, 32'hc1946765},
  {32'h4485d420, 32'h43ae411d, 32'hc2fb5e68},
  {32'hc49b72fa, 32'h426ad464, 32'h43b8e9ee},
  {32'h44b814d7, 32'hc2e352db, 32'hc21cb6c3},
  {32'hc50030d4, 32'h430140b5, 32'h433fba7a},
  {32'h42d10af0, 32'h438fde22, 32'h437b009b},
  {32'hc5066b79, 32'h43c65d00, 32'hc3d21ce2},
  {32'h4449954e, 32'h4369ecbf, 32'h43e616f8},
  {32'hc49cd51c, 32'hc34bda45, 32'hc2c0400a},
  {32'h44965f3a, 32'hc33804c0, 32'hc34682b8},
  {32'hc1be8020, 32'hc2b75246, 32'hc219330c},
  {32'h450a6957, 32'hc31e73cd, 32'hc298f145},
  {32'hc4a3e714, 32'h431e6b22, 32'h42e28c94},
  {32'h450463f7, 32'h4320ca64, 32'h43466ae0},
  {32'hc3bcafe8, 32'hc406f48e, 32'h4418eef3},
  {32'h43b7a1c0, 32'h428640d3, 32'hc3c8b523},
  {32'hc447685c, 32'hc36e3018, 32'hc32ff025},
  {32'h43a1b992, 32'hc3577323, 32'h42959292},
  {32'hc39573b0, 32'h42e04eb1, 32'h440549b8},
  {32'h43f4c3bc, 32'hc29ef6d7, 32'h42a2d748},
  {32'hc41d9e67, 32'hc31b5f7a, 32'h41d0554c},
  {32'h44c61572, 32'hc2aae03c, 32'h4392b309},
  {32'hc4a4d443, 32'h4223799f, 32'h43738c53},
  {32'h44e816aa, 32'hc2a8245d, 32'h41f45738},
  {32'hc4edf288, 32'hc2f2d588, 32'hc34ebf1f},
  {32'h44b861f7, 32'h4347a712, 32'hc378cd07},
  {32'hc4b6ada3, 32'hc194ac18, 32'hc2fd97c5},
  {32'h4517451d, 32'h428b4a70, 32'h43e5bf09},
  {32'hc4c5295c, 32'h4231c4b4, 32'h4308bafa},
  {32'h4439aab0, 32'hc344e44e, 32'h42b16202},
  {32'hc4de2581, 32'h4102b9e4, 32'h428870ef},
  {32'h43b3024e, 32'h437f73b1, 32'h431826f3},
  {32'h42c23ae0, 32'h4336541d, 32'h438d781d},
  {32'h449152d7, 32'hc2a22570, 32'hc00c5fac},
  {32'hc4cf806f, 32'h412508ee, 32'h42502189},
  {32'h4502fbaf, 32'hc3cc65d2, 32'h42a3d0f1},
  {32'hc4863d95, 32'hc3c64de2, 32'hc273d0f3},
  {32'h441d408e, 32'hc38ef573, 32'h43563855},
  {32'hc4d0aee2, 32'hc380c354, 32'hc39b637b},
  {32'h441a60ec, 32'hc202c939, 32'hc380363e},
  {32'hc515a996, 32'hc326e5cf, 32'h440f5145},
  {32'h44855034, 32'h4390553a, 32'hc38410e4},
  {32'hc50e4e68, 32'hc37f82fc, 32'h42e0b806},
  {32'h44e988cd, 32'h431b4567, 32'h43ecfec1},
  {32'hc4964bc2, 32'hc3092378, 32'h4345b5d0},
  {32'h44398416, 32'h43c2dbcd, 32'h4307a372},
  {32'hc4f11128, 32'h417ee7b5, 32'hc3810225},
  {32'h44d24e4d, 32'h438e4025, 32'hc3cd5c0f},
  {32'hc4995163, 32'h43a34b01, 32'h43ddbf4c},
  {32'h421b4488, 32'hc2afbbb0, 32'hc3c4d715},
  {32'hc4c275f4, 32'hc351c6ac, 32'h43af7572},
  {32'h44bae2d5, 32'hc3bbd1d8, 32'h42da9ce3},
  {32'hc410ed88, 32'h439b6333, 32'h439b45bf},
  {32'h44b44f0a, 32'hc2dadd29, 32'h4347d125},
  {32'hc343eb00, 32'hc39e0430, 32'hc3467b00},
  {32'h44c0ca4f, 32'hc317ceb9, 32'hc2bd770f},
  {32'hc50474a0, 32'h4258972b, 32'hc37cb9ee},
  {32'h44c331bf, 32'hc318d67e, 32'hc3876cc3},
  {32'hc3622550, 32'h423881f0, 32'hc3c6bc04},
  {32'h43e3b864, 32'hc24b70fd, 32'hc3c7a122},
  {32'hc3d8bbea, 32'hc25d1021, 32'h42cffd50},
  {32'h41f05cc0, 32'hc2b483d0, 32'h439daca2},
  {32'hc4223f72, 32'hc3cee1ab, 32'h43ad6dd9},
  {32'h43ad959a, 32'h41772202, 32'h42f68c89},
  {32'hc4866c97, 32'hc08f5268, 32'h431bf712},
  {32'h4510f491, 32'hc3965290, 32'h4367406e},
  {32'hc4320575, 32'h43c9a9d6, 32'hc40664ed},
  {32'h44ce5e88, 32'h43ca3926, 32'h42a23f26},
  {32'hc501f32d, 32'h41e78446, 32'h428a1731},
  {32'h43fbea22, 32'hc2c5a099, 32'hc39843fa},
  {32'hc365172c, 32'hc301ac58, 32'hc2d5ed97},
  {32'h450f1b87, 32'hc09501ee, 32'h42c706de},
  {32'hc47ebbd7, 32'hc31a2a84, 32'hc336c848},
  {32'h44944ad8, 32'hc31bde05, 32'hc29c4407},
  {32'hc461f363, 32'hc31afce6, 32'h4330e5ee},
  {32'h43c60e06, 32'h44087aa9, 32'h42ebea78},
  {32'hc3c1a191, 32'h440f9c78, 32'h41c9d35f},
  {32'h448d5147, 32'hc386ba73, 32'h42fd847b},
  {32'hc480d77e, 32'h4307c624, 32'h40482ee8},
  {32'h44502086, 32'hc279c3b1, 32'h438a7d47},
  {32'hc4db0005, 32'hc37c5ad9, 32'h4313b9ed},
  {32'h450117af, 32'h4245bae7, 32'hc2b5cc96},
  {32'hc5081676, 32'h43c728aa, 32'h41b7d307},
  {32'h450b160b, 32'hc3aa4c62, 32'hc3b0ac78},
  {32'hc496187b, 32'h41771afc, 32'h42dcf7f5},
  {32'h446fcef2, 32'hc15a4468, 32'hc34d1cce},
  {32'hc4f186a4, 32'hc39bceaa, 32'hc30d936b},
  {32'h44d21e29, 32'h434536a3, 32'hc4016231},
  {32'hc40f6b68, 32'hc34fc843, 32'hc31c9213},
  {32'h40c6b300, 32'hc2411200, 32'h430c35ad},
  {32'hc4aaeacd, 32'hc2cffd00, 32'hc3367d3e},
  {32'h441d816a, 32'hc2c7811f, 32'h421ef418},
  {32'hc4e90120, 32'hc2a7f9d7, 32'h43eed93a},
  {32'h4510567c, 32'hc2275171, 32'h43314730},
  {32'hc482c5c8, 32'hc2231156, 32'hc2d12d6e},
  {32'h4332f4d8, 32'hc2be5b7d, 32'hc3335a7a},
  {32'hc47b3e1d, 32'h42a408a2, 32'hc38016fe},
  {32'h4369679f, 32'hc2be47b4, 32'h42d3d14a},
  {32'hc469938a, 32'h4378fac0, 32'h439ecfff},
  {32'h448194fc, 32'hc2e588ec, 32'hc1248e4e},
  {32'h41676a7e, 32'h42980792, 32'h4368e446},
  {32'h450b95f2, 32'hc368f514, 32'hc3452546},
  {32'hc4920955, 32'hc393f3bc, 32'h433ae6d7},
  {32'h44a71254, 32'h42e4004c, 32'hc33e6f6a},
  {32'h43c083f6, 32'hc234f6cc, 32'h437ffbb2},
  {32'h438c907c, 32'hc2af44a0, 32'h42988515},
  {32'hc468b220, 32'h43a1fb55, 32'h42e88d98},
  {32'h4501cdd7, 32'hc3c52aaf, 32'hc42767a0},
  {32'hc5121e3f, 32'hc3a6d1ed, 32'h43d5cb66},
  {32'hc2fbe320, 32'hc4021179, 32'h42a899ac},
  {32'hc4d48d18, 32'hc350b1c2, 32'h42a7b3d8},
  {32'h448a56e2, 32'hc32bd5cb, 32'hc3a8b0e5},
  {32'hc5177328, 32'hc2b31ef1, 32'hc2344dda},
  {32'h450ae549, 32'h433d4537, 32'h42cd70e2},
  {32'hc4ea6b2e, 32'h436aa7f8, 32'hc0a9ec46},
  {32'h4503faa0, 32'hc3bf057d, 32'hc30f2de9},
  {32'hc4be7662, 32'hc33a3f60, 32'hc344d923},
  {32'h43601796, 32'h4390cbae, 32'hc3468bbc},
  {32'hc449127c, 32'hc373c727, 32'h4385c8df},
  {32'h450e9af4, 32'hc3824bca, 32'h42d6af9f},
  {32'hc4caabca, 32'hc23552d0, 32'h43423ffc},
  {32'h44974662, 32'hc33c276e, 32'h430b3f87},
  {32'hc4daf4d2, 32'h431427fe, 32'hc3868e68},
  {32'h4382417e, 32'h43badbc7, 32'h41dfa106},
  {32'hc3531776, 32'h4380e095, 32'hc38a1baa},
  {32'h44972ee4, 32'hc25e5a3a, 32'hc3a2d774},
  {32'hc5181310, 32'hc29fb17e, 32'h3f0ca7ba},
  {32'h44458fd9, 32'hc33c094c, 32'h42892189},
  {32'hc49fa839, 32'h40bc7e41, 32'h426ffdc2},
  {32'h450d1b69, 32'hc2b2b707, 32'hc2046a0f},
  {32'hc4d441ed, 32'h4266d11a, 32'h42c3eb67},
  {32'h450409dd, 32'h43a6a6ce, 32'h43c28a66},
  {32'hc4f07058, 32'hc35547b9, 32'hc1fe46ec},
  {32'h4454ef10, 32'hc3c8a472, 32'h4389155e},
  {32'hc4f40aea, 32'h43bf5a06, 32'hc30b6115},
  {32'h44cfe4ca, 32'hc2c45152, 32'hc324451e},
  {32'hc4bf77a2, 32'hc231f178, 32'h42ad9212},
  {32'h44b1ed32, 32'h42c79160, 32'hc2ad353e},
  {32'hc4f589f7, 32'hc33b54fb, 32'h435116c1},
  {32'h4438a002, 32'hc2d76462, 32'h4351f91d},
  {32'hc5001587, 32'h42a88425, 32'h42bacbad},
  {32'h44a42b95, 32'hc2d0d795, 32'hc2c35ae6},
  {32'hc4ed3bda, 32'h420014c8, 32'hc28b1dab},
  {32'h44a03687, 32'h420216f3, 32'h41cdce9e},
  {32'hc4139cbe, 32'h42f678aa, 32'h43ba2357},
  {32'h451462fb, 32'h419f0306, 32'h43c38546},
  {32'hc504a014, 32'hc360cabb, 32'h430a6832},
  {32'h44561f29, 32'hc2d771e5, 32'h4322e31e},
  {32'hc42fb9c0, 32'h428bd55b, 32'hc2adbda6},
  {32'h4343b548, 32'h43634c4c, 32'h424570e6},
  {32'hc509c91c, 32'h42ae9364, 32'hc3446bd9},
  {32'h4496e56e, 32'hc39a0133, 32'h42eac084},
  {32'hc4389046, 32'h41ad9b19, 32'h434ba55b},
  {32'h450d56d6, 32'hc3fe7c41, 32'hc3806299},
  {32'hc4318db2, 32'h4416ac33, 32'hc385080f},
  {32'hc27b5720, 32'hc18381fe, 32'hc16abdc9},
  {32'hc24aeb04, 32'hc2ae6465, 32'hc3eb19ad},
  {32'h4421b32b, 32'h42e7afeb, 32'h435f9bcd},
  {32'hc3b19212, 32'h43601eb2, 32'hc2c81bd3},
  {32'h44d6806c, 32'hbf8ba8dd, 32'hc2df9788},
  {32'hc4a237c8, 32'hc1ad98fd, 32'h436bb57a},
  {32'h441655ea, 32'h41357eb7, 32'h42fa96b8},
  {32'hc2465fc0, 32'hc40f7a2f, 32'h422f090a},
  {32'h4403b0fd, 32'h430f78e6, 32'h432dbe8f},
  {32'hc478585e, 32'h43438299, 32'h42faf0c9},
  {32'h42d245a0, 32'hc37fd5e8, 32'hc36b25b0},
  {32'hc36c6439, 32'hc30a9a65, 32'h432a487a},
  {32'h450341c8, 32'h435ea0ec, 32'h43a78c2a},
  {32'hc408eb07, 32'h40aafc43, 32'h433c02ae},
  {32'h4412d8e6, 32'hc2dd1389, 32'hc309f0bd},
  {32'hc4987ac2, 32'h42e5c6bc, 32'h4318beeb},
  {32'h44eb5127, 32'hc1a1de87, 32'h4303f47b},
  {32'hc4ed5654, 32'h4295837c, 32'h4379cf8d},
  {32'h441d24c0, 32'hc21497ee, 32'h434b345e},
  {32'hc4033cce, 32'h43a60845, 32'h41d19560},
  {32'h43d18703, 32'h42101139, 32'h43dd14b4},
  {32'hc50271ed, 32'hc26d30e0, 32'hc398643c},
  {32'h447d3b36, 32'h429c31cf, 32'h42b972db},
  {32'hc50271c4, 32'h43959dbc, 32'h42ddf5c7},
  {32'h45056573, 32'h43d34ed9, 32'h428dcda1},
  {32'hc497a93c, 32'hc2caf6af, 32'h41a0520c},
  {32'h448faffa, 32'h430ac280, 32'hc319054e},
  {32'hc4c1e7ae, 32'hc1021591, 32'h430d7b75},
  {32'h45198365, 32'h4331116c, 32'h426095ac},
  {32'hc3f927c9, 32'hc37cf2c1, 32'hc19d1b8b},
  {32'h44d7e3ae, 32'h43bad26d, 32'hc2bbea7f},
  {32'hc4bcda4f, 32'hc3e33691, 32'hc3ddeb8e},
  {32'hc2856e50, 32'hc2d12964, 32'hc3b49efa},
  {32'hc4ad374a, 32'h42fabb65, 32'hc2e88d84},
  {32'h448966ba, 32'h432e1a2d, 32'hc4228257},
  {32'hc4988efa, 32'hc2a758d4, 32'hc344ffae},
  {32'h443a3737, 32'hc3862770, 32'h42f017ad},
  {32'hc415ae74, 32'hc224b60b, 32'h43342941},
  {32'h450bf1f0, 32'h42876f31, 32'h4352fc61},
  {32'hc4ae98c6, 32'h433cbb03, 32'hc1fcdfa7},
  {32'h44ac7a66, 32'h429404f5, 32'h42e720e3},
  {32'hc4bbb65c, 32'h428a3404, 32'h43bd98ab},
  {32'h4359bba4, 32'hc2a8793c, 32'hc21b3d6e},
  {32'hc383128a, 32'h41882b3c, 32'h43419907},
  {32'h44e362ef, 32'h424ddd50, 32'hc31ccab8},
  {32'hc31cea34, 32'h433429c9, 32'h434a74bd},
  {32'h444a0185, 32'hc2c49741, 32'h427a4c36},
  {32'hc4ccfe94, 32'hc2cc8cb3, 32'h42da5b9e},
  {32'h44e3c5e1, 32'hc3568dbc, 32'hc380ebd7},
  {32'hc50541af, 32'hc3a1c805, 32'hc26b16d1},
  {32'h441a5252, 32'h43b6c6b3, 32'hc2b2b15c},
  {32'hc283b2f0, 32'h433a2a77, 32'h42ca8044},
  {32'h4483f27d, 32'hc34e10cf, 32'hc39cd639},
  {32'hc4c77de0, 32'hc2b34392, 32'h423db173},
  {32'h450385fc, 32'h4215b007, 32'h436982ae},
  {32'hc4acf2d5, 32'h436939e7, 32'h42ce2ba4},
  {32'h44a34e7e, 32'hc1103d6c, 32'hc318fd6c},
  {32'hc4769198, 32'hc3d45cc9, 32'h42e8ce95},
  {32'h4515b7d5, 32'h42a382a1, 32'hc3442dce},
  {32'h4310afb8, 32'hc37fa23e, 32'h43da4ca0},
  {32'h448e5d33, 32'h437c21ac, 32'hc30d5403},
  {32'hc491549c, 32'h43022324, 32'hc051a2c0},
  {32'h44aefa84, 32'hc3b2171d, 32'hc23295ec},
  {32'hc4e5198e, 32'hc3a791a3, 32'h3fd6b808},
  {32'h42560b08, 32'h431635ea, 32'hc31efa22},
  {32'hc4aef2c4, 32'hc389211d, 32'h43493b37},
  {32'hc18fe480, 32'h434052f5, 32'hc2185a5e},
  {32'hc29bb1e0, 32'h430713eb, 32'hc3191609},
  {32'h449a7bbb, 32'hc37c094b, 32'h4364536e},
  {32'hc4c8cc17, 32'hc39aae51, 32'h434f00eb},
  {32'h449b4a2a, 32'hc39c524e, 32'hc232e7ea},
  {32'hc3e8c418, 32'hc1d92f29, 32'hc2eb87b9},
  {32'h442f4c1e, 32'h436b6190, 32'hc38dd41c},
  {32'hc4f2a3b4, 32'hc2c8e879, 32'h426e2b19},
  {32'h440365d3, 32'h43b0d40d, 32'h438c1e11},
  {32'hc400a7f0, 32'h429151e8, 32'hc0d34766},
  {32'h44dc6980, 32'hc2403612, 32'hc1122f9f},
  {32'hc4b8f71f, 32'hc39f07bf, 32'h4370f1f8},
  {32'h446620f0, 32'hc37ba914, 32'hc286d81e},
  {32'hc48d3af2, 32'hc2d82dcb, 32'hc357589c},
  {32'h44d98b28, 32'h4295c085, 32'hc3a44648},
  {32'hc4aa733e, 32'hc2106b58, 32'hc1a2914c},
  {32'h43ed8120, 32'hc39c563e, 32'h438dac51},
  {32'hc4e17252, 32'h43ac3647, 32'hc3d3610c},
  {32'h45094058, 32'hc39c8620, 32'hc279ddb8},
  {32'hc4e55a77, 32'h43c04374, 32'h42ccd624},
  {32'h4505fc66, 32'hc4049192, 32'hc365d8bf},
  {32'hc4d707d2, 32'hc1ae8cd6, 32'h41ac9860},
  {32'h4268fbd0, 32'hc361ef40, 32'hc38a7ca6},
  {32'hc3aac8d1, 32'hc28fb228, 32'hc3511eaa},
  {32'h44c1f1f8, 32'h4104aff3, 32'hc2e958fe},
  {32'h4183b794, 32'h42c36f05, 32'h42817f1b},
  {32'hc1a42580, 32'hc3a6775c, 32'h423a87c2},
  {32'hc4e817b6, 32'h427fd005, 32'h4363d8dc},
  {32'h44befccc, 32'h43cfe13d, 32'hc2954e0d},
  {32'hc38c11a0, 32'h43e0152a, 32'hc3bb2f49},
  {32'h44628428, 32'h431fb39f, 32'hc317280f},
  {32'hc3b5c3e0, 32'h430a7096, 32'h42c2d7d4},
  {32'hc3a108b6, 32'h436b873a, 32'h430a049a},
  {32'hc4213014, 32'h42bbad66, 32'h42a3d5be},
  {32'h44dd099b, 32'hc3cdbdd0, 32'hc38cfaa2},
  {32'hc514483d, 32'h43b89e02, 32'hc218e674},
  {32'h44a415ae, 32'hc1ed19ee, 32'h4313d0e0},
  {32'hc4031af2, 32'h4222224f, 32'h4386743a},
  {32'h44e695f2, 32'h4302634e, 32'hc2707c38},
  {32'hc414e2e9, 32'h43334ebc, 32'hc2d904f5},
  {32'h442f2718, 32'hc3cf7fb3, 32'h42e79989},
  {32'hc4fe991b, 32'hc2fd2400, 32'h400ba794},
  {32'h44d6386b, 32'h4373d3cd, 32'h424cccb7},
  {32'hc4fc4186, 32'h42c6355d, 32'hc11c1036},
  {32'h44ce7d5a, 32'hc3030214, 32'hc37529a2},
  {32'hc4b08fba, 32'hc2505800, 32'h44146e08},
  {32'h448745b1, 32'hc315158d, 32'hc433d5ca},
  {32'hc50ba428, 32'h433cb670, 32'h43df8af9},
  {32'h444dca75, 32'h42c61884, 32'h413cf4b5},
  {32'hc4132f17, 32'h430e4893, 32'h41df5eb2},
  {32'h44a06df1, 32'h431415cb, 32'hc337b260},
  {32'hc3ba6348, 32'h43a14dda, 32'h4366d169},
  {32'h44910220, 32'h4296fdc8, 32'h4349cb70},
  {32'hc4cc8203, 32'h3ff60b94, 32'h41f1a95b},
  {32'h44a23daf, 32'hc2b25c1f, 32'hc20118cc},
  {32'h428d7e14, 32'h43684b30, 32'h4445db13},
  {32'h44a24b94, 32'hc29896fd, 32'hc27c5cf8},
  {32'hc33bd2b4, 32'hc29d04ea, 32'h40021f06},
  {32'h4511e804, 32'h43b6430d, 32'h43dd937d},
  {32'hc5102251, 32'hc3846ed0, 32'hc29550b4},
  {32'h43f20fd4, 32'hc35c1b03, 32'hc39e498a},
  {32'hc511a3af, 32'h41eb351e, 32'h43f765c9},
  {32'h4478b223, 32'h4316a12a, 32'h41ee5281},
  {32'hc48d295f, 32'h40d6a5c6, 32'h431bde2f},
  {32'h45127251, 32'h4355b6a1, 32'h431498ce},
  {32'hc39c541c, 32'hc36ea692, 32'h4362b9e4},
  {32'h44b3a617, 32'hc331c4dd, 32'h42a87a02},
  {32'hc41048d8, 32'h41c3b649, 32'h42ca284f},
  {32'h443db747, 32'hc3252827, 32'h4210abbe},
  {32'hc4a3a2f4, 32'hc22c2584, 32'hc3ee2d46},
  {32'h42528660, 32'h430b2c04, 32'hc254f282},
  {32'hc496a378, 32'h43192da5, 32'h43434e6a},
  {32'h43ead398, 32'h437fb3a4, 32'hc34345e2},
  {32'hc3924f49, 32'h433d7ef1, 32'hc30d1053},
  {32'h45260b9e, 32'h4358d775, 32'h42f2d8c1},
  {32'h4264ab40, 32'hc2b0674f, 32'h4285617e},
  {32'h44a1c0ed, 32'h43ad3dcb, 32'hc3d2115d},
  {32'hc51d3e90, 32'hc3c669a5, 32'hc193c591},
  {32'h44ca530f, 32'hc1153cc5, 32'h42c81787},
  {32'hc2fb7519, 32'hc3a2e809, 32'hc34bfc71},
  {32'h44cfb7f3, 32'h4320dfe3, 32'hc3702b0f},
  {32'hc50d7591, 32'hc394efd2, 32'hc3d0ef25},
  {32'h44ad0136, 32'hc3ec52da, 32'hc39d99c5},
  {32'hc42614aa, 32'hc388d0bf, 32'h40dafbd8},
  {32'h4500d592, 32'hc2ead6c4, 32'hc248b5ec},
  {32'hc3767664, 32'h432840c4, 32'hc2d64bd7},
  {32'h43cc91f7, 32'h42fded8c, 32'hc23524c3},
  {32'hc50648fc, 32'h426f643c, 32'h42cbd624},
  {32'h4492eb5d, 32'hc325c485, 32'hc2fb657e},
  {32'hc2e2022d, 32'h430277a0, 32'hc283cfd4},
  {32'hc23d9fe0, 32'hc1f9ac10, 32'hc38c2828},
  {32'hc500dda7, 32'h434e5c00, 32'h4385fd5d},
  {32'h44f7fc45, 32'hc2a29d90, 32'hc2ad30e3},
  {32'hc515401a, 32'h43078aa0, 32'h421ec981},
  {32'h451e40f6, 32'h430c6042, 32'hc37f9776},
  {32'hc42d246a, 32'hc23e48c2, 32'hc3a091b7},
  {32'h43f76210, 32'h435c05b3, 32'h44234ec0},
  {32'hc4e9da0c, 32'h43857a08, 32'hc30a09a4},
  {32'h4519f1bc, 32'h42a1eb48, 32'hc3af4afa},
  {32'hc5097891, 32'h428102b1, 32'h42cacacb},
  {32'h442cb22e, 32'hc31f1a72, 32'hc2bf3465},
  {32'hc5156c39, 32'hc3430d4a, 32'h4285e6a5},
  {32'h4486e5bc, 32'h42b69358, 32'h4385a368},
  {32'hc308d630, 32'hc3192a69, 32'h4351d267},
  {32'h4516186e, 32'hc1d0cca6, 32'h42e2019a},
  {32'hc50ae804, 32'h419b8fc6, 32'hc3a9c162},
  {32'h44b4c06b, 32'hc2263680, 32'h4394e080},
  {32'hc51130cc, 32'h436ae92b, 32'h43ab8eca},
  {32'h439239aa, 32'h43fe1b27, 32'hc2e3f38d},
  {32'hc503fd81, 32'hc2d9244e, 32'hc34367a8},
  {32'h441872c8, 32'hc1bbdd6e, 32'h406d5752},
  {32'hc4086a3a, 32'h435194d2, 32'h42867852},
  {32'h44cd5812, 32'hc359cff2, 32'hc36a0680},
  {32'hc4da86c0, 32'hbf9c16ec, 32'hc3cd75eb},
  {32'h444d2875, 32'hc38086bf, 32'h43a94110},
  {32'hc4ed4fb7, 32'h428b36f5, 32'h4264d987},
  {32'h441e5446, 32'hc315ca75, 32'hc31c3e0f},
  {32'hc508cbf9, 32'h42c30d15, 32'h43a6869f},
  {32'h4315bd64, 32'h4415d40c, 32'hc284daba},
  {32'hc4fc7601, 32'h4213a0bc, 32'h43227643},
  {32'h450b4e3b, 32'hc3392d56, 32'hc3954833},
  {32'hc482642c, 32'hc3cf395a, 32'h43e07349},
  {32'h44040f40, 32'h42b70ede, 32'hc30b034f},
  {32'hc4e5bcec, 32'hc2520752, 32'hc3b8315c},
  {32'h44082e18, 32'h4379ce87, 32'hc0244206},
  {32'hc4f03112, 32'hc0958a24, 32'hc16eae8f},
  {32'h42fb76ac, 32'h435464f5, 32'hc3c9742c},
  {32'hc4e2bf4d, 32'h440ca56b, 32'hc2e9cfdc},
  {32'h44edced8, 32'hc2cbdfbf, 32'h41c6736b},
  {32'hc238efb1, 32'h42fa90f9, 32'hc3900b20},
  {32'h451f410f, 32'h4396c555, 32'hc326e2a1},
  {32'hc2fc3458, 32'h42570ccd, 32'hc2e22bb0},
  {32'h45026823, 32'h413689c5, 32'hc17fe1d5},
  {32'hc4fe8ff6, 32'hc2df931b, 32'hc3b38697},
  {32'hc3fc6fd8, 32'h44112efa, 32'h42be5add},
  {32'hc5158c00, 32'hc361f308, 32'h42db3a4c},
  {32'h441cc988, 32'hc2e9d0cb, 32'h431d8b3b},
  {32'hc5078f66, 32'h4211452e, 32'h40a47f42},
  {32'h410ad5a0, 32'h437cab76, 32'h43819b76},
  {32'hc4ad215f, 32'h431dc051, 32'hc207e064},
  {32'h4506aa14, 32'h4286278e, 32'hc08e0592},
  {32'hc5099354, 32'h40670290, 32'h435b194e},
  {32'h44b6adab, 32'h43d76d69, 32'h43321468},
  {32'hc50513fa, 32'hc0b028e2, 32'h4270a8ba},
  {32'h4513428f, 32'hc21e3fd9, 32'hc3caf5ca},
  {32'hc4c70aae, 32'h42fddecf, 32'h42d0d430},
  {32'h44f82e6e, 32'h44003f23, 32'hc1535adb},
  {32'hc4810776, 32'h439ae5a4, 32'hc391abf1},
  {32'h44bf9879, 32'hc3f90f6c, 32'h4328f800},
  {32'hc40fe4e7, 32'h439a9dbb, 32'hc40a235f},
  {32'h42dd5720, 32'h419d2e82, 32'hc34c2a7f},
  {32'hc4d23d70, 32'hc2844a11, 32'h42ee2c80},
  {32'h447d03e7, 32'hc298dac2, 32'h433b024c},
  {32'h436d2c10, 32'h430ef5da, 32'hc2d9146f},
  {32'h44ec17ee, 32'h4354c21d, 32'hc38155d9},
  {32'hc488caee, 32'h40c27e76, 32'h412449a6},
  {32'h42e9dcc0, 32'h439357e2, 32'h4382396e},
  {32'hc3517908, 32'hc406bb93, 32'h432a5217},
  {32'h44f87e7a, 32'hc24d539e, 32'hc0a12faa},
  {32'hc1698e80, 32'h438da546, 32'h419023da},
  {32'hc50daef6, 32'hc2b338bc, 32'h42c161bc},
  {32'h4501adb6, 32'h433ca528, 32'h425b412a},
  {32'hc5158f41, 32'hc2905872, 32'hc2e66f10},
  {32'h43783630, 32'hc273f228, 32'h431ae219},
  {32'hc4b0bc70, 32'hc22b9f93, 32'hc32b600b},
  {32'h44799116, 32'hc39faab2, 32'hc2cc1e0e},
  {32'hc4402948, 32'hc3a27b00, 32'hc21b008e},
  {32'h44d2469c, 32'h418cf90f, 32'hc203a104},
  {32'hc4bf7a77, 32'hc33004c9, 32'h41ae2693},
  {32'h44a3a0b2, 32'h402e3f5c, 32'hc334de41},
  {32'hc4f12648, 32'h4255ec08, 32'hc343faec},
  {32'h45086794, 32'h43577876, 32'h433a8612},
  {32'hc4e0d102, 32'h41db8408, 32'h42b7942b},
  {32'h43f049b4, 32'hc2a23388, 32'hc309694b},
  {32'hc459f48c, 32'h43a9938a, 32'h43ae1e47},
  {32'h441a4526, 32'h433f4dde, 32'h43c0a0e8},
  {32'hc50f64fb, 32'h42e45015, 32'h42951a36},
  {32'h44ea6e50, 32'hc2cecc70, 32'h42b3af03},
  {32'hc4f7be74, 32'h433412ae, 32'h42c28f49},
  {32'h4383a6c0, 32'hc2140a1c, 32'h42e85e88},
  {32'hc5084a3a, 32'h43c9cb50, 32'hc3bd4f59},
  {32'h45088e64, 32'hc19f3c90, 32'h429adee9},
  {32'hc517318b, 32'hc3f228d5, 32'hc2317256},
  {32'h44873d3f, 32'h42569623, 32'h43c0fb95},
  {32'hc4d898ed, 32'h42c57c2c, 32'hc2b833e8},
  {32'h43fe314c, 32'h43233696, 32'h4289cdab},
  {32'hc506eb0a, 32'hc3310d4c, 32'h432810d7},
  {32'h450803a3, 32'h4295d7ad, 32'h42c7d9a6},
  {32'hc52308f4, 32'hc40e47d3, 32'hc3a74b4c},
  {32'h442ab1c2, 32'h432e5c41, 32'h423e5244},
  {32'hc42bf1b8, 32'h4360ad26, 32'h421c4fc2},
  {32'h44cf8af4, 32'hc2a52dd5, 32'hbff833c0},
  {32'h41a94e00, 32'h4363ee67, 32'h43341623},
  {32'h44a05736, 32'hc2acae5e, 32'h43869734},
  {32'hc517279a, 32'hc3148553, 32'h41eb3c1a},
  {32'h428a1080, 32'hc3cc4888, 32'h4358862d},
  {32'hc4d1e164, 32'h43714a63, 32'h43a2cb77},
  {32'h445ab8e3, 32'h4317e7e1, 32'h4390aeb2},
  {32'h42ad09d0, 32'h434279aa, 32'h41e58e9a},
  {32'h44dfaded, 32'h43260d75, 32'h42b40112},
  {32'hc51b0078, 32'h42e820af, 32'hc20247da},
  {32'h4428e43c, 32'hc3989c55, 32'h43deb78d},
  {32'hc483c5d9, 32'hc3a62955, 32'hc29639c0},
  {32'h4460a963, 32'hc38f0d63, 32'h430b9aab},
  {32'hc34f09fc, 32'hc2de5916, 32'hc3157743},
  {32'h44ad56a3, 32'hc28c798d, 32'hc0684ad6},
  {32'hc5021245, 32'h4406e9ef, 32'hc3424610},
  {32'h44ac31c1, 32'h43573b94, 32'h429cd14b},
  {32'hc509dca6, 32'h43173c00, 32'hc33df558},
  {32'h44829ae4, 32'h43e1ddb4, 32'h432cfb70},
  {32'hc45c2246, 32'hc3b4eb0a, 32'hc39aabcd},
  {32'h43228a6c, 32'h43f3a211, 32'hc2b88f97},
  {32'hc4abd375, 32'h42df21c5, 32'hc3b6e4a7},
  {32'h44d101eb, 32'h43b8f583, 32'hc38604f0},
  {32'hc4655dcc, 32'h4385b2f5, 32'hc370a23d},
  {32'hc2122820, 32'hc34a38fb, 32'h4320274c},
  {32'hc494b9e5, 32'hc30f9500, 32'hc3175ca5},
  {32'h448f3404, 32'h43180da2, 32'hc3b775f1},
  {32'hc4f62ff4, 32'hc3d704ce, 32'hc2f3e176},
  {32'hc1ad0120, 32'h428282e0, 32'h42ee6c18},
  {32'hc4c86eab, 32'h43510f1e, 32'h431e5b30},
  {32'h44a642ca, 32'hc2d671b9, 32'h4294e1bb},
  {32'hc49a3254, 32'h42ab5759, 32'hc393e214},
  {32'h4461cd2e, 32'hc354ff95, 32'h4254dc9d},
  {32'hc4af6010, 32'h4310f815, 32'hc2de3f02},
  {32'h447f247f, 32'h43634462, 32'hc3acc302},
  {32'hc502db2e, 32'h4333de54, 32'h42e736f8},
  {32'h436c33ef, 32'h4217778c, 32'hc29e0a93},
  {32'hc447cd0e, 32'h43c88d44, 32'h419ef859},
  {32'h437af538, 32'h40c33d27, 32'hc304587a},
  {32'hc2f79f93, 32'h43203bff, 32'h43282235},
  {32'h44bb9deb, 32'h43079f8c, 32'h43a0f9bf},
  {32'hc4b50cad, 32'h43cd199e, 32'hc3563737},
  {32'h450890f6, 32'hc39ef32c, 32'h4270812c},
  {32'hc4eff5a0, 32'hc0be4bc4, 32'hc3740935},
  {32'h40c8f000, 32'h439d0d82, 32'h42f85e5c},
  {32'hc42a60d9, 32'h432d653b, 32'h42b10789},
  {32'h440b1c9e, 32'h42e7a20b, 32'h3f6ae7e0},
  {32'hc3969a18, 32'h43858122, 32'h430c9a96},
  {32'h44311980, 32'hc3bdb743, 32'h423d7d39},
  {32'hc4e6122e, 32'h42776c69, 32'h42ce1766},
  {32'h44a1eb13, 32'hc3eb6645, 32'h41e3d396},
  {32'hc4eb818b, 32'h42db2a45, 32'hc3bc77da},
  {32'h44c09ebc, 32'h4182c0b2, 32'hc2ea4adb},
  {32'hc2bca920, 32'hc2c8154b, 32'hc30b0fcc},
  {32'h44c5a08e, 32'hc2290e9b, 32'h42eb21e9},
  {32'hc2f1e000, 32'hc3955b7c, 32'h41dbd87e},
  {32'h449fd021, 32'h422b12a0, 32'hc34d46af},
  {32'hc4e27e25, 32'h422b9176, 32'hc3ad29e3},
  {32'h442a6db6, 32'hc32b0093, 32'hc20b6617},
  {32'hc4e2fb74, 32'h43bfb46f, 32'hc326a526},
  {32'h4407086d, 32'h42f150f2, 32'h3fb180ac},
  {32'h43221c5a, 32'hc4118163, 32'hc32fbdff},
  {32'h44620948, 32'hc3c8e4cd, 32'hc34f9d57},
  {32'h413fd400, 32'hc30ceec6, 32'h42ef124f},
  {32'h45145af0, 32'hc236ab05, 32'hc22e6a39},
  {32'hc505ba92, 32'hc36d50cf, 32'hc380a7c4},
  {32'h450f22f9, 32'h425f1fc5, 32'h402daee2},
  {32'hc4d50eae, 32'h4372777b, 32'h430978d6},
  {32'h44cf5edb, 32'hc4271a72, 32'h438ee55f},
  {32'h4327dcc7, 32'h43ea0646, 32'hc2b1cc60},
  {32'h44c933da, 32'h43e44207, 32'h43d14e29},
  {32'hc50fe14d, 32'h438f799a, 32'h42610dec},
  {32'h445143b8, 32'h43b2f79f, 32'h43ef41c8},
  {32'h4380c150, 32'hc2201b35, 32'h428cf73c},
  {32'h43525c35, 32'hc36c7af3, 32'h41e18df0},
  {32'hc4da21bb, 32'h423c91e0, 32'h41924a86},
  {32'h4339ccb6, 32'hc41bffdd, 32'hc3511ba3},
  {32'hc36befb0, 32'h43712fad, 32'hc2de4aae},
  {32'h44ce0433, 32'h44131246, 32'hc3a4ee4c},
  {32'hc4c5b910, 32'h435657c8, 32'h439c8956},
  {32'h44072fa6, 32'h43035ece, 32'h433788d6},
  {32'hc48c5318, 32'h4388c1ce, 32'h4428473a},
  {32'h44ee1058, 32'h428ded76, 32'hc2eee260},
  {32'hc48ef4cc, 32'hc2e624cd, 32'h42ed0913},
  {32'h44d8ac71, 32'h42939569, 32'hc3c24b2e},
  {32'hc464bee4, 32'hc342a4b3, 32'hc3268340},
  {32'h432fa460, 32'h423d4498, 32'h439f4534},
  {32'hc4b8375f, 32'hc30c6e1e, 32'h43d88337},
  {32'h445eda37, 32'hc2991418, 32'hc3a06f5a},
  {32'hc1895540, 32'h4028d104, 32'h437ce4ba},
  {32'h44213618, 32'h4432acb5, 32'h431a47ba},
  {32'hc4e62b41, 32'h43008fea, 32'h42bf465f},
  {32'h42d9b930, 32'hc3900943, 32'h432a771b},
  {32'hc4899874, 32'h414efdb2, 32'h4308898c},
  {32'h45091290, 32'h4353207a, 32'hc333f7d3},
  {32'hc50e72bc, 32'hc0f576a2, 32'h42aad598},
  {32'h442c1d13, 32'hc32e76d3, 32'hc33c80e6},
  {32'hc4979e62, 32'hc23d36ad, 32'hc3a0a2fe},
  {32'h429ea720, 32'h4382826c, 32'h42d659cb},
  {32'hc4aac1da, 32'h4250ccf4, 32'h4365cb55},
  {32'h44b1efd2, 32'hc3221102, 32'h42cfa7d8},
  {32'hc5125e75, 32'h43aa9cab, 32'hc2ada282},
  {32'h44faf0e2, 32'hc334b282, 32'h43188d9a},
  {32'hc4758374, 32'hc32b98eb, 32'h4336bb5e},
  {32'h442cfa82, 32'hc3bad1b8, 32'hc3b9ac1b},
  {32'hc465797b, 32'h42719a5c, 32'hc347d339},
  {32'h4475572e, 32'h439041b1, 32'hc3ebcc0b},
  {32'hc4fb710c, 32'h406336b8, 32'h433397f8},
  {32'h44dd641c, 32'hc2072285, 32'h435fe063},
  {32'hc4afc05a, 32'h43b09ca5, 32'h42098bc6},
  {32'h43bdcc98, 32'hc2cf031b, 32'hc31dad30},
  {32'hc3d241c6, 32'hc365efec, 32'hc31382d0},
  {32'h446a96ce, 32'hbde3d900, 32'h4391977f},
  {32'hc4e00aa2, 32'h437d415b, 32'h4190207f},
  {32'h44d15fdd, 32'hc391f2c1, 32'hc399e3c9},
  {32'hc4940346, 32'h441e066f, 32'h433e4bbb},
  {32'h450ec5b6, 32'h43524066, 32'hc34a8b1a},
  {32'hc50056a4, 32'h439d40f2, 32'h43c0be80},
  {32'h45124050, 32'h4341b7e3, 32'hc186db3d},
  {32'hc496f860, 32'hc395e49b, 32'hc25645e3},
  {32'h4428dff8, 32'h43659126, 32'h43ca3dce},
  {32'hc0285350, 32'hc28ae6e1, 32'hc44c7270},
  {32'h44477676, 32'hc2cf9072, 32'h42a3d978},
  {32'hc4fc7dbc, 32'h424c6af4, 32'hc083815f},
  {32'h440818ca, 32'hc34a3ab8, 32'hc30280a8},
  {32'hc3ac2a28, 32'hc2c9e8f0, 32'h43926100},
  {32'h438b67f1, 32'hc29de198, 32'h435f3388},
  {32'hc4b82a7c, 32'h41983896, 32'h4325b5fb},
  {32'h44357658, 32'hc3895c02, 32'h43ae768c},
  {32'hc3815097, 32'h432b3917, 32'h40d94218},
  {32'h44c40384, 32'hbfeeb83b, 32'hc329da06},
  {32'hc4703e3c, 32'h4282269c, 32'hc3dd3ee0},
  {32'h44349ab7, 32'h43e92cd0, 32'hc2b051fa},
  {32'hc4c3c595, 32'hc224aebe, 32'hc1bd7751},
  {32'h44b778c7, 32'h42164937, 32'h4300ad2e},
  {32'hc4a8e8e7, 32'hc357bb00, 32'hc3e7ced3},
  {32'h44c091ba, 32'hc300ef94, 32'h438a6ff0},
  {32'hc4ae190a, 32'hc3d154ae, 32'hc29f530f},
  {32'h44b8fa08, 32'hc3e9e70e, 32'h43950d76},
  {32'hc3a79a96, 32'hc3791bf7, 32'hc37dea22},
  {32'h44e183b6, 32'hc297d298, 32'hc3592827},
  {32'hc3bbf4e4, 32'h4257dcc8, 32'h43bd3da7},
  {32'h44c8dedf, 32'h430d3b45, 32'h43bf0e42},
  {32'hc4b642bb, 32'h42563686, 32'hc3647684},
  {32'h4394fd20, 32'hc3297e42, 32'hc2c23d8a},
  {32'hc4543954, 32'h42d9ac46, 32'hc317ff38},
  {32'hc370c778, 32'hc3b4266e, 32'h43831ef2},
  {32'hc399dd7c, 32'h436cfc2b, 32'hc3580027},
  {32'h44ae9804, 32'hc2d76b11, 32'hc2ecf872},
  {32'hc50f8f89, 32'hc21287a5, 32'h432ee5b6},
  {32'h44ecddae, 32'h444a4bb8, 32'hc20ed852},
  {32'hc48f3fa3, 32'hc13e87f7, 32'h422a39b0},
  {32'h4436f05a, 32'h431fdb73, 32'hc35d2cd4},
  {32'hc4f18974, 32'hc304a5a9, 32'h435a1e29},
  {32'h44646f99, 32'h426ff738, 32'h438b3c45},
  {32'hc467c38a, 32'h43c54a78, 32'h44222e0e},
  {32'h44ddc52c, 32'hc2eb3370, 32'h4086e99c},
  {32'hc2eaa20a, 32'hc34cb519, 32'h42f6089c},
  {32'h44e78ade, 32'hc366b57f, 32'h41a8dadd},
  {32'hc4068424, 32'hc304290c, 32'h425a985d},
  {32'h44b338aa, 32'h438b90d2, 32'h43f555a0},
  {32'hc3cd57b8, 32'hc28adbee, 32'hc330bd93},
  {32'h44360c20, 32'hc29e5a82, 32'hc26920fc},
  {32'hc4c83955, 32'hc2d3573c, 32'hc3ab1b19},
  {32'h4362a9a9, 32'hc3dc9051, 32'hc2b65d72},
  {32'hc510776d, 32'h43538932, 32'hc2d20205},
  {32'h4417e346, 32'hc35739aa, 32'h439e678c},
  {32'hc481edfb, 32'h430a6009, 32'h434c7d78},
  {32'hc2b39c60, 32'h41d32a9f, 32'h43af3607},
  {32'hc46959c4, 32'hc3c39700, 32'hc30a5d62},
  {32'h4488c94c, 32'h4396d8a1, 32'h428642d8},
  {32'hc4ba4920, 32'hc3ad4427, 32'hc363984d},
  {32'hc3223b78, 32'h432be887, 32'hc3a77899},
  {32'hc4e574b8, 32'hc2be2d55, 32'h438de2a1},
  {32'hc32a3440, 32'hc3b94b60, 32'hc1e7f750},
  {32'hc43f4a62, 32'hc3422364, 32'h43093abb},
  {32'h43c65328, 32'hc2c721b8, 32'hc1b72350},
  {32'hc4e57744, 32'hc1c65070, 32'hc4111f70},
  {32'h44fdf8fe, 32'hc30924d9, 32'hc32780f6},
  {32'hc47b6f66, 32'h41f6d585, 32'h43892a74},
  {32'h4327f59d, 32'hc3737105, 32'hc208a72e},
  {32'hc4c6b651, 32'hc3543731, 32'hc1d091fd},
  {32'h441c9a00, 32'hc40e8a0f, 32'hc2889c70},
  {32'hc5070b07, 32'h43a15fbd, 32'h4291e064},
  {32'h436ab068, 32'hc222603e, 32'h434a08a1},
  {32'hc3e33ffc, 32'hc332fe3f, 32'h3fb8ab58},
  {32'h4439d9ba, 32'h42a6435b, 32'h43e96b5c},
  {32'hc4293c70, 32'hc32833cf, 32'h440fd8a7},
  {32'h4514f39a, 32'hc1ffe382, 32'h438d9dfd},
  {32'hc43d2c1c, 32'h4393ed28, 32'h42dd40e6},
  {32'h440ad9b0, 32'h43125e26, 32'h4300aecd},
  {32'hc399a920, 32'hc0086170, 32'hc1c0be84},
  {32'h4384d430, 32'hc17b0130, 32'h4297a3ec},
  {32'hc48baf3b, 32'hc1cfaa58, 32'h42f18f04},
  {32'h448da538, 32'h439fe263, 32'hc2039cbf},
  {32'hc4f4365e, 32'h40cd20d6, 32'hc2b892b2},
  {32'h44f8edf0, 32'h430f7951, 32'h41071c22},
  {32'hc4f9f481, 32'h42752092, 32'hc222bb1c},
  {32'h42cff496, 32'hc31f9fee, 32'h43856758},
  {32'hc405be30, 32'hc370548f, 32'h4227bc65},
  {32'h44da91e8, 32'h433696dd, 32'h42382266},
  {32'hc49c5b72, 32'h438ea322, 32'hc29b08e5},
  {32'h43e4e718, 32'hc223e2ad, 32'hc2d95a2b},
  {32'hc4bd7504, 32'hc3456b7c, 32'hc2048b6e},
  {32'h4454ba24, 32'hc356951f, 32'h439b8c7c},
  {32'hc4b069ea, 32'hc03ab124, 32'hc2b568f6},
  {32'h43b24014, 32'h4174a3a4, 32'h421f6291},
  {32'hc50ce4ec, 32'hc329d9b2, 32'hc39bb2cd},
  {32'h4292a7e0, 32'h42a01fff, 32'h423d1b40},
  {32'hc5072cd0, 32'h4295bcd0, 32'h424619b1},
  {32'h44930d3b, 32'hc3e1566e, 32'hc2d97cd8},
  {32'hc4ef722e, 32'h4363680a, 32'hc33bb654},
  {32'h44ec8e7b, 32'h41c15b70, 32'hc3e372c3},
  {32'hc4b553ab, 32'hc2a65b45, 32'h41cba045},
  {32'h450c148d, 32'hc31bf56f, 32'hc19d793d},
  {32'hc5042bbd, 32'hc2fd6603, 32'h42606dfe},
  {32'h442e535e, 32'h436c1f4f, 32'h429d3b0d},
  {32'hc4255ec6, 32'h43b1ee75, 32'hc3777051},
  {32'h4387f443, 32'h424aec8f, 32'h432f22cf},
  {32'hc50346b6, 32'h43c8e6b6, 32'hc3c7b3fa},
  {32'h4445132e, 32'hc37a2bfd, 32'h42014d96},
  {32'hc500d863, 32'hc2296be0, 32'h42248f6f},
  {32'h44f27ba0, 32'h430bd495, 32'hc196a7ba},
  {32'hc504a2e8, 32'h42e62223, 32'hc358cb91},
  {32'h44d3c5fc, 32'hc3473b34, 32'hc2a5d6eb},
  {32'hc4f43599, 32'h42b7ba82, 32'hc393f349},
  {32'h44b9b26c, 32'h3ee268f6, 32'hc3974315},
  {32'hc3140460, 32'h4221692e, 32'hc20f6428},
  {32'h44c2ef80, 32'h430f7368, 32'h43dffa54},
  {32'hc3bb4bae, 32'h42be3f0d, 32'hc33bda96},
  {32'h44e7e743, 32'h426967e1, 32'h4304d4cd},
  {32'hc50c24c4, 32'hc3b0283c, 32'h428b8258},
  {32'h44d321a6, 32'h4327d35e, 32'hc3ade5e4},
  {32'h43305014, 32'hc3b453d2, 32'h41785dec},
  {32'h44c773ee, 32'hc361176a, 32'hc2ad1af2},
  {32'hc4da9ed2, 32'hc360cd36, 32'hc3aeee77},
  {32'h44b4e5f8, 32'hc3f69b85, 32'h4377ed4c},
  {32'hc43d01cb, 32'hbfc5738a, 32'hc2291b56},
  {32'h4433c9d4, 32'h4045c650, 32'h42e781d5},
  {32'hc2d58ea0, 32'h43a3b7dd, 32'h42e3cf2e},
  {32'h44f400d0, 32'hc30e6eb6, 32'h42d2846e},
  {32'hc46d5d81, 32'hc2b28e0a, 32'hc405f356},
  {32'hc2c79300, 32'h433ef9cd, 32'h41e4e3ae},
  {32'hc51078fc, 32'h43381828, 32'hc1e641f4},
  {32'h43863b86, 32'hc2fc268d, 32'h430d3beb},
  {32'hc4d63e1e, 32'hc3ba7427, 32'h4376323a},
  {32'h44fc19dc, 32'h428cbb3a, 32'hc1f10653},
  {32'hc4b184bb, 32'hc33b73dd, 32'h42e2668e},
  {32'h4485c5f4, 32'hc3cc9821, 32'h42ec29bd},
  {32'hc400ebf8, 32'hc28ed16f, 32'h439daf2d},
  {32'h44918f3c, 32'hc30f493c, 32'h430c1b7a},
  {32'hc1be294a, 32'h42fc104b, 32'h4397d978},
  {32'h44f078be, 32'hc2e1e140, 32'h4202f8b8},
  {32'hc330ac28, 32'h4386f352, 32'hc1ef2646},
  {32'h447f032c, 32'hc42ea1b4, 32'h430322ef},
  {32'hc50e3f24, 32'h4319eb64, 32'h4324d8c3},
  {32'h4428da52, 32'hc3822640, 32'hc2eab150},
  {32'hc4d65952, 32'h41ed2286, 32'hc223a950},
  {32'h449ad64c, 32'h4310323e, 32'hc295f539},
  {32'hc4310160, 32'hc2ca71e2, 32'h4306863e},
  {32'hc210d4d8, 32'h435a7904, 32'hc2d9c46d},
  {32'hc448c229, 32'h437acc11, 32'h42bfe364},
  {32'h4390c577, 32'h439175ad, 32'hc2c9edd4},
  {32'hc41a61f0, 32'hc304fdc9, 32'hc383f2f2},
  {32'h44d88ea7, 32'hc2134f05, 32'hc41bc0bb},
  {32'hc4e4a82a, 32'hc1bfcaa0, 32'hc352719d},
  {32'h43d12590, 32'hc38c8b4b, 32'h43cadb0a},
  {32'hc41ea2f6, 32'h43bcf3fa, 32'h43538320},
  {32'h441beb7c, 32'hc19cc27c, 32'hc2122a66},
  {32'hc4861e44, 32'h4285dc9b, 32'h43307ead},
  {32'h44cfa96b, 32'h430011bf, 32'h430d05d5},
  {32'hc51ad672, 32'h42366aa9, 32'hc32fc7fa},
  {32'h4504c20d, 32'h41dcef54, 32'hc2f96923},
  {32'hc439af28, 32'hc20fcf35, 32'hc4118ba1},
  {32'h450d9dcf, 32'hc2e5050b, 32'hc2f42c9b},
  {32'hc42d34e6, 32'hc25e0882, 32'hc3a8f921},
  {32'h44af56d2, 32'hc39254c2, 32'h4363be91},
  {32'hc4f44765, 32'hc3368a3b, 32'h40899018},
  {32'h452732ae, 32'h433e5da4, 32'h43fdf8be},
  {32'hc42da4c9, 32'hc28bd48a, 32'hc1c8a4dc},
  {32'hc4ce90c3, 32'hc35c9e2a, 32'hc3c8426b},
  {32'h44b3afb7, 32'hc2fa084c, 32'h437f23b6},
  {32'hc4f2261f, 32'h432c8291, 32'hc3ec8d9a},
  {32'h44a388cc, 32'hc240fda4, 32'hc35a9085},
  {32'hc43dcf5a, 32'hc30a1238, 32'hc2a663b6},
  {32'h44b028e3, 32'h42087706, 32'h42f75da5},
  {32'hc4d42ae5, 32'h43d9b163, 32'hc0825d08},
  {32'h44ef5535, 32'h424b5981, 32'h4292cf0d},
  {32'hc30be81c, 32'hc38771b4, 32'hbf175c07},
  {32'h44874146, 32'hc42d3c99, 32'h43c39e81},
  {32'hc49243c4, 32'hc3a134b0, 32'hc2dc34d2},
  {32'h4491cfb9, 32'hc34d6cf0, 32'hc27f452b},
  {32'hc38a3c47, 32'hc2b6b848, 32'h42ab8393},
  {32'h439cd61c, 32'hc2ee0174, 32'h43827488},
  {32'hc45445ab, 32'h42e3b660, 32'hc2b889c4},
  {32'h444606e8, 32'h42cea062, 32'hc3a5b0fb},
  {32'hc39d89d0, 32'h4288bb4d, 32'h422a04bb},
  {32'h449fda56, 32'h4402ec90, 32'hc16af8e8},
  {32'hc4653a26, 32'hc36ff34a, 32'hc3890619},
  {32'h44ff116b, 32'hc3e262f4, 32'hc39bb2d4},
  {32'hc475a9ca, 32'h422a22f3, 32'h3f11d9ee},
  {32'h440ca519, 32'h43c82e62, 32'hc3467e04},
  {32'hc4ac5807, 32'hc1363e84, 32'hc347fc7e},
  {32'h450e54a2, 32'hc30ad624, 32'hc1b06071},
  {32'hc49539e0, 32'hc3f03f42, 32'h4301fbc5},
  {32'h442520ae, 32'hc32b6146, 32'h427c8120},
  {32'hc4ed7904, 32'h4320f0e5, 32'h4210da4c},
  {32'h44c9988b, 32'hc336eba4, 32'h43668a6e},
  {32'hc463e98a, 32'h4248be1c, 32'h43ce7902},
  {32'h4430718e, 32'h42cc1908, 32'h430c3a96},
  {32'hc5102ed7, 32'h438d919c, 32'h42ac00b1},
  {32'h43f9fa32, 32'h43c25b74, 32'hc2d7529d},
  {32'hc4bb0a5a, 32'hc2b91ca2, 32'h42fe5872},
  {32'h4502df1e, 32'h435de708, 32'hc36b2067},
  {32'hc3656a8a, 32'hc3dd7d15, 32'h3fc93c32},
  {32'h44adf2e8, 32'hc37f4d89, 32'hc402a159},
  {32'hc4828d09, 32'hc28f4b22, 32'hc36e59d6},
  {32'h44c028c2, 32'hc1fff831, 32'h428e87ec},
  {32'hc41bc0b8, 32'h429e8a88, 32'hc3155f31},
  {32'h4503d653, 32'hc34d542e, 32'h42515721},
  {32'hc3008cbf, 32'hc2b690c6, 32'hc329b92e},
  {32'h4431f0ac, 32'hc41944a3, 32'h4312e239},
  {32'hc4894880, 32'h421402ae, 32'hc2972a88},
  {32'h44d26c08, 32'hc3d9257a, 32'h43d197e5},
  {32'hc4a3b7d9, 32'hc227fad4, 32'hc2c68bdb},
  {32'h44c80680, 32'h417c3855, 32'hc25ee0cc},
  {32'hc41bc3b8, 32'h422ec9de, 32'h439808e8},
  {32'h44a7e451, 32'h435ba14b, 32'hc223ea7f},
  {32'hc50f5aee, 32'h4295fef4, 32'h43134038},
  {32'h44d96d38, 32'h43435f46, 32'h41ce7707},
  {32'hc4bc2c64, 32'h427fac85, 32'hc398ca60},
  {32'h44aadf6c, 32'h426d9b87, 32'h43e22782},
  {32'hc417a47c, 32'hc3baa35a, 32'hc34d197b},
  {32'h42fa8160, 32'h433cc4da, 32'hc2ab3a1d},
  {32'hc421d3fd, 32'h43154224, 32'h43b162c2},
  {32'h44daf498, 32'h42fc12af, 32'h431261d2},
  {32'hc40e1709, 32'hc39175f0, 32'hc3502be2},
  {32'h45181587, 32'h4392669e, 32'hc299ea5c},
  {32'hc4d9fd8e, 32'h434dcd67, 32'h42e7663e},
  {32'h4418e234, 32'hc3f1d1d3, 32'hc2101a08},
  {32'hc4bf4114, 32'hc3d6d09c, 32'hc3253834},
  {32'h447b086a, 32'h425c77b0, 32'h43b8a3d2},
  {32'hc4fca562, 32'h4339a3b6, 32'h42393be5},
  {32'h44f9c9d5, 32'h42817d17, 32'hc2d6fbea},
  {32'hc512cb1f, 32'h42726fc8, 32'h43aaaa19},
  {32'h44ff2f97, 32'h435daebc, 32'h437814ee},
  {32'h42de948b, 32'hc33c84ee, 32'h41b00b92},
  {32'h44f8e606, 32'h435d2020, 32'h428890ef},
  {32'hc4f9a253, 32'hc3eee642, 32'hc29f3a73},
  {32'h44444816, 32'h4249b43d, 32'hc2b93412},
  {32'hc508f8dc, 32'hc2b65f7b, 32'hc1b4db59},
  {32'h44d5466f, 32'hc3719db5, 32'hc2c28ccb},
  {32'hc446ca5f, 32'h437e087a, 32'h435269c6},
  {32'h44ff7876, 32'hc3b98ef7, 32'hc30ca99c},
  {32'hc50cb900, 32'h4235c2db, 32'hc36642c0},
  {32'h43ac22bd, 32'hc3200058, 32'hc379d55a},
  {32'hc4d3eb18, 32'h43683342, 32'h4301b445},
  {32'h44da5ed8, 32'h4310e102, 32'h41cf7a8a},
  {32'hc48b7842, 32'h4158eeb2, 32'hc3527d2a},
  {32'h44f6ded1, 32'hc323b622, 32'hc3bd8171},
  {32'hc46438a0, 32'h4305b7d9, 32'h43006562},
  {32'h433e34b0, 32'h4198b370, 32'h42231d5f},
  {32'hc40d1f1e, 32'h431513af, 32'hc33c0e6b},
  {32'h442c02a8, 32'hc2ba8828, 32'hc339788c},
  {32'hc4878932, 32'h43a53ded, 32'hc25e0cef},
  {32'h440b8c32, 32'hc3c22294, 32'hc308f57b},
  {32'hc5126fbc, 32'hc06c0bfa, 32'hc357d754},
  {32'h44a9cbe4, 32'h4388e709, 32'hc3887e51},
  {32'hc5053032, 32'hc24e6077, 32'hc293a653},
  {32'h44e6cb81, 32'h41bb4da8, 32'hc2addca7},
  {32'hc4fda360, 32'hc3273840, 32'hc2934249},
  {32'h451119c8, 32'h43a32f5e, 32'hc36ac88a},
  {32'hc44168c0, 32'hc2d372b2, 32'h438c5144},
  {32'h443b6441, 32'h430d3989, 32'hc3a49ecd},
  {32'hc3de3c5c, 32'hc393dc51, 32'hc27cd781},
  {32'h44218d2e, 32'h42b0cc2d, 32'hc3004fe1},
  {32'hc4a08e27, 32'h4342f17f, 32'hc281a509},
  {32'h444372bc, 32'h42911714, 32'hc276b374},
  {32'hc49b4ef1, 32'hc24799cf, 32'h43700c32},
  {32'h446bfd80, 32'hc3a10c05, 32'hc3b5fbe0},
  {32'h42a37136, 32'hc2583ae3, 32'hc018ed3d},
  {32'h44ab37af, 32'hc2b6d231, 32'h42e66292},
  {32'hc3386c70, 32'h438a5a10, 32'h4421d548},
  {32'h44f1dcd9, 32'hc28375a8, 32'hc2922560},
  {32'hc4bff8aa, 32'h43e0c138, 32'hc31e6404},
  {32'h447e8d3e, 32'hc2fa8fad, 32'h41242da1},
  {32'hc3ef166c, 32'h42a702bf, 32'h434787a4},
  {32'h43a21292, 32'hc308b21a, 32'hc2590598},
  {32'hc503a634, 32'hc3f8a50a, 32'hc2222caa},
  {32'h451495b8, 32'hc2dbb4fb, 32'h431d4988},
  {32'hc4ce8cf8, 32'h43356253, 32'h4340396b},
  {32'h450deed6, 32'h411dc571, 32'hc33dd49b},
  {32'hc44fb96e, 32'hc327352b, 32'h439b5094},
  {32'h4515524e, 32'h3f843ab0, 32'hc2317d7a},
  {32'hc4555fb0, 32'h43161323, 32'hc3045a69},
  {32'h4501b71a, 32'h4235b94e, 32'hc296b2dd},
  {32'hc4bf92b8, 32'h419c8c8f, 32'hc24560ca},
  {32'h4420311c, 32'h434300e8, 32'hbfc74022},
  {32'hc35e8b64, 32'h432b86a9, 32'hc206066e},
  {32'hc30fce70, 32'hc36733e9, 32'hc30798a4},
  {32'h44afcc2a, 32'h43baac10, 32'hc364ce7b},
  {32'hc4e9ba34, 32'hc39a2b96, 32'hc004cf1d},
  {32'h4441b000, 32'h439e9815, 32'hc409fece},
  {32'hc420cd42, 32'h42f8a503, 32'h42a51078},
  {32'h44a1f7ea, 32'hc36a40f0, 32'h43093a38},
  {32'h42080a00, 32'h41d7beff, 32'hc2ff6e00},
  {32'h44ac13f4, 32'hc3a17867, 32'h43bddff9},
  {32'hc502fe41, 32'hc3a398c8, 32'hc195ba1e},
  {32'h44854efe, 32'h42283422, 32'hc3844176},
  {32'hc3b39288, 32'hc351ef4a, 32'h43914043},
  {32'h44b6157c, 32'hc26ccb96, 32'hc39bc7b7},
  {32'hc4997d15, 32'h43a35596, 32'h42356b06},
  {32'h44ed1b44, 32'h428b0c61, 32'hc2d6d652},
  {32'hc397c6f4, 32'h430d385b, 32'hc1f23125},
  {32'h43cb291a, 32'h436a25be, 32'hc3e1ed3f},
  {32'hc3ff6de3, 32'hc33c588e, 32'hc3e6648d},
  {32'h43d14f32, 32'hc2d1b875, 32'hc1ed151f},
  {32'hc4fdaa7a, 32'h43179e98, 32'hc2c88820},
  {32'h450bf3cd, 32'hc39d1da9, 32'hc362ebfd},
  {32'h41845ee0, 32'hc1bf630b, 32'h43297770},
  {32'h45022755, 32'hc2ce9a79, 32'h439dec8a},
  {32'hc3af2d78, 32'hc344413b, 32'hc2d3c5ea},
  {32'h43e33380, 32'hc2d2ffa3, 32'hc342f852},
  {32'hc500e051, 32'hc3983625, 32'h42936170},
  {32'h44bbc625, 32'hc38ea01e, 32'h4144557a},
  {32'hc4a72848, 32'hc33b4d67, 32'hc25cc2f5},
  {32'h44e575b8, 32'h42054d1d, 32'hc34c7a78},
  {32'hc4526a27, 32'hc2ea14ef, 32'hc394035c},
  {32'h4403cd8c, 32'hc298b1a4, 32'hc3290284},
  {32'hc43fb84f, 32'h420d177d, 32'h437cabb7},
  {32'h441a4aa4, 32'h42f2c34f, 32'hc1096095},
  {32'hc4a23727, 32'hc369bff4, 32'hc22dffaa},
  {32'h44593bd1, 32'h434f0cc7, 32'hc36aab52},
  {32'hc4a8ae11, 32'hc309feb7, 32'h4311582d},
  {32'h449e6196, 32'h432621bb, 32'h429c0c36},
  {32'hc4fa7e2f, 32'hc34cd170, 32'h430e71f7},
  {32'h45102d20, 32'h438888b2, 32'hc1a53480},
  {32'hc404a04d, 32'h4396346b, 32'h43d0b5ca},
  {32'h44955b54, 32'h430cc122, 32'h42bef22e},
  {32'hc41c7370, 32'h41f4c16d, 32'hc4333a1a},
  {32'h42bae2c6, 32'hc405f454, 32'hc2cedeb6},
  {32'hc4ed887d, 32'h43cbfc0d, 32'hc3bdc825},
  {32'h44b0c615, 32'hc3ca5d60, 32'h435a6598},
  {32'hc4fe0f07, 32'h42ec2c37, 32'hc2103098},
  {32'h4505c160, 32'h42700971, 32'hc2992dcd},
  {32'hc45437a0, 32'h4311fb0a, 32'h43ff9458},
  {32'h44925dad, 32'hc1227364, 32'h43428698},
  {32'hc4689363, 32'hc29b8c37, 32'hc340cfce},
  {32'h44dddf3a, 32'h43517ae7, 32'h41600e6c},
  {32'hc451175a, 32'hc1cd2c9d, 32'hc2c245c3},
  {32'h4508d45a, 32'h41c92db6, 32'hc357f762},
  {32'hc4ac9f55, 32'h43c9f530, 32'hc31518bd},
  {32'h441d1898, 32'h42da491d, 32'h42ac5469},
  {32'hc4946634, 32'hc22dcc36, 32'hc2d0b8ee},
  {32'h45181fa1, 32'h4182ae61, 32'hc3d434a2},
  {32'hc4bc3fc8, 32'h421ca7b7, 32'hc3aca102},
  {32'h4513f673, 32'h438d597c, 32'hc38ecb21},
  {32'hc3d3d570, 32'h434fb32d, 32'hc315d4fc},
  {32'h449c468c, 32'h43b7ed55, 32'hc23e3556},
  {32'hc4c968de, 32'h4207a0ef, 32'h4384fc96},
  {32'h4510ab25, 32'h422ad13e, 32'h42a4c122},
  {32'hc49cf230, 32'hc28ad370, 32'hc3869a2f},
  {32'h450de169, 32'hc37213c8, 32'hc2a5ad47},
  {32'hc3fce481, 32'hc3536a1d, 32'hc1b7e9de},
  {32'h44b9ea1c, 32'h43e31204, 32'hc38c3f8f},
  {32'hc44d92c2, 32'h4377f792, 32'h441095e4},
  {32'h44d7d981, 32'hc317ce03, 32'hc3d628a0},
  {32'hc4a9f64b, 32'h42b85a5d, 32'hc287b2be},
  {32'h44cd95fd, 32'h437cf894, 32'h42431b9c},
  {32'hc4424db0, 32'hc3439ce4, 32'hc3554027},
  {32'h439d0bc7, 32'h439c65fa, 32'h43b8315c},
  {32'hc4d93d29, 32'h42fb9874, 32'h41c2c7c3},
  {32'h4500c39d, 32'h43d3d1ca, 32'hc388b73c},
  {32'hc514b380, 32'h42a98b7b, 32'hc31bdc45},
  {32'h44b98eca, 32'h43d21a86, 32'h422b2253},
  {32'hc3a8c04c, 32'hc217e820, 32'h42420e46},
  {32'h4489df48, 32'h42a090e2, 32'hc4030e2c},
  {32'hc4751f88, 32'h42ad455c, 32'hc3aa08dc},
  {32'h44c385a6, 32'h41f1a15d, 32'hc333c605},
  {32'hc4a7971f, 32'h43130f69, 32'h42978e99},
  {32'h4452cdd3, 32'h42286a8b, 32'h433545c0},
  {32'hc4bfc918, 32'h42a75fcd, 32'hc2af66aa},
  {32'h443a5fe3, 32'h439858cd, 32'hc205fa68},
  {32'hc509ca27, 32'h43c3bd06, 32'h429e0875},
  {32'h4344b780, 32'hc3a08fb5, 32'hc32a188b},
  {32'hc4090bfe, 32'h418d115b, 32'h429450ce},
  {32'h44005cd5, 32'hc3812950, 32'h40915ba5},
  {32'h43cd8a94, 32'h42b5c335, 32'hc331516a},
  {32'h44652cb8, 32'hc0afc73e, 32'hc322c871},
  {32'hc4c21dcb, 32'hc360315f, 32'h41d0e502},
  {32'h451617c4, 32'h43885b81, 32'h422899d2},
  {32'hc49195d2, 32'h42c1ac20, 32'h43f4b4fa},
  {32'h449f2741, 32'h412920bb, 32'hc382da25},
  {32'hc4f4f2db, 32'h435175f0, 32'hc338d81b},
  {32'h44fb690c, 32'h437d89dd, 32'hc3542f1e},
  {32'hc501e15f, 32'hc325ee47, 32'h42fb0237},
  {32'h44f9a838, 32'h4257ce65, 32'h436d7f04},
  {32'hc502d986, 32'hc330c9ea, 32'hc292995f},
  {32'h44545447, 32'h41fc51a1, 32'h41be3ec4},
  {32'hc4b97770, 32'h42da4b56, 32'h424980db},
  {32'h450eb596, 32'hc23e74f5, 32'hc12bf4be},
  {32'hc50181ae, 32'h4277efc6, 32'hc377bcb2},
  {32'h43e75f19, 32'h435c9193, 32'h4333e427},
  {32'hc4cc7cd6, 32'h42f623b6, 32'h43d7968e},
  {32'h43bcfc84, 32'hc32aaaf6, 32'h43022fa4},
  {32'hc49bc120, 32'hc2a86302, 32'h42a54fe2},
  {32'h44577843, 32'hc3a0be0e, 32'h42cbee4c},
  {32'hc4712b5b, 32'hc3f5fa03, 32'hc280110f},
  {32'h445e1975, 32'hc2fa34d2, 32'h43def1a2},
  {32'hc51e9cd2, 32'hc35e0ffe, 32'hc3319cba},
  {32'h44649708, 32'hc37b4986, 32'h42bcf75d},
  {32'hc42aa244, 32'h43a0b8ca, 32'h434f7d95},
  {32'h4501edeb, 32'h431c6fc1, 32'h43b5d3b8},
  {32'hc4ef9e10, 32'hc38794f6, 32'h43c02e20},
  {32'h4352e620, 32'h43645db8, 32'h4344f256},
  {32'hc407d3a7, 32'h43c46d95, 32'hc20c9883},
  {32'h44dc1f60, 32'hc32a8974, 32'h438599aa},
  {32'hc45bc988, 32'h42825637, 32'hc35b5513},
  {32'h43351090, 32'hc2885489, 32'hc3614bcb},
  {32'hc502316a, 32'hc2dc3e5a, 32'h424d59e5},
  {32'h44e50509, 32'h427f04bd, 32'h4385c3c4},
  {32'hc49fb506, 32'h4235b4e0, 32'h43979c10},
  {32'h44cfd472, 32'h43a9fedc, 32'h43a008d7},
  {32'hc46145c1, 32'hc3d607e2, 32'h43654d67},
  {32'h44448211, 32'h439a3039, 32'hc1069dbe},
  {32'hc4ee5ec6, 32'hc1cee169, 32'h435eda27},
  {32'h44efa5b1, 32'hc26d5351, 32'hc3902c15},
  {32'hc4ce0d53, 32'hc3bebe28, 32'h43acb88d},
  {32'h44790bd2, 32'h42eed2fc, 32'h4318786a},
  {32'hc331fa60, 32'h43465033, 32'h43476bee},
  {32'h4434e42a, 32'hc381f5cd, 32'h425d179f},
  {32'hc5287cf9, 32'h422bac6e, 32'hc31122bc},
  {32'h44b7acad, 32'hc13c0335, 32'h4321f83c},
  {32'hc49a092e, 32'hc351d8ac, 32'h439e8ce5},
  {32'h44205af3, 32'h4380304d, 32'hc2bd5e02},
  {32'hc4c5930b, 32'hc364620e, 32'hc336a42d},
  {32'h44d67756, 32'hc302a795, 32'hc36394b7},
  {32'hc3d0613c, 32'h4329c2c9, 32'h42b285ea},
  {32'h448cc772, 32'hc2831a2a, 32'h439911e2},
  {32'hc502e61c, 32'hc309f08d, 32'h41a03900},
  {32'hc1132600, 32'h43925618, 32'h41806cd0},
  {32'hc32658ba, 32'h42f09ab7, 32'h41a9c7c6},
  {32'h44d12baa, 32'h4347c874, 32'h42ea6af9},
  {32'h41de2400, 32'hc39e4ae9, 32'h43d7c5f8},
  {32'h44fd246f, 32'h42c71bd7, 32'h42dc984b},
  {32'hc5089128, 32'h41cd66ce, 32'hc3383998},
  {32'h43e789b0, 32'hc305135f, 32'h42331dbe},
  {32'hc2ebea80, 32'h4340125a, 32'hc3ec5389},
  {32'h44cbdb98, 32'hc2c7a83b, 32'hc09365fa},
  {32'hc497b012, 32'hc3a51042, 32'h4262b02e},
  {32'h44fc0f76, 32'h4266d0c6, 32'h42228110},
  {32'hc5005bd6, 32'hc3c8f049, 32'hc2a3bacb},
  {32'h4473a19f, 32'h43a0243a, 32'hc33665de},
  {32'hc41e0618, 32'h43961f1c, 32'hc26699ab},
  {32'h44da7e55, 32'h4264c971, 32'hc244deb3},
  {32'hc49e7da5, 32'h42b0f390, 32'hc316322b},
  {32'h44f4be02, 32'hc1c5c1d6, 32'hc2cca956},
  {32'hc480f0ab, 32'hc2d1d29e, 32'h42ce2440},
  {32'h4507b5dc, 32'hc3276ea2, 32'hc33c4853},
  {32'hc4812589, 32'h42879607, 32'h40c3ec44},
  {32'h432fc884, 32'hc3271dff, 32'h430b54b9},
  {32'hc4b120fe, 32'hc2672679, 32'hc3aa2ae8},
  {32'h43edafa8, 32'h43a77bda, 32'hc326ec3e},
  {32'hc502b542, 32'hc342d59b, 32'hc1659d0a},
  {32'h44bae241, 32'hc30529ad, 32'hc34a517f},
  {32'h423b8140, 32'h43a58b2f, 32'hc3c37ed2},
  {32'h4481ca25, 32'hc2cf101e, 32'h423db9aa},
  {32'hc31717a0, 32'hc1ad0e44, 32'h42ce57c7},
  {32'h43c82098, 32'hc181881e, 32'h4222a2c6},
  {32'hc3e97a98, 32'h42a27af8, 32'h42262a29},
  {32'h441e94ec, 32'h42cf7707, 32'h43512e90},
  {32'hc39c4b51, 32'hc28f0503, 32'hc1480d58},
  {32'h43b6e610, 32'h42ef76a7, 32'hc296852e},
  {32'hc498243d, 32'h43405107, 32'hc1fbde37},
  {32'h445929eb, 32'hc3916fc8, 32'h4302520b},
  {32'hc3d39253, 32'h42efd932, 32'hc29d6096},
  {32'h44ee99c2, 32'h432cb5e6, 32'hc2b06e91},
  {32'hc4b59dab, 32'hc33e12bc, 32'hc299f23a},
  {32'h450280c9, 32'h428d2320, 32'hc128765e},
  {32'h434603f0, 32'h41d96cd7, 32'h41bddd40},
  {32'h4386e8e0, 32'h43849a21, 32'h42998249},
  {32'hc4bb54b1, 32'hc3e33a07, 32'hc3036087},
  {32'h42b37278, 32'h438f16d7, 32'hc389d603},
  {32'hc4a1970a, 32'h43998e5b, 32'h438712f5},
  {32'h4514f93c, 32'hc231265f, 32'hc259ae47},
  {32'hc45fea38, 32'hc3a55449, 32'hc2f6aa0c},
  {32'h44e88e8b, 32'hc36c186a, 32'hc2a71c82},
  {32'hc4644d25, 32'h4375fcb5, 32'h4365eec8},
  {32'h448461ca, 32'h432a7824, 32'h4426b842},
  {32'hc516fde9, 32'h43a315ea, 32'hc304a49b},
  {32'h44c685aa, 32'hc3b87a55, 32'h43792254},
  {32'hc50d6a89, 32'h4359d806, 32'h431485b0},
  {32'h44e32040, 32'hc2c7ff11, 32'hc2f8989d},
  {32'hc4544abc, 32'hc4131481, 32'h42869b32},
  {32'h44f7b2ca, 32'hc3238332, 32'h42f04957},
  {32'hc3048b93, 32'hc37a5ff5, 32'h432151bd},
  {32'h44d1aee8, 32'h42df6e09, 32'hc3520ae1},
  {32'hc4ce5a40, 32'hc1134cd4, 32'h41272f76},
  {32'h441f4d20, 32'hc3d9250c, 32'hc0860df8},
  {32'hc4c235b5, 32'hc3ad3b56, 32'h43857f50},
  {32'h4510e9cb, 32'hc2506aaf, 32'h438ee1e9},
  {32'hc4e82dc2, 32'h4382ae5c, 32'h43480ebf},
  {32'h44b0e4be, 32'hc30b6ab3, 32'hc33f45ce},
  {32'hc431e125, 32'h42de4df9, 32'hc2cf880a},
  {32'h44a72aa6, 32'h40eb8700, 32'hc334e31f},
  {32'hc4819c6c, 32'h408bc4ef, 32'h4373da32},
  {32'h442aab20, 32'hc2d35755, 32'hc32f3e09},
  {32'hc49f0f82, 32'hc035b7b4, 32'hc3a7947c},
  {32'h4507933e, 32'hc406b996, 32'hc294cab6},
  {32'hc4ed2bce, 32'hc36962ec, 32'h4308845a},
  {32'h4488534e, 32'h4291d73e, 32'hc33101ea},
  {32'hc4424214, 32'hc2eae8fe, 32'hc2c76c6c},
  {32'h440f3ab4, 32'h42e3cd39, 32'hc35f2cfe},
  {32'hc485ca0f, 32'hc37e0733, 32'h435bb026},
  {32'h4306cc9a, 32'hc13ca59a, 32'h4344f12c},
  {32'hc4f9f87d, 32'hc320e2ed, 32'h4316ed35},
  {32'h44dd3dd3, 32'h433da7af, 32'hc36aaa6d},
  {32'hc4c511c6, 32'h431b5423, 32'hc2b281c7},
  {32'h4510c2b1, 32'h4287bf06, 32'hc2924c76},
  {32'hc4473503, 32'hc2eece86, 32'h4230a17a},
  {32'h4421e1c8, 32'hc39af3f9, 32'hc253098e},
  {32'hc4e7e7ac, 32'h42a6eedf, 32'h42f6c090},
  {32'h443925c1, 32'h430d0ce1, 32'hc1dc0c7c},
  {32'hc5089dbe, 32'h4391a57a, 32'h436770ec},
  {32'h44de40f6, 32'hc2dafbbe, 32'hc2aba638},
  {32'hc4f12f6e, 32'h42826f66, 32'h43563111},
  {32'h4506422f, 32'hc3d50cfc, 32'hc37d2243},
  {32'hc49ca810, 32'h4355626f, 32'h418eab62},
  {32'h44b90080, 32'h427eaca2, 32'hc38a1f03},
  {32'hc4af5ae8, 32'h43eeaee1, 32'hc259917d},
  {32'h44317152, 32'h420f8f3d, 32'h432bcf4f},
  {32'hc4dea8ac, 32'h43ef3887, 32'h421207a9},
  {32'h44db9d54, 32'hc188b6a4, 32'hc288ad6d},
  {32'hc3ffa410, 32'h43aedb8b, 32'hc35ecc69},
  {32'h44a558a0, 32'hc3292401, 32'hc3b1edf1},
  {32'hc4d274aa, 32'hc272ab79, 32'h42871803},
  {32'h450f8568, 32'h432dae6d, 32'h438e30b6},
  {32'hc5095c2e, 32'h434d98f5, 32'h42bed9fc},
  {32'h449ea8ae, 32'hc39e9ed6, 32'hc206f571},
  {32'hc4c4985e, 32'h43b4a037, 32'h439f01b4},
  {32'h434816dc, 32'h439d6550, 32'hc392ee44},
  {32'hc4f0b761, 32'hc2c4ee64, 32'hc37f83bf},
  {32'h450abda1, 32'hc380ca5d, 32'h42dc7c7b},
  {32'hc4922de2, 32'h4396fb62, 32'h4389dc3f},
  {32'h4442fd77, 32'hc36ef3f8, 32'h42c4df46},
  {32'hc2bd2bc0, 32'hc3ab8070, 32'h42ec861e},
  {32'h4495bb56, 32'h43a74ff1, 32'hc379038a},
  {32'hc3631f5e, 32'hc28fc9c5, 32'h437c8767},
  {32'h43253140, 32'hc2aac040, 32'hc358d5e0},
  {32'hc4b24855, 32'hc1e3fb06, 32'h41d476f7},
  {32'hc246bbc0, 32'h42cacfaf, 32'h40f01899},
  {32'hc42c3384, 32'hc3bbfbb1, 32'hc3f663fb},
  {32'h4504b787, 32'h433751ad, 32'h42efaae9},
  {32'hc48c65f6, 32'hc24c9ef2, 32'h4388d4ed},
  {32'h42a30b98, 32'hc3a5291c, 32'hc365ceb8},
  {32'hc4fb79a6, 32'h420781bc, 32'hc356269a},
  {32'h43b4f33c, 32'h426ceffa, 32'h42a5b919},
  {32'hc4bde6de, 32'h4344e7ee, 32'h42f7fbcc},
  {32'h448cf898, 32'h420baf33, 32'h43093fea},
  {32'hc4c2f3be, 32'hc2e4ddb3, 32'h43e137f2},
  {32'h44848516, 32'hc20f1c0c, 32'h434ee5ce},
  {32'hc4ca1318, 32'h43dbc065, 32'h4294fd2b},
  {32'h44fd52ab, 32'h42905c08, 32'hc4020d1f},
  {32'h42bf0ece, 32'hc2e37af0, 32'hc19ad871},
  {32'h44a84708, 32'h416ce377, 32'hc1387c71},
  {32'hc4d69b6b, 32'h43e6a39a, 32'h42fa9ab3},
  {32'h44a0aacd, 32'hc1c15426, 32'h42d318a7},
  {32'hc462da19, 32'hc2f3ceaf, 32'h43f6fdea},
  {32'h44c068f6, 32'h42c81ce9, 32'hc3537f19},
  {32'hc40b49e6, 32'h43a2a0ca, 32'hc23be768},
  {32'h448fed5d, 32'hc2e22a92, 32'hc380f753},
  {32'hc48ab390, 32'hc378448c, 32'hc101d52e},
  {32'h43d4a5a6, 32'hc3008724, 32'hc4127bc3},
  {32'hc3d5358e, 32'hc2ca38ba, 32'h4383f4b3},
  {32'h44a0f540, 32'h434794cf, 32'hc30520ac},
  {32'hc3d311a0, 32'h431df7e6, 32'h42de9b48},
  {32'h450f25b5, 32'h42f8e77d, 32'hc34c9f40},
  {32'hc486b968, 32'h4153ecd8, 32'hc31c86e6},
  {32'h43d69f16, 32'hc29f0ba2, 32'h429943d9},
  {32'hc4c38931, 32'hc3847847, 32'hc0b5dd7a},
  {32'h450760bc, 32'hc1e4d3d7, 32'hc213489b},
  {32'hc4d5c3fe, 32'h4014b82c, 32'h42b3a812},
  {32'h435fce18, 32'h41b3adc5, 32'hc35db3cf},
  {32'hc4cc64ff, 32'h43e81696, 32'h434be7ae},
  {32'h446e5c9a, 32'h43e39f59, 32'hc368f75b},
  {32'hc4f0210b, 32'hc25c566d, 32'hc307904b},
  {32'h44f46d23, 32'hc38703ff, 32'h4272579c},
  {32'hc447a7f8, 32'hc363fa71, 32'h43a503ba},
  {32'h45074358, 32'h42966705, 32'h42e21c84},
  {32'hc517c2ed, 32'hc1b7236e, 32'hc1f2e978},
  {32'h44f8149b, 32'hc2b82ed7, 32'h429063fc},
  {32'hc48f7d56, 32'h4111933a, 32'h4418253d},
  {32'h4443b368, 32'h40b5637e, 32'h43b721c7},
  {32'hc520faba, 32'hc35095ca, 32'h43585b8d},
  {32'h44019a9c, 32'hc3157888, 32'h4308baa6},
  {32'hc504cf02, 32'h41a3336a, 32'hc389a2ab},
  {32'h45082ca6, 32'hc36f1475, 32'h43b889d8},
  {32'hc4a1adcb, 32'hc30903f4, 32'h422a5d50},
  {32'h450330d4, 32'h42a5388b, 32'hc22b5918},
  {32'hc5057548, 32'hc2b75665, 32'hc31ea0c0},
  {32'h43c16e5b, 32'hc32f1ec0, 32'hc2820130},
  {32'hc4e2894e, 32'h4388c30d, 32'h438af0da},
  {32'h44937c5d, 32'hc3754d2b, 32'h4310242b},
  {32'hc425f254, 32'hc34da84d, 32'hc3a8384c},
  {32'h44feb289, 32'hc3ef95f4, 32'h41c40c94},
  {32'hc4b00957, 32'h44128180, 32'h43bdea2e},
  {32'h44c57d48, 32'hc2a9ac05, 32'hc400c085},
  {32'hc3757aa5, 32'h439a886d, 32'hc315bcc8},
  {32'h44f24469, 32'hc28bec92, 32'h43e06ff1},
  {32'hc4fc8aad, 32'hc3888ed1, 32'h443591dc},
  {32'h445806bc, 32'h42853182, 32'hc18e3ddc},
  {32'hc3c6a2b2, 32'hc42331ed, 32'hc2f291eb},
  {32'h45198beb, 32'hc3034983, 32'h430772fd},
  {32'hc4361824, 32'h422ab41e, 32'h439fa498},
  {32'h4265c1b0, 32'hc32eb865, 32'hc3bdfa09},
  {32'hc34e7780, 32'h430e1883, 32'hc33afb06},
  {32'h44e161c6, 32'hc1976a14, 32'h42438582},
  {32'hc508caee, 32'h42801a2a, 32'hc324a3b2},
  {32'h42167f70, 32'h4305a7fb, 32'hc2c8fb8a},
  {32'hc4b8d0ed, 32'h43f071e2, 32'hc3a92283},
  {32'h448e8b3c, 32'h431dad37, 32'hc2fe71d7},
  {32'hc4d89ab5, 32'hc3b623e6, 32'hc3c640b0},
  {32'h44bc0b36, 32'h43fd3269, 32'hc3463adb},
  {32'hc5055d49, 32'hc32b20c3, 32'hc2b830b0},
  {32'h4465500e, 32'hc305b11a, 32'hc30fd202},
  {32'hc507e14a, 32'hc2b5e51b, 32'h4345cbbd},
  {32'h44e2ad4e, 32'h4346a11a, 32'hc3277a1f},
  {32'hc4efd81c, 32'h42e51eda, 32'hc232ce9a},
  {32'h44b4d1a4, 32'hc36cb595, 32'hc38abcaf},
  {32'hc48bfd59, 32'hc28f028f, 32'h4390ea23},
  {32'h44fcbfde, 32'h42da761b, 32'h433922b6},
  {32'h42b6f1b1, 32'h42cd30fc, 32'h437d2628},
  {32'h43de93ac, 32'h435542ba, 32'hc1aa489c},
  {32'hc2340ec0, 32'h423437cd, 32'h4250e55c},
  {32'h449d6a74, 32'hc2d60cc0, 32'h426b614a},
  {32'hc5129174, 32'h4161f02b, 32'hc2047e00},
  {32'h43e0d694, 32'hc2cc209d, 32'h4318ef0f},
  {32'hc4002099, 32'hc347f165, 32'h421f4a41},
  {32'h450dbdeb, 32'hc304bfb9, 32'h429fb900},
  {32'hc39a2bb6, 32'hc208b94f, 32'h41c5b9a6},
  {32'h4485cd96, 32'h430441f9, 32'h40c79dbb},
  {32'hc52530f8, 32'hc281901e, 32'h424a2640},
  {32'h4461f436, 32'h421303e0, 32'hc223d08b},
  {32'hc48f8db5, 32'h433f5428, 32'hc2d9583f},
  {32'h450c25ba, 32'hc3431b3b, 32'h433bb4eb},
  {32'hc5156b0f, 32'hc39f597c, 32'hc30cc4ac},
  {32'hc3be59e8, 32'hc34df716, 32'h42551557},
  {32'hc4ce10e8, 32'h43bc8402, 32'h43755e84},
  {32'h441f8f45, 32'h4294d302, 32'hc1452a5b},
  {32'hc502049c, 32'h433566e9, 32'h435033b8},
  {32'h44c3cf1e, 32'h42060964, 32'h43990e6c},
  {32'hc4610bfa, 32'h4258a0ae, 32'h424abdc0},
  {32'h41f56020, 32'h42b1b0b6, 32'hc35f4d1a},
  {32'hc4b835ec, 32'h4387b692, 32'h4325fcf0},
  {32'h4508df5d, 32'h437cd5e8, 32'h4383ef10},
  {32'hc4e06234, 32'hc32f6a9d, 32'hc2e4957c},
  {32'h442b90c8, 32'hc23f86ee, 32'hc2daa3ac},
  {32'hc502e98d, 32'hc3356712, 32'hc39cb524},
  {32'h44e73f14, 32'hc2f036da, 32'hc2d5f00f},
  {32'hc4a8d380, 32'hc38e806d, 32'hc36f444a},
  {32'h43cc4acc, 32'hc2e2712d, 32'h431dbf4d},
  {32'hc46c55e9, 32'h425f2a82, 32'h4248a6e7},
  {32'h449bd474, 32'hbe197b58, 32'h3ce324df},
  {32'hc4e4cbea, 32'hc3112d75, 32'h42e8bafd},
  {32'h4520b308, 32'hc2b70fa9, 32'hc1beaa95},
  {32'hc5138924, 32'hc2bbdfaf, 32'h41cc2808},
  {32'h4430415a, 32'h41a9b255, 32'h435314b1},
  {32'hc4810381, 32'h42515f8e, 32'hc3837b3b},
  {32'h44af76a4, 32'h42025058, 32'h4246b60e},
  {32'hc4160720, 32'hc36435d1, 32'hc370b708},
  {32'h44958ea4, 32'hc30f91fa, 32'h41623e42},
  {32'hc4d49b72, 32'h41bf0c64, 32'hc30501c2},
  {32'h450b4f42, 32'h43347ee9, 32'h426094d5},
  {32'hc468bc19, 32'h4284c6d5, 32'h43c27f3f},
  {32'h451d2edc, 32'hc4055022, 32'hc333ad0a},
  {32'hc4e5be61, 32'h42b35d3d, 32'hc2ef548c},
  {32'h44a9b8d1, 32'h4392bbde, 32'hc2d4fd2c},
  {32'hc2944fab, 32'h42acb905, 32'hc1731c69},
  {32'h450f12bd, 32'hc2dccec4, 32'h42abdf10},
  {32'hc482d119, 32'hc39c617f, 32'hc2904b13},
  {32'h450c8307, 32'hc2e843b8, 32'hc193f9b1},
  {32'hc484ac68, 32'hc30ad84b, 32'h430bac30},
  {32'h44c9c827, 32'h43651b5b, 32'h42dedcbc},
  {32'hc45df680, 32'h4309ceca, 32'hc325170a},
  {32'h443f8994, 32'hc301218b, 32'h437128fd},
  {32'hc3a256c2, 32'hc1ed7b9e, 32'h4247ddc0},
  {32'h44d87aee, 32'hc2ab1007, 32'hc2d6b95c},
  {32'hc4e4a7e6, 32'h43bb141f, 32'h43f9e6ce},
  {32'h44d0d298, 32'hc3224df4, 32'h439a59b4},
  {32'hc519f5fb, 32'hc32178b8, 32'hc3098dcc},
  {32'h44cc0d70, 32'hc2c0acca, 32'hc380513b},
  {32'hc4c457f3, 32'hc380e3ef, 32'h43334326},
  {32'h442e4c2d, 32'hc3ad6c89, 32'hc389fdff},
  {32'hc4e74dcd, 32'h4343a1d9, 32'hc3276bcb},
  {32'h4419e0d0, 32'h402e80fd, 32'h43453f61},
  {32'hc443fd3f, 32'hc28b44f8, 32'hc2e868b2},
  {32'h4463328c, 32'h40f8bb77, 32'hc3821a7b},
  {32'hc4ac8e39, 32'h437e12cf, 32'hc30ec5f3},
  {32'h43c0e430, 32'h42f9767e, 32'h435f4248},
  {32'hc4a15896, 32'h41b81782, 32'hc36c0945},
  {32'h44c4252c, 32'hc3034564, 32'hc2cb933c},
  {32'hc512cb2b, 32'hc3ac33c8, 32'hc2cc4e6c},
  {32'h44e56ede, 32'h427496a6, 32'hc3756919},
  {32'hc3951e68, 32'h43561966, 32'h43534a91},
  {32'h44be4b31, 32'h433fcf95, 32'h43a1895c},
  {32'hc4156792, 32'hc31a59fb, 32'h41d43f8a},
  {32'h443242f0, 32'hc2d19ec1, 32'h4326b44d},
  {32'hc466612a, 32'hc3811427, 32'hc3498968},
  {32'h44f2d4d7, 32'h43a65e30, 32'h43a08a23},
  {32'hc4585a72, 32'h434b0cb5, 32'h434eb54b},
  {32'h44f54ae3, 32'h431703cc, 32'hc20fc321},
  {32'hc4d3a39a, 32'h42f1cc30, 32'hc28586b4},
  {32'h450463bd, 32'hc3c053e6, 32'h43a8157c},
  {32'hc436e56e, 32'hc37ddbbd, 32'hc346d9c3},
  {32'h448da577, 32'hc38827eb, 32'hc201358b},
  {32'hc425b310, 32'hc1a6f8f1, 32'hc3b0168c},
  {32'h4436b27a, 32'h43c0d96c, 32'hc2ca2f06},
  {32'hc4dcdd84, 32'h434355bb, 32'hc32306e2},
  {32'h450184aa, 32'hc24aa6f8, 32'h40611a58},
  {32'hc4372f04, 32'hc3d43d94, 32'h427c87c6},
  {32'h43955920, 32'h42560a7e, 32'h438c1720},
  {32'h43402533, 32'h4318bc8d, 32'hc3bed128},
  {32'h42ef28a0, 32'hc42a1aab, 32'hc3928eaf},
  {32'hc4a4ff13, 32'hc363373b, 32'hc41d15c6},
  {32'h44a5d09d, 32'h42a3e493, 32'hc3977fa0},
  {32'hc4dbad46, 32'hc20e6b90, 32'hc3986839},
  {32'h42b7a4f0, 32'hc0514ee3, 32'hc3eb291c},
  {32'hc487838e, 32'hc4047682, 32'h3f16a5e4},
  {32'h4417efe3, 32'h43829dae, 32'h4362f13e},
  {32'hc4c92eef, 32'hc2f46c3e, 32'hc3b7b484},
  {32'h448186f8, 32'hc2623caf, 32'hc29f97ec},
  {32'hc3fcfbf4, 32'hc372e39d, 32'hc3bc61e2},
  {32'hc42e3a48, 32'hc2915963, 32'h43397942},
  {32'h42962dd2, 32'h4214cd09, 32'h43ca36d2},
  {32'hc467da43, 32'hc3362ecd, 32'hc2a39e85},
  {32'h4357ad18, 32'h43a251a8, 32'h42f6ae92},
  {32'hc4858f4f, 32'hc2b3035f, 32'h427e45c8},
  {32'h44b45d31, 32'h4374493c, 32'h4270130a},
  {32'hc4194396, 32'h4319a59b, 32'hc1ec237e},
  {32'h4502f9e4, 32'hc3b18692, 32'h433f6cb0},
  {32'hc48495f0, 32'hc20bda60, 32'h43c51f62},
  {32'h44a55d72, 32'hc39be8aa, 32'hc3349d98},
  {32'hc4d2524f, 32'h42bc5290, 32'hc3bbe054},
  {32'h448a4fe7, 32'h430eae72, 32'h42b02aa6},
  {32'hc2c3bf00, 32'h4337b78a, 32'hc39d0a9d},
  {32'h44861604, 32'hc343996e, 32'h4363f4da},
  {32'hc495e702, 32'hc2a81e5c, 32'hc36653ef},
  {32'h44f9c610, 32'hc32dee7f, 32'h421264df},
  {32'hc500b29f, 32'hc3328425, 32'hc3d796e2},
  {32'h44f850ff, 32'h43e548a7, 32'hc27b87f1},
  {32'hc19ba940, 32'h439f1b92, 32'hc39a3b54},
  {32'h444d8ffd, 32'hc35ff458, 32'hc272d07b},
  {32'hc501a0c5, 32'h42cd04fc, 32'hc31c2d8c},
  {32'h44ffe147, 32'h4436d804, 32'hc3205639},
  {32'hc4e24818, 32'hc30a89ea, 32'h4321ecaf},
  {32'h44a1c7b6, 32'h427d4b29, 32'h42285776},
  {32'hc3460180, 32'h4162b5a5, 32'h42d43801},
  {32'h44296000, 32'hc212074f, 32'hc1ad3116},
  {32'hc4ecf291, 32'hc1f6bad4, 32'h42f1add6},
  {32'h449cd722, 32'hc24408a6, 32'h4407e1a5},
  {32'hc41a77d4, 32'h419c8184, 32'hc2495528},
  {32'h44da0102, 32'h4219f2be, 32'hc36e8250},
  {32'hc496ab74, 32'h42b15c09, 32'h43912b60},
  {32'hc354ae44, 32'hc3aab36e, 32'hc3069743},
  {32'hc44e3b02, 32'h41658c01, 32'hc32eef25},
  {32'h43a265b4, 32'hc3442b26, 32'hc338b6b3},
  {32'h42d9b8ba, 32'hc342e2d3, 32'hc35f6c57},
  {32'h44f1cb03, 32'hc3c9d03b, 32'h43478a37},
  {32'hc4204288, 32'hc32f6257, 32'hc3328d93},
  {32'h44fb55fe, 32'hc2adedd1, 32'h42c0bd09},
  {32'hc3b33dd0, 32'hc400a4e3, 32'hc257f0fe},
  {32'h44961dec, 32'h435afea2, 32'hc296bd51},
  {32'hc510ccee, 32'h42cb482a, 32'h438225d9},
  {32'h44b401cc, 32'hc2889933, 32'h43a62666},
  {32'hc4137570, 32'hc37dfa19, 32'h42c5fe35},
  {32'h45063c74, 32'h3fbcc42c, 32'h426403a4},
  {32'hc47deeb8, 32'hc1940efe, 32'h43a6fcd3},
  {32'h42b44670, 32'h42e6365f, 32'hc1f30941},
  {32'hc47ea904, 32'h4190284e, 32'h43198468},
  {32'h44a33c34, 32'h437906d7, 32'h43ec2034},
  {32'hc4e0d95b, 32'hc185fcdc, 32'h429f6262},
  {32'h44a2f16a, 32'hc299059a, 32'hc33e573a},
  {32'hc38f29a0, 32'h439ce298, 32'hc3b44bfd},
  {32'h44229b7a, 32'hc0afa812, 32'h41359616},
  {32'hc4e292a9, 32'hc21c186a, 32'hc28641c6},
  {32'h44c9b0c6, 32'h424e97c0, 32'hc1a674d1},
  {32'hc4174606, 32'h4247790b, 32'hc365b2c9},
  {32'h446e35e2, 32'h4286af03, 32'h43747b09},
  {32'hc4c0905d, 32'h42965d15, 32'hc3045cd5},
  {32'h44a2652f, 32'h42f038e8, 32'h42592eba},
  {32'hc42671d9, 32'hc32f933c, 32'h42fb1c5e},
  {32'h44481f6a, 32'hc33fcfdc, 32'h426b902d},
  {32'hc4959f00, 32'hc3456619, 32'hc3209dd4},
  {32'h44346a48, 32'h42f6e2c0, 32'hc3ec39c3},
  {32'hc4af4a0e, 32'hc2dea738, 32'hc2c2024e},
  {32'h447ed709, 32'h41524e32, 32'h43ce0328},
  {32'hc4fccdc1, 32'h426ee4b1, 32'hc39a4a41},
  {32'h44385454, 32'h41988197, 32'h426e4c71},
  {32'hc46fb325, 32'hc2ca388f, 32'hc2bcbc84},
  {32'h44b7affa, 32'h41d16ee5, 32'h42595fd3},
  {32'hc50aecc9, 32'hc3037955, 32'hc3894b93},
  {32'h44702073, 32'hc32e557a, 32'hbfb81c80},
  {32'hc394a2cc, 32'hc03ae6b8, 32'h42b96595},
  {32'h4509ed98, 32'hc2f6d9ce, 32'h43641057},
  {32'hc49f3e0e, 32'hc2fe391f, 32'h43127219},
  {32'h41e9c800, 32'h42809070, 32'hc31a0d31},
  {32'hc4aaabee, 32'hc3901db7, 32'hc2d644f5},
  {32'h44b81d06, 32'h43509d22, 32'hc3a4e0eb},
  {32'hc356e7d0, 32'hc37c2e92, 32'h41c85274},
  {32'h44383a68, 32'hc1ccce27, 32'h430b0dbb},
  {32'hc5003d84, 32'h43225f4b, 32'h4353be83},
  {32'hc2d0d2f0, 32'hc3afaee2, 32'hc3dc056e},
  {32'hc4d8ef00, 32'hc30a36c6, 32'hc410516c},
  {32'h440943a9, 32'h42a431e9, 32'h439af35f},
  {32'hc50dd8e1, 32'h42a4fd3e, 32'h4328f89d},
  {32'h4428512a, 32'h43538fac, 32'hc2206136},
  {32'hc4d3d2ed, 32'h43a2bfaf, 32'hc2485d75},
  {32'h44e1a81f, 32'h43467249, 32'hc18feb75},
  {32'hc502ae7e, 32'hc3194c96, 32'h41bda990},
  {32'h44eadc38, 32'h4357e729, 32'hc2052bca},
  {32'hc4fdcd50, 32'hc3e40a4e, 32'h43aeed99},
  {32'hc3219568, 32'h43b145b9, 32'hc321f23d},
  {32'hc40c4f61, 32'hc288f37a, 32'hc336a406},
  {32'h451d1560, 32'hc2cbb1a8, 32'hc2bbd17f},
  {32'h41b1adf0, 32'h423a3a3c, 32'hc390e88a},
  {32'h4420f1e2, 32'hc3a40756, 32'h42a36b29},
  {32'hc4e31d0e, 32'h434020a0, 32'hc37ea161},
  {32'h44602831, 32'h43830e7e, 32'h422496e6},
  {32'hc350b9be, 32'hc26dc775, 32'h42957b27},
  {32'h43031130, 32'hc405c7da, 32'hc300a191},
  {32'hc4879ca8, 32'h438a75bf, 32'h438b703f},
  {32'h449ca815, 32'h41c4eed7, 32'hc28ed47c},
  {32'hc40a2e44, 32'hc39e3742, 32'h4365e29e},
  {32'h440767e2, 32'hc3172a27, 32'h431d9d4b},
  {32'hc5054a8b, 32'hc319e618, 32'hc3828de4},
  {32'h44c6bd56, 32'h43526978, 32'h42bc0860},
  {32'hc4710f0f, 32'hc23d3c65, 32'h43adf33a},
  {32'h44a5b52f, 32'hc3402efe, 32'h42fcda70},
  {32'hc4c65c52, 32'hc1ef12ef, 32'h424a38c7},
  {32'h44c64283, 32'hc198b7a3, 32'hc2e3eb6c},
  {32'hc4302824, 32'hc37b6cfe, 32'h43166962},
  {32'h43e962ca, 32'h43ce655d, 32'hc23b1820},
  {32'hc4bc931e, 32'hc2d4bc0d, 32'hc33bf260},
  {32'h44ad1264, 32'hc1710085, 32'h427973bc},
  {32'hc41dad1e, 32'hc35e0ab0, 32'h4388a094},
  {32'h44f58c05, 32'hc1d4dfdf, 32'hc2a9b179},
  {32'hc50626fc, 32'hc3e6592e, 32'h4308022a},
  {32'h43f4f198, 32'hc426f268, 32'hc3a1551d},
  {32'h44c4d0a0, 32'h423ef572, 32'hc377ebb9},
  {32'hc38a4244, 32'hc31d3ee3, 32'h42ec5df0},
  {32'h4505363e, 32'hc3a0b6a5, 32'hc3ff200b},
  {32'hc3cdeab4, 32'h4234b254, 32'h4229a38e},
  {32'h448422f4, 32'h42f0894a, 32'h43eaa87c},
  {32'hc3fa95f0, 32'h433f7e15, 32'h40c4e730},
  {32'h451ed822, 32'hc3dedd0f, 32'h43682a6a},
  {32'hc4c1578b, 32'h4304b37d, 32'hc3c21c35},
  {32'h4420072c, 32'hc18f2d7e, 32'h438e664c},
  {32'hc3dfb54a, 32'h41914fcd, 32'hc34a539a},
  {32'h450450b6, 32'hc4298be6, 32'h42917948},
  {32'hc49b5e6e, 32'h43910ae3, 32'h43a14324},
  {32'h44f0dc99, 32'h4296c890, 32'hc2b5d158},
  {32'hc4434d71, 32'hc2d22163, 32'hc344850a},
  {32'h44f433dc, 32'hc171dd68, 32'h43d523f0},
  {32'hc4127c88, 32'h43c6a8f3, 32'h43a0e89a},
  {32'h442fda1c, 32'hc37d90cd, 32'h43947eac},
  {32'hc48fda6e, 32'hc32a0674, 32'h43c40fe3},
  {32'h43d0a464, 32'hc24e8e47, 32'hc3d637a4},
  {32'hc3e203b0, 32'hc2bb4724, 32'h4367cc00},
  {32'h4495b542, 32'h42a053fa, 32'h425eaa65},
  {32'hc377ff7c, 32'h40f59a4a, 32'h431d3ca1},
  {32'h452351b5, 32'h42b42799, 32'hc0e142b1},
  {32'h4335111a, 32'hc35ae8ba, 32'h4226ab89},
  {32'h44d9c5a3, 32'h4415b691, 32'h434f1aa5},
  {32'hc43aafc4, 32'h42172b61, 32'hc351ef73},
  {32'h449e4c65, 32'hc36f75a6, 32'h42cf5fe5},
  {32'hc4e913e5, 32'hc3992bdc, 32'hc314bde2},
  {32'h439115f4, 32'hc0c733a2, 32'h42dfe329},
  {32'hc49f821d, 32'h4402f1fd, 32'hc31e472c},
  {32'h4415c478, 32'h43882fa2, 32'h426fe07c},
  {32'hc4cdc81c, 32'hc26beb7f, 32'hc2029efb},
  {32'h44f587d2, 32'hc29b6921, 32'h42849d05},
  {32'hc3ec1ade, 32'hc31b5512, 32'hc2811b71},
  {32'h44bffc6b, 32'hc2c9b4f9, 32'hc3a72b98},
  {32'hc31d4cb8, 32'hc38decc1, 32'hc32f4aa8},
  {32'h44a6810a, 32'h4397474a, 32'h43a0c115},
  {32'hc4ed9d92, 32'hc3a616e0, 32'hc290664c},
  {32'h439be62e, 32'h43d55c8f, 32'h42c961c0},
  {32'h42d7f9a0, 32'hc3269d1c, 32'hc2f61200},
  {32'h42c41290, 32'h4288c9d8, 32'h423bbcf3},
  {32'h42b1b732, 32'hc384cf70, 32'hc2d76a0f},
  {32'h4514103c, 32'h4386a58b, 32'hc37b46ed},
  {32'hc28a0189, 32'hc13e7f2a, 32'hc38e6ab3},
  {32'h44e57d36, 32'hc2eb3ed1, 32'hc3b1d9fd},
  {32'hc41fffc0, 32'hc37c2546, 32'h42ac502c},
  {32'h43f50928, 32'h42381902, 32'h41de0efa},
  {32'hc509c6a1, 32'hc37322ca, 32'h42df7011},
  {32'h43ad35b8, 32'hc35cc1b1, 32'hc316f42e},
  {32'hc4650e26, 32'h42ad7b37, 32'h430b9446},
  {32'h44d3a0b8, 32'h42aba40b, 32'hc2c7fee3},
  {32'hc4f8691e, 32'hc2a9d8f9, 32'h41e91cd2},
  {32'h449c6d7a, 32'h4363cb91, 32'h43efb9f1},
  {32'hc379f6a5, 32'h437af853, 32'h43039b95},
  {32'h4495f063, 32'hc3825c4a, 32'hc321cf69},
  {32'hc4a56394, 32'h43c1aab6, 32'h4376c386},
  {32'h447d5b24, 32'hc3ea71af, 32'hc246a7b7},
  {32'hc4e69825, 32'hc2299316, 32'hc383221f},
  {32'h44e09cee, 32'h429a4692, 32'hc287a580},
  {32'hc44bbd8b, 32'h432f81f1, 32'hc311f50f},
  {32'h4499171b, 32'h431e42ae, 32'hc3608574},
  {32'hc48b9a5b, 32'hc2b2e47c, 32'hc34c4305},
  {32'h44966dde, 32'h427b999c, 32'hc3bc083b},
  {32'hc4347ab1, 32'hc311c203, 32'hc3261fb5},
  {32'h44b97ab3, 32'hc33f750b, 32'h3f839f88},
  {32'hc4c4ceb4, 32'hc396fb7a, 32'hc3894cba},
  {32'h4482193f, 32'h43744bac, 32'h4310c60c},
  {32'hc46989ca, 32'h441cc2b2, 32'hc3b1d4ed},
  {32'h43c1e274, 32'hc2927964, 32'hc2f5c079},
  {32'hc508f697, 32'hc392ae24, 32'h41261d48},
  {32'h44027050, 32'h4315adf1, 32'hc2bccf07},
  {32'hc4355cc5, 32'hc2c5d52f, 32'hc2c86589},
  {32'hc284c1a0, 32'h4321f6a6, 32'h428d4724},
  {32'hc2242a8c, 32'h430a77ce, 32'h429a989c},
  {32'h44938129, 32'h43ef5b67, 32'h436587e2},
  {32'hc4aec4c7, 32'h42d60e87, 32'hc2a7cb3e},
  {32'h442169e0, 32'h42318ea8, 32'hc2c6f8ba},
  {32'hc4981df6, 32'h42f55828, 32'hc3250c68},
  {32'h44edc58d, 32'hc3664dc2, 32'hc316d952},
  {32'hc50a7c0e, 32'h4353b4ad, 32'hc314a457},
  {32'h44c680df, 32'hc22fc91b, 32'h4123d3ac},
  {32'hc4d1c95a, 32'hc2239efb, 32'h41e77929},
  {32'h44d355a5, 32'hc3b634e7, 32'h436411c9},
  {32'h43adcd64, 32'h43af510c, 32'h4059be79},
  {32'h451beb14, 32'h434de45f, 32'h44019c66},
  {32'hc4959822, 32'hc369cf18, 32'hc319f6ea},
  {32'h44b9d9be, 32'h4308259b, 32'h429c9319},
  {32'hc471d4a0, 32'h422b842b, 32'h403a8cac},
  {32'h442403f2, 32'h432ce3ec, 32'h42f0cada},
  {32'hc3ddd450, 32'hc2ddef74, 32'hc2eddd41},
  {32'h44bf7914, 32'hc28fb2e5, 32'h4126d056},
  {32'hc4c867ba, 32'h434096b7, 32'hc3c4e535},
  {32'h43f6ac08, 32'h42bb30da, 32'hc3928d10},
  {32'hc3973f18, 32'h436033c4, 32'h432430e7},
  {32'h44676b5e, 32'h430b8721, 32'hc309730f},
  {32'hc48c7bd1, 32'h43619680, 32'h42ae2523},
  {32'h44f30806, 32'h41ae07e3, 32'h42e868d6},
  {32'hc3f2c591, 32'h4307361a, 32'hc3613b6b},
  {32'h4463c8ce, 32'h4353e2b5, 32'h431d717a},
  {32'hc46e7583, 32'hc301f20f, 32'hc3090089},
  {32'hc338eba8, 32'h4332eb8a, 32'h43c78585},
  {32'hc48eee8c, 32'h41aec820, 32'hc0ec4358},
  {32'h44ad78e4, 32'h4185e7f0, 32'h43429cb7},
  {32'hc43dbe92, 32'hc3d864ca, 32'h430e6e07},
  {32'h44366714, 32'h428708a9, 32'hc31bec13},
  {32'hc4e36ff6, 32'h4303cf80, 32'hc3356e7c},
  {32'hc23b3ea0, 32'h43329dbb, 32'h42edb506},
  {32'hc42bd8b6, 32'hc3bb8d79, 32'h4356915e},
  {32'h44a20964, 32'h41bd1fff, 32'hc31e8fd2},
  {32'hc4fb901c, 32'hc309b007, 32'h42f8ce04},
  {32'h44ddc56f, 32'h42f5e5d5, 32'hc38ddee2},
  {32'hc341ca41, 32'hc3bb790b, 32'h4388235d},
  {32'h44624459, 32'h430952a5, 32'hc318cff2},
  {32'hc4f6f5e6, 32'h42b78455, 32'hc284f360},
  {32'h44e53012, 32'hc2b5f266, 32'h4243c417},
  {32'hc4fe92c6, 32'h42a35366, 32'hc318a489},
  {32'h441b078a, 32'hc3672e7d, 32'h418691e8},
  {32'hc328c543, 32'hc1ee1345, 32'hc09f89e2},
  {32'h450b026c, 32'hc3506d94, 32'h439a63a2},
  {32'hc40128fc, 32'h437b58ac, 32'hc399c3b5},
  {32'h449cf77a, 32'h43539e1a, 32'h428c5c39},
  {32'h42b90f72, 32'hc2f0bde4, 32'h42eb030d},
  {32'h448a77bc, 32'hc2ea996b, 32'hc2ff90da},
  {32'h43ce2d78, 32'h430585b6, 32'hc35ee1e5},
  {32'h4485aacf, 32'h428a82a3, 32'h40952470},
  {32'hc4d51022, 32'h435e6991, 32'hc2aaeb5e},
  {32'h4503002f, 32'hc39b9ffe, 32'hc351bf6e},
  {32'h401413c8, 32'hc0fdcd26, 32'h4313d7d8},
  {32'h43c1e790, 32'h4347fc30, 32'h43f40bbe},
  {32'hc50cfcd9, 32'h42c5c542, 32'h437f01d4},
  {32'h44b99ede, 32'hc3ab6ac8, 32'hc311a03e},
  {32'hc4ca8d63, 32'hc34af25f, 32'h429e0b53},
  {32'h44e50847, 32'h43d3d629, 32'hc3828cf9},
  {32'hc4816fd4, 32'hc3461cf3, 32'hc30719cb},
  {32'h44dce87c, 32'h4319ad07, 32'h43848c28},
  {32'h433130c0, 32'hc33f3169, 32'h43622bd6},
  {32'h44c464e4, 32'h42258953, 32'hc36d912c},
  {32'hc458eb16, 32'hc3967df9, 32'h4080d965},
  {32'h439f63c6, 32'h43feb4a3, 32'hc328cb67},
  {32'hc487a26e, 32'hc3856fda, 32'h42ef9750},
  {32'h4314c5dc, 32'h439cf5fe, 32'hc30435de},
  {32'hc4ea80ad, 32'h4379c6f5, 32'hc3d1c7fe},
  {32'h446ae723, 32'h437db353, 32'h43154ce8},
  {32'hc2485440, 32'hc031ba8a, 32'h41a97ae6},
  {32'h44d2af8e, 32'h42be25d4, 32'hc31aca46},
  {32'hc5053752, 32'h42ccb3e4, 32'hc293a5fb},
  {32'h448458a6, 32'h4309dd31, 32'hc2ca0148},
  {32'hc4860724, 32'hc38a8614, 32'h4299a016},
  {32'h44f486d1, 32'h4328b5d4, 32'h439bfca0},
  {32'hc492e93d, 32'h437fb01b, 32'hc3dc5642},
  {32'h45083f05, 32'h439f80bd, 32'h42df721d},
  {32'hc4b97108, 32'hc27e4a9a, 32'hc3866993},
  {32'h41307180, 32'h4387808a, 32'hc25f97a0},
  {32'hc3df4ca2, 32'h42128a62, 32'h42c105a9},
  {32'h44df6350, 32'hc337d518, 32'hc26a1b49},
  {32'hc4fde0b3, 32'hc2b4bae2, 32'h43cce05d},
  {32'h44f766aa, 32'h4264bda0, 32'hc3a81fb0},
  {32'hc460227e, 32'hc23a7630, 32'hc27e0bd0},
  {32'h44d40c09, 32'hc3a7d786, 32'hc31b3780},
  {32'hc4eb1caa, 32'h4323d155, 32'h4381f6f4},
  {32'h44386385, 32'hc27adffa, 32'h413f6b6c},
  {32'hc48c30ee, 32'hc15519b3, 32'hc35e7734},
  {32'h43a2a8ec, 32'hc20abf86, 32'h407af55a},
  {32'hc3c4f880, 32'h430a3139, 32'hc365e673},
  {32'h4506ca7b, 32'h3ff6e1d5, 32'h43970582},
  {32'hc44b6638, 32'hc103964f, 32'h428ca33f},
  {32'h44a2556f, 32'hc30118f4, 32'hc013c3cc},
  {32'hc42af4b4, 32'h43560081, 32'hc31aa866},
  {32'h44bbc04e, 32'hc346fee6, 32'hc37d0699},
  {32'hc4852e2a, 32'hc01d4a40, 32'hc388a86b},
  {32'h448b8fa4, 32'hc2aca392, 32'hc3aedf75},
  {32'hc44d6e4e, 32'h43a0ee81, 32'h40ad63a8},
  {32'h44c413fc, 32'h4386c197, 32'h436cff96},
  {32'hc4aa0ef8, 32'hc3a72721, 32'hc3c5523f},
  {32'h45290d6d, 32'h4380c017, 32'h431861f4},
  {32'hc3d7eada, 32'hc38c2401, 32'h438cd05b},
  {32'h45004323, 32'h42729f9a, 32'h4318af72},
  {32'hc4989d6e, 32'hc29e8982, 32'h42b9e264},
  {32'h4506d22d, 32'hc2ec45d8, 32'h4153c6dc},
  {32'hc3c275a1, 32'hc162fe20, 32'h4311f935},
  {32'h44c7df89, 32'h42e64166, 32'h4396cefc},
  {32'hc4f9f7a5, 32'hc3bb6fc5, 32'h4332081c},
  {32'h4518bed4, 32'h4361159e, 32'hc1e6519f},
  {32'hc2f28c76, 32'hc27ea278, 32'hc3b3689b},
  {32'h443a8da7, 32'h43ad9364, 32'h43c7f89f},
  {32'hc45c53d0, 32'hc2db2255, 32'hc2c4e375},
  {32'h44602100, 32'h435ffd08, 32'hc3505f11},
  {32'hc4eb93a8, 32'h427b2426, 32'h42818270},
  {32'hc3306480, 32'hc2b5f851, 32'h43620300},
  {32'hc506df45, 32'h42c42085, 32'hc3444017},
  {32'h44622231, 32'h431f311d, 32'hc2badcac},
  {32'hc4185c3f, 32'h42f17d31, 32'h433ddd24},
  {32'h43e6055c, 32'h4207ccdb, 32'h4383c310},
  {32'hc4557828, 32'hc3729558, 32'h42d5385f},
  {32'h4456d99c, 32'hc3977fc5, 32'h42aca9dd},
  {32'hc436a1b6, 32'h43dd61de, 32'h436f241e},
  {32'hc37f2470, 32'hc30bb101, 32'hc2a6261a},
  {32'h42d18a80, 32'hc358b687, 32'hc3c8e644},
  {32'h4470e46e, 32'hc241e35b, 32'h42f30eb0},
  {32'hc4e041bf, 32'hc36fec2d, 32'hc2de1ead},
  {32'h44fa74d4, 32'h42ad58ff, 32'h43178879},
  {32'hc19a1040, 32'hc1572ebe, 32'hc3250e45},
  {32'h44a015b2, 32'h438b09c4, 32'h43341437},
  {32'hc4fa0de6, 32'h42d46813, 32'hc3a1f1c7},
  {32'h43331928, 32'hc293faf3, 32'h4357efa7},
  {32'hc4823bc8, 32'h43dfb6dd, 32'hc305f2d1},
  {32'h4501dd16, 32'h43c24dd2, 32'h43e3aa1e},
  {32'hc50f0450, 32'hc2984ea2, 32'h427d15a6},
  {32'h43a6efe6, 32'h428fe824, 32'hc3dd57b5},
  {32'hc4bb8841, 32'h4192d76e, 32'h42b8c32e},
  {32'h44fb30b6, 32'h4387a05b, 32'hc178a69d},
  {32'hc4c497fe, 32'h40a83f6c, 32'h43815080},
  {32'h44fabec1, 32'hc2dd3471, 32'h425048d0},
  {32'hc3e892e0, 32'hc36a6d07, 32'hc2658173},
  {32'h44fe0ed8, 32'h412151c8, 32'h43043891},
  {32'hc3977dd7, 32'hc25fac0f, 32'h43b9d172},
  {32'h43b64b8a, 32'hc21e767c, 32'hc2614189},
  {32'hc4c30f56, 32'h42bcff86, 32'hc2b19a80},
  {32'h44dc70a1, 32'h41e08fc7, 32'h42a169c5},
  {32'hc4b38e64, 32'h43dbfeb4, 32'h42bc0a94},
  {32'h428f7dc0, 32'hc3971e74, 32'h431cebfc},
  {32'hc4f170ec, 32'hc3051f36, 32'h40018e84},
  {32'h44a6cd1e, 32'hc2d0c854, 32'h432e30eb},
  {32'h4504fe22, 32'hc3539ba5, 32'hc3e5964f},
  {32'hc50cd92f, 32'hc1ed2129, 32'hc30a57d4},
  {32'h44954f7b, 32'h4316e7a5, 32'hc38925ff},
  {32'hc38256e7, 32'h430947d8, 32'h421e77bd},
  {32'h44a9ad30, 32'h425bce6c, 32'hc2e787cc},
  {32'hc3e51890, 32'hc292aab0, 32'hc2888d98},
  {32'h437d0f5c, 32'h430d0cc3, 32'hc2b0ac20},
  {32'hc5281e35, 32'hc371e86f, 32'hc323ebe7},
  {32'h438889f7, 32'h416ea068, 32'hc3c11197},
  {32'hc4bcef9c, 32'hc33eb23e, 32'hc32bc505},
  {32'h4501e25f, 32'h4197fa48, 32'h4242854c},
  {32'h42d5ad67, 32'h436a9cf0, 32'hc367ffbd},
  {32'h436b1864, 32'hc31ba2d1, 32'hc3ce12a1},
  {32'hc4c3b657, 32'hc2892386, 32'hc2a51d80},
  {32'h44f1df5e, 32'hc2ef9e5f, 32'hc3d3ad54},
  {32'hc504137c, 32'h4352ccf7, 32'hc3439a8e},
  {32'h44237786, 32'h440f2ebd, 32'h428cd46d},
  {32'hc4ed5e7f, 32'h43171dd3, 32'hc3596fad},
  {32'h4416f9ac, 32'hc240a69e, 32'hc3bd8131},
  {32'hc46dcd9c, 32'hc349ed79, 32'hc382b037},
  {32'h44ff03ba, 32'hc30da62d, 32'h426f4c9c},
  {32'hc5026b99, 32'h43262ba9, 32'hc3324e32},
  {32'h4520182f, 32'hc379e6ec, 32'hc3e8d989},
  {32'hbfb97f60, 32'hc416e4fc, 32'h435aff3d},
  {32'h4511dce6, 32'hc2dacf6c, 32'h437e7576},
  {32'h41885a9a, 32'h431f1b07, 32'hc35c8871},
  {32'h45019082, 32'h433daf86, 32'h423010da},
  {32'hc425b263, 32'hc33bbc89, 32'hc21fd5bc},
  {32'h44669e30, 32'h4348db66, 32'h438644e7},
  {32'hc48c3273, 32'h42cea4d0, 32'h4269892d},
  {32'h4437b1c6, 32'hc335ff35, 32'h4308d2b2},
  {32'hc5023794, 32'h43789c12, 32'hc3931fe8},
  {32'h433c5e08, 32'h421e1dd4, 32'h43fc0f7b},
  {32'hc50e01fa, 32'h43a6e32c, 32'h4384b8cf},
  {32'h44d0d5fb, 32'h437257ff, 32'hc33eaa0c},
  {32'hc500a406, 32'h42e6615b, 32'h4315340e},
  {32'hc301d688, 32'hc08348d4, 32'hc12c40ea},
  {32'hc49b71fa, 32'h43e49415, 32'hc307b2cc},
  {32'h4506c594, 32'h426ad6fa, 32'h4339587b},
  {32'hc492d7e3, 32'h433c938e, 32'hc270619d},
  {32'h450e1406, 32'h44192a94, 32'h42d80af3},
  {32'hc43e4b96, 32'hc39aed8e, 32'h42935c7e},
  {32'h440d0aa9, 32'h420fc74c, 32'h41e76d08},
  {32'hc428fd1c, 32'h41f8fa28, 32'h43ccbc25},
  {32'h446169e6, 32'h434248c8, 32'hc44d3193},
  {32'hc511be72, 32'hc2e4218a, 32'hc20475ef},
  {32'h4519d8f6, 32'h4356dd90, 32'hc2f74730},
  {32'hc4e2f23c, 32'hc3434a4a, 32'hc36a3d88},
  {32'h44d2dbfd, 32'h43cdaa0f, 32'hc336bd62},
  {32'hc4a91dc8, 32'hc3421886, 32'h43d37f01},
  {32'h448f3b05, 32'hc39efa67, 32'h4345f1e3},
  {32'hc3b85e58, 32'h420fed18, 32'hc3a0ae0b},
  {32'h441ebf3c, 32'hc2822e10, 32'hc35e6bfb},
  {32'hc5000bac, 32'hc3529f3b, 32'h43126ea4},
  {32'h442081e6, 32'h43f12dbe, 32'h41c86d00},
  {32'hc34ecbb8, 32'hc38d2863, 32'h43538ce9},
  {32'h432ba808, 32'h43dedd2f, 32'hc3838019},
  {32'hc473bbb2, 32'h4339de2c, 32'h43c214b9},
  {32'h44fc6484, 32'hc210fc4a, 32'h4370862e},
  {32'hc4ac2923, 32'h3f3d4970, 32'hc3ee063b},
  {32'h44aad066, 32'hc398c219, 32'hc410eb87},
  {32'hc4880539, 32'h42a506f3, 32'h42014058},
  {32'h44887e49, 32'hc1afb259, 32'hc3ca10c3},
  {32'hc41773cc, 32'h4254a320, 32'hc3870313},
  {32'h445c2392, 32'hc2390ebe, 32'hc3bfced1},
  {32'hc4a355a7, 32'h439daf4e, 32'hc2c908e4},
  {32'h4501ee94, 32'h42b62190, 32'h4298d4ab},
  {32'hc4f183c0, 32'h411903b8, 32'h43a7ee78},
  {32'h45039fb0, 32'hc3da72fa, 32'hc2486d0b},
  {32'hc4a464fe, 32'h435532a5, 32'h41849aa5},
  {32'h44796f82, 32'h422dd38a, 32'h419212d1},
  {32'hc2a299b0, 32'hc24d2ee5, 32'hc1e36eb8},
  {32'h44de64fc, 32'hc34d6610, 32'hc3809793},
  {32'hc46390e0, 32'hc2963b24, 32'h43554a92},
  {32'h44706685, 32'h4207a82a, 32'hc1271ba8},
  {32'hc47c92c4, 32'h4300cdc2, 32'h4427432e},
  {32'h43c36700, 32'h42d83100, 32'h41b08419},
  {32'h41979d0e, 32'hc324d5de, 32'h43d7c765},
  {32'h44f83cee, 32'h428c3540, 32'h43828201},
  {32'hc4099924, 32'hc34ec67a, 32'h426da1c4},
  {32'h445891dc, 32'hc11d69a3, 32'hc34fb1f7},
  {32'hc4b786da, 32'hc235250b, 32'h4396296b},
  {32'h4416646c, 32'hc3490e7c, 32'hc3f256ab},
  {32'h4309bd4a, 32'h42990ae6, 32'h43cb49f8},
  {32'h449a461e, 32'h43820afd, 32'h42798b9a},
  {32'hc4f06dc2, 32'h42f214bc, 32'h4228e2f2},
  {32'h44aae0d8, 32'h4317e215, 32'hc1aa9211},
  {32'hc3267920, 32'h43504b8c, 32'h4300d904},
  {32'h44e8f175, 32'hc2024321, 32'hc2dfef94},
  {32'hc5038713, 32'h431b1aaa, 32'hc3891ee7},
  {32'h451de5b7, 32'hc38bf022, 32'hc3884b1a},
  {32'h4439c947, 32'hc239df48, 32'hc33577b5},
  {32'hc428f6a0, 32'hc287ea7b, 32'h420fc59d},
  {32'h45004405, 32'hc3110b24, 32'h4385d4d6},
  {32'hc4d16f4c, 32'h42bd5c10, 32'h4288bb79},
  {32'h44424e36, 32'h433d3bb5, 32'hc2ec03aa},
  {32'hc387d3d0, 32'h43b62044, 32'h430510e6},
  {32'h43c0bdc8, 32'hc3bc3f8a, 32'hc4190ac5},
  {32'hc4c8ab61, 32'hc2c96b4a, 32'hc29578d2},
  {32'h4497d719, 32'h4318fae6, 32'hc3108631},
  {32'hc441d304, 32'h4300cfcc, 32'h43020d40},
  {32'h438f3dd4, 32'h4302a801, 32'h41b7caa4},
  {32'hc486c1b9, 32'h42a673d8, 32'h4392b849},
  {32'h4426306d, 32'h43130ea3, 32'hc2d4426b},
  {32'hc4862110, 32'hc23f6d2a, 32'hc1fbcd01},
  {32'h44bab702, 32'hc290bde1, 32'h425c13d7},
  {32'hc4b8966f, 32'h420fdefc, 32'h431f1335},
  {32'h443d4de4, 32'h43ed54a5, 32'hc316e88f},
  {32'hc44196a0, 32'h43371a9a, 32'h430f714d},
  {32'h43400301, 32'h43e0ccbb, 32'h4260c431},
  {32'hc422001e, 32'h431ec8a8, 32'hc21f8e02},
  {32'h444af6e6, 32'hc3d1377e, 32'hc35e49ff},
  {32'hc4318ca8, 32'h4280a200, 32'hc29d5cdb},
  {32'h4458f913, 32'hc1e58849, 32'hc310c990},
  {32'hc4f1c3b5, 32'h4203bb86, 32'h435a3209},
  {32'h441d84ba, 32'hc339cc61, 32'hc33fb657},
  {32'hc4e8db80, 32'hc2f44437, 32'h43199520},
  {32'h44069c3c, 32'hc2185585, 32'hc3a21c03},
  {32'hc4f968c5, 32'hc382b31b, 32'hc3009deb},
  {32'h450e928d, 32'hc2fa9cc4, 32'hc27fb6fb},
  {32'hc4a62888, 32'hc3650eaa, 32'hc3b1ab6c},
  {32'h43ccae10, 32'hc341a4b9, 32'hc3333279},
  {32'hc3762934, 32'hc2333d55, 32'hc237dc72},
  {32'h447d4608, 32'h432e8eba, 32'hc2426892},
  {32'hc4ebef6b, 32'hc34129d4, 32'h42a2adb7},
  {32'h44e172d7, 32'h4256fa03, 32'hc2de85db},
  {32'hc495c0fe, 32'hc35241f8, 32'hc304c6c9},
  {32'h44c35f0d, 32'h418ad0e6, 32'h41a2fdcd},
  {32'hc4a38006, 32'h435bd11e, 32'hc2701ed5},
  {32'h440d7a67, 32'hc3840a7b, 32'h3f6e90b2},
  {32'h43515a50, 32'hc108cc5d, 32'hc304f3c4},
  {32'h45159bb6, 32'h42ce346e, 32'hc18f4ef2},
  {32'hc4662bfc, 32'h43aadcc6, 32'h41fae639},
  {32'h43ce42dc, 32'h4205cffa, 32'hc1af105b},
  {32'hc4fc9049, 32'hc279fa33, 32'h42fafa95},
  {32'h44e6f59d, 32'h41fb2dd0, 32'h42840c42},
  {32'hc4ad88f0, 32'h4401ca82, 32'h4138ac43},
  {32'h450f3365, 32'h4360bc99, 32'hc3102855},
  {32'hc4205648, 32'h42a2692b, 32'hc36e8940},
  {32'h436a9700, 32'hc273d484, 32'h433607f0},
  {32'hc4dc25a4, 32'h42c5fb60, 32'hc22be2eb},
  {32'h4531c310, 32'hc1d8a71f, 32'h419c5064},
  {32'hc486698a, 32'hc30ae46c, 32'hc31eeaee},
  {32'h449d7eec, 32'h431abc7b, 32'h41861580},
  {32'hc508be91, 32'hc2c36c2d, 32'hc2781e12},
  {32'h439e1aa1, 32'hc2cfaef4, 32'hc3ccaec7},
  {32'hc50e694a, 32'hc20588af, 32'hc35720da},
  {32'h4476dcfc, 32'hc39d0f04, 32'hc27502f3},
  {32'hc3201520, 32'h42bb7dac, 32'hc2ff18cc},
  {32'h447e6e66, 32'h43ac2296, 32'h440050ae},
  {32'hc49b352e, 32'hc3961675, 32'h43367275},
  {32'h44ad960e, 32'hc3c4d484, 32'h4323848c},
  {32'hc43e7085, 32'hc30595de, 32'h433fba8c},
  {32'h43dfde96, 32'hc33d57c8, 32'h426fff59},
  {32'hc508ea46, 32'hc03066a8, 32'h43396a05},
  {32'h44f34a9a, 32'hc391217c, 32'hc1968884},
  {32'hc4c53622, 32'hc3834e15, 32'h424f4714},
  {32'h451bccef, 32'hc3f686ed, 32'h436eb657},
  {32'hc42c738e, 32'hc40862cd, 32'h437ee2e1},
  {32'h44f7a532, 32'h43859579, 32'hc34b30d2},
  {32'hc45c04c3, 32'hc27ce3a7, 32'h42f73496},
  {32'h44e465ec, 32'hc2a66902, 32'hc0605514},
  {32'hc4c6369c, 32'h416dd522, 32'h4331bdd7},
  {32'h4455a0b6, 32'h4232b78c, 32'hc316b991},
  {32'hc43f08ce, 32'h4252807f, 32'h4249f024},
  {32'h4480f187, 32'hc287dbf1, 32'hc306b496},
  {32'hc38eb5c8, 32'hc2ad0ee9, 32'hc3a4a9b7},
  {32'h44e2e118, 32'hc36b5055, 32'h420ccd12},
  {32'hc44fab63, 32'h43d31ce8, 32'h4312b6ad},
  {32'h450eadf3, 32'hc202c4f2, 32'h44279f3e},
  {32'hc51e61cb, 32'hc367c22e, 32'hc2eb87d7},
  {32'h44e54d5e, 32'h431491fd, 32'h42a28451},
  {32'hc503db8d, 32'h43582df6, 32'hc330c997},
  {32'h43e1b5cc, 32'h42a6b30e, 32'h41cdd40c},
  {32'hc4ff902a, 32'h42ab365e, 32'h435822db},
  {32'h4506837c, 32'hc3c1b2f3, 32'h4422bfe7},
  {32'hc41635ea, 32'hc366be89, 32'hc29b5628},
  {32'h42e21490, 32'h43f8ff6a, 32'h42d025a7},
  {32'h42812820, 32'h42d42eae, 32'hc38a53a2},
  {32'h444d897c, 32'hc33b4e3b, 32'hc02d3040},
  {32'hc43ec610, 32'h42679be0, 32'hc3b9cfba},
  {32'h44c3579a, 32'hc22091ae, 32'h4316af5f},
  {32'hc4cd4728, 32'h43ab5757, 32'hc2af4d68},
  {32'h427d5ec0, 32'hc367bb12, 32'h4297f7b5},
  {32'hc2caa8ed, 32'hc289d611, 32'hc317455b},
  {32'h44f43391, 32'h431760ee, 32'h4395aa17},
  {32'hc4d67bbd, 32'h435083e2, 32'hc30d5b4c},
  {32'h4378ed4c, 32'h42c12bde, 32'h424ce305},
  {32'hc45abbc4, 32'hc30cfcc9, 32'hc206de1e},
  {32'h450bbf35, 32'hc2b53040, 32'hc369ec98},
  {32'hc4dbebd7, 32'hc3674f8f, 32'h43ec2085},
  {32'h44dc9054, 32'h43b1f981, 32'h433ca37e},
  {32'hc4dd9549, 32'h3fe9e71f, 32'hc24d956c},
  {32'h44ea1aac, 32'h42bca671, 32'h4354c7b4},
  {32'hc487e566, 32'h431ca140, 32'h43b33e4d},
  {32'h43d96c14, 32'h418f7968, 32'h435040b4},
  {32'hc4e95e78, 32'h42b93435, 32'hc379c29e},
  {32'h44acda56, 32'hc2cc4dae, 32'h43417f63},
  {32'hc3324960, 32'h43986fda, 32'h4315bbb2},
  {32'h4468f2b8, 32'hc2d5f488, 32'h42402b98},
  {32'hc4ec454c, 32'hc2bc7b8a, 32'h4368deca},
  {32'h44d1cccd, 32'hc24f30c3, 32'h42a16454},
  {32'hc45f9892, 32'hc36ebea0, 32'hc2c38770},
  {32'h44f4ca0b, 32'h42d68c35, 32'hc328258d},
  {32'hc48fa75c, 32'hc1b85ab8, 32'h43d0dd55},
  {32'h43d64f92, 32'hc35957bd, 32'h4309f453},
  {32'hc3f359d0, 32'hc3df5dcc, 32'hc22fea2a},
  {32'h43e144a8, 32'hc296372a, 32'h43e0e248},
  {32'hc44e4138, 32'h41f8d417, 32'hc2edcc54},
  {32'h446f8a4e, 32'h434e45af, 32'hc38c2fc2},
  {32'hc5106073, 32'h42dbac8e, 32'hc36b60db},
  {32'h4466fa9c, 32'h429adacf, 32'hc31ccc27},
  {32'hc4f016f8, 32'h43d87cb6, 32'h40cb7fc4},
  {32'h451257ed, 32'hc3e7d7a6, 32'hc1bfcbd8},
  {32'hc4866169, 32'h400417f5, 32'hc3020b07},
  {32'h44a81f54, 32'hc32a7f38, 32'h432620f5},
  {32'hc1eb5268, 32'h4341a2c2, 32'h43484e7f},
  {32'h43341338, 32'h426f45e8, 32'h42f32eee},
  {32'hc4a0479e, 32'hc2f26e0c, 32'hc1e809d3},
  {32'h4513634c, 32'h439f9236, 32'h404c7310},
  {32'hc492f6c5, 32'hc1a83790, 32'h42bfd656},
  {32'h440ffd6c, 32'h42144890, 32'hc37648b6},
  {32'hc4b2efa8, 32'hc38838cd, 32'hc2ad6e88},
  {32'h44bd7738, 32'h437cafc7, 32'h4310602f},
  {32'h4367f080, 32'hc3f13a9e, 32'hc1a0f470},
  {32'h44c0223a, 32'h42aa353e, 32'h438fd642},
  {32'h4288b89f, 32'hc228eeca, 32'hc20811ab},
  {32'h44b5157b, 32'h43eddaf7, 32'hc21d4aeb},
  {32'hc4fb9522, 32'hc3b5abc8, 32'hc2e944a6},
  {32'h4442bed8, 32'h42dbfbd7, 32'h42faa31e},
  {32'hc36c54ee, 32'h4327800e, 32'h40410c44},
  {32'h44549ec4, 32'hc2c83cac, 32'hc1c0a854},
  {32'hc41c1e6c, 32'h43cfd77a, 32'h4323eea2},
  {32'h432dfa24, 32'hc3d6d169, 32'hc252367e},
  {32'hc4f5a8fd, 32'h42a4ba9d, 32'h43448edd},
  {32'h4494953f, 32'h3f997709, 32'h43343549},
  {32'h432aec70, 32'h4363183a, 32'hc2412371},
  {32'h444c8fd1, 32'hc30d324e, 32'hc151bd40},
  {32'h436c55e8, 32'h4381d137, 32'hc31f1c2e},
  {32'h45067308, 32'hc3aa927d, 32'h43f599a0},
  {32'hc414ea14, 32'h4117d25e, 32'hc1107b47},
  {32'h44c87c0e, 32'hc3459fb8, 32'h42ae8dc2},
  {32'hc4ea924b, 32'h40c56040, 32'hc2c10a64},
  {32'h44227882, 32'hc37fb4a7, 32'hc2702af5},
  {32'hc4f46cd0, 32'hc3ecf835, 32'hc2770c2b},
  {32'h4487bac4, 32'h430f7061, 32'hc39c5708},
  {32'hc501c490, 32'hc2a92e64, 32'h42b15db2},
  {32'h4508bd04, 32'h4350e869, 32'h4296e65e},
  {32'hc4110bee, 32'hc0bddf41, 32'hc3382cc7},
  {32'h44f150a2, 32'h42a39c36, 32'hc2f425f0},
  {32'hc43dfeb6, 32'h4361b8f0, 32'hc18225e5},
  {32'h44414daf, 32'hc273a725, 32'hc3d90675},
  {32'hc4e87225, 32'hc28d7356, 32'hc20e2363},
  {32'h42f00158, 32'hc32d4d20, 32'h42a8129a},
  {32'hc4363320, 32'hc3bad460, 32'hc28e4f8b},
  {32'h4503d75d, 32'hc28d7e45, 32'h4325637d},
  {32'hc43fcdb8, 32'h43a0f38e, 32'hc14d9c20},
  {32'h43fc14f2, 32'h4375f756, 32'hc3faec8b},
  {32'hc5183681, 32'hc230cc38, 32'hc36ba710},
  {32'h45075c86, 32'hc2900e12, 32'h432e7950},
  {32'hc3dc84fe, 32'hc3696f34, 32'h42e66219},
  {32'h44d2bd29, 32'hc2cb4e0e, 32'hc3760c59},
  {32'hc4a51a3c, 32'h4418bd30, 32'h434a708f},
  {32'h44bc2d26, 32'hc2b64160, 32'h41c03e11},
  {32'hc3a10236, 32'hc2868be5, 32'hc252c3df},
  {32'h43e4e76d, 32'h43847a8b, 32'h43ec4550},
  {32'hc50945ba, 32'h42bfeca4, 32'h4320ef09},
  {32'h44b8ec8e, 32'hc1e5e22f, 32'hc20dd79b},
  {32'hc4baec9a, 32'hc30d4d4d, 32'h42c1adf5},
  {32'h44f209cb, 32'h420642ec, 32'h426604c2},
  {32'hc4921516, 32'h416386f5, 32'h4108144c},
  {32'h44fa26fe, 32'hc2d8303a, 32'h42bed4fa},
  {32'hc4532df1, 32'hc25b9a0d, 32'hc31492c6},
  {32'h43d8b840, 32'h42ee19f0, 32'h4375180e},
  {32'hc4e57c52, 32'hc3525937, 32'hc3a88132},
  {32'h4492d592, 32'hc3a7400e, 32'h41d8fedb},
  {32'hc4b8d704, 32'hc345630f, 32'h434138f1},
  {32'h4428f294, 32'hc2e7df33, 32'hc345211b},
  {32'hc50698fb, 32'h4307f113, 32'hc20efc86},
  {32'h445d9b04, 32'h42874078, 32'hc2c8d235},
  {32'hc5140754, 32'hc38ad938, 32'hc186c5f4},
  {32'hc2679ac0, 32'h43789a7f, 32'hc3517874},
  {32'hc487ad8f, 32'hc384c3b4, 32'h41c75c98},
  {32'h44882f4a, 32'h43806a52, 32'hc1486fb8},
  {32'hc50d7a6a, 32'hc3e1634d, 32'hc1e9272a},
  {32'h44ffe642, 32'h412ce059, 32'h43c07577},
  {32'hc48fb287, 32'h4374e421, 32'h40f761be},
  {32'h443813b8, 32'h431a7714, 32'hc35595be},
  {32'hc4f275e9, 32'hc37469a8, 32'h435221f0},
  {32'h4488c772, 32'h41a50ce3, 32'hc2c58970},
  {32'hc388f640, 32'h431aa3bb, 32'h43a9a667},
  {32'h44b15fce, 32'h432b3915, 32'h42d0617e},
  {32'hc50ffdc9, 32'hc30deaaa, 32'h4333749e},
  {32'h44cd1b7e, 32'h43278490, 32'h42bb960f},
  {32'hc3b14d2e, 32'h41b343f2, 32'hc271b550},
  {32'h43fce360, 32'h434e9f08, 32'hc31d2005},
  {32'hc3f0cd12, 32'h41daf252, 32'hc3a35d7e},
  {32'h449c2708, 32'hc3e6d475, 32'h4261bd68},
  {32'hc4d10c44, 32'h4312b1ab, 32'hc379e530},
  {32'hc0715f00, 32'hc3b018fb, 32'hc2813672},
  {32'hc3c0d896, 32'h434670d7, 32'hbfa183a0},
  {32'h44313fd9, 32'hc2fb9a2c, 32'h4359c937},
  {32'hc4eb31de, 32'hc32f08c6, 32'h43ee6501},
  {32'h4519ec63, 32'h43eec7b4, 32'h4376f7f0},
  {32'hc440dfd4, 32'hc3215df5, 32'hc2cacc73},
  {32'h442b7ad2, 32'hc276b938, 32'h43005284},
  {32'hc4a1cb1c, 32'hc106f422, 32'h42d8239d},
  {32'h439767d6, 32'hc373ae35, 32'hc34c417f},
  {32'hc486f6bb, 32'hc1f455be, 32'hbf833040},
  {32'h44a084b3, 32'hc3110073, 32'hc39e872f},
  {32'hc3891b98, 32'hc10eedda, 32'h43aec788},
  {32'h44fecfdc, 32'hc1a771db, 32'hc303edb4},
  {32'hc46b1b84, 32'h4425783a, 32'h43267001},
  {32'hc29af110, 32'hc29be4b7, 32'h428e7b95},
  {32'hc414255e, 32'hc223d9e3, 32'hc35f7ad1},
  {32'h4445f464, 32'hc34ee043, 32'hc384c881},
  {32'hc51d7d70, 32'h41037ff0, 32'h4235785d},
  {32'hc38b0d44, 32'h43f427a2, 32'h438a66ae},
  {32'hc49085e2, 32'h42d86cdc, 32'hc3073c7c},
  {32'h447effd4, 32'hc20ddc95, 32'hc38f3798},
  {32'hc4f4ed8b, 32'hc2d0c0dc, 32'h431ae0b0},
  {32'h44a9e373, 32'h4320e309, 32'hc305590d},
  {32'hc458a64c, 32'h42906dd7, 32'h41143c31},
  {32'h451f7f92, 32'hc3a558c9, 32'hc28d62d7},
  {32'hc4faf43c, 32'hc19bdf09, 32'h437c59a3},
  {32'h44606dcc, 32'h42320910, 32'hc2e7b218},
  {32'hc4e8a3b0, 32'hc38188e7, 32'hc3cab609},
  {32'h42c8af00, 32'h438b9d54, 32'hc359ec43},
  {32'hc482105f, 32'hc28f31dc, 32'hc347cad5},
  {32'h44f21ef7, 32'h43b69c4e, 32'h435271e5},
  {32'hc5022483, 32'hc1309df7, 32'hc34af45b},
  {32'h444d77e8, 32'hc38dcd0d, 32'hc379f063},
  {32'hc4f86bc8, 32'h42e1ea38, 32'h423e568e},
  {32'h44b75394, 32'hc33926c1, 32'hc231d2bc},
  {32'hc4f0a447, 32'h42e4074b, 32'h42dbd2cc},
  {32'h438a44bd, 32'h42183a4e, 32'h4256c992},
  {32'hc45776e4, 32'h42c56895, 32'hc298cb00},
  {32'h43ef8df4, 32'hc3dc8be6, 32'h42a2c60e},
  {32'hc3b75e90, 32'h40b66ae9, 32'hc3f6c427},
  {32'h44bb0ad5, 32'h42b9645e, 32'hc3578418},
  {32'hc4572c77, 32'h42743268, 32'h43509da1},
  {32'h4491def7, 32'h43059259, 32'h42df9c6b},
  {32'hc4dc5857, 32'h426fe825, 32'h43217b6c},
  {32'h436bbafc, 32'hc3e3160c, 32'hc310ac8e},
  {32'hc4afc862, 32'hc098075c, 32'hc2a60cc2},
  {32'h43e6f548, 32'hc32cf8b9, 32'hc371889d},
  {32'hc3e344c0, 32'h43210bae, 32'h4339cc4c},
  {32'h43dcaec1, 32'hc39cd931, 32'hc296281e},
  {32'hc416f2b9, 32'h41f36be6, 32'h426bde8d},
  {32'h452a7e05, 32'hc24aefd1, 32'hc387337a},
  {32'h4368fa08, 32'h42832796, 32'h43e54650},
  {32'h4442fe16, 32'hc0d4baec, 32'hc3825344},
  {32'hc4dc0809, 32'h43b8848e, 32'hc20dd901},
  {32'h43d8d84b, 32'hc290eed7, 32'h40ea5cf9},
  {32'hc50caee8, 32'h437dcbc3, 32'hc3032e88},
  {32'h45254db0, 32'h428f21a2, 32'h42c3ac78},
  {32'hc46b3e68, 32'hc25e1c78, 32'hc301f21f},
  {32'h44e8eeec, 32'h43085ed9, 32'h415ad8ba},
  {32'hc492579c, 32'hc334dabd, 32'h4027b130},
  {32'h44fd9f26, 32'h42f9792a, 32'hc22df0a5},
  {32'hc489f5d6, 32'hc2da736d, 32'hc24b3fa3},
  {32'h44d41226, 32'h42aa922d, 32'h4231f6e0},
  {32'hc4291796, 32'h437252fe, 32'h4307052a},
  {32'h44a2e015, 32'h42aac434, 32'hc34b174d},
  {32'hc49a67ea, 32'hc2ada3cc, 32'hc1b6554c},
  {32'h442305b4, 32'hc01ff259, 32'hc3c9f612},
  {32'hc4dfa5da, 32'h42fa8b38, 32'hc3331194},
  {32'h44915ca8, 32'hc3277372, 32'hc2a3ea3a},
  {32'hc4d06d1b, 32'h42f34c1d, 32'h429e223d},
  {32'h4405b95c, 32'h43c84ba7, 32'hc255c873},
  {32'hc5070c7d, 32'h42fd4bac, 32'hc386dd05},
  {32'h42d705b0, 32'h43c13077, 32'h43880cd8},
  {32'hc39ced78, 32'h42cc3125, 32'hc0e5f24e},
  {32'h44ec7784, 32'h434d8560, 32'hc3185e37},
  {32'hc4ee157a, 32'hc4156e0b, 32'hc33a32b9},
  {32'h450e41a0, 32'hc2bf01d8, 32'h41e6d4a3},
  {32'h42dbaa62, 32'h42e09589, 32'hc24f4af5},
  {32'h45032fc4, 32'h436de764, 32'h4355ebe5},
  {32'hc4ca1bab, 32'hc38ac6b4, 32'h43048548},
  {32'h44e0794f, 32'hc1f5da13, 32'hc314c5ba},
  {32'hc2bc1ae0, 32'h420d0dc7, 32'h43085d8e},
  {32'h44114f21, 32'h432e15bc, 32'hc390d1ae},
  {32'hc4066546, 32'h438e5a88, 32'hc3dfc5ef},
  {32'h44c8c939, 32'h43305cf1, 32'hc1d557a6},
  {32'hc307c0c0, 32'hc303bf66, 32'h4363cc5c},
  {32'h432a5e90, 32'hc3891756, 32'hc2560d0f},
  {32'hc4e489c7, 32'h40c8f22a, 32'h4363db7c},
  {32'h4405014e, 32'h43b4060e, 32'h43305bea},
  {32'hc443c20c, 32'h43328862, 32'h43713cd2},
  {32'h441a94f6, 32'h421c1f5e, 32'h42a9707c},
  {32'hc4b0b9c6, 32'h431a255d, 32'h43895ceb},
  {32'h45007969, 32'hc374cd06, 32'hc3d43876},
  {32'hc4afa26e, 32'h41e9b96c, 32'h418e3360},
  {32'h44f1651e, 32'h42aa32a6, 32'h413317a4},
  {32'hc484a3ad, 32'hc28c3209, 32'h426a4722},
  {32'h44f29ecd, 32'h42c5cea6, 32'hc18ed453},
  {32'hc47da26f, 32'h40c1e102, 32'h43269594},
  {32'h45158d11, 32'hc30a9d3f, 32'hc2dc335d},
  {32'h429896ee, 32'h41ca62ca, 32'hc26f93db},
  {32'h44ce3b9a, 32'hc2acda2e, 32'h43fdd084},
  {32'hc52335e1, 32'h43e5234c, 32'h40c50d14},
  {32'h450d211a, 32'h4356146a, 32'hc220ea63},
  {32'hc41cd000, 32'h439097df, 32'h430b268c},
  {32'h450ec924, 32'hc28f45d9, 32'hc3178159},
  {32'hc4c09e28, 32'hc3ba180a, 32'h4061369a},
  {32'h44d7061a, 32'hc1da1306, 32'h42966fae},
  {32'hc4ca27d7, 32'h42d38245, 32'hc30ccf12},
  {32'h4496340d, 32'h4363b4df, 32'hc33aa536},
  {32'hc46e84ba, 32'hc34f46da, 32'h439985b2},
  {32'h4502bd8b, 32'hc176f774, 32'hc41888b1},
  {32'hc404d137, 32'hc30cafa5, 32'hc214c33e},
  {32'h4457c2e0, 32'h41af3dee, 32'h425364df},
  {32'hc50eb80d, 32'h43bcbd90, 32'h42ff3508},
  {32'h4485aeb9, 32'hc2797561, 32'h4317f4ad},
  {32'h40ad1b48, 32'h440bce1d, 32'h43c08249},
  {32'h440ee660, 32'hc3359a44, 32'hc39312d6},
  {32'hc3cb6ae7, 32'h436aa2eb, 32'h430ee8ff},
  {32'h444db06a, 32'hc3c1d1d3, 32'h413a316c},
  {32'hc509df79, 32'h41a0aa5a, 32'h4328dccf},
  {32'hc231a168, 32'hc25cc79c, 32'hc3a579f3},
  {32'hc4d88434, 32'h43e83d04, 32'h424ec06a},
  {32'h4441710e, 32'h42061360, 32'hc35cff17},
  {32'hc3ce5174, 32'hc1155c77, 32'h42875997},
  {32'h450b2f06, 32'hc36c4a5d, 32'h425d1a99},
  {32'hc4aa9fd9, 32'h42aa7df0, 32'h42a344e0},
  {32'hc28df854, 32'h4260ede4, 32'h43242104},
  {32'hc30ac697, 32'hc3b5efb8, 32'h43a434e2},
  {32'h44a28059, 32'hc338b3d7, 32'h41ffa9f5},
  {32'hc4d25f78, 32'hc39838f7, 32'hc2ee7178},
  {32'h4519a404, 32'h434f8670, 32'h434b3f3c},
  {32'h431d7dc0, 32'hc3d5097e, 32'h438fca46},
  {32'h44b88f71, 32'hc34358e7, 32'hc12f8c70},
  {32'hc47a630e, 32'hc3362484, 32'hc1df228b},
  {32'h4510050d, 32'hc292b252, 32'h430545b6},
  {32'hc50d1e8a, 32'h432c0c49, 32'hc3045219},
  {32'h44b1435d, 32'hc2b0f55a, 32'hc333197d},
  {32'hc4c7c2e0, 32'h438a86b0, 32'h43aa3702},
  {32'h45039306, 32'hc38c8128, 32'h42067cb9},
  {32'hc4a72609, 32'hc2d1b2f2, 32'h43240088},
  {32'h4518c776, 32'hc2c92ac0, 32'hc3d640a0},
  {32'hc4c6f224, 32'h431842bf, 32'hc22e1618},
  {32'h451f35af, 32'hc26b97c1, 32'hc23960be},
  {32'hc485ee16, 32'hc2294a49, 32'hc2edad82},
  {32'h44cb196f, 32'h43a3cdad, 32'h4002680f},
  {32'h413e8600, 32'hc29eaa72, 32'h42db1d52},
  {32'h44ef66c4, 32'h428967d3, 32'h42561ae0},
  {32'hc4de51da, 32'hc2fe01e7, 32'h41d1a294},
  {32'h44e3e94e, 32'h43111fad, 32'h43c25efa},
  {32'hc4606c78, 32'h42c904e9, 32'h42fd0fc0},
  {32'h4478d5dd, 32'hc26dd828, 32'hc3494aba},
  {32'hc4a838e2, 32'hc1fb168a, 32'h4355a541},
  {32'h4330afac, 32'hc32dd1c1, 32'hc394c540},
  {32'hc2bce062, 32'h43346747, 32'hc3090f67},
  {32'hc3965152, 32'hc33f4dec, 32'hc35a8e7c},
  {32'hc4e41328, 32'h4324a030, 32'h435a0000},
  {32'h4458a5b6, 32'hc3a4de8e, 32'h432917c0},
  {32'hc50bab74, 32'h4367ecbe, 32'hc35b82fa},
  {32'h44b7afb9, 32'h428acc5d, 32'hc3448c35},
  {32'hc4d9b415, 32'h432d60b9, 32'hc3458aa0},
  {32'h44db0888, 32'h41aa73ea, 32'hc3949321},
  {32'hc3ac1a1c, 32'h43b7fa87, 32'hc374ffb7},
  {32'h4519c8ed, 32'h44007229, 32'hc3802e69},
  {32'hc509ab1f, 32'hc188375c, 32'h437f09b6},
  {32'h44b16f03, 32'hc194d993, 32'h439b1195},
  {32'hc4303e1c, 32'hc36a1822, 32'h42420f5a},
  {32'h44a7ddfe, 32'h437e930e, 32'h4305fc6c},
  {32'hc4ca3a35, 32'h432b6e39, 32'h42fbc236},
  {32'h446974bd, 32'hc3671d07, 32'h43f0fc2c},
  {32'hc1fd9d93, 32'h433b6512, 32'hc2339cb9},
  {32'h44278442, 32'h436a7038, 32'hc3bb9c3b},
  {32'hc3eb1067, 32'h43966145, 32'h43869e32},
  {32'h448fd8d9, 32'hc257a1ee, 32'h432ddb1c},
  {32'h434d3ea0, 32'h433c314e, 32'h43efd984},
  {32'h44ccb6d8, 32'hc2f348dd, 32'hc301feea},
  {32'hc4d6f10d, 32'h41ef0e39, 32'hc365271f},
  {32'h444c9529, 32'hc31cb60e, 32'h4391918a},
  {32'hc4fbd8d9, 32'hc362d6d8, 32'h41b26ad4},
  {32'h44b492d7, 32'h432964ac, 32'hc3209025},
  {32'hc3afae9a, 32'hc2f7a7d1, 32'hc3625c26},
  {32'h442bb0d5, 32'hc37df9e6, 32'hc2cb18c0},
  {32'hc5182e73, 32'h4300389e, 32'hc2be1a1b},
  {32'h44f310a1, 32'h43148d5a, 32'hc2e9e511},
  {32'hc50c8f51, 32'h43625539, 32'h43ce6e2f},
  {32'h448b0470, 32'h42695725, 32'h4380c0da},
  {32'hc4d71018, 32'hc1f711e9, 32'hc3fa20e2},
  {32'h44ee5a0a, 32'hc3aacde8, 32'h42c0b1e7},
  {32'hc4f0affb, 32'h435e9aad, 32'hc3967241},
  {32'h441559cc, 32'h4216c4fc, 32'h4381f721},
  {32'hc495a372, 32'h43aa512f, 32'hc1374029},
  {32'h44960752, 32'hc369b35d, 32'h41231aca},
  {32'hc48f9fa5, 32'hc30c8971, 32'hc39fee8c},
  {32'h43683778, 32'h412d49fe, 32'h43cd2521},
  {32'hc3423bf0, 32'h4310380a, 32'hc2fcc020},
  {32'h4513cca2, 32'h4322b48c, 32'hc32e1b4b},
  {32'hc497239d, 32'hc179df8c, 32'hc2dbd1c5},
  {32'h44588569, 32'h43432db7, 32'hc2bb4b27},
  {32'hc40f618a, 32'h43d790c5, 32'hc1e70c07},
  {32'h442800bc, 32'h4380cdfc, 32'h435bc92d},
  {32'hc414aa91, 32'h42903496, 32'hc30a7c20},
  {32'h440c460f, 32'h43301bb5, 32'h43449474},
  {32'hc4c8f64b, 32'h42fe5c57, 32'hc316083e},
  {32'h44b2718f, 32'h422ee055, 32'hc3842123},
  {32'hc489137c, 32'hc2383e71, 32'h437493f3},
  {32'h44cbdcff, 32'hc3ac43aa, 32'hc31ceb51},
  {32'hc485b058, 32'h420108c7, 32'h42bfe3cb},
  {32'h44e5db04, 32'h42ac1d16, 32'h4343b462},
  {32'hc4c1070f, 32'h43ceaacb, 32'hc31a38c8},
  {32'h44b08f2b, 32'hc221df4b, 32'h43a7bc47},
  {32'hc38a2020, 32'h42f48cbb, 32'h42ae228a},
  {32'h441feb37, 32'h40b1cb86, 32'hc34c78d8},
  {32'hc43c4ece, 32'h43614748, 32'hc394725d},
  {32'h440ddcde, 32'hc2db127c, 32'h43a39b28},
  {32'hc4814788, 32'h42bbb337, 32'hc3af8604},
  {32'h43baeadc, 32'h42762ad6, 32'h43216d2d},
  {32'hc4ca1fb8, 32'hc290190a, 32'hc136551a},
  {32'h4430e84c, 32'h413272eb, 32'h43361e21},
  {32'hc4a08016, 32'h43302d43, 32'h427e4e45},
  {32'h44ca4029, 32'hc3347db8, 32'h438786a9},
  {32'hc472acd0, 32'hc24a15c8, 32'h42ad1548},
  {32'h44867016, 32'hc2c95a58, 32'h4288e5f5},
  {32'hc4ced93c, 32'h42a7a96c, 32'h411134ec},
  {32'h4414127e, 32'h42cdd688, 32'h4380f6ca},
  {32'hc42a1d3a, 32'h43db76f9, 32'h42fadd36},
  {32'hc4836e3e, 32'hc3748809, 32'hc303477b},
  {32'h44fecb34, 32'hc1851f5e, 32'h4211ceb8},
  {32'hc3f3bf40, 32'h43d84d7f, 32'hc3843f31},
  {32'h4499c84e, 32'h4324b112, 32'h432056af},
  {32'hc5060309, 32'h42834bd5, 32'hc33d395a},
  {32'h44e0d948, 32'hc2f7d03f, 32'h43c3558f},
  {32'hc45ead9c, 32'hc3c293d6, 32'hc311bc2d},
  {32'h44e118f2, 32'hc3b7a358, 32'hc2921971},
  {32'hc40c1608, 32'h43474a2a, 32'hc32d297c},
  {32'h44c70331, 32'hc308f13d, 32'h41a4fd57},
  {32'hc36f5270, 32'hc1c1b510, 32'hc2a3dfa8},
  {32'h44be89a0, 32'hc321a754, 32'h4381d294},
  {32'hc4d1d06d, 32'h429932ef, 32'h43276478},
  {32'h4490dcc3, 32'h42ced158, 32'hc30503f5},
  {32'hc4ca8f10, 32'hc3951267, 32'hc3152129},
  {32'hc30b387c, 32'h440033d8, 32'hc2f321eb},
  {32'hc3e800f0, 32'h42ac1cfc, 32'h4314f94e},
  {32'h45044b10, 32'hc238b019, 32'h435e1c53},
  {32'hc4b629b4, 32'hc11b2271, 32'hc33efb94},
  {32'hc0711400, 32'h4277c6ac, 32'h40ee832c},
  {32'hc3b035d0, 32'hc389a7cb, 32'hc3c15067},
  {32'h44db6306, 32'hc2b6d2cb, 32'h3f84fc08},
  {32'hc51ad638, 32'hc42d2d5e, 32'hc219364c},
  {32'h44cd77e2, 32'h431b54aa, 32'hc24996e3},
  {32'hc384a89d, 32'hc2fe8d88, 32'h413d6107},
  {32'h44022cb6, 32'h42e8af4a, 32'h42a172c2},
  {32'hc32a22da, 32'hc2dd99b7, 32'h42bd19b4},
  {32'h4240f000, 32'hc393c729, 32'hc102dfb6},
  {32'hc4e6a9f9, 32'hc38c8c13, 32'hc37339db},
  {32'h44dfe49c, 32'hc2983ff7, 32'h43374a3b},
  {32'hc3b1fc18, 32'hc3921b51, 32'hc344abe0},
  {32'h450c5705, 32'hc25ae39f, 32'hc2cf252d},
  {32'hc4829e34, 32'h43ef168f, 32'hc1fa387e},
  {32'h44a083ee, 32'hc1692816, 32'h41eb4f93},
  {32'hc45d2cf6, 32'hc39eeb13, 32'hc29cbda4},
  {32'h442e4f95, 32'hc3c99d14, 32'hc2be8005},
  {32'hc4d72018, 32'hc3139875, 32'hc3e3e50f},
  {32'h44f09060, 32'h4245f8c9, 32'h42d28469},
  {32'hc4ef73b8, 32'h42b8ab0b, 32'h43a8b4e2},
  {32'h4510e188, 32'h4304365c, 32'hc3087bf4},
  {32'hc409e51c, 32'h42f5731d, 32'h43f9cd51},
  {32'h44e2e873, 32'hc3a43588, 32'h432f4360},
  {32'hc425667a, 32'h4391ad49, 32'h437797d9},
  {32'h44bbca82, 32'hc30958d5, 32'hc4244134},
  {32'hc474b860, 32'h43a3ab14, 32'h421934f0},
  {32'h4466484b, 32'h427fcfa6, 32'hc34f8aab},
  {32'hc4585c2c, 32'hc1d9bab0, 32'hc2faef09},
  {32'h44e850eb, 32'hc3a18ff7, 32'hc357990c},
  {32'hc471ae2c, 32'h43b48d41, 32'hc1e0144c},
  {32'h44113b16, 32'h4383a1ce, 32'hc393d3e4},
  {32'hc4dd332f, 32'hc2e6fa89, 32'hc28da9b8},
  {32'h449fc422, 32'hc299f5b1, 32'hc2894a91},
  {32'hc1e3cc80, 32'h438f7471, 32'hc30f5134},
  {32'h450acf64, 32'hc1d9d6c5, 32'h42f38d55},
  {32'hc431fb2c, 32'hc368d131, 32'h434c3623},
  {32'h44dd330f, 32'hc3a20a74, 32'hc2617f70},
  {32'hc50334f8, 32'h42a888ff, 32'h4087e09c},
  {32'h44f30bbe, 32'hc21decaa, 32'hc322a14c},
  {32'hc4347d8a, 32'hc3007dbe, 32'hc2306ae0},
  {32'h438bb7e0, 32'h4350bbb8, 32'hc3fdab0b},
  {32'hc50a7471, 32'h437ee562, 32'hc30637f7},
  {32'h446bb1a3, 32'hc3b30e3e, 32'hc339e5ab},
  {32'hc4ca6f65, 32'h427c0fd9, 32'hc389145e},
  {32'h4406b31b, 32'h4351b51d, 32'hc2a01a98},
  {32'hc3804c23, 32'hc2bc1d38, 32'h43dd922d},
  {32'h429fffb2, 32'h42a8af68, 32'h43587e56},
  {32'hc4d73385, 32'h43a71807, 32'h43973d66},
  {32'h439257ec, 32'h42843dac, 32'hc2d77363},
  {32'hc45f147e, 32'h436f70d5, 32'hc4034c47},
  {32'h44c43326, 32'hc31173cb, 32'hc38a650c},
  {32'hc4b7c627, 32'h42f2c33e, 32'h43822d0d},
  {32'h44fe168d, 32'h431e6e33, 32'h43e60d1b},
  {32'hc49726de, 32'h43af3740, 32'hc3c7aea6},
  {32'h448749d8, 32'h43c3c0a5, 32'hc337bd53},
  {32'hc5015fd9, 32'hc2139c2a, 32'hc30b09e8},
  {32'h451a9e48, 32'h434fea2a, 32'hc244fc8b},
  {32'hc43df3cb, 32'hc36a0a1d, 32'hc33f5b78},
  {32'h43ae437a, 32'hc39bfaef, 32'hc37c8e20},
  {32'hc46d591c, 32'hc21b0c45, 32'hc1f714c6},
  {32'h449f155b, 32'hc39595ca, 32'h4436cb91},
  {32'hc46c2fda, 32'h4359831c, 32'hc2badc81},
  {32'h4515fda8, 32'h425619cb, 32'hc2df5c6b},
  {32'hc3bf603a, 32'hc4206c2b, 32'hc385fc70},
  {32'h442de0f8, 32'hc3dba546, 32'hc30ffc5a},
  {32'hc501e29d, 32'h4225bfab, 32'hc2f4caad},
  {32'h4508531b, 32'h42bd77e9, 32'h42589009},
  {32'hc3c25abe, 32'hc3129e12, 32'hc1e1ffb0},
  {32'h451145c6, 32'hc28ed6d2, 32'h4239d942},
  {32'hc4b0d108, 32'h43383375, 32'h42e1d99e},
  {32'h44f9cf55, 32'hc3918b90, 32'h43950c82},
  {32'hc5139284, 32'h438dd641, 32'hc163e5e9},
  {32'h447ca84b, 32'hc2f06ae1, 32'h431bc7f0},
  {32'hc4621008, 32'h43b8df61, 32'h42fc6e72},
  {32'h4463a6ee, 32'hc2efe67d, 32'h42c51bd5},
  {32'h4372a9be, 32'hc39b4315, 32'h441ab0bc},
  {32'h451add83, 32'h42d5f63f, 32'h41e7a9c8},
  {32'hc4676c08, 32'h431ceb7d, 32'h4261cce3},
  {32'h449d8209, 32'hc33bd08c, 32'hc3107b66},
  {32'hc2a9d330, 32'h425e850a, 32'h4367556a},
  {32'h438504e2, 32'h43707e26, 32'h423fac71},
  {32'hc4fa2c46, 32'hc34b1eea, 32'h428ff888},
  {32'h4510df7b, 32'h436c40cb, 32'hc0e53191},
  {32'hc43daf42, 32'h43c4f3fd, 32'h428fb47e},
  {32'h451045f1, 32'hc3998aeb, 32'h43597556},
  {32'hc1b0e8a0, 32'h4256c566, 32'h437ac84f},
  {32'h44adb73f, 32'hc0ba60a1, 32'h42082d86},
  {32'hc4cda388, 32'hc2abd9c2, 32'h4284f504},
  {32'hc2774de0, 32'hc38769da, 32'h42fb8a95},
  {32'hc494b123, 32'hc19382c5, 32'hc1c34cf8},
  {32'h42add560, 32'h43a4cad4, 32'hc2855e71},
  {32'hc3636560, 32'h4293c924, 32'hc2ef9e95},
  {32'h4504ec98, 32'h43743c4c, 32'h415379fc},
  {32'hc4c8ddf4, 32'h43a652ba, 32'h42636b40},
  {32'h45079872, 32'h4356f136, 32'h42fb3a42},
  {32'hc4939e62, 32'hc339e6fc, 32'h4385f0ea},
  {32'h451da330, 32'hc2a66212, 32'h439d364e},
  {32'hc4bc0c4c, 32'hc3058ae2, 32'h43fd7fb0},
  {32'h448ce375, 32'h42dc0eda, 32'hc2a08c16},
  {32'hc50800a6, 32'hc2cd4ff7, 32'h4343cfb2},
  {32'h43e89b4b, 32'h4294dd13, 32'h424609e6},
  {32'hc48851a1, 32'hc27bd624, 32'h4360a9da},
  {32'h44707d6e, 32'hc37fa901, 32'hc2783097},
  {32'hc41a8574, 32'hc2e88fae, 32'hc32d987b},
  {32'h4497d7e8, 32'h41f2a298, 32'hc25c4b14},
  {32'hc4d123a8, 32'hc32bf543, 32'hc284cc5d},
  {32'hc38acb00, 32'hc33a4008, 32'h435b3523},
  {32'hc3dc4368, 32'h42978002, 32'hc3048c81},
  {32'h451811b2, 32'h4254a6c6, 32'h43f77dc4},
  {32'hc4bc5866, 32'hc39de09c, 32'hc2d1cd2f},
  {32'h44301a30, 32'hc3a3ca66, 32'hc31fd3e3},
  {32'hc49cbe3e, 32'h4392b536, 32'hc271e968},
  {32'h44812844, 32'h435c7981, 32'h4365d58b},
  {32'hc4a1afa0, 32'h42486db0, 32'h43086570},
  {32'h44b72bc5, 32'hc32d59a6, 32'h42730cf8},
  {32'hc3852270, 32'h435348ad, 32'h4309c8ee},
  {32'h446b9ab1, 32'h4344b292, 32'h423808ac},
  {32'hc4f2487f, 32'hc3d7377d, 32'h412df4a8},
  {32'h44117b7f, 32'h4365178f, 32'h438e7748},
  {32'hc4302553, 32'hc27dbb31, 32'h433b02f6},
  {32'h4493ef83, 32'hc389f974, 32'h423a0e8f},
  {32'hc4eec832, 32'hc2bccf89, 32'h43325e3d},
  {32'h43efd418, 32'hc2c048c8, 32'h42fe8412},
  {32'hc4a59653, 32'h422aa0d5, 32'h42983ec0},
  {32'h4294aee8, 32'hc23a27d8, 32'h43443031},
  {32'hc480723a, 32'hc04c31c4, 32'h437bda20},
  {32'h44b0e546, 32'h43a11330, 32'hc35429c0},
  {32'hc4e0c66e, 32'h43e1f7cc, 32'h4380307c},
  {32'h43af07fc, 32'h4361a49c, 32'h43da58a5},
  {32'hc48dd3cb, 32'h429aa6a1, 32'hc390548d},
  {32'h44cb1953, 32'hc36826c4, 32'h42be5e74},
  {32'hc4acb222, 32'h4337125d, 32'h4408e4b9},
  {32'h43a52d66, 32'h4381cbf9, 32'h4289b9af},
  {32'hc49ff134, 32'hc30ce0ea, 32'hc1fb88f0},
  {32'h441aade0, 32'hc3530617, 32'h4366058f},
  {32'hc4e0e820, 32'hc3919804, 32'h426c084a},
  {32'h44ac92cf, 32'hc308ef4a, 32'hc396ce01},
  {32'hc4f73b5d, 32'hc363df2b, 32'h42efcf6c},
  {32'h42128ae0, 32'h4306bca4, 32'hc3332282},
  {32'hc4c909f6, 32'hc2bf5482, 32'h42a9d11c},
  {32'h43f18ac8, 32'hc327ee16, 32'h440772e6},
  {32'hc3ac9414, 32'hc35d129e, 32'h4321f214},
  {32'hc2229940, 32'h43867455, 32'h4356078e},
  {32'hc4e133b5, 32'h42e88a65, 32'hc39854bf},
  {32'h43b35330, 32'h422c12d8, 32'h41bdba6c},
  {32'hc4b2db4d, 32'hc19eb616, 32'h3f8bc4bc},
  {32'h4486de43, 32'hc31919e0, 32'hc0d9d26b},
  {32'h43dba205, 32'hc2c39d09, 32'h3e4f0e71},
  {32'h44fd90af, 32'hc3437c39, 32'h426ea0c0},
  {32'hc45c5973, 32'hc2e86f89, 32'hc2238fb9},
  {32'h436ae4a1, 32'h42a1ab87, 32'h434255b9},
  {32'hc1cce700, 32'h4294c8de, 32'hc3099875},
  {32'h44eb6492, 32'h429cee41, 32'h43cf9b6b},
  {32'hc4893c98, 32'h41d69715, 32'hc25947ee},
  {32'h44d4cdce, 32'h43209f79, 32'h43a64620},
  {32'hc4b229b3, 32'h42ef4e26, 32'hc28f6cdd},
  {32'h44bf9a6d, 32'hc3d10e03, 32'h42d7930b},
  {32'hc4c3c510, 32'h42eee204, 32'h436fcbd6},
  {32'h44af6e3f, 32'hc32605fa, 32'h43362217},
  {32'hc33bee5b, 32'h43179009, 32'h437da9a9},
  {32'h44a59f65, 32'hbffaafe8, 32'h42b13261},
  {32'hc39a9baf, 32'h43f45f71, 32'hc2d438b3},
  {32'h439f83b4, 32'h41429c14, 32'h43b77cab},
  {32'hc4edcc18, 32'hc3148d99, 32'h432ee7ad},
  {32'h44802ca1, 32'h42bc6a0c, 32'hc3985e9c},
  {32'hc41fcb39, 32'hc1e5c0ea, 32'hc307cf17},
  {32'h449e5ea2, 32'h434affc1, 32'h43e7d030},
  {32'hc503b73c, 32'h43efc3ef, 32'h42b46a30},
  {32'h431cccf8, 32'h42b366a0, 32'h43d0fcf0},
  {32'hc50b0df3, 32'h43a1b99c, 32'hc3862e0c},
  {32'h44ef6ca6, 32'h42fdc578, 32'hc3e0fc9d},
  {32'hc4c1b2f3, 32'hc23d88c9, 32'hc2cc925a},
  {32'h44bcb89e, 32'hc33497fd, 32'h43b95dbe},
  {32'hc511ab11, 32'h42859ae4, 32'hc309f588},
  {32'h44480d28, 32'hc2ea6b94, 32'hc371b06d},
  {32'hc4eaea66, 32'h4395d893, 32'hc3774226},
  {32'h43206628, 32'h43857611, 32'h428030ea},
  {32'hc50d4870, 32'h437bdd7d, 32'hc375a801},
  {32'h4498bf50, 32'hc319fa34, 32'h4150dc9a},
  {32'hc4f645d4, 32'h422c3813, 32'h41d57320},
  {32'h43c5f014, 32'hc3af9e76, 32'h4316f5b4},
  {32'hc1332900, 32'hc1811140, 32'hc2f343ca},
  {32'hc20f4bb0, 32'hc3322e18, 32'hc29b4fa6},
  {32'hc4807054, 32'h42202a6e, 32'hc24dea1a},
  {32'hc1258f00, 32'h43fc2a36, 32'h43cafc47},
  {32'hc4f9814c, 32'h429dc249, 32'h4388b795},
  {32'h44433f56, 32'hc3695289, 32'h43166320},
  {32'h4317feca, 32'hc3991ed9, 32'h428c9d03},
  {32'h449c5b8b, 32'hc269b126, 32'h439aa754},
  {32'hc4aef726, 32'h42e753b0, 32'hc3ad5cc6},
  {32'h4486d2ba, 32'hc22d1091, 32'h42d545c0},
  {32'hc4ad3ac7, 32'h433e8da2, 32'hc2c76ee3},
  {32'h440bbc56, 32'hc3974d5e, 32'hc33df360},
  {32'hc2daa6e6, 32'h4382d90d, 32'h41c18a0e},
  {32'h42a867da, 32'hc385d595, 32'hc1e16875},
  {32'hc3df1977, 32'h43daa194, 32'h433f6edf},
  {32'h4502e1a9, 32'h434b6a12, 32'hc23fccbf},
  {32'hc50ddf12, 32'hc3340181, 32'h42e455d6},
  {32'h44e67f5d, 32'hc33c9d5a, 32'hc324fcb9},
  {32'hc50690af, 32'h42974b6b, 32'h43652018},
  {32'h44b7120c, 32'h440d16e0, 32'h4174de32},
  {32'hc3de30c4, 32'h42c9b52c, 32'hc3b67289},
  {32'h4265ca40, 32'h430cce68, 32'h424d65e5},
  {32'hc45e3ee0, 32'h43b11398, 32'h43450f84},
  {32'h43858793, 32'hc3b5ecc6, 32'hc23746f7},
  {32'hc50dfb99, 32'h42f6c531, 32'hc247c08b},
  {32'h450bd4cd, 32'h43964da0, 32'h41ac3976},
  {32'hc5003b5a, 32'h43c3e380, 32'hc35779ef},
  {32'h4518f141, 32'hc3ae09fb, 32'hc39608ce},
  {32'hc39399f8, 32'hc284f3d3, 32'hc260fe42},
  {32'h44b3399a, 32'hc13d0c16, 32'h42bbace3},
  {32'hc3af5800, 32'hc3055286, 32'h42d7df6f},
  {32'hc2a48f80, 32'hc3ca74b4, 32'hc3addeac},
  {32'hc34c6558, 32'hc250b420, 32'h4286703c},
  {32'h44c90627, 32'h43b0bb66, 32'hc322a5fd},
  {32'hc4e42e60, 32'h4390225e, 32'hc28cbfa1},
  {32'hc318b1c8, 32'hc3333b6a, 32'h43da662e},
  {32'hc50247f4, 32'hc1d78c51, 32'h4333dc34},
  {32'h445d60ce, 32'hc3cb07b9, 32'h43151062},
  {32'hc4ddeae0, 32'hc3047d83, 32'hc3a1b3c6},
  {32'h44e7a958, 32'hc390ef00, 32'h42eb8c7c},
  {32'h42f50060, 32'hc2be6e34, 32'h40886c6c},
  {32'h44865c0b, 32'h435994ea, 32'hc2ac06fd},
  {32'hc3c2f840, 32'h42628e20, 32'hbdc19a80},
  {32'h4424b419, 32'hc29656e9, 32'hc222e28b},
  {32'hc4a5bfa3, 32'h436f428b, 32'hc1bc5a11},
  {32'h4513b5df, 32'h427075b2, 32'h4375d9eb},
  {32'hc4bf90c6, 32'hc2da22f0, 32'hc3ae7868},
  {32'h44c90f40, 32'hc34fe574, 32'h4310c90d},
  {32'hc50d02b4, 32'h42acaa0f, 32'h434461c5},
  {32'h4434cd3a, 32'hc3a25231, 32'hc248c3f8},
  {32'hc4e51f5a, 32'h43f1a036, 32'h425b58c0},
  {32'h4453c604, 32'hc36c4e02, 32'h4298a1e7},
  {32'hc508a444, 32'hc30839b0, 32'hc2a51c90},
  {32'h441af641, 32'hc3e81baf, 32'hc3b6fad4},
  {32'hc4a53d3b, 32'hc40122e4, 32'hc38d7662},
  {32'h43d7913c, 32'h435f2148, 32'hc2da084f},
  {32'hc4e0dff1, 32'h43897e27, 32'hc38a60f2},
  {32'h448b6ae2, 32'h433c9ee9, 32'h4103b81e},
  {32'hc3005e2d, 32'hc3118fb4, 32'hc28fef36},
  {32'h44381e6c, 32'h41b4a0d8, 32'hc32cb701},
  {32'hc45385f4, 32'h42f43e10, 32'hc3af3ba6},
  {32'h4508a31b, 32'hc34cd6f0, 32'h432f63a3},
  {32'hc42fd313, 32'hc3403cb0, 32'hc4223d1d},
  {32'h43d3adf4, 32'h43506c5b, 32'h43a8f94f},
  {32'hc4e23ffe, 32'h4388a716, 32'hc388306c},
  {32'h45269f00, 32'h4394bb31, 32'h429b1d08},
  {32'hc4f5a431, 32'hc3a5f214, 32'hc3060daa},
  {32'h446bc7db, 32'h43b24383, 32'h434740af},
  {32'hc504a3cc, 32'hc0318ecc, 32'h43b6ee82},
  {32'h44a54113, 32'hc153c930, 32'h43660167},
  {32'hc4d1841f, 32'h43ec40cb, 32'h436f0aed},
  {32'h43fc1658, 32'hc2bc1c98, 32'hc341cd13},
  {32'hc3462ec0, 32'hc258ac76, 32'hc37aceaf},
  {32'h44827890, 32'hc391aab9, 32'h3d57c700},
  {32'hc4ab9ffa, 32'hc2f7ddeb, 32'hc233b232},
  {32'h43c1d263, 32'hc385cb6f, 32'hc2756dd1},
  {32'hc401bd7b, 32'hc2b2bd9e, 32'hc38c1855},
  {32'h4522ac3a, 32'hc19defc6, 32'hc3509c10},
  {32'hc42914d4, 32'h42c4f1b7, 32'hc3470f99},
  {32'h43d4276a, 32'hc3bdfa35, 32'h428f4cf3},
  {32'hc4dac742, 32'h427ea6c1, 32'hc25d6678},
  {32'h4401d4a8, 32'hc36e9b04, 32'h4215f133},
  {32'hc4d9bb97, 32'h41a360a1, 32'hc3cbe19f},
  {32'h44c56f44, 32'h4322a0d2, 32'hc2908056},
  {32'hc48413d7, 32'h42f21921, 32'hc2e32ab2},
  {32'h437f7b58, 32'h42d87c16, 32'h43aedd34},
  {32'hc4a45cde, 32'h43b923bf, 32'h43b27454},
  {32'h4483eeb3, 32'hc38e83bb, 32'hc22ec392},
  {32'hc4e96d82, 32'h41bddd2f, 32'hc2cc4747},
  {32'h45049735, 32'hc25cee8f, 32'hc3226256},
  {32'h4211d242, 32'hc35139d2, 32'h42fe1bc5},
  {32'hc3071070, 32'hc3a15738, 32'h41925db2},
  {32'hc50d31fc, 32'hc11f0b0e, 32'h4383dc2b},
  {32'h45196e9b, 32'hc36242d3, 32'h434a10c8},
  {32'hc2d0d729, 32'hbfbd180a, 32'hc143c8a4},
  {32'h445c307c, 32'hc1dbc321, 32'hc3c49df8},
  {32'hc50ce8d2, 32'hc1171f61, 32'hc3329f9b},
  {32'h44c356c0, 32'hc20eb65c, 32'h442d24b0},
  {32'h42a5f744, 32'hc32c3d62, 32'h43c1a67b},
  {32'h4431dd49, 32'h426dedca, 32'h430e7ed1},
  {32'hc3bd48e6, 32'hc1eb8dea, 32'hc2eb6867},
  {32'h44b75402, 32'hc37525ed, 32'hc31818f2},
  {32'hc431ac72, 32'hc2b1868a, 32'hc3f5f650},
  {32'h44a0dc95, 32'hc2fbe8d0, 32'hc3e65b7b},
  {32'hc4a400ee, 32'hc2717200, 32'hc2cc96db},
  {32'h44ed8a1d, 32'hc308cc68, 32'hc225fe6e},
  {32'hc507ec3e, 32'hc3996faf, 32'h4281585d},
  {32'h444280dc, 32'h43caae05, 32'hc3c0fb22},
  {32'hc4d79e8c, 32'hc3ad5b95, 32'hc1e780b6},
  {32'h43d26b00, 32'h42cd616f, 32'h433af966},
  {32'hc4f4a22d, 32'hc2ef16a0, 32'h4220b7ef},
  {32'hc4c8433a, 32'hc33b8ce5, 32'h4346aac6},
  {32'h44cab9c3, 32'h4306e9ea, 32'h43559296},
  {32'hc2eaa120, 32'h43519812, 32'hc2f19af5},
  {32'h4506942d, 32'hc34bd18a, 32'hc3717b8e},
  {32'hc4fe46fb, 32'hc40ccbf4, 32'h41d61b7a},
  {32'h4148cf40, 32'h436362a9, 32'h42d13867},
  {32'hc40a2fb0, 32'h43a4f4ae, 32'h4395201a},
  {32'hc3561668, 32'hc356591b, 32'hc3e7445b},
  {32'hc44cd418, 32'h44151688, 32'hc21ecbde},
  {32'h44dc2e9b, 32'h43853ed6, 32'h439d6c7a},
  {32'hc494751d, 32'hc354d6c3, 32'hc3b54c6d},
  {32'h429c36a0, 32'hc36e88a5, 32'h43350bd3},
  {32'hc3d53720, 32'hc328165e, 32'hc341f0e0},
  {32'h43f7d970, 32'h43b2177a, 32'h40f73356},
  {32'hc4fd9c4f, 32'h4279a07c, 32'h43a7d892},
  {32'h43fc5ea4, 32'h4317d77d, 32'h436effc2},
  {32'hc4b01037, 32'hc2d5cafa, 32'hc232c107},
  {32'h4522ab27, 32'h4354e3e9, 32'h42c36305},
  {32'hc494c9c6, 32'h42c93856, 32'h43274645},
  {32'h4482b980, 32'h43a54884, 32'h43f56189},
  {32'hc47d0c74, 32'h420a4782, 32'hc3dbf0bf},
  {32'h44e1592c, 32'h43139698, 32'h42850791},
  {32'hc4a015d8, 32'hc28753f0, 32'hc29d6afc},
  {32'h4512438b, 32'h42a7aa38, 32'h433b747f},
  {32'hc4edecc9, 32'h430596f7, 32'h432c5ed1},
  {32'h451b68f6, 32'hc3e7f031, 32'hc2469ef6},
  {32'hc488a375, 32'hc292680c, 32'h42c58432},
  {32'h450ebc7c, 32'hc3300ed4, 32'h43a4f623},
  {32'hc497e526, 32'h42296cc2, 32'h4416722d},
  {32'h4509125c, 32'h413e75a1, 32'h424f6eab},
  {32'hc4b1aa0e, 32'h42114275, 32'h4340c705},
  {32'h4508b848, 32'hc214bb46, 32'hc3b57049},
  {32'hc406447e, 32'h43ddd91c, 32'h42470ac0},
  {32'h4493cbc1, 32'h43386d6b, 32'hc3289762},
  {32'hc504bdf2, 32'hc3c178ac, 32'hc33aaed0},
  {32'h4484902d, 32'hc31c8f87, 32'h42f3e057},
  {32'hc48dc307, 32'h433af63f, 32'hc3b92333},
  {32'h4389e724, 32'hc2cd42dd, 32'h42299f63},
  {32'hc4f7e80f, 32'hc2e674bc, 32'h41beebe8},
  {32'h449bc513, 32'hc2822ffe, 32'h43571f16},
  {32'hc3963e54, 32'h440ac1e6, 32'hc229a60b},
  {32'h4395fa86, 32'h42a4e274, 32'hc2e52edc},
  {32'hc49ce4f6, 32'h41512f7c, 32'h4374bc50},
  {32'h4505d395, 32'h4113e922, 32'h4261cbae},
  {32'hc4cadf86, 32'h435b9712, 32'hc216d92f},
  {32'h4427a308, 32'hc37ca537, 32'hc256860c},
  {32'h4261d8c0, 32'h42bc2950, 32'h410c3bb2},
  {32'h44fa8113, 32'hc2897857, 32'h42865894},
  {32'hc51ce06c, 32'hc31c40b5, 32'h439a834d},
  {32'h44b3be10, 32'hc29dc223, 32'h435348ab},
  {32'hc4728373, 32'hc375f21d, 32'h44096ce0},
  {32'h43f37ff4, 32'hc1dee47a, 32'hc15f80ab},
  {32'hc40e36ce, 32'hc3a0f690, 32'hc3db5792},
  {32'h44aaaeda, 32'hc3e4b997, 32'hbf1c89f0},
  {32'hc506c270, 32'h4201c2c7, 32'hc3c48622},
  {32'h4509a434, 32'h423a45d0, 32'h438a3874},
  {32'hc4bbebc2, 32'hc3045426, 32'h43bd45a8},
  {32'h4416d8ea, 32'hc3b185d5, 32'hc426e3e7},
  {32'hc4a97860, 32'h412ed87c, 32'hc30730ee},
  {32'h4507a522, 32'hc3011380, 32'h42ff2667},
  {32'hc4640c74, 32'h43fbc8de, 32'h435011d7},
  {32'h44edeb26, 32'hc09f31aa, 32'h43a5ba43},
  {32'hc4d9dee2, 32'h41c75489, 32'hc20d26eb},
  {32'h4494b331, 32'hc2eab778, 32'hc1808d75},
  {32'hc505997d, 32'h43bf360f, 32'hc12a8756},
  {32'h446bdf58, 32'hc3e41d0d, 32'hc31a5d7b},
  {32'hc3af5db8, 32'h43c90a15, 32'h4393d6c6},
  {32'h45261ac4, 32'hc33a6aee, 32'h438da781},
  {32'hc530cff5, 32'h427be0a1, 32'h43ae153b},
  {32'h44a02607, 32'h41a41fa4, 32'h438b4099},
  {32'hc4bad97f, 32'hc2b39907, 32'h4299b641},
  {32'h44dcf08e, 32'hc321dde0, 32'hc2a6a3be},
  {32'hc51ce271, 32'h42a7f366, 32'h4381244b},
  {32'h44c16a8d, 32'h43575e86, 32'h4314f4db},
  {32'h40bd6140, 32'h42b106e4, 32'h425fcacf},
  {32'h43a6e9cd, 32'h426cf44b, 32'h42fce0b8},
  {32'hc4e67a1e, 32'hc2f87cf1, 32'h43c27067},
  {32'h444063c4, 32'hc18d3a0c, 32'hc34d84fa},
  {32'hc504ea6b, 32'hc3772217, 32'hc3da031a},
  {32'h44ff60d4, 32'hc2e8c19b, 32'hc30ff663},
  {32'hc4bef3d3, 32'hc3483ac2, 32'h424e171e},
  {32'h440c4a18, 32'hc39cbad9, 32'hc2550005},
  {32'hc4972589, 32'h42f9a16c, 32'h431e81b1},
  {32'h4512a880, 32'h43a29287, 32'h430cad29},
  {32'hc41509db, 32'hc369680a, 32'h436f87e8},
  {32'h4444b532, 32'hc16aeeb8, 32'h429a4b04},
  {32'hc3cefc53, 32'h435863d5, 32'hc0f16eec},
  {32'h4506a366, 32'h42afbdf7, 32'hc31c085d},
  {32'hc50963b5, 32'h40263030, 32'hc370946c},
  {32'h44d76e75, 32'h42cefb9d, 32'hc301ee88},
  {32'hc40fba54, 32'hc2d48f20, 32'hc33bdcc1},
  {32'h44c1c2c6, 32'h4231e8e9, 32'hc36a51be},
  {32'hc4d31b75, 32'h42985d01, 32'hc213ea18},
  {32'h44c3fc07, 32'hc3ece83f, 32'h432e56e1},
  {32'h416be700, 32'h435ece80, 32'h4369c3d1},
  {32'h44454fca, 32'hc3d49354, 32'hc3e4ff1d},
  {32'hc4769c4c, 32'h43b3231f, 32'h43500684},
  {32'h44ec962a, 32'hc355b47f, 32'hc300cc8b},
  {32'hc451da9a, 32'h43826cd8, 32'hc34e0b26},
  {32'h4471fd20, 32'hc3a2d102, 32'hc33e9304},
  {32'hc506914e, 32'hc3a0107e, 32'h420f14f0},
  {32'h44c716ce, 32'h42b73a5c, 32'h43a65f6e},
  {32'hc4f78ea2, 32'hc327176d, 32'h420c4cbf},
  {32'h442ed22b, 32'hc374e123, 32'hc24a86b1},
  {32'hc43f9f39, 32'hc2bb9227, 32'h43d49f67},
  {32'h441d4c9a, 32'h4388fe0c, 32'hc27a1073},
  {32'hc4971dde, 32'hc210254a, 32'h440955af},
  {32'h44bbfdd4, 32'hc2062556, 32'hc36a8ae2},
  {32'hc4ae5ae6, 32'h43248dfc, 32'h43bfbe17},
  {32'h44cb0e72, 32'hc3855c5f, 32'h425ad892},
  {32'hc4b6e77a, 32'hc32995c8, 32'h43f932c8},
  {32'h44a2ec8b, 32'h42cb08f6, 32'hc2f4dbfc},
  {32'hc435c420, 32'h42cd6dfe, 32'h43599d4d},
  {32'h446d4f7a, 32'hc256b55c, 32'hc3a6d52d},
  {32'hc509d74b, 32'hc2866234, 32'h42a705d7},
  {32'h4506f474, 32'h43906b4a, 32'h42933693},
  {32'hc490ed71, 32'hc1c3f814, 32'hc2de1de5},
  {32'h43c850d0, 32'hc39741e0, 32'h43400cb0},
  {32'hc50340a4, 32'h43f10729, 32'hc0265ce4},
  {32'h450d0bbd, 32'h42bb882e, 32'h43e4d12e},
  {32'h45019e3d, 32'hc2cdf316, 32'hc26767d0},
  {32'hc4d2780c, 32'h4404a185, 32'hc2b32aac},
  {32'h44c6ead5, 32'hc251d235, 32'hc1044a5a},
  {32'hc41880c0, 32'h4283016a, 32'h439325a9},
  {32'h44fa6a57, 32'h423bc210, 32'h43381df7},
  {32'hc4fa73f7, 32'h433f46f3, 32'h4358ed45},
  {32'h44ce1a7c, 32'h42664605, 32'hc390eb01},
  {32'hc4eeda3e, 32'h4404404a, 32'h427929fe},
  {32'h44f672bc, 32'hc2c10cd2, 32'hc245be3e},
  {32'hc4462a18, 32'hc34e589b, 32'h3da21380},
  {32'h44d3293d, 32'h4371a8dd, 32'hc3869f7e},
  {32'hc4bfeb6c, 32'h438c2a44, 32'h43c0955a},
  {32'h445f6c48, 32'hc2377ec6, 32'h4332de39},
  {32'hc50d9736, 32'h432b33b4, 32'hc3c98719},
  {32'h450d26df, 32'hc3455be9, 32'hc3445928},
  {32'hc4cda949, 32'h415f4ea8, 32'hc3ba0208},
  {32'h438042cc, 32'h3f5ee4d0, 32'hc3cc9a01},
  {32'h414f3900, 32'h434d8fde, 32'h4333f728},
  {32'h4463f97a, 32'hc29d19aa, 32'hc311930c},
  {32'hc40105a5, 32'h432601c1, 32'hc30531dc},
  {32'h44b30701, 32'hc2ff4dcb, 32'hc315daa9},
  {32'hc4e9d62d, 32'hc379a0b7, 32'hc2f223f1},
  {32'h45046011, 32'h4307d9ba, 32'hc3016d4c},
  {32'hc2de7c20, 32'hc3618d94, 32'h438999d7},
  {32'h4512d336, 32'hc2ea8168, 32'hc12a39b1},
  {32'hc412a260, 32'hc322950c, 32'hc2a46044},
  {32'h43cc5935, 32'hc3480738, 32'hc2b4b10c},
  {32'hc4092d8f, 32'hc2a02532, 32'hc302f300},
  {32'h44fd9157, 32'hc35df683, 32'h42107ccf},
  {32'hc4985e86, 32'h4311b27a, 32'h42f36b23},
  {32'h450ca50f, 32'h429bd5fd, 32'h423ce204},
  {32'hc4e19e0a, 32'hc3003196, 32'hc2b65b4b},
  {32'h44fa557b, 32'h433ac3cc, 32'hc3a2aec9},
  {32'hc438f9b4, 32'hc313241b, 32'hc17aa838},
  {32'h44768412, 32'hc1b5d737, 32'hc1a3673b},
  {32'hc4c96afc, 32'hc18dc1f6, 32'hc1881323},
  {32'h450c6812, 32'h43a87f9e, 32'hc28f11b8},
  {32'hc4d9f562, 32'h43fd7ab5, 32'h43948e58},
  {32'h45038f5c, 32'h4127d926, 32'hc2b40cde},
  {32'hc4882173, 32'h439a1396, 32'hc3a3a25c},
  {32'h440abc79, 32'hc3c4498d, 32'hc1e2f614},
  {32'hc2b31060, 32'h43c5a17e, 32'h43377ff6},
  {32'h42e2b6d6, 32'hc3c3933f, 32'hc388d82d},
  {32'hc4d37140, 32'hc317be39, 32'hc2b33408},
  {32'h43ee2ec9, 32'h4298c518, 32'h408862c4},
  {32'hc4de8006, 32'h43a63a6a, 32'h42163bd1},
  {32'h44e0e873, 32'h43643833, 32'h42b614c7},
  {32'hc38e9a68, 32'h428595e6, 32'h428235a4},
  {32'h44c2b8dd, 32'h4348637b, 32'h435a01f4},
  {32'hc4ee9140, 32'hc3742fac, 32'hbf705140},
  {32'hc37b9bf4, 32'hc232fa68, 32'h42297ed6},
  {32'hc494f0a6, 32'hc319ebde, 32'hc23afeab},
  {32'h448efea4, 32'hc2b6f38a, 32'hc3ad1fcb},
  {32'hc4c20273, 32'hc167b296, 32'hc361323d},
  {32'h44e0decd, 32'h43891306, 32'hc2d02863},
  {32'hc4a5276b, 32'h42aacc97, 32'h43a6bb53},
  {32'h43dc56d2, 32'h4379435a, 32'h4344e645},
  {32'hc4bc83c3, 32'hc39ea00b, 32'h423322c9},
  {32'h4392306c, 32'hc3c68b1c, 32'hc2ed2970},
  {32'hc4d05568, 32'hc307a0a1, 32'hc36a982e},
  {32'h44bfc1e3, 32'hc2fba203, 32'hc08fc37c},
  {32'hc4f09874, 32'hc33edef6, 32'hc3525bfd},
  {32'h4351c150, 32'h4124d3d7, 32'hc358ebdb},
  {32'hc487e2e1, 32'hc3add0b2, 32'h4210ac66},
  {32'h44ede0d7, 32'h43abc91e, 32'hc34d925c},
  {32'hc40202ae, 32'h43465099, 32'h43c91704},
  {32'h428e8298, 32'hc28dd3c9, 32'hc33f268d},
  {32'hc4e87c9e, 32'h4215a731, 32'h42739248},
  {32'h447cf9e6, 32'h42b8fa90, 32'hc379bbcc},
  {32'hc4c03014, 32'hc3b3e4de, 32'h4311392d},
  {32'h43ee3200, 32'h4309e569, 32'h44045945},
  {32'hc3fb77a2, 32'hc3a260a2, 32'h42c856e9},
  {32'h44219220, 32'h43e6aba2, 32'h43121dd9},
  {32'hc413242c, 32'h42b9d2a2, 32'h42c8a832},
  {32'h448ea328, 32'hc2cd3de3, 32'hc05e27e1},
  {32'hc4e23cf5, 32'h43a8a002, 32'hc403bd75},
  {32'h44efb98d, 32'h43d55f9f, 32'hc3cfff85},
  {32'hc4a76ab7, 32'h43ee551d, 32'h428075e9},
  {32'h4423e36c, 32'h3fd948e0, 32'h43277cf7},
  {32'hc50fb234, 32'h430e60bf, 32'hc2a3e39d},
  {32'h4515c60e, 32'hc3919116, 32'h43dd6d16},
  {32'hc50a55b5, 32'hc377bb33, 32'hc2ef84e4},
  {32'h44224909, 32'h43826fd3, 32'h421594c8},
  {32'hc4de65f7, 32'h43a7534e, 32'hc246b6a5},
  {32'h4415d6bc, 32'h4153945a, 32'hc253e9a8},
  {32'hc5069c90, 32'hc3715150, 32'hc313420d},
  {32'h44085d34, 32'h42df06a5, 32'h42c42db0},
  {32'hc499fcae, 32'hc15dde11, 32'hc2e4c14f},
  {32'h4414d9f5, 32'hc36befcd, 32'h43ca5bad},
  {32'hc4ec70c0, 32'hc322d0f6, 32'hc31c5f62},
  {32'h43a03005, 32'hc289facd, 32'hc2ecfd34},
  {32'hc3ab3ac0, 32'h439d304a, 32'h43193334},
  {32'h44293268, 32'hc34e083f, 32'hc335bd6d},
  {32'hc5183187, 32'h42f4fa1b, 32'h42538a09},
  {32'h45096026, 32'h41e5d031, 32'hc3b4fe22},
  {32'hc4b27d18, 32'hc3f52357, 32'h4343b7a7},
  {32'h444d14a7, 32'h430ba3de, 32'h423d7452},
  {32'hc4c509de, 32'hc3a03043, 32'hc356ee45},
  {32'h43cc8d28, 32'hc097beb0, 32'h41873caa},
  {32'hc4fecaf7, 32'hc27ba3f7, 32'h43b9cb68},
  {32'h44a8e179, 32'h439f651c, 32'hc322fabd},
  {32'hc4b9e102, 32'h433b530c, 32'hc361ede6},
  {32'h43eb7132, 32'h43a0e0a1, 32'h42932ae0},
  {32'hc3ef38d0, 32'h438eadda, 32'h435cd2ef},
  {32'h44d7e99b, 32'hc306ab25, 32'h42233d32},
  {32'hc4b93eb9, 32'hc1d3f6b1, 32'h43157e2b},
  {32'h45100c0f, 32'hc33bc9b2, 32'hc2ad82e4},
  {32'hc3b7f6a1, 32'hc42cd211, 32'h438556a0},
  {32'h4507246c, 32'hc28a3ad5, 32'hc19f4bb4},
  {32'hc41228bc, 32'h43ce7b28, 32'h42f4cc28},
  {32'h44e15a5c, 32'hc1d1e326, 32'h416c28e9},
  {32'hc4e15dd0, 32'hc1a0584f, 32'hc3279b0d},
  {32'h44b97c24, 32'h4345403d, 32'h40d384f4},
  {32'hc4281c85, 32'h427f130c, 32'h4305f978},
  {32'h44cb5ad1, 32'hc385cd55, 32'h4323d5e6},
  {32'hc506b867, 32'h43b41cf3, 32'hbfff2b50},
  {32'h4505af5f, 32'hc3a31606, 32'hc2267ce3},
  {32'hc35ab7c0, 32'hc2002306, 32'hc35dacc7},
  {32'h44cdb22e, 32'h43992754, 32'hc0eb7383},
  {32'hc50374c4, 32'h42221eac, 32'h4392a473},
  {32'h4498978e, 32'h4341f08b, 32'hc34b34a0},
  {32'hc4d8a0c9, 32'hc39fea09, 32'hc29dfbce},
  {32'h44d8f63b, 32'h426c8d09, 32'hc28ebd31},
  {32'hc4d3059e, 32'hc34fb200, 32'h4393fd76},
  {32'h450110a7, 32'h4391c343, 32'hc3881f27},
  {32'hc504e899, 32'hc39f60d4, 32'h4168af88},
  {32'h44c3259f, 32'hc32b53e9, 32'h437f30df},
  {32'hc488b93a, 32'hc1a8dc20, 32'h41ee4b13},
  {32'h45073840, 32'h42adde05, 32'hc328d34f},
  {32'hc4fabaae, 32'h42725a7b, 32'h435ab79e},
  {32'h43d50e0a, 32'h42fbd044, 32'h438e2b25},
  {32'hc4e7a182, 32'h44157c66, 32'hc288adc1},
  {32'h439e3e76, 32'hc384186f, 32'hc22efcdc},
  {32'hc35680f0, 32'hc39decd7, 32'hc35d611c},
  {32'h44b7fba4, 32'h42d3506a, 32'hc2653fc6},
  {32'hc491a759, 32'hc3caf85c, 32'hc1a72331},
  {32'h451488b7, 32'h42de6ca0, 32'h42bfcc35},
  {32'hc4b20cbe, 32'h43bd111b, 32'hc3040037},
  {32'h42f54a20, 32'h43a03f25, 32'hc331e493},
  {32'hc4dcca53, 32'h43aec4d0, 32'h42e43672},
  {32'h450851e6, 32'h42114667, 32'h429fab25},
  {32'h42b6579e, 32'h432b55af, 32'hc1c8ab48},
  {32'h439d3bf2, 32'h43de5f69, 32'h420f85f4},
  {32'hc3d1f5f0, 32'hc36b8714, 32'hc30fb29d},
  {32'h44757f7b, 32'h43136363, 32'h4310694f},
  {32'hc43453c8, 32'hc2d99862, 32'hc3f11a3e},
  {32'h446d581e, 32'h435da483, 32'hc3b69ce1},
  {32'hc442c2b9, 32'hc33d57a8, 32'h43863596},
  {32'h44fad07e, 32'hc31d7e55, 32'h4363555e},
  {32'h42d5c5b0, 32'h431ea0f8, 32'h4339f9fa},
  {32'h427b1850, 32'h42964c99, 32'hc33bd79f},
  {32'hc505c72e, 32'hc305cc1d, 32'hc3168c30},
  {32'h449184c7, 32'hc30f712f, 32'h43c8fe57},
  {32'hc4cbd310, 32'h43954386, 32'hc2ab3630},
  {32'h42bae280, 32'h42ed3b91, 32'h435529a8},
  {32'hc48817ec, 32'h40bf64af, 32'h429bcc8d},
  {32'h44f500ca, 32'hc31b93ec, 32'hc39f3581},
  {32'hc4ede2fb, 32'hc3bca349, 32'hc3dbd3df},
  {32'h450e65da, 32'h422c131c, 32'hc1d43529},
  {32'hc4f298e7, 32'h431a5e7f, 32'h42fcd53f},
  {32'h4492d574, 32'hc28835e4, 32'h42e9958e},
  {32'hc392a48f, 32'hc2208c6d, 32'h428799d5},
  {32'h44c4036a, 32'h4095c3de, 32'h43bfad06},
  {32'hc2ba5e70, 32'h42714b64, 32'hc30511f0},
  {32'h4506fda1, 32'h432742e1, 32'h435277cc},
  {32'h420d033c, 32'h4224ba54, 32'h43995f74},
  {32'h44e620e0, 32'h4386b215, 32'hc3a02f88},
  {32'hc4285b9a, 32'hc2324f86, 32'h436c7532},
  {32'h4476397a, 32'h43154d22, 32'h42e95d3c},
  {32'hc4ef53ec, 32'hc369779d, 32'h43dbcaf8},
  {32'h44a9630b, 32'h42fb79ba, 32'hc1234cca},
  {32'hc4f3e556, 32'h42f8aa4e, 32'hc28916eb},
  {32'h45250b97, 32'hc361c270, 32'h414d5b0a},
  {32'hc423073f, 32'hc1461d0d, 32'hc29abd4c},
  {32'h44802eec, 32'hc3084bc6, 32'h43b1b834},
  {32'hc4e2f976, 32'h439419da, 32'h43649729},
  {32'h44bebfe0, 32'h42a6470e, 32'hc2f57b74},
  {32'hc425928c, 32'hc3a4c281, 32'h43e7afad},
  {32'h42892e48, 32'h4333292e, 32'h4241651d},
  {32'hc4d5b3eb, 32'hc25bc027, 32'h42614307},
  {32'h4482fd72, 32'h4305b6c1, 32'h406e6fbc},
  {32'hc4f9d77c, 32'hc32876f5, 32'hc3052f88},
  {32'h43a10bf0, 32'h420ee46c, 32'hc30b8472},
  {32'hc4dbd326, 32'h4179d31e, 32'h430b3df6},
  {32'h44487ed1, 32'hc3808f8f, 32'hc33b471c},
  {32'hc419481e, 32'h434f179b, 32'hc29bf0ec},
  {32'hc33a29d4, 32'h4384fd35, 32'h4378ef7e},
  {32'hc4d97e46, 32'hc36b95b7, 32'h4358bef6},
  {32'h44a99af4, 32'hc375ea76, 32'h42e27489},
  {32'hc33d38f0, 32'h44290718, 32'h437a995e},
  {32'hc1ab92f8, 32'h4383eeac, 32'hc311199e},
  {32'hc4f39c3c, 32'hc2cc776a, 32'h436bb292},
  {32'h44fa5b1c, 32'hc25967fc, 32'hc2464b25},
  {32'hc4d7bfad, 32'hc27a2ee1, 32'hc398fdfe},
  {32'h4491a0b1, 32'hc1a54ef8, 32'hc26b11f7},
  {32'hc421897a, 32'h42bb6681, 32'hc31c9d6c},
  {32'h447c2516, 32'h4241169a, 32'hc298b1d9},
  {32'hc418669c, 32'hc327e119, 32'h438a5182},
  {32'h4447325b, 32'h437ef485, 32'h43350452},
  {32'h4221e780, 32'hc3a6a27c, 32'hc2b91265},
  {32'h44a2a611, 32'hc3fb46c9, 32'hc28c6a23},
  {32'hc50e6501, 32'h43383f26, 32'h435a5a23},
  {32'h44eeccd2, 32'h437eb1ea, 32'hc3e229e1},
  {32'hc400f4d7, 32'hc1a37069, 32'hc2a7282d},
  {32'h44df0201, 32'hc39a081d, 32'hc2f0fb62},
  {32'hc481cc82, 32'h4283c08b, 32'hc30e6bb7},
  {32'h4478d812, 32'hc20c1f63, 32'h41b3a9f9},
  {32'hc4c0c9bc, 32'hc2a67e68, 32'hc3aee65a},
  {32'h4463a8bb, 32'h42513796, 32'h42be4ba3},
  {32'hc3baf908, 32'h4208af5f, 32'h41d97fc8},
  {32'h439042c0, 32'hc4320f9c, 32'hc33c248b},
  {32'hc496781a, 32'h43af9b22, 32'hc2145cf8},
  {32'h44cfa28b, 32'hc255e700, 32'h4368c83b},
  {32'hc4abbb2c, 32'h435e3bd5, 32'h430c0bab},
  {32'h4431cf40, 32'h437dc8d4, 32'hc34911f1},
  {32'hc4dee671, 32'hc35a0900, 32'h437f724c},
  {32'h44cd6f9b, 32'h42b1381d, 32'hc18de8a7},
  {32'hc4148f89, 32'hc33bcfb3, 32'h433147dc},
  {32'h4449dd70, 32'hc3b93453, 32'h436703eb},
  {32'hc32dfab8, 32'h43068d1c, 32'h42adba22},
  {32'h4492bff1, 32'hc4038b2e, 32'h4400eb57},
  {32'hc4923abe, 32'h422287d2, 32'hc2926fd3},
  {32'h43dfd5b2, 32'h4218c00e, 32'hc20459ea},
  {32'hc44490b0, 32'hc3700e9e, 32'h42812905},
  {32'hc1240ec6, 32'h43f40538, 32'h43adbfdc},
  {32'hc45bb664, 32'h43245b35, 32'hc213ec47},
  {32'h44d5e339, 32'hc350c3af, 32'h4339a5e9},
  {32'hc4d1a574, 32'h43076302, 32'hc338df88},
  {32'h45078e42, 32'hc387fd45, 32'hc39c60ce},
  {32'hc4ecebd4, 32'h42e25bf2, 32'h434c2c8f},
  {32'h450e2926, 32'hc1b7bf18, 32'hc0fbbebf},
  {32'hc4267dc4, 32'h428aed56, 32'hc345b2c3},
  {32'h44f82ff1, 32'hc2d48d1c, 32'h42869a84},
  {32'hc3cc07ec, 32'h43234d12, 32'h43708395},
  {32'h44d1cbe8, 32'h434c218b, 32'hc362f99e},
  {32'hc47c26b8, 32'hbe547dcc, 32'hc31a5e2b},
  {32'h43a3879c, 32'hc28bf192, 32'h43627346},
  {32'hc4fc2ffb, 32'h433771fc, 32'hc2c9fd93},
  {32'h44ea57ae, 32'hc3558ba9, 32'hc3538e18},
  {32'hc42caecc, 32'h429ec332, 32'h42c2599d},
  {32'h44259cae, 32'hc36fe1b9, 32'hc1a384fd},
  {32'hc49aee34, 32'h42cfcb64, 32'hc2e631d5},
  {32'h4452c58c, 32'h4254e5b2, 32'h4355a1d3},
  {32'hc45ea9e6, 32'h429be520, 32'h4386a31d},
  {32'h450f9a1c, 32'hc21d41c3, 32'h434aff2f},
  {32'hc4857d1d, 32'hc3b513fa, 32'hc3bdaf76},
  {32'h43484260, 32'h43d95264, 32'hc388d264},
  {32'h4252f8a0, 32'hc344a504, 32'h43698738},
  {32'h44cb4ba3, 32'h42d65b05, 32'hc380c28a},
  {32'hc4637de3, 32'hc434e506, 32'h42afce11},
  {32'h450cd197, 32'hc37f4a00, 32'hc340771b},
  {32'hc4a260fe, 32'h41816595, 32'h43c03544},
  {32'h437120b0, 32'hc38d465b, 32'h3d9c4780},
  {32'hc4bc9c50, 32'h430922fa, 32'hc3285246},
  {32'h444ffbd8, 32'hc3636217, 32'hc3e928c8},
  {32'hc4ec2e63, 32'h438d523d, 32'hc348d1e7},
  {32'h441db67a, 32'h429b8732, 32'hc3c99467},
  {32'hc407fb29, 32'h422cf329, 32'h418755e2},
  {32'h44c67cbd, 32'h415ecd9f, 32'h418e8a9c},
  {32'hc4ae6f9a, 32'h421ce83d, 32'h43b14a19},
  {32'h4505cc2d, 32'h438d2bd1, 32'h432b8e39},
  {32'hc49a050c, 32'hc356b173, 32'hc1cf43e4},
  {32'h44330751, 32'h431da420, 32'hc4141b9a},
  {32'hc462c036, 32'hc310e322, 32'h435eb0ab},
  {32'h4514cb9d, 32'hc1ea29ab, 32'hc2d032d9},
  {32'hc47ffe30, 32'hc2df9fbc, 32'h41ffb9b2},
  {32'h44b78794, 32'hc211ad2a, 32'h420440de},
  {32'hc4fbf34a, 32'hc3028723, 32'hc3d750e7},
  {32'h43943776, 32'hc2e70e8e, 32'h4296376d},
  {32'hc4d167e4, 32'h44030f0f, 32'h4384b492},
  {32'h45106480, 32'hc3e8ef24, 32'hc2465265},
  {32'hc4f8d4e8, 32'h43b0fd12, 32'hc2ab2f90},
  {32'h44c8d3e4, 32'hc1a5dd0c, 32'hc3ad8094},
  {32'hc4d1d694, 32'hc38a9ad1, 32'h42e8b2ba},
  {32'h44342d2e, 32'hc29fa71d, 32'hc198597a},
  {32'hc4d4f9fd, 32'hc2f97c97, 32'h4320f2e9},
  {32'h450bfe3e, 32'h438a9c18, 32'hc3953ac2},
  {32'hc3cc1422, 32'h41ae0ad7, 32'h43142410},
  {32'h450e3768, 32'hc20365ab, 32'hc30c1048},
  {32'hc43f0626, 32'hc2930e4a, 32'hc387092c},
  {32'h447cabb2, 32'hc35b4b10, 32'hc36ed5d3},
  {32'hc432aeb2, 32'hc0e0cc4a, 32'hc3492a2c},
  {32'h44f7d987, 32'h42636a37, 32'h439e8f69},
  {32'hc4685672, 32'h43313f9b, 32'h42bb542b},
  {32'h4503a467, 32'hc3478ffc, 32'h41e2ee3c},
  {32'hc4ab7791, 32'hc23ebc1a, 32'h41d33dc2},
  {32'h450a687d, 32'hc32bee69, 32'hc1a79cc4},
  {32'hc4ecb37c, 32'hc398cb06, 32'h42515394},
  {32'h447c78a9, 32'h43a6b100, 32'hc28a002a},
  {32'hc47a5f7a, 32'h433cf665, 32'hc2b304d1},
  {32'h44898042, 32'h423d10d4, 32'h431b1b1e},
  {32'hc51050a2, 32'hc2a3559a, 32'hc36c92e5},
  {32'h4479c3e6, 32'hc26ef53f, 32'h42c408f2},
  {32'hc4c6295e, 32'h43f72ac9, 32'h42b4c632},
  {32'h448be9e4, 32'h411d30e0, 32'hc31dac73},
  {32'hc37bb6c8, 32'h4274d76a, 32'h42f74a72},
  {32'h45039c29, 32'hc3842408, 32'h43d5317b},
  {32'hc42c2d82, 32'h413c3f92, 32'h436aebdd},
  {32'h45125de9, 32'hc349c585, 32'h42161a73},
  {32'hc4ea3238, 32'h42c6a68e, 32'h419bb615},
  {32'h44504014, 32'hc33b8ecc, 32'hc32d2c09},
  {32'hc4b27c86, 32'hc3da0e1d, 32'h43890b72},
  {32'h44134665, 32'hc122554f, 32'h42604f77},
  {32'hc3b14760, 32'hc3243724, 32'h437b1251},
  {32'h4330f4ff, 32'h434ac3b6, 32'hc31edaa4},
  {32'hc4d8bdc7, 32'hc1d877da, 32'h41a0237a},
  {32'h441ecc8c, 32'h432262fa, 32'hc3dd7985},
  {32'hc5142a0b, 32'hc31cbd5b, 32'h42f35681},
  {32'h43942d60, 32'hc3782e77, 32'h42b31c3e},
  {32'hc4e5d598, 32'hc2efb973, 32'h43e621ea},
  {32'h4473d388, 32'hc26767e2, 32'h43882a06},
  {32'hc4a1fafa, 32'hc349f39b, 32'hc2008add},
  {32'h437071c0, 32'h42a906cf, 32'h431ef84e},
  {32'hc515e612, 32'h42b0f2d5, 32'h41a4b164},
  {32'h44ab0edd, 32'hc314e096, 32'h42a6d987},
  {32'hc4c9f956, 32'hc372530a, 32'h42a0e6bf},
  {32'h448a5aa7, 32'hc26d7724, 32'hc36135f1},
  {32'hc4a2ccce, 32'h4282eb33, 32'hc302dd47},
  {32'h44666e33, 32'h429ea58b, 32'h43251812},
  {32'hc4dbdb87, 32'h41aa2d29, 32'hc3e5a798},
  {32'h452836c9, 32'h4308ffee, 32'hc31fa87b},
  {32'hc50ac90d, 32'hc40db44c, 32'h42b56aaf},
  {32'h44c30763, 32'h420213ed, 32'h42bb7d4f},
  {32'hc38e5938, 32'hc37bd4d7, 32'h420691d4},
  {32'h447aee9b, 32'h420d151d, 32'h43466527},
  {32'hc4ec153e, 32'h42efde08, 32'h432082a0},
  {32'h4449ba90, 32'hc314554e, 32'hc39b34a5},
  {32'hc4ce152e, 32'hc2d92830, 32'h42588413},
  {32'h44f672b2, 32'h4331d6a2, 32'h42b30a11},
  {32'hc400daf8, 32'hc1f3214a, 32'h43a0c7c3},
  {32'h451571ce, 32'hc39804d7, 32'hc2bd3563},
  {32'hc48b861d, 32'h431af000, 32'hc221108d},
  {32'h445450cb, 32'h4284717e, 32'hc2db0e51},
  {32'hc468c75c, 32'h43d854a3, 32'hc3926e0c},
  {32'h44818e87, 32'h42b55b93, 32'h432523af},
  {32'hc426d93f, 32'hc2f738d2, 32'hc3672f62},
  {32'h44e77fd8, 32'hc3dd7ff8, 32'hc39dfe3d},
  {32'hc2839d48, 32'hc3586ab2, 32'hc1dd1b04},
  {32'h44d006b8, 32'h431d4efd, 32'h433d6a8d},
  {32'hc434e437, 32'h42cd3d35, 32'hc348f3f9},
  {32'hc2ecdab8, 32'hc3a0debc, 32'hc24129c0},
  {32'hc37d7fd8, 32'h42bad29f, 32'hc278974c},
  {32'h44eb663e, 32'h4382b27c, 32'hc24883ec},
  {32'hc514ded5, 32'h40615d10, 32'h42bf27c7},
  {32'h4482d134, 32'hc28baf27, 32'hc1e39339},
  {32'hc4d01d66, 32'hc39196ef, 32'h407405c2},
  {32'h4521cac1, 32'hc3925d81, 32'h4289c7c5},
  {32'hc522b3fa, 32'h43eb1473, 32'hc199d73a},
  {32'h44c348e7, 32'h430459ed, 32'hc4060f3c},
  {32'hc45c097b, 32'h4243e6cb, 32'hc2ca6733},
  {32'h44a2bec2, 32'hc0e11bb5, 32'h4383bad5},
  {32'hc304d37d, 32'h42a72443, 32'h432685ec},
  {32'h44ded18e, 32'hbeb7ce40, 32'hc2d70222},
  {32'hc4288366, 32'hc29f788f, 32'hc239ac32},
  {32'h445a348f, 32'hc2d7de31, 32'hc24ce569},
  {32'hc4f0678e, 32'h431cb904, 32'h4244392d},
  {32'h440623ac, 32'h4203b2cd, 32'hc34fe469},
  {32'hc4bff7d6, 32'hc0a9a6a3, 32'hc30357e7},
  {32'h44d0fae7, 32'h4384b082, 32'hc36934bf},
  {32'hc4a12c92, 32'hc08f0750, 32'hc25b662a},
  {32'h44434184, 32'hc39c216c, 32'hc3294668},
  {32'hc49699fe, 32'hc36bab4b, 32'h4358c232},
  {32'h45128b4a, 32'hbfd5f164, 32'h42d5f1c3},
  {32'hc514f914, 32'h42911091, 32'hc355eb5a},
  {32'h44c7fc50, 32'hc1f9c507, 32'h42cfb87a},
  {32'hc4e44f96, 32'h42997c7d, 32'hc351e0e9},
  {32'h44f18e96, 32'hc38915b1, 32'hc3c2f690},
  {32'hc25b2500, 32'h41f9f205, 32'h439e05c1},
  {32'h44bf0076, 32'hc342cc57, 32'hc319a1ee},
  {32'hc3f00a7d, 32'hc3a0b820, 32'hc2c5556d},
  {32'h450cddc7, 32'h418c8338, 32'h42868ea9},
  {32'hc4cfe76a, 32'hc0ba25d7, 32'h43a29159},
  {32'h4503835b, 32'h43047139, 32'h43b24375},
  {32'h434a1900, 32'hc38f0de5, 32'h424ea67e},
  {32'h43d87ac6, 32'h42f2ac0e, 32'hc3387fec},
  {32'hc4859c82, 32'h432cee27, 32'hc2da7bd9},
  {32'h43adc336, 32'hc33d9f92, 32'h40c78af6},
  {32'hc48915c6, 32'hc25d1078, 32'h43af2363},
  {32'h451e2ad6, 32'h43c8a416, 32'hc1861ba3},
  {32'hc4e5e775, 32'hc321b35e, 32'hc0ff0667},
  {32'h44367145, 32'hc2eca98a, 32'h42a28ca9},
  {32'hc4412114, 32'h43a53835, 32'hc1ef1600},
  {32'h43a852fc, 32'hc227d4c1, 32'hc2e6d645},
  {32'hc3c5d9ca, 32'h41bafbda, 32'hc3c697c3},
  {32'h44f62a8b, 32'h434f1087, 32'hc2f2ee01},
  {32'hc511d4de, 32'hc2ff09fa, 32'h43277892},
  {32'h441a09cc, 32'hc16f7b08, 32'h428a1f27},
  {32'hc4170f46, 32'hc3b01a48, 32'h419070a8},
  {32'h44ed060a, 32'hc2ee7146, 32'h43241f4c},
  {32'hc35e3130, 32'hc384e22f, 32'h421f6173},
  {32'h43e699f4, 32'hc1a7ee0d, 32'h43933e58},
  {32'hc4e0e5a8, 32'hc3c72f52, 32'hc33a2609},
  {32'h442fe67e, 32'hc392cdfa, 32'hc3a787a6},
  {32'hc50a552d, 32'h42ae09fa, 32'h4087a344},
  {32'h44cfcf3c, 32'h432956cf, 32'hc4084bab},
  {32'hc4def39a, 32'hc2f41816, 32'hc417ef88},
  {32'h44aaa8b7, 32'hc332978c, 32'hc18aae61},
  {32'hc3a4b890, 32'h41e2bef5, 32'hc2f33947},
  {32'h43bb4560, 32'h4057e89a, 32'hc20067e7},
  {32'hc4b60c73, 32'h41c1228d, 32'h4352bd3a},
  {32'h44caa8bd, 32'hc2e5e60e, 32'h41acdd61},
  {32'hc42fc8f6, 32'h40fd9c46, 32'hc3502a71},
  {32'h43d0e3ba, 32'hc3846d63, 32'h422abe88},
  {32'hc3b0f7fc, 32'hc2c4e967, 32'hc32df04e},
  {32'h4400f158, 32'hc3a865c8, 32'h4397d144},
  {32'hc48bdbf3, 32'h4297153c, 32'hc38f34a0},
  {32'h44f92cc0, 32'h427a4f17, 32'hc37b4301},
  {32'hc4d6cbf2, 32'h42a88bc0, 32'hc24294c4},
  {32'h449f28b0, 32'hc217cf1b, 32'h4329c022},
  {32'hc52e7a34, 32'h428b8ee8, 32'hc2708f38},
  {32'h43a72138, 32'h42a3031a, 32'h42bc15e4},
  {32'hc4b15724, 32'h43a815f7, 32'hc204f653},
  {32'h4410a853, 32'h4321ad15, 32'h433fcc7a},
  {32'hc4823a36, 32'hc229dbb5, 32'h43f3d252},
  {32'h44937444, 32'hc38af55e, 32'h425303dc},
  {32'hc4e712a2, 32'hc3e38431, 32'h432215d7},
  {32'h44e84864, 32'h42d18d7c, 32'h43cd8507},
  {32'hc49f9215, 32'h42d97900, 32'hc399758f},
  {32'h44cae39b, 32'hc29d5dfc, 32'hc2b0571b},
  {32'hc4b2c982, 32'h42e267c9, 32'h42a7fd16},
  {32'h44d0b64e, 32'h4382fc4c, 32'h42058435},
  {32'hc4aa385f, 32'h3ef38b40, 32'hc43288bf},
  {32'h44c5f4da, 32'h424c70ef, 32'h42dcf767},
  {32'hc5052cb1, 32'hc3628855, 32'h423c3456},
  {32'h45004536, 32'hc32e6fca, 32'h43281e97},
  {32'hc48532d5, 32'hc3871316, 32'hc39ba074},
  {32'h44c529e2, 32'h439f1ef9, 32'hc205c223},
  {32'hc459837d, 32'hc302bebe, 32'hc30feb9f},
  {32'h429780d0, 32'h4382d01d, 32'h434ade74},
  {32'hc49ec43b, 32'hc3279b11, 32'hc3ad4d5a},
  {32'h440e2abe, 32'hc22385d3, 32'h4361a378},
  {32'hc495904c, 32'hc1a5a3e6, 32'hc3af4f81},
  {32'hc3bb138c, 32'h43af1e0a, 32'hc379bb54},
  {32'h44472632, 32'h43a91e07, 32'h43758cf9},
  {32'hc4d04fe2, 32'hc3a4e462, 32'hc237e860},
  {32'h44e4dc84, 32'hc2cc7bb9, 32'hc2a23b5b},
  {32'hc5073066, 32'hc11e89c5, 32'hc28507c9},
  {32'h441484d8, 32'h41eb8f0f, 32'hc37a2b00},
  {32'hc3ceb108, 32'hc110dbc4, 32'hc2ddbb6d},
  {32'h43d61196, 32'hc3751045, 32'h440de954},
  {32'hc512a99d, 32'hc2c3f875, 32'hc23384ca},
  {32'h44872afe, 32'h4341c9be, 32'hc381a029},
  {32'hc35700e0, 32'hc221a0a1, 32'h42dadd40},
  {32'h44c2443b, 32'hc36dfb62, 32'hc18c909a},
  {32'hc4b0de8b, 32'h4371164e, 32'hc2eb2530},
  {32'h448934ea, 32'hc257c0a8, 32'h4364a415},
  {32'hc3a9653c, 32'h4327cc76, 32'h42d79308},
  {32'hc1bb65c0, 32'hc242b275, 32'hc06ec598},
  {32'hc49f954a, 32'h431c6980, 32'hc324e48e},
  {32'h43786944, 32'h42d59ec9, 32'h43b890ca},
  {32'hc4cd432c, 32'hc2176d8b, 32'h43030aab},
  {32'h450166dc, 32'h43bc64d6, 32'h437ccc5e},
  {32'hc413df8e, 32'h42c4d466, 32'hc317bc81},
  {32'h45049ec3, 32'hc32228c2, 32'h433ca8d7},
  {32'hc4a3b492, 32'h42875469, 32'hc2c9d956},
  {32'h429983b0, 32'hbef7b770, 32'h43b456fa},
  {32'hc43938a8, 32'hc31c4598, 32'hc2b051fb},
  {32'h44b55774, 32'hc29a06b1, 32'hc383b91b},
  {32'hc4aae0a7, 32'hc35b5309, 32'h43affced},
  {32'h4504b185, 32'hc386a85a, 32'h42c1bd5e},
  {32'hc4d2fa4c, 32'h40a7450d, 32'hc3906528},
  {32'h4514591d, 32'h408da0b3, 32'hc38dcac7},
  {32'hc50d2be4, 32'hc20b8739, 32'h4315aa5f},
  {32'h44e3aa34, 32'hc29b3d9b, 32'h42c71d64},
  {32'hc4b85e5c, 32'hc3a14317, 32'hc1424d93},
  {32'h44ac5e2e, 32'h4397feca, 32'h42edcb29},
  {32'hc4319782, 32'h42cf272d, 32'hc3873626},
  {32'h444868b4, 32'hc3229a85, 32'hc0b5968d},
  {32'h431b6bc0, 32'hc3170edc, 32'hc36e3296},
  {32'h44154428, 32'h4308a91d, 32'hc33949bd},
  {32'hc4e06b2b, 32'h42c5867d, 32'h432e5d58},
  {32'h4443bb20, 32'h432c51ee, 32'h41244024},
  {32'hc4eb3dc9, 32'hc34823aa, 32'h42b7808b},
  {32'h432cb100, 32'h4309ff9a, 32'h438cc590},
  {32'hc49ea6c9, 32'h433966a5, 32'hc3252be6},
  {32'h44da7b3a, 32'hc40fe8ac, 32'h441b837a},
  {32'hc46d92f8, 32'h413c580e, 32'hc304ba84},
  {32'h4456de8c, 32'hc310b81f, 32'hc2ebb8e6},
  {32'hc4e43b68, 32'hc32152a9, 32'hc25b134f},
  {32'h447be81e, 32'h423e816d, 32'hc400dbbd},
  {32'hc4e536ea, 32'hc2742453, 32'h42af0cf7},
  {32'h44b054db, 32'h4037d55f, 32'h433f95f5},
  {32'hc50f8b80, 32'h43dbc0ee, 32'hc2b9e99b},
  {32'h43a848cc, 32'hc3787161, 32'h4308ddd4},
  {32'hc4f0a160, 32'hc3de7a69, 32'hc393e8c7},
  {32'h43a3bdc8, 32'h41c83767, 32'hc2f074a7},
  {32'hc4db8de8, 32'h431fa75a, 32'hc33e8734},
  {32'h448e53a9, 32'hc227b2be, 32'h4304d71b},
  {32'hc4d7cd30, 32'hc3ae2e5c, 32'h42938367},
  {32'h444dcf6c, 32'hc3f83a5e, 32'h42ddb606},
  {32'hc41ff392, 32'hc368ad5d, 32'hc3691d6d},
  {32'h44929e3c, 32'h428fbdd1, 32'h4227a27e},
  {32'hc324cb74, 32'hc39eb44d, 32'hc1e6ddb9},
  {32'h43be19f0, 32'h432ed5fd, 32'h43e87e32},
  {32'hc4f0a0a0, 32'hc1e30476, 32'h418a816e},
  {32'h442807e9, 32'hc290f330, 32'hc39c53f5},
  {32'hc446ef38, 32'h4184c4ab, 32'h40763708},
  {32'h436d1b2c, 32'hc398c7d7, 32'h42dfca5e},
  {32'hc393fad8, 32'h420cbe5f, 32'h438c3a8f},
  {32'h448f2c67, 32'h431348da, 32'h40950d9e},
  {32'hc3aab544, 32'hc309ac9f, 32'hc266aeba},
  {32'h447ec60e, 32'h4393e4ee, 32'hc22341cc},
  {32'hc4c6edd4, 32'hc2f8fb7c, 32'h424ec620},
  {32'h44db26d1, 32'h4353cb40, 32'h428bbe78},
  {32'hc47d8748, 32'hc3914069, 32'h4251844a},
  {32'h45030a21, 32'h43bc9431, 32'h438e9e28},
  {32'hc2840f40, 32'hc36a0e48, 32'h430a0b3a},
  {32'h443b9088, 32'hc297ad2c, 32'h429c6935},
  {32'hc43ba415, 32'hc4180915, 32'hc2cf7722},
  {32'h449aa986, 32'h42c84975, 32'h4337d4a4},
  {32'hc41bd718, 32'hc28c3a01, 32'hc33c22b6},
  {32'h44d0b8b9, 32'h42d914a1, 32'hc386ec13},
  {32'hc290db2b, 32'h42a75999, 32'h43030a4c},
  {32'h44a98012, 32'h432f63e2, 32'hc3f501f8},
  {32'hc4bed5fd, 32'h437dc2a1, 32'h43539c5d},
  {32'h450bb6b3, 32'h430bdce6, 32'hc2bd85f8},
  {32'hc4d9d0b2, 32'hc353a1bb, 32'hc39fef1b},
  {32'h44ecc259, 32'h4379ad5b, 32'h43d63339},
  {32'h411aa140, 32'h43b43539, 32'hc3cc737f},
  {32'h45033754, 32'hc32c75e9, 32'hc3465752},
  {32'hc3ff9399, 32'h438283b1, 32'hc1c1d2ec},
  {32'h450c94e2, 32'h4373153d, 32'hc402f6ad},
  {32'hc4ee6e1e, 32'hc17828c1, 32'hc04182f0},
  {32'h430d7ad0, 32'h42b3ff07, 32'h410ec072},
  {32'hc5217095, 32'hc2559581, 32'h43611e0a},
  {32'h444c799e, 32'h42668245, 32'hbf70cb64},
  {32'hc395ac96, 32'hc3a7ae33, 32'h425d36e7},
  {32'h44e504b2, 32'hc2da6178, 32'hc36bb7b4},
  {32'hc43fccc8, 32'h43d8e5ed, 32'h437e1f68},
  {32'h4430a994, 32'h42ebaf72, 32'hc2bd919f},
  {32'hc3a8020a, 32'hc0d4ba3c, 32'hc2a656ca},
  {32'h425db8c0, 32'h40922994, 32'h4217371c},
  {32'hc4f7c163, 32'h42071814, 32'h43cf7ee2},
  {32'h41903a80, 32'h43845a7c, 32'hc349bcbb},
  {32'hc2d2cb60, 32'hc2ec89de, 32'h43cb9233},
  {32'h44dd6fb2, 32'hc19e6fda, 32'hc2cff458},
  {32'hc500108b, 32'hc3c155a7, 32'hc1757234},
  {32'h44db890a, 32'h42e335ee, 32'hc2452d04},
  {32'hc43e3495, 32'hc1e08af8, 32'h426d1391},
  {32'hc008ec80, 32'hc3835113, 32'h43238283},
  {32'h431c0b00, 32'h42623b5d, 32'hc30581a6},
  {32'hc184b760, 32'h42f6baff, 32'hc2f3225f},
  {32'h435659f0, 32'hc34160b8, 32'hc37bfe1c},
  {32'hc37daebe, 32'hc335c241, 32'h435346af},
  {32'hc37cf030, 32'hc3853ab1, 32'h43811eba},
  {32'h44588c11, 32'hc2e0c269, 32'hc33a2fd8},
  {32'hc4f0693c, 32'hc25507ac, 32'h44599e8e},
  {32'h4520474c, 32'hc36948c9, 32'hc302be33},
  {32'h43d29406, 32'h42c6f4d6, 32'hc35fd38c},
  {32'hc450112b, 32'h42070978, 32'h42b53a82},
  {32'h4484cf59, 32'hc340a7f6, 32'hc126b7c7},
  {32'hc4a4c50d, 32'h4336cf16, 32'h4358cf0e},
  {32'h4409a272, 32'h4296bb80, 32'h41ac8836},
  {32'hc4802ddf, 32'h4233b00e, 32'h431e6a7a},
  {32'h445c6d06, 32'hc1bc3436, 32'hc306dff4},
  {32'hc4a333a8, 32'h43bb14f0, 32'hc2f1599e},
  {32'h44176980, 32'h424062b0, 32'h431440b3},
  {32'hc499932e, 32'hc32b7307, 32'h42a7297a},
  {32'h4510e893, 32'h42b7712a, 32'hc2bcfefb},
  {32'hc4222d78, 32'h41411d72, 32'hc331eb68},
  {32'h429834d0, 32'h43ee0514, 32'h4291ab40},
  {32'hc3fe4c74, 32'hc34c3375, 32'h43910ac5},
  {32'hc373f900, 32'h42ec8dea, 32'hbde9bb60},
  {32'h4457cb70, 32'hc290f0f5, 32'h41fb58c2},
  {32'hc4fde072, 32'h41e27581, 32'h4379e777},
  {32'h4449b448, 32'hc3a8b4e1, 32'hc30e1b57},
  {32'hc4104fe8, 32'h4302685a, 32'hc2ce4727},
  {32'h44af1d8a, 32'hc37ca3eb, 32'h4377b415},
  {32'hc4f838ff, 32'hc1024dff, 32'h43a741c7},
  {32'h44b270ec, 32'hc20e5582, 32'h42392389},
  {32'hc4d530b8, 32'hc265dd80, 32'h427f8fb1},
  {32'h44127f70, 32'hc280cc7f, 32'hc37b89aa},
  {32'hc449db9a, 32'hc3060dcf, 32'h42687a04},
  {32'h435d6476, 32'h4363343e, 32'h435ab0ea},
  {32'hc469f444, 32'hc379c894, 32'h439a71c2},
  {32'h44e6b164, 32'h4304f717, 32'h43278488},
  {32'hc4cbe177, 32'h40f11e7e, 32'hc268f738},
  {32'h4501ff50, 32'hc26142e3, 32'hc3447734},
  {32'hc450be13, 32'hc344c73f, 32'h4384b4a9},
  {32'h4392a248, 32'h42b00e3a, 32'h4319bb9e},
  {32'hc3eeea58, 32'h4356d751, 32'hc306dee5},
  {32'h44c7cdd0, 32'h41a7113c, 32'hc3bc59d4},
  {32'hc48deb9f, 32'h4335ea00, 32'hc2c57b7e},
  {32'h44141e7c, 32'hc281e5ed, 32'h4313ed03},
  {32'hc4939922, 32'h42340b7e, 32'hc2955c64},
  {32'h44fd2490, 32'h41b42290, 32'h42d5ede5},
  {32'hc4050d78, 32'hc3d8e1ac, 32'h41fa26b6},
  {32'h44aeb7be, 32'hc18d2bcc, 32'h42e52160},
  {32'hc4a73d8c, 32'hc358beeb, 32'hc3473a83},
  {32'hc30a2e7e, 32'hc31d2c8d, 32'hc3c65272},
  {32'h4289ccf0, 32'hc38bd68f, 32'h4390f25b},
  {32'h4521eea2, 32'hc333da52, 32'hc22a02cc},
  {32'hc49bf87b, 32'hc2c8a26d, 32'h41234d37},
  {32'h442cc99e, 32'hc375bb75, 32'hc2ea29cd},
  {32'hc4895d9b, 32'hc2e10e9f, 32'h409968e5},
  {32'h442dee24, 32'hc385b6aa, 32'hc2d8dc3a},
  {32'hc3e908a5, 32'h43105741, 32'h439d1a47},
  {32'h44c3b7b6, 32'h419251f6, 32'hc2df5be9},
  {32'hc511ef36, 32'h419f1b65, 32'hc295d18a},
  {32'h4436e702, 32'h43029bef, 32'h428f979b},
  {32'hc4c2d760, 32'hc350703c, 32'hc3073ce4},
  {32'h44d0f78c, 32'h42c660da, 32'h4306dee9},
  {32'hc4816639, 32'h43a89f2c, 32'hc2d8c0ae},
  {32'h44b74523, 32'hc29065db, 32'hc413deca},
  {32'hc49d60e2, 32'h43170ac6, 32'hc36bcf78},
  {32'h41dbce60, 32'h4357ae53, 32'h419d1b00},
  {32'hc47a6312, 32'h430f4549, 32'hc34adcef},
  {32'h43a471f8, 32'hc311f550, 32'hc340ca0e},
  {32'hc4fa2802, 32'hc31d6770, 32'hc2e7620e},
  {32'h44294eba, 32'h41a854b2, 32'hc3742dde},
  {32'hc4e5f637, 32'h4329404a, 32'h42ed42b6},
  {32'h43f658b4, 32'hc4107548, 32'hc33b6b8e},
  {32'hc4d7db4c, 32'hc2d0f7af, 32'h41f680a6},
  {32'h44964329, 32'hc2ff534d, 32'hc17049a9},
  {32'hc4d6f03d, 32'hc3581f86, 32'h41295b3c},
  {32'h434b89f8, 32'h42116df8, 32'h424c86cc},
  {32'hc43f279a, 32'h438bcf70, 32'h4307542a},
  {32'h446346e2, 32'h43fe226a, 32'h3ffda810},
  {32'hc45cd9d2, 32'h430d3bbf, 32'h4312e7fb},
  {32'h4415b300, 32'hc41c8d4e, 32'h4304056b},
  {32'hc48e2e44, 32'h438ccf60, 32'hc3c9c3dc},
  {32'h444c5def, 32'h430ceec7, 32'hc2f22f90},
  {32'hc4a21a5a, 32'hc3b752b0, 32'h43377397},
  {32'h449f29c3, 32'hc2a7e15c, 32'h431fcbb1},
  {32'hc4b0708f, 32'hc3599c3a, 32'hc352289a},
  {32'h43a7844e, 32'h4288a2d9, 32'h42fb12e3},
  {32'hc4b53d3b, 32'hc0472ca8, 32'hc2ed6950},
  {32'h44982265, 32'hc2c9d725, 32'h42dc0841},
  {32'hc4e26307, 32'hc22ea0c4, 32'h431c0411},
  {32'h44675df7, 32'hc2d5bc42, 32'h43544aef},
  {32'hc514dc82, 32'h43b28bc6, 32'h43e37138},
  {32'h450e9850, 32'hc08edeb0, 32'h42debcdd},
  {32'hc4493f10, 32'hc3b90429, 32'hc18df2ca},
  {32'h44d7eb03, 32'hc3123d52, 32'hc3bb2398},
  {32'hc459b475, 32'h424f7005, 32'h410e3f81},
  {32'h44501655, 32'hc2ae0d10, 32'hc3f2ccdf},
  {32'hc4064a00, 32'hc302814a, 32'h41c1919d},
  {32'h4397f85e, 32'hc3b1fd73, 32'hc33ff994},
  {32'hc396a7b0, 32'hc0a21cc3, 32'h43848d03},
  {32'h4474ac82, 32'h4205332c, 32'h435cf88f},
  {32'hc42477da, 32'hc230af24, 32'h42e2db74},
  {32'h4483fc91, 32'h421b0502, 32'h432b7e09},
  {32'hc284bcb8, 32'h437afebe, 32'hc3b6a231},
  {32'h442ade60, 32'h4341fdbe, 32'h42a537bf},
  {32'hc4d49c0d, 32'hc3817a76, 32'hc3269535},
  {32'h441be0d2, 32'hc3b3d862, 32'hc2cd81cd},
  {32'hc522df18, 32'hc3647161, 32'h4388619a},
  {32'h44b7d78d, 32'hc2ec3aef, 32'hc3267f47},
  {32'hc50b748c, 32'hc199b923, 32'h4310ffac},
  {32'h449eef76, 32'hc3ce7689, 32'h43b85376},
  {32'hc4166422, 32'h4251fdcc, 32'h42b92385},
  {32'h43915eee, 32'h4381ee95, 32'hc37f7c45},
  {32'hc4552dba, 32'h43904f31, 32'hc34537ac},
  {32'h451277ac, 32'h42bfb6b4, 32'h424d6df0},
  {32'hc4a765b4, 32'h4314ca84, 32'h41b454c8},
  {32'h448d3fff, 32'h438216ed, 32'hc2c4406f},
  {32'hc4669042, 32'h437142bf, 32'hc3938f20},
  {32'h450c7f0f, 32'h43076cd1, 32'h430b9102},
  {32'hc4d03070, 32'hc3808111, 32'h42b21d2a},
  {32'h44674e0b, 32'h438d15fc, 32'hc38c59b3},
  {32'hc48e1fd8, 32'hc2b3e4b9, 32'hc32a0097},
  {32'h44ae6f45, 32'h43900b03, 32'hc08f92f0},
  {32'hc497821c, 32'h41f9fcf6, 32'hc0495da2},
  {32'h44d03be2, 32'hc2aba047, 32'hc36aa1f0},
  {32'hc485d09d, 32'h41eba848, 32'hc12bec86},
  {32'hc3766ec8, 32'h41292a78, 32'h42a01420},
  {32'hc42e14c4, 32'h439cdff0, 32'h43a795f1},
  {32'h44adf829, 32'hc05457c4, 32'h438f4d6f},
  {32'hc4795b46, 32'hc36d603a, 32'hc2a75cfe},
  {32'h448be89e, 32'h43cd0aa9, 32'h43d899e0},
  {32'hc46d6efc, 32'h4327a9ad, 32'h42b6bf4c},
  {32'h43fa81fc, 32'h432a7618, 32'hc3e22831},
  {32'hc470f0dc, 32'h42516ab1, 32'h40a529a4},
  {32'h444b9f4d, 32'hc39900d4, 32'h430aade8},
  {32'hc4843faa, 32'h429f4252, 32'hc2a46c79},
  {32'h44a127bb, 32'h431d07b9, 32'hc32923b2},
  {32'hc456855a, 32'h430e48ae, 32'hc380526a},
  {32'h44bc6eb3, 32'hc40c16b0, 32'h439e993f},
  {32'hc3ea2e75, 32'hc3056571, 32'h43905994},
  {32'h44ad6e86, 32'h436e5b9f, 32'hc415ea90},
  {32'hc438331c, 32'hc3c37f5e, 32'h432c8abb},
  {32'h44ec6892, 32'h42f95879, 32'h41b01c5f},
  {32'hc3e91e71, 32'hc294bef3, 32'hc380fcac},
  {32'h44bb5363, 32'h42ac390c, 32'hc24e856e},
  {32'hc48cfb8c, 32'hc3ca2732, 32'h42b223f0},
  {32'h44c466b0, 32'h42a49c71, 32'hc216401e},
  {32'hc39ecaf0, 32'hc33bff72, 32'hc3258a22},
  {32'h44b4185b, 32'h43926413, 32'h441391c8},
  {32'hc3dbcc68, 32'h43ad83da, 32'h43109298},
  {32'h44f21aa7, 32'hc2e96f63, 32'hc33b6e74},
  {32'hc4945f8d, 32'hc35779aa, 32'h437526fa},
  {32'h45130486, 32'h421ff7e6, 32'hc34538a1},
  {32'hc4031e10, 32'hc302fbe6, 32'h42ea0a3b},
  {32'h44bdff8e, 32'hc36210ef, 32'h43a3571c},
  {32'hc4dfd0ee, 32'h42168823, 32'hc35fdcb2},
  {32'h4405d646, 32'h427f920c, 32'h43829c47},
  {32'hc47e5402, 32'hc2c2412e, 32'hc2ed4374},
  {32'h44b7eba7, 32'h4382170d, 32'hc305d539},
  {32'hc4c08307, 32'h423e2e66, 32'hc2915320},
  {32'h450aa2e2, 32'hc317db16, 32'hc3f1c480},
  {32'hc4c62510, 32'h412fa413, 32'hc373b19d},
  {32'h44375473, 32'h430dbde1, 32'h439237c1},
  {32'hc35a511c, 32'h43f660c9, 32'hc071e8ac},
  {32'h4508f3ca, 32'h42ace69d, 32'h42381f24},
  {32'hc483c79c, 32'hc3537d93, 32'hc1b0610d},
  {32'h44fd2752, 32'hc30525e2, 32'h4185e3fb},
  {32'hc4a71f71, 32'h43d0cf1a, 32'hc2b4025e},
  {32'h44b85869, 32'hc28c22a2, 32'hc23e707b},
  {32'hc4dea9ac, 32'h43cc0f0c, 32'h42a8733d},
  {32'h451e5e2c, 32'h433f98da, 32'hc29550b4},
  {32'hc4744780, 32'h439cfdd5, 32'h429c7ee2},
  {32'h43e9c298, 32'h438b28b0, 32'hc3da056e},
  {32'hc3762d40, 32'hc3912125, 32'hc338a8c7},
  {32'h45046ef1, 32'h42511987, 32'h42a06990},
  {32'hc40499bd, 32'h43169b1c, 32'hc1657657},
  {32'h44eadec6, 32'h430c8571, 32'hc38c345b},
  {32'hc3945220, 32'hc22b0dbe, 32'h434f87b5},
  {32'h450e5d23, 32'hc3a93102, 32'hc1ebb576},
  {32'hc4ff395b, 32'hc22249df, 32'hc2a8e85e},
  {32'h448479bd, 32'hc3522c4e, 32'hc2bca549},
  {32'hc4d396e7, 32'hc3486a08, 32'h42158f3f},
  {32'h4479d459, 32'h433ea728, 32'hc2d95927},
  {32'hc4741ec0, 32'h43d205b8, 32'hc3261b34},
  {32'h44707458, 32'h4400b4bd, 32'h43db54e0},
  {32'hc501b7e4, 32'h43b3c730, 32'h42f92d92},
  {32'h4511529f, 32'hc3a1fb23, 32'hc2827276},
  {32'hc4d57822, 32'hc11413de, 32'hc31a5d07},
  {32'h4505c7e5, 32'hc34134c6, 32'h42484271},
  {32'hc47fec97, 32'hc3d54b2b, 32'h43a6c8d5},
  {32'h448d8402, 32'hc391aae3, 32'h42fb7df1},
  {32'hc515f3c5, 32'hc39d0d94, 32'hc345fe39},
  {32'h45213e0a, 32'h443c58c3, 32'h437025d2},
  {32'hc40441fa, 32'hc34bdd21, 32'hc2febcef},
  {32'h44eefded, 32'hc0ef05ce, 32'h436e0e06},
  {32'hc404b0ad, 32'h433d6b30, 32'h43bb46c6},
  {32'h453537e1, 32'h4355d861, 32'h43dcf414},
  {32'hc20b0ca0, 32'hc35738c1, 32'hc39c2f9c},
  {32'h435232e4, 32'h42c24006, 32'hc3bb4e0c},
  {32'hc50e30f2, 32'hc38a35d4, 32'h4184bd38},
  {32'h44bde661, 32'hc38e15e2, 32'h42bd50c4},
  {32'hc408fa79, 32'h43091b88, 32'hc2d2ea31},
  {32'h44768a00, 32'hc354afc7, 32'hc23b61e1},
  {32'hc485c7b2, 32'hc2e39780, 32'h40ff94c6},
  {32'h44c75ab7, 32'hc0615634, 32'h4247a670},
  {32'hc3ca70f0, 32'hc30e3d78, 32'hc20fc98e},
  {32'h43a3ddd8, 32'hc348a653, 32'h43b5cba2},
  {32'hc4f039a3, 32'hc205bdbe, 32'hc417908f},
  {32'h4503f588, 32'hc252ba8b, 32'hc350df66},
  {32'hc4d65bce, 32'h41edb41a, 32'h43234837},
  {32'h44a0d01b, 32'h4326bd7a, 32'h43afcc9b},
  {32'hc3d38afa, 32'h43068473, 32'h43c91508},
  {32'h44095918, 32'hc3e43bff, 32'hc2078461},
  {32'hc4a3bc64, 32'hc25daa6e, 32'h42e81bb8},
  {32'h44adb241, 32'h409a09c1, 32'h4279e492},
  {32'hc3cc6af0, 32'h429972b3, 32'hc39e8e0c},
  {32'h4505b62f, 32'h4356b80e, 32'h4402d423},
  {32'hc4e04c90, 32'hc38e1db3, 32'hc19bfc22},
  {32'h446d2513, 32'h438b6951, 32'hc0eea9df},
  {32'hc484e2af, 32'hc2445ebb, 32'hc1810b79},
  {32'h44cabab8, 32'hc3886c54, 32'hc2fb5ccb},
  {32'hc4a85cb6, 32'hc345e669, 32'h42e41689},
  {32'h451b4dbb, 32'hc2e62d6a, 32'hc3090e87},
  {32'hc3d66528, 32'hc3a4ef18, 32'hc328469b},
  {32'h44d7bc2b, 32'h438ead8b, 32'hc38ea047},
  {32'hc49156f1, 32'h42321d4c, 32'hc3804373},
  {32'h44f69037, 32'hc3486642, 32'h43094a94},
  {32'hc46c88dc, 32'hc3124ceb, 32'h43a2965b},
  {32'h448ea622, 32'hc34ece85, 32'h425bba57},
  {32'hc4f94e2a, 32'h43314202, 32'hc3de3297},
  {32'h44e1c255, 32'h42e376ab, 32'h4262e7e1},
  {32'h4536f544, 32'h4255cf55, 32'hc2b61fa6},
  {32'hc50ffb59, 32'hc30d668a, 32'hc31a8d97},
  {32'h44a0bc9d, 32'h408d82c0, 32'hc2d1b302},
  {32'hc38179ae, 32'hc1d1779c, 32'hc3313d32},
  {32'h44432f64, 32'h43db514b, 32'h433e4303},
  {32'hc5131dff, 32'hc35d4719, 32'hc35e21dc},
  {32'h4418d6f8, 32'hc3031418, 32'hc1dfe3e7},
  {32'hc467c7c8, 32'hc32bbcc4, 32'h435d1700},
  {32'h45049a54, 32'hc2ca3539, 32'h43564536},
  {32'hc5092963, 32'h432c78ce, 32'h4345f08e},
  {32'h451ab6b2, 32'h41eee074, 32'hc25083ab},
  {32'hc46ca3e3, 32'hc389e352, 32'h42f23c71},
  {32'h44acb1ea, 32'h4308111c, 32'hc3ab7a08},
  {32'hc3b50570, 32'hc3b408e4, 32'hc32ee6a1},
  {32'h45217a04, 32'h41db0ee2, 32'h3dc57120},
  {32'hc4971b50, 32'h42d4404e, 32'hc2f9cd97},
  {32'h44f1273f, 32'h434e21a4, 32'hc33f58c6},
  {32'hc4605df4, 32'hc1f85a9f, 32'h43a3774e},
  {32'h45128d5b, 32'hc31e7f3b, 32'hc28d295a},
  {32'hc50c5550, 32'hc2aeb05e, 32'hc29e2a3a},
  {32'h4378a982, 32'h433503f2, 32'hc14cf66c},
  {32'hc43290ff, 32'hc325adf5, 32'hc30ddd8f},
  {32'h451a5ad8, 32'h43ebe050, 32'h43939ebb},
  {32'hc4d34ac8, 32'hc306fed9, 32'hc3bb49b5},
  {32'h44812dd0, 32'h42da1442, 32'hc32cde50},
  {32'hc41323c0, 32'hc3272f33, 32'hc2879514},
  {32'h44f4d0f7, 32'hc2c9d83b, 32'hc3cd0cec},
  {32'hc4869c38, 32'h42324277, 32'h42cacc9a},
  {32'h44ea74cf, 32'hc3529fbb, 32'hc2f865ed},
  {32'hc41651a2, 32'h4393eab2, 32'hc3883be7},
  {32'h45190b7a, 32'h43b17e7d, 32'h432d33f0},
  {32'hc37f5a4c, 32'h430797d6, 32'hc393b33a},
  {32'hc31d9a14, 32'h4253fc58, 32'h43e6d063},
  {32'hc46be214, 32'h439af85a, 32'h438c1eba},
  {32'h44c2a966, 32'h438c71a9, 32'hc11faba8},
  {32'hc4fec295, 32'hc3860198, 32'hbf96ef22},
  {32'h446428b7, 32'hc34dfd72, 32'h43b43d37},
  {32'hc4f718c3, 32'hc23f3831, 32'h436fb4c0},
  {32'h450571bd, 32'h424fc780, 32'hc09acd50},
  {32'hc48d1c76, 32'h42e041a8, 32'hc31474bf},
  {32'h43cb466c, 32'h42de3841, 32'hc264866f},
  {32'hc4e45fc3, 32'h4401705e, 32'h434c96f9},
  {32'h4333d6a0, 32'h426fad05, 32'h42bbcbc3},
  {32'hc4c543f2, 32'hc3998fec, 32'hc31f87dd},
  {32'h4521e6a2, 32'hc326d2dc, 32'h42eaf104},
  {32'hc4ea7db5, 32'hc356c423, 32'h438ef56d},
  {32'h450259b8, 32'hc2f240cb, 32'h411a3127},
  {32'hc4563671, 32'h433a57ab, 32'h43b816d1},
  {32'h42bc34d0, 32'h42fb9916, 32'h42669784},
  {32'hc487ba90, 32'h43269655, 32'h438706ea},
  {32'h4239a385, 32'hc288fab8, 32'hc32a8742},
  {32'hc484ef00, 32'h4368d6ab, 32'h42cf3e51},
  {32'hc2506040, 32'h426a41e5, 32'hc3c208f1},
  {32'hc3d8c17d, 32'hc23c2905, 32'hc2c1f46f},
  {32'h44c7f87c, 32'hc36a7477, 32'hc39b422b},
  {32'hc4b74636, 32'hc39fabd7, 32'hc2904b8d},
  {32'h45127478, 32'h431db34e, 32'hc124fc47},
  {32'hc4bccdee, 32'h438bd64d, 32'hc350414e},
  {32'hc4fdf700, 32'h43509206, 32'hc3337a18},
  {32'h448dbf2c, 32'hc336523d, 32'hc401b706},
  {32'hc4892e1f, 32'hc3191166, 32'hc32a8a97},
  {32'h43c06f9f, 32'hc2ce1568, 32'hc363b8d8},
  {32'hc4ea7c11, 32'hc2bf3cbc, 32'hc3551f51},
  {32'h449a196c, 32'hc15df5ad, 32'hc2f0856e},
  {32'hc4881f11, 32'h435aa599, 32'hc22aa91e},
  {32'h4457d6cc, 32'hc2826eb3, 32'hc3d63814},
  {32'hc427d5a8, 32'hc2d9cdff, 32'hc2e5e96b},
  {32'h436d6d40, 32'hc263b5bf, 32'hc068af70},
  {32'hc40b7f28, 32'h4379247b, 32'h43fdacf8},
  {32'h43b9038c, 32'hc39b19de, 32'h42978bc7},
  {32'hc41a679a, 32'hc3aded6f, 32'h42debabb},
  {32'h44ad92ec, 32'h4283e9fb, 32'hc3521537},
  {32'hc4c763b6, 32'h43276460, 32'h434eaaac},
  {32'h43fe7180, 32'hc1b82460, 32'hc21e320f},
  {32'hc4d01b88, 32'hc31f302a, 32'h4355880c},
  {32'h43b26d9c, 32'h42826459, 32'h42709b7e},
  {32'hc4f2d777, 32'hc2a86533, 32'h426a3c26},
  {32'h445d545f, 32'h42abd0d7, 32'hc3b02a06},
  {32'hc5076406, 32'hc28cf274, 32'h414627f4},
  {32'h447ff6db, 32'h4359a988, 32'h428758b5},
  {32'hc446e1e6, 32'h42e7426f, 32'hc1bcfae7},
  {32'h44a19acf, 32'hc3985305, 32'hc329170d},
  {32'hc4f27af4, 32'h424485e5, 32'h438c3b86},
  {32'h44f6a1fe, 32'h435c0fe6, 32'hc0b42858},
  {32'hc450189f, 32'hc2e1f913, 32'h433c4e12},
  {32'h44b1b818, 32'hc322d024, 32'hc3b695cf},
  {32'hc509c5bc, 32'h432585c2, 32'h429d7d79},
  {32'h44929d8d, 32'hc38e0a73, 32'hc306f7dd},
  {32'hc37c72e0, 32'hc071f550, 32'h439c8c7d},
  {32'h43a374fc, 32'hc2536457, 32'hc2ac0ba7},
  {32'h44758490, 32'hc306c5f0, 32'hc2401397},
  {32'hc36eaef0, 32'h420cfa15, 32'h42ae7567},
  {32'h450b50c8, 32'hc1cf0c7e, 32'hc32e99a2},
  {32'hc43f3963, 32'h420cf10a, 32'h43cefbc1},
  {32'h44de4f03, 32'hc37cacb2, 32'hc3cd4fc5},
  {32'hc39e1419, 32'h43664fc8, 32'h4370d5bc},
  {32'h4286a85c, 32'hc1cc14cd, 32'hc3201be7},
  {32'hc503f400, 32'hc4174dad, 32'h438c7d93},
  {32'h445eae04, 32'h430ec6f2, 32'hc3f71ffb},
  {32'hc4f84446, 32'hc37a4d6c, 32'hc32939ae},
  {32'h44cc11b1, 32'h42512dd5, 32'h429f37a1},
  {32'hc4b364b8, 32'hc2d12647, 32'h4297cd46},
  {32'h44ebfec1, 32'hc13d9343, 32'h43282036},
  {32'hc49c2e2e, 32'h434655b9, 32'hc2c5f867},
  {32'h42200afc, 32'hc2bfa7db, 32'h4301ec14},
  {32'hc48f5a78, 32'hc255cdd1, 32'h43ac0840},
  {32'h44be7e0a, 32'h43e1a2d7, 32'h424f0f1c},
  {32'hc50a5328, 32'h43b24b36, 32'h40c57458},
  {32'h44ac5f79, 32'h43caf385, 32'hc33e2a8e},
  {32'hc5075af2, 32'h43779aa0, 32'hc38ab1d7},
  {32'h44753858, 32'hc3ad564b, 32'hc39f471b},
  {32'hc175dd00, 32'h4368ba42, 32'hc25cc2a6},
  {32'h44995ec2, 32'hc2a196ab, 32'hc2fa8b84},
  {32'hc2c8ec90, 32'h4189ebe3, 32'h43835812},
  {32'h4441c214, 32'h42f9f788, 32'h421f19fa},
  {32'hc51115d2, 32'h43af102e, 32'h43246cda},
  {32'h44d9c88d, 32'h4276c142, 32'hc2633adc},
  {32'hc426d306, 32'h43b8c6d5, 32'h43594795},
  {32'h43bca0b5, 32'hc2490375, 32'hc3cdfe3d},
  {32'hc5045393, 32'hc32f3cfd, 32'h4360980f},
  {32'h448d2422, 32'hc39e1f0f, 32'h4273e483},
  {32'hc48947bc, 32'hc2fc4a62, 32'hc231e40f},
  {32'h447c0668, 32'hc41e4313, 32'hc2a3f73c},
  {32'hc42cfb83, 32'hc4068172, 32'h43409e75},
  {32'h43dcb9d5, 32'hc2d9199a, 32'hc35b49bf},
  {32'hc4f193f2, 32'hc35173dc, 32'h42f4ba48},
  {32'h445670a0, 32'h42661968, 32'h41c57402},
  {32'hc4b35e58, 32'hc3c8bb67, 32'h41999767},
  {32'h451acde3, 32'h426bbd72, 32'hc38304d3},
  {32'hc48525c1, 32'hc2720b3d, 32'h43452622},
  {32'h4480415c, 32'hc3b0f8aa, 32'h43474adf},
  {32'hc4dd556a, 32'h427443f3, 32'hc297ff64},
  {32'h44935990, 32'hc3586c56, 32'h439b7b42},
  {32'hc4e958fb, 32'hc2e5fea1, 32'h41f44244},
  {32'h42fe229c, 32'hc35f4371, 32'h42977aaa},
  {32'h42a3dfb0, 32'hc32baafd, 32'hc197a41f},
  {32'h450612f5, 32'h43636752, 32'h43c0c731},
  {32'h42cb4e00, 32'h4362460c, 32'h43aa6719},
  {32'h4468c1c2, 32'h42896d2b, 32'hc3ff2cba},
  {32'hc5031167, 32'hc3657c62, 32'h42dca640},
  {32'h451edb01, 32'h42c51828, 32'hc2bf2b64},
  {32'hc502bef4, 32'hc29e95d3, 32'hc2cb76aa},
  {32'h44f73b40, 32'h4239dab6, 32'h436209db},
  {32'hc4deeaf6, 32'h41b9d6e2, 32'hbf0f7758},
  {32'h43f708f8, 32'hc20f82a0, 32'hc381913e},
  {32'hc5050f02, 32'h433647f6, 32'hc2a7e854},
  {32'h450e4ef2, 32'hc38a28e5, 32'hc3e6bc6c},
  {32'hc4e810b7, 32'hc1c93d30, 32'hc3f23e06},
  {32'h44e4d872, 32'h437a9858, 32'hc27f1312},
  {32'hc4965985, 32'h4177d6e8, 32'hc1ef6487},
  {32'h438b9260, 32'hc3eee06b, 32'h42304a37},
  {32'hc3ea5d1e, 32'h43b075f0, 32'h41a42485},
  {32'h44f09df5, 32'h4368289c, 32'hc29dd0e4},
  {32'hc50e9817, 32'hc322a0ed, 32'h4122da50},
  {32'h441e11b7, 32'h41aca100, 32'hc2bd8b1c},
  {32'hc5001e1a, 32'hc3c37226, 32'hc1a2b0a7},
  {32'h44252f24, 32'h439652d8, 32'hc33f2262},
  {32'hc48c79a0, 32'hc38abc91, 32'hc203750d},
  {32'h44f3d921, 32'h417fed72, 32'h43261900},
  {32'hc511f372, 32'hc39d6e37, 32'hc2f68c4c},
  {32'h44a57314, 32'h429a57a7, 32'h42b900dd},
  {32'hc420aa86, 32'hc1f2dd66, 32'hc2fd5849},
  {32'h44b0b778, 32'h42a81847, 32'h425236c9},
  {32'hc47ef06c, 32'hc2568bf6, 32'hc204d974},
  {32'hc28650fe, 32'hc328bdb8, 32'hc37acbe4},
  {32'hc49b87ac, 32'h42c3445e, 32'hc3eaf87a},
  {32'h4389f230, 32'h43c69acb, 32'hc30f3053},
  {32'hc35cfd60, 32'hc2ad3758, 32'hc33a1fa4},
  {32'h44094842, 32'hc1d37a10, 32'h42f8aa41},
  {32'hc459f244, 32'hc19319c2, 32'h41e0db39},
  {32'h44380f66, 32'hc3cf542b, 32'h440e10ea},
  {32'hc432e5d0, 32'hc2bd9ad8, 32'h43c46554},
  {32'h43d4fe3a, 32'h41e31362, 32'hc2f470bc},
  {32'hc4b2551f, 32'h42547c2c, 32'h433ff0cc},
  {32'h44b6f062, 32'h42de5965, 32'h41ee3050},
  {32'hc2d6cb20, 32'h42d7fae5, 32'h42412e60},
  {32'h442449f8, 32'h437a2346, 32'h436be85c},
  {32'hc4dbd9f8, 32'hc27d545a, 32'h42e1b336},
  {32'h4490a750, 32'hc3b513ed, 32'h43929ef9},
  {32'hc5116d26, 32'h429a8efd, 32'hc31924e2},
  {32'h4443a410, 32'hc3aa44dd, 32'h42d5633e},
  {32'hc517d1a6, 32'hc33e7ec8, 32'h43eefd8c},
  {32'h43920bf0, 32'hc2ec599b, 32'hc322d215},
  {32'hc4c8f8c4, 32'hc2265531, 32'hc39292c5},
  {32'h450e53a0, 32'h4412cf9b, 32'hc31fc62f},
  {32'hc46fe09e, 32'hc32e9d6a, 32'h4341cf7e},
  {32'h43d7e690, 32'hc2cb4a29, 32'h43f8de95},
  {32'hc50b0a1b, 32'hc28fe146, 32'hc3957563},
  {32'h43e19ff1, 32'hc2ed60c6, 32'hc05ab79e},
  {32'hc4424e70, 32'h4371adbd, 32'h439b39d0},
  {32'h4472e15a, 32'h434be5ad, 32'h438011eb},
  {32'hc4dd26b1, 32'h42be4cdc, 32'h42940245},
  {32'h45181928, 32'h434319d9, 32'h436c3162},
  {32'hc49fddfa, 32'hc31454c7, 32'hc2876a54},
  {32'h4435fe33, 32'hc190cbd5, 32'hc3895562},
  {32'hc31361f0, 32'hc346ff91, 32'hc2c0158e},
  {32'h42a5cca8, 32'h42b0e6e8, 32'h42fb57a9},
  {32'hc411b97f, 32'h41c38603, 32'h4336b342},
  {32'h44d7b549, 32'h4245b911, 32'h42ad661c},
  {32'hc3e97378, 32'hc28dd315, 32'hc2b079b9},
  {32'h444f0847, 32'hc32f63b5, 32'h4330af42},
  {32'hc4b71e5c, 32'hc386d177, 32'hc37d0bef},
  {32'h44f84450, 32'h42babe41, 32'h433ff721},
  {32'hc4354325, 32'hc29fa9ef, 32'h4370c701},
  {32'h44450c33, 32'hc3826849, 32'h42cf3cb1},
  {32'hc43944bd, 32'hc3712d0b, 32'hc394fbcf},
  {32'h44f2bcc1, 32'hc2d81fcf, 32'hc30c7c1b},
  {32'hc4443a62, 32'hc38ed9f7, 32'h439eb16c},
  {32'h4505a815, 32'hc204c3ac, 32'h419477aa},
  {32'hc48407e0, 32'hc274a263, 32'hc3359c80},
  {32'h45133c23, 32'hc3f69632, 32'h4432914d},
  {32'hc44de6c6, 32'h40b34a30, 32'h42f0663c},
  {32'h442ca1e0, 32'h413a300f, 32'h437c4b92},
  {32'hc47ee258, 32'h42d0e5ce, 32'hc35d4e6d},
  {32'h42b86228, 32'hc2c0622f, 32'hc3f24b42},
  {32'hc4fb993e, 32'hc3954509, 32'h43461429},
  {32'h44b05e77, 32'h439dda28, 32'h43b883a4},
  {32'hc1141616, 32'hc32b5c5e, 32'hc1551364},
  {32'h40d670c0, 32'h430ff525, 32'h43e47150},
  {32'hc5141dc9, 32'hc425e301, 32'h44128141},
  {32'h449d8706, 32'h43c37ba7, 32'hc3899eb2},
  {32'hc4ec0b29, 32'hc37dca36, 32'h428569fe},
  {32'h4481a6c1, 32'h4299c472, 32'hc31539e4},
  {32'hc4848a7d, 32'hc2abd761, 32'h436556b0},
  {32'h45009edd, 32'hc3071715, 32'hc30cda90},
  {32'hc4f831cf, 32'hc15727f0, 32'hc29ce155},
  {32'h44b75374, 32'h43d7a01c, 32'hc1eea95e},
  {32'hc516ce1a, 32'h4188633f, 32'h4390e601},
  {32'h44c00938, 32'hc2c51ae0, 32'hc2b752fc},
  {32'hc41c4c13, 32'h437f22b4, 32'h41cea82d},
  {32'h44f268db, 32'hc3c0f59f, 32'hc1b8410c},
  {32'hc48cee9c, 32'h42807016, 32'hc3153024},
  {32'h450b4362, 32'h42f7b3b4, 32'hc2807aa1},
  {32'hc4f75b11, 32'h43064211, 32'h42863558},
  {32'h45015978, 32'h42ab0375, 32'h43b68225},
  {32'hc487c1f6, 32'h4355ad19, 32'h42e2d6f2},
  {32'h44d2542e, 32'h4399e159, 32'hc1e1179b},
  {32'hc41fbacd, 32'hc34214b7, 32'h41f78394},
  {32'h447115d3, 32'hc38fc9ed, 32'h4341f550},
  {32'hc4e9e534, 32'h431403fc, 32'hc348fb6b},
  {32'h4513d7e9, 32'hc2ce5ffe, 32'h43c43fcc},
  {32'hc452e687, 32'hc28fb153, 32'h4371be66},
  {32'h4505c12b, 32'h42bc34ba, 32'h43d00f77},
  {32'hc49ae5cc, 32'h431f17ba, 32'hc3576231},
  {32'h45105552, 32'h4321feb5, 32'hc3c2e16c},
  {32'hc4f2ee30, 32'h43511eda, 32'hc31ea89d},
  {32'h448c3987, 32'hc3701c6a, 32'hc29c639e},
  {32'hc518a4a9, 32'h431be94f, 32'hc22b16f8},
  {32'h44aebf8c, 32'h4399c8a5, 32'h42c465b3},
  {32'hc451beea, 32'hc316842f, 32'h43ac9293},
  {32'h44cdc3ac, 32'h43765127, 32'h4312a05f},
  {32'hc5031253, 32'hc2b64805, 32'hc12dc86e},
  {32'hc2994998, 32'h429badfe, 32'h428e4b9b},
  {32'hc4325b29, 32'h40a3a50f, 32'hc2c0e68e},
  {32'h444c2fc8, 32'h43175888, 32'hc3dbe5dd},
  {32'h426661e0, 32'h42bd95bf, 32'hc1ff7f78},
  {32'h45096d80, 32'h42905594, 32'hbfc2dae0},
  {32'hc4b1207c, 32'hc39715fe, 32'h43d45a40},
  {32'h4411b484, 32'hc248b2dd, 32'h4295868e},
  {32'hc4c77704, 32'hc3079a67, 32'hc2f55d38},
  {32'h44dabc2d, 32'hc3048bb4, 32'hc40b3b5b},
  {32'hc50832e7, 32'hc3a5f5ca, 32'hc19e6f13},
  {32'h4421277a, 32'hc3976798, 32'hc265d0b6},
  {32'hc4d12245, 32'h42d81022, 32'h3f43fda8},
  {32'h44feef5f, 32'h43ea5801, 32'hc3522265},
  {32'hc4b7f429, 32'h43502cbf, 32'h438b64ee},
  {32'h444d5734, 32'h43885096, 32'h4383b926},
  {32'hc4ff9634, 32'h4158ef9c, 32'h41a19db6},
  {32'hc312c6f8, 32'h412fe5a6, 32'h4356d9d1},
  {32'h42beee6a, 32'h42090b33, 32'hc3fd72b0},
  {32'h4449a8d9, 32'hc30ea94f, 32'h42bba5ca},
  {32'hc4d55cc8, 32'h432eb885, 32'hc320b100},
  {32'h44b487e4, 32'hc2f395ed, 32'h43fd2fbd},
  {32'hc4b06df5, 32'hbf2006d8, 32'h42a72c04},
  {32'h44fddc1a, 32'h42ef3e50, 32'h42aff8c5},
  {32'hc4e7280b, 32'h43aede95, 32'h3f653bb6},
  {32'h4457782f, 32'h4261d770, 32'hc3d0df57},
  {32'hc50181d8, 32'h430de3d1, 32'hc30ff311},
  {32'h44fa4b37, 32'h4339c36e, 32'h43112c57},
  {32'hc5025830, 32'hc3c5b0d3, 32'hc2693eb5},
  {32'h44bf9e84, 32'h42865061, 32'h4407218c},
  {32'hc4ec8cfc, 32'h42a430cd, 32'h43be2f5a},
  {32'h43a8c040, 32'h4293bfb2, 32'h43054237},
  {32'hc50302bd, 32'hc22f93eb, 32'hc2abb384},
  {32'h44f54c4e, 32'h43ac7cd7, 32'hc242335e},
  {32'hc41452bc, 32'h42aff2bc, 32'h43862d56},
  {32'h44072146, 32'hc20cbcc9, 32'h41d82c7d},
  {32'hc503dbde, 32'hc406bb7a, 32'h41e7728a},
  {32'h444fd6df, 32'h42951896, 32'h43195221},
  {32'hc3c600b8, 32'h430b31ad, 32'h4347a877},
  {32'h44ea6085, 32'h42d3dbd3, 32'h439c8b18},
  {32'hc519279d, 32'hc3849206, 32'h43ade41c},
  {32'h448bbb3a, 32'hc301ad56, 32'h430ddb06},
  {32'hc3d5154a, 32'hc30232bc, 32'h43c6679a},
  {32'h44ec08e8, 32'h435992a5, 32'h4363914b},
  {32'hc4e98874, 32'h44253ed9, 32'h43722283},
  {32'h44b4802a, 32'hc3894821, 32'hc302e362},
  {32'hc4e35ab0, 32'hc1c8ee39, 32'h411c38a7},
  {32'h44c74d7a, 32'hc375136f, 32'hc0a46f20},
  {32'hc3dc405c, 32'hc395c59d, 32'hc2803f87},
  {32'h44d74aff, 32'hc2954135, 32'h412bfd8f},
  {32'hc4f34e31, 32'h432c1f26, 32'hc2d03be0},
  {32'h4514bbef, 32'h43a67c50, 32'hc36ba0fd},
  {32'hc51411aa, 32'h41b77e46, 32'h4261656d},
  {32'h43bfd3ed, 32'hc314e98d, 32'h4208c707},
  {32'hc4462b30, 32'hc2c9dba9, 32'hc2a01d98},
  {32'h44079292, 32'hc3baede1, 32'hc29b40c9},
  {32'hc4dd546f, 32'h425ef101, 32'hc2f66746},
  {32'hc31812f8, 32'hc162b8ef, 32'h43a50fbd},
  {32'hc4882d28, 32'hc39a8fec, 32'h436efbad},
  {32'h44365edc, 32'hc36590db, 32'h439e9a32},
  {32'hc3e1d98c, 32'h431fbf91, 32'h43c5f149},
  {32'h450912d8, 32'hc328f0c0, 32'h42ca547f},
  {32'h422e8d9c, 32'hc2bf9596, 32'hc3164010},
  {32'h44d44bfe, 32'h4282eb88, 32'hc2b989fb},
  {32'hc428480b, 32'h4268c2a5, 32'h42d2dc91},
  {32'h4290f140, 32'h43ff7868, 32'h43d7d74c},
  {32'hc4aaf327, 32'hc2f8ef06, 32'hc3bb9c11},
  {32'h43ab91dc, 32'hc31ed21e, 32'h42d34086},
  {32'hc4feec01, 32'hc2f8601a, 32'hc35569fe},
  {32'h44b0122d, 32'h4336f05b, 32'hc35fbda7},
  {32'hc51287ef, 32'hc2ca6784, 32'h42e0977b},
  {32'h44deb4f6, 32'h43b416c7, 32'hc28ee834},
  {32'hc500326e, 32'hc23938fd, 32'h43735a05},
  {32'h44e42ce1, 32'h4218c1a4, 32'hc2a22300},
  {32'hc3bcecb4, 32'hc360ffd5, 32'hc2db63fc},
  {32'h44c30da4, 32'hc2676ca9, 32'h41290b44},
  {32'hc4852998, 32'hc3187665, 32'h42d0b039},
  {32'h45152fb8, 32'h435801b5, 32'hc387e13e},
  {32'hc44082ae, 32'h43814f90, 32'h428f1e6b},
  {32'h451442bb, 32'hc2f6c799, 32'hc2a0a373},
  {32'hc4f77b51, 32'hc2dcef7d, 32'hc23418ec},
  {32'h44e30845, 32'hc3c0ff3e, 32'hc2584a10},
  {32'hc435b3e0, 32'h4274dbce, 32'hc3114487},
  {32'h450e7cc9, 32'hc26b11e9, 32'h43093750},
  {32'hc528355f, 32'hc33003d6, 32'h4340540c},
  {32'h44d4971a, 32'hc401f71e, 32'hc203529d},
  {32'hc4b69b86, 32'h43bae9ef, 32'h434c6beb},
  {32'h44ebfc56, 32'h432ad44b, 32'hc37443bf},
  {32'hc395e837, 32'hc31fe73c, 32'h429dfee8},
  {32'h45091935, 32'h438a648f, 32'hc3420afa},
  {32'h415a1e20, 32'hc3687ce6, 32'h3e7a83b0},
  {32'h44ce8844, 32'hc0fba898, 32'hc41eb584},
  {32'hc4ae7d3b, 32'hc34c2a8c, 32'h42715f9a},
  {32'h4286fd60, 32'hc2ad98ce, 32'hc38e9aee},
  {32'hc4e8d0a0, 32'h435e610d, 32'hc35b393f},
  {32'h44aec870, 32'hc2d435d0, 32'hc2eb2dee},
  {32'hc30c55e5, 32'hc35b16e8, 32'h42b89bd6},
  {32'h43d50634, 32'hc39664e9, 32'h43986a88},
  {32'hc2e50fc8, 32'hc394afb3, 32'hc2e7a7c7},
  {32'h448f35b6, 32'h43f26df4, 32'h4375aa8a},
  {32'hc44d559c, 32'h42c456d8, 32'hc3a539e2},
  {32'h42785b70, 32'h42abd305, 32'hc1187719},
  {32'hc509750b, 32'h41e407e9, 32'h4232990a},
  {32'h4404400c, 32'hc239018b, 32'hc341d667},
  {32'hc49cf9e8, 32'h436583bc, 32'hc3829568},
  {32'h446f5657, 32'h42c67a7f, 32'h4386955d},
  {32'hc426a6ec, 32'h42462c12, 32'hc380ce07},
  {32'hc325bd06, 32'h436bff68, 32'h43b2b2bd},
  {32'hc4a7e1f4, 32'h428fbc24, 32'hc30a8e5e},
  {32'h44837344, 32'h4416906d, 32'h430d5232},
  {32'hc4a624b5, 32'h43dc0a72, 32'h43f98585},
  {32'h44baa937, 32'hc332c121, 32'hc3013df4},
  {32'hc3e471e8, 32'h41f0d7be, 32'hc32ab33a},
  {32'h44277c5c, 32'hc1aeba60, 32'hc3bb9120},
  {32'hc51081a5, 32'h429ca17f, 32'hc2e547fd},
  {32'h449b7595, 32'hc382a8fe, 32'hc3d6795f},
  {32'h42372980, 32'h43934c12, 32'h4371be0e},
  {32'h43dccc1c, 32'h4426cd86, 32'hc1c7ba7a},
  {32'hc3870eb4, 32'hc212c9d3, 32'h42b04152},
  {32'h4465d9dc, 32'h42a1e079, 32'hc1558b68},
  {32'hc49620b0, 32'h40a9ab19, 32'hc403b10f},
  {32'h44a24f7e, 32'h4217de78, 32'hbfe42a32},
  {32'hc4a086d4, 32'h42c73a7a, 32'h433b71d1},
  {32'h44911eb0, 32'hc31768b8, 32'hc347dea8},
  {32'hc4fbabca, 32'hc31fbadb, 32'hc3991ab4},
  {32'hc253b980, 32'h42b7d40b, 32'hc27059be},
  {32'hc407049c, 32'hc1edb951, 32'hc35b294c},
  {32'h44bb0f9e, 32'hc268f9aa, 32'h410c3db1},
  {32'h41824330, 32'hc34d7d2a, 32'hc3536f28},
  {32'h44806bf8, 32'hc40ee6d6, 32'hc3045577},
  {32'hc50aefd2, 32'hc30d4f2f, 32'h438ee6c4},
  {32'h44d603f4, 32'hc3209726, 32'h43602238},
  {32'hc4f37579, 32'h431d8ff7, 32'hc30e2805},
  {32'h44e52d7b, 32'h430ada26, 32'hc347480e},
  {32'hc508c280, 32'h437bef32, 32'h42b41123},
  {32'h44115361, 32'h4322199f, 32'h42666029},
  {32'hc4ef80d3, 32'h42dca58e, 32'h4385f8fd},
  {32'hc1d9e500, 32'h421d2437, 32'hc38a4f95},
  {32'hc50e9fc7, 32'hc21f79c4, 32'h42d3eaae},
  {32'h441d0e2a, 32'h438c28d8, 32'hc32958ec},
  {32'hc502c4ac, 32'h4305086b, 32'h40dd011d},
  {32'h44e73c57, 32'h425ec0d0, 32'hc2854272},
  {32'h433214c8, 32'hc1578243, 32'h4361da98},
  {32'h43e4660d, 32'h43e0f1b8, 32'hc2d2dbb8},
  {32'hc50e80b1, 32'hc3ae90f4, 32'h3fecb01a},
  {32'h44d56934, 32'hc135bac4, 32'hc358cfc0},
  {32'hc4ffb0a7, 32'h4322a357, 32'h42a3a1fc},
  {32'h435059e8, 32'h420f5242, 32'hc3016c8a},
  {32'hc5004e7f, 32'h43a42581, 32'h430678c1},
  {32'h444e5941, 32'h4325d3d5, 32'hc2db42f8},
  {32'hc4f53e04, 32'h430efb18, 32'h4224738f},
  {32'h44949273, 32'h4385b5a5, 32'h43aa5b36},
  {32'hc48dd647, 32'hc3613b9d, 32'h433f60f7},
  {32'h44ccbc90, 32'hc37f8ec2, 32'h4382606a},
  {32'hc4d69481, 32'hc2f0a46d, 32'h439c7f3e},
  {32'h43e58eef, 32'hc316b78c, 32'hc36ec75e},
  {32'hc434309c, 32'hc290ea13, 32'h428d09a5},
  {32'h440cd199, 32'h42b628bf, 32'hc3787104},
  {32'hc4cdd958, 32'h4241cb67, 32'h43704c5b},
  {32'h44bfae05, 32'h43141374, 32'h43216bd9},
  {32'hc4ac9264, 32'h42323947, 32'hc33d65bc},
  {32'h44eee48a, 32'h4323c098, 32'h420d79c2},
  {32'hc50a3054, 32'hc366b55f, 32'hc3764c1b},
  {32'h443bdf95, 32'hc3b06274, 32'hc35e5eb0},
  {32'hc48d3e94, 32'h42fb1544, 32'h4304c63a},
  {32'h44bbbdfa, 32'hc2cda0ba, 32'hc2b07553},
  {32'hc50423dd, 32'h430247d1, 32'h424db62d},
  {32'hc4bc3474, 32'h42cc4e2c, 32'h431b75e4},
  {32'h41fd4980, 32'hc1f2125a, 32'h42a02556},
  {32'hc42e9f23, 32'h42ab5b13, 32'h433d1dbe},
  {32'h44946609, 32'hc180dcbc, 32'hc2f92469},
  {32'hc3e0213c, 32'h43892838, 32'hc1b23a9e},
  {32'h44f723fa, 32'h435bce45, 32'h42d5ed52},
  {32'hc4c6b3bc, 32'hc3894db4, 32'h43104798},
  {32'h44bfff3e, 32'h436363e3, 32'hc316c10d},
  {32'hc105e0a0, 32'h436406be, 32'h42dd0afd},
  {32'h45167e9d, 32'hc36eca03, 32'hc29f62ab},
  {32'hc461ec77, 32'h432c82bd, 32'h420ccc1d},
  {32'h44e7410f, 32'hc2e7c446, 32'hc26e81a3},
  {32'hc4b82310, 32'hc16b454a, 32'hc3f53aee},
  {32'h448795ff, 32'h42dc38b5, 32'h433e24a5},
  {32'hc51f919a, 32'hc4201566, 32'hc31a713e},
  {32'h42f59490, 32'hc2f2a52b, 32'hc0d0ac84},
  {32'hc3acd3f8, 32'h43371d66, 32'hc1fc5a1d},
  {32'h43ee2118, 32'hc1878055, 32'h42ed2bff},
  {32'hc4f3ae13, 32'h42cbe02b, 32'h428d3619},
  {32'h444eeab0, 32'h41f98a6f, 32'hc3826dd2},
  {32'hc4f8171e, 32'hc37d4e3e, 32'h439583ae},
  {32'h44d485e0, 32'hc3edec5f, 32'hc2839749},
  {32'hc431ce08, 32'hc3bf3b11, 32'h41e799f9},
  {32'h44ded457, 32'h43140abe, 32'hc3592be1},
  {32'hc465885e, 32'hc35294c3, 32'h438c31bf},
  {32'h450fea06, 32'hc30dcaf1, 32'h430d84de},
  {32'hc41c58d8, 32'hc3d5293c, 32'h42d10cae},
  {32'h43141840, 32'h432fe3f6, 32'h434afdc2},
  {32'hc4f59f06, 32'hc3335337, 32'hc1f39302},
  {32'h43c3f6cf, 32'h432b4000, 32'hc30e981b},
  {32'hc4caa12f, 32'hc331a431, 32'h42aeb846},
  {32'h44b17685, 32'hc2af2045, 32'h431faec1},
  {32'hc49d63be, 32'hc188f7cc, 32'hc241d41c},
  {32'h44595b44, 32'h431a3c26, 32'h43a23407},
  {32'hc51317e5, 32'hc382c898, 32'h432859e6},
  {32'h450f7bcf, 32'hc3c825b5, 32'hc38ec6ea},
  {32'hc40bc549, 32'h43ad0917, 32'hc37037b1},
  {32'h447352bf, 32'h43bdc5df, 32'hc29e9d4f},
  {32'hc4a211dd, 32'h43c4d1db, 32'hc3236b7b},
  {32'h450663cd, 32'hc2aa687a, 32'h434246e7},
  {32'hc4bb7b40, 32'h43120eb2, 32'h4307d30b},
  {32'h446269c3, 32'h42954b36, 32'h43e0bf01},
  {32'hc517a708, 32'hc289ba0c, 32'hc2ba34ff},
  {32'h4506e6fd, 32'h42a60002, 32'hc3422a25},
  {32'hc41d8247, 32'h431d2f37, 32'hc2dd1b9f},
  {32'h44cfd01e, 32'hc12d41f0, 32'h434d5e48},
  {32'hc36ad468, 32'h4082608f, 32'h43accc66},
  {32'h44bc4595, 32'hc3a262f2, 32'h43b249c9},
  {32'h41633f00, 32'hc2b52a17, 32'h43f01a0f},
  {32'h4496b48d, 32'h43cbfd9d, 32'hc30f72c8},
  {32'hc50862b9, 32'h42a29452, 32'h41831302},
  {32'h4286e770, 32'hc3a611ea, 32'hc233f345},
  {32'hc5168233, 32'h430419fc, 32'hc3317945},
  {32'h44b99ead, 32'hc3d159c3, 32'h43302919},
  {32'hc511664b, 32'hc2fe0ed2, 32'h4356be73},
  {32'h44d0af60, 32'hc30b38a7, 32'h436ca500},
  {32'hc4d95299, 32'hc24d8da3, 32'hc3d43345},
  {32'h44ab2769, 32'hc2020235, 32'hc2693223},
  {32'hc40abee2, 32'hc316bf62, 32'h42ac8c9c},
  {32'h4462165d, 32'hc3019eba, 32'hc283d648},
  {32'hc4e7e54b, 32'hc39085a4, 32'hc41270bd},
  {32'h450657ba, 32'h433858b5, 32'hc3769384},
  {32'hc4484ed0, 32'hc34419b6, 32'h4393a76d},
  {32'h448780da, 32'h41aa2669, 32'h4383d448},
  {32'hc42dc1d4, 32'hc2f5765a, 32'h422e179a},
  {32'h444c45b0, 32'hc37939ec, 32'h43308347},
  {32'hc48be7be, 32'h43071480, 32'hc3ae4399},
  {32'h44cb989c, 32'h4314a416, 32'h41f61881},
  {32'hc50f1ce6, 32'h41fdd7ad, 32'hc3898768},
  {32'h44cb47c6, 32'hc303d838, 32'hc2ed3450},
  {32'hc520fea6, 32'h42bdd3a4, 32'h41f7b364},
  {32'h44153927, 32'hc3a4ca71, 32'h4406a550},
  {32'hc3136110, 32'h43992974, 32'hc302ccba},
  {32'h435d9de0, 32'h429e4b96, 32'h438b7133},
  {32'hc3f6516f, 32'h4225c06f, 32'hc30bc51f},
  {32'h4504deca, 32'h43791417, 32'hc1c00edf},
  {32'hc4b0e5a6, 32'h41e90de6, 32'hc3a43270},
  {32'h448a05c9, 32'h42fc2548, 32'hc3bc596b},
  {32'hc41c2390, 32'hc3402b95, 32'hc2180a17},
  {32'h44b00265, 32'hc2965ced, 32'hc304e287},
  {32'hc48c98ac, 32'h428dffe0, 32'h4339cf23},
  {32'h43db1178, 32'h43b95be9, 32'h43a588e7},
  {32'hc4b38dc2, 32'hc104a16e, 32'h42935740},
  {32'h43c4b489, 32'h42d38374, 32'hc36dac10},
  {32'hc4bef9df, 32'hc2d51a77, 32'h43a1cf32},
  {32'h43a0a4d0, 32'h432edc1f, 32'hc2bb4196},
  {32'hc5046605, 32'h410bdbfa, 32'hc31cec30},
  {32'h45180948, 32'hc341fded, 32'hc3b6b608},
  {32'hc4ca2a68, 32'hc370fcda, 32'hc2b45c5c},
  {32'h4402424c, 32'h4338fded, 32'h419fd55f},
  {32'hc4f5908b, 32'hc356c5e8, 32'hc35e6dca},
  {32'h4479f7d8, 32'h433a69df, 32'h438951e0},
  {32'hc337f618, 32'h42a18e50, 32'h424decb6},
  {32'h44dcc62c, 32'hc3d2bcc6, 32'h426656ab},
  {32'hc4c61db8, 32'hc1d7682a, 32'h42a09e97},
  {32'h42ae7278, 32'hc35bff8b, 32'h42a1b1a2},
  {32'hc1cece1c, 32'hc1ba0461, 32'hc38aca43},
  {32'hc3a257dc, 32'hc3dc2fcb, 32'hc2a2669f},
  {32'hc4cf32ee, 32'hc189cded, 32'h433220e7},
  {32'h4474f04c, 32'h42f3cb79, 32'h43078542},
  {32'hc4cce552, 32'hc34773ed, 32'hc405a8a1},
  {32'h44f48c2f, 32'h432fcb00, 32'hc38ecca6},
  {32'hc4d4bdc1, 32'h435e9580, 32'hc2810f04},
  {32'hc4b88724, 32'hc218bf16, 32'hc37a3902},
  {32'h44d619cd, 32'hc223d000, 32'hc31175cc},
  {32'hc44a9440, 32'hc206abb5, 32'hc1002dcd},
  {32'h4504e402, 32'hc14893f1, 32'h43896758},
  {32'hc4db6e66, 32'h421c07b0, 32'hc3c56238},
  {32'h44839437, 32'h433349a1, 32'h43d113c7},
  {32'hc4711fec, 32'h432a17b3, 32'hc36a0210},
  {32'h44a041e8, 32'h42c37142, 32'h421e2bc5},
  {32'hc485b91e, 32'hc363eab3, 32'h40fb11d0},
  {32'h44e95d58, 32'hc34d829e, 32'h41b1ca9c},
  {32'hc4bec639, 32'h43a3d744, 32'hc285e65f},
  {32'h451c6d5d, 32'hc2889022, 32'hc2a5d4c5},
  {32'hc4df169f, 32'hc3fa398e, 32'hc2e28f1e},
  {32'h4502ce7a, 32'h43c37ff0, 32'hc384957c},
  {32'hc4939994, 32'hc1bc9944, 32'h4391713d},
  {32'h450eb940, 32'hc23fe23a, 32'h432a0bf8},
  {32'hc2f47f70, 32'hc23d2811, 32'hc35a0a18},
  {32'h4415625a, 32'hc3743ffa, 32'h435a04c8},
  {32'h43b120bc, 32'hc36a42ab, 32'hc383d9aa},
  {32'h44c95760, 32'h42abf934, 32'h42b1a367},
  {32'hc50ee001, 32'hc2e6d07e, 32'h42e2992e},
  {32'h449b0799, 32'h415967de, 32'h430e53ce},
  {32'hc305c6e4, 32'hc2b0ea97, 32'hc35c1960},
  {32'h438edd40, 32'hc2dd1273, 32'h42caa284},
  {32'hc4408d2f, 32'h431f0f2d, 32'h406f3d71},
  {32'h450282a5, 32'h40e011d1, 32'hc34c88e7},
  {32'hc471d37e, 32'h431485f3, 32'h4262fda7},
  {32'h44336a06, 32'hc3b81015, 32'h43a0b55d},
  {32'hc500d406, 32'hc0b51ce0, 32'hc38a5043},
  {32'h446d1470, 32'h438c23ea, 32'hc2e3412a},
  {32'hc484db9f, 32'hc27e995b, 32'hc391d96e},
  {32'h44db3db5, 32'h4396d447, 32'h43d1776e},
  {32'hc401dd7c, 32'h434eb59c, 32'hc29aafa0},
  {32'h44306d2a, 32'hc3565817, 32'h42c29230},
  {32'hc4958791, 32'hc38f761b, 32'hc388dd78},
  {32'h44dddfaf, 32'h41d6dd65, 32'hc3884b39},
  {32'hc4203381, 32'h4111d746, 32'h4107f903},
  {32'h4492339b, 32'hc38a3fed, 32'h43db4b83},
  {32'hc4e794c2, 32'h42ba4927, 32'hc22212bc},
  {32'h4502108b, 32'hc394a06d, 32'h42a0c737},
  {32'hc4c1ed04, 32'h413c910e, 32'h437d79b4},
  {32'h44a6d053, 32'hc3ee2735, 32'h440adbf7},
  {32'hc41e75b0, 32'h431dee5b, 32'h43779172},
  {32'h43c1ca5e, 32'h431ec7e8, 32'h430fbd4c},
  {32'hc5147d1e, 32'h43a9685d, 32'h42ac92f0},
  {32'h44c55488, 32'hc36cfe9a, 32'hc34ebbea},
  {32'hc460d3a0, 32'hc3877fea, 32'h42178f20},
  {32'h44a4fe9a, 32'hc35ff460, 32'h4357a842},
  {32'hc49924ff, 32'hc21a7dcf, 32'h428af86f},
  {32'h4498f6cf, 32'hc19981eb, 32'hc3698563},
  {32'hc4ec8c82, 32'hc2521c27, 32'h42b8fc7d},
  {32'h4512eb36, 32'h43453edb, 32'hc217d13e},
  {32'hc4b0e142, 32'h42c9d2f2, 32'hc2e9cd3d},
  {32'h45245178, 32'h40b51100, 32'h42a5901f},
  {32'hc4e90c46, 32'h439f8784, 32'h420f4701},
  {32'h44d99bb2, 32'h419b7e3b, 32'hc3619667},
  {32'h430d1210, 32'h434b2794, 32'h4375535d},
  {32'h44d38555, 32'h432c88ca, 32'hc3228733},
  {32'hc45564b8, 32'hc27f8d48, 32'hc39ceec6},
  {32'h431c45f6, 32'hc319b239, 32'h4417340d},
  {32'hc4ef3de0, 32'h4318d5f8, 32'h43b1e5bc},
  {32'h44e47bf8, 32'h42ba3f7c, 32'h42b2338b},
  {32'hc314db8e, 32'h40afc370, 32'h43152165},
  {32'h45189bd5, 32'hc3652e43, 32'hc3b91f85},
  {32'hc510a5ad, 32'hc3641467, 32'hc2873516},
  {32'h42b6fb80, 32'hc219408d, 32'h440ee826},
  {32'hc44ef902, 32'h43b14fb1, 32'hc38a6abe},
  {32'hc2bcca00, 32'h41f30615, 32'hc353020a},
  {32'hc329a9c1, 32'h4307503b, 32'hc396690b},
  {32'hc194c6a0, 32'h43774804, 32'hc31da51e},
  {32'hc45a811b, 32'hc3800f0b, 32'hc2a6d6e9},
  {32'h441c2566, 32'hc22328e3, 32'h4395af15},
  {32'hc4d5ffbc, 32'h4106507e, 32'h438e9131},
  {32'h434ece30, 32'h431b65d6, 32'h42e04276},
  {32'hc4b95a74, 32'h430cc811, 32'h43c7cc8d},
  {32'h445fa488, 32'h42b5af4a, 32'h434ccc5c},
  {32'hc4490ec3, 32'hc2c31833, 32'hc33dee4c},
  {32'h43f1159c, 32'h407d0a30, 32'hc073c65c},
  {32'hc524574a, 32'h429412e6, 32'h41f5cdb4},
  {32'h43bc6e3c, 32'hc39139df, 32'h43b2ffe7},
  {32'hc1223d00, 32'hc2bea21e, 32'hc1a22f4c},
  {32'h447e7566, 32'hc419611f, 32'h4328215f},
  {32'hc4bd8dda, 32'h43af7f9a, 32'hc37508dd},
  {32'h4488192e, 32'hc3c85a31, 32'h4186a960},
  {32'hc4a370d0, 32'h40fa4946, 32'hc284d8ff},
  {32'h45142ae4, 32'h419ac778, 32'hc2b02809},
  {32'hc41b7800, 32'h41b68882, 32'hc390926b},
  {32'h451098b3, 32'hc34613cb, 32'h43209f1b},
  {32'hc43c077a, 32'hc3030c6f, 32'h44002f05},
  {32'h44eb4ebb, 32'h413b20d9, 32'hc3a5ca2f},
  {32'hc430a20c, 32'h43120340, 32'h42935a40},
  {32'h44355a54, 32'h4336db80, 32'h421ee130},
  {32'hc4c7bdb0, 32'h42d933ff, 32'h4399f459},
  {32'h439381b6, 32'h422bb26d, 32'hc381eead},
  {32'hc3ccee74, 32'hc303e427, 32'h42f08e5e},
  {32'h4414d142, 32'hc3ae595b, 32'h433e63ab},
  {32'hc50dca1a, 32'hc0e42489, 32'hc336402b},
  {32'h440bf3da, 32'hc3594a99, 32'hc361e894},
  {32'hc490f553, 32'hc310c734, 32'h4340c413},
  {32'h4339f490, 32'h425169b8, 32'h43017b78},
  {32'hc40adc02, 32'h4323763a, 32'h4162f7de},
  {32'h449ef61a, 32'hc2153c7a, 32'h438f2942},
  {32'hc34ed326, 32'hc37d2b02, 32'hc35c622b},
  {32'h4431d8c2, 32'hc2b5b08a, 32'hc41173c4},
  {32'hc4198bc7, 32'h43f03a03, 32'h43591eb3},
  {32'h4464246c, 32'h4284a55b, 32'hc305600b},
  {32'hc4538bc0, 32'hc22dc29f, 32'h40660926},
  {32'h4454a381, 32'h42a1f3be, 32'hc40ab906},
  {32'h42b3bb12, 32'h435e230e, 32'h4196f3f8},
  {32'h44308912, 32'h4394589b, 32'h42bd6bae},
  {32'hc4d5f4d0, 32'h4325fc2a, 32'h4363d576},
  {32'h445e19df, 32'h434d6489, 32'hc3d4cbc1},
  {32'hc34ee500, 32'h43a9034a, 32'hc1f77e03},
  {32'h4513bc0d, 32'hc31c6300, 32'hc38430cd},
  {32'hc45e5270, 32'h42821ee4, 32'h43e22bda},
  {32'h443338de, 32'h4169f30f, 32'hc3c484e3},
  {32'hc415be08, 32'h431abbc4, 32'hc3f055c3},
  {32'h44c769e6, 32'h43471f96, 32'h43489062},
  {32'hc4ebfb84, 32'h40fb6f1a, 32'h42b895ee},
  {32'h4417f290, 32'hc39f121e, 32'h430ddb55},
  {32'hc4ab31af, 32'h405bc460, 32'hc291569d},
  {32'h44c355fd, 32'hc3a08e19, 32'hc369ea82},
  {32'h43232a9c, 32'h42c56269, 32'h436eceb4},
  {32'h43c44084, 32'hc27ebf65, 32'h43597f90},
  {32'hc48cee26, 32'hc3a5af8f, 32'hc33045e5},
  {32'h44ebf950, 32'h42b1a670, 32'h431a0e10},
  {32'hc44f0404, 32'hc08019d8, 32'h430a4b84},
  {32'h4501a932, 32'hc1f992cf, 32'h4201e01b},
  {32'hc4478bdb, 32'h42a146c2, 32'h43848097},
  {32'h44510afe, 32'h433b90af, 32'hc324ab31},
  {32'hc4ffa710, 32'hc10bf6de, 32'hc3921b9f},
  {32'h44adec67, 32'hc303b40e, 32'h42c34135},
  {32'hc49930ca, 32'h43866db3, 32'h4396b32e},
  {32'h45141c53, 32'hc33e7a2c, 32'hc2d62cda},
  {32'h43b68dce, 32'hc2c52152, 32'hc4133874},
  {32'h44a3ab8e, 32'h426df617, 32'h42a48b70},
  {32'hc30d47d7, 32'h433e3b2c, 32'h43ca8cde},
  {32'h4502a840, 32'h42dd7a5e, 32'hc1b5933b},
  {32'h420f3060, 32'h4405904e, 32'h42998e52},
  {32'h450289ec, 32'hc40ec18c, 32'hbf41bdf8},
  {32'hc4e4fb51, 32'h42ab00c3, 32'h40e2f8c8},
  {32'h43db5670, 32'hc31e5a12, 32'h42a5ef1b},
  {32'hc36b8680, 32'hc1ea4b0a, 32'h43890fe6},
  {32'h44b2615e, 32'hc326eb74, 32'h41e84ef5},
  {32'hc471936c, 32'hc36b3538, 32'h433c6579},
  {32'h450241ce, 32'hc3f25098, 32'hc2b198ad},
  {32'hc4c61a7a, 32'h406f009b, 32'h4332732b},
  {32'h441457a2, 32'h43cd8e7f, 32'hc392d4f6},
  {32'hc499ffb7, 32'hc340b950, 32'h435f5e25},
  {32'h450705bf, 32'hc1a143ad, 32'h4301ceb2},
  {32'hc387f6b8, 32'hc3f5b5a8, 32'hc3b58fcc},
  {32'h446d7e16, 32'h43f0684d, 32'h43ce9ad7},
  {32'h410daaf6, 32'hc25bd30f, 32'hc29d195e},
  {32'h44e59ff6, 32'h423e5df6, 32'hc343f391},
  {32'hc3bea98c, 32'h43ae3325, 32'h421cf768},
  {32'h443a411e, 32'h42b0c712, 32'hc31cbadc},
  {32'hc48026dc, 32'hc30d4346, 32'hc366d212},
  {32'h44e437cf, 32'h43c1bf5e, 32'h435359d1},
  {32'hc394cd8f, 32'h42c33125, 32'hc20fb07b},
  {32'h44310d78, 32'hc24d17b5, 32'h43aaad5e},
  {32'hc3744903, 32'h43f79b30, 32'h41e3a02c},
  {32'h441c7eb5, 32'hc362a995, 32'hc32f3d56},
  {32'hc505eb40, 32'h43513895, 32'hc2c96dc3},
  {32'h450c7056, 32'h43889ad1, 32'h43168011},
  {32'hc4cade53, 32'hc31ece52, 32'hc2a4a494},
  {32'h450cf717, 32'h408324f0, 32'h4329b7e4},
  {32'hc4de623c, 32'h42ec3d7c, 32'hc26f71a1},
  {32'h44f31537, 32'h4404d4fb, 32'h42980582},
  {32'hc480eac2, 32'h434663d4, 32'hc2cabb35},
  {32'h44fe2119, 32'h4296c162, 32'h436a4c94},
  {32'h3e154000, 32'h43b1397e, 32'h4195a329},
  {32'h451ccab6, 32'h43c9475e, 32'h43a45e34},
  {32'hc3d18e12, 32'hc28d0bf8, 32'h4356ec7b},
  {32'h450fa394, 32'h43085f08, 32'h43a16047},
  {32'hc39efbfc, 32'h42efb348, 32'hc2e4bc1a},
  {32'h43c58750, 32'hbfd1af8f, 32'hc2b726e5},
  {32'hc4c0b260, 32'hc0ba9de4, 32'hc3d90f30},
  {32'h44f4fce4, 32'hc2f31e6c, 32'hc3c13b6e},
  {32'hc326d044, 32'hc36f7489, 32'h43b48f1f},
  {32'h43dba7ca, 32'hc32ce2c5, 32'hc3c4b8ad},
  {32'hc4f0d8a1, 32'hc3309ab5, 32'hc1ce115f},
  {32'h44b724d0, 32'h43e0c7e5, 32'h4178502a},
  {32'hc48f0655, 32'hc39950b2, 32'hc39fe583},
  {32'h4439f706, 32'hc266e054, 32'hc3b166b7},
  {32'hc4d19a76, 32'hc30c3875, 32'hc335b59c},
  {32'h45107989, 32'h439f7e21, 32'h4388387a},
  {32'hc4028136, 32'h444cebf1, 32'hc2ec7ea4},
  {32'h44c17250, 32'hc25b1c67, 32'h431cac44},
  {32'hc4f13bba, 32'hc415edae, 32'hc0ecaad6},
  {32'h44e7fa6d, 32'hc32bc512, 32'hc31e0d86},
  {32'hc4b5c55e, 32'h43aecf5e, 32'h4261a379},
  {32'h440fdcee, 32'hc24fb266, 32'h421ca783},
  {32'hc5022e2e, 32'h4373138d, 32'h3fef535c},
  {32'h44b7afc4, 32'hc3e6d64b, 32'h4324765b},
  {32'hc4f9fd6e, 32'h430abf5d, 32'hc26b7f33},
  {32'h43982f73, 32'h43964411, 32'h425aba88},
  {32'hc449f1af, 32'hc25e7aa1, 32'h43293add},
  {32'h44a431ca, 32'h42771ed0, 32'hc3804064},
  {32'h438051d9, 32'hc2fa7d6a, 32'h439281ab},
  {32'h450d084e, 32'h4363be0e, 32'hc279338c},
  {32'hc5019dba, 32'h4372353c, 32'hc36c02d8},
  {32'h450a9993, 32'h4311e154, 32'h43672182},
  {32'hc1713460, 32'hc2ce1e40, 32'hc3180505},
  {32'h449d43f0, 32'h433bfc17, 32'hc3f955c7},
  {32'hc4b01b9d, 32'h3dc39900, 32'h436eb5f2},
  {32'hc308d2b8, 32'hc1c6400e, 32'hc2ab4f10},
  {32'h41627d80, 32'hc3d30821, 32'h42f4bed5},
  {32'h44b3c7f9, 32'hc39842d7, 32'hc3ea2144},
  {32'hc49cbfb4, 32'hc38f0d5a, 32'hc3cdae95},
  {32'h450d85c7, 32'h42dfcb34, 32'hc37aaf90},
  {32'hc4b6d4f2, 32'h434f9164, 32'h4345952b},
  {32'h437aa6a4, 32'hc38666b0, 32'hc3cdcfdb},
  {32'hc3a79d85, 32'hc2c2eefd, 32'hc35a3bfb},
  {32'h44c35f71, 32'hc257d7c1, 32'hc28f09bf},
  {32'hc411c3c4, 32'h42191cc8, 32'h42b58a6e},
  {32'h44c3b901, 32'hc1827364, 32'h43461e0f},
  {32'hc49c42d5, 32'h42aba0d9, 32'hc418e1ff},
  {32'h436029d0, 32'h439dd304, 32'h43d34be8},
  {32'hc29ff8f0, 32'h41949bbd, 32'h432c3c4f},
  {32'h44f38d6f, 32'h430e5f57, 32'h437ae44f},
  {32'hc454f60b, 32'h434514a3, 32'hc327a121},
  {32'h44fc29be, 32'h4327fa2d, 32'h420adb31},
  {32'hc50a6d84, 32'hc2ac4191, 32'hc3a2b246},
  {32'h44d909e2, 32'hc34fc6aa, 32'hc3893321},
  {32'hc447799e, 32'h429e2906, 32'h42f4d821},
  {32'h45082767, 32'hc31be81f, 32'h43825bf7},
  {32'hc4016698, 32'h441ea666, 32'hc3385fa4},
  {32'h43674b70, 32'h43a82a6e, 32'h435fdfbd},
  {32'hc4ded363, 32'h41b89269, 32'h432bdd7b},
  {32'h44238c90, 32'hc30d7dfe, 32'hc3019367},
  {32'hc48e0095, 32'hc3cb87b9, 32'h43862f57},
  {32'h4395686d, 32'hc269c5b4, 32'hc37bbb33},
  {32'hc4f0d43e, 32'h43801296, 32'h424b1424},
  {32'h44220e36, 32'h43331c85, 32'h42d8af12},
  {32'hc437e2f0, 32'hc1bb24c4, 32'h4087aefc},
  {32'h44985e6d, 32'hc36b1f09, 32'h4288a09c},
  {32'hc4fa5632, 32'hc268ad4c, 32'h42d6e055},
  {32'h44eb9d7a, 32'hc22af467, 32'h42d99261},
  {32'hc4accddf, 32'hc373e33e, 32'h43af5b4d},
  {32'h44341032, 32'hc3d43f24, 32'h41ed769d},
  {32'hc50568c7, 32'h43b153a2, 32'h40badffa},
  {32'h44ae2ac8, 32'h43ad10e1, 32'hc2d77140},
  {32'hc434c014, 32'hc2d48968, 32'h4381961d},
  {32'h44fabc6c, 32'hc097124d, 32'h410e291b},
  {32'hc4fcfafe, 32'hc2fb078f, 32'h4306b7fa},
  {32'h439af447, 32'hc31cb5b3, 32'h43736599},
  {32'hc3afe5a0, 32'h43a5b602, 32'hc35ded80},
  {32'h4502bb1e, 32'h43b6f0f8, 32'hc37f45f6},
  {32'hc416765e, 32'hc391f179, 32'hc38b1a5c},
  {32'h44e2b4e7, 32'h42e7b621, 32'h428bcb3f},
  {32'hc49001b7, 32'h441865e2, 32'hc33f14a5},
  {32'h445a85cd, 32'hc2fceea8, 32'h43115d4f},
  {32'hc498137f, 32'h428fe763, 32'hc263b018},
  {32'h451126e8, 32'h429b4131, 32'hc3a6950b},
  {32'hc46941d8, 32'hc202cbd6, 32'hc2c95068},
  {32'h44f96f1c, 32'hc3134171, 32'h42a87a34},
  {32'hc2145c7e, 32'hc11e91a3, 32'h41b14714},
  {32'h44f5fe28, 32'hc1a0452b, 32'h42d3e6c3},
  {32'hc473ae60, 32'h43e698b3, 32'h43710036},
  {32'h44cfc551, 32'h43c27751, 32'h43bd508c},
  {32'hc4bb6a4e, 32'hc3ce5fb3, 32'hc30adb7e},
  {32'h44be9d22, 32'hc2d97e5a, 32'h421681d1},
  {32'hc5045a74, 32'hc21cc135, 32'hc321f768},
  {32'h44b6817f, 32'h431f7e82, 32'hc3ce8ba4},
  {32'hc40ae090, 32'hc2bb3bb5, 32'h43a595b4},
  {32'h44d5c489, 32'hc39cc711, 32'h43854af7},
  {32'hc435cbae, 32'hc1cbf826, 32'hc3b37699},
  {32'h44f6fe70, 32'hc2527184, 32'hc2fa83b3},
  {32'hc42a0aed, 32'h42baaf2b, 32'hc3a2f368},
  {32'h44f6d6f6, 32'hc3bce962, 32'hc3293efc},
  {32'hc4b55d66, 32'hc3197f04, 32'hc2daade4},
  {32'h44ed6c96, 32'hc3420301, 32'h42ab22f0},
  {32'hc0745a00, 32'h436a02fb, 32'hc2f423f8},
  {32'h44b49b78, 32'h43b763c0, 32'hc3afe31a},
  {32'hc3781c2a, 32'hc10d363d, 32'hc24621ba},
  {32'hc0bfee00, 32'hc37431c7, 32'h41ad2824},
  {32'hc3a3d5c8, 32'h41d359e2, 32'h432889e7},
  {32'h4282f350, 32'h4248fdc5, 32'hc09b2156},
  {32'hc51fc741, 32'hc36ff4dd, 32'hc30cc0de},
  {32'h44fc00a9, 32'hc3337340, 32'hc24f2ee1},
  {32'hc35661e0, 32'hc27088ec, 32'h428b5b89},
  {32'h44cfddbf, 32'h422135cc, 32'hc3c158d7},
  {32'hc3b29c2e, 32'h438080d7, 32'h431f71df},
  {32'h42d652d0, 32'hc32bdf2d, 32'h433bc97f},
  {32'hc383a724, 32'h43197fb8, 32'hc3046e79},
  {32'h44f6fa02, 32'hc39e656b, 32'h408ebef6},
  {32'hc502b49e, 32'hc2fb9dcf, 32'hc29a319d},
  {32'hc33aa3f8, 32'h417a8646, 32'h43568410},
  {32'hc4b19e25, 32'h431bfca5, 32'h43ceb20d},
  {32'h4482680b, 32'hc32b5dd2, 32'h4395da1b},
  {32'hc47eecd2, 32'hc205d416, 32'h43207433},
  {32'h44e78a18, 32'h437fc4ad, 32'hc34c8230},
  {32'hc4a405ea, 32'h430f7e0e, 32'hc3cf2757},
  {32'h43a2aa0b, 32'h43ed883a, 32'hc3a8fab6},
  {32'h4127b800, 32'hc2b73bc6, 32'hc37216ee},
  {32'h43b37adc, 32'hc1d97ee1, 32'hc168fc08},
  {32'hc4b84792, 32'h43a1ac74, 32'h4312ac0f},
  {32'h44200da4, 32'h4183a40c, 32'h43423630},
  {32'hc4f9b82e, 32'h4010c2b6, 32'h432923e3},
  {32'h44932bfd, 32'hc30a3f3a, 32'h42abb007},
  {32'hc479ef74, 32'hc2cce1db, 32'hc34d5f62},
  {32'h44a3f0a0, 32'hc1c4b795, 32'h43038550},
  {32'hc4e21606, 32'hc3098605, 32'h434d0daa},
  {32'h43a5030c, 32'hc38ad380, 32'hc34d05bc},
  {32'hc48e3864, 32'hc30b0369, 32'h42ee6dd0},
  {32'h452ae1db, 32'hc3a909d6, 32'hbe463e40},
  {32'hc4b1caca, 32'hc3cd16b3, 32'hc399d7cd},
  {32'h44a24fb7, 32'hc39e2018, 32'h423994b3},
  {32'hc4863997, 32'h41c3a5b6, 32'h41ae1d5d},
  {32'h450e596f, 32'hc282117f, 32'hc3001163},
  {32'h42a6010e, 32'h43259f5b, 32'hc303ba46},
  {32'hc4d5d4c2, 32'hc1c46559, 32'hc347e862},
  {32'h450a1834, 32'hc185ab14, 32'h40dc9fe4},
  {32'hc3acda00, 32'hc350c3b9, 32'hc1a73cfb},
  {32'h453bb0e4, 32'h439f95d0, 32'hc0aa929e},
  {32'hc4591ac9, 32'h43463a76, 32'hc40229da},
  {32'h447648c6, 32'h4348fb81, 32'h42307fa2},
  {32'hc4e2c650, 32'h43196ac2, 32'h43b03f3c},
  {32'hc2a74938, 32'h4346bd2f, 32'hc2c60664},
  {32'hc3b1920c, 32'h4295be76, 32'hc4093ee8},
  {32'h44c6d8cd, 32'hc3df4677, 32'h43d3caca},
  {32'hc4a10034, 32'hc343c415, 32'hc3ff8409},
  {32'h441b52d4, 32'hc3a65c7b, 32'h440017bb},
  {32'hc49dcc92, 32'hc19cfef0, 32'hc2c3ff44},
  {32'h44a6ad34, 32'hc38f258c, 32'h442eafad},
  {32'hc4ef7498, 32'hc3030a8c, 32'h439023c0},
  {32'h44f0a277, 32'hc3a9343d, 32'h428bf951},
  {32'hc507703c, 32'hc3265ceb, 32'h435c3d5c},
  {32'h44c108da, 32'hc380a94d, 32'h43bf4fed},
  {32'hc4b116f6, 32'hc2f3218b, 32'h429e2c6a},
  {32'h43d8b0d2, 32'hc32f9bd0, 32'hc2c1ed39},
  {32'hc41a875c, 32'h42e8594a, 32'h423059fe},
  {32'hc4978d6d, 32'hc355d7d0, 32'hc43ddb30},
  {32'h44558825, 32'hc3968602, 32'hc19564c2},
  {32'hc439bcc4, 32'hc3111b31, 32'hc3c3c68b},
  {32'h44ceea21, 32'hc31f7fd7, 32'hc3260275},
  {32'hc51fa814, 32'h439867e0, 32'hc3ad2851},
  {32'h45035fcf, 32'hc2847b37, 32'h43a04d58},
  {32'hc48f4834, 32'h421b6dec, 32'h43afb969},
  {32'h449a169d, 32'h3eed0d80, 32'h41a5421d},
  {32'hc51afa5f, 32'h428ba6f9, 32'h439c4bda},
  {32'h44e071dd, 32'hc1a0054e, 32'hc2bd62de},
  {32'hc508f0fc, 32'hc2fbb896, 32'hc260d74a},
  {32'h44599ac4, 32'h422918bc, 32'hc39c0a66},
  {32'hc38a45d1, 32'h43bac8ce, 32'h43c3e51a},
  {32'h44c61761, 32'hc3a961b2, 32'hc33c0f60},
  {32'hc4ba7ecb, 32'h42071bef, 32'hc2121201},
  {32'h45143d9b, 32'h434a51c3, 32'h43704145},
  {32'hc29aaaa0, 32'hc269d485, 32'h4393d556},
  {32'h44dcc356, 32'hc35091b9, 32'h428df310},
  {32'h433f3b00, 32'h4310fceb, 32'hc340652e},
  {32'h44b9ad6c, 32'h4267b71b, 32'h4333b30a},
  {32'hc4f696f6, 32'hc2884d0b, 32'h42f58fb3},
  {32'h44e21223, 32'hc25700ff, 32'h4364c9a8},
  {32'hc4aa311e, 32'hc2afc02e, 32'hc26f4235},
  {32'h44d1ea12, 32'hc1de1e2c, 32'h439982f0},
  {32'hc4905ed0, 32'hc33589c4, 32'hc1f9b64a},
  {32'h44e29618, 32'hc26a9e3f, 32'h43522545},
  {32'hc48c7d85, 32'h4258a4c5, 32'h42c38257},
  {32'h4337d090, 32'hc2a4bd2d, 32'hc32a4b01},
  {32'hc4ddd94f, 32'h43f30571, 32'h42959ab6},
  {32'h44af9c0b, 32'h4278226d, 32'hc388b71d},
  {32'hc50b60b3, 32'h408ccf3d, 32'hc38ba625},
  {32'h43854e44, 32'h43b80be0, 32'h43818ab1},
  {32'hc4e1bd5d, 32'hc380f966, 32'h41db3cf0},
  {32'h44b43dfd, 32'h427b7350, 32'h433d5186},
  {32'hc4bcfdc4, 32'h41a93537, 32'h432bce78},
  {32'h448beb14, 32'hc3cbe170, 32'h438f7ba5},
  {32'hc518f3ec, 32'hc2886fd2, 32'hc1c6a2cf},
  {32'h44688a15, 32'hc41e76ba, 32'hc23c7065},
  {32'hc36f1ab8, 32'hc37944ee, 32'h42df52d7},
  {32'h44dc0805, 32'hc38a80b1, 32'h434bf838},
  {32'hc4688bf9, 32'h429dd519, 32'h43b839a8},
  {32'h44fb6710, 32'hc33d3bae, 32'h42cc4c02},
  {32'hc438ff08, 32'h43931171, 32'hc3067754},
  {32'h433fc988, 32'h42422238, 32'hc37a4211},
  {32'hc503c8e1, 32'hc2e6f1be, 32'hc352cc19},
  {32'h4384fcf8, 32'h4384d831, 32'hc28a6fd3},
  {32'hc4e07ded, 32'h43a8b6d3, 32'h42cb663c},
  {32'h43a9105c, 32'h43a64242, 32'hc232b834},
  {32'hc4873b0b, 32'h43a456fc, 32'hc10cf91c},
  {32'h4522a142, 32'hc35f1d60, 32'h4136af50},
  {32'hc4823229, 32'hc32f4799, 32'h43a6746c},
  {32'h43eea9b2, 32'hc3044541, 32'hc3cf4447},
  {32'hc2aef054, 32'hc3419210, 32'hc3a0c7ad},
  {32'h4438bf2a, 32'hc37d9e6d, 32'h4207022d},
  {32'hc50e11e6, 32'h43f15fe1, 32'hc3d6024d},
  {32'h45312262, 32'h42ac3bb7, 32'hc3aa17d4},
  {32'hc4f3e158, 32'hc343dcc9, 32'h42389f0a},
  {32'h429d7880, 32'hc34c4a8a, 32'hc13ba3c2},
  {32'hc3462a80, 32'h439f42c4, 32'hc366b5b4},
  {32'h44c599cb, 32'h42a7e26d, 32'h42aef294},
  {32'hc4caa878, 32'h42f666f8, 32'hc378bcf7},
  {32'h44f25312, 32'h42a5f464, 32'hc2960c35},
  {32'hc5081de6, 32'hc2bddfd8, 32'hc32b90c4},
  {32'h43567ba8, 32'hc3b07e24, 32'hc342461f},
  {32'hc3b8c848, 32'h42c41e84, 32'hc20873f8},
  {32'h443fe7a6, 32'h429303f2, 32'h42c39b10},
  {32'hc4e60cad, 32'h4353c02c, 32'hc3438a1d},
  {32'h44894e39, 32'hc40ef77e, 32'hc3347672},
  {32'hc490e697, 32'hc1e0003c, 32'hc0d7a3e8},
  {32'h44d228f4, 32'hc31ba1c9, 32'h42bfb8fe},
  {32'hc4bd291e, 32'h43203792, 32'h428ab5de},
  {32'h43d78de0, 32'hc2c00707, 32'h40b943ec},
  {32'hc4a23698, 32'h41cd072e, 32'h437312ad},
  {32'h43a051b6, 32'h430ad1bf, 32'hc39550c8},
  {32'hc434471a, 32'hc1b2a027, 32'h4393c3ef},
  {32'h451d8115, 32'h428e703c, 32'h431e8627},
  {32'hc49781c9, 32'h43aeb1dc, 32'hc1819bef},
  {32'h450bfd5f, 32'hc25edce6, 32'h41a4cd0c},
  {32'hc4afed16, 32'h43aa74b5, 32'h41daf4c3},
  {32'h44f8a46a, 32'h4118b71b, 32'hc1d3c255},
  {32'hc46a2e23, 32'hc3748eab, 32'h441e7806},
  {32'h44b8d970, 32'h4226bf2c, 32'h42ffe902},
  {32'hc4624f90, 32'h429dbbe2, 32'h40fc41c5},
  {32'h44996384, 32'h436aa02b, 32'hc382d24b},
  {32'hc4fa629b, 32'hc3f5fe41, 32'h4248255f},
  {32'h42b831e0, 32'hc398742c, 32'h419324d0},
  {32'hc41352d6, 32'h4362b812, 32'hc2b3270a},
  {32'h438cef16, 32'h427b2670, 32'hc156f56d},
  {32'hc515addf, 32'h4348d3ff, 32'h424a483a},
  {32'h43ec4730, 32'h43fc5d37, 32'hc36064b1},
  {32'hc5155fff, 32'hc1fddb32, 32'h4295e92c},
  {32'h4482fb0c, 32'h43b22661, 32'h428b1756},
  {32'hc4d37e1c, 32'h42921c36, 32'h427cc21d},
  {32'h444a31a4, 32'hc314484d, 32'hc3bfd319},
  {32'hc4c2f381, 32'hc29eb786, 32'h41f96dd0},
  {32'h45103df0, 32'hc10949b5, 32'h4314574c},
  {32'hc50803b8, 32'h43de6639, 32'h437d6553},
  {32'h45287771, 32'h42e545c3, 32'hc3269e74},
  {32'h44819c63, 32'hc1845d72, 32'hc2b12e99},
  {32'hc48731bf, 32'h42f1d5db, 32'hc329f4fd},
  {32'h43ec6248, 32'h438c5528, 32'h43778e5d},
  {32'hc327b57c, 32'hc3880b38, 32'h432de8af},
  {32'h44bb2420, 32'h4325f79d, 32'hc399a8bf},
  {32'hc38dca30, 32'hc2c07bec, 32'hc35bd996},
  {32'h44ba035a, 32'hc30ac18e, 32'hc395ff14},
  {32'hc38edd48, 32'h42c2d498, 32'hc1d7f050},
  {32'h44b2a48a, 32'h425b9aaa, 32'hc36e76f2},
  {32'hc4632059, 32'hc26ab5e9, 32'h41ad7dbd},
  {32'h44bb2513, 32'hc34f59a4, 32'hc355620a},
  {32'hc4db8f96, 32'h431a1c70, 32'h435dadf6},
  {32'h43c00998, 32'hc197f970, 32'hc360198e},
  {32'hc4eea24c, 32'h41cf3eb3, 32'hc28ad89d},
  {32'h4466aa28, 32'hc2778720, 32'hc3e3385f},
  {32'hc4bb5eaa, 32'h434d4d31, 32'h43197b9b},
  {32'h442858fc, 32'hc323199b, 32'h4302d0f4},
  {32'hc50c3438, 32'h4036fadc, 32'h422f05bb},
  {32'h4498d50d, 32'hc3a51806, 32'h4380c30c},
  {32'hc45a2106, 32'h432d7687, 32'h43a04f00},
  {32'h42f95598, 32'hc1cb7332, 32'hc2b853d0},
  {32'hc40b03fc, 32'hc2dedb3a, 32'hc2943234},
  {32'h442fe0e4, 32'hc346405a, 32'hc3575c18},
  {32'h43838ea0, 32'hc05643ac, 32'h43370991},
  {32'h432da508, 32'hc329431b, 32'hc2f4b2bb},
  {32'hc50b29cd, 32'hc336fe94, 32'h43c84ce2},
  {32'h44768642, 32'hc38e2b1d, 32'h43d06e76},
  {32'hc5041624, 32'h438f0c97, 32'hc26d5530},
  {32'h44095b56, 32'h42e10d9d, 32'hc379df26},
  {32'hc432bfb6, 32'h4395d49c, 32'h418634e1},
  {32'h449fc977, 32'hc3ffd77f, 32'hc2c7b9ee},
  {32'hc49ab55a, 32'hc3b71f4a, 32'h424b7b64},
  {32'h4404e57a, 32'h43c23238, 32'hc3a661f7},
  {32'hc38cefdd, 32'h440688ad, 32'hc2d456d9},
  {32'h43096756, 32'hc36594c4, 32'hc3415181},
  {32'hc46b35d3, 32'h41600f42, 32'h43a2ce92},
  {32'h447d7edc, 32'h42cebf81, 32'hc38e56fc},
  {32'hc41a86fd, 32'h43fda339, 32'h428dacb7},
  {32'h446443f8, 32'h428f87fe, 32'h43b54251},
  {32'hc51d59a7, 32'h42ca3c8a, 32'h439316a1},
  {32'h44d0c964, 32'h42a15513, 32'hc2fdb7b0},
  {32'hc395007b, 32'h429ff2db, 32'hc38df11c},
  {32'h43983eba, 32'hc2a02851, 32'hc12afa46},
  {32'hc5028f01, 32'hc3d5b8dc, 32'h43316a24},
  {32'h438a8740, 32'hc309e9fe, 32'hc26001ea},
  {32'hc27bcf00, 32'h42a4378e, 32'hc3582722},
  {32'h443f5701, 32'hc385eb35, 32'h42c7a23c},
  {32'hc51f073a, 32'hc30fd176, 32'hc38c91de},
  {32'hc4476f7a, 32'h4217e8f1, 32'h419b2fde},
  {32'h450073ab, 32'h43b2f78c, 32'h4224d92d},
  {32'hc4a60dd1, 32'h4379fd59, 32'hc337260d},
  {32'h43ffeac0, 32'h41995ece, 32'hc20833e5},
  {32'hc512e198, 32'hc384d89f, 32'h4311e918},
  {32'h44aeb1f0, 32'h43795f80, 32'h42b41b76},
  {32'hc40e3ad8, 32'h43b36516, 32'h4206ce72},
  {32'h443a1432, 32'hc0ee4edc, 32'h42ce1a70},
  {32'hc4e7b15d, 32'hc33c661d, 32'hc1f8af20},
  {32'h4406a014, 32'hc3e654cf, 32'hc36a6106},
  {32'hc310a60c, 32'h40ba9b7e, 32'hc316b009},
  {32'h44f9c57d, 32'hc2c001d1, 32'hc368132f},
  {32'hc385eb46, 32'hc37da5e1, 32'hc35c5d17},
  {32'h44d5ae1c, 32'hc3a4d7ff, 32'h42775c9b},
  {32'h44df56e7, 32'h43dba93a, 32'hc346d8fa},
  {32'hc51bf431, 32'h4356d033, 32'hc3878083},
  {32'h442174b4, 32'h416bec0a, 32'hc2b98e3a},
  {32'hc4923d35, 32'h43a6e9eb, 32'hc3b5b5b6},
  {32'h44d2042b, 32'h4314d487, 32'h42910118},
  {32'hc4cb862f, 32'h426d892c, 32'hc29c37b9},
  {32'h439cca04, 32'h43b93766, 32'hc2295f64},
  {32'hc4bab816, 32'h415913f3, 32'hc3d4b4c1},
  {32'h44eb25a8, 32'h43b481b5, 32'h428274c0},
  {32'hc4a60b35, 32'hc2aa7582, 32'h44091568},
  {32'h443ee919, 32'h42fc52d3, 32'hc25b1eb0},
  {32'hc514d6be, 32'hc21538e3, 32'h41051f9e},
  {32'h436d1d2d, 32'hc209fcb6, 32'hc300ce76},
  {32'hc4ca25d6, 32'hc3aee3d5, 32'hc232ffd3},
  {32'h441917cd, 32'h42fee8ea, 32'h4134a93a},
  {32'hc4edb332, 32'h42f83946, 32'hc20226fc},
  {32'h450dbd7a, 32'h427ecdae, 32'h3e839514},
  {32'hc3856d80, 32'h4330db4e, 32'hc355dd84},
  {32'h45268b13, 32'h43b03845, 32'hc37d1c0e},
  {32'hc4632d7a, 32'h440ff57c, 32'hc2615ef0},
  {32'h44e3cf64, 32'hc234d17c, 32'hc3533b06},
  {32'hc511628b, 32'hc407bcab, 32'h42f6cc2f},
  {32'h44fea776, 32'hc3837860, 32'h432e7650},
  {32'hc490eb3e, 32'hc37679bc, 32'hc2196b6d},
  {32'h44e89ca4, 32'h4320c7ab, 32'h433feaac},
  {32'hc4a72e10, 32'h422f57ea, 32'h42f0420c},
  {32'h4327c464, 32'hc36138c2, 32'hc37a882a},
  {32'hc42fd6b5, 32'hc2baede0, 32'h42a7a7ed},
  {32'h43fc3670, 32'hc35b078b, 32'h42b43546},
  {32'hc48778bf, 32'hc34f9285, 32'hc33c02a1},
  {32'h44c36185, 32'h438f775b, 32'hc28016e4},
  {32'hc506a3a3, 32'h4299e542, 32'h42a6a114},
  {32'h4498c1d6, 32'hc2f9913b, 32'h43b127dd},
  {32'hc4781c70, 32'hc2b41d19, 32'hc29d2ae1},
  {32'h44954405, 32'h41e39df7, 32'h43b53159},
  {32'hc4a8ece5, 32'hc2e1ffe1, 32'hc32ed0fa},
  {32'h44b6e4bc, 32'hc35ab6d7, 32'h418443d8},
  {32'hc47494b8, 32'hc369393b, 32'hc32969d2},
  {32'h44d5cd99, 32'h44005320, 32'hc30c4c35},
  {32'hc50f5438, 32'h436c06c8, 32'hc2a32a9b},
  {32'h44b7c985, 32'hc3473dfd, 32'hc34625fe},
  {32'hc4dad7be, 32'hc28c4e37, 32'h43a4080a},
  {32'h4386ce49, 32'hc322864f, 32'h42732fef},
  {32'hc3b70e42, 32'hc37d89aa, 32'hc32403e7},
  {32'h44bf6d45, 32'h43dfc56e, 32'h42214c30},
  {32'hc4ca2fbf, 32'h4257252d, 32'hc2de0c19},
  {32'h4498367d, 32'h4101891f, 32'hc3eed9b4},
  {32'hc48bfe5f, 32'h42efe418, 32'hc359a019},
  {32'h440660bc, 32'hc1438f89, 32'hc11cada2},
  {32'hc3ae4efc, 32'hc2d1863f, 32'hc32de109},
  {32'h44af0924, 32'h43230af0, 32'h42899cf3},
  {32'hc508bdac, 32'hc319ec59, 32'h43f0394b},
  {32'h44527684, 32'hc31b271f, 32'h438e49fd},
  {32'hc50ce87c, 32'hc37d55ed, 32'hc23bb06f},
  {32'h44beea95, 32'hc15208ac, 32'hc291c09e},
  {32'hc4cb5c7a, 32'hc3541ffc, 32'h43cdc5f0},
  {32'h44908aac, 32'hc367a7f0, 32'hc33bc816},
  {32'hc4d85118, 32'hc2dd89b0, 32'h4313dcbe},
  {32'h4422503d, 32'hc3af3041, 32'h42e848dd},
  {32'hc39f5b8e, 32'hc34be977, 32'h432db8a3},
  {32'h450f6ba5, 32'hc16041a2, 32'h436754ab},
  {32'hc4917380, 32'hc0225470, 32'h4354fb4d},
  {32'h44885ec4, 32'hc34e05da, 32'h3ee38520},
  {32'hc46c97c8, 32'hc0c364de, 32'hc394c423},
  {32'h44825f93, 32'h43cb5822, 32'hc3c6f947},
  {32'hc49b7598, 32'h4338345e, 32'h43b4da2c},
  {32'hc3c579fe, 32'h43644359, 32'h43afb036},
  {32'hc429b056, 32'h434b0d43, 32'hc3a3bf4e},
  {32'h44965afd, 32'h42acebb2, 32'h43caaf96},
  {32'hc4c43ad1, 32'hc3b8d7b4, 32'hc405ed7f},
  {32'h4407a454, 32'hc2ab7c06, 32'hc1aa0204},
  {32'hc50f12a8, 32'hc355f99d, 32'hc00b87a9},
  {32'h44ea4cae, 32'h42e9c647, 32'hc2f78ebe},
  {32'hc49ada41, 32'hc346995b, 32'hc3613e1d},
  {32'h439ef618, 32'h434cecc3, 32'hc3ccdb2a},
  {32'hc3d156c8, 32'hc425356b, 32'h4400dc42},
  {32'h44043284, 32'hc342f2a6, 32'h432409bc},
  {32'hc4b95aa5, 32'hc3061970, 32'h42b90625},
  {32'h442b7eae, 32'h43b4d099, 32'hc394a238},
  {32'hc4682f8a, 32'h40907b5e, 32'h433b9993},
  {32'h43df4938, 32'hc28796c0, 32'h4317fe05},
  {32'hc3bea738, 32'hc15d8134, 32'hc39f7349},
  {32'h451d3eab, 32'hc21a63bc, 32'h4315aa29},
  {32'hc48e0dbe, 32'hc2e9268c, 32'h436cca1a},
  {32'h447a7249, 32'h41434c66, 32'hc24885ad},
  {32'hc5003708, 32'h43ebe2bd, 32'h4380041b},
  {32'h430e8f10, 32'h41c5789f, 32'h432b57b8},
  {32'hc4f9c825, 32'h43a73678, 32'h42440735},
  {32'h44e9db14, 32'hc319c9bd, 32'h425c8b4c},
  {32'hc4f3ee7b, 32'hc34bf4c1, 32'hc32d771c},
  {32'h432dc174, 32'h431058a6, 32'hc2d3663e},
  {32'hc4db397b, 32'hc3912692, 32'h4292e1c3},
  {32'h44ed0a4d, 32'h42ae2476, 32'hc2ce52bd},
  {32'hc4970f50, 32'h42d74336, 32'hc2e764cd},
  {32'h44b1bdca, 32'h409a9d18, 32'hc28dd305},
  {32'hc4f28b94, 32'hc390d84a, 32'h4349b3da},
  {32'h45082695, 32'hc377c19f, 32'h43b05361},
  {32'hc4a0a404, 32'hc3de6792, 32'hc3ad5877},
  {32'hc3459710, 32'h430b5e37, 32'hc35e7c31},
  {32'hc4b6c732, 32'h427407d3, 32'hc2ac9cb9},
  {32'h43d2138a, 32'h428692a6, 32'h4218b32f},
  {32'hc4ed8439, 32'hc20554ca, 32'h43c7064b},
  {32'h442804b6, 32'h43014ac6, 32'hc407f353},
  {32'hc4e9eccf, 32'hc3564d2d, 32'hc2fc1ebe},
  {32'h44118392, 32'hc3e26863, 32'h428769ca},
  {32'hc4493655, 32'hc2b6050d, 32'h4385c866},
  {32'h450d28df, 32'h43948a1b, 32'hc40e0968},
  {32'hc4d8384e, 32'h43a759ec, 32'h434821bb},
  {32'h4440fba6, 32'h43414349, 32'hc32e987a},
  {32'hc3159d8e, 32'h4311f5d8, 32'h433b5077},
  {32'h4465e314, 32'h438fd3fa, 32'hc3d353be},
  {32'hc4d370af, 32'hc2edf6e6, 32'hc34bee78},
  {32'h44fb2e8e, 32'hc19bd456, 32'h422c1bf2},
  {32'h4312c078, 32'h41633dfc, 32'hc3804245},
  {32'h4486c07d, 32'h438fec5d, 32'h432c106d},
  {32'hc4b2fd33, 32'h41526f2f, 32'h42b7a4f6},
  {32'h44678968, 32'h43af29da, 32'hc0de546c},
  {32'hc39ac0b0, 32'hc1bcb342, 32'hc3aa7bbf},
  {32'h44ed4730, 32'hc3549ea1, 32'h4393d1f8},
  {32'hc4fe21d7, 32'hc2b89ce8, 32'h42851628},
  {32'h448582b6, 32'hc342bc03, 32'hc3bf5372},
  {32'hc3ffeb2e, 32'h429175f8, 32'h428f0c05},
  {32'h45105aa2, 32'h436e1072, 32'hc2b4a6f3},
  {32'hc496c5cf, 32'h42245991, 32'hc32762bc},
  {32'h44bd131d, 32'hc21cce3a, 32'hc37f8753},
  {32'hc3372d38, 32'h4417b042, 32'h431964e3},
  {32'h4504af66, 32'h42477388, 32'h412310fe},
  {32'hc4f1b610, 32'hc32a6364, 32'h4367ec00},
  {32'h4450db76, 32'hc2f3d6ab, 32'hc36f2d22},
  {32'hc39d9d84, 32'h434b700a, 32'h438d0ff3},
  {32'h444ac257, 32'hc2b23600, 32'hc2ba877c},
  {32'hc3316718, 32'hc2400395, 32'h42b5e46d},
  {32'h450ca3dd, 32'hc3bf058f, 32'hc38c44f2},
  {32'hc45a7dae, 32'hc35b4a9d, 32'h42ff75c8},
  {32'h44eeb507, 32'hc287b6e0, 32'h4323c7a8},
  {32'hc50c6fdc, 32'hc2b17b81, 32'hc1b24dbe},
  {32'h44a4a124, 32'h43b320ae, 32'hc36c4a3d},
  {32'hc43dfad8, 32'h439793d6, 32'h42bed92c},
  {32'h43abb1a6, 32'h438157b8, 32'h4286e03e},
  {32'hc500e98c, 32'h42910ba3, 32'h4165d4c8},
  {32'h43c49d00, 32'h4270c9dd, 32'h44082a34},
  {32'hc40326da, 32'h437861f8, 32'hc3c1c106},
  {32'h44f34a61, 32'h416c44e5, 32'h41edd3be},
  {32'hc4d4c720, 32'hc3c3eea7, 32'hc394b6a6},
  {32'h450af2f8, 32'h42ea8761, 32'h42541c68},
  {32'hc4b8021d, 32'h432eb77d, 32'hc21a7de1},
  {32'h443b5120, 32'h43a67292, 32'h43dcd261},
  {32'hc208eb50, 32'hc3624706, 32'hc37aaf6b},
  {32'h436c2290, 32'hc2020700, 32'hc3de16c2},
  {32'hc40f80f8, 32'hc38380ed, 32'hc2fadae2},
  {32'h449d2232, 32'h43d66071, 32'hc30ce674},
  {32'hc5025708, 32'hc3122ada, 32'hc31043db},
  {32'h442ca7b2, 32'h41cdde68, 32'hc38d50d5},
  {32'hc45f62ac, 32'h4384b55e, 32'h42b71fcf},
  {32'h4361cdd8, 32'hc3cefa59, 32'h42f2b218},
  {32'hc42f923c, 32'hc35cd989, 32'hc12661ad},
  {32'h44cb30df, 32'hc30e25b8, 32'h40363190},
  {32'hc4a5b084, 32'h43e82c3d, 32'h41d4310c},
  {32'h444f6b6e, 32'h4395784e, 32'h423d1518},
  {32'hc44b6aac, 32'h43802fcd, 32'hc333bffd},
  {32'h44b2f42a, 32'hc261b905, 32'hc32310ef},
  {32'hc2c9e140, 32'h433d1856, 32'hc263536c},
  {32'h44d54e2e, 32'h4306ac29, 32'h439338d6},
  {32'hc4aeda10, 32'h434420bd, 32'hc32a250f},
  {32'h4509ada2, 32'h42086f72, 32'hc2908206},
  {32'hc3cc8e1b, 32'hc191e5d9, 32'h43635df6},
  {32'h4502ed72, 32'h42147c9b, 32'h4329f7c8},
  {32'h42d435f2, 32'hc30095b2, 32'hc3b20681},
  {32'h44d48e99, 32'h431adf04, 32'hc0484a18},
  {32'hc4887229, 32'hc2b14340, 32'hc1ca5d3f},
  {32'h4510d1b1, 32'hc3dab7e9, 32'hc2ec38e8},
  {32'hc4a9fcd4, 32'hc388ea73, 32'h432f824a},
  {32'h443e82a4, 32'h417ff3ec, 32'h4344c0ff},
  {32'hc501c2e8, 32'h437f5652, 32'hc320bb07},
  {32'h44f183a7, 32'h43d45be5, 32'h4328935b},
  {32'hc506dbb4, 32'h43147fd6, 32'h43155755},
  {32'h44195e5e, 32'hc33ee921, 32'h439dfd9a},
  {32'hc49777e7, 32'h4392fc36, 32'hc26ea1bf},
  {32'hc2a96bd0, 32'h42893600, 32'h4281b693},
  {32'hc3f87fd0, 32'h42bc638f, 32'h43f729d1},
  {32'h4452afb2, 32'h433f9a17, 32'h40b2ce8b},
  {32'hc510942a, 32'h4339ca3e, 32'hc292a7e9},
  {32'h44dd712f, 32'hc2d17a6b, 32'h425b3037},
  {32'hc4dcfca8, 32'h42d1464f, 32'h425f3f58},
  {32'h44d4ec3e, 32'h432fb6d1, 32'hc347223c},
  {32'hc4dbe5f6, 32'hc1ed7227, 32'hc29f3df3},
  {32'h44e238aa, 32'hc3a4459e, 32'hc1a39413},
  {32'hc501cb18, 32'hc35fb51b, 32'h433be0a7},
  {32'h450c2574, 32'h4390ade9, 32'hc372a453},
  {32'hc47518f4, 32'h438a20ad, 32'h43659f88},
  {32'h44870734, 32'hc382a4a0, 32'h422d0e81},
  {32'hc3c3e53c, 32'hc27b8946, 32'h437be732},
  {32'h44b6dff0, 32'hc3432ff7, 32'hc38916b0},
  {32'hc4f5af17, 32'h432db0f8, 32'h426fe87e},
  {32'h44fd4307, 32'h42fa6715, 32'hc2167f86},
  {32'hc4bfcccd, 32'hc2d5eb4b, 32'h4336475b},
  {32'h4508f54e, 32'h43b3768a, 32'h43970cf2},
  {32'hc2cd7ac0, 32'hc2be0a09, 32'hc18bf622},
  {32'h4488a661, 32'hc31539ec, 32'hc3acb593},
  {32'hc1ae7800, 32'h435921ad, 32'h43071b91},
  {32'h43acd3c8, 32'hc451f6c3, 32'h4307d45a},
  {32'h43a08fa0, 32'h42175840, 32'h431701a3},
  {32'h44ac4d4a, 32'h42aca3de, 32'hc3442734},
  {32'hc4b3a0e3, 32'hc2ff54ba, 32'hc4071d18},
  {32'h450c02b9, 32'h42b7eeed, 32'h431bfc01},
  {32'hc3a99bfa, 32'hc23d1138, 32'hc3772b87},
  {32'h4383b7cd, 32'hc3f0ff9c, 32'h420fffaa},
  {32'hc2eb5b90, 32'hc3f98027, 32'hc266d9cc},
  {32'h43a5db3a, 32'h43d30666, 32'hc354de5d},
  {32'hc4c85c3e, 32'hc314607f, 32'hc38b531e},
  {32'h44393ed8, 32'hc37aee3b, 32'hc42d5e7e},
  {32'hc50da880, 32'h43f9e59b, 32'hc22e02c0},
  {32'h44e301d5, 32'hc3e5b63c, 32'hc3080233},
  {32'hc4e8e0b7, 32'hc351380f, 32'hc350d3ae},
  {32'h4513d2ba, 32'h4194a311, 32'h43546379},
  {32'hc433cce9, 32'h42addb93, 32'h431d38d6},
  {32'h43f1e1c5, 32'hc259d225, 32'h43434f64},
  {32'hc4685a94, 32'hc09ca39c, 32'h43799437},
  {32'h44461ad0, 32'hc4005d59, 32'h440aa560},
  {32'hc3f8a583, 32'hc3fd8772, 32'h43a5e630},
  {32'h44a3f721, 32'h43abf708, 32'hc334fcfa},
  {32'hc4b69f5c, 32'hc2e7fddc, 32'h436122c8},
  {32'h45047f9a, 32'hc2e8a95c, 32'h42f9f3dc},
  {32'hc4490ed2, 32'h438ce864, 32'h4385e6a6},
  {32'h449652bb, 32'h43f5322d, 32'hc24c842e},
  {32'hc43c344f, 32'h43ee0b15, 32'h42485383},
  {32'h43dcf010, 32'hc1f4f274, 32'hc3b900b2},
  {32'hc50e5907, 32'h431145b4, 32'h438ec18e},
  {32'h42b2a59e, 32'h43863252, 32'h43164857},
  {32'hc4b3eedf, 32'h42c7b2e2, 32'h43737319},
  {32'h43b9b4a9, 32'hc3012ac0, 32'hc3939df6},
  {32'hc504401e, 32'h43899905, 32'h43827629},
  {32'h4491fb34, 32'h40f037f5, 32'hc30e49ee},
  {32'hc4f2ca7d, 32'h436bccae, 32'h43f09c75},
  {32'h447b7e6d, 32'h4318ea0b, 32'hc2b9c476},
  {32'hc3fe8a10, 32'hc1c1c2ff, 32'hc3479191},
  {32'h4440be3b, 32'hc28a756e, 32'h42da09c6},
  {32'hc505aa42, 32'h43575d34, 32'hc34fe1ef},
  {32'h42dc48f4, 32'h42623c70, 32'hc337ce5f},
  {32'hc4d210a5, 32'hc3a1f4b3, 32'h423b7f8a},
  {32'h43b1563c, 32'hc2f2e25a, 32'h4251057e},
  {32'hc5061414, 32'hc30abe16, 32'hc2698184},
  {32'h44faf6d6, 32'hc2f9753d, 32'h43623455},
  {32'hc3acd2ea, 32'h4342c3d9, 32'h43837821},
  {32'h443e4efc, 32'h43a8bd66, 32'h437272c4},
  {32'hc4b78006, 32'hc26dc3de, 32'h43f2bd89},
  {32'h447f03dc, 32'hc2f14ca1, 32'h41b51f6b},
  {32'hc3757794, 32'h411d2537, 32'h414fda45},
  {32'h428caa07, 32'h440989e9, 32'h4311f13c},
  {32'hc4d15252, 32'h430059f5, 32'hc26f6eaa},
  {32'h44767130, 32'h431de271, 32'hc219df1a},
  {32'hc3215e87, 32'h43509054, 32'hc2667bc4},
  {32'h4440f5cc, 32'h43a7ab64, 32'hc2c8a62c},
  {32'hc4fe1e42, 32'h43cc8a72, 32'hc3bb4059},
  {32'h449e7651, 32'hc33ee88a, 32'hc3255eea},
  {32'hc3ca76fd, 32'hc3adf997, 32'hc2dc177b},
  {32'h44e97b7d, 32'h42a58e7c, 32'h42ccddb4},
  {32'hc432fcb4, 32'hc2d390fe, 32'h432dce96},
  {32'h441460d8, 32'h4386b428, 32'h4342c555},
  {32'hc4229b1a, 32'h42373670, 32'hc289a701},
  {32'h44f8b076, 32'hc2bf3fc7, 32'h430a08f1},
  {32'hc4ef4727, 32'h434bfacc, 32'hc2ea7366},
  {32'h439b34fa, 32'hc11114e4, 32'hc218c707},
  {32'hc3c46044, 32'h43053611, 32'hc396b7b2},
  {32'h4355023c, 32'h434b8df9, 32'h42fb74f4},
  {32'hc517962f, 32'hc2e001c9, 32'h430a74ed},
  {32'h43c962ad, 32'h4240a1b2, 32'hc31f2b10},
  {32'hc3f94a50, 32'hc37607d1, 32'h4216b4b8},
  {32'h4482b43b, 32'hc380c2ae, 32'hc1e67f86},
  {32'hc5008132, 32'h432bae45, 32'hc2e6beb1},
  {32'h450a5e58, 32'hc3a440b1, 32'hc3ae7d78},
  {32'hc51ee95a, 32'hc33b13d6, 32'hc2dbcc5a},
  {32'h448a54a0, 32'hc399127f, 32'hc2789ab0},
  {32'hc4c7ef6d, 32'hc116c47a, 32'hc367bb45},
  {32'h4502120f, 32'hc345b8cb, 32'h4284f18d},
  {32'hc3b34f8a, 32'hc3330616, 32'hc19725b8},
  {32'h4517652e, 32'h4377e0b9, 32'hc3576b6c},
  {32'hc5030187, 32'h43ad3f87, 32'h4228f8f4},
  {32'h44a2c94e, 32'hc28d139c, 32'h432236ff},
  {32'hc504a8da, 32'h42cd2040, 32'h432cf94f},
  {32'h44da173d, 32'h43738762, 32'hc335cbc7},
  {32'hc4ba7b2e, 32'h4338ada0, 32'hc3c3be2d},
  {32'h4235f000, 32'h42876627, 32'h43fd40c2},
  {32'hc493e593, 32'h43b9bf9a, 32'h424549e1},
  {32'h44bebc93, 32'h418a5b5a, 32'hc420ad21},
  {32'hc4762034, 32'hc23a075f, 32'h411c17f8},
  {32'h45073131, 32'hc2e45c18, 32'hc3b609cb},
  {32'hc5188980, 32'h4396b94e, 32'hc1e7cf0e},
  {32'h43d163e4, 32'hc1d552a3, 32'hc2e981b1},
  {32'hc383f2fb, 32'hc389bd8c, 32'h43b23efe},
  {32'h441c9677, 32'hc33d093f, 32'h4388f018},
  {32'hc398a2f3, 32'hc2bd283b, 32'hc3142844},
  {32'h43b1b888, 32'h436007cf, 32'h43fdcec5},
  {32'hc4ca38bd, 32'hc2828c18, 32'hc23cd377},
  {32'h43f12f38, 32'hc317134a, 32'h430dfc09},
  {32'hc504eb59, 32'hc30fd19c, 32'h42ebfd5b},
  {32'h44a215dc, 32'hc3826bfb, 32'h429867d5},
  {32'hc4a18424, 32'h42e81d63, 32'h40dd2ed4},
  {32'h45045095, 32'hc30eb692, 32'hc3669cdc},
  {32'hc4d0ba48, 32'h431ffd52, 32'h40c7e7e0},
  {32'h43af717a, 32'hc369f34f, 32'hc1f097d4},
  {32'hc50ab38e, 32'hc2847327, 32'hc2f8287b},
  {32'h43acc9e4, 32'h42ffe982, 32'hc33c64c0},
  {32'hc4df1eab, 32'hc2279db0, 32'h434e574c},
  {32'h44760191, 32'h438addff, 32'hc225a398},
  {32'hc4394cca, 32'hc3978be6, 32'h4293af67},
  {32'h43454650, 32'h432fb3c1, 32'h408b2ec6},
  {32'hc41b561c, 32'h43af773c, 32'h42f0e82a},
  {32'h44e37d89, 32'hc350e8f2, 32'hc2c1b19b},
  {32'hc466a210, 32'hc2d49b62, 32'h43fd761f},
  {32'hc3028236, 32'h42c48b24, 32'hc26285d0},
  {32'hc51333c6, 32'h4222c8c0, 32'h439a562a},
  {32'h44bb3634, 32'h43a83900, 32'hc3392556},
  {32'hc4666f05, 32'h42cd30c9, 32'hc2cd09f5},
  {32'h440d336f, 32'h43d428e9, 32'hc3208564},
  {32'hc4aa9c55, 32'h42ba3e7f, 32'h428436aa},
  {32'h439d3648, 32'h436f7728, 32'hc24c7e49},
  {32'hc4bffbb7, 32'hc380534b, 32'h425cae6b},
  {32'h4400a05c, 32'hc2f7cff1, 32'hc2ef183f},
  {32'hc456df01, 32'h411eed2b, 32'hc3f00ff9},
  {32'h43c59516, 32'hc22d82e6, 32'h42ada759},
  {32'hc4b9c9b1, 32'hc36773a1, 32'hc279d464},
  {32'h43b5d648, 32'h421f2d4b, 32'hc38a1681},
  {32'hc48ba04a, 32'h42af3369, 32'hc2be72a5},
  {32'h450de93e, 32'h4293a540, 32'h438300f0},
  {32'hc4ac7d14, 32'h42eb0781, 32'hc2ad3977},
  {32'h4400329a, 32'hc024cc9f, 32'h43f32636},
  {32'hc4d11191, 32'hc3b4e021, 32'h43be1363},
  {32'h4503aa3a, 32'h41477d34, 32'hc3664847},
  {32'hc42de6e8, 32'hc3a7f3da, 32'hc33350af},
  {32'h43809e12, 32'h429b42ef, 32'h42054e9b},
  {32'hc50395b6, 32'hc387718d, 32'hc276b342},
  {32'h43b7d088, 32'hc191e7c9, 32'hc3142151},
  {32'hc4726d42, 32'h43beb127, 32'h41c41cfd},
  {32'h44d87b3d, 32'h42cb0aca, 32'hc3dbd727},
  {32'hc45cd178, 32'hc291c956, 32'h426d93d5},
  {32'h451a222b, 32'hc23d7b7e, 32'h433ed458},
  {32'hc4866589, 32'hc43a6fce, 32'hc2826dc6},
  {32'h44e61ce4, 32'hc35ec69b, 32'h434290dc},
  {32'hc50286f4, 32'hc3411866, 32'h435cfb8c},
  {32'h44481d98, 32'hc13c81f6, 32'h441cab6e},
  {32'hc31f361c, 32'hc271d995, 32'hc343c552},
  {32'h448ed72a, 32'hc253ee86, 32'hc1ccd8b4},
  {32'hbf8a07d0, 32'hc33ea9d6, 32'h432a49c4},
  {32'h44bf3583, 32'h437c4e1a, 32'h43ca54f3},
  {32'hc3d19b48, 32'hc01b9615, 32'hc39b1edb},
  {32'h44e83f6d, 32'hc2e46ca1, 32'h42afa244},
  {32'h422910c0, 32'hc33dd125, 32'h43b5d8e3},
  {32'h44fe7fe5, 32'hc3465a0a, 32'hc31d242d},
  {32'hc4dd3f15, 32'hc2c23d49, 32'hc3720ed5},
  {32'h44641a8a, 32'h42637b88, 32'h43c5ecea},
  {32'hc50195b4, 32'hc3b196e3, 32'h42fdf9c9},
  {32'h43dfcd36, 32'h41c512e2, 32'hc2d5f2e7},
  {32'hc48a005a, 32'hc32a3ae9, 32'hc2257fd8},
  {32'h43ccd30c, 32'hc22ab40e, 32'h43c0dec3},
  {32'hc415bf00, 32'hc0f41c58, 32'hc2fdf687},
  {32'h44ee15d7, 32'h4395af09, 32'h4371b293},
  {32'hc3a84ba0, 32'hc3deca80, 32'h431046d3},
  {32'h44e52179, 32'hc307e239, 32'h429b037e},
  {32'hc4a2643f, 32'hc31928d8, 32'hc39ff3c7},
  {32'h449180f8, 32'h431694b8, 32'hc2c3e4d5},
  {32'hc43840c0, 32'h4386c10c, 32'hc39209ca},
  {32'h45082447, 32'h436c6893, 32'hc3aaeeb8},
  {32'hc3881c18, 32'hc2808f1a, 32'hc3217d7e},
  {32'h44136319, 32'h4347d5fd, 32'h43be0ea7},
  {32'hc48a8dd2, 32'h4271790a, 32'hc327ced5},
  {32'h437dcb84, 32'h430de5ea, 32'h43ce8721},
  {32'hc46a0c8e, 32'hc388f943, 32'hc3adfad6},
  {32'hc41ea7b6, 32'h4331c6f4, 32'hc3454af5},
  {32'h44d41204, 32'h43779500, 32'h429919e7},
  {32'hc4df627e, 32'hc32b38b2, 32'hc36b92c2},
  {32'h444e6d18, 32'hc20e425b, 32'h433c5494},
  {32'hc4918d93, 32'hc219bc56, 32'hc31fec8e},
  {32'h4400bcc4, 32'h420baa93, 32'h43da977a},
  {32'hc5012b24, 32'hc26744ae, 32'hc29f10a7},
  {32'h44000bed, 32'h43d13050, 32'hc337bc34},
  {32'h4365fb70, 32'h41ab8c60, 32'hc3bea598},
  {32'hc303fafa, 32'hc1c4c2ff, 32'hc2c43d63},
  {32'hc5051c36, 32'hc3520c7c, 32'hc402cef0},
  {32'h43caa848, 32'hc338daeb, 32'h4356bb42},
  {32'hc4f8e836, 32'h42e490b8, 32'hc2ff029d},
  {32'h44ce6ef2, 32'hc244970e, 32'h4365591f},
  {32'hc3d81435, 32'h42ca0ca5, 32'hc18e952c},
  {32'h43ceb6da, 32'hc398305c, 32'hc38ef3d6},
  {32'hc49318ce, 32'hc27d4a05, 32'h41844dad},
  {32'h45043cde, 32'h428e0404, 32'h4331ae07},
  {32'hc4dbedb9, 32'hc1e04fde, 32'h420c4b3c},
  {32'h448520f1, 32'hc2ad4f53, 32'h43e402e4},
  {32'hc49b3f6e, 32'hc2236c42, 32'hc22bb850},
  {32'hc0955800, 32'h433ce5e5, 32'hc2bf419c},
  {32'hc506e822, 32'h4370ebd4, 32'h432923bf},
  {32'h44b30d32, 32'hc33684a2, 32'h425303ec},
  {32'hc353d31c, 32'hc3f0e16c, 32'hc281087d},
  {32'h44f30374, 32'hc30b8394, 32'hc36300f2},
  {32'hc4c8e67c, 32'hc3a8213d, 32'hc32224d5},
  {32'h44df2087, 32'hc31ffcdd, 32'h41da2b28},
  {32'hc3a7d0b0, 32'h4346b4b6, 32'hc39f821b},
  {32'h44886778, 32'h41cd8db2, 32'hc33c88fa},
  {32'hc352c900, 32'h43952be3, 32'hc398f8c9},
  {32'h44884cce, 32'hc391d7ea, 32'hc1ce6b26},
  {32'hc4a1c6e5, 32'h422d260e, 32'hc28814e8},
  {32'h4455e7a4, 32'hc25a70e9, 32'h4297eb24},
  {32'hc4ddc0fa, 32'h42cea49e, 32'hc38b34c9},
  {32'h44ff8f80, 32'hc33e0eb6, 32'hc31485e7},
  {32'hc3f3dda6, 32'hc3142c1f, 32'hc3ee6999},
  {32'h44c2804e, 32'h430c81c5, 32'hc2d0d346},
  {32'hc4134202, 32'hc371e35b, 32'h43127fe9},
  {32'h44ab0849, 32'hc2d8abb3, 32'h4344a4c8},
  {32'h44ffeb70, 32'hc348a52a, 32'hc2a41d06},
  {32'hc437aa18, 32'hc2f260d2, 32'h424e1b7c},
  {32'h43117770, 32'hc225cabb, 32'h435a8b76},
  {32'hc520f283, 32'hc399c448, 32'hc372ece5},
  {32'h439eb64e, 32'h440adaf1, 32'hc309a3ec},
  {32'hc51a10b5, 32'h436754a9, 32'h431eb78b},
  {32'h44fb9ead, 32'h438ee506, 32'hc377e3bf},
  {32'hc4f38489, 32'h43616fa3, 32'hc22265bc},
  {32'h44eb8ee6, 32'hc21f2dbb, 32'h41d59583},
  {32'hc4dbab42, 32'h417f9148, 32'h43855bb9},
  {32'h44b2d667, 32'h4382bc15, 32'h43abe4f3},
  {32'hc5145b2a, 32'hc3e1733f, 32'h42ad3893},
  {32'h451aafa6, 32'hc382e271, 32'h42d47ebb},
  {32'h4380728a, 32'hc25ccce5, 32'h43b2952a},
  {32'h44d670b6, 32'h4260150c, 32'hc3b76568},
  {32'hc4594df4, 32'h424c31ad, 32'h43d42be7},
  {32'h4506e059, 32'hc22c32db, 32'hc371f25c},
  {32'hc3d52f08, 32'h43444391, 32'hc3a1a9f5},
  {32'h44eaec4b, 32'hc36aeb07, 32'h4217dcc1},
  {32'hc48d2748, 32'hc323b801, 32'hc3038336},
  {32'h45094ad5, 32'hc39305aa, 32'hc2e64ebd},
  {32'hc5040894, 32'h426d830f, 32'hc260c2c0},
  {32'h446dcbd6, 32'hc304e969, 32'h4193d79f},
  {32'hc503c1af, 32'hc3270a7e, 32'hc2869273},
  {32'h4446d333, 32'hc3cee4e8, 32'h4206fa81},
  {32'hc4f15b1e, 32'hc43663b9, 32'hc27b0100},
  {32'h430bb874, 32'h42294cd2, 32'hc33c9d7b},
  {32'hc513f76d, 32'h435723a7, 32'hc3323364},
  {32'hc35c3830, 32'hc3d04250, 32'h43f38e9c},
  {32'h40a1d100, 32'hc30a7e43, 32'h42e1cd62},
  {32'h44e132db, 32'hc3e2d9ed, 32'h4192c3f6},
  {32'hc4fbd674, 32'h431593d8, 32'hc319be17},
  {32'h44d903fa, 32'hc30af6e5, 32'hc391c5b4},
  {32'hc4c30a0f, 32'hc31559c2, 32'h428ba305},
  {32'h44a2428d, 32'hc296105c, 32'h43512b98},
  {32'hc453b880, 32'hc2450199, 32'hc30db276},
  {32'h4325b1c8, 32'h433a0b1d, 32'h4314c3c9},
  {32'hc49247ba, 32'h439d261a, 32'hc32bca7e},
  {32'h44d7b888, 32'hc394e1d1, 32'hc39b1c67},
  {32'hc50e53f2, 32'hc430f777, 32'h434049f9},
  {32'h4509e7b1, 32'hc21c6524, 32'hc1e726ff},
  {32'hc49fdbf2, 32'hc22393ef, 32'h433e1d0c},
  {32'h44e8262a, 32'h429a2977, 32'h44044dce},
  {32'hc35e5ac2, 32'hc1665282, 32'h4321355f},
  {32'h450100df, 32'hc27d3794, 32'hc3080959},
  {32'hc4a729aa, 32'hc1211795, 32'hc38f4c45},
  {32'h44a1a0f1, 32'h434389d2, 32'h41cb03a6},
  {32'hc4a12a32, 32'hc3dfd563, 32'h439ac7a1},
  {32'h44752518, 32'hc39d469f, 32'hc372957a},
  {32'hc4a0d5bb, 32'hc3793b07, 32'hc2b2a9e6},
  {32'h4496e2e7, 32'h41612720, 32'h4268a5ea},
  {32'hc4afbc17, 32'h429f0bc0, 32'h42d9a542},
  {32'h44a3f3a2, 32'hc370b278, 32'hc26587b4},
  {32'hc496c202, 32'hc35341e3, 32'hc31a3f09},
  {32'h442515fc, 32'h419c7ccd, 32'h42d9364f},
  {32'hc4da3f5f, 32'hc2af98a0, 32'h428ffaac},
  {32'h4483f856, 32'h42e8d038, 32'hc2a98b37},
  {32'hc481b31e, 32'h4296123a, 32'h438db21f},
  {32'h45067aa2, 32'h4329b445, 32'h41d2b3d6},
  {32'hc256dd99, 32'h4362798a, 32'hc3a048cb},
  {32'h44b857d9, 32'hc3372337, 32'hc39c36cb},
  {32'hc42a28ad, 32'h42a1ddb7, 32'h4257beb9},
  {32'h44ad51eb, 32'h44045108, 32'h433f2f9b},
  {32'hc46d49c3, 32'hc3c6961f, 32'hc3cdd445},
  {32'h44767dfd, 32'hc2fe26ef, 32'h432c79f4},
  {32'hc508ad19, 32'hc2494a17, 32'hc330a6ec},
  {32'h4345155c, 32'h425054b0, 32'hc35d31af},
  {32'hc503e4ae, 32'h43b9b503, 32'hc34aa694},
  {32'h44d70cc8, 32'hc325b5ee, 32'hc3a070bf},
  {32'hc2f60e25, 32'hc3040253, 32'hc35c614d},
  {32'h44a37a85, 32'h4313e6d4, 32'hc3046765},
  {32'hc4a19999, 32'hc39455d6, 32'h42df7ae9},
  {32'h444a295e, 32'hc35716f2, 32'h4241fc78},
  {32'hc527a1b8, 32'hc3328e7d, 32'hc14eec86},
  {32'h44165b0c, 32'hc264cc91, 32'hc40150df},
  {32'h43bead62, 32'hc0a7d013, 32'hc3631857},
  {32'hc51bf786, 32'h43ca61a1, 32'hc3ba2f09},
  {32'h450c9e51, 32'h437a2e83, 32'hc227bad7},
  {32'hc476e9b1, 32'hc2a7485f, 32'hc2464e70},
  {32'h448ab601, 32'h42766b1f, 32'h434df3d4},
  {32'hc4a732ea, 32'h41b81ed4, 32'h43a7ae32},
  {32'h449bd48a, 32'hc107ef94, 32'h416d176c},
  {32'hc38acb3a, 32'hc2862942, 32'hc2c145c5},
  {32'h4387c66e, 32'h42a97538, 32'h433998d4},
  {32'hc46c9a23, 32'hc3147ae3, 32'h419726aa},
  {32'h44dc9d53, 32'hc40ff79c, 32'h40a266ab},
  {32'hc4e9a2cf, 32'hc3c53672, 32'h437bbe4f},
  {32'h4453d3c2, 32'hc2160471, 32'hc3191c42},
  {32'hc37b3b70, 32'hc38556ed, 32'h41cc9dc2},
  {32'hc403a84e, 32'h42a193dc, 32'hc386a740},
  {32'h44a23d63, 32'hc30d2ab0, 32'h429a4432},
  {32'hc4dfd362, 32'h434baeb9, 32'hc2dd51c2},
  {32'h4501e0a4, 32'hc3270499, 32'hc369cb78},
  {32'hc5062f19, 32'hc2af5e81, 32'hc2dd3d2c},
  {32'h440b32ab, 32'hc3501067, 32'hc2776ffb},
  {32'hc4398182, 32'hc385ade8, 32'hc3170f1a},
  {32'h448a782f, 32'h42297f32, 32'h41dd8231},
  {32'hc5077a17, 32'hc30999bf, 32'h438cb78a},
  {32'h44fa8a4a, 32'hc2b13cda, 32'h423b9566},
  {32'hc4a77dd1, 32'hc2da385d, 32'h43f02d07},
  {32'h44d586fa, 32'h4364ae0d, 32'hc2a969de},
  {32'hc4927384, 32'h43406a1e, 32'hc0a407a4},
  {32'h445161c3, 32'h433d0f6f, 32'hc3a33100},
  {32'hc5152ee8, 32'hc3aa1125, 32'hc2f1f835},
  {32'hc2ff9790, 32'h438124d5, 32'h41fe4dbd},
  {32'hc4eef8b6, 32'h43abbcbd, 32'h438144f2},
  {32'h44c594a5, 32'h41f81b22, 32'h4387627a},
  {32'hc2596120, 32'hc38620a3, 32'hc31e7562},
  {32'h43bfcba7, 32'hc40aa4c1, 32'hc39ccb83},
  {32'hc3bee4e5, 32'h424ef119, 32'hc0095bef},
  {32'hc34f6ac8, 32'h42cb2a3a, 32'h42f42f3e},
  {32'hc46768ab, 32'hc272e4f2, 32'h434965d3},
  {32'h44ec4e84, 32'h41802a02, 32'h42271372},
  {32'hc47aaa20, 32'hc397d5a4, 32'hc21a76cd},
  {32'h4281d038, 32'hc30d660d, 32'hc2aa14ff},
  {32'hc4dc4960, 32'hc321e6eb, 32'hc3895895},
  {32'h429c0499, 32'hc27ab521, 32'h440c84a6},
  {32'hc42f79cc, 32'hc3e4749c, 32'hc27b9c4e},
  {32'h4381503c, 32'hc231b600, 32'hc2bc1950},
  {32'hc393a668, 32'h42068f48, 32'hc10e6e2e},
  {32'h43cbd0e4, 32'hc3d19e62, 32'hc2fcdb62},
  {32'hc48231a1, 32'h4221aa0a, 32'h4210c867},
  {32'h4328d798, 32'hc34ba235, 32'hc2ea72e6},
  {32'hc47a4f97, 32'hc2863792, 32'h41b43070},
  {32'h44175a15, 32'hc3b00c65, 32'hc27dc73e},
  {32'hc451b0de, 32'h4260b7dd, 32'hc35e47e5},
  {32'h44908372, 32'h436bce04, 32'h42b338fe},
  {32'hc31d1c10, 32'h43a99b39, 32'h43778bbf},
  {32'h44a0a6f3, 32'hc2d9516c, 32'h4362f7d8},
  {32'hc4a4c764, 32'h423dfb94, 32'h4225dc7d},
  {32'h448167d3, 32'hc3580c66, 32'hc4097377},
  {32'hc4bc23be, 32'h428d0ae5, 32'hc2ea50dc},
  {32'h43cf9cb0, 32'h419b6b56, 32'h43b1b001},
  {32'hc25e01c0, 32'h42933ff7, 32'hc35b0176},
  {32'h4507901a, 32'h415752bf, 32'h4255b7b8},
  {32'hc4b14e74, 32'h43974246, 32'hc3018727},
  {32'h437ae8a0, 32'hc2f9dfff, 32'hc3f8c852},
  {32'h43837be4, 32'hc3e87740, 32'h4348c59e},
  {32'h44899c86, 32'hc2149b91, 32'hc32d413b},
  {32'hc3febf23, 32'hc40430fe, 32'h4417044c},
  {32'h448da19c, 32'h4256c69a, 32'h43b82092},
  {32'hc4dbaa10, 32'hc10808bc, 32'h42197472},
  {32'h44a79d73, 32'h4300d81a, 32'h43e6ad0d},
  {32'hc5078819, 32'hc31b6ecf, 32'hc39c0aeb},
  {32'h44862b18, 32'h418e39da, 32'hc2a25827},
  {32'hc506cc36, 32'h420937d6, 32'hc39152c1},
  {32'h44c07f21, 32'hc3529a00, 32'h4255356a},
  {32'hc503921e, 32'hc24b6700, 32'hc34be81c},
  {32'h45071503, 32'h416814c1, 32'h4396cb72},
  {32'hc50c8595, 32'hc235e767, 32'h4381960b},
  {32'h4503d65f, 32'h429c9204, 32'hc16692b7},
  {32'h4263a9e2, 32'h439fad95, 32'hc305034a},
  {32'h44e38f25, 32'h43cba89f, 32'h415ea6ee},
  {32'hc3871230, 32'h4379f222, 32'hc321daf7},
  {32'h44ca6148, 32'hc2b05a66, 32'h419723ca},
  {32'h4311fe98, 32'hc2d20e7c, 32'h42cc002f},
  {32'h448b7995, 32'hc2af38d6, 32'h43761b56},
  {32'hc505ca9b, 32'h43882d5a, 32'hc1ef5d5b},
  {32'h448a33d8, 32'hc1d54aa7, 32'h42c9f103},
  {32'hc34b3af7, 32'hc375f811, 32'h4368b224},
  {32'h44d99ad5, 32'hc24daae8, 32'hc2f71f30},
  {32'hc4c04f07, 32'h4373c825, 32'h426f220e},
  {32'h43b1ae2d, 32'h4340c396, 32'h4299d828},
  {32'h43c75180, 32'h435c65f8, 32'h414644dc},
  {32'h44f8fbf8, 32'hc3d11207, 32'h4357ab6e},
  {32'hc2fec5a2, 32'hc3b550da, 32'h40b3fbd3},
  {32'h42fb9960, 32'hc2265ab0, 32'hc3c194b1},
  {32'hc5124a88, 32'h41421f9e, 32'h433938d0},
  {32'h4303b3af, 32'h42a44c9e, 32'h435dcff0},
  {32'hc3169930, 32'h4317f060, 32'hc39a4f8e},
  {32'h442b32ba, 32'h435bac8d, 32'hbe32db48},
  {32'hc4c1c1e1, 32'hc27cafbd, 32'hc26a793e},
  {32'h4514e678, 32'h413c5dd0, 32'h42556b30},
  {32'hc3c7f80d, 32'hc14b61ff, 32'h424861fc},
  {32'h436e3274, 32'hc2dc028b, 32'h43c16c74},
  {32'hc31a3b1d, 32'hc3650a5d, 32'hc364f811},
  {32'h43f318e8, 32'h44079534, 32'h42bb69af},
  {32'hc4fc288c, 32'h42481b93, 32'hc2f4286b},
  {32'h44efefa3, 32'h436e1160, 32'hc393eb09},
  {32'hc4aef82e, 32'hc37fc81b, 32'hc39c549d},
  {32'h43a62c1e, 32'h42fb223a, 32'hc345ad65},
  {32'hc3f4c094, 32'h4004a12a, 32'hc2b2f6df},
  {32'h44628998, 32'hc2ecb61c, 32'hc346526c},
  {32'hc474b1ea, 32'hc3f88f7c, 32'hc3936a6c},
  {32'h44832987, 32'h43598843, 32'h428b0cfa},
  {32'hc49c7bdc, 32'h4206ca4f, 32'h432bcd41},
  {32'h440aa857, 32'h4340184d, 32'hc365d866},
  {32'hc4869fef, 32'hc3aa2a1d, 32'h43543860},
  {32'h4506a853, 32'h43dba473, 32'h421e7dcb},
  {32'hc3d905c6, 32'hc3232647, 32'hc2fcdaab},
  {32'h43716b1c, 32'hc37a459c, 32'h43bbcce7},
  {32'hc50c12fd, 32'hc37a8920, 32'h4378f6b6},
  {32'hc35f6920, 32'h43578c4e, 32'h428d0918},
  {32'hc50c49a2, 32'h429a7175, 32'h43481315},
  {32'h4500a13b, 32'h43380e11, 32'hc31610f1},
  {32'hc3c02e44, 32'hc3c63459, 32'h43266a93},
  {32'h44a6077c, 32'hc274cc61, 32'h42a10720},
  {32'hc48b843e, 32'hc2484e53, 32'hc3a655ff},
  {32'h44b7e092, 32'h41fdf791, 32'hc2e56c55},
  {32'hc47bc598, 32'h41614ba8, 32'h41bbf808},
  {32'h43296cbd, 32'hc215c601, 32'hc39b8f21},
  {32'hc4d8e8c0, 32'hc37b34b2, 32'h42affae3},
  {32'h44843148, 32'h40e0d604, 32'hc388d4ef},
  {32'hc4e734c8, 32'hc315a19a, 32'h42bcc215},
  {32'h42839e30, 32'hc34d9fcf, 32'hc3bc6ea9},
  {32'hc21ca000, 32'h42d58204, 32'h42bfb09a},
  {32'h44ac7c25, 32'h4300c49a, 32'hc31327bc},
  {32'hc4be51d5, 32'h42e875ae, 32'hc2b69ea8},
  {32'h44cd32a8, 32'h4325e6f7, 32'h43319a7b},
  {32'hc088ea00, 32'hc2ff6836, 32'h430d3878},
  {32'h44a6ae2b, 32'hc2331c56, 32'h4208a092},
  {32'hc283a808, 32'hc0e6ed32, 32'hc2af6f14},
  {32'h4436204f, 32'h43b6ae47, 32'hc2f74eb7},
  {32'hc500145b, 32'hc39ae8d4, 32'hc3e0412b},
  {32'h44b712f5, 32'h43c0e9c8, 32'h40e90428},
  {32'hc4a8f5db, 32'h432a6582, 32'hc311808d},
  {32'h44214f60, 32'h41b16472, 32'h43c43f6e},
  {32'h415c9d00, 32'hc30bcc54, 32'hc384a97c},
  {32'h43d66e10, 32'h4289465f, 32'h433b1b25},
  {32'hc3941c7c, 32'h43078963, 32'h43b2a3a2},
  {32'h450af5fe, 32'hc200a092, 32'h4217a0b3},
  {32'hc4bfd932, 32'h4299ae68, 32'h43347d0f},
  {32'h440d9c92, 32'hc20fc7d8, 32'h43bda64f},
  {32'hc416f4d6, 32'hc328a60c, 32'hc2e4c90e},
  {32'h450a8151, 32'hc326ae08, 32'h4204ac6a},
  {32'hc4728971, 32'hc3489c5f, 32'hc2f28d23},
  {32'h414bb728, 32'hc38075c9, 32'h42856ec5},
  {32'hc4fd0eed, 32'hc39d9269, 32'h4381d57a},
  {32'h44dc1292, 32'h42a9b8be, 32'hc26fd235},
  {32'hc51e1b63, 32'h4319888f, 32'hc2df5ea4},
  {32'h451b1538, 32'hc3b5dfb0, 32'hc3c0bb24},
  {32'hc4a1384b, 32'hc2352d0e, 32'hc32da118},
  {32'h44e52ead, 32'h4408c565, 32'h42ba8bde},
  {32'hc34c4c60, 32'hc3cf96f5, 32'hc369db3c},
  {32'h44e550fd, 32'hc0fd26ec, 32'hc3b0415a},
  {32'hc504b1f9, 32'h433cc371, 32'hc3deaa6b},
  {32'h438c293f, 32'hc32b2baa, 32'hc3061362},
  {32'hc4b7dc36, 32'h43c37e8a, 32'h437acb04},
  {32'h4413c902, 32'hc163e91d, 32'h40ff418c},
  {32'hc4b3d488, 32'hc0f35a4a, 32'hc0457534},
  {32'h44a762fb, 32'hc1d624b8, 32'h4325cc7e},
  {32'hc50744df, 32'h43a33404, 32'h4285101a},
  {32'h44873907, 32'h426a7c4c, 32'hc3176f01},
  {32'hc4106a2c, 32'h4329196a, 32'hc367fe9c},
  {32'h44d0d8de, 32'hc2f6dd17, 32'hc3d79a9a},
  {32'hc42880a8, 32'hc3d0207c, 32'hc37a535f},
  {32'h43b55e18, 32'hc2a27560, 32'hc2eebf10},
  {32'hc42c320e, 32'hc3b3e6fc, 32'h43121165},
  {32'h44a3004d, 32'hc3ca017f, 32'h42e1818e},
  {32'hc4228b40, 32'hc34094a3, 32'hc371c3de},
  {32'h44656d4c, 32'h43860a30, 32'h42f906cc},
  {32'hc4c1bf1a, 32'hc3ba3b68, 32'h42c68974},
  {32'h44a499c0, 32'hc2edef92, 32'h428b801e},
  {32'hc4ad506c, 32'h440cdb44, 32'h4287f55a},
  {32'h43ed95ca, 32'h433b0a51, 32'h410555cc},
  {32'hc481ada7, 32'h41c08a96, 32'h436b9ad2},
  {32'h44a19cab, 32'h4332ea9e, 32'h4303bb2c},
  {32'h427c2d50, 32'h42e8779d, 32'hc32fdf06},
  {32'h44bc3435, 32'hc37b55d8, 32'hc389e540},
  {32'hc5028bb9, 32'h4331c6ac, 32'hc2b5453b},
  {32'h45014468, 32'h427a20e6, 32'hc2dac686},
  {32'hc513d12c, 32'hc270f275, 32'hc38bef8f},
  {32'h43afd627, 32'hc2954b8a, 32'hc1a1f4a4},
  {32'hc4d89b44, 32'hc332e4a1, 32'hc36a4d7e},
  {32'h44ef1ca7, 32'h43a85e17, 32'h42bc6d17},
  {32'hc2cf0e10, 32'h42c315e2, 32'hc2cd87d7},
  {32'h44e489d8, 32'h439b54bf, 32'h43287d9e},
  {32'hc515bd4b, 32'h4402b0c1, 32'h42a40ff8},
  {32'h4426fd77, 32'hc2ac73d7, 32'hc286e58a},
  {32'hc3d24e38, 32'h428d440b, 32'hc350156c},
  {32'h44f69d29, 32'h43d7a534, 32'h438367f0},
  {32'hc443d7e8, 32'hc329dd21, 32'hc33c5391},
  {32'h45106f2a, 32'h439b05b7, 32'h43c1983e},
  {32'hc3050448, 32'h438a3ca0, 32'h4329111f},
  {32'h44e20f0e, 32'hc3a7924b, 32'h430d084e},
  {32'hc2f8f5d8, 32'h42304035, 32'hc3999acc},
  {32'h44eb5a1e, 32'hc3a0a610, 32'hc34ab881},
  {32'hc4a4b78d, 32'h4401d013, 32'h41b81866},
  {32'h452062de, 32'hc3b99c61, 32'h43894d74},
  {32'hc505b659, 32'h435b66c2, 32'h42b9b261},
  {32'h445c9468, 32'h4322bc50, 32'h435ba797},
  {32'hc48178d0, 32'h42676f0f, 32'hc3789341},
  {32'h44b3cbc9, 32'hc2cbd32a, 32'h4308d769},
  {32'hc390d9bb, 32'hc3b29e61, 32'h4343bd6b},
  {32'h4432410a, 32'hc1a066e2, 32'hc2c47d35},
  {32'hc4cb7dee, 32'hc393c572, 32'h44009c8a},
  {32'h44a9129d, 32'h4359e04a, 32'h437b58fc},
  {32'hc4010c4a, 32'hc3a7e9a7, 32'hc2c60982},
  {32'h449b4678, 32'h43167c96, 32'hc387ff0f},
  {32'hc3b1fe4b, 32'hc3957e85, 32'h4241de74},
  {32'h449ec52f, 32'h43a17d8c, 32'h4337ed1f},
  {32'hc49315e8, 32'hc26dffd9, 32'hc1df42f2},
  {32'h440ae638, 32'hc35fce9a, 32'h436d7b57},
  {32'hc3f6f23e, 32'hc3792de8, 32'h432aaf65},
  {32'h44984e55, 32'hc2803e71, 32'hc36729cb},
  {32'hc4b1ba26, 32'hc40ec49e, 32'hc0c6280b},
  {32'h44b58d2a, 32'hc3f82614, 32'h4388e216},
  {32'h44763cc0, 32'h436e3a80, 32'hc27fae6e},
  {32'hc5118388, 32'hc34ff5b9, 32'hc279a95c},
  {32'h44f544f2, 32'h433eda9f, 32'hc2e3fbc4},
  {32'hc48ce265, 32'h4357acec, 32'h43433f2e},
  {32'h4444ed5a, 32'hc2d9648a, 32'hc2a8209e},
  {32'hc50db61a, 32'hc3507717, 32'h43dc6c67},
  {32'h450bc54c, 32'hc3aeb3a8, 32'h427fda3f},
  {32'h420362cc, 32'hc2d45eee, 32'hc35356a1},
  {32'h44e121dd, 32'hc1af23c3, 32'h437d8240},
  {32'hc4f42f8f, 32'hc3950bec, 32'h4386d1c0},
  {32'h4347d6b2, 32'h42bc33dd, 32'hc26e35ff},
  {32'hc4d85dc0, 32'hc231d57d, 32'hc1f213b1},
  {32'h448276dc, 32'h42859e16, 32'hc37f4b47},
  {32'hc4cfa132, 32'h43413d29, 32'hc3873f21},
  {32'h4501d90e, 32'h44025e7c, 32'hc31da3cd},
  {32'hc3e1435c, 32'hc3961146, 32'h4285ecbb},
  {32'h44e369b8, 32'h429d80ab, 32'hc38a7220},
  {32'hc5138bdc, 32'h436c649a, 32'hc37ace97},
  {32'h446c4db8, 32'hc2abe8ea, 32'hc2ad40b1},
  {32'hc503985a, 32'h43107be8, 32'hc31a44fc},
  {32'h44ff51e3, 32'hc35778cf, 32'h42c536ba},
  {32'hc507c90a, 32'h43522c2b, 32'h413c8943},
  {32'h451aa9d2, 32'hc3438add, 32'h42355564},
  {32'hc4e6bc1c, 32'h43fcf9d8, 32'h4146484c},
  {32'h44a45796, 32'h431a7be7, 32'h4233e914},
  {32'hc4fafe41, 32'hc2a865ae, 32'h43450b0a},
  {32'h44587a2f, 32'h42a6dc30, 32'h43165589},
  {32'hc4da5d3a, 32'h43829083, 32'h4336de6c},
  {32'h43b46034, 32'hc379c652, 32'h4343d7bf},
  {32'hc484ee13, 32'hc087dcd8, 32'hc31b83f3},
  {32'h4504a9d3, 32'hc3979506, 32'hc3be2c58},
  {32'hc4a75208, 32'h4309b656, 32'h42d821c2},
  {32'h44af4893, 32'hc23f55dc, 32'hc2d8b939},
  {32'hc3b8a070, 32'h43cfba2b, 32'h430be1b8},
  {32'h451194d8, 32'h429c43bf, 32'hc3863f37},
  {32'hc4f3c576, 32'hc3152c36, 32'h430df1ff},
  {32'h444ce902, 32'h42bf822f, 32'h439bccee},
  {32'hc4ba8fec, 32'h4199cec0, 32'h43636d84},
  {32'h446349ee, 32'h4302566e, 32'h4332335e},
  {32'hc47732e0, 32'hc3220276, 32'h43353059},
  {32'h45076944, 32'h43f15301, 32'h417fd657},
  {32'hc4ef9668, 32'hc36fe4cb, 32'h41919ebb},
  {32'h444d8b1c, 32'h4374d24e, 32'hc31edb7a},
  {32'hc4fd2e33, 32'h42be7bbb, 32'hc3277a2a},
  {32'h44f11fa6, 32'hc3e85b17, 32'hc3008e96},
  {32'hc4f0386e, 32'hc2acb9b5, 32'hc3e2ebb2},
  {32'h449e19fa, 32'h418c3d09, 32'hc3590837},
  {32'hc49bf1a0, 32'h4330478a, 32'hc30c045e},
  {32'h44e00149, 32'h43e04d81, 32'hc3369d94},
  {32'hc5010b4e, 32'h42b5791f, 32'hc268f8b5},
  {32'h439fccc0, 32'hc2cfa546, 32'h42b95880},
  {32'hc3589c38, 32'h429ccec7, 32'h43100389},
  {32'h44eb3b5c, 32'h43e18ffd, 32'h429effa3},
  {32'hc49ec772, 32'h4312884d, 32'hc344c14d},
  {32'h44fbcf0b, 32'hc32c049b, 32'hc344e906},
  {32'hc411c248, 32'h42553105, 32'h4415ea32},
  {32'h44fb715d, 32'hc3b20f73, 32'hc346fc7f},
  {32'hc4f368d7, 32'h4392ebb2, 32'hc1166b11},
  {32'hc4b5b272, 32'hc18cf575, 32'hc3ecbacc},
  {32'h44c3ddfd, 32'hc39a61ad, 32'hc3c6b336},
  {32'hc4c153ea, 32'hc02b848c, 32'hc35f8766},
  {32'h44be339a, 32'h4325e622, 32'h43ab9291},
  {32'hc400f7ff, 32'h42f6cdbb, 32'hc3299ee1},
  {32'h440cfc3e, 32'hc3af6c93, 32'hc33901db},
  {32'hc4fc11d8, 32'h43035978, 32'hc3c0082f},
  {32'h44c01986, 32'h419768c9, 32'hc24da1ea},
  {32'h429a35d3, 32'h42f1c476, 32'hc3844802},
  {32'h44f6df57, 32'h4296d657, 32'h42aa8353},
  {32'hc499ccfd, 32'hc34800db, 32'h42cbdb7b},
  {32'h4496b415, 32'hc359a9e8, 32'hc1f62efd},
  {32'hc4e29c94, 32'hc220abe3, 32'h4330f4da},
  {32'h441009b8, 32'h43f1b4ce, 32'hc34f808e},
  {32'hc3b4648c, 32'h42d5935f, 32'h434d7191},
  {32'h450e5de3, 32'hc2b4462c, 32'hc3e97625},
  {32'hc43449da, 32'h43693c9a, 32'hc27f3702},
  {32'h4506d957, 32'hc3165cbe, 32'hc397b764},
  {32'hc2885114, 32'h4358597a, 32'h4378aa56},
  {32'h44fcc23f, 32'h42d59e79, 32'hc344a648},
  {32'hc4fe5d56, 32'h42ea9a37, 32'h4375570d},
  {32'h443c5c06, 32'hc3832864, 32'h43575c05},
  {32'hc3f24868, 32'hc25607b4, 32'h431a3abb},
  {32'h4453f776, 32'hc3775994, 32'hc38c970a},
  {32'hc429c692, 32'h4308beb1, 32'h42df716d},
  {32'h44ea5612, 32'h41c7e38d, 32'h430ccce9},
  {32'hc469794c, 32'h42654470, 32'hc29f177a},
  {32'h44e60c88, 32'hc357eafc, 32'hc3480bbf},
  {32'hc4dd4f21, 32'h4386b383, 32'h431942f3},
  {32'h44d9d644, 32'hc3b691ee, 32'h439ceed6},
  {32'hc4a0f085, 32'hc330c0b3, 32'hc2e4a040},
  {32'h45091fa5, 32'hc3d182f3, 32'hc39776b8},
  {32'h43356c8c, 32'hc32086f8, 32'h43345bb7},
  {32'hc3bf4e6f, 32'h427f3fd1, 32'h430e461e},
  {32'h44c5aa70, 32'h4331642f, 32'hc26d0f8d},
  {32'hc2a6b9be, 32'h4397524e, 32'h437d5fc5},
  {32'h448d9ccf, 32'hc3851de0, 32'hc2967ab1},
  {32'hc48dd802, 32'h42b1f446, 32'h42de3c8c},
  {32'h4328874c, 32'hc33edd44, 32'hc37b4e1b},
  {32'hc49a6c63, 32'hc390844e, 32'h429ebb57},
  {32'h44d67142, 32'h41e40d66, 32'h4338e31b},
  {32'hc4be8eda, 32'hc23781e2, 32'hc3569ba2},
  {32'h447f07be, 32'hc3539a3b, 32'hc2890748},
  {32'hc3b250a0, 32'hc3a28bed, 32'h42acf6b2},
  {32'h4457c908, 32'hc1b70802, 32'h417f0fea},
  {32'hc4d8eefb, 32'hc320a7f8, 32'h4205cb27},
  {32'h43e01e64, 32'h4225eacb, 32'hc351b52b},
  {32'hc4d06854, 32'hc3bce706, 32'hc24e63df},
  {32'h44b70535, 32'h42d6f422, 32'h42c45ced},
  {32'h431725a8, 32'hc3b466d5, 32'h43209547},
  {32'h44a675f3, 32'h43bd40e9, 32'h4311e8bb},
  {32'hc46a841c, 32'hc3b34dbb, 32'hc31b9797},
  {32'h44fb749d, 32'h4412c2b3, 32'hc1b1e550},
  {32'hc4bf9e3b, 32'hc30467b8, 32'h437402f1},
  {32'h440761ce, 32'h42dd31d5, 32'h4309d383},
  {32'hc3f36882, 32'h43732de6, 32'hc2d85717},
  {32'h452adad8, 32'h43db93ed, 32'h437a1c57},
  {32'hc3b5b671, 32'hc3912037, 32'hc33ca39a},
  {32'h44363008, 32'h4312bd50, 32'h42897ed4},
  {32'hc4335b8d, 32'hc284626e, 32'hc2dcbf0d},
  {32'h44f8e0e4, 32'h435a0768, 32'hc34145f3},
  {32'hc3bfea80, 32'hc320f9b6, 32'hc3423b30},
  {32'h431f3dc0, 32'hc2ba2dc9, 32'hc387aac9},
  {32'hc4a3d4d7, 32'hc1fd4d8d, 32'hc31ef6c6},
  {32'h44e91b44, 32'h43c57915, 32'h43941a7a},
  {32'hc41ee9fc, 32'hc23ce6e6, 32'hc3638b7f},
  {32'h4305fde0, 32'hc2d2b6d5, 32'hc334b69b},
  {32'hc4ab5b17, 32'hc35b5ef9, 32'h42a69ae2},
  {32'h44a0afcf, 32'hc3bf619f, 32'hc21a2851},
  {32'hc4803fb2, 32'h4236c34f, 32'hc414047b},
  {32'h430ebee0, 32'hc2c4ed10, 32'h4396a6ab},
  {32'hc4d2c403, 32'h42fd0936, 32'h4381a36d},
  {32'h44d7f65a, 32'h4216d78e, 32'h436f6537},
  {32'hc4906f15, 32'h4248bb96, 32'h43d0ca4e},
  {32'h442ab1b4, 32'h41ac1fcb, 32'h4369b205},
  {32'hc517fb44, 32'h433870a9, 32'h42a635b2},
  {32'h448d038e, 32'h434a2e20, 32'h42f6f019},
  {32'hc356984b, 32'h4329d173, 32'h4281515e},
  {32'h44af9af1, 32'h4217c71a, 32'h42798444},
  {32'hc4c3303a, 32'h3f9ff8ca, 32'h429affd9},
  {32'h44e64eb5, 32'h43340072, 32'hc3427f6a},
  {32'hc4026680, 32'hc2f85d93, 32'h42a4f5a7},
  {32'h4310451c, 32'h427c300c, 32'h43687f4b},
  {32'hc4e55d80, 32'hc32e86d8, 32'hc386113e},
  {32'h442c1a55, 32'hc2ee50ac, 32'h41337275},
  {32'hc4cd5b98, 32'hc165dc90, 32'h431a467c},
  {32'h4402585c, 32'h43358178, 32'hc067a79b},
  {32'hc4691564, 32'hc26ce39b, 32'h4376f101},
  {32'h4412e12f, 32'h43919633, 32'hc0da9068},
  {32'hc30bbc80, 32'hc37ffb1c, 32'hc2a5482d},
  {32'h43a3aa53, 32'h43487931, 32'hc2ab1acb},
  {32'hc493767f, 32'hc04cd733, 32'h4149072d},
  {32'h43fcdb90, 32'hc4099341, 32'h430ee69b},
  {32'hc3f47be0, 32'hbfda0320, 32'hc14f51ce},
  {32'h440b37a7, 32'hc1ce953a, 32'h423e7de2},
  {32'hc499f0cf, 32'h4350cf38, 32'hc0c4c45c},
  {32'h45100482, 32'hc2f7407c, 32'h43072048},
  {32'hc21b43f7, 32'h42f8d513, 32'hc3a60621},
  {32'h4502c4eb, 32'h4295e9a4, 32'hc3a619e5},
  {32'hc3e051d4, 32'hc29ccae6, 32'hc36588c1},
  {32'h447f65f4, 32'h43fcbfa0, 32'h436fcc59},
  {32'hc4a7be2b, 32'hc223ec53, 32'h438f9564},
  {32'h4507d24e, 32'hc3292772, 32'h4392847d},
  {32'hc40cdc16, 32'hc2ea5551, 32'h436f8215},
  {32'h4434f016, 32'hc3fbdcb2, 32'hc38787ae},
  {32'hc4029249, 32'h42ec1c17, 32'hc3360c42},
  {32'hc2ea3004, 32'hc2fa5ec5, 32'hc39668da},
  {32'hc4a15357, 32'hc30d3ec2, 32'h427ff73c},
  {32'h44c88607, 32'hc192e794, 32'hc36dfb26},
  {32'hc5006bb3, 32'hc3265f50, 32'h4242ec6d},
  {32'h4475256d, 32'h43541e01, 32'hc3025b54},
  {32'hc30029b7, 32'hc37ee1a7, 32'hc1fb54c3},
  {32'h44885ecc, 32'hc339c19c, 32'h434dbca9},
  {32'hc3a94e50, 32'h4342ff9b, 32'hc21dcde8},
  {32'h44edc630, 32'hc296a628, 32'hc3eee150},
  {32'hc4edfb78, 32'h426f922a, 32'hc3175171},
  {32'h446bbef4, 32'hbfd94680, 32'hc2880db6},
  {32'hc5076b99, 32'h436b5b54, 32'h4209c00d},
  {32'h4460fd3c, 32'hc22b0b0f, 32'h43103297},
  {32'hc46aeb28, 32'h424c3f11, 32'hc30e9ccf},
  {32'h442a79f3, 32'h42ff4939, 32'h435677c1},
  {32'hc50d2297, 32'hc33a56ab, 32'h43018491},
  {32'hc476fc9e, 32'hc23ceb34, 32'h43658664},
  {32'h43a73450, 32'h4354fe93, 32'h427b6bf1},
  {32'hc4984107, 32'h429f6bc6, 32'hc349ad4b},
  {32'h43751278, 32'h3efc9e38, 32'h42937593},
  {32'hc4decbef, 32'h4189c049, 32'h43a77774},
  {32'h44fab94a, 32'h4293c23e, 32'hc399a092},
  {32'hc3bfb83e, 32'hc3096cd4, 32'h429790e9},
  {32'h43e128b4, 32'h41ee8a83, 32'hc35f50af},
  {32'hc29ebb40, 32'hc32fe793, 32'hc2b58710},
  {32'h439bf8c4, 32'h430c6420, 32'h43827d5b},
  {32'hc4e5a193, 32'h43137492, 32'h4349722f},
  {32'h44ce586e, 32'hc3a0d3d8, 32'h42eec63e},
  {32'hc4e8ac9a, 32'h4282d591, 32'h430c1bd5},
  {32'h4483a299, 32'hc425ffd0, 32'h41e04b3b},
  {32'hc31b5a28, 32'h4321900b, 32'hc381a31b},
  {32'h436dd748, 32'hc2bf30ab, 32'h42683e21},
  {32'hc4809a07, 32'hc2fb268e, 32'hc34aeb57},
  {32'h4404c3a2, 32'hc2d27112, 32'h43150559},
  {32'hc3cdcf78, 32'h43377b70, 32'h426bed6d},
  {32'h44e92c44, 32'h42ff628d, 32'hc38d6722},
  {32'hc4251475, 32'h42b3e471, 32'h438a2a71},
  {32'h44a9b15a, 32'hc3e7a9b7, 32'hc34055a0},
  {32'hc403e8a4, 32'hc3ec359c, 32'h42494808},
  {32'h44b1bb93, 32'h41f8440d, 32'hc2e66892},
  {32'hc48cb4a7, 32'hc3040ce9, 32'hc34711b6},
  {32'h433221e0, 32'h4408ef3c, 32'hc28735c7},
  {32'hc4e06a33, 32'h4323d25e, 32'h43b09d04},
  {32'h44617964, 32'h43e94311, 32'h43c6d132},
  {32'hc4a089d7, 32'h43082e72, 32'hc331b434},
  {32'h4399c810, 32'h41ff87dc, 32'h4322f098},
  {32'hc2a2db88, 32'h434e5869, 32'hc235c179},
  {32'h445cca3c, 32'h41ee82ec, 32'h43ae2137},
  {32'hc4fc93ea, 32'h43db2e4a, 32'h4298581c},
  {32'h441e53dc, 32'h40e55d31, 32'hc3080749},
  {32'hc4c6742a, 32'h43868d26, 32'h422eb00c},
  {32'h44f8ec22, 32'hc3373e9f, 32'hc3562dc0},
  {32'hc4b41333, 32'hc26d055a, 32'h428f1103},
  {32'h4497488c, 32'hc2a2d2ac, 32'h42a7e537},
  {32'hc4f35444, 32'hc2d0e5ce, 32'h4394e8c8},
  {32'h449b8fba, 32'hc34765dd, 32'h43bec7d0},
  {32'hc451edc9, 32'h4317dac4, 32'h4305caa4},
  {32'h44fe8f5d, 32'h4338d693, 32'h42a52ffa},
  {32'h42b6b4c0, 32'h408302f4, 32'hc342bc85},
  {32'h443fe4ae, 32'hc2cad443, 32'h43b82ade},
  {32'hc481acdc, 32'hc010129f, 32'h424c71a4},
  {32'h44c6573e, 32'h4334722b, 32'hc1ead3ce},
  {32'hc31aaa2a, 32'hc40d9c09, 32'h435083cf},
  {32'h44fcc758, 32'h4371b631, 32'hc194e329},
  {32'hc376864e, 32'h42c959af, 32'h438b14b8},
  {32'h44e2f8ee, 32'hc38d21b5, 32'hc33316d0},
  {32'hc4e25bfd, 32'h432d2209, 32'h435cb601},
  {32'h4042bb00, 32'h439b3933, 32'h43708f26},
  {32'hc4cb9310, 32'h43460833, 32'hc2a9a410},
  {32'hc1c99890, 32'hc331689f, 32'h43704f0d},
  {32'hc4e69a13, 32'h43339f6c, 32'h417a89fb},
  {32'h43c0609f, 32'hc231c5fb, 32'h42d58a11},
  {32'hc400cf5a, 32'h411250bd, 32'hc3b7b48c},
  {32'h44a55830, 32'hc2821fc4, 32'h43e95336},
  {32'hc4283186, 32'h43a7d790, 32'hc1a6a45a},
  {32'h44fb9f9a, 32'hc35363ec, 32'h439d5d20},
  {32'hc4a630f0, 32'hc2fc5a02, 32'h42a0e5e3},
  {32'h43fe4ece, 32'hc313d8be, 32'hc2ce2060},
  {32'hc48bc695, 32'hc3dbee38, 32'h420320eb},
  {32'h443770c7, 32'h434ee431, 32'h438f08cf},
  {32'hc4a33911, 32'h42e10eac, 32'hc102d66f},
  {32'h44e1bf99, 32'h4267aa21, 32'hc34bd3cf},
  {32'hc492a55d, 32'h4235bc4a, 32'hc3aafbc8},
  {32'h44535a86, 32'h42477f95, 32'hc347b27e},
  {32'hc39d8728, 32'h4182c270, 32'h4384167f},
  {32'h43192e44, 32'hc3204441, 32'hc2f87242},
  {32'hc3bb7c88, 32'hc233072c, 32'h42e0625f},
  {32'h44e6055c, 32'h4209e34d, 32'h4214536c},
  {32'hc4f809cc, 32'hc27d4324, 32'h43f283c8},
  {32'h43192f20, 32'hc413985b, 32'h43f6fc6c},
  {32'hc37202dc, 32'hc259836f, 32'h41eafef3},
  {32'h44751fcc, 32'h42c7ecc3, 32'hc1c2c4ba},
  {32'hc4d02b5c, 32'h41e0702c, 32'hc378c443},
  {32'h44d75011, 32'hc3ad7fd8, 32'h4373c81b},
  {32'h403d0f60, 32'h429a832f, 32'hc2186d5d},
  {32'h44b80c0d, 32'h43135e95, 32'hc25e5a23},
  {32'hc36ef950, 32'h42b016fc, 32'h42c4c305},
  {32'h450bb09c, 32'h42e841ad, 32'h433ba3dd},
  {32'hc4ffb665, 32'hc325c0fb, 32'hc37181be},
  {32'h446f370e, 32'h42759204, 32'hc22b385b},
  {32'hc487464f, 32'h43992a3e, 32'h428bb27f},
  {32'h44855ea4, 32'hc2c0c251, 32'h431735c8},
  {32'hc4fa8820, 32'hc3453e19, 32'h4356072a},
  {32'hc012ea00, 32'h42ee9c15, 32'hc3258b09},
  {32'hc50eb7c9, 32'hc356670e, 32'h430b9634},
  {32'h43e578e8, 32'hc382b622, 32'hc32274ff},
  {32'hc47b0ede, 32'h3edd40d0, 32'hc2df7f29},
  {32'h44893bc4, 32'h43892d64, 32'hc2f18412},
  {32'hc49a973c, 32'h42aa891a, 32'h426e2642},
  {32'h44453986, 32'hc2f1ce0e, 32'hc31db691},
  {32'hc4205a22, 32'h42cefe68, 32'hc322944f},
  {32'h44948fee, 32'h43c5e555, 32'h42bfe7e5},
  {32'hc50dd8cc, 32'h431681f8, 32'h42e1bf09},
  {32'h44ea9e8c, 32'hc37319e1, 32'hc3ad567b},
  {32'hc51c557c, 32'hc2c0f6e2, 32'h436747b2},
  {32'h44867069, 32'hc364014d, 32'h43b4244d},
  {32'hc4992a04, 32'hc2b80a5d, 32'h42e15675},
  {32'h443944ff, 32'h435a00b4, 32'hc38545b8},
  {32'hc3ce8eca, 32'hc2eb7b04, 32'h4308fd08},
  {32'h43ea941a, 32'hc1d3add6, 32'h42b51bdd},
  {32'hc4d2f396, 32'hc3a171b5, 32'hc2db83b0},
  {32'h43ba0554, 32'hc2371b0d, 32'h406072d7},
  {32'hc48a0e0d, 32'hc3cdd9f5, 32'hc3988801},
  {32'h4464df60, 32'h42e91b01, 32'h436f5ebf},
  {32'hc3941bac, 32'hc3228150, 32'h41e5d738},
  {32'h452215a5, 32'hc38d7d7e, 32'hc1b165c2},
  {32'hc50fa5d7, 32'hc362a72a, 32'h438537fa},
  {32'h43335cd0, 32'hc34cf48f, 32'h4023efae},
  {32'hc49a4475, 32'hc14b4394, 32'h435f0638},
  {32'h450ab256, 32'hc3ab120c, 32'h44192106},
  {32'hc333d3c8, 32'h423d83ba, 32'h42c09f09},
  {32'h45135f33, 32'hc3100fc4, 32'h43a10c7b},
  {32'hc3ad26e4, 32'hc30d201d, 32'hc3e3e65a},
  {32'h44759b54, 32'h430b5b17, 32'h41fe1106},
  {32'hc524a98a, 32'hc332adf1, 32'h41704cb7},
  {32'h449424a3, 32'h42b1921f, 32'hc279d456},
  {32'hc491a66d, 32'hc327877c, 32'h43a57e20},
  {32'h43ffcda8, 32'h43a43b0f, 32'h434ca72b},
  {32'hc4c07058, 32'hc32d26b9, 32'h429e9ffc},
  {32'h45091cd0, 32'h43af2ba2, 32'hc3288c45},
  {32'hc4c85259, 32'h428adebe, 32'hc39f971e},
  {32'h44e7767b, 32'hc380e9d4, 32'hc2594c02},
  {32'hc4831540, 32'hc294c186, 32'h43abf4cc},
  {32'h450a4d3b, 32'hc38da298, 32'h427f9549},
  {32'hc4ff9f24, 32'h43137acd, 32'h434680d8},
  {32'h43979f6a, 32'hc3756f78, 32'hc2371eb5},
  {32'hc4a329e6, 32'hc211a567, 32'h42903926},
  {32'h44d57315, 32'h41bc6525, 32'h4312947e},
  {32'hc422ff28, 32'hc201a84a, 32'hc32ccc03},
  {32'h44969699, 32'hc3b9c7b8, 32'h4374fb29},
  {32'hc40c9044, 32'h430d26c7, 32'hbfd36fe5},
  {32'h444de1d3, 32'h432c016e, 32'hc11f0ee1},
  {32'hc5054fa1, 32'hc2bb61d4, 32'hc39264da},
  {32'h449e0bec, 32'hc3276648, 32'h42b66d0d},
  {32'h42750cc0, 32'hc3209743, 32'hc0fdd514},
  {32'h442a1714, 32'h4134188d, 32'h42305877},
  {32'hc4551cb0, 32'hc2c061fc, 32'h41d82815},
  {32'h43bf9122, 32'hc3037983, 32'hc36b10db},
  {32'hc49a298a, 32'hc367a0ca, 32'hc332e5f0},
  {32'h451a0d26, 32'hc380db38, 32'hc30d09fa},
  {32'hc48194b7, 32'hc356a72c, 32'hc37dd0f2},
  {32'h44af65c6, 32'h43e179dc, 32'hc2695956},
  {32'hc4b30102, 32'h43a58dea, 32'h41879796},
  {32'h44954e79, 32'h3f10f798, 32'hc3a73550},
  {32'hc4be0e12, 32'h436ff715, 32'h42eeb921},
  {32'h44ff441f, 32'h4401a34d, 32'hc43c11cb},
  {32'hc3f8a70c, 32'h420e5c33, 32'hc2ed8c40},
  {32'h449fb7d8, 32'hc3502e9a, 32'h4299e260},
  {32'hc37bb845, 32'h425d99b3, 32'h4394df48},
  {32'h44bf705c, 32'h430f8dc8, 32'hc3ca1768},
  {32'hc4ea2bd7, 32'hc38f3b14, 32'h41a6570b},
  {32'h418e0840, 32'hc301ae9a, 32'h43a64cf4},
  {32'hc4e6488b, 32'hc36b8325, 32'hc1ebb79f},
  {32'h440b6e6d, 32'h42916950, 32'h43e0b7b0},
  {32'hc4059f52, 32'hc31f6e71, 32'h425bec34},
  {32'h4419deb4, 32'hc1e88855, 32'h4167c98a},
  {32'hc50547c0, 32'h426c2b53, 32'hc27e53a8},
  {32'h449fa0fc, 32'hc3314ceb, 32'hc32e502c},
  {32'hc3ef6676, 32'h4341a94e, 32'h4366d89f},
  {32'h446c065c, 32'hc270a071, 32'hc0a09a71},
  {32'hc3fc040b, 32'h4195ac67, 32'hc3ccefeb},
  {32'h442035ba, 32'hc20fa8c5, 32'h42dc2df7},
  {32'hc3e88754, 32'h433e0e67, 32'hc353ac11},
  {32'h44dcc7c9, 32'hc38c2cad, 32'hc3248640},
  {32'hc3e3644c, 32'hc3c9b50d, 32'h4337a9ff},
  {32'h44912f04, 32'h42eaf904, 32'hc324ea53},
  {32'hc3e99410, 32'h41b34496, 32'h43965f65},
  {32'h44c87812, 32'h41643a8b, 32'hc371d8ad},
  {32'hc514c9dc, 32'h415c30b9, 32'hc1bec41c},
  {32'h451b3bed, 32'hc29fc5b6, 32'h43c7db51},
  {32'hc4af1fd2, 32'hc2c378a0, 32'h416169d1},
  {32'h45263c1f, 32'h43b84c22, 32'h4315c681},
  {32'hc4406488, 32'h43f414a8, 32'h42fc1588},
  {32'h4499026f, 32'h43d10923, 32'h43495d27},
  {32'hc4b95fb7, 32'hc20a9a28, 32'hc0fbe0c4},
  {32'h44d94865, 32'hc2233cc5, 32'hc3864923},
  {32'hc48fc8ee, 32'h4415ed20, 32'h4416c4a9},
  {32'h44892cb2, 32'hc26e6d70, 32'hc2cc1e95},
  {32'hc504bdbf, 32'h42431e46, 32'hc340e067},
  {32'h45099494, 32'hc20fb02f, 32'hc38426da},
  {32'hc512b719, 32'hc0c87b48, 32'h4267cf2a},
  {32'h44deb73a, 32'hc32430c7, 32'h4384a39b},
  {32'hc3fd01e0, 32'hc3075680, 32'hc3800863},
  {32'h44c46684, 32'h42a6dd2c, 32'h438e0d91},
  {32'h430c7d61, 32'hc38f1927, 32'h436b7360},
  {32'h440124e4, 32'h436cd400, 32'h424d5ce1},
  {32'hc512caf8, 32'h425a51fa, 32'h4399c986},
  {32'h4434889a, 32'hc3685ba0, 32'hc2cdd817},
  {32'hc4fc02a5, 32'hc335e519, 32'hc2ce2572},
  {32'h441cc6a6, 32'hc15c6d41, 32'h41704f7a},
  {32'hc43cd2fc, 32'hc329b070, 32'h4409059a},
  {32'h41a5d560, 32'h428c4b8f, 32'hc28f56da},
  {32'hc4f73b05, 32'h4183626f, 32'h43933b63},
  {32'h449f452b, 32'hc2acaece, 32'hc2cef4e0},
  {32'hc2ddc808, 32'hc2ea051a, 32'h42c41655},
  {32'h446349ce, 32'h42e4b7b9, 32'hc31fbe41},
  {32'hc4add8b6, 32'h4416c9dc, 32'h42f057b0},
  {32'h44aec3ec, 32'hc37f0ed7, 32'hc1a3f60e},
  {32'hc46d6cd6, 32'hc3131924, 32'hc34fe4d7},
  {32'h44d21f8c, 32'hc38f2937, 32'h43a8a046},
  {32'hc488dda2, 32'hc30a7830, 32'hc22d3eae},
  {32'h450668b3, 32'hc37ea099, 32'h429d0502},
  {32'hc47a6cf4, 32'h42912036, 32'h4367db9b},
  {32'h44cfcb0a, 32'h43a13c76, 32'hc270909b},
  {32'hc495b87b, 32'hc3966f92, 32'hc38381aa},
  {32'h43943169, 32'h435b14a2, 32'hc328cf3c},
  {32'hc37f3f40, 32'h42935f93, 32'hc2b15bfd},
  {32'h44dc895b, 32'h4216884d, 32'hc368ae98},
  {32'hc512a9a5, 32'h433bcb5b, 32'hc3aec795},
  {32'h43a893c5, 32'hc0fc4909, 32'h4288ea38},
  {32'hc50cf7ad, 32'hc39036ae, 32'h42c72164},
  {32'h451f387c, 32'h4393afeb, 32'hc3e1d53b},
  {32'hc4cd0b00, 32'hc22da7ba, 32'hc2849f0e},
  {32'h444559fa, 32'h41953171, 32'h4380b3e9},
  {32'hc43724f3, 32'h43909429, 32'h42ffc346},
  {32'h44dc2bf2, 32'hc0f22daa, 32'h43051de9},
  {32'hc3fc8fdc, 32'h42f36667, 32'h41b54ac2},
  {32'h451b9a07, 32'h41b00cd5, 32'hc206ae25},
  {32'hc3f05c7d, 32'hc390dc7c, 32'hc2ed91ae},
  {32'h44b1e798, 32'h414f9e90, 32'hc34ab362},
  {32'hc4838b44, 32'hc3761316, 32'h420a44a8},
  {32'h4427896a, 32'hc3538a38, 32'h430b1aca},
  {32'hc4aa8992, 32'h41f7cfda, 32'h4373e13f},
  {32'h450911cc, 32'hc28375f6, 32'hc2f72a8f},
  {32'hc45cf132, 32'hc36eb6bf, 32'hc2b8adf6},
  {32'h44e53dbf, 32'hc302a225, 32'h43d524e9},
  {32'hc5148c6e, 32'hc147707a, 32'hc32cfd52},
  {32'h446acb4c, 32'h4306c7fe, 32'hc179b9ca},
  {32'hc31c5fa4, 32'h440879e3, 32'h423677a5},
  {32'h449ba2da, 32'hc22963b4, 32'h429892f3},
  {32'hc4d66385, 32'hc3140c7a, 32'h42cae0e6},
  {32'h4421462a, 32'hc3941d48, 32'hc35e8001},
  {32'hc490ea0a, 32'hbe29e3c0, 32'h43b4444d},
  {32'hc44888c5, 32'h43d893bd, 32'h41f6b898},
  {32'h44c92be0, 32'h42395f66, 32'h42c6678c},
  {32'hc41041d0, 32'hc18938a4, 32'h438ec3c6},
  {32'h442418a6, 32'hc363abcd, 32'hc3666fd5},
  {32'hc3981d2e, 32'h43a0ffd5, 32'h42b85e36},
  {32'h44c79bd8, 32'hc39fd174, 32'h4204dd05},
  {32'hc503e6d2, 32'hc1b1faab, 32'h416ede78},
  {32'h44649f50, 32'h435ffa3f, 32'h41f44f0e},
  {32'hc4a5f4b2, 32'hc28a1e11, 32'hc281d179},
  {32'h4418df38, 32'h42d2d936, 32'hc2bd0ae6},
  {32'hc344bea0, 32'h428f0e04, 32'hc21b4662},
  {32'h451ed0e1, 32'h438268a9, 32'hc30e04db},
  {32'hc4a49426, 32'h42f94169, 32'hc380bd84},
  {32'h4445c917, 32'h427ba07c, 32'h42eae619},
  {32'hc4eb0dad, 32'h42c8540c, 32'h437c1ff6},
  {32'h450cdae0, 32'h439af6dd, 32'h41eefe8d},
  {32'hc4fb832d, 32'hc25f02b9, 32'h4325c4e7},
  {32'h44fc5a65, 32'h43cf9c51, 32'h42ac359b},
  {32'hc4865906, 32'h41de98e2, 32'hc216eca3},
  {32'h4511d61b, 32'hc3d181e7, 32'h42a10ee5},
  {32'hc50f2370, 32'hc3af315c, 32'h43821d47},
  {32'h44e4f1cc, 32'hc321f3e1, 32'hc3cc7d31},
  {32'hc4fdf8ed, 32'hc287cea7, 32'h4317016e},
  {32'h44a8b967, 32'h418f9025, 32'hc12ac11b},
  {32'hc4f5c95a, 32'hc34d236d, 32'hc2bf789d},
  {32'h44fe5daa, 32'hc44e17e2, 32'hc3082de7},
  {32'hc4c8e016, 32'h42824f96, 32'hc394d425},
  {32'h450067c4, 32'h400eb978, 32'hc304b1f9},
  {32'hc293ade0, 32'h430c0a40, 32'h43076d72},
  {32'h447e66f0, 32'hc3197021, 32'h42ecef73},
  {32'hc45c025c, 32'hc2a9fb28, 32'hc2f2538e},
  {32'h449a67a8, 32'h42ce9ebc, 32'h43807a23},
  {32'hc4c9fd7c, 32'h4229cf69, 32'h42082ebc},
  {32'h44dba566, 32'h41b2c263, 32'hc36a278f},
  {32'hc4db0ca5, 32'h43ecb9d0, 32'hc27d794a},
  {32'h4504c170, 32'hc3150479, 32'hc3882b62},
  {32'hc3a58f40, 32'h43e9b486, 32'hc2f7c68d},
  {32'h44a0cbc3, 32'h43a7da1b, 32'hc29ee545},
  {32'hc30f12d6, 32'h42df2575, 32'hc3f5723f},
  {32'h447405fc, 32'h3fbd0660, 32'h4408f5d8},
  {32'hc3792848, 32'h43f36ad2, 32'h40f9129d},
  {32'h4433e76e, 32'h4272624b, 32'hc29a61fc},
  {32'hc1d94a50, 32'hc30dea5e, 32'hc3645c95},
  {32'h44ea74e9, 32'h42be2ba1, 32'hc350f072},
  {32'hc4c1bc51, 32'h43938a6d, 32'h428790c6},
  {32'h4515598a, 32'hc178e0ec, 32'h438a375f},
  {32'hc4da8a82, 32'h43ae0c52, 32'h408b20e7},
  {32'h44ab23f2, 32'hc25427c8, 32'h42942100},
  {32'hc44c99b4, 32'hc3d362fb, 32'h43015d70},
  {32'h43ea8140, 32'h4306a828, 32'hc306db55},
  {32'hc5023e30, 32'hc2ca5756, 32'hc3a8f96a},
  {32'h43f7c90c, 32'h431b96eb, 32'h426e8166},
  {32'hc346cd1c, 32'h43be2433, 32'hc2c61d3b},
  {32'h419bafc0, 32'hc151a3df, 32'h42fefa59},
  {32'hc39d8f38, 32'h442b991c, 32'h434416dd},
  {32'h4468a250, 32'hc32b2ec0, 32'h4328ec06},
  {32'hc4b865d8, 32'hc29b13e8, 32'hc35fbb88},
  {32'h44efc6c8, 32'h42c1116f, 32'hc32514e0},
  {32'hc4d774ab, 32'hc2eaff75, 32'h43a2dad5},
  {32'h450edc33, 32'h4221bce8, 32'h4367e840},
  {32'hc48f3ce4, 32'hc383e29d, 32'hc342e0dc},
  {32'h434d53fd, 32'h4434c877, 32'h441b45c8},
  {32'hc5153eed, 32'hc305844a, 32'h4387ba5d},
  {32'h45043d6c, 32'hc1a95593, 32'hc3a26318},
  {32'hc49e161f, 32'hc1497928, 32'h43b38382},
  {32'h44ecda41, 32'h436e3714, 32'h43c566e7},
  {32'hc47660ac, 32'hc3a9974e, 32'hc300cf09},
  {32'h44319ca1, 32'hc2806728, 32'h43a0f968},
  {32'hc38ce806, 32'h42dc0331, 32'h42789df9},
  {32'h450e9d54, 32'hc181e5ed, 32'hc3a730f6},
  {32'hc4d3215a, 32'hc32efab1, 32'h430f6025},
  {32'h44d3056a, 32'hc30ce8f0, 32'h430890bf},
  {32'hc17db54c, 32'h43d07216, 32'hc3a4e38c},
  {32'h4408c137, 32'hc2c9d8b7, 32'hc3153985},
  {32'hc2df374e, 32'h43b36570, 32'h42ac58eb},
  {32'h44468130, 32'hc30c8cf6, 32'hc2f2bab8},
  {32'hc342835a, 32'h43bdf25f, 32'hc3717201},
  {32'h44c8f5d6, 32'h4398ea31, 32'h430daed8},
  {32'hc4420d49, 32'hc39b8258, 32'h41f91c62},
  {32'h44e897c7, 32'h4218a3e6, 32'h43ab0581},
  {32'hc50aeea4, 32'h429b2299, 32'hc2888aa6},
  {32'h4415f4ec, 32'hc2f70cd7, 32'h43591904},
  {32'hc4ac915f, 32'h43847ac1, 32'h41c63293},
  {32'h43a7c5d9, 32'h4319e81c, 32'hc2373dcb},
  {32'hc37e1390, 32'hc3ca32fb, 32'h4359d650},
  {32'h44ec9634, 32'h430f268b, 32'hc27fadca},
  {32'h42ca47e0, 32'h42cb918b, 32'h43a21840},
  {32'h44f589b4, 32'h4383b31c, 32'h43f5e7f8},
  {32'hc3b0ff36, 32'h43463785, 32'h4381b507},
  {32'h44ba550a, 32'hc23c1cc6, 32'h430aa6a7},
  {32'hc4a335e9, 32'h43a34de2, 32'hc1690241},
  {32'h44d85d06, 32'hc2a5b203, 32'h43d9eff2},
  {32'hc491dd10, 32'h43314053, 32'hc3677f38},
  {32'h445eff18, 32'hc2675d0e, 32'h4109b184},
  {32'hc31c40d8, 32'hc14350b7, 32'h4280a6df},
  {32'h430f86d8, 32'h42613ab3, 32'h43fdc1fb},
  {32'hc4a446e6, 32'h431ea20a, 32'hc290ad55},
  {32'h444bbde2, 32'h441d6610, 32'hc2da17c3},
  {32'hc4869c73, 32'hc0aeef93, 32'hc340c2b2},
  {32'h4450cea0, 32'hc296e094, 32'h42e60162},
  {32'hc38318f2, 32'hc2ad557c, 32'h42831380},
  {32'h44a5c474, 32'h42c62f4a, 32'h4091a7bd},
  {32'hc4f2be09, 32'hc38bc041, 32'h4315acda},
  {32'hc3c79084, 32'hc33aac96, 32'hc3987e12},
  {32'h44e21e92, 32'hc1326dc4, 32'h4327e2ca},
  {32'hc489b123, 32'h43040dd6, 32'hc2d54174},
  {32'h44ee9c5c, 32'h4309ed9c, 32'h42fc28f4},
  {32'hc5042318, 32'hbfc5391e, 32'hc1da88a8},
  {32'h44fc025b, 32'hc29e5593, 32'hc24b5291},
  {32'hc43087e9, 32'hc1bdd6f1, 32'hc34eb2e5},
  {32'h446b145e, 32'h4341ce69, 32'hc3ab20ad},
  {32'hc4966562, 32'hc23cfee4, 32'hc31a8fa8},
  {32'h45065f0c, 32'hc32b783e, 32'h434cfdf2},
  {32'hc4f10e68, 32'hc323f7dc, 32'hc01d0023},
  {32'h450bca69, 32'hc3b149d0, 32'h43de59f0},
  {32'hc4849242, 32'hc390514a, 32'hc3041694},
  {32'h43393a0c, 32'h4303679d, 32'hc34b9d3f},
  {32'hc49e6f9e, 32'h43233de6, 32'h430262ae},
  {32'h43eb2812, 32'h41587b62, 32'hc4139eff},
  {32'hc30d8d20, 32'hc26dbb66, 32'h42c33456},
  {32'h45218582, 32'hc3a5843a, 32'h4383f9b2},
  {32'hc4250bb0, 32'h42215c39, 32'hc1949cf6},
  {32'h440856f0, 32'hc3207616, 32'hc33f5b59},
  {32'hc4389c9d, 32'h4396ee09, 32'hc33c9ea7},
  {32'h446e7912, 32'h42c7c8ae, 32'h42909a18},
  {32'hc4eaae67, 32'hc41a1d59, 32'h41f0ff67},
  {32'hc2d46cf0, 32'h4321ea8b, 32'h4390d707},
  {32'hc3cca83c, 32'hc37c8e66, 32'hc1eeed34},
  {32'h44cd1d51, 32'hc2c16785, 32'h41a11cb8},
  {32'hc4bda167, 32'h4313a141, 32'h42ecc312},
  {32'h44ea2cda, 32'hc345ed7c, 32'hc224c591},
  {32'hc3f90bb8, 32'h433d5dd3, 32'hc3c0670c},
  {32'hc4ae3d5f, 32'h42f34df0, 32'h438cff0f},
  {32'h441fad44, 32'hc332282f, 32'hc267ed63},
  {32'hc1dde1e0, 32'h419b04c6, 32'h420bca5e},
  {32'h44ed6c58, 32'hc31083f9, 32'hc3038dda},
  {32'hc49ad77d, 32'hc338d6de, 32'hc370a7d5},
  {32'h43fe9fb8, 32'hc243b7e5, 32'h42c19f24},
  {32'hc4ab2522, 32'h41df439a, 32'hc31ebb57},
  {32'h4308472e, 32'h42ad59d2, 32'h42df006c},
  {32'hc4c819a6, 32'h42111fd2, 32'hc312ce1b},
  {32'h44154b32, 32'h4324c46e, 32'hc1350cf1},
  {32'hc4f83035, 32'h4369abeb, 32'hc32bf861},
  {32'h44ae495b, 32'hc32a37c6, 32'hc3ac8cce},
  {32'hc405b390, 32'h435c769b, 32'hc12b6792},
  {32'h45101fb0, 32'h43a8e3c3, 32'hc380667a},
  {32'h420c4405, 32'hc2b4922b, 32'h42fefc5b},
  {32'h443272a8, 32'h42f9bc53, 32'h439fd590},
  {32'hc50db12e, 32'hc278c8f8, 32'h42187c2c},
  {32'h45089a3c, 32'h4367cbac, 32'h43742e67},
  {32'hc3149d60, 32'h426d387a, 32'h42abe524},
  {32'hc2addf14, 32'hc36bf891, 32'hc27d7f89},
  {32'hc5096cbc, 32'h42b98ba1, 32'hc3a8f31c},
  {32'h4354a3f8, 32'h42c73bd0, 32'h440d072c},
  {32'hc51584bf, 32'h430e0127, 32'h4309a544},
  {32'h43eb1429, 32'h42a218a8, 32'h436e87f0},
  {32'hc4e9cfe0, 32'h4325d980, 32'hc2841c8f},
  {32'h44ab526c, 32'hc3309bd1, 32'hc3a65f27},
  {32'hc4469eba, 32'h437869d1, 32'h42b33318},
  {32'h43317d30, 32'h4088dc50, 32'h43ce9859},
  {32'hc4868f67, 32'hc3b7e87d, 32'h42a9fa9a},
  {32'h44d085c7, 32'hc1756b86, 32'hc39f76a2},
  {32'hc3a1ac88, 32'hc290b194, 32'h43021d21},
  {32'h44f257dc, 32'h42dd9140, 32'h439973e5},
  {32'hc50278d8, 32'hc4102bb6, 32'hc3415826},
  {32'h43c6a71a, 32'h4337f5fe, 32'h41e3df07},
  {32'hc45ef853, 32'h43a05183, 32'h42ff88fd},
  {32'h44d63730, 32'h43dfa7d6, 32'hc30cc088},
  {32'hc2480780, 32'hc15391a6, 32'h42496d78},
  {32'h4410e99d, 32'hc2f0c763, 32'hc33438af},
  {32'hc3f35093, 32'h43b1121d, 32'hc395fc71},
  {32'h42463060, 32'hc2ebcadd, 32'hc239ca6d},
  {32'hc453fa0b, 32'h4311f8fe, 32'h43456473},
  {32'h44e6ec37, 32'hc3653064, 32'hc3a6f002},
  {32'h43834460, 32'h440cf2e1, 32'hc2f37ba3},
  {32'h43b40774, 32'h43ada588, 32'hc2d8f608},
  {32'hc4e2c675, 32'hc3067355, 32'h43572668},
  {32'h44b3d160, 32'h42bf8bfa, 32'h4206a854},
  {32'hc42cbbdc, 32'h43159b55, 32'hc249e0a7},
  {32'h45116884, 32'hc3b483fd, 32'h4314907a},
  {32'hc50e6760, 32'hc345dc30, 32'hc34a58fe},
  {32'h4523d9b6, 32'hc333f93e, 32'h43bf83f7},
  {32'hc4917ad4, 32'h420f0c40, 32'hc34fe12a},
  {32'hc4f1f51a, 32'hc3132fd7, 32'h42b1a318},
  {32'h44cf6ee0, 32'h42937a30, 32'h4362ac51},
  {32'hc4883945, 32'hc18eba60, 32'h43181a4b},
  {32'h431f4a1c, 32'h42efb37e, 32'hc30290b0},
  {32'hc28e2cf0, 32'h42c2e6f5, 32'h42fdb346},
  {32'h44901696, 32'hc2e53198, 32'h433aff2a},
  {32'hc52704e1, 32'h437a7047, 32'h423bc094},
  {32'h44b665a4, 32'hc331363d, 32'h42caad2e},
  {32'hc423a8de, 32'h4212bcf8, 32'h4308c85d},
  {32'h44c50334, 32'hc20c3d16, 32'hc3a8d127},
  {32'hc430db72, 32'hbf6d1ff0, 32'h43b373f8},
  {32'h43e417c5, 32'h434f941b, 32'h431750a0},
  {32'hc4d2c1c2, 32'hc336ea81, 32'hc33e7610},
  {32'h42ead830, 32'h42cfcb82, 32'hc36a0d49},
  {32'hc3be876e, 32'hc270d9d3, 32'h43c6097e},
  {32'h447ab052, 32'h429819f9, 32'hc34b8f48},
  {32'h4285ebcc, 32'hc3930fc6, 32'hc31b4e87},
  {32'h440687d6, 32'h43c9282f, 32'hc3cd7810},
  {32'hc3a008a8, 32'hc129c71a, 32'h42ff92bd},
  {32'h44da5f42, 32'h4379e403, 32'hc3af1245},
  {32'hc3c65360, 32'h43b6803a, 32'h4368e197},
  {32'h441fa3fc, 32'h437e69a1, 32'hc18293d2},
  {32'hc4478b8e, 32'h441a6c25, 32'h4374b8ed},
  {32'h448dec3c, 32'h422f57d0, 32'hc0dae077},
  {32'hc4a5ac14, 32'h4122863d, 32'hc2a33600},
  {32'h448d084e, 32'hc39f0c54, 32'hc16fdf30},
  {32'hc2bc6ff4, 32'hc2143f3a, 32'hc32416e6},
  {32'h44dfada3, 32'h4316dcf2, 32'hc3a0c1be},
  {32'hc464b314, 32'h43685ff1, 32'h430ab380},
  {32'h443a0162, 32'h40f0f25a, 32'hc3c5573b},
  {32'hc504ff06, 32'h435c541d, 32'hc15bf6e9},
  {32'h4415ae19, 32'hc2f13614, 32'h42dc820b},
  {32'hc1f47080, 32'h43a63fc1, 32'h4325f2e9},
  {32'h42ae6440, 32'hc2798490, 32'h4308a190},
  {32'hc4954e08, 32'hc1f6cb20, 32'h43b34a99},
  {32'h43d1e530, 32'hc2eba408, 32'h42ac3b3b},
  {32'hc4c23cad, 32'h435f67f9, 32'h430e9012},
  {32'h43cade96, 32'hc2c8e360, 32'hc2931051},
  {32'hc4f482a5, 32'h4326f251, 32'h432238c4},
  {32'h44b39d84, 32'hc37ce5b2, 32'hc3aed37a},
  {32'hc5025ae2, 32'h434c48b8, 32'h42c7d493},
  {32'h44211703, 32'hc23fd0c7, 32'hc30b1607},
  {32'hc4db5736, 32'hc297b112, 32'h4423ef97},
  {32'h44e2ad35, 32'h426c6e0c, 32'h432ae3f0},
  {32'hc32398b3, 32'h426bc646, 32'hc12cecea},
  {32'h43b46ada, 32'hc40e3cf6, 32'h4338f0e7},
  {32'hc4d449a8, 32'h4306c2c8, 32'h4337b580},
  {32'h44c39b80, 32'h439d45c3, 32'hc4127f5b},
  {32'h4328916e, 32'hc36d95bc, 32'h434bcfce},
  {32'hc36efd50, 32'h4312975d, 32'h4397bf13},
  {32'hc502bf59, 32'h4297c1bb, 32'h433e3aef},
  {32'h43d16750, 32'h41a16090, 32'hc33f0d34},
  {32'hc35a5bc4, 32'h42f993e0, 32'h4306a86b},
  {32'h4500147f, 32'h40f920f4, 32'hc35c6e48},
  {32'hc503aed7, 32'hc355d7c3, 32'hc17c1a8e},
  {32'h446a8b1b, 32'h4383660d, 32'h4095bdbf},
  {32'hc4cd6d69, 32'hc36a659d, 32'h438fdfbf},
  {32'h4488ac15, 32'hc3783b1c, 32'hc243f0fb},
  {32'hc4e0dc6d, 32'hc318306f, 32'h43288563},
  {32'h44846f1a, 32'hc38b109c, 32'hc1e05f79},
  {32'hc507d4a8, 32'h42916bae, 32'h443fb32b},
  {32'h449a1048, 32'hc3299965, 32'h438ea69e},
  {32'hc51e8b07, 32'h43413ac7, 32'hc211d7d6},
  {32'h44ece354, 32'h4302ebb0, 32'hc30c56ac},
  {32'hc4b8ea52, 32'h42b6dda5, 32'h43a653eb},
  {32'h443ee904, 32'h436c72db, 32'hc1e62e87},
  {32'hc424363e, 32'hc3b78c19, 32'h4388fe6e},
  {32'h43976e97, 32'hc2ffaf65, 32'h439754e7},
  {32'hc2a9302c, 32'h4343520d, 32'hc33f19dd},
  {32'h44bea35a, 32'h43b11444, 32'h43ce1e70},
  {32'hc48b2719, 32'hc34d0d43, 32'h42c268a2},
  {32'h449e9828, 32'hc212b4bf, 32'h43a57092},
  {32'hc40725c6, 32'hc22c1ce5, 32'h436027bb},
  {32'h4503f53b, 32'h43ada5e3, 32'h4423d599},
  {32'hc4433394, 32'h42895ea2, 32'hc272f1b0},
  {32'h44b3ac6d, 32'hc3d68415, 32'h40aea248},
  {32'hc4c92d28, 32'h431751d5, 32'hc2f180c5},
  {32'h4501bca3, 32'hc239d83f, 32'hc2f8786e},
  {32'hc5182fd2, 32'hc112e73e, 32'h42e1098e},
  {32'h447a9526, 32'h42840a46, 32'hc36464f7},
  {32'h42a24f40, 32'h436b2d2e, 32'hc31ba4d0},
  {32'h44106dc8, 32'h435e1145, 32'h428a023e},
  {32'hc5139d47, 32'hc1dccf13, 32'h404eaee2},
  {32'h44c7d796, 32'h435ae4ea, 32'h437246ed},
  {32'hc5060211, 32'hc31f2758, 32'h43c07e9f},
  {32'h42dd1750, 32'h439ce066, 32'h4345d289},
  {32'hc41f7efa, 32'hc3828730, 32'h433995fd},
  {32'h4496ad0c, 32'hc3426b8c, 32'h42cfb2e4},
  {32'hc4fedc5b, 32'h42da0349, 32'hc1d07227},
  {32'h44b5979c, 32'hc39e9ab8, 32'hc397dbe6},
  {32'hc401f37a, 32'h3fd111cd, 32'hc353998c},
  {32'h44ebd4c9, 32'hc39f4e6e, 32'hc32bd5bc},
  {32'hc4ac0b92, 32'hc2781290, 32'hc322d94c},
  {32'h44f9edad, 32'h41e20c2c, 32'h43acd870},
  {32'hc4da96a6, 32'hc31296eb, 32'hc3a9d863},
  {32'h44c2beef, 32'hc380b5c9, 32'hc25f527b},
  {32'hc4da328a, 32'h42133c5a, 32'hc3ae548e},
  {32'h442b6ec4, 32'h4253ada8, 32'h4332eb29},
  {32'hc46157a1, 32'h431f8394, 32'h42bee425},
  {32'h4402125c, 32'hc2ddd178, 32'hc327d6a1},
  {32'hc49a79aa, 32'hc225430a, 32'hc2203bda},
  {32'h450387d0, 32'hc250c747, 32'h40c4ff4f},
  {32'hc4dfe30a, 32'hc300299b, 32'h42b30047},
  {32'h4502a704, 32'h43162b56, 32'h4366b798},
  {32'hc46968d4, 32'h4403d8dc, 32'hc3833dc9},
  {32'h4394bb64, 32'hc2a15106, 32'hbf9c1f99},
  {32'hc3d8e268, 32'hc381dcfa, 32'h4402cdd5},
  {32'h44e9db79, 32'h4364b4e1, 32'hc28cec24},
  {32'hc4610308, 32'h4393639f, 32'h430c6b1e},
  {32'h448bf1d0, 32'hc38db4f2, 32'h43b2625e},
  {32'hc47af544, 32'hc2f2c578, 32'h435995b3},
  {32'h44820c9a, 32'h430ebda3, 32'h42200341},
  {32'hc4940960, 32'h438ae60d, 32'h430752d0},
  {32'h43667ce2, 32'hc3f86a3b, 32'h3fd2b3b2},
  {32'hc5078de2, 32'h43862a27, 32'hc20a4072},
  {32'h44a80631, 32'h4310d21a, 32'hc216b277},
  {32'hc50065ae, 32'hc30ccd0c, 32'hc3b1c4d2},
  {32'h44829488, 32'h42b15acb, 32'h434383f0},
  {32'hc507dbc6, 32'hc3ec68e1, 32'h438d14cc},
  {32'h45054660, 32'h41670284, 32'h42a17305},
  {32'hc32486c3, 32'h43cc37f4, 32'hc22fa161},
  {32'h45038d8a, 32'h422bb1e0, 32'hc3af8433},
  {32'hc487e9a2, 32'hc28f59f7, 32'h439b27d6},
  {32'h44cc964e, 32'h427b0dd5, 32'hc2af28f6},
  {32'hc45ea50a, 32'hc3810f76, 32'h437b34a6},
  {32'h450c5fb9, 32'hc37c9ed5, 32'hc171ac62},
  {32'hc42d3f04, 32'h437aef82, 32'hc3a71c1c},
  {32'h448ac908, 32'h43629bcb, 32'h437e10bb},
  {32'hc485c67c, 32'h42c1c0e0, 32'h42aa2ec2},
  {32'h44ab8ac8, 32'hc36aa4ed, 32'hc44318ae},
  {32'hc42ef9c8, 32'h429d7c5c, 32'hc1ae0265},
  {32'h4500dfca, 32'hc36a6533, 32'h43ad94e8},
  {32'hc4f3df4d, 32'h433e97b9, 32'hc2c882ba},
  {32'h43d24560, 32'hc38c86ed, 32'hc25d81d7},
  {32'hc4c351d8, 32'h434e3659, 32'hc2acd4a7},
  {32'h43b88644, 32'h432ff63d, 32'h43489dd6},
  {32'hc43d0e9b, 32'h42df8345, 32'h42a90482},
  {32'h449badce, 32'hc368a53d, 32'h4318092a},
  {32'hc47d374b, 32'hc389635f, 32'h43d8239b},
  {32'h414d0b40, 32'h434e7c65, 32'hc2ce7c75},
  {32'hc488d058, 32'h43efce39, 32'h42d141b4},
  {32'h44a7455b, 32'hc41cec29, 32'hbf1a1be0},
  {32'hc5148903, 32'hc3aeb80a, 32'h416fd152},
  {32'h44bca816, 32'h439b0d38, 32'hc368e124},
  {32'hc4ca6582, 32'h43799c4a, 32'h43497af9},
  {32'h43c4fee0, 32'hc33e14de, 32'hc40ad023},
  {32'hc50017f5, 32'hc3aa7f55, 32'h422b58df},
  {32'h44899df4, 32'hc1a8137c, 32'h428d9248},
  {32'hc48b9987, 32'hc38fb125, 32'hbf2f8166},
  {32'h447aedf9, 32'h4362279c, 32'hc38101c9},
  {32'hc4218965, 32'hc209af3b, 32'hbf9a2c10},
  {32'h443f8331, 32'hc400180d, 32'h42331850},
  {32'hc4c08e76, 32'hc2942ed2, 32'h415210a2},
  {32'h44d2b7ca, 32'hc3ba335b, 32'h4363eca8},
  {32'hc427d3ff, 32'hc2f80113, 32'h42c8c08c},
  {32'h444f26d3, 32'h43a1120c, 32'h43789723},
  {32'hc504e507, 32'hc3c0007c, 32'hc321a3c7},
  {32'h431253ee, 32'hc3abac8c, 32'hc2a56bfa},
  {32'hc4f04779, 32'hc2f7855b, 32'hc3e7d09d},
  {32'h44411e0a, 32'hc2c969cd, 32'hc1df2f47},
  {32'hc4f0e3c9, 32'hc12234dc, 32'h4319740e},
  {32'h44b85530, 32'hc37ac98f, 32'hc3810504},
  {32'hc4f91c88, 32'h43f3e500, 32'h43aed857},
  {32'h45173745, 32'hc39e7fed, 32'h4312fa7c},
  {32'hc440dd9c, 32'h43bf8cfa, 32'h42a413a0},
  {32'h4491c884, 32'hc2c9533e, 32'h41c6d5ac},
  {32'h4353375b, 32'h43d41593, 32'hc341012f},
  {32'h442b6814, 32'hc36f49a2, 32'h43360b6c},
  {32'hc49ce142, 32'h431e1a4d, 32'hc3722677},
  {32'h4509f1bc, 32'h43ca3e13, 32'h43a8ed73},
  {32'hc50af7e8, 32'hc3268ad5, 32'h43718dd0},
  {32'h43cb4322, 32'hc2d7805b, 32'hc2949d7c},
  {32'hc50f8397, 32'h42f67c40, 32'h42f80eb2},
  {32'h448abe4a, 32'hc187943a, 32'h4072cf2a},
  {32'hc5020e8a, 32'h431623ac, 32'hc19c6e2c},
  {32'h44fe5f32, 32'h43b60adb, 32'h42aa7393},
  {32'hc5072e48, 32'hc3ba3ef7, 32'hc3a7eb80},
  {32'h447669ae, 32'hc35fd85d, 32'hc14f0521},
  {32'hc4ba4b1e, 32'hc21a4079, 32'h42fa8e2d},
  {32'h4489ab4d, 32'hc20fc792, 32'h4361b024},
  {32'hc5120eb6, 32'h44237825, 32'hc335329e},
  {32'h43b3831a, 32'h43167421, 32'h43ac0c21},
  {32'hc438ca5c, 32'hc4089c85, 32'h42801dcc},
  {32'h451584f6, 32'h4377ca8e, 32'h432f5c43},
  {32'hc4380010, 32'hc0221dc7, 32'h42f8cb4a},
  {32'h43609be4, 32'hc328e325, 32'h43aac3f5},
  {32'hc51e7737, 32'hc369445d, 32'h4329eb53},
  {32'h449f166e, 32'h439c7f59, 32'h42b79947},
  {32'hc516e4c8, 32'h41e80c08, 32'hc2b1b07a},
  {32'h44e8fa7a, 32'h42185664, 32'hc31c3e9a},
  {32'hc2600c80, 32'hc35d8975, 32'hc3406ba8},
  {32'h448900e2, 32'h43b2a3e6, 32'hc3ab2835},
  {32'hc411922c, 32'h43102260, 32'h432eca24},
  {32'h41ff9a10, 32'hc3bd637f, 32'h435ed6c6},
  {32'hc395d4c4, 32'h43de70aa, 32'hc31d6ccf},
  {32'h44c4041f, 32'h44034c07, 32'h43a649d0},
  {32'hc52303f8, 32'h43157c5e, 32'hc38a8c9b},
  {32'h43ac60ce, 32'hc34181e7, 32'hc283e79f},
  {32'h42a0140d, 32'hc3a5f8d8, 32'hc39673eb},
  {32'h444a8a4a, 32'h43a122f7, 32'h43a9c5ba},
  {32'hc4f1a366, 32'h432f34cf, 32'hc3438f48},
  {32'h443d3170, 32'h4321c9a9, 32'hc329b1bd},
  {32'hc34442e0, 32'h429abe78, 32'hc340d1cb},
  {32'h448d87dc, 32'hc3b66e2d, 32'h439404eb},
  {32'hc4a50239, 32'h42979f7c, 32'h4088e888},
  {32'h44210120, 32'hc364c51f, 32'hc28258ec},
  {32'hc1dbc800, 32'hc376ff53, 32'h43532a40},
  {32'h43bc5a92, 32'h44167c70, 32'hc1db259f},
  {32'hc4edde19, 32'hc103d872, 32'hc31911fd},
  {32'h4332c158, 32'hc31e00ae, 32'h4368fe9e},
  {32'hc3e31f22, 32'hc2028b5a, 32'hc30d5497},
  {32'h44dfad87, 32'hc25b5c44, 32'h42f41e00},
  {32'hc4ff7850, 32'hc373f22b, 32'h424452bc},
  {32'h45050fde, 32'h431dfba0, 32'hc341fe4a},
  {32'hc50d69fd, 32'hc3816deb, 32'h430a794d},
  {32'h44d9bf6c, 32'hc3452da3, 32'h43f707e8},
  {32'hc3cdbd94, 32'h4351c7bc, 32'h426943d0},
  {32'h44d8f2b0, 32'hc351dcc0, 32'h43dc9550},
  {32'hc49ac8ab, 32'h4321f1d7, 32'hc272beba},
  {32'h44be13b3, 32'hc32aac7c, 32'hc30c8b8e},
  {32'hc4f5faaf, 32'h4361d7c6, 32'hc28f1033},
  {32'h431f76d4, 32'hc3f07a14, 32'hc32bac44},
  {32'hc3ed120a, 32'hc35ab9c2, 32'h42340869},
  {32'h44ac2f51, 32'hc3e421c6, 32'h42d8a8be},
  {32'hc495abd9, 32'h4339f80c, 32'hc3b1c657},
  {32'h4490e374, 32'hc395d908, 32'h42a5118f},
  {32'hc405e540, 32'hc2a6988f, 32'h43c0c804},
  {32'h440c21f2, 32'h42b6082c, 32'hc2c35176},
  {32'hc46aa5ea, 32'h42bdaf15, 32'hc28f0bc8},
  {32'hc4a5ff1f, 32'hc33a9636, 32'hc2e106ba},
  {32'h444e0303, 32'h43ce202d, 32'h43b3505c},
  {32'hc19bd77c, 32'h440abb44, 32'hc31e419d},
  {32'h443e0238, 32'h41afa062, 32'hc3718f6b},
  {32'hc3cee72c, 32'hc29f00b9, 32'hc3ccebf4},
  {32'h442c1bbc, 32'h4379e869, 32'h4296d0e5},
  {32'hc4c0a6c5, 32'h43d82826, 32'hc31a4a23},
  {32'h444816f2, 32'h429ea3ce, 32'h40aab7ac},
  {32'hc4efcdfd, 32'hc30fcb54, 32'hc3853448},
  {32'h4475e994, 32'hc3b9eac6, 32'hc38509d7},
  {32'hc4464f84, 32'h42f2ea57, 32'hc358a5cf},
  {32'h448c92c4, 32'h433d5f06, 32'h431efc36},
  {32'hc4994c7b, 32'hc36cbbfe, 32'hc3b440dd},
  {32'h44aa863a, 32'hc3319acc, 32'hc3e81609},
  {32'hc4d482da, 32'hc2446adb, 32'hc1c19ad0},
  {32'h44661f1e, 32'h42451dee, 32'h427b6dd8},
  {32'hc3222ab8, 32'hc2a35158, 32'hc3864fd2},
  {32'h450faa09, 32'h4227d3a1, 32'hc302139a},
  {32'hc3ed6227, 32'hc39c2e6b, 32'h43ce5ebd},
  {32'h450e1d10, 32'hc3a96ab7, 32'h42f93775},
  {32'hc4530570, 32'h438b7b5c, 32'hc4236e83},
  {32'hc4d192c3, 32'hbfaa1b01, 32'hc303abea},
  {32'h44650a33, 32'h435c53c0, 32'hc3926654},
  {32'hc47f4d85, 32'hc1c156a6, 32'h42dbfc0a},
  {32'h4389f010, 32'hc2636a83, 32'h438ec546},
  {32'h42efbea8, 32'h43752b65, 32'h437b1d4f},
  {32'h44a70bca, 32'h44266ed0, 32'h43baec4e},
  {32'hc4f787ea, 32'h433c1a8d, 32'h43bdaca0},
  {32'h40456e80, 32'h4343b4ec, 32'hc4150682},
  {32'hc452a6fa, 32'h430e0acb, 32'h433178ec},
  {32'h4470f734, 32'hc1895035, 32'h4053bc44},
  {32'hc512a869, 32'hc334a43c, 32'hc3cff219},
  {32'h450862c4, 32'hc33fe6ea, 32'hc2b84674},
  {32'hc4e774c7, 32'hc340ecb1, 32'hc343773f},
  {32'h43813483, 32'hc2acbb56, 32'h43892794},
  {32'hc4fd2260, 32'hc350c739, 32'hc3524764},
  {32'h444f9a18, 32'hc380d2d4, 32'h43389d34},
  {32'hc3fb1a0b, 32'h4064bcc4, 32'hc30f2c16},
  {32'h44db746e, 32'hc3f1019d, 32'hc3cb2438},
  {32'hc514391c, 32'h434c5c04, 32'hc323831b},
  {32'hc3cee114, 32'h42c2100b, 32'h426d2917},
  {32'hc3cba458, 32'h43bfd8a9, 32'h4200d8ec},
  {32'h4477c4c5, 32'hc2acae57, 32'h41714ed5},
  {32'hc4b507a7, 32'h41f14b2e, 32'hc2f2acc2},
  {32'h44f58a10, 32'h439ecbc7, 32'h43a573ea},
  {32'hc4f7eb58, 32'hc3eac329, 32'h4352ebc8},
  {32'h45044eb3, 32'h4372b92d, 32'h43057f9a},
  {32'hc48eceb0, 32'h42f28f86, 32'hc3587b1d},
  {32'h44a30e12, 32'hc1901b35, 32'hc3c3f78f},
  {32'hc437d33e, 32'h436d7b07, 32'h42c80cce},
  {32'h44254234, 32'hc2c2b504, 32'hc30dc048},
  {32'hc4e398c2, 32'hc3c255ad, 32'hc2a20816},
  {32'h4524921e, 32'hc38ed64f, 32'hc2c2c03b},
  {32'hc4c1dca1, 32'hc26eab0e, 32'hc296056f},
  {32'h4452acb6, 32'hc23f5fb8, 32'h42039a10},
  {32'hc456ffa6, 32'h431c0842, 32'hc3111bcf},
  {32'h44be6fac, 32'hc24efb4e, 32'h435e9e52},
  {32'hc40ac6de, 32'hc36cf7d9, 32'h43c1e739},
  {32'h432b2230, 32'hc3c266c1, 32'hc2635fb7},
  {32'hc447b19b, 32'h436d81c1, 32'hc2563618},
  {32'h44146404, 32'hc2edd6d2, 32'hc2997d8b},
  {32'hc3fea8dc, 32'hc39131ca, 32'h42041145},
  {32'h4526db4e, 32'h4326a813, 32'hc27cb6e0},
  {32'hc393ca5a, 32'h43432056, 32'hc2a4d312},
  {32'h44eaef03, 32'hc3282090, 32'hc38e4dbd},
  {32'hc419b848, 32'hc3af2ad1, 32'h42e28781},
  {32'h43f212bd, 32'h41b72db3, 32'hc38606b8},
  {32'hc476b411, 32'hc3046042, 32'hc3595f9a},
  {32'h44a8a356, 32'h430d6663, 32'hc38db0e6},
  {32'hc46cbe5e, 32'h437924e2, 32'hc24e7f67},
  {32'h451ac405, 32'h42f677ae, 32'h42730e48},
  {32'hc2742a80, 32'hc2ba6256, 32'h43ef5c72},
  {32'h44bb9854, 32'hc3decdc8, 32'hc310c742},
  {32'hc5099586, 32'h42e246e4, 32'hc36a18a8},
  {32'h450c72c7, 32'hc2300ca3, 32'h42ed8257},
  {32'hc43bb958, 32'h427bef34, 32'h432b300a},
  {32'h42219680, 32'h3e2d73c0, 32'hc289e064},
  {32'hc4fdd49f, 32'hc309ebb4, 32'hc371ba1c},
  {32'h443ddadc, 32'h429de66a, 32'h43f3ea1d},
  {32'hc48fc768, 32'h40dca48c, 32'hc3b63850},
  {32'h4420af00, 32'h41a28162, 32'h42c39131},
  {32'h4273d960, 32'h43e7647a, 32'hc3665ef4},
  {32'h44723b30, 32'h438227e4, 32'hc2f0ca84},
  {32'hc3ba6b2a, 32'h439941ff, 32'h4359e21b},
  {32'h44cede0e, 32'h438e52a0, 32'hc3964f8e},
  {32'hc5190d45, 32'h42d9a0e2, 32'h43125f97},
  {32'h450bc06e, 32'h4308dcf0, 32'hc3b3afa8},
  {32'hc4e96b94, 32'h434c53e5, 32'hc3a27a0e},
  {32'h438d8157, 32'h4309689b, 32'hc31d7d57},
  {32'hc4ebb407, 32'h42c62c27, 32'h4244ba8a},
  {32'h4505a541, 32'hc2d8ddc4, 32'h4300df8c},
  {32'hc49d5414, 32'hc31045e1, 32'h433c88be},
  {32'h44556168, 32'h4220a41d, 32'h42a91670},
  {32'hc48a7e8a, 32'h43bd20ab, 32'h40f4a114},
  {32'h43542058, 32'hc3a4e21f, 32'hc36d8405},
  {32'hc4098dde, 32'h43c8ce20, 32'h433e4bcf},
  {32'h4460e716, 32'hc219c3ba, 32'h40d30251},
  {32'hc44f37c4, 32'h431e689d, 32'h43152ce8},
  {32'h444e72ad, 32'h418969e8, 32'h4154cf6e},
  {32'hc49f9343, 32'hc221b87a, 32'h42d988d6},
  {32'h441804f8, 32'hc30e50ee, 32'hc31cbfe5},
  {32'hc4df392d, 32'hc28a5b1e, 32'hc2060057},
  {32'h4423a286, 32'hc38fbae9, 32'hc39f6726},
  {32'hc41be53c, 32'hc310470e, 32'h441c2df5},
  {32'hc3241650, 32'hc14b13bb, 32'h41aeca61},
  {32'h43aea59c, 32'hc2a07f7e, 32'h430b7a9e},
  {32'h448e7517, 32'hc352e60e, 32'hc4049277},
  {32'hc4fd5a68, 32'hc43c4689, 32'h42e515b9},
  {32'h43d2d6a6, 32'h42ef038b, 32'hc307bff6},
  {32'hc3d3afac, 32'hc3a310d6, 32'h438113a8},
  {32'h445b14ec, 32'h43a9f978, 32'h435fa992},
  {32'hc502cdd2, 32'hc177e198, 32'h434d979d},
  {32'h44f9160d, 32'h42973042, 32'hc1842126},
  {32'hc4df4f6d, 32'h420b0f21, 32'h43d13951},
  {32'h44dc01a2, 32'hc34d4ce3, 32'hc322096f},
  {32'hc4f8e586, 32'h418fd37c, 32'h41e8a138},
  {32'h43d4b464, 32'hc376dfd8, 32'hc2cdbc93},
  {32'hc4c433d6, 32'h438ed8ec, 32'h431342ec},
  {32'h44398d38, 32'h4235a010, 32'hc213ed54},
  {32'h43b3ca70, 32'hc2bf53c8, 32'hc26c7896},
  {32'hc4b87017, 32'hc3c61547, 32'h4295bf2e},
  {32'h4421f9d0, 32'h436e0286, 32'hc308cfe0},
  {32'hc49bc5c3, 32'h41c7f2ab, 32'hc355ffae},
  {32'h44cd3d71, 32'hc3c14e71, 32'h431c119a},
  {32'hc43af090, 32'h41c67c81, 32'h43025322},
  {32'h450d7537, 32'hc33d989e, 32'h428977f7},
  {32'hc4e3bc7f, 32'h41c8bc4b, 32'hc2d8ca01},
  {32'h4469844f, 32'h43139c6a, 32'hc2b04c95},
  {32'hc50c3d6e, 32'hc35395b2, 32'h4339404e},
  {32'h44bc57f9, 32'h43cb8a4d, 32'hc39e09ad},
  {32'hc3f941b0, 32'h4304008a, 32'h43aedda1},
  {32'h4352d894, 32'hc1c19c3a, 32'hc1ffd044},
  {32'hc51723ce, 32'hc37a0f5c, 32'hc29232ba},
  {32'h45115539, 32'hc39119d6, 32'h42b66c30},
  {32'hc3603c04, 32'h437ec092, 32'hc200ab5c},
  {32'h43f80b8d, 32'hc30e2067, 32'hc3f81894},
  {32'hc3d57a08, 32'hc3b65a32, 32'h4378eed3},
  {32'h446e071e, 32'hc2fde02a, 32'h439d2293},
  {32'hc4d2b780, 32'hc1bfb09a, 32'h434207fb},
  {32'h43b4802e, 32'h4292d890, 32'hc2a6a45e},
  {32'hc3da42a8, 32'hc1252d50, 32'hc3b4a147},
  {32'h445237f2, 32'hc2d8a4f4, 32'hc3623a44},
  {32'hc51301f3, 32'h424976ca, 32'hc21cb243},
  {32'h450ec158, 32'h42a9bdb8, 32'h4208c969},
  {32'hc40167b4, 32'h43ace19d, 32'h43a4dafb},
  {32'h442a205c, 32'hc3b76fae, 32'h42d64e5c},
  {32'hc4995fd8, 32'hc2baf863, 32'h435e6dd1},
  {32'h43cfbaef, 32'h423074e4, 32'hc36d8d24},
  {32'hc4531770, 32'h41928d88, 32'h43929302},
  {32'h4499acb0, 32'hc35e01d5, 32'hc358892c},
  {32'hc3312bcd, 32'hc381fac0, 32'h424f73c6},
  {32'h444fbc60, 32'h41a2d8fe, 32'h43e07f84},
  {32'hc48a9a9e, 32'hc3ac851b, 32'h4344260f},
  {32'h44f3dd82, 32'hc114c832, 32'h429fa1c1},
  {32'hc4572f47, 32'hc37594eb, 32'h4396f795},
  {32'h4513e0e8, 32'h43258389, 32'h410ecf1b},
  {32'hc3972d30, 32'h4331b8e3, 32'h42e95ac0},
  {32'h43ac9962, 32'h42e494c2, 32'h4336d840},
  {32'hc415e1e8, 32'h43c14f6e, 32'hc37caec1},
  {32'h4501c0af, 32'h43acdf35, 32'hc2c91035},
  {32'hc4a987ba, 32'h4391342d, 32'h4395a179},
  {32'h450771ba, 32'hc24035de, 32'hc2eb63da},
  {32'hc2fc68b4, 32'hc0dfde30, 32'h4323ad7e},
  {32'h453354d1, 32'h4364e2ae, 32'hc3241231},
  {32'hc51ff436, 32'hc3884bf9, 32'hc39e3096},
  {32'h4520f7d8, 32'h4245b1bf, 32'hc0d3f67e},
  {32'hc48af95e, 32'h43244fc4, 32'h4387d287},
  {32'hc4ed3ded, 32'hc3383752, 32'hc153c6e1},
  {32'h449a820c, 32'h4103cea2, 32'hc1838d5f},
  {32'hc3e3753c, 32'h43bc59af, 32'h43b3b756},
  {32'h44178604, 32'hc387bfa4, 32'h43a2a29e},
  {32'hc3d115bc, 32'hc3077591, 32'hc2bd7e67},
  {32'h445ed5de, 32'h4297acda, 32'h438d7bd6},
  {32'hc4479614, 32'hc2eb704a, 32'hc35f731e},
  {32'h435bd4b0, 32'h43b6aa50, 32'hc2e3b69d},
  {32'hc4552e6f, 32'hc2859970, 32'h42da9ef2},
  {32'h45203a8f, 32'h436746eb, 32'h432fb2f1},
  {32'hc4a3eba5, 32'h41699779, 32'hbf257033},
  {32'h44cf183a, 32'hc382e147, 32'hc39616b9},
  {32'hc4fc28e1, 32'hc210098a, 32'h43aa7a74},
  {32'h44a50bf3, 32'h43751fa6, 32'hc383e0ce},
  {32'h4459ed5e, 32'h43154459, 32'hc227d15c},
  {32'hc4c5c1ae, 32'hc3333c3e, 32'hc2fad7fc},
  {32'h45102705, 32'hc37ef1f5, 32'hc37a487d},
  {32'hc442001e, 32'hc34055f0, 32'h42a7bfde},
  {32'h44e2da07, 32'hc3860cda, 32'h437d794c},
  {32'hc4a4ba0e, 32'hc299f51a, 32'hc0d81d32},
  {32'h4433b2db, 32'h42fdf789, 32'h4218fea8},
  {32'hc3e2c5e0, 32'hc36934fe, 32'hc34f70f1},
  {32'h449c8919, 32'hc30167cc, 32'h43540558},
  {32'hc3558c23, 32'h428ec10d, 32'hc3684685},
  {32'h448a3764, 32'hc2c25964, 32'hc2e1f09e},
  {32'hc387db52, 32'h4387e9f0, 32'hc3540411},
  {32'h44f85ac2, 32'hc3967bb9, 32'hc2cb7f11},
  {32'hc419c54d, 32'h44169925, 32'h42b4c703},
  {32'h450fe226, 32'hc33af93c, 32'h43ab52f3},
  {32'hc4b67ddc, 32'hc2913735, 32'hc3243601},
  {32'h4487d40c, 32'h4350a401, 32'h43a7a8ef},
  {32'hc4ba3d17, 32'h435e078a, 32'h41335be7},
  {32'h445f5de8, 32'h43bc68eb, 32'hc401f76d},
  {32'hc3bf1390, 32'h4125c37e, 32'h429512ab},
  {32'h43d17f34, 32'h43645dc5, 32'hc2adeb08},
  {32'hc42c0a5d, 32'hc2bc5747, 32'h42165814},
  {32'h43f76a82, 32'h4214d707, 32'hc3e79163},
  {32'hc38b83c4, 32'h43a78701, 32'h42d866dd},
  {32'h43bbc474, 32'h42213143, 32'h4313f432},
  {32'hc4b4b100, 32'h4343af9a, 32'hc236abd4},
  {32'h448bbd4f, 32'hc31c7bbc, 32'hc398e77a},
  {32'hc4aeb219, 32'hc300d2cb, 32'h437cb146},
  {32'h4432f3b0, 32'hc2bef611, 32'hc3aa0278},
  {32'hc3cb9402, 32'h43e06118, 32'h43506cd2},
  {32'h43fbc184, 32'hc3405187, 32'h4308e9e9},
  {32'h42176840, 32'h4266e903, 32'hc2cf216f},
  {32'h43d3a5cd, 32'h4189ea8e, 32'h43c30538},
  {32'hc4e43f80, 32'h438a8b3e, 32'hc31c369a},
  {32'h4375f690, 32'h430449ad, 32'hc2b595f9},
  {32'hc48722bd, 32'hc4095797, 32'h4362d294},
  {32'h4484c8e0, 32'h42d39560, 32'h43b50512},
  {32'h4297d628, 32'hc2a8e86d, 32'hc2dbf652},
  {32'h441ea964, 32'h42a820e2, 32'h4184cd16},
  {32'hc507f568, 32'h40f6c76d, 32'h42cc9a91},
  {32'h4503d3f2, 32'hc2cb5228, 32'hc38b1e3f},
  {32'hc41fb708, 32'hc394ac80, 32'h438ae97d},
  {32'h4508f347, 32'hc33784c3, 32'h42f381ee},
  {32'hc41c4024, 32'hc268220c, 32'h41ba774a},
  {32'h4472f4e3, 32'h436c6bfa, 32'h42a59411},
  {32'hc2a8eb2e, 32'h422b8e69, 32'h42adba87},
  {32'h44a82eee, 32'hc3b7eb41, 32'hc30de71c},
  {32'hc4859fc2, 32'h4399a6dd, 32'h427d724c},
  {32'h431e7700, 32'h43b6680b, 32'h4345bb48},
  {32'hc4a0ca14, 32'h43392715, 32'h434114d9},
  {32'h44f196e8, 32'h403352a0, 32'hc34e4f96},
  {32'hc4a197cf, 32'hc1dc9370, 32'h43a1eafa},
  {32'h451484e3, 32'h43939410, 32'h4397347d},
  {32'hc51ac966, 32'hc021b3b0, 32'h43b01f53},
  {32'h441b6002, 32'h42ee7449, 32'h436b24e7},
  {32'hc51277bf, 32'h4305a945, 32'h430b1e68},
  {32'h44cb7050, 32'hc2e2c14d, 32'h4310368e},
  {32'hc4ba4cdc, 32'hc3cb4beb, 32'h43a0701c},
  {32'h441a2d94, 32'h43889784, 32'hc37dac82},
  {32'hc4e51c16, 32'h43018583, 32'h43b0832d},
  {32'h44ded0f7, 32'hc348816a, 32'h439b86d6},
  {32'hc4658918, 32'hc29602cd, 32'h43320e00},
  {32'hc32aa5b6, 32'hc2a72e34, 32'h43bcad08},
  {32'hc4878266, 32'h4244827a, 32'hc3473920},
  {32'h44e2bb6d, 32'h435ed0e4, 32'hc2d9257d},
  {32'hc4fcf747, 32'h43f89f7d, 32'h438cf1dd},
  {32'h44f54438, 32'hc3bc915c, 32'h43c7c9d3},
  {32'hc35b3318, 32'h42293e02, 32'hc3056fdd},
  {32'h44ef6241, 32'hc024a284, 32'h41b7763b},
  {32'hc4c16dd1, 32'hc3690406, 32'h43ac0e0f},
  {32'h44ba2f70, 32'h43cb2754, 32'hc36b052e},
  {32'hc4a6a372, 32'hc2dc2b2b, 32'hc3837042},
  {32'h44a714e0, 32'h4324ced5, 32'hc34ebdc9},
  {32'hc37dfb34, 32'hc3bd953f, 32'hc41816a6},
  {32'h44766406, 32'h43aa6f1c, 32'h43559336},
  {32'h42031500, 32'h42d9f854, 32'hc1d4dab5},
  {32'h44d8453b, 32'hc3af8c17, 32'hc156e770},
  {32'hc484c651, 32'hc2f2d71d, 32'h429135e3},
  {32'h44d21089, 32'h430171ff, 32'h4380cd8e},
  {32'hc4e80788, 32'hc313541d, 32'hc2b5bc6a},
  {32'h44a201fa, 32'hc1d004c5, 32'h42de9800},
  {32'hc4e75a06, 32'hc244762c, 32'hc36a6f4e},
  {32'h44148630, 32'h41c20214, 32'h41ce013e},
  {32'hc326b9f8, 32'h425b4dc7, 32'h4413aa8d},
  {32'h441c8952, 32'h423a74a0, 32'h431b4c8b},
  {32'hc4056bc1, 32'h42cb98e9, 32'h42c577c2},
  {32'h446d9c9c, 32'h43210d72, 32'h42842090},
  {32'hc4e3766b, 32'h43ad5edd, 32'hc0003e00},
  {32'h443dcb53, 32'h435d6ab8, 32'hc36cd898},
  {32'h425a76c0, 32'hc3be399a, 32'h41973879},
  {32'h44b8dab9, 32'hc324010c, 32'hc37d5ec6},
  {32'hc410714f, 32'h40436ece, 32'h438a4073},
  {32'h41e979a0, 32'hc3341877, 32'h42d22872},
  {32'hc3bcf501, 32'hc34584fc, 32'hc3be9655},
  {32'h4507d96f, 32'hc3531022, 32'h41db592e},
  {32'hc4a55d4e, 32'h42e3695b, 32'hc30fe586},
  {32'h43f56026, 32'h425f8964, 32'h42dd76e0},
  {32'hc42e71ba, 32'hc2b19dd2, 32'h43cd8a97},
  {32'h44387fd9, 32'hc06afcd2, 32'h4310f0de},
  {32'hc3f033d0, 32'h431f2bf8, 32'hc3644aa3},
  {32'h45141406, 32'h433c47c8, 32'hc33791d5},
  {32'hc512249b, 32'h431712b0, 32'h430c0dac},
  {32'h44582da6, 32'hc328c468, 32'hc29cc690},
  {32'hc50414d8, 32'hc28fcf43, 32'hc2f97b5e},
  {32'h440e56c8, 32'hc354ef66, 32'hc38df102},
  {32'hc3b8b23c, 32'hc397d488, 32'h4301639f},
  {32'h4429a15f, 32'hc3731946, 32'h42a8f554},
  {32'hc51e6834, 32'hc33ae5fc, 32'hc16fc9e6},
  {32'h44021a51, 32'hc2799f24, 32'hc393798b},
  {32'hc480c8ab, 32'h41c87f3b, 32'hc3c84f28},
  {32'h4467aeac, 32'hc2681866, 32'h416acd0c},
  {32'hc4e41098, 32'h42f7ae5a, 32'hc22e2991},
  {32'h44459c20, 32'hc314d9cf, 32'h43823699},
  {32'hc4cdb74d, 32'h43340c2a, 32'hc19b6766},
  {32'h43d8ae58, 32'hc37fa48e, 32'hc356475d},
  {32'hc49d3f44, 32'h41f253f9, 32'h43500dcf},
  {32'h4399f97f, 32'h4205b87d, 32'h42da3cdc},
  {32'hc462ed88, 32'h434f014c, 32'h43184311},
  {32'h44fab288, 32'hc3ad551b, 32'h4329bd3b},
  {32'hc4d31c74, 32'hc2284abb, 32'h4276dad5},
  {32'h43934120, 32'hc2b8fff4, 32'h4316adee},
  {32'hc4b78a07, 32'h43c00527, 32'hc203941f},
  {32'h44630b4e, 32'h43189776, 32'hc1fe4b71},
  {32'hc36fc8f2, 32'hc313cdc5, 32'hc3f9362f},
  {32'h4305a9a2, 32'hc33a5099, 32'h434af270},
  {32'hc382610d, 32'h43846a71, 32'h42e1fd42},
  {32'h43f86bdf, 32'h414bb268, 32'hc2c36ad9},
  {32'hc503751e, 32'hc2ed4291, 32'hc292ec9a},
  {32'h444086c6, 32'h41eea701, 32'hc38ab4e4},
  {32'hc49a249f, 32'h43335b3b, 32'hc2f7c1d8},
  {32'h4466380e, 32'h422e297c, 32'h4281e180},
  {32'hc43b6f1c, 32'hc3c0e741, 32'h4231ffa0},
  {32'h44d819de, 32'h42e1ba24, 32'hc33a2e40},
  {32'hc504d24f, 32'h427f3fb0, 32'h438b60f4},
  {32'h4414a9db, 32'h43f017ec, 32'hc33f65c3},
  {32'h425fbe78, 32'h42da8a44, 32'h43967512},
  {32'h450db30c, 32'hc0f934bc, 32'h42e6386a},
  {32'hc50a2809, 32'hc2bcf475, 32'hc33b4b0d},
  {32'h4493a904, 32'hc2bfd264, 32'h42fc6b43},
  {32'hc3e03a78, 32'h433da22b, 32'h42ea0b69},
  {32'h445ca678, 32'h43f8c63d, 32'h42c2a693},
  {32'hc4b66c21, 32'hc27dfc76, 32'h439144e9},
  {32'h43e5e078, 32'hc37e6ebe, 32'h423cee80},
  {32'hc4c261d0, 32'hc3c0af35, 32'hc1277890},
  {32'h44e0f316, 32'h412f9691, 32'hc1be2247},
  {32'hc2f4c320, 32'hc302562f, 32'hc341c50b},
  {32'h45181e12, 32'hc2d5796a, 32'hc3addd43},
  {32'hc48bd384, 32'hc31ae387, 32'h43e2f7ba},
  {32'h44f2e589, 32'hc2213279, 32'h437c4f99},
  {32'hc4be16ee, 32'h430140cb, 32'h429ba76b},
  {32'h44cfb6d0, 32'h42f05681, 32'h432f01ce},
  {32'hc4e0f13c, 32'hc2e27542, 32'h42780106},
  {32'h44bcb68b, 32'hc3cf4512, 32'h3fdb75dd},
  {32'hc5209433, 32'h434d16b1, 32'h42c064a8},
  {32'h44b6deeb, 32'h4333cb3f, 32'h43c29383},
  {32'hc4b03c05, 32'h433a6a34, 32'h4388f752},
  {32'h43fdcd88, 32'h4320bcc9, 32'hc35eaf18},
  {32'hc2307a80, 32'hbfb07dd0, 32'hc23a2ccf},
  {32'h41f24100, 32'h43d795be, 32'hc327b2a1},
  {32'hc4aae1cc, 32'h41c56d4a, 32'hc3f2bd73},
  {32'h44178ce2, 32'h42515a7e, 32'h43e61804},
  {32'hc40d8ac8, 32'hc300c233, 32'h42acad8a},
  {32'h44bba84e, 32'hc3ca04b7, 32'h434514b8},
  {32'hc320c580, 32'h43ffcaf8, 32'hc28f96c0},
  {32'h450d2be4, 32'h43137ed1, 32'hc4459216},
  {32'hc4de2f47, 32'h42d3f0c4, 32'h4210b645},
  {32'h4509e957, 32'hc322b90c, 32'hc2a18a12},
  {32'hc51a3b4a, 32'h439ebe9b, 32'hc2c447b4},
  {32'h450209fa, 32'h428e1a21, 32'h42ebcfd3},
  {32'hc2dfd2c1, 32'hc1cccf66, 32'h43bcc001},
  {32'h442ef260, 32'h43009a34, 32'hc3f55a85},
  {32'hc1a64280, 32'hc30a5369, 32'h421aa040},
  {32'h431f1d04, 32'h4296b8d5, 32'h4317217b},
  {32'hc4ae28b0, 32'h4268b3c9, 32'h4389e1e1},
  {32'h450f1fc8, 32'hc3c13556, 32'h415e4ca4},
  {32'hc1826280, 32'hc38b2d28, 32'hc1abf8da},
  {32'h44cc2db1, 32'hc2a3f12e, 32'hc33788fd},
  {32'hc485c27d, 32'h42bf6094, 32'hc3a87391},
  {32'h44bf3a42, 32'hc2eaf217, 32'h43f616f9},
  {32'hc51374d4, 32'h424f00ab, 32'h44408de1},
  {32'h448eeb1e, 32'hc390b6d3, 32'hc322b8c7},
  {32'hc483fa4e, 32'hc1d9d19e, 32'h429616fc},
  {32'h44921be0, 32'h40745d13, 32'hc263fe16},
  {32'hc248d136, 32'hc31f4079, 32'h438491db},
  {32'h416b4650, 32'h4187a939, 32'hc29a8a1c},
  {32'hc4431fa0, 32'hc1975d5a, 32'h43382fd9},
  {32'h417d2180, 32'h43bac157, 32'h42937238},
  {32'hc4172c5e, 32'hc31ecb22, 32'h4394cad8},
  {32'hc2328a36, 32'hc301f4f9, 32'hc2a1e8fc},
  {32'h42e3729b, 32'h436901f7, 32'h439eb2f4},
  {32'h44dc2168, 32'hc30c95bd, 32'h43b1ac0d},
  {32'hc4f34930, 32'h44153a79, 32'hc40daf99},
  {32'h4504f43a, 32'h41ba11ed, 32'h422413e7},
  {32'hc3408080, 32'h43aaba81, 32'hc327dad6},
  {32'h44d4e8d7, 32'hc14fd53a, 32'hc1ee0766},
  {32'hc404672c, 32'hc3aa5e7f, 32'hc356ddcb},
  {32'h450c3dfd, 32'hc3a7917e, 32'hc1f46d3a},
  {32'hc50e9adb, 32'hc2cd268d, 32'h4200555c},
  {32'h44c7bbb4, 32'h4182fca8, 32'hc38a5082},
  {32'h43f8f6a0, 32'h43f5c190, 32'hc33cd629},
  {32'h4431bd5e, 32'hc45d76dd, 32'h40e93f30},
  {32'hc4d8f9b6, 32'hc284bd9d, 32'hc30081f4},
  {32'h44435934, 32'hc2ee8e70, 32'hc2ac6179},
  {32'hc3a8e663, 32'h428a869e, 32'h4344a1bc},
  {32'h442cb53e, 32'h4071ae48, 32'hc3654466},
  {32'hc4835d2c, 32'hc36c476d, 32'h432c0e46},
  {32'h443efa8c, 32'hc1e9ac70, 32'h41d94058},
  {32'hc4249df7, 32'hc3bc79e6, 32'hc235073e},
  {32'h4422af92, 32'hc305816d, 32'hc339c14a},
  {32'hc4baf5d6, 32'h41a2db65, 32'hc38bdb5d},
  {32'h437a1290, 32'hc2f267e8, 32'h4101aaec},
  {32'hc4188049, 32'hc3d4c8f4, 32'hc2e88a14},
  {32'h43e5207c, 32'hc31e52f8, 32'hc387e2f2},
  {32'h41bfc8d8, 32'h4313a901, 32'h42864e20},
  {32'h446b4cf6, 32'h4227d0ae, 32'h43c5f43d},
  {32'hc490edb6, 32'h431eb225, 32'h43c47443},
  {32'h44b84ab5, 32'hc3d00efd, 32'hc3259fc6},
  {32'hc4fbddee, 32'hc1c0a94b, 32'h4290f15e},
  {32'h4485bbbf, 32'hc34c47fa, 32'h42ac797d},
  {32'hc4bb8c74, 32'h43076bfd, 32'h441793e2},
  {32'h443653bd, 32'hc2ae7484, 32'h42087370},
  {32'hc4f2962d, 32'hc381281d, 32'hc3365d11},
  {32'h42d27810, 32'hc32a715c, 32'h43195777},
  {32'hc4c6c05c, 32'hc1ede4d7, 32'hc2a77446},
  {32'h4510ff0b, 32'h428272a4, 32'hc32d2474},
  {32'h42ae8da0, 32'hc2ae5d33, 32'h436bdf9f},
  {32'h43d6e040, 32'hc3b0cd2c, 32'hc336b768},
  {32'hc3f8efca, 32'h438f3b4d, 32'h4344cdb9},
  {32'h44cbeffa, 32'hc30d0978, 32'h42b938d5},
  {32'hc4edbdc2, 32'h43ae083d, 32'h429f0521},
  {32'h43aa5d80, 32'hc1dbf93e, 32'hc2ba20da},
  {32'hc42f421c, 32'hc324dcfc, 32'hc219c4a2},
  {32'h44b067b7, 32'hc315a59b, 32'hc2f67084},
  {32'hc51cc2ed, 32'h43531caf, 32'h429af083},
  {32'h44df2b33, 32'h42ba411b, 32'hc2cbeb46},
  {32'hc4a62952, 32'h42eefb7a, 32'hc2fe8e62},
  {32'h4452b4f4, 32'hc3e1db37, 32'hc2aac3be},
  {32'hc509e77f, 32'h43e48221, 32'h42a82729},
  {32'h4453f898, 32'hc38253f0, 32'h431650f1},
  {32'hc4445f5c, 32'hc2fbbc34, 32'hc27a6c94},
  {32'h451bc098, 32'h4381906a, 32'hc2c18ab9},
  {32'hc4cbd63a, 32'h42d91f32, 32'h4356f1a2},
  {32'h450ae5cc, 32'hc2f904b0, 32'h43085ba8},
  {32'hc4cec246, 32'h428cb14c, 32'hc3b503da},
  {32'h44986ced, 32'hc308a9d4, 32'h43205299},
  {32'hc4e5d4d9, 32'h42aae95f, 32'hc301fcd0},
  {32'h447e43e5, 32'hc3817943, 32'h40d4ce54},
  {32'hc40afeca, 32'hc3e90671, 32'hc2eb2812},
  {32'h4469dd72, 32'hc27684e9, 32'h4366f21c},
  {32'hc35b84e4, 32'hc120b7a6, 32'h410a93f3},
  {32'h4441bc72, 32'h428faa87, 32'hc2ea25f4},
  {32'hc48a6fbe, 32'h43c2ffbb, 32'h4381b2bd},
  {32'h43dd93ea, 32'h438c37f6, 32'hc21ae7a8},
  {32'hc491ad7b, 32'h43923196, 32'h439ff083},
  {32'h42edca88, 32'hc3003245, 32'hc3105382},
  {32'hc42308aa, 32'hc243c3ae, 32'hc30f98c4},
  {32'h4513ccf0, 32'hc20c879c, 32'h42a9c451},
  {32'hc4dce1c3, 32'hc3b8485a, 32'h42c81a73},
  {32'h448affe2, 32'h42c67c88, 32'hc31b1c1a},
  {32'hc4764c62, 32'hc3858746, 32'h4362b7c3},
  {32'h4439ddaa, 32'h4320ebba, 32'hc1948ab0},
  {32'hc4b2c47e, 32'h429c8dd9, 32'h43abf7bc},
  {32'h43d0bd34, 32'hc24f01c7, 32'hc3104a52},
  {32'hc50d6c89, 32'hc387ee08, 32'h420bf34e},
  {32'h446a11f8, 32'hc319a9b4, 32'hc21cb4ef},
  {32'hc4df7872, 32'hc3293cff, 32'hc297cdce},
  {32'h44006098, 32'h3f730c38, 32'h4146fc88},
  {32'hc4f7a639, 32'h4301d138, 32'hc3ab9200},
  {32'h449f0e55, 32'h436f7e12, 32'hc333f61e},
  {32'hc2f52ac0, 32'h4359063d, 32'hc3b73717},
  {32'h43dd55fa, 32'h428e724b, 32'hc2c8a562},
  {32'hc51c555f, 32'hc35ac714, 32'h42685f06},
  {32'h43ce1260, 32'hc3849b04, 32'hc2889f48},
  {32'hc5017c06, 32'hc3323223, 32'h41a80eaf},
  {32'h43bc6e4e, 32'hc34a3d22, 32'hc2c6af6b},
  {32'hc3722cf4, 32'h428b5120, 32'hc364a184},
  {32'h452021b2, 32'hc35b1175, 32'h43bc21b5},
  {32'hc3edbf68, 32'h44148f37, 32'h410f29ed},
  {32'h4290a0ec, 32'hc3b4459b, 32'h43b92f7e},
  {32'hc4cf1b92, 32'hc0fdf0c3, 32'hc2b4fa72},
  {32'h44a311b5, 32'h413cea0a, 32'hc33c3428},
  {32'hc500b36f, 32'hc3387481, 32'hc32d1541},
  {32'h440fa0ec, 32'h432af4d4, 32'hc29372f4},
  {32'hc44f8a10, 32'h42c2bfb4, 32'h4306211a},
  {32'h44be3628, 32'hc35b710d, 32'hc34e6adc},
  {32'hc48f9998, 32'h43aac399, 32'h42fe7526},
  {32'h44b445ff, 32'hc38a6df2, 32'h42ea6bf0},
  {32'hc49accce, 32'hc2de5d2a, 32'h43e0f3b4},
  {32'h44a08166, 32'hc204f9e6, 32'h4211379c},
  {32'hc272a708, 32'h43159392, 32'h43a997c3},
  {32'h44c14915, 32'hc39879ad, 32'h438f8f35},
  {32'hc51565f0, 32'h43237cc0, 32'hc0bddc82},
  {32'h448f0190, 32'hc2ea93e4, 32'h4318c31a},
  {32'hc502a127, 32'hc356e00f, 32'h436538df},
  {32'h4507434d, 32'hc25efb04, 32'hc2e5e9be},
  {32'hc50c486e, 32'h42439b1d, 32'h411022a6},
  {32'h45097271, 32'hc2a595eb, 32'hc320b998},
  {32'hc5087b49, 32'h439c3ee4, 32'hc201600d},
  {32'h44d4f992, 32'hc37749de, 32'hc35f25f4},
  {32'hc48ef48e, 32'hc35461ed, 32'h4296d02f},
  {32'h445a3941, 32'h433ce705, 32'h42f35872},
  {32'hc4f2feec, 32'hc355d877, 32'hc30aed27},
  {32'h4492be9a, 32'h432900bd, 32'hc3017c7d},
  {32'h42cd0480, 32'hc3d7227d, 32'h42a3e67c},
  {32'h44994a70, 32'h427bd40a, 32'hc2c95634},
  {32'hc26327c0, 32'hc260dba7, 32'hc316bb92},
  {32'h44c67c2a, 32'h43ae3e6f, 32'hc3c5e1e8},
  {32'hc4f01903, 32'hc2a381e7, 32'h41ed1a3d},
  {32'h44e9872b, 32'h438f65d1, 32'h413d16c8},
  {32'hc5077e64, 32'hc1d6926b, 32'hc31ef8a3},
  {32'h43c984d2, 32'hc3cf6613, 32'h4337b6ca},
  {32'hc44ee680, 32'h421ecd09, 32'h43aeda8a},
  {32'h446a587f, 32'h4390fbc3, 32'hc1b117cd},
  {32'hc49f50f9, 32'hc382f156, 32'hc4016ce5},
  {32'h44a13d2a, 32'hc25ef334, 32'h43f07257},
  {32'hc4f09d65, 32'hc151c5f6, 32'hc269e188},
  {32'h44ebedf0, 32'h4382d4a8, 32'h4268a616},
  {32'hc5036fd8, 32'hc3916d54, 32'h43e2fad2},
  {32'h438bede0, 32'hc301152d, 32'h43951a93},
  {32'hc462740a, 32'h43215942, 32'hc3487c3f},
  {32'h45045140, 32'h40d34c0c, 32'h4349acea},
  {32'hc4fffaa4, 32'h41804a5c, 32'hc2d454d2},
  {32'h4415fecd, 32'hc35b6709, 32'h420bea79},
  {32'hc4d120a4, 32'hc0e9e418, 32'hc38e343c},
  {32'h45146bfa, 32'h436becde, 32'hc26f0071},
  {32'hc4b94ca1, 32'hc31996b3, 32'h43a6e646},
  {32'h44c7b969, 32'hc23bdd70, 32'hc3af0b77},
  {32'hc508be3a, 32'hc2edb172, 32'h441e9e51},
  {32'h44f7ac01, 32'h428a6f08, 32'h41c1193c},
  {32'hc4e13e06, 32'h4327defc, 32'h42696b10},
  {32'h43c5e969, 32'hc39351be, 32'h4318dbda},
  {32'hc4e12ccf, 32'hc1cbd9c2, 32'hc4108a1b},
  {32'h44a73d46, 32'h428adeb3, 32'hc2a89ec0},
  {32'hc3649178, 32'hc3138d37, 32'hc2b451db},
  {32'h44d893a4, 32'h43893222, 32'h421a09c2},
  {32'hc432b83c, 32'hc2020960, 32'hc26c783c},
  {32'h444d49c2, 32'h43a4be04, 32'hbfe34f0e},
  {32'hc2656f80, 32'h43af32b7, 32'hc3a3ee6f},
  {32'h4503fb65, 32'hc34ba228, 32'h4305e7c3},
  {32'hc4f31d6a, 32'hc2dd236b, 32'h418a2a1a},
  {32'h43341300, 32'h42cc05ca, 32'h42865f3c},
  {32'hc4a2b900, 32'hc3abc197, 32'hc3816c1d},
  {32'h44354889, 32'h4216f184, 32'h405e4830},
  {32'hc5020962, 32'hc340dd81, 32'h42154032},
  {32'h451d0e04, 32'h41c10ab8, 32'h43161370},
  {32'hc4c021fd, 32'h42e7d7e6, 32'h4308ee5f},
  {32'h4456364c, 32'hc34ac48d, 32'h4392018d},
  {32'hc4e3c224, 32'h42aa7174, 32'hc21eaa57},
  {32'h449b96ae, 32'hc39199a4, 32'h43024f4d},
  {32'hc4a07aca, 32'hc3319625, 32'h42dae2b8},
  {32'h450cb394, 32'hc1ce11cb, 32'h439340f6},
  {32'hc496cb6d, 32'hc3ce9201, 32'hc34ec39b},
  {32'h44b0eb69, 32'hc2083df4, 32'h4297d780},
  {32'hc3b92980, 32'h42c7a652, 32'hc13272fe},
  {32'h43aef32a, 32'hc2ecf6e4, 32'h436fbb20},
  {32'hc4e90d93, 32'hc2d6fb7d, 32'h4308b151},
  {32'hc01cdc00, 32'hc3296290, 32'hc21ae200},
  {32'hc3932104, 32'hc327d2ec, 32'h4200dd59},
  {32'h451bae47, 32'h4349dc71, 32'hc1ce2615},
  {32'hc4fe2be1, 32'h43acb36c, 32'hc28ee7a4},
  {32'h44d6f53c, 32'h431c980b, 32'h433f8736},
  {32'hc4fdfd18, 32'hc20ed423, 32'hc2b1ce31},
  {32'h44e20351, 32'h429af771, 32'hc3484944},
  {32'hc50c723f, 32'hc3dcd79c, 32'h408445a4},
  {32'h44f51562, 32'hc2868f03, 32'h428dae27},
  {32'hc398885c, 32'hc32d0c04, 32'hc1b59cb0},
  {32'h440e8b71, 32'h438c38c2, 32'h42ec83de},
  {32'hc391a754, 32'hc3a6e799, 32'hc2e4beb2},
  {32'hc4292a06, 32'hc2477db7, 32'hc2d7bbc4},
  {32'h43eb0444, 32'hc1255d08, 32'h43c03dfb},
  {32'hc4769385, 32'hc3cf02e9, 32'hc3ea8f6c},
  {32'h44bbdb34, 32'h4369818d, 32'h432e4a00},
  {32'hc4fce803, 32'hc3e47c8d, 32'hc2e76894},
  {32'h43ee6338, 32'h424057e1, 32'h439d47d5},
  {32'hc488be55, 32'h42d9eaf5, 32'hc2f06ad1},
  {32'h443fabde, 32'hc3d2e3ab, 32'h4393dba9},
  {32'hc4da1573, 32'hc36c7f81, 32'hc387b94d},
  {32'h45000766, 32'h4379d65a, 32'h43597d2e},
  {32'hc5020ffa, 32'hc33ddcf6, 32'hc2a8f988},
  {32'h45031bb0, 32'h43033eaf, 32'hc2560ee1},
  {32'hc39173cc, 32'hc29df5f7, 32'h42d9d080},
  {32'h4361a006, 32'h42b320b2, 32'h426425bf},
  {32'hc4c48c1a, 32'hc0cb0d6e, 32'hc3b9b6a0},
  {32'h45021798, 32'h43c6cf6f, 32'hc36d89b1},
  {32'h434cf532, 32'h4365698c, 32'h425c265a},
  {32'h4419ee2a, 32'hc3b63fa1, 32'h434dad5e},
  {32'hc3bdc430, 32'h43337de8, 32'h429bc9c6},
  {32'h448c3e40, 32'hbfd0dfae, 32'h42d3d8ee},
  {32'hc4054138, 32'h42a847a1, 32'hc368e9f4},
  {32'h44201558, 32'h4271ad00, 32'hc2b82384},
  {32'hc4ecb0fc, 32'h427fa1cd, 32'hc350871d},
  {32'h444d53de, 32'hc2c1ca53, 32'h4383aa23},
  {32'hc4f91fe4, 32'hc24273f0, 32'hc21873cb},
  {32'h4344a805, 32'hc42dda8d, 32'h43312b31},
  {32'hc50f05ae, 32'hc367aa1f, 32'h42a551e5},
  {32'h421e9f7a, 32'h438cf913, 32'h42fbc777},
  {32'hc301c1d0, 32'hc30c7018, 32'hc3f0ba97},
  {32'h44c61f3c, 32'hc40ae31e, 32'h4336d6c3},
  {32'hc46255da, 32'h429dbb38, 32'hc3c992a6},
  {32'h446151f8, 32'hc427932a, 32'hc2f7d37e},
  {32'hc5064d20, 32'h42134063, 32'h43bd4b2f},
  {32'h44b6274a, 32'h43ac60f4, 32'h43063e64},
  {32'hc50f1598, 32'hc1baa674, 32'hc3128771},
  {32'h418c75e0, 32'hc36ba5b7, 32'h4294186e},
  {32'hc4f08088, 32'h40c8e186, 32'hc354731e},
  {32'h443da796, 32'h43efb7ab, 32'hc24932fd},
  {32'hc4ebf5e6, 32'hc3240e57, 32'h43a644bd},
  {32'h44ace81d, 32'hc243bc25, 32'h42958989},
  {32'h444767be, 32'h42378615, 32'hc323bfe5},
  {32'hc48de60e, 32'hc2c2b505, 32'h427430bd},
  {32'h4419c909, 32'hc3ed335e, 32'hc3e5d2ff},
  {32'hc4bff6b2, 32'h42aeaacd, 32'h40850f70},
  {32'h44005a44, 32'hc114127c, 32'h436b3ff8},
  {32'hc4c918b0, 32'h43a220d0, 32'hc2dd496b},
  {32'h4483ea66, 32'h42ed2dbd, 32'h4380a58a},
  {32'hc3cbf44c, 32'h42e678c0, 32'hc322816b},
  {32'h440125cc, 32'h427bc38e, 32'h436c609d},
  {32'hc4811a93, 32'h43015697, 32'hc281075e},
  {32'h44dd35bc, 32'h435eb475, 32'hc370bfb8},
  {32'hc3d4b528, 32'h43bbb4e3, 32'hc3a4acb4},
  {32'h445c8a1e, 32'hc384fe9e, 32'h422e4df7},
  {32'hc4f622cd, 32'h4314fa51, 32'hc3311b4d},
  {32'h44de73b0, 32'hc3140291, 32'hc323bc22},
  {32'hc4818b24, 32'hc36ba2e4, 32'hc3b9b4c8},
  {32'hc515e55f, 32'h4108612e, 32'h438c9a45},
  {32'h44e0a9e2, 32'hc41c3162, 32'hc2e97f50},
  {32'hc30d6908, 32'h430c0e9f, 32'h42b5edde},
  {32'h442806a4, 32'hc322414c, 32'hc31a43bd},
  {32'hc506f039, 32'h4353663c, 32'hc40c6a4a},
  {32'hc51429ac, 32'h42c622f9, 32'h43c6cbeb},
  {32'h42f8722b, 32'h436f2894, 32'hc4059a9b},
  {32'hc4b27a74, 32'h4353cd3b, 32'h41444eec},
  {32'h450045b9, 32'h40b6d7f6, 32'hc2ca13c5},
  {32'hc42c595c, 32'hc3127234, 32'hc3246367},
  {32'h43ebcf78, 32'hc3193dff, 32'h44076789},
  {32'hc4eda949, 32'hc34c9544, 32'h42893871},
  {32'h45100117, 32'hc2fa21b9, 32'h43d00018},
  {32'hc4e8652a, 32'hc2f1bd22, 32'hc12d0364},
  {32'h449471b5, 32'h4380903a, 32'h4215a40c},
  {32'hc4f27d35, 32'hc1b6fc51, 32'hc313d473},
  {32'h4361b868, 32'h41be574e, 32'hc33c2ef8},
  {32'hc4de3c85, 32'h411c1df0, 32'hc22799ca},
  {32'h44a5662b, 32'h431adfae, 32'hc3936913},
  {32'hc511312f, 32'hc38d46f2, 32'h42954912},
  {32'h44dfdb00, 32'hc236c7ce, 32'hc2ade99a},
  {32'hc49bbe39, 32'h40774318, 32'h43401a80},
  {32'h4482cc09, 32'hc3683b70, 32'h44386cc6},
  {32'h42280a05, 32'h42092e77, 32'h42545941},
  {32'h440eff48, 32'h41c900af, 32'hc3e49e7d},
  {32'hc4428897, 32'h431814d8, 32'hc38a624d},
  {32'hc2246480, 32'h4322b654, 32'h43ad2eb2},
  {32'hc4d14abf, 32'hc243f3ef, 32'hc27556f7},
  {32'h442cb7de, 32'hc3b2d423, 32'h42ffbcaf},
  {32'hc4119192, 32'h42293910, 32'hc31abdf9},
  {32'h449d78df, 32'h4374aeee, 32'hc323e726},
  {32'hc50d3d0d, 32'hc360300e, 32'hc2e00f2c},
  {32'h449137d1, 32'hc31759e8, 32'h42d27ee0},
  {32'hc44a7966, 32'h404b2512, 32'h438d4013},
  {32'h4432cb1a, 32'h43465144, 32'hc3d578a6},
  {32'hc3adef68, 32'h434743a2, 32'h4311564c},
  {32'h44c3e1da, 32'h42faf581, 32'h4305b508},
  {32'hc4562d0e, 32'hc3487773, 32'hc33a33ca},
  {32'h448ac336, 32'h43be96db, 32'hc3480edb},
  {32'hc3808b9c, 32'hc315c870, 32'h4312ba76},
  {32'h44237688, 32'h43a3bf2f, 32'h439cb439},
  {32'hc385e762, 32'h43435320, 32'h432c6222},
  {32'h4511695c, 32'h430ae666, 32'h42af213e},
  {32'hc4e3b0e9, 32'hc39e2243, 32'hc20ad7f3},
  {32'h44917a02, 32'hc3118ba2, 32'hc2e385c0},
  {32'hc50944bd, 32'hc2c2ddc5, 32'h423f5589},
  {32'hc2ccee70, 32'hc330e3a9, 32'hc3060d39},
  {32'hc368cbe0, 32'h42e7bd5e, 32'hc173c6f4},
  {32'h4416667c, 32'hc3189833, 32'hc2847364},
  {32'hc426f80e, 32'h430577bd, 32'hc32a3f8e},
  {32'h444aaf00, 32'h43db5433, 32'h4218e5a0},
  {32'hc2d01b70, 32'hc31735e3, 32'hc2974257},
  {32'h450a05e0, 32'hc23a85df, 32'hc2a4c1de},
  {32'h4327a998, 32'hc43e07a2, 32'h430ca885},
  {32'h447b4ee6, 32'hc30e98ff, 32'h429c0150},
  {32'hc4cb95a6, 32'hc3d70a2a, 32'h42c94094},
  {32'h45120f84, 32'h43da6a5f, 32'hc3bc2048},
  {32'h44f82c92, 32'hc1d4eac6, 32'hc3a53405},
  {32'hc4cee1d8, 32'h422900d9, 32'h40f97c9c},
  {32'h4453a14c, 32'h42537d4c, 32'hc3a872a0},
  {32'hc46ea9f6, 32'h422a615c, 32'hbf328a20},
  {32'h443fec3c, 32'hc2659568, 32'h43938acb},
  {32'hc4a0dd1a, 32'hc30c70ed, 32'hc1ab658c},
  {32'h43260650, 32'h41bc372e, 32'hc3b7f467},
  {32'hc4496186, 32'hc280fc56, 32'hc2bc6979},
  {32'h44991b56, 32'h435a4974, 32'hc27f90a0},
  {32'hc3d20013, 32'h437e0df1, 32'h4324890a},
  {32'h43762da8, 32'hc2a61be1, 32'h42ca71be},
  {32'hc4f1db1d, 32'hc29b565c, 32'h431d1067},
  {32'h4487229e, 32'h43894985, 32'hc3bd544d},
  {32'hc3c931e8, 32'hc31deb2e, 32'h43490810},
  {32'hc465ea8a, 32'hc3656bb0, 32'h43685dc7},
  {32'h448653ec, 32'h42a6668a, 32'h436d5900},
  {32'hc2741188, 32'h43859db4, 32'hc39f58be},
  {32'h448937d4, 32'h438d8975, 32'hc2856051},
  {32'h42739600, 32'h4339584a, 32'h43fa9beb},
  {32'h4505f0f2, 32'hc2d5f1aa, 32'h420091a3},
  {32'h42158be8, 32'hc3b0ae03, 32'h435d608a},
  {32'h44b32a19, 32'h4323618e, 32'h43b2cfbb},
  {32'hc4273b9e, 32'hc2442fa0, 32'h439c667b},
  {32'h4384f724, 32'hc2edd673, 32'h43ae1a5a},
  {32'hc3d640a2, 32'hc39e6e72, 32'hc2cdfb3c},
  {32'h44ebd186, 32'h428dbfc0, 32'h43a7dfda},
  {32'hc400d61c, 32'hc335b5f8, 32'h42c608c7},
  {32'h44446d3e, 32'h42df45c5, 32'h429dccae},
  {32'hc36705bc, 32'hc387f2e5, 32'h43a2658e},
  {32'h43d8bf48, 32'h40702050, 32'h42f462ee},
  {32'hc383a030, 32'hc37cb104, 32'hc39ed7f1},
  {32'h44a2fd28, 32'h416c99cd, 32'hc38d0c91},
  {32'hc42be952, 32'h4378be43, 32'h4208e344},
  {32'h44d6770c, 32'hc35d913a, 32'hc37f183b},
  {32'hc4fdf162, 32'h431a6855, 32'hc3738638},
  {32'h44238a13, 32'hc2d759c6, 32'h43a02f67},
  {32'hc3d8b2dc, 32'hc2ebd00c, 32'hc32d96c1},
  {32'h42879678, 32'hc3a5f1dd, 32'hc1fb829b},
  {32'hc4e70413, 32'hc121994c, 32'hc1ec731e},
  {32'h443bcbca, 32'hc3345aac, 32'h420433a8},
  {32'hc50fce72, 32'h434501da, 32'h428969ac},
  {32'hc30e54ec, 32'hc404a6e8, 32'h43ab2ed7},
  {32'hc47d2776, 32'hc3842ff6, 32'hc2fc722d},
  {32'h43cff70e, 32'h42241645, 32'h43ab4c90},
  {32'hc46fac62, 32'hc2d0ac36, 32'h425e1b0d},
  {32'h434436a0, 32'hc3730b8c, 32'hc22e7ebb},
  {32'hc4c3407d, 32'hc2cf6544, 32'hc348e9ab},
  {32'h44d02111, 32'hc2be2b0b, 32'hc335f3cc},
  {32'hc49ec945, 32'h404265b6, 32'hc2e1131c},
  {32'h4515184d, 32'h43be88ff, 32'hc3e13068},
  {32'hc40b7984, 32'h43449502, 32'hc30b0aef},
  {32'h4518b46a, 32'h41ede0c3, 32'hc2d16200},
  {32'hc4c6114d, 32'h44041e8f, 32'h43bda320},
  {32'h44dbd2f6, 32'h43627c56, 32'hc2ebbf0f},
  {32'hc4f2d56d, 32'hc3569cb7, 32'h419ec35f},
  {32'h43a6e290, 32'hc3575a28, 32'hc325ebff},
  {32'hc28f3e40, 32'h42d9b957, 32'hc10a5c9f},
  {32'h449aeaea, 32'h4437a2cd, 32'h43ab217a},
  {32'hc44451b7, 32'h430889a2, 32'hc3191321},
  {32'h44c6d84c, 32'h42ec2d9c, 32'hc128c139},
  {32'hc39ac632, 32'hc398faea, 32'h4256bf7f},
  {32'h4186bb00, 32'h432a9b41, 32'hc3c25fa1},
  {32'hc4ca5c50, 32'h419786d4, 32'h43042147},
  {32'h44924ef3, 32'h4153197c, 32'hc3383702},
  {32'hc445f83e, 32'h41515744, 32'hc2afdf79},
  {32'h446289bc, 32'h429b07df, 32'h429d1795},
  {32'hc4127b97, 32'h4248d557, 32'hc3242e1d},
  {32'h444a6db2, 32'hbea1c690, 32'h40cb7059},
  {32'hc500677f, 32'h4101ee29, 32'h43984cfd},
  {32'h44aceaf5, 32'h439d3bc7, 32'hc3620b82},
  {32'hc50b4f1d, 32'h43be1466, 32'hc3570432},
  {32'h44cb0568, 32'h43dce10a, 32'hc3839cac},
  {32'hc4dd8bba, 32'h432085f0, 32'hc32fbac9},
  {32'h4224ef48, 32'h43e38bed, 32'h4384e4e6},
  {32'hc4d0a17c, 32'hc2fa8757, 32'h42a59397},
  {32'h443c0554, 32'hc3055961, 32'h42e3e5ec},
  {32'hc4103e22, 32'h420d3851, 32'hc32083bb},
  {32'h44f0f126, 32'h4375226a, 32'h4311a0d6},
  {32'hc3f43580, 32'h432e6285, 32'h43aa3e39},
  {32'h44c2c8cf, 32'h43ea1187, 32'h42bb53eb},
  {32'hc2ded700, 32'h4311524d, 32'hc2210f64},
  {32'h451173a0, 32'hc2aee990, 32'hc3984170},
  {32'hc49d8c68, 32'hc3bb5656, 32'h3f800aed},
  {32'h44c47fe1, 32'h42610d39, 32'h3ff72098},
  {32'h4318a990, 32'hc32204b1, 32'hc3a5a5ba},
  {32'hc3059520, 32'hc2a5a128, 32'h43158812},
  {32'hc2647380, 32'h42deb270, 32'h43e21755},
  {32'h439e88b0, 32'h43879bc4, 32'h42b298bb},
  {32'hc4c01517, 32'h420d7305, 32'h42f49529},
  {32'h43ea79d6, 32'hc3bee0c6, 32'hc32b4266},
  {32'hc4dea191, 32'hc1ec9bcc, 32'hc2bb6942},
  {32'hc2bf8190, 32'hc37e3ba7, 32'hc3ac1e48},
  {32'hc485838f, 32'h43893377, 32'hc30173aa},
  {32'h43289d4a, 32'hc3c7aa31, 32'h42fe6d28},
  {32'hc417fb5f, 32'h43c7598a, 32'hc35efe2c},
  {32'h4479ee14, 32'hc32c600b, 32'h43a054d7},
  {32'hc5190f21, 32'h42196438, 32'h4330b03b},
  {32'h4486d735, 32'h4300e8f2, 32'h43555d3e},
  {32'hc3ab994c, 32'h4314d48b, 32'hc3931cd4},
  {32'h43c909b2, 32'h438148c4, 32'h43c8a6b2},
  {32'hc4bbf9c6, 32'hc35bb853, 32'hc2ff783c},
  {32'h43f5b038, 32'hc3a3df89, 32'hc0c54d44},
  {32'hc4c1dd49, 32'hc2219abd, 32'h41720a36},
  {32'h44fb9dee, 32'h4370fa5e, 32'hc37c2094},
  {32'hc4f99011, 32'h44005eea, 32'hc3a5b15b},
  {32'h43cc3340, 32'hc0f49828, 32'h44071d8a},
  {32'hc5010db2, 32'hc2ebbca4, 32'hc3e0efb0},
  {32'h44c75b7d, 32'hc1439b6f, 32'hc3956639},
  {32'hc4521554, 32'hc29ec586, 32'h43aeaeed},
  {32'h44c605c4, 32'h43a6f8f8, 32'hc3580156},
  {32'hc4a47b28, 32'h43d0878c, 32'hc34b1cc1},
  {32'h439fa9b0, 32'hc33f6285, 32'hc3fd7c9a},
  {32'hc4894056, 32'h43afb58f, 32'h43b303ab},
  {32'h44017798, 32'h41be1d60, 32'hc39a8f64},
  {32'hc2c1a190, 32'h43453ad2, 32'hc34c6668},
  {32'h45137b34, 32'h437e3a11, 32'hc2c0d962},
  {32'hc506b08e, 32'hc39a6d90, 32'h43202017},
  {32'h442ed694, 32'h43972711, 32'h424ac1b8},
  {32'hc4236fa6, 32'h435f4fe7, 32'hc33969d8},
  {32'h44d10ac8, 32'h43827834, 32'hc19d4c81},
  {32'hc4227746, 32'hc307e888, 32'hc0455b48},
  {32'h44d5fc2b, 32'h443388e5, 32'hc2480eb9},
  {32'hc4c3b07e, 32'h43688a60, 32'hc3c7a2ef},
  {32'h45127284, 32'h424ab966, 32'hc389fe4b},
  {32'hc21b2288, 32'h429afb46, 32'h4303c8bf},
  {32'h443574ef, 32'hc298ee20, 32'h439a9fbe},
  {32'hc4ea42ca, 32'h43f8f74e, 32'h43a49d45},
  {32'h43fa3ea4, 32'h43d988a4, 32'h43cce46f},
  {32'hc48e9bee, 32'h410a7e73, 32'hc24c18b3},
  {32'h442c685a, 32'hc1673691, 32'h419d1ed8},
  {32'hc4d34a6c, 32'hc2109471, 32'h42f358e5},
  {32'h4458852e, 32'h438b5277, 32'hc2f534ce},
  {32'hc4bb65b3, 32'h43b4aff2, 32'hc30f4201},
  {32'h442c721a, 32'hc31f8e2b, 32'hc0e8e4c9},
  {32'hc3757a68, 32'hc3a856e1, 32'h430ed808},
  {32'h44367d70, 32'h42af3c66, 32'hc303657b},
  {32'hc44099ca, 32'hc306f861, 32'hc31c1556},
  {32'h44b6c664, 32'h42c7c00a, 32'hc1c61eab},
  {32'hc3d946f6, 32'hc2d21905, 32'h42387716},
  {32'h44e9c427, 32'hc1933497, 32'hc22cedb2},
  {32'hc2ac5df1, 32'h4303e601, 32'h439284a3},
  {32'h436e9858, 32'hc2fe23bf, 32'h436f891b},
  {32'hc4ea1c8a, 32'hc31569ef, 32'hc0bb3328},
  {32'h444930c6, 32'h42e7537a, 32'hc300e4d7},
  {32'hc4761543, 32'hc3139cce, 32'hc1773d8f},
  {32'h448db46c, 32'h421c9eef, 32'hc28f23eb},
  {32'hc4e0b8d9, 32'h3e8aa360, 32'hc2806493},
  {32'h452a500d, 32'hc3be7700, 32'h4441388b},
  {32'hc4f0b846, 32'h43387a06, 32'hc2a1196e},
  {32'h44ad7cbf, 32'h4261855b, 32'h42d382e1},
  {32'hc484f02a, 32'hc2ff8b60, 32'h426cb0e1},
  {32'h45084f66, 32'h436c6302, 32'h439332e5},
  {32'hc4a2b2a4, 32'hc34806f9, 32'h436be125},
  {32'h4493ce2a, 32'hc38532ee, 32'h42a3af56},
  {32'hc3a9607a, 32'h43a3b064, 32'hc2c2be57},
  {32'h4510db32, 32'hc1c13f04, 32'h428f44ae},
  {32'hc51ae715, 32'hc361d906, 32'h437e689b},
  {32'h44bcfd5b, 32'hc1f12b7a, 32'hc37109c1},
  {32'hc4133bb6, 32'h42ded2c8, 32'hc190310f},
  {32'h45065d84, 32'hc291cc55, 32'h4265c1f5},
  {32'h4219492e, 32'hc24441dc, 32'hc3dc609b},
  {32'h452a3f48, 32'h4367fd06, 32'h436aad51},
  {32'hc4b5173b, 32'h43cda348, 32'h4382c371},
  {32'h45123fc2, 32'hc34bfbce, 32'hc2e04232},
  {32'hc40de668, 32'hc1838508, 32'h423fc5c8},
  {32'h44d94fcd, 32'h42d8eebe, 32'hc3f024e5},
  {32'hc36ecec0, 32'h42204d87, 32'h43bc58e7},
  {32'h449d2410, 32'hc39566c3, 32'hc1e7a54d},
  {32'hc4fce441, 32'h42825cc9, 32'hc37400e5},
  {32'h414d0900, 32'h436b73ea, 32'hc335a272},
  {32'hc44da933, 32'hc356ed53, 32'hc2eeaa3e},
  {32'h44a6b99a, 32'hc18ca027, 32'hc38825fa},
  {32'hc4ed31bb, 32'h43310eab, 32'hc33fa2e8},
  {32'h444acd26, 32'hc2b94790, 32'hc32ef76c},
  {32'hc4bd7ff0, 32'h433b817a, 32'hc393c05c},
  {32'h44c49c43, 32'hc27eee2d, 32'hc34ba17c},
  {32'hc4dead4f, 32'hc3881d24, 32'hc2f0c542},
  {32'h45158915, 32'hc0f8e7e5, 32'h43113075},
  {32'hc4f2513b, 32'h429e9e87, 32'hc32ac44f},
  {32'h4413e500, 32'hc32cd992, 32'h440ac266},
  {32'hc4dd74f6, 32'h438286c1, 32'h40395f91},
  {32'h4466c476, 32'h43492d4b, 32'h42600323},
  {32'hc329ae00, 32'hc28a42e9, 32'hc3bb91de},
  {32'hc1632380, 32'h441603ab, 32'hc34fec4f},
  {32'hc4c21260, 32'hc410a4cd, 32'hc3c7e7a7},
  {32'h440775f0, 32'hc28fd83a, 32'h420cca5b},
  {32'hc445deba, 32'hc2c9fe78, 32'h432a72a6},
  {32'h431c7c90, 32'hc384ee33, 32'h43b3ed71},
  {32'hc4c019f4, 32'hc30c4847, 32'h43ac745b},
  {32'h44cbf68c, 32'h43b249c7, 32'h4225f55c},
  {32'hc4cc104a, 32'h43109c26, 32'h429650a1},
  {32'h44f20358, 32'hc319d83f, 32'hc3228c9b},
  {32'hc502573c, 32'h4332c652, 32'h423ae8eb},
  {32'hc3ebf59c, 32'hc1e8cc33, 32'h4288eef4},
  {32'hc3a705b8, 32'hc1c0130c, 32'h40ee492d},
  {32'h444eebea, 32'h43bd5707, 32'h43cdfad8},
  {32'hc51f5cb0, 32'hc41e14b1, 32'h42cf64b4},
  {32'h44e63b4d, 32'h435923fc, 32'h43642732},
  {32'hc443204d, 32'hc38e534c, 32'hc399b9ba},
  {32'h44c05496, 32'hc30ab08d, 32'hc2d07beb},
  {32'hc49c00d0, 32'hc3b1da2f, 32'hc367ef35},
  {32'h439170f8, 32'h42d5ab5d, 32'hc28fc5cb},
  {32'hc3d82558, 32'h42a06923, 32'hc3dbbec5},
  {32'h4501e367, 32'h439713ca, 32'hc3b5f735},
  {32'hc2f29ce0, 32'hc225ba39, 32'hc21a2711},
  {32'h445c25a2, 32'hc2ff450d, 32'hc1d2bf46},
  {32'hc44bc9e0, 32'hc318aceb, 32'h42ee9c0b},
  {32'h44d1504a, 32'hc0215c36, 32'hc386a4f1},
  {32'hc43129bc, 32'h426c5c18, 32'hc2b1b8d6},
  {32'h44fb8018, 32'h433f6878, 32'h43631a67},
  {32'hc5043d34, 32'hc39c1f8b, 32'h43c12658},
  {32'h44e0a57f, 32'hc358ed73, 32'hc254c493},
  {32'hc3c16ff0, 32'hc3a8484d, 32'hc30d3ee6},
  {32'h44ad302c, 32'hc3380ddd, 32'hc191cac2},
  {32'hc48b4731, 32'hc1149d40, 32'h4310121c},
  {32'h43ccc448, 32'h42025ae8, 32'h4293b2b0},
  {32'hc50f8ea8, 32'h429ceb96, 32'h44094d91},
  {32'h44d8a8c4, 32'h42ed7c4b, 32'hc291cdfa},
  {32'hc37b05f8, 32'h40ec5966, 32'hc362e054},
  {32'h44ba6db8, 32'hc21c89cf, 32'h42e503d9},
  {32'h42878480, 32'hc2d38390, 32'h437f9174},
  {32'h44be2fde, 32'h42593c7a, 32'h43aef45a},
  {32'h44747392, 32'h431a9f9c, 32'hc1d63651},
  {32'hc4abf7b8, 32'h42514ada, 32'h41b940bc},
  {32'h446a019a, 32'h400cb2f8, 32'h426b2abf},
  {32'hc49ea85f, 32'h432c720e, 32'hc3c5706b},
  {32'h45226c6b, 32'h43880d67, 32'hc3c6256c},
  {32'hc435f092, 32'hc3bc2687, 32'h43ce73f5},
  {32'h44b68815, 32'hc33c14ca, 32'h428240ce},
  {32'hc3a35b76, 32'h432c6c60, 32'hc110f1ca},
  {32'h44e3ca5c, 32'h42784d24, 32'hc2f77e2d},
  {32'hc486f698, 32'h40e94574, 32'h42f57b90},
  {32'hbffe1400, 32'hc32cf245, 32'h432e2fac},
  {32'hc315ae94, 32'h4387c19a, 32'hc34569aa},
  {32'h453185ff, 32'h4395f6ea, 32'h42b27f72},
  {32'hc503932e, 32'h432ffa03, 32'h4234864c},
  {32'h44b93ea8, 32'h41b3a890, 32'hc39c5892},
  {32'hc4b9b8b7, 32'h41b0256c, 32'hc33e3bb7},
  {32'h450211d6, 32'hc29ac636, 32'hc3392d12},
  {32'hc4f80bc0, 32'hc331ea9c, 32'h43eff1ad},
  {32'h438f08c2, 32'hc32489f0, 32'h4316d46d},
  {32'hc330a918, 32'hc3e19161, 32'hc3d6eeb2},
  {32'h44522d3e, 32'h433f6216, 32'hc2d6036e},
  {32'hc4ccab1a, 32'hc40a2443, 32'hc28ad2e9},
  {32'h43d325c8, 32'h43496336, 32'h434a9fb9},
  {32'hc337b1ac, 32'hc38468a6, 32'hc2bbb830},
  {32'h441a7667, 32'hc36b6e44, 32'h433c1e04},
  {32'hc4d83463, 32'h43272062, 32'hc3aa01a2},
  {32'h44b685ba, 32'h4294ce65, 32'h429a30a4},
  {32'hc5180200, 32'h4385bd57, 32'h43d06d92},
  {32'h4481a149, 32'h438366c1, 32'h42d96ad4},
  {32'hc4a7029e, 32'h43e6604b, 32'hc3042444},
  {32'h44ed7225, 32'h4386cfdc, 32'h439fa886},
  {32'hc499e940, 32'h4350e46c, 32'hc2e668af},
  {32'h44f6f7e1, 32'hc29bcc7b, 32'h435b3b2d},
  {32'hc488a528, 32'h4381a2e8, 32'hc36d4f9f},
  {32'h4499fac0, 32'h431eeb2a, 32'h4324e125},
  {32'hc4333846, 32'hc2c5d8fe, 32'h43dc3dd4},
  {32'h44a3eb82, 32'h431bf1b6, 32'hc3a04160},
  {32'hc26dfcc0, 32'hc1d7e1bf, 32'h44081c60},
  {32'h436fe0c2, 32'h431fa3aa, 32'hc329df57},
  {32'hc49c04c4, 32'hc26c53be, 32'h42355753},
  {32'h450a66ad, 32'h43183ce9, 32'h41690b4e},
  {32'hc52d090f, 32'hc3691c09, 32'h43142df2},
  {32'h4505bf59, 32'h42974c20, 32'h412429cd},
  {32'hc4d7d91d, 32'h428e2f9c, 32'hc260fa60},
  {32'h444dc662, 32'h434a0ca7, 32'hc42256af},
  {32'hc4daf273, 32'hc41161ae, 32'hc35bc342},
  {32'h44aeb3f4, 32'h4344a57a, 32'hc283898a},
  {32'hc50bcdf2, 32'h41fa8970, 32'h43ae520e},
  {32'h445ea706, 32'h43990b83, 32'h41816f52},
  {32'hc4b05ec9, 32'hc327c3d2, 32'h42c427a2},
  {32'h444598f8, 32'hc3533276, 32'h43164cd2},
  {32'hc29c91d6, 32'hc35bbca6, 32'h401a030b},
  {32'h446e2a87, 32'hc30f8eec, 32'hc354ec8d},
  {32'hc4f4ede5, 32'hc300c050, 32'h43cbeca8},
  {32'h44b6ee95, 32'h4307aba1, 32'h42950a5f},
  {32'hc2a07f80, 32'hc3a8ca1c, 32'h43cd480c},
  {32'h44b0f7b4, 32'h43fb5b74, 32'hc30c791f},
  {32'hc44b5839, 32'hc395c133, 32'h42ac2f1d},
  {32'hc49177bc, 32'hc387a94c, 32'h42c9d8a6},
  {32'h44e361b4, 32'hc332a947, 32'h42b9b14c},
  {32'hc4ba74e2, 32'hc357484a, 32'h423120e6},
  {32'h44bfbd9a, 32'hc2ca776d, 32'hc3d54ee3},
  {32'hc30b82e3, 32'h42e611d0, 32'h4251c81c},
  {32'h44feff47, 32'hc1a21f46, 32'hc32b2821},
  {32'hc4ff0c37, 32'h4312a5ef, 32'hc39bf0c1},
  {32'h44325028, 32'hc31f1b53, 32'hc3fb6ad4},
  {32'hc3e17204, 32'h42cd58a3, 32'h438681b5},
  {32'h44aab238, 32'hc37d58e4, 32'h41b92bfb},
  {32'hc49267f8, 32'hc3a60f35, 32'h4354df1f},
  {32'h45064498, 32'hc1e230e0, 32'hc2a26dec},
  {32'hc49eb7a3, 32'hc32e56bc, 32'hc3a364b3},
  {32'h44aa528e, 32'h43e02a5f, 32'hc33b62a0},
  {32'hc50813ec, 32'h42e9f4ca, 32'h42eab98c},
  {32'h44b644a1, 32'hc285e679, 32'hc3277810},
  {32'hc2b6d8c2, 32'h440655c2, 32'h43a4a13a},
  {32'h4403a4d4, 32'h42756c63, 32'hc22006f4},
  {32'hc4577dd8, 32'hc27f2c86, 32'h43e13f08},
  {32'h44595df6, 32'h431698e9, 32'hc287ea7b},
  {32'hc45d803b, 32'hc2d20c08, 32'h4338c2b0},
  {32'h44ca14e5, 32'hc2e37711, 32'hc3a06fee},
  {32'hc47f12b7, 32'hc39ca92d, 32'hc294271d},
  {32'h4500f644, 32'hc3afe4b0, 32'hc26a757f},
  {32'hc4d6db5c, 32'hc2e080a6, 32'h42fe4e8f},
  {32'h4454ea70, 32'h43203a9c, 32'hc2add4a0},
  {32'hc40e8c7e, 32'hc31ece5f, 32'hc299f70d},
  {32'h44cd08b6, 32'h41f499a3, 32'hc2512b99},
  {32'hc479a95a, 32'h42da9c61, 32'h4390f264},
  {32'h43a695f0, 32'hc3f3b02f, 32'hc438aa95},
  {32'hc5136eee, 32'h42eb09b4, 32'h438cb1e2},
  {32'h44ea64f0, 32'hc271e614, 32'h441a77c8},
  {32'h44a70741, 32'h43001e51, 32'hc1dc100b},
  {32'hc3c55f98, 32'h41a52044, 32'h43c7a844},
  {32'h447caa0c, 32'hc3964686, 32'hc279419a},
  {32'hc49463fe, 32'h43a319ff, 32'h421e1751},
  {32'h450e0be8, 32'hc37349ed, 32'hc3902ff5},
  {32'hc3f99cf5, 32'h430023f1, 32'h42fe9728},
  {32'h448ffacb, 32'hc3d1f71c, 32'hc32565cc},
  {32'hc3e654c8, 32'hc2ceffe8, 32'h43aa5af7},
  {32'h433a2c10, 32'hc38db44f, 32'hc26e8f5f},
  {32'hc4a5ac22, 32'h3fdca830, 32'hc187516d},
  {32'h444d86de, 32'hc3042f87, 32'h432f6b01},
  {32'hc49b4a76, 32'hc32e7dc4, 32'h43d436da},
  {32'h44f4bc4a, 32'hc33cdaa1, 32'h41b2b9d9},
  {32'hc4a31399, 32'h43dadc81, 32'hc316b8d0},
  {32'h4421a2d2, 32'hc3143946, 32'hc2a6f706},
  {32'hc429271d, 32'hc2fdb8ba, 32'h42b17c15},
  {32'h44b4a552, 32'hc17e4b4b, 32'hc310e7b3},
  {32'hc38bded0, 32'h43a02ae2, 32'h42a3e412},
  {32'h445a2cc0, 32'h43b47532, 32'hc15090da},
  {32'hc49824ac, 32'h42e21259, 32'h432a6eea},
  {32'h4501985e, 32'h440cd52e, 32'hc2c3b094},
  {32'hc4e59b54, 32'hc32c9d82, 32'h434c9333},
  {32'h44838c47, 32'hc2e27227, 32'h410f1ad9},
  {32'hc480a4dd, 32'hc364ee2a, 32'hc228ad82},
  {32'h450dd40e, 32'hc271c25b, 32'hc2b4ff00},
  {32'hc4cbf16a, 32'hc3c23e26, 32'h438bbb05},
  {32'h441b5d23, 32'h42d4ea21, 32'h42cc5c01},
  {32'hc48c53b3, 32'hc28765f7, 32'h4392295d},
  {32'h441ba5de, 32'hc35c2b60, 32'hc40fc391},
  {32'hc3f04090, 32'h4244f6eb, 32'hc37c7e63},
  {32'h44ad9730, 32'hc3a7299b, 32'h4297c886},
  {32'hc43243d2, 32'h4375af48, 32'hc1f9ba4c},
  {32'h4392a4fc, 32'h4323434a, 32'hc3a5be45},
  {32'h42b702c4, 32'hc28fd716, 32'hc2a23f33},
  {32'h4409c84e, 32'h415344cc, 32'hc11f8056},
  {32'hc49bf548, 32'hc1108f3c, 32'h42dec38a},
  {32'h44f0063a, 32'hc3755e80, 32'hc30a2922},
  {32'hc4a394fa, 32'hc1b99abc, 32'hc33e7dcb},
  {32'h44d75e1a, 32'h4327f47b, 32'hc348b706},
  {32'hc4f739ae, 32'h43889520, 32'h436dc312},
  {32'h4482dad5, 32'hc37eb54f, 32'hc3c28ba5},
  {32'hc4ed294b, 32'h43a87d53, 32'h42bcd61c},
  {32'h44af7fa4, 32'hc2fc02ee, 32'h4397b6ac},
  {32'hc4cb6117, 32'hc431ae57, 32'hc1736720},
  {32'h445fdbb6, 32'hc00c5b17, 32'h425f0d74},
  {32'hc50f1a8c, 32'hc4080006, 32'hc3899ddc},
  {32'h450e2428, 32'h43861e14, 32'hc0bc1d1f},
  {32'hc4fefa25, 32'h43d3a653, 32'hc2740e7e},
  {32'h4491fd4b, 32'h43d64e55, 32'hc3196854},
  {32'hc4a7b811, 32'h42e17f3d, 32'hc37a2f98},
  {32'h4484bbe3, 32'h429e1bcf, 32'h43c96776},
  {32'hc4f2f4ed, 32'hc2a27144, 32'h42e49a66},
  {32'h450c803e, 32'h4377cfc2, 32'h425939dc},
  {32'hc496ab3a, 32'h4328d2ab, 32'hc1432194},
  {32'h43cf58d2, 32'hc32f8748, 32'h409c37b4},
  {32'hc3975a82, 32'h43d9b9f8, 32'h42a02fb9},
  {32'h448ba659, 32'h4112f695, 32'h42285d79},
  {32'hc4d36256, 32'hc2003b68, 32'hc3c74981},
  {32'h44e4b330, 32'h42ca1b2a, 32'hc3b33b6a},
  {32'hc46f37fa, 32'hc267d392, 32'h4280144e},
  {32'h44d44654, 32'h42e35dc2, 32'hc272cdfa},
  {32'hc4fb3a18, 32'hc33d7376, 32'hc3b35d26},
  {32'h4448c1ac, 32'h421496ce, 32'hc285a6bb},
  {32'hc4a72e44, 32'h426885df, 32'h429d7674},
  {32'h444ce961, 32'hc3b41b0f, 32'hc3447db5},
  {32'hc480ed0a, 32'hc2e4ff30, 32'h439dcb02},
  {32'h43c8b3d0, 32'h43820877, 32'h43a52e08},
  {32'hc4940bb6, 32'hc3106916, 32'hc39a52e9},
  {32'h429676ba, 32'hc3a4c25c, 32'hc352d121},
  {32'hc4d837b9, 32'hc33d7d38, 32'h4305e486},
  {32'h450401e6, 32'h42edd582, 32'h43a47b6b},
  {32'hc4735460, 32'hc32ec2a9, 32'hc2d7ac80},
  {32'h44e7b710, 32'h434ff8b2, 32'hc35f96d6},
  {32'hc49f8f68, 32'h440644a0, 32'h4398e035},
  {32'h44efb3ed, 32'hc2be94da, 32'hc3a65277},
  {32'hc4c2b23b, 32'h437fd865, 32'hc314e6c2},
  {32'h44c5f0c1, 32'hc3df38e7, 32'hc3ac6b9c},
  {32'hc4a547a3, 32'h436088fb, 32'hc4001975},
  {32'h4516fbf9, 32'h42e12f6f, 32'hc1d2d832},
  {32'hc3b0da3a, 32'hc307c51d, 32'h438c9fa4},
  {32'h44874142, 32'hc3c3121c, 32'hc30f99b6},
  {32'hc4c5f115, 32'h432cfe27, 32'h431d7764},
  {32'h4440ff87, 32'h42fcdb54, 32'h420ee001},
  {32'hc4826e47, 32'h4325c432, 32'h41c3136e},
  {32'h4409bbd8, 32'h43f0b906, 32'h43161979},
  {32'hc50ccd82, 32'h423b7229, 32'hc30de1aa},
  {32'h4452746c, 32'hc2f24030, 32'h442eacf8},
  {32'hc4ff22d0, 32'h423e1a9e, 32'h42bd3213},
  {32'h4506ea0a, 32'hc2f42b83, 32'hc37370a5},
  {32'hc512d1b1, 32'hc36e89a0, 32'hc265be38},
  {32'hc50d9b9e, 32'h43b4b339, 32'h4310071e},
  {32'h4366d558, 32'hc3ae0b8a, 32'h43925514},
  {32'hc3ec1b38, 32'hc0802fb7, 32'hc2a9b083},
  {32'h450a670c, 32'h42893d79, 32'h43c44f8b},
  {32'hc4fe020a, 32'h436d8990, 32'hc29d3a8a},
  {32'h4504d892, 32'h43176d52, 32'hc2142262},
  {32'hc4943df5, 32'hc20a99d7, 32'hc287e404},
  {32'h44eb9c5b, 32'h4223f5e3, 32'h4320d6ea},
  {32'hc4212c5d, 32'hc3079984, 32'h436534e9},
  {32'h440da048, 32'h4297fc49, 32'hc30b8b0d},
  {32'hc4aebacc, 32'h42cf4125, 32'h43358821},
  {32'h44e52871, 32'h4310c363, 32'h43ba5355},
  {32'hc4461726, 32'hc32f02e7, 32'h4321ed39},
  {32'h4453e3fc, 32'hc32aa6a0, 32'hc2f9e152},
  {32'hc3fbfdb2, 32'hc2f3e1fd, 32'h422afce9},
  {32'h44f9b646, 32'hc2bf516d, 32'hc3285296},
  {32'hc40d2fbd, 32'hc2bfb487, 32'hc2d03665},
  {32'h44f930cf, 32'h42270693, 32'h42b10b58},
  {32'hc3a03f55, 32'h43bd8224, 32'h423359aa},
  {32'h449bc700, 32'hc2c7034d, 32'hc384b712},
  {32'hc49ff9d9, 32'h431b6dd1, 32'h42d7dcaa},
  {32'h43d31ed0, 32'hc42d60fb, 32'h4340b71e},
  {32'hc44c475e, 32'hc13f5fde, 32'h432542c5},
  {32'h4408474c, 32'h41ec8944, 32'h44053006},
  {32'hc50baa72, 32'hc395a015, 32'hc2828a26},
  {32'h43bf12e4, 32'h433ebe40, 32'h422bd8a5},
  {32'hc5013273, 32'h43ca2a58, 32'h42cfdde7},
  {32'h449426e2, 32'h43f26252, 32'h4180d3fa},
  {32'hc4ac517d, 32'hc342472e, 32'h42330052},
  {32'h43d36178, 32'h428e8a86, 32'h43a678a1},
  {32'hc44a32c9, 32'h43dd7d77, 32'hc1e96320},
  {32'h450d2f72, 32'hc278c9e3, 32'h424ea055},
  {32'hc4a4af42, 32'h434ef872, 32'h4248bbf7},
  {32'h44af8010, 32'h42ca43d0, 32'hc1806f0b},
  {32'hc4965078, 32'hc393f03e, 32'h43648638},
  {32'h44389974, 32'h4354fe21, 32'h42e1a85d},
  {32'hc4c90f22, 32'hc2ffb0a8, 32'hc1b4ebf1},
  {32'h44b62d3b, 32'hc230990e, 32'h433e5ed9},
  {32'hc501f6a3, 32'hc2bcda7e, 32'h41cee07e},
  {32'h44ba4736, 32'h4201b04f, 32'h441afad7},
  {32'hc4dd04a9, 32'hc350c3df, 32'hc35c46ae},
  {32'h44d90c6e, 32'h435cf938, 32'h424321bc},
  {32'hc49faf31, 32'h4389c47f, 32'h4325855b},
  {32'h4495d13c, 32'hc1299dc4, 32'h4392eeca},
  {32'hc49ae65a, 32'h41d73bff, 32'hc3895fb8},
  {32'h44ec814a, 32'hc3809b8c, 32'h431c4a10},
  {32'hc445a60c, 32'hc35e15ec, 32'h425b12af},
  {32'h4506675d, 32'hc3b1adef, 32'h42310770},
  {32'hc4db2395, 32'hc39c8b1d, 32'hc3f45481},
  {32'h44c6b405, 32'hc2daa62c, 32'hc3a48025},
  {32'hc4e7aeca, 32'hc24efe86, 32'hc33ba352},
  {32'h4437bff8, 32'hc312964c, 32'hc10ad602},
  {32'hc3196e08, 32'hc3748541, 32'h43bf74dc},
  {32'h445734c4, 32'hc23c33e2, 32'h43c57339},
  {32'hc46cb884, 32'hc17030b4, 32'hc2c1b2e0},
  {32'h44a18ef8, 32'h43e75b1a, 32'h430835e0},
  {32'hc4d4d922, 32'hc358e80b, 32'h432f6077},
  {32'h44d14b19, 32'hc3c7bb64, 32'hc3abcfca},
  {32'hc2154830, 32'h4387200d, 32'hc2ecfa14},
  {32'h44bedfe8, 32'h43ab690f, 32'h435981fe},
  {32'h43064b80, 32'hc2eb0df0, 32'hc38d8cd7},
  {32'h43b3b6ae, 32'hc2b23357, 32'hc3057f94},
  {32'hc394612c, 32'hc31017a1, 32'h41a48926},
  {32'h4511a974, 32'hc20f6297, 32'hc3997001},
  {32'h4323f65a, 32'hc2254613, 32'hc2f0d142},
  {32'h44baf9e0, 32'hc2d68f19, 32'h4380b128},
  {32'hc46df7ef, 32'h4182b69e, 32'h433d0d8d},
  {32'h4483a0cb, 32'hc3b88558, 32'hc31b32a1},
  {32'hc44c7dab, 32'h435cc965, 32'h4239d749},
  {32'h445a6ace, 32'h435c1d4d, 32'h4296e0ab},
  {32'hc3be3d50, 32'hc3ca79b3, 32'hc214420f},
  {32'h447c8e52, 32'hc2598dba, 32'hc294a4a7},
  {32'hc4965eee, 32'hc3ab3f5d, 32'h439586db},
  {32'h437483d8, 32'h43078626, 32'h4305990a},
  {32'hc4d6d179, 32'hc1cf573c, 32'h42858dbf},
  {32'h45076c34, 32'hc33b02e6, 32'h42bfc66e},
  {32'hc46a8e82, 32'hc2547804, 32'h42514bec},
  {32'h449a97f8, 32'h43bc7a55, 32'hbe95858d},
  {32'hc4ad3862, 32'h43124f9a, 32'hc3160be8},
  {32'h4505d5d6, 32'h42c5a599, 32'h40be07d2},
  {32'hc40bd244, 32'h43a6e93b, 32'h434faa45},
  {32'h44d4711e, 32'hc044461b, 32'h43f25b00},
  {32'hc4283ee0, 32'hc1030453, 32'h43af03c7},
  {32'h44ad81c4, 32'h41ef0131, 32'hc2b88f89},
  {32'hc4f896a2, 32'hc2e0ad72, 32'h414ddddd},
  {32'h44403896, 32'h4369d8ba, 32'h432295fe},
  {32'hc4deca19, 32'hc3a4970b, 32'hc2e6a780},
  {32'h44522fec, 32'hc44eb701, 32'hc365ba90},
  {32'hc506346c, 32'hc33936d2, 32'h426652f6},
  {32'h4501dfea, 32'hc345dd2f, 32'h42751de6},
  {32'hc4ff26cd, 32'hc379108c, 32'h4283ac9d},
  {32'h44bf40a4, 32'hc3986a0d, 32'hc1bbbac9},
  {32'hc4d9d42f, 32'hc1dd1dcb, 32'hc39242ec},
  {32'h430f8690, 32'h4391686c, 32'hc25f52d8},
  {32'hc3516152, 32'h437419c1, 32'hc351d193},
  {32'h450a6bb1, 32'hc28740ae, 32'hc3d6f564},
  {32'hc4cd8f0a, 32'hc21ff693, 32'h4163c4c8},
  {32'h4400251a, 32'hc22e23bb, 32'hc20a9c6f},
  {32'hc4001a5c, 32'h42be952e, 32'h434dd26d},
  {32'h450ee968, 32'hc13302d0, 32'h4355e0a6},
  {32'hc4e106fa, 32'h440ed368, 32'h4325639e},
  {32'h44d13209, 32'h42f46cc2, 32'h42bb71cc},
  {32'hc5020318, 32'h429345c3, 32'hc37598fd},
  {32'h4419936b, 32'hc331303f, 32'h437b5f81},
  {32'hc4e66499, 32'h42eda1bf, 32'hc248bb53},
  {32'h44afd686, 32'hc34750a3, 32'hc30eda06},
  {32'hc48e5525, 32'hc40ee720, 32'h41ff3331},
  {32'h44da98d6, 32'hc3daefa7, 32'h4378ac9f},
  {32'hc513712c, 32'h432969c5, 32'h42a26102},
  {32'h437ae6b4, 32'hc33c8fb8, 32'h41dc0ad4},
  {32'hc3e9ddd0, 32'hc3598014, 32'h41210ef4},
  {32'h4326ba69, 32'hc31b779e, 32'hc32a276c},
  {32'hc4cab1fe, 32'hc27a8660, 32'hc291d30a},
  {32'h44cdbe9b, 32'h430b5eb9, 32'hc3353f2f},
  {32'hc4e4680b, 32'hc342d736, 32'h43542aad},
  {32'h44b1d9ca, 32'hc3eccd57, 32'h435d5367},
  {32'hc482eedd, 32'hc203e2f1, 32'hc35af03c},
  {32'h450d0882, 32'hc38183bd, 32'h42f178c5},
  {32'hc5198a52, 32'hc1adb776, 32'hc1297790},
  {32'h44b84417, 32'hc34d9c6c, 32'hc1f80a4c},
  {32'hc5042e37, 32'h41752660, 32'h439575c3},
  {32'h41640200, 32'hc2d4b5b0, 32'hc2ebc3d8},
  {32'hc45dd578, 32'hc3def309, 32'h3d314090},
  {32'h450e6c34, 32'h440160fb, 32'hc359aef6},
  {32'hc45088ce, 32'h43c1b304, 32'h42d34e8e},
  {32'h44121054, 32'h4348c2db, 32'hc284e552},
  {32'hc4566e7e, 32'hc302d839, 32'h436f78cf},
  {32'h45048d33, 32'h42d29864, 32'h42cb4ff0},
  {32'h419609e0, 32'hc36a6c8e, 32'h43574b35},
  {32'h44d98ad8, 32'hc3002aba, 32'hc356c93b},
  {32'hc46511dc, 32'h43c3ac86, 32'h438e8f59},
  {32'h44f22fac, 32'h430e0022, 32'hc2853ca0},
  {32'hc4325f4e, 32'hc308554c, 32'h433729b7},
  {32'h449fe02f, 32'hc3ad17a2, 32'hc28416a8},
  {32'hc42c9fe8, 32'hc2c6fae5, 32'h433c9685},
  {32'h452057b5, 32'h44165c4e, 32'h43a5952f},
  {32'hc4670a6c, 32'hc30e3b4c, 32'h43242e85},
  {32'h4441a046, 32'hc28185dc, 32'h436559ff},
  {32'hc4c66b1b, 32'h42e446e4, 32'hc1cb94ca},
  {32'h44c6f53a, 32'hc2d1a480, 32'hc277523b},
  {32'h42ccb452, 32'h43a983d0, 32'hc1e5bdaa},
  {32'h44d7b323, 32'h43daa3e0, 32'h422678ca},
  {32'hc38a9616, 32'hc326b8cf, 32'h431a0302},
  {32'h4513d862, 32'h438d6fd7, 32'hc1b597fb},
  {32'hc40cf41c, 32'hc212e6e9, 32'hc3b22bbc},
  {32'h440e8922, 32'h430738b4, 32'hc2338096},
  {32'hc45b7694, 32'hc12aad12, 32'h4334583e},
  {32'h448064c0, 32'hc108fab3, 32'h43cd0c30},
  {32'hc4effba8, 32'h41188342, 32'h4281ed9b},
  {32'h445de2c6, 32'h42d2f849, 32'hc3d2e91c},
  {32'hc497ad30, 32'h4330d7f6, 32'hc365023f},
  {32'h44ed4e0a, 32'hc3af67af, 32'hc3b66de2},
  {32'hc50d7934, 32'h43dcb34c, 32'hc3a4f8c4},
  {32'h45034f60, 32'h4382c021, 32'hc3dcd8de},
  {32'hc386a06a, 32'h42a66aef, 32'h42c52dec},
  {32'h4450f0e1, 32'hc3890293, 32'h43911995},
  {32'hc3192b82, 32'h42bbeef7, 32'hc391e762},
  {32'h42e4bc24, 32'h43a06e8b, 32'hc30e4eaa},
  {32'h422e25d8, 32'h435305bc, 32'hc32c4fb6},
  {32'h4414ae04, 32'hc12d130c, 32'h41c9b1fe},
  {32'hc465acc6, 32'hc311ade3, 32'h43df2a67},
  {32'h44b2387d, 32'h42c5371c, 32'h43563764},
  {32'hc4e44dcb, 32'h43e8bbdf, 32'h434bd99a},
  {32'h4485cd16, 32'hc23b827c, 32'h431a7df0},
  {32'hc3916908, 32'h43104ec9, 32'h4101cd8c},
  {32'h44855881, 32'hc30c6259, 32'hc24f6b7e},
  {32'hc409985c, 32'h41df6d01, 32'hc0a8c370},
  {32'h44c902f1, 32'hc29fac22, 32'hc3bc418f},
  {32'hc503eaca, 32'hc3840076, 32'h436e3afc},
  {32'h44efdc69, 32'h433857b6, 32'hc30633e0},
  {32'hc4c12b38, 32'h4382b706, 32'hc3c899e2},
  {32'h45117951, 32'h43720ef1, 32'h439d10fb},
  {32'hc489ba16, 32'hc2e1075c, 32'h430a5b99},
  {32'h43e88eb8, 32'h4212f49a, 32'h4306e058},
  {32'hc4fd6526, 32'h437bff00, 32'h42e100fd},
  {32'h4430f5ca, 32'h433611aa, 32'hc32e7ce3},
  {32'hc46e41a9, 32'h43b41fc9, 32'h43b42836},
  {32'h44aec1fe, 32'h43dc1270, 32'hc3a71aaf},
  {32'hc2906f00, 32'hc23ad649, 32'hc3d810d1},
  {32'h44805fcc, 32'h43f0adda, 32'hc14f9158},
  {32'hc4628b48, 32'h43053a78, 32'h4401c6ab},
  {32'h44814d52, 32'hc256fcb7, 32'hc2091965},
  {32'hc519d455, 32'hc36017ab, 32'h43962313},
  {32'h4403fd9a, 32'hc37805b0, 32'hc3988ded},
  {32'hc4947574, 32'h41a49845, 32'h424a7b48},
  {32'h44cf8399, 32'h435976cd, 32'h435ac42f},
  {32'hc4e865b7, 32'h4318d460, 32'hc2fc3565},
  {32'h4358b930, 32'hc0031bb8, 32'h42803299},
  {32'hc4d48808, 32'h43891255, 32'hc26117fa},
  {32'h44113c02, 32'hc3176923, 32'h43c71920},
  {32'hc47f0a98, 32'h4380661b, 32'hc32db1a7},
  {32'h44ab13fa, 32'hc2c07918, 32'hc2bcc579},
  {32'hc443656f, 32'h43a83b5a, 32'hc2203f78},
  {32'h4447ac3a, 32'h43026069, 32'h42688b53},
  {32'hc4c23c96, 32'hc2205a0e, 32'hc2785d69},
  {32'h44a1fd74, 32'h40a1e134, 32'hc3192746},
  {32'hc41a5c32, 32'hc2158413, 32'hc20207d1},
  {32'h448f7c3a, 32'hc3cc26d2, 32'hc24b8020},
  {32'hc314ad30, 32'h428da606, 32'hc2723390},
  {32'h44ca891e, 32'hc32c8ec0, 32'hc2d001c2},
  {32'hc4c1e096, 32'h418c7055, 32'h41fea931},
  {32'hc37ecbc4, 32'h42e6c9a5, 32'hc31317d0},
  {32'hc4f6860e, 32'hc2ac3593, 32'h429df8b8},
  {32'h43d4c648, 32'h434b5ae1, 32'h43699b89},
  {32'hc49298d5, 32'hc1c00811, 32'hc37ab7f4},
  {32'h449c31db, 32'h43061b9a, 32'h433a01aa},
  {32'hc3ae0270, 32'h43922b74, 32'hc367bcd2},
  {32'hc2ce2260, 32'h42f9b273, 32'h433d5825},
  {32'hc39c4b4c, 32'h425e96b8, 32'h428c9fcf},
  {32'h45086479, 32'hc34cc54f, 32'hc3ad6038},
  {32'hc4f0ef1d, 32'h437596ae, 32'hc213e272},
  {32'h44ce1091, 32'hc2f69474, 32'hc29a8bb9},
  {32'hc458e6ab, 32'h424eb4d2, 32'hc211476a},
  {32'h44b8b564, 32'h42dfd5f2, 32'hc284afb8},
  {32'hc4cbb14c, 32'hbfbbbb92, 32'h4314e6a4},
  {32'h447bb49a, 32'h42414e73, 32'hc3aef4a9},
  {32'h43952d96, 32'hc3f86e13, 32'h4270788d},
  {32'h42d6de90, 32'h428907de, 32'hc288a6c4},
  {32'h41198800, 32'h42e81ef9, 32'hc3c755a2},
  {32'h448d3463, 32'h426c226c, 32'h43d372e5},
  {32'hc42908e6, 32'h43c1982f, 32'h43cfcffc},
  {32'h443ecde2, 32'h42a02ed4, 32'h43d9d52e},
  {32'hc4c6344f, 32'hc380e26a, 32'hc2a0bac8},
  {32'h44e68cd6, 32'h438b2db0, 32'h429920b5},
  {32'hc46cafda, 32'hc3535fb4, 32'h40f0292b},
  {32'h4405f871, 32'hc30d834a, 32'hc3abd941},
  {32'hc503f214, 32'h42ac331c, 32'h442413e7},
  {32'h443a152e, 32'h436d86ab, 32'hc22d9c46},
  {32'hc458e193, 32'h431bde3e, 32'hc3717d6a},
  {32'h450fb2f3, 32'h43022768, 32'hc3c64278},
  {32'hc504003b, 32'hc375b3f4, 32'h42c05656},
  {32'h442b0e8a, 32'h43b9a72c, 32'h426755eb},
  {32'hc4839c95, 32'hc3637f9d, 32'hc154944e},
  {32'h4322e6c0, 32'hc305c4d6, 32'h4144b90a},
  {32'hc4f5adf1, 32'h424aaf01, 32'h4286e2a4},
  {32'h44dc8dfd, 32'h4315fbe9, 32'hc32e6e6e},
  {32'hc4b1eaa0, 32'h42c0b1b6, 32'h4347a880},
  {32'hc4372bd2, 32'h43a7ba8b, 32'h432fabd4},
  {32'h44a69d9c, 32'h434aeb6c, 32'hc30208c1},
  {32'hc4c7869a, 32'h43f7d982, 32'hc235dd76},
  {32'h44a76764, 32'h43075e95, 32'h42ee947b},
  {32'hc50edfed, 32'hc31b8580, 32'hc1fc5b44},
  {32'h44712b52, 32'hc2d3b1b0, 32'h43bcb12b},
  {32'h4372e99b, 32'h4249e48d, 32'hc30942f9},
  {32'h44fc8968, 32'h425cbea8, 32'hc2fdcc9a},
  {32'hc5060a4b, 32'hc3941d23, 32'h423c954c},
  {32'h451d516d, 32'h423709a2, 32'hc30d7020},
  {32'hc4d48508, 32'h42356781, 32'hc3a51696},
  {32'h44943956, 32'hc2f6cfba, 32'h4323adc0},
  {32'hc5147ec9, 32'h43710592, 32'hc300a8fb},
  {32'h448bef2f, 32'h434aff9c, 32'hc3b06c4b},
  {32'hc48f5c98, 32'h42fe9a40, 32'hc3803d9c},
  {32'h446c3795, 32'hc0ec5e5d, 32'hc2f8fabb},
  {32'hc4012426, 32'hc21193fa, 32'hc3478369},
  {32'h449d55a5, 32'h436ac2a3, 32'h42b7362d},
  {32'hc4db4fc9, 32'hc2ea1ddc, 32'h431e3fe8},
  {32'h446a6d8b, 32'hc2f01a09, 32'hc2923d2d},
  {32'hc5011ee2, 32'h436e9fe3, 32'hc2380244},
  {32'h44bab936, 32'hc0d0552d, 32'hc32c2cdb},
  {32'hc517a21c, 32'hc28496ee, 32'h43a072a1},
  {32'h450eae38, 32'h421523d5, 32'h43a96a7a},
  {32'hc3afd23e, 32'h43d4b101, 32'h424cf8cb},
  {32'h443a7744, 32'h432a631d, 32'h42d9c882},
  {32'hc48593eb, 32'hc2cde30a, 32'h4349c4ec},
  {32'h4435a114, 32'hc34bdb92, 32'h43783170},
  {32'hc5055b7c, 32'hc126b5b2, 32'h428a30f9},
  {32'h446e4826, 32'hc33d1614, 32'h42775af2},
  {32'hc51ef6d5, 32'h42df82dc, 32'h4351de78},
  {32'h444f2bfc, 32'hc2aace87, 32'hc29b9e95},
  {32'hc44763af, 32'h426fba00, 32'hc3d4c4ec},
  {32'h45011b43, 32'h42abbba2, 32'hc3abc623},
  {32'hc4fc77b0, 32'h43b19ee6, 32'h44017d77},
  {32'h44dc58fe, 32'hc32b090d, 32'h43063d7c},
  {32'hc3b2b1ec, 32'h42385684, 32'h41c415c0},
  {32'h44e8f241, 32'h42a6a274, 32'h431c3a36},
  {32'hc5158862, 32'hc2fdf27b, 32'hc2a1f184},
  {32'h44c78670, 32'h43aef244, 32'h43f71812},
  {32'hc4472eba, 32'h43b26a9d, 32'h4367ef12},
  {32'h4521b536, 32'h43c7e4f6, 32'h432a77e8},
  {32'hc4e51ede, 32'hc3a83b21, 32'hc214745a},
  {32'h44f361b8, 32'hc38b42c3, 32'hc38752d3},
  {32'hc3fefe47, 32'h42b6e91b, 32'hc38ae127},
  {32'h4250f450, 32'h43705887, 32'hc2afd718},
  {32'hc4e178e5, 32'h4378fa9f, 32'hc338f6a1},
  {32'h449d12dc, 32'hc22c4bfc, 32'hc2c005a3},
  {32'hc4001f65, 32'hc26c6330, 32'hc1c67911},
  {32'h44962af3, 32'h434c250f, 32'h434ef0c7},
  {32'hc50d7040, 32'h438f1265, 32'h43e06ea8},
  {32'h45108dcf, 32'hc1a25633, 32'h42defc72},
  {32'hc39ce900, 32'h41b8b3b1, 32'hc301a944},
  {32'h443bbc4c, 32'h41d048b2, 32'h43bfd089},
  {32'hc4d25082, 32'h43c4643c, 32'hc29d0b43},
  {32'h43f8505a, 32'h42fff943, 32'h433fe709},
  {32'hc482184d, 32'h43ef8469, 32'hc3f57545},
  {32'h44a253d8, 32'hc3ddb121, 32'h43138cb1},
  {32'hc485ba68, 32'hc3f1bb1e, 32'h42d9d39d},
  {32'h44381ecc, 32'hc1a903ab, 32'h43176dde},
  {32'hc4ee23cc, 32'hc294d971, 32'hc1045ee2},
  {32'h43d2a746, 32'h43e7e961, 32'h43a75c17},
  {32'hc514dc81, 32'hc3db613e, 32'h430cefb7},
  {32'h447f48db, 32'h432c097b, 32'hc39a0413},
  {32'hc499a35b, 32'hc3be612e, 32'h42a77188},
  {32'h4436cae0, 32'h430fc545, 32'hc1a04f46},
  {32'hc493b83f, 32'hc152b1f4, 32'hc3bbbf8b},
  {32'h43ee571a, 32'h41191e90, 32'h42bfc09f},
  {32'hc4b12672, 32'hc21ca754, 32'h406bbd72},
  {32'h4497ba13, 32'h41fe4d07, 32'hc3942d21},
  {32'hc3339b18, 32'hc31a2a06, 32'hc31e74ca},
  {32'h44b88ca9, 32'hc39788ed, 32'h439c00a7},
  {32'hc40f99b4, 32'hc24a8537, 32'hc064d6e6},
  {32'h44b91634, 32'hc188f6b8, 32'h44222552},
  {32'hc4477cc7, 32'hc35e4064, 32'h431d8f11},
  {32'h450d94c6, 32'h420d860a, 32'hc3a10047},
  {32'hc46cb4b9, 32'h42200b04, 32'hc382cea8},
  {32'h44b4c560, 32'h4175cf3d, 32'h43f0901e},
  {32'hc4c6af29, 32'h41d0a720, 32'hc33e7f2f},
  {32'h451400b6, 32'h429a3f73, 32'h438646f6},
  {32'h4293300c, 32'h431b32d4, 32'h41df09a6},
  {32'h44c08f1c, 32'h4221ebb9, 32'hc3187ea3},
  {32'hc4864058, 32'h42eb3737, 32'hc40d3c26},
  {32'h4418c380, 32'hc3be9ba6, 32'h43388283},
  {32'hc4a32da9, 32'h43c802d4, 32'hc3d80378},
  {32'h44d23129, 32'h4313725f, 32'h42f7572a},
  {32'hc285bfbb, 32'hc12697d7, 32'hc39285aa},
  {32'h443a3dbc, 32'h42730533, 32'h43df4be1},
  {32'hc4da0241, 32'h42e02c94, 32'hc37d1262},
  {32'h443f92ce, 32'h4301261b, 32'h429bb27e},
  {32'hc4c935ab, 32'h43a8c643, 32'h430642d3},
  {32'h44ec1096, 32'hc2814d72, 32'h4373fb11},
  {32'hc43d893f, 32'h42f1a731, 32'h4318923e},
  {32'h44f0be29, 32'hc37921bb, 32'h43195c96},
  {32'hc3b13e30, 32'h42aeb987, 32'hc400f36f},
  {32'h44986b17, 32'hc3348cee, 32'hc22a5f69},
  {32'hc4ef4be4, 32'h42ce0fd6, 32'hc22d39f5},
  {32'h44cff7fa, 32'h42a0a6ac, 32'h4228077e},
  {32'hc4fdb9e7, 32'h42ee96f8, 32'hc1c798fc},
  {32'hc1c1f260, 32'h43afb016, 32'h3f7adcc0},
  {32'hc4317828, 32'h42ad9f19, 32'hc45e224c},
  {32'h44f8d840, 32'hbf06c920, 32'h414516d5},
  {32'hc4df8300, 32'h41d247e8, 32'hc3164fe6},
  {32'hc3f53a10, 32'hc3220ab7, 32'hc3529d85},
  {32'h446f191e, 32'hc36e1a10, 32'hc27b1243},
  {32'hc2b63e30, 32'h43167197, 32'hc2da549d},
  {32'h449938ba, 32'hc3ad45db, 32'h41e8cddc},
  {32'h3f3aa3fe, 32'h43bd3b74, 32'hc1c23d2f},
  {32'h44979450, 32'hc2fc003d, 32'hc3dfff72},
  {32'hc2eb1f64, 32'hc36507a3, 32'hc3393e60},
  {32'h43df1eb4, 32'h430faf4e, 32'h42f69407},
  {32'hc4a85ee1, 32'hc378e256, 32'h425fc186},
  {32'h44513c60, 32'h435a2c0c, 32'hc2420a3d},
  {32'hc4cce840, 32'h42b9229f, 32'hc381e0db},
  {32'h44adf450, 32'hc3860b77, 32'h41e3cf70},
  {32'h439c0394, 32'h43292502, 32'hc3062548},
  {32'h44e252b0, 32'h435f716f, 32'h42d3c6ba},
  {32'hc44a84d1, 32'h43d46440, 32'h436764b1},
  {32'h4267c035, 32'h4405caee, 32'hc3a7fd8d},
  {32'hc5016b05, 32'hc37adf56, 32'h425a8033},
  {32'h43a4f1eb, 32'h43263da3, 32'h431ad229},
  {32'hc483089c, 32'h42906850, 32'hc3905d13},
  {32'h44d5804a, 32'h42f8628c, 32'hc2c79114},
  {32'hc3a25f54, 32'hc20fc8a0, 32'h41345962},
  {32'h43d89b56, 32'hc1746f2c, 32'h433ded58},
  {32'hc4fd3f38, 32'h4356509f, 32'hc32cf955},
  {32'h438ec158, 32'hc2a9af40, 32'h419e0ae0},
  {32'hc4fab717, 32'hc342f029, 32'hc326f636},
  {32'h4505c7ac, 32'h431426f9, 32'hc2b01ec7},
  {32'h432ed5d9, 32'hc3821a9b, 32'hc30af36c},
  {32'h44615b40, 32'hc3ad9285, 32'hc385a2c4},
  {32'hc3265086, 32'hc2d1bf8e, 32'hc32be6c6},
  {32'hc4eb90a6, 32'h3f06db08, 32'hc1f30843},
  {32'h44e1f5de, 32'hc3112b78, 32'h42888c6e},
  {32'hc4feeda4, 32'hc3ebbbbd, 32'hc3d031fe},
  {32'h44d46c3e, 32'h41046f7f, 32'h439aa521},
  {32'hc48ad6e5, 32'hc3913ca9, 32'hc2dcb29e},
  {32'h44a67b28, 32'h4331c45b, 32'hc3857b10},
  {32'hc4a1fbcd, 32'hc384ca55, 32'hc41db921},
  {32'h4446edca, 32'h433fd77f, 32'h42b08c31},
  {32'hc51c84a0, 32'hc274d462, 32'h43084c46},
  {32'h44874644, 32'h42d405fc, 32'hc2f21056},
  {32'hc3bc8f2c, 32'h429a7d8b, 32'h43abf249},
  {32'h445b0b41, 32'hc01fa3a3, 32'h44067471},
  {32'hc411a9a8, 32'hc1ee27b8, 32'hc338bbdf},
  {32'h4341c388, 32'h4323415c, 32'h43d5dbbc},
  {32'hc46cbbac, 32'hc30f1933, 32'hc20d8c97},
  {32'h44ad07c7, 32'h4295ec9b, 32'hc2eebd5b},
  {32'hc4041b58, 32'h4303e9c9, 32'hc3996593},
  {32'h429b57e0, 32'hc30dc2b6, 32'h4297d513},
  {32'hc4ad4d72, 32'h43130cf8, 32'h428613a2},
  {32'h442fb4c8, 32'h42b7ef65, 32'h42900d76},
  {32'hc3e54304, 32'hc2f00880, 32'h4274eb33},
  {32'h44d9a678, 32'hc2489e87, 32'hc30c2a8d},
  {32'hc4f60015, 32'hc2098480, 32'hc31de7f6},
  {32'h44b3396d, 32'h43977933, 32'h42ef6e16},
  {32'hc4e7d140, 32'h429f3ad4, 32'hc2b1c2a7},
  {32'h451dcfb8, 32'h433877a3, 32'hc38765ce},
  {32'hc517b8aa, 32'h4200db67, 32'hc39adb80},
  {32'h4418bcb4, 32'hc3843714, 32'hc31508ac},
  {32'hc50b06d4, 32'hc2a34a93, 32'h420db228},
  {32'h44b0d52c, 32'h43903704, 32'h43633067},
  {32'hc50c2277, 32'h43192c2a, 32'h43636e22},
  {32'h4355b77c, 32'h41c242d8, 32'hc3944815},
  {32'hc50cde84, 32'hc2fe21f3, 32'hc3c4f0d2},
  {32'h44382528, 32'h42724d62, 32'h420c4791},
  {32'hc3f730b8, 32'hc1e45f13, 32'h4331ab3b},
  {32'h42d5dbe4, 32'h423a0352, 32'h43b71edb},
  {32'hc4af10b9, 32'h4312f0ea, 32'hc204d67f},
  {32'h44e99104, 32'hc1cfef98, 32'h437b9c94},
  {32'hc4bcbbe6, 32'hc2838ec6, 32'h4349c03a},
  {32'h449164a8, 32'hc31a3196, 32'hc322c941},
  {32'h42957190, 32'h42f09329, 32'hc11a1926},
  {32'h448ebe41, 32'hc1905bf6, 32'h436e49c8},
  {32'hc4182950, 32'hc32f0bd6, 32'h4396b250},
  {32'h44d31914, 32'hc30ad49d, 32'hc3775c3b},
  {32'hc50123ce, 32'h41ab4fd4, 32'hc387be8f},
  {32'h441ed33a, 32'h42b564fd, 32'hc3546fdb},
  {32'hc4967f87, 32'h43866030, 32'hc3cfbee5},
  {32'h444ca17a, 32'h4203581c, 32'hc3a0c606},
  {32'hc3c34e78, 32'h432b837e, 32'h4225c826},
  {32'h44f57dc7, 32'hc41e6104, 32'h43f027bc},
  {32'hc3abcd98, 32'hc40af3e9, 32'h42584747},
  {32'h43972784, 32'hc39befc6, 32'h432192b9},
  {32'h44f7742c, 32'h4101b31d, 32'h4405a04f},
  {32'hc3bcfcc8, 32'h4403be52, 32'h42f70310},
  {32'h43c9d844, 32'h41cf1810, 32'h43052085},
  {32'hc5082aa2, 32'hc2a8a4f5, 32'hc3507137},
  {32'h42058c60, 32'hc320fa15, 32'hc4074af8},
  {32'hc2993ae2, 32'h4363ccd1, 32'h42d7b7cd},
  {32'h441c6fb9, 32'hc2c41ec8, 32'hc1762180},
  {32'h42f7f480, 32'hc39f7b81, 32'h41abf7cb},
  {32'h44703432, 32'h424ea099, 32'h41a05452},
  {32'hc505f79a, 32'hc282ea03, 32'hc3db7cce},
  {32'hc2c465d4, 32'h43cd4b15, 32'h42175ce2},
  {32'hc444d89c, 32'h426d28dc, 32'h41e70921},
  {32'h44ec9a5f, 32'hc3b2aac4, 32'hc31293d3},
  {32'hc44cec44, 32'hc13dbae6, 32'h43d16b35},
  {32'h445d7712, 32'hc3849964, 32'hc392eecc},
  {32'hc508e3fd, 32'hc3ba39c0, 32'hc37dd7ed},
  {32'h44eb24ea, 32'hc12d00ec, 32'h43cb0638},
  {32'hc4aab99a, 32'h42314287, 32'h4349912f},
  {32'h44ec2da8, 32'h43cc6fdb, 32'h426defa4},
  {32'hc3221090, 32'h42969125, 32'hc3d507dc},
  {32'h4501820f, 32'h42becee0, 32'h43aa46cc},
  {32'hc3ff7ebe, 32'h431c885e, 32'h424317bf},
  {32'hc10e4b10, 32'hc33c473c, 32'h41dcf38b},
  {32'hc4ff0fd3, 32'hc3096f2a, 32'hc3687591},
  {32'h448c2284, 32'hc3a78e46, 32'h41a25350},
  {32'hc4c2f8aa, 32'h431ed5dd, 32'h43945fd1},
  {32'h451bc39c, 32'hc301b4e3, 32'h43930f28},
  {32'hc4e61b56, 32'hbff24948, 32'hc28a8522},
  {32'h4526efb1, 32'hc201e71d, 32'h440b2a1e},
  {32'hc487848f, 32'hc33ca613, 32'hc2de834e},
  {32'h44cbe43d, 32'h43ce67eb, 32'hc2d2017a},
  {32'hc4e7b386, 32'h43bdab6d, 32'h43c9b2b4},
  {32'h43b6eaa8, 32'hc2b06593, 32'h42f3d332},
  {32'hc4abc8ce, 32'h42973e35, 32'hc1faa6e1},
  {32'h44d7a9fa, 32'h428dae30, 32'h4340750f},
  {32'hc4765ff8, 32'hc39be645, 32'h43a62e0f},
  {32'h42deedc0, 32'h438f1591, 32'h43948c0d},
  {32'hc3a09702, 32'hc34bc2b7, 32'hc374ef03},
  {32'h44a153aa, 32'h43c61053, 32'h43f09cf3},
  {32'hc4b6a18c, 32'hc37b8fd2, 32'h43b62ad8},
  {32'h44e20675, 32'hc1b576f8, 32'h430bf5dd},
  {32'hc4984ed6, 32'hc213e87d, 32'hc2288015},
  {32'h44422ea4, 32'h427ae335, 32'h43d2bf8c},
  {32'hc50d2e98, 32'hc00d6e69, 32'h43a301dc},
  {32'h43220bf0, 32'hc3221462, 32'h4404c4a8},
  {32'hc4697a50, 32'h4392c02f, 32'hc30cda19},
  {32'h43e5efc9, 32'h43651f79, 32'hc2915c7b},
  {32'hc4b6cafc, 32'h42ed1bb2, 32'hc3271a35},
  {32'h44964ea1, 32'hc2badba9, 32'hc332a889},
  {32'hc4d69cdb, 32'h42b1a247, 32'hc2b1ed4f},
  {32'h445de0a0, 32'hc24938e8, 32'hc356d124},
  {32'hc4db5dbb, 32'hc333699d, 32'hc2ef1937},
  {32'h43fc3ec8, 32'h4238b16e, 32'h4181c261},
  {32'hc4778a87, 32'h4098fcfb, 32'hc3844cb1},
  {32'h44ebbb40, 32'h42af19ad, 32'h3f4a08b0},
  {32'hc449d740, 32'h4359975a, 32'hc363b4aa},
  {32'h44f8757a, 32'h433ff428, 32'hc405fc47},
  {32'hc4da8b90, 32'hc3594b11, 32'h42faa579},
  {32'h44ce8455, 32'hc35196d8, 32'hc31c3fde},
  {32'hc4e19f10, 32'h43b06eb0, 32'h43787417},
  {32'h44975f56, 32'hc38f44ed, 32'hc30c1138},
  {32'hc439e388, 32'h417de134, 32'h43a91f9c},
  {32'h4297d2c8, 32'hc135ac13, 32'hc3c386ff},
  {32'h44109ddf, 32'hc25102b1, 32'hc284dd6c},
  {32'h448053de, 32'h42e4a269, 32'hc276d5ec},
  {32'hc4c989a6, 32'h43f03c98, 32'hc2be07a4},
  {32'h4323e090, 32'h41a8d546, 32'h43e33bfc},
  {32'hc508d4e3, 32'h42d96c98, 32'h436d7482},
  {32'h44aa2d4d, 32'h42b592f0, 32'hc2ad2760},
  {32'hc502b73f, 32'h429b99cb, 32'hc30752a7},
  {32'h448da915, 32'h43907d03, 32'h439a0253},
  {32'hc445ce96, 32'h42492ec3, 32'hc30075a2},
  {32'h43f7dd4e, 32'h42a242a0, 32'hc32da935},
  {32'hc3c335b4, 32'hc32db877, 32'h440a2b62},
  {32'h43e55448, 32'h42eac062, 32'hc3437b81},
  {32'hc3e4189a, 32'hc26f46eb, 32'hc2fbb090},
  {32'h4398b13c, 32'h429c5625, 32'hc354d907},
  {32'hc3c14594, 32'hc13a50cc, 32'hc2adbf3c},
  {32'h44a3e9ee, 32'h43ea18ce, 32'h3ff1e91b},
  {32'hc5037bba, 32'hc1af0d57, 32'hc38019ae},
  {32'h4431f8b8, 32'h437e9b78, 32'hc37ce9fb},
  {32'hc501e288, 32'hc22dbd2a, 32'h430a3abb},
  {32'h44dc5a00, 32'hc3102f04, 32'h43bbf8bf},
  {32'hc4cd296b, 32'hc17ac8be, 32'hc3a321ae},
  {32'h44d60eb0, 32'hc22beb85, 32'hc2df21a6},
  {32'hc4202008, 32'hc3b7d395, 32'h42dc29fd},
  {32'h44b22073, 32'hc3b861c1, 32'h4386ecd9},
  {32'hc3e2e42c, 32'h43833033, 32'h413372dc},
  {32'h4432a9f7, 32'hc3a0db1d, 32'hc1b4e32e},
  {32'hc3ead0fd, 32'h42d92fdd, 32'h42c461a4},
  {32'h449b97b0, 32'hc36915c3, 32'hc3b51c86},
  {32'hc4ba76b4, 32'hc31dc754, 32'hc2d1799b},
  {32'h444c0d9e, 32'hc385e655, 32'h438286c3},
  {32'hc4a9960a, 32'h439f1b01, 32'hc2ba07a7},
  {32'h45059a49, 32'h3ca51640, 32'hc2b61036},
  {32'hc36e40fb, 32'hc3aaa9f4, 32'h4298117d},
  {32'h447781d4, 32'hc2d78070, 32'h43e981fc},
  {32'hc49d62cd, 32'hc1bcbf5f, 32'hc25eccf4},
  {32'h43e5e1db, 32'h4341bd06, 32'hc2d860d0},
  {32'hc43400a6, 32'hc3aac880, 32'h430a11b0},
  {32'h44c2a134, 32'h4338413c, 32'h42eedbc1},
  {32'hc4531cea, 32'h43201096, 32'hc23b7ad0},
  {32'h44bfed3e, 32'h43becc0f, 32'h43c4d812},
  {32'h43f132da, 32'hc2b6254d, 32'hc2d3d6ed},
  {32'h44399c1c, 32'hc393a871, 32'h4260b1ad},
  {32'hc4ecaba8, 32'h434a2f8a, 32'hc274673e},
  {32'h44deacc2, 32'h42df3d03, 32'hc34d4d37},
  {32'hc3734455, 32'h43a02501, 32'h42d8064c},
  {32'h44f23e6f, 32'hc379c32b, 32'hc297bec9},
  {32'hc49a4a40, 32'hc2b9e8f3, 32'h435e4b99},
  {32'h451431dc, 32'hc34f16a6, 32'h431296e5},
  {32'hc4cf0503, 32'h43920872, 32'h42af7161},
  {32'h42b72a5f, 32'hc39afff4, 32'hc2f8002b},
  {32'hc4e84c44, 32'hc3d94251, 32'h4356b762},
  {32'h4461bc6e, 32'hc1891914, 32'h432af6e3},
  {32'hc4bc4075, 32'h42c9fbda, 32'hc2d030d4},
  {32'h44e3d726, 32'h439cfb41, 32'hc33d3cf6},
  {32'hc50e2bc8, 32'hc3a03783, 32'h42b6be33},
  {32'h438e7c51, 32'h432811be, 32'h437842f5},
  {32'hc317bd80, 32'hc27f73f0, 32'hc41965b4},
  {32'hc3b29f84, 32'hc2680fc8, 32'h42db1427},
  {32'hc4171fc6, 32'hc205b302, 32'h43f57878},
  {32'h447f01f5, 32'hc3e91e6d, 32'hc38ff478},
  {32'hc49ec4a2, 32'hc32a6d86, 32'h439876a0},
  {32'h45046101, 32'h43883e8b, 32'h42c63f3c},
  {32'hc500656c, 32'hc219d538, 32'hc37845ca},
  {32'h44b89ad2, 32'h4198708d, 32'h41b43653},
  {32'hc38e097c, 32'h43a9db74, 32'hc0d17592},
  {32'h422dcbe0, 32'hc3a0ca40, 32'hc3ce5b14},
  {32'hc327fb20, 32'h431eb3be, 32'h43a26851},
  {32'h4414ef9e, 32'hc415d3d3, 32'hc206650d},
  {32'hc5108e57, 32'hc18fe3c3, 32'h43894e80},
  {32'h44d9e271, 32'hc302b4b1, 32'h4103597f},
  {32'hc3e99378, 32'hc301fb08, 32'hc2ecd1c0},
  {32'h44a2f771, 32'hc39daab1, 32'h411c3a26},
  {32'hc3bbfb30, 32'hc25d103d, 32'h43fd374f},
  {32'h446eaa32, 32'h43a72c81, 32'hc3802bf2},
  {32'hc50cc038, 32'hc328feaa, 32'h419505c0},
  {32'h446b4e40, 32'hc39eaea8, 32'hc3a81700},
  {32'hc441010c, 32'h43e720c0, 32'h42ec76fe},
  {32'h43c672f2, 32'h429c6ff5, 32'h434649c1},
  {32'hc4da4683, 32'hc2e81f16, 32'hc11dde1e},
  {32'h450e62ce, 32'h43e13978, 32'hc3cf7e2e},
  {32'hc456ef56, 32'h4416c941, 32'hc2bad397},
  {32'h44a99446, 32'hc27b415b, 32'hc2e1d023},
  {32'hc4dcc47e, 32'hc3dc5fe8, 32'hc2aa8fb4},
  {32'h448cde89, 32'h43a83d89, 32'hc31aaa25},
  {32'hc48f5022, 32'h431ef9e4, 32'h42ad96b3},
  {32'h44b03e7c, 32'hc2a28008, 32'hc397d24c},
  {32'hc413aa18, 32'hc3478ce5, 32'hc31097de},
  {32'h4506f01e, 32'hc3ba472e, 32'h43966b10},
  {32'hc46481f4, 32'h436f3d13, 32'h438bb7d0},
  {32'h44fff561, 32'h424dba45, 32'hc383e6b9},
  {32'hc35066e1, 32'hc37c572f, 32'h4302afc5},
  {32'h44ddd5a1, 32'h42d679d1, 32'h431dff43},
  {32'hc3d07000, 32'hc3c509fe, 32'hc3abc508},
  {32'h44fc4548, 32'h42ec57f3, 32'h43633bdb},
  {32'hc49af456, 32'h42cb72a3, 32'hc32854a7},
  {32'h44838b26, 32'h4326e7bf, 32'hc39e12ca},
  {32'hc508e760, 32'hc29e17a4, 32'hc3a4ad07},
  {32'h45078b60, 32'hc3607ee5, 32'hc36d67dd},
  {32'hc4ce850e, 32'hc33f251c, 32'h43acce44},
  {32'h450adeee, 32'hc3477594, 32'h43d161e5},
  {32'hc4ae8212, 32'hc284428c, 32'hbf73c5b6},
  {32'h44c43bd3, 32'h40ec6789, 32'h43367880},
  {32'hc48121a0, 32'h4351cafb, 32'hc30e25ea},
  {32'h449251f3, 32'hc3b63f06, 32'hc38b1fdd},
  {32'hc4983256, 32'h433a053f, 32'hc19f78c8},
  {32'h43821fa0, 32'h43397952, 32'h4391a4f5},
  {32'hc51156e7, 32'hc0bde37d, 32'h438fd39e},
  {32'h451618ea, 32'h42580cfa, 32'h43c292ed},
  {32'hc4ec8015, 32'h42abc230, 32'hc35e9cd5},
  {32'h44ab0144, 32'hc2ff7ad1, 32'hc2b115b9},
  {32'hc450e0a6, 32'h4344ef0d, 32'h432ddf28},
  {32'h4407e968, 32'hc2553b96, 32'hc36f57fe},
  {32'hc45d1d72, 32'h43024fb0, 32'hc32df0e8},
  {32'h45148fdb, 32'hc343eb0d, 32'h429ad902},
  {32'hc4187004, 32'h434ba6e8, 32'hc283dfdc},
  {32'h44c5bfa5, 32'h427955af, 32'h43135258},
  {32'hc4baed47, 32'h430cd0c3, 32'hc32168fc},
  {32'h44dd3621, 32'h43f25d97, 32'hc310d0f1},
  {32'hc4d8c9be, 32'hc3f06356, 32'hc1cca82b},
  {32'h4421e110, 32'h4121f80c, 32'h41abecf0},
  {32'hc4cdfd28, 32'hc2c67564, 32'hc406fa47},
  {32'h435a9380, 32'hc39fed0c, 32'hc2e9b4a3},
  {32'h43adce90, 32'h43684bd6, 32'h4391e38a},
  {32'h44fc1e3d, 32'hc31382e9, 32'h416de6b5},
  {32'h41f8f780, 32'h438a2f2b, 32'h424faf06},
  {32'h44733503, 32'hc3eb5ae9, 32'hc31ebcbf},
  {32'hc4b14dc9, 32'hc382acd4, 32'h41c3570e},
  {32'h43cd1d88, 32'hc2d022b4, 32'hc223dc8a},
  {32'hc2809640, 32'hc333059d, 32'h4235e3fa},
  {32'h4475d8c8, 32'hc35e1a3e, 32'h431d7e80},
  {32'hc4e1db70, 32'hc34681dc, 32'h439ed0c8},
  {32'h43828240, 32'hc29c9d4b, 32'h3fbe42a0},
  {32'hc4e34efc, 32'hc39af10c, 32'h42911c4f},
  {32'h438852f0, 32'hc2499b5d, 32'h43d8f1e4},
  {32'hc3717816, 32'hc1451675, 32'hc387b01d},
  {32'h4415269c, 32'h4399462b, 32'h43288555},
  {32'hc4aeee12, 32'h42545fde, 32'h43121797},
  {32'h445b018d, 32'h40cfef7f, 32'h42f7bf21},
  {32'hc34ca5be, 32'h43e1442b, 32'h42f376db},
  {32'h4504b5c1, 32'h41e69770, 32'hc29b4dfd},
  {32'hc3fe73ba, 32'h41509351, 32'h43c7390d},
  {32'h44eb5f01, 32'hc339ce28, 32'h4305e731},
  {32'hc44de43e, 32'hc242d9f4, 32'h435a2be1},
  {32'h444c6162, 32'h439eec3e, 32'h4225dd65},
  {32'hc50df4d6, 32'hc30a0113, 32'hc2f750c5},
  {32'h4439e34c, 32'h43b2970b, 32'h434eb711},
  {32'hc409f1b6, 32'h4035f30a, 32'hc2f36216},
  {32'h44b64750, 32'hc0defd26, 32'hc35d09b6},
  {32'hc4f7a046, 32'hc39957b8, 32'h4172e116},
  {32'h45220f0e, 32'hc36dd795, 32'hc2952c44},
  {32'hc3d8a49c, 32'h41d491e4, 32'h4303758c},
  {32'h43f85e13, 32'hc30f1121, 32'hc28c3dce},
  {32'hc43ed594, 32'h43a1ae24, 32'h439a1e47},
  {32'h4425710a, 32'h4259f1f0, 32'hc1d63dd5},
  {32'hc4be3fc8, 32'hc29889ba, 32'hc2adb30b},
  {32'h44145d08, 32'h41de0e53, 32'hc3ba8158},
  {32'hc510e6a0, 32'h42555015, 32'h43586d7a},
  {32'h4511af2c, 32'h43047387, 32'hc3166b77},
  {32'hc52c56ed, 32'h422406fe, 32'hc3962051},
  {32'h44ead53c, 32'hc39aa7b7, 32'h439098a3},
  {32'hc4b85589, 32'hc192df52, 32'hc308ad6f},
  {32'h44b2f491, 32'hc4027dae, 32'h42c5f3c7},
  {32'hc5019f1b, 32'hc237f2bc, 32'hc2b1a633},
  {32'h44177f50, 32'h42b7ed3f, 32'h42bb8e84},
  {32'hc5055d21, 32'h434eaa32, 32'h414c06d6},
  {32'hc4d22b0f, 32'h4123e35c, 32'hc389a9a4},
  {32'h4426499e, 32'h43cb48e2, 32'h4389761c},
  {32'hc4fc3a7e, 32'hc2751be0, 32'hc3db0b4c},
  {32'hc2b8c368, 32'hc3c3423f, 32'hc40f1b71},
  {32'hc4fc732b, 32'h416c9f7c, 32'hc3484bc4},
  {32'h44bf9058, 32'h422b29ba, 32'h437569e2},
  {32'hc4af27d0, 32'h432028b6, 32'hc2c7a6c2},
  {32'h42807018, 32'h4313a288, 32'hc20705c0},
  {32'hc4c049bd, 32'h427390b5, 32'hc38a6348},
  {32'h4446a993, 32'hc3bcde0b, 32'hc36840a9},
  {32'hc2048d94, 32'h40f18f84, 32'hc344bc42},
  {32'h44b04c2e, 32'hc318e92a, 32'h4319f26c},
  {32'hc4f5b7d7, 32'h426dc0bf, 32'h43d3fc92},
  {32'h44a4b4d9, 32'h43bf2519, 32'hc3442de2},
  {32'hc4040273, 32'h4233e475, 32'h41ebd88d},
  {32'h4504f6dd, 32'hc2f53451, 32'h434f4d90},
  {32'hc375b040, 32'h43260a45, 32'h434c80e6},
  {32'h44a141ec, 32'hc2840b7f, 32'hc2d20d8b},
  {32'hc1d4a038, 32'hc2a005d9, 32'h419db2f3},
  {32'h448ad2e5, 32'hc14404c0, 32'h438cbcac},
  {32'hc50f691e, 32'h42c70da3, 32'h42b550c8},
  {32'hc4c8b652, 32'hc3580585, 32'hc349b2f6},
  {32'h446aaa2c, 32'hc2f96ecc, 32'hc26b12da},
  {32'hc5008145, 32'hc2ad3e71, 32'hc3360968},
  {32'h42bac660, 32'h433bb591, 32'h426b6c67},
  {32'hc5052166, 32'hc37fc098, 32'h433f86d1},
  {32'hc1209700, 32'h4285c770, 32'h43280e31},
  {32'hc42a27df, 32'hc3026a2a, 32'hc39e3d8d},
  {32'h450a5974, 32'hc39d4a61, 32'h43c9fac7},
  {32'hc50ac51b, 32'hc20d9e98, 32'hc282d87e},
  {32'h45011ece, 32'h434f65cd, 32'h4313f573},
  {32'hc4fb1a0f, 32'hc27b9175, 32'hc393d6f4},
  {32'h44c03db2, 32'h42ee5414, 32'h41a10c93},
  {32'hc4dc2bd5, 32'hc260a404, 32'h40493adc},
  {32'h4386d406, 32'hc318e2aa, 32'h4352c489},
  {32'hc453928a, 32'h42d3e681, 32'hc36a04c9},
  {32'h43bc91c4, 32'h4215d48b, 32'h439a2e2f},
  {32'hc4832e39, 32'hc3a795db, 32'h432c9947},
  {32'h44b5545a, 32'h4201af98, 32'h42a5289d},
  {32'hc3c52342, 32'h441afb72, 32'hc353b1a8},
  {32'h43f6d575, 32'hc3409b0b, 32'h4384ac3b},
  {32'hc50a8c19, 32'hc3872e15, 32'hc30133b2},
  {32'h43e54164, 32'hc31b4aa3, 32'h423215c1},
  {32'hc30976d0, 32'h435eba15, 32'hc21ef48d},
  {32'h43f5b40d, 32'hc3cd3f92, 32'hc2eac868},
  {32'hc3ab5940, 32'hc36daf5b, 32'h439a6f09},
  {32'h448dce02, 32'hc3996580, 32'hc0676e06},
  {32'hc492ca85, 32'h429a2997, 32'h426e8b16},
  {32'h44e0dd54, 32'h4388eb87, 32'h41fc66f8},
  {32'hc452f3dc, 32'hc2de97ea, 32'h4344c142},
  {32'h449127ca, 32'h4350e4a2, 32'hc1c18170},
  {32'hc4d82748, 32'hc37d82a4, 32'h43812dc4},
  {32'h44b84aba, 32'hc10e1c52, 32'h42f91825},
  {32'hc50364bb, 32'hc3003f90, 32'hc32f1965},
  {32'h449b1d30, 32'h4349070e, 32'hc1345241},
  {32'hc3cfef70, 32'hc1e59924, 32'h421aff94},
  {32'h44d352fa, 32'h42362ee4, 32'hc2d8dcdc},
  {32'hc3636e58, 32'hc28ce55f, 32'h42c31133},
  {32'h44c24e3e, 32'hc27bad99, 32'hc3528c1c},
  {32'hc35ddaf0, 32'h437099d8, 32'hc340201c},
  {32'h435b03b0, 32'hc3aab296, 32'h4309ac27},
  {32'hc498539c, 32'h4326f8ea, 32'hc2b41666},
  {32'h450a175c, 32'hc24399d8, 32'hc3188052},
  {32'hc3135c8e, 32'hc31b7b96, 32'hc3c9d9bc},
  {32'h442fdf0e, 32'h430ea22e, 32'hc3237cb2},
  {32'hc451fd7c, 32'h439626c7, 32'h43302a0c},
  {32'h448a3870, 32'hc1e5d271, 32'hc3a809fa},
  {32'hc46ff2fa, 32'hc30447bc, 32'hc33e22c0},
  {32'h44ec4334, 32'hc2b02f1c, 32'hc2ff261e},
  {32'hc373756c, 32'hc1b59243, 32'h42848c3e},
  {32'h448aad3e, 32'hc21bcaf2, 32'h428f9cf6},
  {32'hc453fdb4, 32'hc1209eb8, 32'h42b1a53a},
  {32'h45064086, 32'hc2f411d0, 32'hc2357444},
  {32'hc4d3a04c, 32'h435346bd, 32'hc3e38e8d},
  {32'h44723352, 32'hc2b163f8, 32'hc3967c1c},
  {32'hc4ed75d8, 32'hc36b9bac, 32'h42d67934},
  {32'h44f1e817, 32'h42fd8ed7, 32'hc1df2942},
  {32'hc48a088e, 32'h41ec236c, 32'hc3208fb9},
  {32'h44d15ed6, 32'hc32b1607, 32'hc238aa66},
  {32'hc458d3b0, 32'h4315fcab, 32'h4422ec40},
  {32'h44f5b00a, 32'hc3d2cc87, 32'h436e38f9},
  {32'hc48eb879, 32'h439d10ca, 32'h42d1e9b7},
  {32'h44a7660a, 32'h432f5e34, 32'hc396d44b},
  {32'hc4b91dc2, 32'hc31894be, 32'h43ae3800},
  {32'h44a9b460, 32'h4343e313, 32'hc28f7cdf},
  {32'hc48f5086, 32'h438101c9, 32'hc2fb0dac},
  {32'h442005df, 32'h4188e341, 32'hc3d9114d},
  {32'hc306c3a4, 32'h4257a1ca, 32'hc190e0a3},
  {32'h4443e81e, 32'h42dcbd35, 32'hc28fbade},
  {32'hc414171e, 32'hc339e9ee, 32'hc1713ae7},
  {32'h44ecf293, 32'hc3a6670c, 32'hc2804b48},
  {32'hc416585f, 32'h40f8368b, 32'h429e7932},
  {32'h44cffd35, 32'hc2deb29e, 32'hc1979d9a},
  {32'hc4b7ea51, 32'h424637c1, 32'h43c5f08d},
  {32'h450ecc28, 32'hc38d71d8, 32'h42264bd3},
  {32'hc3cbd5c0, 32'h430fa547, 32'hc2a5be5f},
  {32'h438c7f9a, 32'h41cad298, 32'hc25aa467},
  {32'hc4514892, 32'h43db4444, 32'h43f8c8b9},
  {32'h44454790, 32'h428b2fe0, 32'h42256122},
  {32'hc4f78371, 32'hc1c5853f, 32'hc36543c9},
  {32'h44e5c983, 32'hc2fa552e, 32'hc3127fea},
  {32'hc5084dad, 32'hc3727019, 32'h429c453e},
  {32'h4331fc10, 32'hc32fe0f0, 32'hc32027a8},
  {32'hc2262080, 32'h418bcd3c, 32'h42c225ac},
  {32'h44d21cef, 32'hc12ae2dc, 32'hc2c7726a},
  {32'hc311aec0, 32'h4228b8b9, 32'h4291f4e2},
  {32'h44743281, 32'h42126bd3, 32'hc2dc15f0},
  {32'hc4e8e2e1, 32'h41e775d4, 32'hc3298b2d},
  {32'h4496a15b, 32'h438765cf, 32'hc2c0df20},
  {32'hc491436b, 32'h415d9b74, 32'h43df4ae8},
  {32'h4486251d, 32'h43371cdf, 32'hc2e9f57b},
  {32'hc46276ca, 32'hc20d0474, 32'hc39b742a},
  {32'h44c7da73, 32'hc1822f7b, 32'hc311d0d4},
  {32'hc4a09668, 32'h42518dc6, 32'h436be99a},
  {32'h43e2a93c, 32'h423d0f19, 32'hc3fc3298},
  {32'hc4e70502, 32'h4352359b, 32'h42ec8b7a},
  {32'h43acbbd9, 32'h434b42c7, 32'hc2d955d1},
  {32'hc4c684e4, 32'h42b6719d, 32'hc31e82a8},
  {32'h44e6dd62, 32'hc405bbd4, 32'h42ab0e33},
  {32'h448051d4, 32'hc31314a7, 32'h42672622},
  {32'hc3bb00b8, 32'h43114691, 32'h43b0ad3e},
  {32'h44be2d11, 32'h42416f7a, 32'h4352e7a0},
  {32'hc2030c80, 32'hc35253f2, 32'h43047b51},
  {32'h451888bf, 32'hc30077d8, 32'hc284d1e8},
  {32'hc453fac2, 32'h42d31ffb, 32'h42b90580},
  {32'h441f26c8, 32'hc00508e0, 32'hc33f0d71},
  {32'hc4835d18, 32'h433e1470, 32'h43dd7bf3},
  {32'h44a8c2b5, 32'hc29fac02, 32'hc19691e6},
  {32'hc4bac906, 32'h42d42ef6, 32'hc1549ac6},
  {32'hc309afbe, 32'h43435e9e, 32'h42cb9aa4},
  {32'hc51e7828, 32'hc2874cc2, 32'h43fae6f4},
  {32'h44a8bfe2, 32'h42c67b11, 32'hc36a35ce},
  {32'hc4a08c52, 32'hc05d4cf8, 32'hc312cefb},
  {32'h444f23d4, 32'h431f631a, 32'hc2b5793c},
  {32'hc467e546, 32'h44064135, 32'hc0b12989},
  {32'h44bd66cc, 32'hc34f5d6a, 32'h42c0e18b},
  {32'hc4a1a2bb, 32'h4318ae2d, 32'hc30c1933},
  {32'h43f8f200, 32'hc332d3fa, 32'h4046867e},
  {32'hc4d2565b, 32'h42fcdfb5, 32'hbfc2ac2c},
  {32'h44f8be6e, 32'hc1f29031, 32'h438aa9b6},
  {32'hc5098219, 32'hc186f81f, 32'hc2b9e5e1},
  {32'h44c2b819, 32'h431bf4fc, 32'hc41a5049},
  {32'hc402e8a0, 32'h418c0cf4, 32'hc2caeca4},
  {32'h44aacd27, 32'h42984c63, 32'hc2e29774},
  {32'hc4fe2350, 32'h43e6d528, 32'h429cd946},
  {32'h44c22ec5, 32'hc2e5fc2c, 32'hc3b3b2aa},
  {32'hc4be61de, 32'hc3c4cc83, 32'h43636a5c},
  {32'h438d5537, 32'h43422032, 32'hc3c3cd41},
  {32'hc411f41a, 32'hc3164563, 32'hc35ef3b1},
  {32'hc3598d08, 32'hc37f5fb0, 32'hc21428ba},
  {32'hc4eb4dfb, 32'hc3fdb5ae, 32'hc3aa6778},
  {32'h4514fc31, 32'h42a288d5, 32'hc329be3e},
  {32'hc46c0816, 32'h42c26ae8, 32'h42c9f358},
  {32'h45098fe1, 32'h43963636, 32'h42ee7c23},
  {32'hc4fc8f02, 32'hc241b2bc, 32'h433703d7},
  {32'h44f6a955, 32'h43ac67ac, 32'hc1c2967c},
  {32'hc48718a7, 32'hc2a3048a, 32'hc3367941},
  {32'h4410fe72, 32'hc31faec2, 32'h4229dacc},
  {32'hc41e02d4, 32'h43453e19, 32'h426338bd},
  {32'h4483f372, 32'h42fb7845, 32'hc311eb54},
  {32'hc48ddab0, 32'h42f59887, 32'hc3439b4e},
  {32'h44def972, 32'h43b51f8d, 32'hc30ad70f},
  {32'hc51c4d9a, 32'hc330c438, 32'hc1b44740},
  {32'h45194d75, 32'hc282094d, 32'hc1e0643e},
  {32'hc45e1294, 32'h43aa61a9, 32'hc38c7eb7},
  {32'h43cde110, 32'h43833620, 32'h409885ba},
  {32'hc513246e, 32'h43508432, 32'h437e9b44},
  {32'hc4da8cc4, 32'hc3178e8a, 32'h41efa805},
  {32'h45094b69, 32'hc38c3274, 32'hc3cdcc0f},
  {32'hc4e68def, 32'h43eb8a83, 32'hc2914a4a},
  {32'h4510eb4b, 32'h4427dece, 32'hc2ee568c},
  {32'hc5145d71, 32'hc25f8454, 32'h42f5ac6c},
  {32'h444448b5, 32'hc2044ee5, 32'hc2cbf2aa},
  {32'hc4a312e2, 32'hc3777864, 32'hc33703d2},
  {32'h43b5fdc8, 32'h42ff486a, 32'h43cf2402},
  {32'h44852343, 32'h436ed35e, 32'hc3dafdce},
  {32'hc45da0ce, 32'h4333c18c, 32'h43c3017f},
  {32'h44c241b0, 32'hc413e0ba, 32'h4317d06a},
  {32'hc389c514, 32'hc384041f, 32'hc3608eef},
  {32'h431fccbc, 32'h4378249a, 32'h43ef89c8},
  {32'h44ce2af8, 32'h441923f3, 32'h41f8e4b3},
  {32'hc42d842a, 32'h41ac433d, 32'h43773adf},
  {32'h45088a12, 32'hc39b3f91, 32'hc342b0bb},
  {32'hc4a50b4b, 32'h42a9613a, 32'hc3732304},
  {32'h4367c572, 32'h43b7572a, 32'hc2868130},
  {32'hc410f714, 32'hc35f0219, 32'hc366ffd6},
  {32'h44b8e147, 32'hc2a40930, 32'h437b2d31},
  {32'hc3545784, 32'hc37cc27b, 32'hc13e7f7b},
  {32'h43852d40, 32'h435af422, 32'hc28d9bd8},
  {32'hc3b77171, 32'h429e051b, 32'h43625fc7},
  {32'h44495769, 32'h4407db06, 32'h43554664},
  {32'hc4be0ea2, 32'h43c2bdd6, 32'h434dfc22},
  {32'h4479466e, 32'h434633ab, 32'hc28d6713},
  {32'hc4bc915a, 32'h4396fb07, 32'h438e813a},
  {32'h44edcac8, 32'h40834185, 32'h43aeab32},
  {32'hc4fb4a8b, 32'hc3f1d582, 32'hc3f7919c},
  {32'h4441fd06, 32'hc31b9495, 32'hc2ff891b},
  {32'hc4a33664, 32'hc34abf27, 32'hc36fbdfa},
  {32'h4513078e, 32'h4307ca64, 32'h420127a5},
  {32'hc5162143, 32'h421df704, 32'hc3b072df},
  {32'h43e4fa60, 32'hc3042560, 32'h4308e716},
  {32'hc4a0ec50, 32'hc3c611fc, 32'h43a2d207},
  {32'h44eb9489, 32'h4339a6c9, 32'hc2a8409d},
  {32'hc4a80df0, 32'hc3b8a588, 32'hc36b0568},
  {32'h44ec7462, 32'h43acba96, 32'h42be58bc},
  {32'hc375c7b6, 32'hc392d6a2, 32'h4307cc49},
  {32'h43e12758, 32'hc308ed7e, 32'h43839627},
  {32'hc48d2ba2, 32'hc331de09, 32'h4326b17a},
  {32'h44041b50, 32'h4354c85b, 32'h43232c12},
  {32'hc40f8f84, 32'h42ed7afe, 32'hc2d52e4a},
  {32'h44e417c2, 32'hc326e4a9, 32'hc2f47126},
  {32'hc3f3bf00, 32'hc37bbf35, 32'h41255eb2},
  {32'h44068ce4, 32'h41c462ab, 32'h43b222e7},
  {32'hc4eab2d4, 32'hc25adfd0, 32'h42fd051e},
  {32'hc0f2c200, 32'h44093fae, 32'hc3571a2a},
  {32'hc3a35a48, 32'hbfd77ee8, 32'hc3b52d36},
  {32'h43aadf1c, 32'h434c4740, 32'hc35e2888},
  {32'hc392512b, 32'hc2ab5182, 32'hc2b4d46a},
  {32'h450fc0ec, 32'hc369d154, 32'h43009a03},
  {32'hc49530bb, 32'h43818a9c, 32'hc246f2bd},
  {32'h43fa8ad4, 32'hc2379ee4, 32'h43034440},
  {32'hc44b7e47, 32'hc3905fe0, 32'hc2c230f8},
  {32'hc1f606b0, 32'h43938374, 32'h43c80e60},
  {32'hc48992e9, 32'hc41789af, 32'hc327d222},
  {32'h450a5883, 32'h42617bfd, 32'h421937f9},
  {32'hc4c93d77, 32'h40a6f16d, 32'h4335ab31},
  {32'h44a6e851, 32'h425a3a73, 32'hc4092b95},
  {32'hc3dfafe0, 32'h438c8ad6, 32'h432b8c75},
  {32'h449050ee, 32'h435c7b5a, 32'hc37db73b},
  {32'hc50a3d84, 32'h4348502c, 32'h439c666f},
  {32'h44a0d0c7, 32'hc180ddd4, 32'h43083957},
  {32'hc49e2ef5, 32'h433404e0, 32'hc1e01c22},
  {32'h4460a346, 32'hc39586e9, 32'h43df7dde},
  {32'hc4ab4438, 32'hc29c8f2c, 32'hc400b6f1},
  {32'h446b4e03, 32'h433ac30a, 32'hc2e5f05a},
  {32'hc48d518a, 32'hc33af90b, 32'h43a5b4ef},
  {32'h44808116, 32'hc2a78864, 32'h436c2a5f},
  {32'h43004464, 32'hc30e6ae2, 32'h4363a893},
  {32'h42f3bbb0, 32'hc1b80269, 32'h431f79ca},
  {32'hc4dfbbfd, 32'hc23d7ca4, 32'h43611ddf},
  {32'h44d997b5, 32'hbf73035e, 32'h4350641c},
  {32'hc4270a7a, 32'hc413e35b, 32'hc38bfed9},
  {32'h44562ff6, 32'hc2d10340, 32'h41d09956},
  {32'hc4ae2ae5, 32'h41406d06, 32'hc1ee7f0a},
  {32'h43f4e720, 32'h432b57d8, 32'hc3bb1593},
  {32'hc4e848a0, 32'hc191875d, 32'hc222a715},
  {32'h44de8133, 32'hc2c50f82, 32'h433bb924},
  {32'hc4e79ac7, 32'h4457219e, 32'h4352865e},
  {32'h44af89f8, 32'hc32a9587, 32'hc387f3ed},
  {32'hc45caeea, 32'hc30b8ceb, 32'hc3945979},
  {32'h45039da9, 32'h4351531d, 32'hc3423f90},
  {32'hc5102f93, 32'hc10aae1a, 32'hc3442f6b},
  {32'h433c62c4, 32'h4307f9ff, 32'h4315b036},
  {32'hc3e5f294, 32'h431b1afd, 32'hc3c6e3e2},
  {32'h44e54248, 32'hc3261948, 32'hc32d5c7b},
  {32'hc4d3d7ba, 32'h43868f35, 32'h41c464b3},
  {32'h44b69c48, 32'h43cefef1, 32'h42978179},
  {32'hc467cfb4, 32'h42b9798e, 32'hc270a8a8},
  {32'h446d99a4, 32'h43bb5c8f, 32'hc321d772},
  {32'hc4e9dc42, 32'hc23c1fe6, 32'hc3af4021},
  {32'h445cac82, 32'h43245dba, 32'hc2a1328c},
  {32'hc517fdb2, 32'h429c3c28, 32'h42fc5a8a},
  {32'hc34e66ea, 32'hc3e6e9bf, 32'h417cbb3d},
  {32'hc3251b70, 32'h43116716, 32'hc39aa2e7},
  {32'h44091262, 32'h4342fa5d, 32'hc1f1517f},
  {32'hc3785a8c, 32'h436fa760, 32'h4383b319},
  {32'h44951224, 32'h43d9c828, 32'h4113c42a},
  {32'hc504172f, 32'hc3275e11, 32'h42c46edc},
  {32'h44d497b9, 32'h4190a117, 32'h42e78888},
  {32'hc3e84178, 32'h4303cd67, 32'hc353dce6},
  {32'h43fa9c90, 32'h433881cf, 32'hc3b89ba8},
  {32'hc4415062, 32'hc39a56d8, 32'h42cbf343},
  {32'h44f5f8bd, 32'hc2c85713, 32'h42c57641},
  {32'hc4397850, 32'hc30d241c, 32'hc3ce7b35},
  {32'h45029012, 32'hc263b31d, 32'hc3cd2d0e},
  {32'hc41eb370, 32'h432a3fdf, 32'h43a50900},
  {32'h44db9f5e, 32'h41bc9129, 32'hc1c93808},
  {32'hc4428708, 32'hc210b284, 32'h428d0e2f},
  {32'h44ca8b77, 32'h42f4196c, 32'h431f9387},
  {32'hc4d314d0, 32'hc4000980, 32'hc28a9567},
  {32'h4511357b, 32'h4344d536, 32'hc30f4d67},
  {32'hc518a5b4, 32'hc37f9159, 32'h438434b7},
  {32'h44d56851, 32'hc2d99c1c, 32'h42d7126a},
  {32'hc4e932fa, 32'hc34bee6a, 32'hc2f77e99},
  {32'h4490ee62, 32'h4340fbe3, 32'h40e6302f},
  {32'hc4e01129, 32'h43e61d89, 32'h43ada48a},
  {32'h45067edc, 32'hc33f617f, 32'h42d310bc},
  {32'hc4e4042e, 32'hc3b018de, 32'h43049efc},
  {32'h4436eafa, 32'h424d4752, 32'h4289a604},
  {32'hc4a989f0, 32'h434ab168, 32'hc313cf58},
  {32'h446452cc, 32'hc39f7093, 32'h4323b9f7},
  {32'hc458a287, 32'h43910226, 32'h42ce8284},
  {32'h439da714, 32'h42c6a068, 32'h411bee02},
  {32'hc36f1530, 32'hc4366d07, 32'hc2e84d7b},
  {32'h428a3628, 32'h430aa6af, 32'h437c22e9},
  {32'hc40a6e60, 32'hc3a85166, 32'hc2e930ca},
  {32'h441c898a, 32'h438072bf, 32'hc2b59d8b},
  {32'hc5020c5c, 32'h42fb258c, 32'hc3623e32},
  {32'h4503d3c8, 32'hc0a51796, 32'h4317ac5f},
  {32'hc42ebdac, 32'h4173853e, 32'h43b2f68e},
  {32'h45130306, 32'h40c0a8c8, 32'hc1baaedc},
  {32'hc472c660, 32'hc03537c4, 32'h40d17d22},
  {32'h448ce0eb, 32'h439602ae, 32'hc38f1eb9},
  {32'hc4c78ee3, 32'h42c9ba5a, 32'h4335d3bf},
  {32'h4256fef8, 32'h429da813, 32'hc2e9ec66},
  {32'hc3f3f360, 32'h439b6571, 32'h438b21ff},
  {32'h44f00267, 32'hc3536223, 32'h4382dcd1},
  {32'hc4199884, 32'h43296533, 32'hc30a031a},
  {32'h44961cc3, 32'hc386cce5, 32'h438b59c5},
  {32'hc32431a0, 32'h437d35b3, 32'h433b1c0a},
  {32'h44d0e641, 32'h4116932a, 32'h43811f40},
  {32'hc336cfa3, 32'hc34e56c7, 32'h4389d277},
  {32'h44c1e0f2, 32'hc30d6678, 32'hc3b9ae63},
  {32'hc49b10d6, 32'hc3c6b843, 32'h3fd687c4},
  {32'h44805230, 32'hc2a2502f, 32'hc0233368},
  {32'hc50324eb, 32'hc308f849, 32'h42ac725c},
  {32'h4472a968, 32'hc2af9f01, 32'h4305f0a0},
  {32'hc50b5a8e, 32'hc27b6e58, 32'h4282444c},
  {32'h4503120e, 32'h42881579, 32'hc2d43f1c},
  {32'hc500dae1, 32'hc3812148, 32'h43d0a1af},
  {32'h44f82ac0, 32'h427ed690, 32'hc220831a},
  {32'hc46bbd7b, 32'hc2bed8b9, 32'hc3888927},
  {32'h44358fa7, 32'h41ce412a, 32'h42b02609},
  {32'hc398df65, 32'h43c5385b, 32'hc291fe8b},
  {32'h40a7bc00, 32'hc275870f, 32'hc183ba92},
  {32'hc4635852, 32'hc398babf, 32'h43a0de61},
  {32'h44f32d8e, 32'h42fe19fb, 32'hc2e90263},
  {32'hc42e07bd, 32'hc3b8716b, 32'h43c8a38f},
  {32'h449a7599, 32'h42934ff2, 32'hc1131072},
  {32'hc3f9ae58, 32'hc328006d, 32'h42337644},
  {32'h449ed5d0, 32'hc1d78ff9, 32'hc219eb20},
  {32'hc4e18085, 32'h40b7619e, 32'hc344c645},
  {32'h44e3f353, 32'hc20854ac, 32'hc38a96e6},
  {32'hc0173cc8, 32'h436e4919, 32'hc2b360d0},
  {32'h444add84, 32'hc230f596, 32'hc333c7e4},
  {32'hc4b50ce1, 32'h42b82feb, 32'h43c39aaf},
  {32'h449ab01c, 32'hc398be25, 32'h4346b4e4},
  {32'hc474d18a, 32'hc33eb49d, 32'h43d5e9a0},
  {32'h44d82436, 32'hc15e0965, 32'hc3c7f09f},
  {32'hc5105388, 32'hc398bdb7, 32'hc2d35aa5},
  {32'h44e87564, 32'hc3523d72, 32'hc372fe15},
  {32'hc43eee45, 32'h42bcfbdc, 32'h43df7b15},
  {32'h4311111c, 32'h435ef2ba, 32'h439ef465},
  {32'hc42e1480, 32'h43cb6342, 32'hc28fd0e0},
  {32'h451538cb, 32'h43b3a294, 32'hc396c2bc},
  {32'hc49466be, 32'hc04dd865, 32'hc3c2782e},
  {32'h44fd8d25, 32'h42dd105b, 32'h42769140},
  {32'hc4fbab84, 32'h418eb04b, 32'h4315173b},
  {32'h436dc722, 32'h4258ac46, 32'hc3c400a5},
  {32'hc42dfeda, 32'h43044e2a, 32'h43378813},
  {32'h45115b4b, 32'hc38a1894, 32'h42c14bc7},
  {32'hc4d6b347, 32'hc224c8e6, 32'hc33a817e},
  {32'h44c8c850, 32'h42c591c4, 32'h431f6f46},
  {32'hc4a7a6f1, 32'h43a59a74, 32'h4295338b},
  {32'h451a88d0, 32'h42e4e4c1, 32'hc395b3a5},
  {32'hc3861074, 32'hc38c92c2, 32'hc2bab8ce},
  {32'h4485dc2c, 32'h4119cf7d, 32'hc396f1ac},
  {32'hc48bc164, 32'h437e98b7, 32'hc3795700},
  {32'h447b4a82, 32'hbfae794d, 32'hc2d9b852},
  {32'hc4be03f6, 32'h4304fcb9, 32'h439ec24e},
  {32'h44d1bc36, 32'hc2f87b7f, 32'hc375deb4},
  {32'hc4cb09c1, 32'hc3397bb5, 32'hc3aa0097},
  {32'h450294e2, 32'hc389e143, 32'h4259497a},
  {32'h420e2133, 32'hc39ffea3, 32'hc17e538d},
  {32'h44efcc4b, 32'hc26cfbae, 32'h4256f91d},
  {32'hc2ab6c5e, 32'hc2f6f0b0, 32'h4322438b},
  {32'h44d30b52, 32'h4281e508, 32'h434676ff},
  {32'hc4f55445, 32'h4270731e, 32'h43666950},
  {32'h4309ede4, 32'hc2ad1dab, 32'h42a4758e},
  {32'hc349fc28, 32'hc3b44fba, 32'hc38fadd8},
  {32'h448f5db3, 32'hc3bb2c91, 32'h4298827a},
  {32'hc399247d, 32'h43181d22, 32'hc38dc43c},
  {32'h427373c0, 32'hc336efa3, 32'hc248764a},
  {32'h4494af9b, 32'h43021c41, 32'hc34d37f3},
  {32'hc3dc12c0, 32'hc198d0a1, 32'h42ada768},
  {32'h45159dee, 32'hc3865283, 32'h43426180},
  {32'hc41dcd80, 32'h433e893b, 32'h4350b32f},
  {32'h45046cad, 32'h419c7f12, 32'hc2cc58ae},
  {32'hc4121e6a, 32'h4323963e, 32'hc2861f05},
  {32'h45180c85, 32'hc31c857f, 32'h4306205e},
  {32'hc47429de, 32'hc34e04e3, 32'hc342f635},
  {32'h441e801b, 32'hc338431a, 32'hc40865af},
  {32'hc49c9589, 32'h440611a1, 32'hc301fdc4},
  {32'h44d0ee7f, 32'h423040f9, 32'h42d82a12},
  {32'hc43ad1a8, 32'h436462f4, 32'hc359ad94},
  {32'h449d3a91, 32'hc385f777, 32'h428e5662},
  {32'hc4db049a, 32'hc349bab5, 32'hc22208db},
  {32'h4390cc7a, 32'h433b9c3d, 32'hc360694b},
  {32'hc4a7372c, 32'hc337c48b, 32'hc36bf558},
  {32'h44a7fb7e, 32'h432849da, 32'hc38e288c},
  {32'hc43522b0, 32'hc0afcdb0, 32'h423aaf6f},
  {32'h4416ab6c, 32'hc26d1df0, 32'hc3db43a7},
  {32'hc4c8fc68, 32'h4330ead7, 32'h4038e8da},
  {32'h4206d040, 32'h43819950, 32'h42bf11e8},
  {32'hc4f83cbb, 32'hc2b62a4b, 32'hc322a76e},
  {32'h43ac93df, 32'hc3ac4205, 32'hc3275be6},
  {32'hc4c9e118, 32'h4225f9f5, 32'h4366adbc},
  {32'h43539670, 32'h430630ea, 32'h42f080cf},
  {32'hc427fd34, 32'h42667052, 32'hc311ca37},
  {32'h44f3dec3, 32'h434edb7a, 32'hc35c48c9},
  {32'hc506d8be, 32'hc37ed6c8, 32'hc2da822b},
  {32'h450eaee8, 32'h438bbe65, 32'h425c54da},
  {32'hc4f171cb, 32'hc360eabf, 32'hc2de8a74},
  {32'h4447e46c, 32'h43f632be, 32'hc2f1aef8},
  {32'hc5078789, 32'h42a2a665, 32'h43538040},
  {32'h44bb287b, 32'h4232ea0f, 32'h43d29ed0},
  {32'hc4a184d8, 32'hc34fb266, 32'hc237fb3d},
  {32'h4500c6b3, 32'hc330f1e3, 32'h438733d1},
  {32'hc47993ce, 32'h42399205, 32'h43aed1f0},
  {32'h44b8ec4c, 32'hc2bc062d, 32'hc35e3d37},
  {32'hc4d122ae, 32'h43a14231, 32'h41eb4bb2},
  {32'h45055f67, 32'h41954c50, 32'hc16b1e84},
  {32'hc3800240, 32'hc2018d20, 32'hc319b303},
  {32'h44e9d450, 32'h4315d2d8, 32'hc1af9ee4},
  {32'hc42247e6, 32'h425ea4e7, 32'h435a9578},
  {32'h44442215, 32'hc3d86607, 32'hc388e9b4},
  {32'hc52471d4, 32'h43199a93, 32'h420bf203},
  {32'h44f67519, 32'h431d2856, 32'hc3ba5cb9},
  {32'hc1f41100, 32'hc426fe8c, 32'hc2d73ce7},
  {32'h450a7c6f, 32'h4248d630, 32'hc2007bd2},
  {32'hc50baf95, 32'h432300ba, 32'h43a9fe62},
  {32'hc329fc3e, 32'hc2843e18, 32'h43334a5b},
  {32'h450aa203, 32'h424671ed, 32'h43733e61},
  {32'hc4a6dd7e, 32'h4324dc0e, 32'hc1c577e4},
  {32'h448804a1, 32'h4266ae6c, 32'h42f2d910},
  {32'hc4b4b146, 32'h429ae874, 32'h439acfac},
  {32'h449fe51a, 32'hc325c9f2, 32'h42d0dfb1},
  {32'hc4f6e1e9, 32'hc259a48c, 32'h42405615},
  {32'h450829df, 32'hc3c2d4fa, 32'hc2958d95},
  {32'hc4bef25b, 32'hc2d2a177, 32'h437144a1},
  {32'h443ed43b, 32'hc374f7b8, 32'hc3bbb0b7},
  {32'hc4e48eee, 32'h438c0d2d, 32'hc2f96266},
  {32'h447cd9d3, 32'h432425b0, 32'h4364a098},
  {32'hc3b808c4, 32'hc1810b7d, 32'hc3446ced},
  {32'h44a1194f, 32'hc393d9a7, 32'hc3849feb},
  {32'hc463bc2c, 32'hc19a69fc, 32'h43732578},
  {32'h44cd6b7c, 32'h43a9aab6, 32'hc36e2d6f},
  {32'hc507dc2f, 32'hc23a9468, 32'hc32d1e91},
  {32'h45040199, 32'h43b5e3a3, 32'hbfe447c1},
  {32'hc41d5916, 32'h423c3272, 32'h4336097f},
  {32'h44aeed2b, 32'h42f1c734, 32'hc1ddfc96},
  {32'hc4b49ab4, 32'h415b0d40, 32'h42ccfc0e},
  {32'h45088e91, 32'h434fb743, 32'hc3b42c8e},
  {32'hc5006f31, 32'h42690b50, 32'h43acfa4d},
  {32'h450b3f04, 32'h4402ae43, 32'h43b29140},
  {32'hc5134e41, 32'hc327e82e, 32'h42176434},
  {32'h4363f670, 32'h421f344c, 32'hc2bc7f86},
  {32'hc313aa88, 32'hc28e7fbf, 32'h42e7e8b8},
  {32'h44c605ed, 32'hc3066c40, 32'hc3ee65b4},
  {32'hc4a1e884, 32'h4292c638, 32'hc2e8d29f},
  {32'h4519d60e, 32'h42b6349f, 32'h3f4a2d37},
  {32'hc4b1099c, 32'hc35801a7, 32'hc3a1d4fa},
  {32'h45140b8d, 32'hc1e444fe, 32'hc33cfac1},
  {32'hc50aaf22, 32'hc1ad2413, 32'h43949d92},
  {32'h445b9bcd, 32'h44090c2a, 32'h430850e6},
  {32'hc325bf16, 32'h42e22a92, 32'hc2586fe0},
  {32'h444aa753, 32'h430df5f8, 32'h42b9f593},
  {32'hc46f3bf2, 32'h43532cd0, 32'h435112cd},
  {32'h452169b8, 32'hc2df9060, 32'hc0b92138},
  {32'hc4c6fd42, 32'h438f6528, 32'hc273c578},
  {32'h44a169c8, 32'hc3fe5ce1, 32'h43cc1500},
  {32'hc3e11080, 32'h4387be5f, 32'h42da0ee1},
  {32'h4514a18c, 32'h43460567, 32'hc3478efe},
  {32'hc425dd00, 32'h4323a5ed, 32'h432bb45b},
  {32'h44a797fe, 32'hc30bdb51, 32'h41c15476},
  {32'hc5043d73, 32'hc2a58653, 32'h43bf165e},
  {32'h42a49a70, 32'h4406ef35, 32'hc3e1740d},
  {32'hc29773a0, 32'hc3cd9179, 32'h4340585d},
  {32'h4491f389, 32'h430ff3b3, 32'hc25e423e},
  {32'hc44b827a, 32'hc40cd645, 32'h41553f58},
  {32'h44f90bac, 32'hc276d43f, 32'h42df04c9},
  {32'hc4a5bd0c, 32'hc3d3b67a, 32'hc3105ace},
  {32'h4328b868, 32'h438f1870, 32'hc3769484},
  {32'hc51c9932, 32'hc35ce698, 32'hc145f98c},
  {32'h44e14f11, 32'h42a6bed4, 32'h436400a2},
  {32'hc4bcd2af, 32'hc2ead98d, 32'h42610160},
  {32'hc50537e9, 32'hc32c6ae0, 32'hc315931d},
  {32'h4421f650, 32'hc3be13af, 32'h43a3305a},
  {32'hc44123dc, 32'hc2457f40, 32'hc3196ee2},
  {32'h44cd7582, 32'hc11a6ffd, 32'hc25d3099},
  {32'hc4bce8df, 32'h43bc375b, 32'hc3fa8532},
  {32'h43334560, 32'h431bfcce, 32'hc3535845},
  {32'hc1df0faf, 32'hc2120b7e, 32'h42ba4456},
  {32'h45149e10, 32'hc1b5c114, 32'hc2d1f3f8},
  {32'hc4a04b6a, 32'h421ed54c, 32'hc39375c0},
  {32'h450d4717, 32'h42df124e, 32'h43bc6711},
  {32'hc2a43040, 32'hc2fb5c32, 32'hc2dc0074},
  {32'h45152b22, 32'hc10cd9f2, 32'hc325256b},
  {32'hc3e4d460, 32'hc344c555, 32'hc3328cab},
  {32'hc2470680, 32'h43a756ec, 32'h43ac8c77},
  {32'hc4822f7d, 32'hc2c5ab47, 32'hc35dae23},
  {32'h45132731, 32'h43277462, 32'hc29067d0},
  {32'hc4567726, 32'h433dd056, 32'h427a46b7},
  {32'h442e6b0c, 32'hc4080c2f, 32'h431174ff},
  {32'hc4849b1e, 32'hc32d30c1, 32'h412c2293},
  {32'h448a5b91, 32'h434de12e, 32'hc3693faa},
  {32'hc4660ed6, 32'hc2fd7722, 32'h423b1bca},
  {32'h44918a22, 32'h417fcddc, 32'hc2dc7205},
  {32'h43de51dc, 32'h43883c1c, 32'hc43ba045},
  {32'h44fa2ce0, 32'hc1946c34, 32'h4269f278},
  {32'hc4425378, 32'hc1799e33, 32'h407b4068},
  {32'h44eb526e, 32'h4345e8fc, 32'h40cc093e},
  {32'hc4c26e6e, 32'hc2b2f5a3, 32'hc3bf5980},
  {32'h44a63560, 32'hc39ba62e, 32'h43f0610b},
  {32'hc4263c23, 32'h429f1497, 32'h42a67094},
  {32'h44d7e50e, 32'h42b4a0cc, 32'hc3e8a245},
  {32'h41c4f5b0, 32'hc2e416ce, 32'hc3a2d1f9},
  {32'h43ac5850, 32'h433fff4f, 32'hc2c31189},
  {32'hc29e942c, 32'hc32e5d15, 32'h42104e3d},
  {32'h44b7654c, 32'hc39a28d0, 32'h4381a888},
  {32'hc4bede3d, 32'h432c4567, 32'h43d82bde},
  {32'h44020e28, 32'hc31dc133, 32'hc2aee1dc},
  {32'hc3c18ba4, 32'hc2b13100, 32'hc3ff0b32},
  {32'h4491e932, 32'hc1ebd432, 32'hc2f8c4a7},
  {32'hc504b0b0, 32'hc23ca8cf, 32'hc3357e72},
  {32'h43fc494d, 32'h40ddd2e2, 32'h447c42ab},
  {32'hc503f5f2, 32'hc3a6fc33, 32'hc2f5cc51},
  {32'h45032493, 32'h438e65c2, 32'h43686187},
  {32'h4486d8bc, 32'hc3b87934, 32'h42f9c3ae},
  {32'hc4893f3e, 32'h4193eadb, 32'hc3680d82},
  {32'h449a8ea2, 32'h437a3374, 32'h43acaea3},
  {32'hc3db4040, 32'h434afcae, 32'hc211de75},
  {32'h43ddd9e1, 32'h4197f4f2, 32'h42f65a90},
  {32'hc4ebd090, 32'hc306cf5f, 32'hc2ed14d7},
  {32'h45009824, 32'hc34c33b2, 32'h42490e0d},
  {32'hc45fe4c5, 32'hc202ebde, 32'h434d3ac8},
  {32'h43c0ffc2, 32'h420ce061, 32'h43b16e4f},
  {32'hc3bf2640, 32'hc2c4982d, 32'hc2902320},
  {32'h44285fb2, 32'hc225f1dc, 32'hc2f5f84f},
  {32'hba000000, 32'hc3a21686, 32'h428b875d},
  {32'h4507789a, 32'hc39eb6bc, 32'h41f818f9},
  {32'hc43d25c7, 32'hc2fb4e87, 32'hc2cfabe3},
  {32'h44f61dd6, 32'h438ace2d, 32'h43a9e972},
  {32'hc503befb, 32'hc318b53a, 32'h41d0e78a},
  {32'h4505347a, 32'h427941da, 32'h43bed92d},
  {32'hc4299139, 32'h43445a91, 32'hc34a2cd4},
  {32'h427dd100, 32'hc2a4a018, 32'h4297fe4f},
  {32'hc4a51a8e, 32'hc3981a71, 32'hc35f9782},
  {32'h45019cdc, 32'hc39ff558, 32'h4301d182},
  {32'hc3d78474, 32'h41c61798, 32'hc343687f},
  {32'h446bca1b, 32'h42f159f1, 32'h43a91087},
  {32'hc41236cb, 32'hc3ea3487, 32'hc382a321},
  {32'h445800a4, 32'h433473af, 32'hc172558c},
  {32'hc4ba5e27, 32'hc2cd1e25, 32'hc2493245},
  {32'hc16a8d9c, 32'hc3689bac, 32'hc2f09920},
  {32'h44e25da2, 32'hc31a5a47, 32'h43794ccb},
  {32'hc4c206b7, 32'hc0a45d60, 32'hc3c1b5b6},
  {32'h44c63910, 32'h4289e5a5, 32'hc3682821},
  {32'hc4ea9181, 32'h4292fcf1, 32'hc3833b33},
  {32'h446c2e7d, 32'hc28e737f, 32'h44119709},
  {32'hc3ab6c68, 32'hc3d1b23c, 32'hc4290cbd},
  {32'h44690406, 32'h43363ceb, 32'h420c6052},
  {32'hc5055c29, 32'hc10f0753, 32'hc36c8897},
  {32'h43677841, 32'hc328197d, 32'hc3af05dd},
  {32'hc47ca8ba, 32'h43358060, 32'h426527f8},
  {32'h43f82780, 32'h43a120e5, 32'h436f7376},
  {32'hc3f37ed6, 32'hc36a39e9, 32'hc3f0dfcc},
  {32'h451589d6, 32'hc40189af, 32'h440e38b1},
  {32'hc4e9f6f4, 32'h4339daf6, 32'hc34a6283},
  {32'h45058102, 32'hc3638bdb, 32'hc2911338},
  {32'hc4f44893, 32'h42f47eec, 32'hbfaf7090},
  {32'h4507decb, 32'h4393822a, 32'hc3ae6963},
  {32'hc4afccf7, 32'h4363eb00, 32'h3ecf8204},
  {32'h4478f08b, 32'hc1d9cffc, 32'h43a7664a},
  {32'hc416ffbc, 32'hc3787e63, 32'hc35a6e52},
  {32'h44ef38a9, 32'h41e65f27, 32'h432d520c},
  {32'hc4e3e7cf, 32'h430cc517, 32'hc31db988},
  {32'h44edc2f3, 32'hc1156c17, 32'h41535e75},
  {32'hc34a6520, 32'hc30c8d30, 32'hc34f1745},
  {32'h43ad99dc, 32'hc3ce9768, 32'h42b72496},
  {32'hc385aa0a, 32'hc2e2c1cc, 32'hc3529558},
  {32'hc3faa3b4, 32'hc3d24925, 32'h43b2cc84},
  {32'hc4c35c66, 32'h423318a4, 32'hc3c04b69},
  {32'h42fc56c0, 32'hc3462a3b, 32'h43955a56},
  {32'hc4ff46d1, 32'hc3326195, 32'h42b505fd},
  {32'h44ead1aa, 32'hc3b537a1, 32'hc3b77584},
  {32'hc4ff3602, 32'h42880eec, 32'hc3ff97b7},
  {32'h44f9783a, 32'hbfedfbfb, 32'hc0c0402c},
  {32'hc3e1a1d0, 32'hc32420a2, 32'hc385df3a},
  {32'h45096884, 32'hc368b63e, 32'hc34dcf55},
  {32'hc4fda006, 32'hc2b53859, 32'h4375a9ad},
  {32'h44eb7f84, 32'h424f44f8, 32'h4302d27f},
  {32'hc480bce4, 32'hc2cf6de6, 32'h42fda7ff},
  {32'h447eb96a, 32'hc38342e5, 32'hc30969ef},
  {32'h4469a818, 32'h4381fd67, 32'hc2d20dd7},
  {32'hc4453f97, 32'h401ecdf3, 32'hc3c65c65},
  {32'h43a34aa0, 32'hc3232f0a, 32'h428d05f6},
  {32'hc4d96f28, 32'hc2cafd46, 32'hc3edc239},
  {32'h441f3bd4, 32'h42fbd5d9, 32'h43af57cb},
  {32'hc2cb4ac0, 32'hc291563c, 32'hc35880dc},
  {32'h4504b019, 32'h42906840, 32'h43b77824},
  {32'h42df2c71, 32'h4390914c, 32'hc3a78f4e},
  {32'h4426c82c, 32'hc3a75b64, 32'h42aa9d3d},
  {32'hc4ed438f, 32'h41cae9ae, 32'h4319ab8b},
  {32'hc2c44d1a, 32'hc398a5b5, 32'h3fc27505},
  {32'hc41eae38, 32'hc4086452, 32'h3e037f80},
  {32'h4435a474, 32'hc287a4fd, 32'h43ec0917},
  {32'hc3cbcdcc, 32'h431a3830, 32'hc1e896d7},
  {32'h44e9f056, 32'hc324c62a, 32'hc4165a1c},
  {32'hc4c2bc0d, 32'hc331606f, 32'h43dfa54b},
  {32'hc4e67ef2, 32'h43982d1d, 32'hc3c764e8},
  {32'h43147720, 32'hc3c76205, 32'hc391ebc9},
  {32'hc465d429, 32'hc3c17c26, 32'hc256410b},
  {32'h450e36af, 32'hc379c007, 32'h43dea243},
  {32'hc4f4b3b9, 32'h42319628, 32'h41895dc3},
  {32'hc50a02da, 32'h432b593f, 32'hc3567dd3},
  {32'h43c345c1, 32'h4383004d, 32'hc26fc0a4},
  {32'hc4bef6b0, 32'h43976b70, 32'h43608eca},
  {32'h44f6b0e4, 32'h41c87c5e, 32'h42c1cb89},
  {32'h43e5325b, 32'h438f3e21, 32'hc2ca62cc},
  {32'h45035a17, 32'hc2e3fd53, 32'h43b442f8},
  {32'hc4c63c89, 32'hc2ab5d39, 32'h425595fc},
  {32'h43e00ab8, 32'hc2dfcfd2, 32'h43169e82},
  {32'hc3d68cc7, 32'hc3ab7d1a, 32'hc3d3ee29},
  {32'h442f9aa6, 32'h431fac90, 32'h41e53d33},
  {32'hc4bdddce, 32'h40dbbb7e, 32'hc328e76c},
  {32'h449b54d0, 32'h42c7d970, 32'h42744bd1},
  {32'hc2fca318, 32'h42c5c661, 32'hc32a72f2},
  {32'h44fea8b4, 32'hc3a726c1, 32'hc2824026},
  {32'hc5011379, 32'hc27888fa, 32'h430258e7},
  {32'h450720f2, 32'hc33cf29f, 32'h442af56d},
  {32'hc3ed02f4, 32'hc2891787, 32'h43084357},
  {32'hc45de45a, 32'hc3897cfa, 32'h43bb917e},
  {32'h44eef3c2, 32'h42f086ae, 32'hbfb183c0},
  {32'hc4fad3d2, 32'h4372b6bc, 32'h40e58f02},
  {32'h45048a50, 32'h41272674, 32'hc2f27f7c},
  {32'h42065f40, 32'h4308be1a, 32'h43a6be3d},
  {32'h4501f479, 32'h4126453c, 32'hc206a942},
  {32'hc488974f, 32'hc422e12b, 32'h43c99c08},
  {32'h44a9959f, 32'h4348f038, 32'hc30953dd},
  {32'hc4f91e0e, 32'hc3be38fb, 32'h43083636},
  {32'h44de521f, 32'hc35722d4, 32'h430e5474},
  {32'hc5134fc6, 32'hc23263e2, 32'hc2e3792a},
  {32'h43f3e5a8, 32'hc34f3c3e, 32'h4216834a},
  {32'hc50fa488, 32'hc321b975, 32'hc4294557},
  {32'hc3415ef2, 32'hc30f6127, 32'h421c5b29},
  {32'hc46b0d80, 32'h43ace5a9, 32'h4320425b},
  {32'h44d542ab, 32'h43262dac, 32'hc225c31c},
  {32'hc47b8bf4, 32'hc409cf28, 32'h433351c7},
  {32'h44bfdbc4, 32'h419d6c92, 32'h43f1e23d},
  {32'hc3a05e98, 32'h43573187, 32'h42db32a7},
  {32'h43d344bb, 32'h42fec698, 32'hc35cad70},
  {32'hc4b5b2e8, 32'hc3789712, 32'hc2a70172},
  {32'h44609e04, 32'h42fd8a18, 32'h42a5dba8},
  {32'hc509bee8, 32'h410c5068, 32'h43cb3001},
  {32'h44df31a8, 32'h42c3d05d, 32'hc31511a0},
  {32'h43a28c13, 32'hc2c9a31a, 32'hc2fcb899},
  {32'hc30145b0, 32'hc30c46b1, 32'h4279be8c},
  {32'hc4a62301, 32'hc205f9d0, 32'hc268295e},
  {32'h4419055a, 32'h43c05a17, 32'hc1dd034d},
  {32'h438516ea, 32'hc4067e66, 32'h43801d6a},
  {32'h4408c088, 32'h438281ee, 32'hc1d24552},
  {32'hc4afa685, 32'h43b00c8c, 32'hc36431a1},
  {32'h44ff7d4a, 32'hc2dd705d, 32'h42f71512},
  {32'hc490bf27, 32'h41fb2803, 32'h4394b48d},
  {32'h44dffab6, 32'hc3a42442, 32'hc2889d8f},
  {32'h4413867a, 32'hc36afc78, 32'hbfb638a8},
  {32'hc44ba226, 32'hc31fcba6, 32'h4311369d},
  {32'h44797b44, 32'h4290a20d, 32'h426c4a52},
  {32'hc4d20805, 32'hc3dfb87a, 32'h42bc5cf9},
  {32'h4427807c, 32'hc382a009, 32'h4320539b},
  {32'hc373c718, 32'h4358508f, 32'h43693cc6},
  {32'h44c521ec, 32'hc3222ea2, 32'hc2297e8a},
  {32'hc3c843a0, 32'h402b389a, 32'h431c0b73},
  {32'h44e66ee2, 32'h43377ffa, 32'h4391c718},
  {32'hc38c6188, 32'h4392bbf4, 32'h43a05c0b},
  {32'h44defa01, 32'hc2acff91, 32'hc11164c5},
  {32'hc48146f4, 32'hc30974d9, 32'h4291d165},
  {32'hc298f580, 32'h4262d883, 32'hc3879e84},
  {32'hc499ef68, 32'h433a280f, 32'hc32ad405},
  {32'hc4098d1c, 32'h431940d1, 32'hc39730f1},
  {32'h434c6318, 32'h41057a4e, 32'hc270dd66},
  {32'hc3e0f7c8, 32'h439fb22a, 32'hc3a3735b},
  {32'h446a46dc, 32'hc21db2ea, 32'hc228056d},
  {32'hc5205cd9, 32'hc1bc8fea, 32'hc407a602},
  {32'h447f0924, 32'h434c2dca, 32'h42aeb750},
  {32'hc4ebbe43, 32'hc3777d07, 32'h43317bb7},
  {32'h44bd34ff, 32'h4387bdc0, 32'h425525bc},
  {32'hc44b2228, 32'hc2e3b05a, 32'hc3518fea},
  {32'h44a60281, 32'h43bb734d, 32'h426f2054},
  {32'hc482a4b0, 32'hc35ec684, 32'h44270468},
  {32'h4501578f, 32'hc3c65a1f, 32'hc3b35e72},
  {32'hc4c2d8c6, 32'hc303c453, 32'h3ff279f8},
  {32'h44933650, 32'h43353fe3, 32'h4316c53a},
  {32'hc46a1acf, 32'hc3ea0288, 32'h44040365},
  {32'h44341621, 32'h43c407fd, 32'hc387e112},
  {32'hc4e5c6d5, 32'hc2dce150, 32'h439786e8},
  {32'h4509b7a8, 32'h43a1ad00, 32'hc1f8a6cd},
  {32'hc48d0dd8, 32'hc301ea8a, 32'h434befdf},
  {32'h43bef4db, 32'hc2c25795, 32'hc2e56432},
  {32'hc5073175, 32'h43a3696a, 32'h43ef048e},
  {32'h451fda69, 32'hc186643e, 32'hc3646683},
  {32'hc4b35cd6, 32'hc201d738, 32'hc2f402cc},
  {32'h44fe2e61, 32'hc3272f8d, 32'h41e6e189},
  {32'h41313e00, 32'h428a722c, 32'h439494f8},
  {32'hc23fb300, 32'h42fc52bd, 32'hc3eb77f6},
  {32'hc497631f, 32'h42856d70, 32'hc3409446},
  {32'h4491d304, 32'h41968718, 32'hc2158f02},
  {32'hc4f47463, 32'h41c72c70, 32'h42d8bcd7},
  {32'h448bffde, 32'hc32169ad, 32'hc33950d1},
  {32'h446657b8, 32'hc29ae58e, 32'hc1e15ad4},
  {32'hc491b4ef, 32'hc251ab22, 32'hc318a322},
  {32'h43bd098a, 32'h42b6557d, 32'hc3082f79},
  {32'h425e39e6, 32'h43d211fd, 32'hc2482d25},
  {32'h445ab172, 32'hc27f2fe6, 32'hc31f656b},
  {32'hc50035fc, 32'hc1089e94, 32'hc2fc1cfb},
  {32'hc3273960, 32'hc28b5506, 32'h42d340f6},
  {32'hc49a2436, 32'hc1fc238c, 32'hc3a40916},
  {32'h44886250, 32'hc37a5ae0, 32'h42eedf28},
  {32'hc48ff132, 32'h439fc84a, 32'h4058d6f8},
  {32'h4470da26, 32'hc335e2e4, 32'hc3173798},
  {32'hc39a4cc0, 32'hc2aef0d9, 32'hc3899578},
  {32'h4504df09, 32'h43544046, 32'h42a6b4c1},
  {32'hc4d9f220, 32'h42a78faf, 32'h408c2313},
  {32'h440a394c, 32'h42eae25e, 32'hc2e8eb8b},
  {32'hc45a9afc, 32'h42fcdce7, 32'h439ebf6b},
  {32'h4430fa56, 32'h43dbd8fd, 32'h41ad5158},
  {32'hc305bbfd, 32'hc380caec, 32'h4224f560},
  {32'h44a46c48, 32'h43cb33a6, 32'hc395e2e9},
  {32'hc49f1400, 32'hc396946f, 32'h425fa4cf},
  {32'h4426a6ab, 32'h42899dee, 32'hc3e3e678},
  {32'hc45bed55, 32'hc337112e, 32'hc35de011},
  {32'h44a7da1d, 32'h425898fc, 32'h43b0b3c0},
  {32'hc502ccc3, 32'hc3163d2d, 32'hc3004b2e},
  {32'h44ec9364, 32'h442a5f6a, 32'h41f7515d},
  {32'hc4a3e119, 32'hc1e5ed02, 32'hc287ce99},
  {32'h437406bb, 32'h405c283f, 32'h43e53084},
  {32'hc4a70d61, 32'hc1f998e0, 32'h43ef66ed},
  {32'h4419d1e0, 32'h42beebf0, 32'hc3a5481b},
  {32'hc5067e29, 32'h41019536, 32'hc342d4a6},
  {32'h44a04b73, 32'hc2eed520, 32'h42a9ba29},
  {32'hc4a5e597, 32'h43676287, 32'h433d15fe},
  {32'h4423ca1c, 32'hc29aa324, 32'h429e49a2},
  {32'hc47c00b9, 32'hc2de2a22, 32'hc249ac42},
  {32'h44e7c010, 32'hc2bd9c10, 32'h436376a7},
  {32'hc38c4fb0, 32'hc2b76600, 32'hc2eabc28},
  {32'h442d0282, 32'h423a0394, 32'h4380455d},
  {32'hc4de08f3, 32'hc40d0a9a, 32'h43451bd1},
  {32'h450cd17d, 32'h43af2c76, 32'hc1ca0130},
  {32'hc4742892, 32'h42fa250c, 32'h41900b12},
  {32'h44e9dbc0, 32'hc275771d, 32'hc3b46bba},
  {32'hc4036659, 32'h428d1778, 32'hc26eb0bd},
  {32'h44ad58a5, 32'h42fd5c06, 32'hc30a51a6},
  {32'hc4535b88, 32'h431c4d67, 32'h433241ff},
  {32'h44b9ee74, 32'hc2ce15d2, 32'h4389d838},
  {32'hc4f29b35, 32'h43cfdbf1, 32'hc3842dda},
  {32'h44e007e2, 32'hc34c232d, 32'hc2a9c765},
  {32'hc4ac3f2b, 32'h4389aab1, 32'hc3b6caca},
  {32'hc3096284, 32'hc313f32d, 32'h40a4167e},
  {32'hc41dc276, 32'h42efd8ce, 32'h40b93696},
  {32'h44c1ce9b, 32'hc18fec1e, 32'hc312b545},
  {32'hc4d2a916, 32'h42994bba, 32'h426d2f31},
  {32'h45085948, 32'h42c637fa, 32'h42f77e0b},
  {32'hc44f5520, 32'hc3ab9185, 32'hc3c9adf8},
  {32'h44f66fd0, 32'hc2d98a1c, 32'hc3260d62},
  {32'hc44a72f6, 32'hc3db6058, 32'h43000ecb},
  {32'h445ad32f, 32'h4271ceb8, 32'hc0847465},
  {32'hc4fe1377, 32'h4248178f, 32'hc3145030},
  {32'h43924335, 32'h43c1679e, 32'hc31ff49a},
  {32'hc482ce28, 32'h438f05b8, 32'h42fd62e1},
  {32'h44b1a240, 32'h431a74cd, 32'hc31d7a1a},
  {32'hc4429e0f, 32'h41e68064, 32'hc2c6a125},
  {32'h450057d1, 32'hc3e88921, 32'hc30c0b89},
  {32'hc4f9b035, 32'h42bceda1, 32'h42b89395},
  {32'h44ac1b49, 32'h430d217f, 32'hc267f4b0},
  {32'hc4d1d224, 32'h42933ce5, 32'hc3c51efd},
  {32'h4491068e, 32'hc3693065, 32'h415668ef},
  {32'hc4aa95ae, 32'hc2e9ce7c, 32'hc2d46de2},
  {32'h445065a1, 32'h428eb8ee, 32'hc2c11462},
  {32'hc430631a, 32'hc3acfb6e, 32'hc12fb133},
  {32'h443c3ca5, 32'h42802716, 32'hc39acbe8},
  {32'hc50bfeed, 32'hc2cbd62f, 32'hc2d3bd4a},
  {32'h44ed1b87, 32'hc2534ae0, 32'h42c233f3},
  {32'hc4227870, 32'h437c0213, 32'h4331de59},
  {32'h4364a736, 32'h43780bfb, 32'h42f03d69},
  {32'hc501aee5, 32'hc3812435, 32'hc35d3b72},
  {32'h44945436, 32'hc3999b86, 32'hc2eb400b},
  {32'hc4a0009a, 32'h425b891e, 32'hc34ed50e},
  {32'h44980b04, 32'hc19e756f, 32'hc3ee4bfb},
  {32'hc4c47700, 32'h436edfe0, 32'h4397809a},
  {32'h44d4a2fa, 32'hc3853038, 32'h431e4069},
  {32'hc3248fc0, 32'hc2ba2cbb, 32'h43be4355},
  {32'h41cb3d80, 32'h439e4b3a, 32'h438924c3},
  {32'hc28abb30, 32'hc38473f9, 32'h42dfe9f3},
  {32'h44e4ab0e, 32'hc424e2ec, 32'hc3a03ce9},
  {32'hc49773f8, 32'hc309d4d8, 32'hc2978898},
  {32'h4462b4f8, 32'h4366b940, 32'hc318d12d},
  {32'hc51060fa, 32'h4247f4cc, 32'h430acd1b},
  {32'h450580c5, 32'h433cf5ca, 32'h43275657},
  {32'hc404ba8e, 32'hc2aa5389, 32'h42d4021c},
  {32'h44fbfc50, 32'h42312717, 32'h437aa13d},
  {32'hc4f8da00, 32'h434d7b3b, 32'hc2da4a2a},
  {32'h44f505ca, 32'h433eac4a, 32'hc17f35f6},
  {32'hc47158ec, 32'hc215cf77, 32'hc323c594},
  {32'h440cbea6, 32'h43735c07, 32'hc335c98e},
  {32'hc4e0a786, 32'hc1ca0f99, 32'h42ed25b0},
  {32'h450704c8, 32'h4220fd28, 32'h420be457},
  {32'hc5148d76, 32'hc2f6f1bf, 32'h41d54b04},
  {32'h45035011, 32'h432258e9, 32'hc36777f6},
  {32'hc4d68f92, 32'hc3dd6bb0, 32'h432d2a9a},
  {32'h43d551ba, 32'hc27c0280, 32'hc13e4a72},
  {32'hc4b74799, 32'hc290437e, 32'hc3580db4},
  {32'h4400043a, 32'h4389a77e, 32'h432abf8c},
  {32'hc4b42ca7, 32'h43953c3a, 32'hc2cca744},
  {32'h4489a1a8, 32'h4392e605, 32'h42aae587},
  {32'hc50b0a5c, 32'hc3a91cf7, 32'h42d6e00c},
  {32'h449e7d70, 32'hc37933da, 32'h429c1256},
  {32'hc44512fc, 32'h42aab6a2, 32'h417db640},
  {32'h443d3d00, 32'h421c311a, 32'hc28e0cd7},
  {32'hc4362218, 32'h42ed63bc, 32'hc3b53eea},
  {32'h4518a9d1, 32'hc24a69fd, 32'hc3613279},
  {32'hc50db3f7, 32'hc2cadeec, 32'h428fd355},
  {32'h450b0e66, 32'hc2752195, 32'h4290abd5},
  {32'hc4b8a726, 32'h43d90671, 32'hc291c8cb},
  {32'h43c97d4d, 32'h438e28e4, 32'h4304f672},
  {32'hc5040e06, 32'h434c7364, 32'hc411895e},
  {32'h43b82626, 32'h434481d7, 32'h422d2c47},
  {32'hc4e99282, 32'h42e6a07d, 32'h40f87308},
  {32'h44f1f534, 32'hc3838fcd, 32'hc32382ba},
  {32'hc401e94d, 32'h435bb70c, 32'hc24031b2},
  {32'h44b7cb84, 32'hc0034d82, 32'hc1fccc1f},
  {32'hc4820478, 32'h43e4923c, 32'h428d74b3},
  {32'h43a4c31a, 32'hc2d095a0, 32'h437990a7},
  {32'hc38db2c0, 32'h43823528, 32'h4323fba8},
  {32'h4414b987, 32'h433b4628, 32'hc3a0795c},
  {32'hc401e6b4, 32'h42d9118e, 32'h4344ebca},
  {32'h43dfa29b, 32'hc2d6d32f, 32'hc34c0897},
  {32'hc3741fb0, 32'h421abad2, 32'hc2a6ffba},
  {32'h445a1214, 32'hc3a9d0af, 32'h423c175e},
  {32'hc478ba1d, 32'hc2d5b6fd, 32'hc356c2d0},
  {32'h44883952, 32'hc12114ac, 32'h43ab2616},
  {32'hc14f4500, 32'hc3365c5c, 32'h4349ce41},
  {32'h4437aa7c, 32'hc014e009, 32'h41d977b8},
  {32'hc47b945c, 32'h43bcee8e, 32'h431404bd},
  {32'h44f7a9bc, 32'h43e94c90, 32'h42df7b4e},
  {32'hc48bb5d1, 32'hc31a599d, 32'hc16483e1},
  {32'h4513635b, 32'h42a11d37, 32'hc3a3ef01},
  {32'hc4c9828b, 32'hc3a77086, 32'h4314057f},
  {32'h44aa1e1c, 32'hc23fae4e, 32'hc37a6d10},
  {32'hc40f6a40, 32'hc326f4d5, 32'hc37f3432},
  {32'h45172f6a, 32'hc2c67ebc, 32'hc32b66e7},
  {32'hc5098fb7, 32'h4231e4e4, 32'hc317ebaa},
  {32'h44e840a9, 32'h43bc2df8, 32'h42f50d90},
  {32'hc4cb5369, 32'h438ca8c1, 32'hc3560dcd},
  {32'h450b6842, 32'h420522b5, 32'hc2e3bdfc},
  {32'hc4c5fe91, 32'h43095ae2, 32'hc24f5f8f},
  {32'h44ac47a8, 32'h437ce2ac, 32'h431fc3ed},
  {32'hc4cee843, 32'hc364eefa, 32'h4316563d},
  {32'h41fcf2a0, 32'h4358a72a, 32'hc2e06e34},
  {32'hc4b5c6ab, 32'h4325285d, 32'hc286cf1a},
  {32'h44f8ec50, 32'hc3e1c708, 32'h439719e9},
  {32'hc4ae6cee, 32'hc325cdd3, 32'h43023103},
  {32'h45007f84, 32'h438ea6e2, 32'h436e19d6},
  {32'h4211f584, 32'h429bde53, 32'h42c3c144},
  {32'h44a6effc, 32'hc383e3a8, 32'h4339aa08},
  {32'hc4137f0a, 32'hc3c0bd6f, 32'hc2d26134},
  {32'h44bb1842, 32'h4311a643, 32'h4389cad7},
  {32'hc49bde6e, 32'h428508f4, 32'hc3940cfe},
  {32'h44bcee47, 32'hc32db808, 32'h44256f58},
  {32'hc48d32e2, 32'h436c1d70, 32'hc2e31018},
  {32'h44f74e1d, 32'hc3d722a7, 32'hc39578a6},
  {32'hc4b9fb50, 32'hc2d5f90a, 32'h431403b5},
  {32'h43cab590, 32'h42ded403, 32'h42cc3463},
  {32'hc4de2fc6, 32'h4339ce4f, 32'h42589a8f},
  {32'h44b9b6e4, 32'h43478314, 32'h42de6381},
  {32'hc4e2d771, 32'h42190cc3, 32'hc2880035},
  {32'h44a91294, 32'h42ec858a, 32'hc23ddb87},
  {32'hc510fad9, 32'hc36ea754, 32'hc31152ad},
  {32'h4497a763, 32'h42a113a3, 32'h429adb48},
  {32'hc278e7ff, 32'hc3b1350d, 32'h43811b7a},
  {32'h448c1037, 32'h434d3497, 32'hc30d7fa8},
  {32'hc4c13abc, 32'hc1f18730, 32'hc32f0a4e},
  {32'h44ffa152, 32'h412b60cb, 32'hc33dd6de},
  {32'hc398cc50, 32'hc23cab96, 32'h4347e1ea},
  {32'h44bb5180, 32'hc3a24ef5, 32'h439ae3f9},
  {32'hc43c8c28, 32'h4365c7d3, 32'h437e8c39},
  {32'h44b134be, 32'h43497050, 32'h430170aa},
  {32'h445d31d9, 32'hc194e56c, 32'hc301fe91},
  {32'hc4650544, 32'hc2ea65de, 32'hc30d29d6},
  {32'h43624140, 32'hc370a27c, 32'h426885c4},
  {32'h448f52d4, 32'h4219f266, 32'hc39c1639},
  {32'hc3768088, 32'hc27d06e9, 32'h42a89f19},
  {32'h43ee3840, 32'h43a49803, 32'h4384cf24},
  {32'hc50977ba, 32'hc1dc90ac, 32'h41e693b5},
  {32'h44334027, 32'hc38413bd, 32'hc35ddc85},
  {32'hc50057c4, 32'h43610ae3, 32'h43d35457},
  {32'h45125b18, 32'h42368c88, 32'h42093610},
  {32'hc4dc9b92, 32'h41d3c916, 32'h439efd52},
  {32'h44828ed6, 32'hc312c3f9, 32'hc3841f6e},
  {32'hc4cd834e, 32'hc221fcbe, 32'h42879ed2},
  {32'h4442c51b, 32'h437c0a94, 32'h3f1c99e8},
  {32'hc470f75c, 32'hc3134558, 32'hc3592a57},
  {32'h4388d78a, 32'hc307d518, 32'h439c0d45},
  {32'hc50b02ac, 32'h43943b96, 32'hc3ace44c},
  {32'h43686f8c, 32'hc39ab712, 32'h43dd2200},
  {32'hc46974ec, 32'h4323fb8e, 32'hbe1a9480},
  {32'h444301b8, 32'h4359e181, 32'hc317ec11},
  {32'hc4ba611e, 32'h42e8612a, 32'hc3a0ec5f},
  {32'h443c32b4, 32'h4386f5ca, 32'h4126c6cd},
  {32'hc42b036c, 32'h436c8253, 32'hc3685c75},
  {32'h443d2034, 32'hc32666c2, 32'h434e22f7},
  {32'hc4e0b66c, 32'hc3990ccb, 32'h432f447a},
  {32'h448977fc, 32'h43565a91, 32'hc2e79af6},
  {32'hc2fae94d, 32'h430d8df5, 32'h43959133},
  {32'h449e9d3e, 32'hc305e3b2, 32'h432c2261},
  {32'hc50bbd86, 32'h4403cb88, 32'hc307156a},
  {32'h44e01dba, 32'hc298a99b, 32'hc1fafe47},
  {32'hc4fb12e2, 32'h4382f4a5, 32'h42fc4728},
  {32'h45166223, 32'hc294e2b2, 32'hc337033a},
  {32'hc4e5b42f, 32'h42d65083, 32'hc30575d3},
  {32'h444ce260, 32'hc27011dd, 32'h43484b54},
  {32'hc3310398, 32'h43d856ab, 32'h4376d46d},
  {32'h4452182c, 32'hc2913481, 32'hc3953fbb},
  {32'hc4c43a3a, 32'hc38040c4, 32'hc162515f},
  {32'h44853a99, 32'h4390f2e4, 32'h440dfa0c},
  {32'hc414f151, 32'hc2c292a5, 32'hc34940db},
  {32'h44e2e89d, 32'h43ab5226, 32'hc34ff63e},
  {32'hc39aba31, 32'hc39a36f3, 32'hc3033745},
  {32'h44ebaab8, 32'hc353e75b, 32'h4267eb34},
  {32'hc4ef0e71, 32'h42567471, 32'h43b863ec},
  {32'h439894dc, 32'hc32335ca, 32'h413d8427},
  {32'hc429d5ee, 32'hc15905e1, 32'h429cbde9},
  {32'h43cdb620, 32'h43c1f303, 32'hc39198c3},
  {32'hc4ba15c1, 32'hc37034d0, 32'hc256805e},
  {32'h446a9848, 32'h430c1bdf, 32'hc3c032d1},
  {32'hc469a164, 32'hc1fc3fad, 32'h434676bd},
  {32'h42452da0, 32'hc2d931e1, 32'hc3959fdd},
  {32'hc2cd12a0, 32'hc2d11c1b, 32'hc39f0d08},
  {32'h449883b4, 32'hc1aafdd3, 32'hc18019a3},
  {32'hc50d69f0, 32'hc25bb294, 32'h42b6248a},
  {32'h44c0c739, 32'h430dc85a, 32'hc29fd86b},
  {32'hc4e4fe18, 32'hc38e3ecb, 32'h444b61f3},
  {32'h448520ea, 32'hc30cf2f5, 32'h41c46a86},
  {32'hc4a174e8, 32'h4377839d, 32'h42bb8fbd},
  {32'hc49fee2c, 32'h42f796cb, 32'hc281095e},
  {32'h439670e0, 32'h427643c4, 32'hc3d9d3d5},
  {32'hc1129b00, 32'h42746efc, 32'h433e349f},
  {32'h44996f74, 32'hc20fff40, 32'hc40128b7},
  {32'hc4f24ed0, 32'hc38a026e, 32'h43ae4062},
  {32'h4400a5a3, 32'hc22d1c05, 32'hc41570cf},
  {32'hc48ecbfd, 32'hc3074040, 32'h43a4a5b3},
  {32'h45154098, 32'h418ac3bf, 32'hc383fa88},
  {32'hc3b9bf4c, 32'h438be3e5, 32'h4313b1a9},
  {32'h44cd1420, 32'hc24b6884, 32'hc23af2d6},
  {32'hc3425e56, 32'h427aa867, 32'hc30b0f5c},
  {32'h45028854, 32'h438f348c, 32'hc1b96769},
  {32'hc37cb540, 32'h43921379, 32'h4383a278},
  {32'h44ac086e, 32'h438f9b90, 32'hc39afe95},
  {32'hc3799618, 32'h43b189c1, 32'h43aae723},
  {32'h4455ee08, 32'h4363b01e, 32'h41a79fef},
  {32'hc4acd120, 32'h42b8d8ca, 32'h43002908},
  {32'h44e31d26, 32'hc233f8d3, 32'hc3104b1c},
  {32'hc4e65450, 32'hc3779222, 32'h433d1459},
  {32'h44e2001c, 32'hc39b1571, 32'hc38b09d7},
  {32'hc49fd5a7, 32'h420014ce, 32'h42b8eebc},
  {32'h450f849d, 32'hc0eb6a55, 32'h42a8a2e4},
  {32'h431f92dd, 32'hc2226323, 32'hc311d395},
  {32'h44b04d9a, 32'hc29e47b8, 32'hc2459d79},
  {32'hc42ad105, 32'hc3336d2c, 32'h43c9142b},
  {32'h44e8eb9e, 32'h42b303ef, 32'hc12c78b4},
  {32'hc4036998, 32'hc3dc579a, 32'h41d0a25a},
  {32'h44ab8968, 32'h4379e99b, 32'hc3bfc120},
  {32'hc390fcfa, 32'h42fbeeae, 32'h4031eba3},
  {32'h44975004, 32'hc3aa4ea8, 32'hc2489130},
  {32'hc3fad820, 32'hc32a30cb, 32'h42bbff13},
  {32'h44fb6467, 32'hc3386125, 32'hc2183771},
  {32'h44d05a6b, 32'h43f24f11, 32'hc3e167cf},
  {32'hc4ddc289, 32'h418f3659, 32'h43034d87},
  {32'h448fba39, 32'hc35c6440, 32'hc393d98a},
  {32'hc49dd1a5, 32'hc375b10c, 32'h42f5cbd8},
  {32'h44d3c4ea, 32'h439e1060, 32'hc369911b},
  {32'hc3d6b394, 32'h44033f95, 32'h43265cd4},
  {32'h450b93df, 32'h42d39c6b, 32'h434b1b58},
  {32'hc40ea4d6, 32'h4398640d, 32'hc3477bec},
  {32'h44ae4b22, 32'hc2e5a647, 32'h43a8610e},
  {32'hc4deaa9b, 32'h42e2b3c9, 32'hc395ee1e},
  {32'h432704ae, 32'h43981c12, 32'hc329c0a0},
  {32'hc3a0bbcc, 32'hc3b2f0fb, 32'hc297043f},
  {32'h449de4e4, 32'h43492653, 32'hc2fda1f7},
  {32'hc3e19014, 32'hc1920325, 32'h4398ba1b},
  {32'h44f6e03c, 32'h435ea25c, 32'hc272ef2e},
  {32'hc4c4354e, 32'h43477d41, 32'hc30ff04e},
  {32'h44bfac97, 32'h4391dfce, 32'h43d14a99},
  {32'h41b8db60, 32'hc3680a33, 32'hc3a5c4a0},
  {32'h44be8e2a, 32'h4338798e, 32'h42cb5bd2},
  {32'hc4bebb77, 32'hc2236fc0, 32'h43725eee},
  {32'h44b0b1b6, 32'hc30c0f45, 32'hc377d5f2},
  {32'hc3cabf7a, 32'hc2cf5747, 32'h42884465},
  {32'h44835501, 32'hc24624bc, 32'h42162864},
  {32'hc33ff596, 32'hc2a6d3c8, 32'h430a724a},
  {32'h448f3d71, 32'h4327e456, 32'hc2ef7ff9},
  {32'hc4a8503d, 32'hc2d4dc58, 32'h43e65522},
  {32'hc3294296, 32'hc2c9553e, 32'hc33ea5ff},
  {32'hc408ef3f, 32'h43728828, 32'h424e0cf6},
  {32'h448590eb, 32'hc2b658bc, 32'h437da709},
  {32'hc3ae5fba, 32'hc36a12c9, 32'h438f9148},
  {32'h4334a3d0, 32'hc29d8ad9, 32'h41b9c610},
  {32'hc42ba5ae, 32'hc3bda87e, 32'h43ed0aa3},
  {32'h44e31026, 32'h439d3ef3, 32'h42311ec0},
  {32'hc4e3f842, 32'hc36ebb6a, 32'h43263e87},
  {32'h430b132e, 32'hc38f3768, 32'hc18e4562},
  {32'hc43defbb, 32'h42b7309f, 32'hc2e09a88},
  {32'h44a3043d, 32'h43ca0ce7, 32'h43ab79d7},
  {32'hc4a6f8a2, 32'h43dfb04b, 32'h42df8e01},
  {32'h44f3b986, 32'hc2576f4d, 32'h4366d937},
  {32'hc48816fd, 32'h431eeeb2, 32'h43a9d9bc},
  {32'h44e6ce1e, 32'h42fac9b7, 32'h427b542d},
  {32'hc4ee2658, 32'h43622630, 32'hc3426e7c},
  {32'h44c33390, 32'h41f46ef0, 32'h4313230d},
  {32'hc4fb817e, 32'hc3bb447b, 32'h41e5b7fa},
  {32'h45080332, 32'h43149946, 32'hc3ac9773},
  {32'hc50411d7, 32'h420a5c07, 32'h421777a6},
  {32'h4502baa2, 32'hc19386bc, 32'h42f9526c},
  {32'hc4e40e19, 32'h4398b81f, 32'hc2b54b8a},
  {32'h4513a4d6, 32'hc391e571, 32'hc0c742d2},
  {32'hc3b61ed8, 32'hc268ee6a, 32'hc32b240d},
  {32'h4493ba62, 32'h4380b6a5, 32'hc32c42ba},
  {32'hc4d768ad, 32'hc3a5ac14, 32'h414b1a24},
  {32'h45086d2c, 32'hc312064a, 32'h4023d9d8},
  {32'hc41f491c, 32'hc28b80f2, 32'h42e614a9},
  {32'h43bd9153, 32'h434a9ccc, 32'hc31c311a},
  {32'hc4d7c028, 32'hc179a818, 32'hc3b057a9},
  {32'h450e4b3c, 32'hc335f11b, 32'h4361d096},
  {32'hc5111d62, 32'hc283bed8, 32'hc396353c},
  {32'h4520a451, 32'hc3a0ced7, 32'hc04233e9},
  {32'hc4e17418, 32'hc39b0e63, 32'hc36122fb},
  {32'h450c9a0b, 32'hc38ed98d, 32'h43170788},
  {32'hc4300010, 32'h43368809, 32'h41c32b22},
  {32'h450140ec, 32'hc3b19d43, 32'h438940ac},
  {32'hc5064078, 32'h426a3bd5, 32'h43913dd2},
  {32'h446e3e18, 32'hc285f755, 32'h4316d920},
  {32'hc31481d0, 32'h43740999, 32'hc32161af},
  {32'h448f5e54, 32'h4302f21a, 32'hc34ee002},
  {32'hc46fce7d, 32'h4401ce11, 32'hc3744cf7},
  {32'h44e11cb9, 32'h4361493a, 32'h435b2aad},
  {32'hc32502ff, 32'h42729196, 32'h429841dc},
  {32'h44a7db91, 32'h43908780, 32'hc12b59c1},
  {32'hc408479e, 32'hc293e007, 32'h4385db59},
  {32'h4519cd63, 32'hc3f1f6af, 32'h438ba6e6},
  {32'hc457940c, 32'h4202f83f, 32'hc21467ce},
  {32'h44d29d33, 32'hc41f1376, 32'hc3799a06},
  {32'hc41583d7, 32'hc28cae6a, 32'hc33d58ec},
  {32'h44ec8554, 32'hc38cc5f0, 32'h4282db99},
  {32'hc4ef0746, 32'h4372cdf6, 32'hc3733dd9},
  {32'h43e13cf9, 32'hc3273f60, 32'hc36510b8},
  {32'hc3b8e380, 32'hc3bf5e12, 32'h42229f73},
  {32'h44e37c74, 32'hc3be8e2d, 32'h42854f54},
  {32'hc40b896c, 32'hc2820996, 32'hc0dad1dd},
  {32'h4450494d, 32'hc330c9a4, 32'hc31577c3},
  {32'hc4a2b745, 32'h42ffb263, 32'hc283e385},
  {32'hc217ac58, 32'h42fc3fa2, 32'h43d7d1f3},
  {32'hc421fe33, 32'hc2b6f971, 32'hc243a296},
  {32'h445132d6, 32'h43480791, 32'hc2899aaa},
  {32'hc4a37305, 32'h41f0d580, 32'hc1f54a09},
  {32'h44c1978a, 32'hc3b4f084, 32'hc23be243},
  {32'hc4993e9c, 32'hc2ef81c9, 32'hc338216e},
  {32'hc4042d22, 32'h4344369a, 32'h43c05cc3},
  {32'h451f80e3, 32'hc28ba4f6, 32'h43c56633},
  {32'hc495d899, 32'hc1e17b73, 32'hc2e05436},
  {32'h43dbed71, 32'h43982603, 32'h436a1f2c},
  {32'hc4b7fa23, 32'h412ad1aa, 32'h438100e4},
  {32'h44cf4efb, 32'hc2fbae24, 32'hc255ed2e},
  {32'hc45e97d4, 32'hc33d43d1, 32'hc3544c6b},
  {32'hc1b46604, 32'h43904fcc, 32'hc38f1657},
  {32'hc4f725de, 32'h43d67307, 32'hc2614104},
  {32'h45110764, 32'h43021d32, 32'h42fe60ac},
  {32'hc44c7046, 32'h43da03a8, 32'hc2f80156},
  {32'h44c48df7, 32'hc3488a79, 32'h42169f79},
  {32'hc4830119, 32'hc3b11e80, 32'h431e76f6},
  {32'h45029359, 32'h42582e5d, 32'h43000503},
  {32'hc4ca1117, 32'hc38288a4, 32'h4355e17f},
  {32'h44e3969b, 32'hc32bfb1e, 32'h43aa537d},
  {32'hc4eabe7c, 32'hc30f55b4, 32'hc24f685a},
  {32'h44e974b3, 32'hc38e4b68, 32'hc33a0c59},
  {32'hc3aa55ac, 32'h427f3ed2, 32'hc2fcbdd1},
  {32'h444c8b27, 32'hc2385a23, 32'hc3854f58},
  {32'hc48aa834, 32'hc2b7c61b, 32'hc39de2f9},
  {32'h446cdb0a, 32'hc37d7195, 32'hc3844143},
  {32'hc4bda45c, 32'hc3090cdf, 32'hc3ab172c},
  {32'h44b1cce5, 32'h43db20c7, 32'h438938a5},
  {32'hc4eb75db, 32'h420e7151, 32'h42bae6c8},
  {32'h44916f28, 32'hc2c95c9d, 32'h42be1d2b},
  {32'hc3e9a434, 32'hc3433e40, 32'hc36d0910},
  {32'h4442800e, 32'hc397798d, 32'h425c0c11},
  {32'hc38d25b8, 32'hc192eb39, 32'hc3366647},
  {32'h44275268, 32'h432b51d7, 32'h4358ed32},
  {32'hc42aa946, 32'h41ed4531, 32'h42379b15},
  {32'h44c21592, 32'h42e8da59, 32'h43dbd33a},
  {32'hc4fa9741, 32'hc319da7d, 32'hc1b4344a},
  {32'h4497805d, 32'hc22d6328, 32'hc30b5c6f},
  {32'hc4821820, 32'hc34c24db, 32'h4359f377},
  {32'h440f342e, 32'hc34a6098, 32'hc2f2c3a2},
  {32'hc44adbcc, 32'hc373054f, 32'hc22648b2},
  {32'h449910bf, 32'h42cc4256, 32'h43e82348},
  {32'hc4f21a54, 32'hc4136236, 32'h4419fc65},
  {32'h445b2bc1, 32'h439d7669, 32'hc17219a4},
  {32'hc48d6b27, 32'hc37c6c5f, 32'hc20cedf6},
  {32'hc2aedc22, 32'h441de099, 32'h42a6a37b},
  {32'hc4988787, 32'h4324e87d, 32'hc2306032},
  {32'h43ee8b74, 32'h42af8f1a, 32'h43855c82},
  {32'hc4820102, 32'h42919df4, 32'h42aeccc9},
  {32'h4510ad12, 32'h43c1427f, 32'h41dc153c},
  {32'hc48e360f, 32'hc2c8d263, 32'h42a0a598},
  {32'h44b4fd6f, 32'hc32180e2, 32'h42f386c3},
  {32'hc4b75d20, 32'h42a5d656, 32'hc2a217fe},
  {32'h44cdef21, 32'h4326da58, 32'h43993212},
  {32'hc41cd934, 32'h432c1ed1, 32'hc2cbc27b},
  {32'h42e35bf8, 32'hc38accd5, 32'h439d9e12},
  {32'hc3e34dba, 32'h43be0cdc, 32'hc34c9aab},
  {32'h44d6878c, 32'h4334f31b, 32'h4322b0d4},
  {32'hc5086dcd, 32'hc3f274f8, 32'hc2ea5867},
  {32'h44a57d47, 32'h439aa5ee, 32'hc2a7da4c},
  {32'hc4b71aa1, 32'h43b0ca77, 32'h43144693},
  {32'h44d901f2, 32'hc3594628, 32'hc28c95c6},
  {32'hc4e19c44, 32'h4448bbca, 32'hc211ca03},
  {32'h44911ffc, 32'h420f98e9, 32'hc31704ad},
  {32'hc45708b6, 32'h42c554ee, 32'h43d82948},
  {32'h449f4cf9, 32'h42a4ddf4, 32'hc1b7093b},
  {32'hc4d9ba64, 32'hc21dd475, 32'h431e3e22},
  {32'hc39aecdb, 32'hc2aa51f0, 32'hc092bb91},
  {32'hc47a90ca, 32'h435a8fd5, 32'hc31e85c2},
  {32'h44a689a8, 32'hc331b37c, 32'hc2dfb4e7},
  {32'hc47d9e74, 32'h43aa82c4, 32'hc28b7a84},
  {32'h441d21cc, 32'hc23c6e0c, 32'hc33b6000},
  {32'hc28a38dc, 32'h430df0a0, 32'h43ea3a64},
  {32'h44582cca, 32'hc1e58bd5, 32'h42c08c13},
  {32'hc4ffea1b, 32'hc3b241b5, 32'hc15cfca4},
  {32'h4430ef52, 32'hc3ad836a, 32'hc2ac204d},
  {32'hc4e7db9b, 32'h433fff8b, 32'hc3479cea},
  {32'h4367f344, 32'hc35fa271, 32'hc3682221},
  {32'hc4a154bf, 32'hc2d7eef2, 32'hc33dec36},
  {32'h44a9c4b8, 32'h43303c1f, 32'hc33382b6},
  {32'hc3ba5e30, 32'hc2fdec60, 32'hc217cfd8},
  {32'h4508dd4e, 32'h43435cdb, 32'h433d4613},
  {32'hc4a43f0a, 32'hc268f674, 32'hc270e127},
  {32'h43a8ec70, 32'hc2dc0745, 32'hc3337a5a},
  {32'hc4945624, 32'h43dbe540, 32'h44041cc1},
  {32'h4509aafb, 32'hc383c4f2, 32'h4312c50e},
  {32'hc4e3bd36, 32'hc38fa0ed, 32'h42d0d00a},
  {32'h43e00d44, 32'hc3044aff, 32'h432f20ab},
  {32'hc346347c, 32'h437d074c, 32'hc36eb5d4},
  {32'h43c5d738, 32'h42b79400, 32'h42c6276a},
  {32'hc4cda743, 32'h4325323a, 32'h4350c229},
  {32'h44e757fc, 32'hc1bfe9bd, 32'hc33fdc60},
  {32'hc43bd55a, 32'hc39ef592, 32'hc2d1fa4d},
  {32'h450c4f32, 32'hc3afd922, 32'hc2ea1546},
  {32'hc48fbeb3, 32'hc2861583, 32'hc39cd81e},
  {32'h44a02028, 32'h43124e98, 32'hc2ad8122},
  {32'hc48f0724, 32'h42cdca3f, 32'hc10a61eb},
  {32'h450549d1, 32'h4339dc36, 32'h4324a64c},
  {32'hc4e126c6, 32'h43942729, 32'h42a89da3},
  {32'h44a2ea9e, 32'h431abef3, 32'hc3376ebd},
  {32'hc4bb8885, 32'h403b3990, 32'hc37eefe6},
  {32'h44b63db1, 32'h430fda78, 32'h4393f5d7},
  {32'hc3a4a638, 32'hc3ad3ae8, 32'h4354f3e8},
  {32'h43b7ddd0, 32'h40a9e9ac, 32'h43e6a4d1},
  {32'hc4b49247, 32'h43f8c6dc, 32'hc3034b23},
  {32'h44dea4ec, 32'h42890acb, 32'hc2e1270f},
  {32'hc4cf486b, 32'hc29f4c92, 32'h41a981ea},
  {32'h45073c65, 32'h43afdb99, 32'hc2552fdd},
  {32'hc5153b19, 32'h42c76dd4, 32'h3f9760b8},
  {32'h440ee731, 32'h43724bd4, 32'h42244809},
  {32'hc49ea8f3, 32'hc321ffff, 32'hc3345ef8},
  {32'h4507614e, 32'hc3bffc47, 32'h428edf8f},
  {32'hc383d86c, 32'hc2cd4525, 32'hc23f0037},
  {32'h45212b03, 32'h43afbb21, 32'h4391a04a},
  {32'hc4625b0a, 32'hc32924f6, 32'h43116aa4},
  {32'h44c81eb4, 32'hc3295cd8, 32'hc3af39b1},
  {32'hc420b860, 32'h436010fe, 32'hc2b7471e},
  {32'h44b3ac9b, 32'h41e1ee1c, 32'h435ccff2},
  {32'hc3bcad64, 32'h433bc8ec, 32'h438f7b9e},
  {32'h4487a08a, 32'hc3aa1330, 32'hc2ad7486},
  {32'h4390c4f5, 32'h42816275, 32'hc4199c84},
  {32'h443e06f9, 32'hc33a1bae, 32'hc1fb9b61},
  {32'hc489a5cd, 32'hc0ca1e3a, 32'hc2b24bbe},
  {32'h45233847, 32'hc1555ad9, 32'hc32dd437},
  {32'hc3e0bc49, 32'hc29ab4fe, 32'h4251b57b},
  {32'h44f73ff6, 32'hc1d749e0, 32'h42e100cb},
  {32'hc4488952, 32'h4277cbd6, 32'h437efee2},
  {32'h42d3f400, 32'h4304d627, 32'h43383cf8},
  {32'hc4de8157, 32'h42759c9e, 32'h432edef8},
  {32'h44d5aba7, 32'h43a5392c, 32'hc2f6352d},
  {32'hc4b0be82, 32'h43d8bac0, 32'hc34bff50},
  {32'h451c014a, 32'h432b44dd, 32'hc35cdade},
  {32'hc4f07202, 32'hc3cc5587, 32'hc20e3238},
  {32'h44d162f7, 32'h43b28ba9, 32'h43b539db},
  {32'hc43fed64, 32'hc2560bd3, 32'h432c6aed},
  {32'h44e1b92c, 32'h42692e83, 32'h43806ac2},
  {32'hc505ef5d, 32'h44022c17, 32'h42c58a17},
  {32'h44f6beaf, 32'h41f8dbf7, 32'hc382127b},
  {32'hc3439c30, 32'h43851475, 32'h4208dce8},
  {32'h440b19f5, 32'hc3be1c6e, 32'h43e05e91},
  {32'hc3f2ee78, 32'hc31280cc, 32'hc3d38a55},
  {32'h44098ced, 32'hc3ba80ad, 32'h42c124c9},
  {32'hc4eb9e69, 32'hc34e6c6c, 32'hc28664e0},
  {32'hc3855840, 32'h42e7f788, 32'h42aa97e1},
  {32'h434714d0, 32'hc18220e5, 32'h431f0f4b},
  {32'h434cbde0, 32'hc38cefc3, 32'hc339e9c7},
  {32'h42dfa060, 32'hc3b03f00, 32'hc204b4ae},
  {32'h430ef4a8, 32'h4372b1d3, 32'hc2a9ab07},
  {32'hc3b59fa5, 32'hc1f1586c, 32'hc3281ee2},
  {32'h4494395c, 32'h42444668, 32'h4162b99a},
  {32'hc4c10420, 32'hc419f2bc, 32'h43022ad1},
  {32'hc49b070c, 32'hc0ed598d, 32'h425815b7},
  {32'h44288b88, 32'hc36f0175, 32'hc39809c5},
  {32'hc4db16fb, 32'hc2b903f6, 32'hc35ddcd8},
  {32'h44ed82e8, 32'hc36d3f63, 32'hc3c87ad9},
  {32'hc4f26e6f, 32'h41749826, 32'h4353b2f0},
  {32'h44d7b47d, 32'hc3455080, 32'h43b520eb},
  {32'hc50db192, 32'h435bc9a4, 32'h3f20f8d2},
  {32'h44e96beb, 32'hc2d4a94b, 32'h4231292c},
  {32'hc506b429, 32'hc41980d0, 32'hc1cd40f7},
  {32'h44eece9c, 32'hc23bc547, 32'hc3a75928},
  {32'hc47a75f7, 32'h439d022d, 32'hc4251da6},
  {32'h44bf3d2e, 32'h43307b88, 32'h43030d4e},
  {32'hc4373004, 32'hc3a5b8fb, 32'h43b00f54},
  {32'h448169a6, 32'hc393ff9d, 32'h435e3224},
  {32'hc4bc1e23, 32'hc297f05d, 32'h42f6ca79},
  {32'h444a80c1, 32'h4362bee6, 32'hc3396ffc},
  {32'hc4da2124, 32'hc23456aa, 32'hc3b97638},
  {32'h43d5a15e, 32'hc3990d68, 32'hc296b11f},
  {32'hc340da48, 32'h44014265, 32'h43a31284},
  {32'h448714da, 32'h43872554, 32'hc268132b},
  {32'hc4c3989a, 32'h430e3ca7, 32'h430bbe9d},
  {32'h44ff495e, 32'h41d3ccf4, 32'hc3ad0603},
  {32'hc3919009, 32'h4372daee, 32'h42725890},
  {32'h43f7f5ed, 32'hc1e565a5, 32'hc1ca74fc},
  {32'hc4dcc6d0, 32'h40547f7e, 32'h438683a5},
  {32'h450e7177, 32'h4282deb3, 32'h43968558},
  {32'hc4dc6a02, 32'hc30de11e, 32'hc3181460},
  {32'h44bb74fd, 32'h424fe0f3, 32'hc3a50cc0},
  {32'hc425d519, 32'h43b7dca4, 32'hc3865327},
  {32'h44d746fd, 32'h42747a13, 32'h422c749e},
  {32'hc49d9634, 32'hc38d4fa3, 32'hc27b070b},
  {32'h44e59f11, 32'h4381028d, 32'h4302dd83},
  {32'hc4e69331, 32'h42c9a229, 32'h43904734},
  {32'h43deb856, 32'h43a07c1e, 32'hc38a155c},
  {32'hc4f6ccfb, 32'hc33132d2, 32'hc38915e1},
  {32'h4490e13e, 32'hc322cbae, 32'hc33bb3f7},
  {32'hc4037b4e, 32'hc396f368, 32'h432418a7},
  {32'h44ff1095, 32'h4022643a, 32'h42c3ff95},
  {32'hc4ab9558, 32'h42ab6f14, 32'hc3ecd81d},
  {32'h44b66c99, 32'hbd8bfc77, 32'hc39795cb},
  {32'hc38cce78, 32'h41831ca4, 32'h42c48c3e},
  {32'hc2f99b18, 32'h42c01eab, 32'h43b80436},
  {32'hc4416442, 32'h42d848ac, 32'hc3bf49b7},
  {32'h449bac4f, 32'h433eb957, 32'h43a5a2d5},
  {32'hc3f3d0b4, 32'hc2d224d7, 32'h435fc241},
  {32'h445d0229, 32'hc2852952, 32'hc2832224},
  {32'hc4a53f86, 32'hc2b1ab15, 32'h439ab135},
  {32'h433375d8, 32'hc2ddb72a, 32'h43ba2362},
  {32'hc45a32b3, 32'hc2b429d0, 32'hc3008cb4},
  {32'h44b13dfa, 32'hc3293fc1, 32'h434487fb},
  {32'hc4419dc1, 32'h434644b9, 32'h421c39ce},
  {32'h429fc640, 32'h42500bba, 32'h42945cb8},
  {32'hc4aacff3, 32'hc38c884e, 32'h42a87bd5},
  {32'h42689640, 32'h4399d1eb, 32'h4318ae5f},
  {32'hc39b64de, 32'hc346062f, 32'h430f7d00},
  {32'h44048c82, 32'hc3bd9339, 32'hc22de6e6},
  {32'hc48ccd7e, 32'hc3529fa3, 32'h423c2189},
  {32'h45042faf, 32'hc3576232, 32'h429f8f7f},
  {32'hc329cdc0, 32'h43946a25, 32'h42d60ab4},
  {32'h4346523f, 32'hc3811e22, 32'h43ae0914},
  {32'hc4640c20, 32'h414974a2, 32'h432d629e},
  {32'h4523a099, 32'h445a821d, 32'h43d1bed0},
  {32'hc4ac8a73, 32'hc3152a10, 32'h42f51ff4},
  {32'h44f72a9f, 32'h42c04de4, 32'h432ff9eb},
  {32'hc49bb1b1, 32'h434efe45, 32'hc39ad773},
  {32'h443f8d68, 32'h4237021b, 32'hc392ac2f},
  {32'hc38adbb2, 32'hc37400b5, 32'h42fe94c7},
  {32'h44bff682, 32'h44049998, 32'hc2ee4f8d},
  {32'hc4f7ef38, 32'hc31bf9d9, 32'hc3822092},
  {32'hc33bb4af, 32'hc2a45e39, 32'h42ef2a5e},
  {32'hc4fae14d, 32'h41dfed58, 32'h430020dd},
  {32'h448f71d2, 32'h43698116, 32'h41b35103},
  {32'hc442cad6, 32'hc33471e0, 32'h43407a62},
  {32'h419bce00, 32'h42f19308, 32'h433bc5ed},
  {32'hc3a455ef, 32'h42159567, 32'h407797f5},
  {32'h4507167e, 32'hc18fb167, 32'h43b7cb34},
  {32'hc411aea0, 32'h42cc68b2, 32'hc3c6c840},
  {32'h44ece66b, 32'h431aa54b, 32'hc2bcf295},
  {32'hc3a43511, 32'hc37194a9, 32'h4302f739},
  {32'h446bbe46, 32'h431e5c4a, 32'hc33ea53f},
  {32'hc488b716, 32'h4317da78, 32'h42c7da8a},
  {32'h44fca456, 32'hc32085c7, 32'hc36c8b9a},
  {32'hc4a5b0b2, 32'h442a9429, 32'hc174e848},
  {32'h4491a29b, 32'hc34b31a1, 32'h438b656a},
  {32'hc4ba268a, 32'hc393df88, 32'h434f8795},
  {32'h44d49c9d, 32'h439e2308, 32'h433ef555},
  {32'hc4ec1ab3, 32'hc3002a94, 32'hbf761e00},
  {32'h445bbd1d, 32'hc2f05062, 32'hc32545d6},
  {32'hc4556760, 32'h4265513f, 32'hc2bfe0c7},
  {32'hc485a35b, 32'h427b6985, 32'h42bcad8c},
  {32'h45042cd1, 32'hc2db0ab1, 32'h423e1a0b},
  {32'hc513d334, 32'hc2b58188, 32'hc2f8a7d2},
  {32'h43e10aa8, 32'h43600401, 32'h43da99fb},
  {32'h41afb380, 32'hc2056790, 32'h43491d3a},
  {32'h44911deb, 32'h4298fd73, 32'h42c81df8},
  {32'hc496f3b8, 32'h42e6dd48, 32'hc296c9f3},
  {32'h44884ae1, 32'hc2623fe3, 32'h431c58e8},
  {32'hc4eb8faa, 32'hc28d259b, 32'h43956465},
  {32'h442a9440, 32'h43043f97, 32'hc38cb604},
  {32'hc23df954, 32'h433e0a7f, 32'h42d803f4},
  {32'h44aa3732, 32'hc2a41839, 32'h4368d80d},
  {32'hc47d95ff, 32'hc34a2714, 32'hc3b95342},
  {32'hc25c3980, 32'hc3bcedc9, 32'hc1b24c1f},
  {32'hc50b3aa9, 32'hc281eccb, 32'hc2d4c766},
  {32'h449ed480, 32'h42b19a15, 32'hc2534e15},
  {32'hc4f5e11f, 32'hc2a1387c, 32'hc28a88bf},
  {32'h4518a1ee, 32'h43467800, 32'hc2d3a345},
  {32'hc3055f0d, 32'h44836f0f, 32'h435fa676},
  {32'h45042904, 32'hc3115cd2, 32'hc1410bdb},
  {32'hc46e4bd4, 32'h4315d0a4, 32'hc3ba6801},
  {32'hc5187746, 32'hc3982ca9, 32'h42db97e5},
  {32'h44d27e07, 32'h433d75d3, 32'hc1b07da1},
  {32'hc4fb0da7, 32'h41c757da, 32'hc337de86},
  {32'h44cc0afc, 32'h41d6b56f, 32'h4348d720},
  {32'hc38898bf, 32'h4263cca1, 32'h429cf1fa},
  {32'h443474ff, 32'h43b3b0aa, 32'hc28cdab0},
  {32'hc493986a, 32'h44028425, 32'h4257ef0e},
  {32'h437f0fa8, 32'hc2bf56b0, 32'hc34799c1},
  {32'hc482e9bf, 32'hc3c653c7, 32'hc296ea9b},
  {32'h44a572d0, 32'hc295dc2a, 32'hc2327879},
  {32'hc4baca04, 32'h426200c8, 32'hc2a22eab},
  {32'h442bc5ec, 32'h428daf48, 32'hc23c4fd4},
  {32'hc3f31cf0, 32'hc234bfa8, 32'hc283cbc6},
  {32'h44b359bc, 32'hc2d51eeb, 32'hc314a90e},
  {32'hc4f1b1a6, 32'h43b0c5f8, 32'hc35f44e7},
  {32'h44aff82a, 32'hc3253701, 32'hc21a1096},
  {32'hc4c64a9f, 32'h43361a88, 32'h4375a7a5},
  {32'h4460a0cb, 32'h43220ea3, 32'h431a3d96},
  {32'hc414f370, 32'h42d0506a, 32'hc2ee6c97},
  {32'h452a72af, 32'h43a320e4, 32'h4334a716},
  {32'hc4cbf5f5, 32'hc367089e, 32'hc3978ca5},
  {32'h44e8c42a, 32'hc31797a7, 32'hc2e9d50a},
  {32'hc4a1faf6, 32'hc38a62ff, 32'h4392c238},
  {32'h44db4fbd, 32'h43b1dbdd, 32'hc31701b3},
  {32'hc45ba0d6, 32'hc20224ca, 32'hc2c9e455},
  {32'h44e5b3df, 32'h4261302c, 32'h42dbbce9},
  {32'hc3d46561, 32'hc321257a, 32'h43d44ecd},
  {32'h4341fc18, 32'h42d90b76, 32'h425c0e8f},
  {32'hc3929aac, 32'h43ad36d6, 32'h430beeed},
  {32'h442ae8c4, 32'h439d0185, 32'hc31cf08c},
  {32'hc528ff0a, 32'hc2b09842, 32'hc258d6ea},
  {32'hc4cc344a, 32'h437cb8a8, 32'hc2756341},
  {32'h450eb386, 32'hc3b5aa4b, 32'h41f376b2},
  {32'hc501509f, 32'hc2ca55cb, 32'hc34f53d4},
  {32'h443bd21b, 32'hc3525068, 32'h43013316},
  {32'hc47072d0, 32'h434e4bda, 32'h43232f61},
  {32'h451058fe, 32'hc1adff4b, 32'h41a83f00},
  {32'hc4a70020, 32'h43ba18ac, 32'h42d7a9f0},
  {32'h43d7738c, 32'hc3bdef30, 32'h4271707b},
  {32'hc43a1b09, 32'hc3206250, 32'hc18595e2},
  {32'h43143630, 32'h433faf42, 32'h4389b11d},
  {32'hc4f4ce67, 32'hc24c414a, 32'h43567252},
  {32'h4461c564, 32'h421673be, 32'h416bd10e},
  {32'hc4994de6, 32'hc39c427a, 32'hc384e1a1},
  {32'h447d6c16, 32'hc2afa294, 32'h43a35991},
  {32'hc480ccd5, 32'h437c07c6, 32'h41d11ef1},
  {32'h44de4882, 32'hc329bc3e, 32'hc300203c},
  {32'hc3bb5bfa, 32'h439f4e09, 32'h4249b7f2},
  {32'h44c4e48c, 32'h4377a9e0, 32'h4304e285},
  {32'hc310324a, 32'h43e267ed, 32'hc3292ddc},
  {32'h43a86c9a, 32'hc2820ecd, 32'h433a8c3a},
  {32'hc45cbbe2, 32'h42abad71, 32'hc20e347b},
  {32'h447eab42, 32'h4277fc96, 32'hbf2e837a},
  {32'hc3a828d0, 32'h433132c9, 32'hc3d9dc0d},
  {32'h4480e04a, 32'h439c9ba4, 32'h43a1123d},
  {32'hc462adfa, 32'hc31f6486, 32'h428a479b},
  {32'h44e33a81, 32'hc3a6e1aa, 32'h42b3262a},
  {32'hc505a98a, 32'hc2b14c3a, 32'h434523b1},
  {32'h446e68bc, 32'hc2693e26, 32'h4183a3be},
  {32'hc4196d5e, 32'hc0b0580e, 32'hc1f21101},
  {32'h450fbe77, 32'h42e3c34c, 32'hc2887a81},
  {32'hc4dfe424, 32'hc1f45dc4, 32'h42a691c8},
  {32'h44ee2f13, 32'hc2caa451, 32'hc30b0b94},
  {32'hc5166982, 32'h430ba86f, 32'h4336d859},
  {32'h43574cf0, 32'h439330bd, 32'h43646f9d},
  {32'h429b7780, 32'hc19f0b86, 32'hc3518dfa},
  {32'h44fe8fb5, 32'hc32991f6, 32'hc35ecc79},
  {32'hc442e852, 32'h434aa58e, 32'hc3dc8692},
  {32'h44aef2dc, 32'hc3feaeae, 32'h4327f139},
  {32'hc4c8532d, 32'h435648c7, 32'hc3474b6f},
  {32'h443a9880, 32'hc1dd6216, 32'h4095aff5},
  {32'hc490318a, 32'h431eb0a1, 32'hc3ed8ba1},
  {32'h44e2f60e, 32'h438ec4d5, 32'hc1ad5112},
  {32'h436a2d80, 32'hc2d464f2, 32'h411ccdfc},
  {32'h44b05ef3, 32'hc29b2ded, 32'h432be16c},
  {32'hc4980606, 32'h42dbe614, 32'h430d3527},
  {32'h44fa2de3, 32'h428015b2, 32'hc1a63220},
  {32'hc2a79ec0, 32'hc3766b5d, 32'hc2c0e237},
  {32'hc50c2a6a, 32'hc1697988, 32'h424105ef},
  {32'hc4804726, 32'h43879f43, 32'hc39b4d84},
  {32'h448dd3d6, 32'hc3f07563, 32'h43e30a85},
  {32'hc48318ac, 32'h43ae31bd, 32'hc229dfe0},
  {32'h44a2a931, 32'h43ba638c, 32'h4151b67b},
  {32'h43237c9c, 32'h41336b6f, 32'h42559ab0},
  {32'h43c70a1c, 32'h43907dfc, 32'h436e64e0},
  {32'hc4a66c2c, 32'h430f2562, 32'hc3a937e3},
  {32'h44e62cc2, 32'hc39a86f8, 32'h4350ced0},
  {32'hc4c408e1, 32'hc2e1afee, 32'hc32fafc1},
  {32'h44694f6a, 32'h4408f8cd, 32'h433a9dcd},
  {32'hc5070bb9, 32'h4378575b, 32'h429c333c},
  {32'h4234c280, 32'hc3566863, 32'h42b519ca},
  {32'hc4aee017, 32'h4292b6bf, 32'hc289a58e},
  {32'h44d78579, 32'hc2d7782b, 32'h43c71a8f},
  {32'hc4fe1515, 32'h4364d0b0, 32'hc3927466},
  {32'h438a5c80, 32'hc3ca5db1, 32'h43967567},
  {32'hc49e6a55, 32'h42215abf, 32'h42fda92f},
  {32'h448b95ad, 32'hc3981bc6, 32'h42ffcc85},
  {32'hc3c4b22c, 32'hc1badac4, 32'hc2fee593},
  {32'hc4714c02, 32'h43ba1025, 32'hc37ee538},
  {32'h4406df59, 32'hc3017636, 32'hc3089c7b},
  {32'hc397a731, 32'h41e62365, 32'hc3807c82},
  {32'h44092405, 32'h42a539c2, 32'h43a5a09f},
  {32'hc501be39, 32'hc36647f3, 32'hc24c7e07},
  {32'h45081917, 32'h43a2adb7, 32'h4384c0a8},
  {32'hc50a7d40, 32'h43d052c0, 32'hc34ad03f},
  {32'h451d3b19, 32'hc358faa8, 32'hc302c92d},
  {32'hc455a27a, 32'h421a7f22, 32'hc40835cb},
  {32'hc39c2a36, 32'hc30c2c8e, 32'h41b5227e},
  {32'h45083851, 32'h4308a12e, 32'h43a717c7},
  {32'hc4a8179c, 32'hc2fb7baf, 32'hc2e46e30},
  {32'h44a686e4, 32'hc29b0998, 32'h41a0f1c0},
  {32'hc4cc2845, 32'h4397a542, 32'h43b4b351},
  {32'h44b5c730, 32'hc2a4b9de, 32'h4390d5c4},
  {32'hc3bb74fa, 32'h423a1925, 32'hc12ce2ff},
  {32'h41b23a40, 32'hc418f3f8, 32'hc252051e},
  {32'hc4c4ad93, 32'h425bb456, 32'h44016c5d},
  {32'hc22fea80, 32'h4212f9e6, 32'hc2f3eac8},
  {32'hc48d20db, 32'h440de4cb, 32'h434f6d77},
  {32'hc1eb7b80, 32'h433aa5b5, 32'hc303c192},
  {32'h439dcc10, 32'h43366d72, 32'hc2d94f8c},
  {32'h4508fdf9, 32'hc383e622, 32'h424d1c83},
  {32'hc48c4c06, 32'hc30139d2, 32'h4292203a},
  {32'h430d6a78, 32'h43e380ac, 32'h43185ab2},
  {32'hc2a74540, 32'hc23ec510, 32'h42d0746a},
  {32'h431cbf2c, 32'hc391ae87, 32'h42caf59a},
  {32'hc4edff62, 32'hc2a0e403, 32'h41bb37ae},
  {32'h44af9642, 32'h43c1b2dd, 32'h42ac88cd},
  {32'hc3f7ea68, 32'hc330b53c, 32'hc39012da},
  {32'h44987440, 32'hc1524873, 32'hc326a780},
  {32'hc4f56713, 32'hc27629c7, 32'hc3ae1f46},
  {32'h44ad89c6, 32'h43b24000, 32'h42f1746c},
  {32'hc48a7855, 32'h440f5806, 32'hc38dfa8f},
  {32'h445e8744, 32'h3f745240, 32'hc35f5041},
  {32'hc37c3228, 32'h43a226e0, 32'h41c6fb31},
  {32'h43c7aa78, 32'hc36e5c8f, 32'h43b9c1fa},
  {32'hc5218fe5, 32'h436084e2, 32'hc39944fc},
  {32'h432bb189, 32'h43886a7b, 32'hc378b022},
  {32'h41d35f00, 32'h434dc074, 32'h42f9d870},
  {32'h4446cf5a, 32'hc3404a58, 32'hc31e54e6},
  {32'hc49e201e, 32'hc1edbd98, 32'hc38171ec},
  {32'h4515e8d2, 32'hc2a41474, 32'h42bad660},
  {32'hc4ef95ec, 32'h431544b6, 32'h4335561c},
  {32'h4512847f, 32'h43f32cc8, 32'h43852c38},
  {32'hc422938e, 32'h42742590, 32'h418946a4},
  {32'h43c40c68, 32'hc346579b, 32'h4262a0b1},
  {32'hc4b4191c, 32'h422e7fb3, 32'h4418718f},
  {32'h41b2f6f0, 32'h43846c1f, 32'h41428749},
  {32'hc4fda328, 32'h43c22085, 32'hc1d4466d},
  {32'h43603e97, 32'hc369f553, 32'h430497bb},
  {32'h435effe0, 32'hc37c7770, 32'hc21aa89b},
  {32'h45098ca6, 32'hc2179e84, 32'hc362e0c2},
  {32'hc3776437, 32'hc1b1ca8d, 32'h43535d5e},
  {32'h44a28011, 32'h43b42ff4, 32'h435898db},
  {32'hc3c920dd, 32'hc29028fe, 32'hc31fee61},
  {32'h44a5eb69, 32'hc2a05801, 32'h4316ba3a},
  {32'hc3d55ac8, 32'h438e9e07, 32'h431bca7a},
  {32'h43e1df20, 32'hc31b1a9a, 32'h43db9760},
  {32'hc49624cb, 32'hc1a741b4, 32'h42f44cfa},
  {32'h43917dca, 32'h4220556a, 32'hc32dc65e},
  {32'h4428bdb6, 32'hc26a2ee5, 32'hc3c2bbf5},
  {32'hc4cad292, 32'hc203e056, 32'hc125e0aa},
  {32'h44c8f84b, 32'hc3be6066, 32'hc2abc1a7},
  {32'hc4fd1c46, 32'hc2e2aa84, 32'hc27f4aa8},
  {32'h44f2c9ca, 32'h42ede9a0, 32'hc2d6299c},
  {32'hc4cdd7c3, 32'h4329256f, 32'hc2abac46},
  {32'h449396fd, 32'hc2eb9bfb, 32'h42511df8},
  {32'h4319bb10, 32'hc1b99d09, 32'hc2526702},
  {32'h44d59e0c, 32'h4321d0da, 32'h42972c9f},
  {32'hc524d823, 32'hc1d53a5b, 32'h4326eeed},
  {32'h439af4bc, 32'h43d97d0b, 32'h43e42c9c},
  {32'hc4e9996e, 32'hc2fb7f3f, 32'hc1398a63},
  {32'h45000fbb, 32'hc2430ad6, 32'hc2c54fd9},
  {32'h42f741bd, 32'h42a0feb4, 32'h43985e62},
  {32'h4505ce14, 32'hc323cf1d, 32'h42dce320},
  {32'hc466f164, 32'h438c73a3, 32'h4285d946},
  {32'h44ada676, 32'h42f3baa5, 32'hc16fd09b},
  {32'hc5016760, 32'hc2ae804a, 32'h4388c88a},
  {32'h44bb1c4e, 32'h43db9aea, 32'h42585d51},
  {32'hc4b8ae86, 32'hc3c98e13, 32'h41229f1c},
  {32'h44280583, 32'h4309ffc8, 32'h431e8dd2},
  {32'hc448f3a0, 32'h44030082, 32'h4343e969},
  {32'h4483e838, 32'h413c1bf1, 32'h4327cc97},
  {32'hc3528348, 32'hc354a358, 32'hc2489218},
  {32'hc4e404c7, 32'hc1e16eda, 32'h428b7141},
  {32'h44cd037f, 32'h4359271e, 32'hc3a20a38},
  {32'hc50293ad, 32'h423d810b, 32'h42308861},
  {32'h4519efff, 32'h4322926c, 32'h43cfda5e},
  {32'hc48ce7aa, 32'hc37bada0, 32'hc2e0c29b},
  {32'h438398a0, 32'h42503dfb, 32'h43bc675b},
  {32'hc47ec0c5, 32'h43d1ebf1, 32'h431616ca},
  {32'h44cf6915, 32'hc30b3aa5, 32'hc3f3e02f},
  {32'hc3da5416, 32'h43790662, 32'hc37f61a3},
  {32'h4395b562, 32'h426131ca, 32'hc33f00fa},
  {32'hc4a68b35, 32'hc380ca6f, 32'hc1d4bd4b},
  {32'h4396cf3e, 32'h43422bec, 32'h43f04bdb},
  {32'hc4d24056, 32'hc2b5bc9e, 32'h430c8bec},
  {32'h4455a28f, 32'h42fefc36, 32'hc277b687},
  {32'hc4004bb9, 32'hc3039167, 32'h430f22b5},
  {32'h44c1e138, 32'hc39003d2, 32'h42a66cf7},
  {32'hc446636c, 32'hc313563b, 32'h427a5334},
  {32'h43ce5dda, 32'hc300927d, 32'h44063790},
  {32'hc4fef686, 32'hc1850801, 32'hc32309da},
  {32'h44fb6160, 32'hc2455560, 32'hc375a36d},
  {32'hc503c7df, 32'h419f4582, 32'hc1cd31b0},
  {32'h44dc7790, 32'h437b7f81, 32'hc204227b},
  {32'hc38d83a8, 32'h4321965e, 32'h4344c8a1},
  {32'h450289c8, 32'hc2cbc95d, 32'hc1d2d88a},
  {32'hc4903b21, 32'hc2f3831c, 32'h43775650},
  {32'h43949588, 32'hc37cf346, 32'hc3839c20},
  {32'hc4fb74ec, 32'hc3a32d68, 32'h43d80c17},
  {32'h44d8ab55, 32'h41972f65, 32'hc250e3a7},
  {32'hc466942d, 32'hc376416b, 32'h43455245},
  {32'h45152d6f, 32'hc2f8f681, 32'h4293a29a},
  {32'h432fe04b, 32'hc2be3657, 32'h42384ea2},
  {32'h449c9cae, 32'hc231787a, 32'h434a1ceb},
  {32'hc49e03ae, 32'h412d266c, 32'h4351bffb},
  {32'h43a19aab, 32'hc39168b7, 32'hc317cb68},
  {32'hc34ec508, 32'h42e69244, 32'hc2cec9d0},
  {32'h44ddace6, 32'h42a58304, 32'hc3994f4b},
  {32'hc4f116f4, 32'hc19ae602, 32'h42a3f93b},
  {32'h4461a5e1, 32'h432720e0, 32'hc34e51b9},
  {32'hc4c4198c, 32'h42b98efc, 32'hc26611b2},
  {32'h451af924, 32'hc35c0446, 32'h43d3b0ef},
  {32'hc439cd6e, 32'h443afba5, 32'hc3332e5d},
  {32'h43ff1470, 32'hc2675853, 32'hc30c54b7},
  {32'hc4cae393, 32'h417b8743, 32'h43322295},
  {32'h43e43172, 32'hc2a8a695, 32'hc3c93bde},
  {32'hc401198c, 32'h43871ad2, 32'h4301d4d7},
  {32'h4474b900, 32'h426f2c77, 32'h43c75b44},
  {32'hc4ef9ba0, 32'h4382e34b, 32'h433725f5},
  {32'h44e9b2c5, 32'hc30b6c77, 32'hc3979156},
  {32'hc3dbfadb, 32'h43975f02, 32'h436abb78},
  {32'h44813058, 32'hc389698d, 32'h4200564a},
  {32'hc501b0d6, 32'hc2fdfcc3, 32'h43563ad9},
  {32'h43e2adfe, 32'h42881a59, 32'h428b5548},
  {32'hc4b19b9f, 32'hc28d0e67, 32'hc433ea21},
  {32'h4468d2e4, 32'h43a3bd49, 32'h42ab8811},
  {32'hc49502b9, 32'h42c7c015, 32'hc22b070e},
  {32'h4462f605, 32'h4385261c, 32'hc2b2b926},
  {32'h42eaeab6, 32'hc2243dc6, 32'h40722957},
  {32'h44544a50, 32'h430edc8a, 32'hc2e610b2},
  {32'hc4bf3cb0, 32'hc2e1ea14, 32'hc2bad715},
  {32'h44ac4a8a, 32'hbe51cb80, 32'h4287a561},
  {32'hc436227c, 32'h43736022, 32'h4310cd7d},
  {32'hc3266940, 32'hc32bef81, 32'h425a76c7},
  {32'hc4f6d734, 32'hc3d2db5e, 32'h43bc0454},
  {32'h44e0e259, 32'h441584f9, 32'h438676b2},
  {32'hc34f8c30, 32'h42da1136, 32'hc40e9467},
  {32'h4472b4b6, 32'hc337167f, 32'hc3ac8c92},
  {32'hc4db90bc, 32'hc2fb2876, 32'hc391db14},
  {32'h4456f611, 32'hc355607a, 32'hc1aa8a44},
  {32'hc385a246, 32'h42d5eb63, 32'hc3163be8},
  {32'hc3213110, 32'hc3d5af82, 32'h430bdf94},
  {32'hc4a58d67, 32'h434a4bfe, 32'hc3a0d142},
  {32'h43744990, 32'hc39d14cd, 32'h422e26e4},
  {32'hc4f1e144, 32'h43492c68, 32'h42df657a},
  {32'h43b3375c, 32'h41f50a9b, 32'h41ea45a3},
  {32'hc3b493bc, 32'hc395c983, 32'h43653f38},
  {32'h4407f689, 32'h4212afb0, 32'h4388e031},
  {32'hc49e0063, 32'hc337ca90, 32'h4134dc5d},
  {32'h4500175a, 32'h4351c899, 32'hc28c71c9},
  {32'hc4bb4bba, 32'h43303b41, 32'h43f7b522},
  {32'h44b7a8e3, 32'hc1b04e48, 32'h43964c56},
  {32'hc503717a, 32'hc430e194, 32'hc1d16f66},
  {32'hc3e25890, 32'h4358f499, 32'hc35a22fb},
  {32'hc4baf27b, 32'hc17b6cb4, 32'hc3490f90},
  {32'h44e25bc1, 32'hc3241ab3, 32'h43b3914c},
  {32'hc447abd3, 32'h4300e86c, 32'hc2bf9f76},
  {32'h449ccf42, 32'hc2b96841, 32'h4396d184},
  {32'hc43fd94c, 32'hc2aa79ee, 32'hc391fcb8},
  {32'h441e40ae, 32'hc3b395e6, 32'hc31dc367},
  {32'hc517293c, 32'hc4254d05, 32'h43626fd6},
  {32'h44b83e62, 32'hc3556c3f, 32'h43495102},
  {32'hc3eb6d7f, 32'hc3d2e4db, 32'h4338f9d2},
  {32'h4407d742, 32'hc3d7b78c, 32'h43a8d96d},
  {32'hc4fec886, 32'hc0d0e06a, 32'h43703d25},
  {32'h44e5958e, 32'h43d37d42, 32'hc39349a5},
  {32'hc4f15604, 32'h43c841b1, 32'hc3b2b06c},
  {32'h43957da4, 32'hc3683b96, 32'hc332ab56},
  {32'hc38cd795, 32'h43609e8d, 32'h426bb497},
  {32'h43e53c7c, 32'h43a96edf, 32'hc369dd43},
  {32'hc502edb0, 32'hc3132626, 32'h435937f9},
  {32'h450d1422, 32'h43b232d7, 32'hc17bad5d},
  {32'hc4a09d49, 32'hc3248288, 32'hc2b2de48},
  {32'h448ee328, 32'h4318ac4e, 32'h413026ea},
  {32'hc4a923a9, 32'hc2d98358, 32'hc153d444},
  {32'h4496ba49, 32'hc3657908, 32'hc3664636},
  {32'hc501a959, 32'h439b0148, 32'h4376c600},
  {32'h439201e8, 32'hc2d2480f, 32'h41af16e1},
  {32'hc476191a, 32'h436c94d4, 32'h4327ff5f},
  {32'h439890e4, 32'hc36de05e, 32'h43122191},
  {32'hc494ba57, 32'hc3779ab2, 32'hc205fdc8},
  {32'h44c0c1d0, 32'hc3417e90, 32'hc3c99e23},
  {32'hc50811be, 32'hc2bea0f8, 32'h43ac5c8f},
  {32'h44b3e471, 32'h43a0e6db, 32'h42fba4a8},
  {32'hc4e7838c, 32'hc41c96d8, 32'h4300425a},
  {32'h4501402c, 32'h437da2f5, 32'h42ceec2a},
  {32'hc481033d, 32'h43651d8b, 32'h438700cf},
  {32'h44a33a36, 32'hc181db4e, 32'hc30cde6c},
  {32'hc4fec709, 32'h42a10743, 32'h4213fa84},
  {32'h4511b1b1, 32'h43c24af2, 32'h429974c8},
  {32'hc5080de1, 32'h43e36b86, 32'h43c52a93},
  {32'h4297aeaa, 32'hc3554b67, 32'h43aa9ed0},
  {32'hc46957fc, 32'h42cd9bc2, 32'h431c8763},
  {32'h444b7cbd, 32'h43483111, 32'hc320b063},
  {32'hc452376c, 32'h42adc6cb, 32'hc25162b4},
  {32'h429a1ac0, 32'hc31b3ecd, 32'hc3ea7ef1},
  {32'hc3c65870, 32'hc29282fc, 32'h43e4f2d1},
  {32'h44ba36dc, 32'hc392565e, 32'h426b8fd7},
  {32'hc4ef5db0, 32'hc2976a66, 32'h434fc472},
  {32'h43805d78, 32'h42562946, 32'h421b2bc6},
  {32'hc30bddba, 32'hc34a7264, 32'h42fb3163},
  {32'h44ef9edc, 32'hc38daa28, 32'hc2bce550},
  {32'hc48ca5ab, 32'hc36d2229, 32'hc381c4f2},
  {32'h43ddd834, 32'hc3ac2918, 32'hc28fe55a},
  {32'hc4e1b4fa, 32'h418448a7, 32'hc387652f},
  {32'h44fece84, 32'h42667161, 32'h43b65c07},
  {32'hc50e4551, 32'h42136bc0, 32'h4333b934},
  {32'h432fc3e0, 32'h43a4e30a, 32'h4283c584},
  {32'hc4af7526, 32'h43f61cb4, 32'h42a2363d},
  {32'h43c1c428, 32'h41d7ca44, 32'hc38b5983},
  {32'hc49ae056, 32'h43859388, 32'h43543dc4},
  {32'h44ac3e56, 32'hc3d1de49, 32'hc1a2acd5},
  {32'hc50e28f8, 32'hc2a89d2b, 32'hc2b07fc5},
  {32'h43cd2cd7, 32'hc3d75164, 32'h41ee4ea8},
  {32'hc3ed96e0, 32'h424280b7, 32'hc18f5391},
  {32'h443c83ee, 32'h430def31, 32'h4260dfab},
  {32'hc50877a0, 32'h42401c98, 32'h429d362d},
  {32'h44617592, 32'hc3b4c3cc, 32'h433a4dce},
  {32'hc4b80f53, 32'h43486911, 32'hc34986fc},
  {32'hc2e17ac0, 32'h42c81c39, 32'hc37877ac},
  {32'hc457b904, 32'h4379da17, 32'h431fb6df},
  {32'h44ec509b, 32'hc2e8d450, 32'h43184aaf},
  {32'hc502dd47, 32'h41bb148d, 32'hc2873dba},
  {32'h429247a0, 32'h42a82258, 32'h434093a1},
  {32'hc50d60b8, 32'hc31cfc07, 32'h439730f9},
  {32'h44f364f2, 32'hc1f69086, 32'h42a19643},
  {32'hc4a62de0, 32'h43ba4864, 32'hc33069ae},
  {32'h43ec2da0, 32'h433894a2, 32'h40ae7350},
  {32'hc4ac7c5c, 32'hc3cba66c, 32'h43a7ec0e},
  {32'h45121a0f, 32'hc30489dd, 32'hc254f9a2},
  {32'hc4d01f9c, 32'h43123a4c, 32'h43551f7e},
  {32'h44b3a64a, 32'h43d6ccda, 32'hc3b0d28a},
  {32'hc3892e30, 32'h42f5d8ff, 32'hc386a02b},
  {32'h4464adf0, 32'h4357c588, 32'hc1f12c04},
  {32'hc43ac2e9, 32'h42b995fe, 32'hc1d40cad},
  {32'h44ec46b2, 32'hc40bf39c, 32'hc39ee099},
  {32'hc4de7f4a, 32'hc209cfe1, 32'hc197390a},
  {32'h43b395b8, 32'hc3089f33, 32'hc3029a78},
  {32'hc4a5f174, 32'hc35b64c0, 32'hc301ebed},
  {32'h44b04721, 32'hc2b443c8, 32'hc3c6f1ee},
  {32'hc48226a2, 32'hc2b44ac5, 32'hc2d8ae5c},
  {32'h44a41d96, 32'h41a78da4, 32'h439a88b3},
  {32'hc4684766, 32'hc206e5bd, 32'h4381ec8f},
  {32'h44df0580, 32'h42c99df1, 32'hc3832aae},
  {32'hc4cad0cb, 32'hc0ba2ca8, 32'h42dc2272},
  {32'h446cf184, 32'hc28a39b7, 32'h4230834c},
  {32'hc3efebe3, 32'h4302e008, 32'h428a26bf},
  {32'h449430ea, 32'hc34712c4, 32'h4237dde0},
  {32'hc4545d16, 32'h4384ac3a, 32'h437709f4},
  {32'h44b20006, 32'h424d25df, 32'h4313902f},
  {32'hc4c26284, 32'h42b0ca94, 32'hbe8b2a60},
  {32'h43be432c, 32'hc1369eb0, 32'h41e893c1},
  {32'hc40699ae, 32'h424e0ac6, 32'hc329d2aa},
  {32'h44846a8d, 32'h43c8d5fc, 32'h42c164d5},
  {32'hc325915e, 32'h4304ebc6, 32'hc3cdf28b},
  {32'h41fd2e18, 32'hc3d4a4ea, 32'h4339d1fa},
  {32'hc1a1b280, 32'hc3108382, 32'h43a5358d},
  {32'h4504bd84, 32'hc392c3d8, 32'h435d4858},
  {32'h42e41b6a, 32'hc2f5fc48, 32'hc3bef28f},
  {32'h44f0cadf, 32'h4327c5f8, 32'h430b9f0f},
  {32'hc324a1c0, 32'hc3802c5f, 32'h426036cc},
  {32'h4472fa7d, 32'h42d4c94a, 32'h432b9f7f},
  {32'hc3a6f563, 32'hc23092ac, 32'h43a1d1a9},
  {32'h44dc4d6c, 32'hc21e3b81, 32'h4107b3ea},
  {32'h413bafd8, 32'hc34b0943, 32'h42c8a723},
  {32'h44e7bdc0, 32'h42995f26, 32'h436c8904},
  {32'hc4c8356a, 32'h44136eca, 32'h43de5172},
  {32'h452328e7, 32'h433878c3, 32'hc327081c},
  {32'hc3306c76, 32'hc3902200, 32'h42901e8c},
  {32'h438ed484, 32'hc31f7d39, 32'h42bd8a61},
  {32'hc4e69632, 32'hc34ec0e6, 32'hc3aeca9a},
  {32'h43b5e5a8, 32'h440ea0d7, 32'hc337599f},
  {32'hc504dfdf, 32'h3fb45b90, 32'h438a965d},
  {32'h4507cfd2, 32'h424af127, 32'h437eb475},
  {32'hc341d8a0, 32'hc13a7f80, 32'hc29e4050},
  {32'hc43864b4, 32'hc36d2c1c, 32'h42b76fe5},
  {32'h445a4848, 32'h422eecfc, 32'h43bb0ca2},
  {32'hc420c4e0, 32'h4354c55b, 32'hc2fb2472},
  {32'h44a649fc, 32'h4329423c, 32'hc216ad8f},
  {32'hc4e7fa7b, 32'h42f098af, 32'hc2f70226},
  {32'h441893d4, 32'h4315f134, 32'h42a4cf79},
  {32'hc48f40ef, 32'hc32785b2, 32'h43b8ce1d},
  {32'h43ccddac, 32'hc2f9081a, 32'hc395fbc1},
  {32'hc4d024e1, 32'h430e29d0, 32'hc4077ee0},
  {32'h4360e3a0, 32'hc390ed48, 32'h42b40063},
  {32'hc21dbc6a, 32'hc3f46e48, 32'hc32cad98},
  {32'h43aeb480, 32'hc3925488, 32'h437111ff},
  {32'hc50c5c4c, 32'hc21facc9, 32'h438b99c2},
  {32'h44325e3e, 32'hc3955bf0, 32'hc21cecff},
  {32'hc5118559, 32'hc3d74078, 32'h4388d736},
  {32'h44b8798f, 32'hc322b0e1, 32'h44059bf3},
  {32'hc43a6833, 32'h429e71fe, 32'hc33d82cb},
  {32'h41859ebc, 32'hc2dc85b7, 32'h43b65ca4},
  {32'hc4791edc, 32'hc2992e80, 32'h43962a86},
  {32'h43f6c12c, 32'h42880165, 32'h41d538f2},
  {32'hc4c75a12, 32'h43ebf9c1, 32'hc35b338c},
  {32'hc4ea3c41, 32'hc2de1fee, 32'hc2939091},
  {32'h42c147da, 32'hc23dd3e9, 32'hc314745d},
  {32'h40395400, 32'h43bd974b, 32'hc302a4b2},
  {32'h434e629e, 32'hc2a6b940, 32'hc1f886ac},
  {32'hc412938a, 32'h429093c8, 32'h432b982a},
  {32'h44ae8faa, 32'hc29629ee, 32'hc2a682c2},
  {32'hc4a52526, 32'h4397d978, 32'h43f03976},
  {32'h444dec0d, 32'h42f107bb, 32'hc2e5f576},
  {32'hc517e8d9, 32'hc188ff92, 32'h43fa5abd},
  {32'h44df631d, 32'h431916cb, 32'hc3000966},
  {32'h434418f0, 32'hc300674a, 32'h3fa85630},
  {32'h440fbf7c, 32'h42d92b8c, 32'hc3aeab1c},
  {32'hc45fdc18, 32'h420187b4, 32'h434a2b8a},
  {32'h436478f8, 32'h434d3337, 32'h43011174},
  {32'hc4cddf7a, 32'hc392fc98, 32'h429353df},
  {32'h44e50698, 32'h42d188fa, 32'hc3fc8287},
  {32'hc48e5b84, 32'hc216e3e4, 32'h43798c48},
  {32'h45177201, 32'hc3a71ea2, 32'hc33ca8bc},
  {32'hc48d3de8, 32'hc329f541, 32'h439bac08},
  {32'h44470c80, 32'hc40f3e9f, 32'h430128f3},
  {32'hc482a87c, 32'h42e3caa0, 32'h41039790},
  {32'h43bc7050, 32'hc2b34517, 32'hc345878e},
  {32'hc4e2c24d, 32'h442c0df4, 32'h43d0330f},
  {32'h4455aaa4, 32'hc3416e1f, 32'hc3d292e0},
  {32'hc4f53bac, 32'h42c87e5a, 32'hc2ba80f4},
  {32'h450bcbc5, 32'hc30e30a0, 32'h433d64d6},
  {32'hc4f4b391, 32'h42446c39, 32'hc3621639},
  {32'h44c11bfc, 32'h43a71acd, 32'hc25473fc},
  {32'hc499323e, 32'hc37094c8, 32'h4343e72d},
  {32'h44e8dbac, 32'h42ef1388, 32'hc2b5f11c},
  {32'hc40afb8f, 32'hc38ac101, 32'hc360d79e},
  {32'h44524344, 32'h42a30f8d, 32'h41f98948},
  {32'h40cc4a00, 32'h43049f75, 32'hc41f3ca6},
  {32'h44957efc, 32'hc2d43a75, 32'hc2616d6e},
  {32'hc268b976, 32'hc2e13b39, 32'h43bcaaea},
  {32'h44e4da76, 32'h4146bab0, 32'h4287d735},
  {32'hc1d37164, 32'h429b9e5d, 32'h42a62fe8},
  {32'h44097f5e, 32'hc2e823a3, 32'h434395b7},
  {32'hc4dbc110, 32'hc23c879a, 32'h43297f01},
  {32'h43116e50, 32'h435c41a3, 32'h432e8a4b},
  {32'hc4e3a01a, 32'h434bd410, 32'h40d0f4a6},
  {32'h45120826, 32'h432c58ad, 32'h43d0372a},
  {32'hc4bd501a, 32'h42bf6c07, 32'h4387b74d},
  {32'h430f6da8, 32'h42dc4d96, 32'hc40e438d},
  {32'hc4b9c8da, 32'h4275fb0d, 32'hc1bc6cc6},
  {32'h4339779f, 32'h42854afd, 32'h418dfc88},
  {32'hc4dd4d8f, 32'h43a0ad25, 32'h42fa4a02},
  {32'h44f8b930, 32'h43a0b436, 32'h43b50345},
  {32'hc52255f8, 32'hc3b0a71b, 32'hc31fab9a},
  {32'h447c53dc, 32'hc3107922, 32'hc2f91bba},
  {32'hc47d79dc, 32'h41a4b8ec, 32'h42d603b9},
  {32'h442cb7a2, 32'hc3d2f1bf, 32'hc1e9f441},
  {32'hc3ac14a8, 32'hc2093f3d, 32'hc3528f1f},
  {32'h44bd203e, 32'h422d580b, 32'hc2df0177},
  {32'hc4eff50e, 32'h43d9d33b, 32'h43a2d2cf},
  {32'h44590a75, 32'hc12ab258, 32'h42e1a9d8},
  {32'hc350f2a0, 32'h42bce9ac, 32'hc2efe921},
  {32'h4518255e, 32'hc24066a2, 32'hc35119c6},
  {32'hc3c42f58, 32'hc3345827, 32'h431bf388},
  {32'h448e5224, 32'h42a6b2f5, 32'hc3920155},
  {32'hc4cd99c7, 32'h4302a97c, 32'h442b8d6a},
  {32'h45186d6b, 32'h430ed31a, 32'hc3a59d55},
  {32'hc3fcd374, 32'h43351119, 32'hc386b883},
  {32'h440b9766, 32'hc3163f22, 32'hc378c956},
  {32'hc4253a69, 32'h410020b9, 32'hc3105d1c},
  {32'hc1602e00, 32'h429bd4b0, 32'hc3aac967},
  {32'hc3a387a0, 32'hc2cf77c5, 32'h4367af0b},
  {32'h449aee86, 32'h422cb13f, 32'hc3a4dd37},
  {32'hc3fa3b10, 32'hc23bdd9b, 32'h42f3f674},
  {32'h44e6de79, 32'h4274393b, 32'hc3c2112d},
  {32'hc4df6e3d, 32'h40d4d6e2, 32'h42c9711a},
  {32'h44bdbc4c, 32'hc412bd63, 32'h436499af},
  {32'hc4bfbeb3, 32'h434607e9, 32'hc3a44591},
  {32'h43b573c6, 32'hc381d220, 32'hc3baa769},
  {32'hc50124a7, 32'h43489088, 32'h43e38d42},
  {32'h442c024e, 32'h43d3d8e6, 32'h42d48ef8},
  {32'hc4d33493, 32'hc36963b5, 32'hc2384343},
  {32'h44b42740, 32'hc295ea3c, 32'h420f502c},
  {32'hc4cebd40, 32'hc3486584, 32'hc1a0874c},
  {32'h44840f2f, 32'hc2333934, 32'h4192c067},
  {32'hc4221746, 32'h42c25980, 32'h43bf8dd1},
  {32'h44fd3258, 32'hc1f6782f, 32'hc358b9a0},
  {32'hc31b34ec, 32'h4371b7ae, 32'hc124a1d0},
  {32'h44383428, 32'hc1fad810, 32'hc26cdb6b},
  {32'hc4251acc, 32'hc3de3802, 32'h4342239f},
  {32'h44fc7cb7, 32'hc08904fe, 32'hc3182c8d},
  {32'hc4b8ee62, 32'hc3358745, 32'h439f3e40},
  {32'h44c53d01, 32'hc1ddc41b, 32'h422d5723},
  {32'h441762c0, 32'hc37fbf73, 32'hc39d1ae8},
  {32'hc4a0acb5, 32'h43b45b8e, 32'h43a19228},
  {32'h4476b221, 32'h433cd7e1, 32'hc32466e6},
  {32'hc2fd7568, 32'hc156ff12, 32'h4395e2ca},
  {32'hc320ba60, 32'hc35138f9, 32'hc2b84e5b},
  {32'hc402b5a8, 32'h41d07078, 32'h4061fb42},
  {32'h443b64c9, 32'h423e5604, 32'hc0ebbd87},
  {32'h43215ba6, 32'h43ce0e7e, 32'hc2c3cb63},
  {32'h438c41d0, 32'hc382cf86, 32'hc2d77461},
  {32'h446fef27, 32'hc3696599, 32'h43937ea6},
  {32'hc4c933ce, 32'hc28eb6f6, 32'hc2a2e80b},
  {32'h44aa83a9, 32'hc2f7da1a, 32'h432f10bb},
  {32'hc4c74bc2, 32'hc288600f, 32'h43ed103e},
  {32'h4492f021, 32'hc36098b7, 32'h42dfaa58},
  {32'hc501173d, 32'h4297607f, 32'h428a9274},
  {32'h442878a8, 32'h437fb75d, 32'hc3ca7d6b},
  {32'hc4eba6d0, 32'h437f750e, 32'hc1bcc2b4},
  {32'h4514d676, 32'hc39eb417, 32'h405acfae},
  {32'hc51dfd29, 32'h4377f6e9, 32'h43250b08},
  {32'h4440b45c, 32'hc22320d7, 32'hc39997c2},
  {32'hc4e4d55c, 32'hc303021e, 32'h437a194e},
  {32'h450c6b86, 32'h43517767, 32'hc20e5cfd},
  {32'hc4b7dc31, 32'hc2c79d37, 32'hc3370e45},
  {32'h430a40fd, 32'hc32e999e, 32'h42c0a4cf},
  {32'hc51646fc, 32'hc3514111, 32'hc32342cb},
  {32'h445df447, 32'hc34f1c71, 32'hc3ad5475},
  {32'hc438198e, 32'h42a201f9, 32'h42607147},
  {32'h44c267be, 32'hc359a94f, 32'hc4031595},
  {32'h42f62ea0, 32'hc308b50c, 32'hc205c8f2},
  {32'h450a4f3c, 32'hc228b116, 32'h431ff3d6},
  {32'hc4b6fbb0, 32'hc335caaf, 32'hc3367b7c},
  {32'h44845446, 32'h43431c44, 32'hc371f65f},
  {32'hc3af3ef0, 32'h42c3657a, 32'hc19e5916},
  {32'h45086100, 32'hc25e8e6d, 32'hc1e34a38},
  {32'hc497bbf8, 32'h420dd219, 32'h438e51f0},
  {32'h444c855c, 32'hc3b1a739, 32'hc2a2e9dc},
  {32'hc4ebfaaf, 32'hc3b6aa63, 32'hc2b11390},
  {32'h44157169, 32'h43344a96, 32'hc3b1bf66},
  {32'hc46f461c, 32'hc387c5be, 32'h41cf6347},
  {32'hc2cb46a8, 32'hc3712b79, 32'hc3741ba6},
  {32'hc3c3146b, 32'h4287740c, 32'h42e7cea2},
  {32'h44790dc6, 32'hc3628b49, 32'h43120e76},
  {32'hc4706adf, 32'hc2ac0bea, 32'h43321ccc},
  {32'h44c11874, 32'hc2089f31, 32'hc303a09f},
  {32'hc439f342, 32'hc31711db, 32'hc3e9f865},
  {32'h44471092, 32'h425028c4, 32'h43b9fe0e},
  {32'hc43f7386, 32'h438a801c, 32'hc4026ec4},
  {32'h44bb1349, 32'h3fbdc27d, 32'hc28343fe},
  {32'hc462daec, 32'h43b64925, 32'hc095eced},
  {32'h43235d0a, 32'hc3251cad, 32'hc3d71d88},
  {32'hc45690a4, 32'hc1ae79f9, 32'hc164b8d4},
  {32'h451c5bf2, 32'h42c69c5f, 32'hc33d0c40},
  {32'hc4ce8e83, 32'h42c01af0, 32'hc27a57d6},
  {32'h4406af06, 32'h4310a011, 32'hc37aee99},
  {32'hc49d32a7, 32'h4352359d, 32'h4233a6fc},
  {32'hc34f481a, 32'hc20c4199, 32'h4377398f},
  {32'hc48a766d, 32'h41d2b285, 32'hc2f263b4},
  {32'hc491a6fa, 32'h429bf8ea, 32'hc24189a5},
  {32'h441b6998, 32'hc2d37f4b, 32'hc2bdc875},
  {32'hc4b84a64, 32'h41c9e423, 32'hc2006a57},
  {32'h44b28e6f, 32'hc362fd63, 32'hc3239790},
  {32'hc4c5a232, 32'h44029ec2, 32'hc36a1a86},
  {32'h448b9546, 32'h43b0be3b, 32'hc29d8257},
  {32'hc41b7095, 32'hc19fa21f, 32'hc2b3c749},
  {32'h451565fd, 32'h4394fd11, 32'hc34cc83c},
  {32'h44841b9b, 32'hc339351a, 32'h4320d785},
  {32'hc47306a8, 32'hc2823817, 32'hc4019285},
  {32'h44d67d58, 32'h42f912eb, 32'hc22904e3},
  {32'hc481d028, 32'hc3814a13, 32'h41c404a3},
  {32'h450e39a4, 32'hc2e30259, 32'h43d29d4a},
  {32'h44fa3ffa, 32'h444db019, 32'hc38914db},
  {32'hc3b08aa8, 32'hc3471ed6, 32'h432eda42},
  {32'h43af4864, 32'h439f0520, 32'hc382888a},
  {32'hc393bff2, 32'hc280e909, 32'hc2877c68},
  {32'h44e20252, 32'hc13eec9e, 32'hc2435102},
  {32'hc4091846, 32'h438b2f0a, 32'h42b1189b},
  {32'h44d329a4, 32'h431e1203, 32'h401296fe},
  {32'hc50eba8f, 32'hc3aedeff, 32'hc323ea2f},
  {32'h44b3f519, 32'h441150e8, 32'hc112783b},
  {32'hc48d6738, 32'h42ca77dd, 32'h432b110e},
  {32'h4470e3bc, 32'h43931922, 32'h43b841f9},
  {32'hc448e036, 32'h440771b0, 32'hc39ca3ee},
  {32'h450388c7, 32'h426dcf39, 32'hc30a0681},
  {32'hc4e14d2d, 32'h43d81b15, 32'h438ebca1},
  {32'h44346665, 32'hc3dbdf45, 32'h431be62a},
  {32'hc50d8043, 32'hc3d56c8b, 32'h4309d904},
  {32'h450f7151, 32'hc23e9449, 32'h43bdd7bf},
  {32'hc4ae06a2, 32'hc2886bcc, 32'hc352e578},
  {32'h44a1bc1a, 32'h440abe59, 32'hc30fa38f},
  {32'hc3a5ded0, 32'h424ed4bc, 32'hc307a40d},
  {32'h43f8ca18, 32'hc3a3ee67, 32'hc0a3166b},
  {32'hc34333f0, 32'hc3e3718c, 32'hc3254f65},
  {32'h44e5c8ee, 32'h42a6d7ab, 32'hc390d1a6},
  {32'hc4fc5468, 32'hc1ab4e26, 32'hc3b02bbd},
  {32'h437a16d8, 32'h431da5d2, 32'h4344ab8c},
  {32'hc412d5b0, 32'h431e57e5, 32'hc3047061},
  {32'h43bb2fc8, 32'h419ddb72, 32'h4237f379},
  {32'hc4730e6f, 32'h43184e62, 32'hc10a3d34},
  {32'h43d244d0, 32'hc35bbfa6, 32'hc2bb5724},
  {32'hc4b7f447, 32'h422fd1b3, 32'hc153abb7},
  {32'h4508efab, 32'hc2ead9a4, 32'h41e23184},
  {32'hc430ac40, 32'h420945ec, 32'h43d4943f},
  {32'h44116b1a, 32'h432e41d4, 32'h4385f5fd},
  {32'hc4ba8fc7, 32'h4397dab9, 32'h43b15b93},
  {32'h44c34bfd, 32'h42ffe6f1, 32'h43337e81},
  {32'hc4d18490, 32'h41844be1, 32'hc3a787f7},
  {32'h450ac798, 32'h43eccfdc, 32'h435b4a3b},
  {32'hc4c6f595, 32'hc354b2bd, 32'h42dc0f33},
  {32'h43bee558, 32'hc34fa23e, 32'hc205f24d},
  {32'hc483a2ea, 32'h43036116, 32'h431de762},
  {32'h4500e8ba, 32'hc1a296cb, 32'hc2cf193f},
  {32'hc408d405, 32'h41286bb0, 32'hc28ec45b},
  {32'hc2d0f6b0, 32'h438e01a6, 32'h43896588},
  {32'hc4837f33, 32'hc2a1429a, 32'hc2f9c090},
  {32'h443e1091, 32'h43b7f3a5, 32'h42f3ed61},
  {32'hc4b857f2, 32'hc3951e5f, 32'hc3209d92},
  {32'h441e4013, 32'hc3cd7912, 32'hc1adf036},
  {32'hc4fe58ee, 32'h432cf9d9, 32'h42cadbf9},
  {32'h450f9df4, 32'h43217932, 32'h42a3ea98},
  {32'hc37d15f0, 32'h4254a3b8, 32'h436b53a4},
  {32'h450ea5c7, 32'h4389f428, 32'h433c13b2},
  {32'hc4be859d, 32'h41ea7bba, 32'h43462da3},
  {32'h44436b72, 32'h40a80f04, 32'h43549c72},
  {32'hc47f78c9, 32'h42509bc9, 32'hc2d65f40},
  {32'h45032057, 32'hc424fdbb, 32'hc06dff40},
  {32'hc5076921, 32'hc3e8a273, 32'h41f7243a},
  {32'h444dba6e, 32'hc2fab8ae, 32'hc2ddd490},
  {32'hc4ab7137, 32'hc2e4f0ab, 32'h4239c1ac},
  {32'h44b707c2, 32'h426c9930, 32'h4272e43c},
  {32'hc3d84018, 32'h438e5281, 32'h430947ee},
  {32'h44e73c5d, 32'h43aa69f7, 32'h3fa34ab0},
  {32'hc4b10f04, 32'h4248a9ff, 32'hc2c75ad2},
  {32'h44e64081, 32'h4212ec32, 32'hc34c5fc1},
  {32'hc48770f6, 32'hc338a2dd, 32'hc2bb7564},
  {32'h43f26990, 32'hc3aaa945, 32'h41f444f3},
  {32'hc45bd277, 32'h43b9b88a, 32'h433e0ce2},
  {32'h4443b13a, 32'hc3976c87, 32'h435ed172},
  {32'hc4b31457, 32'h43a2b860, 32'hc3a77cd5},
  {32'h44416936, 32'hc3024cdb, 32'h422ee60f},
  {32'hc32d9d01, 32'h42ba79e5, 32'h4311aeeb},
  {32'h4458fedb, 32'hc294e806, 32'hc37d8a17},
  {32'hc4c8892f, 32'hc40cb6df, 32'hc37920c0},
  {32'h44c640c4, 32'h4239b79d, 32'hc207b3a1},
  {32'hc52add05, 32'hc242b85a, 32'h4398a8b2},
  {32'h444341a6, 32'hc1f6e57d, 32'hc2df18d7},
  {32'hc41b7db9, 32'hc35fa23e, 32'h42b710ec},
  {32'h446db1b0, 32'h41343174, 32'h434089fc},
  {32'hc4313ed5, 32'hc37a2ec9, 32'h42f0142c},
  {32'hc2e17664, 32'h40bffb5e, 32'h43a42b67},
  {32'hc4203d3e, 32'hc36523f3, 32'h43422fcf},
  {32'h4500d9b0, 32'h418dccf2, 32'h430985cf},
  {32'hc47ee93f, 32'hc2dc3878, 32'hc3e91fa3},
  {32'h448713f8, 32'hc2e77d09, 32'hc20adabb},
  {32'hc4b1c814, 32'hc3612a0f, 32'hc3c902bb},
  {32'h444ec39a, 32'hc345df1f, 32'h3e75a1a0},
  {32'hc30d6924, 32'h4228b8f6, 32'hc37f0621},
  {32'h443554f8, 32'h43947142, 32'h43024ba9},
  {32'hc5158940, 32'h43c3c0de, 32'h433116db},
  {32'h4483d452, 32'h4413e760, 32'hc39d300c},
  {32'hc45b2921, 32'h436662a2, 32'hc364ba43},
  {32'h416b6a80, 32'h429b4e92, 32'h4283ea03},
  {32'hc512beb4, 32'hc2bc844c, 32'h43262d2e},
  {32'h44f027a1, 32'hc2621043, 32'hc2d3f9a3},
  {32'hc500bfef, 32'hc387b697, 32'hc36cabc6},
  {32'h44fc8d4c, 32'h4286bcca, 32'hc3060106},
  {32'hc4efb504, 32'h4411bf64, 32'hc3f2b49f},
  {32'h4475c558, 32'hc1d41983, 32'h441dc350},
  {32'hc4fef916, 32'h43137ea0, 32'hc3175e5a},
  {32'h4406f16a, 32'h422c3dde, 32'h437648fa},
  {32'hc4fd8c8b, 32'hc40b8de1, 32'hc2c09091},
  {32'h44951f7d, 32'hc20436b8, 32'hc3208b47},
  {32'hc4e3bda1, 32'hc3271471, 32'h4324500a},
  {32'h438f8858, 32'hc34053fa, 32'hc2992f84},
  {32'hc4946721, 32'hc2e65d9b, 32'hc227ce29},
  {32'h45004b4d, 32'hc39d151e, 32'h423e8ddf},
  {32'hc4e0ad9c, 32'hc2ecaff9, 32'hc20291b4},
  {32'h44098581, 32'h4367f73c, 32'h43122f99},
  {32'hc4bd808c, 32'h434630fe, 32'hc112ecb2},
  {32'h444597f2, 32'h42c43f3b, 32'h42d49868},
  {32'hc49dc6f0, 32'hc306f021, 32'h41c7c7fb},
  {32'h44bf70a8, 32'h433c5e0d, 32'h41a38224},
  {32'hc4ac0eac, 32'h4325f0a4, 32'hc1740c82},
  {32'h434fdee0, 32'h4212a7f8, 32'h4248b1c3},
  {32'hc42fcd92, 32'hc2b69dff, 32'h437ece9d},
  {32'h4506f804, 32'hbf8c1068, 32'h438986b4},
  {32'hc3d846f8, 32'hc1dbec47, 32'hc382cd75},
  {32'h44af4f4d, 32'h43ed7322, 32'h422e3b2d},
  {32'hc4fc73e6, 32'hc31f4181, 32'hc23f9882},
  {32'h4448961a, 32'hc2536d17, 32'h425ce371},
  {32'hc3c422c0, 32'hc2a19748, 32'h41d7e9b8},
  {32'h44a67647, 32'hc308445c, 32'h4261bdc0},
  {32'hc4b198ef, 32'h430d3bdb, 32'h40d4de00},
  {32'h44feee4a, 32'hc36cf641, 32'h43c61d9b},
  {32'hc3b81068, 32'hc2a9e5b6, 32'hc3461321},
  {32'h44825b4c, 32'h41ad2c64, 32'h42abf38d},
  {32'hc50dcb9a, 32'h411bd9b2, 32'h42722824},
  {32'h44ca30f3, 32'hc2fbd914, 32'hc2e5bad2},
  {32'hc502988d, 32'h42b388c5, 32'hc3f87df4},
  {32'h438541cc, 32'hc3154308, 32'hc1591af1},
  {32'hc4954fcf, 32'hc26e67d5, 32'h4337b12e},
  {32'h45193ca1, 32'hc30e8201, 32'h43955936},
  {32'hc4f3846a, 32'hc3439518, 32'h43155b7e},
  {32'h43dc2d88, 32'h41ae253e, 32'h43756429},
  {32'hc4db1dd9, 32'h42f0505d, 32'h428a6d61},
  {32'h449f3df4, 32'hc1b7eae2, 32'h42e4d00e},
  {32'hc4dd617b, 32'hc3914afa, 32'h4302688e},
  {32'h4466af8c, 32'hc3b56e59, 32'h43f78248},
  {32'hc4bbb1b4, 32'h439a5bf9, 32'h429b5f51},
  {32'h44b24e27, 32'h42ece971, 32'hc13a99c0},
  {32'hc4f0b6a2, 32'h41725b22, 32'h3f10f828},
  {32'h44080f76, 32'hc34cfc96, 32'h43448cf3},
  {32'hc4a89a12, 32'hc34a3697, 32'hc30fb203},
  {32'h447202d0, 32'hc2e2007b, 32'hc21517f1},
  {32'hc4b8fcb4, 32'h43f94e5d, 32'hc3419501},
  {32'h4466e294, 32'hc346a66f, 32'h430e91c4},
  {32'hc3c84080, 32'h437f14c6, 32'h42a791aa},
  {32'h440159f8, 32'h43c9412f, 32'hc3bbd0bd},
  {32'hc48f520b, 32'hc28593f1, 32'h42a20e37},
  {32'h44e215a6, 32'hc2d49770, 32'h4310ea8d},
  {32'hc49bea20, 32'hc36f6ff6, 32'h428bad37},
  {32'h4470bc16, 32'h42e9a0dc, 32'h4227e824},
  {32'hc48aeea9, 32'hc39ddffe, 32'hc29ce350},
  {32'h442ce41f, 32'h420b15bd, 32'hc31c22e8},
  {32'hc51382fc, 32'hc3012fad, 32'h43ef709d},
  {32'h4306c486, 32'hc1026bf4, 32'h43512190},
  {32'hc4b62cce, 32'hc31d9fc4, 32'h40ac1a88},
  {32'h4507b53c, 32'h42eab2d2, 32'h430eca6c},
  {32'hc4cda98d, 32'h42c868c4, 32'hc24d32ae},
  {32'h431ec320, 32'hc36db78f, 32'h40db76e8},
  {32'hc5172370, 32'h42c82098, 32'hc1f7b4d2},
  {32'h450f6002, 32'hc4159a64, 32'h432b78cb},
  {32'hc4c5c815, 32'hc2f7b433, 32'h42abf36a},
  {32'h44b34f1b, 32'hc39a5dc8, 32'h42d14103},
  {32'hc4bd49fa, 32'h43440e16, 32'hc353181d},
  {32'h451eb5f7, 32'hc3087086, 32'h427d3d02},
  {32'hc4cf2ae4, 32'hc3b1dc40, 32'h4353f585},
  {32'h44ed8a0c, 32'h439087b9, 32'hc38a6b2b},
  {32'hc4d36be9, 32'h43461c47, 32'hc30148be},
  {32'h4528926c, 32'hc38d8998, 32'h43989191},
  {32'hc509e40f, 32'hc1ab0c4d, 32'h428d7de5},
  {32'h44289fe4, 32'hc223cc54, 32'h430e480b},
  {32'hc49e275a, 32'h432f2722, 32'h42245eab},
  {32'h44f7b970, 32'h42255ad2, 32'h42332099},
  {32'hc508bedc, 32'h42100c5b, 32'hc2d4583b},
  {32'h450ad8eb, 32'hc322649c, 32'h412b2c97},
  {32'hc4bf9b9c, 32'hc21bfae8, 32'hc2d07e5f},
  {32'h4465bf76, 32'h438900af, 32'hc38a4eac},
  {32'hc37ecc5a, 32'h437b0c6e, 32'hc2eddcb6},
  {32'h43a56944, 32'h430b3710, 32'h42d08d71},
  {32'hc4e67663, 32'h439bc904, 32'h423288da},
  {32'h4463950e, 32'hc2da69da, 32'h430f0f79},
  {32'hc4fa41b0, 32'hc34b0d76, 32'h43b0a333},
  {32'hc28cdacc, 32'h413a3d58, 32'hc2db9ae7},
  {32'hc26fc2d4, 32'h42bca5d7, 32'h420cc769},
  {32'h4419969a, 32'h420624d0, 32'h417ffea7},
  {32'hc4a1300b, 32'h429f9684, 32'hc287f33f},
  {32'h44f1282e, 32'hc319aeec, 32'hc2673b37},
  {32'hc503ef1a, 32'h410477f8, 32'hc38b2a1d},
  {32'h450ad647, 32'h4380840e, 32'h41f1da1c},
  {32'hc4d00154, 32'h42926800, 32'h42733a79},
  {32'h444b33a1, 32'hc3b158ff, 32'hc3be2810},
  {32'hc49c888a, 32'hc187fb5c, 32'hc2e30d3e},
  {32'hc40f03f2, 32'hbfed0c68, 32'hc37e4de6},
  {32'h44b6600a, 32'hc29d4d81, 32'h42d183a2},
  {32'hc464d545, 32'hc37deff4, 32'hc1c17497},
  {32'hc299c92c, 32'h4400a8eb, 32'hc285b44d},
  {32'hc4b76b0c, 32'hc2a5a294, 32'hc3967d7d},
  {32'h42ceae60, 32'hc28e5341, 32'h43804968},
  {32'hc4a592df, 32'h43518f4d, 32'hc2b75805},
  {32'h442d7c31, 32'h431460c5, 32'h43f7b937},
  {32'hc3b48b38, 32'h42f08993, 32'hc2a8e825},
  {32'h4490f95a, 32'h430b3637, 32'hc2a49be1},
  {32'hc5011d53, 32'h426a6cb9, 32'hc2acaafc},
  {32'h4511dd19, 32'hc233a2af, 32'h4293bd77},
  {32'hc3052bf8, 32'hc2df7ec4, 32'h42d26d19},
  {32'h44f7bf5e, 32'h4342e9d0, 32'hc317364a},
  {32'hc49c3701, 32'h4333fabe, 32'hc2fc0a1c},
  {32'h439375dc, 32'hc155a9f3, 32'hc38dc736},
  {32'hc4945119, 32'h41d353c1, 32'hc30a0b6e},
  {32'h44440a72, 32'h43e15515, 32'hc0355cc0},
  {32'hc50e500d, 32'h41a8e875, 32'hc319a0f5},
  {32'h44034e5a, 32'h430ccd47, 32'hc33c2ce7},
  {32'hc3831f00, 32'h4341be0f, 32'h42a70fd7},
  {32'h440cce7c, 32'h4395cb77, 32'hc32f5d50},
  {32'hc4e4e236, 32'h4380546a, 32'h43829fb5},
  {32'h44ff22d3, 32'h42d244d3, 32'hc3948bfa},
  {32'hc424684e, 32'h420c3abd, 32'hc3d9a2d2},
  {32'h44f27a87, 32'hc265aac5, 32'h43b53966},
  {32'hc3acfe69, 32'hc33310cd, 32'h43a345df},
  {32'h4484a9ca, 32'h42374d12, 32'hc3b51d1d},
  {32'hc40620c4, 32'h428613eb, 32'h434e2529},
  {32'h4523d7dc, 32'h433a9a0a, 32'h43d67c52},
  {32'hc40f8c04, 32'h4216a599, 32'hc3931109},
  {32'h43596db0, 32'h438879d7, 32'h4296d5db},
  {32'hc4e7bfc4, 32'h438a38ef, 32'hc2206420},
  {32'h44bbe545, 32'h43a67493, 32'hc296895d},
  {32'hc4a389cc, 32'h44387f04, 32'hc1476387},
  {32'h451c147d, 32'hc3006d04, 32'h42b6031d},
  {32'hc3548540, 32'hc302d30a, 32'h420dd0a7},
  {32'h44fd143f, 32'hc2e60323, 32'hc3048305},
  {32'hc4bdceae, 32'h4270ba7d, 32'hc0a02223},
  {32'h44057382, 32'hc2b82ec5, 32'hc2d8b4d8},
  {32'hc51821df, 32'h41499102, 32'h43c653c4},
  {32'h44f2cbe8, 32'hc2fd0a58, 32'h4211ecf2},
  {32'hc4a1ce1d, 32'h43abbaa8, 32'h432f9d20},
  {32'h43b93de8, 32'hc3f56c47, 32'hc4002a30},
  {32'hc3e7198e, 32'h4328d725, 32'h43480614},
  {32'h44a5d22d, 32'hc3183e1c, 32'hc3c3baeb},
  {32'hc3c9cac0, 32'hc350ee01, 32'h43987eef},
  {32'h43915a14, 32'h42992a2f, 32'hc32d1db7},
  {32'hc478b148, 32'hc3a70bdd, 32'hc37e23aa},
  {32'hc28e69c8, 32'h4397a8bd, 32'hc2d40ae5},
  {32'h445b6460, 32'h428739b5, 32'h438423d8},
  {32'hc500cb89, 32'hc3ac8371, 32'hc31196ca},
  {32'h443e7eb8, 32'hc2422f33, 32'hc2a08070},
  {32'h426acf40, 32'hc2d685a4, 32'hc37bdfd8},
  {32'h44ff12ec, 32'hc34d4cf6, 32'h43a3409f},
  {32'hc5213ad6, 32'h41cfdf08, 32'h424159b3},
  {32'h452bdd80, 32'hc3d682df, 32'hc3b03a0b},
  {32'hc3572a60, 32'hc388db29, 32'h4228035a},
  {32'h43a8de79, 32'h432268b5, 32'hc3236b6e},
  {32'hc4d52f2c, 32'hc29f7400, 32'h43e7386b},
  {32'h44df5a95, 32'hc32e441d, 32'hc318b582},
  {32'hc4cbc7be, 32'hc3ec6adb, 32'hc3e169e8},
  {32'h45264d48, 32'hc3c1156d, 32'hc418dfe4},
  {32'hc403cb5f, 32'hc291a453, 32'h42c0b152},
  {32'h44add1b9, 32'h42005b6b, 32'h40cb28a6},
  {32'hc5087d1c, 32'hc237d31a, 32'hc2da23c1},
  {32'h447a5a9c, 32'hc35cced2, 32'h42e3cc93},
  {32'hc4e8cc21, 32'h42c39ae3, 32'hc3493940},
  {32'h44b11583, 32'h4370447d, 32'h418ae68c},
  {32'hc48c81ba, 32'hc22ae106, 32'h431e2e4f},
  {32'h44f84cfa, 32'hc39f4e66, 32'hc369d61c},
  {32'hc3accb90, 32'h436e383b, 32'h436f1354},
  {32'h443a5ae8, 32'hc29280d8, 32'h41fee78c},
  {32'hc490621a, 32'hc3267db3, 32'h43a4f92b},
  {32'h4406e8d4, 32'h43253e29, 32'hc31bb9fe},
  {32'hc4875886, 32'h43100422, 32'hc31a4738},
  {32'h45063d36, 32'hc230d9b5, 32'hc137375e},
  {32'hc2a4d503, 32'h41105b43, 32'hc398c056},
  {32'h44c5fda6, 32'hc337d179, 32'hc39bf487},
  {32'hc5080eb3, 32'h41a741af, 32'hc22b236b},
  {32'h4381c3bc, 32'hc2136eba, 32'h43955388},
  {32'hc5119e25, 32'hc3418866, 32'hc21edc12},
  {32'h44c6bae6, 32'h42fe9ec3, 32'hc34574f0},
  {32'hc3d49188, 32'h43233031, 32'hc34f4640},
  {32'h4511f53c, 32'hc28d62d5, 32'h43fa4916},
  {32'hc4e0dfa4, 32'hc23a638a, 32'hc297227a},
  {32'h4415e841, 32'h42ff779c, 32'hc2a9017c},
  {32'hc5021720, 32'hc3a4f094, 32'hc334388e},
  {32'h44d15f0f, 32'hc33c4d73, 32'hc2d9e3b5},
  {32'hc4cf769c, 32'h43c7e86f, 32'h434a80ac},
  {32'h45125345, 32'hc3021f6f, 32'hc3c1c917},
  {32'hc516389f, 32'h43812a50, 32'hc209a336},
  {32'h44a5635b, 32'h43101415, 32'h429c4936},
  {32'hc4dd0951, 32'h438a14aa, 32'hc28cdac8},
  {32'h45176a76, 32'hc3a0dd4d, 32'h42481daa},
  {32'hc43ffe67, 32'hc305efa7, 32'hc34a107c},
  {32'h44413eec, 32'hc329faa9, 32'hc3372c96},
  {32'hc4c9ddb9, 32'hc224199c, 32'h421e0884},
  {32'h4489de35, 32'h439bb356, 32'h43806f32},
  {32'hc3f41558, 32'hc43e9fe6, 32'hc2c0bc20},
  {32'h44c271c0, 32'h43474990, 32'hc3946d4f},
  {32'hc36befc8, 32'hc2ec709e, 32'h43b74bc9},
  {32'h44a8ae96, 32'h4221a5e9, 32'h43b535a3},
  {32'hc4c063e8, 32'h428fb1a8, 32'h4302115f},
  {32'hc43820fe, 32'hc235da49, 32'h421ef746},
  {32'h450ed012, 32'hc3b2d414, 32'hc395b504},
  {32'hc4c2f6ce, 32'hc3935247, 32'hc2eb68e5},
  {32'h4499fef9, 32'hc286a536, 32'hc39c5616},
  {32'h42cd0080, 32'hc34e1550, 32'hc31f1fe9},
  {32'h44c3f0d0, 32'h431c3b35, 32'hc409a70a},
  {32'hc493e2bb, 32'h428949ba, 32'hc180292f},
  {32'h450edc16, 32'h43a38eb3, 32'h40ea802c},
  {32'h431b96b0, 32'hc37f85a0, 32'hc34b34ec},
  {32'h446f157a, 32'h42cd0794, 32'hc38cb5fe},
  {32'hc45ada3c, 32'hc3cda820, 32'hc3115fb3},
  {32'h435386e0, 32'hc2cf8fab, 32'hc281e0b8},
  {32'hc2b7b840, 32'hc2291935, 32'h4229c774},
  {32'h44e6c45b, 32'h4383d9a8, 32'hc33b5620},
  {32'hc3b0738c, 32'h4329b51a, 32'h42f8cafc},
  {32'h44b26942, 32'h42d374d5, 32'h429f16f6},
  {32'hc5084fe0, 32'h4385ecbd, 32'hc37d2a73},
  {32'h440c4018, 32'h43302ed7, 32'hc421cdef},
  {32'hc51b40a1, 32'hc3c9ea48, 32'hc3873191},
  {32'h43bdb094, 32'h43283699, 32'hc17941bb},
  {32'hc4a38211, 32'h437579ef, 32'h41e52a33},
  {32'h44f4ade5, 32'h4330deb9, 32'hc22ede19},
  {32'hc4fe4ee5, 32'hc24e562d, 32'h43875c14},
  {32'h44f43fff, 32'hc28228aa, 32'hc31575eb},
  {32'hc45d43a4, 32'h41c241cc, 32'h437d13fd},
  {32'h44d476c7, 32'hc3022dbc, 32'h429290f0},
  {32'hc51c101f, 32'h43d77353, 32'h43571287},
  {32'h44eaa9c9, 32'hc2840818, 32'hc3126305},
  {32'hc47795b2, 32'hc2f5657f, 32'hc307bf9a},
  {32'h45104b1b, 32'hc37b54df, 32'h4345a828},
  {32'hc37b68ba, 32'hc35914f6, 32'hbf385c02},
  {32'h44c57fa0, 32'h438d31a0, 32'hc30214ae},
  {32'hc48ad5a4, 32'hc3bd94af, 32'hc39f05e3},
  {32'h44aa95f6, 32'h43456047, 32'h423dd6b3},
  {32'hc4d59b14, 32'h43701eb7, 32'hc34f8b7d},
  {32'h44de9852, 32'h42ad0044, 32'hc1e21436},
  {32'hc3c25a3c, 32'h4202f7a0, 32'hc2930068},
  {32'h440f0284, 32'hc2d66920, 32'hc294e362},
  {32'hc3278000, 32'h41e2ede7, 32'hc3af71d4},
  {32'h44cd135c, 32'hc2238924, 32'hc28b0b63},
  {32'hc48ae658, 32'h43d92209, 32'h4176087e},
  {32'h43c158f2, 32'h4317215d, 32'h43061578},
  {32'h41d3ec40, 32'h4359cb60, 32'hc0b2263b},
  {32'hc4de7382, 32'hc1ed76b0, 32'h426bfec7},
  {32'h44a9ef14, 32'hc0c655e7, 32'h439ee55a},
  {32'hc44b98b8, 32'hc3a11fab, 32'hc388b77a},
  {32'h44f00c7c, 32'hc2fdf148, 32'hc2002775},
  {32'hc4df8ecf, 32'hc20822a3, 32'h4384b86d},
  {32'h4490a282, 32'hc38f8633, 32'h42fb5fa0},
  {32'hc50a389f, 32'hc30d4ae3, 32'hc31cb7b8},
  {32'h442a4fb6, 32'hc2a16e11, 32'h43bab74f},
  {32'hc48328c8, 32'hc3819dba, 32'h42ad561d},
  {32'h45296c46, 32'h43903fee, 32'hc297c010},
  {32'hc454b512, 32'hc389b01b, 32'hc3844aee},
  {32'h44c62fc1, 32'hc32b3812, 32'hc02e019c},
  {32'hc478c0fe, 32'hc3b9cc58, 32'h42c3916f},
  {32'h443aaac7, 32'h3e735a80, 32'h4018af1b},
  {32'h424e9b38, 32'h3ee73740, 32'hc32d50e3},
  {32'h4443aaa0, 32'hc2538cd6, 32'h41bd1b28},
  {32'hc41a6aa5, 32'h43d55e40, 32'hc3cafd06},
  {32'h45091830, 32'hc16853fb, 32'h41b6030d},
  {32'hc4c8aeda, 32'hc3794b9a, 32'hc3906d19},
  {32'h44df635a, 32'h43ca9660, 32'h41f51b64},
  {32'hc4cd84fc, 32'h40a8c3cc, 32'hc312aa96},
  {32'h444e65ce, 32'h435d0e78, 32'h427c163b},
  {32'hc4c2c442, 32'hc35d8094, 32'h440bed2b},
  {32'h43edf0a2, 32'h434c0906, 32'hc355aa75},
  {32'hc39ac558, 32'hc2cb4cfa, 32'hc38190ef},
  {32'hc420e822, 32'hc29f0887, 32'h4303c1ea},
  {32'h44c3a552, 32'h43aff3b8, 32'hc3516373},
  {32'hc4a2ca6f, 32'h43dc4950, 32'hc393f643},
  {32'h44bb69d4, 32'h42a4d610, 32'h42f53697},
  {32'hc4f90e64, 32'hc245d4f5, 32'hc302d128},
  {32'h4489ad60, 32'h426ef315, 32'h44269d1b},
  {32'hc3978072, 32'hc2532c82, 32'hc340b087},
  {32'h44fe6525, 32'h42a3174a, 32'hc3cec8c9},
  {32'hc43db894, 32'hc381813f, 32'hc2ad17c0},
  {32'h44b36416, 32'h43a8fee6, 32'hc395ffcf},
  {32'hc4517f59, 32'h439f787d, 32'h43218f33},
  {32'h4471717e, 32'hc0b6c8dc, 32'h434f90aa},
  {32'hc3b5f2a8, 32'h4363f740, 32'hc38351ea},
  {32'h45109197, 32'h422aaa16, 32'h42b401eb},
  {32'hc4b080ce, 32'h4239048a, 32'h41e564df},
  {32'h42dedc3a, 32'h43856eb7, 32'h4302cae0},
  {32'hc4afeefb, 32'hc31a3246, 32'h43188152},
  {32'h43d3fad0, 32'hc39d061c, 32'hc29bb703},
  {32'hc4ac92e0, 32'hc2ed87cc, 32'hc210d7a6},
  {32'h42d2eddc, 32'hc2db6229, 32'h4368da4e},
  {32'hc37ea020, 32'hc3f4293c, 32'hc3f81294},
  {32'h440c181a, 32'hc38313bb, 32'hc2a31b87},
  {32'hc4a3d54c, 32'h42b61c65, 32'h43a346d0},
  {32'h448846c3, 32'h4285d073, 32'h43991849},
  {32'hc3ae7ee4, 32'h41f0f275, 32'h436e1352},
  {32'h44d0d0ad, 32'hc40bf7d7, 32'h43f6b307},
  {32'hc50f35b6, 32'hc108fc5d, 32'hc2cf90c5},
  {32'h449cf29e, 32'h43a9496d, 32'h438d8dec},
  {32'hc3925380, 32'hc3427831, 32'h4288caf1},
  {32'h4448b790, 32'hc35efbe0, 32'h42e4c3f1},
  {32'hc3ad41ec, 32'hc33c9971, 32'h42c4bf0b},
  {32'h43533b46, 32'hc3a9cac5, 32'hc29711f1},
  {32'hc4b9ae4b, 32'hc1f12b4c, 32'hc3386cd0},
  {32'h448b1b49, 32'hc2d9dfa9, 32'h42a419d4},
  {32'hc3be1e54, 32'hc30f1afc, 32'hc38c3164},
  {32'h450a769e, 32'hc3d9b1b1, 32'hc2a6d11d},
  {32'hc4452d83, 32'hc328634b, 32'h4328311a},
  {32'h44f48c86, 32'hc34f6175, 32'h4373ac83},
  {32'hc37c5254, 32'hc244a800, 32'hc26ba350},
  {32'hc2a86d88, 32'h41123998, 32'hc276f32a},
  {32'hc3818bc0, 32'h43d88ede, 32'h4370b84f},
  {32'hc50b06a4, 32'h41e1062e, 32'hc3197be3},
  {32'h450f9b77, 32'hc3ef034d, 32'h428336bd},
  {32'h423ebb9d, 32'hc2d61e89, 32'hc375a4e8},
  {32'h43e84248, 32'h3f10d920, 32'hc1640328},
  {32'hc4433e82, 32'hc2229cba, 32'h41a3855b},
  {32'h442cb702, 32'hc20aa567, 32'hc2096625},
  {32'hc31ee630, 32'h432539be, 32'hc2daf1ff},
  {32'h429f370a, 32'hc34325fd, 32'hc1df2b0d},
  {32'hc4020fdc, 32'h42ccac35, 32'hc379829d},
  {32'h4444a9ac, 32'h4102f3a8, 32'h42fdc285},
  {32'hc453b5e8, 32'hc29c1766, 32'hc3814674},
  {32'h44d8248f, 32'hc305d9b1, 32'h42a032b3},
  {32'h4323b894, 32'hc30823ef, 32'h41a3395a},
  {32'h44fbf71e, 32'hc317615f, 32'hc353e17c},
  {32'h43b337cb, 32'hc3e75b4c, 32'h43136a71},
  {32'hc3b3c7ec, 32'hc2028236, 32'hc3a87a16},
  {32'h4491f9db, 32'hc2913d47, 32'h4365eafa},
  {32'hc4b5779a, 32'hc20078bf, 32'h4258f5b7},
  {32'h43ce040c, 32'h41cc8f26, 32'hc3352799},
  {32'hc2ea7200, 32'h43b6c0c0, 32'h425002d6},
  {32'hc38a6010, 32'hc2e5ab12, 32'h436d32e2},
  {32'h4415fff4, 32'hc26fc471, 32'h43351b44},
  {32'hc3604760, 32'hc23cb933, 32'h434d1d1e},
  {32'h4499feb1, 32'hc3da9ff8, 32'h42af4f08},
  {32'hc4f9359e, 32'h433c5bdc, 32'hc28f9024},
  {32'h44ce79b8, 32'h43848e5d, 32'h438bddc6},
  {32'hc50dc191, 32'h428ed85e, 32'hc2045a5c},
  {32'h44f83e9c, 32'hc39359a2, 32'h429801d4},
  {32'hc4f21cb1, 32'hc36998fc, 32'hc1a6608f},
  {32'h445946b4, 32'hc22ef8f0, 32'h438cafe5},
  {32'hc2e06b00, 32'hc33cc574, 32'hc27e3d4c},
  {32'hc34fc405, 32'hc2a05138, 32'h42f3507b},
  {32'hc511197e, 32'hc2890243, 32'h42e0eeee},
  {32'h446e3118, 32'hc32b4473, 32'h42d72a9f},
  {32'hc44324e8, 32'hc3057159, 32'h4295bef7},
  {32'h44273822, 32'h42cdbd88, 32'h4364852e},
  {32'hc31dab30, 32'hc2d88610, 32'h418f0408},
  {32'hc4100274, 32'h4195cf90, 32'h431fb098},
  {32'h44d7ebce, 32'h4325c833, 32'hc33da3fd},
  {32'hc3efd860, 32'h435c88d1, 32'h43c375f4},
  {32'h45032043, 32'hc1953157, 32'h43e22df8},
  {32'hc33a442a, 32'h43981ead, 32'hc032bc39},
  {32'h44e3842e, 32'h437f5c96, 32'hc2ad909c},
  {32'hc42ec66a, 32'hc33805e3, 32'h43d10f68},
  {32'h45117bd7, 32'hc2dcf3c0, 32'hc3012435},
  {32'hc50cd97e, 32'hc343e7e5, 32'h42cc8ca1},
  {32'h43293d32, 32'hc3a55843, 32'hc36be76b},
  {32'hc4b35bac, 32'hc2db42bd, 32'h40f43aea},
  {32'h45047005, 32'h42d3f9d6, 32'h4396be7d},
  {32'hc35984b4, 32'h42b4348c, 32'hc2f1879a},
  {32'h4510b901, 32'hc0dc7c68, 32'hc2fc8db4},
  {32'hc4da9c26, 32'hc2e8c1e9, 32'h4250cf10},
  {32'h44c99e07, 32'h430339c5, 32'hc2b9f823},
  {32'hc3b01b2a, 32'h428180d0, 32'hc295f801},
  {32'h4497ba4a, 32'h431441a0, 32'hc385cd62},
  {32'hc43bb78e, 32'h429275ea, 32'hc3872919},
  {32'hc4f8587a, 32'hc2df0e91, 32'hc36f2cb0},
  {32'h43d9656e, 32'hc2c50064, 32'hc3497299},
  {32'hc4f5da0d, 32'hc2878701, 32'h431c1ebb},
  {32'h431271f7, 32'hc286a3d5, 32'h40ca2076},
  {32'hc501592d, 32'hc3a666af, 32'hc286d939},
  {32'h44b62d7d, 32'h42aff2ca, 32'hc29fe719},
  {32'hc4d90c1e, 32'hc2c61f17, 32'h4100a9eb},
  {32'h422c7320, 32'h43c9a130, 32'h43abda18},
  {32'hc34fb4d8, 32'hc310b748, 32'hc30294c3},
  {32'h432ad3c0, 32'hc2e9b483, 32'h430b228d},
  {32'hc442f283, 32'hc40ea2f9, 32'h44638df9},
  {32'h44968c05, 32'h43cc4022, 32'h42542463},
  {32'hc52110a2, 32'h4328be12, 32'hc19244ce},
  {32'h45089844, 32'hc32aece9, 32'h42602c46},
  {32'h43c517d8, 32'h431be7bb, 32'h43354ad6},
  {32'hc50de0b1, 32'h4425c277, 32'hc3d81648},
  {32'h44223735, 32'h43844f97, 32'h43adba11},
  {32'hc3a7132c, 32'hc2c2ea90, 32'h421f933f},
  {32'h44093cc2, 32'hc32f8718, 32'hc32e5146},
  {32'hc4f4a07a, 32'h42e52542, 32'h43e9fc28},
  {32'h44fdb82c, 32'hc342ceea, 32'h42c867b2},
  {32'h3ff69000, 32'hc1716080, 32'hc2b611d3},
  {32'h44deccc2, 32'h430c22d1, 32'hc30d9113},
  {32'h42dcc9a0, 32'hc2ae304d, 32'h41c20afe},
  {32'h4409ad8c, 32'hc3b00910, 32'hc2e92d1c},
  {32'hc4635f75, 32'h4384d102, 32'h4353fb3a},
  {32'h43541d4c, 32'h436617c5, 32'h43c53fb3},
  {32'h431c03ee, 32'h438fb0ae, 32'h433b6988},
  {32'hc417cb76, 32'h4309af23, 32'hc2aaf621},
  {32'h43a6e492, 32'hc2b4194d, 32'h438fd161},
  {32'hc4f87bf6, 32'h422fd9f4, 32'h43d7a623},
  {32'h4456219c, 32'hc315a80e, 32'hc3bf1200},
  {32'hc4791872, 32'hc258623c, 32'h41a0ca12},
  {32'h450a071b, 32'hc3bb92fe, 32'h4384f409},
  {32'h42e1232b, 32'hc3172baa, 32'h40da8fd9},
  {32'h449ca628, 32'h43c3558b, 32'h42365c01},
  {32'hc4b34c18, 32'hc3173820, 32'h431f58df},
  {32'h449a723c, 32'h446535ad, 32'h43877a06},
  {32'hc4f40dac, 32'h4348ea1b, 32'h43608da0},
  {32'h41e67680, 32'hc3f95f64, 32'hc2422bcf},
  {32'hc47c171a, 32'h42e08ebe, 32'hc20552a6},
  {32'h4506b26b, 32'hc336bd6a, 32'hc30c0a7b},
  {32'hc46b85ac, 32'hc34d7fc9, 32'hc3603930},
  {32'h44d94d42, 32'h43fbbae8, 32'h435cad80},
  {32'hc4b1f3b2, 32'hc3235dd5, 32'h438072db},
  {32'h4381b6a8, 32'h43cb2132, 32'h422bc5bf},
  {32'hc425a110, 32'hc2c3ec5c, 32'hc3401768},
  {32'h44e49d92, 32'h431f970a, 32'h427de201},
  {32'hc4bb157f, 32'hc2ec8cbf, 32'hc0ebd8b3},
  {32'h44c1bfd6, 32'hc2f102c9, 32'hc3205b41},
  {32'hc50d772e, 32'hc33f3d40, 32'hc2d3c591},
  {32'h4478780c, 32'hc32da3db, 32'hc3279110},
  {32'hc457520f, 32'h4203f5d1, 32'hc362ccee},
  {32'hc37cefa4, 32'h43025dba, 32'hc363d7a0},
  {32'hc4246444, 32'h43673a1b, 32'hc3c04ebe},
  {32'h44c6380a, 32'hc384b596, 32'h425cb08c},
  {32'h42f1c400, 32'hc35c98a2, 32'hc3cf2fa7},
  {32'h44f04a56, 32'hc2e97b8f, 32'h4159ea01},
  {32'h44e10f22, 32'hc3807ebb, 32'h41f5281b},
  {32'hc4c58d4f, 32'h4271d6dd, 32'hc36de8db},
  {32'h44651144, 32'h428a7d5c, 32'hc2a5d676},
  {32'hc4ba8934, 32'hc191ef54, 32'h42d506ed},
  {32'h4353c803, 32'hc25fd512, 32'hc1dce667},
  {32'hc3dbcac8, 32'h4419235e, 32'hc2f743fc},
  {32'h437aff40, 32'h42c50964, 32'hc38230eb},
  {32'hc4d7f5c1, 32'h43815ea8, 32'h43beb6d2},
  {32'h441dcb68, 32'hc3423398, 32'hc1552f1c},
  {32'hc43a3997, 32'hc0fa42d6, 32'h4386f3aa},
  {32'h4472c93a, 32'hc309516b, 32'hc3e377f5},
  {32'hc492caf8, 32'h43857536, 32'hc263c292},
  {32'hc22c4d30, 32'h43395260, 32'h42246d93},
  {32'hc4e94234, 32'h4223e406, 32'hc30ba8c3},
  {32'h450202f6, 32'h4312388e, 32'hc2a8211f},
  {32'hc33e44b8, 32'h43afe177, 32'hc4436ac9},
  {32'h43bee08e, 32'hc354718b, 32'h436c9fb5},
  {32'hc42dba2e, 32'hc32b2dec, 32'hc026650b},
  {32'h44a6fdea, 32'h4254e7d3, 32'h40b1eff8},
  {32'hc434741e, 32'h4325a2d3, 32'hc30fe48c},
  {32'h43c655d0, 32'h43d408f2, 32'h440636ab},
  {32'hc4df7cac, 32'hc31d03f5, 32'h4351bf4e},
  {32'h414bf480, 32'hc128a2a4, 32'hc0b4c2d2},
  {32'hc49a9fb2, 32'hc233c876, 32'h42320a4c},
  {32'h45001f34, 32'h422bf087, 32'h425f7dd8},
  {32'hc47a9779, 32'h4321fdc3, 32'h418a5602},
  {32'h44e15d7a, 32'hc34311b3, 32'hc39d5df8},
  {32'hc4dcec12, 32'hc3e3235f, 32'hc3a9c800},
  {32'h44895068, 32'h4396cc6f, 32'hc2e79d18},
  {32'hc3441d33, 32'h42230123, 32'hc30bcd5f},
  {32'h4387e82c, 32'h431f5280, 32'h438a8827},
  {32'hc4c4e95c, 32'hc25f1436, 32'hc312eebb},
  {32'h44d79016, 32'h434f4db4, 32'hc43e3afb},
  {32'hc41b97ae, 32'h42a50957, 32'h437dcedb},
  {32'h44f96b8a, 32'hc3109143, 32'h428add45},
  {32'hc4824721, 32'hc35d1b34, 32'hc37af9d6},
  {32'h446ca48e, 32'h426cdeb2, 32'hc281c9bd},
  {32'hc5020945, 32'h42dcd627, 32'h4284e343},
  {32'h44a93804, 32'h42e1d646, 32'h437abcd3},
  {32'h43739410, 32'hc3cab552, 32'h4349eeaa},
  {32'hc5095130, 32'h4337da6d, 32'h425045a6},
  {32'h44939772, 32'h421280ec, 32'h41fc48ca},
  {32'hc4e50251, 32'hc388f642, 32'h42e85eb8},
  {32'h44cfba78, 32'hc23cba94, 32'hc3853403},
  {32'hc4bc7cbe, 32'h429b66a5, 32'hc31b5fd1},
  {32'h44f527c6, 32'hc2fe5aac, 32'h426c5fba},
  {32'hc4da33ce, 32'hc23eaf7a, 32'h43cfc9a5},
  {32'h448ea3b8, 32'h41dbcdf1, 32'h42481588},
  {32'hc4e6f535, 32'h42c5eac9, 32'h4321b817},
  {32'h43e14221, 32'h431007c0, 32'hc35d2cdc},
  {32'hc5022978, 32'hc1573804, 32'h42871f27},
  {32'h44fc3a5d, 32'h431f5481, 32'hc301de24},
  {32'hc37947d0, 32'hc2763cd0, 32'hc3913f28},
  {32'h4431dd66, 32'hc3868558, 32'h4313cb14},
  {32'hc47eda11, 32'h4162425a, 32'h43582ce2},
  {32'h44eb2c3b, 32'hc29a737e, 32'h42d6d5d5},
  {32'hc45e0fa3, 32'h41a02dd1, 32'hc2f84693},
  {32'h44da6073, 32'hc367872f, 32'hc278de46},
  {32'hc4066b15, 32'h42ea17e7, 32'hc39739e0},
  {32'hc388e9ea, 32'hc3db20bf, 32'h43d69e3f},
  {32'hc4e23ec9, 32'hc2a02a6c, 32'h438f22d1},
  {32'h44d63fea, 32'hc36efe77, 32'h434d55f8},
  {32'hc3f6eb5c, 32'hc371deab, 32'hc340aade},
  {32'h450e2fe8, 32'h44150f6a, 32'hc28bf4bb},
  {32'hc3c19110, 32'hc355b6f2, 32'h436a0a21},
  {32'h4496c7f8, 32'hc3c3ac42, 32'hc381176c},
  {32'hc4180bfe, 32'h43978829, 32'h437a77f8},
  {32'h44a3b550, 32'h4347ed72, 32'hc32252d2},
  {32'hc4440340, 32'hc31a23fb, 32'hc328ba23},
  {32'h44362692, 32'hc375bc56, 32'hc26aa2ba},
  {32'hc508dd2a, 32'hc1a2358f, 32'hc379e0df},
  {32'h43b86627, 32'h43022ee6, 32'h418aaea8},
  {32'hc3eeb378, 32'h4252c82f, 32'hc1eb6354},
  {32'h44b55140, 32'h42f125ce, 32'hc2955915},
  {32'hc42161a6, 32'hc3a23fa5, 32'h41796830},
  {32'h440eb35b, 32'h42ce6b75, 32'h426c3310},
  {32'hc437f080, 32'hc327eb67, 32'hc38a6221},
  {32'h448724bc, 32'h42838d4c, 32'h40c2a11d},
  {32'hc41293c0, 32'hc2b3f594, 32'hc243bfa0},
  {32'h44872a89, 32'h4307da2a, 32'h420672b4},
  {32'hc4f6a055, 32'hc3e3b05b, 32'h43e00471},
  {32'h440aef38, 32'h4387716e, 32'h437c1b7c},
  {32'hc3aba658, 32'hc36e5adb, 32'hc2e0d032},
  {32'h43ba35b0, 32'h42e18710, 32'hc356a936},
  {32'hc221a880, 32'h43342f77, 32'h42a6b09b},
  {32'h44b121c0, 32'h43b0173e, 32'hc33a412e},
  {32'hc3f17a60, 32'hc2560b6e, 32'h4316d963},
  {32'h44a283fa, 32'h41c5116e, 32'h42e33633},
  {32'hc4b83f3e, 32'hc35d7331, 32'hc1abffba},
  {32'h44dc638a, 32'h41ab6c9f, 32'hc2c6751c},
  {32'hc48e5ffb, 32'hbf8a1cfe, 32'h42a398c2},
  {32'h43e27af7, 32'hc3c40e64, 32'h43edda01},
  {32'hc414e733, 32'hc37b4abb, 32'h422be36d},
  {32'h44d17433, 32'h43b3702e, 32'h4331d311},
  {32'hc4db6682, 32'h43e89d99, 32'hc377487f},
  {32'h45079a94, 32'hc2ab3537, 32'h4368f45c},
  {32'hc4bbc1ff, 32'h4288e0ff, 32'h42235322},
  {32'h447a77fe, 32'h435a9159, 32'h432fcd7b},
  {32'hc5022daa, 32'hc1e4da13, 32'h434d78ee},
  {32'h4429da02, 32'hc355137d, 32'h43ba7bb3},
  {32'hc4773943, 32'hc328b4b2, 32'hc3277756},
  {32'h450e1854, 32'h43d6da5a, 32'hc1f0f2eb},
  {32'hc4302fda, 32'h43f516ef, 32'hc34b3921},
  {32'h441a4a44, 32'h43ab8e1c, 32'h4280c8be},
  {32'hc427ea1d, 32'hc32e50fa, 32'h43303c04},
  {32'h44ba769e, 32'hc30cacc4, 32'h43e9bf51},
  {32'hc48afa5f, 32'h42490801, 32'h418fddb8},
  {32'h44a96b73, 32'h43aa998d, 32'h433ce205},
  {32'hc45065dd, 32'h4194eaf1, 32'h438914f1},
  {32'h4494a203, 32'h43322744, 32'hc296f260},
  {32'hc4ad341b, 32'hc399a86a, 32'h4348d34c},
  {32'h4503324c, 32'h42e0d4c0, 32'h422afe5d},
  {32'hc464d34b, 32'hc2664576, 32'hc300b94b},
  {32'h43646a40, 32'hc3a5020b, 32'hc2856656},
  {32'hc497de2c, 32'h430e3d89, 32'hc33f5e5f},
  {32'h44de46f8, 32'h42f8d668, 32'hc2346e0f},
  {32'hc50e1ce6, 32'h439b727c, 32'hc2f5beee},
  {32'h443c703a, 32'hc2843f45, 32'h42d577d0},
  {32'hc4a95464, 32'h426f7baa, 32'hc2ad7b0e},
  {32'h4493981d, 32'hc1b64430, 32'h430c469f},
  {32'hc4ccc6aa, 32'h431e1142, 32'h431504aa},
  {32'h45101631, 32'h4329ed0a, 32'h438e39ae},
  {32'hc4d83b30, 32'hc3033436, 32'h4347319a},
  {32'h45013bf3, 32'h43f16f52, 32'h433efbd2},
  {32'hc501da37, 32'hc345a0a3, 32'h42a280ca},
  {32'h44c11203, 32'hc38dd3e5, 32'h3ff98bc6},
  {32'hc30ea490, 32'hc362453a, 32'h42029d56},
  {32'h44eb8ead, 32'hc254aca8, 32'hc20996cf},
  {32'hc3a372da, 32'hc3510d6a, 32'hc397f6b4},
  {32'h4504c3a8, 32'h438d09f7, 32'h43c4602d},
  {32'hc49b0b5a, 32'h435f6636, 32'h43c3b12b},
  {32'h44f64fd8, 32'hc3ec9626, 32'h4150c0f7},
  {32'hc4ffa636, 32'h41dc7220, 32'hc302765d},
  {32'h44ca83fe, 32'hc28f7cb5, 32'h4384d621},
  {32'hc427e568, 32'h44350107, 32'hc2356ce2},
  {32'h448a74b6, 32'h43340599, 32'hc150eb9b},
  {32'h4348ac60, 32'hc1d3dc7b, 32'h429f3afc},
  {32'h44c3749e, 32'h423411f4, 32'hc3905238},
  {32'hc4ce7b33, 32'h43491342, 32'hc2a11c17},
  {32'h44ce1e4d, 32'h42c89206, 32'hc378719f},
  {32'hc479f86a, 32'h42811171, 32'h42435c0e},
  {32'h445c86bf, 32'hc2c6fae9, 32'h4284c26e},
  {32'hc47463d2, 32'h41c6b3f2, 32'h43589936},
  {32'h43f4c025, 32'hc304fcc2, 32'h42c1665c},
  {32'hc4c4eda1, 32'h42e07939, 32'hc36d4a03},
  {32'h4505e12d, 32'h43ca05fe, 32'h4338a257},
  {32'hc42ed9a2, 32'hc3038fdb, 32'hc35979b6},
  {32'h45174b00, 32'h42d5b56d, 32'hc21aac48},
  {32'hc47ce784, 32'hc1c497ee, 32'hc0b7f353},
  {32'h44c50786, 32'hc39e82ec, 32'hc315d0b6},
  {32'hc40762d2, 32'hc3a50955, 32'hc2b43583},
  {32'h435adea8, 32'hc3cdbe79, 32'h43e8b2d1},
  {32'hc4fcbec3, 32'h42d495eb, 32'hc35eafed},
  {32'h450aea89, 32'hc3925d88, 32'hc306d498},
  {32'hc4a963d0, 32'hc2b05827, 32'hc29983ff},
  {32'h44b2d2a3, 32'hbf95cac8, 32'h41b6ea7d},
  {32'hc3dc9278, 32'h437b7533, 32'h43d6f5f8},
  {32'hc37022aa, 32'h42bb72ae, 32'h4397e5ed},
  {32'hc49f19a2, 32'h428289a6, 32'h421f51d2},
  {32'h44db6db1, 32'hc2112d78, 32'hc233d43f},
  {32'hc4c5d9c2, 32'hc31897a4, 32'hc253a167},
  {32'h44092eca, 32'hc3b2880f, 32'h43c53b8c},
  {32'hc4f82122, 32'hc2a5123f, 32'hc32d20ef},
  {32'h440a9b04, 32'hc24e01da, 32'hc315a696},
  {32'hc4a66164, 32'h430cd533, 32'hc2a09387},
  {32'h44c18df9, 32'h42a76597, 32'h43981eb7},
  {32'hc5087533, 32'hc1286e3e, 32'h42548347},
  {32'h44a01778, 32'h436e39d4, 32'hc232a54e},
  {32'hc4953bd2, 32'hc35b004e, 32'h42cf175b},
  {32'h446213b8, 32'h4266d9a3, 32'h41f18a36},
  {32'hc4990d71, 32'hc3aea223, 32'hc2b9748e},
  {32'h4491078e, 32'h43b4d89e, 32'hc3197e9e},
  {32'hc425f8dc, 32'h42086901, 32'h42f28ab1},
  {32'h445b0f7a, 32'hc2e31f22, 32'h42e4d79a},
  {32'hc31ee230, 32'hc3974482, 32'h438edaf9},
  {32'h44db9067, 32'hc38e907a, 32'h4349f4e3},
  {32'h448488b8, 32'h43b3ba34, 32'hc35e0ccc},
  {32'hc33309bc, 32'h430acf2c, 32'hc36c6d62},
  {32'h44974bc4, 32'hc32bf13a, 32'h428d442c},
  {32'h45190b06, 32'h42f4b220, 32'hc375d9aa},
  {32'hc4af7176, 32'h437a5429, 32'h433e859a},
  {32'h434abdfa, 32'h4391c19a, 32'hc2236f29},
  {32'hc4cd434c, 32'hc34dbe63, 32'h43438dee},
  {32'h4422e896, 32'hc3ba0eac, 32'hc301c628},
  {32'hc3cd0504, 32'h41a269fb, 32'h427617ca},
  {32'h4427ad38, 32'hc2dd0a1e, 32'hc089ad21},
  {32'hc3f646a0, 32'hc2b3522c, 32'h42bb1b11},
  {32'h44d77339, 32'hc35c11b9, 32'h429a0f46},
  {32'hc4cbf047, 32'h4027dd76, 32'h43198011},
  {32'h43bb33c8, 32'hc385e8c5, 32'hc1798879},
  {32'h430334d2, 32'hc395361e, 32'hc3621714},
  {32'h452c0884, 32'h4220f056, 32'hc3c7de50},
  {32'hc4a0f2fa, 32'h41d8a23d, 32'hc319f032},
  {32'h4484f746, 32'hc2ae77c4, 32'h42e7eb6f},
  {32'hc4ebf971, 32'h41d49ba3, 32'hc38ba752},
  {32'h4508bdd7, 32'h43356719, 32'h4326d00f},
  {32'hc50e5645, 32'hc3b8163e, 32'hc29f6889},
  {32'h44eba076, 32'h43346f55, 32'hc16ef157},
  {32'hc4983ccc, 32'h434777da, 32'hc326c0ee},
  {32'h44e38d79, 32'hc271e445, 32'hc2bf6fe4},
  {32'hc435d955, 32'hc21724b2, 32'hc36ceef9},
  {32'h43e25bf2, 32'hc2abc8d9, 32'hc2ee0e69},
  {32'hc3b4267a, 32'h43ac61c0, 32'hc38c6b40},
  {32'h446ae68f, 32'h4237938c, 32'hc361e0fc},
  {32'hc5105450, 32'hc2711942, 32'h4338ec68},
  {32'h4474bd48, 32'h440cadc4, 32'h41af46ac},
  {32'hc5159fd2, 32'h410fd2eb, 32'hc111f27d},
  {32'h445a3006, 32'hc3230b59, 32'hc3a1432f},
  {32'hc4ef3083, 32'h43d4b875, 32'hc1f30a3f},
  {32'h45010143, 32'h4387f306, 32'hc30dbf0d},
  {32'hc4911c93, 32'h420748aa, 32'h43750e27},
  {32'h410a2a00, 32'hc30514c7, 32'hc381a1c6},
  {32'hc4c741b7, 32'h43cb40b1, 32'hc1f7b8b1},
  {32'h435e3460, 32'hc34c0619, 32'h43ae7330},
  {32'hc4948dbe, 32'h43a7bbcb, 32'hc348f84b},
  {32'h451ed684, 32'h43654251, 32'hc3b0bcf2},
  {32'hc44de0d2, 32'hc1fc9814, 32'hc1ffee54},
  {32'h45115bff, 32'h424fdd0a, 32'hc0ee2840},
  {32'hc518d562, 32'hc3000faf, 32'h42d4f468},
  {32'h443466ed, 32'hc2271f1e, 32'hc0ca628b},
  {32'hc3e215f1, 32'hc24f5027, 32'hc3019990},
  {32'h44b611c7, 32'hc25e04bf, 32'hc32635c7},
  {32'hc4b0cc94, 32'h42c57768, 32'h440b8a99},
  {32'h43ce4c28, 32'h42ef7609, 32'hc2cf4e1a},
  {32'hc4b8e57e, 32'h43366822, 32'hc36ea038},
  {32'h4449eaec, 32'h438adc54, 32'h42352a74},
  {32'hc4560af2, 32'hc28e831d, 32'hc22b6919},
  {32'h44b24484, 32'hc30aa63c, 32'hc334b49e},
  {32'hc50207fc, 32'hc3957b4e, 32'h43b31327},
  {32'h4500d20e, 32'hc2fc6234, 32'h40aa8104},
  {32'hc50ae066, 32'hc3d8df39, 32'h440f2178},
  {32'h4471ba5e, 32'hc210722c, 32'h42d944f2},
  {32'hc4c8181e, 32'h43155bec, 32'h41e579b9},
  {32'hc4d6528d, 32'hc2c2ed09, 32'hc4209514},
  {32'h44904225, 32'h42bf25a4, 32'h41ea884d},
  {32'hc3f5e396, 32'h428c4b28, 32'h4383e1e7},
  {32'h44e92909, 32'hc1a5b116, 32'hc3d0d6b4},
  {32'hc526628f, 32'h4380eb6f, 32'hc3742c27},
  {32'h434cadbe, 32'h42c87738, 32'hc3815aec},
  {32'hc48ba27b, 32'h4332960e, 32'h410c0b21},
  {32'h451cebe5, 32'h431c29e8, 32'hbf0bd280},
  {32'hc41b753e, 32'hc23d01af, 32'h4412e6b8},
  {32'h451c954b, 32'h43528ef5, 32'h4352cd0b},
  {32'hc434e0d0, 32'hc306fde6, 32'h43cef728},
  {32'h44fbf383, 32'h429c268e, 32'h42190d66},
  {32'hc3fbc910, 32'hc106e418, 32'hc387f263},
  {32'h44c3c678, 32'hc2a36bca, 32'h42807dad},
  {32'hc4d45526, 32'hc2c20bf2, 32'h43696898},
  {32'h43d1070b, 32'hc21761f3, 32'h4246f9ed},
  {32'hc46446da, 32'hc2e4ec9f, 32'h40fbfcb5},
  {32'h44e8c935, 32'h43402412, 32'h4219cd5d},
  {32'hc49e2594, 32'h422fa69e, 32'h440fae68},
  {32'h44b25354, 32'h42f914df, 32'hc314909b},
  {32'hc4bae0b0, 32'h43303930, 32'h4386857a},
  {32'h43fd686c, 32'h43962bce, 32'h40abc821},
  {32'hc44c697b, 32'h4322bfe1, 32'h42eb720c},
  {32'h44aaedf6, 32'hc2b982b8, 32'h42e52810},
  {32'hc478da0b, 32'h40990e12, 32'h442d139b},
  {32'h436770e8, 32'h43da5744, 32'h4324d197},
  {32'hc45e5b8f, 32'hc42cde92, 32'hc37596d6},
  {32'h446b3f06, 32'h440efb57, 32'hc2534375},
  {32'hc39346fa, 32'hc377bf6d, 32'h4282a24f},
  {32'h4518fada, 32'hc3a88ac4, 32'hc2f079a7},
  {32'hc4b49c42, 32'h430bc609, 32'hc34d43ca},
  {32'h4505957f, 32'hc2b6deff, 32'h431bd1b2},
  {32'h4392dff8, 32'hc2ce6ad7, 32'hc3d40816},
  {32'hc3cae19c, 32'h43bb0f31, 32'h4318cc51},
  {32'h44116fac, 32'hc3bc6d83, 32'hc342cf9b},
  {32'hc4312c56, 32'hc3bbd657, 32'h44243693},
  {32'h44d1deeb, 32'hc31b01c8, 32'h4317af31},
  {32'hc33a756d, 32'h42ffba7d, 32'h436bac4c},
  {32'h4490095e, 32'h43a8aa64, 32'h40a1433f},
  {32'h4235db40, 32'hc27c8cfc, 32'h435863ec},
  {32'h44adb98c, 32'hc3990a62, 32'hc34e3ec3},
  {32'hc4a19dc2, 32'hc330b555, 32'hc258493b},
  {32'h4421c26f, 32'hc23c7152, 32'h4326f218},
  {32'hc2909424, 32'hc2d123f7, 32'hc339c9ce},
  {32'h442a1fba, 32'h42dfb360, 32'h42d840cb},
  {32'hc4c749b5, 32'hc2379236, 32'hc3d3dec8},
  {32'h44851ce2, 32'hc180c6f4, 32'hc2b4ea56},
  {32'hc45d9cdc, 32'h42a7c214, 32'h435d4528},
  {32'h43f8380b, 32'h43251367, 32'hc383e1f3},
  {32'hc3c9d48c, 32'hc2cc6d0b, 32'h4389f166},
  {32'h4502b3f5, 32'hc2c6afde, 32'hc19fd82d},
  {32'hc4bec38e, 32'h43fbdc2f, 32'h4247b989},
  {32'h44d9552a, 32'hc32b57a5, 32'h42a2556b},
  {32'hc449e6f1, 32'hc2db44b6, 32'h43373920},
  {32'h44d02951, 32'h4174c64a, 32'hc37cd687},
  {32'hc49b9984, 32'h4227b32f, 32'hc37147c8},
  {32'h44fdcf35, 32'hc31ae050, 32'h42bcb30d},
  {32'hc3f27370, 32'h43c26811, 32'h41a04c43},
  {32'h45081b5e, 32'h42e2828b, 32'h43241500},
  {32'hc4ee21eb, 32'hc3f5dc03, 32'hc2710bde},
  {32'h44f89e62, 32'hc34222bb, 32'hc2c4ec2c},
  {32'hc3f3ce1a, 32'hc369090c, 32'h42f9e80c},
  {32'h441a5370, 32'h438b98f6, 32'hc3b1a967},
  {32'hc40c7f98, 32'hc291b885, 32'h42993ce3},
  {32'h448db5c6, 32'hc3c5988a, 32'hc2a258f5},
  {32'hc5046cb4, 32'h436062cf, 32'h423e8a76},
  {32'h43bd8638, 32'hc3b17cae, 32'hc2309d2c},
  {32'hc5263dba, 32'hc3869921, 32'h435b9809},
  {32'h44d0cbff, 32'hc3b51bb6, 32'h43c7e3b3},
  {32'hc4900812, 32'h433eb618, 32'hc2fa5ecf},
  {32'h44b0f73a, 32'h433c68b1, 32'h43a71845},
  {32'hc415b0de, 32'h43b3b12a, 32'hc2067f4a},
  {32'h43715b68, 32'hc2aea562, 32'h418713f9},
  {32'hc4949e24, 32'h42622c18, 32'h43434c3e},
  {32'h44ad0baa, 32'hc3bd51fd, 32'h43484f8c},
  {32'hc5008219, 32'hc30edc35, 32'h42cd0c7b},
  {32'h449009f0, 32'hc2b65bc8, 32'h4349550a},
  {32'hc3ca8630, 32'hc32c9134, 32'h43bc7c33},
  {32'h45023b48, 32'h4315966e, 32'hc38a8472},
  {32'hc50d045f, 32'hc40ee2c2, 32'h4303793e},
  {32'h43c8c52c, 32'h4414a506, 32'hc26364c0},
  {32'hc49facf6, 32'hc384dfa5, 32'h41d2ccc0},
  {32'h450b8ddb, 32'h434caa07, 32'h4259561e},
  {32'hc43c78fb, 32'h426c4ceb, 32'h438d80ca},
  {32'hc415d140, 32'h42d74a46, 32'h4265a1b4},
  {32'h439e7f70, 32'hc31328fb, 32'hc32bb522},
  {32'hc4c1f07e, 32'h40e682b8, 32'h438a27fa},
  {32'h44a4a380, 32'hc3a08006, 32'h43474599},
  {32'hc4b3e9f0, 32'hc150737f, 32'hc3839444},
  {32'h4489f61b, 32'h43b01b81, 32'hc37487b1},
  {32'hc4f51584, 32'h4308b5b5, 32'hc2e6b93d},
  {32'h44d4a276, 32'h41a322c2, 32'hc1cb47fa},
  {32'hc4b32c4b, 32'h42ac56b4, 32'hc27450f2},
  {32'h44ad1c7e, 32'hc3d77015, 32'hc3290b79},
  {32'hc465b4a0, 32'h4393658a, 32'h4386c589},
  {32'h44ea92a8, 32'hc307bb65, 32'hc13a93d4},
  {32'hc4d1ec17, 32'hc26b4ad4, 32'hc34bbe7f},
  {32'h44ff9f82, 32'hc298bd73, 32'hc3b75307},
  {32'hc50e19f8, 32'hc3267cef, 32'hc28c423b},
  {32'h44e9d9c1, 32'h4205071b, 32'h43c243d2},
  {32'hc50fe662, 32'h4211bbb8, 32'h43d55aca},
  {32'h44dcfcb9, 32'h42022ae6, 32'h430dd7e0},
  {32'hc46ddfff, 32'hc38f97f7, 32'h42983e0f},
  {32'h4493ed39, 32'hc3bc1ca6, 32'h43ca473a},
  {32'hc4bd6321, 32'hc140917c, 32'h4373c05e},
  {32'h44995b9e, 32'hc2b8a965, 32'h43ea4b25},
  {32'hc4b47774, 32'h428e7e07, 32'hc3dc9339},
  {32'h45064c32, 32'h43a162b5, 32'h43c8c642},
  {32'hc490c62b, 32'h42f00a82, 32'hc341f2a8},
  {32'h44b93aa2, 32'h438556b1, 32'h42d4d30e},
  {32'hc49ffb2b, 32'h421face8, 32'h42fb8442},
  {32'h44f39c0a, 32'hc383982d, 32'h4394e664},
  {32'hc500763b, 32'hc2c3cde8, 32'hc225d41c},
  {32'h44e9085f, 32'h424b56d5, 32'h42a4d7c1},
  {32'hc4405edc, 32'hc33ef62c, 32'hc38dd917},
  {32'h4477118f, 32'h42451719, 32'h42e2df1d},
  {32'hc483d725, 32'h43811e4c, 32'hc38b0459},
  {32'h421b4090, 32'h43a21286, 32'h43d24847},
  {32'hc32ad168, 32'hc3737e06, 32'h424b37d3},
  {32'h441968ae, 32'h42929456, 32'h43cc1e1f},
  {32'hc3ffd194, 32'h429f4237, 32'hc3c03e60},
  {32'hc465a6f5, 32'h42e3a39c, 32'h421f747c},
  {32'h45270ef6, 32'hc3455cb9, 32'h42c22668},
  {32'hc4171132, 32'hc3630d0d, 32'hc3a2b129},
  {32'h44d20968, 32'hc3cb289d, 32'h422a5c24},
  {32'hc442b6ae, 32'hc3028b38, 32'h43039023},
  {32'h44c1d9e2, 32'hc33e474a, 32'hc382e914},
  {32'hc44a9f68, 32'hc3ce233e, 32'hc39a2629},
  {32'h43ad52d5, 32'hc35ae505, 32'hc306d823},
  {32'hc428099e, 32'hc386997c, 32'h436da57b},
  {32'h45155346, 32'h4295faa0, 32'hc3c3c188},
  {32'hc4e21fa2, 32'h4403b13c, 32'h43a3917d},
  {32'h451f94ce, 32'hc3adf9e1, 32'h4365882d},
  {32'hc38b7a5a, 32'h4162165d, 32'h42830ecf},
  {32'h447f51a3, 32'h42001f75, 32'h41588c9d},
  {32'hc3847e80, 32'hc1e718ad, 32'hc30d79ef},
  {32'h41ddc380, 32'hc333551b, 32'h4302284e},
  {32'hc4b279a7, 32'hc09cd3c0, 32'hc295213e},
  {32'h4494ee54, 32'h42e219f7, 32'h429e6f90},
  {32'hc400c5d0, 32'h440659cc, 32'h438600a8},
  {32'h43469668, 32'h434130fe, 32'h43580800},
  {32'hc4e6005c, 32'h4303d637, 32'h42d2faa9},
  {32'h44d8e86e, 32'hc3b6171f, 32'hc227eb9a},
  {32'hc3dbfc10, 32'h41f8e543, 32'hc2a1d335},
  {32'h449c9ead, 32'h4351ed67, 32'h4367cec0},
  {32'hc509e498, 32'h418feff1, 32'h4166f814},
  {32'h43f82221, 32'hc31977c1, 32'h4387556d},
  {32'hc4ee57b2, 32'h43e8b176, 32'hc25f2d02},
  {32'h43c7d216, 32'h437d57fd, 32'h434c50be},
  {32'hc509030d, 32'h42b19de1, 32'hc2b34c99},
  {32'h4252e300, 32'hc382eaf5, 32'h418d3a50},
  {32'hc44f722c, 32'h40dfcd68, 32'hc3b1cccf},
  {32'h43ee83a2, 32'hc0aeb587, 32'hc2f4ebb0},
  {32'hc4e32e44, 32'h43b9e73e, 32'hc15537f2},
  {32'h44b411a0, 32'hc37dad37, 32'hc2a079fd},
  {32'hc3f88f94, 32'h44094444, 32'hc2d737e7},
  {32'h449cc8b7, 32'h42ab272c, 32'hc2ac8f58},
  {32'hc3355998, 32'h42e88e7b, 32'hc2cf9620},
  {32'h43412e4e, 32'hc2ed9286, 32'hc31efc38},
  {32'hc5199e8b, 32'hc1726368, 32'h440f51b6},
  {32'h44de9d99, 32'hc2cb60b2, 32'h4307e566},
  {32'hc44cd394, 32'h4080d5aa, 32'h428cee5d},
  {32'h43b76b20, 32'hc2e9cf46, 32'h42b2cd0e},
  {32'hc509f01a, 32'hc2fe2bd6, 32'h43920e03},
  {32'h44054184, 32'h42a03293, 32'h431b17b7},
  {32'hc4cfb0e7, 32'h42bf5a26, 32'hc2b2a6a4},
  {32'h4488033d, 32'h42d55416, 32'h42d12d71},
  {32'hc3e89c31, 32'hc3a49a5c, 32'h431a92e7},
  {32'h451e3ecd, 32'hc38935df, 32'h439ec556},
  {32'h437836e6, 32'hc18b0c65, 32'hc2abf5cc},
  {32'h44c49440, 32'hc113e955, 32'hc2b74c81},
  {32'hc4fddddd, 32'h43a79729, 32'hc2c299b8},
  {32'h4399ddd4, 32'hc418fba6, 32'hc1ecbe8c},
  {32'hc4ead8c9, 32'hc2d9bf2b, 32'h431b4a6e},
  {32'h445f4f31, 32'hc37c3a0f, 32'hc27fbeea},
  {32'hc4166fff, 32'h4324dca7, 32'h4179aca2},
  {32'h4502863a, 32'hc129b0b8, 32'hc38928e2},
  {32'hc4e1d444, 32'h4334324d, 32'h436427d0},
  {32'h44e86a83, 32'h439b20ea, 32'hc3034789},
  {32'hc49046ae, 32'hc374b410, 32'h425f2054},
  {32'h43b46b41, 32'h4317c12e, 32'h42f87acc},
  {32'hc3bfc922, 32'h4232919e, 32'hc30f7739},
  {32'h44618d72, 32'h4280ca73, 32'hc290c0c0},
  {32'hc50c92c4, 32'h42654c47, 32'h41a2a533},
  {32'h44dac12d, 32'h43843e46, 32'h42024710},
  {32'hc46a6651, 32'h4358ac27, 32'hc393205c},
  {32'h4501accc, 32'h43a8518e, 32'h42e7cbdc},
  {32'hc50a5cb2, 32'h435f6ccb, 32'hc21426c2},
  {32'h4368c3f4, 32'h432ecb7b, 32'hc1a33e97},
  {32'hc485e08c, 32'hc3298e4b, 32'h42db2dea},
  {32'h44a6e81b, 32'hc2d7ab3c, 32'h43fa5acf},
  {32'hc310a77c, 32'hc2a91591, 32'h4282359c},
  {32'h448307a7, 32'hc2f0829d, 32'hc38df43f},
  {32'hc4ffdfec, 32'hc3274a84, 32'hc37efd14},
  {32'h44af63ab, 32'h40927607, 32'hc390b9aa},
  {32'hc4c79a30, 32'hc28c19ce, 32'hc1c4060c},
  {32'h4525babe, 32'hc1853a76, 32'h421bd500},
  {32'hc517d729, 32'hc1919e56, 32'hc34976f6},
  {32'h4467383c, 32'hc2f79b66, 32'h41bdd78c},
  {32'hc49dd7a9, 32'h4361b409, 32'h43641bf9},
  {32'h44a68ed5, 32'hc2a50ed6, 32'hc35ec47f},
  {32'hc49ed788, 32'h4080c202, 32'h436088f5},
  {32'h450dc5a0, 32'h431b5715, 32'hc33e2811},
  {32'hc465d298, 32'h43176ba9, 32'h43283f0e},
  {32'h45054743, 32'hc2fe4d03, 32'hc1405314},
  {32'hc5039a67, 32'h43881f6a, 32'hc3472c5f},
  {32'h4362c4fe, 32'h429962b7, 32'h423a3cbf},
  {32'hc4c70245, 32'hc378350f, 32'h436e4c2e},
  {32'h45081464, 32'hc34837fa, 32'hc2e6de10},
  {32'hc4dd9a9a, 32'h439f6a24, 32'hc3b46e29},
  {32'h42cd3aa0, 32'hc2c4f6e4, 32'h4202b74e},
  {32'hc42430bd, 32'h41c6324e, 32'hc351a4f5},
  {32'h45027129, 32'hc30fc557, 32'hc38264be},
  {32'hc3305ade, 32'h43bf5846, 32'h4161865c},
  {32'h44ec192f, 32'hc40923b9, 32'h420e76ac},
  {32'hc506081a, 32'hc2feae6c, 32'hc1ec1d2a},
  {32'h44f563d6, 32'h439f769a, 32'hc2433bd7},
  {32'hc3296170, 32'hc1c2e7c0, 32'h42a7f46e},
  {32'hc36fa4b0, 32'hc2f2e91e, 32'hc1252ae8},
  {32'hc5063a32, 32'h42cd5793, 32'hc2cfb1f6},
  {32'h44adeb0c, 32'h41c05641, 32'h4385d482},
  {32'hc41e2e62, 32'h42adb919, 32'h42862f96},
  {32'h450d8242, 32'h424cb826, 32'h43adfa99},
  {32'hc4598631, 32'hc3cab839, 32'h43a46a94},
  {32'h43422b44, 32'hc218983c, 32'h427c3ed3},
  {32'hc4ca5011, 32'hc3f627ce, 32'h420d0ebc},
  {32'h441d2d7a, 32'hc3fdaee9, 32'hc2c5ef67},
  {32'hc4ca25bc, 32'h41eda738, 32'hc2e31977},
  {32'h4494920a, 32'h42e2c26a, 32'h43597265},
  {32'hc385a1c0, 32'hc36990bd, 32'h427f0725},
  {32'h441ea7aa, 32'h432966c2, 32'hc2b5a68c},
  {32'hc455d4d6, 32'hc351897c, 32'h4371dd25},
  {32'h448637e5, 32'hc3810cdf, 32'h42dcf88e},
  {32'hc3572a8a, 32'hc321baa1, 32'h423d1a38},
  {32'h44c7f3a5, 32'hc4111248, 32'h43abf8c9},
  {32'hc4034109, 32'h43361379, 32'hc390102c},
  {32'h44d04a8f, 32'hc2bf87de, 32'h4229b68f},
  {32'hc49f8dd5, 32'hc29ecf2f, 32'hc33f4f4d},
  {32'h44ceee7c, 32'h42d3ba69, 32'h436404f5},
  {32'hc4df6fa4, 32'h40b46cf4, 32'hc385ca6c},
  {32'h44770ed2, 32'hc34f997d, 32'hc34faec7},
  {32'hc48b9ef7, 32'h42da1369, 32'h4329c85d},
  {32'hc4ea519a, 32'hc35900c0, 32'h4305cd15},
  {32'h44ee0e72, 32'h42bbfdea, 32'h43180a39},
  {32'hc4335418, 32'hc3050baa, 32'h43556719},
  {32'h44b7b1a0, 32'hc300b4b6, 32'hc39e7f10},
  {32'hc4896d3a, 32'hc209ee83, 32'h4397433e},
  {32'h44e21133, 32'h4307b212, 32'h429bc5ee},
  {32'hc45b02c6, 32'h440b6964, 32'hc24342a6},
  {32'h43d4e16a, 32'hc3a1a38a, 32'hc252fc06},
  {32'hc407745d, 32'hc1a0b14a, 32'hc293e6a0},
  {32'h44d9344c, 32'hc186e227, 32'hc2f839a8},
  {32'hc4ab05ac, 32'h433dc270, 32'hc20cba8c},
  {32'h44b2c54a, 32'h42eda1fb, 32'h43b90db4},
  {32'hc4a923ba, 32'hc22a9338, 32'hc1e37582},
  {32'h446d8b54, 32'h42fab4c6, 32'hc3561030},
  {32'hc3f8b166, 32'h4210a18f, 32'h438bb07d},
  {32'h43b0e4e2, 32'hc3b3d244, 32'hc0b3c3a1},
  {32'hc43c1f6b, 32'hc316d953, 32'hc35177ef},
  {32'h431950b0, 32'h43a87e45, 32'h43100a82},
  {32'hc48a8e29, 32'h41ca8811, 32'hc3312c73},
  {32'h43a5bd60, 32'hc3ba6e1a, 32'h42ce2dbc},
  {32'hc50e835c, 32'hc35e6a1b, 32'h42bfd5ae},
  {32'h43960500, 32'h438835ab, 32'h43706b8e},
  {32'hc4a9ed19, 32'h41b34898, 32'h43203ddd},
  {32'h444c999c, 32'h43a58f66, 32'hc31107f5},
  {32'hc505d8fe, 32'h429ad944, 32'h42261c7e},
  {32'hc514b92a, 32'hc2ba050c, 32'hc286fbb7},
  {32'h44eb7bf8, 32'h427fed74, 32'hc44217ae},
  {32'hc4a539fc, 32'hc27f84c4, 32'hc35d5496},
  {32'h44b4596a, 32'hc3b4f15d, 32'h42d0bbf2},
  {32'hc4dab99b, 32'hc39362c0, 32'h43944ea4},
  {32'h44ede2e2, 32'h42a4612a, 32'h42d58530},
  {32'hc3a0f87b, 32'h430aa103, 32'h433c8cea},
  {32'h44b531ee, 32'hc29dcbd0, 32'hbfb817d4},
  {32'hc4fc193b, 32'hc31603e1, 32'hc341b809},
  {32'h445c63b6, 32'h43bde481, 32'h440a7566},
  {32'hc51b9618, 32'hc32388a1, 32'hc3483722},
  {32'h44aa59a7, 32'h42807621, 32'hc2c55906},
  {32'hc4b9492d, 32'h4396df59, 32'hc33ff612},
  {32'h446737bc, 32'hc4068b80, 32'h422df1cf},
  {32'hc4c6b247, 32'h424eeeb6, 32'hc25552d4},
  {32'h43872c8b, 32'h42473734, 32'hc3307d28},
  {32'hc4abf9d3, 32'hc3b54057, 32'h43b0eaf2},
  {32'h43d11cf8, 32'hc3285c16, 32'h435da5eb},
  {32'hc4dd87ab, 32'h43132e48, 32'hc38adf16},
  {32'h44eae57e, 32'h432a1bf0, 32'h42598de5},
  {32'hc2fa5a78, 32'h43123d6a, 32'h43b9dfd2},
  {32'h441d57b2, 32'h42d7b8df, 32'h42b8d7e2},
  {32'h4361a7b0, 32'h4375dad6, 32'hc38391c4},
  {32'h44a3e69c, 32'hc262da20, 32'hc3a52a0a},
  {32'hc50c44e2, 32'h4362c051, 32'hc380bfd7},
  {32'h43df0c1f, 32'hc22e86fd, 32'hc23bd742},
  {32'h43a12c32, 32'h43aa6cde, 32'hc2796c4e},
  {32'h44d2bd6b, 32'hc308b103, 32'hc396b0be},
  {32'hc4148208, 32'h43525458, 32'h42d0b911},
  {32'h444c1e36, 32'h43f667e6, 32'h43221516},
  {32'hc4fd453c, 32'hc3035a73, 32'hc365b848},
  {32'h451433e2, 32'hc385058a, 32'hc34f1708},
  {32'hc49a105e, 32'h43f8482c, 32'h440878bb},
  {32'h438733d0, 32'h42987c34, 32'hc393db2f},
  {32'hc31ee310, 32'hc1141e0f, 32'hc31d6ccd},
  {32'h44c733a8, 32'h42e5d209, 32'h43d5c828},
  {32'h41d389c0, 32'hc3252b50, 32'h434a5681},
  {32'h44d6a1e7, 32'h438da008, 32'h433a9bd2},
  {32'hc51bbe12, 32'hc2af8561, 32'hc35a4b04},
  {32'hc4f16ede, 32'h43614890, 32'hc305d293},
  {32'h4513cd59, 32'h43f9f9cf, 32'hc318040e},
  {32'hc225b500, 32'h434085a6, 32'hc3daaa76},
  {32'h44a94da0, 32'hc38d653e, 32'hc28c179b},
  {32'hc3c9eeb6, 32'h43540aec, 32'hc19c0bfe},
  {32'h44907eaf, 32'h41c15837, 32'hc2bb4f42},
  {32'hc4927931, 32'h431354b0, 32'h41c59462},
  {32'h43a01274, 32'hc2a11a98, 32'h4334312f},
  {32'hc5006c14, 32'h42a3a7a4, 32'h42d680d8},
  {32'h444322d3, 32'hc34aabb9, 32'hc34a3dd7},
  {32'hc472e0e8, 32'hc007b60b, 32'hc1e063d5},
  {32'h4478e821, 32'h3f632339, 32'h433c3403},
  {32'hc4fae68c, 32'hc33cabf8, 32'hc34b53eb},
  {32'h44acd049, 32'hc2a8c88c, 32'hc2242431},
  {32'hc484ba48, 32'h417e180f, 32'h4295f85a},
  {32'h450f71d6, 32'h4212c913, 32'h43861354},
  {32'hc48525c9, 32'hc280f2cd, 32'h42a9213b},
  {32'h448d0290, 32'h42b2712c, 32'hc2504f8b},
  {32'hc3dd03ae, 32'h43e28ea2, 32'h42da0262},
  {32'h448c7225, 32'h435d7b4a, 32'h42e773ed},
  {32'hc4884a0f, 32'h43034d13, 32'h432ef232},
  {32'h44be9602, 32'h43996aa2, 32'h43558d4a},
  {32'hc435bbad, 32'h42a01526, 32'hc136fcbb},
  {32'h440eff69, 32'hc25d6135, 32'hc12eb7bc},
  {32'hc4092653, 32'hbe0cb548, 32'hc2836d80},
  {32'h4426850a, 32'h435eb0c8, 32'hc34a2015},
  {32'h425e66c0, 32'h42e64e2c, 32'hc1da29ba},
  {32'h4156d200, 32'hc250e8d2, 32'h420be06c},
  {32'hc401460e, 32'h436546f0, 32'h43b304de},
  {32'h43cf31a8, 32'h435ca75f, 32'h41114f85},
  {32'hc4560c5f, 32'h4245ceb2, 32'h434f26f0},
  {32'h444d70e4, 32'h428605c0, 32'h4334b0e0},
  {32'hc4145400, 32'hc3e269a7, 32'hc3190453},
  {32'h451fbca7, 32'hc1bb80d5, 32'h425b974a},
  {32'hc509757e, 32'hc2e1c515, 32'hc29c7828},
  {32'h44c740a0, 32'h43c1b3de, 32'h40c8e72c},
  {32'hc4ed3c51, 32'h43bb66ba, 32'hc367d9df},
  {32'h44b42b75, 32'hc3b6e87d, 32'hc38871be},
  {32'hc3c9a7f8, 32'hc3c32f53, 32'h42041a87},
  {32'h447e96ec, 32'hc3035759, 32'hc3ab76e7},
  {32'hc51416e1, 32'h43bd03de, 32'h439ea319},
  {32'h442ba332, 32'h42ffdd01, 32'hc247f51d},
  {32'hc4832782, 32'hc069fcc0, 32'h41cd4cde},
  {32'h45161ee4, 32'h427f991c, 32'hc37ef0f8},
  {32'hc4803b56, 32'hc2ad8115, 32'h434bad09},
  {32'h450e5a9c, 32'hc36672de, 32'h40d504dd},
  {32'hc2d59120, 32'hc3681c6a, 32'h4327267c},
  {32'h44dbf93d, 32'h431e8e41, 32'h41fa554a},
  {32'hc4d16934, 32'h420e377e, 32'h432507c2},
  {32'hc287ed04, 32'h4310941d, 32'h43606073},
  {32'h44317998, 32'h42744f1b, 32'hc362193f},
  {32'hc488e379, 32'h438ed90b, 32'h428ea29a},
  {32'h44ad9cca, 32'h42a7395f, 32'hc41fa8ee},
  {32'hc515b72c, 32'h4364ae29, 32'hc389a93c},
  {32'h451bdbb2, 32'h43574c37, 32'h43aa005c},
  {32'hc4db3cd9, 32'hc387f59c, 32'hc2c90a04},
  {32'h4511327d, 32'hc2f65b3a, 32'hc33ffda1},
  {32'hc4cb5a3f, 32'hc41ef30b, 32'hc1c9e96d},
  {32'hc1943040, 32'hc287c240, 32'hc26208f2},
  {32'hc4f4cca2, 32'hc2f436f1, 32'h411a58c9},
  {32'h446da092, 32'h42b1d505, 32'h437c5b2c},
  {32'hc49706c5, 32'hc2aef80b, 32'hc3836622},
  {32'hc38568de, 32'hc3ae3616, 32'hc239e07a},
  {32'hc42f7466, 32'hc203e527, 32'hc36e47c5},
  {32'h451e01fd, 32'h42467387, 32'hc404ef1d},
  {32'hc481efa0, 32'h43a61d79, 32'h421d8d90},
  {32'h44d3f228, 32'h4394dd7c, 32'hc358daf9},
  {32'hc49a8842, 32'h436e0d19, 32'h42c1daf6},
  {32'h4476207a, 32'hc3f1d536, 32'hc1314f34},
  {32'hc50974fe, 32'h42a01179, 32'hc36e3fa6},
  {32'hc39402d4, 32'hc2152564, 32'h4102cd97},
  {32'h44785ded, 32'hc29bf639, 32'h43bd567a},
  {32'hc4719110, 32'hc30b85fb, 32'h42a16ee8},
  {32'h45195965, 32'hc38372d2, 32'h42eb8164},
  {32'hc4991983, 32'hc29a9249, 32'hc3395aed},
  {32'h44e7942b, 32'h422c095b, 32'hc2a5ad93},
  {32'hc4d063bd, 32'h41580546, 32'hc2ba8327},
  {32'h4423ec8a, 32'hc1870b23, 32'h42617d20},
  {32'hc5176690, 32'hc40303b4, 32'hc3877d5e},
  {32'h44826d34, 32'h4247e404, 32'h42b3125a},
  {32'hc4589cd9, 32'h4311240d, 32'h435312d9},
  {32'h436df2d2, 32'hc2d53b77, 32'h431e279a},
  {32'hc3ee6794, 32'h4350c45f, 32'h3d355d00},
  {32'h448c6f95, 32'h42de6f96, 32'hc2e146e1},
  {32'hc3e874f0, 32'h435d6d16, 32'hc3b54fbf},
  {32'hc1b41070, 32'h435b2567, 32'hc2575cc5},
  {32'hc4382896, 32'h422e5b82, 32'hc3bc3902},
  {32'h441e8349, 32'h4342d0f4, 32'hc2a7131c},
  {32'hc4c2a220, 32'hc33323ff, 32'h43a990be},
  {32'h43bd2ab3, 32'hc3786c90, 32'hc2f55399},
  {32'hc4df3b3f, 32'hc265e09b, 32'hc3844368},
  {32'h4504323d, 32'hc2a3a1db, 32'hc395065c},
  {32'hc4dacc68, 32'hc28a0e02, 32'hc25266fa},
  {32'h4456cccc, 32'h41a3927c, 32'hc245ee1f},
  {32'hc474827f, 32'h4215cb99, 32'h42e232ef},
  {32'h441bc3b0, 32'hc3d4167c, 32'hc1dbc852},
  {32'hc5059d76, 32'hc33196b7, 32'hc3ff5a12},
  {32'h441420f6, 32'hc3a34cd4, 32'hc365798b},
  {32'h4306ffd0, 32'hc343cd87, 32'hc2c081e6},
  {32'h44d8684e, 32'hc208d33a, 32'hc157d242},
  {32'hc487a232, 32'h42bf7bed, 32'hc392dc23},
  {32'hc50aba8a, 32'h42af3ca2, 32'h434ddb45},
  {32'h43b1f6a4, 32'h426c776c, 32'h43cff48e},
  {32'hc4c21bf6, 32'h43af8996, 32'hc32a3c1e},
  {32'h44275ea0, 32'hc306e809, 32'h43a5847c},
  {32'hc4c7871c, 32'h43053d65, 32'h43a25f78},
  {32'h445599bb, 32'hc3185bb4, 32'hc198c353},
  {32'hc4f2131b, 32'hc30a3b3e, 32'hc3b78e32},
  {32'h4445cdee, 32'h436309c6, 32'h43b1d354},
  {32'hc500664d, 32'hc3246e18, 32'hc1e1c1ba},
  {32'h442d1fe6, 32'h421fc11b, 32'hc37626e1},
  {32'hc43d0efd, 32'hc3d49d5e, 32'hc2e2d7ab},
  {32'hc2448a60, 32'h4320a8f9, 32'hc21e4cee},
  {32'hc5067929, 32'h42dedfb9, 32'hc317bef2},
  {32'h44c26bcf, 32'hc2e14543, 32'hc2a931cc},
  {32'hc3c063e4, 32'h43da1e79, 32'h421a4548},
  {32'h4319dac0, 32'h42a01905, 32'hc31acae7},
  {32'hc4b840b6, 32'h4358ca16, 32'hc34a15bc},
  {32'hc5133835, 32'h4350627f, 32'h43255110},
  {32'h45013ab6, 32'h4418682c, 32'h43bee480},
  {32'hc41fb561, 32'h433b8254, 32'h41c1d60c},
  {32'h44e9766b, 32'h43053086, 32'h4302af8a},
  {32'hc4f46bef, 32'hc32c183b, 32'h42e7e2d6},
  {32'h44f00396, 32'h43ec9051, 32'h437d7452},
  {32'hc4bd8145, 32'hc341289d, 32'h433d8a58},
  {32'h44c9f346, 32'h42b09d0e, 32'h432d3a3e},
  {32'h43881c80, 32'h42767186, 32'hc22cb8f9},
  {32'h40fa3e00, 32'h432f1cd9, 32'h42a86e79},
  {32'hc467a1e4, 32'hc2966033, 32'hc31b2a4a},
  {32'h44f125d3, 32'h43a0705b, 32'h434d7a98},
  {32'hc5084149, 32'hc228e5fb, 32'h42af51d2},
  {32'h4484a6fc, 32'h43536d73, 32'h41253496},
  {32'hc3f18584, 32'hc26bc085, 32'h43c6e4a3},
  {32'hc4b151b0, 32'hc28f8009, 32'h42d71fbb},
  {32'h4444cb5c, 32'h415e89ff, 32'h43e87ffe},
  {32'hc504825a, 32'h434bc23d, 32'hc3a468c5},
  {32'h431a3980, 32'hc1a22dc6, 32'h43aabf1d},
  {32'hc4fee293, 32'h43c45c28, 32'hc38a534c},
  {32'h450475e7, 32'hc401cf79, 32'hc3b1b192},
  {32'hc4a0e591, 32'hc27426ae, 32'hc3e108c6},
  {32'h4504dc0a, 32'h436b49b3, 32'h436ca3e4},
  {32'hc4e6c4fb, 32'h4207150f, 32'hc34cc23e},
  {32'h44f53eb0, 32'h42ceb8d3, 32'h4373788e},
  {32'hc459f759, 32'h423bb2bc, 32'hc232079f},
  {32'h4488d773, 32'h4201daff, 32'h42a331c3},
  {32'hc2e4b070, 32'hc3f8bfa9, 32'hc3ce56bf},
  {32'hc2e8e2c2, 32'h431a9ca2, 32'h43087b59},
  {32'hc376aecc, 32'hc33966db, 32'h42090a1f},
  {32'h43b88c22, 32'hc3665d71, 32'h433f2b31},
  {32'hc4fb7de1, 32'h419bd873, 32'hc227b297},
  {32'h44b46bc2, 32'hc3305e2f, 32'hc18d5684},
  {32'hc50f4def, 32'hc2ad72be, 32'h40c43b08},
  {32'h43eab9f6, 32'hc2db58a5, 32'h4383746e},
  {32'hc43f139a, 32'hc339dc6f, 32'hc3ed86cd},
  {32'h444361cc, 32'h41a0a04f, 32'hc2e8d150},
  {32'hc43746e7, 32'hc2764d72, 32'hc344691c},
  {32'h44c26b16, 32'hc29cb9e7, 32'hc3277786},
  {32'hc4a924c4, 32'hc298e62f, 32'hc3a550ce},
  {32'h45037a2c, 32'hc3fa34f8, 32'h433d0967},
  {32'hc4b3494b, 32'h43580c0c, 32'hc30da3b9},
  {32'h44cb0933, 32'h4306bfe4, 32'h43fc1fc6},
  {32'hc4ee9ed4, 32'hc33ec8d9, 32'h4304ddaf},
  {32'h44194a2c, 32'hc362f17a, 32'h43649e26},
  {32'h42df56c0, 32'hc3a937bb, 32'hc1b2e8a5},
  {32'h448994de, 32'h4309ed48, 32'h4318f0cc},
  {32'hc39287fc, 32'h439a5b70, 32'hc3c52b87},
  {32'hc454aa12, 32'h43a3c6c8, 32'hc2bbae51},
  {32'h44b421cb, 32'hc2df062d, 32'h428ede8b},
  {32'hc4d0be05, 32'hc378ad82, 32'hc35c640d},
  {32'h439353b0, 32'h4180a72c, 32'h4258a92a},
  {32'hc4c1594e, 32'hc230034f, 32'h42ec15a6},
  {32'h44c954fb, 32'hbfb6cba8, 32'hc37616b8},
  {32'hc5071f3d, 32'h4379101e, 32'h418097c6},
  {32'h44a391c0, 32'hc34f07f0, 32'hc30d0c90},
  {32'hc481669b, 32'h41233a32, 32'hc40ca8ff},
  {32'hc4c3fbf5, 32'h434f8bf7, 32'hc396bdd9},
  {32'h44cce73f, 32'h42afa174, 32'hc28e71e5},
  {32'hc49bc589, 32'hc2b09843, 32'hc39a9026},
  {32'h43b5a3f0, 32'h437b70e2, 32'h4382362a},
  {32'hc3eb8bc0, 32'hc3a66c66, 32'hc332b12b},
  {32'h443adcc1, 32'hc3417f9f, 32'h415dc295},
  {32'hc4fb5ea6, 32'hc350aa4c, 32'hc3bc1edb},
  {32'h448c3693, 32'h430b4e3e, 32'hc3ec589c},
  {32'hc4ef0e04, 32'h422105e6, 32'h439503ed},
  {32'h44393053, 32'h4271409a, 32'hc3211bbf},
  {32'hc4c50cca, 32'h41cb7ca0, 32'h421cdb20},
  {32'h43ecf071, 32'hc271e390, 32'h430e1622},
  {32'hc50890b2, 32'h42891aa4, 32'h4330795e},
  {32'h44f898b8, 32'hc36a0223, 32'hc1bf5ccf},
  {32'hc4aa9ba8, 32'hc1e24b52, 32'hc2f37a2c},
  {32'h45090fac, 32'hc3148dba, 32'hc234a88a},
  {32'hc493dd3a, 32'hc2415a36, 32'hc39193b4},
  {32'h42eab608, 32'hc353f545, 32'hc1c11f1c},
  {32'hc424fd35, 32'hc27ded3b, 32'hc33fe5e7},
  {32'h44c907e7, 32'h43bc4825, 32'hc1b75434},
  {32'hc50451f2, 32'hc382a64b, 32'h42cfeb5b},
  {32'hc2d307d0, 32'hc32ea022, 32'h4384976a},
  {32'hc4ea38da, 32'h4332789c, 32'hc372edd2},
  {32'h4501ce72, 32'hc3b24c16, 32'hc375d051},
  {32'hc4d2f5c2, 32'h43827d8c, 32'hc3b092cd},
  {32'h44a58aa1, 32'hbfaf9a14, 32'h422d7a19},
  {32'hc4fb5ee2, 32'h43951c4b, 32'h41bb9300},
  {32'h450cd238, 32'hc2889923, 32'hc3adf97a},
  {32'hc50ad269, 32'hc2fe71da, 32'hc2bed4ee},
  {32'h440d3d3c, 32'h43fb9f34, 32'h40aeab1b},
  {32'hc5146b9f, 32'hc0f5e092, 32'hc2cf9cde},
  {32'h444dfeb8, 32'h428a0459, 32'hc27c4f68},
  {32'hc4e5cffa, 32'hc3ab2d31, 32'hc3bbe05f},
  {32'h44d6d624, 32'h42b8cb44, 32'hc39aa108},
  {32'hc4cb27d4, 32'h42e8762b, 32'hc3413124},
  {32'h44cb401c, 32'h43cf22f7, 32'h4401b992},
  {32'hc338e9ec, 32'h42949863, 32'hc297b3e6},
  {32'h44b3e560, 32'hc2bec04e, 32'h434104c1},
  {32'hc5059e61, 32'hc330f289, 32'hc3ba8b14},
  {32'h44995834, 32'hc36852a6, 32'hc3a838d4},
  {32'hc4ee059c, 32'h42442424, 32'h425e3980},
  {32'h446fbc7e, 32'hc3024603, 32'hc2b88f5d},
  {32'hc40d017d, 32'hc40a48c7, 32'h4400e107},
  {32'h45067a72, 32'hc2b134ce, 32'hc2a76346},
  {32'hc511c8a5, 32'hc2914e3e, 32'h43464e24},
  {32'h449fb9cc, 32'h4325948f, 32'hc307e8cc},
  {32'hc5162786, 32'hc28081ae, 32'hc3b58407},
  {32'h448f43fb, 32'hc2b04faa, 32'h410faf5c},
  {32'h41efd600, 32'h434b88dc, 32'hc2e7d8c5},
  {32'h443becea, 32'h424e687e, 32'h432b2b1e},
  {32'hc50db0cb, 32'hc3c84728, 32'hc1fb9b8c},
  {32'hc1e05e74, 32'h42d61edb, 32'h426230fd},
  {32'h448f5878, 32'hc256f3ed, 32'h4311cbc5},
  {32'hc4599943, 32'h42dc5f08, 32'hc387560f},
  {32'hc283a010, 32'hc2c0e3a6, 32'h44215416},
  {32'hc4b4ebb4, 32'h422250b1, 32'h438a9adf},
  {32'h44ca5b7e, 32'h42951a79, 32'hc38b0b31},
  {32'hc4f76f72, 32'hc18451a4, 32'h40945316},
  {32'h44b6afae, 32'hc38ffb00, 32'h42df5bf9},
  {32'hc5106334, 32'h43000bef, 32'h42d37fee},
  {32'h449321b6, 32'h42326ae5, 32'hc2981442},
  {32'hc386d360, 32'h4130b5ab, 32'h4121185d},
  {32'h43b7eeb0, 32'h4292b55f, 32'hc38b6db1},
  {32'hc485fad5, 32'h43672441, 32'h439396a5},
  {32'h44b2d88d, 32'hc2cd8a25, 32'hc384c8ee},
  {32'hc4f9060f, 32'h435f1743, 32'hc0860dec},
  {32'h42a6cb60, 32'hc2780020, 32'h41ae3b33},
  {32'hc42625c2, 32'h4359b49e, 32'hc299fac2},
  {32'h44f8efb7, 32'hc40b3a4b, 32'hc28ebbf3},
  {32'hc50288bb, 32'hc2715fc9, 32'h43bb91a9},
  {32'h4437161b, 32'h437c6a6c, 32'hc2af0b4a},
  {32'hc4970f17, 32'hc2b2fc41, 32'hc2b27ad6},
  {32'h451b8878, 32'hc30da43c, 32'h439e3153},
  {32'hc4ccdc75, 32'h4387bab0, 32'h430c828e},
  {32'h44c31c87, 32'hc356e493, 32'h43a47fc6},
  {32'h44194cc4, 32'hc3ca7e2c, 32'h437fe6cb},
  {32'hc515a604, 32'h4292cda1, 32'h42d18453},
  {32'h443853a0, 32'h43e7f199, 32'h40dbb870},
  {32'hc447c1ac, 32'hc2383015, 32'h42b36744},
  {32'h44a52cd3, 32'h43ac22b5, 32'hc34bdbc6},
  {32'hc385af8a, 32'h438023cb, 32'h42cf291a},
  {32'h4160a680, 32'h4393e702, 32'h435d719c},
  {32'hbfded800, 32'h43960d0f, 32'hc07b38d4},
  {32'h44bd9d84, 32'hc1d61d0f, 32'hc2cb3259},
  {32'h4357a57d, 32'hc295df98, 32'h43763164},
  {32'hc4762d10, 32'h4336c428, 32'h43027cf5},
  {32'h4422456b, 32'h43e64472, 32'h42dff9c4},
  {32'hc49171e8, 32'h42ba6c6b, 32'hc3095d0e},
  {32'h450914eb, 32'hc381b369, 32'hc2e41d6e},
  {32'hc43596c8, 32'hc25dc0d8, 32'h4319d597},
  {32'h43681760, 32'hc32358f9, 32'hc2a297f3},
  {32'hc4c134e8, 32'hc3495df4, 32'h429a7c06},
  {32'h430498c0, 32'h43d6625c, 32'h4366f3cb},
  {32'hc382ef80, 32'hc2d238a2, 32'hc31254bc},
  {32'h4502ea57, 32'h438fbce0, 32'h42aa4786},
  {32'hc47aca9e, 32'hc292160a, 32'hc23b434e},
  {32'h4508c4f2, 32'h421e788a, 32'hc3af9c03},
  {32'hc4865170, 32'h43f05a49, 32'h420e7b50},
  {32'h44abe88b, 32'h419409f3, 32'h42ab4b05},
  {32'hc4b15787, 32'hc290dca2, 32'hc2eeb6e5},
  {32'h43ab381d, 32'hc3ab7f1a, 32'hc1d8b84e},
  {32'hc47f6f66, 32'h42099246, 32'h436f0507},
  {32'h441c33d9, 32'h4316537e, 32'h41a51a8b},
  {32'hc4a10443, 32'h438e0130, 32'h4346eaa8},
  {32'h43c47f8c, 32'h4336af25, 32'hc38a4bbb},
  {32'hc08f5e50, 32'h441a3201, 32'h431f7008},
  {32'h42af962e, 32'h43bb20de, 32'h42024537},
  {32'hc3287161, 32'h426faef2, 32'h4303b4e0},
  {32'h44397d0e, 32'hc34a9f53, 32'h431a860f},
  {32'hc4e27fc8, 32'h40f77ad7, 32'h43470b6c},
  {32'h44cc5d67, 32'h42d06d62, 32'h4315dd3a},
  {32'hc4e29b6c, 32'h41380728, 32'h432891f2},
  {32'h43da1198, 32'hc27922f4, 32'hc3c85174},
  {32'hc421aaa1, 32'h4432597b, 32'h4239e7f7},
  {32'h447737f6, 32'h440808a3, 32'hc41cacd1},
  {32'hc4eb3398, 32'h415f44c6, 32'hc1be599a},
  {32'h4506d9ef, 32'hc27ce184, 32'hc2b1a199},
  {32'hc42420be, 32'hc35b226b, 32'hc3579150},
  {32'h448f96e5, 32'h43592fe5, 32'h43c33f45},
  {32'hc4b4d728, 32'hc3937f20, 32'h41ea1a7e},
  {32'h448c61e9, 32'h438a1968, 32'hc21267f6},
  {32'hc43130b8, 32'hc3236036, 32'hc32d076d},
  {32'h44ad0d5d, 32'hc35ef6b3, 32'hc30c39c9},
  {32'hc47fcf5b, 32'h41ad69cd, 32'h41c7c030},
  {32'h44c4a96b, 32'hc120943c, 32'hc333533f},
  {32'hc49056ed, 32'hc3897fbd, 32'h434d233a},
  {32'h446e6ca6, 32'h43886c1e, 32'h43bedc03},
  {32'hc20d9398, 32'hc26c0198, 32'hc3871dd5},
  {32'h44c47bf8, 32'h4310a85f, 32'hc3751506},
  {32'hc507b8f8, 32'h4389b6a6, 32'hc3a50b69},
  {32'h4434c0dd, 32'h41d715da, 32'h436a851a},
  {32'hc4ccf13c, 32'hc20c8694, 32'h41e051f1},
  {32'h44c001e3, 32'hc332303f, 32'hc328f3d0},
  {32'hc4fc4232, 32'h43a14816, 32'h438c758f},
  {32'h44c077ec, 32'hc3d147aa, 32'hc39c1e0c},
  {32'hc3e77364, 32'hc32d4d78, 32'hc39a0739},
  {32'h44b5303d, 32'hc3bdf076, 32'h440f065f},
  {32'hc4d499ab, 32'hc3c83104, 32'h419c752f},
  {32'h44a51510, 32'h43bd0244, 32'h43ac83ee},
  {32'hc37d4fd8, 32'hc2a8ceec, 32'h439f40a9},
  {32'h4438f7d4, 32'hc2ab2794, 32'hc3ae7b51},
  {32'hc4a4627f, 32'hc2d6fae4, 32'hc21948b4},
  {32'h45011ded, 32'hc32ed6b4, 32'h43b9a2cb},
  {32'hc390553a, 32'hc1ec066b, 32'hc30f530e},
  {32'h44fc00ee, 32'h422d0d99, 32'hc2c48a25},
  {32'h439a6a31, 32'hc3bf6fb9, 32'h43bc9032},
  {32'h44d9acbc, 32'hc29e4a1b, 32'h411c6f56},
  {32'hc42f4544, 32'h436ac60a, 32'hc3172950},
  {32'h448d43d6, 32'hc33cf7f6, 32'hc2ec9677},
  {32'hc3c24ea8, 32'hc2d8d53e, 32'h433ccfde},
  {32'h4520d442, 32'h432c5637, 32'hc32993d0},
  {32'hc4eec4cc, 32'hc38ffb97, 32'h42d98eee},
  {32'h446b3684, 32'h432f3abd, 32'h43d16b99},
  {32'hc4edeb65, 32'hc3af3f66, 32'h4353ff77},
  {32'h444e6f30, 32'h43259909, 32'hc315f7f0},
  {32'hc5004db3, 32'hc335ea68, 32'h438d8ba6},
  {32'h4490ba50, 32'h4265d715, 32'hc33329a8},
  {32'hc41dbf3a, 32'h43358388, 32'h43d1bd01},
  {32'h44ee0d51, 32'hc2e6bdb1, 32'h439bb767},
  {32'hc434d370, 32'h41b46e15, 32'hc323fca7},
  {32'h44e41d44, 32'h431e21ea, 32'h42d9a48c},
  {32'hc4a2c00d, 32'hc2cb487a, 32'h43046a27},
  {32'h450caf60, 32'hc3d0bf8e, 32'h4276558a},
  {32'hc3e7fac8, 32'h43953b3e, 32'h43e10a66},
  {32'h4513deaa, 32'hc2b3f5e0, 32'h3f74c300},
  {32'hc33d4300, 32'hc30db1d0, 32'h43962091},
  {32'h43605ab4, 32'h425284a7, 32'h439d972a},
  {32'hc443dfc6, 32'hc3f392b3, 32'h42ed704b},
  {32'h43a1427c, 32'hc301f723, 32'h441a6e9f},
  {32'hc3d90e2f, 32'h43a76ea3, 32'hc36301cb},
  {32'h438478c0, 32'h41a4f6bd, 32'hc35c8fb7},
  {32'hc4f6c52c, 32'h43b40964, 32'h43512ebd},
  {32'h44cea06b, 32'h403d0be2, 32'h42f5c29a},
  {32'hc4fbdbf8, 32'hc3acd76a, 32'h436f7dc0},
  {32'h43d6f2cb, 32'hc363571b, 32'h43524c37},
  {32'hc4b9dd02, 32'h4282cf2e, 32'hc34bbaa1},
  {32'h44a4b038, 32'h43dff80c, 32'hc2d65f7e},
  {32'hc4b9cdc7, 32'hc21758cc, 32'h419ba03c},
  {32'h43c71bb4, 32'hc483e09d, 32'hc36ba6b0},
  {32'hc509aade, 32'h4196eddb, 32'h42a2a01c},
  {32'h449afa59, 32'hc39095a1, 32'hc0322444},
  {32'hc504b526, 32'h431b23b1, 32'h44077634},
  {32'h433ce03e, 32'h4357b352, 32'h43871b2e},
  {32'hc50caed0, 32'hc2ea4503, 32'hc30b7ce3},
  {32'h44e160b2, 32'h42f5a652, 32'h42369742},
  {32'hc393e895, 32'hc2cca223, 32'hc23646a5},
  {32'h44108ef1, 32'hc32c2014, 32'hc32087a4},
  {32'hc41a55f6, 32'h4302bc2e, 32'hc3ae0889},
  {32'h42829ed0, 32'h43561998, 32'h43c22820},
  {32'hc2a2fa68, 32'hc296afb9, 32'hc2efc17e},
  {32'h44579224, 32'h4388e8a5, 32'h415dfcfe},
  {32'hc402189e, 32'h4383a1ef, 32'hc2713160},
  {32'h45085e1c, 32'h41b438b1, 32'hc3c0ecac},
  {32'hc4f12275, 32'h43d078d2, 32'hc2193043},
  {32'h45083361, 32'h4310a537, 32'h4380478a},
  {32'hc47e5040, 32'hc39d1677, 32'h43bd6b75},
  {32'h44d72ecb, 32'h42fac6c0, 32'h4170ad41},
  {32'hc40ae58e, 32'hc22804e8, 32'h43a0c84b},
  {32'h44b44638, 32'h42832019, 32'hc1854e06},
  {32'h42a2c213, 32'hc318a102, 32'hc29d579b},
  {32'h44493486, 32'hc1b29b86, 32'hc3736d1d},
  {32'h43219245, 32'h43a5f949, 32'h42a3517e},
  {32'h44be27ed, 32'hc45a7196, 32'h4399c2df},
  {32'hc414b3aa, 32'hc396b11a, 32'h4396783b},
  {32'h44947fd8, 32'hc3d8f0f5, 32'h435d3337},
  {32'hc4d628c1, 32'h42cfb81f, 32'hc31491eb},
  {32'h450f62d8, 32'hc387854a, 32'h4324f677},
  {32'hc49818b9, 32'h425cc990, 32'hc29065f8},
  {32'h447e9540, 32'hc2ff3311, 32'hc326a00f},
  {32'hc4a51bca, 32'hc34bec7a, 32'h43d8c27b},
  {32'h43f9b27c, 32'hc33b2f81, 32'h437f55a2},
  {32'hc4f17fd6, 32'h432916a1, 32'h437b2656},
  {32'h44ab8e67, 32'h43431e5e, 32'h428f1c18},
  {32'hc5012874, 32'h4208870b, 32'hc1461d56},
  {32'h45026462, 32'h41db49e8, 32'h4096543d},
  {32'hc5046a21, 32'hc358f479, 32'hc2945d58},
  {32'h448d85a2, 32'hc2b77a11, 32'hc30b9c21},
  {32'hc43bbb45, 32'h4310c742, 32'hc305535b},
  {32'h44b2043d, 32'hc3bc5173, 32'h422bfdb2},
  {32'hc438e4d8, 32'hc342e22f, 32'h436f48dd},
  {32'h44130fd4, 32'hc38eadd1, 32'hc360cb85},
  {32'hc50e60e8, 32'h42eb0e04, 32'h43454bcb},
  {32'h44d0dc51, 32'hc257e1e1, 32'h42419f77},
  {32'hc4a04fc2, 32'h43538a38, 32'hc3acfda1},
  {32'h450308f8, 32'h41a81072, 32'hc3a670fe},
  {32'hc4586276, 32'h428d9205, 32'hc38601ab},
  {32'h44ad00b3, 32'hc2fd2614, 32'h4389cf8c},
  {32'hc427d6c4, 32'hc1a4ec50, 32'hc3249e72},
  {32'h4494b9a5, 32'hc29023aa, 32'hc3ad469c},
  {32'hc5101433, 32'h43efc98e, 32'hc1d00b22},
  {32'h447e5488, 32'h3fcf0bf0, 32'hc3a93c29},
  {32'hc4adb925, 32'h430efc8e, 32'hc366bbe8},
  {32'h43d7fd10, 32'hc196465a, 32'hc3829340},
  {32'hc4662050, 32'h41b91f34, 32'hc3a9ab96},
  {32'h44d50b7e, 32'h439aa823, 32'h43a98e1f},
  {32'hc41e4534, 32'h43ac3e9e, 32'hc3fef582},
  {32'h43cc5f84, 32'hc307ebd0, 32'h43c2b6a8},
  {32'hc5034cd8, 32'h43cb6e74, 32'h42045eff},
  {32'h44fd8f26, 32'hc38c6fa4, 32'hc327b5be},
  {32'hc4e45071, 32'hc322c5c9, 32'hc358bfef},
  {32'h4486380f, 32'h4377ff67, 32'hc2b60bec},
  {32'hc481e082, 32'hc3590c6e, 32'hc2d65afe},
  {32'h44cfe184, 32'hc37162aa, 32'hc3ae5cd9},
  {32'hc51b42c0, 32'hc229f41f, 32'h4351394c},
  {32'h44b8df66, 32'h43458e8e, 32'h437077a0},
  {32'hc4b9ed10, 32'hc2367270, 32'hc429834e},
  {32'h44c16c95, 32'hc2901097, 32'h431d865f},
  {32'hc508c0fe, 32'hc2731e0a, 32'h439dcbf8},
  {32'h451b5c42, 32'h4259ad03, 32'hc3b14a75},
  {32'hc38218a0, 32'h434604b6, 32'hc2471a96},
  {32'h4504ffac, 32'h41355227, 32'h424c10b9},
  {32'hc4456037, 32'h43d6437f, 32'hc2a63089},
  {32'h436563a8, 32'hc24b6966, 32'h42263b9f},
  {32'hc3ff170b, 32'h426e22b4, 32'h4381b1aa},
  {32'h443327d4, 32'h43131eb9, 32'hc2515ad3},
  {32'hc4a81c59, 32'hc3be011a, 32'h4280520b},
  {32'h44f7050f, 32'h42e896af, 32'h438ac72d},
  {32'hc48cf0a1, 32'h42faed74, 32'hc3579297},
  {32'h44155d9f, 32'hc2525442, 32'hc0cacb23},
  {32'hc4fb9bd5, 32'hc2fe7c71, 32'hc22b21b6},
  {32'h435e24a0, 32'hc3a923d7, 32'hc33fb35c},
  {32'hc510079b, 32'h42348bbb, 32'h42d64bfd},
  {32'h4445f242, 32'hc0d53887, 32'h42d1d8e9},
  {32'hc51434ae, 32'h433dee6f, 32'h41ff046d},
  {32'hc50b3ce2, 32'h4300e248, 32'h4381012b},
  {32'h44dc5317, 32'hc32a5e22, 32'h431131c5},
  {32'hc4a74880, 32'h43640a32, 32'hc351c3fc},
  {32'h42a3fe54, 32'hc3ce7f1d, 32'h43fd2871},
  {32'hc482353a, 32'hc29d01ac, 32'h421e690f},
  {32'h44b9a44e, 32'h43121657, 32'hbfb4526e},
  {32'h4264ae40, 32'h431ce8e0, 32'h4389be24},
  {32'h440c85a4, 32'h44171f6b, 32'hc3b644e9},
  {32'hc4c7011a, 32'hc42b2455, 32'hc2b87e8a},
  {32'h44e6922f, 32'hc1a9f3a0, 32'h42a5504d},
  {32'hc4fdc722, 32'hc371a303, 32'hc18b78bc},
  {32'h451f7fb8, 32'hc2f3f818, 32'h44049929},
  {32'hc50c8e7b, 32'h432cc31f, 32'h42c55e32},
  {32'hc4936aca, 32'h433b7140, 32'hc381ae07},
  {32'h450174d1, 32'h42be9161, 32'h43d15818},
  {32'hc506bcb9, 32'h4395bd2e, 32'hc31718e4},
  {32'h4410676c, 32'hc376fc93, 32'hc34af0ec},
  {32'hc50f75d2, 32'h432e24f8, 32'hc3ca13a7},
  {32'h4489eac9, 32'h4299624f, 32'hc33ac724},
  {32'hc4d603b1, 32'hc3ac9e87, 32'h41c12204},
  {32'h448b18d5, 32'hc33d06b9, 32'hc358a95d},
  {32'hc48778d4, 32'h43987c72, 32'h418713da},
  {32'h445b884c, 32'hc4076b68, 32'h42e3a453},
  {32'hc49e71c6, 32'h43058d8d, 32'hc39fbcb4},
  {32'h44d04457, 32'hc2fa2975, 32'h438c06af},
  {32'hc47766ac, 32'hc3327f83, 32'hc39d0fc5},
  {32'h449f8d8c, 32'hc2eeffae, 32'h43408024},
  {32'h44c3778f, 32'hc2981ca3, 32'h43a9f042},
  {32'hc33c9240, 32'hc340e914, 32'h43d92404},
  {32'h442c1b7c, 32'h43446f2f, 32'h42aeee2e},
  {32'hc44c3c04, 32'hc31e2772, 32'h430317e0},
  {32'h44f407c0, 32'h43678da1, 32'h43c8ac3c},
  {32'hc40e83c6, 32'h41e75e6b, 32'hc2832424},
  {32'h43bec340, 32'h43842793, 32'hc3173a07},
  {32'hc50be55a, 32'hc3539528, 32'hc323f6f5},
  {32'h44f45469, 32'hc341c32d, 32'hc0cc86fb},
  {32'hc4187f59, 32'hc32eab1f, 32'h411316db},
  {32'h44c718c9, 32'h4419094b, 32'hc1b9a9ec},
  {32'hc21d1830, 32'h4300b4dd, 32'hc35d3ee7},
  {32'h4473b9fe, 32'h430e46d2, 32'hc25d2e3b},
  {32'hc454b81e, 32'hc2e8f854, 32'h4186be3d},
  {32'h45068a88, 32'h43906e92, 32'h42c19126},
  {32'hc4ae1ff5, 32'hc3212b74, 32'h40a4cd77},
  {32'h45004be8, 32'hc3039187, 32'hc2c18570},
  {32'hc3bb5cf1, 32'hc39f681f, 32'h42e6a6a3},
  {32'h4531f286, 32'h432a8101, 32'hc37d10e7},
  {32'hc358d528, 32'hc15732cb, 32'hc31d1e09},
  {32'h44ec2a00, 32'h429d50f0, 32'hc2b2afdf},
  {32'hc3ce2044, 32'h424fb30e, 32'hc2ca9720},
  {32'h451143e8, 32'hc38fcea9, 32'hc3332b62},
  {32'hc515cc3c, 32'h410bcbde, 32'h43cbae79},
  {32'h44be00ab, 32'hc2f06bf8, 32'h43330d3c},
  {32'h43aa6463, 32'h4374e193, 32'hc29bb2ac},
  {32'h44c39b6f, 32'hc26cb949, 32'h439d88ed},
  {32'hc49e8d52, 32'hc331405e, 32'hc239e77a},
  {32'h441c7168, 32'hc2aed818, 32'hc3c248f3},
  {32'hc50460d9, 32'h41d79b89, 32'hc10e3a58},
  {32'h4460ca52, 32'hc248bc22, 32'h408cd6a6},
  {32'hc493d87b, 32'hc18c569e, 32'h43a0df35},
  {32'h43ef1f7c, 32'hc2a38195, 32'h42ca4269},
  {32'hc4d2c905, 32'hc2d999d0, 32'hc1d62897},
  {32'h441ca0c6, 32'hc2d1abe7, 32'hc2717dc1},
  {32'hc50daa3d, 32'hc28cd79b, 32'hc2f37212},
  {32'h44ab0e63, 32'hc4282c3d, 32'h408c37d4},
  {32'h43008fca, 32'hc1d56644, 32'hc38db90f},
  {32'h449078f3, 32'hc2b76672, 32'hc252de23},
  {32'hc4b4dc1a, 32'hc384a678, 32'h438b6505},
  {32'h44d31742, 32'hc2b72e74, 32'h42fe902e},
  {32'hc3fd9aa4, 32'h431b4c62, 32'h434f073c},
  {32'h44fdba83, 32'hc359758b, 32'h4274e1f2},
  {32'hc4eb2638, 32'hc2c0559d, 32'h42dce400},
  {32'h43e6437b, 32'h436cefba, 32'h42ae675d},
  {32'hc42be6a8, 32'hc35cfc19, 32'hc3bd8246},
  {32'h45179f54, 32'h40f9afd8, 32'h42ab3e56},
  {32'hc50b2923, 32'h4335ec4a, 32'hc1b5c73a},
  {32'h449d5805, 32'hc1a9df7c, 32'h435c2949},
  {32'hc3caef88, 32'hc39d9dcf, 32'h433ee186},
  {32'hc530312e, 32'hc2150d2e, 32'h43a4940b},
  {32'h44d9556e, 32'hc37f6e64, 32'hc08f5617},
  {32'hc47983a6, 32'hc303fb2a, 32'hc3bd863f},
  {32'h44a69889, 32'h4389acfb, 32'h432a17ef},
  {32'hc20df839, 32'h43bbe96d, 32'h4121dae6},
  {32'h44bba6c7, 32'h419611f3, 32'hc32e6152},
  {32'hc4d4cea6, 32'h4322fd84, 32'hc3b54378},
  {32'h44d9f921, 32'h4270e09f, 32'h4368caa5},
  {32'hc29f62a0, 32'h42f60c77, 32'h43d07f58},
  {32'h44e14dc2, 32'hc2888280, 32'hc38c85d7},
  {32'hc499bf10, 32'hc2d8133a, 32'hc373666a},
  {32'h43dcc5ce, 32'h427d9830, 32'hc29f9eac},
  {32'hc4e1fcdb, 32'hc283d77a, 32'h434b71a7},
  {32'h44f19dc1, 32'hc1458aae, 32'h4371b24f},
  {32'hc4f913ea, 32'hc3e01ce0, 32'hc2934b89},
  {32'h447133f8, 32'hc2a51fc8, 32'h4313986b},
  {32'hc4f2b6cc, 32'hc2263aff, 32'hc26a1e4b},
  {32'h434c8e9c, 32'hc2fa940d, 32'h428414e5},
  {32'hc4d0147d, 32'h433030a8, 32'h4349b43c},
  {32'h42faebe0, 32'hc3059e2d, 32'hc3b33655},
  {32'hc4bfd523, 32'h42c3148c, 32'hc1d3a0b8},
  {32'h44229302, 32'h418e10ef, 32'h4223e6ff},
  {32'hc49f7a4c, 32'h4308f55a, 32'h42f01260},
  {32'h44ffacc4, 32'hc324ff5c, 32'h4230b9e4},
  {32'hc4a17443, 32'h4391b834, 32'h434eced0},
  {32'h44cafdca, 32'hc2128099, 32'hc09eef46},
  {32'hc4a86c5c, 32'h4363a3d8, 32'h43af62be},
  {32'h4432a3e4, 32'h4295fe98, 32'hc361cc29},
  {32'hc3d7cda2, 32'h4354e4c4, 32'h41df052c},
  {32'h4423f56a, 32'h430253a8, 32'hc3777d4b},
  {32'hc4b46ccd, 32'hc18aa6da, 32'h433b0f4e},
  {32'h450a3616, 32'h43a2a877, 32'h40ce5c38},
  {32'hc3cd7b99, 32'h43aa842d, 32'hc35ad01e},
  {32'h4484562a, 32'hc31017a5, 32'hc24ca574},
  {32'hc4efa877, 32'h4386748e, 32'h4396afd6},
  {32'h443e3ef4, 32'h42fcb2d5, 32'hc1448198},
  {32'hc49aefec, 32'h424270c2, 32'hc1fe48de},
  {32'h445337b7, 32'h4324ac6c, 32'hc3523095},
  {32'hc4d6e351, 32'hc302e251, 32'h434c6cdf},
  {32'h44bd2667, 32'hc2a1c358, 32'h42df7eea},
  {32'hc4693000, 32'hc2388d6d, 32'h4324d74c},
  {32'h44ca528c, 32'hc2586d1e, 32'hc0c9e1be},
  {32'h4494ae50, 32'hc22dbaf7, 32'h43d6220b},
  {32'hc444241b, 32'h4388185a, 32'h43b4a801},
  {32'h43b17382, 32'h43f45960, 32'h431eb291},
  {32'hc4bba571, 32'h43b63fab, 32'hc291b86e},
  {32'h4433cb36, 32'hc3f881aa, 32'h42e8d3c5},
  {32'hc4fd019e, 32'hc3bfe257, 32'hc34daf79},
  {32'h44f099b4, 32'h433ae13c, 32'hc356fb06},
  {32'hc468ccde, 32'h431bb637, 32'hc3354db9},
  {32'h450850c3, 32'h440c708d, 32'hc2e77957},
  {32'h44f4408c, 32'h4241a7db, 32'hc1a2b422},
  {32'hc41a3cd0, 32'h43637ec0, 32'h42a60a94},
  {32'h45150746, 32'h4303101c, 32'h43184f8d},
  {32'hc22ef1ad, 32'hc29665df, 32'h4383ab51},
  {32'h45228a6e, 32'hc45d5158, 32'hc37fe419},
  {32'hc4664274, 32'h42a13c00, 32'h438f0e87},
  {32'hc3c1f00a, 32'hc312cedb, 32'hc254084d},
  {32'hc5095bde, 32'h43585652, 32'h42353ac4},
  {32'h45088209, 32'hc2c757e3, 32'hc31ac2a5},
  {32'hc508ef42, 32'hc29dc754, 32'hc352dc98},
  {32'h451f9810, 32'h43338185, 32'h431a9ec5},
  {32'hc3a14e48, 32'hc264d3e8, 32'h43cf8277},
  {32'h43748000, 32'hc314bad3, 32'hc370a154},
  {32'hc47e9b13, 32'h439bd542, 32'hc3281ff5},
  {32'h44a49f51, 32'h4381a20e, 32'hc296c6ae},
  {32'hc464d5fc, 32'hc317d7e8, 32'h42c9488b},
  {32'h43b128bc, 32'hc27252a6, 32'hc3a6b25b},
  {32'hc4313d90, 32'hc33a2e03, 32'h43e6f291},
  {32'h45018d85, 32'h4358c977, 32'hc2bbd981},
  {32'hc432ac9c, 32'h42a50975, 32'hc3bdf612},
  {32'h44c69156, 32'hc3361da6, 32'hc30b6222},
  {32'hc505fa11, 32'hc2a628a8, 32'h429b7a16},
  {32'h44ee9c71, 32'h433ae584, 32'hc28eb984},
  {32'hc3aea9b2, 32'hc1d41331, 32'h41290493},
  {32'h44d859c1, 32'h42e2a116, 32'hc2206530},
  {32'hc442d3fc, 32'h43abe84a, 32'h4318e089},
  {32'h4526d12b, 32'hc413d2d0, 32'h40f21344},
  {32'hc4fb7a6a, 32'h4244711f, 32'hc26834e0},
  {32'h44bf4477, 32'hc21caade, 32'h4392a580},
  {32'hc32b9a6d, 32'h432c337a, 32'h42e247f8},
  {32'h429c4950, 32'h430dbd17, 32'hc2e7006e},
  {32'hc3fe958c, 32'hc39ee870, 32'hc2098de2},
  {32'h4504a9dd, 32'hc3779d25, 32'hc192f86e},
  {32'h43476368, 32'h43d6ac1b, 32'h426b7529},
  {32'h44a14a3b, 32'h42e99623, 32'h4216a24b},
  {32'hc4887cd0, 32'hc2eb8894, 32'h44111a92},
  {32'h4217f360, 32'h42b4d331, 32'hc2c5a42c},
  {32'hc5172c2d, 32'hc12c17b7, 32'hc2a8ec5c},
  {32'h45297e40, 32'h439f0cde, 32'h437ed99c},
  {32'hc5064c58, 32'hc39fd962, 32'h43862ae4},
  {32'h431b53f0, 32'hc209af59, 32'hc3c04bbc},
  {32'hc5171f79, 32'hc3db7287, 32'h4347efe1},
  {32'h44e2d6fe, 32'hc30c61d2, 32'hc26c8fbb},
  {32'hc48f32c9, 32'hc38d17d6, 32'h41ddc721},
  {32'h439a2d34, 32'hc0cb2fde, 32'h411a4172},
  {32'hc43fe047, 32'h433598d3, 32'hc2998f5e},
  {32'h449afa72, 32'hc301e126, 32'h4393e9d5},
  {32'hc4f6b1f7, 32'h430bd55e, 32'hc341cd86},
  {32'hc43f62ce, 32'hc394609b, 32'h42c5bd40},
  {32'h433495ac, 32'hc152286c, 32'h4395d55a},
  {32'hc3415b58, 32'h43ddf7b7, 32'h418cc6ba},
  {32'h445e2ece, 32'h432ad282, 32'h43632654},
  {32'hc4e3b69a, 32'h422e3bcf, 32'hc321bf01},
  {32'h4462cbbe, 32'h42b63b53, 32'h43864a67},
  {32'hc467bdb6, 32'h4319efe8, 32'h426b1da9},
  {32'h44bd0fe0, 32'h4295e394, 32'h4106fa64},
  {32'h43c6b518, 32'hc24aed31, 32'hc29dfded},
  {32'h43d8c718, 32'h438ba13a, 32'hc2dd82a2},
  {32'h44f50c74, 32'h42e86e14, 32'h43282cce},
  {32'h437fdeb8, 32'hc2c5bcb3, 32'hc2f58727},
  {32'h44f9d7d4, 32'hc3e82c32, 32'h421b339f},
  {32'h445d57e0, 32'h43c22e38, 32'h43b27695},
  {32'hc33c34f1, 32'hc32092a7, 32'hc29a57eb},
  {32'h43f2e90c, 32'h430c12ca, 32'h434c20ca},
  {32'hc4cd8b9a, 32'h41f6e7dd, 32'hc29fa7f8},
  {32'h44a33381, 32'h43a63a70, 32'h42689270},
  {32'hc50097a9, 32'hc30ba5e1, 32'hc1dd2e77},
  {32'h445c47b8, 32'h438a54ad, 32'h4341b830},
  {32'hc402463c, 32'hc2f15e34, 32'hc1d76b80},
  {32'h43a9d372, 32'h4355e786, 32'h43afefed},
  {32'hc4725316, 32'h43168623, 32'hc403550e},
  {32'h4517976f, 32'h435e2f22, 32'h43106fbe},
  {32'hc379314c, 32'h43331c33, 32'h428b3e59},
  {32'h451379e2, 32'h4372bdcc, 32'h42459488},
  {32'hc4942e6e, 32'h42374a0f, 32'hc3852201},
  {32'h44d3fd4e, 32'hc2521256, 32'h42dda5f6},
  {32'hc4bd61ae, 32'h42b81c8b, 32'hc2d0a9e0},
  {32'h451a94f5, 32'hc314902e, 32'hc3307842},
  {32'hc507a10a, 32'hc35a2588, 32'hc3b1466b},
  {32'h44b9c945, 32'hc30d8f0e, 32'h431e897a},
  {32'hc372d880, 32'h412d53d0, 32'hc38a99fd},
  {32'h43381868, 32'hc372e54a, 32'hc30ecd6e},
  {32'hc4dc8ef7, 32'h406888d8, 32'hc2b4396f},
  {32'h41528200, 32'h418e6347, 32'hc2aa4452},
  {32'hc36b1421, 32'hc312d72b, 32'h43864cf5},
  {32'h452d9bfd, 32'h43380692, 32'hc1927177},
  {32'hc42b2240, 32'hc2cbfc76, 32'h430a3bd3},
  {32'h4473aa44, 32'hc2e71a0b, 32'hc2d56e9a},
  {32'hc46b576a, 32'h42d0b545, 32'h43dff9dd},
  {32'h44fc630c, 32'hc2b75b6b, 32'hc28add4f},
  {32'hc4fc3560, 32'h43b7cc55, 32'h41dea3ef},
  {32'h443255fb, 32'hc35c5718, 32'h438cfca5},
  {32'hc4c6a169, 32'hc2e46460, 32'hc0d32094},
  {32'h44024a58, 32'hc3b68c72, 32'h423a58a4},
  {32'hc4f7ca5a, 32'h4383cbd4, 32'h434d1397},
  {32'h4506cc88, 32'hc2f7cf95, 32'hc38d27ba},
  {32'hc4ec1104, 32'hc2b1d365, 32'hc2dab61f},
  {32'h43a29c2c, 32'hc3d71591, 32'hc2b0fb67},
  {32'hc50868fd, 32'h42ad7187, 32'h42b6883a},
  {32'h44859eb3, 32'h4331287e, 32'hc303059c},
  {32'hc4a90ebd, 32'h429f331d, 32'h4324eb76},
  {32'h44e96da5, 32'h4252f922, 32'h430716f2},
  {32'hc4e76f44, 32'h43251e86, 32'h4356c963},
  {32'h4411c68c, 32'h43387388, 32'hc2bb6219},
  {32'hc4209d4f, 32'h42aa75b0, 32'h43fbc777},
  {32'h4390172c, 32'h439f58ef, 32'hc3195c61},
  {32'hc45c5fc8, 32'hc2e90153, 32'h4327132e},
  {32'h45234eb7, 32'hc3badf2a, 32'hc259ba76},
  {32'hc3c5d9bf, 32'h425a972b, 32'h42b9f435},
  {32'h4513750e, 32'h430fc814, 32'hc33e745f},
  {32'hc4f18cd6, 32'h43a5e39d, 32'h4277ee4a},
  {32'h44e85913, 32'h43256ad2, 32'hc38b29ea},
  {32'hc4d41880, 32'hc2ede300, 32'h42c15649},
  {32'h4418341c, 32'hc35543a2, 32'hc38ae455},
  {32'hc4ddda80, 32'h43dc7f5d, 32'h430192a4},
  {32'h44f49674, 32'hc2b9d678, 32'h430c2707},
  {32'hc4905a9e, 32'hc32e2050, 32'hc2cb4a4d},
  {32'h44007e22, 32'hc411a665, 32'h41f88b14},
  {32'hc4a655fc, 32'hc18d6cca, 32'h42dfc5b8},
  {32'h44502adf, 32'h432fc502, 32'h41f59b25},
  {32'hc47e4f54, 32'h41c2f983, 32'h43b6142f},
  {32'h44ac6df2, 32'h429dcb97, 32'hc3a2077f},
  {32'hc4078349, 32'hc39357d4, 32'hc36ed64f},
  {32'h4489ea35, 32'hc2c7ca96, 32'hc2143c9e},
  {32'hc491c057, 32'h4388faa7, 32'hc3ead741},
  {32'h4450ed16, 32'h43140fa5, 32'hc301520c},
  {32'hc492ec85, 32'h430868be, 32'h43de9656},
  {32'h44b99ba0, 32'hc39f899d, 32'h43ee89e1},
  {32'hc35802d6, 32'h4395b517, 32'hc2808769},
  {32'h446887b1, 32'hc306aae3, 32'hc4010060},
  {32'hc3cbc21c, 32'hc35b18df, 32'h42b803e4},
  {32'h45056f78, 32'h43c06b66, 32'hc39e484c},
  {32'hc4e4827e, 32'hc2619dae, 32'h415278d7},
  {32'h4324fc20, 32'h420b6e93, 32'h41b83ea5},
  {32'hc3f3fdf6, 32'h4399c6fb, 32'hc2b84d0d},
  {32'h43aaa8be, 32'h424e8076, 32'h43766586},
  {32'hc4cdaa26, 32'h43c974fb, 32'hc188fb26},
  {32'hc227ca48, 32'h4380cb6e, 32'h43bc79ec},
  {32'hc4d07938, 32'hc25b36bd, 32'h430c16a7},
  {32'h448ef7e9, 32'h43a9bae0, 32'h4223fb7e},
  {32'hc4dd40f6, 32'hc31237e0, 32'hc31263c8},
  {32'h442c4f69, 32'hc1894eff, 32'hc37488a0},
  {32'hc500b5ee, 32'hc2b0e59f, 32'hc2ef14f5},
  {32'h44ec6bd7, 32'hc2dfb394, 32'h420eee10},
  {32'hc47cdc88, 32'h4279a4a5, 32'hc34df561},
  {32'h420fa858, 32'h43dafc48, 32'h428888f5},
  {32'hc4f4bac0, 32'hc31dcec0, 32'hc38f1d62},
  {32'h44088bee, 32'hc34e84e1, 32'h42d71833},
  {32'hc2dd1d80, 32'h43b954be, 32'hc28b50ef},
  {32'h44fa9502, 32'h42a194fb, 32'h431853b2},
  {32'hc4a0b3b9, 32'h436a73aa, 32'h43db4a0b},
  {32'h450b1910, 32'h43741c57, 32'h42f45bd2},
  {32'hc39c1ba6, 32'hc33339b3, 32'hc3858dee},
  {32'h44fe420a, 32'hc2a95238, 32'hc29d048a},
  {32'hc4da513f, 32'hc2b05952, 32'h43b7ad6f},
  {32'h44e26cbd, 32'hc3345a3d, 32'hc2a69ae3},
  {32'hc445f968, 32'h42fd0ec8, 32'hc364ef1e},
  {32'h44e64dfe, 32'hc1ac63b4, 32'hc30d6bf8},
  {32'hc406d9dd, 32'h43679b02, 32'h43914b92},
  {32'h4402d1c8, 32'h43a527bf, 32'hc3541cec},
  {32'hc34dad0a, 32'hc39e27d0, 32'hc30299f4},
  {32'h44643ba6, 32'h436ee20e, 32'hc2168ae4},
  {32'hc36847c2, 32'h42ed0b34, 32'hc2f0b704},
  {32'h449084e2, 32'hc34feac7, 32'hc203f582},
  {32'hc4b7e17f, 32'h42a36470, 32'h4337abce},
  {32'h4455bcd2, 32'hc334c9c9, 32'h43127eb8},
  {32'hc4c18069, 32'hc3e2ee28, 32'h42ba5a41},
  {32'h45083ede, 32'h433ef578, 32'hc3589704},
  {32'hc409a7e4, 32'h4394ebf3, 32'h436acf20},
  {32'hc4e6a7de, 32'h431951a5, 32'h4382b1c1},
  {32'h440cff45, 32'h4305cb2d, 32'h42707eb4},
  {32'hc2d86346, 32'hc3b4d3b0, 32'hc386ff28},
  {32'h445e5261, 32'h402ba0f8, 32'hc3a491f6},
  {32'hc4a71311, 32'h429d76be, 32'h42b6a5ef},
  {32'h43c2a280, 32'hc42829ac, 32'hc3ae0090},
  {32'hc41d7672, 32'hc3e05f3d, 32'hc3856256},
  {32'h44bf8a26, 32'hc266baaa, 32'hc3378310},
  {32'h3fc31000, 32'hc260846e, 32'hc38d9b61},
  {32'h43cdae80, 32'hc3693410, 32'hc34158e9},
  {32'hc4f025aa, 32'h41a76636, 32'hc10f3201},
  {32'h450befe6, 32'h439736de, 32'h43efaa0a},
  {32'hc4953e75, 32'h4231aa75, 32'hc1f418cf},
  {32'h43f9e53a, 32'h430b8e29, 32'hc1cac6fb},
  {32'hc48d3a87, 32'h42ba7840, 32'h424d994b},
  {32'h4465e22c, 32'hc3597b95, 32'hc2b5cb3b},
  {32'hc445030a, 32'h43cdc61c, 32'h4380cb27},
  {32'h4492c778, 32'h436eb197, 32'hc3b2c034},
  {32'hc401523f, 32'h415d5f16, 32'hc1493c54},
  {32'h44495d24, 32'hc2b8135b, 32'hc2ae29dc},
  {32'hc50c3f40, 32'h43854453, 32'hc3bfc968},
  {32'hc510cfd0, 32'hc4082cd6, 32'h435d1e74},
  {32'h44a0ef21, 32'hc2a77f85, 32'hc2ddf286},
  {32'hc4491949, 32'hc2c8b808, 32'h43811f4a},
  {32'h44354030, 32'h42d3bf50, 32'h426f9819},
  {32'hc4da5f79, 32'h430c5896, 32'hc33e8155},
  {32'h44a84b34, 32'h429e0107, 32'hc3304ba7},
  {32'hc44f5524, 32'h4301a7c8, 32'h43c76483},
  {32'h44e7875d, 32'hc3322d0f, 32'h435241f4},
  {32'hc4040376, 32'h4303df83, 32'h419ef925},
  {32'h44f464f9, 32'hc2ef2b55, 32'hc342891b},
  {32'hc4d1e0f7, 32'h3f932595, 32'hc34d2474},
  {32'h44c49dd4, 32'hc2b63cf2, 32'hc2830590},
  {32'hc4cdcf15, 32'hc2d0f1b5, 32'h435a05bb},
  {32'h44dd098a, 32'hc4007b23, 32'h434fe482},
  {32'hc389ec08, 32'h4269e79f, 32'hc390ea9d},
  {32'h442048ac, 32'h43a4d9f7, 32'h42eb4bf9},
  {32'h4288970e, 32'hc30ada9c, 32'hc338f9bb},
  {32'h450088c9, 32'hc2cb9dff, 32'h42964100},
  {32'hc3874e3d, 32'hc3b59e80, 32'h43908002},
  {32'h4388cac0, 32'hc02cd77c, 32'h42bcf376},
  {32'hc4186a42, 32'hc3c3d3a4, 32'hc309ed4a},
  {32'h4481083b, 32'h4312d4f4, 32'hc31b48bb},
  {32'hc4d855da, 32'h42d49c75, 32'h43404147},
  {32'h44a38b56, 32'h42014fb3, 32'h42ecb932},
  {32'hc4f8bd81, 32'hc2cb9285, 32'h43279acf},
  {32'h44863ec4, 32'h43bff2a1, 32'h439fbc12},
  {32'hc4755d6d, 32'h41c4eb68, 32'hc2e2e751},
  {32'h4371ea88, 32'hc2acc3c7, 32'h42e376c7},
  {32'hc4b4d0cf, 32'h424727d0, 32'h42758ab9},
  {32'h45147968, 32'hc3af0b14, 32'h428a39a3},
  {32'hc44e340a, 32'h43611a64, 32'hc2e04383},
  {32'h43826849, 32'hc38b2414, 32'h43f7265f},
  {32'hc43c2e01, 32'h4306aa3d, 32'hc32681ba},
  {32'h4511a737, 32'h438abe79, 32'h438b13c3},
  {32'hc502fb02, 32'h42ba1960, 32'hc355c35c},
  {32'h44da96c7, 32'h4326a1d8, 32'h419fefac},
  {32'hc507ef4e, 32'hc38d1e08, 32'h43507c7e},
  {32'h4510d7da, 32'hc2a21526, 32'h438ea9ec},
  {32'hc444d1b1, 32'h42db3399, 32'hc3147b1f},
  {32'h44eb5ab1, 32'h42b7a22f, 32'hc3a7b64a},
  {32'hc3d96d4f, 32'h43404013, 32'h43154ffc},
  {32'h44818d32, 32'hc3024130, 32'hc2e47ad9},
  {32'hc50fe0ff, 32'h43177aee, 32'hc274d3bc},
  {32'h45027bd8, 32'hc307c693, 32'hc29d8d33},
  {32'hc51966ef, 32'hc2888ab5, 32'h43efc196},
  {32'h44f142d8, 32'h4356a29e, 32'h425c5e1e},
  {32'hc460494c, 32'h42b98d77, 32'h42c7bd49},
  {32'h44d30846, 32'h4234631d, 32'h43053bd1},
  {32'hc443cbb3, 32'h426afbe5, 32'h43461d5c},
  {32'h43cd46b8, 32'hc29d825e, 32'hc156e2a2},
  {32'h41e3941e, 32'hc3dc5810, 32'h43141381},
  {32'h4366d4c0, 32'hc2443b16, 32'h43236cce},
  {32'hc4cba02e, 32'hc3af69ea, 32'hc2691c04},
  {32'h448a7758, 32'h420ac28b, 32'h42e4b32f},
  {32'hc5081d8c, 32'hc2f747e3, 32'hc37aefff},
  {32'h44f3912c, 32'hc2193a04, 32'h41cfd97b},
  {32'hc48ea5ba, 32'hc3627c8a, 32'h4365f808},
  {32'h44204ed4, 32'h4281cb8f, 32'h419bb91e},
  {32'hc4ed633d, 32'hc29f950f, 32'hc3672d38},
  {32'h4482cdc8, 32'hc40172f7, 32'h3f02ef12},
  {32'hc404ef23, 32'hc1c3484e, 32'hc156dcfa},
  {32'hc428037b, 32'h43ee42c3, 32'hc2f787c5},
  {32'h451bffdf, 32'h432ff78f, 32'h430a1b1e},
  {32'hc4972304, 32'hc2ad66f4, 32'hc28d4771},
  {32'h44e6200c, 32'hc3333bd5, 32'h43018759},
  {32'hc401b850, 32'h431748a7, 32'h426e90e3},
  {32'h44130cce, 32'h431644fe, 32'hc1cc4887},
  {32'hc4d9c438, 32'h3e683560, 32'h43a06de6},
  {32'h44a38670, 32'hc416b4c6, 32'hc2c07f56},
  {32'hc4990fb8, 32'hc3056120, 32'h42dfc3a5},
  {32'h4510be87, 32'hc3180dea, 32'h438419f3},
  {32'hc4f4ad39, 32'hc363ee3c, 32'hc2f5b69d},
  {32'h44e58d20, 32'hc30e417f, 32'hc34f040a},
  {32'hc4bdc29e, 32'h43fad2fa, 32'h42f9ba40},
  {32'hc394d9b0, 32'hc1db3bde, 32'h429d9fc3},
  {32'hc44683e6, 32'h426452e3, 32'h431701a9},
  {32'h4194a7c8, 32'hc346a5ff, 32'hc3e7b6d0},
  {32'hc40c9c1a, 32'h42a85d58, 32'h4241ac67},
  {32'h4410d7d4, 32'h4373593a, 32'h42369fee},
  {32'hc4400530, 32'h437627ce, 32'hc2a053a3},
  {32'hc276b0d0, 32'h422facc8, 32'hc381553c},
  {32'hc494012e, 32'hc2f81ec1, 32'hc34e56b9},
  {32'h44e3ace9, 32'h43747f8e, 32'hc2166576},
  {32'hc424c67e, 32'hc315a090, 32'hc2397f46},
  {32'h44db7f5d, 32'hc3832822, 32'hc3d13ff9},
  {32'hc4d2face, 32'h422c55bb, 32'h431b5d36},
  {32'h44a6910f, 32'hc35544dc, 32'h431fe022},
  {32'hc4595e14, 32'hc2821ad9, 32'h42bd4608},
  {32'h43b11344, 32'h43158f5e, 32'h41d48276},
  {32'hc49dd340, 32'hc1f9b849, 32'h41a4e612},
  {32'h447dfdaa, 32'hc358c946, 32'h436b0194},
  {32'hc4d7602a, 32'hc29ab3c4, 32'h4351423b},
  {32'h44fa6d4b, 32'h434fab86, 32'h441a3405},
  {32'hc4fd7374, 32'h43114bfa, 32'h4175c78b},
  {32'h44806546, 32'hc30d45e5, 32'hc32a4e0c},
  {32'hc50f992c, 32'h438cf4ab, 32'h42fc421c},
  {32'h43e3db40, 32'h4233554f, 32'h4391029a},
  {32'hc49b9ec5, 32'h432eb8ff, 32'hc2a67b80},
  {32'h44b0b006, 32'h42849df5, 32'hc3569620},
  {32'hc3949750, 32'hc2c4e9de, 32'h42794cd9},
  {32'h45053a11, 32'hc329998d, 32'h437d6437},
  {32'hc214f5e0, 32'hc3a835f1, 32'h4289086e},
  {32'h43cfc486, 32'h43a2aee4, 32'h4280f197},
  {32'hc4f5f177, 32'h4355451c, 32'hc33edd32},
  {32'h44999318, 32'hc3a605dc, 32'hc246c0ef},
  {32'hc51f87ce, 32'h4352748a, 32'h4403a744},
  {32'h4247b6e0, 32'h43702f28, 32'hc37eee30},
  {32'hc3dadbb8, 32'hc43487e8, 32'hc377523a},
  {32'h44f069ca, 32'h4287fa78, 32'hc2959608},
  {32'hc50f33e3, 32'hc3ad12d4, 32'h3f95ab94},
  {32'hc3942474, 32'h43548d83, 32'hc407e0b2},
  {32'h4511a385, 32'h42a5c345, 32'h43947961},
  {32'hc500b7cc, 32'h4366f3b2, 32'hc35413e1},
  {32'h44f5ca16, 32'hc185d471, 32'hc1972f57},
  {32'hc4607278, 32'hc39c5f3a, 32'hc25da038},
  {32'h435f48b0, 32'h43be6aff, 32'h42da581b},
  {32'hc48efadf, 32'h430cdbe9, 32'h4143e95c},
  {32'h45251ce4, 32'hc35fc202, 32'h42b56375},
  {32'hc498897a, 32'h4388fd49, 32'hc3808004},
  {32'h44fbe180, 32'hc36353b5, 32'h402a2844},
  {32'hc389dd58, 32'h42bab0d4, 32'h4313f548},
  {32'hc3209888, 32'h439fdccf, 32'hc2c2c69e},
  {32'hc3c26e80, 32'hc2d47c09, 32'h423f24bf},
  {32'h44fc3cbd, 32'h42c29d48, 32'h431d1164},
  {32'hc4fc9755, 32'hc3e026e4, 32'hc3e261c8},
  {32'h44ffe649, 32'h4298a7a5, 32'h41b1250f},
  {32'hc446b8f2, 32'h4309c04a, 32'h43583bd9},
  {32'h449a96d1, 32'hc33b4d8c, 32'h437ee961},
  {32'hc4d0192c, 32'h4216ba34, 32'h42223948},
  {32'h4430aae8, 32'h43298cf5, 32'h43e660c3},
  {32'hc3820e84, 32'hc328f3c8, 32'h43b94ac5},
  {32'h44b91704, 32'h42b14a43, 32'h42eb82e2},
  {32'hc46fb95c, 32'h42d2f0c6, 32'h43bbd24c},
  {32'hc1028540, 32'hc0fa7667, 32'hc2938323},
  {32'hc506ccf6, 32'hc31a76bb, 32'h4381d70d},
  {32'h44393b8a, 32'hc302b3dd, 32'h43da20e1},
  {32'hc3377e20, 32'hc39299b9, 32'h4369cf5b},
  {32'h44c03530, 32'hc333a2ee, 32'hc1252386},
  {32'hc3563e90, 32'hc2d75ddb, 32'hc3609bfe},
  {32'h44d27edc, 32'hc3bc5b69, 32'h43d935d9},
  {32'hc3d95fa8, 32'h440938a2, 32'hc271b5bf},
  {32'h446a3c30, 32'h4225f742, 32'hc34b283f},
  {32'hc492163c, 32'h42802050, 32'hc374300a},
  {32'h445fe7bd, 32'hc2a077ba, 32'h43384e34},
  {32'hc48bef80, 32'hc1a593ea, 32'hc383560c},
  {32'h450b7c13, 32'hc2b7f4d6, 32'hc3bb9a75},
  {32'hc4d119f2, 32'hc3c4b6a5, 32'hc37d3e3e},
  {32'h451709da, 32'h440b9267, 32'h434dbbdb},
  {32'hc3558558, 32'h4405d036, 32'h42fd3004},
  {32'h441a53eb, 32'hc340b182, 32'hc230e97e},
  {32'hc4e75784, 32'h433dc92c, 32'hc225dea8},
  {32'h44a1559c, 32'h43653225, 32'hc31030e2},
  {32'hc5163f8b, 32'hc28a62ea, 32'h41dbdd58},
  {32'h447ef47e, 32'hc3bcfae6, 32'hc384dae1},
  {32'hc2d06f30, 32'h42eddd49, 32'h4377136d},
  {32'h44cfa471, 32'hc33950a3, 32'hc18934fa},
  {32'hc3cb73e8, 32'h434cdb9b, 32'h42b3a6e6},
  {32'h44907246, 32'hc1800398, 32'hc4028fd3},
  {32'hc4b070a5, 32'hc2af180e, 32'h42920fff},
  {32'h44b09456, 32'h42276cb2, 32'h42c5a4a6},
  {32'hc441e264, 32'hc3e438d2, 32'hc2d6c21f},
  {32'h4489297d, 32'hc26db7fa, 32'h424d7a20},
  {32'hc4180456, 32'hc37da078, 32'hc2c25537},
  {32'h44d0935f, 32'hc38bfb49, 32'h422985a4},
  {32'hc383d046, 32'h431ac607, 32'h437eab64},
  {32'hc4241376, 32'hc2586bde, 32'h4360e79f},
  {32'h450ca259, 32'hc352b009, 32'h43ac0477},
  {32'hc41c6150, 32'hc3979caa, 32'hc371eab7},
  {32'h44f0edda, 32'hc2e8ad27, 32'h42943c62},
  {32'hc453366e, 32'hc30c5e85, 32'hc217bb55},
  {32'h44813c88, 32'hc35aef72, 32'h42e06582},
  {32'hc31d20c4, 32'hc14f5eb2, 32'h43246faa},
  {32'h43847118, 32'hc2f25f72, 32'h43cc471c},
  {32'hc34ca0d8, 32'h4192642a, 32'h43743c94},
  {32'h44be345f, 32'h43056897, 32'hc1941da7},
  {32'hc483ec84, 32'hc218d687, 32'h4310c142},
  {32'h43e173e7, 32'h430667c4, 32'hc32dff7f},
  {32'hc4e79ed6, 32'h436731cb, 32'h4304f9f8},
  {32'h44d5f6db, 32'h4392def6, 32'h438ba2ee},
  {32'hc386f019, 32'h438baa2d, 32'hc3435426},
  {32'h44d5439d, 32'hc39fa883, 32'hc28224ac},
  {32'hc4d70957, 32'hc369a6a6, 32'hc396f141},
  {32'h44fd53da, 32'hc356de4f, 32'hc3563a03},
  {32'hc45238b2, 32'h43b443fa, 32'h419ad14e},
  {32'h4422ece5, 32'hc2dd3f6e, 32'h430a1c34},
  {32'hc4e5c848, 32'h42e4c4db, 32'hc38ec584},
  {32'h451553b7, 32'hc27bb284, 32'h43776401},
  {32'hc4bc9bbe, 32'h43cc1963, 32'hc3a9bcda},
  {32'h44a60bd0, 32'hc2a521d8, 32'hc3b6f55d},
  {32'hc3d25140, 32'h4395ade2, 32'h439f69e0},
  {32'h447b9bb8, 32'hc2e22ebf, 32'h43a5dadb},
  {32'hc4ae5db1, 32'hc310b1a0, 32'h43ed7bf3},
  {32'h4470dc5f, 32'h43b3962d, 32'hc3c6cc12},
  {32'hc3edcf88, 32'hc244aba9, 32'hc2be61fc},
  {32'h44b63db4, 32'hc28e496e, 32'hc2d6e58e},
  {32'hc4512450, 32'h432ff453, 32'hc301959a},
  {32'h450400b2, 32'h4291b17d, 32'h432a3887},
  {32'hc499c697, 32'h4303e796, 32'hbffd8e04},
  {32'h44b04af4, 32'hc1936777, 32'hc2a90b9a},
  {32'hc505f08c, 32'h43c7b259, 32'h430dd26f},
  {32'h44916f43, 32'h43bd2506, 32'h43051c99},
  {32'hc50181a7, 32'hc32d2c3e, 32'hc364c0f9},
  {32'h40b14c00, 32'hc386ff6a, 32'hc4076026},
  {32'hc4af34f8, 32'h43039442, 32'hc3c44769},
  {32'h44f0d141, 32'h4388bd01, 32'h43abd784},
  {32'hc503f89f, 32'h42d3de22, 32'hc33b4184},
  {32'hc2700f20, 32'hc3c21538, 32'h410bfb2a},
  {32'h44401a68, 32'hc1b747ee, 32'h432618c1},
  {32'hc4a1662a, 32'hc261e856, 32'hc2d4203e},
  {32'hc4a0d423, 32'hc2a6eaa6, 32'hc31bb571},
  {32'h44466d04, 32'h42b006df, 32'h429c8c7d},
  {32'hc50fcf76, 32'h43ae8c7b, 32'h429f5e67},
  {32'h437db9f0, 32'h41a97158, 32'h42f0d6b8},
  {32'hc5059fe8, 32'h414840b4, 32'h43b2203c},
  {32'h44d2d583, 32'h42bb0e67, 32'h43cdba92},
  {32'hc4c3a95f, 32'hc254f1fa, 32'hc2091236},
  {32'h44e263c7, 32'h40bbb175, 32'h42904e00},
  {32'hc5049f94, 32'h4336479a, 32'h42b82be8},
  {32'h44059252, 32'hc296c014, 32'hbf6855e0},
  {32'hc506888f, 32'h4209bc04, 32'h42adf395},
  {32'h44b8508c, 32'hc28980b1, 32'h43070b04},
  {32'hc4e82229, 32'hc175127d, 32'h42d3909f},
  {32'h4414842c, 32'hc2b7befe, 32'h430d7c88},
  {32'hc4d872bc, 32'h431a735c, 32'hc3183ca1},
  {32'h44d2bf60, 32'h42681a56, 32'h42e2f7d3},
  {32'hc4dc77ad, 32'h42722c70, 32'hc2fc8388},
  {32'h44d3cf52, 32'hc2bde0ba, 32'hc3c351d9},
  {32'hc4ab5354, 32'hc3939d06, 32'hc348e65a},
  {32'h448840b8, 32'h3fd27f1c, 32'h43b5e76c},
  {32'hc4d779f5, 32'h4392d79a, 32'h42ecf5eb},
  {32'h447ce1f2, 32'h436b2037, 32'h429f5b4c},
  {32'hc4b36064, 32'hc1d2b73e, 32'hc2993c8e}};
