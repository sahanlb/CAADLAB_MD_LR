-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kvulKTwxdM1Y8neRL/980l936+6K30FFtuSyt1aYTGftdTKTkiendsH1c416jcrBfupbejmmekAh
89gTvEqPSNPjdpaTusXNIMhifgfo+eDmACgQKe7oA9rceBQ+aZw8hrp5RSqoHIlhmKjzMdGhoPNw
JisWR08cR8tl2E3wHAo6cTAeUFH/4L77zFOPi1yfITniw3xSezNIDl0bZGUKS6LjQ5CoCRlaYtSY
czeSdeLNM5XxBLubknF1hwGqHwYEQwia8iRfUlGWlOiv2RrCHNjHC4wxwSloDl0UH1idWWtEu0O2
Bwu8sOEPSWsMz5+SIrpgPJWKSjJm6lY9WABvgg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 81696)
`protect data_block
kmTR6nZ8rh5diL598uTKXYj3snYO9onYfRqkhTf6IdHSC30FgE/easjjsFvWD1L844MWZ7ZX+YAT
BEnPkrEx3hVuja3rVoCXLexRRE3t1Pq1lx6oj10lKI4ymmfoTPdBDk+V+CSBtJH3rDnbG4u2En+F
bqVzXz1e8j4dqaapHGFk56ubgHxVPVL8p5TJjKpl4nLiFwKPbG8OCOeBkAmt4o8P5iG9AQTrPBMF
PJGGROemNUw2V6usCr83207faU9lBRkhN1zGNPPU8GYsSG/1AKWwNR4JkOqNGAoDhGQ/IwvgyHB0
R4SrrVseQaqw6gIPKZ4V9UIVlA8QI8D2JP+872tUKQUngiL2pGIe1OG5gmKIuHosooC+L9gO8uZW
wZRjZO5ZeEGZ6X/bCsuBjmRaiqVb9H91XKgNRE98UlDX5aaKTydPVaQlUGghdxWcHtsKFdb85LFK
bfIgwiB0pr8Et8pRFa10Z8L90KUbovEJf2pI5B+0pi+4hZaT1TYIky2hjshK71XcfGDjJjgJ3+9A
5LhqjK7IoeyWNNo2ZDJHhfTDFs42bosi9A8MiaOh6xjQkPLxGtfpg0BGO7PF07EkHDbpdQUB+eGc
057CeDxbnHw6I7+PzXiWLX7aarJ6y01tuJI9+M3h8imtKbi7ybPArtySmvAvBcYPyJeCMQ1yOJN9
ypBJRKUfRvxcBSdpABaVOZMVtl9KmvOvN2/L38cXlEHPqaobWRU3tviWplkgd6oSz3YSF003Rm61
10uRVPCFTEC1wzSIH+fYA7XFpXn2VKsASUyGDpnZWCRUSY7SHQjjP8lMRdmE0Zlbtf8XySvmRzlt
fQ2/BRjocLPyESyZVk+oWXWUIOj83xbUWE+9M6o8JmmTekfZojY2pBqQGAXd95Dp+H4ZFV09Gh25
Nb8Vub5JGgnuHr9gWbmzSRrVdv8H9XGXFriP7NQnarHDDcuPRV1N/6Ii8n4bWR9fTNfn27gTBDeN
AGIFmcA8SzRRXN312lFNA8h5WvXMnP4y018HJkTMzspGCKJvlkcbJWkHA5LB0s4kO6r0NlLmqG2I
iJkqU4Sb2sazPsDdiS193YDcmW5iTwt3p3U5UMtHfHdM9/LnuFtL95ArbK5I92eNJnU7pn5kcMcE
jZzFzRzwbZhoNVb1TiTq7P3o5xM1SufM77Ynx5G90mTbzsPYuGYq56hDv7nVjxDk/Et7Bp7GbxAI
ep2/f4tkNQIvGHZAU6mC5qfqdXF7got625ZqvIGVYyva7hJb7xNo5JMj+R6scYPMqm6+qLWn7OjD
hvhpxinTlPdpZSl5CPDYOJu6XHRK43W85IqGFFUInKh9x1LnUJRcD5Mo9kwmZf5pUcIz4cyFT59N
QqW2+/fiUzCAjS8ryR6+FHyDiUHSHGO1VmuyAbMkl8zVRyWIvMJNHIMqthN6aLZb7xu3/oMCzgqZ
vbHzag29crd6zte1meZSXaWkpCfodnL0jcXRCRsGhb5+oDfJwD7YpfJHcPtJ1cXM/qCJgPAkoTFU
wQx5UDPt8LlfOKsXVT+37hOEpvcC2zq4AjMXR311rPKfQhmHERIU7fKv8lbmYyrHAbnsZxv+cSSQ
xrEpIBLIWxXAN8rHjhF2Gy0QdPnxi4bKYzzLVozOQKX5/QMOMH7Oncn3EIx529t44vzyWVWkbg1P
FfyqpcAxqXzcgmHRspGvcztoODLo/cqD71WIIL4x9Z8BqUR2syasmCTgvBTqgY/9M0UMs23oBOGN
2oxgxpdT/laP9aPiBLn8rdsjZsfSkTybIGQzZc4EvyKDuBerQ7jhq3yiuNlf1C4zc0ZQCEM6p9yc
QwqW3IDjddJXdMOFk33NJVyc697LqB4JVdJJJ36hkgEzTrk0zhdElq+oMPeih4Q5zz+AxDdRtsbD
Ttgm+DLutVVs0vP7Ronfx+BC500Qk5uNXu3nX090O0uoKzdD8cUAyQ2QHn+nUc9o3r2Wbs3ZgpxT
Q4EkKvyQmPILP99c1FVgDKosAum1V6/K8aGB7iQZHGcM6Ez8CC9W2xuqtEPsQpe+TTJygIiCUUOC
go/q8Pg2QU69k78dTj205Xni+EL7EFqNm4p6qoEeZT6IDugICa/wChzHoHRI5Kcavi/3Gt7DOL9F
AflckwMD+iWCq2Zv2OWKts7w0lKF5YkyLWNdIXyzJfJ3gbDr2INN/gVef0xuUsG4lHxTTiwcgrk+
JFc5d3tm5hMVzBkJIDQBCvRrw22e5UWQ/pLrSAurZUdSKy5b/HE5sX7ToaHHarstZblT1kTZP1wD
i2oLZFalt+VuNveSi2UdkSq5ej6KsoaZ1zmj2Li52z4dSZuk5CBQ4nFSv1lbYfeTv7b8fRJDqjEs
KlQrkKcFfpW/2oQqHw8K8x6QQdj28rblcQz7EzfMLM5oNy3c8S/q70qpmetzI1fiAH3F3DKJqSwf
fVMHJGgFzj/xkKFIPDkBG1xGPD75jkYR/0BSn/1YY4bflrQvU96qv2wz6cOObhF0pKSsQAxzJLRc
OxsSFjItBxJHumAuQypSFNBwunna1Vy7yZa7IJLRUVaRYbqqISkWyUPfZ4Lo5jp1vYJWk4ZLjsWG
jgVeOaHlRTDEVX7vr5nB43rjJACpKtgirrIHBMDLviLlLFACLsDn3/o2vVKO0pvRKHC3T43fVANs
g/LR+gjmvab4pQxYunUrCQHRAsKsdE68OvJOW8Od7SosddBfWSr1GXQ4TtizusfgSIQSXn0V/twr
dBhyDdyZWEN9TCb8fh7HGPamXMjsLlNpXhWFEsNQQymrrPEP0F+xEzt45/jDZTbSWYoUxLsJCLSP
pNom4GSa/fd8RlNwXGQDY6zOXs3LM4I3hemklQw3T2ajCB8LqIuD0L3y2tJAZdG2lsb93ehbzIRZ
DCWyRrWR/gj10ChRewaRvOZ12zJl6Phi5J26zYG0Bk+QWOFPzZZBANAhLYd3LHB8hgEu0XW+6Gal
ItRNfMDaV7V1nSQ1hurH07RXZq7zmuLvtpeqPcVuAWDldehKpfy3RTxSHgNV0EAijKOcACscDGK2
PQ3GbF3gxmk6/xISvwcdSOK33VI7stVRiZkBjpuBcpPyXYgOrLsH9hKyfjadcFwOdlSR2Wpt17uM
y8LBpwiQDsDZXoeCfh13xhM4jIQyiG7XQbAKGPipCR1g5S5De2+eGCgZrMSTpB8vFzt/ecUEY1bC
LTlYzs1S0KOQG3pFByVJNHSFJPFWTr0fBizsvx9xlzDPeSSIXlbS6LlKmGWuE5kDpvx6/LgobEpc
I2UWJ9/zeJV8NEB5d3aq41Yq3qTxANLnKwZSm/dqmlL7iHfuthPZjRKtzFwa3lWDqc7/PNDF4nCo
7CdmnyzwvI8vYs7mHntwCL6G6nfvaNKfPG9fy+uB8AtL02/tvDOnjX+sJ025EaQZWaqi8rWWZzeY
y9ihT6BpPL8xRgf9frsWbJWD2RlwhfR0Oo81Czc6i043nJ/TXLiqnsA/6jh6G7h6NugL8XqPW/L9
679IyCvApBVcjCr+THVi2UW58fI3AwdekB+KynJS1gxbjqp4Xq7eyhUkJcwugdH29MSqr44/zDMM
mZuQH3yJ7PGdr1aWza/+zyZmph6K4NDeqZCLdRGXQjvHix6fXYhRYteO/dQzuPDrhc3H5u/ZK1TE
HaSnQSq2xmH6PL+YQ1oshVVLyBveHyVxv8hF9y1BARXzGd6h7+3QCVPr164/391mgwktMLE76dpZ
dDCtelysNk6L/Yh9ZBpj59Ymif5VGNsvAE+4aTbko+mfAK3tq5U6mlSxQnPbpfQez1HecV20UQ8T
9DFTdju79eIvhZ/do/XkHSW2ceXKD3+DrUR3aG7APz7/diyjpNj5Fhv36miKQyYUZHEyMgGTTLWO
doJBum2fWTojOY80ZXCKN8oRChCbTDZiMNH4TLgnkcRokBnKcbcznh+9LxyeItEojWkS/CTJ6YYe
2J2wm0rvjyYKkb9I6Borvpltp+RLCHS6tmhIXeHZk1d8ohE77hzY5Zzck76SFZ4iuiqaArqpK/2i
jyfOFf9MLUfDNlNj07wugeqkeiVcrj1l4owtEcg+/72RytNlJkqb3WrQaRn/K4fclkrqf8AM0Unb
NRIobw2YkncTnoVR7vgpcqKbRCp1KXp4k3YcGGG3uX448FmhXxBvlyh1FNJR0jedIuic8nblz7LH
4VHP13kitoOyZ5krnn0nXYIwvvCF1l+9z+j7bLx7vow2oICvbGnMvS1DlvthFv6gITwg7LBhe1fX
k3UG+rPMiaXt6zWxqzv6pOkgnZuvM75LxtPVD5vJVuxGzJArAQ10dndx2zSSq8bAVfMC8VNHvUr6
NoUV3wYC/LlADlH1fN8peIBnp2y5+PQ1a1HE2dO4l34Qx3XGCBmx+zwom6T4wN5CCW84AOsrr0DX
nIBcmS41bhL3u3alUKg45leKCayqblGserrqwoRovkN0IFsKnNdXRTqWiqZdg7R1lBmZ6Vm0dyRT
fAimHbsQu5Ojaljj34rmbqBpLsaCap637BDzsm5GzOs8sxwHHLryV4t6UPYGmuC0nMrnCwQH8k6T
BTZT/XdO2Ix90BQ89QiZ12TGcFxeUHKs9JGUAFrRySZfoIsTsDLX6IUA6kuWMLHNdJRXe7rvx5Ow
4Z/7eUtXErLgBF7zGPLaAv9JyxFAeVb3trvEhyzRuv+ITBKI3J3CZ4C77BLWLca7rXd0Otm2SSza
F6UUyVLnqzaAQ25cN2gx7vIj2O1Z2DyuLYAauzoznYVcB4HWC2sLCcSDnA4yqpJ0Ndq4iP7yA8vZ
rRdAY/Ku4oWhEBlCNJZDWwgqt2mfrgbdTvAduKmh18YWXDXU4LsebfeL04IXYXqwqXol/9FJT1VS
nLgma03O7Si1wf76pF33uDPMPNrkZ09XbfH2GzcbdPqhXsLIAkFtCCC86N1rpPU8DyNnNSoIoUbJ
FqzADB6gFjc309lerOPUQE/4QJ/jEB520HWfUPJF2GjnSShTejSD3R5TbuKxmaBMM8LHmVyoksUb
xcUbrBzVQ+c02DXQddUiZdW3Oi51jzEunpB6JznZ/eG4/9Gfc4zyBdZJh+dDybwSup4xBhBxHuMY
8SfGsZV4ULYMptOUsy6Mrsk9bQ0V9Ww23RqPprSzZpX8f+GuygaZpBXSJTGGfLyRPDJeCy6dQn0R
DE4ewPNfquCIZ6uNxzzhXa8RPMBwdTtdQbaI40WqUDsrRJtjNqlC+6HFYz+4JDZ9cb2HvkI/vfme
+5bEmvxwsI45ZnQv0VUS8vgYxAsovvrJev/OhHFHsZ+t40VPjAtfEK1tTF6qPlCRk5cbF3c8ikUb
Nx1tes0Ni7SQNbJn0SKCLPhj6ftETSN+TSYZOmCPgAUywFTQ4ft9ymkfK6QTrv9Nc+GQX7oVeGCO
HrmVlVlMjpTL9CVCNHwk/6TKBUb+8FMpVb7EBCqNkwBm60t3cgUkRpdhy4tHxEXH4hfpqcElyqX5
MNgCfZPSsX2m3YZG8Rzx/2eVpbrUc/0KLEWAlNk5C+Jq8kJrW+Ek0v4iyUJpMXHqA0gtDMsqo1Gl
DcoyLHw+4fKV8siOzWtWzDLdo0rtBQ3N3hJ73heVhZ20y9e92FaKdQnAyB8FyxhmT1vLwURjHguT
Ma/sx1kSynliDeL4IShxOD8sQnrKuCzMrdMCI+9a+LDa0PY779PJWTlqrTht9sYc+/Sdal04vTVf
XpTuSVeX2idIMTqiwyC6PSFZOIVR7pwoKE/p/4O/XVzME4STbcViVM5HfPyUSLMUQ/3eS9J7kBiJ
NOxqiAIcOivRio8eGx8FAYXGliGRSeS1XKSv1MdsTelPKKLF3QZLHQGoM5HDUYG9Y2hMcxgC9Fvr
JqyG4PbzLoFT6HGmU8XnP1mLQm3bKipr/iJobY9pUsWVIg6/FNMSMOtf0ldL2lD/jElffaur6vrm
dkMxQznQvYCIM3rcaH8eGYFAje8GvO5ZrsRS+5kwkriiyTEaShfb3Do2kvs8Dvgtm5R+Aeq2J20y
kfW0qku2tWaXoiFFoFg5AlCO49ft/mzUkhOy+lHOqC2qp4e30jD1fjzQP80dHGfFwkBeGZOk6b8x
EKzSuYMcy9uplh219A5if1KB8Y9Wk/NSJj5HEdfbFa5eU0nJCW5Kv4ASybDsJb+8+wSbLCexiVfy
FzYKQGhN2G/oXs4Hpwm3QHDNNIEF16yW1aY33phYm0BqqJw9jdlHKocU7wJ4dQODetDsAidJLrNG
39VDli1MscWzfgfgu/PddW0KyDd0M/rmsxELV9fAdBWFsLX8+eWLFLXltI5zMQBcTSKFw8vS50Fs
yqkUddDhKu/UxqMx1itJ0IGpJgbwWagNN/RO1E+2gDCw82E/HmYYEYGerO4yRypyq6FDEmr6POt3
F6YepXh3wIRjFKkgqXZsB9BwWDzSeu4XFXJG79lweWwzvrJ6L5KU1NFte7IosEZgyaqi3qLsukeh
Yby7XlFFveX2KLbJrT/J8VjYgacPybS8cNV6xiskWNLfy55lD3pgbwU0PXvIa60wp03+2gKd7Lod
+QzQ+IZqxtz0Pea+rq2AIubLEJVQm+0knoIjXcXOcOAfIhD4sriNRmpGNM+PP7TPLQLFhYf0a16d
WxVnOYdsfvkPdZquzXQXvvEpV5ODyXxAMDh7QWr/EMKz9jrQ77qVxU5pIBXVIZHTzsJ6T8+p2wG+
GxJzojZh1TtigVponD4iqZK3ixK2VYVnc7PwW2v+qk1vtyJJ0ioSxeL6qRjIsWv0XpS8/QnaV8l/
MpwmFran3p69/zwLTz+iDk2LGRWbODPVho6GaSgmhZ9+HD6FLbIUUr+6FVDeaaQqdmjZA22yloBp
QKnwmn7wXSVYh6k+WH8ipJqrT92KwQ7AdnEagDvxY8d7v3OzfPYiZnazfWvMU+N8aiIxUs3eBqNH
nRprb6pU12KEZx3O5SnymboplhRhQ5VPEJL0Bdh4zt6cfIRhLBVw0twN7XbaOjwmQmgnQVJr98J5
7P/UIN1WMzRMxAygKj8APKgy4czjZnE+HgyHMPAnSpavAfS8h+o4ggPR9CPxD7l7wjPUqpjA9IDT
dolhxfVweMnvVQe67qWTywKDdemVqm0uqweLfunI24fALbATS4tgdTYGgZ9nKta07MhJX/q/9PWq
0WGEvbgM4aMOu/YW7eAJnMafDWaVIAH8W/jMPQ0tAsegVULesI/wWhm7IjXWym5QXvZEXK3NeQPr
y3ThzjLUxxbCw54f3P3atCQ1+J4YqxG7E+eNXI3iUp74RNLLNx1YlbHil8IpKp8wa9p62aOa2uxk
3dMfBDIgQEipg6PM3Iiskek/3MGuGXuN2ZSe2DE7Uh5gOZewR15HzD3ZuSCFmTzuZJkt/qym569Z
chkQb0M2cEN3rKFUBQFfC+Kt6xmqE8VYOYxOlthvVapxXU5mWxPIIIubA//sgsjzl3IH6hwDWiC0
Dge45hQLel0XmM88hGe9pKFJ5XoeqmbihoTx8FpsLLWNZkH5b7lBNSjlL1ENQi4RDt9HaRzt7vuS
W4k/9MllYxQsOlOpcbnaVmh8UkMofPx33vnyIIhyUD3epezkwIjkXQhQQuaNYtULNwwMQqIF+Iz3
gAWmazEKaCA7GqRxqhLVDy6Dz/xNR5WlPD5cz61bAs5EBqCQcMzY7U6wD/fZ6F/hdFLfAeR9Lcrl
bJTCiQsym+xPsaVMTqIPuA6S9+y3Zw7fgyqJ327icR04f+WPmvX2nhhzE7+We9apVXhUOG7rLj4J
dHub22NjhWZcLvU2EiPRr3nk59k+Sw76rssNRdagxGXJCMwEZAF/TXXcxKBe1mk40FXupV4pQ8R4
782r1l1EtZpw7azZvwJpMOjSt/PdnsbtS9EzPUpcISrpq9G6CqHqKIRZ9ZcvH8ic2bOHaLpWk+m0
qo/aimspUyQTVA4T9FFRg1TWVR7695W606cdIEkV80gCam0QnxT7cLKrqX/7rWX8q8/UuQnY4vEf
1sOdaVouMG8a8QAL7dZGaDrc5MDzZidvsJ+EW5S9BQwQhsNG4mdR3jrVT77UbEMLWMc0O0mVJiX+
6/Mt0ELKGQcQOsW+4H+K2u4NfYZM/12Jrw2jCYMhyTGmGX73lz/LYilNF9BPFwAkDrv8KKNwF/kQ
bGAeXuPswK5GVOydjVoC88cLccMol915Db1xKfMI3IvuXCtcxUkriUEU2mcuO0z7TNlg/9p4Qn6o
mjrOi0vgyY768e/Or10kzENzXogLhinY7BgiwbD+OyJGdq2h6UZP787uJOxCs3njVO8mJhQvS/4P
VvcMeuGcBWU23ynxhUGfWTKoQxSM+cJbLHShlqqlE3ep8tn6Bb+x4G3InykFUD6fZiqXgdYOuj16
huSAGpI7AIgLeWl7q0z7y3WIgwp8g5lrbf7LwLaeLuhwN54OtbcK/2VR9Y79Ky80md2lnwR3xoGZ
EmOd80MW3O7qXUkt7qv5z53xvFv6rUUqI0bztEuwelpRh7S7d9mpk+RFuRRI/5wmxoR6DrZJc+Pp
ZEuO6DTMNLilNHU+F5VOT/CnLFWHDtoTq3YZTtvb6p2mrEXhq4fqaGHfrSiRRHNdE1zeeNg7jvBJ
W3oNoZLcxPKyDnuTON+8Dvud3BlC2Pi8bTRlzLnKg45F52/ArJljs8IeRRqs/QOSrCFOBAF+sYSG
bARtHolNYvfFt878UesaPljazAGM0Ja9hPD3bdGbg8ycMNPvyi27Dd0FhE5iicuSfLBMfZk/Kf+D
OP3nGnDv98/Ey4tvUgLkXsF90Gp3Oj6z8SxTUELKh0gp6dlUZZeefSxSPcKeX2A45Bha/lSYt+cr
EhQATJ5tPKXDQy/NT+rNG6IfyeuOzGyUAlVLXldJqe8WAArQxeVUdP6BWDMb2q0VxqZzQS8ZCrza
sVvpZDFu3wFxeEMKRwEisGrSesupDHbNsUQn1HObZmZDd+EBdFq1A+XDjbpeftpodoSZvndEOLfC
CA81dvJESQiB1Jmg06evG5+jcgG0Kjt3HF+U1X0L2ocMpfsG5PfEzi5KQj5rSH5+NyNaQygrWE7v
92bIuQJyCu+ge1kgPFu/P8XOLlnknx22BP7GjoHjqTPWQfe/7siiihb0MlHOeiRai+h974zgO8oq
kwv2Kv1VRFb6vMwakSno+99S3Q6dR4ll2z4E3wWbRYSorvm6OPJY9vhmXoqCRgrDw+WPP8mWHP8y
UipUIGHZf0vKF6o7mjkYiXQbIEbXn9WA9QOKhC2cRqD2ycqwfHXI1Gua/DTdk/YWiMiatMOgw2n7
JoLve+58VPyFmiiEubwoiyG7JZQZNCTgSHYlDrSZPHHZj1zdAIqzAr/Ul+OZOCrutihtbVvHwBDs
VK9bnPybOtMHwu6DPBRXRpUlPZqQfVwjswSgQlafsjal8Q0/8nNkLZGUi5MNU+7hyplIRAFLTJ2K
CL8FUKjT+vGKrFAft2fY6yBzgvs6OiR/J0MGkVNzAqfoMwFjbiaSHZgvOaLhn+CLmBFLWo74Ffj+
Cr0rEM4DwsLn46szsO+JGzoz3SsOAnNa+4H8qqJIX3/JzNHavzVpbcTnT/T7JxMAUDUnWn62PFvk
E0+f6R33czTkDLi9gX60HF58jQEeKbPK+2B9mzmN4QAy3pcdlSf8IFAKEgY6em81XHISZtBrNq/X
0H6z058JmOlU+fItW+xBf1pNYsUP0shbPKEEJ3RHClQFFhHhJgo9uGY2jueSrhs7gRTRNu9yO1YW
VIQaOXEF2ihvn79NrLRbb+uvUH/DH7gy6kmryqsdW0CeBgCSEYvWrnqZpbJ9NwhjoDWggKzToLbl
mzdMMKuXOtu6k0e2YcfR5UQ1+Gf7Yn0dJPl01sPFXrr5NCyobd3iC5OmXzj+rh1jAEu1CvV0jPEk
YIHchOXnRVBT03GolsEQ/iUHLOd2+ohHSjR49fWFTL8JkoxPCnXnVbpDpXK9T+4ck98EXMCxx1Mm
wF6IucyyLeOK4SPEs/VlLa9eUlJVZSp6OFS5D2afmNK8haubPKvwr0U1qft91gblNGxNR9mEeVuZ
4vKKUX28/xTeeXqOjuoHXAOenUlv9Ma7nlggUqgvJNr+hTww464abzFm+HsJLAO2HbSWOOqDSF2m
ttUaNK6zP/u5jzP2jT/89kT/wQ5ofBkJKl3Ph0kK2mDPzM5uAhBKMeBUmL5wP+z7+/gTH5LNWb/P
C/TEitV8US7BzEBiqOUnbE94s8KG4ZQPwXdYnSEH/WeQgySJUYnICjVYI989jJGs8/vuq8ZoYRDz
3etu2ZEDy53MqD7ptYZke6uLh6cH3SN5ffN6YGe8BAqsAY/DXEToXvcuVaU4KFCp/ShGZ/iSMZdM
Il/vRlnWExlN1LSNcogyvwZ7m92Xw7sDmjVEQ+2q2ylvfOIujSlKcoNjuFt5t7Vv3UdI6Li4/Lv3
MpeDE/k9dgUNuIu6lfVzV5D+P0aBaB3+hGR6U1nb+DZL6o20VJdLMV2ZTwBmLKwmSvfHGcv/khpl
ASqz1k58FWhih9FrOLSaqUqz6RqW9B3fW2zFEe3xNEwcSWD3ANI9SmMK2r7a57j8f3uWpVCr3oSg
pwVst2bPJJHslRX8/KZ0c2+Qa9daJdYXdxiLYZPIWI3mbvWlDNYRcg8DWHIrlxA1lIy0JgH4Ixez
+I82MUrVYZY1WzSJHk8lL23vwdDoyFzzwf6/Jnh2PckJ5fZWJYQQ6F0nTcEINobC3eZ4arpsXyFa
1XGU4YBjATWJsl5jDE4lEqwpiKpaKB6dNgYYqU0eoIsTW34Y9TNm2QoBjlSdxYIpAThR8OQoy7ZL
LkSriMDO/8boQ9qB5e9VxFqqyJNlz/in9ferwau+3HuyGIp1kq729LEoNOl4o48EUl6TeHap+kXd
62ldkwak2s6YQ4qR/pwzP6wrNdl0X5pGev2a6wcSTVYWIVFOPZ6Jtg0n+YS3oLd5X8FxN9tRdJVy
9P0ppo9WFA8p6p4XtSjXzD1Wn9IZIsTTtczR7CGT43L0InW6TJJROFb3t/7wuryD97Zr/fFA9cn7
K+WGNs2fGudwCZy0pwgARvAU2CFBJFEbu0t2h3bfg1L0M12YtjbaSklxilm4NHxK4UbixmmTRx+b
ZNyskjbTaoPSKeJOd1M7n6ri7kYluefajTylPiqpS655Wtrxg53Ae2KZzZgrgVCs0b694LJL9j6n
MpJUAOex1m7Y8bGMhKl9E/f+Favc3Of0uGv2N/PKfplpdqyRgbJSsBBLun90GgNvjTOpGdiP2MoO
uCaSEET8bdyA0YeDzg+ObrPeaYZbAu63G5m2NMpe6GK1QNP4s/tx9DJTamz2N80vrrHdh2KZ8duG
8OtvFr2ExMDkBJ5G/rQbuu2UU8IFrqXZ4oaAjc3gq/+VDk2VabKP4b9LCKej9Q9QsDcYIdcJ61JE
/b2pAACzsHpIvHBmHJcZdFoPcnxQFudfhF6DhB/Y507mLUj/08GmWfV6C4rfoeCxRg2890shEY4d
PGkN1PPkhPTuUOy4D9uxgnXeIpIMkR+muAPFDclrOv6tgXQC/2GBPu06FP9ZHTYbUhW23tvuM7De
5Lcqb4erHgHUzixYVPmclirbTzHBcPP/KrJ4BekxaRrm+qeRe/1V7h/qLCWXQcN4X9jK4iQi8opn
Wia3JCzz2YK1pOCDgCHXYUXZSDXDWQ8PC5dQg0adpTZlxdN597K37FhFtdPQjAmbCB2Tol/tLAHo
kysy9z3l05LUmipB8CUrYnb5ZrK6UUMzjqX5BHYRoW/5ONMfs2/w5PeNukw5AohUH92QD/p9iYav
cwzjYwT46si8X2juSXQTN87GvYa+YVU+p+POFvo8Mys89kmLvQSf+IjdUKKXRYlgTov1tVDJHm8Q
FFVVpKH7jEmAEWQ6gFEaUQk/OCIdO5WQh0ptFtOOGtQhJW5JP3qltsMj2uemmV6FyqKOFUGkJso2
hmci1ve1jzsTK4Oqx9Gc2+kswNeV7xijtzj+m6YeZBCw9hRGeEi4cJzZL9ZJonw7C/6rhzChtyuQ
/HPZJ9mH53FOAiW/smufiDSmh/h6m2IM4EUK0KZf6+QlsVNIE9zYhl3zuYnwyFGEce3O80VhjQDL
uku2Tg7r9C0M3rdxj3iG913HMLsytJVkJOZUkKRO1fnleHOoENqlRL8VtF5WyEC7talAyhVDnT6f
oXbq/hAmSgPsqMd7gfMmLkzIbU83316CwPQC846WF9ZXbF1UnYmOOzRnmZihhKkIXgxSObT6wLGS
oXoCNYvsnWsVUWvwhrd+kmlp6E2KhKXc8yFULJ8P0fSNrrfQLWTA2xg3WoQ0VOqoK8l3thqclQDi
Il9eqnxFlOye1C5edAnrAr/NKSrYQwx7Bd6Fb3LPRu6kjtmz1CNlARTbjP6PEk8OXv3v14C95yVy
0oKMQ7c8llPij4J0YKxrw3OiSodSA/PVZZvadBpBQZnNRnj9ei2JwSCebXEhaS2Oy3u13J0+msIQ
s6zzQP2M/2+sqlcRS+qNLt7EXoyBm5Kp9Ra3U/JjBPJz77bAW9PqexZo/6FhmxNFsMLhmLHM87qA
PsDgjdISvTF7ky/XDOKLgZpJMaWTfXSDwVMqkGUeAKQSzI+/e2Y/afSIm2xRJNrtA8KZcNsj1Ear
Edl95rDujthYpSLJaF1A4wf67PHd7uRfwmrWVR1ZdNNt1bdcXzdcApfqRWAW9DPrZfFj6U5gnG8n
YITmleuWo2jtvO3alxD3rN/jlgRBgIgLb7/ivpdIRWVduRbaV2gNEzKGBy+hGCZXI8QjaaIZt/r3
TDHbOf+Dw5XqrNUQoXm3ygT6Pzj3ureuNIC7qnxalJKEQkwIU5VNUlA/eVHGUTVXB9pFNWKVXk6K
3XoFZNhsUm2cWA0I7PcThuXGPw6qbTZvR2i2xDoArglUhl6JQTVI3Yb4MaTOPcmpDPwc2jmpI0ng
E9jN5FY6NnxmmpoEtLkMhE50UTCiG7Tafa6pYjVlcA6WnbsOnxzV4T4d/Kp80PikMGI1jukzHyOw
3fDAM33ZbuKwnJWiIgluyKIK578+kOsbWJfznEiJ57MEKVq+3mp0i+e9hYF7ld4fSiPhsNil12Me
9wLuBxpFEveCl8M6zbhHcJqtKG/THWLSyAbyvJDHyDsP5ESo3MpOu5/pJGk0tPWjl8tqB7QW0hsQ
Dl3QkbDD+3/EXCCDaDFJcoOwyoCervDKQqVRpyVoHJzRGzKPWAM+pBsnPyvUXlGTT5yy6WZJzjYV
MvP0nAgxLqj79YzPYEbGJKxLqru/CaWQ+1g5nR8CPmD2q8+MbjHmxBsgUg8e9x4t3F2CQIEktsoX
yFABPUTtIuu3JDnncEW4TQ0hQzivHKFQzyhsasf9rGwCpQBDaTlAws73pZZZumoj9iNWY4ypwAS7
PhoXKYdS4gbRjeu2BqaJ2ykulMtshTzzL/5FQriWn8q8+Okf1Wxy5lJLEzwfNV0irBrbKnJjG5Ac
RKER0demOMxv6Nj2uZvS2kkJNdMyZd5I6f07DWVtBG+kro0D93dynjLHqhlDDNyc+5QjfPlDIR24
GhCuw2yuGxpcq64U2JPD0i39/gjOLCX3swxPHXkmioWSIWM1dc8dscKO54yKJ+HOf6FYhUImSTtz
tflHWagbOIquWLcbHIkN9XZslJsfMlU1jwwWVLGO+l5OeRtqfwpD63Sx0a7DNJztMs3FHxO9EfIL
BQt8O5AbjGRAAjxIWqcWnLk1a8LzaZEBLddSvrMREKDI2loy57BRLCx0PO1Y6lC2t2sQLN1DW5ZA
lKuapsRarbaBeFAo1wi2UjT7v/pwovf8xajNbi+oIsHyaYZRk1Z8rYI+1EWJQuOIbG0MSuMUaqzN
MjKjPURC3l83T1ArDAsIGgORmAHVXShEIMRJWjnCIRDYH+C8oW7jlVZPwG2yzNvOhEa9ojOUbcAZ
1g6TYMY+uvIfWwXHBp7zU0X1BKPxzhRM6cMA9c0W964Gs1van4mWQF3uQsU6723xBKf/Bdwj0348
d6t5fIwDdIjccMQwAVYHrB15x40HHTyEc649BOge5dN2/4LxlE1DDKgFVwX3kZKxdCfyUlTTzkUh
zxZuIlb1CzPR+me5YJsT6jH5wtzCuHMpvo5c0UsuG5Rihp5VUDKBW4Fm1OCeSRGIUg/OSUhdg44d
+sR8Zd00dCY/m1jzag9iYXzFjzk3xZCLv/t32NP5KpALY9g4zeNTPQsdESJGv5Ys8n+oQQUHMQjo
Ese88sMmHQBsIIfM4SHea8hHvraPc1filbzOWTWIL21DUdJB1nxDLSR9h1Ql4vsCEllJTEZC3yRw
IDyj+kpKvxyBXC/C3mIk6R7MME3wyRQ9pI2HMr0ndG1Xhh9WjJWJ2bLsxTDAz8iBDOYI51gw+yK0
oWKlakZsnmEYCvXj1pCXlpMzlWCdeSltMBY7PeC4KH10wiUN501tClsb9HYDsDLhUXA1C4H22tl8
mMeLPrR9lTf36BfemZgeYHtlQLI8ClRWceOWNqrlpdF7Hc/rNqkKw9/YNgxsE3qreRAiY8NopqXP
SfL899XpLM9NaI0yx9qjY0pct6bbRuMuXlJU2LenYKkACffXTt786EX+gm3DWJDrfJI2gXE/ODwj
cqvBZm+fx+adVnICICaBV5wYuB//7xKSLmffZu5mBV37D7feLBedBgcAdoFXulPI3VHZeW9LpZSC
oO5u44z1JtFDoDNKAexmoG0D23M9MIBVBKfpe9bu2ndIjnJJm0j7oIvrO0QynJFTzQV+IbFottmy
lO+7qOYOW7D0j66RPtFLZiY+LahrqB4Xrl2jFMH2YGBJwdBeDnUeP6qSXq9zmZDupOECOHqhBCVS
fznnkTXcHbq2KwHPiIQ5JmDWzJbJq56U65gWLlRchZGhtR1KvYHFVjk6QQntn/n6GShJ6wGA5hPZ
51m3lLf36balkUcMcnduoto684zXL1nw8tWy0CuGRnj3nd9AiM5wuOgQ7yekOD25ZBLcaCVNlvs+
R8htfLO+FxlGSeTltMFzjeYb/DhFwqU4UN0AC90XjwReONBXTtDC358JaZsz6v7i5moW8ccntooi
dWGDJMwHgy84VyPzZSo4QuuZUT3qYB+vO5TXENS2Hsf1u++3kaVg98toZQZ+2MRSCuws4uQ5YIsl
t4KFBsORJFo6g9Ran5txe+XkKyb0RPib6fhU+OzAJ5IsaIRwJqGm6kCZCUASa3zKVf+0i7qkUy4g
iPOVDJH/bscTTt3nn5Jgck/GepeARXv+YuRAtYrCl8vablkLIhJvfAto1JNUdi5TptqytvotX+7H
4PdnKZZN633zjO3dSTYoDMmc653PxiWiyfaPVRarA8vgl3AFiiW12EL5UaGY43hZQ3trXLGY2rvU
1vJGRzAHvawH50PqYN+ujdLsBEBGRpXsVIMmHYvyTgg6AWPUruYPYQ276lybvtfIoLs3YufssX4k
o4sEhBY2KIeMVIvnF0UYLUt1YWecxCddQlxI0PelpS/IUdIogfYbjXUGMmYvIV7qHJ7Q3lSCzJcN
UHIwEGXm0p4p7T6Nmy6zxou0IACUg5Pn+fBLwZoxufXsj+j+aacwwoetFbBKrmq+/W0NF/XZZW4z
UQ+dkiQBfsIJTXyzI/GzsBFr9cQcHXhJcz/0vISE/HPGqz0PptmFls2tI7qBNz0sSUv0e2Ie9yq1
6ht0/8IilPMcvc0jdcQrQG13nUkYbwvcX95sLXIuvEnzcelyuyreQe5gxiFBWZ5TXb82JJbM9T2S
c0JPO9BUEckuBV48J8KlKjnFU9qF4PEbhOUtTo4+zFiA71ahMVtmitRz7vQPAnFnG4JMcgTgAxVm
Vx89ap98xzEnba70G3i9DiYHSSukZa/8HZaTirA0ngGmAX+5Yec7UpMfuo+lFrjc+XDzNLcBZJfv
id4f3E2Ub/0epk3ElTONVQAbpfV55T3j/QMjCxjb0RNgv2JIQXe/si1dRKIMKkoxZSEQvhcrj9Rd
D3Lu82Sf9IfS7btud9jAyAv3bGiI+D1ghxwG2fdfwFcwLjpv6Se835TrkexhznWJQtBGnhnRBGua
DTnOBcxwxWW+3DVEnfCjUyc6Uh5F/ylKOJX6tu3qAtQhAHmX6pxBItHHaU+cHJtzG792/6wcy/GR
qot/q6XD51Z4DB4rMCfDPMbdwbE+EQln/FJSOJasy3JCji75njFdo4apnPK1LnAKeDGnXQ7xdWq+
1dVRGuv4ECxtDh3OmhOk+KHh7Y5lHy0mwLAzYesiXwKL9L7BSg7RxBFUES2gbC4IVsEZ4ziDIKpb
i7vCGjjaay15JWiWLrhr+JcbO1YKNjyW389xxJqT4MWIQFHuwg155vKNAt/6fGJtYqqX0fx3GcUY
HuTeChiFshNl1g6FM5Ggvh4eK+MTUOZ/8P6uL3ACcffMJgFouAgHL6RkvY2Ec/1pbVPd0Bdz1hwu
Y+mHFpB2sMyjnp7UAQ0gbiedt/TTgwI5gLivmCEK96PUhMMsUgLmPYPYYOKOcFAXrdWA0H4golgI
heygVt+yZ/zm62nLrRw3HUevQEMWNLA9DEcG7Y5pV7slIEQSlUp/acAE0ldPTJ/HvS6oBNkfLuSH
v6txQoMLhyhvKM6TvN+rdJarTniTcGVHuzYz2eqMH63leUoGCiwcHUWWWC7Ioa0alvqAIORsl4nv
riZhqnfq/dFHXwQKaJajz4Ia+HpF9cG8GojBT0MfO6HcCWaB4x1pHIQTV2oy9mLFqNaJzSNsT0ac
RfP5VBUTMn4zRcM3WHue5h4lvrETC2qZ5MuLY0yxn6h8d5HO4riw8Vbjl/iKZ88QWmIj5LonueTA
3gYdvrnfTAnerWFbBarYd3VgFwaQiC2OQfjkPcI3MGOMP/rQayYHOv64mWrgAPYV9+9HLpTrL2yt
U1USlxsSkVux0gvoRwKlMWMs5/FRGxEahLekFLUJOIr3MjTdGzDcJc/a0T+EpBMQZSEpwFyYby6/
d9AHQ41sJkGN6Pq4CuEIRgIlxOzRYIaEDy+sYEF0ArH1GmR+85U5ft8JcBdwl8Wu7DXIwBJUGVpN
oVT4k6xW0N1wXQyegSl5l+JXUN9XJ5DjWOpoNr37SRBv3Qphmg0XjPtK2WWV1qmPIENaMuPMQnme
/2ShWzfufpW/cpQtMMkXqZmToZeIWhTO1m37vIdSgV7I/S+i/K3TPBYjh2AgLAggy/QQuw5CPX9f
JcFG5dgKD6lQ4Tc6RFsfEux8XReBiJ7M+mwoqgs0CSnmRaqsGggxgZ127q8wpBIkGPacfWau93vc
sFyFWJSTgoIYt+cAJJwiHxoo7x20mDFOfomnAl8Q+MHGxSYSHQJdUG0NPoSwilnWMmcqqArsyYjO
qMmy3RJFGXAPnHy1UPetKF3pmn6tcKJ5lIh+cZC7AeMiWU5LUzFpFS2wxS+YAXNS0stevlcyI8gY
/AAcsRVwQd32PQcqKM07t6WhJO7A5G7HK2orJ4BpUh8KnxiuCEkTQQ+cMaQZ3T8fOZ3GupO6Xu4a
VU6KeS+QE7pztE5YJhFIrF5xZarGLskwX4jNAAHYywVHFy+Mqd5kBP4s06jpvHNV8ZgvfpfnFSKS
Io/uG0jFrBzEPb3dTZbsh3wNisujMB7sbTFaA44Od5bpYl+t9UvsbjzNtj1BaloPst9Bi2WNRc0U
Rbp7xM6mPtQuiPYuCJaeBpXk85AcCnJrCoH6D73LdIh0nhIAZ+BPwtRk84C7AdC3nUPdBRK6Lyca
bTBSOQZEYa35WTptJtGJVroHqRo22JFdYZJgTSx3GfeF150c8trjqjHMmsPpLMWYq7RtzjB4UcAO
74D5gKLfdLBQXmIztDxQQ9uRMoOQKl49e+1N46WhNGxQ10BhGz72belRUvJr8LY/I5x2MdWw3xY/
ge46faSCIiAngU35OzxoGzHhCjtcr6h/G8ZMO20/HCnVBSvZk4/cEodrOi8SjuwzhphSVWHdNnWL
/IKtcEzS/dD1niTmGnhdHm1C0vhKoPyGLt8ceIVWFOSjLh8NHgjn2kBumvLqCc4KLKOMYMbscCFy
Im/Y4SNo9UQ5/2O0dXT+kqNFSTuKphAP+xXtTwxImsoxmAE7oRlWdv9cvzNgY/IEYvbXKDvPkSrp
cunhljtTQwDJ8PxEa8qa/HN/fgTPFItHWl3aveOuGfWda4qG08cIFolq3vxWWdnq5HBxE2UDYDBN
TUrUk9C2VLekLfnbQ0MqWLd9ZyYk9PJCpdb0pcpN9mGWwOah7C1hskUaj2or28fOc4BeFrL8LOKy
FlbQZ2A9oJ4U1FehQGKClPTXiq+QQridbvxnvwfvsMqeNq/iE3plRQ9n/VDGY1py4u4T6TAe7AUM
EgJ46WXWq1Pw4CL1DItnIm+y9vYz+/Y+WzuwAQEeB0xb7FyMUetik4LE+qz8W4NE2y9GfU2zx/nr
oawr+N2DDklG9bL0UYjVx0QJJi5/O+6/XdzJBJZK7aX2Odi2lSQRuXc8mVQA6UlCBrFw6Z4rUafd
OHFTW0C9OR56LvYPEySNWDk5639BVoF+Vm6Y0D00A9If9Ymod4KAyVDOEXc6Be0okwvvg4NIApZT
s2wZdTa/z5bHbUo4kQ/JhHdcWt8U7ZfDpMVWrlD/DjCN/9KHqrKwlk6gaqPKAL0K11pno40lp/lV
zdWw9XMbYvXg7Hvh7BEt5jOjZabyuF8FCojGNcHILO/Nrm3fsBf+pLyX3qghVoDl2QnlA4rhWGzL
nExnPbEb6txt9YEwzjzyEYcNxhFFVULuSFwGBwRxoUTRpGUyWtvAtNjVlwIdviHNgRMtJG2+1/LW
jQ5zTDohQBm445AXxh4rlTocjoF5VhG69j6ZcSs1K3VZaeZIs5HlNzZGRgEdoRwXtZ0gIr4yFwL3
ELa1eNneRTUIryj3i8r2i5Y+frWWw2ORrWWMVmJPc4o1yo59uOVpymNIPONGMKFINc7tFhFY8dRz
1jNjXHfo//U37y9P5X/tA1pewbRnWz3K70f4tNiHHmQ7jigDBFtg9eaWJAyLSVr+m+6ExE/chmsR
K/wgykPNvi08hBmpTR3Bx4F1UG2/aUlj0DvQnhWUq2DhP0Lb/SHuBL5gD58KNTQhKJ9qurMFUuOG
4J90zeLbf24FrICl58+JuVQPh6jrU9awicN5LsEpv9OEMldsGJZTzLyM5DJVd14iMlqFDo6mu8q8
a+QR7V7UnxARhlQH3OvCHinX2bGGyXKxQZfdLO5p7afHbYRVn7KGsJZPR8X0oclHFBGVrpXORAHO
i4kApbTUasctWHBRxYZgDW6nhQ8woKy9TsNzmctvs6tXAv+ZoPTX0yZq3TYii4oB7V95MN2UK/4Y
ph5hAWLjfgON6go2bjGed+AURRz+WQqVN3WCIghCvs+LJ34b6BhjyPRHh/H3xPFHA2sDPqC70a5R
85v3OxK8hnJpDK4vIXDSu9I7sv+GxQ9xhIRE3nCCQjF21pW/cNH2i0GVr4sGbhg7ujYt2C6Ic3qd
fJMSHvHpVJ7UqcbiF1O24ZJ50Det7PgAhr8cIIfM4BPMltaOcSHuuwAbBZ2jyyob9x7DcJmtBZXu
jVAEaL7bS7wgNdRL8QQirVCV4ItFAqrhnBVJyr+x1Qg6k6LvO3FWAtQxbcL+ukwRCqe5YtR7fJXZ
hnBkbXMTOTDE8mL8uun58U3HArK/1d2cxLpMx5NtpXl6DLip8u+cfy0teVVW1RX0evvKZjouTukh
VtspXv7tUyXhWbCBSEjFxLSse5UiNWNfWF9Diccf0IbQsT5gsaJehkiyW9VkTApxgAKUArdL5pAF
KScxcWEvRm8L/f3BAQOg7nru0zGwrA41xew3NtoRdR54QkejmTffT8Qq+Yc+ai41UYsKRUq1SSKU
NyvzYi4Vuqd7APP2XGBpWDbgFAf19wc5bSqc4V9qZn2ToTDNGCzjTUH/2HaUlaT+99RnVcvO7rwy
1PVRY+/+66Fw+suImuFziew/8t7l/LPVHBrZSDxfTmvqAjbq8JNvBLKhXi1nHkTaI7wHAsJTOUcT
Ff0570gKldgXyjSQIhxL66nCz+wRagf2w0YwLZsIydBVinuHfuIzFS7Dyd86iqXwjfRDd9fPeLod
/3gMWalJdlssJIsP3e+7BTN5OTNk2ktBQYlvWZIO9NdmutjNneedq4qZ5hMSrE+dJlUUKiW8/9xL
JjBadVvSEWQnK6MyLwVqioH+Vogq6N5vqKqUgYRBvBT8X+gcGz3iD+OJNgwX/kMyrwGQf//7iIjZ
73AGbnf7xJtLoWxrvUZXgOmk1PJKyZeEU2VWnkAsiM+QUAJ79ROOZzUa5736oxZj4khdu8IXS8yi
8AW9kWWBFdaZlRACUEBSa9j1mYhpWJimG7CgjdmKMqxe7Xahp2HP7ZIM9bSDWYW9m7FIUAmkQJW2
AsPzP2QZ755NI98QEUSF78eUFSyd3w/BWU2BZMU5n6Dy4WpWkBinXJ1K9wiXNLH0kAbW0qSLdEOJ
GmpSc42w9YY0EgXGHH6CznkuX3rTQLmmVUOQhxXDzOyBktcJyw/2DlKqdDnXHw/Ez1GuyrT30L1c
ZhqD9gqFE70tcU7fE88X9e9YxHmcLI3ePrTYPSKDx4F60YpucH0wfA3aqGGRCeUmrRamaC6Cs1lf
EYeHufKV08xGRjcUK0oZiKQ67ZMhRBuiZwbd9fzaaRWw/tJGAwQzRZXKXhk/kEpo/VwjsMaQ484a
YzG2IP/c/PToudMzxIvXQphU3ZvkMQioGLhn9GkrwIAyIlGFz4/fRHTnKXq1TMVn0Y/2X+5kdOIm
BE9NWS4bdGwBe0JTSPMiUEsblnX//Y68Q0eCzjSwD6iwPt60jnfEYRqqJ+vuCfL+nMMgaYk6Q/Lp
XrrEhFUj/g36UvIIHi7hLMESemk2+8njLTDIYYePJ8gAUxGe/FNgf6GuG5Ee9BK5DxgPDkCit9s0
l8jaht5CqhZDYnlVgxTFJ1E5BXi6q6EHCYHautvyxQPvy7FWI7q13XZn9UaUdCzNMOKwpI5zJfQY
KF48EEz3h4yta/ZgcPHD82O2tHVNVpCrxrRjcAqcdb8i//PeH1sorX4U0Qu+lxziPPJ1LuavboGk
rLZkpm6pXub1H8AXOnfJTCNfaKQLGwlw09izLUze0KUaysZlrgdkO6YZj2DspdLlRlQh+SJS1vew
B1VlwEy5ylP21WZ1EzY+EGTc1aZLT6XIxndZFEk1bsv45+JqKweoQEMmmBGOSUUtwDm3kXaSVDwd
vhTP3uibkAWD2xFTgmSODHznXdBCA/H2dm0PTYvOxkOOw4trTP8XUHmJtQZt3XQeJ/wcLWZPteRb
/PvI4cLVNgusfE0JlOVFDoYY+1UlIRhz6nABDLjfRmkbMjNBmKDMcQl1WfICiRdRlCGAGB+AkxyN
J59ODHNE6Jsyk/eykpRSXk4x7BOk/jrPbtPZgsMgZJ/1CAsuW6975NLVh9JhWB8dnvJB1eIBIkDN
QUc8xlO/YUDv9IBBKrS8niSQ+xF/YoAMe6GUUW4NPXEu42g6igEmJqMZN3VDtNXRd0gL5mL/Y7Dz
UPX5UlhLc6jDix8tc9qCw/GFzcFCQvy/m7+ZJHB+RO3+aiLRDbaEyc5KOEIXOaqKFdRUuhYQv+lk
OCNvsEovFAnw30CTa4Ho4SZvskUwiEN6HCVFsuswiL0/O0FAh0bedolOxoAB5DDbY9yxIgBN4wQl
2K0Z3LtUg3RTLOdGj1Hut/SIkHi0cs1MgotEu+M1J2a8ciWPoBqHQNC+mbbMcfbgqcUTk3UFEnxy
sOcpEONt3Pw0XAEbiiy5fcFj1hiYjMjwoOaQGubJz6l6yDSChs6kkgapIw62WVJJGBH5y7/8XRKS
G3WsZ4t4iLPMU8cYtxHNeCsHKyHtqKf87rhzDYwZryDYFxyoWb3OoqtJMwtAclQKdKVOmC/R5XdG
KFMkEcPgOHYYVvMf3+gsmXZcc9Pjxn7AWN5N+30TIoz9FpkT4+nLl1/3YaHaOKh0xOlverEAPl8b
l6a0L+k0KVN8JH3h3b9d5uuuNNNcdBTeEz7x9Q86nm13hiiMgRoozy6B7mkThYbAt/hCj4iDiJC8
cTF8iCN9Kcl1b5vhvqRjSxj2Pln4meCPp8r8Bc7mF2uD61wTx3v4u2muFw90+6W7nJNBYG6umrru
E06EoKBXIgC9wO1enwgqBVLnb0mCSkoPfbrFqlFZ79MpjLXmkV5667uHwqSYYE9X/4mqAx+w31sQ
YzQjvchcS+6JG5xHc5wbaUz3Ti/tPV9ePA1ePcoKWUdOrQd0M4uGUWaqL4Nh6V2YXY0TGdWwZlCY
gcQbZNpACwYSefYOZb0fiG1oIPz4jfUvsjnuuHv1NmXqHRhopqjfMY9UCMTEDRjvIPxlbZYJaeQM
MBPjHsoqSd7V0xSIupRM/BWMJa2d0al8upELvhBFo0EAT/cQIX+4HpkGbNogVWx9/2F0kGRNG2tu
diI7oU9jRdSgWemqDkQzG/4HFr6dgvPy7SDFkLAqsnsYZbsZAD+6xiU8NVNUArZtl9c42D4I8Ohu
BrGYuNbLJpv9dnu8WKXxRazunJ4rrtplMaNyugFP8Jm96u3mmlrENVAOLRn4Y7vnlsC4jdWTwHV0
aOak40m4N8q59y3wXxcNjs0DqG/Il2Cv1Z7n0J0sebo+l7VtABzawKCmYVwYMAvUAXxuD+IVP6hD
w0gCFAb+LQcdQiJLEZC+dNOF5dYel/x+NeBwIka7MBAiNeXGKwoqCwPXyknYZjG9gyVOJcCa4BG8
KtqADnkppN+sSYxEoYNATH3Qmetyc5siEEWBuPE2TL9N4JtJhNBadKTbwwx4XR2ukFaZY5hn09P6
oQ0/Se3kpoWOX82Io5pXzVi3DTBOnTIyB4OXfybIEc6OfbZBPcKaxppli0eHEXLbyBKodxApmanJ
X4izX431aD/j0PaIWf4Uq8NhsZ/BsZXyN7bKKk6In9zlwDYiHtZABsTTs6ejN/FfFHGRDROf0ry1
Biv9R97Fb3/gmBwoiKJLALbc+2cnfY+MzJkxs7oSfrU+gzNjywqltWupBKl1HKDjWDZh1Ma/xQyh
wc4RkXJNb5UtHnmV/dfjqsTKOXiqPFaKl/Ro6mGRXgIAHxCHFicFBbs5sIrJKLNevLKIXaI1qFEz
Rat8ieZnIxfo9wPStna50mP03s/Eitcj+ksiNOq6Ofik0N2nKBnn0IpEFeogZuViWSEPDg2XLFna
cEh3bb2YIfHEsPrYuxaV2S+Q9tE8uJCjjxlFcGMAFKklIEAx+Fwyuj9eHvVcSfMHiXrg000dopTT
dCxA1ca9IaapQ9V2IZoGVdfvpK2PUbwWBb7J+y3u333UXyeILCuNufv5m965DVo5EggPiLdfbKAw
bYdfhGO9zpRJj/8p75zc9s0QPI+qEZPEanLK0PMY7nNrcsmbO2Qkzvw8RW14HiN5uQlFCPWx+6Ab
BeD1jMZAHhw2bP5Ks0hEs0VRoxK0D202gTH7VAjhgAVWGE9c3WJzQkcg73nhUvDNdqLZ0QCPKKkM
i65WKD726/zDpKiLbBMn6iO+6IPkdANhxvwxYCXS5DIC6GtjSObmdkqsfz9nlkhwrfSCaGsnE2A4
rSEg9vPra5i0r2eZFLsX2GlnxhqHee8ZQBdwk3ttsmS5NP95za2zYghqhjPoWLHU4rKc+7fqaegI
Q0oWvjGkekwVJVQ+iWhOtMAXGdqdSm9jnuncqoK47iXOjduXwlyw0TiDyJNaovf+pVUXuZE+ptH+
XIh6wK7a+f9IHZz4hsx67AVuesmSIm1ZPEd17GvzKtzLJEAD5PleB4HAowln8bZM5CakAGvhlepy
N41/SRY3RqBz9vjh5wxwBQKAKkGvg3Pwm3NIDiwAtg8/px2q63VeKaG93pmQnzLHgCDm/m3aqnDc
hH2w3eqXJRXeYLyCDULeQ5B111SIy1eChL6Bl5N5fspBzXsRU07je89FKWbaNzKYt1SNKqnLdJ2n
O4oFWdj6Yha29+qx3iuFrZt3uOaGGAi/ZY8lbyPq+vCTnrJZJdtT+aFZQpGBTbIfabXZsNsxcGt8
dgatyTcS/IjrSl08oI2mH6w6+JBErcmDNEqKTfjx5q+8Dm933wyT5iGmoD8hB59U+KWfTiJ3tdVC
u+kFVWOC2vGc+JaXwADXyEE+LaVDfKeMoewBGel+ppciTdzbBaKrLu+Be+FzeuMutwohSa7OEr62
V/8xYSBi64gRiLzqgzvTDmX+oh21A5NJ9djCTHp6ZsunKJinOkasPTKhdWusG19gsmv9U3mgN4wc
hJyP5AHJM5h/RBgh+vj5fbgZd3TvPnNhJtfMkEyd0FflGlzUUkw2NvE9xyDAsnjuVQKVs5+Wtl/E
X5VMkHGrnSdXOBeLDBeKkHSU0W7Ntn5XXxe5v504+nec5pYwDAq0LArV6/Kc13Cl4w9TyN2fkJ8A
BJXyMH4fP428Tx5iLTaurQn+1Ye0as6/YBTfE6drnKgMGTAW+hlDyMoB8Bc3JbSVfhpMTDadOu/H
MUrpXzFXPw2PMXBdrg6Tc0juSoo/4hYyK53u4JLsUj+kOjfgjgz/Tme+LOk5T7YOB+4hfQLE8O2c
TuAf1cJHmGTV5+0BGOtzj72ez4eFtYqHAzSKM0Tk4N2Oq2NfvaHtZCuf8UElZSiYA2UNn8oYSlRN
5kH+Ih89I12+E9gTom0otm3/CQe8UMZbChBM3y/LX6mxw/44zf6wUS5Ssyz7UM1D4b+x+rrFJf4Q
dnvpn4/BxAP9WgmUonx+BYet3digc16GbXZ4+7llFy7MgPbV4mSS0iy3StFjqLJ0e5AXuOzVvf27
ji1OcdJ/c36+P3GzEg03KppnePuBR1VKqBZgbj+0QyFA8FznoimRN71qquv0n4KVZ89qUUU29KII
OsBf6gUDUNKEgm1/sRvdosQudu5KJyqEVGfRU3880OS8T9MkC2+lAr2DtFSsxuOuHgdpLsz1Flzg
HrDVJZe8Lf7IeP+XJLhKLd//PJ8qfSTBdq9EAC7GbtU+PPZKFHFbvONQkostxazvg8eGx4RyR32h
ywbdCkkNSS2g4YRANmc08YK3VvXu/ZMrXRRTbBSE0StDfNYWM1N5LzNboTmPeCn7UcyHNIjS/rSI
fmBqfnlAuzkVxUcPiMlLnjzW5xgpNdhob0MVFtRvEktQM5zXvuUNQT/OMxxOn81dg8nD9if2lBxD
JYjt2bVeUCY5rkqVhbEp213WgpXcx/brF233HGMdYfZ8wwiEHMFXPcfk16HVtqqMaE8pF2IJS9vQ
UFAjpH0imVgE8xa5641jALZsBi1HD4k+xKqS8kzx3K0XZD+5kC/xu+AQ1frqmauJeDoKVmTl7jOd
6kSzropiepI4XUv8Kn4E6/2hZ9fHTxBzKxgg3FzrGZJnscGfmgwVPMDIemojZgxM/y/xPvG9WvHK
xxf9kOe9FqEUu8DyBQFCrK4hAIyfNqwnXlwlgBLCMO4Vp3xrIcGnCTJvd4TtmQeyBZzFBiircXWu
iHAQU7PifcTGUmGV+NW1qKxBoBU+qjpHIhHLMBt/E3OtSmZ0R9FN8bIF56sbvwfzUN30x6GovvRY
UBEo7iVKgVYFu0VZ080yiFYsyD6ZdYbkQm3T1RVV3vaXbjBxteTj92Ja869HcQH3JuC34x2yVBD7
UmCcT8mCAyyzzieiqbev3apW1hrET9O1Vb9Gpa4Vv7g9BEF+jAq4o3jvQAy0iSH5leoZmxgO/RXB
SvL6XPSZLmkPAcEwJn9tDNRp8XSbvv2rCaI+0w+0cQgBaS+H8Y/hvBqzfYDphj8b6/0exjn+PcdW
wNLhb33q0x7bFwNoYa0j0/XonaGKvDT0N8RmMUGkVkr1AJIFofVVvMkH7ysjRuPYcYKTqVbYz7DD
6wnp2p+f1O9bWJ6at/KF9+ynpIchiMbemIXBakFhenucetoGgmPvnQrxswWggC/d0e2qQjl9TMwn
QZx8ZP93zruxpZL2uxuNoQe5rFuvrWZxuahM6beCk75a/cE/MbTG239KAU02Y5DgmJKK3gkyQoVI
P3BgjBwiRMUa+08KRLSY0Ax1MreFONsy45sUkIz0jApG2GJYSnNqLIycx/5HPIkc/EQm6Va9baiX
4zb7Et2KxuzZ/BV95akBLt+fuixEuJRmE2I5kOyOFVRwYZhRhi6RaXmILCN8ejrBLSrL7ZOEUz0j
IrtU+1OPwYQ1j4qL8CJaNcW7qeNkL5Jz4avyImA98qUS3qfXdSO1QH4iF/8seF3pJvAcYYNUwQH4
23RiWzphFJQcxGdh9kzkBX1+2x53Sppca7MQFjao/fCsh11hfFv3wjtyeJsHQr1wfz7FKUi7OrvO
NFDSQZzDfwhO9FDP0woZQsKzDnj0pr1WEr36kbqjF5EdxlSovJKxOrJTPaNO5mkcnhOGhmbk/af3
vbOQL+4lJGFDsVjQLSTmyyRQQiYGuMAM8RYtgG55ndK2sgs7/EliBbP+lrnjW3fJtiJDIF2HmqMD
cnQas2XqOTw/p60UNm+tn4+tWQwKhWo0nAGr0FdzTpbwRjNIFF2ygkNsD4GtF6iUcMVYBLqwKoQv
fV04+iV9aJaGBhYYTJTeOnN9ISGR+Cv2c0/KOk8Bf8dYkWQaDiJfMGz8OvyzX4UNWo1MQZvtYHsu
qlflDYsCzg7QsT8tsv9ciNjWcfZlnZxrgOdPZcXxAW7WNREhGSipkJFvTnmTWyOW5ZosLxZWTDzj
cCBERKA3HbeHVf6iEy/jN7UhDdsGMyyc2TtU1wx7t9Xrr74umeluqhVZGWyJu++qwp6uKkIru1ll
qzuRR9RKfkYBsu6Ng8prvdwXYyCfqTGVxaHr5bitxgCQNSl0jzjy3fQV3W922noNSYdZlYRYdz9M
hoNx9gkXoy0OPwVPbMo79y/xHBQgdOR9m/QwNgAoU+zxRXpnD/2OjBWDodD2TM8X5Vrz9IDJSn1k
XmLEHi97EQAKkIgOL5lm9n5xMhSYCbjb2NTaZChF1ZgyaDWSbFm4ZHytcEwV2tXNFYaSxNG1Me8j
Fml6NoY7YHXd71rhxelII9G6/O8tjZcS1SaxAjjDOpL3sgM5Cp5RxghaWArThPnYe4aJ2ta6CJzB
QctfUY1BbtNSyc/KJB2h0UgBqr3Pn8TnSmXYHqQWHs9RNEDwJ5LGNMYRR3o7umFdLsmpC4TaE6Ai
iP+Hzw5zVpAMEUgBUmAYwCCq4euQUUhEFJUy7rHP6oqWCmP5iRq8dDgoHNFvI40yfS0B2TOpGfDp
9p2zDoOrchoF+qdIx+txVnR2fjbpYoW67rOr1hUPYjLDxVxL+EzyABZ9aRL1lsfQp27DZVFgjbg2
tHvswQ3Z/b/JU1xnBcRhOkvVBMaJVWAeBrB6maoBFJiAWmZExMaZuoi06EgZGARmMaW4DwaC3QqX
PL0gcAo2IbBsR5YGw/0Ix5u2J0QpVJPKtj/MnwcNUv+6PMqvGgi9URV1oFMtghnGYa8D84T2TV+Z
nSNrSLwf4aRenHxIut9j4ONCBpJ91mkOHvsvUumP1OOWBAI97NXUGWS2biF5aBNmQRHuTVa1T6h9
1FpAPGKwwhuf/irSGZ+qQmgjghTQGL/dStn/rgtexGYxiWcQRt73qCC9SIDRRBthmL0TJVgWAISY
D85QI7qq74nMy9wlQOA2uG/78wqgGmI1OdfwcJQDEGJyHHADdGYjrEIdN1RgvJbyfalr5dex6LV+
fF1ozGW1mYfXASaEWrjTchWW7mWdnqC3BA54NVOn8DLwo2lGD8laLo75bkCSmuHNfDBaaHODwCFl
wMCAVhJzC7jtoo1mlXWpTg6HduQOufjIeDTWvoiS/9xYdHaRWL2/tmZi/4ZB40glvJtt8mz6J4wQ
wc93giAoGxZEvGUQL2wYDI6SI8NaxESMbAtvuC4y1LWpCEBsQ2hpns2ti8DHCeNBBoJYuEc2HFva
nx/nqSXa1SIDB0oCmOqzAM4416jwmcqeBE6xpOsQZXgAEsto22Cszqp9eXiTD2Qv2xljgMlz1pRi
lyEU0bPG+/UXZMaUBDUbvztHArnZfYdWKYk+nVInWcV/k0+UN22N5/McTcOSWmS7J2PMujli7MOI
lqY1MHHdD1Q9gpKsXoNJdTKJhah/pA06E0nXN48tyhFkvCXEer4sDgquTIg+JvM7jf0ZJ9l0nk1x
Mjd1Nq+joAjyr5QgRVhC1kL4jTpF5FTKDCbHzcOGKw0bIg+zy3hF3RcU+dUB2DoamAmv7YfnB6rL
31RdXaabfJ1XV7lnTJ+hlSo6DjonxGGIzHC7PDUpVyzAtovhoQsQ2aU06WCoWXVBghqEsqGQ3SoI
oWbwPdD2tdaQPKZdmdLvR0M8dLyzBDNP+9tOtAO4WX2uPeAh4FAvd8nulaQd93CHaiQKQOljwIpK
IlS7JqM8D3c7hpOFDNN/ieYh1ofr96Pxf3b+bal4Ma2OdPo5FMCeRzQL4vGoMA/T0Off2eKKn/rm
7Y2TNOt4B5Ix4+oVt63j/RhQDzJzzUURwxcqdehZqQDgb5KDeqvnC1kmems4E4CDf6d6Orwtf9TU
CnPOPQFF4OnpmdmCI//1eFDZ9mWvgDJvHjnhyRY1G09hVaCtkBBGyCkfpQn1ALaUQWCNXyORZi3j
ASMwtNh4+lFAJ/Q0og+VssP/4G29kzswmM0odl771IJxJvLJ+UxWz+dT/NmEzVHI954FO5iR6FJz
zap2FPhCBXwBoUNuXViPnsi/PPPQQMURIoZjGShiF48g9p+h1RzAEcBOrz9sSZTGefj63CECGCSU
w4anoP9AQWnxXBn99/a8OSeMxhx50C3KgWl9iPiRYkpCo2S8VQv6Y489z+S0K6yOS2UjP9VJOmTE
BC4+qG5mLKYn/n4tmw3R9kNdmSqEB+0wJs4q4xGd/99wLuBNwq0E2GFt3cndqQt4TH55NecE07qD
KVlDc6ADpyPHbPmBbpYNVLALd+WEtO1PKVzgmL880XjBd2adWDlbfAZY3VfEgKJ/cyvnOEsU8gMe
URotLsrR3arTbed/nOju2sVNrVHWJvnRqg3cVRvzfvfZmQwH8lMwhpNFdBl/61OlI0xFJ0CKDSCr
xyn4KJfqYW1ELxK0AeeWm+XmrOCS5aS/pIJKCi3q1H/yAGzXW06n6PkZNB6puuFu55RNAz1PEQMn
yeyw8Qgnf0FIhTvaIMtxrmiY+LQohP76riMaKAnoAl9tXfmQGp6vrnaxBJo3/EJ5KJ+zaYFSF1ZS
BQLE+1PgWOA4cSMP39kro6BIlc/mtmr3OGs+DF6oPNnkRwbSFCD+hOrQCnM9CwifMMM6rYXpIWsk
r/zBUg2EJRQlTmfQUVIg+Bxic+UT2u7VgXa0zvrw6l54losj1j0aVLZgu1KNh9yAd01B/MDoFUBd
25cvsE8m5O/XTZcpNfP9FGKP3yTGbHtEjY9JAj30W6OlGYsmrFQ5LWEpaaPCK4zoiyEpVI3H7DM5
4AkHIJMBRBbaHqvxwKxwrx0J51keZKalAlOf4PCEfdyF36u/YpJhhQTzue/PjhHQQ3vRVCUhxJKg
a58oZHC+7UIjktW3+Q/ce/oTBGSN9a86qq6FyEViNL0u19TapOcXTUbDMdFa68KbRYwjmDp5HJTL
9AX60HlDI3+3FSEbtEtlEvUDEcdgyNXrs/OlrlnVMoWpqBFyNHE+kv9Q60Mj51k65+ihC04d2QZO
Cw5pDfLR/ZPTUai66YpX+9y2bLX6stjV4bVaLwaQKZJoIb2w8w5sNBZX5Ma6GAB6QSAGHaSKhv6D
Bg9eF9Br9aUxhF5tHzAXNHd0fpna9pJgaG+E9nXZ8xfKOOx3H+aOgRmy0DWS75RVgb+nGUpgso3h
y5Ezo7jMjUEEM8O1P5O45R7MDv+3VVMC8BJSF+kAZpaIPjyswj1R6/M762ml41mx+gfV8wrGIYIa
q2mEr1aPyHGSNPGyv2L4YztlG+KEOfIRsn6chpkvcKJWScP4Lxf+x09UwGrRTifOQjf6hkJtjRbM
8Pa3fTESVWE5iPr164aObqMQRPICVzNxg1bctTCQvWL9lddgfjPL+qIzzE0oqwclu61qH6IG7hTb
wCRgyQ4fu/Mu0fdPOScF8vNOFOCytzwawNe73lxcMr9mJrN+OSocrc74FW+vLpegHmgnNvrRJtS+
X838O0vPl4gNcC2vjk+XRgSR0yLrKlBRPQw4gl7OS0owtL57qKR+w8dGZbtfbyEmirKxxUaYtSkj
auNGho79+aUUrcONKqkJUreeHnn89F20r4Sb1ncidL8LcGuBhSBpRIV1VwGGRofKycu8R+U+VdsU
pWeyqYVE22xJiLwpddJC45Y1eqaZLphoUWOY8pqCJJPzbOrWbre/GBrqtpDvU8zT5ZJhaM9yMwAG
0++/DoRKlSE+qoBPW8NTE9oMmuOw2dqlUrrdhBtgVlMLxLJwBPRMH6G920HQZXhAA/O+5fCl996S
WKC34LgTYte868Nq3F0J+xYTTJL66G2ac10PGpWASRfE/Uyt2f5pNI+eG5acnHSZLdy06JbOzGAT
3tlXQo+6T0GgNSrNGMq+gr9etkDJtUa0TYgdWQqgntO6Y/yx9yvwy0T5tK6A25R0MR/qk1e2sUnN
ddjThQ4tuS3maXbRy4C1aLXgr5CHl9PqSibqys7IEz9xfBFEyUNDgubq1Qyt+u4liSBciLzx1lO+
ZmgeGJFOgrpbHkvdsBOy5dCZ+Dv8y8568S+LmUnM1jW/ZpsVFldHBsrxFNLALO7wrwnmD9/01E0n
EdMG5NkDisg639KeD4mP42HuIS2JiNjLg56HEgeq2dr+x+ZqYW3/JIDNMV1NEZT7olpOK/k3YCu9
/mFUvEXYjOhm9dmOedfO13itLajgwds4yZvDF9l2EyFx+TL6CJOmVipgm6ZUf1SSuZiq41hmUvKw
UerzK2JS+xoNsaBDPdoTOtk/DMFyUVSrWfGSIhk3PtEr/fepArFX5kllpbfz9z24LXhJeqoMfeIX
iCbnTHnd9oibEsgmmknxbekRd1UBKKdpFxfSuW1mwjvLQiHFqsvaypt8SwFzNjDOV5qLyGnR1bx4
ui8ZeeItgfsqmIu1J0SyZpudMboKHJN2KaySzIrpzT3o46pjfixbvSWnTS+D2rvkSZyk/RC2Gj/R
6GuCo9+gXaU1q/HpNLciqk93QCW6O5sD5UnR1F76GvUVZeGqDtBuJYvUChKZw2ToYMlo0MbtCI3t
iAUEM9/fmMgkQuMnx704dSFQjpm44r0nRH5OnS/fOUgyeHbrJlr1tjBdn6j4EMslUhmdahtCgbyW
Vq/mcJfn/j7kpNEWA9YHchtJM+X3C4oRkym77Gt3HX4EcxdEm62iztTSTGf7XMbbSMs2y9op8sdp
8QKXJqM730oENTGV0Lv8SCn7KWq5k2NGXmaYFPnVzZpgCk5anzk0l9Dvtn1hlkmIhJs1AziCxHea
9pyS4JidEEF76M+nzBUbIceAMYGZ0orSqetI21BGCy3Ma4crqiUHKouEdPsFyqVP8n94To9mrGOc
ZU6BruNx/vcO9lzz/OmFUsann5S+5ohjaowkLbunBfI46FdSv1Ur4o3yo+0POgzbPbyHuXVQrxSh
O7aGebrhPCG3kXdT1Mx9wy7ZLhNza7lgrY1+rFW7Tc3rTIpRIG/mvZt6cXlCWtueu/Bq9lZia3BD
lAuO+pnWi+VBQQD5hCbpRJUGNT8dXNJM+w0G56lRVDmwvrxvo84r7glCOxgJIUgTuhh1Bfqhy/WS
zfdjm6TGpvg6QcIsk7cCmiBPkA9+TblZnPPf4lxNXl0Gd/b1/Vj9Kl6CubMHJxNyD4a/7syBHGrn
43VPT7WqBzZVQXbBX2qXzim+mYlJUSyAOhNKL4uuDjaPdmEELgCVKlXQnaoBj4hN1SwfC9vDygpI
bwzb6ksT0UsP4MtmtKykwKymHX9KQi/WE58i0num4RwDHk06silMURsTOAjf7RdKPiL1nTnZD0GG
tgKsK0oJqLWUx386oE60HQ3JQxFqxRvo9IFO+twy6Z4SY3tUsCOiKzLH11WkEUK0Ya/Mcoixo2mG
15gBJfMiEFcDlyujAe26DYAboXmzxoL/wJWmv7QR2n4KpAMZxHntKGvzSaqqxjZMMzzy/tE7T5cm
MyYGTH8zbwAmCJ8o9d7s4mjbLHr3LmC/km3Pj3X/Y8wq9bazs2pkDp66E1RsJsNmXtwBjCEti2PL
sI7Rfss7aW8S2IrEFwUNdF9P6L1H2N+yCDK11QWmNPpkYMxZ9O01CfsfzRKZwMMnF3suE8pOuH7L
cjDAtT+apsVjcQER81TxFvDeJN3/2BYFAi0CNFuKT6wDt8v5yT9fAUZhrFMo5E0Q+8Sp3eXiRFTw
6lNfnljxxK2r2Me7FQ8fEP69/QfoL2db4V1eXfMsQSwwzhI+jsRHJIAmshQ1WoKTt8t4U0GvI5jo
kpL2JzZ+LWup+qD7LFVdX1hePPK8endPpBLX/qI1fN9M+galSDQxStcXWG/4HlFcfL+isf21tjeT
ZGTSO3m2ihSpBS2iIAgVj8acSYA7uBiiTleb57Ux6Kt121fvoi/wUZkNfU/5irg7LjOhnVnXhLCz
RRZn8IxxHp41FwK/2RVF+VTRY7eY6aluuYizdfL4NBYmV2/U6ns/kYVmNxj/6CnhEVufQYaln71u
HuWEl1iELo1902v0c2/jJ/3bWETU6JP9QAy5NHY8yfZgioHqeIlmIXohaXTGtnuhu5nHlU4zbU1p
FcoQ/4O8CuF3hldIIfW4QDM62q8rb08VJ8BYGhxhS677lJ6oqRA8uyu3nn9zWIwSemQA+iyh/Jvg
TavTOv3b+hrrN7gfxKCiuhitsJ2KEh75AnR3w7DisrYib2hD8nFKbJvT0mcntbatuq92deeQKQKi
4ySkKpzltAxjce9kiLBT7deI6CXQ+xi4SgVnvKPgyAWIrc4GgCk48NMO4A8/9OllC/riPGqu0R+c
L+oDzQpjRKsv3X4OciV6aRTRWoYP0CWTJjPogorr6ZcExYE4DpgOo2OmxG1MqsEOT5ybZBa1Cb8u
RcYNrv5ozU70OCyPGkIKFxmGf5WKNTJ/y02Z1+8PsdIc/OluUiqmBq/Kok+ovzrJrQEHhReuqNra
33s6FXy7LpKDp6uy3wf84E0iMK7MSDEJqItbi5dJVLLf779F8VOiP6ygLsTahLIxZGZZFLgJGdHF
FxJoRqLLfrb1wQrzeNErUfqYIdGRoFytE5LH3/nrivLy6Ls/RvNJygSk1kOW7GyyQdKKRpBteTAy
+Eh+ElHQ4KSgCTR8Vg3Hw7NIhGUTSIsKx2AruiicqwVHM/k0IiaGvtkPgBTNE1LqiSTwgpd/PJBt
rCsMKxkdQzx+eXrZ6wjJkFDI6auqDr0T1Md7PzuBx2Bc/iFSAyU7X6T8HiaebxNQavjjuVakAZl9
VCcQF1Fg75iqRtDnEext3CIWoZzsvyIJ3uyr0bQWtppDx7t/LBnXdhScvUFHNteliznJbJ4BcWtX
AY/KR8x47MQ8FMIsbAslzJR1BIR+XoXHY8CUfDkbG597rEGwNISGmCZNVZ8MIqW1vxweDZedvXu7
0v2kesKR/oY5uQIUsBVxRa4tPv7m0cAYX3N9d4Wh4KWRjFmKtSGVfysPChx4y9RhQKUFPOjqhAbm
LVztsEYgc0KkRqOn4ab/m5ONEUsbVZ5MWirHYooeBNNglLdGSpixByUTdupjQnm5V5udUOLntRXK
KqhGVqJkGAwIs884tdlC5VFFQd+IRLBFOKGjKcE+n5xhoB9kqnW1ZKfSPZ3pUpQ9fS9rAR3A1eIj
Cfqp21qGSoXMeqyBNyBn3OpJSP3Yv/Hr0tG01SE4ZUxpLZVgP2tulrsi51fCeSxCBy/M4hiMEbzp
LhInKTWvx8uf9YRHOpmypTBA0soslKN+PE+6VhnCBWumyR5L4EfH8ZmNBNgbayCiqGsA3Z/rOEdp
YBNhRoLenPE0LolO2mYTDyFBiPw10LJuBU/HXtJpvYg/joCBqYBpwp97A01FjHWQb5re9Xu3B52x
kPp40D5f4z2ZFZCIRRVN+2OpUsQAt4g7Bhpf00K7xyGP7mUlcTFHLM/HQfeif0bZC8fdAxXloSZe
s29t9hXntmkMnsxTPz9/j6udxPar0TgXP4QNYzzDNWCvYW746GnC5yGA6fcWvnJ6M0QWCqd8Y3V/
GfW4Kxwv+b5o1ied5/CJiGgCcLidcVShHZSPW4OkBJ9qL8J9i3NayC1/U46N4rLBIpSrVhhVIZwm
SR+qUqYdGtikppUm9K9xFse6RuFjIPYlNz/Vnie3LilPRfmfRWhreyuVvn0/krO16OYIcrX4eJY1
/VrTNh3RolfdtS/VN1bf7W/2siSPCNYhp4YDLrdW6wHPNyBO+DW+mIEb7V5vXn+5e4gzl+sJuMvz
jXWQdL3LDISbK3wHUsVq8WOaipT1oPihX1TKKDDkKtVSAeMB77ksJG8NsCHJZ9Wod5qu6sNaGCf/
78fj5Sb9bww1quOLJQojPdtbtXBjtvtaMc1FHofI7qdqi9+CFzP7nyZHSTqWjWk4Z/D3iIEBWtwO
qenwKs4n/v5EMB2roMmTo7qrYVWFScHa8OimamDOlG3K9uLQo85DNEhg9v7yot41apar/AQ1E7YO
XjLrey157+QIW9UaaZnchiaToe3JLq+5QvE2EBvSmdibYtaMFIRdw0iqbLdrKHoHkLEBMhL92MZG
ML0IqDKdjzfbsfc20MhyBunKC8WB9zOKse2DjrItXWa759dZvo4P86UH2oGOFaTmMREzaKo/+ShZ
3/mPRH+OE71JKSfqwBMx0+jU+Vfe4kX3DbLRwCyv/I/OT5sFRAStDOd/Ial038iHxTpTTV8ZNazp
DZIrIe60M0wy9raPl5eROJb0ncmWqhwkAv/ekTdNKZS3uImaNZZ/XXMfhi0eqgOUSeI0rpvtg+/G
TKzJG1vT5JN696QOko6GxY0FYj+WGsjCwhOb2gKpn7OgRm0HjZkh2i/WfVSpXxkqM4uxxBIuagW8
MciSevNbICS4Rxg0VcGQ3SAteu+LmlMR4DcJwh9rVPbArpVjG2BqvK0OkG3xGeYwtsNedESkpiim
vwOsgyDmPVnMttGekdYI7mWD5NErzqXp/pozJreUP8A/xpZKQLtd7UwsCdbuwpzb1ha2uRw4A4No
923UFb0FSajqOs43II6J0Z9x0+hUwZY/puwQuj0a/EkMgobfdzDEKLY16RKIQ1Mbb6HsAtswufCh
udTf5lOjPHz2xz+0AaFaNffHJH1qzmyNg8JfLKW8R3lwemQ/gUhqPdQ0xnImFFWxR3kSJtSvsyuM
oWC/uA6Xr4rUA1dpygxohx/3OPPuacsfU7RjesCrU3rh4NX1kO+dmkeQp+5zjE0phy77QmcLIxe2
qc+YNfwI+vNmJZwddaX3eyJN4tw/48b+uCpLKH6zD0V0dVFojx+5YKCUBRBFEAOIEbGLiMefaRb5
2IsqUFNGwzhUvMPHnsaM30jFy4vjauO45i6sxa5+/fjGpE7KPke0ouCtminvWvINP1c5176EQ6AL
Uyo7pgtG4H3v1g/UALLfKSeLIWngZljmvqf9USaSG3Ivo4ylhqEgmZQwop/xCYdRvU38t2PPtlLm
MM9mKT0GIsStxS7+NBALpjISYo9ttaH+IehcOAAkRtMLp9NUnvWcUeVQSP5UiDrPZeQwc0eZ4n2V
ePmWm8ong37ISTBmP014WZjqifCrth6OlGOaXN3ZqYVKVOAFMtskg3bNjA746EZ6EyWmqgLzVab7
hiySPGNnhyawbbCHXTxoqboWF07f7DfunRsappGJdpW41O78sP+c+sL+Y5GSucgiYS08UTzW1fNu
JDw06ynCz/TjOMmbX7jXTNS51LqASzorBR7LE29PMJy2OIh933esL6kfREHkvBFLbM+LPyXB6RhH
moctDFg2W4Y8ia+lDpn7/787BGSns6i+UwLfn4Dqyes8ZTOcJn7CAQOnCVjKQoAJmQWuluZvwXGk
uj1mS6ISll1Jl4xZLVJhKZly/Y7ZxkZrDIk6zQ4o4k3+CLIVJHIHkiVG9gKilmYVq7CZcx5wmFuP
RtyKGPKPgFKabf1/sOR1rrlAm9dpKRIrAhlkZGdfxkDAaxiMlyrfV16YoJ1XDpzzsF1NFc2fOPeK
8ADmOaEKTeYq5O6Xr8Ff4gyCnfpbNq71Ujz/ZG6uoJ5eJZVaNJrJ1nF1RI9+47jg2GqoVQ4cjfpA
EVUZvCQvE6Qa0g0SZocrBGiAVT+QSC2hf+2EtEzYlCYDDJfO/tKm62FMmMBmSgViwth9q8AMQqCo
boytAbNRCGRA2VlooQsS/ORHoB2JOEvRh/C3FwHtcFQd+7jZZ7kg7GORX7JvLg6WuEcbjEScsDUx
2XDoFCblADPLmmez/ImzQeQUUek4MIuNg2iVEMR9nyWLWflhx5Boycn3OfbM+Ua3Zm+rMcMd1TXd
AGcP1gmndlkIjgyO1WlHDIbixBxithc2RnsHqOaL8h0wXod6k12ss5BLx5RbeCxn4PlJTpazCjhw
9Tf7EFlwYFer46bQmY3DuNdYMh7mgL5EMqwFMir6Oh2C/DmtZdRvqHSXgvSbTE9DrGjlKNAehZdk
HtSwavMTfPddOskKCnC/VQ5EqY2/wToPlJVMiAB5q/Q6huWGGh9GU8qxjURw+lxUxPXpt9swEcQT
Ka/Wk6AqPybpiQVCdowJELH2vgRc4febVPDHpSRjDcVQbylyqGOFiXjNSseco7h+2/ffh3QBNt3W
2Tgm+Wkew0VawFjkvOXbq3JZyl2apfYRNSpFMoURimj2xHYa7xuZXMnpXh3NZ/4ot4mf2Ek9mPo/
d27Di3gDSeR7IumT8BU9i9tiV1h1hozq1aQQ2F08sEG7iwd3xi79PooK0syERZ7o3boVxsgOmrUy
qykdGTvpXyAJV2VwWkDdu7rJY+rUCPjfulWnVUK1sxGArydsPbEEyLMKVzlsOsPS0sXYtempSeSA
Ksf2ZLiGVu9iFl5AmkZGRFIZaSJP3UdL2gEB3HT09RaJon29Mhid5a5f7IVSyEUBFoi8pQA3TrEf
9eJCC9Zg768sbxuRgX/Hq8pa/WZlwcj7o5eU+ZJweDKB0AsOfy9iMUf1ZKuTM3cOsQSvAhCZeud9
1taV85kCCQwwJuWUWqBSm8oGvHyTUup1qy0XsX7a/16p1VrGtHesKQrcYjhCXaCZsr43YmOroT+i
CNkKiRZVREuyr/omph59HVsByB7iei38HbyqEDz7CX5gBGFW1AY/ZGSFxwI6yjAv8t+twLyNCgtQ
EtIWLsSFe3DbQTsh/Kam6gfRt8iPqKOBb3qkU8LAW/3jeA6lGhm6oBDzGaimzByylAE+HzZiGV6S
vfyoKbXWhBKcMFXjhIYTKjhdKj24QsmoxITfzB7U5iQ3ATzqB/B20f5besb9rMJwjrgL5K67IMPz
pzp6IqW3FjQhG4ahGTLSx7cWSROpquViWDmWTnDtvebYBWjd4enPEbArK3f1dNTKOHVu+xEd5ZE1
756aACyfdOXnKQH7JiOA8YEHePQ0BIT8bi79QCPsX/c9wSPLh0NvQjfZk5QObhotP8o0J+1UbHGS
KRtK474YAXwB80cTSC3Cl2ksTrRfwuG1O1ABWMNHoZ8r/sICa40diV9c5mNLn6MnGY8L892tgfKS
ydoZah1YRrM1UA64a82E0aqldj+1ey7Qun7iBlhHaXy60l2/0y/3UBo9G1sxaQQAhYo8w5a0h/Hj
/pyX7YRY6E7UlyOdv16H6dBGWSOcU2hH5MvDnkW38MbZp30SKmycXfOXOdN8Ss63I9SrMijIelfa
7orVuwz45FDWHXRjk2DJMYagOWsKD+Y8DCATcN9+fNrynyHFXWlrTRc6w33XpQiMV9EZmSB2+cIr
uyyqBZlfzaaImek3glOv0e5YTuHgQ8As/pVMEirO6+OEopuQmHFFfvGWlPw1LX4if4ctN8dZBOdt
MIeuck6L72tXt2BxOMVLrTeRoPoR3QwxuQ7Efo7TQhsRWQZ49Lc9X6L5zwMmaWcK4GW1EGnNFFm4
5xvJtdM3FgL4suHevW9NdksNb/yovEuXUA15XPVdHeWXAgwxU4S+6EBnV7lwBZqV/zHPyyJVRt9Y
I7F0ojGsV34jIB1luX0rdxjTaVOhDWzD14kyAqfnXtXt6mnEBcnbBrtsuYkjc8y6+H4Du62VMLIq
Rv+P85t6wEwGRVXcxfjfhX8onxoDTu9ImypSLs3e7gdafxCFKPDfWbMVQHIqBCZJkmQG51EKa542
Y/G6zfo2cRtdb8sKXGerUE1W/MYYeoQrls5NIwnrx4tDr0gPiEmkfB/XFlkdG4YXFZF56taSAMH4
KlwWlySGAsP6ZM4ZDlc5uon37gKY7Ph84MKJgEdY8gF+/ULM00pGx+JvayulIG0Mry1l3efGzyMp
6eS4p52pjG7qDLngFCK0n+Ei8Kb4mUO3ZpbaSBq2ZG8iYYtJgXTZWafzl0lo4CLKiPH91JWq0Y5P
ExXxDr/gx+ZXixNDG1hzwb//BDWVMfpcQeAhRd5MAr7HmRJepTwcu8ltDTWfuY89yRu5T8eEps1W
Ho+BQ04SnuHL8L96QEw7Mdp5o+ToLzjbGmFYREGcGPs+AkNum5e8xd7qQetgbQy1GuseHtxO3AQC
fEhI1SCZRQiIrRJUTZka8rl1ezBn3yw2tDOOuKOJHaNsyMaRk1r+M8ZPZKa5jeKRLWVH+xYbLl83
OlNMHFl66cVSuHYeUEhT5HUWynmZcRLtxi2Wpaz2Gj2a+0D58H3d8Wq93YjUaAQJtGFLRmIxWgxz
c4GM2q4MDITz0n9PL+hhH8oz77jQl59UGEWrcaaI4MFIntcUyZ0PRz88OQrI/aHqGyF0VeHpXGZR
L6JKS4V7h+VpXL4pxny/1uyZHfCqUqVLZn9Frsy4Xrx2JwDv28eqD4Kh08NMj/bFUHJpjHCxLNud
xmZOyOBLq97eT5WQZc76z9WTmQBYmS1NTvpKkc5b88OvuNSA+gHpvsu+AAWdl79ZOQOlmVOaoXcx
AkF2WnB+FLnVYuEu4E7u+bxQOiUb2RZPXIPI+GJKT4TXdLNOGaOzNzB34cMKydjYjh5OdxzWx446
7/oqc1YvjgIdAUBLaItOtktapJJjmqh2Y8y82bpBKmOWR9AKjd85Rp9U8rKtJauwfso280kdSVEO
R+tpL3NJAwRKTTAapUFS5eP4g5/4Lne5nWQJtsiMyYMvLxp393NfjiurqZd1LjLdx0T8tRUg+a4V
tH8bsQs48UTg24C6S1RqzfXKkGkQle2R86tRp+ofrnfeB9BgOZ4DvodB/cWb3IReVhIQT3y0YAkp
3wBci1zYKmq/pQJfIr3Q3vfwnWLbrWePBxZFx48AoQc5Yl5J8rqAP+KrnhiRoZ7LgPqs0wjIvp0Y
UA6gauTaRCmCHw1BGOZx0mxynTMhXgKuhHtsPm+fu0bQ56EIlj3qExTY/R4O1TzerEHp8IFjEGeN
ie2RenE9olDeqHMWMbkXTLerYr9QS+Unxevow2MZ/6tc40ctmYTmhQ/jq1dKcIoui3V+za4/Ey8k
YcHqET2gkoKTe2hVd6zt07nuXQuA6rKjrXKaVzBxxTDIDJce5RRQK33NznRWZ5Ol/CEpV7s4AzsY
7Im030D+IjYNUiyO6oKkZ2WwVjh2clzChzzfpOIvTvphXZvSlsOX/pSwkVGhEXr81DWCG5xjYduZ
c0CuUO3VJOxuLKF4Ny+GJnTR7vtnT1MSwHlT3YLqMmSEhIRd98RTK7LwV2I/x6B3jgViudqgFpup
n1J6kscmhj5IzprYTSRaOGJd1bhERTLUnGwiYxNPNgFwkBU0wCuHYvU9A4W7zyXtlY/co8eHeJ/+
d+DplOqq/s/T62dE3o16datg6kC9PU67wkBijKYG7mZMdLZCdd2CJ+Oc8Kr2U3nJVGxN++M29sVb
eYMcZHher4CMg9gg20TzF9YoPbhy2IgkNKO0cX1zqgzCLk7zRFDRiIS3z55TRcPELOlIw5PWHuNZ
ndW7tW/HSQva5YW5KdpfB2fV6xokH1pTRsL56c8EPEPXye++V0P8JBYs/zJeAc5jtkBovys/vznC
IPEG4ryQEsCfQnDgB+rCOsFQM1xbhWM0NxanLwiVAZYXvLR1swg3hYVFfRt82fKu6n0DzKtGeevQ
rJRgQKlFNCpqhL6GV572zfbIt2ouj6bYKJUYpes1AwhCielQHFt9Tw155uS4JzsUxvjZVH1c9H9J
PppA9f10oS2ULvnyn1Wxt9AT8edXD5Cjc9MMj/WxYp+8aUe6bCh8VLHOnEcD7Dbigvfq58aYBMl7
jhFUc2LP8k7cqNeE+IpLZ3hcCwQTavimEc981UAaJlnQ2lmCJHnBHVyZQ30XapWGxTjInWDH1eBX
2VkDbOPMhKJ28B3kPl/DpLc/LL7z775nTJnMcEH0pXsPwyLilIiBkWvX7vXa/nCPBU1fDtKkS4ls
LQnJey0SB/HEH9UWaOdUT9hAFcxEZdR+erW1fQ0Y2ujHaiHdluvuEnPkZTYo/kSNDvc675cWW8oD
IdHpJEJrY0KQs+VDwVArwhT6VSkDMDqr/hYwZWXXGX1ArJrm4BkU69x+zwPwh6S6Qi5YU2iuqbQe
N3H3KfnxSDdwtHAtKZ3sV1K9fArYzsgRY5iLuD7nmm8mO2vasi3Nfcv+kc0lqdkz6Dp3pWULFgGT
opGX6UQbKqHoDtVwoTUNAs9PI80BAz5jZqzJ/BJmPMuabEfvsfRDQkPEifctW+pxLq6Or12BFVkF
Lgk0Bm3wKQLphu0jh+Pfdv1xKXrwh0gBQQ33b1gDpm4TqruRDmFFuRjHKpFDsdZo8rApyg/MK45z
1ly2EjEh+tDaoUEt/GEsOANqqG/FuU2VoqdmFLBCSb9T7qcKCevOMjUd+rThKD+k1ntboH5h4Rh7
d7eXwPUwxb8YYBZ3zEvVaanvi7v9kEvEWTYc1tkyAdKOeljc6kZIjVmLdIBlJvuA76QsWVicjiIf
nlDxiUPQrxQFTP8+723SDS1BAOwfviB87XT33RDgQp+8oiM8Ecn/mTf8eLwHcmDD5A0IfOndmGRs
POT1BMWU17fTgN4GJnjvJHBqWgU/24BOhpPkALfv34mMLnvP2VyU1R5gePG41PBLF4C/zUFZw5n6
mfdNKkGTueSwB2m2kUjwsREG3azOtWfFVdObJ4kaP4O3UZoE8V+CrGW7O0SvNON+zYIUwUWVyct1
WMWFN5rHHQbmdbk6wN4wRhaokkm38LZBJjrru9q+tvWWbYhmOHVkwyJp8kNBUUhqFuLpB5Y+/kGv
q6TSxidW0mnEHfxz/8WK39EKZCOzESah4sslxhBC0DbJA3CSBIzgqYjtBnG5AbZ/pF795AKhwbak
f9qPbwgruExx4uQiAYamfQeZqN+ALmabLXtc7chNav0FsxJhmXZH62Ataw7Y5leAHOK+DzNnOFTb
HL4eJOtQXMmMHrWvhSEVJ6q/E0YX/0aNzsDGi3DoKSNi1LoFw/eCJc56MFIHsJI2azc64sEDyas0
2bgNfM52XRHqCC6hZ8WcF4HK75G2BJbcl1wqzHi+FyfiESSMYboylQ44I37ujkfptUXPin7DO7QP
XeEGwfAuUbBBQNWN3u7xoeI7U29uTckMQXyk9KJKCIwnKeHIVQ7Y9qSvHJWN8i2QlMRgRtFkizqL
TLNeYgNMy0YcYGLFDc2t1fRxKFEOCiIvDcIBemQh7FsAHjJ9euffFLkSFtD8pzCGzxzMlsbosCAO
1Jyad7CAuRn9WV2eYzmTRZLIsk5j3DeIS1yx2rxphq1fT3Xt9byksBWyCp+qNLi5ulEhYff8HbZb
NUUvpRG/r3up3rzhx90HJHRj1onCCdZblzr1LV7KYcLUPRR4X6Vk1y3aPK812R7MNiglCAl/93Gt
FSBRWD+HGDS8gURzrZ2zfreyPXEC18BycUE6gx/3C617uqf6N3pdpkZKpQ1KxLv2eIH2hXuuWuym
LHxA0WkNvR1G2p1WIomZP53SLG5LcO8B2Kd0jV5i5PRoY8+l4Xm3GpDqL1A8OHbdXIIW/wEox/yP
tejK7/IRYxRCXHfBBydF/Do4Si6Qlf8sIg++ROHOSd2MoUYx9XXJkN5KDBvuOGlqLz/74MDeWw07
wJltaHL3JsGOrZEeG0/Vxjj9482aYRII0Qt3PXHBGy5yAAB8fPMVWCukDKTz8qLiFcGRfbkX2YwQ
Po4HAyaTPgyn2dPpBV6Rbmgv1iNklNtPfH10Cx+EvuHlUmMRZMDcyIwWiIX+90H+w483tuhTR6kg
TN97mv3IgWxmIjJOzJG8yREcYqu9O6KyTByeAwuLvAJM209L0MYSJTSh83/hlEPe+1iGX3L7KoWi
zkAq+ZpF4bHuii+2NP+3ACDVXdo64fk1D0SObnHeZE0wxU/+GmkPMpJ58pRIXJ/T2s5SgWV7dnVn
wW8PhukMYLjrAbB3X61YzNvdDstp3Z/zGTtZhtHqRgJH5AaH+e6q6JMGpQ10kSdjHNltUptqaJNw
c89lKWqGxKLqUde+Q859J7ZnaKt4ytMKM5n1AkybBUDiIKvBycsFkhuFjq9N0RTQUyVQZgEL3uOe
Gi8NibRYMAw2VqZzfSE4tVnuTpG4OhahobQN5CIFItWrDhgnJIDaoansVYvGjKq+eabYDIRo3QGP
pyYkX77VjBz+ud+/HYzmGL2ZtoUyILHlppdEiIQCbwjbCxq58OJjMwptD83MWHEbThYYk5k/pOWN
FSjLQbB6Wds4kRIhaEcxpgSc2Hh9xe5Q9SCjEREzIAwcrirrxRPRaq2wBOna4LFj5pVaLLznzbVu
mMOr05UOOGBfrjbpALSY8dwphurHUDAmM8JDDFFwzc+6tKpJUBOmkREVNfrm3CBMD0Ag3itK7som
ERBhYo0EpWED3ibOGQnuL0ti1fX/f+d1JiLlte0gBIgnTvr/0cGCBt2QWBFp8Jc8LPoi0lIXnw6/
MSJY7AvvIcUfwIFoRB5tZ3oCFVaF2GCqk/N8o/JK2Zb5ouAomaPpnN90oFuNcvNQLiVyasaolU8d
T+zqZlyyZ98+W6udtPMDVKtyHTQ/H4vlNIT2w1Rf45wipIIlWNhZg+vVN3UvmA3IMBYuDCrjS5DX
SqW4C9DCesJQ1RHd7YhcdgHgr35zW9P45eZtHQvhD1nORWSQuQYEfLrC+Cm2tD4vXnpOatZWSJMC
dzf1RVygxLrS9oWAJI6eNGETqNFnSO0r9HGvkb1eTysugKr6HnaR2kxdezYmbqeUWvYu8GMNoZ6u
oTemvUC/ja7N4WPBIOyd49wl6Mb7e3Dpct8wW5dpPmQX66ETgEybeKT6hADCALDh16veu+r5rATP
CT4a0zg25E2ZxUyPign4gc2Jdvg0APm9wSVcFLiFdkTZJNn4SN2xY7iF9YL/yas2lthhTegr5ud4
ythQpxWgpIqVb6oOrSqDXDmozLBB9eeROZMQgpn8QBaMlbBjNHmQgEapVcIPq9imewDjFjF/OBUH
49JwfpjFrNWhhWJXD9U5PdRgW1IsSotiHoisRezbiYwULIPfWpEdW8c+zMcsMaIw0zzACRY3F6Gc
TpN/mpGGtOXxTjWTNbFIhefNrE3fzsvhTB4kKVi+YQNgAX48J9RtMlG/SkxRIIvGjxdgcVVQQpwT
y9bOwwtOMxjrQAw+WSKihuMDVljGf77nh7zX7hyjIxh/V1MBv3NEX7fgxjt4FVYojWTARDvyBCqo
UL7ZVsrNKdYkxfbW03lBe2GYSRzqGHgWMV570kim+gN7oVjSWOiVb9BnbwKkhLkeul1ZHvm4tV3G
JhYQe69+NoCqQS+Y53w8JwmuQXd/HZMPOsCzkfAa20VPM9ezY3KzHws4P9M+eAPuSJBYA6qAIqW1
eWOXEbGeBRqwCgQcVKCLFjSkkEXy3AljnVN71gJLIRw8Ib7JXsUN8EIs+enewqPK3RhmbX/dUnwc
WeAR1cvTKTy1qgJJupAfPnQgPqUMtA9ByI+NWjKQtWk/I4u98gxJlOQ1ufo8ZZgvSDC85I7jgZIZ
4Q+aTMWYj8fmzz1KKLU7X/zB54hZKuTHhhwQDqxAeXzmLzhHlQPMej+18dAOb6LoMgr3IScp0BUd
42eT4XFACXHlsVS7knjRCI4qD6++pyTWhG/4LxudLgzFKrhiP2xiLU/ytJWIsN0wYJYZPAGy2i6I
AbCNf6SEsPhWRjkX1aWUcoWaGo0cXMje0Vv7+G6IExY6Id5nlQzLdFxwE5Si+gltABZ4ylDvOw8p
xRkJ8+eeyVAGy0rZJBapcc85s45WMT0SbjZfllMwlQ572RYLOOF5kNzeDvpZR7GpbDKUMNSsl4rX
cz3XIvcE/CYXSvIjnww+ZJz1cht7udFfppnXC32WbBh103XnNPqsGuC6PnkwpEEs2s174I6zqnmM
G4FkTmODghsuOyYU7YUV2JBfWTcdh66Se5zdprnQg9PQtHc2m2Mv/fWlvCGn9olPXkmSLZR/fqtN
YllpQs8yHQaMgtB+yX1tL8WvFqy1kHhctHXMvPTV8Vs+IG3RW64Af1KeWYXoxvFGzJpfukk5RY1e
en0eqAVs+02qQTqaSPlr6D2Qghe8iDbNfX2gFNWHEI+LIZMDUVsoEa7wDJRS6HdBEGHbdHdcWfty
jdYXu9iNtgg8jWHgJLnp1pi93EBj016x3oT6B+PcYUJiZ0CnCkve36a/c5i9qVdzNE2dt57Q6Khn
bo38bfEYRKMVpiocNnFglZZbrucYDPClu9scSudC+d32AGg/ahL8J3laHWUn+irdnrir8VR4tTL2
eXlVhZnpoKc5N5pNEL96B5QhZdbMEAo46wwJU7eOKMOHZZZvYr4IUK+aJVMf0EL6eJlGEbAU12k3
aM7QbBw4Rs9MIkWvVdCVSEX6zg2f0Wn5dVUzNEGfQhqDxUi+WMaYTtDrOjJuQ0xmf2L8t8kwKXwM
N6tYatAnq3WjGnqo+oKiPmk7rMigJWVwxTm63eoSwzi1NwKQiFnFz62rX6kDF0mLkscpuY1m6R7o
QYsBPpxWUQPOddwbiKZEjJ2OcLWtb1lzOjIpJEPridoVGTHOvhmS6jRpQWNlXuVDY0+X3JAG0QqI
iS8wTUdAsAyqtKKw8IsHWa9eYRmx+nNwJ1skotGJagHPLu+gSdzZrFNSvbANcfsOGTywP7+2kRG9
Em/C0oTPVjMVzybTs6fsB/VPd0tAdV8qVYBuKoUSG5DxGQPLaVhLUFW8fKNlr0WWPkOYVu0eDMAL
pQvvxZutoJwsaa9YIhPMPfRT1q2iIB3x4XtxpXSfcvDJHWte1mBEn6FCa2kC4AD+t8Z/5D9ZedWI
wjAlROp6HyUVIBJ75FQ5q2hraPFC8wkoDuzih2ncWSkgk0ERyfd1lkJyrTPczaJ9MqA5+sZF7RaJ
DMRlGzxelzsv365mRiuFMiAnIfvKRvtwjUMq2otQqoen4PX8iokyioPlys+jvWDsOEGagJfURJE0
2VNjJeGlsgPEN2XIPN8In8WiKs76r8VacsT9YQyQAKVQLNLjgdrunmRhIL8bOxeDRlx4H3OLV9f7
wgsp4S4NCDaqHeFAkU9kcpyF5bh3lcx+x7wpfz22EOFv4XVCtSrhazlahN40rX4WjqVMlDh/Tip9
Kbg0NhUwfIzJODKnq+vd3oTBgbreqX06dqu3NrFmx7/8T3rAdfscxFwrafDfcScJHctHyUR9+2Gx
tXrr5tLMXHjUh6vVH7GoROe31gZKm+ijtA9L4uaEd1ALPyFDX0F7lmleT7yQgyTeBhlx7nhvndm9
viQ+6ZVdtX6VsPO16q8eCXE5xRSSGf2lTxasRZI2ePk57F6tGLjemzsXhE6eeyzbZHlb8lsaHfIg
OVPUx6vNn2YIuNbd154XTbfjAuq/mW7qry44mPnBENRC7Tv1JK6hLzxMJg64AyKMhZMi71szmtVA
D5EHLTAmJ9e/r9jV2IrTg0lhFLf01qKf//+5kVqFf+K4BKA0LUhAebtBR3KR9Csqq5CqHdxI4y8M
fiBWVSrnb8jXmhYuX/YX3+BL8DV1N01Z/zFsZTJ+cTsnFKLYNsqGuHJXi6ri+5KOxDoNJXqQeMWQ
0H1xXEE3C0xH6o9K+s6YbRivi7qgMJ7FDS5QEuili+EI2+tHDhV8ucZ4J/bBfPiOxzA/+ukFFjEg
dFmxxcUkHHqkmzdBPRBiJQ1te8MZoVAjViyHDvuk7OnjAbqZJaamw+nTvyGwoRySK2VumIDQTxbM
ThV650t0QnDlGo0cQAuhVdNlJ4R5McdiqKOFq7ae28tCNsj7dVseOP4JOpdhNAdg45w0NvM3uHd2
2Ako4VylBrVIsiHcWIfT9WMrb1TS9aE0YwGKk4umTcMCRm/cBQi2VHfSXN0eApG5fT81vTkhYsLW
rRP2BoC+C1qoGdZQHF9dzEhw/Xu3eqoTdZOBXPrUy3yg10I5qdkm3cmOgZUFvrDKQLLJ8dGzqLSA
IbPIby7nDS19Yh83zOYdgnPAgJx5CkY0AzoASHQHC/UFZbDtiR3vYSzge+UpGFDqOsFO5y5p+kVD
x5QtCSCKfTK+nnAgoZZKbookk/OdzYm9LRbfsqmHwjIGAImuYVfxmtRZ8bYL514GQn1STSZIgISy
LMBeSnOciHCtMxmEDvtReMV9kXjoMiC1pIsqwMCuTsUVNQqH4BR3ImC9BT4dAZ08TNYZyZ3oYm+f
nWCK7JzyrNCWl2LARudIVjA+hnxCsFG11zB2cHnKRMnkRq5RY+TbcDNIXgHzlkY6jrBBPtXWgOr+
h+f8zO0T1P/55JgjCYp45y5CpP+zMg31tt3fijRLbpnshEJJmXcKDxlohTKEdet0Ow8lgQ/C5o8x
NLoHgOdNHIZJQGClKjtdIu3lAqopgc17u35w8qzsLZbLhmPB+ZGo2MIrAmKtaNw0k9E+Mv7zgpTR
r7BHs50wVYekYsWy6mWMIDxTxU1oj4DuTXnc8Bp4mjbB1hPXmXDlpNQNoReJo98SdK9BpMEFf01r
Xi6m5El8v2brODnkGwgqQ/DC+7kbVCz4wN0pl7Nzk54EE5wVzhpZYl2f/PsCNGuO+aq6Wrkj/NUv
mMXdG0LooJ036+PhH8mCF26bK9d6mUSvouF6Se3kW/+0W2uOGUj3u5RQKpWlRZdKrBSMQcO0sY0Y
nc5A1Fj0wrYb8bCIeyAdQKXtAeB5c95Cxsiju/tSQQgaA9awVuR6qMI6VTL1Z3ja2yAt5FanSSVT
RuUbxwmCEG1ExHleQj96276Gt6E7tHtppJM+ICMZkkTUCase8Ff7DcWNL/Pf9z40Sza4ORKdoAbL
c7oX/JJYXXHnwlbWXXkI3POiqQloCqroHc4K4ODcOnZnJ9jvBlq2u+EZzbSWUfvC//X4DoVC23Ae
1uu5+fUdndVNwW5ciQAA20BMpFBGcVer34tqGagNonJPgZR4zziUJAQqjtquwZU5XCQEFfPWM5uS
fqtqQ0+gsiow5ZR4ycp91E+Jg+ZHX/OeHPcsCr5gpA4X6OXb8Ffhi4N+J11NE9Sw/uaLZf4Gnk0j
NEy9vHJOW1Oijx2kUDXlaXS9tuCHEdX2H2uKFra0AAmY2ZHxFXCOWUvFI8byr6we5YDBp7hvhIpU
GyK7GB1eNNdiQQBcwgthHJpadbxQ5jAodE7n5ZMVUTbN7b1k+tvVgLIIY9AteXiMEkr0VKhouEEo
DDVoGQLC3uuty+bGPXvX9ewnzGIgUV0WK82io3OloDZ26QXU5LwTrFmX/f3Jd42ja7R+ii5msTBh
q9MmrB/xDdSWonwpzjIBtRiy/Wu58fWmV3RYD1ycEhnva1WI9ww53SCH+FRbz1JjerH5USraUHEx
hjwnK1/54ZDURl/ghbh1jm4rO9uEK3eyn71eyOm+2ISPnbf0gyhpwhvVDQ3vsmS25OkrjyNbr3pG
dkJjROnJ0kQVY1Y+rcPIAs/845eJtJQFpoZAL+cB0uFSkP0sEpaPqp/W/8TCxOtuSnU7sxRv7gyL
Dgf02FyVQ3H8foIWZHNVoO37BqbEwrZ2hskcNn5sKnmSkaCx3+u0p/gUZbQaYH1epP8ac9AlAAfj
2Q8z88dO+q0w7drw+zBwUYNOwMspPEEcMo4SzLJb/ovvXCpv1l7w0hlsyq9FXE1bX1+YTCIxOKgr
5cRa0T0zzzHWIq8NYgY996F5FKQqZak44wIl5lULnj6ZklKla5ssZjRonMA0tvuBEr/3K2pxI15W
nEpx/ta5oiv6ClegTVv1oeh5n4UbhhwGb1m6N8oeQiB7Q2QGJr4WWDud2pSZpczjZI0uRAzz/niS
nXRT3FfAt8hW8L0b5wOyRBepOsJViip8vRZoFliudL78qC3R3VMMjBOOvRXn4DWbENzsHJnSZVzk
VUmRZMNeCIBvPVZ6RIytLkcEZJuwKx1VgOsL/Nz4myILQAHlc0lP5UlkpETX12NEUnmBwuQpQzhS
THuErjDeSsJo8Ja6nl/BWcJmajUBLW+DxsFxe/eFbvXdmSqftF2zcEEw/AszGOQpDSFRx0rSaF8K
mLZvBUwme78Ajegm4Ui27/WwoCWcUo4OwQ/SO69dJqjnQss9aL4yPzSNgb4N5aRC3M77J2+oYiza
Xm6FfkYd+Iu+va9V5KgXHNVPohj9DM3tAdndQcQyE6Aj7CxOlWuItDODRiMeFFOv6nrNHQonPn6v
0djeGALDB46JDOkbQRVHdtnbCc39aAWqQChle1S6uPVN1pS2NgeACLIolM81c9vUKGeMrCliJZQZ
uL/SVWqK0Bh2MWsa55C7GWO99ZxsF3z3JLxUnKxjSg265VPM3Nb+uoh3/Ea4EoUk6vA8RmxiHXfZ
a3QGPN7aA2N77SYtvQfOuYeiE8UewNOcihPq0Wp/e00HoFNslikRsxwY0dfCJ98pEb4GN3W4ae59
4LdbLRyyG8aEBSL2IFVMl7eCkTQ++R1tGlBtlQU8sBAAFzdqPL0X8SuzFJzTV4ttBDLlUkqEhLH1
v3HM5vU0L5/u0KI3aFORPjQCf67Dl4RNJRb+qz0ox/lonm7yCTMJw+wPMv06nAFHnpA4t0UgKoUJ
9qN2Iz8LBQ7vEn40gahankbw5OSmgzfilb6+fJWDFtl4tQ2TheR05rKaMcLGtHuNy8UGjA8jOMFA
ts3nqH5wZLWjHZVDkZFf0N2m4DaPrwEuGW+wYVKsl6aSjcPiNpYaG7JM4/D8VsTVxH6kX5fr8hf5
/mCftAJcd0JxcSVo7LWGrhHpawf/a57mIHIiGFfvRjcdChipkDkfw6FfFqUV+GkC3E5e9Vh/f0qD
WBAGInVEi6+iUSVKstOXkJ52wjGMa8bzUCBESDkFrNLpFHrPvnarnbWkFeLfVpef9IY9fHZRlkGX
Muf/5kSMAX+GYssg+7IKsKJ9vxksfyUlkW3A3q3ruXabXLRBBotPA8hFIL2up5ikC8nfeImOKht/
x6K3rJ6JK+Y7bSvV9b0+AuSVFsvAG/ehlzRiY7j+u0E2X8Z6wLsuhHag9EcxZI4XInyNqWXBoq/T
8MhLUStwwRxZmfqREmqgAAASE4i6cSKxVkQKq1ZqybfHMxT1FWcTCBEfBQSjIje8MYdKUI/amIz0
z80Pm7P2EpGdA2SisrNXWTiBZ0Rhz0rc/7KhOrw/SLl3ncNeyJAdyr7MKnFbE41r/RjdDjNH2I1s
++HVyOK02XvmliaK4nejUwYVVXzIZ3E+VVSJ+V0gk/C3r8lQURJK1SrbYfvm5DVN2CZ4MB2OPZYh
QkPEjhAbeEMfaH/56DKVOEi6p3tyQud9eJUdQ+kA7mXiIcT6RodicnhmbgToT7N5VUmiJAtUv3Pu
Rd3N+Rjv3aMN32v6z+sPTZM+dc54wngLmBEQ4A1n8UY9AZGNQn6AOBc8vewb/KvHxR8n5YXeK5r/
7WY2xdI7XY5jxzMMuPp+lcEPX3mfQUkCHqW63ovmiAYKcoZNmUDQlnERkjwSEcto7xh55dJjOgpS
Of7iroRwCfAmH3GIkV4YT2a7YjMBKGz4P5WZCqKY05cIxs+/+FlAmsSHYH6dYFtHuNNQmnm7FNY3
W7LXFhGFg+YiOf7OsMSL7IeP/Gs8WqccDYFCJ9SiWdEoTUa1mb8MvXyokxvNSCrJ+nNdwn9c20BG
JvnXLKvA5jlAIWfya8kbCa1+KahDrHe2or7I9DdZhvPCMW4BQmIHAysG91AUtvdpJVywT3/hC3FR
sPXICLRYXuZRqjRxgnK77ntrSBpzLDloTJrKVY3UGWFtGKIaBLmr/7oh6VxoEQbRiRoNTWO9bCE+
D0lx4RuI0z5UHV/Xki9yb1ssDuhJa7So+fEukPNY/bmIRVq/5r5usrmvOOUziqD/LMMlkugCx1jo
n5dsT14j2Ji3E0XCQT5iy898ufROI2XtmWFkFzmd8hDavcv5b6js7yVr0IDzCOrHgU3Vs+8ZP8Yp
7JvBaiMd0wMmsX517Slee4kwIWBR41a/n5u9hB+DdWqb675Hzeu2XLHxitRG85Z2wSKQAxf+7SEq
Qzwmm5ubuUbyAiokyIG/wDDzRvrG5UdtR4CeHd5uQ+kU2Acm6K8g1Txp3tEboyX8GPLoCDhZxb0E
4EQw+CJOGMDXCFf3q4/Yf0m9BePs2l0tqE4it2WnXuNcbBTYLvTx3ffR02NGLhOr/Yab90g+RRS8
doPIyQAEZ/9ZGCQKs4dpe3PxGsoXXSMoB6I+Vp1/4Rj3Aj/CIXVLh1pVFpW2cxFz+EJuluMkCGlb
z1gL0ZvzIbUSzW2+brDjIAMQObgHXG2UYsoKHE7qFhi1myL+Iwxyv1CzLHxz0zqqapPqhLjYXPdX
+vJmySNQ4ppZvlbrCFonNvWdWyJNqfixlw5pcH19/6IcdixqoEU71YUKEzrZBLh1sNi3jtesLvUS
WX8B2MG0erxoEi9ppM5K49tIsFTlDedt4e9l1DhsCGM6A1D/VZrWdWJwGxP8ibNcNHmMobP4xol3
IFkJNg7cezMnNDioddbOfGCWHSUch27j/GKUTnUkI7d0oCQeV/rD3Etr3JuTDUbfrptDXAo4+3WD
UkP/m1wu7WTkpqh+CzkbZAYQoES0V4MfIEiiPXQ6F76SO1zzZx7acOWGrayEa9k0eho7xYgueE6l
YvK2ReGFNGQP/+lBHy1BvEQS6GvI4OnAJGBNZ8Jx1OCE5nJBSKWvn/3J5S3IPHYCQunMILzZpIAt
Dp9oq2wcwy/ppTgCWXHxd71plfSfgPO1shTpK6U7jW2kX3Jmp+2I3LzC2gzxwj0C/aqBXr2Bun3n
WGcGyQGcymmsKxjZrPGG3Sd9vkKNgGRUB3ybEpvB8ej980H4Xt7IslPyBFcOdN+Tn9LMdNgB+KlS
7ZKO+vyhqO8CnVIweSqqwYVAZvJTh4pUYsXTBDoyXACeO2kR46Bi0FVgr1iERhsyhY8jGhJDWEK0
Vd6Rtj3/LkHzoXpLkG5rkjUiqd9oOonI/hye/nBdKqYTlfORxW4K5cmkG2vpiB1fGYEhGsBVUuOo
VenW87rjVV4j7eV3SCKeDcgfatRHIqfONchmMTLycfLsyeZTwp6DgKwACmAfrpfJtG+raq0UT6q3
Bk2jG0GIWzhgycUzLcdUbymHQ0Pt+uW4uVZV50PK4Jvr6WdWsGGfsKavZ3yoOO3tg87syqRD7GZt
IANOI23iiZN06KFcKDgfCDdgBVAYeguD+9rHYIXDh0U3P0iC6qPE/ovTIfAmPDKTBG25JAeyDtos
w696mup/KkmzSOwkNWIWuOKA7K6O1nrNs7CtJklmCI7AQY2IimlFVDXHBhDDrcWmFzcNhgTsTZLD
cZg6Mb3CSVHp+hqKN86CfpjG4iAEhIn6eENK8Xj0rFCE5mtovRxXN63KmAUoUFt8KZa3oOH4q1Tj
87KTGB3TAK3j2nXKOo/pu8BCfauuaymgxoUBUxms2rcbR8pA19mlMSnotnlLvV9ElKP8O/N4d/5x
JzMFnqcPDvB7TnRax9p4GMOWS/OHYd0+wljFLYwPXK+lnrUaYf1MAwarPMY3fQVG577yCfxIlg1T
ZDvL7yWFRMQpUmqYP27ZTmyy8fq3CrmbqfJ7WuMPjJpg51YpkkboXjNBbL1/ce4xapMecfb6eo+2
n7uAaYKhAZSCbf+EoANYK03WTtI+wIPsdCfs6kcKp5IcmRUWcuruF/QzST0q2Kw6rA9xRbWSMoKa
XFw7gfYxkeRAuFp20pZLGCGf673i9neql8Rp9HaSB68bJDUExCFc4dd4YnMjGzvEW9hVMVwBs5bP
B591ELgRCoTEHP1ONt0E7Sh94acXVhyw4cpCN/7M1VSLDTzaHPVAKE2N4vJUfqldX+8j3KwUHYEu
et0sXHj4QkuAZu2yxqQMwp51YbNrDqgUZ5FfkmdxkMqXgB/pL38CMhqUTjQx9cAy3mF/Eq0RXv63
S8wcm1nvUh0BXYJ3AZlXJ8jnvHFA1A441PXP3g6Zematd7x4jYnveDxXcyzyV+pj/mKaoefJjK0U
xnGCKqvlWPfscWFGqFlYF1QBjYDFHM9lH9FOFEc07NKwXTlhbxFf8LwR/Kl1aD/jZnS/Hb4PxzQn
O50/5tovIcwgqG676i9uwqHvYyzzn0sv0qGFqweYfW13H/FNRdqYXRAbax05JdgN9xwN7yGXVZSq
P1bbwa0Ug1FJW/bsZ9ymPuip+d0vjjImVBhzlACqLahj+/2AMIUt/haH+c/e2yqGRYNQn7ghxj2D
ArpqJi65dqFgZapxuj/mCCs1tqtuL/+ph1LSmlK4h15YiieRTnie173vFhw6D+Ai/QDcwvNJgZOt
aY/Fnu9Kuc2C00XUa1oQ/eufa1nArwpv1FPECgBghPptcVjsAEuRPiricTnGM2W4KFCwCQkiZKEi
WaGYGhi36unJv7Ya8mkp+Aiz2sa8hzMOjI+Sol2UnBA4aTA7WBOg4EmHeu46AxLCw1mGFPk+Y8/I
kc/TzemsBTusIZQ7vZ4q4BuqNxl9oqSsHXiWfvaCuJee0LrOmzzKlLlS4YKv6GXlKq8avr6VvlIE
nfix1Lom8ixooch4fvt/uqXNQAg/TZpfeZf1UwG3v1toTRvtC4rqP9Jwv4cg6uUOS5OxRUr3sc53
Tfvi0gHdTGvJCwF4ApwXh1a8ElKNtliQyx+nrhmp7eNsenoFvAlDgVSykjD/lJ6qtbB5Y028qVum
RlOs7llXBurGd8ZJ9f87Ja1T1/aL0iZGagVuZqK3ScWKJpBb2qevlz2vGTvvEgmz7VFw5cD1h1S7
mKppiqnEeoYenFhYdhNiPHPuD2bmLTyIDZqELagvxBkgB8q/9iIZuUuTdYjcvGW82qjizXs63gbM
4MZSs530S6tgjSeqlm9m52ReWsThjz/97wzZyTeQYd2tbjHHaRx8yOMWjgYue27eq6BatT4R7m9y
ocPySBnmf3H2ODfYrDFm9ctpXjGwUQYh9tM/nwV5Jg7AqEm78Ahmohihy4/yLGbCqS0DjCqPt/5g
mB9ZVDu1Rf5Yn3KxtqQq5ACGJxLfOjiIIuvBpHta5VnlXP7wcxc5sV5VZUM2Ehn6ZwbFvUPLXUsf
dfRQMe1HLOLDhKODyL/aanzLxLhNcf4xuIP3QZD6Vqz32BDoddA4MDoPaLOXW49qsuzAWqfqqe2p
k7eSnH1uHXrFg2hMcyJrpFTt+eU4vgfjPGelbQ3vd7ZHNsj2N0ht8pvt+AphU7CxgEHQDMwvJkdX
X0P124Xo4i35HAsU19PCxyOdeqseK5SEPF7TINckotKWAZlWjEXeOgO5E+Ec8iRwaTF+4voEL8rT
yzBQsBWZEavuovxmlzkCt6STUGZLeWWaVL437rVh6jlBi1kWk7mIerUI2cTRSSwOusU1A7IN3Dfn
/md0dCZqtpTJghH3u70uIG39d5B3i/n4Jm/BMwNb/PpoPOZuweYITT3K0sifFZJkZpngwpGadjT7
vo92fvBRgZnqMA7XppW3HU1N439MBsHJYlQ1qJp1eIrrXNaPsHGvHdgJTh8zZCqdgyM3kZc9el1D
vIHgZk9xinUqAK0OVAKACXw9G9n8SNc81rKUJeLMSBZmSvrtMMsMiFtwwoUXJ/NP9GD3gxb2B8Lk
N18vmfbBGTiedOdRxu48+cJH7v8fIKG5W5Vo/oK9Jw/MDoYhy4pvNfw0gZ1UKFyDlaMcI/DiECNp
1TXCqpFSjcoxjLpxh0aNnxFVo4mzYYqQjCOcp0wOEkw/YUjy4QOLtSypGiDpqS1fqRpPOspYWyad
9TFW10kHsjkHZd0cpW+WHZicLLrcshZBfe3T7BEwG/eEzx/d6qyj0giFdWmiF8tDS+emjLKjSxtN
P0LMxIIk2TfZVGOmusMmn8PAm6jJKYClqOu1MqP5/muPYEaiW5nf9+7IpCcUD6a9zcOr8Bp5Scj5
mAYKW/IxTwmb63mOuRZsbzl7XaBzsq5AO2ziNce7kHZOZAMUaA7O6qgC6xQwnTZTpHYR2MB/u1wU
6UduqK3CchtDKhoQoOQu+u6g8726FAgGiqrb6C5pPcICWWc5Xcthlm47K6dAmNEni0+yQT713XsR
SStifGe5TevtdW20rzsQMZV5Y1eGI7QMSJFTJC8/HAGbnjU4el/Vh3Swbg1VbSqumMsvAwNwf98b
tgze3Pex/eV/9Nh33f5qzIFym/9hMqA11WLwbPvXIU7vZjFNm9ICBK2UtZNkxhwXTpomyeiSm8Xa
qFFpNRuWhhRpXIBZs35FRR0WCCLgsAlJ7wJvzI1PCN/EMmUc3QhcDaEYyeB2w5Ly4FDtCtQi6hTY
Y6aDKvqo5AaFipebxYym0RA7IxEKT4+CDT4kmVre+ongIwsB7QB0BC8laDGptpD6A3hQERTfgTZ4
1+KLNcsejAmZDR94l3Q/89lE5E9UwsavewTISE5OrBLgVIs55uylw77uFxcvQVJnYjGjI7W/S6wi
Ya+OJRiUtuMEE9NNFlr1ljNmv07aHanOxDwcGBBF6Qf6Ro+aYSTnQZzPQobyOKrqpwLNh5qnrWAB
qNrBasMzxx1/ynhGAgsBykGsxdui8ZfLeZTkXahvFuuMzOrFns1QBmu2fHF758stO5xRzpVGCKLu
mjYe2cfyYiumYvLNtCXvHu3q67UWS40r/rxuofJfMBQYHJRxhVZVbtd25YlEEgUI92w0/PBRVTCj
2ekmMCW3jB4U2CmimxSJPHUsX2q8TEsesGz49GGrV6nxjkUA0rqjEXqxLgJFso2p3FuTfCp15C2G
+tXWvoMKXPyLfeC5YBJyFzK6kmQ7XebVd8Li2Bt9klJ6r0buAztXgLKq8fVKimVZApSh4ZPqQ/Ue
jA+PlK9RL+nXzP0+NOZpSsE0THAfesnyCY94NJXfxNvFo7wlvJQhAFbLxIFK3Vx+NLrhk+n0EkGW
nKjyBourcHp+rVWZOh/GXqVLBepm8ERmLp6KobfBh0SrH+sO0OTGW13hW7NyXaMYRy1j5himr1kk
2OtAaJtMadXb02cZ2a9KkIbM+WBTt4p+8yJ33q4FFx0dP0UloPCQw2QDaPC3xHDPxt+L7dprc5jB
7v5LTPA3YqvJmCEkFv0GhGP1vWZzEy4Uutb8B+ZtfIsFPIKTZTFJlhciXU8CgM7VsFlmczMO8pY/
B+YXOMS6WjxM+VHhnByzMcPf/hCA5084/0yPd42SMR0QMIdHTbjSagWYcg7uFIbIl+ya44FXilzD
p7mNbigPVLONk2G1+V0X6PFya8x76a4zfrHQkFT6Vg1Y8RFxd8eovWAi5v8Mt24WlUA6DDd4NLSP
o0MPnEed/93uVWrRMc2tZETO8fQ8rgfZKeBUSXjBRB16gMyfOU1tUcRq5+b57l9ucWauzOVZ5O34
a0RfcktrN9WLnNOIow90A/Ds8SNbEetCga3rC2qu++Nf98MiPcGdjtFrDpycQ96rzmIZk+X21rFk
uvVqnatd6aGsFwxrLt5+0RaV0noNlf4ZapXdEmoQtuFIqYEInYAopx3Cm56fcy+7HlT4Qwno9f+i
hb3fnbqMhGp/UXmH8tZ0q10SBGUJCMV/yM/1YwSs+rzYFIugYP5y6lDDZv6E7K8ADML10MIs6L10
GGG36USuwJJf1cVORbXCle9msbEodusKGSWsUXby8B83FgxiXwi4iCfXOxs+xcGIaVYeSlrSu6Qy
V1eSEobHcisDAkD9ARPJ+9Em684vc/B62OE++/t59xc160Z2aZbxdJlqA6jNfWjoybqdBmYv2oK+
xtXAzgZWxcm9Zd3Fqev2gBh3wW/vwtRqkC6zGohptetISTWcBhXW9jBwKQLiYNpli94fPxAPRUeU
ptILo9vpvWMBV18H2yJBYsguU9iBwi+TM6UABkDun22TSHWWjRAC6JyKcb5ptYS4eh9k7SDJ8F16
F/lkKcMvzgplcGMg/xuY+8b5HLVhHJiHGUDCaqgcnkKVzx6alDhaOnGtk4w1YkdTK+cbP/tyrrWG
f6R8Fo+xM6pD+5xKoqkdQNd5IKvUupF4R+4HmvMwy+F3xHb9Wd664Sbrk5WSkv0h4fg7QBtpoulz
c/CynoOdb4Uo1BZmd4ut4j6LQ5V9qCfWSUPKVv612epGFGvsuNdJTMfL24dt8aLmCBXb1+7A2ONM
P9NxG0VK9a4RfYOo0P9ZQLKnYw168iQNf7l/vSZJ7ZXxcM1cz6j0zOXbmBhfRc5FSj0YwwOIpDMS
EPq6yafGq0ESL1GYbS1XqF22WQofzYQFm75IJvVXhz+LHo6NbVdF5zrY7F3AB+iGrFUTHoKwbWvC
xPbGXYKMDCdlrLNVtla3kuT0QcLDEZgz/PqE/LMuvImvpPoMlrwN9uDjDEM5kbS0MhnVfUXMNljT
AssGNuMMkIc62+yeBi8TWOoiGluf0V6aoOhaZlc7CN0yUx42JWWjW8ogZ41ckTWWxBaQNkEKUZl/
K3lish0H6SnEkyOn01PxNOsNnc29K0kl+xFkQzdjVUJ1kk7rtCdouKsuLs6QMaZ7ZW9PWNwhsNs0
tgcyppLGBG7X82Ep/cmkj7dzQL59+ah4KfbYp18dkuLCY6LvZfL/gyr6xP0ytRoEZDh+7Y1T9Oxo
f/TH+TyanxwyAYjdju3YKI3QoKoxrcB1bxK71gUTQ/mRPvGBZoPQaK73l722QWbT6wbijpdGPw2y
oTz5Y6tjUq7MLuYgC/IxrGKl0vb6cr57YkpjxHVZ69dfKQBk8rlc9Bko42g9sT9XvoYCrwtzgjQz
P/Koto+R4JNICulFMEbMBmhRhd78bT3oV/GIkNzvDIrIXl3GDlg33xGDnHKgrJiEbPBx2oO4jzOT
obKZ+x8iefWtomHybgMC48nELHc3gqT9oEwBNwjduCohhFEMIFAV3C4IbZ6Y3tnldfBE0CVb8zVC
1z/8zbMfkrZo/E0I4px0L4yv12euxJrvAOJvNyHIXP4OmHsP7Ut5QDyI2VjGSsHbyW1A0TqEgWXa
BctZ20lq8ZBo9rHZMLKUrHLzRfwVV1EWg2qz7ypnF7CGnZGbCPbaedorb8oVfSIb8Rb5XB19t04y
moEI0uEgbDTvLokwY0XY7rsQ58JpJ8V5gFF+4db5qk946jIiOHAJ9EfdAWLXo6x+lHhF26nqaJC0
h7chsmgkGpTv4Mk5eBiqky1LSfyU4rJESFTh/KiIVNmxY9K/Hr/+Mhf8LhDYTfCeP0By+rCZu45N
3QnNN1vgf9kwinC88738/BWmiEEfhyDGFUybQqwvZDBl0u6kRq3p0PUAFVHdYvCv3C+fcHawYv4r
PBzwFSD5SuaYd+4UP9K6/ESBhhOGc2YDzU5IL7l9/WOa6QGDSVxAG8BHRb1B/NW6XYiwSbhkhoGN
rWfafCrE3ZLFPngVLI9ytvANwSvRYO23WffZ3Sqq8jaf9I9Y8i2n9Tk/W3C1OUNeSVZg9sPEPbop
zK6Pf7zkal8ByHQovT8Hmp/B9PLmQwgbwpiMxYFpqcAXUk949A1Ntbio7OXZ9yvFcp8eCem67EHZ
cc98PKSdPzEl+nZRXNAIKF6ZLEy2aC6Msnf6Glexgun3jXyW8Pqc5fxvMf6hXUn0Y62ylQGazBYu
jCcaRE5bLJeHcQXs9cafBgjB/fR3iYSwD725whLE37QFhoAG7xRwdGl0pR41yP/bh2YOtu6CpUs7
4DmSvaDqTRCQp/oD0S7uH8eE5y+ETyaQ5dO/7qVhZK5yxq5WemxBgsEhKZ9VENifPxFcVGj//YxY
DqqTk9DiiwjZo8ah8G9p978iDqqMyftViKxvxyB+G7UCN64A+1/5K3+Pyx+uvzPfcc1/zaQEXDte
1iNQhzc4xvZKCWMHKkMW+nVbpo/JvW4FyTJjPX3gEQLyR2Sh48IfL2Hk2TWQCDsIKkcezYQohYP4
McFTOvcR9eEjPCJSWEKNEnOCfytnaQu9U3MGxHHP4gnbzQhNHX6qbWyP2woj3O6z964REXQPf/Cm
GOd7542jiBaBumDMV24Ko1e6i0HHRswQFNNnBFjssxCnaj8JYF8aXHeRsHkD5eANYygM/Z5BROF/
agJQrJ92qUl1AE7JVqBkTXwtf/LAzw6Ie+c3bdk4SLkbZHmoFbH7F4sAtKB4itB9l3m6rIxkFY2r
lsw4T3pnNl3HatKImSKcQP/qYsCrX+HjgrVQd+JIPXWhU7Cg11udSpDcWe6wryXNqBOAP9JAX5jE
flHCs5MHtx5dM+P5Ri3rAir2AKzznLWrZzqvsSLanNzZ2mOeNXSJ5o4ddizmFm9YK9f0khFVgivp
31koOWNwiyV79jqRJTA2A+nnCl6HPEyGkYxFc4aZb2bjTeca0vHMilUINBJ0E0uDFIHGpunHam+2
h9q8kjG20rHkQA0TTb3bZSFOSbnv4zwHeOlH2LK+bRWtjDaG7gmMX0ut0guFvgde0G7+Zb9d+HA2
kfpbtHio4Y3/0yukXXIUwQKk/7mxyFL4bKitUO5u4NR68CdmiFui+ILwCeddW9eratNuLrwT4a0h
U38+6rfeSKBFYP19n3+Np+4P6vcbgzUaY5OIFuC5cEDXp2rleE/3yBQMuOAOJ961q+knqr52DvaI
25SOaAO2KZ+BNKbPhZKJmufZX6tlWZQcJBsdAQdTDLB0ks2an945zdcmg+e4VYdWrOufOztlGsc/
nGU9xOlt6DHladTHZN2NZoOvtx8WCprwm62VhyOSc1mlbcmIsiw0SpqMsiT2AmrEYvz6dAmUvS0E
sEmfBWQe7jyJMJuBUSmD6ppvUcXqD8twnU9g66P0l9dPG3cQ6gUEQzNCb405Rbao/KpGbZQG+Dcp
qM22tJn/IK2BrlSP/fa/ZWA7pXKiGg3HSaoi+goFDFGzToczP96b1n0bwFm6rdwMDlqrJ+xMteFp
gXFRm0ENx2ix8lhR6IRUOYDXjQMWNjVd6EFxOwICpglaSFFb5MqekxktfoVApzhZbKo+IipIrUIU
UyDLlwQiLNeLJUk2ijSVNNJYdZK3GepHdgG2koB73U7wod57gWEK4uuN1Zd9L2TT9JCZ42TSHcM2
qR9Y4Ww90a4PXy3XjgBD4YtJvl92lGDqvcE5XMyVfEHG13cZHgBamhi+8TAbXDuFqi/UZrlg5ORM
obHpgZqkLXKKlN3ivd40A2rvO+dXBSXeF6QqgDu7rIUpOSqVsH1g8wlleYDijO4FUOCgMPDPF37i
tf9J57lVpwBxJHEnA/bHrVDTM1PLZv+zDH9DE6a0ZEdI+UonsfueeMXXIwCBPFfAyD4ss0Wcuf0L
kDjnXWLkEddUttsWnEPNwEBRJfvNgHTkXTt/xIDGqlBruG0Pg9rYlCU4dympkK7qdhIZBvI4nqK5
JXlziW0wcCs+U1OTqKgntOhGR8/2z14Q5k3oNZMmVEzQuubKDaIWMqLtGhgoj/1WcfFEi1OfW9gj
zP0AmhLXUzXzPC4W0WKgX4BvgxR4DG3SDDfcnnkUWDzuCPvqZWZzrJXWb6h5L8X1W/nFOJLch4jo
qYlDisJIKjvWysYwHrfbl+GX5btwPRUF3kXowzU5eiIpLS/jOOJI1l8qIN91pRZNDrM5E9zmywz0
Ol62bdReZUS1gZ4246TUTh+jTv7Ve/8ikaEujiuzbnYB0eU1YuHyM7ntO2O8s4+kaWY1g6Wb0iaZ
cDv3/03TP0/pxrKxbOXn/fWUgD5GIDuOU+8/7n5dJ1FNcgZWdEkIIRe766d6Qj0V+EpU9fYi3BJ4
K8NoL7AowOSm6sU8ubte3SuivL+3uyf0/QWkSnBmK9Y6i4bBhGjUbt/cwnbVn75R4YT/duD66HKj
9C8ihnAkb/zjR9tVFirujSff6MbwLmC+spRUb/rYHh/VnGO6gLvOqxV5NG9IsoqiUYqOa3vNcOmz
nbmNc/DBWkS6pxjCWWN16Fu2x8rahMcuLR5hIu+87nMPGXQjA8MZvfb2eqKc9Lx9q9zFzN1TjjBm
JGtDNcUIJU4IwE8lyX3HPzyyWDVJ7XLJ+s+YU2PLPOyHz3G2xcl2ivegolTokShxiXnR9nGyv9Ro
EIq2WKCNdt4DdKoAGey7Hu2RyTzzGkaNFoCZUuAa347ebxJu0JzsSN7FO2FMZZN+sndOgstZTU3N
qCY22hh1Z828NR+DPPez9VzmwT1dP9Q/uS6hs7i91NcU69ouKwX7XjUKTKyc5jrfE/RyF1gZWVAr
nFWUpgjhvfMq8MW9d3UkoUn1M71OlAyrWxJYOZKwOpX3ZPKMSPWoGzha8OvehWqRy1eACccwjyyc
fDAxVAwbLVf6C/IqCcwgoZy4Et9o//3tMXCdwm4fnLvyhrucpU/A+VWyYU+WyJjhf94FhRs0AXc8
zpI4og9WJ84UuVzGyxFejiZqrpnJ3sg2xuW04gmQGUf6n2tG4CSL9B058Fq2teYvGibKfViA04mC
8yEF256r2bCKC+iJJrvTcnot0R9JAYwGbOQrywLn+EqaYkapKQ84hdGq8opkAqZjSOfmHvcCfZbf
UrbdgIdrZQX2r2mrmhEf1m+J+a8jOoh6ADSgEP+wKACQyClM2BWqF4cxv7FL88hJ1YGy7wk/Eu2U
BjB5UQ3v5wdl///zLO5hS9YmUdFY5/vq2UlD+SmVyczxzkhFJOeiDFfuPbeb1uQDL+0BWsTB7/xY
DM2T8twtuBDgiz2xaB4LCwEynIf/pluB6iXeBJjjjq2KkPpoRx8c3rvGSaYIqN5X/IUdAtWTZcXh
5GOgzVxKIte2pkKkBRTBm5LKj8f12pXcBos4v9+KbzpTBgHkRHjDptdmwEdP+KvOytdaZ5vfKnCK
1AlgFBZzpxtIyYlhTgm7OmtAG3eTOE/u2PutYwUD9IDZMWsmVuze8fUXhF+wjsw57yN8GB0T9gr0
Unf1rKC3L7M7vMLBmpazvHWMH8vTTB0eMs4F+g4cQxF+qZQVaJo2mNwWt1CT+MuPaf4/QUksVJhl
lnw/9N7gf9wzgPffaMkla2wVmGh815htcmiDkGBBBVgxoekU2CsBNME/W3/vxrP7x6fjfE5wRJyc
3TCfg/thfbxmsSKlOLoQBoyTCIlwhggOnHp9PF4WlKlh6rzX7VlyAFlg9x1v5daeTImMASTwuxuL
l8s7jPAliT4nhXUuxAKw0A5rHni1AV4bycHErecbdC6K3HfEwT7Dm6S2ryl1GIAy1WbIfo1k+Mor
40j06yLg5FGbtj6LU1hckkakb9ft9Mb5czaOj3YV0SYKQ+1KrjiGp3ZPYHxnzcR4jxTGOtuFMiug
+lrI3uxug7ahH3F+uI6QYyAf9M9Di8vRqDg/c2LHHi3Pm0o8+9HZYoc/mHt0iObltGHmPKqhpSUU
p8pYjHufWN7tuOwtMsy+6aYE2dCboHlk2qefGYqCu7FOAAL4pL9iFJNmZRxVER4X63ZvECzm+S7Z
0+nnSF9l1GB7hKaDxpjhPSHQK0EwDC772vKH7YkcvCtHuqaJxg/6w/mijahE1Zs0hjaikzM85o2A
C7dEra2XUHBeKvBWpHcZJ/37ISNXRKhjfGCsdJicPHpccmfr/pSSIwyl3qte8rTgob4W17GIoLDD
21qqb43UehBt0fapvv/8rZWLcy1/ceM4jEJjmX92GOC6lh8RcHONvywGLgvRjN8AuHjO7Z5U304t
Ma77EUh9xBpuo6R32x42usbUwFJUwACsn0ew1FhxQPCeJj8jg1ftwQy5DpAsvTPbu3Dwo9yZSgLD
WTD9CAOwVOnO4atEX+xSKouSZuHEOOXEQALae1Dg5IJ6MDSof/pOBrOcNVoWgv840EoPev/9SesF
FkT5SiPCPQmjwbmqgoX9UW2rQzeE4Z6XYEZaMh3uCP+62g1CKp45/zjoRcenum5FFvvCePUf8CX/
Wl+v0XgXEdnpxxzeNbS3N2Xm26yPKL9O2UEmbwn27/PNtjgrWS2FYAiECSOXD+0H0TLfv1ToUS++
d8rjZQocXLl9nt6tQtCBo8RjdQ1JlDS7FomToWQT7p+iC0enWiuNEacU/B1rvLLU2iiKRJEDaPMy
4J9ge4ENd9W+JJFEL/Lz/jZEfK9e/FfASSSAs0xpoM339NIBc62/XG5xN89F7Hll+PMDEEvxhYum
nsID8jbEfOvpVJi9dOpsYzvWvutx9rY4nvydzxmjM4Y63WPS7AFtnwrc2Wwg6uIuWBVWhqXfyeCG
UEiUimCi6F/0e5ZiZd7a9lEC4hH+0RIUEDchcwzC5s/RPZjZxf0iWrDkg3DaumIKnnihmtY3fiKc
neZBUN1B+i20ACs7ltKiCm1uDdSoWAYgbAKKfnSSCpbsxm3oOTHAv/xlpFPRyBVn9zd+PUL9Wvfv
jXg+XPig4NrysOrd/nljgSAjUWwTVn8232fIHmvIxp7ZUrjV6ZVA+5HJ/W5ixCcZq9i17sffFtkr
yZ5tDdGpJqR+sNYTc8DWhtI1OlxUjeTFksyFn7iVwWtyiYDR7Cwg5UaPpIT9RBO3FlJTIcAH0cDy
pT4WDbYCi579MZGAWT8UaL6AhEfxF52BVBv+B63MtZdoXHECzmFz14JQUgj6jrrkUiPSSi1dUSG9
aNb1rpTWFD+K5LFwqqmeWYBmfUw1CuzX7DwryUeeu3bDYdlOwKCXW0rVqiUXt7Nl6oDe5mTdhuGP
+tQVCl5YAQ2N3MObGXol6xBqTxf+viZqunApvqUIbUxiCh4doF5iMCBKxgOxD2jRWIz8L5VTkjmo
p/5EtXGesTqxrTeyMan2NoSUv9BY1CfnMHQFNKX0XM+ioFsnmrbFFti7IlVgfuyMITaA0omghCV5
LBn3XUpZpB4l6t6ma3dkNnHYoD1YbXHUb+4SyjOBAFCfrN0HiLOmif/+/6KxDB/qU7TYyYiA2f2E
PTfZsGKQRHCCJkZm+ho6X6xkOOzP5cIsOEhSmVozdRUpj+3aF4uk0zbUDxKXkY3TFmw0b53m+O7S
reaF7FVABMgfo/4axXR6ZWa4SAJFoqaLXYVPORiuU8wIfKFtQB+dd0ri6aP+ntdHS/BIgoQWoZLs
8QKBBf/j/KkK/sr32McR4iXAM58bkgtX9CNZXGRAG6KfS1hrD56AMVzEzPEGZqLhhOHTgraZJ129
AqzIymz2w3COj/Bh4Hi5j/9ixDmVt4DraVm3uPJxiYBCUcDL9Jar6GvdTRGGF+EH2O9JJR6J4WO5
XcFJKHDcAnomdEuw6YlK2SzS0bkdq/NC0UjjTDSgtHZuNjdEsf8yFq3JyPULOLnq+ONTcXvB2Xad
3Gc/W2LcPtQ/54m1UrR28GKYnEcNMwt1+GLUglyGVapE8DtHBEXFuWKwgOzJ4oSJpmEP4UV5DCFO
XIHhZ8I/+38HfsEh8ZdbBVSFBBTyTsQ0kaXjLcIzh3LFKJ+I2bbAuctVtSL3jO9NyijG2cRwakTQ
t2ciEbYNtV3FKRXLdX6eRalGqIAffavzxZDuWwzzXuG5IESmZvNY4qAfR33mMMDW6GPuMaMSebdt
2B5zey0lYmUjC3o7T6w6Ah5YsJiONR7SSFQpBdUrJsRfEjxU25EDq7vnNNIegRSEUDzT000OOk7A
5RuFzk2Tag8CCxutR8iHP+LvqM0zPvOGatC/7zfUu4KdxWwE2rdfwzwd0P68Fv87UdNH3GyEThfp
VOOzhEqWZAbH3MSSn9ri8dxOZrJa89HMtyX/CtVG0xWHNe5obBXHA5VNh5jySvIKPZtLt9LzDso3
SkmTLW/CYYoeApPg2D6+tzXPYqRNlIIv1G6eO6IFkLbmCEthHlc6M/KppNlPWlkjc0IHzw+n95HJ
z4c2agSjyo9Aev4UNN8XOH7U1trESGWW70Qz0lRGhRoC5iC5Y2iy5XSBV67poLRo9Nbqmt+Twk2h
fpqUsyzx4Au0rrtMz8dbK07GdGBiJz7hDZdILHqSU4j1Jjoy17nnnP9x8fy53kOQ1OOYSEHKe+f+
UMkbxtS58ATE2eloHcyV53axgOrdJl93GJO5Zysi2wXGa7YfXR9p+ohD/QSuhyTCg53dOOF2mlju
jtgfgZ0qGWEDH3beq4nKm1kX8zT3Vs0nM5VBluZ1CLMNnSUsloy80da00CcAgWNMdCpHkF+iqlnt
9aB5jNpWOqQKBmU1S1k2PIi93XV/fJkNOFpEV0c0EBV3PhCtVVCTgTEK1GwCwy6MM0VHKySliJJm
yq9qqR+fg64LfNX0sM7vj2jSmrJoVtmT0+sFupnGbEKj22TbIln+biplyOZq+lbh7byaZPyQnr7g
4yDLZ9VepjEWdwwj1OmqvVcXxezYTB7bR7oCrkg8TBKlda2hC01jqQ72v4KEKmwW3Ij4qlfJqeqA
myhO8qBuM/5G4+bV3U2LxjnXQPFqU2qZXmuM5ESXfSF/NKagXNIh6KBYHVxNuGFcxD2wesuGSM+Y
42yDXGexjhYNSoOLilAnWsNx1l3SLi8pFbQyzbXhjEzAU3SoA8G61+evQRmlvSgIaygiB0wgOnQb
gkpAvVZgy66KZpD3vntsOsIuqEnp0CpeE8OHD6C0Dtpvhcnqzf7T2Nghm8t528WRYDC4XQqzJdCr
4Q2mxZ3cTSI3WNzh1Zwwhfo6VTG1eDE3oNSF0IcztMewYgS1328ZDNsMAnKG5k2qjPwZIC9ngmT1
I1/Tu6lRyhsnJmNPyk7DZGN2a+kGiOqYpQHSxd0hLRGsALhaoL8EhMZOIThbsRrCMDr3wjo/hNgE
7WBAwPa6f7xImBvs6Sw0GK+gNba4FPT6H92mrHtGuUCciusLR91qbvOl+4FLl8nKYLnfc2gjxAO6
8r7P2xGqfDLKqeHjOFKORZJgZsrULzGUOrCl10Mecuf407p7eS90VzSe3+H7zXBZES16mOLhdDIc
R8YUJi5OnbRrU9WwMoQm1fU7JrOzPMGKnM8tRWkIJnGe5h77xOdkLoGoGFtimHrCNjZOOXjDTJw1
xveuzHSDX164UFfZksdSRaWvVm5tUWtgslauXxorPV5c1rWFwu2g/27ByPbKebn3e9ZehQ5QETTU
QAQCMPzPSXNpsYs0zxKpmWXVD3LlAsde0EdRXhHfz5xSQm5pCOK7zECM5crdK4SSGgwKl8b68rOf
zDWgRkZcFFniiKjeAA2CrbpC9VQ/N0qKKEDMJt8kdTekNVSX6rHaSNPYKdYDvnkYuOP6HuMNj6aT
1SFvFWcwnaG7LApYvEU1QNs82qzbEgNL5ZKVK7Rk2GUNyry5TH4yxVje1FoP+Iet2D70NqeXgEe9
SxZRZzVNM7acmlnWGxm/jxHCAsAvWcgB4Qx/Aiq9O5tIbVD8f9Fptky8ZQd8Wq8SHubPsAgqkxeL
F3vHBs4teQ4D4+FQ7yPGHlN3rvi4kGbcx6qT8pZope8XNqP5J8ZUGo79Ut0WT6TO3MAJy9Z4vmXn
yPoGmx7lYewbWD021gdPxC1UnzOHMIELCQHjoXxH61Vxz7EnTEIfuc43u/YOp/ujO2tZo3oFAUZ4
nApMtMuE0+Td35D4uRbpcdrvxcWdACyGTi4hrwYz0/4IqYIyKTwSKGdPGlT1yohkgooTWMbIEZIH
lvCwyJGvcl7oFvXJxyQ+0My5zviIADzKEGXTnU39LzZjOiKzKjYhM04pyT9Bxog9/Vkjrich0Tnt
mSkj7WiIeS71wSTzijuwS8QwZm1ZfeZWUh2Z7fvMAzb/iyBR2TRYLi+fTg3UdtEHezY3Fr4D48kb
9FxzEnj9SdO0W8JDWqe36O82itR29h5P0RWSoCdlWXudnJL+7YC8LRo3Y/KS7S1o2XRFLdjy3p5U
Jypbv1cN5d0M+PaUvmgs0C6ObZmtx8cM/PMegjIm/4/WeER1rg6cRrddll/YJgOAcefzYmWOTggT
s6J5PdDnf9hfXl0qudKZO7AuE4Lk6XYbibb2fvaKhhzZqLsNxgEc3hub3rt8ekzHvB0ZcuaZ3OTe
V5hZR9lxQtq53l4IVOabaR1Rd7JwRtcTng2IIku3U02XcGFrQxcgSqH46wwgWMYvI1xcpp1NZszC
yTjfB/8YAZjHR3H1NuxtGTRLcRfgfhrl/likqqDT670S1uBTMBayHpW9oprV6Ngb2mRzogrHYBSI
ni/7Vkrp/ajaBNFV54lW6Mz1rAKRML2jWLYV+IYRwkgJZMI/f6JZbBBzjhUnBli+5GcwgtBD1ZZh
ulthVBu8nm9mZGgjCVQvUFaRxPr2bqtwWTKkMygoRcAAKr0rjEn/KLVeP26bVmO6myC/mVArxdPm
yAJ3xC28N2lWaQ/jAJ6hC1uzXrsRYlwNOK1tpTZI9jFue3kfeg7IBExvZ0/Aa+UK+G3Xp+cT3vrt
iJgZ4P39MGreNiQr0J5XWnNxhxppbOUGNqTbFlzm8Lxf9zMdIJZx/Cc03Z1+Bu14PgMb5dqP0d8w
sOyy/Ii9fUtHueYYpxmgatmwaTF72+vnpHWLgZ4bgyxJ99Q7jH0CxVsxQIk4xj47bpb/t7+eiStw
blRK+bRzTA/kjYIYRUMSKTWowhmIEIiA7X5YaHHGRNLT5M0/LtD4PbyTLO9McXRtbABzaa86P8bE
74XGubl4Zbj5rFmzXIpaArJR41Hh4w+Hi/gYp4m9Xw9021ZYP+7ahG2yPJVWtbbJfEE4+zjVvnko
K+roXjjMqa3oMPUwRGUa3gwQMeHU63FpaknKJ4O1lSId37T87re3Dajglw995RtMFDhSNP+LosAg
Iw8RvcT74wSit6IpiEXexvSWSyGLA95pCJXhWFxB/B8uc8McEb90hDYvqpxyKIRIPFFDC3n2PKMu
NsJXLHySzbWpR5IShsgJJX6TEKC5MTl7RFVi+9CW9BQdsCVA9eZvfXZB2ApSYNa99WfxV+iX3Fax
1oAr1nukX5H6JBqqITHTZVfl8J8xS6uCRdVGl20G0MDCISQwtfOEZO3/7IogqmfoQKM7df+loLMo
+Pw6M0euLcuGIik9PFaE4WsyvCZuX1axeeiyiHmzRcujByWzkVFCbm9MTs7JaBvX0NYtvekSEVKl
y78TsU4LHQghqm2q8xgg+onh1kn/7Z45oTt5xdaWl7ePPUT4ZLG8EAjy1NVRL+OdXtqe8idbcf/j
JvQZFrRYOckUJh/S6tMQ3Zt6Ocip8A8S9ffITNb7UGMh2e/BXh5YPG2t1K1ikzA6EIIZsdGLyIYe
u/DrlesgZo1HfiPoR49463EfEQaRLvDGs4jhI7MnamODEUruEzmstB79JIPtqp9ru4wpW/YYER7c
higwuHYMx6vqcKndpM6nPfNTYNxMbQonmFEvfPJIFFwxlVKclU5aKL70aT7rjCUfDzpUREuT77eO
QCjAORHeMGsAivg8HD2m1qqBsSth4OtSAqW7omWCx3Fs6eLXrHDvcsoYbCcK6eAQXAcP+NowAotu
E+EQAi6q/BhA32gfn3flvV3rkaTw3CbbC830g3W55zrGv+aXYd1HFJLhhNX6N9vP/76/THjDKcU0
PiMxY8EDEMwTjitVAv1pSML9KmXTGly/lKi6uWqMzuQgda58GYAtvsDAUR6fb/8cwNrfEeVZ+QiN
w0b+EvHGNStfRgJ4aKZV1O13jKZq3Z1kqN0qIAGP2tGsEchhtWJfBQ3VuQoHKn35CT14fwUMOun7
pMl8PSW/A5Mg1zVdwdNDyhUFKG9/UXtk8J3Jt7xZq0g+dmblc639ZATBBxlIqIW+ZzXMRty9wqhV
LJyyJJa3vF1TW6t3dMIcIXnk9pU3TBfF81pfWDqxte6nc40Uim4mduK8u4oBZvQ/AhtMRK1jnEKg
BOz6SlcsfwwZvEB227mmytKWKUV4hwKf9VMiCHe16sRS771yk0CiJ5HTiqalyHuViyy3+YKKUAtR
tE3WJnMUXB3KR0PhZE2tnEa0T4IgwThb3T3TS918fhsrmsi98v8KQ07MzwgXkke2/0AhXvEYyjlR
3EuUIFkB3LHhpwAbGBnGMpw8PRtTE/5yo0QrNu9xoVAWHr4CuztmqQBG8dBBl41P+w3nrT1Zz33O
q4QbRGVmXY/BiWneaGihV1wUOIujbeOmFu2FpsXMNPIHpNqq9d6/TAVxM9lWg4x7X3LbMZCkZi/3
7OYIRIaRYDUs3GuypoTmkNE5qiAB3SX+OeES0MpPD+aO5MP8lN684/RPB24UkQIPDYOpCjFpy5iY
BfDf0Md15GTK6qNaySfbplb82KUnTPs/lR6J+MNBtdnwhRNoJmAadfEP6stWtY21zLX9flqMGqLq
irEtTXbPN5fSBMyMf83RF8AerhQdIXppDtvxdQVQf8XOKd+y7gSQDJ/bfCbovxdFgaVl/JTj8bqi
GTPe7Ar3YT/z3+Do/Mt4lfHoz9PIzSe3dM7CtPC8JUhfjgvuFyHk9E9RXBjgMHyE7x1NvS/xERFG
sVI0HyXwNLcMmzS+TZwyqbxgjfsZoasEoHpFZjTIJEST7REmpi3Hx0ZSUu8NJzDYHX+ymT9hUs24
UkNNhrqg791iN1DtumeC/Z05WgiFaJ00NlRJOtkYexIsgbzXcOBaZuGS5KUt14ElVdzwE/lL/Wnb
GHItvVxNzYMR8lB05DBOilp7wp/kadP1b3g7aIym7iLtRUgt7TZ8n9wqv9wPtJ7kkNgz42QIteVY
bSI5r3JejFRTxQgrhWkXDi3GcTiT8HFejs+CWC4zAesC0Nsek9jMmR0KK4sNZOJGtiohWnAVzrqd
ey3ESL+i6LQpJq83Ftdzq5PkA0emKkf1Ww4UjO6bO93+yzW3KmM1JjmAUuZYp2U+x6FbMx/egGEI
+SNFtRFbuBeTGAfdH5YOL3uMv04mD5I6LkGB8lBsxci3bh5I3U5amwDURxGNNwoAke6Ocx1Mxd+U
B0iUAC1bYGLAbJHRjfw5qMAgvRphsbHdMUEWIF+ON+XdlfCaqlWrukVWOFlsSU0mkRJElSbFXrIR
NMDsg3gtixQyvsoTLAler2mgBuRz7IVwbpmNJBtqiuY6kWd3lvyXHD8hApXXYT+IMPX6ChlNMzHu
BqoK783KtyxwqFV7age4lwB4noyBDB3YW73QWOTNJGIEy6g6yOpPqTx7+yh64ZwnOxWtx83Zi6Qn
UCK/TvzdckQxzy4KiNINBVcV4wNj/rbDmqw7WNfdI50bN3PIFPtpkr9C2Fpcuc1EhAx/JcUpBPbk
JBH4S6DrUVRnAvzl8Vl0mKvGxbseR41EDVq3VCtl+lpWNjl0nMYOqsbgm/ZJd2Xg68yT5JLP3f9y
1rdxPl35Io1jDgENNyKgKgwiGzu4BZRATF0J9OJ/+KAYWixdPFGGMFrUh4drwNaedoZPozqDtvbV
Yk18T4hli3ZG8YoCzJDx0h3LA8IqkLwzu9pbKMk5XpzlW+YoyJqXIAp2BhAYvDDygrQ5eay1sXUt
+pEjj0oUItMQPLWZsN8nawnMp2B1yQ56bYsVn5crY/tcuwD4Bs6q//2G+F0BZ8/Syscbd3B4gNf2
J6AFMG0pZjsv4oJWkJGv+eN4kbYTGWPsQgK7nMaEL0q2gXjv0bxFs5NGjjI4BrAgMQ7Flxz3eVr1
wB581iHG+3h56yP0bkvWvvDV5xj53Aimr3Zeiw4OOVXYB6r040azoPPuZcVPKJKcysaqHqeE11H6
CFT4ZsHGbeCAukFXpan9lbRRFcIAMcUwSQByiIWaoPiBbV4N6IdsXjLcZxMaen+BRSE106/0Qdb1
B93FAfzQXMfsQd5sZBoL7vSfEjIiZ1vgIzJsIHzvAq5iZvpxGbW56dUBhgd9lV2mZr5zvRUt/aVa
y1PqVft0/cQ2NIFwbh0gyGb0Oj+dUhMSpnjVFmnpOuqxMpNDA8yLvxxITloj8k8bpEVWChDmhbjU
Mw3TPZE5bcR4WVq06Oxfu/jjPeYBN0K9VQhxgv5T8NUPQ5Hgh8iP3qUBZv6Go82pPgewy9kEuuu2
rc65wPKbRFKjFJwt3scMCoWF3NjhnpwkKiLXX/w3DYS0oyebPbHd41FR0jyPlgps6LtfQOARaVPi
Z+zMVc0yhDsrS65OzhvVp+FVsoJ7UTvtaQ2hzx9gAJlt+ZWEocEA98qPwqpndIG9GIVxw1+EsFMe
E4FAWegQNVnvC9XU5py9VG/fFMarEHethrGMs++JSLWZe20qaKoqg2p2qZS0MCV6r6T0XhnHF/WU
glF0zPZG+SyTp9ULVuFSJHEtkGFI2YeFcOPCm2l85+bDcTBOhmgiBovcleU0585fX2aboAU6kwhz
0Z7jY8d/V3Rf9tKxAIeFoWFL6S5RufD2ZYZLk/i22BxCB45j0D/BkAHqxkYzOVoZT1gvcIP9QGA2
airpGWIiiUeBrZytWNEl5A4NcbHHJ/S3lf5TV9eToMEP9vX5aw2a02yCCrD7XyHAIEgdMM2ivLDU
/vSpTWv/eyU5PxT++ichN3/436V0WKpOAmNqoWfL+RNlr7WxmhGM9VC1jhlB18twnuHFcwzakMrv
i5ngfqNC5ZBj8gyMioeBT+ea8o8221GTqYQdIuTigHbhTXx6fZRpZwvyPgT2XtryM1AxPtRjhFGs
zVqQSCoh9QhNVTlD0h4g/CCh4HphzonCbHopzb/A/J2S/xPa8G6t1SklktNSHsPuk8wUnQlrupHN
K4EniQBhNy0fat629DJGbdbD0oTWqd2mA1OXvqUARlWzYaukl5+Kx3CpxRU468K/H3QWfmvH5/nY
GTuyxnPxZY+C78Rc5jmSgb7RUuu7uY8QGUgpow4UvJ6ApennnTk1LYWxK2T+HUvs5lSROVUFR88A
PaLrVtkZR6ki7Au12+L8VQLQN5YvwXJWc8QqNmhNQ8D2x5W8AX5MwHjejJCVEL6L87mZh5JWgP2O
tqPU8Q2sYbLXsaNAHnGdt/lvwALsWPW9xXphSplf7S5jJUIxqrSrAM5Mp9Mgwm+s/OzSDRk4NNk5
mLw33o6IdHmuVMlaPVnHzIEV5Xer8OTi1pS4aSo3aQm22vo+G8zzuDW3UeQiYuW2mL8TUq+PYhqh
oPWbSefPzDo7GfEpVZr7u9aI+Wj5HWas1qYTGr7k9PGG6TwM7Beimg29jZ9B3RX52U5FmM6unDco
sJkmvLKjoEn/6I/l8veZ1SUnXUKEU1bibB6EtkgykRuVaglJ/pK45sSFTN40avNn2BVBosvvncp4
n3ueGWpQ25ZmufXz9eWFSK6UOHVR0Q2IHGJfA4jX38L1xqBM3c5r0+87kKkGPmvpCA2Ahg63Rwkj
xvWKfCl6sCnpanpaQq8pnN1OpP2ZySF6eIDkjxhmTGqA1f7LW1/8qipqMl+zzh2CqLc5ExiP1VwE
2Ytd2YnnnHmCMWzwRv6mvOGNcIy/x47F4e00DsZuiTlp7SawzXjwtbA/sZEDx01VIiGcEjRAFUt7
XmDqPUkQZJWUV+Su1iqKMvSuJSiKVNKmTuY0p9tEyT1U1ROhWEHFdKPUD+sWAtxxbUZei/QEYMOD
B9sTluQrNKSAQQLR5PqizVzvuqORsjLFhpEGc2wagJv5E4We98RlHC2Z1p96Rc2errnS+CZSvKUm
bxKrocrdDhm7GYMbIQJUl5qhzQ+/Df6IEXikwi0Mvt8EU3h5HzPv9v3bEma9Hp7KI1+38o7u5AXr
9y8Rlq2sHfoTorWUDzUOMSYG1A7d6bwNLXEgE0yFqWTW83ERyR63qCS1+a+9+Z2E1N8fdqDl/Tz/
ieHFat8TOTvn6eLC4ENikf8oeNLm5/ZJdlZM+H1wLWDluhnxHSNdmIC9Zf6n7A1q2WS/DUxeq8G+
ScveMB+9XWpTKlkqzxQkMVI2GhZtdppkChJWRQdCawaA+rWIrpk4GAGaXL27x6yNk1wNfUZt/oil
+4mdUgQspTQo2clf2Blmjuu9xpYfBJSVUFAEVWhDfsuByRkChBLsWhuNxFuxyQkmnxSJSgpSOby2
RCWDStJy0KFG53JRggXXmEhYa9MC1wqrY8VJkkEk4e3AE8cYBh9H0WAYvOeaT6eXYUW4w57EodC8
6jL7lsQS7l4PgMu+wfy/Ryq1TDc3zwwVopZ1h1rkRCgNmKY3KdXpyYSUXBSaNN2OwXyBwqVJ2zE9
W2UPWRUDCB9mCvbjtGK9TEhTbERHRFGDt5iDqcWCQjuuMtkoXTLV+uiPKSAUQc41KXR+b25rWvhO
wfAVVrjscUOt+dLGBc16TphRI+dX6yzc90lHHeTh4YU/qbJrOIAq59pBTTnEE13ApgCxC7SLRhEB
0kV+zUwdkm5icJ7HmbflntNqbvdk9iENyH/hGuCIOFz9YI9uRi2CGZvDJ7t78fmUWRYR2WouC7dV
w3YneSlgXbjLuyj4GJO/+b6TQQogz5zvOSLxNpysRmdl115nIA4k2bzEyb7Vq+x69sZplSTrkIzC
gx+3LylIDvdmigBa47BMhAK4KVm+tuD9EtGzLNahnu+FtqMIc+whUHCDV6S9b/QNTx1eeIYPqGd2
Rf6NUeWku9m7SxG0GuqQTabv0wTIYPqvP7teOBk3edrrwE2zCKzOyQynCTzRxdSVmVmC3RjMiHuX
pLxyu5iKtUDfaguWiIjzf9BOY56qH9d8H2CVUWiCJJ+3znt69gAxyLg1TP4IAV/OZboAaqIy4/lm
nxtsCiiotcmqBEP/Dtb7Ss3QNJIGtmwRtO5uxG95sNOO46GYyT/EdJ3ZIC5GhM3BEUnnIF8D9L1Z
odl2n9Z/ly2NqssJO0y+zAF5Gcv1WsyR5+AI/kYnH+fwHgKc6YU7fejkrZkZ0OHl1Y5byXeCSUWW
ZQ6qUn+Fb29PF49FptpJaNy1dbM4XY15I0eW7Nt48WL9dq41gDdHeGZR+4d+Lpl4+bQJjre5hDZ/
ppqtZuCwg9s5jtTAAJFnLrvsAiHvmWvvgL+9IH3J+TNbG8cxJTcQh6ulI1ANV8Dpqbn1hL/aXpdS
d3yL+Wln61ok3f7tHQLAejV/0LkTxeM91ql8EuVzLtQLgjppGmRmScKH2QnobAMBtBt1ivdoaSBW
9tzQrlSccqHD3/Ggb2P+36IDKdNpr6M8z4jlhlW0suEPZLQsUxarg63qXgoQKy4JYUDp9tenApv9
O6VGVuDhmSvCTiugxZ2W3z6lsxkuoA2QI4/Tn+NWG0RGywezvk4BnngF1St274EX4fpB/Nyy1h30
3BGx055U6yU0vVYCWlETls93JQLVe/eldjK73Uj9cwtYozKik5qXqNFbcRjsovudmowGz8F1CfIL
6KcJbbVy2MGZ2jVZ9GEpLtX/J4RcukHZAoh20GRPq9cqGA0n/r7klX6K/tzrGbSmFLTlWAaW6DGQ
L8Cek7/wJkJJBxz4hA13dWkeca0GaAT2TLnBYe1LOgne4sdHUACgU2eorSYaKEHh9xEcThFR084o
iQzviTzogybY1Rlb59yNBC9qESWlwDe7/GvUM1P2374tMd8lymtd55YnZ5hMO77O44o/HWi2ONdd
nBbBmVNNtXKeYs0668+9RuWoMDDlAiYKNleyYEAzLLFMYmApNfwLzlx/zoiiEGGyoZ4j3RbhNYh6
Feg6v1GYiUKsCIOz3CoGlNMC4ZHy/5eMuOhM2hdSZ98uaCujhqH0+xFjJkwutUKlaVzme2OO3YF2
yoadE44iRjE/Blh0PrkGEC7Arq3wBTvNo7iLeBNt8mCorof3RZbov0XShyvL4kW2KQ0IYcXUqwEJ
VSDsZuV4ZLmPm9qK6wglzOVkwJO8Ay/i7bRKWPZU8PXBBtQlSfvh8uh8NAELRriodTNcskaabAIa
uZMRfdNPr/cPsNnrjLlqE/QTvGJgMFjvpj7r1PT1TfADxdC6e6d0/nPZMSXmE+HRJYYwHoA81/ge
SOowDH1rTLKqBloKi1YD4SBjNcWCnP+EpqhU5Q1stHsVjsOGB88My8PFfAMrCX5iOffte8jqPt/q
H6wn82eVZ926jR93hncyzoarJpE4QMFSfvJpEbDJWsFy6jYdj+fsocbHke00EG6+/y1AGekjSBSz
bpNX8EYoSXf+WqKcj2Eqnsh8ahjY6hasmTbDj9uaJNrTSIfMNLiZrs2PhcDkR9KZb03KIyrZhiVN
UnqLKCnVZ8wrYIRvm3sBBbmQF1tCNjMPa2/xwptF82WsVlWRc1w1VY2nPnYIhvNmcdYx55SfmgvW
MOOtH/XYJYiwpKkmTBWIoZA04O1MbHm6m2+qmqiMoMpTDfQQyPhFwpzDVsjDqCdSKMpR40aIt+he
76PPrLuBlqONbGrXCB+521hA5o5iiR7Iit9yOLALDO/uvgQ5IX7+7i9MC70cZkzpKMrDyOK3MOGY
FG5h7j/4EUA7Z6JUnT6JKrDGpiZ1o5zxFhOBR49Zw2THcmVSG+rjp6u+Mrkj3j4G6N7OHvh7XO6a
pGNAiygQYZWReq7ERZ5S+/GiuogfzcSKjCAjgOoYi5u8GuU5eQ5BKxc2MpdqDWdF+eLa2M8KT2kp
l4Vs0guyYWnxBzOqYL43TPden72bs4vVpa6zoJ3oEJKslttbNdoeZaGw8VoSbkYXUAwExckgbB4s
whjOG4R0u2TNhu5dMEl24+EQn+zS17q8teMXWxVI+sBTMbKJOzcOkMa0kcJrxQpcC/1QAixunmPi
5sT+ljVby6/A4tLMrsuKH/gUNv6lXw8Xv6zgdedfIkR3g64S5JIlVL+mnXUvvOQrsp2TjyV9ZD/j
5EaLDq10gs74hkBbBj3w3jXM+TvaHieOOWARhDT85t5gYbROiwP0R5rjzZPC74gmXZ+tsZ2mhIFt
j4ufoN4HGwuRKdJfKckub/gU7hyJJ1P1naWSiqDmgLbmw13SJpAjoHgzZpQwHZ/LHTtpP6NoHKmW
dJSAidenLbkYK252RgCFmdSV469z3qYeh9vxGP0k+idjI+8bdbjokipuawpfYwDhLBlmadZOwaaZ
YJ4QMmxtIb85u1fuJlehD12q+baef0FfWh7fXnc6DsSqD49+o3T+t9VXi1B0bDG+XqbM4kQ3mEnB
ral9KHDe2uhs/v4jREV682FEd3/W5NKnhA1PDJXmxXGpPYZd+DeSeFyEVTpo02XGE6eU7P7Q4KEn
fInXDF3FgZjNdZZomO8GKB33qZguCAuQ8mIt4do+OnqyDqdTcgPDRludg8PCwxjTsooh3M2X3QTX
2ArgLe1tzPE2JYeOCi7yNe0wVDcX4gLhOAdblRRZpBhT1F59ovuPVPnRe5qPsh6qRb0Z+xXUCjaD
F9bxlNIOJ/lbZQwEzxOpSdchF3H3WQeiHPAD/RsmPKvIwHAC+dhk0eN3WCn2YEjeGaaCuM2GJznQ
+nHFLUCxYzwYvQaekL2WGjDllx2Z6FmUDsFt/Xw7uDKcAzSkVMb6bUrdvioaTXT3K+4ihtI2GV6b
u3E9tjf/QkGk9O31UPkFK6u7uhfTWZOeXcoL0CjFAiTM1lCiuDnyHRYLjN/d7zHFvbAEI21WMf6j
87RBWnSa94mUrvw3nC72bQqYoDbz7l19GvO35Se8j0YfbbYbfkNHdpZHNqOsbamF86NDLgMPylW8
6XkFIaGp6PJym8qQDWKNVIjOgrKCyKU1hUQBYKjd4Nd/c26eFLenwPGQ6UHv9HUUe/oXBIxGDWma
3PGDZ1aoPEM3ObqMK7dQnvaxCdvgJj4EX6gBQrZnTPasitrnBcKEDQxpzjOVZVSCLvAAwiQPkrGS
HOeBtiiM/9YlgWS1GPxqbJ6XamiwXzgaYueXzVipwgkfdRw8oLvY3sqD0hgTEfwFth8WRXBYuDxl
+FEq8+tEmLW+W2Lz1rcUdiSzcQNl38P9Y8y5bG76M0AugxjwzUu9kzeMFIxGDkC4nYMAWFv3amGb
m3nZDDNapxd9wFbFoG8JVs3+EVSmlda7OTUPJgNiWg91CXpi78O4F+STxcmMP1xKf7CkyrSZWVZc
kAAp3tWq9YibKlDpTwrbNBvh7oXgRWdwPTbITZ+mAkqea+c0tINymsNXhyb8q9dmUgBzvgmyPBa5
mquK6kZt2/MrybHCzAN8uGEWszs6NncEnNYiOnPod/P2zcYWDOlRY3pJ73PeWFMAgVK0hLvt9LVV
MuCz33o7iQ/oWOL19pwz45pc/dpLY3iYodvR37v9vt4yRfWPku8Ko9eziedZhB17uOtQqyTiuZQ5
HZI0dqwErdZTkGoBhDY3rzqRgaiaF4YYERMOQOcSnJgpJzuHCDvzlI6ahSMfI96KpbIYs5/2z7gf
zl7Yub55bw8ZoKrQlrL+9wOxDCK9cv1rN1vM0rAMn/ZOGut8f7DBzYW4bt7dHLwsqJB6VO1kT+o8
bJTKUDlsF/9t9DtBxz/pUYomYFqU98Hc1zXeE6b/35lZtKh364ocirAO7swItcEiPJJuyMWBqAOb
Kn/Q2XGmYgCmGXLUk+HZfzokUKX067A11PdusNbNNq6pScFEras+OMJjwoOZlDv200bGyrf10w7r
4BIfG2dBroMJ0N0pu+KWtnqRza0TePKofm/4UT2nfnWMzGAABkVzCHwnXQBs4M618zxibPIAxher
itSmNTMGfD3jKdBSBDYYWA1qiLC9TWgSkWNnqwpztjkDFLGS8zmexqx82oyf12Qh0eY/i3reGPeO
pkrdCXZ/KQqf3QxbzVYwte2xqTjj1PIF7LAKOWE6tHd1HQhbwcbdxMyik/G5zL3UH6Fa9doxFVL4
ZDtODGDPsNL58DpAxXwRFz1pCEy7mIOMK5vxOtslIrOl9RE/M1tsvZWRI3HRpt0S/hOYUaTTdGKm
h2qGAuzdWRhp+1xP3H5EEt9QDxjY9vkRgmyeJn5obpqlMYhVxEeHIIWPtncEZDUbcOFsONPF1ddF
M5wPZqdxnDTsSCPg+06wTvIk7IGol/pVX+R1BL7NX98OFLROu8ljk2Dz4ZGALYhO9WyKZUHYc5bL
TwUJGdvUWDq6WZ711xjeVr50c0pjpfkk7o+rzbXHDtMk3/9UCc2ITlls2G3y+f7rMVz1a8tYBP2X
vEthCLvKCOsytpHHORztqXuysroRDoPqgAQJaMPr3CMHNmXCx3cTYjhFH00cPt45S2TS6D4euaSR
qrLP1ihRlgcZjhDjIsYaNs8SmTYsYAPKFeNp8RSGbSDmRg2BGNMxAAevjTfapzmUseNjCBXlQrvk
iWbLLKpA6IdZGnuTIYvIT+PJlcK2MhDTAzmJ1w910jpjSOTkfTm/tfwmzagftRI2lUkqzAt4l75W
3nO/xNHc0FN7nv0JrsPWtVC0dwiMwnorBhcDgPOiN9flsl86NU2uBeeNCbj/HN0qtnwxqSbrNWbL
dxcyEnMAZpB2NDzKHIbivS3ltbhmvRpMX9MlBs6g8aza26p7pNrBhaRhNBdq5Iuia+8yopWwMtOW
dydoV0fDqYVXE2iWob0llEhIGhxaGcY8UDcRdyWpv5p8fTxHVL10sRNIYfe7qDBVuMCbtRPymbY5
0+hBGIo4qsKvcwIJ2VRC+TFbep3EXc30MY2dw9N2Vypy3OqMFijgDmrbhT2h0l13/2rWpVVKxob9
gu/BFo5pJKEbcG00LDqgUTz1JsqMGwZYBMTdIhQv2weNeNfdANbkchJUmpm5fIIhur55INQw+SXT
6lQuz6iBe4WdqeocpHmCUQNJMPLHNvVZdcQlctgSXchAu0508SsgRUz19xgIUt3C1dycg95GAsdg
NO2V4Wd5bgiG9/Q4qSwsAF23H+sdry8XQW3Ug+7u+NPIbmAXii8zkVZ9Q5dYg0OcgmLerKH41HAx
Dpu45sfLE8Bw6dk12rPMstD8Gg7Kt4HqKIX2jim4jhcBEo++j9/LD5JiXpNFAMRSLCOgfzKBsqsw
SE/WanYcmnE1lhEu1xDRDx/gBvtfVKwbZxgFlTwS+7pb8U3z5Q5GCwDKqmOnUqXDgtDN+OWcIBeq
2TqI9ilAjLuFWAe7fSYtdhrkPVlOZh6u3//AowyrMAgOIyij51jFYcWoitJLIuDNVfIpsooPXVH8
womU/SKmQRm9Rp/G90691o9hJRKpq3RyutPFYQhYuLZ3OtD9dWDProN7g+Cj/umJLB+AsD+YX0Tr
CcHRLDsP2Phli3hlY0v50UZXJf6wYd1EiP+87TWZGJPk6FrFsbYsRwEICVpM5pZZS2vKBdC4xm9d
Pl1XKIJUwsyOdSBGx8D5nKWyk+IpeAfNLag0s/h5yzAUldsEDSyRY1q3q/kgDXd7T+8dpP7fpUcx
D0r7fsQgDk9k0SrZhImSIqZHmcAHSRryX+H2MX7h7kYm1OHRL3dMh1nbhJY6pjAWrxI0iis3ALw8
BzLkuK4SmLZ4IHzkGL6shMqnpTWZjXC5uc71gn7FFJ3dgaJ/7O91VwdEKe5Dymbm47h3qT4Fa6H2
R70vjPTlkkFObyBH/ROM4Wj4XL/E3GWAjuvAUNj31MWF8p0TNQScXa5bxns4VJTx7aciJmDTUvU0
fEh1NCwXSNhCVFTjtatx4nvWIxVpsSryJrSNNusAjM2lnZ0AX91lM5hw9Jl8ffEGDLzMqSbl9mFy
ENBzDMAFcQWNOYW+e8ctPd61qSCpu12BgG/Fj320XvdQDYo25PcSBDxeEYoiJ94exkyBF6iUVVE3
9Zvbju4WqJAt2GL0WXsjOXSKzVvN6bF5T6ppE186SqVLKmsYUnDtqV8mqAjbq2xy55ChRdVs4QDA
LNM6upGsTdlXMq4XAKNrzAEozGkXl8k6rwmmBm7mjkuzNpdWRgrMKRRiZcx2FVB9bpwIxbGN8LmJ
zpCRlvoGuFgkbshP+ttivCCKGhoQ8m8R1GQMia1kGPSBdV2/KsKGJL/lbQekn7o3GWCyoiw0bjRv
teQnXM0YoXX0J+e1jx0W26oeUIVh5pItoh//R/x0GYwB3H8j8ewQgEgwSAOljPp36kIM/mA4FUaR
KD0IzrzAKY77U1iBbWtniYphBWA9B57/hknpq8LJxW3b5FmNzLH2L3B/yW5FluMulAfGTOAQczJf
cREatDCzmcL8ZfcUzNHd0XFYZw2/bY4Milnm+RAInwEAqxtQqwu6dntvblkjMqU+Cdc/ch8CSMnS
y91nsFx3y4fMgTw2xL5i9bH4w/hV2uSY7etBRaSF3ZvOJ444d/tfAZx8FvH9fuVQHAYfv5orWrD/
PiDrIiULFUEUu6AQjIEcB5HhZ9chB2kyqEeYY3cAYehqzbl/tdd/vgW/uyeiP0rL8S7kL+L/6xvB
Y2yJvE2TbVAse/F64n+smzWrWzDRVSh7Zo8n0SGO7drXVPSI8ueGz05S603GGSFLISru0Q2ycIfI
nDp+R6MP1zBHIiaPyfDYqi/pMSUhcu6oV4xPRLTi1KO/gcrgA6zfwXyxUxKoGDGujUrppRPWf+wl
cGd76a0nUDSKoYjcq7uxng9Y6fjAJNdRb4qvnA3HUIme6+92JLWirjYqGfzsqnRUlHjBYYx3XMzA
08aI2Ve+wNx3MtGSSmRm4eCqLOFcQWm2XJzacqita+JGDy433k2bLBbx9IRgJjuYyNNHNpD5xVVk
eFsRR3jndpQhoJJW1AqqK2aG2gj0yopRJfqqHqZUmGc8/vdLZyL+QT3r2v52KXFma4WOO2FwRKH9
8/7qI/haZHJQXiS2kmseyiPN3Z6T/6leX0MmZ32SaZXSDoggBovTE473XG8wcX6C6i/ogCk5bEen
DO0rHjC7iDUA8FZDYxyLldMqZs3stTTuXxiIUBS+WvO5aI7v08wclc9z+aaPp6zaOx7QFwsTnAUi
W/mRNIZS04In4dZtdMrDDT00JnWTUxkygEwyBbJJVzwKRoX7JvcVSrz6cu/mG+U2KsRuXntIAmaG
7FXRINcLlKdQG97cX0LOOxpjztKS/NZz+BDMBZPEbZKJuf81P+bypADCzZa/9H8D5+Lz31vSNY2Z
XCmQAl425UoIrZQc82CFU1WWPbpBGqul5x4XnELGzTLp8eXhvyGGQpO4FLl720NtxYZrWpFiNJzy
QfKSWq6DgrRoTBoJ2aUXuk6crPcQLc4INcNmJTwUhSeVsIPZ4vqZeXYo53+nkGWU0p1dKWOFSBsb
m4k629tx5i9QooHsfHtNSOl6iekTlU7P24K2y1gK4GHlvmMLAjhggZKn5zPqn9IzyvYGvpuPRchX
1BsVtR8ptQHJ0eiMO3H1BwORw5bV6wIUINq3KcbUV4DSmrBtfyBzU2Td9o1nLkxF4mIamC351MwW
f0X2Wh2H35nbIgPrVuY2GNQ/4aDk3mXY5dQ3rl1xbzWphKtXiNiKfqIYLaQJYCbAqG5BlCkcFkTC
xWaMlWYSwMwidKWseo+YgEc4qotLKbJYxgyBct9CaSZEZ5QvguP0t36XVMajpoo1Cuq/pswp6Y62
Mm3yHLugEad2zGCOwuSSndRnrdilZQKA21LTPEU94rgunqdKMEnYNvG2Ij7P4VVT1bBqDOIhIsZ9
mB/qj68lBB+uJNQxL591ZpLOc64y53GOcZrk8xrqOsfCvrS1y5qx8sMnrVdElCuqvDhFDIujAzug
lbB0hBZhXXZCObk25H7NSK3OUxLmakSZoLK8VBixKy5b0yeIRZU1pzqBSIJVfE79+bdoUjO39aO8
G2CSEsE7A6hhCI0KLsFHSe0eB/wYvvJ3lNYg76bDk5TbuOo4lmJP5FjjtfoN1dX3gQPekQa568dV
tJNMDvSp8Srzg5WSA9ZfzKpGGI9NWNeCQl6zamsIOg0tQyqsOzYjEKuEvIRKtX03d/o0MKCQYKoo
9qARzMl9GJT5ShjSZj2Y4KYNsfMe2uobEDpNB/9MOJ0QVjafrEh4jkHuaR0P/Ev2PfJujadf4NE2
1zlbma5eVvNOiJdEll+5ViXufRK9T5l5C1ZD4IA8aP4Qq4araL70HFBsdxDgVJc76qPLHy5TK0rl
UYmcScqJfYn+URTDCzkTdZvnna9g6gw0QhHaW6/fgcqVzRn01SvYJwy2bxyRGrlCJ5cD7OhF6N3h
oAJWGb3YOtSTMgkWuVKYKobV/IDUdgvojvDNu/T7HWtamn1Ncb3wkNaPVWf+b4C776PjYqh+O/I6
jW3DnFI4EIDjIUL0XPDfgC4eC4Rca9fESwDDHWWkbxKbIsjXO3wp8+xkF8VSISnOD+j83sFChr5M
A9ps5X8Lq9fxaZQr31bCsBnRSJ7N+h5ABaRDnEyDZ9aIa/NAjF4WmpqFmhczNghhHBvz8A0wUcsl
wqnQuS0K0Kf7f+1uLLZ1JkLzWRrZ84SJIndo6gCReLnPF+dRKyDyKgYKc8cr81JZKvavwvNgPKdM
K+ze8hAQ4OjnUVYrvs2iDJDC2BdFjQVYUsY85zeI1hKOmA/PqknEwoMG5htxTNKuftu+ckk0rQw5
VwGFfao9UIOuVURfMWKy1ERBLZXtJJ7R+AEK50t8Rer+SZDAswtpfdzQAAVplNw9WkeH5ahZoKwc
PwMqp7ZxnOXq1Y7YTjQkH5AnVqruMKDnc9kZ8NSqBontyOY7fsDxFXnUiYq+1547GhMDl0kskrns
vZexYZvBriTFalhC9PbOkYM8sWVgmIH9ENtkES6I9nx6SBFG1Glf31oAyvmgakld3U7RnRyAdCuC
i1TkGeG9MUS8C3TEkYNzd28DGaNVeTkNvwVD84YJwb6p+5VRni0inKLPgO/17txtznxegf0ujbhU
CCtPJka2Si/xDee03sq0p69i4tadvx0jT/Y+TyIhtWHRy6qiM+J8QDqcstH7RcZm8n7Inxbo3cSM
idCzCVPjsZZ0+yNJJAB5QrAczQwg6MbqDhRzKndBucQiffUWjGFLtv/1G++LgPJcm9b7DpK+tDvn
aNnBEbxLDWpooIYneVgl5a/paqSJLKNci6Qygs0fqcNhS55IBmlnRw33pqKBajKroGThfQAtsghh
dXtbSxEEW8lLKettZ18iKvaw72BodFIyZuIUzBhYAAOur6p7Q1LeaHyTJMoZwZCEAhjMO0opy910
0p6n++103ItnffR+iqBd7NvCnBqpJxeIema6MLehTT1vM+uZgwpuK1YHcmFWpqL2CUvNguXoFhwE
Tpbmck1FQPs179Lq1ieZwKxRMvGE9UMRpZGYoNpCpszcPI2V0A0lzOz2J2aV8j+yaJG/4r/7McuK
q0IlHClGNCWuwyngmngBh/RfjtHh48SvLldxeA0/ifHYSiIoHGQ/opiVp6u8Te5F0Ksasxk137nA
iMHkr4eLXPaYCNAioLuPtHCrj44yMwhc3HDxfAuu4dYez2W2kR9qI46lBSwcOc70jzzqDMX6bi/i
cNptmQRroxXMzmlQKxKzKI6d257iPgh0J7/EGuduoR1ZWWyxdKIYjDFK9P5W+E+BsmR41gw0i2mB
4gxwdSRdA+9B/ppuixQKJwDY4lE4POd7CPf6NBV8pe8H0ONSMpA1EJCz3ON6VjYBG0b0Zz1oF1wZ
XgDG4KP3kzVgXAqlqOVcITo3f8+HCpvhpWul+yrjVZBnlXGo9LoQ6RLy79iLt2h/cN2yT8TJ+YET
B8Yg9pdK0MQRgo6Qti1hy7amTK9p6ljHPuu1Fmc6LuAIjYgcZ9exsfVsbMVvlAEJriO0GVDe3/vW
LJior8+75nPVlcU1VsKg7xHJr29jIw+9135KsBRhuH3SokoaAcX3SneW+BkVeH9lZiV5iGwvK+jY
XPI15yecEvvvHh2lrzE3DjZfj9ptSmVFQuTBR8jONxAR33HZ1Lzoe8UDMZokYk1JzFdvBSQSooqb
r2i8lhsQuMheG8gSle0ou0pJaPBVg6NNtZo13gaREDiuGVSR3MAYYFfevP1aCFS1Jli8QtFAQQBp
TdcImLkiZlWEznS4Bj2/TKLQeAEZjcBPN0y02xUK0ZHulrTxxDPNR5orN6ds/Ml/G98dc4jfXnMT
jLJDBfTD/Y/q7UiIQupVLc01/5MhI7Zu6L9Au8l23dtvefMQLgjiFy9nAB0jLuxnZAp+6oaolzgO
t4p8BNDAzYshNdKsl6QhxF/PutitMykqpEynOuRMSftoL3vUhmKkEuHvGvuFh/552WZ1lUFpw7RG
Xy/cKpvTLc663Md/2ZJzr+dkCtPLl9p0HpdyT9XYyYL2yncBWgFHg8htQVQyu7zvWNMrohmXD46d
sTgOXKH1lmBLG1aYuE+Z2SkMm7eLrilcDsRndqUzFsFB38snAMgyXkjC8mOI39YkmG95llmX7cSc
TLzEJCntyV9Z1N1E4HAV6CNk9m2SO1zW3iGxbTZEmVpq+/kl3wcJxwz/Z7D8kq52htlcEaIUpZof
TWfubS0blOMo1GKhyJ5T33Zd8e4MTXgsfUjc16l7V1Ewo3txlGe45L8FOg+bMSHEiCPDdRWJE8t+
AAWlI57KQXwlP/kBipQfcx3KBxYof5HX7iTwYRt7fFiGmjspY0Cy1myNJUePk+XADODIe41QN+g9
7pFsWuv+whEm9otU1USrCgDylJOAHx5mhz/ogkrOWg0LKHQc/QPsVQiH4opAcJU21dxoZOB3IMNi
WX5TXFPgbY4IZ5EAm+W8Mbm3FCO7wZhNDL4TGWsZ19scKQXffkicNZ7Pm/dDx94wJ7K7hK/iaUHd
2O1QDVxiAGnRIRx8yX8qVxFrMrDtTW4lp7VX1nBJcvij+/UZmMynUzZl2hzf8criEMAes+gOQOv3
9bjkAhm9E7D56ng40fVKkSf+iJaAsYyn0KB4EOv+q5FVla1wWxR96JMeffGbhU9mrHqoXXoyfEx9
Czxizd48s55uxQDZRieOs33TDfGFzsZlztDegaB3Nr16oKkC/NHWWIuDMLx3eF7bR/zW5Ye7vbZ7
sDko4HcokfmHuKLIVnhPVhIhbyL9hqcQpZovUqu+dxw1Ck5j7r2EMqKVJ3TgmGloXD8zq78baqgh
mDYz/2fhzbDWuXMLylnZVBng8LtFSYLsLsBnc+n/JafcS03EqiWP/X25Pvz2+PB6zPHJ1BN4aRtc
36xpFmDkM0Q24xUEoX5EBpoQanWCkKdU16F9gh9JGi3n0TrI1+LfYJFAKyTYI09YCheACbP6Lbmz
+Kd656uB2A+6Nf0qab75nW7XsYEOPO5oJQ7IOrSVzgQd6D/XUwXURVCdoScYarHX7zHDYznwYd6q
TZxXOkwn4fxyMzaWoJ0n1Slf2WuMSbbJdao3w41nvA31SaFItNIP1CcTX1rrXzvqGb3Fw5uUVwXD
KT+uhyR2xjvTXgJp93FiuXe/vX5PG1zK8Za+XxCujiVtZctfBYWTb3cOd+60iJ3TSoy54qmfgjjX
0Yt7ANgdK9crz1nGu/MHC5CTEwjmAqUREhR/r8+ry13xeqWntiOy0RE5QodA03Kq9gkC/k9mPpav
p+BYE5ICwg6KQ0Fyv1QJaGCm0uesyKDXV5kpjoxRrDx0WCHmBAC0eQKU5+zJwfMVKAruDCLbGj2M
SXqkZzwKrwWzqckVz6Af6TMHpNjduuoSSImUh1GiqxquWEhmNdpTO2RkEdURFbZvaNVaH3m0pVwR
YpBkg/Klbr6kOF90EmZyplIs+kEXSlkVq+o58G1fAGRbWFHHT1KurVNZCj7KV0uHodHtg5h8ruUi
9fg57/5P+F2FY1gvosaSWwnKvSsW3BB6BR7pJPWdCKgiS+AciyZfd+nK1zxm8Q4WvoKsk1xo13cY
a+D/aLvvN2RTYfz4URab51zL0N8hXqXBK5tLnNDK02MB48q4cLjofgHqEh/ygIY9/dcm6kdLM1+x
lYKOs4lue4cCKkLvVWlpVfTKEAfMOeDTfU4jT0VnHVLmN3V+b4SEwZicVuSsiWaMv2+6IPVZHfeT
wTaBuxhf9iWBAZFyaa9bJS45hYiWQOiE6XxcUzbJ63hB/RjizFY8aT7dF8rL+1X6FXb+hMAyVFpX
DQpfkDHCUPRhsidAEYjuhRyYSW7oXz31xaYVgtkvTupXzxOTUbIDgWksSOM0noTK/aRQw30f/PL5
fKcpglfkzab7LYamfWnkhWEUtABWSG+sznNkmILXQWVDpmExQFa+xHaIKPujnB3FGqmFjsYo+gHw
ple6LzMX30AMJcorEIS+aSjHPgJG08jT3PEEpj9JplzlpbnVDNe8F2PSuo5c+Bkc6fNXAEA5G8T1
iMp2vrSs6MZb+r8HBgtLijkg/kclRc/Z88sEhaGKbpHEjEaowlafUQUWJei7wt51+w7tbGMPscI4
cIK0sb8Rj95Vqvq91GryhXVODtAdrIebEOPTgwCMZVqeHdmmFbM67esvqTn7LGiFf2w4YJfS4eEE
OzQwvEPg0fqmhNm8WPhYHtpTIiYURvI5N1E3TT+oEss7DRd9aNnih83OG/LJh/A2tyvfRfgrXkcJ
ffrGpk0vNgqmAB0DhEUZSxEa3R5XIM04gwUxVVyy91w1rZBX1N1LtNDzUnzxjojXmbGGkUh5NNlG
gJ2tS0BDvmekPaId8vAP/q8NvCPpOC/uQ40m92zvHHfrsL+wLiqS8EUZEUvJH/7oa9PJ9QR/LC8w
DMe6L7UTB2cr8QLOW8FT4LmUKz7LfJLjw7g3JSL5jr7jrElbtL1cXRryp5BFCtSSVxodYebk2bZc
oZmXZKa1p2Zs4O3TxwiiHfEIf9cB1MTMfiiF0c+JUlTVLhiIrR0sdBSYVlx86isQZa6SRoEFWfrz
eI+cIeArcRV7LV/jCY+5sm5ck/H8VScgBDSf3VSJ8tumYLq+me4xqK+7r+nbkTXxi+sx+ixpZutE
MWluW/QMymihj4/y/vQ7WvoVqQ0O2gAMbZ75DnET2QLYdBuNNlt0wOcAAfjUlDJlYW3Ie0IUVN4s
L3QlPQTAFr3sshjqEgfec0H1AiH3Xmz+jK/zQcD5SMkBxYf/YorITYSLDCDYfG4DOFw7tPqdxycc
1dEW9YP07XeoE8vsS6Q/Td2Hi2Wv9AVSX/I/RtdSAeVtY8E4xzGuJ/194iBEv34m8ar/+cwmTEYf
Nc0eZ7tGJ1DXlaPuEHU/Ob661MlChqMGh/4uhqyL06oj26GQ4lfFUX8V1Dvg+tVZRXMkPIls/ThG
dA+iqEfn6a/s22bDZB+Thkme7RWf13OsIBYGeZvuJI5UVmjEsW1cxOU4jnme3mX2pmeOvWBuIsrX
UdTSqSxzGjypr99aZfmAR9YzJyhO+63PXM9BF747+tiCHNLHv0vTGen9EY9Jx+zOXIWiDLGOukS/
3pYOrQZqhxhcGTQgXOxh0zIijP4p1kCOPSJ2bA9bIQ3mNb+1zmwe/dgE/wS/CHsWJRfT3huJlxPh
nzRwWZ8Tl02XBjhIFwAlEwLSfZUnFRDsBcP6unAuh3TwJgYfzow0WTwJqn3M8GCt94hKMOTNdAP+
ZTFVTltVp0s1CN96zHzUpRUnfEChBNvnSqhqwJX1QHHsAnCO/9sMVvMk16Utu48h2jOg9FjmU8Y2
BT7c+f3cLByPcFwNQBEam1rmNsaqUYbydt6ar/EwD8t3Hdz7eIT5Y1HpixFyAZS/gP+75JVr3XFb
/GitF9w/yMpqr6SuXZU1ssAVi4K+AwUR0SihFX3RPmq3btl6o03H1V49c7FaLD7chFr317Nb3QZF
sJ4ed88WqLSV8GvmhDt/yyCLa2S84ZFodQwan7XUFvJTlbQfBsRguyGXRxx1W9EussaZpiHywKbf
UbOJ+lwlAOVB0WiyML/EUhFAZ1MWO3mBVU7Os2qe+sGzkPvY6VQ6UU87NqXFdxRmRoYVc7Dfy2mi
9fkCg+/uGNPigS/DL2WDNtDyiwij0XcrmA78TG4UGJuStX7qw2GICE8B+xl0vV6Qy7O8osG1CAvU
AXZYBqlVqHliDgg/1SzeVHtzrqIrpAZk3WZILgsLAnJqNZFvRGcjEP68wvfpPQBzV4TlzZe1v2Lt
RpwRtkLn31OzT+E89cPWDRksMmLOHwZX7Itb2iug+vnWDQQ/4oxaAwRnpje8W17pzkQ5SGXicw9a
sTsjHNAPtAvnsGmI5nzZeVtDAy3leDSxcK9Hsk2mxmF+ppQbhyjLPZzcXt2ZhbqAGXQYVvOBG8Ka
YI0W5KTdX5AIJNl7QlrM2etz6GWruH8kbe67lLjdAd88eYtGCSH3QOSBt+l7+8IF1wneYYrnA9qK
VM0qhg1Vdq6DJEUnt80Tf2dyrm2IQEgxbWstURyoOndSv8tew56eo8FlJVhVLwej9Z7z3eSHukIq
ujbABoPof+23uzqCO47SoHb2PWHVJiL8HgysjlHPP3FFJP2C5lPgX0x8QH75ebrH+hx9QeJVdF68
TktItJFuVyYSGtP2KKevAugf7XvJAa4rKCcdKugSUk0XnBMxn17pqWyUe053OL3jscav7FqiicXp
KTCTMc1CE+htfn8sQtYQyEYoh/+XpDzU+nJ/mvix3PCRF1eGPG0TvAReki6GYUVlXsP0EI8WXITY
dVPlxsThg6wJhIMSnaWVNN4S4ILAEpcltETJNJUyIvEiBI4CUfcmgwVChQjaByuQ+epOfodyKVf3
1xrVuKkS5lFI857O2mFVRvFNHgDecgPmjKZ5urmDdRE41kYhFKvV4avgZ1pEECfhJWYOw+Mu8Wh8
mQFNyEyGgPJDgWNAP3jzi949uwvt4E5r02FT8kaubhG/A182TAtjyC52iHVJ+fxq4S76wiPwEkno
tIsT/YPWxeH82QEpaT9Cxj9qVnBnfcdteRzjiP2DU3zkx1GHv0l9/9mAIAfEMA++UweXzhGVYUmL
7XNHIha4Pz5xIXL5ckVs0A0jaEFn1qcZVuTQvBOaIOdImwxV9AJxiK35GBp0bky/YAqDWmzy82mf
nSYxMby8ZZPHT1MHpictP01u+e9GmGnAlgI2hYYaAliQ5u9v8bTQdERV0NQ21IyQz6OGC3y4n6yc
GCVPsPGVpmYYEhNRkmlA+dIfM9MQ3PDZaIeu/ml3QQF92zUj3UpWhSHxaN2wBHYD/zLCe1ULJRLN
kiYBJfv2DDF6UGPf6nWVCiSRPUVsO9kD+DYy8c1PrKFFfDgrSEuGJiBntP1f47m15JMADKZSyetI
kfeHvg5B7aNhu+UHI1ub5lfCflfurND+8Ffu9J7/hx76Qf08wS1aOZXsvKYxnzl7/oZQE5MOWMpE
32yhrE5K2c734Zxo2IT/+xN5jMW+zgahBqw3AChJV/Uh3D6/PaQemzam5ddoMsCtq0/DrfMmdRk6
Y1Lh027n0Ws+Xw/r4z96kAd4v9a39PDm8CdwbsNl1d1kTYrIo/PkcL+FTT5qYHlqU+kPpth9lDoM
OX3yvXMg3NxtpAmnmPYMRYAFD+kIt91m9mx3eZ8t/e+3D/p3gPzDsy+qfbckt5Ct6kkC9U3iFNwI
uYKqUAbEnpa+vRXdVd9S0/Xvz1/GIbVTamHTNyofeQoZ4twMuukF7Y6ozdjecT4sO3kfb5IZCLb1
WS9zBqlIu7qVFGWwrBEoOWpkty5kCSAYCU9E4eqSVS0q8d6kOfKisCAYQekWo5Jxc2k2L5nTbfeY
VP9Ns48WBH9ulyOjnY/8SBJcOndRjXCGSAvVAxVmyF/PacJXCjjOPRilJADYBG8YNdKEXA61W1Qv
aeTDknKynzVSeUfXUU7tfws8SlgvygXjdCG3L0sJxQGAGQ2XotfcABjIlqSx8nwtH5TXX7smVMDH
nC7W0cbUdjPayyax0Dyif63gy7MGiV9oRlSoJbh49s0SSWdxiUXFEoO7Kr0pHE/CLAIbLpo6bvqF
TK7TvaVLWGXCjHvhVsC9DD69/KmpQeqwqVg6kLu0RzEMLdng9iD/giT+zYWASFrJTokkkTiA7wDN
6sWpFbMJAdU32RYERbM+dfmV1nOj7hT2Jb+G9kkLeyad6wMCit8sqWWp5isVYk5G851SeVch0gtT
y5WbSh1Y3t2TdDUWUKfHgHlxRLbg4R8qx1kyXs/uFI9bZzz3kMPP/NJKswnsHIAowhHXeFVmVFKC
7nGDIUio1eJEfqqxHpIZkZOzlWmfnymblY/2oH/F2WFtE4jQXjBUoFK/3OEZe4nFW0GjXz2BTsjQ
Y2ZftR35GaPOLxOE9ppxwgNGVU5qvYGK0TADJKBW4YkBHI3+fHA/186tkn0Jcqj3PF86Cv1vYE5H
DdRWM+Ue6NeGf4QatBe9oz5Ww6YVsGpTr1pbo4M01Pf6sEhqzF1fQ12o/O32ybUejWP91ZED1pCr
ttMI6TGKmMRLMYWTfhDsy8sIPKGHc5ckablEyHfooKU2fIOcGtKWC7lHrL6uy06TQju8gDJK9osi
SBVVHUzEpYYqEneVx6J7MaXVh+YFiYO+T7MOtHsIxFCpaDmj4JPr/9mX1vL4Evp5Dvo0ufACG2AS
3GMFqslXGjG+aTTeyUS61fwQJZ4z2GUZ3N2Mx4gpK3iRa2LBl3nxhG2AL1hluW72OWUJengEUGLW
BnY7LBnAOyCGZkatv3cxRReyL4SFskX8HmnOuE3WVp/sceq1FWAj4g9DchM5cYlTQAaZSh0/C3QH
Ej9nIeMgDdBeR5XYVfdj7vT2RGnKNWsi3evaD8cJEgtLZ5k2CmjcSSgHdE4ptUmMeHabJlU4G7Q+
mHF6DhVVo11FkbxalH8/MokqVNZbPs+SnWKcqHOcOcYfgLTObOkotrtpA5eXvfz/5gz3SCadNci0
xjy73JYb6qw+xKiZaX28SBL17euUhQjPXzclJusw4ik24UJ/72OPaVvG979nU6aZoZxPur6ITMVY
vtts2/PVsn7ouYMmY3LHz/WitU7jHE4Ob+WVJ3RaGns3mQH5jTxUDpzzUF35ZQtLJHMMsLSGSnQw
76mHQEqR2wnSg7uWp8Tbo9rQBmXCiPc8aCOFqaGcImqZHqRztMdX8fXz6IWLz2XQlyC0Cam25lsc
AJZoShmHhZkZGo1tSlLlmnVLYY0nnjQr7DTwmZ96ClTiSDTDB/ZxpOpDLG21BSXxINGpjaflYUhd
QwxcqWQvJ555QSIaAfkOwEBSSXXoXkfYDXqdKV538X0HHCHj6XGc4ymjFNBYRVpEj8oF6imDZ1PP
EZYh4uJd997I44o+PB0O+nJSE+e7xOm1j2ljlhypKKnXjzXfIiXQBJTowdQqi7a0wy81+cH70hkf
Jgw3Dh4eNUidVUVXaFsPdFBymXxGs2WXfEfgApk62uAadHOVcs9kx9EKLtLw2EUwoa88z814Q3Ah
eGw8dVX1TrvHHM1E07AWTRvfojLielulKQrpKfZT3y46OgLcmzo7gVW3QFVgfe7JkuThWLzBWbwA
o7NJLYRmtK9W8ZLUGG+teC1D0uqDgVkZCep+phlnGpsDvoCTX7yn15tO7elArIoxbiJ0s5KAikGH
txqMuoIBntMRdwWWOWVAJjx1RIobOK82kfCooPENN9M2DtZCJyzo+vYPQXQRtKyh/J40NR4sIB1h
JTGwWNwilhevGTDCQskAY2oVld56x35U70kfbbUGPpkDZkPVCIfOnHpQgO1eyjQc26SRoKGlCghs
wJsL3Fmy9E2NmlfFXOFFXCCTHis5tKm8DyL/UVZOHugdxaaQD/D1ItRuwBwlp6RBxLySX0rcOm/t
k+HHWeeQ7g74l9TsJsop9RYthXQFy8SdbH4Ki5VI2zQOaE/dAN3ZFfwxuvD3qrvWaZuJOh7XZUwu
ecoda6hagLCrkIAROwaGiQfcfrSrIAF2tsvkwNCP6QdQc+4lGv7v6rdUpBGmz/F5RSKiyTZvOzG5
HQoirSHQzMs4a2W8eCOGagdxxoOnTMCUPOczSDj8eQ3GnoRI29BxBWNcQlyQ33UzhekhkhNM+7hH
h8tIUjLgbFagE+urOrHgu403dI4Rn7f5Tfal2OeA1N5CTHw2LWgq9bbJLfGrQmZ3jFNshLwe0f+p
Bg2/of+hWi1LdCdnCQj/ZrkE6aDKLfCVxXmHkB08eyAsU/UY2b7WoP/NLwkMBnN33kJPwyrjD0aY
mElo90hBQ1G1fdP7u2JbYoRrTm59txojN6Amdv9gV28K/KLMRJu7zLpASkj87/0L2yPG7Xs0BUqc
EZs0+U0fNF+w3feAgRoAagvgdSYP4hiBIJiqPVuKA8Ujp1R5wyp0OggJdH14I29SJNd5B3RwUrqg
NylOwrxB+WfelBvjtR2i3qz7E81pNiN9dsj4oRi7ErgYXEAA9IuUmsAwXdkukum4leQUehuCRPsF
+PnTzfEdNsmRnau3reLDso+b8YLKWTA0JEZbAHrhcGehtrhb0U6rGuQJgfLux4YiCdkk228wG46f
hKemPeAWjBTPfIp1BuVc2Uy4OpwgRIlKHPNQ8MenV1/ewu4un0U7oLNuWMgpu4ww0f/06IWMxuBg
Lv84SxhKBP7sQ68nhzu2/BW/xtx5Er0arf4ZEJplkPx1TjGtMEflWR3Ft5PA7Cs9rTmf42Gmgz5o
0wpmcKi7Sw0lmB56a4wjqDSxLHWwpvcunvRwYxfPG2KpRqUmu6E72h1idjP09VIInXtvL1hWSnf7
mArvaJwNILVxMeOaREj3Tq4SHmNItC7VG6/awpFxqLhq559+YrqCqh5lX1bfuoCGWLrZBTaGo3m7
9fU3X66P7YKjt1tCVrrdPEFpqbC1E9CUQ3/a7eMoC8UHtTzQ/UA/QR3xjYq/ZPaPi8xQ35C0xx0Z
KqYdwnPtyuTv+UD58mAbo4C6tK0HK3+OkPl3G0VEnIr+FF3/pV444ljTag6e3UY5IfC9fagFAoED
M4IImFrM4IWys8C3SGyaHm2pCQv5X7bto0t7eN1ijAPGZalBCQokJ0FSXNIr/zJbLH4vCKGXygJG
9W5tP0BOxSPA6nZEE1LzTXWPDXrn6iFeDdXZu7CvvLKMik0PZZgG/cLQpjICWiJE39VlfY0jaJDw
syjrY8KZUNH6jqCYfMXORnjlrd10NrUyWxnTYZ1syo80Q5kAoI+G7t+FE+te+cxmPIbknuvrzrMs
vtS6AsxaZx+vHo6nmAHxOvA2S9ECA3HFsL5/IXFEnveEbQmX+9aWPiRJ1Z0OYsWYF81S36ubtvVD
xzE0GBpusMwSUt443QE4Zdexg+/gyfFWzOxgXrnr+4dS5ZWlVpfMQVS72D7omAgBG0O9DWTQpt+X
8y4NTXLeIWoQ4EZnHkVdyIeZI3QHuRaGOskelIjMWnTMU//uD3++waR0epIvTBnqt9szhhLn9Ah1
0ZMO9xQ8tCMAwhU2QOy8Hx0SjtPdSkmOc1H+UX3JDYT8E/ETEvpvmFPhjjiyc0NMvzC655jWryFZ
1WbvmymZYw6Gto5O7CLLWp//2wYM1JxJzWrI+Rwyj37/J+OXpskRAxertpYecWdIgYGZ4BC92HY9
PQTMuOSAA3rKKV5SWdCQZjBnUPpEULcSeF1A8e0bPlUYs0PoZLxPMaC35ETNvue+Kmiusno1/EdN
GgBAMKk9uikhmoNMDFwtEUnwLgsUyJeKmGpz3DoNzqgIaVNaRMrG+NM6foNVrwUo+x+e6JgErqWc
moEkaThfGL6qcJAXftTSkXZotLteojfrU4bhg2hyK9IDPRQFe+DlvRhTHHfsudIjM9lyQa555756
vK0lkPzrTI/C+7Z2L+sr9uDE01RAIJVqhaE6DA0tc0bpUsH0h3ZuIuF9UTDXMLZfqA5aKqm41UTz
EfjL90X1wKlXGMhcc+RaXIHqYTraIgSjqhwQvw6x+OkpuzljzCx9elwYow3zomHrwJNXi+b/ERsj
mZNupTU62AXj7fn+6e51+ISPUdbPUsTJdMQQk4QSnJaXQtXNrSr51IKfcgg89KcoTY9r9RtljRR/
vv5wSVQ+hQUVYPKib2AdoKrM4DUb6ndI+x7Lt5nSkw2+kiN8IKoEs0Vvj0HpV8NU4aLlYVHMkbz/
LNG07xuB0NjMT2D69ZrhQczE+iV5vDRCDs0cLO/TsJqRtDrvc/BBHjGd7FOoQ0tGWXjXdGe2EvqE
ZzXlnvv1XshDQDcKpPNB7fyusXfeELQLeIp/RxkVsyPHlJUwykJV/9NDaWiYblVIXcL85/7yMGXy
0+zU9TRQuuQGYpazpiaP5Mh4Ky9UhUTkSWBcaL+z0MhexqMYZB6t95lxWuBgop4NqhqxAhU0OIT9
/pZt9lN4Vbornap6OGVme+/Z2MfNmPtp/VrLIMifB7csN1+qd5g0zWliOF5ss5Q55gKzwHLWTm3w
Lq+I+kf/tFl+ylZEiKq4PEOyl4vn0uoU72JG4HqsQ56v602ZiTR7S7gPByXl/f9wmAFABho9KO4B
4vJxeZtdAZfajqb9u7FJ3rOoAplRQGI7DpazoORjXVDoya9Mo4OuWrvsc70amOleD7S4cABzyYHE
vC22Yg56x4oy+xRlA/S7XIch/MmGLdnJwGm8W0En2FWN/dR8WmvXRq2bDn/imLBPKTaSfiIprVbH
16bMH8Y6LzCJwj4Pdgw8H2PqiPBO2lkF/cYPtivuDLvRi/Tgp16pYQmEud2nMb/ichrhvh+R6IoO
5hyz4WCdUlQshneSn1DK1MiwKvO+Gv8UKC5MCeuLq6k/Tcxh5zjkapmQGUuF7I3XB57SQlbqcRtz
pWd9v6AUKyxtE9V/bG3sZb7SIhYNXaGWSn5Ao8q7QvpKWpOa3ChRsf3QHemW3ZYlnHUjYaBfhaMh
rMUcE5BbbO0JcyO/muMmq31jQdjz0VtouM+lBtN4N+Ruh9uKT8kRYjPn0Duard3VD+w+93XeZtb2
PuZWaOrLomqPxV0M+iTJnHqlKHxEoMLihFfEGAR9sJMWLc1U2gx//fdGhDKKH3xBv9pKZPG5gXLi
Kw54XQtz+YEbXICLwfba3H6eWqPieTZGXWj8+31IzeskVVlsKIiWKoDHuZCX36UnlDfrmPo2fC9k
1B//SDbF938vjM7zY9z+/8Oj3nmKpJdBbhsABzxIyKu1/HVOxYogE5EtvGMYkLIGtuJaE1C8bcnY
DA3gK/FF1C+CGW2k167Goy1Y8xtGuPVN9jVVs/zAz5XhtoHpi1I+nmWRBsSvHgyR56XdqIAuCL5r
pwgEKkOG1nZh3FWzbwcD4AV7gTTje5M6NP4vkW3KRcixkX43A8LcxMW0MZC8J4tNA6Ps7tMof8GO
1zblGWVRjauEQVsq8tnUogIrqhviO+LS9gO0QtJPVFbUZAb5+0T3msB9iMoZ8XxBWWTIlR39/xjl
rXzKt65ux/AAJkU4vlm0Ow6jl78iL+rUt4CFrprBzhYmsFnj/fKfVH3sYHi6qcAtom7uYjtMWloV
PpUL3Lg27CCs+INmxsYi9mif9U2TYmgSjexiEfWFmLqtF+vCYjMo877jjLJuNPJnjK14nwdxFlAz
BI+kKQ8V9OFHP4LTTKZckMBiq83f+GQGFXKP6X4iuKuok/0p8asXRU1OCev5tNH0ygJh3Aj5CywC
KRoBoTt1IZ7AMhHGm8DVjSnLgLxJQBbF4txjQsJDDhWlz/M0O3SKB0arpqADfBOsomgqG0DxaiEf
L82hsdop9hGBu+rk+B5Gwpa1xTa01Kq8LWtp/czBXu5bqphLECIdrvNh4DDUJNhLW2cw4vQlBlcV
KWH5P3RGuJMCR1BAq8wi/2XIUligZKrnpQIh32t0QcLtNtyWvcEXIaFuYRqDPCM+XIVJY4evOWma
/4Gg80oI+rgg31UxAmmlbV3eNeaQDxfZpqIDEPDS8clAiQAuzL3clTnXZFKnIs92W0hftrSg3Stl
SZXj4NRa0HvJkD9Uev/hJJRTxLvl92ZxUJeXwbDRkgb/xdPiae8R9LqC0a9cYVvkjmpMGv9DvpG4
XYY45uO0Apk3tEMuS/zPaM/Q0gRXc+ghP5W26Bt0vCvzbl5PddI/c87bvXqms7ypNUWf5N12KWlJ
BA+DUm3gU/6N7YXXk9TGYZIBQV8fNJZPzzcqS3FoqJTqxA/Iotxdj/HGb6Qxb2Bm/yj/C/f7Gpek
SG52GIAPFfGf+L8hyfEjIeE9nYNK9OMjdLqLDZvRrMtUILxHXVXXwPYznRqImvkDy24D6Qvo2zMV
KbMB53uab9LB9p9xMQVdQ/3hKPvmmYCmjjySBHJ3Fv++cly/eQ5jPw4MwRSFtrmXokmUPUFu0HCJ
q34NH6zuzr2AQ/GABocFnQqds+J1Gh6bxdH7z/PacZvrK49uNB1MoPVlOdyk1EiU5gG6vDKvDB7J
Z5vAPPI6BoC6VQVrzlYQAACn3v3Me4q9pjD2tv42/ULJFLX+5IexHxTojrjPB19rA5LAegEXRv79
aJYma7g0onyAUdVlZ4XUPtj6WY0MW2BdcSd/elR/eOXjne3KNZYze3VRn8zliNXNMHyKAaVyRPJp
bPTZfbGK0B4P/62qzfbA8V6lcIiUpTzZjQt1ghdr9xDPmczRps1qfGLQGPocgvMG5PiTY/MkU+KP
OT6YPE8mtMt8adY0s645mO/skLcXraSAG4BbhQsNYlrsE8S/IypywKNVXT27lqQLkTLBWuIpbTE+
61lgNwajFaYR2y5y8oIutJTZwteBSqaC1NAJpQfvoxw3lCz2/aNuVTJiec8WdtVu2NinFnEUgzJt
V+SHzipqs7Exef4MRNhaPW/i65fusB5o/3ATUvGjYhBr6N0k2vYEwdBVp39ZTPyhOkpVo6znDqi2
I+7VvizzSWJ+ZhexguR25irmkrXKbdt7dQjsUiy4zlOqgg4mrmdBxS6gnqlwInqm33g8Gej89Dm4
oW5Pu71pjjRDOYnsPqA3CckpB1PVgp4wFM9QSwobG7SeYeSoX2YX6REj5L9IcS7/j0Xx4MuNs2JW
1n1sYO+Az4cP5nreXkFdUP5hlTBytd2e1MezzBPzqOJBbhfj+OwrYoyXNw/8gnPT+s2/AkbBbq89
PeEwvjkB36GFyI9GxTAAELoxH5jhgqmHLuGQ23fDY0TIhGTy6PIi9wnOZIKKIP6pGcmB41V9mBBd
zs5q3W1CY66xG/FZeDm3NhgVFjLgvZTX9+IV6anVI9S6zoFsLz94avM5FsYNAuo4dIgcYr15DgCJ
u2X8P599iJA1y8WU2uhcbEjCeHWtllv5v4SymlYCLjoRqF7e83JGHNWnbASsRFUUOF/Lte4UeLz4
iywncETuu+iZ0LfdiRtZ8jp6EpwThQyingErxkdpgRREVgPrCQQmGE7zLebhsdOmyQlzi4GQeWjy
8j7Z/wWKS5r8J0nnUWbkVaSmmJzEQvMJ/HqL6DC1H4pJDmZyt2rdhQH6x3u1rKztexMSfwHgm5Tb
6p5e4P1B2zhC9Luh26T2zyUR7KTWEsJQMAO+zBleknVnauHjQArOnPo+Z7T8RWU/P4+rDvkyhUwa
cXncDlQwYLLIRGwx03YUqcnTUq/pbtkW+XpodywdDpx6zmI6UXHKZIud6yEDwruT9bPetMW3lLun
aZSyb/k7ZJpXlUJrf3iV22DDg+vTJxl7fdxTFxpQPLy54qA4JcqQMRFsk1SeQ4YqNh/1T5pyQIqg
P95ljWZLGfSpJtFFXdLToMeUf4KWRYYynoybzZMuerhY/tPVmXvwPkiEu/uT2H79nRLEqy/VCU/+
4w7mVKaZ8n/GSdMtr7xIPwKj6cEwLgR2cshVIM0zZWheCPW73/pML2Q4Dcpb8RLs1nvUi4QIKELZ
lpuVoochaT7eq1PEXk4fml5pSnDFCxOEmpJM3aq83UipDLXpguUE/OK/uNtBrFE6kDFnLFTjOwi9
VBZDH76qGa6RgQEDliuneGB/9gBEbkDEYC/Pti3XBmdxirQdaSsVQZVe9sSblz+yVhSQ5Sr7+jsC
ynL01dtTr+LEc9KxtyIF1TJDTO0LoD+h0rMezqbErkfLmz9mv4tyLFt0itXgUpdrBUEvyMy4n7FI
S/Fu5tXkMXRX8L+lfQ1N1G0Auhr5Snvvo+47+Mzi0H2NZLgWPbHIN9VLtoxfYMLKDttXjy6eQKh0
AsL3+/nBWhS1i8ZlbjldfYiIdSSwHA4OcEMgiKHOaOS+4LixrKme+GW5xbMyJ4yTFV4tbCs2KLnW
/amN866yCD7VurVKRLPWvbafLW0gL5+WrR+r5rAJwJEC1VxNkQJbLOzPt+4vC3oeYiMbiymwKYD2
rYxOAch0GU85cX5uxdljllKD9T6ASHTosfg1939Ph46wNdfFb9c8a56BLCucByS65yV1bKca7TiN
aG3qY7j7pi8b66yFAP98iqAMfFTEU6V5jp2x5yPBCm3zD+gA3NmGc9I16riY4gBr89ghM9kURksj
citf2+TqAh8zOhLKr1H9j0lGCenvVepDcrP1va0OuMWXg41lvbcWXGh0xZQRaf95kxHrU9Hsz52Y
J7TNaDjdoyCRMAdkGQYZwkuJavnTU0DKmEaGqaV1g+ymkiZGSLT9NLDi24owIWW1li7+uu0az1Gp
W9i5WZtZVBM/Gc7HBOhbaY7agvy3P08rZ15EpR2RgG2XCjyblUPzP9FF8HfIXs9EO1CnDUaK/U/W
WLQ1Ym19if8UNLh/bG6jRqD4awWDUVHUWtBrUVFjXCHNoQsJZDjjclmnIglqC88a0CrZ/wsh80cZ
GoEfyDjw7LOZZiwAIzBCPZ/To5Bqbw0zgu/TArfGlotdrDIvu44sWiVDb+XdJLdRexpMMWllXjQt
86HExFOkrvhmvcOiIsBNiyFy8VeOcFGPE4dOo100KKXUnPdOYU2Fl1S9W4rrdR6gUfxX0x5URJ8l
yiobthc6aiaGUjFRTr39k7VPOTKa1utKiBUM4KtjniBUM9DCTliiHdKeboZAduXZhJugvQ3DZ7/l
EHKP92VRjWvbl+NEg8EdEqvgDjA1iCDTYXYn9zFo9lUJXig8iPB8568M3nyqt8UkoF1gqJ/MvgCW
IjMLOQ/DMh/HYjtaDswOadt5HE9zOkeP0Hz7pM9hoz06yX9e0N2qsqwkzFscSMCIWWfe7CVtl+Ak
mlG9vShUbksm03I5CQWpvD+VISx9e6M4Z6UOwiaguG31BTzRMp5KFZs0DHO8RccW11afn3/gDIKe
dUs9EO1hWAPbxrUgHfbrzs05Hn0rqzRYApOgrfBi02LheSxV2y4Jp+rkyZXIBZn2axCovk+ZYFTN
ZdMfubwmD9AacZ5ByewukuZ+BS0eu710nUuo1lqd0lhEVe1z++Y4A6urfFB9UAmhKAVgs1/a5YCr
kah7YsbYVnnEFu7tnl1GTA8SDkLnCGqdE1DU56OdgGJd4VlsN4HeWxQh65ZE9TJXFfSNOfOJ5OAI
SCREtLjhgT2wg0PvK9wT/lkKnSRETA2XilzeyUewTRY5HIVxcIwJsNwHZjRACrI8FmGw9R4fhWaR
DzrgSNDMBb2GdX8ao8OTJnobCo8dNp7mmw24mLAKcbZlU4tuAdR7HIckxMOv2I7hzCf82O85kJ59
b8lGWg4LfccuzU0pA+tMJQ91a0/NKBApULoVPKc7YCV/ymkG669owKi8Jv4IxwWHZgSbYdxC+pD+
J1Nm88mjL6GxBPBWnihx67nzGJhNSUkDmB1McqaP+lySo7zh8GX/he5tnrHGeo22onFp6KJkd6L0
jsMk8mE38CP2Tiw4qPcSXalT/hF0yrH0Gqhh1FQfws19K9nDIzw6nXB2j5iFynj/CO8O+lXbDlk/
HiUhe1sLqrNuVhAC+yrhpJ3f4YSiQ3EPQ+DlE6Q5Xy47z2jFxoIUWQ8fjpORWhfwlUeif2eKYVrD
FihTTRerx9xeiBXllSuVS+H1ZaL9I5zGtTlETXKmI8qFWdAPsaxa5iQC9p6PCvs4+X9ZgD53MTSd
Pva8id5B36p5aQu6e3HJs53X3j0dvpUgcSSKXsRGhu74mlaAQy1YYhIeHS2eGGHREqdOnHGENHVa
skdIRdExjVyQagphZ+Gp/fUgmbsUCAnoFJFt4982z+CcMAPmEeLaH9k4vT3CXnWSwhpDMtH4A48a
CpzVRuEDCQyLytktALIebuYIyFGNoOk5yBJkTM7uYLb/Ri8XKie6gtsXmYiY/AOsXcFChkcUxTS3
Tke2megqvLsAwQX4qbhGISaw0Ay9DoVD8lgiAKw88Cx8mTvRDYEsoOTSUiSaq+MIkcJYbF7Ce/fX
EQ67xQkiLpWL42rWaPq64gPdsoLfo/5cEORDdUO6FwD04tnmNwb3akDZ+mbbOD7fwUsUuasTPDY0
WUyFEq+aB1uPzkK6AYJemct8Er3MLrgrTMXhv25tk/VzMLJC6KjerORpv4rPAt7riJFJTusmApu7
sNKLsvHh5p2RY0vcp+ft4naLkMDWFzCg2YHzSo+0IN+AzD39Beada2ARoxCEw++uc7DkDObsLA1K
FYu7QnsQ77ATbzzAQQ08MMBB36deLbDb6JdT3rIUoI+2SriSz9J1QF7B3KVIuVyBf4CxAPwt6HP6
zA0kIE77/LBFI4UpDbAVBWaQg7aQLCaQP8u+80mvEBs1fE8em2K14QK+CpEoUGtMb2WGZBtf+vVa
gJN4EHjhypsgFe4V2rfIubA+ylUqA6nba+7HlZSjO4VBNwnX6sN04NmwLDxbu1Qu/+zS1pg4DZfI
vDksrvvtEKWE9ndM569+R74NmIZOgIpf8lSJe/SZqzdLBTC0Qhw95ixUn7Xfr3PdSolDy2R6Cc77
mrJ2Vzk3UEwKS0r28yF4KFREw2nAj/uheOEXF9vVdqHBa+UG7DpkP7+IXX57nr1AK/cnTClvq+k0
CfdNVkvXeS/ZAmydZXSnlfbdKaEhSzQEiGIsWmLW/+OF2OThbVFj+L9k66shnuTBX4gOevDbhd80
L1opq5mqbyGXquC9Cj70YjdPkHRaeDYGv/akx8O7q5yRSTAiCl36Xm5yPFZL3EcbP3e9edvK8f6I
JFqlR214rrfjoI44t5gaQPqF6QqtHikdlB9wYkDygxQ5S/PbvFWjtnEoqXO34s8n83RPd283MA80
QRXUiE8yBCK8Gtc2hvLwiI9BoqQG/OlE7BEz4DuS+WriNHpNRPLkXchB0Y1D52NEnDyUwtXZDy5h
HOoIl6q4Q5eJOee//f3LNZkQhSRw4jmbiZi+TlzCb7NgKeE5SvJQtw09oKhi3B/9KynLWanreRvx
lkHUS0RpWMNMjnkgzkZgs/leL0Z1HOq4fsBEyL56IbIKzUsYDnqJd55Kogmf9D29PWw6guQf6TIt
SKaN6qwJmDmXkvtxzYXpMoFwXYXMyH7p8nCLx5kgDN6xfohVjBS5rAKLLE8Erw0OvfbOHqwY3pnB
2X+82G2za6a3JXbi3H9Oi8rKFvMeGKQ2liEvVALMUW3mjMSV6Jog2gozeas2Dn8uT+TbJ0iAWEvN
fl5oDEo+jKIYCdR2FZUnEbjZhuzxcqI1OtoquGA6zv2I5S6ilv4n+Qzx/EvTbD+xY8lSajt4uCm5
jEUL0oSyFyYyFT4wjvgKMMb430o0hAzafjMCTaToi1uLAEU3FGaN11M3rWFbfEmXjp+47pRsMImd
U49oHFoCU/khOt2F24cxuEHTwSyhKW7CGJeVkwbmUF0qLadmR84CuFQEHQEpn3SvSE7e1LKW99er
VpR/TDZszTNeMgSIuaW1Y2MWFuKPVyOWqajXMv4Bvc+pfTimCpnoEKdVSXUtPxx85IkaaglO1IRk
RhNJqAai7Wq8GqMOgcNUSzHyODkF5zv+FZDUGdwJkMk8JWlYmmyz2/ASYwZG0AFdMRGbetiZWGcW
oCMhz5iYYutPgyegVw8HnD9+Ff+CSyv7g5dp1RHnz3f4B+/TuFECiIhhZ31CA/nAROu/86JzNP8K
RiC0+uDRBQ3QlrYzNHZmvH/99R2bsoAWHWfe4Mq8gA8vdMR7dR1GBSylRSndX1+Nw0mBLACqDBCI
M0XbclFtm5AttTfzg2RYUyv5U2LahoodeI5y2BURlau1EFJLZeY2xnpe4nPBm7w3NWlR6E0lHcp8
DmdeFQ07oXG9CF/ixAm5gVqO88/w6hGajlhvydo81furMKO+BNhMx2nRJmPAn5JlpeiDSWGOUsAM
dY61CgzfN+148yf+vNTdjTNa8MX84Hd/56zOaBDLlJ2yLqESB6zXfLnU/Yt+r6AGo4DCw5Mq+Jaa
XQZvYlnNWsoAGdV3ZVSpabp7ENjyH1ICleTYzwITWmO1gpyELf7/26CkdtRuhwUvuM8XzBUsZLXi
v9F9XQV5VutzLGlS31aZ7DRfYrLde0uCuHDXhKkujZrXA+YgFGcBcHklxIOjQttAyjUeiJ5TYZx9
+stJuTfv1uAEoVWS9eQS8HJNg525iVHIojYsX3VFdE/E1QV7ORsjzsq7WePqeC/Q8PZqkdWjei0t
cmZoynJMWMiP8O9Wq2JA+MlSTUtmD818aPpFSJyQ5vM0+r3hCUy/86sX5Ov2Rib7g0FGzrZ20748
d2yrL2CFC9Thv+wU4FBmq7oZey9sWPlCDOue6GLdE4dsbLqhz79/PUUl1MNgsDvpLLIzW9xcPTGp
Zc2v1OkzQmV3T15n9sv42QaZLtYnJFX4tty6ZFZC1lQmY1cSSeFRpp9VH+2bIF6wIL30yAIgqY9q
1j7OkVANd9mv52WnIs+nrUDtcXemQcf6Jhe/6HRnWATByvqEx0fOvCV82sgOD58MM8TW6JulQeis
x9g0nmN74lXi6kMY6KmlYGdTO/SeoiZ6xBs1uY8blfjfw6uSaDLVf+jk5uUyT1PsfeuraFOBE1hi
kpDrUjF/DdIr0EDIFjQ2v6CHF6zBVLvNbsYAsuQ3h141ooXL9w0KmWYf+7s0AjGnFiJokZsYNBYg
yI2663aDtYyYpyKdxWUCmfd++OC4hbIDn9NVGTP/S59L0QV9wHU3ajYS7M6hvbp8S16cxK3cLK0H
DM44TQTXykAiEPUCd5f462rkzNMgThRX3WyPWWJG43n8MPt0adB77Yunvh9LsS42Wup4TQ8Rgsoi
hLk/epxrGYLajB0s8mvfuKJM1ajn7+n6bFemr43LpmIrhh+mS0r4pcILj5tCA+pe0OBbWxzvke/i
CFlreF4LdNamZAaeOFJKncHfTSEbBKMFqbNk7H5eQcR2hGob/V7QeT8jeBT+7VJ8niKELQdzSvYd
nuH+psRkJXr4ClPvLOeF2cHyTw3SoNJIMJzpe/DP4GC9qJm9mBjgARf+YT+YeHPcpKGXu1n+TSGG
GpmFdoI7HjGSnl+K1+h1xbAxrsuKv52pyGjIAKjfRyhdO7X/HrXYSM0FH+mfuOzTb/84xqnfFrXd
jmcs4rKBazqUwJeH7O71oGEII6ooo669a/myhZurpEXEx/FbtEcjU9a/P3xDrTNtv2zLOnw/0u+6
eQ+qDGezeU/I5sRWebNNr5vzi/SM8QdUfkq6/W7hEK+oWnMue1GqTs43aRoNvB5SMDrxQij6kuKK
RT670jD08W9qjIBFp4kbG4zJy+bvmgQMm9vuPEv0M1L9QAD2HCxUZw3+D/yZlrZPQPWwkE1r6CQY
v0pgPxKcwLCsp4ItfBQ+acT7LXZ1+YEzAVnAJBE+dW7PsOk6Gm29CU71knuFxiS1MlqKwm7xRu0X
4nol9vmzveWtpMOhuHlcVWg+TLuxVGvmfyRefo4DfI9alVRbIQUUWUE5LlDiY/kw/6X0XYgFbWO5
J18jfcqQnbG6f7gehFGj5oXQ+AHcQZ3K30zmR4D8W3hqvD1UOps/D9Ah7gcF3s0HcOoKboJ9Pr4o
OcPcxTqC7RTLdRA6JXaRCGKvrmGJ1U18V9vX4dOPx1Y2wDmL3uzsUJ51GnsEmc+mtHuXpBQYL3nQ
wgMKMXba7dJQ9hhCC7/g1w+HFmYg/+y4xHtyqI/QUqnRUrsorZPlwhPgnmgaJdjqNh0hfX9mhi1K
kgP3sEEDcEbySnr+PrHqphfNzimEUytE6YFEyGnwAiDvN3KjL2ghXz4iu4qsdvGz1M3aLO5BZuw4
HTVX2+dDePIYDDrnt8odlN0bY0V7fL7wbcNljU96I3eBvPD8IBt4yHor2lpBGnGrKX4AvKKn/nWW
rllN0BFTa2r86OmHNuGyV+Oqegs5SuEB/jT7zGhdQOtrvmF5OTkBOJ5yTqYg/78vjaWwwTn1Cicf
4kOZvBppHGD1mBvWK01caIRsoo1gPJ5gfZr6BsMZ6PDCYdLSRsg+bMmZzPA9TTrcvD5BcBpuxa/0
kAx6u3nlb3K/iSGAWFEG9UFxhXveA5UbDFloe2ZGC/C0j20HF7w7DyPN6o8Y2B7x+ZHFoMJxDTM5
2wFxc9DYnLI+9dALGhVsUM0L+5L7lxTEJozSO7b1/jUqd72AggeyxXypXxDz6p7Spocg0Vwbwj1s
0yeCoVu7cXsxI6dxtyf/fmRH9OdgTnSstIyw45BV3zvTaHqaFUUwLfLWSbdduo7IHJwGfDzapE7b
C9SaME61s2DkCcRUX+qUHTOSrBJtfXC06qYnT5qn4Nr8qJdJHvYCX0DvUjFhte+wMJ8lNnUuosyK
S7cyuJrv+HJr8Mp4BoKxabCRz29nFFZr7zoXAl4AK3sxZarvfzAbtRSwL2IY0dU8ADXNbwXxEHNK
fGnGkhu2Q6HwhnO2N/So/czbPpjOj2kEsW9fnnvxPpMTvCMsw6Z3nTvfr7GeEVRmISbatDurIurv
MVwQ9jqC9MhInykP2bJnIYXRj5+VRs5IUyCkxIDZp+9uHOvxKM+1Ztu6StkRpiTn3T3OYTl9UO4W
mq8Lw+u/EjNhMT4+v1F95cXZkRSQtoM8ezT/SgZn5ZP9TVCTRy7bMSR1hs7YiIiwgImmYK1r3oAE
jEAw2bugPv97n5Q4f4pGH4L3tGcMxC51AmK/BU0M9LBjh3Q4815m2yfUh2t5To0fp6DZo95Pi77c
VW3VEcvvNpIK8amgncGicSUGUoxbZR7CkTeaYCCCnYaalR3hizdCFVK29c3o7CefNdVRk/THnBfX
4DbY9T7cjzY38z5YQqzd60Vp7h2jbdo+qOqRL0ARbMd5A7ZhFEoaSF9wpKv1ysTeqj1T8+1auOZo
D+3kH5mxygrk4IC0t8NTFBIY5CQXCqU9QaHEXycLs1rFgnQkOO7ALxOvxkOxLpewn+BqXF1lmGoz
FWYTbHVc4Dbij8snKzaWs85aGlB2WZMfH4XqhgBxpfA+qb0t83BHv/B8piPyqJeD4yEGmXkYyUQm
l4+imTEG3K7aWDYcZT98qNldkV5szPQmB1gyb9nRV5EL0xXXpCQcauKyWJqyQgdO93U6oN6kzphz
rajZTLI7nrJW2dWE+yZLFWprfyXrzWX/v84687xSfFy+2kbHif0vDcF4afI4OMRpx/JK/V72STHk
2eU+E2EG1AKLpAi05jdDR1Wn2xKhAsCFaJInKubU82xgMtYqxAEBKWe0MjvLsedEvL2t4o0isy40
me87oAdyz6tG8226xlzNNV741h6aZLLI/xQ1BQ5wscXBs8RPb87zhPn0LLja+Y1/ofMuve7hIPqB
MrdBVlBoWA4f19Dz6fAf4Mgz9+M27Gn2wntw6Xq/1FiVumOANjAxuwoeemIzC7d6Y8rGFteDjsSI
YJ9ENiXmJfo3L9BFIDT63oQP3i174eU+xd3DGt5jQazbH5b0F3+4JB2HvARdAlvChCFEKBNQ3Ayp
xA0YsWAZsklVGAyvp7ayldYIAbI2Hc4yi7Y6MKmcSw1BYOLjcAWfO+b2T7TIq3IrMH4ly8tlh3G8
m9DCvD4P7mPcg//PDNGTmzu/RIHwXFViEhwsFDKIsnOF43l654kYdu9XCFIQZrcB2UGHBfRNMyB2
Acy5064g3hlaHgi/4sPmlG4R6MT4YPONbunlPHsr0F57ZgiZSFeO6VjiQ9vpExtmIw0bnJia9w40
2snvg7q9Xg5DXwCjesmNL3qVr7X++kWkZPWMEJ0YGl1SWKq6fQDV50cozCtFOUIVD4FFXDh4vFq+
aPapC+75mU7fi02zhbg12dV9EJNzWXKE87kAg8+NEJxSZvt/8ER4qysOyp4u1/zc+vpPktxR9D8G
TH8Q6hfR3lb4YwLh7HUvO5i7CaUvJKHVQ4JmLphpvWbsXtdog/7mAzzKPprpdifw6W7dKHe8fa0d
bH89LZQBUIXtqUJlIu+PCVFGrBt7JtEV9rNLtaHlJ6y5bs4iIVMDsS8j2eeFE6OsfEzzSkFoD9l/
ZONKknk1vNo5FKAPJ9LeeS2Wuae0LSQOUyOnVwXTftnqCS7D3P8KmNZXqWQaSNVDgWwLaYd1BM+d
+zWAe3LHttD7q+H8HRsrbrsVw7faNiUvQ/gziYMlq2yJ1vXnDZuot0Gy/8+XjN2PNkyXU4YGEf+3
6MJDOdmSql8LsrVFXCG87Wlvm3xcJpIfCjW72vYatgY79Rzh7DioLnUHuwQs0m+gBswWR1LBZZf5
LpPl3WnmGoPYBr85lgOG/8G6miCg0+VRlcUtiFlOKLbHguTBRBKAPHPdlhGrBWfFdmfxA9b5yF6n
AtSpblM2O3wsi5if0Wr3bPH8BSKd8BqAI+2pARNKkh2dwEZM23jgaUqU7XnEzY4yzhGa0noCtagm
35PgCDQakKGwsVda4fab8WX9u5jM+u4AZ4LOJerzu1xgp4Be4n2JmN2EKHUXQ1LlicfxDwAJOM5t
/wU2yZLzevLeOreoXoe0myZuaVVZFI3suvyDNOKz6XdwRFrG48HOiNxDk0ezhLjQfeIS7aO152Bi
DqL60yxv576CYAWuyM2otHJOR2iHs9rrR07T6Bv/Dt8nfqRKV9k6kMYH4+B/ytpmbgBkT4alS9BU
0+aQMu/MMMw+9R6H67cYLf/85fKp1zegIuhqXarU3qHXQF6IyA8d7AcpmqW3ito9d6YjM6G/4kP/
Pvy64fKnYuiwnvQik1m79RmesvjzLci79A0HOXMkSPHkQ9uxtdv+aMPpLBkK4f2KiwnbC6rUiwzO
d+H66+EdZCSBFMER5OYD+oQKaOPX12Ue4TNsq4gklfZ/7mG/0CpYxdSJDhQwcVHhuJjQNjyXp4ZA
Xtv6hNXZepvJtaIUPYljF2l72KSe9ayhahMmAOk3oUqm+9/bwoxLw93C7h327HfDiFZJJ3eLDOZO
rhbE6XtN21wArG5qoxPWH5vSd+sJnOzXLQXsvlmqXqCpVbNDWL3cQGhg2DVym19ztg+SmZNANRz+
Ykwhdu/QanB4d0GwNIMw9qmZdqnJW3JpWnyHIRNEeomWi68iRxheFXs2N+nxRYT/Z7jkx4YgUx+E
95kA4hIfO5mWmLOV62ubNWGBLjA7xDe0Iq+RR964B11YsCZ9sGAe3NS3p9wYXjm2O7VZPQh6ujEM
dogZH3LqK85qZ+zXR/0riukyHDwn6kWAXO51T/XPmHs19awd3kAtE43lSSpcClXt722uEPBGB0RK
ZevoEcWnJ73P/96bJxTSglwADClzVUPAgy65xZu4a3XlSzMr+1kR/8JppNpEtL7F5UbHAT4FsnCr
VqHKy3CXlgnY63n8jpEZ79fXCdR1e8f0Y5/F05zaIPocpon++truX2NwyPHc/TQVctAK+yiZpDaJ
TWA8v7nKgt8kMteRoXfXSU6VlDUHRWz31x05nGwnDXENqzSopnmDtN55uOJ7ywLZlWKxbHBgie9d
9RM05ymiiFxqIYsBSTy4VTyLerlPmvAnfBqUKTcpIFzb3tK4Y280lUYjk89jw/reLZVGo+Hz2g/z
1gj65/Vh/6RpQnW2k2odFgc0RKS3nOExiAdxeSN8+3v8JgYWS+V+CuITiHa5DL6yjnq7msIwtgDo
Txmg5BdVDvvYEiGmSXW69iH5EFoRDrlxM7eA24vBQ59aGWPP/dxhjiTqNhYxwnNBZsp4Z+BMRdRH
Vlba5g9OsVm5c6qlsRjVAyMlyomqPbFS//hDEgU0uOCW8x+4eeRiDNWSV83cs9CJe1RFr4yvXLM3
xh3PtF2RY2mLn+8sxrbCS9HsQvLnwkoYzfxgm/1qEwnpMp/mG1C3TrdgXnCcA2A74GR6xRHMgZJ3
7GOMCm/JVtdmelysNnbeLAUzXd2NuPr+NdZlA2o03gbT8xliEtjo+/mYYeUuwQEK8hi/akgFGWQx
TfK5UB6k3hdIIOt51GXmj+Qx4pYP4MCkQPcRNSzN5frniSQeuhHGTWcILMIAlKKdpd3w5p/KSj3c
jZ3+v2GuaT4Syc2ODbGvmxOxAg+sn+P9PJwS6VjqsBxfpcid4T/BUg8SB9oMwTnBreYVY2QpOusi
duB9boZWHlqnSDi+P5GJIxBP+zZyumK/0QNMfuXzeyvRVvkU+PoecGWUtftWFc672LCq/zjdPHFz
LOxGf7JcqLcxLfRQO/4IcpyNrly41FC2dQr3DsolFaBwFQY7jith2ZKnsS+EcFhaSMiQ/CGYha5P
5lDu8pRIMj/o+1ngNKT79sWFRNGYincvAMNnIpmrBg/+rf7NbuoKxJ/rx4K3UIZpw1EP4ZTi7K4h
e/SBNHsShDEUA0mzC1bxnnBNqpfr+KKmKTqOIgxtEDbGrI6uLZaaJYB+OSklqxL8jcWFEtOh58zf
RJycxJqCocyvDj4TC4q6jW1YC5ysmA8SwJyFWOfHBIn5sJxpu8Tqo/avLl2lm9FqY9IpMIpeCEZ6
NRK7ad+aEwJYcbLInMmupf7ZhZCedCKYBbfm8ZfmsSzaWKxKyWfvycqC1HCbSHnZP69xLVPB7VEk
KySp5ExTM+ewPS5sVN1U0Sk6OHxqV8yQdRprxVZx/tKeksix3nPaL3tS4kkStvHOy/Y5IDYeHGBP
7R3gPCr/jvptw05hQwNJ0F7wGa3tkJERAPRGjo3FbVFm/AJriqWh1RXofVa+F0WgP7UzIe2P5N6U
xnCxfsFvfYa4+r6tbMeqWp1hfdP/BwbZCaDRlGQLaGMbwheOSCBUT5PwBZk6uJlqebnOVrmMP+Q5
BwEuAIousylOeFJRGWAEKbIswbS0eENAHDQguMNPlc4g2dgIB4F+UkC8+bThBftNcZEGQ34mP/J8
bPb5INsxNdkHlAYy08p16gDZFZB2ukojuf9wvKP9rsfELoQFFywLUVTKthFMK/GyAKeedn97SDN/
qe2Gxd+fgY1SSu+Z3m++EtlZ/qG5yUiSFELZzapFfM8l+Wo8AGpXW4/WIMuuiGbGQxCv4SMXmnAL
4NoeHy5BT3SP+6r+V5E1lIsO8UeeNwv+r9Qhq9Qnk7x2fklfP2RH/9eLlx95cc5DZoVJ1yrjQhYq
grylIJ7R2tsQL3ZW39kx4L72GBhVRouQhLmtX9n4oABj14U4fU1qW0XzCWLTnAAwU7P3ejd2oJ5S
Gj8SDxrrvZo5bHI79ebilP9SkTTsMPBCNflWloFlgt6u+IjJzER617bUO2Tmn4MXpMjPor5T7x+a
obNTEg09lMr1u99ogZS6MH5mPsS0ItTN8Q/IjPaVQf5eqrgA2YAZ4hTcbKCTTQA5InGhOY4alK2H
mBjSb9x1jtYDRMl28eGlo03pH6Vh4lLNhX/xEVFIE9VPWbgm9XAlBobr0uz9vGSXdjPqBit1T9Gt
1W2mASfzhMe5Jj4Eh5Odo0Ugqy06DCM+czS6xuI99AwC+JJNMPdF6c1CyzO/lKiUyP5TloCoktJ5
JVWBkv2glwdKOW/+76gc6+Sa3qbRH8vMyi/xxZW7VhJarcT5Fs1RovAjM8L2XB6U1vnLQ63D67YW
RgQyv7dojT0hGGO5LqJ7k3yLpiMtnszhWoiYabEte8zj4ZGGzlALv3wD5UayrzKMvUBZtlANDPwf
Ry13tYLq7sqX4xZ3g0LT+HWjesps3B1HoVnnEylbDndC6/eXPPdK72xUvwKT6uxhCP1ieV74adtv
O6Wv+uls1YHRFy7vGVLzdQFVkyCexxfL5R9BJrx6Ahf2Uy1X64Goidv5nr2Yr9dZkdgUf58jrKmv
mIuiy56YDiWUxuIVdp1TPMxYtP8oBKNJRCoopZED9/rChjECSvcwG7HxO5w4pGfJgVSx9pWphv+w
26htCpBh1DxTSv3YKVkm
`protect end_protected
