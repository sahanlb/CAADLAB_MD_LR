-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QKgf06Jeui+vhnslwsUlE9yUtifw0Jihmyhze0uMJ+P3Y7xzRJG0KbmcQQftlSJcN2iHm43cMPtx
YvZd8JjjM+e660e+X+Bw4QlSqZ51lAlRLljYhcS6MOo5a706ZhnwbsT40nzLI5y2oDmaijWf4BvO
lJ/TG7INMfph5YlpPNjkSSTeqTCwa7h60yeKgGivf1hrnCr+MBZE2vVBfVj44PN42pSS74WBupYg
QkhTV+7QlgMo3nO037nKCh8F+lERpZSfDl8yX7bimXKBQ+S8Fc7bm1KY0jI6m7SAyGpvH5jalJSh
nIvbquJEmq1ZWWudx6UFw/uyAHgChg2GF0Wx2w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24944)
`protect data_block
fRdaobf770BiISIa4BBLgGdXirVukph2vPfMlXffHL0i4c6Fuy9C/+mftLTdOfE6jh/m8yAal+Vj
5f6H/LLMOA5Q9Swslp0Ra1198R9J0m0zR5Wb+hgXn75iSRdr7Qn7jQA+L/7SB9bVEo8mJfgjBrwD
HonPw7ky4Eg578kkLeUc2MN0D6rzxNJRZHfeoNiT3ZcxMycAUmB8ameyt5Jnx6Whlozo0YYR7+La
/lAdX2SDIAD5SzvYGSmnGHbG/UluZwr1QowU/u5gscrTuXsLFojHKqaca6iHXVIj0v92goMz79im
FbAP7JJO76rB2WDO3qU3BRcfygKO4tMHsajKd7Fs5Zuk6VxcGLHT9oWGyvLPQ1/Uj+AKbSU55ZG5
kDTp9r7579hrBd3POSxOa4u8ZWFs4TvPxs+jiSQk18Rdga23exCcJOq0IDxP4gE7Ul5s9sTuHCEA
WvmNgsPAuwLQ0rGHimRZ+JxhbHXAUVsZpA61b5iaKFZpqLP5PHjSTT+0p2iwV8soxY3UnBOsiWW2
0ybI9NKt3uIM5JXO7I6sPo1OM/zX+90SbgghCtURnS6NfbRAZFL6cJsAvWLhc99Url9iSix/5CSa
Oo5VOVWnNLFYQZvU9SbXegMk9jvhPKVQsSWEFqMYDYWRecZGjVhoPRrVkHsnfL/TzHNTbqz78ISo
ZNqGCMoF4MfRLjWS1Ff/sRyIfV1pY4rft1LnDfNc5PkDnf6bBS7Wr5CZKu6pzB/0JVVbke7cXzLg
eiDVe5ghxZXymcfzMkz+QW2LuQdf/4r7m1GbEsXViCzcHNJePCzS91vw9iAIhzX6MJx6KQI8bCXI
VwqM5qB3iklkEqoykJueGJViACwWbI3U9xfF0HESUid2Ok37CEyrOi9m9aGpdSsDExptpe4rNEuN
/8Q7zccgHgKh/FMgdRkBW9pxaMIMDHkYBbBYG+8b9CMdA9ex3c71HPyLzTxuKnA3wBh9LIVShpZp
F8o6pSN+wPDzMdyZGTW4fmPt/29wn7E4kkpicwhyqd4YQ8YhcvDU9P/6YDzIE1i3AAZ7X8pR0Z0C
ziYuN8+JqndvrStN2+2ma2gY+BWWp+cRMVvx/iq3i19cS8vv+yB9sVclnw39pbPGNVZsk6NSf193
7g+ggxhwO7C9v1sbpquoBYYJF6kAAL6mnVEIimkyPm2pw2kQAR48ylxpqNMK4eP1g2wc6FtXKykd
8Xo1uS3OME8EuJXSSsqOHP7Uf8oB2MHz5UYx9JFRtEZhWMk5CEp5CADwvZQemiLEoxI/f+aubYJj
Ynd9gGD/Dj9Dv1fB7ZLzPhiL88R3ckbuv3Ek0G74L0cUV3V+YgcLvGaTFd53WKYkYztuOXs2696C
MueM4Banb3++CO8sisNiWBq+d0M2UE+eYDdGYChtP3aB4rMP6lGSM/mNZl3mUHpIbl6tGGkmnCu2
QMIqb/4Rs2RAiB0YrJlMT/hoR3ALEdjEUY9fZnazcQPWmxxNidU5T58xy6x6cTJWXY76670g+EwD
e0U9oQyjOdAyBH79lVy0jVKuHmjB/RxmfqlwMx6MnfNeaBbvTcSxp7CabFtmIYOkwBTWfBIlUjJe
TMUy7YjqQsBhPJTGGtg1/0Go3kxR30t9829TxoqaxjXAVH97uXI5yxbYEeIbEvwQ8gF05AaFOwij
zCaduQoEOiOyRPBLSjMZodmF5n1E4PUJdJAXRDcLY9QJtw2X2uvGjtn7+AP8rUdCSNdAPCVRBNsz
isXHhD8gw8RTsIXOJo3clOuZfkrjrLfNmhnxT10UcruxPNy6MxGGJdkga1oSebhdXrHrPRNHawGl
FV5gv0J0mpOoZbNQQinDDcntZDAE2cuknykuHrSniEWG+lLwUw42nTEUkEF1AzOB8cIslzKZqinn
OAHR+Xc3ktoVswgFenpPVu8jq85z1Xzl6jyDnYj4/UthUFKdW92ZkhburleWKiQScH/zjL/jh1qV
ann2bx/PzFEDbrr178QAH2VvP6wi9E8x3vLwfmk9GZ3pOn4KDaDK1HlBZZV8Mtx9dvXAb/RNnhrV
9cf00CuWQ0lDaJ3cO1xNVkiPMiqq7SMmbxOjVblKBQwI3O0PIl7768R2WKnvyMHvLLBKTpmW6Edy
Iqu3tYJHMmg6lq7iQLsEL2eQKhdZ0q71hHWvSXRX3IAj25UabQED5SEj43bcBJ4hgQP9Yq+18+QN
Q+Kw/mZ2NQ68+aMbGRckamXeR/xD6Aw5yZrVt3+Y52QFElUKQmoKnOvi8N7lI1w/zS41Mdi6qFOs
HZQZtZGXiqJrlOca1DKgtGgrMse+sX4wEZgVYNNEHrxO5Y9sOYAJFlDcrXVX2K5lo/2qSHbYUyil
FmyuT23cDprtz7ncjJlqF7UNuTHPGtAuR8SkIYc36Wud12KWl8JQbXnnkd4MiWLMIhyle3wr05y8
jk8ep4A+CRnlrQqYzkfUaJr6ZCQKNKi4gag2TWucQNuORNIWnOSmPPLKAqDER1ZN1AU3F/d9baEj
opfwaO3NWJs00sAWhDqEFgcxnPfR94qI5s2rI9yMmVa5MNjn4T4F0tKKoru/fBTUbmE3JrbZWRED
GMkyZPVsinZqs1p/O9bULfyW6SE/1uvVW4tR5aTEmZscfBoWMjbctJVbZZ6ml6igN8NY+DKP2JIG
d2O0WZgQsuJ35UGuyfXN7PCfnBGvmfv5ErIsq5NOfdHSr2Fo3C/dWzpYCTinPLHUbyVNERzHT6y3
NV4dwMLTVY6nM/vHdQdGkztFMADVMl87jtjkgrmfIpT0QZ0LL546W9Uf77AMRDmhtDQlVE66NY5P
DlHEZ7gYioiEv14P9NphmrTsEX+jbOY4HHsElCLE4CXzwBOLDn45GkagX+UG3zJ5MhE2p8BAHvww
v0V3rtymstj9i3bHC7jRIvTyAbLpnyCCyJ7uD+/mW9YeNvCakf4mpOjUQRUuBGrj4SAvHQwzwGg4
1RrJWQtW2PDgXWmQAge6aFiZmzPpHOQbYVA7owecsShP0M/h3WoH1PFl9Yzhoe/Zmw5xovDIbnfg
22keMlH85N+I/ubBZ4OPfwWLbvA/OI8hglBx4cCpeY01FWg5wsBbFDNt/r274+NwokN+/zj+plCO
sbcju+BNbcxFl+BU4neyHi8Yb7cwZCFZJeeBLIibDVKavYaxmk8CQJDTMBfhH475zPqT/CkZoeKQ
0UenY940uEgzMeV/wDZGj+YobufJ9ar5Ym9cZoLMM6I5GgX0ea48+4Vc3Ek0/6kx6HltPmuIf5li
Oe/nElVGJqBPm7ElxYFnKvxKo31JwOz6CNI31Vd8sNXDooBUeV4qhsUWbfEWuRjmk6luFNrLYRup
exnCvpDSzZaWq41g74Jf/1tSd1n9e4boY2lx4s7l2BVOm7y9OKpAG7cxK+qgKTOWuc9NBq1TDISS
Wk6LOmZM9Y0ipNRlKmgVUchaAGg641ypigdrVjPBN8rvL9h5q1+V0hGc3JVOdJBJfeFN1rAbuowA
OZlPLW62Gnu5ipAsxAnqThYHeLGHmLTCufqbTn6veYnc9qXwG88ARK1/NLKYI2qNozyltl1qnUz6
2nzTPHxO3QqSU8eZRFA0CrC+zuxYp1toooGg2lXNe21KLPPp9mR7ctXIcjpO9yXhH9YFa0BCYfa9
OUa861m3GDMzlQDhaCdI/Tadikx4Cr9J1tSjC+pAxYnK0Q2omv0fgk5IABqJjIfSVGr9o3z0YstV
KVh75HzNH4cV44Gf+nQj6vfZT/+VjJzfsMkCGjuhnh+KXfpQzcjD+3e1f8BkAJz5Xm+H6Pdck7Jl
yXdXWc3RlZ+tIFwW1kZbPd9F7cMIuMJ30kmIo1v/cqIHSWxGHAAK0twXwWfcdIkRrdkIUFXWeOtR
TZWLC3DO3VMxOp7ugmTScqhqMlPFAvzpAdZCTcrNcet5FCtf9hyp/R9qvDoUXScn2EhlYYYO1VS5
jXIUkWG5lfp7o1VoW2OuQPf58GcF1pEKeNDTQ+AbbOgTioGABXXWdbz1djf9SNd1603hw9edA+F8
lHJcZvBE4kMpHWwIFe8LeGmPZB9Qs+rUzYADb/2ACsQGEKBCebrovj9aTJ384u7dKbcV7+WH7PrW
wjCzq13SGSTzIuLTebkYqK/5zSay+qzVBWe+VvzT38Ej1usTR2jerabv5dFmQRSv8DauhB5iDiXy
s+OUKTHWY0S85HAZms+lwth6DF0sa6MUY+2Ba8sJ866xy5bkYfNtT4ZRAGk/0Y9KVjabhGVOdZbA
sMA51S8Ih81Wt96U/o3KXNs/fn/OwinLUJ4BFkKC8ZXrzf/QTQubDPZXVlFg83UmjO7O+h3nIDub
oRe7XIEARA6leJnEAxJyxKBA5gc9jSmB2QV9V9I6xAVdWPJymixp4LPCV//3mT7vU0k7FQb3UH/w
bi7cqDn7VbFk9RH47uHCD5JHXCu31tSMv5vPAatOcfZf9jnJ7u++AIHJiBPbGlkluUIjTgvsMBoG
vFAc/8wZxy+47SC6MhvdcdDJfpQB4JUigpZ5w307l0TODETxiLjgn4on9aXXEaj33PzsGkWhjk+r
Db+gavbddeV2HP4SLw7bKNYeAF+lQqJJHOQ8c4RAzrP1niitXetTO+5W7u2mD1DaPIAvvX9cpzzQ
ehe0evoXG+zAMRErurfJYBd0Qu9tKSFH38UJKkJ0nb9+b+9t4B26SgCw6Cr/suFrje/5JWrqsAMz
SWMn/+kdfrRBay65Yd6kYURlvZVb5MQL3VxYxGxVu1akKIcmtXdzuJALLAykwGlkWxdgBy67yICq
f/avGt73biN9CxreGq+FubMkL4iz/BUNDINhVGc+5GWhTf8t2gUQ7eVvxKjOFJu8fVOCQ8VqNOCW
1xgOiUobSYuH+edOfRGRWMpa509NHfJsUUWvWO/y9jBv/H1qejmbjBPFVjLozuKEnbX7+vWFpFv/
rD9dIptIioH8+uVTiMgGgONX5O6Vm8U0mGN66TvP8TLBdvJSV2fu0YRZgqYgzQuvKz1QN35M74Xn
1YfhYlcYwHgafN4PIhreWRYUddjHmvN/FMd/TZ9rLaBHn7y7yc7OSxbr8dUO/D6iew+J937BI0jF
x2IqoZ6ZG6DHBPrQ6gVkxeIXNzNEoCKURCDDQxz8r48VSFwTeLypKti5gZAs8/zfkg6lpnQvPICp
LZiCcZCGfUGu1lUWXV/Mxgwyywl9SWDkDIeobyoPQeVT1QF/05iG2arHesTTosEj8IpBaILI1ojQ
P2Rd7utJ1ui3/B7H5Dde4SF2KMSDO/sA9UXpEocNTYa2UU5n30SHaSYbiKD7O5W73JkYSo/0ghZa
p87v7ie2TSCkIwpL9pBrh9HyO9bPlTdXBVswG3IG+SmKwQLb2+jb+ELKI+TcDaOTJfPTtG8vAiQZ
H3wohJO/fM1TCinuul9n3vLDc5FGxw8jO+ywnX3eNvvHbOlVeymnIZEqcfvBnR+EC9EZb+QNQo/T
0gouDVsDcQwiiyQ2ACqM0SCPSLViKUxoPmXMJHOxjY6BJbJjt/j6NPYvxNfLI0P6r7LDp8WpbTee
iRevMAed/TBdURZymZERDOwpzsScAUfggBhz9KiT5i1du2jxfehRJWrcAUWBT2JKMoVctzyGpwyu
LtguMrKB5IWHebHOAF3nTnvlsH//i0zoVIN5hroqzNmTKff1zRh8Cfbps/3JViNO2G9hd1Yo1fyK
pEpj32hqFZBjbAYn571C9poQnttjEQvO6gcjFIvmLi4MhpqOV3Nf97KYG2wtb+9OZUj6p/C6lKTF
2LfBs8MLdGmYZ53tIMU7C2CKOlOu0SjbaR7iymdLJ79FhNrzqdWI+h2B3Ks1nUJvM9F7bYguF/NB
R0qhqOTWxUAygVyFzjdxwb6YNfHjJYl9g5hOC1UOftOwXtftmaqXf8z9aUaqDEdjQPaYVE0FOYGH
m8UK2vICo45u/gN4BspvWXhww+6WFVA2+OZEBL+kqWYyoNFwKlZ9i4ItKhGYiYZZa8nrZZe7cZew
MmWX8pGcZ8++I+87X48M1NxZ8xWXvQmVG55sj9bcqYSrdd2w78SehWSFPTmKjB9Ib9Zj8z2jKp/a
gHlg/98xzRrqfikQrpNy3zXsaoqcUhOjcT6Jz1Yv4wCNXwBOeqnIC8kqODsw4K/08e9LgB5iZx9I
lHv7/UgaHwb9t88hK1V/0C/hJ0P8XzidwlyO05tPe8NCzWELVfqdvo7oHBcOlYLN2ruLpR93TAGl
+Kgp+CCXiPkrhTgft36OoxpigwNVv1BOItYqt6yLz9JeQbGtOx+rnTie0VKD/Ryo1MRScPdcgTJk
yxc+r15wVmYp+wxk6j07u8sFr25vNCD3KGRaHmLLkDjP66xuR5A5sDtkyM+Z6WC2v/K6hHMJVxxE
+9IBxU4vccHJ3RjkOF8iKoFAX2dUVBef3HGdZ2lPLPW6SgcTby9gLb/rtsIITDKl1qvpnsoDUj7p
OUsB8PTrUJI1mynj79J6Nd+n2RlQZNgkucbs9PybJ25sFyEpRP1jmonKtqAA72FU1oeWQwiKYDls
VzN+toNxWfJsXVYw81xTW6JWCp/d+t0f64dEWy45tOlaAu7UZEODoguAFkDODWuQ/TKfHUgaG3d0
v8GVTy+7gP03EuePQuBqAasJEgbOh1//sIqyM1ox/tThWZTAkQoNDns0VlaCdfGSgaw9x4sJpgYm
gEDuX1yMOGaS0V9eyhkb+VFLwSe8Cswjcwe8+e66I0NuTxVZl5QnfPF2wzmlXMnRP3QIWry+t3+W
55cKRt/pa8qR5/CieFgDbS2yOp5pky+gaAn0RN6/5YSNZuv1HtqUUF0j7V8I9s1TdlCAg8nvBYav
k0PArGKCw9DhoIQ2zbk+8Vd+s8gOZUUb0/5ZpjxQAZog1Tz9NS8JWCvVOBToIPFNgbX9Tq2B+ydf
uVWlD8NBusBppPA5ZbEC0bOotFZWyV1c7BugHaRAQ6LGo8fEvF6WyrEZ84jyAEvuowwqtXO2g1rj
XfJRZuZQTyW/ieK2y50HuHWtwRJvazI4NjlAjPeZUOgCQI7vQc+lrrabivZ53xSBTZeXIXx7+ZRc
dXaqOouzAzVwHPH2uH5Jvycd83HrQXR72PQJoVGkre6oB0Fb26hdYzXDzQbgdQMGpsBgG78G3OSG
w6/+YoktlB4oeUR6ktUOCmQbDOLjyqN3ckefM7SG91n6k09IxdYFjRC1D7qh3BFD5Eth2ufgJLPp
bdGDdJWMwjPsosD0Zv/1BaUHEqH77mXa+KMYTsLyTHTCiPyae7025gi2OhAP0FwWFt9YYW8rEGlu
4pEAqF/m1+liJJp5Nj+DQDbXnDUeOXNAW2DNfJLMUQ4mWcCZt+zRx7dxsiwfRYNBdOkFKMOpJDNm
yEQhQwMXYu2A8PzLjSGidROPJK07DDzAWXAY1VeE4CDwmc07obPxyw7F3dWR37AqxRHsnpzaN3Ne
8G3ZbOG9f/KSqgNhof1Lk3RPqilwmd5FdYoxnkm52nV6OEARMBAEbf560v33Wjwnqv5L4Oysdldr
OhdsdwvRMLeaZnZZ/TzDfKTfAZVrihchcVfAFsqgvlZNvGkNjuzfgN4tBGGhTIEJ2BzZjANuWjsg
8s8/Az7Q3gsxh6krm0nXZ26zQIpDMgtN/rYbCc+XwLjSNCleOPtfFwFJq2Z8OmUmZXSpodm1QIpd
piZbjutXfhxljAevCn1LXZGJf4vUqNsbZcIRUm1GiwG4t6N+Q7y6f4V4wfBRaxC4heeIB8Aq/bz4
LvgUO+XLvQZWQNcZFR00mnzGvSpjxW1BGUFVtsy9FBy/5P+APfLU8GV/TkpYkUiY4R+Hp0Km0XT7
HD0dq1e78ihBZbweKi0qemdKH66DIEeLnB8yklzbYtDbLOn+4+3UtDbXnn4Me02GsE5IlqgPSor9
XLlCltWrahy2wcDTtYDwwDb/eOZlWpmTE5MxVLVJTy8oh7xwM3JCOPjZzwO3xsFhzZho9YH+hIvB
4cq/DcMs8yKoAZf4ScSCfD6OhdpeS2mTI28QnUkqajx8lCRfykcShJVI1RYi0WWi8LCoAC1hnKf/
BFaIJzprvJvUInM4GiMJyBz+aKOLCSuUBUtlKw2CtutgSam6XCTxlflLB4kCN8hdSsbu4iqnB+Vv
wyu6t4KEZSokL1NL34WrmVBUs1cjQP+CXWA3lbHzYNIR7gfTBdrr3I1ZIi2r/LMCqrpTNrmPAm52
9aPMelJ+/e9MYzuzNiOLAqH6SYkZ4KsSDaFpljKeSMDv7XnWcrO0/unfX/oKJaqTnHPNjFsIjWs5
ECiTslcs8+K4P05/MA5o9EEmE2YDtVxmaoEtC71iqd4M05Ja1nRLxH3wm7F0kkqFDcq5aHWBJycn
t0XbYemViNbTNrolUmC8tlee8AgcpIONqCY1oWnoD1h2J9IAzsbWdm1y0/Q2slVhsP9RG5OKIEHS
ygdKomWVQkGU04Pijb+mDxr1pMPT9Q+hWJPe1btwglJDSRMdSDg8zPQTBc1xwiXjmQoSlzhuPxrB
+CG53jGHeJinsi1sJBUQ760i49AtL9UJ203lPUPKEz+aeffdeb7J575KBgjLHfBcN2IKewWpj4KC
Z2HuXYgAF16s972Ows+hbKLPtTcc29SxxDtu6Yg6rwFZuij5s2NfjbGo0kAt8hqJKvVs6KRbWpYh
YnwW8ELJArgwkC9U9SqAsbiy3NnjeuwUhAY7GdO1+aJpBQLIlO+0L5l6UudzfF6FmaxeXvU8zvj1
3fsTMNAKSJu+5FaGXVrvCK/+IbyYIyCQ4LcWpdLwzPNsHZKlyhiGUPqOpZ0ymBUJ7GWapBc2bJpg
cM3sfvDfGfsIVMp+cCtSm33wCu5oK/WPHHfGvKuvzfEfts0a/WDOAqu6frnprMTzZTJLumxZzzjn
jxT/SDEAtCP0UZqn9e0Re0E8wfQKrBziEc8FNOBPjBJm9CN4PGwF3IeCYy55ns3Y/KPG8bzZ3KVk
F88hSXeHhA/sXSY1MkDUi8FC6c/21fL0vv+L+/1fgNxzRHJlajyDrFLRJ0SyPpdi0znVH1QM/Uzz
sMf1QvF71J2scjU28WQ1uVhmAWRniEKhxn/Cz+pvq2jqCyYZL/MQsuZcyBgos6Oo4LlBNA6e5Rxw
j5vlTv30xPCNO+Fhqsvej6+jdGgJUT5DOFalxaRipVS5/F9ac20MxUwAhvy/eJM5WTZfnh4/C9iA
G1vl08f0SlCJoHNWi1wfyz1mzokXrrxI9TkGtAyLhtxLgLMV/4gDGMsBSL5f8kgqKRAWqzRtUXba
rpm43EsLya9St6VSZytRkl9NzwuLkhrOvmA8UXhf0SNZOqk4KUi04NXIiY1BDg65Z17hJ9xwX32u
KUZHqFIePF6rJppvIxbUlMNN5juEQDMzMZDuUuvRVsgMpSuLAPhfRci8QxXv+Qe476GvHBaRDUXH
lov407lapL5zlvycD7HJDkqpq1d/AslXxsz7cD+wSWPLaWYBR6y0Y8UFWI8GFBb2wJ13rdD7cXvS
wmBWBJrZDd+icMxqeGCzO00cBaQ2ZqD7sInwUzPjj3MBvumlPhGwQJIktMY2kr7pjKs/SzzUR5tn
+u04Ryoyhd07OxB9KOaf9mhNc/jmJYHRWu3W0q8lg+ZunP9GGwgRa0eMTw1eGwyF6/kjIRl4e4oq
zLUBihU8TElUWtrLkZNq2+6oKn3Lh1TYzUKn67IipU15VdBx0+IbVEI7stfDYNO5qoVGplHesXj9
UncMaEeYWlwC6E90xDlDka9NEv0i5IB8uaG/Bw2UqKezHLpRb8mPjt2CZRZT0SjxZDIr2l6ESGJa
+MPR1vCbrVhVSKYMupyANmNkjcQQeSPYaRRLrKqcKiGG6dL969d/WIM+VDgbEhXwoORwhvA7HCSb
uBF8Ub250kOek9pdLlGqjBmL7I008zWswB+6hUYKuo36mWAGgyIxaWmNXOSFqmObrAryv6K4oCnV
8Zmfeig4bSZ1eByrkHjEvl9TbtAEKG6cKE2oAYAo2RoBG4UvABf8ZRNOfQqWX7+KFk2xzTgO4eYv
hl9BVh8WlWAhB22+eminc4OIqR86hfP6bgK91OxkiBfVr+Pc7KojWrckBp67tVDIR1sg6pNK2Mkj
zZ9zBOJ0oymMNGgU9Iv/uV3siwod0LxQgOZfQ2/X2n4oolc+UBT90bPJZ/E7rCScFbUaiSkW+l9F
mJhYWPbf1ltp3Wnuz1XO0+yDpN4guVmNBy/TGqCIgFelX7v9yrBnXzccGvr9e+xWNl5Gj+cFnK7K
t+LU6gkk1TXBsF+apOMq2VU/TGN4pl2b3/HUXPIDS8hJdEdxtGhuU8aRhqzrYyq41ETcPK6g6pEk
Cbt9r3pn1jWqSjD8iZYFEPTB56lo77mkaZFLYRZZyh3EIxJNPw4MXGr3zXYhc6KtliTLvjlnvyJH
EZjAPtNFalb2GRHUuXOgOFz+J9PCmcRnqoK45fticKlpsrcR0HxzDMBiyj57vlQjEtz6DSTGV9J+
TTeZPW8CnjCL4nCiBAMbVN6+G8uix4j0o58Mm86kq7muCqEA09ky4M8UbC2CTXOeJGJqfxZ9gY6U
qP7dqClfKEhgXywexbT1p7jZIZ27lW0ImtyaoHNj0EokJ0tFDOqCK2TopJF271y9MWjpI2wztWnW
+V2WfCjRWz9dstvRUx96BoDKxnknUesgvOFufC3cBCcyDbsm4+pa4uPtOnxcqIjhj+evkamRKyL+
pTyOEBN4vSSBj3Oec89lYMzwko36NrI2rdKrnB7bpGNgqHxPwE5tUEHDik8e/Ciw0QOMljEFfiR4
I0oEUI+meVrFUKniyVBdcteNux0FOHkm1J7Ft+5f/46diR+m/MDKk1NEgNthLY/o8Bn9b6uqgfwk
5+fWiqpm5ioHVfj+6YEMSo3itGnt+pPz1jkN6BrQzj0dXErUu/XANA7nOY93/4ihmR6YtC3jmhRy
rItfRC43S0AdrTiTHq/FESWPD5WT+cjOQr835U3QJYM3fciMfjQ+sUKaymJoz7uerZ3A7PVD2tvV
S/RAoLSNIG+4mQCoj7z2sFRqVfq0p9vSBg6bg259XrUFB5/bybrooQIvm/+pVo/GcvkyqciYPuRW
fLNQy6Z615hwlrlU143eXc9B8yZeja1zxZnYjBZIffKbn5w6eGjOqwbWttH/IJWTCX4kFW7b+d/w
40rjKfBjsPSYolIXqWTzHTN8qu+lrve98o7i6LR7ceIe0MX7QbYtIaqoOXdj8tMKbr4FHkkw45HJ
XkVDHqOQ+WbmyfhRSO9FmHKHGh/lV+vmMERh1TEWX9v7Gj0OWzEWcg+d1wRbyPnzpKrk/tkeFP//
iR6JkFIhhfd/ya1i83+Ms6UI2VPm8jrYhdanxcq2m8dofryJASFB4FD8TeLivtGM5NsWPgUeXlwl
do2Ov1MUiRew0lsbHPOwwppf3oyWc2Bws/0uWydKmFerBv0Kbs2xX9fQePQxGArE2DndGs1RF5HA
DFpRZDQeAJS1nwohEJaPwvjrUla7LaZn+W93b0MiCDr1/N4YMw2XxehC4GSUPUBKRrK7YzVhc6ti
lGt2AX+LN4kDdCOr4r4SrkYeHWYdwCOIcW2/eoNczVo5wVLV2N6sKTx8GfxrCGUD/QxD91xazk3H
FFNpwrEtcmOH1qS0LVzH+5XDyIbZkXDPG/ct8CQigmnW27mk5Bq49tNaMGpwQE0zD09N7TeRn+Gm
WKVGqb76lh+zUU+BXqPpOSHA/hxQTZX/APra3NIN+1l3vTKkLvGyphN1Qb0VPEzzpHOTmSnfQz3x
jR7el0BsK/nv/KWktsyUigUeETbEU8RCtFGZ4Z3bhmZNjLNMT0yt1JCogfLINKqn+6TU1bf9kOaL
UdvWDNHEFFM7+wHGICmu9tMrB2WVhEuCBZl/gfUv+ZP85bFvEU9v1YhxFpE8Sv+MnLWFeQ8SE1XU
LtbCJsAZyGZSbJ1Z0jgVX0jAhivzAPL+eZncQ7GYwqTVCsW57EGmz6+hsc9rhYzDl08w/kijDDHa
mYfHcLnuRiCN+3VX8gwJ1xyzroJnojM2qvKv8wvtlSaDAwrxdsbjFM7D9g7aKFUZOdOyp15hMCJB
XiqluE0Notl1Ig30sbqmw0DbIw6wo7iIkaWNvNe6yF11EGsm/PZvHU9ohwYKAFsj3ArwwDD5X7eV
PtgNV1wGDlourn6+qeBHAbN/ANOPdBs8A8qGXOGJX9kmul7wOF9++v3IoOaI8alcaxAWoPHa5XMe
CAAP3A+Q1Lix/AjTyLUEJ/KdZwjSGpmyUvuYcLWET8cs/eScG/klzEXnmvjTlyulqKRAv3AK2hDd
yglRCtbF53XJQrova6OISRbU+gjQeLc5dLmDxH+4kKo2+4qeyw3dhRmCXh9e2abc7GBlqC7p91pG
WsHB3E/PzRHps5TB0YZqkEQg66pAx9EVd2KP7NgFfhW4Ylme0IqPCiAg1ZA/7medluokBLwHSuux
PT/9jqyqyn5A8S2FSnUBXlNcNxoTkIUc5eeh11tbVtYx+rStMqVh81mKhpOI/CeQusyWHJCHRNtA
eH5fELvv5CxqehEjza11DeBzN1oDQEqJMljz0HJdt7ExoTpFloSxV3tWfQBo6Nu7nKUAxG5PzAh5
kOb+SD09Xe/5PkORNsFdpVfoujACGup/DcjAqainUWPjERVMQccGRGm72tec63c8LSbR4V1dXmSc
zuEZNV/Q1CEPsep58ZF8mdKA5oz9enfZL673baKDN0qf4GSbdphBUwyZNmj1B+YqNEjqDvA+eCev
p9GIY9LsYx1cfbXiiD7UKKmxwtb2X86nwr2rFp3vvgNJAhO9enmqoT9svp1hZeJiBxAV8sjrQWnY
5Lo8XUXkweCGl4JpzozdDFsa1SRk9gOjGbtM8RejwjCFNd0ZWQWHKE3CFNAkwJ6HiEqctYufFjuG
F6eN80u5YVygl+fcjFAXzxqC5OaHnCPJvOxD5geHy21foR4ZRyTHeISE2YZ4S5NnZdrzSOjcc2IX
s/1BON87HnHfgx2v+2IaSWeEt+arWvzXiOSW2ZG0R1U0rKWM5psdY5gKIjHc0yVRc1TV0dl1uMGn
S4X8PJI/XYF+qEUEEPbcSN5xvCMun28xOQXIks3HD9Ms60bxlcInAw73tZYa5DMZoMMK/3nDscHk
NktAGuJ5NAsvohU/ijFX6Xz1duvSDljiqGFB4/nmgN9YZi+Vxz/YVdEmtUwieUq/eWJi5gv6mdt3
iYoBPYQecNDphBhMY53WVdCF2FSdcEP/uK0udrYWwTNze68hcQaDYsE8u102eT/e0eWwAZK1++VV
oQVwVhIgUpKCNbn0KAHYrXvscj8RwptPwN9qQQTsIDh3hGQ6Zai4EgW91x3xtImj4HAdbVNsymWb
iElfNvCUiJtMBQCxruIu+26GisIlaK8bbD0ON7gP6M6YslpFEbcsqzCiufmqjELv7rdXbeIvyi6Y
EjA62Nn6tImxBnMwxVLEw4VQfrzCXyQHiQqQr0pedaVJSiOhS0I6T0R9RZ6WOIw34Oob79d1TciU
ph+vMWgU7O4sp/CaY4DZK9p9E9nr8eXZjolEApzQs7/yPIDQuI/tNVYkxS4YyvJmuo6voWgvB4Yc
pn95ebHtA84GwitW9vwGUe649CjM1bx8ZlGVYFNVaL6QcPEGBVXEicUZ6Ks+OZT6xmneeVCzEIF7
TqmqWVqdrGAcaJt72I7ksH/zaobSsufiR2FV8CwOy8Ujet05RTJ3Zx2hl78Zg0q7sM8vdThui2x5
eiMfALMPFHOc0CrgQnf47voNa7zBAMvZy5uF8DL149rgEY9hP5MPuGvWYQy7tPhOlP3Wz3k5+ErH
PhWQ3046ZVbqhl+S6o1xvz0I7omtbE1Jl7NGUWeDUK5QW81wVXDh5MXqhRTIQY+sNsbKJq12iHjp
JZ36+R62iUrYoCUX9ynEduDJ+pd5BTd9cOFlWYDUWG7RHZeSgWPlodSSblInBhsJXOsnWoJV3iiK
PQDiWVpsojOGc2hp7oqZ02Z9uMb/Jt9AntlWo0OSL9EoI8MskjeLvDG/XiBrzBZGZAx16Ks8kY4N
8JV7zoMyEx4DMKohQ5/NwQCyo70VgqeEITNueg8XvHQtSvZ+7av5lxCwP4fARYdMr3KzTqs4wzc/
8Mh7HRwpc1S0i3QHrloxuYe6QBDK7KnzEo3xWSe7rktLpF9oDNS9kbbaOjY0GT6uO+zktBuFzNwP
SZ/gLyz6xgOXbx029GBlTq3W6SX5O8bbUqB23xr4etkl7byd6tsUARFERdA/btm7mNU8nkAntbqT
yUHPS2Gzq4twnjldmwl/er9CCyFE9YH+AcQRibHD4xYKFuQQb2pnf4Een9raCDkxzfmxbAWhcaDN
AlSkTBbPdFDtzWH6ldxRJoDw1MXn79eGYBjEUDyCdUvCkrXHkyBUkKmbJvkKHhIn+U3jtTZfBm2t
8zOZkX06EbyiYa/NM4mBckE3c0eAyLGFTTO8+RuxNPQDQ8Qxu1xvb5MbOJ1WhTklWncB3JHfpybx
DHxJhPCGsucJbXTYo9X4w5K149nVZkneiFc4QJsfWuqt0X9mxYBBp2aIYAtbkGPIj/kSYN+KOxSN
d4b23VBLKkMaI3jArMwDVrFYRt0Umllt0vYIULw9gOssWQfh0ljCro53sy+bi3bjkQjBu8kySpfK
Zor+wHVLI3H3cb6307qmkzO9wi187AbLTgMVdfTZ4feiDnDQ2qbanYMMPYnNeToUgTV1NjcTCCaW
C5RWWDP7Yi3lg8SXiny98O8YCleNkQTCt9UGlEFYAr6G4e7kNBKdysokeoo1WvYde+FfEqictACi
aNax0B0nlK9fANiyoM4Ku2uJfoieUYcSlRUnuAKSZgoCdTCrtoGmJKP2FW0F66drUwPR3tFX3aS7
LLitXktVibcEnklJgccpr2YCyRrqcYa3SIOpZt1GLrxg8ja/y4GgQbsHKrPT0Z83/DudqUTN3+1t
xuCCG+M11y0GMk8I4POjaxM9Knl58hlCMAn8EXj5Pp3wqcXmtVYi7m7PEkMbjNrKH+c2Gl+d40m6
RK2DcHmxi+i1E3cNZqB6KQcVtVCx5Vje1lc5P7boHmHOdlZNeGW6u4BR3FUoE/1cSkMPYHRUvitU
+59OAmbcGdAtTt7oXTkUzj505/akctkmVMS5xwic+iU8IZoSBGePbYRTxhFjkhRPgpgC4QLJAHDn
N2hBL5lcylx99ZB8uC0RYkxDBzDvzbAcr6bVl+beP3mgb9WB6Y1slDf0hpZb2hwumVbf9iO0YpGF
yiAqiNhrDM2AUUh/vd5iiBPsLpAubNY+gz8TuJjSHdu5ZppBp+VPGKd9VxLvwzfgwoYvGluZ9AlW
/cPQDiPztRSydT4BdrsMvHvXXqST9MAspf2/8pJVqt08iF4j3Haf0KAXy0SNslI8ltiWnJfafnoY
e6CqWZC83jPwVqElV4WYxyQvBe4LNnnqsTvhU1tZHU4fijIzXTlhsqXdyqSYzvTxKV9S6IG4eIep
Quiwp0CV7FGZnhUV0/wJZhfznBTijYeLL8BU1Mi6GqBb1sHoj6gi9U+kt1aWwpnoc9nQgmp7PGRl
Tul0NPlg/ylUROtOpuBbwiHi6/ZlRQB7AjQiyrEf6tjpjjO01zES9AHDrMNtiXlV7/GngE2iH4cN
BopBCusCpN/2y7k5oJt59J+w3rvYSEQAHR+uY3lnP7R/9OUwUSKqRqdjOC2jTThLviz/HucGYQat
sLMZsvozKHLIQ+A/TvxFI67O8Uiiy/T9AGwwazMNjEwrNgmY4lS+K/+ysji4FEb9yOuRb3LQF59Q
fklwy2LOIhgRQiadsx/5mkuJM6eXNFryOZzVkUeMrJxmk1iKIzW7jDc06vzVu1H2G54VSupSiV1Q
UTB+yol/apxVpwt+p220Uqa95oh6mKbo4D631+EYjw/EoYgozT23l4wBmXHishcols5gNEYH9i59
oiwwntG5FJ2QT6+lVykOjMPfblxv32oJK5aj/GCuM6Wd/7qmkm5K9nGUC9gc4ZvLNeJ45EEEDZmP
kIO1ywEfHNB2Xn2+SUmnDyxYUzo1i/GAqFNxdpBGhqViLVn8vVLznpN9aahkROfrMbkJW3WF2zuq
RgIqPEXEOVN0r1RK7iXASzGHSHYKPeaiEIpuRep4zuNoap2wSq4EEG4cJsqihsKzsfewxd+oj1Po
Cvrl9bRWCkyx0eCCvhWboe1Oy7k3Wh3i6vOcJ8H2Bwi5TyejSCISSICeyX/+8wyuRX+bnftJ85dA
uo6KnkUMiryVJamfw+sEhs5af2J5MlOkiRPWSU5opOdJZYsRpQbgLAXWUdyokN80TwjHOXqZtsII
gLDrToww1fPhOdFY2NBH9QaBAFBV9/L2b+urTCLaBJBj3xnLoxMs+3902TxPBRqGSsOAvc+Et9pG
XvsYb/4WEnz6znttK9Go+mtLNK4SjCyONJfyEAWyaaQAQFngGYUZ/ciOMxcCRhtJA8jv40jpzEMb
PQH+DP/EK+tg79vxhyUP2fbLPMITuEKnrEfbtuqQfWgSl5DP2IkM/ny4L5OGhPkQp57jwUZ0x26F
ErButNGgj72LhOkn07YiWSnaZK4d6cS6cxdCsoV6g9EtjG8shEc0x+/rqha8pjcBEnjHwwlRKOZO
8QHSUntmeQhxfLN8dCzTpFDQbIEk4CXJtPIMcdiK2n/6PiuYhD7AjV+Ep7XIzqTR9yNSmDLHMXG/
c+/JPIUbGWlZOc7crpemIb5gI3aI0TJSr6AuTuezvdCtUSpDUlXFUvbLo1ckcuJOyaAKvOM2j5ev
HaBh0Dco2lj9tewxvawLJKRXsr+d1WibK4R6ZhsQqTx0HJ4nGl2An/jUTArecNn05miR7AJhlR7G
fsUA0PTXdgbJx5wYlf6e5cBnKJ/fKo3TCkY83wmn+VY9wNkGWz76KgNdUEoAvzE1M+kNFsyOgHip
jYqDxR2Pi3bULeKcK+jfvgkI1f5aq2pVtZPM2dUXqxm2SWFMrzRr0Fv+8gmQDnLzKakNxfProHif
Q3ydAPgNWGdijV4KJxNU5y/ONCTkUkH0yhgNX2496efBIPCD6K6kETUs6ka/hqorHQFv2Y3aBoGM
JIjb9LZutLA/noZ+l3L2nqDHEC3388W89AReESrIFekm57wt0N42BfX9f43Cus1K8xFWT3GVzNtm
YZjkgfyRyEDvrOFnO9aUrhobHFyBHsQxlevi6hdHVTQAOy88QPTiPm7Sxfm4g2PgVpA8jpAG78Vv
Czjs339r/XKCVoHViNg+O2XVmB6fF3R7wwVf1uvHvBH6nWO8rbysWI5v5eG1hKW0SQPeQX0JilDr
62Fa4bo5ReemvbCUpjMsTADjCFNLLogwaF4+VWM0wkr72lwHY2m2vvUsoOmmF8voIEUTTJICbAPB
wkBexvDNB8DKlkd9TZ6UZTJtR+nlLFk1Hj7Qlb4g3fpOFUHqxPKZkT2m7he5yZcv4CV1HUbBKiYy
qFG2WFWTUMtu7g/FnXWHgLRzeGowEsG0JZiWhSdxMu9Qy6K/ZAvbxm/lA4dc1FoelpBi17njbt4d
tLzs4ng+Rz6vd4QHjRq3uV/dnVCgRihNsisk9AN8uhPJfmP3oUV82DLvX94OAIOY7+sao9+TLM47
MX8WggVitEh0a2//ETXnGoobm/wb1ebPiahtE+ZO1ulasqaaLAV10yYOfevQXxKhmMOJhS2yR1lN
/hClizqq4wJ3OfTo6++xX8ejPBWuhE0V/rwUaarn0vL38wNAMr3Q+u41xRSjVJMKk6A5LQzKO5eN
ccndWLdb+FgrV5tof6sOT1vc8qslAOV6TahstRbO1WUcoc1dHvx9G5CXMqVrfBm+gqA+sKm1kgzn
NR1Ga5LtlWlkv9QWwZaSjqOR+HOlX1QC70g0niLtjB/XkNjob4RQ7k5l2oZ3uqM9MBBto+1bmGXm
HTZUfuqlxHslblIw0K0ctnEskj3LbXapj2xMUQrT+OlRAIQJnC5PmUqzS4O1f7zjRtSmwoPxkuEo
6PkDZaALWmwo3055D5xE6SpLbnNAxpuoXHkbAGc7lKF+kqsrzGdfOYgJwzYBS+Qe9d68xSEdmDH5
IUN5h7vYADGhnZ5vtvk2H5Y+YEnJj/+5vCjPHjDJ1Kh8r6SnGzbuNth+hvPhWi3UIOjtCCzqk3gl
h7J8+8IF6oZZ9VyMcyNtFCAiwAyytYbpr9zt6n9cQbD2WVbVggdKq/FcJqsBGHuHhl6AG04LK1Gb
FVIRqDuZ5IusTBhkwkZpUTIe2q2e458Rd71Cz8IkaWKgKZR7m+5gH0EWfCcUiG7zGhRpxK2A41c0
+2JiBLwWyMajE1NVAO30oMhzlqfKIINUY9dXcFvoi+Aa7My9POmEXhZXBoZE4HyKl0Q1TPn9tnhX
A2+KhHbcEOwjX+RFC6i0wKd8Xqy9J/8V9Zh2F7zu2GXcKLc7onZiwRSLgzbmofaI+lOGYt4xM3R5
dColurHNOASgu1wS1Oh6n4Rls6Ky7O03xO9ATqaj8D48tCIGo/ZkeahTx3SFLy7ibSJoWClBv/QI
IzjRZycewzsS6q+4BYPzSAdeN7wVAkolTZG0L0YK3sywzYqhiJjvEI75QqjJnv2adQY4WhZSKDru
zJwEf0ZGfTuOBBa7Rnjc6w+xhLLplwH5wwy4pZEsbmixtgkFIzg3wSChsI36FjQ+HWpzIZbEzG+d
YsFXMrCmCaDiH8rNp+S9Ts69yXptJ6zU424sawe8gB5m0rN9A3H2ibDXt13Pa+yuV82jyukvTmCx
VC2zVeiDt/kKnII9m1+GdaPWd96IkPnxl0y4r2B0tV+mll4hUHsMn12nyJsB7Cwwnm3ceqCz1gfy
dqhlL0QAk8DZownD1DcYPFvjCQgUoRSXR8D+S31YyfHRDPxX/yFaDWEKLSjvJQkdjrBzFypg6Dtq
X0kx5WCpU9H+Ekc3T8PR08+8BRXCeKZxCNp+r/FYyExOjO3p4Cwd9Ey1FHo59zdwdKeZpEBJRsCK
QwdV1m+aOyAcyqcMU9c41aUKJkHvzC/4VkaJPhsrWTPGsS+72USHB6iR9ZyR5eyxZXKjkW+1kwYI
GHX/JLCFHDgMgwFeQzv7bnjN2BJfGGt7+XL34jB2DE9Xo5zHF1IP2sdigb99X8YTeQvDtmvgxDd6
Cc+5QpY5AbcoVE1QEj6kSDgi59YuNl6DVAILCBOM60/2Gd6GLVmdC9XwR/AuCogVYF+d7EG8/KMa
9DviJvPpX9sAALBeYlliBhlXV3FKYI++luN4dTqfPTfbWCFryc4/l1lxHtC5IjdaRiBCxACM9BzN
espQgnpcC9K06Z80YG8Bd+/5Jo7zQNlUYwezdna3UsKoaBV6nQabgLGcr8Sz+KvRutjfqtYv5x1r
Zh/WpGtYpPRFDfDGOL4WkhjEYN6By/28xhI7+DbS3fz/idgYnkhMCWY8qDMDvLYEPLntCXyMjrgN
uHzDcKLY+sOg5+ObGEv81dWgJsCBeMUfn+nmTT6z+nJBirT/BAPlj0pjPVuLlHFIqMmDNOGrjEbr
2xYI25OYTM2FwPOVBx1enjC9yxdkrXcF2RnfPO/frufV7EhH8Vwxi/MlA22KJ9XGM6KCrgdZ0rJz
7Qrm2MIMOLKDkDcCMo6u/+lIc76m0mPJJ1NTiZdVeZ5ssLKe3MbK1ykBk7O3ubfRKBJcdcDkOGcs
vCqZisXm3UA6H0lyqQw9Hegju42TPKXL0VebC6hDx9jQNUnpZEmxVsM4qDddBFLJxOcccXiPxhiQ
HcF1Nk4sNA84piF7bcU76Hs9ufvjLsfETFfpIt0wP2cb2heQ6C7vFMcol+nrYlaBHnj3gwzvMFr0
Jgfmit9Ogvsojw9BQ4UHhX1AOkbwVrK62sIe/RldN5wbBKFbq6hcCc4O5rDsCB191O8hUqrjsgiQ
4A2tsk8IIhOhT15wPQ/jNQ/NI/36cASZz+ygaSc7b6WmrsRkSQvPmuq0ipt9wa2muWAXDkppeoCM
exgGSHQjLkQvdsbkOhsiw1FNxT9PWnfFuk6gmKKiYbgad07zHpATixnk0fznpFdTQsAnn52bf1Il
C0sXTTLtO+Ryxobysctuu1GPiuHzAenRtsHhR6cJ0og/9fIdVWz/e6NBdgucnbrGiPDWhUu5coln
yKW2VhFH8RqqFaopLWPBq7CYUTQrbEgJJ0N7arDogX9LQBghoBfOtEjiVG6KH6KAZN483sVVEJXA
l7tpd4npINLTf8p/2099G4ZvRN1NPgLphHhqMck3GF8QdcFj1q21RMiqLLLUO9Sdh0ebY0g0z7Qj
7t2ZTgWQr1TML1GoWrsGWIZGMcev6Zkvda+15FMc+ENjzsUhlef6a7xv/7cXLL/YtIovtZQPk1K7
EcucPyUePl1KwIzonl66gh9ORdC46kZIPJJawo+0+NE7ggY/UQ3cB78z9kY5JowhmhHfxhQVgcGD
zY9e3qXWbpa86U+w9JI4f5RYG01rom8IC9Hvkje9lk/bjvU9pISoy2URsHVxfQZ0YlamUsJXe2Fy
IVxHQppJ7IlJ2QKxFe7GxDFPt2EJmRyau/Nr6omhQdFoNxr7rbhCzTdk6eE40ayi5i+1+IjXiFWl
+i9UsBgXuYhc1eMsOCRnNvNo5KknR3cyMdwhcPWs+IEgcvWkBprcuSNHPxqsPJoKSMGpqV3YO4h6
eO7vaD1yNS6mQmWKUv8w8j01G9ypEF+3DPHBcOqTr8MqMEbpRYrri362hjHoirG6lcc38FqINO2+
gQ/k3wAkQDOqfWWnhuudqtRe3Cknot+GP+mpqFuVDB7hIANUD+zWenFw2NROxivz6k6ZqmJA3f+u
qy7HoJ7cyyt96pbfM6y8Ytg5nyW2qkSX/Q82PvFQYsY9/UK6WoK57i1sYqHamjdHO8eDOAv0ne+o
gM2NtrOgnVCAMRpNp1ezhGXxyHv7KPAUPy/yGT+EsuC6FttLIP1n+enmcaGSt2HSOyihOAdHtbfI
CmAwnDTx3b4FcakUY6UsZy5P/rMZ95voehpmxH85I0ns0wHgTPf2P90WA9zI+0I08VYsHzEeMpQW
8JVvOvee++A8a6HCIvpp03FwkZuQjizMzMc75cmjT1KK+6WTdj7cR5Ck9PPuDKkKrinMcEtFxBSS
8F4GuP62hXtc078sXTWcDfZT+molnDCurW2zjVP1ZS+yQb13t89TN9BQf5Q1a90qDPQC6DS29Uhe
xU6LdQ23ZtJqKN4+uJ4Y1d21OCpNbYulszFrgNj7Zjbsz6OCcwiHTblPiqRkvxkgj23gpYmjlG+Q
AHvBlgScdOTFzxg8TEOZXcjTasKvluEpFhrEKmoa0XT3S3h2J3K2cGEymaE2LtOMmgGAhhGUkaZQ
jBb051wZk/tAEu0plSge5bsaeKe3GncORvBPxE5aSEtpwMPTWX/ovvQMnJBKoBdx+9KyR3ErvnbJ
sJcOkaKlOR2KIHyFT9F1wm0ThdQoZ0XWfeL4VbUiZ+NRDx+XnMKHb9MHPXUkQ+mOuFeXPS3Fi5ZZ
7UZh4AkRj8M+DRcTgh0U5dK5C0yUiLrqW6tzF/7oiNjhq9IotshTny25oyvmxk2NGaYA8Ewxjzbt
R3jxXt6A54Taq4z2AAhOPGUxdP9eaSsGB9MHKOUZUgeVWTH2kkkxItVTBynB0lygF/khyczBJsq0
7JvdrfB4vGjVKewYkKjO7IbEMXp+8W13Y/aQ+9X6s29VEWMc6LJ+OAsktEiLxdaX0vqO7lipiecB
emvVkwrPsxVMuOsVnvQt5HraVEU2VojtTS1MKP6fCe2N0mVERZfNy8QSkcjwyQ0zYEhsqOns6w43
lq0sJw8s7d/E0HtrIFrTRLaoTIRCFJ+YOswtPJcIysVR2kpsXnTn8DBle+q2Esqb0k7JaeaxaNV2
OPXt/XFC+ViWrML5+mVuoEUa0LMEerRhvFuclYnAvM5YW5uww8O3qlNndCc+YQwKMlqLytMPmCmI
n+7w5xsbvG0JYs91/+5n/0Ez4Yu4SHMx23tgvQmgebHh0GsVEH+Dh2ecZ7BN8IgNPrpNyX0/I3zR
hJS2TneC7L5aVnvDSXLWpooBk2MLlgg99I0QjDMU9q+GaKBqw1p/bwiFoOZG0qmELgmt+u5a7L0+
vptgKrNDXpaVFDvX9RtR3mFGblOjtbERRqKo581sDPCHSE4h9O2IDWXV2Fo3kBYRjynlpKrrJdm6
h2/DuVD5I7WenSIyZE7O4W5xAxmCR1qHwv7RGWXRdfHkBrRNXulWquk9SS0TrMl4pNMacO8HZGdM
xsNOlbD8eg+BZv1/gqvc5QGb5t1PH7lI2n/ntyI6V6yg8K1GBI9Da1Vs26RoVWKreOJVmKxJQpbs
R1j15ySh8lAmIRYWR7deYyw1b3zYEvkWZ4VOLetjbO039R9NT01Ej/59F9SxUbXoFdqUZ8vXgAlO
RIRR8MDW9APDEVqU3Ljsg8+sfGRjXCySzUOLDzNn9KYuqPN+alDvEx8zaQ6FSJBE59h2mvmtqxlv
0BX+K62rE2L71YJy228NySW3HCbvorlb49C7K9Ui8kh2VVptUE6E4QcGUynL4JQu/RBxGN+KJfRb
sT4YEtJUukndsLVQhDu0Bxf/z/bAdGAyZ0ws9Pz4JJK8Ghm1bp5sSVsNZC0kWaxtnM1nx6FHJ9Gp
fzbMj2I4rysj7TaH+EXnLSFX1qr3kEqU83Gs565zwK6cNGFR8Lx1bm96DTbNu11auTqv7Ye0TBfg
nz9IKosRT6xjVmejn98RGPvSchtaHYQ3bmD5CnFGw4ILY/wpEnNNcEWjhk1Qn80uyXmMdwApdLyg
d9LTPQdX9cya6MrbPztXvQMEK1x7u/X9UMUU8OkJ9zioYt2wGGbAG6gJd7dZ2FgDvgcQi+0i+M69
WRHFshEsfmPFJ7zlecBKF85hDqLAQKJsQ2GLsATOvZFQ5vAgNVagIfQkqgzfcTNXdMdYJzeDL+vF
2+66VfhW+5BpWr3tXl9hXoc4YRbozkAgQ0RyyrlZ4N9IXKuol7l5DlFeQQO7ZTMDrPfsxJ6x/MZD
SoqCEL9VLMDdRA8BPp9dFQAOik6HVNuPh/Eb5DR+mHHDTru3H3oTB5H6YJsYakHoPZd+Pb7YMLZ+
ti7wxRf5ZBLgtCAUTKQiGdT84deqeq1x15xddOb3zIEGYD0GS3ODiT7gIq8+zfqMWx5n5Wrk6cJQ
8TGAfq88or6Bz4DbehLMeYAMxRKOf7lSQ3GRwMlPBmzVso6y8xfp5QpiVP0l2uwqm8ZZu/hmvdr7
Bt4QhJwns1nnZ1qEoIQQ4N+aDFdvLc8/4ZQ56JhykOG0gru8S8sBOCB1Zj/reu216BWMlC4d39Ck
hXhsH3gYGP5iX6+i1At7AEt2xlO7KVHXUc72R1ig6dGSEghSZYoft7zOSAoXWeNyfwQ0PFqvty61
nloFJWcDQDgMBNDEk44Y932RPiST4/I7/lbcY+Q5LIiF7p/BtLBrWAGl1wYtIX9Hz1huBs++rcm4
vdUnD/wO3Y1OGYbTibEjizWu8PD09ZJkXqLpeopTzyqrP5vv4UpvRNFaC+UNnLUl7OKaqrPSGKIH
FaJRF5uth5QPeE7gZI/uDOsL8kwdW7QG7cxnmbabyRvqrEnZr0qzszTVcJe/0veTHNrPYdFKCSjq
Pkas/b/mewMvFun06KDqjTuL7inKgc+NiPf4NNdgYaUhdZSrnDZUGqwP5G//jOkT+7DJdgJdS5qh
PHFPfePHolc7oQBCx33O7MyP+ZJnXvKI+yv6K9XycsuygYqu9Vbrw/H/RPC6DBF7CXvHUqYRlUqt
evmwtEd0JRPBPKv1S0QQgiloFWnjBHElHwJit3q8T4tnJYTqo56tvGPyMNCNUZs7Xhrmlp5flInA
I6bVJu6I8nQohwV5B0eU4hzOi3jwl6Am5HfOvK3NTsqVihJ7oa6cjoMW314L7K9IsSiZ9WlbqXkT
AnTQR+3OQ9s90zBlJehxxLDGk/dhA6a5uGtwc/6Pw0N/Vb5PQYcmlJ2sbyI3jEcctikB/jDcbvIu
ypvR4PHFO7yNkuqTBvPGnl6wc68zfi6HamRKyVtTmR/xk+zMzS2Rf7OUXb1YAehp0xkv1f36V6hc
WzZCxft0e9oMywvks9XX+BaQOuB6ocIM4/WYgR7E/Zzssh9ywwQ7ZS2lyEdsvuDC3Fro+8z3R0tP
KsKmeyOHUeYD06D/5X3RtL8iXMEdnT/CaTIjmT/xt/hlASIu2Q7O7F4sZuIEjMruCWluiofKVxK6
lzFm4ECjZ7oTCEs3+kq+IzSUQ2olYupDNjqkxLgj2lsnSQCq22UegQQlSXPHejLGSutvLFutrqqj
98QhwKu05RXUhir9uia2DlU1esoEXL8BFn5J0ErQvNvWoI3Z43tddXKWU1YPxoMRSPfnHP13tacf
gKwcjF88ZVMrwS6YTGG/ydyjspkvz7Muq3WGwNi9ePx6AGAWt6u4pCvajRh9bc/PfNsZ/jsJNAAl
ybg89xHdhKecm5lg+Kpn6DUiHkkUwxUkiuXl8M8Dgw0OPFsQmBynV2hvzOyndzrCzKoPGP+Pek1M
lJkjD2UI7hgj/noWrMduHoDe0NINx62lt6zOgDzdGkohD4TUhHGKrC2RxQDRZGPJepBkzWlcK0to
nUJSJ5fU4zDlxjt35XwT54LoCtV4lYPdvZGJRCVJWmGUCBl6s6CAzZ7/Bt0sII3Y8dwJ1/XZ9XN9
3kKFcLLcmryuzMBk2wfxyDHtKorXAXFLQ2Ax36btdX/GpU9zwYEWg8xTYV8FhqyoN30Q0WnXXvye
Yhj6crtFk/ml2cQoagg0q1kNLAwyzHZCQQo28q8/z7uJBs5gOUJk97BgCW/HkOUBileYBpEOCLV0
Q7lzy5v25MpCTXWQ59s+h6coB3SGMN60L57xyuIk44Em+9c1ie8KFu+RqVx8/fIfVQq+l5Xm6R/4
07zHFOASJM/cf1GeajootKsxKlDAgLl6orK43zx0u0g7XBPV9fCZ1EXEvWG0jgXcA5rFBFK27/Sm
pZ2BS+aU6SzUYqOAwglxBh+bppu+sx+0d4S/4U4Ky/KoqTMQJ5RFeb8OyA46eYdmnPnYqfO626+6
+l9gXuQVXZXKYplDEY7t3qOst8571Rvn3bsD8LGpv6s6Z5ym3bhbPmQN5HbCfqbVQeEz3qi0m85C
iLw8XsLNs9eEZ+8yhkL1tlIabHAS/Kx0xdiJMa2+x3FBGzzGkT9rx8FRCaeGbixvg5eSzOaCfPFb
bwBdRUQ6VVxsr42qE+v62UGwRPLi5pvC8CSt+YKaBp1Hbrfm1kSF17y4b/+b/kVagwZeRTwP1TP1
oLeMNOwP0MYIsKuyIEJ2kGLEv3rObPdr0SaBEBvONCMXQHnYxVTBijtfI3Wm5PLM6wIw7dyRY1wu
onA/ph+woXXw0fO+DLkKBKYFuTCVeyLkfjRZOQYaG4qJZysYH3mC7cg3TkIGBIRvnOaFLlnjcMTq
LilQLwluKToYprC681EayWGHgBydhNLQx2Cj5T/bzpW1DEQ2AHnNIWunl0Xtg2aN9DofRATWFD+T
UDdMre6HyzziQypKh86luZySqbqanESGHAFkTBH0J+NttAQ0iRxl9zltkXX+2Plj8TojzSdczaZX
Dktb6eOtpp7M0JCXBV5N9086ZtjfL4HUYNRAUO7T0iSb6N7IE6KSJQ4B3lZIJiFal3TIzrKNFy0U
+0cNUniFX29H5OWh1szu4PxspizVUSwlx5O0DgDYgS0XTHwXtUdQEGxG6ENovqUxoPwK5CfKuShy
EwJj+/9zy02w4I+NV2cHaemvvV2VQGz8XTvfxh3n5hm8goSaMC7vHtcl3cq3nK4OHVN/jdc9ODxY
HOx/xE3WT5TTY8HuFh/ewVxtqEs9Qx3UCsGyr/FQx+4aY2voOWqcYfWEN/NabVei3PtRzvdhMC0O
bKieI7xpugXvo4PUwZZds3bSBulYsj+IbYgSAs7BnsHK9ATXEqa+VrgKqdEopKfOvZMPJze5VTKo
nxPX5j465aDZJhlDAuU1yuEjKz80epHXHtkUcTUNO7Ms5aolqY6DZmLsmBggSq3/p98+vXBN1Blt
CEl/BGGhsXMY1kca+Za8E+Sg34UKQQX356fxc3ZI9GWzrVy1eXx8vKvLIXpYqtgnSpdKkLJbYVnr
HoUL5gAD0KfF2jve5ZMi8yesvRKTuE2MkL+GpOilJfX/A6HgAdfu31Qobr21s0v09EZhqzapIOHh
RR8LrFRh/eNMwFBn8o4H5tE17gSBiavxnEK3AJYJxO10JETV3R65vqgfgkAWzV6zQZg+x2rO1nYL
r0XnWTNFFVF7z9C8JrWZk6Pf3GVsZqCd52suv0cVLD4ne/898do4Sa10qrafCHRZ0ih4LBN/OE5r
XJPWirkfSE+36yy+4Jkio6cMOR4qG501BFaDM+4ybOgQalRyE9ZiiMmJwN/h1ujzB2Q0HBilhs5O
lQzkM2SONqgfF27yBxRr189ovPyLBMr3DmfR/QqefSK90Q5jBDhvm27I4hQXPDN8JVLf0HiDowCn
XO3T98fEF7xjQn+RmLf9Xgzjt7wftQV/cJx34xNz75MAuqHmyEy67ojgGoTMIylQtSoD/y8OBx4/
Ahhjei/asAF/G4YvQFkxJpwck3afDWdbQ3V7UUyUdycpp9LtMiSJV3os0itSeIEuwRmGFNoIgl3u
TbboM+P6KDAdutMzXEjACZEBtjuu2SY0Ya8oDfg6F9LzWdLhtOG7rxLG5Y4Mpj+tQwuq+Umq6efW
TGuIRz/9U9iafNrspCdgbwyBnfn+/i1muBhQ7HliTRDg9wLyOyoEtVXspFoszpJPKE2tZbZkaF/2
MLIcpH0muxh/vkgl7KVpgvdRkrWY3yE0flzOHfzb+kkTPsKTGiIx8LNQxdi5br/l8vCZdNIe53ae
Aldih7UpwWgbj0B/wUGzYEbs06WEhKaDiP1MfZmStP7dJWcdYksyqMuPwO0G/wZHFoig841kPeYr
FzWDAkoKnySNIUUCo3xl0l+Lqctcj3PJTl243+X67zY06UtoOvmjSkLESFctF8IBkkY6Fo4SzY1U
6uawOepBSJO2LherClJYDfuZNCM98GF1Oa2Wi/7t6Wqq0ooCxFFoEYQsWoGIUkOaw7Fiqmu9+l3z
fDUTQZXGZVuiq3UfszdR4y1N0QXA1eNaQia3FV3oEi8v+hS/XYgNWj6zIK/PyZm4lappvPyH7VVK
+HRwg/TCuZZ+gDD81AFxN4kooNgYbZSxyK8PblGI00VMobp4+6dE/Lg/ITnB6wp6eRN1zFUveT6p
InLSVsAZUOaNq0YDhq7KnvX/K8BpvZ8UNenTeaac2ZfcdvO4bzN853smCaau1UtYXiGB9vOLR9gj
OWgwZGqrToUsEcVyQ40a1eaiRdZR9K18PRZTzCZbP4f1+Wa1veU3kbO3QBsTJUcqr5T8dVf0SfmM
WXsRbkrMpzyLBHXbr49jJ2x1C3OsLsN9YSFU+G2VM94KQI/UjdOCd1eCR8xymnfnMv3Ugy4/PRUo
FD+TV4xjE8Te/FvBjODB1ED9G07i7O3lGzIT7EFyyNTRmK32Tuf7QpDWVME5WXoF3NTRBAqoCwhG
V+zK4itn77vR7cmR8FprfhX3ykT24VFYaM6t3/YgWzj/2eOKv2b99fdU+Vx9C9osSXqOZUohhlEL
N2/1Ak1VgUkX4zRwyRl/Mo1EBYN6FVKi8lfczBu54ZbNek1YOaPAFcM+eTxGNIR2/RHIKyAoDsJ8
80CfWaLOjaCYKc/CfrKTuNexOgAuB9mNXU/iKsv83GTc2ZvD+lL0rQnsyfiuQcFnAzK+gBcaGIiN
KiXR4lenuXIfiQvWoQrmYqQfQ1np4Jj4sewSnFcdbNZ4bhGwD+NLggpHh5T2aKa+ok57zn3rZQ+4
sTEYuJQDNy7PKt8E+74wrExnQEj6G9b13S8XX2VgyEt1pbVk3/M2t+Us0ldi3TsliVs0uYj0PEgo
malGp1hBoX2Yri9bIk8eybP6891VKnI+x+Nld5hbHIfhpJChMSCINLavi/IS4hkjL5za4abhdUGC
bIC2AwnRBvFckG8HFd8w1eR+ZRCBLYyju25MtymYz1H+tb1ezwbEpBoZeoSIwVjaZeqDze/334x8
JW3fVim1L91qt51svGLxKcJwF1VasYuVkiN3VbZRBPplovQ2zilOHx4zz+GxrZ/ZGjoIJvO2504+
WKAyG9xv2d48sW2MbhujIENOfgIbTfybPlBQTJYaBNE/R0wHi57NhczxvmQork8lb5sP9IzUjhwC
foYTu2Wz6/JCOBWFuda4i6aeRfkKt+fMyD1zZIdedBxWjN0iPX10EVVXxm5n9EY/v9PbzzvL1cT1
aPMYVPFJT0Pf5wwdmGbeCv9P5JGjJzAy72Y6RoIbcsXsJ/DRgrBnqULkn6QeZx47txQPEEFLCcaJ
eOhZqL0ktjkML7zdikT4/R5eY2kKspRCt6IdtyHM0o236oEr5QXrps5bESVniXIjoR2lHoIFvdut
TAIjQWDpRg22tzxEkRFA10B4zn2o6+oVKwy0MID9veeRowrwWvfJiVqD3wqrXkwLlywTYLVp3V4l
lVC5r45MzTqsww1vCRvYSr4FA+NkatgKviML3ZWZE3vm8ydR0VQJHjYCz/nR32E1I2y0zyDExJSC
1I+G50n20ac9HTrfiPs+0OyJhVUEmpAAdMml247lZkHJMt5/mvPP1Jfn8s6W+FdRFRDwK1YuJJOr
uCBYoCQqq9wu9rfvSMaxAfCylcTvFHERrtBBSTCUSF61bRTl40DD88nHexaSnj31rvC8EnAbajuK
ylqo2VB18VtzsVhwOBN3J571ZLw2Pic99j8Du7LIzFLEr1tgsyTfKNKoZumWmEzjBuOUQRlSRHm1
tzWVkN2PUtzTCutidcAPDz+gt2f4BxgsdomKDWcI2rEgWFLpfWwLVaEM+Fy26/g8JRNyj0dgqxGN
i0T1uMZEekt2/dntGhX4NzvIz9xLWrUARgwdEg5OF6MerptluTDEHsxikrtgljlbjO70bCVT1kvQ
4oYNi0jd1Y4zvCpT3Qui5YbyFPDx8tWFdAcMZFQKwH41H82hleCa3LNLT9c8zXLXagzV71+X2J4p
Epf0cgZsYzdb7iJoctJROj4S800m4zH7WzaWlYBgwvNxKOXIpsHk4AGCMYfNB/0ALGj0f+TlRYYn
G8Ji/EPXoU00jBMuAbzPMsKCKPAUVYTX0/CYf6JKaJY9AUl9nskGu8F/tJtLqD6fMLGy34UDc7sN
xqFMD9Df7LY0myerBs7JJ0spUjwSLWeUz8ySnJxou7RxrPQ0ftNwQttxij8daAyJHitRFyP/wm4Z
Dp6DPxPjGpaFho89WQFeMy7ryBb9jlD4/A1/xm6dxonuKAaYmG6iuM8uRShAng42Ch6c+oV5z1AW
RsSgvEbx9gp0y4HxcZhlDSK/X2TIp3Drh7sl8y+5wIJPNR/IArqmxWkII0EoiOWYPMShKGrNAG04
m4Eg+SX97x1kVjtoCEiR49WdDeWhh3eU5CUSEm/RBpT7LLtCB2IPGFTpvoDqsKXwLNhttjrr0AFw
fVgdaViYYzM451nEnGkRXgr/n1OgekpIMc/bc/ot6RXz8mnPd29e4m2Ycti3/A12uvFgr+ccl6Re
Fr67YoqEnFFSxOPwoDpWx4zU0M7F6iY9YK2Me2egS3F54rKmB3HspKv1ueFHtFzfnlKccqE+V5mM
+2WY0/VmH+zd0ccHiN4RRGbkwHp+WxfEpwGN4B7DmCzjIjTbUUOlbhaCrv/TIfOiHMqgK6LLuNoX
MVqigKsrWVnEmcYIZuL+G/W0RgoHorihDk7erH00HgZzie5Z9n/DDen2QAjzW0wvAjfoi2JrjjcN
NyngC8aV8+Hv5QL2mRhQwhlWmUtJwcbby8hvF0Tbs8ojBWMLtsxyYdDjged8EssqtKXDWPm6ciHk
zfA9RgkQAjqvp4SvfVDqEd0IHJviWftVwJrYrEL7yTWZY0OnmUn+CQrf9IffSUNE83/s+qw/S3Dh
4PKgdW2NFbdQEQkpaK3lelaJFHTQlfIJHIYxnZnKfvxEHY1ETFPfRI568cDy0LpJ4piuTmS+SXWr
N3nI7/Jha0G68EWVqiKcc0RhpJLt/VTl/R938Qv0NHiZwV/QoaHgVTjaPnwhU/as/edL1OV6bUoG
TRyYiIZ+/tJsaAHecebM6Ol58hQVi0cEyOd5NJu+dapX3CPupt2zI3sG2OIpg3OF77AswGVm1ZyP
IHxlfPAkxGPvKCJS094AoIZ5gGh915C88Cui6KwN53FQ48V9jpEgsIn/ap/ibpb61y69wps5grTr
6C9s1O7zDhN54b/04PqY1LDMNMIwIDUvcYo+yqMYaYrDKrK2R4NO49cMZ6o/r+pKU7f+9MoTumaY
J6PBzIrOBU9FADHlprKfc6X5aqtxBUVezgiUpAIckqJYFzA+X13MeAXRsBc7MNQLAOjjhXFb5cRY
uBBV3rEj0Z9JGpAOGNomBGYOMNtkhgd4pavWadWYVVt4bj+TRtOinYOxq0gt9PqN4lpzB3E8iJl7
LqgHWu6ob/dclLJEgz1ZdViZMvdpA/SOhhoaXKMeqn21ufCYFIuHNS0vhBjUWITeR+lMKGP7evA5
HBsPwapZPem5l8NKEMkm2YPJWyXKP17vwACGp4DLgvpm6VjDb1ZrA1ObZYCFtSUE59QRpKQ9eGJX
QRS/5UNDdO8RJl280+Td/6WgwoXMwqNhRMV4ur6fo36GIl+UasgEdZRqVZjROq6kio+xuK4XS9OD
2OdkcNmEfoOhXmQA6y4644CHAwvHZD5LyHyHGul5XfZsk8HGC25VkGCO0ArCwN776Gc3M8ble+dh
gHfrCeQ7H/ULqRe4PumVadmbbqL654sNTm2B2AqCXLibAw8wcdmBJ/mhOHYmY5dbzrl60r5ODb6u
ZXSoijnGrrK1ffW6IL0gezTeD2W+6/FaMnH8bILAhtekCPRt0NAnT3L8msWTajkayfrwXj/hGuUt
94gzZKiuwzfUOtK7HL29zOBWTiF/jegxpFnYxWipozbmNdCJOoeKzRlq7KWom0yomk8gU5xgKa8X
MpO00Cxrphmtex7J74Zp4R3AZwswEXUr59HpjgcGxBb99WBQ7338tDdX/xjlJSlocl1Yl6DHVkik
fCfIwDxwXbeN9qoo/gx8iCrzWtW+wQybZxap3Tkd6/W27B9ouYNHz5Y2rLYrxFTudfQIqQNey3Nt
MYTBVUoxwMIClvYKD1g/2edQphe4AJ0jNYBc5gHrAopmy+7xtX9+nS6OcuBlhZjkms/y27Fxrc9e
0uwspxHCTq7l0I6aZ9aWFO66XclTORpiQqOcEG6s5s50BF4qhbp3YUfe2uARbatciNqRhPIwJdIk
a7bHo71aJiCYZ02zk48c4h+hyppMBmxmWX/dGEfM2/jd3T3l0baPWzYOMR1gRL8lia9R8hGJ5eKV
bFn7xNvqHTFqTU5aQcFx/snz1hNcRXffx37JoXZ86UyhpMkd7EaK2bgwSJBZdxZEqipultHDC8x0
GEOkbtYpbE9098VFoHnBGTksrifNrNtaA/wtvW9WDj/Au2I18kMsIDOriHqhfInGJWADDcAOFFI0
2UyN50RII/52NPcXuLTU4IB5G+Dq0wDFjIxyoOmvYvVs0l/drLU5QQzekd32uVqSAw29eDi6AUJ4
wi8RUhzW3mYcPhUv7k96oDr20tjc2XYnhcjRrjdkVkJ2vKrTnpADSGXim5bms9VvUj9TgUmVWqWb
M9bVEFa4IQqwk6KC78/EFyreOD9PeqBL4iNReCJBO9ZOcmFgNCaSxQNg6FTTtBKz1rdw58Okuqiu
haff5K5RL7+fVX/WrLEEM0yOULQCIS+S6zvZR6bkCPpoTrDzQcANc2WyV3n3W5eO1h7qVr2L2P+R
Y49X1oZcbh6xFI5rmTzgGxl4Xs6fnGnQdJPguiiS8GbjZ13wHyqwv9jl7YG1/owwueBGIIaV9VEG
nMTdMtGhjfG8PpD4Bdq+b/a8GrSmz22UbilmhjLlZXqDBUvUFsmNOJuHNbMv0koy3kNNpdNlw5VA
ipFlTdc5TACLERj/ZsviOBHzG/XFR1NhV/gs+kog9N1eBxwBKccC43MSv69iXm1SsIbrUEHVMTLZ
PyOA1ZTEwtPVOcxpoMY4zTNgdkcURIHb07MX01eku1M8rI203nXdznHi7llU9Yw1dQwpiVoZjo4p
Pg2YoyJStPDIKke3890lYF6nhK0e8epvvmO93Z3xoul7VbAeA5J/dS30jgPbYqpNnKnRHiGaUffS
6V3lNMgddwuxwzsDclaNtaMEUabgHgeNkefxYXXOYGdy9Ktn0I2UNRLv1/kCsvzKd5KPnKwQJCFq
J0DSKes/0Td7UGbWZwItLm0f8QDUO6eddXuXcq6HRHDXh5AZZXwJVTecusgspK+tOgqw0MssYDQn
q+RsctFXw0WXOm9V0vc410kT/7/RP1AVa6tZMD4/j1EXvc3DDHz8yjbfK5lP9vfxvT9fySbTsZiU
OrgXc10uaraf4H0LMK4J1saPOTm6+LB2dGXEmfpfzQ09dbr1ZvHPubl5WZu9xIFvaGUOknxxnwd7
PBk1dD+R8vTaiznh8ZQCihqE0+ZsQRTpE2yHuIKnX3cfy37Cc4CIFqUJFsPbQnSuHhrcADo98hEL
8X5UE/NPbqt8COnSC1VAVVjH3+Ec44i/66DfOoP5WC3ulbQILuiRoh+3bSwybe1w27uYSHX2nF/Q
L0fceh807nnmFTleSNuo0f3rUcs2BqH6L5P6fKrhcaTmMeqkBF8cdt01xjm1+pk7pf/oxxUcuavT
ysq8lw43fFxP/DR6OISo1yrm3O7tEF9soCaAmWQ0xi4wtT0Q2DAR2YHvnvzPfaG8diO2QxSsGfC2
lfVCdI1frZoAjd5p6RfJtKguYsAgMXa7UGn0DgN1ID1uL6dc2rrDiIf49aFI0jKzQcECtj5HPF16
+iFKTwIomyF9ogyT5uaybvYQ9VgOghUfLom1WlQXwH9O3rG8qF/m2rcYZar042NDiT+X4f4Ep6zE
1sWdY6ppvpHRCXUtU27kYwhrMTyrf0i9youc6RpgvDxh0igyAllmG8c/rEicK2FIiTlC3v7LJxFj
HtdHz5x2TOQCj84WoMIo0vRGml1xJTRty6O7nyv4Fcn1+cXJVRKVzxN2lZqod7heCWU6T2K7odw/
lSWmTPedSUHM9g3C5odiULsDllvmnvewqytKwWfHrFIZTV8=
`protect end_protected
