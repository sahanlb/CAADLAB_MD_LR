-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PGFY4a+sBYxslj9eLWlhFgvaQKQYHdp1qXEBmfRpXbsGpDpVwLoSgXPLTkHtjoVq1Rck4LLMGM0R
Qd6sqQdUaSY9fF+yfCttsMSAks75dh0Ks0iSOGq65zy9V3dsTHFRpV/iHea9tKXDgrJ5EBA5UJJB
ONY27CwOG2Y6EZVhDI9NS9S5FKEgyym4Rp+qSN6A78mBeecq0Gj0io4VIh7hfSNstRiXccdawG3C
hcD5bOH+d8hAdLWiu7RGBaPmJUrkq66ZJASjhXx9VNLc+24oiDJdJJjCROq71IHi6uEGKuUIFpZN
bU7MwOv7dUNu5H4Mj5SXVhRH/4YgEIPLdw1Qlw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
qhRPI2JG07ENAaGTudbGftozAFE+TRlNOC2c9027H7jrS9butMWBBGeDUx4oU7gt672jABxPNQ3v
7ApxnNazpDQNpEeF0Kr964XnvtJlNAXfMtOeLJrCkSBoFjgBpIuIjA0psO7UMtt9JwEFNEa1E8hb
qGXcflfVOYjvtMDxvKof/EXBuZJnjnMfok7LL2QpiNgjNyS0E/cmoDRYcIkcXc5bJxwfrapFz72I
I9sKFN8na1U51wzIIvlTtd5QKo5e/2Y2NbUMS9h75Plzq5611z/JWF6Q2rYDXbx6Rj3o6zuJR6fa
X3DBtAFRZtOqDB8UkV0a1efnjOF43bfjwfZQREfaU+WulRGt6RdRMLuT50hPaqOnViUZ/Y6qXp23
D2C3h3sCQ/dJ80OKdZ7xvYI+KCtWDCGvdMv5ThXbinIJjil4FHgUAAYzNzzzSaqoil7mJ8y1bfxQ
2fSWp65XamSkgz4cH6/oaSN4D7MmJKxuWR3o0Z4Gsn8e5lrR0wh0YinCPB7JeYKtHFEP7QxXLUNE
qjBwDvSHhmXLwzE4R/a2RAQMB+vFL3tfmwY5W81Nz0ndrXEjIkaKJsiqrBosC8WiONA/tfauHF+2
PdYrwPGYqveoriGU6mhtJDU04RzVTzmwyKbTJS5NukKx2MRDiBLpxVSNQmgGwGtTZKPjTjcNkOE4
LXIGQDsCZMizpmCkweGQWVvVSkpWQy5rmcjLMOb74RUVbGBl/EU712lXzpXL9RR0Fy7HzO67eslu
y1BLhm8zTaZozwY0P8oEFVOH/iwGqup1Ejcq+uf2bfbiBmju6TC2BVB7YPHkIWuRL/jn8aDP4nu9
v6fsqCJMzqBV67ZHTfiA/i7QyzL52HbwYbgtIIvROSXOPC1gIWjWfocBpcA+oZVrFyFZcexJS7u9
PD1jCDm0G0w+OG2xoZcMVkpuHjTN0anKsZggL7YaG68i0xxAikEfgLZxJoSWV2xb4MREuMuM4TwQ
F1DORIVpiCKZSlwWudY6EJ8fqfw3AwrtqifmBXZ4xvJr7AylyvRWmzso95vW6uaP2JuuuvhZp9n9
EM3v5iWMfrTU34OaPdJADfrVAc3npJmZ2/SaoM2ZEY9E3zCfzpgnkxiQKgVuqU9EOXzgnBCG2fE5
INo4tREM/ompLsI/N7lzP6GwMZQEV7zw4G3s0z8KvVXoKvSBScmMdaZRRje3GnKSaBNjai/w8qOM
xi+kXoE/7UYkekdmim4rhW7//VDSxg4EqUmOKx/FLNnRnOMMs77GeIOicBXE0oDtsHpPSrqpSzkh
o7MULpvDfO9NG569QPr12sGH2eJMQOilZGwufvDk0czM4xmA/00Y4VUb14TrX8y1Qc2NtUNl+JK4
/3mMXBjRCwN78mopSw+KGpgTl0AZyxYlTEq+GzYXM8OXi3Z3bPVFGAKkZStPQPlZgzAQeXX6p6ca
yQAZ0FILm/2eD2wklL7VvauFrAnUagwIlrMtdTPrfIDm1/mxFqQjFjPtJazQcbsb0AkAWwpQF1Iz
0f29zRKB63oGGHqlB6OehWEBo7/69CZX6jlXqq45hLfDLiZd1VFd/lUXFBci9fqGK0HcZZo0h2Yy
mW8Y0w2TUKbIf34o8HOK6DFWM/oYMcQJ7WoxXn50S2jqSMfWA4VA5nV1DjWLrZ3qqoHMezTwtWZq
+zoz8aN+BH5hLWl0XR8jfdy54eR1FQ1vYWpQPNjKDtZdXdOXjc6n56N98isdvwerdSR2RNcMfMuR
AgAmKnQCL9r01gOYHmSzMHOCxP4HlOENB33geeQrdHURcXk8FvtIi4CUHRuw5Vfhz4+6gunSRW3z
SydAARiMslWTPYH1P0qiIMsm38nIOIkBAzWlkaoX9PMvr+/NeX5mHx+lT4X6itT5cxaurVSOt5vg
LaKqLQfjTTEGOUXC8uOyH7bqWjN0YXKWp55sfKsWh1UZg97Ky+otrcbtoEILChJGK2XlD9ADKGsQ
HFpDes37k+DhLMENZdvEzlgIp2KO4ZXKHKb2iX5A1SECCEVL+fhUF8wAsCc5tc3/6a3TWoSmkwaC
TTOY3GAden/BjwWXLpEsXYj/dJ5yRD2iDCUZCWUMjwk7u57mEHshhtbErZKXsMQEFIolyNXrWdo7
biXSlmRMNHjQHQPIz2ypr/diQeRsRCvbZmbafIPVWQ4bvohvqXssHGc/AnUrVYwk2krmh+3Gl1NQ
CD3u8vCzL13K+hrVxr9QsYUgnxvYbvUhRRvSe9EVSFHnvn34OAU3VKaHTsJxRS/u5baz2VAW9hWt
X0yanjJKsQmMwd4vt/HgYy7K15FPAvnbkG7Kuh2/vbxFL+bJMoPs6x4ktIrXf4UFNDLD8B6je4gG
Ib6GxgCsvDtt2NniUtXxN8vgX9w5LuS1uyWtJJb+PrP/XgX6g2iI3v4oM/YEV0fLce4flScA1kWw
+0JAKN3Gf6GRz1YRegdrpEZ0wKson3CGMhUos/epZXzFZcbOqepjAoddKgkydDVHCuAaAgq+g3F3
ohuRBBA/enOdD8y+jWJFK58RhB0OjbCY3O2uVxrFetycaaZLkY3ya5R8ujIZqRKuWzDEx2TMIkTs
naWFuC9TdXIW3ETPFigfs/vusg453Wbo4L1rQZpx4Sxefxc6fMVGz6IzRRetMYK8zjGjVsbvsO4K
Xn+eIxEGi6umXgX3JK+nwW/VqnutwEfzxkPFjs4pXwyvhIJ+ukU4qClICeS3VOsFhr8pvJnpNPz9
Eql6vz4uqm4Q0Jqo/Uob4VWHsMs42yO6QyAodVhe+RsK8KWpW1A6XGlkFs2Mb0KGVZPH2JxLX5nK
k7dOw9sQWbJcVW4eyeqTLhix20bnRTRlkURAUTBGM5awC3zG00BVYrvYiRQ2fw/FK138rEbDJrKh
tfLVZaYYY4UZ+UDQ/NfUGLmkOqhGdjuc0B51Opr97rf3PSpSOVG/Yg7r218I41AixpnQEjHk+S6n
tyiRhowjpBFce+AEewXtMMx8zMyEYhxuotM8idyU3v5lVKM47RHowmb3+plj0JToK9LhSzT8s7h6
iWhc1EcUZ7O8aU1f9fGuvK3QllKr+YdK7IQfEIxAEiolmhYXht6yt/1na6YH7XZ948v0Hr/JFzmQ
AKZeCvwAmDOyU0JeqhHEDB5kGRJOoMN4u7f/8dnjraiO86Lh+0DSACxmYKZjUcd2kVKgKyxuvm7M
B4AgaUWwOTMiQUH3b0shqYhWqwxkO4iHstEopQFNHM2b6I7z2TQkccDM8xtdh1T4IPIrq5kCEbOc
B0lf1JwUdlApYiypdvvPreeNiSIxy0CBK2Sa6KvyqyMx5KY1ESx3tTDpyAJssKMYoNjDvRHOFWoV
j8uMqMmCAbjZI9ypHD9UL8qdy6QbzhdOWBO9pcqS1b/j+gg1jo7QJH+UZRv0NFEE7C7AeIJzMlJ2
360eFzcTS9ObpWrrQXxisQTPD7UU0dnJ441uKi2udgr2twvsQZm5rjgE7K55d9K1Nr/rGtr5o3aY
pX1evu3HeRNH4HMhHd2cd7tX0FblWxpqPNlzIBkZvc+740NJbxUyjYjk5f981PVPy2/PV+i6PwXd
v8mWsVNhGHv/7GtYavKwPmbdzxmcU2NydrArO3mx5Xb63lvqocU06mbHPKz5Hqg2jdL+o1Nj7vCR
XAZWu5d8ylK+ZWRTNp5Hh9ZkBIwW3Zv17B/qGy6YerlahE4mGsMGqFarWqPNFRciH+Hjbitdyt1n
v58IRxhJlknMdmR3EYXWfskr6JClwZ3tmlv+kPGaty2/zsteUyJoXEDWyGoV1cLXkeHG8MnxVOE3
/9F/afr6f0hPGuISrWEzmCcATwptH/q+gED7wdgj3y6LDF5HWMepCzl87WyvOJBYm3TvM6ktyf4k
9LeobHzI1peZjuUOtc9leHr9o7UFL02K2BgnlRcMpF1v/uwVYmFMAwJZIwCDOHfccBFB5LtiQACU
UclVxjfUJPDpUolryYlY9E4IY1EKz5aGoaD04nvyyOX+mR+1X/1DFff33VJuw2nYfeBW+BvPEweU
VXnXKOp7wW8971dJQ0RcmoTTPwymkp8Em25LX60famQhy/petVRY4Yub3+VYCySVI0xf3c0Z7qXX
2QCmwX8FmwKFzyibJlwfVBU5ZxuD693B2nYZ478+7IHU81h2LL+4mWXw9i9Tode3cMp1HsbMT8dK
BRtyTz5bW4OShNg9ypB3hcLwFBCVltcaNPWk6ED2rthPO6MguL4LxiFPqT2rEmUZZij4wGE8sM8g
zAxJio76JOXemhAMJ0KNGQ0qoAhpycQw9ynYtI/SwQL1yONDxdWhKXQbnRQca3oM9zyHeRKoPExt
WG3KL5by8aqSO/XX9N442bw68GFxBTa97nzAjqetD3nXQ5cz+p1b1d2STcp6+dTMbrw+3dQ/ENrJ
uOmqL/mu5Sa8e5YBwE60PKisbOk3P7BFMNY+/+MhvEQOVkg6rmwc7WE/NZPRFGjUoCb2+mBCtRj9
YILHXk64YITWdfxUnct7HCOmWW/yMHRYcHczsrTKrhMqXDjttL7dXtg5lfhoXRTXWd8sNXewXaGG
MmyBuqXIxS8+3Zx2wZPXvojXz4bxlrDJczVB8gpSM2EXAebArFILhbGYzD2FGRCrxeRNj71BXJhs
Q/C6tNkdGYAKIruaEijwDvQ5o3+kCpb/BgHfdUhxCpHpc7SYG5YkvwFIFn8SJpTl8rkhXZCvtki3
o6Zk7Ok5IOgvZtho1FrfpGvgIE7v64cEVrTs43NX2sHyGSPJjf/re5LqZGsMkz5IzWk1V1VAz5ET
2SkCneFSdvYkHstHuiwJZIkdwmVVaLwMv9FngUnnlPpGaQk0/KhkcN9zLiAdlUjyVhOuIhToEVeX
XWPbr3IaAqQmoNoH2+YLK/QiWWRXKB5Hkj9Xxr96MUkPbM4EIhN5Rvvha+osDsnTunLfclCtd42R
E0Pd9WAsswE48X/9QLWTHHKUnyleTm/XQ6B6HMbZquwhduqqi9dNgBVGV1n9Ig8su9445E/tHb4l
CKQk+87KP4cxl0XTBs5vOmhWXKxVxDnxcPXxTm7tmmZ/lB6V08UI3X6fqq8SqYn5XY6unE5rHcxa
CWMi4tr44IZPaA3b5YHFvM1QgUM5cdsaTigdEfqB1ogMV+dRyarZL/3FHbB0keWZ5G4Y2o18yqMS
AO0YekM0t+7nCSbAEzRJWezITLck7N7oayUG0K638HQf1PaTHtbDKN93fgj9cfztQBO13nrsxQtN
v/ulcDgM7QNBuR2sPGxs8hIh9q9v3NYqZ2HTk5iSKTXDjsfUNbymM/7NBuSY0VN2IWCvhb2CD7W6
+FXNM9qeHT7ecaSdbGzubj9ShGcIIFoCHQcCIgwuKafkOBENp1wpMuPGustdZgRCu8Ha7NfnoRfz
gebLouNtZH5dUMT8+e9kdKUombqni8R8bl9wQMa3SIw9XqKthwVvGUamJM9Icrtq+LnDxWKlwcHC
J4P+rAHCGAI94r3UWMRGB3ZyGHNFDO5YJC5RVc99zcXAHFSUxPPNpCbycx5MF19U4UsHAQmkUV1L
unJ5MR/FeMorSshV1UdnvN8w0/3upLQTtAQ/h+l1gDJ6DE82Xi+C1XKE/iIkClNyrgDoip8vKYDq
Y8AxC/QM8J0A/7xr7V3GVMt/DGgfipb5+ivyvLNLpxWiKPNr8PQwdG1ivtsJNB0xjEdD8CcInnny
OODXNqv1dlJwfA4XuiPdkD1ivFZFkDd5GEJyJdUIOaGcY0WweoUZMtcT39ilmcXS/86jmSKayhO/
JYBNVBwrPcjl1rg9+5vNIZPbJNpnuNSEiUHFh8sd7ie9DpHQTva/GxIvFHUcQRKrXdKBCO3u8+jx
oO95KnmH8qVy1D/tSEddonUvwmeaXiJObbOtr7fXwF0RECPpK8juXxQQRrEFPuoMxsqQtxB87lgp
k3F9nbAvekZvvnggOkvJLsFXW+ZXWxSV7SoTCVDPfcYQTTSmSJ63mCSF3DjFk/95WfJY7ZRYDR3E
ORn7QzFp9KivKmC4P0yqR887eY8iA2c5d49zcJaqbL7ae2Jk3+oRey50sOilj1Ho/1+vZfNvSaE9
nqX+lO1H2F4nBb5qh5W1ErrspfKzTPLX+T4KxNMFumKewTc9qhXhcDJfgIMIRCrG5tETUXKpISoH
m8kEY10AU4wmV5z8vqvbJQ3clfDeyt/k1yJZZLXknN9whwOGzFYGOH9CTuCxDiPyLjEexMkMLSdT
EgKXW7vK3kqTAjHh8ntIq8me0I+zRWxba0eX8PJV/SawoZPibkLwllpXZ8SuyC4irTfbcyZxFvUw
J+BxtWRC0noWdlVTVIXyzXoLRKFSQIfI6aeYnHjeVGwESWUE8pFlz+JFhEGVIuxPXbVHPu2box/m
J09pYmaX06+5gwEDOyrB8Q80sewW+OeRtgJTZjX1eVmgv6dSb5130G69OE7Y9A37OpFiciGFtBud
XXGnvmZZC4kZQ9h7d4CFtYrtfrPDX4OJPe1o4l3krFWLIGNro9zv7WHIxFBD/aH1DoQdySGv6Lj1
46DpNCVnoKob6gHY4GsJiiRfHHOrxDYYkBCtrdma/szTnYIeP08K9G93rOV/uKJR2erq5KHSTWz3
AEu2q0UVzjvZEmm6oIqv4fzNw6Nb8AvBPTJDft+8ZXEWgKVxOK+ggciVktv9oHjw0woHU5n0r86P
pUmoYHxxUbIkDS3anwnJiPQynlLDc2cRFaZ9JPcw5eTY/sHI6xzHFsbk69qK/dSie36JJ1E5XmnR
Jclsmf3mSnAW2XOkMkHRohjg6WCysQOp7BfBflBtpCo/R1+RmysF6IidZc4+Q2CdUnX7EAAWyU9r
rElQsMW08QDG5V7KNiV4cOtd3IvmSXazDx5TfVQSCo/eL8D0z8RF9wr6BuWadACvajVvfrzN+gZ6
WPgSCnw71Nhda0g5dgdQDd1QyB212ZXuYvMO699QPHPF/qOw7+WdqqoKY57jLNcXnmXhiD8g0KK5
/jy4TzlJk+mI8scHJfP5Z8ApWqPFpr/RDSJck1DOau19jCzibDKT70Y9d+mjuhdxYEo21es++fgo
D50qt0FJrtOUWm/RzGMZL+lhLgUgm97FYIdiOe/SZA4MCRqLq3fbHVTU4YbkbY58sMLxsFewqLfK
nRLMXrRpjNjxS8/Hm+usFCowpXLLaXP09u8eGEZiY87V7uIVQIITTEvysRADSIz0Kh+74mXXMKVI
gfvrKRB2v3F75RNvoRPulisUnQnwZVqeBjoZrjZfg8m0o8JobIf3vNRfWp/1ZBBof89nYGdHk4HT
UlNDKagRF9MMiTI8rp7EN7tcsSNEXGi6oXMo/wU/xrn57+Ys7+WWCw6Y2nSvub+Dr3P1aICFP5LO
qiml35kyjni7cVNMIZJ8knLW4zwwh+ee6TG43TZ+uVa1xeKLOuJjmHridktL7lqgIkMUbkDctgNu
Xt4y28xy8O7Y4O38RDUACf2XqnzaIR8XFx2akb8duFf2kNlEC3p2aMb+Ye/wTp4trYMXianNenBn
w18Qoju1s+wEb4/DILJswGq/Pc1HnIoz5roMP5quZwUcqMqVp0E7NuBp0mCyM/qqsPDsRKsfGZ67
g3NxgkwZNyYlDC2DqmW1IFDYNbzH8Zn3m6V7BmmD0q8G5Sm4+OZWBRax1r20ZCbgZbcEPEbV8jg+
c3NbXb2d6Ma/9L+LW56O5Qzj2YoV8Uf7B9KloDauUU1yKjX4j19Q4BfqGLTHafnLK79iLJfLxWaG
9lDm6t8BpAT5xMS3ST/7w4KOwxN4gZYcUySo3k14Kr5NMwbWb1aDhsXf+zeJvkfwTL//7/zhngwK
4ETi8uY0I8P+RAuLlzLDS5d5iF+q452lX5Zp0hoV/DZnipZHGKaGca/FpXGkDpxgasHn6gp+wY/K
qEMiG519EM1KIma/Z6cih2axHzjmJbkfpF4kJ1W+2g8et0U0gajnASTHCj15Om+JC50wpe5+7ZF3
HecA8ABJ1SM27FFf5DlrBmuAl6dZmABy1hIEmKNKgCQD44g3DYwJbwv9jhb+2MuuDY8tw2QypwPs
c3U/7MM5kYS3ad4rRI2+qtTe13+/sbuBXY8BOJ32bH4kEHtyvcUtNv5Rje0vo7q8DSeNT1scpegD
mONvQXGNGzh6xcLfiU3PKm2w0dlPif55mgQjRyP+G1j+fnBzwsYlShs6kLyRrppTa2NJVf6mT9xZ
DdNtnT7SfwWFm5ccaIV4oA5Ma9ENrvB160Y7agTEi5upxj6y4RwsDpSEvKrkjYJH84JoqIQQcr/h
Qh2W+Jy5gkSDEyOSOfk8d2z8yhUwxruMqYBoQjUfLY5CDpu19nyzkfZDy9iVHb87qSD0RMjiv2/j
GAeJwdlStctjrkEwHr5faX8dQccvJN1TSWQS6XUDuCARsP3SQuDen+H7ugWs/6IbEbWmLjVMRWuY
Sg0JcbcAPEV+T4dorrNAKbyg5E2lzCWDLWEfHUcHTxL0mrKV8ARg/2p7yD9sVfUrpTrxQo1x5L+B
ZoA05n6sjfTwBgtibpcfjsX2Fkd7TLFn9sX3DW3ql0APm3YwxqhZ3v92HLl5WFTqyunJbVmsGK0Z
53ZHjxfoFGX9Czq74eHAhuzlfK36QmAtI/fJA6wglazvjNrcwxkx6zi7sWoESr6hKOYF7z8Fvr+r
WpAVwTa5x3N+a4sbMbfNEJ+Uu83GUoPh2JUWCCrdK2Aul0gzloPyFjI/BUkDWYGZboKW+vY3jBvQ
lgaaJyRB1Ehxro18qH9naPbkBbpeWdiSvp9Vr/Q4AGQMV6jteXghp2ts2GILF4UvM9a/Xymjsg2Y
cyNNI7wvT1Y+cKxBFSIYXgX99jb//0AmHAo/ZZFnDiVbyWWbreAMqCnGAUArxlJ97pMmMpf/YWP4
aVPauvPZTA3W4FP4MGqXEtNf6AK7CONdgkQA/4Rc7Q7rl+qDdUPLPclAeOcv5pxxHYaktowguJ5h
JBik/pJBs3fCkXqNbEs7BPcOdeIeThYZT93HozRxPx69g+v+k5epS2ppS3+UcTrzYcSHo26iN+dF
Y6RH8Cx/GPL3ym4efm9yTPk+xnRcGk/RbWVFmz1qBbi4ngb2MrXTJhPZ3TnB3IO8NlQEIfVUXtj7
tAHaxQEgqdU52ulpY7xyI11DWUxpP5Bc0cc2Jzq0qRrJQuAEw19nRNrP/7+sbk2CbXOpcyhSQSQj
RGbzzje3RcdaTq08Tzkj49sRw4fbxSOJ2euEkb9uAoL4MjfNzN2i6/gEnQtGQ6jUHkG7enUJdui0
hGSmguOy8Np92d1KyxdB8IFMK0th53lKV6nQkmKQRpt7DHwVw2SH2twivFozJ5L9YSqr3LG7ZRP8
H9oNTxe4tu1NBW6BXIQ9vyuNl4Tt9L7+D4SWDNSzp1JiyTchsXoSEy892whtyjvUWBj/e41G4v6+
F2EMIlWzlg/cA/BGkA5Ug0PY4wdAsP9nMg7RJzd32mI/2hJZP4CdV44QmPXvHmyd5idnW/0vuzqA
AHrFdcjht6buUSBEAVvAl+2oTPaq4wuH9rHHOysKUbUsMgFHI/Uo6zkmvDy0rjXskFBQyBub8iGv
EHE1kmvJpArh5JGSS950W/u1LrF4TIP9bVeAVQTf9wPftH3KruTVXDoPPZTRJaF/0KVrylZh7ukA
Eqekqx+2I/5B+6A/QZ4awMjynq/9j4coqpX/V2TNzo12yynWLBMY7Z/JKQ16JxZPF6uAM9bXBOvn
+cdTKzJyTrorI4n5cuN2qDpNbyQ4+X0CAtk/tm1Pfha51ESUZXrG7tNubSGRvXI3d8zqj05Ou6ZD
NTF/LNBLUVl9s6wEg/AjW0ewNn6UBkHw53e7cjfE4WnRQaQgbI3ylqqpFjfEJbSijZxkZHSBMvhn
AO8CpfxM5yHCE56050VA9BBx89IfPWb9W3hxNgUX9MLCOWdtb08ei6JjCHsn2Hvy/QIsOLuBWo35
Xyk9JIzn3sL8F9GQUbRkQ5eXtksdFnrFGb8Jf+KlMC8C02oqOGZOAxi6iLWe2IIna5LKo/MHeKE8
bcfeJj67C+b5Fq7h9wcsoXG6z2BsYdaXBnPytqTrQb1Kog0EjI7FPlBWaVhmN2NosdD7unKHc7eZ
TyovBZrWPjzfUZGypQi49wQ/+/TU+ThcZ8jo+Do/I5JsToiWeAKKfbaq961NOjChKILIzDcjkhOt
/cgtMCZKe9iuRfs2WuWJKIOJ49Pu1P2DJrY5mE1OkolIG9tyPgHHiKTAxeMY0wS1Y1ZeiRz8N+E5
vdeHJy2I+GuAZ6nu4wjyqBE=
`protect end_protected
