-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SRnwPxour2JG6gJwrsbXiN75AZk+hW5nMVB6Z10aNp5OOezwkHx7pfPjuM8uVkLP01HRUQYz6xT6
R7z5bLs6TmGqC0sl8Q7E0QHf8Em2s7G6OkDP8m/oWHy5hl8YuR0sCPJDxmDx/e/0vyr23ZaIWy9R
lfvufzjmiy8gOblcfW2TdR4EMjr8cDm+BJpiJjRPlmhxuILruciYe7+6BLpFa53d/gBMJZfOaSgP
ozt6JvWvu+k+gL8dy9IRKj9AeL6YTfnkCuORV4kcqL2qwCEAcsy9ln6xPmWkLtZQed9z0qTvc+8o
PVDLNB8YsazvotSTfApX++3Ncq2qDyM57zu1Xw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30000)
`protect data_block
BJUXSTZ9rbjaGmq0QywHNP7O557uO1NalHmMX+Tz+zVlzqzvinfGkFgTMxbBPkhbEIEGMvOLNQk6
WGliExFQvccqAuKaxdGlqg0h+1ZhbpT0WPwrqLZ4vOM+WnOVNC5u1tmd5mfoLMdZSLlGaStkB/Q+
QpKHSZGlAtAm4YlK9b1Fgu51UCOxSRTMz3gJaRgGOp74FTEexIB/5oyzWj/gheCaAKz2dyHg0c09
bWxf/MYmqGohVciHzyEVEtcHkAa0dAGiDfcHMDQJYjwWNs/10uQaerRV56TDNDz0rqzdIgfmJFnz
H5ruP8BSNrXr36jsyakQJpuy7++Z8eyr6Vjf5zIj/CMiVRacAFP7NVZHUC2AK9hC6CjuK78TFTFu
SPkwfloAhw9EdrZgYsFnRIa06vqmKpPf+hfh2J/HbpbpyKvYVzsqsJ0q3bV65zV3Hbm1muj+5/Em
WeBlzQuBZi5mwLKweiKeWlClQpLwhpYYIT+qwXG7DQfrdHe1cBEYmWLsZoH4ARZtwmpfqlm+cOh9
ImhbhQHVzXSdm2OCyv2yxVto9oNErY8rY8kJg59v5VAXL8xtbuDok+n5DqODtJ2VxHEbkrqwe0CW
+pqR2tr9RC+Te7ZcfBL6J0qZMwUv2wHeDtLEOrSUCAhvJzol961eCIkjbgxoB1JKeYz7G06p7fW2
ZtC9EJO7c4zv+DOxOVNGa0JYcXF7fmKw4Suojq5h2BqrnIrpLy+tTLzqUtr5MNmfeePKul/Hvwlj
nuKz0tj1J9cDhMv/V+dOfubDmW+XXljyZomwyZ3p4O03qcL+NVSbzI+WRi/WWWBNI93syjmUE0/g
QjJCTDEzCSEuKTqf6+gRbW/eYDpyEtQhLGFsJkUDSUcqrOL9v5zNATlHY/iiEFIIzPn4KP3uA7+x
I3IJiDfn7phuLn2nWAGA7IF0qxrJrojNWbn5mnBKEDyUXaX4Gkx8PbOU7f6kjWY8wIWkrRsGVqY+
8FqV8SAFFdw1GXAM0uCpyVGluIOrJTO9U5m2jp3JaVvKxcAZE/qYKiw3YRuZdd72UiGnJc0NEkpG
GFZML7m35SkB4CLDi4ZHULUggWpIJVJoCGX14D9dnhsYnKbwarFNvdOtY64LOSspN5nec0KV+pJl
hGwUlPMqzwVma3OihX8ZorpaWrIVvZBKqbuOHnXBrQr+pGn7kCQqxUBl1ZFKLdCXbi9gRRRnSkD0
VNQPLIJriInzod+EmBxXJZd0PAw8LWyMv6MaS5lcb+a5K3D8hoiFxMXlkMmqiMjG38JiHS8FEaKO
Ouim6kh//I6JZO1ldvnVpcjvFnJttlv8CCiWgDMuEaqsENGCc6apdsTeU66eqUXWoyhN6yMMbm8D
WOVyLrwpOjeWjTaEAE7p5cMT7n4Z2/vXdBOdtd7cGK0h9eNVISSTy/du9uXq+F8PsLROcty9Kg4D
46/eqq9TxcCjR4o9lH0xo+tvUvjZwdBDZcLZ1/QO2Csc2gS1HMa6jW03MefMZktjEyyXMq/R3jXd
AnbQ46qX2RrFAk1CgHh7qflVuT2yb6Y24/fis8jNP64AzGnmWd8RLvVq28sNQPTxACowN0qMiu8z
uJOKYRiNoK5LWUqQRPvNJC13Q0R3OmWfUC/JmMZS+2dGdS6PKhOthG/wxkrG9Ix/wlm0U5+wvvhf
05cFx2AOsWxag0j6IEOQY6criptrTqjBD0ViHDgMGg7Wsr29oqt9L6NHJ47MrVerK2XQYPHet7TM
yc6cV0AVvyrVxxfoL0xx1hAHm1h7/abFJkN7xgwXjD2Ijwk2DakDhTlpeBiIV7ZP7Qv/peFDY5kJ
WEjDLafJQYvSoEQjLhcnWsjW3grXa/uC0Mjh+i0BN9z558jn+b9Q9/DAkPUnOvkueuenDZ1TNnLt
r1POto7VMklMXaUfd4zir+J0asW+1nsW40eKaAFUjhkGCex5wzCQsG8v1ABDGMjhvup5f1pSY2PW
TmpfddesTNdS/Cb+q7BGAWSUp3chpYymMAgLQELIeiR44z5+2VaAJAzslQ4MR442O2CINTO4dR7s
4LJ1wLU+oRu1AWC96JsjqY2Ftkp8BkXRbITmsQYG41MAcLD0kuxH4PVAjphTLrV9643360NBQ+sP
BVCc9ZxUns9ARFH8tIcOVAWriBph8X0uvGIowPqgaCbyRpkQ7Awv4Dr50fNFR5KjZmjr7qD3cvEK
9+aoGDg7Y0GI6169FtJ8P/FIkjQYWmc8DTd1tl7Gu4jcnSYU0t9A+3RA7cgNpU6VI1PfdmAVJM/d
2hTadWurR2D1qIHzQ6NbgcpxqeyfRFFbqAVxw+61kOZYmp4RV66C9WvzP4KdK5OdZj87oMHAW1YO
JA1Cr3jwwIITJFaZ6mNDBxpCFXe8xx8Uy0sOtpGJu6UoZ4TzQp1Xt4499UIyJZJxy4DCxHv6QsL4
LrI270K2wjlvu3j37RSwzeM7+CFqFEDBU7D+wIFVYTpbIPBocWd8OzfXMDRUYufGn9jPYJpnI9ba
N7ZXBgG/xfjODk7dl0IPaHIs2W7eI4xWryTnu3uWTbLYEZFTrHV0WsadbeWHnqgKqojUgucDORa8
2v7d9ATIqZtFjH2OCynM743zpIDjBEMmVui/g6ytussGTUCsQl3v4SocY5ua1/7koabRb5NHnX7d
jBesi/4s56joK481pGqOxGbVZMZqd1YE0mr8rHPNzyiRUYz0i8ranmQ27s8j3bEhVfjf+K1ig0rO
8UGiMo+l/U0eWAvLD/uov+dCc0h7VRgFIhWMJI3mPVC1IgaBIfR2dFjZJ7Z2QtiEQFPs+dvca3av
gvGyVI1TMgniHbL1v7UDoIvwQgvrLvxaAG4Tj+x6MS/pEeHQ0tLQdy0KjjhFheXNohMsyJWsGMDS
SJ5LkGLgisMUuoemoG67GK8aEOnY3+0Z7HtCVR62zY69ZxiCPEf6nuJSDgFpAp3YsFFUngzISq2O
DI/kttF3lDszt5jpPvZRieLX5nyjlCaSkFCd/6C8F26ftIpD6N3I9+IhAjGcojnZfWdYc5HUeMo3
nJnY6cC0qX9a/Cdy3KGTwkx9E15A0beWsUT23cRnSWRzN9+luvMiP7jHvO2AL+PvM4d9zGWSYFhD
IM/6pjvekTSf5mvktwUmO/le4sJvfIe+OllWY/2hszrJ0rOmHlRBmh7wpA7yQju8nMGMAXhcY4oR
CI81qhlACBQjoqPZ97+c6LxvMduRPmwOxISdRx3iX6F4e7onFnrXtWGaiiOLXD5zfPNoGeEbAfr/
7OFU3+Nx+GsOWYPc+thl8Eqwsheksvk2UXL8rbUAQrsvPLHPeJXDNkOhm6f+Tu77GPRmhUXUkUQ8
35dt6anxC/Qu6iU+HPrZypszSom2l2E9bxvVNpFoU4TvsyYZVhBBSliCgaEzSLTca94Yc2xw7wER
c7SR8eFL2bsuYTwy7WagOfn++D0wmx+3vdOKzWhRLoltV8T+pzouVnmCMV14f3PuElv9HL7tQ+fF
PDRGyvu2Zk1y+mSn8AS57YCK0X9m8rgKGhrAHluzvFBaTd31sP6w0PDTF9LG9SyveTpPOF27IcVV
uM/B7vnDZrvCGh4kmMNSvvfkEfNN9soU6y9Ob6K9fIBqO0dqDoVDJCZfrEyo7OeJKQrMGC54wcSd
m9Vg61Cnf1kPq0PK5Oz5pjzH/LI0UOq0wEoCy74uXAqWpiu/y0WgpyvJRKnF3scs2auWP+PyXDCf
OrlzLor2T3m4gwQE1gRFcQ16M/AUgzbA9kAQ5Bkyl4QVNXoOyprVE/rxQbvSEEJ2WX4H0KbnRJqP
jL/WuN16wXGpGUqZYHWR1jOi+DYSbSO1OkQVJTGv3eq7xrePXDPozVts+IMRWmFuOc1TCRo9de9x
cpHqNFxvoRbDv1HPoy+y6pU7B0gAVss0cr8aPHm6UhtQEIlhTgh06mGgt5JYaW+e5Q9QACr674Q1
F60hBZ1WLTO2/JacwkYymRl3u+s3+8JZMOFETr3yEKwT/ATd2u+YuyDB+GKi/ax6Lryt771aqYtz
sDd+b+8Rk2kczV/JLkwE6vT9dDr8HVB/PDkbGZ6rGpbmlYEHhfO3etwqx/yzchnbv3gZYDqogPt3
jPzo7CMc7l3qF1KrlSF6Oc/aQ4TaQKQSIemx6ZpK8f+VbYL/NEHOBX2ZYyQsFRB/cWhFpYJPOnuj
diLLiWe9ptyXEhP/9XcghuwtD5vqwkh9dDzh7z7bd8bgQawm8aFYLg69+nvrEcWjx+7SyvCOHFkB
TIWGFszPndRy1t2ZSdvmapi1dV0RkxNZ903YtwY3PHc7bSzDzx6A6KfN57QvzwyqjafBCx2OLh14
wt9L6YTkrsWEOl4YfmBKzaE3IqrQK30/GS3ru7zI+Wfmx4jas+6hJsQgYEOI10omLDcp0FM2/2tw
tCMwxECvYMwXype1cBp5QdCFmJbyGab9jEnfqG5D0KtvzsBIHjvPvZUlJl6HqpMqTI+j63c7lt6C
eoS5AG2t5XFlkJhJmYde0f407aY60uspoymXwS8zyCneHOFUedSOtlJv8ka8jtvBbqLmC1CsPSmJ
4BB1gr7UBS6akHx6IhEwYItNEQMbKXBZzKpwhWLfbV/HFyKyS7dnVctuDjPdvWHoqL0gsNbHpb1i
yfUNKcYar9k9CMQSQueO+QHUoFNqvlHRqbMts09RiUjWiG13UzsgQVcexlqqF3w+M7a1Vaqi/pc+
pvBTE10RCFVcLEYBZD7d7nW3RSqOpgGUAJWvmMywZ8UpuYpGCfsrB9dLEFO2Au99C4Ug6oE+2NtU
1MG45oOVg3cxnRrmLEM6y8uoM+Ip0yJdLToSGpU7wt7bf0MF85x+vtarPSq1Hl2c1+bSNvtVkXfc
6aeXxJHpsl+fnZXNzhh6Xfx01cPGd8RRye5tilf1XyaGTU603zQoyczzUEX5FzZOhsxKpfyI0wqp
i5SBkczK5ipaGljOmf6uYjnsk8Kee/cEMYO6HYstGfmRETVNdzzpZ03ndinnnqrRweMpByRenU9c
crEtiziT/bF9n/LMOWsL/rTlhRFBGrab3UVXpZ2RfeVd4ahXKuqRRPkxXHpuG71PY0Oq+CZfO08V
sBNxa3/uQgNPXc5zAR2TJ+Fxn9DrYoRnvDur+CDxWnZKNlL5hjvl1Udrd1C39cS9lbKoqXm6jBxn
buJTXXwjT22FkmrwnkUb01xRwnthfuQW/jhSZudODOE6KShTpkCQkD/slZEiDFfjJPyYxutJD5pL
vblP4u9kLO52JMRZW0iy5MxARsffGAJPg0UzjJy+zOFFXETx8sMAs9icn5cylZZF1AX/VzKHOMCJ
tMa91APoEJmKkGZl/TobJ3eFxaVytohQtnki/upf2OP57IGd5B+WNtavvh211bhlZpRuijWVBiEc
727s8J0+9z2Lk84Onz2+QR111y0VzSaHDzIiXWrCl6/fvyzu4GcEyGHbuwkaJW5rfYJJx8Z7VVeu
my3aBeI0z+LXm8FKu+PnlE+5xEp3QnhLn+w6gVQqYJ0oSiG8uROhaXuNycCL/swshZfO6zbK/9M4
Z6xZa5/2hOqEDUnJoJZHGhzXpNOkKmbd2Te7MemSoHMF55ZZS6lZVNxPx3kOxEklwR+2KvKmWmzv
DHKPSSj7T+CqkeHr2iztweTdaMA4z5DfJRXl4/8mloe1WvU+6Wi8KpHNWVr1gR0B1ZQp8MAz0n4k
MdvZhcXA/3frwCBI6b/vif5SrTOEptcAqvzdr0rP0AAgudpjl6VnI+80nlbs1eT7Rn8nRTMDwZ2C
Vz4RnieIyIaJPKg/YBhCm6lrEEFVjj4b6hjsZFuCddAVcnEEydFmq1VyVHEV1Ms20I4jU5hWiyGA
1+0reXaTOfLiFwIC3RFcFv/O7Hl0CGEPl2+SCAJm7uTXeRjLXfdm6ULfFhcSxSl4iDNrEDOb8SM9
vNOSAFcFsSV5ohhdfqmOIMl9Fc884oCMtTjPvwxUbuCM+I+En60GYZJxx2unoSXPTVYRmInptKBu
WvLZG7owfAcGslKPR6xPnbYlkGFJ5Tw0aKwrPGVgQ5+jntjVr3tv84Bo/WD5dpCBuRMJOOQRr6TC
0FXNqnjV+4YxX8/VqMS+H3L5+bgNKuUBOmQ2M5imKPxVpkikt83iNVmanGROa3psagP1bLBZtlJN
OIpS2sd+btAGJGCTD69qwdNE2jusSHm+PRgHJah9noZdeoRNW/H3QPkhi3m+fwS1kE9Ys6n2J1Sa
RlrolZJFs1qUf9PUj1oS/COxb+ZSd2BLYgoe/y/pMoJBXNJL2BphDIjKLlY7a/dBhcspYH55+UKV
1S0/PDToDyUpySklmxhelziFJoiwJUM8L+8YRiS6EP+f4IkFy2Hezy6SjrdxnuWzZXBgnlIaLm6o
1qJsbdxln89zyKJhnlD1ql+USr5OrP6ziJhizWgmpuslPVMVpqgbqyRSsfuVCEODaaac44D8DyDp
rNS0/+jdnigOZLCHhKK02R6arvPiSIxEOf3tImPuLeHIKtKjQmBR5aPzxKS0wwnscCwCp6JOfCG9
nU13TyVPscVrInHmqOMXgVr0VpGKLtjzIBafrhE/yuPuDR8tH37gXFe2NhK3qcKm20aRrYbmem/L
gWAFDM2kbns+2aIB+yBFhsEX1CY6VL0nvJlrp+Lb5IQFzFNBJJM9Ejuv9ZRyoyhn3Zo0OUFbtMGW
hwhHFOhG8u5/AOGziqoDF2KF+vp9H1b6xwA5Gq9U+NDG21g3kGygYedd8jxRBastzR227rXZ8kVe
z6+T+K2LBRY4+bVbE0+t6f+njwGE34+E4BliunlRa0QYa0S+m0ykp1+u3Q9y3f+m4JEKUOAIj8tt
a9Pad6DyuFFH2iKJQq9dIZuiqWLnE+pOKXObfw0HHrwfRyeYDyVCQYdkwW2ojsh6dt/GWttE48a1
HclymM2TZ2LPav8ZlCdJAEyNLJmQ8FKwZJaPhNyA3YeCxjelG2Y4+ks8Eg9UId2rAUfIKuIHgzm3
nhWyrIDoOl43HPGvFdMINWAFmO+ITYYnM/6K9HEshylGPIJ0qW9wn7sr8r2ELsuvbfmZVA0RvxBM
pOAzwEfFnnUiOvRW1ci2c+2CwQDFXKjkK7BFpbWEST0IzBtqAD6Kcz5WwS/S2qf7I6WcgC4ke6dq
pUWx6YqhW2FDe0vwJBxuZ3rKlFUevyOPEBvCC95Gyh67yIG2hAua3NTvmC6c9SP/doFYUN9DxWDH
6WsGJGDqq+9ad7BPy5nS1Jji/mS+gWbD0TkI59V7gINwUY2S+Lqs6UAmC4sW74zPmCauaaZzmJRY
5kSvA43ydf8B2EnPyudsiGwwbXRvgadI4pehAY5u9MgrRgyO5n0f25M/0rTjjc+VdCfw/0O5+UuL
SLRrHgUMv1mols29l2DS+L+9wiWJeyUf2EsopPvT/hhFIT758EQhMRnn1ndMRpcxs+paV20+kvB5
MWTVrnGreabTfe3+U+j8ikkLdZKOTdNOFJVUGeymMxumVS3cE69ylbOqCnFmj6GSoox9qMMojLTT
jnK1pTSJ6pZYVdSW/zgjFwwMFL1DeBYubjnDKqqDjP9cZAjTZ0OEkTsAUQICgTCNjnXCfQSeleqf
uNHpVs2dEeuD622ml2I8JNhwBBy9uTMKUNjCxZ8WEJ6sDR4U+y+Zfb0GlKbNb4pdhzA66uyfxLB6
nL/sPG30jy/BxxC2mDqJg/XnJWx/idaj70YOX/N+F2m42fi5LoivyDgIigQde1/UuBRDfDxMTwq5
v6oynCui4ihpWX2KQrBtqFhNcXADkNcc+gmudc3B/HLmXdgA+hHuES11/d2v3E5ZsGJkO5jzPiR8
t8qXjW1p8CyD2OOV+hpKYMN9qwqk8w5X9jxeWEygggU5P+3prw4iLwvea80PcHyERV/fmtk4l8iB
dTuytoKUMWKXVUNzKzGZdU0mWoglFU2hc3y6pmMcJ+tAEhVtJO2FVjjIwBVg3cNVsoJYT1wKljL3
WxKFFuE0FlR1jAmuUhB9kEoTQvpqNxH4mmH4lbHhm0B4Mf38Uqw3AjS4GLBZYNMHNgn7D7qQ81F0
BijFqcY0ksd4uRbYZhQEpskjfMnlYBkvNbMmdBBAt/60BZMizek3Wu4XyPCObhwPoB0ggsBkNGyE
tlC/twmVUb9GIOYWXtg+tr3eRoYKFaEyt8ZXiBH0n8ljHufugtq3QFc0fWgRImzsSydOv9KJZXHn
D65BPzapHc79tBLBb6Vh/cnSAyOnqbO4Wyfgly1mMU5LPzt6sNJ1sRnuFK1M11OSBu59ennO6aij
f0FyDdfrIP7jHsf1yUYN3RdsSd/7NXDiyuFpKivb+671Pz40l+ABo6kYnBSDcb+zcxDclTTYmzB/
/jwC2KGm4eCw2ALA4zPqhhSU7xIc1LZg5qRo1lbbuFmokLUKUb9bfi3A2tch8HpGgOvPqH3u71K0
xlTGKwao6bISd8ThsRble6cU7jfsIIbhUXnUxEj+e9BDaobTm67Hnw+JHIH//UHXjdejrQLI5k/e
3HTnyhhm0mYCBvWsf/kdC7U97inLmXVYnxd4dfUhm7jLTuGhSmnYDJIvhZNbeM+FCF6kjy2pi/Lj
IeZ0Tu68xLyGl68kr8etHqqp9cTLHI/oJCVfjkVNKDdV5DSJb0UHLJ7dDz5+p5oE94UPT/0WLWT5
4VrTV1wEimkC+PwuUTLG0ZPVtyek5d+I+9cq8KIKjZiF8EyTuA/GHBtiRWKp11+rHgV9AQv3hAh9
inqhyuuevvT0RGKuQCJZFsty3bWN7ofyQs26HtdxaePQUI2Wgnyd+5TIFXZwCtAV3pqs2mkohuu/
JMA4sjGdH7w51AuFDx8HgcNE4CuR4XyeSTMqGOHJAqVE9mwv20wJLuPYDbtJpw0kCtcFkcgoxguc
5C0pP28+iuiOKyAAh2qD9pB91xs3Ov9BumpDwUP4T/oyJOTxu2X6di3BOULyfEgzv/FHVK1Kblaj
/OMoepKC1EjKC0XJX37APo71rKi1BzsFAxSW+jC8ZHarYOZcsSYT/OhwURfOI4+tjAorjnJwu/yd
0+6DOropZVoHezJyNjDKPF8oVgQCYiEYC7zBFqIwm5TClepoY0htuHcJBYCyKZSWLQRjhFAX7c2B
MSSwUkF7Pk3e+xza02R8s7c/ZIRAJdmxyA9wcsE2XLiN0L2C5Fw05nB2I9f7y+Rg/tk5cgE7Wf8d
AI/LtkmbAv8wr8q3CaT7NJUNX5DXOYQMJMLQGdrw1JoLvvBmbFCBTvBAB0mZ6TwQJRcbUpHsuKEp
xLCvZ+nIjPjPVzIHcVY/ErJL0BXJZCG3mxnbZ3Quu6ouB5iBSIM+w62lt2hkp0F6HWpDGhdiiDcc
EsS/Yeyi/Wi0pzsTev/tYnK4JwDHh9Eb7e69t/iHB7AgvPoS0i950TaW97mYNNBavByxaS3FcKCv
K05YjdmILmOfjWwF934dOn4si9mLvqWyTVo6PrwKjF2lj2gwpfUMzI/JNxd/amP1Ll76RXegaVn4
YyrzMIGyG+A6HVki5V3BX8Zr+ErMXoaTXTiEKfuUDgndlmwBr3qtDMSxpekPN4gorQ9Kz8Qh91pr
6kthRtNxZeDWb/fdMWBlM/suNHEh+qzPoFDvCnTlT6H8UdshnQiETn6mj6qGhbYartxX+1YyU1AU
uBHzQNFnVOJq8jouGJiMsHMw2KeLypuEOs+WbydIm9grfR6+6GsxtADsp0kFx7aCNameEhKKQVUO
pvANvVWFwKbnqXZQz3TssV4dRSklL9Yy1kGPu0Zk9iEWTWbxuDwnus8SJstNbSbZ9mWbIbz08yek
4GBTJGNcu4WFWDytwdboTrc9qzImtOrNC7Rr0tMpPUJwmOG8gF8vf6j66j4Uddrp35jDbu7KY2ht
gVQFa9Y/JwNAOBp9KDiTLLr5v72hrjT5emgzw1f/gweNoi5c3JFIE6/mK0XJvH3qsFKy6SZoydug
LYg85hyAJ8cipmRwYr7EiAlX1AiCzDqK260Llt/SPE7R2+1etfLA0B2rNZv1rrZd82nzrlB7qj1d
0jSdurOYUQS+a5sVh9sxD8EybQ0v050uBV7xlFdBQZMOCOueNOVMG7aTbBID/fGT+ohBMS+cGNxP
QtIhRVi6Kk3sKzTuvjpusmWRYa4sKqLPgu55AiifALSMRGr8YOnm1wRSpDbuvU71Yd0YykOyC+mE
CDQVYTEkxgZpBvzooxfuC1hcIMFiWkq7UjfVVlhMAA+fBf2CBWVJIK1ynortIgFowrfbg+IwTFHg
5o3Ww6nA+11cVBZ6i6tZLgoqp25SO92ztLaWCzW8dSAMgZYB6T+9L+yzifSIxtI9jG/rz5n+fS6X
XWFyofOmOe+odjQ9FHdRy8d4A4y+Cvq7D7ObuuxKwZf9isvOj6dFTJiUhq5gBazx7zJap0VXi1/l
laG9X3rw0bXqJpmFt1r7fwAqBSJt/MbUuVz3vP44L6fpQ6zJEJyOYBle1N60CCTQ0/oS0QrVS7FA
0EayC/bg65Rb0CMstGknQsNA08ELlgQ03dkcK3fmLolJkCOEslSuZnoqS8thsSGnlkEQghSb1qqn
8z6E/Nbc2Ov4XYbDcGof+Wtjnmdh7egkhBHSMH6KivrUoVzEZToUZ2YReqg/zrgEBQE8pFompeXW
zeJj5GWMdxf5awe8GmYUONLjn9+XHT5YiusXgQyT2DtYUqEnG/qYYwKOnv2UNamkV8XoajpBj4cd
SRPpau0AgfLd9p28hCv9KHC58vnoyzQpaBgFJ8nbZx5V+axPsN5K6bECGluVw1mcfK1gEuQ437KU
B14oGDlQO8NsfStkjk1JZ9eFHW3wdfEfjBRuubUUwajqBCE2O21fmibdMjRcD0X/a+u++1aF2PKO
j8jXIC0pJfpsuH0PV3mf3SThaab2bzThOsvTKCJWetnYLMwF25DXNnJ3YGCuF5HY4N4bOsXsQgsG
jR7l7Nu4OuIeqw5WEX8gV0CrEObCvYDZju0Gmv67O8XMuxXNAp+PCbFYgpJIx5nQXbBZA/oHS0lI
pX2t3SWB96BnEEVVc56tw6VErnIOv7G0SXYCVWAchZvq5yFksC0mRjyBmWYWgIhzerqwkWLIN1eM
nn91st6IAtwnye755Nd4tETEfQ/EdB7qBbg7xU7I8/wsOJsVthzsVB2LCFWcWmJ7jGtKshe5lgie
9T7QKNvomBLVff/0ez4B4xjPZZjwcMDn/w1ZkbFfJ3gEWYSryJUSGT9C5mFd0x8ALsLZF+EkKms0
V87UkKfzTjNXmz9+3YZcQAxYZsAuAkYt9zytfIPEgonpGjlpBi/q5cxMMOI9gl+XPODPI3zxuxdN
diW8SAeV9mz+QvSmWAe0GhTg6qVuRgwk3UbqpV+tnbpsXI6tWAdmCQjOQIhzD/cX7P6CtHvsWags
MUV0+qw3TFSIx2pf2loPZj3ObjIeoxC1FsQXCwmE7fvNd3RH1IEfXkuBpdly6+14imNNjL16zyOO
2saqsk98Q7I+Me/pzbhVusKdsFZZijWJqiTG+b5JvIUMqXMw9CGpWQKgJ7e09e5SGkVzs64oR0X8
OI4B2Lixe7wlpE8SDM2T6hcHtDNGML6/TQnfi1doIZrTZdDW1e9W/LfC2LlAXYZ0Ay9fiaJ75qGO
PaXnWh+KjvJ2yRD1b3qY67NI9Z6pg6tdN1pj5j8Ac+oIPUWH1DTGf7nlk5EGJQJrMR75cBJ2Tzxs
xOLhIy9hHkuIpCOwjg/kkBOcjTL6JtoFaHrg7VS0HihTvH4nvGbMuDlGRykfWk094cmsaaCpSaND
U6eHJVjp1w554OCnnEH+ouhQXY8mgLpnLTwS9wHxoCJSihuemL5949krx0KjSLafARRocxB5sLZV
uNif2k78HE6eb/cjhgHOZcfMzE8oqRZTsK0E+XCvULdEpxrQU7qeOcvlWhGGIhiWoVopGdyHtpBO
2zTDknfKQiNEn5O2Itf90dDI0VVxjhG1/YXBpm0rdhBwLYmswSKJmPzyxC+L40B+4194LN5Omg+j
NG8qpvghqHyJRA/EiOQCEM8f0FltVnToa0lNJK4a04qkGEEm0z6DcwjUzKEfXlKF7ZojrcbCplIm
20RB6YZsIyZdQ3v9NoKdgSLiGoDVBKBIXo4sAWbH3WPa1oyyp7Xxw0ueWS1cey/e6EOHDJokZXtH
+wpVIPYeLVu9bsYi7sO5YTqRYUD0dHqR6jqTKWWAK2dy9YWz5kNSf/r/Ghcw9XNy/AZbA3iGD7Eh
oKM+0CVDQHSGQeenGlEKHCg4gkv7qeZOTtWzcsnn9Ph38U4t09zoXhzill7n5BjGY2oYGPsmd5+g
q92hC3GJHxR4fJ/UVfcLBp5YVTWku3TFSWPE1x7lYrm6fR+2szjtlkSg5RwfNrhw0IhK/QrCXkuv
HjYTQDSzMsp5BMmeMFGItRHEp1OQTwG357Cc+9RqOrfOfZkrn3Ll8QXOw7C1gGd9dz99r1eSK6MR
JW7K/sP5N2lDGEwRh6tYhcmD84DIFU0pCue5ovsORU0uSAoE2C/fTwuVuFsQJ8O8VU7rbw2VxYsF
XFD8DxSbW00WCjhizIHsExdra8XxHRitX2+TJ+z1UOhW2BbV8SeLIM3lGvz6NsVFTjTp6r0VEu1N
bdo3msMnteCj8h3EQ1FXgcZEl3cwUc7HweQN3MvNzLLFKmjkOq+42DBcypKiHZC5C1D3NTwt2E1J
aqXCVUDDxpkI1btkKyeHKv7m9anv1kzv/nsk3kruDGlRLzYSUFDtgr1YDLo/RM2/LONjBOAF9CZ4
KxzLyRKMCpLa3gDXpefXVOsY/jCOYazE4QEl96wljN0/oY+wYZFfadfnMYXYFrQ25U3UK9TtraIY
cDedN+Z6QSaUgtdt67XpylFDPiERYVZBiPni4rVBBpKm0CNp2ExlP+vKVMe19eyIRkR+8lReIJFQ
O+GFbS47VXZnGSYGSId/NdgycvuTdHJ2WOBg3yepw7fJAMZ2AshE6NqxJtQne1RGkMXf9Dh/OiJ2
wRNTLS6/ORxlKJzAsx8pPaoU+L4Bftfx/lzdMotHYkv4a7m23bOvhZB97yVD2dCg6qlJTSE6T7LM
1dD9IqQPOfQrGdRIvydIc4UgT7mHTc/AbQoxZma9XHQW3Zq3nr7SDsfKFdYfjlBK8lQAfVMpFb/j
XSPwevkk2EdjdlyXY2Lj9LSrLc2frF9GgvZ46yi/Dy1+/LDT7bATPzF1aX30ncR06CJWSEdVyYTP
eIgl+XmTSDblPWxQWKfBhfwB8vL8cU83aIDx7At1J8a95DbssrK8lINsgcQ39GuBx2IF8buac8S3
AhyPv+j/J1OWFUfG04RhIJBot4+PwsOevtBFgAomQaRN4ugefKrtDnzjwFe5TFrLq7WsJdn9g8dd
WlHY5xftoi4xbmo1XfgZ/jJVrNhBj5/JMZk1BOTaJUEBfilqgZitt12Vph2Pdle996krGgpBkfrw
4xXgyNvi5UBxLh2m+RWLc/cFgLUnLYGEFsXz/io1kf1ikzbc5swY8SPhM9YzXTZ6liU05ABKwf9v
XFIJyYKf8WnGvnmPDeXggJ1CPym49evTNwf5O/KOBjDDZNn6j1EV1NHFvPIi1RtYCOxs13hwuBY2
3tu2XRnDTt1UX43QvDW+DDaYkVmikCcZmxplE1kiuN5IOetGNz6D4epAsFT8KMJU45e3qXGmj3IJ
/XKi/q2+RdK1eJ2sY5XvuReKZbAoNjsjWkjYTQSi3yA7XoP7ry5Q17s5vUO9dpIXqDXNL7X4I6HI
iSWH/ZO89RfBPFJ85lZvkSBwTWmULfQGqH/lkR1osF9eKJaF4QHbNnoD5PA3fTxtoeZe1sRfIgvj
StcKjYxQYGhvfCBmBuoCYwy6TPHnAJorGWPJcZpU39IEGqdOhCObG7GvD6tZAjNKmb7Jb91w6Zvc
JLne2MO4ov8GLl1ImKkOWYw5MDkRTpl9Nl9R0UVbCgMNR7VIOvi2IQtHr6H6zrWvB5pzROLV3kIS
RTeclYgryqvJk4Tus0rIhKJOP3D9TfxhawkJj6kWXVHBsuhA3aIpPkCLmHzKjba5J9BLMZ1GZOYB
h8PWOSoFTB2yW4l8EBXA8Z2eIUWv+2RecTxGUkBGuAlkGYZD/g+kkFM8HHm27o33+FkQQqOuUNO4
NeGMRJ7qW1kZP8jdx/h3nnM3fc17V+1D9/3oUa2sRjiFj3vNfrHVZhDEu0zUDsFyJMDBHBzlZ+at
ReBBtCytYunrrblyVbrhCE4DfZ5E9ewYenqvM3DiLE/+P+o4hxIljthC48qNci7kalZ0nR/mOTc0
2V9od6qP74garN4FqwJd7g+CppWKhCd48N87p+ZA1/gDD0g0Zma7IB/r+KxUqcQGutYOKhtghVmq
AVUji6LoGn0Rogw6/eaI761eXsV1QDIpYrkKU/OemHVNHk7Ha/6KQEf0us5vx+yMwYzosGtdcNl7
4bqCRfULepDTIFkJqXnGC+mEZ4tP02o30vLEq2+qsIAqHOyRw7OiWQ2lj3oD4ktXfqixhNUg19Jm
XGkkFtGvdhti7sdbkWIlU0nAIEDt6N1K3jOhwh8Tkg8vhnd1mVDr/nlK0U8ParekZO1ArfqADhaX
gppK+WF2iIersLOP6LcmSf2lEoDpQojhuUH7mgs75wmwAHmcKBvZ/izx7bDGxf67c1eEEPZdbAhO
hRBZElyRVAp1yc1KlUUkG6Zab4WGLrXH9Cnx2x+qeTbOnLm3IDsQA32ho1auCHgta8q/SN6oapzp
LdzAJcg0hrTbWIPnQYkhZNBB9RJJ8Nx09A0B6QY+y2Ip3mzSyoozctIKL/SBDVszoYtcb8+dQg5Q
hhvGavwimxd+SjQ6EVLtkPGUD0ucv0mBe+hYgCGMZ+Xhd3yZ2ywRik57bTk/kKkG7Xb8jOXpKX5D
CdwXp6v/qkvVXHm+KNX9TrDCLFwkUG3EoC0EJ26QUdxfz2/rQLi0TbPsJ+aFuOjLMXhd53tGKO6M
BYFcUmufut4dzY5Nk/xUZ1CJIXngSo6TkOBPfgTKVjpw4Hfa/iQkR7O8avjXzevBXAv9vSQRVzMQ
X7GCT80bzoIbfqW95r2DNT2K515H8Bk975zOFjlXLgJesr9aLE9ezB4x8zxXwCslu/x9VBISE2Y1
h1aw6hqYRVAEkBqjp+Lr9n5DyN7XDVF2B5HOQFl0sv5XQdr+rVJyAUfKp8dOSZXPsRd8ml6ZOtQw
vh+gChDDCb6wVB6DhinJmhQ/d+Zf2i9aNG5Dl5QMBSlR3OxTpjk9XWVsBBFBkXY4EyA2yV6REwbc
w3h2dqTLMmU8Aaqvn7FRi1m9JvtNynX7hEaOZJAN0Paf+QUI3QePCTu3KlBmUD+/eVN2rnVLIdyb
ArzzJt//kHlipxRk6rJ/As0/MlxvN20g0JfJODKUHeryFqR34MIZ0+fLPA7jWcFys0VHEVh/yTbv
4Kt+nZAYcGjX+zO0nqZPLbbEgynotAU/Oc+P29oF1IYjn79+QvSV0dozdLQTYtfekylP+fZL3HuJ
AewcDl7RmnfXWQ/obd7HqBuEv074jW5Dyo8cwQkssICgHb48BxVDB6vS6Q2M2HNhK/D4xEICpvxW
kvWhfN6jWKg49DJKYsMGa6fbtEfy8T9DV/tpLurpc/nvttaLZ6ZRKob89zz3rGrZS8zC8sMoYT4j
dulOS2WmFu+3AS5bVDb1N1iyWmykWLANorY5/7/BwqrhNY2gFSOPs1dqWfbGU4xHz33d2P65SESt
5MstD1miKGeEASoyJIcvXGMxvnJ/U7XPFYmTFhXkN7bGJV9W7Yl0H4Ach1JoeKQovX6+7ZaWKqdG
dhH5lnDpBOgej3h5g9H3WUMJCoiv6Yza6KV9+DnaNGF7ZmPpRyH/dvZWp9ygFdQLO3G6VN81Es9U
CSd15N5IibAWU7cVnPP5SgNa/k9Y19btzhM9hSvvI5955rI6Is8UG5JOiFUO5AYzwEafGabmmGMI
WOMAlFJEa0PHC8oS5MWSH5RwIjnemi5n1zSuHCA68t218f9HBjaWbwqp8dziBMuF4i4nwrHZP/Eo
TPzR1SLZt3/dhdxy/3B14AC+EEmQPs/CXMO35+4I2sMvg1wHmE182EGOG3WfN6dkTeAlfvtCeTeL
NZ91FI8WjFhuotqfQMwWXBM3dPoLaolGnzsNKpUd4QA6BR6wee3gR1fX3hqE8GQ/Do2/tJVgosYX
jAN1mB5q9Fi5u3wWrWAHDuJzb6SjWYgR9Feoivw0UGLADaxoDuuWi+OfOY0yvx+YIGgaYulNl6wR
04IxAqubFgGarXGj8SD6u/xca92WzI/AMDDpK4PAINidUZICSOE3bzyjPql8y2/9pKO014INHBT1
a8620PumzixQS5tfSnl8+Zkj4fUpeRIcw96RQV/hGNTLzkdZFRef/F7JtHmxQF+PjQFXeQauhqXW
65EDQRue/t8pzRH9btCeF5dcjEJG08C8zNfuh+ow0R84eouNdndDpVNqEInvLniJydheWZhnyeuo
NqfSd27KOb61yNVumA90olUE8SJOxnd7Ftn41Aa8z7clnuudDHEr6kFIHc34/x1YBJ1Few1CuzsZ
JHsAfl1DzDJt2FYHx4ZPx0hHksYctv9CEekEGCd1xAGnzGfguQL3QJBjQTGg3FWq3wz/gjumWrOi
qk5Hh/rJJXQcuLenxaABRPlrFF1oCqPdwDrifR8wCNj9QF9RKRnqI40Bg6hJBcMyapgACGF1v9tM
YZBGNgFYwR1JT4JJTC/IZza++wyzuTrLhwydQ29klO7OavEQ0sv/D1Ix2befELcMaF8CFsD0wTNn
HwWGop2v+J+34u0NWZngDUmMja5G5D8HEVOLpHoyxhx6IVZpHndiK+Sf4WznTFRKSU0jTECxjSgl
4hab5ws2JYMEuZEdY4q9mTyqanRrGdnD6saMEYeJBYHS+JOxdvya7Y8gWpuL/ILZp3EZzjV6UeaH
KsCWbRSdQjib1DVPrxoVhc6WkznWrziSWgzXt6GiENcT6k1J+kbfA8t4s+vlwbzd00HGg6IPDgF7
5wca3nIN9uf+dAIl8KUdvJ7vbE9BUY7+OLWaAJfUMyStO86BIJrPqIv42zDXVN1zLmgpBpminghQ
zIzisXufG3seckKdFrNe6f41TAlkS94G8cg2UnvUJ2/Mh9DDkpUQVih3gxM4MgCIsuXKjkNKR3zR
0AUgp4OJk1MHnzUwgJnJIfEsV92pojUSTebvceR6oXpPUmR6+N0+XkfmpqSeNwOvhgz482qYzcdS
8CEf2eSizZ7h6l+gD4fKNfzzvy67ZNvMFpxwbh/zLbFng4BuHbSgRplOAd/X1jQYqxt3q7AIiNzo
9nRkYQpyBrPKA66fZostRLEER2S/0K0BW1QFfmH3PDB6HwoEHrf8LI7aAJgIOoO6f78vzlKZFIfX
eAOvRDl2E1fLfFHGQ6QUtW/7mAyicl9XVgyv3KjeWPRahB+A20OihV7xj12HoqvF3x1si7UUvLA0
RbpmeU16aab2rAmlFEDhP80Kq/xZtqkM0EvDLDx2g5XQtIXHkzxDrhQ2iErcCqAIun7mO8yGX9Bj
BkFZm0S8CAuWYD6aS9OGDjOufa6TdwEDKTdHEXoQZj3hY1ISN2cs9s8Sr9dlvHe4+AXFERkLzGHu
ZyDRDL6ybMqS4Ut6dGyrZuY9ec4lUhaFQ62fv47u9ZtDu1vDcQCe+dqvwNjK7VTf6PNPfp8dUtqb
lw7Okj33WkptdvuGb08boe9eMhxzLDJnwqzIPgxt2l7yIdphvB3PJ7Xye4CNz5fjNAZsd6anJbkp
9FtB8D5StKy5tzk2aBMd3xg18Bhe3o+T7PKS5WwZzHUkuhfdsYlJnPhGnH8Y59d4E8bzf8ivV7Bt
cwr/mQtdlTQ2ppOzjdOtW/oq8NFXYoDihdqQUB5RU6FwDzEhyRposJ187H/ahzgTZFSSHgGAWa02
A21PWkTHlJ7Vg5grzM+y6m6jXGyACJ/2Xqt9tuMEziRPhbBa2AIyy3aYHxpHGSKc7lqzJjmmXLuf
3tFAziabVxFR0NMUN0Do7bPloKRsqMOB2cgho8Sn8jpmNoKO4D0RAn5zH+/iA1Q9EdsGMmwiyPxO
uSaUI+Md1KDGLyj7e2gCb2YTpOedmJy5EJ+LXH9RsvWX94wH4PqnHtgHLd688Cibbi5SDYbeDUbR
CAMBb6i6jYzmY+heV8jj/dx3gBQnZ0+QoCTxZrXLa/c6HkDgebEKz+ZUEqgorNRaN2PrP8oxjzcn
+WAfNV8MqHDWSpm9uicOjb9jcr7zUhfI3bIRrGKR4IlT+E2LbqcY5pxXCm7EQogJJnOmA9Sm5t0r
8ogVUMKqYY1b4G2cN27fy+i6H2keVAb0BCTeXscjW9Gk85xndJbgGq1XgzavxbggIAW2r52T+FyH
c7gdvwiuoDLh22hIA7FfDSgtezNznj5kmma64P/bpt+TmMffPjSJK4Xve16A9HvOedHWAm9jCkHJ
2UJoKbxMaTXs0fWBG5hP7aP8OcpKHkYeSmIUgL0rTAHrphlH5k76Zkjj19OnRcTMkxGsPXGjB+1f
BrnPfu0t0GBJE3Qaha4Jvrmd+SlQBKxgJEhuuWmynCE58HqOshKlxE2p3Vl0FcaZYE/96+Wdvb/0
m3ypkEgFJ5gQJtPFdJanLp78y0WVgpxVVwgfi1HNtByQpbvRH7uKMjXkE3LAON0ePackNKwuVsmm
yS0GFAR0jQnspfHz4DWg8A5RuP7ZjyYA2KYVsjhpmQKqjGHGReaarM/Fv4VMX2Cx7y/7m2bJLsJZ
2RNcV7ewNe0ES7SOYFFiG+ZVc6OHvc48ktWYhpSV9icBtxfq9Gy9cqFYKA4JOqZX66Cmmz/cENZE
1RPdHcP4MVEds4OS3/7ROFlZFQsnwPYsG2KJdHhhdD2bvT1txt0DZNvG3BcRCqp8xuKyxO2+AanB
p8wN1zMp0+4+hfADsv91jRZZ39PUiExZKbvxsKdai1aC7L+XK0pdoYyBEPosvt2b9dUqD+Skmzke
0BUI50OXZ+5248Xggj2uxN+tPtxfGmBrXzQnMkBusmBgBvbOi4M+EAHN4+Tb5EMVgQIdZUhK2Jg4
ALqmkRomB32o8yGw5JDYW7tikOTvNRYQAnM32fkokICkfXJeFDpoAhZygOHyXYhLsmyWeBpzEDDL
TM3BexQjRleboJbHuRVMosenQoh3G4N3t4Gn8VX5Bb+n7n3pwPY61hXY7SiO6mhcOxM0cHamPUnM
53nm5QGbT09Un3iTUOLMRN0cq1S3sMC4uKpvxEeyl6KmxSvc00/wKjVUfGNkigbEC/wvdXv5OG5j
utyqpQem6C8k/tcF0byK8kK1RediJ32wUAyOqWjCqXMVQfoe69PqMUZmEMP/ucJuy4z1zWdaGvIN
JnLy7lqwOejVl/R0B1MGa40y9hlzu7iLmI2j3Z9bSg1BNLnVUZkag+DAWUwSZactypbzcezf/bG0
10Qbg5KmXQBusuofC6PYtL1C6W1yj4trIg5nqw2FQhIS78GFrs2AguXGbcoRqgzT/WJDQRG6LuU8
E2/7ynyj6FZ2vBH/rKb4Qch0ur5+Ea52jAlN8hRmlvLUJxahTzWx6ayRi2XcLqPQbYGrJCMnlEIF
pI3ITdFzTqsfBFqxa/9EmveK4yDuBYRuKJ0v5avdzksQzDrCDT0vexdyj8dLkVhxKxbEtK/zpcA+
CfJfW0Z9y1OUuidAmX6J/SXOaUzuKcDabUHQGOwtMPADf2Jvv+IGqAGylMOpa/7uvmgFKjUHbUCB
NjvSkh3FTqQJrHGP9Ogz93V/UwxGGwe3oewcc8ZoFaBMkniOqHtDEhqmZcNCEGfAa0KB1cKsHHqY
t+VkuVV9LfbrUFXC4+PRH306QmL+tx0Sf/xGiv4R+Jxt7sWbUkG89SILSdEqkLjkY2ZVuTT5UrYD
lR+m0RyMoxQSbO09C4oefaM2/EjYnQMGJdeW4ZUHFBgrI1tfNlg4qIjHaprQMdFt6reH2KGXe1qc
bw9kBjvWlVDMs2wtlNMwIh6sFuncgUJrsGyOcbw71w5Vmy0QeGTLe59a4cTeJ7E6iqi6qynrAHLW
e5H4hg7vnRAYKezoTMYiGMsx9JR0OCPYuJddiyqMHzp1+d9vxczEhuAk26uENQ/p4keC+5xizLDp
qpKUfC/S+HnJfbTeLNUK6IjKzDcyZt3jYKsVhrLCkkwBiNiQO7nG9OUUX5ir025pOfKXSVrJInNV
okdeRW+4oYMF98gn4U8O/fOtOAv6ig+kJpFtw7CUuyHaxVZQ0kglabXPT2AaQKhIB9ebLuCTcU2X
v52eCwXI5S3a2RyYpl4mtxehp1pidmDfeO3Fhc3VhBWG5AB/v04sS8YHc59YNAtKVbTia0Nm9xH4
Wph5Dcv/8QKrtTNELHlksYNueM8LzWn+lyQSCZK2MtJJlXyGXa2NpDHtj9AUQjvqWjC9t+cl3x1L
S90Y/W+M7LSfYdpAPER0aGWOU2FPSl2wBI6gSOG9PA1GZ02+0d9QPlYH4Pvi87WxqaxAuV7B3oUI
BhNltYyJCdYuO/3y2+dB8J4OroFkhta8i7yQTvG1sADvbiTOYuBiln4ES3NEcceZabvHfSRuKL5d
HLzAa7PxeVO6A3wBHWOpZIKteG7gg8/wRZUxpPk8BwbeavJkOwUZqgxjZI6ff+gJ2nr9jek6PcTo
eRGhPHJD/YAog69Nj2bHfm4c5/val4MQ4Qdx2yt3abpDMta/xZj4BWWbF8hZ2oyRr5by9xO6drvs
gEjCKMolHiJiMGoc+GNGMsy4drZKm12HLRPaD7TotHvI5H+I/oyHE5THPR6OEIXPmJvOR5flVbep
W26dS+T2nBxR5T0Q+26UFZkaEAYrUiGBfvIXMRt4VJKy/hEsQ4iGUthpz0Qwhcm7dNisMARkDBpr
mkWvGfEw5ouoiIa9RZsExvhjicosX7vFgmdAb/Apla0olc36gXQ3GUrmVj7IeZ+0Ac4dvs2y+xo5
sFWdtIhFbZzBHu6nk9vaubWcDpThlt9PsDJWs9Tj9v6abidK1bbqFDnP3xof8EVXUnLtqCn8lW5N
dENmeQXWfIEc1PXVgIGqLmoc0cQL56vDC/HhIzwem19StP2cW/oAZ7RHnOnyGXT10DWF80ewirqb
vawKHecIDYbhNGM3tqk2gsdYSsgK8VygcUbNr+ZAt35CNNuQCMvToy+ClcIf0N26sIOjlaQdt5TB
VMPo5/a8jRYP54iMswZBG/uN2lN4nw7oiih9GZRxftd8DsC8hcUe6PmAC6PViokxp1mCXDEha7UB
EEOelnHHWyJhedxyPrbEus6IMAH1/VyKUxjLXY9LwKI68LP+ZwY+29adKR1fFpI5XNrGFWFl14du
ZPPiGZae2yXXYGfQ6B6e79yq3ql49mxfpTL5gF3ImiU4szVkbDQK7goYtp/CUcYmv2Aa18oXn3is
KlztfvhaUi6zBDPKLDyQ9S0F16N0RHOnvoJ/9bXlFDj9nEQN7Ps2APQcbLCpd1wat6AwwA5ixay/
qeIiq3SOk6hA7vo3EVE/Ah/FYNOrUZwWClwWQmrVmjKeh7zoez+nnJYv1iNrKCuEOMQsExf1yeFU
72mjhyHrxnNZTcD6zDt+cfq2IVeky9cq71lnoHWSxHiaQ3IUO/iqNydI62m1Cx9n/vXRzTVNbaes
oF2Nx5ieNEx3eOPK3Ce4ZroVuMYOTXgBqClyYEogyDpOwhiToGUDJ5evp56EXA/RxXypjnXKBlK+
aeXOqUv3PuWhGjqwKuGmGV8wIHvJ9/B7hE5u632dub6+iT5wHe6JaeHoNQoxAek88IP0DeJp8rhn
SRUUhEH3AgYzF57dFnD1nb3cc2yqIAeGyKTQ4ffhnn6OSHwihNdAZYgLZtDf9VGuLBEaBUyLHC08
fbkdETHz4PO527TecaiIN5Mza55mmXU3HQgbRv69bq+9B2EMSvAwNpLVrPC9VmGvJwyfe29t7B8a
QFnV+mGtbV62UtMHS4+gC6K1L8sWutmyO8UAH3dvOaBs0rcetp7X2I8l3AleE0uG/zd2MlKclaWh
ZurzYcira/4zRI4iDLklp2OR6yd5FzgEs/JFzAOXL8qCMKG9SbqZFTpfQhakqTmlzqT7k522GIvX
n75Qeu6TwsWnsjlGIKqWJ8YtkO8w1t5qebyG6KLKh6UZ5RlxymsZhEOtO4MonJAMUvX/DSnd8GCJ
68RkzLcrL5yESL0tLSaSmWg8YYt5hcI2BxH2mfuBEx1KdUoix9RnvOWjGyVo3VijRWolMglgLmEK
Q2BAVWRm3te2JAQTj/vZwl81iAu5lyuAIJ8fIt1TxqYe7eWnR7ejfbv0f8YO7WGrnvjJgx+HEffs
Ri3uTccLwCjZ9NAUopr09o5TfoBU3ryLjSFVqGEGzm5XICPSqbO0U9/R7ZEMR6tCVeSDExItvI/2
FNnQCapKcIoOMheCPaQY+mntOYb+OG4c8wwVfy1RoEp9iLbyBvTqztwVO9gES98cHvS2+zxMJA4o
S9Ng9SDWLmkzSglSPcOIKYsIrlZRXgGNFHp32mOyUxeVuhUS0d2vakJUUYt5b35nxHhtMKNjkRdn
fdJM/4moccBciOOxwc2OlfDYiFooWS9a5UuU8Fh/R238WelwtwYOrNmM0TozYLtX2k5E5ffvswdg
w/7h29Y9rSvP3gOcX+i414AAe5Rg2MIYlM7+53CNepOWcr0uOXQ9Sv64t57+JR0XnYWWU+C1qnLv
hSjy+gky6S02W5rbvUkqZF/kNVxMZZSM06LAIrr+vkhqRCck+kRNesQ15vB/j52wv/ZtwJZif7uy
sO8NnFBlTrATmRAgv14BkWB9wVkHaJScAjVaZGD0u90ECD1khj2fvHO/kmOtofpl1GGPKLIViqt3
+v8D8FNRtgUuizrExrxczMYqHZC+GLyxtn/hNDq5Ai1D8kAx/bqpg1M6FyTLAMTD1qen7tlwlzf0
JzZJLxPOIizQTUknZGspOvQrLEvNy3juuYVjq06C/OKARXgxsgbIVz4t7KxjV8egLkDWY4HmUlyh
4BZTXVGgtJ9jM3xQDrKncrqu4ZT2cAMPHf2OCXJ08IKNBZDr9L3xBI/OQvqOyPanOHyU3/uXFqke
LUp/XYqR6fTAm9kdm/UOTmAlAfKxSLI+q3RgxAQijp9rR2X91k8X1CgxJyvhWEc0pPJqlc5SKISW
fY3glP0aJibZNwm6zSlg0jak/3N1rHPsgYDf3VAhK4rWnQB9/IlxpCJTxYnjra2OfNHc50zcFzKJ
wEEOrLYQSQUkPth6DGQimLHcPT5V/gFnPZuZ9c28Ow6Uc1QU2dZUBaopBC3o7bbjxVkRGyun2lfB
G9HqToHrMEljn0iBzF75t6Il1kBJ2mk4jCDlqCNiazYUqghMiZTsCXdKOMJbi/gZqKLTenOJkUIx
CzqGluxeue47yNkuNPd4YC6h8+RjbHgxGY2DRHdLuufdrEP0DKW7aWUkk1mYtpHkMRx3tb8Yu/vi
7xsRSWSzdohns9u6oiGX0j13ivX6ACiJFt43M26Jd7Hztw8UGtJtNRLn9PWgi2AfWUxZ5rOpB3zV
t0wFhHe424LPghBm5AW4OpkjlYZP6KWlzak25X5Fr0ehwd2hNDAfTx+vDA9y2dOfT1kkbvS+W6+Q
f0BS9YQJrrMPFfeiLy6T3iJLK/ZMJEVIkQnbCYSKxr2yasZdxntjCNOu5OIVFCwK8xszem6lx/n5
vArmxmFOVSvW5Hsd5o+CyUFZQ6pZCEQ9xYTaG9Fc3sJGMh+Upk8M5vZ7i4gY2272eixIHaI7hqKL
Q79QTR1jKrfYOLKybBl4aJQcaDDLKmVaJMmqLTKTfynorX1eisQ9Qikwsj8L0UGZL8+CzR6LxiBV
6VvEIuLiGTxcNlSGti/H/phuyqvbXbquY8nZjPJt3Gf32BfPfH4+JjHJYCajWT+u3FBH5ukOxtmt
5k21GhsDRQZnCFN7b8aZg4ha9rF9y0KNM1MHdkmzspE3QHXTNlx4bZeKgp3EqNlVHcib6Bi2IaVb
z2qGAe5X0tairY88kah6cMD8appoUjw3f3e7fjKCMGToz30WHII1pKnf9phfq7g1bOY3aCgqzS9v
7J3OaRO52+5R7FBJYkeWdcYbgvAaWrAO3N6xExTBzHyVjoi43SycIM/40vFuJyMpRsWzMexpvSZS
7VUMIGD9yy7D/WW3SF7rSomJnYIQM546z/88+Nx964SGxYZV1AMYRv/WApCbUV9gRr6tbmnklNsj
M4G59bUPJ/NOemson/2GsKaCoVz1J3JIH8OGTJN9YGbsh8KoL7pKWIdHXXxEKJODPQDTy45aVm7H
v5G/sSoqTqzoUsD88JjtkHAqRtW/jRSquNSyhOGdVMBhIUhWdyhC8BIk6YmFFU9/xcG5uIN3arkF
Ky9+z1awKaViamHDy904jMCpQKg/6ompqUTebEa0rLGiGEUmFl1eXQ06LeX9LkUOXvAR/ellpqkF
3+QnIav3CqEvuTShVFkDn2ZtqNKHgp00BypZeXN7xCFxmugzijh2rkZJ05S46jrJUqNUCOcYB54J
jV95ju/w8nvNgWAFANJmoCiBtD19nRNzsETilqFaPsbUrFKJnJtZT7HbknHa2Nl5rsWqUlXiJq0o
CjL8Iom6mFTgfY19MMkK4IMj2NaJArFhVcx6bsedFwvrn+E/kpWcwA2jyBU+vvcmFInVvYzFNKAs
7GUH4HWMy894kw8aPeV3QjSlXQU9jRVTCB7oCx/E59BXQ3O239y30wAzP3ofN+AGoNza5LNqpTqH
Nr2PhS2Q3gjrEcrbnnfqOfKz2O5Em2t5RSQpHIvzc6u5DaP4jYq/AfEykHVaTy04aPD1DmvHhmnR
QrtUnzAmGOvduaeTg4Mml+VcdapUy7PV7UCrtVjfzmp5PenevUbImboW+2BNgmxxDAYDul2uCUBQ
IcBI8DI8CIwnemZhxDqk2cMNBEl4XXNNdzZ+2pKqY0Myny2+pduZZHzUaDf3OHfYuogn829BUXif
0ATlXekZMflgVOK2K/2E4yJOd7lOk7bLFcPIX9mXFjVwwdcl3wWk+toWNAWBim+naQ4d8DOkQr3X
Q79Mn/+I9FLwupqhGaEVcJWRozV79Y9Gy5ZYgEQ/AxrQq9jul7mvU/Jd1iL2L+HUfnq3mHBB3Q5R
665cAJn1wJCXKJqrZiQTsjn9Z7snB7fhxmP31gwl1Fldgp6Z2Y8FPiGdnrxFEAEEULuoax/kLgjr
mo+tB3pblWPBDaKoqp8z3LUFBnbQOkrHZBnennI0eWOfMNrNl6j3PVG7lOOe+md8cUeG0xQCYeZR
eyGz/XqYqASkbzsL5AqoT2dL3WuUMHSnz6Q9ne6TSKSOHKvb70oQ/X3tCzvmQtGxD2kPNc9SG76T
jylHhHdKS/iusE8DsVfKym48F3o7ypIrO/Ol+ZCBUBaP3Rlln0vkXa1ARv9LQIUiqP+b5e10pvwT
korvUAMG18IOMeRZp3/I/Eu30bsMrvhjRxSZ+mAVJcwnHCn5y7QS1VlB6zZmo8cGCRtPt9q9szs8
7fUG7OJcO6Ln2KMfxkjvSZskPsc/l8RgYHeqE5B6t9vIbhIJGvPwVP9LaVuaYYgBAhT9laMiAYLD
ZUttepRBUPxelTq+5+8aUkNYR3Wsf1r/xThvCC9uDSN3iLlWBeXXYHFyf+7FUgTBJr6mVPos1L+3
XjtgAO0mpW44GLo8pAfIei2w9ROjg3VITaLlBsYSiGYk4L+cNLM7ivVdAHjMCvJ/QnggEPvFmmFB
wIvoX9/MFFGDCP4DQulPFzfFbc5AmonlgsqgmtO5nYBKKw6WE1cQsUFYODkz6bdmPsiLb9xVyxUI
XjYrsygyMrxciYGa2gi/jKp947to1DIhOjpcF3xmrHWu2wQP4MHCElmn3WNcJ6pU+UIu5Wd4Lcq0
OB6MwiSeWKAmIEjPJB4CUR9kHF6WBHQU0U2ORJ6gjAPf9x/ZrMtNsMhPJgM4V20vIKAow1RXik6Q
C01z9V0S/hafO9jiLYIxiKUz8VqbsLX+HN38iuoc5kGvSMLKMHo28OSg0micg3Z8H8BfdF3iB7gJ
IkO1qYgWxuBlNOwoXRT2THQu2AB+zyXifGozaUq+2hK8oQa6vYMxNF5SO5QpWPhRRTHPCF+vqqIY
vOS8GA0yQVZStrttqmuxGe5r6Io7QZ4QQpSryZOmRVgmRvPnDhf00WcHnN0c35hJ8UUqiT3TzDci
v339Xa4uvtFvD+gpIRO1rpLbCs6+Zfz7LFWL4qxWXIThSp9eHI6hdLzmd4lU9CLQ0nBwaonDocuh
skmTLbISCnyyZenu3n5kBVyrEBCaHBLigLxOjeyqlpg+sueG1Y7FDHKNgfo2sci16ievgCr+ozA/
OqlQ1V+4Gv8xXahzn5QY1tnO2F4JXob0c96TqUT6uITFlwdSjep1/UhNSHX945o3+PiJi6jfR/TV
AH8Npqiu9b4K7TSTMkoqqHMYwAmx8k0UAVd7lMBh2+dYf92QjNubd+QXTqJW1GRjeSnk9dRavtzy
csz6i1gYrS66PhJk/11ajqE+AyLZuRW3LA6FnxHMoLCWODOoSKH4cNLbdRcY40v5GK+cnNEvGPpX
p4JyIcA7wmNIzvsriZ8ok4rcSH67j+typLVAYyhVr8dhZeOF6VvbSFtb6itNJ3rcfLihg7zOSfbP
h7QHbUgaKJcm1bwknVpfJNlNRkq4pivfHyzdBY+2g/Yfq6tW/N3y1k1pGC1QcVAZa0WlcUCpOnWO
7OkyiCX6yaQHH2ncMz49mBOvdcJdERpOFpoCU8pi37DaOk2YiOd2QV9yjcNuml0Soc4njfg+8+yn
G/ZaJw9wA4ySzNJ+5E2pHPdjbPpYF1tRVyky5g0V9pcw6ZUayAd6LoU3zRo2fu9yh21q4vHuKeqP
YYeNXyFTw+H6PVUn9idkGCeYEj97b5P2Z9X7TWo1EAyRnaiezmioDITl4xZw9MHId6MVbnvAJ8Nh
nLMHQu143vQB7jD5+U6MDKN7LvCkkq977peX8tPCI2WXpO8Z4i2afoejfmiryp5OvgC4DuFHY34K
B6eZ5yu+Lnf7I3v0YAmAo6QldQuBFB/DGm3cSAM0aqn7a61afI7CSdgsIeherAawoKSy6N0dpIBv
MFdT/r3YeAfgvk9VsLiixt4ILOEXcKJ8Or8UDN1eEZQrDsPl5DtsZau3qRJXriQNsjmZJ2sapLsc
zeAUiG1fcIlwy4OVOHuH2ML1Gv5GDE4jFXj28aNx+4ZtR6o1RaK1yFdR0BARLtCleWbDsDyUITly
hMxgqlOWlGr5sbFWq6KSVpQPBsngte7GXWToyJid9PC7QA9G6ZmrGVmsjYgjE9Jk65EghBeFldV+
pALtseNgsvPIUV9f1UKIhXWf40Hg3QHiRlsY37bngNaUK3f/bY6Vgu9Hom5+8XkD4D6CtroqhTY4
1JXa2jsx/ec2jPLxrWXrtd9v8OwV3hsV4gtBhSkMn5w/ZcoGZkRXGy90KlBav84DyJrtfZKjlpUZ
0Qe1BLMVd+bcFIYf9T4H+P80cfy99qIFrNdLyu29Fbz3LBlFL4yHr1dn9q8LuSFDSaiq8nfUNV5y
mxbhFT4OweMD7h32zSXB47pZUKbmY2AK5afZkFeHRYBWIRT8r+xbFBXQ13BWiFxo+nBPARioJ0BN
gZntOD1Ge1k93zcOGB1OvnWVY6lGTdgHfOewE7JHtSG+pXImWe8q+EyGjQYxg19ksCXC3quDHrqS
Ny4OLdpU7DvXqgcr5yj9FpxMpYe4Bvl1ssUqlf7/hTDWMvmjotiQ+HEsZdvTDxttDc6O7NJN3Xd+
c2VN9g3r8ZujuhqLWS4/UItRCNWT8F9Dv8CKRaWA72oBqk3lrUQAgC37M060YU4+IMEpRFN/SRyM
vTWU9b0xMEOJ4bz8bkQtRTQL6dn224ycFUeYsBvWaMu6TcGEyri3s9xwWDLq9tOzNbflM+LMmRR0
OWfuwZDfbWF9eejO4OmAQCd11HHgHTWUEes3GwoMFwYd9CBCkwbv470Zvh8X1A5V9vkJIY1TNf+w
tXFyvb9nyHBcHrNtxd+Q+IQJ+7THWB6VcBeph3mdyZYRvAfsgDD9BzZyNPLlYY8gotK89lQVf0cW
wIHWQMj8juwW9Pa2tIR6cOLuspGeSHk43MxSmQC+8J4G1HELHfzwFKPy6qlGWtMkmTgo9ZvpC8MD
Ov9nvbSv+XcgXxqLAOMFmE/dpsJcVBdkx4im6VFR2hVBWYg00/mAMyM2TPHAnoBA/97S0G9QbDrN
o51iUI8gH8WXMb6rfAsQacllC0asEWxMEF/QNgjjkr3RZ3VD7HvK4DDZOsS07jiNJrvHegGdkI0l
IADDgHA0jdZRRD4ux0T6Q9FO1Nu1FZcMWdbuNm1rGV2k3nYg9NUUlCWfSWxQ5293tB42YKlqhwVC
WBx/39pNShqQdTQYhYn/cgZr9L3YaiB+DYqSJTOhtWN2RN5Tm67XHh/XgCuu7HgVDazmph8+lK2f
JiRaNucOHr0ZTgBPrMUSHfbczs8Wl0XmdntKFUSiYyTPMHU7mVisJj0Z1CumnQRk/po7D+7YoE0w
VejOkR9cofhDlyF67/qfz9UvTK3cHgv7uya4UMGWDLpYkzIHJb1Cvv3O78tSb6q2zFin7fRQ1KCm
c4Z68CeSXR1IofNU77uMNc0o4zw4TsxwWmrQ1vuvjsxjQbU5rORK7qS5n2LDFPCEk2U6FafaDgu+
s9fVbdb2WLa2gM4QJYePD4VaVkdpl7UWGM7ZLKZp+EmI1NLAVna20NbkddrUr6WuEvpMJzzhS6GZ
X0DzdiMeTZ8wMlm6YDFfYqjkbShGU/3m2aOagbntCR2ruzOtQUe+nUqdewWD6vQvXGOKp07u8EAo
VRtPU+VVSyrIHqVcvI6aDumUvWa1a220CWlWfWlmkETtvIsTroba8AOA0+rcbcrxB6MzSaKnidJg
1duVZHVYGg+OKRGz/2z7+Sp2ipIb/S9djni5PymD6BkJ3AvQuzJ9f7myT8C0Dmj382hteNo8NFkS
FbYC88YSFU+hKAmjYWiOmaJndmHTs17Jiv5Ej9ZhVUfazZzQAPp920o1o07/FH/lW8lPpS4qtfYy
LCCqaiZQ1FHkAMkXcy/wCoa1ToE3Jbtuf24iLSb80pliz8Efg9Hxq2/XmI9BdUOmoTeV71U1iA5O
gyTcQb3Wzds2z05fnvwnXCEUXN7B0lDgAn643q+LTRAxadV2Smhw2357cCwnjvQIFi6Sv4hDxoj1
Tkp5iIa8m/vZucml3EgmgK2pZ8tI3ZN6sJAsQfS5qbxD6S887sKCOKqdsLkbC1vUajYJAGxPh4HE
zD+7lxf3EmyNI56OBvSxjHgaJFlEtnJP8x3C8g+nlcoa6t2kGvIB12ndsdvHNcT0xw4K1pj6AJj1
IoQsAnhyy3mbBKBgqRSCdAWi804IyP7G6E5VlIy7eq3JsprCQh5vbjZhy80PJy58qbjwqPl9CltH
cfJlh5yjYrPrxiCrYvqKIO4/xukzPpqA2RIrgLv76Eexf1K1qrAvrSIbiGkNn/nOC+qXEdv5/RG6
Ny/rz+u7fPInbAq09K7jrLNQO3qNVgP2GPx+1dyGG0EUI8N5/pSJQH5obZ4z+KlUd1FKt3d+g54F
KqnGhYsa4d4M2nRwNJS/hwcTN3aTDZhnEsG4Cgcji5j8R9m3T5qUZBmUFLeEP0YnrCnvTG1XAlye
QUp0bxdexEF4Eke7bM7TPZHXhZbVmT8OX55Go5uNW9xF+5qW6HzpCBrAPCU4u/EbbrQeFOmzLI5Q
FtRLMw2UNG1WM+B3siH3NT+lLqKrXkj+qzHKC3M6E8fXsv0j/FTxm0FxhA2VhUidsTPZRYROl0uZ
hmY3ucgBWcm51nlmPDNstrRyuIDbNJ1qwrdEAbEVxgDtScQSY6Y+8uYVnBvacn1V8orlXsoIDFk1
sv4Jmtj6ebnRe0Fz52syfvY8OhEnIMnQVs5ysGcdTaPDppMkqpFqfVzZFO785S7Fe6+LPTs28zfU
ELUiPlNwMmR9dFdVrxACT5U5u63E9OEO7deT+nHfHRwej0Z2q66/uLbQ6+kZKiXZMHgmFKqb47t6
W2V8ZCr/VykHZjRTvrUDUUagYPZ7bRQWgiKouBgzJSUp3RRaZEoHV8+iYtFI3MDyNYdxt9nTUKnL
3iC1+o08RVmIi4EXhwjCudbn8+6mG2Ij6s6ULV0tEzDUMVz7gyOTG9WkZnnaWlToEUVLvvgwtsul
h7S3ZTgpd11Du8CA5W8GeRoHkY2B48nWEZEHH6kfFerMaXp9ioAiILP4lQP57LOtBMYlTaO7lY3J
2MdMFXra/yHuz+1E3ttndIzvYr5wB2o2jBdXoF02k9jItPz1wNKvmivP3XrHwW+bw4P+6Vsg6inU
aGxPGEpdsVZRjlEgefhJNLtDoeTAlC292Ur/hMKJzmKEau+2P+71guYywUmTCPGZ+gR7bZI3r4d3
S5XKxrVibBOZCH0AOST1h4hpUqEX/cc77EIWizIWwwbt+XHMzp0s4hhK9C2rXK2N5jBGAkonjcHz
26X0SkTKs+cxPFcWQ0AtTOioueJ7iJ+1tpAXJCiLTuHNweC9+FYfb/W6AdoM9gVkxYJw5G5W1GY0
ITNB09ZcTKmK/gFnr6JM4lhVmGjJfodeVqV/Y4EIEiii8ICACYLxbNIEA8UHiwdhxNqwBqg73hOB
42JxI7xB6gyWR7pdAYwpOd6m09///ttmwUNkFcprL/h6mcEFA8WhMQCGbIvUaN1/HVoTgOOslONy
+DKhxAEYsuJc8+75SjXcqWuQyVa1LbAfHbSAYHAB1i6qv5GeIrm2h/7yJg6AVoVIIOQXY3oY5tF3
4FpZHw//hw5TpDeOCRDzSsXKNuF4mHV3tUUhRduXR156p1+F864ODR6k3cktMb6Ph0ryr44REZRv
/lRbn6sQnjIkxUJ2PcCBUlV7ep7DxayUt/5IL/CV2tchL5dnjQb1jrBJcFXA8vYOB50Is2Zi5wvS
JKdHQqhS3MRo3Ma6I9T+KihUGNVkXZX1ei4cZoa46SQSXS5o8eCEWElirNhJC102K4WWZHmLwMsK
EEuWAPndRnWJ3tF64ORyGe7Ej8XPdrVxhOWRjAC++7AjrKrMWniazKKqEYTmFs09X73caaw+0ol4
Y7i/Gk6rwzLsV1rmdFny0ueXcw8z62RymrWb94y5lL+jBlTF+s7ARj/3f0qIWVFnOt2/+j9h4B2w
Ea/SmUAuI+5Oi+cqVkqM1JlJkjICx57KEWktwUrdtISIQGhOkS31Oty+WGMegbn5DO/MZynGDJ2s
X3h74gSyP8bil+e1BJmnmIpu2YNxRWjdaKRqgtS6hu82w4bQ7l/Ldri5XPdC8XYdkwUJ/PIU9i0n
qyn8L/xoNjsw1l/8362ugHKqU+YL2auyeXE51yC1d+510hLkSK+0gec0R20+cSBNbwm58iSfJHPs
CjO4DW0zC2G8poapzDIsDRklYWvCVGtaCWuHmEGE8jX5y6+w+g9TVvoCnqHG3dnRjYQAhQxARill
JPmzEEc3T17XqRGAUtPNK+NFfq8lLh32Wytu6Q1yKr9+9iQ6HjuppfskThP3UdvewJtCVkKZbnVD
vfrHykZ/sn5UkBhqPP3RrzPNYWoT1whGrMVNm2y7FeeJuLFBc8wJwFIB1eWXd2p1NG/kvkWUTI/g
f/FdiXlbNLoxipRlmIbFF/azJXFM4KVRIe9vxOM8ol/CkIwORTHfnnYj/+sU9T3fH2jL99thgzwy
CM0AhZ4FbXKBD80EBABc+v2+5TVyWJ0mMBTHJbHba/X/vZg4DCYIPWvb0UCP8YJj7jvCc+lOm/tA
8GKAfkNagpIwXEw8mhCc6lW5ObGmj139hgFb277JKu0151ol/agc8UcC3D32jObjxn6oPTWdJnHY
+G6Iz6/6Vhc2zGwTm4/tO3TskbkXbnUvFZFS8U4P/CN4W1p1aZChhKNJZZLvhTR4XlBYxp2m/Lcr
wh78j+0lybCux1TCTtKeYAr/WddvK4eYF+NH9otuA2b9LCyY/EyRkczDHQ4s7tOpgBef+XC3OmOm
AZha3CRfGlYSuUmp3ky64Ul9fgpbgVHUz6c1WDZETKaSMoD3WiiyKfVYUpwBrkXd5nRv2Yf/IRMY
t+hsAJ4wAawqtcUekT0k2FHeuz8SNh6uPyWktHejnKIwIafMElPTwgHLZYGUffLh4ouUW2reuAtI
nDFYnTrjjYVuzqzl19slAAXCu9vQX9hHkAeUidoFTJ5hS/pS5OyxRMQpmHDRZp04UyyLs7CS0Hlg
dX0amKlKS034geOQGiF3OE6MJXFxly2giuLbKUTkyd+poZnfiyKmCyX2O35TSO36NEGOTyIRfxik
ahlOXdIhNGdGPQo3fC0J4Vtv3SA0oyhedGFUnKNjuhBVQauEGocOWS+tOLCeE0LnqspHD7DTDmXX
siLP7X9pauzg9NEWiG+JQw9SOpk+ziFyB5O26Omf1o+TsgUB0T7hVbSdI5VBpb2vGdr/1a1rPTqf
l22Hsjoyn37pradickUEeXXAO9lOgktHfpOmfnMpqWE7XBLhZGQ+N0Cr1OS6nSwp8MFt3hcrT2D4
OXuKMza/oswqhEJtAIlVoknG6dYipdsGNAGqKQFAni0pltK9BM9HNS5DLRydp9igit6VHZn4NUlG
NAd1q6eP0ffInXly5VFjip6lV/4M39t8R11zAcGydmkj2h+zuwSORzlaK7DstTNWs+dsDLSQM9SH
Ra1K1Mc5ML7JXpc0C0j+gXCzhCl4D3R4jos4Ep0M3m7sEMH8izphoeHls2rG6cmYbb+S7XL2zKKO
Rp2yfg8CTTbo5H9zaHVcn+NeIBVYklbmMnLSqtKtA0zjewFdJxrW0VVyEN5qkwWuwVCkrvlBGxJx
ij3ORvrpF++IEe1B4G+gd9uud0vBmL8HXGknnI4V7rqaFezyqtGINaBs8ARjvAT9EeJx1T5y9YDG
JEF/AwPXBEUI+VaMNjshJ/cdBR6cc4t4OJKRiviAGQTqLJNkdi1GiNCBTlVLkSw1MOJIo5iR1J3S
Nka/EEtnncOwr1Ek9KzI3C+Re/96wpgZZosjz6kokjIA6b0dzJFBCerHNuBGdrWCie9U2T1KNrlj
+toYzOr0cewKyX02fm1YWx78/nFrQfx0FEWqPUcMccDtLhAFSV4oxFBBwSPV/DMGet52mtPjJ+4k
FnuDQGUJOu+wihi3mD/3+u/Uz7ZuDf/2pk63m7VN+g6BmenL0nCJfZ07sVk3QryhkJOlZrJ+oEJ4
A8oYDVkIS6FpRihrapKDNqvsyfKobC3spObCkeFf8YTjjGA0Lxx4FQbFPFHDMU7SjR8oimJCeWn6
RvtA9402mcagqwv1CRfBEo7Ta2wKkBAFrxqMz3vuB2WOrydnECLGakg+Xc7+83hu0guJAm/kVckI
KgMcs4hhoPTIjyXuKcRNnHOjFdiiNlLBE7xZqP4IWlIAfEakPu4KeXOS31lImDfYyJnL36QwEzmW
8yHJFcN86nfFJxco/0jvTv8+sTba7LYMUpv0cgB6QdBvtvybOyTA/Ghdednx7DZdP4YYTxys0HSy
b+M1E8ul7JU9Xbz/kNweeGZe73F37upgjzSr7FE9k9RU84JwagHbOgQ5OCeFszIayRdsILK8+qXC
9Fc/jFyaaWLStRYYFEau07FWLU4uUH8b+7uG5EsfYTnvAN58RNmlJuTzLbHbxIRvRn1UIZtOTDtq
PyKc0Cnub/2MfaBUYsag+59uWMiCNhIp80NYtEwzPu7Qj5OFx4uG743vJYHOjT6esw3KQ4wARUqr
cmjsWjPYyh8GHMCjAUeMJ9x08oYnjkXarPh+hTvq+pzwrVl40mXN/A/mSb6+3Gxd6WXtHtIa9LmE
Ng1mHZZY+44gHS3vwBx1C98fznPqNHcKsq8Hhgl5sbTY9bXmyK/kNhd7EglKE00c6roj0jbVvzk5
nRTwYkrU2qGvuYVw0DdXk9UY4M49PCwR8jeIxzHS9uSzaIAzQnzvJxeEv9hXtjJ/kr/Q2dGbobnZ
PsvQzNfKL5S/yNo8ym0VVDQzmeomMBwKwY/KabYwslqkOTG4DYM8gRw5mjJ+LE5X5YSnTS4myf8A
CytMiSBxSDN4ToBh373CqB+Eug9owfEG9E9AK4R1FuagHLvBI0d7cCmx6IrUx2J6w4+ot+VtEXzW
o97gZkvAQ/e511ylSEcPTsuhdkiojQy5m6x04bATk2WqdxC8QgiL4fmnXB2Iix4wuAq86wakREJh
B6AVVc54E04i8cYG8seiknNmI0i3TeLhVmoCippNy66y9lTpnOvsErLW+Lb35yEU+aqzB1Fgh5xU
W9dX29sREBdjW8YnsX3TweTdcLEXun0WTEFyDbBAQ2QGBg45MbhQqzaRTZdc2FzbGTVXEjghq6ZX
bNyTVxeyZ0qhUC/gp/bPhAzFagusM00Cc0hjZR2uSLzTi+h8R30sKP+AI2U2Xay6y4XEWauV4lpP
Bz5zSt84zY/cgftKqayHYw0vjCm2CCijTWBmP6/6//WURjmEtz2hjUzWxkF2OG3pza5icPM2oYVh
vs1Kjhqv02ArZph0Mr6PH3s39ojWpjBroUnc3zSkCG9sqjw7VoT0dAmEDcP4vCKVb0XG18yK6MmG
L9MJ8ORqm0v52VC0ug/itTErdGq3Het01jMneu3YCQ6MHMfMkFp3GH6Z0my5VQ5sokjXRvB+hpB8
l4soUboUyi/P4vWQE7ZMrUmpWLyMzA+Gc4svmEDLUoa33bnxqZ/pWBU01QXPAvyw9Rjp4R3eGGtj
FEilyHCyQ7cHvbspa3V8SAka9uE/9RzG4F4uyZXLQDU7FGXpSxoLJLGXZljXokLcM1Tk7avgUcTv
gP0E2sdCaG3oYg6dXvKZS/fV5TjIBXqpX4EEuFgv1Ncz0qER00wDtPG7Fk79HLzlhwxAcsqnpIpM
QAC8XTX27qgKSkwMyZfE5YNmex7Lj5vKmGMLkX35ANBq7+6/God+QJDxHfpdT3KvZyMHQSIRmij3
neRiXjvp4CAFGt9D4dqHq9h63RF5NulZZdfDVaLiXzKhr2bnX1wERdGVYrG8kcJhlC/MyeNSWYnC
AypEckVOGDe7PWo/zUlG0nMin+ZblPfzkf4NIgLJnBhqqiESjjkKM3xrCs79U8K0d48bzImH/Rum
AKuFubqx3bRiMPxJlQz6VOwyrNEoor+Ssn+gnmtnOuDFOPb+FUiLNnVuwndxK/2OU5JJ58sR174e
OTYkgSzSvJy3cyNnML50z8HNzbcVjN/ffSVTFFD9qenwNqb7Grv8krajzxfsnpQQQuT+BXbYMZzC
rGNdLzRyO5GIaSj4jyUI5cMIix74wSaakTcBqgvqmBMFyz0Cb9/x/wXn/kDzGGSSiIWhZlHtx9fB
3mSXks/Z/Xi8esQ3wm2lKg7iweDKi2efeW+SlQmRL8OHtx6Bf9Di/jJh7SWvRyKs9YleqrwaiY58
2DKfw0DarTL/Z8DEp4RpjR3E63cGxwAIMFEBryuJw1j+UPicbtwjvRRSTzIJDFtJQMl8iRqUyzJV
yzfxpKvq7WroFOfS+ob5dyFw/WHVk0a/wqX9RLNe6hocOs4Gr2ei6OHUOPCGNcguWpY5axEZHcDs
eAq5BIBkLXTAKfcF6YBuKSKltzGQUoDVw+zji1lWrXksQ+q81PoXXDLec4HNSwMx9FX0Lxpzvb2c
fIll+j/kEw0eyda92sKt5UozEh4sgajba/GpPtENUKxNW6HC5pYkXyQrx7kyA/Z1xLdDvphT0VSg
Fqeppn1ikEtxWfvKSkAXmi+sWMy6EO/MBYRo8zVRl1H4L9x79b1RXKBbug8CjppBnLDOiiTWCxhl
5TO9q/jKCJYmFNp9VBRWUmLU3g4yEH0dOszi9kyPl8N+qjUvvU5cebwDFCEBZKbBhRcVXJGNsa/z
d86ca56M6UDwTOEMs2Fqptl6QHAlX6COR6p9N1Ms7QdB1IWLJ7GWBam1YZV7nuJefJMR50q/2a1D
kpDjT92Glya4PHtSMwZhVConywviNUlg7vs1U/Fp5MPujJtNlL4BQGx6ss+DxPhSSKn8JNxokiId
IAjsETT9NasWiS+fOMpe6IpsqE5bj7r29QnouVOqiBk5QX/9c+lNj+XXRzQctLjSZMmKCDMhmilz
T8+1xtwcCUaTZRpAopPNwLL3ElXlWXEFMcCSW5EOkrQbexKZTnnYWSPhil3LeNBBiL4eHMYHZdsz
U+oUwpelTbgqLCqSLvm6LXVDIScKsIWGDfNVQc3/HeEcTbG/boM/WHCFHh26l/cjD9OkNJZePn5C
V34UJLw0BQypIjs+Cqm7ptSx1eMHCBXcxG1v5t03ZechnX76OgfauY4/hEnr7Z6X/BiEeKLRsLWn
jWKXGR41+VAxSjsbV2CZLara2WMycRTptJL2o3purjSLc+Jr/ZOpFuovJl0qV2rdQoQ64Tzwk5v+
FL/1yeUMLWrbX7tJ8ZXqLqIakTTFZd8u+t6eGHRx4mu+qjDb6dhSL9Szm+eUckbyRQQRVCOGfgHU
Ti6VJzDUfgCm7IHwvnettXgGjRXzkphRKAO2NQZOXBy9ZOlKKgYf76kPBuur0NrHC3aUeX/WdZ34
kHm/UmgNO8jLrWKSNvDQdJ5/yuldbS/OHoRZXirqnGyep+YwqAuLh9rn1jzyCPtYSNwiRQVSP3MM
F1tkiG25bqi/eia/JuVivBiSSY5J3IjDIidO8WWKqwUREqHGhG6k3UuTbGAw5AzCBeMmz5E+0OTt
5xn+5+E+UxZyw4OFMIm/tuwnC4ecalLDOJ3RGMv48WPhHxuY8c0y6qGz1KVS11tCw7M6c5Bjjw8L
4xDfVf2PzkOA3d6YQXKbcJWrZ1KRJYNOv8VcdtjHp5tB2vPeAGsc5buHl/tITB5G/H0Xl59044fK
wd1MCGeKf8DnZS7klEWTRNaPHU3eGb1BT4k6ulZjVld9OyWT+qol6ZS9EnHIXYsoihiv09Xw6zBT
GEKC7CDV/N9I1LsDgA4XA/23sCkvZK5o0nP7iIB4GQ1Fb+nc9LREfV2ZD5WMCd4uDUbwkJqaYcJ+
K4YEaCqhYBQ2YydzcunO1OKpNyohsM9qnqcrA88sZYqFO5X+FmB1C+6vBb9/MYRH3dj2akBYM7D4
ZICPAA7yMI4RlxSZCzOrWaNYmsdN9ZSuimONlgzGA+jbSsGuLgcakxBGKYr/wr4jygrdurx/jhQv
5QuZdeq5at9miO0A7sftnZhppt4MqXvVmYwaDy2YeFraQ6h5iaV629EekGqiqW5iS3etKLNBJUoy
NK19SCMboG1L3V6gKGUHDy9f6q5HdJvVLVEhq3AWSG4+S0EWUqYHAsirVrW1Rqcim/Xnovi6skw2
sN+UMS1lqU88mhYq6PzOyqeUps629l/hRcKgDFvwGpdpf1hbVhDguvrfEO/+s6UZe2C41//nlSu2
9HXSosCJNRSGTz11YquA1J9Xg7XPvLFW5fyY4qyOnQ/BiGJHJaJ5/WRSfidscQurphx4wIkOPnZR
CvzRUm3Ealsrd2aOvXIn65DvBlLhI59528fIndtsosr0lhqXrViXFdV+3/qfHQyhOUAg2JvFS7P/
cCzlVCeQJR1/DDPn1vOy2kZe0zlA69KEWcFliRoPYtYBGb1lMgZ+PegaeAzw8bo0cNBTBTluEL8F
4Ek/HgCoYDJ96KP6WqXevRFR2fW2NHsdSErGBl/Ub78/xI3kfaiUt36XNRRF8YuJRtwH/zBWW6Zl
7s1/NGgD4OtHAH/VtRPvJqgQZ8pCwdolbRS/d3VBULV1wAImWVTZb+1+1zWJRBwkKo4y581EiMdh
iTigg4dVqeUtOQF8RXpHyTwX9ttaRKOOLLbuViXVLR25sy3HmvqyrcqX3EJBxtRGDNt/oS+C/jYj
cwQ8Eykoex0gEiufd2KLB/M/5Ec5DoXLaypnmybFcNlixjDEWgo5lHG9he1qEfca1yTgQ2KFWEYo
pUREMSoaAbsy5PTdRwmmskF2VfPPdqUC56qmmQIJmyZWtvyEJbYn0BzAlydJTOa6cuYR5hHHXovX
TJkWNpx+wmSohj/wYj5+1mfZbXQo/6B/FB1+beW0Ja9B6uS8wFAOungI99/EQqk+CAzm2im87cBi
lLpmXNCQXPivdsstdN2g0eX5AZyiQzVWLPsyuLnWhBinq+pPpgYkO2phlwhpxypKYs6vGgUlyFjA
3cA7zt0eOly4QC76xp9migIpOCqS8uqOKqSCW6G4FbSy0MKcEMZJig7tpMIFXgIbIgihY5YXBj/f
KF3DIFdD4U8jeeQ7W58A4krJ4pwQB+a38TSfbFmVuIhmD1ZCYJJVsj9DFuPHK9ooKu+Jc0Q+5ycL
c/inm/S9USB3IbiXrGqYgqVBqJv2zNgpf7ZBp6P42Iz24YsPwaqits/lqOH1Mt7wnW+btR6zQxKF
mgTBVPUN0XcYhPRAc4RpigD+buA8xhzye56YHyldLl6lelDGNJNy06ClJQknn9AfZisq+VoLyfUH
7jW5nDpN0226iDfObf98PIS2V895NmyF+1fc83Kxa/5DbPNa1jlbD8VEylKvKzqKDd24K7fZ8hIX
v5Mi04C8DqcrtWpUqtcz+CV0GJdTB5blFgKvTwtpMLRYUirisFin/QDieNExgjnvYeVlQrCto1st
3JApUe/QL9oaP01yOP8KELk/4VmAzQJdtWdZlXgB8H+0I3WPe2rl9P4bVbH5naWSED3eOEDtSVxR
xNg681t07XkICIJlG13mkWUs3PU4+vfNpkXLgqF6ES8rXWS9g5FwRUrgeah//Z3modHVKQnGM4DC
hdRBLqsErhXiqrkoEtidaIBSZtDWbL1OUI4MwuEFp+tiiwFwvAQHL37ohja1WZXt2ON5o1sOxU/1
vT2yqebGKGmgb5K9x/NsB2ucfhna6LKgboJHDUozi7FkIrK5kOfKf0r1GgRERPHDOSF7/6pmgOpy
RYoURBRgZgkPPqtZ+AyLkA7imoGAfqicwhoVa7FfFr3mrP3SxbRzJipZ3694940iPyIVuO6jGNyy
yoVvV+1HaBETVT1j5zPBH3s8OUofngkN/Ly1o8gwMC3YebwNaDr8fOjRrbAtAd5PJiTPQXvzgAFc
a7rSSPfzmkuu7OXrX//Aptmc/PUi/5WPmKu4T/OuyLT9BemBW+r8wQOUKyeXgRblob4RyOvTrYTK
e1m24hLEFjoAHVrO4knqycrEW5yNIzO4CTBjr3z2ao+6IuR1AlXe79NmrzbNRZKKABefbDpxxr+M
M4SS7lueeEAC2B3X++C+Kb0oLsRMZrF30nR5ATfkHpRDkCbvNZxwWvS0FWg//hTdAxGjEnGk+62l
AbGY2d1YMYJrDgP/pfBvqifnlkVMSyWWTRhawpsnxSJMmTNOeRveOrTK0rim7UVSV5+981hN1pet
yAcbLaBytyCgR3nflUjERSrfchP7YuWYHabxNbfVvaXhRYSl6l/LmqkVzGrP7Iz085hy9/WLavti
yOadr5laoXFG4qcEWRP+I0WGN/Q2378EtAZEWZx+NuvTf25Cjix6nvO0Kh+p0BqgXINhQzJscJ2l
bU2fkuAVkoML1qw/8hphG+JeySHQhKt3DEtn39iK3itcmSjPqAH25a2ZGVJzzNa2gBfkP+vzRj6f
HUAZMW83u+29dAARUxldAQhNChn6bzvUESDfBwkuYZ92GnjH9ohIFAgVurqJrOqZVi1+v91H43TP
swaoLMp6vPN2dfAQruoN191yZmVBFGCH1yQ4id6etQjn95S2G4PwHh+Or9lL6dbRYAt4+a8TZus4
S68Yc02EhfrhVAfHFRUP5bJlczLHfT7SnTJTK/cNHJ9iBI4K/fioOZOStfng1B0wcRoUxzC92t/3
Hlj9vVPBX/k93SvIFNwYVL1vzMBxs3CS0WRwzSFyPfMNAAXl6IFXouD65lVMOAN4+PerbragoPmw
Lvo5MQdqV521siiW7n6dpflp
`protect end_protected
