localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTX_CHK = {
  {32'h411dee52, 32'hc0138702} /* (31, 31, 31) {real, imag} */,
  {32'hc08daf0d, 32'h40b2027c} /* (31, 31, 30) {real, imag} */,
  {32'h3eb62f1c, 32'hbf93848f} /* (31, 31, 29) {real, imag} */,
  {32'h3f919b1d, 32'h3f257278} /* (31, 31, 28) {real, imag} */,
  {32'hbf419ccd, 32'h3f1e7756} /* (31, 31, 27) {real, imag} */,
  {32'hbe7abd28, 32'h3dd31204} /* (31, 31, 26) {real, imag} */,
  {32'h3db4c462, 32'hbf2033b4} /* (31, 31, 25) {real, imag} */,
  {32'h3e2eb782, 32'h3f5d0b00} /* (31, 31, 24) {real, imag} */,
  {32'h3e3efc4c, 32'h3eeeb4a8} /* (31, 31, 23) {real, imag} */,
  {32'hbe21aa6b, 32'h3d688044} /* (31, 31, 22) {real, imag} */,
  {32'hbebe7cb9, 32'hbd7c6964} /* (31, 31, 21) {real, imag} */,
  {32'h3e39e30e, 32'hbe54cb9f} /* (31, 31, 20) {real, imag} */,
  {32'h3df54597, 32'hbf120d4f} /* (31, 31, 19) {real, imag} */,
  {32'hbe93965f, 32'h3e9959cb} /* (31, 31, 18) {real, imag} */,
  {32'h3d4e1af4, 32'hbeb59f0a} /* (31, 31, 17) {real, imag} */,
  {32'hbe156dda, 32'hbde8c794} /* (31, 31, 16) {real, imag} */,
  {32'hbdb376be, 32'hbe6bb03b} /* (31, 31, 15) {real, imag} */,
  {32'h3d1663be, 32'hbe3f7cac} /* (31, 31, 14) {real, imag} */,
  {32'hbf0ff067, 32'hbe9a0dd8} /* (31, 31, 13) {real, imag} */,
  {32'h3ee2982f, 32'hbf04c0fc} /* (31, 31, 12) {real, imag} */,
  {32'hbe347e5f, 32'hbe540cf9} /* (31, 31, 11) {real, imag} */,
  {32'h3db0aed2, 32'h3d5ba0ce} /* (31, 31, 10) {real, imag} */,
  {32'hbf0af551, 32'h3d1eae88} /* (31, 31, 9) {real, imag} */,
  {32'hbf006408, 32'h3e4e4434} /* (31, 31, 8) {real, imag} */,
  {32'h3e1b413c, 32'h3ee214f5} /* (31, 31, 7) {real, imag} */,
  {32'hbd3810a0, 32'hbd7fde38} /* (31, 31, 6) {real, imag} */,
  {32'hbf580064, 32'hbdda9e8c} /* (31, 31, 5) {real, imag} */,
  {32'h3f9a1c02, 32'h3e8caad7} /* (31, 31, 4) {real, imag} */,
  {32'hbe9bf57e, 32'hbea5fb3a} /* (31, 31, 3) {real, imag} */,
  {32'hc06f09e9, 32'hbe982aed} /* (31, 31, 2) {real, imag} */,
  {32'h410493cc, 32'h40380d32} /* (31, 31, 1) {real, imag} */,
  {32'h40a6c852, 32'hc03b7234} /* (31, 31, 0) {real, imag} */,
  {32'hc0c99a5c, 32'hc03d7840} /* (31, 30, 31) {real, imag} */,
  {32'h405d3696, 32'hbe5124e8} /* (31, 30, 30) {real, imag} */,
  {32'hbf20ac18, 32'h3f80c31b} /* (31, 30, 29) {real, imag} */,
  {32'hbf36511c, 32'hbea337df} /* (31, 30, 28) {real, imag} */,
  {32'h3ed30186, 32'hbdf37260} /* (31, 30, 27) {real, imag} */,
  {32'h3e097e56, 32'hbeaed806} /* (31, 30, 26) {real, imag} */,
  {32'hbeabb2f7, 32'h3ecb5111} /* (31, 30, 25) {real, imag} */,
  {32'h3f6f2bee, 32'hbe52222c} /* (31, 30, 24) {real, imag} */,
  {32'hbe98dfc2, 32'hbeb158fd} /* (31, 30, 23) {real, imag} */,
  {32'hbd59caf4, 32'hbb1b3b10} /* (31, 30, 22) {real, imag} */,
  {32'hbd34c15e, 32'hbe69df0e} /* (31, 30, 21) {real, imag} */,
  {32'h3e5c355c, 32'hbe4dd14b} /* (31, 30, 20) {real, imag} */,
  {32'h3dc09b1c, 32'h3d4f5d8a} /* (31, 30, 19) {real, imag} */,
  {32'h3e895751, 32'hbec8427a} /* (31, 30, 18) {real, imag} */,
  {32'hbe86fac4, 32'h3d9b8682} /* (31, 30, 17) {real, imag} */,
  {32'hbc631124, 32'h3ccd4240} /* (31, 30, 16) {real, imag} */,
  {32'h3e89e9f6, 32'h3d44be64} /* (31, 30, 15) {real, imag} */,
  {32'hbdeba101, 32'h3d66c780} /* (31, 30, 14) {real, imag} */,
  {32'h3ee2f04c, 32'hbe019754} /* (31, 30, 13) {real, imag} */,
  {32'hbd23ec68, 32'hbd2e130e} /* (31, 30, 12) {real, imag} */,
  {32'h3ee2f668, 32'h3e61515c} /* (31, 30, 11) {real, imag} */,
  {32'hbef2f0ec, 32'h3c8e8310} /* (31, 30, 10) {real, imag} */,
  {32'h3eab479c, 32'hbd8c3dfa} /* (31, 30, 9) {real, imag} */,
  {32'h3f1b96c1, 32'h3e7b7fe6} /* (31, 30, 8) {real, imag} */,
  {32'hbe0a9e1e, 32'h3e1fd663} /* (31, 30, 7) {real, imag} */,
  {32'h3e6a6cf8, 32'hbe838de6} /* (31, 30, 6) {real, imag} */,
  {32'h3f6d2bd4, 32'hbd0c53b0} /* (31, 30, 5) {real, imag} */,
  {32'hbfbfda9e, 32'hbfcd1a50} /* (31, 30, 4) {real, imag} */,
  {32'h3d2cdf70, 32'hbe2eaf80} /* (31, 30, 3) {real, imag} */,
  {32'h40819d18, 32'h40149812} /* (31, 30, 2) {real, imag} */,
  {32'hc0ef6960, 32'h3fc168f2} /* (31, 30, 1) {real, imag} */,
  {32'hc0a76984, 32'h3f2d4ce4} /* (31, 30, 0) {real, imag} */,
  {32'h3f9bedbb, 32'h3cae9a40} /* (31, 29, 31) {real, imag} */,
  {32'hbf3bf5ae, 32'h3f343a34} /* (31, 29, 30) {real, imag} */,
  {32'h3f3d52ca, 32'h3eb569dc} /* (31, 29, 29) {real, imag} */,
  {32'hbe4f0708, 32'hbe4fc6d6} /* (31, 29, 28) {real, imag} */,
  {32'hbf4fc8b4, 32'hbefdcb73} /* (31, 29, 27) {real, imag} */,
  {32'hbe0a434c, 32'hbe34a165} /* (31, 29, 26) {real, imag} */,
  {32'hbe9072bd, 32'hbe03d25f} /* (31, 29, 25) {real, imag} */,
  {32'h3e93b4ba, 32'h3ec30222} /* (31, 29, 24) {real, imag} */,
  {32'hbdd561a2, 32'hbe477273} /* (31, 29, 23) {real, imag} */,
  {32'hbebe0bff, 32'h3e7308ea} /* (31, 29, 22) {real, imag} */,
  {32'h3df7c029, 32'h3e9e2e57} /* (31, 29, 21) {real, imag} */,
  {32'hbe9260de, 32'h3df6e638} /* (31, 29, 20) {real, imag} */,
  {32'hbe667c76, 32'h3e49adce} /* (31, 29, 19) {real, imag} */,
  {32'h3e8b7d17, 32'hbeb81d17} /* (31, 29, 18) {real, imag} */,
  {32'hbd7bca76, 32'h3daced04} /* (31, 29, 17) {real, imag} */,
  {32'hbdbd577a, 32'hbe031819} /* (31, 29, 16) {real, imag} */,
  {32'h3e239150, 32'h3de1ab12} /* (31, 29, 15) {real, imag} */,
  {32'h3efcc18b, 32'h3ed345b8} /* (31, 29, 14) {real, imag} */,
  {32'h3d7eee6c, 32'h3d1dff84} /* (31, 29, 13) {real, imag} */,
  {32'hbda9770b, 32'hbd6b5224} /* (31, 29, 12) {real, imag} */,
  {32'h3c10a1b8, 32'h3f0a7893} /* (31, 29, 11) {real, imag} */,
  {32'h3ddce6d2, 32'hbe4b54ff} /* (31, 29, 10) {real, imag} */,
  {32'hbe81ca50, 32'hbd797fac} /* (31, 29, 9) {real, imag} */,
  {32'h3dd299b0, 32'hbe56086c} /* (31, 29, 8) {real, imag} */,
  {32'h3df30f8c, 32'h3d2cd130} /* (31, 29, 7) {real, imag} */,
  {32'hbd828ff6, 32'h3e01c2d8} /* (31, 29, 6) {real, imag} */,
  {32'hbe2dcfd6, 32'h3e9d4a9e} /* (31, 29, 5) {real, imag} */,
  {32'h3e4e45fe, 32'hbf07ec76} /* (31, 29, 4) {real, imag} */,
  {32'h3f68cefa, 32'hbd0fbcf8} /* (31, 29, 3) {real, imag} */,
  {32'h3f33963e, 32'h3f8d7a5d} /* (31, 29, 2) {real, imag} */,
  {32'hbfb608b6, 32'hbf772bdf} /* (31, 29, 1) {real, imag} */,
  {32'h3e0c0d34, 32'hbf25b2a1} /* (31, 29, 0) {real, imag} */,
  {32'h400b97f5, 32'hbfdb3f8b} /* (31, 28, 31) {real, imag} */,
  {32'hbf9d270a, 32'h3f8f271f} /* (31, 28, 30) {real, imag} */,
  {32'h3e44b08c, 32'hbf00d07c} /* (31, 28, 29) {real, imag} */,
  {32'hbc6ed220, 32'hbf4e1884} /* (31, 28, 28) {real, imag} */,
  {32'h3ec9c876, 32'h3f3f98cf} /* (31, 28, 27) {real, imag} */,
  {32'hbd5b1d20, 32'hbe85cabc} /* (31, 28, 26) {real, imag} */,
  {32'h3ebc07ec, 32'hbeb46270} /* (31, 28, 25) {real, imag} */,
  {32'hbe8fa1f5, 32'hbddddcf8} /* (31, 28, 24) {real, imag} */,
  {32'hbdfd92de, 32'hbe72a6ac} /* (31, 28, 23) {real, imag} */,
  {32'hbec83aa2, 32'hbe082314} /* (31, 28, 22) {real, imag} */,
  {32'h3ea55d38, 32'h3dfb0a90} /* (31, 28, 21) {real, imag} */,
  {32'h3e64a678, 32'h3ec49646} /* (31, 28, 20) {real, imag} */,
  {32'h3eedec7a, 32'h3d99efa9} /* (31, 28, 19) {real, imag} */,
  {32'h3e34afc2, 32'hbdc3539c} /* (31, 28, 18) {real, imag} */,
  {32'hbdac984a, 32'h3e209fa2} /* (31, 28, 17) {real, imag} */,
  {32'h3c0a9b1c, 32'h3ddee748} /* (31, 28, 16) {real, imag} */,
  {32'h3de45e95, 32'hbed0588b} /* (31, 28, 15) {real, imag} */,
  {32'h3e0576ca, 32'h3e15ebf1} /* (31, 28, 14) {real, imag} */,
  {32'h3e4b28c2, 32'h3c8655f8} /* (31, 28, 13) {real, imag} */,
  {32'h3f1eb55e, 32'h3eb29cf9} /* (31, 28, 12) {real, imag} */,
  {32'hbeae4620, 32'hbe40408f} /* (31, 28, 11) {real, imag} */,
  {32'h3e7950e0, 32'hbee09340} /* (31, 28, 10) {real, imag} */,
  {32'hbe8443ac, 32'hbd53453e} /* (31, 28, 9) {real, imag} */,
  {32'hbd8fe500, 32'h3e456b6c} /* (31, 28, 8) {real, imag} */,
  {32'hbe87ea4e, 32'hbd626a54} /* (31, 28, 7) {real, imag} */,
  {32'hbea1d585, 32'h3e7b82a8} /* (31, 28, 6) {real, imag} */,
  {32'hbf0bfcda, 32'h3f051f03} /* (31, 28, 5) {real, imag} */,
  {32'h3f6042af, 32'hbe7156a7} /* (31, 28, 4) {real, imag} */,
  {32'hbe8fbb80, 32'hbb366200} /* (31, 28, 3) {real, imag} */,
  {32'hc00cd4ce, 32'h3e024a68} /* (31, 28, 2) {real, imag} */,
  {32'h3f1c4ad8, 32'hbfb11866} /* (31, 28, 1) {real, imag} */,
  {32'h3ff929bb, 32'hbef78e14} /* (31, 28, 0) {real, imag} */,
  {32'hbf9ae460, 32'h3f8d72c8} /* (31, 27, 31) {real, imag} */,
  {32'h3f9e150c, 32'hbf22426c} /* (31, 27, 30) {real, imag} */,
  {32'hbf36e6c7, 32'h3e59bee6} /* (31, 27, 29) {real, imag} */,
  {32'hbf4dd508, 32'h3e33407b} /* (31, 27, 28) {real, imag} */,
  {32'h3d47fd20, 32'hbea3aa34} /* (31, 27, 27) {real, imag} */,
  {32'h3f05fe23, 32'hbe69b1fe} /* (31, 27, 26) {real, imag} */,
  {32'h3ec64126, 32'h3f25b9b8} /* (31, 27, 25) {real, imag} */,
  {32'hbd31666c, 32'hbebe995e} /* (31, 27, 24) {real, imag} */,
  {32'h3d5a6cb6, 32'hbeae0e2d} /* (31, 27, 23) {real, imag} */,
  {32'h3dd06fff, 32'hbe83cb71} /* (31, 27, 22) {real, imag} */,
  {32'hbedaee64, 32'h3e2a447c} /* (31, 27, 21) {real, imag} */,
  {32'h3e1ad9ac, 32'hbe2615b6} /* (31, 27, 20) {real, imag} */,
  {32'hbdf78f8c, 32'hbe107087} /* (31, 27, 19) {real, imag} */,
  {32'hbe714d14, 32'hbe14ddf8} /* (31, 27, 18) {real, imag} */,
  {32'hbdf0d2ba, 32'h3e4fe692} /* (31, 27, 17) {real, imag} */,
  {32'hbebeb538, 32'h3ade6d00} /* (31, 27, 16) {real, imag} */,
  {32'hbdc538e9, 32'h3db481fc} /* (31, 27, 15) {real, imag} */,
  {32'h3cc8afe8, 32'hbe0b4f34} /* (31, 27, 14) {real, imag} */,
  {32'h3e776658, 32'h3d89a787} /* (31, 27, 13) {real, imag} */,
  {32'h3edb75a4, 32'h3eb22510} /* (31, 27, 12) {real, imag} */,
  {32'hbdf44fbb, 32'hbec768a9} /* (31, 27, 11) {real, imag} */,
  {32'h3e489cda, 32'h3e9036b4} /* (31, 27, 10) {real, imag} */,
  {32'h3d9d31ad, 32'hbd635210} /* (31, 27, 9) {real, imag} */,
  {32'hbe050512, 32'h3c2b8fb0} /* (31, 27, 8) {real, imag} */,
  {32'hbe9f7293, 32'hbec6d03c} /* (31, 27, 7) {real, imag} */,
  {32'h3dda5d36, 32'hbddd2658} /* (31, 27, 6) {real, imag} */,
  {32'h3f35ed08, 32'h3da19d04} /* (31, 27, 5) {real, imag} */,
  {32'hbd78d7b2, 32'h3f13d560} /* (31, 27, 4) {real, imag} */,
  {32'hbd8cb030, 32'h3e5ec44c} /* (31, 27, 3) {real, imag} */,
  {32'h3e8b8b90, 32'h3f094173} /* (31, 27, 2) {real, imag} */,
  {32'hbfcaf712, 32'h3dd0c9e2} /* (31, 27, 1) {real, imag} */,
  {32'hbfb893cf, 32'hbe52dc80} /* (31, 27, 0) {real, imag} */,
  {32'hbf0981a3, 32'h3e08c332} /* (31, 26, 31) {real, imag} */,
  {32'hbd742db6, 32'h3f3a80eb} /* (31, 26, 30) {real, imag} */,
  {32'h3e203cb0, 32'hbdb1741e} /* (31, 26, 29) {real, imag} */,
  {32'hbd9133dc, 32'hbe443be0} /* (31, 26, 28) {real, imag} */,
  {32'h3ebe0844, 32'hbeb9b7c6} /* (31, 26, 27) {real, imag} */,
  {32'hbe69ead0, 32'h3cae1798} /* (31, 26, 26) {real, imag} */,
  {32'hbeeb66f3, 32'hbeb550c5} /* (31, 26, 25) {real, imag} */,
  {32'h3edcb0f2, 32'hbe89e8af} /* (31, 26, 24) {real, imag} */,
  {32'h3e094cfb, 32'h3b9c0a00} /* (31, 26, 23) {real, imag} */,
  {32'hbe541c83, 32'h3e81bad7} /* (31, 26, 22) {real, imag} */,
  {32'hbcf641e8, 32'hbb9e9700} /* (31, 26, 21) {real, imag} */,
  {32'hbe992283, 32'hbc83d8ac} /* (31, 26, 20) {real, imag} */,
  {32'hbe88d089, 32'h3ea82d26} /* (31, 26, 19) {real, imag} */,
  {32'h3da81c76, 32'h3ec47cdf} /* (31, 26, 18) {real, imag} */,
  {32'h3e2cefb7, 32'hbe5b3ad6} /* (31, 26, 17) {real, imag} */,
  {32'h3de3b9c0, 32'hbd528bf4} /* (31, 26, 16) {real, imag} */,
  {32'hbe310418, 32'h3ea579d2} /* (31, 26, 15) {real, imag} */,
  {32'h3cabda52, 32'hbe784644} /* (31, 26, 14) {real, imag} */,
  {32'hbeb00fbd, 32'h3cdb33f8} /* (31, 26, 13) {real, imag} */,
  {32'hbeb1d34a, 32'h3c80427a} /* (31, 26, 12) {real, imag} */,
  {32'h3ea2b3a2, 32'h3ec95768} /* (31, 26, 11) {real, imag} */,
  {32'h3d239282, 32'h3ea10a6a} /* (31, 26, 10) {real, imag} */,
  {32'hbe1a798c, 32'h3ee5a3df} /* (31, 26, 9) {real, imag} */,
  {32'h3e2e60dc, 32'hbe595abe} /* (31, 26, 8) {real, imag} */,
  {32'hbd673422, 32'h3df3e94a} /* (31, 26, 7) {real, imag} */,
  {32'h3e73b8d0, 32'hbf05d8c4} /* (31, 26, 6) {real, imag} */,
  {32'hbe240e4c, 32'hbe478610} /* (31, 26, 5) {real, imag} */,
  {32'hbdb79818, 32'hbdd32e6a} /* (31, 26, 4) {real, imag} */,
  {32'h3ed501e8, 32'hbc9024a0} /* (31, 26, 3) {real, imag} */,
  {32'hbef93ef2, 32'h3f12f0bd} /* (31, 26, 2) {real, imag} */,
  {32'hbe9e14ac, 32'hbf190a00} /* (31, 26, 1) {real, imag} */,
  {32'h3f0b9ecc, 32'h3e894da7} /* (31, 26, 0) {real, imag} */,
  {32'hbe7ba278, 32'hbd5f8b58} /* (31, 25, 31) {real, imag} */,
  {32'h3ea93268, 32'h3e965ef5} /* (31, 25, 30) {real, imag} */,
  {32'h3e9f2e3e, 32'hbc3c42c0} /* (31, 25, 29) {real, imag} */,
  {32'h3e1e1d5e, 32'h3ca80c30} /* (31, 25, 28) {real, imag} */,
  {32'h3e89c6b4, 32'h3c2c5f60} /* (31, 25, 27) {real, imag} */,
  {32'h3e41bab5, 32'h3db31082} /* (31, 25, 26) {real, imag} */,
  {32'h3d1a2034, 32'h3d3470e4} /* (31, 25, 25) {real, imag} */,
  {32'hbe378ca5, 32'hbe2c7309} /* (31, 25, 24) {real, imag} */,
  {32'hbe54eccd, 32'h3e90d042} /* (31, 25, 23) {real, imag} */,
  {32'h3e78dbc1, 32'hba941200} /* (31, 25, 22) {real, imag} */,
  {32'h3eb6823c, 32'hbd750374} /* (31, 25, 21) {real, imag} */,
  {32'hbd719626, 32'h3e31cac9} /* (31, 25, 20) {real, imag} */,
  {32'hbe4dd438, 32'h3db2e3e0} /* (31, 25, 19) {real, imag} */,
  {32'hbe739be6, 32'hbe910df6} /* (31, 25, 18) {real, imag} */,
  {32'h3d99860d, 32'hbe30dd6d} /* (31, 25, 17) {real, imag} */,
  {32'h3d85a819, 32'h3db4fd79} /* (31, 25, 16) {real, imag} */,
  {32'h3ee6fd63, 32'hbe38346a} /* (31, 25, 15) {real, imag} */,
  {32'hbe20c473, 32'hbe40fea0} /* (31, 25, 14) {real, imag} */,
  {32'hbd683328, 32'hbe644fbc} /* (31, 25, 13) {real, imag} */,
  {32'hbe8a01ef, 32'h3e1af006} /* (31, 25, 12) {real, imag} */,
  {32'hbd08a6e0, 32'hbea3dc38} /* (31, 25, 11) {real, imag} */,
  {32'hbe0df467, 32'hbc9b1934} /* (31, 25, 10) {real, imag} */,
  {32'h3e9f2d74, 32'hbdcb695e} /* (31, 25, 9) {real, imag} */,
  {32'hbe42e356, 32'hbebc8bcd} /* (31, 25, 8) {real, imag} */,
  {32'h3e479370, 32'h3d6b8a66} /* (31, 25, 7) {real, imag} */,
  {32'h3e8a5bc2, 32'hbe582780} /* (31, 25, 6) {real, imag} */,
  {32'hbe7785e5, 32'h3e4e5842} /* (31, 25, 5) {real, imag} */,
  {32'hbedbaf1b, 32'hbd49e580} /* (31, 25, 4) {real, imag} */,
  {32'h3d67df34, 32'h3cf80128} /* (31, 25, 3) {real, imag} */,
  {32'hbe313a1e, 32'h3e2653c2} /* (31, 25, 2) {real, imag} */,
  {32'h3e67ff8e, 32'hbbda9460} /* (31, 25, 1) {real, imag} */,
  {32'h3f3c68b9, 32'hbeddbf4f} /* (31, 25, 0) {real, imag} */,
  {32'hbf1a969c, 32'h3eedb412} /* (31, 24, 31) {real, imag} */,
  {32'h3ed94f0e, 32'hbf94167c} /* (31, 24, 30) {real, imag} */,
  {32'hbf44b78b, 32'h3d6e5298} /* (31, 24, 29) {real, imag} */,
  {32'h3e42184c, 32'hbe49c841} /* (31, 24, 28) {real, imag} */,
  {32'h3d66175a, 32'hbe6e92c0} /* (31, 24, 27) {real, imag} */,
  {32'h3eaf152f, 32'hbe174dd7} /* (31, 24, 26) {real, imag} */,
  {32'hbd945f40, 32'h3ebbd7cf} /* (31, 24, 25) {real, imag} */,
  {32'h3d570de0, 32'h3e756abe} /* (31, 24, 24) {real, imag} */,
  {32'h3da8504e, 32'h3e078ba2} /* (31, 24, 23) {real, imag} */,
  {32'hbd2b4bc4, 32'hbe915521} /* (31, 24, 22) {real, imag} */,
  {32'hbe549f56, 32'hbe4cf1b2} /* (31, 24, 21) {real, imag} */,
  {32'hbc036b80, 32'hbe915e94} /* (31, 24, 20) {real, imag} */,
  {32'h3e08d7d6, 32'h3d60e870} /* (31, 24, 19) {real, imag} */,
  {32'h3d691e8c, 32'hbd8c5802} /* (31, 24, 18) {real, imag} */,
  {32'hbd0ba3a0, 32'h3d2a554a} /* (31, 24, 17) {real, imag} */,
  {32'hbd452614, 32'h3dd26313} /* (31, 24, 16) {real, imag} */,
  {32'h3e8095c5, 32'hbedd26c9} /* (31, 24, 15) {real, imag} */,
  {32'hbe390fcc, 32'hbe1af45e} /* (31, 24, 14) {real, imag} */,
  {32'hbdb9c6be, 32'hbdb1a2e4} /* (31, 24, 13) {real, imag} */,
  {32'hbd7dd8d0, 32'hbdf5aaaa} /* (31, 24, 12) {real, imag} */,
  {32'hbe64b441, 32'hbd17b2cf} /* (31, 24, 11) {real, imag} */,
  {32'h3e1babf0, 32'h3e5466b6} /* (31, 24, 10) {real, imag} */,
  {32'h3db7007c, 32'hbe8f0ba4} /* (31, 24, 9) {real, imag} */,
  {32'hbe492ac2, 32'h3db77b80} /* (31, 24, 8) {real, imag} */,
  {32'h3e72cd22, 32'h3bceb150} /* (31, 24, 7) {real, imag} */,
  {32'hbedea0ef, 32'h3d17d3d0} /* (31, 24, 6) {real, imag} */,
  {32'h3e1bef4b, 32'hbde0721f} /* (31, 24, 5) {real, imag} */,
  {32'hbedf86e0, 32'hbe9cb912} /* (31, 24, 4) {real, imag} */,
  {32'hbe6482e0, 32'hbcece152} /* (31, 24, 3) {real, imag} */,
  {32'h3f884781, 32'h3df5c13c} /* (31, 24, 2) {real, imag} */,
  {32'hbf50e843, 32'h3f24fb94} /* (31, 24, 1) {real, imag} */,
  {32'hbf114c26, 32'hba421600} /* (31, 24, 0) {real, imag} */,
  {32'h3e4c622c, 32'h3d185c98} /* (31, 23, 31) {real, imag} */,
  {32'hbdff7808, 32'h3f04fa9e} /* (31, 23, 30) {real, imag} */,
  {32'hbf521346, 32'hbe096349} /* (31, 23, 29) {real, imag} */,
  {32'h3f18b11b, 32'h3cce8150} /* (31, 23, 28) {real, imag} */,
  {32'hbdf3cc42, 32'h3b8c8420} /* (31, 23, 27) {real, imag} */,
  {32'hbea282da, 32'h3dfe8882} /* (31, 23, 26) {real, imag} */,
  {32'h3ef12da5, 32'h3e48d34e} /* (31, 23, 25) {real, imag} */,
  {32'hbe70dc44, 32'h3ebd8d9c} /* (31, 23, 24) {real, imag} */,
  {32'h3de8b5d8, 32'h3eb5b0c7} /* (31, 23, 23) {real, imag} */,
  {32'h3dcac83a, 32'hbd9e7aaa} /* (31, 23, 22) {real, imag} */,
  {32'h3e0f7852, 32'h3ca32ec4} /* (31, 23, 21) {real, imag} */,
  {32'hbd7bc24e, 32'h3ec22173} /* (31, 23, 20) {real, imag} */,
  {32'h3f05fe52, 32'h3bb170a0} /* (31, 23, 19) {real, imag} */,
  {32'h3e663a16, 32'h3d42c578} /* (31, 23, 18) {real, imag} */,
  {32'h3d6fa734, 32'h3db7f21d} /* (31, 23, 17) {real, imag} */,
  {32'h3d6b3254, 32'h3d606e7c} /* (31, 23, 16) {real, imag} */,
  {32'h3e994d99, 32'h3dbecb92} /* (31, 23, 15) {real, imag} */,
  {32'hbe472524, 32'h3d368b96} /* (31, 23, 14) {real, imag} */,
  {32'hbec8ab2c, 32'h3e148950} /* (31, 23, 13) {real, imag} */,
  {32'h3d2d2ad0, 32'h3e0c6ea8} /* (31, 23, 12) {real, imag} */,
  {32'h3e64eb5c, 32'h3e6de0ce} /* (31, 23, 11) {real, imag} */,
  {32'h3b21e380, 32'hbe128605} /* (31, 23, 10) {real, imag} */,
  {32'hbd974a9c, 32'hbd3cfafe} /* (31, 23, 9) {real, imag} */,
  {32'h3d8aae08, 32'h3d6de7f4} /* (31, 23, 8) {real, imag} */,
  {32'h3daeeba3, 32'hbaa42480} /* (31, 23, 7) {real, imag} */,
  {32'h3e08c8e4, 32'hbe67a1cc} /* (31, 23, 6) {real, imag} */,
  {32'h3e75c4d8, 32'h3e7e20d1} /* (31, 23, 5) {real, imag} */,
  {32'h3f0b52f8, 32'hbe8fa040} /* (31, 23, 4) {real, imag} */,
  {32'h3ed3cc2b, 32'hbda51eb4} /* (31, 23, 3) {real, imag} */,
  {32'h3dbbd282, 32'hbe75aaae} /* (31, 23, 2) {real, imag} */,
  {32'hbd151e64, 32'hbf306eab} /* (31, 23, 1) {real, imag} */,
  {32'h3c6423a0, 32'hbea98906} /* (31, 23, 0) {real, imag} */,
  {32'h3efb2137, 32'h3de2948a} /* (31, 22, 31) {real, imag} */,
  {32'h3ca92820, 32'h3e899ad6} /* (31, 22, 30) {real, imag} */,
  {32'h3eefcaff, 32'h3e1234fb} /* (31, 22, 29) {real, imag} */,
  {32'hbd021650, 32'hbe504090} /* (31, 22, 28) {real, imag} */,
  {32'h3c417f20, 32'h3e2459bc} /* (31, 22, 27) {real, imag} */,
  {32'hbe32ae8a, 32'h3ea80efc} /* (31, 22, 26) {real, imag} */,
  {32'h3e8499a7, 32'hbe9ac8ae} /* (31, 22, 25) {real, imag} */,
  {32'hbdcb8329, 32'h3e1ed2ac} /* (31, 22, 24) {real, imag} */,
  {32'h3e499dcc, 32'hbea66e8c} /* (31, 22, 23) {real, imag} */,
  {32'hbe9be0ba, 32'h3ca67df0} /* (31, 22, 22) {real, imag} */,
  {32'hbe20c3c1, 32'h3e04d479} /* (31, 22, 21) {real, imag} */,
  {32'hbe5003ac, 32'hbec2e57a} /* (31, 22, 20) {real, imag} */,
  {32'h3c9332f0, 32'hbed26b2c} /* (31, 22, 19) {real, imag} */,
  {32'hbd3eac1c, 32'h3c958a18} /* (31, 22, 18) {real, imag} */,
  {32'hbc8d18d3, 32'h3c95a1f8} /* (31, 22, 17) {real, imag} */,
  {32'hbdc78fae, 32'hbdbb0c29} /* (31, 22, 16) {real, imag} */,
  {32'hbe383a84, 32'h3dabd4e2} /* (31, 22, 15) {real, imag} */,
  {32'h3e49545a, 32'h3e7fc24c} /* (31, 22, 14) {real, imag} */,
  {32'h3d729148, 32'h3eb5247e} /* (31, 22, 13) {real, imag} */,
  {32'hbe4dc24c, 32'hbee1f6d6} /* (31, 22, 12) {real, imag} */,
  {32'hbed91886, 32'h3e357960} /* (31, 22, 11) {real, imag} */,
  {32'h3eb605f8, 32'h3da8a82e} /* (31, 22, 10) {real, imag} */,
  {32'hbf0732e3, 32'hbe92e901} /* (31, 22, 9) {real, imag} */,
  {32'hbdd65b06, 32'h3d305448} /* (31, 22, 8) {real, imag} */,
  {32'hbdbf5fa4, 32'h3e6bcc2c} /* (31, 22, 7) {real, imag} */,
  {32'hbd6d302c, 32'hbe873d2c} /* (31, 22, 6) {real, imag} */,
  {32'hbdcce049, 32'h3ed29c58} /* (31, 22, 5) {real, imag} */,
  {32'h3efaab8a, 32'h3ddd56f4} /* (31, 22, 4) {real, imag} */,
  {32'hbc95a9f0, 32'hbdf6f8b6} /* (31, 22, 3) {real, imag} */,
  {32'h3d485468, 32'hbdc09008} /* (31, 22, 2) {real, imag} */,
  {32'hbdb7182e, 32'hbed5751c} /* (31, 22, 1) {real, imag} */,
  {32'hbe9b69de, 32'hbd716ea6} /* (31, 22, 0) {real, imag} */,
  {32'hbda1a8e4, 32'hbdca40bc} /* (31, 21, 31) {real, imag} */,
  {32'hbe433bf4, 32'hbdeb53c8} /* (31, 21, 30) {real, imag} */,
  {32'h3e08b553, 32'h3d42f370} /* (31, 21, 29) {real, imag} */,
  {32'h3e25fa2a, 32'hbed776c7} /* (31, 21, 28) {real, imag} */,
  {32'h3e87d1fd, 32'h3e7b2ea3} /* (31, 21, 27) {real, imag} */,
  {32'h3d6bae20, 32'hbe1bf936} /* (31, 21, 26) {real, imag} */,
  {32'hbe631f3a, 32'h3e93480f} /* (31, 21, 25) {real, imag} */,
  {32'h3e41b487, 32'h3cadbd94} /* (31, 21, 24) {real, imag} */,
  {32'hbdac9ad2, 32'h3d7942dc} /* (31, 21, 23) {real, imag} */,
  {32'h3f1546ee, 32'hbe7efc90} /* (31, 21, 22) {real, imag} */,
  {32'h3e31c0c8, 32'hbefdb588} /* (31, 21, 21) {real, imag} */,
  {32'hbe68ec32, 32'h3f4ddde0} /* (31, 21, 20) {real, imag} */,
  {32'hbea4ae6e, 32'h3e43f882} /* (31, 21, 19) {real, imag} */,
  {32'hbec6cd51, 32'h3d02daf4} /* (31, 21, 18) {real, imag} */,
  {32'h3c9997e4, 32'h3d8a0578} /* (31, 21, 17) {real, imag} */,
  {32'h3cfb1668, 32'hbd05a969} /* (31, 21, 16) {real, imag} */,
  {32'h3d66146c, 32'hbdd5fabb} /* (31, 21, 15) {real, imag} */,
  {32'hbc40bd30, 32'h3e86079f} /* (31, 21, 14) {real, imag} */,
  {32'hbdfdc950, 32'h3ef6c5f8} /* (31, 21, 13) {real, imag} */,
  {32'hbe3e6374, 32'hbe5bb608} /* (31, 21, 12) {real, imag} */,
  {32'h3e92f17d, 32'hbee39db0} /* (31, 21, 11) {real, imag} */,
  {32'hbc509060, 32'h3cfaff60} /* (31, 21, 10) {real, imag} */,
  {32'h3d4f8258, 32'hbf02107c} /* (31, 21, 9) {real, imag} */,
  {32'h3e0376c0, 32'h3e80dec2} /* (31, 21, 8) {real, imag} */,
  {32'hbf014fd7, 32'hbe088f4e} /* (31, 21, 7) {real, imag} */,
  {32'hbdc356a4, 32'h3e023a46} /* (31, 21, 6) {real, imag} */,
  {32'hbce0ec54, 32'hbbfca8c0} /* (31, 21, 5) {real, imag} */,
  {32'hbe85a598, 32'hbe954e42} /* (31, 21, 4) {real, imag} */,
  {32'h3da0c944, 32'hbe2d8e7a} /* (31, 21, 3) {real, imag} */,
  {32'hbde53658, 32'hbec37cfc} /* (31, 21, 2) {real, imag} */,
  {32'h3da8efb0, 32'h3e4c6be4} /* (31, 21, 1) {real, imag} */,
  {32'h3d8acf98, 32'h3e302c98} /* (31, 21, 0) {real, imag} */,
  {32'hbdd43cf8, 32'hbebf0ac8} /* (31, 20, 31) {real, imag} */,
  {32'hbed89a43, 32'h3d24cdc4} /* (31, 20, 30) {real, imag} */,
  {32'hbe564c01, 32'hbc06f570} /* (31, 20, 29) {real, imag} */,
  {32'h3d580b50, 32'h3e04a77d} /* (31, 20, 28) {real, imag} */,
  {32'h3c69c1c0, 32'h3d809b30} /* (31, 20, 27) {real, imag} */,
  {32'h3c358d80, 32'h3e3a8861} /* (31, 20, 26) {real, imag} */,
  {32'hbe88fbc3, 32'h3ea4c18d} /* (31, 20, 25) {real, imag} */,
  {32'h3dff55dc, 32'hbe9a0719} /* (31, 20, 24) {real, imag} */,
  {32'hbb0d6120, 32'h3ee156ec} /* (31, 20, 23) {real, imag} */,
  {32'h3e3589ae, 32'hbe956562} /* (31, 20, 22) {real, imag} */,
  {32'h3e4ceeb6, 32'h3e1d76f5} /* (31, 20, 21) {real, imag} */,
  {32'hbe24d572, 32'hbe1b5ac0} /* (31, 20, 20) {real, imag} */,
  {32'hbef8413e, 32'hbe1d2f8d} /* (31, 20, 19) {real, imag} */,
  {32'h3da7b070, 32'hbe8028b7} /* (31, 20, 18) {real, imag} */,
  {32'hbe792e4c, 32'hbe15de98} /* (31, 20, 17) {real, imag} */,
  {32'h3e0742f1, 32'h3db11834} /* (31, 20, 16) {real, imag} */,
  {32'h3e3de3ee, 32'h3e168084} /* (31, 20, 15) {real, imag} */,
  {32'hbeede012, 32'h3c974a9c} /* (31, 20, 14) {real, imag} */,
  {32'hbf050658, 32'h3df63ff8} /* (31, 20, 13) {real, imag} */,
  {32'hbe645933, 32'hbea1384f} /* (31, 20, 12) {real, imag} */,
  {32'h3e98e874, 32'hbe89367a} /* (31, 20, 11) {real, imag} */,
  {32'hbd03b0a0, 32'hbe878050} /* (31, 20, 10) {real, imag} */,
  {32'h3d4cdd22, 32'h3d1f3a48} /* (31, 20, 9) {real, imag} */,
  {32'hbe50279e, 32'h3eb709e2} /* (31, 20, 8) {real, imag} */,
  {32'h3c95e1c8, 32'hbee82ee6} /* (31, 20, 7) {real, imag} */,
  {32'hbc094928, 32'h3e16d987} /* (31, 20, 6) {real, imag} */,
  {32'h3e1d1826, 32'h3e5b0090} /* (31, 20, 5) {real, imag} */,
  {32'hbe8a7620, 32'h3ef3d52d} /* (31, 20, 4) {real, imag} */,
  {32'h3e2ad024, 32'h3d6399a8} /* (31, 20, 3) {real, imag} */,
  {32'h3e9c4160, 32'hbe8a4e9d} /* (31, 20, 2) {real, imag} */,
  {32'h3d80ec8a, 32'h3e21efa1} /* (31, 20, 1) {real, imag} */,
  {32'h3dec86e8, 32'hbd5ee5a0} /* (31, 20, 0) {real, imag} */,
  {32'h3e581b6a, 32'h3d31fd74} /* (31, 19, 31) {real, imag} */,
  {32'h3d2b63d0, 32'h3ce2140e} /* (31, 19, 30) {real, imag} */,
  {32'hbdc64b7b, 32'hbe2b7c00} /* (31, 19, 29) {real, imag} */,
  {32'hbe6f1cd4, 32'hbc49b078} /* (31, 19, 28) {real, imag} */,
  {32'hbe9c26dd, 32'h3d24c24c} /* (31, 19, 27) {real, imag} */,
  {32'hbdb47838, 32'hbd2bb318} /* (31, 19, 26) {real, imag} */,
  {32'h3e97f0f1, 32'h3c992d38} /* (31, 19, 25) {real, imag} */,
  {32'hbebc521a, 32'h3d7faf34} /* (31, 19, 24) {real, imag} */,
  {32'h3ea51077, 32'h3e23cb33} /* (31, 19, 23) {real, imag} */,
  {32'h3d1e061c, 32'hbd97175f} /* (31, 19, 22) {real, imag} */,
  {32'hbe9ccd3e, 32'hbe1bca84} /* (31, 19, 21) {real, imag} */,
  {32'hbe03d163, 32'hbc01be44} /* (31, 19, 20) {real, imag} */,
  {32'hbec929d3, 32'h3dc2d611} /* (31, 19, 19) {real, imag} */,
  {32'h3e260478, 32'hbc04a4ac} /* (31, 19, 18) {real, imag} */,
  {32'hbe2d712a, 32'h3c8bea74} /* (31, 19, 17) {real, imag} */,
  {32'hbd2e0778, 32'hbea66b70} /* (31, 19, 16) {real, imag} */,
  {32'h3e166334, 32'h3e827db3} /* (31, 19, 15) {real, imag} */,
  {32'h3f171075, 32'h3e4809a3} /* (31, 19, 14) {real, imag} */,
  {32'h3ee9b856, 32'hbe557d13} /* (31, 19, 13) {real, imag} */,
  {32'h3e12d966, 32'h3cb3c830} /* (31, 19, 12) {real, imag} */,
  {32'hbd8bea62, 32'h3e9ebb67} /* (31, 19, 11) {real, imag} */,
  {32'hbb682a60, 32'h3df0add0} /* (31, 19, 10) {real, imag} */,
  {32'h3dae39ce, 32'h3d9df376} /* (31, 19, 9) {real, imag} */,
  {32'hbde4bd6c, 32'h3e6d93fc} /* (31, 19, 8) {real, imag} */,
  {32'hbc7d8678, 32'h3d637ce8} /* (31, 19, 7) {real, imag} */,
  {32'h3e1b2502, 32'h3ea7c662} /* (31, 19, 6) {real, imag} */,
  {32'h3ce8bb7a, 32'h3e9442a4} /* (31, 19, 5) {real, imag} */,
  {32'h3b2664c0, 32'hbda0a082} /* (31, 19, 4) {real, imag} */,
  {32'h3e9e1c76, 32'h3b8577a8} /* (31, 19, 3) {real, imag} */,
  {32'hbee6f562, 32'hbdcfa33c} /* (31, 19, 2) {real, imag} */,
  {32'hbe580b49, 32'h3e24a311} /* (31, 19, 1) {real, imag} */,
  {32'hbe7e0ebe, 32'h3d1b3684} /* (31, 19, 0) {real, imag} */,
  {32'h3e81bf84, 32'h3e0b7d9b} /* (31, 18, 31) {real, imag} */,
  {32'h3e293009, 32'hbd7e9298} /* (31, 18, 30) {real, imag} */,
  {32'h3e83903f, 32'hbe2cb238} /* (31, 18, 29) {real, imag} */,
  {32'h3d4a79ae, 32'h3e6f80ca} /* (31, 18, 28) {real, imag} */,
  {32'h3eab6264, 32'hbe97f7ec} /* (31, 18, 27) {real, imag} */,
  {32'hbebb58ff, 32'hbd4cc574} /* (31, 18, 26) {real, imag} */,
  {32'hbeb3f133, 32'hbf3296e0} /* (31, 18, 25) {real, imag} */,
  {32'h3e3b7a3a, 32'h3c817220} /* (31, 18, 24) {real, imag} */,
  {32'h3eaf36b2, 32'hbde82970} /* (31, 18, 23) {real, imag} */,
  {32'h3e9751a8, 32'hbdb1307c} /* (31, 18, 22) {real, imag} */,
  {32'hbe1bceac, 32'h3d63da30} /* (31, 18, 21) {real, imag} */,
  {32'h3b31bcc0, 32'hbda7ea2e} /* (31, 18, 20) {real, imag} */,
  {32'h3dd01aa2, 32'hbee3deb6} /* (31, 18, 19) {real, imag} */,
  {32'h3c7086c0, 32'h3eceb670} /* (31, 18, 18) {real, imag} */,
  {32'hbe17802f, 32'h3d47bf90} /* (31, 18, 17) {real, imag} */,
  {32'hbda0b9a0, 32'hbe84032c} /* (31, 18, 16) {real, imag} */,
  {32'hbe37c90e, 32'h3d8fe72c} /* (31, 18, 15) {real, imag} */,
  {32'hbe125510, 32'hbb3a12a0} /* (31, 18, 14) {real, imag} */,
  {32'hbdcca990, 32'hbef35c1c} /* (31, 18, 13) {real, imag} */,
  {32'hbe91509c, 32'hbd88059a} /* (31, 18, 12) {real, imag} */,
  {32'h3d1be65a, 32'h3e23716b} /* (31, 18, 11) {real, imag} */,
  {32'h3eba0946, 32'hbef8b440} /* (31, 18, 10) {real, imag} */,
  {32'hbe874454, 32'hbdc751d2} /* (31, 18, 9) {real, imag} */,
  {32'h3d9acde2, 32'h3e727ffb} /* (31, 18, 8) {real, imag} */,
  {32'h3dde656c, 32'hbe060b01} /* (31, 18, 7) {real, imag} */,
  {32'h3eee40ac, 32'hbe32cdec} /* (31, 18, 6) {real, imag} */,
  {32'hbee1b329, 32'hbe417294} /* (31, 18, 5) {real, imag} */,
  {32'hbeb65b50, 32'h3d99b62d} /* (31, 18, 4) {real, imag} */,
  {32'hbe2c0c12, 32'h3da76470} /* (31, 18, 3) {real, imag} */,
  {32'h3e3c42c3, 32'hbe3b78df} /* (31, 18, 2) {real, imag} */,
  {32'hbe735f1a, 32'h3da968e9} /* (31, 18, 1) {real, imag} */,
  {32'hbdcce2f7, 32'h3df42a7a} /* (31, 18, 0) {real, imag} */,
  {32'h3df4a53b, 32'hbe04cc7a} /* (31, 17, 31) {real, imag} */,
  {32'hbbdbfb60, 32'h3dfef370} /* (31, 17, 30) {real, imag} */,
  {32'h3d014068, 32'hbda5de1e} /* (31, 17, 29) {real, imag} */,
  {32'h3cd3b3e0, 32'hbdee7580} /* (31, 17, 28) {real, imag} */,
  {32'h3d9487ef, 32'hbd43c96c} /* (31, 17, 27) {real, imag} */,
  {32'h3e2e9c56, 32'hbdaf9e12} /* (31, 17, 26) {real, imag} */,
  {32'h3e29fbe4, 32'h3e922d20} /* (31, 17, 25) {real, imag} */,
  {32'hbe6f167a, 32'hbc7a0940} /* (31, 17, 24) {real, imag} */,
  {32'h3e220942, 32'hbddf8dbe} /* (31, 17, 23) {real, imag} */,
  {32'hbe0b75ea, 32'h3d1200e4} /* (31, 17, 22) {real, imag} */,
  {32'h3e85b139, 32'h3da74b7c} /* (31, 17, 21) {real, imag} */,
  {32'h3deae666, 32'hbe95cad1} /* (31, 17, 20) {real, imag} */,
  {32'hbe0f8b84, 32'h3e181a4e} /* (31, 17, 19) {real, imag} */,
  {32'h3d80daef, 32'hbec26d7a} /* (31, 17, 18) {real, imag} */,
  {32'hbcb18148, 32'h3df88808} /* (31, 17, 17) {real, imag} */,
  {32'h3c8a84ac, 32'hbd6cb748} /* (31, 17, 16) {real, imag} */,
  {32'h3dc5f59a, 32'h3e78547c} /* (31, 17, 15) {real, imag} */,
  {32'hbe1f0069, 32'hbe83ae12} /* (31, 17, 14) {real, imag} */,
  {32'h3b4e6b00, 32'h3e0753f7} /* (31, 17, 13) {real, imag} */,
  {32'h3d523c7f, 32'hbe8f67df} /* (31, 17, 12) {real, imag} */,
  {32'h3e4bbabb, 32'h3e3b11bf} /* (31, 17, 11) {real, imag} */,
  {32'h3d5d7938, 32'hbe5890eb} /* (31, 17, 10) {real, imag} */,
  {32'h3ddad27c, 32'h3e6f4fdd} /* (31, 17, 9) {real, imag} */,
  {32'hbd5bea20, 32'hbd30d2f8} /* (31, 17, 8) {real, imag} */,
  {32'hbe25a7ee, 32'h3e0fa31e} /* (31, 17, 7) {real, imag} */,
  {32'h3e6c48b5, 32'hbe033c0f} /* (31, 17, 6) {real, imag} */,
  {32'h3d991868, 32'hbdc42bb2} /* (31, 17, 5) {real, imag} */,
  {32'h3daf87ac, 32'h3e05e8a5} /* (31, 17, 4) {real, imag} */,
  {32'hbd3e9c4c, 32'h3e9a840d} /* (31, 17, 3) {real, imag} */,
  {32'h3ce19fd8, 32'h3d9e5058} /* (31, 17, 2) {real, imag} */,
  {32'hbe92b414, 32'hbd8fe061} /* (31, 17, 1) {real, imag} */,
  {32'hbe0948b2, 32'h3e1a678d} /* (31, 17, 0) {real, imag} */,
  {32'h3db35242, 32'h3db35c43} /* (31, 16, 31) {real, imag} */,
  {32'hbe3771b3, 32'h3d842732} /* (31, 16, 30) {real, imag} */,
  {32'h3e801190, 32'h3da8a1b2} /* (31, 16, 29) {real, imag} */,
  {32'h3daa207f, 32'h3e3b70a8} /* (31, 16, 28) {real, imag} */,
  {32'h3ce87118, 32'h3ca5d780} /* (31, 16, 27) {real, imag} */,
  {32'h3e1c574a, 32'hbd39b54e} /* (31, 16, 26) {real, imag} */,
  {32'h3d90fa58, 32'hbe092f70} /* (31, 16, 25) {real, imag} */,
  {32'h3e2255bf, 32'h3eac6e22} /* (31, 16, 24) {real, imag} */,
  {32'hbdaeae0c, 32'hbe497008} /* (31, 16, 23) {real, imag} */,
  {32'hbe52f68a, 32'h3dfcd688} /* (31, 16, 22) {real, imag} */,
  {32'h3d47a490, 32'hbe12958d} /* (31, 16, 21) {real, imag} */,
  {32'h3dc599f2, 32'h3d7a860c} /* (31, 16, 20) {real, imag} */,
  {32'h3df1a6bb, 32'hbd9ccfed} /* (31, 16, 19) {real, imag} */,
  {32'h3e7c737d, 32'h3cdcece8} /* (31, 16, 18) {real, imag} */,
  {32'hbe2b9d15, 32'hbd949a13} /* (31, 16, 17) {real, imag} */,
  {32'hbe2670fc, 32'h00000000} /* (31, 16, 16) {real, imag} */,
  {32'hbe2b9d15, 32'h3d949a13} /* (31, 16, 15) {real, imag} */,
  {32'h3e7c737d, 32'hbcdcece8} /* (31, 16, 14) {real, imag} */,
  {32'h3df1a6bb, 32'h3d9ccfed} /* (31, 16, 13) {real, imag} */,
  {32'h3dc599f2, 32'hbd7a860c} /* (31, 16, 12) {real, imag} */,
  {32'h3d47a490, 32'h3e12958d} /* (31, 16, 11) {real, imag} */,
  {32'hbe52f68a, 32'hbdfcd688} /* (31, 16, 10) {real, imag} */,
  {32'hbdaeae0c, 32'h3e497008} /* (31, 16, 9) {real, imag} */,
  {32'h3e2255bf, 32'hbeac6e22} /* (31, 16, 8) {real, imag} */,
  {32'h3d90fa58, 32'h3e092f70} /* (31, 16, 7) {real, imag} */,
  {32'h3e1c574a, 32'h3d39b54e} /* (31, 16, 6) {real, imag} */,
  {32'h3ce87118, 32'hbca5d780} /* (31, 16, 5) {real, imag} */,
  {32'h3daa207f, 32'hbe3b70a8} /* (31, 16, 4) {real, imag} */,
  {32'h3e801190, 32'hbda8a1b2} /* (31, 16, 3) {real, imag} */,
  {32'hbe3771b3, 32'hbd842732} /* (31, 16, 2) {real, imag} */,
  {32'h3db35242, 32'hbdb35c43} /* (31, 16, 1) {real, imag} */,
  {32'hbee215fa, 32'h00000000} /* (31, 16, 0) {real, imag} */,
  {32'hbe92b414, 32'h3d8fe061} /* (31, 15, 31) {real, imag} */,
  {32'h3ce19fd8, 32'hbd9e5058} /* (31, 15, 30) {real, imag} */,
  {32'hbd3e9c4c, 32'hbe9a840d} /* (31, 15, 29) {real, imag} */,
  {32'h3daf87ac, 32'hbe05e8a5} /* (31, 15, 28) {real, imag} */,
  {32'h3d991868, 32'h3dc42bb2} /* (31, 15, 27) {real, imag} */,
  {32'h3e6c48b5, 32'h3e033c0f} /* (31, 15, 26) {real, imag} */,
  {32'hbe25a7ee, 32'hbe0fa31e} /* (31, 15, 25) {real, imag} */,
  {32'hbd5bea20, 32'h3d30d2f8} /* (31, 15, 24) {real, imag} */,
  {32'h3ddad27c, 32'hbe6f4fdd} /* (31, 15, 23) {real, imag} */,
  {32'h3d5d7938, 32'h3e5890eb} /* (31, 15, 22) {real, imag} */,
  {32'h3e4bbabb, 32'hbe3b11bf} /* (31, 15, 21) {real, imag} */,
  {32'h3d523c7f, 32'h3e8f67df} /* (31, 15, 20) {real, imag} */,
  {32'h3b4e6b00, 32'hbe0753f7} /* (31, 15, 19) {real, imag} */,
  {32'hbe1f0069, 32'h3e83ae12} /* (31, 15, 18) {real, imag} */,
  {32'h3dc5f59a, 32'hbe78547c} /* (31, 15, 17) {real, imag} */,
  {32'h3c8a84ac, 32'h3d6cb748} /* (31, 15, 16) {real, imag} */,
  {32'hbcb18148, 32'hbdf88808} /* (31, 15, 15) {real, imag} */,
  {32'h3d80daef, 32'h3ec26d7a} /* (31, 15, 14) {real, imag} */,
  {32'hbe0f8b84, 32'hbe181a4e} /* (31, 15, 13) {real, imag} */,
  {32'h3deae666, 32'h3e95cad1} /* (31, 15, 12) {real, imag} */,
  {32'h3e85b139, 32'hbda74b7c} /* (31, 15, 11) {real, imag} */,
  {32'hbe0b75ea, 32'hbd1200e4} /* (31, 15, 10) {real, imag} */,
  {32'h3e220942, 32'h3ddf8dbe} /* (31, 15, 9) {real, imag} */,
  {32'hbe6f167a, 32'h3c7a0940} /* (31, 15, 8) {real, imag} */,
  {32'h3e29fbe4, 32'hbe922d20} /* (31, 15, 7) {real, imag} */,
  {32'h3e2e9c56, 32'h3daf9e12} /* (31, 15, 6) {real, imag} */,
  {32'h3d9487ef, 32'h3d43c96c} /* (31, 15, 5) {real, imag} */,
  {32'h3cd3b3e0, 32'h3dee7580} /* (31, 15, 4) {real, imag} */,
  {32'h3d014068, 32'h3da5de1e} /* (31, 15, 3) {real, imag} */,
  {32'hbbdbfb60, 32'hbdfef370} /* (31, 15, 2) {real, imag} */,
  {32'h3df4a53b, 32'h3e04cc7a} /* (31, 15, 1) {real, imag} */,
  {32'hbe0948b2, 32'hbe1a678d} /* (31, 15, 0) {real, imag} */,
  {32'hbe735f1a, 32'hbda968e9} /* (31, 14, 31) {real, imag} */,
  {32'h3e3c42c3, 32'h3e3b78df} /* (31, 14, 30) {real, imag} */,
  {32'hbe2c0c12, 32'hbda76470} /* (31, 14, 29) {real, imag} */,
  {32'hbeb65b50, 32'hbd99b62d} /* (31, 14, 28) {real, imag} */,
  {32'hbee1b329, 32'h3e417294} /* (31, 14, 27) {real, imag} */,
  {32'h3eee40ac, 32'h3e32cdec} /* (31, 14, 26) {real, imag} */,
  {32'h3dde656c, 32'h3e060b01} /* (31, 14, 25) {real, imag} */,
  {32'h3d9acde2, 32'hbe727ffb} /* (31, 14, 24) {real, imag} */,
  {32'hbe874454, 32'h3dc751d2} /* (31, 14, 23) {real, imag} */,
  {32'h3eba0946, 32'h3ef8b440} /* (31, 14, 22) {real, imag} */,
  {32'h3d1be65a, 32'hbe23716b} /* (31, 14, 21) {real, imag} */,
  {32'hbe91509c, 32'h3d88059a} /* (31, 14, 20) {real, imag} */,
  {32'hbdcca990, 32'h3ef35c1c} /* (31, 14, 19) {real, imag} */,
  {32'hbe125510, 32'h3b3a12a0} /* (31, 14, 18) {real, imag} */,
  {32'hbe37c90e, 32'hbd8fe72c} /* (31, 14, 17) {real, imag} */,
  {32'hbda0b9a0, 32'h3e84032c} /* (31, 14, 16) {real, imag} */,
  {32'hbe17802f, 32'hbd47bf90} /* (31, 14, 15) {real, imag} */,
  {32'h3c7086c0, 32'hbeceb670} /* (31, 14, 14) {real, imag} */,
  {32'h3dd01aa2, 32'h3ee3deb6} /* (31, 14, 13) {real, imag} */,
  {32'h3b31bcc0, 32'h3da7ea2e} /* (31, 14, 12) {real, imag} */,
  {32'hbe1bceac, 32'hbd63da30} /* (31, 14, 11) {real, imag} */,
  {32'h3e9751a8, 32'h3db1307c} /* (31, 14, 10) {real, imag} */,
  {32'h3eaf36b2, 32'h3de82970} /* (31, 14, 9) {real, imag} */,
  {32'h3e3b7a3a, 32'hbc817220} /* (31, 14, 8) {real, imag} */,
  {32'hbeb3f133, 32'h3f3296e0} /* (31, 14, 7) {real, imag} */,
  {32'hbebb58ff, 32'h3d4cc574} /* (31, 14, 6) {real, imag} */,
  {32'h3eab6264, 32'h3e97f7ec} /* (31, 14, 5) {real, imag} */,
  {32'h3d4a79ae, 32'hbe6f80ca} /* (31, 14, 4) {real, imag} */,
  {32'h3e83903f, 32'h3e2cb238} /* (31, 14, 3) {real, imag} */,
  {32'h3e293009, 32'h3d7e9298} /* (31, 14, 2) {real, imag} */,
  {32'h3e81bf84, 32'hbe0b7d9b} /* (31, 14, 1) {real, imag} */,
  {32'hbdcce2f7, 32'hbdf42a7a} /* (31, 14, 0) {real, imag} */,
  {32'hbe580b49, 32'hbe24a311} /* (31, 13, 31) {real, imag} */,
  {32'hbee6f562, 32'h3dcfa33c} /* (31, 13, 30) {real, imag} */,
  {32'h3e9e1c76, 32'hbb8577a8} /* (31, 13, 29) {real, imag} */,
  {32'h3b2664c0, 32'h3da0a082} /* (31, 13, 28) {real, imag} */,
  {32'h3ce8bb7a, 32'hbe9442a4} /* (31, 13, 27) {real, imag} */,
  {32'h3e1b2502, 32'hbea7c662} /* (31, 13, 26) {real, imag} */,
  {32'hbc7d8678, 32'hbd637ce8} /* (31, 13, 25) {real, imag} */,
  {32'hbde4bd6c, 32'hbe6d93fc} /* (31, 13, 24) {real, imag} */,
  {32'h3dae39ce, 32'hbd9df376} /* (31, 13, 23) {real, imag} */,
  {32'hbb682a60, 32'hbdf0add0} /* (31, 13, 22) {real, imag} */,
  {32'hbd8bea62, 32'hbe9ebb67} /* (31, 13, 21) {real, imag} */,
  {32'h3e12d966, 32'hbcb3c830} /* (31, 13, 20) {real, imag} */,
  {32'h3ee9b856, 32'h3e557d13} /* (31, 13, 19) {real, imag} */,
  {32'h3f171075, 32'hbe4809a3} /* (31, 13, 18) {real, imag} */,
  {32'h3e166334, 32'hbe827db3} /* (31, 13, 17) {real, imag} */,
  {32'hbd2e0778, 32'h3ea66b70} /* (31, 13, 16) {real, imag} */,
  {32'hbe2d712a, 32'hbc8bea74} /* (31, 13, 15) {real, imag} */,
  {32'h3e260478, 32'h3c04a4ac} /* (31, 13, 14) {real, imag} */,
  {32'hbec929d3, 32'hbdc2d611} /* (31, 13, 13) {real, imag} */,
  {32'hbe03d163, 32'h3c01be44} /* (31, 13, 12) {real, imag} */,
  {32'hbe9ccd3e, 32'h3e1bca84} /* (31, 13, 11) {real, imag} */,
  {32'h3d1e061c, 32'h3d97175f} /* (31, 13, 10) {real, imag} */,
  {32'h3ea51077, 32'hbe23cb33} /* (31, 13, 9) {real, imag} */,
  {32'hbebc521a, 32'hbd7faf34} /* (31, 13, 8) {real, imag} */,
  {32'h3e97f0f1, 32'hbc992d38} /* (31, 13, 7) {real, imag} */,
  {32'hbdb47838, 32'h3d2bb318} /* (31, 13, 6) {real, imag} */,
  {32'hbe9c26dd, 32'hbd24c24c} /* (31, 13, 5) {real, imag} */,
  {32'hbe6f1cd4, 32'h3c49b078} /* (31, 13, 4) {real, imag} */,
  {32'hbdc64b7b, 32'h3e2b7c00} /* (31, 13, 3) {real, imag} */,
  {32'h3d2b63d0, 32'hbce2140e} /* (31, 13, 2) {real, imag} */,
  {32'h3e581b6a, 32'hbd31fd74} /* (31, 13, 1) {real, imag} */,
  {32'hbe7e0ebe, 32'hbd1b3684} /* (31, 13, 0) {real, imag} */,
  {32'h3d80ec8a, 32'hbe21efa1} /* (31, 12, 31) {real, imag} */,
  {32'h3e9c4160, 32'h3e8a4e9d} /* (31, 12, 30) {real, imag} */,
  {32'h3e2ad024, 32'hbd6399a8} /* (31, 12, 29) {real, imag} */,
  {32'hbe8a7620, 32'hbef3d52d} /* (31, 12, 28) {real, imag} */,
  {32'h3e1d1826, 32'hbe5b0090} /* (31, 12, 27) {real, imag} */,
  {32'hbc094928, 32'hbe16d987} /* (31, 12, 26) {real, imag} */,
  {32'h3c95e1c8, 32'h3ee82ee6} /* (31, 12, 25) {real, imag} */,
  {32'hbe50279e, 32'hbeb709e2} /* (31, 12, 24) {real, imag} */,
  {32'h3d4cdd22, 32'hbd1f3a48} /* (31, 12, 23) {real, imag} */,
  {32'hbd03b0a0, 32'h3e878050} /* (31, 12, 22) {real, imag} */,
  {32'h3e98e874, 32'h3e89367a} /* (31, 12, 21) {real, imag} */,
  {32'hbe645933, 32'h3ea1384f} /* (31, 12, 20) {real, imag} */,
  {32'hbf050658, 32'hbdf63ff8} /* (31, 12, 19) {real, imag} */,
  {32'hbeede012, 32'hbc974a9c} /* (31, 12, 18) {real, imag} */,
  {32'h3e3de3ee, 32'hbe168084} /* (31, 12, 17) {real, imag} */,
  {32'h3e0742f1, 32'hbdb11834} /* (31, 12, 16) {real, imag} */,
  {32'hbe792e4c, 32'h3e15de98} /* (31, 12, 15) {real, imag} */,
  {32'h3da7b070, 32'h3e8028b7} /* (31, 12, 14) {real, imag} */,
  {32'hbef8413e, 32'h3e1d2f8d} /* (31, 12, 13) {real, imag} */,
  {32'hbe24d572, 32'h3e1b5ac0} /* (31, 12, 12) {real, imag} */,
  {32'h3e4ceeb6, 32'hbe1d76f5} /* (31, 12, 11) {real, imag} */,
  {32'h3e3589ae, 32'h3e956562} /* (31, 12, 10) {real, imag} */,
  {32'hbb0d6120, 32'hbee156ec} /* (31, 12, 9) {real, imag} */,
  {32'h3dff55dc, 32'h3e9a0719} /* (31, 12, 8) {real, imag} */,
  {32'hbe88fbc3, 32'hbea4c18d} /* (31, 12, 7) {real, imag} */,
  {32'h3c358d80, 32'hbe3a8861} /* (31, 12, 6) {real, imag} */,
  {32'h3c69c1c0, 32'hbd809b30} /* (31, 12, 5) {real, imag} */,
  {32'h3d580b50, 32'hbe04a77d} /* (31, 12, 4) {real, imag} */,
  {32'hbe564c01, 32'h3c06f570} /* (31, 12, 3) {real, imag} */,
  {32'hbed89a43, 32'hbd24cdc4} /* (31, 12, 2) {real, imag} */,
  {32'hbdd43cf8, 32'h3ebf0ac8} /* (31, 12, 1) {real, imag} */,
  {32'h3dec86e8, 32'h3d5ee5a0} /* (31, 12, 0) {real, imag} */,
  {32'h3da8efb0, 32'hbe4c6be4} /* (31, 11, 31) {real, imag} */,
  {32'hbde53658, 32'h3ec37cfc} /* (31, 11, 30) {real, imag} */,
  {32'h3da0c944, 32'h3e2d8e7a} /* (31, 11, 29) {real, imag} */,
  {32'hbe85a598, 32'h3e954e42} /* (31, 11, 28) {real, imag} */,
  {32'hbce0ec54, 32'h3bfca8c0} /* (31, 11, 27) {real, imag} */,
  {32'hbdc356a4, 32'hbe023a46} /* (31, 11, 26) {real, imag} */,
  {32'hbf014fd7, 32'h3e088f4e} /* (31, 11, 25) {real, imag} */,
  {32'h3e0376c0, 32'hbe80dec2} /* (31, 11, 24) {real, imag} */,
  {32'h3d4f8258, 32'h3f02107c} /* (31, 11, 23) {real, imag} */,
  {32'hbc509060, 32'hbcfaff60} /* (31, 11, 22) {real, imag} */,
  {32'h3e92f17d, 32'h3ee39db0} /* (31, 11, 21) {real, imag} */,
  {32'hbe3e6374, 32'h3e5bb608} /* (31, 11, 20) {real, imag} */,
  {32'hbdfdc950, 32'hbef6c5f8} /* (31, 11, 19) {real, imag} */,
  {32'hbc40bd30, 32'hbe86079f} /* (31, 11, 18) {real, imag} */,
  {32'h3d66146c, 32'h3dd5fabb} /* (31, 11, 17) {real, imag} */,
  {32'h3cfb1668, 32'h3d05a969} /* (31, 11, 16) {real, imag} */,
  {32'h3c9997e4, 32'hbd8a0578} /* (31, 11, 15) {real, imag} */,
  {32'hbec6cd51, 32'hbd02daf4} /* (31, 11, 14) {real, imag} */,
  {32'hbea4ae6e, 32'hbe43f882} /* (31, 11, 13) {real, imag} */,
  {32'hbe68ec32, 32'hbf4ddde0} /* (31, 11, 12) {real, imag} */,
  {32'h3e31c0c8, 32'h3efdb588} /* (31, 11, 11) {real, imag} */,
  {32'h3f1546ee, 32'h3e7efc90} /* (31, 11, 10) {real, imag} */,
  {32'hbdac9ad2, 32'hbd7942dc} /* (31, 11, 9) {real, imag} */,
  {32'h3e41b487, 32'hbcadbd94} /* (31, 11, 8) {real, imag} */,
  {32'hbe631f3a, 32'hbe93480f} /* (31, 11, 7) {real, imag} */,
  {32'h3d6bae20, 32'h3e1bf936} /* (31, 11, 6) {real, imag} */,
  {32'h3e87d1fd, 32'hbe7b2ea3} /* (31, 11, 5) {real, imag} */,
  {32'h3e25fa2a, 32'h3ed776c7} /* (31, 11, 4) {real, imag} */,
  {32'h3e08b553, 32'hbd42f370} /* (31, 11, 3) {real, imag} */,
  {32'hbe433bf4, 32'h3deb53c8} /* (31, 11, 2) {real, imag} */,
  {32'hbda1a8e4, 32'h3dca40bc} /* (31, 11, 1) {real, imag} */,
  {32'h3d8acf98, 32'hbe302c98} /* (31, 11, 0) {real, imag} */,
  {32'hbdb7182e, 32'h3ed5751c} /* (31, 10, 31) {real, imag} */,
  {32'h3d485468, 32'h3dc09008} /* (31, 10, 30) {real, imag} */,
  {32'hbc95a9f0, 32'h3df6f8b6} /* (31, 10, 29) {real, imag} */,
  {32'h3efaab8a, 32'hbddd56f4} /* (31, 10, 28) {real, imag} */,
  {32'hbdcce049, 32'hbed29c58} /* (31, 10, 27) {real, imag} */,
  {32'hbd6d302c, 32'h3e873d2c} /* (31, 10, 26) {real, imag} */,
  {32'hbdbf5fa4, 32'hbe6bcc2c} /* (31, 10, 25) {real, imag} */,
  {32'hbdd65b06, 32'hbd305448} /* (31, 10, 24) {real, imag} */,
  {32'hbf0732e3, 32'h3e92e901} /* (31, 10, 23) {real, imag} */,
  {32'h3eb605f8, 32'hbda8a82e} /* (31, 10, 22) {real, imag} */,
  {32'hbed91886, 32'hbe357960} /* (31, 10, 21) {real, imag} */,
  {32'hbe4dc24c, 32'h3ee1f6d6} /* (31, 10, 20) {real, imag} */,
  {32'h3d729148, 32'hbeb5247e} /* (31, 10, 19) {real, imag} */,
  {32'h3e49545a, 32'hbe7fc24c} /* (31, 10, 18) {real, imag} */,
  {32'hbe383a84, 32'hbdabd4e2} /* (31, 10, 17) {real, imag} */,
  {32'hbdc78fae, 32'h3dbb0c29} /* (31, 10, 16) {real, imag} */,
  {32'hbc8d18d3, 32'hbc95a1f8} /* (31, 10, 15) {real, imag} */,
  {32'hbd3eac1c, 32'hbc958a18} /* (31, 10, 14) {real, imag} */,
  {32'h3c9332f0, 32'h3ed26b2c} /* (31, 10, 13) {real, imag} */,
  {32'hbe5003ac, 32'h3ec2e57a} /* (31, 10, 12) {real, imag} */,
  {32'hbe20c3c1, 32'hbe04d479} /* (31, 10, 11) {real, imag} */,
  {32'hbe9be0ba, 32'hbca67df0} /* (31, 10, 10) {real, imag} */,
  {32'h3e499dcc, 32'h3ea66e8c} /* (31, 10, 9) {real, imag} */,
  {32'hbdcb8329, 32'hbe1ed2ac} /* (31, 10, 8) {real, imag} */,
  {32'h3e8499a7, 32'h3e9ac8ae} /* (31, 10, 7) {real, imag} */,
  {32'hbe32ae8a, 32'hbea80efc} /* (31, 10, 6) {real, imag} */,
  {32'h3c417f20, 32'hbe2459bc} /* (31, 10, 5) {real, imag} */,
  {32'hbd021650, 32'h3e504090} /* (31, 10, 4) {real, imag} */,
  {32'h3eefcaff, 32'hbe1234fb} /* (31, 10, 3) {real, imag} */,
  {32'h3ca92820, 32'hbe899ad6} /* (31, 10, 2) {real, imag} */,
  {32'h3efb2137, 32'hbde2948a} /* (31, 10, 1) {real, imag} */,
  {32'hbe9b69de, 32'h3d716ea6} /* (31, 10, 0) {real, imag} */,
  {32'hbd151e64, 32'h3f306eab} /* (31, 9, 31) {real, imag} */,
  {32'h3dbbd282, 32'h3e75aaae} /* (31, 9, 30) {real, imag} */,
  {32'h3ed3cc2b, 32'h3da51eb4} /* (31, 9, 29) {real, imag} */,
  {32'h3f0b52f8, 32'h3e8fa040} /* (31, 9, 28) {real, imag} */,
  {32'h3e75c4d8, 32'hbe7e20d1} /* (31, 9, 27) {real, imag} */,
  {32'h3e08c8e4, 32'h3e67a1cc} /* (31, 9, 26) {real, imag} */,
  {32'h3daeeba3, 32'h3aa42480} /* (31, 9, 25) {real, imag} */,
  {32'h3d8aae08, 32'hbd6de7f4} /* (31, 9, 24) {real, imag} */,
  {32'hbd974a9c, 32'h3d3cfafe} /* (31, 9, 23) {real, imag} */,
  {32'h3b21e380, 32'h3e128605} /* (31, 9, 22) {real, imag} */,
  {32'h3e64eb5c, 32'hbe6de0ce} /* (31, 9, 21) {real, imag} */,
  {32'h3d2d2ad0, 32'hbe0c6ea8} /* (31, 9, 20) {real, imag} */,
  {32'hbec8ab2c, 32'hbe148950} /* (31, 9, 19) {real, imag} */,
  {32'hbe472524, 32'hbd368b96} /* (31, 9, 18) {real, imag} */,
  {32'h3e994d99, 32'hbdbecb92} /* (31, 9, 17) {real, imag} */,
  {32'h3d6b3254, 32'hbd606e7c} /* (31, 9, 16) {real, imag} */,
  {32'h3d6fa734, 32'hbdb7f21d} /* (31, 9, 15) {real, imag} */,
  {32'h3e663a16, 32'hbd42c578} /* (31, 9, 14) {real, imag} */,
  {32'h3f05fe52, 32'hbbb170a0} /* (31, 9, 13) {real, imag} */,
  {32'hbd7bc24e, 32'hbec22173} /* (31, 9, 12) {real, imag} */,
  {32'h3e0f7852, 32'hbca32ec4} /* (31, 9, 11) {real, imag} */,
  {32'h3dcac83a, 32'h3d9e7aaa} /* (31, 9, 10) {real, imag} */,
  {32'h3de8b5d8, 32'hbeb5b0c7} /* (31, 9, 9) {real, imag} */,
  {32'hbe70dc44, 32'hbebd8d9c} /* (31, 9, 8) {real, imag} */,
  {32'h3ef12da5, 32'hbe48d34e} /* (31, 9, 7) {real, imag} */,
  {32'hbea282da, 32'hbdfe8882} /* (31, 9, 6) {real, imag} */,
  {32'hbdf3cc42, 32'hbb8c8420} /* (31, 9, 5) {real, imag} */,
  {32'h3f18b11b, 32'hbcce8150} /* (31, 9, 4) {real, imag} */,
  {32'hbf521346, 32'h3e096349} /* (31, 9, 3) {real, imag} */,
  {32'hbdff7808, 32'hbf04fa9e} /* (31, 9, 2) {real, imag} */,
  {32'h3e4c622c, 32'hbd185c98} /* (31, 9, 1) {real, imag} */,
  {32'h3c6423a0, 32'h3ea98906} /* (31, 9, 0) {real, imag} */,
  {32'hbf50e843, 32'hbf24fb94} /* (31, 8, 31) {real, imag} */,
  {32'h3f884781, 32'hbdf5c13c} /* (31, 8, 30) {real, imag} */,
  {32'hbe6482e0, 32'h3cece152} /* (31, 8, 29) {real, imag} */,
  {32'hbedf86e0, 32'h3e9cb912} /* (31, 8, 28) {real, imag} */,
  {32'h3e1bef4b, 32'h3de0721f} /* (31, 8, 27) {real, imag} */,
  {32'hbedea0ef, 32'hbd17d3d0} /* (31, 8, 26) {real, imag} */,
  {32'h3e72cd22, 32'hbbceb150} /* (31, 8, 25) {real, imag} */,
  {32'hbe492ac2, 32'hbdb77b80} /* (31, 8, 24) {real, imag} */,
  {32'h3db7007c, 32'h3e8f0ba4} /* (31, 8, 23) {real, imag} */,
  {32'h3e1babf0, 32'hbe5466b6} /* (31, 8, 22) {real, imag} */,
  {32'hbe64b441, 32'h3d17b2cf} /* (31, 8, 21) {real, imag} */,
  {32'hbd7dd8d0, 32'h3df5aaaa} /* (31, 8, 20) {real, imag} */,
  {32'hbdb9c6be, 32'h3db1a2e4} /* (31, 8, 19) {real, imag} */,
  {32'hbe390fcc, 32'h3e1af45e} /* (31, 8, 18) {real, imag} */,
  {32'h3e8095c5, 32'h3edd26c9} /* (31, 8, 17) {real, imag} */,
  {32'hbd452614, 32'hbdd26313} /* (31, 8, 16) {real, imag} */,
  {32'hbd0ba3a0, 32'hbd2a554a} /* (31, 8, 15) {real, imag} */,
  {32'h3d691e8c, 32'h3d8c5802} /* (31, 8, 14) {real, imag} */,
  {32'h3e08d7d6, 32'hbd60e870} /* (31, 8, 13) {real, imag} */,
  {32'hbc036b80, 32'h3e915e94} /* (31, 8, 12) {real, imag} */,
  {32'hbe549f56, 32'h3e4cf1b2} /* (31, 8, 11) {real, imag} */,
  {32'hbd2b4bc4, 32'h3e915521} /* (31, 8, 10) {real, imag} */,
  {32'h3da8504e, 32'hbe078ba2} /* (31, 8, 9) {real, imag} */,
  {32'h3d570de0, 32'hbe756abe} /* (31, 8, 8) {real, imag} */,
  {32'hbd945f40, 32'hbebbd7cf} /* (31, 8, 7) {real, imag} */,
  {32'h3eaf152f, 32'h3e174dd7} /* (31, 8, 6) {real, imag} */,
  {32'h3d66175a, 32'h3e6e92c0} /* (31, 8, 5) {real, imag} */,
  {32'h3e42184c, 32'h3e49c841} /* (31, 8, 4) {real, imag} */,
  {32'hbf44b78b, 32'hbd6e5298} /* (31, 8, 3) {real, imag} */,
  {32'h3ed94f0e, 32'h3f94167c} /* (31, 8, 2) {real, imag} */,
  {32'hbf1a969c, 32'hbeedb412} /* (31, 8, 1) {real, imag} */,
  {32'hbf114c26, 32'h3a421600} /* (31, 8, 0) {real, imag} */,
  {32'h3e67ff8e, 32'h3bda9460} /* (31, 7, 31) {real, imag} */,
  {32'hbe313a1e, 32'hbe2653c2} /* (31, 7, 30) {real, imag} */,
  {32'h3d67df34, 32'hbcf80128} /* (31, 7, 29) {real, imag} */,
  {32'hbedbaf1b, 32'h3d49e580} /* (31, 7, 28) {real, imag} */,
  {32'hbe7785e5, 32'hbe4e5842} /* (31, 7, 27) {real, imag} */,
  {32'h3e8a5bc2, 32'h3e582780} /* (31, 7, 26) {real, imag} */,
  {32'h3e479370, 32'hbd6b8a66} /* (31, 7, 25) {real, imag} */,
  {32'hbe42e356, 32'h3ebc8bcd} /* (31, 7, 24) {real, imag} */,
  {32'h3e9f2d74, 32'h3dcb695e} /* (31, 7, 23) {real, imag} */,
  {32'hbe0df467, 32'h3c9b1934} /* (31, 7, 22) {real, imag} */,
  {32'hbd08a6e0, 32'h3ea3dc38} /* (31, 7, 21) {real, imag} */,
  {32'hbe8a01ef, 32'hbe1af006} /* (31, 7, 20) {real, imag} */,
  {32'hbd683328, 32'h3e644fbc} /* (31, 7, 19) {real, imag} */,
  {32'hbe20c473, 32'h3e40fea0} /* (31, 7, 18) {real, imag} */,
  {32'h3ee6fd63, 32'h3e38346a} /* (31, 7, 17) {real, imag} */,
  {32'h3d85a819, 32'hbdb4fd79} /* (31, 7, 16) {real, imag} */,
  {32'h3d99860d, 32'h3e30dd6d} /* (31, 7, 15) {real, imag} */,
  {32'hbe739be6, 32'h3e910df6} /* (31, 7, 14) {real, imag} */,
  {32'hbe4dd438, 32'hbdb2e3e0} /* (31, 7, 13) {real, imag} */,
  {32'hbd719626, 32'hbe31cac9} /* (31, 7, 12) {real, imag} */,
  {32'h3eb6823c, 32'h3d750374} /* (31, 7, 11) {real, imag} */,
  {32'h3e78dbc1, 32'h3a941200} /* (31, 7, 10) {real, imag} */,
  {32'hbe54eccd, 32'hbe90d042} /* (31, 7, 9) {real, imag} */,
  {32'hbe378ca5, 32'h3e2c7309} /* (31, 7, 8) {real, imag} */,
  {32'h3d1a2034, 32'hbd3470e4} /* (31, 7, 7) {real, imag} */,
  {32'h3e41bab5, 32'hbdb31082} /* (31, 7, 6) {real, imag} */,
  {32'h3e89c6b4, 32'hbc2c5f60} /* (31, 7, 5) {real, imag} */,
  {32'h3e1e1d5e, 32'hbca80c30} /* (31, 7, 4) {real, imag} */,
  {32'h3e9f2e3e, 32'h3c3c42c0} /* (31, 7, 3) {real, imag} */,
  {32'h3ea93268, 32'hbe965ef5} /* (31, 7, 2) {real, imag} */,
  {32'hbe7ba278, 32'h3d5f8b58} /* (31, 7, 1) {real, imag} */,
  {32'h3f3c68b9, 32'h3eddbf4f} /* (31, 7, 0) {real, imag} */,
  {32'hbe9e14ac, 32'h3f190a00} /* (31, 6, 31) {real, imag} */,
  {32'hbef93ef2, 32'hbf12f0bd} /* (31, 6, 30) {real, imag} */,
  {32'h3ed501e8, 32'h3c9024a0} /* (31, 6, 29) {real, imag} */,
  {32'hbdb79818, 32'h3dd32e6a} /* (31, 6, 28) {real, imag} */,
  {32'hbe240e4c, 32'h3e478610} /* (31, 6, 27) {real, imag} */,
  {32'h3e73b8d0, 32'h3f05d8c4} /* (31, 6, 26) {real, imag} */,
  {32'hbd673422, 32'hbdf3e94a} /* (31, 6, 25) {real, imag} */,
  {32'h3e2e60dc, 32'h3e595abe} /* (31, 6, 24) {real, imag} */,
  {32'hbe1a798c, 32'hbee5a3df} /* (31, 6, 23) {real, imag} */,
  {32'h3d239282, 32'hbea10a6a} /* (31, 6, 22) {real, imag} */,
  {32'h3ea2b3a2, 32'hbec95768} /* (31, 6, 21) {real, imag} */,
  {32'hbeb1d34a, 32'hbc80427a} /* (31, 6, 20) {real, imag} */,
  {32'hbeb00fbd, 32'hbcdb33f8} /* (31, 6, 19) {real, imag} */,
  {32'h3cabda52, 32'h3e784644} /* (31, 6, 18) {real, imag} */,
  {32'hbe310418, 32'hbea579d2} /* (31, 6, 17) {real, imag} */,
  {32'h3de3b9c0, 32'h3d528bf4} /* (31, 6, 16) {real, imag} */,
  {32'h3e2cefb7, 32'h3e5b3ad6} /* (31, 6, 15) {real, imag} */,
  {32'h3da81c76, 32'hbec47cdf} /* (31, 6, 14) {real, imag} */,
  {32'hbe88d089, 32'hbea82d26} /* (31, 6, 13) {real, imag} */,
  {32'hbe992283, 32'h3c83d8ac} /* (31, 6, 12) {real, imag} */,
  {32'hbcf641e8, 32'h3b9e9700} /* (31, 6, 11) {real, imag} */,
  {32'hbe541c83, 32'hbe81bad7} /* (31, 6, 10) {real, imag} */,
  {32'h3e094cfb, 32'hbb9c0a00} /* (31, 6, 9) {real, imag} */,
  {32'h3edcb0f2, 32'h3e89e8af} /* (31, 6, 8) {real, imag} */,
  {32'hbeeb66f3, 32'h3eb550c5} /* (31, 6, 7) {real, imag} */,
  {32'hbe69ead0, 32'hbcae1798} /* (31, 6, 6) {real, imag} */,
  {32'h3ebe0844, 32'h3eb9b7c6} /* (31, 6, 5) {real, imag} */,
  {32'hbd9133dc, 32'h3e443be0} /* (31, 6, 4) {real, imag} */,
  {32'h3e203cb0, 32'h3db1741e} /* (31, 6, 3) {real, imag} */,
  {32'hbd742db6, 32'hbf3a80eb} /* (31, 6, 2) {real, imag} */,
  {32'hbf0981a3, 32'hbe08c332} /* (31, 6, 1) {real, imag} */,
  {32'h3f0b9ecc, 32'hbe894da7} /* (31, 6, 0) {real, imag} */,
  {32'hbfcaf712, 32'hbdd0c9e2} /* (31, 5, 31) {real, imag} */,
  {32'h3e8b8b90, 32'hbf094173} /* (31, 5, 30) {real, imag} */,
  {32'hbd8cb030, 32'hbe5ec44c} /* (31, 5, 29) {real, imag} */,
  {32'hbd78d7b2, 32'hbf13d560} /* (31, 5, 28) {real, imag} */,
  {32'h3f35ed08, 32'hbda19d04} /* (31, 5, 27) {real, imag} */,
  {32'h3dda5d36, 32'h3ddd2658} /* (31, 5, 26) {real, imag} */,
  {32'hbe9f7293, 32'h3ec6d03c} /* (31, 5, 25) {real, imag} */,
  {32'hbe050512, 32'hbc2b8fb0} /* (31, 5, 24) {real, imag} */,
  {32'h3d9d31ad, 32'h3d635210} /* (31, 5, 23) {real, imag} */,
  {32'h3e489cda, 32'hbe9036b4} /* (31, 5, 22) {real, imag} */,
  {32'hbdf44fbb, 32'h3ec768a9} /* (31, 5, 21) {real, imag} */,
  {32'h3edb75a4, 32'hbeb22510} /* (31, 5, 20) {real, imag} */,
  {32'h3e776658, 32'hbd89a787} /* (31, 5, 19) {real, imag} */,
  {32'h3cc8afe8, 32'h3e0b4f34} /* (31, 5, 18) {real, imag} */,
  {32'hbdc538e9, 32'hbdb481fc} /* (31, 5, 17) {real, imag} */,
  {32'hbebeb538, 32'hbade6d00} /* (31, 5, 16) {real, imag} */,
  {32'hbdf0d2ba, 32'hbe4fe692} /* (31, 5, 15) {real, imag} */,
  {32'hbe714d14, 32'h3e14ddf8} /* (31, 5, 14) {real, imag} */,
  {32'hbdf78f8c, 32'h3e107087} /* (31, 5, 13) {real, imag} */,
  {32'h3e1ad9ac, 32'h3e2615b6} /* (31, 5, 12) {real, imag} */,
  {32'hbedaee64, 32'hbe2a447c} /* (31, 5, 11) {real, imag} */,
  {32'h3dd06fff, 32'h3e83cb71} /* (31, 5, 10) {real, imag} */,
  {32'h3d5a6cb6, 32'h3eae0e2d} /* (31, 5, 9) {real, imag} */,
  {32'hbd31666c, 32'h3ebe995e} /* (31, 5, 8) {real, imag} */,
  {32'h3ec64126, 32'hbf25b9b8} /* (31, 5, 7) {real, imag} */,
  {32'h3f05fe23, 32'h3e69b1fe} /* (31, 5, 6) {real, imag} */,
  {32'h3d47fd20, 32'h3ea3aa34} /* (31, 5, 5) {real, imag} */,
  {32'hbf4dd508, 32'hbe33407b} /* (31, 5, 4) {real, imag} */,
  {32'hbf36e6c7, 32'hbe59bee6} /* (31, 5, 3) {real, imag} */,
  {32'h3f9e150c, 32'h3f22426c} /* (31, 5, 2) {real, imag} */,
  {32'hbf9ae460, 32'hbf8d72c8} /* (31, 5, 1) {real, imag} */,
  {32'hbfb893cf, 32'h3e52dc80} /* (31, 5, 0) {real, imag} */,
  {32'h3f1c4ad8, 32'h3fb11866} /* (31, 4, 31) {real, imag} */,
  {32'hc00cd4ce, 32'hbe024a68} /* (31, 4, 30) {real, imag} */,
  {32'hbe8fbb80, 32'h3b366200} /* (31, 4, 29) {real, imag} */,
  {32'h3f6042af, 32'h3e7156a7} /* (31, 4, 28) {real, imag} */,
  {32'hbf0bfcda, 32'hbf051f03} /* (31, 4, 27) {real, imag} */,
  {32'hbea1d585, 32'hbe7b82a8} /* (31, 4, 26) {real, imag} */,
  {32'hbe87ea4e, 32'h3d626a54} /* (31, 4, 25) {real, imag} */,
  {32'hbd8fe500, 32'hbe456b6c} /* (31, 4, 24) {real, imag} */,
  {32'hbe8443ac, 32'h3d53453e} /* (31, 4, 23) {real, imag} */,
  {32'h3e7950e0, 32'h3ee09340} /* (31, 4, 22) {real, imag} */,
  {32'hbeae4620, 32'h3e40408f} /* (31, 4, 21) {real, imag} */,
  {32'h3f1eb55e, 32'hbeb29cf9} /* (31, 4, 20) {real, imag} */,
  {32'h3e4b28c2, 32'hbc8655f8} /* (31, 4, 19) {real, imag} */,
  {32'h3e0576ca, 32'hbe15ebf1} /* (31, 4, 18) {real, imag} */,
  {32'h3de45e95, 32'h3ed0588b} /* (31, 4, 17) {real, imag} */,
  {32'h3c0a9b1c, 32'hbddee748} /* (31, 4, 16) {real, imag} */,
  {32'hbdac984a, 32'hbe209fa2} /* (31, 4, 15) {real, imag} */,
  {32'h3e34afc2, 32'h3dc3539c} /* (31, 4, 14) {real, imag} */,
  {32'h3eedec7a, 32'hbd99efa9} /* (31, 4, 13) {real, imag} */,
  {32'h3e64a678, 32'hbec49646} /* (31, 4, 12) {real, imag} */,
  {32'h3ea55d38, 32'hbdfb0a90} /* (31, 4, 11) {real, imag} */,
  {32'hbec83aa2, 32'h3e082314} /* (31, 4, 10) {real, imag} */,
  {32'hbdfd92de, 32'h3e72a6ac} /* (31, 4, 9) {real, imag} */,
  {32'hbe8fa1f5, 32'h3ddddcf8} /* (31, 4, 8) {real, imag} */,
  {32'h3ebc07ec, 32'h3eb46270} /* (31, 4, 7) {real, imag} */,
  {32'hbd5b1d20, 32'h3e85cabc} /* (31, 4, 6) {real, imag} */,
  {32'h3ec9c876, 32'hbf3f98cf} /* (31, 4, 5) {real, imag} */,
  {32'hbc6ed220, 32'h3f4e1884} /* (31, 4, 4) {real, imag} */,
  {32'h3e44b08c, 32'h3f00d07c} /* (31, 4, 3) {real, imag} */,
  {32'hbf9d270a, 32'hbf8f271f} /* (31, 4, 2) {real, imag} */,
  {32'h400b97f5, 32'h3fdb3f8b} /* (31, 4, 1) {real, imag} */,
  {32'h3ff929bb, 32'h3ef78e14} /* (31, 4, 0) {real, imag} */,
  {32'hbfb608b6, 32'h3f772bdf} /* (31, 3, 31) {real, imag} */,
  {32'h3f33963e, 32'hbf8d7a5d} /* (31, 3, 30) {real, imag} */,
  {32'h3f68cefa, 32'h3d0fbcf8} /* (31, 3, 29) {real, imag} */,
  {32'h3e4e45fe, 32'h3f07ec76} /* (31, 3, 28) {real, imag} */,
  {32'hbe2dcfd6, 32'hbe9d4a9e} /* (31, 3, 27) {real, imag} */,
  {32'hbd828ff6, 32'hbe01c2d8} /* (31, 3, 26) {real, imag} */,
  {32'h3df30f8c, 32'hbd2cd130} /* (31, 3, 25) {real, imag} */,
  {32'h3dd299b0, 32'h3e56086c} /* (31, 3, 24) {real, imag} */,
  {32'hbe81ca50, 32'h3d797fac} /* (31, 3, 23) {real, imag} */,
  {32'h3ddce6d2, 32'h3e4b54ff} /* (31, 3, 22) {real, imag} */,
  {32'h3c10a1b8, 32'hbf0a7893} /* (31, 3, 21) {real, imag} */,
  {32'hbda9770b, 32'h3d6b5224} /* (31, 3, 20) {real, imag} */,
  {32'h3d7eee6c, 32'hbd1dff84} /* (31, 3, 19) {real, imag} */,
  {32'h3efcc18b, 32'hbed345b8} /* (31, 3, 18) {real, imag} */,
  {32'h3e239150, 32'hbde1ab12} /* (31, 3, 17) {real, imag} */,
  {32'hbdbd577a, 32'h3e031819} /* (31, 3, 16) {real, imag} */,
  {32'hbd7bca76, 32'hbdaced04} /* (31, 3, 15) {real, imag} */,
  {32'h3e8b7d17, 32'h3eb81d17} /* (31, 3, 14) {real, imag} */,
  {32'hbe667c76, 32'hbe49adce} /* (31, 3, 13) {real, imag} */,
  {32'hbe9260de, 32'hbdf6e638} /* (31, 3, 12) {real, imag} */,
  {32'h3df7c029, 32'hbe9e2e57} /* (31, 3, 11) {real, imag} */,
  {32'hbebe0bff, 32'hbe7308ea} /* (31, 3, 10) {real, imag} */,
  {32'hbdd561a2, 32'h3e477273} /* (31, 3, 9) {real, imag} */,
  {32'h3e93b4ba, 32'hbec30222} /* (31, 3, 8) {real, imag} */,
  {32'hbe9072bd, 32'h3e03d25f} /* (31, 3, 7) {real, imag} */,
  {32'hbe0a434c, 32'h3e34a165} /* (31, 3, 6) {real, imag} */,
  {32'hbf4fc8b4, 32'h3efdcb73} /* (31, 3, 5) {real, imag} */,
  {32'hbe4f0708, 32'h3e4fc6d6} /* (31, 3, 4) {real, imag} */,
  {32'h3f3d52ca, 32'hbeb569dc} /* (31, 3, 3) {real, imag} */,
  {32'hbf3bf5ae, 32'hbf343a34} /* (31, 3, 2) {real, imag} */,
  {32'h3f9bedbb, 32'hbcae9a40} /* (31, 3, 1) {real, imag} */,
  {32'h3e0c0d34, 32'h3f25b2a1} /* (31, 3, 0) {real, imag} */,
  {32'hc0ef6960, 32'hbfc168f2} /* (31, 2, 31) {real, imag} */,
  {32'h40819d18, 32'hc0149812} /* (31, 2, 30) {real, imag} */,
  {32'h3d2cdf70, 32'h3e2eaf80} /* (31, 2, 29) {real, imag} */,
  {32'hbfbfda9e, 32'h3fcd1a50} /* (31, 2, 28) {real, imag} */,
  {32'h3f6d2bd4, 32'h3d0c53b0} /* (31, 2, 27) {real, imag} */,
  {32'h3e6a6cf8, 32'h3e838de6} /* (31, 2, 26) {real, imag} */,
  {32'hbe0a9e1e, 32'hbe1fd663} /* (31, 2, 25) {real, imag} */,
  {32'h3f1b96c1, 32'hbe7b7fe6} /* (31, 2, 24) {real, imag} */,
  {32'h3eab479c, 32'h3d8c3dfa} /* (31, 2, 23) {real, imag} */,
  {32'hbef2f0ec, 32'hbc8e8310} /* (31, 2, 22) {real, imag} */,
  {32'h3ee2f668, 32'hbe61515c} /* (31, 2, 21) {real, imag} */,
  {32'hbd23ec68, 32'h3d2e130e} /* (31, 2, 20) {real, imag} */,
  {32'h3ee2f04c, 32'h3e019754} /* (31, 2, 19) {real, imag} */,
  {32'hbdeba101, 32'hbd66c780} /* (31, 2, 18) {real, imag} */,
  {32'h3e89e9f6, 32'hbd44be64} /* (31, 2, 17) {real, imag} */,
  {32'hbc631124, 32'hbccd4240} /* (31, 2, 16) {real, imag} */,
  {32'hbe86fac4, 32'hbd9b8682} /* (31, 2, 15) {real, imag} */,
  {32'h3e895751, 32'h3ec8427a} /* (31, 2, 14) {real, imag} */,
  {32'h3dc09b1c, 32'hbd4f5d8a} /* (31, 2, 13) {real, imag} */,
  {32'h3e5c355c, 32'h3e4dd14b} /* (31, 2, 12) {real, imag} */,
  {32'hbd34c15e, 32'h3e69df0e} /* (31, 2, 11) {real, imag} */,
  {32'hbd59caf4, 32'h3b1b3b10} /* (31, 2, 10) {real, imag} */,
  {32'hbe98dfc2, 32'h3eb158fd} /* (31, 2, 9) {real, imag} */,
  {32'h3f6f2bee, 32'h3e52222c} /* (31, 2, 8) {real, imag} */,
  {32'hbeabb2f7, 32'hbecb5111} /* (31, 2, 7) {real, imag} */,
  {32'h3e097e56, 32'h3eaed806} /* (31, 2, 6) {real, imag} */,
  {32'h3ed30186, 32'h3df37260} /* (31, 2, 5) {real, imag} */,
  {32'hbf36511c, 32'h3ea337df} /* (31, 2, 4) {real, imag} */,
  {32'hbf20ac18, 32'hbf80c31b} /* (31, 2, 3) {real, imag} */,
  {32'h405d3696, 32'h3e5124e8} /* (31, 2, 2) {real, imag} */,
  {32'hc0c99a5c, 32'h403d7840} /* (31, 2, 1) {real, imag} */,
  {32'hc0a76984, 32'hbf2d4ce4} /* (31, 2, 0) {real, imag} */,
  {32'h410493cc, 32'hc0380d32} /* (31, 1, 31) {real, imag} */,
  {32'hc06f09e9, 32'h3e982aed} /* (31, 1, 30) {real, imag} */,
  {32'hbe9bf57e, 32'h3ea5fb3a} /* (31, 1, 29) {real, imag} */,
  {32'h3f9a1c02, 32'hbe8caad7} /* (31, 1, 28) {real, imag} */,
  {32'hbf580064, 32'h3dda9e8c} /* (31, 1, 27) {real, imag} */,
  {32'hbd3810a0, 32'h3d7fde38} /* (31, 1, 26) {real, imag} */,
  {32'h3e1b413c, 32'hbee214f5} /* (31, 1, 25) {real, imag} */,
  {32'hbf006408, 32'hbe4e4434} /* (31, 1, 24) {real, imag} */,
  {32'hbf0af551, 32'hbd1eae88} /* (31, 1, 23) {real, imag} */,
  {32'h3db0aed2, 32'hbd5ba0ce} /* (31, 1, 22) {real, imag} */,
  {32'hbe347e5f, 32'h3e540cf9} /* (31, 1, 21) {real, imag} */,
  {32'h3ee2982f, 32'h3f04c0fc} /* (31, 1, 20) {real, imag} */,
  {32'hbf0ff067, 32'h3e9a0dd8} /* (31, 1, 19) {real, imag} */,
  {32'h3d1663be, 32'h3e3f7cac} /* (31, 1, 18) {real, imag} */,
  {32'hbdb376be, 32'h3e6bb03b} /* (31, 1, 17) {real, imag} */,
  {32'hbe156dda, 32'h3de8c794} /* (31, 1, 16) {real, imag} */,
  {32'h3d4e1af4, 32'h3eb59f0a} /* (31, 1, 15) {real, imag} */,
  {32'hbe93965f, 32'hbe9959cb} /* (31, 1, 14) {real, imag} */,
  {32'h3df54597, 32'h3f120d4f} /* (31, 1, 13) {real, imag} */,
  {32'h3e39e30e, 32'h3e54cb9f} /* (31, 1, 12) {real, imag} */,
  {32'hbebe7cb9, 32'h3d7c6964} /* (31, 1, 11) {real, imag} */,
  {32'hbe21aa6b, 32'hbd688044} /* (31, 1, 10) {real, imag} */,
  {32'h3e3efc4c, 32'hbeeeb4a8} /* (31, 1, 9) {real, imag} */,
  {32'h3e2eb782, 32'hbf5d0b00} /* (31, 1, 8) {real, imag} */,
  {32'h3db4c462, 32'h3f2033b4} /* (31, 1, 7) {real, imag} */,
  {32'hbe7abd28, 32'hbdd31204} /* (31, 1, 6) {real, imag} */,
  {32'hbf419ccd, 32'hbf1e7756} /* (31, 1, 5) {real, imag} */,
  {32'h3f919b1d, 32'hbf257278} /* (31, 1, 4) {real, imag} */,
  {32'h3eb62f1c, 32'h3f93848f} /* (31, 1, 3) {real, imag} */,
  {32'hc08daf0d, 32'hc0b2027c} /* (31, 1, 2) {real, imag} */,
  {32'h411dee52, 32'h40138702} /* (31, 1, 1) {real, imag} */,
  {32'h40a6c852, 32'h403b7234} /* (31, 1, 0) {real, imag} */,
  {32'h406591e2, 32'hc082af47} /* (31, 0, 31) {real, imag} */,
  {32'hc0139901, 32'h40735c40} /* (31, 0, 30) {real, imag} */,
  {32'hbdf28870, 32'h3f1941c4} /* (31, 0, 29) {real, imag} */,
  {32'hbf00970b, 32'h3e0278d0} /* (31, 0, 28) {real, imag} */,
  {32'h3da6e590, 32'hbd0108d8} /* (31, 0, 27) {real, imag} */,
  {32'hbefc997b, 32'h3db82b37} /* (31, 0, 26) {real, imag} */,
  {32'hbe905c1e, 32'hbf4942cd} /* (31, 0, 25) {real, imag} */,
  {32'h3dfe83b0, 32'h3d8c4b38} /* (31, 0, 24) {real, imag} */,
  {32'hbec60724, 32'h3e69cb32} /* (31, 0, 23) {real, imag} */,
  {32'h3e17e8f4, 32'hbead2e0a} /* (31, 0, 22) {real, imag} */,
  {32'hbf081b3d, 32'h3d94ba00} /* (31, 0, 21) {real, imag} */,
  {32'hbeaedbb8, 32'hbcf8b388} /* (31, 0, 20) {real, imag} */,
  {32'hbddcd052, 32'hbeb145fc} /* (31, 0, 19) {real, imag} */,
  {32'h3e7135b3, 32'h3da4c5c0} /* (31, 0, 18) {real, imag} */,
  {32'h3ccba7d8, 32'h3e649236} /* (31, 0, 17) {real, imag} */,
  {32'h3e4c8415, 32'h00000000} /* (31, 0, 16) {real, imag} */,
  {32'h3ccba7d8, 32'hbe649236} /* (31, 0, 15) {real, imag} */,
  {32'h3e7135b3, 32'hbda4c5c0} /* (31, 0, 14) {real, imag} */,
  {32'hbddcd052, 32'h3eb145fc} /* (31, 0, 13) {real, imag} */,
  {32'hbeaedbb8, 32'h3cf8b388} /* (31, 0, 12) {real, imag} */,
  {32'hbf081b3d, 32'hbd94ba00} /* (31, 0, 11) {real, imag} */,
  {32'h3e17e8f4, 32'h3ead2e0a} /* (31, 0, 10) {real, imag} */,
  {32'hbec60724, 32'hbe69cb32} /* (31, 0, 9) {real, imag} */,
  {32'h3dfe83b0, 32'hbd8c4b38} /* (31, 0, 8) {real, imag} */,
  {32'hbe905c1e, 32'h3f4942cd} /* (31, 0, 7) {real, imag} */,
  {32'hbefc997b, 32'hbdb82b37} /* (31, 0, 6) {real, imag} */,
  {32'h3da6e590, 32'h3d0108d8} /* (31, 0, 5) {real, imag} */,
  {32'hbf00970b, 32'hbe0278d0} /* (31, 0, 4) {real, imag} */,
  {32'hbdf28870, 32'hbf1941c4} /* (31, 0, 3) {real, imag} */,
  {32'hc0139901, 32'hc0735c40} /* (31, 0, 2) {real, imag} */,
  {32'h406591e2, 32'h4082af47} /* (31, 0, 1) {real, imag} */,
  {32'h3d282280, 32'h00000000} /* (31, 0, 0) {real, imag} */,
  {32'h41c21f17, 32'hc1227cc4} /* (30, 31, 31) {real, imag} */,
  {32'hc11e4521, 32'h4130ccd0} /* (30, 31, 30) {real, imag} */,
  {32'hbf5471d1, 32'hbfe25256} /* (30, 31, 29) {real, imag} */,
  {32'h3f99e16e, 32'hbdc17f90} /* (30, 31, 28) {real, imag} */,
  {32'hc038d91a, 32'h3f93a988} /* (30, 31, 27) {real, imag} */,
  {32'hbf32c782, 32'hbf359bb4} /* (30, 31, 26) {real, imag} */,
  {32'hbef184f2, 32'hbf13b1cb} /* (30, 31, 25) {real, imag} */,
  {32'h3d063858, 32'h3fd27a4a} /* (30, 31, 24) {real, imag} */,
  {32'h3f18db4c, 32'hbeb9a8f2} /* (30, 31, 23) {real, imag} */,
  {32'hbebf4064, 32'hbdfe9342} /* (30, 31, 22) {real, imag} */,
  {32'hbcb25a50, 32'h3ea9db26} /* (30, 31, 21) {real, imag} */,
  {32'h3ef9c11e, 32'h3e1b6199} /* (30, 31, 20) {real, imag} */,
  {32'h3e0fc74a, 32'hbf15c9ad} /* (30, 31, 19) {real, imag} */,
  {32'hbdf9a088, 32'h3e66a9ed} /* (30, 31, 18) {real, imag} */,
  {32'hbed89c5c, 32'h3d08bd24} /* (30, 31, 17) {real, imag} */,
  {32'h3d6a57ea, 32'hbc116758} /* (30, 31, 16) {real, imag} */,
  {32'h3de3144b, 32'h3e25d5b4} /* (30, 31, 15) {real, imag} */,
  {32'hbec54006, 32'hbf0c791b} /* (30, 31, 14) {real, imag} */,
  {32'h3e24a62a, 32'hbda07b78} /* (30, 31, 13) {real, imag} */,
  {32'h3eaf6794, 32'hbc9b6f90} /* (30, 31, 12) {real, imag} */,
  {32'hbe77277c, 32'hbf95520f} /* (30, 31, 11) {real, imag} */,
  {32'h3ea65ee8, 32'h3ed41d05} /* (30, 31, 10) {real, imag} */,
  {32'hbee073d7, 32'h3d66efc4} /* (30, 31, 9) {real, imag} */,
  {32'hbea44c3c, 32'hbf8901d8} /* (30, 31, 8) {real, imag} */,
  {32'h3f016a50, 32'h3f875831} /* (30, 31, 7) {real, imag} */,
  {32'hbf096380, 32'h3f193bbc} /* (30, 31, 6) {real, imag} */,
  {32'hc01085d0, 32'h3dd918e3} /* (30, 31, 5) {real, imag} */,
  {32'h3fd8ebff, 32'hbeda0434} /* (30, 31, 4) {real, imag} */,
  {32'hbf3856be, 32'hbd8f5720} /* (30, 31, 3) {real, imag} */,
  {32'hc0e8e09c, 32'hbf46c33f} /* (30, 31, 2) {real, imag} */,
  {32'h418cc7f4, 32'h409c48f1} /* (30, 31, 1) {real, imag} */,
  {32'h416a7508, 32'hc05c2030} /* (30, 31, 0) {real, imag} */,
  {32'hc14c7bde, 32'hc094ae16} /* (30, 30, 31) {real, imag} */,
  {32'h40e04551, 32'h3f27d804} /* (30, 30, 30) {real, imag} */,
  {32'hbf93b24c, 32'h3f9ef420} /* (30, 30, 29) {real, imag} */,
  {32'hbfca1882, 32'hbe81c8f0} /* (30, 30, 28) {real, imag} */,
  {32'h3fcc8b2c, 32'hbec4d83c} /* (30, 30, 27) {real, imag} */,
  {32'h3db3ab24, 32'hbeca03fe} /* (30, 30, 26) {real, imag} */,
  {32'h3e613ed8, 32'h3f2ea44b} /* (30, 30, 25) {real, imag} */,
  {32'h3e94623a, 32'hbdcc80cc} /* (30, 30, 24) {real, imag} */,
  {32'h3f10a162, 32'hbd80af9b} /* (30, 30, 23) {real, imag} */,
  {32'h3a81ad00, 32'h3ea88ab8} /* (30, 30, 22) {real, imag} */,
  {32'h3f5159aa, 32'hbf8343f8} /* (30, 30, 21) {real, imag} */,
  {32'h3c95ef50, 32'h3ec91cc6} /* (30, 30, 20) {real, imag} */,
  {32'hbea96c5a, 32'h3cb6d1be} /* (30, 30, 19) {real, imag} */,
  {32'hbc7f0570, 32'h3d11b640} /* (30, 30, 18) {real, imag} */,
  {32'hbe8ddf8d, 32'hbda48edc} /* (30, 30, 17) {real, imag} */,
  {32'h3daf37a3, 32'hbdf8583c} /* (30, 30, 16) {real, imag} */,
  {32'h3e9e51fd, 32'h3e6ce93b} /* (30, 30, 15) {real, imag} */,
  {32'hbe11d9f6, 32'h3efa90a0} /* (30, 30, 14) {real, imag} */,
  {32'hbd9dc810, 32'h3e2fe492} /* (30, 30, 13) {real, imag} */,
  {32'hbdcd99d1, 32'hbef07dc8} /* (30, 30, 12) {real, imag} */,
  {32'hbe2974d3, 32'h3ef3507e} /* (30, 30, 11) {real, imag} */,
  {32'hbea5b02e, 32'hbe0b10c2} /* (30, 30, 10) {real, imag} */,
  {32'h3cca5ee0, 32'hbe4d3253} /* (30, 30, 9) {real, imag} */,
  {32'h3fae19b9, 32'h3ea64456} /* (30, 30, 8) {real, imag} */,
  {32'hbeb5bba6, 32'h3e6836ca} /* (30, 30, 7) {real, imag} */,
  {32'h3f0ee529, 32'hbe8e4f4a} /* (30, 30, 6) {real, imag} */,
  {32'h3fb6c4f6, 32'h3e9f778e} /* (30, 30, 5) {real, imag} */,
  {32'hbfcc6cd7, 32'hc035afd4} /* (30, 30, 4) {real, imag} */,
  {32'h3f971962, 32'hbdbe4ad4} /* (30, 30, 3) {real, imag} */,
  {32'h411c9632, 32'h4072ba10} /* (30, 30, 2) {real, imag} */,
  {32'hc19425c8, 32'h400b522d} /* (30, 30, 1) {real, imag} */,
  {32'hc126596a, 32'h3f816126} /* (30, 30, 0) {real, imag} */,
  {32'h3fe21b78, 32'hbfdd548c} /* (30, 29, 31) {real, imag} */,
  {32'hbe539334, 32'h400bb6a3} /* (30, 29, 30) {real, imag} */,
  {32'h3f54574d, 32'hbdc10af0} /* (30, 29, 29) {real, imag} */,
  {32'hbe68d1cc, 32'hbf15f5e1} /* (30, 29, 28) {real, imag} */,
  {32'hbf5df5c5, 32'hbf0f1870} /* (30, 29, 27) {real, imag} */,
  {32'hbcfa5d40, 32'hbe18577e} /* (30, 29, 26) {real, imag} */,
  {32'h3f3d5a26, 32'hbe85a390} /* (30, 29, 25) {real, imag} */,
  {32'hbde25cf7, 32'h3e2beb4c} /* (30, 29, 24) {real, imag} */,
  {32'h3e15c2aa, 32'hbe47d443} /* (30, 29, 23) {real, imag} */,
  {32'hbf11b68a, 32'h3efe70c3} /* (30, 29, 22) {real, imag} */,
  {32'hbe964c3f, 32'hbec198a1} /* (30, 29, 21) {real, imag} */,
  {32'hbe22c39c, 32'h3e608925} /* (30, 29, 20) {real, imag} */,
  {32'h3ecd5ac8, 32'hbe9b256e} /* (30, 29, 19) {real, imag} */,
  {32'hbd04a0f0, 32'h3d325bc0} /* (30, 29, 18) {real, imag} */,
  {32'h3da5959d, 32'hbdeb5d44} /* (30, 29, 17) {real, imag} */,
  {32'hbad1b640, 32'h3effa722} /* (30, 29, 16) {real, imag} */,
  {32'h3e320d94, 32'h3e1062ce} /* (30, 29, 15) {real, imag} */,
  {32'h3d7a41db, 32'hbd30baf8} /* (30, 29, 14) {real, imag} */,
  {32'hbe2dddc2, 32'hbe66501a} /* (30, 29, 13) {real, imag} */,
  {32'hbefad778, 32'hbd9371e4} /* (30, 29, 12) {real, imag} */,
  {32'hbecdbfc9, 32'hbe0d0915} /* (30, 29, 11) {real, imag} */,
  {32'hb9fcf580, 32'hbeac0f0b} /* (30, 29, 10) {real, imag} */,
  {32'h3cdd1d40, 32'hbdc0569c} /* (30, 29, 9) {real, imag} */,
  {32'hbe9da3a4, 32'h3c6de760} /* (30, 29, 8) {real, imag} */,
  {32'hbe9fd18d, 32'hbe977b6e} /* (30, 29, 7) {real, imag} */,
  {32'h3dacf338, 32'h3e1d30f0} /* (30, 29, 6) {real, imag} */,
  {32'h3e3148a3, 32'h3f1bf8b4} /* (30, 29, 5) {real, imag} */,
  {32'h3dadb324, 32'hbf2cd2ee} /* (30, 29, 4) {real, imag} */,
  {32'h3eb8d2b4, 32'hbeb8d840} /* (30, 29, 3) {real, imag} */,
  {32'h3fe322f8, 32'h401a2415} /* (30, 29, 2) {real, imag} */,
  {32'hc036eec5, 32'hc01606d2} /* (30, 29, 1) {real, imag} */,
  {32'hbebfa95e, 32'hbf17dbf8} /* (30, 29, 0) {real, imag} */,
  {32'h4080b95a, 32'hc00a6147} /* (30, 28, 31) {real, imag} */,
  {32'hbfa12f4a, 32'h40118674} /* (30, 28, 30) {real, imag} */,
  {32'h3e43c42e, 32'hbf06919d} /* (30, 28, 29) {real, imag} */,
  {32'hbd8600f4, 32'hbf6cb9e9} /* (30, 28, 28) {real, imag} */,
  {32'h3efdf056, 32'h3f58f569} /* (30, 28, 27) {real, imag} */,
  {32'hbc4a2cf0, 32'h3e8da080} /* (30, 28, 26) {real, imag} */,
  {32'h3f279a69, 32'hbf604ac4} /* (30, 28, 25) {real, imag} */,
  {32'hbd11c210, 32'hbe7111a4} /* (30, 28, 24) {real, imag} */,
  {32'h3f1798d1, 32'h3cf54592} /* (30, 28, 23) {real, imag} */,
  {32'hbf1261bf, 32'hbf450aba} /* (30, 28, 22) {real, imag} */,
  {32'h3eb51043, 32'h3e70734c} /* (30, 28, 21) {real, imag} */,
  {32'hbbf523d0, 32'h3eb2ec21} /* (30, 28, 20) {real, imag} */,
  {32'h3e843fae, 32'h3e01e9d0} /* (30, 28, 19) {real, imag} */,
  {32'hbdecddf0, 32'h3daf1f6c} /* (30, 28, 18) {real, imag} */,
  {32'h3df835ca, 32'h3cf7d3c0} /* (30, 28, 17) {real, imag} */,
  {32'hbeaf5a5c, 32'h3cd0cb5e} /* (30, 28, 16) {real, imag} */,
  {32'h3e24b966, 32'h3da3b0fc} /* (30, 28, 15) {real, imag} */,
  {32'h3dbb39a8, 32'hbea7093e} /* (30, 28, 14) {real, imag} */,
  {32'h3df3f710, 32'hbddb3409} /* (30, 28, 13) {real, imag} */,
  {32'h3dd2ee7b, 32'h3eaa1db6} /* (30, 28, 12) {real, imag} */,
  {32'hbf0f906e, 32'hbe91c2d4} /* (30, 28, 11) {real, imag} */,
  {32'h3efcc0b4, 32'h3d8e9a2c} /* (30, 28, 10) {real, imag} */,
  {32'h3eb88d6a, 32'hbe2ed6cc} /* (30, 28, 9) {real, imag} */,
  {32'hbd947ad1, 32'h3dc0b6f4} /* (30, 28, 8) {real, imag} */,
  {32'hbee70735, 32'h3e055dcf} /* (30, 28, 7) {real, imag} */,
  {32'hbb556980, 32'hbc6bd640} /* (30, 28, 6) {real, imag} */,
  {32'hbf731231, 32'h3ecc2f3e} /* (30, 28, 5) {real, imag} */,
  {32'h3f8456f6, 32'hbf3fa27a} /* (30, 28, 4) {real, imag} */,
  {32'hbe743d2a, 32'hbf6aa4fc} /* (30, 28, 3) {real, imag} */,
  {32'hc03e70cc, 32'h3de8fcf0} /* (30, 28, 2) {real, imag} */,
  {32'h3fe08b95, 32'hc0020672} /* (30, 28, 1) {real, imag} */,
  {32'h4008bf4e, 32'hbf29079d} /* (30, 28, 0) {real, imag} */,
  {32'hbfe85825, 32'h4004576e} /* (30, 27, 31) {real, imag} */,
  {32'h3fc840ea, 32'hbf997758} /* (30, 27, 30) {real, imag} */,
  {32'hbe07ca4c, 32'h3b714fc0} /* (30, 27, 29) {real, imag} */,
  {32'hbf1401c5, 32'h3f1075ac} /* (30, 27, 28) {real, imag} */,
  {32'hbeeecd65, 32'hbf0397dc} /* (30, 27, 27) {real, imag} */,
  {32'h3f08efa0, 32'h3d5322ec} /* (30, 27, 26) {real, imag} */,
  {32'h3ed540df, 32'h3ef60a79} /* (30, 27, 25) {real, imag} */,
  {32'hbe9cf8d5, 32'hbedde052} /* (30, 27, 24) {real, imag} */,
  {32'h3e04106e, 32'hbf056184} /* (30, 27, 23) {real, imag} */,
  {32'hbd581dea, 32'hbdf22fb6} /* (30, 27, 22) {real, imag} */,
  {32'hbf29fc6d, 32'hbdac69c4} /* (30, 27, 21) {real, imag} */,
  {32'hbdbc5990, 32'hbef987d1} /* (30, 27, 20) {real, imag} */,
  {32'h3e7a1402, 32'hbc44d0c0} /* (30, 27, 19) {real, imag} */,
  {32'h3d4183de, 32'hbe6235ca} /* (30, 27, 18) {real, imag} */,
  {32'hbe1e57c3, 32'hbd45a6f4} /* (30, 27, 17) {real, imag} */,
  {32'hbdc4c6d9, 32'hbdd97a15} /* (30, 27, 16) {real, imag} */,
  {32'hbe020c95, 32'h3d5b1ac2} /* (30, 27, 15) {real, imag} */,
  {32'hbe87ba82, 32'h3cb7e630} /* (30, 27, 14) {real, imag} */,
  {32'h3e124e91, 32'h3ddb4768} /* (30, 27, 13) {real, imag} */,
  {32'hbe1a1fad, 32'h3dfe8696} /* (30, 27, 12) {real, imag} */,
  {32'h3e39d914, 32'h3ce69868} /* (30, 27, 11) {real, imag} */,
  {32'h3d4e1470, 32'h3f686c70} /* (30, 27, 10) {real, imag} */,
  {32'hbed13b06, 32'h3e88c0c7} /* (30, 27, 9) {real, imag} */,
  {32'hbda01f6e, 32'hbf0ab02e} /* (30, 27, 8) {real, imag} */,
  {32'hbf376f45, 32'hbeb0e778} /* (30, 27, 7) {real, imag} */,
  {32'hbe784284, 32'hbd9ea044} /* (30, 27, 6) {real, imag} */,
  {32'h3f55bf3b, 32'h3d8f45c6} /* (30, 27, 5) {real, imag} */,
  {32'h3ea4fc64, 32'hbed45c23} /* (30, 27, 4) {real, imag} */,
  {32'h3e12d792, 32'h3e128776} /* (30, 27, 3) {real, imag} */,
  {32'h3f382820, 32'h3f8b0019} /* (30, 27, 2) {real, imag} */,
  {32'hc01f0a5e, 32'h3ed0e478} /* (30, 27, 1) {real, imag} */,
  {32'hc011a4a3, 32'hbe6b5d26} /* (30, 27, 0) {real, imag} */,
  {32'hbf9b5ed5, 32'h3e92e702} /* (30, 26, 31) {real, imag} */,
  {32'h3db392c0, 32'h3ecb219a} /* (30, 26, 30) {real, imag} */,
  {32'hbe9d94b9, 32'hbe84dd62} /* (30, 26, 29) {real, imag} */,
  {32'h3ed8ef52, 32'hbd02cc2c} /* (30, 26, 28) {real, imag} */,
  {32'h3f3200d6, 32'hbeae0121} /* (30, 26, 27) {real, imag} */,
  {32'hbf00f4e0, 32'hbee6e546} /* (30, 26, 26) {real, imag} */,
  {32'h3d93c534, 32'hbea3cba9} /* (30, 26, 25) {real, imag} */,
  {32'h3e10d4ec, 32'hbde4432c} /* (30, 26, 24) {real, imag} */,
  {32'hbeec06c4, 32'hbe88b9da} /* (30, 26, 23) {real, imag} */,
  {32'h3df23bd8, 32'h3f08211b} /* (30, 26, 22) {real, imag} */,
  {32'h3db62000, 32'h3e5e3954} /* (30, 26, 21) {real, imag} */,
  {32'hbed475ce, 32'h3e3759a2} /* (30, 26, 20) {real, imag} */,
  {32'h3e09b9b2, 32'hbe52a89b} /* (30, 26, 19) {real, imag} */,
  {32'h3dbd65c1, 32'hbe1ffa9c} /* (30, 26, 18) {real, imag} */,
  {32'hbe4f65f8, 32'hbe065fbc} /* (30, 26, 17) {real, imag} */,
  {32'h3e806c63, 32'h3e4b91b6} /* (30, 26, 16) {real, imag} */,
  {32'hbd8535b6, 32'h3ea8c4b4} /* (30, 26, 15) {real, imag} */,
  {32'h3f013200, 32'hbead4bfe} /* (30, 26, 14) {real, imag} */,
  {32'hbf24ee8c, 32'h3eeaadce} /* (30, 26, 13) {real, imag} */,
  {32'hbf02fe59, 32'hbe4346d2} /* (30, 26, 12) {real, imag} */,
  {32'hbe960f55, 32'hbd7131b8} /* (30, 26, 11) {real, imag} */,
  {32'h3de41684, 32'h3d66d9a0} /* (30, 26, 10) {real, imag} */,
  {32'hbd0a9284, 32'h3e0fc940} /* (30, 26, 9) {real, imag} */,
  {32'h3f0ad94a, 32'h3ee9030b} /* (30, 26, 8) {real, imag} */,
  {32'h3d0cef84, 32'h3d259848} /* (30, 26, 7) {real, imag} */,
  {32'h3eb1d327, 32'hbf2e08e8} /* (30, 26, 6) {real, imag} */,
  {32'h3d3770f2, 32'hbe8c30b1} /* (30, 26, 5) {real, imag} */,
  {32'hbd580430, 32'h3d6085c0} /* (30, 26, 4) {real, imag} */,
  {32'h3ddb73e8, 32'h3f28213e} /* (30, 26, 3) {real, imag} */,
  {32'hbf1e0e33, 32'hbe33dfed} /* (30, 26, 2) {real, imag} */,
  {32'hbf287fe7, 32'hbf97ef32} /* (30, 26, 1) {real, imag} */,
  {32'h3f3b76e3, 32'hbdc5bf5b} /* (30, 26, 0) {real, imag} */,
  {32'hbe3d6db2, 32'hbeeef9e3} /* (30, 25, 31) {real, imag} */,
  {32'h3f1e2ee1, 32'h3ef9c2d0} /* (30, 25, 30) {real, imag} */,
  {32'h3e050b90, 32'h3e92043d} /* (30, 25, 29) {real, imag} */,
  {32'h3dd01f4c, 32'hbdbcfb98} /* (30, 25, 28) {real, imag} */,
  {32'h3ed786f6, 32'hbe9063f8} /* (30, 25, 27) {real, imag} */,
  {32'h3e043dea, 32'h3e464d82} /* (30, 25, 26) {real, imag} */,
  {32'h3db1f4d7, 32'h3e15bfd4} /* (30, 25, 25) {real, imag} */,
  {32'h3eb1bb08, 32'hbd92e5c4} /* (30, 25, 24) {real, imag} */,
  {32'h3d8fd6ac, 32'h3d67c2e8} /* (30, 25, 23) {real, imag} */,
  {32'h3ead0b25, 32'hbe95a868} /* (30, 25, 22) {real, imag} */,
  {32'h3dc641d6, 32'hbd91d657} /* (30, 25, 21) {real, imag} */,
  {32'h3dcc8518, 32'h3dd75962} /* (30, 25, 20) {real, imag} */,
  {32'h3e9ceef9, 32'h3d726084} /* (30, 25, 19) {real, imag} */,
  {32'hbe9ff05d, 32'hbd478734} /* (30, 25, 18) {real, imag} */,
  {32'hbdfa5d28, 32'h3dd66ab7} /* (30, 25, 17) {real, imag} */,
  {32'h3eb1ac6d, 32'h3d56d25a} /* (30, 25, 16) {real, imag} */,
  {32'hbe9caaf4, 32'hbca28cfc} /* (30, 25, 15) {real, imag} */,
  {32'h3df5cd34, 32'hbd7a7830} /* (30, 25, 14) {real, imag} */,
  {32'h3e3cceba, 32'h3e83d585} /* (30, 25, 13) {real, imag} */,
  {32'hbef1bda8, 32'hbd4918b8} /* (30, 25, 12) {real, imag} */,
  {32'h3ee23703, 32'hbdb635cb} /* (30, 25, 11) {real, imag} */,
  {32'hbe09818a, 32'h3e0bd4d5} /* (30, 25, 10) {real, imag} */,
  {32'h3e9dc2e9, 32'hbeabfa4d} /* (30, 25, 9) {real, imag} */,
  {32'hbddc959c, 32'hbcd6a23c} /* (30, 25, 8) {real, imag} */,
  {32'hbf0697da, 32'h3d739020} /* (30, 25, 7) {real, imag} */,
  {32'h3ec798e6, 32'hbf2581d0} /* (30, 25, 6) {real, imag} */,
  {32'hbec4aa52, 32'h3ea34d83} /* (30, 25, 5) {real, imag} */,
  {32'hbf444bba, 32'h3c1fae30} /* (30, 25, 4) {real, imag} */,
  {32'h3e6e91b0, 32'hbea55a68} /* (30, 25, 3) {real, imag} */,
  {32'hbf0689a4, 32'h3eea6674} /* (30, 25, 2) {real, imag} */,
  {32'h3e51cba9, 32'hbeb5a8d2} /* (30, 25, 1) {real, imag} */,
  {32'h3f46a4ad, 32'hbe35171e} /* (30, 25, 0) {real, imag} */,
  {32'hbf332438, 32'h3f6df06f} /* (30, 24, 31) {real, imag} */,
  {32'h3f1b5584, 32'hbfa504e6} /* (30, 24, 30) {real, imag} */,
  {32'hbeb001c4, 32'hbef02912} /* (30, 24, 29) {real, imag} */,
  {32'hbf1471d2, 32'hbe878619} /* (30, 24, 28) {real, imag} */,
  {32'h3eac15fa, 32'hbe007bad} /* (30, 24, 27) {real, imag} */,
  {32'h3da52170, 32'hbea6649a} /* (30, 24, 26) {real, imag} */,
  {32'hbe795c26, 32'hbede36ea} /* (30, 24, 25) {real, imag} */,
  {32'hbe84fe0f, 32'h3d7b56b6} /* (30, 24, 24) {real, imag} */,
  {32'hbe965bf5, 32'h3ecaefe6} /* (30, 24, 23) {real, imag} */,
  {32'h3dc26b7e, 32'hbf0358a9} /* (30, 24, 22) {real, imag} */,
  {32'hbca0c910, 32'hbdce748c} /* (30, 24, 21) {real, imag} */,
  {32'hbee3c9f2, 32'hbe0388ee} /* (30, 24, 20) {real, imag} */,
  {32'hbd937ce0, 32'h3e8a1193} /* (30, 24, 19) {real, imag} */,
  {32'hbd8e7770, 32'h3f01f9c7} /* (30, 24, 18) {real, imag} */,
  {32'hbe7ce68a, 32'h3d7bb210} /* (30, 24, 17) {real, imag} */,
  {32'hbeb82322, 32'hbe170fcc} /* (30, 24, 16) {real, imag} */,
  {32'h3f0c39fe, 32'hbddd06e5} /* (30, 24, 15) {real, imag} */,
  {32'hbd6e6366, 32'hbe6dcf2f} /* (30, 24, 14) {real, imag} */,
  {32'h3ea380d8, 32'hbd2f3668} /* (30, 24, 13) {real, imag} */,
  {32'h3de492b8, 32'h3e2bb85a} /* (30, 24, 12) {real, imag} */,
  {32'h3dba114e, 32'h3ecb43ca} /* (30, 24, 11) {real, imag} */,
  {32'h3dfc39da, 32'h3eba9878} /* (30, 24, 10) {real, imag} */,
  {32'hbe084798, 32'hbdb48eb0} /* (30, 24, 9) {real, imag} */,
  {32'h3e0cefeb, 32'h3dac7548} /* (30, 24, 8) {real, imag} */,
  {32'h3d8a2bb4, 32'h3ece5c8b} /* (30, 24, 7) {real, imag} */,
  {32'h3d9f7754, 32'hbe9d7536} /* (30, 24, 6) {real, imag} */,
  {32'hbe1ae594, 32'hbe7f5602} /* (30, 24, 5) {real, imag} */,
  {32'hbd958e38, 32'hbed515d3} /* (30, 24, 4) {real, imag} */,
  {32'hbebf5af0, 32'h3f187ff3} /* (30, 24, 3) {real, imag} */,
  {32'h3f90b064, 32'hbc2c1720} /* (30, 24, 2) {real, imag} */,
  {32'hbf8c8f3f, 32'h3f322d7c} /* (30, 24, 1) {real, imag} */,
  {32'hbf9f2882, 32'hbd6d2c20} /* (30, 24, 0) {real, imag} */,
  {32'h3f545051, 32'hbe1e398e} /* (30, 23, 31) {real, imag} */,
  {32'hbf7117be, 32'h3f42bc3e} /* (30, 23, 30) {real, imag} */,
  {32'hbf437583, 32'h3ecabf67} /* (30, 23, 29) {real, imag} */,
  {32'h3df4c8e1, 32'hbebd72f0} /* (30, 23, 28) {real, imag} */,
  {32'h3e45e35f, 32'hbf01f461} /* (30, 23, 27) {real, imag} */,
  {32'hbd4e00d2, 32'h3de30438} /* (30, 23, 26) {real, imag} */,
  {32'h3e5e55f9, 32'h3f0ce627} /* (30, 23, 25) {real, imag} */,
  {32'hbd8fb214, 32'hbe03d40c} /* (30, 23, 24) {real, imag} */,
  {32'h3eaf055c, 32'hbd958a74} /* (30, 23, 23) {real, imag} */,
  {32'hbe2a0f40, 32'h3e9abc9b} /* (30, 23, 22) {real, imag} */,
  {32'hbe677c3a, 32'hbcf765c0} /* (30, 23, 21) {real, imag} */,
  {32'h3e727e2a, 32'h3f07b336} /* (30, 23, 20) {real, imag} */,
  {32'hbe83398a, 32'h3ce5778c} /* (30, 23, 19) {real, imag} */,
  {32'hbef8098c, 32'hbea64943} /* (30, 23, 18) {real, imag} */,
  {32'hbe03cfec, 32'hbd510ef0} /* (30, 23, 17) {real, imag} */,
  {32'h3e3c6a7a, 32'h3c04cc40} /* (30, 23, 16) {real, imag} */,
  {32'h3dc1f254, 32'hbcba6898} /* (30, 23, 15) {real, imag} */,
  {32'h3e373258, 32'h3f0cbd82} /* (30, 23, 14) {real, imag} */,
  {32'hbe997830, 32'h3de0e2ab} /* (30, 23, 13) {real, imag} */,
  {32'h3f07d16d, 32'h3e9eea4b} /* (30, 23, 12) {real, imag} */,
  {32'h3e84c942, 32'hbebee5ad} /* (30, 23, 11) {real, imag} */,
  {32'h3e259cd6, 32'hbea737c6} /* (30, 23, 10) {real, imag} */,
  {32'hbdd75508, 32'h3e7ba745} /* (30, 23, 9) {real, imag} */,
  {32'hbef965c9, 32'h3f3694d7} /* (30, 23, 8) {real, imag} */,
  {32'h3df8e610, 32'h3e984bdd} /* (30, 23, 7) {real, imag} */,
  {32'h3eb1e7da, 32'hbe94b30d} /* (30, 23, 6) {real, imag} */,
  {32'hbede196a, 32'h3ed292ae} /* (30, 23, 5) {real, imag} */,
  {32'hbd75d16e, 32'hbe52beca} /* (30, 23, 4) {real, imag} */,
  {32'hbf0f4920, 32'hbf31f972} /* (30, 23, 3) {real, imag} */,
  {32'h3e4232de, 32'h3dc39528} /* (30, 23, 2) {real, imag} */,
  {32'hbf0ed06e, 32'hbeb8c11c} /* (30, 23, 1) {real, imag} */,
  {32'h3dda2068, 32'hbe7c53fe} /* (30, 23, 0) {real, imag} */,
  {32'hbe95bedf, 32'hbd5a6bac} /* (30, 22, 31) {real, imag} */,
  {32'hbeeef0b4, 32'h3f127529} /* (30, 22, 30) {real, imag} */,
  {32'h3e1b1c70, 32'hbe86a8e6} /* (30, 22, 29) {real, imag} */,
  {32'hbe479b4a, 32'hb829a000} /* (30, 22, 28) {real, imag} */,
  {32'hbe88b1d6, 32'h3e80da76} /* (30, 22, 27) {real, imag} */,
  {32'hbdfea1aa, 32'h3f28ad98} /* (30, 22, 26) {real, imag} */,
  {32'h3eb9ce38, 32'hbedd0a30} /* (30, 22, 25) {real, imag} */,
  {32'h3e4f3be3, 32'h3ea20cc7} /* (30, 22, 24) {real, imag} */,
  {32'h3e874a44, 32'hbd547fa0} /* (30, 22, 23) {real, imag} */,
  {32'hbe66cd6b, 32'hbec84332} /* (30, 22, 22) {real, imag} */,
  {32'h3e0059c2, 32'hbe042ad2} /* (30, 22, 21) {real, imag} */,
  {32'hbf1ec2e5, 32'hbe3aa276} /* (30, 22, 20) {real, imag} */,
  {32'h3f71c158, 32'h3e957f1e} /* (30, 22, 19) {real, imag} */,
  {32'hbd82409c, 32'hbe04bffa} /* (30, 22, 18) {real, imag} */,
  {32'hbe07a3f2, 32'hbe8cb621} /* (30, 22, 17) {real, imag} */,
  {32'hbe60bd61, 32'hbcd47bb8} /* (30, 22, 16) {real, imag} */,
  {32'h3d331994, 32'hbdf661a1} /* (30, 22, 15) {real, imag} */,
  {32'h3e61b281, 32'h3ecb7c42} /* (30, 22, 14) {real, imag} */,
  {32'h3f360d69, 32'hbe1ea928} /* (30, 22, 13) {real, imag} */,
  {32'h3e40898e, 32'hbf21188e} /* (30, 22, 12) {real, imag} */,
  {32'hbf3b61aa, 32'h3d33b9c8} /* (30, 22, 11) {real, imag} */,
  {32'h3df562e6, 32'h3f3db0e8} /* (30, 22, 10) {real, imag} */,
  {32'hbe8af730, 32'h3de47bf4} /* (30, 22, 9) {real, imag} */,
  {32'hbeef821e, 32'h3e0b15bb} /* (30, 22, 8) {real, imag} */,
  {32'hbd9d5bce, 32'h3e872227} /* (30, 22, 7) {real, imag} */,
  {32'h3dde485a, 32'h3e16c279} /* (30, 22, 6) {real, imag} */,
  {32'h3e37f15a, 32'hbdd20ca5} /* (30, 22, 5) {real, imag} */,
  {32'h3e4bc290, 32'h3ebc59b2} /* (30, 22, 4) {real, imag} */,
  {32'h3e5fc0dd, 32'h3cf1c478} /* (30, 22, 3) {real, imag} */,
  {32'h3efe9c1b, 32'h3e8fdf20} /* (30, 22, 2) {real, imag} */,
  {32'hbc837ded, 32'hbf244a5a} /* (30, 22, 1) {real, imag} */,
  {32'hbd9c8662, 32'h3ec188d2} /* (30, 22, 0) {real, imag} */,
  {32'hbe286b2d, 32'h3eae839f} /* (30, 21, 31) {real, imag} */,
  {32'hbeb06b0b, 32'hbef655dd} /* (30, 21, 30) {real, imag} */,
  {32'h3ee6c75a, 32'h3e95b272} /* (30, 21, 29) {real, imag} */,
  {32'h3e0902ec, 32'h3e6d00c0} /* (30, 21, 28) {real, imag} */,
  {32'h3e15f5da, 32'hbcbe0370} /* (30, 21, 27) {real, imag} */,
  {32'hbe7b842a, 32'h3e030f5e} /* (30, 21, 26) {real, imag} */,
  {32'h3e94cd2e, 32'h3e22297d} /* (30, 21, 25) {real, imag} */,
  {32'hbda822ee, 32'h3e6f4c10} /* (30, 21, 24) {real, imag} */,
  {32'hbf065044, 32'hbe573561} /* (30, 21, 23) {real, imag} */,
  {32'h3ea996e6, 32'hbe14882b} /* (30, 21, 22) {real, imag} */,
  {32'h3e6e4c9c, 32'h3eaa0132} /* (30, 21, 21) {real, imag} */,
  {32'hbbfda970, 32'hbea2ba80} /* (30, 21, 20) {real, imag} */,
  {32'h3e174a51, 32'hbe0229ca} /* (30, 21, 19) {real, imag} */,
  {32'hbe8a1767, 32'hbc6da5a0} /* (30, 21, 18) {real, imag} */,
  {32'h3ea225ef, 32'h3e77a1cf} /* (30, 21, 17) {real, imag} */,
  {32'hbea1d6bd, 32'hbdde3d58} /* (30, 21, 16) {real, imag} */,
  {32'h3d32293a, 32'hbea0ddea} /* (30, 21, 15) {real, imag} */,
  {32'h3eb2d10a, 32'h3e3726ca} /* (30, 21, 14) {real, imag} */,
  {32'hbf05f5ac, 32'hbde96e77} /* (30, 21, 13) {real, imag} */,
  {32'h3edc7672, 32'hbe92ad82} /* (30, 21, 12) {real, imag} */,
  {32'h3eaabc1b, 32'hbe89efe8} /* (30, 21, 11) {real, imag} */,
  {32'hbf1c0043, 32'h3e3f8a0a} /* (30, 21, 10) {real, imag} */,
  {32'hbd0bba78, 32'h3ed8f721} /* (30, 21, 9) {real, imag} */,
  {32'hbdd17870, 32'hbecf13ea} /* (30, 21, 8) {real, imag} */,
  {32'hbd58f9c0, 32'h3c800590} /* (30, 21, 7) {real, imag} */,
  {32'hbec121f4, 32'hbed07525} /* (30, 21, 6) {real, imag} */,
  {32'hbdf6c9ca, 32'h3dd341f0} /* (30, 21, 5) {real, imag} */,
  {32'h3ec7f48e, 32'h3dee1e7c} /* (30, 21, 4) {real, imag} */,
  {32'h3e91fee8, 32'hbe807700} /* (30, 21, 3) {real, imag} */,
  {32'h3eef55f6, 32'hbef8a8f4} /* (30, 21, 2) {real, imag} */,
  {32'hbe00c062, 32'h3eda124a} /* (30, 21, 1) {real, imag} */,
  {32'hbde5903f, 32'h3f44ca47} /* (30, 21, 0) {real, imag} */,
  {32'h3e174fb8, 32'hbe7ff5ea} /* (30, 20, 31) {real, imag} */,
  {32'hbd0edd60, 32'h3d2b7942} /* (30, 20, 30) {real, imag} */,
  {32'h3ea6259e, 32'hbdf5d25e} /* (30, 20, 29) {real, imag} */,
  {32'h3c0a7468, 32'h3e22f9da} /* (30, 20, 28) {real, imag} */,
  {32'hbeb419bb, 32'h3e745c2b} /* (30, 20, 27) {real, imag} */,
  {32'h3f00dc04, 32'hbca81340} /* (30, 20, 26) {real, imag} */,
  {32'h38e09000, 32'hbe61ea44} /* (30, 20, 25) {real, imag} */,
  {32'hbe8e824e, 32'hbe63533d} /* (30, 20, 24) {real, imag} */,
  {32'hbe23d86e, 32'hbcb5e280} /* (30, 20, 23) {real, imag} */,
  {32'hbe883ca8, 32'h3c97b748} /* (30, 20, 22) {real, imag} */,
  {32'hbe91c2c6, 32'hbe9d05c4} /* (30, 20, 21) {real, imag} */,
  {32'h3ed9882a, 32'hbe122226} /* (30, 20, 20) {real, imag} */,
  {32'hbe8e083b, 32'hbc9470a0} /* (30, 20, 19) {real, imag} */,
  {32'hbd6756a8, 32'hbd8a09d8} /* (30, 20, 18) {real, imag} */,
  {32'h3de2f340, 32'hbde5f8f4} /* (30, 20, 17) {real, imag} */,
  {32'h3cf2f122, 32'hbe8aa61c} /* (30, 20, 16) {real, imag} */,
  {32'h3e9949e6, 32'hbeb9ea26} /* (30, 20, 15) {real, imag} */,
  {32'hbe96e3ec, 32'h3ec224ac} /* (30, 20, 14) {real, imag} */,
  {32'hbf0527cb, 32'h3ef3b049} /* (30, 20, 13) {real, imag} */,
  {32'hbed3098a, 32'h3cf88d78} /* (30, 20, 12) {real, imag} */,
  {32'h3eee7ce5, 32'hbdb9e252} /* (30, 20, 11) {real, imag} */,
  {32'h3ef2e13f, 32'hbe1bed08} /* (30, 20, 10) {real, imag} */,
  {32'hbc7258e8, 32'hbe5a4104} /* (30, 20, 9) {real, imag} */,
  {32'h3d539486, 32'h3e2d0cbe} /* (30, 20, 8) {real, imag} */,
  {32'hbe1df638, 32'hbc2424e0} /* (30, 20, 7) {real, imag} */,
  {32'h3d687a52, 32'h3f27dd56} /* (30, 20, 6) {real, imag} */,
  {32'hbe3879f2, 32'hbe7347be} /* (30, 20, 5) {real, imag} */,
  {32'hbe1e51a3, 32'hbe78a863} /* (30, 20, 4) {real, imag} */,
  {32'h3e83396c, 32'h3ed5d77a} /* (30, 20, 3) {real, imag} */,
  {32'hbd84b48c, 32'hbf0d2cd6} /* (30, 20, 2) {real, imag} */,
  {32'hbc18e780, 32'h3d4a38d0} /* (30, 20, 1) {real, imag} */,
  {32'hbd731310, 32'h3e808ecd} /* (30, 20, 0) {real, imag} */,
  {32'h3f1f5b05, 32'hbdc1d768} /* (30, 19, 31) {real, imag} */,
  {32'hbeb997fa, 32'h3d8ecb58} /* (30, 19, 30) {real, imag} */,
  {32'h3ea02240, 32'h3d4ee400} /* (30, 19, 29) {real, imag} */,
  {32'hbdb5ec2c, 32'h3f0124ab} /* (30, 19, 28) {real, imag} */,
  {32'hbed5d369, 32'hbecd0fc2} /* (30, 19, 27) {real, imag} */,
  {32'h3eea3900, 32'hbd2f1604} /* (30, 19, 26) {real, imag} */,
  {32'h3e0516c0, 32'hbefc4d68} /* (30, 19, 25) {real, imag} */,
  {32'hbeb30781, 32'hbc7d7ff0} /* (30, 19, 24) {real, imag} */,
  {32'hbe275752, 32'h3d124640} /* (30, 19, 23) {real, imag} */,
  {32'hbda2d9c8, 32'h3e6d85c4} /* (30, 19, 22) {real, imag} */,
  {32'hbe9393e8, 32'hbe975cd8} /* (30, 19, 21) {real, imag} */,
  {32'hbf0d1bd9, 32'hbda20d74} /* (30, 19, 20) {real, imag} */,
  {32'hbc41b110, 32'hbe2a2195} /* (30, 19, 19) {real, imag} */,
  {32'h3e855c05, 32'h3d9b5b10} /* (30, 19, 18) {real, imag} */,
  {32'h3ed5e640, 32'h3f10fc78} /* (30, 19, 17) {real, imag} */,
  {32'h3e7074f6, 32'h3c9f3a9e} /* (30, 19, 16) {real, imag} */,
  {32'hbedaf2d2, 32'h3e8300fe} /* (30, 19, 15) {real, imag} */,
  {32'hbf1cba2f, 32'h3c457a50} /* (30, 19, 14) {real, imag} */,
  {32'hbe98983d, 32'h3d9c37c0} /* (30, 19, 13) {real, imag} */,
  {32'hbdfd7d3d, 32'h3e3a843c} /* (30, 19, 12) {real, imag} */,
  {32'h3e1cdb3c, 32'h3e053084} /* (30, 19, 11) {real, imag} */,
  {32'h3e980f00, 32'h3cc5b310} /* (30, 19, 10) {real, imag} */,
  {32'hbd11fa60, 32'hbe07d1c2} /* (30, 19, 9) {real, imag} */,
  {32'hbca45f10, 32'hbe0f7e29} /* (30, 19, 8) {real, imag} */,
  {32'h3c3ed5e0, 32'hbe9aa37d} /* (30, 19, 7) {real, imag} */,
  {32'h3d8fd739, 32'h3f3d360d} /* (30, 19, 6) {real, imag} */,
  {32'hbea56ae2, 32'h3e2f55e4} /* (30, 19, 5) {real, imag} */,
  {32'h3e781470, 32'h3e146000} /* (30, 19, 4) {real, imag} */,
  {32'h3e209dc6, 32'h3def6e92} /* (30, 19, 3) {real, imag} */,
  {32'hbec9915e, 32'hbc93b010} /* (30, 19, 2) {real, imag} */,
  {32'hbe92dc48, 32'h3ea2d0d4} /* (30, 19, 1) {real, imag} */,
  {32'h3ded2d6f, 32'hbe34e4e6} /* (30, 19, 0) {real, imag} */,
  {32'hbc290890, 32'h3ec5f24a} /* (30, 18, 31) {real, imag} */,
  {32'hbd730368, 32'hbdb5d37e} /* (30, 18, 30) {real, imag} */,
  {32'hbd12ac84, 32'hbe45b661} /* (30, 18, 29) {real, imag} */,
  {32'hbefd7086, 32'h3f03fc4b} /* (30, 18, 28) {real, imag} */,
  {32'h3e87fc74, 32'hbd95fe68} /* (30, 18, 27) {real, imag} */,
  {32'h3f08589a, 32'hbe59d81e} /* (30, 18, 26) {real, imag} */,
  {32'h3e155823, 32'h3d8630e8} /* (30, 18, 25) {real, imag} */,
  {32'h3ef43b75, 32'hbe5e26dc} /* (30, 18, 24) {real, imag} */,
  {32'hbe35e323, 32'h3eae52a5} /* (30, 18, 23) {real, imag} */,
  {32'hbefee23c, 32'h3d40d8c5} /* (30, 18, 22) {real, imag} */,
  {32'hbcfdbfe0, 32'h3da8926c} /* (30, 18, 21) {real, imag} */,
  {32'hbe41b471, 32'h3d464d88} /* (30, 18, 20) {real, imag} */,
  {32'hbea19672, 32'h3e0ee620} /* (30, 18, 19) {real, imag} */,
  {32'h3ee2530a, 32'h3e0bf508} /* (30, 18, 18) {real, imag} */,
  {32'h3db8d8b5, 32'hbe304b3c} /* (30, 18, 17) {real, imag} */,
  {32'h3e7f8645, 32'h3e7e86b8} /* (30, 18, 16) {real, imag} */,
  {32'h3dbcad34, 32'h3dc08fb1} /* (30, 18, 15) {real, imag} */,
  {32'hbee271c9, 32'hbf06eee4} /* (30, 18, 14) {real, imag} */,
  {32'hbc454308, 32'hbf183775} /* (30, 18, 13) {real, imag} */,
  {32'hbe7eadc7, 32'h3e147ffa} /* (30, 18, 12) {real, imag} */,
  {32'hbd5960a5, 32'h3ddc0ab0} /* (30, 18, 11) {real, imag} */,
  {32'hbe6f2772, 32'hbdae0dee} /* (30, 18, 10) {real, imag} */,
  {32'hbe56e280, 32'hbd938d8c} /* (30, 18, 9) {real, imag} */,
  {32'h3f0c7b1b, 32'hbbdaddb0} /* (30, 18, 8) {real, imag} */,
  {32'h3e94ddde, 32'hbd07ef20} /* (30, 18, 7) {real, imag} */,
  {32'h3f091ebe, 32'h3e0c3e6d} /* (30, 18, 6) {real, imag} */,
  {32'h3b2b6fc0, 32'hbe5ddc99} /* (30, 18, 5) {real, imag} */,
  {32'hbd875a94, 32'h3da29434} /* (30, 18, 4) {real, imag} */,
  {32'h3ccc1550, 32'hbd9afcd6} /* (30, 18, 3) {real, imag} */,
  {32'h3dbdbca2, 32'hbd626840} /* (30, 18, 2) {real, imag} */,
  {32'h3c34dc6e, 32'h3f15ee2a} /* (30, 18, 1) {real, imag} */,
  {32'h3ec3c66e, 32'h3f0cb16e} /* (30, 18, 0) {real, imag} */,
  {32'h3c75d9e8, 32'hbe3e077b} /* (30, 17, 31) {real, imag} */,
  {32'hb9ad1c00, 32'h3edbc9cc} /* (30, 17, 30) {real, imag} */,
  {32'hbeb2531d, 32'h3d5c54fd} /* (30, 17, 29) {real, imag} */,
  {32'h3e922e44, 32'hbd5a470e} /* (30, 17, 28) {real, imag} */,
  {32'hbe3f6420, 32'hbe5b4af5} /* (30, 17, 27) {real, imag} */,
  {32'h3dc05ef0, 32'hbe19a0b0} /* (30, 17, 26) {real, imag} */,
  {32'hbe8ccc96, 32'h3e127e63} /* (30, 17, 25) {real, imag} */,
  {32'hbec6ef75, 32'hbeedb41a} /* (30, 17, 24) {real, imag} */,
  {32'h3d908484, 32'hbd4f85f6} /* (30, 17, 23) {real, imag} */,
  {32'hbd9d41be, 32'h3e8236cf} /* (30, 17, 22) {real, imag} */,
  {32'h3f240fa8, 32'hbe4c3151} /* (30, 17, 21) {real, imag} */,
  {32'h3e63ff33, 32'hbdc66fc9} /* (30, 17, 20) {real, imag} */,
  {32'hbd43c7b0, 32'h3e0ce660} /* (30, 17, 19) {real, imag} */,
  {32'hbe88d9e7, 32'h3d90f5da} /* (30, 17, 18) {real, imag} */,
  {32'h3daa6ccf, 32'h3db6414a} /* (30, 17, 17) {real, imag} */,
  {32'h3e730b59, 32'h3e4a2682} /* (30, 17, 16) {real, imag} */,
  {32'hbd3c9c93, 32'hbe48a377} /* (30, 17, 15) {real, imag} */,
  {32'h3d135bfa, 32'hbdf79ed0} /* (30, 17, 14) {real, imag} */,
  {32'hbeeb7a1c, 32'h3e2ca59c} /* (30, 17, 13) {real, imag} */,
  {32'h3e69525c, 32'h3e40ca8b} /* (30, 17, 12) {real, imag} */,
  {32'hbde71c92, 32'hbe0017d3} /* (30, 17, 11) {real, imag} */,
  {32'h3df92392, 32'hbe99945e} /* (30, 17, 10) {real, imag} */,
  {32'hbcdcac5c, 32'h3c3a2900} /* (30, 17, 9) {real, imag} */,
  {32'h3e902d09, 32'h3df1bdab} /* (30, 17, 8) {real, imag} */,
  {32'hbdd9c5ae, 32'hbea2ab8c} /* (30, 17, 7) {real, imag} */,
  {32'h3e8b9547, 32'hbd0c4bfa} /* (30, 17, 6) {real, imag} */,
  {32'h3df8cdac, 32'h3d29b848} /* (30, 17, 5) {real, imag} */,
  {32'h3d28eb47, 32'hbe3d9e08} /* (30, 17, 4) {real, imag} */,
  {32'h3dbb9036, 32'hbdd3a2a5} /* (30, 17, 3) {real, imag} */,
  {32'h3d9b0bc8, 32'h3f307e06} /* (30, 17, 2) {real, imag} */,
  {32'hbd5137f0, 32'hbe1cd7f2} /* (30, 17, 1) {real, imag} */,
  {32'h3c89f38c, 32'h3e55801a} /* (30, 17, 0) {real, imag} */,
  {32'h3e055a50, 32'hbdd820f9} /* (30, 16, 31) {real, imag} */,
  {32'hbded626a, 32'h3d978731} /* (30, 16, 30) {real, imag} */,
  {32'hbd98b504, 32'hbe721dd4} /* (30, 16, 29) {real, imag} */,
  {32'hbd14f03c, 32'hbe72a4c2} /* (30, 16, 28) {real, imag} */,
  {32'hbde7764c, 32'hbc62a50c} /* (30, 16, 27) {real, imag} */,
  {32'h3d5310e4, 32'h3eac6029} /* (30, 16, 26) {real, imag} */,
  {32'hbe82bbac, 32'h3c26c600} /* (30, 16, 25) {real, imag} */,
  {32'h3e103a62, 32'h3d1cd470} /* (30, 16, 24) {real, imag} */,
  {32'hbcbec850, 32'h3e020317} /* (30, 16, 23) {real, imag} */,
  {32'h3ed4fde2, 32'hbe88832a} /* (30, 16, 22) {real, imag} */,
  {32'h3e72aa30, 32'h3e1a1ede} /* (30, 16, 21) {real, imag} */,
  {32'h3e256bb6, 32'h3e8877d8} /* (30, 16, 20) {real, imag} */,
  {32'hbe936893, 32'h3f08f6b7} /* (30, 16, 19) {real, imag} */,
  {32'hbdae362e, 32'h3e1d9e36} /* (30, 16, 18) {real, imag} */,
  {32'hbe414c16, 32'hbe302e4e} /* (30, 16, 17) {real, imag} */,
  {32'hbd7ce92c, 32'h00000000} /* (30, 16, 16) {real, imag} */,
  {32'hbe414c16, 32'h3e302e4e} /* (30, 16, 15) {real, imag} */,
  {32'hbdae362e, 32'hbe1d9e36} /* (30, 16, 14) {real, imag} */,
  {32'hbe936893, 32'hbf08f6b7} /* (30, 16, 13) {real, imag} */,
  {32'h3e256bb6, 32'hbe8877d8} /* (30, 16, 12) {real, imag} */,
  {32'h3e72aa30, 32'hbe1a1ede} /* (30, 16, 11) {real, imag} */,
  {32'h3ed4fde2, 32'h3e88832a} /* (30, 16, 10) {real, imag} */,
  {32'hbcbec850, 32'hbe020317} /* (30, 16, 9) {real, imag} */,
  {32'h3e103a62, 32'hbd1cd470} /* (30, 16, 8) {real, imag} */,
  {32'hbe82bbac, 32'hbc26c600} /* (30, 16, 7) {real, imag} */,
  {32'h3d5310e4, 32'hbeac6029} /* (30, 16, 6) {real, imag} */,
  {32'hbde7764c, 32'h3c62a50c} /* (30, 16, 5) {real, imag} */,
  {32'hbd14f03c, 32'h3e72a4c2} /* (30, 16, 4) {real, imag} */,
  {32'hbd98b504, 32'h3e721dd4} /* (30, 16, 3) {real, imag} */,
  {32'hbded626a, 32'hbd978731} /* (30, 16, 2) {real, imag} */,
  {32'h3e055a50, 32'h3dd820f9} /* (30, 16, 1) {real, imag} */,
  {32'hbc0f9638, 32'h00000000} /* (30, 16, 0) {real, imag} */,
  {32'hbd5137f0, 32'h3e1cd7f2} /* (30, 15, 31) {real, imag} */,
  {32'h3d9b0bc8, 32'hbf307e06} /* (30, 15, 30) {real, imag} */,
  {32'h3dbb9036, 32'h3dd3a2a5} /* (30, 15, 29) {real, imag} */,
  {32'h3d28eb47, 32'h3e3d9e08} /* (30, 15, 28) {real, imag} */,
  {32'h3df8cdac, 32'hbd29b848} /* (30, 15, 27) {real, imag} */,
  {32'h3e8b9547, 32'h3d0c4bfa} /* (30, 15, 26) {real, imag} */,
  {32'hbdd9c5ae, 32'h3ea2ab8c} /* (30, 15, 25) {real, imag} */,
  {32'h3e902d09, 32'hbdf1bdab} /* (30, 15, 24) {real, imag} */,
  {32'hbcdcac5c, 32'hbc3a2900} /* (30, 15, 23) {real, imag} */,
  {32'h3df92392, 32'h3e99945e} /* (30, 15, 22) {real, imag} */,
  {32'hbde71c92, 32'h3e0017d3} /* (30, 15, 21) {real, imag} */,
  {32'h3e69525c, 32'hbe40ca8b} /* (30, 15, 20) {real, imag} */,
  {32'hbeeb7a1c, 32'hbe2ca59c} /* (30, 15, 19) {real, imag} */,
  {32'h3d135bfa, 32'h3df79ed0} /* (30, 15, 18) {real, imag} */,
  {32'hbd3c9c93, 32'h3e48a377} /* (30, 15, 17) {real, imag} */,
  {32'h3e730b59, 32'hbe4a2682} /* (30, 15, 16) {real, imag} */,
  {32'h3daa6ccf, 32'hbdb6414a} /* (30, 15, 15) {real, imag} */,
  {32'hbe88d9e7, 32'hbd90f5da} /* (30, 15, 14) {real, imag} */,
  {32'hbd43c7b0, 32'hbe0ce660} /* (30, 15, 13) {real, imag} */,
  {32'h3e63ff33, 32'h3dc66fc9} /* (30, 15, 12) {real, imag} */,
  {32'h3f240fa8, 32'h3e4c3151} /* (30, 15, 11) {real, imag} */,
  {32'hbd9d41be, 32'hbe8236cf} /* (30, 15, 10) {real, imag} */,
  {32'h3d908484, 32'h3d4f85f6} /* (30, 15, 9) {real, imag} */,
  {32'hbec6ef75, 32'h3eedb41a} /* (30, 15, 8) {real, imag} */,
  {32'hbe8ccc96, 32'hbe127e63} /* (30, 15, 7) {real, imag} */,
  {32'h3dc05ef0, 32'h3e19a0b0} /* (30, 15, 6) {real, imag} */,
  {32'hbe3f6420, 32'h3e5b4af5} /* (30, 15, 5) {real, imag} */,
  {32'h3e922e44, 32'h3d5a470e} /* (30, 15, 4) {real, imag} */,
  {32'hbeb2531d, 32'hbd5c54fd} /* (30, 15, 3) {real, imag} */,
  {32'hb9ad1c00, 32'hbedbc9cc} /* (30, 15, 2) {real, imag} */,
  {32'h3c75d9e8, 32'h3e3e077b} /* (30, 15, 1) {real, imag} */,
  {32'h3c89f38c, 32'hbe55801a} /* (30, 15, 0) {real, imag} */,
  {32'h3c34dc6e, 32'hbf15ee2a} /* (30, 14, 31) {real, imag} */,
  {32'h3dbdbca2, 32'h3d626840} /* (30, 14, 30) {real, imag} */,
  {32'h3ccc1550, 32'h3d9afcd6} /* (30, 14, 29) {real, imag} */,
  {32'hbd875a94, 32'hbda29434} /* (30, 14, 28) {real, imag} */,
  {32'h3b2b6fc0, 32'h3e5ddc99} /* (30, 14, 27) {real, imag} */,
  {32'h3f091ebe, 32'hbe0c3e6d} /* (30, 14, 26) {real, imag} */,
  {32'h3e94ddde, 32'h3d07ef20} /* (30, 14, 25) {real, imag} */,
  {32'h3f0c7b1b, 32'h3bdaddb0} /* (30, 14, 24) {real, imag} */,
  {32'hbe56e280, 32'h3d938d8c} /* (30, 14, 23) {real, imag} */,
  {32'hbe6f2772, 32'h3dae0dee} /* (30, 14, 22) {real, imag} */,
  {32'hbd5960a5, 32'hbddc0ab0} /* (30, 14, 21) {real, imag} */,
  {32'hbe7eadc7, 32'hbe147ffa} /* (30, 14, 20) {real, imag} */,
  {32'hbc454308, 32'h3f183775} /* (30, 14, 19) {real, imag} */,
  {32'hbee271c9, 32'h3f06eee4} /* (30, 14, 18) {real, imag} */,
  {32'h3dbcad34, 32'hbdc08fb1} /* (30, 14, 17) {real, imag} */,
  {32'h3e7f8645, 32'hbe7e86b8} /* (30, 14, 16) {real, imag} */,
  {32'h3db8d8b5, 32'h3e304b3c} /* (30, 14, 15) {real, imag} */,
  {32'h3ee2530a, 32'hbe0bf508} /* (30, 14, 14) {real, imag} */,
  {32'hbea19672, 32'hbe0ee620} /* (30, 14, 13) {real, imag} */,
  {32'hbe41b471, 32'hbd464d88} /* (30, 14, 12) {real, imag} */,
  {32'hbcfdbfe0, 32'hbda8926c} /* (30, 14, 11) {real, imag} */,
  {32'hbefee23c, 32'hbd40d8c5} /* (30, 14, 10) {real, imag} */,
  {32'hbe35e323, 32'hbeae52a5} /* (30, 14, 9) {real, imag} */,
  {32'h3ef43b75, 32'h3e5e26dc} /* (30, 14, 8) {real, imag} */,
  {32'h3e155823, 32'hbd8630e8} /* (30, 14, 7) {real, imag} */,
  {32'h3f08589a, 32'h3e59d81e} /* (30, 14, 6) {real, imag} */,
  {32'h3e87fc74, 32'h3d95fe68} /* (30, 14, 5) {real, imag} */,
  {32'hbefd7086, 32'hbf03fc4b} /* (30, 14, 4) {real, imag} */,
  {32'hbd12ac84, 32'h3e45b661} /* (30, 14, 3) {real, imag} */,
  {32'hbd730368, 32'h3db5d37e} /* (30, 14, 2) {real, imag} */,
  {32'hbc290890, 32'hbec5f24a} /* (30, 14, 1) {real, imag} */,
  {32'h3ec3c66e, 32'hbf0cb16e} /* (30, 14, 0) {real, imag} */,
  {32'hbe92dc48, 32'hbea2d0d4} /* (30, 13, 31) {real, imag} */,
  {32'hbec9915e, 32'h3c93b010} /* (30, 13, 30) {real, imag} */,
  {32'h3e209dc6, 32'hbdef6e92} /* (30, 13, 29) {real, imag} */,
  {32'h3e781470, 32'hbe146000} /* (30, 13, 28) {real, imag} */,
  {32'hbea56ae2, 32'hbe2f55e4} /* (30, 13, 27) {real, imag} */,
  {32'h3d8fd739, 32'hbf3d360d} /* (30, 13, 26) {real, imag} */,
  {32'h3c3ed5e0, 32'h3e9aa37d} /* (30, 13, 25) {real, imag} */,
  {32'hbca45f10, 32'h3e0f7e29} /* (30, 13, 24) {real, imag} */,
  {32'hbd11fa60, 32'h3e07d1c2} /* (30, 13, 23) {real, imag} */,
  {32'h3e980f00, 32'hbcc5b310} /* (30, 13, 22) {real, imag} */,
  {32'h3e1cdb3c, 32'hbe053084} /* (30, 13, 21) {real, imag} */,
  {32'hbdfd7d3d, 32'hbe3a843c} /* (30, 13, 20) {real, imag} */,
  {32'hbe98983d, 32'hbd9c37c0} /* (30, 13, 19) {real, imag} */,
  {32'hbf1cba2f, 32'hbc457a50} /* (30, 13, 18) {real, imag} */,
  {32'hbedaf2d2, 32'hbe8300fe} /* (30, 13, 17) {real, imag} */,
  {32'h3e7074f6, 32'hbc9f3a9e} /* (30, 13, 16) {real, imag} */,
  {32'h3ed5e640, 32'hbf10fc78} /* (30, 13, 15) {real, imag} */,
  {32'h3e855c05, 32'hbd9b5b10} /* (30, 13, 14) {real, imag} */,
  {32'hbc41b110, 32'h3e2a2195} /* (30, 13, 13) {real, imag} */,
  {32'hbf0d1bd9, 32'h3da20d74} /* (30, 13, 12) {real, imag} */,
  {32'hbe9393e8, 32'h3e975cd8} /* (30, 13, 11) {real, imag} */,
  {32'hbda2d9c8, 32'hbe6d85c4} /* (30, 13, 10) {real, imag} */,
  {32'hbe275752, 32'hbd124640} /* (30, 13, 9) {real, imag} */,
  {32'hbeb30781, 32'h3c7d7ff0} /* (30, 13, 8) {real, imag} */,
  {32'h3e0516c0, 32'h3efc4d68} /* (30, 13, 7) {real, imag} */,
  {32'h3eea3900, 32'h3d2f1604} /* (30, 13, 6) {real, imag} */,
  {32'hbed5d369, 32'h3ecd0fc2} /* (30, 13, 5) {real, imag} */,
  {32'hbdb5ec2c, 32'hbf0124ab} /* (30, 13, 4) {real, imag} */,
  {32'h3ea02240, 32'hbd4ee400} /* (30, 13, 3) {real, imag} */,
  {32'hbeb997fa, 32'hbd8ecb58} /* (30, 13, 2) {real, imag} */,
  {32'h3f1f5b05, 32'h3dc1d768} /* (30, 13, 1) {real, imag} */,
  {32'h3ded2d6f, 32'h3e34e4e6} /* (30, 13, 0) {real, imag} */,
  {32'hbc18e780, 32'hbd4a38d0} /* (30, 12, 31) {real, imag} */,
  {32'hbd84b48c, 32'h3f0d2cd6} /* (30, 12, 30) {real, imag} */,
  {32'h3e83396c, 32'hbed5d77a} /* (30, 12, 29) {real, imag} */,
  {32'hbe1e51a3, 32'h3e78a863} /* (30, 12, 28) {real, imag} */,
  {32'hbe3879f2, 32'h3e7347be} /* (30, 12, 27) {real, imag} */,
  {32'h3d687a52, 32'hbf27dd56} /* (30, 12, 26) {real, imag} */,
  {32'hbe1df638, 32'h3c2424e0} /* (30, 12, 25) {real, imag} */,
  {32'h3d539486, 32'hbe2d0cbe} /* (30, 12, 24) {real, imag} */,
  {32'hbc7258e8, 32'h3e5a4104} /* (30, 12, 23) {real, imag} */,
  {32'h3ef2e13f, 32'h3e1bed08} /* (30, 12, 22) {real, imag} */,
  {32'h3eee7ce5, 32'h3db9e252} /* (30, 12, 21) {real, imag} */,
  {32'hbed3098a, 32'hbcf88d78} /* (30, 12, 20) {real, imag} */,
  {32'hbf0527cb, 32'hbef3b049} /* (30, 12, 19) {real, imag} */,
  {32'hbe96e3ec, 32'hbec224ac} /* (30, 12, 18) {real, imag} */,
  {32'h3e9949e6, 32'h3eb9ea26} /* (30, 12, 17) {real, imag} */,
  {32'h3cf2f122, 32'h3e8aa61c} /* (30, 12, 16) {real, imag} */,
  {32'h3de2f340, 32'h3de5f8f4} /* (30, 12, 15) {real, imag} */,
  {32'hbd6756a8, 32'h3d8a09d8} /* (30, 12, 14) {real, imag} */,
  {32'hbe8e083b, 32'h3c9470a0} /* (30, 12, 13) {real, imag} */,
  {32'h3ed9882a, 32'h3e122226} /* (30, 12, 12) {real, imag} */,
  {32'hbe91c2c6, 32'h3e9d05c4} /* (30, 12, 11) {real, imag} */,
  {32'hbe883ca8, 32'hbc97b748} /* (30, 12, 10) {real, imag} */,
  {32'hbe23d86e, 32'h3cb5e280} /* (30, 12, 9) {real, imag} */,
  {32'hbe8e824e, 32'h3e63533d} /* (30, 12, 8) {real, imag} */,
  {32'h38e09000, 32'h3e61ea44} /* (30, 12, 7) {real, imag} */,
  {32'h3f00dc04, 32'h3ca81340} /* (30, 12, 6) {real, imag} */,
  {32'hbeb419bb, 32'hbe745c2b} /* (30, 12, 5) {real, imag} */,
  {32'h3c0a7468, 32'hbe22f9da} /* (30, 12, 4) {real, imag} */,
  {32'h3ea6259e, 32'h3df5d25e} /* (30, 12, 3) {real, imag} */,
  {32'hbd0edd60, 32'hbd2b7942} /* (30, 12, 2) {real, imag} */,
  {32'h3e174fb8, 32'h3e7ff5ea} /* (30, 12, 1) {real, imag} */,
  {32'hbd731310, 32'hbe808ecd} /* (30, 12, 0) {real, imag} */,
  {32'hbe00c062, 32'hbeda124a} /* (30, 11, 31) {real, imag} */,
  {32'h3eef55f6, 32'h3ef8a8f4} /* (30, 11, 30) {real, imag} */,
  {32'h3e91fee8, 32'h3e807700} /* (30, 11, 29) {real, imag} */,
  {32'h3ec7f48e, 32'hbdee1e7c} /* (30, 11, 28) {real, imag} */,
  {32'hbdf6c9ca, 32'hbdd341f0} /* (30, 11, 27) {real, imag} */,
  {32'hbec121f4, 32'h3ed07525} /* (30, 11, 26) {real, imag} */,
  {32'hbd58f9c0, 32'hbc800590} /* (30, 11, 25) {real, imag} */,
  {32'hbdd17870, 32'h3ecf13ea} /* (30, 11, 24) {real, imag} */,
  {32'hbd0bba78, 32'hbed8f721} /* (30, 11, 23) {real, imag} */,
  {32'hbf1c0043, 32'hbe3f8a0a} /* (30, 11, 22) {real, imag} */,
  {32'h3eaabc1b, 32'h3e89efe8} /* (30, 11, 21) {real, imag} */,
  {32'h3edc7672, 32'h3e92ad82} /* (30, 11, 20) {real, imag} */,
  {32'hbf05f5ac, 32'h3de96e77} /* (30, 11, 19) {real, imag} */,
  {32'h3eb2d10a, 32'hbe3726ca} /* (30, 11, 18) {real, imag} */,
  {32'h3d32293a, 32'h3ea0ddea} /* (30, 11, 17) {real, imag} */,
  {32'hbea1d6bd, 32'h3dde3d58} /* (30, 11, 16) {real, imag} */,
  {32'h3ea225ef, 32'hbe77a1cf} /* (30, 11, 15) {real, imag} */,
  {32'hbe8a1767, 32'h3c6da5a0} /* (30, 11, 14) {real, imag} */,
  {32'h3e174a51, 32'h3e0229ca} /* (30, 11, 13) {real, imag} */,
  {32'hbbfda970, 32'h3ea2ba80} /* (30, 11, 12) {real, imag} */,
  {32'h3e6e4c9c, 32'hbeaa0132} /* (30, 11, 11) {real, imag} */,
  {32'h3ea996e6, 32'h3e14882b} /* (30, 11, 10) {real, imag} */,
  {32'hbf065044, 32'h3e573561} /* (30, 11, 9) {real, imag} */,
  {32'hbda822ee, 32'hbe6f4c10} /* (30, 11, 8) {real, imag} */,
  {32'h3e94cd2e, 32'hbe22297d} /* (30, 11, 7) {real, imag} */,
  {32'hbe7b842a, 32'hbe030f5e} /* (30, 11, 6) {real, imag} */,
  {32'h3e15f5da, 32'h3cbe0370} /* (30, 11, 5) {real, imag} */,
  {32'h3e0902ec, 32'hbe6d00c0} /* (30, 11, 4) {real, imag} */,
  {32'h3ee6c75a, 32'hbe95b272} /* (30, 11, 3) {real, imag} */,
  {32'hbeb06b0b, 32'h3ef655dd} /* (30, 11, 2) {real, imag} */,
  {32'hbe286b2d, 32'hbeae839f} /* (30, 11, 1) {real, imag} */,
  {32'hbde5903f, 32'hbf44ca47} /* (30, 11, 0) {real, imag} */,
  {32'hbc837ded, 32'h3f244a5a} /* (30, 10, 31) {real, imag} */,
  {32'h3efe9c1b, 32'hbe8fdf20} /* (30, 10, 30) {real, imag} */,
  {32'h3e5fc0dd, 32'hbcf1c478} /* (30, 10, 29) {real, imag} */,
  {32'h3e4bc290, 32'hbebc59b2} /* (30, 10, 28) {real, imag} */,
  {32'h3e37f15a, 32'h3dd20ca5} /* (30, 10, 27) {real, imag} */,
  {32'h3dde485a, 32'hbe16c279} /* (30, 10, 26) {real, imag} */,
  {32'hbd9d5bce, 32'hbe872227} /* (30, 10, 25) {real, imag} */,
  {32'hbeef821e, 32'hbe0b15bb} /* (30, 10, 24) {real, imag} */,
  {32'hbe8af730, 32'hbde47bf4} /* (30, 10, 23) {real, imag} */,
  {32'h3df562e6, 32'hbf3db0e8} /* (30, 10, 22) {real, imag} */,
  {32'hbf3b61aa, 32'hbd33b9c8} /* (30, 10, 21) {real, imag} */,
  {32'h3e40898e, 32'h3f21188e} /* (30, 10, 20) {real, imag} */,
  {32'h3f360d69, 32'h3e1ea928} /* (30, 10, 19) {real, imag} */,
  {32'h3e61b281, 32'hbecb7c42} /* (30, 10, 18) {real, imag} */,
  {32'h3d331994, 32'h3df661a1} /* (30, 10, 17) {real, imag} */,
  {32'hbe60bd61, 32'h3cd47bb8} /* (30, 10, 16) {real, imag} */,
  {32'hbe07a3f2, 32'h3e8cb621} /* (30, 10, 15) {real, imag} */,
  {32'hbd82409c, 32'h3e04bffa} /* (30, 10, 14) {real, imag} */,
  {32'h3f71c158, 32'hbe957f1e} /* (30, 10, 13) {real, imag} */,
  {32'hbf1ec2e5, 32'h3e3aa276} /* (30, 10, 12) {real, imag} */,
  {32'h3e0059c2, 32'h3e042ad2} /* (30, 10, 11) {real, imag} */,
  {32'hbe66cd6b, 32'h3ec84332} /* (30, 10, 10) {real, imag} */,
  {32'h3e874a44, 32'h3d547fa0} /* (30, 10, 9) {real, imag} */,
  {32'h3e4f3be3, 32'hbea20cc7} /* (30, 10, 8) {real, imag} */,
  {32'h3eb9ce38, 32'h3edd0a30} /* (30, 10, 7) {real, imag} */,
  {32'hbdfea1aa, 32'hbf28ad98} /* (30, 10, 6) {real, imag} */,
  {32'hbe88b1d6, 32'hbe80da76} /* (30, 10, 5) {real, imag} */,
  {32'hbe479b4a, 32'h3829a000} /* (30, 10, 4) {real, imag} */,
  {32'h3e1b1c70, 32'h3e86a8e6} /* (30, 10, 3) {real, imag} */,
  {32'hbeeef0b4, 32'hbf127529} /* (30, 10, 2) {real, imag} */,
  {32'hbe95bedf, 32'h3d5a6bac} /* (30, 10, 1) {real, imag} */,
  {32'hbd9c8662, 32'hbec188d2} /* (30, 10, 0) {real, imag} */,
  {32'hbf0ed06e, 32'h3eb8c11c} /* (30, 9, 31) {real, imag} */,
  {32'h3e4232de, 32'hbdc39528} /* (30, 9, 30) {real, imag} */,
  {32'hbf0f4920, 32'h3f31f972} /* (30, 9, 29) {real, imag} */,
  {32'hbd75d16e, 32'h3e52beca} /* (30, 9, 28) {real, imag} */,
  {32'hbede196a, 32'hbed292ae} /* (30, 9, 27) {real, imag} */,
  {32'h3eb1e7da, 32'h3e94b30d} /* (30, 9, 26) {real, imag} */,
  {32'h3df8e610, 32'hbe984bdd} /* (30, 9, 25) {real, imag} */,
  {32'hbef965c9, 32'hbf3694d7} /* (30, 9, 24) {real, imag} */,
  {32'hbdd75508, 32'hbe7ba745} /* (30, 9, 23) {real, imag} */,
  {32'h3e259cd6, 32'h3ea737c6} /* (30, 9, 22) {real, imag} */,
  {32'h3e84c942, 32'h3ebee5ad} /* (30, 9, 21) {real, imag} */,
  {32'h3f07d16d, 32'hbe9eea4b} /* (30, 9, 20) {real, imag} */,
  {32'hbe997830, 32'hbde0e2ab} /* (30, 9, 19) {real, imag} */,
  {32'h3e373258, 32'hbf0cbd82} /* (30, 9, 18) {real, imag} */,
  {32'h3dc1f254, 32'h3cba6898} /* (30, 9, 17) {real, imag} */,
  {32'h3e3c6a7a, 32'hbc04cc40} /* (30, 9, 16) {real, imag} */,
  {32'hbe03cfec, 32'h3d510ef0} /* (30, 9, 15) {real, imag} */,
  {32'hbef8098c, 32'h3ea64943} /* (30, 9, 14) {real, imag} */,
  {32'hbe83398a, 32'hbce5778c} /* (30, 9, 13) {real, imag} */,
  {32'h3e727e2a, 32'hbf07b336} /* (30, 9, 12) {real, imag} */,
  {32'hbe677c3a, 32'h3cf765c0} /* (30, 9, 11) {real, imag} */,
  {32'hbe2a0f40, 32'hbe9abc9b} /* (30, 9, 10) {real, imag} */,
  {32'h3eaf055c, 32'h3d958a74} /* (30, 9, 9) {real, imag} */,
  {32'hbd8fb214, 32'h3e03d40c} /* (30, 9, 8) {real, imag} */,
  {32'h3e5e55f9, 32'hbf0ce627} /* (30, 9, 7) {real, imag} */,
  {32'hbd4e00d2, 32'hbde30438} /* (30, 9, 6) {real, imag} */,
  {32'h3e45e35f, 32'h3f01f461} /* (30, 9, 5) {real, imag} */,
  {32'h3df4c8e1, 32'h3ebd72f0} /* (30, 9, 4) {real, imag} */,
  {32'hbf437583, 32'hbecabf67} /* (30, 9, 3) {real, imag} */,
  {32'hbf7117be, 32'hbf42bc3e} /* (30, 9, 2) {real, imag} */,
  {32'h3f545051, 32'h3e1e398e} /* (30, 9, 1) {real, imag} */,
  {32'h3dda2068, 32'h3e7c53fe} /* (30, 9, 0) {real, imag} */,
  {32'hbf8c8f3f, 32'hbf322d7c} /* (30, 8, 31) {real, imag} */,
  {32'h3f90b064, 32'h3c2c1720} /* (30, 8, 30) {real, imag} */,
  {32'hbebf5af0, 32'hbf187ff3} /* (30, 8, 29) {real, imag} */,
  {32'hbd958e38, 32'h3ed515d3} /* (30, 8, 28) {real, imag} */,
  {32'hbe1ae594, 32'h3e7f5602} /* (30, 8, 27) {real, imag} */,
  {32'h3d9f7754, 32'h3e9d7536} /* (30, 8, 26) {real, imag} */,
  {32'h3d8a2bb4, 32'hbece5c8b} /* (30, 8, 25) {real, imag} */,
  {32'h3e0cefeb, 32'hbdac7548} /* (30, 8, 24) {real, imag} */,
  {32'hbe084798, 32'h3db48eb0} /* (30, 8, 23) {real, imag} */,
  {32'h3dfc39da, 32'hbeba9878} /* (30, 8, 22) {real, imag} */,
  {32'h3dba114e, 32'hbecb43ca} /* (30, 8, 21) {real, imag} */,
  {32'h3de492b8, 32'hbe2bb85a} /* (30, 8, 20) {real, imag} */,
  {32'h3ea380d8, 32'h3d2f3668} /* (30, 8, 19) {real, imag} */,
  {32'hbd6e6366, 32'h3e6dcf2f} /* (30, 8, 18) {real, imag} */,
  {32'h3f0c39fe, 32'h3ddd06e5} /* (30, 8, 17) {real, imag} */,
  {32'hbeb82322, 32'h3e170fcc} /* (30, 8, 16) {real, imag} */,
  {32'hbe7ce68a, 32'hbd7bb210} /* (30, 8, 15) {real, imag} */,
  {32'hbd8e7770, 32'hbf01f9c7} /* (30, 8, 14) {real, imag} */,
  {32'hbd937ce0, 32'hbe8a1193} /* (30, 8, 13) {real, imag} */,
  {32'hbee3c9f2, 32'h3e0388ee} /* (30, 8, 12) {real, imag} */,
  {32'hbca0c910, 32'h3dce748c} /* (30, 8, 11) {real, imag} */,
  {32'h3dc26b7e, 32'h3f0358a9} /* (30, 8, 10) {real, imag} */,
  {32'hbe965bf5, 32'hbecaefe6} /* (30, 8, 9) {real, imag} */,
  {32'hbe84fe0f, 32'hbd7b56b6} /* (30, 8, 8) {real, imag} */,
  {32'hbe795c26, 32'h3ede36ea} /* (30, 8, 7) {real, imag} */,
  {32'h3da52170, 32'h3ea6649a} /* (30, 8, 6) {real, imag} */,
  {32'h3eac15fa, 32'h3e007bad} /* (30, 8, 5) {real, imag} */,
  {32'hbf1471d2, 32'h3e878619} /* (30, 8, 4) {real, imag} */,
  {32'hbeb001c4, 32'h3ef02912} /* (30, 8, 3) {real, imag} */,
  {32'h3f1b5584, 32'h3fa504e6} /* (30, 8, 2) {real, imag} */,
  {32'hbf332438, 32'hbf6df06f} /* (30, 8, 1) {real, imag} */,
  {32'hbf9f2882, 32'h3d6d2c20} /* (30, 8, 0) {real, imag} */,
  {32'h3e51cba9, 32'h3eb5a8d2} /* (30, 7, 31) {real, imag} */,
  {32'hbf0689a4, 32'hbeea6674} /* (30, 7, 30) {real, imag} */,
  {32'h3e6e91b0, 32'h3ea55a68} /* (30, 7, 29) {real, imag} */,
  {32'hbf444bba, 32'hbc1fae30} /* (30, 7, 28) {real, imag} */,
  {32'hbec4aa52, 32'hbea34d83} /* (30, 7, 27) {real, imag} */,
  {32'h3ec798e6, 32'h3f2581d0} /* (30, 7, 26) {real, imag} */,
  {32'hbf0697da, 32'hbd739020} /* (30, 7, 25) {real, imag} */,
  {32'hbddc959c, 32'h3cd6a23c} /* (30, 7, 24) {real, imag} */,
  {32'h3e9dc2e9, 32'h3eabfa4d} /* (30, 7, 23) {real, imag} */,
  {32'hbe09818a, 32'hbe0bd4d5} /* (30, 7, 22) {real, imag} */,
  {32'h3ee23703, 32'h3db635cb} /* (30, 7, 21) {real, imag} */,
  {32'hbef1bda8, 32'h3d4918b8} /* (30, 7, 20) {real, imag} */,
  {32'h3e3cceba, 32'hbe83d585} /* (30, 7, 19) {real, imag} */,
  {32'h3df5cd34, 32'h3d7a7830} /* (30, 7, 18) {real, imag} */,
  {32'hbe9caaf4, 32'h3ca28cfc} /* (30, 7, 17) {real, imag} */,
  {32'h3eb1ac6d, 32'hbd56d25a} /* (30, 7, 16) {real, imag} */,
  {32'hbdfa5d28, 32'hbdd66ab7} /* (30, 7, 15) {real, imag} */,
  {32'hbe9ff05d, 32'h3d478734} /* (30, 7, 14) {real, imag} */,
  {32'h3e9ceef9, 32'hbd726084} /* (30, 7, 13) {real, imag} */,
  {32'h3dcc8518, 32'hbdd75962} /* (30, 7, 12) {real, imag} */,
  {32'h3dc641d6, 32'h3d91d657} /* (30, 7, 11) {real, imag} */,
  {32'h3ead0b25, 32'h3e95a868} /* (30, 7, 10) {real, imag} */,
  {32'h3d8fd6ac, 32'hbd67c2e8} /* (30, 7, 9) {real, imag} */,
  {32'h3eb1bb08, 32'h3d92e5c4} /* (30, 7, 8) {real, imag} */,
  {32'h3db1f4d7, 32'hbe15bfd4} /* (30, 7, 7) {real, imag} */,
  {32'h3e043dea, 32'hbe464d82} /* (30, 7, 6) {real, imag} */,
  {32'h3ed786f6, 32'h3e9063f8} /* (30, 7, 5) {real, imag} */,
  {32'h3dd01f4c, 32'h3dbcfb98} /* (30, 7, 4) {real, imag} */,
  {32'h3e050b90, 32'hbe92043d} /* (30, 7, 3) {real, imag} */,
  {32'h3f1e2ee1, 32'hbef9c2d0} /* (30, 7, 2) {real, imag} */,
  {32'hbe3d6db2, 32'h3eeef9e3} /* (30, 7, 1) {real, imag} */,
  {32'h3f46a4ad, 32'h3e35171e} /* (30, 7, 0) {real, imag} */,
  {32'hbf287fe7, 32'h3f97ef32} /* (30, 6, 31) {real, imag} */,
  {32'hbf1e0e33, 32'h3e33dfed} /* (30, 6, 30) {real, imag} */,
  {32'h3ddb73e8, 32'hbf28213e} /* (30, 6, 29) {real, imag} */,
  {32'hbd580430, 32'hbd6085c0} /* (30, 6, 28) {real, imag} */,
  {32'h3d3770f2, 32'h3e8c30b1} /* (30, 6, 27) {real, imag} */,
  {32'h3eb1d327, 32'h3f2e08e8} /* (30, 6, 26) {real, imag} */,
  {32'h3d0cef84, 32'hbd259848} /* (30, 6, 25) {real, imag} */,
  {32'h3f0ad94a, 32'hbee9030b} /* (30, 6, 24) {real, imag} */,
  {32'hbd0a9284, 32'hbe0fc940} /* (30, 6, 23) {real, imag} */,
  {32'h3de41684, 32'hbd66d9a0} /* (30, 6, 22) {real, imag} */,
  {32'hbe960f55, 32'h3d7131b8} /* (30, 6, 21) {real, imag} */,
  {32'hbf02fe59, 32'h3e4346d2} /* (30, 6, 20) {real, imag} */,
  {32'hbf24ee8c, 32'hbeeaadce} /* (30, 6, 19) {real, imag} */,
  {32'h3f013200, 32'h3ead4bfe} /* (30, 6, 18) {real, imag} */,
  {32'hbd8535b6, 32'hbea8c4b4} /* (30, 6, 17) {real, imag} */,
  {32'h3e806c63, 32'hbe4b91b6} /* (30, 6, 16) {real, imag} */,
  {32'hbe4f65f8, 32'h3e065fbc} /* (30, 6, 15) {real, imag} */,
  {32'h3dbd65c1, 32'h3e1ffa9c} /* (30, 6, 14) {real, imag} */,
  {32'h3e09b9b2, 32'h3e52a89b} /* (30, 6, 13) {real, imag} */,
  {32'hbed475ce, 32'hbe3759a2} /* (30, 6, 12) {real, imag} */,
  {32'h3db62000, 32'hbe5e3954} /* (30, 6, 11) {real, imag} */,
  {32'h3df23bd8, 32'hbf08211b} /* (30, 6, 10) {real, imag} */,
  {32'hbeec06c4, 32'h3e88b9da} /* (30, 6, 9) {real, imag} */,
  {32'h3e10d4ec, 32'h3de4432c} /* (30, 6, 8) {real, imag} */,
  {32'h3d93c534, 32'h3ea3cba9} /* (30, 6, 7) {real, imag} */,
  {32'hbf00f4e0, 32'h3ee6e546} /* (30, 6, 6) {real, imag} */,
  {32'h3f3200d6, 32'h3eae0121} /* (30, 6, 5) {real, imag} */,
  {32'h3ed8ef52, 32'h3d02cc2c} /* (30, 6, 4) {real, imag} */,
  {32'hbe9d94b9, 32'h3e84dd62} /* (30, 6, 3) {real, imag} */,
  {32'h3db392c0, 32'hbecb219a} /* (30, 6, 2) {real, imag} */,
  {32'hbf9b5ed5, 32'hbe92e702} /* (30, 6, 1) {real, imag} */,
  {32'h3f3b76e3, 32'h3dc5bf5b} /* (30, 6, 0) {real, imag} */,
  {32'hc01f0a5e, 32'hbed0e478} /* (30, 5, 31) {real, imag} */,
  {32'h3f382820, 32'hbf8b0019} /* (30, 5, 30) {real, imag} */,
  {32'h3e12d792, 32'hbe128776} /* (30, 5, 29) {real, imag} */,
  {32'h3ea4fc64, 32'h3ed45c23} /* (30, 5, 28) {real, imag} */,
  {32'h3f55bf3b, 32'hbd8f45c6} /* (30, 5, 27) {real, imag} */,
  {32'hbe784284, 32'h3d9ea044} /* (30, 5, 26) {real, imag} */,
  {32'hbf376f45, 32'h3eb0e778} /* (30, 5, 25) {real, imag} */,
  {32'hbda01f6e, 32'h3f0ab02e} /* (30, 5, 24) {real, imag} */,
  {32'hbed13b06, 32'hbe88c0c7} /* (30, 5, 23) {real, imag} */,
  {32'h3d4e1470, 32'hbf686c70} /* (30, 5, 22) {real, imag} */,
  {32'h3e39d914, 32'hbce69868} /* (30, 5, 21) {real, imag} */,
  {32'hbe1a1fad, 32'hbdfe8696} /* (30, 5, 20) {real, imag} */,
  {32'h3e124e91, 32'hbddb4768} /* (30, 5, 19) {real, imag} */,
  {32'hbe87ba82, 32'hbcb7e630} /* (30, 5, 18) {real, imag} */,
  {32'hbe020c95, 32'hbd5b1ac2} /* (30, 5, 17) {real, imag} */,
  {32'hbdc4c6d9, 32'h3dd97a15} /* (30, 5, 16) {real, imag} */,
  {32'hbe1e57c3, 32'h3d45a6f4} /* (30, 5, 15) {real, imag} */,
  {32'h3d4183de, 32'h3e6235ca} /* (30, 5, 14) {real, imag} */,
  {32'h3e7a1402, 32'h3c44d0c0} /* (30, 5, 13) {real, imag} */,
  {32'hbdbc5990, 32'h3ef987d1} /* (30, 5, 12) {real, imag} */,
  {32'hbf29fc6d, 32'h3dac69c4} /* (30, 5, 11) {real, imag} */,
  {32'hbd581dea, 32'h3df22fb6} /* (30, 5, 10) {real, imag} */,
  {32'h3e04106e, 32'h3f056184} /* (30, 5, 9) {real, imag} */,
  {32'hbe9cf8d5, 32'h3edde052} /* (30, 5, 8) {real, imag} */,
  {32'h3ed540df, 32'hbef60a79} /* (30, 5, 7) {real, imag} */,
  {32'h3f08efa0, 32'hbd5322ec} /* (30, 5, 6) {real, imag} */,
  {32'hbeeecd65, 32'h3f0397dc} /* (30, 5, 5) {real, imag} */,
  {32'hbf1401c5, 32'hbf1075ac} /* (30, 5, 4) {real, imag} */,
  {32'hbe07ca4c, 32'hbb714fc0} /* (30, 5, 3) {real, imag} */,
  {32'h3fc840ea, 32'h3f997758} /* (30, 5, 2) {real, imag} */,
  {32'hbfe85825, 32'hc004576e} /* (30, 5, 1) {real, imag} */,
  {32'hc011a4a3, 32'h3e6b5d26} /* (30, 5, 0) {real, imag} */,
  {32'h3fe08b95, 32'h40020672} /* (30, 4, 31) {real, imag} */,
  {32'hc03e70cc, 32'hbde8fcf0} /* (30, 4, 30) {real, imag} */,
  {32'hbe743d2a, 32'h3f6aa4fc} /* (30, 4, 29) {real, imag} */,
  {32'h3f8456f6, 32'h3f3fa27a} /* (30, 4, 28) {real, imag} */,
  {32'hbf731231, 32'hbecc2f3e} /* (30, 4, 27) {real, imag} */,
  {32'hbb556980, 32'h3c6bd640} /* (30, 4, 26) {real, imag} */,
  {32'hbee70735, 32'hbe055dcf} /* (30, 4, 25) {real, imag} */,
  {32'hbd947ad1, 32'hbdc0b6f4} /* (30, 4, 24) {real, imag} */,
  {32'h3eb88d6a, 32'h3e2ed6cc} /* (30, 4, 23) {real, imag} */,
  {32'h3efcc0b4, 32'hbd8e9a2c} /* (30, 4, 22) {real, imag} */,
  {32'hbf0f906e, 32'h3e91c2d4} /* (30, 4, 21) {real, imag} */,
  {32'h3dd2ee7b, 32'hbeaa1db6} /* (30, 4, 20) {real, imag} */,
  {32'h3df3f710, 32'h3ddb3409} /* (30, 4, 19) {real, imag} */,
  {32'h3dbb39a8, 32'h3ea7093e} /* (30, 4, 18) {real, imag} */,
  {32'h3e24b966, 32'hbda3b0fc} /* (30, 4, 17) {real, imag} */,
  {32'hbeaf5a5c, 32'hbcd0cb5e} /* (30, 4, 16) {real, imag} */,
  {32'h3df835ca, 32'hbcf7d3c0} /* (30, 4, 15) {real, imag} */,
  {32'hbdecddf0, 32'hbdaf1f6c} /* (30, 4, 14) {real, imag} */,
  {32'h3e843fae, 32'hbe01e9d0} /* (30, 4, 13) {real, imag} */,
  {32'hbbf523d0, 32'hbeb2ec21} /* (30, 4, 12) {real, imag} */,
  {32'h3eb51043, 32'hbe70734c} /* (30, 4, 11) {real, imag} */,
  {32'hbf1261bf, 32'h3f450aba} /* (30, 4, 10) {real, imag} */,
  {32'h3f1798d1, 32'hbcf54592} /* (30, 4, 9) {real, imag} */,
  {32'hbd11c210, 32'h3e7111a4} /* (30, 4, 8) {real, imag} */,
  {32'h3f279a69, 32'h3f604ac4} /* (30, 4, 7) {real, imag} */,
  {32'hbc4a2cf0, 32'hbe8da080} /* (30, 4, 6) {real, imag} */,
  {32'h3efdf056, 32'hbf58f569} /* (30, 4, 5) {real, imag} */,
  {32'hbd8600f4, 32'h3f6cb9e9} /* (30, 4, 4) {real, imag} */,
  {32'h3e43c42e, 32'h3f06919d} /* (30, 4, 3) {real, imag} */,
  {32'hbfa12f4a, 32'hc0118674} /* (30, 4, 2) {real, imag} */,
  {32'h4080b95a, 32'h400a6147} /* (30, 4, 1) {real, imag} */,
  {32'h4008bf4e, 32'h3f29079d} /* (30, 4, 0) {real, imag} */,
  {32'hc036eec5, 32'h401606d2} /* (30, 3, 31) {real, imag} */,
  {32'h3fe322f8, 32'hc01a2415} /* (30, 3, 30) {real, imag} */,
  {32'h3eb8d2b4, 32'h3eb8d840} /* (30, 3, 29) {real, imag} */,
  {32'h3dadb324, 32'h3f2cd2ee} /* (30, 3, 28) {real, imag} */,
  {32'h3e3148a3, 32'hbf1bf8b4} /* (30, 3, 27) {real, imag} */,
  {32'h3dacf338, 32'hbe1d30f0} /* (30, 3, 26) {real, imag} */,
  {32'hbe9fd18d, 32'h3e977b6e} /* (30, 3, 25) {real, imag} */,
  {32'hbe9da3a4, 32'hbc6de760} /* (30, 3, 24) {real, imag} */,
  {32'h3cdd1d40, 32'h3dc0569c} /* (30, 3, 23) {real, imag} */,
  {32'hb9fcf580, 32'h3eac0f0b} /* (30, 3, 22) {real, imag} */,
  {32'hbecdbfc9, 32'h3e0d0915} /* (30, 3, 21) {real, imag} */,
  {32'hbefad778, 32'h3d9371e4} /* (30, 3, 20) {real, imag} */,
  {32'hbe2dddc2, 32'h3e66501a} /* (30, 3, 19) {real, imag} */,
  {32'h3d7a41db, 32'h3d30baf8} /* (30, 3, 18) {real, imag} */,
  {32'h3e320d94, 32'hbe1062ce} /* (30, 3, 17) {real, imag} */,
  {32'hbad1b640, 32'hbeffa722} /* (30, 3, 16) {real, imag} */,
  {32'h3da5959d, 32'h3deb5d44} /* (30, 3, 15) {real, imag} */,
  {32'hbd04a0f0, 32'hbd325bc0} /* (30, 3, 14) {real, imag} */,
  {32'h3ecd5ac8, 32'h3e9b256e} /* (30, 3, 13) {real, imag} */,
  {32'hbe22c39c, 32'hbe608925} /* (30, 3, 12) {real, imag} */,
  {32'hbe964c3f, 32'h3ec198a1} /* (30, 3, 11) {real, imag} */,
  {32'hbf11b68a, 32'hbefe70c3} /* (30, 3, 10) {real, imag} */,
  {32'h3e15c2aa, 32'h3e47d443} /* (30, 3, 9) {real, imag} */,
  {32'hbde25cf7, 32'hbe2beb4c} /* (30, 3, 8) {real, imag} */,
  {32'h3f3d5a26, 32'h3e85a390} /* (30, 3, 7) {real, imag} */,
  {32'hbcfa5d40, 32'h3e18577e} /* (30, 3, 6) {real, imag} */,
  {32'hbf5df5c5, 32'h3f0f1870} /* (30, 3, 5) {real, imag} */,
  {32'hbe68d1cc, 32'h3f15f5e1} /* (30, 3, 4) {real, imag} */,
  {32'h3f54574d, 32'h3dc10af0} /* (30, 3, 3) {real, imag} */,
  {32'hbe539334, 32'hc00bb6a3} /* (30, 3, 2) {real, imag} */,
  {32'h3fe21b78, 32'h3fdd548c} /* (30, 3, 1) {real, imag} */,
  {32'hbebfa95e, 32'h3f17dbf8} /* (30, 3, 0) {real, imag} */,
  {32'hc19425c8, 32'hc00b522d} /* (30, 2, 31) {real, imag} */,
  {32'h411c9632, 32'hc072ba10} /* (30, 2, 30) {real, imag} */,
  {32'h3f971962, 32'h3dbe4ad4} /* (30, 2, 29) {real, imag} */,
  {32'hbfcc6cd7, 32'h4035afd4} /* (30, 2, 28) {real, imag} */,
  {32'h3fb6c4f6, 32'hbe9f778e} /* (30, 2, 27) {real, imag} */,
  {32'h3f0ee529, 32'h3e8e4f4a} /* (30, 2, 26) {real, imag} */,
  {32'hbeb5bba6, 32'hbe6836ca} /* (30, 2, 25) {real, imag} */,
  {32'h3fae19b9, 32'hbea64456} /* (30, 2, 24) {real, imag} */,
  {32'h3cca5ee0, 32'h3e4d3253} /* (30, 2, 23) {real, imag} */,
  {32'hbea5b02e, 32'h3e0b10c2} /* (30, 2, 22) {real, imag} */,
  {32'hbe2974d3, 32'hbef3507e} /* (30, 2, 21) {real, imag} */,
  {32'hbdcd99d1, 32'h3ef07dc8} /* (30, 2, 20) {real, imag} */,
  {32'hbd9dc810, 32'hbe2fe492} /* (30, 2, 19) {real, imag} */,
  {32'hbe11d9f6, 32'hbefa90a0} /* (30, 2, 18) {real, imag} */,
  {32'h3e9e51fd, 32'hbe6ce93b} /* (30, 2, 17) {real, imag} */,
  {32'h3daf37a3, 32'h3df8583c} /* (30, 2, 16) {real, imag} */,
  {32'hbe8ddf8d, 32'h3da48edc} /* (30, 2, 15) {real, imag} */,
  {32'hbc7f0570, 32'hbd11b640} /* (30, 2, 14) {real, imag} */,
  {32'hbea96c5a, 32'hbcb6d1be} /* (30, 2, 13) {real, imag} */,
  {32'h3c95ef50, 32'hbec91cc6} /* (30, 2, 12) {real, imag} */,
  {32'h3f5159aa, 32'h3f8343f8} /* (30, 2, 11) {real, imag} */,
  {32'h3a81ad00, 32'hbea88ab8} /* (30, 2, 10) {real, imag} */,
  {32'h3f10a162, 32'h3d80af9b} /* (30, 2, 9) {real, imag} */,
  {32'h3e94623a, 32'h3dcc80cc} /* (30, 2, 8) {real, imag} */,
  {32'h3e613ed8, 32'hbf2ea44b} /* (30, 2, 7) {real, imag} */,
  {32'h3db3ab24, 32'h3eca03fe} /* (30, 2, 6) {real, imag} */,
  {32'h3fcc8b2c, 32'h3ec4d83c} /* (30, 2, 5) {real, imag} */,
  {32'hbfca1882, 32'h3e81c8f0} /* (30, 2, 4) {real, imag} */,
  {32'hbf93b24c, 32'hbf9ef420} /* (30, 2, 3) {real, imag} */,
  {32'h40e04551, 32'hbf27d804} /* (30, 2, 2) {real, imag} */,
  {32'hc14c7bde, 32'h4094ae16} /* (30, 2, 1) {real, imag} */,
  {32'hc126596a, 32'hbf816126} /* (30, 2, 0) {real, imag} */,
  {32'h418cc7f4, 32'hc09c48f1} /* (30, 1, 31) {real, imag} */,
  {32'hc0e8e09c, 32'h3f46c33f} /* (30, 1, 30) {real, imag} */,
  {32'hbf3856be, 32'h3d8f5720} /* (30, 1, 29) {real, imag} */,
  {32'h3fd8ebff, 32'h3eda0434} /* (30, 1, 28) {real, imag} */,
  {32'hc01085d0, 32'hbdd918e3} /* (30, 1, 27) {real, imag} */,
  {32'hbf096380, 32'hbf193bbc} /* (30, 1, 26) {real, imag} */,
  {32'h3f016a50, 32'hbf875831} /* (30, 1, 25) {real, imag} */,
  {32'hbea44c3c, 32'h3f8901d8} /* (30, 1, 24) {real, imag} */,
  {32'hbee073d7, 32'hbd66efc4} /* (30, 1, 23) {real, imag} */,
  {32'h3ea65ee8, 32'hbed41d05} /* (30, 1, 22) {real, imag} */,
  {32'hbe77277c, 32'h3f95520f} /* (30, 1, 21) {real, imag} */,
  {32'h3eaf6794, 32'h3c9b6f90} /* (30, 1, 20) {real, imag} */,
  {32'h3e24a62a, 32'h3da07b78} /* (30, 1, 19) {real, imag} */,
  {32'hbec54006, 32'h3f0c791b} /* (30, 1, 18) {real, imag} */,
  {32'h3de3144b, 32'hbe25d5b4} /* (30, 1, 17) {real, imag} */,
  {32'h3d6a57ea, 32'h3c116758} /* (30, 1, 16) {real, imag} */,
  {32'hbed89c5c, 32'hbd08bd24} /* (30, 1, 15) {real, imag} */,
  {32'hbdf9a088, 32'hbe66a9ed} /* (30, 1, 14) {real, imag} */,
  {32'h3e0fc74a, 32'h3f15c9ad} /* (30, 1, 13) {real, imag} */,
  {32'h3ef9c11e, 32'hbe1b6199} /* (30, 1, 12) {real, imag} */,
  {32'hbcb25a50, 32'hbea9db26} /* (30, 1, 11) {real, imag} */,
  {32'hbebf4064, 32'h3dfe9342} /* (30, 1, 10) {real, imag} */,
  {32'h3f18db4c, 32'h3eb9a8f2} /* (30, 1, 9) {real, imag} */,
  {32'h3d063858, 32'hbfd27a4a} /* (30, 1, 8) {real, imag} */,
  {32'hbef184f2, 32'h3f13b1cb} /* (30, 1, 7) {real, imag} */,
  {32'hbf32c782, 32'h3f359bb4} /* (30, 1, 6) {real, imag} */,
  {32'hc038d91a, 32'hbf93a988} /* (30, 1, 5) {real, imag} */,
  {32'h3f99e16e, 32'h3dc17f90} /* (30, 1, 4) {real, imag} */,
  {32'hbf5471d1, 32'h3fe25256} /* (30, 1, 3) {real, imag} */,
  {32'hc11e4521, 32'hc130ccd0} /* (30, 1, 2) {real, imag} */,
  {32'h41c21f17, 32'h41227cc4} /* (30, 1, 1) {real, imag} */,
  {32'h416a7508, 32'h405c2030} /* (30, 1, 0) {real, imag} */,
  {32'h4116b5b5, 32'hc107eb1d} /* (30, 0, 31) {real, imag} */,
  {32'hc023310d, 32'h40d9e4c2} /* (30, 0, 30) {real, imag} */,
  {32'hbf0f67ac, 32'h3e33bea8} /* (30, 0, 29) {real, imag} */,
  {32'hbe279b62, 32'h3f983828} /* (30, 0, 28) {real, imag} */,
  {32'hbf84d0e0, 32'hbe88d736} /* (30, 0, 27) {real, imag} */,
  {32'hbed5bc83, 32'hbe73985c} /* (30, 0, 26) {real, imag} */,
  {32'hbf3f91c0, 32'hbf25d6ba} /* (30, 0, 25) {real, imag} */,
  {32'hbf200882, 32'h3f57d573} /* (30, 0, 24) {real, imag} */,
  {32'hbdb93eb2, 32'h3f2244c4} /* (30, 0, 23) {real, imag} */,
  {32'h3e171eed, 32'hbe0b66a1} /* (30, 0, 22) {real, imag} */,
  {32'hbd3b1660, 32'hbd9b0dd0} /* (30, 0, 21) {real, imag} */,
  {32'hbd355350, 32'hbea081c7} /* (30, 0, 20) {real, imag} */,
  {32'h3d37e9bc, 32'hbdb7545b} /* (30, 0, 19) {real, imag} */,
  {32'h3e4f8ec4, 32'h3e17dd0a} /* (30, 0, 18) {real, imag} */,
  {32'h3eea8982, 32'h3d328282} /* (30, 0, 17) {real, imag} */,
  {32'hbea72180, 32'h00000000} /* (30, 0, 16) {real, imag} */,
  {32'h3eea8982, 32'hbd328282} /* (30, 0, 15) {real, imag} */,
  {32'h3e4f8ec4, 32'hbe17dd0a} /* (30, 0, 14) {real, imag} */,
  {32'h3d37e9bc, 32'h3db7545b} /* (30, 0, 13) {real, imag} */,
  {32'hbd355350, 32'h3ea081c7} /* (30, 0, 12) {real, imag} */,
  {32'hbd3b1660, 32'h3d9b0dd0} /* (30, 0, 11) {real, imag} */,
  {32'h3e171eed, 32'h3e0b66a1} /* (30, 0, 10) {real, imag} */,
  {32'hbdb93eb2, 32'hbf2244c4} /* (30, 0, 9) {real, imag} */,
  {32'hbf200882, 32'hbf57d573} /* (30, 0, 8) {real, imag} */,
  {32'hbf3f91c0, 32'h3f25d6ba} /* (30, 0, 7) {real, imag} */,
  {32'hbed5bc83, 32'h3e73985c} /* (30, 0, 6) {real, imag} */,
  {32'hbf84d0e0, 32'h3e88d736} /* (30, 0, 5) {real, imag} */,
  {32'hbe279b62, 32'hbf983828} /* (30, 0, 4) {real, imag} */,
  {32'hbf0f67ac, 32'hbe33bea8} /* (30, 0, 3) {real, imag} */,
  {32'hc023310d, 32'hc0d9e4c2} /* (30, 0, 2) {real, imag} */,
  {32'h4116b5b5, 32'h4107eb1d} /* (30, 0, 1) {real, imag} */,
  {32'h402338ba, 32'h00000000} /* (30, 0, 0) {real, imag} */,
  {32'h41e981a4, 32'hc1456bdc} /* (29, 31, 31) {real, imag} */,
  {32'hc140cccc, 32'h4163363a} /* (29, 31, 30) {real, imag} */,
  {32'hbf46232c, 32'hbfc49552} /* (29, 31, 29) {real, imag} */,
  {32'h3fbcf852, 32'hbf8e7a8a} /* (29, 31, 28) {real, imag} */,
  {32'hc00d7d19, 32'h3f862d79} /* (29, 31, 27) {real, imag} */,
  {32'hbea3bcfc, 32'hbed5cc87} /* (29, 31, 26) {real, imag} */,
  {32'hbeb03fd2, 32'hbe80b5bc} /* (29, 31, 25) {real, imag} */,
  {32'hbe53e927, 32'h3f62fc62} /* (29, 31, 24) {real, imag} */,
  {32'hbeac2cae, 32'hbe58be7f} /* (29, 31, 23) {real, imag} */,
  {32'hbf5014ec, 32'hbcefafe0} /* (29, 31, 22) {real, imag} */,
  {32'h3e22a97c, 32'h3ef7e64d} /* (29, 31, 21) {real, imag} */,
  {32'h3e218aee, 32'hbe1d66f0} /* (29, 31, 20) {real, imag} */,
  {32'h3de37cec, 32'h3e746b4a} /* (29, 31, 19) {real, imag} */,
  {32'h3e8d20a3, 32'h3ebc3204} /* (29, 31, 18) {real, imag} */,
  {32'h3de8306e, 32'hbdb09a0e} /* (29, 31, 17) {real, imag} */,
  {32'hbe6a626f, 32'h3e90d995} /* (29, 31, 16) {real, imag} */,
  {32'h3d23cfd8, 32'hbd0d225c} /* (29, 31, 15) {real, imag} */,
  {32'hbf0de0e5, 32'hbe341b40} /* (29, 31, 14) {real, imag} */,
  {32'h3ebf87fc, 32'hbdb9c239} /* (29, 31, 13) {real, imag} */,
  {32'hbe35c04e, 32'hbe327d7b} /* (29, 31, 12) {real, imag} */,
  {32'hbe1a43f6, 32'hbf32db66} /* (29, 31, 11) {real, imag} */,
  {32'h3eb5fd69, 32'h3e6b686f} /* (29, 31, 10) {real, imag} */,
  {32'h3e1f221c, 32'h3dbc9a68} /* (29, 31, 9) {real, imag} */,
  {32'h3de0bee0, 32'hbf4062bd} /* (29, 31, 8) {real, imag} */,
  {32'h3ced8b00, 32'h3fba28f8} /* (29, 31, 7) {real, imag} */,
  {32'hbf166796, 32'hbdfde660} /* (29, 31, 6) {real, imag} */,
  {32'hc069e5bc, 32'hbfb4c304} /* (29, 31, 5) {real, imag} */,
  {32'h3fc5a46a, 32'hc0000d1f} /* (29, 31, 4) {real, imag} */,
  {32'hbe34d694, 32'h3f06f9a0} /* (29, 31, 3) {real, imag} */,
  {32'hc10976e2, 32'hbdf29c18} /* (29, 31, 2) {real, imag} */,
  {32'h41a0b567, 32'h40c716e8} /* (29, 31, 1) {real, imag} */,
  {32'h418e6846, 32'hc03994f4} /* (29, 31, 0) {real, imag} */,
  {32'hc164ca54, 32'hc083ee06} /* (29, 30, 31) {real, imag} */,
  {32'h4108fdd2, 32'h401f5e9c} /* (29, 30, 30) {real, imag} */,
  {32'hbf3d1c38, 32'h3f23899d} /* (29, 30, 29) {real, imag} */,
  {32'hbfe3036c, 32'h3ef5a0d6} /* (29, 30, 28) {real, imag} */,
  {32'h3f9b7092, 32'hbebf1c97} /* (29, 30, 27) {real, imag} */,
  {32'h3d0e2640, 32'hbef25786} /* (29, 30, 26) {real, imag} */,
  {32'h3ed4c7f0, 32'h3e9d8360} /* (29, 30, 25) {real, imag} */,
  {32'hbe2d2634, 32'hbe8bf4a1} /* (29, 30, 24) {real, imag} */,
  {32'h3ee98acd, 32'hbe22cc1f} /* (29, 30, 23) {real, imag} */,
  {32'hbf001f2f, 32'hbf0c7bd0} /* (29, 30, 22) {real, imag} */,
  {32'h3ed28e85, 32'hbea6298e} /* (29, 30, 21) {real, imag} */,
  {32'h3d67d760, 32'hbeabaf6c} /* (29, 30, 20) {real, imag} */,
  {32'h3e17fee6, 32'h3efc5bf3} /* (29, 30, 19) {real, imag} */,
  {32'h3df1c924, 32'hbe58a92f} /* (29, 30, 18) {real, imag} */,
  {32'hbe1ed663, 32'h3e6248c8} /* (29, 30, 17) {real, imag} */,
  {32'h3e561933, 32'h3e5684e9} /* (29, 30, 16) {real, imag} */,
  {32'hbd1e136e, 32'hbe503fb5} /* (29, 30, 15) {real, imag} */,
  {32'h3e87b257, 32'h3bf42080} /* (29, 30, 14) {real, imag} */,
  {32'hbdb966c4, 32'h3eb68f86} /* (29, 30, 13) {real, imag} */,
  {32'hbf0e3ab9, 32'hbee1cc11} /* (29, 30, 12) {real, imag} */,
  {32'h3ebaccce, 32'h3eb2d43e} /* (29, 30, 11) {real, imag} */,
  {32'h3ea2f6ad, 32'hbf1941f3} /* (29, 30, 10) {real, imag} */,
  {32'hbe6dcd34, 32'h3dba5248} /* (29, 30, 9) {real, imag} */,
  {32'h3f99f172, 32'h3f2b32ee} /* (29, 30, 8) {real, imag} */,
  {32'hbda7b968, 32'hbf73f13f} /* (29, 30, 7) {real, imag} */,
  {32'h3e8ebeba, 32'hbe9c4232} /* (29, 30, 6) {real, imag} */,
  {32'h3fcbd6e6, 32'h3f4d27c1} /* (29, 30, 5) {real, imag} */,
  {32'hbf8df8e2, 32'hc01fef6e} /* (29, 30, 4) {real, imag} */,
  {32'h3e7bede4, 32'h3ed50b5a} /* (29, 30, 3) {real, imag} */,
  {32'h414cf7ac, 32'h40903bce} /* (29, 30, 2) {real, imag} */,
  {32'hc1b5e489, 32'h3f480b8a} /* (29, 30, 1) {real, imag} */,
  {32'hc13e597d, 32'h3fe894af} /* (29, 30, 0) {real, imag} */,
  {32'h400333fa, 32'hc0713afc} /* (29, 29, 31) {real, imag} */,
  {32'hbdc5ee4c, 32'h401b7f9e} /* (29, 29, 30) {real, imag} */,
  {32'h3f003b05, 32'hbee188aa} /* (29, 29, 29) {real, imag} */,
  {32'hbec2324c, 32'hbf7b9454} /* (29, 29, 28) {real, imag} */,
  {32'hbc547b00, 32'hbe02952c} /* (29, 29, 27) {real, imag} */,
  {32'hbf4935f0, 32'h3f253013} /* (29, 29, 26) {real, imag} */,
  {32'h3f5a5811, 32'hbe1c433c} /* (29, 29, 25) {real, imag} */,
  {32'hbe0a70d2, 32'h3c8cb730} /* (29, 29, 24) {real, imag} */,
  {32'h3e5c5bac, 32'h3d03dc8a} /* (29, 29, 23) {real, imag} */,
  {32'h3dea5ab8, 32'h3e401e90} /* (29, 29, 22) {real, imag} */,
  {32'hbd52d808, 32'h3ce89cf0} /* (29, 29, 21) {real, imag} */,
  {32'h3eb6dc91, 32'hbf013486} /* (29, 29, 20) {real, imag} */,
  {32'h3e55aaa8, 32'h3da87e92} /* (29, 29, 19) {real, imag} */,
  {32'h3d6a1162, 32'hbe316024} /* (29, 29, 18) {real, imag} */,
  {32'h3e3cc4aa, 32'h3e8420a1} /* (29, 29, 17) {real, imag} */,
  {32'hbdb9534a, 32'h3dd8d5d9} /* (29, 29, 16) {real, imag} */,
  {32'h3d807b5c, 32'hbdc77155} /* (29, 29, 15) {real, imag} */,
  {32'hbe14c728, 32'h3b194f20} /* (29, 29, 14) {real, imag} */,
  {32'hbeb35c07, 32'hbe861542} /* (29, 29, 13) {real, imag} */,
  {32'h3e2cb71a, 32'hbeb36d6a} /* (29, 29, 12) {real, imag} */,
  {32'hbf6f964a, 32'hbd334a00} /* (29, 29, 11) {real, imag} */,
  {32'h3e37213a, 32'h3ccccad8} /* (29, 29, 10) {real, imag} */,
  {32'h3e92f84d, 32'hbd57fa70} /* (29, 29, 9) {real, imag} */,
  {32'hbecbbb9a, 32'h3f35f5b2} /* (29, 29, 8) {real, imag} */,
  {32'hbe843f86, 32'hbe9607ae} /* (29, 29, 7) {real, imag} */,
  {32'hbe311c4a, 32'hbe843564} /* (29, 29, 6) {real, imag} */,
  {32'hbe3b6a7c, 32'h3f9dc348} /* (29, 29, 5) {real, imag} */,
  {32'h3efd76fd, 32'hbf646c6a} /* (29, 29, 4) {real, imag} */,
  {32'h3d9a5a4c, 32'hbefa681b} /* (29, 29, 3) {real, imag} */,
  {32'h4005dcc3, 32'h401d31b6} /* (29, 29, 2) {real, imag} */,
  {32'hc0754d4c, 32'hc01403bf} /* (29, 29, 1) {real, imag} */,
  {32'h3e839992, 32'h3d112a38} /* (29, 29, 0) {real, imag} */,
  {32'h40a04205, 32'hc00c80a3} /* (29, 28, 31) {real, imag} */,
  {32'hbf92ba78, 32'h3ffea0c2} /* (29, 28, 30) {real, imag} */,
  {32'h3e76001b, 32'h3e349028} /* (29, 28, 29) {real, imag} */,
  {32'h3f4d952e, 32'hbecac78e} /* (29, 28, 28) {real, imag} */,
  {32'h3d27d09a, 32'h3f582390} /* (29, 28, 27) {real, imag} */,
  {32'hbdcdb624, 32'hbec7aaed} /* (29, 28, 26) {real, imag} */,
  {32'h3e8d7a3c, 32'h3eb88083} /* (29, 28, 25) {real, imag} */,
  {32'hbe9b468f, 32'h3ebe9f39} /* (29, 28, 24) {real, imag} */,
  {32'h3e40acc6, 32'h3efff297} /* (29, 28, 23) {real, imag} */,
  {32'hbd68f344, 32'hbe9e8616} /* (29, 28, 22) {real, imag} */,
  {32'h3da0e28b, 32'hbee666ec} /* (29, 28, 21) {real, imag} */,
  {32'hbead7468, 32'h3ea3988c} /* (29, 28, 20) {real, imag} */,
  {32'h3e301119, 32'h3ef8d3d8} /* (29, 28, 19) {real, imag} */,
  {32'hbe1c403e, 32'hbdfcb684} /* (29, 28, 18) {real, imag} */,
  {32'hbea14475, 32'h3c81c6e8} /* (29, 28, 17) {real, imag} */,
  {32'hbe228a79, 32'h3d175a39} /* (29, 28, 16) {real, imag} */,
  {32'h3eadada3, 32'h3cf2dfa8} /* (29, 28, 15) {real, imag} */,
  {32'hbf3b638d, 32'h3dd35941} /* (29, 28, 14) {real, imag} */,
  {32'h3e80ccfc, 32'h3eb86b56} /* (29, 28, 13) {real, imag} */,
  {32'hbe096b6e, 32'h3e855abe} /* (29, 28, 12) {real, imag} */,
  {32'h3d77d138, 32'h3e5ed278} /* (29, 28, 11) {real, imag} */,
  {32'h3daa60fc, 32'h3e3751f0} /* (29, 28, 10) {real, imag} */,
  {32'hbf021620, 32'h3f1be7ae} /* (29, 28, 9) {real, imag} */,
  {32'hbec31488, 32'hbcdd0a88} /* (29, 28, 8) {real, imag} */,
  {32'hbe6ea136, 32'hbc7c1050} /* (29, 28, 7) {real, imag} */,
  {32'h3e352336, 32'hbec5bc19} /* (29, 28, 6) {real, imag} */,
  {32'hbfe983fa, 32'hbf25379e} /* (29, 28, 5) {real, imag} */,
  {32'h3f8c07fc, 32'h3db6ad34} /* (29, 28, 4) {real, imag} */,
  {32'hbf89de3a, 32'hbfee653c} /* (29, 28, 3) {real, imag} */,
  {32'hc019d5af, 32'h3f7d2350} /* (29, 28, 2) {real, imag} */,
  {32'h402757d7, 32'hc01cd0ce} /* (29, 28, 1) {real, imag} */,
  {32'h3fd3fc1a, 32'hbf871e66} /* (29, 28, 0) {real, imag} */,
  {32'hc011ac68, 32'h3fde705c} /* (29, 27, 31) {real, imag} */,
  {32'h3fa46168, 32'h3c94cae0} /* (29, 27, 30) {real, imag} */,
  {32'h3e4611ae, 32'h3ec938be} /* (29, 27, 29) {real, imag} */,
  {32'hbefe69bd, 32'h3e838b41} /* (29, 27, 28) {real, imag} */,
  {32'hbce208c0, 32'hbf97000c} /* (29, 27, 27) {real, imag} */,
  {32'hbe321746, 32'h3ebccb46} /* (29, 27, 26) {real, imag} */,
  {32'h3e2ea345, 32'hbdc49fa8} /* (29, 27, 25) {real, imag} */,
  {32'h3e5950e5, 32'hbcf51580} /* (29, 27, 24) {real, imag} */,
  {32'hbd912d60, 32'hbd13a558} /* (29, 27, 23) {real, imag} */,
  {32'hbf06ab3e, 32'h3e54db47} /* (29, 27, 22) {real, imag} */,
  {32'h3d8a1da1, 32'h3e5ddeef} /* (29, 27, 21) {real, imag} */,
  {32'h3d92dcda, 32'h3c2b1660} /* (29, 27, 20) {real, imag} */,
  {32'hbe33532a, 32'h3de486fe} /* (29, 27, 19) {real, imag} */,
  {32'h3d86e269, 32'h3e238b44} /* (29, 27, 18) {real, imag} */,
  {32'hbd6742d0, 32'hbe1da836} /* (29, 27, 17) {real, imag} */,
  {32'h3db405a2, 32'h3e223b46} /* (29, 27, 16) {real, imag} */,
  {32'h3e35f004, 32'hbe1008ce} /* (29, 27, 15) {real, imag} */,
  {32'h3dd646e2, 32'hbd8d6d65} /* (29, 27, 14) {real, imag} */,
  {32'h3e5bbbea, 32'hbc722748} /* (29, 27, 13) {real, imag} */,
  {32'hbdda8138, 32'hbe365176} /* (29, 27, 12) {real, imag} */,
  {32'h3f1ed5c1, 32'h3dc07660} /* (29, 27, 11) {real, imag} */,
  {32'h3de93fec, 32'hbf4e8117} /* (29, 27, 10) {real, imag} */,
  {32'hbe6b3758, 32'h3e8f080e} /* (29, 27, 9) {real, imag} */,
  {32'hbe59e0a2, 32'hbbd9dd10} /* (29, 27, 8) {real, imag} */,
  {32'hbf1da539, 32'hbea1be85} /* (29, 27, 7) {real, imag} */,
  {32'h3e346253, 32'h3eff8d9c} /* (29, 27, 6) {real, imag} */,
  {32'h3f94df07, 32'hbeb15bc9} /* (29, 27, 5) {real, imag} */,
  {32'hbf2b6320, 32'hbee612d7} /* (29, 27, 4) {real, imag} */,
  {32'h3ed74e96, 32'h3f3ddeb1} /* (29, 27, 3) {real, imag} */,
  {32'h3e65522e, 32'h3f581c36} /* (29, 27, 2) {real, imag} */,
  {32'hc05a22bc, 32'h3f1b92e9} /* (29, 27, 1) {real, imag} */,
  {32'hbff9715a, 32'h3f86368c} /* (29, 27, 0) {real, imag} */,
  {32'hbf580c40, 32'hbede2120} /* (29, 26, 31) {real, imag} */,
  {32'hb920a800, 32'h3da5bc9c} /* (29, 26, 30) {real, imag} */,
  {32'h3e0fcf25, 32'h3b4405c0} /* (29, 26, 29) {real, imag} */,
  {32'h3f024f82, 32'h3e4bf979} /* (29, 26, 28) {real, imag} */,
  {32'h3e7182c8, 32'hbd741818} /* (29, 26, 27) {real, imag} */,
  {32'hbc0aae40, 32'hbdf0b19c} /* (29, 26, 26) {real, imag} */,
  {32'h3f43cc15, 32'hbeaf472b} /* (29, 26, 25) {real, imag} */,
  {32'h3d6a60de, 32'hbdee0e0c} /* (29, 26, 24) {real, imag} */,
  {32'h3e0476ac, 32'hbe00ba64} /* (29, 26, 23) {real, imag} */,
  {32'h3e47ee34, 32'h3df9e334} /* (29, 26, 22) {real, imag} */,
  {32'h3d68176c, 32'hbf026d5e} /* (29, 26, 21) {real, imag} */,
  {32'h3ee00a5e, 32'hbeeb9e9c} /* (29, 26, 20) {real, imag} */,
  {32'h3ed92c34, 32'hbe7c256f} /* (29, 26, 19) {real, imag} */,
  {32'hbf080b34, 32'hbe635262} /* (29, 26, 18) {real, imag} */,
  {32'hbeb061fd, 32'h3e8a2db6} /* (29, 26, 17) {real, imag} */,
  {32'h3d23ecf0, 32'hbe807e58} /* (29, 26, 16) {real, imag} */,
  {32'hbe83dbce, 32'hbe6069c6} /* (29, 26, 15) {real, imag} */,
  {32'h3ec33878, 32'hbe199570} /* (29, 26, 14) {real, imag} */,
  {32'h3eba5d3a, 32'h3f4160c0} /* (29, 26, 13) {real, imag} */,
  {32'hbd6aee8c, 32'h3e295d83} /* (29, 26, 12) {real, imag} */,
  {32'hbf17e075, 32'h3e9f4a16} /* (29, 26, 11) {real, imag} */,
  {32'hbe8d7024, 32'hbe2ee5ef} /* (29, 26, 10) {real, imag} */,
  {32'h3f0e5da6, 32'h3e72fce8} /* (29, 26, 9) {real, imag} */,
  {32'hbe946fa1, 32'hbf5fc1da} /* (29, 26, 8) {real, imag} */,
  {32'h3edd6bcc, 32'hbf6f1faa} /* (29, 26, 7) {real, imag} */,
  {32'hbebce9f8, 32'h3de5b973} /* (29, 26, 6) {real, imag} */,
  {32'hbf87fe74, 32'hbdefb05f} /* (29, 26, 5) {real, imag} */,
  {32'hbdc20a48, 32'h3f32fc21} /* (29, 26, 4) {real, imag} */,
  {32'h3b3bb3a0, 32'hbd06d348} /* (29, 26, 3) {real, imag} */,
  {32'h3f00d86e, 32'hbf22ee15} /* (29, 26, 2) {real, imag} */,
  {32'h3ede14bc, 32'hbf4a7d0e} /* (29, 26, 1) {real, imag} */,
  {32'h3e9ef882, 32'hbeb8a253} /* (29, 26, 0) {real, imag} */,
  {32'h3fb7f53c, 32'hbd291360} /* (29, 25, 31) {real, imag} */,
  {32'h3ec08744, 32'h3e715334} /* (29, 25, 30) {real, imag} */,
  {32'hbf3fa8c2, 32'h3eb6ea50} /* (29, 25, 29) {real, imag} */,
  {32'h3ccacd60, 32'h3e0a06cd} /* (29, 25, 28) {real, imag} */,
  {32'h3e0c9a26, 32'h3f592f99} /* (29, 25, 27) {real, imag} */,
  {32'h3f4d13f4, 32'h3ee7a1ca} /* (29, 25, 26) {real, imag} */,
  {32'hbde95e04, 32'h3eaa0862} /* (29, 25, 25) {real, imag} */,
  {32'hbe2d8f49, 32'h3dd4b929} /* (29, 25, 24) {real, imag} */,
  {32'h3ec6f770, 32'hbece263c} /* (29, 25, 23) {real, imag} */,
  {32'hbe80e071, 32'h3de4a56b} /* (29, 25, 22) {real, imag} */,
  {32'hbe8b6491, 32'hbf022dce} /* (29, 25, 21) {real, imag} */,
  {32'h3e0b8dea, 32'h3d5e3984} /* (29, 25, 20) {real, imag} */,
  {32'hbee84bb8, 32'hbdecff98} /* (29, 25, 19) {real, imag} */,
  {32'hbd2ad8a4, 32'h3e44e83c} /* (29, 25, 18) {real, imag} */,
  {32'hbc37fe10, 32'h3d97c0e0} /* (29, 25, 17) {real, imag} */,
  {32'h3dbb379a, 32'h3e86b1d8} /* (29, 25, 16) {real, imag} */,
  {32'hbf013f4c, 32'h3ea64641} /* (29, 25, 15) {real, imag} */,
  {32'h3ea7c3a6, 32'hbe0110bc} /* (29, 25, 14) {real, imag} */,
  {32'h3ea60a35, 32'hbe3efc9a} /* (29, 25, 13) {real, imag} */,
  {32'h3e7e2e4d, 32'hbc891f00} /* (29, 25, 12) {real, imag} */,
  {32'hbdf2c9fc, 32'hbeaa4c4f} /* (29, 25, 11) {real, imag} */,
  {32'hbe4eef20, 32'hbf28d10e} /* (29, 25, 10) {real, imag} */,
  {32'h3afd6300, 32'h3eaa06d7} /* (29, 25, 9) {real, imag} */,
  {32'hbc88042a, 32'h3e38d04b} /* (29, 25, 8) {real, imag} */,
  {32'hbefdf12b, 32'hbe5aeb8b} /* (29, 25, 7) {real, imag} */,
  {32'hbe39af4a, 32'hbabe1700} /* (29, 25, 6) {real, imag} */,
  {32'h3ea85846, 32'hbf30d7c9} /* (29, 25, 5) {real, imag} */,
  {32'hbf21fc78, 32'h3e34d244} /* (29, 25, 4) {real, imag} */,
  {32'hbea2feaf, 32'hbd27a23c} /* (29, 25, 3) {real, imag} */,
  {32'hbf138f1c, 32'hbf5c0515} /* (29, 25, 2) {real, imag} */,
  {32'hbde7bc7e, 32'h3e8ce8fa} /* (29, 25, 1) {real, imag} */,
  {32'h3f9315c2, 32'h3dd5a24c} /* (29, 25, 0) {real, imag} */,
  {32'hbf0c2148, 32'h3faca212} /* (29, 24, 31) {real, imag} */,
  {32'hbe2afe14, 32'h3ee3f56f} /* (29, 24, 30) {real, imag} */,
  {32'h3f5554d8, 32'hbf22e601} /* (29, 24, 29) {real, imag} */,
  {32'hbe3e2ea7, 32'h3e87af7c} /* (29, 24, 28) {real, imag} */,
  {32'h3e8896a8, 32'hbef5af81} /* (29, 24, 27) {real, imag} */,
  {32'hbebd9f33, 32'hbeecfabc} /* (29, 24, 26) {real, imag} */,
  {32'hbeef64fa, 32'hbd940df7} /* (29, 24, 25) {real, imag} */,
  {32'h3df3bfb0, 32'hbe3aa950} /* (29, 24, 24) {real, imag} */,
  {32'hbe99ed08, 32'h3e75475e} /* (29, 24, 23) {real, imag} */,
  {32'h3e9fbc46, 32'h3eaf67fa} /* (29, 24, 22) {real, imag} */,
  {32'hbc8bec78, 32'hbf52b48e} /* (29, 24, 21) {real, imag} */,
  {32'hbde07c02, 32'hbe6b9c1a} /* (29, 24, 20) {real, imag} */,
  {32'h3f3cf1e7, 32'hbe0f413a} /* (29, 24, 19) {real, imag} */,
  {32'hbcd52eb0, 32'h3e82907d} /* (29, 24, 18) {real, imag} */,
  {32'h3e863393, 32'hbbcd4fc0} /* (29, 24, 17) {real, imag} */,
  {32'h3e9d3ae3, 32'hbe6db3e6} /* (29, 24, 16) {real, imag} */,
  {32'hbb96f480, 32'hbde86fa6} /* (29, 24, 15) {real, imag} */,
  {32'h3ed324bd, 32'h3edadac9} /* (29, 24, 14) {real, imag} */,
  {32'hbeb528bb, 32'hbe010c29} /* (29, 24, 13) {real, imag} */,
  {32'hbe7d21e6, 32'h3e607c79} /* (29, 24, 12) {real, imag} */,
  {32'h3ef8ce4c, 32'hbee47cee} /* (29, 24, 11) {real, imag} */,
  {32'h3f2f30de, 32'h3ea20684} /* (29, 24, 10) {real, imag} */,
  {32'hbe678150, 32'h3d8e0fab} /* (29, 24, 9) {real, imag} */,
  {32'h3d140f90, 32'hbd1534b0} /* (29, 24, 8) {real, imag} */,
  {32'hbead3a13, 32'h3f3215bc} /* (29, 24, 7) {real, imag} */,
  {32'h3ec51a58, 32'h3e81e3a0} /* (29, 24, 6) {real, imag} */,
  {32'hbeebd34d, 32'h3e054d50} /* (29, 24, 5) {real, imag} */,
  {32'h3e9dc24c, 32'h3e62ce16} /* (29, 24, 4) {real, imag} */,
  {32'hbd555d70, 32'h3f3ddbb4} /* (29, 24, 3) {real, imag} */,
  {32'h3f544fbc, 32'hbf1a93fd} /* (29, 24, 2) {real, imag} */,
  {32'hbff3bd9a, 32'h3fa6fe51} /* (29, 24, 1) {real, imag} */,
  {32'hbf066be3, 32'h3e6cc587} /* (29, 24, 0) {real, imag} */,
  {32'h3f4e3aae, 32'h3da618c0} /* (29, 23, 31) {real, imag} */,
  {32'hbf402127, 32'h3f034bcc} /* (29, 23, 30) {real, imag} */,
  {32'hbec8c264, 32'hbdbee9ba} /* (29, 23, 29) {real, imag} */,
  {32'h3d36dd06, 32'h3d49c147} /* (29, 23, 28) {real, imag} */,
  {32'h3e1fd260, 32'hbf4d0b14} /* (29, 23, 27) {real, imag} */,
  {32'h3e6d125e, 32'h3d322ba9} /* (29, 23, 26) {real, imag} */,
  {32'hbde05c1a, 32'h3e7a94a6} /* (29, 23, 25) {real, imag} */,
  {32'h3ee32176, 32'h3e607702} /* (29, 23, 24) {real, imag} */,
  {32'hbe8b4b9e, 32'h3b2d58c0} /* (29, 23, 23) {real, imag} */,
  {32'hbf3aa175, 32'hbdd6bba8} /* (29, 23, 22) {real, imag} */,
  {32'h3bba46b0, 32'h3e5a6d4f} /* (29, 23, 21) {real, imag} */,
  {32'h3e9cbcc0, 32'hbea104bd} /* (29, 23, 20) {real, imag} */,
  {32'hbede9694, 32'hbf054fae} /* (29, 23, 19) {real, imag} */,
  {32'hbe6d99bb, 32'hbf085a56} /* (29, 23, 18) {real, imag} */,
  {32'hbdee75a7, 32'hbe59ecc3} /* (29, 23, 17) {real, imag} */,
  {32'h3edf7688, 32'h3e7ac36d} /* (29, 23, 16) {real, imag} */,
  {32'hbe8b350c, 32'h3e87cac0} /* (29, 23, 15) {real, imag} */,
  {32'h3ec9cf49, 32'hbe2e3d66} /* (29, 23, 14) {real, imag} */,
  {32'h3ed3fefe, 32'hbf2b96ae} /* (29, 23, 13) {real, imag} */,
  {32'hbe579ffe, 32'h3f0e8cc6} /* (29, 23, 12) {real, imag} */,
  {32'hbecf2d0e, 32'h3e89a696} /* (29, 23, 11) {real, imag} */,
  {32'hbf704259, 32'h3ebd588e} /* (29, 23, 10) {real, imag} */,
  {32'hbe553f06, 32'hbed5ebef} /* (29, 23, 9) {real, imag} */,
  {32'h3e03e961, 32'h3e8b2d18} /* (29, 23, 8) {real, imag} */,
  {32'hbeb92f02, 32'hbddce680} /* (29, 23, 7) {real, imag} */,
  {32'hbdaa9e82, 32'hbeddbb75} /* (29, 23, 6) {real, imag} */,
  {32'hbed1f940, 32'hbe14e59e} /* (29, 23, 5) {real, imag} */,
  {32'hbce141d8, 32'hbf6fc942} /* (29, 23, 4) {real, imag} */,
  {32'h3e80e1f9, 32'h3b9a2040} /* (29, 23, 3) {real, imag} */,
  {32'h3f700e87, 32'h3dfb6408} /* (29, 23, 2) {real, imag} */,
  {32'hbf9d4b78, 32'hbeafedfd} /* (29, 23, 1) {real, imag} */,
  {32'hbedb22aa, 32'h3f133602} /* (29, 23, 0) {real, imag} */,
  {32'h3cf4b9b0, 32'h3d7ec1f8} /* (29, 22, 31) {real, imag} */,
  {32'h3d7663b8, 32'hbdedcbda} /* (29, 22, 30) {real, imag} */,
  {32'hbf28222c, 32'h3d082e0e} /* (29, 22, 29) {real, imag} */,
  {32'hbf25fbab, 32'h3f0ca5de} /* (29, 22, 28) {real, imag} */,
  {32'hbea42e18, 32'hbd8cda36} /* (29, 22, 27) {real, imag} */,
  {32'h3e965c5e, 32'h3ecad827} /* (29, 22, 26) {real, imag} */,
  {32'h3ec935dc, 32'h3ed38068} /* (29, 22, 25) {real, imag} */,
  {32'hbe598cdb, 32'hbe8b345d} /* (29, 22, 24) {real, imag} */,
  {32'hbe8ad5a8, 32'hbdfea94f} /* (29, 22, 23) {real, imag} */,
  {32'h3e096bcc, 32'hbeb8ed01} /* (29, 22, 22) {real, imag} */,
  {32'h3efb1dd4, 32'hbe06643c} /* (29, 22, 21) {real, imag} */,
  {32'h3e2c7e6a, 32'hbefc905a} /* (29, 22, 20) {real, imag} */,
  {32'hbf1a7738, 32'hbdb57cd4} /* (29, 22, 19) {real, imag} */,
  {32'h3f2c238a, 32'h3c86ee38} /* (29, 22, 18) {real, imag} */,
  {32'h3ef0d46d, 32'h3e5c259e} /* (29, 22, 17) {real, imag} */,
  {32'hbecfa086, 32'hbe53c999} /* (29, 22, 16) {real, imag} */,
  {32'h3c6dba88, 32'hbdfe5fa2} /* (29, 22, 15) {real, imag} */,
  {32'h3d8a3a04, 32'hbe5e0e08} /* (29, 22, 14) {real, imag} */,
  {32'h3e80663a, 32'h3ecd31a0} /* (29, 22, 13) {real, imag} */,
  {32'h3ea5c536, 32'h3e951ed2} /* (29, 22, 12) {real, imag} */,
  {32'h3e0d77a2, 32'h3e77c95c} /* (29, 22, 11) {real, imag} */,
  {32'h3d86baee, 32'hbf2bb94a} /* (29, 22, 10) {real, imag} */,
  {32'hbef49658, 32'hbe399fe2} /* (29, 22, 9) {real, imag} */,
  {32'hbdcc0f8a, 32'h3f31cc43} /* (29, 22, 8) {real, imag} */,
  {32'h3e8fb50b, 32'hbe947ef8} /* (29, 22, 7) {real, imag} */,
  {32'h3e0dd4ca, 32'h3ee1c73e} /* (29, 22, 6) {real, imag} */,
  {32'h3f02ceb2, 32'h3ed45c67} /* (29, 22, 5) {real, imag} */,
  {32'h3dbd040a, 32'hbccf1120} /* (29, 22, 4) {real, imag} */,
  {32'h3e9fd5c0, 32'hbec31c44} /* (29, 22, 3) {real, imag} */,
  {32'h3e08d53f, 32'h3e8a0253} /* (29, 22, 2) {real, imag} */,
  {32'h3f093280, 32'hbe6251be} /* (29, 22, 1) {real, imag} */,
  {32'hbf040ff1, 32'hbe42fdb9} /* (29, 22, 0) {real, imag} */,
  {32'hbdad1db6, 32'h3f68f050} /* (29, 21, 31) {real, imag} */,
  {32'hbe0ca481, 32'hbf81279d} /* (29, 21, 30) {real, imag} */,
  {32'hbdb1742e, 32'hbe25b40a} /* (29, 21, 29) {real, imag} */,
  {32'hbefe4fe0, 32'hbf0673a6} /* (29, 21, 28) {real, imag} */,
  {32'hbe90ef5f, 32'hbf0a923c} /* (29, 21, 27) {real, imag} */,
  {32'hbeea89be, 32'hbedf8912} /* (29, 21, 26) {real, imag} */,
  {32'hbd314d3e, 32'hbe32f829} /* (29, 21, 25) {real, imag} */,
  {32'h3e2e3a98, 32'hbeafe429} /* (29, 21, 24) {real, imag} */,
  {32'h3f4d18fc, 32'hbda2d232} /* (29, 21, 23) {real, imag} */,
  {32'h3f0d3517, 32'h3db5bba6} /* (29, 21, 22) {real, imag} */,
  {32'hbe79ada9, 32'h3d8e350a} /* (29, 21, 21) {real, imag} */,
  {32'h3e709d21, 32'h3e64a33d} /* (29, 21, 20) {real, imag} */,
  {32'hbe94815e, 32'h3db09f50} /* (29, 21, 19) {real, imag} */,
  {32'hbdd38ea9, 32'h3f010ee0} /* (29, 21, 18) {real, imag} */,
  {32'hbf0a0f4c, 32'hbe1d8042} /* (29, 21, 17) {real, imag} */,
  {32'hbe274d4e, 32'h3dc7046c} /* (29, 21, 16) {real, imag} */,
  {32'h3cb4fd70, 32'hbe268cac} /* (29, 21, 15) {real, imag} */,
  {32'hbeb5e27a, 32'h3e9b7e1e} /* (29, 21, 14) {real, imag} */,
  {32'h3ee1e42e, 32'h3c968420} /* (29, 21, 13) {real, imag} */,
  {32'h3e815a29, 32'h3e7cdc92} /* (29, 21, 12) {real, imag} */,
  {32'h3e871699, 32'h3f08a7f0} /* (29, 21, 11) {real, imag} */,
  {32'hbf302278, 32'hbe51fb2a} /* (29, 21, 10) {real, imag} */,
  {32'hbe3b9e5e, 32'hbe9154d4} /* (29, 21, 9) {real, imag} */,
  {32'hbe998ce8, 32'h3dd8c814} /* (29, 21, 8) {real, imag} */,
  {32'h3ec08d4c, 32'hbe457db5} /* (29, 21, 7) {real, imag} */,
  {32'hbec0c734, 32'hbe9f8e09} /* (29, 21, 6) {real, imag} */,
  {32'h3d8de658, 32'h3f00de65} /* (29, 21, 5) {real, imag} */,
  {32'h3edfd46e, 32'hbdb78fbf} /* (29, 21, 4) {real, imag} */,
  {32'h3eb57124, 32'h3dad3ed4} /* (29, 21, 3) {real, imag} */,
  {32'h3e01b80b, 32'hbed5cd53} /* (29, 21, 2) {real, imag} */,
  {32'hbe71669e, 32'h3eb7be2a} /* (29, 21, 1) {real, imag} */,
  {32'hbf48c8d5, 32'h3f6190a6} /* (29, 21, 0) {real, imag} */,
  {32'h3e047005, 32'h3d89a964} /* (29, 20, 31) {real, imag} */,
  {32'hbf167eae, 32'h3c968e10} /* (29, 20, 30) {real, imag} */,
  {32'h3d81bb26, 32'hbe19f5d0} /* (29, 20, 29) {real, imag} */,
  {32'hbdc6f93c, 32'h3ebbc80d} /* (29, 20, 28) {real, imag} */,
  {32'h3c3310d8, 32'hbe810fb9} /* (29, 20, 27) {real, imag} */,
  {32'h3e1ad192, 32'h3d7c850e} /* (29, 20, 26) {real, imag} */,
  {32'hbeac6ea6, 32'h3eb6ffd2} /* (29, 20, 25) {real, imag} */,
  {32'hbf1d60be, 32'hbd2f4ba0} /* (29, 20, 24) {real, imag} */,
  {32'h3e199126, 32'h3d8b8296} /* (29, 20, 23) {real, imag} */,
  {32'hbed48e53, 32'hbd859a5c} /* (29, 20, 22) {real, imag} */,
  {32'h3ea1d2d3, 32'h3f05c4bf} /* (29, 20, 21) {real, imag} */,
  {32'hbe113716, 32'hbee658ad} /* (29, 20, 20) {real, imag} */,
  {32'h3e332ed5, 32'h3e7687fc} /* (29, 20, 19) {real, imag} */,
  {32'hbe87228e, 32'h3e1da82e} /* (29, 20, 18) {real, imag} */,
  {32'h3e1fb6de, 32'hbdc34418} /* (29, 20, 17) {real, imag} */,
  {32'hbe20e8e4, 32'hbc3c7b30} /* (29, 20, 16) {real, imag} */,
  {32'hbd71b190, 32'h3d690a0c} /* (29, 20, 15) {real, imag} */,
  {32'h3e7f429a, 32'hbe6ea53f} /* (29, 20, 14) {real, imag} */,
  {32'h3ca2587f, 32'hbe658bcc} /* (29, 20, 13) {real, imag} */,
  {32'h3ddaa03d, 32'hbe6c6b61} /* (29, 20, 12) {real, imag} */,
  {32'hbec51336, 32'hbeb1647c} /* (29, 20, 11) {real, imag} */,
  {32'hbe0abd26, 32'h3f1835cc} /* (29, 20, 10) {real, imag} */,
  {32'hbf0be8cd, 32'h3d57e876} /* (29, 20, 9) {real, imag} */,
  {32'h3daa7c00, 32'hbde8fc05} /* (29, 20, 8) {real, imag} */,
  {32'hbe758c0c, 32'h3ec1bfd4} /* (29, 20, 7) {real, imag} */,
  {32'h3dcdbab0, 32'hbe896148} /* (29, 20, 6) {real, imag} */,
  {32'h3d37ef96, 32'h3ead2b92} /* (29, 20, 5) {real, imag} */,
  {32'h3f397dd8, 32'h3cbfae98} /* (29, 20, 4) {real, imag} */,
  {32'hbe1eff65, 32'hbf041617} /* (29, 20, 3) {real, imag} */,
  {32'h3e4f02d0, 32'hbe04ae80} /* (29, 20, 2) {real, imag} */,
  {32'h3e6cb2d6, 32'hbea11ae9} /* (29, 20, 1) {real, imag} */,
  {32'hbe056e92, 32'h3e2ffb60} /* (29, 20, 0) {real, imag} */,
  {32'h3e54a2ee, 32'hbe97d557} /* (29, 19, 31) {real, imag} */,
  {32'h3c5770fc, 32'h3f0ba3cd} /* (29, 19, 30) {real, imag} */,
  {32'h3eacb908, 32'h3e5e57a6} /* (29, 19, 29) {real, imag} */,
  {32'h3ea547c9, 32'hbc59a290} /* (29, 19, 28) {real, imag} */,
  {32'hbf0caf56, 32'h3ea6147f} /* (29, 19, 27) {real, imag} */,
  {32'h3e067b7c, 32'hbd51cc44} /* (29, 19, 26) {real, imag} */,
  {32'h3d9b16a4, 32'h3da99531} /* (29, 19, 25) {real, imag} */,
  {32'hbe6ba2e8, 32'hbd124400} /* (29, 19, 24) {real, imag} */,
  {32'hbefe61ae, 32'h3d7ce973} /* (29, 19, 23) {real, imag} */,
  {32'hbe80cf90, 32'hbe29573e} /* (29, 19, 22) {real, imag} */,
  {32'hbdfd5ab4, 32'h3e0848ca} /* (29, 19, 21) {real, imag} */,
  {32'h3e969ef8, 32'h3eb40c84} /* (29, 19, 20) {real, imag} */,
  {32'h3e4973af, 32'h3e44c7bb} /* (29, 19, 19) {real, imag} */,
  {32'h3f049638, 32'h3df1d478} /* (29, 19, 18) {real, imag} */,
  {32'hbd3505dc, 32'hbf254efe} /* (29, 19, 17) {real, imag} */,
  {32'hbd50d4c0, 32'h3de6795e} /* (29, 19, 16) {real, imag} */,
  {32'hbe00ecc7, 32'h3e9a0e5c} /* (29, 19, 15) {real, imag} */,
  {32'hbe71bd1f, 32'h3df28fd4} /* (29, 19, 14) {real, imag} */,
  {32'h3dde8208, 32'h3c406b20} /* (29, 19, 13) {real, imag} */,
  {32'hbd3dbbd4, 32'hbe86436c} /* (29, 19, 12) {real, imag} */,
  {32'h3ee98bfc, 32'hbe9ae316} /* (29, 19, 11) {real, imag} */,
  {32'hbe0feb33, 32'h3eb3276c} /* (29, 19, 10) {real, imag} */,
  {32'h3ec8dc6a, 32'hbf1cab74} /* (29, 19, 9) {real, imag} */,
  {32'h3e387803, 32'h3dff2c93} /* (29, 19, 8) {real, imag} */,
  {32'hbde5fabc, 32'h3e8e6d62} /* (29, 19, 7) {real, imag} */,
  {32'h3f07376e, 32'h3e0685e3} /* (29, 19, 6) {real, imag} */,
  {32'h3dd1b777, 32'hbdbb4199} /* (29, 19, 5) {real, imag} */,
  {32'h3ddb3e8a, 32'h3d8be55c} /* (29, 19, 4) {real, imag} */,
  {32'hbeeaabeb, 32'hbee35331} /* (29, 19, 3) {real, imag} */,
  {32'h3ee358bc, 32'h3e6ed2cc} /* (29, 19, 2) {real, imag} */,
  {32'hbca2fcb0, 32'hbd595910} /* (29, 19, 1) {real, imag} */,
  {32'h3f212d44, 32'hbec45c50} /* (29, 19, 0) {real, imag} */,
  {32'hbe7a2e6d, 32'h3e8707ee} /* (29, 18, 31) {real, imag} */,
  {32'hbd2467bc, 32'hbe7f90b0} /* (29, 18, 30) {real, imag} */,
  {32'hbea32008, 32'hbeb6105d} /* (29, 18, 29) {real, imag} */,
  {32'hbed2f3f5, 32'hbec8d664} /* (29, 18, 28) {real, imag} */,
  {32'hbef24c12, 32'hbe4658ea} /* (29, 18, 27) {real, imag} */,
  {32'h3e2d07bc, 32'hbe72cf76} /* (29, 18, 26) {real, imag} */,
  {32'hbf1ef27f, 32'hbeb63de2} /* (29, 18, 25) {real, imag} */,
  {32'h3e2d8112, 32'h3e2af467} /* (29, 18, 24) {real, imag} */,
  {32'h3f48eb5d, 32'h3f01a58b} /* (29, 18, 23) {real, imag} */,
  {32'hbe560cb1, 32'h3f1a111f} /* (29, 18, 22) {real, imag} */,
  {32'hbe53f290, 32'hbea15912} /* (29, 18, 21) {real, imag} */,
  {32'hbf006a97, 32'h3e805194} /* (29, 18, 20) {real, imag} */,
  {32'h3e9b7695, 32'h3e9f1686} /* (29, 18, 19) {real, imag} */,
  {32'hbe5af0ef, 32'h3e004178} /* (29, 18, 18) {real, imag} */,
  {32'hbd3157b4, 32'h3e79927c} /* (29, 18, 17) {real, imag} */,
  {32'h3e8a6f9c, 32'h3e1b0381} /* (29, 18, 16) {real, imag} */,
  {32'hbd21cfba, 32'hbdfbf516} /* (29, 18, 15) {real, imag} */,
  {32'h3e847f12, 32'h3d3fbe30} /* (29, 18, 14) {real, imag} */,
  {32'hbd32b52e, 32'h3d6e57c8} /* (29, 18, 13) {real, imag} */,
  {32'h3d923474, 32'h3e6cdd78} /* (29, 18, 12) {real, imag} */,
  {32'hbd1302e3, 32'h3f2f83af} /* (29, 18, 11) {real, imag} */,
  {32'h3ea00cc8, 32'h3d434d1a} /* (29, 18, 10) {real, imag} */,
  {32'hbd02a664, 32'h3b3603d0} /* (29, 18, 9) {real, imag} */,
  {32'h3e02645b, 32'h3d04a8a0} /* (29, 18, 8) {real, imag} */,
  {32'hbe368c7a, 32'hbe16c349} /* (29, 18, 7) {real, imag} */,
  {32'hbe874b84, 32'h3eaba979} /* (29, 18, 6) {real, imag} */,
  {32'h3e8dbc0c, 32'hbe9b8340} /* (29, 18, 5) {real, imag} */,
  {32'h3c9bf610, 32'h3d122038} /* (29, 18, 4) {real, imag} */,
  {32'h3e28f0e9, 32'h3f06260c} /* (29, 18, 3) {real, imag} */,
  {32'hbdb16950, 32'h3df46d44} /* (29, 18, 2) {real, imag} */,
  {32'hbe3acb3a, 32'h3e476a52} /* (29, 18, 1) {real, imag} */,
  {32'hbe2a0964, 32'h3ee009d4} /* (29, 18, 0) {real, imag} */,
  {32'h3e2b920e, 32'hbe373a0e} /* (29, 17, 31) {real, imag} */,
  {32'h3d438797, 32'h3dad04a4} /* (29, 17, 30) {real, imag} */,
  {32'h3e482168, 32'h3cfba950} /* (29, 17, 29) {real, imag} */,
  {32'hbd6184d4, 32'h3e705478} /* (29, 17, 28) {real, imag} */,
  {32'hbe935174, 32'hba0d9140} /* (29, 17, 27) {real, imag} */,
  {32'hbe8c1689, 32'hbdca48bc} /* (29, 17, 26) {real, imag} */,
  {32'h3dd1e19f, 32'h3dad99e6} /* (29, 17, 25) {real, imag} */,
  {32'h3cf41c9a, 32'h3e952ed5} /* (29, 17, 24) {real, imag} */,
  {32'hbe5b7497, 32'h3e5fe5a6} /* (29, 17, 23) {real, imag} */,
  {32'hbe6c8c82, 32'hbc9f1510} /* (29, 17, 22) {real, imag} */,
  {32'h3f02d0aa, 32'hbdcda594} /* (29, 17, 21) {real, imag} */,
  {32'h3ebc3036, 32'h3f0f8754} /* (29, 17, 20) {real, imag} */,
  {32'hbd0cd7e4, 32'h3e3e1c3a} /* (29, 17, 19) {real, imag} */,
  {32'h3d0800bc, 32'h3daf6958} /* (29, 17, 18) {real, imag} */,
  {32'hbe15f09a, 32'h3d105943} /* (29, 17, 17) {real, imag} */,
  {32'hbdc23242, 32'h3e57c8c1} /* (29, 17, 16) {real, imag} */,
  {32'hbb955bc0, 32'h3d5c3074} /* (29, 17, 15) {real, imag} */,
  {32'h3e91214b, 32'h3df0ae3d} /* (29, 17, 14) {real, imag} */,
  {32'h3e970064, 32'h3e36ba7e} /* (29, 17, 13) {real, imag} */,
  {32'hbe9e7f3b, 32'hbe2c8158} /* (29, 17, 12) {real, imag} */,
  {32'h3ebfc9da, 32'hbbbc8950} /* (29, 17, 11) {real, imag} */,
  {32'hbe3c3cca, 32'hbe1ab975} /* (29, 17, 10) {real, imag} */,
  {32'hbd708154, 32'h3ea79397} /* (29, 17, 9) {real, imag} */,
  {32'h3ea5993c, 32'hbf16bb08} /* (29, 17, 8) {real, imag} */,
  {32'h3ed1aa62, 32'h3dc45adf} /* (29, 17, 7) {real, imag} */,
  {32'h3e36eef4, 32'hbf1484af} /* (29, 17, 6) {real, imag} */,
  {32'h3dbea870, 32'h3c3ab560} /* (29, 17, 5) {real, imag} */,
  {32'hbe881ff2, 32'h3e8713df} /* (29, 17, 4) {real, imag} */,
  {32'h3e28ab0c, 32'hbec1c69a} /* (29, 17, 3) {real, imag} */,
  {32'h3ecdaac1, 32'h3dcbfdf2} /* (29, 17, 2) {real, imag} */,
  {32'hbdf8e9f0, 32'hbe88e117} /* (29, 17, 1) {real, imag} */,
  {32'h3e0800ae, 32'hbd831845} /* (29, 17, 0) {real, imag} */,
  {32'hbc955428, 32'hbdb9a658} /* (29, 16, 31) {real, imag} */,
  {32'h3e9e2693, 32'h3e15f4bc} /* (29, 16, 30) {real, imag} */,
  {32'hbcff918e, 32'hbe5f2856} /* (29, 16, 29) {real, imag} */,
  {32'hbce50b2c, 32'hbdd59718} /* (29, 16, 28) {real, imag} */,
  {32'h3ea0a2a8, 32'h3e637287} /* (29, 16, 27) {real, imag} */,
  {32'hbe0276d9, 32'hbd1b1aa8} /* (29, 16, 26) {real, imag} */,
  {32'hbd3d5c3f, 32'h3e9015cc} /* (29, 16, 25) {real, imag} */,
  {32'hbe95e63a, 32'hbdbb1ea2} /* (29, 16, 24) {real, imag} */,
  {32'h3ee812e0, 32'h3ed865a5} /* (29, 16, 23) {real, imag} */,
  {32'hbe7a732f, 32'h3d2336c4} /* (29, 16, 22) {real, imag} */,
  {32'hbeb05132, 32'hbe833e4f} /* (29, 16, 21) {real, imag} */,
  {32'hbd2e88b0, 32'hbe6a9dac} /* (29, 16, 20) {real, imag} */,
  {32'hbe1d1c89, 32'h3dba2b30} /* (29, 16, 19) {real, imag} */,
  {32'h3f0ec182, 32'hbdf39af2} /* (29, 16, 18) {real, imag} */,
  {32'h3d99de53, 32'hbde537fe} /* (29, 16, 17) {real, imag} */,
  {32'hbd41b8d5, 32'h00000000} /* (29, 16, 16) {real, imag} */,
  {32'h3d99de53, 32'h3de537fe} /* (29, 16, 15) {real, imag} */,
  {32'h3f0ec182, 32'h3df39af2} /* (29, 16, 14) {real, imag} */,
  {32'hbe1d1c89, 32'hbdba2b30} /* (29, 16, 13) {real, imag} */,
  {32'hbd2e88b0, 32'h3e6a9dac} /* (29, 16, 12) {real, imag} */,
  {32'hbeb05132, 32'h3e833e4f} /* (29, 16, 11) {real, imag} */,
  {32'hbe7a732f, 32'hbd2336c4} /* (29, 16, 10) {real, imag} */,
  {32'h3ee812e0, 32'hbed865a5} /* (29, 16, 9) {real, imag} */,
  {32'hbe95e63a, 32'h3dbb1ea2} /* (29, 16, 8) {real, imag} */,
  {32'hbd3d5c3f, 32'hbe9015cc} /* (29, 16, 7) {real, imag} */,
  {32'hbe0276d9, 32'h3d1b1aa8} /* (29, 16, 6) {real, imag} */,
  {32'h3ea0a2a8, 32'hbe637287} /* (29, 16, 5) {real, imag} */,
  {32'hbce50b2c, 32'h3dd59718} /* (29, 16, 4) {real, imag} */,
  {32'hbcff918e, 32'h3e5f2856} /* (29, 16, 3) {real, imag} */,
  {32'h3e9e2693, 32'hbe15f4bc} /* (29, 16, 2) {real, imag} */,
  {32'hbc955428, 32'h3db9a658} /* (29, 16, 1) {real, imag} */,
  {32'h3e9952a2, 32'h00000000} /* (29, 16, 0) {real, imag} */,
  {32'hbdf8e9f0, 32'h3e88e117} /* (29, 15, 31) {real, imag} */,
  {32'h3ecdaac1, 32'hbdcbfdf2} /* (29, 15, 30) {real, imag} */,
  {32'h3e28ab0c, 32'h3ec1c69a} /* (29, 15, 29) {real, imag} */,
  {32'hbe881ff2, 32'hbe8713df} /* (29, 15, 28) {real, imag} */,
  {32'h3dbea870, 32'hbc3ab560} /* (29, 15, 27) {real, imag} */,
  {32'h3e36eef4, 32'h3f1484af} /* (29, 15, 26) {real, imag} */,
  {32'h3ed1aa62, 32'hbdc45adf} /* (29, 15, 25) {real, imag} */,
  {32'h3ea5993c, 32'h3f16bb08} /* (29, 15, 24) {real, imag} */,
  {32'hbd708154, 32'hbea79397} /* (29, 15, 23) {real, imag} */,
  {32'hbe3c3cca, 32'h3e1ab975} /* (29, 15, 22) {real, imag} */,
  {32'h3ebfc9da, 32'h3bbc8950} /* (29, 15, 21) {real, imag} */,
  {32'hbe9e7f3b, 32'h3e2c8158} /* (29, 15, 20) {real, imag} */,
  {32'h3e970064, 32'hbe36ba7e} /* (29, 15, 19) {real, imag} */,
  {32'h3e91214b, 32'hbdf0ae3d} /* (29, 15, 18) {real, imag} */,
  {32'hbb955bc0, 32'hbd5c3074} /* (29, 15, 17) {real, imag} */,
  {32'hbdc23242, 32'hbe57c8c1} /* (29, 15, 16) {real, imag} */,
  {32'hbe15f09a, 32'hbd105943} /* (29, 15, 15) {real, imag} */,
  {32'h3d0800bc, 32'hbdaf6958} /* (29, 15, 14) {real, imag} */,
  {32'hbd0cd7e4, 32'hbe3e1c3a} /* (29, 15, 13) {real, imag} */,
  {32'h3ebc3036, 32'hbf0f8754} /* (29, 15, 12) {real, imag} */,
  {32'h3f02d0aa, 32'h3dcda594} /* (29, 15, 11) {real, imag} */,
  {32'hbe6c8c82, 32'h3c9f1510} /* (29, 15, 10) {real, imag} */,
  {32'hbe5b7497, 32'hbe5fe5a6} /* (29, 15, 9) {real, imag} */,
  {32'h3cf41c9a, 32'hbe952ed5} /* (29, 15, 8) {real, imag} */,
  {32'h3dd1e19f, 32'hbdad99e6} /* (29, 15, 7) {real, imag} */,
  {32'hbe8c1689, 32'h3dca48bc} /* (29, 15, 6) {real, imag} */,
  {32'hbe935174, 32'h3a0d9140} /* (29, 15, 5) {real, imag} */,
  {32'hbd6184d4, 32'hbe705478} /* (29, 15, 4) {real, imag} */,
  {32'h3e482168, 32'hbcfba950} /* (29, 15, 3) {real, imag} */,
  {32'h3d438797, 32'hbdad04a4} /* (29, 15, 2) {real, imag} */,
  {32'h3e2b920e, 32'h3e373a0e} /* (29, 15, 1) {real, imag} */,
  {32'h3e0800ae, 32'h3d831845} /* (29, 15, 0) {real, imag} */,
  {32'hbe3acb3a, 32'hbe476a52} /* (29, 14, 31) {real, imag} */,
  {32'hbdb16950, 32'hbdf46d44} /* (29, 14, 30) {real, imag} */,
  {32'h3e28f0e9, 32'hbf06260c} /* (29, 14, 29) {real, imag} */,
  {32'h3c9bf610, 32'hbd122038} /* (29, 14, 28) {real, imag} */,
  {32'h3e8dbc0c, 32'h3e9b8340} /* (29, 14, 27) {real, imag} */,
  {32'hbe874b84, 32'hbeaba979} /* (29, 14, 26) {real, imag} */,
  {32'hbe368c7a, 32'h3e16c349} /* (29, 14, 25) {real, imag} */,
  {32'h3e02645b, 32'hbd04a8a0} /* (29, 14, 24) {real, imag} */,
  {32'hbd02a664, 32'hbb3603d0} /* (29, 14, 23) {real, imag} */,
  {32'h3ea00cc8, 32'hbd434d1a} /* (29, 14, 22) {real, imag} */,
  {32'hbd1302e3, 32'hbf2f83af} /* (29, 14, 21) {real, imag} */,
  {32'h3d923474, 32'hbe6cdd78} /* (29, 14, 20) {real, imag} */,
  {32'hbd32b52e, 32'hbd6e57c8} /* (29, 14, 19) {real, imag} */,
  {32'h3e847f12, 32'hbd3fbe30} /* (29, 14, 18) {real, imag} */,
  {32'hbd21cfba, 32'h3dfbf516} /* (29, 14, 17) {real, imag} */,
  {32'h3e8a6f9c, 32'hbe1b0381} /* (29, 14, 16) {real, imag} */,
  {32'hbd3157b4, 32'hbe79927c} /* (29, 14, 15) {real, imag} */,
  {32'hbe5af0ef, 32'hbe004178} /* (29, 14, 14) {real, imag} */,
  {32'h3e9b7695, 32'hbe9f1686} /* (29, 14, 13) {real, imag} */,
  {32'hbf006a97, 32'hbe805194} /* (29, 14, 12) {real, imag} */,
  {32'hbe53f290, 32'h3ea15912} /* (29, 14, 11) {real, imag} */,
  {32'hbe560cb1, 32'hbf1a111f} /* (29, 14, 10) {real, imag} */,
  {32'h3f48eb5d, 32'hbf01a58b} /* (29, 14, 9) {real, imag} */,
  {32'h3e2d8112, 32'hbe2af467} /* (29, 14, 8) {real, imag} */,
  {32'hbf1ef27f, 32'h3eb63de2} /* (29, 14, 7) {real, imag} */,
  {32'h3e2d07bc, 32'h3e72cf76} /* (29, 14, 6) {real, imag} */,
  {32'hbef24c12, 32'h3e4658ea} /* (29, 14, 5) {real, imag} */,
  {32'hbed2f3f5, 32'h3ec8d664} /* (29, 14, 4) {real, imag} */,
  {32'hbea32008, 32'h3eb6105d} /* (29, 14, 3) {real, imag} */,
  {32'hbd2467bc, 32'h3e7f90b0} /* (29, 14, 2) {real, imag} */,
  {32'hbe7a2e6d, 32'hbe8707ee} /* (29, 14, 1) {real, imag} */,
  {32'hbe2a0964, 32'hbee009d4} /* (29, 14, 0) {real, imag} */,
  {32'hbca2fcb0, 32'h3d595910} /* (29, 13, 31) {real, imag} */,
  {32'h3ee358bc, 32'hbe6ed2cc} /* (29, 13, 30) {real, imag} */,
  {32'hbeeaabeb, 32'h3ee35331} /* (29, 13, 29) {real, imag} */,
  {32'h3ddb3e8a, 32'hbd8be55c} /* (29, 13, 28) {real, imag} */,
  {32'h3dd1b777, 32'h3dbb4199} /* (29, 13, 27) {real, imag} */,
  {32'h3f07376e, 32'hbe0685e3} /* (29, 13, 26) {real, imag} */,
  {32'hbde5fabc, 32'hbe8e6d62} /* (29, 13, 25) {real, imag} */,
  {32'h3e387803, 32'hbdff2c93} /* (29, 13, 24) {real, imag} */,
  {32'h3ec8dc6a, 32'h3f1cab74} /* (29, 13, 23) {real, imag} */,
  {32'hbe0feb33, 32'hbeb3276c} /* (29, 13, 22) {real, imag} */,
  {32'h3ee98bfc, 32'h3e9ae316} /* (29, 13, 21) {real, imag} */,
  {32'hbd3dbbd4, 32'h3e86436c} /* (29, 13, 20) {real, imag} */,
  {32'h3dde8208, 32'hbc406b20} /* (29, 13, 19) {real, imag} */,
  {32'hbe71bd1f, 32'hbdf28fd4} /* (29, 13, 18) {real, imag} */,
  {32'hbe00ecc7, 32'hbe9a0e5c} /* (29, 13, 17) {real, imag} */,
  {32'hbd50d4c0, 32'hbde6795e} /* (29, 13, 16) {real, imag} */,
  {32'hbd3505dc, 32'h3f254efe} /* (29, 13, 15) {real, imag} */,
  {32'h3f049638, 32'hbdf1d478} /* (29, 13, 14) {real, imag} */,
  {32'h3e4973af, 32'hbe44c7bb} /* (29, 13, 13) {real, imag} */,
  {32'h3e969ef8, 32'hbeb40c84} /* (29, 13, 12) {real, imag} */,
  {32'hbdfd5ab4, 32'hbe0848ca} /* (29, 13, 11) {real, imag} */,
  {32'hbe80cf90, 32'h3e29573e} /* (29, 13, 10) {real, imag} */,
  {32'hbefe61ae, 32'hbd7ce973} /* (29, 13, 9) {real, imag} */,
  {32'hbe6ba2e8, 32'h3d124400} /* (29, 13, 8) {real, imag} */,
  {32'h3d9b16a4, 32'hbda99531} /* (29, 13, 7) {real, imag} */,
  {32'h3e067b7c, 32'h3d51cc44} /* (29, 13, 6) {real, imag} */,
  {32'hbf0caf56, 32'hbea6147f} /* (29, 13, 5) {real, imag} */,
  {32'h3ea547c9, 32'h3c59a290} /* (29, 13, 4) {real, imag} */,
  {32'h3eacb908, 32'hbe5e57a6} /* (29, 13, 3) {real, imag} */,
  {32'h3c5770fc, 32'hbf0ba3cd} /* (29, 13, 2) {real, imag} */,
  {32'h3e54a2ee, 32'h3e97d557} /* (29, 13, 1) {real, imag} */,
  {32'h3f212d44, 32'h3ec45c50} /* (29, 13, 0) {real, imag} */,
  {32'h3e6cb2d6, 32'h3ea11ae9} /* (29, 12, 31) {real, imag} */,
  {32'h3e4f02d0, 32'h3e04ae80} /* (29, 12, 30) {real, imag} */,
  {32'hbe1eff65, 32'h3f041617} /* (29, 12, 29) {real, imag} */,
  {32'h3f397dd8, 32'hbcbfae98} /* (29, 12, 28) {real, imag} */,
  {32'h3d37ef96, 32'hbead2b92} /* (29, 12, 27) {real, imag} */,
  {32'h3dcdbab0, 32'h3e896148} /* (29, 12, 26) {real, imag} */,
  {32'hbe758c0c, 32'hbec1bfd4} /* (29, 12, 25) {real, imag} */,
  {32'h3daa7c00, 32'h3de8fc05} /* (29, 12, 24) {real, imag} */,
  {32'hbf0be8cd, 32'hbd57e876} /* (29, 12, 23) {real, imag} */,
  {32'hbe0abd26, 32'hbf1835cc} /* (29, 12, 22) {real, imag} */,
  {32'hbec51336, 32'h3eb1647c} /* (29, 12, 21) {real, imag} */,
  {32'h3ddaa03d, 32'h3e6c6b61} /* (29, 12, 20) {real, imag} */,
  {32'h3ca2587f, 32'h3e658bcc} /* (29, 12, 19) {real, imag} */,
  {32'h3e7f429a, 32'h3e6ea53f} /* (29, 12, 18) {real, imag} */,
  {32'hbd71b190, 32'hbd690a0c} /* (29, 12, 17) {real, imag} */,
  {32'hbe20e8e4, 32'h3c3c7b30} /* (29, 12, 16) {real, imag} */,
  {32'h3e1fb6de, 32'h3dc34418} /* (29, 12, 15) {real, imag} */,
  {32'hbe87228e, 32'hbe1da82e} /* (29, 12, 14) {real, imag} */,
  {32'h3e332ed5, 32'hbe7687fc} /* (29, 12, 13) {real, imag} */,
  {32'hbe113716, 32'h3ee658ad} /* (29, 12, 12) {real, imag} */,
  {32'h3ea1d2d3, 32'hbf05c4bf} /* (29, 12, 11) {real, imag} */,
  {32'hbed48e53, 32'h3d859a5c} /* (29, 12, 10) {real, imag} */,
  {32'h3e199126, 32'hbd8b8296} /* (29, 12, 9) {real, imag} */,
  {32'hbf1d60be, 32'h3d2f4ba0} /* (29, 12, 8) {real, imag} */,
  {32'hbeac6ea6, 32'hbeb6ffd2} /* (29, 12, 7) {real, imag} */,
  {32'h3e1ad192, 32'hbd7c850e} /* (29, 12, 6) {real, imag} */,
  {32'h3c3310d8, 32'h3e810fb9} /* (29, 12, 5) {real, imag} */,
  {32'hbdc6f93c, 32'hbebbc80d} /* (29, 12, 4) {real, imag} */,
  {32'h3d81bb26, 32'h3e19f5d0} /* (29, 12, 3) {real, imag} */,
  {32'hbf167eae, 32'hbc968e10} /* (29, 12, 2) {real, imag} */,
  {32'h3e047005, 32'hbd89a964} /* (29, 12, 1) {real, imag} */,
  {32'hbe056e92, 32'hbe2ffb60} /* (29, 12, 0) {real, imag} */,
  {32'hbe71669e, 32'hbeb7be2a} /* (29, 11, 31) {real, imag} */,
  {32'h3e01b80b, 32'h3ed5cd53} /* (29, 11, 30) {real, imag} */,
  {32'h3eb57124, 32'hbdad3ed4} /* (29, 11, 29) {real, imag} */,
  {32'h3edfd46e, 32'h3db78fbf} /* (29, 11, 28) {real, imag} */,
  {32'h3d8de658, 32'hbf00de65} /* (29, 11, 27) {real, imag} */,
  {32'hbec0c734, 32'h3e9f8e09} /* (29, 11, 26) {real, imag} */,
  {32'h3ec08d4c, 32'h3e457db5} /* (29, 11, 25) {real, imag} */,
  {32'hbe998ce8, 32'hbdd8c814} /* (29, 11, 24) {real, imag} */,
  {32'hbe3b9e5e, 32'h3e9154d4} /* (29, 11, 23) {real, imag} */,
  {32'hbf302278, 32'h3e51fb2a} /* (29, 11, 22) {real, imag} */,
  {32'h3e871699, 32'hbf08a7f0} /* (29, 11, 21) {real, imag} */,
  {32'h3e815a29, 32'hbe7cdc92} /* (29, 11, 20) {real, imag} */,
  {32'h3ee1e42e, 32'hbc968420} /* (29, 11, 19) {real, imag} */,
  {32'hbeb5e27a, 32'hbe9b7e1e} /* (29, 11, 18) {real, imag} */,
  {32'h3cb4fd70, 32'h3e268cac} /* (29, 11, 17) {real, imag} */,
  {32'hbe274d4e, 32'hbdc7046c} /* (29, 11, 16) {real, imag} */,
  {32'hbf0a0f4c, 32'h3e1d8042} /* (29, 11, 15) {real, imag} */,
  {32'hbdd38ea9, 32'hbf010ee0} /* (29, 11, 14) {real, imag} */,
  {32'hbe94815e, 32'hbdb09f50} /* (29, 11, 13) {real, imag} */,
  {32'h3e709d21, 32'hbe64a33d} /* (29, 11, 12) {real, imag} */,
  {32'hbe79ada9, 32'hbd8e350a} /* (29, 11, 11) {real, imag} */,
  {32'h3f0d3517, 32'hbdb5bba6} /* (29, 11, 10) {real, imag} */,
  {32'h3f4d18fc, 32'h3da2d232} /* (29, 11, 9) {real, imag} */,
  {32'h3e2e3a98, 32'h3eafe429} /* (29, 11, 8) {real, imag} */,
  {32'hbd314d3e, 32'h3e32f829} /* (29, 11, 7) {real, imag} */,
  {32'hbeea89be, 32'h3edf8912} /* (29, 11, 6) {real, imag} */,
  {32'hbe90ef5f, 32'h3f0a923c} /* (29, 11, 5) {real, imag} */,
  {32'hbefe4fe0, 32'h3f0673a6} /* (29, 11, 4) {real, imag} */,
  {32'hbdb1742e, 32'h3e25b40a} /* (29, 11, 3) {real, imag} */,
  {32'hbe0ca481, 32'h3f81279d} /* (29, 11, 2) {real, imag} */,
  {32'hbdad1db6, 32'hbf68f050} /* (29, 11, 1) {real, imag} */,
  {32'hbf48c8d5, 32'hbf6190a6} /* (29, 11, 0) {real, imag} */,
  {32'h3f093280, 32'h3e6251be} /* (29, 10, 31) {real, imag} */,
  {32'h3e08d53f, 32'hbe8a0253} /* (29, 10, 30) {real, imag} */,
  {32'h3e9fd5c0, 32'h3ec31c44} /* (29, 10, 29) {real, imag} */,
  {32'h3dbd040a, 32'h3ccf1120} /* (29, 10, 28) {real, imag} */,
  {32'h3f02ceb2, 32'hbed45c67} /* (29, 10, 27) {real, imag} */,
  {32'h3e0dd4ca, 32'hbee1c73e} /* (29, 10, 26) {real, imag} */,
  {32'h3e8fb50b, 32'h3e947ef8} /* (29, 10, 25) {real, imag} */,
  {32'hbdcc0f8a, 32'hbf31cc43} /* (29, 10, 24) {real, imag} */,
  {32'hbef49658, 32'h3e399fe2} /* (29, 10, 23) {real, imag} */,
  {32'h3d86baee, 32'h3f2bb94a} /* (29, 10, 22) {real, imag} */,
  {32'h3e0d77a2, 32'hbe77c95c} /* (29, 10, 21) {real, imag} */,
  {32'h3ea5c536, 32'hbe951ed2} /* (29, 10, 20) {real, imag} */,
  {32'h3e80663a, 32'hbecd31a0} /* (29, 10, 19) {real, imag} */,
  {32'h3d8a3a04, 32'h3e5e0e08} /* (29, 10, 18) {real, imag} */,
  {32'h3c6dba88, 32'h3dfe5fa2} /* (29, 10, 17) {real, imag} */,
  {32'hbecfa086, 32'h3e53c999} /* (29, 10, 16) {real, imag} */,
  {32'h3ef0d46d, 32'hbe5c259e} /* (29, 10, 15) {real, imag} */,
  {32'h3f2c238a, 32'hbc86ee38} /* (29, 10, 14) {real, imag} */,
  {32'hbf1a7738, 32'h3db57cd4} /* (29, 10, 13) {real, imag} */,
  {32'h3e2c7e6a, 32'h3efc905a} /* (29, 10, 12) {real, imag} */,
  {32'h3efb1dd4, 32'h3e06643c} /* (29, 10, 11) {real, imag} */,
  {32'h3e096bcc, 32'h3eb8ed01} /* (29, 10, 10) {real, imag} */,
  {32'hbe8ad5a8, 32'h3dfea94f} /* (29, 10, 9) {real, imag} */,
  {32'hbe598cdb, 32'h3e8b345d} /* (29, 10, 8) {real, imag} */,
  {32'h3ec935dc, 32'hbed38068} /* (29, 10, 7) {real, imag} */,
  {32'h3e965c5e, 32'hbecad827} /* (29, 10, 6) {real, imag} */,
  {32'hbea42e18, 32'h3d8cda36} /* (29, 10, 5) {real, imag} */,
  {32'hbf25fbab, 32'hbf0ca5de} /* (29, 10, 4) {real, imag} */,
  {32'hbf28222c, 32'hbd082e0e} /* (29, 10, 3) {real, imag} */,
  {32'h3d7663b8, 32'h3dedcbda} /* (29, 10, 2) {real, imag} */,
  {32'h3cf4b9b0, 32'hbd7ec1f8} /* (29, 10, 1) {real, imag} */,
  {32'hbf040ff1, 32'h3e42fdb9} /* (29, 10, 0) {real, imag} */,
  {32'hbf9d4b78, 32'h3eafedfd} /* (29, 9, 31) {real, imag} */,
  {32'h3f700e87, 32'hbdfb6408} /* (29, 9, 30) {real, imag} */,
  {32'h3e80e1f9, 32'hbb9a2040} /* (29, 9, 29) {real, imag} */,
  {32'hbce141d8, 32'h3f6fc942} /* (29, 9, 28) {real, imag} */,
  {32'hbed1f940, 32'h3e14e59e} /* (29, 9, 27) {real, imag} */,
  {32'hbdaa9e82, 32'h3eddbb75} /* (29, 9, 26) {real, imag} */,
  {32'hbeb92f02, 32'h3ddce680} /* (29, 9, 25) {real, imag} */,
  {32'h3e03e961, 32'hbe8b2d18} /* (29, 9, 24) {real, imag} */,
  {32'hbe553f06, 32'h3ed5ebef} /* (29, 9, 23) {real, imag} */,
  {32'hbf704259, 32'hbebd588e} /* (29, 9, 22) {real, imag} */,
  {32'hbecf2d0e, 32'hbe89a696} /* (29, 9, 21) {real, imag} */,
  {32'hbe579ffe, 32'hbf0e8cc6} /* (29, 9, 20) {real, imag} */,
  {32'h3ed3fefe, 32'h3f2b96ae} /* (29, 9, 19) {real, imag} */,
  {32'h3ec9cf49, 32'h3e2e3d66} /* (29, 9, 18) {real, imag} */,
  {32'hbe8b350c, 32'hbe87cac0} /* (29, 9, 17) {real, imag} */,
  {32'h3edf7688, 32'hbe7ac36d} /* (29, 9, 16) {real, imag} */,
  {32'hbdee75a7, 32'h3e59ecc3} /* (29, 9, 15) {real, imag} */,
  {32'hbe6d99bb, 32'h3f085a56} /* (29, 9, 14) {real, imag} */,
  {32'hbede9694, 32'h3f054fae} /* (29, 9, 13) {real, imag} */,
  {32'h3e9cbcc0, 32'h3ea104bd} /* (29, 9, 12) {real, imag} */,
  {32'h3bba46b0, 32'hbe5a6d4f} /* (29, 9, 11) {real, imag} */,
  {32'hbf3aa175, 32'h3dd6bba8} /* (29, 9, 10) {real, imag} */,
  {32'hbe8b4b9e, 32'hbb2d58c0} /* (29, 9, 9) {real, imag} */,
  {32'h3ee32176, 32'hbe607702} /* (29, 9, 8) {real, imag} */,
  {32'hbde05c1a, 32'hbe7a94a6} /* (29, 9, 7) {real, imag} */,
  {32'h3e6d125e, 32'hbd322ba9} /* (29, 9, 6) {real, imag} */,
  {32'h3e1fd260, 32'h3f4d0b14} /* (29, 9, 5) {real, imag} */,
  {32'h3d36dd06, 32'hbd49c147} /* (29, 9, 4) {real, imag} */,
  {32'hbec8c264, 32'h3dbee9ba} /* (29, 9, 3) {real, imag} */,
  {32'hbf402127, 32'hbf034bcc} /* (29, 9, 2) {real, imag} */,
  {32'h3f4e3aae, 32'hbda618c0} /* (29, 9, 1) {real, imag} */,
  {32'hbedb22aa, 32'hbf133602} /* (29, 9, 0) {real, imag} */,
  {32'hbff3bd9a, 32'hbfa6fe51} /* (29, 8, 31) {real, imag} */,
  {32'h3f544fbc, 32'h3f1a93fd} /* (29, 8, 30) {real, imag} */,
  {32'hbd555d70, 32'hbf3ddbb4} /* (29, 8, 29) {real, imag} */,
  {32'h3e9dc24c, 32'hbe62ce16} /* (29, 8, 28) {real, imag} */,
  {32'hbeebd34d, 32'hbe054d50} /* (29, 8, 27) {real, imag} */,
  {32'h3ec51a58, 32'hbe81e3a0} /* (29, 8, 26) {real, imag} */,
  {32'hbead3a13, 32'hbf3215bc} /* (29, 8, 25) {real, imag} */,
  {32'h3d140f90, 32'h3d1534b0} /* (29, 8, 24) {real, imag} */,
  {32'hbe678150, 32'hbd8e0fab} /* (29, 8, 23) {real, imag} */,
  {32'h3f2f30de, 32'hbea20684} /* (29, 8, 22) {real, imag} */,
  {32'h3ef8ce4c, 32'h3ee47cee} /* (29, 8, 21) {real, imag} */,
  {32'hbe7d21e6, 32'hbe607c79} /* (29, 8, 20) {real, imag} */,
  {32'hbeb528bb, 32'h3e010c29} /* (29, 8, 19) {real, imag} */,
  {32'h3ed324bd, 32'hbedadac9} /* (29, 8, 18) {real, imag} */,
  {32'hbb96f480, 32'h3de86fa6} /* (29, 8, 17) {real, imag} */,
  {32'h3e9d3ae3, 32'h3e6db3e6} /* (29, 8, 16) {real, imag} */,
  {32'h3e863393, 32'h3bcd4fc0} /* (29, 8, 15) {real, imag} */,
  {32'hbcd52eb0, 32'hbe82907d} /* (29, 8, 14) {real, imag} */,
  {32'h3f3cf1e7, 32'h3e0f413a} /* (29, 8, 13) {real, imag} */,
  {32'hbde07c02, 32'h3e6b9c1a} /* (29, 8, 12) {real, imag} */,
  {32'hbc8bec78, 32'h3f52b48e} /* (29, 8, 11) {real, imag} */,
  {32'h3e9fbc46, 32'hbeaf67fa} /* (29, 8, 10) {real, imag} */,
  {32'hbe99ed08, 32'hbe75475e} /* (29, 8, 9) {real, imag} */,
  {32'h3df3bfb0, 32'h3e3aa950} /* (29, 8, 8) {real, imag} */,
  {32'hbeef64fa, 32'h3d940df7} /* (29, 8, 7) {real, imag} */,
  {32'hbebd9f33, 32'h3eecfabc} /* (29, 8, 6) {real, imag} */,
  {32'h3e8896a8, 32'h3ef5af81} /* (29, 8, 5) {real, imag} */,
  {32'hbe3e2ea7, 32'hbe87af7c} /* (29, 8, 4) {real, imag} */,
  {32'h3f5554d8, 32'h3f22e601} /* (29, 8, 3) {real, imag} */,
  {32'hbe2afe14, 32'hbee3f56f} /* (29, 8, 2) {real, imag} */,
  {32'hbf0c2148, 32'hbfaca212} /* (29, 8, 1) {real, imag} */,
  {32'hbf066be3, 32'hbe6cc587} /* (29, 8, 0) {real, imag} */,
  {32'hbde7bc7e, 32'hbe8ce8fa} /* (29, 7, 31) {real, imag} */,
  {32'hbf138f1c, 32'h3f5c0515} /* (29, 7, 30) {real, imag} */,
  {32'hbea2feaf, 32'h3d27a23c} /* (29, 7, 29) {real, imag} */,
  {32'hbf21fc78, 32'hbe34d244} /* (29, 7, 28) {real, imag} */,
  {32'h3ea85846, 32'h3f30d7c9} /* (29, 7, 27) {real, imag} */,
  {32'hbe39af4a, 32'h3abe1700} /* (29, 7, 26) {real, imag} */,
  {32'hbefdf12b, 32'h3e5aeb8b} /* (29, 7, 25) {real, imag} */,
  {32'hbc88042a, 32'hbe38d04b} /* (29, 7, 24) {real, imag} */,
  {32'h3afd6300, 32'hbeaa06d7} /* (29, 7, 23) {real, imag} */,
  {32'hbe4eef20, 32'h3f28d10e} /* (29, 7, 22) {real, imag} */,
  {32'hbdf2c9fc, 32'h3eaa4c4f} /* (29, 7, 21) {real, imag} */,
  {32'h3e7e2e4d, 32'h3c891f00} /* (29, 7, 20) {real, imag} */,
  {32'h3ea60a35, 32'h3e3efc9a} /* (29, 7, 19) {real, imag} */,
  {32'h3ea7c3a6, 32'h3e0110bc} /* (29, 7, 18) {real, imag} */,
  {32'hbf013f4c, 32'hbea64641} /* (29, 7, 17) {real, imag} */,
  {32'h3dbb379a, 32'hbe86b1d8} /* (29, 7, 16) {real, imag} */,
  {32'hbc37fe10, 32'hbd97c0e0} /* (29, 7, 15) {real, imag} */,
  {32'hbd2ad8a4, 32'hbe44e83c} /* (29, 7, 14) {real, imag} */,
  {32'hbee84bb8, 32'h3decff98} /* (29, 7, 13) {real, imag} */,
  {32'h3e0b8dea, 32'hbd5e3984} /* (29, 7, 12) {real, imag} */,
  {32'hbe8b6491, 32'h3f022dce} /* (29, 7, 11) {real, imag} */,
  {32'hbe80e071, 32'hbde4a56b} /* (29, 7, 10) {real, imag} */,
  {32'h3ec6f770, 32'h3ece263c} /* (29, 7, 9) {real, imag} */,
  {32'hbe2d8f49, 32'hbdd4b929} /* (29, 7, 8) {real, imag} */,
  {32'hbde95e04, 32'hbeaa0862} /* (29, 7, 7) {real, imag} */,
  {32'h3f4d13f4, 32'hbee7a1ca} /* (29, 7, 6) {real, imag} */,
  {32'h3e0c9a26, 32'hbf592f99} /* (29, 7, 5) {real, imag} */,
  {32'h3ccacd60, 32'hbe0a06cd} /* (29, 7, 4) {real, imag} */,
  {32'hbf3fa8c2, 32'hbeb6ea50} /* (29, 7, 3) {real, imag} */,
  {32'h3ec08744, 32'hbe715334} /* (29, 7, 2) {real, imag} */,
  {32'h3fb7f53c, 32'h3d291360} /* (29, 7, 1) {real, imag} */,
  {32'h3f9315c2, 32'hbdd5a24c} /* (29, 7, 0) {real, imag} */,
  {32'h3ede14bc, 32'h3f4a7d0e} /* (29, 6, 31) {real, imag} */,
  {32'h3f00d86e, 32'h3f22ee15} /* (29, 6, 30) {real, imag} */,
  {32'h3b3bb3a0, 32'h3d06d348} /* (29, 6, 29) {real, imag} */,
  {32'hbdc20a48, 32'hbf32fc21} /* (29, 6, 28) {real, imag} */,
  {32'hbf87fe74, 32'h3defb05f} /* (29, 6, 27) {real, imag} */,
  {32'hbebce9f8, 32'hbde5b973} /* (29, 6, 26) {real, imag} */,
  {32'h3edd6bcc, 32'h3f6f1faa} /* (29, 6, 25) {real, imag} */,
  {32'hbe946fa1, 32'h3f5fc1da} /* (29, 6, 24) {real, imag} */,
  {32'h3f0e5da6, 32'hbe72fce8} /* (29, 6, 23) {real, imag} */,
  {32'hbe8d7024, 32'h3e2ee5ef} /* (29, 6, 22) {real, imag} */,
  {32'hbf17e075, 32'hbe9f4a16} /* (29, 6, 21) {real, imag} */,
  {32'hbd6aee8c, 32'hbe295d83} /* (29, 6, 20) {real, imag} */,
  {32'h3eba5d3a, 32'hbf4160c0} /* (29, 6, 19) {real, imag} */,
  {32'h3ec33878, 32'h3e199570} /* (29, 6, 18) {real, imag} */,
  {32'hbe83dbce, 32'h3e6069c6} /* (29, 6, 17) {real, imag} */,
  {32'h3d23ecf0, 32'h3e807e58} /* (29, 6, 16) {real, imag} */,
  {32'hbeb061fd, 32'hbe8a2db6} /* (29, 6, 15) {real, imag} */,
  {32'hbf080b34, 32'h3e635262} /* (29, 6, 14) {real, imag} */,
  {32'h3ed92c34, 32'h3e7c256f} /* (29, 6, 13) {real, imag} */,
  {32'h3ee00a5e, 32'h3eeb9e9c} /* (29, 6, 12) {real, imag} */,
  {32'h3d68176c, 32'h3f026d5e} /* (29, 6, 11) {real, imag} */,
  {32'h3e47ee34, 32'hbdf9e334} /* (29, 6, 10) {real, imag} */,
  {32'h3e0476ac, 32'h3e00ba64} /* (29, 6, 9) {real, imag} */,
  {32'h3d6a60de, 32'h3dee0e0c} /* (29, 6, 8) {real, imag} */,
  {32'h3f43cc15, 32'h3eaf472b} /* (29, 6, 7) {real, imag} */,
  {32'hbc0aae40, 32'h3df0b19c} /* (29, 6, 6) {real, imag} */,
  {32'h3e7182c8, 32'h3d741818} /* (29, 6, 5) {real, imag} */,
  {32'h3f024f82, 32'hbe4bf979} /* (29, 6, 4) {real, imag} */,
  {32'h3e0fcf25, 32'hbb4405c0} /* (29, 6, 3) {real, imag} */,
  {32'hb920a800, 32'hbda5bc9c} /* (29, 6, 2) {real, imag} */,
  {32'hbf580c40, 32'h3ede2120} /* (29, 6, 1) {real, imag} */,
  {32'h3e9ef882, 32'h3eb8a253} /* (29, 6, 0) {real, imag} */,
  {32'hc05a22bc, 32'hbf1b92e9} /* (29, 5, 31) {real, imag} */,
  {32'h3e65522e, 32'hbf581c36} /* (29, 5, 30) {real, imag} */,
  {32'h3ed74e96, 32'hbf3ddeb1} /* (29, 5, 29) {real, imag} */,
  {32'hbf2b6320, 32'h3ee612d7} /* (29, 5, 28) {real, imag} */,
  {32'h3f94df07, 32'h3eb15bc9} /* (29, 5, 27) {real, imag} */,
  {32'h3e346253, 32'hbeff8d9c} /* (29, 5, 26) {real, imag} */,
  {32'hbf1da539, 32'h3ea1be85} /* (29, 5, 25) {real, imag} */,
  {32'hbe59e0a2, 32'h3bd9dd10} /* (29, 5, 24) {real, imag} */,
  {32'hbe6b3758, 32'hbe8f080e} /* (29, 5, 23) {real, imag} */,
  {32'h3de93fec, 32'h3f4e8117} /* (29, 5, 22) {real, imag} */,
  {32'h3f1ed5c1, 32'hbdc07660} /* (29, 5, 21) {real, imag} */,
  {32'hbdda8138, 32'h3e365176} /* (29, 5, 20) {real, imag} */,
  {32'h3e5bbbea, 32'h3c722748} /* (29, 5, 19) {real, imag} */,
  {32'h3dd646e2, 32'h3d8d6d65} /* (29, 5, 18) {real, imag} */,
  {32'h3e35f004, 32'h3e1008ce} /* (29, 5, 17) {real, imag} */,
  {32'h3db405a2, 32'hbe223b46} /* (29, 5, 16) {real, imag} */,
  {32'hbd6742d0, 32'h3e1da836} /* (29, 5, 15) {real, imag} */,
  {32'h3d86e269, 32'hbe238b44} /* (29, 5, 14) {real, imag} */,
  {32'hbe33532a, 32'hbde486fe} /* (29, 5, 13) {real, imag} */,
  {32'h3d92dcda, 32'hbc2b1660} /* (29, 5, 12) {real, imag} */,
  {32'h3d8a1da1, 32'hbe5ddeef} /* (29, 5, 11) {real, imag} */,
  {32'hbf06ab3e, 32'hbe54db47} /* (29, 5, 10) {real, imag} */,
  {32'hbd912d60, 32'h3d13a558} /* (29, 5, 9) {real, imag} */,
  {32'h3e5950e5, 32'h3cf51580} /* (29, 5, 8) {real, imag} */,
  {32'h3e2ea345, 32'h3dc49fa8} /* (29, 5, 7) {real, imag} */,
  {32'hbe321746, 32'hbebccb46} /* (29, 5, 6) {real, imag} */,
  {32'hbce208c0, 32'h3f97000c} /* (29, 5, 5) {real, imag} */,
  {32'hbefe69bd, 32'hbe838b41} /* (29, 5, 4) {real, imag} */,
  {32'h3e4611ae, 32'hbec938be} /* (29, 5, 3) {real, imag} */,
  {32'h3fa46168, 32'hbc94cae0} /* (29, 5, 2) {real, imag} */,
  {32'hc011ac68, 32'hbfde705c} /* (29, 5, 1) {real, imag} */,
  {32'hbff9715a, 32'hbf86368c} /* (29, 5, 0) {real, imag} */,
  {32'h402757d7, 32'h401cd0ce} /* (29, 4, 31) {real, imag} */,
  {32'hc019d5af, 32'hbf7d2350} /* (29, 4, 30) {real, imag} */,
  {32'hbf89de3a, 32'h3fee653c} /* (29, 4, 29) {real, imag} */,
  {32'h3f8c07fc, 32'hbdb6ad34} /* (29, 4, 28) {real, imag} */,
  {32'hbfe983fa, 32'h3f25379e} /* (29, 4, 27) {real, imag} */,
  {32'h3e352336, 32'h3ec5bc19} /* (29, 4, 26) {real, imag} */,
  {32'hbe6ea136, 32'h3c7c1050} /* (29, 4, 25) {real, imag} */,
  {32'hbec31488, 32'h3cdd0a88} /* (29, 4, 24) {real, imag} */,
  {32'hbf021620, 32'hbf1be7ae} /* (29, 4, 23) {real, imag} */,
  {32'h3daa60fc, 32'hbe3751f0} /* (29, 4, 22) {real, imag} */,
  {32'h3d77d138, 32'hbe5ed278} /* (29, 4, 21) {real, imag} */,
  {32'hbe096b6e, 32'hbe855abe} /* (29, 4, 20) {real, imag} */,
  {32'h3e80ccfc, 32'hbeb86b56} /* (29, 4, 19) {real, imag} */,
  {32'hbf3b638d, 32'hbdd35941} /* (29, 4, 18) {real, imag} */,
  {32'h3eadada3, 32'hbcf2dfa8} /* (29, 4, 17) {real, imag} */,
  {32'hbe228a79, 32'hbd175a39} /* (29, 4, 16) {real, imag} */,
  {32'hbea14475, 32'hbc81c6e8} /* (29, 4, 15) {real, imag} */,
  {32'hbe1c403e, 32'h3dfcb684} /* (29, 4, 14) {real, imag} */,
  {32'h3e301119, 32'hbef8d3d8} /* (29, 4, 13) {real, imag} */,
  {32'hbead7468, 32'hbea3988c} /* (29, 4, 12) {real, imag} */,
  {32'h3da0e28b, 32'h3ee666ec} /* (29, 4, 11) {real, imag} */,
  {32'hbd68f344, 32'h3e9e8616} /* (29, 4, 10) {real, imag} */,
  {32'h3e40acc6, 32'hbefff297} /* (29, 4, 9) {real, imag} */,
  {32'hbe9b468f, 32'hbebe9f39} /* (29, 4, 8) {real, imag} */,
  {32'h3e8d7a3c, 32'hbeb88083} /* (29, 4, 7) {real, imag} */,
  {32'hbdcdb624, 32'h3ec7aaed} /* (29, 4, 6) {real, imag} */,
  {32'h3d27d09a, 32'hbf582390} /* (29, 4, 5) {real, imag} */,
  {32'h3f4d952e, 32'h3ecac78e} /* (29, 4, 4) {real, imag} */,
  {32'h3e76001b, 32'hbe349028} /* (29, 4, 3) {real, imag} */,
  {32'hbf92ba78, 32'hbffea0c2} /* (29, 4, 2) {real, imag} */,
  {32'h40a04205, 32'h400c80a3} /* (29, 4, 1) {real, imag} */,
  {32'h3fd3fc1a, 32'h3f871e66} /* (29, 4, 0) {real, imag} */,
  {32'hc0754d4c, 32'h401403bf} /* (29, 3, 31) {real, imag} */,
  {32'h4005dcc3, 32'hc01d31b6} /* (29, 3, 30) {real, imag} */,
  {32'h3d9a5a4c, 32'h3efa681b} /* (29, 3, 29) {real, imag} */,
  {32'h3efd76fd, 32'h3f646c6a} /* (29, 3, 28) {real, imag} */,
  {32'hbe3b6a7c, 32'hbf9dc348} /* (29, 3, 27) {real, imag} */,
  {32'hbe311c4a, 32'h3e843564} /* (29, 3, 26) {real, imag} */,
  {32'hbe843f86, 32'h3e9607ae} /* (29, 3, 25) {real, imag} */,
  {32'hbecbbb9a, 32'hbf35f5b2} /* (29, 3, 24) {real, imag} */,
  {32'h3e92f84d, 32'h3d57fa70} /* (29, 3, 23) {real, imag} */,
  {32'h3e37213a, 32'hbccccad8} /* (29, 3, 22) {real, imag} */,
  {32'hbf6f964a, 32'h3d334a00} /* (29, 3, 21) {real, imag} */,
  {32'h3e2cb71a, 32'h3eb36d6a} /* (29, 3, 20) {real, imag} */,
  {32'hbeb35c07, 32'h3e861542} /* (29, 3, 19) {real, imag} */,
  {32'hbe14c728, 32'hbb194f20} /* (29, 3, 18) {real, imag} */,
  {32'h3d807b5c, 32'h3dc77155} /* (29, 3, 17) {real, imag} */,
  {32'hbdb9534a, 32'hbdd8d5d9} /* (29, 3, 16) {real, imag} */,
  {32'h3e3cc4aa, 32'hbe8420a1} /* (29, 3, 15) {real, imag} */,
  {32'h3d6a1162, 32'h3e316024} /* (29, 3, 14) {real, imag} */,
  {32'h3e55aaa8, 32'hbda87e92} /* (29, 3, 13) {real, imag} */,
  {32'h3eb6dc91, 32'h3f013486} /* (29, 3, 12) {real, imag} */,
  {32'hbd52d808, 32'hbce89cf0} /* (29, 3, 11) {real, imag} */,
  {32'h3dea5ab8, 32'hbe401e90} /* (29, 3, 10) {real, imag} */,
  {32'h3e5c5bac, 32'hbd03dc8a} /* (29, 3, 9) {real, imag} */,
  {32'hbe0a70d2, 32'hbc8cb730} /* (29, 3, 8) {real, imag} */,
  {32'h3f5a5811, 32'h3e1c433c} /* (29, 3, 7) {real, imag} */,
  {32'hbf4935f0, 32'hbf253013} /* (29, 3, 6) {real, imag} */,
  {32'hbc547b00, 32'h3e02952c} /* (29, 3, 5) {real, imag} */,
  {32'hbec2324c, 32'h3f7b9454} /* (29, 3, 4) {real, imag} */,
  {32'h3f003b05, 32'h3ee188aa} /* (29, 3, 3) {real, imag} */,
  {32'hbdc5ee4c, 32'hc01b7f9e} /* (29, 3, 2) {real, imag} */,
  {32'h400333fa, 32'h40713afc} /* (29, 3, 1) {real, imag} */,
  {32'h3e839992, 32'hbd112a38} /* (29, 3, 0) {real, imag} */,
  {32'hc1b5e489, 32'hbf480b8a} /* (29, 2, 31) {real, imag} */,
  {32'h414cf7ac, 32'hc0903bce} /* (29, 2, 30) {real, imag} */,
  {32'h3e7bede4, 32'hbed50b5a} /* (29, 2, 29) {real, imag} */,
  {32'hbf8df8e2, 32'h401fef6e} /* (29, 2, 28) {real, imag} */,
  {32'h3fcbd6e6, 32'hbf4d27c1} /* (29, 2, 27) {real, imag} */,
  {32'h3e8ebeba, 32'h3e9c4232} /* (29, 2, 26) {real, imag} */,
  {32'hbda7b968, 32'h3f73f13f} /* (29, 2, 25) {real, imag} */,
  {32'h3f99f172, 32'hbf2b32ee} /* (29, 2, 24) {real, imag} */,
  {32'hbe6dcd34, 32'hbdba5248} /* (29, 2, 23) {real, imag} */,
  {32'h3ea2f6ad, 32'h3f1941f3} /* (29, 2, 22) {real, imag} */,
  {32'h3ebaccce, 32'hbeb2d43e} /* (29, 2, 21) {real, imag} */,
  {32'hbf0e3ab9, 32'h3ee1cc11} /* (29, 2, 20) {real, imag} */,
  {32'hbdb966c4, 32'hbeb68f86} /* (29, 2, 19) {real, imag} */,
  {32'h3e87b257, 32'hbbf42080} /* (29, 2, 18) {real, imag} */,
  {32'hbd1e136e, 32'h3e503fb5} /* (29, 2, 17) {real, imag} */,
  {32'h3e561933, 32'hbe5684e9} /* (29, 2, 16) {real, imag} */,
  {32'hbe1ed663, 32'hbe6248c8} /* (29, 2, 15) {real, imag} */,
  {32'h3df1c924, 32'h3e58a92f} /* (29, 2, 14) {real, imag} */,
  {32'h3e17fee6, 32'hbefc5bf3} /* (29, 2, 13) {real, imag} */,
  {32'h3d67d760, 32'h3eabaf6c} /* (29, 2, 12) {real, imag} */,
  {32'h3ed28e85, 32'h3ea6298e} /* (29, 2, 11) {real, imag} */,
  {32'hbf001f2f, 32'h3f0c7bd0} /* (29, 2, 10) {real, imag} */,
  {32'h3ee98acd, 32'h3e22cc1f} /* (29, 2, 9) {real, imag} */,
  {32'hbe2d2634, 32'h3e8bf4a1} /* (29, 2, 8) {real, imag} */,
  {32'h3ed4c7f0, 32'hbe9d8360} /* (29, 2, 7) {real, imag} */,
  {32'h3d0e2640, 32'h3ef25786} /* (29, 2, 6) {real, imag} */,
  {32'h3f9b7092, 32'h3ebf1c97} /* (29, 2, 5) {real, imag} */,
  {32'hbfe3036c, 32'hbef5a0d6} /* (29, 2, 4) {real, imag} */,
  {32'hbf3d1c38, 32'hbf23899d} /* (29, 2, 3) {real, imag} */,
  {32'h4108fdd2, 32'hc01f5e9c} /* (29, 2, 2) {real, imag} */,
  {32'hc164ca54, 32'h4083ee06} /* (29, 2, 1) {real, imag} */,
  {32'hc13e597d, 32'hbfe894af} /* (29, 2, 0) {real, imag} */,
  {32'h41a0b567, 32'hc0c716e8} /* (29, 1, 31) {real, imag} */,
  {32'hc10976e2, 32'h3df29c18} /* (29, 1, 30) {real, imag} */,
  {32'hbe34d694, 32'hbf06f9a0} /* (29, 1, 29) {real, imag} */,
  {32'h3fc5a46a, 32'h40000d1f} /* (29, 1, 28) {real, imag} */,
  {32'hc069e5bc, 32'h3fb4c304} /* (29, 1, 27) {real, imag} */,
  {32'hbf166796, 32'h3dfde660} /* (29, 1, 26) {real, imag} */,
  {32'h3ced8b00, 32'hbfba28f8} /* (29, 1, 25) {real, imag} */,
  {32'h3de0bee0, 32'h3f4062bd} /* (29, 1, 24) {real, imag} */,
  {32'h3e1f221c, 32'hbdbc9a68} /* (29, 1, 23) {real, imag} */,
  {32'h3eb5fd69, 32'hbe6b686f} /* (29, 1, 22) {real, imag} */,
  {32'hbe1a43f6, 32'h3f32db66} /* (29, 1, 21) {real, imag} */,
  {32'hbe35c04e, 32'h3e327d7b} /* (29, 1, 20) {real, imag} */,
  {32'h3ebf87fc, 32'h3db9c239} /* (29, 1, 19) {real, imag} */,
  {32'hbf0de0e5, 32'h3e341b40} /* (29, 1, 18) {real, imag} */,
  {32'h3d23cfd8, 32'h3d0d225c} /* (29, 1, 17) {real, imag} */,
  {32'hbe6a626f, 32'hbe90d995} /* (29, 1, 16) {real, imag} */,
  {32'h3de8306e, 32'h3db09a0e} /* (29, 1, 15) {real, imag} */,
  {32'h3e8d20a3, 32'hbebc3204} /* (29, 1, 14) {real, imag} */,
  {32'h3de37cec, 32'hbe746b4a} /* (29, 1, 13) {real, imag} */,
  {32'h3e218aee, 32'h3e1d66f0} /* (29, 1, 12) {real, imag} */,
  {32'h3e22a97c, 32'hbef7e64d} /* (29, 1, 11) {real, imag} */,
  {32'hbf5014ec, 32'h3cefafe0} /* (29, 1, 10) {real, imag} */,
  {32'hbeac2cae, 32'h3e58be7f} /* (29, 1, 9) {real, imag} */,
  {32'hbe53e927, 32'hbf62fc62} /* (29, 1, 8) {real, imag} */,
  {32'hbeb03fd2, 32'h3e80b5bc} /* (29, 1, 7) {real, imag} */,
  {32'hbea3bcfc, 32'h3ed5cc87} /* (29, 1, 6) {real, imag} */,
  {32'hc00d7d19, 32'hbf862d79} /* (29, 1, 5) {real, imag} */,
  {32'h3fbcf852, 32'h3f8e7a8a} /* (29, 1, 4) {real, imag} */,
  {32'hbf46232c, 32'h3fc49552} /* (29, 1, 3) {real, imag} */,
  {32'hc140cccc, 32'hc163363a} /* (29, 1, 2) {real, imag} */,
  {32'h41e981a4, 32'h41456bdc} /* (29, 1, 1) {real, imag} */,
  {32'h418e6846, 32'h403994f4} /* (29, 1, 0) {real, imag} */,
  {32'h410603c2, 32'hc10835c3} /* (29, 0, 31) {real, imag} */,
  {32'hc0432d0d, 32'h40f73eef} /* (29, 0, 30) {real, imag} */,
  {32'hbf95baf1, 32'hbf0c93e8} /* (29, 0, 29) {real, imag} */,
  {32'h3e13818c, 32'h3f615320} /* (29, 0, 28) {real, imag} */,
  {32'hbfe6f9e6, 32'hbf6a217b} /* (29, 0, 27) {real, imag} */,
  {32'hbe41a960, 32'hbf1ed9b6} /* (29, 0, 26) {real, imag} */,
  {32'hbf0267a2, 32'hbf864156} /* (29, 0, 25) {real, imag} */,
  {32'h3e3b7ca4, 32'h3f1cadc1} /* (29, 0, 24) {real, imag} */,
  {32'h3cf47f40, 32'h3efc8a75} /* (29, 0, 23) {real, imag} */,
  {32'h3ee1b7ee, 32'h3e8fcec0} /* (29, 0, 22) {real, imag} */,
  {32'h3e31375c, 32'h3eab3296} /* (29, 0, 21) {real, imag} */,
  {32'hbceff390, 32'hbe27ebdb} /* (29, 0, 20) {real, imag} */,
  {32'hbe27f065, 32'hbe84b613} /* (29, 0, 19) {real, imag} */,
  {32'h3d3d8f28, 32'h3dfe152c} /* (29, 0, 18) {real, imag} */,
  {32'h3e27850e, 32'hbecebffe} /* (29, 0, 17) {real, imag} */,
  {32'hbcd2eae4, 32'h00000000} /* (29, 0, 16) {real, imag} */,
  {32'h3e27850e, 32'h3ecebffe} /* (29, 0, 15) {real, imag} */,
  {32'h3d3d8f28, 32'hbdfe152c} /* (29, 0, 14) {real, imag} */,
  {32'hbe27f065, 32'h3e84b613} /* (29, 0, 13) {real, imag} */,
  {32'hbceff390, 32'h3e27ebdb} /* (29, 0, 12) {real, imag} */,
  {32'h3e31375c, 32'hbeab3296} /* (29, 0, 11) {real, imag} */,
  {32'h3ee1b7ee, 32'hbe8fcec0} /* (29, 0, 10) {real, imag} */,
  {32'h3cf47f40, 32'hbefc8a75} /* (29, 0, 9) {real, imag} */,
  {32'h3e3b7ca4, 32'hbf1cadc1} /* (29, 0, 8) {real, imag} */,
  {32'hbf0267a2, 32'h3f864156} /* (29, 0, 7) {real, imag} */,
  {32'hbe41a960, 32'h3f1ed9b6} /* (29, 0, 6) {real, imag} */,
  {32'hbfe6f9e6, 32'h3f6a217b} /* (29, 0, 5) {real, imag} */,
  {32'h3e13818c, 32'hbf615320} /* (29, 0, 4) {real, imag} */,
  {32'hbf95baf1, 32'h3f0c93e8} /* (29, 0, 3) {real, imag} */,
  {32'hc0432d0d, 32'hc0f73eef} /* (29, 0, 2) {real, imag} */,
  {32'h410603c2, 32'h410835c3} /* (29, 0, 1) {real, imag} */,
  {32'h3fbd556c, 32'h00000000} /* (29, 0, 0) {real, imag} */,
  {32'h41cdec3a, 32'hc12fa2b3} /* (28, 31, 31) {real, imag} */,
  {32'hc13d1793, 32'h4149ec43} /* (28, 31, 30) {real, imag} */,
  {32'hc002ece5, 32'h3c8ac020} /* (28, 31, 29) {real, imag} */,
  {32'h3fb9a870, 32'hbe89da7e} /* (28, 31, 28) {real, imag} */,
  {32'hc000a52d, 32'h3f6dc7c4} /* (28, 31, 27) {real, imag} */,
  {32'hbcef8a40, 32'h3eba8ec6} /* (28, 31, 26) {real, imag} */,
  {32'hbefcf2b4, 32'hbf44bdc6} /* (28, 31, 25) {real, imag} */,
  {32'h3d11aba8, 32'h3f3c0a80} /* (28, 31, 24) {real, imag} */,
  {32'hbdba5e10, 32'h3e9e695c} /* (28, 31, 23) {real, imag} */,
  {32'hbea8a226, 32'hbd9808ef} /* (28, 31, 22) {real, imag} */,
  {32'hbe9b96d6, 32'hbe7ef79c} /* (28, 31, 21) {real, imag} */,
  {32'h3e1ef4c2, 32'h3e053a7b} /* (28, 31, 20) {real, imag} */,
  {32'hbcbe7d64, 32'hbe8294c1} /* (28, 31, 19) {real, imag} */,
  {32'h3edc89a0, 32'h3f29389a} /* (28, 31, 18) {real, imag} */,
  {32'h3e121178, 32'hbea50ee0} /* (28, 31, 17) {real, imag} */,
  {32'h3d965326, 32'h3e2ed598} /* (28, 31, 16) {real, imag} */,
  {32'h3d6a361c, 32'hbe3c4fa0} /* (28, 31, 15) {real, imag} */,
  {32'h3dc34f80, 32'hbdc0008a} /* (28, 31, 14) {real, imag} */,
  {32'hbea21359, 32'hbc05bf20} /* (28, 31, 13) {real, imag} */,
  {32'h3d8e97fe, 32'h3e1e0274} /* (28, 31, 12) {real, imag} */,
  {32'hbee114bc, 32'hbd983bde} /* (28, 31, 11) {real, imag} */,
  {32'hbf1a26a2, 32'hbeb75566} /* (28, 31, 10) {real, imag} */,
  {32'h3a521e00, 32'hbebaa354} /* (28, 31, 9) {real, imag} */,
  {32'hbefdf928, 32'hbe7519ed} /* (28, 31, 8) {real, imag} */,
  {32'hbd1710c0, 32'h3f095d26} /* (28, 31, 7) {real, imag} */,
  {32'hbf05e7f1, 32'hbdc1ae04} /* (28, 31, 6) {real, imag} */,
  {32'hc05fa512, 32'hbf8113ad} /* (28, 31, 5) {real, imag} */,
  {32'h3fc26a2e, 32'hbf984bf4} /* (28, 31, 4) {real, imag} */,
  {32'h3e17c6c0, 32'hbea07c5e} /* (28, 31, 3) {real, imag} */,
  {32'hc1036f90, 32'hbf9e4a7b} /* (28, 31, 2) {real, imag} */,
  {32'h418cc812, 32'h40be7672} /* (28, 31, 1) {real, imag} */,
  {32'h415cc76e, 32'hbff21544} /* (28, 31, 0) {real, imag} */,
  {32'hc141e4c5, 32'hc04a20c0} /* (28, 30, 31) {real, imag} */,
  {32'h4117c4b4, 32'h4077ff4a} /* (28, 30, 30) {real, imag} */,
  {32'hbf0954e4, 32'h3d6781ec} /* (28, 30, 29) {real, imag} */,
  {32'hc033813b, 32'h3f89fa5c} /* (28, 30, 28) {real, imag} */,
  {32'h3fb2b837, 32'hbf5b6217} /* (28, 30, 27) {real, imag} */,
  {32'hbdf7b184, 32'h3db1178c} /* (28, 30, 26) {real, imag} */,
  {32'hbeb7df7c, 32'h3e600a9f} /* (28, 30, 25) {real, imag} */,
  {32'h3f39549f, 32'hbf2bbf56} /* (28, 30, 24) {real, imag} */,
  {32'h3e5d10dc, 32'hbf351a8e} /* (28, 30, 23) {real, imag} */,
  {32'hbef9d68c, 32'h3e5814a0} /* (28, 30, 22) {real, imag} */,
  {32'h3cdf00b8, 32'hbe40afd6} /* (28, 30, 21) {real, imag} */,
  {32'hbe990331, 32'h3e3d0ec8} /* (28, 30, 20) {real, imag} */,
  {32'hbdfcbe84, 32'hbe438fe1} /* (28, 30, 19) {real, imag} */,
  {32'h3d53b17e, 32'hbecb86f1} /* (28, 30, 18) {real, imag} */,
  {32'hbe2e6e97, 32'hbe786131} /* (28, 30, 17) {real, imag} */,
  {32'h3e82a39e, 32'h3df3909e} /* (28, 30, 16) {real, imag} */,
  {32'hbe22ff02, 32'hbef7f5b3} /* (28, 30, 15) {real, imag} */,
  {32'h3e90b6a0, 32'h3ee3d349} /* (28, 30, 14) {real, imag} */,
  {32'hbe5d4be1, 32'hbe987722} /* (28, 30, 13) {real, imag} */,
  {32'h3e3fd038, 32'h3e762b38} /* (28, 30, 12) {real, imag} */,
  {32'h3c113890, 32'h3f76fb7c} /* (28, 30, 11) {real, imag} */,
  {32'h3f384a46, 32'hbdb5454a} /* (28, 30, 10) {real, imag} */,
  {32'h3e0152ed, 32'h3e668edf} /* (28, 30, 9) {real, imag} */,
  {32'h3e19aa95, 32'h3fa48af4} /* (28, 30, 8) {real, imag} */,
  {32'hbd3658fa, 32'hbfac00c3} /* (28, 30, 7) {real, imag} */,
  {32'h3f31fa1a, 32'hbf3fc7c6} /* (28, 30, 6) {real, imag} */,
  {32'h3f591d94, 32'h3f688b18} /* (28, 30, 5) {real, imag} */,
  {32'hbf485007, 32'hc02efa3a} /* (28, 30, 4) {real, imag} */,
  {32'hbf0fec69, 32'h3e764a62} /* (28, 30, 3) {real, imag} */,
  {32'h4145513e, 32'h409b8fb2} /* (28, 30, 2) {real, imag} */,
  {32'hc1a5e041, 32'hbf51e393} /* (28, 30, 1) {real, imag} */,
  {32'hc12f5eb5, 32'h40199eaa} /* (28, 30, 0) {real, imag} */,
  {32'h4013bb0d, 32'hc0998610} /* (28, 29, 31) {real, imag} */,
  {32'hbefb7dbb, 32'h40477516} /* (28, 29, 30) {real, imag} */,
  {32'h3f6276c6, 32'hbf00af85} /* (28, 29, 29) {real, imag} */,
  {32'hbd84ecfc, 32'hbfacba7a} /* (28, 29, 28) {real, imag} */,
  {32'h3f5510a9, 32'h3dd698e0} /* (28, 29, 27) {real, imag} */,
  {32'hbfd6890a, 32'h3f2326ad} /* (28, 29, 26) {real, imag} */,
  {32'h3f0c29a3, 32'hbe854129} /* (28, 29, 25) {real, imag} */,
  {32'h3d8e7b46, 32'h3e5e8a86} /* (28, 29, 24) {real, imag} */,
  {32'hbe1ac983, 32'hbeea7ee3} /* (28, 29, 23) {real, imag} */,
  {32'hbddabf1e, 32'hbe3b725c} /* (28, 29, 22) {real, imag} */,
  {32'h3ed7585b, 32'h3ef86ded} /* (28, 29, 21) {real, imag} */,
  {32'hbe52c720, 32'h3f03d950} /* (28, 29, 20) {real, imag} */,
  {32'hbeeeccb0, 32'h3f22567f} /* (28, 29, 19) {real, imag} */,
  {32'hbe0e4213, 32'h3d921e58} /* (28, 29, 18) {real, imag} */,
  {32'h3e61b17c, 32'hbd4854e0} /* (28, 29, 17) {real, imag} */,
  {32'hbe8146e2, 32'hbc26fa20} /* (28, 29, 16) {real, imag} */,
  {32'hbe2c6ec9, 32'h3e9f7e50} /* (28, 29, 15) {real, imag} */,
  {32'h3df06cdc, 32'h3ebfeffc} /* (28, 29, 14) {real, imag} */,
  {32'hbe732a1b, 32'h3e32d14f} /* (28, 29, 13) {real, imag} */,
  {32'h3ed013f8, 32'h3d6a8bca} /* (28, 29, 12) {real, imag} */,
  {32'hbf1f03d1, 32'h3c75abc0} /* (28, 29, 11) {real, imag} */,
  {32'h3f72ea15, 32'hbf877ad3} /* (28, 29, 10) {real, imag} */,
  {32'h3e8de770, 32'hbf02c896} /* (28, 29, 9) {real, imag} */,
  {32'hbdf943ea, 32'h3f69089a} /* (28, 29, 8) {real, imag} */,
  {32'hbefa7386, 32'hbed16e46} /* (28, 29, 7) {real, imag} */,
  {32'h3f09f571, 32'h3d8f7f58} /* (28, 29, 6) {real, imag} */,
  {32'hbea83e50, 32'h3f69021b} /* (28, 29, 5) {real, imag} */,
  {32'h3ebdf34d, 32'hbf4e12ce} /* (28, 29, 4) {real, imag} */,
  {32'hbf215212, 32'hbe6c96c6} /* (28, 29, 3) {real, imag} */,
  {32'h4015b366, 32'h403f95c8} /* (28, 29, 2) {real, imag} */,
  {32'hc0930f7f, 32'hbfa2f434} /* (28, 29, 1) {real, imag} */,
  {32'h3f2fc724, 32'h3f037278} /* (28, 29, 0) {real, imag} */,
  {32'h40649c41, 32'hc018f1ba} /* (28, 28, 31) {real, imag} */,
  {32'hbfe7b92e, 32'h40171cfb} /* (28, 28, 30) {real, imag} */,
  {32'h3f4aaf5d, 32'h3f867e75} /* (28, 28, 29) {real, imag} */,
  {32'h3fbcd1c2, 32'h3f5339ac} /* (28, 28, 28) {real, imag} */,
  {32'h3e519af8, 32'h3eac549a} /* (28, 28, 27) {real, imag} */,
  {32'hbd3f92e0, 32'hbf2b8bc5} /* (28, 28, 26) {real, imag} */,
  {32'hbf09befe, 32'hbd907e14} /* (28, 28, 25) {real, imag} */,
  {32'h3d5705cf, 32'h3e842c3c} /* (28, 28, 24) {real, imag} */,
  {32'hbef840ee, 32'h3eab2690} /* (28, 28, 23) {real, imag} */,
  {32'hbd84ea30, 32'hbe024f41} /* (28, 28, 22) {real, imag} */,
  {32'h3ddbd804, 32'hbecf20ad} /* (28, 28, 21) {real, imag} */,
  {32'h3e021d9c, 32'h3f1e1e44} /* (28, 28, 20) {real, imag} */,
  {32'h3deeec6e, 32'hbe4a7927} /* (28, 28, 19) {real, imag} */,
  {32'hbe3d3b40, 32'hbd9d4bc6} /* (28, 28, 18) {real, imag} */,
  {32'hbea14080, 32'hbea3fe6d} /* (28, 28, 17) {real, imag} */,
  {32'h3db2c1a2, 32'h3dab470d} /* (28, 28, 16) {real, imag} */,
  {32'hbdbbc62e, 32'hbde235a0} /* (28, 28, 15) {real, imag} */,
  {32'h3ca8abe8, 32'hbe089076} /* (28, 28, 14) {real, imag} */,
  {32'hbcff2968, 32'h3d8e6de5} /* (28, 28, 13) {real, imag} */,
  {32'h3f3b9cca, 32'h3ebc2635} /* (28, 28, 12) {real, imag} */,
  {32'hbf236ae0, 32'hbe4daa93} /* (28, 28, 11) {real, imag} */,
  {32'hbe8ad9fd, 32'hbe141e22} /* (28, 28, 10) {real, imag} */,
  {32'hbefeac1b, 32'hbe2930be} /* (28, 28, 9) {real, imag} */,
  {32'hbeca3c29, 32'hbd9d77fb} /* (28, 28, 8) {real, imag} */,
  {32'h3e8cca1c, 32'h3eab05ac} /* (28, 28, 7) {real, imag} */,
  {32'h3f02e4c3, 32'hbef4cc02} /* (28, 28, 6) {real, imag} */,
  {32'hbde7cb7f, 32'hbe272a54} /* (28, 28, 5) {real, imag} */,
  {32'h3f813465, 32'h3e94d7c5} /* (28, 28, 4) {real, imag} */,
  {32'h3e3e0f14, 32'h3d9291f4} /* (28, 28, 3) {real, imag} */,
  {32'hc0085c64, 32'h3fba225d} /* (28, 28, 2) {real, imag} */,
  {32'h4002ba56, 32'hc00cc1ba} /* (28, 28, 1) {real, imag} */,
  {32'h3f8b550a, 32'hbfcf361d} /* (28, 28, 0) {real, imag} */,
  {32'hc0142d54, 32'h3fd087b0} /* (28, 27, 31) {real, imag} */,
  {32'h3f5d4471, 32'h3f594585} /* (28, 27, 30) {real, imag} */,
  {32'hbeb86856, 32'h3f2153dc} /* (28, 27, 29) {real, imag} */,
  {32'h3ddeccb8, 32'hbf21b553} /* (28, 27, 28) {real, imag} */,
  {32'h3f21eb24, 32'hbf4e45cd} /* (28, 27, 27) {real, imag} */,
  {32'hbdba380e, 32'hbd9d063c} /* (28, 27, 26) {real, imag} */,
  {32'h3d359c66, 32'hbe9f0d35} /* (28, 27, 25) {real, imag} */,
  {32'h3c279cbc, 32'hbeb82bf8} /* (28, 27, 24) {real, imag} */,
  {32'h3e947aa6, 32'h3f00c0eb} /* (28, 27, 23) {real, imag} */,
  {32'hbe5ccc51, 32'h3ee532ad} /* (28, 27, 22) {real, imag} */,
  {32'hbdec5adc, 32'hbe68cee0} /* (28, 27, 21) {real, imag} */,
  {32'h3e75ef3b, 32'h3e5d6a0a} /* (28, 27, 20) {real, imag} */,
  {32'hbd89a5ca, 32'h3dafa0cc} /* (28, 27, 19) {real, imag} */,
  {32'hbdf51552, 32'hbe0ff4c6} /* (28, 27, 18) {real, imag} */,
  {32'hbd985527, 32'hbe8e20b4} /* (28, 27, 17) {real, imag} */,
  {32'hbd6690c3, 32'h3e302633} /* (28, 27, 16) {real, imag} */,
  {32'hbd1b95e8, 32'h3f031d68} /* (28, 27, 15) {real, imag} */,
  {32'hbd7ada94, 32'hbe98b7c9} /* (28, 27, 14) {real, imag} */,
  {32'hbe969420, 32'hbd5c67a0} /* (28, 27, 13) {real, imag} */,
  {32'h3c2a8f78, 32'h3d427362} /* (28, 27, 12) {real, imag} */,
  {32'h3eae30f6, 32'h3ecc6f27} /* (28, 27, 11) {real, imag} */,
  {32'h3e91e984, 32'hbd6cf340} /* (28, 27, 10) {real, imag} */,
  {32'h3e84279e, 32'hbe3016d9} /* (28, 27, 9) {real, imag} */,
  {32'h3d925730, 32'h3db9732f} /* (28, 27, 8) {real, imag} */,
  {32'h3ee5f15d, 32'hbf27feae} /* (28, 27, 7) {real, imag} */,
  {32'h3ecba2aa, 32'h3f2832d4} /* (28, 27, 6) {real, imag} */,
  {32'h3f94909c, 32'hbe5d58af} /* (28, 27, 5) {real, imag} */,
  {32'hbf1e8c5a, 32'hbe08a5c8} /* (28, 27, 4) {real, imag} */,
  {32'h3e136b43, 32'h3f4181aa} /* (28, 27, 3) {real, imag} */,
  {32'h3f05815e, 32'h3e87527e} /* (28, 27, 2) {real, imag} */,
  {32'hc055b67a, 32'h3f3b7554} /* (28, 27, 1) {real, imag} */,
  {32'hbff36a56, 32'h3f9e2570} /* (28, 27, 0) {real, imag} */,
  {32'hbf0b3c59, 32'h3ea1aa63} /* (28, 26, 31) {real, imag} */,
  {32'h3e4a8dbc, 32'h3c051f08} /* (28, 26, 30) {real, imag} */,
  {32'h3e927e10, 32'hbe5a764b} /* (28, 26, 29) {real, imag} */,
  {32'h3e6370ce, 32'hbdb416b8} /* (28, 26, 28) {real, imag} */,
  {32'hbe0edf2f, 32'h3af837c0} /* (28, 26, 27) {real, imag} */,
  {32'hbea8d14f, 32'hbeb1d618} /* (28, 26, 26) {real, imag} */,
  {32'h3f433aa0, 32'hbf03f672} /* (28, 26, 25) {real, imag} */,
  {32'hbd5aa980, 32'h3f1d89ba} /* (28, 26, 24) {real, imag} */,
  {32'h3ead0edc, 32'h3ed1388c} /* (28, 26, 23) {real, imag} */,
  {32'hbefe4aae, 32'hbec43ff2} /* (28, 26, 22) {real, imag} */,
  {32'h3f064051, 32'h3d548410} /* (28, 26, 21) {real, imag} */,
  {32'h3e39fe10, 32'h3dbd548c} /* (28, 26, 20) {real, imag} */,
  {32'hbdfcedd8, 32'hbee60a54} /* (28, 26, 19) {real, imag} */,
  {32'hbdbb76bc, 32'h3debca14} /* (28, 26, 18) {real, imag} */,
  {32'h3dd0d53f, 32'hbe2819f4} /* (28, 26, 17) {real, imag} */,
  {32'hbd8b5341, 32'h3ee8dd12} /* (28, 26, 16) {real, imag} */,
  {32'h3e7e5a48, 32'hbddd92d4} /* (28, 26, 15) {real, imag} */,
  {32'hbe944c0e, 32'hbd62ea7a} /* (28, 26, 14) {real, imag} */,
  {32'h3e0e56cb, 32'h3ebd70b8} /* (28, 26, 13) {real, imag} */,
  {32'h3ea4a72c, 32'hbdc8d146} /* (28, 26, 12) {real, imag} */,
  {32'h3c2e24d0, 32'h3df44f74} /* (28, 26, 11) {real, imag} */,
  {32'h3ddd1eb2, 32'hbe9a2f64} /* (28, 26, 10) {real, imag} */,
  {32'h3d54e3c4, 32'h3dd95322} /* (28, 26, 9) {real, imag} */,
  {32'h3e588c08, 32'hbf2ba1e5} /* (28, 26, 8) {real, imag} */,
  {32'h3e53b6f0, 32'hbefd03bc} /* (28, 26, 7) {real, imag} */,
  {32'h3eaf2d98, 32'h3d77fc68} /* (28, 26, 6) {real, imag} */,
  {32'hbf311803, 32'h3e5403c1} /* (28, 26, 5) {real, imag} */,
  {32'hbe128b16, 32'h3eceb5da} /* (28, 26, 4) {real, imag} */,
  {32'h3ebc8296, 32'hbea5708d} /* (28, 26, 3) {real, imag} */,
  {32'h3f244c66, 32'hbf262a9c} /* (28, 26, 2) {real, imag} */,
  {32'hbf251b2e, 32'h3c8f16f0} /* (28, 26, 1) {real, imag} */,
  {32'hbda41964, 32'hbee3cbaa} /* (28, 26, 0) {real, imag} */,
  {32'h3f754ef2, 32'hbea3ccd3} /* (28, 25, 31) {real, imag} */,
  {32'hbecc56b0, 32'hbe6f60a3} /* (28, 25, 30) {real, imag} */,
  {32'hbf0ea72a, 32'hbf04f07a} /* (28, 25, 29) {real, imag} */,
  {32'hbde310c4, 32'hbe84a790} /* (28, 25, 28) {real, imag} */,
  {32'h3e63469c, 32'h3d1adb18} /* (28, 25, 27) {real, imag} */,
  {32'hbe6f16e4, 32'h3dc5746b} /* (28, 25, 26) {real, imag} */,
  {32'h3eec5cd6, 32'hbeb5bfe3} /* (28, 25, 25) {real, imag} */,
  {32'hbe95c0fa, 32'h3f0f20e6} /* (28, 25, 24) {real, imag} */,
  {32'hbe4789c4, 32'h3d852f2a} /* (28, 25, 23) {real, imag} */,
  {32'hbcffb334, 32'h3e365b9e} /* (28, 25, 22) {real, imag} */,
  {32'hbdbe3264, 32'h3ee19751} /* (28, 25, 21) {real, imag} */,
  {32'hbdf46f60, 32'hbd7d9f48} /* (28, 25, 20) {real, imag} */,
  {32'hbee5cd5a, 32'hbd696304} /* (28, 25, 19) {real, imag} */,
  {32'h3ebd555a, 32'h3e703682} /* (28, 25, 18) {real, imag} */,
  {32'h3e9ca8a7, 32'h3c57fce0} /* (28, 25, 17) {real, imag} */,
  {32'hbdaaf9b4, 32'hbe94efc2} /* (28, 25, 16) {real, imag} */,
  {32'hbd69ef76, 32'h3da527be} /* (28, 25, 15) {real, imag} */,
  {32'hbe70a5b5, 32'hbe2f31b5} /* (28, 25, 14) {real, imag} */,
  {32'h3ef5da1a, 32'hbdfecdee} /* (28, 25, 13) {real, imag} */,
  {32'hbdd8a26f, 32'h3efdacbf} /* (28, 25, 12) {real, imag} */,
  {32'h3cdefc88, 32'hbedc7ef8} /* (28, 25, 11) {real, imag} */,
  {32'hbe90217d, 32'h3f22ab31} /* (28, 25, 10) {real, imag} */,
  {32'hbe0868c6, 32'h3e9e684c} /* (28, 25, 9) {real, imag} */,
  {32'hbedcaef2, 32'hbe046b15} /* (28, 25, 8) {real, imag} */,
  {32'hbe35d977, 32'hbec61cc3} /* (28, 25, 7) {real, imag} */,
  {32'hbe8809b7, 32'h3eccea20} /* (28, 25, 6) {real, imag} */,
  {32'hbf253250, 32'hbf0ad63f} /* (28, 25, 5) {real, imag} */,
  {32'hbe2946a7, 32'h3ee97dd1} /* (28, 25, 4) {real, imag} */,
  {32'hbd13d1a0, 32'h3e0f31f1} /* (28, 25, 3) {real, imag} */,
  {32'hbeaab9d3, 32'hbef4c624} /* (28, 25, 2) {real, imag} */,
  {32'hbee2a2c5, 32'hbdc49763} /* (28, 25, 1) {real, imag} */,
  {32'h3fa2f657, 32'hbdfc1c54} /* (28, 25, 0) {real, imag} */,
  {32'hbf1f16fe, 32'h3f406398} /* (28, 24, 31) {real, imag} */,
  {32'h3d822cd4, 32'h3d89635e} /* (28, 24, 30) {real, imag} */,
  {32'h3b95a910, 32'hbf0b78fe} /* (28, 24, 29) {real, imag} */,
  {32'h3f13f97d, 32'h3f01ebd8} /* (28, 24, 28) {real, imag} */,
  {32'h3edeb9fe, 32'hbd90fe70} /* (28, 24, 27) {real, imag} */,
  {32'h3e8acda3, 32'h3ea5ba40} /* (28, 24, 26) {real, imag} */,
  {32'hbe1e2ad4, 32'h3f567ca9} /* (28, 24, 25) {real, imag} */,
  {32'h3d52e5f0, 32'h3e346c7a} /* (28, 24, 24) {real, imag} */,
  {32'hbdfdb988, 32'hbe514cc2} /* (28, 24, 23) {real, imag} */,
  {32'h3ed9a0b2, 32'hbeb92e61} /* (28, 24, 22) {real, imag} */,
  {32'h3e8ad7be, 32'hbe1bf843} /* (28, 24, 21) {real, imag} */,
  {32'hbe529a4c, 32'hbea1a934} /* (28, 24, 20) {real, imag} */,
  {32'hbe3697b5, 32'h3e098519} /* (28, 24, 19) {real, imag} */,
  {32'h3dcd34de, 32'hbe675e9c} /* (28, 24, 18) {real, imag} */,
  {32'h3e3d625e, 32'hbe2f0488} /* (28, 24, 17) {real, imag} */,
  {32'hbc7180fc, 32'h3ead6cde} /* (28, 24, 16) {real, imag} */,
  {32'hbec94cd6, 32'hbddbf3aa} /* (28, 24, 15) {real, imag} */,
  {32'h3e26b263, 32'hbd579c27} /* (28, 24, 14) {real, imag} */,
  {32'h3eea423c, 32'h3eebf5fe} /* (28, 24, 13) {real, imag} */,
  {32'h3d414118, 32'h3e5df628} /* (28, 24, 12) {real, imag} */,
  {32'h3ec581e2, 32'h3e06f76a} /* (28, 24, 11) {real, imag} */,
  {32'hbc040640, 32'hbdc5824e} /* (28, 24, 10) {real, imag} */,
  {32'h3da86ea0, 32'h3f097cde} /* (28, 24, 9) {real, imag} */,
  {32'hbe830f86, 32'hbe4daa41} /* (28, 24, 8) {real, imag} */,
  {32'h3da34b92, 32'h3ea6f9ba} /* (28, 24, 7) {real, imag} */,
  {32'h3cac371c, 32'hbd7a7c24} /* (28, 24, 6) {real, imag} */,
  {32'hbf728792, 32'h3e4e4eb0} /* (28, 24, 5) {real, imag} */,
  {32'hbf19b2ab, 32'h3c215aec} /* (28, 24, 4) {real, imag} */,
  {32'h3f5ca3b4, 32'h3f086d6e} /* (28, 24, 3) {real, imag} */,
  {32'h3f95138a, 32'hbf1dfc39} /* (28, 24, 2) {real, imag} */,
  {32'hbff28c1c, 32'h3ecb2b93} /* (28, 24, 1) {real, imag} */,
  {32'hbf1e7bf5, 32'h3f063c77} /* (28, 24, 0) {real, imag} */,
  {32'h3eae7387, 32'hbd5e6f48} /* (28, 23, 31) {real, imag} */,
  {32'h3f6c98a6, 32'h3e7add06} /* (28, 23, 30) {real, imag} */,
  {32'hbe35698b, 32'h3df3ca38} /* (28, 23, 29) {real, imag} */,
  {32'h3edb7e9a, 32'h3dea473e} /* (28, 23, 28) {real, imag} */,
  {32'hbe220c90, 32'hbee63c13} /* (28, 23, 27) {real, imag} */,
  {32'hbe766202, 32'hbd4d4cb6} /* (28, 23, 26) {real, imag} */,
  {32'h3e5606be, 32'hbde74f8c} /* (28, 23, 25) {real, imag} */,
  {32'h3e3fa574, 32'h3f12cbe6} /* (28, 23, 24) {real, imag} */,
  {32'hbcb38978, 32'hbe17d866} /* (28, 23, 23) {real, imag} */,
  {32'h3d70f540, 32'hbddaf5aa} /* (28, 23, 22) {real, imag} */,
  {32'hbe9ce7f6, 32'h3e9794a5} /* (28, 23, 21) {real, imag} */,
  {32'hbd2f8006, 32'hbdf5dfb2} /* (28, 23, 20) {real, imag} */,
  {32'h3ded1168, 32'h3e085f9a} /* (28, 23, 19) {real, imag} */,
  {32'hbd704682, 32'hbe862cf3} /* (28, 23, 18) {real, imag} */,
  {32'h3e943200, 32'hbe173744} /* (28, 23, 17) {real, imag} */,
  {32'h3ed77184, 32'hbecdd3be} /* (28, 23, 16) {real, imag} */,
  {32'hbdefb6fa, 32'h3e14fd19} /* (28, 23, 15) {real, imag} */,
  {32'h3e547c06, 32'hbe593c95} /* (28, 23, 14) {real, imag} */,
  {32'hbee5df9b, 32'hbee59258} /* (28, 23, 13) {real, imag} */,
  {32'h3e3b1284, 32'h3dd632d6} /* (28, 23, 12) {real, imag} */,
  {32'hbf3f00f3, 32'h3ef95fbb} /* (28, 23, 11) {real, imag} */,
  {32'hbe0bd5e4, 32'h3ddbab9c} /* (28, 23, 10) {real, imag} */,
  {32'h3e278eea, 32'hbe7b8fc8} /* (28, 23, 9) {real, imag} */,
  {32'hbdf8260a, 32'hbec16772} /* (28, 23, 8) {real, imag} */,
  {32'h3e4e2565, 32'hbe69ab3e} /* (28, 23, 7) {real, imag} */,
  {32'hbe949a26, 32'hbee75a9c} /* (28, 23, 6) {real, imag} */,
  {32'hbeb69914, 32'h3f0782b7} /* (28, 23, 5) {real, imag} */,
  {32'h3ca10a2c, 32'hbe4e5360} /* (28, 23, 4) {real, imag} */,
  {32'hbe1988fe, 32'h3df2de1c} /* (28, 23, 3) {real, imag} */,
  {32'h3f4342b2, 32'h3f7bff59} /* (28, 23, 2) {real, imag} */,
  {32'hbf32bf8d, 32'hbf66e5c8} /* (28, 23, 1) {real, imag} */,
  {32'hbf2c50ea, 32'hbee0da6f} /* (28, 23, 0) {real, imag} */,
  {32'h3e0a17ea, 32'hbdca38fb} /* (28, 22, 31) {real, imag} */,
  {32'hbf032239, 32'h3cc8a720} /* (28, 22, 30) {real, imag} */,
  {32'hbc224bc0, 32'h3e56acd9} /* (28, 22, 29) {real, imag} */,
  {32'h3ed0bca4, 32'hbe32b845} /* (28, 22, 28) {real, imag} */,
  {32'hbef0a6ab, 32'h3e965dbe} /* (28, 22, 27) {real, imag} */,
  {32'hbd904988, 32'hbc4a9fa0} /* (28, 22, 26) {real, imag} */,
  {32'h3e176aba, 32'hbe387c6e} /* (28, 22, 25) {real, imag} */,
  {32'hbf46edfa, 32'hbe280a21} /* (28, 22, 24) {real, imag} */,
  {32'h3e9fa5d4, 32'hbe6e7f0d} /* (28, 22, 23) {real, imag} */,
  {32'hbd04cebc, 32'hbe9e74a2} /* (28, 22, 22) {real, imag} */,
  {32'hbe82966a, 32'hbcfde54c} /* (28, 22, 21) {real, imag} */,
  {32'h3be39680, 32'h3ef092d8} /* (28, 22, 20) {real, imag} */,
  {32'h3e37d593, 32'h3e07cb1c} /* (28, 22, 19) {real, imag} */,
  {32'hbf07b31a, 32'h3e1a5459} /* (28, 22, 18) {real, imag} */,
  {32'hbdafd18c, 32'h3e611de1} /* (28, 22, 17) {real, imag} */,
  {32'h3e1000c8, 32'hbe0d82e0} /* (28, 22, 16) {real, imag} */,
  {32'h3e680d20, 32'h3e429620} /* (28, 22, 15) {real, imag} */,
  {32'h3ee99b1a, 32'h3e4758ca} /* (28, 22, 14) {real, imag} */,
  {32'hbe4f6344, 32'hbe897bf8} /* (28, 22, 13) {real, imag} */,
  {32'h3da0534c, 32'h3e786116} /* (28, 22, 12) {real, imag} */,
  {32'h3d8d501c, 32'h3f066cbb} /* (28, 22, 11) {real, imag} */,
  {32'hbd9ce48a, 32'hbe92992f} /* (28, 22, 10) {real, imag} */,
  {32'h3e81690e, 32'hbcbe9c3e} /* (28, 22, 9) {real, imag} */,
  {32'hbea3c06b, 32'h3d837fd8} /* (28, 22, 8) {real, imag} */,
  {32'h3c3798e0, 32'h3edd496d} /* (28, 22, 7) {real, imag} */,
  {32'h3eb4f770, 32'hbe06a1a8} /* (28, 22, 6) {real, imag} */,
  {32'hbee0849e, 32'h3e781126} /* (28, 22, 5) {real, imag} */,
  {32'h3d90ffc2, 32'h3eb59732} /* (28, 22, 4) {real, imag} */,
  {32'hbdcbed66, 32'hbdfd8934} /* (28, 22, 3) {real, imag} */,
  {32'h3dd4083f, 32'h3f087439} /* (28, 22, 2) {real, imag} */,
  {32'h3ea06018, 32'hbeae1fc9} /* (28, 22, 1) {real, imag} */,
  {32'h3d7cfb4c, 32'hbec6fb89} /* (28, 22, 0) {real, imag} */,
  {32'hbe3c8e69, 32'h3f16f4b7} /* (28, 21, 31) {real, imag} */,
  {32'hbe9dbfd5, 32'hbf6d76ae} /* (28, 21, 30) {real, imag} */,
  {32'h3e5abaf9, 32'hbf17473b} /* (28, 21, 29) {real, imag} */,
  {32'hbeab68c8, 32'h3f15e4b6} /* (28, 21, 28) {real, imag} */,
  {32'h3f499cfc, 32'hbde58230} /* (28, 21, 27) {real, imag} */,
  {32'hbea449da, 32'hbf36cd14} /* (28, 21, 26) {real, imag} */,
  {32'hbabbbb00, 32'h3e4c2418} /* (28, 21, 25) {real, imag} */,
  {32'h3e3482b0, 32'h3ebfd110} /* (28, 21, 24) {real, imag} */,
  {32'h3ee42a99, 32'hbe7c7356} /* (28, 21, 23) {real, imag} */,
  {32'h3ea021d5, 32'hbea3b569} /* (28, 21, 22) {real, imag} */,
  {32'hbe4e6e32, 32'hbeaba89a} /* (28, 21, 21) {real, imag} */,
  {32'hbcd3d770, 32'hbcef0cc0} /* (28, 21, 20) {real, imag} */,
  {32'h3e03f9e7, 32'hbde232f8} /* (28, 21, 19) {real, imag} */,
  {32'h3f0b6103, 32'hbcbf0444} /* (28, 21, 18) {real, imag} */,
  {32'h3e9f2511, 32'hbe030764} /* (28, 21, 17) {real, imag} */,
  {32'hbe070568, 32'hbe5ee0f6} /* (28, 21, 16) {real, imag} */,
  {32'h3db9cd71, 32'hbd5cb90c} /* (28, 21, 15) {real, imag} */,
  {32'hbe8105b2, 32'h3e1a19e0} /* (28, 21, 14) {real, imag} */,
  {32'hbe4c8d13, 32'hbd645ddc} /* (28, 21, 13) {real, imag} */,
  {32'hbf1a5bae, 32'h3cc7b6d0} /* (28, 21, 12) {real, imag} */,
  {32'h3e70c3a4, 32'hbea40018} /* (28, 21, 11) {real, imag} */,
  {32'h3e1a2862, 32'hbe1e350c} /* (28, 21, 10) {real, imag} */,
  {32'hbe59b0f4, 32'h3ef4ea66} /* (28, 21, 9) {real, imag} */,
  {32'h3e57fcaa, 32'hbd5a859a} /* (28, 21, 8) {real, imag} */,
  {32'h3e867dec, 32'h3caecfe0} /* (28, 21, 7) {real, imag} */,
  {32'h3ee653ef, 32'hbd83885c} /* (28, 21, 6) {real, imag} */,
  {32'hbe2a9407, 32'hbf1a0495} /* (28, 21, 5) {real, imag} */,
  {32'hbdf3d62b, 32'hbe018fd1} /* (28, 21, 4) {real, imag} */,
  {32'h3de9f634, 32'h3cee5c8e} /* (28, 21, 3) {real, imag} */,
  {32'h3f0549c1, 32'h3c88c9d0} /* (28, 21, 2) {real, imag} */,
  {32'hbe68a1d9, 32'hbde4f526} /* (28, 21, 1) {real, imag} */,
  {32'hbf08439a, 32'h3eaabdb3} /* (28, 21, 0) {real, imag} */,
  {32'hbe221920, 32'hbed9fe70} /* (28, 20, 31) {real, imag} */,
  {32'h3c6fbf28, 32'h3ea4a17e} /* (28, 20, 30) {real, imag} */,
  {32'h3eb07ed0, 32'hbe484cc3} /* (28, 20, 29) {real, imag} */,
  {32'h3e23df49, 32'hbbbeadc0} /* (28, 20, 28) {real, imag} */,
  {32'hbe1331ac, 32'hbe8a04b6} /* (28, 20, 27) {real, imag} */,
  {32'h3e61bf44, 32'h3d10e632} /* (28, 20, 26) {real, imag} */,
  {32'hbd39de94, 32'h3ed253af} /* (28, 20, 25) {real, imag} */,
  {32'h3d5f4fb0, 32'hbe36bcd2} /* (28, 20, 24) {real, imag} */,
  {32'hbe7648f0, 32'h3ea89fe2} /* (28, 20, 23) {real, imag} */,
  {32'h3ee4d32f, 32'h3f1ca5da} /* (28, 20, 22) {real, imag} */,
  {32'hbda9e5ee, 32'hbea0e548} /* (28, 20, 21) {real, imag} */,
  {32'hbf037018, 32'h3d0196e8} /* (28, 20, 20) {real, imag} */,
  {32'h3f3e8bbf, 32'h3e1393d8} /* (28, 20, 19) {real, imag} */,
  {32'hbe64d25e, 32'h3ec78131} /* (28, 20, 18) {real, imag} */,
  {32'h3ddf60a0, 32'hbd455b34} /* (28, 20, 17) {real, imag} */,
  {32'hbeb6c43d, 32'hbe026191} /* (28, 20, 16) {real, imag} */,
  {32'hbdab66a6, 32'h3e8622f7} /* (28, 20, 15) {real, imag} */,
  {32'hbf171273, 32'h3dad14f3} /* (28, 20, 14) {real, imag} */,
  {32'h3e5e9f3a, 32'hbe425b30} /* (28, 20, 13) {real, imag} */,
  {32'hbdc4dc2f, 32'hbeca3908} /* (28, 20, 12) {real, imag} */,
  {32'hbeaf4610, 32'hbea09d9d} /* (28, 20, 11) {real, imag} */,
  {32'h3ecd3a36, 32'hbdb8b6b4} /* (28, 20, 10) {real, imag} */,
  {32'h3d95f4e6, 32'h3e11ce18} /* (28, 20, 9) {real, imag} */,
  {32'h3cbe4140, 32'hbee89164} /* (28, 20, 8) {real, imag} */,
  {32'hbf2009cc, 32'hbb02e100} /* (28, 20, 7) {real, imag} */,
  {32'hbebb795e, 32'h3dd48769} /* (28, 20, 6) {real, imag} */,
  {32'h3dbe4863, 32'hbf4e03cc} /* (28, 20, 5) {real, imag} */,
  {32'hbdb12e36, 32'hbebd2ac6} /* (28, 20, 4) {real, imag} */,
  {32'hbf62b6ec, 32'h3eb1ed29} /* (28, 20, 3) {real, imag} */,
  {32'h3d7fe810, 32'h3e2970a9} /* (28, 20, 2) {real, imag} */,
  {32'h3f4fa8a3, 32'hbd400996} /* (28, 20, 1) {real, imag} */,
  {32'h3dfd4b44, 32'h3eef620a} /* (28, 20, 0) {real, imag} */,
  {32'h3e0d3a78, 32'hbe863a06} /* (28, 19, 31) {real, imag} */,
  {32'h3dde71e0, 32'h3e8040d4} /* (28, 19, 30) {real, imag} */,
  {32'h3c9eecd8, 32'hbeab474a} /* (28, 19, 29) {real, imag} */,
  {32'hbdb74272, 32'hbe1ae311} /* (28, 19, 28) {real, imag} */,
  {32'hbe377ac0, 32'hbe51b29d} /* (28, 19, 27) {real, imag} */,
  {32'h3cba14b0, 32'h3e66befe} /* (28, 19, 26) {real, imag} */,
  {32'h3e1d9b08, 32'h3f22e6d6} /* (28, 19, 25) {real, imag} */,
  {32'h3eb87566, 32'hbe06c0f0} /* (28, 19, 24) {real, imag} */,
  {32'hbe17e621, 32'hbe12536a} /* (28, 19, 23) {real, imag} */,
  {32'hbed63aca, 32'h3e82af7e} /* (28, 19, 22) {real, imag} */,
  {32'hbd5082fa, 32'h3ea15a0a} /* (28, 19, 21) {real, imag} */,
  {32'h3eadba6f, 32'hbe3aad72} /* (28, 19, 20) {real, imag} */,
  {32'h3e9e1d8f, 32'hbeb3b659} /* (28, 19, 19) {real, imag} */,
  {32'h3e559864, 32'hbd6b6f02} /* (28, 19, 18) {real, imag} */,
  {32'hbe957eda, 32'h3ea9ff9a} /* (28, 19, 17) {real, imag} */,
  {32'h3de9ca40, 32'hbec6c9fa} /* (28, 19, 16) {real, imag} */,
  {32'h3e5b3344, 32'hbe355246} /* (28, 19, 15) {real, imag} */,
  {32'h3ee613ae, 32'hbe628aca} /* (28, 19, 14) {real, imag} */,
  {32'h3eebb879, 32'hbe13f7f5} /* (28, 19, 13) {real, imag} */,
  {32'hbe1f0147, 32'hbdcd2f90} /* (28, 19, 12) {real, imag} */,
  {32'hbe88f832, 32'h3ec9641b} /* (28, 19, 11) {real, imag} */,
  {32'hbcf9578c, 32'h3f13229c} /* (28, 19, 10) {real, imag} */,
  {32'hbe0a5a5c, 32'hbd349414} /* (28, 19, 9) {real, imag} */,
  {32'hbe32aa70, 32'hbc98a0c4} /* (28, 19, 8) {real, imag} */,
  {32'h3da4e457, 32'hbe916ccd} /* (28, 19, 7) {real, imag} */,
  {32'hbddab0fe, 32'h3ed108c0} /* (28, 19, 6) {real, imag} */,
  {32'h3f41c11e, 32'hbe0ac749} /* (28, 19, 5) {real, imag} */,
  {32'hbcb23af9, 32'h3e56ca14} /* (28, 19, 4) {real, imag} */,
  {32'h3ea2bed2, 32'h3e10b919} /* (28, 19, 3) {real, imag} */,
  {32'hbd0ed94e, 32'h3e0f3965} /* (28, 19, 2) {real, imag} */,
  {32'hbe9f1ae9, 32'hbd8f2fd2} /* (28, 19, 1) {real, imag} */,
  {32'h3e918098, 32'h3eb1f4a3} /* (28, 19, 0) {real, imag} */,
  {32'h3ddc2658, 32'h3d2b087c} /* (28, 18, 31) {real, imag} */,
  {32'hbe918f1e, 32'hbf3a58fb} /* (28, 18, 30) {real, imag} */,
  {32'h3d228614, 32'h3e0f1b03} /* (28, 18, 29) {real, imag} */,
  {32'hbe518b4f, 32'h3e8e4f0e} /* (28, 18, 28) {real, imag} */,
  {32'hbe8f9c2a, 32'hbe320a0b} /* (28, 18, 27) {real, imag} */,
  {32'hbe817e8d, 32'hbe966dd2} /* (28, 18, 26) {real, imag} */,
  {32'h3d3732b8, 32'h3e791b1c} /* (28, 18, 25) {real, imag} */,
  {32'hbe071a18, 32'h3ea90686} /* (28, 18, 24) {real, imag} */,
  {32'h3d739b58, 32'hbf557fb4} /* (28, 18, 23) {real, imag} */,
  {32'h3efe18b4, 32'hbdf2dca6} /* (28, 18, 22) {real, imag} */,
  {32'hbe486722, 32'hbdc48dbe} /* (28, 18, 21) {real, imag} */,
  {32'h3f1f44db, 32'h3deac9f2} /* (28, 18, 20) {real, imag} */,
  {32'hbdd098f6, 32'hbd65ad98} /* (28, 18, 19) {real, imag} */,
  {32'h3ed11c71, 32'hbda2535d} /* (28, 18, 18) {real, imag} */,
  {32'h3d962df0, 32'h3cfdbd04} /* (28, 18, 17) {real, imag} */,
  {32'hbe606173, 32'h3e8287bc} /* (28, 18, 16) {real, imag} */,
  {32'hbe81735f, 32'hbea5ebb0} /* (28, 18, 15) {real, imag} */,
  {32'h3e264842, 32'hbd680748} /* (28, 18, 14) {real, imag} */,
  {32'hbd93fd5c, 32'hbe4cec14} /* (28, 18, 13) {real, imag} */,
  {32'h3d05d6ab, 32'h3e304824} /* (28, 18, 12) {real, imag} */,
  {32'hbdbfc7a3, 32'hbea75896} /* (28, 18, 11) {real, imag} */,
  {32'hbdc6ca6b, 32'hbe507bf6} /* (28, 18, 10) {real, imag} */,
  {32'hbe2f2148, 32'h3e936113} /* (28, 18, 9) {real, imag} */,
  {32'h3dfcd028, 32'hbe25f1c1} /* (28, 18, 8) {real, imag} */,
  {32'h3e4e1ce9, 32'h3e1b572c} /* (28, 18, 7) {real, imag} */,
  {32'hbeaa1c5b, 32'h3ef3b9bf} /* (28, 18, 6) {real, imag} */,
  {32'h3f036424, 32'h3df98898} /* (28, 18, 5) {real, imag} */,
  {32'h3dee56ad, 32'h3f060f6a} /* (28, 18, 4) {real, imag} */,
  {32'hbe1584cd, 32'hbe45b62a} /* (28, 18, 3) {real, imag} */,
  {32'h3e9b33b2, 32'hbebba2b4} /* (28, 18, 2) {real, imag} */,
  {32'hbeb6aadc, 32'h3e899395} /* (28, 18, 1) {real, imag} */,
  {32'h3de381dc, 32'h3d78e32c} /* (28, 18, 0) {real, imag} */,
  {32'h3e0908d2, 32'hbd8da668} /* (28, 17, 31) {real, imag} */,
  {32'hbe874bc4, 32'h3e7547c6} /* (28, 17, 30) {real, imag} */,
  {32'h3e14472c, 32'h3e2e3736} /* (28, 17, 29) {real, imag} */,
  {32'hbed104ca, 32'hbe236437} /* (28, 17, 28) {real, imag} */,
  {32'hbc90eef0, 32'h3e8c0ca0} /* (28, 17, 27) {real, imag} */,
  {32'hbe1bd671, 32'hbf1a731e} /* (28, 17, 26) {real, imag} */,
  {32'h3ec959c3, 32'hbe222f77} /* (28, 17, 25) {real, imag} */,
  {32'h3efb4853, 32'h3e8018c5} /* (28, 17, 24) {real, imag} */,
  {32'hbe31b805, 32'h3e1ad822} /* (28, 17, 23) {real, imag} */,
  {32'hbe88d1dc, 32'hbe373272} /* (28, 17, 22) {real, imag} */,
  {32'hbe9b3bf7, 32'h3f14a21c} /* (28, 17, 21) {real, imag} */,
  {32'hbebda522, 32'h3e30127e} /* (28, 17, 20) {real, imag} */,
  {32'hbf0522dd, 32'hbe61e2f0} /* (28, 17, 19) {real, imag} */,
  {32'hbe4b0ac8, 32'h3e8626a3} /* (28, 17, 18) {real, imag} */,
  {32'h3de7165e, 32'hbe44fd14} /* (28, 17, 17) {real, imag} */,
  {32'h3e1b76cf, 32'h3e19b4ee} /* (28, 17, 16) {real, imag} */,
  {32'h3d183244, 32'h3cb886e8} /* (28, 17, 15) {real, imag} */,
  {32'hbe18aa4a, 32'h3cccf570} /* (28, 17, 14) {real, imag} */,
  {32'h3eacaf2e, 32'hbd138580} /* (28, 17, 13) {real, imag} */,
  {32'h3e8937a7, 32'hbd797b1a} /* (28, 17, 12) {real, imag} */,
  {32'h3eaf8660, 32'h3e291fad} /* (28, 17, 11) {real, imag} */,
  {32'hbd50c22c, 32'hbe70c642} /* (28, 17, 10) {real, imag} */,
  {32'h3d5179da, 32'hbd887cd8} /* (28, 17, 9) {real, imag} */,
  {32'h3e34c0a0, 32'h3cd9a21c} /* (28, 17, 8) {real, imag} */,
  {32'hbe822c66, 32'h3bf7f2a0} /* (28, 17, 7) {real, imag} */,
  {32'hbe89d54a, 32'hbdd4e458} /* (28, 17, 6) {real, imag} */,
  {32'h3d90aa27, 32'hbe347747} /* (28, 17, 5) {real, imag} */,
  {32'h3e0a2911, 32'h3dd1ed2a} /* (28, 17, 4) {real, imag} */,
  {32'h3ec54c12, 32'hbddc7b18} /* (28, 17, 3) {real, imag} */,
  {32'hbed7db43, 32'hbe105df3} /* (28, 17, 2) {real, imag} */,
  {32'h3dc91b52, 32'h3d4a728c} /* (28, 17, 1) {real, imag} */,
  {32'hbeaad55c, 32'h3e564d9d} /* (28, 17, 0) {real, imag} */,
  {32'hbc760160, 32'h3e93fac9} /* (28, 16, 31) {real, imag} */,
  {32'hbe9abf5c, 32'hbcfe3586} /* (28, 16, 30) {real, imag} */,
  {32'h3ea3fd33, 32'hbe248845} /* (28, 16, 29) {real, imag} */,
  {32'h3e200579, 32'h3e1cd382} /* (28, 16, 28) {real, imag} */,
  {32'h3d49b8f0, 32'hbe8e7545} /* (28, 16, 27) {real, imag} */,
  {32'h3e0912be, 32'hbe80fcd6} /* (28, 16, 26) {real, imag} */,
  {32'h3d7ef057, 32'hbd153c70} /* (28, 16, 25) {real, imag} */,
  {32'h3d161dda, 32'hbe9e1836} /* (28, 16, 24) {real, imag} */,
  {32'hbf027b7f, 32'hbe702b0f} /* (28, 16, 23) {real, imag} */,
  {32'h3f33d4e0, 32'h3e305d22} /* (28, 16, 22) {real, imag} */,
  {32'h3d91a196, 32'h3df4239c} /* (28, 16, 21) {real, imag} */,
  {32'h3e17510a, 32'h3e4404c9} /* (28, 16, 20) {real, imag} */,
  {32'h3e2dc39d, 32'h3d9ebd9a} /* (28, 16, 19) {real, imag} */,
  {32'hbdd9b85a, 32'hbdfcebc6} /* (28, 16, 18) {real, imag} */,
  {32'hbdab466c, 32'hbd499ec8} /* (28, 16, 17) {real, imag} */,
  {32'h3e843b32, 32'h00000000} /* (28, 16, 16) {real, imag} */,
  {32'hbdab466c, 32'h3d499ec8} /* (28, 16, 15) {real, imag} */,
  {32'hbdd9b85a, 32'h3dfcebc6} /* (28, 16, 14) {real, imag} */,
  {32'h3e2dc39d, 32'hbd9ebd9a} /* (28, 16, 13) {real, imag} */,
  {32'h3e17510a, 32'hbe4404c9} /* (28, 16, 12) {real, imag} */,
  {32'h3d91a196, 32'hbdf4239c} /* (28, 16, 11) {real, imag} */,
  {32'h3f33d4e0, 32'hbe305d22} /* (28, 16, 10) {real, imag} */,
  {32'hbf027b7f, 32'h3e702b0f} /* (28, 16, 9) {real, imag} */,
  {32'h3d161dda, 32'h3e9e1836} /* (28, 16, 8) {real, imag} */,
  {32'h3d7ef057, 32'h3d153c70} /* (28, 16, 7) {real, imag} */,
  {32'h3e0912be, 32'h3e80fcd6} /* (28, 16, 6) {real, imag} */,
  {32'h3d49b8f0, 32'h3e8e7545} /* (28, 16, 5) {real, imag} */,
  {32'h3e200579, 32'hbe1cd382} /* (28, 16, 4) {real, imag} */,
  {32'h3ea3fd33, 32'h3e248845} /* (28, 16, 3) {real, imag} */,
  {32'hbe9abf5c, 32'h3cfe3586} /* (28, 16, 2) {real, imag} */,
  {32'hbc760160, 32'hbe93fac9} /* (28, 16, 1) {real, imag} */,
  {32'hbeb0b84b, 32'h00000000} /* (28, 16, 0) {real, imag} */,
  {32'h3dc91b52, 32'hbd4a728c} /* (28, 15, 31) {real, imag} */,
  {32'hbed7db43, 32'h3e105df3} /* (28, 15, 30) {real, imag} */,
  {32'h3ec54c12, 32'h3ddc7b18} /* (28, 15, 29) {real, imag} */,
  {32'h3e0a2911, 32'hbdd1ed2a} /* (28, 15, 28) {real, imag} */,
  {32'h3d90aa27, 32'h3e347747} /* (28, 15, 27) {real, imag} */,
  {32'hbe89d54a, 32'h3dd4e458} /* (28, 15, 26) {real, imag} */,
  {32'hbe822c66, 32'hbbf7f2a0} /* (28, 15, 25) {real, imag} */,
  {32'h3e34c0a0, 32'hbcd9a21c} /* (28, 15, 24) {real, imag} */,
  {32'h3d5179da, 32'h3d887cd8} /* (28, 15, 23) {real, imag} */,
  {32'hbd50c22c, 32'h3e70c642} /* (28, 15, 22) {real, imag} */,
  {32'h3eaf8660, 32'hbe291fad} /* (28, 15, 21) {real, imag} */,
  {32'h3e8937a7, 32'h3d797b1a} /* (28, 15, 20) {real, imag} */,
  {32'h3eacaf2e, 32'h3d138580} /* (28, 15, 19) {real, imag} */,
  {32'hbe18aa4a, 32'hbcccf570} /* (28, 15, 18) {real, imag} */,
  {32'h3d183244, 32'hbcb886e8} /* (28, 15, 17) {real, imag} */,
  {32'h3e1b76cf, 32'hbe19b4ee} /* (28, 15, 16) {real, imag} */,
  {32'h3de7165e, 32'h3e44fd14} /* (28, 15, 15) {real, imag} */,
  {32'hbe4b0ac8, 32'hbe8626a3} /* (28, 15, 14) {real, imag} */,
  {32'hbf0522dd, 32'h3e61e2f0} /* (28, 15, 13) {real, imag} */,
  {32'hbebda522, 32'hbe30127e} /* (28, 15, 12) {real, imag} */,
  {32'hbe9b3bf7, 32'hbf14a21c} /* (28, 15, 11) {real, imag} */,
  {32'hbe88d1dc, 32'h3e373272} /* (28, 15, 10) {real, imag} */,
  {32'hbe31b805, 32'hbe1ad822} /* (28, 15, 9) {real, imag} */,
  {32'h3efb4853, 32'hbe8018c5} /* (28, 15, 8) {real, imag} */,
  {32'h3ec959c3, 32'h3e222f77} /* (28, 15, 7) {real, imag} */,
  {32'hbe1bd671, 32'h3f1a731e} /* (28, 15, 6) {real, imag} */,
  {32'hbc90eef0, 32'hbe8c0ca0} /* (28, 15, 5) {real, imag} */,
  {32'hbed104ca, 32'h3e236437} /* (28, 15, 4) {real, imag} */,
  {32'h3e14472c, 32'hbe2e3736} /* (28, 15, 3) {real, imag} */,
  {32'hbe874bc4, 32'hbe7547c6} /* (28, 15, 2) {real, imag} */,
  {32'h3e0908d2, 32'h3d8da668} /* (28, 15, 1) {real, imag} */,
  {32'hbeaad55c, 32'hbe564d9d} /* (28, 15, 0) {real, imag} */,
  {32'hbeb6aadc, 32'hbe899395} /* (28, 14, 31) {real, imag} */,
  {32'h3e9b33b2, 32'h3ebba2b4} /* (28, 14, 30) {real, imag} */,
  {32'hbe1584cd, 32'h3e45b62a} /* (28, 14, 29) {real, imag} */,
  {32'h3dee56ad, 32'hbf060f6a} /* (28, 14, 28) {real, imag} */,
  {32'h3f036424, 32'hbdf98898} /* (28, 14, 27) {real, imag} */,
  {32'hbeaa1c5b, 32'hbef3b9bf} /* (28, 14, 26) {real, imag} */,
  {32'h3e4e1ce9, 32'hbe1b572c} /* (28, 14, 25) {real, imag} */,
  {32'h3dfcd028, 32'h3e25f1c1} /* (28, 14, 24) {real, imag} */,
  {32'hbe2f2148, 32'hbe936113} /* (28, 14, 23) {real, imag} */,
  {32'hbdc6ca6b, 32'h3e507bf6} /* (28, 14, 22) {real, imag} */,
  {32'hbdbfc7a3, 32'h3ea75896} /* (28, 14, 21) {real, imag} */,
  {32'h3d05d6ab, 32'hbe304824} /* (28, 14, 20) {real, imag} */,
  {32'hbd93fd5c, 32'h3e4cec14} /* (28, 14, 19) {real, imag} */,
  {32'h3e264842, 32'h3d680748} /* (28, 14, 18) {real, imag} */,
  {32'hbe81735f, 32'h3ea5ebb0} /* (28, 14, 17) {real, imag} */,
  {32'hbe606173, 32'hbe8287bc} /* (28, 14, 16) {real, imag} */,
  {32'h3d962df0, 32'hbcfdbd04} /* (28, 14, 15) {real, imag} */,
  {32'h3ed11c71, 32'h3da2535d} /* (28, 14, 14) {real, imag} */,
  {32'hbdd098f6, 32'h3d65ad98} /* (28, 14, 13) {real, imag} */,
  {32'h3f1f44db, 32'hbdeac9f2} /* (28, 14, 12) {real, imag} */,
  {32'hbe486722, 32'h3dc48dbe} /* (28, 14, 11) {real, imag} */,
  {32'h3efe18b4, 32'h3df2dca6} /* (28, 14, 10) {real, imag} */,
  {32'h3d739b58, 32'h3f557fb4} /* (28, 14, 9) {real, imag} */,
  {32'hbe071a18, 32'hbea90686} /* (28, 14, 8) {real, imag} */,
  {32'h3d3732b8, 32'hbe791b1c} /* (28, 14, 7) {real, imag} */,
  {32'hbe817e8d, 32'h3e966dd2} /* (28, 14, 6) {real, imag} */,
  {32'hbe8f9c2a, 32'h3e320a0b} /* (28, 14, 5) {real, imag} */,
  {32'hbe518b4f, 32'hbe8e4f0e} /* (28, 14, 4) {real, imag} */,
  {32'h3d228614, 32'hbe0f1b03} /* (28, 14, 3) {real, imag} */,
  {32'hbe918f1e, 32'h3f3a58fb} /* (28, 14, 2) {real, imag} */,
  {32'h3ddc2658, 32'hbd2b087c} /* (28, 14, 1) {real, imag} */,
  {32'h3de381dc, 32'hbd78e32c} /* (28, 14, 0) {real, imag} */,
  {32'hbe9f1ae9, 32'h3d8f2fd2} /* (28, 13, 31) {real, imag} */,
  {32'hbd0ed94e, 32'hbe0f3965} /* (28, 13, 30) {real, imag} */,
  {32'h3ea2bed2, 32'hbe10b919} /* (28, 13, 29) {real, imag} */,
  {32'hbcb23af9, 32'hbe56ca14} /* (28, 13, 28) {real, imag} */,
  {32'h3f41c11e, 32'h3e0ac749} /* (28, 13, 27) {real, imag} */,
  {32'hbddab0fe, 32'hbed108c0} /* (28, 13, 26) {real, imag} */,
  {32'h3da4e457, 32'h3e916ccd} /* (28, 13, 25) {real, imag} */,
  {32'hbe32aa70, 32'h3c98a0c4} /* (28, 13, 24) {real, imag} */,
  {32'hbe0a5a5c, 32'h3d349414} /* (28, 13, 23) {real, imag} */,
  {32'hbcf9578c, 32'hbf13229c} /* (28, 13, 22) {real, imag} */,
  {32'hbe88f832, 32'hbec9641b} /* (28, 13, 21) {real, imag} */,
  {32'hbe1f0147, 32'h3dcd2f90} /* (28, 13, 20) {real, imag} */,
  {32'h3eebb879, 32'h3e13f7f5} /* (28, 13, 19) {real, imag} */,
  {32'h3ee613ae, 32'h3e628aca} /* (28, 13, 18) {real, imag} */,
  {32'h3e5b3344, 32'h3e355246} /* (28, 13, 17) {real, imag} */,
  {32'h3de9ca40, 32'h3ec6c9fa} /* (28, 13, 16) {real, imag} */,
  {32'hbe957eda, 32'hbea9ff9a} /* (28, 13, 15) {real, imag} */,
  {32'h3e559864, 32'h3d6b6f02} /* (28, 13, 14) {real, imag} */,
  {32'h3e9e1d8f, 32'h3eb3b659} /* (28, 13, 13) {real, imag} */,
  {32'h3eadba6f, 32'h3e3aad72} /* (28, 13, 12) {real, imag} */,
  {32'hbd5082fa, 32'hbea15a0a} /* (28, 13, 11) {real, imag} */,
  {32'hbed63aca, 32'hbe82af7e} /* (28, 13, 10) {real, imag} */,
  {32'hbe17e621, 32'h3e12536a} /* (28, 13, 9) {real, imag} */,
  {32'h3eb87566, 32'h3e06c0f0} /* (28, 13, 8) {real, imag} */,
  {32'h3e1d9b08, 32'hbf22e6d6} /* (28, 13, 7) {real, imag} */,
  {32'h3cba14b0, 32'hbe66befe} /* (28, 13, 6) {real, imag} */,
  {32'hbe377ac0, 32'h3e51b29d} /* (28, 13, 5) {real, imag} */,
  {32'hbdb74272, 32'h3e1ae311} /* (28, 13, 4) {real, imag} */,
  {32'h3c9eecd8, 32'h3eab474a} /* (28, 13, 3) {real, imag} */,
  {32'h3dde71e0, 32'hbe8040d4} /* (28, 13, 2) {real, imag} */,
  {32'h3e0d3a78, 32'h3e863a06} /* (28, 13, 1) {real, imag} */,
  {32'h3e918098, 32'hbeb1f4a3} /* (28, 13, 0) {real, imag} */,
  {32'h3f4fa8a3, 32'h3d400996} /* (28, 12, 31) {real, imag} */,
  {32'h3d7fe810, 32'hbe2970a9} /* (28, 12, 30) {real, imag} */,
  {32'hbf62b6ec, 32'hbeb1ed29} /* (28, 12, 29) {real, imag} */,
  {32'hbdb12e36, 32'h3ebd2ac6} /* (28, 12, 28) {real, imag} */,
  {32'h3dbe4863, 32'h3f4e03cc} /* (28, 12, 27) {real, imag} */,
  {32'hbebb795e, 32'hbdd48769} /* (28, 12, 26) {real, imag} */,
  {32'hbf2009cc, 32'h3b02e100} /* (28, 12, 25) {real, imag} */,
  {32'h3cbe4140, 32'h3ee89164} /* (28, 12, 24) {real, imag} */,
  {32'h3d95f4e6, 32'hbe11ce18} /* (28, 12, 23) {real, imag} */,
  {32'h3ecd3a36, 32'h3db8b6b4} /* (28, 12, 22) {real, imag} */,
  {32'hbeaf4610, 32'h3ea09d9d} /* (28, 12, 21) {real, imag} */,
  {32'hbdc4dc2f, 32'h3eca3908} /* (28, 12, 20) {real, imag} */,
  {32'h3e5e9f3a, 32'h3e425b30} /* (28, 12, 19) {real, imag} */,
  {32'hbf171273, 32'hbdad14f3} /* (28, 12, 18) {real, imag} */,
  {32'hbdab66a6, 32'hbe8622f7} /* (28, 12, 17) {real, imag} */,
  {32'hbeb6c43d, 32'h3e026191} /* (28, 12, 16) {real, imag} */,
  {32'h3ddf60a0, 32'h3d455b34} /* (28, 12, 15) {real, imag} */,
  {32'hbe64d25e, 32'hbec78131} /* (28, 12, 14) {real, imag} */,
  {32'h3f3e8bbf, 32'hbe1393d8} /* (28, 12, 13) {real, imag} */,
  {32'hbf037018, 32'hbd0196e8} /* (28, 12, 12) {real, imag} */,
  {32'hbda9e5ee, 32'h3ea0e548} /* (28, 12, 11) {real, imag} */,
  {32'h3ee4d32f, 32'hbf1ca5da} /* (28, 12, 10) {real, imag} */,
  {32'hbe7648f0, 32'hbea89fe2} /* (28, 12, 9) {real, imag} */,
  {32'h3d5f4fb0, 32'h3e36bcd2} /* (28, 12, 8) {real, imag} */,
  {32'hbd39de94, 32'hbed253af} /* (28, 12, 7) {real, imag} */,
  {32'h3e61bf44, 32'hbd10e632} /* (28, 12, 6) {real, imag} */,
  {32'hbe1331ac, 32'h3e8a04b6} /* (28, 12, 5) {real, imag} */,
  {32'h3e23df49, 32'h3bbeadc0} /* (28, 12, 4) {real, imag} */,
  {32'h3eb07ed0, 32'h3e484cc3} /* (28, 12, 3) {real, imag} */,
  {32'h3c6fbf28, 32'hbea4a17e} /* (28, 12, 2) {real, imag} */,
  {32'hbe221920, 32'h3ed9fe70} /* (28, 12, 1) {real, imag} */,
  {32'h3dfd4b44, 32'hbeef620a} /* (28, 12, 0) {real, imag} */,
  {32'hbe68a1d9, 32'h3de4f526} /* (28, 11, 31) {real, imag} */,
  {32'h3f0549c1, 32'hbc88c9d0} /* (28, 11, 30) {real, imag} */,
  {32'h3de9f634, 32'hbcee5c8e} /* (28, 11, 29) {real, imag} */,
  {32'hbdf3d62b, 32'h3e018fd1} /* (28, 11, 28) {real, imag} */,
  {32'hbe2a9407, 32'h3f1a0495} /* (28, 11, 27) {real, imag} */,
  {32'h3ee653ef, 32'h3d83885c} /* (28, 11, 26) {real, imag} */,
  {32'h3e867dec, 32'hbcaecfe0} /* (28, 11, 25) {real, imag} */,
  {32'h3e57fcaa, 32'h3d5a859a} /* (28, 11, 24) {real, imag} */,
  {32'hbe59b0f4, 32'hbef4ea66} /* (28, 11, 23) {real, imag} */,
  {32'h3e1a2862, 32'h3e1e350c} /* (28, 11, 22) {real, imag} */,
  {32'h3e70c3a4, 32'h3ea40018} /* (28, 11, 21) {real, imag} */,
  {32'hbf1a5bae, 32'hbcc7b6d0} /* (28, 11, 20) {real, imag} */,
  {32'hbe4c8d13, 32'h3d645ddc} /* (28, 11, 19) {real, imag} */,
  {32'hbe8105b2, 32'hbe1a19e0} /* (28, 11, 18) {real, imag} */,
  {32'h3db9cd71, 32'h3d5cb90c} /* (28, 11, 17) {real, imag} */,
  {32'hbe070568, 32'h3e5ee0f6} /* (28, 11, 16) {real, imag} */,
  {32'h3e9f2511, 32'h3e030764} /* (28, 11, 15) {real, imag} */,
  {32'h3f0b6103, 32'h3cbf0444} /* (28, 11, 14) {real, imag} */,
  {32'h3e03f9e7, 32'h3de232f8} /* (28, 11, 13) {real, imag} */,
  {32'hbcd3d770, 32'h3cef0cc0} /* (28, 11, 12) {real, imag} */,
  {32'hbe4e6e32, 32'h3eaba89a} /* (28, 11, 11) {real, imag} */,
  {32'h3ea021d5, 32'h3ea3b569} /* (28, 11, 10) {real, imag} */,
  {32'h3ee42a99, 32'h3e7c7356} /* (28, 11, 9) {real, imag} */,
  {32'h3e3482b0, 32'hbebfd110} /* (28, 11, 8) {real, imag} */,
  {32'hbabbbb00, 32'hbe4c2418} /* (28, 11, 7) {real, imag} */,
  {32'hbea449da, 32'h3f36cd14} /* (28, 11, 6) {real, imag} */,
  {32'h3f499cfc, 32'h3de58230} /* (28, 11, 5) {real, imag} */,
  {32'hbeab68c8, 32'hbf15e4b6} /* (28, 11, 4) {real, imag} */,
  {32'h3e5abaf9, 32'h3f17473b} /* (28, 11, 3) {real, imag} */,
  {32'hbe9dbfd5, 32'h3f6d76ae} /* (28, 11, 2) {real, imag} */,
  {32'hbe3c8e69, 32'hbf16f4b7} /* (28, 11, 1) {real, imag} */,
  {32'hbf08439a, 32'hbeaabdb3} /* (28, 11, 0) {real, imag} */,
  {32'h3ea06018, 32'h3eae1fc9} /* (28, 10, 31) {real, imag} */,
  {32'h3dd4083f, 32'hbf087439} /* (28, 10, 30) {real, imag} */,
  {32'hbdcbed66, 32'h3dfd8934} /* (28, 10, 29) {real, imag} */,
  {32'h3d90ffc2, 32'hbeb59732} /* (28, 10, 28) {real, imag} */,
  {32'hbee0849e, 32'hbe781126} /* (28, 10, 27) {real, imag} */,
  {32'h3eb4f770, 32'h3e06a1a8} /* (28, 10, 26) {real, imag} */,
  {32'h3c3798e0, 32'hbedd496d} /* (28, 10, 25) {real, imag} */,
  {32'hbea3c06b, 32'hbd837fd8} /* (28, 10, 24) {real, imag} */,
  {32'h3e81690e, 32'h3cbe9c3e} /* (28, 10, 23) {real, imag} */,
  {32'hbd9ce48a, 32'h3e92992f} /* (28, 10, 22) {real, imag} */,
  {32'h3d8d501c, 32'hbf066cbb} /* (28, 10, 21) {real, imag} */,
  {32'h3da0534c, 32'hbe786116} /* (28, 10, 20) {real, imag} */,
  {32'hbe4f6344, 32'h3e897bf8} /* (28, 10, 19) {real, imag} */,
  {32'h3ee99b1a, 32'hbe4758ca} /* (28, 10, 18) {real, imag} */,
  {32'h3e680d20, 32'hbe429620} /* (28, 10, 17) {real, imag} */,
  {32'h3e1000c8, 32'h3e0d82e0} /* (28, 10, 16) {real, imag} */,
  {32'hbdafd18c, 32'hbe611de1} /* (28, 10, 15) {real, imag} */,
  {32'hbf07b31a, 32'hbe1a5459} /* (28, 10, 14) {real, imag} */,
  {32'h3e37d593, 32'hbe07cb1c} /* (28, 10, 13) {real, imag} */,
  {32'h3be39680, 32'hbef092d8} /* (28, 10, 12) {real, imag} */,
  {32'hbe82966a, 32'h3cfde54c} /* (28, 10, 11) {real, imag} */,
  {32'hbd04cebc, 32'h3e9e74a2} /* (28, 10, 10) {real, imag} */,
  {32'h3e9fa5d4, 32'h3e6e7f0d} /* (28, 10, 9) {real, imag} */,
  {32'hbf46edfa, 32'h3e280a21} /* (28, 10, 8) {real, imag} */,
  {32'h3e176aba, 32'h3e387c6e} /* (28, 10, 7) {real, imag} */,
  {32'hbd904988, 32'h3c4a9fa0} /* (28, 10, 6) {real, imag} */,
  {32'hbef0a6ab, 32'hbe965dbe} /* (28, 10, 5) {real, imag} */,
  {32'h3ed0bca4, 32'h3e32b845} /* (28, 10, 4) {real, imag} */,
  {32'hbc224bc0, 32'hbe56acd9} /* (28, 10, 3) {real, imag} */,
  {32'hbf032239, 32'hbcc8a720} /* (28, 10, 2) {real, imag} */,
  {32'h3e0a17ea, 32'h3dca38fb} /* (28, 10, 1) {real, imag} */,
  {32'h3d7cfb4c, 32'h3ec6fb89} /* (28, 10, 0) {real, imag} */,
  {32'hbf32bf8d, 32'h3f66e5c8} /* (28, 9, 31) {real, imag} */,
  {32'h3f4342b2, 32'hbf7bff59} /* (28, 9, 30) {real, imag} */,
  {32'hbe1988fe, 32'hbdf2de1c} /* (28, 9, 29) {real, imag} */,
  {32'h3ca10a2c, 32'h3e4e5360} /* (28, 9, 28) {real, imag} */,
  {32'hbeb69914, 32'hbf0782b7} /* (28, 9, 27) {real, imag} */,
  {32'hbe949a26, 32'h3ee75a9c} /* (28, 9, 26) {real, imag} */,
  {32'h3e4e2565, 32'h3e69ab3e} /* (28, 9, 25) {real, imag} */,
  {32'hbdf8260a, 32'h3ec16772} /* (28, 9, 24) {real, imag} */,
  {32'h3e278eea, 32'h3e7b8fc8} /* (28, 9, 23) {real, imag} */,
  {32'hbe0bd5e4, 32'hbddbab9c} /* (28, 9, 22) {real, imag} */,
  {32'hbf3f00f3, 32'hbef95fbb} /* (28, 9, 21) {real, imag} */,
  {32'h3e3b1284, 32'hbdd632d6} /* (28, 9, 20) {real, imag} */,
  {32'hbee5df9b, 32'h3ee59258} /* (28, 9, 19) {real, imag} */,
  {32'h3e547c06, 32'h3e593c95} /* (28, 9, 18) {real, imag} */,
  {32'hbdefb6fa, 32'hbe14fd19} /* (28, 9, 17) {real, imag} */,
  {32'h3ed77184, 32'h3ecdd3be} /* (28, 9, 16) {real, imag} */,
  {32'h3e943200, 32'h3e173744} /* (28, 9, 15) {real, imag} */,
  {32'hbd704682, 32'h3e862cf3} /* (28, 9, 14) {real, imag} */,
  {32'h3ded1168, 32'hbe085f9a} /* (28, 9, 13) {real, imag} */,
  {32'hbd2f8006, 32'h3df5dfb2} /* (28, 9, 12) {real, imag} */,
  {32'hbe9ce7f6, 32'hbe9794a5} /* (28, 9, 11) {real, imag} */,
  {32'h3d70f540, 32'h3ddaf5aa} /* (28, 9, 10) {real, imag} */,
  {32'hbcb38978, 32'h3e17d866} /* (28, 9, 9) {real, imag} */,
  {32'h3e3fa574, 32'hbf12cbe6} /* (28, 9, 8) {real, imag} */,
  {32'h3e5606be, 32'h3de74f8c} /* (28, 9, 7) {real, imag} */,
  {32'hbe766202, 32'h3d4d4cb6} /* (28, 9, 6) {real, imag} */,
  {32'hbe220c90, 32'h3ee63c13} /* (28, 9, 5) {real, imag} */,
  {32'h3edb7e9a, 32'hbdea473e} /* (28, 9, 4) {real, imag} */,
  {32'hbe35698b, 32'hbdf3ca38} /* (28, 9, 3) {real, imag} */,
  {32'h3f6c98a6, 32'hbe7add06} /* (28, 9, 2) {real, imag} */,
  {32'h3eae7387, 32'h3d5e6f48} /* (28, 9, 1) {real, imag} */,
  {32'hbf2c50ea, 32'h3ee0da6f} /* (28, 9, 0) {real, imag} */,
  {32'hbff28c1c, 32'hbecb2b93} /* (28, 8, 31) {real, imag} */,
  {32'h3f95138a, 32'h3f1dfc39} /* (28, 8, 30) {real, imag} */,
  {32'h3f5ca3b4, 32'hbf086d6e} /* (28, 8, 29) {real, imag} */,
  {32'hbf19b2ab, 32'hbc215aec} /* (28, 8, 28) {real, imag} */,
  {32'hbf728792, 32'hbe4e4eb0} /* (28, 8, 27) {real, imag} */,
  {32'h3cac371c, 32'h3d7a7c24} /* (28, 8, 26) {real, imag} */,
  {32'h3da34b92, 32'hbea6f9ba} /* (28, 8, 25) {real, imag} */,
  {32'hbe830f86, 32'h3e4daa41} /* (28, 8, 24) {real, imag} */,
  {32'h3da86ea0, 32'hbf097cde} /* (28, 8, 23) {real, imag} */,
  {32'hbc040640, 32'h3dc5824e} /* (28, 8, 22) {real, imag} */,
  {32'h3ec581e2, 32'hbe06f76a} /* (28, 8, 21) {real, imag} */,
  {32'h3d414118, 32'hbe5df628} /* (28, 8, 20) {real, imag} */,
  {32'h3eea423c, 32'hbeebf5fe} /* (28, 8, 19) {real, imag} */,
  {32'h3e26b263, 32'h3d579c27} /* (28, 8, 18) {real, imag} */,
  {32'hbec94cd6, 32'h3ddbf3aa} /* (28, 8, 17) {real, imag} */,
  {32'hbc7180fc, 32'hbead6cde} /* (28, 8, 16) {real, imag} */,
  {32'h3e3d625e, 32'h3e2f0488} /* (28, 8, 15) {real, imag} */,
  {32'h3dcd34de, 32'h3e675e9c} /* (28, 8, 14) {real, imag} */,
  {32'hbe3697b5, 32'hbe098519} /* (28, 8, 13) {real, imag} */,
  {32'hbe529a4c, 32'h3ea1a934} /* (28, 8, 12) {real, imag} */,
  {32'h3e8ad7be, 32'h3e1bf843} /* (28, 8, 11) {real, imag} */,
  {32'h3ed9a0b2, 32'h3eb92e61} /* (28, 8, 10) {real, imag} */,
  {32'hbdfdb988, 32'h3e514cc2} /* (28, 8, 9) {real, imag} */,
  {32'h3d52e5f0, 32'hbe346c7a} /* (28, 8, 8) {real, imag} */,
  {32'hbe1e2ad4, 32'hbf567ca9} /* (28, 8, 7) {real, imag} */,
  {32'h3e8acda3, 32'hbea5ba40} /* (28, 8, 6) {real, imag} */,
  {32'h3edeb9fe, 32'h3d90fe70} /* (28, 8, 5) {real, imag} */,
  {32'h3f13f97d, 32'hbf01ebd8} /* (28, 8, 4) {real, imag} */,
  {32'h3b95a910, 32'h3f0b78fe} /* (28, 8, 3) {real, imag} */,
  {32'h3d822cd4, 32'hbd89635e} /* (28, 8, 2) {real, imag} */,
  {32'hbf1f16fe, 32'hbf406398} /* (28, 8, 1) {real, imag} */,
  {32'hbf1e7bf5, 32'hbf063c77} /* (28, 8, 0) {real, imag} */,
  {32'hbee2a2c5, 32'h3dc49763} /* (28, 7, 31) {real, imag} */,
  {32'hbeaab9d3, 32'h3ef4c624} /* (28, 7, 30) {real, imag} */,
  {32'hbd13d1a0, 32'hbe0f31f1} /* (28, 7, 29) {real, imag} */,
  {32'hbe2946a7, 32'hbee97dd1} /* (28, 7, 28) {real, imag} */,
  {32'hbf253250, 32'h3f0ad63f} /* (28, 7, 27) {real, imag} */,
  {32'hbe8809b7, 32'hbeccea20} /* (28, 7, 26) {real, imag} */,
  {32'hbe35d977, 32'h3ec61cc3} /* (28, 7, 25) {real, imag} */,
  {32'hbedcaef2, 32'h3e046b15} /* (28, 7, 24) {real, imag} */,
  {32'hbe0868c6, 32'hbe9e684c} /* (28, 7, 23) {real, imag} */,
  {32'hbe90217d, 32'hbf22ab31} /* (28, 7, 22) {real, imag} */,
  {32'h3cdefc88, 32'h3edc7ef8} /* (28, 7, 21) {real, imag} */,
  {32'hbdd8a26f, 32'hbefdacbf} /* (28, 7, 20) {real, imag} */,
  {32'h3ef5da1a, 32'h3dfecdee} /* (28, 7, 19) {real, imag} */,
  {32'hbe70a5b5, 32'h3e2f31b5} /* (28, 7, 18) {real, imag} */,
  {32'hbd69ef76, 32'hbda527be} /* (28, 7, 17) {real, imag} */,
  {32'hbdaaf9b4, 32'h3e94efc2} /* (28, 7, 16) {real, imag} */,
  {32'h3e9ca8a7, 32'hbc57fce0} /* (28, 7, 15) {real, imag} */,
  {32'h3ebd555a, 32'hbe703682} /* (28, 7, 14) {real, imag} */,
  {32'hbee5cd5a, 32'h3d696304} /* (28, 7, 13) {real, imag} */,
  {32'hbdf46f60, 32'h3d7d9f48} /* (28, 7, 12) {real, imag} */,
  {32'hbdbe3264, 32'hbee19751} /* (28, 7, 11) {real, imag} */,
  {32'hbcffb334, 32'hbe365b9e} /* (28, 7, 10) {real, imag} */,
  {32'hbe4789c4, 32'hbd852f2a} /* (28, 7, 9) {real, imag} */,
  {32'hbe95c0fa, 32'hbf0f20e6} /* (28, 7, 8) {real, imag} */,
  {32'h3eec5cd6, 32'h3eb5bfe3} /* (28, 7, 7) {real, imag} */,
  {32'hbe6f16e4, 32'hbdc5746b} /* (28, 7, 6) {real, imag} */,
  {32'h3e63469c, 32'hbd1adb18} /* (28, 7, 5) {real, imag} */,
  {32'hbde310c4, 32'h3e84a790} /* (28, 7, 4) {real, imag} */,
  {32'hbf0ea72a, 32'h3f04f07a} /* (28, 7, 3) {real, imag} */,
  {32'hbecc56b0, 32'h3e6f60a3} /* (28, 7, 2) {real, imag} */,
  {32'h3f754ef2, 32'h3ea3ccd3} /* (28, 7, 1) {real, imag} */,
  {32'h3fa2f657, 32'h3dfc1c54} /* (28, 7, 0) {real, imag} */,
  {32'hbf251b2e, 32'hbc8f16f0} /* (28, 6, 31) {real, imag} */,
  {32'h3f244c66, 32'h3f262a9c} /* (28, 6, 30) {real, imag} */,
  {32'h3ebc8296, 32'h3ea5708d} /* (28, 6, 29) {real, imag} */,
  {32'hbe128b16, 32'hbeceb5da} /* (28, 6, 28) {real, imag} */,
  {32'hbf311803, 32'hbe5403c1} /* (28, 6, 27) {real, imag} */,
  {32'h3eaf2d98, 32'hbd77fc68} /* (28, 6, 26) {real, imag} */,
  {32'h3e53b6f0, 32'h3efd03bc} /* (28, 6, 25) {real, imag} */,
  {32'h3e588c08, 32'h3f2ba1e5} /* (28, 6, 24) {real, imag} */,
  {32'h3d54e3c4, 32'hbdd95322} /* (28, 6, 23) {real, imag} */,
  {32'h3ddd1eb2, 32'h3e9a2f64} /* (28, 6, 22) {real, imag} */,
  {32'h3c2e24d0, 32'hbdf44f74} /* (28, 6, 21) {real, imag} */,
  {32'h3ea4a72c, 32'h3dc8d146} /* (28, 6, 20) {real, imag} */,
  {32'h3e0e56cb, 32'hbebd70b8} /* (28, 6, 19) {real, imag} */,
  {32'hbe944c0e, 32'h3d62ea7a} /* (28, 6, 18) {real, imag} */,
  {32'h3e7e5a48, 32'h3ddd92d4} /* (28, 6, 17) {real, imag} */,
  {32'hbd8b5341, 32'hbee8dd12} /* (28, 6, 16) {real, imag} */,
  {32'h3dd0d53f, 32'h3e2819f4} /* (28, 6, 15) {real, imag} */,
  {32'hbdbb76bc, 32'hbdebca14} /* (28, 6, 14) {real, imag} */,
  {32'hbdfcedd8, 32'h3ee60a54} /* (28, 6, 13) {real, imag} */,
  {32'h3e39fe10, 32'hbdbd548c} /* (28, 6, 12) {real, imag} */,
  {32'h3f064051, 32'hbd548410} /* (28, 6, 11) {real, imag} */,
  {32'hbefe4aae, 32'h3ec43ff2} /* (28, 6, 10) {real, imag} */,
  {32'h3ead0edc, 32'hbed1388c} /* (28, 6, 9) {real, imag} */,
  {32'hbd5aa980, 32'hbf1d89ba} /* (28, 6, 8) {real, imag} */,
  {32'h3f433aa0, 32'h3f03f672} /* (28, 6, 7) {real, imag} */,
  {32'hbea8d14f, 32'h3eb1d618} /* (28, 6, 6) {real, imag} */,
  {32'hbe0edf2f, 32'hbaf837c0} /* (28, 6, 5) {real, imag} */,
  {32'h3e6370ce, 32'h3db416b8} /* (28, 6, 4) {real, imag} */,
  {32'h3e927e10, 32'h3e5a764b} /* (28, 6, 3) {real, imag} */,
  {32'h3e4a8dbc, 32'hbc051f08} /* (28, 6, 2) {real, imag} */,
  {32'hbf0b3c59, 32'hbea1aa63} /* (28, 6, 1) {real, imag} */,
  {32'hbda41964, 32'h3ee3cbaa} /* (28, 6, 0) {real, imag} */,
  {32'hc055b67a, 32'hbf3b7554} /* (28, 5, 31) {real, imag} */,
  {32'h3f05815e, 32'hbe87527e} /* (28, 5, 30) {real, imag} */,
  {32'h3e136b43, 32'hbf4181aa} /* (28, 5, 29) {real, imag} */,
  {32'hbf1e8c5a, 32'h3e08a5c8} /* (28, 5, 28) {real, imag} */,
  {32'h3f94909c, 32'h3e5d58af} /* (28, 5, 27) {real, imag} */,
  {32'h3ecba2aa, 32'hbf2832d4} /* (28, 5, 26) {real, imag} */,
  {32'h3ee5f15d, 32'h3f27feae} /* (28, 5, 25) {real, imag} */,
  {32'h3d925730, 32'hbdb9732f} /* (28, 5, 24) {real, imag} */,
  {32'h3e84279e, 32'h3e3016d9} /* (28, 5, 23) {real, imag} */,
  {32'h3e91e984, 32'h3d6cf340} /* (28, 5, 22) {real, imag} */,
  {32'h3eae30f6, 32'hbecc6f27} /* (28, 5, 21) {real, imag} */,
  {32'h3c2a8f78, 32'hbd427362} /* (28, 5, 20) {real, imag} */,
  {32'hbe969420, 32'h3d5c67a0} /* (28, 5, 19) {real, imag} */,
  {32'hbd7ada94, 32'h3e98b7c9} /* (28, 5, 18) {real, imag} */,
  {32'hbd1b95e8, 32'hbf031d68} /* (28, 5, 17) {real, imag} */,
  {32'hbd6690c3, 32'hbe302633} /* (28, 5, 16) {real, imag} */,
  {32'hbd985527, 32'h3e8e20b4} /* (28, 5, 15) {real, imag} */,
  {32'hbdf51552, 32'h3e0ff4c6} /* (28, 5, 14) {real, imag} */,
  {32'hbd89a5ca, 32'hbdafa0cc} /* (28, 5, 13) {real, imag} */,
  {32'h3e75ef3b, 32'hbe5d6a0a} /* (28, 5, 12) {real, imag} */,
  {32'hbdec5adc, 32'h3e68cee0} /* (28, 5, 11) {real, imag} */,
  {32'hbe5ccc51, 32'hbee532ad} /* (28, 5, 10) {real, imag} */,
  {32'h3e947aa6, 32'hbf00c0eb} /* (28, 5, 9) {real, imag} */,
  {32'h3c279cbc, 32'h3eb82bf8} /* (28, 5, 8) {real, imag} */,
  {32'h3d359c66, 32'h3e9f0d35} /* (28, 5, 7) {real, imag} */,
  {32'hbdba380e, 32'h3d9d063c} /* (28, 5, 6) {real, imag} */,
  {32'h3f21eb24, 32'h3f4e45cd} /* (28, 5, 5) {real, imag} */,
  {32'h3ddeccb8, 32'h3f21b553} /* (28, 5, 4) {real, imag} */,
  {32'hbeb86856, 32'hbf2153dc} /* (28, 5, 3) {real, imag} */,
  {32'h3f5d4471, 32'hbf594585} /* (28, 5, 2) {real, imag} */,
  {32'hc0142d54, 32'hbfd087b0} /* (28, 5, 1) {real, imag} */,
  {32'hbff36a56, 32'hbf9e2570} /* (28, 5, 0) {real, imag} */,
  {32'h4002ba56, 32'h400cc1ba} /* (28, 4, 31) {real, imag} */,
  {32'hc0085c64, 32'hbfba225d} /* (28, 4, 30) {real, imag} */,
  {32'h3e3e0f14, 32'hbd9291f4} /* (28, 4, 29) {real, imag} */,
  {32'h3f813465, 32'hbe94d7c5} /* (28, 4, 28) {real, imag} */,
  {32'hbde7cb7f, 32'h3e272a54} /* (28, 4, 27) {real, imag} */,
  {32'h3f02e4c3, 32'h3ef4cc02} /* (28, 4, 26) {real, imag} */,
  {32'h3e8cca1c, 32'hbeab05ac} /* (28, 4, 25) {real, imag} */,
  {32'hbeca3c29, 32'h3d9d77fb} /* (28, 4, 24) {real, imag} */,
  {32'hbefeac1b, 32'h3e2930be} /* (28, 4, 23) {real, imag} */,
  {32'hbe8ad9fd, 32'h3e141e22} /* (28, 4, 22) {real, imag} */,
  {32'hbf236ae0, 32'h3e4daa93} /* (28, 4, 21) {real, imag} */,
  {32'h3f3b9cca, 32'hbebc2635} /* (28, 4, 20) {real, imag} */,
  {32'hbcff2968, 32'hbd8e6de5} /* (28, 4, 19) {real, imag} */,
  {32'h3ca8abe8, 32'h3e089076} /* (28, 4, 18) {real, imag} */,
  {32'hbdbbc62e, 32'h3de235a0} /* (28, 4, 17) {real, imag} */,
  {32'h3db2c1a2, 32'hbdab470d} /* (28, 4, 16) {real, imag} */,
  {32'hbea14080, 32'h3ea3fe6d} /* (28, 4, 15) {real, imag} */,
  {32'hbe3d3b40, 32'h3d9d4bc6} /* (28, 4, 14) {real, imag} */,
  {32'h3deeec6e, 32'h3e4a7927} /* (28, 4, 13) {real, imag} */,
  {32'h3e021d9c, 32'hbf1e1e44} /* (28, 4, 12) {real, imag} */,
  {32'h3ddbd804, 32'h3ecf20ad} /* (28, 4, 11) {real, imag} */,
  {32'hbd84ea30, 32'h3e024f41} /* (28, 4, 10) {real, imag} */,
  {32'hbef840ee, 32'hbeab2690} /* (28, 4, 9) {real, imag} */,
  {32'h3d5705cf, 32'hbe842c3c} /* (28, 4, 8) {real, imag} */,
  {32'hbf09befe, 32'h3d907e14} /* (28, 4, 7) {real, imag} */,
  {32'hbd3f92e0, 32'h3f2b8bc5} /* (28, 4, 6) {real, imag} */,
  {32'h3e519af8, 32'hbeac549a} /* (28, 4, 5) {real, imag} */,
  {32'h3fbcd1c2, 32'hbf5339ac} /* (28, 4, 4) {real, imag} */,
  {32'h3f4aaf5d, 32'hbf867e75} /* (28, 4, 3) {real, imag} */,
  {32'hbfe7b92e, 32'hc0171cfb} /* (28, 4, 2) {real, imag} */,
  {32'h40649c41, 32'h4018f1ba} /* (28, 4, 1) {real, imag} */,
  {32'h3f8b550a, 32'h3fcf361d} /* (28, 4, 0) {real, imag} */,
  {32'hc0930f7f, 32'h3fa2f434} /* (28, 3, 31) {real, imag} */,
  {32'h4015b366, 32'hc03f95c8} /* (28, 3, 30) {real, imag} */,
  {32'hbf215212, 32'h3e6c96c6} /* (28, 3, 29) {real, imag} */,
  {32'h3ebdf34d, 32'h3f4e12ce} /* (28, 3, 28) {real, imag} */,
  {32'hbea83e50, 32'hbf69021b} /* (28, 3, 27) {real, imag} */,
  {32'h3f09f571, 32'hbd8f7f58} /* (28, 3, 26) {real, imag} */,
  {32'hbefa7386, 32'h3ed16e46} /* (28, 3, 25) {real, imag} */,
  {32'hbdf943ea, 32'hbf69089a} /* (28, 3, 24) {real, imag} */,
  {32'h3e8de770, 32'h3f02c896} /* (28, 3, 23) {real, imag} */,
  {32'h3f72ea15, 32'h3f877ad3} /* (28, 3, 22) {real, imag} */,
  {32'hbf1f03d1, 32'hbc75abc0} /* (28, 3, 21) {real, imag} */,
  {32'h3ed013f8, 32'hbd6a8bca} /* (28, 3, 20) {real, imag} */,
  {32'hbe732a1b, 32'hbe32d14f} /* (28, 3, 19) {real, imag} */,
  {32'h3df06cdc, 32'hbebfeffc} /* (28, 3, 18) {real, imag} */,
  {32'hbe2c6ec9, 32'hbe9f7e50} /* (28, 3, 17) {real, imag} */,
  {32'hbe8146e2, 32'h3c26fa20} /* (28, 3, 16) {real, imag} */,
  {32'h3e61b17c, 32'h3d4854e0} /* (28, 3, 15) {real, imag} */,
  {32'hbe0e4213, 32'hbd921e58} /* (28, 3, 14) {real, imag} */,
  {32'hbeeeccb0, 32'hbf22567f} /* (28, 3, 13) {real, imag} */,
  {32'hbe52c720, 32'hbf03d950} /* (28, 3, 12) {real, imag} */,
  {32'h3ed7585b, 32'hbef86ded} /* (28, 3, 11) {real, imag} */,
  {32'hbddabf1e, 32'h3e3b725c} /* (28, 3, 10) {real, imag} */,
  {32'hbe1ac983, 32'h3eea7ee3} /* (28, 3, 9) {real, imag} */,
  {32'h3d8e7b46, 32'hbe5e8a86} /* (28, 3, 8) {real, imag} */,
  {32'h3f0c29a3, 32'h3e854129} /* (28, 3, 7) {real, imag} */,
  {32'hbfd6890a, 32'hbf2326ad} /* (28, 3, 6) {real, imag} */,
  {32'h3f5510a9, 32'hbdd698e0} /* (28, 3, 5) {real, imag} */,
  {32'hbd84ecfc, 32'h3facba7a} /* (28, 3, 4) {real, imag} */,
  {32'h3f6276c6, 32'h3f00af85} /* (28, 3, 3) {real, imag} */,
  {32'hbefb7dbb, 32'hc0477516} /* (28, 3, 2) {real, imag} */,
  {32'h4013bb0d, 32'h40998610} /* (28, 3, 1) {real, imag} */,
  {32'h3f2fc724, 32'hbf037278} /* (28, 3, 0) {real, imag} */,
  {32'hc1a5e041, 32'h3f51e393} /* (28, 2, 31) {real, imag} */,
  {32'h4145513e, 32'hc09b8fb2} /* (28, 2, 30) {real, imag} */,
  {32'hbf0fec69, 32'hbe764a62} /* (28, 2, 29) {real, imag} */,
  {32'hbf485007, 32'h402efa3a} /* (28, 2, 28) {real, imag} */,
  {32'h3f591d94, 32'hbf688b18} /* (28, 2, 27) {real, imag} */,
  {32'h3f31fa1a, 32'h3f3fc7c6} /* (28, 2, 26) {real, imag} */,
  {32'hbd3658fa, 32'h3fac00c3} /* (28, 2, 25) {real, imag} */,
  {32'h3e19aa95, 32'hbfa48af4} /* (28, 2, 24) {real, imag} */,
  {32'h3e0152ed, 32'hbe668edf} /* (28, 2, 23) {real, imag} */,
  {32'h3f384a46, 32'h3db5454a} /* (28, 2, 22) {real, imag} */,
  {32'h3c113890, 32'hbf76fb7c} /* (28, 2, 21) {real, imag} */,
  {32'h3e3fd038, 32'hbe762b38} /* (28, 2, 20) {real, imag} */,
  {32'hbe5d4be1, 32'h3e987722} /* (28, 2, 19) {real, imag} */,
  {32'h3e90b6a0, 32'hbee3d349} /* (28, 2, 18) {real, imag} */,
  {32'hbe22ff02, 32'h3ef7f5b3} /* (28, 2, 17) {real, imag} */,
  {32'h3e82a39e, 32'hbdf3909e} /* (28, 2, 16) {real, imag} */,
  {32'hbe2e6e97, 32'h3e786131} /* (28, 2, 15) {real, imag} */,
  {32'h3d53b17e, 32'h3ecb86f1} /* (28, 2, 14) {real, imag} */,
  {32'hbdfcbe84, 32'h3e438fe1} /* (28, 2, 13) {real, imag} */,
  {32'hbe990331, 32'hbe3d0ec8} /* (28, 2, 12) {real, imag} */,
  {32'h3cdf00b8, 32'h3e40afd6} /* (28, 2, 11) {real, imag} */,
  {32'hbef9d68c, 32'hbe5814a0} /* (28, 2, 10) {real, imag} */,
  {32'h3e5d10dc, 32'h3f351a8e} /* (28, 2, 9) {real, imag} */,
  {32'h3f39549f, 32'h3f2bbf56} /* (28, 2, 8) {real, imag} */,
  {32'hbeb7df7c, 32'hbe600a9f} /* (28, 2, 7) {real, imag} */,
  {32'hbdf7b184, 32'hbdb1178c} /* (28, 2, 6) {real, imag} */,
  {32'h3fb2b837, 32'h3f5b6217} /* (28, 2, 5) {real, imag} */,
  {32'hc033813b, 32'hbf89fa5c} /* (28, 2, 4) {real, imag} */,
  {32'hbf0954e4, 32'hbd6781ec} /* (28, 2, 3) {real, imag} */,
  {32'h4117c4b4, 32'hc077ff4a} /* (28, 2, 2) {real, imag} */,
  {32'hc141e4c5, 32'h404a20c0} /* (28, 2, 1) {real, imag} */,
  {32'hc12f5eb5, 32'hc0199eaa} /* (28, 2, 0) {real, imag} */,
  {32'h418cc812, 32'hc0be7672} /* (28, 1, 31) {real, imag} */,
  {32'hc1036f90, 32'h3f9e4a7b} /* (28, 1, 30) {real, imag} */,
  {32'h3e17c6c0, 32'h3ea07c5e} /* (28, 1, 29) {real, imag} */,
  {32'h3fc26a2e, 32'h3f984bf4} /* (28, 1, 28) {real, imag} */,
  {32'hc05fa512, 32'h3f8113ad} /* (28, 1, 27) {real, imag} */,
  {32'hbf05e7f1, 32'h3dc1ae04} /* (28, 1, 26) {real, imag} */,
  {32'hbd1710c0, 32'hbf095d26} /* (28, 1, 25) {real, imag} */,
  {32'hbefdf928, 32'h3e7519ed} /* (28, 1, 24) {real, imag} */,
  {32'h3a521e00, 32'h3ebaa354} /* (28, 1, 23) {real, imag} */,
  {32'hbf1a26a2, 32'h3eb75566} /* (28, 1, 22) {real, imag} */,
  {32'hbee114bc, 32'h3d983bde} /* (28, 1, 21) {real, imag} */,
  {32'h3d8e97fe, 32'hbe1e0274} /* (28, 1, 20) {real, imag} */,
  {32'hbea21359, 32'h3c05bf20} /* (28, 1, 19) {real, imag} */,
  {32'h3dc34f80, 32'h3dc0008a} /* (28, 1, 18) {real, imag} */,
  {32'h3d6a361c, 32'h3e3c4fa0} /* (28, 1, 17) {real, imag} */,
  {32'h3d965326, 32'hbe2ed598} /* (28, 1, 16) {real, imag} */,
  {32'h3e121178, 32'h3ea50ee0} /* (28, 1, 15) {real, imag} */,
  {32'h3edc89a0, 32'hbf29389a} /* (28, 1, 14) {real, imag} */,
  {32'hbcbe7d64, 32'h3e8294c1} /* (28, 1, 13) {real, imag} */,
  {32'h3e1ef4c2, 32'hbe053a7b} /* (28, 1, 12) {real, imag} */,
  {32'hbe9b96d6, 32'h3e7ef79c} /* (28, 1, 11) {real, imag} */,
  {32'hbea8a226, 32'h3d9808ef} /* (28, 1, 10) {real, imag} */,
  {32'hbdba5e10, 32'hbe9e695c} /* (28, 1, 9) {real, imag} */,
  {32'h3d11aba8, 32'hbf3c0a80} /* (28, 1, 8) {real, imag} */,
  {32'hbefcf2b4, 32'h3f44bdc6} /* (28, 1, 7) {real, imag} */,
  {32'hbcef8a40, 32'hbeba8ec6} /* (28, 1, 6) {real, imag} */,
  {32'hc000a52d, 32'hbf6dc7c4} /* (28, 1, 5) {real, imag} */,
  {32'h3fb9a870, 32'h3e89da7e} /* (28, 1, 4) {real, imag} */,
  {32'hc002ece5, 32'hbc8ac020} /* (28, 1, 3) {real, imag} */,
  {32'hc13d1793, 32'hc149ec43} /* (28, 1, 2) {real, imag} */,
  {32'h41cdec3a, 32'h412fa2b3} /* (28, 1, 1) {real, imag} */,
  {32'h415cc76e, 32'h3ff21544} /* (28, 1, 0) {real, imag} */,
  {32'h40991d40, 32'hc0b37a0d} /* (28, 0, 31) {real, imag} */,
  {32'hc06e5408, 32'h40dd99ac} /* (28, 0, 30) {real, imag} */,
  {32'hbea5f894, 32'hbf3c5b31} /* (28, 0, 29) {real, imag} */,
  {32'hbdc2034c, 32'h3eff8618} /* (28, 0, 28) {real, imag} */,
  {32'hc01a31d0, 32'h3ed1935a} /* (28, 0, 27) {real, imag} */,
  {32'hbdc4d628, 32'hbe86606f} /* (28, 0, 26) {real, imag} */,
  {32'h3e6a5be4, 32'hbfaa1411} /* (28, 0, 25) {real, imag} */,
  {32'h3ee591a7, 32'h3e2e1464} /* (28, 0, 24) {real, imag} */,
  {32'h3dbdef34, 32'hbe8677e0} /* (28, 0, 23) {real, imag} */,
  {32'h3c053cf0, 32'hbd9a6088} /* (28, 0, 22) {real, imag} */,
  {32'hbee93342, 32'h3ee55b4c} /* (28, 0, 21) {real, imag} */,
  {32'h3ea23e35, 32'hbf01a746} /* (28, 0, 20) {real, imag} */,
  {32'hbe6bddfa, 32'hbea2b86e} /* (28, 0, 19) {real, imag} */,
  {32'hbd473d10, 32'hbe7ae38b} /* (28, 0, 18) {real, imag} */,
  {32'hbe257334, 32'h3e51bd7f} /* (28, 0, 17) {real, imag} */,
  {32'hbe4f6430, 32'h00000000} /* (28, 0, 16) {real, imag} */,
  {32'hbe257334, 32'hbe51bd7f} /* (28, 0, 15) {real, imag} */,
  {32'hbd473d10, 32'h3e7ae38b} /* (28, 0, 14) {real, imag} */,
  {32'hbe6bddfa, 32'h3ea2b86e} /* (28, 0, 13) {real, imag} */,
  {32'h3ea23e35, 32'h3f01a746} /* (28, 0, 12) {real, imag} */,
  {32'hbee93342, 32'hbee55b4c} /* (28, 0, 11) {real, imag} */,
  {32'h3c053cf0, 32'h3d9a6088} /* (28, 0, 10) {real, imag} */,
  {32'h3dbdef34, 32'h3e8677e0} /* (28, 0, 9) {real, imag} */,
  {32'h3ee591a7, 32'hbe2e1464} /* (28, 0, 8) {real, imag} */,
  {32'h3e6a5be4, 32'h3faa1411} /* (28, 0, 7) {real, imag} */,
  {32'hbdc4d628, 32'h3e86606f} /* (28, 0, 6) {real, imag} */,
  {32'hc01a31d0, 32'hbed1935a} /* (28, 0, 5) {real, imag} */,
  {32'hbdc2034c, 32'hbeff8618} /* (28, 0, 4) {real, imag} */,
  {32'hbea5f894, 32'h3f3c5b31} /* (28, 0, 3) {real, imag} */,
  {32'hc06e5408, 32'hc0dd99ac} /* (28, 0, 2) {real, imag} */,
  {32'h40991d40, 32'h40b37a0d} /* (28, 0, 1) {real, imag} */,
  {32'hc0678278, 32'h00000000} /* (28, 0, 0) {real, imag} */,
  {32'h4150e7c2, 32'hc0b24765} /* (27, 31, 31) {real, imag} */,
  {32'hc10eb0ba, 32'h410aeec8} /* (27, 31, 30) {real, imag} */,
  {32'hbfc2ca0c, 32'h3e9fcc40} /* (27, 31, 29) {real, imag} */,
  {32'h3f77485f, 32'hbf1830e3} /* (27, 31, 28) {real, imag} */,
  {32'hbfe28a12, 32'h3f61ba4d} /* (27, 31, 27) {real, imag} */,
  {32'hbe46a3e6, 32'h3ec1f8f7} /* (27, 31, 26) {real, imag} */,
  {32'hbf1960fd, 32'hbe8c7ef0} /* (27, 31, 25) {real, imag} */,
  {32'hbedb6946, 32'h3f7c1033} /* (27, 31, 24) {real, imag} */,
  {32'hbf3191f8, 32'h3ed74fff} /* (27, 31, 23) {real, imag} */,
  {32'hbc844ed0, 32'hbf32fc27} /* (27, 31, 22) {real, imag} */,
  {32'hbf0df652, 32'h3ecde1ac} /* (27, 31, 21) {real, imag} */,
  {32'hbeb213de, 32'hbd6b1ff4} /* (27, 31, 20) {real, imag} */,
  {32'h3f0823dd, 32'h3d10da8c} /* (27, 31, 19) {real, imag} */,
  {32'h3ed3acdd, 32'h3ef1b2f5} /* (27, 31, 18) {real, imag} */,
  {32'hbe9017c2, 32'hbeefa48c} /* (27, 31, 17) {real, imag} */,
  {32'hbe04dd01, 32'h3e05ad3f} /* (27, 31, 16) {real, imag} */,
  {32'hbc94e0e8, 32'hbe0538c1} /* (27, 31, 15) {real, imag} */,
  {32'h3ebbf42a, 32'hbe750aae} /* (27, 31, 14) {real, imag} */,
  {32'h3d3e4c1e, 32'h3f057a26} /* (27, 31, 13) {real, imag} */,
  {32'hbdc4237e, 32'hbf2d64e8} /* (27, 31, 12) {real, imag} */,
  {32'hbf816acc, 32'hbe9163da} /* (27, 31, 11) {real, imag} */,
  {32'hbdd1c792, 32'h3e10aebb} /* (27, 31, 10) {real, imag} */,
  {32'hbe735c0a, 32'h3f1dab4e} /* (27, 31, 9) {real, imag} */,
  {32'h3d3b9ab8, 32'hbebad6a3} /* (27, 31, 8) {real, imag} */,
  {32'h3e99fb76, 32'hbeb57ac6} /* (27, 31, 7) {real, imag} */,
  {32'hbea5eea1, 32'h3f0ea87b} /* (27, 31, 6) {real, imag} */,
  {32'hc049c86f, 32'hbe74bf50} /* (27, 31, 5) {real, imag} */,
  {32'h3ec18f7f, 32'hbf6d56af} /* (27, 31, 4) {real, imag} */,
  {32'h3e41b018, 32'hbe45ff42} /* (27, 31, 3) {real, imag} */,
  {32'hc0a180c4, 32'hc0062957} /* (27, 31, 2) {real, imag} */,
  {32'h411803d0, 32'h407c004e} /* (27, 31, 1) {real, imag} */,
  {32'h4083ac36, 32'h3e197190} /* (27, 31, 0) {real, imag} */,
  {32'hc10244db, 32'hc06b4504} /* (27, 30, 31) {real, imag} */,
  {32'h410100c2, 32'h40563fb4} /* (27, 30, 30) {real, imag} */,
  {32'h3d8c2e84, 32'h3eefbccf} /* (27, 30, 29) {real, imag} */,
  {32'hc008be87, 32'h3fdc77a4} /* (27, 30, 28) {real, imag} */,
  {32'h3f5c2f2b, 32'hbf94c5a7} /* (27, 30, 27) {real, imag} */,
  {32'hbd24b296, 32'h3e067122} /* (27, 30, 26) {real, imag} */,
  {32'hbe847546, 32'h3ddc2ea0} /* (27, 30, 25) {real, imag} */,
  {32'h3f1939e4, 32'hbf3e9ff9} /* (27, 30, 24) {real, imag} */,
  {32'h3e330e99, 32'hbd179090} /* (27, 30, 23) {real, imag} */,
  {32'hbea6da20, 32'h3f07c0b5} /* (27, 30, 22) {real, imag} */,
  {32'hbea115d8, 32'hbf318e1e} /* (27, 30, 21) {real, imag} */,
  {32'hbee6fa1c, 32'hbe19587e} /* (27, 30, 20) {real, imag} */,
  {32'h3cfffe46, 32'h3ebd37d2} /* (27, 30, 19) {real, imag} */,
  {32'h3e1c1d65, 32'h3d105c88} /* (27, 30, 18) {real, imag} */,
  {32'h3d002f60, 32'hbb4af2e0} /* (27, 30, 17) {real, imag} */,
  {32'hbe88eb1d, 32'h3d0bdd5c} /* (27, 30, 16) {real, imag} */,
  {32'h3f00a813, 32'hbe7d52f0} /* (27, 30, 15) {real, imag} */,
  {32'h3ea31dcf, 32'h3e90e1da} /* (27, 30, 14) {real, imag} */,
  {32'hbdb78b54, 32'h3d9c10a8} /* (27, 30, 13) {real, imag} */,
  {32'h3e9c30e8, 32'hbe49bfb0} /* (27, 30, 12) {real, imag} */,
  {32'h3d6adc14, 32'h3e581515} /* (27, 30, 11) {real, imag} */,
  {32'hbe801b4f, 32'h3eb7e102} /* (27, 30, 10) {real, imag} */,
  {32'h3eecfb96, 32'hbdb3add3} /* (27, 30, 9) {real, imag} */,
  {32'h3ee2d8ce, 32'h3f1d7c5a} /* (27, 30, 8) {real, imag} */,
  {32'hbd5e9688, 32'hbf818f7b} /* (27, 30, 7) {real, imag} */,
  {32'h3e84fa0c, 32'h3e6894fb} /* (27, 30, 6) {real, imag} */,
  {32'h3f8615a2, 32'h3fadbd5b} /* (27, 30, 5) {real, imag} */,
  {32'hbf1e34d9, 32'hc0275e12} /* (27, 30, 4) {real, imag} */,
  {32'hbf3458b2, 32'hbd1d2510} /* (27, 30, 3) {real, imag} */,
  {32'h411da3ec, 32'h40659e92} /* (27, 30, 2) {real, imag} */,
  {32'hc15b2dce, 32'hbfbd744f} /* (27, 30, 1) {real, imag} */,
  {32'hc0ce7eff, 32'h4059d8f0} /* (27, 30, 0) {real, imag} */,
  {32'h3fdc4ef9, 32'hc06695fb} /* (27, 29, 31) {real, imag} */,
  {32'hbd4388a0, 32'h4025c636} /* (27, 29, 30) {real, imag} */,
  {32'hbde9513e, 32'hbe87f9b4} /* (27, 29, 29) {real, imag} */,
  {32'hbd435610, 32'hbf763c0a} /* (27, 29, 28) {real, imag} */,
  {32'h3ea33c8c, 32'hbdb2b51a} /* (27, 29, 27) {real, imag} */,
  {32'hbf6cf93a, 32'h3e2967a6} /* (27, 29, 26) {real, imag} */,
  {32'h3e2bba19, 32'hbeccc0e3} /* (27, 29, 25) {real, imag} */,
  {32'hbeb5d000, 32'hbb6ec340} /* (27, 29, 24) {real, imag} */,
  {32'h3ec9c73a, 32'hbf1171e1} /* (27, 29, 23) {real, imag} */,
  {32'hbec95b6c, 32'h3e988ab9} /* (27, 29, 22) {real, imag} */,
  {32'h3ed26b56, 32'h3de91f9e} /* (27, 29, 21) {real, imag} */,
  {32'h3d2ebc9c, 32'h3f58b63c} /* (27, 29, 20) {real, imag} */,
  {32'h3d9c88a8, 32'hbd97533e} /* (27, 29, 19) {real, imag} */,
  {32'hbe14ea3a, 32'hbe0d50fe} /* (27, 29, 18) {real, imag} */,
  {32'h3d93461c, 32'hbde3caee} /* (27, 29, 17) {real, imag} */,
  {32'h3e2d2138, 32'h3e9748c6} /* (27, 29, 16) {real, imag} */,
  {32'hbe8ebf6e, 32'h3ec66ba6} /* (27, 29, 15) {real, imag} */,
  {32'h3d24de4a, 32'h3cdcf09c} /* (27, 29, 14) {real, imag} */,
  {32'hbd490cee, 32'hbe7ecc16} /* (27, 29, 13) {real, imag} */,
  {32'hbe2d0f9e, 32'h3f400362} /* (27, 29, 12) {real, imag} */,
  {32'hbd895674, 32'hbeac2759} /* (27, 29, 11) {real, imag} */,
  {32'h3f1c31b4, 32'hbed30580} /* (27, 29, 10) {real, imag} */,
  {32'h3ecb6aba, 32'hbeb03d49} /* (27, 29, 9) {real, imag} */,
  {32'hbf5d36f2, 32'h3ef60dec} /* (27, 29, 8) {real, imag} */,
  {32'h3ef0100a, 32'hbe221a1b} /* (27, 29, 7) {real, imag} */,
  {32'h3eafb106, 32'hbf350600} /* (27, 29, 6) {real, imag} */,
  {32'hbf11d7a0, 32'h3f210e02} /* (27, 29, 5) {real, imag} */,
  {32'h3f3e1560, 32'hbf003889} /* (27, 29, 4) {real, imag} */,
  {32'hbede59b8, 32'hbdb0fc20} /* (27, 29, 3) {real, imag} */,
  {32'h401e489b, 32'h400c9735} /* (27, 29, 2) {real, imag} */,
  {32'hc053fafa, 32'hbf3d7322} /* (27, 29, 1) {real, imag} */,
  {32'h3fde5ea8, 32'hbe9ca644} /* (27, 29, 0) {real, imag} */,
  {32'h403881f6, 32'hc02adb38} /* (27, 28, 31) {real, imag} */,
  {32'hbfca82ad, 32'h4014c728} /* (27, 28, 30) {real, imag} */,
  {32'h3f32c8af, 32'h3e242fba} /* (27, 28, 29) {real, imag} */,
  {32'h3fd8aefe, 32'h3e524ab0} /* (27, 28, 28) {real, imag} */,
  {32'hbda0e50c, 32'h3f4530cf} /* (27, 28, 27) {real, imag} */,
  {32'hbec9695b, 32'hbcb10b48} /* (27, 28, 26) {real, imag} */,
  {32'h3e6f767e, 32'hbeb01302} /* (27, 28, 25) {real, imag} */,
  {32'hbeb351e2, 32'hbe7245e2} /* (27, 28, 24) {real, imag} */,
  {32'h3da63342, 32'h3e9a8b7e} /* (27, 28, 23) {real, imag} */,
  {32'hbe430bf0, 32'hbe80a57e} /* (27, 28, 22) {real, imag} */,
  {32'hbf2dde9c, 32'hbea5efe1} /* (27, 28, 21) {real, imag} */,
  {32'hbd52a578, 32'h3eae5a12} /* (27, 28, 20) {real, imag} */,
  {32'h3e3e8789, 32'hbeb24175} /* (27, 28, 19) {real, imag} */,
  {32'hbec4270c, 32'hbe4e4517} /* (27, 28, 18) {real, imag} */,
  {32'hbe0d67d3, 32'hbe1d99a1} /* (27, 28, 17) {real, imag} */,
  {32'h3d5f4456, 32'h3e00512e} /* (27, 28, 16) {real, imag} */,
  {32'h3e0cd94e, 32'h3d9bc627} /* (27, 28, 15) {real, imag} */,
  {32'hbbd947c0, 32'h3e67ec8a} /* (27, 28, 14) {real, imag} */,
  {32'hbdc56931, 32'hbebcbc25} /* (27, 28, 13) {real, imag} */,
  {32'h3e00a630, 32'h3d48b968} /* (27, 28, 12) {real, imag} */,
  {32'hbf01b231, 32'hbe8bb5a0} /* (27, 28, 11) {real, imag} */,
  {32'h3f6e405b, 32'h3e8c89a5} /* (27, 28, 10) {real, imag} */,
  {32'hbdec8c0b, 32'hbe93aad8} /* (27, 28, 9) {real, imag} */,
  {32'h3e4db023, 32'h3d985976} /* (27, 28, 8) {real, imag} */,
  {32'hbef703d0, 32'h3eb294b3} /* (27, 28, 7) {real, imag} */,
  {32'hbd0aef70, 32'hbf5a1ab0} /* (27, 28, 6) {real, imag} */,
  {32'h3eba01b6, 32'h3e51a504} /* (27, 28, 5) {real, imag} */,
  {32'h3d4e1194, 32'h3e72622f} /* (27, 28, 4) {real, imag} */,
  {32'h3dde9a15, 32'h3f031010} /* (27, 28, 3) {real, imag} */,
  {32'hbfd5cf0f, 32'h3fded96c} /* (27, 28, 2) {real, imag} */,
  {32'h3f2732f9, 32'hbf9a1c8a} /* (27, 28, 1) {real, imag} */,
  {32'h3de97564, 32'hbe61ba87} /* (27, 28, 0) {real, imag} */,
  {32'hbfda1798, 32'h3f8e8ee7} /* (27, 27, 31) {real, imag} */,
  {32'h3f1fb4a0, 32'h3eaefa44} /* (27, 27, 30) {real, imag} */,
  {32'hbccc2f50, 32'h3f47fc55} /* (27, 27, 29) {real, imag} */,
  {32'h3ec4d278, 32'hbe62403d} /* (27, 27, 28) {real, imag} */,
  {32'h3f4d1ee8, 32'hbe8f1eb2} /* (27, 27, 27) {real, imag} */,
  {32'h3eb8836a, 32'hbe84c585} /* (27, 27, 26) {real, imag} */,
  {32'hbee55151, 32'h3d506f30} /* (27, 27, 25) {real, imag} */,
  {32'hbd7e3914, 32'hbdf2bafd} /* (27, 27, 24) {real, imag} */,
  {32'h3dcaa73a, 32'h3ebfe0e8} /* (27, 27, 23) {real, imag} */,
  {32'h3ed97fe0, 32'hbd8e5348} /* (27, 27, 22) {real, imag} */,
  {32'hbec16ad7, 32'h3e981a95} /* (27, 27, 21) {real, imag} */,
  {32'hbde847af, 32'h3f0ca2c5} /* (27, 27, 20) {real, imag} */,
  {32'h3dbdeddc, 32'hbdfd825c} /* (27, 27, 19) {real, imag} */,
  {32'hbe628b64, 32'hbe3a13d0} /* (27, 27, 18) {real, imag} */,
  {32'hbe7d9e44, 32'hbe8e523d} /* (27, 27, 17) {real, imag} */,
  {32'h3d726c78, 32'h3cf65758} /* (27, 27, 16) {real, imag} */,
  {32'hbe18dda3, 32'hbdb67f37} /* (27, 27, 15) {real, imag} */,
  {32'h3e72a8cc, 32'h3ef98082} /* (27, 27, 14) {real, imag} */,
  {32'hbf255147, 32'hbe087ca9} /* (27, 27, 13) {real, imag} */,
  {32'h3eb4bb18, 32'h3f156e16} /* (27, 27, 12) {real, imag} */,
  {32'hbdb9d608, 32'h3e16789c} /* (27, 27, 11) {real, imag} */,
  {32'hbda7b7aa, 32'h3e90f9b8} /* (27, 27, 10) {real, imag} */,
  {32'hbc662460, 32'hbf13db7a} /* (27, 27, 9) {real, imag} */,
  {32'hbe32a3d4, 32'hbf2a7853} /* (27, 27, 8) {real, imag} */,
  {32'h3e4886c4, 32'hbdbfbf6a} /* (27, 27, 7) {real, imag} */,
  {32'hbd67b4c8, 32'h3d40e1a8} /* (27, 27, 6) {real, imag} */,
  {32'h3f49df62, 32'h3f14b7b2} /* (27, 27, 5) {real, imag} */,
  {32'hbec237e1, 32'hbf824c48} /* (27, 27, 4) {real, imag} */,
  {32'h3e267210, 32'h3e530ea5} /* (27, 27, 3) {real, imag} */,
  {32'h3f9b5eb8, 32'h3f0bbabe} /* (27, 27, 2) {real, imag} */,
  {32'hc01fef84, 32'h3f8af04b} /* (27, 27, 1) {real, imag} */,
  {32'hc00feb59, 32'h3ec8c32b} /* (27, 27, 0) {real, imag} */,
  {32'hbdadfe14, 32'h3f257130} /* (27, 26, 31) {real, imag} */,
  {32'h3f50a624, 32'h3e523582} /* (27, 26, 30) {real, imag} */,
  {32'hbd3c99b0, 32'h3ebbc695} /* (27, 26, 29) {real, imag} */,
  {32'hbe370dd0, 32'hb9d81700} /* (27, 26, 28) {real, imag} */,
  {32'h3e2d7e68, 32'hbc96f7c8} /* (27, 26, 27) {real, imag} */,
  {32'h3c0d50f0, 32'hbe2f6564} /* (27, 26, 26) {real, imag} */,
  {32'h3ea00e0c, 32'h3e1209d7} /* (27, 26, 25) {real, imag} */,
  {32'hbf4fe459, 32'hbe7ff674} /* (27, 26, 24) {real, imag} */,
  {32'hbcc66a14, 32'h3da6e71a} /* (27, 26, 23) {real, imag} */,
  {32'hbf16a01e, 32'hbe4b4284} /* (27, 26, 22) {real, imag} */,
  {32'hbe1a86a8, 32'hbe4f2ee0} /* (27, 26, 21) {real, imag} */,
  {32'hbdc4c442, 32'h3ea5c871} /* (27, 26, 20) {real, imag} */,
  {32'h3e3d97ee, 32'hbe08c70e} /* (27, 26, 19) {real, imag} */,
  {32'hbe7e628b, 32'h3eaa3c5b} /* (27, 26, 18) {real, imag} */,
  {32'hbe16725e, 32'h3f034f5e} /* (27, 26, 17) {real, imag} */,
  {32'hbe001044, 32'hbea69c66} /* (27, 26, 16) {real, imag} */,
  {32'h3c1a4610, 32'hbe2894ec} /* (27, 26, 15) {real, imag} */,
  {32'h3eaac7ee, 32'h3c42f100} /* (27, 26, 14) {real, imag} */,
  {32'hbe055830, 32'h3eb23663} /* (27, 26, 13) {real, imag} */,
  {32'hbe864031, 32'h3ec0714a} /* (27, 26, 12) {real, imag} */,
  {32'h3e63a359, 32'hbecee442} /* (27, 26, 11) {real, imag} */,
  {32'h3e7ed69b, 32'h3bb6ce20} /* (27, 26, 10) {real, imag} */,
  {32'hbd88924e, 32'h3e29088c} /* (27, 26, 9) {real, imag} */,
  {32'hbe9ed2bc, 32'h3e4e50cd} /* (27, 26, 8) {real, imag} */,
  {32'hbe46cf9a, 32'hbe48b9d2} /* (27, 26, 7) {real, imag} */,
  {32'h3ec2f739, 32'h3f2e63fe} /* (27, 26, 6) {real, imag} */,
  {32'h3f0388ae, 32'h3c56be50} /* (27, 26, 5) {real, imag} */,
  {32'h3dea3b5c, 32'hbde3e24e} /* (27, 26, 4) {real, imag} */,
  {32'h3ef9c22e, 32'h3e88c7c0} /* (27, 26, 3) {real, imag} */,
  {32'hbe187bb3, 32'hbd9b9a10} /* (27, 26, 2) {real, imag} */,
  {32'hbf1d2f18, 32'h3d821646} /* (27, 26, 1) {real, imag} */,
  {32'h3e35af1c, 32'h3f3e8495} /* (27, 26, 0) {real, imag} */,
  {32'h3f4de80b, 32'hbebe775e} /* (27, 25, 31) {real, imag} */,
  {32'hbe80fd82, 32'hbeb5baad} /* (27, 25, 30) {real, imag} */,
  {32'h3f084e1e, 32'h3d80a54a} /* (27, 25, 29) {real, imag} */,
  {32'h3ec92ff8, 32'h3d4d6d6e} /* (27, 25, 28) {real, imag} */,
  {32'hbe0a9d38, 32'h3e5f83dc} /* (27, 25, 27) {real, imag} */,
  {32'h3eead942, 32'hbe07d093} /* (27, 25, 26) {real, imag} */,
  {32'h3dc2be7e, 32'hbca9c564} /* (27, 25, 25) {real, imag} */,
  {32'hbe748170, 32'h3ea56cbc} /* (27, 25, 24) {real, imag} */,
  {32'h3eeedafe, 32'hbe398fa0} /* (27, 25, 23) {real, imag} */,
  {32'h3e083331, 32'hbee7915d} /* (27, 25, 22) {real, imag} */,
  {32'hbf04fb42, 32'h3ecb0d4d} /* (27, 25, 21) {real, imag} */,
  {32'h3e21d508, 32'hbdc33947} /* (27, 25, 20) {real, imag} */,
  {32'hbdbf72a4, 32'h3e7728e0} /* (27, 25, 19) {real, imag} */,
  {32'h3e9a993a, 32'hbd9ab95e} /* (27, 25, 18) {real, imag} */,
  {32'h3e2effb7, 32'h3e60b5f2} /* (27, 25, 17) {real, imag} */,
  {32'h3f0b3f1e, 32'hbe80ab4d} /* (27, 25, 16) {real, imag} */,
  {32'hbea712ad, 32'h3e8b232f} /* (27, 25, 15) {real, imag} */,
  {32'hbe6ea909, 32'h3e1c1046} /* (27, 25, 14) {real, imag} */,
  {32'h3ec5b795, 32'hbe72fd00} /* (27, 25, 13) {real, imag} */,
  {32'hbea29f3d, 32'h3d793b08} /* (27, 25, 12) {real, imag} */,
  {32'h3f6a6e13, 32'hbe375baa} /* (27, 25, 11) {real, imag} */,
  {32'h3f337304, 32'h3ea6109f} /* (27, 25, 10) {real, imag} */,
  {32'h3d916ea4, 32'hbef87966} /* (27, 25, 9) {real, imag} */,
  {32'hbe459762, 32'hbe8510f9} /* (27, 25, 8) {real, imag} */,
  {32'h3c0f2600, 32'hbf252522} /* (27, 25, 7) {real, imag} */,
  {32'h3e999720, 32'hbd86b660} /* (27, 25, 6) {real, imag} */,
  {32'hbef1542f, 32'h3cb4f114} /* (27, 25, 5) {real, imag} */,
  {32'hbf009cec, 32'h3f14cf23} /* (27, 25, 4) {real, imag} */,
  {32'h3e254207, 32'hbd6918a5} /* (27, 25, 3) {real, imag} */,
  {32'hbde63b04, 32'h3f27f2e8} /* (27, 25, 2) {real, imag} */,
  {32'hbe16fd6c, 32'hbf26946b} /* (27, 25, 1) {real, imag} */,
  {32'h3f210288, 32'h3ed520ba} /* (27, 25, 0) {real, imag} */,
  {32'hbf4e83cc, 32'h3eedeb44} /* (27, 24, 31) {real, imag} */,
  {32'h3e501873, 32'hbd779b60} /* (27, 24, 30) {real, imag} */,
  {32'h3c915460, 32'hbea5c898} /* (27, 24, 29) {real, imag} */,
  {32'hbf3d9314, 32'h3e0971d7} /* (27, 24, 28) {real, imag} */,
  {32'h3e96684c, 32'hbf1fa76a} /* (27, 24, 27) {real, imag} */,
  {32'hbee254e2, 32'h3e75d222} /* (27, 24, 26) {real, imag} */,
  {32'h3f54cc58, 32'hbeccb8aa} /* (27, 24, 25) {real, imag} */,
  {32'hbe8ab63c, 32'hbd7df6e0} /* (27, 24, 24) {real, imag} */,
  {32'hbe62b0da, 32'hbbade280} /* (27, 24, 23) {real, imag} */,
  {32'hbda67ba8, 32'h3f2d71d9} /* (27, 24, 22) {real, imag} */,
  {32'h3f0929a5, 32'hbec24e7e} /* (27, 24, 21) {real, imag} */,
  {32'h3e3e398a, 32'h3e4178c4} /* (27, 24, 20) {real, imag} */,
  {32'h3daced20, 32'h3c313930} /* (27, 24, 19) {real, imag} */,
  {32'hbe95a0a0, 32'hbf0d1dce} /* (27, 24, 18) {real, imag} */,
  {32'hbecde61a, 32'h3d9654ba} /* (27, 24, 17) {real, imag} */,
  {32'hbcd5a6a0, 32'hbd60e4e4} /* (27, 24, 16) {real, imag} */,
  {32'h3e85f180, 32'hbea2f7e2} /* (27, 24, 15) {real, imag} */,
  {32'hbe727e90, 32'hbdfdec6f} /* (27, 24, 14) {real, imag} */,
  {32'hbd57a99f, 32'hbe24f782} /* (27, 24, 13) {real, imag} */,
  {32'h3f1d05d8, 32'h3eb25e51} /* (27, 24, 12) {real, imag} */,
  {32'h3ec81968, 32'hbe529627} /* (27, 24, 11) {real, imag} */,
  {32'hbf076675, 32'h3dcccf44} /* (27, 24, 10) {real, imag} */,
  {32'hbeb90367, 32'h3ebe830e} /* (27, 24, 9) {real, imag} */,
  {32'h3e23bfb7, 32'hbec072d8} /* (27, 24, 8) {real, imag} */,
  {32'hbd92005e, 32'h3ec512d8} /* (27, 24, 7) {real, imag} */,
  {32'hbe48d23e, 32'h3c19a310} /* (27, 24, 6) {real, imag} */,
  {32'hbf2be020, 32'h3ec8f104} /* (27, 24, 5) {real, imag} */,
  {32'h3e8f8e1e, 32'h3eb70c9c} /* (27, 24, 4) {real, imag} */,
  {32'h3ddce6f8, 32'h3f0dd46b} /* (27, 24, 3) {real, imag} */,
  {32'h3f0709a5, 32'hbc04b248} /* (27, 24, 2) {real, imag} */,
  {32'hbfb2bee8, 32'h3f0b7f20} /* (27, 24, 1) {real, imag} */,
  {32'hbf1d2840, 32'h3e881326} /* (27, 24, 0) {real, imag} */,
  {32'h3e8d731a, 32'h3f4bc9ec} /* (27, 23, 31) {real, imag} */,
  {32'h3edfb0f0, 32'h3edd2c93} /* (27, 23, 30) {real, imag} */,
  {32'hbe971a36, 32'h3f04ea97} /* (27, 23, 29) {real, imag} */,
  {32'h3cd2f5f2, 32'hbed8fce9} /* (27, 23, 28) {real, imag} */,
  {32'h3ebe9468, 32'hbf47569e} /* (27, 23, 27) {real, imag} */,
  {32'hbecd7231, 32'hbf01192a} /* (27, 23, 26) {real, imag} */,
  {32'hbc6800d0, 32'hbedbdae4} /* (27, 23, 25) {real, imag} */,
  {32'h3ebd17e1, 32'hbc026b10} /* (27, 23, 24) {real, imag} */,
  {32'h3e820308, 32'h3ebab4fb} /* (27, 23, 23) {real, imag} */,
  {32'hbe878ed7, 32'h3e9bf1e8} /* (27, 23, 22) {real, imag} */,
  {32'h3e7d792e, 32'hbe9b2fc2} /* (27, 23, 21) {real, imag} */,
  {32'h3aadc9c0, 32'hbe4d9232} /* (27, 23, 20) {real, imag} */,
  {32'h3da80d1c, 32'h3e86218f} /* (27, 23, 19) {real, imag} */,
  {32'h3f076bce, 32'hbd00aef6} /* (27, 23, 18) {real, imag} */,
  {32'hbd736f0c, 32'h3e0941e4} /* (27, 23, 17) {real, imag} */,
  {32'hbe0b0f88, 32'hbec40f96} /* (27, 23, 16) {real, imag} */,
  {32'h3e198766, 32'hbd4df3f8} /* (27, 23, 15) {real, imag} */,
  {32'hbd9b5548, 32'h3e25ba98} /* (27, 23, 14) {real, imag} */,
  {32'h3e2bc49f, 32'h3ee530a8} /* (27, 23, 13) {real, imag} */,
  {32'h3eb0fde5, 32'h3e8ebb2e} /* (27, 23, 12) {real, imag} */,
  {32'h3e9f7095, 32'hbeb837c8} /* (27, 23, 11) {real, imag} */,
  {32'hbe2cc7e7, 32'h3efae98a} /* (27, 23, 10) {real, imag} */,
  {32'hbe1ffffe, 32'h3ed94c78} /* (27, 23, 9) {real, imag} */,
  {32'hbebb681f, 32'h3ef6dccd} /* (27, 23, 8) {real, imag} */,
  {32'h3e9669b3, 32'hbe752374} /* (27, 23, 7) {real, imag} */,
  {32'hbf067d48, 32'hbebadc64} /* (27, 23, 6) {real, imag} */,
  {32'hbe4c44fb, 32'hbcf5c978} /* (27, 23, 5) {real, imag} */,
  {32'hbeeaa86f, 32'hbe5a38d2} /* (27, 23, 4) {real, imag} */,
  {32'hbd491df2, 32'h3e01f6a6} /* (27, 23, 3) {real, imag} */,
  {32'h3f27efe4, 32'h3e6709a8} /* (27, 23, 2) {real, imag} */,
  {32'hbf42a1a4, 32'hbf0c3b53} /* (27, 23, 1) {real, imag} */,
  {32'hbe4d061c, 32'hbecb7d4a} /* (27, 23, 0) {real, imag} */,
  {32'h3f1c6399, 32'h3b972d50} /* (27, 22, 31) {real, imag} */,
  {32'hbf45f5bc, 32'h3dd51794} /* (27, 22, 30) {real, imag} */,
  {32'hbe5db25c, 32'hbe5d5135} /* (27, 22, 29) {real, imag} */,
  {32'h3edd2c9e, 32'hbf1bff3e} /* (27, 22, 28) {real, imag} */,
  {32'h3de6c88f, 32'h3cc33bca} /* (27, 22, 27) {real, imag} */,
  {32'hbd89b1bd, 32'h3e54eb28} /* (27, 22, 26) {real, imag} */,
  {32'h3f01cd56, 32'h3f227cf8} /* (27, 22, 25) {real, imag} */,
  {32'h3ed18eed, 32'hbea0a4e4} /* (27, 22, 24) {real, imag} */,
  {32'h3d1e4088, 32'h3ea21fe0} /* (27, 22, 23) {real, imag} */,
  {32'hbde3eb06, 32'h3e474d36} /* (27, 22, 22) {real, imag} */,
  {32'hbe0effdb, 32'hbd0cce0e} /* (27, 22, 21) {real, imag} */,
  {32'hbd892b94, 32'hbda2aac0} /* (27, 22, 20) {real, imag} */,
  {32'hbe4dbe4c, 32'h3e961ae9} /* (27, 22, 19) {real, imag} */,
  {32'h3d2e4342, 32'h3e256d52} /* (27, 22, 18) {real, imag} */,
  {32'hbeab0677, 32'hbe770448} /* (27, 22, 17) {real, imag} */,
  {32'h3ea05302, 32'h3e079754} /* (27, 22, 16) {real, imag} */,
  {32'hbe7dff40, 32'hbeeb16ee} /* (27, 22, 15) {real, imag} */,
  {32'hbe804ccd, 32'hbe03822a} /* (27, 22, 14) {real, imag} */,
  {32'h3d14931c, 32'h3ea37553} /* (27, 22, 13) {real, imag} */,
  {32'hbd47bd32, 32'hbed3485e} /* (27, 22, 12) {real, imag} */,
  {32'hbea6840c, 32'hbe769cf0} /* (27, 22, 11) {real, imag} */,
  {32'hbe898f61, 32'h3f308573} /* (27, 22, 10) {real, imag} */,
  {32'h3e289623, 32'hbf04a87f} /* (27, 22, 9) {real, imag} */,
  {32'h3c8f5db0, 32'h3ea46940} /* (27, 22, 8) {real, imag} */,
  {32'hbeefb57a, 32'h3e808186} /* (27, 22, 7) {real, imag} */,
  {32'h3ea888bc, 32'h3ea2990f} /* (27, 22, 6) {real, imag} */,
  {32'hbe97dcc3, 32'h3ea68340} /* (27, 22, 5) {real, imag} */,
  {32'hbe5aede9, 32'h3e1f6cfd} /* (27, 22, 4) {real, imag} */,
  {32'h3e0d0f72, 32'hbed940e9} /* (27, 22, 3) {real, imag} */,
  {32'h3e4a4acb, 32'h3ea4678a} /* (27, 22, 2) {real, imag} */,
  {32'hbf09b75c, 32'hbee880b5} /* (27, 22, 1) {real, imag} */,
  {32'h3e0778b5, 32'hbd87ef2a} /* (27, 22, 0) {real, imag} */,
  {32'hbe29e3a4, 32'h3f1fc7aa} /* (27, 21, 31) {real, imag} */,
  {32'hbe1755b1, 32'hbec47bc0} /* (27, 21, 30) {real, imag} */,
  {32'h3ea1b13e, 32'hbe536579} /* (27, 21, 29) {real, imag} */,
  {32'hbd28ca58, 32'h3ea445a9} /* (27, 21, 28) {real, imag} */,
  {32'hbf257f29, 32'hbec8af01} /* (27, 21, 27) {real, imag} */,
  {32'hbf00d48d, 32'hbe3c325e} /* (27, 21, 26) {real, imag} */,
  {32'h3e2d90ee, 32'h3dca204a} /* (27, 21, 25) {real, imag} */,
  {32'h3db8c6ce, 32'hbc4ad680} /* (27, 21, 24) {real, imag} */,
  {32'h3ea24d76, 32'hbe12147a} /* (27, 21, 23) {real, imag} */,
  {32'h3d0fd1d0, 32'h3e8aad94} /* (27, 21, 22) {real, imag} */,
  {32'h3e5bdbf4, 32'hbdd903d5} /* (27, 21, 21) {real, imag} */,
  {32'h3e867e8a, 32'hbe0a8792} /* (27, 21, 20) {real, imag} */,
  {32'hbf252468, 32'hbe92b7a6} /* (27, 21, 19) {real, imag} */,
  {32'h3e34ed21, 32'h3e95d0de} /* (27, 21, 18) {real, imag} */,
  {32'hbb835540, 32'hbe2204b0} /* (27, 21, 17) {real, imag} */,
  {32'hbeab08aa, 32'hbed5fdfc} /* (27, 21, 16) {real, imag} */,
  {32'hbe8537b9, 32'h3ed1906f} /* (27, 21, 15) {real, imag} */,
  {32'h3e2e2d20, 32'h3eaab526} /* (27, 21, 14) {real, imag} */,
  {32'h3e826210, 32'hbe024daa} /* (27, 21, 13) {real, imag} */,
  {32'h3e98261c, 32'hbec9e26c} /* (27, 21, 12) {real, imag} */,
  {32'h3e8c05bd, 32'hbe84c589} /* (27, 21, 11) {real, imag} */,
  {32'h3bf4cab0, 32'hbeeb50cc} /* (27, 21, 10) {real, imag} */,
  {32'h3d6ea392, 32'h3e848896} /* (27, 21, 9) {real, imag} */,
  {32'hbdbfb646, 32'h3b23ccd0} /* (27, 21, 8) {real, imag} */,
  {32'h3e341e2e, 32'h3eec93ba} /* (27, 21, 7) {real, imag} */,
  {32'hbde59877, 32'h3d7206f2} /* (27, 21, 6) {real, imag} */,
  {32'hbd302ef3, 32'hbedee18c} /* (27, 21, 5) {real, imag} */,
  {32'h3c884b40, 32'hbecfc47e} /* (27, 21, 4) {real, imag} */,
  {32'h3ee8edf2, 32'h3e939a3f} /* (27, 21, 3) {real, imag} */,
  {32'h3d3e9d90, 32'h3e3b317e} /* (27, 21, 2) {real, imag} */,
  {32'hbe7de776, 32'h3eb517f0} /* (27, 21, 1) {real, imag} */,
  {32'hbe417977, 32'h3eb12387} /* (27, 21, 0) {real, imag} */,
  {32'hbd91d5f4, 32'hbe8be7ae} /* (27, 20, 31) {real, imag} */,
  {32'hbebc4246, 32'h3e0ed098} /* (27, 20, 30) {real, imag} */,
  {32'h3eada972, 32'hbe6dff76} /* (27, 20, 29) {real, imag} */,
  {32'hbf1ac1e2, 32'hbd6d672c} /* (27, 20, 28) {real, imag} */,
  {32'h3f36285e, 32'h3ec5493f} /* (27, 20, 27) {real, imag} */,
  {32'hbcb1ab08, 32'h3e971c61} /* (27, 20, 26) {real, imag} */,
  {32'hbddf7f08, 32'hbcc03350} /* (27, 20, 25) {real, imag} */,
  {32'hbdfc5e08, 32'h3e30e956} /* (27, 20, 24) {real, imag} */,
  {32'h3e640f44, 32'h3e813058} /* (27, 20, 23) {real, imag} */,
  {32'h3ee8baa3, 32'hbe880b69} /* (27, 20, 22) {real, imag} */,
  {32'h3e9a296c, 32'h3e8abab5} /* (27, 20, 21) {real, imag} */,
  {32'hbe01e657, 32'h3ec89d02} /* (27, 20, 20) {real, imag} */,
  {32'h3d78e6f4, 32'h3dda2499} /* (27, 20, 19) {real, imag} */,
  {32'hbf465766, 32'h3dc90880} /* (27, 20, 18) {real, imag} */,
  {32'hbc177a20, 32'hbe061c9c} /* (27, 20, 17) {real, imag} */,
  {32'h3b9d0ff8, 32'hbde08d0d} /* (27, 20, 16) {real, imag} */,
  {32'h3e0cd60b, 32'hbe95634f} /* (27, 20, 15) {real, imag} */,
  {32'hbe874e0c, 32'h3c76e430} /* (27, 20, 14) {real, imag} */,
  {32'h3d4d6dce, 32'h3e4c42d7} /* (27, 20, 13) {real, imag} */,
  {32'hbdcda95c, 32'hbf0bae9b} /* (27, 20, 12) {real, imag} */,
  {32'h3ebcba34, 32'h3eb12f9c} /* (27, 20, 11) {real, imag} */,
  {32'h3f172d4c, 32'h3e7fa70e} /* (27, 20, 10) {real, imag} */,
  {32'h3efa1ee6, 32'h3f08e680} /* (27, 20, 9) {real, imag} */,
  {32'hbe6269ae, 32'hbf160bc8} /* (27, 20, 8) {real, imag} */,
  {32'h3e7fba5c, 32'h3e556326} /* (27, 20, 7) {real, imag} */,
  {32'hbe90f92a, 32'h3f08bec2} /* (27, 20, 6) {real, imag} */,
  {32'hbddda597, 32'hbf118175} /* (27, 20, 5) {real, imag} */,
  {32'hbf0bb2f2, 32'h3e97753b} /* (27, 20, 4) {real, imag} */,
  {32'hbe5670c4, 32'h3c8a6b70} /* (27, 20, 3) {real, imag} */,
  {32'hbe9cd02b, 32'h3efe1bc4} /* (27, 20, 2) {real, imag} */,
  {32'hbbd57330, 32'h3d4036ba} /* (27, 20, 1) {real, imag} */,
  {32'h3e9361ef, 32'h3e42fb8f} /* (27, 20, 0) {real, imag} */,
  {32'h3e864276, 32'hbdb2e441} /* (27, 19, 31) {real, imag} */,
  {32'hbdabdde8, 32'hbe306b6e} /* (27, 19, 30) {real, imag} */,
  {32'hbdb56b96, 32'h3d68faf1} /* (27, 19, 29) {real, imag} */,
  {32'hbd98aab2, 32'h3e1d2958} /* (27, 19, 28) {real, imag} */,
  {32'h3e7ddfa5, 32'hbe47a856} /* (27, 19, 27) {real, imag} */,
  {32'hbf013305, 32'h3dfda0e0} /* (27, 19, 26) {real, imag} */,
  {32'h3df73c98, 32'hbd910c4e} /* (27, 19, 25) {real, imag} */,
  {32'h3d38f49d, 32'hbf40be6e} /* (27, 19, 24) {real, imag} */,
  {32'h3e40cd73, 32'hbd23b7f0} /* (27, 19, 23) {real, imag} */,
  {32'h3e9b9e66, 32'h3dfe4d13} /* (27, 19, 22) {real, imag} */,
  {32'hbe25734f, 32'hbe69659a} /* (27, 19, 21) {real, imag} */,
  {32'h3e999484, 32'hbd3d785c} /* (27, 19, 20) {real, imag} */,
  {32'h3e8a1e5c, 32'h3f08737e} /* (27, 19, 19) {real, imag} */,
  {32'h3e5cb82a, 32'h3db719e2} /* (27, 19, 18) {real, imag} */,
  {32'h3e843b58, 32'h3e38e938} /* (27, 19, 17) {real, imag} */,
  {32'h3d9cc122, 32'h3e5bd0b1} /* (27, 19, 16) {real, imag} */,
  {32'h3c8774c0, 32'hbc5c8a10} /* (27, 19, 15) {real, imag} */,
  {32'hbed83360, 32'h3e69be91} /* (27, 19, 14) {real, imag} */,
  {32'hbe51e522, 32'h3da2e74b} /* (27, 19, 13) {real, imag} */,
  {32'hbd722630, 32'h3e05faa2} /* (27, 19, 12) {real, imag} */,
  {32'hbdab8e10, 32'hbe7acb24} /* (27, 19, 11) {real, imag} */,
  {32'h3e97cafb, 32'hbed797ca} /* (27, 19, 10) {real, imag} */,
  {32'h3eff2d3a, 32'hbf1924c0} /* (27, 19, 9) {real, imag} */,
  {32'h3d13b004, 32'hbe058018} /* (27, 19, 8) {real, imag} */,
  {32'hbe23d391, 32'h3e4d9c03} /* (27, 19, 7) {real, imag} */,
  {32'hbe93c571, 32'hbd5a251a} /* (27, 19, 6) {real, imag} */,
  {32'h3c4ef4f8, 32'hbe0fd09d} /* (27, 19, 5) {real, imag} */,
  {32'h3db0d64e, 32'h3ea2c536} /* (27, 19, 4) {real, imag} */,
  {32'hbea1d018, 32'hbcff2b80} /* (27, 19, 3) {real, imag} */,
  {32'hbdce7bc8, 32'h3e1a3993} /* (27, 19, 2) {real, imag} */,
  {32'hbe8af6b6, 32'h3c902060} /* (27, 19, 1) {real, imag} */,
  {32'hbe5ee5a4, 32'h3dd58886} /* (27, 19, 0) {real, imag} */,
  {32'hbe8ee311, 32'h3ef68990} /* (27, 18, 31) {real, imag} */,
  {32'hbd8a0a90, 32'hbf0b5d9a} /* (27, 18, 30) {real, imag} */,
  {32'h3f13c229, 32'h3dc324a4} /* (27, 18, 29) {real, imag} */,
  {32'hbeca559e, 32'h3ee228e5} /* (27, 18, 28) {real, imag} */,
  {32'hbe4f82e6, 32'h3e29b716} /* (27, 18, 27) {real, imag} */,
  {32'hbc81252c, 32'hbb2fa3c0} /* (27, 18, 26) {real, imag} */,
  {32'hbdf1704c, 32'hbdae672c} /* (27, 18, 25) {real, imag} */,
  {32'hbd8126e0, 32'hbf2ebdf9} /* (27, 18, 24) {real, imag} */,
  {32'hbe10af1d, 32'hbb0d4530} /* (27, 18, 23) {real, imag} */,
  {32'hbe42350a, 32'hbe89fc9f} /* (27, 18, 22) {real, imag} */,
  {32'h3caacc80, 32'h3e624622} /* (27, 18, 21) {real, imag} */,
  {32'hbdea5e24, 32'hbf336762} /* (27, 18, 20) {real, imag} */,
  {32'hbe091777, 32'h3e52db22} /* (27, 18, 19) {real, imag} */,
  {32'h3e825519, 32'hbe941e88} /* (27, 18, 18) {real, imag} */,
  {32'h3e552249, 32'h3ea0b8dd} /* (27, 18, 17) {real, imag} */,
  {32'hbccf8fa4, 32'hbdff9f6c} /* (27, 18, 16) {real, imag} */,
  {32'h3db2c3fd, 32'hbe5c9c16} /* (27, 18, 15) {real, imag} */,
  {32'h3e61d3d8, 32'h3d73a24f} /* (27, 18, 14) {real, imag} */,
  {32'h3e0e9f8d, 32'h3b0812e0} /* (27, 18, 13) {real, imag} */,
  {32'h3e2e15e0, 32'h3f11e91b} /* (27, 18, 12) {real, imag} */,
  {32'h3d55ffbc, 32'h3e040742} /* (27, 18, 11) {real, imag} */,
  {32'hbf21104c, 32'h3f240f65} /* (27, 18, 10) {real, imag} */,
  {32'hbe51663f, 32'h3e94efb4} /* (27, 18, 9) {real, imag} */,
  {32'h3e912acf, 32'hbd49619e} /* (27, 18, 8) {real, imag} */,
  {32'h3e8305a2, 32'h3e648712} /* (27, 18, 7) {real, imag} */,
  {32'hbede7f45, 32'hbd9800a4} /* (27, 18, 6) {real, imag} */,
  {32'h3a89d720, 32'h3e5ed89d} /* (27, 18, 5) {real, imag} */,
  {32'hbe6da60c, 32'h3d35b7a8} /* (27, 18, 4) {real, imag} */,
  {32'h3e127422, 32'h3da77b3b} /* (27, 18, 3) {real, imag} */,
  {32'hbe308450, 32'hbe743798} /* (27, 18, 2) {real, imag} */,
  {32'hbf128b0b, 32'h3e9e58c6} /* (27, 18, 1) {real, imag} */,
  {32'hbbef9ae0, 32'h3eb83e98} /* (27, 18, 0) {real, imag} */,
  {32'h3e34d318, 32'h3d650fac} /* (27, 17, 31) {real, imag} */,
  {32'h3e09e59f, 32'h3ec456e7} /* (27, 17, 30) {real, imag} */,
  {32'hbe0c0707, 32'h3e1cc1ac} /* (27, 17, 29) {real, imag} */,
  {32'hbda53772, 32'h3e965f16} /* (27, 17, 28) {real, imag} */,
  {32'h3dc72588, 32'hbe3042c8} /* (27, 17, 27) {real, imag} */,
  {32'h3e19e31a, 32'h3da1f763} /* (27, 17, 26) {real, imag} */,
  {32'h3dd1f98e, 32'hbdae7634} /* (27, 17, 25) {real, imag} */,
  {32'hbddf820a, 32'hbd9f9ab3} /* (27, 17, 24) {real, imag} */,
  {32'hbe8c098a, 32'hbe5eccc6} /* (27, 17, 23) {real, imag} */,
  {32'h3e2d94cb, 32'hbdbf4b96} /* (27, 17, 22) {real, imag} */,
  {32'h3ed1b982, 32'hbdd03464} /* (27, 17, 21) {real, imag} */,
  {32'hb982cc00, 32'h3e644f8e} /* (27, 17, 20) {real, imag} */,
  {32'hbdd93cf6, 32'hbe006df2} /* (27, 17, 19) {real, imag} */,
  {32'hbdf04285, 32'h3f300cb4} /* (27, 17, 18) {real, imag} */,
  {32'h3d016a12, 32'h3ec9ed56} /* (27, 17, 17) {real, imag} */,
  {32'hbe2dd904, 32'h3db9c482} /* (27, 17, 16) {real, imag} */,
  {32'hbd8aff41, 32'hbec0f3d8} /* (27, 17, 15) {real, imag} */,
  {32'h3db60d2e, 32'h3ea61f7c} /* (27, 17, 14) {real, imag} */,
  {32'h3e477900, 32'hbe154ebd} /* (27, 17, 13) {real, imag} */,
  {32'hbec88ac1, 32'hbec5a090} /* (27, 17, 12) {real, imag} */,
  {32'h3cd81940, 32'h3eca2758} /* (27, 17, 11) {real, imag} */,
  {32'hbcd7ddce, 32'hbf43271c} /* (27, 17, 10) {real, imag} */,
  {32'h3e311d6d, 32'hbbfe9d00} /* (27, 17, 9) {real, imag} */,
  {32'hbc4cc010, 32'hbe01902a} /* (27, 17, 8) {real, imag} */,
  {32'h3e8a0aa6, 32'hbd864ec0} /* (27, 17, 7) {real, imag} */,
  {32'h3e669813, 32'h3d53dd20} /* (27, 17, 6) {real, imag} */,
  {32'hbec5fb9a, 32'h3e9e791a} /* (27, 17, 5) {real, imag} */,
  {32'h3eb6a53a, 32'hbde1b1aa} /* (27, 17, 4) {real, imag} */,
  {32'h3e103185, 32'h3ea26822} /* (27, 17, 3) {real, imag} */,
  {32'hbed9ad6a, 32'h3ea6d0ba} /* (27, 17, 2) {real, imag} */,
  {32'hbea4414e, 32'hbd9a3934} /* (27, 17, 1) {real, imag} */,
  {32'hbe2842ad, 32'hbe8c4bf7} /* (27, 17, 0) {real, imag} */,
  {32'h3cae38e4, 32'h3e9dddea} /* (27, 16, 31) {real, imag} */,
  {32'hbe17342c, 32'h3e6d45ba} /* (27, 16, 30) {real, imag} */,
  {32'h3d3bdc92, 32'h3ddc73c0} /* (27, 16, 29) {real, imag} */,
  {32'h3e199264, 32'hbe1d4dec} /* (27, 16, 28) {real, imag} */,
  {32'hbe1c746c, 32'h3e8b8a02} /* (27, 16, 27) {real, imag} */,
  {32'h3d8f6aa2, 32'h3e375278} /* (27, 16, 26) {real, imag} */,
  {32'h3a03eb40, 32'hbea97fe4} /* (27, 16, 25) {real, imag} */,
  {32'hbd21b6d4, 32'h3e80af56} /* (27, 16, 24) {real, imag} */,
  {32'hbdb59594, 32'h3d288632} /* (27, 16, 23) {real, imag} */,
  {32'h3c8e2ba0, 32'hbcda3ebe} /* (27, 16, 22) {real, imag} */,
  {32'h3e94c1e3, 32'h3d732876} /* (27, 16, 21) {real, imag} */,
  {32'h3de65a8d, 32'hbebfb4ae} /* (27, 16, 20) {real, imag} */,
  {32'hbec0241b, 32'hbf14932e} /* (27, 16, 19) {real, imag} */,
  {32'h3d9f567c, 32'h3eb30c22} /* (27, 16, 18) {real, imag} */,
  {32'hbe3bacbb, 32'h3e44b335} /* (27, 16, 17) {real, imag} */,
  {32'hbccf940c, 32'h00000000} /* (27, 16, 16) {real, imag} */,
  {32'hbe3bacbb, 32'hbe44b335} /* (27, 16, 15) {real, imag} */,
  {32'h3d9f567c, 32'hbeb30c22} /* (27, 16, 14) {real, imag} */,
  {32'hbec0241b, 32'h3f14932e} /* (27, 16, 13) {real, imag} */,
  {32'h3de65a8d, 32'h3ebfb4ae} /* (27, 16, 12) {real, imag} */,
  {32'h3e94c1e3, 32'hbd732876} /* (27, 16, 11) {real, imag} */,
  {32'h3c8e2ba0, 32'h3cda3ebe} /* (27, 16, 10) {real, imag} */,
  {32'hbdb59594, 32'hbd288632} /* (27, 16, 9) {real, imag} */,
  {32'hbd21b6d4, 32'hbe80af56} /* (27, 16, 8) {real, imag} */,
  {32'h3a03eb40, 32'h3ea97fe4} /* (27, 16, 7) {real, imag} */,
  {32'h3d8f6aa2, 32'hbe375278} /* (27, 16, 6) {real, imag} */,
  {32'hbe1c746c, 32'hbe8b8a02} /* (27, 16, 5) {real, imag} */,
  {32'h3e199264, 32'h3e1d4dec} /* (27, 16, 4) {real, imag} */,
  {32'h3d3bdc92, 32'hbddc73c0} /* (27, 16, 3) {real, imag} */,
  {32'hbe17342c, 32'hbe6d45ba} /* (27, 16, 2) {real, imag} */,
  {32'h3cae38e4, 32'hbe9dddea} /* (27, 16, 1) {real, imag} */,
  {32'hbee5da4f, 32'h00000000} /* (27, 16, 0) {real, imag} */,
  {32'hbea4414e, 32'h3d9a3934} /* (27, 15, 31) {real, imag} */,
  {32'hbed9ad6a, 32'hbea6d0ba} /* (27, 15, 30) {real, imag} */,
  {32'h3e103185, 32'hbea26822} /* (27, 15, 29) {real, imag} */,
  {32'h3eb6a53a, 32'h3de1b1aa} /* (27, 15, 28) {real, imag} */,
  {32'hbec5fb9a, 32'hbe9e791a} /* (27, 15, 27) {real, imag} */,
  {32'h3e669813, 32'hbd53dd20} /* (27, 15, 26) {real, imag} */,
  {32'h3e8a0aa6, 32'h3d864ec0} /* (27, 15, 25) {real, imag} */,
  {32'hbc4cc010, 32'h3e01902a} /* (27, 15, 24) {real, imag} */,
  {32'h3e311d6d, 32'h3bfe9d00} /* (27, 15, 23) {real, imag} */,
  {32'hbcd7ddce, 32'h3f43271c} /* (27, 15, 22) {real, imag} */,
  {32'h3cd81940, 32'hbeca2758} /* (27, 15, 21) {real, imag} */,
  {32'hbec88ac1, 32'h3ec5a090} /* (27, 15, 20) {real, imag} */,
  {32'h3e477900, 32'h3e154ebd} /* (27, 15, 19) {real, imag} */,
  {32'h3db60d2e, 32'hbea61f7c} /* (27, 15, 18) {real, imag} */,
  {32'hbd8aff41, 32'h3ec0f3d8} /* (27, 15, 17) {real, imag} */,
  {32'hbe2dd904, 32'hbdb9c482} /* (27, 15, 16) {real, imag} */,
  {32'h3d016a12, 32'hbec9ed56} /* (27, 15, 15) {real, imag} */,
  {32'hbdf04285, 32'hbf300cb4} /* (27, 15, 14) {real, imag} */,
  {32'hbdd93cf6, 32'h3e006df2} /* (27, 15, 13) {real, imag} */,
  {32'hb982cc00, 32'hbe644f8e} /* (27, 15, 12) {real, imag} */,
  {32'h3ed1b982, 32'h3dd03464} /* (27, 15, 11) {real, imag} */,
  {32'h3e2d94cb, 32'h3dbf4b96} /* (27, 15, 10) {real, imag} */,
  {32'hbe8c098a, 32'h3e5eccc6} /* (27, 15, 9) {real, imag} */,
  {32'hbddf820a, 32'h3d9f9ab3} /* (27, 15, 8) {real, imag} */,
  {32'h3dd1f98e, 32'h3dae7634} /* (27, 15, 7) {real, imag} */,
  {32'h3e19e31a, 32'hbda1f763} /* (27, 15, 6) {real, imag} */,
  {32'h3dc72588, 32'h3e3042c8} /* (27, 15, 5) {real, imag} */,
  {32'hbda53772, 32'hbe965f16} /* (27, 15, 4) {real, imag} */,
  {32'hbe0c0707, 32'hbe1cc1ac} /* (27, 15, 3) {real, imag} */,
  {32'h3e09e59f, 32'hbec456e7} /* (27, 15, 2) {real, imag} */,
  {32'h3e34d318, 32'hbd650fac} /* (27, 15, 1) {real, imag} */,
  {32'hbe2842ad, 32'h3e8c4bf7} /* (27, 15, 0) {real, imag} */,
  {32'hbf128b0b, 32'hbe9e58c6} /* (27, 14, 31) {real, imag} */,
  {32'hbe308450, 32'h3e743798} /* (27, 14, 30) {real, imag} */,
  {32'h3e127422, 32'hbda77b3b} /* (27, 14, 29) {real, imag} */,
  {32'hbe6da60c, 32'hbd35b7a8} /* (27, 14, 28) {real, imag} */,
  {32'h3a89d720, 32'hbe5ed89d} /* (27, 14, 27) {real, imag} */,
  {32'hbede7f45, 32'h3d9800a4} /* (27, 14, 26) {real, imag} */,
  {32'h3e8305a2, 32'hbe648712} /* (27, 14, 25) {real, imag} */,
  {32'h3e912acf, 32'h3d49619e} /* (27, 14, 24) {real, imag} */,
  {32'hbe51663f, 32'hbe94efb4} /* (27, 14, 23) {real, imag} */,
  {32'hbf21104c, 32'hbf240f65} /* (27, 14, 22) {real, imag} */,
  {32'h3d55ffbc, 32'hbe040742} /* (27, 14, 21) {real, imag} */,
  {32'h3e2e15e0, 32'hbf11e91b} /* (27, 14, 20) {real, imag} */,
  {32'h3e0e9f8d, 32'hbb0812e0} /* (27, 14, 19) {real, imag} */,
  {32'h3e61d3d8, 32'hbd73a24f} /* (27, 14, 18) {real, imag} */,
  {32'h3db2c3fd, 32'h3e5c9c16} /* (27, 14, 17) {real, imag} */,
  {32'hbccf8fa4, 32'h3dff9f6c} /* (27, 14, 16) {real, imag} */,
  {32'h3e552249, 32'hbea0b8dd} /* (27, 14, 15) {real, imag} */,
  {32'h3e825519, 32'h3e941e88} /* (27, 14, 14) {real, imag} */,
  {32'hbe091777, 32'hbe52db22} /* (27, 14, 13) {real, imag} */,
  {32'hbdea5e24, 32'h3f336762} /* (27, 14, 12) {real, imag} */,
  {32'h3caacc80, 32'hbe624622} /* (27, 14, 11) {real, imag} */,
  {32'hbe42350a, 32'h3e89fc9f} /* (27, 14, 10) {real, imag} */,
  {32'hbe10af1d, 32'h3b0d4530} /* (27, 14, 9) {real, imag} */,
  {32'hbd8126e0, 32'h3f2ebdf9} /* (27, 14, 8) {real, imag} */,
  {32'hbdf1704c, 32'h3dae672c} /* (27, 14, 7) {real, imag} */,
  {32'hbc81252c, 32'h3b2fa3c0} /* (27, 14, 6) {real, imag} */,
  {32'hbe4f82e6, 32'hbe29b716} /* (27, 14, 5) {real, imag} */,
  {32'hbeca559e, 32'hbee228e5} /* (27, 14, 4) {real, imag} */,
  {32'h3f13c229, 32'hbdc324a4} /* (27, 14, 3) {real, imag} */,
  {32'hbd8a0a90, 32'h3f0b5d9a} /* (27, 14, 2) {real, imag} */,
  {32'hbe8ee311, 32'hbef68990} /* (27, 14, 1) {real, imag} */,
  {32'hbbef9ae0, 32'hbeb83e98} /* (27, 14, 0) {real, imag} */,
  {32'hbe8af6b6, 32'hbc902060} /* (27, 13, 31) {real, imag} */,
  {32'hbdce7bc8, 32'hbe1a3993} /* (27, 13, 30) {real, imag} */,
  {32'hbea1d018, 32'h3cff2b80} /* (27, 13, 29) {real, imag} */,
  {32'h3db0d64e, 32'hbea2c536} /* (27, 13, 28) {real, imag} */,
  {32'h3c4ef4f8, 32'h3e0fd09d} /* (27, 13, 27) {real, imag} */,
  {32'hbe93c571, 32'h3d5a251a} /* (27, 13, 26) {real, imag} */,
  {32'hbe23d391, 32'hbe4d9c03} /* (27, 13, 25) {real, imag} */,
  {32'h3d13b004, 32'h3e058018} /* (27, 13, 24) {real, imag} */,
  {32'h3eff2d3a, 32'h3f1924c0} /* (27, 13, 23) {real, imag} */,
  {32'h3e97cafb, 32'h3ed797ca} /* (27, 13, 22) {real, imag} */,
  {32'hbdab8e10, 32'h3e7acb24} /* (27, 13, 21) {real, imag} */,
  {32'hbd722630, 32'hbe05faa2} /* (27, 13, 20) {real, imag} */,
  {32'hbe51e522, 32'hbda2e74b} /* (27, 13, 19) {real, imag} */,
  {32'hbed83360, 32'hbe69be91} /* (27, 13, 18) {real, imag} */,
  {32'h3c8774c0, 32'h3c5c8a10} /* (27, 13, 17) {real, imag} */,
  {32'h3d9cc122, 32'hbe5bd0b1} /* (27, 13, 16) {real, imag} */,
  {32'h3e843b58, 32'hbe38e938} /* (27, 13, 15) {real, imag} */,
  {32'h3e5cb82a, 32'hbdb719e2} /* (27, 13, 14) {real, imag} */,
  {32'h3e8a1e5c, 32'hbf08737e} /* (27, 13, 13) {real, imag} */,
  {32'h3e999484, 32'h3d3d785c} /* (27, 13, 12) {real, imag} */,
  {32'hbe25734f, 32'h3e69659a} /* (27, 13, 11) {real, imag} */,
  {32'h3e9b9e66, 32'hbdfe4d13} /* (27, 13, 10) {real, imag} */,
  {32'h3e40cd73, 32'h3d23b7f0} /* (27, 13, 9) {real, imag} */,
  {32'h3d38f49d, 32'h3f40be6e} /* (27, 13, 8) {real, imag} */,
  {32'h3df73c98, 32'h3d910c4e} /* (27, 13, 7) {real, imag} */,
  {32'hbf013305, 32'hbdfda0e0} /* (27, 13, 6) {real, imag} */,
  {32'h3e7ddfa5, 32'h3e47a856} /* (27, 13, 5) {real, imag} */,
  {32'hbd98aab2, 32'hbe1d2958} /* (27, 13, 4) {real, imag} */,
  {32'hbdb56b96, 32'hbd68faf1} /* (27, 13, 3) {real, imag} */,
  {32'hbdabdde8, 32'h3e306b6e} /* (27, 13, 2) {real, imag} */,
  {32'h3e864276, 32'h3db2e441} /* (27, 13, 1) {real, imag} */,
  {32'hbe5ee5a4, 32'hbdd58886} /* (27, 13, 0) {real, imag} */,
  {32'hbbd57330, 32'hbd4036ba} /* (27, 12, 31) {real, imag} */,
  {32'hbe9cd02b, 32'hbefe1bc4} /* (27, 12, 30) {real, imag} */,
  {32'hbe5670c4, 32'hbc8a6b70} /* (27, 12, 29) {real, imag} */,
  {32'hbf0bb2f2, 32'hbe97753b} /* (27, 12, 28) {real, imag} */,
  {32'hbddda597, 32'h3f118175} /* (27, 12, 27) {real, imag} */,
  {32'hbe90f92a, 32'hbf08bec2} /* (27, 12, 26) {real, imag} */,
  {32'h3e7fba5c, 32'hbe556326} /* (27, 12, 25) {real, imag} */,
  {32'hbe6269ae, 32'h3f160bc8} /* (27, 12, 24) {real, imag} */,
  {32'h3efa1ee6, 32'hbf08e680} /* (27, 12, 23) {real, imag} */,
  {32'h3f172d4c, 32'hbe7fa70e} /* (27, 12, 22) {real, imag} */,
  {32'h3ebcba34, 32'hbeb12f9c} /* (27, 12, 21) {real, imag} */,
  {32'hbdcda95c, 32'h3f0bae9b} /* (27, 12, 20) {real, imag} */,
  {32'h3d4d6dce, 32'hbe4c42d7} /* (27, 12, 19) {real, imag} */,
  {32'hbe874e0c, 32'hbc76e430} /* (27, 12, 18) {real, imag} */,
  {32'h3e0cd60b, 32'h3e95634f} /* (27, 12, 17) {real, imag} */,
  {32'h3b9d0ff8, 32'h3de08d0d} /* (27, 12, 16) {real, imag} */,
  {32'hbc177a20, 32'h3e061c9c} /* (27, 12, 15) {real, imag} */,
  {32'hbf465766, 32'hbdc90880} /* (27, 12, 14) {real, imag} */,
  {32'h3d78e6f4, 32'hbdda2499} /* (27, 12, 13) {real, imag} */,
  {32'hbe01e657, 32'hbec89d02} /* (27, 12, 12) {real, imag} */,
  {32'h3e9a296c, 32'hbe8abab5} /* (27, 12, 11) {real, imag} */,
  {32'h3ee8baa3, 32'h3e880b69} /* (27, 12, 10) {real, imag} */,
  {32'h3e640f44, 32'hbe813058} /* (27, 12, 9) {real, imag} */,
  {32'hbdfc5e08, 32'hbe30e956} /* (27, 12, 8) {real, imag} */,
  {32'hbddf7f08, 32'h3cc03350} /* (27, 12, 7) {real, imag} */,
  {32'hbcb1ab08, 32'hbe971c61} /* (27, 12, 6) {real, imag} */,
  {32'h3f36285e, 32'hbec5493f} /* (27, 12, 5) {real, imag} */,
  {32'hbf1ac1e2, 32'h3d6d672c} /* (27, 12, 4) {real, imag} */,
  {32'h3eada972, 32'h3e6dff76} /* (27, 12, 3) {real, imag} */,
  {32'hbebc4246, 32'hbe0ed098} /* (27, 12, 2) {real, imag} */,
  {32'hbd91d5f4, 32'h3e8be7ae} /* (27, 12, 1) {real, imag} */,
  {32'h3e9361ef, 32'hbe42fb8f} /* (27, 12, 0) {real, imag} */,
  {32'hbe7de776, 32'hbeb517f0} /* (27, 11, 31) {real, imag} */,
  {32'h3d3e9d90, 32'hbe3b317e} /* (27, 11, 30) {real, imag} */,
  {32'h3ee8edf2, 32'hbe939a3f} /* (27, 11, 29) {real, imag} */,
  {32'h3c884b40, 32'h3ecfc47e} /* (27, 11, 28) {real, imag} */,
  {32'hbd302ef3, 32'h3edee18c} /* (27, 11, 27) {real, imag} */,
  {32'hbde59877, 32'hbd7206f2} /* (27, 11, 26) {real, imag} */,
  {32'h3e341e2e, 32'hbeec93ba} /* (27, 11, 25) {real, imag} */,
  {32'hbdbfb646, 32'hbb23ccd0} /* (27, 11, 24) {real, imag} */,
  {32'h3d6ea392, 32'hbe848896} /* (27, 11, 23) {real, imag} */,
  {32'h3bf4cab0, 32'h3eeb50cc} /* (27, 11, 22) {real, imag} */,
  {32'h3e8c05bd, 32'h3e84c589} /* (27, 11, 21) {real, imag} */,
  {32'h3e98261c, 32'h3ec9e26c} /* (27, 11, 20) {real, imag} */,
  {32'h3e826210, 32'h3e024daa} /* (27, 11, 19) {real, imag} */,
  {32'h3e2e2d20, 32'hbeaab526} /* (27, 11, 18) {real, imag} */,
  {32'hbe8537b9, 32'hbed1906f} /* (27, 11, 17) {real, imag} */,
  {32'hbeab08aa, 32'h3ed5fdfc} /* (27, 11, 16) {real, imag} */,
  {32'hbb835540, 32'h3e2204b0} /* (27, 11, 15) {real, imag} */,
  {32'h3e34ed21, 32'hbe95d0de} /* (27, 11, 14) {real, imag} */,
  {32'hbf252468, 32'h3e92b7a6} /* (27, 11, 13) {real, imag} */,
  {32'h3e867e8a, 32'h3e0a8792} /* (27, 11, 12) {real, imag} */,
  {32'h3e5bdbf4, 32'h3dd903d5} /* (27, 11, 11) {real, imag} */,
  {32'h3d0fd1d0, 32'hbe8aad94} /* (27, 11, 10) {real, imag} */,
  {32'h3ea24d76, 32'h3e12147a} /* (27, 11, 9) {real, imag} */,
  {32'h3db8c6ce, 32'h3c4ad680} /* (27, 11, 8) {real, imag} */,
  {32'h3e2d90ee, 32'hbdca204a} /* (27, 11, 7) {real, imag} */,
  {32'hbf00d48d, 32'h3e3c325e} /* (27, 11, 6) {real, imag} */,
  {32'hbf257f29, 32'h3ec8af01} /* (27, 11, 5) {real, imag} */,
  {32'hbd28ca58, 32'hbea445a9} /* (27, 11, 4) {real, imag} */,
  {32'h3ea1b13e, 32'h3e536579} /* (27, 11, 3) {real, imag} */,
  {32'hbe1755b1, 32'h3ec47bc0} /* (27, 11, 2) {real, imag} */,
  {32'hbe29e3a4, 32'hbf1fc7aa} /* (27, 11, 1) {real, imag} */,
  {32'hbe417977, 32'hbeb12387} /* (27, 11, 0) {real, imag} */,
  {32'hbf09b75c, 32'h3ee880b5} /* (27, 10, 31) {real, imag} */,
  {32'h3e4a4acb, 32'hbea4678a} /* (27, 10, 30) {real, imag} */,
  {32'h3e0d0f72, 32'h3ed940e9} /* (27, 10, 29) {real, imag} */,
  {32'hbe5aede9, 32'hbe1f6cfd} /* (27, 10, 28) {real, imag} */,
  {32'hbe97dcc3, 32'hbea68340} /* (27, 10, 27) {real, imag} */,
  {32'h3ea888bc, 32'hbea2990f} /* (27, 10, 26) {real, imag} */,
  {32'hbeefb57a, 32'hbe808186} /* (27, 10, 25) {real, imag} */,
  {32'h3c8f5db0, 32'hbea46940} /* (27, 10, 24) {real, imag} */,
  {32'h3e289623, 32'h3f04a87f} /* (27, 10, 23) {real, imag} */,
  {32'hbe898f61, 32'hbf308573} /* (27, 10, 22) {real, imag} */,
  {32'hbea6840c, 32'h3e769cf0} /* (27, 10, 21) {real, imag} */,
  {32'hbd47bd32, 32'h3ed3485e} /* (27, 10, 20) {real, imag} */,
  {32'h3d14931c, 32'hbea37553} /* (27, 10, 19) {real, imag} */,
  {32'hbe804ccd, 32'h3e03822a} /* (27, 10, 18) {real, imag} */,
  {32'hbe7dff40, 32'h3eeb16ee} /* (27, 10, 17) {real, imag} */,
  {32'h3ea05302, 32'hbe079754} /* (27, 10, 16) {real, imag} */,
  {32'hbeab0677, 32'h3e770448} /* (27, 10, 15) {real, imag} */,
  {32'h3d2e4342, 32'hbe256d52} /* (27, 10, 14) {real, imag} */,
  {32'hbe4dbe4c, 32'hbe961ae9} /* (27, 10, 13) {real, imag} */,
  {32'hbd892b94, 32'h3da2aac0} /* (27, 10, 12) {real, imag} */,
  {32'hbe0effdb, 32'h3d0cce0e} /* (27, 10, 11) {real, imag} */,
  {32'hbde3eb06, 32'hbe474d36} /* (27, 10, 10) {real, imag} */,
  {32'h3d1e4088, 32'hbea21fe0} /* (27, 10, 9) {real, imag} */,
  {32'h3ed18eed, 32'h3ea0a4e4} /* (27, 10, 8) {real, imag} */,
  {32'h3f01cd56, 32'hbf227cf8} /* (27, 10, 7) {real, imag} */,
  {32'hbd89b1bd, 32'hbe54eb28} /* (27, 10, 6) {real, imag} */,
  {32'h3de6c88f, 32'hbcc33bca} /* (27, 10, 5) {real, imag} */,
  {32'h3edd2c9e, 32'h3f1bff3e} /* (27, 10, 4) {real, imag} */,
  {32'hbe5db25c, 32'h3e5d5135} /* (27, 10, 3) {real, imag} */,
  {32'hbf45f5bc, 32'hbdd51794} /* (27, 10, 2) {real, imag} */,
  {32'h3f1c6399, 32'hbb972d50} /* (27, 10, 1) {real, imag} */,
  {32'h3e0778b5, 32'h3d87ef2a} /* (27, 10, 0) {real, imag} */,
  {32'hbf42a1a4, 32'h3f0c3b53} /* (27, 9, 31) {real, imag} */,
  {32'h3f27efe4, 32'hbe6709a8} /* (27, 9, 30) {real, imag} */,
  {32'hbd491df2, 32'hbe01f6a6} /* (27, 9, 29) {real, imag} */,
  {32'hbeeaa86f, 32'h3e5a38d2} /* (27, 9, 28) {real, imag} */,
  {32'hbe4c44fb, 32'h3cf5c978} /* (27, 9, 27) {real, imag} */,
  {32'hbf067d48, 32'h3ebadc64} /* (27, 9, 26) {real, imag} */,
  {32'h3e9669b3, 32'h3e752374} /* (27, 9, 25) {real, imag} */,
  {32'hbebb681f, 32'hbef6dccd} /* (27, 9, 24) {real, imag} */,
  {32'hbe1ffffe, 32'hbed94c78} /* (27, 9, 23) {real, imag} */,
  {32'hbe2cc7e7, 32'hbefae98a} /* (27, 9, 22) {real, imag} */,
  {32'h3e9f7095, 32'h3eb837c8} /* (27, 9, 21) {real, imag} */,
  {32'h3eb0fde5, 32'hbe8ebb2e} /* (27, 9, 20) {real, imag} */,
  {32'h3e2bc49f, 32'hbee530a8} /* (27, 9, 19) {real, imag} */,
  {32'hbd9b5548, 32'hbe25ba98} /* (27, 9, 18) {real, imag} */,
  {32'h3e198766, 32'h3d4df3f8} /* (27, 9, 17) {real, imag} */,
  {32'hbe0b0f88, 32'h3ec40f96} /* (27, 9, 16) {real, imag} */,
  {32'hbd736f0c, 32'hbe0941e4} /* (27, 9, 15) {real, imag} */,
  {32'h3f076bce, 32'h3d00aef6} /* (27, 9, 14) {real, imag} */,
  {32'h3da80d1c, 32'hbe86218f} /* (27, 9, 13) {real, imag} */,
  {32'h3aadc9c0, 32'h3e4d9232} /* (27, 9, 12) {real, imag} */,
  {32'h3e7d792e, 32'h3e9b2fc2} /* (27, 9, 11) {real, imag} */,
  {32'hbe878ed7, 32'hbe9bf1e8} /* (27, 9, 10) {real, imag} */,
  {32'h3e820308, 32'hbebab4fb} /* (27, 9, 9) {real, imag} */,
  {32'h3ebd17e1, 32'h3c026b10} /* (27, 9, 8) {real, imag} */,
  {32'hbc6800d0, 32'h3edbdae4} /* (27, 9, 7) {real, imag} */,
  {32'hbecd7231, 32'h3f01192a} /* (27, 9, 6) {real, imag} */,
  {32'h3ebe9468, 32'h3f47569e} /* (27, 9, 5) {real, imag} */,
  {32'h3cd2f5f2, 32'h3ed8fce9} /* (27, 9, 4) {real, imag} */,
  {32'hbe971a36, 32'hbf04ea97} /* (27, 9, 3) {real, imag} */,
  {32'h3edfb0f0, 32'hbedd2c93} /* (27, 9, 2) {real, imag} */,
  {32'h3e8d731a, 32'hbf4bc9ec} /* (27, 9, 1) {real, imag} */,
  {32'hbe4d061c, 32'h3ecb7d4a} /* (27, 9, 0) {real, imag} */,
  {32'hbfb2bee8, 32'hbf0b7f20} /* (27, 8, 31) {real, imag} */,
  {32'h3f0709a5, 32'h3c04b248} /* (27, 8, 30) {real, imag} */,
  {32'h3ddce6f8, 32'hbf0dd46b} /* (27, 8, 29) {real, imag} */,
  {32'h3e8f8e1e, 32'hbeb70c9c} /* (27, 8, 28) {real, imag} */,
  {32'hbf2be020, 32'hbec8f104} /* (27, 8, 27) {real, imag} */,
  {32'hbe48d23e, 32'hbc19a310} /* (27, 8, 26) {real, imag} */,
  {32'hbd92005e, 32'hbec512d8} /* (27, 8, 25) {real, imag} */,
  {32'h3e23bfb7, 32'h3ec072d8} /* (27, 8, 24) {real, imag} */,
  {32'hbeb90367, 32'hbebe830e} /* (27, 8, 23) {real, imag} */,
  {32'hbf076675, 32'hbdcccf44} /* (27, 8, 22) {real, imag} */,
  {32'h3ec81968, 32'h3e529627} /* (27, 8, 21) {real, imag} */,
  {32'h3f1d05d8, 32'hbeb25e51} /* (27, 8, 20) {real, imag} */,
  {32'hbd57a99f, 32'h3e24f782} /* (27, 8, 19) {real, imag} */,
  {32'hbe727e90, 32'h3dfdec6f} /* (27, 8, 18) {real, imag} */,
  {32'h3e85f180, 32'h3ea2f7e2} /* (27, 8, 17) {real, imag} */,
  {32'hbcd5a6a0, 32'h3d60e4e4} /* (27, 8, 16) {real, imag} */,
  {32'hbecde61a, 32'hbd9654ba} /* (27, 8, 15) {real, imag} */,
  {32'hbe95a0a0, 32'h3f0d1dce} /* (27, 8, 14) {real, imag} */,
  {32'h3daced20, 32'hbc313930} /* (27, 8, 13) {real, imag} */,
  {32'h3e3e398a, 32'hbe4178c4} /* (27, 8, 12) {real, imag} */,
  {32'h3f0929a5, 32'h3ec24e7e} /* (27, 8, 11) {real, imag} */,
  {32'hbda67ba8, 32'hbf2d71d9} /* (27, 8, 10) {real, imag} */,
  {32'hbe62b0da, 32'h3bade280} /* (27, 8, 9) {real, imag} */,
  {32'hbe8ab63c, 32'h3d7df6e0} /* (27, 8, 8) {real, imag} */,
  {32'h3f54cc58, 32'h3eccb8aa} /* (27, 8, 7) {real, imag} */,
  {32'hbee254e2, 32'hbe75d222} /* (27, 8, 6) {real, imag} */,
  {32'h3e96684c, 32'h3f1fa76a} /* (27, 8, 5) {real, imag} */,
  {32'hbf3d9314, 32'hbe0971d7} /* (27, 8, 4) {real, imag} */,
  {32'h3c915460, 32'h3ea5c898} /* (27, 8, 3) {real, imag} */,
  {32'h3e501873, 32'h3d779b60} /* (27, 8, 2) {real, imag} */,
  {32'hbf4e83cc, 32'hbeedeb44} /* (27, 8, 1) {real, imag} */,
  {32'hbf1d2840, 32'hbe881326} /* (27, 8, 0) {real, imag} */,
  {32'hbe16fd6c, 32'h3f26946b} /* (27, 7, 31) {real, imag} */,
  {32'hbde63b04, 32'hbf27f2e8} /* (27, 7, 30) {real, imag} */,
  {32'h3e254207, 32'h3d6918a5} /* (27, 7, 29) {real, imag} */,
  {32'hbf009cec, 32'hbf14cf23} /* (27, 7, 28) {real, imag} */,
  {32'hbef1542f, 32'hbcb4f114} /* (27, 7, 27) {real, imag} */,
  {32'h3e999720, 32'h3d86b660} /* (27, 7, 26) {real, imag} */,
  {32'h3c0f2600, 32'h3f252522} /* (27, 7, 25) {real, imag} */,
  {32'hbe459762, 32'h3e8510f9} /* (27, 7, 24) {real, imag} */,
  {32'h3d916ea4, 32'h3ef87966} /* (27, 7, 23) {real, imag} */,
  {32'h3f337304, 32'hbea6109f} /* (27, 7, 22) {real, imag} */,
  {32'h3f6a6e13, 32'h3e375baa} /* (27, 7, 21) {real, imag} */,
  {32'hbea29f3d, 32'hbd793b08} /* (27, 7, 20) {real, imag} */,
  {32'h3ec5b795, 32'h3e72fd00} /* (27, 7, 19) {real, imag} */,
  {32'hbe6ea909, 32'hbe1c1046} /* (27, 7, 18) {real, imag} */,
  {32'hbea712ad, 32'hbe8b232f} /* (27, 7, 17) {real, imag} */,
  {32'h3f0b3f1e, 32'h3e80ab4d} /* (27, 7, 16) {real, imag} */,
  {32'h3e2effb7, 32'hbe60b5f2} /* (27, 7, 15) {real, imag} */,
  {32'h3e9a993a, 32'h3d9ab95e} /* (27, 7, 14) {real, imag} */,
  {32'hbdbf72a4, 32'hbe7728e0} /* (27, 7, 13) {real, imag} */,
  {32'h3e21d508, 32'h3dc33947} /* (27, 7, 12) {real, imag} */,
  {32'hbf04fb42, 32'hbecb0d4d} /* (27, 7, 11) {real, imag} */,
  {32'h3e083331, 32'h3ee7915d} /* (27, 7, 10) {real, imag} */,
  {32'h3eeedafe, 32'h3e398fa0} /* (27, 7, 9) {real, imag} */,
  {32'hbe748170, 32'hbea56cbc} /* (27, 7, 8) {real, imag} */,
  {32'h3dc2be7e, 32'h3ca9c564} /* (27, 7, 7) {real, imag} */,
  {32'h3eead942, 32'h3e07d093} /* (27, 7, 6) {real, imag} */,
  {32'hbe0a9d38, 32'hbe5f83dc} /* (27, 7, 5) {real, imag} */,
  {32'h3ec92ff8, 32'hbd4d6d6e} /* (27, 7, 4) {real, imag} */,
  {32'h3f084e1e, 32'hbd80a54a} /* (27, 7, 3) {real, imag} */,
  {32'hbe80fd82, 32'h3eb5baad} /* (27, 7, 2) {real, imag} */,
  {32'h3f4de80b, 32'h3ebe775e} /* (27, 7, 1) {real, imag} */,
  {32'h3f210288, 32'hbed520ba} /* (27, 7, 0) {real, imag} */,
  {32'hbf1d2f18, 32'hbd821646} /* (27, 6, 31) {real, imag} */,
  {32'hbe187bb3, 32'h3d9b9a10} /* (27, 6, 30) {real, imag} */,
  {32'h3ef9c22e, 32'hbe88c7c0} /* (27, 6, 29) {real, imag} */,
  {32'h3dea3b5c, 32'h3de3e24e} /* (27, 6, 28) {real, imag} */,
  {32'h3f0388ae, 32'hbc56be50} /* (27, 6, 27) {real, imag} */,
  {32'h3ec2f739, 32'hbf2e63fe} /* (27, 6, 26) {real, imag} */,
  {32'hbe46cf9a, 32'h3e48b9d2} /* (27, 6, 25) {real, imag} */,
  {32'hbe9ed2bc, 32'hbe4e50cd} /* (27, 6, 24) {real, imag} */,
  {32'hbd88924e, 32'hbe29088c} /* (27, 6, 23) {real, imag} */,
  {32'h3e7ed69b, 32'hbbb6ce20} /* (27, 6, 22) {real, imag} */,
  {32'h3e63a359, 32'h3ecee442} /* (27, 6, 21) {real, imag} */,
  {32'hbe864031, 32'hbec0714a} /* (27, 6, 20) {real, imag} */,
  {32'hbe055830, 32'hbeb23663} /* (27, 6, 19) {real, imag} */,
  {32'h3eaac7ee, 32'hbc42f100} /* (27, 6, 18) {real, imag} */,
  {32'h3c1a4610, 32'h3e2894ec} /* (27, 6, 17) {real, imag} */,
  {32'hbe001044, 32'h3ea69c66} /* (27, 6, 16) {real, imag} */,
  {32'hbe16725e, 32'hbf034f5e} /* (27, 6, 15) {real, imag} */,
  {32'hbe7e628b, 32'hbeaa3c5b} /* (27, 6, 14) {real, imag} */,
  {32'h3e3d97ee, 32'h3e08c70e} /* (27, 6, 13) {real, imag} */,
  {32'hbdc4c442, 32'hbea5c871} /* (27, 6, 12) {real, imag} */,
  {32'hbe1a86a8, 32'h3e4f2ee0} /* (27, 6, 11) {real, imag} */,
  {32'hbf16a01e, 32'h3e4b4284} /* (27, 6, 10) {real, imag} */,
  {32'hbcc66a14, 32'hbda6e71a} /* (27, 6, 9) {real, imag} */,
  {32'hbf4fe459, 32'h3e7ff674} /* (27, 6, 8) {real, imag} */,
  {32'h3ea00e0c, 32'hbe1209d7} /* (27, 6, 7) {real, imag} */,
  {32'h3c0d50f0, 32'h3e2f6564} /* (27, 6, 6) {real, imag} */,
  {32'h3e2d7e68, 32'h3c96f7c8} /* (27, 6, 5) {real, imag} */,
  {32'hbe370dd0, 32'h39d81700} /* (27, 6, 4) {real, imag} */,
  {32'hbd3c99b0, 32'hbebbc695} /* (27, 6, 3) {real, imag} */,
  {32'h3f50a624, 32'hbe523582} /* (27, 6, 2) {real, imag} */,
  {32'hbdadfe14, 32'hbf257130} /* (27, 6, 1) {real, imag} */,
  {32'h3e35af1c, 32'hbf3e8495} /* (27, 6, 0) {real, imag} */,
  {32'hc01fef84, 32'hbf8af04b} /* (27, 5, 31) {real, imag} */,
  {32'h3f9b5eb8, 32'hbf0bbabe} /* (27, 5, 30) {real, imag} */,
  {32'h3e267210, 32'hbe530ea5} /* (27, 5, 29) {real, imag} */,
  {32'hbec237e1, 32'h3f824c48} /* (27, 5, 28) {real, imag} */,
  {32'h3f49df62, 32'hbf14b7b2} /* (27, 5, 27) {real, imag} */,
  {32'hbd67b4c8, 32'hbd40e1a8} /* (27, 5, 26) {real, imag} */,
  {32'h3e4886c4, 32'h3dbfbf6a} /* (27, 5, 25) {real, imag} */,
  {32'hbe32a3d4, 32'h3f2a7853} /* (27, 5, 24) {real, imag} */,
  {32'hbc662460, 32'h3f13db7a} /* (27, 5, 23) {real, imag} */,
  {32'hbda7b7aa, 32'hbe90f9b8} /* (27, 5, 22) {real, imag} */,
  {32'hbdb9d608, 32'hbe16789c} /* (27, 5, 21) {real, imag} */,
  {32'h3eb4bb18, 32'hbf156e16} /* (27, 5, 20) {real, imag} */,
  {32'hbf255147, 32'h3e087ca9} /* (27, 5, 19) {real, imag} */,
  {32'h3e72a8cc, 32'hbef98082} /* (27, 5, 18) {real, imag} */,
  {32'hbe18dda3, 32'h3db67f37} /* (27, 5, 17) {real, imag} */,
  {32'h3d726c78, 32'hbcf65758} /* (27, 5, 16) {real, imag} */,
  {32'hbe7d9e44, 32'h3e8e523d} /* (27, 5, 15) {real, imag} */,
  {32'hbe628b64, 32'h3e3a13d0} /* (27, 5, 14) {real, imag} */,
  {32'h3dbdeddc, 32'h3dfd825c} /* (27, 5, 13) {real, imag} */,
  {32'hbde847af, 32'hbf0ca2c5} /* (27, 5, 12) {real, imag} */,
  {32'hbec16ad7, 32'hbe981a95} /* (27, 5, 11) {real, imag} */,
  {32'h3ed97fe0, 32'h3d8e5348} /* (27, 5, 10) {real, imag} */,
  {32'h3dcaa73a, 32'hbebfe0e8} /* (27, 5, 9) {real, imag} */,
  {32'hbd7e3914, 32'h3df2bafd} /* (27, 5, 8) {real, imag} */,
  {32'hbee55151, 32'hbd506f30} /* (27, 5, 7) {real, imag} */,
  {32'h3eb8836a, 32'h3e84c585} /* (27, 5, 6) {real, imag} */,
  {32'h3f4d1ee8, 32'h3e8f1eb2} /* (27, 5, 5) {real, imag} */,
  {32'h3ec4d278, 32'h3e62403d} /* (27, 5, 4) {real, imag} */,
  {32'hbccc2f50, 32'hbf47fc55} /* (27, 5, 3) {real, imag} */,
  {32'h3f1fb4a0, 32'hbeaefa44} /* (27, 5, 2) {real, imag} */,
  {32'hbfda1798, 32'hbf8e8ee7} /* (27, 5, 1) {real, imag} */,
  {32'hc00feb59, 32'hbec8c32b} /* (27, 5, 0) {real, imag} */,
  {32'h3f2732f9, 32'h3f9a1c8a} /* (27, 4, 31) {real, imag} */,
  {32'hbfd5cf0f, 32'hbfded96c} /* (27, 4, 30) {real, imag} */,
  {32'h3dde9a15, 32'hbf031010} /* (27, 4, 29) {real, imag} */,
  {32'h3d4e1194, 32'hbe72622f} /* (27, 4, 28) {real, imag} */,
  {32'h3eba01b6, 32'hbe51a504} /* (27, 4, 27) {real, imag} */,
  {32'hbd0aef70, 32'h3f5a1ab0} /* (27, 4, 26) {real, imag} */,
  {32'hbef703d0, 32'hbeb294b3} /* (27, 4, 25) {real, imag} */,
  {32'h3e4db023, 32'hbd985976} /* (27, 4, 24) {real, imag} */,
  {32'hbdec8c0b, 32'h3e93aad8} /* (27, 4, 23) {real, imag} */,
  {32'h3f6e405b, 32'hbe8c89a5} /* (27, 4, 22) {real, imag} */,
  {32'hbf01b231, 32'h3e8bb5a0} /* (27, 4, 21) {real, imag} */,
  {32'h3e00a630, 32'hbd48b968} /* (27, 4, 20) {real, imag} */,
  {32'hbdc56931, 32'h3ebcbc25} /* (27, 4, 19) {real, imag} */,
  {32'hbbd947c0, 32'hbe67ec8a} /* (27, 4, 18) {real, imag} */,
  {32'h3e0cd94e, 32'hbd9bc627} /* (27, 4, 17) {real, imag} */,
  {32'h3d5f4456, 32'hbe00512e} /* (27, 4, 16) {real, imag} */,
  {32'hbe0d67d3, 32'h3e1d99a1} /* (27, 4, 15) {real, imag} */,
  {32'hbec4270c, 32'h3e4e4517} /* (27, 4, 14) {real, imag} */,
  {32'h3e3e8789, 32'h3eb24175} /* (27, 4, 13) {real, imag} */,
  {32'hbd52a578, 32'hbeae5a12} /* (27, 4, 12) {real, imag} */,
  {32'hbf2dde9c, 32'h3ea5efe1} /* (27, 4, 11) {real, imag} */,
  {32'hbe430bf0, 32'h3e80a57e} /* (27, 4, 10) {real, imag} */,
  {32'h3da63342, 32'hbe9a8b7e} /* (27, 4, 9) {real, imag} */,
  {32'hbeb351e2, 32'h3e7245e2} /* (27, 4, 8) {real, imag} */,
  {32'h3e6f767e, 32'h3eb01302} /* (27, 4, 7) {real, imag} */,
  {32'hbec9695b, 32'h3cb10b48} /* (27, 4, 6) {real, imag} */,
  {32'hbda0e50c, 32'hbf4530cf} /* (27, 4, 5) {real, imag} */,
  {32'h3fd8aefe, 32'hbe524ab0} /* (27, 4, 4) {real, imag} */,
  {32'h3f32c8af, 32'hbe242fba} /* (27, 4, 3) {real, imag} */,
  {32'hbfca82ad, 32'hc014c728} /* (27, 4, 2) {real, imag} */,
  {32'h403881f6, 32'h402adb38} /* (27, 4, 1) {real, imag} */,
  {32'h3de97564, 32'h3e61ba87} /* (27, 4, 0) {real, imag} */,
  {32'hc053fafa, 32'h3f3d7322} /* (27, 3, 31) {real, imag} */,
  {32'h401e489b, 32'hc00c9735} /* (27, 3, 30) {real, imag} */,
  {32'hbede59b8, 32'h3db0fc20} /* (27, 3, 29) {real, imag} */,
  {32'h3f3e1560, 32'h3f003889} /* (27, 3, 28) {real, imag} */,
  {32'hbf11d7a0, 32'hbf210e02} /* (27, 3, 27) {real, imag} */,
  {32'h3eafb106, 32'h3f350600} /* (27, 3, 26) {real, imag} */,
  {32'h3ef0100a, 32'h3e221a1b} /* (27, 3, 25) {real, imag} */,
  {32'hbf5d36f2, 32'hbef60dec} /* (27, 3, 24) {real, imag} */,
  {32'h3ecb6aba, 32'h3eb03d49} /* (27, 3, 23) {real, imag} */,
  {32'h3f1c31b4, 32'h3ed30580} /* (27, 3, 22) {real, imag} */,
  {32'hbd895674, 32'h3eac2759} /* (27, 3, 21) {real, imag} */,
  {32'hbe2d0f9e, 32'hbf400362} /* (27, 3, 20) {real, imag} */,
  {32'hbd490cee, 32'h3e7ecc16} /* (27, 3, 19) {real, imag} */,
  {32'h3d24de4a, 32'hbcdcf09c} /* (27, 3, 18) {real, imag} */,
  {32'hbe8ebf6e, 32'hbec66ba6} /* (27, 3, 17) {real, imag} */,
  {32'h3e2d2138, 32'hbe9748c6} /* (27, 3, 16) {real, imag} */,
  {32'h3d93461c, 32'h3de3caee} /* (27, 3, 15) {real, imag} */,
  {32'hbe14ea3a, 32'h3e0d50fe} /* (27, 3, 14) {real, imag} */,
  {32'h3d9c88a8, 32'h3d97533e} /* (27, 3, 13) {real, imag} */,
  {32'h3d2ebc9c, 32'hbf58b63c} /* (27, 3, 12) {real, imag} */,
  {32'h3ed26b56, 32'hbde91f9e} /* (27, 3, 11) {real, imag} */,
  {32'hbec95b6c, 32'hbe988ab9} /* (27, 3, 10) {real, imag} */,
  {32'h3ec9c73a, 32'h3f1171e1} /* (27, 3, 9) {real, imag} */,
  {32'hbeb5d000, 32'h3b6ec340} /* (27, 3, 8) {real, imag} */,
  {32'h3e2bba19, 32'h3eccc0e3} /* (27, 3, 7) {real, imag} */,
  {32'hbf6cf93a, 32'hbe2967a6} /* (27, 3, 6) {real, imag} */,
  {32'h3ea33c8c, 32'h3db2b51a} /* (27, 3, 5) {real, imag} */,
  {32'hbd435610, 32'h3f763c0a} /* (27, 3, 4) {real, imag} */,
  {32'hbde9513e, 32'h3e87f9b4} /* (27, 3, 3) {real, imag} */,
  {32'hbd4388a0, 32'hc025c636} /* (27, 3, 2) {real, imag} */,
  {32'h3fdc4ef9, 32'h406695fb} /* (27, 3, 1) {real, imag} */,
  {32'h3fde5ea8, 32'h3e9ca644} /* (27, 3, 0) {real, imag} */,
  {32'hc15b2dce, 32'h3fbd744f} /* (27, 2, 31) {real, imag} */,
  {32'h411da3ec, 32'hc0659e92} /* (27, 2, 30) {real, imag} */,
  {32'hbf3458b2, 32'h3d1d2510} /* (27, 2, 29) {real, imag} */,
  {32'hbf1e34d9, 32'h40275e12} /* (27, 2, 28) {real, imag} */,
  {32'h3f8615a2, 32'hbfadbd5b} /* (27, 2, 27) {real, imag} */,
  {32'h3e84fa0c, 32'hbe6894fb} /* (27, 2, 26) {real, imag} */,
  {32'hbd5e9688, 32'h3f818f7b} /* (27, 2, 25) {real, imag} */,
  {32'h3ee2d8ce, 32'hbf1d7c5a} /* (27, 2, 24) {real, imag} */,
  {32'h3eecfb96, 32'h3db3add3} /* (27, 2, 23) {real, imag} */,
  {32'hbe801b4f, 32'hbeb7e102} /* (27, 2, 22) {real, imag} */,
  {32'h3d6adc14, 32'hbe581515} /* (27, 2, 21) {real, imag} */,
  {32'h3e9c30e8, 32'h3e49bfb0} /* (27, 2, 20) {real, imag} */,
  {32'hbdb78b54, 32'hbd9c10a8} /* (27, 2, 19) {real, imag} */,
  {32'h3ea31dcf, 32'hbe90e1da} /* (27, 2, 18) {real, imag} */,
  {32'h3f00a813, 32'h3e7d52f0} /* (27, 2, 17) {real, imag} */,
  {32'hbe88eb1d, 32'hbd0bdd5c} /* (27, 2, 16) {real, imag} */,
  {32'h3d002f60, 32'h3b4af2e0} /* (27, 2, 15) {real, imag} */,
  {32'h3e1c1d65, 32'hbd105c88} /* (27, 2, 14) {real, imag} */,
  {32'h3cfffe46, 32'hbebd37d2} /* (27, 2, 13) {real, imag} */,
  {32'hbee6fa1c, 32'h3e19587e} /* (27, 2, 12) {real, imag} */,
  {32'hbea115d8, 32'h3f318e1e} /* (27, 2, 11) {real, imag} */,
  {32'hbea6da20, 32'hbf07c0b5} /* (27, 2, 10) {real, imag} */,
  {32'h3e330e99, 32'h3d179090} /* (27, 2, 9) {real, imag} */,
  {32'h3f1939e4, 32'h3f3e9ff9} /* (27, 2, 8) {real, imag} */,
  {32'hbe847546, 32'hbddc2ea0} /* (27, 2, 7) {real, imag} */,
  {32'hbd24b296, 32'hbe067122} /* (27, 2, 6) {real, imag} */,
  {32'h3f5c2f2b, 32'h3f94c5a7} /* (27, 2, 5) {real, imag} */,
  {32'hc008be87, 32'hbfdc77a4} /* (27, 2, 4) {real, imag} */,
  {32'h3d8c2e84, 32'hbeefbccf} /* (27, 2, 3) {real, imag} */,
  {32'h410100c2, 32'hc0563fb4} /* (27, 2, 2) {real, imag} */,
  {32'hc10244db, 32'h406b4504} /* (27, 2, 1) {real, imag} */,
  {32'hc0ce7eff, 32'hc059d8f0} /* (27, 2, 0) {real, imag} */,
  {32'h411803d0, 32'hc07c004e} /* (27, 1, 31) {real, imag} */,
  {32'hc0a180c4, 32'h40062957} /* (27, 1, 30) {real, imag} */,
  {32'h3e41b018, 32'h3e45ff42} /* (27, 1, 29) {real, imag} */,
  {32'h3ec18f7f, 32'h3f6d56af} /* (27, 1, 28) {real, imag} */,
  {32'hc049c86f, 32'h3e74bf50} /* (27, 1, 27) {real, imag} */,
  {32'hbea5eea1, 32'hbf0ea87b} /* (27, 1, 26) {real, imag} */,
  {32'h3e99fb76, 32'h3eb57ac6} /* (27, 1, 25) {real, imag} */,
  {32'h3d3b9ab8, 32'h3ebad6a3} /* (27, 1, 24) {real, imag} */,
  {32'hbe735c0a, 32'hbf1dab4e} /* (27, 1, 23) {real, imag} */,
  {32'hbdd1c792, 32'hbe10aebb} /* (27, 1, 22) {real, imag} */,
  {32'hbf816acc, 32'h3e9163da} /* (27, 1, 21) {real, imag} */,
  {32'hbdc4237e, 32'h3f2d64e8} /* (27, 1, 20) {real, imag} */,
  {32'h3d3e4c1e, 32'hbf057a26} /* (27, 1, 19) {real, imag} */,
  {32'h3ebbf42a, 32'h3e750aae} /* (27, 1, 18) {real, imag} */,
  {32'hbc94e0e8, 32'h3e0538c1} /* (27, 1, 17) {real, imag} */,
  {32'hbe04dd01, 32'hbe05ad3f} /* (27, 1, 16) {real, imag} */,
  {32'hbe9017c2, 32'h3eefa48c} /* (27, 1, 15) {real, imag} */,
  {32'h3ed3acdd, 32'hbef1b2f5} /* (27, 1, 14) {real, imag} */,
  {32'h3f0823dd, 32'hbd10da8c} /* (27, 1, 13) {real, imag} */,
  {32'hbeb213de, 32'h3d6b1ff4} /* (27, 1, 12) {real, imag} */,
  {32'hbf0df652, 32'hbecde1ac} /* (27, 1, 11) {real, imag} */,
  {32'hbc844ed0, 32'h3f32fc27} /* (27, 1, 10) {real, imag} */,
  {32'hbf3191f8, 32'hbed74fff} /* (27, 1, 9) {real, imag} */,
  {32'hbedb6946, 32'hbf7c1033} /* (27, 1, 8) {real, imag} */,
  {32'hbf1960fd, 32'h3e8c7ef0} /* (27, 1, 7) {real, imag} */,
  {32'hbe46a3e6, 32'hbec1f8f7} /* (27, 1, 6) {real, imag} */,
  {32'hbfe28a12, 32'hbf61ba4d} /* (27, 1, 5) {real, imag} */,
  {32'h3f77485f, 32'h3f1830e3} /* (27, 1, 4) {real, imag} */,
  {32'hbfc2ca0c, 32'hbe9fcc40} /* (27, 1, 3) {real, imag} */,
  {32'hc10eb0ba, 32'hc10aeec8} /* (27, 1, 2) {real, imag} */,
  {32'h4150e7c2, 32'h40b24765} /* (27, 1, 1) {real, imag} */,
  {32'h4083ac36, 32'hbe197190} /* (27, 1, 0) {real, imag} */,
  {32'hbfa2ca40, 32'h3f7603d8} /* (27, 0, 31) {real, imag} */,
  {32'hc01db0b6, 32'h40b591de} /* (27, 0, 30) {real, imag} */,
  {32'hbea0984c, 32'hbfbb3c02} /* (27, 0, 29) {real, imag} */,
  {32'h3f82a9ba, 32'h3f285bdc} /* (27, 0, 28) {real, imag} */,
  {32'hbfea827e, 32'h3f82a4ca} /* (27, 0, 27) {real, imag} */,
  {32'h3f315af5, 32'h3e173e8e} /* (27, 0, 26) {real, imag} */,
  {32'h3f178ccf, 32'hbf947a70} /* (27, 0, 25) {real, imag} */,
  {32'hbe300df0, 32'h3f9a87bc} /* (27, 0, 24) {real, imag} */,
  {32'hbecba551, 32'hbd37a948} /* (27, 0, 23) {real, imag} */,
  {32'hbec93bda, 32'h3ed58b32} /* (27, 0, 22) {real, imag} */,
  {32'h3dc72106, 32'h3ea5794e} /* (27, 0, 21) {real, imag} */,
  {32'h3e8588f8, 32'h3d555a2c} /* (27, 0, 20) {real, imag} */,
  {32'h3e3bcdfd, 32'hbdc2d058} /* (27, 0, 19) {real, imag} */,
  {32'h3ed73f26, 32'h3e55ec14} /* (27, 0, 18) {real, imag} */,
  {32'h3e5d1e78, 32'hbd31b466} /* (27, 0, 17) {real, imag} */,
  {32'hbeafdd7c, 32'h00000000} /* (27, 0, 16) {real, imag} */,
  {32'h3e5d1e78, 32'h3d31b466} /* (27, 0, 15) {real, imag} */,
  {32'h3ed73f26, 32'hbe55ec14} /* (27, 0, 14) {real, imag} */,
  {32'h3e3bcdfd, 32'h3dc2d058} /* (27, 0, 13) {real, imag} */,
  {32'h3e8588f8, 32'hbd555a2c} /* (27, 0, 12) {real, imag} */,
  {32'h3dc72106, 32'hbea5794e} /* (27, 0, 11) {real, imag} */,
  {32'hbec93bda, 32'hbed58b32} /* (27, 0, 10) {real, imag} */,
  {32'hbecba551, 32'h3d37a948} /* (27, 0, 9) {real, imag} */,
  {32'hbe300df0, 32'hbf9a87bc} /* (27, 0, 8) {real, imag} */,
  {32'h3f178ccf, 32'h3f947a70} /* (27, 0, 7) {real, imag} */,
  {32'h3f315af5, 32'hbe173e8e} /* (27, 0, 6) {real, imag} */,
  {32'hbfea827e, 32'hbf82a4ca} /* (27, 0, 5) {real, imag} */,
  {32'h3f82a9ba, 32'hbf285bdc} /* (27, 0, 4) {real, imag} */,
  {32'hbea0984c, 32'h3fbb3c02} /* (27, 0, 3) {real, imag} */,
  {32'hc01db0b6, 32'hc0b591de} /* (27, 0, 2) {real, imag} */,
  {32'hbfa2ca40, 32'hbf7603d8} /* (27, 0, 1) {real, imag} */,
  {32'hc15271ac, 32'h00000000} /* (27, 0, 0) {real, imag} */,
  {32'hc1110940, 32'h40dc801d} /* (26, 31, 31) {real, imag} */,
  {32'hbf7ce798, 32'h3f8169f4} /* (26, 31, 30) {real, imag} */,
  {32'h3be7c600, 32'h3f330c6c} /* (26, 31, 29) {real, imag} */,
  {32'hbf12dc72, 32'h3f00c656} /* (26, 31, 28) {real, imag} */,
  {32'h3d6f3620, 32'hbea47a2e} /* (26, 31, 27) {real, imag} */,
  {32'h3eef0c36, 32'h3daae662} /* (26, 31, 26) {real, imag} */,
  {32'h3eb69168, 32'hbf26c130} /* (26, 31, 25) {real, imag} */,
  {32'hbeab1098, 32'h3f1a6005} /* (26, 31, 24) {real, imag} */,
  {32'hbf2e7514, 32'hbd143fe0} /* (26, 31, 23) {real, imag} */,
  {32'hbf5ccbee, 32'hbc483278} /* (26, 31, 22) {real, imag} */,
  {32'hbf1d1598, 32'hbd032e10} /* (26, 31, 21) {real, imag} */,
  {32'h3e8907c2, 32'hbeca5faa} /* (26, 31, 20) {real, imag} */,
  {32'h3f595d35, 32'hbe129d18} /* (26, 31, 19) {real, imag} */,
  {32'h3dfe397a, 32'h3e23ba98} /* (26, 31, 18) {real, imag} */,
  {32'hbb64a4c0, 32'h3d080bcc} /* (26, 31, 17) {real, imag} */,
  {32'hbe7f199a, 32'h3d6a115d} /* (26, 31, 16) {real, imag} */,
  {32'h3e03bd20, 32'h3e7c0667} /* (26, 31, 15) {real, imag} */,
  {32'h3eb03ef8, 32'hbd35c9a4} /* (26, 31, 14) {real, imag} */,
  {32'h3f050d11, 32'h3e3e3764} /* (26, 31, 13) {real, imag} */,
  {32'h3eb9e5a6, 32'hbf08db82} /* (26, 31, 12) {real, imag} */,
  {32'hbd65da08, 32'h3eb55303} /* (26, 31, 11) {real, imag} */,
  {32'h3d813678, 32'hbe2848ee} /* (26, 31, 10) {real, imag} */,
  {32'h3e8e2b92, 32'hbbf921c0} /* (26, 31, 9) {real, imag} */,
  {32'h3e857d44, 32'h3e0516f1} /* (26, 31, 8) {real, imag} */,
  {32'hbe4ce52e, 32'h3ea8f8e9} /* (26, 31, 7) {real, imag} */,
  {32'hbf560d2d, 32'h3e81b218} /* (26, 31, 6) {real, imag} */,
  {32'hbf147850, 32'h3bc16300} /* (26, 31, 5) {real, imag} */,
  {32'hbee9817a, 32'hbf141052} /* (26, 31, 4) {real, imag} */,
  {32'h3e6986d4, 32'h3d490a00} /* (26, 31, 3) {real, imag} */,
  {32'h3efa1570, 32'hc058bf26} /* (26, 31, 2) {real, imag} */,
  {32'hc0d6de14, 32'hbd8695e0} /* (26, 31, 1) {real, imag} */,
  {32'hc168fd6c, 32'h4053370a} /* (26, 31, 0) {real, imag} */,
  {32'h3e359680, 32'hc008b118} /* (26, 30, 31) {real, imag} */,
  {32'h40061f12, 32'h3f5c8ee8} /* (26, 30, 30) {real, imag} */,
  {32'hbf7537d2, 32'h3eb5a3bb} /* (26, 30, 29) {real, imag} */,
  {32'hbf114d0c, 32'h3f94c973} /* (26, 30, 28) {real, imag} */,
  {32'hbf13011d, 32'hbfa263f2} /* (26, 30, 27) {real, imag} */,
  {32'h3ee09cbe, 32'hbe43c967} /* (26, 30, 26) {real, imag} */,
  {32'h3e4ef612, 32'hbf4366d6} /* (26, 30, 25) {real, imag} */,
  {32'hbe145796, 32'hbf28f5c5} /* (26, 30, 24) {real, imag} */,
  {32'hbf14259f, 32'h3ed2f550} /* (26, 30, 23) {real, imag} */,
  {32'h3c5b00b0, 32'hbd99b554} /* (26, 30, 22) {real, imag} */,
  {32'h3edede48, 32'hbe8115e9} /* (26, 30, 21) {real, imag} */,
  {32'h3e3793f8, 32'hbd879494} /* (26, 30, 20) {real, imag} */,
  {32'hbdefe79e, 32'hbd790ac2} /* (26, 30, 19) {real, imag} */,
  {32'hbe026a38, 32'h3e6aaffa} /* (26, 30, 18) {real, imag} */,
  {32'hbceed506, 32'h3e448894} /* (26, 30, 17) {real, imag} */,
  {32'h3d9e675e, 32'hbe39f76d} /* (26, 30, 16) {real, imag} */,
  {32'h3e9aa0ae, 32'hbe7dfd77} /* (26, 30, 15) {real, imag} */,
  {32'h3e9b1964, 32'hbec0c8cf} /* (26, 30, 14) {real, imag} */,
  {32'hbe766dda, 32'h3d0b2cb8} /* (26, 30, 13) {real, imag} */,
  {32'hbe70bd3f, 32'h3c738940} /* (26, 30, 12) {real, imag} */,
  {32'h3e039c7c, 32'hbd3ffd80} /* (26, 30, 11) {real, imag} */,
  {32'hbec06eb2, 32'h3db6331e} /* (26, 30, 10) {real, imag} */,
  {32'h3f65fcf9, 32'h3eeee2d3} /* (26, 30, 9) {real, imag} */,
  {32'h3f2afec6, 32'hbea8d31d} /* (26, 30, 8) {real, imag} */,
  {32'hbe3ffe56, 32'hbfa1b930} /* (26, 30, 7) {real, imag} */,
  {32'h3e34bb75, 32'hbedf0e50} /* (26, 30, 6) {real, imag} */,
  {32'h3f6b715f, 32'h3f3ef157} /* (26, 30, 5) {real, imag} */,
  {32'hbec1df94, 32'hbeb3531a} /* (26, 30, 4) {real, imag} */,
  {32'hbeb4a8ec, 32'h3e68e93e} /* (26, 30, 3) {real, imag} */,
  {32'h3fe2fe10, 32'h3ff918f2} /* (26, 30, 2) {real, imag} */,
  {32'h3f35c9e0, 32'hbff760bc} /* (26, 30, 1) {real, imag} */,
  {32'h3fd3d7cc, 32'h400b7808} /* (26, 30, 0) {real, imag} */,
  {32'hbde03680, 32'hc014a578} /* (26, 29, 31) {real, imag} */,
  {32'h3f52df75, 32'h3e75bf94} /* (26, 29, 30) {real, imag} */,
  {32'hbf029350, 32'h3cd002e0} /* (26, 29, 29) {real, imag} */,
  {32'hbe3efcea, 32'hbee4205d} /* (26, 29, 28) {real, imag} */,
  {32'hbef03418, 32'hbed9f036} /* (26, 29, 27) {real, imag} */,
  {32'hbee8f290, 32'hbedbf076} /* (26, 29, 26) {real, imag} */,
  {32'hbdf6243c, 32'hbeea9a5a} /* (26, 29, 25) {real, imag} */,
  {32'hbe6ee221, 32'h3ecd4281} /* (26, 29, 24) {real, imag} */,
  {32'hbe0c4b2c, 32'h3e7e9390} /* (26, 29, 23) {real, imag} */,
  {32'hbe88d650, 32'h3dc4720a} /* (26, 29, 22) {real, imag} */,
  {32'h3d801bc2, 32'h3e236302} /* (26, 29, 21) {real, imag} */,
  {32'h3e7e260e, 32'h3e972ce0} /* (26, 29, 20) {real, imag} */,
  {32'h3ea11535, 32'h3f0d7278} /* (26, 29, 19) {real, imag} */,
  {32'h3dcc7684, 32'hbf0498f4} /* (26, 29, 18) {real, imag} */,
  {32'hbe10ab61, 32'h3e4e1dc2} /* (26, 29, 17) {real, imag} */,
  {32'h3e076e9e, 32'hbe8184ef} /* (26, 29, 16) {real, imag} */,
  {32'h3f1344da, 32'hbe52d840} /* (26, 29, 15) {real, imag} */,
  {32'hbea8e9d6, 32'h3f1d1ad3} /* (26, 29, 14) {real, imag} */,
  {32'h3ec3a574, 32'h3e4c9c4c} /* (26, 29, 13) {real, imag} */,
  {32'hbeb7af6a, 32'h3df3e51a} /* (26, 29, 12) {real, imag} */,
  {32'h3c9af8c0, 32'hbe29174a} /* (26, 29, 11) {real, imag} */,
  {32'hbd83b432, 32'hbe2bd33f} /* (26, 29, 10) {real, imag} */,
  {32'h3e4392fb, 32'h3e9680ba} /* (26, 29, 9) {real, imag} */,
  {32'hbe60c97e, 32'h3eba0988} /* (26, 29, 8) {real, imag} */,
  {32'hbf2f19f9, 32'hbd0f2c90} /* (26, 29, 7) {real, imag} */,
  {32'hbea94fdf, 32'hbedd9480} /* (26, 29, 6) {real, imag} */,
  {32'hbd96b900, 32'h3e7044af} /* (26, 29, 5) {real, imag} */,
  {32'h3f1f5ad8, 32'hbf0a913f} /* (26, 29, 4) {real, imag} */,
  {32'h3eabdac1, 32'hbd84177e} /* (26, 29, 3) {real, imag} */,
  {32'h3fc90e17, 32'h3edf3e10} /* (26, 29, 2) {real, imag} */,
  {32'hbf57bc14, 32'hbe117fc8} /* (26, 29, 1) {real, imag} */,
  {32'h401e92db, 32'hbf7d20d5} /* (26, 29, 0) {real, imag} */,
  {32'h3ed80fc8, 32'hbeb5c77a} /* (26, 28, 31) {real, imag} */,
  {32'hbee73dec, 32'h3e08d008} /* (26, 28, 30) {real, imag} */,
  {32'hbdc716f6, 32'h3e0587e6} /* (26, 28, 29) {real, imag} */,
  {32'h3f2e8843, 32'h3f6872be} /* (26, 28, 28) {real, imag} */,
  {32'h3edaaf09, 32'h3d2faf24} /* (26, 28, 27) {real, imag} */,
  {32'hbf178266, 32'hbe9c6e08} /* (26, 28, 26) {real, imag} */,
  {32'hbda0d54c, 32'hbeca25f4} /* (26, 28, 25) {real, imag} */,
  {32'h3d8c760c, 32'h3e908507} /* (26, 28, 24) {real, imag} */,
  {32'hbe3a6adf, 32'hbdc6e62c} /* (26, 28, 23) {real, imag} */,
  {32'h3e056319, 32'h3e261476} /* (26, 28, 22) {real, imag} */,
  {32'h3f255f87, 32'hbe992c14} /* (26, 28, 21) {real, imag} */,
  {32'hbebca03f, 32'h3e97b227} /* (26, 28, 20) {real, imag} */,
  {32'h3dc4e50e, 32'hbeb86426} /* (26, 28, 19) {real, imag} */,
  {32'hbe835352, 32'hbd3cd410} /* (26, 28, 18) {real, imag} */,
  {32'hbef50474, 32'h3e058686} /* (26, 28, 17) {real, imag} */,
  {32'hbe15c904, 32'h3d3ce1d4} /* (26, 28, 16) {real, imag} */,
  {32'h3e3946b8, 32'h3d4985fc} /* (26, 28, 15) {real, imag} */,
  {32'hbf1eec98, 32'h3e903573} /* (26, 28, 14) {real, imag} */,
  {32'hbc54757e, 32'h3e4b3a8b} /* (26, 28, 13) {real, imag} */,
  {32'h3e203a5c, 32'hbd9e0994} /* (26, 28, 12) {real, imag} */,
  {32'hbe271056, 32'hbf22e4f0} /* (26, 28, 11) {real, imag} */,
  {32'h3f3acb31, 32'hbe8cd3cf} /* (26, 28, 10) {real, imag} */,
  {32'hbb3ba040, 32'hbe8e73ad} /* (26, 28, 9) {real, imag} */,
  {32'h3db5ab34, 32'h3eb27150} /* (26, 28, 8) {real, imag} */,
  {32'hbd3bdcce, 32'hbf96858b} /* (26, 28, 7) {real, imag} */,
  {32'hbf405772, 32'h3ed577c5} /* (26, 28, 6) {real, imag} */,
  {32'h3cfb8754, 32'hbe0909d3} /* (26, 28, 5) {real, imag} */,
  {32'h3cb463f0, 32'h3eaaf775} /* (26, 28, 4) {real, imag} */,
  {32'hbf44089d, 32'hbda2a804} /* (26, 28, 3) {real, imag} */,
  {32'hbeb5daee, 32'h3e0d1a58} /* (26, 28, 2) {real, imag} */,
  {32'hbec5a5e2, 32'h3d869b28} /* (26, 28, 1) {real, imag} */,
  {32'hbf2c42ca, 32'h3f7c5812} /* (26, 28, 0) {real, imag} */,
  {32'hbf8a3bc1, 32'hbea24b98} /* (26, 27, 31) {real, imag} */,
  {32'hbf1275bd, 32'h3eb67f6a} /* (26, 27, 30) {real, imag} */,
  {32'hbee61926, 32'h3f3aee14} /* (26, 27, 29) {real, imag} */,
  {32'hbdf14a65, 32'h3e80f6d3} /* (26, 27, 28) {real, imag} */,
  {32'h3ef9b22f, 32'hbd3681c0} /* (26, 27, 27) {real, imag} */,
  {32'hbf3b1a1a, 32'hbee1ca44} /* (26, 27, 26) {real, imag} */,
  {32'h3f1a4e22, 32'hbeead4a6} /* (26, 27, 25) {real, imag} */,
  {32'h3f53f6e6, 32'h3e5b83d6} /* (26, 27, 24) {real, imag} */,
  {32'h3ebbe2b8, 32'h3c82f2b0} /* (26, 27, 23) {real, imag} */,
  {32'h3e9af272, 32'hbde562d2} /* (26, 27, 22) {real, imag} */,
  {32'h3dde159d, 32'hbf0b5dbe} /* (26, 27, 21) {real, imag} */,
  {32'hbe086714, 32'hbcb91f70} /* (26, 27, 20) {real, imag} */,
  {32'hbeb8e9fa, 32'hbef44ae4} /* (26, 27, 19) {real, imag} */,
  {32'hbe04cea8, 32'h3c732e20} /* (26, 27, 18) {real, imag} */,
  {32'hbdd9c69c, 32'hbd8683e4} /* (26, 27, 17) {real, imag} */,
  {32'hbec34b38, 32'h3efb725a} /* (26, 27, 16) {real, imag} */,
  {32'h3d15362c, 32'h3e8950ce} /* (26, 27, 15) {real, imag} */,
  {32'h3e5b013e, 32'h3ea715ae} /* (26, 27, 14) {real, imag} */,
  {32'h3e8ab40e, 32'hbefecbca} /* (26, 27, 13) {real, imag} */,
  {32'h3f1e6ae0, 32'hbe1c0209} /* (26, 27, 12) {real, imag} */,
  {32'h3ddbec2a, 32'h3ece430a} /* (26, 27, 11) {real, imag} */,
  {32'h3ee173d6, 32'h3b224080} /* (26, 27, 10) {real, imag} */,
  {32'hbed80ee4, 32'hbed8e888} /* (26, 27, 9) {real, imag} */,
  {32'h3d78d904, 32'h3e2b74c9} /* (26, 27, 8) {real, imag} */,
  {32'h3d523fa2, 32'h3eb11360} /* (26, 27, 7) {real, imag} */,
  {32'h3e067d77, 32'h3d1902e2} /* (26, 27, 6) {real, imag} */,
  {32'hbef5a32e, 32'h3ea2b9dc} /* (26, 27, 5) {real, imag} */,
  {32'hbebbbcf3, 32'hbf2e4bd0} /* (26, 27, 4) {real, imag} */,
  {32'h3f57bcd2, 32'hbd84fff4} /* (26, 27, 3) {real, imag} */,
  {32'h3f0ed5a4, 32'h3ea4b4dc} /* (26, 27, 2) {real, imag} */,
  {32'hbdd94940, 32'h3f9dd99e} /* (26, 27, 1) {real, imag} */,
  {32'hbfd69100, 32'hbf24f675} /* (26, 27, 0) {real, imag} */,
  {32'hbe4004ec, 32'hbe857943} /* (26, 26, 31) {real, imag} */,
  {32'h3e8e4984, 32'hbd80b062} /* (26, 26, 30) {real, imag} */,
  {32'h3f2137d9, 32'h3ee20997} /* (26, 26, 29) {real, imag} */,
  {32'hbe436798, 32'h3ee14baa} /* (26, 26, 28) {real, imag} */,
  {32'h3d1778f8, 32'hbed8a6c5} /* (26, 26, 27) {real, imag} */,
  {32'h3f108912, 32'h3f01811d} /* (26, 26, 26) {real, imag} */,
  {32'h3ea518f8, 32'hbd13e8c0} /* (26, 26, 25) {real, imag} */,
  {32'h3f0e19d2, 32'hbea38252} /* (26, 26, 24) {real, imag} */,
  {32'h3f22bcbd, 32'h3ed876c0} /* (26, 26, 23) {real, imag} */,
  {32'hbe1d473b, 32'hbd7eb7f8} /* (26, 26, 22) {real, imag} */,
  {32'h3ef8b646, 32'h3e127c61} /* (26, 26, 21) {real, imag} */,
  {32'hbedb3124, 32'hbed31ff6} /* (26, 26, 20) {real, imag} */,
  {32'h3ecaf7d5, 32'h3ecb920b} /* (26, 26, 19) {real, imag} */,
  {32'h3e0e04ee, 32'h3bffcf08} /* (26, 26, 18) {real, imag} */,
  {32'h3e46ad99, 32'hbe0c0473} /* (26, 26, 17) {real, imag} */,
  {32'h3e582811, 32'hbda58bd4} /* (26, 26, 16) {real, imag} */,
  {32'hbe8e9852, 32'h3ed5e600} /* (26, 26, 15) {real, imag} */,
  {32'h3dc01351, 32'hbeaecd0c} /* (26, 26, 14) {real, imag} */,
  {32'hbe6f3dc3, 32'h3eb6cda9} /* (26, 26, 13) {real, imag} */,
  {32'h3e90852e, 32'hbe604f39} /* (26, 26, 12) {real, imag} */,
  {32'h3e2a9500, 32'h3db7bd48} /* (26, 26, 11) {real, imag} */,
  {32'h3f0a8a17, 32'hbe9c2d76} /* (26, 26, 10) {real, imag} */,
  {32'h3ce2ac38, 32'h3dbb0c4a} /* (26, 26, 9) {real, imag} */,
  {32'h3e69228a, 32'hbf7cf696} /* (26, 26, 8) {real, imag} */,
  {32'hbed5871f, 32'h3ec97a98} /* (26, 26, 7) {real, imag} */,
  {32'h3d76b1a8, 32'hbf2d71cd} /* (26, 26, 6) {real, imag} */,
  {32'hbd59ea4c, 32'hbd38ed48} /* (26, 26, 5) {real, imag} */,
  {32'h3eb56916, 32'h3ee319dd} /* (26, 26, 4) {real, imag} */,
  {32'hbd91ce2a, 32'hbe1b32d6} /* (26, 26, 3) {real, imag} */,
  {32'hbf2f530d, 32'hbd97ec3c} /* (26, 26, 2) {real, imag} */,
  {32'hbed6d6fe, 32'hbda291d0} /* (26, 26, 1) {real, imag} */,
  {32'h3ed62ce8, 32'h3efb96c0} /* (26, 26, 0) {real, imag} */,
  {32'h3f819004, 32'hbe811cea} /* (26, 25, 31) {real, imag} */,
  {32'h3ea7aad6, 32'hbf24ae94} /* (26, 25, 30) {real, imag} */,
  {32'h3f361906, 32'h3e015854} /* (26, 25, 29) {real, imag} */,
  {32'h3e911ffa, 32'h3f8d3dca} /* (26, 25, 28) {real, imag} */,
  {32'hbeb16552, 32'h3f0c6381} /* (26, 25, 27) {real, imag} */,
  {32'h3f23e214, 32'hbee52827} /* (26, 25, 26) {real, imag} */,
  {32'hbea10d75, 32'h3e893c50} /* (26, 25, 25) {real, imag} */,
  {32'h3e9baaf6, 32'h3f1c95f7} /* (26, 25, 24) {real, imag} */,
  {32'h3ef15f48, 32'hbeb859de} /* (26, 25, 23) {real, imag} */,
  {32'hbf55f7ba, 32'h3ec8deb6} /* (26, 25, 22) {real, imag} */,
  {32'hbe4a93f0, 32'hbf00c998} /* (26, 25, 21) {real, imag} */,
  {32'h3cad3028, 32'h3e8aeb84} /* (26, 25, 20) {real, imag} */,
  {32'hbe145503, 32'h3d6e6d0a} /* (26, 25, 19) {real, imag} */,
  {32'hbf0daa64, 32'h3d66ab3b} /* (26, 25, 18) {real, imag} */,
  {32'h3d8bc6b4, 32'hbd14ae44} /* (26, 25, 17) {real, imag} */,
  {32'hbea66cd6, 32'h3db9db67} /* (26, 25, 16) {real, imag} */,
  {32'hbdac6782, 32'hbd028cae} /* (26, 25, 15) {real, imag} */,
  {32'hbece3674, 32'hbe904ae8} /* (26, 25, 14) {real, imag} */,
  {32'hbe839bfe, 32'hbea33ede} /* (26, 25, 13) {real, imag} */,
  {32'h3f21a452, 32'hbeb8a6ea} /* (26, 25, 12) {real, imag} */,
  {32'h3c597660, 32'h3f1b5a6c} /* (26, 25, 11) {real, imag} */,
  {32'hbd4caf44, 32'hbf058e57} /* (26, 25, 10) {real, imag} */,
  {32'hbe8405ea, 32'hbf093669} /* (26, 25, 9) {real, imag} */,
  {32'h3eb70ab3, 32'h3f5c250c} /* (26, 25, 8) {real, imag} */,
  {32'h3c85bd58, 32'h3dc3c430} /* (26, 25, 7) {real, imag} */,
  {32'hbdc2a6e4, 32'hbf1a4a94} /* (26, 25, 6) {real, imag} */,
  {32'h3eff5eab, 32'hbf1a7957} /* (26, 25, 5) {real, imag} */,
  {32'hbe212fc0, 32'hbe024eb0} /* (26, 25, 4) {real, imag} */,
  {32'h3de5c368, 32'h3f0bdd00} /* (26, 25, 3) {real, imag} */,
  {32'hbe2568ea, 32'h3e3e00ce} /* (26, 25, 2) {real, imag} */,
  {32'hbf4d02ca, 32'hbe31503e} /* (26, 25, 1) {real, imag} */,
  {32'hbf1c5b62, 32'hbd009baa} /* (26, 25, 0) {real, imag} */,
  {32'hbdec2ee0, 32'h3e154f88} /* (26, 24, 31) {real, imag} */,
  {32'hbf19902f, 32'h3e316dec} /* (26, 24, 30) {real, imag} */,
  {32'h3f4b5d50, 32'hbf664b8a} /* (26, 24, 29) {real, imag} */,
  {32'hbf2edd4e, 32'hbeedd199} /* (26, 24, 28) {real, imag} */,
  {32'h3ecffc8f, 32'hbc0a0828} /* (26, 24, 27) {real, imag} */,
  {32'h3dfa1a24, 32'hbc7a93c8} /* (26, 24, 26) {real, imag} */,
  {32'h3f285fdd, 32'h3dc430ba} /* (26, 24, 25) {real, imag} */,
  {32'hbf0c4e9a, 32'h3f0c6f4e} /* (26, 24, 24) {real, imag} */,
  {32'h3e2edc9c, 32'hbe654afa} /* (26, 24, 23) {real, imag} */,
  {32'hbee556d4, 32'h3eac036a} /* (26, 24, 22) {real, imag} */,
  {32'h3eb2fe28, 32'h3e5cb0d9} /* (26, 24, 21) {real, imag} */,
  {32'h3cfdd9de, 32'h3d558734} /* (26, 24, 20) {real, imag} */,
  {32'h3e9836aa, 32'hbe11c576} /* (26, 24, 19) {real, imag} */,
  {32'h3dcf2a30, 32'hbe31f37a} /* (26, 24, 18) {real, imag} */,
  {32'h3e7442d3, 32'hbd48c350} /* (26, 24, 17) {real, imag} */,
  {32'h3dfe6c3e, 32'hbdd3c554} /* (26, 24, 16) {real, imag} */,
  {32'h3d7d60b4, 32'hbeb09f67} /* (26, 24, 15) {real, imag} */,
  {32'hbe222ae0, 32'hbdbc2d25} /* (26, 24, 14) {real, imag} */,
  {32'hbf147d64, 32'h3d4f93d4} /* (26, 24, 13) {real, imag} */,
  {32'h3e3fa957, 32'hbeb2b9f2} /* (26, 24, 12) {real, imag} */,
  {32'h3bc45880, 32'h3ed75176} /* (26, 24, 11) {real, imag} */,
  {32'h3c3970e0, 32'h3dc515ec} /* (26, 24, 10) {real, imag} */,
  {32'hbe68adf0, 32'h3e83859c} /* (26, 24, 9) {real, imag} */,
  {32'h3f72ee4d, 32'hbe60e254} /* (26, 24, 8) {real, imag} */,
  {32'h3e37418c, 32'h3e915e8f} /* (26, 24, 7) {real, imag} */,
  {32'hbf14bf92, 32'hbf2135f8} /* (26, 24, 6) {real, imag} */,
  {32'hbef31677, 32'hbe8b9ed2} /* (26, 24, 5) {real, imag} */,
  {32'hbd7c5cf0, 32'hbe8ba91c} /* (26, 24, 4) {real, imag} */,
  {32'hbe6586c8, 32'h3ea37e35} /* (26, 24, 3) {real, imag} */,
  {32'h3e8146c1, 32'h3cd93bc4} /* (26, 24, 2) {real, imag} */,
  {32'h3d34f5b8, 32'h3f20619d} /* (26, 24, 1) {real, imag} */,
  {32'hbe7b99ca, 32'h3dd622e0} /* (26, 24, 0) {real, imag} */,
  {32'h3e766a80, 32'h3f03b103} /* (26, 23, 31) {real, imag} */,
  {32'h3e9e6240, 32'h3f01b1d4} /* (26, 23, 30) {real, imag} */,
  {32'hbe6035e4, 32'h3e738ef4} /* (26, 23, 29) {real, imag} */,
  {32'h3d6d7868, 32'hbeaac05d} /* (26, 23, 28) {real, imag} */,
  {32'h3ed886c1, 32'hbf496e64} /* (26, 23, 27) {real, imag} */,
  {32'h3ee18bc8, 32'hbe7cef79} /* (26, 23, 26) {real, imag} */,
  {32'h3e135104, 32'hbec91233} /* (26, 23, 25) {real, imag} */,
  {32'h3d337f60, 32'h3f2ee746} /* (26, 23, 24) {real, imag} */,
  {32'h3c151d80, 32'hbe202954} /* (26, 23, 23) {real, imag} */,
  {32'hbdc2a731, 32'hbddc49b8} /* (26, 23, 22) {real, imag} */,
  {32'h3dccd736, 32'hbed71efe} /* (26, 23, 21) {real, imag} */,
  {32'h3e0249d4, 32'hbd607770} /* (26, 23, 20) {real, imag} */,
  {32'h3c309090, 32'hbe320f2b} /* (26, 23, 19) {real, imag} */,
  {32'hbe195e93, 32'hbe184899} /* (26, 23, 18) {real, imag} */,
  {32'hbb716f80, 32'h3ed8731b} /* (26, 23, 17) {real, imag} */,
  {32'h3dfd3eb4, 32'hbe25602d} /* (26, 23, 16) {real, imag} */,
  {32'h3d01eb24, 32'h3e1f4ecd} /* (26, 23, 15) {real, imag} */,
  {32'hbae87780, 32'h3d6918f8} /* (26, 23, 14) {real, imag} */,
  {32'h3e6027b4, 32'hbd3d7e40} /* (26, 23, 13) {real, imag} */,
  {32'hbef98553, 32'hbeb64fd9} /* (26, 23, 12) {real, imag} */,
  {32'hbebb3944, 32'hbd5f0024} /* (26, 23, 11) {real, imag} */,
  {32'hbe5000e1, 32'hbe41fcca} /* (26, 23, 10) {real, imag} */,
  {32'hbe2a95a7, 32'hbf1e7c0c} /* (26, 23, 9) {real, imag} */,
  {32'h3d4043ca, 32'h3e37dd09} /* (26, 23, 8) {real, imag} */,
  {32'h3d8853bc, 32'hbd889768} /* (26, 23, 7) {real, imag} */,
  {32'hbe233e48, 32'h3ebf418b} /* (26, 23, 6) {real, imag} */,
  {32'h3e3887cc, 32'hbdedfe79} /* (26, 23, 5) {real, imag} */,
  {32'hbec2b5a2, 32'h3e0fe7a8} /* (26, 23, 4) {real, imag} */,
  {32'h3ea7ad28, 32'h3de0f3ba} /* (26, 23, 3) {real, imag} */,
  {32'hbd7d1028, 32'hbf4dfbde} /* (26, 23, 2) {real, imag} */,
  {32'hbe64b64f, 32'hbf64d6a6} /* (26, 23, 1) {real, imag} */,
  {32'h3dbe6910, 32'hbee234a0} /* (26, 23, 0) {real, imag} */,
  {32'h3d737ea0, 32'hbe30a3f2} /* (26, 22, 31) {real, imag} */,
  {32'hbf11351a, 32'h3cb82150} /* (26, 22, 30) {real, imag} */,
  {32'hbe556b5a, 32'hbe23f062} /* (26, 22, 29) {real, imag} */,
  {32'hbe01c794, 32'hbe766728} /* (26, 22, 28) {real, imag} */,
  {32'hbcccb45c, 32'hbee67a43} /* (26, 22, 27) {real, imag} */,
  {32'h3e99c96f, 32'hbf04ff1d} /* (26, 22, 26) {real, imag} */,
  {32'h3f120d6b, 32'hbc9a1684} /* (26, 22, 25) {real, imag} */,
  {32'h3f09e765, 32'hbdf944a6} /* (26, 22, 24) {real, imag} */,
  {32'hbef351c7, 32'h3ed43188} /* (26, 22, 23) {real, imag} */,
  {32'hbed0e269, 32'hbd7f0b48} /* (26, 22, 22) {real, imag} */,
  {32'hbdc76a06, 32'hbed38315} /* (26, 22, 21) {real, imag} */,
  {32'hbe166510, 32'hbe74c794} /* (26, 22, 20) {real, imag} */,
  {32'hbd367f98, 32'h3f31b2a9} /* (26, 22, 19) {real, imag} */,
  {32'h3f60c595, 32'hbe312660} /* (26, 22, 18) {real, imag} */,
  {32'hbcb34160, 32'h3d25b0a4} /* (26, 22, 17) {real, imag} */,
  {32'h3e96159a, 32'hbdb56529} /* (26, 22, 16) {real, imag} */,
  {32'h3e8358ba, 32'h3c95447a} /* (26, 22, 15) {real, imag} */,
  {32'hbd47d13e, 32'hbe1ceebe} /* (26, 22, 14) {real, imag} */,
  {32'h3ef0d5be, 32'hbe9826d9} /* (26, 22, 13) {real, imag} */,
  {32'hbe9c7097, 32'hbd664184} /* (26, 22, 12) {real, imag} */,
  {32'h3e7a354a, 32'h3e973496} /* (26, 22, 11) {real, imag} */,
  {32'h3f13a47a, 32'h3ed3c15d} /* (26, 22, 10) {real, imag} */,
  {32'hbe1d1f16, 32'hbf76c6fc} /* (26, 22, 9) {real, imag} */,
  {32'hbecd5566, 32'h3e835672} /* (26, 22, 8) {real, imag} */,
  {32'hbe898e7b, 32'h3e64c5fb} /* (26, 22, 7) {real, imag} */,
  {32'hbf07f7a3, 32'h3e5a04f0} /* (26, 22, 6) {real, imag} */,
  {32'h3e6af63f, 32'h3e3891b7} /* (26, 22, 5) {real, imag} */,
  {32'hbe522fe0, 32'hbdb79ad2} /* (26, 22, 4) {real, imag} */,
  {32'h3d88df6e, 32'hbeb13864} /* (26, 22, 3) {real, imag} */,
  {32'h3eb66c73, 32'hbcb79950} /* (26, 22, 2) {real, imag} */,
  {32'hbe6b6042, 32'hbe955927} /* (26, 22, 1) {real, imag} */,
  {32'h3e714cac, 32'hbe59a308} /* (26, 22, 0) {real, imag} */,
  {32'hbe293c00, 32'hbe81dd33} /* (26, 21, 31) {real, imag} */,
  {32'h3e3cddbe, 32'hbd2d04f8} /* (26, 21, 30) {real, imag} */,
  {32'hbf324d69, 32'hbe1889c9} /* (26, 21, 29) {real, imag} */,
  {32'hbdd944df, 32'hbf307906} /* (26, 21, 28) {real, imag} */,
  {32'h3d7f6f32, 32'h3ef98328} /* (26, 21, 27) {real, imag} */,
  {32'hbd927096, 32'hbe6d5f42} /* (26, 21, 26) {real, imag} */,
  {32'hbeba0d38, 32'hbc84f020} /* (26, 21, 25) {real, imag} */,
  {32'hbebe31cf, 32'hbe9df5b9} /* (26, 21, 24) {real, imag} */,
  {32'h3e24d760, 32'hbe0b940b} /* (26, 21, 23) {real, imag} */,
  {32'hbeda5cca, 32'hbd539c68} /* (26, 21, 22) {real, imag} */,
  {32'hbd79c260, 32'hbf1a1442} /* (26, 21, 21) {real, imag} */,
  {32'h3e84884c, 32'h3e895928} /* (26, 21, 20) {real, imag} */,
  {32'hbf1d9f5a, 32'hbe8dd217} /* (26, 21, 19) {real, imag} */,
  {32'h3e92566b, 32'hbcc887d4} /* (26, 21, 18) {real, imag} */,
  {32'h3e1a359a, 32'h3e8ef6a6} /* (26, 21, 17) {real, imag} */,
  {32'h3c3cc8d8, 32'h3ed125d2} /* (26, 21, 16) {real, imag} */,
  {32'h3eae67c8, 32'hbee7d40b} /* (26, 21, 15) {real, imag} */,
  {32'hbf23239a, 32'h3eee5c2d} /* (26, 21, 14) {real, imag} */,
  {32'h3e2af216, 32'h3d887f90} /* (26, 21, 13) {real, imag} */,
  {32'hbec735f2, 32'h3f0ff434} /* (26, 21, 12) {real, imag} */,
  {32'hbd97cdd8, 32'h3e4f0da7} /* (26, 21, 11) {real, imag} */,
  {32'hbee118dc, 32'h3e4fce8c} /* (26, 21, 10) {real, imag} */,
  {32'h3da963d4, 32'hbe205b54} /* (26, 21, 9) {real, imag} */,
  {32'hbec5db78, 32'h3d6c2614} /* (26, 21, 8) {real, imag} */,
  {32'h3e941c1c, 32'hbdd02d52} /* (26, 21, 7) {real, imag} */,
  {32'hbedadd87, 32'h3f567cd0} /* (26, 21, 6) {real, imag} */,
  {32'hbed59f8f, 32'h3e363809} /* (26, 21, 5) {real, imag} */,
  {32'hbd1cd748, 32'hbed94964} /* (26, 21, 4) {real, imag} */,
  {32'h3ebe9fb4, 32'h3e2824ca} /* (26, 21, 3) {real, imag} */,
  {32'h3d9b8fa9, 32'hbd470910} /* (26, 21, 2) {real, imag} */,
  {32'hbe7dd766, 32'h3ef97d7f} /* (26, 21, 1) {real, imag} */,
  {32'hbf1cf981, 32'h3ee8ead4} /* (26, 21, 0) {real, imag} */,
  {32'hbdb005fa, 32'hbde7c8e0} /* (26, 20, 31) {real, imag} */,
  {32'h3d233438, 32'hbe1f0cc6} /* (26, 20, 30) {real, imag} */,
  {32'h3d84af28, 32'hbf0577a6} /* (26, 20, 29) {real, imag} */,
  {32'hbdeb1312, 32'hbd2efb1e} /* (26, 20, 28) {real, imag} */,
  {32'h3d71b10e, 32'hbd579170} /* (26, 20, 27) {real, imag} */,
  {32'hbf1193ea, 32'hbe772b32} /* (26, 20, 26) {real, imag} */,
  {32'h3e9cf298, 32'hbe708f68} /* (26, 20, 25) {real, imag} */,
  {32'h3d9b7768, 32'h3d55a208} /* (26, 20, 24) {real, imag} */,
  {32'hbefe8487, 32'h3ef087a2} /* (26, 20, 23) {real, imag} */,
  {32'hbe095ed2, 32'hbe276729} /* (26, 20, 22) {real, imag} */,
  {32'h3e1e5f59, 32'hbde5074e} /* (26, 20, 21) {real, imag} */,
  {32'hbcff40ca, 32'h3e3d7112} /* (26, 20, 20) {real, imag} */,
  {32'h3e0877b3, 32'h3e1ada38} /* (26, 20, 19) {real, imag} */,
  {32'h3e81f634, 32'hbda2d0bf} /* (26, 20, 18) {real, imag} */,
  {32'hbdc3800c, 32'hbe8c50be} /* (26, 20, 17) {real, imag} */,
  {32'hbdae036a, 32'h3ecca1e7} /* (26, 20, 16) {real, imag} */,
  {32'hbf220a3a, 32'hbec6b939} /* (26, 20, 15) {real, imag} */,
  {32'h3df0a5ea, 32'hbdd9479d} /* (26, 20, 14) {real, imag} */,
  {32'h3e475e6c, 32'hbef52ca6} /* (26, 20, 13) {real, imag} */,
  {32'hbdd8794e, 32'hbd68e140} /* (26, 20, 12) {real, imag} */,
  {32'hbece872e, 32'hbdfd3d3c} /* (26, 20, 11) {real, imag} */,
  {32'h3bbc67a0, 32'h3e230ca4} /* (26, 20, 10) {real, imag} */,
  {32'h3e152f68, 32'h3f360888} /* (26, 20, 9) {real, imag} */,
  {32'hbf11d211, 32'h3e6dda89} /* (26, 20, 8) {real, imag} */,
  {32'hbe7a6148, 32'hbf1210ca} /* (26, 20, 7) {real, imag} */,
  {32'h3d926fce, 32'h3e8fd298} /* (26, 20, 6) {real, imag} */,
  {32'hbd371670, 32'hbdbe3716} /* (26, 20, 5) {real, imag} */,
  {32'hbe2a7129, 32'hbe724096} /* (26, 20, 4) {real, imag} */,
  {32'h3e2e339e, 32'h3ebb52aa} /* (26, 20, 3) {real, imag} */,
  {32'hbccc53d0, 32'hbebfb70e} /* (26, 20, 2) {real, imag} */,
  {32'hbd055e90, 32'hbeb91d7f} /* (26, 20, 1) {real, imag} */,
  {32'h3f2336c3, 32'h3f636d4a} /* (26, 20, 0) {real, imag} */,
  {32'hbd85bd0e, 32'hbdf0c2a4} /* (26, 19, 31) {real, imag} */,
  {32'hbdd83bba, 32'hbe880ca9} /* (26, 19, 30) {real, imag} */,
  {32'h3ec9ae4b, 32'hbd817432} /* (26, 19, 29) {real, imag} */,
  {32'hbe9a84e1, 32'hbef5018c} /* (26, 19, 28) {real, imag} */,
  {32'hbcc51770, 32'h3eaa72f2} /* (26, 19, 27) {real, imag} */,
  {32'hbeda23b0, 32'h3e7d65ea} /* (26, 19, 26) {real, imag} */,
  {32'h3e9c2a31, 32'h3e1e92d8} /* (26, 19, 25) {real, imag} */,
  {32'h3ed1ef5d, 32'h3dd1f536} /* (26, 19, 24) {real, imag} */,
  {32'hbe811c5f, 32'h3c09d5a0} /* (26, 19, 23) {real, imag} */,
  {32'h3eb709d4, 32'hbd65ffb2} /* (26, 19, 22) {real, imag} */,
  {32'h3e83ad80, 32'hbeb0b11e} /* (26, 19, 21) {real, imag} */,
  {32'hbe9a8176, 32'hbd7a4ec8} /* (26, 19, 20) {real, imag} */,
  {32'hbee5feea, 32'h3ef95524} /* (26, 19, 19) {real, imag} */,
  {32'h3e644d9e, 32'h3ea800a5} /* (26, 19, 18) {real, imag} */,
  {32'h3e1383ec, 32'hbda863d4} /* (26, 19, 17) {real, imag} */,
  {32'h3dabd8ba, 32'h3da58bcd} /* (26, 19, 16) {real, imag} */,
  {32'hbed1fb1a, 32'hbd9413d5} /* (26, 19, 15) {real, imag} */,
  {32'hbe396370, 32'hbda7344d} /* (26, 19, 14) {real, imag} */,
  {32'hbe4f78b8, 32'hbe88d67c} /* (26, 19, 13) {real, imag} */,
  {32'hbd6076a0, 32'hbf073aac} /* (26, 19, 12) {real, imag} */,
  {32'hbc69a530, 32'hbe0256db} /* (26, 19, 11) {real, imag} */,
  {32'h3eb01879, 32'hbf13a284} /* (26, 19, 10) {real, imag} */,
  {32'h3df93d04, 32'h3c175860} /* (26, 19, 9) {real, imag} */,
  {32'h3dfb26fb, 32'h3f157fb6} /* (26, 19, 8) {real, imag} */,
  {32'h3e82169a, 32'hbe2c4182} /* (26, 19, 7) {real, imag} */,
  {32'h3ec9183e, 32'h3d3ecd1e} /* (26, 19, 6) {real, imag} */,
  {32'hbde81048, 32'hbeaa3c4f} /* (26, 19, 5) {real, imag} */,
  {32'h3e4a08f7, 32'hbe7b802c} /* (26, 19, 4) {real, imag} */,
  {32'hbbd07aa0, 32'h3d1f8452} /* (26, 19, 3) {real, imag} */,
  {32'h3e23a817, 32'h3d8f4338} /* (26, 19, 2) {real, imag} */,
  {32'h3d7efd8c, 32'h3ee5a5f2} /* (26, 19, 1) {real, imag} */,
  {32'hbdc69110, 32'hbe1656f6} /* (26, 19, 0) {real, imag} */,
  {32'hbec3cb49, 32'hbddac8d6} /* (26, 18, 31) {real, imag} */,
  {32'h3e4a0ec2, 32'h3f13cfbe} /* (26, 18, 30) {real, imag} */,
  {32'h3eb1eb71, 32'hbec72c37} /* (26, 18, 29) {real, imag} */,
  {32'hbeab4235, 32'hbe5a2794} /* (26, 18, 28) {real, imag} */,
  {32'h3e442bb2, 32'h3eb6e976} /* (26, 18, 27) {real, imag} */,
  {32'hbead0114, 32'hbde7e7ec} /* (26, 18, 26) {real, imag} */,
  {32'hbe8f1161, 32'h3ea72c00} /* (26, 18, 25) {real, imag} */,
  {32'hbdc208fd, 32'hbe072640} /* (26, 18, 24) {real, imag} */,
  {32'h3e0ef6a6, 32'hbe600c2a} /* (26, 18, 23) {real, imag} */,
  {32'hbce53800, 32'h3ee97c82} /* (26, 18, 22) {real, imag} */,
  {32'hbd91098c, 32'h3ec74949} /* (26, 18, 21) {real, imag} */,
  {32'hbed580c5, 32'h3e7173b4} /* (26, 18, 20) {real, imag} */,
  {32'h3e465278, 32'hbe1704b2} /* (26, 18, 19) {real, imag} */,
  {32'hbe28d713, 32'h3f082daa} /* (26, 18, 18) {real, imag} */,
  {32'hbea8db21, 32'hbe015976} /* (26, 18, 17) {real, imag} */,
  {32'h3e18af1f, 32'h3e471ac2} /* (26, 18, 16) {real, imag} */,
  {32'h3ef145d2, 32'h3ef22df8} /* (26, 18, 15) {real, imag} */,
  {32'hbe4c740e, 32'hbdc78f79} /* (26, 18, 14) {real, imag} */,
  {32'h3d6b9ff0, 32'h3df2dc74} /* (26, 18, 13) {real, imag} */,
  {32'h3e6a8b87, 32'h3d47c508} /* (26, 18, 12) {real, imag} */,
  {32'h3ee06ae2, 32'h3dcc6106} /* (26, 18, 11) {real, imag} */,
  {32'h3e53dd1c, 32'hbdf2ef80} /* (26, 18, 10) {real, imag} */,
  {32'h3e86b58a, 32'hbdeba05c} /* (26, 18, 9) {real, imag} */,
  {32'hbde7cada, 32'hbe926c1b} /* (26, 18, 8) {real, imag} */,
  {32'h3df82f88, 32'hbe3569c8} /* (26, 18, 7) {real, imag} */,
  {32'h3e8ed0be, 32'hbc7c9568} /* (26, 18, 6) {real, imag} */,
  {32'hbe365743, 32'h3e060ad2} /* (26, 18, 5) {real, imag} */,
  {32'hbe8b1bf2, 32'h3e835dad} /* (26, 18, 4) {real, imag} */,
  {32'h3e8ac57c, 32'h3dd02ac0} /* (26, 18, 3) {real, imag} */,
  {32'h3edd557a, 32'hbe5d732d} /* (26, 18, 2) {real, imag} */,
  {32'hbe3f0f6c, 32'h3e00fe24} /* (26, 18, 1) {real, imag} */,
  {32'h3e74d8d0, 32'hbee3b734} /* (26, 18, 0) {real, imag} */,
  {32'hbddec7e8, 32'hbd8d8f37} /* (26, 17, 31) {real, imag} */,
  {32'hbd37c612, 32'hbca82a30} /* (26, 17, 30) {real, imag} */,
  {32'h3e31db82, 32'h3e13d620} /* (26, 17, 29) {real, imag} */,
  {32'hbe111d3e, 32'h3b51ad00} /* (26, 17, 28) {real, imag} */,
  {32'h3ea37628, 32'hbe64be64} /* (26, 17, 27) {real, imag} */,
  {32'hbc243bd4, 32'hbeda4351} /* (26, 17, 26) {real, imag} */,
  {32'h3e373414, 32'hbd359324} /* (26, 17, 25) {real, imag} */,
  {32'hbe956468, 32'h3e1e94a9} /* (26, 17, 24) {real, imag} */,
  {32'hbe17db80, 32'h3d86d8fa} /* (26, 17, 23) {real, imag} */,
  {32'hbea37d38, 32'hbefaee83} /* (26, 17, 22) {real, imag} */,
  {32'h3e6ab226, 32'h3effba3a} /* (26, 17, 21) {real, imag} */,
  {32'hbea396bc, 32'hbe084e6a} /* (26, 17, 20) {real, imag} */,
  {32'hbd150dae, 32'h3dc38a91} /* (26, 17, 19) {real, imag} */,
  {32'hbcbc803c, 32'hbec1f766} /* (26, 17, 18) {real, imag} */,
  {32'hbe620a90, 32'hbe6d94f8} /* (26, 17, 17) {real, imag} */,
  {32'h3e0f8928, 32'h3c7af228} /* (26, 17, 16) {real, imag} */,
  {32'h3e9716d6, 32'h3dded3e0} /* (26, 17, 15) {real, imag} */,
  {32'h3d20c60a, 32'h3e8fc3c4} /* (26, 17, 14) {real, imag} */,
  {32'hbeb79f5a, 32'hbe0cf49a} /* (26, 17, 13) {real, imag} */,
  {32'h3e5626b0, 32'hbc0d8ec8} /* (26, 17, 12) {real, imag} */,
  {32'h3e0fc810, 32'h3e2fdcae} /* (26, 17, 11) {real, imag} */,
  {32'hbb107780, 32'hbef743cf} /* (26, 17, 10) {real, imag} */,
  {32'hbe4090db, 32'h3e9c79b2} /* (26, 17, 9) {real, imag} */,
  {32'hbe3daafa, 32'hbe708194} /* (26, 17, 8) {real, imag} */,
  {32'hbd9ed18a, 32'h3d805a88} /* (26, 17, 7) {real, imag} */,
  {32'h3e8c5cf3, 32'hbe603ef3} /* (26, 17, 6) {real, imag} */,
  {32'hbe8133ac, 32'h3d0fbfe0} /* (26, 17, 5) {real, imag} */,
  {32'h3e4f4178, 32'h3eb98e5c} /* (26, 17, 4) {real, imag} */,
  {32'hbe0abd77, 32'hb9210300} /* (26, 17, 3) {real, imag} */,
  {32'hbe37f41a, 32'hbe02a19f} /* (26, 17, 2) {real, imag} */,
  {32'hbee18874, 32'h3e9424c0} /* (26, 17, 1) {real, imag} */,
  {32'hbdf39cd6, 32'hbd0a1d90} /* (26, 17, 0) {real, imag} */,
  {32'h3d2f9696, 32'hbe762ab7} /* (26, 16, 31) {real, imag} */,
  {32'h3e22568c, 32'hbdf3ffa2} /* (26, 16, 30) {real, imag} */,
  {32'h3b2718a0, 32'hbe49c2d9} /* (26, 16, 29) {real, imag} */,
  {32'h3db3067c, 32'hbe50a902} /* (26, 16, 28) {real, imag} */,
  {32'hbe29a95c, 32'hbe7ce2b2} /* (26, 16, 27) {real, imag} */,
  {32'hbe68ac0c, 32'hbc33d5ee} /* (26, 16, 26) {real, imag} */,
  {32'hbd49f16e, 32'hbd39f718} /* (26, 16, 25) {real, imag} */,
  {32'hbe62eb82, 32'h3e948576} /* (26, 16, 24) {real, imag} */,
  {32'h3e7b631d, 32'h3c9f1e38} /* (26, 16, 23) {real, imag} */,
  {32'h3cfcf498, 32'hbda3e0ac} /* (26, 16, 22) {real, imag} */,
  {32'h3e635c66, 32'hbd584a12} /* (26, 16, 21) {real, imag} */,
  {32'hbe4c3f01, 32'hbe87aa71} /* (26, 16, 20) {real, imag} */,
  {32'hbb9ac210, 32'h3e45c16c} /* (26, 16, 19) {real, imag} */,
  {32'h3d9bbbd6, 32'hbea46c62} /* (26, 16, 18) {real, imag} */,
  {32'h3e5a3487, 32'hbdcd0cea} /* (26, 16, 17) {real, imag} */,
  {32'h3c96db44, 32'h00000000} /* (26, 16, 16) {real, imag} */,
  {32'h3e5a3487, 32'h3dcd0cea} /* (26, 16, 15) {real, imag} */,
  {32'h3d9bbbd6, 32'h3ea46c62} /* (26, 16, 14) {real, imag} */,
  {32'hbb9ac210, 32'hbe45c16c} /* (26, 16, 13) {real, imag} */,
  {32'hbe4c3f01, 32'h3e87aa71} /* (26, 16, 12) {real, imag} */,
  {32'h3e635c66, 32'h3d584a12} /* (26, 16, 11) {real, imag} */,
  {32'h3cfcf498, 32'h3da3e0ac} /* (26, 16, 10) {real, imag} */,
  {32'h3e7b631d, 32'hbc9f1e38} /* (26, 16, 9) {real, imag} */,
  {32'hbe62eb82, 32'hbe948576} /* (26, 16, 8) {real, imag} */,
  {32'hbd49f16e, 32'h3d39f718} /* (26, 16, 7) {real, imag} */,
  {32'hbe68ac0c, 32'h3c33d5ee} /* (26, 16, 6) {real, imag} */,
  {32'hbe29a95c, 32'h3e7ce2b2} /* (26, 16, 5) {real, imag} */,
  {32'h3db3067c, 32'h3e50a902} /* (26, 16, 4) {real, imag} */,
  {32'h3b2718a0, 32'h3e49c2d9} /* (26, 16, 3) {real, imag} */,
  {32'h3e22568c, 32'h3df3ffa2} /* (26, 16, 2) {real, imag} */,
  {32'h3d2f9696, 32'h3e762ab7} /* (26, 16, 1) {real, imag} */,
  {32'h3e3dbece, 32'h00000000} /* (26, 16, 0) {real, imag} */,
  {32'hbee18874, 32'hbe9424c0} /* (26, 15, 31) {real, imag} */,
  {32'hbe37f41a, 32'h3e02a19f} /* (26, 15, 30) {real, imag} */,
  {32'hbe0abd77, 32'h39210300} /* (26, 15, 29) {real, imag} */,
  {32'h3e4f4178, 32'hbeb98e5c} /* (26, 15, 28) {real, imag} */,
  {32'hbe8133ac, 32'hbd0fbfe0} /* (26, 15, 27) {real, imag} */,
  {32'h3e8c5cf3, 32'h3e603ef3} /* (26, 15, 26) {real, imag} */,
  {32'hbd9ed18a, 32'hbd805a88} /* (26, 15, 25) {real, imag} */,
  {32'hbe3daafa, 32'h3e708194} /* (26, 15, 24) {real, imag} */,
  {32'hbe4090db, 32'hbe9c79b2} /* (26, 15, 23) {real, imag} */,
  {32'hbb107780, 32'h3ef743cf} /* (26, 15, 22) {real, imag} */,
  {32'h3e0fc810, 32'hbe2fdcae} /* (26, 15, 21) {real, imag} */,
  {32'h3e5626b0, 32'h3c0d8ec8} /* (26, 15, 20) {real, imag} */,
  {32'hbeb79f5a, 32'h3e0cf49a} /* (26, 15, 19) {real, imag} */,
  {32'h3d20c60a, 32'hbe8fc3c4} /* (26, 15, 18) {real, imag} */,
  {32'h3e9716d6, 32'hbdded3e0} /* (26, 15, 17) {real, imag} */,
  {32'h3e0f8928, 32'hbc7af228} /* (26, 15, 16) {real, imag} */,
  {32'hbe620a90, 32'h3e6d94f8} /* (26, 15, 15) {real, imag} */,
  {32'hbcbc803c, 32'h3ec1f766} /* (26, 15, 14) {real, imag} */,
  {32'hbd150dae, 32'hbdc38a91} /* (26, 15, 13) {real, imag} */,
  {32'hbea396bc, 32'h3e084e6a} /* (26, 15, 12) {real, imag} */,
  {32'h3e6ab226, 32'hbeffba3a} /* (26, 15, 11) {real, imag} */,
  {32'hbea37d38, 32'h3efaee83} /* (26, 15, 10) {real, imag} */,
  {32'hbe17db80, 32'hbd86d8fa} /* (26, 15, 9) {real, imag} */,
  {32'hbe956468, 32'hbe1e94a9} /* (26, 15, 8) {real, imag} */,
  {32'h3e373414, 32'h3d359324} /* (26, 15, 7) {real, imag} */,
  {32'hbc243bd4, 32'h3eda4351} /* (26, 15, 6) {real, imag} */,
  {32'h3ea37628, 32'h3e64be64} /* (26, 15, 5) {real, imag} */,
  {32'hbe111d3e, 32'hbb51ad00} /* (26, 15, 4) {real, imag} */,
  {32'h3e31db82, 32'hbe13d620} /* (26, 15, 3) {real, imag} */,
  {32'hbd37c612, 32'h3ca82a30} /* (26, 15, 2) {real, imag} */,
  {32'hbddec7e8, 32'h3d8d8f37} /* (26, 15, 1) {real, imag} */,
  {32'hbdf39cd6, 32'h3d0a1d90} /* (26, 15, 0) {real, imag} */,
  {32'hbe3f0f6c, 32'hbe00fe24} /* (26, 14, 31) {real, imag} */,
  {32'h3edd557a, 32'h3e5d732d} /* (26, 14, 30) {real, imag} */,
  {32'h3e8ac57c, 32'hbdd02ac0} /* (26, 14, 29) {real, imag} */,
  {32'hbe8b1bf2, 32'hbe835dad} /* (26, 14, 28) {real, imag} */,
  {32'hbe365743, 32'hbe060ad2} /* (26, 14, 27) {real, imag} */,
  {32'h3e8ed0be, 32'h3c7c9568} /* (26, 14, 26) {real, imag} */,
  {32'h3df82f88, 32'h3e3569c8} /* (26, 14, 25) {real, imag} */,
  {32'hbde7cada, 32'h3e926c1b} /* (26, 14, 24) {real, imag} */,
  {32'h3e86b58a, 32'h3deba05c} /* (26, 14, 23) {real, imag} */,
  {32'h3e53dd1c, 32'h3df2ef80} /* (26, 14, 22) {real, imag} */,
  {32'h3ee06ae2, 32'hbdcc6106} /* (26, 14, 21) {real, imag} */,
  {32'h3e6a8b87, 32'hbd47c508} /* (26, 14, 20) {real, imag} */,
  {32'h3d6b9ff0, 32'hbdf2dc74} /* (26, 14, 19) {real, imag} */,
  {32'hbe4c740e, 32'h3dc78f79} /* (26, 14, 18) {real, imag} */,
  {32'h3ef145d2, 32'hbef22df8} /* (26, 14, 17) {real, imag} */,
  {32'h3e18af1f, 32'hbe471ac2} /* (26, 14, 16) {real, imag} */,
  {32'hbea8db21, 32'h3e015976} /* (26, 14, 15) {real, imag} */,
  {32'hbe28d713, 32'hbf082daa} /* (26, 14, 14) {real, imag} */,
  {32'h3e465278, 32'h3e1704b2} /* (26, 14, 13) {real, imag} */,
  {32'hbed580c5, 32'hbe7173b4} /* (26, 14, 12) {real, imag} */,
  {32'hbd91098c, 32'hbec74949} /* (26, 14, 11) {real, imag} */,
  {32'hbce53800, 32'hbee97c82} /* (26, 14, 10) {real, imag} */,
  {32'h3e0ef6a6, 32'h3e600c2a} /* (26, 14, 9) {real, imag} */,
  {32'hbdc208fd, 32'h3e072640} /* (26, 14, 8) {real, imag} */,
  {32'hbe8f1161, 32'hbea72c00} /* (26, 14, 7) {real, imag} */,
  {32'hbead0114, 32'h3de7e7ec} /* (26, 14, 6) {real, imag} */,
  {32'h3e442bb2, 32'hbeb6e976} /* (26, 14, 5) {real, imag} */,
  {32'hbeab4235, 32'h3e5a2794} /* (26, 14, 4) {real, imag} */,
  {32'h3eb1eb71, 32'h3ec72c37} /* (26, 14, 3) {real, imag} */,
  {32'h3e4a0ec2, 32'hbf13cfbe} /* (26, 14, 2) {real, imag} */,
  {32'hbec3cb49, 32'h3ddac8d6} /* (26, 14, 1) {real, imag} */,
  {32'h3e74d8d0, 32'h3ee3b734} /* (26, 14, 0) {real, imag} */,
  {32'h3d7efd8c, 32'hbee5a5f2} /* (26, 13, 31) {real, imag} */,
  {32'h3e23a817, 32'hbd8f4338} /* (26, 13, 30) {real, imag} */,
  {32'hbbd07aa0, 32'hbd1f8452} /* (26, 13, 29) {real, imag} */,
  {32'h3e4a08f7, 32'h3e7b802c} /* (26, 13, 28) {real, imag} */,
  {32'hbde81048, 32'h3eaa3c4f} /* (26, 13, 27) {real, imag} */,
  {32'h3ec9183e, 32'hbd3ecd1e} /* (26, 13, 26) {real, imag} */,
  {32'h3e82169a, 32'h3e2c4182} /* (26, 13, 25) {real, imag} */,
  {32'h3dfb26fb, 32'hbf157fb6} /* (26, 13, 24) {real, imag} */,
  {32'h3df93d04, 32'hbc175860} /* (26, 13, 23) {real, imag} */,
  {32'h3eb01879, 32'h3f13a284} /* (26, 13, 22) {real, imag} */,
  {32'hbc69a530, 32'h3e0256db} /* (26, 13, 21) {real, imag} */,
  {32'hbd6076a0, 32'h3f073aac} /* (26, 13, 20) {real, imag} */,
  {32'hbe4f78b8, 32'h3e88d67c} /* (26, 13, 19) {real, imag} */,
  {32'hbe396370, 32'h3da7344d} /* (26, 13, 18) {real, imag} */,
  {32'hbed1fb1a, 32'h3d9413d5} /* (26, 13, 17) {real, imag} */,
  {32'h3dabd8ba, 32'hbda58bcd} /* (26, 13, 16) {real, imag} */,
  {32'h3e1383ec, 32'h3da863d4} /* (26, 13, 15) {real, imag} */,
  {32'h3e644d9e, 32'hbea800a5} /* (26, 13, 14) {real, imag} */,
  {32'hbee5feea, 32'hbef95524} /* (26, 13, 13) {real, imag} */,
  {32'hbe9a8176, 32'h3d7a4ec8} /* (26, 13, 12) {real, imag} */,
  {32'h3e83ad80, 32'h3eb0b11e} /* (26, 13, 11) {real, imag} */,
  {32'h3eb709d4, 32'h3d65ffb2} /* (26, 13, 10) {real, imag} */,
  {32'hbe811c5f, 32'hbc09d5a0} /* (26, 13, 9) {real, imag} */,
  {32'h3ed1ef5d, 32'hbdd1f536} /* (26, 13, 8) {real, imag} */,
  {32'h3e9c2a31, 32'hbe1e92d8} /* (26, 13, 7) {real, imag} */,
  {32'hbeda23b0, 32'hbe7d65ea} /* (26, 13, 6) {real, imag} */,
  {32'hbcc51770, 32'hbeaa72f2} /* (26, 13, 5) {real, imag} */,
  {32'hbe9a84e1, 32'h3ef5018c} /* (26, 13, 4) {real, imag} */,
  {32'h3ec9ae4b, 32'h3d817432} /* (26, 13, 3) {real, imag} */,
  {32'hbdd83bba, 32'h3e880ca9} /* (26, 13, 2) {real, imag} */,
  {32'hbd85bd0e, 32'h3df0c2a4} /* (26, 13, 1) {real, imag} */,
  {32'hbdc69110, 32'h3e1656f6} /* (26, 13, 0) {real, imag} */,
  {32'hbd055e90, 32'h3eb91d7f} /* (26, 12, 31) {real, imag} */,
  {32'hbccc53d0, 32'h3ebfb70e} /* (26, 12, 30) {real, imag} */,
  {32'h3e2e339e, 32'hbebb52aa} /* (26, 12, 29) {real, imag} */,
  {32'hbe2a7129, 32'h3e724096} /* (26, 12, 28) {real, imag} */,
  {32'hbd371670, 32'h3dbe3716} /* (26, 12, 27) {real, imag} */,
  {32'h3d926fce, 32'hbe8fd298} /* (26, 12, 26) {real, imag} */,
  {32'hbe7a6148, 32'h3f1210ca} /* (26, 12, 25) {real, imag} */,
  {32'hbf11d211, 32'hbe6dda89} /* (26, 12, 24) {real, imag} */,
  {32'h3e152f68, 32'hbf360888} /* (26, 12, 23) {real, imag} */,
  {32'h3bbc67a0, 32'hbe230ca4} /* (26, 12, 22) {real, imag} */,
  {32'hbece872e, 32'h3dfd3d3c} /* (26, 12, 21) {real, imag} */,
  {32'hbdd8794e, 32'h3d68e140} /* (26, 12, 20) {real, imag} */,
  {32'h3e475e6c, 32'h3ef52ca6} /* (26, 12, 19) {real, imag} */,
  {32'h3df0a5ea, 32'h3dd9479d} /* (26, 12, 18) {real, imag} */,
  {32'hbf220a3a, 32'h3ec6b939} /* (26, 12, 17) {real, imag} */,
  {32'hbdae036a, 32'hbecca1e7} /* (26, 12, 16) {real, imag} */,
  {32'hbdc3800c, 32'h3e8c50be} /* (26, 12, 15) {real, imag} */,
  {32'h3e81f634, 32'h3da2d0bf} /* (26, 12, 14) {real, imag} */,
  {32'h3e0877b3, 32'hbe1ada38} /* (26, 12, 13) {real, imag} */,
  {32'hbcff40ca, 32'hbe3d7112} /* (26, 12, 12) {real, imag} */,
  {32'h3e1e5f59, 32'h3de5074e} /* (26, 12, 11) {real, imag} */,
  {32'hbe095ed2, 32'h3e276729} /* (26, 12, 10) {real, imag} */,
  {32'hbefe8487, 32'hbef087a2} /* (26, 12, 9) {real, imag} */,
  {32'h3d9b7768, 32'hbd55a208} /* (26, 12, 8) {real, imag} */,
  {32'h3e9cf298, 32'h3e708f68} /* (26, 12, 7) {real, imag} */,
  {32'hbf1193ea, 32'h3e772b32} /* (26, 12, 6) {real, imag} */,
  {32'h3d71b10e, 32'h3d579170} /* (26, 12, 5) {real, imag} */,
  {32'hbdeb1312, 32'h3d2efb1e} /* (26, 12, 4) {real, imag} */,
  {32'h3d84af28, 32'h3f0577a6} /* (26, 12, 3) {real, imag} */,
  {32'h3d233438, 32'h3e1f0cc6} /* (26, 12, 2) {real, imag} */,
  {32'hbdb005fa, 32'h3de7c8e0} /* (26, 12, 1) {real, imag} */,
  {32'h3f2336c3, 32'hbf636d4a} /* (26, 12, 0) {real, imag} */,
  {32'hbe7dd766, 32'hbef97d7f} /* (26, 11, 31) {real, imag} */,
  {32'h3d9b8fa9, 32'h3d470910} /* (26, 11, 30) {real, imag} */,
  {32'h3ebe9fb4, 32'hbe2824ca} /* (26, 11, 29) {real, imag} */,
  {32'hbd1cd748, 32'h3ed94964} /* (26, 11, 28) {real, imag} */,
  {32'hbed59f8f, 32'hbe363809} /* (26, 11, 27) {real, imag} */,
  {32'hbedadd87, 32'hbf567cd0} /* (26, 11, 26) {real, imag} */,
  {32'h3e941c1c, 32'h3dd02d52} /* (26, 11, 25) {real, imag} */,
  {32'hbec5db78, 32'hbd6c2614} /* (26, 11, 24) {real, imag} */,
  {32'h3da963d4, 32'h3e205b54} /* (26, 11, 23) {real, imag} */,
  {32'hbee118dc, 32'hbe4fce8c} /* (26, 11, 22) {real, imag} */,
  {32'hbd97cdd8, 32'hbe4f0da7} /* (26, 11, 21) {real, imag} */,
  {32'hbec735f2, 32'hbf0ff434} /* (26, 11, 20) {real, imag} */,
  {32'h3e2af216, 32'hbd887f90} /* (26, 11, 19) {real, imag} */,
  {32'hbf23239a, 32'hbeee5c2d} /* (26, 11, 18) {real, imag} */,
  {32'h3eae67c8, 32'h3ee7d40b} /* (26, 11, 17) {real, imag} */,
  {32'h3c3cc8d8, 32'hbed125d2} /* (26, 11, 16) {real, imag} */,
  {32'h3e1a359a, 32'hbe8ef6a6} /* (26, 11, 15) {real, imag} */,
  {32'h3e92566b, 32'h3cc887d4} /* (26, 11, 14) {real, imag} */,
  {32'hbf1d9f5a, 32'h3e8dd217} /* (26, 11, 13) {real, imag} */,
  {32'h3e84884c, 32'hbe895928} /* (26, 11, 12) {real, imag} */,
  {32'hbd79c260, 32'h3f1a1442} /* (26, 11, 11) {real, imag} */,
  {32'hbeda5cca, 32'h3d539c68} /* (26, 11, 10) {real, imag} */,
  {32'h3e24d760, 32'h3e0b940b} /* (26, 11, 9) {real, imag} */,
  {32'hbebe31cf, 32'h3e9df5b9} /* (26, 11, 8) {real, imag} */,
  {32'hbeba0d38, 32'h3c84f020} /* (26, 11, 7) {real, imag} */,
  {32'hbd927096, 32'h3e6d5f42} /* (26, 11, 6) {real, imag} */,
  {32'h3d7f6f32, 32'hbef98328} /* (26, 11, 5) {real, imag} */,
  {32'hbdd944df, 32'h3f307906} /* (26, 11, 4) {real, imag} */,
  {32'hbf324d69, 32'h3e1889c9} /* (26, 11, 3) {real, imag} */,
  {32'h3e3cddbe, 32'h3d2d04f8} /* (26, 11, 2) {real, imag} */,
  {32'hbe293c00, 32'h3e81dd33} /* (26, 11, 1) {real, imag} */,
  {32'hbf1cf981, 32'hbee8ead4} /* (26, 11, 0) {real, imag} */,
  {32'hbe6b6042, 32'h3e955927} /* (26, 10, 31) {real, imag} */,
  {32'h3eb66c73, 32'h3cb79950} /* (26, 10, 30) {real, imag} */,
  {32'h3d88df6e, 32'h3eb13864} /* (26, 10, 29) {real, imag} */,
  {32'hbe522fe0, 32'h3db79ad2} /* (26, 10, 28) {real, imag} */,
  {32'h3e6af63f, 32'hbe3891b7} /* (26, 10, 27) {real, imag} */,
  {32'hbf07f7a3, 32'hbe5a04f0} /* (26, 10, 26) {real, imag} */,
  {32'hbe898e7b, 32'hbe64c5fb} /* (26, 10, 25) {real, imag} */,
  {32'hbecd5566, 32'hbe835672} /* (26, 10, 24) {real, imag} */,
  {32'hbe1d1f16, 32'h3f76c6fc} /* (26, 10, 23) {real, imag} */,
  {32'h3f13a47a, 32'hbed3c15d} /* (26, 10, 22) {real, imag} */,
  {32'h3e7a354a, 32'hbe973496} /* (26, 10, 21) {real, imag} */,
  {32'hbe9c7097, 32'h3d664184} /* (26, 10, 20) {real, imag} */,
  {32'h3ef0d5be, 32'h3e9826d9} /* (26, 10, 19) {real, imag} */,
  {32'hbd47d13e, 32'h3e1ceebe} /* (26, 10, 18) {real, imag} */,
  {32'h3e8358ba, 32'hbc95447a} /* (26, 10, 17) {real, imag} */,
  {32'h3e96159a, 32'h3db56529} /* (26, 10, 16) {real, imag} */,
  {32'hbcb34160, 32'hbd25b0a4} /* (26, 10, 15) {real, imag} */,
  {32'h3f60c595, 32'h3e312660} /* (26, 10, 14) {real, imag} */,
  {32'hbd367f98, 32'hbf31b2a9} /* (26, 10, 13) {real, imag} */,
  {32'hbe166510, 32'h3e74c794} /* (26, 10, 12) {real, imag} */,
  {32'hbdc76a06, 32'h3ed38315} /* (26, 10, 11) {real, imag} */,
  {32'hbed0e269, 32'h3d7f0b48} /* (26, 10, 10) {real, imag} */,
  {32'hbef351c7, 32'hbed43188} /* (26, 10, 9) {real, imag} */,
  {32'h3f09e765, 32'h3df944a6} /* (26, 10, 8) {real, imag} */,
  {32'h3f120d6b, 32'h3c9a1684} /* (26, 10, 7) {real, imag} */,
  {32'h3e99c96f, 32'h3f04ff1d} /* (26, 10, 6) {real, imag} */,
  {32'hbcccb45c, 32'h3ee67a43} /* (26, 10, 5) {real, imag} */,
  {32'hbe01c794, 32'h3e766728} /* (26, 10, 4) {real, imag} */,
  {32'hbe556b5a, 32'h3e23f062} /* (26, 10, 3) {real, imag} */,
  {32'hbf11351a, 32'hbcb82150} /* (26, 10, 2) {real, imag} */,
  {32'h3d737ea0, 32'h3e30a3f2} /* (26, 10, 1) {real, imag} */,
  {32'h3e714cac, 32'h3e59a308} /* (26, 10, 0) {real, imag} */,
  {32'hbe64b64f, 32'h3f64d6a6} /* (26, 9, 31) {real, imag} */,
  {32'hbd7d1028, 32'h3f4dfbde} /* (26, 9, 30) {real, imag} */,
  {32'h3ea7ad28, 32'hbde0f3ba} /* (26, 9, 29) {real, imag} */,
  {32'hbec2b5a2, 32'hbe0fe7a8} /* (26, 9, 28) {real, imag} */,
  {32'h3e3887cc, 32'h3dedfe79} /* (26, 9, 27) {real, imag} */,
  {32'hbe233e48, 32'hbebf418b} /* (26, 9, 26) {real, imag} */,
  {32'h3d8853bc, 32'h3d889768} /* (26, 9, 25) {real, imag} */,
  {32'h3d4043ca, 32'hbe37dd09} /* (26, 9, 24) {real, imag} */,
  {32'hbe2a95a7, 32'h3f1e7c0c} /* (26, 9, 23) {real, imag} */,
  {32'hbe5000e1, 32'h3e41fcca} /* (26, 9, 22) {real, imag} */,
  {32'hbebb3944, 32'h3d5f0024} /* (26, 9, 21) {real, imag} */,
  {32'hbef98553, 32'h3eb64fd9} /* (26, 9, 20) {real, imag} */,
  {32'h3e6027b4, 32'h3d3d7e40} /* (26, 9, 19) {real, imag} */,
  {32'hbae87780, 32'hbd6918f8} /* (26, 9, 18) {real, imag} */,
  {32'h3d01eb24, 32'hbe1f4ecd} /* (26, 9, 17) {real, imag} */,
  {32'h3dfd3eb4, 32'h3e25602d} /* (26, 9, 16) {real, imag} */,
  {32'hbb716f80, 32'hbed8731b} /* (26, 9, 15) {real, imag} */,
  {32'hbe195e93, 32'h3e184899} /* (26, 9, 14) {real, imag} */,
  {32'h3c309090, 32'h3e320f2b} /* (26, 9, 13) {real, imag} */,
  {32'h3e0249d4, 32'h3d607770} /* (26, 9, 12) {real, imag} */,
  {32'h3dccd736, 32'h3ed71efe} /* (26, 9, 11) {real, imag} */,
  {32'hbdc2a731, 32'h3ddc49b8} /* (26, 9, 10) {real, imag} */,
  {32'h3c151d80, 32'h3e202954} /* (26, 9, 9) {real, imag} */,
  {32'h3d337f60, 32'hbf2ee746} /* (26, 9, 8) {real, imag} */,
  {32'h3e135104, 32'h3ec91233} /* (26, 9, 7) {real, imag} */,
  {32'h3ee18bc8, 32'h3e7cef79} /* (26, 9, 6) {real, imag} */,
  {32'h3ed886c1, 32'h3f496e64} /* (26, 9, 5) {real, imag} */,
  {32'h3d6d7868, 32'h3eaac05d} /* (26, 9, 4) {real, imag} */,
  {32'hbe6035e4, 32'hbe738ef4} /* (26, 9, 3) {real, imag} */,
  {32'h3e9e6240, 32'hbf01b1d4} /* (26, 9, 2) {real, imag} */,
  {32'h3e766a80, 32'hbf03b103} /* (26, 9, 1) {real, imag} */,
  {32'h3dbe6910, 32'h3ee234a0} /* (26, 9, 0) {real, imag} */,
  {32'h3d34f5b8, 32'hbf20619d} /* (26, 8, 31) {real, imag} */,
  {32'h3e8146c1, 32'hbcd93bc4} /* (26, 8, 30) {real, imag} */,
  {32'hbe6586c8, 32'hbea37e35} /* (26, 8, 29) {real, imag} */,
  {32'hbd7c5cf0, 32'h3e8ba91c} /* (26, 8, 28) {real, imag} */,
  {32'hbef31677, 32'h3e8b9ed2} /* (26, 8, 27) {real, imag} */,
  {32'hbf14bf92, 32'h3f2135f8} /* (26, 8, 26) {real, imag} */,
  {32'h3e37418c, 32'hbe915e8f} /* (26, 8, 25) {real, imag} */,
  {32'h3f72ee4d, 32'h3e60e254} /* (26, 8, 24) {real, imag} */,
  {32'hbe68adf0, 32'hbe83859c} /* (26, 8, 23) {real, imag} */,
  {32'h3c3970e0, 32'hbdc515ec} /* (26, 8, 22) {real, imag} */,
  {32'h3bc45880, 32'hbed75176} /* (26, 8, 21) {real, imag} */,
  {32'h3e3fa957, 32'h3eb2b9f2} /* (26, 8, 20) {real, imag} */,
  {32'hbf147d64, 32'hbd4f93d4} /* (26, 8, 19) {real, imag} */,
  {32'hbe222ae0, 32'h3dbc2d25} /* (26, 8, 18) {real, imag} */,
  {32'h3d7d60b4, 32'h3eb09f67} /* (26, 8, 17) {real, imag} */,
  {32'h3dfe6c3e, 32'h3dd3c554} /* (26, 8, 16) {real, imag} */,
  {32'h3e7442d3, 32'h3d48c350} /* (26, 8, 15) {real, imag} */,
  {32'h3dcf2a30, 32'h3e31f37a} /* (26, 8, 14) {real, imag} */,
  {32'h3e9836aa, 32'h3e11c576} /* (26, 8, 13) {real, imag} */,
  {32'h3cfdd9de, 32'hbd558734} /* (26, 8, 12) {real, imag} */,
  {32'h3eb2fe28, 32'hbe5cb0d9} /* (26, 8, 11) {real, imag} */,
  {32'hbee556d4, 32'hbeac036a} /* (26, 8, 10) {real, imag} */,
  {32'h3e2edc9c, 32'h3e654afa} /* (26, 8, 9) {real, imag} */,
  {32'hbf0c4e9a, 32'hbf0c6f4e} /* (26, 8, 8) {real, imag} */,
  {32'h3f285fdd, 32'hbdc430ba} /* (26, 8, 7) {real, imag} */,
  {32'h3dfa1a24, 32'h3c7a93c8} /* (26, 8, 6) {real, imag} */,
  {32'h3ecffc8f, 32'h3c0a0828} /* (26, 8, 5) {real, imag} */,
  {32'hbf2edd4e, 32'h3eedd199} /* (26, 8, 4) {real, imag} */,
  {32'h3f4b5d50, 32'h3f664b8a} /* (26, 8, 3) {real, imag} */,
  {32'hbf19902f, 32'hbe316dec} /* (26, 8, 2) {real, imag} */,
  {32'hbdec2ee0, 32'hbe154f88} /* (26, 8, 1) {real, imag} */,
  {32'hbe7b99ca, 32'hbdd622e0} /* (26, 8, 0) {real, imag} */,
  {32'hbf4d02ca, 32'h3e31503e} /* (26, 7, 31) {real, imag} */,
  {32'hbe2568ea, 32'hbe3e00ce} /* (26, 7, 30) {real, imag} */,
  {32'h3de5c368, 32'hbf0bdd00} /* (26, 7, 29) {real, imag} */,
  {32'hbe212fc0, 32'h3e024eb0} /* (26, 7, 28) {real, imag} */,
  {32'h3eff5eab, 32'h3f1a7957} /* (26, 7, 27) {real, imag} */,
  {32'hbdc2a6e4, 32'h3f1a4a94} /* (26, 7, 26) {real, imag} */,
  {32'h3c85bd58, 32'hbdc3c430} /* (26, 7, 25) {real, imag} */,
  {32'h3eb70ab3, 32'hbf5c250c} /* (26, 7, 24) {real, imag} */,
  {32'hbe8405ea, 32'h3f093669} /* (26, 7, 23) {real, imag} */,
  {32'hbd4caf44, 32'h3f058e57} /* (26, 7, 22) {real, imag} */,
  {32'h3c597660, 32'hbf1b5a6c} /* (26, 7, 21) {real, imag} */,
  {32'h3f21a452, 32'h3eb8a6ea} /* (26, 7, 20) {real, imag} */,
  {32'hbe839bfe, 32'h3ea33ede} /* (26, 7, 19) {real, imag} */,
  {32'hbece3674, 32'h3e904ae8} /* (26, 7, 18) {real, imag} */,
  {32'hbdac6782, 32'h3d028cae} /* (26, 7, 17) {real, imag} */,
  {32'hbea66cd6, 32'hbdb9db67} /* (26, 7, 16) {real, imag} */,
  {32'h3d8bc6b4, 32'h3d14ae44} /* (26, 7, 15) {real, imag} */,
  {32'hbf0daa64, 32'hbd66ab3b} /* (26, 7, 14) {real, imag} */,
  {32'hbe145503, 32'hbd6e6d0a} /* (26, 7, 13) {real, imag} */,
  {32'h3cad3028, 32'hbe8aeb84} /* (26, 7, 12) {real, imag} */,
  {32'hbe4a93f0, 32'h3f00c998} /* (26, 7, 11) {real, imag} */,
  {32'hbf55f7ba, 32'hbec8deb6} /* (26, 7, 10) {real, imag} */,
  {32'h3ef15f48, 32'h3eb859de} /* (26, 7, 9) {real, imag} */,
  {32'h3e9baaf6, 32'hbf1c95f7} /* (26, 7, 8) {real, imag} */,
  {32'hbea10d75, 32'hbe893c50} /* (26, 7, 7) {real, imag} */,
  {32'h3f23e214, 32'h3ee52827} /* (26, 7, 6) {real, imag} */,
  {32'hbeb16552, 32'hbf0c6381} /* (26, 7, 5) {real, imag} */,
  {32'h3e911ffa, 32'hbf8d3dca} /* (26, 7, 4) {real, imag} */,
  {32'h3f361906, 32'hbe015854} /* (26, 7, 3) {real, imag} */,
  {32'h3ea7aad6, 32'h3f24ae94} /* (26, 7, 2) {real, imag} */,
  {32'h3f819004, 32'h3e811cea} /* (26, 7, 1) {real, imag} */,
  {32'hbf1c5b62, 32'h3d009baa} /* (26, 7, 0) {real, imag} */,
  {32'hbed6d6fe, 32'h3da291d0} /* (26, 6, 31) {real, imag} */,
  {32'hbf2f530d, 32'h3d97ec3c} /* (26, 6, 30) {real, imag} */,
  {32'hbd91ce2a, 32'h3e1b32d6} /* (26, 6, 29) {real, imag} */,
  {32'h3eb56916, 32'hbee319dd} /* (26, 6, 28) {real, imag} */,
  {32'hbd59ea4c, 32'h3d38ed48} /* (26, 6, 27) {real, imag} */,
  {32'h3d76b1a8, 32'h3f2d71cd} /* (26, 6, 26) {real, imag} */,
  {32'hbed5871f, 32'hbec97a98} /* (26, 6, 25) {real, imag} */,
  {32'h3e69228a, 32'h3f7cf696} /* (26, 6, 24) {real, imag} */,
  {32'h3ce2ac38, 32'hbdbb0c4a} /* (26, 6, 23) {real, imag} */,
  {32'h3f0a8a17, 32'h3e9c2d76} /* (26, 6, 22) {real, imag} */,
  {32'h3e2a9500, 32'hbdb7bd48} /* (26, 6, 21) {real, imag} */,
  {32'h3e90852e, 32'h3e604f39} /* (26, 6, 20) {real, imag} */,
  {32'hbe6f3dc3, 32'hbeb6cda9} /* (26, 6, 19) {real, imag} */,
  {32'h3dc01351, 32'h3eaecd0c} /* (26, 6, 18) {real, imag} */,
  {32'hbe8e9852, 32'hbed5e600} /* (26, 6, 17) {real, imag} */,
  {32'h3e582811, 32'h3da58bd4} /* (26, 6, 16) {real, imag} */,
  {32'h3e46ad99, 32'h3e0c0473} /* (26, 6, 15) {real, imag} */,
  {32'h3e0e04ee, 32'hbbffcf08} /* (26, 6, 14) {real, imag} */,
  {32'h3ecaf7d5, 32'hbecb920b} /* (26, 6, 13) {real, imag} */,
  {32'hbedb3124, 32'h3ed31ff6} /* (26, 6, 12) {real, imag} */,
  {32'h3ef8b646, 32'hbe127c61} /* (26, 6, 11) {real, imag} */,
  {32'hbe1d473b, 32'h3d7eb7f8} /* (26, 6, 10) {real, imag} */,
  {32'h3f22bcbd, 32'hbed876c0} /* (26, 6, 9) {real, imag} */,
  {32'h3f0e19d2, 32'h3ea38252} /* (26, 6, 8) {real, imag} */,
  {32'h3ea518f8, 32'h3d13e8c0} /* (26, 6, 7) {real, imag} */,
  {32'h3f108912, 32'hbf01811d} /* (26, 6, 6) {real, imag} */,
  {32'h3d1778f8, 32'h3ed8a6c5} /* (26, 6, 5) {real, imag} */,
  {32'hbe436798, 32'hbee14baa} /* (26, 6, 4) {real, imag} */,
  {32'h3f2137d9, 32'hbee20997} /* (26, 6, 3) {real, imag} */,
  {32'h3e8e4984, 32'h3d80b062} /* (26, 6, 2) {real, imag} */,
  {32'hbe4004ec, 32'h3e857943} /* (26, 6, 1) {real, imag} */,
  {32'h3ed62ce8, 32'hbefb96c0} /* (26, 6, 0) {real, imag} */,
  {32'hbdd94940, 32'hbf9dd99e} /* (26, 5, 31) {real, imag} */,
  {32'h3f0ed5a4, 32'hbea4b4dc} /* (26, 5, 30) {real, imag} */,
  {32'h3f57bcd2, 32'h3d84fff4} /* (26, 5, 29) {real, imag} */,
  {32'hbebbbcf3, 32'h3f2e4bd0} /* (26, 5, 28) {real, imag} */,
  {32'hbef5a32e, 32'hbea2b9dc} /* (26, 5, 27) {real, imag} */,
  {32'h3e067d77, 32'hbd1902e2} /* (26, 5, 26) {real, imag} */,
  {32'h3d523fa2, 32'hbeb11360} /* (26, 5, 25) {real, imag} */,
  {32'h3d78d904, 32'hbe2b74c9} /* (26, 5, 24) {real, imag} */,
  {32'hbed80ee4, 32'h3ed8e888} /* (26, 5, 23) {real, imag} */,
  {32'h3ee173d6, 32'hbb224080} /* (26, 5, 22) {real, imag} */,
  {32'h3ddbec2a, 32'hbece430a} /* (26, 5, 21) {real, imag} */,
  {32'h3f1e6ae0, 32'h3e1c0209} /* (26, 5, 20) {real, imag} */,
  {32'h3e8ab40e, 32'h3efecbca} /* (26, 5, 19) {real, imag} */,
  {32'h3e5b013e, 32'hbea715ae} /* (26, 5, 18) {real, imag} */,
  {32'h3d15362c, 32'hbe8950ce} /* (26, 5, 17) {real, imag} */,
  {32'hbec34b38, 32'hbefb725a} /* (26, 5, 16) {real, imag} */,
  {32'hbdd9c69c, 32'h3d8683e4} /* (26, 5, 15) {real, imag} */,
  {32'hbe04cea8, 32'hbc732e20} /* (26, 5, 14) {real, imag} */,
  {32'hbeb8e9fa, 32'h3ef44ae4} /* (26, 5, 13) {real, imag} */,
  {32'hbe086714, 32'h3cb91f70} /* (26, 5, 12) {real, imag} */,
  {32'h3dde159d, 32'h3f0b5dbe} /* (26, 5, 11) {real, imag} */,
  {32'h3e9af272, 32'h3de562d2} /* (26, 5, 10) {real, imag} */,
  {32'h3ebbe2b8, 32'hbc82f2b0} /* (26, 5, 9) {real, imag} */,
  {32'h3f53f6e6, 32'hbe5b83d6} /* (26, 5, 8) {real, imag} */,
  {32'h3f1a4e22, 32'h3eead4a6} /* (26, 5, 7) {real, imag} */,
  {32'hbf3b1a1a, 32'h3ee1ca44} /* (26, 5, 6) {real, imag} */,
  {32'h3ef9b22f, 32'h3d3681c0} /* (26, 5, 5) {real, imag} */,
  {32'hbdf14a65, 32'hbe80f6d3} /* (26, 5, 4) {real, imag} */,
  {32'hbee61926, 32'hbf3aee14} /* (26, 5, 3) {real, imag} */,
  {32'hbf1275bd, 32'hbeb67f6a} /* (26, 5, 2) {real, imag} */,
  {32'hbf8a3bc1, 32'h3ea24b98} /* (26, 5, 1) {real, imag} */,
  {32'hbfd69100, 32'h3f24f675} /* (26, 5, 0) {real, imag} */,
  {32'hbec5a5e2, 32'hbd869b28} /* (26, 4, 31) {real, imag} */,
  {32'hbeb5daee, 32'hbe0d1a58} /* (26, 4, 30) {real, imag} */,
  {32'hbf44089d, 32'h3da2a804} /* (26, 4, 29) {real, imag} */,
  {32'h3cb463f0, 32'hbeaaf775} /* (26, 4, 28) {real, imag} */,
  {32'h3cfb8754, 32'h3e0909d3} /* (26, 4, 27) {real, imag} */,
  {32'hbf405772, 32'hbed577c5} /* (26, 4, 26) {real, imag} */,
  {32'hbd3bdcce, 32'h3f96858b} /* (26, 4, 25) {real, imag} */,
  {32'h3db5ab34, 32'hbeb27150} /* (26, 4, 24) {real, imag} */,
  {32'hbb3ba040, 32'h3e8e73ad} /* (26, 4, 23) {real, imag} */,
  {32'h3f3acb31, 32'h3e8cd3cf} /* (26, 4, 22) {real, imag} */,
  {32'hbe271056, 32'h3f22e4f0} /* (26, 4, 21) {real, imag} */,
  {32'h3e203a5c, 32'h3d9e0994} /* (26, 4, 20) {real, imag} */,
  {32'hbc54757e, 32'hbe4b3a8b} /* (26, 4, 19) {real, imag} */,
  {32'hbf1eec98, 32'hbe903573} /* (26, 4, 18) {real, imag} */,
  {32'h3e3946b8, 32'hbd4985fc} /* (26, 4, 17) {real, imag} */,
  {32'hbe15c904, 32'hbd3ce1d4} /* (26, 4, 16) {real, imag} */,
  {32'hbef50474, 32'hbe058686} /* (26, 4, 15) {real, imag} */,
  {32'hbe835352, 32'h3d3cd410} /* (26, 4, 14) {real, imag} */,
  {32'h3dc4e50e, 32'h3eb86426} /* (26, 4, 13) {real, imag} */,
  {32'hbebca03f, 32'hbe97b227} /* (26, 4, 12) {real, imag} */,
  {32'h3f255f87, 32'h3e992c14} /* (26, 4, 11) {real, imag} */,
  {32'h3e056319, 32'hbe261476} /* (26, 4, 10) {real, imag} */,
  {32'hbe3a6adf, 32'h3dc6e62c} /* (26, 4, 9) {real, imag} */,
  {32'h3d8c760c, 32'hbe908507} /* (26, 4, 8) {real, imag} */,
  {32'hbda0d54c, 32'h3eca25f4} /* (26, 4, 7) {real, imag} */,
  {32'hbf178266, 32'h3e9c6e08} /* (26, 4, 6) {real, imag} */,
  {32'h3edaaf09, 32'hbd2faf24} /* (26, 4, 5) {real, imag} */,
  {32'h3f2e8843, 32'hbf6872be} /* (26, 4, 4) {real, imag} */,
  {32'hbdc716f6, 32'hbe0587e6} /* (26, 4, 3) {real, imag} */,
  {32'hbee73dec, 32'hbe08d008} /* (26, 4, 2) {real, imag} */,
  {32'h3ed80fc8, 32'h3eb5c77a} /* (26, 4, 1) {real, imag} */,
  {32'hbf2c42ca, 32'hbf7c5812} /* (26, 4, 0) {real, imag} */,
  {32'hbf57bc14, 32'h3e117fc8} /* (26, 3, 31) {real, imag} */,
  {32'h3fc90e17, 32'hbedf3e10} /* (26, 3, 30) {real, imag} */,
  {32'h3eabdac1, 32'h3d84177e} /* (26, 3, 29) {real, imag} */,
  {32'h3f1f5ad8, 32'h3f0a913f} /* (26, 3, 28) {real, imag} */,
  {32'hbd96b900, 32'hbe7044af} /* (26, 3, 27) {real, imag} */,
  {32'hbea94fdf, 32'h3edd9480} /* (26, 3, 26) {real, imag} */,
  {32'hbf2f19f9, 32'h3d0f2c90} /* (26, 3, 25) {real, imag} */,
  {32'hbe60c97e, 32'hbeba0988} /* (26, 3, 24) {real, imag} */,
  {32'h3e4392fb, 32'hbe9680ba} /* (26, 3, 23) {real, imag} */,
  {32'hbd83b432, 32'h3e2bd33f} /* (26, 3, 22) {real, imag} */,
  {32'h3c9af8c0, 32'h3e29174a} /* (26, 3, 21) {real, imag} */,
  {32'hbeb7af6a, 32'hbdf3e51a} /* (26, 3, 20) {real, imag} */,
  {32'h3ec3a574, 32'hbe4c9c4c} /* (26, 3, 19) {real, imag} */,
  {32'hbea8e9d6, 32'hbf1d1ad3} /* (26, 3, 18) {real, imag} */,
  {32'h3f1344da, 32'h3e52d840} /* (26, 3, 17) {real, imag} */,
  {32'h3e076e9e, 32'h3e8184ef} /* (26, 3, 16) {real, imag} */,
  {32'hbe10ab61, 32'hbe4e1dc2} /* (26, 3, 15) {real, imag} */,
  {32'h3dcc7684, 32'h3f0498f4} /* (26, 3, 14) {real, imag} */,
  {32'h3ea11535, 32'hbf0d7278} /* (26, 3, 13) {real, imag} */,
  {32'h3e7e260e, 32'hbe972ce0} /* (26, 3, 12) {real, imag} */,
  {32'h3d801bc2, 32'hbe236302} /* (26, 3, 11) {real, imag} */,
  {32'hbe88d650, 32'hbdc4720a} /* (26, 3, 10) {real, imag} */,
  {32'hbe0c4b2c, 32'hbe7e9390} /* (26, 3, 9) {real, imag} */,
  {32'hbe6ee221, 32'hbecd4281} /* (26, 3, 8) {real, imag} */,
  {32'hbdf6243c, 32'h3eea9a5a} /* (26, 3, 7) {real, imag} */,
  {32'hbee8f290, 32'h3edbf076} /* (26, 3, 6) {real, imag} */,
  {32'hbef03418, 32'h3ed9f036} /* (26, 3, 5) {real, imag} */,
  {32'hbe3efcea, 32'h3ee4205d} /* (26, 3, 4) {real, imag} */,
  {32'hbf029350, 32'hbcd002e0} /* (26, 3, 3) {real, imag} */,
  {32'h3f52df75, 32'hbe75bf94} /* (26, 3, 2) {real, imag} */,
  {32'hbde03680, 32'h4014a578} /* (26, 3, 1) {real, imag} */,
  {32'h401e92db, 32'h3f7d20d5} /* (26, 3, 0) {real, imag} */,
  {32'h3f35c9e0, 32'h3ff760bc} /* (26, 2, 31) {real, imag} */,
  {32'h3fe2fe10, 32'hbff918f2} /* (26, 2, 30) {real, imag} */,
  {32'hbeb4a8ec, 32'hbe68e93e} /* (26, 2, 29) {real, imag} */,
  {32'hbec1df94, 32'h3eb3531a} /* (26, 2, 28) {real, imag} */,
  {32'h3f6b715f, 32'hbf3ef157} /* (26, 2, 27) {real, imag} */,
  {32'h3e34bb75, 32'h3edf0e50} /* (26, 2, 26) {real, imag} */,
  {32'hbe3ffe56, 32'h3fa1b930} /* (26, 2, 25) {real, imag} */,
  {32'h3f2afec6, 32'h3ea8d31d} /* (26, 2, 24) {real, imag} */,
  {32'h3f65fcf9, 32'hbeeee2d3} /* (26, 2, 23) {real, imag} */,
  {32'hbec06eb2, 32'hbdb6331e} /* (26, 2, 22) {real, imag} */,
  {32'h3e039c7c, 32'h3d3ffd80} /* (26, 2, 21) {real, imag} */,
  {32'hbe70bd3f, 32'hbc738940} /* (26, 2, 20) {real, imag} */,
  {32'hbe766dda, 32'hbd0b2cb8} /* (26, 2, 19) {real, imag} */,
  {32'h3e9b1964, 32'h3ec0c8cf} /* (26, 2, 18) {real, imag} */,
  {32'h3e9aa0ae, 32'h3e7dfd77} /* (26, 2, 17) {real, imag} */,
  {32'h3d9e675e, 32'h3e39f76d} /* (26, 2, 16) {real, imag} */,
  {32'hbceed506, 32'hbe448894} /* (26, 2, 15) {real, imag} */,
  {32'hbe026a38, 32'hbe6aaffa} /* (26, 2, 14) {real, imag} */,
  {32'hbdefe79e, 32'h3d790ac2} /* (26, 2, 13) {real, imag} */,
  {32'h3e3793f8, 32'h3d879494} /* (26, 2, 12) {real, imag} */,
  {32'h3edede48, 32'h3e8115e9} /* (26, 2, 11) {real, imag} */,
  {32'h3c5b00b0, 32'h3d99b554} /* (26, 2, 10) {real, imag} */,
  {32'hbf14259f, 32'hbed2f550} /* (26, 2, 9) {real, imag} */,
  {32'hbe145796, 32'h3f28f5c5} /* (26, 2, 8) {real, imag} */,
  {32'h3e4ef612, 32'h3f4366d6} /* (26, 2, 7) {real, imag} */,
  {32'h3ee09cbe, 32'h3e43c967} /* (26, 2, 6) {real, imag} */,
  {32'hbf13011d, 32'h3fa263f2} /* (26, 2, 5) {real, imag} */,
  {32'hbf114d0c, 32'hbf94c973} /* (26, 2, 4) {real, imag} */,
  {32'hbf7537d2, 32'hbeb5a3bb} /* (26, 2, 3) {real, imag} */,
  {32'h40061f12, 32'hbf5c8ee8} /* (26, 2, 2) {real, imag} */,
  {32'h3e359680, 32'h4008b118} /* (26, 2, 1) {real, imag} */,
  {32'h3fd3d7cc, 32'hc00b7808} /* (26, 2, 0) {real, imag} */,
  {32'hc0d6de14, 32'h3d8695e0} /* (26, 1, 31) {real, imag} */,
  {32'h3efa1570, 32'h4058bf26} /* (26, 1, 30) {real, imag} */,
  {32'h3e6986d4, 32'hbd490a00} /* (26, 1, 29) {real, imag} */,
  {32'hbee9817a, 32'h3f141052} /* (26, 1, 28) {real, imag} */,
  {32'hbf147850, 32'hbbc16300} /* (26, 1, 27) {real, imag} */,
  {32'hbf560d2d, 32'hbe81b218} /* (26, 1, 26) {real, imag} */,
  {32'hbe4ce52e, 32'hbea8f8e9} /* (26, 1, 25) {real, imag} */,
  {32'h3e857d44, 32'hbe0516f1} /* (26, 1, 24) {real, imag} */,
  {32'h3e8e2b92, 32'h3bf921c0} /* (26, 1, 23) {real, imag} */,
  {32'h3d813678, 32'h3e2848ee} /* (26, 1, 22) {real, imag} */,
  {32'hbd65da08, 32'hbeb55303} /* (26, 1, 21) {real, imag} */,
  {32'h3eb9e5a6, 32'h3f08db82} /* (26, 1, 20) {real, imag} */,
  {32'h3f050d11, 32'hbe3e3764} /* (26, 1, 19) {real, imag} */,
  {32'h3eb03ef8, 32'h3d35c9a4} /* (26, 1, 18) {real, imag} */,
  {32'h3e03bd20, 32'hbe7c0667} /* (26, 1, 17) {real, imag} */,
  {32'hbe7f199a, 32'hbd6a115d} /* (26, 1, 16) {real, imag} */,
  {32'hbb64a4c0, 32'hbd080bcc} /* (26, 1, 15) {real, imag} */,
  {32'h3dfe397a, 32'hbe23ba98} /* (26, 1, 14) {real, imag} */,
  {32'h3f595d35, 32'h3e129d18} /* (26, 1, 13) {real, imag} */,
  {32'h3e8907c2, 32'h3eca5faa} /* (26, 1, 12) {real, imag} */,
  {32'hbf1d1598, 32'h3d032e10} /* (26, 1, 11) {real, imag} */,
  {32'hbf5ccbee, 32'h3c483278} /* (26, 1, 10) {real, imag} */,
  {32'hbf2e7514, 32'h3d143fe0} /* (26, 1, 9) {real, imag} */,
  {32'hbeab1098, 32'hbf1a6005} /* (26, 1, 8) {real, imag} */,
  {32'h3eb69168, 32'h3f26c130} /* (26, 1, 7) {real, imag} */,
  {32'h3eef0c36, 32'hbdaae662} /* (26, 1, 6) {real, imag} */,
  {32'h3d6f3620, 32'h3ea47a2e} /* (26, 1, 5) {real, imag} */,
  {32'hbf12dc72, 32'hbf00c656} /* (26, 1, 4) {real, imag} */,
  {32'h3be7c600, 32'hbf330c6c} /* (26, 1, 3) {real, imag} */,
  {32'hbf7ce798, 32'hbf8169f4} /* (26, 1, 2) {real, imag} */,
  {32'hc1110940, 32'hc0dc801d} /* (26, 1, 1) {real, imag} */,
  {32'hc168fd6c, 32'hc053370a} /* (26, 1, 0) {real, imag} */,
  {32'hc15295f2, 32'h412ab656} /* (26, 0, 31) {real, imag} */,
  {32'hbf2f3b58, 32'h40248ee9} /* (26, 0, 30) {real, imag} */,
  {32'h3eef01e6, 32'hbfb0bae8} /* (26, 0, 29) {real, imag} */,
  {32'h3fa1e952, 32'hbebe3a2c} /* (26, 0, 28) {real, imag} */,
  {32'hbdc04dc0, 32'h3e74e91e} /* (26, 0, 27) {real, imag} */,
  {32'h3f28150f, 32'hbe0dcab4} /* (26, 0, 26) {real, imag} */,
  {32'h3e9e15f6, 32'hbe82dc65} /* (26, 0, 25) {real, imag} */,
  {32'h3e18ebc2, 32'hbf5b92e7} /* (26, 0, 24) {real, imag} */,
  {32'hbf1a73f1, 32'hbdf1062f} /* (26, 0, 23) {real, imag} */,
  {32'hbebf310c, 32'h3ed0c886} /* (26, 0, 22) {real, imag} */,
  {32'hbdc88daa, 32'h3f23c9df} /* (26, 0, 21) {real, imag} */,
  {32'hbc7053d0, 32'hbea51f12} /* (26, 0, 20) {real, imag} */,
  {32'hbe646985, 32'hbdb2e116} /* (26, 0, 19) {real, imag} */,
  {32'h3e199450, 32'h3e115b58} /* (26, 0, 18) {real, imag} */,
  {32'h3e11214c, 32'h3d55a837} /* (26, 0, 17) {real, imag} */,
  {32'h3f3fb9f6, 32'h00000000} /* (26, 0, 16) {real, imag} */,
  {32'h3e11214c, 32'hbd55a837} /* (26, 0, 15) {real, imag} */,
  {32'h3e199450, 32'hbe115b58} /* (26, 0, 14) {real, imag} */,
  {32'hbe646985, 32'h3db2e116} /* (26, 0, 13) {real, imag} */,
  {32'hbc7053d0, 32'h3ea51f12} /* (26, 0, 12) {real, imag} */,
  {32'hbdc88daa, 32'hbf23c9df} /* (26, 0, 11) {real, imag} */,
  {32'hbebf310c, 32'hbed0c886} /* (26, 0, 10) {real, imag} */,
  {32'hbf1a73f1, 32'h3df1062f} /* (26, 0, 9) {real, imag} */,
  {32'h3e18ebc2, 32'h3f5b92e7} /* (26, 0, 8) {real, imag} */,
  {32'h3e9e15f6, 32'h3e82dc65} /* (26, 0, 7) {real, imag} */,
  {32'h3f28150f, 32'h3e0dcab4} /* (26, 0, 6) {real, imag} */,
  {32'hbdc04dc0, 32'hbe74e91e} /* (26, 0, 5) {real, imag} */,
  {32'h3fa1e952, 32'h3ebe3a2c} /* (26, 0, 4) {real, imag} */,
  {32'h3eef01e6, 32'h3fb0bae8} /* (26, 0, 3) {real, imag} */,
  {32'hbf2f3b58, 32'hc0248ee9} /* (26, 0, 2) {real, imag} */,
  {32'hc15295f2, 32'hc12ab656} /* (26, 0, 1) {real, imag} */,
  {32'hc1ec0ae3, 32'h00000000} /* (26, 0, 0) {real, imag} */,
  {32'hc2124069, 32'h41aea98b} /* (25, 31, 31) {real, imag} */,
  {32'h410543ce, 32'hc10875b1} /* (25, 31, 30) {real, imag} */,
  {32'h3f9710a7, 32'h3d25f380} /* (25, 31, 29) {real, imag} */,
  {32'hbd8a35c0, 32'h3ff53126} /* (25, 31, 28) {real, imag} */,
  {32'h3fc05e16, 32'hbfb57b70} /* (25, 31, 27) {real, imag} */,
  {32'h3eef6cb3, 32'hbefe8b53} /* (25, 31, 26) {real, imag} */,
  {32'hbe01714b, 32'hbdb48370} /* (25, 31, 25) {real, imag} */,
  {32'h3e83e51f, 32'hbf7b5807} /* (25, 31, 24) {real, imag} */,
  {32'h3e8b0e3d, 32'h3e8b89ba} /* (25, 31, 23) {real, imag} */,
  {32'h3e389066, 32'hbd2bb4a8} /* (25, 31, 22) {real, imag} */,
  {32'h3ec42a38, 32'hbf483c00} /* (25, 31, 21) {real, imag} */,
  {32'hbd374e4e, 32'hbd64efcc} /* (25, 31, 20) {real, imag} */,
  {32'h3e569b90, 32'h3e6a93da} /* (25, 31, 19) {real, imag} */,
  {32'hbebaaa8d, 32'hbef0d1e0} /* (25, 31, 18) {real, imag} */,
  {32'hbea3ad74, 32'h3eeb3d5f} /* (25, 31, 17) {real, imag} */,
  {32'h3d9de935, 32'hbeacee39} /* (25, 31, 16) {real, imag} */,
  {32'hbddd30c6, 32'hbe1e5d68} /* (25, 31, 15) {real, imag} */,
  {32'h3e4e2313, 32'h3f07981c} /* (25, 31, 14) {real, imag} */,
  {32'hbe3bd3fd, 32'h3ce73428} /* (25, 31, 13) {real, imag} */,
  {32'h3ecf9a2e, 32'h3df55af7} /* (25, 31, 12) {real, imag} */,
  {32'h3f412222, 32'h3ef21ba8} /* (25, 31, 11) {real, imag} */,
  {32'hbd68b750, 32'h3f07fb38} /* (25, 31, 10) {real, imag} */,
  {32'h3d8856a9, 32'hbef2155e} /* (25, 31, 9) {real, imag} */,
  {32'h3d6e04f0, 32'h3d3b3408} /* (25, 31, 8) {real, imag} */,
  {32'hbf00ef26, 32'hbea83732} /* (25, 31, 7) {real, imag} */,
  {32'hbf3494fb, 32'h3e2bd18c} /* (25, 31, 6) {real, imag} */,
  {32'h40078014, 32'h3ece00d6} /* (25, 31, 5) {real, imag} */,
  {32'hbfa3353e, 32'h3f48d99e} /* (25, 31, 4) {real, imag} */,
  {32'h3f5217c5, 32'h3f2fe7c8} /* (25, 31, 3) {real, imag} */,
  {32'h40bc3442, 32'hc05fe528} /* (25, 31, 2) {real, imag} */,
  {32'hc1c64ef4, 32'hc0b23f18} /* (25, 31, 1) {real, imag} */,
  {32'hc213f352, 32'h40bfcf31} /* (25, 31, 0) {real, imag} */,
  {32'h4131396f, 32'hbf0b3d40} /* (25, 30, 31) {real, imag} */,
  {32'hc0ab65b9, 32'hbf935d2d} /* (25, 30, 30) {real, imag} */,
  {32'hbf1386fb, 32'h3e7806b4} /* (25, 30, 29) {real, imag} */,
  {32'h3fc30485, 32'h3dce70f4} /* (25, 30, 28) {real, imag} */,
  {32'hc00778e3, 32'h3f8769b3} /* (25, 30, 27) {real, imag} */,
  {32'hbe22a9fe, 32'h3ec3250d} /* (25, 30, 26) {real, imag} */,
  {32'h3f6a4924, 32'hbee9d390} /* (25, 30, 25) {real, imag} */,
  {32'hbf07854d, 32'h3e587b6e} /* (25, 30, 24) {real, imag} */,
  {32'hbd2b8274, 32'h3eecc5f6} /* (25, 30, 23) {real, imag} */,
  {32'h3edf2f14, 32'hbe860087} /* (25, 30, 22) {real, imag} */,
  {32'hbe5a26df, 32'h3f6ec50f} /* (25, 30, 21) {real, imag} */,
  {32'hbd33a4a8, 32'h3f15536b} /* (25, 30, 20) {real, imag} */,
  {32'h3e89a426, 32'hbd17197c} /* (25, 30, 19) {real, imag} */,
  {32'hbd67cd48, 32'hbed03225} /* (25, 30, 18) {real, imag} */,
  {32'h3e60c574, 32'hbe1a5ed1} /* (25, 30, 17) {real, imag} */,
  {32'hbe6a1156, 32'hbe4d9fe1} /* (25, 30, 16) {real, imag} */,
  {32'hbe548374, 32'h3ecddffa} /* (25, 30, 15) {real, imag} */,
  {32'hbe23d4f4, 32'hbe7016c0} /* (25, 30, 14) {real, imag} */,
  {32'h3ca437cc, 32'hbd7024f4} /* (25, 30, 13) {real, imag} */,
  {32'hbc0bf2b0, 32'h3e739ca0} /* (25, 30, 12) {real, imag} */,
  {32'hbdb7db4a, 32'h3e96d028} /* (25, 30, 11) {real, imag} */,
  {32'h3e707241, 32'h3f487158} /* (25, 30, 10) {real, imag} */,
  {32'h3e8fe85f, 32'hbca23f38} /* (25, 30, 9) {real, imag} */,
  {32'hbecca1ad, 32'hbf822582} /* (25, 30, 8) {real, imag} */,
  {32'hb92f1800, 32'hbf792af4} /* (25, 30, 7) {real, imag} */,
  {32'h3e48d3e0, 32'hbcc123f0} /* (25, 30, 6) {real, imag} */,
  {32'h3d18c7f0, 32'h3ed2c160} /* (25, 30, 5) {real, imag} */,
  {32'h3f80646f, 32'h3f9d9bb9} /* (25, 30, 4) {real, imag} */,
  {32'h3f4b205e, 32'h3f652d8e} /* (25, 30, 3) {real, imag} */,
  {32'hc10b0d3a, 32'hbfcb1585} /* (25, 30, 2) {real, imag} */,
  {32'h41924ac2, 32'hc0174649} /* (25, 30, 1) {real, imag} */,
  {32'h412f9197, 32'hbf21350c} /* (25, 30, 0) {real, imag} */,
  {32'hc03703a1, 32'h3fbc75bf} /* (25, 29, 31) {real, imag} */,
  {32'h3e43a557, 32'hc03cd155} /* (25, 29, 30) {real, imag} */,
  {32'hbd8c1486, 32'h3f0dcfcd} /* (25, 29, 29) {real, imag} */,
  {32'h3f45d2e2, 32'h3e2516c8} /* (25, 29, 28) {real, imag} */,
  {32'hbf52fc5e, 32'h3ef5dcd8} /* (25, 29, 27) {real, imag} */,
  {32'hbdb549d8, 32'hbf0e9266} /* (25, 29, 26) {real, imag} */,
  {32'hbe42ff4c, 32'hbd0d42be} /* (25, 29, 25) {real, imag} */,
  {32'hbebb0c1e, 32'h3e84cd56} /* (25, 29, 24) {real, imag} */,
  {32'hbd883f66, 32'h3e6a6a4a} /* (25, 29, 23) {real, imag} */,
  {32'hbd6a2caa, 32'hbdbe7304} /* (25, 29, 22) {real, imag} */,
  {32'hbf0a8f00, 32'h3dd29ac4} /* (25, 29, 21) {real, imag} */,
  {32'h3ec8094d, 32'h3e25df7a} /* (25, 29, 20) {real, imag} */,
  {32'h3dbf0a54, 32'hbe83a276} /* (25, 29, 19) {real, imag} */,
  {32'hbee609ca, 32'h3dd111b2} /* (25, 29, 18) {real, imag} */,
  {32'h3de1958c, 32'hbda6a4b7} /* (25, 29, 17) {real, imag} */,
  {32'hbe59fbd5, 32'hbe4ecdf1} /* (25, 29, 16) {real, imag} */,
  {32'h3b8c44b8, 32'h3e346f5d} /* (25, 29, 15) {real, imag} */,
  {32'h3e991012, 32'hbe39eeae} /* (25, 29, 14) {real, imag} */,
  {32'h3ec8745a, 32'h3e2fd396} /* (25, 29, 13) {real, imag} */,
  {32'hbdbf1ab9, 32'hbeaed7a0} /* (25, 29, 12) {real, imag} */,
  {32'hbd0d6c22, 32'hbe4910e0} /* (25, 29, 11) {real, imag} */,
  {32'hbe0e16be, 32'hbe69ba4a} /* (25, 29, 10) {real, imag} */,
  {32'h3df369b4, 32'h3ee92c34} /* (25, 29, 9) {real, imag} */,
  {32'h3ede588d, 32'hbf5b916c} /* (25, 29, 8) {real, imag} */,
  {32'h3e49f958, 32'hbe89e0fa} /* (25, 29, 7) {real, imag} */,
  {32'hbcab5230, 32'hbe54ba12} /* (25, 29, 6) {real, imag} */,
  {32'h3eeabea8, 32'h3d9821e8} /* (25, 29, 5) {real, imag} */,
  {32'hbf4e4370, 32'h3f208bd4} /* (25, 29, 4) {real, imag} */,
  {32'h3f2ddf9e, 32'hbed80e26} /* (25, 29, 3) {real, imag} */,
  {32'hbea3e0a8, 32'hbfebde3d} /* (25, 29, 2) {real, imag} */,
  {32'h400d6642, 32'h401f3f28} /* (25, 29, 1) {real, imag} */,
  {32'h401cc1ef, 32'hbf1c36dc} /* (25, 29, 0) {real, imag} */,
  {32'hc06053b4, 32'h3f01c330} /* (25, 28, 31) {real, imag} */,
  {32'h3fe4ec3e, 32'hbfc350b5} /* (25, 28, 30) {real, imag} */,
  {32'hbe24025c, 32'h3dfdc67a} /* (25, 28, 29) {real, imag} */,
  {32'h3e91834b, 32'h3ffeae9b} /* (25, 28, 28) {real, imag} */,
  {32'h3e96da0c, 32'hbb918b80} /* (25, 28, 27) {real, imag} */,
  {32'hbf4d1b52, 32'hbf536dd4} /* (25, 28, 26) {real, imag} */,
  {32'hbf37d815, 32'hbe9fd46d} /* (25, 28, 25) {real, imag} */,
  {32'h3efb6267, 32'hbf7982f6} /* (25, 28, 24) {real, imag} */,
  {32'hbe74b68c, 32'hbebc036e} /* (25, 28, 23) {real, imag} */,
  {32'h3d980685, 32'h3e1312d3} /* (25, 28, 22) {real, imag} */,
  {32'h3eaafa78, 32'hbf2e7fa2} /* (25, 28, 21) {real, imag} */,
  {32'h3da51f20, 32'h3cdf4f30} /* (25, 28, 20) {real, imag} */,
  {32'h3e8253f6, 32'hbe61c37c} /* (25, 28, 19) {real, imag} */,
  {32'h3d73a3e0, 32'h3dff2100} /* (25, 28, 18) {real, imag} */,
  {32'hbe341313, 32'h3d2bce2c} /* (25, 28, 17) {real, imag} */,
  {32'hbc7c99fe, 32'hbe3ab18a} /* (25, 28, 16) {real, imag} */,
  {32'h3d45be7c, 32'hbe68a313} /* (25, 28, 15) {real, imag} */,
  {32'h3f0e9bee, 32'h3e13e7d0} /* (25, 28, 14) {real, imag} */,
  {32'hbe653144, 32'hbe867ab2} /* (25, 28, 13) {real, imag} */,
  {32'h3d696b78, 32'h3c433560} /* (25, 28, 12) {real, imag} */,
  {32'h3e62c443, 32'hbf053101} /* (25, 28, 11) {real, imag} */,
  {32'hbeba97a6, 32'h3e2cdbc0} /* (25, 28, 10) {real, imag} */,
  {32'hbe10bfea, 32'h3e66ab51} /* (25, 28, 9) {real, imag} */,
  {32'h3c90c830, 32'hbde8e8d0} /* (25, 28, 8) {real, imag} */,
  {32'h3e8a4d82, 32'hbe9e4403} /* (25, 28, 7) {real, imag} */,
  {32'hbdf8bcd8, 32'h3f579b3c} /* (25, 28, 6) {real, imag} */,
  {32'h3e4167df, 32'h3c4b2e10} /* (25, 28, 5) {real, imag} */,
  {32'hbf89d772, 32'h3f9a93f5} /* (25, 28, 4) {real, imag} */,
  {32'hbf1e76c3, 32'h3e755a6e} /* (25, 28, 3) {real, imag} */,
  {32'h3fabde28, 32'hc012508d} /* (25, 28, 2) {real, imag} */,
  {32'hbf8b4cb0, 32'h400ba980} /* (25, 28, 1) {real, imag} */,
  {32'hbfca60d6, 32'h3f974fad} /* (25, 28, 0) {real, imag} */,
  {32'h3fb88489, 32'hc01edf1e} /* (25, 27, 31) {real, imag} */,
  {32'hbf8556c6, 32'h3fa8ec60} /* (25, 27, 30) {real, imag} */,
  {32'h3cf11870, 32'h3f82c8a4} /* (25, 27, 29) {real, imag} */,
  {32'hbeb81486, 32'hbed95528} /* (25, 27, 28) {real, imag} */,
  {32'h3f65cf84, 32'h3e976e91} /* (25, 27, 27) {real, imag} */,
  {32'hbdc0d3c8, 32'hbe1cdadc} /* (25, 27, 26) {real, imag} */,
  {32'h3e97b582, 32'hbe827211} /* (25, 27, 25) {real, imag} */,
  {32'hbda8b09c, 32'h3d838a04} /* (25, 27, 24) {real, imag} */,
  {32'hbf0dab18, 32'h3ebfb2b6} /* (25, 27, 23) {real, imag} */,
  {32'h3d5e39b0, 32'h3eed6cd6} /* (25, 27, 22) {real, imag} */,
  {32'hbdcce098, 32'h3f3890b6} /* (25, 27, 21) {real, imag} */,
  {32'h3d1fd11a, 32'hbe7f99e8} /* (25, 27, 20) {real, imag} */,
  {32'hbb969f78, 32'hbe5badc2} /* (25, 27, 19) {real, imag} */,
  {32'h3e28aa02, 32'hbe804d78} /* (25, 27, 18) {real, imag} */,
  {32'hbdd8e84e, 32'hbec93f97} /* (25, 27, 17) {real, imag} */,
  {32'h3d4f91ec, 32'hbc8a0bb8} /* (25, 27, 16) {real, imag} */,
  {32'hbee69352, 32'h3d8d9da0} /* (25, 27, 15) {real, imag} */,
  {32'hbda05594, 32'hbed6eca8} /* (25, 27, 14) {real, imag} */,
  {32'h3eb5ffe8, 32'hbdc797a1} /* (25, 27, 13) {real, imag} */,
  {32'h3ee4da6b, 32'hbe175e26} /* (25, 27, 12) {real, imag} */,
  {32'hbef1087e, 32'h3cbe75d8} /* (25, 27, 11) {real, imag} */,
  {32'h3e2c70bd, 32'hbe53b53e} /* (25, 27, 10) {real, imag} */,
  {32'hbe086c84, 32'h3e89edc8} /* (25, 27, 9) {real, imag} */,
  {32'hbe208e68, 32'hbec77fd0} /* (25, 27, 8) {real, imag} */,
  {32'h3f1d87ad, 32'h3eec0be0} /* (25, 27, 7) {real, imag} */,
  {32'h3f3a2781, 32'h3ecdc8c2} /* (25, 27, 6) {real, imag} */,
  {32'hbfa3f762, 32'hbe6e848c} /* (25, 27, 5) {real, imag} */,
  {32'h3e141bb5, 32'hbefb89ec} /* (25, 27, 4) {real, imag} */,
  {32'h3eb91df4, 32'h3e63ff62} /* (25, 27, 3) {real, imag} */,
  {32'hbf879cda, 32'h3f587950} /* (25, 27, 2) {real, imag} */,
  {32'h4028f802, 32'h3f04a4e4} /* (25, 27, 1) {real, imag} */,
  {32'h3f89b2dc, 32'hbfcb057a} /* (25, 27, 0) {real, imag} */,
  {32'hbe1640a1, 32'hbe398f75} /* (25, 26, 31) {real, imag} */,
  {32'h3f432d6e, 32'h3e04b04c} /* (25, 26, 30) {real, imag} */,
  {32'h3e25fac4, 32'h3e080ab0} /* (25, 26, 29) {real, imag} */,
  {32'h3e49778e, 32'h3f3c6d8d} /* (25, 26, 28) {real, imag} */,
  {32'h3e14659c, 32'h3cb9a474} /* (25, 26, 27) {real, imag} */,
  {32'h3edf8948, 32'h3eb474fc} /* (25, 26, 26) {real, imag} */,
  {32'hbf16d020, 32'h3e5a20bc} /* (25, 26, 25) {real, imag} */,
  {32'h3f08e4c9, 32'hbe8a2690} /* (25, 26, 24) {real, imag} */,
  {32'h3e95293a, 32'hbd51856e} /* (25, 26, 23) {real, imag} */,
  {32'h3f0a54e5, 32'hbe4cf76c} /* (25, 26, 22) {real, imag} */,
  {32'hbe528e72, 32'h3dbeab44} /* (25, 26, 21) {real, imag} */,
  {32'hbcc89ac8, 32'hbd20caa0} /* (25, 26, 20) {real, imag} */,
  {32'h3ed8a848, 32'h3e7042f2} /* (25, 26, 19) {real, imag} */,
  {32'hbe5180a6, 32'hbdee0796} /* (25, 26, 18) {real, imag} */,
  {32'hbc000178, 32'hbece1e4e} /* (25, 26, 17) {real, imag} */,
  {32'h3efb1526, 32'hbc79ddf0} /* (25, 26, 16) {real, imag} */,
  {32'h3e1b5be2, 32'h3d829d40} /* (25, 26, 15) {real, imag} */,
  {32'hbe617fd8, 32'hbc917988} /* (25, 26, 14) {real, imag} */,
  {32'hbe525501, 32'h3e24ee69} /* (25, 26, 13) {real, imag} */,
  {32'h3ea6afd0, 32'h3db3dab0} /* (25, 26, 12) {real, imag} */,
  {32'h3e151cbb, 32'h3e212a8a} /* (25, 26, 11) {real, imag} */,
  {32'h3e25008c, 32'hbeb060ff} /* (25, 26, 10) {real, imag} */,
  {32'h3e67204d, 32'hbf041b3f} /* (25, 26, 9) {real, imag} */,
  {32'h3e14aca2, 32'h3e233576} /* (25, 26, 8) {real, imag} */,
  {32'hbe26f290, 32'hbe983f23} /* (25, 26, 7) {real, imag} */,
  {32'hbe2827f4, 32'hbf79ee26} /* (25, 26, 6) {real, imag} */,
  {32'hbe2ad513, 32'h3ec1be39} /* (25, 26, 5) {real, imag} */,
  {32'h3f4482ea, 32'h3f3cf13c} /* (25, 26, 4) {real, imag} */,
  {32'hbe7522e7, 32'hbdfe53f2} /* (25, 26, 3) {real, imag} */,
  {32'hbef89a47, 32'hbee784f3} /* (25, 26, 2) {real, imag} */,
  {32'h3ea161d2, 32'h3ec95ee7} /* (25, 26, 1) {real, imag} */,
  {32'h3d89d972, 32'hbcd20d00} /* (25, 26, 0) {real, imag} */,
  {32'hbf5708f7, 32'h3f20f6b1} /* (25, 25, 31) {real, imag} */,
  {32'h3d8180a4, 32'hbf514108} /* (25, 25, 30) {real, imag} */,
  {32'h3e7e936a, 32'hbf5584cc} /* (25, 25, 29) {real, imag} */,
  {32'h3f22fe4c, 32'h3f3202f3} /* (25, 25, 28) {real, imag} */,
  {32'hbf0c5bf6, 32'hbed28bfe} /* (25, 25, 27) {real, imag} */,
  {32'hbec5a902, 32'h3c27a840} /* (25, 25, 26) {real, imag} */,
  {32'h3dd22f0c, 32'h3ec0a940} /* (25, 25, 25) {real, imag} */,
  {32'h3e1f565b, 32'hbe74d1f4} /* (25, 25, 24) {real, imag} */,
  {32'hbe1ce534, 32'h3eb50910} /* (25, 25, 23) {real, imag} */,
  {32'hbf32401c, 32'h3ed68c1b} /* (25, 25, 22) {real, imag} */,
  {32'h3e5e08b8, 32'h3eb76f92} /* (25, 25, 21) {real, imag} */,
  {32'hbe11ff30, 32'hbedac813} /* (25, 25, 20) {real, imag} */,
  {32'h3f04969e, 32'hbeac9750} /* (25, 25, 19) {real, imag} */,
  {32'hbca0a488, 32'h3dce5f6d} /* (25, 25, 18) {real, imag} */,
  {32'hbe54377c, 32'hbe52e07a} /* (25, 25, 17) {real, imag} */,
  {32'hbdad7ade, 32'hbd627d44} /* (25, 25, 16) {real, imag} */,
  {32'h3dd2ab41, 32'hbea081d8} /* (25, 25, 15) {real, imag} */,
  {32'h3e343fe1, 32'h3e745803} /* (25, 25, 14) {real, imag} */,
  {32'hbedda76d, 32'h3ef15148} /* (25, 25, 13) {real, imag} */,
  {32'hbc1a2168, 32'hbdecdbb9} /* (25, 25, 12) {real, imag} */,
  {32'hbde62472, 32'h3ef2fa71} /* (25, 25, 11) {real, imag} */,
  {32'hbec378fe, 32'hbe023dcc} /* (25, 25, 10) {real, imag} */,
  {32'h3e587688, 32'hbead5b1f} /* (25, 25, 9) {real, imag} */,
  {32'h3db0ec86, 32'h3f849174} /* (25, 25, 8) {real, imag} */,
  {32'h3e582542, 32'h3eb27b17} /* (25, 25, 7) {real, imag} */,
  {32'hbe984002, 32'h3ea415e0} /* (25, 25, 6) {real, imag} */,
  {32'h3ce9e68c, 32'hbe34e45e} /* (25, 25, 5) {real, imag} */,
  {32'hbe9fbb24, 32'hbe48adcc} /* (25, 25, 4) {real, imag} */,
  {32'hbdfe4b14, 32'h3f3347a6} /* (25, 25, 3) {real, imag} */,
  {32'h3e2f3e3c, 32'h3e7aa3a0} /* (25, 25, 2) {real, imag} */,
  {32'hbf0ad48b, 32'h3eb54daa} /* (25, 25, 1) {real, imag} */,
  {32'hbf83d5fe, 32'h3da9c4ca} /* (25, 25, 0) {real, imag} */,
  {32'h3fb3094d, 32'hbecf4c7a} /* (25, 24, 31) {real, imag} */,
  {32'hbf739902, 32'h3e883a64} /* (25, 24, 30) {real, imag} */,
  {32'hbf5ff362, 32'hbe9297d6} /* (25, 24, 29) {real, imag} */,
  {32'hbe75d92a, 32'hbf6e730f} /* (25, 24, 28) {real, imag} */,
  {32'hbd1c7080, 32'hbd75b8fc} /* (25, 24, 27) {real, imag} */,
  {32'hbef54518, 32'h3e42cf94} /* (25, 24, 26) {real, imag} */,
  {32'hbdad0482, 32'h3ece6344} /* (25, 24, 25) {real, imag} */,
  {32'hbe2e9970, 32'h3f189e30} /* (25, 24, 24) {real, imag} */,
  {32'h3e1e7b40, 32'hbd9a89b4} /* (25, 24, 23) {real, imag} */,
  {32'h3e9aab6a, 32'hbde98a8a} /* (25, 24, 22) {real, imag} */,
  {32'h3ebd8652, 32'h3ea9b408} /* (25, 24, 21) {real, imag} */,
  {32'hbecd2d90, 32'hbeb43660} /* (25, 24, 20) {real, imag} */,
  {32'h3d4591d8, 32'h3f1cc25b} /* (25, 24, 19) {real, imag} */,
  {32'h3dd383a8, 32'h3f0d106b} /* (25, 24, 18) {real, imag} */,
  {32'h3e7d077a, 32'hbef7d72c} /* (25, 24, 17) {real, imag} */,
  {32'h3ea9fbac, 32'h3e8bc557} /* (25, 24, 16) {real, imag} */,
  {32'hbe195df7, 32'h3d9e6d7a} /* (25, 24, 15) {real, imag} */,
  {32'hbed6d18a, 32'hbe24b51e} /* (25, 24, 14) {real, imag} */,
  {32'hbe74286e, 32'hbe800618} /* (25, 24, 13) {real, imag} */,
  {32'h3c5fb9a8, 32'hbe8a896a} /* (25, 24, 12) {real, imag} */,
  {32'hbdc136c6, 32'h3e94641c} /* (25, 24, 11) {real, imag} */,
  {32'h3e38494c, 32'h3df17172} /* (25, 24, 10) {real, imag} */,
  {32'h3f1a0ad0, 32'h3f0a2d84} /* (25, 24, 9) {real, imag} */,
  {32'h3e6836ea, 32'h3d101770} /* (25, 24, 8) {real, imag} */,
  {32'h3f29f621, 32'h3de67b06} /* (25, 24, 7) {real, imag} */,
  {32'hbbd4f1a0, 32'h3d4c1ee8} /* (25, 24, 6) {real, imag} */,
  {32'hbef33594, 32'hbd257604} /* (25, 24, 5) {real, imag} */,
  {32'hbdcf6da0, 32'h3d494e4c} /* (25, 24, 4) {real, imag} */,
  {32'h3f12d514, 32'hbdcf0906} /* (25, 24, 3) {real, imag} */,
  {32'hbf170cdf, 32'hbe98abe0} /* (25, 24, 2) {real, imag} */,
  {32'h3fc9ab45, 32'hbed213d0} /* (25, 24, 1) {real, imag} */,
  {32'h3efdf5fa, 32'hbdfe68ee} /* (25, 24, 0) {real, imag} */,
  {32'hbe533190, 32'h3f03e02d} /* (25, 23, 31) {real, imag} */,
  {32'h3dd3a19e, 32'h3e91e0a8} /* (25, 23, 30) {real, imag} */,
  {32'h3d5ddd02, 32'h3f3c249c} /* (25, 23, 29) {real, imag} */,
  {32'hbe92c907, 32'h3ed0214c} /* (25, 23, 28) {real, imag} */,
  {32'hbda9d784, 32'hbf113a2c} /* (25, 23, 27) {real, imag} */,
  {32'h3f2ac6b4, 32'hbdb7de98} /* (25, 23, 26) {real, imag} */,
  {32'hbdf42fda, 32'h3eacaaec} /* (25, 23, 25) {real, imag} */,
  {32'h3ec2affe, 32'h3e72ef23} /* (25, 23, 24) {real, imag} */,
  {32'hbe40a2df, 32'hbd4fef68} /* (25, 23, 23) {real, imag} */,
  {32'hbe863128, 32'h3da739f4} /* (25, 23, 22) {real, imag} */,
  {32'hbe01ad3c, 32'hbeee45a4} /* (25, 23, 21) {real, imag} */,
  {32'hbe79a1a6, 32'hbdbb3bba} /* (25, 23, 20) {real, imag} */,
  {32'hbed747d5, 32'hbe4b3a78} /* (25, 23, 19) {real, imag} */,
  {32'h3e92ffa8, 32'h3cffacc4} /* (25, 23, 18) {real, imag} */,
  {32'hbe2d79e2, 32'h3e6a9c48} /* (25, 23, 17) {real, imag} */,
  {32'h3d3790d9, 32'hbc9ef7a8} /* (25, 23, 16) {real, imag} */,
  {32'hbe6928b7, 32'hbeff7810} /* (25, 23, 15) {real, imag} */,
  {32'hbe2bb44e, 32'hbcc55a28} /* (25, 23, 14) {real, imag} */,
  {32'h3e510ebc, 32'hbe84d225} /* (25, 23, 13) {real, imag} */,
  {32'h3ed7b1c0, 32'hbe876b61} /* (25, 23, 12) {real, imag} */,
  {32'h3ed7b435, 32'hbd49b99e} /* (25, 23, 11) {real, imag} */,
  {32'hbe633bbe, 32'h3d4171ec} /* (25, 23, 10) {real, imag} */,
  {32'h3ebdbab7, 32'hbedbd3b3} /* (25, 23, 9) {real, imag} */,
  {32'h3ea2a3cc, 32'h3ca92728} /* (25, 23, 8) {real, imag} */,
  {32'h3d44f110, 32'h3e812b9a} /* (25, 23, 7) {real, imag} */,
  {32'hbf318670, 32'h3e79ba44} /* (25, 23, 6) {real, imag} */,
  {32'h3f2550b6, 32'hbeb17aed} /* (25, 23, 5) {real, imag} */,
  {32'hbe84af65, 32'h3e2da943} /* (25, 23, 4) {real, imag} */,
  {32'h3eebdb40, 32'hbe220095} /* (25, 23, 3) {real, imag} */,
  {32'hbe281d80, 32'hbe1aaea2} /* (25, 23, 2) {real, imag} */,
  {32'h3ee9b67c, 32'h3e926a5e} /* (25, 23, 1) {real, imag} */,
  {32'hbf20a077, 32'h3e00c449} /* (25, 23, 0) {real, imag} */,
  {32'h3de8e4d0, 32'h3f31cc26} /* (25, 22, 31) {real, imag} */,
  {32'hbf031662, 32'h3ddefbe2} /* (25, 22, 30) {real, imag} */,
  {32'h3ec3f4f0, 32'hbec022e4} /* (25, 22, 29) {real, imag} */,
  {32'h3dbc37fb, 32'h3f0996aa} /* (25, 22, 28) {real, imag} */,
  {32'hbe834ea6, 32'hbf1342b2} /* (25, 22, 27) {real, imag} */,
  {32'h3e67ffde, 32'h3ddb69ea} /* (25, 22, 26) {real, imag} */,
  {32'h3e8bb1b5, 32'h3d7c65c4} /* (25, 22, 25) {real, imag} */,
  {32'h3eac89a0, 32'h3e4682a1} /* (25, 22, 24) {real, imag} */,
  {32'h3eb2273e, 32'hbe2fc0b5} /* (25, 22, 23) {real, imag} */,
  {32'hbdba60c6, 32'hbe1c273f} /* (25, 22, 22) {real, imag} */,
  {32'h3c0399f8, 32'h3ea21763} /* (25, 22, 21) {real, imag} */,
  {32'hbed0a59a, 32'h3f0bc40f} /* (25, 22, 20) {real, imag} */,
  {32'h3d7c87ec, 32'h3f2cf721} /* (25, 22, 19) {real, imag} */,
  {32'hbe9451c1, 32'hbead13b5} /* (25, 22, 18) {real, imag} */,
  {32'hbc385f72, 32'h3e1e581e} /* (25, 22, 17) {real, imag} */,
  {32'hbe1873c9, 32'hbe9087e1} /* (25, 22, 16) {real, imag} */,
  {32'h3e29db15, 32'hbe90168c} /* (25, 22, 15) {real, imag} */,
  {32'h3ed6773b, 32'hbef1ac66} /* (25, 22, 14) {real, imag} */,
  {32'h3de5bfd2, 32'hbdcf5b94} /* (25, 22, 13) {real, imag} */,
  {32'h3d3418e0, 32'h3c333c70} /* (25, 22, 12) {real, imag} */,
  {32'hbd2cd130, 32'h3d6014a0} /* (25, 22, 11) {real, imag} */,
  {32'h3ee4a091, 32'hbeef449a} /* (25, 22, 10) {real, imag} */,
  {32'h3f0d794f, 32'h3ee5bb35} /* (25, 22, 9) {real, imag} */,
  {32'hbf3d6904, 32'h3d88373d} /* (25, 22, 8) {real, imag} */,
  {32'h3ebd357a, 32'hbddf23e2} /* (25, 22, 7) {real, imag} */,
  {32'hbeaca2f7, 32'h3e9d6012} /* (25, 22, 6) {real, imag} */,
  {32'h3e92f74a, 32'h3eab7c2d} /* (25, 22, 5) {real, imag} */,
  {32'hbe2ccca0, 32'h3e300e5c} /* (25, 22, 4) {real, imag} */,
  {32'hbe621b00, 32'h3e831b2d} /* (25, 22, 3) {real, imag} */,
  {32'h3ebece1c, 32'hbf33439e} /* (25, 22, 2) {real, imag} */,
  {32'hbd3efed0, 32'h3ecb8bde} /* (25, 22, 1) {real, imag} */,
  {32'h3e922290, 32'h3e291a48} /* (25, 22, 0) {real, imag} */,
  {32'h3ecc079a, 32'hbe85b702} /* (25, 21, 31) {real, imag} */,
  {32'hbde9898a, 32'h3f12a943} /* (25, 21, 30) {real, imag} */,
  {32'h3e5f8e7d, 32'h3e97befa} /* (25, 21, 29) {real, imag} */,
  {32'h3e4d3f70, 32'hbf2a1eb6} /* (25, 21, 28) {real, imag} */,
  {32'h3e3966d0, 32'hbd908cf2} /* (25, 21, 27) {real, imag} */,
  {32'hbd8b932a, 32'h3ea8040f} /* (25, 21, 26) {real, imag} */,
  {32'hbe7c8673, 32'h3c445fa0} /* (25, 21, 25) {real, imag} */,
  {32'h3e6483ee, 32'hbe2a05ba} /* (25, 21, 24) {real, imag} */,
  {32'hbe8e420a, 32'h3e35bd45} /* (25, 21, 23) {real, imag} */,
  {32'hbe8d809c, 32'hbd301eb8} /* (25, 21, 22) {real, imag} */,
  {32'h3f2afa01, 32'hbe4c6831} /* (25, 21, 21) {real, imag} */,
  {32'h3eb20440, 32'h3d17d278} /* (25, 21, 20) {real, imag} */,
  {32'hbe60986c, 32'h3e36cf51} /* (25, 21, 19) {real, imag} */,
  {32'h3dcf0028, 32'h3e74c5d4} /* (25, 21, 18) {real, imag} */,
  {32'hbe5182a8, 32'h3d1758b4} /* (25, 21, 17) {real, imag} */,
  {32'h3d0b2e0c, 32'h3dfa8964} /* (25, 21, 16) {real, imag} */,
  {32'hbd6b65e4, 32'h3de2fe4a} /* (25, 21, 15) {real, imag} */,
  {32'h3e237ab6, 32'hbef88787} /* (25, 21, 14) {real, imag} */,
  {32'h3e76fae2, 32'h3e6dea47} /* (25, 21, 13) {real, imag} */,
  {32'h3cbc1a70, 32'h3d6b1292} /* (25, 21, 12) {real, imag} */,
  {32'hbef25a01, 32'hbc32cb30} /* (25, 21, 11) {real, imag} */,
  {32'hbea073df, 32'hbf1aa84a} /* (25, 21, 10) {real, imag} */,
  {32'hbe351fde, 32'h3d3a5b38} /* (25, 21, 9) {real, imag} */,
  {32'h3efd159b, 32'hbeebdcee} /* (25, 21, 8) {real, imag} */,
  {32'h3e99293c, 32'hbb1ff450} /* (25, 21, 7) {real, imag} */,
  {32'hbde742dd, 32'hbe1c8d6b} /* (25, 21, 6) {real, imag} */,
  {32'hbeef310f, 32'h3e40eec4} /* (25, 21, 5) {real, imag} */,
  {32'h3d122b7c, 32'h3cba48a0} /* (25, 21, 4) {real, imag} */,
  {32'h3ec5181c, 32'h3e37cff4} /* (25, 21, 3) {real, imag} */,
  {32'hbe71983e, 32'h3f41dd03} /* (25, 21, 2) {real, imag} */,
  {32'h3f1d9d56, 32'hbe4f2a3a} /* (25, 21, 1) {real, imag} */,
  {32'hbd2aafa8, 32'hbf19c7ce} /* (25, 21, 0) {real, imag} */,
  {32'h3eab1cef, 32'hbd5a24b2} /* (25, 20, 31) {real, imag} */,
  {32'h3f0c0c6e, 32'hbda22958} /* (25, 20, 30) {real, imag} */,
  {32'hbe2d9835, 32'h3e2cce55} /* (25, 20, 29) {real, imag} */,
  {32'hbe0998f7, 32'hbead6d65} /* (25, 20, 28) {real, imag} */,
  {32'hbf08a032, 32'hbdae0780} /* (25, 20, 27) {real, imag} */,
  {32'hbe50c6fa, 32'hbd65dc40} /* (25, 20, 26) {real, imag} */,
  {32'h3da46c70, 32'h3d7d2e80} /* (25, 20, 25) {real, imag} */,
  {32'hbee7e9c6, 32'hbea7a1c8} /* (25, 20, 24) {real, imag} */,
  {32'hbe9d7e38, 32'h3f1e1bb4} /* (25, 20, 23) {real, imag} */,
  {32'h3bb1d5a0, 32'h3e4a8346} /* (25, 20, 22) {real, imag} */,
  {32'hbe6fda4e, 32'hbe6e98b6} /* (25, 20, 21) {real, imag} */,
  {32'h3ef449a3, 32'hbdd70608} /* (25, 20, 20) {real, imag} */,
  {32'hbea78d47, 32'h3eb105ef} /* (25, 20, 19) {real, imag} */,
  {32'h3eaffccd, 32'h3d4191f4} /* (25, 20, 18) {real, imag} */,
  {32'h3ed75087, 32'hbf21c4cc} /* (25, 20, 17) {real, imag} */,
  {32'hbdeda0d9, 32'hbecc3502} /* (25, 20, 16) {real, imag} */,
  {32'h3e94f071, 32'hbeabf2d4} /* (25, 20, 15) {real, imag} */,
  {32'h3c9f7fb8, 32'h3e706742} /* (25, 20, 14) {real, imag} */,
  {32'h3f09b32d, 32'h3d3cb7fc} /* (25, 20, 13) {real, imag} */,
  {32'hbe8067a2, 32'h3ddf0a12} /* (25, 20, 12) {real, imag} */,
  {32'hbec3b987, 32'hbe50aeb2} /* (25, 20, 11) {real, imag} */,
  {32'h3eab4d47, 32'hbe29c37c} /* (25, 20, 10) {real, imag} */,
  {32'h3f1ea32f, 32'hbe6eff41} /* (25, 20, 9) {real, imag} */,
  {32'h3f0af56f, 32'h3d85e7b9} /* (25, 20, 8) {real, imag} */,
  {32'h3e860159, 32'hbe1f15c4} /* (25, 20, 7) {real, imag} */,
  {32'h3e3ac52a, 32'hbec254f3} /* (25, 20, 6) {real, imag} */,
  {32'h3f1b422c, 32'h3e20b1bf} /* (25, 20, 5) {real, imag} */,
  {32'h3c273450, 32'h3ed17c7a} /* (25, 20, 4) {real, imag} */,
  {32'hbf07dcf2, 32'h3eb64248} /* (25, 20, 3) {real, imag} */,
  {32'hbe2b25fe, 32'hbe28e3ac} /* (25, 20, 2) {real, imag} */,
  {32'hbe39d765, 32'h3da7b078} /* (25, 20, 1) {real, imag} */,
  {32'h3e890201, 32'h3e4060c6} /* (25, 20, 0) {real, imag} */,
  {32'hbf150b53, 32'hbe97c71a} /* (25, 19, 31) {real, imag} */,
  {32'hbe66c07d, 32'hbe822e14} /* (25, 19, 30) {real, imag} */,
  {32'h3e5f3386, 32'hbea0a616} /* (25, 19, 29) {real, imag} */,
  {32'hbe46f82a, 32'hbdbdb487} /* (25, 19, 28) {real, imag} */,
  {32'hbe44ddbb, 32'hbec521b4} /* (25, 19, 27) {real, imag} */,
  {32'h3d1342eb, 32'hbe592c34} /* (25, 19, 26) {real, imag} */,
  {32'h3e728d39, 32'hbe97c3c9} /* (25, 19, 25) {real, imag} */,
  {32'h3e94ef65, 32'h3d387d64} /* (25, 19, 24) {real, imag} */,
  {32'hbe7044ca, 32'hbe4e8fd1} /* (25, 19, 23) {real, imag} */,
  {32'h3cb6d9e0, 32'hbe670eec} /* (25, 19, 22) {real, imag} */,
  {32'hbe95ba59, 32'h3e281f8c} /* (25, 19, 21) {real, imag} */,
  {32'h3e469097, 32'hbedcefdc} /* (25, 19, 20) {real, imag} */,
  {32'hbde135a6, 32'h3de0d2df} /* (25, 19, 19) {real, imag} */,
  {32'h3f23cc90, 32'h3da040ac} /* (25, 19, 18) {real, imag} */,
  {32'hbd762f48, 32'hbddfeff9} /* (25, 19, 17) {real, imag} */,
  {32'hbf062a87, 32'h3e45ccb6} /* (25, 19, 16) {real, imag} */,
  {32'h3eae70ed, 32'h3d807f52} /* (25, 19, 15) {real, imag} */,
  {32'h3e620a0a, 32'h3ec8ad99} /* (25, 19, 14) {real, imag} */,
  {32'h3c5e60c0, 32'hbda20898} /* (25, 19, 13) {real, imag} */,
  {32'hbdc5d75c, 32'h3ec7b3c2} /* (25, 19, 12) {real, imag} */,
  {32'hbee15d7d, 32'hbf172ed8} /* (25, 19, 11) {real, imag} */,
  {32'h3e387ae3, 32'hbf13ad19} /* (25, 19, 10) {real, imag} */,
  {32'hbeb68fe2, 32'h3e445710} /* (25, 19, 9) {real, imag} */,
  {32'hbb522040, 32'hbd1771c0} /* (25, 19, 8) {real, imag} */,
  {32'hbee00281, 32'h3d637da9} /* (25, 19, 7) {real, imag} */,
  {32'h3e92cef3, 32'hbebe07ea} /* (25, 19, 6) {real, imag} */,
  {32'h3dec640a, 32'h3e467d6e} /* (25, 19, 5) {real, imag} */,
  {32'hbbd40c20, 32'hbe08cfa4} /* (25, 19, 4) {real, imag} */,
  {32'h3de3864f, 32'h3eeeccf5} /* (25, 19, 3) {real, imag} */,
  {32'h3d5c20b4, 32'h3ec10978} /* (25, 19, 2) {real, imag} */,
  {32'hbeaeb6ef, 32'h3d798054} /* (25, 19, 1) {real, imag} */,
  {32'hbe362b90, 32'h3ea7397e} /* (25, 19, 0) {real, imag} */,
  {32'hbdd18b5f, 32'hbf132681} /* (25, 18, 31) {real, imag} */,
  {32'h3ee0ff0a, 32'h3e85905a} /* (25, 18, 30) {real, imag} */,
  {32'hbdbf135b, 32'hbe2d08d8} /* (25, 18, 29) {real, imag} */,
  {32'hbdb1aace, 32'hbeae7b2e} /* (25, 18, 28) {real, imag} */,
  {32'h3f05f016, 32'hbde469fe} /* (25, 18, 27) {real, imag} */,
  {32'h3ee79860, 32'hbe5ab92f} /* (25, 18, 26) {real, imag} */,
  {32'hbea2a343, 32'h3c5d65c2} /* (25, 18, 25) {real, imag} */,
  {32'h3efaadd8, 32'hbd73837c} /* (25, 18, 24) {real, imag} */,
  {32'h3ebd7af6, 32'hbe4e879d} /* (25, 18, 23) {real, imag} */,
  {32'h3e6200aa, 32'hbebbd6ed} /* (25, 18, 22) {real, imag} */,
  {32'h3e0cc244, 32'hbdf48534} /* (25, 18, 21) {real, imag} */,
  {32'h3dc6891a, 32'h3eaafca9} /* (25, 18, 20) {real, imag} */,
  {32'h3e4187b2, 32'h3eba611e} /* (25, 18, 19) {real, imag} */,
  {32'h3dc0642c, 32'h3d351e48} /* (25, 18, 18) {real, imag} */,
  {32'h3c4677e0, 32'hbc1b29fc} /* (25, 18, 17) {real, imag} */,
  {32'h3d9c77f0, 32'hbc45eee0} /* (25, 18, 16) {real, imag} */,
  {32'h3dc50272, 32'h3e2390cf} /* (25, 18, 15) {real, imag} */,
  {32'h3e191a0a, 32'hbe6fd804} /* (25, 18, 14) {real, imag} */,
  {32'hbee12b79, 32'h3e26d64b} /* (25, 18, 13) {real, imag} */,
  {32'hbf02d1d0, 32'hbe429d54} /* (25, 18, 12) {real, imag} */,
  {32'h3e5c8888, 32'hbddd2e98} /* (25, 18, 11) {real, imag} */,
  {32'h3ef673a9, 32'h3df0cfa2} /* (25, 18, 10) {real, imag} */,
  {32'hbefe280a, 32'h3f2a4a28} /* (25, 18, 9) {real, imag} */,
  {32'hbe9d24a9, 32'hbec68f3e} /* (25, 18, 8) {real, imag} */,
  {32'hbf7bcbc4, 32'hbea0a711} /* (25, 18, 7) {real, imag} */,
  {32'hbd75f708, 32'h3e54fdcb} /* (25, 18, 6) {real, imag} */,
  {32'h3e5eb84c, 32'hbea122a4} /* (25, 18, 5) {real, imag} */,
  {32'h3f02ba72, 32'h3ea67177} /* (25, 18, 4) {real, imag} */,
  {32'hbe58397a, 32'hbe5f44ce} /* (25, 18, 3) {real, imag} */,
  {32'hbc184c38, 32'hbddbd707} /* (25, 18, 2) {real, imag} */,
  {32'h3de6c5ee, 32'hbf2df588} /* (25, 18, 1) {real, imag} */,
  {32'hbe435684, 32'hbf302eb2} /* (25, 18, 0) {real, imag} */,
  {32'hbe46f8d6, 32'h3d5d3a00} /* (25, 17, 31) {real, imag} */,
  {32'hbd715749, 32'hbf220e93} /* (25, 17, 30) {real, imag} */,
  {32'hbcb3ccf4, 32'h3e2b5640} /* (25, 17, 29) {real, imag} */,
  {32'hbe272e3e, 32'hbd8c06ba} /* (25, 17, 28) {real, imag} */,
  {32'hbe0f430e, 32'h3ecf686c} /* (25, 17, 27) {real, imag} */,
  {32'hbd8613d7, 32'hbe2e916a} /* (25, 17, 26) {real, imag} */,
  {32'h3e33e910, 32'h3e60b1c0} /* (25, 17, 25) {real, imag} */,
  {32'h3ec59995, 32'hbe341c65} /* (25, 17, 24) {real, imag} */,
  {32'h3cc57f8c, 32'h3e5c8569} /* (25, 17, 23) {real, imag} */,
  {32'h3e801151, 32'h3dbf5674} /* (25, 17, 22) {real, imag} */,
  {32'hbeb9e1aa, 32'h3e8c63d8} /* (25, 17, 21) {real, imag} */,
  {32'h3dd552f0, 32'h3e7ea7fc} /* (25, 17, 20) {real, imag} */,
  {32'hbd6d5b72, 32'hbe8fb30b} /* (25, 17, 19) {real, imag} */,
  {32'h3eee9a46, 32'h3ec14abc} /* (25, 17, 18) {real, imag} */,
  {32'h3e2a1482, 32'h3d0abe26} /* (25, 17, 17) {real, imag} */,
  {32'h3d3264dc, 32'h3e1d6b44} /* (25, 17, 16) {real, imag} */,
  {32'hbe96ac7a, 32'hbe94fbde} /* (25, 17, 15) {real, imag} */,
  {32'hbe95c3e4, 32'hbe5b70d0} /* (25, 17, 14) {real, imag} */,
  {32'h3e0d0f65, 32'hbdf1b0c5} /* (25, 17, 13) {real, imag} */,
  {32'h3e575a82, 32'h3e20c56e} /* (25, 17, 12) {real, imag} */,
  {32'h3e3fd4cc, 32'hbe538299} /* (25, 17, 11) {real, imag} */,
  {32'h3e0e87f4, 32'h3f237046} /* (25, 17, 10) {real, imag} */,
  {32'h3e6b9aa3, 32'hbdd0f03b} /* (25, 17, 9) {real, imag} */,
  {32'h3d032d3a, 32'hbd027390} /* (25, 17, 8) {real, imag} */,
  {32'hbe40d2e0, 32'h3f347ef0} /* (25, 17, 7) {real, imag} */,
  {32'h3e13d434, 32'hbe075b0d} /* (25, 17, 6) {real, imag} */,
  {32'hbe6740f8, 32'h3d17c9d0} /* (25, 17, 5) {real, imag} */,
  {32'h3cbe7a24, 32'h3cda9a2e} /* (25, 17, 4) {real, imag} */,
  {32'hbaea9f40, 32'hbdd93240} /* (25, 17, 3) {real, imag} */,
  {32'hbd08695c, 32'hbe3499cd} /* (25, 17, 2) {real, imag} */,
  {32'hbe981c16, 32'h3ee0ad96} /* (25, 17, 1) {real, imag} */,
  {32'h3f04a911, 32'hbd77fe70} /* (25, 17, 0) {real, imag} */,
  {32'h3e2f8c82, 32'h3e37c0fa} /* (25, 16, 31) {real, imag} */,
  {32'h3e02b66c, 32'hbcf5b7d4} /* (25, 16, 30) {real, imag} */,
  {32'hbe454254, 32'hbcf49246} /* (25, 16, 29) {real, imag} */,
  {32'h3e2ad96e, 32'h3ea87ee1} /* (25, 16, 28) {real, imag} */,
  {32'h3dbfbe34, 32'h3dbc30e2} /* (25, 16, 27) {real, imag} */,
  {32'h3ea35f08, 32'h3e83eb6c} /* (25, 16, 26) {real, imag} */,
  {32'hbe2e39b8, 32'hbe4b99ce} /* (25, 16, 25) {real, imag} */,
  {32'hbe46da56, 32'h3d6fcd16} /* (25, 16, 24) {real, imag} */,
  {32'hbedf2bba, 32'hbcedff00} /* (25, 16, 23) {real, imag} */,
  {32'hbdab4bee, 32'hbe1ad0b5} /* (25, 16, 22) {real, imag} */,
  {32'hbd26ddd2, 32'h3e629ec8} /* (25, 16, 21) {real, imag} */,
  {32'h3c803798, 32'h3ee70a12} /* (25, 16, 20) {real, imag} */,
  {32'hbe95297a, 32'h3bf9b650} /* (25, 16, 19) {real, imag} */,
  {32'hbe01a8fe, 32'h3c83c3e7} /* (25, 16, 18) {real, imag} */,
  {32'hbdc67dd8, 32'hbe4cec62} /* (25, 16, 17) {real, imag} */,
  {32'h3cb443c8, 32'h00000000} /* (25, 16, 16) {real, imag} */,
  {32'hbdc67dd8, 32'h3e4cec62} /* (25, 16, 15) {real, imag} */,
  {32'hbe01a8fe, 32'hbc83c3e7} /* (25, 16, 14) {real, imag} */,
  {32'hbe95297a, 32'hbbf9b650} /* (25, 16, 13) {real, imag} */,
  {32'h3c803798, 32'hbee70a12} /* (25, 16, 12) {real, imag} */,
  {32'hbd26ddd2, 32'hbe629ec8} /* (25, 16, 11) {real, imag} */,
  {32'hbdab4bee, 32'h3e1ad0b5} /* (25, 16, 10) {real, imag} */,
  {32'hbedf2bba, 32'h3cedff00} /* (25, 16, 9) {real, imag} */,
  {32'hbe46da56, 32'hbd6fcd16} /* (25, 16, 8) {real, imag} */,
  {32'hbe2e39b8, 32'h3e4b99ce} /* (25, 16, 7) {real, imag} */,
  {32'h3ea35f08, 32'hbe83eb6c} /* (25, 16, 6) {real, imag} */,
  {32'h3dbfbe34, 32'hbdbc30e2} /* (25, 16, 5) {real, imag} */,
  {32'h3e2ad96e, 32'hbea87ee1} /* (25, 16, 4) {real, imag} */,
  {32'hbe454254, 32'h3cf49246} /* (25, 16, 3) {real, imag} */,
  {32'h3e02b66c, 32'h3cf5b7d4} /* (25, 16, 2) {real, imag} */,
  {32'h3e2f8c82, 32'hbe37c0fa} /* (25, 16, 1) {real, imag} */,
  {32'h3ed64851, 32'h00000000} /* (25, 16, 0) {real, imag} */,
  {32'hbe981c16, 32'hbee0ad96} /* (25, 15, 31) {real, imag} */,
  {32'hbd08695c, 32'h3e3499cd} /* (25, 15, 30) {real, imag} */,
  {32'hbaea9f40, 32'h3dd93240} /* (25, 15, 29) {real, imag} */,
  {32'h3cbe7a24, 32'hbcda9a2e} /* (25, 15, 28) {real, imag} */,
  {32'hbe6740f8, 32'hbd17c9d0} /* (25, 15, 27) {real, imag} */,
  {32'h3e13d434, 32'h3e075b0d} /* (25, 15, 26) {real, imag} */,
  {32'hbe40d2e0, 32'hbf347ef0} /* (25, 15, 25) {real, imag} */,
  {32'h3d032d3a, 32'h3d027390} /* (25, 15, 24) {real, imag} */,
  {32'h3e6b9aa3, 32'h3dd0f03b} /* (25, 15, 23) {real, imag} */,
  {32'h3e0e87f4, 32'hbf237046} /* (25, 15, 22) {real, imag} */,
  {32'h3e3fd4cc, 32'h3e538299} /* (25, 15, 21) {real, imag} */,
  {32'h3e575a82, 32'hbe20c56e} /* (25, 15, 20) {real, imag} */,
  {32'h3e0d0f65, 32'h3df1b0c5} /* (25, 15, 19) {real, imag} */,
  {32'hbe95c3e4, 32'h3e5b70d0} /* (25, 15, 18) {real, imag} */,
  {32'hbe96ac7a, 32'h3e94fbde} /* (25, 15, 17) {real, imag} */,
  {32'h3d3264dc, 32'hbe1d6b44} /* (25, 15, 16) {real, imag} */,
  {32'h3e2a1482, 32'hbd0abe26} /* (25, 15, 15) {real, imag} */,
  {32'h3eee9a46, 32'hbec14abc} /* (25, 15, 14) {real, imag} */,
  {32'hbd6d5b72, 32'h3e8fb30b} /* (25, 15, 13) {real, imag} */,
  {32'h3dd552f0, 32'hbe7ea7fc} /* (25, 15, 12) {real, imag} */,
  {32'hbeb9e1aa, 32'hbe8c63d8} /* (25, 15, 11) {real, imag} */,
  {32'h3e801151, 32'hbdbf5674} /* (25, 15, 10) {real, imag} */,
  {32'h3cc57f8c, 32'hbe5c8569} /* (25, 15, 9) {real, imag} */,
  {32'h3ec59995, 32'h3e341c65} /* (25, 15, 8) {real, imag} */,
  {32'h3e33e910, 32'hbe60b1c0} /* (25, 15, 7) {real, imag} */,
  {32'hbd8613d7, 32'h3e2e916a} /* (25, 15, 6) {real, imag} */,
  {32'hbe0f430e, 32'hbecf686c} /* (25, 15, 5) {real, imag} */,
  {32'hbe272e3e, 32'h3d8c06ba} /* (25, 15, 4) {real, imag} */,
  {32'hbcb3ccf4, 32'hbe2b5640} /* (25, 15, 3) {real, imag} */,
  {32'hbd715749, 32'h3f220e93} /* (25, 15, 2) {real, imag} */,
  {32'hbe46f8d6, 32'hbd5d3a00} /* (25, 15, 1) {real, imag} */,
  {32'h3f04a911, 32'h3d77fe70} /* (25, 15, 0) {real, imag} */,
  {32'h3de6c5ee, 32'h3f2df588} /* (25, 14, 31) {real, imag} */,
  {32'hbc184c38, 32'h3ddbd707} /* (25, 14, 30) {real, imag} */,
  {32'hbe58397a, 32'h3e5f44ce} /* (25, 14, 29) {real, imag} */,
  {32'h3f02ba72, 32'hbea67177} /* (25, 14, 28) {real, imag} */,
  {32'h3e5eb84c, 32'h3ea122a4} /* (25, 14, 27) {real, imag} */,
  {32'hbd75f708, 32'hbe54fdcb} /* (25, 14, 26) {real, imag} */,
  {32'hbf7bcbc4, 32'h3ea0a711} /* (25, 14, 25) {real, imag} */,
  {32'hbe9d24a9, 32'h3ec68f3e} /* (25, 14, 24) {real, imag} */,
  {32'hbefe280a, 32'hbf2a4a28} /* (25, 14, 23) {real, imag} */,
  {32'h3ef673a9, 32'hbdf0cfa2} /* (25, 14, 22) {real, imag} */,
  {32'h3e5c8888, 32'h3ddd2e98} /* (25, 14, 21) {real, imag} */,
  {32'hbf02d1d0, 32'h3e429d54} /* (25, 14, 20) {real, imag} */,
  {32'hbee12b79, 32'hbe26d64b} /* (25, 14, 19) {real, imag} */,
  {32'h3e191a0a, 32'h3e6fd804} /* (25, 14, 18) {real, imag} */,
  {32'h3dc50272, 32'hbe2390cf} /* (25, 14, 17) {real, imag} */,
  {32'h3d9c77f0, 32'h3c45eee0} /* (25, 14, 16) {real, imag} */,
  {32'h3c4677e0, 32'h3c1b29fc} /* (25, 14, 15) {real, imag} */,
  {32'h3dc0642c, 32'hbd351e48} /* (25, 14, 14) {real, imag} */,
  {32'h3e4187b2, 32'hbeba611e} /* (25, 14, 13) {real, imag} */,
  {32'h3dc6891a, 32'hbeaafca9} /* (25, 14, 12) {real, imag} */,
  {32'h3e0cc244, 32'h3df48534} /* (25, 14, 11) {real, imag} */,
  {32'h3e6200aa, 32'h3ebbd6ed} /* (25, 14, 10) {real, imag} */,
  {32'h3ebd7af6, 32'h3e4e879d} /* (25, 14, 9) {real, imag} */,
  {32'h3efaadd8, 32'h3d73837c} /* (25, 14, 8) {real, imag} */,
  {32'hbea2a343, 32'hbc5d65c2} /* (25, 14, 7) {real, imag} */,
  {32'h3ee79860, 32'h3e5ab92f} /* (25, 14, 6) {real, imag} */,
  {32'h3f05f016, 32'h3de469fe} /* (25, 14, 5) {real, imag} */,
  {32'hbdb1aace, 32'h3eae7b2e} /* (25, 14, 4) {real, imag} */,
  {32'hbdbf135b, 32'h3e2d08d8} /* (25, 14, 3) {real, imag} */,
  {32'h3ee0ff0a, 32'hbe85905a} /* (25, 14, 2) {real, imag} */,
  {32'hbdd18b5f, 32'h3f132681} /* (25, 14, 1) {real, imag} */,
  {32'hbe435684, 32'h3f302eb2} /* (25, 14, 0) {real, imag} */,
  {32'hbeaeb6ef, 32'hbd798054} /* (25, 13, 31) {real, imag} */,
  {32'h3d5c20b4, 32'hbec10978} /* (25, 13, 30) {real, imag} */,
  {32'h3de3864f, 32'hbeeeccf5} /* (25, 13, 29) {real, imag} */,
  {32'hbbd40c20, 32'h3e08cfa4} /* (25, 13, 28) {real, imag} */,
  {32'h3dec640a, 32'hbe467d6e} /* (25, 13, 27) {real, imag} */,
  {32'h3e92cef3, 32'h3ebe07ea} /* (25, 13, 26) {real, imag} */,
  {32'hbee00281, 32'hbd637da9} /* (25, 13, 25) {real, imag} */,
  {32'hbb522040, 32'h3d1771c0} /* (25, 13, 24) {real, imag} */,
  {32'hbeb68fe2, 32'hbe445710} /* (25, 13, 23) {real, imag} */,
  {32'h3e387ae3, 32'h3f13ad19} /* (25, 13, 22) {real, imag} */,
  {32'hbee15d7d, 32'h3f172ed8} /* (25, 13, 21) {real, imag} */,
  {32'hbdc5d75c, 32'hbec7b3c2} /* (25, 13, 20) {real, imag} */,
  {32'h3c5e60c0, 32'h3da20898} /* (25, 13, 19) {real, imag} */,
  {32'h3e620a0a, 32'hbec8ad99} /* (25, 13, 18) {real, imag} */,
  {32'h3eae70ed, 32'hbd807f52} /* (25, 13, 17) {real, imag} */,
  {32'hbf062a87, 32'hbe45ccb6} /* (25, 13, 16) {real, imag} */,
  {32'hbd762f48, 32'h3ddfeff9} /* (25, 13, 15) {real, imag} */,
  {32'h3f23cc90, 32'hbda040ac} /* (25, 13, 14) {real, imag} */,
  {32'hbde135a6, 32'hbde0d2df} /* (25, 13, 13) {real, imag} */,
  {32'h3e469097, 32'h3edcefdc} /* (25, 13, 12) {real, imag} */,
  {32'hbe95ba59, 32'hbe281f8c} /* (25, 13, 11) {real, imag} */,
  {32'h3cb6d9e0, 32'h3e670eec} /* (25, 13, 10) {real, imag} */,
  {32'hbe7044ca, 32'h3e4e8fd1} /* (25, 13, 9) {real, imag} */,
  {32'h3e94ef65, 32'hbd387d64} /* (25, 13, 8) {real, imag} */,
  {32'h3e728d39, 32'h3e97c3c9} /* (25, 13, 7) {real, imag} */,
  {32'h3d1342eb, 32'h3e592c34} /* (25, 13, 6) {real, imag} */,
  {32'hbe44ddbb, 32'h3ec521b4} /* (25, 13, 5) {real, imag} */,
  {32'hbe46f82a, 32'h3dbdb487} /* (25, 13, 4) {real, imag} */,
  {32'h3e5f3386, 32'h3ea0a616} /* (25, 13, 3) {real, imag} */,
  {32'hbe66c07d, 32'h3e822e14} /* (25, 13, 2) {real, imag} */,
  {32'hbf150b53, 32'h3e97c71a} /* (25, 13, 1) {real, imag} */,
  {32'hbe362b90, 32'hbea7397e} /* (25, 13, 0) {real, imag} */,
  {32'hbe39d765, 32'hbda7b078} /* (25, 12, 31) {real, imag} */,
  {32'hbe2b25fe, 32'h3e28e3ac} /* (25, 12, 30) {real, imag} */,
  {32'hbf07dcf2, 32'hbeb64248} /* (25, 12, 29) {real, imag} */,
  {32'h3c273450, 32'hbed17c7a} /* (25, 12, 28) {real, imag} */,
  {32'h3f1b422c, 32'hbe20b1bf} /* (25, 12, 27) {real, imag} */,
  {32'h3e3ac52a, 32'h3ec254f3} /* (25, 12, 26) {real, imag} */,
  {32'h3e860159, 32'h3e1f15c4} /* (25, 12, 25) {real, imag} */,
  {32'h3f0af56f, 32'hbd85e7b9} /* (25, 12, 24) {real, imag} */,
  {32'h3f1ea32f, 32'h3e6eff41} /* (25, 12, 23) {real, imag} */,
  {32'h3eab4d47, 32'h3e29c37c} /* (25, 12, 22) {real, imag} */,
  {32'hbec3b987, 32'h3e50aeb2} /* (25, 12, 21) {real, imag} */,
  {32'hbe8067a2, 32'hbddf0a12} /* (25, 12, 20) {real, imag} */,
  {32'h3f09b32d, 32'hbd3cb7fc} /* (25, 12, 19) {real, imag} */,
  {32'h3c9f7fb8, 32'hbe706742} /* (25, 12, 18) {real, imag} */,
  {32'h3e94f071, 32'h3eabf2d4} /* (25, 12, 17) {real, imag} */,
  {32'hbdeda0d9, 32'h3ecc3502} /* (25, 12, 16) {real, imag} */,
  {32'h3ed75087, 32'h3f21c4cc} /* (25, 12, 15) {real, imag} */,
  {32'h3eaffccd, 32'hbd4191f4} /* (25, 12, 14) {real, imag} */,
  {32'hbea78d47, 32'hbeb105ef} /* (25, 12, 13) {real, imag} */,
  {32'h3ef449a3, 32'h3dd70608} /* (25, 12, 12) {real, imag} */,
  {32'hbe6fda4e, 32'h3e6e98b6} /* (25, 12, 11) {real, imag} */,
  {32'h3bb1d5a0, 32'hbe4a8346} /* (25, 12, 10) {real, imag} */,
  {32'hbe9d7e38, 32'hbf1e1bb4} /* (25, 12, 9) {real, imag} */,
  {32'hbee7e9c6, 32'h3ea7a1c8} /* (25, 12, 8) {real, imag} */,
  {32'h3da46c70, 32'hbd7d2e80} /* (25, 12, 7) {real, imag} */,
  {32'hbe50c6fa, 32'h3d65dc40} /* (25, 12, 6) {real, imag} */,
  {32'hbf08a032, 32'h3dae0780} /* (25, 12, 5) {real, imag} */,
  {32'hbe0998f7, 32'h3ead6d65} /* (25, 12, 4) {real, imag} */,
  {32'hbe2d9835, 32'hbe2cce55} /* (25, 12, 3) {real, imag} */,
  {32'h3f0c0c6e, 32'h3da22958} /* (25, 12, 2) {real, imag} */,
  {32'h3eab1cef, 32'h3d5a24b2} /* (25, 12, 1) {real, imag} */,
  {32'h3e890201, 32'hbe4060c6} /* (25, 12, 0) {real, imag} */,
  {32'h3f1d9d56, 32'h3e4f2a3a} /* (25, 11, 31) {real, imag} */,
  {32'hbe71983e, 32'hbf41dd03} /* (25, 11, 30) {real, imag} */,
  {32'h3ec5181c, 32'hbe37cff4} /* (25, 11, 29) {real, imag} */,
  {32'h3d122b7c, 32'hbcba48a0} /* (25, 11, 28) {real, imag} */,
  {32'hbeef310f, 32'hbe40eec4} /* (25, 11, 27) {real, imag} */,
  {32'hbde742dd, 32'h3e1c8d6b} /* (25, 11, 26) {real, imag} */,
  {32'h3e99293c, 32'h3b1ff450} /* (25, 11, 25) {real, imag} */,
  {32'h3efd159b, 32'h3eebdcee} /* (25, 11, 24) {real, imag} */,
  {32'hbe351fde, 32'hbd3a5b38} /* (25, 11, 23) {real, imag} */,
  {32'hbea073df, 32'h3f1aa84a} /* (25, 11, 22) {real, imag} */,
  {32'hbef25a01, 32'h3c32cb30} /* (25, 11, 21) {real, imag} */,
  {32'h3cbc1a70, 32'hbd6b1292} /* (25, 11, 20) {real, imag} */,
  {32'h3e76fae2, 32'hbe6dea47} /* (25, 11, 19) {real, imag} */,
  {32'h3e237ab6, 32'h3ef88787} /* (25, 11, 18) {real, imag} */,
  {32'hbd6b65e4, 32'hbde2fe4a} /* (25, 11, 17) {real, imag} */,
  {32'h3d0b2e0c, 32'hbdfa8964} /* (25, 11, 16) {real, imag} */,
  {32'hbe5182a8, 32'hbd1758b4} /* (25, 11, 15) {real, imag} */,
  {32'h3dcf0028, 32'hbe74c5d4} /* (25, 11, 14) {real, imag} */,
  {32'hbe60986c, 32'hbe36cf51} /* (25, 11, 13) {real, imag} */,
  {32'h3eb20440, 32'hbd17d278} /* (25, 11, 12) {real, imag} */,
  {32'h3f2afa01, 32'h3e4c6831} /* (25, 11, 11) {real, imag} */,
  {32'hbe8d809c, 32'h3d301eb8} /* (25, 11, 10) {real, imag} */,
  {32'hbe8e420a, 32'hbe35bd45} /* (25, 11, 9) {real, imag} */,
  {32'h3e6483ee, 32'h3e2a05ba} /* (25, 11, 8) {real, imag} */,
  {32'hbe7c8673, 32'hbc445fa0} /* (25, 11, 7) {real, imag} */,
  {32'hbd8b932a, 32'hbea8040f} /* (25, 11, 6) {real, imag} */,
  {32'h3e3966d0, 32'h3d908cf2} /* (25, 11, 5) {real, imag} */,
  {32'h3e4d3f70, 32'h3f2a1eb6} /* (25, 11, 4) {real, imag} */,
  {32'h3e5f8e7d, 32'hbe97befa} /* (25, 11, 3) {real, imag} */,
  {32'hbde9898a, 32'hbf12a943} /* (25, 11, 2) {real, imag} */,
  {32'h3ecc079a, 32'h3e85b702} /* (25, 11, 1) {real, imag} */,
  {32'hbd2aafa8, 32'h3f19c7ce} /* (25, 11, 0) {real, imag} */,
  {32'hbd3efed0, 32'hbecb8bde} /* (25, 10, 31) {real, imag} */,
  {32'h3ebece1c, 32'h3f33439e} /* (25, 10, 30) {real, imag} */,
  {32'hbe621b00, 32'hbe831b2d} /* (25, 10, 29) {real, imag} */,
  {32'hbe2ccca0, 32'hbe300e5c} /* (25, 10, 28) {real, imag} */,
  {32'h3e92f74a, 32'hbeab7c2d} /* (25, 10, 27) {real, imag} */,
  {32'hbeaca2f7, 32'hbe9d6012} /* (25, 10, 26) {real, imag} */,
  {32'h3ebd357a, 32'h3ddf23e2} /* (25, 10, 25) {real, imag} */,
  {32'hbf3d6904, 32'hbd88373d} /* (25, 10, 24) {real, imag} */,
  {32'h3f0d794f, 32'hbee5bb35} /* (25, 10, 23) {real, imag} */,
  {32'h3ee4a091, 32'h3eef449a} /* (25, 10, 22) {real, imag} */,
  {32'hbd2cd130, 32'hbd6014a0} /* (25, 10, 21) {real, imag} */,
  {32'h3d3418e0, 32'hbc333c70} /* (25, 10, 20) {real, imag} */,
  {32'h3de5bfd2, 32'h3dcf5b94} /* (25, 10, 19) {real, imag} */,
  {32'h3ed6773b, 32'h3ef1ac66} /* (25, 10, 18) {real, imag} */,
  {32'h3e29db15, 32'h3e90168c} /* (25, 10, 17) {real, imag} */,
  {32'hbe1873c9, 32'h3e9087e1} /* (25, 10, 16) {real, imag} */,
  {32'hbc385f72, 32'hbe1e581e} /* (25, 10, 15) {real, imag} */,
  {32'hbe9451c1, 32'h3ead13b5} /* (25, 10, 14) {real, imag} */,
  {32'h3d7c87ec, 32'hbf2cf721} /* (25, 10, 13) {real, imag} */,
  {32'hbed0a59a, 32'hbf0bc40f} /* (25, 10, 12) {real, imag} */,
  {32'h3c0399f8, 32'hbea21763} /* (25, 10, 11) {real, imag} */,
  {32'hbdba60c6, 32'h3e1c273f} /* (25, 10, 10) {real, imag} */,
  {32'h3eb2273e, 32'h3e2fc0b5} /* (25, 10, 9) {real, imag} */,
  {32'h3eac89a0, 32'hbe4682a1} /* (25, 10, 8) {real, imag} */,
  {32'h3e8bb1b5, 32'hbd7c65c4} /* (25, 10, 7) {real, imag} */,
  {32'h3e67ffde, 32'hbddb69ea} /* (25, 10, 6) {real, imag} */,
  {32'hbe834ea6, 32'h3f1342b2} /* (25, 10, 5) {real, imag} */,
  {32'h3dbc37fb, 32'hbf0996aa} /* (25, 10, 4) {real, imag} */,
  {32'h3ec3f4f0, 32'h3ec022e4} /* (25, 10, 3) {real, imag} */,
  {32'hbf031662, 32'hbddefbe2} /* (25, 10, 2) {real, imag} */,
  {32'h3de8e4d0, 32'hbf31cc26} /* (25, 10, 1) {real, imag} */,
  {32'h3e922290, 32'hbe291a48} /* (25, 10, 0) {real, imag} */,
  {32'h3ee9b67c, 32'hbe926a5e} /* (25, 9, 31) {real, imag} */,
  {32'hbe281d80, 32'h3e1aaea2} /* (25, 9, 30) {real, imag} */,
  {32'h3eebdb40, 32'h3e220095} /* (25, 9, 29) {real, imag} */,
  {32'hbe84af65, 32'hbe2da943} /* (25, 9, 28) {real, imag} */,
  {32'h3f2550b6, 32'h3eb17aed} /* (25, 9, 27) {real, imag} */,
  {32'hbf318670, 32'hbe79ba44} /* (25, 9, 26) {real, imag} */,
  {32'h3d44f110, 32'hbe812b9a} /* (25, 9, 25) {real, imag} */,
  {32'h3ea2a3cc, 32'hbca92728} /* (25, 9, 24) {real, imag} */,
  {32'h3ebdbab7, 32'h3edbd3b3} /* (25, 9, 23) {real, imag} */,
  {32'hbe633bbe, 32'hbd4171ec} /* (25, 9, 22) {real, imag} */,
  {32'h3ed7b435, 32'h3d49b99e} /* (25, 9, 21) {real, imag} */,
  {32'h3ed7b1c0, 32'h3e876b61} /* (25, 9, 20) {real, imag} */,
  {32'h3e510ebc, 32'h3e84d225} /* (25, 9, 19) {real, imag} */,
  {32'hbe2bb44e, 32'h3cc55a28} /* (25, 9, 18) {real, imag} */,
  {32'hbe6928b7, 32'h3eff7810} /* (25, 9, 17) {real, imag} */,
  {32'h3d3790d9, 32'h3c9ef7a8} /* (25, 9, 16) {real, imag} */,
  {32'hbe2d79e2, 32'hbe6a9c48} /* (25, 9, 15) {real, imag} */,
  {32'h3e92ffa8, 32'hbcffacc4} /* (25, 9, 14) {real, imag} */,
  {32'hbed747d5, 32'h3e4b3a78} /* (25, 9, 13) {real, imag} */,
  {32'hbe79a1a6, 32'h3dbb3bba} /* (25, 9, 12) {real, imag} */,
  {32'hbe01ad3c, 32'h3eee45a4} /* (25, 9, 11) {real, imag} */,
  {32'hbe863128, 32'hbda739f4} /* (25, 9, 10) {real, imag} */,
  {32'hbe40a2df, 32'h3d4fef68} /* (25, 9, 9) {real, imag} */,
  {32'h3ec2affe, 32'hbe72ef23} /* (25, 9, 8) {real, imag} */,
  {32'hbdf42fda, 32'hbeacaaec} /* (25, 9, 7) {real, imag} */,
  {32'h3f2ac6b4, 32'h3db7de98} /* (25, 9, 6) {real, imag} */,
  {32'hbda9d784, 32'h3f113a2c} /* (25, 9, 5) {real, imag} */,
  {32'hbe92c907, 32'hbed0214c} /* (25, 9, 4) {real, imag} */,
  {32'h3d5ddd02, 32'hbf3c249c} /* (25, 9, 3) {real, imag} */,
  {32'h3dd3a19e, 32'hbe91e0a8} /* (25, 9, 2) {real, imag} */,
  {32'hbe533190, 32'hbf03e02d} /* (25, 9, 1) {real, imag} */,
  {32'hbf20a077, 32'hbe00c449} /* (25, 9, 0) {real, imag} */,
  {32'h3fc9ab45, 32'h3ed213d0} /* (25, 8, 31) {real, imag} */,
  {32'hbf170cdf, 32'h3e98abe0} /* (25, 8, 30) {real, imag} */,
  {32'h3f12d514, 32'h3dcf0906} /* (25, 8, 29) {real, imag} */,
  {32'hbdcf6da0, 32'hbd494e4c} /* (25, 8, 28) {real, imag} */,
  {32'hbef33594, 32'h3d257604} /* (25, 8, 27) {real, imag} */,
  {32'hbbd4f1a0, 32'hbd4c1ee8} /* (25, 8, 26) {real, imag} */,
  {32'h3f29f621, 32'hbde67b06} /* (25, 8, 25) {real, imag} */,
  {32'h3e6836ea, 32'hbd101770} /* (25, 8, 24) {real, imag} */,
  {32'h3f1a0ad0, 32'hbf0a2d84} /* (25, 8, 23) {real, imag} */,
  {32'h3e38494c, 32'hbdf17172} /* (25, 8, 22) {real, imag} */,
  {32'hbdc136c6, 32'hbe94641c} /* (25, 8, 21) {real, imag} */,
  {32'h3c5fb9a8, 32'h3e8a896a} /* (25, 8, 20) {real, imag} */,
  {32'hbe74286e, 32'h3e800618} /* (25, 8, 19) {real, imag} */,
  {32'hbed6d18a, 32'h3e24b51e} /* (25, 8, 18) {real, imag} */,
  {32'hbe195df7, 32'hbd9e6d7a} /* (25, 8, 17) {real, imag} */,
  {32'h3ea9fbac, 32'hbe8bc557} /* (25, 8, 16) {real, imag} */,
  {32'h3e7d077a, 32'h3ef7d72c} /* (25, 8, 15) {real, imag} */,
  {32'h3dd383a8, 32'hbf0d106b} /* (25, 8, 14) {real, imag} */,
  {32'h3d4591d8, 32'hbf1cc25b} /* (25, 8, 13) {real, imag} */,
  {32'hbecd2d90, 32'h3eb43660} /* (25, 8, 12) {real, imag} */,
  {32'h3ebd8652, 32'hbea9b408} /* (25, 8, 11) {real, imag} */,
  {32'h3e9aab6a, 32'h3de98a8a} /* (25, 8, 10) {real, imag} */,
  {32'h3e1e7b40, 32'h3d9a89b4} /* (25, 8, 9) {real, imag} */,
  {32'hbe2e9970, 32'hbf189e30} /* (25, 8, 8) {real, imag} */,
  {32'hbdad0482, 32'hbece6344} /* (25, 8, 7) {real, imag} */,
  {32'hbef54518, 32'hbe42cf94} /* (25, 8, 6) {real, imag} */,
  {32'hbd1c7080, 32'h3d75b8fc} /* (25, 8, 5) {real, imag} */,
  {32'hbe75d92a, 32'h3f6e730f} /* (25, 8, 4) {real, imag} */,
  {32'hbf5ff362, 32'h3e9297d6} /* (25, 8, 3) {real, imag} */,
  {32'hbf739902, 32'hbe883a64} /* (25, 8, 2) {real, imag} */,
  {32'h3fb3094d, 32'h3ecf4c7a} /* (25, 8, 1) {real, imag} */,
  {32'h3efdf5fa, 32'h3dfe68ee} /* (25, 8, 0) {real, imag} */,
  {32'hbf0ad48b, 32'hbeb54daa} /* (25, 7, 31) {real, imag} */,
  {32'h3e2f3e3c, 32'hbe7aa3a0} /* (25, 7, 30) {real, imag} */,
  {32'hbdfe4b14, 32'hbf3347a6} /* (25, 7, 29) {real, imag} */,
  {32'hbe9fbb24, 32'h3e48adcc} /* (25, 7, 28) {real, imag} */,
  {32'h3ce9e68c, 32'h3e34e45e} /* (25, 7, 27) {real, imag} */,
  {32'hbe984002, 32'hbea415e0} /* (25, 7, 26) {real, imag} */,
  {32'h3e582542, 32'hbeb27b17} /* (25, 7, 25) {real, imag} */,
  {32'h3db0ec86, 32'hbf849174} /* (25, 7, 24) {real, imag} */,
  {32'h3e587688, 32'h3ead5b1f} /* (25, 7, 23) {real, imag} */,
  {32'hbec378fe, 32'h3e023dcc} /* (25, 7, 22) {real, imag} */,
  {32'hbde62472, 32'hbef2fa71} /* (25, 7, 21) {real, imag} */,
  {32'hbc1a2168, 32'h3decdbb9} /* (25, 7, 20) {real, imag} */,
  {32'hbedda76d, 32'hbef15148} /* (25, 7, 19) {real, imag} */,
  {32'h3e343fe1, 32'hbe745803} /* (25, 7, 18) {real, imag} */,
  {32'h3dd2ab41, 32'h3ea081d8} /* (25, 7, 17) {real, imag} */,
  {32'hbdad7ade, 32'h3d627d44} /* (25, 7, 16) {real, imag} */,
  {32'hbe54377c, 32'h3e52e07a} /* (25, 7, 15) {real, imag} */,
  {32'hbca0a488, 32'hbdce5f6d} /* (25, 7, 14) {real, imag} */,
  {32'h3f04969e, 32'h3eac9750} /* (25, 7, 13) {real, imag} */,
  {32'hbe11ff30, 32'h3edac813} /* (25, 7, 12) {real, imag} */,
  {32'h3e5e08b8, 32'hbeb76f92} /* (25, 7, 11) {real, imag} */,
  {32'hbf32401c, 32'hbed68c1b} /* (25, 7, 10) {real, imag} */,
  {32'hbe1ce534, 32'hbeb50910} /* (25, 7, 9) {real, imag} */,
  {32'h3e1f565b, 32'h3e74d1f4} /* (25, 7, 8) {real, imag} */,
  {32'h3dd22f0c, 32'hbec0a940} /* (25, 7, 7) {real, imag} */,
  {32'hbec5a902, 32'hbc27a840} /* (25, 7, 6) {real, imag} */,
  {32'hbf0c5bf6, 32'h3ed28bfe} /* (25, 7, 5) {real, imag} */,
  {32'h3f22fe4c, 32'hbf3202f3} /* (25, 7, 4) {real, imag} */,
  {32'h3e7e936a, 32'h3f5584cc} /* (25, 7, 3) {real, imag} */,
  {32'h3d8180a4, 32'h3f514108} /* (25, 7, 2) {real, imag} */,
  {32'hbf5708f7, 32'hbf20f6b1} /* (25, 7, 1) {real, imag} */,
  {32'hbf83d5fe, 32'hbda9c4ca} /* (25, 7, 0) {real, imag} */,
  {32'h3ea161d2, 32'hbec95ee7} /* (25, 6, 31) {real, imag} */,
  {32'hbef89a47, 32'h3ee784f3} /* (25, 6, 30) {real, imag} */,
  {32'hbe7522e7, 32'h3dfe53f2} /* (25, 6, 29) {real, imag} */,
  {32'h3f4482ea, 32'hbf3cf13c} /* (25, 6, 28) {real, imag} */,
  {32'hbe2ad513, 32'hbec1be39} /* (25, 6, 27) {real, imag} */,
  {32'hbe2827f4, 32'h3f79ee26} /* (25, 6, 26) {real, imag} */,
  {32'hbe26f290, 32'h3e983f23} /* (25, 6, 25) {real, imag} */,
  {32'h3e14aca2, 32'hbe233576} /* (25, 6, 24) {real, imag} */,
  {32'h3e67204d, 32'h3f041b3f} /* (25, 6, 23) {real, imag} */,
  {32'h3e25008c, 32'h3eb060ff} /* (25, 6, 22) {real, imag} */,
  {32'h3e151cbb, 32'hbe212a8a} /* (25, 6, 21) {real, imag} */,
  {32'h3ea6afd0, 32'hbdb3dab0} /* (25, 6, 20) {real, imag} */,
  {32'hbe525501, 32'hbe24ee69} /* (25, 6, 19) {real, imag} */,
  {32'hbe617fd8, 32'h3c917988} /* (25, 6, 18) {real, imag} */,
  {32'h3e1b5be2, 32'hbd829d40} /* (25, 6, 17) {real, imag} */,
  {32'h3efb1526, 32'h3c79ddf0} /* (25, 6, 16) {real, imag} */,
  {32'hbc000178, 32'h3ece1e4e} /* (25, 6, 15) {real, imag} */,
  {32'hbe5180a6, 32'h3dee0796} /* (25, 6, 14) {real, imag} */,
  {32'h3ed8a848, 32'hbe7042f2} /* (25, 6, 13) {real, imag} */,
  {32'hbcc89ac8, 32'h3d20caa0} /* (25, 6, 12) {real, imag} */,
  {32'hbe528e72, 32'hbdbeab44} /* (25, 6, 11) {real, imag} */,
  {32'h3f0a54e5, 32'h3e4cf76c} /* (25, 6, 10) {real, imag} */,
  {32'h3e95293a, 32'h3d51856e} /* (25, 6, 9) {real, imag} */,
  {32'h3f08e4c9, 32'h3e8a2690} /* (25, 6, 8) {real, imag} */,
  {32'hbf16d020, 32'hbe5a20bc} /* (25, 6, 7) {real, imag} */,
  {32'h3edf8948, 32'hbeb474fc} /* (25, 6, 6) {real, imag} */,
  {32'h3e14659c, 32'hbcb9a474} /* (25, 6, 5) {real, imag} */,
  {32'h3e49778e, 32'hbf3c6d8d} /* (25, 6, 4) {real, imag} */,
  {32'h3e25fac4, 32'hbe080ab0} /* (25, 6, 3) {real, imag} */,
  {32'h3f432d6e, 32'hbe04b04c} /* (25, 6, 2) {real, imag} */,
  {32'hbe1640a1, 32'h3e398f75} /* (25, 6, 1) {real, imag} */,
  {32'h3d89d972, 32'h3cd20d00} /* (25, 6, 0) {real, imag} */,
  {32'h4028f802, 32'hbf04a4e4} /* (25, 5, 31) {real, imag} */,
  {32'hbf879cda, 32'hbf587950} /* (25, 5, 30) {real, imag} */,
  {32'h3eb91df4, 32'hbe63ff62} /* (25, 5, 29) {real, imag} */,
  {32'h3e141bb5, 32'h3efb89ec} /* (25, 5, 28) {real, imag} */,
  {32'hbfa3f762, 32'h3e6e848c} /* (25, 5, 27) {real, imag} */,
  {32'h3f3a2781, 32'hbecdc8c2} /* (25, 5, 26) {real, imag} */,
  {32'h3f1d87ad, 32'hbeec0be0} /* (25, 5, 25) {real, imag} */,
  {32'hbe208e68, 32'h3ec77fd0} /* (25, 5, 24) {real, imag} */,
  {32'hbe086c84, 32'hbe89edc8} /* (25, 5, 23) {real, imag} */,
  {32'h3e2c70bd, 32'h3e53b53e} /* (25, 5, 22) {real, imag} */,
  {32'hbef1087e, 32'hbcbe75d8} /* (25, 5, 21) {real, imag} */,
  {32'h3ee4da6b, 32'h3e175e26} /* (25, 5, 20) {real, imag} */,
  {32'h3eb5ffe8, 32'h3dc797a1} /* (25, 5, 19) {real, imag} */,
  {32'hbda05594, 32'h3ed6eca8} /* (25, 5, 18) {real, imag} */,
  {32'hbee69352, 32'hbd8d9da0} /* (25, 5, 17) {real, imag} */,
  {32'h3d4f91ec, 32'h3c8a0bb8} /* (25, 5, 16) {real, imag} */,
  {32'hbdd8e84e, 32'h3ec93f97} /* (25, 5, 15) {real, imag} */,
  {32'h3e28aa02, 32'h3e804d78} /* (25, 5, 14) {real, imag} */,
  {32'hbb969f78, 32'h3e5badc2} /* (25, 5, 13) {real, imag} */,
  {32'h3d1fd11a, 32'h3e7f99e8} /* (25, 5, 12) {real, imag} */,
  {32'hbdcce098, 32'hbf3890b6} /* (25, 5, 11) {real, imag} */,
  {32'h3d5e39b0, 32'hbeed6cd6} /* (25, 5, 10) {real, imag} */,
  {32'hbf0dab18, 32'hbebfb2b6} /* (25, 5, 9) {real, imag} */,
  {32'hbda8b09c, 32'hbd838a04} /* (25, 5, 8) {real, imag} */,
  {32'h3e97b582, 32'h3e827211} /* (25, 5, 7) {real, imag} */,
  {32'hbdc0d3c8, 32'h3e1cdadc} /* (25, 5, 6) {real, imag} */,
  {32'h3f65cf84, 32'hbe976e91} /* (25, 5, 5) {real, imag} */,
  {32'hbeb81486, 32'h3ed95528} /* (25, 5, 4) {real, imag} */,
  {32'h3cf11870, 32'hbf82c8a4} /* (25, 5, 3) {real, imag} */,
  {32'hbf8556c6, 32'hbfa8ec60} /* (25, 5, 2) {real, imag} */,
  {32'h3fb88489, 32'h401edf1e} /* (25, 5, 1) {real, imag} */,
  {32'h3f89b2dc, 32'h3fcb057a} /* (25, 5, 0) {real, imag} */,
  {32'hbf8b4cb0, 32'hc00ba980} /* (25, 4, 31) {real, imag} */,
  {32'h3fabde28, 32'h4012508d} /* (25, 4, 30) {real, imag} */,
  {32'hbf1e76c3, 32'hbe755a6e} /* (25, 4, 29) {real, imag} */,
  {32'hbf89d772, 32'hbf9a93f5} /* (25, 4, 28) {real, imag} */,
  {32'h3e4167df, 32'hbc4b2e10} /* (25, 4, 27) {real, imag} */,
  {32'hbdf8bcd8, 32'hbf579b3c} /* (25, 4, 26) {real, imag} */,
  {32'h3e8a4d82, 32'h3e9e4403} /* (25, 4, 25) {real, imag} */,
  {32'h3c90c830, 32'h3de8e8d0} /* (25, 4, 24) {real, imag} */,
  {32'hbe10bfea, 32'hbe66ab51} /* (25, 4, 23) {real, imag} */,
  {32'hbeba97a6, 32'hbe2cdbc0} /* (25, 4, 22) {real, imag} */,
  {32'h3e62c443, 32'h3f053101} /* (25, 4, 21) {real, imag} */,
  {32'h3d696b78, 32'hbc433560} /* (25, 4, 20) {real, imag} */,
  {32'hbe653144, 32'h3e867ab2} /* (25, 4, 19) {real, imag} */,
  {32'h3f0e9bee, 32'hbe13e7d0} /* (25, 4, 18) {real, imag} */,
  {32'h3d45be7c, 32'h3e68a313} /* (25, 4, 17) {real, imag} */,
  {32'hbc7c99fe, 32'h3e3ab18a} /* (25, 4, 16) {real, imag} */,
  {32'hbe341313, 32'hbd2bce2c} /* (25, 4, 15) {real, imag} */,
  {32'h3d73a3e0, 32'hbdff2100} /* (25, 4, 14) {real, imag} */,
  {32'h3e8253f6, 32'h3e61c37c} /* (25, 4, 13) {real, imag} */,
  {32'h3da51f20, 32'hbcdf4f30} /* (25, 4, 12) {real, imag} */,
  {32'h3eaafa78, 32'h3f2e7fa2} /* (25, 4, 11) {real, imag} */,
  {32'h3d980685, 32'hbe1312d3} /* (25, 4, 10) {real, imag} */,
  {32'hbe74b68c, 32'h3ebc036e} /* (25, 4, 9) {real, imag} */,
  {32'h3efb6267, 32'h3f7982f6} /* (25, 4, 8) {real, imag} */,
  {32'hbf37d815, 32'h3e9fd46d} /* (25, 4, 7) {real, imag} */,
  {32'hbf4d1b52, 32'h3f536dd4} /* (25, 4, 6) {real, imag} */,
  {32'h3e96da0c, 32'h3b918b80} /* (25, 4, 5) {real, imag} */,
  {32'h3e91834b, 32'hbffeae9b} /* (25, 4, 4) {real, imag} */,
  {32'hbe24025c, 32'hbdfdc67a} /* (25, 4, 3) {real, imag} */,
  {32'h3fe4ec3e, 32'h3fc350b5} /* (25, 4, 2) {real, imag} */,
  {32'hc06053b4, 32'hbf01c330} /* (25, 4, 1) {real, imag} */,
  {32'hbfca60d6, 32'hbf974fad} /* (25, 4, 0) {real, imag} */,
  {32'h400d6642, 32'hc01f3f28} /* (25, 3, 31) {real, imag} */,
  {32'hbea3e0a8, 32'h3febde3d} /* (25, 3, 30) {real, imag} */,
  {32'h3f2ddf9e, 32'h3ed80e26} /* (25, 3, 29) {real, imag} */,
  {32'hbf4e4370, 32'hbf208bd4} /* (25, 3, 28) {real, imag} */,
  {32'h3eeabea8, 32'hbd9821e8} /* (25, 3, 27) {real, imag} */,
  {32'hbcab5230, 32'h3e54ba12} /* (25, 3, 26) {real, imag} */,
  {32'h3e49f958, 32'h3e89e0fa} /* (25, 3, 25) {real, imag} */,
  {32'h3ede588d, 32'h3f5b916c} /* (25, 3, 24) {real, imag} */,
  {32'h3df369b4, 32'hbee92c34} /* (25, 3, 23) {real, imag} */,
  {32'hbe0e16be, 32'h3e69ba4a} /* (25, 3, 22) {real, imag} */,
  {32'hbd0d6c22, 32'h3e4910e0} /* (25, 3, 21) {real, imag} */,
  {32'hbdbf1ab9, 32'h3eaed7a0} /* (25, 3, 20) {real, imag} */,
  {32'h3ec8745a, 32'hbe2fd396} /* (25, 3, 19) {real, imag} */,
  {32'h3e991012, 32'h3e39eeae} /* (25, 3, 18) {real, imag} */,
  {32'h3b8c44b8, 32'hbe346f5d} /* (25, 3, 17) {real, imag} */,
  {32'hbe59fbd5, 32'h3e4ecdf1} /* (25, 3, 16) {real, imag} */,
  {32'h3de1958c, 32'h3da6a4b7} /* (25, 3, 15) {real, imag} */,
  {32'hbee609ca, 32'hbdd111b2} /* (25, 3, 14) {real, imag} */,
  {32'h3dbf0a54, 32'h3e83a276} /* (25, 3, 13) {real, imag} */,
  {32'h3ec8094d, 32'hbe25df7a} /* (25, 3, 12) {real, imag} */,
  {32'hbf0a8f00, 32'hbdd29ac4} /* (25, 3, 11) {real, imag} */,
  {32'hbd6a2caa, 32'h3dbe7304} /* (25, 3, 10) {real, imag} */,
  {32'hbd883f66, 32'hbe6a6a4a} /* (25, 3, 9) {real, imag} */,
  {32'hbebb0c1e, 32'hbe84cd56} /* (25, 3, 8) {real, imag} */,
  {32'hbe42ff4c, 32'h3d0d42be} /* (25, 3, 7) {real, imag} */,
  {32'hbdb549d8, 32'h3f0e9266} /* (25, 3, 6) {real, imag} */,
  {32'hbf52fc5e, 32'hbef5dcd8} /* (25, 3, 5) {real, imag} */,
  {32'h3f45d2e2, 32'hbe2516c8} /* (25, 3, 4) {real, imag} */,
  {32'hbd8c1486, 32'hbf0dcfcd} /* (25, 3, 3) {real, imag} */,
  {32'h3e43a557, 32'h403cd155} /* (25, 3, 2) {real, imag} */,
  {32'hc03703a1, 32'hbfbc75bf} /* (25, 3, 1) {real, imag} */,
  {32'h401cc1ef, 32'h3f1c36dc} /* (25, 3, 0) {real, imag} */,
  {32'h41924ac2, 32'h40174649} /* (25, 2, 31) {real, imag} */,
  {32'hc10b0d3a, 32'h3fcb1585} /* (25, 2, 30) {real, imag} */,
  {32'h3f4b205e, 32'hbf652d8e} /* (25, 2, 29) {real, imag} */,
  {32'h3f80646f, 32'hbf9d9bb9} /* (25, 2, 28) {real, imag} */,
  {32'h3d18c7f0, 32'hbed2c160} /* (25, 2, 27) {real, imag} */,
  {32'h3e48d3e0, 32'h3cc123f0} /* (25, 2, 26) {real, imag} */,
  {32'hb92f1800, 32'h3f792af4} /* (25, 2, 25) {real, imag} */,
  {32'hbecca1ad, 32'h3f822582} /* (25, 2, 24) {real, imag} */,
  {32'h3e8fe85f, 32'h3ca23f38} /* (25, 2, 23) {real, imag} */,
  {32'h3e707241, 32'hbf487158} /* (25, 2, 22) {real, imag} */,
  {32'hbdb7db4a, 32'hbe96d028} /* (25, 2, 21) {real, imag} */,
  {32'hbc0bf2b0, 32'hbe739ca0} /* (25, 2, 20) {real, imag} */,
  {32'h3ca437cc, 32'h3d7024f4} /* (25, 2, 19) {real, imag} */,
  {32'hbe23d4f4, 32'h3e7016c0} /* (25, 2, 18) {real, imag} */,
  {32'hbe548374, 32'hbecddffa} /* (25, 2, 17) {real, imag} */,
  {32'hbe6a1156, 32'h3e4d9fe1} /* (25, 2, 16) {real, imag} */,
  {32'h3e60c574, 32'h3e1a5ed1} /* (25, 2, 15) {real, imag} */,
  {32'hbd67cd48, 32'h3ed03225} /* (25, 2, 14) {real, imag} */,
  {32'h3e89a426, 32'h3d17197c} /* (25, 2, 13) {real, imag} */,
  {32'hbd33a4a8, 32'hbf15536b} /* (25, 2, 12) {real, imag} */,
  {32'hbe5a26df, 32'hbf6ec50f} /* (25, 2, 11) {real, imag} */,
  {32'h3edf2f14, 32'h3e860087} /* (25, 2, 10) {real, imag} */,
  {32'hbd2b8274, 32'hbeecc5f6} /* (25, 2, 9) {real, imag} */,
  {32'hbf07854d, 32'hbe587b6e} /* (25, 2, 8) {real, imag} */,
  {32'h3f6a4924, 32'h3ee9d390} /* (25, 2, 7) {real, imag} */,
  {32'hbe22a9fe, 32'hbec3250d} /* (25, 2, 6) {real, imag} */,
  {32'hc00778e3, 32'hbf8769b3} /* (25, 2, 5) {real, imag} */,
  {32'h3fc30485, 32'hbdce70f4} /* (25, 2, 4) {real, imag} */,
  {32'hbf1386fb, 32'hbe7806b4} /* (25, 2, 3) {real, imag} */,
  {32'hc0ab65b9, 32'h3f935d2d} /* (25, 2, 2) {real, imag} */,
  {32'h4131396f, 32'h3f0b3d40} /* (25, 2, 1) {real, imag} */,
  {32'h412f9197, 32'h3f21350c} /* (25, 2, 0) {real, imag} */,
  {32'hc1c64ef4, 32'h40b23f18} /* (25, 1, 31) {real, imag} */,
  {32'h40bc3442, 32'h405fe528} /* (25, 1, 30) {real, imag} */,
  {32'h3f5217c5, 32'hbf2fe7c8} /* (25, 1, 29) {real, imag} */,
  {32'hbfa3353e, 32'hbf48d99e} /* (25, 1, 28) {real, imag} */,
  {32'h40078014, 32'hbece00d6} /* (25, 1, 27) {real, imag} */,
  {32'hbf3494fb, 32'hbe2bd18c} /* (25, 1, 26) {real, imag} */,
  {32'hbf00ef26, 32'h3ea83732} /* (25, 1, 25) {real, imag} */,
  {32'h3d6e04f0, 32'hbd3b3408} /* (25, 1, 24) {real, imag} */,
  {32'h3d8856a9, 32'h3ef2155e} /* (25, 1, 23) {real, imag} */,
  {32'hbd68b750, 32'hbf07fb38} /* (25, 1, 22) {real, imag} */,
  {32'h3f412222, 32'hbef21ba8} /* (25, 1, 21) {real, imag} */,
  {32'h3ecf9a2e, 32'hbdf55af7} /* (25, 1, 20) {real, imag} */,
  {32'hbe3bd3fd, 32'hbce73428} /* (25, 1, 19) {real, imag} */,
  {32'h3e4e2313, 32'hbf07981c} /* (25, 1, 18) {real, imag} */,
  {32'hbddd30c6, 32'h3e1e5d68} /* (25, 1, 17) {real, imag} */,
  {32'h3d9de935, 32'h3eacee39} /* (25, 1, 16) {real, imag} */,
  {32'hbea3ad74, 32'hbeeb3d5f} /* (25, 1, 15) {real, imag} */,
  {32'hbebaaa8d, 32'h3ef0d1e0} /* (25, 1, 14) {real, imag} */,
  {32'h3e569b90, 32'hbe6a93da} /* (25, 1, 13) {real, imag} */,
  {32'hbd374e4e, 32'h3d64efcc} /* (25, 1, 12) {real, imag} */,
  {32'h3ec42a38, 32'h3f483c00} /* (25, 1, 11) {real, imag} */,
  {32'h3e389066, 32'h3d2bb4a8} /* (25, 1, 10) {real, imag} */,
  {32'h3e8b0e3d, 32'hbe8b89ba} /* (25, 1, 9) {real, imag} */,
  {32'h3e83e51f, 32'h3f7b5807} /* (25, 1, 8) {real, imag} */,
  {32'hbe01714b, 32'h3db48370} /* (25, 1, 7) {real, imag} */,
  {32'h3eef6cb3, 32'h3efe8b53} /* (25, 1, 6) {real, imag} */,
  {32'h3fc05e16, 32'h3fb57b70} /* (25, 1, 5) {real, imag} */,
  {32'hbd8a35c0, 32'hbff53126} /* (25, 1, 4) {real, imag} */,
  {32'h3f9710a7, 32'hbd25f380} /* (25, 1, 3) {real, imag} */,
  {32'h410543ce, 32'h410875b1} /* (25, 1, 2) {real, imag} */,
  {32'hc2124069, 32'hc1aea98b} /* (25, 1, 1) {real, imag} */,
  {32'hc213f352, 32'hc0bfcf31} /* (25, 1, 0) {real, imag} */,
  {32'hc1e3a334, 32'h41ad9fb2} /* (25, 0, 31) {real, imag} */,
  {32'h3ff4f99d, 32'hbfb3c9a4} /* (25, 0, 30) {real, imag} */,
  {32'h3f51fbc1, 32'hbf5782d7} /* (25, 0, 29) {real, imag} */,
  {32'h3f442766, 32'hc0101663} /* (25, 0, 28) {real, imag} */,
  {32'h40085bc8, 32'hbea13bfc} /* (25, 0, 27) {real, imag} */,
  {32'hbe14cec5, 32'h3ef17d91} /* (25, 0, 26) {real, imag} */,
  {32'hbc90e378, 32'h3b611400} /* (25, 0, 25) {real, imag} */,
  {32'hbf26ce92, 32'hbfde0c8a} /* (25, 0, 24) {real, imag} */,
  {32'h3eb84fc4, 32'hbf2e4e71} /* (25, 0, 23) {real, imag} */,
  {32'h3d63dd04, 32'hbc106d68} /* (25, 0, 22) {real, imag} */,
  {32'h3edfcbac, 32'hbe665d57} /* (25, 0, 21) {real, imag} */,
  {32'hbed7e5f8, 32'hbec1688c} /* (25, 0, 20) {real, imag} */,
  {32'h3e80d74c, 32'h3e212a80} /* (25, 0, 19) {real, imag} */,
  {32'hbe386dc6, 32'hbf34cefd} /* (25, 0, 18) {real, imag} */,
  {32'h3e29387c, 32'h3cbff458} /* (25, 0, 17) {real, imag} */,
  {32'h3f1c8272, 32'h00000000} /* (25, 0, 16) {real, imag} */,
  {32'h3e29387c, 32'hbcbff458} /* (25, 0, 15) {real, imag} */,
  {32'hbe386dc6, 32'h3f34cefd} /* (25, 0, 14) {real, imag} */,
  {32'h3e80d74c, 32'hbe212a80} /* (25, 0, 13) {real, imag} */,
  {32'hbed7e5f8, 32'h3ec1688c} /* (25, 0, 12) {real, imag} */,
  {32'h3edfcbac, 32'h3e665d57} /* (25, 0, 11) {real, imag} */,
  {32'h3d63dd04, 32'h3c106d68} /* (25, 0, 10) {real, imag} */,
  {32'h3eb84fc4, 32'h3f2e4e71} /* (25, 0, 9) {real, imag} */,
  {32'hbf26ce92, 32'h3fde0c8a} /* (25, 0, 8) {real, imag} */,
  {32'hbc90e378, 32'hbb611400} /* (25, 0, 7) {real, imag} */,
  {32'hbe14cec5, 32'hbef17d91} /* (25, 0, 6) {real, imag} */,
  {32'h40085bc8, 32'h3ea13bfc} /* (25, 0, 5) {real, imag} */,
  {32'h3f442766, 32'h40101663} /* (25, 0, 4) {real, imag} */,
  {32'h3f51fbc1, 32'h3f5782d7} /* (25, 0, 3) {real, imag} */,
  {32'h3ff4f99d, 32'h3fb3c9a4} /* (25, 0, 2) {real, imag} */,
  {32'hc1e3a334, 32'hc1ad9fb2} /* (25, 0, 1) {real, imag} */,
  {32'hc23bf222, 32'h00000000} /* (25, 0, 0) {real, imag} */,
  {32'hc25a1b49, 32'h41fba9e1} /* (24, 31, 31) {real, imag} */,
  {32'h4153f596, 32'hc14c952c} /* (24, 31, 30) {real, imag} */,
  {32'h3f2cdc58, 32'hbef6266a} /* (24, 31, 29) {real, imag} */,
  {32'hbf48c5bc, 32'h3fc0efb0} /* (24, 31, 28) {real, imag} */,
  {32'h4006aabc, 32'hbfbd260a} /* (24, 31, 27) {real, imag} */,
  {32'h3efa6cdc, 32'h3d201aa8} /* (24, 31, 26) {real, imag} */,
  {32'hbec65812, 32'h3eeb890a} /* (24, 31, 25) {real, imag} */,
  {32'h3f497c17, 32'hbf59d703} /* (24, 31, 24) {real, imag} */,
  {32'hbaf3f480, 32'hbe7dbbe6} /* (24, 31, 23) {real, imag} */,
  {32'hbe57a006, 32'h3e76db3a} /* (24, 31, 22) {real, imag} */,
  {32'h3e4c3c0d, 32'hbf011cc6} /* (24, 31, 21) {real, imag} */,
  {32'hbddc2fc6, 32'h3cb40ca0} /* (24, 31, 20) {real, imag} */,
  {32'hbb3b4ba0, 32'h3ecefacc} /* (24, 31, 19) {real, imag} */,
  {32'hbe69c1a8, 32'hbefd4c14} /* (24, 31, 18) {real, imag} */,
  {32'hbc3d1c00, 32'h3ddc9e08} /* (24, 31, 17) {real, imag} */,
  {32'h3cc46fc8, 32'h3dc209b4} /* (24, 31, 16) {real, imag} */,
  {32'h3d9bd268, 32'hbe5fb4ea} /* (24, 31, 15) {real, imag} */,
  {32'hbd587bf8, 32'h3f0aa1f2} /* (24, 31, 14) {real, imag} */,
  {32'h3e17426a, 32'h3f11c677} /* (24, 31, 13) {real, imag} */,
  {32'hbf23941a, 32'hbe8842c2} /* (24, 31, 12) {real, imag} */,
  {32'h3e9b3418, 32'h3f4e1184} /* (24, 31, 11) {real, imag} */,
  {32'h3e2d67a2, 32'h3f221b46} /* (24, 31, 10) {real, imag} */,
  {32'h3edfb864, 32'hbe1fab2d} /* (24, 31, 9) {real, imag} */,
  {32'h3f6df247, 32'h3f756b36} /* (24, 31, 8) {real, imag} */,
  {32'hbf2995b9, 32'hbf171191} /* (24, 31, 7) {real, imag} */,
  {32'hbf64ff74, 32'h3e5e3bb6} /* (24, 31, 6) {real, imag} */,
  {32'h403d1066, 32'h3e9dc783} /* (24, 31, 5) {real, imag} */,
  {32'hc031d835, 32'h3f0f146e} /* (24, 31, 4) {real, imag} */,
  {32'h3fbcef3e, 32'h3f5067d0} /* (24, 31, 3) {real, imag} */,
  {32'h410a21ab, 32'hc0355130} /* (24, 31, 2) {real, imag} */,
  {32'hc2177b8b, 32'hc117591a} /* (24, 31, 1) {real, imag} */,
  {32'hc24ea4af, 32'h40dbd352} /* (24, 31, 0) {real, imag} */,
  {32'h4183bf18, 32'h3f8b6cb7} /* (24, 30, 31) {real, imag} */,
  {32'hc104b84e, 32'hbfa1f5cc} /* (24, 30, 30) {real, imag} */,
  {32'h3e8689ce, 32'h3fa4e195} /* (24, 30, 29) {real, imag} */,
  {32'h40349c5c, 32'hbf28ef62} /* (24, 30, 28) {real, imag} */,
  {32'hc01e93f2, 32'h3f9c20fb} /* (24, 30, 27) {real, imag} */,
  {32'h3f485b5a, 32'hbb0a57c0} /* (24, 30, 26) {real, imag} */,
  {32'h3ef633d0, 32'hbe60b594} /* (24, 30, 25) {real, imag} */,
  {32'hbf0d9b6e, 32'hbe51e0cf} /* (24, 30, 24) {real, imag} */,
  {32'h3e79165d, 32'hbc51be70} /* (24, 30, 23) {real, imag} */,
  {32'h3ea1e90f, 32'h3f0abe24} /* (24, 30, 22) {real, imag} */,
  {32'hbe86951e, 32'h3f0a8943} /* (24, 30, 21) {real, imag} */,
  {32'h3e9e9f07, 32'hbebeb63c} /* (24, 30, 20) {real, imag} */,
  {32'hbe129db8, 32'h3eecd54e} /* (24, 30, 19) {real, imag} */,
  {32'hbd376e04, 32'h3e1ec6f6} /* (24, 30, 18) {real, imag} */,
  {32'h3dc35ade, 32'h3e450d37} /* (24, 30, 17) {real, imag} */,
  {32'hbe32c55c, 32'hbdfb3631} /* (24, 30, 16) {real, imag} */,
  {32'hbe3c473e, 32'hbcbf3598} /* (24, 30, 15) {real, imag} */,
  {32'h3d681c4a, 32'hbe61a8ff} /* (24, 30, 14) {real, imag} */,
  {32'hbe367834, 32'hbea4fbdf} /* (24, 30, 13) {real, imag} */,
  {32'hbd8870b4, 32'h3ef43f38} /* (24, 30, 12) {real, imag} */,
  {32'h3f6617f8, 32'hbed8d9fe} /* (24, 30, 11) {real, imag} */,
  {32'hbe9f356f, 32'h3ee11de0} /* (24, 30, 10) {real, imag} */,
  {32'h3f0916ba, 32'hbdb6bbbe} /* (24, 30, 9) {real, imag} */,
  {32'h3c4d80c0, 32'hbf9581f2} /* (24, 30, 8) {real, imag} */,
  {32'hbeaa64c7, 32'hbea798e2} /* (24, 30, 7) {real, imag} */,
  {32'hbf41d6bc, 32'hbea976a5} /* (24, 30, 6) {real, imag} */,
  {32'hbf7e4eb0, 32'hbea7d3d1} /* (24, 30, 5) {real, imag} */,
  {32'h3fcc8c7c, 32'h3fc4b9aa} /* (24, 30, 4) {real, imag} */,
  {32'h3fb71b66, 32'h3f604c0a} /* (24, 30, 3) {real, imag} */,
  {32'hc15475c7, 32'hc0491990} /* (24, 30, 2) {real, imag} */,
  {32'h41e1eb34, 32'hbfe216af} /* (24, 30, 1) {real, imag} */,
  {32'h4170ba5e, 32'hc0121bb6} /* (24, 30, 0) {real, imag} */,
  {32'hc06a3ab7, 32'h402e5ab6} /* (24, 29, 31) {real, imag} */,
  {32'hbf3d8f3c, 32'hc07b3b78} /* (24, 29, 30) {real, imag} */,
  {32'h3be41d40, 32'h3df2ac48} /* (24, 29, 29) {real, imag} */,
  {32'h3fb53f41, 32'h3f1c749e} /* (24, 29, 28) {real, imag} */,
  {32'hbe74c42d, 32'h3f174d74} /* (24, 29, 27) {real, imag} */,
  {32'hbef947b9, 32'hbf7b27a8} /* (24, 29, 26) {real, imag} */,
  {32'hbec0b7c2, 32'h3cea4a60} /* (24, 29, 25) {real, imag} */,
  {32'h3dce781c, 32'hbdff605e} /* (24, 29, 24) {real, imag} */,
  {32'h3ea37a9c, 32'h3db111da} /* (24, 29, 23) {real, imag} */,
  {32'h3e3fb824, 32'h3c1e5a58} /* (24, 29, 22) {real, imag} */,
  {32'h3e7486fe, 32'hbcb0a94c} /* (24, 29, 21) {real, imag} */,
  {32'hbd6feac8, 32'h3d297c70} /* (24, 29, 20) {real, imag} */,
  {32'hbf47c258, 32'h3df57863} /* (24, 29, 19) {real, imag} */,
  {32'hbc0f6978, 32'hbd91da00} /* (24, 29, 18) {real, imag} */,
  {32'h3d21a4e8, 32'h3d4732c0} /* (24, 29, 17) {real, imag} */,
  {32'h3e4e5534, 32'h3dd980f4} /* (24, 29, 16) {real, imag} */,
  {32'hbdbd6eac, 32'hbd9c51d3} /* (24, 29, 15) {real, imag} */,
  {32'h3e99eda7, 32'hbf370f59} /* (24, 29, 14) {real, imag} */,
  {32'hbd8d48ac, 32'h3f181ee6} /* (24, 29, 13) {real, imag} */,
  {32'h3d688362, 32'hbe4514c1} /* (24, 29, 12) {real, imag} */,
  {32'hbe0808b6, 32'h3f0ab045} /* (24, 29, 11) {real, imag} */,
  {32'h3e507c55, 32'hbe8b42fe} /* (24, 29, 10) {real, imag} */,
  {32'hbf1c1dc0, 32'hbe197d6d} /* (24, 29, 9) {real, imag} */,
  {32'hbe9ddd94, 32'hbf2bcb94} /* (24, 29, 8) {real, imag} */,
  {32'hbe30bddc, 32'h3ede12ca} /* (24, 29, 7) {real, imag} */,
  {32'hbe324cc2, 32'hbea762ec} /* (24, 29, 6) {real, imag} */,
  {32'h3f99523e, 32'hbe89de0d} /* (24, 29, 5) {real, imag} */,
  {32'hbf30c5a2, 32'h3f7cc259} /* (24, 29, 4) {real, imag} */,
  {32'h3eae0e67, 32'hbf6e17d9} /* (24, 29, 3) {real, imag} */,
  {32'hc00909d8, 32'hc02a7b68} /* (24, 29, 2) {real, imag} */,
  {32'h406e42f4, 32'h403b5b5c} /* (24, 29, 1) {real, imag} */,
  {32'h403aac1c, 32'hbeb32833} /* (24, 29, 0) {real, imag} */,
  {32'hc08f7771, 32'h3f8d80e7} /* (24, 28, 31) {real, imag} */,
  {32'h40769f0c, 32'hbfce413e} /* (24, 28, 30) {real, imag} */,
  {32'h3f2cbf7c, 32'h3ec4c790} /* (24, 28, 29) {real, imag} */,
  {32'h3f59b7e6, 32'h3fdd0dee} /* (24, 28, 28) {real, imag} */,
  {32'hbe9622e1, 32'hbf2dfb16} /* (24, 28, 27) {real, imag} */,
  {32'hbf512acd, 32'hbddb0574} /* (24, 28, 26) {real, imag} */,
  {32'hbf291dd4, 32'hbe5561fc} /* (24, 28, 25) {real, imag} */,
  {32'hbe1c8886, 32'hbed58dee} /* (24, 28, 24) {real, imag} */,
  {32'h3ef24d46, 32'hbe3ee805} /* (24, 28, 23) {real, imag} */,
  {32'h3eb8bd7f, 32'h3f008031} /* (24, 28, 22) {real, imag} */,
  {32'hbda9feda, 32'hbf0213d6} /* (24, 28, 21) {real, imag} */,
  {32'hbe9711e0, 32'h3e96043e} /* (24, 28, 20) {real, imag} */,
  {32'h3e46e964, 32'h3ea15006} /* (24, 28, 19) {real, imag} */,
  {32'h3e0160ae, 32'hbe926220} /* (24, 28, 18) {real, imag} */,
  {32'hbb4d8680, 32'h3e76ca73} /* (24, 28, 17) {real, imag} */,
  {32'hbe5567d2, 32'hbdbc08e7} /* (24, 28, 16) {real, imag} */,
  {32'h3e6572e8, 32'hbee99fd0} /* (24, 28, 15) {real, imag} */,
  {32'h3e272405, 32'h3e3c16ea} /* (24, 28, 14) {real, imag} */,
  {32'hbe260275, 32'h3e7022ee} /* (24, 28, 13) {real, imag} */,
  {32'hbd67ece0, 32'h3d6e9530} /* (24, 28, 12) {real, imag} */,
  {32'h3eaf6748, 32'hbe377b8e} /* (24, 28, 11) {real, imag} */,
  {32'hbf085499, 32'hbe5b455c} /* (24, 28, 10) {real, imag} */,
  {32'h3f2c2990, 32'h3ee13998} /* (24, 28, 9) {real, imag} */,
  {32'h3f0adde4, 32'hbec2ceab} /* (24, 28, 8) {real, imag} */,
  {32'hbd718830, 32'hbdba8748} /* (24, 28, 7) {real, imag} */,
  {32'h3f2dbcfe, 32'h3f1a5c43} /* (24, 28, 6) {real, imag} */,
  {32'h3ec795a8, 32'h3eef6cb8} /* (24, 28, 5) {real, imag} */,
  {32'hbfe3deca, 32'h3f923c7d} /* (24, 28, 4) {real, imag} */,
  {32'h3d181108, 32'h3f6a39f2} /* (24, 28, 3) {real, imag} */,
  {32'h4012366f, 32'hc0499c03} /* (24, 28, 2) {real, imag} */,
  {32'hbfaf51f3, 32'h403b7c9e} /* (24, 28, 1) {real, imag} */,
  {32'hc0170c33, 32'h3f7776a4} /* (24, 28, 0) {real, imag} */,
  {32'h3fd43057, 32'hc027e872} /* (24, 27, 31) {real, imag} */,
  {32'hbf85c5e0, 32'h3fb14f54} /* (24, 27, 30) {real, imag} */,
  {32'h3ee4cd44, 32'h3e9e4582} /* (24, 27, 29) {real, imag} */,
  {32'h3dd0ba0c, 32'hbf8157cc} /* (24, 27, 28) {real, imag} */,
  {32'h3d67c470, 32'h3f0a69a6} /* (24, 27, 27) {real, imag} */,
  {32'hbebfe688, 32'h3bd9b380} /* (24, 27, 26) {real, imag} */,
  {32'h3ec1b58c, 32'hbe756444} /* (24, 27, 25) {real, imag} */,
  {32'h3da801d8, 32'h3f049e9a} /* (24, 27, 24) {real, imag} */,
  {32'hbf0812e2, 32'hbe41b86e} /* (24, 27, 23) {real, imag} */,
  {32'h3e8477ec, 32'h3e4158ee} /* (24, 27, 22) {real, imag} */,
  {32'h3dbc3e9b, 32'hbde423d4} /* (24, 27, 21) {real, imag} */,
  {32'h3e5be933, 32'h3d42e406} /* (24, 27, 20) {real, imag} */,
  {32'hbefb5636, 32'h3eb8926b} /* (24, 27, 19) {real, imag} */,
  {32'hbe3c3010, 32'h3ed183d1} /* (24, 27, 18) {real, imag} */,
  {32'hbe93444c, 32'h3df26188} /* (24, 27, 17) {real, imag} */,
  {32'h3e5ccb34, 32'hbdd0c612} /* (24, 27, 16) {real, imag} */,
  {32'hbe2de89a, 32'hbc9ff5e6} /* (24, 27, 15) {real, imag} */,
  {32'hbe425a2a, 32'hbe029510} /* (24, 27, 14) {real, imag} */,
  {32'h3e81c6c8, 32'h3e9be939} /* (24, 27, 13) {real, imag} */,
  {32'hbdc875de, 32'hbd629874} /* (24, 27, 12) {real, imag} */,
  {32'hbe5a5e72, 32'h3c8fa0a0} /* (24, 27, 11) {real, imag} */,
  {32'hbe80da3d, 32'hbea23213} /* (24, 27, 10) {real, imag} */,
  {32'h3d7d82fa, 32'hbcf80d18} /* (24, 27, 9) {real, imag} */,
  {32'hbe403cbc, 32'h3e94f407} /* (24, 27, 8) {real, imag} */,
  {32'hbec06f0a, 32'h3ebcb7fe} /* (24, 27, 7) {real, imag} */,
  {32'h3f248003, 32'hbd45ef68} /* (24, 27, 6) {real, imag} */,
  {32'hbf7cc1ae, 32'hbf35833a} /* (24, 27, 5) {real, imag} */,
  {32'h3e37cb82, 32'hbdbeeb96} /* (24, 27, 4) {real, imag} */,
  {32'h3e7c0ebd, 32'h3f0639f2} /* (24, 27, 3) {real, imag} */,
  {32'hbfe2499d, 32'hbce20c40} /* (24, 27, 2) {real, imag} */,
  {32'h406763bc, 32'hbef0a48d} /* (24, 27, 1) {real, imag} */,
  {32'h3fc1438a, 32'hbf76d6c1} /* (24, 27, 0) {real, imag} */,
  {32'hbe911978, 32'h3e09fe5b} /* (24, 26, 31) {real, imag} */,
  {32'h3f90c538, 32'h3ddc70aa} /* (24, 26, 30) {real, imag} */,
  {32'h3d15d6bc, 32'hbde17376} /* (24, 26, 29) {real, imag} */,
  {32'h3ecc1193, 32'hbeb7ad74} /* (24, 26, 28) {real, imag} */,
  {32'h3f370c02, 32'hbd6556f8} /* (24, 26, 27) {real, imag} */,
  {32'h3afd6880, 32'h3f533a36} /* (24, 26, 26) {real, imag} */,
  {32'hbeb7e425, 32'hbe613e98} /* (24, 26, 25) {real, imag} */,
  {32'hbe86aba6, 32'h3e953478} /* (24, 26, 24) {real, imag} */,
  {32'h3f3fcafa, 32'h3ea2c0ca} /* (24, 26, 23) {real, imag} */,
  {32'hbec9e764, 32'hbe8ac272} /* (24, 26, 22) {real, imag} */,
  {32'hbf346da8, 32'hbc06fa20} /* (24, 26, 21) {real, imag} */,
  {32'hbdf60737, 32'h3f14597c} /* (24, 26, 20) {real, imag} */,
  {32'hbe8f0e0a, 32'h3d89e157} /* (24, 26, 19) {real, imag} */,
  {32'h3e988a54, 32'hbe44a596} /* (24, 26, 18) {real, imag} */,
  {32'h3e05609e, 32'h3df81e8c} /* (24, 26, 17) {real, imag} */,
  {32'hbbe9df00, 32'h3d471596} /* (24, 26, 16) {real, imag} */,
  {32'h3b5aefb0, 32'hbea713a1} /* (24, 26, 15) {real, imag} */,
  {32'h3d4f319c, 32'h3e8f6c61} /* (24, 26, 14) {real, imag} */,
  {32'h3f310193, 32'h3e764879} /* (24, 26, 13) {real, imag} */,
  {32'h3ee9c9fc, 32'h3d0576c0} /* (24, 26, 12) {real, imag} */,
  {32'hbec15463, 32'hbe5d6df0} /* (24, 26, 11) {real, imag} */,
  {32'hbea0375e, 32'h3e4233b3} /* (24, 26, 10) {real, imag} */,
  {32'hbed46a88, 32'hbc0d88c0} /* (24, 26, 9) {real, imag} */,
  {32'hbcb72104, 32'h3f394bda} /* (24, 26, 8) {real, imag} */,
  {32'hbdaaef31, 32'hbf10c9a1} /* (24, 26, 7) {real, imag} */,
  {32'hbf65bf77, 32'hbee318a0} /* (24, 26, 6) {real, imag} */,
  {32'hbd11848c, 32'h3cb3a7c0} /* (24, 26, 5) {real, imag} */,
  {32'h3f21d446, 32'hbf29c722} /* (24, 26, 4) {real, imag} */,
  {32'hbe828e68, 32'h3ec39cf5} /* (24, 26, 3) {real, imag} */,
  {32'hbe628d1e, 32'hbef450aa} /* (24, 26, 2) {real, imag} */,
  {32'h3ea7404c, 32'h3e1de668} /* (24, 26, 1) {real, imag} */,
  {32'hbd94d688, 32'h3e0ee3cc} /* (24, 26, 0) {real, imag} */,
  {32'hbf4e74de, 32'h3f7477c7} /* (24, 25, 31) {real, imag} */,
  {32'hbc7c3f30, 32'hbf83b6c0} /* (24, 25, 30) {real, imag} */,
  {32'hbf0363fa, 32'hbf304c2c} /* (24, 25, 29) {real, imag} */,
  {32'h3e84a084, 32'h3d5c8cab} /* (24, 25, 28) {real, imag} */,
  {32'hbe95c452, 32'hbed4f8c1} /* (24, 25, 27) {real, imag} */,
  {32'h3cba2f40, 32'h3e075817} /* (24, 25, 26) {real, imag} */,
  {32'hbe6b2600, 32'h3ecde22a} /* (24, 25, 25) {real, imag} */,
  {32'h3e7c305a, 32'hbf826b74} /* (24, 25, 24) {real, imag} */,
  {32'h3f010876, 32'h3d7a1908} /* (24, 25, 23) {real, imag} */,
  {32'hbeb6deb8, 32'hbf331fa9} /* (24, 25, 22) {real, imag} */,
  {32'hbe0d0b2b, 32'hbdda5912} /* (24, 25, 21) {real, imag} */,
  {32'h3eba12ba, 32'hbe9800a2} /* (24, 25, 20) {real, imag} */,
  {32'h3ed4befa, 32'h3d55d662} /* (24, 25, 19) {real, imag} */,
  {32'h3f11d8fa, 32'hbecaea74} /* (24, 25, 18) {real, imag} */,
  {32'hbe2d6530, 32'hbe772870} /* (24, 25, 17) {real, imag} */,
  {32'hbe1015ad, 32'h3e3c8549} /* (24, 25, 16) {real, imag} */,
  {32'h3e97384d, 32'h3e673fb3} /* (24, 25, 15) {real, imag} */,
  {32'hbeff155e, 32'hbd2da0f4} /* (24, 25, 14) {real, imag} */,
  {32'hbe654f6c, 32'hbe339b78} /* (24, 25, 13) {real, imag} */,
  {32'h3d90c83f, 32'hbede7e2c} /* (24, 25, 12) {real, imag} */,
  {32'hbf131e78, 32'h3db83abc} /* (24, 25, 11) {real, imag} */,
  {32'hbd8f8e96, 32'h3df1a820} /* (24, 25, 10) {real, imag} */,
  {32'h3f2675bf, 32'hbeb15da0} /* (24, 25, 9) {real, imag} */,
  {32'h3ea68770, 32'hbeab7aa4} /* (24, 25, 8) {real, imag} */,
  {32'h3e47b414, 32'hbedec1aa} /* (24, 25, 7) {real, imag} */,
  {32'hbe6d6f4d, 32'h3f6afd46} /* (24, 25, 6) {real, imag} */,
  {32'hbec289f5, 32'hbda42070} /* (24, 25, 5) {real, imag} */,
  {32'hbf00d10b, 32'h3ec4eefd} /* (24, 25, 4) {real, imag} */,
  {32'hbea31d50, 32'hbe275ee3} /* (24, 25, 3) {real, imag} */,
  {32'h3e026bdc, 32'hbe98e15e} /* (24, 25, 2) {real, imag} */,
  {32'hbf76203b, 32'hbc4a1e40} /* (24, 25, 1) {real, imag} */,
  {32'hbf182442, 32'h3ea70262} /* (24, 25, 0) {real, imag} */,
  {32'h3f92f4bd, 32'hbf1e7531} /* (24, 24, 31) {real, imag} */,
  {32'hbf75980a, 32'h3ef83853} /* (24, 24, 30) {real, imag} */,
  {32'hbef48a33, 32'h3eb8e8c0} /* (24, 24, 29) {real, imag} */,
  {32'h3f1a0965, 32'h3cd1fdf0} /* (24, 24, 28) {real, imag} */,
  {32'hbf1fe7d8, 32'h3e2c280d} /* (24, 24, 27) {real, imag} */,
  {32'h3eef4b3e, 32'h3eff90bd} /* (24, 24, 26) {real, imag} */,
  {32'h3d415558, 32'h3ed9cfe2} /* (24, 24, 25) {real, imag} */,
  {32'hbebc57cc, 32'h3eb5a0d7} /* (24, 24, 24) {real, imag} */,
  {32'hbe1808df, 32'hbe762e16} /* (24, 24, 23) {real, imag} */,
  {32'hbdc4c118, 32'hbd96ab60} /* (24, 24, 22) {real, imag} */,
  {32'h3dd3779f, 32'hbe39c296} /* (24, 24, 21) {real, imag} */,
  {32'h3ea455d0, 32'h3e65f22e} /* (24, 24, 20) {real, imag} */,
  {32'h3e834d81, 32'h3d6d91fc} /* (24, 24, 19) {real, imag} */,
  {32'hbda20cf6, 32'hbe870902} /* (24, 24, 18) {real, imag} */,
  {32'h3e0fbca5, 32'hbe17b9b1} /* (24, 24, 17) {real, imag} */,
  {32'hbc301240, 32'h3ea5a4be} /* (24, 24, 16) {real, imag} */,
  {32'h3da1087a, 32'hbd9e3d86} /* (24, 24, 15) {real, imag} */,
  {32'h3d3dc57c, 32'hbcd27c88} /* (24, 24, 14) {real, imag} */,
  {32'hbe16cfd5, 32'hbe16372a} /* (24, 24, 13) {real, imag} */,
  {32'h3e6d8fe1, 32'hbec9a799} /* (24, 24, 12) {real, imag} */,
  {32'h3cea3504, 32'hbf00678e} /* (24, 24, 11) {real, imag} */,
  {32'hbc943b35, 32'hbee9c6b8} /* (24, 24, 10) {real, imag} */,
  {32'h3c2a2c7c, 32'hbebf9592} /* (24, 24, 9) {real, imag} */,
  {32'hbde12076, 32'h3ee6ae6b} /* (24, 24, 8) {real, imag} */,
  {32'h3f13ccb2, 32'h3f423c84} /* (24, 24, 7) {real, imag} */,
  {32'h3e940d74, 32'h3f15afd0} /* (24, 24, 6) {real, imag} */,
  {32'hbefcf1e8, 32'hbec6e3bc} /* (24, 24, 5) {real, imag} */,
  {32'h3ec94199, 32'h3e325374} /* (24, 24, 4) {real, imag} */,
  {32'h3e0c7710, 32'hbdf48fed} /* (24, 24, 3) {real, imag} */,
  {32'hbf4f68e0, 32'h3e91f9a2} /* (24, 24, 2) {real, imag} */,
  {32'h3fbea0ad, 32'hbf37e9ca} /* (24, 24, 1) {real, imag} */,
  {32'h3dbe2992, 32'hbea422e0} /* (24, 24, 0) {real, imag} */,
  {32'hbf94bd6a, 32'hbcafb200} /* (24, 23, 31) {real, imag} */,
  {32'h39c09d00, 32'hbdd6d3b0} /* (24, 23, 30) {real, imag} */,
  {32'h3b1a5fa0, 32'h3f1945a3} /* (24, 23, 29) {real, imag} */,
  {32'hbe06f494, 32'h3e3ea6ca} /* (24, 23, 28) {real, imag} */,
  {32'h3e981b3f, 32'hbe478497} /* (24, 23, 27) {real, imag} */,
  {32'h3eb0991c, 32'hbdc4bb36} /* (24, 23, 26) {real, imag} */,
  {32'hbefa4be0, 32'hbe2b0c5c} /* (24, 23, 25) {real, imag} */,
  {32'hbe79c855, 32'hbe1f3391} /* (24, 23, 24) {real, imag} */,
  {32'hbe303e2e, 32'h3cb2c678} /* (24, 23, 23) {real, imag} */,
  {32'hbe31215f, 32'hbef2cc30} /* (24, 23, 22) {real, imag} */,
  {32'hbea29b35, 32'h3a9032c0} /* (24, 23, 21) {real, imag} */,
  {32'hbdd08558, 32'h3e12f3f2} /* (24, 23, 20) {real, imag} */,
  {32'hbe55b216, 32'h3daae604} /* (24, 23, 19) {real, imag} */,
  {32'hbeb15790, 32'hbe717428} /* (24, 23, 18) {real, imag} */,
  {32'h3db5411c, 32'h3d8f8e60} /* (24, 23, 17) {real, imag} */,
  {32'hbd923430, 32'h3f09b418} /* (24, 23, 16) {real, imag} */,
  {32'hbde6dbc3, 32'h3e7c1b06} /* (24, 23, 15) {real, imag} */,
  {32'hbbfd56c0, 32'hbed7e0d0} /* (24, 23, 14) {real, imag} */,
  {32'h3ea109a5, 32'hbe854a9e} /* (24, 23, 13) {real, imag} */,
  {32'h3dc8896c, 32'h3e0274a1} /* (24, 23, 12) {real, imag} */,
  {32'h3ce0a6fc, 32'h3ea9ac20} /* (24, 23, 11) {real, imag} */,
  {32'h3e7fd569, 32'h3dfebdc9} /* (24, 23, 10) {real, imag} */,
  {32'hbf0c6f1b, 32'h3e7a9d9c} /* (24, 23, 9) {real, imag} */,
  {32'hbd823e49, 32'hbd81099c} /* (24, 23, 8) {real, imag} */,
  {32'hbd1be4ca, 32'h3d7a5898} /* (24, 23, 7) {real, imag} */,
  {32'hbecc16d0, 32'hbddb5f3e} /* (24, 23, 6) {real, imag} */,
  {32'h3f1e404f, 32'hbf42193e} /* (24, 23, 5) {real, imag} */,
  {32'h3e7b9904, 32'hbd1bc604} /* (24, 23, 4) {real, imag} */,
  {32'h3e75eb89, 32'h3edaff92} /* (24, 23, 3) {real, imag} */,
  {32'hbeb66cbe, 32'hbf1d4058} /* (24, 23, 2) {real, imag} */,
  {32'h3dee9c08, 32'h3eab8bb6} /* (24, 23, 1) {real, imag} */,
  {32'h3cb079d0, 32'h3dfe9448} /* (24, 23, 0) {real, imag} */,
  {32'hbe92045a, 32'h3f1c347a} /* (24, 22, 31) {real, imag} */,
  {32'h3e928ae3, 32'h3e001d62} /* (24, 22, 30) {real, imag} */,
  {32'hbeaa3755, 32'h3d456079} /* (24, 22, 29) {real, imag} */,
  {32'h3dde68da, 32'h3e70e17a} /* (24, 22, 28) {real, imag} */,
  {32'h3cced038, 32'hbeaaccb4} /* (24, 22, 27) {real, imag} */,
  {32'hbf0d138d, 32'hbe857efa} /* (24, 22, 26) {real, imag} */,
  {32'h3ebadd4a, 32'h3e44a7b2} /* (24, 22, 25) {real, imag} */,
  {32'h3ec3f3cc, 32'h3f189c6b} /* (24, 22, 24) {real, imag} */,
  {32'hbdfddb80, 32'hbe0b1a43} /* (24, 22, 23) {real, imag} */,
  {32'hbedad57f, 32'h3e00304a} /* (24, 22, 22) {real, imag} */,
  {32'h3e178dae, 32'h3eacc08a} /* (24, 22, 21) {real, imag} */,
  {32'hbe839f4d, 32'hbefa25c8} /* (24, 22, 20) {real, imag} */,
  {32'h3e8ea27a, 32'hbeab0729} /* (24, 22, 19) {real, imag} */,
  {32'h3e3b774b, 32'h3ef0863e} /* (24, 22, 18) {real, imag} */,
  {32'hbe041bec, 32'hbf073266} /* (24, 22, 17) {real, imag} */,
  {32'hbd99db70, 32'h3e05d796} /* (24, 22, 16) {real, imag} */,
  {32'h3e1a63ba, 32'h3ed1e6ac} /* (24, 22, 15) {real, imag} */,
  {32'hbf32ed17, 32'hbd3eea62} /* (24, 22, 14) {real, imag} */,
  {32'hbe9a1510, 32'hbc6a5550} /* (24, 22, 13) {real, imag} */,
  {32'hbea4e66b, 32'hbe8b6dd9} /* (24, 22, 12) {real, imag} */,
  {32'h3eb40d0a, 32'h3f36ec60} /* (24, 22, 11) {real, imag} */,
  {32'hbc68ca30, 32'hbe1f082f} /* (24, 22, 10) {real, imag} */,
  {32'h3f001bfe, 32'h3ed5eefe} /* (24, 22, 9) {real, imag} */,
  {32'hbec43eb8, 32'h3dd89574} /* (24, 22, 8) {real, imag} */,
  {32'h3dcd92a8, 32'h3e31b27f} /* (24, 22, 7) {real, imag} */,
  {32'hbdfaa384, 32'h3f0583b0} /* (24, 22, 6) {real, imag} */,
  {32'h3e16cd40, 32'hbe9e5ace} /* (24, 22, 5) {real, imag} */,
  {32'hbf24bd3b, 32'h3e8d3c4a} /* (24, 22, 4) {real, imag} */,
  {32'hbf01d08a, 32'h3e4eeb42} /* (24, 22, 3) {real, imag} */,
  {32'hbce04be0, 32'hbf982f52} /* (24, 22, 2) {real, imag} */,
  {32'hbec80bb6, 32'h3f5e4132} /* (24, 22, 1) {real, imag} */,
  {32'hbe54c971, 32'h3f1ec9d3} /* (24, 22, 0) {real, imag} */,
  {32'h3db858b0, 32'hbf04702a} /* (24, 21, 31) {real, imag} */,
  {32'h3f124f42, 32'h3ebc856a} /* (24, 21, 30) {real, imag} */,
  {32'h3f5909b0, 32'hbd8aa81f} /* (24, 21, 29) {real, imag} */,
  {32'hbd90a0b0, 32'hbcb1699c} /* (24, 21, 28) {real, imag} */,
  {32'hbe69af4c, 32'h3e11bbc0} /* (24, 21, 27) {real, imag} */,
  {32'hbee11a50, 32'h3dee5f47} /* (24, 21, 26) {real, imag} */,
  {32'hbd20e374, 32'hbf5fc24e} /* (24, 21, 25) {real, imag} */,
  {32'hbe52021f, 32'h3ebea240} /* (24, 21, 24) {real, imag} */,
  {32'h3ecf2bc4, 32'h3eb94251} /* (24, 21, 23) {real, imag} */,
  {32'hbe3e1c88, 32'hbecbdd49} /* (24, 21, 22) {real, imag} */,
  {32'h3df0e3f9, 32'hbda5747e} /* (24, 21, 21) {real, imag} */,
  {32'h3e331fa0, 32'h3eb93168} /* (24, 21, 20) {real, imag} */,
  {32'hbb0c6f00, 32'h3ef2f065} /* (24, 21, 19) {real, imag} */,
  {32'h3ebd2ec0, 32'hbd945c36} /* (24, 21, 18) {real, imag} */,
  {32'hbe979c04, 32'hbeb384e4} /* (24, 21, 17) {real, imag} */,
  {32'h3f01bfa4, 32'hbe775f83} /* (24, 21, 16) {real, imag} */,
  {32'hbedf703c, 32'h3c9c2f38} /* (24, 21, 15) {real, imag} */,
  {32'h3dbd91c3, 32'h3d43caf6} /* (24, 21, 14) {real, imag} */,
  {32'hbd692e8a, 32'h3c723de0} /* (24, 21, 13) {real, imag} */,
  {32'h3c7c5250, 32'hbe61488e} /* (24, 21, 12) {real, imag} */,
  {32'h3e11b849, 32'hbf45bf44} /* (24, 21, 11) {real, imag} */,
  {32'h3e952c3b, 32'h3e29a86a} /* (24, 21, 10) {real, imag} */,
  {32'hbd7cd69b, 32'h3e004dc2} /* (24, 21, 9) {real, imag} */,
  {32'h3e3b12f7, 32'hbe7ca492} /* (24, 21, 8) {real, imag} */,
  {32'h3f158501, 32'h3ed470b2} /* (24, 21, 7) {real, imag} */,
  {32'hbd28ba10, 32'h3e882fd8} /* (24, 21, 6) {real, imag} */,
  {32'h3e654d04, 32'h3d4316dc} /* (24, 21, 5) {real, imag} */,
  {32'hbd37d342, 32'hbd248180} /* (24, 21, 4) {real, imag} */,
  {32'hbeb5840e, 32'hbdcb3a98} /* (24, 21, 3) {real, imag} */,
  {32'hbe7e4dd2, 32'h3f30a015} /* (24, 21, 2) {real, imag} */,
  {32'h3f4c71ec, 32'hbe81c8a6} /* (24, 21, 1) {real, imag} */,
  {32'h3e601e50, 32'hbed3983a} /* (24, 21, 0) {real, imag} */,
  {32'h3d3a5a0c, 32'hbd9db146} /* (24, 20, 31) {real, imag} */,
  {32'hbe447a34, 32'h3c8b6c00} /* (24, 20, 30) {real, imag} */,
  {32'h3d3b02e1, 32'h3e3fb4d6} /* (24, 20, 29) {real, imag} */,
  {32'hbb324e80, 32'hbed422d8} /* (24, 20, 28) {real, imag} */,
  {32'h3d5aa0f8, 32'h3e4704f2} /* (24, 20, 27) {real, imag} */,
  {32'h3e48a023, 32'hbdc22a38} /* (24, 20, 26) {real, imag} */,
  {32'h3ef0bbe9, 32'hbe806952} /* (24, 20, 25) {real, imag} */,
  {32'hbe0c6f30, 32'hbe4c0da4} /* (24, 20, 24) {real, imag} */,
  {32'hbe8ac9ab, 32'h3ec0faec} /* (24, 20, 23) {real, imag} */,
  {32'hbf1cc2d6, 32'hbd8b2156} /* (24, 20, 22) {real, imag} */,
  {32'hbe547caf, 32'h3f0ace78} /* (24, 20, 21) {real, imag} */,
  {32'hbde876ca, 32'h3e26e40a} /* (24, 20, 20) {real, imag} */,
  {32'hbd89b3e4, 32'hbdfb5132} /* (24, 20, 19) {real, imag} */,
  {32'h3d49a7b6, 32'h3e2c6563} /* (24, 20, 18) {real, imag} */,
  {32'h3aa35d80, 32'h3edab6dc} /* (24, 20, 17) {real, imag} */,
  {32'h3d7a75b4, 32'hbd68f5df} /* (24, 20, 16) {real, imag} */,
  {32'h3e5c1436, 32'h3d1f7b66} /* (24, 20, 15) {real, imag} */,
  {32'hbe1e1ba4, 32'h3ecc7dd2} /* (24, 20, 14) {real, imag} */,
  {32'h3e575c7d, 32'hbd8908de} /* (24, 20, 13) {real, imag} */,
  {32'h3f476918, 32'h3e28039c} /* (24, 20, 12) {real, imag} */,
  {32'hbe4ed349, 32'hbda8e81e} /* (24, 20, 11) {real, imag} */,
  {32'h3d5ffd58, 32'hbedf1668} /* (24, 20, 10) {real, imag} */,
  {32'hbea4f667, 32'hbc923bc8} /* (24, 20, 9) {real, imag} */,
  {32'hbec681c4, 32'hbf122c55} /* (24, 20, 8) {real, imag} */,
  {32'hbb0d5e00, 32'h3e966a26} /* (24, 20, 7) {real, imag} */,
  {32'h3c2a48b0, 32'hbedfa9d0} /* (24, 20, 6) {real, imag} */,
  {32'hbec780ae, 32'h3f2b1b8c} /* (24, 20, 5) {real, imag} */,
  {32'h3ea64843, 32'h3e9d08ec} /* (24, 20, 4) {real, imag} */,
  {32'h3d1deb16, 32'h3dc06e2c} /* (24, 20, 3) {real, imag} */,
  {32'h3dfa99e0, 32'hbd839e31} /* (24, 20, 2) {real, imag} */,
  {32'hbebfa884, 32'hbeb5012d} /* (24, 20, 1) {real, imag} */,
  {32'h3f1b8a8c, 32'hbe73ea75} /* (24, 20, 0) {real, imag} */,
  {32'hbd9b6f24, 32'hbf0d3268} /* (24, 19, 31) {real, imag} */,
  {32'h3e5499b4, 32'h3ededa4a} /* (24, 19, 30) {real, imag} */,
  {32'h3e22bde8, 32'h3d097c98} /* (24, 19, 29) {real, imag} */,
  {32'hbefa2577, 32'h3f138afa} /* (24, 19, 28) {real, imag} */,
  {32'h3ef83d75, 32'h3ca4dd90} /* (24, 19, 27) {real, imag} */,
  {32'h3ec097b6, 32'hbe2d6860} /* (24, 19, 26) {real, imag} */,
  {32'h3e912ef1, 32'hbdd1b588} /* (24, 19, 25) {real, imag} */,
  {32'h3e6bb7d3, 32'hbdf559b2} /* (24, 19, 24) {real, imag} */,
  {32'h3df6a91a, 32'hbea295bb} /* (24, 19, 23) {real, imag} */,
  {32'h3e1f7ae2, 32'h3e1a3e78} /* (24, 19, 22) {real, imag} */,
  {32'h3dd16af3, 32'h3e7299a0} /* (24, 19, 21) {real, imag} */,
  {32'h3d2fb2de, 32'hbded7b4b} /* (24, 19, 20) {real, imag} */,
  {32'hbe461f6b, 32'hbcc1e5c0} /* (24, 19, 19) {real, imag} */,
  {32'hbeda21b4, 32'h3e75dd28} /* (24, 19, 18) {real, imag} */,
  {32'hbeb64b66, 32'hbd34bc6c} /* (24, 19, 17) {real, imag} */,
  {32'hbdeb5159, 32'hbe6b1194} /* (24, 19, 16) {real, imag} */,
  {32'h3e9a3447, 32'h3ea00188} /* (24, 19, 15) {real, imag} */,
  {32'hbddc5277, 32'hbbb2f610} /* (24, 19, 14) {real, imag} */,
  {32'h3ed3f967, 32'hbe968564} /* (24, 19, 13) {real, imag} */,
  {32'hbdb1b2ec, 32'h3f04923c} /* (24, 19, 12) {real, imag} */,
  {32'h3e72e8d2, 32'h3e490523} /* (24, 19, 11) {real, imag} */,
  {32'hbe9bed9a, 32'hbebb4c50} /* (24, 19, 10) {real, imag} */,
  {32'hbec973f2, 32'h3e4c1806} /* (24, 19, 9) {real, imag} */,
  {32'hbddbeb4e, 32'h3d6aa68e} /* (24, 19, 8) {real, imag} */,
  {32'hbe346cef, 32'hbf04a811} /* (24, 19, 7) {real, imag} */,
  {32'hbe29392e, 32'hbedb2eea} /* (24, 19, 6) {real, imag} */,
  {32'hbe1dda8e, 32'hbe672e82} /* (24, 19, 5) {real, imag} */,
  {32'hbe9db17d, 32'hbe594316} /* (24, 19, 4) {real, imag} */,
  {32'h3eab4f9f, 32'hbd82339c} /* (24, 19, 3) {real, imag} */,
  {32'hbe441cc4, 32'h3eaa2aca} /* (24, 19, 2) {real, imag} */,
  {32'hbf095488, 32'hbe405505} /* (24, 19, 1) {real, imag} */,
  {32'hbd58b280, 32'h3e48c809} /* (24, 19, 0) {real, imag} */,
  {32'hbd9fd9de, 32'hbe983f5e} /* (24, 18, 31) {real, imag} */,
  {32'hbe77994a, 32'h3ebbb441} /* (24, 18, 30) {real, imag} */,
  {32'h3db159f1, 32'hbd86dbae} /* (24, 18, 29) {real, imag} */,
  {32'h3b172f50, 32'hbc9a0cdc} /* (24, 18, 28) {real, imag} */,
  {32'hbea0df2b, 32'h3ed5225e} /* (24, 18, 27) {real, imag} */,
  {32'h3e4834e6, 32'h3d10435c} /* (24, 18, 26) {real, imag} */,
  {32'hbf06390e, 32'hbd8c8741} /* (24, 18, 25) {real, imag} */,
  {32'hbdd6c781, 32'h3ea9e3dc} /* (24, 18, 24) {real, imag} */,
  {32'h3ec095e9, 32'hbeba99ef} /* (24, 18, 23) {real, imag} */,
  {32'hbecafcfd, 32'hbe78f612} /* (24, 18, 22) {real, imag} */,
  {32'h3ea14010, 32'hbe518f34} /* (24, 18, 21) {real, imag} */,
  {32'hbdadbc2f, 32'hbcc881a8} /* (24, 18, 20) {real, imag} */,
  {32'hbe1f94f3, 32'hbd2cb50c} /* (24, 18, 19) {real, imag} */,
  {32'h3cb497b0, 32'h3d13ca24} /* (24, 18, 18) {real, imag} */,
  {32'hbd9486d8, 32'hbd295fc4} /* (24, 18, 17) {real, imag} */,
  {32'h3ea43521, 32'h3dd527f4} /* (24, 18, 16) {real, imag} */,
  {32'hbe863afc, 32'hbdf92380} /* (24, 18, 15) {real, imag} */,
  {32'hbe70f6d8, 32'hbec78d2c} /* (24, 18, 14) {real, imag} */,
  {32'h3e42a475, 32'h3e3eeb0a} /* (24, 18, 13) {real, imag} */,
  {32'hbe2a265c, 32'h3e038755} /* (24, 18, 12) {real, imag} */,
  {32'hbf0661a3, 32'h3dbc3f86} /* (24, 18, 11) {real, imag} */,
  {32'h3e369508, 32'h3d5da50c} /* (24, 18, 10) {real, imag} */,
  {32'h3ec5852e, 32'hbd1116f8} /* (24, 18, 9) {real, imag} */,
  {32'hbeba5d0a, 32'hbe17aa42} /* (24, 18, 8) {real, imag} */,
  {32'h3d8dc1ee, 32'h3a0531c0} /* (24, 18, 7) {real, imag} */,
  {32'hbe2332c8, 32'hbed106bc} /* (24, 18, 6) {real, imag} */,
  {32'h3db6262e, 32'h3d597088} /* (24, 18, 5) {real, imag} */,
  {32'h3f08c6b2, 32'h3ece6208} /* (24, 18, 4) {real, imag} */,
  {32'h3ee21400, 32'hbd113834} /* (24, 18, 3) {real, imag} */,
  {32'hbf20a493, 32'h3e2abf5c} /* (24, 18, 2) {real, imag} */,
  {32'h3e3b989f, 32'hbedc8a74} /* (24, 18, 1) {real, imag} */,
  {32'h3e8356ea, 32'hbdfd10e6} /* (24, 18, 0) {real, imag} */,
  {32'hbb2a5e90, 32'hbd23c850} /* (24, 17, 31) {real, imag} */,
  {32'hbe2c079f, 32'hbe4fe5fd} /* (24, 17, 30) {real, imag} */,
  {32'hbe975e34, 32'hbe3ec5bc} /* (24, 17, 29) {real, imag} */,
  {32'h3e87c13c, 32'h3e828813} /* (24, 17, 28) {real, imag} */,
  {32'h3aaa4100, 32'hbc3ca7a0} /* (24, 17, 27) {real, imag} */,
  {32'hbcb35200, 32'h3e8b3ba2} /* (24, 17, 26) {real, imag} */,
  {32'hbe30e526, 32'hbecb15b2} /* (24, 17, 25) {real, imag} */,
  {32'h3e550642, 32'hbd277960} /* (24, 17, 24) {real, imag} */,
  {32'hbf09185a, 32'hbe0d4442} /* (24, 17, 23) {real, imag} */,
  {32'hbe836360, 32'h3e93a241} /* (24, 17, 22) {real, imag} */,
  {32'h3ebafad6, 32'hbf046e95} /* (24, 17, 21) {real, imag} */,
  {32'hbc80a88c, 32'h3daedbe0} /* (24, 17, 20) {real, imag} */,
  {32'h3e5850ce, 32'hbbde4040} /* (24, 17, 19) {real, imag} */,
  {32'h3e9200d2, 32'h3e0dff4b} /* (24, 17, 18) {real, imag} */,
  {32'hbdb17624, 32'hbdea5802} /* (24, 17, 17) {real, imag} */,
  {32'hbcf07d60, 32'h3d8e501e} /* (24, 17, 16) {real, imag} */,
  {32'hbd3760b8, 32'h3cdc0a40} /* (24, 17, 15) {real, imag} */,
  {32'hbe08a77a, 32'h3e1425b8} /* (24, 17, 14) {real, imag} */,
  {32'h3d9eb17f, 32'hbe0cd7f0} /* (24, 17, 13) {real, imag} */,
  {32'h3c63eaa8, 32'hbdac11ad} /* (24, 17, 12) {real, imag} */,
  {32'hbd835fc2, 32'hbe566a77} /* (24, 17, 11) {real, imag} */,
  {32'hbc8275d0, 32'h3e43c394} /* (24, 17, 10) {real, imag} */,
  {32'h3ec9335f, 32'h3e570928} /* (24, 17, 9) {real, imag} */,
  {32'h3e1dee31, 32'h3dc32bba} /* (24, 17, 8) {real, imag} */,
  {32'h3d3f76d4, 32'hbf148829} /* (24, 17, 7) {real, imag} */,
  {32'h3e16b012, 32'hbea43290} /* (24, 17, 6) {real, imag} */,
  {32'hbc1a3fa4, 32'h3d9df903} /* (24, 17, 5) {real, imag} */,
  {32'hbe19ee8c, 32'h3d3c5b47} /* (24, 17, 4) {real, imag} */,
  {32'hbea01314, 32'h3e19370c} /* (24, 17, 3) {real, imag} */,
  {32'h3e81e38f, 32'hbd3fed4c} /* (24, 17, 2) {real, imag} */,
  {32'hbd0315e7, 32'h3d076098} /* (24, 17, 1) {real, imag} */,
  {32'hbd9ac802, 32'h3e61093a} /* (24, 17, 0) {real, imag} */,
  {32'h3e58811a, 32'hbb4f2c60} /* (24, 16, 31) {real, imag} */,
  {32'h3df460aa, 32'hbd943ba8} /* (24, 16, 30) {real, imag} */,
  {32'hbe30b48b, 32'h3dd32096} /* (24, 16, 29) {real, imag} */,
  {32'h3d42c97c, 32'h3d3a561a} /* (24, 16, 28) {real, imag} */,
  {32'hbe622ab7, 32'hbe6badab} /* (24, 16, 27) {real, imag} */,
  {32'h3dd16367, 32'hbec57bd1} /* (24, 16, 26) {real, imag} */,
  {32'h3e9c54a8, 32'h3e0a0896} /* (24, 16, 25) {real, imag} */,
  {32'h3e6310f4, 32'h3eb55262} /* (24, 16, 24) {real, imag} */,
  {32'h3cfd5e40, 32'h3ee49adc} /* (24, 16, 23) {real, imag} */,
  {32'hbeccf9fb, 32'hbe1ce1fe} /* (24, 16, 22) {real, imag} */,
  {32'hba31cd00, 32'h3e032f6d} /* (24, 16, 21) {real, imag} */,
  {32'h3e01ce9a, 32'hbe198052} /* (24, 16, 20) {real, imag} */,
  {32'h3dd642a4, 32'hbdcc8054} /* (24, 16, 19) {real, imag} */,
  {32'hbdc7aa54, 32'hbe082b0f} /* (24, 16, 18) {real, imag} */,
  {32'hbe807c81, 32'hbe2383f8} /* (24, 16, 17) {real, imag} */,
  {32'hbe2a69bc, 32'h00000000} /* (24, 16, 16) {real, imag} */,
  {32'hbe807c81, 32'h3e2383f8} /* (24, 16, 15) {real, imag} */,
  {32'hbdc7aa54, 32'h3e082b0f} /* (24, 16, 14) {real, imag} */,
  {32'h3dd642a4, 32'h3dcc8054} /* (24, 16, 13) {real, imag} */,
  {32'h3e01ce9a, 32'h3e198052} /* (24, 16, 12) {real, imag} */,
  {32'hba31cd00, 32'hbe032f6d} /* (24, 16, 11) {real, imag} */,
  {32'hbeccf9fb, 32'h3e1ce1fe} /* (24, 16, 10) {real, imag} */,
  {32'h3cfd5e40, 32'hbee49adc} /* (24, 16, 9) {real, imag} */,
  {32'h3e6310f4, 32'hbeb55262} /* (24, 16, 8) {real, imag} */,
  {32'h3e9c54a8, 32'hbe0a0896} /* (24, 16, 7) {real, imag} */,
  {32'h3dd16367, 32'h3ec57bd1} /* (24, 16, 6) {real, imag} */,
  {32'hbe622ab7, 32'h3e6badab} /* (24, 16, 5) {real, imag} */,
  {32'h3d42c97c, 32'hbd3a561a} /* (24, 16, 4) {real, imag} */,
  {32'hbe30b48b, 32'hbdd32096} /* (24, 16, 3) {real, imag} */,
  {32'h3df460aa, 32'h3d943ba8} /* (24, 16, 2) {real, imag} */,
  {32'h3e58811a, 32'h3b4f2c60} /* (24, 16, 1) {real, imag} */,
  {32'hbdab64c0, 32'h00000000} /* (24, 16, 0) {real, imag} */,
  {32'hbd0315e7, 32'hbd076098} /* (24, 15, 31) {real, imag} */,
  {32'h3e81e38f, 32'h3d3fed4c} /* (24, 15, 30) {real, imag} */,
  {32'hbea01314, 32'hbe19370c} /* (24, 15, 29) {real, imag} */,
  {32'hbe19ee8c, 32'hbd3c5b47} /* (24, 15, 28) {real, imag} */,
  {32'hbc1a3fa4, 32'hbd9df903} /* (24, 15, 27) {real, imag} */,
  {32'h3e16b012, 32'h3ea43290} /* (24, 15, 26) {real, imag} */,
  {32'h3d3f76d4, 32'h3f148829} /* (24, 15, 25) {real, imag} */,
  {32'h3e1dee31, 32'hbdc32bba} /* (24, 15, 24) {real, imag} */,
  {32'h3ec9335f, 32'hbe570928} /* (24, 15, 23) {real, imag} */,
  {32'hbc8275d0, 32'hbe43c394} /* (24, 15, 22) {real, imag} */,
  {32'hbd835fc2, 32'h3e566a77} /* (24, 15, 21) {real, imag} */,
  {32'h3c63eaa8, 32'h3dac11ad} /* (24, 15, 20) {real, imag} */,
  {32'h3d9eb17f, 32'h3e0cd7f0} /* (24, 15, 19) {real, imag} */,
  {32'hbe08a77a, 32'hbe1425b8} /* (24, 15, 18) {real, imag} */,
  {32'hbd3760b8, 32'hbcdc0a40} /* (24, 15, 17) {real, imag} */,
  {32'hbcf07d60, 32'hbd8e501e} /* (24, 15, 16) {real, imag} */,
  {32'hbdb17624, 32'h3dea5802} /* (24, 15, 15) {real, imag} */,
  {32'h3e9200d2, 32'hbe0dff4b} /* (24, 15, 14) {real, imag} */,
  {32'h3e5850ce, 32'h3bde4040} /* (24, 15, 13) {real, imag} */,
  {32'hbc80a88c, 32'hbdaedbe0} /* (24, 15, 12) {real, imag} */,
  {32'h3ebafad6, 32'h3f046e95} /* (24, 15, 11) {real, imag} */,
  {32'hbe836360, 32'hbe93a241} /* (24, 15, 10) {real, imag} */,
  {32'hbf09185a, 32'h3e0d4442} /* (24, 15, 9) {real, imag} */,
  {32'h3e550642, 32'h3d277960} /* (24, 15, 8) {real, imag} */,
  {32'hbe30e526, 32'h3ecb15b2} /* (24, 15, 7) {real, imag} */,
  {32'hbcb35200, 32'hbe8b3ba2} /* (24, 15, 6) {real, imag} */,
  {32'h3aaa4100, 32'h3c3ca7a0} /* (24, 15, 5) {real, imag} */,
  {32'h3e87c13c, 32'hbe828813} /* (24, 15, 4) {real, imag} */,
  {32'hbe975e34, 32'h3e3ec5bc} /* (24, 15, 3) {real, imag} */,
  {32'hbe2c079f, 32'h3e4fe5fd} /* (24, 15, 2) {real, imag} */,
  {32'hbb2a5e90, 32'h3d23c850} /* (24, 15, 1) {real, imag} */,
  {32'hbd9ac802, 32'hbe61093a} /* (24, 15, 0) {real, imag} */,
  {32'h3e3b989f, 32'h3edc8a74} /* (24, 14, 31) {real, imag} */,
  {32'hbf20a493, 32'hbe2abf5c} /* (24, 14, 30) {real, imag} */,
  {32'h3ee21400, 32'h3d113834} /* (24, 14, 29) {real, imag} */,
  {32'h3f08c6b2, 32'hbece6208} /* (24, 14, 28) {real, imag} */,
  {32'h3db6262e, 32'hbd597088} /* (24, 14, 27) {real, imag} */,
  {32'hbe2332c8, 32'h3ed106bc} /* (24, 14, 26) {real, imag} */,
  {32'h3d8dc1ee, 32'hba0531c0} /* (24, 14, 25) {real, imag} */,
  {32'hbeba5d0a, 32'h3e17aa42} /* (24, 14, 24) {real, imag} */,
  {32'h3ec5852e, 32'h3d1116f8} /* (24, 14, 23) {real, imag} */,
  {32'h3e369508, 32'hbd5da50c} /* (24, 14, 22) {real, imag} */,
  {32'hbf0661a3, 32'hbdbc3f86} /* (24, 14, 21) {real, imag} */,
  {32'hbe2a265c, 32'hbe038755} /* (24, 14, 20) {real, imag} */,
  {32'h3e42a475, 32'hbe3eeb0a} /* (24, 14, 19) {real, imag} */,
  {32'hbe70f6d8, 32'h3ec78d2c} /* (24, 14, 18) {real, imag} */,
  {32'hbe863afc, 32'h3df92380} /* (24, 14, 17) {real, imag} */,
  {32'h3ea43521, 32'hbdd527f4} /* (24, 14, 16) {real, imag} */,
  {32'hbd9486d8, 32'h3d295fc4} /* (24, 14, 15) {real, imag} */,
  {32'h3cb497b0, 32'hbd13ca24} /* (24, 14, 14) {real, imag} */,
  {32'hbe1f94f3, 32'h3d2cb50c} /* (24, 14, 13) {real, imag} */,
  {32'hbdadbc2f, 32'h3cc881a8} /* (24, 14, 12) {real, imag} */,
  {32'h3ea14010, 32'h3e518f34} /* (24, 14, 11) {real, imag} */,
  {32'hbecafcfd, 32'h3e78f612} /* (24, 14, 10) {real, imag} */,
  {32'h3ec095e9, 32'h3eba99ef} /* (24, 14, 9) {real, imag} */,
  {32'hbdd6c781, 32'hbea9e3dc} /* (24, 14, 8) {real, imag} */,
  {32'hbf06390e, 32'h3d8c8741} /* (24, 14, 7) {real, imag} */,
  {32'h3e4834e6, 32'hbd10435c} /* (24, 14, 6) {real, imag} */,
  {32'hbea0df2b, 32'hbed5225e} /* (24, 14, 5) {real, imag} */,
  {32'h3b172f50, 32'h3c9a0cdc} /* (24, 14, 4) {real, imag} */,
  {32'h3db159f1, 32'h3d86dbae} /* (24, 14, 3) {real, imag} */,
  {32'hbe77994a, 32'hbebbb441} /* (24, 14, 2) {real, imag} */,
  {32'hbd9fd9de, 32'h3e983f5e} /* (24, 14, 1) {real, imag} */,
  {32'h3e8356ea, 32'h3dfd10e6} /* (24, 14, 0) {real, imag} */,
  {32'hbf095488, 32'h3e405505} /* (24, 13, 31) {real, imag} */,
  {32'hbe441cc4, 32'hbeaa2aca} /* (24, 13, 30) {real, imag} */,
  {32'h3eab4f9f, 32'h3d82339c} /* (24, 13, 29) {real, imag} */,
  {32'hbe9db17d, 32'h3e594316} /* (24, 13, 28) {real, imag} */,
  {32'hbe1dda8e, 32'h3e672e82} /* (24, 13, 27) {real, imag} */,
  {32'hbe29392e, 32'h3edb2eea} /* (24, 13, 26) {real, imag} */,
  {32'hbe346cef, 32'h3f04a811} /* (24, 13, 25) {real, imag} */,
  {32'hbddbeb4e, 32'hbd6aa68e} /* (24, 13, 24) {real, imag} */,
  {32'hbec973f2, 32'hbe4c1806} /* (24, 13, 23) {real, imag} */,
  {32'hbe9bed9a, 32'h3ebb4c50} /* (24, 13, 22) {real, imag} */,
  {32'h3e72e8d2, 32'hbe490523} /* (24, 13, 21) {real, imag} */,
  {32'hbdb1b2ec, 32'hbf04923c} /* (24, 13, 20) {real, imag} */,
  {32'h3ed3f967, 32'h3e968564} /* (24, 13, 19) {real, imag} */,
  {32'hbddc5277, 32'h3bb2f610} /* (24, 13, 18) {real, imag} */,
  {32'h3e9a3447, 32'hbea00188} /* (24, 13, 17) {real, imag} */,
  {32'hbdeb5159, 32'h3e6b1194} /* (24, 13, 16) {real, imag} */,
  {32'hbeb64b66, 32'h3d34bc6c} /* (24, 13, 15) {real, imag} */,
  {32'hbeda21b4, 32'hbe75dd28} /* (24, 13, 14) {real, imag} */,
  {32'hbe461f6b, 32'h3cc1e5c0} /* (24, 13, 13) {real, imag} */,
  {32'h3d2fb2de, 32'h3ded7b4b} /* (24, 13, 12) {real, imag} */,
  {32'h3dd16af3, 32'hbe7299a0} /* (24, 13, 11) {real, imag} */,
  {32'h3e1f7ae2, 32'hbe1a3e78} /* (24, 13, 10) {real, imag} */,
  {32'h3df6a91a, 32'h3ea295bb} /* (24, 13, 9) {real, imag} */,
  {32'h3e6bb7d3, 32'h3df559b2} /* (24, 13, 8) {real, imag} */,
  {32'h3e912ef1, 32'h3dd1b588} /* (24, 13, 7) {real, imag} */,
  {32'h3ec097b6, 32'h3e2d6860} /* (24, 13, 6) {real, imag} */,
  {32'h3ef83d75, 32'hbca4dd90} /* (24, 13, 5) {real, imag} */,
  {32'hbefa2577, 32'hbf138afa} /* (24, 13, 4) {real, imag} */,
  {32'h3e22bde8, 32'hbd097c98} /* (24, 13, 3) {real, imag} */,
  {32'h3e5499b4, 32'hbededa4a} /* (24, 13, 2) {real, imag} */,
  {32'hbd9b6f24, 32'h3f0d3268} /* (24, 13, 1) {real, imag} */,
  {32'hbd58b280, 32'hbe48c809} /* (24, 13, 0) {real, imag} */,
  {32'hbebfa884, 32'h3eb5012d} /* (24, 12, 31) {real, imag} */,
  {32'h3dfa99e0, 32'h3d839e31} /* (24, 12, 30) {real, imag} */,
  {32'h3d1deb16, 32'hbdc06e2c} /* (24, 12, 29) {real, imag} */,
  {32'h3ea64843, 32'hbe9d08ec} /* (24, 12, 28) {real, imag} */,
  {32'hbec780ae, 32'hbf2b1b8c} /* (24, 12, 27) {real, imag} */,
  {32'h3c2a48b0, 32'h3edfa9d0} /* (24, 12, 26) {real, imag} */,
  {32'hbb0d5e00, 32'hbe966a26} /* (24, 12, 25) {real, imag} */,
  {32'hbec681c4, 32'h3f122c55} /* (24, 12, 24) {real, imag} */,
  {32'hbea4f667, 32'h3c923bc8} /* (24, 12, 23) {real, imag} */,
  {32'h3d5ffd58, 32'h3edf1668} /* (24, 12, 22) {real, imag} */,
  {32'hbe4ed349, 32'h3da8e81e} /* (24, 12, 21) {real, imag} */,
  {32'h3f476918, 32'hbe28039c} /* (24, 12, 20) {real, imag} */,
  {32'h3e575c7d, 32'h3d8908de} /* (24, 12, 19) {real, imag} */,
  {32'hbe1e1ba4, 32'hbecc7dd2} /* (24, 12, 18) {real, imag} */,
  {32'h3e5c1436, 32'hbd1f7b66} /* (24, 12, 17) {real, imag} */,
  {32'h3d7a75b4, 32'h3d68f5df} /* (24, 12, 16) {real, imag} */,
  {32'h3aa35d80, 32'hbedab6dc} /* (24, 12, 15) {real, imag} */,
  {32'h3d49a7b6, 32'hbe2c6563} /* (24, 12, 14) {real, imag} */,
  {32'hbd89b3e4, 32'h3dfb5132} /* (24, 12, 13) {real, imag} */,
  {32'hbde876ca, 32'hbe26e40a} /* (24, 12, 12) {real, imag} */,
  {32'hbe547caf, 32'hbf0ace78} /* (24, 12, 11) {real, imag} */,
  {32'hbf1cc2d6, 32'h3d8b2156} /* (24, 12, 10) {real, imag} */,
  {32'hbe8ac9ab, 32'hbec0faec} /* (24, 12, 9) {real, imag} */,
  {32'hbe0c6f30, 32'h3e4c0da4} /* (24, 12, 8) {real, imag} */,
  {32'h3ef0bbe9, 32'h3e806952} /* (24, 12, 7) {real, imag} */,
  {32'h3e48a023, 32'h3dc22a38} /* (24, 12, 6) {real, imag} */,
  {32'h3d5aa0f8, 32'hbe4704f2} /* (24, 12, 5) {real, imag} */,
  {32'hbb324e80, 32'h3ed422d8} /* (24, 12, 4) {real, imag} */,
  {32'h3d3b02e1, 32'hbe3fb4d6} /* (24, 12, 3) {real, imag} */,
  {32'hbe447a34, 32'hbc8b6c00} /* (24, 12, 2) {real, imag} */,
  {32'h3d3a5a0c, 32'h3d9db146} /* (24, 12, 1) {real, imag} */,
  {32'h3f1b8a8c, 32'h3e73ea75} /* (24, 12, 0) {real, imag} */,
  {32'h3f4c71ec, 32'h3e81c8a6} /* (24, 11, 31) {real, imag} */,
  {32'hbe7e4dd2, 32'hbf30a015} /* (24, 11, 30) {real, imag} */,
  {32'hbeb5840e, 32'h3dcb3a98} /* (24, 11, 29) {real, imag} */,
  {32'hbd37d342, 32'h3d248180} /* (24, 11, 28) {real, imag} */,
  {32'h3e654d04, 32'hbd4316dc} /* (24, 11, 27) {real, imag} */,
  {32'hbd28ba10, 32'hbe882fd8} /* (24, 11, 26) {real, imag} */,
  {32'h3f158501, 32'hbed470b2} /* (24, 11, 25) {real, imag} */,
  {32'h3e3b12f7, 32'h3e7ca492} /* (24, 11, 24) {real, imag} */,
  {32'hbd7cd69b, 32'hbe004dc2} /* (24, 11, 23) {real, imag} */,
  {32'h3e952c3b, 32'hbe29a86a} /* (24, 11, 22) {real, imag} */,
  {32'h3e11b849, 32'h3f45bf44} /* (24, 11, 21) {real, imag} */,
  {32'h3c7c5250, 32'h3e61488e} /* (24, 11, 20) {real, imag} */,
  {32'hbd692e8a, 32'hbc723de0} /* (24, 11, 19) {real, imag} */,
  {32'h3dbd91c3, 32'hbd43caf6} /* (24, 11, 18) {real, imag} */,
  {32'hbedf703c, 32'hbc9c2f38} /* (24, 11, 17) {real, imag} */,
  {32'h3f01bfa4, 32'h3e775f83} /* (24, 11, 16) {real, imag} */,
  {32'hbe979c04, 32'h3eb384e4} /* (24, 11, 15) {real, imag} */,
  {32'h3ebd2ec0, 32'h3d945c36} /* (24, 11, 14) {real, imag} */,
  {32'hbb0c6f00, 32'hbef2f065} /* (24, 11, 13) {real, imag} */,
  {32'h3e331fa0, 32'hbeb93168} /* (24, 11, 12) {real, imag} */,
  {32'h3df0e3f9, 32'h3da5747e} /* (24, 11, 11) {real, imag} */,
  {32'hbe3e1c88, 32'h3ecbdd49} /* (24, 11, 10) {real, imag} */,
  {32'h3ecf2bc4, 32'hbeb94251} /* (24, 11, 9) {real, imag} */,
  {32'hbe52021f, 32'hbebea240} /* (24, 11, 8) {real, imag} */,
  {32'hbd20e374, 32'h3f5fc24e} /* (24, 11, 7) {real, imag} */,
  {32'hbee11a50, 32'hbdee5f47} /* (24, 11, 6) {real, imag} */,
  {32'hbe69af4c, 32'hbe11bbc0} /* (24, 11, 5) {real, imag} */,
  {32'hbd90a0b0, 32'h3cb1699c} /* (24, 11, 4) {real, imag} */,
  {32'h3f5909b0, 32'h3d8aa81f} /* (24, 11, 3) {real, imag} */,
  {32'h3f124f42, 32'hbebc856a} /* (24, 11, 2) {real, imag} */,
  {32'h3db858b0, 32'h3f04702a} /* (24, 11, 1) {real, imag} */,
  {32'h3e601e50, 32'h3ed3983a} /* (24, 11, 0) {real, imag} */,
  {32'hbec80bb6, 32'hbf5e4132} /* (24, 10, 31) {real, imag} */,
  {32'hbce04be0, 32'h3f982f52} /* (24, 10, 30) {real, imag} */,
  {32'hbf01d08a, 32'hbe4eeb42} /* (24, 10, 29) {real, imag} */,
  {32'hbf24bd3b, 32'hbe8d3c4a} /* (24, 10, 28) {real, imag} */,
  {32'h3e16cd40, 32'h3e9e5ace} /* (24, 10, 27) {real, imag} */,
  {32'hbdfaa384, 32'hbf0583b0} /* (24, 10, 26) {real, imag} */,
  {32'h3dcd92a8, 32'hbe31b27f} /* (24, 10, 25) {real, imag} */,
  {32'hbec43eb8, 32'hbdd89574} /* (24, 10, 24) {real, imag} */,
  {32'h3f001bfe, 32'hbed5eefe} /* (24, 10, 23) {real, imag} */,
  {32'hbc68ca30, 32'h3e1f082f} /* (24, 10, 22) {real, imag} */,
  {32'h3eb40d0a, 32'hbf36ec60} /* (24, 10, 21) {real, imag} */,
  {32'hbea4e66b, 32'h3e8b6dd9} /* (24, 10, 20) {real, imag} */,
  {32'hbe9a1510, 32'h3c6a5550} /* (24, 10, 19) {real, imag} */,
  {32'hbf32ed17, 32'h3d3eea62} /* (24, 10, 18) {real, imag} */,
  {32'h3e1a63ba, 32'hbed1e6ac} /* (24, 10, 17) {real, imag} */,
  {32'hbd99db70, 32'hbe05d796} /* (24, 10, 16) {real, imag} */,
  {32'hbe041bec, 32'h3f073266} /* (24, 10, 15) {real, imag} */,
  {32'h3e3b774b, 32'hbef0863e} /* (24, 10, 14) {real, imag} */,
  {32'h3e8ea27a, 32'h3eab0729} /* (24, 10, 13) {real, imag} */,
  {32'hbe839f4d, 32'h3efa25c8} /* (24, 10, 12) {real, imag} */,
  {32'h3e178dae, 32'hbeacc08a} /* (24, 10, 11) {real, imag} */,
  {32'hbedad57f, 32'hbe00304a} /* (24, 10, 10) {real, imag} */,
  {32'hbdfddb80, 32'h3e0b1a43} /* (24, 10, 9) {real, imag} */,
  {32'h3ec3f3cc, 32'hbf189c6b} /* (24, 10, 8) {real, imag} */,
  {32'h3ebadd4a, 32'hbe44a7b2} /* (24, 10, 7) {real, imag} */,
  {32'hbf0d138d, 32'h3e857efa} /* (24, 10, 6) {real, imag} */,
  {32'h3cced038, 32'h3eaaccb4} /* (24, 10, 5) {real, imag} */,
  {32'h3dde68da, 32'hbe70e17a} /* (24, 10, 4) {real, imag} */,
  {32'hbeaa3755, 32'hbd456079} /* (24, 10, 3) {real, imag} */,
  {32'h3e928ae3, 32'hbe001d62} /* (24, 10, 2) {real, imag} */,
  {32'hbe92045a, 32'hbf1c347a} /* (24, 10, 1) {real, imag} */,
  {32'hbe54c971, 32'hbf1ec9d3} /* (24, 10, 0) {real, imag} */,
  {32'h3dee9c08, 32'hbeab8bb6} /* (24, 9, 31) {real, imag} */,
  {32'hbeb66cbe, 32'h3f1d4058} /* (24, 9, 30) {real, imag} */,
  {32'h3e75eb89, 32'hbedaff92} /* (24, 9, 29) {real, imag} */,
  {32'h3e7b9904, 32'h3d1bc604} /* (24, 9, 28) {real, imag} */,
  {32'h3f1e404f, 32'h3f42193e} /* (24, 9, 27) {real, imag} */,
  {32'hbecc16d0, 32'h3ddb5f3e} /* (24, 9, 26) {real, imag} */,
  {32'hbd1be4ca, 32'hbd7a5898} /* (24, 9, 25) {real, imag} */,
  {32'hbd823e49, 32'h3d81099c} /* (24, 9, 24) {real, imag} */,
  {32'hbf0c6f1b, 32'hbe7a9d9c} /* (24, 9, 23) {real, imag} */,
  {32'h3e7fd569, 32'hbdfebdc9} /* (24, 9, 22) {real, imag} */,
  {32'h3ce0a6fc, 32'hbea9ac20} /* (24, 9, 21) {real, imag} */,
  {32'h3dc8896c, 32'hbe0274a1} /* (24, 9, 20) {real, imag} */,
  {32'h3ea109a5, 32'h3e854a9e} /* (24, 9, 19) {real, imag} */,
  {32'hbbfd56c0, 32'h3ed7e0d0} /* (24, 9, 18) {real, imag} */,
  {32'hbde6dbc3, 32'hbe7c1b06} /* (24, 9, 17) {real, imag} */,
  {32'hbd923430, 32'hbf09b418} /* (24, 9, 16) {real, imag} */,
  {32'h3db5411c, 32'hbd8f8e60} /* (24, 9, 15) {real, imag} */,
  {32'hbeb15790, 32'h3e717428} /* (24, 9, 14) {real, imag} */,
  {32'hbe55b216, 32'hbdaae604} /* (24, 9, 13) {real, imag} */,
  {32'hbdd08558, 32'hbe12f3f2} /* (24, 9, 12) {real, imag} */,
  {32'hbea29b35, 32'hba9032c0} /* (24, 9, 11) {real, imag} */,
  {32'hbe31215f, 32'h3ef2cc30} /* (24, 9, 10) {real, imag} */,
  {32'hbe303e2e, 32'hbcb2c678} /* (24, 9, 9) {real, imag} */,
  {32'hbe79c855, 32'h3e1f3391} /* (24, 9, 8) {real, imag} */,
  {32'hbefa4be0, 32'h3e2b0c5c} /* (24, 9, 7) {real, imag} */,
  {32'h3eb0991c, 32'h3dc4bb36} /* (24, 9, 6) {real, imag} */,
  {32'h3e981b3f, 32'h3e478497} /* (24, 9, 5) {real, imag} */,
  {32'hbe06f494, 32'hbe3ea6ca} /* (24, 9, 4) {real, imag} */,
  {32'h3b1a5fa0, 32'hbf1945a3} /* (24, 9, 3) {real, imag} */,
  {32'h39c09d00, 32'h3dd6d3b0} /* (24, 9, 2) {real, imag} */,
  {32'hbf94bd6a, 32'h3cafb200} /* (24, 9, 1) {real, imag} */,
  {32'h3cb079d0, 32'hbdfe9448} /* (24, 9, 0) {real, imag} */,
  {32'h3fbea0ad, 32'h3f37e9ca} /* (24, 8, 31) {real, imag} */,
  {32'hbf4f68e0, 32'hbe91f9a2} /* (24, 8, 30) {real, imag} */,
  {32'h3e0c7710, 32'h3df48fed} /* (24, 8, 29) {real, imag} */,
  {32'h3ec94199, 32'hbe325374} /* (24, 8, 28) {real, imag} */,
  {32'hbefcf1e8, 32'h3ec6e3bc} /* (24, 8, 27) {real, imag} */,
  {32'h3e940d74, 32'hbf15afd0} /* (24, 8, 26) {real, imag} */,
  {32'h3f13ccb2, 32'hbf423c84} /* (24, 8, 25) {real, imag} */,
  {32'hbde12076, 32'hbee6ae6b} /* (24, 8, 24) {real, imag} */,
  {32'h3c2a2c7c, 32'h3ebf9592} /* (24, 8, 23) {real, imag} */,
  {32'hbc943b35, 32'h3ee9c6b8} /* (24, 8, 22) {real, imag} */,
  {32'h3cea3504, 32'h3f00678e} /* (24, 8, 21) {real, imag} */,
  {32'h3e6d8fe1, 32'h3ec9a799} /* (24, 8, 20) {real, imag} */,
  {32'hbe16cfd5, 32'h3e16372a} /* (24, 8, 19) {real, imag} */,
  {32'h3d3dc57c, 32'h3cd27c88} /* (24, 8, 18) {real, imag} */,
  {32'h3da1087a, 32'h3d9e3d86} /* (24, 8, 17) {real, imag} */,
  {32'hbc301240, 32'hbea5a4be} /* (24, 8, 16) {real, imag} */,
  {32'h3e0fbca5, 32'h3e17b9b1} /* (24, 8, 15) {real, imag} */,
  {32'hbda20cf6, 32'h3e870902} /* (24, 8, 14) {real, imag} */,
  {32'h3e834d81, 32'hbd6d91fc} /* (24, 8, 13) {real, imag} */,
  {32'h3ea455d0, 32'hbe65f22e} /* (24, 8, 12) {real, imag} */,
  {32'h3dd3779f, 32'h3e39c296} /* (24, 8, 11) {real, imag} */,
  {32'hbdc4c118, 32'h3d96ab60} /* (24, 8, 10) {real, imag} */,
  {32'hbe1808df, 32'h3e762e16} /* (24, 8, 9) {real, imag} */,
  {32'hbebc57cc, 32'hbeb5a0d7} /* (24, 8, 8) {real, imag} */,
  {32'h3d415558, 32'hbed9cfe2} /* (24, 8, 7) {real, imag} */,
  {32'h3eef4b3e, 32'hbeff90bd} /* (24, 8, 6) {real, imag} */,
  {32'hbf1fe7d8, 32'hbe2c280d} /* (24, 8, 5) {real, imag} */,
  {32'h3f1a0965, 32'hbcd1fdf0} /* (24, 8, 4) {real, imag} */,
  {32'hbef48a33, 32'hbeb8e8c0} /* (24, 8, 3) {real, imag} */,
  {32'hbf75980a, 32'hbef83853} /* (24, 8, 2) {real, imag} */,
  {32'h3f92f4bd, 32'h3f1e7531} /* (24, 8, 1) {real, imag} */,
  {32'h3dbe2992, 32'h3ea422e0} /* (24, 8, 0) {real, imag} */,
  {32'hbf76203b, 32'h3c4a1e40} /* (24, 7, 31) {real, imag} */,
  {32'h3e026bdc, 32'h3e98e15e} /* (24, 7, 30) {real, imag} */,
  {32'hbea31d50, 32'h3e275ee3} /* (24, 7, 29) {real, imag} */,
  {32'hbf00d10b, 32'hbec4eefd} /* (24, 7, 28) {real, imag} */,
  {32'hbec289f5, 32'h3da42070} /* (24, 7, 27) {real, imag} */,
  {32'hbe6d6f4d, 32'hbf6afd46} /* (24, 7, 26) {real, imag} */,
  {32'h3e47b414, 32'h3edec1aa} /* (24, 7, 25) {real, imag} */,
  {32'h3ea68770, 32'h3eab7aa4} /* (24, 7, 24) {real, imag} */,
  {32'h3f2675bf, 32'h3eb15da0} /* (24, 7, 23) {real, imag} */,
  {32'hbd8f8e96, 32'hbdf1a820} /* (24, 7, 22) {real, imag} */,
  {32'hbf131e78, 32'hbdb83abc} /* (24, 7, 21) {real, imag} */,
  {32'h3d90c83f, 32'h3ede7e2c} /* (24, 7, 20) {real, imag} */,
  {32'hbe654f6c, 32'h3e339b78} /* (24, 7, 19) {real, imag} */,
  {32'hbeff155e, 32'h3d2da0f4} /* (24, 7, 18) {real, imag} */,
  {32'h3e97384d, 32'hbe673fb3} /* (24, 7, 17) {real, imag} */,
  {32'hbe1015ad, 32'hbe3c8549} /* (24, 7, 16) {real, imag} */,
  {32'hbe2d6530, 32'h3e772870} /* (24, 7, 15) {real, imag} */,
  {32'h3f11d8fa, 32'h3ecaea74} /* (24, 7, 14) {real, imag} */,
  {32'h3ed4befa, 32'hbd55d662} /* (24, 7, 13) {real, imag} */,
  {32'h3eba12ba, 32'h3e9800a2} /* (24, 7, 12) {real, imag} */,
  {32'hbe0d0b2b, 32'h3dda5912} /* (24, 7, 11) {real, imag} */,
  {32'hbeb6deb8, 32'h3f331fa9} /* (24, 7, 10) {real, imag} */,
  {32'h3f010876, 32'hbd7a1908} /* (24, 7, 9) {real, imag} */,
  {32'h3e7c305a, 32'h3f826b74} /* (24, 7, 8) {real, imag} */,
  {32'hbe6b2600, 32'hbecde22a} /* (24, 7, 7) {real, imag} */,
  {32'h3cba2f40, 32'hbe075817} /* (24, 7, 6) {real, imag} */,
  {32'hbe95c452, 32'h3ed4f8c1} /* (24, 7, 5) {real, imag} */,
  {32'h3e84a084, 32'hbd5c8cab} /* (24, 7, 4) {real, imag} */,
  {32'hbf0363fa, 32'h3f304c2c} /* (24, 7, 3) {real, imag} */,
  {32'hbc7c3f30, 32'h3f83b6c0} /* (24, 7, 2) {real, imag} */,
  {32'hbf4e74de, 32'hbf7477c7} /* (24, 7, 1) {real, imag} */,
  {32'hbf182442, 32'hbea70262} /* (24, 7, 0) {real, imag} */,
  {32'h3ea7404c, 32'hbe1de668} /* (24, 6, 31) {real, imag} */,
  {32'hbe628d1e, 32'h3ef450aa} /* (24, 6, 30) {real, imag} */,
  {32'hbe828e68, 32'hbec39cf5} /* (24, 6, 29) {real, imag} */,
  {32'h3f21d446, 32'h3f29c722} /* (24, 6, 28) {real, imag} */,
  {32'hbd11848c, 32'hbcb3a7c0} /* (24, 6, 27) {real, imag} */,
  {32'hbf65bf77, 32'h3ee318a0} /* (24, 6, 26) {real, imag} */,
  {32'hbdaaef31, 32'h3f10c9a1} /* (24, 6, 25) {real, imag} */,
  {32'hbcb72104, 32'hbf394bda} /* (24, 6, 24) {real, imag} */,
  {32'hbed46a88, 32'h3c0d88c0} /* (24, 6, 23) {real, imag} */,
  {32'hbea0375e, 32'hbe4233b3} /* (24, 6, 22) {real, imag} */,
  {32'hbec15463, 32'h3e5d6df0} /* (24, 6, 21) {real, imag} */,
  {32'h3ee9c9fc, 32'hbd0576c0} /* (24, 6, 20) {real, imag} */,
  {32'h3f310193, 32'hbe764879} /* (24, 6, 19) {real, imag} */,
  {32'h3d4f319c, 32'hbe8f6c61} /* (24, 6, 18) {real, imag} */,
  {32'h3b5aefb0, 32'h3ea713a1} /* (24, 6, 17) {real, imag} */,
  {32'hbbe9df00, 32'hbd471596} /* (24, 6, 16) {real, imag} */,
  {32'h3e05609e, 32'hbdf81e8c} /* (24, 6, 15) {real, imag} */,
  {32'h3e988a54, 32'h3e44a596} /* (24, 6, 14) {real, imag} */,
  {32'hbe8f0e0a, 32'hbd89e157} /* (24, 6, 13) {real, imag} */,
  {32'hbdf60737, 32'hbf14597c} /* (24, 6, 12) {real, imag} */,
  {32'hbf346da8, 32'h3c06fa20} /* (24, 6, 11) {real, imag} */,
  {32'hbec9e764, 32'h3e8ac272} /* (24, 6, 10) {real, imag} */,
  {32'h3f3fcafa, 32'hbea2c0ca} /* (24, 6, 9) {real, imag} */,
  {32'hbe86aba6, 32'hbe953478} /* (24, 6, 8) {real, imag} */,
  {32'hbeb7e425, 32'h3e613e98} /* (24, 6, 7) {real, imag} */,
  {32'h3afd6880, 32'hbf533a36} /* (24, 6, 6) {real, imag} */,
  {32'h3f370c02, 32'h3d6556f8} /* (24, 6, 5) {real, imag} */,
  {32'h3ecc1193, 32'h3eb7ad74} /* (24, 6, 4) {real, imag} */,
  {32'h3d15d6bc, 32'h3de17376} /* (24, 6, 3) {real, imag} */,
  {32'h3f90c538, 32'hbddc70aa} /* (24, 6, 2) {real, imag} */,
  {32'hbe911978, 32'hbe09fe5b} /* (24, 6, 1) {real, imag} */,
  {32'hbd94d688, 32'hbe0ee3cc} /* (24, 6, 0) {real, imag} */,
  {32'h406763bc, 32'h3ef0a48d} /* (24, 5, 31) {real, imag} */,
  {32'hbfe2499d, 32'h3ce20c40} /* (24, 5, 30) {real, imag} */,
  {32'h3e7c0ebd, 32'hbf0639f2} /* (24, 5, 29) {real, imag} */,
  {32'h3e37cb82, 32'h3dbeeb96} /* (24, 5, 28) {real, imag} */,
  {32'hbf7cc1ae, 32'h3f35833a} /* (24, 5, 27) {real, imag} */,
  {32'h3f248003, 32'h3d45ef68} /* (24, 5, 26) {real, imag} */,
  {32'hbec06f0a, 32'hbebcb7fe} /* (24, 5, 25) {real, imag} */,
  {32'hbe403cbc, 32'hbe94f407} /* (24, 5, 24) {real, imag} */,
  {32'h3d7d82fa, 32'h3cf80d18} /* (24, 5, 23) {real, imag} */,
  {32'hbe80da3d, 32'h3ea23213} /* (24, 5, 22) {real, imag} */,
  {32'hbe5a5e72, 32'hbc8fa0a0} /* (24, 5, 21) {real, imag} */,
  {32'hbdc875de, 32'h3d629874} /* (24, 5, 20) {real, imag} */,
  {32'h3e81c6c8, 32'hbe9be939} /* (24, 5, 19) {real, imag} */,
  {32'hbe425a2a, 32'h3e029510} /* (24, 5, 18) {real, imag} */,
  {32'hbe2de89a, 32'h3c9ff5e6} /* (24, 5, 17) {real, imag} */,
  {32'h3e5ccb34, 32'h3dd0c612} /* (24, 5, 16) {real, imag} */,
  {32'hbe93444c, 32'hbdf26188} /* (24, 5, 15) {real, imag} */,
  {32'hbe3c3010, 32'hbed183d1} /* (24, 5, 14) {real, imag} */,
  {32'hbefb5636, 32'hbeb8926b} /* (24, 5, 13) {real, imag} */,
  {32'h3e5be933, 32'hbd42e406} /* (24, 5, 12) {real, imag} */,
  {32'h3dbc3e9b, 32'h3de423d4} /* (24, 5, 11) {real, imag} */,
  {32'h3e8477ec, 32'hbe4158ee} /* (24, 5, 10) {real, imag} */,
  {32'hbf0812e2, 32'h3e41b86e} /* (24, 5, 9) {real, imag} */,
  {32'h3da801d8, 32'hbf049e9a} /* (24, 5, 8) {real, imag} */,
  {32'h3ec1b58c, 32'h3e756444} /* (24, 5, 7) {real, imag} */,
  {32'hbebfe688, 32'hbbd9b380} /* (24, 5, 6) {real, imag} */,
  {32'h3d67c470, 32'hbf0a69a6} /* (24, 5, 5) {real, imag} */,
  {32'h3dd0ba0c, 32'h3f8157cc} /* (24, 5, 4) {real, imag} */,
  {32'h3ee4cd44, 32'hbe9e4582} /* (24, 5, 3) {real, imag} */,
  {32'hbf85c5e0, 32'hbfb14f54} /* (24, 5, 2) {real, imag} */,
  {32'h3fd43057, 32'h4027e872} /* (24, 5, 1) {real, imag} */,
  {32'h3fc1438a, 32'h3f76d6c1} /* (24, 5, 0) {real, imag} */,
  {32'hbfaf51f3, 32'hc03b7c9e} /* (24, 4, 31) {real, imag} */,
  {32'h4012366f, 32'h40499c03} /* (24, 4, 30) {real, imag} */,
  {32'h3d181108, 32'hbf6a39f2} /* (24, 4, 29) {real, imag} */,
  {32'hbfe3deca, 32'hbf923c7d} /* (24, 4, 28) {real, imag} */,
  {32'h3ec795a8, 32'hbeef6cb8} /* (24, 4, 27) {real, imag} */,
  {32'h3f2dbcfe, 32'hbf1a5c43} /* (24, 4, 26) {real, imag} */,
  {32'hbd718830, 32'h3dba8748} /* (24, 4, 25) {real, imag} */,
  {32'h3f0adde4, 32'h3ec2ceab} /* (24, 4, 24) {real, imag} */,
  {32'h3f2c2990, 32'hbee13998} /* (24, 4, 23) {real, imag} */,
  {32'hbf085499, 32'h3e5b455c} /* (24, 4, 22) {real, imag} */,
  {32'h3eaf6748, 32'h3e377b8e} /* (24, 4, 21) {real, imag} */,
  {32'hbd67ece0, 32'hbd6e9530} /* (24, 4, 20) {real, imag} */,
  {32'hbe260275, 32'hbe7022ee} /* (24, 4, 19) {real, imag} */,
  {32'h3e272405, 32'hbe3c16ea} /* (24, 4, 18) {real, imag} */,
  {32'h3e6572e8, 32'h3ee99fd0} /* (24, 4, 17) {real, imag} */,
  {32'hbe5567d2, 32'h3dbc08e7} /* (24, 4, 16) {real, imag} */,
  {32'hbb4d8680, 32'hbe76ca73} /* (24, 4, 15) {real, imag} */,
  {32'h3e0160ae, 32'h3e926220} /* (24, 4, 14) {real, imag} */,
  {32'h3e46e964, 32'hbea15006} /* (24, 4, 13) {real, imag} */,
  {32'hbe9711e0, 32'hbe96043e} /* (24, 4, 12) {real, imag} */,
  {32'hbda9feda, 32'h3f0213d6} /* (24, 4, 11) {real, imag} */,
  {32'h3eb8bd7f, 32'hbf008031} /* (24, 4, 10) {real, imag} */,
  {32'h3ef24d46, 32'h3e3ee805} /* (24, 4, 9) {real, imag} */,
  {32'hbe1c8886, 32'h3ed58dee} /* (24, 4, 8) {real, imag} */,
  {32'hbf291dd4, 32'h3e5561fc} /* (24, 4, 7) {real, imag} */,
  {32'hbf512acd, 32'h3ddb0574} /* (24, 4, 6) {real, imag} */,
  {32'hbe9622e1, 32'h3f2dfb16} /* (24, 4, 5) {real, imag} */,
  {32'h3f59b7e6, 32'hbfdd0dee} /* (24, 4, 4) {real, imag} */,
  {32'h3f2cbf7c, 32'hbec4c790} /* (24, 4, 3) {real, imag} */,
  {32'h40769f0c, 32'h3fce413e} /* (24, 4, 2) {real, imag} */,
  {32'hc08f7771, 32'hbf8d80e7} /* (24, 4, 1) {real, imag} */,
  {32'hc0170c33, 32'hbf7776a4} /* (24, 4, 0) {real, imag} */,
  {32'h406e42f4, 32'hc03b5b5c} /* (24, 3, 31) {real, imag} */,
  {32'hc00909d8, 32'h402a7b68} /* (24, 3, 30) {real, imag} */,
  {32'h3eae0e67, 32'h3f6e17d9} /* (24, 3, 29) {real, imag} */,
  {32'hbf30c5a2, 32'hbf7cc259} /* (24, 3, 28) {real, imag} */,
  {32'h3f99523e, 32'h3e89de0d} /* (24, 3, 27) {real, imag} */,
  {32'hbe324cc2, 32'h3ea762ec} /* (24, 3, 26) {real, imag} */,
  {32'hbe30bddc, 32'hbede12ca} /* (24, 3, 25) {real, imag} */,
  {32'hbe9ddd94, 32'h3f2bcb94} /* (24, 3, 24) {real, imag} */,
  {32'hbf1c1dc0, 32'h3e197d6d} /* (24, 3, 23) {real, imag} */,
  {32'h3e507c55, 32'h3e8b42fe} /* (24, 3, 22) {real, imag} */,
  {32'hbe0808b6, 32'hbf0ab045} /* (24, 3, 21) {real, imag} */,
  {32'h3d688362, 32'h3e4514c1} /* (24, 3, 20) {real, imag} */,
  {32'hbd8d48ac, 32'hbf181ee6} /* (24, 3, 19) {real, imag} */,
  {32'h3e99eda7, 32'h3f370f59} /* (24, 3, 18) {real, imag} */,
  {32'hbdbd6eac, 32'h3d9c51d3} /* (24, 3, 17) {real, imag} */,
  {32'h3e4e5534, 32'hbdd980f4} /* (24, 3, 16) {real, imag} */,
  {32'h3d21a4e8, 32'hbd4732c0} /* (24, 3, 15) {real, imag} */,
  {32'hbc0f6978, 32'h3d91da00} /* (24, 3, 14) {real, imag} */,
  {32'hbf47c258, 32'hbdf57863} /* (24, 3, 13) {real, imag} */,
  {32'hbd6feac8, 32'hbd297c70} /* (24, 3, 12) {real, imag} */,
  {32'h3e7486fe, 32'h3cb0a94c} /* (24, 3, 11) {real, imag} */,
  {32'h3e3fb824, 32'hbc1e5a58} /* (24, 3, 10) {real, imag} */,
  {32'h3ea37a9c, 32'hbdb111da} /* (24, 3, 9) {real, imag} */,
  {32'h3dce781c, 32'h3dff605e} /* (24, 3, 8) {real, imag} */,
  {32'hbec0b7c2, 32'hbcea4a60} /* (24, 3, 7) {real, imag} */,
  {32'hbef947b9, 32'h3f7b27a8} /* (24, 3, 6) {real, imag} */,
  {32'hbe74c42d, 32'hbf174d74} /* (24, 3, 5) {real, imag} */,
  {32'h3fb53f41, 32'hbf1c749e} /* (24, 3, 4) {real, imag} */,
  {32'h3be41d40, 32'hbdf2ac48} /* (24, 3, 3) {real, imag} */,
  {32'hbf3d8f3c, 32'h407b3b78} /* (24, 3, 2) {real, imag} */,
  {32'hc06a3ab7, 32'hc02e5ab6} /* (24, 3, 1) {real, imag} */,
  {32'h403aac1c, 32'h3eb32833} /* (24, 3, 0) {real, imag} */,
  {32'h41e1eb34, 32'h3fe216af} /* (24, 2, 31) {real, imag} */,
  {32'hc15475c7, 32'h40491990} /* (24, 2, 30) {real, imag} */,
  {32'h3fb71b66, 32'hbf604c0a} /* (24, 2, 29) {real, imag} */,
  {32'h3fcc8c7c, 32'hbfc4b9aa} /* (24, 2, 28) {real, imag} */,
  {32'hbf7e4eb0, 32'h3ea7d3d1} /* (24, 2, 27) {real, imag} */,
  {32'hbf41d6bc, 32'h3ea976a5} /* (24, 2, 26) {real, imag} */,
  {32'hbeaa64c7, 32'h3ea798e2} /* (24, 2, 25) {real, imag} */,
  {32'h3c4d80c0, 32'h3f9581f2} /* (24, 2, 24) {real, imag} */,
  {32'h3f0916ba, 32'h3db6bbbe} /* (24, 2, 23) {real, imag} */,
  {32'hbe9f356f, 32'hbee11de0} /* (24, 2, 22) {real, imag} */,
  {32'h3f6617f8, 32'h3ed8d9fe} /* (24, 2, 21) {real, imag} */,
  {32'hbd8870b4, 32'hbef43f38} /* (24, 2, 20) {real, imag} */,
  {32'hbe367834, 32'h3ea4fbdf} /* (24, 2, 19) {real, imag} */,
  {32'h3d681c4a, 32'h3e61a8ff} /* (24, 2, 18) {real, imag} */,
  {32'hbe3c473e, 32'h3cbf3598} /* (24, 2, 17) {real, imag} */,
  {32'hbe32c55c, 32'h3dfb3631} /* (24, 2, 16) {real, imag} */,
  {32'h3dc35ade, 32'hbe450d37} /* (24, 2, 15) {real, imag} */,
  {32'hbd376e04, 32'hbe1ec6f6} /* (24, 2, 14) {real, imag} */,
  {32'hbe129db8, 32'hbeecd54e} /* (24, 2, 13) {real, imag} */,
  {32'h3e9e9f07, 32'h3ebeb63c} /* (24, 2, 12) {real, imag} */,
  {32'hbe86951e, 32'hbf0a8943} /* (24, 2, 11) {real, imag} */,
  {32'h3ea1e90f, 32'hbf0abe24} /* (24, 2, 10) {real, imag} */,
  {32'h3e79165d, 32'h3c51be70} /* (24, 2, 9) {real, imag} */,
  {32'hbf0d9b6e, 32'h3e51e0cf} /* (24, 2, 8) {real, imag} */,
  {32'h3ef633d0, 32'h3e60b594} /* (24, 2, 7) {real, imag} */,
  {32'h3f485b5a, 32'h3b0a57c0} /* (24, 2, 6) {real, imag} */,
  {32'hc01e93f2, 32'hbf9c20fb} /* (24, 2, 5) {real, imag} */,
  {32'h40349c5c, 32'h3f28ef62} /* (24, 2, 4) {real, imag} */,
  {32'h3e8689ce, 32'hbfa4e195} /* (24, 2, 3) {real, imag} */,
  {32'hc104b84e, 32'h3fa1f5cc} /* (24, 2, 2) {real, imag} */,
  {32'h4183bf18, 32'hbf8b6cb7} /* (24, 2, 1) {real, imag} */,
  {32'h4170ba5e, 32'h40121bb6} /* (24, 2, 0) {real, imag} */,
  {32'hc2177b8b, 32'h4117591a} /* (24, 1, 31) {real, imag} */,
  {32'h410a21ab, 32'h40355130} /* (24, 1, 30) {real, imag} */,
  {32'h3fbcef3e, 32'hbf5067d0} /* (24, 1, 29) {real, imag} */,
  {32'hc031d835, 32'hbf0f146e} /* (24, 1, 28) {real, imag} */,
  {32'h403d1066, 32'hbe9dc783} /* (24, 1, 27) {real, imag} */,
  {32'hbf64ff74, 32'hbe5e3bb6} /* (24, 1, 26) {real, imag} */,
  {32'hbf2995b9, 32'h3f171191} /* (24, 1, 25) {real, imag} */,
  {32'h3f6df247, 32'hbf756b36} /* (24, 1, 24) {real, imag} */,
  {32'h3edfb864, 32'h3e1fab2d} /* (24, 1, 23) {real, imag} */,
  {32'h3e2d67a2, 32'hbf221b46} /* (24, 1, 22) {real, imag} */,
  {32'h3e9b3418, 32'hbf4e1184} /* (24, 1, 21) {real, imag} */,
  {32'hbf23941a, 32'h3e8842c2} /* (24, 1, 20) {real, imag} */,
  {32'h3e17426a, 32'hbf11c677} /* (24, 1, 19) {real, imag} */,
  {32'hbd587bf8, 32'hbf0aa1f2} /* (24, 1, 18) {real, imag} */,
  {32'h3d9bd268, 32'h3e5fb4ea} /* (24, 1, 17) {real, imag} */,
  {32'h3cc46fc8, 32'hbdc209b4} /* (24, 1, 16) {real, imag} */,
  {32'hbc3d1c00, 32'hbddc9e08} /* (24, 1, 15) {real, imag} */,
  {32'hbe69c1a8, 32'h3efd4c14} /* (24, 1, 14) {real, imag} */,
  {32'hbb3b4ba0, 32'hbecefacc} /* (24, 1, 13) {real, imag} */,
  {32'hbddc2fc6, 32'hbcb40ca0} /* (24, 1, 12) {real, imag} */,
  {32'h3e4c3c0d, 32'h3f011cc6} /* (24, 1, 11) {real, imag} */,
  {32'hbe57a006, 32'hbe76db3a} /* (24, 1, 10) {real, imag} */,
  {32'hbaf3f480, 32'h3e7dbbe6} /* (24, 1, 9) {real, imag} */,
  {32'h3f497c17, 32'h3f59d703} /* (24, 1, 8) {real, imag} */,
  {32'hbec65812, 32'hbeeb890a} /* (24, 1, 7) {real, imag} */,
  {32'h3efa6cdc, 32'hbd201aa8} /* (24, 1, 6) {real, imag} */,
  {32'h4006aabc, 32'h3fbd260a} /* (24, 1, 5) {real, imag} */,
  {32'hbf48c5bc, 32'hbfc0efb0} /* (24, 1, 4) {real, imag} */,
  {32'h3f2cdc58, 32'h3ef6266a} /* (24, 1, 3) {real, imag} */,
  {32'h4153f596, 32'h414c952c} /* (24, 1, 2) {real, imag} */,
  {32'hc25a1b49, 32'hc1fba9e1} /* (24, 1, 1) {real, imag} */,
  {32'hc24ea4af, 32'hc0dbd352} /* (24, 1, 0) {real, imag} */,
  {32'hc218aeef, 32'h41eece01} /* (24, 0, 31) {real, imag} */,
  {32'h40836024, 32'hc09e667a} /* (24, 0, 30) {real, imag} */,
  {32'h3f82c1d0, 32'h3f2e93e5} /* (24, 0, 29) {real, imag} */,
  {32'h3f8c1c00, 32'hc02fa9ed} /* (24, 0, 28) {real, imag} */,
  {32'h3fda5078, 32'hbf18fd08} /* (24, 0, 27) {real, imag} */,
  {32'h3f2f62fa, 32'h3db15f7c} /* (24, 0, 26) {real, imag} */,
  {32'h3f398a10, 32'h3e582484} /* (24, 0, 25) {real, imag} */,
  {32'h3e377c1e, 32'hbea07ca8} /* (24, 0, 24) {real, imag} */,
  {32'hbf325277, 32'hbea78586} /* (24, 0, 23) {real, imag} */,
  {32'hbdfa43db, 32'hbe7d8f1c} /* (24, 0, 22) {real, imag} */,
  {32'hbc81da88, 32'hbc1a1e60} /* (24, 0, 21) {real, imag} */,
  {32'hbf144378, 32'hbdb78edc} /* (24, 0, 20) {real, imag} */,
  {32'hbdb1880c, 32'h3d1b49fb} /* (24, 0, 19) {real, imag} */,
  {32'h3ef74a8e, 32'hbd6a3550} /* (24, 0, 18) {real, imag} */,
  {32'hbdc83e7f, 32'h3cf20684} /* (24, 0, 17) {real, imag} */,
  {32'h3ede1625, 32'h00000000} /* (24, 0, 16) {real, imag} */,
  {32'hbdc83e7f, 32'hbcf20684} /* (24, 0, 15) {real, imag} */,
  {32'h3ef74a8e, 32'h3d6a3550} /* (24, 0, 14) {real, imag} */,
  {32'hbdb1880c, 32'hbd1b49fb} /* (24, 0, 13) {real, imag} */,
  {32'hbf144378, 32'h3db78edc} /* (24, 0, 12) {real, imag} */,
  {32'hbc81da88, 32'h3c1a1e60} /* (24, 0, 11) {real, imag} */,
  {32'hbdfa43db, 32'h3e7d8f1c} /* (24, 0, 10) {real, imag} */,
  {32'hbf325277, 32'h3ea78586} /* (24, 0, 9) {real, imag} */,
  {32'h3e377c1e, 32'h3ea07ca8} /* (24, 0, 8) {real, imag} */,
  {32'h3f398a10, 32'hbe582484} /* (24, 0, 7) {real, imag} */,
  {32'h3f2f62fa, 32'hbdb15f7c} /* (24, 0, 6) {real, imag} */,
  {32'h3fda5078, 32'h3f18fd08} /* (24, 0, 5) {real, imag} */,
  {32'h3f8c1c00, 32'h402fa9ed} /* (24, 0, 4) {real, imag} */,
  {32'h3f82c1d0, 32'hbf2e93e5} /* (24, 0, 3) {real, imag} */,
  {32'h40836024, 32'h409e667a} /* (24, 0, 2) {real, imag} */,
  {32'hc218aeef, 32'hc1eece01} /* (24, 0, 1) {real, imag} */,
  {32'hc2708769, 32'h00000000} /* (24, 0, 0) {real, imag} */,
  {32'hc2868bfc, 32'h4217fdc2} /* (23, 31, 31) {real, imag} */,
  {32'h4183b620, 32'hc174792e} /* (23, 31, 30) {real, imag} */,
  {32'h3fe795ba, 32'hbf117c12} /* (23, 31, 29) {real, imag} */,
  {32'hbff79290, 32'h3fce75d0} /* (23, 31, 28) {real, imag} */,
  {32'h4009667e, 32'hbfbc3ea8} /* (23, 31, 27) {real, imag} */,
  {32'h3f7a9161, 32'h3f1f313e} /* (23, 31, 26) {real, imag} */,
  {32'hbf1b6a79, 32'h3ef13484} /* (23, 31, 25) {real, imag} */,
  {32'h3f08e354, 32'hbf047db0} /* (23, 31, 24) {real, imag} */,
  {32'h3f22d8b8, 32'hbe560520} /* (23, 31, 23) {real, imag} */,
  {32'h3e8a7593, 32'h3da5abe0} /* (23, 31, 22) {real, imag} */,
  {32'hbe157f2a, 32'hbf49ef1c} /* (23, 31, 21) {real, imag} */,
  {32'h3d9276c0, 32'h3d8b597a} /* (23, 31, 20) {real, imag} */,
  {32'h3d412f58, 32'h3e9cd642} /* (23, 31, 19) {real, imag} */,
  {32'hbb7af530, 32'hbe711340} /* (23, 31, 18) {real, imag} */,
  {32'h3e157fdf, 32'h3dc5ed62} /* (23, 31, 17) {real, imag} */,
  {32'hbcc096e4, 32'hbd37c518} /* (23, 31, 16) {real, imag} */,
  {32'h3da61db8, 32'h3ecb530e} /* (23, 31, 15) {real, imag} */,
  {32'hbe95d8c3, 32'h3e81f154} /* (23, 31, 14) {real, imag} */,
  {32'h3cc31cb4, 32'hbe2416b5} /* (23, 31, 13) {real, imag} */,
  {32'hbdb680a9, 32'hbd271c0e} /* (23, 31, 12) {real, imag} */,
  {32'h3ed4f591, 32'h3e626385} /* (23, 31, 11) {real, imag} */,
  {32'hbeb5a73e, 32'h3bf46030} /* (23, 31, 10) {real, imag} */,
  {32'h3e8b3e58, 32'h3f02ef78} /* (23, 31, 9) {real, imag} */,
  {32'h3ee4f898, 32'h3f18423e} /* (23, 31, 8) {real, imag} */,
  {32'hbf08bbaa, 32'hbf32af03} /* (23, 31, 7) {real, imag} */,
  {32'h3f000e6c, 32'hbe0ba27f} /* (23, 31, 6) {real, imag} */,
  {32'h40835292, 32'h3e8a4b87} /* (23, 31, 5) {real, imag} */,
  {32'hc07497c3, 32'h3f3b464a} /* (23, 31, 4) {real, imag} */,
  {32'h3fbed4c7, 32'h3f917ce6} /* (23, 31, 3) {real, imag} */,
  {32'h41397e08, 32'hc047a4af} /* (23, 31, 2) {real, imag} */,
  {32'hc23ef642, 32'hc1464375} /* (23, 31, 1) {real, imag} */,
  {32'hc277c643, 32'h40f49fae} /* (23, 31, 0) {real, imag} */,
  {32'h41a3b111, 32'h400030bb} /* (23, 30, 31) {real, imag} */,
  {32'hc13782d9, 32'hbfe039dd} /* (23, 30, 30) {real, imag} */,
  {32'h3e3051ae, 32'h3f84bbfa} /* (23, 30, 29) {real, imag} */,
  {32'h403ae243, 32'hbfef8566} /* (23, 30, 28) {real, imag} */,
  {32'hc01969ca, 32'h40095e65} /* (23, 30, 27) {real, imag} */,
  {32'hbd5b9b90, 32'hbe14fb42} /* (23, 30, 26) {real, imag} */,
  {32'h3f12a0e2, 32'hbe98f4de} /* (23, 30, 25) {real, imag} */,
  {32'hbf47eb87, 32'hbf40f53e} /* (23, 30, 24) {real, imag} */,
  {32'h3eb4e1ee, 32'hbec9d1cb} /* (23, 30, 23) {real, imag} */,
  {32'h3df705b6, 32'hbebf5da4} /* (23, 30, 22) {real, imag} */,
  {32'hbea8cdde, 32'h3ee9f938} /* (23, 30, 21) {real, imag} */,
  {32'hbe101495, 32'hbe03563e} /* (23, 30, 20) {real, imag} */,
  {32'hbe0d3392, 32'h3cc36538} /* (23, 30, 19) {real, imag} */,
  {32'hbe5dafee, 32'h3d7c2230} /* (23, 30, 18) {real, imag} */,
  {32'h3ecd39ba, 32'hbe840d6c} /* (23, 30, 17) {real, imag} */,
  {32'hbe8054e7, 32'hbeccd86c} /* (23, 30, 16) {real, imag} */,
  {32'hbe96f083, 32'h3eca5172} /* (23, 30, 15) {real, imag} */,
  {32'h3cf7215d, 32'hbcc684e0} /* (23, 30, 14) {real, imag} */,
  {32'h3e681410, 32'hbe8996f8} /* (23, 30, 13) {real, imag} */,
  {32'h3e349ca0, 32'hbe835139} /* (23, 30, 12) {real, imag} */,
  {32'hbda19e03, 32'h3c9d9d76} /* (23, 30, 11) {real, imag} */,
  {32'h3dca5c8e, 32'hbe8e57a6} /* (23, 30, 10) {real, imag} */,
  {32'hbe92a177, 32'hbe6a2e14} /* (23, 30, 9) {real, imag} */,
  {32'hbe0e63de, 32'hbf075939} /* (23, 30, 8) {real, imag} */,
  {32'h3e1d8022, 32'hbe49aef5} /* (23, 30, 7) {real, imag} */,
  {32'hbecdc896, 32'hbf2648f5} /* (23, 30, 6) {real, imag} */,
  {32'hbfef603e, 32'hbef0b745} /* (23, 30, 5) {real, imag} */,
  {32'h3f90b104, 32'h4026d48d} /* (23, 30, 4) {real, imag} */,
  {32'h3f85622a, 32'h3f7e6136} /* (23, 30, 3) {real, imag} */,
  {32'hc1804dd6, 32'hc098de2e} /* (23, 30, 2) {real, imag} */,
  {32'h420d8d54, 32'hc00929ed} /* (23, 30, 1) {real, imag} */,
  {32'h41936f1d, 32'hc05ebdb6} /* (23, 30, 0) {real, imag} */,
  {32'hc07a0378, 32'h400b5b6e} /* (23, 29, 31) {real, imag} */,
  {32'hbf0fba7a, 32'hc094b7e2} /* (23, 29, 30) {real, imag} */,
  {32'hbe898167, 32'h3e72d87c} /* (23, 29, 29) {real, imag} */,
  {32'h3f99a45a, 32'h3f971346} /* (23, 29, 28) {real, imag} */,
  {32'hbeff5bf6, 32'h3f18e7ab} /* (23, 29, 27) {real, imag} */,
  {32'hbec75569, 32'hbf2ba4e3} /* (23, 29, 26) {real, imag} */,
  {32'hbeb5a23a, 32'h3f2fadc0} /* (23, 29, 25) {real, imag} */,
  {32'hbe860738, 32'hbee1a9de} /* (23, 29, 24) {real, imag} */,
  {32'h3d847a64, 32'hbc170c38} /* (23, 29, 23) {real, imag} */,
  {32'hbe328a51, 32'hbe6fe7f5} /* (23, 29, 22) {real, imag} */,
  {32'h3e9452f5, 32'h3e5fc04f} /* (23, 29, 21) {real, imag} */,
  {32'hbf060867, 32'h3efbb03a} /* (23, 29, 20) {real, imag} */,
  {32'h3dbbc1ae, 32'hbd89c567} /* (23, 29, 19) {real, imag} */,
  {32'h3ceab118, 32'hbea1dce6} /* (23, 29, 18) {real, imag} */,
  {32'h3e11f61f, 32'h3ddaf65c} /* (23, 29, 17) {real, imag} */,
  {32'h3f09be82, 32'hbd0e9e6c} /* (23, 29, 16) {real, imag} */,
  {32'hbe9b4e51, 32'hbdf626b0} /* (23, 29, 15) {real, imag} */,
  {32'h3e661327, 32'hbe42aa06} /* (23, 29, 14) {real, imag} */,
  {32'hbe75e146, 32'hbeaf8656} /* (23, 29, 13) {real, imag} */,
  {32'hbe8803fc, 32'h3ed798a4} /* (23, 29, 12) {real, imag} */,
  {32'h3d734252, 32'h3e5d369b} /* (23, 29, 11) {real, imag} */,
  {32'hbdc4a30c, 32'h3d8b2673} /* (23, 29, 10) {real, imag} */,
  {32'hbeba70ab, 32'h3ee9f307} /* (23, 29, 9) {real, imag} */,
  {32'hbe7842c4, 32'hbed18260} /* (23, 29, 8) {real, imag} */,
  {32'hbc51c5c0, 32'h3f7302c2} /* (23, 29, 7) {real, imag} */,
  {32'hbea10dfb, 32'hbe3854ed} /* (23, 29, 6) {real, imag} */,
  {32'h3fbe318e, 32'hbdc4c28c} /* (23, 29, 5) {real, imag} */,
  {32'hbf9632bb, 32'h3f538c60} /* (23, 29, 4) {real, imag} */,
  {32'hbeeb201a, 32'hbea2248a} /* (23, 29, 3) {real, imag} */,
  {32'hc004e30c, 32'hc04ca452} /* (23, 29, 2) {real, imag} */,
  {32'h4087fc76, 32'h402ade2e} /* (23, 29, 1) {real, imag} */,
  {32'h403289dc, 32'hbe8fab8d} /* (23, 29, 0) {real, imag} */,
  {32'hc084c3d7, 32'h3fef1274} /* (23, 28, 31) {real, imag} */,
  {32'h406c2057, 32'hbfe18a3b} /* (23, 28, 30) {real, imag} */,
  {32'h3ef02ed0, 32'h3f449130} /* (23, 28, 29) {real, imag} */,
  {32'h3f86d6d6, 32'h3fa65bf0} /* (23, 28, 28) {real, imag} */,
  {32'h3e8a241c, 32'hbda70af4} /* (23, 28, 27) {real, imag} */,
  {32'hbf1cb234, 32'hbe24a876} /* (23, 28, 26) {real, imag} */,
  {32'hbf439506, 32'h3e849418} /* (23, 28, 25) {real, imag} */,
  {32'h3e0b4bbe, 32'h3ecc0111} /* (23, 28, 24) {real, imag} */,
  {32'hbe6f21ae, 32'h3eaf7851} /* (23, 28, 23) {real, imag} */,
  {32'h3e7dbe28, 32'hbe8a49f0} /* (23, 28, 22) {real, imag} */,
  {32'hbee21ae0, 32'hbec690a3} /* (23, 28, 21) {real, imag} */,
  {32'hbdef15c8, 32'hbd14386c} /* (23, 28, 20) {real, imag} */,
  {32'hbdb3f2ec, 32'hbe72c11e} /* (23, 28, 19) {real, imag} */,
  {32'h3c1399c8, 32'hbedb53d6} /* (23, 28, 18) {real, imag} */,
  {32'h3eafde39, 32'h3e2dc509} /* (23, 28, 17) {real, imag} */,
  {32'hbd97fd9a, 32'hbdd39c0b} /* (23, 28, 16) {real, imag} */,
  {32'h3ca57258, 32'h3eb4ff53} /* (23, 28, 15) {real, imag} */,
  {32'h3d56d6cc, 32'hbe95c101} /* (23, 28, 14) {real, imag} */,
  {32'h3ee15fd6, 32'h3e4b687f} /* (23, 28, 13) {real, imag} */,
  {32'h3e8448f0, 32'hbed5fba0} /* (23, 28, 12) {real, imag} */,
  {32'h3c442a58, 32'h3e8d2907} /* (23, 28, 11) {real, imag} */,
  {32'hbef1ffd4, 32'hbe827f1a} /* (23, 28, 10) {real, imag} */,
  {32'hbdb9c4ba, 32'h3bd00048} /* (23, 28, 9) {real, imag} */,
  {32'h3fca805e, 32'hbe0fce1c} /* (23, 28, 8) {real, imag} */,
  {32'hbece9410, 32'h3d8da686} /* (23, 28, 7) {real, imag} */,
  {32'hbe142418, 32'h3e2e4926} /* (23, 28, 6) {real, imag} */,
  {32'h3f512176, 32'h3f54c085} /* (23, 28, 5) {real, imag} */,
  {32'hbfc33705, 32'h3ef77f69} /* (23, 28, 4) {real, imag} */,
  {32'h3e7356ad, 32'h3dc57254} /* (23, 28, 3) {real, imag} */,
  {32'h403e3f20, 32'hc036ddde} /* (23, 28, 2) {real, imag} */,
  {32'hbfcc40d1, 32'h40423c90} /* (23, 28, 1) {real, imag} */,
  {32'hc01b529e, 32'hbf218e94} /* (23, 28, 0) {real, imag} */,
  {32'h400039a0, 32'hc024d11e} /* (23, 27, 31) {real, imag} */,
  {32'hbefae3ee, 32'h3f8f6100} /* (23, 27, 30) {real, imag} */,
  {32'h3e1f5de4, 32'h3f11ecb0} /* (23, 27, 29) {real, imag} */,
  {32'h3e741b86, 32'hbfbd769c} /* (23, 27, 28) {real, imag} */,
  {32'h3c9a0680, 32'h3f61f99c} /* (23, 27, 27) {real, imag} */,
  {32'h3c6b3bc0, 32'hbeff234c} /* (23, 27, 26) {real, imag} */,
  {32'h3b9a4540, 32'h3d370114} /* (23, 27, 25) {real, imag} */,
  {32'h3f46e1f5, 32'hbd3bcd28} /* (23, 27, 24) {real, imag} */,
  {32'hbaa25580, 32'h3dabb5bf} /* (23, 27, 23) {real, imag} */,
  {32'hbed18ac2, 32'h3c5c3ec0} /* (23, 27, 22) {real, imag} */,
  {32'hbeb41078, 32'h3f04a428} /* (23, 27, 21) {real, imag} */,
  {32'hbd9814bd, 32'hbab827e0} /* (23, 27, 20) {real, imag} */,
  {32'hbdac6413, 32'h3e397878} /* (23, 27, 19) {real, imag} */,
  {32'hbc8a9cc0, 32'h3da3d4dd} /* (23, 27, 18) {real, imag} */,
  {32'hbd117420, 32'h3e099dbe} /* (23, 27, 17) {real, imag} */,
  {32'h3db46ed0, 32'hbe9f71ca} /* (23, 27, 16) {real, imag} */,
  {32'hbe34298b, 32'h3d4744bc} /* (23, 27, 15) {real, imag} */,
  {32'h3cc5fcf8, 32'hbe0d26e2} /* (23, 27, 14) {real, imag} */,
  {32'h3e43a10c, 32'hbf00a834} /* (23, 27, 13) {real, imag} */,
  {32'h3d852f14, 32'hbd9a7d22} /* (23, 27, 12) {real, imag} */,
  {32'h3e1c1f36, 32'h3eb7d366} /* (23, 27, 11) {real, imag} */,
  {32'hbe9e4626, 32'h3dbba524} /* (23, 27, 10) {real, imag} */,
  {32'h3f15c50e, 32'hbd98f537} /* (23, 27, 9) {real, imag} */,
  {32'hbd978cf6, 32'hbe57d9aa} /* (23, 27, 8) {real, imag} */,
  {32'h3d83c90d, 32'h3f049993} /* (23, 27, 7) {real, imag} */,
  {32'hbecb39b2, 32'h3dd9ee3c} /* (23, 27, 6) {real, imag} */,
  {32'hbf98a6e6, 32'h3e9e20a0} /* (23, 27, 5) {real, imag} */,
  {32'h3e7b3e3a, 32'h3f4b11bb} /* (23, 27, 4) {real, imag} */,
  {32'h3f51db1b, 32'h3ed32b5d} /* (23, 27, 3) {real, imag} */,
  {32'hbffd2036, 32'hbec5ac7f} /* (23, 27, 2) {real, imag} */,
  {32'h40584026, 32'hbf89b5bd} /* (23, 27, 1) {real, imag} */,
  {32'h40179ddc, 32'hbf8a2077} /* (23, 27, 0) {real, imag} */,
  {32'h3ee78306, 32'hbec1db32} /* (23, 26, 31) {real, imag} */,
  {32'hbec15c35, 32'h3da81fbc} /* (23, 26, 30) {real, imag} */,
  {32'h3eac603a, 32'h3e95a49c} /* (23, 26, 29) {real, imag} */,
  {32'h3f1b5aee, 32'h3ee49fc4} /* (23, 26, 28) {real, imag} */,
  {32'hb96f5e00, 32'hbeebf90a} /* (23, 26, 27) {real, imag} */,
  {32'hbf499020, 32'hbc802df0} /* (23, 26, 26) {real, imag} */,
  {32'hbe8ddbfb, 32'hbedfafae} /* (23, 26, 25) {real, imag} */,
  {32'hbf020dad, 32'h3e2ebc9c} /* (23, 26, 24) {real, imag} */,
  {32'hbd4de19c, 32'hbe4d831d} /* (23, 26, 23) {real, imag} */,
  {32'hbe2fed9e, 32'hbe2e63c2} /* (23, 26, 22) {real, imag} */,
  {32'hbebebffc, 32'hbed59f47} /* (23, 26, 21) {real, imag} */,
  {32'h3d6a1554, 32'h3d6d0980} /* (23, 26, 20) {real, imag} */,
  {32'hbddccd0a, 32'hbdd15180} /* (23, 26, 19) {real, imag} */,
  {32'h3d5b7960, 32'hbe8335c0} /* (23, 26, 18) {real, imag} */,
  {32'h3e317006, 32'hbd300cce} /* (23, 26, 17) {real, imag} */,
  {32'h3da053c4, 32'h3ec5b694} /* (23, 26, 16) {real, imag} */,
  {32'h3e0fde06, 32'h3d4b38dc} /* (23, 26, 15) {real, imag} */,
  {32'h3ed20c32, 32'h3e20bb34} /* (23, 26, 14) {real, imag} */,
  {32'hbeb264af, 32'hbe29ad21} /* (23, 26, 13) {real, imag} */,
  {32'h3ec671de, 32'h3e10ceb2} /* (23, 26, 12) {real, imag} */,
  {32'hbef292ee, 32'h3c1ab3a0} /* (23, 26, 11) {real, imag} */,
  {32'hbec57b56, 32'h3f305815} /* (23, 26, 10) {real, imag} */,
  {32'h3e1e337f, 32'hbe6419b8} /* (23, 26, 9) {real, imag} */,
  {32'hbd1a8b74, 32'hbddf09be} /* (23, 26, 8) {real, imag} */,
  {32'h3e60ce3c, 32'h3dd513eb} /* (23, 26, 7) {real, imag} */,
  {32'hbf668903, 32'hbd8c0338} /* (23, 26, 6) {real, imag} */,
  {32'hbe1f516d, 32'hbf38e9c2} /* (23, 26, 5) {real, imag} */,
  {32'hbba909c0, 32'hbf565081} /* (23, 26, 4) {real, imag} */,
  {32'hbebc4c1c, 32'h3f2384bc} /* (23, 26, 3) {real, imag} */,
  {32'hbdb34f8c, 32'h3e04adf7} /* (23, 26, 2) {real, imag} */,
  {32'h3eb43a3f, 32'h3f479094} /* (23, 26, 1) {real, imag} */,
  {32'h3e2102da, 32'h3e2e895c} /* (23, 26, 0) {real, imag} */,
  {32'hbeb629ee, 32'h3f8501b4} /* (23, 25, 31) {real, imag} */,
  {32'h3f4b8a6c, 32'h3cb32fb0} /* (23, 25, 30) {real, imag} */,
  {32'hbec1d150, 32'hbf2a09f7} /* (23, 25, 29) {real, imag} */,
  {32'h3e8ef746, 32'hbd0f6750} /* (23, 25, 28) {real, imag} */,
  {32'h3d82a37c, 32'hbe127f6f} /* (23, 25, 27) {real, imag} */,
  {32'h3f19dc3c, 32'hbe68b651} /* (23, 25, 26) {real, imag} */,
  {32'h3ec93031, 32'h3e27d049} /* (23, 25, 25) {real, imag} */,
  {32'h3ef68fcc, 32'h3b1bca20} /* (23, 25, 24) {real, imag} */,
  {32'hbe5697fa, 32'h3e8e8c3e} /* (23, 25, 23) {real, imag} */,
  {32'hbe7a8098, 32'hbebe5339} /* (23, 25, 22) {real, imag} */,
  {32'h3e2cb3e1, 32'h3ed78a4d} /* (23, 25, 21) {real, imag} */,
  {32'hbef12f4b, 32'h3e10fb74} /* (23, 25, 20) {real, imag} */,
  {32'h3e720ba2, 32'hbd74b1e0} /* (23, 25, 19) {real, imag} */,
  {32'hbe6ac151, 32'h3d951972} /* (23, 25, 18) {real, imag} */,
  {32'h3de1d248, 32'h3d917d8a} /* (23, 25, 17) {real, imag} */,
  {32'h3e6efa2a, 32'h3ef4e8a6} /* (23, 25, 16) {real, imag} */,
  {32'h3e8ab6e3, 32'h3eff4848} /* (23, 25, 15) {real, imag} */,
  {32'hbe4cd845, 32'hbdb0765c} /* (23, 25, 14) {real, imag} */,
  {32'h3d3e6590, 32'h3d6422bc} /* (23, 25, 13) {real, imag} */,
  {32'h3ea84ace, 32'h3ec451a2} /* (23, 25, 12) {real, imag} */,
  {32'hbd82eabe, 32'hbd2ed48a} /* (23, 25, 11) {real, imag} */,
  {32'h3e811315, 32'hbdca9ef2} /* (23, 25, 10) {real, imag} */,
  {32'h3e95f174, 32'hbdf0079c} /* (23, 25, 9) {real, imag} */,
  {32'h3eef2485, 32'hbeb4965f} /* (23, 25, 8) {real, imag} */,
  {32'hbebd1f38, 32'hbd7c6c08} /* (23, 25, 7) {real, imag} */,
  {32'hbe26fd25, 32'hbf4db741} /* (23, 25, 6) {real, imag} */,
  {32'hbf308a3a, 32'hbdd9bd1e} /* (23, 25, 5) {real, imag} */,
  {32'h3f0a148e, 32'h3d6f9068} /* (23, 25, 4) {real, imag} */,
  {32'h3eb01304, 32'hbedbe9bf} /* (23, 25, 3) {real, imag} */,
  {32'hbe6d11b6, 32'hbeb3f151} /* (23, 25, 2) {real, imag} */,
  {32'hbf91e3b0, 32'h3e949aa7} /* (23, 25, 1) {real, imag} */,
  {32'h3e1e47b3, 32'h3f6edda0} /* (23, 25, 0) {real, imag} */,
  {32'h3d83f8d6, 32'hbf1e10c6} /* (23, 24, 31) {real, imag} */,
  {32'hbf0ff9e0, 32'h3e27689c} /* (23, 24, 30) {real, imag} */,
  {32'h3e6b53a0, 32'h3f13cd37} /* (23, 24, 29) {real, imag} */,
  {32'h3e3057c6, 32'hbe11b212} /* (23, 24, 28) {real, imag} */,
  {32'hbe70d0f6, 32'h3f8079c3} /* (23, 24, 27) {real, imag} */,
  {32'h3c975200, 32'hbf03ea75} /* (23, 24, 26) {real, imag} */,
  {32'h3f8d0358, 32'h3e1775a0} /* (23, 24, 25) {real, imag} */,
  {32'hbef5b386, 32'h3ea563c2} /* (23, 24, 24) {real, imag} */,
  {32'hbd5a6674, 32'h3eac4477} /* (23, 24, 23) {real, imag} */,
  {32'h3f4740e4, 32'hbed5221a} /* (23, 24, 22) {real, imag} */,
  {32'h3e8c3290, 32'h3ea8ac84} /* (23, 24, 21) {real, imag} */,
  {32'hbec14446, 32'hbdf02e25} /* (23, 24, 20) {real, imag} */,
  {32'hbeed2f37, 32'hbec47da2} /* (23, 24, 19) {real, imag} */,
  {32'hbd49f93c, 32'h3e8ae0e8} /* (23, 24, 18) {real, imag} */,
  {32'h3de46d53, 32'hbe06d88c} /* (23, 24, 17) {real, imag} */,
  {32'h3e91cdc1, 32'h3e658322} /* (23, 24, 16) {real, imag} */,
  {32'h3db065b1, 32'h3e516526} /* (23, 24, 15) {real, imag} */,
  {32'hbde4c3f6, 32'hbdb825d6} /* (23, 24, 14) {real, imag} */,
  {32'h3e8944f9, 32'hbe16ae51} /* (23, 24, 13) {real, imag} */,
  {32'hbe5312e0, 32'h3e173606} /* (23, 24, 12) {real, imag} */,
  {32'h3ea64767, 32'h3e5fe905} /* (23, 24, 11) {real, imag} */,
  {32'h3e42664c, 32'h3ed3b718} /* (23, 24, 10) {real, imag} */,
  {32'hbe0f55d2, 32'hbebd71e5} /* (23, 24, 9) {real, imag} */,
  {32'hbf07091e, 32'hbdc0aa8c} /* (23, 24, 8) {real, imag} */,
  {32'h3e77a234, 32'h3f0a31ef} /* (23, 24, 7) {real, imag} */,
  {32'h3e39efba, 32'h3e4b6392} /* (23, 24, 6) {real, imag} */,
  {32'hbec2072e, 32'hbeb3d818} /* (23, 24, 5) {real, imag} */,
  {32'h3e5534c3, 32'h3eeb2516} /* (23, 24, 4) {real, imag} */,
  {32'h3dc6c4c9, 32'hbe4d7145} /* (23, 24, 3) {real, imag} */,
  {32'hbf28028d, 32'h3e1ca0f0} /* (23, 24, 2) {real, imag} */,
  {32'h3fcaaac8, 32'hbf0862db} /* (23, 24, 1) {real, imag} */,
  {32'h3e7f9ee4, 32'hbf26abbc} /* (23, 24, 0) {real, imag} */,
  {32'hbf5e8423, 32'h3f244a91} /* (23, 23, 31) {real, imag} */,
  {32'hbf0c1a68, 32'h3d821c94} /* (23, 23, 30) {real, imag} */,
  {32'hbddf7302, 32'hbdbc2280} /* (23, 23, 29) {real, imag} */,
  {32'hbcde0670, 32'hbe8e6080} /* (23, 23, 28) {real, imag} */,
  {32'hbf08db91, 32'hbdc45ba8} /* (23, 23, 27) {real, imag} */,
  {32'h3dcf040f, 32'h3e017a2d} /* (23, 23, 26) {real, imag} */,
  {32'h3e3dd510, 32'hbe9b9214} /* (23, 23, 25) {real, imag} */,
  {32'h3f3163be, 32'hbf0497e0} /* (23, 23, 24) {real, imag} */,
  {32'hbe4c66d6, 32'hbec1e3a6} /* (23, 23, 23) {real, imag} */,
  {32'h3f50fd49, 32'h3d5a12e8} /* (23, 23, 22) {real, imag} */,
  {32'hbe39bf76, 32'h3e0da08b} /* (23, 23, 21) {real, imag} */,
  {32'h3ef44ef3, 32'hbeecb563} /* (23, 23, 20) {real, imag} */,
  {32'h3e53b34e, 32'h3e4a94c4} /* (23, 23, 19) {real, imag} */,
  {32'h3df436f0, 32'h3df4dd01} /* (23, 23, 18) {real, imag} */,
  {32'h3e96dabc, 32'h3e8f19d0} /* (23, 23, 17) {real, imag} */,
  {32'h3e8fe848, 32'h3e4f384c} /* (23, 23, 16) {real, imag} */,
  {32'hbe958493, 32'h3e151e47} /* (23, 23, 15) {real, imag} */,
  {32'hbe41c57c, 32'hbea4b509} /* (23, 23, 14) {real, imag} */,
  {32'h3e84e7d6, 32'h3ec691ab} /* (23, 23, 13) {real, imag} */,
  {32'h3ed98078, 32'h3e9193e7} /* (23, 23, 12) {real, imag} */,
  {32'hbe6603e4, 32'hbe906264} /* (23, 23, 11) {real, imag} */,
  {32'hbd2a2e0a, 32'hbd428fb4} /* (23, 23, 10) {real, imag} */,
  {32'h3ef49e88, 32'hbe1ccc58} /* (23, 23, 9) {real, imag} */,
  {32'h3df5787c, 32'hbee52dac} /* (23, 23, 8) {real, imag} */,
  {32'h3ccbdd30, 32'hbd88146d} /* (23, 23, 7) {real, imag} */,
  {32'h3edc1db0, 32'h3d51f408} /* (23, 23, 6) {real, imag} */,
  {32'hbd24d36a, 32'hbeeabbab} /* (23, 23, 5) {real, imag} */,
  {32'h3e10384c, 32'hbece81ca} /* (23, 23, 4) {real, imag} */,
  {32'hbf32f509, 32'h3f40a547} /* (23, 23, 3) {real, imag} */,
  {32'h3f1a071a, 32'hbd9d9124} /* (23, 23, 2) {real, imag} */,
  {32'h3f210013, 32'h3f4ba5f4} /* (23, 23, 1) {real, imag} */,
  {32'h3d3e8112, 32'h3e53e839} /* (23, 23, 0) {real, imag} */,
  {32'hbf1fc695, 32'h3cf45190} /* (23, 22, 31) {real, imag} */,
  {32'h3cc9d92c, 32'hbce2e834} /* (23, 22, 30) {real, imag} */,
  {32'h3eae8545, 32'h3e683a47} /* (23, 22, 29) {real, imag} */,
  {32'h3b7c5d00, 32'h3eb66238} /* (23, 22, 28) {real, imag} */,
  {32'h3d489800, 32'hbc24ac40} /* (23, 22, 27) {real, imag} */,
  {32'hbda47d03, 32'hbeefec30} /* (23, 22, 26) {real, imag} */,
  {32'h3e45d82a, 32'hbe6a8747} /* (23, 22, 25) {real, imag} */,
  {32'hbe98212b, 32'h3c363370} /* (23, 22, 24) {real, imag} */,
  {32'h3eb51d48, 32'h3f52cad0} /* (23, 22, 23) {real, imag} */,
  {32'h3f17c04d, 32'hbeb261e2} /* (23, 22, 22) {real, imag} */,
  {32'hbe9551a2, 32'hbe109df8} /* (23, 22, 21) {real, imag} */,
  {32'h3f06a381, 32'h3e298d43} /* (23, 22, 20) {real, imag} */,
  {32'h3deb2684, 32'hbf01aac9} /* (23, 22, 19) {real, imag} */,
  {32'hbe4a4faa, 32'h3cd85c40} /* (23, 22, 18) {real, imag} */,
  {32'hbde0f2a2, 32'h3e5a4a65} /* (23, 22, 17) {real, imag} */,
  {32'hbeeccbdc, 32'h3e4d517e} /* (23, 22, 16) {real, imag} */,
  {32'hbbcc13d0, 32'hbe3605a7} /* (23, 22, 15) {real, imag} */,
  {32'hbe1a2e02, 32'hbe7e8862} /* (23, 22, 14) {real, imag} */,
  {32'h3f1ff176, 32'h3eaf7e65} /* (23, 22, 13) {real, imag} */,
  {32'h3d84956e, 32'hbd5c7180} /* (23, 22, 12) {real, imag} */,
  {32'hbd82cf88, 32'hbe6375e2} /* (23, 22, 11) {real, imag} */,
  {32'hbf0efa9a, 32'h3e0e1bf4} /* (23, 22, 10) {real, imag} */,
  {32'hbd065ba4, 32'h3d892bce} /* (23, 22, 9) {real, imag} */,
  {32'h3f16431c, 32'h3e756f04} /* (23, 22, 8) {real, imag} */,
  {32'hbdb80269, 32'hbeb63736} /* (23, 22, 7) {real, imag} */,
  {32'h3e67568a, 32'hbe49614d} /* (23, 22, 6) {real, imag} */,
  {32'hbf0ed951, 32'hbe919af3} /* (23, 22, 5) {real, imag} */,
  {32'hbeb1ce43, 32'h3f425cd3} /* (23, 22, 4) {real, imag} */,
  {32'hbf374276, 32'h3f2a6572} /* (23, 22, 3) {real, imag} */,
  {32'h3dc528ef, 32'hbf580256} /* (23, 22, 2) {real, imag} */,
  {32'hbada6a00, 32'h3efa9897} /* (23, 22, 1) {real, imag} */,
  {32'h3eff8c26, 32'h3e0da9b5} /* (23, 22, 0) {real, imag} */,
  {32'h3e9bcc05, 32'hbe36a45c} /* (23, 21, 31) {real, imag} */,
  {32'hbe213562, 32'h3e864a30} /* (23, 21, 30) {real, imag} */,
  {32'hbda1b0fc, 32'h3e89bf44} /* (23, 21, 29) {real, imag} */,
  {32'hbcf83680, 32'h3ed0c79f} /* (23, 21, 28) {real, imag} */,
  {32'hbef49d32, 32'h3e8df234} /* (23, 21, 27) {real, imag} */,
  {32'hbe8801de, 32'h3e3f5433} /* (23, 21, 26) {real, imag} */,
  {32'h3e273f40, 32'hbec24341} /* (23, 21, 25) {real, imag} */,
  {32'hbeffd908, 32'hbe23317f} /* (23, 21, 24) {real, imag} */,
  {32'hbe27df44, 32'h3e388676} /* (23, 21, 23) {real, imag} */,
  {32'hbea814f7, 32'h3b9ba020} /* (23, 21, 22) {real, imag} */,
  {32'h3f2629bc, 32'hbe8f51e8} /* (23, 21, 21) {real, imag} */,
  {32'h3e9d9f72, 32'h3e0c48a0} /* (23, 21, 20) {real, imag} */,
  {32'h3ef686ea, 32'hbe185315} /* (23, 21, 19) {real, imag} */,
  {32'hbf246324, 32'h3f3071cf} /* (23, 21, 18) {real, imag} */,
  {32'hbe1d5ed1, 32'hbedd00a4} /* (23, 21, 17) {real, imag} */,
  {32'hbdedcba7, 32'h3dba8d5e} /* (23, 21, 16) {real, imag} */,
  {32'hbd14be2c, 32'hbd27a26f} /* (23, 21, 15) {real, imag} */,
  {32'hbf05a0c4, 32'hbf18019c} /* (23, 21, 14) {real, imag} */,
  {32'hbed2d5b3, 32'hbea1684a} /* (23, 21, 13) {real, imag} */,
  {32'hbdf70446, 32'h3e500d26} /* (23, 21, 12) {real, imag} */,
  {32'hbe96f9c2, 32'hbdd746dc} /* (23, 21, 11) {real, imag} */,
  {32'h3e928706, 32'h3e021792} /* (23, 21, 10) {real, imag} */,
  {32'h3f01ebcc, 32'h3ece4f21} /* (23, 21, 9) {real, imag} */,
  {32'hbeb7d229, 32'h3cd56248} /* (23, 21, 8) {real, imag} */,
  {32'hbe29b6fb, 32'h3d5e8bc0} /* (23, 21, 7) {real, imag} */,
  {32'hbd452294, 32'h3f346e8d} /* (23, 21, 6) {real, imag} */,
  {32'hbedec663, 32'h3e0475e2} /* (23, 21, 5) {real, imag} */,
  {32'h3dd08d85, 32'h3e92469a} /* (23, 21, 4) {real, imag} */,
  {32'hbe51b5aa, 32'hbeb81fb4} /* (23, 21, 3) {real, imag} */,
  {32'hbe07d698, 32'h3eb67c3a} /* (23, 21, 2) {real, imag} */,
  {32'h3f154da5, 32'hbf3c4463} /* (23, 21, 1) {real, imag} */,
  {32'h3dd03828, 32'hbea3d91e} /* (23, 21, 0) {real, imag} */,
  {32'hbe6d7d63, 32'hbe615068} /* (23, 20, 31) {real, imag} */,
  {32'hbe112fae, 32'hbda2d708} /* (23, 20, 30) {real, imag} */,
  {32'hbdeabfcc, 32'h3e92214f} /* (23, 20, 29) {real, imag} */,
  {32'h3e70ad78, 32'hbcd70f3c} /* (23, 20, 28) {real, imag} */,
  {32'hbf0bd314, 32'hbdb435c0} /* (23, 20, 27) {real, imag} */,
  {32'hbe5f2638, 32'hbd544f78} /* (23, 20, 26) {real, imag} */,
  {32'h3e8c3f7c, 32'h3de04710} /* (23, 20, 25) {real, imag} */,
  {32'h3ede61be, 32'h3f1f1f38} /* (23, 20, 24) {real, imag} */,
  {32'hbec64232, 32'hbd882819} /* (23, 20, 23) {real, imag} */,
  {32'h3e52286a, 32'h3e06b5f2} /* (23, 20, 22) {real, imag} */,
  {32'hbbc299d8, 32'hbf1a112d} /* (23, 20, 21) {real, imag} */,
  {32'hbdccac5a, 32'hbeb0dbf5} /* (23, 20, 20) {real, imag} */,
  {32'hbe8b13a8, 32'hbe893162} /* (23, 20, 19) {real, imag} */,
  {32'h3c86de9c, 32'hbe9d5994} /* (23, 20, 18) {real, imag} */,
  {32'hbe85fefd, 32'hbe60b11c} /* (23, 20, 17) {real, imag} */,
  {32'h3db65234, 32'h3e6ed2a4} /* (23, 20, 16) {real, imag} */,
  {32'hbd2319ae, 32'h3e4bf318} /* (23, 20, 15) {real, imag} */,
  {32'hbca50280, 32'h3e93ba91} /* (23, 20, 14) {real, imag} */,
  {32'h3e4b35d0, 32'hbe95cff6} /* (23, 20, 13) {real, imag} */,
  {32'hbeed116e, 32'hbebbe564} /* (23, 20, 12) {real, imag} */,
  {32'hbf1edfd8, 32'hbeb581f4} /* (23, 20, 11) {real, imag} */,
  {32'hbeae0e46, 32'h3ebc00e9} /* (23, 20, 10) {real, imag} */,
  {32'h3e51b3c3, 32'hbe32b777} /* (23, 20, 9) {real, imag} */,
  {32'hbf0c1934, 32'h3eb04854} /* (23, 20, 8) {real, imag} */,
  {32'hbcf7ee30, 32'hbe07bc00} /* (23, 20, 7) {real, imag} */,
  {32'h3ed20aa8, 32'h3ca30a9c} /* (23, 20, 6) {real, imag} */,
  {32'h3d502188, 32'h3f6adbe4} /* (23, 20, 5) {real, imag} */,
  {32'hbdd888d1, 32'hbe913f30} /* (23, 20, 4) {real, imag} */,
  {32'h3e6faa7a, 32'hbdc229b1} /* (23, 20, 3) {real, imag} */,
  {32'hbd8db6be, 32'h3dc66e59} /* (23, 20, 2) {real, imag} */,
  {32'hbf0ed755, 32'h3e839ec7} /* (23, 20, 1) {real, imag} */,
  {32'h3d40d6f8, 32'h3f240fbd} /* (23, 20, 0) {real, imag} */,
  {32'h3e9b5912, 32'hbea66dfc} /* (23, 19, 31) {real, imag} */,
  {32'h3e705f88, 32'hbf322541} /* (23, 19, 30) {real, imag} */,
  {32'hbe453d6a, 32'hbe4a8099} /* (23, 19, 29) {real, imag} */,
  {32'h3cbee2be, 32'hbe8de438} /* (23, 19, 28) {real, imag} */,
  {32'h3dafe6c2, 32'h3cd767cc} /* (23, 19, 27) {real, imag} */,
  {32'h3cb2712e, 32'h3e3dc21c} /* (23, 19, 26) {real, imag} */,
  {32'hbef47bac, 32'hbe732a11} /* (23, 19, 25) {real, imag} */,
  {32'h3c3933d0, 32'h3b3b0000} /* (23, 19, 24) {real, imag} */,
  {32'hbe40e140, 32'h3ec7743c} /* (23, 19, 23) {real, imag} */,
  {32'h3e7c0caf, 32'hbea27a52} /* (23, 19, 22) {real, imag} */,
  {32'hbe774a92, 32'hbd5d8e6a} /* (23, 19, 21) {real, imag} */,
  {32'h3edc92d4, 32'hbc9fb838} /* (23, 19, 20) {real, imag} */,
  {32'hbdaeab08, 32'h3e68d470} /* (23, 19, 19) {real, imag} */,
  {32'hbd372488, 32'h3e86d63b} /* (23, 19, 18) {real, imag} */,
  {32'hbd290e36, 32'hbe2d8f02} /* (23, 19, 17) {real, imag} */,
  {32'h3e3b5e0d, 32'hbe265a76} /* (23, 19, 16) {real, imag} */,
  {32'hbd9611eb, 32'hbdae3254} /* (23, 19, 15) {real, imag} */,
  {32'hbe97e093, 32'hbe2941d2} /* (23, 19, 14) {real, imag} */,
  {32'hbe79cc84, 32'hbc77ba78} /* (23, 19, 13) {real, imag} */,
  {32'h3ece3db2, 32'hbe9f7e3a} /* (23, 19, 12) {real, imag} */,
  {32'hbee262cf, 32'h3f07098a} /* (23, 19, 11) {real, imag} */,
  {32'h3d8b25b8, 32'h3e4a0a27} /* (23, 19, 10) {real, imag} */,
  {32'h3f0e5b4e, 32'hbe7d20e2} /* (23, 19, 9) {real, imag} */,
  {32'h3d169b5d, 32'hbd8453f1} /* (23, 19, 8) {real, imag} */,
  {32'h3e224622, 32'hbeb52820} /* (23, 19, 7) {real, imag} */,
  {32'h3ec2abae, 32'h3effef97} /* (23, 19, 6) {real, imag} */,
  {32'h3f172d9b, 32'hbe880e04} /* (23, 19, 5) {real, imag} */,
  {32'h3eaea246, 32'h3ce833f4} /* (23, 19, 4) {real, imag} */,
  {32'h3e395e8d, 32'h3e35e2c3} /* (23, 19, 3) {real, imag} */,
  {32'hbf4e7c2c, 32'hbd516718} /* (23, 19, 2) {real, imag} */,
  {32'h3e6a26fc, 32'hbebd4e17} /* (23, 19, 1) {real, imag} */,
  {32'hbe537e0a, 32'h3ee70947} /* (23, 19, 0) {real, imag} */,
  {32'hbe0b98d2, 32'hbea0d4e4} /* (23, 18, 31) {real, imag} */,
  {32'hbce30540, 32'h3ea8b452} /* (23, 18, 30) {real, imag} */,
  {32'hbbfb7ff0, 32'h3c727740} /* (23, 18, 29) {real, imag} */,
  {32'h3dd79092, 32'hbd9cfe96} /* (23, 18, 28) {real, imag} */,
  {32'hbe0510b3, 32'h3ecf0666} /* (23, 18, 27) {real, imag} */,
  {32'h3eb379a0, 32'h3deb35fe} /* (23, 18, 26) {real, imag} */,
  {32'h3e4b054c, 32'hbe927deb} /* (23, 18, 25) {real, imag} */,
  {32'hbe1c417e, 32'h3e83bfaa} /* (23, 18, 24) {real, imag} */,
  {32'hbd9deeff, 32'hbdab4268} /* (23, 18, 23) {real, imag} */,
  {32'h3ea488a7, 32'h3ea16c4a} /* (23, 18, 22) {real, imag} */,
  {32'h3e9351dc, 32'hbe09c932} /* (23, 18, 21) {real, imag} */,
  {32'hbd4b00c2, 32'hbb9001d8} /* (23, 18, 20) {real, imag} */,
  {32'h3eb19ea8, 32'h3ed7ce84} /* (23, 18, 19) {real, imag} */,
  {32'hbeb24eb7, 32'hbe23b68e} /* (23, 18, 18) {real, imag} */,
  {32'hbe943a89, 32'h3eb0bf8e} /* (23, 18, 17) {real, imag} */,
  {32'hbe322127, 32'h3e30743b} /* (23, 18, 16) {real, imag} */,
  {32'h3e6d2533, 32'hbd15cce8} /* (23, 18, 15) {real, imag} */,
  {32'h3ea45ecd, 32'h3df65cb0} /* (23, 18, 14) {real, imag} */,
  {32'hbe920387, 32'h3e72f14b} /* (23, 18, 13) {real, imag} */,
  {32'h3e88e2c9, 32'hbe9304ad} /* (23, 18, 12) {real, imag} */,
  {32'hbef8b687, 32'hbe192e73} /* (23, 18, 11) {real, imag} */,
  {32'hbe36d886, 32'hbf21a630} /* (23, 18, 10) {real, imag} */,
  {32'h3e986e84, 32'hbe84b105} /* (23, 18, 9) {real, imag} */,
  {32'h3db8c3dc, 32'h3d760cfa} /* (23, 18, 8) {real, imag} */,
  {32'h3e81a9e6, 32'hbd86ff0e} /* (23, 18, 7) {real, imag} */,
  {32'hbefbe4ec, 32'hbde1bb52} /* (23, 18, 6) {real, imag} */,
  {32'h3cb090a0, 32'hbc17b1c0} /* (23, 18, 5) {real, imag} */,
  {32'h3d932bd4, 32'h3e3a927f} /* (23, 18, 4) {real, imag} */,
  {32'h3cf57172, 32'h3d0a25b4} /* (23, 18, 3) {real, imag} */,
  {32'h3e34f5e6, 32'hbe0eb254} /* (23, 18, 2) {real, imag} */,
  {32'h3e3ad86f, 32'hbf022e1e} /* (23, 18, 1) {real, imag} */,
  {32'hbe4d8886, 32'hbe0b148e} /* (23, 18, 0) {real, imag} */,
  {32'h3e6ab760, 32'h3e5a3be8} /* (23, 17, 31) {real, imag} */,
  {32'h3e9efce7, 32'hbe692ebc} /* (23, 17, 30) {real, imag} */,
  {32'hbe72e244, 32'hbe4c8a80} /* (23, 17, 29) {real, imag} */,
  {32'h3d34be6c, 32'hbe5d1c41} /* (23, 17, 28) {real, imag} */,
  {32'h3d8c6cb3, 32'hbec87ca6} /* (23, 17, 27) {real, imag} */,
  {32'h3f3947fd, 32'h3d57bc60} /* (23, 17, 26) {real, imag} */,
  {32'h3cbcbeb0, 32'hbdb2224c} /* (23, 17, 25) {real, imag} */,
  {32'hbd895e00, 32'hbe6bd61a} /* (23, 17, 24) {real, imag} */,
  {32'h3e14cfb4, 32'h3ec3ee50} /* (23, 17, 23) {real, imag} */,
  {32'hbe75f204, 32'hbe167312} /* (23, 17, 22) {real, imag} */,
  {32'hbe94d7e4, 32'h3d7fff34} /* (23, 17, 21) {real, imag} */,
  {32'hbe93adf6, 32'h3e8b053e} /* (23, 17, 20) {real, imag} */,
  {32'hbedbc0d9, 32'hbd0dee46} /* (23, 17, 19) {real, imag} */,
  {32'h3de92bb7, 32'h3dae3c02} /* (23, 17, 18) {real, imag} */,
  {32'h3e45c55f, 32'h3d97ffad} /* (23, 17, 17) {real, imag} */,
  {32'h3d265b1a, 32'hbdc47d06} /* (23, 17, 16) {real, imag} */,
  {32'hbdc299e3, 32'h3d24a818} /* (23, 17, 15) {real, imag} */,
  {32'h3ed49fc6, 32'h3e46df48} /* (23, 17, 14) {real, imag} */,
  {32'hbe914fbd, 32'hbdd1cbe9} /* (23, 17, 13) {real, imag} */,
  {32'h3e84eb9b, 32'hbe7d426b} /* (23, 17, 12) {real, imag} */,
  {32'h3e11b278, 32'h3e316cbd} /* (23, 17, 11) {real, imag} */,
  {32'h3eb85939, 32'hbd7d8700} /* (23, 17, 10) {real, imag} */,
  {32'hbe5f5f71, 32'h3f0e477a} /* (23, 17, 9) {real, imag} */,
  {32'hbea75328, 32'h3e3ab348} /* (23, 17, 8) {real, imag} */,
  {32'h3ebb9648, 32'hbe04a71e} /* (23, 17, 7) {real, imag} */,
  {32'hbd0d911c, 32'h3d864c8e} /* (23, 17, 6) {real, imag} */,
  {32'h3dad8f47, 32'hbe83e321} /* (23, 17, 5) {real, imag} */,
  {32'hbe76ad3a, 32'hbcedacda} /* (23, 17, 4) {real, imag} */,
  {32'hbeaf631d, 32'hbe21e4dc} /* (23, 17, 3) {real, imag} */,
  {32'h3ed9de60, 32'hbebc52d5} /* (23, 17, 2) {real, imag} */,
  {32'hbd334d9c, 32'h3ecd2207} /* (23, 17, 1) {real, imag} */,
  {32'hbf18aa52, 32'h3e8d3607} /* (23, 17, 0) {real, imag} */,
  {32'h3e12e74a, 32'h3ebf1b57} /* (23, 16, 31) {real, imag} */,
  {32'hbd8ea486, 32'hbea5a2ab} /* (23, 16, 30) {real, imag} */,
  {32'h3e3565a6, 32'h3d7079c7} /* (23, 16, 29) {real, imag} */,
  {32'h3e02fe6e, 32'h3d9b0f1e} /* (23, 16, 28) {real, imag} */,
  {32'hbe09acdb, 32'hbe2718b0} /* (23, 16, 27) {real, imag} */,
  {32'h3d0e4a22, 32'hbe8e3582} /* (23, 16, 26) {real, imag} */,
  {32'hbebda1bb, 32'h3e5075bd} /* (23, 16, 25) {real, imag} */,
  {32'h3c89fa46, 32'h3ed55777} /* (23, 16, 24) {real, imag} */,
  {32'hbe6be3ea, 32'h3e1c8bf6} /* (23, 16, 23) {real, imag} */,
  {32'hbbdb23c0, 32'hbdfc8240} /* (23, 16, 22) {real, imag} */,
  {32'hbeb06a22, 32'h3e8fd13c} /* (23, 16, 21) {real, imag} */,
  {32'hbdff98e8, 32'hbeb8a13c} /* (23, 16, 20) {real, imag} */,
  {32'h3ec548ce, 32'h3f053cce} /* (23, 16, 19) {real, imag} */,
  {32'h3e8f0366, 32'h3d8dc819} /* (23, 16, 18) {real, imag} */,
  {32'hbd1aa0a3, 32'hbe2511e0} /* (23, 16, 17) {real, imag} */,
  {32'h3f060335, 32'h00000000} /* (23, 16, 16) {real, imag} */,
  {32'hbd1aa0a3, 32'h3e2511e0} /* (23, 16, 15) {real, imag} */,
  {32'h3e8f0366, 32'hbd8dc819} /* (23, 16, 14) {real, imag} */,
  {32'h3ec548ce, 32'hbf053cce} /* (23, 16, 13) {real, imag} */,
  {32'hbdff98e8, 32'h3eb8a13c} /* (23, 16, 12) {real, imag} */,
  {32'hbeb06a22, 32'hbe8fd13c} /* (23, 16, 11) {real, imag} */,
  {32'hbbdb23c0, 32'h3dfc8240} /* (23, 16, 10) {real, imag} */,
  {32'hbe6be3ea, 32'hbe1c8bf6} /* (23, 16, 9) {real, imag} */,
  {32'h3c89fa46, 32'hbed55777} /* (23, 16, 8) {real, imag} */,
  {32'hbebda1bb, 32'hbe5075bd} /* (23, 16, 7) {real, imag} */,
  {32'h3d0e4a22, 32'h3e8e3582} /* (23, 16, 6) {real, imag} */,
  {32'hbe09acdb, 32'h3e2718b0} /* (23, 16, 5) {real, imag} */,
  {32'h3e02fe6e, 32'hbd9b0f1e} /* (23, 16, 4) {real, imag} */,
  {32'h3e3565a6, 32'hbd7079c7} /* (23, 16, 3) {real, imag} */,
  {32'hbd8ea486, 32'h3ea5a2ab} /* (23, 16, 2) {real, imag} */,
  {32'h3e12e74a, 32'hbebf1b57} /* (23, 16, 1) {real, imag} */,
  {32'h3e8a6e47, 32'h00000000} /* (23, 16, 0) {real, imag} */,
  {32'hbd334d9c, 32'hbecd2207} /* (23, 15, 31) {real, imag} */,
  {32'h3ed9de60, 32'h3ebc52d5} /* (23, 15, 30) {real, imag} */,
  {32'hbeaf631d, 32'h3e21e4dc} /* (23, 15, 29) {real, imag} */,
  {32'hbe76ad3a, 32'h3cedacda} /* (23, 15, 28) {real, imag} */,
  {32'h3dad8f47, 32'h3e83e321} /* (23, 15, 27) {real, imag} */,
  {32'hbd0d911c, 32'hbd864c8e} /* (23, 15, 26) {real, imag} */,
  {32'h3ebb9648, 32'h3e04a71e} /* (23, 15, 25) {real, imag} */,
  {32'hbea75328, 32'hbe3ab348} /* (23, 15, 24) {real, imag} */,
  {32'hbe5f5f71, 32'hbf0e477a} /* (23, 15, 23) {real, imag} */,
  {32'h3eb85939, 32'h3d7d8700} /* (23, 15, 22) {real, imag} */,
  {32'h3e11b278, 32'hbe316cbd} /* (23, 15, 21) {real, imag} */,
  {32'h3e84eb9b, 32'h3e7d426b} /* (23, 15, 20) {real, imag} */,
  {32'hbe914fbd, 32'h3dd1cbe9} /* (23, 15, 19) {real, imag} */,
  {32'h3ed49fc6, 32'hbe46df48} /* (23, 15, 18) {real, imag} */,
  {32'hbdc299e3, 32'hbd24a818} /* (23, 15, 17) {real, imag} */,
  {32'h3d265b1a, 32'h3dc47d06} /* (23, 15, 16) {real, imag} */,
  {32'h3e45c55f, 32'hbd97ffad} /* (23, 15, 15) {real, imag} */,
  {32'h3de92bb7, 32'hbdae3c02} /* (23, 15, 14) {real, imag} */,
  {32'hbedbc0d9, 32'h3d0dee46} /* (23, 15, 13) {real, imag} */,
  {32'hbe93adf6, 32'hbe8b053e} /* (23, 15, 12) {real, imag} */,
  {32'hbe94d7e4, 32'hbd7fff34} /* (23, 15, 11) {real, imag} */,
  {32'hbe75f204, 32'h3e167312} /* (23, 15, 10) {real, imag} */,
  {32'h3e14cfb4, 32'hbec3ee50} /* (23, 15, 9) {real, imag} */,
  {32'hbd895e00, 32'h3e6bd61a} /* (23, 15, 8) {real, imag} */,
  {32'h3cbcbeb0, 32'h3db2224c} /* (23, 15, 7) {real, imag} */,
  {32'h3f3947fd, 32'hbd57bc60} /* (23, 15, 6) {real, imag} */,
  {32'h3d8c6cb3, 32'h3ec87ca6} /* (23, 15, 5) {real, imag} */,
  {32'h3d34be6c, 32'h3e5d1c41} /* (23, 15, 4) {real, imag} */,
  {32'hbe72e244, 32'h3e4c8a80} /* (23, 15, 3) {real, imag} */,
  {32'h3e9efce7, 32'h3e692ebc} /* (23, 15, 2) {real, imag} */,
  {32'h3e6ab760, 32'hbe5a3be8} /* (23, 15, 1) {real, imag} */,
  {32'hbf18aa52, 32'hbe8d3607} /* (23, 15, 0) {real, imag} */,
  {32'h3e3ad86f, 32'h3f022e1e} /* (23, 14, 31) {real, imag} */,
  {32'h3e34f5e6, 32'h3e0eb254} /* (23, 14, 30) {real, imag} */,
  {32'h3cf57172, 32'hbd0a25b4} /* (23, 14, 29) {real, imag} */,
  {32'h3d932bd4, 32'hbe3a927f} /* (23, 14, 28) {real, imag} */,
  {32'h3cb090a0, 32'h3c17b1c0} /* (23, 14, 27) {real, imag} */,
  {32'hbefbe4ec, 32'h3de1bb52} /* (23, 14, 26) {real, imag} */,
  {32'h3e81a9e6, 32'h3d86ff0e} /* (23, 14, 25) {real, imag} */,
  {32'h3db8c3dc, 32'hbd760cfa} /* (23, 14, 24) {real, imag} */,
  {32'h3e986e84, 32'h3e84b105} /* (23, 14, 23) {real, imag} */,
  {32'hbe36d886, 32'h3f21a630} /* (23, 14, 22) {real, imag} */,
  {32'hbef8b687, 32'h3e192e73} /* (23, 14, 21) {real, imag} */,
  {32'h3e88e2c9, 32'h3e9304ad} /* (23, 14, 20) {real, imag} */,
  {32'hbe920387, 32'hbe72f14b} /* (23, 14, 19) {real, imag} */,
  {32'h3ea45ecd, 32'hbdf65cb0} /* (23, 14, 18) {real, imag} */,
  {32'h3e6d2533, 32'h3d15cce8} /* (23, 14, 17) {real, imag} */,
  {32'hbe322127, 32'hbe30743b} /* (23, 14, 16) {real, imag} */,
  {32'hbe943a89, 32'hbeb0bf8e} /* (23, 14, 15) {real, imag} */,
  {32'hbeb24eb7, 32'h3e23b68e} /* (23, 14, 14) {real, imag} */,
  {32'h3eb19ea8, 32'hbed7ce84} /* (23, 14, 13) {real, imag} */,
  {32'hbd4b00c2, 32'h3b9001d8} /* (23, 14, 12) {real, imag} */,
  {32'h3e9351dc, 32'h3e09c932} /* (23, 14, 11) {real, imag} */,
  {32'h3ea488a7, 32'hbea16c4a} /* (23, 14, 10) {real, imag} */,
  {32'hbd9deeff, 32'h3dab4268} /* (23, 14, 9) {real, imag} */,
  {32'hbe1c417e, 32'hbe83bfaa} /* (23, 14, 8) {real, imag} */,
  {32'h3e4b054c, 32'h3e927deb} /* (23, 14, 7) {real, imag} */,
  {32'h3eb379a0, 32'hbdeb35fe} /* (23, 14, 6) {real, imag} */,
  {32'hbe0510b3, 32'hbecf0666} /* (23, 14, 5) {real, imag} */,
  {32'h3dd79092, 32'h3d9cfe96} /* (23, 14, 4) {real, imag} */,
  {32'hbbfb7ff0, 32'hbc727740} /* (23, 14, 3) {real, imag} */,
  {32'hbce30540, 32'hbea8b452} /* (23, 14, 2) {real, imag} */,
  {32'hbe0b98d2, 32'h3ea0d4e4} /* (23, 14, 1) {real, imag} */,
  {32'hbe4d8886, 32'h3e0b148e} /* (23, 14, 0) {real, imag} */,
  {32'h3e6a26fc, 32'h3ebd4e17} /* (23, 13, 31) {real, imag} */,
  {32'hbf4e7c2c, 32'h3d516718} /* (23, 13, 30) {real, imag} */,
  {32'h3e395e8d, 32'hbe35e2c3} /* (23, 13, 29) {real, imag} */,
  {32'h3eaea246, 32'hbce833f4} /* (23, 13, 28) {real, imag} */,
  {32'h3f172d9b, 32'h3e880e04} /* (23, 13, 27) {real, imag} */,
  {32'h3ec2abae, 32'hbeffef97} /* (23, 13, 26) {real, imag} */,
  {32'h3e224622, 32'h3eb52820} /* (23, 13, 25) {real, imag} */,
  {32'h3d169b5d, 32'h3d8453f1} /* (23, 13, 24) {real, imag} */,
  {32'h3f0e5b4e, 32'h3e7d20e2} /* (23, 13, 23) {real, imag} */,
  {32'h3d8b25b8, 32'hbe4a0a27} /* (23, 13, 22) {real, imag} */,
  {32'hbee262cf, 32'hbf07098a} /* (23, 13, 21) {real, imag} */,
  {32'h3ece3db2, 32'h3e9f7e3a} /* (23, 13, 20) {real, imag} */,
  {32'hbe79cc84, 32'h3c77ba78} /* (23, 13, 19) {real, imag} */,
  {32'hbe97e093, 32'h3e2941d2} /* (23, 13, 18) {real, imag} */,
  {32'hbd9611eb, 32'h3dae3254} /* (23, 13, 17) {real, imag} */,
  {32'h3e3b5e0d, 32'h3e265a76} /* (23, 13, 16) {real, imag} */,
  {32'hbd290e36, 32'h3e2d8f02} /* (23, 13, 15) {real, imag} */,
  {32'hbd372488, 32'hbe86d63b} /* (23, 13, 14) {real, imag} */,
  {32'hbdaeab08, 32'hbe68d470} /* (23, 13, 13) {real, imag} */,
  {32'h3edc92d4, 32'h3c9fb838} /* (23, 13, 12) {real, imag} */,
  {32'hbe774a92, 32'h3d5d8e6a} /* (23, 13, 11) {real, imag} */,
  {32'h3e7c0caf, 32'h3ea27a52} /* (23, 13, 10) {real, imag} */,
  {32'hbe40e140, 32'hbec7743c} /* (23, 13, 9) {real, imag} */,
  {32'h3c3933d0, 32'hbb3b0000} /* (23, 13, 8) {real, imag} */,
  {32'hbef47bac, 32'h3e732a11} /* (23, 13, 7) {real, imag} */,
  {32'h3cb2712e, 32'hbe3dc21c} /* (23, 13, 6) {real, imag} */,
  {32'h3dafe6c2, 32'hbcd767cc} /* (23, 13, 5) {real, imag} */,
  {32'h3cbee2be, 32'h3e8de438} /* (23, 13, 4) {real, imag} */,
  {32'hbe453d6a, 32'h3e4a8099} /* (23, 13, 3) {real, imag} */,
  {32'h3e705f88, 32'h3f322541} /* (23, 13, 2) {real, imag} */,
  {32'h3e9b5912, 32'h3ea66dfc} /* (23, 13, 1) {real, imag} */,
  {32'hbe537e0a, 32'hbee70947} /* (23, 13, 0) {real, imag} */,
  {32'hbf0ed755, 32'hbe839ec7} /* (23, 12, 31) {real, imag} */,
  {32'hbd8db6be, 32'hbdc66e59} /* (23, 12, 30) {real, imag} */,
  {32'h3e6faa7a, 32'h3dc229b1} /* (23, 12, 29) {real, imag} */,
  {32'hbdd888d1, 32'h3e913f30} /* (23, 12, 28) {real, imag} */,
  {32'h3d502188, 32'hbf6adbe4} /* (23, 12, 27) {real, imag} */,
  {32'h3ed20aa8, 32'hbca30a9c} /* (23, 12, 26) {real, imag} */,
  {32'hbcf7ee30, 32'h3e07bc00} /* (23, 12, 25) {real, imag} */,
  {32'hbf0c1934, 32'hbeb04854} /* (23, 12, 24) {real, imag} */,
  {32'h3e51b3c3, 32'h3e32b777} /* (23, 12, 23) {real, imag} */,
  {32'hbeae0e46, 32'hbebc00e9} /* (23, 12, 22) {real, imag} */,
  {32'hbf1edfd8, 32'h3eb581f4} /* (23, 12, 21) {real, imag} */,
  {32'hbeed116e, 32'h3ebbe564} /* (23, 12, 20) {real, imag} */,
  {32'h3e4b35d0, 32'h3e95cff6} /* (23, 12, 19) {real, imag} */,
  {32'hbca50280, 32'hbe93ba91} /* (23, 12, 18) {real, imag} */,
  {32'hbd2319ae, 32'hbe4bf318} /* (23, 12, 17) {real, imag} */,
  {32'h3db65234, 32'hbe6ed2a4} /* (23, 12, 16) {real, imag} */,
  {32'hbe85fefd, 32'h3e60b11c} /* (23, 12, 15) {real, imag} */,
  {32'h3c86de9c, 32'h3e9d5994} /* (23, 12, 14) {real, imag} */,
  {32'hbe8b13a8, 32'h3e893162} /* (23, 12, 13) {real, imag} */,
  {32'hbdccac5a, 32'h3eb0dbf5} /* (23, 12, 12) {real, imag} */,
  {32'hbbc299d8, 32'h3f1a112d} /* (23, 12, 11) {real, imag} */,
  {32'h3e52286a, 32'hbe06b5f2} /* (23, 12, 10) {real, imag} */,
  {32'hbec64232, 32'h3d882819} /* (23, 12, 9) {real, imag} */,
  {32'h3ede61be, 32'hbf1f1f38} /* (23, 12, 8) {real, imag} */,
  {32'h3e8c3f7c, 32'hbde04710} /* (23, 12, 7) {real, imag} */,
  {32'hbe5f2638, 32'h3d544f78} /* (23, 12, 6) {real, imag} */,
  {32'hbf0bd314, 32'h3db435c0} /* (23, 12, 5) {real, imag} */,
  {32'h3e70ad78, 32'h3cd70f3c} /* (23, 12, 4) {real, imag} */,
  {32'hbdeabfcc, 32'hbe92214f} /* (23, 12, 3) {real, imag} */,
  {32'hbe112fae, 32'h3da2d708} /* (23, 12, 2) {real, imag} */,
  {32'hbe6d7d63, 32'h3e615068} /* (23, 12, 1) {real, imag} */,
  {32'h3d40d6f8, 32'hbf240fbd} /* (23, 12, 0) {real, imag} */,
  {32'h3f154da5, 32'h3f3c4463} /* (23, 11, 31) {real, imag} */,
  {32'hbe07d698, 32'hbeb67c3a} /* (23, 11, 30) {real, imag} */,
  {32'hbe51b5aa, 32'h3eb81fb4} /* (23, 11, 29) {real, imag} */,
  {32'h3dd08d85, 32'hbe92469a} /* (23, 11, 28) {real, imag} */,
  {32'hbedec663, 32'hbe0475e2} /* (23, 11, 27) {real, imag} */,
  {32'hbd452294, 32'hbf346e8d} /* (23, 11, 26) {real, imag} */,
  {32'hbe29b6fb, 32'hbd5e8bc0} /* (23, 11, 25) {real, imag} */,
  {32'hbeb7d229, 32'hbcd56248} /* (23, 11, 24) {real, imag} */,
  {32'h3f01ebcc, 32'hbece4f21} /* (23, 11, 23) {real, imag} */,
  {32'h3e928706, 32'hbe021792} /* (23, 11, 22) {real, imag} */,
  {32'hbe96f9c2, 32'h3dd746dc} /* (23, 11, 21) {real, imag} */,
  {32'hbdf70446, 32'hbe500d26} /* (23, 11, 20) {real, imag} */,
  {32'hbed2d5b3, 32'h3ea1684a} /* (23, 11, 19) {real, imag} */,
  {32'hbf05a0c4, 32'h3f18019c} /* (23, 11, 18) {real, imag} */,
  {32'hbd14be2c, 32'h3d27a26f} /* (23, 11, 17) {real, imag} */,
  {32'hbdedcba7, 32'hbdba8d5e} /* (23, 11, 16) {real, imag} */,
  {32'hbe1d5ed1, 32'h3edd00a4} /* (23, 11, 15) {real, imag} */,
  {32'hbf246324, 32'hbf3071cf} /* (23, 11, 14) {real, imag} */,
  {32'h3ef686ea, 32'h3e185315} /* (23, 11, 13) {real, imag} */,
  {32'h3e9d9f72, 32'hbe0c48a0} /* (23, 11, 12) {real, imag} */,
  {32'h3f2629bc, 32'h3e8f51e8} /* (23, 11, 11) {real, imag} */,
  {32'hbea814f7, 32'hbb9ba020} /* (23, 11, 10) {real, imag} */,
  {32'hbe27df44, 32'hbe388676} /* (23, 11, 9) {real, imag} */,
  {32'hbeffd908, 32'h3e23317f} /* (23, 11, 8) {real, imag} */,
  {32'h3e273f40, 32'h3ec24341} /* (23, 11, 7) {real, imag} */,
  {32'hbe8801de, 32'hbe3f5433} /* (23, 11, 6) {real, imag} */,
  {32'hbef49d32, 32'hbe8df234} /* (23, 11, 5) {real, imag} */,
  {32'hbcf83680, 32'hbed0c79f} /* (23, 11, 4) {real, imag} */,
  {32'hbda1b0fc, 32'hbe89bf44} /* (23, 11, 3) {real, imag} */,
  {32'hbe213562, 32'hbe864a30} /* (23, 11, 2) {real, imag} */,
  {32'h3e9bcc05, 32'h3e36a45c} /* (23, 11, 1) {real, imag} */,
  {32'h3dd03828, 32'h3ea3d91e} /* (23, 11, 0) {real, imag} */,
  {32'hbada6a00, 32'hbefa9897} /* (23, 10, 31) {real, imag} */,
  {32'h3dc528ef, 32'h3f580256} /* (23, 10, 30) {real, imag} */,
  {32'hbf374276, 32'hbf2a6572} /* (23, 10, 29) {real, imag} */,
  {32'hbeb1ce43, 32'hbf425cd3} /* (23, 10, 28) {real, imag} */,
  {32'hbf0ed951, 32'h3e919af3} /* (23, 10, 27) {real, imag} */,
  {32'h3e67568a, 32'h3e49614d} /* (23, 10, 26) {real, imag} */,
  {32'hbdb80269, 32'h3eb63736} /* (23, 10, 25) {real, imag} */,
  {32'h3f16431c, 32'hbe756f04} /* (23, 10, 24) {real, imag} */,
  {32'hbd065ba4, 32'hbd892bce} /* (23, 10, 23) {real, imag} */,
  {32'hbf0efa9a, 32'hbe0e1bf4} /* (23, 10, 22) {real, imag} */,
  {32'hbd82cf88, 32'h3e6375e2} /* (23, 10, 21) {real, imag} */,
  {32'h3d84956e, 32'h3d5c7180} /* (23, 10, 20) {real, imag} */,
  {32'h3f1ff176, 32'hbeaf7e65} /* (23, 10, 19) {real, imag} */,
  {32'hbe1a2e02, 32'h3e7e8862} /* (23, 10, 18) {real, imag} */,
  {32'hbbcc13d0, 32'h3e3605a7} /* (23, 10, 17) {real, imag} */,
  {32'hbeeccbdc, 32'hbe4d517e} /* (23, 10, 16) {real, imag} */,
  {32'hbde0f2a2, 32'hbe5a4a65} /* (23, 10, 15) {real, imag} */,
  {32'hbe4a4faa, 32'hbcd85c40} /* (23, 10, 14) {real, imag} */,
  {32'h3deb2684, 32'h3f01aac9} /* (23, 10, 13) {real, imag} */,
  {32'h3f06a381, 32'hbe298d43} /* (23, 10, 12) {real, imag} */,
  {32'hbe9551a2, 32'h3e109df8} /* (23, 10, 11) {real, imag} */,
  {32'h3f17c04d, 32'h3eb261e2} /* (23, 10, 10) {real, imag} */,
  {32'h3eb51d48, 32'hbf52cad0} /* (23, 10, 9) {real, imag} */,
  {32'hbe98212b, 32'hbc363370} /* (23, 10, 8) {real, imag} */,
  {32'h3e45d82a, 32'h3e6a8747} /* (23, 10, 7) {real, imag} */,
  {32'hbda47d03, 32'h3eefec30} /* (23, 10, 6) {real, imag} */,
  {32'h3d489800, 32'h3c24ac40} /* (23, 10, 5) {real, imag} */,
  {32'h3b7c5d00, 32'hbeb66238} /* (23, 10, 4) {real, imag} */,
  {32'h3eae8545, 32'hbe683a47} /* (23, 10, 3) {real, imag} */,
  {32'h3cc9d92c, 32'h3ce2e834} /* (23, 10, 2) {real, imag} */,
  {32'hbf1fc695, 32'hbcf45190} /* (23, 10, 1) {real, imag} */,
  {32'h3eff8c26, 32'hbe0da9b5} /* (23, 10, 0) {real, imag} */,
  {32'h3f210013, 32'hbf4ba5f4} /* (23, 9, 31) {real, imag} */,
  {32'h3f1a071a, 32'h3d9d9124} /* (23, 9, 30) {real, imag} */,
  {32'hbf32f509, 32'hbf40a547} /* (23, 9, 29) {real, imag} */,
  {32'h3e10384c, 32'h3ece81ca} /* (23, 9, 28) {real, imag} */,
  {32'hbd24d36a, 32'h3eeabbab} /* (23, 9, 27) {real, imag} */,
  {32'h3edc1db0, 32'hbd51f408} /* (23, 9, 26) {real, imag} */,
  {32'h3ccbdd30, 32'h3d88146d} /* (23, 9, 25) {real, imag} */,
  {32'h3df5787c, 32'h3ee52dac} /* (23, 9, 24) {real, imag} */,
  {32'h3ef49e88, 32'h3e1ccc58} /* (23, 9, 23) {real, imag} */,
  {32'hbd2a2e0a, 32'h3d428fb4} /* (23, 9, 22) {real, imag} */,
  {32'hbe6603e4, 32'h3e906264} /* (23, 9, 21) {real, imag} */,
  {32'h3ed98078, 32'hbe9193e7} /* (23, 9, 20) {real, imag} */,
  {32'h3e84e7d6, 32'hbec691ab} /* (23, 9, 19) {real, imag} */,
  {32'hbe41c57c, 32'h3ea4b509} /* (23, 9, 18) {real, imag} */,
  {32'hbe958493, 32'hbe151e47} /* (23, 9, 17) {real, imag} */,
  {32'h3e8fe848, 32'hbe4f384c} /* (23, 9, 16) {real, imag} */,
  {32'h3e96dabc, 32'hbe8f19d0} /* (23, 9, 15) {real, imag} */,
  {32'h3df436f0, 32'hbdf4dd01} /* (23, 9, 14) {real, imag} */,
  {32'h3e53b34e, 32'hbe4a94c4} /* (23, 9, 13) {real, imag} */,
  {32'h3ef44ef3, 32'h3eecb563} /* (23, 9, 12) {real, imag} */,
  {32'hbe39bf76, 32'hbe0da08b} /* (23, 9, 11) {real, imag} */,
  {32'h3f50fd49, 32'hbd5a12e8} /* (23, 9, 10) {real, imag} */,
  {32'hbe4c66d6, 32'h3ec1e3a6} /* (23, 9, 9) {real, imag} */,
  {32'h3f3163be, 32'h3f0497e0} /* (23, 9, 8) {real, imag} */,
  {32'h3e3dd510, 32'h3e9b9214} /* (23, 9, 7) {real, imag} */,
  {32'h3dcf040f, 32'hbe017a2d} /* (23, 9, 6) {real, imag} */,
  {32'hbf08db91, 32'h3dc45ba8} /* (23, 9, 5) {real, imag} */,
  {32'hbcde0670, 32'h3e8e6080} /* (23, 9, 4) {real, imag} */,
  {32'hbddf7302, 32'h3dbc2280} /* (23, 9, 3) {real, imag} */,
  {32'hbf0c1a68, 32'hbd821c94} /* (23, 9, 2) {real, imag} */,
  {32'hbf5e8423, 32'hbf244a91} /* (23, 9, 1) {real, imag} */,
  {32'h3d3e8112, 32'hbe53e839} /* (23, 9, 0) {real, imag} */,
  {32'h3fcaaac8, 32'h3f0862db} /* (23, 8, 31) {real, imag} */,
  {32'hbf28028d, 32'hbe1ca0f0} /* (23, 8, 30) {real, imag} */,
  {32'h3dc6c4c9, 32'h3e4d7145} /* (23, 8, 29) {real, imag} */,
  {32'h3e5534c3, 32'hbeeb2516} /* (23, 8, 28) {real, imag} */,
  {32'hbec2072e, 32'h3eb3d818} /* (23, 8, 27) {real, imag} */,
  {32'h3e39efba, 32'hbe4b6392} /* (23, 8, 26) {real, imag} */,
  {32'h3e77a234, 32'hbf0a31ef} /* (23, 8, 25) {real, imag} */,
  {32'hbf07091e, 32'h3dc0aa8c} /* (23, 8, 24) {real, imag} */,
  {32'hbe0f55d2, 32'h3ebd71e5} /* (23, 8, 23) {real, imag} */,
  {32'h3e42664c, 32'hbed3b718} /* (23, 8, 22) {real, imag} */,
  {32'h3ea64767, 32'hbe5fe905} /* (23, 8, 21) {real, imag} */,
  {32'hbe5312e0, 32'hbe173606} /* (23, 8, 20) {real, imag} */,
  {32'h3e8944f9, 32'h3e16ae51} /* (23, 8, 19) {real, imag} */,
  {32'hbde4c3f6, 32'h3db825d6} /* (23, 8, 18) {real, imag} */,
  {32'h3db065b1, 32'hbe516526} /* (23, 8, 17) {real, imag} */,
  {32'h3e91cdc1, 32'hbe658322} /* (23, 8, 16) {real, imag} */,
  {32'h3de46d53, 32'h3e06d88c} /* (23, 8, 15) {real, imag} */,
  {32'hbd49f93c, 32'hbe8ae0e8} /* (23, 8, 14) {real, imag} */,
  {32'hbeed2f37, 32'h3ec47da2} /* (23, 8, 13) {real, imag} */,
  {32'hbec14446, 32'h3df02e25} /* (23, 8, 12) {real, imag} */,
  {32'h3e8c3290, 32'hbea8ac84} /* (23, 8, 11) {real, imag} */,
  {32'h3f4740e4, 32'h3ed5221a} /* (23, 8, 10) {real, imag} */,
  {32'hbd5a6674, 32'hbeac4477} /* (23, 8, 9) {real, imag} */,
  {32'hbef5b386, 32'hbea563c2} /* (23, 8, 8) {real, imag} */,
  {32'h3f8d0358, 32'hbe1775a0} /* (23, 8, 7) {real, imag} */,
  {32'h3c975200, 32'h3f03ea75} /* (23, 8, 6) {real, imag} */,
  {32'hbe70d0f6, 32'hbf8079c3} /* (23, 8, 5) {real, imag} */,
  {32'h3e3057c6, 32'h3e11b212} /* (23, 8, 4) {real, imag} */,
  {32'h3e6b53a0, 32'hbf13cd37} /* (23, 8, 3) {real, imag} */,
  {32'hbf0ff9e0, 32'hbe27689c} /* (23, 8, 2) {real, imag} */,
  {32'h3d83f8d6, 32'h3f1e10c6} /* (23, 8, 1) {real, imag} */,
  {32'h3e7f9ee4, 32'h3f26abbc} /* (23, 8, 0) {real, imag} */,
  {32'hbf91e3b0, 32'hbe949aa7} /* (23, 7, 31) {real, imag} */,
  {32'hbe6d11b6, 32'h3eb3f151} /* (23, 7, 30) {real, imag} */,
  {32'h3eb01304, 32'h3edbe9bf} /* (23, 7, 29) {real, imag} */,
  {32'h3f0a148e, 32'hbd6f9068} /* (23, 7, 28) {real, imag} */,
  {32'hbf308a3a, 32'h3dd9bd1e} /* (23, 7, 27) {real, imag} */,
  {32'hbe26fd25, 32'h3f4db741} /* (23, 7, 26) {real, imag} */,
  {32'hbebd1f38, 32'h3d7c6c08} /* (23, 7, 25) {real, imag} */,
  {32'h3eef2485, 32'h3eb4965f} /* (23, 7, 24) {real, imag} */,
  {32'h3e95f174, 32'h3df0079c} /* (23, 7, 23) {real, imag} */,
  {32'h3e811315, 32'h3dca9ef2} /* (23, 7, 22) {real, imag} */,
  {32'hbd82eabe, 32'h3d2ed48a} /* (23, 7, 21) {real, imag} */,
  {32'h3ea84ace, 32'hbec451a2} /* (23, 7, 20) {real, imag} */,
  {32'h3d3e6590, 32'hbd6422bc} /* (23, 7, 19) {real, imag} */,
  {32'hbe4cd845, 32'h3db0765c} /* (23, 7, 18) {real, imag} */,
  {32'h3e8ab6e3, 32'hbeff4848} /* (23, 7, 17) {real, imag} */,
  {32'h3e6efa2a, 32'hbef4e8a6} /* (23, 7, 16) {real, imag} */,
  {32'h3de1d248, 32'hbd917d8a} /* (23, 7, 15) {real, imag} */,
  {32'hbe6ac151, 32'hbd951972} /* (23, 7, 14) {real, imag} */,
  {32'h3e720ba2, 32'h3d74b1e0} /* (23, 7, 13) {real, imag} */,
  {32'hbef12f4b, 32'hbe10fb74} /* (23, 7, 12) {real, imag} */,
  {32'h3e2cb3e1, 32'hbed78a4d} /* (23, 7, 11) {real, imag} */,
  {32'hbe7a8098, 32'h3ebe5339} /* (23, 7, 10) {real, imag} */,
  {32'hbe5697fa, 32'hbe8e8c3e} /* (23, 7, 9) {real, imag} */,
  {32'h3ef68fcc, 32'hbb1bca20} /* (23, 7, 8) {real, imag} */,
  {32'h3ec93031, 32'hbe27d049} /* (23, 7, 7) {real, imag} */,
  {32'h3f19dc3c, 32'h3e68b651} /* (23, 7, 6) {real, imag} */,
  {32'h3d82a37c, 32'h3e127f6f} /* (23, 7, 5) {real, imag} */,
  {32'h3e8ef746, 32'h3d0f6750} /* (23, 7, 4) {real, imag} */,
  {32'hbec1d150, 32'h3f2a09f7} /* (23, 7, 3) {real, imag} */,
  {32'h3f4b8a6c, 32'hbcb32fb0} /* (23, 7, 2) {real, imag} */,
  {32'hbeb629ee, 32'hbf8501b4} /* (23, 7, 1) {real, imag} */,
  {32'h3e1e47b3, 32'hbf6edda0} /* (23, 7, 0) {real, imag} */,
  {32'h3eb43a3f, 32'hbf479094} /* (23, 6, 31) {real, imag} */,
  {32'hbdb34f8c, 32'hbe04adf7} /* (23, 6, 30) {real, imag} */,
  {32'hbebc4c1c, 32'hbf2384bc} /* (23, 6, 29) {real, imag} */,
  {32'hbba909c0, 32'h3f565081} /* (23, 6, 28) {real, imag} */,
  {32'hbe1f516d, 32'h3f38e9c2} /* (23, 6, 27) {real, imag} */,
  {32'hbf668903, 32'h3d8c0338} /* (23, 6, 26) {real, imag} */,
  {32'h3e60ce3c, 32'hbdd513eb} /* (23, 6, 25) {real, imag} */,
  {32'hbd1a8b74, 32'h3ddf09be} /* (23, 6, 24) {real, imag} */,
  {32'h3e1e337f, 32'h3e6419b8} /* (23, 6, 23) {real, imag} */,
  {32'hbec57b56, 32'hbf305815} /* (23, 6, 22) {real, imag} */,
  {32'hbef292ee, 32'hbc1ab3a0} /* (23, 6, 21) {real, imag} */,
  {32'h3ec671de, 32'hbe10ceb2} /* (23, 6, 20) {real, imag} */,
  {32'hbeb264af, 32'h3e29ad21} /* (23, 6, 19) {real, imag} */,
  {32'h3ed20c32, 32'hbe20bb34} /* (23, 6, 18) {real, imag} */,
  {32'h3e0fde06, 32'hbd4b38dc} /* (23, 6, 17) {real, imag} */,
  {32'h3da053c4, 32'hbec5b694} /* (23, 6, 16) {real, imag} */,
  {32'h3e317006, 32'h3d300cce} /* (23, 6, 15) {real, imag} */,
  {32'h3d5b7960, 32'h3e8335c0} /* (23, 6, 14) {real, imag} */,
  {32'hbddccd0a, 32'h3dd15180} /* (23, 6, 13) {real, imag} */,
  {32'h3d6a1554, 32'hbd6d0980} /* (23, 6, 12) {real, imag} */,
  {32'hbebebffc, 32'h3ed59f47} /* (23, 6, 11) {real, imag} */,
  {32'hbe2fed9e, 32'h3e2e63c2} /* (23, 6, 10) {real, imag} */,
  {32'hbd4de19c, 32'h3e4d831d} /* (23, 6, 9) {real, imag} */,
  {32'hbf020dad, 32'hbe2ebc9c} /* (23, 6, 8) {real, imag} */,
  {32'hbe8ddbfb, 32'h3edfafae} /* (23, 6, 7) {real, imag} */,
  {32'hbf499020, 32'h3c802df0} /* (23, 6, 6) {real, imag} */,
  {32'hb96f5e00, 32'h3eebf90a} /* (23, 6, 5) {real, imag} */,
  {32'h3f1b5aee, 32'hbee49fc4} /* (23, 6, 4) {real, imag} */,
  {32'h3eac603a, 32'hbe95a49c} /* (23, 6, 3) {real, imag} */,
  {32'hbec15c35, 32'hbda81fbc} /* (23, 6, 2) {real, imag} */,
  {32'h3ee78306, 32'h3ec1db32} /* (23, 6, 1) {real, imag} */,
  {32'h3e2102da, 32'hbe2e895c} /* (23, 6, 0) {real, imag} */,
  {32'h40584026, 32'h3f89b5bd} /* (23, 5, 31) {real, imag} */,
  {32'hbffd2036, 32'h3ec5ac7f} /* (23, 5, 30) {real, imag} */,
  {32'h3f51db1b, 32'hbed32b5d} /* (23, 5, 29) {real, imag} */,
  {32'h3e7b3e3a, 32'hbf4b11bb} /* (23, 5, 28) {real, imag} */,
  {32'hbf98a6e6, 32'hbe9e20a0} /* (23, 5, 27) {real, imag} */,
  {32'hbecb39b2, 32'hbdd9ee3c} /* (23, 5, 26) {real, imag} */,
  {32'h3d83c90d, 32'hbf049993} /* (23, 5, 25) {real, imag} */,
  {32'hbd978cf6, 32'h3e57d9aa} /* (23, 5, 24) {real, imag} */,
  {32'h3f15c50e, 32'h3d98f537} /* (23, 5, 23) {real, imag} */,
  {32'hbe9e4626, 32'hbdbba524} /* (23, 5, 22) {real, imag} */,
  {32'h3e1c1f36, 32'hbeb7d366} /* (23, 5, 21) {real, imag} */,
  {32'h3d852f14, 32'h3d9a7d22} /* (23, 5, 20) {real, imag} */,
  {32'h3e43a10c, 32'h3f00a834} /* (23, 5, 19) {real, imag} */,
  {32'h3cc5fcf8, 32'h3e0d26e2} /* (23, 5, 18) {real, imag} */,
  {32'hbe34298b, 32'hbd4744bc} /* (23, 5, 17) {real, imag} */,
  {32'h3db46ed0, 32'h3e9f71ca} /* (23, 5, 16) {real, imag} */,
  {32'hbd117420, 32'hbe099dbe} /* (23, 5, 15) {real, imag} */,
  {32'hbc8a9cc0, 32'hbda3d4dd} /* (23, 5, 14) {real, imag} */,
  {32'hbdac6413, 32'hbe397878} /* (23, 5, 13) {real, imag} */,
  {32'hbd9814bd, 32'h3ab827e0} /* (23, 5, 12) {real, imag} */,
  {32'hbeb41078, 32'hbf04a428} /* (23, 5, 11) {real, imag} */,
  {32'hbed18ac2, 32'hbc5c3ec0} /* (23, 5, 10) {real, imag} */,
  {32'hbaa25580, 32'hbdabb5bf} /* (23, 5, 9) {real, imag} */,
  {32'h3f46e1f5, 32'h3d3bcd28} /* (23, 5, 8) {real, imag} */,
  {32'h3b9a4540, 32'hbd370114} /* (23, 5, 7) {real, imag} */,
  {32'h3c6b3bc0, 32'h3eff234c} /* (23, 5, 6) {real, imag} */,
  {32'h3c9a0680, 32'hbf61f99c} /* (23, 5, 5) {real, imag} */,
  {32'h3e741b86, 32'h3fbd769c} /* (23, 5, 4) {real, imag} */,
  {32'h3e1f5de4, 32'hbf11ecb0} /* (23, 5, 3) {real, imag} */,
  {32'hbefae3ee, 32'hbf8f6100} /* (23, 5, 2) {real, imag} */,
  {32'h400039a0, 32'h4024d11e} /* (23, 5, 1) {real, imag} */,
  {32'h40179ddc, 32'h3f8a2077} /* (23, 5, 0) {real, imag} */,
  {32'hbfcc40d1, 32'hc0423c90} /* (23, 4, 31) {real, imag} */,
  {32'h403e3f20, 32'h4036ddde} /* (23, 4, 30) {real, imag} */,
  {32'h3e7356ad, 32'hbdc57254} /* (23, 4, 29) {real, imag} */,
  {32'hbfc33705, 32'hbef77f69} /* (23, 4, 28) {real, imag} */,
  {32'h3f512176, 32'hbf54c085} /* (23, 4, 27) {real, imag} */,
  {32'hbe142418, 32'hbe2e4926} /* (23, 4, 26) {real, imag} */,
  {32'hbece9410, 32'hbd8da686} /* (23, 4, 25) {real, imag} */,
  {32'h3fca805e, 32'h3e0fce1c} /* (23, 4, 24) {real, imag} */,
  {32'hbdb9c4ba, 32'hbbd00048} /* (23, 4, 23) {real, imag} */,
  {32'hbef1ffd4, 32'h3e827f1a} /* (23, 4, 22) {real, imag} */,
  {32'h3c442a58, 32'hbe8d2907} /* (23, 4, 21) {real, imag} */,
  {32'h3e8448f0, 32'h3ed5fba0} /* (23, 4, 20) {real, imag} */,
  {32'h3ee15fd6, 32'hbe4b687f} /* (23, 4, 19) {real, imag} */,
  {32'h3d56d6cc, 32'h3e95c101} /* (23, 4, 18) {real, imag} */,
  {32'h3ca57258, 32'hbeb4ff53} /* (23, 4, 17) {real, imag} */,
  {32'hbd97fd9a, 32'h3dd39c0b} /* (23, 4, 16) {real, imag} */,
  {32'h3eafde39, 32'hbe2dc509} /* (23, 4, 15) {real, imag} */,
  {32'h3c1399c8, 32'h3edb53d6} /* (23, 4, 14) {real, imag} */,
  {32'hbdb3f2ec, 32'h3e72c11e} /* (23, 4, 13) {real, imag} */,
  {32'hbdef15c8, 32'h3d14386c} /* (23, 4, 12) {real, imag} */,
  {32'hbee21ae0, 32'h3ec690a3} /* (23, 4, 11) {real, imag} */,
  {32'h3e7dbe28, 32'h3e8a49f0} /* (23, 4, 10) {real, imag} */,
  {32'hbe6f21ae, 32'hbeaf7851} /* (23, 4, 9) {real, imag} */,
  {32'h3e0b4bbe, 32'hbecc0111} /* (23, 4, 8) {real, imag} */,
  {32'hbf439506, 32'hbe849418} /* (23, 4, 7) {real, imag} */,
  {32'hbf1cb234, 32'h3e24a876} /* (23, 4, 6) {real, imag} */,
  {32'h3e8a241c, 32'h3da70af4} /* (23, 4, 5) {real, imag} */,
  {32'h3f86d6d6, 32'hbfa65bf0} /* (23, 4, 4) {real, imag} */,
  {32'h3ef02ed0, 32'hbf449130} /* (23, 4, 3) {real, imag} */,
  {32'h406c2057, 32'h3fe18a3b} /* (23, 4, 2) {real, imag} */,
  {32'hc084c3d7, 32'hbfef1274} /* (23, 4, 1) {real, imag} */,
  {32'hc01b529e, 32'h3f218e94} /* (23, 4, 0) {real, imag} */,
  {32'h4087fc76, 32'hc02ade2e} /* (23, 3, 31) {real, imag} */,
  {32'hc004e30c, 32'h404ca452} /* (23, 3, 30) {real, imag} */,
  {32'hbeeb201a, 32'h3ea2248a} /* (23, 3, 29) {real, imag} */,
  {32'hbf9632bb, 32'hbf538c60} /* (23, 3, 28) {real, imag} */,
  {32'h3fbe318e, 32'h3dc4c28c} /* (23, 3, 27) {real, imag} */,
  {32'hbea10dfb, 32'h3e3854ed} /* (23, 3, 26) {real, imag} */,
  {32'hbc51c5c0, 32'hbf7302c2} /* (23, 3, 25) {real, imag} */,
  {32'hbe7842c4, 32'h3ed18260} /* (23, 3, 24) {real, imag} */,
  {32'hbeba70ab, 32'hbee9f307} /* (23, 3, 23) {real, imag} */,
  {32'hbdc4a30c, 32'hbd8b2673} /* (23, 3, 22) {real, imag} */,
  {32'h3d734252, 32'hbe5d369b} /* (23, 3, 21) {real, imag} */,
  {32'hbe8803fc, 32'hbed798a4} /* (23, 3, 20) {real, imag} */,
  {32'hbe75e146, 32'h3eaf8656} /* (23, 3, 19) {real, imag} */,
  {32'h3e661327, 32'h3e42aa06} /* (23, 3, 18) {real, imag} */,
  {32'hbe9b4e51, 32'h3df626b0} /* (23, 3, 17) {real, imag} */,
  {32'h3f09be82, 32'h3d0e9e6c} /* (23, 3, 16) {real, imag} */,
  {32'h3e11f61f, 32'hbddaf65c} /* (23, 3, 15) {real, imag} */,
  {32'h3ceab118, 32'h3ea1dce6} /* (23, 3, 14) {real, imag} */,
  {32'h3dbbc1ae, 32'h3d89c567} /* (23, 3, 13) {real, imag} */,
  {32'hbf060867, 32'hbefbb03a} /* (23, 3, 12) {real, imag} */,
  {32'h3e9452f5, 32'hbe5fc04f} /* (23, 3, 11) {real, imag} */,
  {32'hbe328a51, 32'h3e6fe7f5} /* (23, 3, 10) {real, imag} */,
  {32'h3d847a64, 32'h3c170c38} /* (23, 3, 9) {real, imag} */,
  {32'hbe860738, 32'h3ee1a9de} /* (23, 3, 8) {real, imag} */,
  {32'hbeb5a23a, 32'hbf2fadc0} /* (23, 3, 7) {real, imag} */,
  {32'hbec75569, 32'h3f2ba4e3} /* (23, 3, 6) {real, imag} */,
  {32'hbeff5bf6, 32'hbf18e7ab} /* (23, 3, 5) {real, imag} */,
  {32'h3f99a45a, 32'hbf971346} /* (23, 3, 4) {real, imag} */,
  {32'hbe898167, 32'hbe72d87c} /* (23, 3, 3) {real, imag} */,
  {32'hbf0fba7a, 32'h4094b7e2} /* (23, 3, 2) {real, imag} */,
  {32'hc07a0378, 32'hc00b5b6e} /* (23, 3, 1) {real, imag} */,
  {32'h403289dc, 32'h3e8fab8d} /* (23, 3, 0) {real, imag} */,
  {32'h420d8d54, 32'h400929ed} /* (23, 2, 31) {real, imag} */,
  {32'hc1804dd6, 32'h4098de2e} /* (23, 2, 30) {real, imag} */,
  {32'h3f85622a, 32'hbf7e6136} /* (23, 2, 29) {real, imag} */,
  {32'h3f90b104, 32'hc026d48d} /* (23, 2, 28) {real, imag} */,
  {32'hbfef603e, 32'h3ef0b745} /* (23, 2, 27) {real, imag} */,
  {32'hbecdc896, 32'h3f2648f5} /* (23, 2, 26) {real, imag} */,
  {32'h3e1d8022, 32'h3e49aef5} /* (23, 2, 25) {real, imag} */,
  {32'hbe0e63de, 32'h3f075939} /* (23, 2, 24) {real, imag} */,
  {32'hbe92a177, 32'h3e6a2e14} /* (23, 2, 23) {real, imag} */,
  {32'h3dca5c8e, 32'h3e8e57a6} /* (23, 2, 22) {real, imag} */,
  {32'hbda19e03, 32'hbc9d9d76} /* (23, 2, 21) {real, imag} */,
  {32'h3e349ca0, 32'h3e835139} /* (23, 2, 20) {real, imag} */,
  {32'h3e681410, 32'h3e8996f8} /* (23, 2, 19) {real, imag} */,
  {32'h3cf7215d, 32'h3cc684e0} /* (23, 2, 18) {real, imag} */,
  {32'hbe96f083, 32'hbeca5172} /* (23, 2, 17) {real, imag} */,
  {32'hbe8054e7, 32'h3eccd86c} /* (23, 2, 16) {real, imag} */,
  {32'h3ecd39ba, 32'h3e840d6c} /* (23, 2, 15) {real, imag} */,
  {32'hbe5dafee, 32'hbd7c2230} /* (23, 2, 14) {real, imag} */,
  {32'hbe0d3392, 32'hbcc36538} /* (23, 2, 13) {real, imag} */,
  {32'hbe101495, 32'h3e03563e} /* (23, 2, 12) {real, imag} */,
  {32'hbea8cdde, 32'hbee9f938} /* (23, 2, 11) {real, imag} */,
  {32'h3df705b6, 32'h3ebf5da4} /* (23, 2, 10) {real, imag} */,
  {32'h3eb4e1ee, 32'h3ec9d1cb} /* (23, 2, 9) {real, imag} */,
  {32'hbf47eb87, 32'h3f40f53e} /* (23, 2, 8) {real, imag} */,
  {32'h3f12a0e2, 32'h3e98f4de} /* (23, 2, 7) {real, imag} */,
  {32'hbd5b9b90, 32'h3e14fb42} /* (23, 2, 6) {real, imag} */,
  {32'hc01969ca, 32'hc0095e65} /* (23, 2, 5) {real, imag} */,
  {32'h403ae243, 32'h3fef8566} /* (23, 2, 4) {real, imag} */,
  {32'h3e3051ae, 32'hbf84bbfa} /* (23, 2, 3) {real, imag} */,
  {32'hc13782d9, 32'h3fe039dd} /* (23, 2, 2) {real, imag} */,
  {32'h41a3b111, 32'hc00030bb} /* (23, 2, 1) {real, imag} */,
  {32'h41936f1d, 32'h405ebdb6} /* (23, 2, 0) {real, imag} */,
  {32'hc23ef642, 32'h41464375} /* (23, 1, 31) {real, imag} */,
  {32'h41397e08, 32'h4047a4af} /* (23, 1, 30) {real, imag} */,
  {32'h3fbed4c7, 32'hbf917ce6} /* (23, 1, 29) {real, imag} */,
  {32'hc07497c3, 32'hbf3b464a} /* (23, 1, 28) {real, imag} */,
  {32'h40835292, 32'hbe8a4b87} /* (23, 1, 27) {real, imag} */,
  {32'h3f000e6c, 32'h3e0ba27f} /* (23, 1, 26) {real, imag} */,
  {32'hbf08bbaa, 32'h3f32af03} /* (23, 1, 25) {real, imag} */,
  {32'h3ee4f898, 32'hbf18423e} /* (23, 1, 24) {real, imag} */,
  {32'h3e8b3e58, 32'hbf02ef78} /* (23, 1, 23) {real, imag} */,
  {32'hbeb5a73e, 32'hbbf46030} /* (23, 1, 22) {real, imag} */,
  {32'h3ed4f591, 32'hbe626385} /* (23, 1, 21) {real, imag} */,
  {32'hbdb680a9, 32'h3d271c0e} /* (23, 1, 20) {real, imag} */,
  {32'h3cc31cb4, 32'h3e2416b5} /* (23, 1, 19) {real, imag} */,
  {32'hbe95d8c3, 32'hbe81f154} /* (23, 1, 18) {real, imag} */,
  {32'h3da61db8, 32'hbecb530e} /* (23, 1, 17) {real, imag} */,
  {32'hbcc096e4, 32'h3d37c518} /* (23, 1, 16) {real, imag} */,
  {32'h3e157fdf, 32'hbdc5ed62} /* (23, 1, 15) {real, imag} */,
  {32'hbb7af530, 32'h3e711340} /* (23, 1, 14) {real, imag} */,
  {32'h3d412f58, 32'hbe9cd642} /* (23, 1, 13) {real, imag} */,
  {32'h3d9276c0, 32'hbd8b597a} /* (23, 1, 12) {real, imag} */,
  {32'hbe157f2a, 32'h3f49ef1c} /* (23, 1, 11) {real, imag} */,
  {32'h3e8a7593, 32'hbda5abe0} /* (23, 1, 10) {real, imag} */,
  {32'h3f22d8b8, 32'h3e560520} /* (23, 1, 9) {real, imag} */,
  {32'h3f08e354, 32'h3f047db0} /* (23, 1, 8) {real, imag} */,
  {32'hbf1b6a79, 32'hbef13484} /* (23, 1, 7) {real, imag} */,
  {32'h3f7a9161, 32'hbf1f313e} /* (23, 1, 6) {real, imag} */,
  {32'h4009667e, 32'h3fbc3ea8} /* (23, 1, 5) {real, imag} */,
  {32'hbff79290, 32'hbfce75d0} /* (23, 1, 4) {real, imag} */,
  {32'h3fe795ba, 32'h3f117c12} /* (23, 1, 3) {real, imag} */,
  {32'h4183b620, 32'h4174792e} /* (23, 1, 2) {real, imag} */,
  {32'hc2868bfc, 32'hc217fdc2} /* (23, 1, 1) {real, imag} */,
  {32'hc277c643, 32'hc0f49fae} /* (23, 1, 0) {real, imag} */,
  {32'hc2317406, 32'h420d2b08} /* (23, 0, 31) {real, imag} */,
  {32'h40b96d4a, 32'hc0dbc84f} /* (23, 0, 30) {real, imag} */,
  {32'h3eef21d6, 32'h3eb9f254} /* (23, 0, 29) {real, imag} */,
  {32'h3fcd64b2, 32'hc01f7024} /* (23, 0, 28) {real, imag} */,
  {32'h3fe8e6b6, 32'hbe08d3c1} /* (23, 0, 27) {real, imag} */,
  {32'h3e8d7894, 32'h3e66c979} /* (23, 0, 26) {real, imag} */,
  {32'h3f5dd128, 32'h3f0128b3} /* (23, 0, 25) {real, imag} */,
  {32'hbd8af342, 32'h3e1b05bc} /* (23, 0, 24) {real, imag} */,
  {32'h3ea3112e, 32'h3eadb5c9} /* (23, 0, 23) {real, imag} */,
  {32'hbf07c69d, 32'hbd9a0468} /* (23, 0, 22) {real, imag} */,
  {32'h3f045376, 32'h3ac5ec80} /* (23, 0, 21) {real, imag} */,
  {32'hbebdec88, 32'h3e4aa794} /* (23, 0, 20) {real, imag} */,
  {32'hbf136f7e, 32'hbd7e52d0} /* (23, 0, 19) {real, imag} */,
  {32'h3d3da822, 32'hbdedac72} /* (23, 0, 18) {real, imag} */,
  {32'h3d11129c, 32'h3d1982a4} /* (23, 0, 17) {real, imag} */,
  {32'hbe10722e, 32'h00000000} /* (23, 0, 16) {real, imag} */,
  {32'h3d11129c, 32'hbd1982a4} /* (23, 0, 15) {real, imag} */,
  {32'h3d3da822, 32'h3dedac72} /* (23, 0, 14) {real, imag} */,
  {32'hbf136f7e, 32'h3d7e52d0} /* (23, 0, 13) {real, imag} */,
  {32'hbebdec88, 32'hbe4aa794} /* (23, 0, 12) {real, imag} */,
  {32'h3f045376, 32'hbac5ec80} /* (23, 0, 11) {real, imag} */,
  {32'hbf07c69d, 32'h3d9a0468} /* (23, 0, 10) {real, imag} */,
  {32'h3ea3112e, 32'hbeadb5c9} /* (23, 0, 9) {real, imag} */,
  {32'hbd8af342, 32'hbe1b05bc} /* (23, 0, 8) {real, imag} */,
  {32'h3f5dd128, 32'hbf0128b3} /* (23, 0, 7) {real, imag} */,
  {32'h3e8d7894, 32'hbe66c979} /* (23, 0, 6) {real, imag} */,
  {32'h3fe8e6b6, 32'h3e08d3c1} /* (23, 0, 5) {real, imag} */,
  {32'h3fcd64b2, 32'h401f7024} /* (23, 0, 4) {real, imag} */,
  {32'h3eef21d6, 32'hbeb9f254} /* (23, 0, 3) {real, imag} */,
  {32'h40b96d4a, 32'h40dbc84f} /* (23, 0, 2) {real, imag} */,
  {32'hc2317406, 32'hc20d2b08} /* (23, 0, 1) {real, imag} */,
  {32'hc28b5d50, 32'h00000000} /* (23, 0, 0) {real, imag} */,
  {32'hc2988d2b, 32'h4223f327} /* (22, 31, 31) {real, imag} */,
  {32'h41900e9d, 32'hc18e30d7} /* (22, 31, 30) {real, imag} */,
  {32'h40056b01, 32'hbf410cc4} /* (22, 31, 29) {real, imag} */,
  {32'hbfd493e2, 32'h400f9744} /* (22, 31, 28) {real, imag} */,
  {32'h40087c97, 32'hbfe006c1} /* (22, 31, 27) {real, imag} */,
  {32'hbe01a2c4, 32'h3e4959ba} /* (22, 31, 26) {real, imag} */,
  {32'hbec586a9, 32'h3fadcd14} /* (22, 31, 25) {real, imag} */,
  {32'h3e19a629, 32'hbfbcd0a4} /* (22, 31, 24) {real, imag} */,
  {32'h3e4c8ed1, 32'h3ec5d99d} /* (22, 31, 23) {real, imag} */,
  {32'hbeb9412a, 32'hbecf3ee7} /* (22, 31, 22) {real, imag} */,
  {32'h3f03ab84, 32'hbe4cfb0d} /* (22, 31, 21) {real, imag} */,
  {32'h3e98f52a, 32'hbe10004c} /* (22, 31, 20) {real, imag} */,
  {32'hbeeed590, 32'h3e406d60} /* (22, 31, 19) {real, imag} */,
  {32'h3c543330, 32'hbee28776} /* (22, 31, 18) {real, imag} */,
  {32'hbe10964e, 32'hbea3f154} /* (22, 31, 17) {real, imag} */,
  {32'h3e2d62ce, 32'h3e18e40c} /* (22, 31, 16) {real, imag} */,
  {32'hbe0e4226, 32'hbdf2ac55} /* (22, 31, 15) {real, imag} */,
  {32'h3e1ab3ec, 32'hbe89683a} /* (22, 31, 14) {real, imag} */,
  {32'h3da08910, 32'h3e51ebb4} /* (22, 31, 13) {real, imag} */,
  {32'h3e4dcde5, 32'h3e5a1ffa} /* (22, 31, 12) {real, imag} */,
  {32'h3e7e650b, 32'hbe791436} /* (22, 31, 11) {real, imag} */,
  {32'h3eaeb0bd, 32'h3e8304c3} /* (22, 31, 10) {real, imag} */,
  {32'h3ef1c55c, 32'h3f4fefc6} /* (22, 31, 9) {real, imag} */,
  {32'h3ef9f2c4, 32'h3edd731e} /* (22, 31, 8) {real, imag} */,
  {32'hbf0ec39c, 32'h3ec895c4} /* (22, 31, 7) {real, imag} */,
  {32'h3f56bc25, 32'h3dd42674} /* (22, 31, 6) {real, imag} */,
  {32'h408f695e, 32'h3e9fe67f} /* (22, 31, 5) {real, imag} */,
  {32'hc08cdf8f, 32'h4002e392} /* (22, 31, 4) {real, imag} */,
  {32'h3f5c9d48, 32'h40092b77} /* (22, 31, 3) {real, imag} */,
  {32'h41649f0c, 32'hc02a096e} /* (22, 31, 2) {real, imag} */,
  {32'hc255cc2b, 32'hc1659299} /* (22, 31, 1) {real, imag} */,
  {32'hc286879a, 32'h41171b6c} /* (22, 31, 0) {real, imag} */,
  {32'h41b39153, 32'h40262180} /* (22, 30, 31) {real, imag} */,
  {32'hc14d8aca, 32'hc0361d12} /* (22, 30, 30) {real, imag} */,
  {32'h3e26fc6c, 32'h3fb6204b} /* (22, 30, 29) {real, imag} */,
  {32'h40403adf, 32'hc00b6ee7} /* (22, 30, 28) {real, imag} */,
  {32'hc0234c60, 32'h40103032} /* (22, 30, 27) {real, imag} */,
  {32'hbe62859a, 32'hbedce178} /* (22, 30, 26) {real, imag} */,
  {32'h3cdf1538, 32'h3dc9f334} /* (22, 30, 25) {real, imag} */,
  {32'hbf2b67ca, 32'h3f105571} /* (22, 30, 24) {real, imag} */,
  {32'h3e09fac1, 32'h3d48fcfc} /* (22, 30, 23) {real, imag} */,
  {32'h3ed9f63e, 32'hbf3283f3} /* (22, 30, 22) {real, imag} */,
  {32'hbe12b6b3, 32'h3f296855} /* (22, 30, 21) {real, imag} */,
  {32'hbedb1b2a, 32'h3f07bac5} /* (22, 30, 20) {real, imag} */,
  {32'h3ebd8a8e, 32'hbe3a691a} /* (22, 30, 19) {real, imag} */,
  {32'h3edc3672, 32'hbd9cd974} /* (22, 30, 18) {real, imag} */,
  {32'hbd1b4978, 32'hbdb2ef32} /* (22, 30, 17) {real, imag} */,
  {32'h3d216b7e, 32'h3c01b444} /* (22, 30, 16) {real, imag} */,
  {32'h37368000, 32'h3e5d188a} /* (22, 30, 15) {real, imag} */,
  {32'hbdd2c0c6, 32'hbedf3a92} /* (22, 30, 14) {real, imag} */,
  {32'hbf126ad2, 32'hbee30a28} /* (22, 30, 13) {real, imag} */,
  {32'h3ea646c0, 32'hbea78714} /* (22, 30, 12) {real, imag} */,
  {32'h3d7429b4, 32'hbe906ed8} /* (22, 30, 11) {real, imag} */,
  {32'hbdde7c60, 32'hbeacb5f8} /* (22, 30, 10) {real, imag} */,
  {32'hbe886ef7, 32'h3e858c64} /* (22, 30, 9) {real, imag} */,
  {32'hbeabd461, 32'hbe8ba84c} /* (22, 30, 8) {real, imag} */,
  {32'h3f623c04, 32'h3ee20bc2} /* (22, 30, 7) {real, imag} */,
  {32'hbf9428ad, 32'h3e343f0c} /* (22, 30, 6) {real, imag} */,
  {32'hbfde244b, 32'hbf69443b} /* (22, 30, 5) {real, imag} */,
  {32'h3f8fa701, 32'h40443e52} /* (22, 30, 4) {real, imag} */,
  {32'hbe05e878, 32'h3f31d48c} /* (22, 30, 3) {real, imag} */,
  {32'hc18ac138, 32'hc0d04f88} /* (22, 30, 2) {real, imag} */,
  {32'h421cedcb, 32'hbf999956} /* (22, 30, 1) {real, imag} */,
  {32'h419f47b8, 32'hc089dc98} /* (22, 30, 0) {real, imag} */,
  {32'hc084234c, 32'h402bcd6e} /* (22, 29, 31) {real, imag} */,
  {32'hbf0e3b76, 32'hc08959f0} /* (22, 29, 30) {real, imag} */,
  {32'h3db09af0, 32'h3f26b081} /* (22, 29, 29) {real, imag} */,
  {32'h3f5c5fce, 32'h3ff481d2} /* (22, 29, 28) {real, imag} */,
  {32'hbf3d52a3, 32'h3e61d01e} /* (22, 29, 27) {real, imag} */,
  {32'h3ef16600, 32'hbdc16bda} /* (22, 29, 26) {real, imag} */,
  {32'h3e6f066d, 32'h3e80565c} /* (22, 29, 25) {real, imag} */,
  {32'hbed8a89a, 32'hbef847e9} /* (22, 29, 24) {real, imag} */,
  {32'hbeac692c, 32'h3f0d3c98} /* (22, 29, 23) {real, imag} */,
  {32'hbe98ca58, 32'hbf2b1016} /* (22, 29, 22) {real, imag} */,
  {32'hbe8190a6, 32'hbd60d310} /* (22, 29, 21) {real, imag} */,
  {32'h3f20bde2, 32'h3e158254} /* (22, 29, 20) {real, imag} */,
  {32'h3dd60d7b, 32'hbea3a702} /* (22, 29, 19) {real, imag} */,
  {32'hbea88d5a, 32'hbd56ae3c} /* (22, 29, 18) {real, imag} */,
  {32'hbead7de3, 32'h3d795bc0} /* (22, 29, 17) {real, imag} */,
  {32'h3e252e0e, 32'h3e3c638a} /* (22, 29, 16) {real, imag} */,
  {32'hbe3893e3, 32'hbe124c06} /* (22, 29, 15) {real, imag} */,
  {32'h3ec84e6e, 32'hbdaa3cf0} /* (22, 29, 14) {real, imag} */,
  {32'h3e9e469c, 32'hbe97baa7} /* (22, 29, 13) {real, imag} */,
  {32'h3eacb868, 32'h3ea4bee4} /* (22, 29, 12) {real, imag} */,
  {32'hbbfd4e98, 32'hbe5f7e68} /* (22, 29, 11) {real, imag} */,
  {32'hbec0f862, 32'h3eb9b9e8} /* (22, 29, 10) {real, imag} */,
  {32'hbdf14d3c, 32'h3ef7f472} /* (22, 29, 9) {real, imag} */,
  {32'h3f494744, 32'hbe434ee3} /* (22, 29, 8) {real, imag} */,
  {32'h3e931b8f, 32'h3f19069b} /* (22, 29, 7) {real, imag} */,
  {32'h3e13ddb4, 32'h3e0605e2} /* (22, 29, 6) {real, imag} */,
  {32'h3f299642, 32'hbe7385f4} /* (22, 29, 5) {real, imag} */,
  {32'hbfeafca8, 32'h3f7a9d50} /* (22, 29, 4) {real, imag} */,
  {32'hbda16f84, 32'h3e0ddfa6} /* (22, 29, 3) {real, imag} */,
  {32'hc03e7f5b, 32'hc05b40fa} /* (22, 29, 2) {real, imag} */,
  {32'h40928d49, 32'h400e305d} /* (22, 29, 1) {real, imag} */,
  {32'h40050126, 32'h3c845a60} /* (22, 29, 0) {real, imag} */,
  {32'hc068461e, 32'h3f94eb4a} /* (22, 28, 31) {real, imag} */,
  {32'h4059f190, 32'hc004598b} /* (22, 28, 30) {real, imag} */,
  {32'h3ea73f7a, 32'h3e87b3df} /* (22, 28, 29) {real, imag} */,
  {32'h3f0fd021, 32'h3f9d48d5} /* (22, 28, 28) {real, imag} */,
  {32'h3daf07ec, 32'hbd8149b0} /* (22, 28, 27) {real, imag} */,
  {32'hbef1bdc2, 32'h3db0a72c} /* (22, 28, 26) {real, imag} */,
  {32'hbe1adeb2, 32'h3c5728f0} /* (22, 28, 25) {real, imag} */,
  {32'h3f0529ee, 32'h3e2c7a72} /* (22, 28, 24) {real, imag} */,
  {32'h3e6cd5c7, 32'h3e4956e1} /* (22, 28, 23) {real, imag} */,
  {32'hbcd12900, 32'hbefdd395} /* (22, 28, 22) {real, imag} */,
  {32'h3eb88ff7, 32'hbef30493} /* (22, 28, 21) {real, imag} */,
  {32'hbe462c98, 32'h3f1dd60a} /* (22, 28, 20) {real, imag} */,
  {32'hbe7d0c50, 32'hbe4b30e0} /* (22, 28, 19) {real, imag} */,
  {32'h3ece3398, 32'hbde42fb5} /* (22, 28, 18) {real, imag} */,
  {32'hbe0239bd, 32'hbda717d0} /* (22, 28, 17) {real, imag} */,
  {32'hbdf0b3f8, 32'hbd999a83} /* (22, 28, 16) {real, imag} */,
  {32'hbb212eb8, 32'h3c9a0f30} /* (22, 28, 15) {real, imag} */,
  {32'h3ef568e6, 32'h3e79c769} /* (22, 28, 14) {real, imag} */,
  {32'hbca40991, 32'hbddc9c43} /* (22, 28, 13) {real, imag} */,
  {32'h3cf9ade8, 32'h3ddf8728} /* (22, 28, 12) {real, imag} */,
  {32'hbea99460, 32'hbeb26464} /* (22, 28, 11) {real, imag} */,
  {32'hbe056abc, 32'hbe3277ee} /* (22, 28, 10) {real, imag} */,
  {32'hbe99c65e, 32'h3eead1b3} /* (22, 28, 9) {real, imag} */,
  {32'h3f142800, 32'hbed4c1ee} /* (22, 28, 8) {real, imag} */,
  {32'h3e9272a0, 32'h3e24770b} /* (22, 28, 7) {real, imag} */,
  {32'h3e1b4b7e, 32'h3ea30b76} /* (22, 28, 6) {real, imag} */,
  {32'h3ecc0331, 32'h3ebe7112} /* (22, 28, 5) {real, imag} */,
  {32'hbf27e602, 32'h3e431b48} /* (22, 28, 4) {real, imag} */,
  {32'hbf56fa5a, 32'hbe4f89b1} /* (22, 28, 3) {real, imag} */,
  {32'h402cce27, 32'hc0258a7e} /* (22, 28, 2) {real, imag} */,
  {32'hbf8ac486, 32'h404aa144} /* (22, 28, 1) {real, imag} */,
  {32'hc02687b2, 32'hbf523d72} /* (22, 28, 0) {real, imag} */,
  {32'h4043ee42, 32'hc03cd575} /* (22, 27, 31) {real, imag} */,
  {32'h3e577095, 32'h3fa206a0} /* (22, 27, 30) {real, imag} */,
  {32'hbda7484b, 32'h3e2225be} /* (22, 27, 29) {real, imag} */,
  {32'hbea60f44, 32'hbfbf19b2} /* (22, 27, 28) {real, imag} */,
  {32'hbe98e420, 32'h3f3a9662} /* (22, 27, 27) {real, imag} */,
  {32'h3ec3ae9a, 32'hbd89e92a} /* (22, 27, 26) {real, imag} */,
  {32'h3e9ca0d2, 32'h3d15b224} /* (22, 27, 25) {real, imag} */,
  {32'hbd348140, 32'h3bd47800} /* (22, 27, 24) {real, imag} */,
  {32'h3e45c1b3, 32'h3c2eb738} /* (22, 27, 23) {real, imag} */,
  {32'hbe291a7e, 32'h3eb4a42a} /* (22, 27, 22) {real, imag} */,
  {32'hbe2da160, 32'h3f016d7c} /* (22, 27, 21) {real, imag} */,
  {32'hbed6c29c, 32'h3e58ed0f} /* (22, 27, 20) {real, imag} */,
  {32'h3ece23aa, 32'h3e2b34ff} /* (22, 27, 19) {real, imag} */,
  {32'h3eb1207a, 32'h3e404c78} /* (22, 27, 18) {real, imag} */,
  {32'hbd9ba87c, 32'hbe4240c8} /* (22, 27, 17) {real, imag} */,
  {32'hbeea741c, 32'h3e943956} /* (22, 27, 16) {real, imag} */,
  {32'h3d4bfbe1, 32'h3daad196} /* (22, 27, 15) {real, imag} */,
  {32'h3ec05570, 32'hbc010700} /* (22, 27, 14) {real, imag} */,
  {32'h3e345590, 32'h3e277a51} /* (22, 27, 13) {real, imag} */,
  {32'h3e863ef1, 32'h3f012952} /* (22, 27, 12) {real, imag} */,
  {32'hbda1cc62, 32'hbd771508} /* (22, 27, 11) {real, imag} */,
  {32'hbf2aa39b, 32'hbe6bd3de} /* (22, 27, 10) {real, imag} */,
  {32'h3e894d30, 32'h3f0040d8} /* (22, 27, 9) {real, imag} */,
  {32'hbec9f456, 32'hbd5bddd0} /* (22, 27, 8) {real, imag} */,
  {32'hbe39983c, 32'h3e4ead34} /* (22, 27, 7) {real, imag} */,
  {32'hbd53cf8a, 32'hbf348a86} /* (22, 27, 6) {real, imag} */,
  {32'hbf981e7b, 32'h3dca6d3a} /* (22, 27, 5) {real, imag} */,
  {32'hbef7b875, 32'h3df0f3e8} /* (22, 27, 4) {real, imag} */,
  {32'hbd921dbf, 32'h3e332cc4} /* (22, 27, 3) {real, imag} */,
  {32'hbff955d3, 32'h3ef0a908} /* (22, 27, 2) {real, imag} */,
  {32'h40421804, 32'hbf4d22ba} /* (22, 27, 1) {real, imag} */,
  {32'h400e3266, 32'hbfa1a283} /* (22, 27, 0) {real, imag} */,
  {32'h3ec6bbf4, 32'hbe59f576} /* (22, 26, 31) {real, imag} */,
  {32'hbf1c8e86, 32'hbdb8636c} /* (22, 26, 30) {real, imag} */,
  {32'h3f3e9294, 32'h3f8208b2} /* (22, 26, 29) {real, imag} */,
  {32'h3e845c35, 32'hbd2dbb34} /* (22, 26, 28) {real, imag} */,
  {32'hbf48a185, 32'hbe7bd728} /* (22, 26, 27) {real, imag} */,
  {32'hbe285a07, 32'h3f023415} /* (22, 26, 26) {real, imag} */,
  {32'hbef03075, 32'h3e735a2e} /* (22, 26, 25) {real, imag} */,
  {32'h3e348b03, 32'h3e9f0ce4} /* (22, 26, 24) {real, imag} */,
  {32'h3e0b95f7, 32'h3dacae22} /* (22, 26, 23) {real, imag} */,
  {32'hbf1c00b5, 32'hbcc3dbf0} /* (22, 26, 22) {real, imag} */,
  {32'hbea37747, 32'hbe4a14f6} /* (22, 26, 21) {real, imag} */,
  {32'h3e8f0d5f, 32'hbeeb3741} /* (22, 26, 20) {real, imag} */,
  {32'h3e88d128, 32'hbd96f279} /* (22, 26, 19) {real, imag} */,
  {32'hbe7934d4, 32'hbea1719e} /* (22, 26, 18) {real, imag} */,
  {32'hbe3d2b0a, 32'hbe62332f} /* (22, 26, 17) {real, imag} */,
  {32'hbe1e9fb3, 32'hbda735e0} /* (22, 26, 16) {real, imag} */,
  {32'h3d389124, 32'h3e70202a} /* (22, 26, 15) {real, imag} */,
  {32'hbdaa1d7a, 32'hbe1ca880} /* (22, 26, 14) {real, imag} */,
  {32'hbd8ff1e4, 32'hbec6abe1} /* (22, 26, 13) {real, imag} */,
  {32'hbe031127, 32'h3e761efd} /* (22, 26, 12) {real, imag} */,
  {32'hbc8a1560, 32'h3e4fb4f0} /* (22, 26, 11) {real, imag} */,
  {32'hbe1d2bd2, 32'hbf00d7e6} /* (22, 26, 10) {real, imag} */,
  {32'hbedec086, 32'hbdc27e68} /* (22, 26, 9) {real, imag} */,
  {32'h3e827f05, 32'h3ee3b4f2} /* (22, 26, 8) {real, imag} */,
  {32'hbe8cae06, 32'h3c558d18} /* (22, 26, 7) {real, imag} */,
  {32'hbf155776, 32'hbe845686} /* (22, 26, 6) {real, imag} */,
  {32'hbdd5aec8, 32'h3e3d3122} /* (22, 26, 5) {real, imag} */,
  {32'hbd8926ec, 32'h3f2c5217} /* (22, 26, 4) {real, imag} */,
  {32'h3e5784e1, 32'hbedbcf7c} /* (22, 26, 3) {real, imag} */,
  {32'hbe5aba98, 32'h3e5e9f77} /* (22, 26, 2) {real, imag} */,
  {32'h3e9730e6, 32'hbe70ccd4} /* (22, 26, 1) {real, imag} */,
  {32'h3cd057f0, 32'hbeae6960} /* (22, 26, 0) {real, imag} */,
  {32'hbdfe6088, 32'h3f1a0693} /* (22, 25, 31) {real, imag} */,
  {32'hbe98243d, 32'h3e923a1f} /* (22, 25, 30) {real, imag} */,
  {32'h3eba04ed, 32'hbf97fc00} /* (22, 25, 29) {real, imag} */,
  {32'h3cd47e88, 32'h3ed56654} /* (22, 25, 28) {real, imag} */,
  {32'h3e1be992, 32'hbe8778ad} /* (22, 25, 27) {real, imag} */,
  {32'h3e8207e4, 32'hbe2dbc15} /* (22, 25, 26) {real, imag} */,
  {32'hbe23cd84, 32'h3f7b595c} /* (22, 25, 25) {real, imag} */,
  {32'h3e469615, 32'h3eda709b} /* (22, 25, 24) {real, imag} */,
  {32'hbdd8415e, 32'h3d284cfc} /* (22, 25, 23) {real, imag} */,
  {32'hbea41624, 32'hbea44048} /* (22, 25, 22) {real, imag} */,
  {32'hbf412ec4, 32'hbcf9bcb8} /* (22, 25, 21) {real, imag} */,
  {32'hbe0dfb04, 32'hbe62de5c} /* (22, 25, 20) {real, imag} */,
  {32'h3dbf3eb6, 32'hbdb9a450} /* (22, 25, 19) {real, imag} */,
  {32'hbe531a67, 32'hbb82df40} /* (22, 25, 18) {real, imag} */,
  {32'h3d3da130, 32'hbe8cc1ed} /* (22, 25, 17) {real, imag} */,
  {32'h3e09a110, 32'hbe2fb7e3} /* (22, 25, 16) {real, imag} */,
  {32'h3e8df84d, 32'h3e653efa} /* (22, 25, 15) {real, imag} */,
  {32'h3e8a371e, 32'h3d5a6f24} /* (22, 25, 14) {real, imag} */,
  {32'hbeff67d8, 32'hbe6a6ede} /* (22, 25, 13) {real, imag} */,
  {32'h3d1dd128, 32'h3f0737ad} /* (22, 25, 12) {real, imag} */,
  {32'h3ed25f6f, 32'h3d322162} /* (22, 25, 11) {real, imag} */,
  {32'hbe733b7f, 32'h3dca8c68} /* (22, 25, 10) {real, imag} */,
  {32'h3eecc39c, 32'hbe9bb4c1} /* (22, 25, 9) {real, imag} */,
  {32'hbf7ede80, 32'hbdd8fada} /* (22, 25, 8) {real, imag} */,
  {32'h3e351048, 32'hbc5960d0} /* (22, 25, 7) {real, imag} */,
  {32'hbeb23ec0, 32'hbec8946c} /* (22, 25, 6) {real, imag} */,
  {32'hbd8dff9c, 32'hbdd11860} /* (22, 25, 5) {real, imag} */,
  {32'h3f18ee7e, 32'hbec4ac83} /* (22, 25, 4) {real, imag} */,
  {32'h3f2ccc00, 32'hbe6c65aa} /* (22, 25, 3) {real, imag} */,
  {32'h3e938f8e, 32'hbdccb8a4} /* (22, 25, 2) {real, imag} */,
  {32'hbf2b9732, 32'h3f194f12} /* (22, 25, 1) {real, imag} */,
  {32'hbe1c0135, 32'h3f086aca} /* (22, 25, 0) {real, imag} */,
  {32'h3d309408, 32'hbe80b8d0} /* (22, 24, 31) {real, imag} */,
  {32'hbe0acbbc, 32'hbdb25fbc} /* (22, 24, 30) {real, imag} */,
  {32'h3d175e78, 32'h3ec1ca30} /* (22, 24, 29) {real, imag} */,
  {32'h3ee855cc, 32'hbf174d68} /* (22, 24, 28) {real, imag} */,
  {32'hbf43f168, 32'h3e94d480} /* (22, 24, 27) {real, imag} */,
  {32'h3d8450a6, 32'hbdc45bfa} /* (22, 24, 26) {real, imag} */,
  {32'h3f08fee8, 32'h3e958c42} /* (22, 24, 25) {real, imag} */,
  {32'hbed614ca, 32'h3ece72d1} /* (22, 24, 24) {real, imag} */,
  {32'hbce01f88, 32'hbe9013b2} /* (22, 24, 23) {real, imag} */,
  {32'hbd059606, 32'hbf0c7c12} /* (22, 24, 22) {real, imag} */,
  {32'h3f282a69, 32'h3e489583} /* (22, 24, 21) {real, imag} */,
  {32'hbeb9c91a, 32'hbcc4632c} /* (22, 24, 20) {real, imag} */,
  {32'hbec99845, 32'h3e923204} /* (22, 24, 19) {real, imag} */,
  {32'h3e3c1594, 32'h3f05fac3} /* (22, 24, 18) {real, imag} */,
  {32'hbd74420c, 32'hbd28dc81} /* (22, 24, 17) {real, imag} */,
  {32'hbeda6224, 32'hbd82520a} /* (22, 24, 16) {real, imag} */,
  {32'hbbb0d948, 32'h3db51b24} /* (22, 24, 15) {real, imag} */,
  {32'hbdf5c764, 32'h3e5db011} /* (22, 24, 14) {real, imag} */,
  {32'hbea76f60, 32'h3e65f2ac} /* (22, 24, 13) {real, imag} */,
  {32'hbe317df2, 32'hbdd72944} /* (22, 24, 12) {real, imag} */,
  {32'hbe6f5480, 32'hbeb44aa6} /* (22, 24, 11) {real, imag} */,
  {32'hbed1c784, 32'h3e988649} /* (22, 24, 10) {real, imag} */,
  {32'h3ed59cda, 32'hbd1fd8fa} /* (22, 24, 9) {real, imag} */,
  {32'hbe648a0e, 32'h3e959480} /* (22, 24, 8) {real, imag} */,
  {32'h3e988029, 32'hbf23d7ea} /* (22, 24, 7) {real, imag} */,
  {32'h3cc58ecc, 32'h3e0f167a} /* (22, 24, 6) {real, imag} */,
  {32'hbf7767f4, 32'h3e7d2656} /* (22, 24, 5) {real, imag} */,
  {32'h3e4234ba, 32'h3e96adec} /* (22, 24, 4) {real, imag} */,
  {32'hbbd8e480, 32'hbeaa1da8} /* (22, 24, 3) {real, imag} */,
  {32'hbf265f70, 32'h3de2ef98} /* (22, 24, 2) {real, imag} */,
  {32'h3fa1e523, 32'hbf2ccf87} /* (22, 24, 1) {real, imag} */,
  {32'h3f4836bc, 32'h3cce39f0} /* (22, 24, 0) {real, imag} */,
  {32'hbeb668f0, 32'h3f341f1c} /* (22, 23, 31) {real, imag} */,
  {32'h3e5ea2d2, 32'hbe726056} /* (22, 23, 30) {real, imag} */,
  {32'h3e5be485, 32'hbf3a0f44} /* (22, 23, 29) {real, imag} */,
  {32'h3eeceb87, 32'h3dad917e} /* (22, 23, 28) {real, imag} */,
  {32'hbd163938, 32'h3c457f20} /* (22, 23, 27) {real, imag} */,
  {32'hbf5bf7b6, 32'h3e79aab9} /* (22, 23, 26) {real, imag} */,
  {32'h3ef88d0a, 32'hbd007fa8} /* (22, 23, 25) {real, imag} */,
  {32'h3f0d77de, 32'hbf1e6f9a} /* (22, 23, 24) {real, imag} */,
  {32'h3f14c7b8, 32'h3f11d592} /* (22, 23, 23) {real, imag} */,
  {32'hbdbe2834, 32'hbe5a4ff6} /* (22, 23, 22) {real, imag} */,
  {32'h3ded52fa, 32'hbce9c8f8} /* (22, 23, 21) {real, imag} */,
  {32'h3e846a88, 32'h3f03578a} /* (22, 23, 20) {real, imag} */,
  {32'hbee8021e, 32'hbd53443c} /* (22, 23, 19) {real, imag} */,
  {32'h3c836740, 32'h3e94e742} /* (22, 23, 18) {real, imag} */,
  {32'h3f16e4d8, 32'hbcfe2078} /* (22, 23, 17) {real, imag} */,
  {32'hbdf4b04e, 32'hbd1cc73a} /* (22, 23, 16) {real, imag} */,
  {32'hbe19be2f, 32'hbeb4fd80} /* (22, 23, 15) {real, imag} */,
  {32'hbdce4362, 32'hbe567db9} /* (22, 23, 14) {real, imag} */,
  {32'h3da17952, 32'h3ecb4666} /* (22, 23, 13) {real, imag} */,
  {32'h3e2544ea, 32'hbdf6113c} /* (22, 23, 12) {real, imag} */,
  {32'hbe850f30, 32'hbe2b1c36} /* (22, 23, 11) {real, imag} */,
  {32'h3e8717e4, 32'hbf12538c} /* (22, 23, 10) {real, imag} */,
  {32'hbe0c2066, 32'h3dbf9dd8} /* (22, 23, 9) {real, imag} */,
  {32'h3e83cfa6, 32'h3df4f100} /* (22, 23, 8) {real, imag} */,
  {32'hbec7a8e8, 32'h3f02cae7} /* (22, 23, 7) {real, imag} */,
  {32'hbeb526f1, 32'hbe8a7080} /* (22, 23, 6) {real, imag} */,
  {32'h3edd8f46, 32'hbcd4d198} /* (22, 23, 5) {real, imag} */,
  {32'h3cc4a8c0, 32'hbf69db56} /* (22, 23, 4) {real, imag} */,
  {32'h3afa0bc0, 32'h3e5a0497} /* (22, 23, 3) {real, imag} */,
  {32'h3eb617ae, 32'hbf26955a} /* (22, 23, 2) {real, imag} */,
  {32'h3ee0f5a0, 32'h3e771154} /* (22, 23, 1) {real, imag} */,
  {32'h3a44c380, 32'hbf0778a3} /* (22, 23, 0) {real, imag} */,
  {32'hbef5f9f3, 32'h3f26a64c} /* (22, 22, 31) {real, imag} */,
  {32'h3dcd29c4, 32'hbf20ae24} /* (22, 22, 30) {real, imag} */,
  {32'h3eb9e037, 32'h3ed1bce4} /* (22, 22, 29) {real, imag} */,
  {32'h3d6e6e53, 32'h3e5b33ef} /* (22, 22, 28) {real, imag} */,
  {32'hbeb3cdb6, 32'hbee6d7e3} /* (22, 22, 27) {real, imag} */,
  {32'h3c3146a0, 32'hbf063872} /* (22, 22, 26) {real, imag} */,
  {32'hbe23abc2, 32'h3e57ceb0} /* (22, 22, 25) {real, imag} */,
  {32'hbe3ae46b, 32'hbe17de57} /* (22, 22, 24) {real, imag} */,
  {32'hbe04a6f4, 32'hbe82639c} /* (22, 22, 23) {real, imag} */,
  {32'hbf1b12a4, 32'hbd7c0af0} /* (22, 22, 22) {real, imag} */,
  {32'hbe92c0aa, 32'h3e43c5e1} /* (22, 22, 21) {real, imag} */,
  {32'hbe652cec, 32'h3eb0e0db} /* (22, 22, 20) {real, imag} */,
  {32'h3eb9aa2b, 32'hbf19c92d} /* (22, 22, 19) {real, imag} */,
  {32'hbd403668, 32'hbaecd400} /* (22, 22, 18) {real, imag} */,
  {32'h3c979c48, 32'h3e28a8a4} /* (22, 22, 17) {real, imag} */,
  {32'hbd98b262, 32'h3d93c91f} /* (22, 22, 16) {real, imag} */,
  {32'hbe847320, 32'h3d7136c2} /* (22, 22, 15) {real, imag} */,
  {32'h3d82ef9a, 32'hbe83d3db} /* (22, 22, 14) {real, imag} */,
  {32'hbe3d6bb0, 32'hbbe26800} /* (22, 22, 13) {real, imag} */,
  {32'h3f409cb0, 32'hbd9956f0} /* (22, 22, 12) {real, imag} */,
  {32'hbe9ffd89, 32'h3e32bc9e} /* (22, 22, 11) {real, imag} */,
  {32'h3e014a0c, 32'h3ebc4d40} /* (22, 22, 10) {real, imag} */,
  {32'hbd5300a0, 32'hbd2c69a0} /* (22, 22, 9) {real, imag} */,
  {32'h3ea85826, 32'h3b107600} /* (22, 22, 8) {real, imag} */,
  {32'hbe436150, 32'h3df7c867} /* (22, 22, 7) {real, imag} */,
  {32'hbde0b63e, 32'h3dd9f8fc} /* (22, 22, 6) {real, imag} */,
  {32'h3d708c98, 32'h3f031928} /* (22, 22, 5) {real, imag} */,
  {32'hbea44114, 32'h3eb32a8a} /* (22, 22, 4) {real, imag} */,
  {32'hbdb28002, 32'h3f2cd678} /* (22, 22, 3) {real, imag} */,
  {32'hbe868551, 32'hbe43a112} /* (22, 22, 2) {real, imag} */,
  {32'h3d9e6ff8, 32'h3efa19cb} /* (22, 22, 1) {real, imag} */,
  {32'hbd184f34, 32'h3ed5420c} /* (22, 22, 0) {real, imag} */,
  {32'hbd1a2989, 32'hbf624284} /* (22, 21, 31) {real, imag} */,
  {32'h3d5c9170, 32'h3de5075c} /* (22, 21, 30) {real, imag} */,
  {32'hbda07cf0, 32'h3e30bf5f} /* (22, 21, 29) {real, imag} */,
  {32'h3e846f58, 32'hbf190675} /* (22, 21, 28) {real, imag} */,
  {32'hbed951da, 32'hbef686e0} /* (22, 21, 27) {real, imag} */,
  {32'hbf555511, 32'hbe37e8a2} /* (22, 21, 26) {real, imag} */,
  {32'hbde2cce0, 32'h3e1dc849} /* (22, 21, 25) {real, imag} */,
  {32'hbdb36229, 32'h3e9e395e} /* (22, 21, 24) {real, imag} */,
  {32'hbe09ca3e, 32'hbf85e66c} /* (22, 21, 23) {real, imag} */,
  {32'hbd756f12, 32'hbe28c722} /* (22, 21, 22) {real, imag} */,
  {32'hbf078182, 32'h3e098eb0} /* (22, 21, 21) {real, imag} */,
  {32'h3eadb0d6, 32'hbf30bc9a} /* (22, 21, 20) {real, imag} */,
  {32'hbe72b125, 32'hbedbb445} /* (22, 21, 19) {real, imag} */,
  {32'h3e4881dd, 32'hbe41d402} /* (22, 21, 18) {real, imag} */,
  {32'hbd56a005, 32'h3c5bad90} /* (22, 21, 17) {real, imag} */,
  {32'hbc4119d0, 32'hbe5ca602} /* (22, 21, 16) {real, imag} */,
  {32'h3e9f54d3, 32'h3db3f33e} /* (22, 21, 15) {real, imag} */,
  {32'hbe9df448, 32'hbecf0619} /* (22, 21, 14) {real, imag} */,
  {32'h3dbcd7b1, 32'h3c8a09f8} /* (22, 21, 13) {real, imag} */,
  {32'h3e58c2f0, 32'hbcdf94f8} /* (22, 21, 12) {real, imag} */,
  {32'hbe378b1d, 32'h3e086bf8} /* (22, 21, 11) {real, imag} */,
  {32'hbf2eded1, 32'h3daa374c} /* (22, 21, 10) {real, imag} */,
  {32'hbedc7b3b, 32'hbf0aaa5a} /* (22, 21, 9) {real, imag} */,
  {32'h3e845016, 32'hbd23fe18} /* (22, 21, 8) {real, imag} */,
  {32'hbe35202e, 32'hbf14c302} /* (22, 21, 7) {real, imag} */,
  {32'h3c769840, 32'hbea47110} /* (22, 21, 6) {real, imag} */,
  {32'hbcc8fa24, 32'h3f1ed968} /* (22, 21, 5) {real, imag} */,
  {32'hbe59efb1, 32'h3e0aa936} /* (22, 21, 4) {real, imag} */,
  {32'h3e0ed08e, 32'h3d6e7294} /* (22, 21, 3) {real, imag} */,
  {32'hbe4746e0, 32'h3f44c023} /* (22, 21, 2) {real, imag} */,
  {32'h3e803910, 32'hbe90caa4} /* (22, 21, 1) {real, imag} */,
  {32'h3e5a7052, 32'hbebe6be2} /* (22, 21, 0) {real, imag} */,
  {32'hbcbf298e, 32'hbda31ea6} /* (22, 20, 31) {real, imag} */,
  {32'h3e3aa854, 32'h3e18a69a} /* (22, 20, 30) {real, imag} */,
  {32'hbad2b340, 32'h3e80f2cc} /* (22, 20, 29) {real, imag} */,
  {32'h3d946c24, 32'h3e0905b5} /* (22, 20, 28) {real, imag} */,
  {32'h3e5b55b6, 32'hbf47d110} /* (22, 20, 27) {real, imag} */,
  {32'h3e10c3e9, 32'h3d8b20bb} /* (22, 20, 26) {real, imag} */,
  {32'hbe4a6606, 32'hbe9005a0} /* (22, 20, 25) {real, imag} */,
  {32'hbe6120ba, 32'hbea137f2} /* (22, 20, 24) {real, imag} */,
  {32'h3ebbdccc, 32'h3c35eb60} /* (22, 20, 23) {real, imag} */,
  {32'h3e9349cc, 32'hbd269958} /* (22, 20, 22) {real, imag} */,
  {32'h3dd847ee, 32'hbe7963ff} /* (22, 20, 21) {real, imag} */,
  {32'h3ee59c80, 32'h3ea70fd3} /* (22, 20, 20) {real, imag} */,
  {32'hbd1a288c, 32'hbeb23004} /* (22, 20, 19) {real, imag} */,
  {32'h3e489104, 32'h3f0a4ec4} /* (22, 20, 18) {real, imag} */,
  {32'hbd84ee7e, 32'hbdfd8a6d} /* (22, 20, 17) {real, imag} */,
  {32'hbe0b9f53, 32'hbbe770a0} /* (22, 20, 16) {real, imag} */,
  {32'hbc81b850, 32'hbdac93da} /* (22, 20, 15) {real, imag} */,
  {32'hbf041030, 32'h3cdbb260} /* (22, 20, 14) {real, imag} */,
  {32'h3e3f90a8, 32'h3f0066df} /* (22, 20, 13) {real, imag} */,
  {32'hbe932aa9, 32'hbe91ab0d} /* (22, 20, 12) {real, imag} */,
  {32'h3d3aa90e, 32'h3dbef578} /* (22, 20, 11) {real, imag} */,
  {32'h3f2d47d4, 32'hbe8d8bab} /* (22, 20, 10) {real, imag} */,
  {32'h3ea64c5f, 32'hbda74ef4} /* (22, 20, 9) {real, imag} */,
  {32'hbebb331b, 32'hbd3ac208} /* (22, 20, 8) {real, imag} */,
  {32'h3ea6b59c, 32'hbc852550} /* (22, 20, 7) {real, imag} */,
  {32'hbd12a0ab, 32'hbe287980} /* (22, 20, 6) {real, imag} */,
  {32'h3d74ae70, 32'hbe1f767e} /* (22, 20, 5) {real, imag} */,
  {32'hbe0ab043, 32'h3e86a182} /* (22, 20, 4) {real, imag} */,
  {32'h3e8d3a37, 32'hbe0e0852} /* (22, 20, 3) {real, imag} */,
  {32'h3e92e6c2, 32'hbea48bdd} /* (22, 20, 2) {real, imag} */,
  {32'hbf114350, 32'h3e4a5c70} /* (22, 20, 1) {real, imag} */,
  {32'hbd78ad4c, 32'h3e470210} /* (22, 20, 0) {real, imag} */,
  {32'hbe314100, 32'h3e8f3d34} /* (22, 19, 31) {real, imag} */,
  {32'h3eb1538c, 32'h3ec4299c} /* (22, 19, 30) {real, imag} */,
  {32'h3ef31b75, 32'h3dae944b} /* (22, 19, 29) {real, imag} */,
  {32'hbc15eb20, 32'hbed858fd} /* (22, 19, 28) {real, imag} */,
  {32'hbf1d1002, 32'h3f0f1c1a} /* (22, 19, 27) {real, imag} */,
  {32'h3e7c1072, 32'hbd9cc652} /* (22, 19, 26) {real, imag} */,
  {32'hbd987574, 32'h3ddfab3e} /* (22, 19, 25) {real, imag} */,
  {32'hbeb14535, 32'hbe0bf5d7} /* (22, 19, 24) {real, imag} */,
  {32'h3e6f804a, 32'hbed5309f} /* (22, 19, 23) {real, imag} */,
  {32'h3da4dc1e, 32'hbd907e38} /* (22, 19, 22) {real, imag} */,
  {32'hbf08bc3a, 32'hbdc9dec6} /* (22, 19, 21) {real, imag} */,
  {32'hbe89523c, 32'h3d4e48a8} /* (22, 19, 20) {real, imag} */,
  {32'hbe94d4be, 32'h3e42a0b3} /* (22, 19, 19) {real, imag} */,
  {32'hbee0ce38, 32'hbe800e17} /* (22, 19, 18) {real, imag} */,
  {32'hbce2bf8c, 32'hbebe36c6} /* (22, 19, 17) {real, imag} */,
  {32'h3d68508d, 32'h3e897fa4} /* (22, 19, 16) {real, imag} */,
  {32'hbe1520c0, 32'hbdaff77c} /* (22, 19, 15) {real, imag} */,
  {32'h3d975ead, 32'h3eb473ad} /* (22, 19, 14) {real, imag} */,
  {32'hbdcd6036, 32'h3ea6c6cc} /* (22, 19, 13) {real, imag} */,
  {32'hbdf9fca0, 32'hbd06846a} /* (22, 19, 12) {real, imag} */,
  {32'h3eeb47ea, 32'hbdc71e26} /* (22, 19, 11) {real, imag} */,
  {32'hbe091f76, 32'hbed1736a} /* (22, 19, 10) {real, imag} */,
  {32'h3ec8e99e, 32'h3efa423e} /* (22, 19, 9) {real, imag} */,
  {32'h3e87601c, 32'hbc763180} /* (22, 19, 8) {real, imag} */,
  {32'hbc59d370, 32'hbf036c9f} /* (22, 19, 7) {real, imag} */,
  {32'hbe331ccc, 32'hbeb19a3f} /* (22, 19, 6) {real, imag} */,
  {32'h3ead9cec, 32'h3ec8f865} /* (22, 19, 5) {real, imag} */,
  {32'hbed7fe86, 32'hbe6e942a} /* (22, 19, 4) {real, imag} */,
  {32'hbf02b3ad, 32'h3e2d6a6c} /* (22, 19, 3) {real, imag} */,
  {32'hbeb08ebf, 32'h3e8850e4} /* (22, 19, 2) {real, imag} */,
  {32'h3ed9f7e2, 32'h3e9ecddb} /* (22, 19, 1) {real, imag} */,
  {32'hbe014c90, 32'hbe93c642} /* (22, 19, 0) {real, imag} */,
  {32'hbee3b868, 32'hbf144b45} /* (22, 18, 31) {real, imag} */,
  {32'hbe9d4bed, 32'hbe0aa5ef} /* (22, 18, 30) {real, imag} */,
  {32'h3e854de0, 32'h3e223bc4} /* (22, 18, 29) {real, imag} */,
  {32'hbccbf5bc, 32'hbe5fd2fe} /* (22, 18, 28) {real, imag} */,
  {32'h3df61a04, 32'h3e999bf6} /* (22, 18, 27) {real, imag} */,
  {32'hbe4dd18e, 32'h3eecdec0} /* (22, 18, 26) {real, imag} */,
  {32'hbed0af6e, 32'h3e2ad8f6} /* (22, 18, 25) {real, imag} */,
  {32'h3ec3ccd7, 32'h3cb23337} /* (22, 18, 24) {real, imag} */,
  {32'h3c913e6c, 32'hbe58c696} /* (22, 18, 23) {real, imag} */,
  {32'hbec35194, 32'h3de6e04c} /* (22, 18, 22) {real, imag} */,
  {32'hbdf042ec, 32'hbd3c0da8} /* (22, 18, 21) {real, imag} */,
  {32'hbe8c66ec, 32'h3f241999} /* (22, 18, 20) {real, imag} */,
  {32'hbeb07f3c, 32'hbec777f2} /* (22, 18, 19) {real, imag} */,
  {32'h3e2a3b1b, 32'hbea3939a} /* (22, 18, 18) {real, imag} */,
  {32'h3e834ab7, 32'hbeb53bd4} /* (22, 18, 17) {real, imag} */,
  {32'h3dd2a88a, 32'hbdf3e58a} /* (22, 18, 16) {real, imag} */,
  {32'hbdc6e2b8, 32'h3e1c3470} /* (22, 18, 15) {real, imag} */,
  {32'hbd0f83c4, 32'hbc703258} /* (22, 18, 14) {real, imag} */,
  {32'hbe914e7d, 32'h3dc43ffa} /* (22, 18, 13) {real, imag} */,
  {32'h3dd5e85a, 32'hbed6bdcd} /* (22, 18, 12) {real, imag} */,
  {32'hbcd10c30, 32'hbdda6584} /* (22, 18, 11) {real, imag} */,
  {32'h3ee19a92, 32'h3e9c7aa4} /* (22, 18, 10) {real, imag} */,
  {32'hbe6af2e9, 32'h3e12c309} /* (22, 18, 9) {real, imag} */,
  {32'hbeef6275, 32'hbcf507b4} /* (22, 18, 8) {real, imag} */,
  {32'h3ed7cdca, 32'h3f3f3b3a} /* (22, 18, 7) {real, imag} */,
  {32'h3e982fe2, 32'h3ec071b4} /* (22, 18, 6) {real, imag} */,
  {32'h3d7aea97, 32'h3ebaca4a} /* (22, 18, 5) {real, imag} */,
  {32'h3da348eb, 32'hbe3079c0} /* (22, 18, 4) {real, imag} */,
  {32'h3da0255c, 32'h3e6f72f5} /* (22, 18, 3) {real, imag} */,
  {32'hbea58f32, 32'h3f032756} /* (22, 18, 2) {real, imag} */,
  {32'h3d1ff0c4, 32'hbe13cfda} /* (22, 18, 1) {real, imag} */,
  {32'hbebd81dd, 32'hbf03976a} /* (22, 18, 0) {real, imag} */,
  {32'hbea5d50e, 32'h3eb65aa2} /* (22, 17, 31) {real, imag} */,
  {32'h3e79d3c4, 32'h3df57818} /* (22, 17, 30) {real, imag} */,
  {32'hbc678170, 32'hbd473a22} /* (22, 17, 29) {real, imag} */,
  {32'hbd3b6932, 32'h3ea1daeb} /* (22, 17, 28) {real, imag} */,
  {32'hbe37cda5, 32'h3ee10e3c} /* (22, 17, 27) {real, imag} */,
  {32'hbd3f0512, 32'hbe1e947e} /* (22, 17, 26) {real, imag} */,
  {32'h3e052eb8, 32'hbe4b68c7} /* (22, 17, 25) {real, imag} */,
  {32'h3ec25e20, 32'h3db9bcb2} /* (22, 17, 24) {real, imag} */,
  {32'hbe57633f, 32'hbd214494} /* (22, 17, 23) {real, imag} */,
  {32'hbf4b4da4, 32'hbeb10cfd} /* (22, 17, 22) {real, imag} */,
  {32'hbe51cd00, 32'h3d7a89d8} /* (22, 17, 21) {real, imag} */,
  {32'h3f1e4bf4, 32'hbd7d180b} /* (22, 17, 20) {real, imag} */,
  {32'h3e2f5f65, 32'hbe4535e4} /* (22, 17, 19) {real, imag} */,
  {32'h3e1e5804, 32'hbedcb78e} /* (22, 17, 18) {real, imag} */,
  {32'h3e0ced19, 32'h3cbeae18} /* (22, 17, 17) {real, imag} */,
  {32'h3d165807, 32'h3dff78ce} /* (22, 17, 16) {real, imag} */,
  {32'h3d919180, 32'h3cb8dc98} /* (22, 17, 15) {real, imag} */,
  {32'h3dab4fc7, 32'h3df959e8} /* (22, 17, 14) {real, imag} */,
  {32'h3cef723c, 32'hbf277284} /* (22, 17, 13) {real, imag} */,
  {32'hbef454c0, 32'h3e82299e} /* (22, 17, 12) {real, imag} */,
  {32'h3ed572b2, 32'hbdbf4ede} /* (22, 17, 11) {real, imag} */,
  {32'hbe566142, 32'h3dd24d18} /* (22, 17, 10) {real, imag} */,
  {32'h3e9dfe92, 32'h3c3f0700} /* (22, 17, 9) {real, imag} */,
  {32'h3ea7402d, 32'hbda49580} /* (22, 17, 8) {real, imag} */,
  {32'h3e6e22dd, 32'h3f00adbe} /* (22, 17, 7) {real, imag} */,
  {32'hbe183b81, 32'h3a9f4d80} /* (22, 17, 6) {real, imag} */,
  {32'hbe71bd51, 32'hbd340f08} /* (22, 17, 5) {real, imag} */,
  {32'hbdece1e4, 32'hbc7e66d0} /* (22, 17, 4) {real, imag} */,
  {32'hbe87bf94, 32'hbdb80996} /* (22, 17, 3) {real, imag} */,
  {32'hbe4d3e52, 32'hbef7e92c} /* (22, 17, 2) {real, imag} */,
  {32'h3e2ae46a, 32'hbc10d380} /* (22, 17, 1) {real, imag} */,
  {32'hbdf3f2b1, 32'hbc7a2a88} /* (22, 17, 0) {real, imag} */,
  {32'h3e45dad2, 32'hbdf4aee8} /* (22, 16, 31) {real, imag} */,
  {32'h3e29db77, 32'h3e508986} /* (22, 16, 30) {real, imag} */,
  {32'hbdc3fad8, 32'h3e94e719} /* (22, 16, 29) {real, imag} */,
  {32'hbdd3a227, 32'h3dace7da} /* (22, 16, 28) {real, imag} */,
  {32'h3af556c0, 32'hbc24b968} /* (22, 16, 27) {real, imag} */,
  {32'h3e0d85a8, 32'h3c82b89a} /* (22, 16, 26) {real, imag} */,
  {32'hbe020115, 32'hbd7b7207} /* (22, 16, 25) {real, imag} */,
  {32'h3d62e398, 32'hbe6306ad} /* (22, 16, 24) {real, imag} */,
  {32'hbe1dceaa, 32'h3dab25c6} /* (22, 16, 23) {real, imag} */,
  {32'hbec93698, 32'h3d9755ac} /* (22, 16, 22) {real, imag} */,
  {32'h3e454cd6, 32'hbe6a132a} /* (22, 16, 21) {real, imag} */,
  {32'hbe4db665, 32'h3e8704b5} /* (22, 16, 20) {real, imag} */,
  {32'h3dd5ba7b, 32'h3e23d5f0} /* (22, 16, 19) {real, imag} */,
  {32'h3ed3d9d6, 32'h3e9ab7be} /* (22, 16, 18) {real, imag} */,
  {32'hbcb83838, 32'h3cde4ca4} /* (22, 16, 17) {real, imag} */,
  {32'hbe581f1d, 32'h00000000} /* (22, 16, 16) {real, imag} */,
  {32'hbcb83838, 32'hbcde4ca4} /* (22, 16, 15) {real, imag} */,
  {32'h3ed3d9d6, 32'hbe9ab7be} /* (22, 16, 14) {real, imag} */,
  {32'h3dd5ba7b, 32'hbe23d5f0} /* (22, 16, 13) {real, imag} */,
  {32'hbe4db665, 32'hbe8704b5} /* (22, 16, 12) {real, imag} */,
  {32'h3e454cd6, 32'h3e6a132a} /* (22, 16, 11) {real, imag} */,
  {32'hbec93698, 32'hbd9755ac} /* (22, 16, 10) {real, imag} */,
  {32'hbe1dceaa, 32'hbdab25c6} /* (22, 16, 9) {real, imag} */,
  {32'h3d62e398, 32'h3e6306ad} /* (22, 16, 8) {real, imag} */,
  {32'hbe020115, 32'h3d7b7207} /* (22, 16, 7) {real, imag} */,
  {32'h3e0d85a8, 32'hbc82b89a} /* (22, 16, 6) {real, imag} */,
  {32'h3af556c0, 32'h3c24b968} /* (22, 16, 5) {real, imag} */,
  {32'hbdd3a227, 32'hbdace7da} /* (22, 16, 4) {real, imag} */,
  {32'hbdc3fad8, 32'hbe94e719} /* (22, 16, 3) {real, imag} */,
  {32'h3e29db77, 32'hbe508986} /* (22, 16, 2) {real, imag} */,
  {32'h3e45dad2, 32'h3df4aee8} /* (22, 16, 1) {real, imag} */,
  {32'h3ef7ec54, 32'h00000000} /* (22, 16, 0) {real, imag} */,
  {32'h3e2ae46a, 32'h3c10d380} /* (22, 15, 31) {real, imag} */,
  {32'hbe4d3e52, 32'h3ef7e92c} /* (22, 15, 30) {real, imag} */,
  {32'hbe87bf94, 32'h3db80996} /* (22, 15, 29) {real, imag} */,
  {32'hbdece1e4, 32'h3c7e66d0} /* (22, 15, 28) {real, imag} */,
  {32'hbe71bd51, 32'h3d340f08} /* (22, 15, 27) {real, imag} */,
  {32'hbe183b81, 32'hba9f4d80} /* (22, 15, 26) {real, imag} */,
  {32'h3e6e22dd, 32'hbf00adbe} /* (22, 15, 25) {real, imag} */,
  {32'h3ea7402d, 32'h3da49580} /* (22, 15, 24) {real, imag} */,
  {32'h3e9dfe92, 32'hbc3f0700} /* (22, 15, 23) {real, imag} */,
  {32'hbe566142, 32'hbdd24d18} /* (22, 15, 22) {real, imag} */,
  {32'h3ed572b2, 32'h3dbf4ede} /* (22, 15, 21) {real, imag} */,
  {32'hbef454c0, 32'hbe82299e} /* (22, 15, 20) {real, imag} */,
  {32'h3cef723c, 32'h3f277284} /* (22, 15, 19) {real, imag} */,
  {32'h3dab4fc7, 32'hbdf959e8} /* (22, 15, 18) {real, imag} */,
  {32'h3d919180, 32'hbcb8dc98} /* (22, 15, 17) {real, imag} */,
  {32'h3d165807, 32'hbdff78ce} /* (22, 15, 16) {real, imag} */,
  {32'h3e0ced19, 32'hbcbeae18} /* (22, 15, 15) {real, imag} */,
  {32'h3e1e5804, 32'h3edcb78e} /* (22, 15, 14) {real, imag} */,
  {32'h3e2f5f65, 32'h3e4535e4} /* (22, 15, 13) {real, imag} */,
  {32'h3f1e4bf4, 32'h3d7d180b} /* (22, 15, 12) {real, imag} */,
  {32'hbe51cd00, 32'hbd7a89d8} /* (22, 15, 11) {real, imag} */,
  {32'hbf4b4da4, 32'h3eb10cfd} /* (22, 15, 10) {real, imag} */,
  {32'hbe57633f, 32'h3d214494} /* (22, 15, 9) {real, imag} */,
  {32'h3ec25e20, 32'hbdb9bcb2} /* (22, 15, 8) {real, imag} */,
  {32'h3e052eb8, 32'h3e4b68c7} /* (22, 15, 7) {real, imag} */,
  {32'hbd3f0512, 32'h3e1e947e} /* (22, 15, 6) {real, imag} */,
  {32'hbe37cda5, 32'hbee10e3c} /* (22, 15, 5) {real, imag} */,
  {32'hbd3b6932, 32'hbea1daeb} /* (22, 15, 4) {real, imag} */,
  {32'hbc678170, 32'h3d473a22} /* (22, 15, 3) {real, imag} */,
  {32'h3e79d3c4, 32'hbdf57818} /* (22, 15, 2) {real, imag} */,
  {32'hbea5d50e, 32'hbeb65aa2} /* (22, 15, 1) {real, imag} */,
  {32'hbdf3f2b1, 32'h3c7a2a88} /* (22, 15, 0) {real, imag} */,
  {32'h3d1ff0c4, 32'h3e13cfda} /* (22, 14, 31) {real, imag} */,
  {32'hbea58f32, 32'hbf032756} /* (22, 14, 30) {real, imag} */,
  {32'h3da0255c, 32'hbe6f72f5} /* (22, 14, 29) {real, imag} */,
  {32'h3da348eb, 32'h3e3079c0} /* (22, 14, 28) {real, imag} */,
  {32'h3d7aea97, 32'hbebaca4a} /* (22, 14, 27) {real, imag} */,
  {32'h3e982fe2, 32'hbec071b4} /* (22, 14, 26) {real, imag} */,
  {32'h3ed7cdca, 32'hbf3f3b3a} /* (22, 14, 25) {real, imag} */,
  {32'hbeef6275, 32'h3cf507b4} /* (22, 14, 24) {real, imag} */,
  {32'hbe6af2e9, 32'hbe12c309} /* (22, 14, 23) {real, imag} */,
  {32'h3ee19a92, 32'hbe9c7aa4} /* (22, 14, 22) {real, imag} */,
  {32'hbcd10c30, 32'h3dda6584} /* (22, 14, 21) {real, imag} */,
  {32'h3dd5e85a, 32'h3ed6bdcd} /* (22, 14, 20) {real, imag} */,
  {32'hbe914e7d, 32'hbdc43ffa} /* (22, 14, 19) {real, imag} */,
  {32'hbd0f83c4, 32'h3c703258} /* (22, 14, 18) {real, imag} */,
  {32'hbdc6e2b8, 32'hbe1c3470} /* (22, 14, 17) {real, imag} */,
  {32'h3dd2a88a, 32'h3df3e58a} /* (22, 14, 16) {real, imag} */,
  {32'h3e834ab7, 32'h3eb53bd4} /* (22, 14, 15) {real, imag} */,
  {32'h3e2a3b1b, 32'h3ea3939a} /* (22, 14, 14) {real, imag} */,
  {32'hbeb07f3c, 32'h3ec777f2} /* (22, 14, 13) {real, imag} */,
  {32'hbe8c66ec, 32'hbf241999} /* (22, 14, 12) {real, imag} */,
  {32'hbdf042ec, 32'h3d3c0da8} /* (22, 14, 11) {real, imag} */,
  {32'hbec35194, 32'hbde6e04c} /* (22, 14, 10) {real, imag} */,
  {32'h3c913e6c, 32'h3e58c696} /* (22, 14, 9) {real, imag} */,
  {32'h3ec3ccd7, 32'hbcb23337} /* (22, 14, 8) {real, imag} */,
  {32'hbed0af6e, 32'hbe2ad8f6} /* (22, 14, 7) {real, imag} */,
  {32'hbe4dd18e, 32'hbeecdec0} /* (22, 14, 6) {real, imag} */,
  {32'h3df61a04, 32'hbe999bf6} /* (22, 14, 5) {real, imag} */,
  {32'hbccbf5bc, 32'h3e5fd2fe} /* (22, 14, 4) {real, imag} */,
  {32'h3e854de0, 32'hbe223bc4} /* (22, 14, 3) {real, imag} */,
  {32'hbe9d4bed, 32'h3e0aa5ef} /* (22, 14, 2) {real, imag} */,
  {32'hbee3b868, 32'h3f144b45} /* (22, 14, 1) {real, imag} */,
  {32'hbebd81dd, 32'h3f03976a} /* (22, 14, 0) {real, imag} */,
  {32'h3ed9f7e2, 32'hbe9ecddb} /* (22, 13, 31) {real, imag} */,
  {32'hbeb08ebf, 32'hbe8850e4} /* (22, 13, 30) {real, imag} */,
  {32'hbf02b3ad, 32'hbe2d6a6c} /* (22, 13, 29) {real, imag} */,
  {32'hbed7fe86, 32'h3e6e942a} /* (22, 13, 28) {real, imag} */,
  {32'h3ead9cec, 32'hbec8f865} /* (22, 13, 27) {real, imag} */,
  {32'hbe331ccc, 32'h3eb19a3f} /* (22, 13, 26) {real, imag} */,
  {32'hbc59d370, 32'h3f036c9f} /* (22, 13, 25) {real, imag} */,
  {32'h3e87601c, 32'h3c763180} /* (22, 13, 24) {real, imag} */,
  {32'h3ec8e99e, 32'hbefa423e} /* (22, 13, 23) {real, imag} */,
  {32'hbe091f76, 32'h3ed1736a} /* (22, 13, 22) {real, imag} */,
  {32'h3eeb47ea, 32'h3dc71e26} /* (22, 13, 21) {real, imag} */,
  {32'hbdf9fca0, 32'h3d06846a} /* (22, 13, 20) {real, imag} */,
  {32'hbdcd6036, 32'hbea6c6cc} /* (22, 13, 19) {real, imag} */,
  {32'h3d975ead, 32'hbeb473ad} /* (22, 13, 18) {real, imag} */,
  {32'hbe1520c0, 32'h3daff77c} /* (22, 13, 17) {real, imag} */,
  {32'h3d68508d, 32'hbe897fa4} /* (22, 13, 16) {real, imag} */,
  {32'hbce2bf8c, 32'h3ebe36c6} /* (22, 13, 15) {real, imag} */,
  {32'hbee0ce38, 32'h3e800e17} /* (22, 13, 14) {real, imag} */,
  {32'hbe94d4be, 32'hbe42a0b3} /* (22, 13, 13) {real, imag} */,
  {32'hbe89523c, 32'hbd4e48a8} /* (22, 13, 12) {real, imag} */,
  {32'hbf08bc3a, 32'h3dc9dec6} /* (22, 13, 11) {real, imag} */,
  {32'h3da4dc1e, 32'h3d907e38} /* (22, 13, 10) {real, imag} */,
  {32'h3e6f804a, 32'h3ed5309f} /* (22, 13, 9) {real, imag} */,
  {32'hbeb14535, 32'h3e0bf5d7} /* (22, 13, 8) {real, imag} */,
  {32'hbd987574, 32'hbddfab3e} /* (22, 13, 7) {real, imag} */,
  {32'h3e7c1072, 32'h3d9cc652} /* (22, 13, 6) {real, imag} */,
  {32'hbf1d1002, 32'hbf0f1c1a} /* (22, 13, 5) {real, imag} */,
  {32'hbc15eb20, 32'h3ed858fd} /* (22, 13, 4) {real, imag} */,
  {32'h3ef31b75, 32'hbdae944b} /* (22, 13, 3) {real, imag} */,
  {32'h3eb1538c, 32'hbec4299c} /* (22, 13, 2) {real, imag} */,
  {32'hbe314100, 32'hbe8f3d34} /* (22, 13, 1) {real, imag} */,
  {32'hbe014c90, 32'h3e93c642} /* (22, 13, 0) {real, imag} */,
  {32'hbf114350, 32'hbe4a5c70} /* (22, 12, 31) {real, imag} */,
  {32'h3e92e6c2, 32'h3ea48bdd} /* (22, 12, 30) {real, imag} */,
  {32'h3e8d3a37, 32'h3e0e0852} /* (22, 12, 29) {real, imag} */,
  {32'hbe0ab043, 32'hbe86a182} /* (22, 12, 28) {real, imag} */,
  {32'h3d74ae70, 32'h3e1f767e} /* (22, 12, 27) {real, imag} */,
  {32'hbd12a0ab, 32'h3e287980} /* (22, 12, 26) {real, imag} */,
  {32'h3ea6b59c, 32'h3c852550} /* (22, 12, 25) {real, imag} */,
  {32'hbebb331b, 32'h3d3ac208} /* (22, 12, 24) {real, imag} */,
  {32'h3ea64c5f, 32'h3da74ef4} /* (22, 12, 23) {real, imag} */,
  {32'h3f2d47d4, 32'h3e8d8bab} /* (22, 12, 22) {real, imag} */,
  {32'h3d3aa90e, 32'hbdbef578} /* (22, 12, 21) {real, imag} */,
  {32'hbe932aa9, 32'h3e91ab0d} /* (22, 12, 20) {real, imag} */,
  {32'h3e3f90a8, 32'hbf0066df} /* (22, 12, 19) {real, imag} */,
  {32'hbf041030, 32'hbcdbb260} /* (22, 12, 18) {real, imag} */,
  {32'hbc81b850, 32'h3dac93da} /* (22, 12, 17) {real, imag} */,
  {32'hbe0b9f53, 32'h3be770a0} /* (22, 12, 16) {real, imag} */,
  {32'hbd84ee7e, 32'h3dfd8a6d} /* (22, 12, 15) {real, imag} */,
  {32'h3e489104, 32'hbf0a4ec4} /* (22, 12, 14) {real, imag} */,
  {32'hbd1a288c, 32'h3eb23004} /* (22, 12, 13) {real, imag} */,
  {32'h3ee59c80, 32'hbea70fd3} /* (22, 12, 12) {real, imag} */,
  {32'h3dd847ee, 32'h3e7963ff} /* (22, 12, 11) {real, imag} */,
  {32'h3e9349cc, 32'h3d269958} /* (22, 12, 10) {real, imag} */,
  {32'h3ebbdccc, 32'hbc35eb60} /* (22, 12, 9) {real, imag} */,
  {32'hbe6120ba, 32'h3ea137f2} /* (22, 12, 8) {real, imag} */,
  {32'hbe4a6606, 32'h3e9005a0} /* (22, 12, 7) {real, imag} */,
  {32'h3e10c3e9, 32'hbd8b20bb} /* (22, 12, 6) {real, imag} */,
  {32'h3e5b55b6, 32'h3f47d110} /* (22, 12, 5) {real, imag} */,
  {32'h3d946c24, 32'hbe0905b5} /* (22, 12, 4) {real, imag} */,
  {32'hbad2b340, 32'hbe80f2cc} /* (22, 12, 3) {real, imag} */,
  {32'h3e3aa854, 32'hbe18a69a} /* (22, 12, 2) {real, imag} */,
  {32'hbcbf298e, 32'h3da31ea6} /* (22, 12, 1) {real, imag} */,
  {32'hbd78ad4c, 32'hbe470210} /* (22, 12, 0) {real, imag} */,
  {32'h3e803910, 32'h3e90caa4} /* (22, 11, 31) {real, imag} */,
  {32'hbe4746e0, 32'hbf44c023} /* (22, 11, 30) {real, imag} */,
  {32'h3e0ed08e, 32'hbd6e7294} /* (22, 11, 29) {real, imag} */,
  {32'hbe59efb1, 32'hbe0aa936} /* (22, 11, 28) {real, imag} */,
  {32'hbcc8fa24, 32'hbf1ed968} /* (22, 11, 27) {real, imag} */,
  {32'h3c769840, 32'h3ea47110} /* (22, 11, 26) {real, imag} */,
  {32'hbe35202e, 32'h3f14c302} /* (22, 11, 25) {real, imag} */,
  {32'h3e845016, 32'h3d23fe18} /* (22, 11, 24) {real, imag} */,
  {32'hbedc7b3b, 32'h3f0aaa5a} /* (22, 11, 23) {real, imag} */,
  {32'hbf2eded1, 32'hbdaa374c} /* (22, 11, 22) {real, imag} */,
  {32'hbe378b1d, 32'hbe086bf8} /* (22, 11, 21) {real, imag} */,
  {32'h3e58c2f0, 32'h3cdf94f8} /* (22, 11, 20) {real, imag} */,
  {32'h3dbcd7b1, 32'hbc8a09f8} /* (22, 11, 19) {real, imag} */,
  {32'hbe9df448, 32'h3ecf0619} /* (22, 11, 18) {real, imag} */,
  {32'h3e9f54d3, 32'hbdb3f33e} /* (22, 11, 17) {real, imag} */,
  {32'hbc4119d0, 32'h3e5ca602} /* (22, 11, 16) {real, imag} */,
  {32'hbd56a005, 32'hbc5bad90} /* (22, 11, 15) {real, imag} */,
  {32'h3e4881dd, 32'h3e41d402} /* (22, 11, 14) {real, imag} */,
  {32'hbe72b125, 32'h3edbb445} /* (22, 11, 13) {real, imag} */,
  {32'h3eadb0d6, 32'h3f30bc9a} /* (22, 11, 12) {real, imag} */,
  {32'hbf078182, 32'hbe098eb0} /* (22, 11, 11) {real, imag} */,
  {32'hbd756f12, 32'h3e28c722} /* (22, 11, 10) {real, imag} */,
  {32'hbe09ca3e, 32'h3f85e66c} /* (22, 11, 9) {real, imag} */,
  {32'hbdb36229, 32'hbe9e395e} /* (22, 11, 8) {real, imag} */,
  {32'hbde2cce0, 32'hbe1dc849} /* (22, 11, 7) {real, imag} */,
  {32'hbf555511, 32'h3e37e8a2} /* (22, 11, 6) {real, imag} */,
  {32'hbed951da, 32'h3ef686e0} /* (22, 11, 5) {real, imag} */,
  {32'h3e846f58, 32'h3f190675} /* (22, 11, 4) {real, imag} */,
  {32'hbda07cf0, 32'hbe30bf5f} /* (22, 11, 3) {real, imag} */,
  {32'h3d5c9170, 32'hbde5075c} /* (22, 11, 2) {real, imag} */,
  {32'hbd1a2989, 32'h3f624284} /* (22, 11, 1) {real, imag} */,
  {32'h3e5a7052, 32'h3ebe6be2} /* (22, 11, 0) {real, imag} */,
  {32'h3d9e6ff8, 32'hbefa19cb} /* (22, 10, 31) {real, imag} */,
  {32'hbe868551, 32'h3e43a112} /* (22, 10, 30) {real, imag} */,
  {32'hbdb28002, 32'hbf2cd678} /* (22, 10, 29) {real, imag} */,
  {32'hbea44114, 32'hbeb32a8a} /* (22, 10, 28) {real, imag} */,
  {32'h3d708c98, 32'hbf031928} /* (22, 10, 27) {real, imag} */,
  {32'hbde0b63e, 32'hbdd9f8fc} /* (22, 10, 26) {real, imag} */,
  {32'hbe436150, 32'hbdf7c867} /* (22, 10, 25) {real, imag} */,
  {32'h3ea85826, 32'hbb107600} /* (22, 10, 24) {real, imag} */,
  {32'hbd5300a0, 32'h3d2c69a0} /* (22, 10, 23) {real, imag} */,
  {32'h3e014a0c, 32'hbebc4d40} /* (22, 10, 22) {real, imag} */,
  {32'hbe9ffd89, 32'hbe32bc9e} /* (22, 10, 21) {real, imag} */,
  {32'h3f409cb0, 32'h3d9956f0} /* (22, 10, 20) {real, imag} */,
  {32'hbe3d6bb0, 32'h3be26800} /* (22, 10, 19) {real, imag} */,
  {32'h3d82ef9a, 32'h3e83d3db} /* (22, 10, 18) {real, imag} */,
  {32'hbe847320, 32'hbd7136c2} /* (22, 10, 17) {real, imag} */,
  {32'hbd98b262, 32'hbd93c91f} /* (22, 10, 16) {real, imag} */,
  {32'h3c979c48, 32'hbe28a8a4} /* (22, 10, 15) {real, imag} */,
  {32'hbd403668, 32'h3aecd400} /* (22, 10, 14) {real, imag} */,
  {32'h3eb9aa2b, 32'h3f19c92d} /* (22, 10, 13) {real, imag} */,
  {32'hbe652cec, 32'hbeb0e0db} /* (22, 10, 12) {real, imag} */,
  {32'hbe92c0aa, 32'hbe43c5e1} /* (22, 10, 11) {real, imag} */,
  {32'hbf1b12a4, 32'h3d7c0af0} /* (22, 10, 10) {real, imag} */,
  {32'hbe04a6f4, 32'h3e82639c} /* (22, 10, 9) {real, imag} */,
  {32'hbe3ae46b, 32'h3e17de57} /* (22, 10, 8) {real, imag} */,
  {32'hbe23abc2, 32'hbe57ceb0} /* (22, 10, 7) {real, imag} */,
  {32'h3c3146a0, 32'h3f063872} /* (22, 10, 6) {real, imag} */,
  {32'hbeb3cdb6, 32'h3ee6d7e3} /* (22, 10, 5) {real, imag} */,
  {32'h3d6e6e53, 32'hbe5b33ef} /* (22, 10, 4) {real, imag} */,
  {32'h3eb9e037, 32'hbed1bce4} /* (22, 10, 3) {real, imag} */,
  {32'h3dcd29c4, 32'h3f20ae24} /* (22, 10, 2) {real, imag} */,
  {32'hbef5f9f3, 32'hbf26a64c} /* (22, 10, 1) {real, imag} */,
  {32'hbd184f34, 32'hbed5420c} /* (22, 10, 0) {real, imag} */,
  {32'h3ee0f5a0, 32'hbe771154} /* (22, 9, 31) {real, imag} */,
  {32'h3eb617ae, 32'h3f26955a} /* (22, 9, 30) {real, imag} */,
  {32'h3afa0bc0, 32'hbe5a0497} /* (22, 9, 29) {real, imag} */,
  {32'h3cc4a8c0, 32'h3f69db56} /* (22, 9, 28) {real, imag} */,
  {32'h3edd8f46, 32'h3cd4d198} /* (22, 9, 27) {real, imag} */,
  {32'hbeb526f1, 32'h3e8a7080} /* (22, 9, 26) {real, imag} */,
  {32'hbec7a8e8, 32'hbf02cae7} /* (22, 9, 25) {real, imag} */,
  {32'h3e83cfa6, 32'hbdf4f100} /* (22, 9, 24) {real, imag} */,
  {32'hbe0c2066, 32'hbdbf9dd8} /* (22, 9, 23) {real, imag} */,
  {32'h3e8717e4, 32'h3f12538c} /* (22, 9, 22) {real, imag} */,
  {32'hbe850f30, 32'h3e2b1c36} /* (22, 9, 21) {real, imag} */,
  {32'h3e2544ea, 32'h3df6113c} /* (22, 9, 20) {real, imag} */,
  {32'h3da17952, 32'hbecb4666} /* (22, 9, 19) {real, imag} */,
  {32'hbdce4362, 32'h3e567db9} /* (22, 9, 18) {real, imag} */,
  {32'hbe19be2f, 32'h3eb4fd80} /* (22, 9, 17) {real, imag} */,
  {32'hbdf4b04e, 32'h3d1cc73a} /* (22, 9, 16) {real, imag} */,
  {32'h3f16e4d8, 32'h3cfe2078} /* (22, 9, 15) {real, imag} */,
  {32'h3c836740, 32'hbe94e742} /* (22, 9, 14) {real, imag} */,
  {32'hbee8021e, 32'h3d53443c} /* (22, 9, 13) {real, imag} */,
  {32'h3e846a88, 32'hbf03578a} /* (22, 9, 12) {real, imag} */,
  {32'h3ded52fa, 32'h3ce9c8f8} /* (22, 9, 11) {real, imag} */,
  {32'hbdbe2834, 32'h3e5a4ff6} /* (22, 9, 10) {real, imag} */,
  {32'h3f14c7b8, 32'hbf11d592} /* (22, 9, 9) {real, imag} */,
  {32'h3f0d77de, 32'h3f1e6f9a} /* (22, 9, 8) {real, imag} */,
  {32'h3ef88d0a, 32'h3d007fa8} /* (22, 9, 7) {real, imag} */,
  {32'hbf5bf7b6, 32'hbe79aab9} /* (22, 9, 6) {real, imag} */,
  {32'hbd163938, 32'hbc457f20} /* (22, 9, 5) {real, imag} */,
  {32'h3eeceb87, 32'hbdad917e} /* (22, 9, 4) {real, imag} */,
  {32'h3e5be485, 32'h3f3a0f44} /* (22, 9, 3) {real, imag} */,
  {32'h3e5ea2d2, 32'h3e726056} /* (22, 9, 2) {real, imag} */,
  {32'hbeb668f0, 32'hbf341f1c} /* (22, 9, 1) {real, imag} */,
  {32'h3a44c380, 32'h3f0778a3} /* (22, 9, 0) {real, imag} */,
  {32'h3fa1e523, 32'h3f2ccf87} /* (22, 8, 31) {real, imag} */,
  {32'hbf265f70, 32'hbde2ef98} /* (22, 8, 30) {real, imag} */,
  {32'hbbd8e480, 32'h3eaa1da8} /* (22, 8, 29) {real, imag} */,
  {32'h3e4234ba, 32'hbe96adec} /* (22, 8, 28) {real, imag} */,
  {32'hbf7767f4, 32'hbe7d2656} /* (22, 8, 27) {real, imag} */,
  {32'h3cc58ecc, 32'hbe0f167a} /* (22, 8, 26) {real, imag} */,
  {32'h3e988029, 32'h3f23d7ea} /* (22, 8, 25) {real, imag} */,
  {32'hbe648a0e, 32'hbe959480} /* (22, 8, 24) {real, imag} */,
  {32'h3ed59cda, 32'h3d1fd8fa} /* (22, 8, 23) {real, imag} */,
  {32'hbed1c784, 32'hbe988649} /* (22, 8, 22) {real, imag} */,
  {32'hbe6f5480, 32'h3eb44aa6} /* (22, 8, 21) {real, imag} */,
  {32'hbe317df2, 32'h3dd72944} /* (22, 8, 20) {real, imag} */,
  {32'hbea76f60, 32'hbe65f2ac} /* (22, 8, 19) {real, imag} */,
  {32'hbdf5c764, 32'hbe5db011} /* (22, 8, 18) {real, imag} */,
  {32'hbbb0d948, 32'hbdb51b24} /* (22, 8, 17) {real, imag} */,
  {32'hbeda6224, 32'h3d82520a} /* (22, 8, 16) {real, imag} */,
  {32'hbd74420c, 32'h3d28dc81} /* (22, 8, 15) {real, imag} */,
  {32'h3e3c1594, 32'hbf05fac3} /* (22, 8, 14) {real, imag} */,
  {32'hbec99845, 32'hbe923204} /* (22, 8, 13) {real, imag} */,
  {32'hbeb9c91a, 32'h3cc4632c} /* (22, 8, 12) {real, imag} */,
  {32'h3f282a69, 32'hbe489583} /* (22, 8, 11) {real, imag} */,
  {32'hbd059606, 32'h3f0c7c12} /* (22, 8, 10) {real, imag} */,
  {32'hbce01f88, 32'h3e9013b2} /* (22, 8, 9) {real, imag} */,
  {32'hbed614ca, 32'hbece72d1} /* (22, 8, 8) {real, imag} */,
  {32'h3f08fee8, 32'hbe958c42} /* (22, 8, 7) {real, imag} */,
  {32'h3d8450a6, 32'h3dc45bfa} /* (22, 8, 6) {real, imag} */,
  {32'hbf43f168, 32'hbe94d480} /* (22, 8, 5) {real, imag} */,
  {32'h3ee855cc, 32'h3f174d68} /* (22, 8, 4) {real, imag} */,
  {32'h3d175e78, 32'hbec1ca30} /* (22, 8, 3) {real, imag} */,
  {32'hbe0acbbc, 32'h3db25fbc} /* (22, 8, 2) {real, imag} */,
  {32'h3d309408, 32'h3e80b8d0} /* (22, 8, 1) {real, imag} */,
  {32'h3f4836bc, 32'hbcce39f0} /* (22, 8, 0) {real, imag} */,
  {32'hbf2b9732, 32'hbf194f12} /* (22, 7, 31) {real, imag} */,
  {32'h3e938f8e, 32'h3dccb8a4} /* (22, 7, 30) {real, imag} */,
  {32'h3f2ccc00, 32'h3e6c65aa} /* (22, 7, 29) {real, imag} */,
  {32'h3f18ee7e, 32'h3ec4ac83} /* (22, 7, 28) {real, imag} */,
  {32'hbd8dff9c, 32'h3dd11860} /* (22, 7, 27) {real, imag} */,
  {32'hbeb23ec0, 32'h3ec8946c} /* (22, 7, 26) {real, imag} */,
  {32'h3e351048, 32'h3c5960d0} /* (22, 7, 25) {real, imag} */,
  {32'hbf7ede80, 32'h3dd8fada} /* (22, 7, 24) {real, imag} */,
  {32'h3eecc39c, 32'h3e9bb4c1} /* (22, 7, 23) {real, imag} */,
  {32'hbe733b7f, 32'hbdca8c68} /* (22, 7, 22) {real, imag} */,
  {32'h3ed25f6f, 32'hbd322162} /* (22, 7, 21) {real, imag} */,
  {32'h3d1dd128, 32'hbf0737ad} /* (22, 7, 20) {real, imag} */,
  {32'hbeff67d8, 32'h3e6a6ede} /* (22, 7, 19) {real, imag} */,
  {32'h3e8a371e, 32'hbd5a6f24} /* (22, 7, 18) {real, imag} */,
  {32'h3e8df84d, 32'hbe653efa} /* (22, 7, 17) {real, imag} */,
  {32'h3e09a110, 32'h3e2fb7e3} /* (22, 7, 16) {real, imag} */,
  {32'h3d3da130, 32'h3e8cc1ed} /* (22, 7, 15) {real, imag} */,
  {32'hbe531a67, 32'h3b82df40} /* (22, 7, 14) {real, imag} */,
  {32'h3dbf3eb6, 32'h3db9a450} /* (22, 7, 13) {real, imag} */,
  {32'hbe0dfb04, 32'h3e62de5c} /* (22, 7, 12) {real, imag} */,
  {32'hbf412ec4, 32'h3cf9bcb8} /* (22, 7, 11) {real, imag} */,
  {32'hbea41624, 32'h3ea44048} /* (22, 7, 10) {real, imag} */,
  {32'hbdd8415e, 32'hbd284cfc} /* (22, 7, 9) {real, imag} */,
  {32'h3e469615, 32'hbeda709b} /* (22, 7, 8) {real, imag} */,
  {32'hbe23cd84, 32'hbf7b595c} /* (22, 7, 7) {real, imag} */,
  {32'h3e8207e4, 32'h3e2dbc15} /* (22, 7, 6) {real, imag} */,
  {32'h3e1be992, 32'h3e8778ad} /* (22, 7, 5) {real, imag} */,
  {32'h3cd47e88, 32'hbed56654} /* (22, 7, 4) {real, imag} */,
  {32'h3eba04ed, 32'h3f97fc00} /* (22, 7, 3) {real, imag} */,
  {32'hbe98243d, 32'hbe923a1f} /* (22, 7, 2) {real, imag} */,
  {32'hbdfe6088, 32'hbf1a0693} /* (22, 7, 1) {real, imag} */,
  {32'hbe1c0135, 32'hbf086aca} /* (22, 7, 0) {real, imag} */,
  {32'h3e9730e6, 32'h3e70ccd4} /* (22, 6, 31) {real, imag} */,
  {32'hbe5aba98, 32'hbe5e9f77} /* (22, 6, 30) {real, imag} */,
  {32'h3e5784e1, 32'h3edbcf7c} /* (22, 6, 29) {real, imag} */,
  {32'hbd8926ec, 32'hbf2c5217} /* (22, 6, 28) {real, imag} */,
  {32'hbdd5aec8, 32'hbe3d3122} /* (22, 6, 27) {real, imag} */,
  {32'hbf155776, 32'h3e845686} /* (22, 6, 26) {real, imag} */,
  {32'hbe8cae06, 32'hbc558d18} /* (22, 6, 25) {real, imag} */,
  {32'h3e827f05, 32'hbee3b4f2} /* (22, 6, 24) {real, imag} */,
  {32'hbedec086, 32'h3dc27e68} /* (22, 6, 23) {real, imag} */,
  {32'hbe1d2bd2, 32'h3f00d7e6} /* (22, 6, 22) {real, imag} */,
  {32'hbc8a1560, 32'hbe4fb4f0} /* (22, 6, 21) {real, imag} */,
  {32'hbe031127, 32'hbe761efd} /* (22, 6, 20) {real, imag} */,
  {32'hbd8ff1e4, 32'h3ec6abe1} /* (22, 6, 19) {real, imag} */,
  {32'hbdaa1d7a, 32'h3e1ca880} /* (22, 6, 18) {real, imag} */,
  {32'h3d389124, 32'hbe70202a} /* (22, 6, 17) {real, imag} */,
  {32'hbe1e9fb3, 32'h3da735e0} /* (22, 6, 16) {real, imag} */,
  {32'hbe3d2b0a, 32'h3e62332f} /* (22, 6, 15) {real, imag} */,
  {32'hbe7934d4, 32'h3ea1719e} /* (22, 6, 14) {real, imag} */,
  {32'h3e88d128, 32'h3d96f279} /* (22, 6, 13) {real, imag} */,
  {32'h3e8f0d5f, 32'h3eeb3741} /* (22, 6, 12) {real, imag} */,
  {32'hbea37747, 32'h3e4a14f6} /* (22, 6, 11) {real, imag} */,
  {32'hbf1c00b5, 32'h3cc3dbf0} /* (22, 6, 10) {real, imag} */,
  {32'h3e0b95f7, 32'hbdacae22} /* (22, 6, 9) {real, imag} */,
  {32'h3e348b03, 32'hbe9f0ce4} /* (22, 6, 8) {real, imag} */,
  {32'hbef03075, 32'hbe735a2e} /* (22, 6, 7) {real, imag} */,
  {32'hbe285a07, 32'hbf023415} /* (22, 6, 6) {real, imag} */,
  {32'hbf48a185, 32'h3e7bd728} /* (22, 6, 5) {real, imag} */,
  {32'h3e845c35, 32'h3d2dbb34} /* (22, 6, 4) {real, imag} */,
  {32'h3f3e9294, 32'hbf8208b2} /* (22, 6, 3) {real, imag} */,
  {32'hbf1c8e86, 32'h3db8636c} /* (22, 6, 2) {real, imag} */,
  {32'h3ec6bbf4, 32'h3e59f576} /* (22, 6, 1) {real, imag} */,
  {32'h3cd057f0, 32'h3eae6960} /* (22, 6, 0) {real, imag} */,
  {32'h40421804, 32'h3f4d22ba} /* (22, 5, 31) {real, imag} */,
  {32'hbff955d3, 32'hbef0a908} /* (22, 5, 30) {real, imag} */,
  {32'hbd921dbf, 32'hbe332cc4} /* (22, 5, 29) {real, imag} */,
  {32'hbef7b875, 32'hbdf0f3e8} /* (22, 5, 28) {real, imag} */,
  {32'hbf981e7b, 32'hbdca6d3a} /* (22, 5, 27) {real, imag} */,
  {32'hbd53cf8a, 32'h3f348a86} /* (22, 5, 26) {real, imag} */,
  {32'hbe39983c, 32'hbe4ead34} /* (22, 5, 25) {real, imag} */,
  {32'hbec9f456, 32'h3d5bddd0} /* (22, 5, 24) {real, imag} */,
  {32'h3e894d30, 32'hbf0040d8} /* (22, 5, 23) {real, imag} */,
  {32'hbf2aa39b, 32'h3e6bd3de} /* (22, 5, 22) {real, imag} */,
  {32'hbda1cc62, 32'h3d771508} /* (22, 5, 21) {real, imag} */,
  {32'h3e863ef1, 32'hbf012952} /* (22, 5, 20) {real, imag} */,
  {32'h3e345590, 32'hbe277a51} /* (22, 5, 19) {real, imag} */,
  {32'h3ec05570, 32'h3c010700} /* (22, 5, 18) {real, imag} */,
  {32'h3d4bfbe1, 32'hbdaad196} /* (22, 5, 17) {real, imag} */,
  {32'hbeea741c, 32'hbe943956} /* (22, 5, 16) {real, imag} */,
  {32'hbd9ba87c, 32'h3e4240c8} /* (22, 5, 15) {real, imag} */,
  {32'h3eb1207a, 32'hbe404c78} /* (22, 5, 14) {real, imag} */,
  {32'h3ece23aa, 32'hbe2b34ff} /* (22, 5, 13) {real, imag} */,
  {32'hbed6c29c, 32'hbe58ed0f} /* (22, 5, 12) {real, imag} */,
  {32'hbe2da160, 32'hbf016d7c} /* (22, 5, 11) {real, imag} */,
  {32'hbe291a7e, 32'hbeb4a42a} /* (22, 5, 10) {real, imag} */,
  {32'h3e45c1b3, 32'hbc2eb738} /* (22, 5, 9) {real, imag} */,
  {32'hbd348140, 32'hbbd47800} /* (22, 5, 8) {real, imag} */,
  {32'h3e9ca0d2, 32'hbd15b224} /* (22, 5, 7) {real, imag} */,
  {32'h3ec3ae9a, 32'h3d89e92a} /* (22, 5, 6) {real, imag} */,
  {32'hbe98e420, 32'hbf3a9662} /* (22, 5, 5) {real, imag} */,
  {32'hbea60f44, 32'h3fbf19b2} /* (22, 5, 4) {real, imag} */,
  {32'hbda7484b, 32'hbe2225be} /* (22, 5, 3) {real, imag} */,
  {32'h3e577095, 32'hbfa206a0} /* (22, 5, 2) {real, imag} */,
  {32'h4043ee42, 32'h403cd575} /* (22, 5, 1) {real, imag} */,
  {32'h400e3266, 32'h3fa1a283} /* (22, 5, 0) {real, imag} */,
  {32'hbf8ac486, 32'hc04aa144} /* (22, 4, 31) {real, imag} */,
  {32'h402cce27, 32'h40258a7e} /* (22, 4, 30) {real, imag} */,
  {32'hbf56fa5a, 32'h3e4f89b1} /* (22, 4, 29) {real, imag} */,
  {32'hbf27e602, 32'hbe431b48} /* (22, 4, 28) {real, imag} */,
  {32'h3ecc0331, 32'hbebe7112} /* (22, 4, 27) {real, imag} */,
  {32'h3e1b4b7e, 32'hbea30b76} /* (22, 4, 26) {real, imag} */,
  {32'h3e9272a0, 32'hbe24770b} /* (22, 4, 25) {real, imag} */,
  {32'h3f142800, 32'h3ed4c1ee} /* (22, 4, 24) {real, imag} */,
  {32'hbe99c65e, 32'hbeead1b3} /* (22, 4, 23) {real, imag} */,
  {32'hbe056abc, 32'h3e3277ee} /* (22, 4, 22) {real, imag} */,
  {32'hbea99460, 32'h3eb26464} /* (22, 4, 21) {real, imag} */,
  {32'h3cf9ade8, 32'hbddf8728} /* (22, 4, 20) {real, imag} */,
  {32'hbca40991, 32'h3ddc9c43} /* (22, 4, 19) {real, imag} */,
  {32'h3ef568e6, 32'hbe79c769} /* (22, 4, 18) {real, imag} */,
  {32'hbb212eb8, 32'hbc9a0f30} /* (22, 4, 17) {real, imag} */,
  {32'hbdf0b3f8, 32'h3d999a83} /* (22, 4, 16) {real, imag} */,
  {32'hbe0239bd, 32'h3da717d0} /* (22, 4, 15) {real, imag} */,
  {32'h3ece3398, 32'h3de42fb5} /* (22, 4, 14) {real, imag} */,
  {32'hbe7d0c50, 32'h3e4b30e0} /* (22, 4, 13) {real, imag} */,
  {32'hbe462c98, 32'hbf1dd60a} /* (22, 4, 12) {real, imag} */,
  {32'h3eb88ff7, 32'h3ef30493} /* (22, 4, 11) {real, imag} */,
  {32'hbcd12900, 32'h3efdd395} /* (22, 4, 10) {real, imag} */,
  {32'h3e6cd5c7, 32'hbe4956e1} /* (22, 4, 9) {real, imag} */,
  {32'h3f0529ee, 32'hbe2c7a72} /* (22, 4, 8) {real, imag} */,
  {32'hbe1adeb2, 32'hbc5728f0} /* (22, 4, 7) {real, imag} */,
  {32'hbef1bdc2, 32'hbdb0a72c} /* (22, 4, 6) {real, imag} */,
  {32'h3daf07ec, 32'h3d8149b0} /* (22, 4, 5) {real, imag} */,
  {32'h3f0fd021, 32'hbf9d48d5} /* (22, 4, 4) {real, imag} */,
  {32'h3ea73f7a, 32'hbe87b3df} /* (22, 4, 3) {real, imag} */,
  {32'h4059f190, 32'h4004598b} /* (22, 4, 2) {real, imag} */,
  {32'hc068461e, 32'hbf94eb4a} /* (22, 4, 1) {real, imag} */,
  {32'hc02687b2, 32'h3f523d72} /* (22, 4, 0) {real, imag} */,
  {32'h40928d49, 32'hc00e305d} /* (22, 3, 31) {real, imag} */,
  {32'hc03e7f5b, 32'h405b40fa} /* (22, 3, 30) {real, imag} */,
  {32'hbda16f84, 32'hbe0ddfa6} /* (22, 3, 29) {real, imag} */,
  {32'hbfeafca8, 32'hbf7a9d50} /* (22, 3, 28) {real, imag} */,
  {32'h3f299642, 32'h3e7385f4} /* (22, 3, 27) {real, imag} */,
  {32'h3e13ddb4, 32'hbe0605e2} /* (22, 3, 26) {real, imag} */,
  {32'h3e931b8f, 32'hbf19069b} /* (22, 3, 25) {real, imag} */,
  {32'h3f494744, 32'h3e434ee3} /* (22, 3, 24) {real, imag} */,
  {32'hbdf14d3c, 32'hbef7f472} /* (22, 3, 23) {real, imag} */,
  {32'hbec0f862, 32'hbeb9b9e8} /* (22, 3, 22) {real, imag} */,
  {32'hbbfd4e98, 32'h3e5f7e68} /* (22, 3, 21) {real, imag} */,
  {32'h3eacb868, 32'hbea4bee4} /* (22, 3, 20) {real, imag} */,
  {32'h3e9e469c, 32'h3e97baa7} /* (22, 3, 19) {real, imag} */,
  {32'h3ec84e6e, 32'h3daa3cf0} /* (22, 3, 18) {real, imag} */,
  {32'hbe3893e3, 32'h3e124c06} /* (22, 3, 17) {real, imag} */,
  {32'h3e252e0e, 32'hbe3c638a} /* (22, 3, 16) {real, imag} */,
  {32'hbead7de3, 32'hbd795bc0} /* (22, 3, 15) {real, imag} */,
  {32'hbea88d5a, 32'h3d56ae3c} /* (22, 3, 14) {real, imag} */,
  {32'h3dd60d7b, 32'h3ea3a702} /* (22, 3, 13) {real, imag} */,
  {32'h3f20bde2, 32'hbe158254} /* (22, 3, 12) {real, imag} */,
  {32'hbe8190a6, 32'h3d60d310} /* (22, 3, 11) {real, imag} */,
  {32'hbe98ca58, 32'h3f2b1016} /* (22, 3, 10) {real, imag} */,
  {32'hbeac692c, 32'hbf0d3c98} /* (22, 3, 9) {real, imag} */,
  {32'hbed8a89a, 32'h3ef847e9} /* (22, 3, 8) {real, imag} */,
  {32'h3e6f066d, 32'hbe80565c} /* (22, 3, 7) {real, imag} */,
  {32'h3ef16600, 32'h3dc16bda} /* (22, 3, 6) {real, imag} */,
  {32'hbf3d52a3, 32'hbe61d01e} /* (22, 3, 5) {real, imag} */,
  {32'h3f5c5fce, 32'hbff481d2} /* (22, 3, 4) {real, imag} */,
  {32'h3db09af0, 32'hbf26b081} /* (22, 3, 3) {real, imag} */,
  {32'hbf0e3b76, 32'h408959f0} /* (22, 3, 2) {real, imag} */,
  {32'hc084234c, 32'hc02bcd6e} /* (22, 3, 1) {real, imag} */,
  {32'h40050126, 32'hbc845a60} /* (22, 3, 0) {real, imag} */,
  {32'h421cedcb, 32'h3f999956} /* (22, 2, 31) {real, imag} */,
  {32'hc18ac138, 32'h40d04f88} /* (22, 2, 30) {real, imag} */,
  {32'hbe05e878, 32'hbf31d48c} /* (22, 2, 29) {real, imag} */,
  {32'h3f8fa701, 32'hc0443e52} /* (22, 2, 28) {real, imag} */,
  {32'hbfde244b, 32'h3f69443b} /* (22, 2, 27) {real, imag} */,
  {32'hbf9428ad, 32'hbe343f0c} /* (22, 2, 26) {real, imag} */,
  {32'h3f623c04, 32'hbee20bc2} /* (22, 2, 25) {real, imag} */,
  {32'hbeabd461, 32'h3e8ba84c} /* (22, 2, 24) {real, imag} */,
  {32'hbe886ef7, 32'hbe858c64} /* (22, 2, 23) {real, imag} */,
  {32'hbdde7c60, 32'h3eacb5f8} /* (22, 2, 22) {real, imag} */,
  {32'h3d7429b4, 32'h3e906ed8} /* (22, 2, 21) {real, imag} */,
  {32'h3ea646c0, 32'h3ea78714} /* (22, 2, 20) {real, imag} */,
  {32'hbf126ad2, 32'h3ee30a28} /* (22, 2, 19) {real, imag} */,
  {32'hbdd2c0c6, 32'h3edf3a92} /* (22, 2, 18) {real, imag} */,
  {32'h37368000, 32'hbe5d188a} /* (22, 2, 17) {real, imag} */,
  {32'h3d216b7e, 32'hbc01b444} /* (22, 2, 16) {real, imag} */,
  {32'hbd1b4978, 32'h3db2ef32} /* (22, 2, 15) {real, imag} */,
  {32'h3edc3672, 32'h3d9cd974} /* (22, 2, 14) {real, imag} */,
  {32'h3ebd8a8e, 32'h3e3a691a} /* (22, 2, 13) {real, imag} */,
  {32'hbedb1b2a, 32'hbf07bac5} /* (22, 2, 12) {real, imag} */,
  {32'hbe12b6b3, 32'hbf296855} /* (22, 2, 11) {real, imag} */,
  {32'h3ed9f63e, 32'h3f3283f3} /* (22, 2, 10) {real, imag} */,
  {32'h3e09fac1, 32'hbd48fcfc} /* (22, 2, 9) {real, imag} */,
  {32'hbf2b67ca, 32'hbf105571} /* (22, 2, 8) {real, imag} */,
  {32'h3cdf1538, 32'hbdc9f334} /* (22, 2, 7) {real, imag} */,
  {32'hbe62859a, 32'h3edce178} /* (22, 2, 6) {real, imag} */,
  {32'hc0234c60, 32'hc0103032} /* (22, 2, 5) {real, imag} */,
  {32'h40403adf, 32'h400b6ee7} /* (22, 2, 4) {real, imag} */,
  {32'h3e26fc6c, 32'hbfb6204b} /* (22, 2, 3) {real, imag} */,
  {32'hc14d8aca, 32'h40361d12} /* (22, 2, 2) {real, imag} */,
  {32'h41b39153, 32'hc0262180} /* (22, 2, 1) {real, imag} */,
  {32'h419f47b8, 32'h4089dc98} /* (22, 2, 0) {real, imag} */,
  {32'hc255cc2b, 32'h41659299} /* (22, 1, 31) {real, imag} */,
  {32'h41649f0c, 32'h402a096e} /* (22, 1, 30) {real, imag} */,
  {32'h3f5c9d48, 32'hc0092b77} /* (22, 1, 29) {real, imag} */,
  {32'hc08cdf8f, 32'hc002e392} /* (22, 1, 28) {real, imag} */,
  {32'h408f695e, 32'hbe9fe67f} /* (22, 1, 27) {real, imag} */,
  {32'h3f56bc25, 32'hbdd42674} /* (22, 1, 26) {real, imag} */,
  {32'hbf0ec39c, 32'hbec895c4} /* (22, 1, 25) {real, imag} */,
  {32'h3ef9f2c4, 32'hbedd731e} /* (22, 1, 24) {real, imag} */,
  {32'h3ef1c55c, 32'hbf4fefc6} /* (22, 1, 23) {real, imag} */,
  {32'h3eaeb0bd, 32'hbe8304c3} /* (22, 1, 22) {real, imag} */,
  {32'h3e7e650b, 32'h3e791436} /* (22, 1, 21) {real, imag} */,
  {32'h3e4dcde5, 32'hbe5a1ffa} /* (22, 1, 20) {real, imag} */,
  {32'h3da08910, 32'hbe51ebb4} /* (22, 1, 19) {real, imag} */,
  {32'h3e1ab3ec, 32'h3e89683a} /* (22, 1, 18) {real, imag} */,
  {32'hbe0e4226, 32'h3df2ac55} /* (22, 1, 17) {real, imag} */,
  {32'h3e2d62ce, 32'hbe18e40c} /* (22, 1, 16) {real, imag} */,
  {32'hbe10964e, 32'h3ea3f154} /* (22, 1, 15) {real, imag} */,
  {32'h3c543330, 32'h3ee28776} /* (22, 1, 14) {real, imag} */,
  {32'hbeeed590, 32'hbe406d60} /* (22, 1, 13) {real, imag} */,
  {32'h3e98f52a, 32'h3e10004c} /* (22, 1, 12) {real, imag} */,
  {32'h3f03ab84, 32'h3e4cfb0d} /* (22, 1, 11) {real, imag} */,
  {32'hbeb9412a, 32'h3ecf3ee7} /* (22, 1, 10) {real, imag} */,
  {32'h3e4c8ed1, 32'hbec5d99d} /* (22, 1, 9) {real, imag} */,
  {32'h3e19a629, 32'h3fbcd0a4} /* (22, 1, 8) {real, imag} */,
  {32'hbec586a9, 32'hbfadcd14} /* (22, 1, 7) {real, imag} */,
  {32'hbe01a2c4, 32'hbe4959ba} /* (22, 1, 6) {real, imag} */,
  {32'h40087c97, 32'h3fe006c1} /* (22, 1, 5) {real, imag} */,
  {32'hbfd493e2, 32'hc00f9744} /* (22, 1, 4) {real, imag} */,
  {32'h40056b01, 32'h3f410cc4} /* (22, 1, 3) {real, imag} */,
  {32'h41900e9d, 32'h418e30d7} /* (22, 1, 2) {real, imag} */,
  {32'hc2988d2b, 32'hc223f327} /* (22, 1, 1) {real, imag} */,
  {32'hc286879a, 32'hc1171b6c} /* (22, 1, 0) {real, imag} */,
  {32'hc2403ee8, 32'h42195acc} /* (22, 0, 31) {real, imag} */,
  {32'h40b32310, 32'hc10b3bc4} /* (22, 0, 30) {real, imag} */,
  {32'h3bbb6500, 32'hbeb52c96} /* (22, 0, 29) {real, imag} */,
  {32'h3f849fdf, 32'hc0090194} /* (22, 0, 28) {real, imag} */,
  {32'h401772d6, 32'h3d7d81d8} /* (22, 0, 27) {real, imag} */,
  {32'hbec6c26a, 32'hbeed4910} /* (22, 0, 26) {real, imag} */,
  {32'h3f32a2ce, 32'hbd025010} /* (22, 0, 25) {real, imag} */,
  {32'h3d9d9b94, 32'hbf88ff76} /* (22, 0, 24) {real, imag} */,
  {32'h3ee0a356, 32'hbe204a88} /* (22, 0, 23) {real, imag} */,
  {32'h3e973167, 32'h3e8021ce} /* (22, 0, 22) {real, imag} */,
  {32'h3e4919b8, 32'hbf03c30f} /* (22, 0, 21) {real, imag} */,
  {32'hbe6850fd, 32'h3dfce99f} /* (22, 0, 20) {real, imag} */,
  {32'h3d7bcaf1, 32'hbe6eb7ee} /* (22, 0, 19) {real, imag} */,
  {32'hbed193f8, 32'hbda7ad29} /* (22, 0, 18) {real, imag} */,
  {32'h3d85fbec, 32'h3e893e9a} /* (22, 0, 17) {real, imag} */,
  {32'h3db29ff8, 32'h00000000} /* (22, 0, 16) {real, imag} */,
  {32'h3d85fbec, 32'hbe893e9a} /* (22, 0, 15) {real, imag} */,
  {32'hbed193f8, 32'h3da7ad29} /* (22, 0, 14) {real, imag} */,
  {32'h3d7bcaf1, 32'h3e6eb7ee} /* (22, 0, 13) {real, imag} */,
  {32'hbe6850fd, 32'hbdfce99f} /* (22, 0, 12) {real, imag} */,
  {32'h3e4919b8, 32'h3f03c30f} /* (22, 0, 11) {real, imag} */,
  {32'h3e973167, 32'hbe8021ce} /* (22, 0, 10) {real, imag} */,
  {32'h3ee0a356, 32'h3e204a88} /* (22, 0, 9) {real, imag} */,
  {32'h3d9d9b94, 32'h3f88ff76} /* (22, 0, 8) {real, imag} */,
  {32'h3f32a2ce, 32'h3d025010} /* (22, 0, 7) {real, imag} */,
  {32'hbec6c26a, 32'h3eed4910} /* (22, 0, 6) {real, imag} */,
  {32'h401772d6, 32'hbd7d81d8} /* (22, 0, 5) {real, imag} */,
  {32'h3f849fdf, 32'h40090194} /* (22, 0, 4) {real, imag} */,
  {32'h3bbb6500, 32'h3eb52c96} /* (22, 0, 3) {real, imag} */,
  {32'h40b32310, 32'h410b3bc4} /* (22, 0, 2) {real, imag} */,
  {32'hc2403ee8, 32'hc2195acc} /* (22, 0, 1) {real, imag} */,
  {32'hc29598fc, 32'h00000000} /* (22, 0, 0) {real, imag} */,
  {32'hc29ee7a3, 32'h422a4da7} /* (21, 31, 31) {real, imag} */,
  {32'h418f4c17, 32'hc1904db4} /* (21, 31, 30) {real, imag} */,
  {32'h3fe163fa, 32'hbf2846d6} /* (21, 31, 29) {real, imag} */,
  {32'hbf467fe8, 32'h401162c8} /* (21, 31, 28) {real, imag} */,
  {32'h40054e6c, 32'hc000f509} /* (21, 31, 27) {real, imag} */,
  {32'hbe95ca7d, 32'h3e57d8f4} /* (21, 31, 26) {real, imag} */,
  {32'h3de1fdc8, 32'h3f4e4f79} /* (21, 31, 25) {real, imag} */,
  {32'h3e577b58, 32'hbfb4bb8a} /* (21, 31, 24) {real, imag} */,
  {32'h3f98a2bd, 32'hbe9d4159} /* (21, 31, 23) {real, imag} */,
  {32'hbef27c7c, 32'h3de7abec} /* (21, 31, 22) {real, imag} */,
  {32'h3e43dd87, 32'hbf559e6a} /* (21, 31, 21) {real, imag} */,
  {32'h3dcd9fd2, 32'hbf2121f0} /* (21, 31, 20) {real, imag} */,
  {32'hbd07e6e0, 32'h3efb8434} /* (21, 31, 19) {real, imag} */,
  {32'hbe90b2e6, 32'hbe9142ca} /* (21, 31, 18) {real, imag} */,
  {32'hbe07d492, 32'h3e6822ca} /* (21, 31, 17) {real, imag} */,
  {32'hbcd8c234, 32'h3e4da5c6} /* (21, 31, 16) {real, imag} */,
  {32'h3f063785, 32'hbd05abc0} /* (21, 31, 15) {real, imag} */,
  {32'h3e0bc460, 32'hbe221341} /* (21, 31, 14) {real, imag} */,
  {32'hbd34d968, 32'h3eaac105} /* (21, 31, 13) {real, imag} */,
  {32'h3ebec4fc, 32'hbdb892db} /* (21, 31, 12) {real, imag} */,
  {32'h3f7002f3, 32'hbe528a8b} /* (21, 31, 11) {real, imag} */,
  {32'h3f7fed07, 32'h3dd4a3f8} /* (21, 31, 10) {real, imag} */,
  {32'h3f287ea4, 32'h3ef6d706} /* (21, 31, 9) {real, imag} */,
  {32'h3dca2924, 32'h3f080721} /* (21, 31, 8) {real, imag} */,
  {32'h3e3c3e07, 32'h3f166f83} /* (21, 31, 7) {real, imag} */,
  {32'h3e934a2f, 32'h3f60eaff} /* (21, 31, 6) {real, imag} */,
  {32'h40876ed6, 32'h3ee832f8} /* (21, 31, 5) {real, imag} */,
  {32'hc05c6d9a, 32'h4049a8ce} /* (21, 31, 4) {real, imag} */,
  {32'h3df047d0, 32'h3fe920f2} /* (21, 31, 3) {real, imag} */,
  {32'h417436ba, 32'hbf2b5ccb} /* (21, 31, 2) {real, imag} */,
  {32'hc2615558, 32'hc173fda5} /* (21, 31, 1) {real, imag} */,
  {32'hc28a002c, 32'h412856a6} /* (21, 31, 0) {real, imag} */,
  {32'h41c3ca46, 32'h40546b7e} /* (21, 30, 31) {real, imag} */,
  {32'hc1492148, 32'hc03bd477} /* (21, 30, 30) {real, imag} */,
  {32'h3dd090d0, 32'h3f558fc4} /* (21, 30, 29) {real, imag} */,
  {32'h40442db8, 32'hbf283ce5} /* (21, 30, 28) {real, imag} */,
  {32'hc02dfe11, 32'h3fe9ac94} /* (21, 30, 27) {real, imag} */,
  {32'h3dfb8667, 32'hbeb2b07d} /* (21, 30, 26) {real, imag} */,
  {32'h3d68248e, 32'h3eb86ddf} /* (21, 30, 25) {real, imag} */,
  {32'hbef29192, 32'h3f764f98} /* (21, 30, 24) {real, imag} */,
  {32'h3ee83a34, 32'h3e26cceb} /* (21, 30, 23) {real, imag} */,
  {32'h3eb76366, 32'h3dfcbe30} /* (21, 30, 22) {real, imag} */,
  {32'h3c9ecd74, 32'h3f119470} /* (21, 30, 21) {real, imag} */,
  {32'h3e85be9e, 32'hbd98c694} /* (21, 30, 20) {real, imag} */,
  {32'hbe1167ec, 32'hbea0187a} /* (21, 30, 19) {real, imag} */,
  {32'h3e62beec, 32'h3f415f93} /* (21, 30, 18) {real, imag} */,
  {32'hbdd3f85c, 32'hbe34ccda} /* (21, 30, 17) {real, imag} */,
  {32'hbe80017b, 32'hbd373352} /* (21, 30, 16) {real, imag} */,
  {32'h3d0e6650, 32'h3ec1acdc} /* (21, 30, 15) {real, imag} */,
  {32'hbf1d12a0, 32'hbe4620c8} /* (21, 30, 14) {real, imag} */,
  {32'hbd97e177, 32'h3e061f04} /* (21, 30, 13) {real, imag} */,
  {32'h3e93a82e, 32'h3e149d28} /* (21, 30, 12) {real, imag} */,
  {32'h3d3ad3fc, 32'hbe1abe48} /* (21, 30, 11) {real, imag} */,
  {32'hbee0899b, 32'h3c00c098} /* (21, 30, 10) {real, imag} */,
  {32'hbeed993a, 32'hbda33836} /* (21, 30, 9) {real, imag} */,
  {32'hbf790397, 32'hbfbaeb5f} /* (21, 30, 8) {real, imag} */,
  {32'h3f40fc76, 32'h3f1a725e} /* (21, 30, 7) {real, imag} */,
  {32'hbd3db5d8, 32'hbee74c88} /* (21, 30, 6) {real, imag} */,
  {32'hbfa76feb, 32'hbf6ac712} /* (21, 30, 5) {real, imag} */,
  {32'h3e232870, 32'h3ffe464c} /* (21, 30, 4) {real, imag} */,
  {32'hbca50508, 32'hbe6d6e25} /* (21, 30, 3) {real, imag} */,
  {32'hc1943477, 32'hc0e680f3} /* (21, 30, 2) {real, imag} */,
  {32'h42246bad, 32'hbf075c0a} /* (21, 30, 1) {real, imag} */,
  {32'h41a4705c, 32'hc0873b9c} /* (21, 30, 0) {real, imag} */,
  {32'hc088adde, 32'h4037548c} /* (21, 29, 31) {real, imag} */,
  {32'hbe852833, 32'hc06586ac} /* (21, 29, 30) {real, imag} */,
  {32'h3fcac748, 32'hbe9a2c5a} /* (21, 29, 29) {real, imag} */,
  {32'h3fb12b07, 32'h3fb24670} /* (21, 29, 28) {real, imag} */,
  {32'hbe8b83c6, 32'h3de39be2} /* (21, 29, 27) {real, imag} */,
  {32'hbd249684, 32'h3d9a418a} /* (21, 29, 26) {real, imag} */,
  {32'h3f1dc7dc, 32'h3eb52d3f} /* (21, 29, 25) {real, imag} */,
  {32'hbf03c27e, 32'hbed92208} /* (21, 29, 24) {real, imag} */,
  {32'hbf5a58ce, 32'hbd6c76c4} /* (21, 29, 23) {real, imag} */,
  {32'h3e51a864, 32'hbebd6069} /* (21, 29, 22) {real, imag} */,
  {32'hbdee3a9a, 32'hbe3f8c20} /* (21, 29, 21) {real, imag} */,
  {32'hbd373850, 32'hbeab0e13} /* (21, 29, 20) {real, imag} */,
  {32'h3dcfdacc, 32'h3ca3a002} /* (21, 29, 19) {real, imag} */,
  {32'hbc7c3aa0, 32'hbec73263} /* (21, 29, 18) {real, imag} */,
  {32'h3e9a784b, 32'hbc865550} /* (21, 29, 17) {real, imag} */,
  {32'h3f0005d1, 32'hbdaf0124} /* (21, 29, 16) {real, imag} */,
  {32'h3cf6f1b8, 32'hbd28d270} /* (21, 29, 15) {real, imag} */,
  {32'hbe61615e, 32'h3ec73e02} /* (21, 29, 14) {real, imag} */,
  {32'h3efcfb7d, 32'h3e9d4fff} /* (21, 29, 13) {real, imag} */,
  {32'h3f0a5966, 32'hbf15f017} /* (21, 29, 12) {real, imag} */,
  {32'h3eb1061a, 32'hbf200dd0} /* (21, 29, 11) {real, imag} */,
  {32'hbe6fc6db, 32'h3f4b9a10} /* (21, 29, 10) {real, imag} */,
  {32'hbd152e9c, 32'h3f2d83df} /* (21, 29, 9) {real, imag} */,
  {32'h3f36d850, 32'hbe5d6283} /* (21, 29, 8) {real, imag} */,
  {32'hbf53e032, 32'h3e1bda4a} /* (21, 29, 7) {real, imag} */,
  {32'h3e8e44fc, 32'h3f5a7e81} /* (21, 29, 6) {real, imag} */,
  {32'h3effad59, 32'h3df20d54} /* (21, 29, 5) {real, imag} */,
  {32'hbfc47536, 32'h3f9809de} /* (21, 29, 4) {real, imag} */,
  {32'hbe9a8dcb, 32'hbdf924b9} /* (21, 29, 3) {real, imag} */,
  {32'hc04f5563, 32'hc045f0e9} /* (21, 29, 2) {real, imag} */,
  {32'h4093f214, 32'h402111e1} /* (21, 29, 1) {real, imag} */,
  {32'h3fc0fea0, 32'hbeb207d2} /* (21, 29, 0) {real, imag} */,
  {32'hc08e25c0, 32'h3fec4de8} /* (21, 28, 31) {real, imag} */,
  {32'h40736fd0, 32'hbff0705c} /* (21, 28, 30) {real, imag} */,
  {32'hbdeaabe0, 32'h3f98af4a} /* (21, 28, 29) {real, imag} */,
  {32'h3f4f7a63, 32'h3f8587ad} /* (21, 28, 28) {real, imag} */,
  {32'h3f3cfe58, 32'hbe90531e} /* (21, 28, 27) {real, imag} */,
  {32'hbd0863c8, 32'hbd182d08} /* (21, 28, 26) {real, imag} */,
  {32'hbf10d2e4, 32'hbe1e8fe7} /* (21, 28, 25) {real, imag} */,
  {32'h3f319a4d, 32'hbebb8a99} /* (21, 28, 24) {real, imag} */,
  {32'h3dba87e8, 32'hbd614bb4} /* (21, 28, 23) {real, imag} */,
  {32'h3e1cdff2, 32'h3e0616f5} /* (21, 28, 22) {real, imag} */,
  {32'h3f18bac7, 32'hbe079407} /* (21, 28, 21) {real, imag} */,
  {32'hbe639be7, 32'hbd375a0f} /* (21, 28, 20) {real, imag} */,
  {32'hbe8e3c3a, 32'h3f315bb6} /* (21, 28, 19) {real, imag} */,
  {32'h3baaf9e0, 32'h3e81ceea} /* (21, 28, 18) {real, imag} */,
  {32'h3dca15a4, 32'h3bc53428} /* (21, 28, 17) {real, imag} */,
  {32'hbe3700a2, 32'hbd5dcf24} /* (21, 28, 16) {real, imag} */,
  {32'h3d31349c, 32'hbdd29ae4} /* (21, 28, 15) {real, imag} */,
  {32'h3f0a62ac, 32'hbee02be6} /* (21, 28, 14) {real, imag} */,
  {32'hbe41e5b0, 32'hbf1a8f9a} /* (21, 28, 13) {real, imag} */,
  {32'h3f0a8a6d, 32'hbf0f7464} /* (21, 28, 12) {real, imag} */,
  {32'hbf0c8005, 32'h3e855968} /* (21, 28, 11) {real, imag} */,
  {32'hbe957701, 32'hbd9548d7} /* (21, 28, 10) {real, imag} */,
  {32'hbe950669, 32'h3e063eb5} /* (21, 28, 9) {real, imag} */,
  {32'h3ecf046c, 32'hbe753f05} /* (21, 28, 8) {real, imag} */,
  {32'h3e96f032, 32'hbf1d6c32} /* (21, 28, 7) {real, imag} */,
  {32'h3ea04934, 32'h3f2774f2} /* (21, 28, 6) {real, imag} */,
  {32'h3ddffa2e, 32'h3f47ef34} /* (21, 28, 5) {real, imag} */,
  {32'hbf126db6, 32'hbf3739ac} /* (21, 28, 4) {real, imag} */,
  {32'h3e3570c2, 32'hbc145e20} /* (21, 28, 3) {real, imag} */,
  {32'h4041bff3, 32'hbfe864da} /* (21, 28, 2) {real, imag} */,
  {32'hbf76f992, 32'h4059fc9f} /* (21, 28, 1) {real, imag} */,
  {32'hc003df29, 32'hbfa80a95} /* (21, 28, 0) {real, imag} */,
  {32'h4001da38, 32'hc00106c8} /* (21, 27, 31) {real, imag} */,
  {32'hbeff4f69, 32'h3fbca04f} /* (21, 27, 30) {real, imag} */,
  {32'h3e923773, 32'hbe94306c} /* (21, 27, 29) {real, imag} */,
  {32'hbee3baf0, 32'hbf14d418} /* (21, 27, 28) {real, imag} */,
  {32'hbf139dd8, 32'h3f01563d} /* (21, 27, 27) {real, imag} */,
  {32'h3e79787c, 32'h3ea36fe8} /* (21, 27, 26) {real, imag} */,
  {32'h3f874d8c, 32'hbecd9639} /* (21, 27, 25) {real, imag} */,
  {32'hbe4da84b, 32'h3dc12ed0} /* (21, 27, 24) {real, imag} */,
  {32'h3e7e9a15, 32'h3efa41a2} /* (21, 27, 23) {real, imag} */,
  {32'h3e867b40, 32'hbe47d274} /* (21, 27, 22) {real, imag} */,
  {32'hbe8f9e70, 32'h3f12d404} /* (21, 27, 21) {real, imag} */,
  {32'hbe2a43d0, 32'h3e840ba6} /* (21, 27, 20) {real, imag} */,
  {32'h3e262d48, 32'h3caa5670} /* (21, 27, 19) {real, imag} */,
  {32'hbe933b91, 32'h3da13344} /* (21, 27, 18) {real, imag} */,
  {32'hbe4ee78c, 32'hbb369a00} /* (21, 27, 17) {real, imag} */,
  {32'hbe2c0092, 32'hbdcb97be} /* (21, 27, 16) {real, imag} */,
  {32'h3e2b4179, 32'h3e9c60db} /* (21, 27, 15) {real, imag} */,
  {32'hbd449b52, 32'hbde0551e} /* (21, 27, 14) {real, imag} */,
  {32'hbd8e23e8, 32'hbd6db4dc} /* (21, 27, 13) {real, imag} */,
  {32'h3ea5506a, 32'hbe82bb36} /* (21, 27, 12) {real, imag} */,
  {32'hbc50e568, 32'h3e57b5ce} /* (21, 27, 11) {real, imag} */,
  {32'hbe3d7857, 32'h3ac04700} /* (21, 27, 10) {real, imag} */,
  {32'h3d75a488, 32'hbe532f05} /* (21, 27, 9) {real, imag} */,
  {32'hbe2a8644, 32'hbe247504} /* (21, 27, 8) {real, imag} */,
  {32'h3e8d6142, 32'hbd28dfde} /* (21, 27, 7) {real, imag} */,
  {32'hbf59b72e, 32'hbdb7449e} /* (21, 27, 6) {real, imag} */,
  {32'hbf738dee, 32'h3dc7c98c} /* (21, 27, 5) {real, imag} */,
  {32'h3f15423c, 32'h3e62c888} /* (21, 27, 4) {real, imag} */,
  {32'h3d674b80, 32'hbecf53e4} /* (21, 27, 3) {real, imag} */,
  {32'hbf83cf70, 32'h3ed3c5f0} /* (21, 27, 2) {real, imag} */,
  {32'h403d67e2, 32'hbee18323} /* (21, 27, 1) {real, imag} */,
  {32'h3f962774, 32'hc015cd98} /* (21, 27, 0) {real, imag} */,
  {32'hbdd0f7c8, 32'hbeac6f77} /* (21, 26, 31) {real, imag} */,
  {32'h3e0e3884, 32'hbf383a26} /* (21, 26, 30) {real, imag} */,
  {32'h3f1b20b3, 32'h3f250a81} /* (21, 26, 29) {real, imag} */,
  {32'hbe0c1600, 32'hbd9647d1} /* (21, 26, 28) {real, imag} */,
  {32'hbf387360, 32'hbe3ee95d} /* (21, 26, 27) {real, imag} */,
  {32'hbed0a914, 32'h3f10b2ee} /* (21, 26, 26) {real, imag} */,
  {32'hbe765d1e, 32'h3d95ea8a} /* (21, 26, 25) {real, imag} */,
  {32'hbe052d8a, 32'h3f2f788c} /* (21, 26, 24) {real, imag} */,
  {32'h3cc64030, 32'hbee2f9c7} /* (21, 26, 23) {real, imag} */,
  {32'h3bd6bf00, 32'hbf18492c} /* (21, 26, 22) {real, imag} */,
  {32'hbf11e8c2, 32'h3f0066cb} /* (21, 26, 21) {real, imag} */,
  {32'hbe9b616e, 32'hbe05f412} /* (21, 26, 20) {real, imag} */,
  {32'hbd2d5b67, 32'h3ef3bb01} /* (21, 26, 19) {real, imag} */,
  {32'h3e4125ea, 32'hbe18adb0} /* (21, 26, 18) {real, imag} */,
  {32'h3af40f60, 32'hbd796d5e} /* (21, 26, 17) {real, imag} */,
  {32'hbe423fd4, 32'h3e562aad} /* (21, 26, 16) {real, imag} */,
  {32'h3f0630e9, 32'hbe6e77d2} /* (21, 26, 15) {real, imag} */,
  {32'hbe03c696, 32'hbefdb580} /* (21, 26, 14) {real, imag} */,
  {32'hbe8adb2e, 32'h3eaa702b} /* (21, 26, 13) {real, imag} */,
  {32'hbeec2d95, 32'h3c354f10} /* (21, 26, 12) {real, imag} */,
  {32'hbe6038eb, 32'h3d660c80} /* (21, 26, 11) {real, imag} */,
  {32'h3d9c7640, 32'h3eb69056} /* (21, 26, 10) {real, imag} */,
  {32'hbe8dd212, 32'hbef7ff78} /* (21, 26, 9) {real, imag} */,
  {32'hbe8009c6, 32'hbe66a97b} /* (21, 26, 8) {real, imag} */,
  {32'hbe1f4018, 32'h3ea1a559} /* (21, 26, 7) {real, imag} */,
  {32'h3eca7d0e, 32'h3f02638a} /* (21, 26, 6) {real, imag} */,
  {32'hbe7e644c, 32'h3f3aaf9d} /* (21, 26, 5) {real, imag} */,
  {32'h3f2de48c, 32'h3f20a7f5} /* (21, 26, 4) {real, imag} */,
  {32'h3e7e0aa5, 32'hbe04667a} /* (21, 26, 3) {real, imag} */,
  {32'h3d05c200, 32'h3e070388} /* (21, 26, 2) {real, imag} */,
  {32'hbe8be10a, 32'hbf829357} /* (21, 26, 1) {real, imag} */,
  {32'hbe533a47, 32'hbe15f1e1} /* (21, 26, 0) {real, imag} */,
  {32'h3e505b28, 32'h3de05b6f} /* (21, 25, 31) {real, imag} */,
  {32'h3e9c4d14, 32'hbe5ef07c} /* (21, 25, 30) {real, imag} */,
  {32'h3f56105b, 32'hbee26cce} /* (21, 25, 29) {real, imag} */,
  {32'h3c4e6d40, 32'h3eb5830d} /* (21, 25, 28) {real, imag} */,
  {32'h3f55ed6c, 32'h3e85035a} /* (21, 25, 27) {real, imag} */,
  {32'hbe630ddf, 32'hbf15c674} /* (21, 25, 26) {real, imag} */,
  {32'hbf3968ae, 32'h3cf55d90} /* (21, 25, 25) {real, imag} */,
  {32'hbe7139bd, 32'hbc3eeef8} /* (21, 25, 24) {real, imag} */,
  {32'hbe14d9b7, 32'hbdc7f028} /* (21, 25, 23) {real, imag} */,
  {32'hbe4d5d66, 32'h3e510976} /* (21, 25, 22) {real, imag} */,
  {32'hbf2f4b36, 32'hbee2ea48} /* (21, 25, 21) {real, imag} */,
  {32'hbe043ab3, 32'h3e4be7ea} /* (21, 25, 20) {real, imag} */,
  {32'hbd92808e, 32'hbe4ae15b} /* (21, 25, 19) {real, imag} */,
  {32'hbeed2434, 32'hbdc0cdb8} /* (21, 25, 18) {real, imag} */,
  {32'h3c09fca4, 32'hbdb591fe} /* (21, 25, 17) {real, imag} */,
  {32'hbde39f69, 32'h3ed0b56d} /* (21, 25, 16) {real, imag} */,
  {32'hbe9b595c, 32'hbe13efb4} /* (21, 25, 15) {real, imag} */,
  {32'h3d704e38, 32'h3e330e13} /* (21, 25, 14) {real, imag} */,
  {32'h3dbb437c, 32'hbebcbfeb} /* (21, 25, 13) {real, imag} */,
  {32'hbe177cb0, 32'h3c3dbeac} /* (21, 25, 12) {real, imag} */,
  {32'h3cc43f28, 32'h3f1437f4} /* (21, 25, 11) {real, imag} */,
  {32'hbf1df8cb, 32'hbe2a2584} /* (21, 25, 10) {real, imag} */,
  {32'hbe174642, 32'h3e41b15f} /* (21, 25, 9) {real, imag} */,
  {32'hbe1a5dd2, 32'hbf012ca6} /* (21, 25, 8) {real, imag} */,
  {32'hbeae164c, 32'hbee0b147} /* (21, 25, 7) {real, imag} */,
  {32'hbe9b75ba, 32'hbf3209f8} /* (21, 25, 6) {real, imag} */,
  {32'hbeb75d73, 32'hbe201ec5} /* (21, 25, 5) {real, imag} */,
  {32'h3f1e85c6, 32'hbe00a594} /* (21, 25, 4) {real, imag} */,
  {32'h3dd9f536, 32'h3e088e9b} /* (21, 25, 3) {real, imag} */,
  {32'h3f0d938f, 32'h3f47321b} /* (21, 25, 2) {real, imag} */,
  {32'h3c523780, 32'h3ee7c94c} /* (21, 25, 1) {real, imag} */,
  {32'hbf46c9e7, 32'h3f6c1c8e} /* (21, 25, 0) {real, imag} */,
  {32'h3f186e44, 32'hbec9bbf2} /* (21, 24, 31) {real, imag} */,
  {32'hbf1bbb3f, 32'h3e6784d0} /* (21, 24, 30) {real, imag} */,
  {32'h3ef20080, 32'h3e60fefd} /* (21, 24, 29) {real, imag} */,
  {32'h3f0738b9, 32'h3dfbc962} /* (21, 24, 28) {real, imag} */,
  {32'hbf887754, 32'h3deac1d4} /* (21, 24, 27) {real, imag} */,
  {32'h3db5b7cc, 32'hbcabac00} /* (21, 24, 26) {real, imag} */,
  {32'hbd9552f4, 32'h3e4aac96} /* (21, 24, 25) {real, imag} */,
  {32'hbcca14e0, 32'hbd8cafc2} /* (21, 24, 24) {real, imag} */,
  {32'hbd71f840, 32'h3d8c10d8} /* (21, 24, 23) {real, imag} */,
  {32'hbf0db8f6, 32'hbf42438e} /* (21, 24, 22) {real, imag} */,
  {32'hbba99a40, 32'h3f49d051} /* (21, 24, 21) {real, imag} */,
  {32'h3e44c29a, 32'h3eb4c39a} /* (21, 24, 20) {real, imag} */,
  {32'h3c90f380, 32'h3e781da0} /* (21, 24, 19) {real, imag} */,
  {32'hbe6bb5b3, 32'hbd851572} /* (21, 24, 18) {real, imag} */,
  {32'hbe5d22dc, 32'hbe2c4711} /* (21, 24, 17) {real, imag} */,
  {32'h3d07269c, 32'h3e0a9782} /* (21, 24, 16) {real, imag} */,
  {32'h3d84d4cc, 32'hbc977110} /* (21, 24, 15) {real, imag} */,
  {32'hbdd0c5dc, 32'hbeaa805a} /* (21, 24, 14) {real, imag} */,
  {32'h3de2e398, 32'h3ed41651} /* (21, 24, 13) {real, imag} */,
  {32'h3e23eb8b, 32'hbd3fc9b4} /* (21, 24, 12) {real, imag} */,
  {32'hbdf09a8e, 32'hbf495788} /* (21, 24, 11) {real, imag} */,
  {32'hbb878d80, 32'h3dbab0d8} /* (21, 24, 10) {real, imag} */,
  {32'h3e9c3a13, 32'hbe9e78b7} /* (21, 24, 9) {real, imag} */,
  {32'hbe198693, 32'h3f028a0c} /* (21, 24, 8) {real, imag} */,
  {32'h3e7742b3, 32'h3df803d0} /* (21, 24, 7) {real, imag} */,
  {32'h3f73339a, 32'h3be41a00} /* (21, 24, 6) {real, imag} */,
  {32'hbf54a9fe, 32'h3f11bb49} /* (21, 24, 5) {real, imag} */,
  {32'h3df5ec40, 32'hbe93132b} /* (21, 24, 4) {real, imag} */,
  {32'h3e8451b2, 32'hbcfc6b18} /* (21, 24, 3) {real, imag} */,
  {32'hbf3b04cd, 32'h3ed1d501} /* (21, 24, 2) {real, imag} */,
  {32'h3f956bc1, 32'hbf852325} /* (21, 24, 1) {real, imag} */,
  {32'h3e9e3e58, 32'h3e424b1c} /* (21, 24, 0) {real, imag} */,
  {32'hbf2c64f8, 32'h3dbde9dc} /* (21, 23, 31) {real, imag} */,
  {32'hbd082fbc, 32'hbeb2c967} /* (21, 23, 30) {real, imag} */,
  {32'h3ed28adf, 32'h3eb1aa87} /* (21, 23, 29) {real, imag} */,
  {32'hbef36f04, 32'hbd9dd7ef} /* (21, 23, 28) {real, imag} */,
  {32'h3f3dea61, 32'hbe289747} /* (21, 23, 27) {real, imag} */,
  {32'hbec96e07, 32'h3f516a40} /* (21, 23, 26) {real, imag} */,
  {32'h3e415b7c, 32'h3f223ddc} /* (21, 23, 25) {real, imag} */,
  {32'hbefb1608, 32'hbe4ae552} /* (21, 23, 24) {real, imag} */,
  {32'h3f34f97a, 32'h3e551398} /* (21, 23, 23) {real, imag} */,
  {32'h3e9e3e20, 32'h3e5701c7} /* (21, 23, 22) {real, imag} */,
  {32'h3c211430, 32'hbee3c516} /* (21, 23, 21) {real, imag} */,
  {32'hbf25acbf, 32'hbdd41d60} /* (21, 23, 20) {real, imag} */,
  {32'hbe2c8392, 32'hbe60bb37} /* (21, 23, 19) {real, imag} */,
  {32'h3c1be448, 32'hbebab478} /* (21, 23, 18) {real, imag} */,
  {32'h3e07eb8a, 32'h3dc02015} /* (21, 23, 17) {real, imag} */,
  {32'hbb75cd40, 32'hbe11f94f} /* (21, 23, 16) {real, imag} */,
  {32'hbe0b4b3c, 32'h3f1cc79e} /* (21, 23, 15) {real, imag} */,
  {32'h3ea5d6c7, 32'hbde8cd36} /* (21, 23, 14) {real, imag} */,
  {32'hbd8c7c80, 32'h3da45668} /* (21, 23, 13) {real, imag} */,
  {32'h3d8e5c44, 32'hbe1bce5e} /* (21, 23, 12) {real, imag} */,
  {32'hbe8307d3, 32'hbdba3544} /* (21, 23, 11) {real, imag} */,
  {32'hbe33ce7f, 32'h3f07346a} /* (21, 23, 10) {real, imag} */,
  {32'hbc9f4ce4, 32'h3b8e1080} /* (21, 23, 9) {real, imag} */,
  {32'hbe0f7c11, 32'hbf052dbd} /* (21, 23, 8) {real, imag} */,
  {32'hbe4ae2a4, 32'hbe1009c5} /* (21, 23, 7) {real, imag} */,
  {32'hbdf84c4c, 32'hbd377e14} /* (21, 23, 6) {real, imag} */,
  {32'h3dce0378, 32'h3e56bc65} /* (21, 23, 5) {real, imag} */,
  {32'hbd5625e8, 32'h3f1cf116} /* (21, 23, 4) {real, imag} */,
  {32'hbea6acbc, 32'h3ef48036} /* (21, 23, 3) {real, imag} */,
  {32'hbdf6b3be, 32'hbe9d2e84} /* (21, 23, 2) {real, imag} */,
  {32'h3ef1b561, 32'hbefe8fca} /* (21, 23, 1) {real, imag} */,
  {32'h3f06b3e3, 32'hbea28e66} /* (21, 23, 0) {real, imag} */,
  {32'hbf70e694, 32'h3ee93db2} /* (21, 22, 31) {real, imag} */,
  {32'h3e591e1a, 32'h3d369548} /* (21, 22, 30) {real, imag} */,
  {32'h3d7b40cc, 32'h3c96cf28} /* (21, 22, 29) {real, imag} */,
  {32'h3dd41328, 32'hbec5d2b8} /* (21, 22, 28) {real, imag} */,
  {32'hbef3fd64, 32'h3ee80ed3} /* (21, 22, 27) {real, imag} */,
  {32'h3edc72fa, 32'h3f036d7c} /* (21, 22, 26) {real, imag} */,
  {32'hbe7fe706, 32'hbdee3219} /* (21, 22, 25) {real, imag} */,
  {32'hbe742492, 32'h3e8457b8} /* (21, 22, 24) {real, imag} */,
  {32'hbd33ded0, 32'h3d3ab364} /* (21, 22, 23) {real, imag} */,
  {32'h3ed2a866, 32'hbeefb632} /* (21, 22, 22) {real, imag} */,
  {32'hbde1d9e0, 32'hbd8c6cec} /* (21, 22, 21) {real, imag} */,
  {32'hbdb8167c, 32'hbf0d67e8} /* (21, 22, 20) {real, imag} */,
  {32'hbde85b45, 32'h3d428370} /* (21, 22, 19) {real, imag} */,
  {32'hbd6102ce, 32'h3e469c80} /* (21, 22, 18) {real, imag} */,
  {32'h3e48acb2, 32'h3c4bd1d0} /* (21, 22, 17) {real, imag} */,
  {32'h3f090f35, 32'h3e53e9ba} /* (21, 22, 16) {real, imag} */,
  {32'hbe91b11a, 32'hbecb3cc0} /* (21, 22, 15) {real, imag} */,
  {32'h3a781c40, 32'h3e71a102} /* (21, 22, 14) {real, imag} */,
  {32'hbe5cbcd7, 32'h3e04ae55} /* (21, 22, 13) {real, imag} */,
  {32'hbc94d074, 32'h3eefb11a} /* (21, 22, 12) {real, imag} */,
  {32'h3f224b53, 32'h3e7abfb4} /* (21, 22, 11) {real, imag} */,
  {32'h3bdd9fb0, 32'h3e8d12f5} /* (21, 22, 10) {real, imag} */,
  {32'hbed39aa6, 32'h3e463d94} /* (21, 22, 9) {real, imag} */,
  {32'h3eafb52a, 32'hbe26163e} /* (21, 22, 8) {real, imag} */,
  {32'hbf0b2b00, 32'h3dead684} /* (21, 22, 7) {real, imag} */,
  {32'h3ea03376, 32'hbebe7db1} /* (21, 22, 6) {real, imag} */,
  {32'h3e906aeb, 32'hbe24f73b} /* (21, 22, 5) {real, imag} */,
  {32'hbea29643, 32'hbdddb6ef} /* (21, 22, 4) {real, imag} */,
  {32'h3dbc7839, 32'h3d2de910} /* (21, 22, 3) {real, imag} */,
  {32'h3ed1c0ef, 32'hbf289d7b} /* (21, 22, 2) {real, imag} */,
  {32'h3ebd8b1c, 32'h3f760b3e} /* (21, 22, 1) {real, imag} */,
  {32'hbf5ad4c8, 32'h3e4ac227} /* (21, 22, 0) {real, imag} */,
  {32'h3d7a5853, 32'hbf19bf30} /* (21, 21, 31) {real, imag} */,
  {32'h3e78aa08, 32'h3ea54854} /* (21, 21, 30) {real, imag} */,
  {32'h3eb31ef5, 32'h3f038600} /* (21, 21, 29) {real, imag} */,
  {32'hbe95f8b0, 32'hbe0c445e} /* (21, 21, 28) {real, imag} */,
  {32'h3ed35014, 32'h3d54a4b0} /* (21, 21, 27) {real, imag} */,
  {32'h3ec5a0c2, 32'hbe6652a7} /* (21, 21, 26) {real, imag} */,
  {32'h3e91a605, 32'h3d4bac38} /* (21, 21, 25) {real, imag} */,
  {32'h3eedbfbf, 32'h3b5c8180} /* (21, 21, 24) {real, imag} */,
  {32'h3ecbaa62, 32'h3e9a7108} /* (21, 21, 23) {real, imag} */,
  {32'h3e0a3b45, 32'h3d5722d8} /* (21, 21, 22) {real, imag} */,
  {32'hbf064264, 32'h3ca99afc} /* (21, 21, 21) {real, imag} */,
  {32'hbec4da70, 32'hbeabc2bd} /* (21, 21, 20) {real, imag} */,
  {32'hbd997313, 32'hbde049f6} /* (21, 21, 19) {real, imag} */,
  {32'h3b789b40, 32'hbe16a9c6} /* (21, 21, 18) {real, imag} */,
  {32'h3d883876, 32'h3e84a76e} /* (21, 21, 17) {real, imag} */,
  {32'hbedcaec6, 32'hbe9c11e5} /* (21, 21, 16) {real, imag} */,
  {32'hbe03a6ec, 32'h3e2f1030} /* (21, 21, 15) {real, imag} */,
  {32'h3ee84bbe, 32'h3f113ff1} /* (21, 21, 14) {real, imag} */,
  {32'h3eb4ea39, 32'hbe6f7f97} /* (21, 21, 13) {real, imag} */,
  {32'h3e321faa, 32'hbc4e1ec0} /* (21, 21, 12) {real, imag} */,
  {32'hbe7ccd98, 32'hbe9b2a41} /* (21, 21, 11) {real, imag} */,
  {32'h3ed79ee8, 32'h3e78d3b0} /* (21, 21, 10) {real, imag} */,
  {32'h3d079a6c, 32'h3d424928} /* (21, 21, 9) {real, imag} */,
  {32'h3ea5f604, 32'h3de6f3b2} /* (21, 21, 8) {real, imag} */,
  {32'hbe7a8bf8, 32'hbde00e0c} /* (21, 21, 7) {real, imag} */,
  {32'hbef904e3, 32'h3e4d8ff0} /* (21, 21, 6) {real, imag} */,
  {32'hbda072f2, 32'hbeb0e5fe} /* (21, 21, 5) {real, imag} */,
  {32'hbf273d46, 32'hbe0f4f5f} /* (21, 21, 4) {real, imag} */,
  {32'h3d91d856, 32'hbe00797b} /* (21, 21, 3) {real, imag} */,
  {32'hbf4ade5b, 32'hbd9c217d} /* (21, 21, 2) {real, imag} */,
  {32'h3ea01852, 32'hbde9af7e} /* (21, 21, 1) {real, imag} */,
  {32'h3ebecdfb, 32'hbf2917ed} /* (21, 21, 0) {real, imag} */,
  {32'h3dd0d53d, 32'h3e228556} /* (21, 20, 31) {real, imag} */,
  {32'h3dd416f6, 32'h3e4470b4} /* (21, 20, 30) {real, imag} */,
  {32'hbe55dadd, 32'hbe22dad7} /* (21, 20, 29) {real, imag} */,
  {32'h3e888516, 32'h3dc4c705} /* (21, 20, 28) {real, imag} */,
  {32'h3e83ad56, 32'h3d9a7554} /* (21, 20, 27) {real, imag} */,
  {32'h3e8e0ffa, 32'hbdbb274c} /* (21, 20, 26) {real, imag} */,
  {32'hbf2023c8, 32'hbdb72dbc} /* (21, 20, 25) {real, imag} */,
  {32'hbec3acc6, 32'hbeb351a6} /* (21, 20, 24) {real, imag} */,
  {32'h3e5a209b, 32'h3e6fd856} /* (21, 20, 23) {real, imag} */,
  {32'hbdafe40e, 32'hbe6b3ab6} /* (21, 20, 22) {real, imag} */,
  {32'hbf0bdb46, 32'hbd9bb139} /* (21, 20, 21) {real, imag} */,
  {32'h3ef54a2c, 32'hbef0b9b0} /* (21, 20, 20) {real, imag} */,
  {32'h3e5bc5a7, 32'hbdbb9e45} /* (21, 20, 19) {real, imag} */,
  {32'h3e39a501, 32'hbd1eb0f8} /* (21, 20, 18) {real, imag} */,
  {32'h3e5a2d46, 32'h3ebb5ea0} /* (21, 20, 17) {real, imag} */,
  {32'hbe51ea52, 32'hbe4f51a4} /* (21, 20, 16) {real, imag} */,
  {32'h3ee22385, 32'hbeae5653} /* (21, 20, 15) {real, imag} */,
  {32'h3e81ce7e, 32'h3ee28062} /* (21, 20, 14) {real, imag} */,
  {32'h3d9a5cd7, 32'h3d8409fe} /* (21, 20, 13) {real, imag} */,
  {32'h3e554c5c, 32'h3f12df42} /* (21, 20, 12) {real, imag} */,
  {32'h3f6fbce0, 32'hbe22bd34} /* (21, 20, 11) {real, imag} */,
  {32'h3dcd7a84, 32'hbc4c0a0c} /* (21, 20, 10) {real, imag} */,
  {32'h3ef6d3e8, 32'h3db7c210} /* (21, 20, 9) {real, imag} */,
  {32'h3da81c7c, 32'hbeadca3f} /* (21, 20, 8) {real, imag} */,
  {32'h3e9e026b, 32'h3bccf3e0} /* (21, 20, 7) {real, imag} */,
  {32'hbf38cb9c, 32'hbe3c2390} /* (21, 20, 6) {real, imag} */,
  {32'h3d019ee2, 32'h3ec1e1db} /* (21, 20, 5) {real, imag} */,
  {32'hbe273185, 32'hbe50b578} /* (21, 20, 4) {real, imag} */,
  {32'h3cbf81d4, 32'h3eaa7a2a} /* (21, 20, 3) {real, imag} */,
  {32'hbeeef9f8, 32'h3df8f5c0} /* (21, 20, 2) {real, imag} */,
  {32'hbe0aa9d4, 32'hbcf815f8} /* (21, 20, 1) {real, imag} */,
  {32'h3f49bc09, 32'hbea9d1c4} /* (21, 20, 0) {real, imag} */,
  {32'hbf392bb0, 32'h3e964d96} /* (21, 19, 31) {real, imag} */,
  {32'hbece4ac1, 32'h3bcef6c0} /* (21, 19, 30) {real, imag} */,
  {32'hbe932e18, 32'h3d5078b6} /* (21, 19, 29) {real, imag} */,
  {32'h3ebde89d, 32'h3e8b7ac3} /* (21, 19, 28) {real, imag} */,
  {32'h3ea3eeb4, 32'h3f10c37e} /* (21, 19, 27) {real, imag} */,
  {32'hbeb2b89e, 32'hbf3fb61a} /* (21, 19, 26) {real, imag} */,
  {32'hb9fe5c00, 32'h3e3f9283} /* (21, 19, 25) {real, imag} */,
  {32'h3f0fc9c8, 32'hbec4021e} /* (21, 19, 24) {real, imag} */,
  {32'hbdcf3b62, 32'h3dc1f490} /* (21, 19, 23) {real, imag} */,
  {32'hbed8e6e0, 32'hbe554c50} /* (21, 19, 22) {real, imag} */,
  {32'h3ea1ccf5, 32'h3f26c184} /* (21, 19, 21) {real, imag} */,
  {32'hbe8cef3e, 32'hbec56134} /* (21, 19, 20) {real, imag} */,
  {32'h3eb0e958, 32'h3d5fa6d0} /* (21, 19, 19) {real, imag} */,
  {32'h3f1cff7f, 32'hbe42c5f0} /* (21, 19, 18) {real, imag} */,
  {32'h3caa46b6, 32'h3d5bb3c0} /* (21, 19, 17) {real, imag} */,
  {32'hbeb792a9, 32'h3db834fc} /* (21, 19, 16) {real, imag} */,
  {32'hbe224e52, 32'h3e5cc876} /* (21, 19, 15) {real, imag} */,
  {32'h3e8453f5, 32'hbe87564b} /* (21, 19, 14) {real, imag} */,
  {32'hbeab57ff, 32'hbe65f7ca} /* (21, 19, 13) {real, imag} */,
  {32'h3df77974, 32'hbdb11f74} /* (21, 19, 12) {real, imag} */,
  {32'h3d6d0438, 32'hbe29e829} /* (21, 19, 11) {real, imag} */,
  {32'h3eb43332, 32'hbca834a8} /* (21, 19, 10) {real, imag} */,
  {32'h3e462d96, 32'h3e24c1a2} /* (21, 19, 9) {real, imag} */,
  {32'h3e600d04, 32'h3efde83a} /* (21, 19, 8) {real, imag} */,
  {32'hbe272ef9, 32'hbefcd96e} /* (21, 19, 7) {real, imag} */,
  {32'hbf299d4e, 32'h3e1f4bd1} /* (21, 19, 6) {real, imag} */,
  {32'hbdd68c1b, 32'h3e0c65f3} /* (21, 19, 5) {real, imag} */,
  {32'hbe125ba1, 32'h3e447b43} /* (21, 19, 4) {real, imag} */,
  {32'h3ea05238, 32'hbf0398e4} /* (21, 19, 3) {real, imag} */,
  {32'hbf1653eb, 32'h3dcccd78} /* (21, 19, 2) {real, imag} */,
  {32'h3e8e1954, 32'hbdd7b80c} /* (21, 19, 1) {real, imag} */,
  {32'hbe85b42f, 32'h3d7ff12c} /* (21, 19, 0) {real, imag} */,
  {32'hbe63447a, 32'hbb98d2c0} /* (21, 18, 31) {real, imag} */,
  {32'hbe38d353, 32'hbd8094ff} /* (21, 18, 30) {real, imag} */,
  {32'h3de0e670, 32'h3d359948} /* (21, 18, 29) {real, imag} */,
  {32'h3db81b2c, 32'hbdad413c} /* (21, 18, 28) {real, imag} */,
  {32'hbe6a76c5, 32'h3e57e048} /* (21, 18, 27) {real, imag} */,
  {32'hbe7b3f8d, 32'h3c41cd4c} /* (21, 18, 26) {real, imag} */,
  {32'hbeec80f0, 32'hbe56b64c} /* (21, 18, 25) {real, imag} */,
  {32'h3ebdd722, 32'h3bb0f320} /* (21, 18, 24) {real, imag} */,
  {32'hbe8debd2, 32'hbf0ec8ed} /* (21, 18, 23) {real, imag} */,
  {32'h3dced554, 32'hbed1d598} /* (21, 18, 22) {real, imag} */,
  {32'h3e9e0c5a, 32'hbddc9eb8} /* (21, 18, 21) {real, imag} */,
  {32'h3f30c67d, 32'h3ed087e4} /* (21, 18, 20) {real, imag} */,
  {32'h3dbf3104, 32'hbe541ce2} /* (21, 18, 19) {real, imag} */,
  {32'hbdc91cd0, 32'h3e66abbb} /* (21, 18, 18) {real, imag} */,
  {32'h3df1874a, 32'h3ef703d2} /* (21, 18, 17) {real, imag} */,
  {32'hbd0dd91c, 32'h3e1b7f06} /* (21, 18, 16) {real, imag} */,
  {32'hbf03cd7d, 32'h3d1548a8} /* (21, 18, 15) {real, imag} */,
  {32'h3e86f027, 32'hbdd75cda} /* (21, 18, 14) {real, imag} */,
  {32'hbdb1b4a2, 32'hbecfdd0b} /* (21, 18, 13) {real, imag} */,
  {32'hbeae6808, 32'h3dfdc60b} /* (21, 18, 12) {real, imag} */,
  {32'hbedb3e08, 32'hbe5d6808} /* (21, 18, 11) {real, imag} */,
  {32'hbee7251c, 32'hbd90e9d8} /* (21, 18, 10) {real, imag} */,
  {32'hbd97d881, 32'h3e496d20} /* (21, 18, 9) {real, imag} */,
  {32'hbedf24ac, 32'h3e7cdbc3} /* (21, 18, 8) {real, imag} */,
  {32'h3c246134, 32'hbee0f968} /* (21, 18, 7) {real, imag} */,
  {32'hbcfb7c78, 32'hbed517f9} /* (21, 18, 6) {real, imag} */,
  {32'hbdb6d4b6, 32'h3d914870} /* (21, 18, 5) {real, imag} */,
  {32'h3ec26593, 32'h3cf1c950} /* (21, 18, 4) {real, imag} */,
  {32'h3e9e0726, 32'h3e11b13e} /* (21, 18, 3) {real, imag} */,
  {32'hbe8add00, 32'h3d949a74} /* (21, 18, 2) {real, imag} */,
  {32'h3e72a63a, 32'hbf079689} /* (21, 18, 1) {real, imag} */,
  {32'hbe6848e2, 32'hbef97276} /* (21, 18, 0) {real, imag} */,
  {32'h3e266ace, 32'hbe6e319a} /* (21, 17, 31) {real, imag} */,
  {32'h3e829f17, 32'hbe8edd29} /* (21, 17, 30) {real, imag} */,
  {32'h3ceeedf8, 32'h3e1cd37a} /* (21, 17, 29) {real, imag} */,
  {32'hbed2df54, 32'hbe2a5e72} /* (21, 17, 28) {real, imag} */,
  {32'hbebef61c, 32'h3e452c81} /* (21, 17, 27) {real, imag} */,
  {32'hbc90627c, 32'h3d412628} /* (21, 17, 26) {real, imag} */,
  {32'hbd12ed96, 32'h3d054af0} /* (21, 17, 25) {real, imag} */,
  {32'hbe89b7d9, 32'h3df3c8f9} /* (21, 17, 24) {real, imag} */,
  {32'hbe30f7ce, 32'hbe1caaa6} /* (21, 17, 23) {real, imag} */,
  {32'h3f00b474, 32'h3e18440f} /* (21, 17, 22) {real, imag} */,
  {32'h3e1745dd, 32'hbefdb58e} /* (21, 17, 21) {real, imag} */,
  {32'h3e831d19, 32'h3e0bd5c3} /* (21, 17, 20) {real, imag} */,
  {32'hbd8a344a, 32'h3e3b83fa} /* (21, 17, 19) {real, imag} */,
  {32'hbdefac64, 32'h3e665399} /* (21, 17, 18) {real, imag} */,
  {32'h3d980bc4, 32'hbecb03f1} /* (21, 17, 17) {real, imag} */,
  {32'hbe8fdc35, 32'h3e9bf7d1} /* (21, 17, 16) {real, imag} */,
  {32'h3e79a65b, 32'hbee8c672} /* (21, 17, 15) {real, imag} */,
  {32'h3d6bcdf8, 32'hbdff792c} /* (21, 17, 14) {real, imag} */,
  {32'hbd2ca420, 32'h3e3d52ca} /* (21, 17, 13) {real, imag} */,
  {32'h3d967124, 32'h3da34208} /* (21, 17, 12) {real, imag} */,
  {32'hbf0968f4, 32'hbec85712} /* (21, 17, 11) {real, imag} */,
  {32'hbed3e3bc, 32'h3e6794e5} /* (21, 17, 10) {real, imag} */,
  {32'h3e8e07b5, 32'h3c3f8bb0} /* (21, 17, 9) {real, imag} */,
  {32'hbe9c109c, 32'h3e025cec} /* (21, 17, 8) {real, imag} */,
  {32'hbd1c5f84, 32'h3e2e5b57} /* (21, 17, 7) {real, imag} */,
  {32'hbe28ffbd, 32'hbdc037ad} /* (21, 17, 6) {real, imag} */,
  {32'hbdf89d30, 32'h3e323947} /* (21, 17, 5) {real, imag} */,
  {32'h3df96fe4, 32'hbafc8a40} /* (21, 17, 4) {real, imag} */,
  {32'h3e14546c, 32'hbde21393} /* (21, 17, 3) {real, imag} */,
  {32'hbddd4069, 32'h3dd2980f} /* (21, 17, 2) {real, imag} */,
  {32'h3e94ec56, 32'h3dbf8abc} /* (21, 17, 1) {real, imag} */,
  {32'h3e5e4622, 32'h3e68eed8} /* (21, 17, 0) {real, imag} */,
  {32'h3ddcb700, 32'h3d253ea5} /* (21, 16, 31) {real, imag} */,
  {32'h3dc26d33, 32'hbe4fed72} /* (21, 16, 30) {real, imag} */,
  {32'hbd3037fd, 32'hbe3099b7} /* (21, 16, 29) {real, imag} */,
  {32'hbed4b3ee, 32'hbe083c57} /* (21, 16, 28) {real, imag} */,
  {32'hbcc9ad3c, 32'hbeaf6c18} /* (21, 16, 27) {real, imag} */,
  {32'hbe66b13d, 32'hbd8f2c91} /* (21, 16, 26) {real, imag} */,
  {32'hbca6ee7a, 32'hbe004ccc} /* (21, 16, 25) {real, imag} */,
  {32'h3dac2e4c, 32'h3b8f2390} /* (21, 16, 24) {real, imag} */,
  {32'hbc903a08, 32'h3e47bc36} /* (21, 16, 23) {real, imag} */,
  {32'h3e7bdecb, 32'hbc6a0fae} /* (21, 16, 22) {real, imag} */,
  {32'hbd8cfb3c, 32'hbde4e78c} /* (21, 16, 21) {real, imag} */,
  {32'h3dffbb09, 32'hbe842226} /* (21, 16, 20) {real, imag} */,
  {32'hbe5da24e, 32'hbe7caad3} /* (21, 16, 19) {real, imag} */,
  {32'h3db4d51c, 32'hbdc5ca76} /* (21, 16, 18) {real, imag} */,
  {32'h3d1d5bb5, 32'hbceeead0} /* (21, 16, 17) {real, imag} */,
  {32'hbdd87578, 32'h00000000} /* (21, 16, 16) {real, imag} */,
  {32'h3d1d5bb5, 32'h3ceeead0} /* (21, 16, 15) {real, imag} */,
  {32'h3db4d51c, 32'h3dc5ca76} /* (21, 16, 14) {real, imag} */,
  {32'hbe5da24e, 32'h3e7caad3} /* (21, 16, 13) {real, imag} */,
  {32'h3dffbb09, 32'h3e842226} /* (21, 16, 12) {real, imag} */,
  {32'hbd8cfb3c, 32'h3de4e78c} /* (21, 16, 11) {real, imag} */,
  {32'h3e7bdecb, 32'h3c6a0fae} /* (21, 16, 10) {real, imag} */,
  {32'hbc903a08, 32'hbe47bc36} /* (21, 16, 9) {real, imag} */,
  {32'h3dac2e4c, 32'hbb8f2390} /* (21, 16, 8) {real, imag} */,
  {32'hbca6ee7a, 32'h3e004ccc} /* (21, 16, 7) {real, imag} */,
  {32'hbe66b13d, 32'h3d8f2c91} /* (21, 16, 6) {real, imag} */,
  {32'hbcc9ad3c, 32'h3eaf6c18} /* (21, 16, 5) {real, imag} */,
  {32'hbed4b3ee, 32'h3e083c57} /* (21, 16, 4) {real, imag} */,
  {32'hbd3037fd, 32'h3e3099b7} /* (21, 16, 3) {real, imag} */,
  {32'h3dc26d33, 32'h3e4fed72} /* (21, 16, 2) {real, imag} */,
  {32'h3ddcb700, 32'hbd253ea5} /* (21, 16, 1) {real, imag} */,
  {32'h3e8d583c, 32'h00000000} /* (21, 16, 0) {real, imag} */,
  {32'h3e94ec56, 32'hbdbf8abc} /* (21, 15, 31) {real, imag} */,
  {32'hbddd4069, 32'hbdd2980f} /* (21, 15, 30) {real, imag} */,
  {32'h3e14546c, 32'h3de21393} /* (21, 15, 29) {real, imag} */,
  {32'h3df96fe4, 32'h3afc8a40} /* (21, 15, 28) {real, imag} */,
  {32'hbdf89d30, 32'hbe323947} /* (21, 15, 27) {real, imag} */,
  {32'hbe28ffbd, 32'h3dc037ad} /* (21, 15, 26) {real, imag} */,
  {32'hbd1c5f84, 32'hbe2e5b57} /* (21, 15, 25) {real, imag} */,
  {32'hbe9c109c, 32'hbe025cec} /* (21, 15, 24) {real, imag} */,
  {32'h3e8e07b5, 32'hbc3f8bb0} /* (21, 15, 23) {real, imag} */,
  {32'hbed3e3bc, 32'hbe6794e5} /* (21, 15, 22) {real, imag} */,
  {32'hbf0968f4, 32'h3ec85712} /* (21, 15, 21) {real, imag} */,
  {32'h3d967124, 32'hbda34208} /* (21, 15, 20) {real, imag} */,
  {32'hbd2ca420, 32'hbe3d52ca} /* (21, 15, 19) {real, imag} */,
  {32'h3d6bcdf8, 32'h3dff792c} /* (21, 15, 18) {real, imag} */,
  {32'h3e79a65b, 32'h3ee8c672} /* (21, 15, 17) {real, imag} */,
  {32'hbe8fdc35, 32'hbe9bf7d1} /* (21, 15, 16) {real, imag} */,
  {32'h3d980bc4, 32'h3ecb03f1} /* (21, 15, 15) {real, imag} */,
  {32'hbdefac64, 32'hbe665399} /* (21, 15, 14) {real, imag} */,
  {32'hbd8a344a, 32'hbe3b83fa} /* (21, 15, 13) {real, imag} */,
  {32'h3e831d19, 32'hbe0bd5c3} /* (21, 15, 12) {real, imag} */,
  {32'h3e1745dd, 32'h3efdb58e} /* (21, 15, 11) {real, imag} */,
  {32'h3f00b474, 32'hbe18440f} /* (21, 15, 10) {real, imag} */,
  {32'hbe30f7ce, 32'h3e1caaa6} /* (21, 15, 9) {real, imag} */,
  {32'hbe89b7d9, 32'hbdf3c8f9} /* (21, 15, 8) {real, imag} */,
  {32'hbd12ed96, 32'hbd054af0} /* (21, 15, 7) {real, imag} */,
  {32'hbc90627c, 32'hbd412628} /* (21, 15, 6) {real, imag} */,
  {32'hbebef61c, 32'hbe452c81} /* (21, 15, 5) {real, imag} */,
  {32'hbed2df54, 32'h3e2a5e72} /* (21, 15, 4) {real, imag} */,
  {32'h3ceeedf8, 32'hbe1cd37a} /* (21, 15, 3) {real, imag} */,
  {32'h3e829f17, 32'h3e8edd29} /* (21, 15, 2) {real, imag} */,
  {32'h3e266ace, 32'h3e6e319a} /* (21, 15, 1) {real, imag} */,
  {32'h3e5e4622, 32'hbe68eed8} /* (21, 15, 0) {real, imag} */,
  {32'h3e72a63a, 32'h3f079689} /* (21, 14, 31) {real, imag} */,
  {32'hbe8add00, 32'hbd949a74} /* (21, 14, 30) {real, imag} */,
  {32'h3e9e0726, 32'hbe11b13e} /* (21, 14, 29) {real, imag} */,
  {32'h3ec26593, 32'hbcf1c950} /* (21, 14, 28) {real, imag} */,
  {32'hbdb6d4b6, 32'hbd914870} /* (21, 14, 27) {real, imag} */,
  {32'hbcfb7c78, 32'h3ed517f9} /* (21, 14, 26) {real, imag} */,
  {32'h3c246134, 32'h3ee0f968} /* (21, 14, 25) {real, imag} */,
  {32'hbedf24ac, 32'hbe7cdbc3} /* (21, 14, 24) {real, imag} */,
  {32'hbd97d881, 32'hbe496d20} /* (21, 14, 23) {real, imag} */,
  {32'hbee7251c, 32'h3d90e9d8} /* (21, 14, 22) {real, imag} */,
  {32'hbedb3e08, 32'h3e5d6808} /* (21, 14, 21) {real, imag} */,
  {32'hbeae6808, 32'hbdfdc60b} /* (21, 14, 20) {real, imag} */,
  {32'hbdb1b4a2, 32'h3ecfdd0b} /* (21, 14, 19) {real, imag} */,
  {32'h3e86f027, 32'h3dd75cda} /* (21, 14, 18) {real, imag} */,
  {32'hbf03cd7d, 32'hbd1548a8} /* (21, 14, 17) {real, imag} */,
  {32'hbd0dd91c, 32'hbe1b7f06} /* (21, 14, 16) {real, imag} */,
  {32'h3df1874a, 32'hbef703d2} /* (21, 14, 15) {real, imag} */,
  {32'hbdc91cd0, 32'hbe66abbb} /* (21, 14, 14) {real, imag} */,
  {32'h3dbf3104, 32'h3e541ce2} /* (21, 14, 13) {real, imag} */,
  {32'h3f30c67d, 32'hbed087e4} /* (21, 14, 12) {real, imag} */,
  {32'h3e9e0c5a, 32'h3ddc9eb8} /* (21, 14, 11) {real, imag} */,
  {32'h3dced554, 32'h3ed1d598} /* (21, 14, 10) {real, imag} */,
  {32'hbe8debd2, 32'h3f0ec8ed} /* (21, 14, 9) {real, imag} */,
  {32'h3ebdd722, 32'hbbb0f320} /* (21, 14, 8) {real, imag} */,
  {32'hbeec80f0, 32'h3e56b64c} /* (21, 14, 7) {real, imag} */,
  {32'hbe7b3f8d, 32'hbc41cd4c} /* (21, 14, 6) {real, imag} */,
  {32'hbe6a76c5, 32'hbe57e048} /* (21, 14, 5) {real, imag} */,
  {32'h3db81b2c, 32'h3dad413c} /* (21, 14, 4) {real, imag} */,
  {32'h3de0e670, 32'hbd359948} /* (21, 14, 3) {real, imag} */,
  {32'hbe38d353, 32'h3d8094ff} /* (21, 14, 2) {real, imag} */,
  {32'hbe63447a, 32'h3b98d2c0} /* (21, 14, 1) {real, imag} */,
  {32'hbe6848e2, 32'h3ef97276} /* (21, 14, 0) {real, imag} */,
  {32'h3e8e1954, 32'h3dd7b80c} /* (21, 13, 31) {real, imag} */,
  {32'hbf1653eb, 32'hbdcccd78} /* (21, 13, 30) {real, imag} */,
  {32'h3ea05238, 32'h3f0398e4} /* (21, 13, 29) {real, imag} */,
  {32'hbe125ba1, 32'hbe447b43} /* (21, 13, 28) {real, imag} */,
  {32'hbdd68c1b, 32'hbe0c65f3} /* (21, 13, 27) {real, imag} */,
  {32'hbf299d4e, 32'hbe1f4bd1} /* (21, 13, 26) {real, imag} */,
  {32'hbe272ef9, 32'h3efcd96e} /* (21, 13, 25) {real, imag} */,
  {32'h3e600d04, 32'hbefde83a} /* (21, 13, 24) {real, imag} */,
  {32'h3e462d96, 32'hbe24c1a2} /* (21, 13, 23) {real, imag} */,
  {32'h3eb43332, 32'h3ca834a8} /* (21, 13, 22) {real, imag} */,
  {32'h3d6d0438, 32'h3e29e829} /* (21, 13, 21) {real, imag} */,
  {32'h3df77974, 32'h3db11f74} /* (21, 13, 20) {real, imag} */,
  {32'hbeab57ff, 32'h3e65f7ca} /* (21, 13, 19) {real, imag} */,
  {32'h3e8453f5, 32'h3e87564b} /* (21, 13, 18) {real, imag} */,
  {32'hbe224e52, 32'hbe5cc876} /* (21, 13, 17) {real, imag} */,
  {32'hbeb792a9, 32'hbdb834fc} /* (21, 13, 16) {real, imag} */,
  {32'h3caa46b6, 32'hbd5bb3c0} /* (21, 13, 15) {real, imag} */,
  {32'h3f1cff7f, 32'h3e42c5f0} /* (21, 13, 14) {real, imag} */,
  {32'h3eb0e958, 32'hbd5fa6d0} /* (21, 13, 13) {real, imag} */,
  {32'hbe8cef3e, 32'h3ec56134} /* (21, 13, 12) {real, imag} */,
  {32'h3ea1ccf5, 32'hbf26c184} /* (21, 13, 11) {real, imag} */,
  {32'hbed8e6e0, 32'h3e554c50} /* (21, 13, 10) {real, imag} */,
  {32'hbdcf3b62, 32'hbdc1f490} /* (21, 13, 9) {real, imag} */,
  {32'h3f0fc9c8, 32'h3ec4021e} /* (21, 13, 8) {real, imag} */,
  {32'hb9fe5c00, 32'hbe3f9283} /* (21, 13, 7) {real, imag} */,
  {32'hbeb2b89e, 32'h3f3fb61a} /* (21, 13, 6) {real, imag} */,
  {32'h3ea3eeb4, 32'hbf10c37e} /* (21, 13, 5) {real, imag} */,
  {32'h3ebde89d, 32'hbe8b7ac3} /* (21, 13, 4) {real, imag} */,
  {32'hbe932e18, 32'hbd5078b6} /* (21, 13, 3) {real, imag} */,
  {32'hbece4ac1, 32'hbbcef6c0} /* (21, 13, 2) {real, imag} */,
  {32'hbf392bb0, 32'hbe964d96} /* (21, 13, 1) {real, imag} */,
  {32'hbe85b42f, 32'hbd7ff12c} /* (21, 13, 0) {real, imag} */,
  {32'hbe0aa9d4, 32'h3cf815f8} /* (21, 12, 31) {real, imag} */,
  {32'hbeeef9f8, 32'hbdf8f5c0} /* (21, 12, 30) {real, imag} */,
  {32'h3cbf81d4, 32'hbeaa7a2a} /* (21, 12, 29) {real, imag} */,
  {32'hbe273185, 32'h3e50b578} /* (21, 12, 28) {real, imag} */,
  {32'h3d019ee2, 32'hbec1e1db} /* (21, 12, 27) {real, imag} */,
  {32'hbf38cb9c, 32'h3e3c2390} /* (21, 12, 26) {real, imag} */,
  {32'h3e9e026b, 32'hbbccf3e0} /* (21, 12, 25) {real, imag} */,
  {32'h3da81c7c, 32'h3eadca3f} /* (21, 12, 24) {real, imag} */,
  {32'h3ef6d3e8, 32'hbdb7c210} /* (21, 12, 23) {real, imag} */,
  {32'h3dcd7a84, 32'h3c4c0a0c} /* (21, 12, 22) {real, imag} */,
  {32'h3f6fbce0, 32'h3e22bd34} /* (21, 12, 21) {real, imag} */,
  {32'h3e554c5c, 32'hbf12df42} /* (21, 12, 20) {real, imag} */,
  {32'h3d9a5cd7, 32'hbd8409fe} /* (21, 12, 19) {real, imag} */,
  {32'h3e81ce7e, 32'hbee28062} /* (21, 12, 18) {real, imag} */,
  {32'h3ee22385, 32'h3eae5653} /* (21, 12, 17) {real, imag} */,
  {32'hbe51ea52, 32'h3e4f51a4} /* (21, 12, 16) {real, imag} */,
  {32'h3e5a2d46, 32'hbebb5ea0} /* (21, 12, 15) {real, imag} */,
  {32'h3e39a501, 32'h3d1eb0f8} /* (21, 12, 14) {real, imag} */,
  {32'h3e5bc5a7, 32'h3dbb9e45} /* (21, 12, 13) {real, imag} */,
  {32'h3ef54a2c, 32'h3ef0b9b0} /* (21, 12, 12) {real, imag} */,
  {32'hbf0bdb46, 32'h3d9bb139} /* (21, 12, 11) {real, imag} */,
  {32'hbdafe40e, 32'h3e6b3ab6} /* (21, 12, 10) {real, imag} */,
  {32'h3e5a209b, 32'hbe6fd856} /* (21, 12, 9) {real, imag} */,
  {32'hbec3acc6, 32'h3eb351a6} /* (21, 12, 8) {real, imag} */,
  {32'hbf2023c8, 32'h3db72dbc} /* (21, 12, 7) {real, imag} */,
  {32'h3e8e0ffa, 32'h3dbb274c} /* (21, 12, 6) {real, imag} */,
  {32'h3e83ad56, 32'hbd9a7554} /* (21, 12, 5) {real, imag} */,
  {32'h3e888516, 32'hbdc4c705} /* (21, 12, 4) {real, imag} */,
  {32'hbe55dadd, 32'h3e22dad7} /* (21, 12, 3) {real, imag} */,
  {32'h3dd416f6, 32'hbe4470b4} /* (21, 12, 2) {real, imag} */,
  {32'h3dd0d53d, 32'hbe228556} /* (21, 12, 1) {real, imag} */,
  {32'h3f49bc09, 32'h3ea9d1c4} /* (21, 12, 0) {real, imag} */,
  {32'h3ea01852, 32'h3de9af7e} /* (21, 11, 31) {real, imag} */,
  {32'hbf4ade5b, 32'h3d9c217d} /* (21, 11, 30) {real, imag} */,
  {32'h3d91d856, 32'h3e00797b} /* (21, 11, 29) {real, imag} */,
  {32'hbf273d46, 32'h3e0f4f5f} /* (21, 11, 28) {real, imag} */,
  {32'hbda072f2, 32'h3eb0e5fe} /* (21, 11, 27) {real, imag} */,
  {32'hbef904e3, 32'hbe4d8ff0} /* (21, 11, 26) {real, imag} */,
  {32'hbe7a8bf8, 32'h3de00e0c} /* (21, 11, 25) {real, imag} */,
  {32'h3ea5f604, 32'hbde6f3b2} /* (21, 11, 24) {real, imag} */,
  {32'h3d079a6c, 32'hbd424928} /* (21, 11, 23) {real, imag} */,
  {32'h3ed79ee8, 32'hbe78d3b0} /* (21, 11, 22) {real, imag} */,
  {32'hbe7ccd98, 32'h3e9b2a41} /* (21, 11, 21) {real, imag} */,
  {32'h3e321faa, 32'h3c4e1ec0} /* (21, 11, 20) {real, imag} */,
  {32'h3eb4ea39, 32'h3e6f7f97} /* (21, 11, 19) {real, imag} */,
  {32'h3ee84bbe, 32'hbf113ff1} /* (21, 11, 18) {real, imag} */,
  {32'hbe03a6ec, 32'hbe2f1030} /* (21, 11, 17) {real, imag} */,
  {32'hbedcaec6, 32'h3e9c11e5} /* (21, 11, 16) {real, imag} */,
  {32'h3d883876, 32'hbe84a76e} /* (21, 11, 15) {real, imag} */,
  {32'h3b789b40, 32'h3e16a9c6} /* (21, 11, 14) {real, imag} */,
  {32'hbd997313, 32'h3de049f6} /* (21, 11, 13) {real, imag} */,
  {32'hbec4da70, 32'h3eabc2bd} /* (21, 11, 12) {real, imag} */,
  {32'hbf064264, 32'hbca99afc} /* (21, 11, 11) {real, imag} */,
  {32'h3e0a3b45, 32'hbd5722d8} /* (21, 11, 10) {real, imag} */,
  {32'h3ecbaa62, 32'hbe9a7108} /* (21, 11, 9) {real, imag} */,
  {32'h3eedbfbf, 32'hbb5c8180} /* (21, 11, 8) {real, imag} */,
  {32'h3e91a605, 32'hbd4bac38} /* (21, 11, 7) {real, imag} */,
  {32'h3ec5a0c2, 32'h3e6652a7} /* (21, 11, 6) {real, imag} */,
  {32'h3ed35014, 32'hbd54a4b0} /* (21, 11, 5) {real, imag} */,
  {32'hbe95f8b0, 32'h3e0c445e} /* (21, 11, 4) {real, imag} */,
  {32'h3eb31ef5, 32'hbf038600} /* (21, 11, 3) {real, imag} */,
  {32'h3e78aa08, 32'hbea54854} /* (21, 11, 2) {real, imag} */,
  {32'h3d7a5853, 32'h3f19bf30} /* (21, 11, 1) {real, imag} */,
  {32'h3ebecdfb, 32'h3f2917ed} /* (21, 11, 0) {real, imag} */,
  {32'h3ebd8b1c, 32'hbf760b3e} /* (21, 10, 31) {real, imag} */,
  {32'h3ed1c0ef, 32'h3f289d7b} /* (21, 10, 30) {real, imag} */,
  {32'h3dbc7839, 32'hbd2de910} /* (21, 10, 29) {real, imag} */,
  {32'hbea29643, 32'h3dddb6ef} /* (21, 10, 28) {real, imag} */,
  {32'h3e906aeb, 32'h3e24f73b} /* (21, 10, 27) {real, imag} */,
  {32'h3ea03376, 32'h3ebe7db1} /* (21, 10, 26) {real, imag} */,
  {32'hbf0b2b00, 32'hbdead684} /* (21, 10, 25) {real, imag} */,
  {32'h3eafb52a, 32'h3e26163e} /* (21, 10, 24) {real, imag} */,
  {32'hbed39aa6, 32'hbe463d94} /* (21, 10, 23) {real, imag} */,
  {32'h3bdd9fb0, 32'hbe8d12f5} /* (21, 10, 22) {real, imag} */,
  {32'h3f224b53, 32'hbe7abfb4} /* (21, 10, 21) {real, imag} */,
  {32'hbc94d074, 32'hbeefb11a} /* (21, 10, 20) {real, imag} */,
  {32'hbe5cbcd7, 32'hbe04ae55} /* (21, 10, 19) {real, imag} */,
  {32'h3a781c40, 32'hbe71a102} /* (21, 10, 18) {real, imag} */,
  {32'hbe91b11a, 32'h3ecb3cc0} /* (21, 10, 17) {real, imag} */,
  {32'h3f090f35, 32'hbe53e9ba} /* (21, 10, 16) {real, imag} */,
  {32'h3e48acb2, 32'hbc4bd1d0} /* (21, 10, 15) {real, imag} */,
  {32'hbd6102ce, 32'hbe469c80} /* (21, 10, 14) {real, imag} */,
  {32'hbde85b45, 32'hbd428370} /* (21, 10, 13) {real, imag} */,
  {32'hbdb8167c, 32'h3f0d67e8} /* (21, 10, 12) {real, imag} */,
  {32'hbde1d9e0, 32'h3d8c6cec} /* (21, 10, 11) {real, imag} */,
  {32'h3ed2a866, 32'h3eefb632} /* (21, 10, 10) {real, imag} */,
  {32'hbd33ded0, 32'hbd3ab364} /* (21, 10, 9) {real, imag} */,
  {32'hbe742492, 32'hbe8457b8} /* (21, 10, 8) {real, imag} */,
  {32'hbe7fe706, 32'h3dee3219} /* (21, 10, 7) {real, imag} */,
  {32'h3edc72fa, 32'hbf036d7c} /* (21, 10, 6) {real, imag} */,
  {32'hbef3fd64, 32'hbee80ed3} /* (21, 10, 5) {real, imag} */,
  {32'h3dd41328, 32'h3ec5d2b8} /* (21, 10, 4) {real, imag} */,
  {32'h3d7b40cc, 32'hbc96cf28} /* (21, 10, 3) {real, imag} */,
  {32'h3e591e1a, 32'hbd369548} /* (21, 10, 2) {real, imag} */,
  {32'hbf70e694, 32'hbee93db2} /* (21, 10, 1) {real, imag} */,
  {32'hbf5ad4c8, 32'hbe4ac227} /* (21, 10, 0) {real, imag} */,
  {32'h3ef1b561, 32'h3efe8fca} /* (21, 9, 31) {real, imag} */,
  {32'hbdf6b3be, 32'h3e9d2e84} /* (21, 9, 30) {real, imag} */,
  {32'hbea6acbc, 32'hbef48036} /* (21, 9, 29) {real, imag} */,
  {32'hbd5625e8, 32'hbf1cf116} /* (21, 9, 28) {real, imag} */,
  {32'h3dce0378, 32'hbe56bc65} /* (21, 9, 27) {real, imag} */,
  {32'hbdf84c4c, 32'h3d377e14} /* (21, 9, 26) {real, imag} */,
  {32'hbe4ae2a4, 32'h3e1009c5} /* (21, 9, 25) {real, imag} */,
  {32'hbe0f7c11, 32'h3f052dbd} /* (21, 9, 24) {real, imag} */,
  {32'hbc9f4ce4, 32'hbb8e1080} /* (21, 9, 23) {real, imag} */,
  {32'hbe33ce7f, 32'hbf07346a} /* (21, 9, 22) {real, imag} */,
  {32'hbe8307d3, 32'h3dba3544} /* (21, 9, 21) {real, imag} */,
  {32'h3d8e5c44, 32'h3e1bce5e} /* (21, 9, 20) {real, imag} */,
  {32'hbd8c7c80, 32'hbda45668} /* (21, 9, 19) {real, imag} */,
  {32'h3ea5d6c7, 32'h3de8cd36} /* (21, 9, 18) {real, imag} */,
  {32'hbe0b4b3c, 32'hbf1cc79e} /* (21, 9, 17) {real, imag} */,
  {32'hbb75cd40, 32'h3e11f94f} /* (21, 9, 16) {real, imag} */,
  {32'h3e07eb8a, 32'hbdc02015} /* (21, 9, 15) {real, imag} */,
  {32'h3c1be448, 32'h3ebab478} /* (21, 9, 14) {real, imag} */,
  {32'hbe2c8392, 32'h3e60bb37} /* (21, 9, 13) {real, imag} */,
  {32'hbf25acbf, 32'h3dd41d60} /* (21, 9, 12) {real, imag} */,
  {32'h3c211430, 32'h3ee3c516} /* (21, 9, 11) {real, imag} */,
  {32'h3e9e3e20, 32'hbe5701c7} /* (21, 9, 10) {real, imag} */,
  {32'h3f34f97a, 32'hbe551398} /* (21, 9, 9) {real, imag} */,
  {32'hbefb1608, 32'h3e4ae552} /* (21, 9, 8) {real, imag} */,
  {32'h3e415b7c, 32'hbf223ddc} /* (21, 9, 7) {real, imag} */,
  {32'hbec96e07, 32'hbf516a40} /* (21, 9, 6) {real, imag} */,
  {32'h3f3dea61, 32'h3e289747} /* (21, 9, 5) {real, imag} */,
  {32'hbef36f04, 32'h3d9dd7ef} /* (21, 9, 4) {real, imag} */,
  {32'h3ed28adf, 32'hbeb1aa87} /* (21, 9, 3) {real, imag} */,
  {32'hbd082fbc, 32'h3eb2c967} /* (21, 9, 2) {real, imag} */,
  {32'hbf2c64f8, 32'hbdbde9dc} /* (21, 9, 1) {real, imag} */,
  {32'h3f06b3e3, 32'h3ea28e66} /* (21, 9, 0) {real, imag} */,
  {32'h3f956bc1, 32'h3f852325} /* (21, 8, 31) {real, imag} */,
  {32'hbf3b04cd, 32'hbed1d501} /* (21, 8, 30) {real, imag} */,
  {32'h3e8451b2, 32'h3cfc6b18} /* (21, 8, 29) {real, imag} */,
  {32'h3df5ec40, 32'h3e93132b} /* (21, 8, 28) {real, imag} */,
  {32'hbf54a9fe, 32'hbf11bb49} /* (21, 8, 27) {real, imag} */,
  {32'h3f73339a, 32'hbbe41a00} /* (21, 8, 26) {real, imag} */,
  {32'h3e7742b3, 32'hbdf803d0} /* (21, 8, 25) {real, imag} */,
  {32'hbe198693, 32'hbf028a0c} /* (21, 8, 24) {real, imag} */,
  {32'h3e9c3a13, 32'h3e9e78b7} /* (21, 8, 23) {real, imag} */,
  {32'hbb878d80, 32'hbdbab0d8} /* (21, 8, 22) {real, imag} */,
  {32'hbdf09a8e, 32'h3f495788} /* (21, 8, 21) {real, imag} */,
  {32'h3e23eb8b, 32'h3d3fc9b4} /* (21, 8, 20) {real, imag} */,
  {32'h3de2e398, 32'hbed41651} /* (21, 8, 19) {real, imag} */,
  {32'hbdd0c5dc, 32'h3eaa805a} /* (21, 8, 18) {real, imag} */,
  {32'h3d84d4cc, 32'h3c977110} /* (21, 8, 17) {real, imag} */,
  {32'h3d07269c, 32'hbe0a9782} /* (21, 8, 16) {real, imag} */,
  {32'hbe5d22dc, 32'h3e2c4711} /* (21, 8, 15) {real, imag} */,
  {32'hbe6bb5b3, 32'h3d851572} /* (21, 8, 14) {real, imag} */,
  {32'h3c90f380, 32'hbe781da0} /* (21, 8, 13) {real, imag} */,
  {32'h3e44c29a, 32'hbeb4c39a} /* (21, 8, 12) {real, imag} */,
  {32'hbba99a40, 32'hbf49d051} /* (21, 8, 11) {real, imag} */,
  {32'hbf0db8f6, 32'h3f42438e} /* (21, 8, 10) {real, imag} */,
  {32'hbd71f840, 32'hbd8c10d8} /* (21, 8, 9) {real, imag} */,
  {32'hbcca14e0, 32'h3d8cafc2} /* (21, 8, 8) {real, imag} */,
  {32'hbd9552f4, 32'hbe4aac96} /* (21, 8, 7) {real, imag} */,
  {32'h3db5b7cc, 32'h3cabac00} /* (21, 8, 6) {real, imag} */,
  {32'hbf887754, 32'hbdeac1d4} /* (21, 8, 5) {real, imag} */,
  {32'h3f0738b9, 32'hbdfbc962} /* (21, 8, 4) {real, imag} */,
  {32'h3ef20080, 32'hbe60fefd} /* (21, 8, 3) {real, imag} */,
  {32'hbf1bbb3f, 32'hbe6784d0} /* (21, 8, 2) {real, imag} */,
  {32'h3f186e44, 32'h3ec9bbf2} /* (21, 8, 1) {real, imag} */,
  {32'h3e9e3e58, 32'hbe424b1c} /* (21, 8, 0) {real, imag} */,
  {32'h3c523780, 32'hbee7c94c} /* (21, 7, 31) {real, imag} */,
  {32'h3f0d938f, 32'hbf47321b} /* (21, 7, 30) {real, imag} */,
  {32'h3dd9f536, 32'hbe088e9b} /* (21, 7, 29) {real, imag} */,
  {32'h3f1e85c6, 32'h3e00a594} /* (21, 7, 28) {real, imag} */,
  {32'hbeb75d73, 32'h3e201ec5} /* (21, 7, 27) {real, imag} */,
  {32'hbe9b75ba, 32'h3f3209f8} /* (21, 7, 26) {real, imag} */,
  {32'hbeae164c, 32'h3ee0b147} /* (21, 7, 25) {real, imag} */,
  {32'hbe1a5dd2, 32'h3f012ca6} /* (21, 7, 24) {real, imag} */,
  {32'hbe174642, 32'hbe41b15f} /* (21, 7, 23) {real, imag} */,
  {32'hbf1df8cb, 32'h3e2a2584} /* (21, 7, 22) {real, imag} */,
  {32'h3cc43f28, 32'hbf1437f4} /* (21, 7, 21) {real, imag} */,
  {32'hbe177cb0, 32'hbc3dbeac} /* (21, 7, 20) {real, imag} */,
  {32'h3dbb437c, 32'h3ebcbfeb} /* (21, 7, 19) {real, imag} */,
  {32'h3d704e38, 32'hbe330e13} /* (21, 7, 18) {real, imag} */,
  {32'hbe9b595c, 32'h3e13efb4} /* (21, 7, 17) {real, imag} */,
  {32'hbde39f69, 32'hbed0b56d} /* (21, 7, 16) {real, imag} */,
  {32'h3c09fca4, 32'h3db591fe} /* (21, 7, 15) {real, imag} */,
  {32'hbeed2434, 32'h3dc0cdb8} /* (21, 7, 14) {real, imag} */,
  {32'hbd92808e, 32'h3e4ae15b} /* (21, 7, 13) {real, imag} */,
  {32'hbe043ab3, 32'hbe4be7ea} /* (21, 7, 12) {real, imag} */,
  {32'hbf2f4b36, 32'h3ee2ea48} /* (21, 7, 11) {real, imag} */,
  {32'hbe4d5d66, 32'hbe510976} /* (21, 7, 10) {real, imag} */,
  {32'hbe14d9b7, 32'h3dc7f028} /* (21, 7, 9) {real, imag} */,
  {32'hbe7139bd, 32'h3c3eeef8} /* (21, 7, 8) {real, imag} */,
  {32'hbf3968ae, 32'hbcf55d90} /* (21, 7, 7) {real, imag} */,
  {32'hbe630ddf, 32'h3f15c674} /* (21, 7, 6) {real, imag} */,
  {32'h3f55ed6c, 32'hbe85035a} /* (21, 7, 5) {real, imag} */,
  {32'h3c4e6d40, 32'hbeb5830d} /* (21, 7, 4) {real, imag} */,
  {32'h3f56105b, 32'h3ee26cce} /* (21, 7, 3) {real, imag} */,
  {32'h3e9c4d14, 32'h3e5ef07c} /* (21, 7, 2) {real, imag} */,
  {32'h3e505b28, 32'hbde05b6f} /* (21, 7, 1) {real, imag} */,
  {32'hbf46c9e7, 32'hbf6c1c8e} /* (21, 7, 0) {real, imag} */,
  {32'hbe8be10a, 32'h3f829357} /* (21, 6, 31) {real, imag} */,
  {32'h3d05c200, 32'hbe070388} /* (21, 6, 30) {real, imag} */,
  {32'h3e7e0aa5, 32'h3e04667a} /* (21, 6, 29) {real, imag} */,
  {32'h3f2de48c, 32'hbf20a7f5} /* (21, 6, 28) {real, imag} */,
  {32'hbe7e644c, 32'hbf3aaf9d} /* (21, 6, 27) {real, imag} */,
  {32'h3eca7d0e, 32'hbf02638a} /* (21, 6, 26) {real, imag} */,
  {32'hbe1f4018, 32'hbea1a559} /* (21, 6, 25) {real, imag} */,
  {32'hbe8009c6, 32'h3e66a97b} /* (21, 6, 24) {real, imag} */,
  {32'hbe8dd212, 32'h3ef7ff78} /* (21, 6, 23) {real, imag} */,
  {32'h3d9c7640, 32'hbeb69056} /* (21, 6, 22) {real, imag} */,
  {32'hbe6038eb, 32'hbd660c80} /* (21, 6, 21) {real, imag} */,
  {32'hbeec2d95, 32'hbc354f10} /* (21, 6, 20) {real, imag} */,
  {32'hbe8adb2e, 32'hbeaa702b} /* (21, 6, 19) {real, imag} */,
  {32'hbe03c696, 32'h3efdb580} /* (21, 6, 18) {real, imag} */,
  {32'h3f0630e9, 32'h3e6e77d2} /* (21, 6, 17) {real, imag} */,
  {32'hbe423fd4, 32'hbe562aad} /* (21, 6, 16) {real, imag} */,
  {32'h3af40f60, 32'h3d796d5e} /* (21, 6, 15) {real, imag} */,
  {32'h3e4125ea, 32'h3e18adb0} /* (21, 6, 14) {real, imag} */,
  {32'hbd2d5b67, 32'hbef3bb01} /* (21, 6, 13) {real, imag} */,
  {32'hbe9b616e, 32'h3e05f412} /* (21, 6, 12) {real, imag} */,
  {32'hbf11e8c2, 32'hbf0066cb} /* (21, 6, 11) {real, imag} */,
  {32'h3bd6bf00, 32'h3f18492c} /* (21, 6, 10) {real, imag} */,
  {32'h3cc64030, 32'h3ee2f9c7} /* (21, 6, 9) {real, imag} */,
  {32'hbe052d8a, 32'hbf2f788c} /* (21, 6, 8) {real, imag} */,
  {32'hbe765d1e, 32'hbd95ea8a} /* (21, 6, 7) {real, imag} */,
  {32'hbed0a914, 32'hbf10b2ee} /* (21, 6, 6) {real, imag} */,
  {32'hbf387360, 32'h3e3ee95d} /* (21, 6, 5) {real, imag} */,
  {32'hbe0c1600, 32'h3d9647d1} /* (21, 6, 4) {real, imag} */,
  {32'h3f1b20b3, 32'hbf250a81} /* (21, 6, 3) {real, imag} */,
  {32'h3e0e3884, 32'h3f383a26} /* (21, 6, 2) {real, imag} */,
  {32'hbdd0f7c8, 32'h3eac6f77} /* (21, 6, 1) {real, imag} */,
  {32'hbe533a47, 32'h3e15f1e1} /* (21, 6, 0) {real, imag} */,
  {32'h403d67e2, 32'h3ee18323} /* (21, 5, 31) {real, imag} */,
  {32'hbf83cf70, 32'hbed3c5f0} /* (21, 5, 30) {real, imag} */,
  {32'h3d674b80, 32'h3ecf53e4} /* (21, 5, 29) {real, imag} */,
  {32'h3f15423c, 32'hbe62c888} /* (21, 5, 28) {real, imag} */,
  {32'hbf738dee, 32'hbdc7c98c} /* (21, 5, 27) {real, imag} */,
  {32'hbf59b72e, 32'h3db7449e} /* (21, 5, 26) {real, imag} */,
  {32'h3e8d6142, 32'h3d28dfde} /* (21, 5, 25) {real, imag} */,
  {32'hbe2a8644, 32'h3e247504} /* (21, 5, 24) {real, imag} */,
  {32'h3d75a488, 32'h3e532f05} /* (21, 5, 23) {real, imag} */,
  {32'hbe3d7857, 32'hbac04700} /* (21, 5, 22) {real, imag} */,
  {32'hbc50e568, 32'hbe57b5ce} /* (21, 5, 21) {real, imag} */,
  {32'h3ea5506a, 32'h3e82bb36} /* (21, 5, 20) {real, imag} */,
  {32'hbd8e23e8, 32'h3d6db4dc} /* (21, 5, 19) {real, imag} */,
  {32'hbd449b52, 32'h3de0551e} /* (21, 5, 18) {real, imag} */,
  {32'h3e2b4179, 32'hbe9c60db} /* (21, 5, 17) {real, imag} */,
  {32'hbe2c0092, 32'h3dcb97be} /* (21, 5, 16) {real, imag} */,
  {32'hbe4ee78c, 32'h3b369a00} /* (21, 5, 15) {real, imag} */,
  {32'hbe933b91, 32'hbda13344} /* (21, 5, 14) {real, imag} */,
  {32'h3e262d48, 32'hbcaa5670} /* (21, 5, 13) {real, imag} */,
  {32'hbe2a43d0, 32'hbe840ba6} /* (21, 5, 12) {real, imag} */,
  {32'hbe8f9e70, 32'hbf12d404} /* (21, 5, 11) {real, imag} */,
  {32'h3e867b40, 32'h3e47d274} /* (21, 5, 10) {real, imag} */,
  {32'h3e7e9a15, 32'hbefa41a2} /* (21, 5, 9) {real, imag} */,
  {32'hbe4da84b, 32'hbdc12ed0} /* (21, 5, 8) {real, imag} */,
  {32'h3f874d8c, 32'h3ecd9639} /* (21, 5, 7) {real, imag} */,
  {32'h3e79787c, 32'hbea36fe8} /* (21, 5, 6) {real, imag} */,
  {32'hbf139dd8, 32'hbf01563d} /* (21, 5, 5) {real, imag} */,
  {32'hbee3baf0, 32'h3f14d418} /* (21, 5, 4) {real, imag} */,
  {32'h3e923773, 32'h3e94306c} /* (21, 5, 3) {real, imag} */,
  {32'hbeff4f69, 32'hbfbca04f} /* (21, 5, 2) {real, imag} */,
  {32'h4001da38, 32'h400106c8} /* (21, 5, 1) {real, imag} */,
  {32'h3f962774, 32'h4015cd98} /* (21, 5, 0) {real, imag} */,
  {32'hbf76f992, 32'hc059fc9f} /* (21, 4, 31) {real, imag} */,
  {32'h4041bff3, 32'h3fe864da} /* (21, 4, 30) {real, imag} */,
  {32'h3e3570c2, 32'h3c145e20} /* (21, 4, 29) {real, imag} */,
  {32'hbf126db6, 32'h3f3739ac} /* (21, 4, 28) {real, imag} */,
  {32'h3ddffa2e, 32'hbf47ef34} /* (21, 4, 27) {real, imag} */,
  {32'h3ea04934, 32'hbf2774f2} /* (21, 4, 26) {real, imag} */,
  {32'h3e96f032, 32'h3f1d6c32} /* (21, 4, 25) {real, imag} */,
  {32'h3ecf046c, 32'h3e753f05} /* (21, 4, 24) {real, imag} */,
  {32'hbe950669, 32'hbe063eb5} /* (21, 4, 23) {real, imag} */,
  {32'hbe957701, 32'h3d9548d7} /* (21, 4, 22) {real, imag} */,
  {32'hbf0c8005, 32'hbe855968} /* (21, 4, 21) {real, imag} */,
  {32'h3f0a8a6d, 32'h3f0f7464} /* (21, 4, 20) {real, imag} */,
  {32'hbe41e5b0, 32'h3f1a8f9a} /* (21, 4, 19) {real, imag} */,
  {32'h3f0a62ac, 32'h3ee02be6} /* (21, 4, 18) {real, imag} */,
  {32'h3d31349c, 32'h3dd29ae4} /* (21, 4, 17) {real, imag} */,
  {32'hbe3700a2, 32'h3d5dcf24} /* (21, 4, 16) {real, imag} */,
  {32'h3dca15a4, 32'hbbc53428} /* (21, 4, 15) {real, imag} */,
  {32'h3baaf9e0, 32'hbe81ceea} /* (21, 4, 14) {real, imag} */,
  {32'hbe8e3c3a, 32'hbf315bb6} /* (21, 4, 13) {real, imag} */,
  {32'hbe639be7, 32'h3d375a0f} /* (21, 4, 12) {real, imag} */,
  {32'h3f18bac7, 32'h3e079407} /* (21, 4, 11) {real, imag} */,
  {32'h3e1cdff2, 32'hbe0616f5} /* (21, 4, 10) {real, imag} */,
  {32'h3dba87e8, 32'h3d614bb4} /* (21, 4, 9) {real, imag} */,
  {32'h3f319a4d, 32'h3ebb8a99} /* (21, 4, 8) {real, imag} */,
  {32'hbf10d2e4, 32'h3e1e8fe7} /* (21, 4, 7) {real, imag} */,
  {32'hbd0863c8, 32'h3d182d08} /* (21, 4, 6) {real, imag} */,
  {32'h3f3cfe58, 32'h3e90531e} /* (21, 4, 5) {real, imag} */,
  {32'h3f4f7a63, 32'hbf8587ad} /* (21, 4, 4) {real, imag} */,
  {32'hbdeaabe0, 32'hbf98af4a} /* (21, 4, 3) {real, imag} */,
  {32'h40736fd0, 32'h3ff0705c} /* (21, 4, 2) {real, imag} */,
  {32'hc08e25c0, 32'hbfec4de8} /* (21, 4, 1) {real, imag} */,
  {32'hc003df29, 32'h3fa80a95} /* (21, 4, 0) {real, imag} */,
  {32'h4093f214, 32'hc02111e1} /* (21, 3, 31) {real, imag} */,
  {32'hc04f5563, 32'h4045f0e9} /* (21, 3, 30) {real, imag} */,
  {32'hbe9a8dcb, 32'h3df924b9} /* (21, 3, 29) {real, imag} */,
  {32'hbfc47536, 32'hbf9809de} /* (21, 3, 28) {real, imag} */,
  {32'h3effad59, 32'hbdf20d54} /* (21, 3, 27) {real, imag} */,
  {32'h3e8e44fc, 32'hbf5a7e81} /* (21, 3, 26) {real, imag} */,
  {32'hbf53e032, 32'hbe1bda4a} /* (21, 3, 25) {real, imag} */,
  {32'h3f36d850, 32'h3e5d6283} /* (21, 3, 24) {real, imag} */,
  {32'hbd152e9c, 32'hbf2d83df} /* (21, 3, 23) {real, imag} */,
  {32'hbe6fc6db, 32'hbf4b9a10} /* (21, 3, 22) {real, imag} */,
  {32'h3eb1061a, 32'h3f200dd0} /* (21, 3, 21) {real, imag} */,
  {32'h3f0a5966, 32'h3f15f017} /* (21, 3, 20) {real, imag} */,
  {32'h3efcfb7d, 32'hbe9d4fff} /* (21, 3, 19) {real, imag} */,
  {32'hbe61615e, 32'hbec73e02} /* (21, 3, 18) {real, imag} */,
  {32'h3cf6f1b8, 32'h3d28d270} /* (21, 3, 17) {real, imag} */,
  {32'h3f0005d1, 32'h3daf0124} /* (21, 3, 16) {real, imag} */,
  {32'h3e9a784b, 32'h3c865550} /* (21, 3, 15) {real, imag} */,
  {32'hbc7c3aa0, 32'h3ec73263} /* (21, 3, 14) {real, imag} */,
  {32'h3dcfdacc, 32'hbca3a002} /* (21, 3, 13) {real, imag} */,
  {32'hbd373850, 32'h3eab0e13} /* (21, 3, 12) {real, imag} */,
  {32'hbdee3a9a, 32'h3e3f8c20} /* (21, 3, 11) {real, imag} */,
  {32'h3e51a864, 32'h3ebd6069} /* (21, 3, 10) {real, imag} */,
  {32'hbf5a58ce, 32'h3d6c76c4} /* (21, 3, 9) {real, imag} */,
  {32'hbf03c27e, 32'h3ed92208} /* (21, 3, 8) {real, imag} */,
  {32'h3f1dc7dc, 32'hbeb52d3f} /* (21, 3, 7) {real, imag} */,
  {32'hbd249684, 32'hbd9a418a} /* (21, 3, 6) {real, imag} */,
  {32'hbe8b83c6, 32'hbde39be2} /* (21, 3, 5) {real, imag} */,
  {32'h3fb12b07, 32'hbfb24670} /* (21, 3, 4) {real, imag} */,
  {32'h3fcac748, 32'h3e9a2c5a} /* (21, 3, 3) {real, imag} */,
  {32'hbe852833, 32'h406586ac} /* (21, 3, 2) {real, imag} */,
  {32'hc088adde, 32'hc037548c} /* (21, 3, 1) {real, imag} */,
  {32'h3fc0fea0, 32'h3eb207d2} /* (21, 3, 0) {real, imag} */,
  {32'h42246bad, 32'h3f075c0a} /* (21, 2, 31) {real, imag} */,
  {32'hc1943477, 32'h40e680f3} /* (21, 2, 30) {real, imag} */,
  {32'hbca50508, 32'h3e6d6e25} /* (21, 2, 29) {real, imag} */,
  {32'h3e232870, 32'hbffe464c} /* (21, 2, 28) {real, imag} */,
  {32'hbfa76feb, 32'h3f6ac712} /* (21, 2, 27) {real, imag} */,
  {32'hbd3db5d8, 32'h3ee74c88} /* (21, 2, 26) {real, imag} */,
  {32'h3f40fc76, 32'hbf1a725e} /* (21, 2, 25) {real, imag} */,
  {32'hbf790397, 32'h3fbaeb5f} /* (21, 2, 24) {real, imag} */,
  {32'hbeed993a, 32'h3da33836} /* (21, 2, 23) {real, imag} */,
  {32'hbee0899b, 32'hbc00c098} /* (21, 2, 22) {real, imag} */,
  {32'h3d3ad3fc, 32'h3e1abe48} /* (21, 2, 21) {real, imag} */,
  {32'h3e93a82e, 32'hbe149d28} /* (21, 2, 20) {real, imag} */,
  {32'hbd97e177, 32'hbe061f04} /* (21, 2, 19) {real, imag} */,
  {32'hbf1d12a0, 32'h3e4620c8} /* (21, 2, 18) {real, imag} */,
  {32'h3d0e6650, 32'hbec1acdc} /* (21, 2, 17) {real, imag} */,
  {32'hbe80017b, 32'h3d373352} /* (21, 2, 16) {real, imag} */,
  {32'hbdd3f85c, 32'h3e34ccda} /* (21, 2, 15) {real, imag} */,
  {32'h3e62beec, 32'hbf415f93} /* (21, 2, 14) {real, imag} */,
  {32'hbe1167ec, 32'h3ea0187a} /* (21, 2, 13) {real, imag} */,
  {32'h3e85be9e, 32'h3d98c694} /* (21, 2, 12) {real, imag} */,
  {32'h3c9ecd74, 32'hbf119470} /* (21, 2, 11) {real, imag} */,
  {32'h3eb76366, 32'hbdfcbe30} /* (21, 2, 10) {real, imag} */,
  {32'h3ee83a34, 32'hbe26cceb} /* (21, 2, 9) {real, imag} */,
  {32'hbef29192, 32'hbf764f98} /* (21, 2, 8) {real, imag} */,
  {32'h3d68248e, 32'hbeb86ddf} /* (21, 2, 7) {real, imag} */,
  {32'h3dfb8667, 32'h3eb2b07d} /* (21, 2, 6) {real, imag} */,
  {32'hc02dfe11, 32'hbfe9ac94} /* (21, 2, 5) {real, imag} */,
  {32'h40442db8, 32'h3f283ce5} /* (21, 2, 4) {real, imag} */,
  {32'h3dd090d0, 32'hbf558fc4} /* (21, 2, 3) {real, imag} */,
  {32'hc1492148, 32'h403bd477} /* (21, 2, 2) {real, imag} */,
  {32'h41c3ca46, 32'hc0546b7e} /* (21, 2, 1) {real, imag} */,
  {32'h41a4705c, 32'h40873b9c} /* (21, 2, 0) {real, imag} */,
  {32'hc2615558, 32'h4173fda5} /* (21, 1, 31) {real, imag} */,
  {32'h417436ba, 32'h3f2b5ccb} /* (21, 1, 30) {real, imag} */,
  {32'h3df047d0, 32'hbfe920f2} /* (21, 1, 29) {real, imag} */,
  {32'hc05c6d9a, 32'hc049a8ce} /* (21, 1, 28) {real, imag} */,
  {32'h40876ed6, 32'hbee832f8} /* (21, 1, 27) {real, imag} */,
  {32'h3e934a2f, 32'hbf60eaff} /* (21, 1, 26) {real, imag} */,
  {32'h3e3c3e07, 32'hbf166f83} /* (21, 1, 25) {real, imag} */,
  {32'h3dca2924, 32'hbf080721} /* (21, 1, 24) {real, imag} */,
  {32'h3f287ea4, 32'hbef6d706} /* (21, 1, 23) {real, imag} */,
  {32'h3f7fed07, 32'hbdd4a3f8} /* (21, 1, 22) {real, imag} */,
  {32'h3f7002f3, 32'h3e528a8b} /* (21, 1, 21) {real, imag} */,
  {32'h3ebec4fc, 32'h3db892db} /* (21, 1, 20) {real, imag} */,
  {32'hbd34d968, 32'hbeaac105} /* (21, 1, 19) {real, imag} */,
  {32'h3e0bc460, 32'h3e221341} /* (21, 1, 18) {real, imag} */,
  {32'h3f063785, 32'h3d05abc0} /* (21, 1, 17) {real, imag} */,
  {32'hbcd8c234, 32'hbe4da5c6} /* (21, 1, 16) {real, imag} */,
  {32'hbe07d492, 32'hbe6822ca} /* (21, 1, 15) {real, imag} */,
  {32'hbe90b2e6, 32'h3e9142ca} /* (21, 1, 14) {real, imag} */,
  {32'hbd07e6e0, 32'hbefb8434} /* (21, 1, 13) {real, imag} */,
  {32'h3dcd9fd2, 32'h3f2121f0} /* (21, 1, 12) {real, imag} */,
  {32'h3e43dd87, 32'h3f559e6a} /* (21, 1, 11) {real, imag} */,
  {32'hbef27c7c, 32'hbde7abec} /* (21, 1, 10) {real, imag} */,
  {32'h3f98a2bd, 32'h3e9d4159} /* (21, 1, 9) {real, imag} */,
  {32'h3e577b58, 32'h3fb4bb8a} /* (21, 1, 8) {real, imag} */,
  {32'h3de1fdc8, 32'hbf4e4f79} /* (21, 1, 7) {real, imag} */,
  {32'hbe95ca7d, 32'hbe57d8f4} /* (21, 1, 6) {real, imag} */,
  {32'h40054e6c, 32'h4000f509} /* (21, 1, 5) {real, imag} */,
  {32'hbf467fe8, 32'hc01162c8} /* (21, 1, 4) {real, imag} */,
  {32'h3fe163fa, 32'h3f2846d6} /* (21, 1, 3) {real, imag} */,
  {32'h418f4c17, 32'h41904db4} /* (21, 1, 2) {real, imag} */,
  {32'hc29ee7a3, 32'hc22a4da7} /* (21, 1, 1) {real, imag} */,
  {32'hc28a002c, 32'hc12856a6} /* (21, 1, 0) {real, imag} */,
  {32'hc244a908, 32'h421a1a0d} /* (21, 0, 31) {real, imag} */,
  {32'h40c3e9a1, 32'hc1210a2c} /* (21, 0, 30) {real, imag} */,
  {32'hbe31fe24, 32'hbdf38e28} /* (21, 0, 29) {real, imag} */,
  {32'hbbdd2e00, 32'hc0035dc0} /* (21, 0, 28) {real, imag} */,
  {32'h40200ea0, 32'hbe00cdd4} /* (21, 0, 27) {real, imag} */,
  {32'hbec2f0fe, 32'hbec368f9} /* (21, 0, 26) {real, imag} */,
  {32'h3eebdc93, 32'h3f68391c} /* (21, 0, 25) {real, imag} */,
  {32'h3e50c002, 32'hbf2a21d3} /* (21, 0, 24) {real, imag} */,
  {32'h3e4cff6e, 32'h3f513dec} /* (21, 0, 23) {real, imag} */,
  {32'h3ec7efb0, 32'hbeb65d92} /* (21, 0, 22) {real, imag} */,
  {32'hbee9e5da, 32'hbd5f9992} /* (21, 0, 21) {real, imag} */,
  {32'hbe7e1e0f, 32'hbecedc24} /* (21, 0, 20) {real, imag} */,
  {32'h3e361723, 32'h3d57c418} /* (21, 0, 19) {real, imag} */,
  {32'h3e362747, 32'hbe4656ad} /* (21, 0, 18) {real, imag} */,
  {32'hbebbfcb5, 32'h3da05f4e} /* (21, 0, 17) {real, imag} */,
  {32'h3ee21bba, 32'h00000000} /* (21, 0, 16) {real, imag} */,
  {32'hbebbfcb5, 32'hbda05f4e} /* (21, 0, 15) {real, imag} */,
  {32'h3e362747, 32'h3e4656ad} /* (21, 0, 14) {real, imag} */,
  {32'h3e361723, 32'hbd57c418} /* (21, 0, 13) {real, imag} */,
  {32'hbe7e1e0f, 32'h3ecedc24} /* (21, 0, 12) {real, imag} */,
  {32'hbee9e5da, 32'h3d5f9992} /* (21, 0, 11) {real, imag} */,
  {32'h3ec7efb0, 32'h3eb65d92} /* (21, 0, 10) {real, imag} */,
  {32'h3e4cff6e, 32'hbf513dec} /* (21, 0, 9) {real, imag} */,
  {32'h3e50c002, 32'h3f2a21d3} /* (21, 0, 8) {real, imag} */,
  {32'h3eebdc93, 32'hbf68391c} /* (21, 0, 7) {real, imag} */,
  {32'hbec2f0fe, 32'h3ec368f9} /* (21, 0, 6) {real, imag} */,
  {32'h40200ea0, 32'h3e00cdd4} /* (21, 0, 5) {real, imag} */,
  {32'hbbdd2e00, 32'h40035dc0} /* (21, 0, 4) {real, imag} */,
  {32'hbe31fe24, 32'h3df38e28} /* (21, 0, 3) {real, imag} */,
  {32'h40c3e9a1, 32'h41210a2c} /* (21, 0, 2) {real, imag} */,
  {32'hc244a908, 32'hc21a1a0d} /* (21, 0, 1) {real, imag} */,
  {32'hc294e715, 32'h00000000} /* (21, 0, 0) {real, imag} */,
  {32'hc29b5d9d, 32'h422444ab} /* (20, 31, 31) {real, imag} */,
  {32'h418b9b13, 32'hc194fd1c} /* (20, 31, 30) {real, imag} */,
  {32'h3fee8cc4, 32'hbf4b97e1} /* (20, 31, 29) {real, imag} */,
  {32'hbf47bd5a, 32'h4024b38c} /* (20, 31, 28) {real, imag} */,
  {32'h3ff0ad2f, 32'hbfc5485f} /* (20, 31, 27) {real, imag} */,
  {32'h3d46d2f0, 32'hbe3bc3fa} /* (20, 31, 26) {real, imag} */,
  {32'hbf9a6639, 32'h3f0c1a32} /* (20, 31, 25) {real, imag} */,
  {32'h3f0a1dde, 32'hbf6990b1} /* (20, 31, 24) {real, imag} */,
  {32'h3dccb25f, 32'h3c63c4f0} /* (20, 31, 23) {real, imag} */,
  {32'h3f3470f4, 32'hbe0a0fe3} /* (20, 31, 22) {real, imag} */,
  {32'hbe0c7bdc, 32'hbf3df1d7} /* (20, 31, 21) {real, imag} */,
  {32'hbe8e1ace, 32'hbe57b255} /* (20, 31, 20) {real, imag} */,
  {32'hbe084d52, 32'hbe80f278} /* (20, 31, 19) {real, imag} */,
  {32'h3d487e42, 32'hbed8a142} /* (20, 31, 18) {real, imag} */,
  {32'h3e7e1e08, 32'h3e0d20ab} /* (20, 31, 17) {real, imag} */,
  {32'hbc42fef8, 32'h3e051dc0} /* (20, 31, 16) {real, imag} */,
  {32'hbe4defa8, 32'h3e369388} /* (20, 31, 15) {real, imag} */,
  {32'h3e23aa64, 32'h3efa716a} /* (20, 31, 14) {real, imag} */,
  {32'h3d545798, 32'h3d2dc170} /* (20, 31, 13) {real, imag} */,
  {32'hbe5ddfab, 32'hbe1de5f7} /* (20, 31, 12) {real, imag} */,
  {32'h3eab1f1e, 32'hbe0791f8} /* (20, 31, 11) {real, imag} */,
  {32'h3e223ff6, 32'h3eef6e2e} /* (20, 31, 10) {real, imag} */,
  {32'h3bd7de40, 32'h3d9a6e88} /* (20, 31, 9) {real, imag} */,
  {32'hbe89d17b, 32'h3f42817c} /* (20, 31, 8) {real, imag} */,
  {32'hbef38d96, 32'hbf0c1ed6} /* (20, 31, 7) {real, imag} */,
  {32'h3f55c249, 32'h3ea39f03} /* (20, 31, 6) {real, imag} */,
  {32'h4087550d, 32'hbe916d18} /* (20, 31, 5) {real, imag} */,
  {32'hc0134257, 32'h4038bb86} /* (20, 31, 4) {real, imag} */,
  {32'hbf60731e, 32'h3f659471} /* (20, 31, 3) {real, imag} */,
  {32'h416dbc2f, 32'hbf1f65a7} /* (20, 31, 2) {real, imag} */,
  {32'hc25b3350, 32'hc1756ab8} /* (20, 31, 1) {real, imag} */,
  {32'hc2857347, 32'h412791d7} /* (20, 31, 0) {real, imag} */,
  {32'h41c48726, 32'h406e840f} /* (20, 30, 31) {real, imag} */,
  {32'hc150d7c1, 32'hc02ce058} /* (20, 30, 30) {real, imag} */,
  {32'h3e9c25e9, 32'h3dc395a6} /* (20, 30, 29) {real, imag} */,
  {32'h407f0aeb, 32'hbe5426f8} /* (20, 30, 28) {real, imag} */,
  {32'hc0203008, 32'h4031db17} /* (20, 30, 27) {real, imag} */,
  {32'hbe8ce8cd, 32'h3edd3819} /* (20, 30, 26) {real, imag} */,
  {32'h3e9e8ae0, 32'hbe130a32} /* (20, 30, 25) {real, imag} */,
  {32'hbf565898, 32'h3f9925f4} /* (20, 30, 24) {real, imag} */,
  {32'hbd0ac0e0, 32'hbead17b2} /* (20, 30, 23) {real, imag} */,
  {32'h3ed7d422, 32'hbebee3ac} /* (20, 30, 22) {real, imag} */,
  {32'h3ea6570a, 32'h3ea930d0} /* (20, 30, 21) {real, imag} */,
  {32'h3d5586a4, 32'hbdab00d8} /* (20, 30, 20) {real, imag} */,
  {32'hbe84a2fa, 32'h3e552e63} /* (20, 30, 19) {real, imag} */,
  {32'hbee530b4, 32'h3d88d8ac} /* (20, 30, 18) {real, imag} */,
  {32'h3eb014c1, 32'h3e6d1a6a} /* (20, 30, 17) {real, imag} */,
  {32'hbcfaeb0e, 32'h3e22dc2a} /* (20, 30, 16) {real, imag} */,
  {32'hbe7b4408, 32'h3ecf9bee} /* (20, 30, 15) {real, imag} */,
  {32'hbc716b12, 32'h3e3be3d3} /* (20, 30, 14) {real, imag} */,
  {32'hbe89cf30, 32'hbccc6fc4} /* (20, 30, 13) {real, imag} */,
  {32'h3e79e3a8, 32'h3dd43d10} /* (20, 30, 12) {real, imag} */,
  {32'h3cc91000, 32'hbee8af79} /* (20, 30, 11) {real, imag} */,
  {32'hbf0ec44e, 32'h3ed6af92} /* (20, 30, 10) {real, imag} */,
  {32'h3d1ca65c, 32'h3e48728b} /* (20, 30, 9) {real, imag} */,
  {32'hbea00584, 32'hbfa43d57} /* (20, 30, 8) {real, imag} */,
  {32'h3f01bcec, 32'h3f2f8576} /* (20, 30, 7) {real, imag} */,
  {32'h3f14ceed, 32'hbec11471} /* (20, 30, 6) {real, imag} */,
  {32'hbfe226ad, 32'hbd961cf0} /* (20, 30, 5) {real, imag} */,
  {32'h3f2a320d, 32'h3fcb2e18} /* (20, 30, 4) {real, imag} */,
  {32'h3f924ba8, 32'h3ee193bb} /* (20, 30, 3) {real, imag} */,
  {32'hc197a590, 32'hc0d7c390} /* (20, 30, 2) {real, imag} */,
  {32'h4220d4b0, 32'hbe193e6e} /* (20, 30, 1) {real, imag} */,
  {32'h41a75dce, 32'hc06cb550} /* (20, 30, 0) {real, imag} */,
  {32'hc098e2c7, 32'h402891b5} /* (20, 29, 31) {real, imag} */,
  {32'h3f48b5de, 32'hc089d2aa} /* (20, 29, 30) {real, imag} */,
  {32'h3f9f48b2, 32'hbf08b819} /* (20, 29, 29) {real, imag} */,
  {32'h3f98e171, 32'h3e858c4c} /* (20, 29, 28) {real, imag} */,
  {32'hbf214155, 32'h3ce2f0e0} /* (20, 29, 27) {real, imag} */,
  {32'h3c3fbb60, 32'h3e9544ba} /* (20, 29, 26) {real, imag} */,
  {32'h3f1d71f9, 32'hbd5d5c38} /* (20, 29, 25) {real, imag} */,
  {32'hbe81bb3a, 32'hbf0aabef} /* (20, 29, 24) {real, imag} */,
  {32'hbeff68e8, 32'h3e65a600} /* (20, 29, 23) {real, imag} */,
  {32'h3eec316a, 32'hbe82bb29} /* (20, 29, 22) {real, imag} */,
  {32'hbdbe104c, 32'hbe0d39ee} /* (20, 29, 21) {real, imag} */,
  {32'h3ece70ba, 32'hbdc4cb48} /* (20, 29, 20) {real, imag} */,
  {32'hbd9e7d7e, 32'hbe9596ec} /* (20, 29, 19) {real, imag} */,
  {32'h3e46d120, 32'h3c836050} /* (20, 29, 18) {real, imag} */,
  {32'hbe8762ae, 32'hbc7098e0} /* (20, 29, 17) {real, imag} */,
  {32'hbc47b3fa, 32'h3dafec0c} /* (20, 29, 16) {real, imag} */,
  {32'hbcb2d772, 32'h3defcf01} /* (20, 29, 15) {real, imag} */,
  {32'hbde1520e, 32'hbdb6ab12} /* (20, 29, 14) {real, imag} */,
  {32'hbe92c8d0, 32'hbe108d64} /* (20, 29, 13) {real, imag} */,
  {32'h3e234a6a, 32'hbdf7d575} /* (20, 29, 12) {real, imag} */,
  {32'hbe701982, 32'hbe22894e} /* (20, 29, 11) {real, imag} */,
  {32'hbdbdf5ce, 32'h3e2c98f4} /* (20, 29, 10) {real, imag} */,
  {32'hbd6b2830, 32'h3ec616a7} /* (20, 29, 9) {real, imag} */,
  {32'hbe5a3a72, 32'h3dd60d08} /* (20, 29, 8) {real, imag} */,
  {32'hbf428a8f, 32'hbe3b0f46} /* (20, 29, 7) {real, imag} */,
  {32'hbc966be4, 32'h3df09e5c} /* (20, 29, 6) {real, imag} */,
  {32'hbdd8f320, 32'h3e9bab82} /* (20, 29, 5) {real, imag} */,
  {32'hbf5d0ef2, 32'h3f94668c} /* (20, 29, 4) {real, imag} */,
  {32'hbf29dbc1, 32'h3e07c5f6} /* (20, 29, 3) {real, imag} */,
  {32'hc006b455, 32'hc0849385} /* (20, 29, 2) {real, imag} */,
  {32'h4068e9b9, 32'h405e163e} /* (20, 29, 1) {real, imag} */,
  {32'h3ea447d1, 32'hbef4ecd2} /* (20, 29, 0) {real, imag} */,
  {32'hc0866ec0, 32'h3ff90c92} /* (20, 28, 31) {real, imag} */,
  {32'h408011c4, 32'hc0210ec4} /* (20, 28, 30) {real, imag} */,
  {32'hbf58ac38, 32'h3fa305c0} /* (20, 28, 29) {real, imag} */,
  {32'h3d8116ac, 32'h3f09d6f4} /* (20, 28, 28) {real, imag} */,
  {32'h3f3ea895, 32'hbf6192d6} /* (20, 28, 27) {real, imag} */,
  {32'hbf057b17, 32'hbf15999a} /* (20, 28, 26) {real, imag} */,
  {32'hbe13965c, 32'h3f634184} /* (20, 28, 25) {real, imag} */,
  {32'h3d7b73e3, 32'hbbfdf100} /* (20, 28, 24) {real, imag} */,
  {32'hbc7fff20, 32'h3eaed022} /* (20, 28, 23) {real, imag} */,
  {32'hbe838bb5, 32'h3e0a5a56} /* (20, 28, 22) {real, imag} */,
  {32'hbef686de, 32'hbe78d113} /* (20, 28, 21) {real, imag} */,
  {32'hbe97bc6a, 32'hbf01bf96} /* (20, 28, 20) {real, imag} */,
  {32'h3e69202a, 32'h3c101850} /* (20, 28, 19) {real, imag} */,
  {32'hbe00aefa, 32'hbec15543} /* (20, 28, 18) {real, imag} */,
  {32'hbde1d383, 32'h3e9fb0e2} /* (20, 28, 17) {real, imag} */,
  {32'h3db57c39, 32'hbe4b8f34} /* (20, 28, 16) {real, imag} */,
  {32'hbe94ea90, 32'hbec22195} /* (20, 28, 15) {real, imag} */,
  {32'hbe87f912, 32'hbe217f4c} /* (20, 28, 14) {real, imag} */,
  {32'h3ee4f95c, 32'h3ef10963} /* (20, 28, 13) {real, imag} */,
  {32'hbe1231e4, 32'hbe6dc38c} /* (20, 28, 12) {real, imag} */,
  {32'h3ec5f0c8, 32'h3eb85300} /* (20, 28, 11) {real, imag} */,
  {32'h3e972054, 32'h3d3e34d6} /* (20, 28, 10) {real, imag} */,
  {32'hbe871c90, 32'h3e59c3c8} /* (20, 28, 9) {real, imag} */,
  {32'h3f4e0c7c, 32'h3e395d3c} /* (20, 28, 8) {real, imag} */,
  {32'h3e5f4006, 32'hbef40a7e} /* (20, 28, 7) {real, imag} */,
  {32'hbf57da59, 32'h3f67de52} /* (20, 28, 6) {real, imag} */,
  {32'h3f3765e3, 32'h3f4e5344} /* (20, 28, 5) {real, imag} */,
  {32'hbf55c348, 32'h3c6a1da8} /* (20, 28, 4) {real, imag} */,
  {32'hbd9be250, 32'hbe13553a} /* (20, 28, 3) {real, imag} */,
  {32'h40015489, 32'hc00ed1b3} /* (20, 28, 2) {real, imag} */,
  {32'hbf7c09eb, 32'h4080e973} /* (20, 28, 1) {real, imag} */,
  {32'hc0068616, 32'h3e15598b} /* (20, 28, 0) {real, imag} */,
  {32'h3f9a6ddc, 32'hc03178a3} /* (20, 27, 31) {real, imag} */,
  {32'hbf60b282, 32'h3fc99bde} /* (20, 27, 30) {real, imag} */,
  {32'h3f0625f8, 32'hbe9b65bc} /* (20, 27, 29) {real, imag} */,
  {32'h3f3d3304, 32'hbdeb6e60} /* (20, 27, 28) {real, imag} */,
  {32'hbea55955, 32'h3ebc26ca} /* (20, 27, 27) {real, imag} */,
  {32'h3f34610c, 32'h3de7c73b} /* (20, 27, 26) {real, imag} */,
  {32'h3d90dc34, 32'hbef30297} /* (20, 27, 25) {real, imag} */,
  {32'h3e9aa1d9, 32'hbe9c5f98} /* (20, 27, 24) {real, imag} */,
  {32'hbe85d81a, 32'h3f0468f1} /* (20, 27, 23) {real, imag} */,
  {32'h3ed3f76e, 32'hbec6893e} /* (20, 27, 22) {real, imag} */,
  {32'h3ec5ee58, 32'h3f4fcdd4} /* (20, 27, 21) {real, imag} */,
  {32'hbe0a4af9, 32'h3f0a0554} /* (20, 27, 20) {real, imag} */,
  {32'hbe0c5f61, 32'h3d336870} /* (20, 27, 19) {real, imag} */,
  {32'hbe190c06, 32'hbd90121c} /* (20, 27, 18) {real, imag} */,
  {32'h3db5c1a8, 32'hbd9208f5} /* (20, 27, 17) {real, imag} */,
  {32'h3da2dbc4, 32'hbe6fe0ca} /* (20, 27, 16) {real, imag} */,
  {32'hbe87e1d6, 32'hbdd2079c} /* (20, 27, 15) {real, imag} */,
  {32'hbe1e455f, 32'hbe2d570c} /* (20, 27, 14) {real, imag} */,
  {32'hbe9acfd9, 32'h3ec750d3} /* (20, 27, 13) {real, imag} */,
  {32'h3e2519d0, 32'h3d302335} /* (20, 27, 12) {real, imag} */,
  {32'h3e01416a, 32'hbdd805d9} /* (20, 27, 11) {real, imag} */,
  {32'hbf83a9a4, 32'h3d1cbb0c} /* (20, 27, 10) {real, imag} */,
  {32'hbecaae46, 32'hbe879192} /* (20, 27, 9) {real, imag} */,
  {32'hbe703c4d, 32'hbf4bfb54} /* (20, 27, 8) {real, imag} */,
  {32'hbd5ba644, 32'hbeb9b508} /* (20, 27, 7) {real, imag} */,
  {32'hbe45aa50, 32'h3d050c74} /* (20, 27, 6) {real, imag} */,
  {32'hbf2160f1, 32'h3d2d75a8} /* (20, 27, 5) {real, imag} */,
  {32'hbdbdee38, 32'hbe123b9c} /* (20, 27, 4) {real, imag} */,
  {32'h3f47ef15, 32'hbf57e91f} /* (20, 27, 3) {real, imag} */,
  {32'hbfd56600, 32'hbe3fd076} /* (20, 27, 2) {real, imag} */,
  {32'h403a0310, 32'h3de24920} /* (20, 27, 1) {real, imag} */,
  {32'h3fcaa5ed, 32'hc00a429f} /* (20, 27, 0) {real, imag} */,
  {32'hbf36c592, 32'h3be10f00} /* (20, 26, 31) {real, imag} */,
  {32'h3e645a5f, 32'hbe692969} /* (20, 26, 30) {real, imag} */,
  {32'h3e110e23, 32'h3f74a99a} /* (20, 26, 29) {real, imag} */,
  {32'hbe7fce53, 32'hbefd8094} /* (20, 26, 28) {real, imag} */,
  {32'h3e2565ee, 32'h3e7b9868} /* (20, 26, 27) {real, imag} */,
  {32'h3e0559c4, 32'h3ed35b39} /* (20, 26, 26) {real, imag} */,
  {32'hbf5075bc, 32'hbefe7a82} /* (20, 26, 25) {real, imag} */,
  {32'hbdb3aaf6, 32'h3d72ef68} /* (20, 26, 24) {real, imag} */,
  {32'hbe82f89e, 32'hbeecf436} /* (20, 26, 23) {real, imag} */,
  {32'h3b7f7b80, 32'hbe63bbb7} /* (20, 26, 22) {real, imag} */,
  {32'h3dd634a1, 32'hbd7de8e2} /* (20, 26, 21) {real, imag} */,
  {32'h3e85b0c4, 32'h3e254d4b} /* (20, 26, 20) {real, imag} */,
  {32'h3e4fc910, 32'h3f1489d4} /* (20, 26, 19) {real, imag} */,
  {32'hbeb5d137, 32'hbea8f46a} /* (20, 26, 18) {real, imag} */,
  {32'h3e2c34dc, 32'h3ea9451f} /* (20, 26, 17) {real, imag} */,
  {32'h3c0752e0, 32'h3d1f5c36} /* (20, 26, 16) {real, imag} */,
  {32'hbe04114e, 32'h3ede10e1} /* (20, 26, 15) {real, imag} */,
  {32'h3dd8208e, 32'hbe298e76} /* (20, 26, 14) {real, imag} */,
  {32'hbe8cc962, 32'h3e7dca5c} /* (20, 26, 13) {real, imag} */,
  {32'h3ef412c6, 32'hbe3cb469} /* (20, 26, 12) {real, imag} */,
  {32'hbea6caae, 32'h3e0cb0e0} /* (20, 26, 11) {real, imag} */,
  {32'hbe1890a2, 32'h3f3b9990} /* (20, 26, 10) {real, imag} */,
  {32'h3ebc6376, 32'hbf11d0f9} /* (20, 26, 9) {real, imag} */,
  {32'hbf15c302, 32'h3eb9b449} /* (20, 26, 8) {real, imag} */,
  {32'hbed83296, 32'h3ea8ae2c} /* (20, 26, 7) {real, imag} */,
  {32'h3e2d2e0f, 32'h3f0fbd76} /* (20, 26, 6) {real, imag} */,
  {32'h3cd80858, 32'h3e953ec2} /* (20, 26, 5) {real, imag} */,
  {32'h3ec383ac, 32'hbea1ed42} /* (20, 26, 4) {real, imag} */,
  {32'hbe5fb65a, 32'h3b881540} /* (20, 26, 3) {real, imag} */,
  {32'hbd962bd0, 32'h3cf56dc8} /* (20, 26, 2) {real, imag} */,
  {32'hbd739f8c, 32'hbe991200} /* (20, 26, 1) {real, imag} */,
  {32'h3f19724f, 32'h3de5857e} /* (20, 26, 0) {real, imag} */,
  {32'h3eed0924, 32'h3f1174d8} /* (20, 25, 31) {real, imag} */,
  {32'hbdca37b0, 32'hbe44d278} /* (20, 25, 30) {real, imag} */,
  {32'h3f0dde7a, 32'hbe223f08} /* (20, 25, 29) {real, imag} */,
  {32'h3f2e3b3a, 32'hbea19f87} /* (20, 25, 28) {real, imag} */,
  {32'h3d7a5e7c, 32'hbeeab43b} /* (20, 25, 27) {real, imag} */,
  {32'h3e448faa, 32'h3f148d34} /* (20, 25, 26) {real, imag} */,
  {32'hbf37ba0b, 32'hbe0fbeb4} /* (20, 25, 25) {real, imag} */,
  {32'hbe9fde34, 32'hbe6be86f} /* (20, 25, 24) {real, imag} */,
  {32'h3f006bbd, 32'h3e26c641} /* (20, 25, 23) {real, imag} */,
  {32'h3eebfdc6, 32'h3e9d07d0} /* (20, 25, 22) {real, imag} */,
  {32'hbecd1408, 32'hbe8425f6} /* (20, 25, 21) {real, imag} */,
  {32'h3e992869, 32'hbe91330f} /* (20, 25, 20) {real, imag} */,
  {32'hbdde5b02, 32'h3d26a740} /* (20, 25, 19) {real, imag} */,
  {32'hbea4b591, 32'hbe271608} /* (20, 25, 18) {real, imag} */,
  {32'hbdfc8079, 32'hbea5d4f3} /* (20, 25, 17) {real, imag} */,
  {32'h3d8ad124, 32'hbe232f4a} /* (20, 25, 16) {real, imag} */,
  {32'h3e2a63db, 32'hbe7d1d1a} /* (20, 25, 15) {real, imag} */,
  {32'h3e11360c, 32'h3e85fe47} /* (20, 25, 14) {real, imag} */,
  {32'hbd898602, 32'hbe1bc936} /* (20, 25, 13) {real, imag} */,
  {32'hbea63f12, 32'hbca17af8} /* (20, 25, 12) {real, imag} */,
  {32'hbee11412, 32'hbbd4ade0} /* (20, 25, 11) {real, imag} */,
  {32'h3e365848, 32'h3dd5844c} /* (20, 25, 10) {real, imag} */,
  {32'hbc3a6850, 32'hbecda967} /* (20, 25, 9) {real, imag} */,
  {32'h3f0aa836, 32'hbe95f140} /* (20, 25, 8) {real, imag} */,
  {32'h3cffd1e0, 32'hbf43b334} /* (20, 25, 7) {real, imag} */,
  {32'hbd0d60a7, 32'hbdc99b02} /* (20, 25, 6) {real, imag} */,
  {32'hbeadf262, 32'hbea7e1a2} /* (20, 25, 5) {real, imag} */,
  {32'hbed30690, 32'h3e9aa057} /* (20, 25, 4) {real, imag} */,
  {32'h3ed274b2, 32'h3e86fd42} /* (20, 25, 3) {real, imag} */,
  {32'hbc84b02c, 32'h3d2b59c0} /* (20, 25, 2) {real, imag} */,
  {32'hbf14538c, 32'h3f847887} /* (20, 25, 1) {real, imag} */,
  {32'hbe6b5726, 32'h3eac5a7c} /* (20, 25, 0) {real, imag} */,
  {32'h3f328eb0, 32'hbf3d2269} /* (20, 24, 31) {real, imag} */,
  {32'hbf9bd865, 32'h3ee32e1e} /* (20, 24, 30) {real, imag} */,
  {32'hbf152b94, 32'hbe7efd92} /* (20, 24, 29) {real, imag} */,
  {32'h3d59e370, 32'hbe23b2f8} /* (20, 24, 28) {real, imag} */,
  {32'hbf2d4317, 32'h3f26517e} /* (20, 24, 27) {real, imag} */,
  {32'hbd5b9698, 32'hbe126f15} /* (20, 24, 26) {real, imag} */,
  {32'hbf0fd401, 32'hbe46e073} /* (20, 24, 25) {real, imag} */,
  {32'hbf274173, 32'h3c090f20} /* (20, 24, 24) {real, imag} */,
  {32'hbed65319, 32'hbe487fce} /* (20, 24, 23) {real, imag} */,
  {32'hbe99c774, 32'hbf602b54} /* (20, 24, 22) {real, imag} */,
  {32'h3e837d76, 32'h3d4ab458} /* (20, 24, 21) {real, imag} */,
  {32'hbdb085c3, 32'h3e9250c0} /* (20, 24, 20) {real, imag} */,
  {32'h3e0b5016, 32'hbe7f4639} /* (20, 24, 19) {real, imag} */,
  {32'h3b1b65c0, 32'hbdeaafba} /* (20, 24, 18) {real, imag} */,
  {32'hbe92b41e, 32'hbcb3b8e8} /* (20, 24, 17) {real, imag} */,
  {32'hbdca899b, 32'hbdd8e90e} /* (20, 24, 16) {real, imag} */,
  {32'hbd876cdd, 32'hbd3af460} /* (20, 24, 15) {real, imag} */,
  {32'hbdd10810, 32'hbbe5fe24} /* (20, 24, 14) {real, imag} */,
  {32'h3ef08ddc, 32'hbdc6578a} /* (20, 24, 13) {real, imag} */,
  {32'hbf366b68, 32'hbdf9e564} /* (20, 24, 12) {real, imag} */,
  {32'hbebc547c, 32'h3e81a1d0} /* (20, 24, 11) {real, imag} */,
  {32'hbd950460, 32'hbf3d0c72} /* (20, 24, 10) {real, imag} */,
  {32'hbc3f0c20, 32'h3ed7cc25} /* (20, 24, 9) {real, imag} */,
  {32'h3e68dfb5, 32'h3ee9b4fd} /* (20, 24, 8) {real, imag} */,
  {32'h3d9bd033, 32'h3e7893ec} /* (20, 24, 7) {real, imag} */,
  {32'h3e241e9d, 32'h3ec34443} /* (20, 24, 6) {real, imag} */,
  {32'hbf89ad76, 32'h3da8b10b} /* (20, 24, 5) {real, imag} */,
  {32'h3e3aa97f, 32'hbe551a45} /* (20, 24, 4) {real, imag} */,
  {32'h3ebdb43e, 32'h3eda03ea} /* (20, 24, 3) {real, imag} */,
  {32'hbe52b89c, 32'h3e470603} /* (20, 24, 2) {real, imag} */,
  {32'h3fd576b6, 32'hbfaa2995} /* (20, 24, 1) {real, imag} */,
  {32'h3f196922, 32'h3e893043} /* (20, 24, 0) {real, imag} */,
  {32'hbf1e807e, 32'h3f143045} /* (20, 23, 31) {real, imag} */,
  {32'hbf59495c, 32'hbe749d68} /* (20, 23, 30) {real, imag} */,
  {32'h3eac8f42, 32'h3ed1eab5} /* (20, 23, 29) {real, imag} */,
  {32'hbdd7d4b7, 32'hbdc998da} /* (20, 23, 28) {real, imag} */,
  {32'hbe19fd8a, 32'hbe05e56e} /* (20, 23, 27) {real, imag} */,
  {32'hbc0ec480, 32'hbea3e896} /* (20, 23, 26) {real, imag} */,
  {32'h3ddf0ea6, 32'h3dab067d} /* (20, 23, 25) {real, imag} */,
  {32'h3eada96f, 32'hbec4532d} /* (20, 23, 24) {real, imag} */,
  {32'h3e484159, 32'hbf3abc62} /* (20, 23, 23) {real, imag} */,
  {32'hbe2cc0fc, 32'h3e6f74b1} /* (20, 23, 22) {real, imag} */,
  {32'h3f00427d, 32'h3e1b8a6b} /* (20, 23, 21) {real, imag} */,
  {32'h3ed8f37f, 32'h3e427bc4} /* (20, 23, 20) {real, imag} */,
  {32'hbe922090, 32'h3e8dd33c} /* (20, 23, 19) {real, imag} */,
  {32'h3c9a3024, 32'h3f161592} /* (20, 23, 18) {real, imag} */,
  {32'h3d90260b, 32'hbdb25d72} /* (20, 23, 17) {real, imag} */,
  {32'hbed77ccb, 32'h3dd2d33d} /* (20, 23, 16) {real, imag} */,
  {32'hbc5e0b84, 32'h3e38d622} /* (20, 23, 15) {real, imag} */,
  {32'hbed4b4d6, 32'hbdddb367} /* (20, 23, 14) {real, imag} */,
  {32'hbe58d528, 32'hbe8f312d} /* (20, 23, 13) {real, imag} */,
  {32'h3ee0ada0, 32'h3eaec94c} /* (20, 23, 12) {real, imag} */,
  {32'hbe0f57c5, 32'h3da1eb32} /* (20, 23, 11) {real, imag} */,
  {32'hbee76224, 32'hbf2b7b67} /* (20, 23, 10) {real, imag} */,
  {32'hbda7bc41, 32'h3d995d68} /* (20, 23, 9) {real, imag} */,
  {32'h3dcb6008, 32'h3c178a40} /* (20, 23, 8) {real, imag} */,
  {32'h3eb878ec, 32'hbe42edf5} /* (20, 23, 7) {real, imag} */,
  {32'hbec3f1db, 32'hbf044168} /* (20, 23, 6) {real, imag} */,
  {32'hbe768727, 32'hbe6b5e42} /* (20, 23, 5) {real, imag} */,
  {32'hbef7257c, 32'h3dc1e740} /* (20, 23, 4) {real, imag} */,
  {32'h3e562968, 32'h3e6d1324} /* (20, 23, 3) {real, imag} */,
  {32'hbe7ed538, 32'h3d8b0454} /* (20, 23, 2) {real, imag} */,
  {32'h3ef2084f, 32'hbedd4f54} /* (20, 23, 1) {real, imag} */,
  {32'h3f0f1d57, 32'h3e5fec7e} /* (20, 23, 0) {real, imag} */,
  {32'hbdf79cbc, 32'hbe97fe50} /* (20, 22, 31) {real, imag} */,
  {32'h3ce14158, 32'hbe797ec8} /* (20, 22, 30) {real, imag} */,
  {32'h3f13f7bf, 32'hbf103d2e} /* (20, 22, 29) {real, imag} */,
  {32'hbd9c89e8, 32'h3f4eb1e9} /* (20, 22, 28) {real, imag} */,
  {32'hbeb42ffc, 32'h3e26b3cb} /* (20, 22, 27) {real, imag} */,
  {32'hbe5481f9, 32'hbc01b310} /* (20, 22, 26) {real, imag} */,
  {32'h3e1aa905, 32'hbc629f20} /* (20, 22, 25) {real, imag} */,
  {32'h3e3b37fe, 32'hbeb3f34c} /* (20, 22, 24) {real, imag} */,
  {32'hbf023fed, 32'hbcb1f9d8} /* (20, 22, 23) {real, imag} */,
  {32'h3e3d58e9, 32'hbd477aa8} /* (20, 22, 22) {real, imag} */,
  {32'h3f1d25e4, 32'hbe211c13} /* (20, 22, 21) {real, imag} */,
  {32'hbf4e18f8, 32'h3d48fda4} /* (20, 22, 20) {real, imag} */,
  {32'hbdbfa56e, 32'hbe9b6206} /* (20, 22, 19) {real, imag} */,
  {32'h3e197842, 32'hbed8fe88} /* (20, 22, 18) {real, imag} */,
  {32'hbc3d8420, 32'hbe0ad5d5} /* (20, 22, 17) {real, imag} */,
  {32'h3d5564f0, 32'hbe0ea540} /* (20, 22, 16) {real, imag} */,
  {32'hbcc09cee, 32'h3ea7f827} /* (20, 22, 15) {real, imag} */,
  {32'hbe5cab4e, 32'hbe6a10af} /* (20, 22, 14) {real, imag} */,
  {32'h3e164507, 32'hbe27cb7c} /* (20, 22, 13) {real, imag} */,
  {32'h3e106be9, 32'hbe29207a} /* (20, 22, 12) {real, imag} */,
  {32'hbcb61020, 32'hbf273318} /* (20, 22, 11) {real, imag} */,
  {32'h3e03457b, 32'h3e8925e2} /* (20, 22, 10) {real, imag} */,
  {32'hbe0fce1e, 32'hbf2cafbd} /* (20, 22, 9) {real, imag} */,
  {32'h3f323d2e, 32'h3e1741af} /* (20, 22, 8) {real, imag} */,
  {32'h3e191872, 32'h3dbe4b28} /* (20, 22, 7) {real, imag} */,
  {32'hbeeb6b10, 32'h3eab28e6} /* (20, 22, 6) {real, imag} */,
  {32'h3eb93084, 32'h3f1b80df} /* (20, 22, 5) {real, imag} */,
  {32'hbe9a9840, 32'h3f0a06da} /* (20, 22, 4) {real, imag} */,
  {32'hbf16c596, 32'h3c9de3f4} /* (20, 22, 3) {real, imag} */,
  {32'hbeac9115, 32'hbec46e40} /* (20, 22, 2) {real, imag} */,
  {32'h3dd5ffce, 32'h3c79ff20} /* (20, 22, 1) {real, imag} */,
  {32'h3e81d95e, 32'h3e773817} /* (20, 22, 0) {real, imag} */,
  {32'h3effc744, 32'hbef8a518} /* (20, 21, 31) {real, imag} */,
  {32'hbf037d69, 32'h3ee1abf5} /* (20, 21, 30) {real, imag} */,
  {32'hbd859f30, 32'h3ee73b40} /* (20, 21, 29) {real, imag} */,
  {32'hbec9f244, 32'h3d9f8b90} /* (20, 21, 28) {real, imag} */,
  {32'hbea904f1, 32'h3d7ffeb4} /* (20, 21, 27) {real, imag} */,
  {32'h3e1c2eb3, 32'h3e56ea06} /* (20, 21, 26) {real, imag} */,
  {32'h3e020afa, 32'hbf250bb4} /* (20, 21, 25) {real, imag} */,
  {32'hbef49eee, 32'h3e3329c9} /* (20, 21, 24) {real, imag} */,
  {32'hbefa0ea9, 32'h3f1616c6} /* (20, 21, 23) {real, imag} */,
  {32'hbe6ebb33, 32'h3dd41ac4} /* (20, 21, 22) {real, imag} */,
  {32'h3e3694b9, 32'h3e2f870a} /* (20, 21, 21) {real, imag} */,
  {32'hbde44378, 32'h3cfe0750} /* (20, 21, 20) {real, imag} */,
  {32'hbb66ddb0, 32'hbdb73a3c} /* (20, 21, 19) {real, imag} */,
  {32'hbe7d1eaa, 32'h3e919cea} /* (20, 21, 18) {real, imag} */,
  {32'h3e999130, 32'hbd1e4172} /* (20, 21, 17) {real, imag} */,
  {32'hbdf20fc0, 32'hbd1c089a} /* (20, 21, 16) {real, imag} */,
  {32'hbe878307, 32'hbf21241f} /* (20, 21, 15) {real, imag} */,
  {32'h3ecdb8c8, 32'h3c8ee064} /* (20, 21, 14) {real, imag} */,
  {32'hbba56840, 32'h3e6731a8} /* (20, 21, 13) {real, imag} */,
  {32'hbe133330, 32'h3de8cdfa} /* (20, 21, 12) {real, imag} */,
  {32'h3d82f1c0, 32'h3ebf757c} /* (20, 21, 11) {real, imag} */,
  {32'hbe0e4b82, 32'h3e8d0ce1} /* (20, 21, 10) {real, imag} */,
  {32'h3eea664f, 32'h3eddc5cf} /* (20, 21, 9) {real, imag} */,
  {32'hbea17a93, 32'h3dbcc7a1} /* (20, 21, 8) {real, imag} */,
  {32'hbf32b481, 32'h3db5a5c0} /* (20, 21, 7) {real, imag} */,
  {32'hbf034b62, 32'h3ee25048} /* (20, 21, 6) {real, imag} */,
  {32'hbcb7e13c, 32'hbd9d215a} /* (20, 21, 5) {real, imag} */,
  {32'hbe56eb4a, 32'h3f16368c} /* (20, 21, 4) {real, imag} */,
  {32'hbe73ffdc, 32'hbd143577} /* (20, 21, 3) {real, imag} */,
  {32'hbcef5630, 32'hbc66d300} /* (20, 21, 2) {real, imag} */,
  {32'h3f0e061a, 32'hbf263a66} /* (20, 21, 1) {real, imag} */,
  {32'h3ee73e20, 32'hbec16aeb} /* (20, 21, 0) {real, imag} */,
  {32'hbde0d1f5, 32'hbe6199c4} /* (20, 20, 31) {real, imag} */,
  {32'h3cebbc38, 32'hbf180fda} /* (20, 20, 30) {real, imag} */,
  {32'hbedaed6e, 32'h3efbcee9} /* (20, 20, 29) {real, imag} */,
  {32'h3d676ecb, 32'h3e855e21} /* (20, 20, 28) {real, imag} */,
  {32'hbe52581a, 32'h3e10eca0} /* (20, 20, 27) {real, imag} */,
  {32'hbea425aa, 32'hbe122e48} /* (20, 20, 26) {real, imag} */,
  {32'h3f4c3823, 32'h3e540565} /* (20, 20, 25) {real, imag} */,
  {32'h3e92ea43, 32'hbf2d8baf} /* (20, 20, 24) {real, imag} */,
  {32'hbe5d6814, 32'hbe98d146} /* (20, 20, 23) {real, imag} */,
  {32'hbd59c428, 32'h3ed03b95} /* (20, 20, 22) {real, imag} */,
  {32'hbe0fc422, 32'hbbd5ab40} /* (20, 20, 21) {real, imag} */,
  {32'hbe270450, 32'hbf06fa40} /* (20, 20, 20) {real, imag} */,
  {32'h3e5f5084, 32'hbe08f9f3} /* (20, 20, 19) {real, imag} */,
  {32'h3dd36183, 32'hbd725a7c} /* (20, 20, 18) {real, imag} */,
  {32'h3e2996a4, 32'h3da71970} /* (20, 20, 17) {real, imag} */,
  {32'hbdd892e6, 32'h3ea7d392} /* (20, 20, 16) {real, imag} */,
  {32'h3eb64af0, 32'hbde03a0f} /* (20, 20, 15) {real, imag} */,
  {32'hbc9232d8, 32'h3dc15230} /* (20, 20, 14) {real, imag} */,
  {32'hbce0cc28, 32'hbead475f} /* (20, 20, 13) {real, imag} */,
  {32'h3ec4a79c, 32'hbe783d26} /* (20, 20, 12) {real, imag} */,
  {32'hbe8dfcec, 32'h3dd0d9d5} /* (20, 20, 11) {real, imag} */,
  {32'hbeaec521, 32'h3eef0b4c} /* (20, 20, 10) {real, imag} */,
  {32'h3ea87d1e, 32'hbedc99c8} /* (20, 20, 9) {real, imag} */,
  {32'h3eb1b9d6, 32'hbd8d8ce5} /* (20, 20, 8) {real, imag} */,
  {32'h3e7f4545, 32'hbf31ac6d} /* (20, 20, 7) {real, imag} */,
  {32'h3e2d4968, 32'hbe9869a1} /* (20, 20, 6) {real, imag} */,
  {32'hbe5778ca, 32'hbc99d0d8} /* (20, 20, 5) {real, imag} */,
  {32'h3f067514, 32'h3db071f9} /* (20, 20, 4) {real, imag} */,
  {32'h3dfb1c18, 32'hbe1d0008} /* (20, 20, 3) {real, imag} */,
  {32'hbf195553, 32'h3e5e776a} /* (20, 20, 2) {real, imag} */,
  {32'hbe913700, 32'hbd7e883c} /* (20, 20, 1) {real, imag} */,
  {32'hbd7fd774, 32'h3df03531} /* (20, 20, 0) {real, imag} */,
  {32'hbe84051e, 32'h3c9d0394} /* (20, 19, 31) {real, imag} */,
  {32'h3e918f1f, 32'h3e92943a} /* (20, 19, 30) {real, imag} */,
  {32'h3d2ae097, 32'hbe9fc451} /* (20, 19, 29) {real, imag} */,
  {32'h3e0a9e38, 32'h3d80fa7c} /* (20, 19, 28) {real, imag} */,
  {32'hbe69cc58, 32'hbed60b12} /* (20, 19, 27) {real, imag} */,
  {32'h3ecf681e, 32'hbd77ceca} /* (20, 19, 26) {real, imag} */,
  {32'hbeb905bb, 32'hbea872f5} /* (20, 19, 25) {real, imag} */,
  {32'h3ea8bb3c, 32'hbe808b09} /* (20, 19, 24) {real, imag} */,
  {32'h3e573663, 32'hbe26e9d2} /* (20, 19, 23) {real, imag} */,
  {32'h3e47dbd1, 32'h3e7312c6} /* (20, 19, 22) {real, imag} */,
  {32'hbf2dbe52, 32'h3ed3e8b4} /* (20, 19, 21) {real, imag} */,
  {32'hbe672b62, 32'h3ea5ff9d} /* (20, 19, 20) {real, imag} */,
  {32'hbe26722d, 32'h3c7c5280} /* (20, 19, 19) {real, imag} */,
  {32'h3e7c8e6e, 32'h3e8cdacb} /* (20, 19, 18) {real, imag} */,
  {32'hbecf404a, 32'h3e8cef46} /* (20, 19, 17) {real, imag} */,
  {32'h3ea802fa, 32'h3e7b73f8} /* (20, 19, 16) {real, imag} */,
  {32'h3e552468, 32'hbd6fcfa9} /* (20, 19, 15) {real, imag} */,
  {32'hbe6d47b8, 32'h3edff0ac} /* (20, 19, 14) {real, imag} */,
  {32'h3e16fd16, 32'h3df2d863} /* (20, 19, 13) {real, imag} */,
  {32'hbf24757d, 32'h3f513359} /* (20, 19, 12) {real, imag} */,
  {32'h3e061072, 32'h3eb68904} /* (20, 19, 11) {real, imag} */,
  {32'hbeb5112e, 32'hbde92d3c} /* (20, 19, 10) {real, imag} */,
  {32'h3e82b7da, 32'hbe30d6cd} /* (20, 19, 9) {real, imag} */,
  {32'hbe5b4e72, 32'hbed77998} /* (20, 19, 8) {real, imag} */,
  {32'h3dbfc495, 32'h3ec0f357} /* (20, 19, 7) {real, imag} */,
  {32'hbe201a77, 32'hbcaf6ca2} /* (20, 19, 6) {real, imag} */,
  {32'h3e21eec7, 32'h3e828af7} /* (20, 19, 5) {real, imag} */,
  {32'hbe9d89e4, 32'h3e8052a6} /* (20, 19, 4) {real, imag} */,
  {32'h3e6a6a76, 32'hbe029b20} /* (20, 19, 3) {real, imag} */,
  {32'hbe0ce87f, 32'hbe30bfaf} /* (20, 19, 2) {real, imag} */,
  {32'h3c32c170, 32'h3e5f20b9} /* (20, 19, 1) {real, imag} */,
  {32'hbe95487a, 32'h3e7aca54} /* (20, 19, 0) {real, imag} */,
  {32'hbeef8674, 32'hbe958c69} /* (20, 18, 31) {real, imag} */,
  {32'hbb972930, 32'h3e311de0} /* (20, 18, 30) {real, imag} */,
  {32'h3e6c414d, 32'h3c597940} /* (20, 18, 29) {real, imag} */,
  {32'hbd1aabc0, 32'h3ef4bf74} /* (20, 18, 28) {real, imag} */,
  {32'h3e851322, 32'hbe2de898} /* (20, 18, 27) {real, imag} */,
  {32'hbe8f1d4c, 32'h3e549906} /* (20, 18, 26) {real, imag} */,
  {32'h3e81c1c3, 32'hbe91b35f} /* (20, 18, 25) {real, imag} */,
  {32'h3ea5e9f1, 32'h3d2291c5} /* (20, 18, 24) {real, imag} */,
  {32'h3d7e3a64, 32'h3ec28b8c} /* (20, 18, 23) {real, imag} */,
  {32'h3f04259a, 32'hbe0f0c70} /* (20, 18, 22) {real, imag} */,
  {32'hbd998e22, 32'hbe51ac39} /* (20, 18, 21) {real, imag} */,
  {32'h3da4dfde, 32'hbebf9972} /* (20, 18, 20) {real, imag} */,
  {32'h3dcdc0ac, 32'hbdb08fe2} /* (20, 18, 19) {real, imag} */,
  {32'h3cb5f0ac, 32'h3e1cfb83} /* (20, 18, 18) {real, imag} */,
  {32'hbc856176, 32'hbe78f2c6} /* (20, 18, 17) {real, imag} */,
  {32'h3e1fd6d5, 32'hbe4e4c56} /* (20, 18, 16) {real, imag} */,
  {32'h3ea8fe52, 32'h3e296904} /* (20, 18, 15) {real, imag} */,
  {32'h3dbea7e0, 32'h3e93e2b4} /* (20, 18, 14) {real, imag} */,
  {32'hbf103e28, 32'hbee2024c} /* (20, 18, 13) {real, imag} */,
  {32'h3ee82fd3, 32'hbedc606e} /* (20, 18, 12) {real, imag} */,
  {32'h3e07be00, 32'h3dcbaf9a} /* (20, 18, 11) {real, imag} */,
  {32'hbea2efe9, 32'h3df16341} /* (20, 18, 10) {real, imag} */,
  {32'h3e94f344, 32'hbe4206e0} /* (20, 18, 9) {real, imag} */,
  {32'hbe8e90de, 32'h3eebb45c} /* (20, 18, 8) {real, imag} */,
  {32'h3e5c5094, 32'hbbd24020} /* (20, 18, 7) {real, imag} */,
  {32'hbc7f05d0, 32'h3d9374db} /* (20, 18, 6) {real, imag} */,
  {32'h3ae23f00, 32'h3d9beff0} /* (20, 18, 5) {real, imag} */,
  {32'h3ecd78d5, 32'h3e1544ec} /* (20, 18, 4) {real, imag} */,
  {32'hbb91d4b4, 32'hbd19f54b} /* (20, 18, 3) {real, imag} */,
  {32'hbeaca460, 32'h3d2717a0} /* (20, 18, 2) {real, imag} */,
  {32'hbd230144, 32'hbedafaef} /* (20, 18, 1) {real, imag} */,
  {32'hbb4ec550, 32'hbef09d26} /* (20, 18, 0) {real, imag} */,
  {32'h3e640a98, 32'h3d97ff4a} /* (20, 17, 31) {real, imag} */,
  {32'h3ece845e, 32'h3c3e7f38} /* (20, 17, 30) {real, imag} */,
  {32'h3d8ee998, 32'h3e667586} /* (20, 17, 29) {real, imag} */,
  {32'h3d48fd87, 32'hbe2a93e6} /* (20, 17, 28) {real, imag} */,
  {32'hbd56296e, 32'hbc494e88} /* (20, 17, 27) {real, imag} */,
  {32'hbebe5cea, 32'h3e8ea8aa} /* (20, 17, 26) {real, imag} */,
  {32'hbe3386e2, 32'hbc2441e0} /* (20, 17, 25) {real, imag} */,
  {32'h3ce8d978, 32'hbe996046} /* (20, 17, 24) {real, imag} */,
  {32'hbde4446e, 32'h3cf8ea00} /* (20, 17, 23) {real, imag} */,
  {32'h3e62f4ee, 32'h3c8e7364} /* (20, 17, 22) {real, imag} */,
  {32'h3e096802, 32'hbdb5da11} /* (20, 17, 21) {real, imag} */,
  {32'hbe8846b9, 32'hbeb5d999} /* (20, 17, 20) {real, imag} */,
  {32'hbcc1552c, 32'hbe26d6a1} /* (20, 17, 19) {real, imag} */,
  {32'hbcd36e50, 32'h3d830168} /* (20, 17, 18) {real, imag} */,
  {32'hbe6c6d02, 32'h3e8511a4} /* (20, 17, 17) {real, imag} */,
  {32'hbd8078b1, 32'h3e84c500} /* (20, 17, 16) {real, imag} */,
  {32'hbec7b25d, 32'hbe0b29c1} /* (20, 17, 15) {real, imag} */,
  {32'hbed1ea94, 32'h3e2e1372} /* (20, 17, 14) {real, imag} */,
  {32'hbeaf8a34, 32'h3e9253df} /* (20, 17, 13) {real, imag} */,
  {32'hbe14c5a0, 32'hbcb8d480} /* (20, 17, 12) {real, imag} */,
  {32'h3e9860da, 32'h3ea4e572} /* (20, 17, 11) {real, imag} */,
  {32'hbeffea06, 32'hbe9f9b9f} /* (20, 17, 10) {real, imag} */,
  {32'hbe84903e, 32'hbec417f3} /* (20, 17, 9) {real, imag} */,
  {32'hbea4cfd0, 32'hbed3f637} /* (20, 17, 8) {real, imag} */,
  {32'h3c5d0950, 32'h3e266c38} /* (20, 17, 7) {real, imag} */,
  {32'hbe2bfff4, 32'h3eb1c06c} /* (20, 17, 6) {real, imag} */,
  {32'hbdb890be, 32'hbd5a4717} /* (20, 17, 5) {real, imag} */,
  {32'hbe90d1b0, 32'hbeb2e37f} /* (20, 17, 4) {real, imag} */,
  {32'hbf101476, 32'hbeac9f35} /* (20, 17, 3) {real, imag} */,
  {32'h3e07cca0, 32'hbd699f40} /* (20, 17, 2) {real, imag} */,
  {32'hbde53982, 32'h3e5fd27f} /* (20, 17, 1) {real, imag} */,
  {32'h3d5790b8, 32'h3e88c6cd} /* (20, 17, 0) {real, imag} */,
  {32'hbec93c4d, 32'h3ca7cfda} /* (20, 16, 31) {real, imag} */,
  {32'h3e803c0a, 32'hbbbdc870} /* (20, 16, 30) {real, imag} */,
  {32'h3b6731a0, 32'hbe41c9cf} /* (20, 16, 29) {real, imag} */,
  {32'hbda40029, 32'hbd8fde18} /* (20, 16, 28) {real, imag} */,
  {32'h3d91d80a, 32'hbdd7d4aa} /* (20, 16, 27) {real, imag} */,
  {32'h3e821b04, 32'hbeb2cd78} /* (20, 16, 26) {real, imag} */,
  {32'hbe8cb490, 32'h3e258422} /* (20, 16, 25) {real, imag} */,
  {32'hbd2a080c, 32'h39e9ab00} /* (20, 16, 24) {real, imag} */,
  {32'h3c6c1548, 32'h3dfcfe5e} /* (20, 16, 23) {real, imag} */,
  {32'hbe97ab87, 32'h3e0fb979} /* (20, 16, 22) {real, imag} */,
  {32'hbe0afeea, 32'h3e810373} /* (20, 16, 21) {real, imag} */,
  {32'h3d10979f, 32'hbf153760} /* (20, 16, 20) {real, imag} */,
  {32'h3e9b3d96, 32'h3e43294e} /* (20, 16, 19) {real, imag} */,
  {32'hbe0ddc74, 32'h3e88f533} /* (20, 16, 18) {real, imag} */,
  {32'h3d7ff234, 32'hbd701c47} /* (20, 16, 17) {real, imag} */,
  {32'hbdf66ca0, 32'h00000000} /* (20, 16, 16) {real, imag} */,
  {32'h3d7ff234, 32'h3d701c47} /* (20, 16, 15) {real, imag} */,
  {32'hbe0ddc74, 32'hbe88f533} /* (20, 16, 14) {real, imag} */,
  {32'h3e9b3d96, 32'hbe43294e} /* (20, 16, 13) {real, imag} */,
  {32'h3d10979f, 32'h3f153760} /* (20, 16, 12) {real, imag} */,
  {32'hbe0afeea, 32'hbe810373} /* (20, 16, 11) {real, imag} */,
  {32'hbe97ab87, 32'hbe0fb979} /* (20, 16, 10) {real, imag} */,
  {32'h3c6c1548, 32'hbdfcfe5e} /* (20, 16, 9) {real, imag} */,
  {32'hbd2a080c, 32'hb9e9ab00} /* (20, 16, 8) {real, imag} */,
  {32'hbe8cb490, 32'hbe258422} /* (20, 16, 7) {real, imag} */,
  {32'h3e821b04, 32'h3eb2cd78} /* (20, 16, 6) {real, imag} */,
  {32'h3d91d80a, 32'h3dd7d4aa} /* (20, 16, 5) {real, imag} */,
  {32'hbda40029, 32'h3d8fde18} /* (20, 16, 4) {real, imag} */,
  {32'h3b6731a0, 32'h3e41c9cf} /* (20, 16, 3) {real, imag} */,
  {32'h3e803c0a, 32'h3bbdc870} /* (20, 16, 2) {real, imag} */,
  {32'hbec93c4d, 32'hbca7cfda} /* (20, 16, 1) {real, imag} */,
  {32'h3d5ad272, 32'h00000000} /* (20, 16, 0) {real, imag} */,
  {32'hbde53982, 32'hbe5fd27f} /* (20, 15, 31) {real, imag} */,
  {32'h3e07cca0, 32'h3d699f40} /* (20, 15, 30) {real, imag} */,
  {32'hbf101476, 32'h3eac9f35} /* (20, 15, 29) {real, imag} */,
  {32'hbe90d1b0, 32'h3eb2e37f} /* (20, 15, 28) {real, imag} */,
  {32'hbdb890be, 32'h3d5a4717} /* (20, 15, 27) {real, imag} */,
  {32'hbe2bfff4, 32'hbeb1c06c} /* (20, 15, 26) {real, imag} */,
  {32'h3c5d0950, 32'hbe266c38} /* (20, 15, 25) {real, imag} */,
  {32'hbea4cfd0, 32'h3ed3f637} /* (20, 15, 24) {real, imag} */,
  {32'hbe84903e, 32'h3ec417f3} /* (20, 15, 23) {real, imag} */,
  {32'hbeffea06, 32'h3e9f9b9f} /* (20, 15, 22) {real, imag} */,
  {32'h3e9860da, 32'hbea4e572} /* (20, 15, 21) {real, imag} */,
  {32'hbe14c5a0, 32'h3cb8d480} /* (20, 15, 20) {real, imag} */,
  {32'hbeaf8a34, 32'hbe9253df} /* (20, 15, 19) {real, imag} */,
  {32'hbed1ea94, 32'hbe2e1372} /* (20, 15, 18) {real, imag} */,
  {32'hbec7b25d, 32'h3e0b29c1} /* (20, 15, 17) {real, imag} */,
  {32'hbd8078b1, 32'hbe84c500} /* (20, 15, 16) {real, imag} */,
  {32'hbe6c6d02, 32'hbe8511a4} /* (20, 15, 15) {real, imag} */,
  {32'hbcd36e50, 32'hbd830168} /* (20, 15, 14) {real, imag} */,
  {32'hbcc1552c, 32'h3e26d6a1} /* (20, 15, 13) {real, imag} */,
  {32'hbe8846b9, 32'h3eb5d999} /* (20, 15, 12) {real, imag} */,
  {32'h3e096802, 32'h3db5da11} /* (20, 15, 11) {real, imag} */,
  {32'h3e62f4ee, 32'hbc8e7364} /* (20, 15, 10) {real, imag} */,
  {32'hbde4446e, 32'hbcf8ea00} /* (20, 15, 9) {real, imag} */,
  {32'h3ce8d978, 32'h3e996046} /* (20, 15, 8) {real, imag} */,
  {32'hbe3386e2, 32'h3c2441e0} /* (20, 15, 7) {real, imag} */,
  {32'hbebe5cea, 32'hbe8ea8aa} /* (20, 15, 6) {real, imag} */,
  {32'hbd56296e, 32'h3c494e88} /* (20, 15, 5) {real, imag} */,
  {32'h3d48fd87, 32'h3e2a93e6} /* (20, 15, 4) {real, imag} */,
  {32'h3d8ee998, 32'hbe667586} /* (20, 15, 3) {real, imag} */,
  {32'h3ece845e, 32'hbc3e7f38} /* (20, 15, 2) {real, imag} */,
  {32'h3e640a98, 32'hbd97ff4a} /* (20, 15, 1) {real, imag} */,
  {32'h3d5790b8, 32'hbe88c6cd} /* (20, 15, 0) {real, imag} */,
  {32'hbd230144, 32'h3edafaef} /* (20, 14, 31) {real, imag} */,
  {32'hbeaca460, 32'hbd2717a0} /* (20, 14, 30) {real, imag} */,
  {32'hbb91d4b4, 32'h3d19f54b} /* (20, 14, 29) {real, imag} */,
  {32'h3ecd78d5, 32'hbe1544ec} /* (20, 14, 28) {real, imag} */,
  {32'h3ae23f00, 32'hbd9beff0} /* (20, 14, 27) {real, imag} */,
  {32'hbc7f05d0, 32'hbd9374db} /* (20, 14, 26) {real, imag} */,
  {32'h3e5c5094, 32'h3bd24020} /* (20, 14, 25) {real, imag} */,
  {32'hbe8e90de, 32'hbeebb45c} /* (20, 14, 24) {real, imag} */,
  {32'h3e94f344, 32'h3e4206e0} /* (20, 14, 23) {real, imag} */,
  {32'hbea2efe9, 32'hbdf16341} /* (20, 14, 22) {real, imag} */,
  {32'h3e07be00, 32'hbdcbaf9a} /* (20, 14, 21) {real, imag} */,
  {32'h3ee82fd3, 32'h3edc606e} /* (20, 14, 20) {real, imag} */,
  {32'hbf103e28, 32'h3ee2024c} /* (20, 14, 19) {real, imag} */,
  {32'h3dbea7e0, 32'hbe93e2b4} /* (20, 14, 18) {real, imag} */,
  {32'h3ea8fe52, 32'hbe296904} /* (20, 14, 17) {real, imag} */,
  {32'h3e1fd6d5, 32'h3e4e4c56} /* (20, 14, 16) {real, imag} */,
  {32'hbc856176, 32'h3e78f2c6} /* (20, 14, 15) {real, imag} */,
  {32'h3cb5f0ac, 32'hbe1cfb83} /* (20, 14, 14) {real, imag} */,
  {32'h3dcdc0ac, 32'h3db08fe2} /* (20, 14, 13) {real, imag} */,
  {32'h3da4dfde, 32'h3ebf9972} /* (20, 14, 12) {real, imag} */,
  {32'hbd998e22, 32'h3e51ac39} /* (20, 14, 11) {real, imag} */,
  {32'h3f04259a, 32'h3e0f0c70} /* (20, 14, 10) {real, imag} */,
  {32'h3d7e3a64, 32'hbec28b8c} /* (20, 14, 9) {real, imag} */,
  {32'h3ea5e9f1, 32'hbd2291c5} /* (20, 14, 8) {real, imag} */,
  {32'h3e81c1c3, 32'h3e91b35f} /* (20, 14, 7) {real, imag} */,
  {32'hbe8f1d4c, 32'hbe549906} /* (20, 14, 6) {real, imag} */,
  {32'h3e851322, 32'h3e2de898} /* (20, 14, 5) {real, imag} */,
  {32'hbd1aabc0, 32'hbef4bf74} /* (20, 14, 4) {real, imag} */,
  {32'h3e6c414d, 32'hbc597940} /* (20, 14, 3) {real, imag} */,
  {32'hbb972930, 32'hbe311de0} /* (20, 14, 2) {real, imag} */,
  {32'hbeef8674, 32'h3e958c69} /* (20, 14, 1) {real, imag} */,
  {32'hbb4ec550, 32'h3ef09d26} /* (20, 14, 0) {real, imag} */,
  {32'h3c32c170, 32'hbe5f20b9} /* (20, 13, 31) {real, imag} */,
  {32'hbe0ce87f, 32'h3e30bfaf} /* (20, 13, 30) {real, imag} */,
  {32'h3e6a6a76, 32'h3e029b20} /* (20, 13, 29) {real, imag} */,
  {32'hbe9d89e4, 32'hbe8052a6} /* (20, 13, 28) {real, imag} */,
  {32'h3e21eec7, 32'hbe828af7} /* (20, 13, 27) {real, imag} */,
  {32'hbe201a77, 32'h3caf6ca2} /* (20, 13, 26) {real, imag} */,
  {32'h3dbfc495, 32'hbec0f357} /* (20, 13, 25) {real, imag} */,
  {32'hbe5b4e72, 32'h3ed77998} /* (20, 13, 24) {real, imag} */,
  {32'h3e82b7da, 32'h3e30d6cd} /* (20, 13, 23) {real, imag} */,
  {32'hbeb5112e, 32'h3de92d3c} /* (20, 13, 22) {real, imag} */,
  {32'h3e061072, 32'hbeb68904} /* (20, 13, 21) {real, imag} */,
  {32'hbf24757d, 32'hbf513359} /* (20, 13, 20) {real, imag} */,
  {32'h3e16fd16, 32'hbdf2d863} /* (20, 13, 19) {real, imag} */,
  {32'hbe6d47b8, 32'hbedff0ac} /* (20, 13, 18) {real, imag} */,
  {32'h3e552468, 32'h3d6fcfa9} /* (20, 13, 17) {real, imag} */,
  {32'h3ea802fa, 32'hbe7b73f8} /* (20, 13, 16) {real, imag} */,
  {32'hbecf404a, 32'hbe8cef46} /* (20, 13, 15) {real, imag} */,
  {32'h3e7c8e6e, 32'hbe8cdacb} /* (20, 13, 14) {real, imag} */,
  {32'hbe26722d, 32'hbc7c5280} /* (20, 13, 13) {real, imag} */,
  {32'hbe672b62, 32'hbea5ff9d} /* (20, 13, 12) {real, imag} */,
  {32'hbf2dbe52, 32'hbed3e8b4} /* (20, 13, 11) {real, imag} */,
  {32'h3e47dbd1, 32'hbe7312c6} /* (20, 13, 10) {real, imag} */,
  {32'h3e573663, 32'h3e26e9d2} /* (20, 13, 9) {real, imag} */,
  {32'h3ea8bb3c, 32'h3e808b09} /* (20, 13, 8) {real, imag} */,
  {32'hbeb905bb, 32'h3ea872f5} /* (20, 13, 7) {real, imag} */,
  {32'h3ecf681e, 32'h3d77ceca} /* (20, 13, 6) {real, imag} */,
  {32'hbe69cc58, 32'h3ed60b12} /* (20, 13, 5) {real, imag} */,
  {32'h3e0a9e38, 32'hbd80fa7c} /* (20, 13, 4) {real, imag} */,
  {32'h3d2ae097, 32'h3e9fc451} /* (20, 13, 3) {real, imag} */,
  {32'h3e918f1f, 32'hbe92943a} /* (20, 13, 2) {real, imag} */,
  {32'hbe84051e, 32'hbc9d0394} /* (20, 13, 1) {real, imag} */,
  {32'hbe95487a, 32'hbe7aca54} /* (20, 13, 0) {real, imag} */,
  {32'hbe913700, 32'h3d7e883c} /* (20, 12, 31) {real, imag} */,
  {32'hbf195553, 32'hbe5e776a} /* (20, 12, 30) {real, imag} */,
  {32'h3dfb1c18, 32'h3e1d0008} /* (20, 12, 29) {real, imag} */,
  {32'h3f067514, 32'hbdb071f9} /* (20, 12, 28) {real, imag} */,
  {32'hbe5778ca, 32'h3c99d0d8} /* (20, 12, 27) {real, imag} */,
  {32'h3e2d4968, 32'h3e9869a1} /* (20, 12, 26) {real, imag} */,
  {32'h3e7f4545, 32'h3f31ac6d} /* (20, 12, 25) {real, imag} */,
  {32'h3eb1b9d6, 32'h3d8d8ce5} /* (20, 12, 24) {real, imag} */,
  {32'h3ea87d1e, 32'h3edc99c8} /* (20, 12, 23) {real, imag} */,
  {32'hbeaec521, 32'hbeef0b4c} /* (20, 12, 22) {real, imag} */,
  {32'hbe8dfcec, 32'hbdd0d9d5} /* (20, 12, 21) {real, imag} */,
  {32'h3ec4a79c, 32'h3e783d26} /* (20, 12, 20) {real, imag} */,
  {32'hbce0cc28, 32'h3ead475f} /* (20, 12, 19) {real, imag} */,
  {32'hbc9232d8, 32'hbdc15230} /* (20, 12, 18) {real, imag} */,
  {32'h3eb64af0, 32'h3de03a0f} /* (20, 12, 17) {real, imag} */,
  {32'hbdd892e6, 32'hbea7d392} /* (20, 12, 16) {real, imag} */,
  {32'h3e2996a4, 32'hbda71970} /* (20, 12, 15) {real, imag} */,
  {32'h3dd36183, 32'h3d725a7c} /* (20, 12, 14) {real, imag} */,
  {32'h3e5f5084, 32'h3e08f9f3} /* (20, 12, 13) {real, imag} */,
  {32'hbe270450, 32'h3f06fa40} /* (20, 12, 12) {real, imag} */,
  {32'hbe0fc422, 32'h3bd5ab40} /* (20, 12, 11) {real, imag} */,
  {32'hbd59c428, 32'hbed03b95} /* (20, 12, 10) {real, imag} */,
  {32'hbe5d6814, 32'h3e98d146} /* (20, 12, 9) {real, imag} */,
  {32'h3e92ea43, 32'h3f2d8baf} /* (20, 12, 8) {real, imag} */,
  {32'h3f4c3823, 32'hbe540565} /* (20, 12, 7) {real, imag} */,
  {32'hbea425aa, 32'h3e122e48} /* (20, 12, 6) {real, imag} */,
  {32'hbe52581a, 32'hbe10eca0} /* (20, 12, 5) {real, imag} */,
  {32'h3d676ecb, 32'hbe855e21} /* (20, 12, 4) {real, imag} */,
  {32'hbedaed6e, 32'hbefbcee9} /* (20, 12, 3) {real, imag} */,
  {32'h3cebbc38, 32'h3f180fda} /* (20, 12, 2) {real, imag} */,
  {32'hbde0d1f5, 32'h3e6199c4} /* (20, 12, 1) {real, imag} */,
  {32'hbd7fd774, 32'hbdf03531} /* (20, 12, 0) {real, imag} */,
  {32'h3f0e061a, 32'h3f263a66} /* (20, 11, 31) {real, imag} */,
  {32'hbcef5630, 32'h3c66d300} /* (20, 11, 30) {real, imag} */,
  {32'hbe73ffdc, 32'h3d143577} /* (20, 11, 29) {real, imag} */,
  {32'hbe56eb4a, 32'hbf16368c} /* (20, 11, 28) {real, imag} */,
  {32'hbcb7e13c, 32'h3d9d215a} /* (20, 11, 27) {real, imag} */,
  {32'hbf034b62, 32'hbee25048} /* (20, 11, 26) {real, imag} */,
  {32'hbf32b481, 32'hbdb5a5c0} /* (20, 11, 25) {real, imag} */,
  {32'hbea17a93, 32'hbdbcc7a1} /* (20, 11, 24) {real, imag} */,
  {32'h3eea664f, 32'hbeddc5cf} /* (20, 11, 23) {real, imag} */,
  {32'hbe0e4b82, 32'hbe8d0ce1} /* (20, 11, 22) {real, imag} */,
  {32'h3d82f1c0, 32'hbebf757c} /* (20, 11, 21) {real, imag} */,
  {32'hbe133330, 32'hbde8cdfa} /* (20, 11, 20) {real, imag} */,
  {32'hbba56840, 32'hbe6731a8} /* (20, 11, 19) {real, imag} */,
  {32'h3ecdb8c8, 32'hbc8ee064} /* (20, 11, 18) {real, imag} */,
  {32'hbe878307, 32'h3f21241f} /* (20, 11, 17) {real, imag} */,
  {32'hbdf20fc0, 32'h3d1c089a} /* (20, 11, 16) {real, imag} */,
  {32'h3e999130, 32'h3d1e4172} /* (20, 11, 15) {real, imag} */,
  {32'hbe7d1eaa, 32'hbe919cea} /* (20, 11, 14) {real, imag} */,
  {32'hbb66ddb0, 32'h3db73a3c} /* (20, 11, 13) {real, imag} */,
  {32'hbde44378, 32'hbcfe0750} /* (20, 11, 12) {real, imag} */,
  {32'h3e3694b9, 32'hbe2f870a} /* (20, 11, 11) {real, imag} */,
  {32'hbe6ebb33, 32'hbdd41ac4} /* (20, 11, 10) {real, imag} */,
  {32'hbefa0ea9, 32'hbf1616c6} /* (20, 11, 9) {real, imag} */,
  {32'hbef49eee, 32'hbe3329c9} /* (20, 11, 8) {real, imag} */,
  {32'h3e020afa, 32'h3f250bb4} /* (20, 11, 7) {real, imag} */,
  {32'h3e1c2eb3, 32'hbe56ea06} /* (20, 11, 6) {real, imag} */,
  {32'hbea904f1, 32'hbd7ffeb4} /* (20, 11, 5) {real, imag} */,
  {32'hbec9f244, 32'hbd9f8b90} /* (20, 11, 4) {real, imag} */,
  {32'hbd859f30, 32'hbee73b40} /* (20, 11, 3) {real, imag} */,
  {32'hbf037d69, 32'hbee1abf5} /* (20, 11, 2) {real, imag} */,
  {32'h3effc744, 32'h3ef8a518} /* (20, 11, 1) {real, imag} */,
  {32'h3ee73e20, 32'h3ec16aeb} /* (20, 11, 0) {real, imag} */,
  {32'h3dd5ffce, 32'hbc79ff20} /* (20, 10, 31) {real, imag} */,
  {32'hbeac9115, 32'h3ec46e40} /* (20, 10, 30) {real, imag} */,
  {32'hbf16c596, 32'hbc9de3f4} /* (20, 10, 29) {real, imag} */,
  {32'hbe9a9840, 32'hbf0a06da} /* (20, 10, 28) {real, imag} */,
  {32'h3eb93084, 32'hbf1b80df} /* (20, 10, 27) {real, imag} */,
  {32'hbeeb6b10, 32'hbeab28e6} /* (20, 10, 26) {real, imag} */,
  {32'h3e191872, 32'hbdbe4b28} /* (20, 10, 25) {real, imag} */,
  {32'h3f323d2e, 32'hbe1741af} /* (20, 10, 24) {real, imag} */,
  {32'hbe0fce1e, 32'h3f2cafbd} /* (20, 10, 23) {real, imag} */,
  {32'h3e03457b, 32'hbe8925e2} /* (20, 10, 22) {real, imag} */,
  {32'hbcb61020, 32'h3f273318} /* (20, 10, 21) {real, imag} */,
  {32'h3e106be9, 32'h3e29207a} /* (20, 10, 20) {real, imag} */,
  {32'h3e164507, 32'h3e27cb7c} /* (20, 10, 19) {real, imag} */,
  {32'hbe5cab4e, 32'h3e6a10af} /* (20, 10, 18) {real, imag} */,
  {32'hbcc09cee, 32'hbea7f827} /* (20, 10, 17) {real, imag} */,
  {32'h3d5564f0, 32'h3e0ea540} /* (20, 10, 16) {real, imag} */,
  {32'hbc3d8420, 32'h3e0ad5d5} /* (20, 10, 15) {real, imag} */,
  {32'h3e197842, 32'h3ed8fe88} /* (20, 10, 14) {real, imag} */,
  {32'hbdbfa56e, 32'h3e9b6206} /* (20, 10, 13) {real, imag} */,
  {32'hbf4e18f8, 32'hbd48fda4} /* (20, 10, 12) {real, imag} */,
  {32'h3f1d25e4, 32'h3e211c13} /* (20, 10, 11) {real, imag} */,
  {32'h3e3d58e9, 32'h3d477aa8} /* (20, 10, 10) {real, imag} */,
  {32'hbf023fed, 32'h3cb1f9d8} /* (20, 10, 9) {real, imag} */,
  {32'h3e3b37fe, 32'h3eb3f34c} /* (20, 10, 8) {real, imag} */,
  {32'h3e1aa905, 32'h3c629f20} /* (20, 10, 7) {real, imag} */,
  {32'hbe5481f9, 32'h3c01b310} /* (20, 10, 6) {real, imag} */,
  {32'hbeb42ffc, 32'hbe26b3cb} /* (20, 10, 5) {real, imag} */,
  {32'hbd9c89e8, 32'hbf4eb1e9} /* (20, 10, 4) {real, imag} */,
  {32'h3f13f7bf, 32'h3f103d2e} /* (20, 10, 3) {real, imag} */,
  {32'h3ce14158, 32'h3e797ec8} /* (20, 10, 2) {real, imag} */,
  {32'hbdf79cbc, 32'h3e97fe50} /* (20, 10, 1) {real, imag} */,
  {32'h3e81d95e, 32'hbe773817} /* (20, 10, 0) {real, imag} */,
  {32'h3ef2084f, 32'h3edd4f54} /* (20, 9, 31) {real, imag} */,
  {32'hbe7ed538, 32'hbd8b0454} /* (20, 9, 30) {real, imag} */,
  {32'h3e562968, 32'hbe6d1324} /* (20, 9, 29) {real, imag} */,
  {32'hbef7257c, 32'hbdc1e740} /* (20, 9, 28) {real, imag} */,
  {32'hbe768727, 32'h3e6b5e42} /* (20, 9, 27) {real, imag} */,
  {32'hbec3f1db, 32'h3f044168} /* (20, 9, 26) {real, imag} */,
  {32'h3eb878ec, 32'h3e42edf5} /* (20, 9, 25) {real, imag} */,
  {32'h3dcb6008, 32'hbc178a40} /* (20, 9, 24) {real, imag} */,
  {32'hbda7bc41, 32'hbd995d68} /* (20, 9, 23) {real, imag} */,
  {32'hbee76224, 32'h3f2b7b67} /* (20, 9, 22) {real, imag} */,
  {32'hbe0f57c5, 32'hbda1eb32} /* (20, 9, 21) {real, imag} */,
  {32'h3ee0ada0, 32'hbeaec94c} /* (20, 9, 20) {real, imag} */,
  {32'hbe58d528, 32'h3e8f312d} /* (20, 9, 19) {real, imag} */,
  {32'hbed4b4d6, 32'h3dddb367} /* (20, 9, 18) {real, imag} */,
  {32'hbc5e0b84, 32'hbe38d622} /* (20, 9, 17) {real, imag} */,
  {32'hbed77ccb, 32'hbdd2d33d} /* (20, 9, 16) {real, imag} */,
  {32'h3d90260b, 32'h3db25d72} /* (20, 9, 15) {real, imag} */,
  {32'h3c9a3024, 32'hbf161592} /* (20, 9, 14) {real, imag} */,
  {32'hbe922090, 32'hbe8dd33c} /* (20, 9, 13) {real, imag} */,
  {32'h3ed8f37f, 32'hbe427bc4} /* (20, 9, 12) {real, imag} */,
  {32'h3f00427d, 32'hbe1b8a6b} /* (20, 9, 11) {real, imag} */,
  {32'hbe2cc0fc, 32'hbe6f74b1} /* (20, 9, 10) {real, imag} */,
  {32'h3e484159, 32'h3f3abc62} /* (20, 9, 9) {real, imag} */,
  {32'h3eada96f, 32'h3ec4532d} /* (20, 9, 8) {real, imag} */,
  {32'h3ddf0ea6, 32'hbdab067d} /* (20, 9, 7) {real, imag} */,
  {32'hbc0ec480, 32'h3ea3e896} /* (20, 9, 6) {real, imag} */,
  {32'hbe19fd8a, 32'h3e05e56e} /* (20, 9, 5) {real, imag} */,
  {32'hbdd7d4b7, 32'h3dc998da} /* (20, 9, 4) {real, imag} */,
  {32'h3eac8f42, 32'hbed1eab5} /* (20, 9, 3) {real, imag} */,
  {32'hbf59495c, 32'h3e749d68} /* (20, 9, 2) {real, imag} */,
  {32'hbf1e807e, 32'hbf143045} /* (20, 9, 1) {real, imag} */,
  {32'h3f0f1d57, 32'hbe5fec7e} /* (20, 9, 0) {real, imag} */,
  {32'h3fd576b6, 32'h3faa2995} /* (20, 8, 31) {real, imag} */,
  {32'hbe52b89c, 32'hbe470603} /* (20, 8, 30) {real, imag} */,
  {32'h3ebdb43e, 32'hbeda03ea} /* (20, 8, 29) {real, imag} */,
  {32'h3e3aa97f, 32'h3e551a45} /* (20, 8, 28) {real, imag} */,
  {32'hbf89ad76, 32'hbda8b10b} /* (20, 8, 27) {real, imag} */,
  {32'h3e241e9d, 32'hbec34443} /* (20, 8, 26) {real, imag} */,
  {32'h3d9bd033, 32'hbe7893ec} /* (20, 8, 25) {real, imag} */,
  {32'h3e68dfb5, 32'hbee9b4fd} /* (20, 8, 24) {real, imag} */,
  {32'hbc3f0c20, 32'hbed7cc25} /* (20, 8, 23) {real, imag} */,
  {32'hbd950460, 32'h3f3d0c72} /* (20, 8, 22) {real, imag} */,
  {32'hbebc547c, 32'hbe81a1d0} /* (20, 8, 21) {real, imag} */,
  {32'hbf366b68, 32'h3df9e564} /* (20, 8, 20) {real, imag} */,
  {32'h3ef08ddc, 32'h3dc6578a} /* (20, 8, 19) {real, imag} */,
  {32'hbdd10810, 32'h3be5fe24} /* (20, 8, 18) {real, imag} */,
  {32'hbd876cdd, 32'h3d3af460} /* (20, 8, 17) {real, imag} */,
  {32'hbdca899b, 32'h3dd8e90e} /* (20, 8, 16) {real, imag} */,
  {32'hbe92b41e, 32'h3cb3b8e8} /* (20, 8, 15) {real, imag} */,
  {32'h3b1b65c0, 32'h3deaafba} /* (20, 8, 14) {real, imag} */,
  {32'h3e0b5016, 32'h3e7f4639} /* (20, 8, 13) {real, imag} */,
  {32'hbdb085c3, 32'hbe9250c0} /* (20, 8, 12) {real, imag} */,
  {32'h3e837d76, 32'hbd4ab458} /* (20, 8, 11) {real, imag} */,
  {32'hbe99c774, 32'h3f602b54} /* (20, 8, 10) {real, imag} */,
  {32'hbed65319, 32'h3e487fce} /* (20, 8, 9) {real, imag} */,
  {32'hbf274173, 32'hbc090f20} /* (20, 8, 8) {real, imag} */,
  {32'hbf0fd401, 32'h3e46e073} /* (20, 8, 7) {real, imag} */,
  {32'hbd5b9698, 32'h3e126f15} /* (20, 8, 6) {real, imag} */,
  {32'hbf2d4317, 32'hbf26517e} /* (20, 8, 5) {real, imag} */,
  {32'h3d59e370, 32'h3e23b2f8} /* (20, 8, 4) {real, imag} */,
  {32'hbf152b94, 32'h3e7efd92} /* (20, 8, 3) {real, imag} */,
  {32'hbf9bd865, 32'hbee32e1e} /* (20, 8, 2) {real, imag} */,
  {32'h3f328eb0, 32'h3f3d2269} /* (20, 8, 1) {real, imag} */,
  {32'h3f196922, 32'hbe893043} /* (20, 8, 0) {real, imag} */,
  {32'hbf14538c, 32'hbf847887} /* (20, 7, 31) {real, imag} */,
  {32'hbc84b02c, 32'hbd2b59c0} /* (20, 7, 30) {real, imag} */,
  {32'h3ed274b2, 32'hbe86fd42} /* (20, 7, 29) {real, imag} */,
  {32'hbed30690, 32'hbe9aa057} /* (20, 7, 28) {real, imag} */,
  {32'hbeadf262, 32'h3ea7e1a2} /* (20, 7, 27) {real, imag} */,
  {32'hbd0d60a7, 32'h3dc99b02} /* (20, 7, 26) {real, imag} */,
  {32'h3cffd1e0, 32'h3f43b334} /* (20, 7, 25) {real, imag} */,
  {32'h3f0aa836, 32'h3e95f140} /* (20, 7, 24) {real, imag} */,
  {32'hbc3a6850, 32'h3ecda967} /* (20, 7, 23) {real, imag} */,
  {32'h3e365848, 32'hbdd5844c} /* (20, 7, 22) {real, imag} */,
  {32'hbee11412, 32'h3bd4ade0} /* (20, 7, 21) {real, imag} */,
  {32'hbea63f12, 32'h3ca17af8} /* (20, 7, 20) {real, imag} */,
  {32'hbd898602, 32'h3e1bc936} /* (20, 7, 19) {real, imag} */,
  {32'h3e11360c, 32'hbe85fe47} /* (20, 7, 18) {real, imag} */,
  {32'h3e2a63db, 32'h3e7d1d1a} /* (20, 7, 17) {real, imag} */,
  {32'h3d8ad124, 32'h3e232f4a} /* (20, 7, 16) {real, imag} */,
  {32'hbdfc8079, 32'h3ea5d4f3} /* (20, 7, 15) {real, imag} */,
  {32'hbea4b591, 32'h3e271608} /* (20, 7, 14) {real, imag} */,
  {32'hbdde5b02, 32'hbd26a740} /* (20, 7, 13) {real, imag} */,
  {32'h3e992869, 32'h3e91330f} /* (20, 7, 12) {real, imag} */,
  {32'hbecd1408, 32'h3e8425f6} /* (20, 7, 11) {real, imag} */,
  {32'h3eebfdc6, 32'hbe9d07d0} /* (20, 7, 10) {real, imag} */,
  {32'h3f006bbd, 32'hbe26c641} /* (20, 7, 9) {real, imag} */,
  {32'hbe9fde34, 32'h3e6be86f} /* (20, 7, 8) {real, imag} */,
  {32'hbf37ba0b, 32'h3e0fbeb4} /* (20, 7, 7) {real, imag} */,
  {32'h3e448faa, 32'hbf148d34} /* (20, 7, 6) {real, imag} */,
  {32'h3d7a5e7c, 32'h3eeab43b} /* (20, 7, 5) {real, imag} */,
  {32'h3f2e3b3a, 32'h3ea19f87} /* (20, 7, 4) {real, imag} */,
  {32'h3f0dde7a, 32'h3e223f08} /* (20, 7, 3) {real, imag} */,
  {32'hbdca37b0, 32'h3e44d278} /* (20, 7, 2) {real, imag} */,
  {32'h3eed0924, 32'hbf1174d8} /* (20, 7, 1) {real, imag} */,
  {32'hbe6b5726, 32'hbeac5a7c} /* (20, 7, 0) {real, imag} */,
  {32'hbd739f8c, 32'h3e991200} /* (20, 6, 31) {real, imag} */,
  {32'hbd962bd0, 32'hbcf56dc8} /* (20, 6, 30) {real, imag} */,
  {32'hbe5fb65a, 32'hbb881540} /* (20, 6, 29) {real, imag} */,
  {32'h3ec383ac, 32'h3ea1ed42} /* (20, 6, 28) {real, imag} */,
  {32'h3cd80858, 32'hbe953ec2} /* (20, 6, 27) {real, imag} */,
  {32'h3e2d2e0f, 32'hbf0fbd76} /* (20, 6, 26) {real, imag} */,
  {32'hbed83296, 32'hbea8ae2c} /* (20, 6, 25) {real, imag} */,
  {32'hbf15c302, 32'hbeb9b449} /* (20, 6, 24) {real, imag} */,
  {32'h3ebc6376, 32'h3f11d0f9} /* (20, 6, 23) {real, imag} */,
  {32'hbe1890a2, 32'hbf3b9990} /* (20, 6, 22) {real, imag} */,
  {32'hbea6caae, 32'hbe0cb0e0} /* (20, 6, 21) {real, imag} */,
  {32'h3ef412c6, 32'h3e3cb469} /* (20, 6, 20) {real, imag} */,
  {32'hbe8cc962, 32'hbe7dca5c} /* (20, 6, 19) {real, imag} */,
  {32'h3dd8208e, 32'h3e298e76} /* (20, 6, 18) {real, imag} */,
  {32'hbe04114e, 32'hbede10e1} /* (20, 6, 17) {real, imag} */,
  {32'h3c0752e0, 32'hbd1f5c36} /* (20, 6, 16) {real, imag} */,
  {32'h3e2c34dc, 32'hbea9451f} /* (20, 6, 15) {real, imag} */,
  {32'hbeb5d137, 32'h3ea8f46a} /* (20, 6, 14) {real, imag} */,
  {32'h3e4fc910, 32'hbf1489d4} /* (20, 6, 13) {real, imag} */,
  {32'h3e85b0c4, 32'hbe254d4b} /* (20, 6, 12) {real, imag} */,
  {32'h3dd634a1, 32'h3d7de8e2} /* (20, 6, 11) {real, imag} */,
  {32'h3b7f7b80, 32'h3e63bbb7} /* (20, 6, 10) {real, imag} */,
  {32'hbe82f89e, 32'h3eecf436} /* (20, 6, 9) {real, imag} */,
  {32'hbdb3aaf6, 32'hbd72ef68} /* (20, 6, 8) {real, imag} */,
  {32'hbf5075bc, 32'h3efe7a82} /* (20, 6, 7) {real, imag} */,
  {32'h3e0559c4, 32'hbed35b39} /* (20, 6, 6) {real, imag} */,
  {32'h3e2565ee, 32'hbe7b9868} /* (20, 6, 5) {real, imag} */,
  {32'hbe7fce53, 32'h3efd8094} /* (20, 6, 4) {real, imag} */,
  {32'h3e110e23, 32'hbf74a99a} /* (20, 6, 3) {real, imag} */,
  {32'h3e645a5f, 32'h3e692969} /* (20, 6, 2) {real, imag} */,
  {32'hbf36c592, 32'hbbe10f00} /* (20, 6, 1) {real, imag} */,
  {32'h3f19724f, 32'hbde5857e} /* (20, 6, 0) {real, imag} */,
  {32'h403a0310, 32'hbde24920} /* (20, 5, 31) {real, imag} */,
  {32'hbfd56600, 32'h3e3fd076} /* (20, 5, 30) {real, imag} */,
  {32'h3f47ef15, 32'h3f57e91f} /* (20, 5, 29) {real, imag} */,
  {32'hbdbdee38, 32'h3e123b9c} /* (20, 5, 28) {real, imag} */,
  {32'hbf2160f1, 32'hbd2d75a8} /* (20, 5, 27) {real, imag} */,
  {32'hbe45aa50, 32'hbd050c74} /* (20, 5, 26) {real, imag} */,
  {32'hbd5ba644, 32'h3eb9b508} /* (20, 5, 25) {real, imag} */,
  {32'hbe703c4d, 32'h3f4bfb54} /* (20, 5, 24) {real, imag} */,
  {32'hbecaae46, 32'h3e879192} /* (20, 5, 23) {real, imag} */,
  {32'hbf83a9a4, 32'hbd1cbb0c} /* (20, 5, 22) {real, imag} */,
  {32'h3e01416a, 32'h3dd805d9} /* (20, 5, 21) {real, imag} */,
  {32'h3e2519d0, 32'hbd302335} /* (20, 5, 20) {real, imag} */,
  {32'hbe9acfd9, 32'hbec750d3} /* (20, 5, 19) {real, imag} */,
  {32'hbe1e455f, 32'h3e2d570c} /* (20, 5, 18) {real, imag} */,
  {32'hbe87e1d6, 32'h3dd2079c} /* (20, 5, 17) {real, imag} */,
  {32'h3da2dbc4, 32'h3e6fe0ca} /* (20, 5, 16) {real, imag} */,
  {32'h3db5c1a8, 32'h3d9208f5} /* (20, 5, 15) {real, imag} */,
  {32'hbe190c06, 32'h3d90121c} /* (20, 5, 14) {real, imag} */,
  {32'hbe0c5f61, 32'hbd336870} /* (20, 5, 13) {real, imag} */,
  {32'hbe0a4af9, 32'hbf0a0554} /* (20, 5, 12) {real, imag} */,
  {32'h3ec5ee58, 32'hbf4fcdd4} /* (20, 5, 11) {real, imag} */,
  {32'h3ed3f76e, 32'h3ec6893e} /* (20, 5, 10) {real, imag} */,
  {32'hbe85d81a, 32'hbf0468f1} /* (20, 5, 9) {real, imag} */,
  {32'h3e9aa1d9, 32'h3e9c5f98} /* (20, 5, 8) {real, imag} */,
  {32'h3d90dc34, 32'h3ef30297} /* (20, 5, 7) {real, imag} */,
  {32'h3f34610c, 32'hbde7c73b} /* (20, 5, 6) {real, imag} */,
  {32'hbea55955, 32'hbebc26ca} /* (20, 5, 5) {real, imag} */,
  {32'h3f3d3304, 32'h3deb6e60} /* (20, 5, 4) {real, imag} */,
  {32'h3f0625f8, 32'h3e9b65bc} /* (20, 5, 3) {real, imag} */,
  {32'hbf60b282, 32'hbfc99bde} /* (20, 5, 2) {real, imag} */,
  {32'h3f9a6ddc, 32'h403178a3} /* (20, 5, 1) {real, imag} */,
  {32'h3fcaa5ed, 32'h400a429f} /* (20, 5, 0) {real, imag} */,
  {32'hbf7c09eb, 32'hc080e973} /* (20, 4, 31) {real, imag} */,
  {32'h40015489, 32'h400ed1b3} /* (20, 4, 30) {real, imag} */,
  {32'hbd9be250, 32'h3e13553a} /* (20, 4, 29) {real, imag} */,
  {32'hbf55c348, 32'hbc6a1da8} /* (20, 4, 28) {real, imag} */,
  {32'h3f3765e3, 32'hbf4e5344} /* (20, 4, 27) {real, imag} */,
  {32'hbf57da59, 32'hbf67de52} /* (20, 4, 26) {real, imag} */,
  {32'h3e5f4006, 32'h3ef40a7e} /* (20, 4, 25) {real, imag} */,
  {32'h3f4e0c7c, 32'hbe395d3c} /* (20, 4, 24) {real, imag} */,
  {32'hbe871c90, 32'hbe59c3c8} /* (20, 4, 23) {real, imag} */,
  {32'h3e972054, 32'hbd3e34d6} /* (20, 4, 22) {real, imag} */,
  {32'h3ec5f0c8, 32'hbeb85300} /* (20, 4, 21) {real, imag} */,
  {32'hbe1231e4, 32'h3e6dc38c} /* (20, 4, 20) {real, imag} */,
  {32'h3ee4f95c, 32'hbef10963} /* (20, 4, 19) {real, imag} */,
  {32'hbe87f912, 32'h3e217f4c} /* (20, 4, 18) {real, imag} */,
  {32'hbe94ea90, 32'h3ec22195} /* (20, 4, 17) {real, imag} */,
  {32'h3db57c39, 32'h3e4b8f34} /* (20, 4, 16) {real, imag} */,
  {32'hbde1d383, 32'hbe9fb0e2} /* (20, 4, 15) {real, imag} */,
  {32'hbe00aefa, 32'h3ec15543} /* (20, 4, 14) {real, imag} */,
  {32'h3e69202a, 32'hbc101850} /* (20, 4, 13) {real, imag} */,
  {32'hbe97bc6a, 32'h3f01bf96} /* (20, 4, 12) {real, imag} */,
  {32'hbef686de, 32'h3e78d113} /* (20, 4, 11) {real, imag} */,
  {32'hbe838bb5, 32'hbe0a5a56} /* (20, 4, 10) {real, imag} */,
  {32'hbc7fff20, 32'hbeaed022} /* (20, 4, 9) {real, imag} */,
  {32'h3d7b73e3, 32'h3bfdf100} /* (20, 4, 8) {real, imag} */,
  {32'hbe13965c, 32'hbf634184} /* (20, 4, 7) {real, imag} */,
  {32'hbf057b17, 32'h3f15999a} /* (20, 4, 6) {real, imag} */,
  {32'h3f3ea895, 32'h3f6192d6} /* (20, 4, 5) {real, imag} */,
  {32'h3d8116ac, 32'hbf09d6f4} /* (20, 4, 4) {real, imag} */,
  {32'hbf58ac38, 32'hbfa305c0} /* (20, 4, 3) {real, imag} */,
  {32'h408011c4, 32'h40210ec4} /* (20, 4, 2) {real, imag} */,
  {32'hc0866ec0, 32'hbff90c92} /* (20, 4, 1) {real, imag} */,
  {32'hc0068616, 32'hbe15598b} /* (20, 4, 0) {real, imag} */,
  {32'h4068e9b9, 32'hc05e163e} /* (20, 3, 31) {real, imag} */,
  {32'hc006b455, 32'h40849385} /* (20, 3, 30) {real, imag} */,
  {32'hbf29dbc1, 32'hbe07c5f6} /* (20, 3, 29) {real, imag} */,
  {32'hbf5d0ef2, 32'hbf94668c} /* (20, 3, 28) {real, imag} */,
  {32'hbdd8f320, 32'hbe9bab82} /* (20, 3, 27) {real, imag} */,
  {32'hbc966be4, 32'hbdf09e5c} /* (20, 3, 26) {real, imag} */,
  {32'hbf428a8f, 32'h3e3b0f46} /* (20, 3, 25) {real, imag} */,
  {32'hbe5a3a72, 32'hbdd60d08} /* (20, 3, 24) {real, imag} */,
  {32'hbd6b2830, 32'hbec616a7} /* (20, 3, 23) {real, imag} */,
  {32'hbdbdf5ce, 32'hbe2c98f4} /* (20, 3, 22) {real, imag} */,
  {32'hbe701982, 32'h3e22894e} /* (20, 3, 21) {real, imag} */,
  {32'h3e234a6a, 32'h3df7d575} /* (20, 3, 20) {real, imag} */,
  {32'hbe92c8d0, 32'h3e108d64} /* (20, 3, 19) {real, imag} */,
  {32'hbde1520e, 32'h3db6ab12} /* (20, 3, 18) {real, imag} */,
  {32'hbcb2d772, 32'hbdefcf01} /* (20, 3, 17) {real, imag} */,
  {32'hbc47b3fa, 32'hbdafec0c} /* (20, 3, 16) {real, imag} */,
  {32'hbe8762ae, 32'h3c7098e0} /* (20, 3, 15) {real, imag} */,
  {32'h3e46d120, 32'hbc836050} /* (20, 3, 14) {real, imag} */,
  {32'hbd9e7d7e, 32'h3e9596ec} /* (20, 3, 13) {real, imag} */,
  {32'h3ece70ba, 32'h3dc4cb48} /* (20, 3, 12) {real, imag} */,
  {32'hbdbe104c, 32'h3e0d39ee} /* (20, 3, 11) {real, imag} */,
  {32'h3eec316a, 32'h3e82bb29} /* (20, 3, 10) {real, imag} */,
  {32'hbeff68e8, 32'hbe65a600} /* (20, 3, 9) {real, imag} */,
  {32'hbe81bb3a, 32'h3f0aabef} /* (20, 3, 8) {real, imag} */,
  {32'h3f1d71f9, 32'h3d5d5c38} /* (20, 3, 7) {real, imag} */,
  {32'h3c3fbb60, 32'hbe9544ba} /* (20, 3, 6) {real, imag} */,
  {32'hbf214155, 32'hbce2f0e0} /* (20, 3, 5) {real, imag} */,
  {32'h3f98e171, 32'hbe858c4c} /* (20, 3, 4) {real, imag} */,
  {32'h3f9f48b2, 32'h3f08b819} /* (20, 3, 3) {real, imag} */,
  {32'h3f48b5de, 32'h4089d2aa} /* (20, 3, 2) {real, imag} */,
  {32'hc098e2c7, 32'hc02891b5} /* (20, 3, 1) {real, imag} */,
  {32'h3ea447d1, 32'h3ef4ecd2} /* (20, 3, 0) {real, imag} */,
  {32'h4220d4b0, 32'h3e193e6e} /* (20, 2, 31) {real, imag} */,
  {32'hc197a590, 32'h40d7c390} /* (20, 2, 30) {real, imag} */,
  {32'h3f924ba8, 32'hbee193bb} /* (20, 2, 29) {real, imag} */,
  {32'h3f2a320d, 32'hbfcb2e18} /* (20, 2, 28) {real, imag} */,
  {32'hbfe226ad, 32'h3d961cf0} /* (20, 2, 27) {real, imag} */,
  {32'h3f14ceed, 32'h3ec11471} /* (20, 2, 26) {real, imag} */,
  {32'h3f01bcec, 32'hbf2f8576} /* (20, 2, 25) {real, imag} */,
  {32'hbea00584, 32'h3fa43d57} /* (20, 2, 24) {real, imag} */,
  {32'h3d1ca65c, 32'hbe48728b} /* (20, 2, 23) {real, imag} */,
  {32'hbf0ec44e, 32'hbed6af92} /* (20, 2, 22) {real, imag} */,
  {32'h3cc91000, 32'h3ee8af79} /* (20, 2, 21) {real, imag} */,
  {32'h3e79e3a8, 32'hbdd43d10} /* (20, 2, 20) {real, imag} */,
  {32'hbe89cf30, 32'h3ccc6fc4} /* (20, 2, 19) {real, imag} */,
  {32'hbc716b12, 32'hbe3be3d3} /* (20, 2, 18) {real, imag} */,
  {32'hbe7b4408, 32'hbecf9bee} /* (20, 2, 17) {real, imag} */,
  {32'hbcfaeb0e, 32'hbe22dc2a} /* (20, 2, 16) {real, imag} */,
  {32'h3eb014c1, 32'hbe6d1a6a} /* (20, 2, 15) {real, imag} */,
  {32'hbee530b4, 32'hbd88d8ac} /* (20, 2, 14) {real, imag} */,
  {32'hbe84a2fa, 32'hbe552e63} /* (20, 2, 13) {real, imag} */,
  {32'h3d5586a4, 32'h3dab00d8} /* (20, 2, 12) {real, imag} */,
  {32'h3ea6570a, 32'hbea930d0} /* (20, 2, 11) {real, imag} */,
  {32'h3ed7d422, 32'h3ebee3ac} /* (20, 2, 10) {real, imag} */,
  {32'hbd0ac0e0, 32'h3ead17b2} /* (20, 2, 9) {real, imag} */,
  {32'hbf565898, 32'hbf9925f4} /* (20, 2, 8) {real, imag} */,
  {32'h3e9e8ae0, 32'h3e130a32} /* (20, 2, 7) {real, imag} */,
  {32'hbe8ce8cd, 32'hbedd3819} /* (20, 2, 6) {real, imag} */,
  {32'hc0203008, 32'hc031db17} /* (20, 2, 5) {real, imag} */,
  {32'h407f0aeb, 32'h3e5426f8} /* (20, 2, 4) {real, imag} */,
  {32'h3e9c25e9, 32'hbdc395a6} /* (20, 2, 3) {real, imag} */,
  {32'hc150d7c1, 32'h402ce058} /* (20, 2, 2) {real, imag} */,
  {32'h41c48726, 32'hc06e840f} /* (20, 2, 1) {real, imag} */,
  {32'h41a75dce, 32'h406cb550} /* (20, 2, 0) {real, imag} */,
  {32'hc25b3350, 32'h41756ab8} /* (20, 1, 31) {real, imag} */,
  {32'h416dbc2f, 32'h3f1f65a7} /* (20, 1, 30) {real, imag} */,
  {32'hbf60731e, 32'hbf659471} /* (20, 1, 29) {real, imag} */,
  {32'hc0134257, 32'hc038bb86} /* (20, 1, 28) {real, imag} */,
  {32'h4087550d, 32'h3e916d18} /* (20, 1, 27) {real, imag} */,
  {32'h3f55c249, 32'hbea39f03} /* (20, 1, 26) {real, imag} */,
  {32'hbef38d96, 32'h3f0c1ed6} /* (20, 1, 25) {real, imag} */,
  {32'hbe89d17b, 32'hbf42817c} /* (20, 1, 24) {real, imag} */,
  {32'h3bd7de40, 32'hbd9a6e88} /* (20, 1, 23) {real, imag} */,
  {32'h3e223ff6, 32'hbeef6e2e} /* (20, 1, 22) {real, imag} */,
  {32'h3eab1f1e, 32'h3e0791f8} /* (20, 1, 21) {real, imag} */,
  {32'hbe5ddfab, 32'h3e1de5f7} /* (20, 1, 20) {real, imag} */,
  {32'h3d545798, 32'hbd2dc170} /* (20, 1, 19) {real, imag} */,
  {32'h3e23aa64, 32'hbefa716a} /* (20, 1, 18) {real, imag} */,
  {32'hbe4defa8, 32'hbe369388} /* (20, 1, 17) {real, imag} */,
  {32'hbc42fef8, 32'hbe051dc0} /* (20, 1, 16) {real, imag} */,
  {32'h3e7e1e08, 32'hbe0d20ab} /* (20, 1, 15) {real, imag} */,
  {32'h3d487e42, 32'h3ed8a142} /* (20, 1, 14) {real, imag} */,
  {32'hbe084d52, 32'h3e80f278} /* (20, 1, 13) {real, imag} */,
  {32'hbe8e1ace, 32'h3e57b255} /* (20, 1, 12) {real, imag} */,
  {32'hbe0c7bdc, 32'h3f3df1d7} /* (20, 1, 11) {real, imag} */,
  {32'h3f3470f4, 32'h3e0a0fe3} /* (20, 1, 10) {real, imag} */,
  {32'h3dccb25f, 32'hbc63c4f0} /* (20, 1, 9) {real, imag} */,
  {32'h3f0a1dde, 32'h3f6990b1} /* (20, 1, 8) {real, imag} */,
  {32'hbf9a6639, 32'hbf0c1a32} /* (20, 1, 7) {real, imag} */,
  {32'h3d46d2f0, 32'h3e3bc3fa} /* (20, 1, 6) {real, imag} */,
  {32'h3ff0ad2f, 32'h3fc5485f} /* (20, 1, 5) {real, imag} */,
  {32'hbf47bd5a, 32'hc024b38c} /* (20, 1, 4) {real, imag} */,
  {32'h3fee8cc4, 32'h3f4b97e1} /* (20, 1, 3) {real, imag} */,
  {32'h418b9b13, 32'h4194fd1c} /* (20, 1, 2) {real, imag} */,
  {32'hc29b5d9d, 32'hc22444ab} /* (20, 1, 1) {real, imag} */,
  {32'hc2857347, 32'hc12791d7} /* (20, 1, 0) {real, imag} */,
  {32'hc240efc0, 32'h42146c9f} /* (20, 0, 31) {real, imag} */,
  {32'h40ccd765, 32'hc1211e89} /* (20, 0, 30) {real, imag} */,
  {32'h3ebec3b8, 32'hbf081810} /* (20, 0, 29) {real, imag} */,
  {32'hbe86c05e, 32'hbfc93621} /* (20, 0, 28) {real, imag} */,
  {32'h400202fd, 32'h3f1238cb} /* (20, 0, 27) {real, imag} */,
  {32'h3cb142a0, 32'hbf440874} /* (20, 0, 26) {real, imag} */,
  {32'hbc8cb324, 32'h3e44b2b8} /* (20, 0, 25) {real, imag} */,
  {32'hbebdc6d5, 32'hbee5ec6d} /* (20, 0, 24) {real, imag} */,
  {32'hbe829b1c, 32'h3f19dd94} /* (20, 0, 23) {real, imag} */,
  {32'hbebd798e, 32'hbeca37b4} /* (20, 0, 22) {real, imag} */,
  {32'h3ec4a080, 32'h3e330d8c} /* (20, 0, 21) {real, imag} */,
  {32'h3bbd4480, 32'hbe7e0af6} /* (20, 0, 20) {real, imag} */,
  {32'hbe0a194e, 32'hbe92fc40} /* (20, 0, 19) {real, imag} */,
  {32'h3e7ae526, 32'h3d8c5816} /* (20, 0, 18) {real, imag} */,
  {32'hbda2c801, 32'hbdaf9340} /* (20, 0, 17) {real, imag} */,
  {32'hbe723924, 32'h00000000} /* (20, 0, 16) {real, imag} */,
  {32'hbda2c801, 32'h3daf9340} /* (20, 0, 15) {real, imag} */,
  {32'h3e7ae526, 32'hbd8c5816} /* (20, 0, 14) {real, imag} */,
  {32'hbe0a194e, 32'h3e92fc40} /* (20, 0, 13) {real, imag} */,
  {32'h3bbd4480, 32'h3e7e0af6} /* (20, 0, 12) {real, imag} */,
  {32'h3ec4a080, 32'hbe330d8c} /* (20, 0, 11) {real, imag} */,
  {32'hbebd798e, 32'h3eca37b4} /* (20, 0, 10) {real, imag} */,
  {32'hbe829b1c, 32'hbf19dd94} /* (20, 0, 9) {real, imag} */,
  {32'hbebdc6d5, 32'h3ee5ec6d} /* (20, 0, 8) {real, imag} */,
  {32'hbc8cb324, 32'hbe44b2b8} /* (20, 0, 7) {real, imag} */,
  {32'h3cb142a0, 32'h3f440874} /* (20, 0, 6) {real, imag} */,
  {32'h400202fd, 32'hbf1238cb} /* (20, 0, 5) {real, imag} */,
  {32'hbe86c05e, 32'h3fc93621} /* (20, 0, 4) {real, imag} */,
  {32'h3ebec3b8, 32'h3f081810} /* (20, 0, 3) {real, imag} */,
  {32'h40ccd765, 32'h41211e89} /* (20, 0, 2) {real, imag} */,
  {32'hc240efc0, 32'hc2146c9f} /* (20, 0, 1) {real, imag} */,
  {32'hc28dc6b6, 32'h00000000} /* (20, 0, 0) {real, imag} */,
  {32'hc28d96c0, 32'h42126cb8} /* (19, 31, 31) {real, imag} */,
  {32'h418653f0, 32'hc1949d4d} /* (19, 31, 30) {real, imag} */,
  {32'h3fa7ab86, 32'h3c7ca780} /* (19, 31, 29) {real, imag} */,
  {32'hbfdac26a, 32'h3ff89b00} /* (19, 31, 28) {real, imag} */,
  {32'h3fdc707a, 32'hbf974044} /* (19, 31, 27) {real, imag} */,
  {32'h3e8db760, 32'hbdb9a8d8} /* (19, 31, 26) {real, imag} */,
  {32'hbefe6a95, 32'h3e1779ab} /* (19, 31, 25) {real, imag} */,
  {32'h3f38fbac, 32'hbf2399dc} /* (19, 31, 24) {real, imag} */,
  {32'hbf6a3b3f, 32'hbd3a1744} /* (19, 31, 23) {real, imag} */,
  {32'h3f07e204, 32'hbd271c4a} /* (19, 31, 22) {real, imag} */,
  {32'h3f46c586, 32'hbedba026} /* (19, 31, 21) {real, imag} */,
  {32'hbdfa8334, 32'hbe0d6764} /* (19, 31, 20) {real, imag} */,
  {32'hbd6172eb, 32'hbdebe5f8} /* (19, 31, 19) {real, imag} */,
  {32'hbe099036, 32'hbecc92ce} /* (19, 31, 18) {real, imag} */,
  {32'h3e48eaea, 32'h3d7c2fa4} /* (19, 31, 17) {real, imag} */,
  {32'hbdd52879, 32'h3a011980} /* (19, 31, 16) {real, imag} */,
  {32'hbe7e3945, 32'hbd2f1cfc} /* (19, 31, 15) {real, imag} */,
  {32'h3eb7e1e0, 32'h3f33eae0} /* (19, 31, 14) {real, imag} */,
  {32'h3eb263bc, 32'hbd6b920c} /* (19, 31, 13) {real, imag} */,
  {32'hbd1cf1f2, 32'hbe9e022b} /* (19, 31, 12) {real, imag} */,
  {32'h3eaaef27, 32'h3f498c38} /* (19, 31, 11) {real, imag} */,
  {32'h3e27127e, 32'hbea95a08} /* (19, 31, 10) {real, imag} */,
  {32'h3f4fccd1, 32'h3e6a1754} /* (19, 31, 9) {real, imag} */,
  {32'h3dac82e0, 32'h3ede57fb} /* (19, 31, 8) {real, imag} */,
  {32'hbec2ad45, 32'hbf763974} /* (19, 31, 7) {real, imag} */,
  {32'h3f615250, 32'h3f90711c} /* (19, 31, 6) {real, imag} */,
  {32'h4078108b, 32'hbf12529f} /* (19, 31, 5) {real, imag} */,
  {32'hc0189234, 32'h40196fae} /* (19, 31, 4) {real, imag} */,
  {32'hbf21674d, 32'h3fae63c3} /* (19, 31, 3) {real, imag} */,
  {32'h41545f5f, 32'hbf22f934} /* (19, 31, 2) {real, imag} */,
  {32'hc24755b8, 32'hc14ef1e9} /* (19, 31, 1) {real, imag} */,
  {32'hc2706f6a, 32'h411e44bc} /* (19, 31, 0) {real, imag} */,
  {32'h41b41a12, 32'h408a4c11} /* (19, 30, 31) {real, imag} */,
  {32'hc15a912f, 32'hc06f188a} /* (19, 30, 30) {real, imag} */,
  {32'h3f146dcd, 32'hbf250ed3} /* (19, 30, 29) {real, imag} */,
  {32'h4068a60e, 32'h3e8d23c2} /* (19, 30, 28) {real, imag} */,
  {32'hc017ab95, 32'h4022e8c7} /* (19, 30, 27) {real, imag} */,
  {32'h3e82c26a, 32'h3db9af58} /* (19, 30, 26) {real, imag} */,
  {32'h3e6cdc44, 32'h3ebb3f66} /* (19, 30, 25) {real, imag} */,
  {32'hbe486bd4, 32'h3fc4d424} /* (19, 30, 24) {real, imag} */,
  {32'h3e8f7533, 32'hbeab22eb} /* (19, 30, 23) {real, imag} */,
  {32'hbd66ad3e, 32'hbe8125ef} /* (19, 30, 22) {real, imag} */,
  {32'hbed3d6a8, 32'h3f4e17d4} /* (19, 30, 21) {real, imag} */,
  {32'hbeb4704e, 32'hbcfe7e2c} /* (19, 30, 20) {real, imag} */,
  {32'h3d138489, 32'hbebd4e69} /* (19, 30, 19) {real, imag} */,
  {32'h3de14566, 32'h3e325b9e} /* (19, 30, 18) {real, imag} */,
  {32'h3d3426c4, 32'hbd16e272} /* (19, 30, 17) {real, imag} */,
  {32'h3e90cbfe, 32'hbcd516bc} /* (19, 30, 16) {real, imag} */,
  {32'h3c4cef60, 32'h3ebb548b} /* (19, 30, 15) {real, imag} */,
  {32'h3e5bca44, 32'hbcf3fe7c} /* (19, 30, 14) {real, imag} */,
  {32'hbe9aa231, 32'hbd71d848} /* (19, 30, 13) {real, imag} */,
  {32'h3ecf24ed, 32'h3e9fc726} /* (19, 30, 12) {real, imag} */,
  {32'hbf3cb7f9, 32'hbf504bce} /* (19, 30, 11) {real, imag} */,
  {32'h3cf39674, 32'h3e8c3be0} /* (19, 30, 10) {real, imag} */,
  {32'hbea4df02, 32'h3f13f618} /* (19, 30, 9) {real, imag} */,
  {32'hbdce87c0, 32'hbf66da45} /* (19, 30, 8) {real, imag} */,
  {32'h3ed43815, 32'h3f931c38} /* (19, 30, 7) {real, imag} */,
  {32'hbe87fc44, 32'hbef5a83e} /* (19, 30, 6) {real, imag} */,
  {32'hbf9d8382, 32'hbe9546e2} /* (19, 30, 5) {real, imag} */,
  {32'h401139d3, 32'h4025bd74} /* (19, 30, 4) {real, imag} */,
  {32'h3fe4ebc4, 32'hbe9d3bea} /* (19, 30, 3) {real, imag} */,
  {32'hc1a00bf6, 32'hc09783a5} /* (19, 30, 2) {real, imag} */,
  {32'h42183966, 32'h3f6e873e} /* (19, 30, 1) {real, imag} */,
  {32'h41a2870c, 32'hc0527fe6} /* (19, 30, 0) {real, imag} */,
  {32'hc0787158, 32'h407fa6a3} /* (19, 29, 31) {real, imag} */,
  {32'h4010e6d0, 32'hc0844652} /* (19, 29, 30) {real, imag} */,
  {32'h3f9b4812, 32'h3e3d9077} /* (19, 29, 29) {real, imag} */,
  {32'h3f703abd, 32'hbe81f997} /* (19, 29, 28) {real, imag} */,
  {32'hbee6997b, 32'hbc8d14a0} /* (19, 29, 27) {real, imag} */,
  {32'h3ec32411, 32'h3d22c94e} /* (19, 29, 26) {real, imag} */,
  {32'hbf010248, 32'h3e27daac} /* (19, 29, 25) {real, imag} */,
  {32'h3d3f5a18, 32'hbe537ff8} /* (19, 29, 24) {real, imag} */,
  {32'h3e835da2, 32'h3f1bf923} /* (19, 29, 23) {real, imag} */,
  {32'h3e9baff1, 32'hbea13286} /* (19, 29, 22) {real, imag} */,
  {32'hbef4f227, 32'h3e99d71f} /* (19, 29, 21) {real, imag} */,
  {32'h3f27e896, 32'h3d1a2588} /* (19, 29, 20) {real, imag} */,
  {32'hbe77d880, 32'hbe7becfa} /* (19, 29, 19) {real, imag} */,
  {32'hbe872c9f, 32'hbe0b7e99} /* (19, 29, 18) {real, imag} */,
  {32'hbe9571a9, 32'h3de2bc94} /* (19, 29, 17) {real, imag} */,
  {32'hbdad0c22, 32'h3e1b5293} /* (19, 29, 16) {real, imag} */,
  {32'h3dcb5068, 32'hbe2c92ba} /* (19, 29, 15) {real, imag} */,
  {32'h3f055cd6, 32'h3e63d4e6} /* (19, 29, 14) {real, imag} */,
  {32'hbe9ef57c, 32'hbf12f3f4} /* (19, 29, 13) {real, imag} */,
  {32'h3e9ec64f, 32'h3ede5611} /* (19, 29, 12) {real, imag} */,
  {32'h3e16ccc1, 32'h3d463cec} /* (19, 29, 11) {real, imag} */,
  {32'hbf8aa34c, 32'h3f54624a} /* (19, 29, 10) {real, imag} */,
  {32'h3e31fb91, 32'hbef89852} /* (19, 29, 9) {real, imag} */,
  {32'h3eb4f57c, 32'h3d076960} /* (19, 29, 8) {real, imag} */,
  {32'hbf302a8e, 32'hbf7556e4} /* (19, 29, 7) {real, imag} */,
  {32'h3e847d8a, 32'h3e5f2cc2} /* (19, 29, 6) {real, imag} */,
  {32'hbde4b90c, 32'h3f643918} /* (19, 29, 5) {real, imag} */,
  {32'hbf373c64, 32'h3eba94d5} /* (19, 29, 4) {real, imag} */,
  {32'hbf8c2a7e, 32'h3e4bd342} /* (19, 29, 3) {real, imag} */,
  {32'hc00324c7, 32'hc0c0b34e} /* (19, 29, 2) {real, imag} */,
  {32'h406d1552, 32'h407f18b3} /* (19, 29, 1) {real, imag} */,
  {32'hbf2a1f56, 32'hbf92d83e} /* (19, 29, 0) {real, imag} */,
  {32'hc0a0ee6b, 32'h4015057c} /* (19, 28, 31) {real, imag} */,
  {32'h405b3682, 32'hc00b5a9b} /* (19, 28, 30) {real, imag} */,
  {32'hbf8c1000, 32'h3f5e74b8} /* (19, 28, 29) {real, imag} */,
  {32'h3ed42306, 32'h3ed5c51a} /* (19, 28, 28) {real, imag} */,
  {32'hbd70d1aa, 32'hbf6b6441} /* (19, 28, 27) {real, imag} */,
  {32'hbe93bf44, 32'hbe63ede6} /* (19, 28, 26) {real, imag} */,
  {32'hbe4d0f69, 32'h3dd2922e} /* (19, 28, 25) {real, imag} */,
  {32'h3e0a7c58, 32'hbe957658} /* (19, 28, 24) {real, imag} */,
  {32'h3bf547a0, 32'h3ebf77df} /* (19, 28, 23) {real, imag} */,
  {32'hbea6453a, 32'hbb74a2c0} /* (19, 28, 22) {real, imag} */,
  {32'hbeb31862, 32'hbe7c18d2} /* (19, 28, 21) {real, imag} */,
  {32'hbdc1d393, 32'h3cc1d5e0} /* (19, 28, 20) {real, imag} */,
  {32'h3f034280, 32'hbde0beea} /* (19, 28, 19) {real, imag} */,
  {32'hbe4b3354, 32'hbedff7bb} /* (19, 28, 18) {real, imag} */,
  {32'hbd0834a0, 32'h3ee555d2} /* (19, 28, 17) {real, imag} */,
  {32'hbe92da76, 32'hbd9e26ea} /* (19, 28, 16) {real, imag} */,
  {32'h3dc861d9, 32'h3e332eac} /* (19, 28, 15) {real, imag} */,
  {32'hbea641d6, 32'h3c67a820} /* (19, 28, 14) {real, imag} */,
  {32'hbe572b2e, 32'h3f538093} /* (19, 28, 13) {real, imag} */,
  {32'hbf2636ce, 32'h3e85043f} /* (19, 28, 12) {real, imag} */,
  {32'h3f1d38f9, 32'hbd8b214c} /* (19, 28, 11) {real, imag} */,
  {32'hbc955dc4, 32'hbd06a6a4} /* (19, 28, 10) {real, imag} */,
  {32'h3cbb57d0, 32'hbdf7d6aa} /* (19, 28, 9) {real, imag} */,
  {32'h3f049765, 32'h3daf96cc} /* (19, 28, 8) {real, imag} */,
  {32'h3e84e112, 32'hbf24b92a} /* (19, 28, 7) {real, imag} */,
  {32'hbf94282e, 32'h3f183514} /* (19, 28, 6) {real, imag} */,
  {32'h3fc071c9, 32'h3f806161} /* (19, 28, 5) {real, imag} */,
  {32'hbfacd552, 32'h3eb024ae} /* (19, 28, 4) {real, imag} */,
  {32'hbf0e63e5, 32'h3dc84d1e} /* (19, 28, 3) {real, imag} */,
  {32'h3fedd8de, 32'hbfeca51b} /* (19, 28, 2) {real, imag} */,
  {32'hbfa6b5c0, 32'h406efdb4} /* (19, 28, 1) {real, imag} */,
  {32'hc0119f9c, 32'h3f271882} /* (19, 28, 0) {real, imag} */,
  {32'h40026cc2, 32'hc01ceb15} /* (19, 27, 31) {real, imag} */,
  {32'hbf9a71aa, 32'h3f98a112} /* (19, 27, 30) {real, imag} */,
  {32'h3e411250, 32'hbe31ee9b} /* (19, 27, 29) {real, imag} */,
  {32'h3f38956d, 32'hbdfae328} /* (19, 27, 28) {real, imag} */,
  {32'hbfa977b9, 32'hbde36958} /* (19, 27, 27) {real, imag} */,
  {32'hbe1c9743, 32'h3f16bcec} /* (19, 27, 26) {real, imag} */,
  {32'h3fab8570, 32'h3e0b872d} /* (19, 27, 25) {real, imag} */,
  {32'hbe88b8a8, 32'h3e139f89} /* (19, 27, 24) {real, imag} */,
  {32'hbe353ed3, 32'hbf1724c7} /* (19, 27, 23) {real, imag} */,
  {32'hbe8855ff, 32'hbeeb3dec} /* (19, 27, 22) {real, imag} */,
  {32'h3e465874, 32'h3e3832c1} /* (19, 27, 21) {real, imag} */,
  {32'h3ed87bc4, 32'hbda61588} /* (19, 27, 20) {real, imag} */,
  {32'hbdcea606, 32'hbb62ff40} /* (19, 27, 19) {real, imag} */,
  {32'hba0b9d60, 32'h3e288c9d} /* (19, 27, 18) {real, imag} */,
  {32'h3e8973a9, 32'h3e4c8f5a} /* (19, 27, 17) {real, imag} */,
  {32'hbe00d748, 32'hbe9e8bc0} /* (19, 27, 16) {real, imag} */,
  {32'h3f1c751e, 32'hbe129ff2} /* (19, 27, 15) {real, imag} */,
  {32'h3e96676a, 32'hbef33c61} /* (19, 27, 14) {real, imag} */,
  {32'hbe46b7c4, 32'hbdc8c093} /* (19, 27, 13) {real, imag} */,
  {32'hbe65bf52, 32'h3ccf7918} /* (19, 27, 12) {real, imag} */,
  {32'hbe4e5fbe, 32'hbe94128f} /* (19, 27, 11) {real, imag} */,
  {32'h3d035870, 32'hbf0c5db3} /* (19, 27, 10) {real, imag} */,
  {32'hbe0496bc, 32'hbedfb443} /* (19, 27, 9) {real, imag} */,
  {32'hbeb3fd88, 32'h3f108162} /* (19, 27, 8) {real, imag} */,
  {32'h3e90cc68, 32'hbe9f1b4e} /* (19, 27, 7) {real, imag} */,
  {32'h3e5cde93, 32'hbf01fbd1} /* (19, 27, 6) {real, imag} */,
  {32'hbed45832, 32'h3e961d6b} /* (19, 27, 5) {real, imag} */,
  {32'hbf0d3c62, 32'h3e11bd70} /* (19, 27, 4) {real, imag} */,
  {32'h3f0f7300, 32'hbf872e5d} /* (19, 27, 3) {real, imag} */,
  {32'hbfc5716e, 32'hbe5b76a2} /* (19, 27, 2) {real, imag} */,
  {32'h40527f34, 32'h3ebbb466} /* (19, 27, 1) {real, imag} */,
  {32'h3fb35bde, 32'hbfa6520e} /* (19, 27, 0) {real, imag} */,
  {32'hbea0fc08, 32'h3cc87840} /* (19, 26, 31) {real, imag} */,
  {32'hbe882679, 32'h3ec602e8} /* (19, 26, 30) {real, imag} */,
  {32'h3f609a3d, 32'h3f0d7073} /* (19, 26, 29) {real, imag} */,
  {32'hbe59d17a, 32'hbf5601fe} /* (19, 26, 28) {real, imag} */,
  {32'hbef2708c, 32'h3f06b3a2} /* (19, 26, 27) {real, imag} */,
  {32'h3f74b90e, 32'h3e9c5459} /* (19, 26, 26) {real, imag} */,
  {32'h3dbf0f70, 32'hbc9d3310} /* (19, 26, 25) {real, imag} */,
  {32'hbf071d73, 32'hbf3f1688} /* (19, 26, 24) {real, imag} */,
  {32'hbf837597, 32'h3e1db860} /* (19, 26, 23) {real, imag} */,
  {32'h3e752360, 32'h3e00ff0c} /* (19, 26, 22) {real, imag} */,
  {32'hbd63397c, 32'hbe12e3d2} /* (19, 26, 21) {real, imag} */,
  {32'h3ddaf764, 32'hbb2dd860} /* (19, 26, 20) {real, imag} */,
  {32'h3de6c008, 32'hbe676597} /* (19, 26, 19) {real, imag} */,
  {32'h3e3cbb34, 32'h3f50c56e} /* (19, 26, 18) {real, imag} */,
  {32'hbe708ee4, 32'hbedaa2e1} /* (19, 26, 17) {real, imag} */,
  {32'hbd63e088, 32'hbd6bac5c} /* (19, 26, 16) {real, imag} */,
  {32'hbd5dfaa6, 32'h3e888d8c} /* (19, 26, 15) {real, imag} */,
  {32'hbecdbfe4, 32'h3f0c723a} /* (19, 26, 14) {real, imag} */,
  {32'h3e1c54c4, 32'hbd06321c} /* (19, 26, 13) {real, imag} */,
  {32'hbd24e76d, 32'h3dfb9ce0} /* (19, 26, 12) {real, imag} */,
  {32'hbe38b133, 32'hbe0e468d} /* (19, 26, 11) {real, imag} */,
  {32'h3f5c604b, 32'hbde37ecc} /* (19, 26, 10) {real, imag} */,
  {32'hbe04bc76, 32'hbecf28f3} /* (19, 26, 9) {real, imag} */,
  {32'hbefeb02c, 32'h3f2d7a0a} /* (19, 26, 8) {real, imag} */,
  {32'hbe3d4447, 32'h3db92c38} /* (19, 26, 7) {real, imag} */,
  {32'hbde91fc0, 32'h3e70c93a} /* (19, 26, 6) {real, imag} */,
  {32'hbe905c0d, 32'h3e8a4c61} /* (19, 26, 5) {real, imag} */,
  {32'h3e6eb21e, 32'hbe9007f9} /* (19, 26, 4) {real, imag} */,
  {32'hbf35c7ff, 32'hbe5e49fc} /* (19, 26, 3) {real, imag} */,
  {32'hbe72464c, 32'hbda2b9f8} /* (19, 26, 2) {real, imag} */,
  {32'hbe7efcf3, 32'h3da4e73e} /* (19, 26, 1) {real, imag} */,
  {32'hbdb0cfbc, 32'hbec8823a} /* (19, 26, 0) {real, imag} */,
  {32'hb9de3400, 32'h3f3658aa} /* (19, 25, 31) {real, imag} */,
  {32'h3eae4796, 32'hbc69cb20} /* (19, 25, 30) {real, imag} */,
  {32'h3f24558c, 32'hbe8649d7} /* (19, 25, 29) {real, imag} */,
  {32'h3e89e116, 32'h3df3b504} /* (19, 25, 28) {real, imag} */,
  {32'h3daa3790, 32'h3dba3962} /* (19, 25, 27) {real, imag} */,
  {32'h3ea3b9dc, 32'h3ea3cba5} /* (19, 25, 26) {real, imag} */,
  {32'hbf363d96, 32'hbda78ce7} /* (19, 25, 25) {real, imag} */,
  {32'hbd10fbc0, 32'hbe6ac096} /* (19, 25, 24) {real, imag} */,
  {32'h3ecaccc2, 32'h3e085364} /* (19, 25, 23) {real, imag} */,
  {32'hbeab28ca, 32'h3e1dd2fa} /* (19, 25, 22) {real, imag} */,
  {32'hbe32ef24, 32'hbdcecb51} /* (19, 25, 21) {real, imag} */,
  {32'hbd02c1f8, 32'hbce0e020} /* (19, 25, 20) {real, imag} */,
  {32'h3ec57595, 32'hbe59b97a} /* (19, 25, 19) {real, imag} */,
  {32'hbd928e4e, 32'h3e491ca8} /* (19, 25, 18) {real, imag} */,
  {32'hbdbe668a, 32'hbeb0bbc6} /* (19, 25, 17) {real, imag} */,
  {32'h3e8e8ce2, 32'h3ed90632} /* (19, 25, 16) {real, imag} */,
  {32'h3e542d9d, 32'hbe650067} /* (19, 25, 15) {real, imag} */,
  {32'h3db6562e, 32'h3e6e3590} /* (19, 25, 14) {real, imag} */,
  {32'h3be06de0, 32'h3e4839f4} /* (19, 25, 13) {real, imag} */,
  {32'hbdcd48fc, 32'hbe91f961} /* (19, 25, 12) {real, imag} */,
  {32'h3ebb2285, 32'hbd364ee0} /* (19, 25, 11) {real, imag} */,
  {32'h3e101794, 32'hbd020dd0} /* (19, 25, 10) {real, imag} */,
  {32'h3bac7680, 32'hbf603940} /* (19, 25, 9) {real, imag} */,
  {32'h3dad9db2, 32'h3ea85522} /* (19, 25, 8) {real, imag} */,
  {32'hbe8228bb, 32'h3dd179f6} /* (19, 25, 7) {real, imag} */,
  {32'hbe82eae2, 32'h3f310672} /* (19, 25, 6) {real, imag} */,
  {32'h3f374788, 32'hbef3e716} /* (19, 25, 5) {real, imag} */,
  {32'h3e36d0a4, 32'hbe93d83a} /* (19, 25, 4) {real, imag} */,
  {32'hbe9991c4, 32'h3cc21b70} /* (19, 25, 3) {real, imag} */,
  {32'h3dcfc71f, 32'hbda4536e} /* (19, 25, 2) {real, imag} */,
  {32'hbf6b5acd, 32'h3f01bdf6} /* (19, 25, 1) {real, imag} */,
  {32'hbc7b8bd0, 32'h3f5d3b81} /* (19, 25, 0) {real, imag} */,
  {32'h3f0e2444, 32'hbf8255e2} /* (19, 24, 31) {real, imag} */,
  {32'hbf882f95, 32'h3f0ed096} /* (19, 24, 30) {real, imag} */,
  {32'hbe383e9a, 32'hbe8fd540} /* (19, 24, 29) {real, imag} */,
  {32'h3f0efa06, 32'hbebd6898} /* (19, 24, 28) {real, imag} */,
  {32'h3e98e6b8, 32'h3f832d05} /* (19, 24, 27) {real, imag} */,
  {32'h3f3f9aa8, 32'h3eda923e} /* (19, 24, 26) {real, imag} */,
  {32'hbee2a11d, 32'hbb503fa0} /* (19, 24, 25) {real, imag} */,
  {32'hbf3b8c2a, 32'hbea0f158} /* (19, 24, 24) {real, imag} */,
  {32'hbe03ac35, 32'h3eb711f3} /* (19, 24, 23) {real, imag} */,
  {32'hbe5f8de7, 32'hbdf10b67} /* (19, 24, 22) {real, imag} */,
  {32'h3ea9bcd4, 32'hbebfcb1f} /* (19, 24, 21) {real, imag} */,
  {32'h3e10a3c2, 32'h3e796b16} /* (19, 24, 20) {real, imag} */,
  {32'h3d5997f6, 32'h3f24acdd} /* (19, 24, 19) {real, imag} */,
  {32'h3e4a2d5c, 32'hbeaa7baa} /* (19, 24, 18) {real, imag} */,
  {32'h3eaad4a5, 32'h3e431586} /* (19, 24, 17) {real, imag} */,
  {32'h3e5acbba, 32'hbe02309a} /* (19, 24, 16) {real, imag} */,
  {32'hbed8cf56, 32'h3e1c29ca} /* (19, 24, 15) {real, imag} */,
  {32'hbd4710e4, 32'hbe1a98fe} /* (19, 24, 14) {real, imag} */,
  {32'hbe89fffc, 32'h3e4104a2} /* (19, 24, 13) {real, imag} */,
  {32'hbe191e02, 32'h3d50f430} /* (19, 24, 12) {real, imag} */,
  {32'h3e2f03c4, 32'h3e52aca8} /* (19, 24, 11) {real, imag} */,
  {32'hbe785b2e, 32'h3d9dc874} /* (19, 24, 10) {real, imag} */,
  {32'hbedce57a, 32'hbedac673} /* (19, 24, 9) {real, imag} */,
  {32'hbeb6478e, 32'h3e64f9fc} /* (19, 24, 8) {real, imag} */,
  {32'h3e5e8cba, 32'hbdb12ed8} /* (19, 24, 7) {real, imag} */,
  {32'hbee0f108, 32'h3e1a4e03} /* (19, 24, 6) {real, imag} */,
  {32'hbf12b746, 32'hbda9de03} /* (19, 24, 5) {real, imag} */,
  {32'hbf02e730, 32'hbf5eaad3} /* (19, 24, 4) {real, imag} */,
  {32'h3c1d9940, 32'h3f2d1e17} /* (19, 24, 3) {real, imag} */,
  {32'hbf37d7d7, 32'hbe883db0} /* (19, 24, 2) {real, imag} */,
  {32'h3f8fd2ad, 32'hbf80de7d} /* (19, 24, 1) {real, imag} */,
  {32'h3f375556, 32'hbf05c36d} /* (19, 24, 0) {real, imag} */,
  {32'h3d22150c, 32'h3f4f3c73} /* (19, 23, 31) {real, imag} */,
  {32'hbe12671b, 32'hbf5122ed} /* (19, 23, 30) {real, imag} */,
  {32'hbd1e958a, 32'h3f463506} /* (19, 23, 29) {real, imag} */,
  {32'hbe8bd3ae, 32'h3e8d9e7a} /* (19, 23, 28) {real, imag} */,
  {32'h3e407476, 32'hbf24fd1e} /* (19, 23, 27) {real, imag} */,
  {32'hbb583880, 32'hbdc0b226} /* (19, 23, 26) {real, imag} */,
  {32'h3d33125a, 32'hbe01d186} /* (19, 23, 25) {real, imag} */,
  {32'hbedf6d73, 32'h3ebda109} /* (19, 23, 24) {real, imag} */,
  {32'h3d0b709c, 32'hbe8bd287} /* (19, 23, 23) {real, imag} */,
  {32'h3eced0bc, 32'h3e46b75f} /* (19, 23, 22) {real, imag} */,
  {32'h3e491ae4, 32'hbe8cbd70} /* (19, 23, 21) {real, imag} */,
  {32'hbe0bc99b, 32'h3e5b371a} /* (19, 23, 20) {real, imag} */,
  {32'hbd69368b, 32'h3edf3e17} /* (19, 23, 19) {real, imag} */,
  {32'h3e184ac4, 32'hbf0e23a2} /* (19, 23, 18) {real, imag} */,
  {32'h3e8b6aa5, 32'h3ee9c7f0} /* (19, 23, 17) {real, imag} */,
  {32'hbc9c2870, 32'hba7bc500} /* (19, 23, 16) {real, imag} */,
  {32'h3f14be80, 32'hbd5b16d0} /* (19, 23, 15) {real, imag} */,
  {32'h3cfa4d00, 32'h3e8b650e} /* (19, 23, 14) {real, imag} */,
  {32'h3e82fed6, 32'hbf2c3f02} /* (19, 23, 13) {real, imag} */,
  {32'hbd9b5161, 32'hbddf0c02} /* (19, 23, 12) {real, imag} */,
  {32'hbec97cb8, 32'hbdbe4d07} /* (19, 23, 11) {real, imag} */,
  {32'h3e85b66a, 32'hbe5e516d} /* (19, 23, 10) {real, imag} */,
  {32'hbeb53168, 32'hbe68211a} /* (19, 23, 9) {real, imag} */,
  {32'h3d9b55b6, 32'hbe9fa0e4} /* (19, 23, 8) {real, imag} */,
  {32'h3e4a7542, 32'hbe2a42b0} /* (19, 23, 7) {real, imag} */,
  {32'hbf5f7430, 32'h3e0778e4} /* (19, 23, 6) {real, imag} */,
  {32'h3e0beff2, 32'h3f6e5048} /* (19, 23, 5) {real, imag} */,
  {32'hbeae0c91, 32'h3ec9a753} /* (19, 23, 4) {real, imag} */,
  {32'h3f3acf45, 32'hbe5119b8} /* (19, 23, 3) {real, imag} */,
  {32'hbef692ab, 32'hbfaa495c} /* (19, 23, 2) {real, imag} */,
  {32'h3e10293b, 32'hbf0540ae} /* (19, 23, 1) {real, imag} */,
  {32'hbd26ea9e, 32'h3d917f98} /* (19, 23, 0) {real, imag} */,
  {32'hbe93c848, 32'h3f0630c8} /* (19, 22, 31) {real, imag} */,
  {32'h3f4464da, 32'hbec8e6c6} /* (19, 22, 30) {real, imag} */,
  {32'hbee9cde8, 32'hbe572f88} /* (19, 22, 29) {real, imag} */,
  {32'hbe903e9c, 32'h3e588846} /* (19, 22, 28) {real, imag} */,
  {32'hbee21516, 32'hbe74c836} /* (19, 22, 27) {real, imag} */,
  {32'hbf3bf721, 32'h3eb31880} /* (19, 22, 26) {real, imag} */,
  {32'hbecd1e7e, 32'h3cdc1a44} /* (19, 22, 25) {real, imag} */,
  {32'hbe13a8c0, 32'hbf631878} /* (19, 22, 24) {real, imag} */,
  {32'hbf30ae04, 32'hbe61269a} /* (19, 22, 23) {real, imag} */,
  {32'h3d132238, 32'h3e16dc3c} /* (19, 22, 22) {real, imag} */,
  {32'h3e5afb14, 32'h3e86175c} /* (19, 22, 21) {real, imag} */,
  {32'hbeef9ab0, 32'hbd7ef1d2} /* (19, 22, 20) {real, imag} */,
  {32'h3dba5e96, 32'h3e08427f} /* (19, 22, 19) {real, imag} */,
  {32'h3e9c551c, 32'hbe8002b2} /* (19, 22, 18) {real, imag} */,
  {32'hbd13924a, 32'h3aae1100} /* (19, 22, 17) {real, imag} */,
  {32'hbea60e08, 32'h3f2dfa22} /* (19, 22, 16) {real, imag} */,
  {32'hbe6b27d0, 32'h3ea61bdd} /* (19, 22, 15) {real, imag} */,
  {32'h3e88a17a, 32'hbd5410aa} /* (19, 22, 14) {real, imag} */,
  {32'h3df042b0, 32'h3df8cc50} /* (19, 22, 13) {real, imag} */,
  {32'h3ea02b04, 32'h3e097b70} /* (19, 22, 12) {real, imag} */,
  {32'h3d7ad38c, 32'hbeb37604} /* (19, 22, 11) {real, imag} */,
  {32'hbe7dce1b, 32'hbe51e272} /* (19, 22, 10) {real, imag} */,
  {32'h3c624598, 32'h3e4e695e} /* (19, 22, 9) {real, imag} */,
  {32'hbeefbf22, 32'hbee53d36} /* (19, 22, 8) {real, imag} */,
  {32'h3f1a9af9, 32'h3efff782} /* (19, 22, 7) {real, imag} */,
  {32'hbe740fc9, 32'hbe5017c7} /* (19, 22, 6) {real, imag} */,
  {32'h3e2f24ce, 32'hbcf65330} /* (19, 22, 5) {real, imag} */,
  {32'h3ed3451c, 32'hbec21426} /* (19, 22, 4) {real, imag} */,
  {32'hbeddab3e, 32'h3e796596} /* (19, 22, 3) {real, imag} */,
  {32'h3ded9b02, 32'h3f45759b} /* (19, 22, 2) {real, imag} */,
  {32'h3d4b0c1e, 32'h3e94554b} /* (19, 22, 1) {real, imag} */,
  {32'hbe553874, 32'hbb5c6040} /* (19, 22, 0) {real, imag} */,
  {32'h3c45b620, 32'hbf0eeb9d} /* (19, 21, 31) {real, imag} */,
  {32'h3e50a15e, 32'h3f00ffda} /* (19, 21, 30) {real, imag} */,
  {32'hbe95948f, 32'hbc4b1660} /* (19, 21, 29) {real, imag} */,
  {32'h3e885c22, 32'h3edb53cd} /* (19, 21, 28) {real, imag} */,
  {32'hbe2b207c, 32'h3e4a96d3} /* (19, 21, 27) {real, imag} */,
  {32'hbdc05a93, 32'h3e83153a} /* (19, 21, 26) {real, imag} */,
  {32'hbef81009, 32'hbe9ebf7a} /* (19, 21, 25) {real, imag} */,
  {32'hbe9934e6, 32'hbdf375c9} /* (19, 21, 24) {real, imag} */,
  {32'hbe78aba4, 32'h3cc3a260} /* (19, 21, 23) {real, imag} */,
  {32'hbecf4687, 32'h3e8ae2ba} /* (19, 21, 22) {real, imag} */,
  {32'h3e1ea468, 32'h3e8b0e46} /* (19, 21, 21) {real, imag} */,
  {32'hbeac722d, 32'hbeebb1d0} /* (19, 21, 20) {real, imag} */,
  {32'h3edf15b9, 32'h3e470dc6} /* (19, 21, 19) {real, imag} */,
  {32'hbea4eb35, 32'hbe59ae24} /* (19, 21, 18) {real, imag} */,
  {32'hbe7ef14d, 32'hbdb01e43} /* (19, 21, 17) {real, imag} */,
  {32'h3e7ba3b2, 32'h3e3c76c0} /* (19, 21, 16) {real, imag} */,
  {32'h3d822cc6, 32'hbc948f30} /* (19, 21, 15) {real, imag} */,
  {32'h3e9d989d, 32'h3e7d79bb} /* (19, 21, 14) {real, imag} */,
  {32'h3e23408c, 32'h3e6a76a5} /* (19, 21, 13) {real, imag} */,
  {32'h3dc2a75a, 32'h3d2bf698} /* (19, 21, 12) {real, imag} */,
  {32'h3ef910c4, 32'hbed94d54} /* (19, 21, 11) {real, imag} */,
  {32'hbe954bfb, 32'hbed3250b} /* (19, 21, 10) {real, imag} */,
  {32'h3e818724, 32'hbdd8510e} /* (19, 21, 9) {real, imag} */,
  {32'hbf292de6, 32'hbdb4740c} /* (19, 21, 8) {real, imag} */,
  {32'h3e82406f, 32'h3e9c57a1} /* (19, 21, 7) {real, imag} */,
  {32'hbe69b0ae, 32'h3e0ec48e} /* (19, 21, 6) {real, imag} */,
  {32'hbdf4f630, 32'hbeacb6a4} /* (19, 21, 5) {real, imag} */,
  {32'hbe086e32, 32'h3ead8b2a} /* (19, 21, 4) {real, imag} */,
  {32'h3ea96676, 32'h3d8f6bca} /* (19, 21, 3) {real, imag} */,
  {32'hbd7b843c, 32'h3efd4829} /* (19, 21, 2) {real, imag} */,
  {32'h3f1c2b15, 32'h3d80c507} /* (19, 21, 1) {real, imag} */,
  {32'h3f82f94f, 32'hbec3a0b4} /* (19, 21, 0) {real, imag} */,
  {32'h3ebf7ec1, 32'hbea35db8} /* (19, 20, 31) {real, imag} */,
  {32'hbd07ed54, 32'hbe2077ee} /* (19, 20, 30) {real, imag} */,
  {32'hbe829364, 32'h38d3a000} /* (19, 20, 29) {real, imag} */,
  {32'h3d95eb6a, 32'h3d72ab98} /* (19, 20, 28) {real, imag} */,
  {32'hbe380d84, 32'hbeab46f3} /* (19, 20, 27) {real, imag} */,
  {32'hbe625868, 32'h3def186a} /* (19, 20, 26) {real, imag} */,
  {32'hbe8a6874, 32'h3ea61034} /* (19, 20, 25) {real, imag} */,
  {32'h3f0247a4, 32'h3e93a01f} /* (19, 20, 24) {real, imag} */,
  {32'h3f57366f, 32'hbefd28d4} /* (19, 20, 23) {real, imag} */,
  {32'hbed6247a, 32'hbf470862} /* (19, 20, 22) {real, imag} */,
  {32'h3e8c9a4b, 32'hbe495302} /* (19, 20, 21) {real, imag} */,
  {32'h3d5c6560, 32'h3f071036} /* (19, 20, 20) {real, imag} */,
  {32'hbf2ac912, 32'hbc8183b0} /* (19, 20, 19) {real, imag} */,
  {32'h3f00672c, 32'hbd83813c} /* (19, 20, 18) {real, imag} */,
  {32'h3d6d7f40, 32'hbd8e19b7} /* (19, 20, 17) {real, imag} */,
  {32'h3e8edefb, 32'h3bbcc500} /* (19, 20, 16) {real, imag} */,
  {32'h3ecc618e, 32'hbe4adde0} /* (19, 20, 15) {real, imag} */,
  {32'hbf008b60, 32'hbeba3ac0} /* (19, 20, 14) {real, imag} */,
  {32'hbe1e240a, 32'h3f1e8a29} /* (19, 20, 13) {real, imag} */,
  {32'hbe088e42, 32'h3e05edf6} /* (19, 20, 12) {real, imag} */,
  {32'hbf477b87, 32'hbf1dc757} /* (19, 20, 11) {real, imag} */,
  {32'hbe4c6f88, 32'hbe3da914} /* (19, 20, 10) {real, imag} */,
  {32'hbd0fdcf4, 32'h3e97167d} /* (19, 20, 9) {real, imag} */,
  {32'hbe392cf4, 32'hbe546292} /* (19, 20, 8) {real, imag} */,
  {32'hbe45851e, 32'h3f0e0760} /* (19, 20, 7) {real, imag} */,
  {32'h3f19a17b, 32'hbec50c56} /* (19, 20, 6) {real, imag} */,
  {32'hbe8fc47e, 32'hbe70278f} /* (19, 20, 5) {real, imag} */,
  {32'hbf14e264, 32'h3ea8cfbc} /* (19, 20, 4) {real, imag} */,
  {32'h3e45de43, 32'hbe3fcbcd} /* (19, 20, 3) {real, imag} */,
  {32'h3e12902c, 32'h3ecc86b2} /* (19, 20, 2) {real, imag} */,
  {32'h3e3cbe93, 32'h3e62f348} /* (19, 20, 1) {real, imag} */,
  {32'h3e926f9b, 32'h3b8b3dc0} /* (19, 20, 0) {real, imag} */,
  {32'hbef4069e, 32'h3dd76d11} /* (19, 19, 31) {real, imag} */,
  {32'hbe4d7ffc, 32'h3e6f10de} /* (19, 19, 30) {real, imag} */,
  {32'h3ee9f39f, 32'hbe41722a} /* (19, 19, 29) {real, imag} */,
  {32'hbeb39fa4, 32'h3ec0c668} /* (19, 19, 28) {real, imag} */,
  {32'h3ec8ef50, 32'h3ea65b3f} /* (19, 19, 27) {real, imag} */,
  {32'h3f19d886, 32'h3c58c64e} /* (19, 19, 26) {real, imag} */,
  {32'hbd761604, 32'h3e5213ca} /* (19, 19, 25) {real, imag} */,
  {32'h3e69bb28, 32'h3d93d4eb} /* (19, 19, 24) {real, imag} */,
  {32'hbdf60be2, 32'hbeb3f26b} /* (19, 19, 23) {real, imag} */,
  {32'h3f23fbe8, 32'h3e6778da} /* (19, 19, 22) {real, imag} */,
  {32'hbda9fcf6, 32'hbf711246} /* (19, 19, 21) {real, imag} */,
  {32'h3ed7234c, 32'hbe679836} /* (19, 19, 20) {real, imag} */,
  {32'hbeb6eeb0, 32'h3ef71af0} /* (19, 19, 19) {real, imag} */,
  {32'hbec705fc, 32'h3f75cff7} /* (19, 19, 18) {real, imag} */,
  {32'h3e86cb08, 32'hbece5517} /* (19, 19, 17) {real, imag} */,
  {32'h3e0f7d66, 32'hbd86aa52} /* (19, 19, 16) {real, imag} */,
  {32'hbe6ea98c, 32'h3e3653ea} /* (19, 19, 15) {real, imag} */,
  {32'hbd7f933f, 32'h3ec43bd1} /* (19, 19, 14) {real, imag} */,
  {32'h3e901b56, 32'hbe9aa538} /* (19, 19, 13) {real, imag} */,
  {32'hbdfd495e, 32'h3e60e038} /* (19, 19, 12) {real, imag} */,
  {32'h3e31dbc8, 32'hbdeda332} /* (19, 19, 11) {real, imag} */,
  {32'h3e66ecc3, 32'hbec0c643} /* (19, 19, 10) {real, imag} */,
  {32'hbe9551e1, 32'hbd17b210} /* (19, 19, 9) {real, imag} */,
  {32'hbe874d72, 32'h3e0ddad0} /* (19, 19, 8) {real, imag} */,
  {32'h3e614886, 32'hbd6561ac} /* (19, 19, 7) {real, imag} */,
  {32'hbd3f44ae, 32'hbe8731d8} /* (19, 19, 6) {real, imag} */,
  {32'hbedd52f0, 32'hbe3fde90} /* (19, 19, 5) {real, imag} */,
  {32'hbc3b3d08, 32'h3ea53688} /* (19, 19, 4) {real, imag} */,
  {32'hbf3069ae, 32'h3eeb45ca} /* (19, 19, 3) {real, imag} */,
  {32'hbe3f7f7d, 32'hbe580e9a} /* (19, 19, 2) {real, imag} */,
  {32'h3eac7cee, 32'hbdc5dff3} /* (19, 19, 1) {real, imag} */,
  {32'h3e1a0125, 32'h3d83fafd} /* (19, 19, 0) {real, imag} */,
  {32'hbeb57247, 32'hbd304d28} /* (19, 18, 31) {real, imag} */,
  {32'h3d9843d8, 32'hbc734b48} /* (19, 18, 30) {real, imag} */,
  {32'hbd23ae4b, 32'h3d6ed308} /* (19, 18, 29) {real, imag} */,
  {32'h3e48f3aa, 32'h3dcaa9fc} /* (19, 18, 28) {real, imag} */,
  {32'hbe6e3b2d, 32'h3e59e419} /* (19, 18, 27) {real, imag} */,
  {32'hbe5af0d6, 32'h3e92f4e4} /* (19, 18, 26) {real, imag} */,
  {32'h3e999d62, 32'h3d66bb97} /* (19, 18, 25) {real, imag} */,
  {32'h3dee1f74, 32'hbe2bb1ab} /* (19, 18, 24) {real, imag} */,
  {32'hbee08d97, 32'hbdadf0c3} /* (19, 18, 23) {real, imag} */,
  {32'h3e96bcbe, 32'hbdbc2b37} /* (19, 18, 22) {real, imag} */,
  {32'h3d68795f, 32'h3e58fa54} /* (19, 18, 21) {real, imag} */,
  {32'h3dde2570, 32'h3e0b5eeb} /* (19, 18, 20) {real, imag} */,
  {32'hbe013f30, 32'hbdc1b21f} /* (19, 18, 19) {real, imag} */,
  {32'h3e4f743b, 32'h3d8d81b6} /* (19, 18, 18) {real, imag} */,
  {32'h3e8cbdbc, 32'hbd54fcae} /* (19, 18, 17) {real, imag} */,
  {32'hbe722b6a, 32'hbe71c34c} /* (19, 18, 16) {real, imag} */,
  {32'hbe27455c, 32'hbd8d88f6} /* (19, 18, 15) {real, imag} */,
  {32'hbeb25591, 32'h3d3ff004} /* (19, 18, 14) {real, imag} */,
  {32'h3e4212f8, 32'hbe64065a} /* (19, 18, 13) {real, imag} */,
  {32'h3e1cb895, 32'hbeb80ae4} /* (19, 18, 12) {real, imag} */,
  {32'h3ea856d8, 32'hbc53d1a0} /* (19, 18, 11) {real, imag} */,
  {32'h3ef521f8, 32'h3e920d88} /* (19, 18, 10) {real, imag} */,
  {32'h3eb63802, 32'h3e6430e2} /* (19, 18, 9) {real, imag} */,
  {32'h3daf73e6, 32'hbe1df35e} /* (19, 18, 8) {real, imag} */,
  {32'hbdb0162c, 32'hbe1c3e66} /* (19, 18, 7) {real, imag} */,
  {32'h3c8fb6c8, 32'hbe293c5b} /* (19, 18, 6) {real, imag} */,
  {32'h3c25df38, 32'h3d29d734} /* (19, 18, 5) {real, imag} */,
  {32'h3e26146e, 32'hbf189c20} /* (19, 18, 4) {real, imag} */,
  {32'hbdb0dc3a, 32'h3e754b02} /* (19, 18, 3) {real, imag} */,
  {32'hbb7d4c00, 32'h3e9573d5} /* (19, 18, 2) {real, imag} */,
  {32'h3ec49c92, 32'hbf231b12} /* (19, 18, 1) {real, imag} */,
  {32'hbe67542b, 32'hbcb12158} /* (19, 18, 0) {real, imag} */,
  {32'h3d3064fa, 32'h3e078794} /* (19, 17, 31) {real, imag} */,
  {32'h3da78f08, 32'hbe173695} /* (19, 17, 30) {real, imag} */,
  {32'h3d01b110, 32'hbd5e3349} /* (19, 17, 29) {real, imag} */,
  {32'h3e2baa5a, 32'h3e51f4e8} /* (19, 17, 28) {real, imag} */,
  {32'h3e420878, 32'hbdb998e2} /* (19, 17, 27) {real, imag} */,
  {32'h3ee1ea51, 32'h3f157bf0} /* (19, 17, 26) {real, imag} */,
  {32'hbd3ba038, 32'hbf10edf4} /* (19, 17, 25) {real, imag} */,
  {32'h3dbed2ff, 32'hbe144502} /* (19, 17, 24) {real, imag} */,
  {32'h3e5e79a4, 32'hbcfc9c0c} /* (19, 17, 23) {real, imag} */,
  {32'hbd35f49c, 32'h3edd87d8} /* (19, 17, 22) {real, imag} */,
  {32'h3e1b3052, 32'hbe2219ff} /* (19, 17, 21) {real, imag} */,
  {32'h3d8fd86c, 32'h3e425aef} /* (19, 17, 20) {real, imag} */,
  {32'hbd6423ac, 32'h3d018b88} /* (19, 17, 19) {real, imag} */,
  {32'hbe7e841e, 32'hbee35da4} /* (19, 17, 18) {real, imag} */,
  {32'h3e15fe80, 32'hbe978ccc} /* (19, 17, 17) {real, imag} */,
  {32'h3eaf5a5c, 32'hbdac2f82} /* (19, 17, 16) {real, imag} */,
  {32'h3dbd99cc, 32'hbe3c8a48} /* (19, 17, 15) {real, imag} */,
  {32'h3e89c8f8, 32'h3d5ad057} /* (19, 17, 14) {real, imag} */,
  {32'h3edbd79a, 32'h3e3a56e6} /* (19, 17, 13) {real, imag} */,
  {32'hbcbbd7f2, 32'h3d9dddc4} /* (19, 17, 12) {real, imag} */,
  {32'h3dec1814, 32'h3e350942} /* (19, 17, 11) {real, imag} */,
  {32'hbe220322, 32'hbe6a4a74} /* (19, 17, 10) {real, imag} */,
  {32'hbe88a09a, 32'hbe6832e6} /* (19, 17, 9) {real, imag} */,
  {32'hbd055962, 32'hbf0daf75} /* (19, 17, 8) {real, imag} */,
  {32'h3e3f5a72, 32'hbea34bd8} /* (19, 17, 7) {real, imag} */,
  {32'hbe0468b2, 32'h3e237b84} /* (19, 17, 6) {real, imag} */,
  {32'hbef2a6ff, 32'hbe68368a} /* (19, 17, 5) {real, imag} */,
  {32'h3d94dcd7, 32'h3f070ced} /* (19, 17, 4) {real, imag} */,
  {32'hbd15748d, 32'hbd3924f0} /* (19, 17, 3) {real, imag} */,
  {32'h3e4e91d1, 32'hbc23f680} /* (19, 17, 2) {real, imag} */,
  {32'h3e0547af, 32'hbd044619} /* (19, 17, 1) {real, imag} */,
  {32'h3ea67450, 32'h3e852775} /* (19, 17, 0) {real, imag} */,
  {32'hbd0a387c, 32'hbd126228} /* (19, 16, 31) {real, imag} */,
  {32'hbe2760ba, 32'h3e999406} /* (19, 16, 30) {real, imag} */,
  {32'h3dcdf51e, 32'h3de8e6dc} /* (19, 16, 29) {real, imag} */,
  {32'h3c974d75, 32'hbe0ce4a0} /* (19, 16, 28) {real, imag} */,
  {32'hbd12f174, 32'hbe1793c6} /* (19, 16, 27) {real, imag} */,
  {32'hbd78a327, 32'hbec903ac} /* (19, 16, 26) {real, imag} */,
  {32'h3e26d7d3, 32'h3e2e8fda} /* (19, 16, 25) {real, imag} */,
  {32'hbe918ea6, 32'h3deb9f25} /* (19, 16, 24) {real, imag} */,
  {32'hbd8b0f53, 32'hbea1f3cb} /* (19, 16, 23) {real, imag} */,
  {32'h3e0c08e6, 32'hbe2925d5} /* (19, 16, 22) {real, imag} */,
  {32'hbe913fc5, 32'h3d85a732} /* (19, 16, 21) {real, imag} */,
  {32'hbd808007, 32'h3da52550} /* (19, 16, 20) {real, imag} */,
  {32'hbe9777f4, 32'hbe4fd009} /* (19, 16, 19) {real, imag} */,
  {32'h3e2f2db4, 32'hbe522232} /* (19, 16, 18) {real, imag} */,
  {32'hbe912631, 32'hbcf403fa} /* (19, 16, 17) {real, imag} */,
  {32'hbe29cc10, 32'h00000000} /* (19, 16, 16) {real, imag} */,
  {32'hbe912631, 32'h3cf403fa} /* (19, 16, 15) {real, imag} */,
  {32'h3e2f2db4, 32'h3e522232} /* (19, 16, 14) {real, imag} */,
  {32'hbe9777f4, 32'h3e4fd009} /* (19, 16, 13) {real, imag} */,
  {32'hbd808007, 32'hbda52550} /* (19, 16, 12) {real, imag} */,
  {32'hbe913fc5, 32'hbd85a732} /* (19, 16, 11) {real, imag} */,
  {32'h3e0c08e6, 32'h3e2925d5} /* (19, 16, 10) {real, imag} */,
  {32'hbd8b0f53, 32'h3ea1f3cb} /* (19, 16, 9) {real, imag} */,
  {32'hbe918ea6, 32'hbdeb9f25} /* (19, 16, 8) {real, imag} */,
  {32'h3e26d7d3, 32'hbe2e8fda} /* (19, 16, 7) {real, imag} */,
  {32'hbd78a327, 32'h3ec903ac} /* (19, 16, 6) {real, imag} */,
  {32'hbd12f174, 32'h3e1793c6} /* (19, 16, 5) {real, imag} */,
  {32'h3c974d75, 32'h3e0ce4a0} /* (19, 16, 4) {real, imag} */,
  {32'h3dcdf51e, 32'hbde8e6dc} /* (19, 16, 3) {real, imag} */,
  {32'hbe2760ba, 32'hbe999406} /* (19, 16, 2) {real, imag} */,
  {32'hbd0a387c, 32'h3d126228} /* (19, 16, 1) {real, imag} */,
  {32'hbea1e5d3, 32'h00000000} /* (19, 16, 0) {real, imag} */,
  {32'h3e0547af, 32'h3d044619} /* (19, 15, 31) {real, imag} */,
  {32'h3e4e91d1, 32'h3c23f680} /* (19, 15, 30) {real, imag} */,
  {32'hbd15748d, 32'h3d3924f0} /* (19, 15, 29) {real, imag} */,
  {32'h3d94dcd7, 32'hbf070ced} /* (19, 15, 28) {real, imag} */,
  {32'hbef2a6ff, 32'h3e68368a} /* (19, 15, 27) {real, imag} */,
  {32'hbe0468b2, 32'hbe237b84} /* (19, 15, 26) {real, imag} */,
  {32'h3e3f5a72, 32'h3ea34bd8} /* (19, 15, 25) {real, imag} */,
  {32'hbd055962, 32'h3f0daf75} /* (19, 15, 24) {real, imag} */,
  {32'hbe88a09a, 32'h3e6832e6} /* (19, 15, 23) {real, imag} */,
  {32'hbe220322, 32'h3e6a4a74} /* (19, 15, 22) {real, imag} */,
  {32'h3dec1814, 32'hbe350942} /* (19, 15, 21) {real, imag} */,
  {32'hbcbbd7f2, 32'hbd9dddc4} /* (19, 15, 20) {real, imag} */,
  {32'h3edbd79a, 32'hbe3a56e6} /* (19, 15, 19) {real, imag} */,
  {32'h3e89c8f8, 32'hbd5ad057} /* (19, 15, 18) {real, imag} */,
  {32'h3dbd99cc, 32'h3e3c8a48} /* (19, 15, 17) {real, imag} */,
  {32'h3eaf5a5c, 32'h3dac2f82} /* (19, 15, 16) {real, imag} */,
  {32'h3e15fe80, 32'h3e978ccc} /* (19, 15, 15) {real, imag} */,
  {32'hbe7e841e, 32'h3ee35da4} /* (19, 15, 14) {real, imag} */,
  {32'hbd6423ac, 32'hbd018b88} /* (19, 15, 13) {real, imag} */,
  {32'h3d8fd86c, 32'hbe425aef} /* (19, 15, 12) {real, imag} */,
  {32'h3e1b3052, 32'h3e2219ff} /* (19, 15, 11) {real, imag} */,
  {32'hbd35f49c, 32'hbedd87d8} /* (19, 15, 10) {real, imag} */,
  {32'h3e5e79a4, 32'h3cfc9c0c} /* (19, 15, 9) {real, imag} */,
  {32'h3dbed2ff, 32'h3e144502} /* (19, 15, 8) {real, imag} */,
  {32'hbd3ba038, 32'h3f10edf4} /* (19, 15, 7) {real, imag} */,
  {32'h3ee1ea51, 32'hbf157bf0} /* (19, 15, 6) {real, imag} */,
  {32'h3e420878, 32'h3db998e2} /* (19, 15, 5) {real, imag} */,
  {32'h3e2baa5a, 32'hbe51f4e8} /* (19, 15, 4) {real, imag} */,
  {32'h3d01b110, 32'h3d5e3349} /* (19, 15, 3) {real, imag} */,
  {32'h3da78f08, 32'h3e173695} /* (19, 15, 2) {real, imag} */,
  {32'h3d3064fa, 32'hbe078794} /* (19, 15, 1) {real, imag} */,
  {32'h3ea67450, 32'hbe852775} /* (19, 15, 0) {real, imag} */,
  {32'h3ec49c92, 32'h3f231b12} /* (19, 14, 31) {real, imag} */,
  {32'hbb7d4c00, 32'hbe9573d5} /* (19, 14, 30) {real, imag} */,
  {32'hbdb0dc3a, 32'hbe754b02} /* (19, 14, 29) {real, imag} */,
  {32'h3e26146e, 32'h3f189c20} /* (19, 14, 28) {real, imag} */,
  {32'h3c25df38, 32'hbd29d734} /* (19, 14, 27) {real, imag} */,
  {32'h3c8fb6c8, 32'h3e293c5b} /* (19, 14, 26) {real, imag} */,
  {32'hbdb0162c, 32'h3e1c3e66} /* (19, 14, 25) {real, imag} */,
  {32'h3daf73e6, 32'h3e1df35e} /* (19, 14, 24) {real, imag} */,
  {32'h3eb63802, 32'hbe6430e2} /* (19, 14, 23) {real, imag} */,
  {32'h3ef521f8, 32'hbe920d88} /* (19, 14, 22) {real, imag} */,
  {32'h3ea856d8, 32'h3c53d1a0} /* (19, 14, 21) {real, imag} */,
  {32'h3e1cb895, 32'h3eb80ae4} /* (19, 14, 20) {real, imag} */,
  {32'h3e4212f8, 32'h3e64065a} /* (19, 14, 19) {real, imag} */,
  {32'hbeb25591, 32'hbd3ff004} /* (19, 14, 18) {real, imag} */,
  {32'hbe27455c, 32'h3d8d88f6} /* (19, 14, 17) {real, imag} */,
  {32'hbe722b6a, 32'h3e71c34c} /* (19, 14, 16) {real, imag} */,
  {32'h3e8cbdbc, 32'h3d54fcae} /* (19, 14, 15) {real, imag} */,
  {32'h3e4f743b, 32'hbd8d81b6} /* (19, 14, 14) {real, imag} */,
  {32'hbe013f30, 32'h3dc1b21f} /* (19, 14, 13) {real, imag} */,
  {32'h3dde2570, 32'hbe0b5eeb} /* (19, 14, 12) {real, imag} */,
  {32'h3d68795f, 32'hbe58fa54} /* (19, 14, 11) {real, imag} */,
  {32'h3e96bcbe, 32'h3dbc2b37} /* (19, 14, 10) {real, imag} */,
  {32'hbee08d97, 32'h3dadf0c3} /* (19, 14, 9) {real, imag} */,
  {32'h3dee1f74, 32'h3e2bb1ab} /* (19, 14, 8) {real, imag} */,
  {32'h3e999d62, 32'hbd66bb97} /* (19, 14, 7) {real, imag} */,
  {32'hbe5af0d6, 32'hbe92f4e4} /* (19, 14, 6) {real, imag} */,
  {32'hbe6e3b2d, 32'hbe59e419} /* (19, 14, 5) {real, imag} */,
  {32'h3e48f3aa, 32'hbdcaa9fc} /* (19, 14, 4) {real, imag} */,
  {32'hbd23ae4b, 32'hbd6ed308} /* (19, 14, 3) {real, imag} */,
  {32'h3d9843d8, 32'h3c734b48} /* (19, 14, 2) {real, imag} */,
  {32'hbeb57247, 32'h3d304d28} /* (19, 14, 1) {real, imag} */,
  {32'hbe67542b, 32'h3cb12158} /* (19, 14, 0) {real, imag} */,
  {32'h3eac7cee, 32'h3dc5dff3} /* (19, 13, 31) {real, imag} */,
  {32'hbe3f7f7d, 32'h3e580e9a} /* (19, 13, 30) {real, imag} */,
  {32'hbf3069ae, 32'hbeeb45ca} /* (19, 13, 29) {real, imag} */,
  {32'hbc3b3d08, 32'hbea53688} /* (19, 13, 28) {real, imag} */,
  {32'hbedd52f0, 32'h3e3fde90} /* (19, 13, 27) {real, imag} */,
  {32'hbd3f44ae, 32'h3e8731d8} /* (19, 13, 26) {real, imag} */,
  {32'h3e614886, 32'h3d6561ac} /* (19, 13, 25) {real, imag} */,
  {32'hbe874d72, 32'hbe0ddad0} /* (19, 13, 24) {real, imag} */,
  {32'hbe9551e1, 32'h3d17b210} /* (19, 13, 23) {real, imag} */,
  {32'h3e66ecc3, 32'h3ec0c643} /* (19, 13, 22) {real, imag} */,
  {32'h3e31dbc8, 32'h3deda332} /* (19, 13, 21) {real, imag} */,
  {32'hbdfd495e, 32'hbe60e038} /* (19, 13, 20) {real, imag} */,
  {32'h3e901b56, 32'h3e9aa538} /* (19, 13, 19) {real, imag} */,
  {32'hbd7f933f, 32'hbec43bd1} /* (19, 13, 18) {real, imag} */,
  {32'hbe6ea98c, 32'hbe3653ea} /* (19, 13, 17) {real, imag} */,
  {32'h3e0f7d66, 32'h3d86aa52} /* (19, 13, 16) {real, imag} */,
  {32'h3e86cb08, 32'h3ece5517} /* (19, 13, 15) {real, imag} */,
  {32'hbec705fc, 32'hbf75cff7} /* (19, 13, 14) {real, imag} */,
  {32'hbeb6eeb0, 32'hbef71af0} /* (19, 13, 13) {real, imag} */,
  {32'h3ed7234c, 32'h3e679836} /* (19, 13, 12) {real, imag} */,
  {32'hbda9fcf6, 32'h3f711246} /* (19, 13, 11) {real, imag} */,
  {32'h3f23fbe8, 32'hbe6778da} /* (19, 13, 10) {real, imag} */,
  {32'hbdf60be2, 32'h3eb3f26b} /* (19, 13, 9) {real, imag} */,
  {32'h3e69bb28, 32'hbd93d4eb} /* (19, 13, 8) {real, imag} */,
  {32'hbd761604, 32'hbe5213ca} /* (19, 13, 7) {real, imag} */,
  {32'h3f19d886, 32'hbc58c64e} /* (19, 13, 6) {real, imag} */,
  {32'h3ec8ef50, 32'hbea65b3f} /* (19, 13, 5) {real, imag} */,
  {32'hbeb39fa4, 32'hbec0c668} /* (19, 13, 4) {real, imag} */,
  {32'h3ee9f39f, 32'h3e41722a} /* (19, 13, 3) {real, imag} */,
  {32'hbe4d7ffc, 32'hbe6f10de} /* (19, 13, 2) {real, imag} */,
  {32'hbef4069e, 32'hbdd76d11} /* (19, 13, 1) {real, imag} */,
  {32'h3e1a0125, 32'hbd83fafd} /* (19, 13, 0) {real, imag} */,
  {32'h3e3cbe93, 32'hbe62f348} /* (19, 12, 31) {real, imag} */,
  {32'h3e12902c, 32'hbecc86b2} /* (19, 12, 30) {real, imag} */,
  {32'h3e45de43, 32'h3e3fcbcd} /* (19, 12, 29) {real, imag} */,
  {32'hbf14e264, 32'hbea8cfbc} /* (19, 12, 28) {real, imag} */,
  {32'hbe8fc47e, 32'h3e70278f} /* (19, 12, 27) {real, imag} */,
  {32'h3f19a17b, 32'h3ec50c56} /* (19, 12, 26) {real, imag} */,
  {32'hbe45851e, 32'hbf0e0760} /* (19, 12, 25) {real, imag} */,
  {32'hbe392cf4, 32'h3e546292} /* (19, 12, 24) {real, imag} */,
  {32'hbd0fdcf4, 32'hbe97167d} /* (19, 12, 23) {real, imag} */,
  {32'hbe4c6f88, 32'h3e3da914} /* (19, 12, 22) {real, imag} */,
  {32'hbf477b87, 32'h3f1dc757} /* (19, 12, 21) {real, imag} */,
  {32'hbe088e42, 32'hbe05edf6} /* (19, 12, 20) {real, imag} */,
  {32'hbe1e240a, 32'hbf1e8a29} /* (19, 12, 19) {real, imag} */,
  {32'hbf008b60, 32'h3eba3ac0} /* (19, 12, 18) {real, imag} */,
  {32'h3ecc618e, 32'h3e4adde0} /* (19, 12, 17) {real, imag} */,
  {32'h3e8edefb, 32'hbbbcc500} /* (19, 12, 16) {real, imag} */,
  {32'h3d6d7f40, 32'h3d8e19b7} /* (19, 12, 15) {real, imag} */,
  {32'h3f00672c, 32'h3d83813c} /* (19, 12, 14) {real, imag} */,
  {32'hbf2ac912, 32'h3c8183b0} /* (19, 12, 13) {real, imag} */,
  {32'h3d5c6560, 32'hbf071036} /* (19, 12, 12) {real, imag} */,
  {32'h3e8c9a4b, 32'h3e495302} /* (19, 12, 11) {real, imag} */,
  {32'hbed6247a, 32'h3f470862} /* (19, 12, 10) {real, imag} */,
  {32'h3f57366f, 32'h3efd28d4} /* (19, 12, 9) {real, imag} */,
  {32'h3f0247a4, 32'hbe93a01f} /* (19, 12, 8) {real, imag} */,
  {32'hbe8a6874, 32'hbea61034} /* (19, 12, 7) {real, imag} */,
  {32'hbe625868, 32'hbdef186a} /* (19, 12, 6) {real, imag} */,
  {32'hbe380d84, 32'h3eab46f3} /* (19, 12, 5) {real, imag} */,
  {32'h3d95eb6a, 32'hbd72ab98} /* (19, 12, 4) {real, imag} */,
  {32'hbe829364, 32'hb8d3a000} /* (19, 12, 3) {real, imag} */,
  {32'hbd07ed54, 32'h3e2077ee} /* (19, 12, 2) {real, imag} */,
  {32'h3ebf7ec1, 32'h3ea35db8} /* (19, 12, 1) {real, imag} */,
  {32'h3e926f9b, 32'hbb8b3dc0} /* (19, 12, 0) {real, imag} */,
  {32'h3f1c2b15, 32'hbd80c507} /* (19, 11, 31) {real, imag} */,
  {32'hbd7b843c, 32'hbefd4829} /* (19, 11, 30) {real, imag} */,
  {32'h3ea96676, 32'hbd8f6bca} /* (19, 11, 29) {real, imag} */,
  {32'hbe086e32, 32'hbead8b2a} /* (19, 11, 28) {real, imag} */,
  {32'hbdf4f630, 32'h3eacb6a4} /* (19, 11, 27) {real, imag} */,
  {32'hbe69b0ae, 32'hbe0ec48e} /* (19, 11, 26) {real, imag} */,
  {32'h3e82406f, 32'hbe9c57a1} /* (19, 11, 25) {real, imag} */,
  {32'hbf292de6, 32'h3db4740c} /* (19, 11, 24) {real, imag} */,
  {32'h3e818724, 32'h3dd8510e} /* (19, 11, 23) {real, imag} */,
  {32'hbe954bfb, 32'h3ed3250b} /* (19, 11, 22) {real, imag} */,
  {32'h3ef910c4, 32'h3ed94d54} /* (19, 11, 21) {real, imag} */,
  {32'h3dc2a75a, 32'hbd2bf698} /* (19, 11, 20) {real, imag} */,
  {32'h3e23408c, 32'hbe6a76a5} /* (19, 11, 19) {real, imag} */,
  {32'h3e9d989d, 32'hbe7d79bb} /* (19, 11, 18) {real, imag} */,
  {32'h3d822cc6, 32'h3c948f30} /* (19, 11, 17) {real, imag} */,
  {32'h3e7ba3b2, 32'hbe3c76c0} /* (19, 11, 16) {real, imag} */,
  {32'hbe7ef14d, 32'h3db01e43} /* (19, 11, 15) {real, imag} */,
  {32'hbea4eb35, 32'h3e59ae24} /* (19, 11, 14) {real, imag} */,
  {32'h3edf15b9, 32'hbe470dc6} /* (19, 11, 13) {real, imag} */,
  {32'hbeac722d, 32'h3eebb1d0} /* (19, 11, 12) {real, imag} */,
  {32'h3e1ea468, 32'hbe8b0e46} /* (19, 11, 11) {real, imag} */,
  {32'hbecf4687, 32'hbe8ae2ba} /* (19, 11, 10) {real, imag} */,
  {32'hbe78aba4, 32'hbcc3a260} /* (19, 11, 9) {real, imag} */,
  {32'hbe9934e6, 32'h3df375c9} /* (19, 11, 8) {real, imag} */,
  {32'hbef81009, 32'h3e9ebf7a} /* (19, 11, 7) {real, imag} */,
  {32'hbdc05a93, 32'hbe83153a} /* (19, 11, 6) {real, imag} */,
  {32'hbe2b207c, 32'hbe4a96d3} /* (19, 11, 5) {real, imag} */,
  {32'h3e885c22, 32'hbedb53cd} /* (19, 11, 4) {real, imag} */,
  {32'hbe95948f, 32'h3c4b1660} /* (19, 11, 3) {real, imag} */,
  {32'h3e50a15e, 32'hbf00ffda} /* (19, 11, 2) {real, imag} */,
  {32'h3c45b620, 32'h3f0eeb9d} /* (19, 11, 1) {real, imag} */,
  {32'h3f82f94f, 32'h3ec3a0b4} /* (19, 11, 0) {real, imag} */,
  {32'h3d4b0c1e, 32'hbe94554b} /* (19, 10, 31) {real, imag} */,
  {32'h3ded9b02, 32'hbf45759b} /* (19, 10, 30) {real, imag} */,
  {32'hbeddab3e, 32'hbe796596} /* (19, 10, 29) {real, imag} */,
  {32'h3ed3451c, 32'h3ec21426} /* (19, 10, 28) {real, imag} */,
  {32'h3e2f24ce, 32'h3cf65330} /* (19, 10, 27) {real, imag} */,
  {32'hbe740fc9, 32'h3e5017c7} /* (19, 10, 26) {real, imag} */,
  {32'h3f1a9af9, 32'hbefff782} /* (19, 10, 25) {real, imag} */,
  {32'hbeefbf22, 32'h3ee53d36} /* (19, 10, 24) {real, imag} */,
  {32'h3c624598, 32'hbe4e695e} /* (19, 10, 23) {real, imag} */,
  {32'hbe7dce1b, 32'h3e51e272} /* (19, 10, 22) {real, imag} */,
  {32'h3d7ad38c, 32'h3eb37604} /* (19, 10, 21) {real, imag} */,
  {32'h3ea02b04, 32'hbe097b70} /* (19, 10, 20) {real, imag} */,
  {32'h3df042b0, 32'hbdf8cc50} /* (19, 10, 19) {real, imag} */,
  {32'h3e88a17a, 32'h3d5410aa} /* (19, 10, 18) {real, imag} */,
  {32'hbe6b27d0, 32'hbea61bdd} /* (19, 10, 17) {real, imag} */,
  {32'hbea60e08, 32'hbf2dfa22} /* (19, 10, 16) {real, imag} */,
  {32'hbd13924a, 32'hbaae1100} /* (19, 10, 15) {real, imag} */,
  {32'h3e9c551c, 32'h3e8002b2} /* (19, 10, 14) {real, imag} */,
  {32'h3dba5e96, 32'hbe08427f} /* (19, 10, 13) {real, imag} */,
  {32'hbeef9ab0, 32'h3d7ef1d2} /* (19, 10, 12) {real, imag} */,
  {32'h3e5afb14, 32'hbe86175c} /* (19, 10, 11) {real, imag} */,
  {32'h3d132238, 32'hbe16dc3c} /* (19, 10, 10) {real, imag} */,
  {32'hbf30ae04, 32'h3e61269a} /* (19, 10, 9) {real, imag} */,
  {32'hbe13a8c0, 32'h3f631878} /* (19, 10, 8) {real, imag} */,
  {32'hbecd1e7e, 32'hbcdc1a44} /* (19, 10, 7) {real, imag} */,
  {32'hbf3bf721, 32'hbeb31880} /* (19, 10, 6) {real, imag} */,
  {32'hbee21516, 32'h3e74c836} /* (19, 10, 5) {real, imag} */,
  {32'hbe903e9c, 32'hbe588846} /* (19, 10, 4) {real, imag} */,
  {32'hbee9cde8, 32'h3e572f88} /* (19, 10, 3) {real, imag} */,
  {32'h3f4464da, 32'h3ec8e6c6} /* (19, 10, 2) {real, imag} */,
  {32'hbe93c848, 32'hbf0630c8} /* (19, 10, 1) {real, imag} */,
  {32'hbe553874, 32'h3b5c6040} /* (19, 10, 0) {real, imag} */,
  {32'h3e10293b, 32'h3f0540ae} /* (19, 9, 31) {real, imag} */,
  {32'hbef692ab, 32'h3faa495c} /* (19, 9, 30) {real, imag} */,
  {32'h3f3acf45, 32'h3e5119b8} /* (19, 9, 29) {real, imag} */,
  {32'hbeae0c91, 32'hbec9a753} /* (19, 9, 28) {real, imag} */,
  {32'h3e0beff2, 32'hbf6e5048} /* (19, 9, 27) {real, imag} */,
  {32'hbf5f7430, 32'hbe0778e4} /* (19, 9, 26) {real, imag} */,
  {32'h3e4a7542, 32'h3e2a42b0} /* (19, 9, 25) {real, imag} */,
  {32'h3d9b55b6, 32'h3e9fa0e4} /* (19, 9, 24) {real, imag} */,
  {32'hbeb53168, 32'h3e68211a} /* (19, 9, 23) {real, imag} */,
  {32'h3e85b66a, 32'h3e5e516d} /* (19, 9, 22) {real, imag} */,
  {32'hbec97cb8, 32'h3dbe4d07} /* (19, 9, 21) {real, imag} */,
  {32'hbd9b5161, 32'h3ddf0c02} /* (19, 9, 20) {real, imag} */,
  {32'h3e82fed6, 32'h3f2c3f02} /* (19, 9, 19) {real, imag} */,
  {32'h3cfa4d00, 32'hbe8b650e} /* (19, 9, 18) {real, imag} */,
  {32'h3f14be80, 32'h3d5b16d0} /* (19, 9, 17) {real, imag} */,
  {32'hbc9c2870, 32'h3a7bc500} /* (19, 9, 16) {real, imag} */,
  {32'h3e8b6aa5, 32'hbee9c7f0} /* (19, 9, 15) {real, imag} */,
  {32'h3e184ac4, 32'h3f0e23a2} /* (19, 9, 14) {real, imag} */,
  {32'hbd69368b, 32'hbedf3e17} /* (19, 9, 13) {real, imag} */,
  {32'hbe0bc99b, 32'hbe5b371a} /* (19, 9, 12) {real, imag} */,
  {32'h3e491ae4, 32'h3e8cbd70} /* (19, 9, 11) {real, imag} */,
  {32'h3eced0bc, 32'hbe46b75f} /* (19, 9, 10) {real, imag} */,
  {32'h3d0b709c, 32'h3e8bd287} /* (19, 9, 9) {real, imag} */,
  {32'hbedf6d73, 32'hbebda109} /* (19, 9, 8) {real, imag} */,
  {32'h3d33125a, 32'h3e01d186} /* (19, 9, 7) {real, imag} */,
  {32'hbb583880, 32'h3dc0b226} /* (19, 9, 6) {real, imag} */,
  {32'h3e407476, 32'h3f24fd1e} /* (19, 9, 5) {real, imag} */,
  {32'hbe8bd3ae, 32'hbe8d9e7a} /* (19, 9, 4) {real, imag} */,
  {32'hbd1e958a, 32'hbf463506} /* (19, 9, 3) {real, imag} */,
  {32'hbe12671b, 32'h3f5122ed} /* (19, 9, 2) {real, imag} */,
  {32'h3d22150c, 32'hbf4f3c73} /* (19, 9, 1) {real, imag} */,
  {32'hbd26ea9e, 32'hbd917f98} /* (19, 9, 0) {real, imag} */,
  {32'h3f8fd2ad, 32'h3f80de7d} /* (19, 8, 31) {real, imag} */,
  {32'hbf37d7d7, 32'h3e883db0} /* (19, 8, 30) {real, imag} */,
  {32'h3c1d9940, 32'hbf2d1e17} /* (19, 8, 29) {real, imag} */,
  {32'hbf02e730, 32'h3f5eaad3} /* (19, 8, 28) {real, imag} */,
  {32'hbf12b746, 32'h3da9de03} /* (19, 8, 27) {real, imag} */,
  {32'hbee0f108, 32'hbe1a4e03} /* (19, 8, 26) {real, imag} */,
  {32'h3e5e8cba, 32'h3db12ed8} /* (19, 8, 25) {real, imag} */,
  {32'hbeb6478e, 32'hbe64f9fc} /* (19, 8, 24) {real, imag} */,
  {32'hbedce57a, 32'h3edac673} /* (19, 8, 23) {real, imag} */,
  {32'hbe785b2e, 32'hbd9dc874} /* (19, 8, 22) {real, imag} */,
  {32'h3e2f03c4, 32'hbe52aca8} /* (19, 8, 21) {real, imag} */,
  {32'hbe191e02, 32'hbd50f430} /* (19, 8, 20) {real, imag} */,
  {32'hbe89fffc, 32'hbe4104a2} /* (19, 8, 19) {real, imag} */,
  {32'hbd4710e4, 32'h3e1a98fe} /* (19, 8, 18) {real, imag} */,
  {32'hbed8cf56, 32'hbe1c29ca} /* (19, 8, 17) {real, imag} */,
  {32'h3e5acbba, 32'h3e02309a} /* (19, 8, 16) {real, imag} */,
  {32'h3eaad4a5, 32'hbe431586} /* (19, 8, 15) {real, imag} */,
  {32'h3e4a2d5c, 32'h3eaa7baa} /* (19, 8, 14) {real, imag} */,
  {32'h3d5997f6, 32'hbf24acdd} /* (19, 8, 13) {real, imag} */,
  {32'h3e10a3c2, 32'hbe796b16} /* (19, 8, 12) {real, imag} */,
  {32'h3ea9bcd4, 32'h3ebfcb1f} /* (19, 8, 11) {real, imag} */,
  {32'hbe5f8de7, 32'h3df10b67} /* (19, 8, 10) {real, imag} */,
  {32'hbe03ac35, 32'hbeb711f3} /* (19, 8, 9) {real, imag} */,
  {32'hbf3b8c2a, 32'h3ea0f158} /* (19, 8, 8) {real, imag} */,
  {32'hbee2a11d, 32'h3b503fa0} /* (19, 8, 7) {real, imag} */,
  {32'h3f3f9aa8, 32'hbeda923e} /* (19, 8, 6) {real, imag} */,
  {32'h3e98e6b8, 32'hbf832d05} /* (19, 8, 5) {real, imag} */,
  {32'h3f0efa06, 32'h3ebd6898} /* (19, 8, 4) {real, imag} */,
  {32'hbe383e9a, 32'h3e8fd540} /* (19, 8, 3) {real, imag} */,
  {32'hbf882f95, 32'hbf0ed096} /* (19, 8, 2) {real, imag} */,
  {32'h3f0e2444, 32'h3f8255e2} /* (19, 8, 1) {real, imag} */,
  {32'h3f375556, 32'h3f05c36d} /* (19, 8, 0) {real, imag} */,
  {32'hbf6b5acd, 32'hbf01bdf6} /* (19, 7, 31) {real, imag} */,
  {32'h3dcfc71f, 32'h3da4536e} /* (19, 7, 30) {real, imag} */,
  {32'hbe9991c4, 32'hbcc21b70} /* (19, 7, 29) {real, imag} */,
  {32'h3e36d0a4, 32'h3e93d83a} /* (19, 7, 28) {real, imag} */,
  {32'h3f374788, 32'h3ef3e716} /* (19, 7, 27) {real, imag} */,
  {32'hbe82eae2, 32'hbf310672} /* (19, 7, 26) {real, imag} */,
  {32'hbe8228bb, 32'hbdd179f6} /* (19, 7, 25) {real, imag} */,
  {32'h3dad9db2, 32'hbea85522} /* (19, 7, 24) {real, imag} */,
  {32'h3bac7680, 32'h3f603940} /* (19, 7, 23) {real, imag} */,
  {32'h3e101794, 32'h3d020dd0} /* (19, 7, 22) {real, imag} */,
  {32'h3ebb2285, 32'h3d364ee0} /* (19, 7, 21) {real, imag} */,
  {32'hbdcd48fc, 32'h3e91f961} /* (19, 7, 20) {real, imag} */,
  {32'h3be06de0, 32'hbe4839f4} /* (19, 7, 19) {real, imag} */,
  {32'h3db6562e, 32'hbe6e3590} /* (19, 7, 18) {real, imag} */,
  {32'h3e542d9d, 32'h3e650067} /* (19, 7, 17) {real, imag} */,
  {32'h3e8e8ce2, 32'hbed90632} /* (19, 7, 16) {real, imag} */,
  {32'hbdbe668a, 32'h3eb0bbc6} /* (19, 7, 15) {real, imag} */,
  {32'hbd928e4e, 32'hbe491ca8} /* (19, 7, 14) {real, imag} */,
  {32'h3ec57595, 32'h3e59b97a} /* (19, 7, 13) {real, imag} */,
  {32'hbd02c1f8, 32'h3ce0e020} /* (19, 7, 12) {real, imag} */,
  {32'hbe32ef24, 32'h3dcecb51} /* (19, 7, 11) {real, imag} */,
  {32'hbeab28ca, 32'hbe1dd2fa} /* (19, 7, 10) {real, imag} */,
  {32'h3ecaccc2, 32'hbe085364} /* (19, 7, 9) {real, imag} */,
  {32'hbd10fbc0, 32'h3e6ac096} /* (19, 7, 8) {real, imag} */,
  {32'hbf363d96, 32'h3da78ce7} /* (19, 7, 7) {real, imag} */,
  {32'h3ea3b9dc, 32'hbea3cba5} /* (19, 7, 6) {real, imag} */,
  {32'h3daa3790, 32'hbdba3962} /* (19, 7, 5) {real, imag} */,
  {32'h3e89e116, 32'hbdf3b504} /* (19, 7, 4) {real, imag} */,
  {32'h3f24558c, 32'h3e8649d7} /* (19, 7, 3) {real, imag} */,
  {32'h3eae4796, 32'h3c69cb20} /* (19, 7, 2) {real, imag} */,
  {32'hb9de3400, 32'hbf3658aa} /* (19, 7, 1) {real, imag} */,
  {32'hbc7b8bd0, 32'hbf5d3b81} /* (19, 7, 0) {real, imag} */,
  {32'hbe7efcf3, 32'hbda4e73e} /* (19, 6, 31) {real, imag} */,
  {32'hbe72464c, 32'h3da2b9f8} /* (19, 6, 30) {real, imag} */,
  {32'hbf35c7ff, 32'h3e5e49fc} /* (19, 6, 29) {real, imag} */,
  {32'h3e6eb21e, 32'h3e9007f9} /* (19, 6, 28) {real, imag} */,
  {32'hbe905c0d, 32'hbe8a4c61} /* (19, 6, 27) {real, imag} */,
  {32'hbde91fc0, 32'hbe70c93a} /* (19, 6, 26) {real, imag} */,
  {32'hbe3d4447, 32'hbdb92c38} /* (19, 6, 25) {real, imag} */,
  {32'hbefeb02c, 32'hbf2d7a0a} /* (19, 6, 24) {real, imag} */,
  {32'hbe04bc76, 32'h3ecf28f3} /* (19, 6, 23) {real, imag} */,
  {32'h3f5c604b, 32'h3de37ecc} /* (19, 6, 22) {real, imag} */,
  {32'hbe38b133, 32'h3e0e468d} /* (19, 6, 21) {real, imag} */,
  {32'hbd24e76d, 32'hbdfb9ce0} /* (19, 6, 20) {real, imag} */,
  {32'h3e1c54c4, 32'h3d06321c} /* (19, 6, 19) {real, imag} */,
  {32'hbecdbfe4, 32'hbf0c723a} /* (19, 6, 18) {real, imag} */,
  {32'hbd5dfaa6, 32'hbe888d8c} /* (19, 6, 17) {real, imag} */,
  {32'hbd63e088, 32'h3d6bac5c} /* (19, 6, 16) {real, imag} */,
  {32'hbe708ee4, 32'h3edaa2e1} /* (19, 6, 15) {real, imag} */,
  {32'h3e3cbb34, 32'hbf50c56e} /* (19, 6, 14) {real, imag} */,
  {32'h3de6c008, 32'h3e676597} /* (19, 6, 13) {real, imag} */,
  {32'h3ddaf764, 32'h3b2dd860} /* (19, 6, 12) {real, imag} */,
  {32'hbd63397c, 32'h3e12e3d2} /* (19, 6, 11) {real, imag} */,
  {32'h3e752360, 32'hbe00ff0c} /* (19, 6, 10) {real, imag} */,
  {32'hbf837597, 32'hbe1db860} /* (19, 6, 9) {real, imag} */,
  {32'hbf071d73, 32'h3f3f1688} /* (19, 6, 8) {real, imag} */,
  {32'h3dbf0f70, 32'h3c9d3310} /* (19, 6, 7) {real, imag} */,
  {32'h3f74b90e, 32'hbe9c5459} /* (19, 6, 6) {real, imag} */,
  {32'hbef2708c, 32'hbf06b3a2} /* (19, 6, 5) {real, imag} */,
  {32'hbe59d17a, 32'h3f5601fe} /* (19, 6, 4) {real, imag} */,
  {32'h3f609a3d, 32'hbf0d7073} /* (19, 6, 3) {real, imag} */,
  {32'hbe882679, 32'hbec602e8} /* (19, 6, 2) {real, imag} */,
  {32'hbea0fc08, 32'hbcc87840} /* (19, 6, 1) {real, imag} */,
  {32'hbdb0cfbc, 32'h3ec8823a} /* (19, 6, 0) {real, imag} */,
  {32'h40527f34, 32'hbebbb466} /* (19, 5, 31) {real, imag} */,
  {32'hbfc5716e, 32'h3e5b76a2} /* (19, 5, 30) {real, imag} */,
  {32'h3f0f7300, 32'h3f872e5d} /* (19, 5, 29) {real, imag} */,
  {32'hbf0d3c62, 32'hbe11bd70} /* (19, 5, 28) {real, imag} */,
  {32'hbed45832, 32'hbe961d6b} /* (19, 5, 27) {real, imag} */,
  {32'h3e5cde93, 32'h3f01fbd1} /* (19, 5, 26) {real, imag} */,
  {32'h3e90cc68, 32'h3e9f1b4e} /* (19, 5, 25) {real, imag} */,
  {32'hbeb3fd88, 32'hbf108162} /* (19, 5, 24) {real, imag} */,
  {32'hbe0496bc, 32'h3edfb443} /* (19, 5, 23) {real, imag} */,
  {32'h3d035870, 32'h3f0c5db3} /* (19, 5, 22) {real, imag} */,
  {32'hbe4e5fbe, 32'h3e94128f} /* (19, 5, 21) {real, imag} */,
  {32'hbe65bf52, 32'hbccf7918} /* (19, 5, 20) {real, imag} */,
  {32'hbe46b7c4, 32'h3dc8c093} /* (19, 5, 19) {real, imag} */,
  {32'h3e96676a, 32'h3ef33c61} /* (19, 5, 18) {real, imag} */,
  {32'h3f1c751e, 32'h3e129ff2} /* (19, 5, 17) {real, imag} */,
  {32'hbe00d748, 32'h3e9e8bc0} /* (19, 5, 16) {real, imag} */,
  {32'h3e8973a9, 32'hbe4c8f5a} /* (19, 5, 15) {real, imag} */,
  {32'hba0b9d60, 32'hbe288c9d} /* (19, 5, 14) {real, imag} */,
  {32'hbdcea606, 32'h3b62ff40} /* (19, 5, 13) {real, imag} */,
  {32'h3ed87bc4, 32'h3da61588} /* (19, 5, 12) {real, imag} */,
  {32'h3e465874, 32'hbe3832c1} /* (19, 5, 11) {real, imag} */,
  {32'hbe8855ff, 32'h3eeb3dec} /* (19, 5, 10) {real, imag} */,
  {32'hbe353ed3, 32'h3f1724c7} /* (19, 5, 9) {real, imag} */,
  {32'hbe88b8a8, 32'hbe139f89} /* (19, 5, 8) {real, imag} */,
  {32'h3fab8570, 32'hbe0b872d} /* (19, 5, 7) {real, imag} */,
  {32'hbe1c9743, 32'hbf16bcec} /* (19, 5, 6) {real, imag} */,
  {32'hbfa977b9, 32'h3de36958} /* (19, 5, 5) {real, imag} */,
  {32'h3f38956d, 32'h3dfae328} /* (19, 5, 4) {real, imag} */,
  {32'h3e411250, 32'h3e31ee9b} /* (19, 5, 3) {real, imag} */,
  {32'hbf9a71aa, 32'hbf98a112} /* (19, 5, 2) {real, imag} */,
  {32'h40026cc2, 32'h401ceb15} /* (19, 5, 1) {real, imag} */,
  {32'h3fb35bde, 32'h3fa6520e} /* (19, 5, 0) {real, imag} */,
  {32'hbfa6b5c0, 32'hc06efdb4} /* (19, 4, 31) {real, imag} */,
  {32'h3fedd8de, 32'h3feca51b} /* (19, 4, 30) {real, imag} */,
  {32'hbf0e63e5, 32'hbdc84d1e} /* (19, 4, 29) {real, imag} */,
  {32'hbfacd552, 32'hbeb024ae} /* (19, 4, 28) {real, imag} */,
  {32'h3fc071c9, 32'hbf806161} /* (19, 4, 27) {real, imag} */,
  {32'hbf94282e, 32'hbf183514} /* (19, 4, 26) {real, imag} */,
  {32'h3e84e112, 32'h3f24b92a} /* (19, 4, 25) {real, imag} */,
  {32'h3f049765, 32'hbdaf96cc} /* (19, 4, 24) {real, imag} */,
  {32'h3cbb57d0, 32'h3df7d6aa} /* (19, 4, 23) {real, imag} */,
  {32'hbc955dc4, 32'h3d06a6a4} /* (19, 4, 22) {real, imag} */,
  {32'h3f1d38f9, 32'h3d8b214c} /* (19, 4, 21) {real, imag} */,
  {32'hbf2636ce, 32'hbe85043f} /* (19, 4, 20) {real, imag} */,
  {32'hbe572b2e, 32'hbf538093} /* (19, 4, 19) {real, imag} */,
  {32'hbea641d6, 32'hbc67a820} /* (19, 4, 18) {real, imag} */,
  {32'h3dc861d9, 32'hbe332eac} /* (19, 4, 17) {real, imag} */,
  {32'hbe92da76, 32'h3d9e26ea} /* (19, 4, 16) {real, imag} */,
  {32'hbd0834a0, 32'hbee555d2} /* (19, 4, 15) {real, imag} */,
  {32'hbe4b3354, 32'h3edff7bb} /* (19, 4, 14) {real, imag} */,
  {32'h3f034280, 32'h3de0beea} /* (19, 4, 13) {real, imag} */,
  {32'hbdc1d393, 32'hbcc1d5e0} /* (19, 4, 12) {real, imag} */,
  {32'hbeb31862, 32'h3e7c18d2} /* (19, 4, 11) {real, imag} */,
  {32'hbea6453a, 32'h3b74a2c0} /* (19, 4, 10) {real, imag} */,
  {32'h3bf547a0, 32'hbebf77df} /* (19, 4, 9) {real, imag} */,
  {32'h3e0a7c58, 32'h3e957658} /* (19, 4, 8) {real, imag} */,
  {32'hbe4d0f69, 32'hbdd2922e} /* (19, 4, 7) {real, imag} */,
  {32'hbe93bf44, 32'h3e63ede6} /* (19, 4, 6) {real, imag} */,
  {32'hbd70d1aa, 32'h3f6b6441} /* (19, 4, 5) {real, imag} */,
  {32'h3ed42306, 32'hbed5c51a} /* (19, 4, 4) {real, imag} */,
  {32'hbf8c1000, 32'hbf5e74b8} /* (19, 4, 3) {real, imag} */,
  {32'h405b3682, 32'h400b5a9b} /* (19, 4, 2) {real, imag} */,
  {32'hc0a0ee6b, 32'hc015057c} /* (19, 4, 1) {real, imag} */,
  {32'hc0119f9c, 32'hbf271882} /* (19, 4, 0) {real, imag} */,
  {32'h406d1552, 32'hc07f18b3} /* (19, 3, 31) {real, imag} */,
  {32'hc00324c7, 32'h40c0b34e} /* (19, 3, 30) {real, imag} */,
  {32'hbf8c2a7e, 32'hbe4bd342} /* (19, 3, 29) {real, imag} */,
  {32'hbf373c64, 32'hbeba94d5} /* (19, 3, 28) {real, imag} */,
  {32'hbde4b90c, 32'hbf643918} /* (19, 3, 27) {real, imag} */,
  {32'h3e847d8a, 32'hbe5f2cc2} /* (19, 3, 26) {real, imag} */,
  {32'hbf302a8e, 32'h3f7556e4} /* (19, 3, 25) {real, imag} */,
  {32'h3eb4f57c, 32'hbd076960} /* (19, 3, 24) {real, imag} */,
  {32'h3e31fb91, 32'h3ef89852} /* (19, 3, 23) {real, imag} */,
  {32'hbf8aa34c, 32'hbf54624a} /* (19, 3, 22) {real, imag} */,
  {32'h3e16ccc1, 32'hbd463cec} /* (19, 3, 21) {real, imag} */,
  {32'h3e9ec64f, 32'hbede5611} /* (19, 3, 20) {real, imag} */,
  {32'hbe9ef57c, 32'h3f12f3f4} /* (19, 3, 19) {real, imag} */,
  {32'h3f055cd6, 32'hbe63d4e6} /* (19, 3, 18) {real, imag} */,
  {32'h3dcb5068, 32'h3e2c92ba} /* (19, 3, 17) {real, imag} */,
  {32'hbdad0c22, 32'hbe1b5293} /* (19, 3, 16) {real, imag} */,
  {32'hbe9571a9, 32'hbde2bc94} /* (19, 3, 15) {real, imag} */,
  {32'hbe872c9f, 32'h3e0b7e99} /* (19, 3, 14) {real, imag} */,
  {32'hbe77d880, 32'h3e7becfa} /* (19, 3, 13) {real, imag} */,
  {32'h3f27e896, 32'hbd1a2588} /* (19, 3, 12) {real, imag} */,
  {32'hbef4f227, 32'hbe99d71f} /* (19, 3, 11) {real, imag} */,
  {32'h3e9baff1, 32'h3ea13286} /* (19, 3, 10) {real, imag} */,
  {32'h3e835da2, 32'hbf1bf923} /* (19, 3, 9) {real, imag} */,
  {32'h3d3f5a18, 32'h3e537ff8} /* (19, 3, 8) {real, imag} */,
  {32'hbf010248, 32'hbe27daac} /* (19, 3, 7) {real, imag} */,
  {32'h3ec32411, 32'hbd22c94e} /* (19, 3, 6) {real, imag} */,
  {32'hbee6997b, 32'h3c8d14a0} /* (19, 3, 5) {real, imag} */,
  {32'h3f703abd, 32'h3e81f997} /* (19, 3, 4) {real, imag} */,
  {32'h3f9b4812, 32'hbe3d9077} /* (19, 3, 3) {real, imag} */,
  {32'h4010e6d0, 32'h40844652} /* (19, 3, 2) {real, imag} */,
  {32'hc0787158, 32'hc07fa6a3} /* (19, 3, 1) {real, imag} */,
  {32'hbf2a1f56, 32'h3f92d83e} /* (19, 3, 0) {real, imag} */,
  {32'h42183966, 32'hbf6e873e} /* (19, 2, 31) {real, imag} */,
  {32'hc1a00bf6, 32'h409783a5} /* (19, 2, 30) {real, imag} */,
  {32'h3fe4ebc4, 32'h3e9d3bea} /* (19, 2, 29) {real, imag} */,
  {32'h401139d3, 32'hc025bd74} /* (19, 2, 28) {real, imag} */,
  {32'hbf9d8382, 32'h3e9546e2} /* (19, 2, 27) {real, imag} */,
  {32'hbe87fc44, 32'h3ef5a83e} /* (19, 2, 26) {real, imag} */,
  {32'h3ed43815, 32'hbf931c38} /* (19, 2, 25) {real, imag} */,
  {32'hbdce87c0, 32'h3f66da45} /* (19, 2, 24) {real, imag} */,
  {32'hbea4df02, 32'hbf13f618} /* (19, 2, 23) {real, imag} */,
  {32'h3cf39674, 32'hbe8c3be0} /* (19, 2, 22) {real, imag} */,
  {32'hbf3cb7f9, 32'h3f504bce} /* (19, 2, 21) {real, imag} */,
  {32'h3ecf24ed, 32'hbe9fc726} /* (19, 2, 20) {real, imag} */,
  {32'hbe9aa231, 32'h3d71d848} /* (19, 2, 19) {real, imag} */,
  {32'h3e5bca44, 32'h3cf3fe7c} /* (19, 2, 18) {real, imag} */,
  {32'h3c4cef60, 32'hbebb548b} /* (19, 2, 17) {real, imag} */,
  {32'h3e90cbfe, 32'h3cd516bc} /* (19, 2, 16) {real, imag} */,
  {32'h3d3426c4, 32'h3d16e272} /* (19, 2, 15) {real, imag} */,
  {32'h3de14566, 32'hbe325b9e} /* (19, 2, 14) {real, imag} */,
  {32'h3d138489, 32'h3ebd4e69} /* (19, 2, 13) {real, imag} */,
  {32'hbeb4704e, 32'h3cfe7e2c} /* (19, 2, 12) {real, imag} */,
  {32'hbed3d6a8, 32'hbf4e17d4} /* (19, 2, 11) {real, imag} */,
  {32'hbd66ad3e, 32'h3e8125ef} /* (19, 2, 10) {real, imag} */,
  {32'h3e8f7533, 32'h3eab22eb} /* (19, 2, 9) {real, imag} */,
  {32'hbe486bd4, 32'hbfc4d424} /* (19, 2, 8) {real, imag} */,
  {32'h3e6cdc44, 32'hbebb3f66} /* (19, 2, 7) {real, imag} */,
  {32'h3e82c26a, 32'hbdb9af58} /* (19, 2, 6) {real, imag} */,
  {32'hc017ab95, 32'hc022e8c7} /* (19, 2, 5) {real, imag} */,
  {32'h4068a60e, 32'hbe8d23c2} /* (19, 2, 4) {real, imag} */,
  {32'h3f146dcd, 32'h3f250ed3} /* (19, 2, 3) {real, imag} */,
  {32'hc15a912f, 32'h406f188a} /* (19, 2, 2) {real, imag} */,
  {32'h41b41a12, 32'hc08a4c11} /* (19, 2, 1) {real, imag} */,
  {32'h41a2870c, 32'h40527fe6} /* (19, 2, 0) {real, imag} */,
  {32'hc24755b8, 32'h414ef1e9} /* (19, 1, 31) {real, imag} */,
  {32'h41545f5f, 32'h3f22f934} /* (19, 1, 30) {real, imag} */,
  {32'hbf21674d, 32'hbfae63c3} /* (19, 1, 29) {real, imag} */,
  {32'hc0189234, 32'hc0196fae} /* (19, 1, 28) {real, imag} */,
  {32'h4078108b, 32'h3f12529f} /* (19, 1, 27) {real, imag} */,
  {32'h3f615250, 32'hbf90711c} /* (19, 1, 26) {real, imag} */,
  {32'hbec2ad45, 32'h3f763974} /* (19, 1, 25) {real, imag} */,
  {32'h3dac82e0, 32'hbede57fb} /* (19, 1, 24) {real, imag} */,
  {32'h3f4fccd1, 32'hbe6a1754} /* (19, 1, 23) {real, imag} */,
  {32'h3e27127e, 32'h3ea95a08} /* (19, 1, 22) {real, imag} */,
  {32'h3eaaef27, 32'hbf498c38} /* (19, 1, 21) {real, imag} */,
  {32'hbd1cf1f2, 32'h3e9e022b} /* (19, 1, 20) {real, imag} */,
  {32'h3eb263bc, 32'h3d6b920c} /* (19, 1, 19) {real, imag} */,
  {32'h3eb7e1e0, 32'hbf33eae0} /* (19, 1, 18) {real, imag} */,
  {32'hbe7e3945, 32'h3d2f1cfc} /* (19, 1, 17) {real, imag} */,
  {32'hbdd52879, 32'hba011980} /* (19, 1, 16) {real, imag} */,
  {32'h3e48eaea, 32'hbd7c2fa4} /* (19, 1, 15) {real, imag} */,
  {32'hbe099036, 32'h3ecc92ce} /* (19, 1, 14) {real, imag} */,
  {32'hbd6172eb, 32'h3debe5f8} /* (19, 1, 13) {real, imag} */,
  {32'hbdfa8334, 32'h3e0d6764} /* (19, 1, 12) {real, imag} */,
  {32'h3f46c586, 32'h3edba026} /* (19, 1, 11) {real, imag} */,
  {32'h3f07e204, 32'h3d271c4a} /* (19, 1, 10) {real, imag} */,
  {32'hbf6a3b3f, 32'h3d3a1744} /* (19, 1, 9) {real, imag} */,
  {32'h3f38fbac, 32'h3f2399dc} /* (19, 1, 8) {real, imag} */,
  {32'hbefe6a95, 32'hbe1779ab} /* (19, 1, 7) {real, imag} */,
  {32'h3e8db760, 32'h3db9a8d8} /* (19, 1, 6) {real, imag} */,
  {32'h3fdc707a, 32'h3f974044} /* (19, 1, 5) {real, imag} */,
  {32'hbfdac26a, 32'hbff89b00} /* (19, 1, 4) {real, imag} */,
  {32'h3fa7ab86, 32'hbc7ca780} /* (19, 1, 3) {real, imag} */,
  {32'h418653f0, 32'h41949d4d} /* (19, 1, 2) {real, imag} */,
  {32'hc28d96c0, 32'hc2126cb8} /* (19, 1, 1) {real, imag} */,
  {32'hc2706f6a, 32'hc11e44bc} /* (19, 1, 0) {real, imag} */,
  {32'hc234955a, 32'h42071047} /* (19, 0, 31) {real, imag} */,
  {32'h40a469c7, 32'hc11d60a3} /* (19, 0, 30) {real, imag} */,
  {32'hbecb3016, 32'hbf9247de} /* (19, 0, 29) {real, imag} */,
  {32'hbeb92829, 32'hbf82596a} /* (19, 0, 28) {real, imag} */,
  {32'h3fe7ff0e, 32'h3f686c4d} /* (19, 0, 27) {real, imag} */,
  {32'h3eec0766, 32'hbf3951c8} /* (19, 0, 26) {real, imag} */,
  {32'hbeace883, 32'h3e6f5ebe} /* (19, 0, 25) {real, imag} */,
  {32'h3e1f3d16, 32'hbf16d38e} /* (19, 0, 24) {real, imag} */,
  {32'h3f854f34, 32'hbee7621a} /* (19, 0, 23) {real, imag} */,
  {32'hbe45dd6c, 32'hbec1b8fc} /* (19, 0, 22) {real, imag} */,
  {32'h3e08e23c, 32'hbe0f130f} /* (19, 0, 21) {real, imag} */,
  {32'h3e0a0bc8, 32'h3d713f6e} /* (19, 0, 20) {real, imag} */,
  {32'h3ec35fa0, 32'h3dbf9ba4} /* (19, 0, 19) {real, imag} */,
  {32'h3ea5f34e, 32'hbdf3fffa} /* (19, 0, 18) {real, imag} */,
  {32'hbd4fa002, 32'hbd7072d8} /* (19, 0, 17) {real, imag} */,
  {32'h3f54992e, 32'h00000000} /* (19, 0, 16) {real, imag} */,
  {32'hbd4fa002, 32'h3d7072d8} /* (19, 0, 15) {real, imag} */,
  {32'h3ea5f34e, 32'h3df3fffa} /* (19, 0, 14) {real, imag} */,
  {32'h3ec35fa0, 32'hbdbf9ba4} /* (19, 0, 13) {real, imag} */,
  {32'h3e0a0bc8, 32'hbd713f6e} /* (19, 0, 12) {real, imag} */,
  {32'h3e08e23c, 32'h3e0f130f} /* (19, 0, 11) {real, imag} */,
  {32'hbe45dd6c, 32'h3ec1b8fc} /* (19, 0, 10) {real, imag} */,
  {32'h3f854f34, 32'h3ee7621a} /* (19, 0, 9) {real, imag} */,
  {32'h3e1f3d16, 32'h3f16d38e} /* (19, 0, 8) {real, imag} */,
  {32'hbeace883, 32'hbe6f5ebe} /* (19, 0, 7) {real, imag} */,
  {32'h3eec0766, 32'h3f3951c8} /* (19, 0, 6) {real, imag} */,
  {32'h3fe7ff0e, 32'hbf686c4d} /* (19, 0, 5) {real, imag} */,
  {32'hbeb92829, 32'h3f82596a} /* (19, 0, 4) {real, imag} */,
  {32'hbecb3016, 32'h3f9247de} /* (19, 0, 3) {real, imag} */,
  {32'h40a469c7, 32'h411d60a3} /* (19, 0, 2) {real, imag} */,
  {32'hc234955a, 32'hc2071047} /* (19, 0, 1) {real, imag} */,
  {32'hc282a720, 32'h00000000} /* (19, 0, 0) {real, imag} */,
  {32'hc26e823b, 32'h41f00eda} /* (18, 31, 31) {real, imag} */,
  {32'h416a29e0, 32'hc1866126} /* (18, 31, 30) {real, imag} */,
  {32'hbe802ec0, 32'h3fb26612} /* (18, 31, 29) {real, imag} */,
  {32'hc00ec0fb, 32'h3f73042b} /* (18, 31, 28) {real, imag} */,
  {32'h3ff0565c, 32'hbfa6304d} /* (18, 31, 27) {real, imag} */,
  {32'h3ebd99f9, 32'h3ebb9e74} /* (18, 31, 26) {real, imag} */,
  {32'h3e933642, 32'h3ebe826c} /* (18, 31, 25) {real, imag} */,
  {32'h3f559114, 32'hbfa5812a} /* (18, 31, 24) {real, imag} */,
  {32'h3d77aa80, 32'hbda0195d} /* (18, 31, 23) {real, imag} */,
  {32'hbdcc2398, 32'hbeac2ff1} /* (18, 31, 22) {real, imag} */,
  {32'hbe46b422, 32'hbef97b76} /* (18, 31, 21) {real, imag} */,
  {32'h3efd21e6, 32'hbe2ad8a0} /* (18, 31, 20) {real, imag} */,
  {32'hbdcd6980, 32'hbdc2d80e} /* (18, 31, 19) {real, imag} */,
  {32'h3dd53931, 32'hbf2eca0a} /* (18, 31, 18) {real, imag} */,
  {32'hbea8bc65, 32'h3d9fcaa5} /* (18, 31, 17) {real, imag} */,
  {32'h3e99ee35, 32'hbcd78718} /* (18, 31, 16) {real, imag} */,
  {32'h3eb162c4, 32'hbdcf189d} /* (18, 31, 15) {real, imag} */,
  {32'h3e034555, 32'hbd9f2735} /* (18, 31, 14) {real, imag} */,
  {32'h3f011eda, 32'h3dafd45c} /* (18, 31, 13) {real, imag} */,
  {32'hbf63cc12, 32'hbe38bb6e} /* (18, 31, 12) {real, imag} */,
  {32'h3f5bea6d, 32'h3f3b826a} /* (18, 31, 11) {real, imag} */,
  {32'hbd58b9ca, 32'hbeb9152c} /* (18, 31, 10) {real, imag} */,
  {32'hbe06d7d4, 32'h3f651a0b} /* (18, 31, 9) {real, imag} */,
  {32'h3eeafe8a, 32'h3ef06d21} /* (18, 31, 8) {real, imag} */,
  {32'hbeb43e0d, 32'hbf7a1f54} /* (18, 31, 7) {real, imag} */,
  {32'h3fbf9e19, 32'h3f8297ce} /* (18, 31, 6) {real, imag} */,
  {32'h4074b350, 32'h3e988ef4} /* (18, 31, 5) {real, imag} */,
  {32'hc01c0b24, 32'h3fe34bbd} /* (18, 31, 4) {real, imag} */,
  {32'hbeabd25c, 32'hbdc813e0} /* (18, 31, 3) {real, imag} */,
  {32'h4130f2ea, 32'h3fc8d7d4} /* (18, 31, 2) {real, imag} */,
  {32'hc2259ac8, 32'hc116bdb0} /* (18, 31, 1) {real, imag} */,
  {32'hc24974b6, 32'h410889b4} /* (18, 31, 0) {real, imag} */,
  {32'h419ef118, 32'h40863630} /* (18, 30, 31) {real, imag} */,
  {32'hc13fb06a, 32'hc060251e} /* (18, 30, 30) {real, imag} */,
  {32'h3f9f44af, 32'hbf3e5dcc} /* (18, 30, 29) {real, imag} */,
  {32'h40476c6e, 32'h3f9b6e10} /* (18, 30, 28) {real, imag} */,
  {32'hbff9d368, 32'h402cbb2f} /* (18, 30, 27) {real, imag} */,
  {32'h3f33f47c, 32'hbf3c609f} /* (18, 30, 26) {real, imag} */,
  {32'h3f155588, 32'h3e82905a} /* (18, 30, 25) {real, imag} */,
  {32'hbec253be, 32'h3fa34232} /* (18, 30, 24) {real, imag} */,
  {32'h3f0eae98, 32'h3c34d750} /* (18, 30, 23) {real, imag} */,
  {32'hbdf8c564, 32'h3dfa6448} /* (18, 30, 22) {real, imag} */,
  {32'hbf1b09f2, 32'h3f421458} /* (18, 30, 21) {real, imag} */,
  {32'h3e52f316, 32'hbe818188} /* (18, 30, 20) {real, imag} */,
  {32'h3d30d500, 32'h3e6b0c05} /* (18, 30, 19) {real, imag} */,
  {32'hbdb61690, 32'h3dbc9606} /* (18, 30, 18) {real, imag} */,
  {32'h3e54502c, 32'h3e13f18a} /* (18, 30, 17) {real, imag} */,
  {32'hbd710c6a, 32'h3dd3ddd4} /* (18, 30, 16) {real, imag} */,
  {32'h3e62e486, 32'h3e087311} /* (18, 30, 15) {real, imag} */,
  {32'hbd96983f, 32'hbed174bd} /* (18, 30, 14) {real, imag} */,
  {32'hbe946b9f, 32'hbdbd1d20} /* (18, 30, 13) {real, imag} */,
  {32'h3d1b9b18, 32'h3e868819} /* (18, 30, 12) {real, imag} */,
  {32'hbda4dd75, 32'hbf32dc6b} /* (18, 30, 11) {real, imag} */,
  {32'hbd17b9c4, 32'hbe8d62d1} /* (18, 30, 10) {real, imag} */,
  {32'h3e0cdc66, 32'hbd4faa3c} /* (18, 30, 9) {real, imag} */,
  {32'hbee13b0a, 32'hbed8ef14} /* (18, 30, 8) {real, imag} */,
  {32'h3f21c464, 32'h3f023f05} /* (18, 30, 7) {real, imag} */,
  {32'hbeb30a2d, 32'hbece353d} /* (18, 30, 6) {real, imag} */,
  {32'hbfc9ea44, 32'hbf9c15e2} /* (18, 30, 5) {real, imag} */,
  {32'h40115d30, 32'h40201cde} /* (18, 30, 4) {real, imag} */,
  {32'h3f8b143d, 32'hbf7e5615} /* (18, 30, 3) {real, imag} */,
  {32'hc1875d3a, 32'hc0686d00} /* (18, 30, 2) {real, imag} */,
  {32'h4205513a, 32'h3ea712a0} /* (18, 30, 1) {real, imag} */,
  {32'h418dcf57, 32'hc0425e41} /* (18, 30, 0) {real, imag} */,
  {32'hc0348fa7, 32'h40a60828} /* (18, 29, 31) {real, imag} */,
  {32'h3fb20704, 32'hc041a831} /* (18, 29, 30) {real, imag} */,
  {32'h3f600ead, 32'h3fc026d7} /* (18, 29, 29) {real, imag} */,
  {32'h3f2ea328, 32'hbf83dfa6} /* (18, 29, 28) {real, imag} */,
  {32'hbdce3ad8, 32'hbd332a90} /* (18, 29, 27) {real, imag} */,
  {32'h3f07f5fd, 32'h3e599b5c} /* (18, 29, 26) {real, imag} */,
  {32'hbf1fffc0, 32'hbed67e7a} /* (18, 29, 25) {real, imag} */,
  {32'hbf1246d0, 32'h3f152422} /* (18, 29, 24) {real, imag} */,
  {32'h3eb13a2d, 32'h3d852554} /* (18, 29, 23) {real, imag} */,
  {32'h3f00f45e, 32'h3e574fba} /* (18, 29, 22) {real, imag} */,
  {32'hbe8973dc, 32'h3ddd9b4a} /* (18, 29, 21) {real, imag} */,
  {32'hbefe97ae, 32'hbd5f5a00} /* (18, 29, 20) {real, imag} */,
  {32'h3e49e798, 32'h3f0954a7} /* (18, 29, 19) {real, imag} */,
  {32'hbe7f1c46, 32'hbb1e5300} /* (18, 29, 18) {real, imag} */,
  {32'h3e2d0e2a, 32'hbde96407} /* (18, 29, 17) {real, imag} */,
  {32'hbdbbc42b, 32'h3db77460} /* (18, 29, 16) {real, imag} */,
  {32'h3d4abcba, 32'h3e8934a2} /* (18, 29, 15) {real, imag} */,
  {32'h3dc32a18, 32'hbe909a89} /* (18, 29, 14) {real, imag} */,
  {32'h3e9cdb5d, 32'h3b319480} /* (18, 29, 13) {real, imag} */,
  {32'hbdc8c2fe, 32'h3ed8738c} /* (18, 29, 12) {real, imag} */,
  {32'h3e225c72, 32'h3f3862d6} /* (18, 29, 11) {real, imag} */,
  {32'hbe1011e6, 32'h3f59080b} /* (18, 29, 10) {real, imag} */,
  {32'h3e3d12dc, 32'hbe177c17} /* (18, 29, 9) {real, imag} */,
  {32'h3f2a120c, 32'h3dd93a4e} /* (18, 29, 8) {real, imag} */,
  {32'hbe8b909a, 32'hbf0302ce} /* (18, 29, 7) {real, imag} */,
  {32'hbf2ac12a, 32'h3f158560} /* (18, 29, 6) {real, imag} */,
  {32'h3f51bb1e, 32'h3f970d95} /* (18, 29, 5) {real, imag} */,
  {32'hbf64befe, 32'h3c205de0} /* (18, 29, 4) {real, imag} */,
  {32'hbf8aa8e9, 32'hbee5ffcf} /* (18, 29, 3) {real, imag} */,
  {32'hbfee0f18, 32'hc0c74fde} /* (18, 29, 2) {real, imag} */,
  {32'h404a9d42, 32'h407edc80} /* (18, 29, 1) {real, imag} */,
  {32'hbcba5bc0, 32'h3e826d97} /* (18, 29, 0) {real, imag} */,
  {32'hc07fc6c7, 32'h3fb10953} /* (18, 28, 31) {real, imag} */,
  {32'h4057928a, 32'hbfe7c8c7} /* (18, 28, 30) {real, imag} */,
  {32'hbd9b8cb8, 32'h3f018fab} /* (18, 28, 29) {real, imag} */,
  {32'h3f18c316, 32'hbe065ea4} /* (18, 28, 28) {real, imag} */,
  {32'hbe91795a, 32'hbf63db25} /* (18, 28, 27) {real, imag} */,
  {32'hbe977314, 32'hbf9ae2a6} /* (18, 28, 26) {real, imag} */,
  {32'hbde2813a, 32'h3d8ff1f4} /* (18, 28, 25) {real, imag} */,
  {32'h3ea3e1be, 32'hbecf356b} /* (18, 28, 24) {real, imag} */,
  {32'h3e0f3ca8, 32'h3e5e4f87} /* (18, 28, 23) {real, imag} */,
  {32'h3f19d7af, 32'h3f10b966} /* (18, 28, 22) {real, imag} */,
  {32'h3eac9bbe, 32'h3d3bda16} /* (18, 28, 21) {real, imag} */,
  {32'h3def3f67, 32'h3f231d7a} /* (18, 28, 20) {real, imag} */,
  {32'hbde1f4be, 32'hbec34b59} /* (18, 28, 19) {real, imag} */,
  {32'h3d881b3e, 32'hbd30f1d0} /* (18, 28, 18) {real, imag} */,
  {32'h3e370e60, 32'h3d3275e0} /* (18, 28, 17) {real, imag} */,
  {32'hbeb37658, 32'h3e2d2a68} /* (18, 28, 16) {real, imag} */,
  {32'hbe015f50, 32'h3d6c8440} /* (18, 28, 15) {real, imag} */,
  {32'hbe43cd48, 32'h3eac2125} /* (18, 28, 14) {real, imag} */,
  {32'hbcc49070, 32'hbebd046b} /* (18, 28, 13) {real, imag} */,
  {32'h3edac598, 32'hbd00cf73} /* (18, 28, 12) {real, imag} */,
  {32'h3bacb390, 32'h3e63109e} /* (18, 28, 11) {real, imag} */,
  {32'hbea4f1a0, 32'hbf0bb399} /* (18, 28, 10) {real, imag} */,
  {32'hbe5f0bd2, 32'hbe670ad4} /* (18, 28, 9) {real, imag} */,
  {32'h3df4bd7e, 32'h3c648ba8} /* (18, 28, 8) {real, imag} */,
  {32'hbe06c778, 32'hbeaa01ba} /* (18, 28, 7) {real, imag} */,
  {32'hbe5c34f6, 32'hbe88da1c} /* (18, 28, 6) {real, imag} */,
  {32'h3f3aaf6e, 32'h3f1bf6e0} /* (18, 28, 5) {real, imag} */,
  {32'hbfecaaf3, 32'h3f4335ad} /* (18, 28, 4) {real, imag} */,
  {32'h3db908ea, 32'h3e5ff103} /* (18, 28, 3) {real, imag} */,
  {32'h3f05754b, 32'hbfe609b9} /* (18, 28, 2) {real, imag} */,
  {32'hbfc84ff7, 32'h4083b242} /* (18, 28, 1) {real, imag} */,
  {32'hc0018090, 32'h3f49ca12} /* (18, 28, 0) {real, imag} */,
  {32'h3fe81686, 32'hc010e72e} /* (18, 27, 31) {real, imag} */,
  {32'hbf4e6b93, 32'h3fb8f374} /* (18, 27, 30) {real, imag} */,
  {32'hbdad2e56, 32'hbe7e8db4} /* (18, 27, 29) {real, imag} */,
  {32'hbdf25112, 32'hbf0b0a0d} /* (18, 27, 28) {real, imag} */,
  {32'hbf585a34, 32'hbe9973f2} /* (18, 27, 27) {real, imag} */,
  {32'hbf2a97f4, 32'h3e922791} /* (18, 27, 26) {real, imag} */,
  {32'h3f951339, 32'hbe836c77} /* (18, 27, 25) {real, imag} */,
  {32'h3f226e57, 32'hbed79de6} /* (18, 27, 24) {real, imag} */,
  {32'h3b82aa08, 32'h3f3ec104} /* (18, 27, 23) {real, imag} */,
  {32'h3d91fe8f, 32'h3e23906a} /* (18, 27, 22) {real, imag} */,
  {32'hbe4a4efa, 32'h3f5c728b} /* (18, 27, 21) {real, imag} */,
  {32'h3bc0e900, 32'h3f0f6592} /* (18, 27, 20) {real, imag} */,
  {32'h3ed6e875, 32'hbe92d87e} /* (18, 27, 19) {real, imag} */,
  {32'h3e235792, 32'hbe692dcb} /* (18, 27, 18) {real, imag} */,
  {32'h3cab2268, 32'h3c72d4d0} /* (18, 27, 17) {real, imag} */,
  {32'h3e515a50, 32'h3de72d15} /* (18, 27, 16) {real, imag} */,
  {32'h3cbc89f6, 32'hbedf9d38} /* (18, 27, 15) {real, imag} */,
  {32'hbe2d566b, 32'hbf214a7d} /* (18, 27, 14) {real, imag} */,
  {32'hbd92765a, 32'h3cf4d978} /* (18, 27, 13) {real, imag} */,
  {32'hbeaf27a1, 32'h3dc9164c} /* (18, 27, 12) {real, imag} */,
  {32'hbef4a2a4, 32'h3e08ed37} /* (18, 27, 11) {real, imag} */,
  {32'h3e78e11f, 32'h3e3c4a4f} /* (18, 27, 10) {real, imag} */,
  {32'h3eb31538, 32'h3d342315} /* (18, 27, 9) {real, imag} */,
  {32'h3c926c1e, 32'h3f11838e} /* (18, 27, 8) {real, imag} */,
  {32'h3decad1c, 32'hbe9a1fc5} /* (18, 27, 7) {real, imag} */,
  {32'hbe2002d5, 32'hbee68fd7} /* (18, 27, 6) {real, imag} */,
  {32'h3dddbc1c, 32'hbe4b5269} /* (18, 27, 5) {real, imag} */,
  {32'hbe3acc79, 32'h3e8a7920} /* (18, 27, 4) {real, imag} */,
  {32'h3f0f9346, 32'h3db64c78} /* (18, 27, 3) {real, imag} */,
  {32'hbfbc1b42, 32'hbefefceb} /* (18, 27, 2) {real, imag} */,
  {32'h4029d441, 32'hbf686370} /* (18, 27, 1) {real, imag} */,
  {32'h3fa6e5e7, 32'hbfc1347b} /* (18, 27, 0) {real, imag} */,
  {32'h3de6e11c, 32'h3e7fd4f3} /* (18, 26, 31) {real, imag} */,
  {32'h3ea298d6, 32'hbebc2be4} /* (18, 26, 30) {real, imag} */,
  {32'h3e7251d8, 32'hbe921351} /* (18, 26, 29) {real, imag} */,
  {32'h3e0373e5, 32'hbd09fb8c} /* (18, 26, 28) {real, imag} */,
  {32'hbef02ad4, 32'hbe6f7bb1} /* (18, 26, 27) {real, imag} */,
  {32'h3e7ec143, 32'h3eb32e32} /* (18, 26, 26) {real, imag} */,
  {32'h3f3f3470, 32'hbe8dacb0} /* (18, 26, 25) {real, imag} */,
  {32'hbe9717f0, 32'h3c2e02a0} /* (18, 26, 24) {real, imag} */,
  {32'hbd82bc54, 32'hbe816721} /* (18, 26, 23) {real, imag} */,
  {32'hbe2b5943, 32'hbdacfa27} /* (18, 26, 22) {real, imag} */,
  {32'hbda43448, 32'h3f1c3c45} /* (18, 26, 21) {real, imag} */,
  {32'h3e9896b4, 32'hbe1ecee4} /* (18, 26, 20) {real, imag} */,
  {32'hbed4feee, 32'hbe33c034} /* (18, 26, 19) {real, imag} */,
  {32'h3dae67ae, 32'hbdaf15df} /* (18, 26, 18) {real, imag} */,
  {32'h3e18106e, 32'hbe7758b0} /* (18, 26, 17) {real, imag} */,
  {32'h3db8221c, 32'hbe4ca0a8} /* (18, 26, 16) {real, imag} */,
  {32'h3d95121b, 32'h3dbe7b92} /* (18, 26, 15) {real, imag} */,
  {32'hbd34dcfc, 32'hbe5702ce} /* (18, 26, 14) {real, imag} */,
  {32'h3e26c33e, 32'h3dbc9148} /* (18, 26, 13) {real, imag} */,
  {32'h3ea85615, 32'hbe15f74e} /* (18, 26, 12) {real, imag} */,
  {32'hbd5d5c6d, 32'h3e1d9944} /* (18, 26, 11) {real, imag} */,
  {32'h3e9a3e71, 32'hbe96a9f1} /* (18, 26, 10) {real, imag} */,
  {32'h3efc95d0, 32'h3e4ed53d} /* (18, 26, 9) {real, imag} */,
  {32'hbd8431c4, 32'hbd0d5e38} /* (18, 26, 8) {real, imag} */,
  {32'hbe27696a, 32'h3ec4d52e} /* (18, 26, 7) {real, imag} */,
  {32'h3cc52a8c, 32'h3e664c6c} /* (18, 26, 6) {real, imag} */,
  {32'hbf03ae76, 32'hbe162556} /* (18, 26, 5) {real, imag} */,
  {32'hbe8bdb60, 32'hbda2d910} /* (18, 26, 4) {real, imag} */,
  {32'hbf7947a8, 32'hbe1bfaea} /* (18, 26, 3) {real, imag} */,
  {32'hbec7e3fb, 32'h3f34bcdb} /* (18, 26, 2) {real, imag} */,
  {32'h3e968407, 32'h3e4a0da9} /* (18, 26, 1) {real, imag} */,
  {32'hbe1ea980, 32'h3e967201} /* (18, 26, 0) {real, imag} */,
  {32'hbe889c61, 32'h3edefa54} /* (18, 25, 31) {real, imag} */,
  {32'h3e99782c, 32'hbf4ac280} /* (18, 25, 30) {real, imag} */,
  {32'h3da74128, 32'hbdc0ae17} /* (18, 25, 29) {real, imag} */,
  {32'h3f015c3c, 32'hbf09f8f7} /* (18, 25, 28) {real, imag} */,
  {32'hbede64c0, 32'h3e90fce9} /* (18, 25, 27) {real, imag} */,
  {32'h3e894ff2, 32'hbdb37177} /* (18, 25, 26) {real, imag} */,
  {32'hbeff0cb9, 32'hbf032600} /* (18, 25, 25) {real, imag} */,
  {32'hbee6ffde, 32'h3f4397ce} /* (18, 25, 24) {real, imag} */,
  {32'hbf16f172, 32'hbe3d4130} /* (18, 25, 23) {real, imag} */,
  {32'hbedb5c64, 32'hbc2f7600} /* (18, 25, 22) {real, imag} */,
  {32'h3e2df2c6, 32'hbeafe1f8} /* (18, 25, 21) {real, imag} */,
  {32'h3e9c2a00, 32'hbd7769c0} /* (18, 25, 20) {real, imag} */,
  {32'hbe752dd1, 32'h3deb7948} /* (18, 25, 19) {real, imag} */,
  {32'h3c447380, 32'hbf124975} /* (18, 25, 18) {real, imag} */,
  {32'hbe0cf666, 32'h3e438f80} /* (18, 25, 17) {real, imag} */,
  {32'hbdeee27a, 32'hbd0887fc} /* (18, 25, 16) {real, imag} */,
  {32'hbdaf4798, 32'h3eb0e194} /* (18, 25, 15) {real, imag} */,
  {32'h3e9cc670, 32'hbee57840} /* (18, 25, 14) {real, imag} */,
  {32'hbee0bc04, 32'h3db54315} /* (18, 25, 13) {real, imag} */,
  {32'h3e76a654, 32'hbd7f5270} /* (18, 25, 12) {real, imag} */,
  {32'hbe461a6a, 32'hbeb12c68} /* (18, 25, 11) {real, imag} */,
  {32'hbed53b6e, 32'h3d4d63ab} /* (18, 25, 10) {real, imag} */,
  {32'h3ea69425, 32'hbedf2b09} /* (18, 25, 9) {real, imag} */,
  {32'hbd26c28c, 32'h3e2a817a} /* (18, 25, 8) {real, imag} */,
  {32'hbf2a3959, 32'h3f40d96e} /* (18, 25, 7) {real, imag} */,
  {32'h3eca1bd6, 32'h3eae77c7} /* (18, 25, 6) {real, imag} */,
  {32'h3f11ff38, 32'hbde129e4} /* (18, 25, 5) {real, imag} */,
  {32'h3ebce270, 32'hbe576006} /* (18, 25, 4) {real, imag} */,
  {32'hbe9937b0, 32'h3e65547d} /* (18, 25, 3) {real, imag} */,
  {32'h3f426626, 32'h3dd72550} /* (18, 25, 2) {real, imag} */,
  {32'hbe44742c, 32'h3f13fe1e} /* (18, 25, 1) {real, imag} */,
  {32'hbe865c86, 32'h3ee8a097} /* (18, 25, 0) {real, imag} */,
  {32'h3f24a274, 32'hbf3bd90e} /* (18, 24, 31) {real, imag} */,
  {32'hbf2e4f33, 32'h3f279fd2} /* (18, 24, 30) {real, imag} */,
  {32'hbda844fa, 32'hbd1fa0ba} /* (18, 24, 29) {real, imag} */,
  {32'h3e1db65a, 32'hbd9c4b41} /* (18, 24, 28) {real, imag} */,
  {32'h3d895815, 32'h3d382808} /* (18, 24, 27) {real, imag} */,
  {32'h3e723594, 32'h3e369b9d} /* (18, 24, 26) {real, imag} */,
  {32'hbca587d0, 32'h3ac17440} /* (18, 24, 25) {real, imag} */,
  {32'hbe67807a, 32'hbe817f57} /* (18, 24, 24) {real, imag} */,
  {32'h3e05f377, 32'h3e24cfda} /* (18, 24, 23) {real, imag} */,
  {32'h3e309488, 32'h3f19dc28} /* (18, 24, 22) {real, imag} */,
  {32'h3f0360e8, 32'hbd473e58} /* (18, 24, 21) {real, imag} */,
  {32'h3e88072e, 32'hbcdab0d0} /* (18, 24, 20) {real, imag} */,
  {32'hbeb787b9, 32'h3e7c9629} /* (18, 24, 19) {real, imag} */,
  {32'h3e06e7fa, 32'h3d7c4b12} /* (18, 24, 18) {real, imag} */,
  {32'hbded8e70, 32'hbca67500} /* (18, 24, 17) {real, imag} */,
  {32'hbe693a5a, 32'hbe00ea24} /* (18, 24, 16) {real, imag} */,
  {32'hbe3e9580, 32'h3e0e6074} /* (18, 24, 15) {real, imag} */,
  {32'h3e4aa6c5, 32'h3d9e00e6} /* (18, 24, 14) {real, imag} */,
  {32'h3f03e79c, 32'hbe04c6cd} /* (18, 24, 13) {real, imag} */,
  {32'h3e9f8ebc, 32'h3ebf807a} /* (18, 24, 12) {real, imag} */,
  {32'hbf02fa47, 32'hbe2c5295} /* (18, 24, 11) {real, imag} */,
  {32'hbf2bd018, 32'hbdadbc82} /* (18, 24, 10) {real, imag} */,
  {32'hbed357be, 32'hbebdadf3} /* (18, 24, 9) {real, imag} */,
  {32'hbdf0c720, 32'h3e8e75bc} /* (18, 24, 8) {real, imag} */,
  {32'h3ef4a263, 32'h3ea1575e} /* (18, 24, 7) {real, imag} */,
  {32'hbe428a4a, 32'h3e8ef21a} /* (18, 24, 6) {real, imag} */,
  {32'hbed8047c, 32'h3db3f9b5} /* (18, 24, 5) {real, imag} */,
  {32'h3e466a80, 32'hbf1a2a99} /* (18, 24, 4) {real, imag} */,
  {32'h3c8ac2b0, 32'h3e79037a} /* (18, 24, 3) {real, imag} */,
  {32'hbf9f0f48, 32'hbe0cdccf} /* (18, 24, 2) {real, imag} */,
  {32'h3fccb150, 32'hbf8c0d71} /* (18, 24, 1) {real, imag} */,
  {32'h3f0bae06, 32'hbf8b0557} /* (18, 24, 0) {real, imag} */,
  {32'hbd0c24c0, 32'h3ec2a79b} /* (18, 23, 31) {real, imag} */,
  {32'hbdbf16a6, 32'hbef7edee} /* (18, 23, 30) {real, imag} */,
  {32'hbe4cf12d, 32'hbdf65444} /* (18, 23, 29) {real, imag} */,
  {32'h3d873d34, 32'h3f53ee12} /* (18, 23, 28) {real, imag} */,
  {32'hbeb5dedb, 32'hbe2eca4a} /* (18, 23, 27) {real, imag} */,
  {32'h3e7ad470, 32'h3e67c5b1} /* (18, 23, 26) {real, imag} */,
  {32'hbea29d3d, 32'hbc807ea0} /* (18, 23, 25) {real, imag} */,
  {32'hbe70c392, 32'h3d5ada28} /* (18, 23, 24) {real, imag} */,
  {32'hbecf78c0, 32'h3f1289ae} /* (18, 23, 23) {real, imag} */,
  {32'h3cba56f8, 32'hbf28a20a} /* (18, 23, 22) {real, imag} */,
  {32'hbf623c80, 32'hbf1eb781} /* (18, 23, 21) {real, imag} */,
  {32'hbea57953, 32'h3e02c6f6} /* (18, 23, 20) {real, imag} */,
  {32'h3e147e26, 32'hbed8895c} /* (18, 23, 19) {real, imag} */,
  {32'hbe327778, 32'hbd821d5f} /* (18, 23, 18) {real, imag} */,
  {32'h3d2f3662, 32'hbe1891d4} /* (18, 23, 17) {real, imag} */,
  {32'h3ef09a9a, 32'h3e33cd96} /* (18, 23, 16) {real, imag} */,
  {32'h3e02275e, 32'hbf1f6ffe} /* (18, 23, 15) {real, imag} */,
  {32'h3e4d74d0, 32'h3ee29c12} /* (18, 23, 14) {real, imag} */,
  {32'hbe4e54b8, 32'h3e86b5ed} /* (18, 23, 13) {real, imag} */,
  {32'hbe60aa19, 32'hbefd1e83} /* (18, 23, 12) {real, imag} */,
  {32'h3eba3d79, 32'hbe4a3648} /* (18, 23, 11) {real, imag} */,
  {32'h3ee022a2, 32'h3f32e552} /* (18, 23, 10) {real, imag} */,
  {32'hbe5fe69c, 32'hbf2127d8} /* (18, 23, 9) {real, imag} */,
  {32'h3f07a1f6, 32'h3ea7810c} /* (18, 23, 8) {real, imag} */,
  {32'hbecea782, 32'hbf28d47c} /* (18, 23, 7) {real, imag} */,
  {32'hbe1638e5, 32'h3f170567} /* (18, 23, 6) {real, imag} */,
  {32'h3e2ed934, 32'h3edc8344} /* (18, 23, 5) {real, imag} */,
  {32'hbf068147, 32'h3eaa71f0} /* (18, 23, 4) {real, imag} */,
  {32'h3f0dcb36, 32'hbd9c2207} /* (18, 23, 3) {real, imag} */,
  {32'hbbe86ec0, 32'hbf9fe30a} /* (18, 23, 2) {real, imag} */,
  {32'h3e478cdb, 32'h3e5d63b0} /* (18, 23, 1) {real, imag} */,
  {32'h3e5b0059, 32'h3dc55da4} /* (18, 23, 0) {real, imag} */,
  {32'hbf115382, 32'h3eaa47fe} /* (18, 22, 31) {real, imag} */,
  {32'h3f023b0a, 32'hbf58cadc} /* (18, 22, 30) {real, imag} */,
  {32'hbf78cd7c, 32'h3e8b0f55} /* (18, 22, 29) {real, imag} */,
  {32'hbed135be, 32'h3f0c9a5a} /* (18, 22, 28) {real, imag} */,
  {32'hbedc4ef8, 32'hbea7c67e} /* (18, 22, 27) {real, imag} */,
  {32'hbf09c652, 32'h3ef0b666} /* (18, 22, 26) {real, imag} */,
  {32'hbc3373b0, 32'hbb8b2b70} /* (18, 22, 25) {real, imag} */,
  {32'h3d800aec, 32'hbde84340} /* (18, 22, 24) {real, imag} */,
  {32'hbe1a4fbf, 32'hbd0395a0} /* (18, 22, 23) {real, imag} */,
  {32'h3e09aa15, 32'hbef4da06} /* (18, 22, 22) {real, imag} */,
  {32'h3f04e3d5, 32'hbebafa88} /* (18, 22, 21) {real, imag} */,
  {32'h3e8fedc9, 32'h3dab1f58} /* (18, 22, 20) {real, imag} */,
  {32'hbed67cb2, 32'hbe0aca7a} /* (18, 22, 19) {real, imag} */,
  {32'h3e590ee0, 32'h3e894de2} /* (18, 22, 18) {real, imag} */,
  {32'hbe37933e, 32'h3ed0bcde} /* (18, 22, 17) {real, imag} */,
  {32'h3d151248, 32'hbdf41b0d} /* (18, 22, 16) {real, imag} */,
  {32'hbd8d049e, 32'h3e1d2cdc} /* (18, 22, 15) {real, imag} */,
  {32'hbd85bf93, 32'h3e97de0c} /* (18, 22, 14) {real, imag} */,
  {32'h3dcb12f6, 32'h3e79e3d5} /* (18, 22, 13) {real, imag} */,
  {32'hbd916647, 32'h3e718d64} /* (18, 22, 12) {real, imag} */,
  {32'hbe0763cf, 32'h3d914954} /* (18, 22, 11) {real, imag} */,
  {32'hbe1e4ee4, 32'h3f146131} /* (18, 22, 10) {real, imag} */,
  {32'hbe8687d9, 32'hbf281e12} /* (18, 22, 9) {real, imag} */,
  {32'hbe50b588, 32'h3d0f53dc} /* (18, 22, 8) {real, imag} */,
  {32'hbc7aac60, 32'h3d9c2600} /* (18, 22, 7) {real, imag} */,
  {32'h3d9aabf8, 32'hbd76384c} /* (18, 22, 6) {real, imag} */,
  {32'h3e271518, 32'hbdbddb87} /* (18, 22, 5) {real, imag} */,
  {32'hbd7ea7b0, 32'hbe09e608} /* (18, 22, 4) {real, imag} */,
  {32'hbe5a7cd1, 32'h3e99c3af} /* (18, 22, 3) {real, imag} */,
  {32'h3e62a9d2, 32'h3ed4acbc} /* (18, 22, 2) {real, imag} */,
  {32'h3d217b12, 32'hbaf9db00} /* (18, 22, 1) {real, imag} */,
  {32'h3f051758, 32'hbd10f790} /* (18, 22, 0) {real, imag} */,
  {32'hbcf75106, 32'hbf616006} /* (18, 21, 31) {real, imag} */,
  {32'h3d568bd0, 32'h3ec01b0b} /* (18, 21, 30) {real, imag} */,
  {32'hbef3c868, 32'hbf343d52} /* (18, 21, 29) {real, imag} */,
  {32'hbd4c9dab, 32'hbf0aad2d} /* (18, 21, 28) {real, imag} */,
  {32'h3de65f6a, 32'h3f54a1aa} /* (18, 21, 27) {real, imag} */,
  {32'h3e912699, 32'hbe8ea340} /* (18, 21, 26) {real, imag} */,
  {32'h3ea42938, 32'h3e5ce20e} /* (18, 21, 25) {real, imag} */,
  {32'h3f283fa8, 32'hbd30e27a} /* (18, 21, 24) {real, imag} */,
  {32'hbe38f910, 32'h3bcff0e0} /* (18, 21, 23) {real, imag} */,
  {32'h3e966274, 32'h3dc3d304} /* (18, 21, 22) {real, imag} */,
  {32'h3f383316, 32'h3e5a4636} /* (18, 21, 21) {real, imag} */,
  {32'hbef453a6, 32'h3e6b7c6a} /* (18, 21, 20) {real, imag} */,
  {32'hbe9898c2, 32'h3ea02b0a} /* (18, 21, 19) {real, imag} */,
  {32'h3db18192, 32'h3ec55b0f} /* (18, 21, 18) {real, imag} */,
  {32'hbf15541a, 32'hbeaa9232} /* (18, 21, 17) {real, imag} */,
  {32'hbe04fb12, 32'hbe7f6a4e} /* (18, 21, 16) {real, imag} */,
  {32'h3e177e5a, 32'h3db3235f} /* (18, 21, 15) {real, imag} */,
  {32'h3dc32bd9, 32'h3dc6f8c0} /* (18, 21, 14) {real, imag} */,
  {32'h3ec11eba, 32'h3dfc059d} /* (18, 21, 13) {real, imag} */,
  {32'h3ca4a95c, 32'h3ecb7288} /* (18, 21, 12) {real, imag} */,
  {32'hbe910e78, 32'h3e5f91bc} /* (18, 21, 11) {real, imag} */,
  {32'h3f175be4, 32'hbd84661f} /* (18, 21, 10) {real, imag} */,
  {32'hbec86ea6, 32'h3f1eb80c} /* (18, 21, 9) {real, imag} */,
  {32'hbe567d52, 32'h3eb5009c} /* (18, 21, 8) {real, imag} */,
  {32'h3f4eef9f, 32'h3e3fd62d} /* (18, 21, 7) {real, imag} */,
  {32'h3ee88b53, 32'hbeb5c210} /* (18, 21, 6) {real, imag} */,
  {32'h3e7dd55c, 32'hbcf30590} /* (18, 21, 5) {real, imag} */,
  {32'h3b3e9a60, 32'hbe2240e0} /* (18, 21, 4) {real, imag} */,
  {32'hbea242b6, 32'h3ee70ba4} /* (18, 21, 3) {real, imag} */,
  {32'hbee54173, 32'h3eb051e9} /* (18, 21, 2) {real, imag} */,
  {32'h3e27949a, 32'hbdb2d392} /* (18, 21, 1) {real, imag} */,
  {32'h3e920752, 32'hbedcedeb} /* (18, 21, 0) {real, imag} */,
  {32'hbdc71fb0, 32'hbeb29c2f} /* (18, 20, 31) {real, imag} */,
  {32'hbf1ab664, 32'hbd494cb4} /* (18, 20, 30) {real, imag} */,
  {32'hbe0ff586, 32'h3e8bad8c} /* (18, 20, 29) {real, imag} */,
  {32'h3d9091fa, 32'h3e22173d} /* (18, 20, 28) {real, imag} */,
  {32'h3de8e0ec, 32'hbc64886c} /* (18, 20, 27) {real, imag} */,
  {32'hbea62a54, 32'h3db508e0} /* (18, 20, 26) {real, imag} */,
  {32'hbe824209, 32'h3f2a681b} /* (18, 20, 25) {real, imag} */,
  {32'h3be5a7a0, 32'h3ed97184} /* (18, 20, 24) {real, imag} */,
  {32'hbe73b0b3, 32'hbe1bdef0} /* (18, 20, 23) {real, imag} */,
  {32'hbcbd1448, 32'hbdb7bd7e} /* (18, 20, 22) {real, imag} */,
  {32'hbe3d57c4, 32'hbd821a76} /* (18, 20, 21) {real, imag} */,
  {32'h3e8646c0, 32'hbef13927} /* (18, 20, 20) {real, imag} */,
  {32'h3c995ed2, 32'h3deb5256} /* (18, 20, 19) {real, imag} */,
  {32'hbecc83f8, 32'h3ea0a826} /* (18, 20, 18) {real, imag} */,
  {32'h3eb32505, 32'hbe1bcb72} /* (18, 20, 17) {real, imag} */,
  {32'hbe6976dd, 32'h3df85484} /* (18, 20, 16) {real, imag} */,
  {32'hbe54ca73, 32'h3de2dc40} /* (18, 20, 15) {real, imag} */,
  {32'h3e424968, 32'h3bed0740} /* (18, 20, 14) {real, imag} */,
  {32'hbec3d6e6, 32'h3e5ff217} /* (18, 20, 13) {real, imag} */,
  {32'h3f38c16e, 32'hbe0f9ed5} /* (18, 20, 12) {real, imag} */,
  {32'hbe9adb9e, 32'hbe99041b} /* (18, 20, 11) {real, imag} */,
  {32'hbf2a1811, 32'h3e75b4d7} /* (18, 20, 10) {real, imag} */,
  {32'hbe58aa39, 32'hbd887955} /* (18, 20, 9) {real, imag} */,
  {32'hbd146d18, 32'hbf1e2ac6} /* (18, 20, 8) {real, imag} */,
  {32'h3dba321f, 32'hbe6459f0} /* (18, 20, 7) {real, imag} */,
  {32'hbe94985f, 32'hbe12654c} /* (18, 20, 6) {real, imag} */,
  {32'hbdf11a41, 32'h3e6b947e} /* (18, 20, 5) {real, imag} */,
  {32'h3d6ba57a, 32'h3dcf0cfa} /* (18, 20, 4) {real, imag} */,
  {32'h3d8ae748, 32'hbe7336c7} /* (18, 20, 3) {real, imag} */,
  {32'hbe781319, 32'h3e6fbd08} /* (18, 20, 2) {real, imag} */,
  {32'h3d78cbd0, 32'hbe9b588f} /* (18, 20, 1) {real, imag} */,
  {32'h3efbc074, 32'h3ed2bdb5} /* (18, 20, 0) {real, imag} */,
  {32'hbe03c684, 32'hbe0e70d8} /* (18, 19, 31) {real, imag} */,
  {32'h3eb084b8, 32'h3e8921ad} /* (18, 19, 30) {real, imag} */,
  {32'hbdff4f14, 32'h3eb1926f} /* (18, 19, 29) {real, imag} */,
  {32'hbdab3816, 32'hbea2c0ce} /* (18, 19, 28) {real, imag} */,
  {32'h3edf3f63, 32'h3ef40757} /* (18, 19, 27) {real, imag} */,
  {32'hbe9c215b, 32'hbebebe92} /* (18, 19, 26) {real, imag} */,
  {32'hbe99f602, 32'h3d054184} /* (18, 19, 25) {real, imag} */,
  {32'h3e5074e3, 32'h3ecf0f0c} /* (18, 19, 24) {real, imag} */,
  {32'hbe6b9820, 32'hbe72172a} /* (18, 19, 23) {real, imag} */,
  {32'hbea436ca, 32'hbe48202a} /* (18, 19, 22) {real, imag} */,
  {32'hbcb32020, 32'hbe48243f} /* (18, 19, 21) {real, imag} */,
  {32'hbe2afaee, 32'hbe553c9d} /* (18, 19, 20) {real, imag} */,
  {32'h3ea75bd6, 32'h3e141bd3} /* (18, 19, 19) {real, imag} */,
  {32'hbe913be8, 32'h3d2e6a68} /* (18, 19, 18) {real, imag} */,
  {32'h3defe730, 32'hbd81d07a} /* (18, 19, 17) {real, imag} */,
  {32'h3e193c56, 32'hbe486cae} /* (18, 19, 16) {real, imag} */,
  {32'h3e269095, 32'hbe01ee48} /* (18, 19, 15) {real, imag} */,
  {32'h3f2afe95, 32'hbe4e76b1} /* (18, 19, 14) {real, imag} */,
  {32'h3f4f8df6, 32'h3d046b88} /* (18, 19, 13) {real, imag} */,
  {32'h3f12a5e3, 32'hbd62fe00} /* (18, 19, 12) {real, imag} */,
  {32'h3db2cf65, 32'h3dce84bc} /* (18, 19, 11) {real, imag} */,
  {32'h3ee394e4, 32'hbea617c9} /* (18, 19, 10) {real, imag} */,
  {32'h3efcd9a4, 32'h3e90f20f} /* (18, 19, 9) {real, imag} */,
  {32'h3da0dfe9, 32'h3ed2fd32} /* (18, 19, 8) {real, imag} */,
  {32'hbd560818, 32'h3dd782c8} /* (18, 19, 7) {real, imag} */,
  {32'hbf5ca231, 32'h3e8aa398} /* (18, 19, 6) {real, imag} */,
  {32'hbe495cec, 32'h3ecdfaf8} /* (18, 19, 5) {real, imag} */,
  {32'hbe83f294, 32'hbd20c7d2} /* (18, 19, 4) {real, imag} */,
  {32'h3d90c27f, 32'hbd0a0c3e} /* (18, 19, 3) {real, imag} */,
  {32'h3db3000b, 32'hbf28271a} /* (18, 19, 2) {real, imag} */,
  {32'h3e785c80, 32'h3b59b580} /* (18, 19, 1) {real, imag} */,
  {32'h3d023ba0, 32'h3e6707f2} /* (18, 19, 0) {real, imag} */,
  {32'hbe914320, 32'hbe0db4d8} /* (18, 18, 31) {real, imag} */,
  {32'h3da740c4, 32'h3e3fd1aa} /* (18, 18, 30) {real, imag} */,
  {32'hbc997858, 32'hbe5aba38} /* (18, 18, 29) {real, imag} */,
  {32'h3e15b7ab, 32'hbeea5468} /* (18, 18, 28) {real, imag} */,
  {32'hbe547126, 32'hbdab1363} /* (18, 18, 27) {real, imag} */,
  {32'h3cede2a0, 32'h3e902074} /* (18, 18, 26) {real, imag} */,
  {32'hbcd527f8, 32'hb907a800} /* (18, 18, 25) {real, imag} */,
  {32'hbd903bba, 32'hbcd71880} /* (18, 18, 24) {real, imag} */,
  {32'hbdf47b00, 32'h3e727f1e} /* (18, 18, 23) {real, imag} */,
  {32'hbdd46084, 32'hbec10882} /* (18, 18, 22) {real, imag} */,
  {32'h3dbb5c68, 32'hbe328fdc} /* (18, 18, 21) {real, imag} */,
  {32'h3e0c9a88, 32'h3e9b8521} /* (18, 18, 20) {real, imag} */,
  {32'h3eaf04f0, 32'hbe0fe660} /* (18, 18, 19) {real, imag} */,
  {32'hbdfcbbf8, 32'h3ed48273} /* (18, 18, 18) {real, imag} */,
  {32'hbd5d1d06, 32'hbdd49b76} /* (18, 18, 17) {real, imag} */,
  {32'hbe2fcc62, 32'hbc7c52a0} /* (18, 18, 16) {real, imag} */,
  {32'h3e1c0bea, 32'h3c09dd08} /* (18, 18, 15) {real, imag} */,
  {32'h3e193e0e, 32'hbd5a3282} /* (18, 18, 14) {real, imag} */,
  {32'h3ef118d8, 32'hbea488ee} /* (18, 18, 13) {real, imag} */,
  {32'hbb6e5fa0, 32'h3f0146bb} /* (18, 18, 12) {real, imag} */,
  {32'hbd37d1c4, 32'h3f30feae} /* (18, 18, 11) {real, imag} */,
  {32'h3e4be98c, 32'h3d9e1ef2} /* (18, 18, 10) {real, imag} */,
  {32'hbc976348, 32'hbe94b996} /* (18, 18, 9) {real, imag} */,
  {32'h3d3f8f1c, 32'h3eca5870} /* (18, 18, 8) {real, imag} */,
  {32'hbee9c87e, 32'h3c09d020} /* (18, 18, 7) {real, imag} */,
  {32'hbec1ed54, 32'hbcb23ae6} /* (18, 18, 6) {real, imag} */,
  {32'hbe4c7bb3, 32'h3eba3adc} /* (18, 18, 5) {real, imag} */,
  {32'hbe4818e0, 32'hbe583ee0} /* (18, 18, 4) {real, imag} */,
  {32'h3e8229c5, 32'hbd05c548} /* (18, 18, 3) {real, imag} */,
  {32'hbddb84a6, 32'h3e17f9b6} /* (18, 18, 2) {real, imag} */,
  {32'h3e7468b1, 32'hbecf1a22} /* (18, 18, 1) {real, imag} */,
  {32'h3ed72fe8, 32'hbeafd0ac} /* (18, 18, 0) {real, imag} */,
  {32'hbd90ab79, 32'h3f047832} /* (18, 17, 31) {real, imag} */,
  {32'hbd818330, 32'h3e537c10} /* (18, 17, 30) {real, imag} */,
  {32'hbe5f6b56, 32'hbd1f5236} /* (18, 17, 29) {real, imag} */,
  {32'hbd2438ee, 32'h3db9b613} /* (18, 17, 28) {real, imag} */,
  {32'h3e777f08, 32'hbeebef3c} /* (18, 17, 27) {real, imag} */,
  {32'hbd289141, 32'h3e075d0a} /* (18, 17, 26) {real, imag} */,
  {32'h3eb1ab08, 32'hbc3a9880} /* (18, 17, 25) {real, imag} */,
  {32'h3e1d44fa, 32'hbf05dc2f} /* (18, 17, 24) {real, imag} */,
  {32'h3e0a41d4, 32'h3d0c85e4} /* (18, 17, 23) {real, imag} */,
  {32'hbd4317b0, 32'hbecb2fed} /* (18, 17, 22) {real, imag} */,
  {32'hbe4b8611, 32'h3dab6fa6} /* (18, 17, 21) {real, imag} */,
  {32'h3e913122, 32'hbb15dac0} /* (18, 17, 20) {real, imag} */,
  {32'hbd0f7988, 32'h3ea15de0} /* (18, 17, 19) {real, imag} */,
  {32'h3c981a3a, 32'h3e9b3cef} /* (18, 17, 18) {real, imag} */,
  {32'h3d04c8a2, 32'h3e435e68} /* (18, 17, 17) {real, imag} */,
  {32'hbbe33367, 32'hbe236c66} /* (18, 17, 16) {real, imag} */,
  {32'hbe0d5c5a, 32'h3dd6d4d2} /* (18, 17, 15) {real, imag} */,
  {32'h3e7e5e06, 32'h3e4747d7} /* (18, 17, 14) {real, imag} */,
  {32'h3ecca010, 32'hbe8f3f06} /* (18, 17, 13) {real, imag} */,
  {32'hbea40fc0, 32'h3e8b41c7} /* (18, 17, 12) {real, imag} */,
  {32'h3da8f351, 32'hbdd58d10} /* (18, 17, 11) {real, imag} */,
  {32'h3ebf876f, 32'hbcda6edc} /* (18, 17, 10) {real, imag} */,
  {32'h3ee2d4c5, 32'h3d51513c} /* (18, 17, 9) {real, imag} */,
  {32'hbd95a1db, 32'h3de41724} /* (18, 17, 8) {real, imag} */,
  {32'hbe3f6779, 32'hbe8c2d3c} /* (18, 17, 7) {real, imag} */,
  {32'hbe78e602, 32'hbe18da7c} /* (18, 17, 6) {real, imag} */,
  {32'h3d36a354, 32'hbe530de6} /* (18, 17, 5) {real, imag} */,
  {32'h3cd2481e, 32'hbe3a9d16} /* (18, 17, 4) {real, imag} */,
  {32'hbdcf0e2a, 32'hbe295ce9} /* (18, 17, 3) {real, imag} */,
  {32'h3ce31588, 32'h3d028b10} /* (18, 17, 2) {real, imag} */,
  {32'hbdf217f4, 32'hbd1854ee} /* (18, 17, 1) {real, imag} */,
  {32'h3e09569a, 32'h3cced984} /* (18, 17, 0) {real, imag} */,
  {32'hbd9f8ef4, 32'h3e1d9620} /* (18, 16, 31) {real, imag} */,
  {32'hbe86bc9f, 32'hbe62ce3a} /* (18, 16, 30) {real, imag} */,
  {32'hbc048458, 32'hbda47f48} /* (18, 16, 29) {real, imag} */,
  {32'h3ee1b9ed, 32'h3e64aa08} /* (18, 16, 28) {real, imag} */,
  {32'h3d9608c0, 32'h3e12739a} /* (18, 16, 27) {real, imag} */,
  {32'hbe25423e, 32'hbe9d1af2} /* (18, 16, 26) {real, imag} */,
  {32'hbd2a88e6, 32'hbed23414} /* (18, 16, 25) {real, imag} */,
  {32'hbcb464c8, 32'h3d6c91d0} /* (18, 16, 24) {real, imag} */,
  {32'h3db6db4e, 32'h3e1fccb9} /* (18, 16, 23) {real, imag} */,
  {32'hbe01086b, 32'h3e9766cc} /* (18, 16, 22) {real, imag} */,
  {32'h3d701a48, 32'hbe5d3282} /* (18, 16, 21) {real, imag} */,
  {32'h3d5a77be, 32'h3e6240a3} /* (18, 16, 20) {real, imag} */,
  {32'h3e40f6eb, 32'h3d0cc7a8} /* (18, 16, 19) {real, imag} */,
  {32'hbdac5b1f, 32'h3c552300} /* (18, 16, 18) {real, imag} */,
  {32'hbd815bff, 32'hbe4456f6} /* (18, 16, 17) {real, imag} */,
  {32'hbeb61599, 32'h00000000} /* (18, 16, 16) {real, imag} */,
  {32'hbd815bff, 32'h3e4456f6} /* (18, 16, 15) {real, imag} */,
  {32'hbdac5b1f, 32'hbc552300} /* (18, 16, 14) {real, imag} */,
  {32'h3e40f6eb, 32'hbd0cc7a8} /* (18, 16, 13) {real, imag} */,
  {32'h3d5a77be, 32'hbe6240a3} /* (18, 16, 12) {real, imag} */,
  {32'h3d701a48, 32'h3e5d3282} /* (18, 16, 11) {real, imag} */,
  {32'hbe01086b, 32'hbe9766cc} /* (18, 16, 10) {real, imag} */,
  {32'h3db6db4e, 32'hbe1fccb9} /* (18, 16, 9) {real, imag} */,
  {32'hbcb464c8, 32'hbd6c91d0} /* (18, 16, 8) {real, imag} */,
  {32'hbd2a88e6, 32'h3ed23414} /* (18, 16, 7) {real, imag} */,
  {32'hbe25423e, 32'h3e9d1af2} /* (18, 16, 6) {real, imag} */,
  {32'h3d9608c0, 32'hbe12739a} /* (18, 16, 5) {real, imag} */,
  {32'h3ee1b9ed, 32'hbe64aa08} /* (18, 16, 4) {real, imag} */,
  {32'hbc048458, 32'h3da47f48} /* (18, 16, 3) {real, imag} */,
  {32'hbe86bc9f, 32'h3e62ce3a} /* (18, 16, 2) {real, imag} */,
  {32'hbd9f8ef4, 32'hbe1d9620} /* (18, 16, 1) {real, imag} */,
  {32'hbd890c88, 32'h00000000} /* (18, 16, 0) {real, imag} */,
  {32'hbdf217f4, 32'h3d1854ee} /* (18, 15, 31) {real, imag} */,
  {32'h3ce31588, 32'hbd028b10} /* (18, 15, 30) {real, imag} */,
  {32'hbdcf0e2a, 32'h3e295ce9} /* (18, 15, 29) {real, imag} */,
  {32'h3cd2481e, 32'h3e3a9d16} /* (18, 15, 28) {real, imag} */,
  {32'h3d36a354, 32'h3e530de6} /* (18, 15, 27) {real, imag} */,
  {32'hbe78e602, 32'h3e18da7c} /* (18, 15, 26) {real, imag} */,
  {32'hbe3f6779, 32'h3e8c2d3c} /* (18, 15, 25) {real, imag} */,
  {32'hbd95a1db, 32'hbde41724} /* (18, 15, 24) {real, imag} */,
  {32'h3ee2d4c5, 32'hbd51513c} /* (18, 15, 23) {real, imag} */,
  {32'h3ebf876f, 32'h3cda6edc} /* (18, 15, 22) {real, imag} */,
  {32'h3da8f351, 32'h3dd58d10} /* (18, 15, 21) {real, imag} */,
  {32'hbea40fc0, 32'hbe8b41c7} /* (18, 15, 20) {real, imag} */,
  {32'h3ecca010, 32'h3e8f3f06} /* (18, 15, 19) {real, imag} */,
  {32'h3e7e5e06, 32'hbe4747d7} /* (18, 15, 18) {real, imag} */,
  {32'hbe0d5c5a, 32'hbdd6d4d2} /* (18, 15, 17) {real, imag} */,
  {32'hbbe33367, 32'h3e236c66} /* (18, 15, 16) {real, imag} */,
  {32'h3d04c8a2, 32'hbe435e68} /* (18, 15, 15) {real, imag} */,
  {32'h3c981a3a, 32'hbe9b3cef} /* (18, 15, 14) {real, imag} */,
  {32'hbd0f7988, 32'hbea15de0} /* (18, 15, 13) {real, imag} */,
  {32'h3e913122, 32'h3b15dac0} /* (18, 15, 12) {real, imag} */,
  {32'hbe4b8611, 32'hbdab6fa6} /* (18, 15, 11) {real, imag} */,
  {32'hbd4317b0, 32'h3ecb2fed} /* (18, 15, 10) {real, imag} */,
  {32'h3e0a41d4, 32'hbd0c85e4} /* (18, 15, 9) {real, imag} */,
  {32'h3e1d44fa, 32'h3f05dc2f} /* (18, 15, 8) {real, imag} */,
  {32'h3eb1ab08, 32'h3c3a9880} /* (18, 15, 7) {real, imag} */,
  {32'hbd289141, 32'hbe075d0a} /* (18, 15, 6) {real, imag} */,
  {32'h3e777f08, 32'h3eebef3c} /* (18, 15, 5) {real, imag} */,
  {32'hbd2438ee, 32'hbdb9b613} /* (18, 15, 4) {real, imag} */,
  {32'hbe5f6b56, 32'h3d1f5236} /* (18, 15, 3) {real, imag} */,
  {32'hbd818330, 32'hbe537c10} /* (18, 15, 2) {real, imag} */,
  {32'hbd90ab79, 32'hbf047832} /* (18, 15, 1) {real, imag} */,
  {32'h3e09569a, 32'hbcced984} /* (18, 15, 0) {real, imag} */,
  {32'h3e7468b1, 32'h3ecf1a22} /* (18, 14, 31) {real, imag} */,
  {32'hbddb84a6, 32'hbe17f9b6} /* (18, 14, 30) {real, imag} */,
  {32'h3e8229c5, 32'h3d05c548} /* (18, 14, 29) {real, imag} */,
  {32'hbe4818e0, 32'h3e583ee0} /* (18, 14, 28) {real, imag} */,
  {32'hbe4c7bb3, 32'hbeba3adc} /* (18, 14, 27) {real, imag} */,
  {32'hbec1ed54, 32'h3cb23ae6} /* (18, 14, 26) {real, imag} */,
  {32'hbee9c87e, 32'hbc09d020} /* (18, 14, 25) {real, imag} */,
  {32'h3d3f8f1c, 32'hbeca5870} /* (18, 14, 24) {real, imag} */,
  {32'hbc976348, 32'h3e94b996} /* (18, 14, 23) {real, imag} */,
  {32'h3e4be98c, 32'hbd9e1ef2} /* (18, 14, 22) {real, imag} */,
  {32'hbd37d1c4, 32'hbf30feae} /* (18, 14, 21) {real, imag} */,
  {32'hbb6e5fa0, 32'hbf0146bb} /* (18, 14, 20) {real, imag} */,
  {32'h3ef118d8, 32'h3ea488ee} /* (18, 14, 19) {real, imag} */,
  {32'h3e193e0e, 32'h3d5a3282} /* (18, 14, 18) {real, imag} */,
  {32'h3e1c0bea, 32'hbc09dd08} /* (18, 14, 17) {real, imag} */,
  {32'hbe2fcc62, 32'h3c7c52a0} /* (18, 14, 16) {real, imag} */,
  {32'hbd5d1d06, 32'h3dd49b76} /* (18, 14, 15) {real, imag} */,
  {32'hbdfcbbf8, 32'hbed48273} /* (18, 14, 14) {real, imag} */,
  {32'h3eaf04f0, 32'h3e0fe660} /* (18, 14, 13) {real, imag} */,
  {32'h3e0c9a88, 32'hbe9b8521} /* (18, 14, 12) {real, imag} */,
  {32'h3dbb5c68, 32'h3e328fdc} /* (18, 14, 11) {real, imag} */,
  {32'hbdd46084, 32'h3ec10882} /* (18, 14, 10) {real, imag} */,
  {32'hbdf47b00, 32'hbe727f1e} /* (18, 14, 9) {real, imag} */,
  {32'hbd903bba, 32'h3cd71880} /* (18, 14, 8) {real, imag} */,
  {32'hbcd527f8, 32'h3907a800} /* (18, 14, 7) {real, imag} */,
  {32'h3cede2a0, 32'hbe902074} /* (18, 14, 6) {real, imag} */,
  {32'hbe547126, 32'h3dab1363} /* (18, 14, 5) {real, imag} */,
  {32'h3e15b7ab, 32'h3eea5468} /* (18, 14, 4) {real, imag} */,
  {32'hbc997858, 32'h3e5aba38} /* (18, 14, 3) {real, imag} */,
  {32'h3da740c4, 32'hbe3fd1aa} /* (18, 14, 2) {real, imag} */,
  {32'hbe914320, 32'h3e0db4d8} /* (18, 14, 1) {real, imag} */,
  {32'h3ed72fe8, 32'h3eafd0ac} /* (18, 14, 0) {real, imag} */,
  {32'h3e785c80, 32'hbb59b580} /* (18, 13, 31) {real, imag} */,
  {32'h3db3000b, 32'h3f28271a} /* (18, 13, 30) {real, imag} */,
  {32'h3d90c27f, 32'h3d0a0c3e} /* (18, 13, 29) {real, imag} */,
  {32'hbe83f294, 32'h3d20c7d2} /* (18, 13, 28) {real, imag} */,
  {32'hbe495cec, 32'hbecdfaf8} /* (18, 13, 27) {real, imag} */,
  {32'hbf5ca231, 32'hbe8aa398} /* (18, 13, 26) {real, imag} */,
  {32'hbd560818, 32'hbdd782c8} /* (18, 13, 25) {real, imag} */,
  {32'h3da0dfe9, 32'hbed2fd32} /* (18, 13, 24) {real, imag} */,
  {32'h3efcd9a4, 32'hbe90f20f} /* (18, 13, 23) {real, imag} */,
  {32'h3ee394e4, 32'h3ea617c9} /* (18, 13, 22) {real, imag} */,
  {32'h3db2cf65, 32'hbdce84bc} /* (18, 13, 21) {real, imag} */,
  {32'h3f12a5e3, 32'h3d62fe00} /* (18, 13, 20) {real, imag} */,
  {32'h3f4f8df6, 32'hbd046b88} /* (18, 13, 19) {real, imag} */,
  {32'h3f2afe95, 32'h3e4e76b1} /* (18, 13, 18) {real, imag} */,
  {32'h3e269095, 32'h3e01ee48} /* (18, 13, 17) {real, imag} */,
  {32'h3e193c56, 32'h3e486cae} /* (18, 13, 16) {real, imag} */,
  {32'h3defe730, 32'h3d81d07a} /* (18, 13, 15) {real, imag} */,
  {32'hbe913be8, 32'hbd2e6a68} /* (18, 13, 14) {real, imag} */,
  {32'h3ea75bd6, 32'hbe141bd3} /* (18, 13, 13) {real, imag} */,
  {32'hbe2afaee, 32'h3e553c9d} /* (18, 13, 12) {real, imag} */,
  {32'hbcb32020, 32'h3e48243f} /* (18, 13, 11) {real, imag} */,
  {32'hbea436ca, 32'h3e48202a} /* (18, 13, 10) {real, imag} */,
  {32'hbe6b9820, 32'h3e72172a} /* (18, 13, 9) {real, imag} */,
  {32'h3e5074e3, 32'hbecf0f0c} /* (18, 13, 8) {real, imag} */,
  {32'hbe99f602, 32'hbd054184} /* (18, 13, 7) {real, imag} */,
  {32'hbe9c215b, 32'h3ebebe92} /* (18, 13, 6) {real, imag} */,
  {32'h3edf3f63, 32'hbef40757} /* (18, 13, 5) {real, imag} */,
  {32'hbdab3816, 32'h3ea2c0ce} /* (18, 13, 4) {real, imag} */,
  {32'hbdff4f14, 32'hbeb1926f} /* (18, 13, 3) {real, imag} */,
  {32'h3eb084b8, 32'hbe8921ad} /* (18, 13, 2) {real, imag} */,
  {32'hbe03c684, 32'h3e0e70d8} /* (18, 13, 1) {real, imag} */,
  {32'h3d023ba0, 32'hbe6707f2} /* (18, 13, 0) {real, imag} */,
  {32'h3d78cbd0, 32'h3e9b588f} /* (18, 12, 31) {real, imag} */,
  {32'hbe781319, 32'hbe6fbd08} /* (18, 12, 30) {real, imag} */,
  {32'h3d8ae748, 32'h3e7336c7} /* (18, 12, 29) {real, imag} */,
  {32'h3d6ba57a, 32'hbdcf0cfa} /* (18, 12, 28) {real, imag} */,
  {32'hbdf11a41, 32'hbe6b947e} /* (18, 12, 27) {real, imag} */,
  {32'hbe94985f, 32'h3e12654c} /* (18, 12, 26) {real, imag} */,
  {32'h3dba321f, 32'h3e6459f0} /* (18, 12, 25) {real, imag} */,
  {32'hbd146d18, 32'h3f1e2ac6} /* (18, 12, 24) {real, imag} */,
  {32'hbe58aa39, 32'h3d887955} /* (18, 12, 23) {real, imag} */,
  {32'hbf2a1811, 32'hbe75b4d7} /* (18, 12, 22) {real, imag} */,
  {32'hbe9adb9e, 32'h3e99041b} /* (18, 12, 21) {real, imag} */,
  {32'h3f38c16e, 32'h3e0f9ed5} /* (18, 12, 20) {real, imag} */,
  {32'hbec3d6e6, 32'hbe5ff217} /* (18, 12, 19) {real, imag} */,
  {32'h3e424968, 32'hbbed0740} /* (18, 12, 18) {real, imag} */,
  {32'hbe54ca73, 32'hbde2dc40} /* (18, 12, 17) {real, imag} */,
  {32'hbe6976dd, 32'hbdf85484} /* (18, 12, 16) {real, imag} */,
  {32'h3eb32505, 32'h3e1bcb72} /* (18, 12, 15) {real, imag} */,
  {32'hbecc83f8, 32'hbea0a826} /* (18, 12, 14) {real, imag} */,
  {32'h3c995ed2, 32'hbdeb5256} /* (18, 12, 13) {real, imag} */,
  {32'h3e8646c0, 32'h3ef13927} /* (18, 12, 12) {real, imag} */,
  {32'hbe3d57c4, 32'h3d821a76} /* (18, 12, 11) {real, imag} */,
  {32'hbcbd1448, 32'h3db7bd7e} /* (18, 12, 10) {real, imag} */,
  {32'hbe73b0b3, 32'h3e1bdef0} /* (18, 12, 9) {real, imag} */,
  {32'h3be5a7a0, 32'hbed97184} /* (18, 12, 8) {real, imag} */,
  {32'hbe824209, 32'hbf2a681b} /* (18, 12, 7) {real, imag} */,
  {32'hbea62a54, 32'hbdb508e0} /* (18, 12, 6) {real, imag} */,
  {32'h3de8e0ec, 32'h3c64886c} /* (18, 12, 5) {real, imag} */,
  {32'h3d9091fa, 32'hbe22173d} /* (18, 12, 4) {real, imag} */,
  {32'hbe0ff586, 32'hbe8bad8c} /* (18, 12, 3) {real, imag} */,
  {32'hbf1ab664, 32'h3d494cb4} /* (18, 12, 2) {real, imag} */,
  {32'hbdc71fb0, 32'h3eb29c2f} /* (18, 12, 1) {real, imag} */,
  {32'h3efbc074, 32'hbed2bdb5} /* (18, 12, 0) {real, imag} */,
  {32'h3e27949a, 32'h3db2d392} /* (18, 11, 31) {real, imag} */,
  {32'hbee54173, 32'hbeb051e9} /* (18, 11, 30) {real, imag} */,
  {32'hbea242b6, 32'hbee70ba4} /* (18, 11, 29) {real, imag} */,
  {32'h3b3e9a60, 32'h3e2240e0} /* (18, 11, 28) {real, imag} */,
  {32'h3e7dd55c, 32'h3cf30590} /* (18, 11, 27) {real, imag} */,
  {32'h3ee88b53, 32'h3eb5c210} /* (18, 11, 26) {real, imag} */,
  {32'h3f4eef9f, 32'hbe3fd62d} /* (18, 11, 25) {real, imag} */,
  {32'hbe567d52, 32'hbeb5009c} /* (18, 11, 24) {real, imag} */,
  {32'hbec86ea6, 32'hbf1eb80c} /* (18, 11, 23) {real, imag} */,
  {32'h3f175be4, 32'h3d84661f} /* (18, 11, 22) {real, imag} */,
  {32'hbe910e78, 32'hbe5f91bc} /* (18, 11, 21) {real, imag} */,
  {32'h3ca4a95c, 32'hbecb7288} /* (18, 11, 20) {real, imag} */,
  {32'h3ec11eba, 32'hbdfc059d} /* (18, 11, 19) {real, imag} */,
  {32'h3dc32bd9, 32'hbdc6f8c0} /* (18, 11, 18) {real, imag} */,
  {32'h3e177e5a, 32'hbdb3235f} /* (18, 11, 17) {real, imag} */,
  {32'hbe04fb12, 32'h3e7f6a4e} /* (18, 11, 16) {real, imag} */,
  {32'hbf15541a, 32'h3eaa9232} /* (18, 11, 15) {real, imag} */,
  {32'h3db18192, 32'hbec55b0f} /* (18, 11, 14) {real, imag} */,
  {32'hbe9898c2, 32'hbea02b0a} /* (18, 11, 13) {real, imag} */,
  {32'hbef453a6, 32'hbe6b7c6a} /* (18, 11, 12) {real, imag} */,
  {32'h3f383316, 32'hbe5a4636} /* (18, 11, 11) {real, imag} */,
  {32'h3e966274, 32'hbdc3d304} /* (18, 11, 10) {real, imag} */,
  {32'hbe38f910, 32'hbbcff0e0} /* (18, 11, 9) {real, imag} */,
  {32'h3f283fa8, 32'h3d30e27a} /* (18, 11, 8) {real, imag} */,
  {32'h3ea42938, 32'hbe5ce20e} /* (18, 11, 7) {real, imag} */,
  {32'h3e912699, 32'h3e8ea340} /* (18, 11, 6) {real, imag} */,
  {32'h3de65f6a, 32'hbf54a1aa} /* (18, 11, 5) {real, imag} */,
  {32'hbd4c9dab, 32'h3f0aad2d} /* (18, 11, 4) {real, imag} */,
  {32'hbef3c868, 32'h3f343d52} /* (18, 11, 3) {real, imag} */,
  {32'h3d568bd0, 32'hbec01b0b} /* (18, 11, 2) {real, imag} */,
  {32'hbcf75106, 32'h3f616006} /* (18, 11, 1) {real, imag} */,
  {32'h3e920752, 32'h3edcedeb} /* (18, 11, 0) {real, imag} */,
  {32'h3d217b12, 32'h3af9db00} /* (18, 10, 31) {real, imag} */,
  {32'h3e62a9d2, 32'hbed4acbc} /* (18, 10, 30) {real, imag} */,
  {32'hbe5a7cd1, 32'hbe99c3af} /* (18, 10, 29) {real, imag} */,
  {32'hbd7ea7b0, 32'h3e09e608} /* (18, 10, 28) {real, imag} */,
  {32'h3e271518, 32'h3dbddb87} /* (18, 10, 27) {real, imag} */,
  {32'h3d9aabf8, 32'h3d76384c} /* (18, 10, 26) {real, imag} */,
  {32'hbc7aac60, 32'hbd9c2600} /* (18, 10, 25) {real, imag} */,
  {32'hbe50b588, 32'hbd0f53dc} /* (18, 10, 24) {real, imag} */,
  {32'hbe8687d9, 32'h3f281e12} /* (18, 10, 23) {real, imag} */,
  {32'hbe1e4ee4, 32'hbf146131} /* (18, 10, 22) {real, imag} */,
  {32'hbe0763cf, 32'hbd914954} /* (18, 10, 21) {real, imag} */,
  {32'hbd916647, 32'hbe718d64} /* (18, 10, 20) {real, imag} */,
  {32'h3dcb12f6, 32'hbe79e3d5} /* (18, 10, 19) {real, imag} */,
  {32'hbd85bf93, 32'hbe97de0c} /* (18, 10, 18) {real, imag} */,
  {32'hbd8d049e, 32'hbe1d2cdc} /* (18, 10, 17) {real, imag} */,
  {32'h3d151248, 32'h3df41b0d} /* (18, 10, 16) {real, imag} */,
  {32'hbe37933e, 32'hbed0bcde} /* (18, 10, 15) {real, imag} */,
  {32'h3e590ee0, 32'hbe894de2} /* (18, 10, 14) {real, imag} */,
  {32'hbed67cb2, 32'h3e0aca7a} /* (18, 10, 13) {real, imag} */,
  {32'h3e8fedc9, 32'hbdab1f58} /* (18, 10, 12) {real, imag} */,
  {32'h3f04e3d5, 32'h3ebafa88} /* (18, 10, 11) {real, imag} */,
  {32'h3e09aa15, 32'h3ef4da06} /* (18, 10, 10) {real, imag} */,
  {32'hbe1a4fbf, 32'h3d0395a0} /* (18, 10, 9) {real, imag} */,
  {32'h3d800aec, 32'h3de84340} /* (18, 10, 8) {real, imag} */,
  {32'hbc3373b0, 32'h3b8b2b70} /* (18, 10, 7) {real, imag} */,
  {32'hbf09c652, 32'hbef0b666} /* (18, 10, 6) {real, imag} */,
  {32'hbedc4ef8, 32'h3ea7c67e} /* (18, 10, 5) {real, imag} */,
  {32'hbed135be, 32'hbf0c9a5a} /* (18, 10, 4) {real, imag} */,
  {32'hbf78cd7c, 32'hbe8b0f55} /* (18, 10, 3) {real, imag} */,
  {32'h3f023b0a, 32'h3f58cadc} /* (18, 10, 2) {real, imag} */,
  {32'hbf115382, 32'hbeaa47fe} /* (18, 10, 1) {real, imag} */,
  {32'h3f051758, 32'h3d10f790} /* (18, 10, 0) {real, imag} */,
  {32'h3e478cdb, 32'hbe5d63b0} /* (18, 9, 31) {real, imag} */,
  {32'hbbe86ec0, 32'h3f9fe30a} /* (18, 9, 30) {real, imag} */,
  {32'h3f0dcb36, 32'h3d9c2207} /* (18, 9, 29) {real, imag} */,
  {32'hbf068147, 32'hbeaa71f0} /* (18, 9, 28) {real, imag} */,
  {32'h3e2ed934, 32'hbedc8344} /* (18, 9, 27) {real, imag} */,
  {32'hbe1638e5, 32'hbf170567} /* (18, 9, 26) {real, imag} */,
  {32'hbecea782, 32'h3f28d47c} /* (18, 9, 25) {real, imag} */,
  {32'h3f07a1f6, 32'hbea7810c} /* (18, 9, 24) {real, imag} */,
  {32'hbe5fe69c, 32'h3f2127d8} /* (18, 9, 23) {real, imag} */,
  {32'h3ee022a2, 32'hbf32e552} /* (18, 9, 22) {real, imag} */,
  {32'h3eba3d79, 32'h3e4a3648} /* (18, 9, 21) {real, imag} */,
  {32'hbe60aa19, 32'h3efd1e83} /* (18, 9, 20) {real, imag} */,
  {32'hbe4e54b8, 32'hbe86b5ed} /* (18, 9, 19) {real, imag} */,
  {32'h3e4d74d0, 32'hbee29c12} /* (18, 9, 18) {real, imag} */,
  {32'h3e02275e, 32'h3f1f6ffe} /* (18, 9, 17) {real, imag} */,
  {32'h3ef09a9a, 32'hbe33cd96} /* (18, 9, 16) {real, imag} */,
  {32'h3d2f3662, 32'h3e1891d4} /* (18, 9, 15) {real, imag} */,
  {32'hbe327778, 32'h3d821d5f} /* (18, 9, 14) {real, imag} */,
  {32'h3e147e26, 32'h3ed8895c} /* (18, 9, 13) {real, imag} */,
  {32'hbea57953, 32'hbe02c6f6} /* (18, 9, 12) {real, imag} */,
  {32'hbf623c80, 32'h3f1eb781} /* (18, 9, 11) {real, imag} */,
  {32'h3cba56f8, 32'h3f28a20a} /* (18, 9, 10) {real, imag} */,
  {32'hbecf78c0, 32'hbf1289ae} /* (18, 9, 9) {real, imag} */,
  {32'hbe70c392, 32'hbd5ada28} /* (18, 9, 8) {real, imag} */,
  {32'hbea29d3d, 32'h3c807ea0} /* (18, 9, 7) {real, imag} */,
  {32'h3e7ad470, 32'hbe67c5b1} /* (18, 9, 6) {real, imag} */,
  {32'hbeb5dedb, 32'h3e2eca4a} /* (18, 9, 5) {real, imag} */,
  {32'h3d873d34, 32'hbf53ee12} /* (18, 9, 4) {real, imag} */,
  {32'hbe4cf12d, 32'h3df65444} /* (18, 9, 3) {real, imag} */,
  {32'hbdbf16a6, 32'h3ef7edee} /* (18, 9, 2) {real, imag} */,
  {32'hbd0c24c0, 32'hbec2a79b} /* (18, 9, 1) {real, imag} */,
  {32'h3e5b0059, 32'hbdc55da4} /* (18, 9, 0) {real, imag} */,
  {32'h3fccb150, 32'h3f8c0d71} /* (18, 8, 31) {real, imag} */,
  {32'hbf9f0f48, 32'h3e0cdccf} /* (18, 8, 30) {real, imag} */,
  {32'h3c8ac2b0, 32'hbe79037a} /* (18, 8, 29) {real, imag} */,
  {32'h3e466a80, 32'h3f1a2a99} /* (18, 8, 28) {real, imag} */,
  {32'hbed8047c, 32'hbdb3f9b5} /* (18, 8, 27) {real, imag} */,
  {32'hbe428a4a, 32'hbe8ef21a} /* (18, 8, 26) {real, imag} */,
  {32'h3ef4a263, 32'hbea1575e} /* (18, 8, 25) {real, imag} */,
  {32'hbdf0c720, 32'hbe8e75bc} /* (18, 8, 24) {real, imag} */,
  {32'hbed357be, 32'h3ebdadf3} /* (18, 8, 23) {real, imag} */,
  {32'hbf2bd018, 32'h3dadbc82} /* (18, 8, 22) {real, imag} */,
  {32'hbf02fa47, 32'h3e2c5295} /* (18, 8, 21) {real, imag} */,
  {32'h3e9f8ebc, 32'hbebf807a} /* (18, 8, 20) {real, imag} */,
  {32'h3f03e79c, 32'h3e04c6cd} /* (18, 8, 19) {real, imag} */,
  {32'h3e4aa6c5, 32'hbd9e00e6} /* (18, 8, 18) {real, imag} */,
  {32'hbe3e9580, 32'hbe0e6074} /* (18, 8, 17) {real, imag} */,
  {32'hbe693a5a, 32'h3e00ea24} /* (18, 8, 16) {real, imag} */,
  {32'hbded8e70, 32'h3ca67500} /* (18, 8, 15) {real, imag} */,
  {32'h3e06e7fa, 32'hbd7c4b12} /* (18, 8, 14) {real, imag} */,
  {32'hbeb787b9, 32'hbe7c9629} /* (18, 8, 13) {real, imag} */,
  {32'h3e88072e, 32'h3cdab0d0} /* (18, 8, 12) {real, imag} */,
  {32'h3f0360e8, 32'h3d473e58} /* (18, 8, 11) {real, imag} */,
  {32'h3e309488, 32'hbf19dc28} /* (18, 8, 10) {real, imag} */,
  {32'h3e05f377, 32'hbe24cfda} /* (18, 8, 9) {real, imag} */,
  {32'hbe67807a, 32'h3e817f57} /* (18, 8, 8) {real, imag} */,
  {32'hbca587d0, 32'hbac17440} /* (18, 8, 7) {real, imag} */,
  {32'h3e723594, 32'hbe369b9d} /* (18, 8, 6) {real, imag} */,
  {32'h3d895815, 32'hbd382808} /* (18, 8, 5) {real, imag} */,
  {32'h3e1db65a, 32'h3d9c4b41} /* (18, 8, 4) {real, imag} */,
  {32'hbda844fa, 32'h3d1fa0ba} /* (18, 8, 3) {real, imag} */,
  {32'hbf2e4f33, 32'hbf279fd2} /* (18, 8, 2) {real, imag} */,
  {32'h3f24a274, 32'h3f3bd90e} /* (18, 8, 1) {real, imag} */,
  {32'h3f0bae06, 32'h3f8b0557} /* (18, 8, 0) {real, imag} */,
  {32'hbe44742c, 32'hbf13fe1e} /* (18, 7, 31) {real, imag} */,
  {32'h3f426626, 32'hbdd72550} /* (18, 7, 30) {real, imag} */,
  {32'hbe9937b0, 32'hbe65547d} /* (18, 7, 29) {real, imag} */,
  {32'h3ebce270, 32'h3e576006} /* (18, 7, 28) {real, imag} */,
  {32'h3f11ff38, 32'h3de129e4} /* (18, 7, 27) {real, imag} */,
  {32'h3eca1bd6, 32'hbeae77c7} /* (18, 7, 26) {real, imag} */,
  {32'hbf2a3959, 32'hbf40d96e} /* (18, 7, 25) {real, imag} */,
  {32'hbd26c28c, 32'hbe2a817a} /* (18, 7, 24) {real, imag} */,
  {32'h3ea69425, 32'h3edf2b09} /* (18, 7, 23) {real, imag} */,
  {32'hbed53b6e, 32'hbd4d63ab} /* (18, 7, 22) {real, imag} */,
  {32'hbe461a6a, 32'h3eb12c68} /* (18, 7, 21) {real, imag} */,
  {32'h3e76a654, 32'h3d7f5270} /* (18, 7, 20) {real, imag} */,
  {32'hbee0bc04, 32'hbdb54315} /* (18, 7, 19) {real, imag} */,
  {32'h3e9cc670, 32'h3ee57840} /* (18, 7, 18) {real, imag} */,
  {32'hbdaf4798, 32'hbeb0e194} /* (18, 7, 17) {real, imag} */,
  {32'hbdeee27a, 32'h3d0887fc} /* (18, 7, 16) {real, imag} */,
  {32'hbe0cf666, 32'hbe438f80} /* (18, 7, 15) {real, imag} */,
  {32'h3c447380, 32'h3f124975} /* (18, 7, 14) {real, imag} */,
  {32'hbe752dd1, 32'hbdeb7948} /* (18, 7, 13) {real, imag} */,
  {32'h3e9c2a00, 32'h3d7769c0} /* (18, 7, 12) {real, imag} */,
  {32'h3e2df2c6, 32'h3eafe1f8} /* (18, 7, 11) {real, imag} */,
  {32'hbedb5c64, 32'h3c2f7600} /* (18, 7, 10) {real, imag} */,
  {32'hbf16f172, 32'h3e3d4130} /* (18, 7, 9) {real, imag} */,
  {32'hbee6ffde, 32'hbf4397ce} /* (18, 7, 8) {real, imag} */,
  {32'hbeff0cb9, 32'h3f032600} /* (18, 7, 7) {real, imag} */,
  {32'h3e894ff2, 32'h3db37177} /* (18, 7, 6) {real, imag} */,
  {32'hbede64c0, 32'hbe90fce9} /* (18, 7, 5) {real, imag} */,
  {32'h3f015c3c, 32'h3f09f8f7} /* (18, 7, 4) {real, imag} */,
  {32'h3da74128, 32'h3dc0ae17} /* (18, 7, 3) {real, imag} */,
  {32'h3e99782c, 32'h3f4ac280} /* (18, 7, 2) {real, imag} */,
  {32'hbe889c61, 32'hbedefa54} /* (18, 7, 1) {real, imag} */,
  {32'hbe865c86, 32'hbee8a097} /* (18, 7, 0) {real, imag} */,
  {32'h3e968407, 32'hbe4a0da9} /* (18, 6, 31) {real, imag} */,
  {32'hbec7e3fb, 32'hbf34bcdb} /* (18, 6, 30) {real, imag} */,
  {32'hbf7947a8, 32'h3e1bfaea} /* (18, 6, 29) {real, imag} */,
  {32'hbe8bdb60, 32'h3da2d910} /* (18, 6, 28) {real, imag} */,
  {32'hbf03ae76, 32'h3e162556} /* (18, 6, 27) {real, imag} */,
  {32'h3cc52a8c, 32'hbe664c6c} /* (18, 6, 26) {real, imag} */,
  {32'hbe27696a, 32'hbec4d52e} /* (18, 6, 25) {real, imag} */,
  {32'hbd8431c4, 32'h3d0d5e38} /* (18, 6, 24) {real, imag} */,
  {32'h3efc95d0, 32'hbe4ed53d} /* (18, 6, 23) {real, imag} */,
  {32'h3e9a3e71, 32'h3e96a9f1} /* (18, 6, 22) {real, imag} */,
  {32'hbd5d5c6d, 32'hbe1d9944} /* (18, 6, 21) {real, imag} */,
  {32'h3ea85615, 32'h3e15f74e} /* (18, 6, 20) {real, imag} */,
  {32'h3e26c33e, 32'hbdbc9148} /* (18, 6, 19) {real, imag} */,
  {32'hbd34dcfc, 32'h3e5702ce} /* (18, 6, 18) {real, imag} */,
  {32'h3d95121b, 32'hbdbe7b92} /* (18, 6, 17) {real, imag} */,
  {32'h3db8221c, 32'h3e4ca0a8} /* (18, 6, 16) {real, imag} */,
  {32'h3e18106e, 32'h3e7758b0} /* (18, 6, 15) {real, imag} */,
  {32'h3dae67ae, 32'h3daf15df} /* (18, 6, 14) {real, imag} */,
  {32'hbed4feee, 32'h3e33c034} /* (18, 6, 13) {real, imag} */,
  {32'h3e9896b4, 32'h3e1ecee4} /* (18, 6, 12) {real, imag} */,
  {32'hbda43448, 32'hbf1c3c45} /* (18, 6, 11) {real, imag} */,
  {32'hbe2b5943, 32'h3dacfa27} /* (18, 6, 10) {real, imag} */,
  {32'hbd82bc54, 32'h3e816721} /* (18, 6, 9) {real, imag} */,
  {32'hbe9717f0, 32'hbc2e02a0} /* (18, 6, 8) {real, imag} */,
  {32'h3f3f3470, 32'h3e8dacb0} /* (18, 6, 7) {real, imag} */,
  {32'h3e7ec143, 32'hbeb32e32} /* (18, 6, 6) {real, imag} */,
  {32'hbef02ad4, 32'h3e6f7bb1} /* (18, 6, 5) {real, imag} */,
  {32'h3e0373e5, 32'h3d09fb8c} /* (18, 6, 4) {real, imag} */,
  {32'h3e7251d8, 32'h3e921351} /* (18, 6, 3) {real, imag} */,
  {32'h3ea298d6, 32'h3ebc2be4} /* (18, 6, 2) {real, imag} */,
  {32'h3de6e11c, 32'hbe7fd4f3} /* (18, 6, 1) {real, imag} */,
  {32'hbe1ea980, 32'hbe967201} /* (18, 6, 0) {real, imag} */,
  {32'h4029d441, 32'h3f686370} /* (18, 5, 31) {real, imag} */,
  {32'hbfbc1b42, 32'h3efefceb} /* (18, 5, 30) {real, imag} */,
  {32'h3f0f9346, 32'hbdb64c78} /* (18, 5, 29) {real, imag} */,
  {32'hbe3acc79, 32'hbe8a7920} /* (18, 5, 28) {real, imag} */,
  {32'h3dddbc1c, 32'h3e4b5269} /* (18, 5, 27) {real, imag} */,
  {32'hbe2002d5, 32'h3ee68fd7} /* (18, 5, 26) {real, imag} */,
  {32'h3decad1c, 32'h3e9a1fc5} /* (18, 5, 25) {real, imag} */,
  {32'h3c926c1e, 32'hbf11838e} /* (18, 5, 24) {real, imag} */,
  {32'h3eb31538, 32'hbd342315} /* (18, 5, 23) {real, imag} */,
  {32'h3e78e11f, 32'hbe3c4a4f} /* (18, 5, 22) {real, imag} */,
  {32'hbef4a2a4, 32'hbe08ed37} /* (18, 5, 21) {real, imag} */,
  {32'hbeaf27a1, 32'hbdc9164c} /* (18, 5, 20) {real, imag} */,
  {32'hbd92765a, 32'hbcf4d978} /* (18, 5, 19) {real, imag} */,
  {32'hbe2d566b, 32'h3f214a7d} /* (18, 5, 18) {real, imag} */,
  {32'h3cbc89f6, 32'h3edf9d38} /* (18, 5, 17) {real, imag} */,
  {32'h3e515a50, 32'hbde72d15} /* (18, 5, 16) {real, imag} */,
  {32'h3cab2268, 32'hbc72d4d0} /* (18, 5, 15) {real, imag} */,
  {32'h3e235792, 32'h3e692dcb} /* (18, 5, 14) {real, imag} */,
  {32'h3ed6e875, 32'h3e92d87e} /* (18, 5, 13) {real, imag} */,
  {32'h3bc0e900, 32'hbf0f6592} /* (18, 5, 12) {real, imag} */,
  {32'hbe4a4efa, 32'hbf5c728b} /* (18, 5, 11) {real, imag} */,
  {32'h3d91fe8f, 32'hbe23906a} /* (18, 5, 10) {real, imag} */,
  {32'h3b82aa08, 32'hbf3ec104} /* (18, 5, 9) {real, imag} */,
  {32'h3f226e57, 32'h3ed79de6} /* (18, 5, 8) {real, imag} */,
  {32'h3f951339, 32'h3e836c77} /* (18, 5, 7) {real, imag} */,
  {32'hbf2a97f4, 32'hbe922791} /* (18, 5, 6) {real, imag} */,
  {32'hbf585a34, 32'h3e9973f2} /* (18, 5, 5) {real, imag} */,
  {32'hbdf25112, 32'h3f0b0a0d} /* (18, 5, 4) {real, imag} */,
  {32'hbdad2e56, 32'h3e7e8db4} /* (18, 5, 3) {real, imag} */,
  {32'hbf4e6b93, 32'hbfb8f374} /* (18, 5, 2) {real, imag} */,
  {32'h3fe81686, 32'h4010e72e} /* (18, 5, 1) {real, imag} */,
  {32'h3fa6e5e7, 32'h3fc1347b} /* (18, 5, 0) {real, imag} */,
  {32'hbfc84ff7, 32'hc083b242} /* (18, 4, 31) {real, imag} */,
  {32'h3f05754b, 32'h3fe609b9} /* (18, 4, 30) {real, imag} */,
  {32'h3db908ea, 32'hbe5ff103} /* (18, 4, 29) {real, imag} */,
  {32'hbfecaaf3, 32'hbf4335ad} /* (18, 4, 28) {real, imag} */,
  {32'h3f3aaf6e, 32'hbf1bf6e0} /* (18, 4, 27) {real, imag} */,
  {32'hbe5c34f6, 32'h3e88da1c} /* (18, 4, 26) {real, imag} */,
  {32'hbe06c778, 32'h3eaa01ba} /* (18, 4, 25) {real, imag} */,
  {32'h3df4bd7e, 32'hbc648ba8} /* (18, 4, 24) {real, imag} */,
  {32'hbe5f0bd2, 32'h3e670ad4} /* (18, 4, 23) {real, imag} */,
  {32'hbea4f1a0, 32'h3f0bb399} /* (18, 4, 22) {real, imag} */,
  {32'h3bacb390, 32'hbe63109e} /* (18, 4, 21) {real, imag} */,
  {32'h3edac598, 32'h3d00cf73} /* (18, 4, 20) {real, imag} */,
  {32'hbcc49070, 32'h3ebd046b} /* (18, 4, 19) {real, imag} */,
  {32'hbe43cd48, 32'hbeac2125} /* (18, 4, 18) {real, imag} */,
  {32'hbe015f50, 32'hbd6c8440} /* (18, 4, 17) {real, imag} */,
  {32'hbeb37658, 32'hbe2d2a68} /* (18, 4, 16) {real, imag} */,
  {32'h3e370e60, 32'hbd3275e0} /* (18, 4, 15) {real, imag} */,
  {32'h3d881b3e, 32'h3d30f1d0} /* (18, 4, 14) {real, imag} */,
  {32'hbde1f4be, 32'h3ec34b59} /* (18, 4, 13) {real, imag} */,
  {32'h3def3f67, 32'hbf231d7a} /* (18, 4, 12) {real, imag} */,
  {32'h3eac9bbe, 32'hbd3bda16} /* (18, 4, 11) {real, imag} */,
  {32'h3f19d7af, 32'hbf10b966} /* (18, 4, 10) {real, imag} */,
  {32'h3e0f3ca8, 32'hbe5e4f87} /* (18, 4, 9) {real, imag} */,
  {32'h3ea3e1be, 32'h3ecf356b} /* (18, 4, 8) {real, imag} */,
  {32'hbde2813a, 32'hbd8ff1f4} /* (18, 4, 7) {real, imag} */,
  {32'hbe977314, 32'h3f9ae2a6} /* (18, 4, 6) {real, imag} */,
  {32'hbe91795a, 32'h3f63db25} /* (18, 4, 5) {real, imag} */,
  {32'h3f18c316, 32'h3e065ea4} /* (18, 4, 4) {real, imag} */,
  {32'hbd9b8cb8, 32'hbf018fab} /* (18, 4, 3) {real, imag} */,
  {32'h4057928a, 32'h3fe7c8c7} /* (18, 4, 2) {real, imag} */,
  {32'hc07fc6c7, 32'hbfb10953} /* (18, 4, 1) {real, imag} */,
  {32'hc0018090, 32'hbf49ca12} /* (18, 4, 0) {real, imag} */,
  {32'h404a9d42, 32'hc07edc80} /* (18, 3, 31) {real, imag} */,
  {32'hbfee0f18, 32'h40c74fde} /* (18, 3, 30) {real, imag} */,
  {32'hbf8aa8e9, 32'h3ee5ffcf} /* (18, 3, 29) {real, imag} */,
  {32'hbf64befe, 32'hbc205de0} /* (18, 3, 28) {real, imag} */,
  {32'h3f51bb1e, 32'hbf970d95} /* (18, 3, 27) {real, imag} */,
  {32'hbf2ac12a, 32'hbf158560} /* (18, 3, 26) {real, imag} */,
  {32'hbe8b909a, 32'h3f0302ce} /* (18, 3, 25) {real, imag} */,
  {32'h3f2a120c, 32'hbdd93a4e} /* (18, 3, 24) {real, imag} */,
  {32'h3e3d12dc, 32'h3e177c17} /* (18, 3, 23) {real, imag} */,
  {32'hbe1011e6, 32'hbf59080b} /* (18, 3, 22) {real, imag} */,
  {32'h3e225c72, 32'hbf3862d6} /* (18, 3, 21) {real, imag} */,
  {32'hbdc8c2fe, 32'hbed8738c} /* (18, 3, 20) {real, imag} */,
  {32'h3e9cdb5d, 32'hbb319480} /* (18, 3, 19) {real, imag} */,
  {32'h3dc32a18, 32'h3e909a89} /* (18, 3, 18) {real, imag} */,
  {32'h3d4abcba, 32'hbe8934a2} /* (18, 3, 17) {real, imag} */,
  {32'hbdbbc42b, 32'hbdb77460} /* (18, 3, 16) {real, imag} */,
  {32'h3e2d0e2a, 32'h3de96407} /* (18, 3, 15) {real, imag} */,
  {32'hbe7f1c46, 32'h3b1e5300} /* (18, 3, 14) {real, imag} */,
  {32'h3e49e798, 32'hbf0954a7} /* (18, 3, 13) {real, imag} */,
  {32'hbefe97ae, 32'h3d5f5a00} /* (18, 3, 12) {real, imag} */,
  {32'hbe8973dc, 32'hbddd9b4a} /* (18, 3, 11) {real, imag} */,
  {32'h3f00f45e, 32'hbe574fba} /* (18, 3, 10) {real, imag} */,
  {32'h3eb13a2d, 32'hbd852554} /* (18, 3, 9) {real, imag} */,
  {32'hbf1246d0, 32'hbf152422} /* (18, 3, 8) {real, imag} */,
  {32'hbf1fffc0, 32'h3ed67e7a} /* (18, 3, 7) {real, imag} */,
  {32'h3f07f5fd, 32'hbe599b5c} /* (18, 3, 6) {real, imag} */,
  {32'hbdce3ad8, 32'h3d332a90} /* (18, 3, 5) {real, imag} */,
  {32'h3f2ea328, 32'h3f83dfa6} /* (18, 3, 4) {real, imag} */,
  {32'h3f600ead, 32'hbfc026d7} /* (18, 3, 3) {real, imag} */,
  {32'h3fb20704, 32'h4041a831} /* (18, 3, 2) {real, imag} */,
  {32'hc0348fa7, 32'hc0a60828} /* (18, 3, 1) {real, imag} */,
  {32'hbcba5bc0, 32'hbe826d97} /* (18, 3, 0) {real, imag} */,
  {32'h4205513a, 32'hbea712a0} /* (18, 2, 31) {real, imag} */,
  {32'hc1875d3a, 32'h40686d00} /* (18, 2, 30) {real, imag} */,
  {32'h3f8b143d, 32'h3f7e5615} /* (18, 2, 29) {real, imag} */,
  {32'h40115d30, 32'hc0201cde} /* (18, 2, 28) {real, imag} */,
  {32'hbfc9ea44, 32'h3f9c15e2} /* (18, 2, 27) {real, imag} */,
  {32'hbeb30a2d, 32'h3ece353d} /* (18, 2, 26) {real, imag} */,
  {32'h3f21c464, 32'hbf023f05} /* (18, 2, 25) {real, imag} */,
  {32'hbee13b0a, 32'h3ed8ef14} /* (18, 2, 24) {real, imag} */,
  {32'h3e0cdc66, 32'h3d4faa3c} /* (18, 2, 23) {real, imag} */,
  {32'hbd17b9c4, 32'h3e8d62d1} /* (18, 2, 22) {real, imag} */,
  {32'hbda4dd75, 32'h3f32dc6b} /* (18, 2, 21) {real, imag} */,
  {32'h3d1b9b18, 32'hbe868819} /* (18, 2, 20) {real, imag} */,
  {32'hbe946b9f, 32'h3dbd1d20} /* (18, 2, 19) {real, imag} */,
  {32'hbd96983f, 32'h3ed174bd} /* (18, 2, 18) {real, imag} */,
  {32'h3e62e486, 32'hbe087311} /* (18, 2, 17) {real, imag} */,
  {32'hbd710c6a, 32'hbdd3ddd4} /* (18, 2, 16) {real, imag} */,
  {32'h3e54502c, 32'hbe13f18a} /* (18, 2, 15) {real, imag} */,
  {32'hbdb61690, 32'hbdbc9606} /* (18, 2, 14) {real, imag} */,
  {32'h3d30d500, 32'hbe6b0c05} /* (18, 2, 13) {real, imag} */,
  {32'h3e52f316, 32'h3e818188} /* (18, 2, 12) {real, imag} */,
  {32'hbf1b09f2, 32'hbf421458} /* (18, 2, 11) {real, imag} */,
  {32'hbdf8c564, 32'hbdfa6448} /* (18, 2, 10) {real, imag} */,
  {32'h3f0eae98, 32'hbc34d750} /* (18, 2, 9) {real, imag} */,
  {32'hbec253be, 32'hbfa34232} /* (18, 2, 8) {real, imag} */,
  {32'h3f155588, 32'hbe82905a} /* (18, 2, 7) {real, imag} */,
  {32'h3f33f47c, 32'h3f3c609f} /* (18, 2, 6) {real, imag} */,
  {32'hbff9d368, 32'hc02cbb2f} /* (18, 2, 5) {real, imag} */,
  {32'h40476c6e, 32'hbf9b6e10} /* (18, 2, 4) {real, imag} */,
  {32'h3f9f44af, 32'h3f3e5dcc} /* (18, 2, 3) {real, imag} */,
  {32'hc13fb06a, 32'h4060251e} /* (18, 2, 2) {real, imag} */,
  {32'h419ef118, 32'hc0863630} /* (18, 2, 1) {real, imag} */,
  {32'h418dcf57, 32'h40425e41} /* (18, 2, 0) {real, imag} */,
  {32'hc2259ac8, 32'h4116bdb0} /* (18, 1, 31) {real, imag} */,
  {32'h4130f2ea, 32'hbfc8d7d4} /* (18, 1, 30) {real, imag} */,
  {32'hbeabd25c, 32'h3dc813e0} /* (18, 1, 29) {real, imag} */,
  {32'hc01c0b24, 32'hbfe34bbd} /* (18, 1, 28) {real, imag} */,
  {32'h4074b350, 32'hbe988ef4} /* (18, 1, 27) {real, imag} */,
  {32'h3fbf9e19, 32'hbf8297ce} /* (18, 1, 26) {real, imag} */,
  {32'hbeb43e0d, 32'h3f7a1f54} /* (18, 1, 25) {real, imag} */,
  {32'h3eeafe8a, 32'hbef06d21} /* (18, 1, 24) {real, imag} */,
  {32'hbe06d7d4, 32'hbf651a0b} /* (18, 1, 23) {real, imag} */,
  {32'hbd58b9ca, 32'h3eb9152c} /* (18, 1, 22) {real, imag} */,
  {32'h3f5bea6d, 32'hbf3b826a} /* (18, 1, 21) {real, imag} */,
  {32'hbf63cc12, 32'h3e38bb6e} /* (18, 1, 20) {real, imag} */,
  {32'h3f011eda, 32'hbdafd45c} /* (18, 1, 19) {real, imag} */,
  {32'h3e034555, 32'h3d9f2735} /* (18, 1, 18) {real, imag} */,
  {32'h3eb162c4, 32'h3dcf189d} /* (18, 1, 17) {real, imag} */,
  {32'h3e99ee35, 32'h3cd78718} /* (18, 1, 16) {real, imag} */,
  {32'hbea8bc65, 32'hbd9fcaa5} /* (18, 1, 15) {real, imag} */,
  {32'h3dd53931, 32'h3f2eca0a} /* (18, 1, 14) {real, imag} */,
  {32'hbdcd6980, 32'h3dc2d80e} /* (18, 1, 13) {real, imag} */,
  {32'h3efd21e6, 32'h3e2ad8a0} /* (18, 1, 12) {real, imag} */,
  {32'hbe46b422, 32'h3ef97b76} /* (18, 1, 11) {real, imag} */,
  {32'hbdcc2398, 32'h3eac2ff1} /* (18, 1, 10) {real, imag} */,
  {32'h3d77aa80, 32'h3da0195d} /* (18, 1, 9) {real, imag} */,
  {32'h3f559114, 32'h3fa5812a} /* (18, 1, 8) {real, imag} */,
  {32'h3e933642, 32'hbebe826c} /* (18, 1, 7) {real, imag} */,
  {32'h3ebd99f9, 32'hbebb9e74} /* (18, 1, 6) {real, imag} */,
  {32'h3ff0565c, 32'h3fa6304d} /* (18, 1, 5) {real, imag} */,
  {32'hc00ec0fb, 32'hbf73042b} /* (18, 1, 4) {real, imag} */,
  {32'hbe802ec0, 32'hbfb26612} /* (18, 1, 3) {real, imag} */,
  {32'h416a29e0, 32'h41866126} /* (18, 1, 2) {real, imag} */,
  {32'hc26e823b, 32'hc1f00eda} /* (18, 1, 1) {real, imag} */,
  {32'hc24974b6, 32'hc10889b4} /* (18, 1, 0) {real, imag} */,
  {32'hc2197341, 32'h41e2c249} /* (18, 0, 31) {real, imag} */,
  {32'h4084c9ac, 32'hc107f00f} /* (18, 0, 30) {real, imag} */,
  {32'h3f99ebdc, 32'hbf20da9c} /* (18, 0, 29) {real, imag} */,
  {32'h3f10b979, 32'hbf7b6b00} /* (18, 0, 28) {real, imag} */,
  {32'h3f99ae56, 32'h3eec8ae2} /* (18, 0, 27) {real, imag} */,
  {32'h3ed92cee, 32'h3f2169f5} /* (18, 0, 26) {real, imag} */,
  {32'hbdc3118a, 32'h3dfe040c} /* (18, 0, 25) {real, imag} */,
  {32'h3f058355, 32'hbf8d6550} /* (18, 0, 24) {real, imag} */,
  {32'hbe2b37da, 32'hbdcf3dce} /* (18, 0, 23) {real, imag} */,
  {32'h3d29c570, 32'hbe8bfc0a} /* (18, 0, 22) {real, imag} */,
  {32'h3e38d772, 32'hbbaafda0} /* (18, 0, 21) {real, imag} */,
  {32'h3d144520, 32'hbe01e762} /* (18, 0, 20) {real, imag} */,
  {32'h3e8f81ce, 32'h3e15d0fc} /* (18, 0, 19) {real, imag} */,
  {32'hbc87fff0, 32'hbe18d6d0} /* (18, 0, 18) {real, imag} */,
  {32'h3e645abb, 32'h3ea3f8e2} /* (18, 0, 17) {real, imag} */,
  {32'hbd225886, 32'h00000000} /* (18, 0, 16) {real, imag} */,
  {32'h3e645abb, 32'hbea3f8e2} /* (18, 0, 15) {real, imag} */,
  {32'hbc87fff0, 32'h3e18d6d0} /* (18, 0, 14) {real, imag} */,
  {32'h3e8f81ce, 32'hbe15d0fc} /* (18, 0, 13) {real, imag} */,
  {32'h3d144520, 32'h3e01e762} /* (18, 0, 12) {real, imag} */,
  {32'h3e38d772, 32'h3baafda0} /* (18, 0, 11) {real, imag} */,
  {32'h3d29c570, 32'h3e8bfc0a} /* (18, 0, 10) {real, imag} */,
  {32'hbe2b37da, 32'h3dcf3dce} /* (18, 0, 9) {real, imag} */,
  {32'h3f058355, 32'h3f8d6550} /* (18, 0, 8) {real, imag} */,
  {32'hbdc3118a, 32'hbdfe040c} /* (18, 0, 7) {real, imag} */,
  {32'h3ed92cee, 32'hbf2169f5} /* (18, 0, 6) {real, imag} */,
  {32'h3f99ae56, 32'hbeec8ae2} /* (18, 0, 5) {real, imag} */,
  {32'h3f10b979, 32'h3f7b6b00} /* (18, 0, 4) {real, imag} */,
  {32'h3f99ebdc, 32'h3f20da9c} /* (18, 0, 3) {real, imag} */,
  {32'h4084c9ac, 32'h4107f00f} /* (18, 0, 2) {real, imag} */,
  {32'hc2197341, 32'hc1e2c249} /* (18, 0, 1) {real, imag} */,
  {32'hc2563932, 32'h00000000} /* (18, 0, 0) {real, imag} */,
  {32'hc22af334, 32'h41a50cfc} /* (17, 31, 31) {real, imag} */,
  {32'h413119ae, 32'hc15a851f} /* (17, 31, 30) {real, imag} */,
  {32'hbfad1d2b, 32'h3fd736df} /* (17, 31, 29) {real, imag} */,
  {32'hbfad22e4, 32'h3f7e4f6d} /* (17, 31, 28) {real, imag} */,
  {32'h3fef34bc, 32'hbf99facb} /* (17, 31, 27) {real, imag} */,
  {32'h3eaa8dda, 32'h3d908c04} /* (17, 31, 26) {real, imag} */,
  {32'hbe882fea, 32'h3eaa350a} /* (17, 31, 25) {real, imag} */,
  {32'h3f250ad9, 32'hc00df75e} /* (17, 31, 24) {real, imag} */,
  {32'hbdd9dcbc, 32'h3e143fb1} /* (17, 31, 23) {real, imag} */,
  {32'h3e3e94db, 32'h3c99d878} /* (17, 31, 22) {real, imag} */,
  {32'h3cf015e0, 32'hbf525396} /* (17, 31, 21) {real, imag} */,
  {32'h3ee6d210, 32'h3ece21ae} /* (17, 31, 20) {real, imag} */,
  {32'hbf0a5661, 32'h3e2ad338} /* (17, 31, 19) {real, imag} */,
  {32'hbf02c1b2, 32'h3deb45f4} /* (17, 31, 18) {real, imag} */,
  {32'h3eb8029a, 32'hbd31f370} /* (17, 31, 17) {real, imag} */,
  {32'hbe994d8e, 32'h3ea9aef1} /* (17, 31, 16) {real, imag} */,
  {32'h3e3e2cb7, 32'hbf05e109} /* (17, 31, 15) {real, imag} */,
  {32'hbd202454, 32'hbdf379a5} /* (17, 31, 14) {real, imag} */,
  {32'hbd877376, 32'hbd87e550} /* (17, 31, 13) {real, imag} */,
  {32'h3ebb49f7, 32'hbebe1108} /* (17, 31, 12) {real, imag} */,
  {32'hbdbe8df6, 32'h3f126f32} /* (17, 31, 11) {real, imag} */,
  {32'hbdd1f9b6, 32'h3e9254de} /* (17, 31, 10) {real, imag} */,
  {32'hbc0ac650, 32'h3ea6c95f} /* (17, 31, 9) {real, imag} */,
  {32'h3f1f9115, 32'h3f8c2e6e} /* (17, 31, 8) {real, imag} */,
  {32'hbedea69c, 32'hbee6a351} /* (17, 31, 7) {real, imag} */,
  {32'h3fb476a8, 32'hbe7d81b3} /* (17, 31, 6) {real, imag} */,
  {32'h409a21f0, 32'hbec962a4} /* (17, 31, 5) {real, imag} */,
  {32'hbff98756, 32'h400e2986} /* (17, 31, 4) {real, imag} */,
  {32'hbd578d70, 32'hbf29f710} /* (17, 31, 3) {real, imag} */,
  {32'h410723ca, 32'h3fd07471} /* (17, 31, 2) {real, imag} */,
  {32'hc1e325b8, 32'hc0a04e43} /* (17, 31, 1) {real, imag} */,
  {32'hc20ef3c0, 32'h40fde829} /* (17, 31, 0) {real, imag} */,
  {32'h41645dc9, 32'h408390fb} /* (17, 30, 31) {real, imag} */,
  {32'hc10e17b0, 32'hc04cefe8} /* (17, 30, 30) {real, imag} */,
  {32'h3fa4a4b4, 32'h3e43785f} /* (17, 30, 29) {real, imag} */,
  {32'h404df940, 32'h3facdad9} /* (17, 30, 28) {real, imag} */,
  {32'hc02a10a1, 32'h401e6237} /* (17, 30, 27) {real, imag} */,
  {32'hbbe44850, 32'hbf8a2d36} /* (17, 30, 26) {real, imag} */,
  {32'h3d6bc9e9, 32'h3e8136c6} /* (17, 30, 25) {real, imag} */,
  {32'hbea299bb, 32'h3ec456ab} /* (17, 30, 24) {real, imag} */,
  {32'hbe737bc8, 32'hbe5d08d7} /* (17, 30, 23) {real, imag} */,
  {32'h3ea99585, 32'hbe4b4fe4} /* (17, 30, 22) {real, imag} */,
  {32'hbdbd5ae1, 32'h3d5e1358} /* (17, 30, 21) {real, imag} */,
  {32'h3db3c1d0, 32'h3e682340} /* (17, 30, 20) {real, imag} */,
  {32'h3d211f96, 32'h3d835031} /* (17, 30, 19) {real, imag} */,
  {32'hbec5a022, 32'h3e93a118} /* (17, 30, 18) {real, imag} */,
  {32'h3e034f7e, 32'hbe0eedc6} /* (17, 30, 17) {real, imag} */,
  {32'h3e52c800, 32'h3dde694c} /* (17, 30, 16) {real, imag} */,
  {32'h3c97f04c, 32'h3ec619fc} /* (17, 30, 15) {real, imag} */,
  {32'h3e493973, 32'hbea248c7} /* (17, 30, 14) {real, imag} */,
  {32'h3d6dae26, 32'hbdaff8d8} /* (17, 30, 13) {real, imag} */,
  {32'h3c1d8ac0, 32'h3eb2476c} /* (17, 30, 12) {real, imag} */,
  {32'hbe14a283, 32'hbed995c9} /* (17, 30, 11) {real, imag} */,
  {32'hbe19dee0, 32'hbeab02f3} /* (17, 30, 10) {real, imag} */,
  {32'hbe47ef9d, 32'hbe5e6cc8} /* (17, 30, 9) {real, imag} */,
  {32'hbfcba448, 32'hbf286196} /* (17, 30, 8) {real, imag} */,
  {32'h3f828a66, 32'h3ece0f40} /* (17, 30, 7) {real, imag} */,
  {32'hbbaa4e00, 32'h3e8a4aee} /* (17, 30, 6) {real, imag} */,
  {32'hbffacdea, 32'hbfa8e65a} /* (17, 30, 5) {real, imag} */,
  {32'h3f99df6a, 32'h400263c2} /* (17, 30, 4) {real, imag} */,
  {32'h400fef67, 32'hbd801cd8} /* (17, 30, 3) {real, imag} */,
  {32'hc13d1670, 32'hc0234ecf} /* (17, 30, 2) {real, imag} */,
  {32'h41c7915e, 32'hbe99cbf4} /* (17, 30, 1) {real, imag} */,
  {32'h4153456d, 32'hc02fd54d} /* (17, 30, 0) {real, imag} */,
  {32'hbfe54387, 32'h4085d28e} /* (17, 29, 31) {real, imag} */,
  {32'h3fb0f8ea, 32'hc02b433c} /* (17, 29, 30) {real, imag} */,
  {32'h3f350749, 32'h3ff7ab50} /* (17, 29, 29) {real, imag} */,
  {32'h3f41ccfe, 32'hbf930496} /* (17, 29, 28) {real, imag} */,
  {32'hbf24350a, 32'hbf3986f0} /* (17, 29, 27) {real, imag} */,
  {32'h3e72105a, 32'hbec9a48d} /* (17, 29, 26) {real, imag} */,
  {32'hbe8c2bab, 32'hbe4fd531} /* (17, 29, 25) {real, imag} */,
  {32'h3e72efa9, 32'h3e9ce4fc} /* (17, 29, 24) {real, imag} */,
  {32'h3e423098, 32'h3e580a4e} /* (17, 29, 23) {real, imag} */,
  {32'hbdbcd734, 32'hbeae8d2a} /* (17, 29, 22) {real, imag} */,
  {32'h3e8364bd, 32'h3cbcf810} /* (17, 29, 21) {real, imag} */,
  {32'hbe25bd73, 32'h3f0432b4} /* (17, 29, 20) {real, imag} */,
  {32'h3e0c8fbc, 32'h3c8b82b0} /* (17, 29, 19) {real, imag} */,
  {32'h3dd68e6d, 32'h3ab3d740} /* (17, 29, 18) {real, imag} */,
  {32'h3d400922, 32'h3e1ff018} /* (17, 29, 17) {real, imag} */,
  {32'hbeba2fd4, 32'hbe8eb359} /* (17, 29, 16) {real, imag} */,
  {32'h3ea62c02, 32'h3eb7b195} /* (17, 29, 15) {real, imag} */,
  {32'hbf118005, 32'hbea35f08} /* (17, 29, 14) {real, imag} */,
  {32'hbd63a8d2, 32'hbe9d670a} /* (17, 29, 13) {real, imag} */,
  {32'hbe1537ba, 32'hbdb317b0} /* (17, 29, 12) {real, imag} */,
  {32'hbefbe565, 32'hbe8eb270} /* (17, 29, 11) {real, imag} */,
  {32'hbdcbfca9, 32'hbe17cc30} /* (17, 29, 10) {real, imag} */,
  {32'hbee9063c, 32'h3e8bc7a0} /* (17, 29, 9) {real, imag} */,
  {32'hbdc9598c, 32'hbe2b2d17} /* (17, 29, 8) {real, imag} */,
  {32'hbe22b79c, 32'hbf1ba0c9} /* (17, 29, 7) {real, imag} */,
  {32'hbf6db4db, 32'h3e7f7a40} /* (17, 29, 6) {real, imag} */,
  {32'h3fa07314, 32'h3ecb5c9e} /* (17, 29, 5) {real, imag} */,
  {32'hbfa6d3fa, 32'h3f41aa41} /* (17, 29, 4) {real, imag} */,
  {32'h3e8b0521, 32'h3e732a60} /* (17, 29, 3) {real, imag} */,
  {32'hbfb89607, 32'hc098522a} /* (17, 29, 2) {real, imag} */,
  {32'h4080dd57, 32'h403579f5} /* (17, 29, 1) {real, imag} */,
  {32'h3f8341ba, 32'h3e033f42} /* (17, 29, 0) {real, imag} */,
  {32'hc0404ae0, 32'h3f9d6da8} /* (17, 28, 31) {real, imag} */,
  {32'h40229447, 32'hc0239302} /* (17, 28, 30) {real, imag} */,
  {32'hbf5bbaa7, 32'h3f696c84} /* (17, 28, 29) {real, imag} */,
  {32'h3f35a3fe, 32'hbe431bfa} /* (17, 28, 28) {real, imag} */,
  {32'hbf4d42d7, 32'hbf226184} /* (17, 28, 27) {real, imag} */,
  {32'hbd580170, 32'hbf688f71} /* (17, 28, 26) {real, imag} */,
  {32'hbf10ec04, 32'h3f22e694} /* (17, 28, 25) {real, imag} */,
  {32'h3ec98354, 32'h3dcf3887} /* (17, 28, 24) {real, imag} */,
  {32'h3db46804, 32'hbe543eeb} /* (17, 28, 23) {real, imag} */,
  {32'h3eb36582, 32'h3ddea772} /* (17, 28, 22) {real, imag} */,
  {32'h3ea1376b, 32'h3ea198e2} /* (17, 28, 21) {real, imag} */,
  {32'hbe6daac3, 32'h3dd18c38} /* (17, 28, 20) {real, imag} */,
  {32'h3c0c3c60, 32'hbf04eb5d} /* (17, 28, 19) {real, imag} */,
  {32'h3e2066c8, 32'hbc9062b8} /* (17, 28, 18) {real, imag} */,
  {32'h3e25e585, 32'hbe2cc103} /* (17, 28, 17) {real, imag} */,
  {32'h3ec1e00c, 32'hbe802555} /* (17, 28, 16) {real, imag} */,
  {32'hbeb1be4a, 32'h3ea6acea} /* (17, 28, 15) {real, imag} */,
  {32'h3ecba620, 32'h3e2414c0} /* (17, 28, 14) {real, imag} */,
  {32'h3dd6db14, 32'h3dba0161} /* (17, 28, 13) {real, imag} */,
  {32'h3e69525a, 32'h3e0ec5d9} /* (17, 28, 12) {real, imag} */,
  {32'hbd12ed97, 32'hbef4f120} /* (17, 28, 11) {real, imag} */,
  {32'hbdfe56e3, 32'hbecd006c} /* (17, 28, 10) {real, imag} */,
  {32'hbed7e283, 32'hbd06e4ee} /* (17, 28, 9) {real, imag} */,
  {32'h3f67814d, 32'h3f67e69c} /* (17, 28, 8) {real, imag} */,
  {32'h3db9665a, 32'hbe8e25e2} /* (17, 28, 7) {real, imag} */,
  {32'hbef57136, 32'hbe57b64c} /* (17, 28, 6) {real, imag} */,
  {32'h3f1ea620, 32'h3bbb7ad0} /* (17, 28, 5) {real, imag} */,
  {32'hbff15196, 32'h3f527f96} /* (17, 28, 4) {real, imag} */,
  {32'h3ee60558, 32'h3f489c82} /* (17, 28, 3) {real, imag} */,
  {32'h3ecae830, 32'hbfd911df} /* (17, 28, 2) {real, imag} */,
  {32'hbf44f2d4, 32'h405419ba} /* (17, 28, 1) {real, imag} */,
  {32'hc01cbe58, 32'h3ff3c19b} /* (17, 28, 0) {real, imag} */,
  {32'h3fb1115a, 32'hc0215aad} /* (17, 27, 31) {real, imag} */,
  {32'h3e88be06, 32'h3fa2e1ac} /* (17, 27, 30) {real, imag} */,
  {32'hbda52f50, 32'hbed50cb8} /* (17, 27, 29) {real, imag} */,
  {32'hbe35fc26, 32'hbe672f2d} /* (17, 27, 28) {real, imag} */,
  {32'hbf265d44, 32'hbf370752} /* (17, 27, 27) {real, imag} */,
  {32'h3d1257b0, 32'h3f8a1da8} /* (17, 27, 26) {real, imag} */,
  {32'hbf4bb574, 32'hbf5393a4} /* (17, 27, 25) {real, imag} */,
  {32'h3ec7e471, 32'h3ebbc81a} /* (17, 27, 24) {real, imag} */,
  {32'h3f145d6e, 32'h3f014249} /* (17, 27, 23) {real, imag} */,
  {32'h3ede8afb, 32'h3df27918} /* (17, 27, 22) {real, imag} */,
  {32'hbeade120, 32'hbd837aac} /* (17, 27, 21) {real, imag} */,
  {32'hbc85c15a, 32'h3eeacd4c} /* (17, 27, 20) {real, imag} */,
  {32'h3e891c18, 32'hbed8718e} /* (17, 27, 19) {real, imag} */,
  {32'h3e4522ca, 32'hbe174341} /* (17, 27, 18) {real, imag} */,
  {32'h3d9578f2, 32'h3e460530} /* (17, 27, 17) {real, imag} */,
  {32'h3e9e0188, 32'h3de20910} /* (17, 27, 16) {real, imag} */,
  {32'h3d802650, 32'h3e46687d} /* (17, 27, 15) {real, imag} */,
  {32'h3e1ccafe, 32'h3dbc30ce} /* (17, 27, 14) {real, imag} */,
  {32'hbddeed69, 32'h3c99238c} /* (17, 27, 13) {real, imag} */,
  {32'h3ee78729, 32'h3ea76fc6} /* (17, 27, 12) {real, imag} */,
  {32'hbe2357ce, 32'hbe0fc2e4} /* (17, 27, 11) {real, imag} */,
  {32'hbf133d1e, 32'h3ef7daf8} /* (17, 27, 10) {real, imag} */,
  {32'hbce78388, 32'h3e27a49a} /* (17, 27, 9) {real, imag} */,
  {32'hbe7a2238, 32'hbe839ad4} /* (17, 27, 8) {real, imag} */,
  {32'h3e875cea, 32'hbe1e30c0} /* (17, 27, 7) {real, imag} */,
  {32'h3c886558, 32'hbee84462} /* (17, 27, 6) {real, imag} */,
  {32'h3e83344e, 32'hbdaaacb8} /* (17, 27, 5) {real, imag} */,
  {32'hbf0c3c2e, 32'hbe806192} /* (17, 27, 4) {real, imag} */,
  {32'h3e69ee35, 32'hbe1f5d45} /* (17, 27, 3) {real, imag} */,
  {32'hbf9b94ba, 32'h3e184324} /* (17, 27, 2) {real, imag} */,
  {32'h403c336d, 32'hbf7a391f} /* (17, 27, 1) {real, imag} */,
  {32'h3f6caa0f, 32'hbfb53dfb} /* (17, 27, 0) {real, imag} */,
  {32'h3f1c0ad1, 32'h3d4c1b98} /* (17, 26, 31) {real, imag} */,
  {32'h3e5750d2, 32'h3d8beeda} /* (17, 26, 30) {real, imag} */,
  {32'hbef01db7, 32'h3e1f5cb3} /* (17, 26, 29) {real, imag} */,
  {32'h3e8975f8, 32'hbe655a7e} /* (17, 26, 28) {real, imag} */,
  {32'hbc571f40, 32'hbe276230} /* (17, 26, 27) {real, imag} */,
  {32'hbe02fb68, 32'hbd40043c} /* (17, 26, 26) {real, imag} */,
  {32'h3f461766, 32'hbda31105} /* (17, 26, 25) {real, imag} */,
  {32'hbf876142, 32'h3e29f186} /* (17, 26, 24) {real, imag} */,
  {32'h3f143509, 32'h3ed89656} /* (17, 26, 23) {real, imag} */,
  {32'hbf35e78a, 32'h3e6ab484} /* (17, 26, 22) {real, imag} */,
  {32'h3e257003, 32'hbe89045d} /* (17, 26, 21) {real, imag} */,
  {32'h3eac306e, 32'h3e464b40} /* (17, 26, 20) {real, imag} */,
  {32'h3dd797f8, 32'h3eef3ecf} /* (17, 26, 19) {real, imag} */,
  {32'hbd6c8da4, 32'h3f0a70fb} /* (17, 26, 18) {real, imag} */,
  {32'hbeb017bf, 32'h3e56c220} /* (17, 26, 17) {real, imag} */,
  {32'hbc9d27c0, 32'h3e4a5d24} /* (17, 26, 16) {real, imag} */,
  {32'hbcb5d0c0, 32'hbe9a1159} /* (17, 26, 15) {real, imag} */,
  {32'h3e9a0c3a, 32'hbefcdda0} /* (17, 26, 14) {real, imag} */,
  {32'hbdaa7715, 32'h3dfe474b} /* (17, 26, 13) {real, imag} */,
  {32'h3cef84b0, 32'hbd01144f} /* (17, 26, 12) {real, imag} */,
  {32'h3e669aeb, 32'h3d219564} /* (17, 26, 11) {real, imag} */,
  {32'hbeea9c85, 32'hbe9d64d6} /* (17, 26, 10) {real, imag} */,
  {32'h3e989e84, 32'h3e71d3dc} /* (17, 26, 9) {real, imag} */,
  {32'hbebbb20f, 32'h3dd64e42} /* (17, 26, 8) {real, imag} */,
  {32'h3eacca39, 32'hbecb0fe8} /* (17, 26, 7) {real, imag} */,
  {32'h3f0258de, 32'hbda1d861} /* (17, 26, 6) {real, imag} */,
  {32'hbe461f40, 32'h3ecab8e0} /* (17, 26, 5) {real, imag} */,
  {32'hbe09a4bb, 32'hbef99f9f} /* (17, 26, 4) {real, imag} */,
  {32'hbbcafc70, 32'h3f8252a7} /* (17, 26, 3) {real, imag} */,
  {32'hbf40960e, 32'h3e570cfb} /* (17, 26, 2) {real, imag} */,
  {32'h3f547d58, 32'hbe2f9170} /* (17, 26, 1) {real, imag} */,
  {32'hbec8770f, 32'h3e244bb6} /* (17, 26, 0) {real, imag} */,
  {32'hbe221d4c, 32'h3e4ea690} /* (17, 25, 31) {real, imag} */,
  {32'hbe8ebeae, 32'hbe316189} /* (17, 25, 30) {real, imag} */,
  {32'hbed97566, 32'h3c76a980} /* (17, 25, 29) {real, imag} */,
  {32'h3f41ce0c, 32'hbe350339} /* (17, 25, 28) {real, imag} */,
  {32'hbebfece6, 32'h3e8e8190} /* (17, 25, 27) {real, imag} */,
  {32'h3d3bdd50, 32'h3f6220a0} /* (17, 25, 26) {real, imag} */,
  {32'h3dc8af70, 32'hbbef15e0} /* (17, 25, 25) {real, imag} */,
  {32'hbe1af406, 32'h3e968f58} /* (17, 25, 24) {real, imag} */,
  {32'h3df8df06, 32'hbf191d74} /* (17, 25, 23) {real, imag} */,
  {32'hbe58cdf1, 32'h3e54c8af} /* (17, 25, 22) {real, imag} */,
  {32'h3e87033d, 32'h3e1d59a7} /* (17, 25, 21) {real, imag} */,
  {32'h3ce3693f, 32'hbe984337} /* (17, 25, 20) {real, imag} */,
  {32'hbdf2bbff, 32'h3e8825d2} /* (17, 25, 19) {real, imag} */,
  {32'hbeaba945, 32'hbdc3fee1} /* (17, 25, 18) {real, imag} */,
  {32'h3e6334c6, 32'h3c96d614} /* (17, 25, 17) {real, imag} */,
  {32'h3ebb7d54, 32'hbef5c08d} /* (17, 25, 16) {real, imag} */,
  {32'hbe04ceb0, 32'h3ea90fe5} /* (17, 25, 15) {real, imag} */,
  {32'hbbf2a660, 32'h3e9f8c56} /* (17, 25, 14) {real, imag} */,
  {32'h3e34fda5, 32'hbe2c22c6} /* (17, 25, 13) {real, imag} */,
  {32'h3e0c5b15, 32'h3da22e3d} /* (17, 25, 12) {real, imag} */,
  {32'h3efef63c, 32'hbedc15f4} /* (17, 25, 11) {real, imag} */,
  {32'h3f00cf70, 32'hbea0d1c0} /* (17, 25, 10) {real, imag} */,
  {32'hbd38e294, 32'hbec162b1} /* (17, 25, 9) {real, imag} */,
  {32'hbd2d47c4, 32'hbd6c9560} /* (17, 25, 8) {real, imag} */,
  {32'hbd64f840, 32'h3ee8819b} /* (17, 25, 7) {real, imag} */,
  {32'hbf2202aa, 32'h3e0be56c} /* (17, 25, 6) {real, imag} */,
  {32'hbefce140, 32'h3e7574e4} /* (17, 25, 5) {real, imag} */,
  {32'hbe4e81b4, 32'hbf3440e0} /* (17, 25, 4) {real, imag} */,
  {32'hbe01af26, 32'hbdac7d13} /* (17, 25, 3) {real, imag} */,
  {32'h3f928712, 32'h3eb8a2b3} /* (17, 25, 2) {real, imag} */,
  {32'hbe4306d4, 32'hbddd9518} /* (17, 25, 1) {real, imag} */,
  {32'hbea8a444, 32'hbf2dcd86} /* (17, 25, 0) {real, imag} */,
  {32'h3ecdd8a0, 32'hbedcee6c} /* (17, 24, 31) {real, imag} */,
  {32'hbf2a00ee, 32'h3f0a558c} /* (17, 24, 30) {real, imag} */,
  {32'hbe2060ec, 32'hbf4d3f04} /* (17, 24, 29) {real, imag} */,
  {32'h3f8c2766, 32'hbe0dfe6b} /* (17, 24, 28) {real, imag} */,
  {32'hbd584030, 32'hbee69dc0} /* (17, 24, 27) {real, imag} */,
  {32'hbe667990, 32'hbdd67dc8} /* (17, 24, 26) {real, imag} */,
  {32'hbe99ae6f, 32'hbede18c8} /* (17, 24, 25) {real, imag} */,
  {32'h3e3b8bc0, 32'h3efa636e} /* (17, 24, 24) {real, imag} */,
  {32'h3ebb2c56, 32'hbdfca8a8} /* (17, 24, 23) {real, imag} */,
  {32'hbdb0ee0c, 32'hbe2f83d2} /* (17, 24, 22) {real, imag} */,
  {32'h3e82b87e, 32'hbc8a9212} /* (17, 24, 21) {real, imag} */,
  {32'h3f010d72, 32'hbed0abe0} /* (17, 24, 20) {real, imag} */,
  {32'hbe822c74, 32'hbe4fe76a} /* (17, 24, 19) {real, imag} */,
  {32'h3d804c33, 32'h3e93c6d4} /* (17, 24, 18) {real, imag} */,
  {32'hbdec6594, 32'h3af4cac0} /* (17, 24, 17) {real, imag} */,
  {32'h3e9e2791, 32'h3dfbcc8e} /* (17, 24, 16) {real, imag} */,
  {32'hbe0e1725, 32'hbe318f24} /* (17, 24, 15) {real, imag} */,
  {32'h3dc1a8ad, 32'hbe8ea972} /* (17, 24, 14) {real, imag} */,
  {32'hbd16165c, 32'h3d2933ea} /* (17, 24, 13) {real, imag} */,
  {32'h3d93278c, 32'hbe835490} /* (17, 24, 12) {real, imag} */,
  {32'hbea855cd, 32'hbe80491f} /* (17, 24, 11) {real, imag} */,
  {32'hbe099b3c, 32'h3f00d8d6} /* (17, 24, 10) {real, imag} */,
  {32'h3e5ac23a, 32'hbe7c370a} /* (17, 24, 9) {real, imag} */,
  {32'hbf80aa9b, 32'hbe380978} /* (17, 24, 8) {real, imag} */,
  {32'h3e068c50, 32'hbe4993a6} /* (17, 24, 7) {real, imag} */,
  {32'hbea66aad, 32'h3d0f2d20} /* (17, 24, 6) {real, imag} */,
  {32'h3dfdc456, 32'h3e82f736} /* (17, 24, 5) {real, imag} */,
  {32'h3ebbb5cf, 32'hbe079bc4} /* (17, 24, 4) {real, imag} */,
  {32'hbd17a4b8, 32'h3ebf32e1} /* (17, 24, 3) {real, imag} */,
  {32'hbf94bc10, 32'hbf18df3c} /* (17, 24, 2) {real, imag} */,
  {32'h3f8d1468, 32'hbf534360} /* (17, 24, 1) {real, imag} */,
  {32'h3ef73b30, 32'hbe844b34} /* (17, 24, 0) {real, imag} */,
  {32'h3f18da5b, 32'h3fa81a51} /* (17, 23, 31) {real, imag} */,
  {32'hbe0d153b, 32'hbe254723} /* (17, 23, 30) {real, imag} */,
  {32'hbf09cd7c, 32'h3cbd12b8} /* (17, 23, 29) {real, imag} */,
  {32'h3dae1ac0, 32'h3f0eff12} /* (17, 23, 28) {real, imag} */,
  {32'hbec210fb, 32'h3dd85528} /* (17, 23, 27) {real, imag} */,
  {32'hbc8e1b20, 32'hbe6c2828} /* (17, 23, 26) {real, imag} */,
  {32'h3dad7d54, 32'h38e5d000} /* (17, 23, 25) {real, imag} */,
  {32'hbe44eec0, 32'hbe30efe3} /* (17, 23, 24) {real, imag} */,
  {32'h3ef99966, 32'hbd191808} /* (17, 23, 23) {real, imag} */,
  {32'hbe309bec, 32'hbd8d69c6} /* (17, 23, 22) {real, imag} */,
  {32'hbf19ec52, 32'h3e94cfab} /* (17, 23, 21) {real, imag} */,
  {32'hbecce0ae, 32'h3dc0ada8} /* (17, 23, 20) {real, imag} */,
  {32'h3e3d236a, 32'hbf2863c0} /* (17, 23, 19) {real, imag} */,
  {32'h3db88cda, 32'h3ed5a87f} /* (17, 23, 18) {real, imag} */,
  {32'hbdb2a35c, 32'hbf0435f1} /* (17, 23, 17) {real, imag} */,
  {32'hbe1918e8, 32'hbd997d02} /* (17, 23, 16) {real, imag} */,
  {32'hbe719f4c, 32'hbe8ddd42} /* (17, 23, 15) {real, imag} */,
  {32'h3e6d8a8b, 32'h3ed66c2f} /* (17, 23, 14) {real, imag} */,
  {32'hbe92c012, 32'hbe178e79} /* (17, 23, 13) {real, imag} */,
  {32'h3daa86de, 32'h3f2df0fa} /* (17, 23, 12) {real, imag} */,
  {32'h3f16fe56, 32'h3dd33273} /* (17, 23, 11) {real, imag} */,
  {32'hbd013480, 32'h3ef88e89} /* (17, 23, 10) {real, imag} */,
  {32'hbd036b64, 32'hbe8b2c9b} /* (17, 23, 9) {real, imag} */,
  {32'h3eb8baf2, 32'hbf878aeb} /* (17, 23, 8) {real, imag} */,
  {32'hbe73f890, 32'hbe314db8} /* (17, 23, 7) {real, imag} */,
  {32'h3d6b3690, 32'hbf42f3c1} /* (17, 23, 6) {real, imag} */,
  {32'h3e650ac4, 32'hbe4d9ea1} /* (17, 23, 5) {real, imag} */,
  {32'hbefde05c, 32'h3eb6d576} /* (17, 23, 4) {real, imag} */,
  {32'h3e802016, 32'hbe8e551f} /* (17, 23, 3) {real, imag} */,
  {32'hbe4c6edd, 32'hbe2d3992} /* (17, 23, 2) {real, imag} */,
  {32'hbe4ceeb8, 32'h3e2e5b4b} /* (17, 23, 1) {real, imag} */,
  {32'h3eaf1767, 32'hbdd3ac8f} /* (17, 23, 0) {real, imag} */,
  {32'hbf0fa6c2, 32'hbd2cf8a4} /* (17, 22, 31) {real, imag} */,
  {32'h3db88076, 32'hbe2547a2} /* (17, 22, 30) {real, imag} */,
  {32'h3e4b7de6, 32'h3e7b7685} /* (17, 22, 29) {real, imag} */,
  {32'h3d395c30, 32'h3e14ce7c} /* (17, 22, 28) {real, imag} */,
  {32'h3e69b0a4, 32'h3e76a8a3} /* (17, 22, 27) {real, imag} */,
  {32'h3e3aa6a7, 32'hbd8e9be2} /* (17, 22, 26) {real, imag} */,
  {32'hbe4d2042, 32'h3d01d4d8} /* (17, 22, 25) {real, imag} */,
  {32'h3d73ce9b, 32'hbe6be44e} /* (17, 22, 24) {real, imag} */,
  {32'h3e2cb65c, 32'h3e85ca6f} /* (17, 22, 23) {real, imag} */,
  {32'hbe059ff2, 32'hbe4b940c} /* (17, 22, 22) {real, imag} */,
  {32'hbf2f96b2, 32'hbe96a26e} /* (17, 22, 21) {real, imag} */,
  {32'hbea77e70, 32'h3e2db817} /* (17, 22, 20) {real, imag} */,
  {32'hbd291a20, 32'h3e5343b5} /* (17, 22, 19) {real, imag} */,
  {32'hbe55f370, 32'h3d65c40c} /* (17, 22, 18) {real, imag} */,
  {32'hbf011be2, 32'h3d407cd4} /* (17, 22, 17) {real, imag} */,
  {32'h3e6a7ebf, 32'h3e58a490} /* (17, 22, 16) {real, imag} */,
  {32'h3e99d7ec, 32'hbd75f7a1} /* (17, 22, 15) {real, imag} */,
  {32'h3e9cdc65, 32'hbd0a3280} /* (17, 22, 14) {real, imag} */,
  {32'hbd2ad272, 32'h3ce25340} /* (17, 22, 13) {real, imag} */,
  {32'hbd9a3807, 32'h3cb962f0} /* (17, 22, 12) {real, imag} */,
  {32'h3ed8b25c, 32'hbeaf70b3} /* (17, 22, 11) {real, imag} */,
  {32'hbea5bba4, 32'hbedf96c4} /* (17, 22, 10) {real, imag} */,
  {32'hbd8a0ac0, 32'h3d713bf8} /* (17, 22, 9) {real, imag} */,
  {32'h3eaee91c, 32'h3eacaccb} /* (17, 22, 8) {real, imag} */,
  {32'h3c500878, 32'h3deed1b3} /* (17, 22, 7) {real, imag} */,
  {32'h3e8f5a86, 32'hbdd9e5d8} /* (17, 22, 6) {real, imag} */,
  {32'h3e77faf8, 32'h3ec87f2c} /* (17, 22, 5) {real, imag} */,
  {32'hbe4aaec9, 32'hbe32594e} /* (17, 22, 4) {real, imag} */,
  {32'hbdfe838d, 32'h3e0178df} /* (17, 22, 3) {real, imag} */,
  {32'hbd78e098, 32'hbe306d2b} /* (17, 22, 2) {real, imag} */,
  {32'hbe910f01, 32'h3e07f32a} /* (17, 22, 1) {real, imag} */,
  {32'hbd72ea9c, 32'hbeca36b5} /* (17, 22, 0) {real, imag} */,
  {32'hbd72801e, 32'hbed4d49a} /* (17, 21, 31) {real, imag} */,
  {32'h3eb24fb6, 32'h3ef599c8} /* (17, 21, 30) {real, imag} */,
  {32'hbe1f4d2b, 32'hbc632680} /* (17, 21, 29) {real, imag} */,
  {32'hbeb28e41, 32'hbe54dd6a} /* (17, 21, 28) {real, imag} */,
  {32'hbe310a90, 32'h3f1c3618} /* (17, 21, 27) {real, imag} */,
  {32'h3bf82a00, 32'hbf263c00} /* (17, 21, 26) {real, imag} */,
  {32'h3e2d3175, 32'h3eb747b5} /* (17, 21, 25) {real, imag} */,
  {32'hbec47703, 32'h3f10c22a} /* (17, 21, 24) {real, imag} */,
  {32'hbeba246c, 32'hbeaf0e9e} /* (17, 21, 23) {real, imag} */,
  {32'h3f0e55f2, 32'hbc45ab98} /* (17, 21, 22) {real, imag} */,
  {32'hbd8f27de, 32'h3e20fe62} /* (17, 21, 21) {real, imag} */,
  {32'hbe79b023, 32'hbe58a404} /* (17, 21, 20) {real, imag} */,
  {32'h3e0d9400, 32'h3e6268e3} /* (17, 21, 19) {real, imag} */,
  {32'hbcdf3688, 32'h3d8e6000} /* (17, 21, 18) {real, imag} */,
  {32'h3e0bebf4, 32'hbeca09c8} /* (17, 21, 17) {real, imag} */,
  {32'hbe8a8dcb, 32'h3ecd4039} /* (17, 21, 16) {real, imag} */,
  {32'h3d19d877, 32'h3c2dedd0} /* (17, 21, 15) {real, imag} */,
  {32'hbebf9209, 32'h3de6121e} /* (17, 21, 14) {real, imag} */,
  {32'h3cbf65d8, 32'h3e5c9527} /* (17, 21, 13) {real, imag} */,
  {32'hbe54670d, 32'h3d3a9a28} /* (17, 21, 12) {real, imag} */,
  {32'hbf21fd78, 32'h3da264ec} /* (17, 21, 11) {real, imag} */,
  {32'hbe39becc, 32'h3d295646} /* (17, 21, 10) {real, imag} */,
  {32'hbed40c5d, 32'h3ecdecb1} /* (17, 21, 9) {real, imag} */,
  {32'hbf00efde, 32'h3e35cbc5} /* (17, 21, 8) {real, imag} */,
  {32'h3d3d3ca4, 32'h3da0099c} /* (17, 21, 7) {real, imag} */,
  {32'hbea99cd2, 32'hbe527574} /* (17, 21, 6) {real, imag} */,
  {32'hbde02a24, 32'h3f100bb5} /* (17, 21, 5) {real, imag} */,
  {32'h3f2cadd4, 32'hbe689f4e} /* (17, 21, 4) {real, imag} */,
  {32'hbd9afcd4, 32'hbecd3cc9} /* (17, 21, 3) {real, imag} */,
  {32'h3ec9ad6c, 32'h3d481ba4} /* (17, 21, 2) {real, imag} */,
  {32'h3e80dc11, 32'hbf28e124} /* (17, 21, 1) {real, imag} */,
  {32'h3f0f4503, 32'hbede391e} /* (17, 21, 0) {real, imag} */,
  {32'h3e0c9bd3, 32'h3cdabd40} /* (17, 20, 31) {real, imag} */,
  {32'h3ece66cb, 32'h3e4dc575} /* (17, 20, 30) {real, imag} */,
  {32'hbe174c49, 32'hbcc86100} /* (17, 20, 29) {real, imag} */,
  {32'hbed81e80, 32'h3e6a5f77} /* (17, 20, 28) {real, imag} */,
  {32'hbd844804, 32'h3ddc6832} /* (17, 20, 27) {real, imag} */,
  {32'h3e4fcb68, 32'h3e6b6705} /* (17, 20, 26) {real, imag} */,
  {32'hbe2c0e33, 32'h3e0b3d4e} /* (17, 20, 25) {real, imag} */,
  {32'h3f54b99d, 32'h3e91c7c4} /* (17, 20, 24) {real, imag} */,
  {32'hbed15e18, 32'h3e81ad04} /* (17, 20, 23) {real, imag} */,
  {32'hbdf78612, 32'h3e3b4604} /* (17, 20, 22) {real, imag} */,
  {32'h3f2fcb32, 32'hbd8b2c34} /* (17, 20, 21) {real, imag} */,
  {32'hbe17f504, 32'h3e9b02ba} /* (17, 20, 20) {real, imag} */,
  {32'hbdd78119, 32'h3e5a9e42} /* (17, 20, 19) {real, imag} */,
  {32'h3ea050d4, 32'hbe5f58a6} /* (17, 20, 18) {real, imag} */,
  {32'hbe07cd1a, 32'hbd4b69da} /* (17, 20, 17) {real, imag} */,
  {32'hbedb3e13, 32'hbe02220a} /* (17, 20, 16) {real, imag} */,
  {32'hbe73db29, 32'h3d90e2a4} /* (17, 20, 15) {real, imag} */,
  {32'h3e6082ec, 32'h3e0bcb99} /* (17, 20, 14) {real, imag} */,
  {32'h3de33af2, 32'h3d139b08} /* (17, 20, 13) {real, imag} */,
  {32'hbedcae30, 32'hbcf2747c} /* (17, 20, 12) {real, imag} */,
  {32'hbdd35182, 32'h3f3be6aa} /* (17, 20, 11) {real, imag} */,
  {32'h3ee6520b, 32'hbece9606} /* (17, 20, 10) {real, imag} */,
  {32'h3dc5d9b2, 32'h3e96ae00} /* (17, 20, 9) {real, imag} */,
  {32'h3ed816f0, 32'hbec63ce0} /* (17, 20, 8) {real, imag} */,
  {32'hbe698e8f, 32'hbe85bb29} /* (17, 20, 7) {real, imag} */,
  {32'h3ea7604a, 32'hbe8c6d31} /* (17, 20, 6) {real, imag} */,
  {32'h3dc55e1d, 32'h3d895ad8} /* (17, 20, 5) {real, imag} */,
  {32'h3d533122, 32'hbb616880} /* (17, 20, 4) {real, imag} */,
  {32'hbe9b1de2, 32'hbe7b5b28} /* (17, 20, 3) {real, imag} */,
  {32'h3dcad6d8, 32'hbd7ebe30} /* (17, 20, 2) {real, imag} */,
  {32'hbe89324e, 32'h3e059769} /* (17, 20, 1) {real, imag} */,
  {32'hbeeacf5f, 32'h3dea3d4d} /* (17, 20, 0) {real, imag} */,
  {32'hbf3e1052, 32'hbbe17b00} /* (17, 19, 31) {real, imag} */,
  {32'hbe3e6fd4, 32'hbeb4ef6e} /* (17, 19, 30) {real, imag} */,
  {32'h3e3952c8, 32'h3e4ac8fc} /* (17, 19, 29) {real, imag} */,
  {32'h3e4876d9, 32'h3f1909d6} /* (17, 19, 28) {real, imag} */,
  {32'hbeec1018, 32'hbeab8c44} /* (17, 19, 27) {real, imag} */,
  {32'h3efbef96, 32'h3e8d9675} /* (17, 19, 26) {real, imag} */,
  {32'h3d2a3b16, 32'hbe30ba8d} /* (17, 19, 25) {real, imag} */,
  {32'h3e969f2c, 32'hbe7c5f0a} /* (17, 19, 24) {real, imag} */,
  {32'hbea08dab, 32'hbe179400} /* (17, 19, 23) {real, imag} */,
  {32'h3ec313a0, 32'h3c9451d4} /* (17, 19, 22) {real, imag} */,
  {32'hbed633d4, 32'h3f196611} /* (17, 19, 21) {real, imag} */,
  {32'h3e24d978, 32'h3e565c8a} /* (17, 19, 20) {real, imag} */,
  {32'h3e26db87, 32'h3c9d6fe8} /* (17, 19, 19) {real, imag} */,
  {32'hbf4451f6, 32'hbd0267c0} /* (17, 19, 18) {real, imag} */,
  {32'h3ec4cb66, 32'h3e1c3fe5} /* (17, 19, 17) {real, imag} */,
  {32'h3dc0acb6, 32'h3ee645cb} /* (17, 19, 16) {real, imag} */,
  {32'hbc848c84, 32'hbe8f0438} /* (17, 19, 15) {real, imag} */,
  {32'h3e1aab95, 32'hbe56ec5c} /* (17, 19, 14) {real, imag} */,
  {32'hbdaf3610, 32'hbeb68f5e} /* (17, 19, 13) {real, imag} */,
  {32'h3dd196dc, 32'hbdb3c7ee} /* (17, 19, 12) {real, imag} */,
  {32'h3de84efd, 32'hbee70bc3} /* (17, 19, 11) {real, imag} */,
  {32'hbe904ffb, 32'h3e556177} /* (17, 19, 10) {real, imag} */,
  {32'h3e004424, 32'hbe64d601} /* (17, 19, 9) {real, imag} */,
  {32'hbde53648, 32'h3e6cff59} /* (17, 19, 8) {real, imag} */,
  {32'hbcc93148, 32'h3eb218cd} /* (17, 19, 7) {real, imag} */,
  {32'hbe4c7117, 32'h3e918d62} /* (17, 19, 6) {real, imag} */,
  {32'h3ebb7ff4, 32'h3eead9cf} /* (17, 19, 5) {real, imag} */,
  {32'hbea48862, 32'hbe129fc4} /* (17, 19, 4) {real, imag} */,
  {32'hbe2a8b6c, 32'h3e62929f} /* (17, 19, 3) {real, imag} */,
  {32'hbe82c924, 32'h3e612d4e} /* (17, 19, 2) {real, imag} */,
  {32'hbd782350, 32'hbef32dbc} /* (17, 19, 1) {real, imag} */,
  {32'h3e23d74e, 32'h3e582467} /* (17, 19, 0) {real, imag} */,
  {32'h3e6d0667, 32'hbeb0c6c2} /* (17, 18, 31) {real, imag} */,
  {32'h3da79a74, 32'h3cd30870} /* (17, 18, 30) {real, imag} */,
  {32'hbedb4b0b, 32'h3eac01ca} /* (17, 18, 29) {real, imag} */,
  {32'h3eb21590, 32'h3ec48864} /* (17, 18, 28) {real, imag} */,
  {32'h3e2d6630, 32'hbe00be6a} /* (17, 18, 27) {real, imag} */,
  {32'h3dc50325, 32'h3e491538} /* (17, 18, 26) {real, imag} */,
  {32'h3e994eca, 32'h3d2c8d20} /* (17, 18, 25) {real, imag} */,
  {32'h3e717687, 32'h3e4a629f} /* (17, 18, 24) {real, imag} */,
  {32'h3ed4ea1e, 32'h3ebd6ff1} /* (17, 18, 23) {real, imag} */,
  {32'hbef088ef, 32'hbd0cfee0} /* (17, 18, 22) {real, imag} */,
  {32'hbd18b7e4, 32'hbc027688} /* (17, 18, 21) {real, imag} */,
  {32'hbda6fda2, 32'h3db064b0} /* (17, 18, 20) {real, imag} */,
  {32'hbe82173a, 32'hb8a0a000} /* (17, 18, 19) {real, imag} */,
  {32'h3e1ceb31, 32'hbf0bcb12} /* (17, 18, 18) {real, imag} */,
  {32'hbe2dfd30, 32'h3e817bea} /* (17, 18, 17) {real, imag} */,
  {32'h3dc52e56, 32'hbdcdb3ee} /* (17, 18, 16) {real, imag} */,
  {32'h3d87dc44, 32'hbe20e004} /* (17, 18, 15) {real, imag} */,
  {32'h3eb8cbb6, 32'h3b0e5010} /* (17, 18, 14) {real, imag} */,
  {32'hbe7d348f, 32'hbda29696} /* (17, 18, 13) {real, imag} */,
  {32'hbe225da8, 32'hbe926155} /* (17, 18, 12) {real, imag} */,
  {32'hbaf1d3c0, 32'hbddafa8e} /* (17, 18, 11) {real, imag} */,
  {32'hbca58e6c, 32'hbce18e0c} /* (17, 18, 10) {real, imag} */,
  {32'h3ed8cdb4, 32'hbd25252a} /* (17, 18, 9) {real, imag} */,
  {32'hbda29df6, 32'hbd34ba26} /* (17, 18, 8) {real, imag} */,
  {32'hbe87678e, 32'h3a86dc80} /* (17, 18, 7) {real, imag} */,
  {32'h3e979b82, 32'hbe0a4d0d} /* (17, 18, 6) {real, imag} */,
  {32'hbe93475a, 32'h3dea50e3} /* (17, 18, 5) {real, imag} */,
  {32'hbd2c0ee4, 32'hbe3dc1bc} /* (17, 18, 4) {real, imag} */,
  {32'h3f0c9aa0, 32'h3e712a4a} /* (17, 18, 3) {real, imag} */,
  {32'hbe93c92d, 32'hbd3af65a} /* (17, 18, 2) {real, imag} */,
  {32'h3e8cad42, 32'hbddb3113} /* (17, 18, 1) {real, imag} */,
  {32'hbcaf4e0c, 32'hbec22354} /* (17, 18, 0) {real, imag} */,
  {32'hbe3ca8e2, 32'h3e7b5a8a} /* (17, 17, 31) {real, imag} */,
  {32'hbd780b84, 32'h3e8f7e34} /* (17, 17, 30) {real, imag} */,
  {32'h3eaf1d5a, 32'hbdfc75e2} /* (17, 17, 29) {real, imag} */,
  {32'hbe845b82, 32'hbd79c2d8} /* (17, 17, 28) {real, imag} */,
  {32'h3e6e596e, 32'hbd98bfc0} /* (17, 17, 27) {real, imag} */,
  {32'hbe507d69, 32'hbf2b83e0} /* (17, 17, 26) {real, imag} */,
  {32'h3dcd42b7, 32'h3ec68410} /* (17, 17, 25) {real, imag} */,
  {32'hbe5b715d, 32'hbdf1bf78} /* (17, 17, 24) {real, imag} */,
  {32'hbe14baaf, 32'h3ed1ab7b} /* (17, 17, 23) {real, imag} */,
  {32'hbdd449b2, 32'hbd7e1262} /* (17, 17, 22) {real, imag} */,
  {32'hbdc33d74, 32'h3e805223} /* (17, 17, 21) {real, imag} */,
  {32'h3e5c69a2, 32'hbebb82b7} /* (17, 17, 20) {real, imag} */,
  {32'h3ebd5295, 32'hbdca6d2c} /* (17, 17, 19) {real, imag} */,
  {32'h3e319da0, 32'h3e7be7a8} /* (17, 17, 18) {real, imag} */,
  {32'h3e3ac9aa, 32'h3de6cae8} /* (17, 17, 17) {real, imag} */,
  {32'hb9201700, 32'hbe36763c} /* (17, 17, 16) {real, imag} */,
  {32'hbdd8f06e, 32'h3ed25fbe} /* (17, 17, 15) {real, imag} */,
  {32'h3e8ee659, 32'h3c256da0} /* (17, 17, 14) {real, imag} */,
  {32'hbe26f4e4, 32'hbe80ddce} /* (17, 17, 13) {real, imag} */,
  {32'h3f1b78e5, 32'h3d0d6686} /* (17, 17, 12) {real, imag} */,
  {32'hbf01ba7b, 32'h3f02a412} /* (17, 17, 11) {real, imag} */,
  {32'h3d8c9224, 32'hbebc7caa} /* (17, 17, 10) {real, imag} */,
  {32'hbe21f79f, 32'hbe8a9d60} /* (17, 17, 9) {real, imag} */,
  {32'h3ed9017b, 32'hbe001d84} /* (17, 17, 8) {real, imag} */,
  {32'h3e88ab06, 32'h3d1f537c} /* (17, 17, 7) {real, imag} */,
  {32'hbeb4ea22, 32'h3e5cd3b6} /* (17, 17, 6) {real, imag} */,
  {32'h3e8d91c2, 32'hbda50d3a} /* (17, 17, 5) {real, imag} */,
  {32'hbd215940, 32'h3e05a064} /* (17, 17, 4) {real, imag} */,
  {32'hbd40fdb0, 32'hbdb18fbc} /* (17, 17, 3) {real, imag} */,
  {32'hbe885406, 32'hbeb97d34} /* (17, 17, 2) {real, imag} */,
  {32'h3e4ac849, 32'h3ebd4283} /* (17, 17, 1) {real, imag} */,
  {32'h3ec2f7eb, 32'h3d92f6a5} /* (17, 17, 0) {real, imag} */,
  {32'h3e2ed0ab, 32'hbea9c1f9} /* (17, 16, 31) {real, imag} */,
  {32'hbccea908, 32'hbda040ec} /* (17, 16, 30) {real, imag} */,
  {32'hbe05a32c, 32'hbe1ff758} /* (17, 16, 29) {real, imag} */,
  {32'hbb87cbc0, 32'hbeab8cdd} /* (17, 16, 28) {real, imag} */,
  {32'hbdd2e95f, 32'hbe7a5344} /* (17, 16, 27) {real, imag} */,
  {32'h3e4ef036, 32'h3eb5d13c} /* (17, 16, 26) {real, imag} */,
  {32'hbe440955, 32'h3d148c04} /* (17, 16, 25) {real, imag} */,
  {32'h3dcf15af, 32'hbe113aaa} /* (17, 16, 24) {real, imag} */,
  {32'hbe10e126, 32'h3c019e30} /* (17, 16, 23) {real, imag} */,
  {32'h3d7a9095, 32'hbe09bebc} /* (17, 16, 22) {real, imag} */,
  {32'hbda61b84, 32'h3e95ba92} /* (17, 16, 21) {real, imag} */,
  {32'hbb7e10c0, 32'h3ebae6a8} /* (17, 16, 20) {real, imag} */,
  {32'hbe0fc8ee, 32'hbcbecb1c} /* (17, 16, 19) {real, imag} */,
  {32'h3da999f8, 32'hbe53fba1} /* (17, 16, 18) {real, imag} */,
  {32'hbee11614, 32'h3e880314} /* (17, 16, 17) {real, imag} */,
  {32'hbdb4025c, 32'h00000000} /* (17, 16, 16) {real, imag} */,
  {32'hbee11614, 32'hbe880314} /* (17, 16, 15) {real, imag} */,
  {32'h3da999f8, 32'h3e53fba1} /* (17, 16, 14) {real, imag} */,
  {32'hbe0fc8ee, 32'h3cbecb1c} /* (17, 16, 13) {real, imag} */,
  {32'hbb7e10c0, 32'hbebae6a8} /* (17, 16, 12) {real, imag} */,
  {32'hbda61b84, 32'hbe95ba92} /* (17, 16, 11) {real, imag} */,
  {32'h3d7a9095, 32'h3e09bebc} /* (17, 16, 10) {real, imag} */,
  {32'hbe10e126, 32'hbc019e30} /* (17, 16, 9) {real, imag} */,
  {32'h3dcf15af, 32'h3e113aaa} /* (17, 16, 8) {real, imag} */,
  {32'hbe440955, 32'hbd148c04} /* (17, 16, 7) {real, imag} */,
  {32'h3e4ef036, 32'hbeb5d13c} /* (17, 16, 6) {real, imag} */,
  {32'hbdd2e95f, 32'h3e7a5344} /* (17, 16, 5) {real, imag} */,
  {32'hbb87cbc0, 32'h3eab8cdd} /* (17, 16, 4) {real, imag} */,
  {32'hbe05a32c, 32'h3e1ff758} /* (17, 16, 3) {real, imag} */,
  {32'hbccea908, 32'h3da040ec} /* (17, 16, 2) {real, imag} */,
  {32'h3e2ed0ab, 32'h3ea9c1f9} /* (17, 16, 1) {real, imag} */,
  {32'hbe16b4c2, 32'h00000000} /* (17, 16, 0) {real, imag} */,
  {32'h3e4ac849, 32'hbebd4283} /* (17, 15, 31) {real, imag} */,
  {32'hbe885406, 32'h3eb97d34} /* (17, 15, 30) {real, imag} */,
  {32'hbd40fdb0, 32'h3db18fbc} /* (17, 15, 29) {real, imag} */,
  {32'hbd215940, 32'hbe05a064} /* (17, 15, 28) {real, imag} */,
  {32'h3e8d91c2, 32'h3da50d3a} /* (17, 15, 27) {real, imag} */,
  {32'hbeb4ea22, 32'hbe5cd3b6} /* (17, 15, 26) {real, imag} */,
  {32'h3e88ab06, 32'hbd1f537c} /* (17, 15, 25) {real, imag} */,
  {32'h3ed9017b, 32'h3e001d84} /* (17, 15, 24) {real, imag} */,
  {32'hbe21f79f, 32'h3e8a9d60} /* (17, 15, 23) {real, imag} */,
  {32'h3d8c9224, 32'h3ebc7caa} /* (17, 15, 22) {real, imag} */,
  {32'hbf01ba7b, 32'hbf02a412} /* (17, 15, 21) {real, imag} */,
  {32'h3f1b78e5, 32'hbd0d6686} /* (17, 15, 20) {real, imag} */,
  {32'hbe26f4e4, 32'h3e80ddce} /* (17, 15, 19) {real, imag} */,
  {32'h3e8ee659, 32'hbc256da0} /* (17, 15, 18) {real, imag} */,
  {32'hbdd8f06e, 32'hbed25fbe} /* (17, 15, 17) {real, imag} */,
  {32'hb9201700, 32'h3e36763c} /* (17, 15, 16) {real, imag} */,
  {32'h3e3ac9aa, 32'hbde6cae8} /* (17, 15, 15) {real, imag} */,
  {32'h3e319da0, 32'hbe7be7a8} /* (17, 15, 14) {real, imag} */,
  {32'h3ebd5295, 32'h3dca6d2c} /* (17, 15, 13) {real, imag} */,
  {32'h3e5c69a2, 32'h3ebb82b7} /* (17, 15, 12) {real, imag} */,
  {32'hbdc33d74, 32'hbe805223} /* (17, 15, 11) {real, imag} */,
  {32'hbdd449b2, 32'h3d7e1262} /* (17, 15, 10) {real, imag} */,
  {32'hbe14baaf, 32'hbed1ab7b} /* (17, 15, 9) {real, imag} */,
  {32'hbe5b715d, 32'h3df1bf78} /* (17, 15, 8) {real, imag} */,
  {32'h3dcd42b7, 32'hbec68410} /* (17, 15, 7) {real, imag} */,
  {32'hbe507d69, 32'h3f2b83e0} /* (17, 15, 6) {real, imag} */,
  {32'h3e6e596e, 32'h3d98bfc0} /* (17, 15, 5) {real, imag} */,
  {32'hbe845b82, 32'h3d79c2d8} /* (17, 15, 4) {real, imag} */,
  {32'h3eaf1d5a, 32'h3dfc75e2} /* (17, 15, 3) {real, imag} */,
  {32'hbd780b84, 32'hbe8f7e34} /* (17, 15, 2) {real, imag} */,
  {32'hbe3ca8e2, 32'hbe7b5a8a} /* (17, 15, 1) {real, imag} */,
  {32'h3ec2f7eb, 32'hbd92f6a5} /* (17, 15, 0) {real, imag} */,
  {32'h3e8cad42, 32'h3ddb3113} /* (17, 14, 31) {real, imag} */,
  {32'hbe93c92d, 32'h3d3af65a} /* (17, 14, 30) {real, imag} */,
  {32'h3f0c9aa0, 32'hbe712a4a} /* (17, 14, 29) {real, imag} */,
  {32'hbd2c0ee4, 32'h3e3dc1bc} /* (17, 14, 28) {real, imag} */,
  {32'hbe93475a, 32'hbdea50e3} /* (17, 14, 27) {real, imag} */,
  {32'h3e979b82, 32'h3e0a4d0d} /* (17, 14, 26) {real, imag} */,
  {32'hbe87678e, 32'hba86dc80} /* (17, 14, 25) {real, imag} */,
  {32'hbda29df6, 32'h3d34ba26} /* (17, 14, 24) {real, imag} */,
  {32'h3ed8cdb4, 32'h3d25252a} /* (17, 14, 23) {real, imag} */,
  {32'hbca58e6c, 32'h3ce18e0c} /* (17, 14, 22) {real, imag} */,
  {32'hbaf1d3c0, 32'h3ddafa8e} /* (17, 14, 21) {real, imag} */,
  {32'hbe225da8, 32'h3e926155} /* (17, 14, 20) {real, imag} */,
  {32'hbe7d348f, 32'h3da29696} /* (17, 14, 19) {real, imag} */,
  {32'h3eb8cbb6, 32'hbb0e5010} /* (17, 14, 18) {real, imag} */,
  {32'h3d87dc44, 32'h3e20e004} /* (17, 14, 17) {real, imag} */,
  {32'h3dc52e56, 32'h3dcdb3ee} /* (17, 14, 16) {real, imag} */,
  {32'hbe2dfd30, 32'hbe817bea} /* (17, 14, 15) {real, imag} */,
  {32'h3e1ceb31, 32'h3f0bcb12} /* (17, 14, 14) {real, imag} */,
  {32'hbe82173a, 32'h38a0a000} /* (17, 14, 13) {real, imag} */,
  {32'hbda6fda2, 32'hbdb064b0} /* (17, 14, 12) {real, imag} */,
  {32'hbd18b7e4, 32'h3c027688} /* (17, 14, 11) {real, imag} */,
  {32'hbef088ef, 32'h3d0cfee0} /* (17, 14, 10) {real, imag} */,
  {32'h3ed4ea1e, 32'hbebd6ff1} /* (17, 14, 9) {real, imag} */,
  {32'h3e717687, 32'hbe4a629f} /* (17, 14, 8) {real, imag} */,
  {32'h3e994eca, 32'hbd2c8d20} /* (17, 14, 7) {real, imag} */,
  {32'h3dc50325, 32'hbe491538} /* (17, 14, 6) {real, imag} */,
  {32'h3e2d6630, 32'h3e00be6a} /* (17, 14, 5) {real, imag} */,
  {32'h3eb21590, 32'hbec48864} /* (17, 14, 4) {real, imag} */,
  {32'hbedb4b0b, 32'hbeac01ca} /* (17, 14, 3) {real, imag} */,
  {32'h3da79a74, 32'hbcd30870} /* (17, 14, 2) {real, imag} */,
  {32'h3e6d0667, 32'h3eb0c6c2} /* (17, 14, 1) {real, imag} */,
  {32'hbcaf4e0c, 32'h3ec22354} /* (17, 14, 0) {real, imag} */,
  {32'hbd782350, 32'h3ef32dbc} /* (17, 13, 31) {real, imag} */,
  {32'hbe82c924, 32'hbe612d4e} /* (17, 13, 30) {real, imag} */,
  {32'hbe2a8b6c, 32'hbe62929f} /* (17, 13, 29) {real, imag} */,
  {32'hbea48862, 32'h3e129fc4} /* (17, 13, 28) {real, imag} */,
  {32'h3ebb7ff4, 32'hbeead9cf} /* (17, 13, 27) {real, imag} */,
  {32'hbe4c7117, 32'hbe918d62} /* (17, 13, 26) {real, imag} */,
  {32'hbcc93148, 32'hbeb218cd} /* (17, 13, 25) {real, imag} */,
  {32'hbde53648, 32'hbe6cff59} /* (17, 13, 24) {real, imag} */,
  {32'h3e004424, 32'h3e64d601} /* (17, 13, 23) {real, imag} */,
  {32'hbe904ffb, 32'hbe556177} /* (17, 13, 22) {real, imag} */,
  {32'h3de84efd, 32'h3ee70bc3} /* (17, 13, 21) {real, imag} */,
  {32'h3dd196dc, 32'h3db3c7ee} /* (17, 13, 20) {real, imag} */,
  {32'hbdaf3610, 32'h3eb68f5e} /* (17, 13, 19) {real, imag} */,
  {32'h3e1aab95, 32'h3e56ec5c} /* (17, 13, 18) {real, imag} */,
  {32'hbc848c84, 32'h3e8f0438} /* (17, 13, 17) {real, imag} */,
  {32'h3dc0acb6, 32'hbee645cb} /* (17, 13, 16) {real, imag} */,
  {32'h3ec4cb66, 32'hbe1c3fe5} /* (17, 13, 15) {real, imag} */,
  {32'hbf4451f6, 32'h3d0267c0} /* (17, 13, 14) {real, imag} */,
  {32'h3e26db87, 32'hbc9d6fe8} /* (17, 13, 13) {real, imag} */,
  {32'h3e24d978, 32'hbe565c8a} /* (17, 13, 12) {real, imag} */,
  {32'hbed633d4, 32'hbf196611} /* (17, 13, 11) {real, imag} */,
  {32'h3ec313a0, 32'hbc9451d4} /* (17, 13, 10) {real, imag} */,
  {32'hbea08dab, 32'h3e179400} /* (17, 13, 9) {real, imag} */,
  {32'h3e969f2c, 32'h3e7c5f0a} /* (17, 13, 8) {real, imag} */,
  {32'h3d2a3b16, 32'h3e30ba8d} /* (17, 13, 7) {real, imag} */,
  {32'h3efbef96, 32'hbe8d9675} /* (17, 13, 6) {real, imag} */,
  {32'hbeec1018, 32'h3eab8c44} /* (17, 13, 5) {real, imag} */,
  {32'h3e4876d9, 32'hbf1909d6} /* (17, 13, 4) {real, imag} */,
  {32'h3e3952c8, 32'hbe4ac8fc} /* (17, 13, 3) {real, imag} */,
  {32'hbe3e6fd4, 32'h3eb4ef6e} /* (17, 13, 2) {real, imag} */,
  {32'hbf3e1052, 32'h3be17b00} /* (17, 13, 1) {real, imag} */,
  {32'h3e23d74e, 32'hbe582467} /* (17, 13, 0) {real, imag} */,
  {32'hbe89324e, 32'hbe059769} /* (17, 12, 31) {real, imag} */,
  {32'h3dcad6d8, 32'h3d7ebe30} /* (17, 12, 30) {real, imag} */,
  {32'hbe9b1de2, 32'h3e7b5b28} /* (17, 12, 29) {real, imag} */,
  {32'h3d533122, 32'h3b616880} /* (17, 12, 28) {real, imag} */,
  {32'h3dc55e1d, 32'hbd895ad8} /* (17, 12, 27) {real, imag} */,
  {32'h3ea7604a, 32'h3e8c6d31} /* (17, 12, 26) {real, imag} */,
  {32'hbe698e8f, 32'h3e85bb29} /* (17, 12, 25) {real, imag} */,
  {32'h3ed816f0, 32'h3ec63ce0} /* (17, 12, 24) {real, imag} */,
  {32'h3dc5d9b2, 32'hbe96ae00} /* (17, 12, 23) {real, imag} */,
  {32'h3ee6520b, 32'h3ece9606} /* (17, 12, 22) {real, imag} */,
  {32'hbdd35182, 32'hbf3be6aa} /* (17, 12, 21) {real, imag} */,
  {32'hbedcae30, 32'h3cf2747c} /* (17, 12, 20) {real, imag} */,
  {32'h3de33af2, 32'hbd139b08} /* (17, 12, 19) {real, imag} */,
  {32'h3e6082ec, 32'hbe0bcb99} /* (17, 12, 18) {real, imag} */,
  {32'hbe73db29, 32'hbd90e2a4} /* (17, 12, 17) {real, imag} */,
  {32'hbedb3e13, 32'h3e02220a} /* (17, 12, 16) {real, imag} */,
  {32'hbe07cd1a, 32'h3d4b69da} /* (17, 12, 15) {real, imag} */,
  {32'h3ea050d4, 32'h3e5f58a6} /* (17, 12, 14) {real, imag} */,
  {32'hbdd78119, 32'hbe5a9e42} /* (17, 12, 13) {real, imag} */,
  {32'hbe17f504, 32'hbe9b02ba} /* (17, 12, 12) {real, imag} */,
  {32'h3f2fcb32, 32'h3d8b2c34} /* (17, 12, 11) {real, imag} */,
  {32'hbdf78612, 32'hbe3b4604} /* (17, 12, 10) {real, imag} */,
  {32'hbed15e18, 32'hbe81ad04} /* (17, 12, 9) {real, imag} */,
  {32'h3f54b99d, 32'hbe91c7c4} /* (17, 12, 8) {real, imag} */,
  {32'hbe2c0e33, 32'hbe0b3d4e} /* (17, 12, 7) {real, imag} */,
  {32'h3e4fcb68, 32'hbe6b6705} /* (17, 12, 6) {real, imag} */,
  {32'hbd844804, 32'hbddc6832} /* (17, 12, 5) {real, imag} */,
  {32'hbed81e80, 32'hbe6a5f77} /* (17, 12, 4) {real, imag} */,
  {32'hbe174c49, 32'h3cc86100} /* (17, 12, 3) {real, imag} */,
  {32'h3ece66cb, 32'hbe4dc575} /* (17, 12, 2) {real, imag} */,
  {32'h3e0c9bd3, 32'hbcdabd40} /* (17, 12, 1) {real, imag} */,
  {32'hbeeacf5f, 32'hbdea3d4d} /* (17, 12, 0) {real, imag} */,
  {32'h3e80dc11, 32'h3f28e124} /* (17, 11, 31) {real, imag} */,
  {32'h3ec9ad6c, 32'hbd481ba4} /* (17, 11, 30) {real, imag} */,
  {32'hbd9afcd4, 32'h3ecd3cc9} /* (17, 11, 29) {real, imag} */,
  {32'h3f2cadd4, 32'h3e689f4e} /* (17, 11, 28) {real, imag} */,
  {32'hbde02a24, 32'hbf100bb5} /* (17, 11, 27) {real, imag} */,
  {32'hbea99cd2, 32'h3e527574} /* (17, 11, 26) {real, imag} */,
  {32'h3d3d3ca4, 32'hbda0099c} /* (17, 11, 25) {real, imag} */,
  {32'hbf00efde, 32'hbe35cbc5} /* (17, 11, 24) {real, imag} */,
  {32'hbed40c5d, 32'hbecdecb1} /* (17, 11, 23) {real, imag} */,
  {32'hbe39becc, 32'hbd295646} /* (17, 11, 22) {real, imag} */,
  {32'hbf21fd78, 32'hbda264ec} /* (17, 11, 21) {real, imag} */,
  {32'hbe54670d, 32'hbd3a9a28} /* (17, 11, 20) {real, imag} */,
  {32'h3cbf65d8, 32'hbe5c9527} /* (17, 11, 19) {real, imag} */,
  {32'hbebf9209, 32'hbde6121e} /* (17, 11, 18) {real, imag} */,
  {32'h3d19d877, 32'hbc2dedd0} /* (17, 11, 17) {real, imag} */,
  {32'hbe8a8dcb, 32'hbecd4039} /* (17, 11, 16) {real, imag} */,
  {32'h3e0bebf4, 32'h3eca09c8} /* (17, 11, 15) {real, imag} */,
  {32'hbcdf3688, 32'hbd8e6000} /* (17, 11, 14) {real, imag} */,
  {32'h3e0d9400, 32'hbe6268e3} /* (17, 11, 13) {real, imag} */,
  {32'hbe79b023, 32'h3e58a404} /* (17, 11, 12) {real, imag} */,
  {32'hbd8f27de, 32'hbe20fe62} /* (17, 11, 11) {real, imag} */,
  {32'h3f0e55f2, 32'h3c45ab98} /* (17, 11, 10) {real, imag} */,
  {32'hbeba246c, 32'h3eaf0e9e} /* (17, 11, 9) {real, imag} */,
  {32'hbec47703, 32'hbf10c22a} /* (17, 11, 8) {real, imag} */,
  {32'h3e2d3175, 32'hbeb747b5} /* (17, 11, 7) {real, imag} */,
  {32'h3bf82a00, 32'h3f263c00} /* (17, 11, 6) {real, imag} */,
  {32'hbe310a90, 32'hbf1c3618} /* (17, 11, 5) {real, imag} */,
  {32'hbeb28e41, 32'h3e54dd6a} /* (17, 11, 4) {real, imag} */,
  {32'hbe1f4d2b, 32'h3c632680} /* (17, 11, 3) {real, imag} */,
  {32'h3eb24fb6, 32'hbef599c8} /* (17, 11, 2) {real, imag} */,
  {32'hbd72801e, 32'h3ed4d49a} /* (17, 11, 1) {real, imag} */,
  {32'h3f0f4503, 32'h3ede391e} /* (17, 11, 0) {real, imag} */,
  {32'hbe910f01, 32'hbe07f32a} /* (17, 10, 31) {real, imag} */,
  {32'hbd78e098, 32'h3e306d2b} /* (17, 10, 30) {real, imag} */,
  {32'hbdfe838d, 32'hbe0178df} /* (17, 10, 29) {real, imag} */,
  {32'hbe4aaec9, 32'h3e32594e} /* (17, 10, 28) {real, imag} */,
  {32'h3e77faf8, 32'hbec87f2c} /* (17, 10, 27) {real, imag} */,
  {32'h3e8f5a86, 32'h3dd9e5d8} /* (17, 10, 26) {real, imag} */,
  {32'h3c500878, 32'hbdeed1b3} /* (17, 10, 25) {real, imag} */,
  {32'h3eaee91c, 32'hbeacaccb} /* (17, 10, 24) {real, imag} */,
  {32'hbd8a0ac0, 32'hbd713bf8} /* (17, 10, 23) {real, imag} */,
  {32'hbea5bba4, 32'h3edf96c4} /* (17, 10, 22) {real, imag} */,
  {32'h3ed8b25c, 32'h3eaf70b3} /* (17, 10, 21) {real, imag} */,
  {32'hbd9a3807, 32'hbcb962f0} /* (17, 10, 20) {real, imag} */,
  {32'hbd2ad272, 32'hbce25340} /* (17, 10, 19) {real, imag} */,
  {32'h3e9cdc65, 32'h3d0a3280} /* (17, 10, 18) {real, imag} */,
  {32'h3e99d7ec, 32'h3d75f7a1} /* (17, 10, 17) {real, imag} */,
  {32'h3e6a7ebf, 32'hbe58a490} /* (17, 10, 16) {real, imag} */,
  {32'hbf011be2, 32'hbd407cd4} /* (17, 10, 15) {real, imag} */,
  {32'hbe55f370, 32'hbd65c40c} /* (17, 10, 14) {real, imag} */,
  {32'hbd291a20, 32'hbe5343b5} /* (17, 10, 13) {real, imag} */,
  {32'hbea77e70, 32'hbe2db817} /* (17, 10, 12) {real, imag} */,
  {32'hbf2f96b2, 32'h3e96a26e} /* (17, 10, 11) {real, imag} */,
  {32'hbe059ff2, 32'h3e4b940c} /* (17, 10, 10) {real, imag} */,
  {32'h3e2cb65c, 32'hbe85ca6f} /* (17, 10, 9) {real, imag} */,
  {32'h3d73ce9b, 32'h3e6be44e} /* (17, 10, 8) {real, imag} */,
  {32'hbe4d2042, 32'hbd01d4d8} /* (17, 10, 7) {real, imag} */,
  {32'h3e3aa6a7, 32'h3d8e9be2} /* (17, 10, 6) {real, imag} */,
  {32'h3e69b0a4, 32'hbe76a8a3} /* (17, 10, 5) {real, imag} */,
  {32'h3d395c30, 32'hbe14ce7c} /* (17, 10, 4) {real, imag} */,
  {32'h3e4b7de6, 32'hbe7b7685} /* (17, 10, 3) {real, imag} */,
  {32'h3db88076, 32'h3e2547a2} /* (17, 10, 2) {real, imag} */,
  {32'hbf0fa6c2, 32'h3d2cf8a4} /* (17, 10, 1) {real, imag} */,
  {32'hbd72ea9c, 32'h3eca36b5} /* (17, 10, 0) {real, imag} */,
  {32'hbe4ceeb8, 32'hbe2e5b4b} /* (17, 9, 31) {real, imag} */,
  {32'hbe4c6edd, 32'h3e2d3992} /* (17, 9, 30) {real, imag} */,
  {32'h3e802016, 32'h3e8e551f} /* (17, 9, 29) {real, imag} */,
  {32'hbefde05c, 32'hbeb6d576} /* (17, 9, 28) {real, imag} */,
  {32'h3e650ac4, 32'h3e4d9ea1} /* (17, 9, 27) {real, imag} */,
  {32'h3d6b3690, 32'h3f42f3c1} /* (17, 9, 26) {real, imag} */,
  {32'hbe73f890, 32'h3e314db8} /* (17, 9, 25) {real, imag} */,
  {32'h3eb8baf2, 32'h3f878aeb} /* (17, 9, 24) {real, imag} */,
  {32'hbd036b64, 32'h3e8b2c9b} /* (17, 9, 23) {real, imag} */,
  {32'hbd013480, 32'hbef88e89} /* (17, 9, 22) {real, imag} */,
  {32'h3f16fe56, 32'hbdd33273} /* (17, 9, 21) {real, imag} */,
  {32'h3daa86de, 32'hbf2df0fa} /* (17, 9, 20) {real, imag} */,
  {32'hbe92c012, 32'h3e178e79} /* (17, 9, 19) {real, imag} */,
  {32'h3e6d8a8b, 32'hbed66c2f} /* (17, 9, 18) {real, imag} */,
  {32'hbe719f4c, 32'h3e8ddd42} /* (17, 9, 17) {real, imag} */,
  {32'hbe1918e8, 32'h3d997d02} /* (17, 9, 16) {real, imag} */,
  {32'hbdb2a35c, 32'h3f0435f1} /* (17, 9, 15) {real, imag} */,
  {32'h3db88cda, 32'hbed5a87f} /* (17, 9, 14) {real, imag} */,
  {32'h3e3d236a, 32'h3f2863c0} /* (17, 9, 13) {real, imag} */,
  {32'hbecce0ae, 32'hbdc0ada8} /* (17, 9, 12) {real, imag} */,
  {32'hbf19ec52, 32'hbe94cfab} /* (17, 9, 11) {real, imag} */,
  {32'hbe309bec, 32'h3d8d69c6} /* (17, 9, 10) {real, imag} */,
  {32'h3ef99966, 32'h3d191808} /* (17, 9, 9) {real, imag} */,
  {32'hbe44eec0, 32'h3e30efe3} /* (17, 9, 8) {real, imag} */,
  {32'h3dad7d54, 32'hb8e5d000} /* (17, 9, 7) {real, imag} */,
  {32'hbc8e1b20, 32'h3e6c2828} /* (17, 9, 6) {real, imag} */,
  {32'hbec210fb, 32'hbdd85528} /* (17, 9, 5) {real, imag} */,
  {32'h3dae1ac0, 32'hbf0eff12} /* (17, 9, 4) {real, imag} */,
  {32'hbf09cd7c, 32'hbcbd12b8} /* (17, 9, 3) {real, imag} */,
  {32'hbe0d153b, 32'h3e254723} /* (17, 9, 2) {real, imag} */,
  {32'h3f18da5b, 32'hbfa81a51} /* (17, 9, 1) {real, imag} */,
  {32'h3eaf1767, 32'h3dd3ac8f} /* (17, 9, 0) {real, imag} */,
  {32'h3f8d1468, 32'h3f534360} /* (17, 8, 31) {real, imag} */,
  {32'hbf94bc10, 32'h3f18df3c} /* (17, 8, 30) {real, imag} */,
  {32'hbd17a4b8, 32'hbebf32e1} /* (17, 8, 29) {real, imag} */,
  {32'h3ebbb5cf, 32'h3e079bc4} /* (17, 8, 28) {real, imag} */,
  {32'h3dfdc456, 32'hbe82f736} /* (17, 8, 27) {real, imag} */,
  {32'hbea66aad, 32'hbd0f2d20} /* (17, 8, 26) {real, imag} */,
  {32'h3e068c50, 32'h3e4993a6} /* (17, 8, 25) {real, imag} */,
  {32'hbf80aa9b, 32'h3e380978} /* (17, 8, 24) {real, imag} */,
  {32'h3e5ac23a, 32'h3e7c370a} /* (17, 8, 23) {real, imag} */,
  {32'hbe099b3c, 32'hbf00d8d6} /* (17, 8, 22) {real, imag} */,
  {32'hbea855cd, 32'h3e80491f} /* (17, 8, 21) {real, imag} */,
  {32'h3d93278c, 32'h3e835490} /* (17, 8, 20) {real, imag} */,
  {32'hbd16165c, 32'hbd2933ea} /* (17, 8, 19) {real, imag} */,
  {32'h3dc1a8ad, 32'h3e8ea972} /* (17, 8, 18) {real, imag} */,
  {32'hbe0e1725, 32'h3e318f24} /* (17, 8, 17) {real, imag} */,
  {32'h3e9e2791, 32'hbdfbcc8e} /* (17, 8, 16) {real, imag} */,
  {32'hbdec6594, 32'hbaf4cac0} /* (17, 8, 15) {real, imag} */,
  {32'h3d804c33, 32'hbe93c6d4} /* (17, 8, 14) {real, imag} */,
  {32'hbe822c74, 32'h3e4fe76a} /* (17, 8, 13) {real, imag} */,
  {32'h3f010d72, 32'h3ed0abe0} /* (17, 8, 12) {real, imag} */,
  {32'h3e82b87e, 32'h3c8a9212} /* (17, 8, 11) {real, imag} */,
  {32'hbdb0ee0c, 32'h3e2f83d2} /* (17, 8, 10) {real, imag} */,
  {32'h3ebb2c56, 32'h3dfca8a8} /* (17, 8, 9) {real, imag} */,
  {32'h3e3b8bc0, 32'hbefa636e} /* (17, 8, 8) {real, imag} */,
  {32'hbe99ae6f, 32'h3ede18c8} /* (17, 8, 7) {real, imag} */,
  {32'hbe667990, 32'h3dd67dc8} /* (17, 8, 6) {real, imag} */,
  {32'hbd584030, 32'h3ee69dc0} /* (17, 8, 5) {real, imag} */,
  {32'h3f8c2766, 32'h3e0dfe6b} /* (17, 8, 4) {real, imag} */,
  {32'hbe2060ec, 32'h3f4d3f04} /* (17, 8, 3) {real, imag} */,
  {32'hbf2a00ee, 32'hbf0a558c} /* (17, 8, 2) {real, imag} */,
  {32'h3ecdd8a0, 32'h3edcee6c} /* (17, 8, 1) {real, imag} */,
  {32'h3ef73b30, 32'h3e844b34} /* (17, 8, 0) {real, imag} */,
  {32'hbe4306d4, 32'h3ddd9518} /* (17, 7, 31) {real, imag} */,
  {32'h3f928712, 32'hbeb8a2b3} /* (17, 7, 30) {real, imag} */,
  {32'hbe01af26, 32'h3dac7d13} /* (17, 7, 29) {real, imag} */,
  {32'hbe4e81b4, 32'h3f3440e0} /* (17, 7, 28) {real, imag} */,
  {32'hbefce140, 32'hbe7574e4} /* (17, 7, 27) {real, imag} */,
  {32'hbf2202aa, 32'hbe0be56c} /* (17, 7, 26) {real, imag} */,
  {32'hbd64f840, 32'hbee8819b} /* (17, 7, 25) {real, imag} */,
  {32'hbd2d47c4, 32'h3d6c9560} /* (17, 7, 24) {real, imag} */,
  {32'hbd38e294, 32'h3ec162b1} /* (17, 7, 23) {real, imag} */,
  {32'h3f00cf70, 32'h3ea0d1c0} /* (17, 7, 22) {real, imag} */,
  {32'h3efef63c, 32'h3edc15f4} /* (17, 7, 21) {real, imag} */,
  {32'h3e0c5b15, 32'hbda22e3d} /* (17, 7, 20) {real, imag} */,
  {32'h3e34fda5, 32'h3e2c22c6} /* (17, 7, 19) {real, imag} */,
  {32'hbbf2a660, 32'hbe9f8c56} /* (17, 7, 18) {real, imag} */,
  {32'hbe04ceb0, 32'hbea90fe5} /* (17, 7, 17) {real, imag} */,
  {32'h3ebb7d54, 32'h3ef5c08d} /* (17, 7, 16) {real, imag} */,
  {32'h3e6334c6, 32'hbc96d614} /* (17, 7, 15) {real, imag} */,
  {32'hbeaba945, 32'h3dc3fee1} /* (17, 7, 14) {real, imag} */,
  {32'hbdf2bbff, 32'hbe8825d2} /* (17, 7, 13) {real, imag} */,
  {32'h3ce3693f, 32'h3e984337} /* (17, 7, 12) {real, imag} */,
  {32'h3e87033d, 32'hbe1d59a7} /* (17, 7, 11) {real, imag} */,
  {32'hbe58cdf1, 32'hbe54c8af} /* (17, 7, 10) {real, imag} */,
  {32'h3df8df06, 32'h3f191d74} /* (17, 7, 9) {real, imag} */,
  {32'hbe1af406, 32'hbe968f58} /* (17, 7, 8) {real, imag} */,
  {32'h3dc8af70, 32'h3bef15e0} /* (17, 7, 7) {real, imag} */,
  {32'h3d3bdd50, 32'hbf6220a0} /* (17, 7, 6) {real, imag} */,
  {32'hbebfece6, 32'hbe8e8190} /* (17, 7, 5) {real, imag} */,
  {32'h3f41ce0c, 32'h3e350339} /* (17, 7, 4) {real, imag} */,
  {32'hbed97566, 32'hbc76a980} /* (17, 7, 3) {real, imag} */,
  {32'hbe8ebeae, 32'h3e316189} /* (17, 7, 2) {real, imag} */,
  {32'hbe221d4c, 32'hbe4ea690} /* (17, 7, 1) {real, imag} */,
  {32'hbea8a444, 32'h3f2dcd86} /* (17, 7, 0) {real, imag} */,
  {32'h3f547d58, 32'h3e2f9170} /* (17, 6, 31) {real, imag} */,
  {32'hbf40960e, 32'hbe570cfb} /* (17, 6, 30) {real, imag} */,
  {32'hbbcafc70, 32'hbf8252a7} /* (17, 6, 29) {real, imag} */,
  {32'hbe09a4bb, 32'h3ef99f9f} /* (17, 6, 28) {real, imag} */,
  {32'hbe461f40, 32'hbecab8e0} /* (17, 6, 27) {real, imag} */,
  {32'h3f0258de, 32'h3da1d861} /* (17, 6, 26) {real, imag} */,
  {32'h3eacca39, 32'h3ecb0fe8} /* (17, 6, 25) {real, imag} */,
  {32'hbebbb20f, 32'hbdd64e42} /* (17, 6, 24) {real, imag} */,
  {32'h3e989e84, 32'hbe71d3dc} /* (17, 6, 23) {real, imag} */,
  {32'hbeea9c85, 32'h3e9d64d6} /* (17, 6, 22) {real, imag} */,
  {32'h3e669aeb, 32'hbd219564} /* (17, 6, 21) {real, imag} */,
  {32'h3cef84b0, 32'h3d01144f} /* (17, 6, 20) {real, imag} */,
  {32'hbdaa7715, 32'hbdfe474b} /* (17, 6, 19) {real, imag} */,
  {32'h3e9a0c3a, 32'h3efcdda0} /* (17, 6, 18) {real, imag} */,
  {32'hbcb5d0c0, 32'h3e9a1159} /* (17, 6, 17) {real, imag} */,
  {32'hbc9d27c0, 32'hbe4a5d24} /* (17, 6, 16) {real, imag} */,
  {32'hbeb017bf, 32'hbe56c220} /* (17, 6, 15) {real, imag} */,
  {32'hbd6c8da4, 32'hbf0a70fb} /* (17, 6, 14) {real, imag} */,
  {32'h3dd797f8, 32'hbeef3ecf} /* (17, 6, 13) {real, imag} */,
  {32'h3eac306e, 32'hbe464b40} /* (17, 6, 12) {real, imag} */,
  {32'h3e257003, 32'h3e89045d} /* (17, 6, 11) {real, imag} */,
  {32'hbf35e78a, 32'hbe6ab484} /* (17, 6, 10) {real, imag} */,
  {32'h3f143509, 32'hbed89656} /* (17, 6, 9) {real, imag} */,
  {32'hbf876142, 32'hbe29f186} /* (17, 6, 8) {real, imag} */,
  {32'h3f461766, 32'h3da31105} /* (17, 6, 7) {real, imag} */,
  {32'hbe02fb68, 32'h3d40043c} /* (17, 6, 6) {real, imag} */,
  {32'hbc571f40, 32'h3e276230} /* (17, 6, 5) {real, imag} */,
  {32'h3e8975f8, 32'h3e655a7e} /* (17, 6, 4) {real, imag} */,
  {32'hbef01db7, 32'hbe1f5cb3} /* (17, 6, 3) {real, imag} */,
  {32'h3e5750d2, 32'hbd8beeda} /* (17, 6, 2) {real, imag} */,
  {32'h3f1c0ad1, 32'hbd4c1b98} /* (17, 6, 1) {real, imag} */,
  {32'hbec8770f, 32'hbe244bb6} /* (17, 6, 0) {real, imag} */,
  {32'h403c336d, 32'h3f7a391f} /* (17, 5, 31) {real, imag} */,
  {32'hbf9b94ba, 32'hbe184324} /* (17, 5, 30) {real, imag} */,
  {32'h3e69ee35, 32'h3e1f5d45} /* (17, 5, 29) {real, imag} */,
  {32'hbf0c3c2e, 32'h3e806192} /* (17, 5, 28) {real, imag} */,
  {32'h3e83344e, 32'h3daaacb8} /* (17, 5, 27) {real, imag} */,
  {32'h3c886558, 32'h3ee84462} /* (17, 5, 26) {real, imag} */,
  {32'h3e875cea, 32'h3e1e30c0} /* (17, 5, 25) {real, imag} */,
  {32'hbe7a2238, 32'h3e839ad4} /* (17, 5, 24) {real, imag} */,
  {32'hbce78388, 32'hbe27a49a} /* (17, 5, 23) {real, imag} */,
  {32'hbf133d1e, 32'hbef7daf8} /* (17, 5, 22) {real, imag} */,
  {32'hbe2357ce, 32'h3e0fc2e4} /* (17, 5, 21) {real, imag} */,
  {32'h3ee78729, 32'hbea76fc6} /* (17, 5, 20) {real, imag} */,
  {32'hbddeed69, 32'hbc99238c} /* (17, 5, 19) {real, imag} */,
  {32'h3e1ccafe, 32'hbdbc30ce} /* (17, 5, 18) {real, imag} */,
  {32'h3d802650, 32'hbe46687d} /* (17, 5, 17) {real, imag} */,
  {32'h3e9e0188, 32'hbde20910} /* (17, 5, 16) {real, imag} */,
  {32'h3d9578f2, 32'hbe460530} /* (17, 5, 15) {real, imag} */,
  {32'h3e4522ca, 32'h3e174341} /* (17, 5, 14) {real, imag} */,
  {32'h3e891c18, 32'h3ed8718e} /* (17, 5, 13) {real, imag} */,
  {32'hbc85c15a, 32'hbeeacd4c} /* (17, 5, 12) {real, imag} */,
  {32'hbeade120, 32'h3d837aac} /* (17, 5, 11) {real, imag} */,
  {32'h3ede8afb, 32'hbdf27918} /* (17, 5, 10) {real, imag} */,
  {32'h3f145d6e, 32'hbf014249} /* (17, 5, 9) {real, imag} */,
  {32'h3ec7e471, 32'hbebbc81a} /* (17, 5, 8) {real, imag} */,
  {32'hbf4bb574, 32'h3f5393a4} /* (17, 5, 7) {real, imag} */,
  {32'h3d1257b0, 32'hbf8a1da8} /* (17, 5, 6) {real, imag} */,
  {32'hbf265d44, 32'h3f370752} /* (17, 5, 5) {real, imag} */,
  {32'hbe35fc26, 32'h3e672f2d} /* (17, 5, 4) {real, imag} */,
  {32'hbda52f50, 32'h3ed50cb8} /* (17, 5, 3) {real, imag} */,
  {32'h3e88be06, 32'hbfa2e1ac} /* (17, 5, 2) {real, imag} */,
  {32'h3fb1115a, 32'h40215aad} /* (17, 5, 1) {real, imag} */,
  {32'h3f6caa0f, 32'h3fb53dfb} /* (17, 5, 0) {real, imag} */,
  {32'hbf44f2d4, 32'hc05419ba} /* (17, 4, 31) {real, imag} */,
  {32'h3ecae830, 32'h3fd911df} /* (17, 4, 30) {real, imag} */,
  {32'h3ee60558, 32'hbf489c82} /* (17, 4, 29) {real, imag} */,
  {32'hbff15196, 32'hbf527f96} /* (17, 4, 28) {real, imag} */,
  {32'h3f1ea620, 32'hbbbb7ad0} /* (17, 4, 27) {real, imag} */,
  {32'hbef57136, 32'h3e57b64c} /* (17, 4, 26) {real, imag} */,
  {32'h3db9665a, 32'h3e8e25e2} /* (17, 4, 25) {real, imag} */,
  {32'h3f67814d, 32'hbf67e69c} /* (17, 4, 24) {real, imag} */,
  {32'hbed7e283, 32'h3d06e4ee} /* (17, 4, 23) {real, imag} */,
  {32'hbdfe56e3, 32'h3ecd006c} /* (17, 4, 22) {real, imag} */,
  {32'hbd12ed97, 32'h3ef4f120} /* (17, 4, 21) {real, imag} */,
  {32'h3e69525a, 32'hbe0ec5d9} /* (17, 4, 20) {real, imag} */,
  {32'h3dd6db14, 32'hbdba0161} /* (17, 4, 19) {real, imag} */,
  {32'h3ecba620, 32'hbe2414c0} /* (17, 4, 18) {real, imag} */,
  {32'hbeb1be4a, 32'hbea6acea} /* (17, 4, 17) {real, imag} */,
  {32'h3ec1e00c, 32'h3e802555} /* (17, 4, 16) {real, imag} */,
  {32'h3e25e585, 32'h3e2cc103} /* (17, 4, 15) {real, imag} */,
  {32'h3e2066c8, 32'h3c9062b8} /* (17, 4, 14) {real, imag} */,
  {32'h3c0c3c60, 32'h3f04eb5d} /* (17, 4, 13) {real, imag} */,
  {32'hbe6daac3, 32'hbdd18c38} /* (17, 4, 12) {real, imag} */,
  {32'h3ea1376b, 32'hbea198e2} /* (17, 4, 11) {real, imag} */,
  {32'h3eb36582, 32'hbddea772} /* (17, 4, 10) {real, imag} */,
  {32'h3db46804, 32'h3e543eeb} /* (17, 4, 9) {real, imag} */,
  {32'h3ec98354, 32'hbdcf3887} /* (17, 4, 8) {real, imag} */,
  {32'hbf10ec04, 32'hbf22e694} /* (17, 4, 7) {real, imag} */,
  {32'hbd580170, 32'h3f688f71} /* (17, 4, 6) {real, imag} */,
  {32'hbf4d42d7, 32'h3f226184} /* (17, 4, 5) {real, imag} */,
  {32'h3f35a3fe, 32'h3e431bfa} /* (17, 4, 4) {real, imag} */,
  {32'hbf5bbaa7, 32'hbf696c84} /* (17, 4, 3) {real, imag} */,
  {32'h40229447, 32'h40239302} /* (17, 4, 2) {real, imag} */,
  {32'hc0404ae0, 32'hbf9d6da8} /* (17, 4, 1) {real, imag} */,
  {32'hc01cbe58, 32'hbff3c19b} /* (17, 4, 0) {real, imag} */,
  {32'h4080dd57, 32'hc03579f5} /* (17, 3, 31) {real, imag} */,
  {32'hbfb89607, 32'h4098522a} /* (17, 3, 30) {real, imag} */,
  {32'h3e8b0521, 32'hbe732a60} /* (17, 3, 29) {real, imag} */,
  {32'hbfa6d3fa, 32'hbf41aa41} /* (17, 3, 28) {real, imag} */,
  {32'h3fa07314, 32'hbecb5c9e} /* (17, 3, 27) {real, imag} */,
  {32'hbf6db4db, 32'hbe7f7a40} /* (17, 3, 26) {real, imag} */,
  {32'hbe22b79c, 32'h3f1ba0c9} /* (17, 3, 25) {real, imag} */,
  {32'hbdc9598c, 32'h3e2b2d17} /* (17, 3, 24) {real, imag} */,
  {32'hbee9063c, 32'hbe8bc7a0} /* (17, 3, 23) {real, imag} */,
  {32'hbdcbfca9, 32'h3e17cc30} /* (17, 3, 22) {real, imag} */,
  {32'hbefbe565, 32'h3e8eb270} /* (17, 3, 21) {real, imag} */,
  {32'hbe1537ba, 32'h3db317b0} /* (17, 3, 20) {real, imag} */,
  {32'hbd63a8d2, 32'h3e9d670a} /* (17, 3, 19) {real, imag} */,
  {32'hbf118005, 32'h3ea35f08} /* (17, 3, 18) {real, imag} */,
  {32'h3ea62c02, 32'hbeb7b195} /* (17, 3, 17) {real, imag} */,
  {32'hbeba2fd4, 32'h3e8eb359} /* (17, 3, 16) {real, imag} */,
  {32'h3d400922, 32'hbe1ff018} /* (17, 3, 15) {real, imag} */,
  {32'h3dd68e6d, 32'hbab3d740} /* (17, 3, 14) {real, imag} */,
  {32'h3e0c8fbc, 32'hbc8b82b0} /* (17, 3, 13) {real, imag} */,
  {32'hbe25bd73, 32'hbf0432b4} /* (17, 3, 12) {real, imag} */,
  {32'h3e8364bd, 32'hbcbcf810} /* (17, 3, 11) {real, imag} */,
  {32'hbdbcd734, 32'h3eae8d2a} /* (17, 3, 10) {real, imag} */,
  {32'h3e423098, 32'hbe580a4e} /* (17, 3, 9) {real, imag} */,
  {32'h3e72efa9, 32'hbe9ce4fc} /* (17, 3, 8) {real, imag} */,
  {32'hbe8c2bab, 32'h3e4fd531} /* (17, 3, 7) {real, imag} */,
  {32'h3e72105a, 32'h3ec9a48d} /* (17, 3, 6) {real, imag} */,
  {32'hbf24350a, 32'h3f3986f0} /* (17, 3, 5) {real, imag} */,
  {32'h3f41ccfe, 32'h3f930496} /* (17, 3, 4) {real, imag} */,
  {32'h3f350749, 32'hbff7ab50} /* (17, 3, 3) {real, imag} */,
  {32'h3fb0f8ea, 32'h402b433c} /* (17, 3, 2) {real, imag} */,
  {32'hbfe54387, 32'hc085d28e} /* (17, 3, 1) {real, imag} */,
  {32'h3f8341ba, 32'hbe033f42} /* (17, 3, 0) {real, imag} */,
  {32'h41c7915e, 32'h3e99cbf4} /* (17, 2, 31) {real, imag} */,
  {32'hc13d1670, 32'h40234ecf} /* (17, 2, 30) {real, imag} */,
  {32'h400fef67, 32'h3d801cd8} /* (17, 2, 29) {real, imag} */,
  {32'h3f99df6a, 32'hc00263c2} /* (17, 2, 28) {real, imag} */,
  {32'hbffacdea, 32'h3fa8e65a} /* (17, 2, 27) {real, imag} */,
  {32'hbbaa4e00, 32'hbe8a4aee} /* (17, 2, 26) {real, imag} */,
  {32'h3f828a66, 32'hbece0f40} /* (17, 2, 25) {real, imag} */,
  {32'hbfcba448, 32'h3f286196} /* (17, 2, 24) {real, imag} */,
  {32'hbe47ef9d, 32'h3e5e6cc8} /* (17, 2, 23) {real, imag} */,
  {32'hbe19dee0, 32'h3eab02f3} /* (17, 2, 22) {real, imag} */,
  {32'hbe14a283, 32'h3ed995c9} /* (17, 2, 21) {real, imag} */,
  {32'h3c1d8ac0, 32'hbeb2476c} /* (17, 2, 20) {real, imag} */,
  {32'h3d6dae26, 32'h3daff8d8} /* (17, 2, 19) {real, imag} */,
  {32'h3e493973, 32'h3ea248c7} /* (17, 2, 18) {real, imag} */,
  {32'h3c97f04c, 32'hbec619fc} /* (17, 2, 17) {real, imag} */,
  {32'h3e52c800, 32'hbdde694c} /* (17, 2, 16) {real, imag} */,
  {32'h3e034f7e, 32'h3e0eedc6} /* (17, 2, 15) {real, imag} */,
  {32'hbec5a022, 32'hbe93a118} /* (17, 2, 14) {real, imag} */,
  {32'h3d211f96, 32'hbd835031} /* (17, 2, 13) {real, imag} */,
  {32'h3db3c1d0, 32'hbe682340} /* (17, 2, 12) {real, imag} */,
  {32'hbdbd5ae1, 32'hbd5e1358} /* (17, 2, 11) {real, imag} */,
  {32'h3ea99585, 32'h3e4b4fe4} /* (17, 2, 10) {real, imag} */,
  {32'hbe737bc8, 32'h3e5d08d7} /* (17, 2, 9) {real, imag} */,
  {32'hbea299bb, 32'hbec456ab} /* (17, 2, 8) {real, imag} */,
  {32'h3d6bc9e9, 32'hbe8136c6} /* (17, 2, 7) {real, imag} */,
  {32'hbbe44850, 32'h3f8a2d36} /* (17, 2, 6) {real, imag} */,
  {32'hc02a10a1, 32'hc01e6237} /* (17, 2, 5) {real, imag} */,
  {32'h404df940, 32'hbfacdad9} /* (17, 2, 4) {real, imag} */,
  {32'h3fa4a4b4, 32'hbe43785f} /* (17, 2, 3) {real, imag} */,
  {32'hc10e17b0, 32'h404cefe8} /* (17, 2, 2) {real, imag} */,
  {32'h41645dc9, 32'hc08390fb} /* (17, 2, 1) {real, imag} */,
  {32'h4153456d, 32'h402fd54d} /* (17, 2, 0) {real, imag} */,
  {32'hc1e325b8, 32'h40a04e43} /* (17, 1, 31) {real, imag} */,
  {32'h410723ca, 32'hbfd07471} /* (17, 1, 30) {real, imag} */,
  {32'hbd578d70, 32'h3f29f710} /* (17, 1, 29) {real, imag} */,
  {32'hbff98756, 32'hc00e2986} /* (17, 1, 28) {real, imag} */,
  {32'h409a21f0, 32'h3ec962a4} /* (17, 1, 27) {real, imag} */,
  {32'h3fb476a8, 32'h3e7d81b3} /* (17, 1, 26) {real, imag} */,
  {32'hbedea69c, 32'h3ee6a351} /* (17, 1, 25) {real, imag} */,
  {32'h3f1f9115, 32'hbf8c2e6e} /* (17, 1, 24) {real, imag} */,
  {32'hbc0ac650, 32'hbea6c95f} /* (17, 1, 23) {real, imag} */,
  {32'hbdd1f9b6, 32'hbe9254de} /* (17, 1, 22) {real, imag} */,
  {32'hbdbe8df6, 32'hbf126f32} /* (17, 1, 21) {real, imag} */,
  {32'h3ebb49f7, 32'h3ebe1108} /* (17, 1, 20) {real, imag} */,
  {32'hbd877376, 32'h3d87e550} /* (17, 1, 19) {real, imag} */,
  {32'hbd202454, 32'h3df379a5} /* (17, 1, 18) {real, imag} */,
  {32'h3e3e2cb7, 32'h3f05e109} /* (17, 1, 17) {real, imag} */,
  {32'hbe994d8e, 32'hbea9aef1} /* (17, 1, 16) {real, imag} */,
  {32'h3eb8029a, 32'h3d31f370} /* (17, 1, 15) {real, imag} */,
  {32'hbf02c1b2, 32'hbdeb45f4} /* (17, 1, 14) {real, imag} */,
  {32'hbf0a5661, 32'hbe2ad338} /* (17, 1, 13) {real, imag} */,
  {32'h3ee6d210, 32'hbece21ae} /* (17, 1, 12) {real, imag} */,
  {32'h3cf015e0, 32'h3f525396} /* (17, 1, 11) {real, imag} */,
  {32'h3e3e94db, 32'hbc99d878} /* (17, 1, 10) {real, imag} */,
  {32'hbdd9dcbc, 32'hbe143fb1} /* (17, 1, 9) {real, imag} */,
  {32'h3f250ad9, 32'h400df75e} /* (17, 1, 8) {real, imag} */,
  {32'hbe882fea, 32'hbeaa350a} /* (17, 1, 7) {real, imag} */,
  {32'h3eaa8dda, 32'hbd908c04} /* (17, 1, 6) {real, imag} */,
  {32'h3fef34bc, 32'h3f99facb} /* (17, 1, 5) {real, imag} */,
  {32'hbfad22e4, 32'hbf7e4f6d} /* (17, 1, 4) {real, imag} */,
  {32'hbfad1d2b, 32'hbfd736df} /* (17, 1, 3) {real, imag} */,
  {32'h413119ae, 32'h415a851f} /* (17, 1, 2) {real, imag} */,
  {32'hc22af334, 32'hc1a50cfc} /* (17, 1, 1) {real, imag} */,
  {32'hc20ef3c0, 32'hc0fde829} /* (17, 1, 0) {real, imag} */,
  {32'hc1e71599, 32'h41a2213a} /* (17, 0, 31) {real, imag} */,
  {32'h4025bd79, 32'hc0e3558b} /* (17, 0, 30) {real, imag} */,
  {32'h3ff1d857, 32'h3f652f40} /* (17, 0, 29) {real, imag} */,
  {32'h3e93d84e, 32'hbf48ef74} /* (17, 0, 28) {real, imag} */,
  {32'h3f74c91c, 32'h3fab5e56} /* (17, 0, 27) {real, imag} */,
  {32'h3d793b08, 32'hbe595845} /* (17, 0, 26) {real, imag} */,
  {32'hbe7aba63, 32'h3efda962} /* (17, 0, 25) {real, imag} */,
  {32'h3f7c9351, 32'hbebbb64e} /* (17, 0, 24) {real, imag} */,
  {32'h3e2a1894, 32'hbeee5358} /* (17, 0, 23) {real, imag} */,
  {32'h3e42ac6e, 32'h3e0ee08e} /* (17, 0, 22) {real, imag} */,
  {32'h3f0b1072, 32'hbf30c811} /* (17, 0, 21) {real, imag} */,
  {32'h3d9fcefa, 32'h3e1b7fb2} /* (17, 0, 20) {real, imag} */,
  {32'h3e97bee2, 32'h3ea95176} /* (17, 0, 19) {real, imag} */,
  {32'hbea8fa80, 32'hbe6c2939} /* (17, 0, 18) {real, imag} */,
  {32'hbdb3dc7f, 32'h3e84f2a3} /* (17, 0, 17) {real, imag} */,
  {32'hbec448a2, 32'h00000000} /* (17, 0, 16) {real, imag} */,
  {32'hbdb3dc7f, 32'hbe84f2a3} /* (17, 0, 15) {real, imag} */,
  {32'hbea8fa80, 32'h3e6c2939} /* (17, 0, 14) {real, imag} */,
  {32'h3e97bee2, 32'hbea95176} /* (17, 0, 13) {real, imag} */,
  {32'h3d9fcefa, 32'hbe1b7fb2} /* (17, 0, 12) {real, imag} */,
  {32'h3f0b1072, 32'h3f30c811} /* (17, 0, 11) {real, imag} */,
  {32'h3e42ac6e, 32'hbe0ee08e} /* (17, 0, 10) {real, imag} */,
  {32'h3e2a1894, 32'h3eee5358} /* (17, 0, 9) {real, imag} */,
  {32'h3f7c9351, 32'h3ebbb64e} /* (17, 0, 8) {real, imag} */,
  {32'hbe7aba63, 32'hbefda962} /* (17, 0, 7) {real, imag} */,
  {32'h3d793b08, 32'h3e595845} /* (17, 0, 6) {real, imag} */,
  {32'h3f74c91c, 32'hbfab5e56} /* (17, 0, 5) {real, imag} */,
  {32'h3e93d84e, 32'h3f48ef74} /* (17, 0, 4) {real, imag} */,
  {32'h3ff1d857, 32'hbf652f40} /* (17, 0, 3) {real, imag} */,
  {32'h4025bd79, 32'h40e3558b} /* (17, 0, 2) {real, imag} */,
  {32'hc1e71599, 32'hc1a2213a} /* (17, 0, 1) {real, imag} */,
  {32'hc20c0ae0, 32'h00000000} /* (17, 0, 0) {real, imag} */,
  {32'hc196a040, 32'h40f0ba5d} /* (16, 31, 31) {real, imag} */,
  {32'h40803086, 32'hc0d42f73} /* (16, 31, 30) {real, imag} */,
  {32'hbf7ee1ff, 32'hbeba5880} /* (16, 31, 29) {real, imag} */,
  {32'hbfba5c66, 32'h3ea49777} /* (16, 31, 28) {real, imag} */,
  {32'h3ff660e2, 32'hbf7518ce} /* (16, 31, 27) {real, imag} */,
  {32'hbe10c21a, 32'hbf1679ee} /* (16, 31, 26) {real, imag} */,
  {32'hbd8f8e26, 32'h3f20ac28} /* (16, 31, 25) {real, imag} */,
  {32'h3e7e7128, 32'hbf3d5189} /* (16, 31, 24) {real, imag} */,
  {32'h3e928433, 32'hbe7fd64c} /* (16, 31, 23) {real, imag} */,
  {32'h3e078c98, 32'hbde1d634} /* (16, 31, 22) {real, imag} */,
  {32'h3df54fc6, 32'hbf4f6f50} /* (16, 31, 21) {real, imag} */,
  {32'hbe8bd5c4, 32'h3f2a38c2} /* (16, 31, 20) {real, imag} */,
  {32'h3c3a93a8, 32'hbdd7d8c8} /* (16, 31, 19) {real, imag} */,
  {32'hbcac29cc, 32'hbe64d42a} /* (16, 31, 18) {real, imag} */,
  {32'hbcb8b92c, 32'hbe152676} /* (16, 31, 17) {real, imag} */,
  {32'hbe443076, 32'hbeb151b0} /* (16, 31, 16) {real, imag} */,
  {32'hbebd88f8, 32'h3de59aef} /* (16, 31, 15) {real, imag} */,
  {32'h3d8488e8, 32'hbe44c194} /* (16, 31, 14) {real, imag} */,
  {32'h3bd71d80, 32'hbed0cc18} /* (16, 31, 13) {real, imag} */,
  {32'h3e4597a8, 32'h3ec96438} /* (16, 31, 12) {real, imag} */,
  {32'hbd005608, 32'h3f304976} /* (16, 31, 11) {real, imag} */,
  {32'hbe15f084, 32'hbe565155} /* (16, 31, 10) {real, imag} */,
  {32'hbec7fb94, 32'hbee1bd66} /* (16, 31, 9) {real, imag} */,
  {32'hbc1a22b0, 32'h3ecca71f} /* (16, 31, 8) {real, imag} */,
  {32'hbea2288c, 32'hbeb17902} /* (16, 31, 7) {real, imag} */,
  {32'h3f9fb484, 32'h3cbe6d20} /* (16, 31, 6) {real, imag} */,
  {32'h402c0bc7, 32'h3def9e22} /* (16, 31, 5) {real, imag} */,
  {32'hbf67daa7, 32'h3fffb5b5} /* (16, 31, 4) {real, imag} */,
  {32'hbe262fb2, 32'hbf961134} /* (16, 31, 3) {real, imag} */,
  {32'h404eb9cb, 32'h3fad3df8} /* (16, 31, 2) {real, imag} */,
  {32'hc129e471, 32'hbf77d62e} /* (16, 31, 1) {real, imag} */,
  {32'hc15bf39e, 32'h40d6e162} /* (16, 31, 0) {real, imag} */,
  {32'h40d25d58, 32'h40074e32} /* (16, 30, 31) {real, imag} */,
  {32'hc0935ae8, 32'hbfd57096} /* (16, 30, 30) {real, imag} */,
  {32'h3fce23a5, 32'h3f88953e} /* (16, 30, 29) {real, imag} */,
  {32'h400cd20f, 32'h3ffba005} /* (16, 30, 28) {real, imag} */,
  {32'hbfa7d671, 32'h3f85cc47} /* (16, 30, 27) {real, imag} */,
  {32'h3ec60f24, 32'hbf886788} /* (16, 30, 26) {real, imag} */,
  {32'h3e815ed4, 32'h3f28dbae} /* (16, 30, 25) {real, imag} */,
  {32'hbd089ec0, 32'h3f1e9816} /* (16, 30, 24) {real, imag} */,
  {32'hbeb75fee, 32'hbec13fc8} /* (16, 30, 23) {real, imag} */,
  {32'hbe69d6d9, 32'hbe9f7780} /* (16, 30, 22) {real, imag} */,
  {32'h3cece7e8, 32'h3eb3794e} /* (16, 30, 21) {real, imag} */,
  {32'hbf32f796, 32'hbe8b6330} /* (16, 30, 20) {real, imag} */,
  {32'h3e083189, 32'hbea95024} /* (16, 30, 19) {real, imag} */,
  {32'hbe80a7b6, 32'h3eb63e1f} /* (16, 30, 18) {real, imag} */,
  {32'hbec2b1cf, 32'hbdaeceec} /* (16, 30, 17) {real, imag} */,
  {32'hbdb2db5d, 32'hbe2ae302} /* (16, 30, 16) {real, imag} */,
  {32'hbe854dc6, 32'h3dcb1777} /* (16, 30, 15) {real, imag} */,
  {32'hbda9ca0b, 32'h3c43d998} /* (16, 30, 14) {real, imag} */,
  {32'hbeb4a8cc, 32'h3cb6c77e} /* (16, 30, 13) {real, imag} */,
  {32'h3e36fcaa, 32'h3e07d80a} /* (16, 30, 12) {real, imag} */,
  {32'h3b824e20, 32'hbf40d919} /* (16, 30, 11) {real, imag} */,
  {32'hbdcedfa3, 32'h3e4a6495} /* (16, 30, 10) {real, imag} */,
  {32'hbecc89d3, 32'hbf0cc3a5} /* (16, 30, 9) {real, imag} */,
  {32'hbf885792, 32'hbed66ed8} /* (16, 30, 8) {real, imag} */,
  {32'h3f535b7e, 32'h3f944c77} /* (16, 30, 7) {real, imag} */,
  {32'h3e0f1896, 32'hbee4c2ed} /* (16, 30, 6) {real, imag} */,
  {32'hbf7d5c0e, 32'hbf16de1c} /* (16, 30, 5) {real, imag} */,
  {32'h3f453ad6, 32'h3f3337ce} /* (16, 30, 4) {real, imag} */,
  {32'h4010f9ee, 32'hbf26bee2} /* (16, 30, 3) {real, imag} */,
  {32'hc0ab9d67, 32'hbf96c7cd} /* (16, 30, 2) {real, imag} */,
  {32'h4135b55c, 32'h3f882d55} /* (16, 30, 1) {real, imag} */,
  {32'h40a463d3, 32'hc009471a} /* (16, 30, 0) {real, imag} */,
  {32'hbf826ac2, 32'h4023f852} /* (16, 29, 31) {real, imag} */,
  {32'h40171188, 32'hbf96f3d0} /* (16, 29, 30) {real, imag} */,
  {32'h3e8cfc1b, 32'h3efdfa0d} /* (16, 29, 29) {real, imag} */,
  {32'h3f10803e, 32'hbf1d0864} /* (16, 29, 28) {real, imag} */,
  {32'hbf0e1e02, 32'hbe802733} /* (16, 29, 27) {real, imag} */,
  {32'hbf0005d0, 32'hbe0311c2} /* (16, 29, 26) {real, imag} */,
  {32'hbe50444c, 32'h3e9b23b6} /* (16, 29, 25) {real, imag} */,
  {32'h3d82eb04, 32'h3f0226a3} /* (16, 29, 24) {real, imag} */,
  {32'hbf0f8df1, 32'hbe687389} /* (16, 29, 23) {real, imag} */,
  {32'h3c6acb50, 32'h3f08e3c5} /* (16, 29, 22) {real, imag} */,
  {32'h3ee7c226, 32'h3e1fbefd} /* (16, 29, 21) {real, imag} */,
  {32'hbeb16220, 32'h3e7ecc8b} /* (16, 29, 20) {real, imag} */,
  {32'hbecd823d, 32'h3e3a483a} /* (16, 29, 19) {real, imag} */,
  {32'h3ecd49bd, 32'h3d7c036a} /* (16, 29, 18) {real, imag} */,
  {32'h3ec8a698, 32'hbeaf8729} /* (16, 29, 17) {real, imag} */,
  {32'h3e14aec2, 32'hbe5777d5} /* (16, 29, 16) {real, imag} */,
  {32'hbe1ac3ce, 32'h3db295e6} /* (16, 29, 15) {real, imag} */,
  {32'hbcb5b548, 32'h3e323e14} /* (16, 29, 14) {real, imag} */,
  {32'hbd7f8368, 32'h3e81c5aa} /* (16, 29, 13) {real, imag} */,
  {32'hbc218910, 32'hbdeab9b7} /* (16, 29, 12) {real, imag} */,
  {32'h3ed02bdd, 32'hbd1431be} /* (16, 29, 11) {real, imag} */,
  {32'h3c16ec70, 32'h3e40ba5d} /* (16, 29, 10) {real, imag} */,
  {32'hbed12ec5, 32'hbd978b56} /* (16, 29, 9) {real, imag} */,
  {32'hbe5cea7a, 32'h3d758794} /* (16, 29, 8) {real, imag} */,
  {32'hbf3aa252, 32'hbf2bb9e5} /* (16, 29, 7) {real, imag} */,
  {32'hbd988f58, 32'hbd2196b6} /* (16, 29, 6) {real, imag} */,
  {32'h3ee191b8, 32'hbde68ad4} /* (16, 29, 5) {real, imag} */,
  {32'hbec6e227, 32'hbd3f4d74} /* (16, 29, 4) {real, imag} */,
  {32'hbf48b58a, 32'hbf179098} /* (16, 29, 3) {real, imag} */,
  {32'h3f2b2c82, 32'hc0246962} /* (16, 29, 2) {real, imag} */,
  {32'h4055e0dc, 32'h3fd0b5ec} /* (16, 29, 1) {real, imag} */,
  {32'h3f105f7a, 32'hbf24b14b} /* (16, 29, 0) {real, imag} */,
  {32'hbf8ce2be, 32'h3f95a388} /* (16, 28, 31) {real, imag} */,
  {32'h3f976092, 32'hbff8c2f9} /* (16, 28, 30) {real, imag} */,
  {32'hbefd33a6, 32'h3e0b24d8} /* (16, 28, 29) {real, imag} */,
  {32'hbe83fc49, 32'h3f57fa27} /* (16, 28, 28) {real, imag} */,
  {32'hbf0aae12, 32'hbe8239a2} /* (16, 28, 27) {real, imag} */,
  {32'hbea3d011, 32'h3ea4bb9c} /* (16, 28, 26) {real, imag} */,
  {32'hbf5b095a, 32'h3e160a48} /* (16, 28, 25) {real, imag} */,
  {32'h3f11f692, 32'hbead68be} /* (16, 28, 24) {real, imag} */,
  {32'hbe9930da, 32'hbf01ad64} /* (16, 28, 23) {real, imag} */,
  {32'h3f238449, 32'hbd894c7c} /* (16, 28, 22) {real, imag} */,
  {32'hbe4b16fe, 32'h3e9ec8b7} /* (16, 28, 21) {real, imag} */,
  {32'h3df07691, 32'hbd8a6a56} /* (16, 28, 20) {real, imag} */,
  {32'hbecb4da3, 32'hbe85ef57} /* (16, 28, 19) {real, imag} */,
  {32'hbe241c75, 32'hbe4e2ff2} /* (16, 28, 18) {real, imag} */,
  {32'h3e946a74, 32'h3dca939e} /* (16, 28, 17) {real, imag} */,
  {32'hbe1e3c68, 32'h3e1ae6a6} /* (16, 28, 16) {real, imag} */,
  {32'hbe8576e6, 32'hbd0c59a6} /* (16, 28, 15) {real, imag} */,
  {32'h3e12e2e9, 32'hbda7d58e} /* (16, 28, 14) {real, imag} */,
  {32'h3d24c4b0, 32'hbde4b6d6} /* (16, 28, 13) {real, imag} */,
  {32'hbd853f98, 32'hbe4c0c12} /* (16, 28, 12) {real, imag} */,
  {32'hbce4ad36, 32'h3e3aa582} /* (16, 28, 11) {real, imag} */,
  {32'h3de1fc82, 32'hbe05ff20} /* (16, 28, 10) {real, imag} */,
  {32'h3dacfae6, 32'hbce9bf10} /* (16, 28, 9) {real, imag} */,
  {32'h3f899a8e, 32'h3f38d4ff} /* (16, 28, 8) {real, imag} */,
  {32'hbf1cb690, 32'hbab17400} /* (16, 28, 7) {real, imag} */,
  {32'hbea59ff8, 32'hbe0d4d5f} /* (16, 28, 6) {real, imag} */,
  {32'h3f14e39b, 32'hbe289d65} /* (16, 28, 5) {real, imag} */,
  {32'hbf9c27aa, 32'hbe7c8e5e} /* (16, 28, 4) {real, imag} */,
  {32'hbda0bf02, 32'h3f9ae6e1} /* (16, 28, 3) {real, imag} */,
  {32'h3f8f346b, 32'hbf47f420} /* (16, 28, 2) {real, imag} */,
  {32'hbe7ef748, 32'h400e53ee} /* (16, 28, 1) {real, imag} */,
  {32'hc00acaa1, 32'h4016486a} /* (16, 28, 0) {real, imag} */,
  {32'h3f20dc8e, 32'hbfdc1706} /* (16, 27, 31) {real, imag} */,
  {32'hbdc6f4b8, 32'h3fb66d87} /* (16, 27, 30) {real, imag} */,
  {32'hbea489dd, 32'h3d324d8c} /* (16, 27, 29) {real, imag} */,
  {32'h3ed4b8f5, 32'hbce32e98} /* (16, 27, 28) {real, imag} */,
  {32'hbf600008, 32'hbf5cbb5b} /* (16, 27, 27) {real, imag} */,
  {32'hbdcf8582, 32'hbe4f2bf4} /* (16, 27, 26) {real, imag} */,
  {32'hbd1854b8, 32'hbf06caac} /* (16, 27, 25) {real, imag} */,
  {32'h3e4e175e, 32'hbe9a4fe6} /* (16, 27, 24) {real, imag} */,
  {32'hbef8c88c, 32'hbd9e1b2a} /* (16, 27, 23) {real, imag} */,
  {32'hbe841c64, 32'h3f4378ea} /* (16, 27, 22) {real, imag} */,
  {32'h3f0f13c0, 32'hbe818f4d} /* (16, 27, 21) {real, imag} */,
  {32'h3eee77ad, 32'hbe98a145} /* (16, 27, 20) {real, imag} */,
  {32'hbd851cda, 32'h3dea0f04} /* (16, 27, 19) {real, imag} */,
  {32'h3e893b1a, 32'h3deac28b} /* (16, 27, 18) {real, imag} */,
  {32'hbe9c228f, 32'hbeabbf3b} /* (16, 27, 17) {real, imag} */,
  {32'hbeae3380, 32'hbe8d46b1} /* (16, 27, 16) {real, imag} */,
  {32'h3d484a76, 32'hbd00c8e1} /* (16, 27, 15) {real, imag} */,
  {32'h3daf3984, 32'h3d2b52b8} /* (16, 27, 14) {real, imag} */,
  {32'h3bfdb080, 32'h3eb0760e} /* (16, 27, 13) {real, imag} */,
  {32'hbeab2d92, 32'hbd0b64e0} /* (16, 27, 12) {real, imag} */,
  {32'hbe0bab9e, 32'h3e514531} /* (16, 27, 11) {real, imag} */,
  {32'h3c9b9680, 32'hbebb0653} /* (16, 27, 10) {real, imag} */,
  {32'hbe83a542, 32'hbd58a9e8} /* (16, 27, 9) {real, imag} */,
  {32'hbf394790, 32'hbec29a9f} /* (16, 27, 8) {real, imag} */,
  {32'hbe54e649, 32'h3e434098} /* (16, 27, 7) {real, imag} */,
  {32'hbde144db, 32'hbf05ebf2} /* (16, 27, 6) {real, imag} */,
  {32'h3dddb322, 32'hbf26a638} /* (16, 27, 5) {real, imag} */,
  {32'h3d9dce72, 32'hbedb7df2} /* (16, 27, 4) {real, imag} */,
  {32'h3eb18f0c, 32'hbf52cc37} /* (16, 27, 3) {real, imag} */,
  {32'hbf5de820, 32'h3f5ae196} /* (16, 27, 2) {real, imag} */,
  {32'h3fd146f0, 32'hbf6ab79a} /* (16, 27, 1) {real, imag} */,
  {32'h3eb619bc, 32'hbfa4ad66} /* (16, 27, 0) {real, imag} */,
  {32'h3f1c7b22, 32'hbdbcc0b0} /* (16, 26, 31) {real, imag} */,
  {32'h3ec9149e, 32'h3dfbba58} /* (16, 26, 30) {real, imag} */,
  {32'h3e160241, 32'hbe6e1746} /* (16, 26, 29) {real, imag} */,
  {32'h3d2327c0, 32'hbf30f047} /* (16, 26, 28) {real, imag} */,
  {32'hbdb50853, 32'h3e1c36f4} /* (16, 26, 27) {real, imag} */,
  {32'h3df8c06a, 32'hbb89c6b0} /* (16, 26, 26) {real, imag} */,
  {32'h3f2f4862, 32'hbd6719f8} /* (16, 26, 25) {real, imag} */,
  {32'hbd91c108, 32'h3f003afc} /* (16, 26, 24) {real, imag} */,
  {32'h3bac44e0, 32'h3d2d4c3c} /* (16, 26, 23) {real, imag} */,
  {32'hbf248c5d, 32'hbdadc1ac} /* (16, 26, 22) {real, imag} */,
  {32'hbeddf51b, 32'hbe98e706} /* (16, 26, 21) {real, imag} */,
  {32'h3ec3dae3, 32'h3c315270} /* (16, 26, 20) {real, imag} */,
  {32'h3ebacf5e, 32'h3f043cfb} /* (16, 26, 19) {real, imag} */,
  {32'h3ecf250a, 32'hbe2e7ffe} /* (16, 26, 18) {real, imag} */,
  {32'h3e2bb11d, 32'hbe81672d} /* (16, 26, 17) {real, imag} */,
  {32'hbd8b14c0, 32'h3d703d4a} /* (16, 26, 16) {real, imag} */,
  {32'h3e47ac93, 32'hbc9e9f4a} /* (16, 26, 15) {real, imag} */,
  {32'hbda05ba6, 32'h3f101716} /* (16, 26, 14) {real, imag} */,
  {32'h3e78964e, 32'hbd2533bf} /* (16, 26, 13) {real, imag} */,
  {32'hbd35a018, 32'h3f385db2} /* (16, 26, 12) {real, imag} */,
  {32'hbc2f36b0, 32'hbe0860fc} /* (16, 26, 11) {real, imag} */,
  {32'h3e5c52dc, 32'h3d73cbfc} /* (16, 26, 10) {real, imag} */,
  {32'hbe6b0490, 32'hbd319bc0} /* (16, 26, 9) {real, imag} */,
  {32'h3d9fc3c1, 32'h3ee846a6} /* (16, 26, 8) {real, imag} */,
  {32'h3dde029e, 32'hbf0cbda7} /* (16, 26, 7) {real, imag} */,
  {32'hbd9ebc74, 32'h3dd12764} /* (16, 26, 6) {real, imag} */,
  {32'hb9c17c00, 32'hbdeafc42} /* (16, 26, 5) {real, imag} */,
  {32'hbe839244, 32'hbeb650b5} /* (16, 26, 4) {real, imag} */,
  {32'h3cecebe4, 32'h3f46318b} /* (16, 26, 3) {real, imag} */,
  {32'hbf634a9f, 32'hbdd31000} /* (16, 26, 2) {real, imag} */,
  {32'h3eea83e1, 32'hbd8e69cc} /* (16, 26, 1) {real, imag} */,
  {32'hbee4373a, 32'h3f47785a} /* (16, 26, 0) {real, imag} */,
  {32'hbf8e2258, 32'hbec12336} /* (16, 25, 31) {real, imag} */,
  {32'h3e95fb1a, 32'h3ee41866} /* (16, 25, 30) {real, imag} */,
  {32'hbda5b60c, 32'h3de97c23} /* (16, 25, 29) {real, imag} */,
  {32'h3f1a940c, 32'hbe3e27ed} /* (16, 25, 28) {real, imag} */,
  {32'h3e454229, 32'hbe87814e} /* (16, 25, 27) {real, imag} */,
  {32'hbe74ca63, 32'h3e788243} /* (16, 25, 26) {real, imag} */,
  {32'h3db8b28d, 32'h3d4c36d8} /* (16, 25, 25) {real, imag} */,
  {32'hbec81bec, 32'h3d1ca6bc} /* (16, 25, 24) {real, imag} */,
  {32'hbe348c16, 32'h3e9f5a90} /* (16, 25, 23) {real, imag} */,
  {32'h3d664f44, 32'hbec6108e} /* (16, 25, 22) {real, imag} */,
  {32'h3e9cb243, 32'h3eedec23} /* (16, 25, 21) {real, imag} */,
  {32'hbe67da49, 32'h3cebe698} /* (16, 25, 20) {real, imag} */,
  {32'hbe967886, 32'h3ed72bce} /* (16, 25, 19) {real, imag} */,
  {32'h3e8f3f86, 32'hbd5f0ce2} /* (16, 25, 18) {real, imag} */,
  {32'hbef7365a, 32'hbe763554} /* (16, 25, 17) {real, imag} */,
  {32'h3e691d02, 32'h3e283555} /* (16, 25, 16) {real, imag} */,
  {32'hbe6a4d8c, 32'h3d891450} /* (16, 25, 15) {real, imag} */,
  {32'hbe3cd34b, 32'h3e5c146b} /* (16, 25, 14) {real, imag} */,
  {32'h3e0fc175, 32'h3f3d2980} /* (16, 25, 13) {real, imag} */,
  {32'hbf2d22ab, 32'hbe0904e0} /* (16, 25, 12) {real, imag} */,
  {32'h3e8dc0ac, 32'hbe36abdc} /* (16, 25, 11) {real, imag} */,
  {32'h3e4c6de2, 32'h3e747b89} /* (16, 25, 10) {real, imag} */,
  {32'h3ef3b8a2, 32'hbe6d1bb8} /* (16, 25, 9) {real, imag} */,
  {32'hbd81e20f, 32'hbb2cad80} /* (16, 25, 8) {real, imag} */,
  {32'hbe5da323, 32'h3dbba25a} /* (16, 25, 7) {real, imag} */,
  {32'h3e1d4e34, 32'h3e0a75e8} /* (16, 25, 6) {real, imag} */,
  {32'hbdac55ef, 32'h3cc2a76c} /* (16, 25, 5) {real, imag} */,
  {32'hbefebc5e, 32'hbe617932} /* (16, 25, 4) {real, imag} */,
  {32'hbf3d531a, 32'h3c708240} /* (16, 25, 3) {real, imag} */,
  {32'h3ed938be, 32'h3f3f75e4} /* (16, 25, 2) {real, imag} */,
  {32'h3d73a648, 32'hbf83c1b0} /* (16, 25, 1) {real, imag} */,
  {32'hbdab7490, 32'h3eb21a3c} /* (16, 25, 0) {real, imag} */,
  {32'h3f3afc54, 32'hbf719911} /* (16, 24, 31) {real, imag} */,
  {32'hbe62054c, 32'hbd675f36} /* (16, 24, 30) {real, imag} */,
  {32'hbe900690, 32'hbeaa6a21} /* (16, 24, 29) {real, imag} */,
  {32'h3d475044, 32'h3f20916d} /* (16, 24, 28) {real, imag} */,
  {32'h3ebde063, 32'h3efb5a17} /* (16, 24, 27) {real, imag} */,
  {32'h3ee302e4, 32'h3f1518b9} /* (16, 24, 26) {real, imag} */,
  {32'hbe999166, 32'hbf081508} /* (16, 24, 25) {real, imag} */,
  {32'hbd9cbd02, 32'h3ef0eb11} /* (16, 24, 24) {real, imag} */,
  {32'h3eb1c973, 32'hbda1db98} /* (16, 24, 23) {real, imag} */,
  {32'hbec03fbe, 32'hbe4652de} /* (16, 24, 22) {real, imag} */,
  {32'hbedff4e4, 32'hbebcdc1a} /* (16, 24, 21) {real, imag} */,
  {32'h3ec6f27e, 32'hbd893d4e} /* (16, 24, 20) {real, imag} */,
  {32'hbe2bf8c2, 32'hbccaca60} /* (16, 24, 19) {real, imag} */,
  {32'hbe09583c, 32'hbe99f0ed} /* (16, 24, 18) {real, imag} */,
  {32'h3ee36aee, 32'hbe3147ac} /* (16, 24, 17) {real, imag} */,
  {32'hbd75c088, 32'hbe6756d5} /* (16, 24, 16) {real, imag} */,
  {32'h3da51ffb, 32'h3cc16e2a} /* (16, 24, 15) {real, imag} */,
  {32'h3e49b438, 32'hbea4083c} /* (16, 24, 14) {real, imag} */,
  {32'hbf0f07fa, 32'h3eef5374} /* (16, 24, 13) {real, imag} */,
  {32'hbdedd372, 32'hbdfafdcc} /* (16, 24, 12) {real, imag} */,
  {32'h3b831f10, 32'hbe8b4763} /* (16, 24, 11) {real, imag} */,
  {32'hbeb4f0c2, 32'h3f0589df} /* (16, 24, 10) {real, imag} */,
  {32'h3f152c9a, 32'h3e04102d} /* (16, 24, 9) {real, imag} */,
  {32'hbf3b4e97, 32'h3d617ca0} /* (16, 24, 8) {real, imag} */,
  {32'h3b95fc60, 32'h3e96bd29} /* (16, 24, 7) {real, imag} */,
  {32'hbf88a4fb, 32'hbf0385de} /* (16, 24, 6) {real, imag} */,
  {32'hbe97b41f, 32'hbcad34ac} /* (16, 24, 5) {real, imag} */,
  {32'h3e5f0298, 32'h3f01a8fe} /* (16, 24, 4) {real, imag} */,
  {32'hbee85e3a, 32'h3c69b080} /* (16, 24, 3) {real, imag} */,
  {32'hbf3e68b2, 32'h3eefd801} /* (16, 24, 2) {real, imag} */,
  {32'h3e792d32, 32'hbf8e7938} /* (16, 24, 1) {real, imag} */,
  {32'h3ef4daed, 32'hbe96a838} /* (16, 24, 0) {real, imag} */,
  {32'hbe8f69c9, 32'h3e61725c} /* (16, 23, 31) {real, imag} */,
  {32'hbed95fe8, 32'hbf594b4e} /* (16, 23, 30) {real, imag} */,
  {32'h3d9851d6, 32'h3b9e1d80} /* (16, 23, 29) {real, imag} */,
  {32'hbea93bb8, 32'hbeac3dab} /* (16, 23, 28) {real, imag} */,
  {32'h3d49154b, 32'h3c094d40} /* (16, 23, 27) {real, imag} */,
  {32'h3f0ab3b2, 32'h3f389c90} /* (16, 23, 26) {real, imag} */,
  {32'h3f1af1cb, 32'hbe4793c6} /* (16, 23, 25) {real, imag} */,
  {32'hbebe5da1, 32'hbe23af6b} /* (16, 23, 24) {real, imag} */,
  {32'h3eb43dc9, 32'hbec405ae} /* (16, 23, 23) {real, imag} */,
  {32'hbf21ca96, 32'h3e999872} /* (16, 23, 22) {real, imag} */,
  {32'h3e8ed7ec, 32'hbe99cf89} /* (16, 23, 21) {real, imag} */,
  {32'h3e3a1339, 32'hbe34a265} /* (16, 23, 20) {real, imag} */,
  {32'hbe233aa7, 32'hbce2496c} /* (16, 23, 19) {real, imag} */,
  {32'h3e795a54, 32'h3cf59184} /* (16, 23, 18) {real, imag} */,
  {32'h3e601d24, 32'hbe8dc252} /* (16, 23, 17) {real, imag} */,
  {32'hbcaeb338, 32'hbe913a07} /* (16, 23, 16) {real, imag} */,
  {32'h3e92a36e, 32'hbe872ae6} /* (16, 23, 15) {real, imag} */,
  {32'h3e7c7b59, 32'hbeb81228} /* (16, 23, 14) {real, imag} */,
  {32'hbd77874a, 32'h3e20cb22} /* (16, 23, 13) {real, imag} */,
  {32'h3e69cf4b, 32'hbec4b732} /* (16, 23, 12) {real, imag} */,
  {32'hbe8d8e04, 32'h3e973746} /* (16, 23, 11) {real, imag} */,
  {32'hbe88ef1f, 32'hbedb6b3a} /* (16, 23, 10) {real, imag} */,
  {32'hbeb81999, 32'hbeed484c} /* (16, 23, 9) {real, imag} */,
  {32'h3c7e5800, 32'hbdf7aa8b} /* (16, 23, 8) {real, imag} */,
  {32'h3d7b3ede, 32'h3ed6a950} /* (16, 23, 7) {real, imag} */,
  {32'h3f322a8b, 32'hbe87132c} /* (16, 23, 6) {real, imag} */,
  {32'h3e9325f2, 32'h3e23b785} /* (16, 23, 5) {real, imag} */,
  {32'hbe8fdbb2, 32'hbdb330c0} /* (16, 23, 4) {real, imag} */,
  {32'h3e87e81b, 32'h3e84da68} /* (16, 23, 3) {real, imag} */,
  {32'hbebaf3aa, 32'hbe066a1b} /* (16, 23, 2) {real, imag} */,
  {32'hbe6ced88, 32'hbef91898} /* (16, 23, 1) {real, imag} */,
  {32'h3e81cf3d, 32'h3f00fb34} /* (16, 23, 0) {real, imag} */,
  {32'h3c81f0b0, 32'h3e9a3298} /* (16, 22, 31) {real, imag} */,
  {32'h3ea1afc8, 32'h3e02d55a} /* (16, 22, 30) {real, imag} */,
  {32'hbe365c0e, 32'h3e7121a2} /* (16, 22, 29) {real, imag} */,
  {32'h3e9b498c, 32'h3f4a9b39} /* (16, 22, 28) {real, imag} */,
  {32'h3e6f9d00, 32'hbdc67517} /* (16, 22, 27) {real, imag} */,
  {32'h3dc61b26, 32'hbecc05a0} /* (16, 22, 26) {real, imag} */,
  {32'h3dcf9478, 32'h3ddf3462} /* (16, 22, 25) {real, imag} */,
  {32'hbe9d4e97, 32'hbeb23c9e} /* (16, 22, 24) {real, imag} */,
  {32'h3e240f4c, 32'hbdb0f870} /* (16, 22, 23) {real, imag} */,
  {32'h3f125ae8, 32'hbe10f0c3} /* (16, 22, 22) {real, imag} */,
  {32'h3e994178, 32'hbb4b8a30} /* (16, 22, 21) {real, imag} */,
  {32'hbef410a0, 32'hbe3c72d6} /* (16, 22, 20) {real, imag} */,
  {32'h3de387d8, 32'h3eef5fb5} /* (16, 22, 19) {real, imag} */,
  {32'hbf01e9fd, 32'hbed701d3} /* (16, 22, 18) {real, imag} */,
  {32'h3e4e2324, 32'h3e3528d7} /* (16, 22, 17) {real, imag} */,
  {32'hbeb5ff1a, 32'hbea9d092} /* (16, 22, 16) {real, imag} */,
  {32'h3d59e73a, 32'hbf3bc68c} /* (16, 22, 15) {real, imag} */,
  {32'h3d9cbb54, 32'hbdcd690d} /* (16, 22, 14) {real, imag} */,
  {32'h3f35f964, 32'hbea13ff7} /* (16, 22, 13) {real, imag} */,
  {32'h3eec0107, 32'h3f02ad62} /* (16, 22, 12) {real, imag} */,
  {32'hbdbe9554, 32'h3f567618} /* (16, 22, 11) {real, imag} */,
  {32'hbe48a849, 32'hbebe0c27} /* (16, 22, 10) {real, imag} */,
  {32'h3ed0d99f, 32'h3e844364} /* (16, 22, 9) {real, imag} */,
  {32'hbe4e1d87, 32'hbe0491ee} /* (16, 22, 8) {real, imag} */,
  {32'hbefdbe89, 32'hbe1fb19a} /* (16, 22, 7) {real, imag} */,
  {32'hbe8ffbaa, 32'hbf005166} /* (16, 22, 6) {real, imag} */,
  {32'hbf10de90, 32'hbe1d5560} /* (16, 22, 5) {real, imag} */,
  {32'hbf061950, 32'h3d4a81b8} /* (16, 22, 4) {real, imag} */,
  {32'hbe91d38c, 32'hbde8439f} /* (16, 22, 3) {real, imag} */,
  {32'h3f03e306, 32'hbf0dbfdc} /* (16, 22, 2) {real, imag} */,
  {32'h3c992688, 32'h3e93b20e} /* (16, 22, 1) {real, imag} */,
  {32'hbe0ae0e6, 32'h3c243d30} /* (16, 22, 0) {real, imag} */,
  {32'h3e742859, 32'hbe7ae46d} /* (16, 21, 31) {real, imag} */,
  {32'h3e85a62b, 32'h3ea579a7} /* (16, 21, 30) {real, imag} */,
  {32'hbe57c77b, 32'h3e990f94} /* (16, 21, 29) {real, imag} */,
  {32'hbec75cd6, 32'h3df20474} /* (16, 21, 28) {real, imag} */,
  {32'h3ce1d300, 32'h3e93e7ba} /* (16, 21, 27) {real, imag} */,
  {32'hbe03fc47, 32'hbdfc1e84} /* (16, 21, 26) {real, imag} */,
  {32'hbf6e11e8, 32'h3d4c8fc3} /* (16, 21, 25) {real, imag} */,
  {32'h3f08b7f1, 32'hbf2eef45} /* (16, 21, 24) {real, imag} */,
  {32'hbd4309dc, 32'hbed4321c} /* (16, 21, 23) {real, imag} */,
  {32'hbe09cb2e, 32'h3d899941} /* (16, 21, 22) {real, imag} */,
  {32'h3ed0d457, 32'h3e7b1054} /* (16, 21, 21) {real, imag} */,
  {32'hbe8a1ba6, 32'h3e42a748} /* (16, 21, 20) {real, imag} */,
  {32'hbed13d12, 32'hbeed0ef4} /* (16, 21, 19) {real, imag} */,
  {32'hbec9ad96, 32'h3d09afc4} /* (16, 21, 18) {real, imag} */,
  {32'h3ec7d4fa, 32'hb9048200} /* (16, 21, 17) {real, imag} */,
  {32'hbb392540, 32'hbee37ff1} /* (16, 21, 16) {real, imag} */,
  {32'hbe37c2ca, 32'h3e1bbdef} /* (16, 21, 15) {real, imag} */,
  {32'h3eaeeffc, 32'hbd708ddc} /* (16, 21, 14) {real, imag} */,
  {32'hbe4b0ea8, 32'hbce4ab00} /* (16, 21, 13) {real, imag} */,
  {32'hbf0e24ad, 32'hbf482e02} /* (16, 21, 12) {real, imag} */,
  {32'hbd110e58, 32'h3dfa6f0c} /* (16, 21, 11) {real, imag} */,
  {32'h3eba6004, 32'hbdc9f90c} /* (16, 21, 10) {real, imag} */,
  {32'h3f2d8660, 32'h3dfc98f8} /* (16, 21, 9) {real, imag} */,
  {32'hbcba0f00, 32'hbd892e5a} /* (16, 21, 8) {real, imag} */,
  {32'h3d8d3cc7, 32'hbe811628} /* (16, 21, 7) {real, imag} */,
  {32'h3ed31dfa, 32'h3f5812b5} /* (16, 21, 6) {real, imag} */,
  {32'hbe50c494, 32'h3f17f5dc} /* (16, 21, 5) {real, imag} */,
  {32'h3e94ca48, 32'hbeae70a4} /* (16, 21, 4) {real, imag} */,
  {32'h3f11ae65, 32'h3e3218b5} /* (16, 21, 3) {real, imag} */,
  {32'hbd932f28, 32'h3c45c718} /* (16, 21, 2) {real, imag} */,
  {32'hbcadca90, 32'h3deb2840} /* (16, 21, 1) {real, imag} */,
  {32'h3f1acd5a, 32'hbea1ac34} /* (16, 21, 0) {real, imag} */,
  {32'hbd0ca0dc, 32'hbdd30146} /* (16, 20, 31) {real, imag} */,
  {32'hbbad8900, 32'h3d9baf21} /* (16, 20, 30) {real, imag} */,
  {32'hbeaa3deb, 32'hbe94651a} /* (16, 20, 29) {real, imag} */,
  {32'hbdec15a6, 32'h3e149879} /* (16, 20, 28) {real, imag} */,
  {32'hbe57f7b3, 32'h3e1e2778} /* (16, 20, 27) {real, imag} */,
  {32'h3e3ec7d0, 32'h3e930070} /* (16, 20, 26) {real, imag} */,
  {32'h3e3749ad, 32'h3bdddd20} /* (16, 20, 25) {real, imag} */,
  {32'hbd1d72a8, 32'hbf0fad80} /* (16, 20, 24) {real, imag} */,
  {32'h3d85e55c, 32'hbd1eed0c} /* (16, 20, 23) {real, imag} */,
  {32'h3e64edbe, 32'hbec10586} /* (16, 20, 22) {real, imag} */,
  {32'hbe4aa815, 32'hbdc6dcb2} /* (16, 20, 21) {real, imag} */,
  {32'h3da80910, 32'h3f09a76c} /* (16, 20, 20) {real, imag} */,
  {32'hbe3e43cf, 32'h3db9cea8} /* (16, 20, 19) {real, imag} */,
  {32'hbe8a1115, 32'h3ea5a04c} /* (16, 20, 18) {real, imag} */,
  {32'hbd535114, 32'hbdd2ff1c} /* (16, 20, 17) {real, imag} */,
  {32'h3c4de2d4, 32'hbd33ede2} /* (16, 20, 16) {real, imag} */,
  {32'hbe6543b2, 32'h3f1aa1a3} /* (16, 20, 15) {real, imag} */,
  {32'hbe15ef9b, 32'hbf123193} /* (16, 20, 14) {real, imag} */,
  {32'h3f0b5523, 32'hbd830112} /* (16, 20, 13) {real, imag} */,
  {32'hbe443a97, 32'h3e04b8fa} /* (16, 20, 12) {real, imag} */,
  {32'hbf0064a2, 32'h3e83663b} /* (16, 20, 11) {real, imag} */,
  {32'hbd77669f, 32'hbf0f40c2} /* (16, 20, 10) {real, imag} */,
  {32'hbea9cab9, 32'hbe4de0b5} /* (16, 20, 9) {real, imag} */,
  {32'h3e4091df, 32'h3e27a6a6} /* (16, 20, 8) {real, imag} */,
  {32'h3d655f20, 32'hbc320b78} /* (16, 20, 7) {real, imag} */,
  {32'h3df5486d, 32'h3ee90f70} /* (16, 20, 6) {real, imag} */,
  {32'hbe8237f4, 32'h3e0fa772} /* (16, 20, 5) {real, imag} */,
  {32'h39462200, 32'h3c640a20} /* (16, 20, 4) {real, imag} */,
  {32'hbdcd876b, 32'h3e872dcc} /* (16, 20, 3) {real, imag} */,
  {32'h3efa5444, 32'hbe1e1ca2} /* (16, 20, 2) {real, imag} */,
  {32'hbea7b835, 32'hbbdbeec0} /* (16, 20, 1) {real, imag} */,
  {32'h3db53da6, 32'h3e0e11fc} /* (16, 20, 0) {real, imag} */,
  {32'hbe9735f4, 32'h3eb67d3e} /* (16, 19, 31) {real, imag} */,
  {32'hbe353adb, 32'h3d2ebf2e} /* (16, 19, 30) {real, imag} */,
  {32'hbde03aec, 32'hbefda553} /* (16, 19, 29) {real, imag} */,
  {32'hbd651d88, 32'h3eb46ff9} /* (16, 19, 28) {real, imag} */,
  {32'h3d2107b1, 32'h3e3fe432} /* (16, 19, 27) {real, imag} */,
  {32'h3d711356, 32'hbf5b34e6} /* (16, 19, 26) {real, imag} */,
  {32'hbec14d4a, 32'h3e8f7559} /* (16, 19, 25) {real, imag} */,
  {32'h3f1d685c, 32'hbd673930} /* (16, 19, 24) {real, imag} */,
  {32'hbb1de940, 32'hbeb24954} /* (16, 19, 23) {real, imag} */,
  {32'h3f095a34, 32'hbeccc114} /* (16, 19, 22) {real, imag} */,
  {32'hbe33a8a6, 32'hbe6c4cc1} /* (16, 19, 21) {real, imag} */,
  {32'h3e65dda4, 32'h3ece5280} /* (16, 19, 20) {real, imag} */,
  {32'hbde2405c, 32'h3d0cb371} /* (16, 19, 19) {real, imag} */,
  {32'h3e2dba14, 32'hbdae1069} /* (16, 19, 18) {real, imag} */,
  {32'h3ea014d6, 32'h3e1e61aa} /* (16, 19, 17) {real, imag} */,
  {32'hbe8de0fd, 32'h3e82b515} /* (16, 19, 16) {real, imag} */,
  {32'h3d982cd0, 32'hbdfe1861} /* (16, 19, 15) {real, imag} */,
  {32'h3dc5b92c, 32'hbd393ff4} /* (16, 19, 14) {real, imag} */,
  {32'h3e92908a, 32'hbde599de} /* (16, 19, 13) {real, imag} */,
  {32'hbd81eda8, 32'hbdeca543} /* (16, 19, 12) {real, imag} */,
  {32'h3daedf42, 32'h3d9d035f} /* (16, 19, 11) {real, imag} */,
  {32'hbbd9cc30, 32'h3e1a80e6} /* (16, 19, 10) {real, imag} */,
  {32'hbdfd5580, 32'hbda00c42} /* (16, 19, 9) {real, imag} */,
  {32'hbf02e43f, 32'h3e70c816} /* (16, 19, 8) {real, imag} */,
  {32'h3cfdd340, 32'hbf04f1ee} /* (16, 19, 7) {real, imag} */,
  {32'hbf01fd21, 32'hbe9db568} /* (16, 19, 6) {real, imag} */,
  {32'h3edbb36b, 32'hbd3e834c} /* (16, 19, 5) {real, imag} */,
  {32'hb9eee680, 32'hbdf87ed6} /* (16, 19, 4) {real, imag} */,
  {32'h3e025cf3, 32'hbea73b38} /* (16, 19, 3) {real, imag} */,
  {32'h3e08a2e3, 32'h3e3dccd6} /* (16, 19, 2) {real, imag} */,
  {32'hbbcd4aa0, 32'h3dc89c7c} /* (16, 19, 1) {real, imag} */,
  {32'h3e94ef5e, 32'h3e535019} /* (16, 19, 0) {real, imag} */,
  {32'h3e4e0811, 32'hbd9d3cce} /* (16, 18, 31) {real, imag} */,
  {32'hbe0258b4, 32'h3e8b9474} /* (16, 18, 30) {real, imag} */,
  {32'h3e3b583d, 32'h3ea64ab4} /* (16, 18, 29) {real, imag} */,
  {32'h3e27a766, 32'hbe5ea23b} /* (16, 18, 28) {real, imag} */,
  {32'h3c98bf38, 32'h3e126c6e} /* (16, 18, 27) {real, imag} */,
  {32'hbeb00030, 32'h3e0ca6fa} /* (16, 18, 26) {real, imag} */,
  {32'hbd0c1a3c, 32'h3f09a076} /* (16, 18, 25) {real, imag} */,
  {32'hbe9262e9, 32'hbda0357c} /* (16, 18, 24) {real, imag} */,
  {32'h3c63f160, 32'h3e37537a} /* (16, 18, 23) {real, imag} */,
  {32'hbd432a34, 32'h3f1cadaa} /* (16, 18, 22) {real, imag} */,
  {32'h3deb5a4a, 32'h3c9b6af0} /* (16, 18, 21) {real, imag} */,
  {32'hbd95d314, 32'hbf077534} /* (16, 18, 20) {real, imag} */,
  {32'h3e2b97e1, 32'h3e8e0940} /* (16, 18, 19) {real, imag} */,
  {32'h3bf22fe8, 32'hbea7de98} /* (16, 18, 18) {real, imag} */,
  {32'h3e8966b6, 32'h3d2aa1aa} /* (16, 18, 17) {real, imag} */,
  {32'hbeb4376f, 32'h3d59a214} /* (16, 18, 16) {real, imag} */,
  {32'hbe912859, 32'hbedfe9f0} /* (16, 18, 15) {real, imag} */,
  {32'hbe915e02, 32'h3bce7360} /* (16, 18, 14) {real, imag} */,
  {32'hbda9e36c, 32'h3e04f060} /* (16, 18, 13) {real, imag} */,
  {32'hbd97e7e0, 32'hbe34aeed} /* (16, 18, 12) {real, imag} */,
  {32'h3e860fbe, 32'hbdc98b72} /* (16, 18, 11) {real, imag} */,
  {32'hbea966ee, 32'h3e6463ce} /* (16, 18, 10) {real, imag} */,
  {32'h3d7be2ea, 32'h3f115462} /* (16, 18, 9) {real, imag} */,
  {32'h3e98d928, 32'h3e8de5a4} /* (16, 18, 8) {real, imag} */,
  {32'h3e4580cf, 32'hbeac0560} /* (16, 18, 7) {real, imag} */,
  {32'h3eac316c, 32'h3e0a96f7} /* (16, 18, 6) {real, imag} */,
  {32'h3e0d79e8, 32'hbeb07d21} /* (16, 18, 5) {real, imag} */,
  {32'h3ee98586, 32'h3e8ef6af} /* (16, 18, 4) {real, imag} */,
  {32'h3dbfdb2b, 32'hbd531278} /* (16, 18, 3) {real, imag} */,
  {32'h3e168743, 32'h3db2cf72} /* (16, 18, 2) {real, imag} */,
  {32'h3e32b50b, 32'hbeb4ad20} /* (16, 18, 1) {real, imag} */,
  {32'hbe6b84a3, 32'hbf0a40de} /* (16, 18, 0) {real, imag} */,
  {32'hbdc62245, 32'h3e8e5ac6} /* (16, 17, 31) {real, imag} */,
  {32'h3e0c0c53, 32'h3c89c638} /* (16, 17, 30) {real, imag} */,
  {32'h3d7fac28, 32'hbeb882e0} /* (16, 17, 29) {real, imag} */,
  {32'hbca63296, 32'hbe2ce88e} /* (16, 17, 28) {real, imag} */,
  {32'hbe32ce8a, 32'hbcebbd3a} /* (16, 17, 27) {real, imag} */,
  {32'h3c505840, 32'h3ea960f6} /* (16, 17, 26) {real, imag} */,
  {32'h3d4a4774, 32'hbe0dc8b8} /* (16, 17, 25) {real, imag} */,
  {32'hbdfcc876, 32'h3e4c1fb2} /* (16, 17, 24) {real, imag} */,
  {32'h3eaf9704, 32'h3eb012d3} /* (16, 17, 23) {real, imag} */,
  {32'hbe4944b3, 32'hbe0e94a8} /* (16, 17, 22) {real, imag} */,
  {32'h3e399cd5, 32'h3f2f28b6} /* (16, 17, 21) {real, imag} */,
  {32'hbdc43202, 32'h3ee906b5} /* (16, 17, 20) {real, imag} */,
  {32'h3bdcc100, 32'hbdba909b} /* (16, 17, 19) {real, imag} */,
  {32'hbe90e5da, 32'h3eae1f53} /* (16, 17, 18) {real, imag} */,
  {32'hbd888ea8, 32'h3e738a42} /* (16, 17, 17) {real, imag} */,
  {32'h3d3078d0, 32'hbb392270} /* (16, 17, 16) {real, imag} */,
  {32'hbca2c0b8, 32'hbe9075a8} /* (16, 17, 15) {real, imag} */,
  {32'h3eb94087, 32'hbe27001b} /* (16, 17, 14) {real, imag} */,
  {32'hbe26816c, 32'hbec575b7} /* (16, 17, 13) {real, imag} */,
  {32'hbdf8e5f0, 32'hbe08d284} /* (16, 17, 12) {real, imag} */,
  {32'hbefbdc8f, 32'h3e40e90e} /* (16, 17, 11) {real, imag} */,
  {32'h3eb3e1bb, 32'h3e8b7ff0} /* (16, 17, 10) {real, imag} */,
  {32'h3e647389, 32'h3d88c577} /* (16, 17, 9) {real, imag} */,
  {32'h3e663b2c, 32'hbd82450b} /* (16, 17, 8) {real, imag} */,
  {32'h3e80fd1a, 32'h3e927b78} /* (16, 17, 7) {real, imag} */,
  {32'h3e51320d, 32'hbeafc0bc} /* (16, 17, 6) {real, imag} */,
  {32'hbe1ccfb2, 32'h3ea44556} /* (16, 17, 5) {real, imag} */,
  {32'hbcac2cdc, 32'h3df7b260} /* (16, 17, 4) {real, imag} */,
  {32'h3e73a6d0, 32'h3e3f046a} /* (16, 17, 3) {real, imag} */,
  {32'hbe73aedc, 32'h3cbcb940} /* (16, 17, 2) {real, imag} */,
  {32'h3e1e6998, 32'hbdeee26a} /* (16, 17, 1) {real, imag} */,
  {32'h3d816c62, 32'hbde18c12} /* (16, 17, 0) {real, imag} */,
  {32'h3c0f7344, 32'hbdfd1b94} /* (16, 16, 31) {real, imag} */,
  {32'hbc908d80, 32'hbe58f684} /* (16, 16, 30) {real, imag} */,
  {32'hbe4e884f, 32'h3df95643} /* (16, 16, 29) {real, imag} */,
  {32'hbd1853d7, 32'hbea03216} /* (16, 16, 28) {real, imag} */,
  {32'hbe67b5a0, 32'hbe48bc34} /* (16, 16, 27) {real, imag} */,
  {32'hbe217485, 32'h3e2f8b28} /* (16, 16, 26) {real, imag} */,
  {32'h3e8202a0, 32'h3e85954a} /* (16, 16, 25) {real, imag} */,
  {32'hbeb80873, 32'hbe2575bb} /* (16, 16, 24) {real, imag} */,
  {32'hbe20b7f8, 32'hbc18c8c8} /* (16, 16, 23) {real, imag} */,
  {32'hbe278fec, 32'h3e408f7a} /* (16, 16, 22) {real, imag} */,
  {32'h3d75c469, 32'hbe2329dc} /* (16, 16, 21) {real, imag} */,
  {32'h3ecabf08, 32'hbea5bf3a} /* (16, 16, 20) {real, imag} */,
  {32'hbb8c6f88, 32'h3e924a00} /* (16, 16, 19) {real, imag} */,
  {32'h3e023e92, 32'hbe6392b6} /* (16, 16, 18) {real, imag} */,
  {32'h3d9bc844, 32'h39de4e00} /* (16, 16, 17) {real, imag} */,
  {32'h3dc8067c, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h3d9bc844, 32'hb9de4e00} /* (16, 16, 15) {real, imag} */,
  {32'h3e023e92, 32'h3e6392b6} /* (16, 16, 14) {real, imag} */,
  {32'hbb8c6f88, 32'hbe924a00} /* (16, 16, 13) {real, imag} */,
  {32'h3ecabf08, 32'h3ea5bf3a} /* (16, 16, 12) {real, imag} */,
  {32'h3d75c469, 32'h3e2329dc} /* (16, 16, 11) {real, imag} */,
  {32'hbe278fec, 32'hbe408f7a} /* (16, 16, 10) {real, imag} */,
  {32'hbe20b7f8, 32'h3c18c8c8} /* (16, 16, 9) {real, imag} */,
  {32'hbeb80873, 32'h3e2575bb} /* (16, 16, 8) {real, imag} */,
  {32'h3e8202a0, 32'hbe85954a} /* (16, 16, 7) {real, imag} */,
  {32'hbe217485, 32'hbe2f8b28} /* (16, 16, 6) {real, imag} */,
  {32'hbe67b5a0, 32'h3e48bc34} /* (16, 16, 5) {real, imag} */,
  {32'hbd1853d7, 32'h3ea03216} /* (16, 16, 4) {real, imag} */,
  {32'hbe4e884f, 32'hbdf95643} /* (16, 16, 3) {real, imag} */,
  {32'hbc908d80, 32'h3e58f684} /* (16, 16, 2) {real, imag} */,
  {32'h3c0f7344, 32'h3dfd1b94} /* (16, 16, 1) {real, imag} */,
  {32'hbe1eef1f, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h3e1e6998, 32'h3deee26a} /* (16, 15, 31) {real, imag} */,
  {32'hbe73aedc, 32'hbcbcb940} /* (16, 15, 30) {real, imag} */,
  {32'h3e73a6d0, 32'hbe3f046a} /* (16, 15, 29) {real, imag} */,
  {32'hbcac2cdc, 32'hbdf7b260} /* (16, 15, 28) {real, imag} */,
  {32'hbe1ccfb2, 32'hbea44556} /* (16, 15, 27) {real, imag} */,
  {32'h3e51320d, 32'h3eafc0bc} /* (16, 15, 26) {real, imag} */,
  {32'h3e80fd1a, 32'hbe927b78} /* (16, 15, 25) {real, imag} */,
  {32'h3e663b2c, 32'h3d82450b} /* (16, 15, 24) {real, imag} */,
  {32'h3e647389, 32'hbd88c577} /* (16, 15, 23) {real, imag} */,
  {32'h3eb3e1bb, 32'hbe8b7ff0} /* (16, 15, 22) {real, imag} */,
  {32'hbefbdc8f, 32'hbe40e90e} /* (16, 15, 21) {real, imag} */,
  {32'hbdf8e5f0, 32'h3e08d284} /* (16, 15, 20) {real, imag} */,
  {32'hbe26816c, 32'h3ec575b7} /* (16, 15, 19) {real, imag} */,
  {32'h3eb94087, 32'h3e27001b} /* (16, 15, 18) {real, imag} */,
  {32'hbca2c0b8, 32'h3e9075a8} /* (16, 15, 17) {real, imag} */,
  {32'h3d3078d0, 32'h3b392270} /* (16, 15, 16) {real, imag} */,
  {32'hbd888ea8, 32'hbe738a42} /* (16, 15, 15) {real, imag} */,
  {32'hbe90e5da, 32'hbeae1f53} /* (16, 15, 14) {real, imag} */,
  {32'h3bdcc100, 32'h3dba909b} /* (16, 15, 13) {real, imag} */,
  {32'hbdc43202, 32'hbee906b5} /* (16, 15, 12) {real, imag} */,
  {32'h3e399cd5, 32'hbf2f28b6} /* (16, 15, 11) {real, imag} */,
  {32'hbe4944b3, 32'h3e0e94a8} /* (16, 15, 10) {real, imag} */,
  {32'h3eaf9704, 32'hbeb012d3} /* (16, 15, 9) {real, imag} */,
  {32'hbdfcc876, 32'hbe4c1fb2} /* (16, 15, 8) {real, imag} */,
  {32'h3d4a4774, 32'h3e0dc8b8} /* (16, 15, 7) {real, imag} */,
  {32'h3c505840, 32'hbea960f6} /* (16, 15, 6) {real, imag} */,
  {32'hbe32ce8a, 32'h3cebbd3a} /* (16, 15, 5) {real, imag} */,
  {32'hbca63296, 32'h3e2ce88e} /* (16, 15, 4) {real, imag} */,
  {32'h3d7fac28, 32'h3eb882e0} /* (16, 15, 3) {real, imag} */,
  {32'h3e0c0c53, 32'hbc89c638} /* (16, 15, 2) {real, imag} */,
  {32'hbdc62245, 32'hbe8e5ac6} /* (16, 15, 1) {real, imag} */,
  {32'h3d816c62, 32'h3de18c12} /* (16, 15, 0) {real, imag} */,
  {32'h3e32b50b, 32'h3eb4ad20} /* (16, 14, 31) {real, imag} */,
  {32'h3e168743, 32'hbdb2cf72} /* (16, 14, 30) {real, imag} */,
  {32'h3dbfdb2b, 32'h3d531278} /* (16, 14, 29) {real, imag} */,
  {32'h3ee98586, 32'hbe8ef6af} /* (16, 14, 28) {real, imag} */,
  {32'h3e0d79e8, 32'h3eb07d21} /* (16, 14, 27) {real, imag} */,
  {32'h3eac316c, 32'hbe0a96f7} /* (16, 14, 26) {real, imag} */,
  {32'h3e4580cf, 32'h3eac0560} /* (16, 14, 25) {real, imag} */,
  {32'h3e98d928, 32'hbe8de5a4} /* (16, 14, 24) {real, imag} */,
  {32'h3d7be2ea, 32'hbf115462} /* (16, 14, 23) {real, imag} */,
  {32'hbea966ee, 32'hbe6463ce} /* (16, 14, 22) {real, imag} */,
  {32'h3e860fbe, 32'h3dc98b72} /* (16, 14, 21) {real, imag} */,
  {32'hbd97e7e0, 32'h3e34aeed} /* (16, 14, 20) {real, imag} */,
  {32'hbda9e36c, 32'hbe04f060} /* (16, 14, 19) {real, imag} */,
  {32'hbe915e02, 32'hbbce7360} /* (16, 14, 18) {real, imag} */,
  {32'hbe912859, 32'h3edfe9f0} /* (16, 14, 17) {real, imag} */,
  {32'hbeb4376f, 32'hbd59a214} /* (16, 14, 16) {real, imag} */,
  {32'h3e8966b6, 32'hbd2aa1aa} /* (16, 14, 15) {real, imag} */,
  {32'h3bf22fe8, 32'h3ea7de98} /* (16, 14, 14) {real, imag} */,
  {32'h3e2b97e1, 32'hbe8e0940} /* (16, 14, 13) {real, imag} */,
  {32'hbd95d314, 32'h3f077534} /* (16, 14, 12) {real, imag} */,
  {32'h3deb5a4a, 32'hbc9b6af0} /* (16, 14, 11) {real, imag} */,
  {32'hbd432a34, 32'hbf1cadaa} /* (16, 14, 10) {real, imag} */,
  {32'h3c63f160, 32'hbe37537a} /* (16, 14, 9) {real, imag} */,
  {32'hbe9262e9, 32'h3da0357c} /* (16, 14, 8) {real, imag} */,
  {32'hbd0c1a3c, 32'hbf09a076} /* (16, 14, 7) {real, imag} */,
  {32'hbeb00030, 32'hbe0ca6fa} /* (16, 14, 6) {real, imag} */,
  {32'h3c98bf38, 32'hbe126c6e} /* (16, 14, 5) {real, imag} */,
  {32'h3e27a766, 32'h3e5ea23b} /* (16, 14, 4) {real, imag} */,
  {32'h3e3b583d, 32'hbea64ab4} /* (16, 14, 3) {real, imag} */,
  {32'hbe0258b4, 32'hbe8b9474} /* (16, 14, 2) {real, imag} */,
  {32'h3e4e0811, 32'h3d9d3cce} /* (16, 14, 1) {real, imag} */,
  {32'hbe6b84a3, 32'h3f0a40de} /* (16, 14, 0) {real, imag} */,
  {32'hbbcd4aa0, 32'hbdc89c7c} /* (16, 13, 31) {real, imag} */,
  {32'h3e08a2e3, 32'hbe3dccd6} /* (16, 13, 30) {real, imag} */,
  {32'h3e025cf3, 32'h3ea73b38} /* (16, 13, 29) {real, imag} */,
  {32'hb9eee680, 32'h3df87ed6} /* (16, 13, 28) {real, imag} */,
  {32'h3edbb36b, 32'h3d3e834c} /* (16, 13, 27) {real, imag} */,
  {32'hbf01fd21, 32'h3e9db568} /* (16, 13, 26) {real, imag} */,
  {32'h3cfdd340, 32'h3f04f1ee} /* (16, 13, 25) {real, imag} */,
  {32'hbf02e43f, 32'hbe70c816} /* (16, 13, 24) {real, imag} */,
  {32'hbdfd5580, 32'h3da00c42} /* (16, 13, 23) {real, imag} */,
  {32'hbbd9cc30, 32'hbe1a80e6} /* (16, 13, 22) {real, imag} */,
  {32'h3daedf42, 32'hbd9d035f} /* (16, 13, 21) {real, imag} */,
  {32'hbd81eda8, 32'h3deca543} /* (16, 13, 20) {real, imag} */,
  {32'h3e92908a, 32'h3de599de} /* (16, 13, 19) {real, imag} */,
  {32'h3dc5b92c, 32'h3d393ff4} /* (16, 13, 18) {real, imag} */,
  {32'h3d982cd0, 32'h3dfe1861} /* (16, 13, 17) {real, imag} */,
  {32'hbe8de0fd, 32'hbe82b515} /* (16, 13, 16) {real, imag} */,
  {32'h3ea014d6, 32'hbe1e61aa} /* (16, 13, 15) {real, imag} */,
  {32'h3e2dba14, 32'h3dae1069} /* (16, 13, 14) {real, imag} */,
  {32'hbde2405c, 32'hbd0cb371} /* (16, 13, 13) {real, imag} */,
  {32'h3e65dda4, 32'hbece5280} /* (16, 13, 12) {real, imag} */,
  {32'hbe33a8a6, 32'h3e6c4cc1} /* (16, 13, 11) {real, imag} */,
  {32'h3f095a34, 32'h3eccc114} /* (16, 13, 10) {real, imag} */,
  {32'hbb1de940, 32'h3eb24954} /* (16, 13, 9) {real, imag} */,
  {32'h3f1d685c, 32'h3d673930} /* (16, 13, 8) {real, imag} */,
  {32'hbec14d4a, 32'hbe8f7559} /* (16, 13, 7) {real, imag} */,
  {32'h3d711356, 32'h3f5b34e6} /* (16, 13, 6) {real, imag} */,
  {32'h3d2107b1, 32'hbe3fe432} /* (16, 13, 5) {real, imag} */,
  {32'hbd651d88, 32'hbeb46ff9} /* (16, 13, 4) {real, imag} */,
  {32'hbde03aec, 32'h3efda553} /* (16, 13, 3) {real, imag} */,
  {32'hbe353adb, 32'hbd2ebf2e} /* (16, 13, 2) {real, imag} */,
  {32'hbe9735f4, 32'hbeb67d3e} /* (16, 13, 1) {real, imag} */,
  {32'h3e94ef5e, 32'hbe535019} /* (16, 13, 0) {real, imag} */,
  {32'hbea7b835, 32'h3bdbeec0} /* (16, 12, 31) {real, imag} */,
  {32'h3efa5444, 32'h3e1e1ca2} /* (16, 12, 30) {real, imag} */,
  {32'hbdcd876b, 32'hbe872dcc} /* (16, 12, 29) {real, imag} */,
  {32'h39462200, 32'hbc640a20} /* (16, 12, 28) {real, imag} */,
  {32'hbe8237f4, 32'hbe0fa772} /* (16, 12, 27) {real, imag} */,
  {32'h3df5486d, 32'hbee90f70} /* (16, 12, 26) {real, imag} */,
  {32'h3d655f20, 32'h3c320b78} /* (16, 12, 25) {real, imag} */,
  {32'h3e4091df, 32'hbe27a6a6} /* (16, 12, 24) {real, imag} */,
  {32'hbea9cab9, 32'h3e4de0b5} /* (16, 12, 23) {real, imag} */,
  {32'hbd77669f, 32'h3f0f40c2} /* (16, 12, 22) {real, imag} */,
  {32'hbf0064a2, 32'hbe83663b} /* (16, 12, 21) {real, imag} */,
  {32'hbe443a97, 32'hbe04b8fa} /* (16, 12, 20) {real, imag} */,
  {32'h3f0b5523, 32'h3d830112} /* (16, 12, 19) {real, imag} */,
  {32'hbe15ef9b, 32'h3f123193} /* (16, 12, 18) {real, imag} */,
  {32'hbe6543b2, 32'hbf1aa1a3} /* (16, 12, 17) {real, imag} */,
  {32'h3c4de2d4, 32'h3d33ede2} /* (16, 12, 16) {real, imag} */,
  {32'hbd535114, 32'h3dd2ff1c} /* (16, 12, 15) {real, imag} */,
  {32'hbe8a1115, 32'hbea5a04c} /* (16, 12, 14) {real, imag} */,
  {32'hbe3e43cf, 32'hbdb9cea8} /* (16, 12, 13) {real, imag} */,
  {32'h3da80910, 32'hbf09a76c} /* (16, 12, 12) {real, imag} */,
  {32'hbe4aa815, 32'h3dc6dcb2} /* (16, 12, 11) {real, imag} */,
  {32'h3e64edbe, 32'h3ec10586} /* (16, 12, 10) {real, imag} */,
  {32'h3d85e55c, 32'h3d1eed0c} /* (16, 12, 9) {real, imag} */,
  {32'hbd1d72a8, 32'h3f0fad80} /* (16, 12, 8) {real, imag} */,
  {32'h3e3749ad, 32'hbbdddd20} /* (16, 12, 7) {real, imag} */,
  {32'h3e3ec7d0, 32'hbe930070} /* (16, 12, 6) {real, imag} */,
  {32'hbe57f7b3, 32'hbe1e2778} /* (16, 12, 5) {real, imag} */,
  {32'hbdec15a6, 32'hbe149879} /* (16, 12, 4) {real, imag} */,
  {32'hbeaa3deb, 32'h3e94651a} /* (16, 12, 3) {real, imag} */,
  {32'hbbad8900, 32'hbd9baf21} /* (16, 12, 2) {real, imag} */,
  {32'hbd0ca0dc, 32'h3dd30146} /* (16, 12, 1) {real, imag} */,
  {32'h3db53da6, 32'hbe0e11fc} /* (16, 12, 0) {real, imag} */,
  {32'hbcadca90, 32'hbdeb2840} /* (16, 11, 31) {real, imag} */,
  {32'hbd932f28, 32'hbc45c718} /* (16, 11, 30) {real, imag} */,
  {32'h3f11ae65, 32'hbe3218b5} /* (16, 11, 29) {real, imag} */,
  {32'h3e94ca48, 32'h3eae70a4} /* (16, 11, 28) {real, imag} */,
  {32'hbe50c494, 32'hbf17f5dc} /* (16, 11, 27) {real, imag} */,
  {32'h3ed31dfa, 32'hbf5812b5} /* (16, 11, 26) {real, imag} */,
  {32'h3d8d3cc7, 32'h3e811628} /* (16, 11, 25) {real, imag} */,
  {32'hbcba0f00, 32'h3d892e5a} /* (16, 11, 24) {real, imag} */,
  {32'h3f2d8660, 32'hbdfc98f8} /* (16, 11, 23) {real, imag} */,
  {32'h3eba6004, 32'h3dc9f90c} /* (16, 11, 22) {real, imag} */,
  {32'hbd110e58, 32'hbdfa6f0c} /* (16, 11, 21) {real, imag} */,
  {32'hbf0e24ad, 32'h3f482e02} /* (16, 11, 20) {real, imag} */,
  {32'hbe4b0ea8, 32'h3ce4ab00} /* (16, 11, 19) {real, imag} */,
  {32'h3eaeeffc, 32'h3d708ddc} /* (16, 11, 18) {real, imag} */,
  {32'hbe37c2ca, 32'hbe1bbdef} /* (16, 11, 17) {real, imag} */,
  {32'hbb392540, 32'h3ee37ff1} /* (16, 11, 16) {real, imag} */,
  {32'h3ec7d4fa, 32'h39048200} /* (16, 11, 15) {real, imag} */,
  {32'hbec9ad96, 32'hbd09afc4} /* (16, 11, 14) {real, imag} */,
  {32'hbed13d12, 32'h3eed0ef4} /* (16, 11, 13) {real, imag} */,
  {32'hbe8a1ba6, 32'hbe42a748} /* (16, 11, 12) {real, imag} */,
  {32'h3ed0d457, 32'hbe7b1054} /* (16, 11, 11) {real, imag} */,
  {32'hbe09cb2e, 32'hbd899941} /* (16, 11, 10) {real, imag} */,
  {32'hbd4309dc, 32'h3ed4321c} /* (16, 11, 9) {real, imag} */,
  {32'h3f08b7f1, 32'h3f2eef45} /* (16, 11, 8) {real, imag} */,
  {32'hbf6e11e8, 32'hbd4c8fc3} /* (16, 11, 7) {real, imag} */,
  {32'hbe03fc47, 32'h3dfc1e84} /* (16, 11, 6) {real, imag} */,
  {32'h3ce1d300, 32'hbe93e7ba} /* (16, 11, 5) {real, imag} */,
  {32'hbec75cd6, 32'hbdf20474} /* (16, 11, 4) {real, imag} */,
  {32'hbe57c77b, 32'hbe990f94} /* (16, 11, 3) {real, imag} */,
  {32'h3e85a62b, 32'hbea579a7} /* (16, 11, 2) {real, imag} */,
  {32'h3e742859, 32'h3e7ae46d} /* (16, 11, 1) {real, imag} */,
  {32'h3f1acd5a, 32'h3ea1ac34} /* (16, 11, 0) {real, imag} */,
  {32'h3c992688, 32'hbe93b20e} /* (16, 10, 31) {real, imag} */,
  {32'h3f03e306, 32'h3f0dbfdc} /* (16, 10, 30) {real, imag} */,
  {32'hbe91d38c, 32'h3de8439f} /* (16, 10, 29) {real, imag} */,
  {32'hbf061950, 32'hbd4a81b8} /* (16, 10, 28) {real, imag} */,
  {32'hbf10de90, 32'h3e1d5560} /* (16, 10, 27) {real, imag} */,
  {32'hbe8ffbaa, 32'h3f005166} /* (16, 10, 26) {real, imag} */,
  {32'hbefdbe89, 32'h3e1fb19a} /* (16, 10, 25) {real, imag} */,
  {32'hbe4e1d87, 32'h3e0491ee} /* (16, 10, 24) {real, imag} */,
  {32'h3ed0d99f, 32'hbe844364} /* (16, 10, 23) {real, imag} */,
  {32'hbe48a849, 32'h3ebe0c27} /* (16, 10, 22) {real, imag} */,
  {32'hbdbe9554, 32'hbf567618} /* (16, 10, 21) {real, imag} */,
  {32'h3eec0107, 32'hbf02ad62} /* (16, 10, 20) {real, imag} */,
  {32'h3f35f964, 32'h3ea13ff7} /* (16, 10, 19) {real, imag} */,
  {32'h3d9cbb54, 32'h3dcd690d} /* (16, 10, 18) {real, imag} */,
  {32'h3d59e73a, 32'h3f3bc68c} /* (16, 10, 17) {real, imag} */,
  {32'hbeb5ff1a, 32'h3ea9d092} /* (16, 10, 16) {real, imag} */,
  {32'h3e4e2324, 32'hbe3528d7} /* (16, 10, 15) {real, imag} */,
  {32'hbf01e9fd, 32'h3ed701d3} /* (16, 10, 14) {real, imag} */,
  {32'h3de387d8, 32'hbeef5fb5} /* (16, 10, 13) {real, imag} */,
  {32'hbef410a0, 32'h3e3c72d6} /* (16, 10, 12) {real, imag} */,
  {32'h3e994178, 32'h3b4b8a30} /* (16, 10, 11) {real, imag} */,
  {32'h3f125ae8, 32'h3e10f0c3} /* (16, 10, 10) {real, imag} */,
  {32'h3e240f4c, 32'h3db0f870} /* (16, 10, 9) {real, imag} */,
  {32'hbe9d4e97, 32'h3eb23c9e} /* (16, 10, 8) {real, imag} */,
  {32'h3dcf9478, 32'hbddf3462} /* (16, 10, 7) {real, imag} */,
  {32'h3dc61b26, 32'h3ecc05a0} /* (16, 10, 6) {real, imag} */,
  {32'h3e6f9d00, 32'h3dc67517} /* (16, 10, 5) {real, imag} */,
  {32'h3e9b498c, 32'hbf4a9b39} /* (16, 10, 4) {real, imag} */,
  {32'hbe365c0e, 32'hbe7121a2} /* (16, 10, 3) {real, imag} */,
  {32'h3ea1afc8, 32'hbe02d55a} /* (16, 10, 2) {real, imag} */,
  {32'h3c81f0b0, 32'hbe9a3298} /* (16, 10, 1) {real, imag} */,
  {32'hbe0ae0e6, 32'hbc243d30} /* (16, 10, 0) {real, imag} */,
  {32'hbe6ced88, 32'h3ef91898} /* (16, 9, 31) {real, imag} */,
  {32'hbebaf3aa, 32'h3e066a1b} /* (16, 9, 30) {real, imag} */,
  {32'h3e87e81b, 32'hbe84da68} /* (16, 9, 29) {real, imag} */,
  {32'hbe8fdbb2, 32'h3db330c0} /* (16, 9, 28) {real, imag} */,
  {32'h3e9325f2, 32'hbe23b785} /* (16, 9, 27) {real, imag} */,
  {32'h3f322a8b, 32'h3e87132c} /* (16, 9, 26) {real, imag} */,
  {32'h3d7b3ede, 32'hbed6a950} /* (16, 9, 25) {real, imag} */,
  {32'h3c7e5800, 32'h3df7aa8b} /* (16, 9, 24) {real, imag} */,
  {32'hbeb81999, 32'h3eed484c} /* (16, 9, 23) {real, imag} */,
  {32'hbe88ef1f, 32'h3edb6b3a} /* (16, 9, 22) {real, imag} */,
  {32'hbe8d8e04, 32'hbe973746} /* (16, 9, 21) {real, imag} */,
  {32'h3e69cf4b, 32'h3ec4b732} /* (16, 9, 20) {real, imag} */,
  {32'hbd77874a, 32'hbe20cb22} /* (16, 9, 19) {real, imag} */,
  {32'h3e7c7b59, 32'h3eb81228} /* (16, 9, 18) {real, imag} */,
  {32'h3e92a36e, 32'h3e872ae6} /* (16, 9, 17) {real, imag} */,
  {32'hbcaeb338, 32'h3e913a07} /* (16, 9, 16) {real, imag} */,
  {32'h3e601d24, 32'h3e8dc252} /* (16, 9, 15) {real, imag} */,
  {32'h3e795a54, 32'hbcf59184} /* (16, 9, 14) {real, imag} */,
  {32'hbe233aa7, 32'h3ce2496c} /* (16, 9, 13) {real, imag} */,
  {32'h3e3a1339, 32'h3e34a265} /* (16, 9, 12) {real, imag} */,
  {32'h3e8ed7ec, 32'h3e99cf89} /* (16, 9, 11) {real, imag} */,
  {32'hbf21ca96, 32'hbe999872} /* (16, 9, 10) {real, imag} */,
  {32'h3eb43dc9, 32'h3ec405ae} /* (16, 9, 9) {real, imag} */,
  {32'hbebe5da1, 32'h3e23af6b} /* (16, 9, 8) {real, imag} */,
  {32'h3f1af1cb, 32'h3e4793c6} /* (16, 9, 7) {real, imag} */,
  {32'h3f0ab3b2, 32'hbf389c90} /* (16, 9, 6) {real, imag} */,
  {32'h3d49154b, 32'hbc094d40} /* (16, 9, 5) {real, imag} */,
  {32'hbea93bb8, 32'h3eac3dab} /* (16, 9, 4) {real, imag} */,
  {32'h3d9851d6, 32'hbb9e1d80} /* (16, 9, 3) {real, imag} */,
  {32'hbed95fe8, 32'h3f594b4e} /* (16, 9, 2) {real, imag} */,
  {32'hbe8f69c9, 32'hbe61725c} /* (16, 9, 1) {real, imag} */,
  {32'h3e81cf3d, 32'hbf00fb34} /* (16, 9, 0) {real, imag} */,
  {32'h3e792d32, 32'h3f8e7938} /* (16, 8, 31) {real, imag} */,
  {32'hbf3e68b2, 32'hbeefd801} /* (16, 8, 30) {real, imag} */,
  {32'hbee85e3a, 32'hbc69b080} /* (16, 8, 29) {real, imag} */,
  {32'h3e5f0298, 32'hbf01a8fe} /* (16, 8, 28) {real, imag} */,
  {32'hbe97b41f, 32'h3cad34ac} /* (16, 8, 27) {real, imag} */,
  {32'hbf88a4fb, 32'h3f0385de} /* (16, 8, 26) {real, imag} */,
  {32'h3b95fc60, 32'hbe96bd29} /* (16, 8, 25) {real, imag} */,
  {32'hbf3b4e97, 32'hbd617ca0} /* (16, 8, 24) {real, imag} */,
  {32'h3f152c9a, 32'hbe04102d} /* (16, 8, 23) {real, imag} */,
  {32'hbeb4f0c2, 32'hbf0589df} /* (16, 8, 22) {real, imag} */,
  {32'h3b831f10, 32'h3e8b4763} /* (16, 8, 21) {real, imag} */,
  {32'hbdedd372, 32'h3dfafdcc} /* (16, 8, 20) {real, imag} */,
  {32'hbf0f07fa, 32'hbeef5374} /* (16, 8, 19) {real, imag} */,
  {32'h3e49b438, 32'h3ea4083c} /* (16, 8, 18) {real, imag} */,
  {32'h3da51ffb, 32'hbcc16e2a} /* (16, 8, 17) {real, imag} */,
  {32'hbd75c088, 32'h3e6756d5} /* (16, 8, 16) {real, imag} */,
  {32'h3ee36aee, 32'h3e3147ac} /* (16, 8, 15) {real, imag} */,
  {32'hbe09583c, 32'h3e99f0ed} /* (16, 8, 14) {real, imag} */,
  {32'hbe2bf8c2, 32'h3ccaca60} /* (16, 8, 13) {real, imag} */,
  {32'h3ec6f27e, 32'h3d893d4e} /* (16, 8, 12) {real, imag} */,
  {32'hbedff4e4, 32'h3ebcdc1a} /* (16, 8, 11) {real, imag} */,
  {32'hbec03fbe, 32'h3e4652de} /* (16, 8, 10) {real, imag} */,
  {32'h3eb1c973, 32'h3da1db98} /* (16, 8, 9) {real, imag} */,
  {32'hbd9cbd02, 32'hbef0eb11} /* (16, 8, 8) {real, imag} */,
  {32'hbe999166, 32'h3f081508} /* (16, 8, 7) {real, imag} */,
  {32'h3ee302e4, 32'hbf1518b9} /* (16, 8, 6) {real, imag} */,
  {32'h3ebde063, 32'hbefb5a17} /* (16, 8, 5) {real, imag} */,
  {32'h3d475044, 32'hbf20916d} /* (16, 8, 4) {real, imag} */,
  {32'hbe900690, 32'h3eaa6a21} /* (16, 8, 3) {real, imag} */,
  {32'hbe62054c, 32'h3d675f36} /* (16, 8, 2) {real, imag} */,
  {32'h3f3afc54, 32'h3f719911} /* (16, 8, 1) {real, imag} */,
  {32'h3ef4daed, 32'h3e96a838} /* (16, 8, 0) {real, imag} */,
  {32'h3d73a648, 32'h3f83c1b0} /* (16, 7, 31) {real, imag} */,
  {32'h3ed938be, 32'hbf3f75e4} /* (16, 7, 30) {real, imag} */,
  {32'hbf3d531a, 32'hbc708240} /* (16, 7, 29) {real, imag} */,
  {32'hbefebc5e, 32'h3e617932} /* (16, 7, 28) {real, imag} */,
  {32'hbdac55ef, 32'hbcc2a76c} /* (16, 7, 27) {real, imag} */,
  {32'h3e1d4e34, 32'hbe0a75e8} /* (16, 7, 26) {real, imag} */,
  {32'hbe5da323, 32'hbdbba25a} /* (16, 7, 25) {real, imag} */,
  {32'hbd81e20f, 32'h3b2cad80} /* (16, 7, 24) {real, imag} */,
  {32'h3ef3b8a2, 32'h3e6d1bb8} /* (16, 7, 23) {real, imag} */,
  {32'h3e4c6de2, 32'hbe747b89} /* (16, 7, 22) {real, imag} */,
  {32'h3e8dc0ac, 32'h3e36abdc} /* (16, 7, 21) {real, imag} */,
  {32'hbf2d22ab, 32'h3e0904e0} /* (16, 7, 20) {real, imag} */,
  {32'h3e0fc175, 32'hbf3d2980} /* (16, 7, 19) {real, imag} */,
  {32'hbe3cd34b, 32'hbe5c146b} /* (16, 7, 18) {real, imag} */,
  {32'hbe6a4d8c, 32'hbd891450} /* (16, 7, 17) {real, imag} */,
  {32'h3e691d02, 32'hbe283555} /* (16, 7, 16) {real, imag} */,
  {32'hbef7365a, 32'h3e763554} /* (16, 7, 15) {real, imag} */,
  {32'h3e8f3f86, 32'h3d5f0ce2} /* (16, 7, 14) {real, imag} */,
  {32'hbe967886, 32'hbed72bce} /* (16, 7, 13) {real, imag} */,
  {32'hbe67da49, 32'hbcebe698} /* (16, 7, 12) {real, imag} */,
  {32'h3e9cb243, 32'hbeedec23} /* (16, 7, 11) {real, imag} */,
  {32'h3d664f44, 32'h3ec6108e} /* (16, 7, 10) {real, imag} */,
  {32'hbe348c16, 32'hbe9f5a90} /* (16, 7, 9) {real, imag} */,
  {32'hbec81bec, 32'hbd1ca6bc} /* (16, 7, 8) {real, imag} */,
  {32'h3db8b28d, 32'hbd4c36d8} /* (16, 7, 7) {real, imag} */,
  {32'hbe74ca63, 32'hbe788243} /* (16, 7, 6) {real, imag} */,
  {32'h3e454229, 32'h3e87814e} /* (16, 7, 5) {real, imag} */,
  {32'h3f1a940c, 32'h3e3e27ed} /* (16, 7, 4) {real, imag} */,
  {32'hbda5b60c, 32'hbde97c23} /* (16, 7, 3) {real, imag} */,
  {32'h3e95fb1a, 32'hbee41866} /* (16, 7, 2) {real, imag} */,
  {32'hbf8e2258, 32'h3ec12336} /* (16, 7, 1) {real, imag} */,
  {32'hbdab7490, 32'hbeb21a3c} /* (16, 7, 0) {real, imag} */,
  {32'h3eea83e1, 32'h3d8e69cc} /* (16, 6, 31) {real, imag} */,
  {32'hbf634a9f, 32'h3dd31000} /* (16, 6, 30) {real, imag} */,
  {32'h3cecebe4, 32'hbf46318b} /* (16, 6, 29) {real, imag} */,
  {32'hbe839244, 32'h3eb650b5} /* (16, 6, 28) {real, imag} */,
  {32'hb9c17c00, 32'h3deafc42} /* (16, 6, 27) {real, imag} */,
  {32'hbd9ebc74, 32'hbdd12764} /* (16, 6, 26) {real, imag} */,
  {32'h3dde029e, 32'h3f0cbda7} /* (16, 6, 25) {real, imag} */,
  {32'h3d9fc3c1, 32'hbee846a6} /* (16, 6, 24) {real, imag} */,
  {32'hbe6b0490, 32'h3d319bc0} /* (16, 6, 23) {real, imag} */,
  {32'h3e5c52dc, 32'hbd73cbfc} /* (16, 6, 22) {real, imag} */,
  {32'hbc2f36b0, 32'h3e0860fc} /* (16, 6, 21) {real, imag} */,
  {32'hbd35a018, 32'hbf385db2} /* (16, 6, 20) {real, imag} */,
  {32'h3e78964e, 32'h3d2533bf} /* (16, 6, 19) {real, imag} */,
  {32'hbda05ba6, 32'hbf101716} /* (16, 6, 18) {real, imag} */,
  {32'h3e47ac93, 32'h3c9e9f4a} /* (16, 6, 17) {real, imag} */,
  {32'hbd8b14c0, 32'hbd703d4a} /* (16, 6, 16) {real, imag} */,
  {32'h3e2bb11d, 32'h3e81672d} /* (16, 6, 15) {real, imag} */,
  {32'h3ecf250a, 32'h3e2e7ffe} /* (16, 6, 14) {real, imag} */,
  {32'h3ebacf5e, 32'hbf043cfb} /* (16, 6, 13) {real, imag} */,
  {32'h3ec3dae3, 32'hbc315270} /* (16, 6, 12) {real, imag} */,
  {32'hbeddf51b, 32'h3e98e706} /* (16, 6, 11) {real, imag} */,
  {32'hbf248c5d, 32'h3dadc1ac} /* (16, 6, 10) {real, imag} */,
  {32'h3bac44e0, 32'hbd2d4c3c} /* (16, 6, 9) {real, imag} */,
  {32'hbd91c108, 32'hbf003afc} /* (16, 6, 8) {real, imag} */,
  {32'h3f2f4862, 32'h3d6719f8} /* (16, 6, 7) {real, imag} */,
  {32'h3df8c06a, 32'h3b89c6b0} /* (16, 6, 6) {real, imag} */,
  {32'hbdb50853, 32'hbe1c36f4} /* (16, 6, 5) {real, imag} */,
  {32'h3d2327c0, 32'h3f30f047} /* (16, 6, 4) {real, imag} */,
  {32'h3e160241, 32'h3e6e1746} /* (16, 6, 3) {real, imag} */,
  {32'h3ec9149e, 32'hbdfbba58} /* (16, 6, 2) {real, imag} */,
  {32'h3f1c7b22, 32'h3dbcc0b0} /* (16, 6, 1) {real, imag} */,
  {32'hbee4373a, 32'hbf47785a} /* (16, 6, 0) {real, imag} */,
  {32'h3fd146f0, 32'h3f6ab79a} /* (16, 5, 31) {real, imag} */,
  {32'hbf5de820, 32'hbf5ae196} /* (16, 5, 30) {real, imag} */,
  {32'h3eb18f0c, 32'h3f52cc37} /* (16, 5, 29) {real, imag} */,
  {32'h3d9dce72, 32'h3edb7df2} /* (16, 5, 28) {real, imag} */,
  {32'h3dddb322, 32'h3f26a638} /* (16, 5, 27) {real, imag} */,
  {32'hbde144db, 32'h3f05ebf2} /* (16, 5, 26) {real, imag} */,
  {32'hbe54e649, 32'hbe434098} /* (16, 5, 25) {real, imag} */,
  {32'hbf394790, 32'h3ec29a9f} /* (16, 5, 24) {real, imag} */,
  {32'hbe83a542, 32'h3d58a9e8} /* (16, 5, 23) {real, imag} */,
  {32'h3c9b9680, 32'h3ebb0653} /* (16, 5, 22) {real, imag} */,
  {32'hbe0bab9e, 32'hbe514531} /* (16, 5, 21) {real, imag} */,
  {32'hbeab2d92, 32'h3d0b64e0} /* (16, 5, 20) {real, imag} */,
  {32'h3bfdb080, 32'hbeb0760e} /* (16, 5, 19) {real, imag} */,
  {32'h3daf3984, 32'hbd2b52b8} /* (16, 5, 18) {real, imag} */,
  {32'h3d484a76, 32'h3d00c8e1} /* (16, 5, 17) {real, imag} */,
  {32'hbeae3380, 32'h3e8d46b1} /* (16, 5, 16) {real, imag} */,
  {32'hbe9c228f, 32'h3eabbf3b} /* (16, 5, 15) {real, imag} */,
  {32'h3e893b1a, 32'hbdeac28b} /* (16, 5, 14) {real, imag} */,
  {32'hbd851cda, 32'hbdea0f04} /* (16, 5, 13) {real, imag} */,
  {32'h3eee77ad, 32'h3e98a145} /* (16, 5, 12) {real, imag} */,
  {32'h3f0f13c0, 32'h3e818f4d} /* (16, 5, 11) {real, imag} */,
  {32'hbe841c64, 32'hbf4378ea} /* (16, 5, 10) {real, imag} */,
  {32'hbef8c88c, 32'h3d9e1b2a} /* (16, 5, 9) {real, imag} */,
  {32'h3e4e175e, 32'h3e9a4fe6} /* (16, 5, 8) {real, imag} */,
  {32'hbd1854b8, 32'h3f06caac} /* (16, 5, 7) {real, imag} */,
  {32'hbdcf8582, 32'h3e4f2bf4} /* (16, 5, 6) {real, imag} */,
  {32'hbf600008, 32'h3f5cbb5b} /* (16, 5, 5) {real, imag} */,
  {32'h3ed4b8f5, 32'h3ce32e98} /* (16, 5, 4) {real, imag} */,
  {32'hbea489dd, 32'hbd324d8c} /* (16, 5, 3) {real, imag} */,
  {32'hbdc6f4b8, 32'hbfb66d87} /* (16, 5, 2) {real, imag} */,
  {32'h3f20dc8e, 32'h3fdc1706} /* (16, 5, 1) {real, imag} */,
  {32'h3eb619bc, 32'h3fa4ad66} /* (16, 5, 0) {real, imag} */,
  {32'hbe7ef748, 32'hc00e53ee} /* (16, 4, 31) {real, imag} */,
  {32'h3f8f346b, 32'h3f47f420} /* (16, 4, 30) {real, imag} */,
  {32'hbda0bf02, 32'hbf9ae6e1} /* (16, 4, 29) {real, imag} */,
  {32'hbf9c27aa, 32'h3e7c8e5e} /* (16, 4, 28) {real, imag} */,
  {32'h3f14e39b, 32'h3e289d65} /* (16, 4, 27) {real, imag} */,
  {32'hbea59ff8, 32'h3e0d4d5f} /* (16, 4, 26) {real, imag} */,
  {32'hbf1cb690, 32'h3ab17400} /* (16, 4, 25) {real, imag} */,
  {32'h3f899a8e, 32'hbf38d4ff} /* (16, 4, 24) {real, imag} */,
  {32'h3dacfae6, 32'h3ce9bf10} /* (16, 4, 23) {real, imag} */,
  {32'h3de1fc82, 32'h3e05ff20} /* (16, 4, 22) {real, imag} */,
  {32'hbce4ad36, 32'hbe3aa582} /* (16, 4, 21) {real, imag} */,
  {32'hbd853f98, 32'h3e4c0c12} /* (16, 4, 20) {real, imag} */,
  {32'h3d24c4b0, 32'h3de4b6d6} /* (16, 4, 19) {real, imag} */,
  {32'h3e12e2e9, 32'h3da7d58e} /* (16, 4, 18) {real, imag} */,
  {32'hbe8576e6, 32'h3d0c59a6} /* (16, 4, 17) {real, imag} */,
  {32'hbe1e3c68, 32'hbe1ae6a6} /* (16, 4, 16) {real, imag} */,
  {32'h3e946a74, 32'hbdca939e} /* (16, 4, 15) {real, imag} */,
  {32'hbe241c75, 32'h3e4e2ff2} /* (16, 4, 14) {real, imag} */,
  {32'hbecb4da3, 32'h3e85ef57} /* (16, 4, 13) {real, imag} */,
  {32'h3df07691, 32'h3d8a6a56} /* (16, 4, 12) {real, imag} */,
  {32'hbe4b16fe, 32'hbe9ec8b7} /* (16, 4, 11) {real, imag} */,
  {32'h3f238449, 32'h3d894c7c} /* (16, 4, 10) {real, imag} */,
  {32'hbe9930da, 32'h3f01ad64} /* (16, 4, 9) {real, imag} */,
  {32'h3f11f692, 32'h3ead68be} /* (16, 4, 8) {real, imag} */,
  {32'hbf5b095a, 32'hbe160a48} /* (16, 4, 7) {real, imag} */,
  {32'hbea3d011, 32'hbea4bb9c} /* (16, 4, 6) {real, imag} */,
  {32'hbf0aae12, 32'h3e8239a2} /* (16, 4, 5) {real, imag} */,
  {32'hbe83fc49, 32'hbf57fa27} /* (16, 4, 4) {real, imag} */,
  {32'hbefd33a6, 32'hbe0b24d8} /* (16, 4, 3) {real, imag} */,
  {32'h3f976092, 32'h3ff8c2f9} /* (16, 4, 2) {real, imag} */,
  {32'hbf8ce2be, 32'hbf95a388} /* (16, 4, 1) {real, imag} */,
  {32'hc00acaa1, 32'hc016486a} /* (16, 4, 0) {real, imag} */,
  {32'h4055e0dc, 32'hbfd0b5ec} /* (16, 3, 31) {real, imag} */,
  {32'h3f2b2c82, 32'h40246962} /* (16, 3, 30) {real, imag} */,
  {32'hbf48b58a, 32'h3f179098} /* (16, 3, 29) {real, imag} */,
  {32'hbec6e227, 32'h3d3f4d74} /* (16, 3, 28) {real, imag} */,
  {32'h3ee191b8, 32'h3de68ad4} /* (16, 3, 27) {real, imag} */,
  {32'hbd988f58, 32'h3d2196b6} /* (16, 3, 26) {real, imag} */,
  {32'hbf3aa252, 32'h3f2bb9e5} /* (16, 3, 25) {real, imag} */,
  {32'hbe5cea7a, 32'hbd758794} /* (16, 3, 24) {real, imag} */,
  {32'hbed12ec5, 32'h3d978b56} /* (16, 3, 23) {real, imag} */,
  {32'h3c16ec70, 32'hbe40ba5d} /* (16, 3, 22) {real, imag} */,
  {32'h3ed02bdd, 32'h3d1431be} /* (16, 3, 21) {real, imag} */,
  {32'hbc218910, 32'h3deab9b7} /* (16, 3, 20) {real, imag} */,
  {32'hbd7f8368, 32'hbe81c5aa} /* (16, 3, 19) {real, imag} */,
  {32'hbcb5b548, 32'hbe323e14} /* (16, 3, 18) {real, imag} */,
  {32'hbe1ac3ce, 32'hbdb295e6} /* (16, 3, 17) {real, imag} */,
  {32'h3e14aec2, 32'h3e5777d5} /* (16, 3, 16) {real, imag} */,
  {32'h3ec8a698, 32'h3eaf8729} /* (16, 3, 15) {real, imag} */,
  {32'h3ecd49bd, 32'hbd7c036a} /* (16, 3, 14) {real, imag} */,
  {32'hbecd823d, 32'hbe3a483a} /* (16, 3, 13) {real, imag} */,
  {32'hbeb16220, 32'hbe7ecc8b} /* (16, 3, 12) {real, imag} */,
  {32'h3ee7c226, 32'hbe1fbefd} /* (16, 3, 11) {real, imag} */,
  {32'h3c6acb50, 32'hbf08e3c5} /* (16, 3, 10) {real, imag} */,
  {32'hbf0f8df1, 32'h3e687389} /* (16, 3, 9) {real, imag} */,
  {32'h3d82eb04, 32'hbf0226a3} /* (16, 3, 8) {real, imag} */,
  {32'hbe50444c, 32'hbe9b23b6} /* (16, 3, 7) {real, imag} */,
  {32'hbf0005d0, 32'h3e0311c2} /* (16, 3, 6) {real, imag} */,
  {32'hbf0e1e02, 32'h3e802733} /* (16, 3, 5) {real, imag} */,
  {32'h3f10803e, 32'h3f1d0864} /* (16, 3, 4) {real, imag} */,
  {32'h3e8cfc1b, 32'hbefdfa0d} /* (16, 3, 3) {real, imag} */,
  {32'h40171188, 32'h3f96f3d0} /* (16, 3, 2) {real, imag} */,
  {32'hbf826ac2, 32'hc023f852} /* (16, 3, 1) {real, imag} */,
  {32'h3f105f7a, 32'h3f24b14b} /* (16, 3, 0) {real, imag} */,
  {32'h4135b55c, 32'hbf882d55} /* (16, 2, 31) {real, imag} */,
  {32'hc0ab9d67, 32'h3f96c7cd} /* (16, 2, 30) {real, imag} */,
  {32'h4010f9ee, 32'h3f26bee2} /* (16, 2, 29) {real, imag} */,
  {32'h3f453ad6, 32'hbf3337ce} /* (16, 2, 28) {real, imag} */,
  {32'hbf7d5c0e, 32'h3f16de1c} /* (16, 2, 27) {real, imag} */,
  {32'h3e0f1896, 32'h3ee4c2ed} /* (16, 2, 26) {real, imag} */,
  {32'h3f535b7e, 32'hbf944c77} /* (16, 2, 25) {real, imag} */,
  {32'hbf885792, 32'h3ed66ed8} /* (16, 2, 24) {real, imag} */,
  {32'hbecc89d3, 32'h3f0cc3a5} /* (16, 2, 23) {real, imag} */,
  {32'hbdcedfa3, 32'hbe4a6495} /* (16, 2, 22) {real, imag} */,
  {32'h3b824e20, 32'h3f40d919} /* (16, 2, 21) {real, imag} */,
  {32'h3e36fcaa, 32'hbe07d80a} /* (16, 2, 20) {real, imag} */,
  {32'hbeb4a8cc, 32'hbcb6c77e} /* (16, 2, 19) {real, imag} */,
  {32'hbda9ca0b, 32'hbc43d998} /* (16, 2, 18) {real, imag} */,
  {32'hbe854dc6, 32'hbdcb1777} /* (16, 2, 17) {real, imag} */,
  {32'hbdb2db5d, 32'h3e2ae302} /* (16, 2, 16) {real, imag} */,
  {32'hbec2b1cf, 32'h3daeceec} /* (16, 2, 15) {real, imag} */,
  {32'hbe80a7b6, 32'hbeb63e1f} /* (16, 2, 14) {real, imag} */,
  {32'h3e083189, 32'h3ea95024} /* (16, 2, 13) {real, imag} */,
  {32'hbf32f796, 32'h3e8b6330} /* (16, 2, 12) {real, imag} */,
  {32'h3cece7e8, 32'hbeb3794e} /* (16, 2, 11) {real, imag} */,
  {32'hbe69d6d9, 32'h3e9f7780} /* (16, 2, 10) {real, imag} */,
  {32'hbeb75fee, 32'h3ec13fc8} /* (16, 2, 9) {real, imag} */,
  {32'hbd089ec0, 32'hbf1e9816} /* (16, 2, 8) {real, imag} */,
  {32'h3e815ed4, 32'hbf28dbae} /* (16, 2, 7) {real, imag} */,
  {32'h3ec60f24, 32'h3f886788} /* (16, 2, 6) {real, imag} */,
  {32'hbfa7d671, 32'hbf85cc47} /* (16, 2, 5) {real, imag} */,
  {32'h400cd20f, 32'hbffba005} /* (16, 2, 4) {real, imag} */,
  {32'h3fce23a5, 32'hbf88953e} /* (16, 2, 3) {real, imag} */,
  {32'hc0935ae8, 32'h3fd57096} /* (16, 2, 2) {real, imag} */,
  {32'h40d25d58, 32'hc0074e32} /* (16, 2, 1) {real, imag} */,
  {32'h40a463d3, 32'h4009471a} /* (16, 2, 0) {real, imag} */,
  {32'hc129e471, 32'h3f77d62e} /* (16, 1, 31) {real, imag} */,
  {32'h404eb9cb, 32'hbfad3df8} /* (16, 1, 30) {real, imag} */,
  {32'hbe262fb2, 32'h3f961134} /* (16, 1, 29) {real, imag} */,
  {32'hbf67daa7, 32'hbfffb5b5} /* (16, 1, 28) {real, imag} */,
  {32'h402c0bc7, 32'hbdef9e22} /* (16, 1, 27) {real, imag} */,
  {32'h3f9fb484, 32'hbcbe6d20} /* (16, 1, 26) {real, imag} */,
  {32'hbea2288c, 32'h3eb17902} /* (16, 1, 25) {real, imag} */,
  {32'hbc1a22b0, 32'hbecca71f} /* (16, 1, 24) {real, imag} */,
  {32'hbec7fb94, 32'h3ee1bd66} /* (16, 1, 23) {real, imag} */,
  {32'hbe15f084, 32'h3e565155} /* (16, 1, 22) {real, imag} */,
  {32'hbd005608, 32'hbf304976} /* (16, 1, 21) {real, imag} */,
  {32'h3e4597a8, 32'hbec96438} /* (16, 1, 20) {real, imag} */,
  {32'h3bd71d80, 32'h3ed0cc18} /* (16, 1, 19) {real, imag} */,
  {32'h3d8488e8, 32'h3e44c194} /* (16, 1, 18) {real, imag} */,
  {32'hbebd88f8, 32'hbde59aef} /* (16, 1, 17) {real, imag} */,
  {32'hbe443076, 32'h3eb151b0} /* (16, 1, 16) {real, imag} */,
  {32'hbcb8b92c, 32'h3e152676} /* (16, 1, 15) {real, imag} */,
  {32'hbcac29cc, 32'h3e64d42a} /* (16, 1, 14) {real, imag} */,
  {32'h3c3a93a8, 32'h3dd7d8c8} /* (16, 1, 13) {real, imag} */,
  {32'hbe8bd5c4, 32'hbf2a38c2} /* (16, 1, 12) {real, imag} */,
  {32'h3df54fc6, 32'h3f4f6f50} /* (16, 1, 11) {real, imag} */,
  {32'h3e078c98, 32'h3de1d634} /* (16, 1, 10) {real, imag} */,
  {32'h3e928433, 32'h3e7fd64c} /* (16, 1, 9) {real, imag} */,
  {32'h3e7e7128, 32'h3f3d5189} /* (16, 1, 8) {real, imag} */,
  {32'hbd8f8e26, 32'hbf20ac28} /* (16, 1, 7) {real, imag} */,
  {32'hbe10c21a, 32'h3f1679ee} /* (16, 1, 6) {real, imag} */,
  {32'h3ff660e2, 32'h3f7518ce} /* (16, 1, 5) {real, imag} */,
  {32'hbfba5c66, 32'hbea49777} /* (16, 1, 4) {real, imag} */,
  {32'hbf7ee1ff, 32'h3eba5880} /* (16, 1, 3) {real, imag} */,
  {32'h40803086, 32'h40d42f73} /* (16, 1, 2) {real, imag} */,
  {32'hc196a040, 32'hc0f0ba5d} /* (16, 1, 1) {real, imag} */,
  {32'hc15bf39e, 32'hc0d6e162} /* (16, 1, 0) {real, imag} */,
  {32'hc1620ab6, 32'h4110a64a} /* (16, 0, 31) {real, imag} */,
  {32'h3f742fc5, 32'hc0473f5d} /* (16, 0, 30) {real, imag} */,
  {32'h3f7e0f7d, 32'h3e8ad063} /* (16, 0, 29) {real, imag} */,
  {32'hbf37660c, 32'hbf8cbb86} /* (16, 0, 28) {real, imag} */,
  {32'h3ec6f808, 32'h3da514b8} /* (16, 0, 27) {real, imag} */,
  {32'h3edda8ad, 32'hbed62bfb} /* (16, 0, 26) {real, imag} */,
  {32'h3e0ac698, 32'hbe5b7eea} /* (16, 0, 25) {real, imag} */,
  {32'h3e552678, 32'hbe2db9b2} /* (16, 0, 24) {real, imag} */,
  {32'h3f145767, 32'hbe464972} /* (16, 0, 23) {real, imag} */,
  {32'hbcd8ca10, 32'h3c749bc0} /* (16, 0, 22) {real, imag} */,
  {32'h3d80c83c, 32'hbe4cbe07} /* (16, 0, 21) {real, imag} */,
  {32'h3e55eba4, 32'h3c5eb5b0} /* (16, 0, 20) {real, imag} */,
  {32'hbe045d26, 32'h3d063b3b} /* (16, 0, 19) {real, imag} */,
  {32'hbec611c8, 32'h3d3b0930} /* (16, 0, 18) {real, imag} */,
  {32'h3dd03e54, 32'hbe6ab21c} /* (16, 0, 17) {real, imag} */,
  {32'hbd8d19a7, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h3dd03e54, 32'h3e6ab21c} /* (16, 0, 15) {real, imag} */,
  {32'hbec611c8, 32'hbd3b0930} /* (16, 0, 14) {real, imag} */,
  {32'hbe045d26, 32'hbd063b3b} /* (16, 0, 13) {real, imag} */,
  {32'h3e55eba4, 32'hbc5eb5b0} /* (16, 0, 12) {real, imag} */,
  {32'h3d80c83c, 32'h3e4cbe07} /* (16, 0, 11) {real, imag} */,
  {32'hbcd8ca10, 32'hbc749bc0} /* (16, 0, 10) {real, imag} */,
  {32'h3f145767, 32'h3e464972} /* (16, 0, 9) {real, imag} */,
  {32'h3e552678, 32'h3e2db9b2} /* (16, 0, 8) {real, imag} */,
  {32'h3e0ac698, 32'h3e5b7eea} /* (16, 0, 7) {real, imag} */,
  {32'h3edda8ad, 32'h3ed62bfb} /* (16, 0, 6) {real, imag} */,
  {32'h3ec6f808, 32'hbda514b8} /* (16, 0, 5) {real, imag} */,
  {32'hbf37660c, 32'h3f8cbb86} /* (16, 0, 4) {real, imag} */,
  {32'h3f7e0f7d, 32'hbe8ad063} /* (16, 0, 3) {real, imag} */,
  {32'h3f742fc5, 32'h40473f5d} /* (16, 0, 2) {real, imag} */,
  {32'hc1620ab6, 32'hc110a64a} /* (16, 0, 1) {real, imag} */,
  {32'hc1420fa8, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h415eba7e, 32'hc1276652} /* (15, 31, 31) {real, imag} */,
  {32'hc0d82234, 32'h40879866} /* (15, 31, 30) {real, imag} */,
  {32'hbffe0c61, 32'hbe6f4938} /* (15, 31, 29) {real, imag} */,
  {32'hbf40ee98, 32'hbfb0abe2} /* (15, 31, 28) {real, imag} */,
  {32'hbec70a0a, 32'h3ea39f68} /* (15, 31, 27) {real, imag} */,
  {32'h3edd400e, 32'h3ef7816f} /* (15, 31, 26) {real, imag} */,
  {32'h3f636749, 32'hbeb3a78e} /* (15, 31, 25) {real, imag} */,
  {32'hbf1c2dfb, 32'h3f215b96} /* (15, 31, 24) {real, imag} */,
  {32'h3caa78da, 32'hbe32ed53} /* (15, 31, 23) {real, imag} */,
  {32'h3d8bcd7e, 32'h3e8aad7a} /* (15, 31, 22) {real, imag} */,
  {32'hbe7318b2, 32'h3cd2feb0} /* (15, 31, 21) {real, imag} */,
  {32'hbe862490, 32'h3f133f61} /* (15, 31, 20) {real, imag} */,
  {32'h3ef7cc9e, 32'h3d10055a} /* (15, 31, 19) {real, imag} */,
  {32'h3ebef1c5, 32'h3e6f4662} /* (15, 31, 18) {real, imag} */,
  {32'hbe7a9b04, 32'hbe8faaf0} /* (15, 31, 17) {real, imag} */,
  {32'h3e2a6adf, 32'h3f0bfdf0} /* (15, 31, 16) {real, imag} */,
  {32'h3eaa92c4, 32'h3dd62f48} /* (15, 31, 15) {real, imag} */,
  {32'hbdd63de8, 32'hbe8bc191} /* (15, 31, 14) {real, imag} */,
  {32'h3e426fe1, 32'hbf187dd0} /* (15, 31, 13) {real, imag} */,
  {32'h3ee0bff3, 32'h3d4bd704} /* (15, 31, 12) {real, imag} */,
  {32'hbef64074, 32'hbe83b3d4} /* (15, 31, 11) {real, imag} */,
  {32'h3f07daa9, 32'h3e27086c} /* (15, 31, 10) {real, imag} */,
  {32'hbec3235a, 32'hbf07b618} /* (15, 31, 9) {real, imag} */,
  {32'hbec9a74e, 32'hbeb5d01a} /* (15, 31, 8) {real, imag} */,
  {32'hbd90a002, 32'hbeea7351} /* (15, 31, 7) {real, imag} */,
  {32'h3f573571, 32'h3ef115ce} /* (15, 31, 6) {real, imag} */,
  {32'hbfb10238, 32'hbf34d6e6} /* (15, 31, 5) {real, imag} */,
  {32'h3fc58192, 32'h3f199196} /* (15, 31, 4) {real, imag} */,
  {32'hbe40fadc, 32'hbfff0978} /* (15, 31, 3) {real, imag} */,
  {32'hc0904efa, 32'h3f98cc8b} /* (15, 31, 2) {real, imag} */,
  {32'h41560f50, 32'h40886eb9} /* (15, 31, 1) {real, imag} */,
  {32'h4154b47b, 32'h404e2f16} /* (15, 31, 0) {real, imag} */,
  {32'hc09dbeae, 32'h3f2a6c18} /* (15, 30, 31) {real, imag} */,
  {32'h406c5e68, 32'h3eb12d1c} /* (15, 30, 30) {real, imag} */,
  {32'h3f2b8b3f, 32'h3e8a9278} /* (15, 30, 29) {real, imag} */,
  {32'h3e69a620, 32'h3ffa85c9} /* (15, 30, 28) {real, imag} */,
  {32'h3f3fdd0d, 32'hbfa79d04} /* (15, 30, 27) {real, imag} */,
  {32'h3da0a6df, 32'hbee4eab7} /* (15, 30, 26) {real, imag} */,
  {32'hbbaab738, 32'hbe532c30} /* (15, 30, 25) {real, imag} */,
  {32'h3f718c62, 32'hbd718db0} /* (15, 30, 24) {real, imag} */,
  {32'hbe8bf8c0, 32'hbe805efe} /* (15, 30, 23) {real, imag} */,
  {32'hbf0bedac, 32'h3e865a68} /* (15, 30, 22) {real, imag} */,
  {32'hbead1c62, 32'hbe90aedd} /* (15, 30, 21) {real, imag} */,
  {32'h3e0e462c, 32'hbec86628} /* (15, 30, 20) {real, imag} */,
  {32'h3e140144, 32'h3d30bfba} /* (15, 30, 19) {real, imag} */,
  {32'h3e3c4161, 32'hbef96a64} /* (15, 30, 18) {real, imag} */,
  {32'h3c63c278, 32'h3e0d37ae} /* (15, 30, 17) {real, imag} */,
  {32'hbe3b5706, 32'h3e5d9872} /* (15, 30, 16) {real, imag} */,
  {32'hbd766c02, 32'h3dc8f7fe} /* (15, 30, 15) {real, imag} */,
  {32'h3d422708, 32'hbe0be652} /* (15, 30, 14) {real, imag} */,
  {32'hbe4ee376, 32'hbea2f9d4} /* (15, 30, 13) {real, imag} */,
  {32'hbe7b40f8, 32'h3c309e00} /* (15, 30, 12) {real, imag} */,
  {32'h3cee42e8, 32'h3e7aeb06} /* (15, 30, 11) {real, imag} */,
  {32'h3e5e441a, 32'h3e44be1e} /* (15, 30, 10) {real, imag} */,
  {32'hbed177fa, 32'hbef1ec78} /* (15, 30, 9) {real, imag} */,
  {32'h3f012e38, 32'h3fb8869f} /* (15, 30, 8) {real, imag} */,
  {32'hbe36ed96, 32'hbe156dc5} /* (15, 30, 7) {real, imag} */,
  {32'hbf3bffd0, 32'hbf8c132a} /* (15, 30, 6) {real, imag} */,
  {32'h3e83ec76, 32'h3e696154} /* (15, 30, 5) {real, imag} */,
  {32'hbf23d818, 32'hbfd85694} /* (15, 30, 4) {real, imag} */,
  {32'h3f80f102, 32'hbf8c7ea2} /* (15, 30, 3) {real, imag} */,
  {32'h40ba0394, 32'h3f94978c} /* (15, 30, 2) {real, imag} */,
  {32'hc11cc5a7, 32'h401cc922} /* (15, 30, 1) {real, imag} */,
  {32'hc0c446ee, 32'hbde18e20} /* (15, 30, 0) {real, imag} */,
  {32'h3fe87e13, 32'hbe20f4f0} /* (15, 29, 31) {real, imag} */,
  {32'h3ec5a74e, 32'h3fa00cd7} /* (15, 29, 30) {real, imag} */,
  {32'h3e1d4050, 32'hbef75db8} /* (15, 29, 29) {real, imag} */,
  {32'hbf12c4f2, 32'hbf6c8acc} /* (15, 29, 28) {real, imag} */,
  {32'h3ebb5d54, 32'hbec3e139} /* (15, 29, 27) {real, imag} */,
  {32'hbe0373ec, 32'hbe4f5ec6} /* (15, 29, 26) {real, imag} */,
  {32'hbea05b99, 32'h3e81857c} /* (15, 29, 25) {real, imag} */,
  {32'h3e073249, 32'h3e54793f} /* (15, 29, 24) {real, imag} */,
  {32'hbeb71e38, 32'hbcf0825c} /* (15, 29, 23) {real, imag} */,
  {32'hbe179c0c, 32'hbe199ac6} /* (15, 29, 22) {real, imag} */,
  {32'hbea7e2a5, 32'hbe9a2dd3} /* (15, 29, 21) {real, imag} */,
  {32'h3e11e365, 32'h3e3995d2} /* (15, 29, 20) {real, imag} */,
  {32'h3e88c562, 32'hbeb3722d} /* (15, 29, 19) {real, imag} */,
  {32'hbca1b824, 32'hbd0a287a} /* (15, 29, 18) {real, imag} */,
  {32'hbe617484, 32'h3de14d6d} /* (15, 29, 17) {real, imag} */,
  {32'hbcd99f38, 32'h3e0d8b9c} /* (15, 29, 16) {real, imag} */,
  {32'h3d42587c, 32'hbef8e007} /* (15, 29, 15) {real, imag} */,
  {32'h3dd418f0, 32'h3ed54048} /* (15, 29, 14) {real, imag} */,
  {32'hbd585dc6, 32'h3ee7f592} /* (15, 29, 13) {real, imag} */,
  {32'hbe60f4ea, 32'hbf38a196} /* (15, 29, 12) {real, imag} */,
  {32'hbdd7112c, 32'h3e95ea64} /* (15, 29, 11) {real, imag} */,
  {32'h3eabe82a, 32'h3e26f92a} /* (15, 29, 10) {real, imag} */,
  {32'hbf0bfd10, 32'hbe530932} /* (15, 29, 9) {real, imag} */,
  {32'hbef76c19, 32'h3ebfae00} /* (15, 29, 8) {real, imag} */,
  {32'hbf2fa7cf, 32'hbcee18a0} /* (15, 29, 7) {real, imag} */,
  {32'hbc49b4c0, 32'hbf387748} /* (15, 29, 6) {real, imag} */,
  {32'hbe5d8e40, 32'hbeac4008} /* (15, 29, 5) {real, imag} */,
  {32'h3f4f13ec, 32'hbef940f6} /* (15, 29, 4) {real, imag} */,
  {32'hbf571ca0, 32'h3e8c5562} /* (15, 29, 3) {real, imag} */,
  {32'h3fb7d485, 32'h3f1d1ab0} /* (15, 29, 2) {real, imag} */,
  {32'h3f035fde, 32'h3ab97800} /* (15, 29, 1) {real, imag} */,
  {32'h3ead938e, 32'hbf745722} /* (15, 29, 0) {real, imag} */,
  {32'h4047996a, 32'hbf1f55d5} /* (15, 28, 31) {real, imag} */,
  {32'hbebdcab8, 32'h3fb6e4eb} /* (15, 28, 30) {real, imag} */,
  {32'hbf0ee141, 32'hbf3c9308} /* (15, 28, 29) {real, imag} */,
  {32'hbf04f422, 32'hbeac464b} /* (15, 28, 28) {real, imag} */,
  {32'hbf3be5f9, 32'h3ed232e4} /* (15, 28, 27) {real, imag} */,
  {32'hbf413c7e, 32'h3f3b5633} /* (15, 28, 26) {real, imag} */,
  {32'h3ebdc926, 32'hbf673398} /* (15, 28, 25) {real, imag} */,
  {32'hbec52cb2, 32'h3e4349f0} /* (15, 28, 24) {real, imag} */,
  {32'h3e34424c, 32'h3e454cbd} /* (15, 28, 23) {real, imag} */,
  {32'h3ef0a6e2, 32'h3f06eef5} /* (15, 28, 22) {real, imag} */,
  {32'h3ec0b383, 32'hbe36149a} /* (15, 28, 21) {real, imag} */,
  {32'h3d0ee8b4, 32'hbdaaff94} /* (15, 28, 20) {real, imag} */,
  {32'h3ec316b5, 32'hbd707f50} /* (15, 28, 19) {real, imag} */,
  {32'hbe63e2d4, 32'h3e3d7ebd} /* (15, 28, 18) {real, imag} */,
  {32'hbe02eb07, 32'hbf0e0cb9} /* (15, 28, 17) {real, imag} */,
  {32'hbe591c69, 32'h3e36950c} /* (15, 28, 16) {real, imag} */,
  {32'h3d92a4c6, 32'h3e2a39e5} /* (15, 28, 15) {real, imag} */,
  {32'h3e4b6a14, 32'h3e4a8c5e} /* (15, 28, 14) {real, imag} */,
  {32'hbeee9b47, 32'hbe2cf6d6} /* (15, 28, 13) {real, imag} */,
  {32'hbbac5b70, 32'h3e4ebf23} /* (15, 28, 12) {real, imag} */,
  {32'h3cab2f62, 32'h3e28e580} /* (15, 28, 11) {real, imag} */,
  {32'hbd074bb6, 32'h3e47aa4c} /* (15, 28, 10) {real, imag} */,
  {32'hbe234b2e, 32'h3d684f6e} /* (15, 28, 9) {real, imag} */,
  {32'h3de33658, 32'h3c19cdc0} /* (15, 28, 8) {real, imag} */,
  {32'hbe8e1cb0, 32'hbf94df92} /* (15, 28, 7) {real, imag} */,
  {32'hbe910838, 32'hbf0d1f41} /* (15, 28, 6) {real, imag} */,
  {32'hbf220fc4, 32'hbe229844} /* (15, 28, 5) {real, imag} */,
  {32'h3f806e5c, 32'hbf14af2e} /* (15, 28, 4) {real, imag} */,
  {32'h3db725e0, 32'h3f1e83b8} /* (15, 28, 3) {real, imag} */,
  {32'hbf1e6d60, 32'h3f16f5ba} /* (15, 28, 2) {real, imag} */,
  {32'h3f9d9fbc, 32'hbd372c80} /* (15, 28, 1) {real, imag} */,
  {32'hbf5c134a, 32'h3f98548b} /* (15, 28, 0) {real, imag} */,
  {32'hbfd54f7e, 32'h3eb74c58} /* (15, 27, 31) {real, imag} */,
  {32'h3e9b8e68, 32'hbf1f5f70} /* (15, 27, 30) {real, imag} */,
  {32'h3f1041b0, 32'h3f15d2e4} /* (15, 27, 29) {real, imag} */,
  {32'h3f229328, 32'h3eb1d82c} /* (15, 27, 28) {real, imag} */,
  {32'h3e94528c, 32'hbe7739e2} /* (15, 27, 27) {real, imag} */,
  {32'h3e7ec830, 32'h3cf07600} /* (15, 27, 26) {real, imag} */,
  {32'hbe0fb8ea, 32'h3da0ec10} /* (15, 27, 25) {real, imag} */,
  {32'h3e237cce, 32'hbf4a2ad7} /* (15, 27, 24) {real, imag} */,
  {32'hbea5f42a, 32'h3ed96398} /* (15, 27, 23) {real, imag} */,
  {32'hbe1a2fca, 32'h3ec9022a} /* (15, 27, 22) {real, imag} */,
  {32'hbd93142e, 32'hbe6e9bb6} /* (15, 27, 21) {real, imag} */,
  {32'hbe0d3b8b, 32'h3e09d9dc} /* (15, 27, 20) {real, imag} */,
  {32'hbe9c9fae, 32'h3d23f114} /* (15, 27, 19) {real, imag} */,
  {32'hbeaa67df, 32'h3e23a5d1} /* (15, 27, 18) {real, imag} */,
  {32'h3efcbc4c, 32'hbd821428} /* (15, 27, 17) {real, imag} */,
  {32'hbe7eeb64, 32'h3d8219f4} /* (15, 27, 16) {real, imag} */,
  {32'hbe59b8a8, 32'h3ee9f82a} /* (15, 27, 15) {real, imag} */,
  {32'h3e456958, 32'h3d0869b4} /* (15, 27, 14) {real, imag} */,
  {32'hbd85f2a7, 32'h3d84c9bf} /* (15, 27, 13) {real, imag} */,
  {32'hbdb0c4dc, 32'h3e35ca5f} /* (15, 27, 12) {real, imag} */,
  {32'h3c258570, 32'hbd3f9576} /* (15, 27, 11) {real, imag} */,
  {32'h3e386be6, 32'h3ee881ec} /* (15, 27, 10) {real, imag} */,
  {32'hbea1cadc, 32'hbdc791d8} /* (15, 27, 9) {real, imag} */,
  {32'hbec6b8e2, 32'h3d65e3b4} /* (15, 27, 8) {real, imag} */,
  {32'hbfa48c64, 32'hbe42bd64} /* (15, 27, 7) {real, imag} */,
  {32'hbd14ffb4, 32'h3ea86480} /* (15, 27, 6) {real, imag} */,
  {32'h3ec65102, 32'hbf62d8af} /* (15, 27, 5) {real, imag} */,
  {32'h3dcd1a90, 32'hbcf79cb8} /* (15, 27, 4) {real, imag} */,
  {32'h3d3fdc1c, 32'hbf20c403} /* (15, 27, 3) {real, imag} */,
  {32'h3df7cc00, 32'h3edb8776} /* (15, 27, 2) {real, imag} */,
  {32'hbf91640a, 32'hbfbdcea6} /* (15, 27, 1) {real, imag} */,
  {32'hbfc179e4, 32'h3db8dc30} /* (15, 27, 0) {real, imag} */,
  {32'h3f277bff, 32'hbf55ce2e} /* (15, 26, 31) {real, imag} */,
  {32'h3f2767b2, 32'hbf034c19} /* (15, 26, 30) {real, imag} */,
  {32'h3ed64445, 32'hbe27c6c5} /* (15, 26, 29) {real, imag} */,
  {32'hbec32d5e, 32'hbe0defba} /* (15, 26, 28) {real, imag} */,
  {32'h3ec72324, 32'h3e80d02c} /* (15, 26, 27) {real, imag} */,
  {32'hbe3e2efe, 32'hbe97208e} /* (15, 26, 26) {real, imag} */,
  {32'hbe18c8d2, 32'hbcd44c94} /* (15, 26, 25) {real, imag} */,
  {32'hbf013df1, 32'h3e9cedeb} /* (15, 26, 24) {real, imag} */,
  {32'h3e9a7126, 32'hbe821f3a} /* (15, 26, 23) {real, imag} */,
  {32'hbe8c38f6, 32'hbf16ef9e} /* (15, 26, 22) {real, imag} */,
  {32'h3e32ad73, 32'hbe3177f8} /* (15, 26, 21) {real, imag} */,
  {32'h3da2c340, 32'hbe6fb8be} /* (15, 26, 20) {real, imag} */,
  {32'h3aba1ce0, 32'hbd559a68} /* (15, 26, 19) {real, imag} */,
  {32'h3d990b4e, 32'hbeb86f18} /* (15, 26, 18) {real, imag} */,
  {32'h3e80214b, 32'h3e1a8350} /* (15, 26, 17) {real, imag} */,
  {32'h3dafa00a, 32'hbef42f66} /* (15, 26, 16) {real, imag} */,
  {32'h3e2fda9a, 32'h3e3c33da} /* (15, 26, 15) {real, imag} */,
  {32'h3eaa8d6e, 32'h3e09ad78} /* (15, 26, 14) {real, imag} */,
  {32'hbe9133e3, 32'h3e215578} /* (15, 26, 13) {real, imag} */,
  {32'hbf2d6aca, 32'hbdecd050} /* (15, 26, 12) {real, imag} */,
  {32'hbe05623b, 32'hbe96834e} /* (15, 26, 11) {real, imag} */,
  {32'h3deb982c, 32'hbe3f6acd} /* (15, 26, 10) {real, imag} */,
  {32'h3eb916e0, 32'h3e39addc} /* (15, 26, 9) {real, imag} */,
  {32'h3d2ab5d8, 32'h3ed2285a} /* (15, 26, 8) {real, imag} */,
  {32'hbf179a1a, 32'hbe32b79d} /* (15, 26, 7) {real, imag} */,
  {32'hbe92b338, 32'h3d64f512} /* (15, 26, 6) {real, imag} */,
  {32'hbf05bbba, 32'hbd97e1ae} /* (15, 26, 5) {real, imag} */,
  {32'hbe197bfb, 32'hbdfe0b64} /* (15, 26, 4) {real, imag} */,
  {32'hbe14832c, 32'hbb1fe200} /* (15, 26, 3) {real, imag} */,
  {32'hbe8c4c8c, 32'hbdaaa0e2} /* (15, 26, 2) {real, imag} */,
  {32'hbdae55e0, 32'hbe000aec} /* (15, 26, 1) {real, imag} */,
  {32'hbf4276ba, 32'h3e7f1662} /* (15, 26, 0) {real, imag} */,
  {32'hbef3f4ce, 32'hbfbbc676} /* (15, 25, 31) {real, imag} */,
  {32'h3d865af0, 32'h3e64b8f3} /* (15, 25, 30) {real, imag} */,
  {32'hbe38fe40, 32'h3f1afd12} /* (15, 25, 29) {real, imag} */,
  {32'h3e2a9560, 32'h3d8d7d96} /* (15, 25, 28) {real, imag} */,
  {32'hbe8381b0, 32'hbd036770} /* (15, 25, 27) {real, imag} */,
  {32'hbf376059, 32'hbd8575c0} /* (15, 25, 26) {real, imag} */,
  {32'h3ee723e0, 32'hbef2931c} /* (15, 25, 25) {real, imag} */,
  {32'h3dc734d8, 32'h3f43afac} /* (15, 25, 24) {real, imag} */,
  {32'hbee65b4a, 32'hbe1e1e08} /* (15, 25, 23) {real, imag} */,
  {32'hbe5579bb, 32'hbea2093c} /* (15, 25, 22) {real, imag} */,
  {32'h3e5cd702, 32'hbe6b1839} /* (15, 25, 21) {real, imag} */,
  {32'h3d5b1f98, 32'hbdda05a8} /* (15, 25, 20) {real, imag} */,
  {32'hbddf3f45, 32'h3e271ed0} /* (15, 25, 19) {real, imag} */,
  {32'h3e3721ee, 32'hbe619244} /* (15, 25, 18) {real, imag} */,
  {32'hbf24a7f4, 32'h3e7d1a4a} /* (15, 25, 17) {real, imag} */,
  {32'h3e338f60, 32'h3d95410c} /* (15, 25, 16) {real, imag} */,
  {32'h3dd3c8d6, 32'h3de792b3} /* (15, 25, 15) {real, imag} */,
  {32'hbe1891b0, 32'h3d8ecda0} /* (15, 25, 14) {real, imag} */,
  {32'h3d056e3c, 32'h3ea966a8} /* (15, 25, 13) {real, imag} */,
  {32'h3c77a16c, 32'h3e7d5cd6} /* (15, 25, 12) {real, imag} */,
  {32'hbd8b7bd2, 32'hbe83f200} /* (15, 25, 11) {real, imag} */,
  {32'h3d06d1ec, 32'hbd86a0d2} /* (15, 25, 10) {real, imag} */,
  {32'hbe9a118a, 32'hbd6632f0} /* (15, 25, 9) {real, imag} */,
  {32'hbe86301e, 32'hbd271cc0} /* (15, 25, 8) {real, imag} */,
  {32'hbd7dae48, 32'h3e99eca1} /* (15, 25, 7) {real, imag} */,
  {32'hbe512498, 32'h3d7655cf} /* (15, 25, 6) {real, imag} */,
  {32'hbd6d4d60, 32'h3e083c28} /* (15, 25, 5) {real, imag} */,
  {32'hbed74ada, 32'h3eb9a3a9} /* (15, 25, 4) {real, imag} */,
  {32'hbea15c1a, 32'h3d820f95} /* (15, 25, 3) {real, imag} */,
  {32'hbe24f2e0, 32'h3f52b5d8} /* (15, 25, 2) {real, imag} */,
  {32'h3e0f8f94, 32'hbf530667} /* (15, 25, 1) {real, imag} */,
  {32'hbe9173b2, 32'h3e33d8de} /* (15, 25, 0) {real, imag} */,
  {32'hbea135f8, 32'hbd203034} /* (15, 24, 31) {real, imag} */,
  {32'h3e5942dc, 32'hbeacadc0} /* (15, 24, 30) {real, imag} */,
  {32'hbea3cc91, 32'hbe432fc6} /* (15, 24, 29) {real, imag} */,
  {32'hbf1eede4, 32'h3e55b193} /* (15, 24, 28) {real, imag} */,
  {32'hbee1fe98, 32'hbc20e3d0} /* (15, 24, 27) {real, imag} */,
  {32'hbdd3ecc0, 32'h3f2d07a5} /* (15, 24, 26) {real, imag} */,
  {32'hbe3beffe, 32'h3e5624d1} /* (15, 24, 25) {real, imag} */,
  {32'h3f398e6d, 32'h3ea0452c} /* (15, 24, 24) {real, imag} */,
  {32'hbe40f554, 32'hbf317861} /* (15, 24, 23) {real, imag} */,
  {32'h3f0c8918, 32'hbe0277b6} /* (15, 24, 22) {real, imag} */,
  {32'h3e8946a8, 32'hbd7df039} /* (15, 24, 21) {real, imag} */,
  {32'hbf5b646c, 32'hbedcfacc} /* (15, 24, 20) {real, imag} */,
  {32'hbe28b95b, 32'hbe2ac47c} /* (15, 24, 19) {real, imag} */,
  {32'h3e45ee66, 32'h3c4625b0} /* (15, 24, 18) {real, imag} */,
  {32'hbcf32558, 32'hbcd0199c} /* (15, 24, 17) {real, imag} */,
  {32'h3df25459, 32'h3db2c0e6} /* (15, 24, 16) {real, imag} */,
  {32'h3b601b00, 32'h3f0f4e94} /* (15, 24, 15) {real, imag} */,
  {32'hbd7a0596, 32'hbe780001} /* (15, 24, 14) {real, imag} */,
  {32'hbeb127b6, 32'h3e8deb73} /* (15, 24, 13) {real, imag} */,
  {32'h3d69cbd0, 32'hbf4eaec4} /* (15, 24, 12) {real, imag} */,
  {32'h3eaf2227, 32'hbe09b929} /* (15, 24, 11) {real, imag} */,
  {32'h3f19e225, 32'hbd85f594} /* (15, 24, 10) {real, imag} */,
  {32'h3b568e60, 32'hbdda2ef9} /* (15, 24, 9) {real, imag} */,
  {32'h3ea266ed, 32'h3f29dcbd} /* (15, 24, 8) {real, imag} */,
  {32'hbea88eda, 32'h3f143f6a} /* (15, 24, 7) {real, imag} */,
  {32'h3edab47d, 32'hbefb1ad0} /* (15, 24, 6) {real, imag} */,
  {32'h3e3e9d01, 32'h3c1cc868} /* (15, 24, 5) {real, imag} */,
  {32'h3e94b431, 32'hbc6a31c8} /* (15, 24, 4) {real, imag} */,
  {32'h3ea6f42d, 32'hbd96e0b0} /* (15, 24, 3) {real, imag} */,
  {32'h3e864daf, 32'h3e5b79ee} /* (15, 24, 2) {real, imag} */,
  {32'hbfc29f92, 32'h3f66403c} /* (15, 24, 1) {real, imag} */,
  {32'hbede19bc, 32'hbef8a85e} /* (15, 24, 0) {real, imag} */,
  {32'h3e0861eb, 32'hbefa34c4} /* (15, 23, 31) {real, imag} */,
  {32'h3d63c11d, 32'h3e9d3a9a} /* (15, 23, 30) {real, imag} */,
  {32'h3e10f282, 32'hbd7b17ec} /* (15, 23, 29) {real, imag} */,
  {32'h3e033f1e, 32'hbe17cd32} /* (15, 23, 28) {real, imag} */,
  {32'hbebdd375, 32'h3d2f994c} /* (15, 23, 27) {real, imag} */,
  {32'h3ea2def8, 32'h3ce5c474} /* (15, 23, 26) {real, imag} */,
  {32'hbf0507d4, 32'hbeac7ce9} /* (15, 23, 25) {real, imag} */,
  {32'hbdc10ae4, 32'hbc33cff0} /* (15, 23, 24) {real, imag} */,
  {32'h3f73e339, 32'hbe7880e8} /* (15, 23, 23) {real, imag} */,
  {32'hbebfeab6, 32'h3ef933fa} /* (15, 23, 22) {real, imag} */,
  {32'hbe36edc6, 32'h3e4e0796} /* (15, 23, 21) {real, imag} */,
  {32'h3b0b9040, 32'h3e07c416} /* (15, 23, 20) {real, imag} */,
  {32'h3f0da9e6, 32'hbea1560c} /* (15, 23, 19) {real, imag} */,
  {32'hbec7de34, 32'hbd616fb8} /* (15, 23, 18) {real, imag} */,
  {32'h3db1e910, 32'h3e98f60c} /* (15, 23, 17) {real, imag} */,
  {32'h3d00c388, 32'hbe31c279} /* (15, 23, 16) {real, imag} */,
  {32'hbe48a230, 32'h3e9b818a} /* (15, 23, 15) {real, imag} */,
  {32'hbf2d5a77, 32'h3e8be229} /* (15, 23, 14) {real, imag} */,
  {32'h3ea232a6, 32'hbdd7059e} /* (15, 23, 13) {real, imag} */,
  {32'h3e1d0e71, 32'hbd0ff480} /* (15, 23, 12) {real, imag} */,
  {32'h3f049ac8, 32'hbea20442} /* (15, 23, 11) {real, imag} */,
  {32'hbe83ef04, 32'hbe8f584f} /* (15, 23, 10) {real, imag} */,
  {32'h3c37cfc8, 32'hbd2db888} /* (15, 23, 9) {real, imag} */,
  {32'h3de60bdc, 32'h3ee97ce5} /* (15, 23, 8) {real, imag} */,
  {32'h3eaa85e2, 32'h3e958ec2} /* (15, 23, 7) {real, imag} */,
  {32'h3ea614f0, 32'hbd9b0288} /* (15, 23, 6) {real, imag} */,
  {32'h3e8848ce, 32'h3ead4a82} /* (15, 23, 5) {real, imag} */,
  {32'hbdeb7816, 32'hbf5003c5} /* (15, 23, 4) {real, imag} */,
  {32'h3ec6c516, 32'h3cc4f5d0} /* (15, 23, 3) {real, imag} */,
  {32'h3c9ffb38, 32'h3dc05d1c} /* (15, 23, 2) {real, imag} */,
  {32'hbf4bdbc6, 32'h3d684b0c} /* (15, 23, 1) {real, imag} */,
  {32'h3ebcd3ad, 32'hbde6b44f} /* (15, 23, 0) {real, imag} */,
  {32'h3eabde19, 32'h3e9414fa} /* (15, 22, 31) {real, imag} */,
  {32'hbdba73da, 32'h3b8d84c0} /* (15, 22, 30) {real, imag} */,
  {32'h3e8a500b, 32'h3dfb16ae} /* (15, 22, 29) {real, imag} */,
  {32'hbe825d3b, 32'h3e3ca1ac} /* (15, 22, 28) {real, imag} */,
  {32'hbe70a26c, 32'h3ebd3b98} /* (15, 22, 27) {real, imag} */,
  {32'h3e88a96e, 32'hbe7d1cd7} /* (15, 22, 26) {real, imag} */,
  {32'h3e1cabba, 32'hbf0ba758} /* (15, 22, 25) {real, imag} */,
  {32'h3d5c6887, 32'hbeb171a3} /* (15, 22, 24) {real, imag} */,
  {32'h3e9f1e9a, 32'h3f164328} /* (15, 22, 23) {real, imag} */,
  {32'h3de602cf, 32'hbedc5e9a} /* (15, 22, 22) {real, imag} */,
  {32'hbdc45f7c, 32'hbf41c0e9} /* (15, 22, 21) {real, imag} */,
  {32'hbea3e690, 32'hbf141c16} /* (15, 22, 20) {real, imag} */,
  {32'h3f1e5785, 32'h3f2dbe84} /* (15, 22, 19) {real, imag} */,
  {32'h3ddcd0fb, 32'h3ef66fb0} /* (15, 22, 18) {real, imag} */,
  {32'hbf198c8e, 32'h3e5d692d} /* (15, 22, 17) {real, imag} */,
  {32'hbde8569a, 32'hbefc4d5c} /* (15, 22, 16) {real, imag} */,
  {32'hbd44aabc, 32'hbe2700cb} /* (15, 22, 15) {real, imag} */,
  {32'h3ce90b00, 32'hbe94e6cc} /* (15, 22, 14) {real, imag} */,
  {32'h3bb2f770, 32'h3f4bf15e} /* (15, 22, 13) {real, imag} */,
  {32'hbe835ca8, 32'h3eaebba8} /* (15, 22, 12) {real, imag} */,
  {32'hbe69f173, 32'h3f1c912c} /* (15, 22, 11) {real, imag} */,
  {32'h3e2338dd, 32'hbc2cda70} /* (15, 22, 10) {real, imag} */,
  {32'h3e2c5b3e, 32'h3db1c224} /* (15, 22, 9) {real, imag} */,
  {32'hbcf9b418, 32'hbe284e32} /* (15, 22, 8) {real, imag} */,
  {32'h3e2ee686, 32'hbe9b754f} /* (15, 22, 7) {real, imag} */,
  {32'hbf2baf52, 32'hbe4df8bc} /* (15, 22, 6) {real, imag} */,
  {32'h3dccde35, 32'hbe4b1294} /* (15, 22, 5) {real, imag} */,
  {32'hbe67dabf, 32'h3d8ce26c} /* (15, 22, 4) {real, imag} */,
  {32'h3d62c3ba, 32'h3e20a785} /* (15, 22, 3) {real, imag} */,
  {32'hbc435770, 32'h3f05b75f} /* (15, 22, 2) {real, imag} */,
  {32'h3e749bf6, 32'hbf5cd624} /* (15, 22, 1) {real, imag} */,
  {32'hbe43cad9, 32'hbf463b8a} /* (15, 22, 0) {real, imag} */,
  {32'hbda1a531, 32'h3edb11f4} /* (15, 21, 31) {real, imag} */,
  {32'hbe02e6dc, 32'h3d0c62d0} /* (15, 21, 30) {real, imag} */,
  {32'hbe9f5f3c, 32'h3f438fd4} /* (15, 21, 29) {real, imag} */,
  {32'hbf0eb5bc, 32'h3d7ad968} /* (15, 21, 28) {real, imag} */,
  {32'h3e3388e8, 32'hbec8e47d} /* (15, 21, 27) {real, imag} */,
  {32'hbe30b8c0, 32'h3e9f6d71} /* (15, 21, 26) {real, imag} */,
  {32'hbe9943d2, 32'h3d204028} /* (15, 21, 25) {real, imag} */,
  {32'hbe88699d, 32'hbeb2c9db} /* (15, 21, 24) {real, imag} */,
  {32'h3d37a4dc, 32'hbca1c018} /* (15, 21, 23) {real, imag} */,
  {32'h3eb21d83, 32'h3d0d9cb6} /* (15, 21, 22) {real, imag} */,
  {32'h3d395fd4, 32'h3e8c0ef5} /* (15, 21, 21) {real, imag} */,
  {32'hbe0184f5, 32'hbe8cf2aa} /* (15, 21, 20) {real, imag} */,
  {32'hbe8b3301, 32'hbe1979b1} /* (15, 21, 19) {real, imag} */,
  {32'h3dda1854, 32'h3c1d7444} /* (15, 21, 18) {real, imag} */,
  {32'h3e9577a3, 32'hbe244eec} /* (15, 21, 17) {real, imag} */,
  {32'hbdda2314, 32'hbe39968e} /* (15, 21, 16) {real, imag} */,
  {32'h3b87aae8, 32'hbeece434} /* (15, 21, 15) {real, imag} */,
  {32'h3f07fe86, 32'h3e67af1f} /* (15, 21, 14) {real, imag} */,
  {32'hbea7ee3e, 32'h3eda8a1c} /* (15, 21, 13) {real, imag} */,
  {32'hbdee7e66, 32'h3d3be098} /* (15, 21, 12) {real, imag} */,
  {32'h3c30a4a0, 32'hbf00f1b8} /* (15, 21, 11) {real, imag} */,
  {32'h3dbcbd70, 32'h3e096aba} /* (15, 21, 10) {real, imag} */,
  {32'h3d959004, 32'h3eac0643} /* (15, 21, 9) {real, imag} */,
  {32'h3f6039f2, 32'h3e704595} /* (15, 21, 8) {real, imag} */,
  {32'hbeac963e, 32'h3ee786d5} /* (15, 21, 7) {real, imag} */,
  {32'h3f6cd4a3, 32'h3cd82c9c} /* (15, 21, 6) {real, imag} */,
  {32'hbbeba950, 32'h3ed1fac0} /* (15, 21, 5) {real, imag} */,
  {32'hbeb02108, 32'hbe418964} /* (15, 21, 4) {real, imag} */,
  {32'h3d8d0332, 32'h3decf89c} /* (15, 21, 3) {real, imag} */,
  {32'hbe53ba79, 32'hbecf0f14} /* (15, 21, 2) {real, imag} */,
  {32'hbf4a16f4, 32'h3eae927c} /* (15, 21, 1) {real, imag} */,
  {32'hbe25f738, 32'h3e9b1666} /* (15, 21, 0) {real, imag} */,
  {32'h3d086f98, 32'hbed9220e} /* (15, 20, 31) {real, imag} */,
  {32'hbe8618a3, 32'h3e5ab32b} /* (15, 20, 30) {real, imag} */,
  {32'hbe9189f4, 32'h3f0f905a} /* (15, 20, 29) {real, imag} */,
  {32'hbe63f197, 32'h3e8f6d50} /* (15, 20, 28) {real, imag} */,
  {32'h3eb5a953, 32'h3e4e7f21} /* (15, 20, 27) {real, imag} */,
  {32'hbd8d799f, 32'hbea81c38} /* (15, 20, 26) {real, imag} */,
  {32'h3e6c6529, 32'hbdd2fa2d} /* (15, 20, 25) {real, imag} */,
  {32'h3e4b38d4, 32'h3e8b3488} /* (15, 20, 24) {real, imag} */,
  {32'hbeaa70f6, 32'hbea63754} /* (15, 20, 23) {real, imag} */,
  {32'hbea7e9e8, 32'hbecebe68} /* (15, 20, 22) {real, imag} */,
  {32'h3f201eba, 32'h3e9a93d3} /* (15, 20, 21) {real, imag} */,
  {32'h3dad81bf, 32'hbd2657d0} /* (15, 20, 20) {real, imag} */,
  {32'hbe7314ba, 32'h3cf681d0} /* (15, 20, 19) {real, imag} */,
  {32'hbdcf24b9, 32'hbeae4e73} /* (15, 20, 18) {real, imag} */,
  {32'h3eae5410, 32'h3dbaf877} /* (15, 20, 17) {real, imag} */,
  {32'h3e316a32, 32'h3dbd4aa8} /* (15, 20, 16) {real, imag} */,
  {32'h3eb449dc, 32'hbd0e7644} /* (15, 20, 15) {real, imag} */,
  {32'h3e07b404, 32'hbec7c534} /* (15, 20, 14) {real, imag} */,
  {32'h3e669179, 32'hbeb9619e} /* (15, 20, 13) {real, imag} */,
  {32'h3e9687ae, 32'hbdb5ca75} /* (15, 20, 12) {real, imag} */,
  {32'hbee318b4, 32'hbe637422} /* (15, 20, 11) {real, imag} */,
  {32'hbdd6d7dc, 32'h3e34075d} /* (15, 20, 10) {real, imag} */,
  {32'hbe39ad3b, 32'h3dfa429a} /* (15, 20, 9) {real, imag} */,
  {32'hbf07132c, 32'hbe26ce30} /* (15, 20, 8) {real, imag} */,
  {32'h3e9179e0, 32'hbe3e7a02} /* (15, 20, 7) {real, imag} */,
  {32'hbd940c78, 32'h3f206f24} /* (15, 20, 6) {real, imag} */,
  {32'h3e489ffa, 32'h3eadb6fe} /* (15, 20, 5) {real, imag} */,
  {32'h3da40939, 32'h3ea981e3} /* (15, 20, 4) {real, imag} */,
  {32'h3eaf42f4, 32'h3ef22d10} /* (15, 20, 3) {real, imag} */,
  {32'h3d4754a7, 32'hbe86c7c3} /* (15, 20, 2) {real, imag} */,
  {32'h3e5ed52e, 32'hbf13c004} /* (15, 20, 1) {real, imag} */,
  {32'hbe0fafb2, 32'hbcfb80ac} /* (15, 20, 0) {real, imag} */,
  {32'h3ec4528c, 32'h3e155aa4} /* (15, 19, 31) {real, imag} */,
  {32'h3db1b308, 32'hbd9e3a76} /* (15, 19, 30) {real, imag} */,
  {32'hbe40a7b6, 32'hbe24349a} /* (15, 19, 29) {real, imag} */,
  {32'hbcd318f8, 32'hbe40d10a} /* (15, 19, 28) {real, imag} */,
  {32'hbe643194, 32'hbbc2eae0} /* (15, 19, 27) {real, imag} */,
  {32'h3ee5323c, 32'h3e8ad525} /* (15, 19, 26) {real, imag} */,
  {32'hbe8b226f, 32'h3dc5673a} /* (15, 19, 25) {real, imag} */,
  {32'h3e4d01c0, 32'h3e15d680} /* (15, 19, 24) {real, imag} */,
  {32'hbea5cd7f, 32'h3f38d614} /* (15, 19, 23) {real, imag} */,
  {32'hbf2356d8, 32'hbd5235ba} /* (15, 19, 22) {real, imag} */,
  {32'hbdfec47e, 32'hbf0bcb15} /* (15, 19, 21) {real, imag} */,
  {32'hbeab972b, 32'h3e9f006b} /* (15, 19, 20) {real, imag} */,
  {32'hbdd8563a, 32'hbeba4796} /* (15, 19, 19) {real, imag} */,
  {32'h3ed24dfb, 32'hbe3b23a0} /* (15, 19, 18) {real, imag} */,
  {32'hbcfa7318, 32'hbe357bfd} /* (15, 19, 17) {real, imag} */,
  {32'h3de90f9c, 32'hbe5999f2} /* (15, 19, 16) {real, imag} */,
  {32'hbdcbcfd7, 32'hbd931e2a} /* (15, 19, 15) {real, imag} */,
  {32'hbea27eaa, 32'hbe1567e0} /* (15, 19, 14) {real, imag} */,
  {32'h3ddf08a4, 32'hbebe7b5a} /* (15, 19, 13) {real, imag} */,
  {32'h3d3465ac, 32'h3eeeab58} /* (15, 19, 12) {real, imag} */,
  {32'hbdf5d3b7, 32'h3ebd1e8f} /* (15, 19, 11) {real, imag} */,
  {32'hbe13b956, 32'hbe1a813b} /* (15, 19, 10) {real, imag} */,
  {32'h3e75b232, 32'h3ea8ca22} /* (15, 19, 9) {real, imag} */,
  {32'h3ef62936, 32'hbf01c546} /* (15, 19, 8) {real, imag} */,
  {32'hbe24ad6b, 32'h3e60c0e2} /* (15, 19, 7) {real, imag} */,
  {32'hbf00c296, 32'hbde61c9a} /* (15, 19, 6) {real, imag} */,
  {32'h3ea59ff4, 32'h3df03cdc} /* (15, 19, 5) {real, imag} */,
  {32'h3e8cc830, 32'hbc908a60} /* (15, 19, 4) {real, imag} */,
  {32'hbe00e214, 32'h3dbe024a} /* (15, 19, 3) {real, imag} */,
  {32'hbe4d178f, 32'hbdd89e20} /* (15, 19, 2) {real, imag} */,
  {32'h3e5d3e34, 32'hbdf4e2be} /* (15, 19, 1) {real, imag} */,
  {32'h3e42cfda, 32'hbe0ba94b} /* (15, 19, 0) {real, imag} */,
  {32'hbd83656a, 32'h3ecfaaf2} /* (15, 18, 31) {real, imag} */,
  {32'hbdb3ae70, 32'hbd2f0228} /* (15, 18, 30) {real, imag} */,
  {32'h3d553af8, 32'hbc549d80} /* (15, 18, 29) {real, imag} */,
  {32'h3ef7e942, 32'h3eaa45b4} /* (15, 18, 28) {real, imag} */,
  {32'hbe5b0aa2, 32'hbf31f232} /* (15, 18, 27) {real, imag} */,
  {32'h3d5a10ca, 32'hbe30575a} /* (15, 18, 26) {real, imag} */,
  {32'h3e96a9f6, 32'h3e935385} /* (15, 18, 25) {real, imag} */,
  {32'h3ecf6ace, 32'hbe15b549} /* (15, 18, 24) {real, imag} */,
  {32'hbd33c8a8, 32'hbce667c0} /* (15, 18, 23) {real, imag} */,
  {32'hbe87b5cd, 32'h3f27f712} /* (15, 18, 22) {real, imag} */,
  {32'h3dc3aa1e, 32'hbcd8423c} /* (15, 18, 21) {real, imag} */,
  {32'hba80b140, 32'h3dc471b8} /* (15, 18, 20) {real, imag} */,
  {32'hbeddd190, 32'h3e6f3170} /* (15, 18, 19) {real, imag} */,
  {32'h3d9d9f54, 32'h3d8f7c14} /* (15, 18, 18) {real, imag} */,
  {32'hbeb1bfd2, 32'h3ec12d76} /* (15, 18, 17) {real, imag} */,
  {32'hbe0acefc, 32'hbe1b3a0b} /* (15, 18, 16) {real, imag} */,
  {32'h3ebe4f8b, 32'h3d7c58d7} /* (15, 18, 15) {real, imag} */,
  {32'hbe26253c, 32'hbdc0c25a} /* (15, 18, 14) {real, imag} */,
  {32'h3e686bc9, 32'h3e68fd21} /* (15, 18, 13) {real, imag} */,
  {32'hbc4cd440, 32'hbdcb3b60} /* (15, 18, 12) {real, imag} */,
  {32'hbe26f1e6, 32'h3ed98f3c} /* (15, 18, 11) {real, imag} */,
  {32'h3db1f5cf, 32'h3e1b42ce} /* (15, 18, 10) {real, imag} */,
  {32'h3e8844a0, 32'hbe0f9ec6} /* (15, 18, 9) {real, imag} */,
  {32'hbda81da0, 32'hbe15893a} /* (15, 18, 8) {real, imag} */,
  {32'h3e7461e5, 32'hbe194466} /* (15, 18, 7) {real, imag} */,
  {32'h3f23e6bf, 32'h3eae205e} /* (15, 18, 6) {real, imag} */,
  {32'h3dd7fe4e, 32'h3e71a578} /* (15, 18, 5) {real, imag} */,
  {32'hbeaf7bae, 32'hbdb3095f} /* (15, 18, 4) {real, imag} */,
  {32'hbdd3b760, 32'hbe0d280e} /* (15, 18, 3) {real, imag} */,
  {32'h3e25dd2c, 32'hbe66d80c} /* (15, 18, 2) {real, imag} */,
  {32'hbe080169, 32'hbdb690b9} /* (15, 18, 1) {real, imag} */,
  {32'h3e28a740, 32'h3d1f55e4} /* (15, 18, 0) {real, imag} */,
  {32'hbda6252f, 32'h3d80d59b} /* (15, 17, 31) {real, imag} */,
  {32'h3ea52b5a, 32'h3e2d5fb1} /* (15, 17, 30) {real, imag} */,
  {32'hbeb1fade, 32'h3dc8657e} /* (15, 17, 29) {real, imag} */,
  {32'h3eb58e42, 32'hbeb11a27} /* (15, 17, 28) {real, imag} */,
  {32'hbe11406a, 32'h3e9507f7} /* (15, 17, 27) {real, imag} */,
  {32'hbe3a2af7, 32'hbe9aced4} /* (15, 17, 26) {real, imag} */,
  {32'h3ceef134, 32'h3ef5fd4e} /* (15, 17, 25) {real, imag} */,
  {32'h3eaad374, 32'h3d84b860} /* (15, 17, 24) {real, imag} */,
  {32'hbe507215, 32'h3e3bfc12} /* (15, 17, 23) {real, imag} */,
  {32'h3e89bea6, 32'hbe9060d2} /* (15, 17, 22) {real, imag} */,
  {32'h3e349f28, 32'hbec1f8df} /* (15, 17, 21) {real, imag} */,
  {32'h3e32e04a, 32'hbeb4f209} /* (15, 17, 20) {real, imag} */,
  {32'hbe9f98cf, 32'hbddf9378} /* (15, 17, 19) {real, imag} */,
  {32'h3edc3b28, 32'h3e0131de} /* (15, 17, 18) {real, imag} */,
  {32'h3d1441ba, 32'hbe8d8e0b} /* (15, 17, 17) {real, imag} */,
  {32'hbd82a65a, 32'h3e2c95c4} /* (15, 17, 16) {real, imag} */,
  {32'hbe799d2d, 32'hbe5d0174} /* (15, 17, 15) {real, imag} */,
  {32'hbe974deb, 32'hbf25ad7a} /* (15, 17, 14) {real, imag} */,
  {32'h3eab3ea4, 32'hbe83531c} /* (15, 17, 13) {real, imag} */,
  {32'h3e8fcba6, 32'hbd446a22} /* (15, 17, 12) {real, imag} */,
  {32'hbd71460c, 32'hbe18ff62} /* (15, 17, 11) {real, imag} */,
  {32'hbe9d3b2b, 32'h3ec94846} /* (15, 17, 10) {real, imag} */,
  {32'h3db7f27a, 32'hbd9c7d9e} /* (15, 17, 9) {real, imag} */,
  {32'hbefd3c97, 32'h3efd9056} /* (15, 17, 8) {real, imag} */,
  {32'hbe8466fe, 32'hbd2be760} /* (15, 17, 7) {real, imag} */,
  {32'hbdb43282, 32'hbedb0ea9} /* (15, 17, 6) {real, imag} */,
  {32'hbe8d420a, 32'hbec23128} /* (15, 17, 5) {real, imag} */,
  {32'h3f106119, 32'h3e03ec6c} /* (15, 17, 4) {real, imag} */,
  {32'hbe213ff2, 32'hbdbe2f7a} /* (15, 17, 3) {real, imag} */,
  {32'hbc928ba8, 32'h3ee68018} /* (15, 17, 2) {real, imag} */,
  {32'hbddc69da, 32'h3e05c3aa} /* (15, 17, 1) {real, imag} */,
  {32'h3deaf4fc, 32'hbd41a4ce} /* (15, 17, 0) {real, imag} */,
  {32'hbe83b388, 32'h3e5a5796} /* (15, 16, 31) {real, imag} */,
  {32'h3df05b42, 32'h3cae0c0e} /* (15, 16, 30) {real, imag} */,
  {32'h3e71de90, 32'h3e80c47c} /* (15, 16, 29) {real, imag} */,
  {32'h3d72695a, 32'h3e6b6686} /* (15, 16, 28) {real, imag} */,
  {32'hbdbe4145, 32'h3e06af9e} /* (15, 16, 27) {real, imag} */,
  {32'h3d91fb45, 32'h3c4db650} /* (15, 16, 26) {real, imag} */,
  {32'h3c9c9398, 32'h3bbd38fc} /* (15, 16, 25) {real, imag} */,
  {32'hbd95c203, 32'hbdbf1795} /* (15, 16, 24) {real, imag} */,
  {32'hbe6af1f2, 32'hbd772e90} /* (15, 16, 23) {real, imag} */,
  {32'h3e221f8d, 32'hbd18d14a} /* (15, 16, 22) {real, imag} */,
  {32'h3e875eb5, 32'h3dda4cce} /* (15, 16, 21) {real, imag} */,
  {32'hbdce479a, 32'hbe6e0dd7} /* (15, 16, 20) {real, imag} */,
  {32'h3f0a2272, 32'h3e0c061a} /* (15, 16, 19) {real, imag} */,
  {32'hbe05e722, 32'h3e378ef1} /* (15, 16, 18) {real, imag} */,
  {32'h3e779cfc, 32'hbeb83e36} /* (15, 16, 17) {real, imag} */,
  {32'h3ef81d5d, 32'h00000000} /* (15, 16, 16) {real, imag} */,
  {32'h3e779cfc, 32'h3eb83e36} /* (15, 16, 15) {real, imag} */,
  {32'hbe05e722, 32'hbe378ef1} /* (15, 16, 14) {real, imag} */,
  {32'h3f0a2272, 32'hbe0c061a} /* (15, 16, 13) {real, imag} */,
  {32'hbdce479a, 32'h3e6e0dd7} /* (15, 16, 12) {real, imag} */,
  {32'h3e875eb5, 32'hbdda4cce} /* (15, 16, 11) {real, imag} */,
  {32'h3e221f8d, 32'h3d18d14a} /* (15, 16, 10) {real, imag} */,
  {32'hbe6af1f2, 32'h3d772e90} /* (15, 16, 9) {real, imag} */,
  {32'hbd95c203, 32'h3dbf1795} /* (15, 16, 8) {real, imag} */,
  {32'h3c9c9398, 32'hbbbd38fc} /* (15, 16, 7) {real, imag} */,
  {32'h3d91fb45, 32'hbc4db650} /* (15, 16, 6) {real, imag} */,
  {32'hbdbe4145, 32'hbe06af9e} /* (15, 16, 5) {real, imag} */,
  {32'h3d72695a, 32'hbe6b6686} /* (15, 16, 4) {real, imag} */,
  {32'h3e71de90, 32'hbe80c47c} /* (15, 16, 3) {real, imag} */,
  {32'h3df05b42, 32'hbcae0c0e} /* (15, 16, 2) {real, imag} */,
  {32'hbe83b388, 32'hbe5a5796} /* (15, 16, 1) {real, imag} */,
  {32'h3daf705b, 32'h00000000} /* (15, 16, 0) {real, imag} */,
  {32'hbddc69da, 32'hbe05c3aa} /* (15, 15, 31) {real, imag} */,
  {32'hbc928ba8, 32'hbee68018} /* (15, 15, 30) {real, imag} */,
  {32'hbe213ff2, 32'h3dbe2f7a} /* (15, 15, 29) {real, imag} */,
  {32'h3f106119, 32'hbe03ec6c} /* (15, 15, 28) {real, imag} */,
  {32'hbe8d420a, 32'h3ec23128} /* (15, 15, 27) {real, imag} */,
  {32'hbdb43282, 32'h3edb0ea9} /* (15, 15, 26) {real, imag} */,
  {32'hbe8466fe, 32'h3d2be760} /* (15, 15, 25) {real, imag} */,
  {32'hbefd3c97, 32'hbefd9056} /* (15, 15, 24) {real, imag} */,
  {32'h3db7f27a, 32'h3d9c7d9e} /* (15, 15, 23) {real, imag} */,
  {32'hbe9d3b2b, 32'hbec94846} /* (15, 15, 22) {real, imag} */,
  {32'hbd71460c, 32'h3e18ff62} /* (15, 15, 21) {real, imag} */,
  {32'h3e8fcba6, 32'h3d446a22} /* (15, 15, 20) {real, imag} */,
  {32'h3eab3ea4, 32'h3e83531c} /* (15, 15, 19) {real, imag} */,
  {32'hbe974deb, 32'h3f25ad7a} /* (15, 15, 18) {real, imag} */,
  {32'hbe799d2d, 32'h3e5d0174} /* (15, 15, 17) {real, imag} */,
  {32'hbd82a65a, 32'hbe2c95c4} /* (15, 15, 16) {real, imag} */,
  {32'h3d1441ba, 32'h3e8d8e0b} /* (15, 15, 15) {real, imag} */,
  {32'h3edc3b28, 32'hbe0131de} /* (15, 15, 14) {real, imag} */,
  {32'hbe9f98cf, 32'h3ddf9378} /* (15, 15, 13) {real, imag} */,
  {32'h3e32e04a, 32'h3eb4f209} /* (15, 15, 12) {real, imag} */,
  {32'h3e349f28, 32'h3ec1f8df} /* (15, 15, 11) {real, imag} */,
  {32'h3e89bea6, 32'h3e9060d2} /* (15, 15, 10) {real, imag} */,
  {32'hbe507215, 32'hbe3bfc12} /* (15, 15, 9) {real, imag} */,
  {32'h3eaad374, 32'hbd84b860} /* (15, 15, 8) {real, imag} */,
  {32'h3ceef134, 32'hbef5fd4e} /* (15, 15, 7) {real, imag} */,
  {32'hbe3a2af7, 32'h3e9aced4} /* (15, 15, 6) {real, imag} */,
  {32'hbe11406a, 32'hbe9507f7} /* (15, 15, 5) {real, imag} */,
  {32'h3eb58e42, 32'h3eb11a27} /* (15, 15, 4) {real, imag} */,
  {32'hbeb1fade, 32'hbdc8657e} /* (15, 15, 3) {real, imag} */,
  {32'h3ea52b5a, 32'hbe2d5fb1} /* (15, 15, 2) {real, imag} */,
  {32'hbda6252f, 32'hbd80d59b} /* (15, 15, 1) {real, imag} */,
  {32'h3deaf4fc, 32'h3d41a4ce} /* (15, 15, 0) {real, imag} */,
  {32'hbe080169, 32'h3db690b9} /* (15, 14, 31) {real, imag} */,
  {32'h3e25dd2c, 32'h3e66d80c} /* (15, 14, 30) {real, imag} */,
  {32'hbdd3b760, 32'h3e0d280e} /* (15, 14, 29) {real, imag} */,
  {32'hbeaf7bae, 32'h3db3095f} /* (15, 14, 28) {real, imag} */,
  {32'h3dd7fe4e, 32'hbe71a578} /* (15, 14, 27) {real, imag} */,
  {32'h3f23e6bf, 32'hbeae205e} /* (15, 14, 26) {real, imag} */,
  {32'h3e7461e5, 32'h3e194466} /* (15, 14, 25) {real, imag} */,
  {32'hbda81da0, 32'h3e15893a} /* (15, 14, 24) {real, imag} */,
  {32'h3e8844a0, 32'h3e0f9ec6} /* (15, 14, 23) {real, imag} */,
  {32'h3db1f5cf, 32'hbe1b42ce} /* (15, 14, 22) {real, imag} */,
  {32'hbe26f1e6, 32'hbed98f3c} /* (15, 14, 21) {real, imag} */,
  {32'hbc4cd440, 32'h3dcb3b60} /* (15, 14, 20) {real, imag} */,
  {32'h3e686bc9, 32'hbe68fd21} /* (15, 14, 19) {real, imag} */,
  {32'hbe26253c, 32'h3dc0c25a} /* (15, 14, 18) {real, imag} */,
  {32'h3ebe4f8b, 32'hbd7c58d7} /* (15, 14, 17) {real, imag} */,
  {32'hbe0acefc, 32'h3e1b3a0b} /* (15, 14, 16) {real, imag} */,
  {32'hbeb1bfd2, 32'hbec12d76} /* (15, 14, 15) {real, imag} */,
  {32'h3d9d9f54, 32'hbd8f7c14} /* (15, 14, 14) {real, imag} */,
  {32'hbeddd190, 32'hbe6f3170} /* (15, 14, 13) {real, imag} */,
  {32'hba80b140, 32'hbdc471b8} /* (15, 14, 12) {real, imag} */,
  {32'h3dc3aa1e, 32'h3cd8423c} /* (15, 14, 11) {real, imag} */,
  {32'hbe87b5cd, 32'hbf27f712} /* (15, 14, 10) {real, imag} */,
  {32'hbd33c8a8, 32'h3ce667c0} /* (15, 14, 9) {real, imag} */,
  {32'h3ecf6ace, 32'h3e15b549} /* (15, 14, 8) {real, imag} */,
  {32'h3e96a9f6, 32'hbe935385} /* (15, 14, 7) {real, imag} */,
  {32'h3d5a10ca, 32'h3e30575a} /* (15, 14, 6) {real, imag} */,
  {32'hbe5b0aa2, 32'h3f31f232} /* (15, 14, 5) {real, imag} */,
  {32'h3ef7e942, 32'hbeaa45b4} /* (15, 14, 4) {real, imag} */,
  {32'h3d553af8, 32'h3c549d80} /* (15, 14, 3) {real, imag} */,
  {32'hbdb3ae70, 32'h3d2f0228} /* (15, 14, 2) {real, imag} */,
  {32'hbd83656a, 32'hbecfaaf2} /* (15, 14, 1) {real, imag} */,
  {32'h3e28a740, 32'hbd1f55e4} /* (15, 14, 0) {real, imag} */,
  {32'h3e5d3e34, 32'h3df4e2be} /* (15, 13, 31) {real, imag} */,
  {32'hbe4d178f, 32'h3dd89e20} /* (15, 13, 30) {real, imag} */,
  {32'hbe00e214, 32'hbdbe024a} /* (15, 13, 29) {real, imag} */,
  {32'h3e8cc830, 32'h3c908a60} /* (15, 13, 28) {real, imag} */,
  {32'h3ea59ff4, 32'hbdf03cdc} /* (15, 13, 27) {real, imag} */,
  {32'hbf00c296, 32'h3de61c9a} /* (15, 13, 26) {real, imag} */,
  {32'hbe24ad6b, 32'hbe60c0e2} /* (15, 13, 25) {real, imag} */,
  {32'h3ef62936, 32'h3f01c546} /* (15, 13, 24) {real, imag} */,
  {32'h3e75b232, 32'hbea8ca22} /* (15, 13, 23) {real, imag} */,
  {32'hbe13b956, 32'h3e1a813b} /* (15, 13, 22) {real, imag} */,
  {32'hbdf5d3b7, 32'hbebd1e8f} /* (15, 13, 21) {real, imag} */,
  {32'h3d3465ac, 32'hbeeeab58} /* (15, 13, 20) {real, imag} */,
  {32'h3ddf08a4, 32'h3ebe7b5a} /* (15, 13, 19) {real, imag} */,
  {32'hbea27eaa, 32'h3e1567e0} /* (15, 13, 18) {real, imag} */,
  {32'hbdcbcfd7, 32'h3d931e2a} /* (15, 13, 17) {real, imag} */,
  {32'h3de90f9c, 32'h3e5999f2} /* (15, 13, 16) {real, imag} */,
  {32'hbcfa7318, 32'h3e357bfd} /* (15, 13, 15) {real, imag} */,
  {32'h3ed24dfb, 32'h3e3b23a0} /* (15, 13, 14) {real, imag} */,
  {32'hbdd8563a, 32'h3eba4796} /* (15, 13, 13) {real, imag} */,
  {32'hbeab972b, 32'hbe9f006b} /* (15, 13, 12) {real, imag} */,
  {32'hbdfec47e, 32'h3f0bcb15} /* (15, 13, 11) {real, imag} */,
  {32'hbf2356d8, 32'h3d5235ba} /* (15, 13, 10) {real, imag} */,
  {32'hbea5cd7f, 32'hbf38d614} /* (15, 13, 9) {real, imag} */,
  {32'h3e4d01c0, 32'hbe15d680} /* (15, 13, 8) {real, imag} */,
  {32'hbe8b226f, 32'hbdc5673a} /* (15, 13, 7) {real, imag} */,
  {32'h3ee5323c, 32'hbe8ad525} /* (15, 13, 6) {real, imag} */,
  {32'hbe643194, 32'h3bc2eae0} /* (15, 13, 5) {real, imag} */,
  {32'hbcd318f8, 32'h3e40d10a} /* (15, 13, 4) {real, imag} */,
  {32'hbe40a7b6, 32'h3e24349a} /* (15, 13, 3) {real, imag} */,
  {32'h3db1b308, 32'h3d9e3a76} /* (15, 13, 2) {real, imag} */,
  {32'h3ec4528c, 32'hbe155aa4} /* (15, 13, 1) {real, imag} */,
  {32'h3e42cfda, 32'h3e0ba94b} /* (15, 13, 0) {real, imag} */,
  {32'h3e5ed52e, 32'h3f13c004} /* (15, 12, 31) {real, imag} */,
  {32'h3d4754a7, 32'h3e86c7c3} /* (15, 12, 30) {real, imag} */,
  {32'h3eaf42f4, 32'hbef22d10} /* (15, 12, 29) {real, imag} */,
  {32'h3da40939, 32'hbea981e3} /* (15, 12, 28) {real, imag} */,
  {32'h3e489ffa, 32'hbeadb6fe} /* (15, 12, 27) {real, imag} */,
  {32'hbd940c78, 32'hbf206f24} /* (15, 12, 26) {real, imag} */,
  {32'h3e9179e0, 32'h3e3e7a02} /* (15, 12, 25) {real, imag} */,
  {32'hbf07132c, 32'h3e26ce30} /* (15, 12, 24) {real, imag} */,
  {32'hbe39ad3b, 32'hbdfa429a} /* (15, 12, 23) {real, imag} */,
  {32'hbdd6d7dc, 32'hbe34075d} /* (15, 12, 22) {real, imag} */,
  {32'hbee318b4, 32'h3e637422} /* (15, 12, 21) {real, imag} */,
  {32'h3e9687ae, 32'h3db5ca75} /* (15, 12, 20) {real, imag} */,
  {32'h3e669179, 32'h3eb9619e} /* (15, 12, 19) {real, imag} */,
  {32'h3e07b404, 32'h3ec7c534} /* (15, 12, 18) {real, imag} */,
  {32'h3eb449dc, 32'h3d0e7644} /* (15, 12, 17) {real, imag} */,
  {32'h3e316a32, 32'hbdbd4aa8} /* (15, 12, 16) {real, imag} */,
  {32'h3eae5410, 32'hbdbaf877} /* (15, 12, 15) {real, imag} */,
  {32'hbdcf24b9, 32'h3eae4e73} /* (15, 12, 14) {real, imag} */,
  {32'hbe7314ba, 32'hbcf681d0} /* (15, 12, 13) {real, imag} */,
  {32'h3dad81bf, 32'h3d2657d0} /* (15, 12, 12) {real, imag} */,
  {32'h3f201eba, 32'hbe9a93d3} /* (15, 12, 11) {real, imag} */,
  {32'hbea7e9e8, 32'h3ecebe68} /* (15, 12, 10) {real, imag} */,
  {32'hbeaa70f6, 32'h3ea63754} /* (15, 12, 9) {real, imag} */,
  {32'h3e4b38d4, 32'hbe8b3488} /* (15, 12, 8) {real, imag} */,
  {32'h3e6c6529, 32'h3dd2fa2d} /* (15, 12, 7) {real, imag} */,
  {32'hbd8d799f, 32'h3ea81c38} /* (15, 12, 6) {real, imag} */,
  {32'h3eb5a953, 32'hbe4e7f21} /* (15, 12, 5) {real, imag} */,
  {32'hbe63f197, 32'hbe8f6d50} /* (15, 12, 4) {real, imag} */,
  {32'hbe9189f4, 32'hbf0f905a} /* (15, 12, 3) {real, imag} */,
  {32'hbe8618a3, 32'hbe5ab32b} /* (15, 12, 2) {real, imag} */,
  {32'h3d086f98, 32'h3ed9220e} /* (15, 12, 1) {real, imag} */,
  {32'hbe0fafb2, 32'h3cfb80ac} /* (15, 12, 0) {real, imag} */,
  {32'hbf4a16f4, 32'hbeae927c} /* (15, 11, 31) {real, imag} */,
  {32'hbe53ba79, 32'h3ecf0f14} /* (15, 11, 30) {real, imag} */,
  {32'h3d8d0332, 32'hbdecf89c} /* (15, 11, 29) {real, imag} */,
  {32'hbeb02108, 32'h3e418964} /* (15, 11, 28) {real, imag} */,
  {32'hbbeba950, 32'hbed1fac0} /* (15, 11, 27) {real, imag} */,
  {32'h3f6cd4a3, 32'hbcd82c9c} /* (15, 11, 26) {real, imag} */,
  {32'hbeac963e, 32'hbee786d5} /* (15, 11, 25) {real, imag} */,
  {32'h3f6039f2, 32'hbe704595} /* (15, 11, 24) {real, imag} */,
  {32'h3d959004, 32'hbeac0643} /* (15, 11, 23) {real, imag} */,
  {32'h3dbcbd70, 32'hbe096aba} /* (15, 11, 22) {real, imag} */,
  {32'h3c30a4a0, 32'h3f00f1b8} /* (15, 11, 21) {real, imag} */,
  {32'hbdee7e66, 32'hbd3be098} /* (15, 11, 20) {real, imag} */,
  {32'hbea7ee3e, 32'hbeda8a1c} /* (15, 11, 19) {real, imag} */,
  {32'h3f07fe86, 32'hbe67af1f} /* (15, 11, 18) {real, imag} */,
  {32'h3b87aae8, 32'h3eece434} /* (15, 11, 17) {real, imag} */,
  {32'hbdda2314, 32'h3e39968e} /* (15, 11, 16) {real, imag} */,
  {32'h3e9577a3, 32'h3e244eec} /* (15, 11, 15) {real, imag} */,
  {32'h3dda1854, 32'hbc1d7444} /* (15, 11, 14) {real, imag} */,
  {32'hbe8b3301, 32'h3e1979b1} /* (15, 11, 13) {real, imag} */,
  {32'hbe0184f5, 32'h3e8cf2aa} /* (15, 11, 12) {real, imag} */,
  {32'h3d395fd4, 32'hbe8c0ef5} /* (15, 11, 11) {real, imag} */,
  {32'h3eb21d83, 32'hbd0d9cb6} /* (15, 11, 10) {real, imag} */,
  {32'h3d37a4dc, 32'h3ca1c018} /* (15, 11, 9) {real, imag} */,
  {32'hbe88699d, 32'h3eb2c9db} /* (15, 11, 8) {real, imag} */,
  {32'hbe9943d2, 32'hbd204028} /* (15, 11, 7) {real, imag} */,
  {32'hbe30b8c0, 32'hbe9f6d71} /* (15, 11, 6) {real, imag} */,
  {32'h3e3388e8, 32'h3ec8e47d} /* (15, 11, 5) {real, imag} */,
  {32'hbf0eb5bc, 32'hbd7ad968} /* (15, 11, 4) {real, imag} */,
  {32'hbe9f5f3c, 32'hbf438fd4} /* (15, 11, 3) {real, imag} */,
  {32'hbe02e6dc, 32'hbd0c62d0} /* (15, 11, 2) {real, imag} */,
  {32'hbda1a531, 32'hbedb11f4} /* (15, 11, 1) {real, imag} */,
  {32'hbe25f738, 32'hbe9b1666} /* (15, 11, 0) {real, imag} */,
  {32'h3e749bf6, 32'h3f5cd624} /* (15, 10, 31) {real, imag} */,
  {32'hbc435770, 32'hbf05b75f} /* (15, 10, 30) {real, imag} */,
  {32'h3d62c3ba, 32'hbe20a785} /* (15, 10, 29) {real, imag} */,
  {32'hbe67dabf, 32'hbd8ce26c} /* (15, 10, 28) {real, imag} */,
  {32'h3dccde35, 32'h3e4b1294} /* (15, 10, 27) {real, imag} */,
  {32'hbf2baf52, 32'h3e4df8bc} /* (15, 10, 26) {real, imag} */,
  {32'h3e2ee686, 32'h3e9b754f} /* (15, 10, 25) {real, imag} */,
  {32'hbcf9b418, 32'h3e284e32} /* (15, 10, 24) {real, imag} */,
  {32'h3e2c5b3e, 32'hbdb1c224} /* (15, 10, 23) {real, imag} */,
  {32'h3e2338dd, 32'h3c2cda70} /* (15, 10, 22) {real, imag} */,
  {32'hbe69f173, 32'hbf1c912c} /* (15, 10, 21) {real, imag} */,
  {32'hbe835ca8, 32'hbeaebba8} /* (15, 10, 20) {real, imag} */,
  {32'h3bb2f770, 32'hbf4bf15e} /* (15, 10, 19) {real, imag} */,
  {32'h3ce90b00, 32'h3e94e6cc} /* (15, 10, 18) {real, imag} */,
  {32'hbd44aabc, 32'h3e2700cb} /* (15, 10, 17) {real, imag} */,
  {32'hbde8569a, 32'h3efc4d5c} /* (15, 10, 16) {real, imag} */,
  {32'hbf198c8e, 32'hbe5d692d} /* (15, 10, 15) {real, imag} */,
  {32'h3ddcd0fb, 32'hbef66fb0} /* (15, 10, 14) {real, imag} */,
  {32'h3f1e5785, 32'hbf2dbe84} /* (15, 10, 13) {real, imag} */,
  {32'hbea3e690, 32'h3f141c16} /* (15, 10, 12) {real, imag} */,
  {32'hbdc45f7c, 32'h3f41c0e9} /* (15, 10, 11) {real, imag} */,
  {32'h3de602cf, 32'h3edc5e9a} /* (15, 10, 10) {real, imag} */,
  {32'h3e9f1e9a, 32'hbf164328} /* (15, 10, 9) {real, imag} */,
  {32'h3d5c6887, 32'h3eb171a3} /* (15, 10, 8) {real, imag} */,
  {32'h3e1cabba, 32'h3f0ba758} /* (15, 10, 7) {real, imag} */,
  {32'h3e88a96e, 32'h3e7d1cd7} /* (15, 10, 6) {real, imag} */,
  {32'hbe70a26c, 32'hbebd3b98} /* (15, 10, 5) {real, imag} */,
  {32'hbe825d3b, 32'hbe3ca1ac} /* (15, 10, 4) {real, imag} */,
  {32'h3e8a500b, 32'hbdfb16ae} /* (15, 10, 3) {real, imag} */,
  {32'hbdba73da, 32'hbb8d84c0} /* (15, 10, 2) {real, imag} */,
  {32'h3eabde19, 32'hbe9414fa} /* (15, 10, 1) {real, imag} */,
  {32'hbe43cad9, 32'h3f463b8a} /* (15, 10, 0) {real, imag} */,
  {32'hbf4bdbc6, 32'hbd684b0c} /* (15, 9, 31) {real, imag} */,
  {32'h3c9ffb38, 32'hbdc05d1c} /* (15, 9, 30) {real, imag} */,
  {32'h3ec6c516, 32'hbcc4f5d0} /* (15, 9, 29) {real, imag} */,
  {32'hbdeb7816, 32'h3f5003c5} /* (15, 9, 28) {real, imag} */,
  {32'h3e8848ce, 32'hbead4a82} /* (15, 9, 27) {real, imag} */,
  {32'h3ea614f0, 32'h3d9b0288} /* (15, 9, 26) {real, imag} */,
  {32'h3eaa85e2, 32'hbe958ec2} /* (15, 9, 25) {real, imag} */,
  {32'h3de60bdc, 32'hbee97ce5} /* (15, 9, 24) {real, imag} */,
  {32'h3c37cfc8, 32'h3d2db888} /* (15, 9, 23) {real, imag} */,
  {32'hbe83ef04, 32'h3e8f584f} /* (15, 9, 22) {real, imag} */,
  {32'h3f049ac8, 32'h3ea20442} /* (15, 9, 21) {real, imag} */,
  {32'h3e1d0e71, 32'h3d0ff480} /* (15, 9, 20) {real, imag} */,
  {32'h3ea232a6, 32'h3dd7059e} /* (15, 9, 19) {real, imag} */,
  {32'hbf2d5a77, 32'hbe8be229} /* (15, 9, 18) {real, imag} */,
  {32'hbe48a230, 32'hbe9b818a} /* (15, 9, 17) {real, imag} */,
  {32'h3d00c388, 32'h3e31c279} /* (15, 9, 16) {real, imag} */,
  {32'h3db1e910, 32'hbe98f60c} /* (15, 9, 15) {real, imag} */,
  {32'hbec7de34, 32'h3d616fb8} /* (15, 9, 14) {real, imag} */,
  {32'h3f0da9e6, 32'h3ea1560c} /* (15, 9, 13) {real, imag} */,
  {32'h3b0b9040, 32'hbe07c416} /* (15, 9, 12) {real, imag} */,
  {32'hbe36edc6, 32'hbe4e0796} /* (15, 9, 11) {real, imag} */,
  {32'hbebfeab6, 32'hbef933fa} /* (15, 9, 10) {real, imag} */,
  {32'h3f73e339, 32'h3e7880e8} /* (15, 9, 9) {real, imag} */,
  {32'hbdc10ae4, 32'h3c33cff0} /* (15, 9, 8) {real, imag} */,
  {32'hbf0507d4, 32'h3eac7ce9} /* (15, 9, 7) {real, imag} */,
  {32'h3ea2def8, 32'hbce5c474} /* (15, 9, 6) {real, imag} */,
  {32'hbebdd375, 32'hbd2f994c} /* (15, 9, 5) {real, imag} */,
  {32'h3e033f1e, 32'h3e17cd32} /* (15, 9, 4) {real, imag} */,
  {32'h3e10f282, 32'h3d7b17ec} /* (15, 9, 3) {real, imag} */,
  {32'h3d63c11d, 32'hbe9d3a9a} /* (15, 9, 2) {real, imag} */,
  {32'h3e0861eb, 32'h3efa34c4} /* (15, 9, 1) {real, imag} */,
  {32'h3ebcd3ad, 32'h3de6b44f} /* (15, 9, 0) {real, imag} */,
  {32'hbfc29f92, 32'hbf66403c} /* (15, 8, 31) {real, imag} */,
  {32'h3e864daf, 32'hbe5b79ee} /* (15, 8, 30) {real, imag} */,
  {32'h3ea6f42d, 32'h3d96e0b0} /* (15, 8, 29) {real, imag} */,
  {32'h3e94b431, 32'h3c6a31c8} /* (15, 8, 28) {real, imag} */,
  {32'h3e3e9d01, 32'hbc1cc868} /* (15, 8, 27) {real, imag} */,
  {32'h3edab47d, 32'h3efb1ad0} /* (15, 8, 26) {real, imag} */,
  {32'hbea88eda, 32'hbf143f6a} /* (15, 8, 25) {real, imag} */,
  {32'h3ea266ed, 32'hbf29dcbd} /* (15, 8, 24) {real, imag} */,
  {32'h3b568e60, 32'h3dda2ef9} /* (15, 8, 23) {real, imag} */,
  {32'h3f19e225, 32'h3d85f594} /* (15, 8, 22) {real, imag} */,
  {32'h3eaf2227, 32'h3e09b929} /* (15, 8, 21) {real, imag} */,
  {32'h3d69cbd0, 32'h3f4eaec4} /* (15, 8, 20) {real, imag} */,
  {32'hbeb127b6, 32'hbe8deb73} /* (15, 8, 19) {real, imag} */,
  {32'hbd7a0596, 32'h3e780001} /* (15, 8, 18) {real, imag} */,
  {32'h3b601b00, 32'hbf0f4e94} /* (15, 8, 17) {real, imag} */,
  {32'h3df25459, 32'hbdb2c0e6} /* (15, 8, 16) {real, imag} */,
  {32'hbcf32558, 32'h3cd0199c} /* (15, 8, 15) {real, imag} */,
  {32'h3e45ee66, 32'hbc4625b0} /* (15, 8, 14) {real, imag} */,
  {32'hbe28b95b, 32'h3e2ac47c} /* (15, 8, 13) {real, imag} */,
  {32'hbf5b646c, 32'h3edcfacc} /* (15, 8, 12) {real, imag} */,
  {32'h3e8946a8, 32'h3d7df039} /* (15, 8, 11) {real, imag} */,
  {32'h3f0c8918, 32'h3e0277b6} /* (15, 8, 10) {real, imag} */,
  {32'hbe40f554, 32'h3f317861} /* (15, 8, 9) {real, imag} */,
  {32'h3f398e6d, 32'hbea0452c} /* (15, 8, 8) {real, imag} */,
  {32'hbe3beffe, 32'hbe5624d1} /* (15, 8, 7) {real, imag} */,
  {32'hbdd3ecc0, 32'hbf2d07a5} /* (15, 8, 6) {real, imag} */,
  {32'hbee1fe98, 32'h3c20e3d0} /* (15, 8, 5) {real, imag} */,
  {32'hbf1eede4, 32'hbe55b193} /* (15, 8, 4) {real, imag} */,
  {32'hbea3cc91, 32'h3e432fc6} /* (15, 8, 3) {real, imag} */,
  {32'h3e5942dc, 32'h3eacadc0} /* (15, 8, 2) {real, imag} */,
  {32'hbea135f8, 32'h3d203034} /* (15, 8, 1) {real, imag} */,
  {32'hbede19bc, 32'h3ef8a85e} /* (15, 8, 0) {real, imag} */,
  {32'h3e0f8f94, 32'h3f530667} /* (15, 7, 31) {real, imag} */,
  {32'hbe24f2e0, 32'hbf52b5d8} /* (15, 7, 30) {real, imag} */,
  {32'hbea15c1a, 32'hbd820f95} /* (15, 7, 29) {real, imag} */,
  {32'hbed74ada, 32'hbeb9a3a9} /* (15, 7, 28) {real, imag} */,
  {32'hbd6d4d60, 32'hbe083c28} /* (15, 7, 27) {real, imag} */,
  {32'hbe512498, 32'hbd7655cf} /* (15, 7, 26) {real, imag} */,
  {32'hbd7dae48, 32'hbe99eca1} /* (15, 7, 25) {real, imag} */,
  {32'hbe86301e, 32'h3d271cc0} /* (15, 7, 24) {real, imag} */,
  {32'hbe9a118a, 32'h3d6632f0} /* (15, 7, 23) {real, imag} */,
  {32'h3d06d1ec, 32'h3d86a0d2} /* (15, 7, 22) {real, imag} */,
  {32'hbd8b7bd2, 32'h3e83f200} /* (15, 7, 21) {real, imag} */,
  {32'h3c77a16c, 32'hbe7d5cd6} /* (15, 7, 20) {real, imag} */,
  {32'h3d056e3c, 32'hbea966a8} /* (15, 7, 19) {real, imag} */,
  {32'hbe1891b0, 32'hbd8ecda0} /* (15, 7, 18) {real, imag} */,
  {32'h3dd3c8d6, 32'hbde792b3} /* (15, 7, 17) {real, imag} */,
  {32'h3e338f60, 32'hbd95410c} /* (15, 7, 16) {real, imag} */,
  {32'hbf24a7f4, 32'hbe7d1a4a} /* (15, 7, 15) {real, imag} */,
  {32'h3e3721ee, 32'h3e619244} /* (15, 7, 14) {real, imag} */,
  {32'hbddf3f45, 32'hbe271ed0} /* (15, 7, 13) {real, imag} */,
  {32'h3d5b1f98, 32'h3dda05a8} /* (15, 7, 12) {real, imag} */,
  {32'h3e5cd702, 32'h3e6b1839} /* (15, 7, 11) {real, imag} */,
  {32'hbe5579bb, 32'h3ea2093c} /* (15, 7, 10) {real, imag} */,
  {32'hbee65b4a, 32'h3e1e1e08} /* (15, 7, 9) {real, imag} */,
  {32'h3dc734d8, 32'hbf43afac} /* (15, 7, 8) {real, imag} */,
  {32'h3ee723e0, 32'h3ef2931c} /* (15, 7, 7) {real, imag} */,
  {32'hbf376059, 32'h3d8575c0} /* (15, 7, 6) {real, imag} */,
  {32'hbe8381b0, 32'h3d036770} /* (15, 7, 5) {real, imag} */,
  {32'h3e2a9560, 32'hbd8d7d96} /* (15, 7, 4) {real, imag} */,
  {32'hbe38fe40, 32'hbf1afd12} /* (15, 7, 3) {real, imag} */,
  {32'h3d865af0, 32'hbe64b8f3} /* (15, 7, 2) {real, imag} */,
  {32'hbef3f4ce, 32'h3fbbc676} /* (15, 7, 1) {real, imag} */,
  {32'hbe9173b2, 32'hbe33d8de} /* (15, 7, 0) {real, imag} */,
  {32'hbdae55e0, 32'h3e000aec} /* (15, 6, 31) {real, imag} */,
  {32'hbe8c4c8c, 32'h3daaa0e2} /* (15, 6, 30) {real, imag} */,
  {32'hbe14832c, 32'h3b1fe200} /* (15, 6, 29) {real, imag} */,
  {32'hbe197bfb, 32'h3dfe0b64} /* (15, 6, 28) {real, imag} */,
  {32'hbf05bbba, 32'h3d97e1ae} /* (15, 6, 27) {real, imag} */,
  {32'hbe92b338, 32'hbd64f512} /* (15, 6, 26) {real, imag} */,
  {32'hbf179a1a, 32'h3e32b79d} /* (15, 6, 25) {real, imag} */,
  {32'h3d2ab5d8, 32'hbed2285a} /* (15, 6, 24) {real, imag} */,
  {32'h3eb916e0, 32'hbe39addc} /* (15, 6, 23) {real, imag} */,
  {32'h3deb982c, 32'h3e3f6acd} /* (15, 6, 22) {real, imag} */,
  {32'hbe05623b, 32'h3e96834e} /* (15, 6, 21) {real, imag} */,
  {32'hbf2d6aca, 32'h3decd050} /* (15, 6, 20) {real, imag} */,
  {32'hbe9133e3, 32'hbe215578} /* (15, 6, 19) {real, imag} */,
  {32'h3eaa8d6e, 32'hbe09ad78} /* (15, 6, 18) {real, imag} */,
  {32'h3e2fda9a, 32'hbe3c33da} /* (15, 6, 17) {real, imag} */,
  {32'h3dafa00a, 32'h3ef42f66} /* (15, 6, 16) {real, imag} */,
  {32'h3e80214b, 32'hbe1a8350} /* (15, 6, 15) {real, imag} */,
  {32'h3d990b4e, 32'h3eb86f18} /* (15, 6, 14) {real, imag} */,
  {32'h3aba1ce0, 32'h3d559a68} /* (15, 6, 13) {real, imag} */,
  {32'h3da2c340, 32'h3e6fb8be} /* (15, 6, 12) {real, imag} */,
  {32'h3e32ad73, 32'h3e3177f8} /* (15, 6, 11) {real, imag} */,
  {32'hbe8c38f6, 32'h3f16ef9e} /* (15, 6, 10) {real, imag} */,
  {32'h3e9a7126, 32'h3e821f3a} /* (15, 6, 9) {real, imag} */,
  {32'hbf013df1, 32'hbe9cedeb} /* (15, 6, 8) {real, imag} */,
  {32'hbe18c8d2, 32'h3cd44c94} /* (15, 6, 7) {real, imag} */,
  {32'hbe3e2efe, 32'h3e97208e} /* (15, 6, 6) {real, imag} */,
  {32'h3ec72324, 32'hbe80d02c} /* (15, 6, 5) {real, imag} */,
  {32'hbec32d5e, 32'h3e0defba} /* (15, 6, 4) {real, imag} */,
  {32'h3ed64445, 32'h3e27c6c5} /* (15, 6, 3) {real, imag} */,
  {32'h3f2767b2, 32'h3f034c19} /* (15, 6, 2) {real, imag} */,
  {32'h3f277bff, 32'h3f55ce2e} /* (15, 6, 1) {real, imag} */,
  {32'hbf4276ba, 32'hbe7f1662} /* (15, 6, 0) {real, imag} */,
  {32'hbf91640a, 32'h3fbdcea6} /* (15, 5, 31) {real, imag} */,
  {32'h3df7cc00, 32'hbedb8776} /* (15, 5, 30) {real, imag} */,
  {32'h3d3fdc1c, 32'h3f20c403} /* (15, 5, 29) {real, imag} */,
  {32'h3dcd1a90, 32'h3cf79cb8} /* (15, 5, 28) {real, imag} */,
  {32'h3ec65102, 32'h3f62d8af} /* (15, 5, 27) {real, imag} */,
  {32'hbd14ffb4, 32'hbea86480} /* (15, 5, 26) {real, imag} */,
  {32'hbfa48c64, 32'h3e42bd64} /* (15, 5, 25) {real, imag} */,
  {32'hbec6b8e2, 32'hbd65e3b4} /* (15, 5, 24) {real, imag} */,
  {32'hbea1cadc, 32'h3dc791d8} /* (15, 5, 23) {real, imag} */,
  {32'h3e386be6, 32'hbee881ec} /* (15, 5, 22) {real, imag} */,
  {32'h3c258570, 32'h3d3f9576} /* (15, 5, 21) {real, imag} */,
  {32'hbdb0c4dc, 32'hbe35ca5f} /* (15, 5, 20) {real, imag} */,
  {32'hbd85f2a7, 32'hbd84c9bf} /* (15, 5, 19) {real, imag} */,
  {32'h3e456958, 32'hbd0869b4} /* (15, 5, 18) {real, imag} */,
  {32'hbe59b8a8, 32'hbee9f82a} /* (15, 5, 17) {real, imag} */,
  {32'hbe7eeb64, 32'hbd8219f4} /* (15, 5, 16) {real, imag} */,
  {32'h3efcbc4c, 32'h3d821428} /* (15, 5, 15) {real, imag} */,
  {32'hbeaa67df, 32'hbe23a5d1} /* (15, 5, 14) {real, imag} */,
  {32'hbe9c9fae, 32'hbd23f114} /* (15, 5, 13) {real, imag} */,
  {32'hbe0d3b8b, 32'hbe09d9dc} /* (15, 5, 12) {real, imag} */,
  {32'hbd93142e, 32'h3e6e9bb6} /* (15, 5, 11) {real, imag} */,
  {32'hbe1a2fca, 32'hbec9022a} /* (15, 5, 10) {real, imag} */,
  {32'hbea5f42a, 32'hbed96398} /* (15, 5, 9) {real, imag} */,
  {32'h3e237cce, 32'h3f4a2ad7} /* (15, 5, 8) {real, imag} */,
  {32'hbe0fb8ea, 32'hbda0ec10} /* (15, 5, 7) {real, imag} */,
  {32'h3e7ec830, 32'hbcf07600} /* (15, 5, 6) {real, imag} */,
  {32'h3e94528c, 32'h3e7739e2} /* (15, 5, 5) {real, imag} */,
  {32'h3f229328, 32'hbeb1d82c} /* (15, 5, 4) {real, imag} */,
  {32'h3f1041b0, 32'hbf15d2e4} /* (15, 5, 3) {real, imag} */,
  {32'h3e9b8e68, 32'h3f1f5f70} /* (15, 5, 2) {real, imag} */,
  {32'hbfd54f7e, 32'hbeb74c58} /* (15, 5, 1) {real, imag} */,
  {32'hbfc179e4, 32'hbdb8dc30} /* (15, 5, 0) {real, imag} */,
  {32'h3f9d9fbc, 32'h3d372c80} /* (15, 4, 31) {real, imag} */,
  {32'hbf1e6d60, 32'hbf16f5ba} /* (15, 4, 30) {real, imag} */,
  {32'h3db725e0, 32'hbf1e83b8} /* (15, 4, 29) {real, imag} */,
  {32'h3f806e5c, 32'h3f14af2e} /* (15, 4, 28) {real, imag} */,
  {32'hbf220fc4, 32'h3e229844} /* (15, 4, 27) {real, imag} */,
  {32'hbe910838, 32'h3f0d1f41} /* (15, 4, 26) {real, imag} */,
  {32'hbe8e1cb0, 32'h3f94df92} /* (15, 4, 25) {real, imag} */,
  {32'h3de33658, 32'hbc19cdc0} /* (15, 4, 24) {real, imag} */,
  {32'hbe234b2e, 32'hbd684f6e} /* (15, 4, 23) {real, imag} */,
  {32'hbd074bb6, 32'hbe47aa4c} /* (15, 4, 22) {real, imag} */,
  {32'h3cab2f62, 32'hbe28e580} /* (15, 4, 21) {real, imag} */,
  {32'hbbac5b70, 32'hbe4ebf23} /* (15, 4, 20) {real, imag} */,
  {32'hbeee9b47, 32'h3e2cf6d6} /* (15, 4, 19) {real, imag} */,
  {32'h3e4b6a14, 32'hbe4a8c5e} /* (15, 4, 18) {real, imag} */,
  {32'h3d92a4c6, 32'hbe2a39e5} /* (15, 4, 17) {real, imag} */,
  {32'hbe591c69, 32'hbe36950c} /* (15, 4, 16) {real, imag} */,
  {32'hbe02eb07, 32'h3f0e0cb9} /* (15, 4, 15) {real, imag} */,
  {32'hbe63e2d4, 32'hbe3d7ebd} /* (15, 4, 14) {real, imag} */,
  {32'h3ec316b5, 32'h3d707f50} /* (15, 4, 13) {real, imag} */,
  {32'h3d0ee8b4, 32'h3daaff94} /* (15, 4, 12) {real, imag} */,
  {32'h3ec0b383, 32'h3e36149a} /* (15, 4, 11) {real, imag} */,
  {32'h3ef0a6e2, 32'hbf06eef5} /* (15, 4, 10) {real, imag} */,
  {32'h3e34424c, 32'hbe454cbd} /* (15, 4, 9) {real, imag} */,
  {32'hbec52cb2, 32'hbe4349f0} /* (15, 4, 8) {real, imag} */,
  {32'h3ebdc926, 32'h3f673398} /* (15, 4, 7) {real, imag} */,
  {32'hbf413c7e, 32'hbf3b5633} /* (15, 4, 6) {real, imag} */,
  {32'hbf3be5f9, 32'hbed232e4} /* (15, 4, 5) {real, imag} */,
  {32'hbf04f422, 32'h3eac464b} /* (15, 4, 4) {real, imag} */,
  {32'hbf0ee141, 32'h3f3c9308} /* (15, 4, 3) {real, imag} */,
  {32'hbebdcab8, 32'hbfb6e4eb} /* (15, 4, 2) {real, imag} */,
  {32'h4047996a, 32'h3f1f55d5} /* (15, 4, 1) {real, imag} */,
  {32'hbf5c134a, 32'hbf98548b} /* (15, 4, 0) {real, imag} */,
  {32'h3f035fde, 32'hbab97800} /* (15, 3, 31) {real, imag} */,
  {32'h3fb7d485, 32'hbf1d1ab0} /* (15, 3, 30) {real, imag} */,
  {32'hbf571ca0, 32'hbe8c5562} /* (15, 3, 29) {real, imag} */,
  {32'h3f4f13ec, 32'h3ef940f6} /* (15, 3, 28) {real, imag} */,
  {32'hbe5d8e40, 32'h3eac4008} /* (15, 3, 27) {real, imag} */,
  {32'hbc49b4c0, 32'h3f387748} /* (15, 3, 26) {real, imag} */,
  {32'hbf2fa7cf, 32'h3cee18a0} /* (15, 3, 25) {real, imag} */,
  {32'hbef76c19, 32'hbebfae00} /* (15, 3, 24) {real, imag} */,
  {32'hbf0bfd10, 32'h3e530932} /* (15, 3, 23) {real, imag} */,
  {32'h3eabe82a, 32'hbe26f92a} /* (15, 3, 22) {real, imag} */,
  {32'hbdd7112c, 32'hbe95ea64} /* (15, 3, 21) {real, imag} */,
  {32'hbe60f4ea, 32'h3f38a196} /* (15, 3, 20) {real, imag} */,
  {32'hbd585dc6, 32'hbee7f592} /* (15, 3, 19) {real, imag} */,
  {32'h3dd418f0, 32'hbed54048} /* (15, 3, 18) {real, imag} */,
  {32'h3d42587c, 32'h3ef8e007} /* (15, 3, 17) {real, imag} */,
  {32'hbcd99f38, 32'hbe0d8b9c} /* (15, 3, 16) {real, imag} */,
  {32'hbe617484, 32'hbde14d6d} /* (15, 3, 15) {real, imag} */,
  {32'hbca1b824, 32'h3d0a287a} /* (15, 3, 14) {real, imag} */,
  {32'h3e88c562, 32'h3eb3722d} /* (15, 3, 13) {real, imag} */,
  {32'h3e11e365, 32'hbe3995d2} /* (15, 3, 12) {real, imag} */,
  {32'hbea7e2a5, 32'h3e9a2dd3} /* (15, 3, 11) {real, imag} */,
  {32'hbe179c0c, 32'h3e199ac6} /* (15, 3, 10) {real, imag} */,
  {32'hbeb71e38, 32'h3cf0825c} /* (15, 3, 9) {real, imag} */,
  {32'h3e073249, 32'hbe54793f} /* (15, 3, 8) {real, imag} */,
  {32'hbea05b99, 32'hbe81857c} /* (15, 3, 7) {real, imag} */,
  {32'hbe0373ec, 32'h3e4f5ec6} /* (15, 3, 6) {real, imag} */,
  {32'h3ebb5d54, 32'h3ec3e139} /* (15, 3, 5) {real, imag} */,
  {32'hbf12c4f2, 32'h3f6c8acc} /* (15, 3, 4) {real, imag} */,
  {32'h3e1d4050, 32'h3ef75db8} /* (15, 3, 3) {real, imag} */,
  {32'h3ec5a74e, 32'hbfa00cd7} /* (15, 3, 2) {real, imag} */,
  {32'h3fe87e13, 32'h3e20f4f0} /* (15, 3, 1) {real, imag} */,
  {32'h3ead938e, 32'h3f745722} /* (15, 3, 0) {real, imag} */,
  {32'hc11cc5a7, 32'hc01cc922} /* (15, 2, 31) {real, imag} */,
  {32'h40ba0394, 32'hbf94978c} /* (15, 2, 30) {real, imag} */,
  {32'h3f80f102, 32'h3f8c7ea2} /* (15, 2, 29) {real, imag} */,
  {32'hbf23d818, 32'h3fd85694} /* (15, 2, 28) {real, imag} */,
  {32'h3e83ec76, 32'hbe696154} /* (15, 2, 27) {real, imag} */,
  {32'hbf3bffd0, 32'h3f8c132a} /* (15, 2, 26) {real, imag} */,
  {32'hbe36ed96, 32'h3e156dc5} /* (15, 2, 25) {real, imag} */,
  {32'h3f012e38, 32'hbfb8869f} /* (15, 2, 24) {real, imag} */,
  {32'hbed177fa, 32'h3ef1ec78} /* (15, 2, 23) {real, imag} */,
  {32'h3e5e441a, 32'hbe44be1e} /* (15, 2, 22) {real, imag} */,
  {32'h3cee42e8, 32'hbe7aeb06} /* (15, 2, 21) {real, imag} */,
  {32'hbe7b40f8, 32'hbc309e00} /* (15, 2, 20) {real, imag} */,
  {32'hbe4ee376, 32'h3ea2f9d4} /* (15, 2, 19) {real, imag} */,
  {32'h3d422708, 32'h3e0be652} /* (15, 2, 18) {real, imag} */,
  {32'hbd766c02, 32'hbdc8f7fe} /* (15, 2, 17) {real, imag} */,
  {32'hbe3b5706, 32'hbe5d9872} /* (15, 2, 16) {real, imag} */,
  {32'h3c63c278, 32'hbe0d37ae} /* (15, 2, 15) {real, imag} */,
  {32'h3e3c4161, 32'h3ef96a64} /* (15, 2, 14) {real, imag} */,
  {32'h3e140144, 32'hbd30bfba} /* (15, 2, 13) {real, imag} */,
  {32'h3e0e462c, 32'h3ec86628} /* (15, 2, 12) {real, imag} */,
  {32'hbead1c62, 32'h3e90aedd} /* (15, 2, 11) {real, imag} */,
  {32'hbf0bedac, 32'hbe865a68} /* (15, 2, 10) {real, imag} */,
  {32'hbe8bf8c0, 32'h3e805efe} /* (15, 2, 9) {real, imag} */,
  {32'h3f718c62, 32'h3d718db0} /* (15, 2, 8) {real, imag} */,
  {32'hbbaab738, 32'h3e532c30} /* (15, 2, 7) {real, imag} */,
  {32'h3da0a6df, 32'h3ee4eab7} /* (15, 2, 6) {real, imag} */,
  {32'h3f3fdd0d, 32'h3fa79d04} /* (15, 2, 5) {real, imag} */,
  {32'h3e69a620, 32'hbffa85c9} /* (15, 2, 4) {real, imag} */,
  {32'h3f2b8b3f, 32'hbe8a9278} /* (15, 2, 3) {real, imag} */,
  {32'h406c5e68, 32'hbeb12d1c} /* (15, 2, 2) {real, imag} */,
  {32'hc09dbeae, 32'hbf2a6c18} /* (15, 2, 1) {real, imag} */,
  {32'hc0c446ee, 32'h3de18e20} /* (15, 2, 0) {real, imag} */,
  {32'h41560f50, 32'hc0886eb9} /* (15, 1, 31) {real, imag} */,
  {32'hc0904efa, 32'hbf98cc8b} /* (15, 1, 30) {real, imag} */,
  {32'hbe40fadc, 32'h3fff0978} /* (15, 1, 29) {real, imag} */,
  {32'h3fc58192, 32'hbf199196} /* (15, 1, 28) {real, imag} */,
  {32'hbfb10238, 32'h3f34d6e6} /* (15, 1, 27) {real, imag} */,
  {32'h3f573571, 32'hbef115ce} /* (15, 1, 26) {real, imag} */,
  {32'hbd90a002, 32'h3eea7351} /* (15, 1, 25) {real, imag} */,
  {32'hbec9a74e, 32'h3eb5d01a} /* (15, 1, 24) {real, imag} */,
  {32'hbec3235a, 32'h3f07b618} /* (15, 1, 23) {real, imag} */,
  {32'h3f07daa9, 32'hbe27086c} /* (15, 1, 22) {real, imag} */,
  {32'hbef64074, 32'h3e83b3d4} /* (15, 1, 21) {real, imag} */,
  {32'h3ee0bff3, 32'hbd4bd704} /* (15, 1, 20) {real, imag} */,
  {32'h3e426fe1, 32'h3f187dd0} /* (15, 1, 19) {real, imag} */,
  {32'hbdd63de8, 32'h3e8bc191} /* (15, 1, 18) {real, imag} */,
  {32'h3eaa92c4, 32'hbdd62f48} /* (15, 1, 17) {real, imag} */,
  {32'h3e2a6adf, 32'hbf0bfdf0} /* (15, 1, 16) {real, imag} */,
  {32'hbe7a9b04, 32'h3e8faaf0} /* (15, 1, 15) {real, imag} */,
  {32'h3ebef1c5, 32'hbe6f4662} /* (15, 1, 14) {real, imag} */,
  {32'h3ef7cc9e, 32'hbd10055a} /* (15, 1, 13) {real, imag} */,
  {32'hbe862490, 32'hbf133f61} /* (15, 1, 12) {real, imag} */,
  {32'hbe7318b2, 32'hbcd2feb0} /* (15, 1, 11) {real, imag} */,
  {32'h3d8bcd7e, 32'hbe8aad7a} /* (15, 1, 10) {real, imag} */,
  {32'h3caa78da, 32'h3e32ed53} /* (15, 1, 9) {real, imag} */,
  {32'hbf1c2dfb, 32'hbf215b96} /* (15, 1, 8) {real, imag} */,
  {32'h3f636749, 32'h3eb3a78e} /* (15, 1, 7) {real, imag} */,
  {32'h3edd400e, 32'hbef7816f} /* (15, 1, 6) {real, imag} */,
  {32'hbec70a0a, 32'hbea39f68} /* (15, 1, 5) {real, imag} */,
  {32'hbf40ee98, 32'h3fb0abe2} /* (15, 1, 4) {real, imag} */,
  {32'hbffe0c61, 32'h3e6f4938} /* (15, 1, 3) {real, imag} */,
  {32'hc0d82234, 32'hc0879866} /* (15, 1, 2) {real, imag} */,
  {32'h415eba7e, 32'h41276652} /* (15, 1, 1) {real, imag} */,
  {32'h4154b47b, 32'hc04e2f16} /* (15, 1, 0) {real, imag} */,
  {32'h4093a5c4, 32'hc0afeab8} /* (15, 0, 31) {real, imag} */,
  {32'hbf856028, 32'h405e8106} /* (15, 0, 30) {real, imag} */,
  {32'h3f5d4a56, 32'hbeba5708} /* (15, 0, 29) {real, imag} */,
  {32'hbfc5168a, 32'hbef64408} /* (15, 0, 28) {real, imag} */,
  {32'hbfb84eee, 32'hbe8f2b3e} /* (15, 0, 27) {real, imag} */,
  {32'h3e5598be, 32'h3e0df1cb} /* (15, 0, 26) {real, imag} */,
  {32'h3ee7edae, 32'hbf1d35cb} /* (15, 0, 25) {real, imag} */,
  {32'h3c3cd880, 32'h3eee44c6} /* (15, 0, 24) {real, imag} */,
  {32'hbda26794, 32'h3ba2be00} /* (15, 0, 23) {real, imag} */,
  {32'hbf0e0b00, 32'hbe1b5c34} /* (15, 0, 22) {real, imag} */,
  {32'hbe8fec97, 32'h3e60fa74} /* (15, 0, 21) {real, imag} */,
  {32'h3ee3f586, 32'hbc926744} /* (15, 0, 20) {real, imag} */,
  {32'hbee89efa, 32'h3e86d76a} /* (15, 0, 19) {real, imag} */,
  {32'h3d60407c, 32'h3f2086e4} /* (15, 0, 18) {real, imag} */,
  {32'h3dbabbb5, 32'h3ee647dd} /* (15, 0, 17) {real, imag} */,
  {32'h3ef51cb0, 32'h00000000} /* (15, 0, 16) {real, imag} */,
  {32'h3dbabbb5, 32'hbee647dd} /* (15, 0, 15) {real, imag} */,
  {32'h3d60407c, 32'hbf2086e4} /* (15, 0, 14) {real, imag} */,
  {32'hbee89efa, 32'hbe86d76a} /* (15, 0, 13) {real, imag} */,
  {32'h3ee3f586, 32'h3c926744} /* (15, 0, 12) {real, imag} */,
  {32'hbe8fec97, 32'hbe60fa74} /* (15, 0, 11) {real, imag} */,
  {32'hbf0e0b00, 32'h3e1b5c34} /* (15, 0, 10) {real, imag} */,
  {32'hbda26794, 32'hbba2be00} /* (15, 0, 9) {real, imag} */,
  {32'h3c3cd880, 32'hbeee44c6} /* (15, 0, 8) {real, imag} */,
  {32'h3ee7edae, 32'h3f1d35cb} /* (15, 0, 7) {real, imag} */,
  {32'h3e5598be, 32'hbe0df1cb} /* (15, 0, 6) {real, imag} */,
  {32'hbfb84eee, 32'h3e8f2b3e} /* (15, 0, 5) {real, imag} */,
  {32'hbfc5168a, 32'h3ef64408} /* (15, 0, 4) {real, imag} */,
  {32'h3f5d4a56, 32'h3eba5708} /* (15, 0, 3) {real, imag} */,
  {32'hbf856028, 32'hc05e8106} /* (15, 0, 2) {real, imag} */,
  {32'h4093a5c4, 32'h40afeab8} /* (15, 0, 1) {real, imag} */,
  {32'h4163b4ba, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h421b9faf, 32'hc1c42c5e} /* (14, 31, 31) {real, imag} */,
  {32'hc144f800, 32'h412c851c} /* (14, 31, 30) {real, imag} */,
  {32'hc05292c6, 32'h3eb46ae2} /* (14, 31, 29) {real, imag} */,
  {32'hbf81c90a, 32'hc00b4e7f} /* (14, 31, 28) {real, imag} */,
  {32'hbf8e2118, 32'h3f7e0fc7} /* (14, 31, 27) {real, imag} */,
  {32'h3dc62b18, 32'h3fc28469} /* (14, 31, 26) {real, imag} */,
  {32'h3f3ba0cb, 32'hbf75aa6e} /* (14, 31, 25) {real, imag} */,
  {32'hbf0d17b2, 32'h3ecc599e} /* (14, 31, 24) {real, imag} */,
  {32'hbd7adf00, 32'hbe706a1c} /* (14, 31, 23) {real, imag} */,
  {32'hbd8ad7d8, 32'h3e91c863} /* (14, 31, 22) {real, imag} */,
  {32'h3c49ea30, 32'h3f1c8435} /* (14, 31, 21) {real, imag} */,
  {32'h3e66d3df, 32'h3e4ee9a6} /* (14, 31, 20) {real, imag} */,
  {32'h3f25bc2e, 32'hbb26aab0} /* (14, 31, 19) {real, imag} */,
  {32'hbd90b127, 32'h3ef1a5a8} /* (14, 31, 18) {real, imag} */,
  {32'hbe37a2e6, 32'hbe169be0} /* (14, 31, 17) {real, imag} */,
  {32'h3e4fc513, 32'h3e05c5da} /* (14, 31, 16) {real, imag} */,
  {32'hbdea6e9e, 32'hbe6b499e} /* (14, 31, 15) {real, imag} */,
  {32'hbd614204, 32'hbea444f4} /* (14, 31, 14) {real, imag} */,
  {32'hbd548f88, 32'h3e0c41e0} /* (14, 31, 13) {real, imag} */,
  {32'hbe0537a0, 32'h3e0bb386} /* (14, 31, 12) {real, imag} */,
  {32'hbeeb1256, 32'hbf7b4b94} /* (14, 31, 11) {real, imag} */,
  {32'h3e8330a7, 32'h3dcfd346} /* (14, 31, 10) {real, imag} */,
  {32'hbebd07ec, 32'h3ddcc148} /* (14, 31, 9) {real, imag} */,
  {32'hbf8962fe, 32'hbd8a0b3c} /* (14, 31, 8) {real, imag} */,
  {32'h3b342880, 32'hbf6734e8} /* (14, 31, 7) {real, imag} */,
  {32'h3f3c57f6, 32'h3e36ba80} /* (14, 31, 6) {real, imag} */,
  {32'hc021f3d4, 32'hbf173340} /* (14, 31, 5) {real, imag} */,
  {32'h400bda14, 32'h3e32bcd8} /* (14, 31, 4) {real, imag} */,
  {32'h3de25e82, 32'hbff86364} /* (14, 31, 3) {real, imag} */,
  {32'hc10f225e, 32'h3f0fbbcb} /* (14, 31, 2) {real, imag} */,
  {32'h41f54011, 32'h41019160} /* (14, 31, 1) {real, imag} */,
  {32'h420aa966, 32'h3effab80} /* (14, 31, 0) {real, imag} */,
  {32'hc15ce4b0, 32'hbf9bfa32} /* (14, 30, 31) {real, imag} */,
  {32'h40fef71b, 32'h3f5b8362} /* (14, 30, 30) {real, imag} */,
  {32'h3e3e1bd8, 32'hbe26f602} /* (14, 30, 29) {real, imag} */,
  {32'hbfba6fd8, 32'h3ff90b6e} /* (14, 30, 28) {real, imag} */,
  {32'h3fd387d8, 32'hc01dad09} /* (14, 30, 27) {real, imag} */,
  {32'hbecbac48, 32'hbf9a9d6f} /* (14, 30, 26) {real, imag} */,
  {32'hbcb66040, 32'hbe1e00c3} /* (14, 30, 25) {real, imag} */,
  {32'h3fc0d158, 32'hbeee1d02} /* (14, 30, 24) {real, imag} */,
  {32'h3d0ca328, 32'hbec5aa72} /* (14, 30, 23) {real, imag} */,
  {32'hbcf19170, 32'hbdf8a7ac} /* (14, 30, 22) {real, imag} */,
  {32'h3e7ab9d2, 32'hbf01fa44} /* (14, 30, 21) {real, imag} */,
  {32'hbd71e780, 32'h3e95bf64} /* (14, 30, 20) {real, imag} */,
  {32'hbf130e4a, 32'hbea8162b} /* (14, 30, 19) {real, imag} */,
  {32'h3f3ce754, 32'hbdd52982} /* (14, 30, 18) {real, imag} */,
  {32'hbce46878, 32'hbd6e0fb6} /* (14, 30, 17) {real, imag} */,
  {32'h3d5507f8, 32'h3e323628} /* (14, 30, 16) {real, imag} */,
  {32'h3e798700, 32'hbf04d02c} /* (14, 30, 15) {real, imag} */,
  {32'h3e492458, 32'h3f103a1c} /* (14, 30, 14) {real, imag} */,
  {32'hbe9fbfbf, 32'hbea6809e} /* (14, 30, 13) {real, imag} */,
  {32'h3e626fd6, 32'h3eb8df83} /* (14, 30, 12) {real, imag} */,
  {32'h3debe5cd, 32'h3e0c533c} /* (14, 30, 11) {real, imag} */,
  {32'h3e2e2cb8, 32'hbef7ca5b} /* (14, 30, 10) {real, imag} */,
  {32'h3db2944b, 32'h3edeecb2} /* (14, 30, 9) {real, imag} */,
  {32'h3e1c9cd3, 32'h3ee373d8} /* (14, 30, 8) {real, imag} */,
  {32'hbf4cc744, 32'hbe95f5cf} /* (14, 30, 7) {real, imag} */,
  {32'h3ddfc6a8, 32'h3f390066} /* (14, 30, 6) {real, imag} */,
  {32'h3fbbefd2, 32'h3efe4132} /* (14, 30, 5) {real, imag} */,
  {32'hbfcfb7b5, 32'hc0296ac6} /* (14, 30, 4) {real, imag} */,
  {32'h3eb84045, 32'hbed4297a} /* (14, 30, 3) {real, imag} */,
  {32'h414a1049, 32'h409496c6} /* (14, 30, 2) {real, imag} */,
  {32'hc1c04433, 32'h40000be0} /* (14, 30, 1) {real, imag} */,
  {32'hc14edef5, 32'h3ff91f82} /* (14, 30, 0) {real, imag} */,
  {32'h405aa10d, 32'hc00aa287} /* (14, 29, 31) {real, imag} */,
  {32'hbf57d97b, 32'h3ffeee7a} /* (14, 29, 30) {real, imag} */,
  {32'h3f10bc2d, 32'hbec550dc} /* (14, 29, 29) {real, imag} */,
  {32'hbe744766, 32'hbf22b238} /* (14, 29, 28) {real, imag} */,
  {32'h3e2551f8, 32'hbf8a92a0} /* (14, 29, 27) {real, imag} */,
  {32'h3c9e43c0, 32'h3e274f0c} /* (14, 29, 26) {real, imag} */,
  {32'h3f45b8bc, 32'h3e43492c} /* (14, 29, 25) {real, imag} */,
  {32'h3ebe50a5, 32'hbcc78ec0} /* (14, 29, 24) {real, imag} */,
  {32'hbe5f326e, 32'h3f6ef5bc} /* (14, 29, 23) {real, imag} */,
  {32'hbd9a3350, 32'hbe1a661c} /* (14, 29, 22) {real, imag} */,
  {32'h3ebf6950, 32'hbf0759ef} /* (14, 29, 21) {real, imag} */,
  {32'h3da80470, 32'hbda5163c} /* (14, 29, 20) {real, imag} */,
  {32'hbd039296, 32'h3d641104} /* (14, 29, 19) {real, imag} */,
  {32'h3e9e6c95, 32'hbdd18254} /* (14, 29, 18) {real, imag} */,
  {32'hbe56e812, 32'hbe8848bc} /* (14, 29, 17) {real, imag} */,
  {32'hbe050566, 32'hbd4aaae0} /* (14, 29, 16) {real, imag} */,
  {32'hbdc96dfb, 32'hbd26038c} /* (14, 29, 15) {real, imag} */,
  {32'hbd762d7f, 32'h3e2ea436} /* (14, 29, 14) {real, imag} */,
  {32'h3eac1c13, 32'h3e1b2ac4} /* (14, 29, 13) {real, imag} */,
  {32'h3e9a6fe2, 32'hbeba8d5e} /* (14, 29, 12) {real, imag} */,
  {32'hbeb6a7db, 32'h3ebb18dc} /* (14, 29, 11) {real, imag} */,
  {32'hbe9849e9, 32'hbf3f51fd} /* (14, 29, 10) {real, imag} */,
  {32'hbf259772, 32'h3e695803} /* (14, 29, 9) {real, imag} */,
  {32'hbebdad1d, 32'h3e8d8afe} /* (14, 29, 8) {real, imag} */,
  {32'hbde11cb9, 32'h3e719618} /* (14, 29, 7) {real, imag} */,
  {32'hbe8bb090, 32'h3dd29ec8} /* (14, 29, 6) {real, imag} */,
  {32'hbf181f2e, 32'h3e848d60} /* (14, 29, 5) {real, imag} */,
  {32'h3f4bba10, 32'hbf0aeab8} /* (14, 29, 4) {real, imag} */,
  {32'hbe9d9938, 32'hbf794558} /* (14, 29, 3) {real, imag} */,
  {32'h400c3096, 32'h3fd49870} /* (14, 29, 2) {real, imag} */,
  {32'hc0204d1c, 32'hbfb015a3} /* (14, 29, 1) {real, imag} */,
  {32'h3f23d1be, 32'hbe522f1e} /* (14, 29, 0) {real, imag} */,
  {32'h40a1860a, 32'hbf5fed02} /* (14, 28, 31) {real, imag} */,
  {32'hbffd71c0, 32'h4000cfd4} /* (14, 28, 30) {real, imag} */,
  {32'hbecc4708, 32'hbf36cea1} /* (14, 28, 29) {real, imag} */,
  {32'h3efd4c94, 32'hbf6268e5} /* (14, 28, 28) {real, imag} */,
  {32'hbf204ab9, 32'h3ed4b97a} /* (14, 28, 27) {real, imag} */,
  {32'hbf245d95, 32'hbf15fbc3} /* (14, 28, 26) {real, imag} */,
  {32'hbe22d18d, 32'hbdd598ec} /* (14, 28, 25) {real, imag} */,
  {32'hbe0b8abd, 32'hbe76d71a} /* (14, 28, 24) {real, imag} */,
  {32'h3f95c679, 32'h3e5725db} /* (14, 28, 23) {real, imag} */,
  {32'h3e9ff1de, 32'hbf2cefd6} /* (14, 28, 22) {real, imag} */,
  {32'hbe723ae4, 32'h3de38603} /* (14, 28, 21) {real, imag} */,
  {32'h3ce7cb54, 32'h3ddc865c} /* (14, 28, 20) {real, imag} */,
  {32'hbe4545e5, 32'hbe1355fe} /* (14, 28, 19) {real, imag} */,
  {32'hbe2ec4c5, 32'h3ef42284} /* (14, 28, 18) {real, imag} */,
  {32'hbd5a3196, 32'h3eeed944} /* (14, 28, 17) {real, imag} */,
  {32'h3dd3392a, 32'h3c219e58} /* (14, 28, 16) {real, imag} */,
  {32'hbe9c6e6b, 32'hbe951f59} /* (14, 28, 15) {real, imag} */,
  {32'hbe4ca6f4, 32'hbdd820bd} /* (14, 28, 14) {real, imag} */,
  {32'hbede1de1, 32'h3f07f8f1} /* (14, 28, 13) {real, imag} */,
  {32'h3d417eec, 32'hbde6af62} /* (14, 28, 12) {real, imag} */,
  {32'hbe796f88, 32'hbdfa4d25} /* (14, 28, 11) {real, imag} */,
  {32'hbe3a6203, 32'hbdd15d70} /* (14, 28, 10) {real, imag} */,
  {32'hbdaf57e4, 32'h3e942478} /* (14, 28, 9) {real, imag} */,
  {32'hbec1fbbe, 32'hbe7e98f2} /* (14, 28, 8) {real, imag} */,
  {32'hbe7e5b74, 32'hbf8cc61a} /* (14, 28, 7) {real, imag} */,
  {32'hbdcecff4, 32'hbee4c278} /* (14, 28, 6) {real, imag} */,
  {32'hbf144570, 32'hbf3fcf1e} /* (14, 28, 5) {real, imag} */,
  {32'h3f528d42, 32'hbfb1772c} /* (14, 28, 4) {real, imag} */,
  {32'hbefd9df8, 32'h3e927616} /* (14, 28, 3) {real, imag} */,
  {32'hbfcf7cae, 32'h401f0bce} /* (14, 28, 2) {real, imag} */,
  {32'h400f529d, 32'hbf5443c0} /* (14, 28, 1) {real, imag} */,
  {32'hbdd038b8, 32'h3f363da8} /* (14, 28, 0) {real, imag} */,
  {32'hc04d3d71, 32'h3f248e40} /* (14, 27, 31) {real, imag} */,
  {32'hbb06c500, 32'hbede278c} /* (14, 27, 30) {real, imag} */,
  {32'hbddc9e28, 32'hbd8d9280} /* (14, 27, 29) {real, imag} */,
  {32'h3e72bc27, 32'h3ef0e036} /* (14, 27, 28) {real, imag} */,
  {32'h3eda6178, 32'hbf2e6b49} /* (14, 27, 27) {real, imag} */,
  {32'h3ec5672d, 32'h3c915b80} /* (14, 27, 26) {real, imag} */,
  {32'hbe59279e, 32'hbc641dd8} /* (14, 27, 25) {real, imag} */,
  {32'hbeebae52, 32'hbec67e9e} /* (14, 27, 24) {real, imag} */,
  {32'h3d87d2b4, 32'h3d8eb2d8} /* (14, 27, 23) {real, imag} */,
  {32'h3d725186, 32'hbef725a7} /* (14, 27, 22) {real, imag} */,
  {32'hbd016d0e, 32'h3ce85bc0} /* (14, 27, 21) {real, imag} */,
  {32'hbea1158d, 32'hbe037c86} /* (14, 27, 20) {real, imag} */,
  {32'h3ebf3c45, 32'h3e17a45a} /* (14, 27, 19) {real, imag} */,
  {32'h3bb56860, 32'hbefcd092} /* (14, 27, 18) {real, imag} */,
  {32'h3e5b2fab, 32'h3d5b4002} /* (14, 27, 17) {real, imag} */,
  {32'hbd53ad4e, 32'h3e08e3d4} /* (14, 27, 16) {real, imag} */,
  {32'h3e1313db, 32'hbdb6a100} /* (14, 27, 15) {real, imag} */,
  {32'h3e974fbe, 32'h3e6312c4} /* (14, 27, 14) {real, imag} */,
  {32'hbc5a2e8a, 32'hbdc2ad0c} /* (14, 27, 13) {real, imag} */,
  {32'hbe2c88ba, 32'h3d5e12dc} /* (14, 27, 12) {real, imag} */,
  {32'h3e8b0d2c, 32'h3caa6d28} /* (14, 27, 11) {real, imag} */,
  {32'hbbdedee0, 32'h3d73fd54} /* (14, 27, 10) {real, imag} */,
  {32'h3daf7814, 32'h3d4058d5} /* (14, 27, 9) {real, imag} */,
  {32'h3e0be2f0, 32'hbd0f8218} /* (14, 27, 8) {real, imag} */,
  {32'hbe17b01e, 32'hbe83c661} /* (14, 27, 7) {real, imag} */,
  {32'hbe85c78e, 32'hbe395292} /* (14, 27, 6) {real, imag} */,
  {32'h3f212148, 32'h3e857d60} /* (14, 27, 5) {real, imag} */,
  {32'hbe83166e, 32'h3e101be0} /* (14, 27, 4) {real, imag} */,
  {32'hbe9bf32b, 32'hbf213c4d} /* (14, 27, 3) {real, imag} */,
  {32'h3e3f196c, 32'hbe99df2d} /* (14, 27, 2) {real, imag} */,
  {32'hc00a8fb9, 32'hbf906b62} /* (14, 27, 1) {real, imag} */,
  {32'hc002f9fd, 32'h3fa03f75} /* (14, 27, 0) {real, imag} */,
  {32'hbee50a4d, 32'h3b9fa320} /* (14, 26, 31) {real, imag} */,
  {32'h3f64a15d, 32'hbe87f3d8} /* (14, 26, 30) {real, imag} */,
  {32'h3e103f6c, 32'hbf1dd5dc} /* (14, 26, 29) {real, imag} */,
  {32'hbea4bb72, 32'hbe41714b} /* (14, 26, 28) {real, imag} */,
  {32'h3cc130a8, 32'h3f268dfc} /* (14, 26, 27) {real, imag} */,
  {32'hbecdae02, 32'hbe070fd2} /* (14, 26, 26) {real, imag} */,
  {32'hbd15af88, 32'h3ea3e626} /* (14, 26, 25) {real, imag} */,
  {32'h3e5c6480, 32'hbe9f0860} /* (14, 26, 24) {real, imag} */,
  {32'hbeaabd29, 32'hbe80f859} /* (14, 26, 23) {real, imag} */,
  {32'h3f11b883, 32'hbd7ffbc2} /* (14, 26, 22) {real, imag} */,
  {32'h3ed0c398, 32'h3e8f4176} /* (14, 26, 21) {real, imag} */,
  {32'h3e773050, 32'h3e4a2770} /* (14, 26, 20) {real, imag} */,
  {32'h3da955b4, 32'h3d87b2a4} /* (14, 26, 19) {real, imag} */,
  {32'hbedfa61c, 32'hbc2e2298} /* (14, 26, 18) {real, imag} */,
  {32'h3e87bd8f, 32'hbdae5980} /* (14, 26, 17) {real, imag} */,
  {32'hbbcb79b8, 32'h3ce26804} /* (14, 26, 16) {real, imag} */,
  {32'hbdaf6a21, 32'h3efe59a8} /* (14, 26, 15) {real, imag} */,
  {32'h3d9cf1fa, 32'h3e998f25} /* (14, 26, 14) {real, imag} */,
  {32'h3e577f42, 32'h3ed26a7a} /* (14, 26, 13) {real, imag} */,
  {32'hbd58aac8, 32'hbf1249e2} /* (14, 26, 12) {real, imag} */,
  {32'hbe08f2e9, 32'hbe9cdd25} /* (14, 26, 11) {real, imag} */,
  {32'hbe293bda, 32'h3f09bc72} /* (14, 26, 10) {real, imag} */,
  {32'h3e6789e5, 32'hbf103725} /* (14, 26, 9) {real, imag} */,
  {32'hbd877de8, 32'hbe8768ad} /* (14, 26, 8) {real, imag} */,
  {32'hbf293a68, 32'h3f7e66ad} /* (14, 26, 7) {real, imag} */,
  {32'h3e5abdea, 32'hbf3663df} /* (14, 26, 6) {real, imag} */,
  {32'hbe94de72, 32'hbe5e7216} /* (14, 26, 5) {real, imag} */,
  {32'hbeccac08, 32'h3e83f7fe} /* (14, 26, 4) {real, imag} */,
  {32'hbf8a773c, 32'h3f070b6e} /* (14, 26, 3) {real, imag} */,
  {32'h3f493076, 32'hbe254934} /* (14, 26, 2) {real, imag} */,
  {32'h3eac37d9, 32'hbe93cbb8} /* (14, 26, 1) {real, imag} */,
  {32'hbeb24388, 32'hbdf0aaa4} /* (14, 26, 0) {real, imag} */,
  {32'hbe751c4e, 32'hbf636c2e} /* (14, 25, 31) {real, imag} */,
  {32'h3e156b2c, 32'h3f1833ce} /* (14, 25, 30) {real, imag} */,
  {32'hbe08a118, 32'h3e7f7a2c} /* (14, 25, 29) {real, imag} */,
  {32'hbf6e6cac, 32'hbf04a701} /* (14, 25, 28) {real, imag} */,
  {32'hbe89f044, 32'h3e16c99a} /* (14, 25, 27) {real, imag} */,
  {32'h3eabf63a, 32'h3eac81a8} /* (14, 25, 26) {real, imag} */,
  {32'hbe6db2b6, 32'h3eda94f4} /* (14, 25, 25) {real, imag} */,
  {32'h3e95c152, 32'h3f30954c} /* (14, 25, 24) {real, imag} */,
  {32'hbea9c79b, 32'h3f1a7a14} /* (14, 25, 23) {real, imag} */,
  {32'hbd337cac, 32'hbf33a45c} /* (14, 25, 22) {real, imag} */,
  {32'hbe1670a6, 32'hbe05bc8b} /* (14, 25, 21) {real, imag} */,
  {32'hbf0a9490, 32'hbeff0658} /* (14, 25, 20) {real, imag} */,
  {32'h3d4d5a2c, 32'hbf432e6d} /* (14, 25, 19) {real, imag} */,
  {32'hbe26c378, 32'hbc15b040} /* (14, 25, 18) {real, imag} */,
  {32'h3e83890f, 32'hbe25e198} /* (14, 25, 17) {real, imag} */,
  {32'h3ea9d26c, 32'hbee68c96} /* (14, 25, 16) {real, imag} */,
  {32'h3ea04da6, 32'h3d20e598} /* (14, 25, 15) {real, imag} */,
  {32'hbe0fd3ed, 32'h3d71fa00} /* (14, 25, 14) {real, imag} */,
  {32'h3eab7bc6, 32'hbe98d94d} /* (14, 25, 13) {real, imag} */,
  {32'h3f369b24, 32'h3f5b02b9} /* (14, 25, 12) {real, imag} */,
  {32'h3eacba39, 32'h3e3c2ff9} /* (14, 25, 11) {real, imag} */,
  {32'h3e884198, 32'hbdc70696} /* (14, 25, 10) {real, imag} */,
  {32'hbe8ee0e5, 32'hbe859fef} /* (14, 25, 9) {real, imag} */,
  {32'hbcdffd68, 32'h3d5b750a} /* (14, 25, 8) {real, imag} */,
  {32'hbe9c5816, 32'hbe00fda0} /* (14, 25, 7) {real, imag} */,
  {32'hbf28b55b, 32'h3d7f4468} /* (14, 25, 6) {real, imag} */,
  {32'hbf07d4d8, 32'hbf6bc854} /* (14, 25, 5) {real, imag} */,
  {32'hbe8eef98, 32'h3ea59c4d} /* (14, 25, 4) {real, imag} */,
  {32'h3df65ea0, 32'h3e00ace5} /* (14, 25, 3) {real, imag} */,
  {32'hbe210d46, 32'h3f6a0730} /* (14, 25, 2) {real, imag} */,
  {32'h3f664b91, 32'h3f28ec68} /* (14, 25, 1) {real, imag} */,
  {32'hbd71350c, 32'hbf9d80aa} /* (14, 25, 0) {real, imag} */,
  {32'hbf2ea470, 32'h3f8a9226} /* (14, 24, 31) {real, imag} */,
  {32'h3f365f51, 32'hbdee5a60} /* (14, 24, 30) {real, imag} */,
  {32'hbe30765f, 32'hbe41c104} /* (14, 24, 29) {real, imag} */,
  {32'hbf4c9cd6, 32'hbd887159} /* (14, 24, 28) {real, imag} */,
  {32'hbd7f0ef6, 32'hbf488ef6} /* (14, 24, 27) {real, imag} */,
  {32'h3d9923af, 32'hbd3254ec} /* (14, 24, 26) {real, imag} */,
  {32'h3e88f3c7, 32'hbe46f734} /* (14, 24, 25) {real, imag} */,
  {32'hbcadb8c0, 32'hbb8b3bc0} /* (14, 24, 24) {real, imag} */,
  {32'hbe4f55fd, 32'hbdc4726f} /* (14, 24, 23) {real, imag} */,
  {32'hbf63d422, 32'hbe46dfd0} /* (14, 24, 22) {real, imag} */,
  {32'h3f10ff78, 32'h3e6c41ea} /* (14, 24, 21) {real, imag} */,
  {32'hbeb784c2, 32'h3eb50657} /* (14, 24, 20) {real, imag} */,
  {32'hbcac4510, 32'h3e3c17f3} /* (14, 24, 19) {real, imag} */,
  {32'h3e19a760, 32'hbe1b7eae} /* (14, 24, 18) {real, imag} */,
  {32'hbe994266, 32'h3ef160dd} /* (14, 24, 17) {real, imag} */,
  {32'hbe5b26aa, 32'hbe53c248} /* (14, 24, 16) {real, imag} */,
  {32'hbe06c192, 32'hbeaa9510} /* (14, 24, 15) {real, imag} */,
  {32'h3cb1ff88, 32'h3d26cf1c} /* (14, 24, 14) {real, imag} */,
  {32'h3dd579c4, 32'hbea86238} /* (14, 24, 13) {real, imag} */,
  {32'hbec012a8, 32'hbe33907d} /* (14, 24, 12) {real, imag} */,
  {32'h3ed0918c, 32'h3cc4b998} /* (14, 24, 11) {real, imag} */,
  {32'h3e30e129, 32'h3f11a2dc} /* (14, 24, 10) {real, imag} */,
  {32'hbdbe9ce8, 32'h3ed26e8f} /* (14, 24, 9) {real, imag} */,
  {32'h3b8a84e8, 32'h3e4b9b90} /* (14, 24, 8) {real, imag} */,
  {32'h3ecd44c3, 32'hbe0da6a8} /* (14, 24, 7) {real, imag} */,
  {32'h3ee1e62d, 32'hbd27a084} /* (14, 24, 6) {real, imag} */,
  {32'h3f404486, 32'h3d06343a} /* (14, 24, 5) {real, imag} */,
  {32'hbeb93fa0, 32'hbe9ca426} /* (14, 24, 4) {real, imag} */,
  {32'h3ebf9e15, 32'h3e6f409a} /* (14, 24, 3) {real, imag} */,
  {32'h3f2eaa56, 32'hbf198e3b} /* (14, 24, 2) {real, imag} */,
  {32'hc00b4cde, 32'h3f9379d5} /* (14, 24, 1) {real, imag} */,
  {32'hbf3a0d4e, 32'h3e64e9e6} /* (14, 24, 0) {real, imag} */,
  {32'h3d1144c0, 32'h3d72ffb8} /* (14, 23, 31) {real, imag} */,
  {32'h3e16cdaf, 32'h3e57fdf8} /* (14, 23, 30) {real, imag} */,
  {32'hbe727797, 32'hbe9d50a5} /* (14, 23, 29) {real, imag} */,
  {32'hbe3b1f17, 32'hbec99d1d} /* (14, 23, 28) {real, imag} */,
  {32'h3ebdc41b, 32'h3ebab2c3} /* (14, 23, 27) {real, imag} */,
  {32'hbe21a11a, 32'h3f1afbba} /* (14, 23, 26) {real, imag} */,
  {32'hbf3582ae, 32'hbe91940a} /* (14, 23, 25) {real, imag} */,
  {32'hbed8d8f3, 32'hbec7ad17} /* (14, 23, 24) {real, imag} */,
  {32'h3e5a1cc1, 32'h3d8b4bec} /* (14, 23, 23) {real, imag} */,
  {32'hbe00633b, 32'hbeefc54c} /* (14, 23, 22) {real, imag} */,
  {32'hbe91e473, 32'hbec988be} /* (14, 23, 21) {real, imag} */,
  {32'hbe941b13, 32'h3e41febe} /* (14, 23, 20) {real, imag} */,
  {32'h3e4d795c, 32'h3e980da8} /* (14, 23, 19) {real, imag} */,
  {32'hbea31163, 32'hbcfc4b64} /* (14, 23, 18) {real, imag} */,
  {32'hbd000f72, 32'h3f06e588} /* (14, 23, 17) {real, imag} */,
  {32'hbe1735ab, 32'hbdae30ec} /* (14, 23, 16) {real, imag} */,
  {32'hbea7d911, 32'h3e6a68e0} /* (14, 23, 15) {real, imag} */,
  {32'h3f2a6e97, 32'h3f172b7f} /* (14, 23, 14) {real, imag} */,
  {32'h3f115c1c, 32'h3ede164f} /* (14, 23, 13) {real, imag} */,
  {32'hbdcf694a, 32'hbc5b8520} /* (14, 23, 12) {real, imag} */,
  {32'hbf361464, 32'hbea6f738} /* (14, 23, 11) {real, imag} */,
  {32'hbeb91550, 32'hbe7a17ce} /* (14, 23, 10) {real, imag} */,
  {32'hbe83d0fb, 32'h3db8e3e4} /* (14, 23, 9) {real, imag} */,
  {32'h3e49773a, 32'h3e9ecf6c} /* (14, 23, 8) {real, imag} */,
  {32'h3f4c817f, 32'hbe963ba8} /* (14, 23, 7) {real, imag} */,
  {32'h3e833108, 32'h3dc45c80} /* (14, 23, 6) {real, imag} */,
  {32'hbf261ebf, 32'h3eb8b3c8} /* (14, 23, 5) {real, imag} */,
  {32'h3ec414a9, 32'hbe5fa954} /* (14, 23, 4) {real, imag} */,
  {32'h3e809193, 32'hbdea286f} /* (14, 23, 3) {real, imag} */,
  {32'hbd97aa20, 32'h3eeeec56} /* (14, 23, 2) {real, imag} */,
  {32'hbe259db5, 32'hbf05d1b4} /* (14, 23, 1) {real, imag} */,
  {32'h3e6f8717, 32'hbe34ceba} /* (14, 23, 0) {real, imag} */,
  {32'h3f670a46, 32'hbe0f2d3b} /* (14, 22, 31) {real, imag} */,
  {32'hbe389566, 32'h3d08d198} /* (14, 22, 30) {real, imag} */,
  {32'hbe094436, 32'hbe197633} /* (14, 22, 29) {real, imag} */,
  {32'hbd14d510, 32'h3f1810cc} /* (14, 22, 28) {real, imag} */,
  {32'h3ef8faf0, 32'h3b217f00} /* (14, 22, 27) {real, imag} */,
  {32'h3e8955ea, 32'hbd7669ec} /* (14, 22, 26) {real, imag} */,
  {32'h3ea36ee6, 32'hbdb3e555} /* (14, 22, 25) {real, imag} */,
  {32'hbd7b5fc8, 32'h3d3ef619} /* (14, 22, 24) {real, imag} */,
  {32'h3e02e1b3, 32'h3f04af94} /* (14, 22, 23) {real, imag} */,
  {32'h3da70212, 32'h3ee86cb2} /* (14, 22, 22) {real, imag} */,
  {32'h3f148a6d, 32'h3d9fa698} /* (14, 22, 21) {real, imag} */,
  {32'h3c6a5ca0, 32'hbeb39646} /* (14, 22, 20) {real, imag} */,
  {32'hbde25868, 32'h3ee45687} /* (14, 22, 19) {real, imag} */,
  {32'h3d663f28, 32'hbe38e038} /* (14, 22, 18) {real, imag} */,
  {32'hbf0e4ea6, 32'hbed1fe88} /* (14, 22, 17) {real, imag} */,
  {32'hbe82234b, 32'h3e990e8d} /* (14, 22, 16) {real, imag} */,
  {32'h3e248a77, 32'h3f25e7c5} /* (14, 22, 15) {real, imag} */,
  {32'h3e01dda2, 32'h3d81bd8e} /* (14, 22, 14) {real, imag} */,
  {32'hbe60b663, 32'hbda56ee2} /* (14, 22, 13) {real, imag} */,
  {32'hbb5116e0, 32'h3ea2dc9c} /* (14, 22, 12) {real, imag} */,
  {32'h3e0b2ac3, 32'h3ee69055} /* (14, 22, 11) {real, imag} */,
  {32'h3cf6f910, 32'hbdfcdb92} /* (14, 22, 10) {real, imag} */,
  {32'h3e955a53, 32'hbf3c4af6} /* (14, 22, 9) {real, imag} */,
  {32'hbeaa9ed4, 32'hbe9acb56} /* (14, 22, 8) {real, imag} */,
  {32'h3f2ea7ae, 32'hbf42a69e} /* (14, 22, 7) {real, imag} */,
  {32'h3f3985d9, 32'hbe1a9b70} /* (14, 22, 6) {real, imag} */,
  {32'hbe81bdd8, 32'h3e5d8994} /* (14, 22, 5) {real, imag} */,
  {32'hbf2a1715, 32'hbe1f50f4} /* (14, 22, 4) {real, imag} */,
  {32'hbdae4d7a, 32'hbcb60260} /* (14, 22, 3) {real, imag} */,
  {32'h3dd79e20, 32'h3f30250c} /* (14, 22, 2) {real, imag} */,
  {32'hbe12e34a, 32'hbe8f28c3} /* (14, 22, 1) {real, imag} */,
  {32'h3ea29090, 32'hbf4efe2b} /* (14, 22, 0) {real, imag} */,
  {32'h3cab12da, 32'h3f7baf2a} /* (14, 21, 31) {real, imag} */,
  {32'hbd945138, 32'hbed5eb35} /* (14, 21, 30) {real, imag} */,
  {32'hbe1daa61, 32'hbe8076b6} /* (14, 21, 29) {real, imag} */,
  {32'h3d7baf97, 32'h3e904fba} /* (14, 21, 28) {real, imag} */,
  {32'hbe1754a3, 32'hbe642ca6} /* (14, 21, 27) {real, imag} */,
  {32'h3f02d79c, 32'hbedc5786} /* (14, 21, 26) {real, imag} */,
  {32'h3ed775a8, 32'hbefafa1b} /* (14, 21, 25) {real, imag} */,
  {32'h3dc5fc20, 32'hbe1d54b8} /* (14, 21, 24) {real, imag} */,
  {32'hbe2aeb46, 32'h3ce00658} /* (14, 21, 23) {real, imag} */,
  {32'h3df9b8a2, 32'h3f3622c2} /* (14, 21, 22) {real, imag} */,
  {32'hbe5aef2a, 32'h3eed6f43} /* (14, 21, 21) {real, imag} */,
  {32'h3e703928, 32'h3ddddc29} /* (14, 21, 20) {real, imag} */,
  {32'h3eea0856, 32'h3d8f1dea} /* (14, 21, 19) {real, imag} */,
  {32'h3ef90ef0, 32'hbee2ec17} /* (14, 21, 18) {real, imag} */,
  {32'h3e84cf07, 32'hbd68e494} /* (14, 21, 17) {real, imag} */,
  {32'hbefab361, 32'h3d40e98a} /* (14, 21, 16) {real, imag} */,
  {32'hbe3f3d1a, 32'hbd8ee391} /* (14, 21, 15) {real, imag} */,
  {32'h3dd86fe5, 32'h3c90166e} /* (14, 21, 14) {real, imag} */,
  {32'hbf018b8d, 32'hbe89ce17} /* (14, 21, 13) {real, imag} */,
  {32'hbe352ea2, 32'hbe171131} /* (14, 21, 12) {real, imag} */,
  {32'h3eb30e8a, 32'hbf39a82d} /* (14, 21, 11) {real, imag} */,
  {32'hbc7fe100, 32'h3e22f092} /* (14, 21, 10) {real, imag} */,
  {32'h3eed133e, 32'h3ee5aad3} /* (14, 21, 9) {real, imag} */,
  {32'h3ed44e2f, 32'h3f0e26d8} /* (14, 21, 8) {real, imag} */,
  {32'h3e9027f2, 32'h3ee1efce} /* (14, 21, 7) {real, imag} */,
  {32'hbd91eb64, 32'h3e310b6b} /* (14, 21, 6) {real, imag} */,
  {32'h3f44d613, 32'hbf0eda24} /* (14, 21, 5) {real, imag} */,
  {32'hbcfdeb44, 32'hbe8658b2} /* (14, 21, 4) {real, imag} */,
  {32'hbf0ca28e, 32'hbcf8ba58} /* (14, 21, 3) {real, imag} */,
  {32'hbdb0a0e4, 32'hbf18fa90} /* (14, 21, 2) {real, imag} */,
  {32'hbf443bc0, 32'h3dead3be} /* (14, 21, 1) {real, imag} */,
  {32'hbf106db5, 32'h3f766e78} /* (14, 21, 0) {real, imag} */,
  {32'h3f00fceb, 32'hbdcc4d48} /* (14, 20, 31) {real, imag} */,
  {32'h3e05882c, 32'hbcd641f0} /* (14, 20, 30) {real, imag} */,
  {32'hbde8c3eb, 32'hbea5ac4a} /* (14, 20, 29) {real, imag} */,
  {32'h3ec6ac00, 32'h3e33d437} /* (14, 20, 28) {real, imag} */,
  {32'hbe119b36, 32'hbd11d10d} /* (14, 20, 27) {real, imag} */,
  {32'h3df1a94f, 32'h3eb914c1} /* (14, 20, 26) {real, imag} */,
  {32'h3ed09ac1, 32'hbd4c4e50} /* (14, 20, 25) {real, imag} */,
  {32'hbeabab96, 32'h3e9a2f5c} /* (14, 20, 24) {real, imag} */,
  {32'hbe8fed94, 32'hbf1568eb} /* (14, 20, 23) {real, imag} */,
  {32'hbe22390f, 32'hbe394af9} /* (14, 20, 22) {real, imag} */,
  {32'hbe977a16, 32'hbdeecae2} /* (14, 20, 21) {real, imag} */,
  {32'hbebc2880, 32'h3e7daffe} /* (14, 20, 20) {real, imag} */,
  {32'hbbc50088, 32'h3e584515} /* (14, 20, 19) {real, imag} */,
  {32'hbe2d15f8, 32'h3da3df9a} /* (14, 20, 18) {real, imag} */,
  {32'hbec24eaf, 32'h3d95fac4} /* (14, 20, 17) {real, imag} */,
  {32'hbd43a4ec, 32'h3dbd1d18} /* (14, 20, 16) {real, imag} */,
  {32'hbe9fa2d2, 32'h3cc1ef8e} /* (14, 20, 15) {real, imag} */,
  {32'hbdeef3c0, 32'h3e8befa5} /* (14, 20, 14) {real, imag} */,
  {32'h3e9e32d6, 32'hbefd7a7e} /* (14, 20, 13) {real, imag} */,
  {32'hbeeac9f4, 32'hbdad35da} /* (14, 20, 12) {real, imag} */,
  {32'h3e6b8024, 32'h3e5726a7} /* (14, 20, 11) {real, imag} */,
  {32'h3e82973a, 32'h3d5213bc} /* (14, 20, 10) {real, imag} */,
  {32'hbe7be71f, 32'hbe0b31d6} /* (14, 20, 9) {real, imag} */,
  {32'h3ec091b1, 32'hbe6bd58c} /* (14, 20, 8) {real, imag} */,
  {32'h3d1cfaae, 32'h3e9ec116} /* (14, 20, 7) {real, imag} */,
  {32'hbe94b019, 32'hbe016204} /* (14, 20, 6) {real, imag} */,
  {32'h3d6c36fe, 32'h3ec7e1b3} /* (14, 20, 5) {real, imag} */,
  {32'h3db4dfe9, 32'h3e8d1f42} /* (14, 20, 4) {real, imag} */,
  {32'h3cedff10, 32'h3dd7e6ee} /* (14, 20, 3) {real, imag} */,
  {32'h3e11835f, 32'hbf14468e} /* (14, 20, 2) {real, imag} */,
  {32'hbe64bf90, 32'hbd30e358} /* (14, 20, 1) {real, imag} */,
  {32'h3ed0862e, 32'h3e24bb46} /* (14, 20, 0) {real, imag} */,
  {32'h3e850d3c, 32'hbecbedda} /* (14, 19, 31) {real, imag} */,
  {32'h3e31d12c, 32'hbe6a931b} /* (14, 19, 30) {real, imag} */,
  {32'h3ad5cbe0, 32'hbe6c8c86} /* (14, 19, 29) {real, imag} */,
  {32'hbe4ff28f, 32'hbd5b15a0} /* (14, 19, 28) {real, imag} */,
  {32'hbdcbd2c4, 32'hbe9a3d0f} /* (14, 19, 27) {real, imag} */,
  {32'h3e564742, 32'h3e6a1520} /* (14, 19, 26) {real, imag} */,
  {32'hbd44980c, 32'h3d65c6ac} /* (14, 19, 25) {real, imag} */,
  {32'hbe1f361f, 32'hbe3ad620} /* (14, 19, 24) {real, imag} */,
  {32'hbe4296f8, 32'hbe1212bc} /* (14, 19, 23) {real, imag} */,
  {32'h3e5d079c, 32'h3e00f852} /* (14, 19, 22) {real, imag} */,
  {32'hbd3345d0, 32'h3eaad11c} /* (14, 19, 21) {real, imag} */,
  {32'hbceedd6c, 32'hbf061bb1} /* (14, 19, 20) {real, imag} */,
  {32'h3c7d4a70, 32'hbe259fc9} /* (14, 19, 19) {real, imag} */,
  {32'h3efe3368, 32'h3e825e56} /* (14, 19, 18) {real, imag} */,
  {32'hbf45d546, 32'hbe0c5787} /* (14, 19, 17) {real, imag} */,
  {32'h3dd8d8ac, 32'hbe1ae742} /* (14, 19, 16) {real, imag} */,
  {32'h3d987ce6, 32'hbe6c2d28} /* (14, 19, 15) {real, imag} */,
  {32'hbf063cd1, 32'h3ea7723e} /* (14, 19, 14) {real, imag} */,
  {32'hbee9dcd9, 32'h3e6c664a} /* (14, 19, 13) {real, imag} */,
  {32'h3edfb897, 32'h3efab5b4} /* (14, 19, 12) {real, imag} */,
  {32'h3dedafc9, 32'hbde580c8} /* (14, 19, 11) {real, imag} */,
  {32'hbe013e79, 32'hbe5ce3de} /* (14, 19, 10) {real, imag} */,
  {32'hbe6248c9, 32'hbe894285} /* (14, 19, 9) {real, imag} */,
  {32'hbd90cd97, 32'hbb9dace0} /* (14, 19, 8) {real, imag} */,
  {32'h3ecc208f, 32'hbcaedd70} /* (14, 19, 7) {real, imag} */,
  {32'hbee75cca, 32'h3f18c5a4} /* (14, 19, 6) {real, imag} */,
  {32'hbf092253, 32'h3e096ad0} /* (14, 19, 5) {real, imag} */,
  {32'h3dd3c1f5, 32'h3e37be22} /* (14, 19, 4) {real, imag} */,
  {32'h3d74d69e, 32'h3e3bfe9a} /* (14, 19, 3) {real, imag} */,
  {32'hbd73304a, 32'hbe69b071} /* (14, 19, 2) {real, imag} */,
  {32'h39d2d700, 32'h3eae2e74} /* (14, 19, 1) {real, imag} */,
  {32'hbf046821, 32'hbe7289fa} /* (14, 19, 0) {real, imag} */,
  {32'hbcc08828, 32'h3ebd712e} /* (14, 18, 31) {real, imag} */,
  {32'hbeae7ff9, 32'hbf1a24c6} /* (14, 18, 30) {real, imag} */,
  {32'h3ea96f4a, 32'h3dbf4790} /* (14, 18, 29) {real, imag} */,
  {32'hbe070ba9, 32'h3dcf86c6} /* (14, 18, 28) {real, imag} */,
  {32'hbdc3c230, 32'h3e52649e} /* (14, 18, 27) {real, imag} */,
  {32'h3ea61c82, 32'hbec6b524} /* (14, 18, 26) {real, imag} */,
  {32'hbeb9afc6, 32'h3cd3f450} /* (14, 18, 25) {real, imag} */,
  {32'hbe481cf9, 32'h3ea58db0} /* (14, 18, 24) {real, imag} */,
  {32'hbe8e67cd, 32'h3d9d5d0c} /* (14, 18, 23) {real, imag} */,
  {32'h3f38424a, 32'h3e89969e} /* (14, 18, 22) {real, imag} */,
  {32'h3eadd80a, 32'h3e99cafa} /* (14, 18, 21) {real, imag} */,
  {32'h3e9af5d1, 32'h3d9286ac} /* (14, 18, 20) {real, imag} */,
  {32'h3e1ef2a2, 32'h3f08ca88} /* (14, 18, 19) {real, imag} */,
  {32'h3eff1194, 32'h3d3d0df8} /* (14, 18, 18) {real, imag} */,
  {32'h3e95d91b, 32'hbcab82e0} /* (14, 18, 17) {real, imag} */,
  {32'h3d5dbe32, 32'hbd95ec8c} /* (14, 18, 16) {real, imag} */,
  {32'h3f550c56, 32'hbe21e6bc} /* (14, 18, 15) {real, imag} */,
  {32'h3f1a3c40, 32'hbe872e9e} /* (14, 18, 14) {real, imag} */,
  {32'hbd8bcdf0, 32'hbeb705a2} /* (14, 18, 13) {real, imag} */,
  {32'h3df7ff15, 32'hbe66a297} /* (14, 18, 12) {real, imag} */,
  {32'h3dcd408e, 32'h3e829b12} /* (14, 18, 11) {real, imag} */,
  {32'hbef181a8, 32'h3dfbab6e} /* (14, 18, 10) {real, imag} */,
  {32'hbde2104e, 32'h3ed0b406} /* (14, 18, 9) {real, imag} */,
  {32'hbed52756, 32'h3e4d9b58} /* (14, 18, 8) {real, imag} */,
  {32'hbe56ff30, 32'h3eab995e} /* (14, 18, 7) {real, imag} */,
  {32'h3f38f986, 32'hbd6978b1} /* (14, 18, 6) {real, imag} */,
  {32'hbd8f7a2e, 32'h3ebb15d4} /* (14, 18, 5) {real, imag} */,
  {32'h3e31745c, 32'hbe8f3ab9} /* (14, 18, 4) {real, imag} */,
  {32'hbd6d6c8a, 32'hbdd85e70} /* (14, 18, 3) {real, imag} */,
  {32'hbe416bf7, 32'h3c29f5f8} /* (14, 18, 2) {real, imag} */,
  {32'hbe73e3a1, 32'h3ea97002} /* (14, 18, 1) {real, imag} */,
  {32'hbd320d0c, 32'h3dd66b82} /* (14, 18, 0) {real, imag} */,
  {32'h3e225ee0, 32'hbe65b531} /* (14, 17, 31) {real, imag} */,
  {32'hbd48ffee, 32'h3d6cc0c0} /* (14, 17, 30) {real, imag} */,
  {32'h3ed5405b, 32'hbe0b2d48} /* (14, 17, 29) {real, imag} */,
  {32'hbd53dc0a, 32'h3e01c56d} /* (14, 17, 28) {real, imag} */,
  {32'hbe6c9e2c, 32'h3e9cbcd4} /* (14, 17, 27) {real, imag} */,
  {32'hbe093268, 32'hbe5566c8} /* (14, 17, 26) {real, imag} */,
  {32'hbc94fe98, 32'hbe2f02a1} /* (14, 17, 25) {real, imag} */,
  {32'h3edc1589, 32'hbdf0f942} /* (14, 17, 24) {real, imag} */,
  {32'h3eb6a390, 32'hbe7d3f63} /* (14, 17, 23) {real, imag} */,
  {32'h3e1f2fe8, 32'h3d929914} /* (14, 17, 22) {real, imag} */,
  {32'hbb3f4ec0, 32'hbde04242} /* (14, 17, 21) {real, imag} */,
  {32'h3ce32658, 32'h3eadbed0} /* (14, 17, 20) {real, imag} */,
  {32'h3c726280, 32'h3d4db3d0} /* (14, 17, 19) {real, imag} */,
  {32'hbdc719b6, 32'h3e9d8547} /* (14, 17, 18) {real, imag} */,
  {32'hbdd3e797, 32'h3d021152} /* (14, 17, 17) {real, imag} */,
  {32'h3c063834, 32'h3e9e5da7} /* (14, 17, 16) {real, imag} */,
  {32'h3c232620, 32'h3eb24c42} /* (14, 17, 15) {real, imag} */,
  {32'hbe788386, 32'h3d66e62c} /* (14, 17, 14) {real, imag} */,
  {32'hbef27710, 32'h3e00cd18} /* (14, 17, 13) {real, imag} */,
  {32'hbe3eaf50, 32'hbd790bd0} /* (14, 17, 12) {real, imag} */,
  {32'h3e338b8a, 32'hbec55026} /* (14, 17, 11) {real, imag} */,
  {32'h3e837e0b, 32'hbdd314e5} /* (14, 17, 10) {real, imag} */,
  {32'hbdc1941c, 32'hbca176b0} /* (14, 17, 9) {real, imag} */,
  {32'hbcd33504, 32'h3eba0931} /* (14, 17, 8) {real, imag} */,
  {32'hbe3bf4e1, 32'h3db81332} /* (14, 17, 7) {real, imag} */,
  {32'hbe8fadc1, 32'h3ed99cc6} /* (14, 17, 6) {real, imag} */,
  {32'hbddce9c6, 32'hbdb7ac25} /* (14, 17, 5) {real, imag} */,
  {32'hbd6f5589, 32'hbeb8e043} /* (14, 17, 4) {real, imag} */,
  {32'h3e85718e, 32'hbe8b85cb} /* (14, 17, 3) {real, imag} */,
  {32'hbdd54486, 32'hbd5ef4d0} /* (14, 17, 2) {real, imag} */,
  {32'h3ddd73f4, 32'hbe23013e} /* (14, 17, 1) {real, imag} */,
  {32'hbea65459, 32'hbe4861aa} /* (14, 17, 0) {real, imag} */,
  {32'h3d9825b8, 32'h3dde34c7} /* (14, 16, 31) {real, imag} */,
  {32'hbe957375, 32'hbdd68c54} /* (14, 16, 30) {real, imag} */,
  {32'hbe5670b2, 32'hbd41e020} /* (14, 16, 29) {real, imag} */,
  {32'h3e5b552e, 32'h3e5d02f8} /* (14, 16, 28) {real, imag} */,
  {32'h3d14c8e1, 32'h3dd4dc5a} /* (14, 16, 27) {real, imag} */,
  {32'hbd81aa3d, 32'h3e02d6d8} /* (14, 16, 26) {real, imag} */,
  {32'h3db5329d, 32'hbd4867c0} /* (14, 16, 25) {real, imag} */,
  {32'hbdcf12f6, 32'hbd491dfc} /* (14, 16, 24) {real, imag} */,
  {32'h3d2a85ad, 32'hbd268b9c} /* (14, 16, 23) {real, imag} */,
  {32'h3e7f0d25, 32'h3ee018b0} /* (14, 16, 22) {real, imag} */,
  {32'h3e354561, 32'hbec7adcf} /* (14, 16, 21) {real, imag} */,
  {32'hbe1039f0, 32'hbdafbb12} /* (14, 16, 20) {real, imag} */,
  {32'hbe8a03c6, 32'h3e858d41} /* (14, 16, 19) {real, imag} */,
  {32'h3c996eec, 32'hbe06b67c} /* (14, 16, 18) {real, imag} */,
  {32'hbe1f3ff2, 32'hbea14de1} /* (14, 16, 17) {real, imag} */,
  {32'hbe768552, 32'h00000000} /* (14, 16, 16) {real, imag} */,
  {32'hbe1f3ff2, 32'h3ea14de1} /* (14, 16, 15) {real, imag} */,
  {32'h3c996eec, 32'h3e06b67c} /* (14, 16, 14) {real, imag} */,
  {32'hbe8a03c6, 32'hbe858d41} /* (14, 16, 13) {real, imag} */,
  {32'hbe1039f0, 32'h3dafbb12} /* (14, 16, 12) {real, imag} */,
  {32'h3e354561, 32'h3ec7adcf} /* (14, 16, 11) {real, imag} */,
  {32'h3e7f0d25, 32'hbee018b0} /* (14, 16, 10) {real, imag} */,
  {32'h3d2a85ad, 32'h3d268b9c} /* (14, 16, 9) {real, imag} */,
  {32'hbdcf12f6, 32'h3d491dfc} /* (14, 16, 8) {real, imag} */,
  {32'h3db5329d, 32'h3d4867c0} /* (14, 16, 7) {real, imag} */,
  {32'hbd81aa3d, 32'hbe02d6d8} /* (14, 16, 6) {real, imag} */,
  {32'h3d14c8e1, 32'hbdd4dc5a} /* (14, 16, 5) {real, imag} */,
  {32'h3e5b552e, 32'hbe5d02f8} /* (14, 16, 4) {real, imag} */,
  {32'hbe5670b2, 32'h3d41e020} /* (14, 16, 3) {real, imag} */,
  {32'hbe957375, 32'h3dd68c54} /* (14, 16, 2) {real, imag} */,
  {32'h3d9825b8, 32'hbdde34c7} /* (14, 16, 1) {real, imag} */,
  {32'h3e699a4c, 32'h00000000} /* (14, 16, 0) {real, imag} */,
  {32'h3ddd73f4, 32'h3e23013e} /* (14, 15, 31) {real, imag} */,
  {32'hbdd54486, 32'h3d5ef4d0} /* (14, 15, 30) {real, imag} */,
  {32'h3e85718e, 32'h3e8b85cb} /* (14, 15, 29) {real, imag} */,
  {32'hbd6f5589, 32'h3eb8e043} /* (14, 15, 28) {real, imag} */,
  {32'hbddce9c6, 32'h3db7ac25} /* (14, 15, 27) {real, imag} */,
  {32'hbe8fadc1, 32'hbed99cc6} /* (14, 15, 26) {real, imag} */,
  {32'hbe3bf4e1, 32'hbdb81332} /* (14, 15, 25) {real, imag} */,
  {32'hbcd33504, 32'hbeba0931} /* (14, 15, 24) {real, imag} */,
  {32'hbdc1941c, 32'h3ca176b0} /* (14, 15, 23) {real, imag} */,
  {32'h3e837e0b, 32'h3dd314e5} /* (14, 15, 22) {real, imag} */,
  {32'h3e338b8a, 32'h3ec55026} /* (14, 15, 21) {real, imag} */,
  {32'hbe3eaf50, 32'h3d790bd0} /* (14, 15, 20) {real, imag} */,
  {32'hbef27710, 32'hbe00cd18} /* (14, 15, 19) {real, imag} */,
  {32'hbe788386, 32'hbd66e62c} /* (14, 15, 18) {real, imag} */,
  {32'h3c232620, 32'hbeb24c42} /* (14, 15, 17) {real, imag} */,
  {32'h3c063834, 32'hbe9e5da7} /* (14, 15, 16) {real, imag} */,
  {32'hbdd3e797, 32'hbd021152} /* (14, 15, 15) {real, imag} */,
  {32'hbdc719b6, 32'hbe9d8547} /* (14, 15, 14) {real, imag} */,
  {32'h3c726280, 32'hbd4db3d0} /* (14, 15, 13) {real, imag} */,
  {32'h3ce32658, 32'hbeadbed0} /* (14, 15, 12) {real, imag} */,
  {32'hbb3f4ec0, 32'h3de04242} /* (14, 15, 11) {real, imag} */,
  {32'h3e1f2fe8, 32'hbd929914} /* (14, 15, 10) {real, imag} */,
  {32'h3eb6a390, 32'h3e7d3f63} /* (14, 15, 9) {real, imag} */,
  {32'h3edc1589, 32'h3df0f942} /* (14, 15, 8) {real, imag} */,
  {32'hbc94fe98, 32'h3e2f02a1} /* (14, 15, 7) {real, imag} */,
  {32'hbe093268, 32'h3e5566c8} /* (14, 15, 6) {real, imag} */,
  {32'hbe6c9e2c, 32'hbe9cbcd4} /* (14, 15, 5) {real, imag} */,
  {32'hbd53dc0a, 32'hbe01c56d} /* (14, 15, 4) {real, imag} */,
  {32'h3ed5405b, 32'h3e0b2d48} /* (14, 15, 3) {real, imag} */,
  {32'hbd48ffee, 32'hbd6cc0c0} /* (14, 15, 2) {real, imag} */,
  {32'h3e225ee0, 32'h3e65b531} /* (14, 15, 1) {real, imag} */,
  {32'hbea65459, 32'h3e4861aa} /* (14, 15, 0) {real, imag} */,
  {32'hbe73e3a1, 32'hbea97002} /* (14, 14, 31) {real, imag} */,
  {32'hbe416bf7, 32'hbc29f5f8} /* (14, 14, 30) {real, imag} */,
  {32'hbd6d6c8a, 32'h3dd85e70} /* (14, 14, 29) {real, imag} */,
  {32'h3e31745c, 32'h3e8f3ab9} /* (14, 14, 28) {real, imag} */,
  {32'hbd8f7a2e, 32'hbebb15d4} /* (14, 14, 27) {real, imag} */,
  {32'h3f38f986, 32'h3d6978b1} /* (14, 14, 26) {real, imag} */,
  {32'hbe56ff30, 32'hbeab995e} /* (14, 14, 25) {real, imag} */,
  {32'hbed52756, 32'hbe4d9b58} /* (14, 14, 24) {real, imag} */,
  {32'hbde2104e, 32'hbed0b406} /* (14, 14, 23) {real, imag} */,
  {32'hbef181a8, 32'hbdfbab6e} /* (14, 14, 22) {real, imag} */,
  {32'h3dcd408e, 32'hbe829b12} /* (14, 14, 21) {real, imag} */,
  {32'h3df7ff15, 32'h3e66a297} /* (14, 14, 20) {real, imag} */,
  {32'hbd8bcdf0, 32'h3eb705a2} /* (14, 14, 19) {real, imag} */,
  {32'h3f1a3c40, 32'h3e872e9e} /* (14, 14, 18) {real, imag} */,
  {32'h3f550c56, 32'h3e21e6bc} /* (14, 14, 17) {real, imag} */,
  {32'h3d5dbe32, 32'h3d95ec8c} /* (14, 14, 16) {real, imag} */,
  {32'h3e95d91b, 32'h3cab82e0} /* (14, 14, 15) {real, imag} */,
  {32'h3eff1194, 32'hbd3d0df8} /* (14, 14, 14) {real, imag} */,
  {32'h3e1ef2a2, 32'hbf08ca88} /* (14, 14, 13) {real, imag} */,
  {32'h3e9af5d1, 32'hbd9286ac} /* (14, 14, 12) {real, imag} */,
  {32'h3eadd80a, 32'hbe99cafa} /* (14, 14, 11) {real, imag} */,
  {32'h3f38424a, 32'hbe89969e} /* (14, 14, 10) {real, imag} */,
  {32'hbe8e67cd, 32'hbd9d5d0c} /* (14, 14, 9) {real, imag} */,
  {32'hbe481cf9, 32'hbea58db0} /* (14, 14, 8) {real, imag} */,
  {32'hbeb9afc6, 32'hbcd3f450} /* (14, 14, 7) {real, imag} */,
  {32'h3ea61c82, 32'h3ec6b524} /* (14, 14, 6) {real, imag} */,
  {32'hbdc3c230, 32'hbe52649e} /* (14, 14, 5) {real, imag} */,
  {32'hbe070ba9, 32'hbdcf86c6} /* (14, 14, 4) {real, imag} */,
  {32'h3ea96f4a, 32'hbdbf4790} /* (14, 14, 3) {real, imag} */,
  {32'hbeae7ff9, 32'h3f1a24c6} /* (14, 14, 2) {real, imag} */,
  {32'hbcc08828, 32'hbebd712e} /* (14, 14, 1) {real, imag} */,
  {32'hbd320d0c, 32'hbdd66b82} /* (14, 14, 0) {real, imag} */,
  {32'h39d2d700, 32'hbeae2e74} /* (14, 13, 31) {real, imag} */,
  {32'hbd73304a, 32'h3e69b071} /* (14, 13, 30) {real, imag} */,
  {32'h3d74d69e, 32'hbe3bfe9a} /* (14, 13, 29) {real, imag} */,
  {32'h3dd3c1f5, 32'hbe37be22} /* (14, 13, 28) {real, imag} */,
  {32'hbf092253, 32'hbe096ad0} /* (14, 13, 27) {real, imag} */,
  {32'hbee75cca, 32'hbf18c5a4} /* (14, 13, 26) {real, imag} */,
  {32'h3ecc208f, 32'h3caedd70} /* (14, 13, 25) {real, imag} */,
  {32'hbd90cd97, 32'h3b9dace0} /* (14, 13, 24) {real, imag} */,
  {32'hbe6248c9, 32'h3e894285} /* (14, 13, 23) {real, imag} */,
  {32'hbe013e79, 32'h3e5ce3de} /* (14, 13, 22) {real, imag} */,
  {32'h3dedafc9, 32'h3de580c8} /* (14, 13, 21) {real, imag} */,
  {32'h3edfb897, 32'hbefab5b4} /* (14, 13, 20) {real, imag} */,
  {32'hbee9dcd9, 32'hbe6c664a} /* (14, 13, 19) {real, imag} */,
  {32'hbf063cd1, 32'hbea7723e} /* (14, 13, 18) {real, imag} */,
  {32'h3d987ce6, 32'h3e6c2d28} /* (14, 13, 17) {real, imag} */,
  {32'h3dd8d8ac, 32'h3e1ae742} /* (14, 13, 16) {real, imag} */,
  {32'hbf45d546, 32'h3e0c5787} /* (14, 13, 15) {real, imag} */,
  {32'h3efe3368, 32'hbe825e56} /* (14, 13, 14) {real, imag} */,
  {32'h3c7d4a70, 32'h3e259fc9} /* (14, 13, 13) {real, imag} */,
  {32'hbceedd6c, 32'h3f061bb1} /* (14, 13, 12) {real, imag} */,
  {32'hbd3345d0, 32'hbeaad11c} /* (14, 13, 11) {real, imag} */,
  {32'h3e5d079c, 32'hbe00f852} /* (14, 13, 10) {real, imag} */,
  {32'hbe4296f8, 32'h3e1212bc} /* (14, 13, 9) {real, imag} */,
  {32'hbe1f361f, 32'h3e3ad620} /* (14, 13, 8) {real, imag} */,
  {32'hbd44980c, 32'hbd65c6ac} /* (14, 13, 7) {real, imag} */,
  {32'h3e564742, 32'hbe6a1520} /* (14, 13, 6) {real, imag} */,
  {32'hbdcbd2c4, 32'h3e9a3d0f} /* (14, 13, 5) {real, imag} */,
  {32'hbe4ff28f, 32'h3d5b15a0} /* (14, 13, 4) {real, imag} */,
  {32'h3ad5cbe0, 32'h3e6c8c86} /* (14, 13, 3) {real, imag} */,
  {32'h3e31d12c, 32'h3e6a931b} /* (14, 13, 2) {real, imag} */,
  {32'h3e850d3c, 32'h3ecbedda} /* (14, 13, 1) {real, imag} */,
  {32'hbf046821, 32'h3e7289fa} /* (14, 13, 0) {real, imag} */,
  {32'hbe64bf90, 32'h3d30e358} /* (14, 12, 31) {real, imag} */,
  {32'h3e11835f, 32'h3f14468e} /* (14, 12, 30) {real, imag} */,
  {32'h3cedff10, 32'hbdd7e6ee} /* (14, 12, 29) {real, imag} */,
  {32'h3db4dfe9, 32'hbe8d1f42} /* (14, 12, 28) {real, imag} */,
  {32'h3d6c36fe, 32'hbec7e1b3} /* (14, 12, 27) {real, imag} */,
  {32'hbe94b019, 32'h3e016204} /* (14, 12, 26) {real, imag} */,
  {32'h3d1cfaae, 32'hbe9ec116} /* (14, 12, 25) {real, imag} */,
  {32'h3ec091b1, 32'h3e6bd58c} /* (14, 12, 24) {real, imag} */,
  {32'hbe7be71f, 32'h3e0b31d6} /* (14, 12, 23) {real, imag} */,
  {32'h3e82973a, 32'hbd5213bc} /* (14, 12, 22) {real, imag} */,
  {32'h3e6b8024, 32'hbe5726a7} /* (14, 12, 21) {real, imag} */,
  {32'hbeeac9f4, 32'h3dad35da} /* (14, 12, 20) {real, imag} */,
  {32'h3e9e32d6, 32'h3efd7a7e} /* (14, 12, 19) {real, imag} */,
  {32'hbdeef3c0, 32'hbe8befa5} /* (14, 12, 18) {real, imag} */,
  {32'hbe9fa2d2, 32'hbcc1ef8e} /* (14, 12, 17) {real, imag} */,
  {32'hbd43a4ec, 32'hbdbd1d18} /* (14, 12, 16) {real, imag} */,
  {32'hbec24eaf, 32'hbd95fac4} /* (14, 12, 15) {real, imag} */,
  {32'hbe2d15f8, 32'hbda3df9a} /* (14, 12, 14) {real, imag} */,
  {32'hbbc50088, 32'hbe584515} /* (14, 12, 13) {real, imag} */,
  {32'hbebc2880, 32'hbe7daffe} /* (14, 12, 12) {real, imag} */,
  {32'hbe977a16, 32'h3deecae2} /* (14, 12, 11) {real, imag} */,
  {32'hbe22390f, 32'h3e394af9} /* (14, 12, 10) {real, imag} */,
  {32'hbe8fed94, 32'h3f1568eb} /* (14, 12, 9) {real, imag} */,
  {32'hbeabab96, 32'hbe9a2f5c} /* (14, 12, 8) {real, imag} */,
  {32'h3ed09ac1, 32'h3d4c4e50} /* (14, 12, 7) {real, imag} */,
  {32'h3df1a94f, 32'hbeb914c1} /* (14, 12, 6) {real, imag} */,
  {32'hbe119b36, 32'h3d11d10d} /* (14, 12, 5) {real, imag} */,
  {32'h3ec6ac00, 32'hbe33d437} /* (14, 12, 4) {real, imag} */,
  {32'hbde8c3eb, 32'h3ea5ac4a} /* (14, 12, 3) {real, imag} */,
  {32'h3e05882c, 32'h3cd641f0} /* (14, 12, 2) {real, imag} */,
  {32'h3f00fceb, 32'h3dcc4d48} /* (14, 12, 1) {real, imag} */,
  {32'h3ed0862e, 32'hbe24bb46} /* (14, 12, 0) {real, imag} */,
  {32'hbf443bc0, 32'hbdead3be} /* (14, 11, 31) {real, imag} */,
  {32'hbdb0a0e4, 32'h3f18fa90} /* (14, 11, 30) {real, imag} */,
  {32'hbf0ca28e, 32'h3cf8ba58} /* (14, 11, 29) {real, imag} */,
  {32'hbcfdeb44, 32'h3e8658b2} /* (14, 11, 28) {real, imag} */,
  {32'h3f44d613, 32'h3f0eda24} /* (14, 11, 27) {real, imag} */,
  {32'hbd91eb64, 32'hbe310b6b} /* (14, 11, 26) {real, imag} */,
  {32'h3e9027f2, 32'hbee1efce} /* (14, 11, 25) {real, imag} */,
  {32'h3ed44e2f, 32'hbf0e26d8} /* (14, 11, 24) {real, imag} */,
  {32'h3eed133e, 32'hbee5aad3} /* (14, 11, 23) {real, imag} */,
  {32'hbc7fe100, 32'hbe22f092} /* (14, 11, 22) {real, imag} */,
  {32'h3eb30e8a, 32'h3f39a82d} /* (14, 11, 21) {real, imag} */,
  {32'hbe352ea2, 32'h3e171131} /* (14, 11, 20) {real, imag} */,
  {32'hbf018b8d, 32'h3e89ce17} /* (14, 11, 19) {real, imag} */,
  {32'h3dd86fe5, 32'hbc90166e} /* (14, 11, 18) {real, imag} */,
  {32'hbe3f3d1a, 32'h3d8ee391} /* (14, 11, 17) {real, imag} */,
  {32'hbefab361, 32'hbd40e98a} /* (14, 11, 16) {real, imag} */,
  {32'h3e84cf07, 32'h3d68e494} /* (14, 11, 15) {real, imag} */,
  {32'h3ef90ef0, 32'h3ee2ec17} /* (14, 11, 14) {real, imag} */,
  {32'h3eea0856, 32'hbd8f1dea} /* (14, 11, 13) {real, imag} */,
  {32'h3e703928, 32'hbddddc29} /* (14, 11, 12) {real, imag} */,
  {32'hbe5aef2a, 32'hbeed6f43} /* (14, 11, 11) {real, imag} */,
  {32'h3df9b8a2, 32'hbf3622c2} /* (14, 11, 10) {real, imag} */,
  {32'hbe2aeb46, 32'hbce00658} /* (14, 11, 9) {real, imag} */,
  {32'h3dc5fc20, 32'h3e1d54b8} /* (14, 11, 8) {real, imag} */,
  {32'h3ed775a8, 32'h3efafa1b} /* (14, 11, 7) {real, imag} */,
  {32'h3f02d79c, 32'h3edc5786} /* (14, 11, 6) {real, imag} */,
  {32'hbe1754a3, 32'h3e642ca6} /* (14, 11, 5) {real, imag} */,
  {32'h3d7baf97, 32'hbe904fba} /* (14, 11, 4) {real, imag} */,
  {32'hbe1daa61, 32'h3e8076b6} /* (14, 11, 3) {real, imag} */,
  {32'hbd945138, 32'h3ed5eb35} /* (14, 11, 2) {real, imag} */,
  {32'h3cab12da, 32'hbf7baf2a} /* (14, 11, 1) {real, imag} */,
  {32'hbf106db5, 32'hbf766e78} /* (14, 11, 0) {real, imag} */,
  {32'hbe12e34a, 32'h3e8f28c3} /* (14, 10, 31) {real, imag} */,
  {32'h3dd79e20, 32'hbf30250c} /* (14, 10, 30) {real, imag} */,
  {32'hbdae4d7a, 32'h3cb60260} /* (14, 10, 29) {real, imag} */,
  {32'hbf2a1715, 32'h3e1f50f4} /* (14, 10, 28) {real, imag} */,
  {32'hbe81bdd8, 32'hbe5d8994} /* (14, 10, 27) {real, imag} */,
  {32'h3f3985d9, 32'h3e1a9b70} /* (14, 10, 26) {real, imag} */,
  {32'h3f2ea7ae, 32'h3f42a69e} /* (14, 10, 25) {real, imag} */,
  {32'hbeaa9ed4, 32'h3e9acb56} /* (14, 10, 24) {real, imag} */,
  {32'h3e955a53, 32'h3f3c4af6} /* (14, 10, 23) {real, imag} */,
  {32'h3cf6f910, 32'h3dfcdb92} /* (14, 10, 22) {real, imag} */,
  {32'h3e0b2ac3, 32'hbee69055} /* (14, 10, 21) {real, imag} */,
  {32'hbb5116e0, 32'hbea2dc9c} /* (14, 10, 20) {real, imag} */,
  {32'hbe60b663, 32'h3da56ee2} /* (14, 10, 19) {real, imag} */,
  {32'h3e01dda2, 32'hbd81bd8e} /* (14, 10, 18) {real, imag} */,
  {32'h3e248a77, 32'hbf25e7c5} /* (14, 10, 17) {real, imag} */,
  {32'hbe82234b, 32'hbe990e8d} /* (14, 10, 16) {real, imag} */,
  {32'hbf0e4ea6, 32'h3ed1fe88} /* (14, 10, 15) {real, imag} */,
  {32'h3d663f28, 32'h3e38e038} /* (14, 10, 14) {real, imag} */,
  {32'hbde25868, 32'hbee45687} /* (14, 10, 13) {real, imag} */,
  {32'h3c6a5ca0, 32'h3eb39646} /* (14, 10, 12) {real, imag} */,
  {32'h3f148a6d, 32'hbd9fa698} /* (14, 10, 11) {real, imag} */,
  {32'h3da70212, 32'hbee86cb2} /* (14, 10, 10) {real, imag} */,
  {32'h3e02e1b3, 32'hbf04af94} /* (14, 10, 9) {real, imag} */,
  {32'hbd7b5fc8, 32'hbd3ef619} /* (14, 10, 8) {real, imag} */,
  {32'h3ea36ee6, 32'h3db3e555} /* (14, 10, 7) {real, imag} */,
  {32'h3e8955ea, 32'h3d7669ec} /* (14, 10, 6) {real, imag} */,
  {32'h3ef8faf0, 32'hbb217f00} /* (14, 10, 5) {real, imag} */,
  {32'hbd14d510, 32'hbf1810cc} /* (14, 10, 4) {real, imag} */,
  {32'hbe094436, 32'h3e197633} /* (14, 10, 3) {real, imag} */,
  {32'hbe389566, 32'hbd08d198} /* (14, 10, 2) {real, imag} */,
  {32'h3f670a46, 32'h3e0f2d3b} /* (14, 10, 1) {real, imag} */,
  {32'h3ea29090, 32'h3f4efe2b} /* (14, 10, 0) {real, imag} */,
  {32'hbe259db5, 32'h3f05d1b4} /* (14, 9, 31) {real, imag} */,
  {32'hbd97aa20, 32'hbeeeec56} /* (14, 9, 30) {real, imag} */,
  {32'h3e809193, 32'h3dea286f} /* (14, 9, 29) {real, imag} */,
  {32'h3ec414a9, 32'h3e5fa954} /* (14, 9, 28) {real, imag} */,
  {32'hbf261ebf, 32'hbeb8b3c8} /* (14, 9, 27) {real, imag} */,
  {32'h3e833108, 32'hbdc45c80} /* (14, 9, 26) {real, imag} */,
  {32'h3f4c817f, 32'h3e963ba8} /* (14, 9, 25) {real, imag} */,
  {32'h3e49773a, 32'hbe9ecf6c} /* (14, 9, 24) {real, imag} */,
  {32'hbe83d0fb, 32'hbdb8e3e4} /* (14, 9, 23) {real, imag} */,
  {32'hbeb91550, 32'h3e7a17ce} /* (14, 9, 22) {real, imag} */,
  {32'hbf361464, 32'h3ea6f738} /* (14, 9, 21) {real, imag} */,
  {32'hbdcf694a, 32'h3c5b8520} /* (14, 9, 20) {real, imag} */,
  {32'h3f115c1c, 32'hbede164f} /* (14, 9, 19) {real, imag} */,
  {32'h3f2a6e97, 32'hbf172b7f} /* (14, 9, 18) {real, imag} */,
  {32'hbea7d911, 32'hbe6a68e0} /* (14, 9, 17) {real, imag} */,
  {32'hbe1735ab, 32'h3dae30ec} /* (14, 9, 16) {real, imag} */,
  {32'hbd000f72, 32'hbf06e588} /* (14, 9, 15) {real, imag} */,
  {32'hbea31163, 32'h3cfc4b64} /* (14, 9, 14) {real, imag} */,
  {32'h3e4d795c, 32'hbe980da8} /* (14, 9, 13) {real, imag} */,
  {32'hbe941b13, 32'hbe41febe} /* (14, 9, 12) {real, imag} */,
  {32'hbe91e473, 32'h3ec988be} /* (14, 9, 11) {real, imag} */,
  {32'hbe00633b, 32'h3eefc54c} /* (14, 9, 10) {real, imag} */,
  {32'h3e5a1cc1, 32'hbd8b4bec} /* (14, 9, 9) {real, imag} */,
  {32'hbed8d8f3, 32'h3ec7ad17} /* (14, 9, 8) {real, imag} */,
  {32'hbf3582ae, 32'h3e91940a} /* (14, 9, 7) {real, imag} */,
  {32'hbe21a11a, 32'hbf1afbba} /* (14, 9, 6) {real, imag} */,
  {32'h3ebdc41b, 32'hbebab2c3} /* (14, 9, 5) {real, imag} */,
  {32'hbe3b1f17, 32'h3ec99d1d} /* (14, 9, 4) {real, imag} */,
  {32'hbe727797, 32'h3e9d50a5} /* (14, 9, 3) {real, imag} */,
  {32'h3e16cdaf, 32'hbe57fdf8} /* (14, 9, 2) {real, imag} */,
  {32'h3d1144c0, 32'hbd72ffb8} /* (14, 9, 1) {real, imag} */,
  {32'h3e6f8717, 32'h3e34ceba} /* (14, 9, 0) {real, imag} */,
  {32'hc00b4cde, 32'hbf9379d5} /* (14, 8, 31) {real, imag} */,
  {32'h3f2eaa56, 32'h3f198e3b} /* (14, 8, 30) {real, imag} */,
  {32'h3ebf9e15, 32'hbe6f409a} /* (14, 8, 29) {real, imag} */,
  {32'hbeb93fa0, 32'h3e9ca426} /* (14, 8, 28) {real, imag} */,
  {32'h3f404486, 32'hbd06343a} /* (14, 8, 27) {real, imag} */,
  {32'h3ee1e62d, 32'h3d27a084} /* (14, 8, 26) {real, imag} */,
  {32'h3ecd44c3, 32'h3e0da6a8} /* (14, 8, 25) {real, imag} */,
  {32'h3b8a84e8, 32'hbe4b9b90} /* (14, 8, 24) {real, imag} */,
  {32'hbdbe9ce8, 32'hbed26e8f} /* (14, 8, 23) {real, imag} */,
  {32'h3e30e129, 32'hbf11a2dc} /* (14, 8, 22) {real, imag} */,
  {32'h3ed0918c, 32'hbcc4b998} /* (14, 8, 21) {real, imag} */,
  {32'hbec012a8, 32'h3e33907d} /* (14, 8, 20) {real, imag} */,
  {32'h3dd579c4, 32'h3ea86238} /* (14, 8, 19) {real, imag} */,
  {32'h3cb1ff88, 32'hbd26cf1c} /* (14, 8, 18) {real, imag} */,
  {32'hbe06c192, 32'h3eaa9510} /* (14, 8, 17) {real, imag} */,
  {32'hbe5b26aa, 32'h3e53c248} /* (14, 8, 16) {real, imag} */,
  {32'hbe994266, 32'hbef160dd} /* (14, 8, 15) {real, imag} */,
  {32'h3e19a760, 32'h3e1b7eae} /* (14, 8, 14) {real, imag} */,
  {32'hbcac4510, 32'hbe3c17f3} /* (14, 8, 13) {real, imag} */,
  {32'hbeb784c2, 32'hbeb50657} /* (14, 8, 12) {real, imag} */,
  {32'h3f10ff78, 32'hbe6c41ea} /* (14, 8, 11) {real, imag} */,
  {32'hbf63d422, 32'h3e46dfd0} /* (14, 8, 10) {real, imag} */,
  {32'hbe4f55fd, 32'h3dc4726f} /* (14, 8, 9) {real, imag} */,
  {32'hbcadb8c0, 32'h3b8b3bc0} /* (14, 8, 8) {real, imag} */,
  {32'h3e88f3c7, 32'h3e46f734} /* (14, 8, 7) {real, imag} */,
  {32'h3d9923af, 32'h3d3254ec} /* (14, 8, 6) {real, imag} */,
  {32'hbd7f0ef6, 32'h3f488ef6} /* (14, 8, 5) {real, imag} */,
  {32'hbf4c9cd6, 32'h3d887159} /* (14, 8, 4) {real, imag} */,
  {32'hbe30765f, 32'h3e41c104} /* (14, 8, 3) {real, imag} */,
  {32'h3f365f51, 32'h3dee5a60} /* (14, 8, 2) {real, imag} */,
  {32'hbf2ea470, 32'hbf8a9226} /* (14, 8, 1) {real, imag} */,
  {32'hbf3a0d4e, 32'hbe64e9e6} /* (14, 8, 0) {real, imag} */,
  {32'h3f664b91, 32'hbf28ec68} /* (14, 7, 31) {real, imag} */,
  {32'hbe210d46, 32'hbf6a0730} /* (14, 7, 30) {real, imag} */,
  {32'h3df65ea0, 32'hbe00ace5} /* (14, 7, 29) {real, imag} */,
  {32'hbe8eef98, 32'hbea59c4d} /* (14, 7, 28) {real, imag} */,
  {32'hbf07d4d8, 32'h3f6bc854} /* (14, 7, 27) {real, imag} */,
  {32'hbf28b55b, 32'hbd7f4468} /* (14, 7, 26) {real, imag} */,
  {32'hbe9c5816, 32'h3e00fda0} /* (14, 7, 25) {real, imag} */,
  {32'hbcdffd68, 32'hbd5b750a} /* (14, 7, 24) {real, imag} */,
  {32'hbe8ee0e5, 32'h3e859fef} /* (14, 7, 23) {real, imag} */,
  {32'h3e884198, 32'h3dc70696} /* (14, 7, 22) {real, imag} */,
  {32'h3eacba39, 32'hbe3c2ff9} /* (14, 7, 21) {real, imag} */,
  {32'h3f369b24, 32'hbf5b02b9} /* (14, 7, 20) {real, imag} */,
  {32'h3eab7bc6, 32'h3e98d94d} /* (14, 7, 19) {real, imag} */,
  {32'hbe0fd3ed, 32'hbd71fa00} /* (14, 7, 18) {real, imag} */,
  {32'h3ea04da6, 32'hbd20e598} /* (14, 7, 17) {real, imag} */,
  {32'h3ea9d26c, 32'h3ee68c96} /* (14, 7, 16) {real, imag} */,
  {32'h3e83890f, 32'h3e25e198} /* (14, 7, 15) {real, imag} */,
  {32'hbe26c378, 32'h3c15b040} /* (14, 7, 14) {real, imag} */,
  {32'h3d4d5a2c, 32'h3f432e6d} /* (14, 7, 13) {real, imag} */,
  {32'hbf0a9490, 32'h3eff0658} /* (14, 7, 12) {real, imag} */,
  {32'hbe1670a6, 32'h3e05bc8b} /* (14, 7, 11) {real, imag} */,
  {32'hbd337cac, 32'h3f33a45c} /* (14, 7, 10) {real, imag} */,
  {32'hbea9c79b, 32'hbf1a7a14} /* (14, 7, 9) {real, imag} */,
  {32'h3e95c152, 32'hbf30954c} /* (14, 7, 8) {real, imag} */,
  {32'hbe6db2b6, 32'hbeda94f4} /* (14, 7, 7) {real, imag} */,
  {32'h3eabf63a, 32'hbeac81a8} /* (14, 7, 6) {real, imag} */,
  {32'hbe89f044, 32'hbe16c99a} /* (14, 7, 5) {real, imag} */,
  {32'hbf6e6cac, 32'h3f04a701} /* (14, 7, 4) {real, imag} */,
  {32'hbe08a118, 32'hbe7f7a2c} /* (14, 7, 3) {real, imag} */,
  {32'h3e156b2c, 32'hbf1833ce} /* (14, 7, 2) {real, imag} */,
  {32'hbe751c4e, 32'h3f636c2e} /* (14, 7, 1) {real, imag} */,
  {32'hbd71350c, 32'h3f9d80aa} /* (14, 7, 0) {real, imag} */,
  {32'h3eac37d9, 32'h3e93cbb8} /* (14, 6, 31) {real, imag} */,
  {32'h3f493076, 32'h3e254934} /* (14, 6, 30) {real, imag} */,
  {32'hbf8a773c, 32'hbf070b6e} /* (14, 6, 29) {real, imag} */,
  {32'hbeccac08, 32'hbe83f7fe} /* (14, 6, 28) {real, imag} */,
  {32'hbe94de72, 32'h3e5e7216} /* (14, 6, 27) {real, imag} */,
  {32'h3e5abdea, 32'h3f3663df} /* (14, 6, 26) {real, imag} */,
  {32'hbf293a68, 32'hbf7e66ad} /* (14, 6, 25) {real, imag} */,
  {32'hbd877de8, 32'h3e8768ad} /* (14, 6, 24) {real, imag} */,
  {32'h3e6789e5, 32'h3f103725} /* (14, 6, 23) {real, imag} */,
  {32'hbe293bda, 32'hbf09bc72} /* (14, 6, 22) {real, imag} */,
  {32'hbe08f2e9, 32'h3e9cdd25} /* (14, 6, 21) {real, imag} */,
  {32'hbd58aac8, 32'h3f1249e2} /* (14, 6, 20) {real, imag} */,
  {32'h3e577f42, 32'hbed26a7a} /* (14, 6, 19) {real, imag} */,
  {32'h3d9cf1fa, 32'hbe998f25} /* (14, 6, 18) {real, imag} */,
  {32'hbdaf6a21, 32'hbefe59a8} /* (14, 6, 17) {real, imag} */,
  {32'hbbcb79b8, 32'hbce26804} /* (14, 6, 16) {real, imag} */,
  {32'h3e87bd8f, 32'h3dae5980} /* (14, 6, 15) {real, imag} */,
  {32'hbedfa61c, 32'h3c2e2298} /* (14, 6, 14) {real, imag} */,
  {32'h3da955b4, 32'hbd87b2a4} /* (14, 6, 13) {real, imag} */,
  {32'h3e773050, 32'hbe4a2770} /* (14, 6, 12) {real, imag} */,
  {32'h3ed0c398, 32'hbe8f4176} /* (14, 6, 11) {real, imag} */,
  {32'h3f11b883, 32'h3d7ffbc2} /* (14, 6, 10) {real, imag} */,
  {32'hbeaabd29, 32'h3e80f859} /* (14, 6, 9) {real, imag} */,
  {32'h3e5c6480, 32'h3e9f0860} /* (14, 6, 8) {real, imag} */,
  {32'hbd15af88, 32'hbea3e626} /* (14, 6, 7) {real, imag} */,
  {32'hbecdae02, 32'h3e070fd2} /* (14, 6, 6) {real, imag} */,
  {32'h3cc130a8, 32'hbf268dfc} /* (14, 6, 5) {real, imag} */,
  {32'hbea4bb72, 32'h3e41714b} /* (14, 6, 4) {real, imag} */,
  {32'h3e103f6c, 32'h3f1dd5dc} /* (14, 6, 3) {real, imag} */,
  {32'h3f64a15d, 32'h3e87f3d8} /* (14, 6, 2) {real, imag} */,
  {32'hbee50a4d, 32'hbb9fa320} /* (14, 6, 1) {real, imag} */,
  {32'hbeb24388, 32'h3df0aaa4} /* (14, 6, 0) {real, imag} */,
  {32'hc00a8fb9, 32'h3f906b62} /* (14, 5, 31) {real, imag} */,
  {32'h3e3f196c, 32'h3e99df2d} /* (14, 5, 30) {real, imag} */,
  {32'hbe9bf32b, 32'h3f213c4d} /* (14, 5, 29) {real, imag} */,
  {32'hbe83166e, 32'hbe101be0} /* (14, 5, 28) {real, imag} */,
  {32'h3f212148, 32'hbe857d60} /* (14, 5, 27) {real, imag} */,
  {32'hbe85c78e, 32'h3e395292} /* (14, 5, 26) {real, imag} */,
  {32'hbe17b01e, 32'h3e83c661} /* (14, 5, 25) {real, imag} */,
  {32'h3e0be2f0, 32'h3d0f8218} /* (14, 5, 24) {real, imag} */,
  {32'h3daf7814, 32'hbd4058d5} /* (14, 5, 23) {real, imag} */,
  {32'hbbdedee0, 32'hbd73fd54} /* (14, 5, 22) {real, imag} */,
  {32'h3e8b0d2c, 32'hbcaa6d28} /* (14, 5, 21) {real, imag} */,
  {32'hbe2c88ba, 32'hbd5e12dc} /* (14, 5, 20) {real, imag} */,
  {32'hbc5a2e8a, 32'h3dc2ad0c} /* (14, 5, 19) {real, imag} */,
  {32'h3e974fbe, 32'hbe6312c4} /* (14, 5, 18) {real, imag} */,
  {32'h3e1313db, 32'h3db6a100} /* (14, 5, 17) {real, imag} */,
  {32'hbd53ad4e, 32'hbe08e3d4} /* (14, 5, 16) {real, imag} */,
  {32'h3e5b2fab, 32'hbd5b4002} /* (14, 5, 15) {real, imag} */,
  {32'h3bb56860, 32'h3efcd092} /* (14, 5, 14) {real, imag} */,
  {32'h3ebf3c45, 32'hbe17a45a} /* (14, 5, 13) {real, imag} */,
  {32'hbea1158d, 32'h3e037c86} /* (14, 5, 12) {real, imag} */,
  {32'hbd016d0e, 32'hbce85bc0} /* (14, 5, 11) {real, imag} */,
  {32'h3d725186, 32'h3ef725a7} /* (14, 5, 10) {real, imag} */,
  {32'h3d87d2b4, 32'hbd8eb2d8} /* (14, 5, 9) {real, imag} */,
  {32'hbeebae52, 32'h3ec67e9e} /* (14, 5, 8) {real, imag} */,
  {32'hbe59279e, 32'h3c641dd8} /* (14, 5, 7) {real, imag} */,
  {32'h3ec5672d, 32'hbc915b80} /* (14, 5, 6) {real, imag} */,
  {32'h3eda6178, 32'h3f2e6b49} /* (14, 5, 5) {real, imag} */,
  {32'h3e72bc27, 32'hbef0e036} /* (14, 5, 4) {real, imag} */,
  {32'hbddc9e28, 32'h3d8d9280} /* (14, 5, 3) {real, imag} */,
  {32'hbb06c500, 32'h3ede278c} /* (14, 5, 2) {real, imag} */,
  {32'hc04d3d71, 32'hbf248e40} /* (14, 5, 1) {real, imag} */,
  {32'hc002f9fd, 32'hbfa03f75} /* (14, 5, 0) {real, imag} */,
  {32'h400f529d, 32'h3f5443c0} /* (14, 4, 31) {real, imag} */,
  {32'hbfcf7cae, 32'hc01f0bce} /* (14, 4, 30) {real, imag} */,
  {32'hbefd9df8, 32'hbe927616} /* (14, 4, 29) {real, imag} */,
  {32'h3f528d42, 32'h3fb1772c} /* (14, 4, 28) {real, imag} */,
  {32'hbf144570, 32'h3f3fcf1e} /* (14, 4, 27) {real, imag} */,
  {32'hbdcecff4, 32'h3ee4c278} /* (14, 4, 26) {real, imag} */,
  {32'hbe7e5b74, 32'h3f8cc61a} /* (14, 4, 25) {real, imag} */,
  {32'hbec1fbbe, 32'h3e7e98f2} /* (14, 4, 24) {real, imag} */,
  {32'hbdaf57e4, 32'hbe942478} /* (14, 4, 23) {real, imag} */,
  {32'hbe3a6203, 32'h3dd15d70} /* (14, 4, 22) {real, imag} */,
  {32'hbe796f88, 32'h3dfa4d25} /* (14, 4, 21) {real, imag} */,
  {32'h3d417eec, 32'h3de6af62} /* (14, 4, 20) {real, imag} */,
  {32'hbede1de1, 32'hbf07f8f1} /* (14, 4, 19) {real, imag} */,
  {32'hbe4ca6f4, 32'h3dd820bd} /* (14, 4, 18) {real, imag} */,
  {32'hbe9c6e6b, 32'h3e951f59} /* (14, 4, 17) {real, imag} */,
  {32'h3dd3392a, 32'hbc219e58} /* (14, 4, 16) {real, imag} */,
  {32'hbd5a3196, 32'hbeeed944} /* (14, 4, 15) {real, imag} */,
  {32'hbe2ec4c5, 32'hbef42284} /* (14, 4, 14) {real, imag} */,
  {32'hbe4545e5, 32'h3e1355fe} /* (14, 4, 13) {real, imag} */,
  {32'h3ce7cb54, 32'hbddc865c} /* (14, 4, 12) {real, imag} */,
  {32'hbe723ae4, 32'hbde38603} /* (14, 4, 11) {real, imag} */,
  {32'h3e9ff1de, 32'h3f2cefd6} /* (14, 4, 10) {real, imag} */,
  {32'h3f95c679, 32'hbe5725db} /* (14, 4, 9) {real, imag} */,
  {32'hbe0b8abd, 32'h3e76d71a} /* (14, 4, 8) {real, imag} */,
  {32'hbe22d18d, 32'h3dd598ec} /* (14, 4, 7) {real, imag} */,
  {32'hbf245d95, 32'h3f15fbc3} /* (14, 4, 6) {real, imag} */,
  {32'hbf204ab9, 32'hbed4b97a} /* (14, 4, 5) {real, imag} */,
  {32'h3efd4c94, 32'h3f6268e5} /* (14, 4, 4) {real, imag} */,
  {32'hbecc4708, 32'h3f36cea1} /* (14, 4, 3) {real, imag} */,
  {32'hbffd71c0, 32'hc000cfd4} /* (14, 4, 2) {real, imag} */,
  {32'h40a1860a, 32'h3f5fed02} /* (14, 4, 1) {real, imag} */,
  {32'hbdd038b8, 32'hbf363da8} /* (14, 4, 0) {real, imag} */,
  {32'hc0204d1c, 32'h3fb015a3} /* (14, 3, 31) {real, imag} */,
  {32'h400c3096, 32'hbfd49870} /* (14, 3, 30) {real, imag} */,
  {32'hbe9d9938, 32'h3f794558} /* (14, 3, 29) {real, imag} */,
  {32'h3f4bba10, 32'h3f0aeab8} /* (14, 3, 28) {real, imag} */,
  {32'hbf181f2e, 32'hbe848d60} /* (14, 3, 27) {real, imag} */,
  {32'hbe8bb090, 32'hbdd29ec8} /* (14, 3, 26) {real, imag} */,
  {32'hbde11cb9, 32'hbe719618} /* (14, 3, 25) {real, imag} */,
  {32'hbebdad1d, 32'hbe8d8afe} /* (14, 3, 24) {real, imag} */,
  {32'hbf259772, 32'hbe695803} /* (14, 3, 23) {real, imag} */,
  {32'hbe9849e9, 32'h3f3f51fd} /* (14, 3, 22) {real, imag} */,
  {32'hbeb6a7db, 32'hbebb18dc} /* (14, 3, 21) {real, imag} */,
  {32'h3e9a6fe2, 32'h3eba8d5e} /* (14, 3, 20) {real, imag} */,
  {32'h3eac1c13, 32'hbe1b2ac4} /* (14, 3, 19) {real, imag} */,
  {32'hbd762d7f, 32'hbe2ea436} /* (14, 3, 18) {real, imag} */,
  {32'hbdc96dfb, 32'h3d26038c} /* (14, 3, 17) {real, imag} */,
  {32'hbe050566, 32'h3d4aaae0} /* (14, 3, 16) {real, imag} */,
  {32'hbe56e812, 32'h3e8848bc} /* (14, 3, 15) {real, imag} */,
  {32'h3e9e6c95, 32'h3dd18254} /* (14, 3, 14) {real, imag} */,
  {32'hbd039296, 32'hbd641104} /* (14, 3, 13) {real, imag} */,
  {32'h3da80470, 32'h3da5163c} /* (14, 3, 12) {real, imag} */,
  {32'h3ebf6950, 32'h3f0759ef} /* (14, 3, 11) {real, imag} */,
  {32'hbd9a3350, 32'h3e1a661c} /* (14, 3, 10) {real, imag} */,
  {32'hbe5f326e, 32'hbf6ef5bc} /* (14, 3, 9) {real, imag} */,
  {32'h3ebe50a5, 32'h3cc78ec0} /* (14, 3, 8) {real, imag} */,
  {32'h3f45b8bc, 32'hbe43492c} /* (14, 3, 7) {real, imag} */,
  {32'h3c9e43c0, 32'hbe274f0c} /* (14, 3, 6) {real, imag} */,
  {32'h3e2551f8, 32'h3f8a92a0} /* (14, 3, 5) {real, imag} */,
  {32'hbe744766, 32'h3f22b238} /* (14, 3, 4) {real, imag} */,
  {32'h3f10bc2d, 32'h3ec550dc} /* (14, 3, 3) {real, imag} */,
  {32'hbf57d97b, 32'hbffeee7a} /* (14, 3, 2) {real, imag} */,
  {32'h405aa10d, 32'h400aa287} /* (14, 3, 1) {real, imag} */,
  {32'h3f23d1be, 32'h3e522f1e} /* (14, 3, 0) {real, imag} */,
  {32'hc1c04433, 32'hc0000be0} /* (14, 2, 31) {real, imag} */,
  {32'h414a1049, 32'hc09496c6} /* (14, 2, 30) {real, imag} */,
  {32'h3eb84045, 32'h3ed4297a} /* (14, 2, 29) {real, imag} */,
  {32'hbfcfb7b5, 32'h40296ac6} /* (14, 2, 28) {real, imag} */,
  {32'h3fbbefd2, 32'hbefe4132} /* (14, 2, 27) {real, imag} */,
  {32'h3ddfc6a8, 32'hbf390066} /* (14, 2, 26) {real, imag} */,
  {32'hbf4cc744, 32'h3e95f5cf} /* (14, 2, 25) {real, imag} */,
  {32'h3e1c9cd3, 32'hbee373d8} /* (14, 2, 24) {real, imag} */,
  {32'h3db2944b, 32'hbedeecb2} /* (14, 2, 23) {real, imag} */,
  {32'h3e2e2cb8, 32'h3ef7ca5b} /* (14, 2, 22) {real, imag} */,
  {32'h3debe5cd, 32'hbe0c533c} /* (14, 2, 21) {real, imag} */,
  {32'h3e626fd6, 32'hbeb8df83} /* (14, 2, 20) {real, imag} */,
  {32'hbe9fbfbf, 32'h3ea6809e} /* (14, 2, 19) {real, imag} */,
  {32'h3e492458, 32'hbf103a1c} /* (14, 2, 18) {real, imag} */,
  {32'h3e798700, 32'h3f04d02c} /* (14, 2, 17) {real, imag} */,
  {32'h3d5507f8, 32'hbe323628} /* (14, 2, 16) {real, imag} */,
  {32'hbce46878, 32'h3d6e0fb6} /* (14, 2, 15) {real, imag} */,
  {32'h3f3ce754, 32'h3dd52982} /* (14, 2, 14) {real, imag} */,
  {32'hbf130e4a, 32'h3ea8162b} /* (14, 2, 13) {real, imag} */,
  {32'hbd71e780, 32'hbe95bf64} /* (14, 2, 12) {real, imag} */,
  {32'h3e7ab9d2, 32'h3f01fa44} /* (14, 2, 11) {real, imag} */,
  {32'hbcf19170, 32'h3df8a7ac} /* (14, 2, 10) {real, imag} */,
  {32'h3d0ca328, 32'h3ec5aa72} /* (14, 2, 9) {real, imag} */,
  {32'h3fc0d158, 32'h3eee1d02} /* (14, 2, 8) {real, imag} */,
  {32'hbcb66040, 32'h3e1e00c3} /* (14, 2, 7) {real, imag} */,
  {32'hbecbac48, 32'h3f9a9d6f} /* (14, 2, 6) {real, imag} */,
  {32'h3fd387d8, 32'h401dad09} /* (14, 2, 5) {real, imag} */,
  {32'hbfba6fd8, 32'hbff90b6e} /* (14, 2, 4) {real, imag} */,
  {32'h3e3e1bd8, 32'h3e26f602} /* (14, 2, 3) {real, imag} */,
  {32'h40fef71b, 32'hbf5b8362} /* (14, 2, 2) {real, imag} */,
  {32'hc15ce4b0, 32'h3f9bfa32} /* (14, 2, 1) {real, imag} */,
  {32'hc14edef5, 32'hbff91f82} /* (14, 2, 0) {real, imag} */,
  {32'h41f54011, 32'hc1019160} /* (14, 1, 31) {real, imag} */,
  {32'hc10f225e, 32'hbf0fbbcb} /* (14, 1, 30) {real, imag} */,
  {32'h3de25e82, 32'h3ff86364} /* (14, 1, 29) {real, imag} */,
  {32'h400bda14, 32'hbe32bcd8} /* (14, 1, 28) {real, imag} */,
  {32'hc021f3d4, 32'h3f173340} /* (14, 1, 27) {real, imag} */,
  {32'h3f3c57f6, 32'hbe36ba80} /* (14, 1, 26) {real, imag} */,
  {32'h3b342880, 32'h3f6734e8} /* (14, 1, 25) {real, imag} */,
  {32'hbf8962fe, 32'h3d8a0b3c} /* (14, 1, 24) {real, imag} */,
  {32'hbebd07ec, 32'hbddcc148} /* (14, 1, 23) {real, imag} */,
  {32'h3e8330a7, 32'hbdcfd346} /* (14, 1, 22) {real, imag} */,
  {32'hbeeb1256, 32'h3f7b4b94} /* (14, 1, 21) {real, imag} */,
  {32'hbe0537a0, 32'hbe0bb386} /* (14, 1, 20) {real, imag} */,
  {32'hbd548f88, 32'hbe0c41e0} /* (14, 1, 19) {real, imag} */,
  {32'hbd614204, 32'h3ea444f4} /* (14, 1, 18) {real, imag} */,
  {32'hbdea6e9e, 32'h3e6b499e} /* (14, 1, 17) {real, imag} */,
  {32'h3e4fc513, 32'hbe05c5da} /* (14, 1, 16) {real, imag} */,
  {32'hbe37a2e6, 32'h3e169be0} /* (14, 1, 15) {real, imag} */,
  {32'hbd90b127, 32'hbef1a5a8} /* (14, 1, 14) {real, imag} */,
  {32'h3f25bc2e, 32'h3b26aab0} /* (14, 1, 13) {real, imag} */,
  {32'h3e66d3df, 32'hbe4ee9a6} /* (14, 1, 12) {real, imag} */,
  {32'h3c49ea30, 32'hbf1c8435} /* (14, 1, 11) {real, imag} */,
  {32'hbd8ad7d8, 32'hbe91c863} /* (14, 1, 10) {real, imag} */,
  {32'hbd7adf00, 32'h3e706a1c} /* (14, 1, 9) {real, imag} */,
  {32'hbf0d17b2, 32'hbecc599e} /* (14, 1, 8) {real, imag} */,
  {32'h3f3ba0cb, 32'h3f75aa6e} /* (14, 1, 7) {real, imag} */,
  {32'h3dc62b18, 32'hbfc28469} /* (14, 1, 6) {real, imag} */,
  {32'hbf8e2118, 32'hbf7e0fc7} /* (14, 1, 5) {real, imag} */,
  {32'hbf81c90a, 32'h400b4e7f} /* (14, 1, 4) {real, imag} */,
  {32'hc05292c6, 32'hbeb46ae2} /* (14, 1, 3) {real, imag} */,
  {32'hc144f800, 32'hc12c851c} /* (14, 1, 2) {real, imag} */,
  {32'h421b9faf, 32'h41c42c5e} /* (14, 1, 1) {real, imag} */,
  {32'h420aa966, 32'hbeffab80} /* (14, 1, 0) {real, imag} */,
  {32'h41a1fa34, 32'hc18d8503} /* (14, 0, 31) {real, imag} */,
  {32'hc073e1ad, 32'h40ce8f90} /* (14, 0, 30) {real, imag} */,
  {32'h3ea8c798, 32'h3e0f08a0} /* (14, 0, 29) {real, imag} */,
  {32'hbf0721a9, 32'h3edd747f} /* (14, 0, 28) {real, imag} */,
  {32'hbff36b84, 32'h3ec1dbec} /* (14, 0, 27) {real, imag} */,
  {32'h3c620210, 32'hbe7c444c} /* (14, 0, 26) {real, imag} */,
  {32'hbe95e2c2, 32'hbe752606} /* (14, 0, 25) {real, imag} */,
  {32'h3f289dfb, 32'h3f0819f4} /* (14, 0, 24) {real, imag} */,
  {32'hbee6cc03, 32'h3e588449} /* (14, 0, 23) {real, imag} */,
  {32'hbef44116, 32'hbf4f10b5} /* (14, 0, 22) {real, imag} */,
  {32'hbee1921f, 32'h3c409550} /* (14, 0, 21) {real, imag} */,
  {32'h3f0c5a07, 32'h3eabcc18} /* (14, 0, 20) {real, imag} */,
  {32'h3c92ab38, 32'hbe37d640} /* (14, 0, 19) {real, imag} */,
  {32'hbee08057, 32'h3ea2d0d7} /* (14, 0, 18) {real, imag} */,
  {32'hbde81d9e, 32'h3e9bcf86} /* (14, 0, 17) {real, imag} */,
  {32'h3df6c459, 32'h00000000} /* (14, 0, 16) {real, imag} */,
  {32'hbde81d9e, 32'hbe9bcf86} /* (14, 0, 15) {real, imag} */,
  {32'hbee08057, 32'hbea2d0d7} /* (14, 0, 14) {real, imag} */,
  {32'h3c92ab38, 32'h3e37d640} /* (14, 0, 13) {real, imag} */,
  {32'h3f0c5a07, 32'hbeabcc18} /* (14, 0, 12) {real, imag} */,
  {32'hbee1921f, 32'hbc409550} /* (14, 0, 11) {real, imag} */,
  {32'hbef44116, 32'h3f4f10b5} /* (14, 0, 10) {real, imag} */,
  {32'hbee6cc03, 32'hbe588449} /* (14, 0, 9) {real, imag} */,
  {32'h3f289dfb, 32'hbf0819f4} /* (14, 0, 8) {real, imag} */,
  {32'hbe95e2c2, 32'h3e752606} /* (14, 0, 7) {real, imag} */,
  {32'h3c620210, 32'h3e7c444c} /* (14, 0, 6) {real, imag} */,
  {32'hbff36b84, 32'hbec1dbec} /* (14, 0, 5) {real, imag} */,
  {32'hbf0721a9, 32'hbedd747f} /* (14, 0, 4) {real, imag} */,
  {32'h3ea8c798, 32'hbe0f08a0} /* (14, 0, 3) {real, imag} */,
  {32'hc073e1ad, 32'hc0ce8f90} /* (14, 0, 2) {real, imag} */,
  {32'h41a1fa34, 32'h418d8503} /* (14, 0, 1) {real, imag} */,
  {32'h420f1b02, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h4261b185, 32'hc2086478} /* (13, 31, 31) {real, imag} */,
  {32'hc182e8c4, 32'h416c369e} /* (13, 31, 30) {real, imag} */,
  {32'hc034c27d, 32'h3e5ada78} /* (13, 31, 29) {real, imag} */,
  {32'hbf2e13db, 32'hc023767e} /* (13, 31, 28) {real, imag} */,
  {32'hbfdabc92, 32'h3f27d83a} /* (13, 31, 27) {real, imag} */,
  {32'hbea6abd0, 32'h3fbc441e} /* (13, 31, 26) {real, imag} */,
  {32'h3f84747f, 32'hbe6777a5} /* (13, 31, 25) {real, imag} */,
  {32'hbe787749, 32'h3fba3654} /* (13, 31, 24) {real, imag} */,
  {32'h3dacbf30, 32'hbe23a6f9} /* (13, 31, 23) {real, imag} */,
  {32'h3e55f99e, 32'h3e5461a2} /* (13, 31, 22) {real, imag} */,
  {32'hbee84b84, 32'hbe587810} /* (13, 31, 21) {real, imag} */,
  {32'h3f032e1e, 32'h3da09c45} /* (13, 31, 20) {real, imag} */,
  {32'hbd891a82, 32'h3e127560} /* (13, 31, 19) {real, imag} */,
  {32'h3e5aa498, 32'hbec2f752} /* (13, 31, 18) {real, imag} */,
  {32'hbe15677c, 32'h3e504219} /* (13, 31, 17) {real, imag} */,
  {32'h3d1e4d7a, 32'hbdeb9c43} /* (13, 31, 16) {real, imag} */,
  {32'hbe6b603b, 32'h3eb797e4} /* (13, 31, 15) {real, imag} */,
  {32'hbcf6c148, 32'hbe9373e6} /* (13, 31, 14) {real, imag} */,
  {32'h3dba2386, 32'h3e880944} /* (13, 31, 13) {real, imag} */,
  {32'hbe4962ea, 32'h3e16c8ee} /* (13, 31, 12) {real, imag} */,
  {32'h3e77833e, 32'hbf5130c4} /* (13, 31, 11) {real, imag} */,
  {32'h3ed6a2ef, 32'hbee7e2aa} /* (13, 31, 10) {real, imag} */,
  {32'hbf665271, 32'hbe9d0d82} /* (13, 31, 9) {real, imag} */,
  {32'hbf45ff5d, 32'hbf673836} /* (13, 31, 8) {real, imag} */,
  {32'h3e4f47b6, 32'hbe0a0662} /* (13, 31, 7) {real, imag} */,
  {32'h3f715cf4, 32'hbcf31240} /* (13, 31, 6) {real, imag} */,
  {32'hc050536d, 32'hbf139335} /* (13, 31, 5) {real, imag} */,
  {32'h400aae68, 32'hbf0e8612} /* (13, 31, 4) {real, imag} */,
  {32'h3dfb94b8, 32'hbfc90d33} /* (13, 31, 3) {real, imag} */,
  {32'hc13454ff, 32'h3b5bd280} /* (13, 31, 2) {real, imag} */,
  {32'h422a3b02, 32'h411bc8b7} /* (13, 31, 1) {real, imag} */,
  {32'h4250d69a, 32'hc009118f} /* (13, 31, 0) {real, imag} */,
  {32'hc19114de, 32'hc0028f76} /* (13, 30, 31) {real, imag} */,
  {32'h411f13b5, 32'h40325670} /* (13, 30, 30) {real, imag} */,
  {32'h3eb0d0ee, 32'hbe976950} /* (13, 30, 29) {real, imag} */,
  {32'hc0294460, 32'h4000e95a} /* (13, 30, 28) {real, imag} */,
  {32'h3fad1202, 32'hc012c31d} /* (13, 30, 27) {real, imag} */,
  {32'h3e42dbcf, 32'hbf20b9a9} /* (13, 30, 26) {real, imag} */,
  {32'hbf04c831, 32'h3ec8bc52} /* (13, 30, 25) {real, imag} */,
  {32'h3f320941, 32'h3e489240} /* (13, 30, 24) {real, imag} */,
  {32'hbea9a519, 32'h3e9a11d5} /* (13, 30, 23) {real, imag} */,
  {32'hbdf3e737, 32'hbdaed053} /* (13, 30, 22) {real, imag} */,
  {32'h3d8a8dfa, 32'hbe8e0133} /* (13, 30, 21) {real, imag} */,
  {32'h3ec4da32, 32'h3d19dd4a} /* (13, 30, 20) {real, imag} */,
  {32'hbdc41c38, 32'h3d727df8} /* (13, 30, 19) {real, imag} */,
  {32'h3e06d73e, 32'h3cc77020} /* (13, 30, 18) {real, imag} */,
  {32'hbdfa6fe6, 32'hbd80c659} /* (13, 30, 17) {real, imag} */,
  {32'h3dc048ba, 32'h3e89ff00} /* (13, 30, 16) {real, imag} */,
  {32'h3e271e94, 32'h3df1e27c} /* (13, 30, 15) {real, imag} */,
  {32'h3e52eaa6, 32'h3e39d64a} /* (13, 30, 14) {real, imag} */,
  {32'hbebd2edf, 32'hbebdddff} /* (13, 30, 13) {real, imag} */,
  {32'hbe88a3c5, 32'h3d023a6c} /* (13, 30, 12) {real, imag} */,
  {32'h3f45c5b7, 32'h3f165722} /* (13, 30, 11) {real, imag} */,
  {32'h3d7be8a6, 32'hbe451894} /* (13, 30, 10) {real, imag} */,
  {32'hbf2a734e, 32'hbd9195c8} /* (13, 30, 9) {real, imag} */,
  {32'h3f0a2f20, 32'h3f9cc432} /* (13, 30, 8) {real, imag} */,
  {32'hbf3f6962, 32'hbea68bfe} /* (13, 30, 7) {real, imag} */,
  {32'h3f71b084, 32'h3f164333} /* (13, 30, 6) {real, imag} */,
  {32'h3fd2dfd8, 32'h3faeb7d0} /* (13, 30, 5) {real, imag} */,
  {32'hbffc727d, 32'hc01aa5a0} /* (13, 30, 4) {real, imag} */,
  {32'h3f0ee477, 32'hbfb6c940} /* (13, 30, 3) {real, imag} */,
  {32'h4180fd8c, 32'h40bc423d} /* (13, 30, 2) {real, imag} */,
  {32'hc2015e68, 32'h3f818fb5} /* (13, 30, 1) {real, imag} */,
  {32'hc180e086, 32'h4001dfa2} /* (13, 30, 0) {real, imag} */,
  {32'h409fb372, 32'hc03e16a3} /* (13, 29, 31) {real, imag} */,
  {32'hbf7e4c2e, 32'h400f0f16} /* (13, 29, 30) {real, imag} */,
  {32'h3d881768, 32'hbee725fc} /* (13, 29, 29) {real, imag} */,
  {32'hbe71406c, 32'hbe9adfc1} /* (13, 29, 28) {real, imag} */,
  {32'h3e12de62, 32'hbf815ec2} /* (13, 29, 27) {real, imag} */,
  {32'h3e1ada3e, 32'h3e5748a0} /* (13, 29, 26) {real, imag} */,
  {32'h3f073f7e, 32'hbe545d4e} /* (13, 29, 25) {real, imag} */,
  {32'h3ed44653, 32'h3e632b28} /* (13, 29, 24) {real, imag} */,
  {32'hbf2665ad, 32'h3f45a785} /* (13, 29, 23) {real, imag} */,
  {32'hbeb55213, 32'hbe48641c} /* (13, 29, 22) {real, imag} */,
  {32'h3f1c4002, 32'h3e2ebbca} /* (13, 29, 21) {real, imag} */,
  {32'h3e8734c1, 32'h3ebae193} /* (13, 29, 20) {real, imag} */,
  {32'hbd628a90, 32'hbe5394ce} /* (13, 29, 19) {real, imag} */,
  {32'hbe940fbd, 32'hbe5fb95f} /* (13, 29, 18) {real, imag} */,
  {32'h3e862dcb, 32'h3ef59eb1} /* (13, 29, 17) {real, imag} */,
  {32'h3e0c217f, 32'h3d97d838} /* (13, 29, 16) {real, imag} */,
  {32'hbe1b4100, 32'hbeb06c75} /* (13, 29, 15) {real, imag} */,
  {32'hbdd19008, 32'hbe79caa6} /* (13, 29, 14) {real, imag} */,
  {32'hbe176c15, 32'h3ea2b43e} /* (13, 29, 13) {real, imag} */,
  {32'hbe8bb8bf, 32'h3ec4d7fd} /* (13, 29, 12) {real, imag} */,
  {32'hbe2ea28d, 32'h3e353435} /* (13, 29, 11) {real, imag} */,
  {32'h3dd4200c, 32'hbf1f8cf4} /* (13, 29, 10) {real, imag} */,
  {32'h3ae40c80, 32'hbe68fc8d} /* (13, 29, 9) {real, imag} */,
  {32'h3e92f958, 32'h3f1f822c} /* (13, 29, 8) {real, imag} */,
  {32'h3ef954ec, 32'hbe845988} /* (13, 29, 7) {real, imag} */,
  {32'hbf5ef5ef, 32'hbc8bc6b0} /* (13, 29, 6) {real, imag} */,
  {32'hbe966041, 32'hbe8d634d} /* (13, 29, 5) {real, imag} */,
  {32'h3f819c62, 32'hbf610618} /* (13, 29, 4) {real, imag} */,
  {32'hbec42026, 32'hbf2e3352} /* (13, 29, 3) {real, imag} */,
  {32'h4031e709, 32'h401ad8bc} /* (13, 29, 2) {real, imag} */,
  {32'hc0a3e835, 32'hbfb61e82} /* (13, 29, 1) {real, imag} */,
  {32'h3d2660e0, 32'h3eeacc22} /* (13, 29, 0) {real, imag} */,
  {32'h40c134bb, 32'hbf23fbe6} /* (13, 28, 31) {real, imag} */,
  {32'hbff38a88, 32'h4014fddf} /* (13, 28, 30) {real, imag} */,
  {32'hbebd5dd2, 32'hbf466230} /* (13, 28, 29) {real, imag} */,
  {32'hbe95f132, 32'hbf150263} /* (13, 28, 28) {real, imag} */,
  {32'hbe95d4a8, 32'h3f92b3a1} /* (13, 28, 27) {real, imag} */,
  {32'hbeb4e8dc, 32'hbe95d063} /* (13, 28, 26) {real, imag} */,
  {32'hbeb8111a, 32'h3e6f40a5} /* (13, 28, 25) {real, imag} */,
  {32'h3c08b118, 32'h3f2796ce} /* (13, 28, 24) {real, imag} */,
  {32'h3eabf314, 32'hbc1fd3e0} /* (13, 28, 23) {real, imag} */,
  {32'hbef2e426, 32'hbd537064} /* (13, 28, 22) {real, imag} */,
  {32'h3ee72d82, 32'hbddc4be5} /* (13, 28, 21) {real, imag} */,
  {32'hbdbc8419, 32'hbeb5cf08} /* (13, 28, 20) {real, imag} */,
  {32'h3e8f1810, 32'h3e982688} /* (13, 28, 19) {real, imag} */,
  {32'hbd732c70, 32'h3ecbbd1f} /* (13, 28, 18) {real, imag} */,
  {32'h3e5e528c, 32'h3d861a46} /* (13, 28, 17) {real, imag} */,
  {32'h3d5ec480, 32'hbe3f1d7d} /* (13, 28, 16) {real, imag} */,
  {32'h3e97c6a2, 32'h3ca10444} /* (13, 28, 15) {real, imag} */,
  {32'h3e2b6e14, 32'hbeeace81} /* (13, 28, 14) {real, imag} */,
  {32'h3ebc092b, 32'h3ecbc68e} /* (13, 28, 13) {real, imag} */,
  {32'hbed910d7, 32'h3ed22389} /* (13, 28, 12) {real, imag} */,
  {32'hbee2338a, 32'hbe964ae7} /* (13, 28, 11) {real, imag} */,
  {32'h3e275a64, 32'h3b933c00} /* (13, 28, 10) {real, imag} */,
  {32'h3e0589ea, 32'h3f0d8598} /* (13, 28, 9) {real, imag} */,
  {32'h3d5d60bc, 32'h3f3f91f0} /* (13, 28, 8) {real, imag} */,
  {32'h3e360ff3, 32'hbe7eea37} /* (13, 28, 7) {real, imag} */,
  {32'hbe5001d2, 32'h3e48ca52} /* (13, 28, 6) {real, imag} */,
  {32'hbf1a2cce, 32'h3e81cccb} /* (13, 28, 5) {real, imag} */,
  {32'h3fd8e3ca, 32'hbf7fa87d} /* (13, 28, 4) {real, imag} */,
  {32'hbf2e96af, 32'h3ec08be4} /* (13, 28, 3) {real, imag} */,
  {32'hc02e7a55, 32'h402671e1} /* (13, 28, 2) {real, imag} */,
  {32'h3ff63424, 32'hbffeb9e1} /* (13, 28, 1) {real, imag} */,
  {32'h3eb80e20, 32'h3eaec639} /* (13, 28, 0) {real, imag} */,
  {32'hc046f1cc, 32'h3faf97c2} /* (13, 27, 31) {real, imag} */,
  {32'h3e65bdfc, 32'hbf962bd2} /* (13, 27, 30) {real, imag} */,
  {32'hbd944124, 32'hbed24846} /* (13, 27, 29) {real, imag} */,
  {32'h3e973b86, 32'h3ec777c2} /* (13, 27, 28) {real, imag} */,
  {32'h3eaeb203, 32'h3bdf9100} /* (13, 27, 27) {real, imag} */,
  {32'hbe36526f, 32'hbf847398} /* (13, 27, 26) {real, imag} */,
  {32'h3e9c90d6, 32'h3edb972a} /* (13, 27, 25) {real, imag} */,
  {32'hbe5c47e2, 32'hbe4b32e7} /* (13, 27, 24) {real, imag} */,
  {32'h3ef5407a, 32'h3c8607c0} /* (13, 27, 23) {real, imag} */,
  {32'hbd775528, 32'hbd81d2b2} /* (13, 27, 22) {real, imag} */,
  {32'h3e2cc1d8, 32'hbf00485e} /* (13, 27, 21) {real, imag} */,
  {32'h3f29452e, 32'h3f5bfb07} /* (13, 27, 20) {real, imag} */,
  {32'hbe967bc6, 32'h3eac0b6e} /* (13, 27, 19) {real, imag} */,
  {32'h3d529ed2, 32'hbe1929b3} /* (13, 27, 18) {real, imag} */,
  {32'hbf39ec88, 32'hbe1ed446} /* (13, 27, 17) {real, imag} */,
  {32'hbe0e8f1e, 32'h3ea1450c} /* (13, 27, 16) {real, imag} */,
  {32'h3e4bab56, 32'hbc957c20} /* (13, 27, 15) {real, imag} */,
  {32'h3e2dddfe, 32'h3e68ec86} /* (13, 27, 14) {real, imag} */,
  {32'hbebad052, 32'h3e559138} /* (13, 27, 13) {real, imag} */,
  {32'hbee795e5, 32'hbe708931} /* (13, 27, 12) {real, imag} */,
  {32'h3f078da4, 32'h3e70f856} /* (13, 27, 11) {real, imag} */,
  {32'h3e91f752, 32'hbdc2755a} /* (13, 27, 10) {real, imag} */,
  {32'h3c489760, 32'hbf8c54eb} /* (13, 27, 9) {real, imag} */,
  {32'hbd7696ac, 32'h3f239c88} /* (13, 27, 8) {real, imag} */,
  {32'h3e61e970, 32'h3eaf145e} /* (13, 27, 7) {real, imag} */,
  {32'h3ea384c4, 32'hbe81ae72} /* (13, 27, 6) {real, imag} */,
  {32'h3f83f2be, 32'hbe9c3dfb} /* (13, 27, 5) {real, imag} */,
  {32'hbf172e40, 32'hbe86de6e} /* (13, 27, 4) {real, imag} */,
  {32'h3e5c56b6, 32'hbf2d358a} /* (13, 27, 3) {real, imag} */,
  {32'h3f013790, 32'hbeb8a0b9} /* (13, 27, 2) {real, imag} */,
  {32'hc0363146, 32'h3e01a5b4} /* (13, 27, 1) {real, imag} */,
  {32'hbfef3a4c, 32'h3f92d780} /* (13, 27, 0) {real, imag} */,
  {32'hbf4455c4, 32'h3f32da9a} /* (13, 26, 31) {real, imag} */,
  {32'h3f77b36e, 32'hbec9b3ee} /* (13, 26, 30) {real, imag} */,
  {32'hbd739ad0, 32'hbe7469ec} /* (13, 26, 29) {real, imag} */,
  {32'hbf2f4012, 32'hbe05c350} /* (13, 26, 28) {real, imag} */,
  {32'hbf2c545c, 32'h3f22170a} /* (13, 26, 27) {real, imag} */,
  {32'hbed43b88, 32'h3f2f63c4} /* (13, 26, 26) {real, imag} */,
  {32'hbeefb5fe, 32'hbe411700} /* (13, 26, 25) {real, imag} */,
  {32'h3f3aa759, 32'hbd1bdf78} /* (13, 26, 24) {real, imag} */,
  {32'hbeb16944, 32'hbedc55bc} /* (13, 26, 23) {real, imag} */,
  {32'hbd91fb8b, 32'h3f22e4eb} /* (13, 26, 22) {real, imag} */,
  {32'hbcce3ed0, 32'hbf5a7a4e} /* (13, 26, 21) {real, imag} */,
  {32'h3df64150, 32'h3d959ac3} /* (13, 26, 20) {real, imag} */,
  {32'h3f035f85, 32'hbddc0136} /* (13, 26, 19) {real, imag} */,
  {32'h3e83e04a, 32'h3ea80c0f} /* (13, 26, 18) {real, imag} */,
  {32'h3e38ad38, 32'h3e8f9a67} /* (13, 26, 17) {real, imag} */,
  {32'hbeb3c81d, 32'h3d24bdec} /* (13, 26, 16) {real, imag} */,
  {32'hbe1c5098, 32'hbd03a1c8} /* (13, 26, 15) {real, imag} */,
  {32'h3e9bf044, 32'h3eb7df40} /* (13, 26, 14) {real, imag} */,
  {32'h3e895335, 32'hbebec5c2} /* (13, 26, 13) {real, imag} */,
  {32'hbe1db331, 32'hbd919c30} /* (13, 26, 12) {real, imag} */,
  {32'hbc848af8, 32'h3daa0f5e} /* (13, 26, 11) {real, imag} */,
  {32'h3dd5be40, 32'hbf18c41e} /* (13, 26, 10) {real, imag} */,
  {32'h3d8229a9, 32'h3e4e1962} /* (13, 26, 9) {real, imag} */,
  {32'h3d049590, 32'hbccf6850} /* (13, 26, 8) {real, imag} */,
  {32'h3d7944b4, 32'h3edb0ebc} /* (13, 26, 7) {real, imag} */,
  {32'h3edbfc44, 32'hbe479ad8} /* (13, 26, 6) {real, imag} */,
  {32'h3f2c914a, 32'hbd6336be} /* (13, 26, 5) {real, imag} */,
  {32'hbe6e3792, 32'h3e957319} /* (13, 26, 4) {real, imag} */,
  {32'h3df57450, 32'h3f1817bb} /* (13, 26, 3) {real, imag} */,
  {32'h3fa9db9c, 32'h3f476efd} /* (13, 26, 2) {real, imag} */,
  {32'hbee64e1a, 32'h3e0adba3} /* (13, 26, 1) {real, imag} */,
  {32'h3e76795a, 32'hbf360a7b} /* (13, 26, 0) {real, imag} */,
  {32'h3ee9c74d, 32'hbfbf104b} /* (13, 25, 31) {real, imag} */,
  {32'h3ee7deae, 32'h3ee6f549} /* (13, 25, 30) {real, imag} */,
  {32'hbdc46cfc, 32'hbed43637} /* (13, 25, 29) {real, imag} */,
  {32'hbf286111, 32'hbe0cb928} /* (13, 25, 28) {real, imag} */,
  {32'h3ee1087c, 32'h3d9e804a} /* (13, 25, 27) {real, imag} */,
  {32'h3ec50506, 32'h3d2df2d8} /* (13, 25, 26) {real, imag} */,
  {32'h3d7833a8, 32'h3da34031} /* (13, 25, 25) {real, imag} */,
  {32'hbefe0184, 32'h3e35bd42} /* (13, 25, 24) {real, imag} */,
  {32'hbe1566b0, 32'hbe8e7455} /* (13, 25, 23) {real, imag} */,
  {32'hbe25bddc, 32'hbeaae05d} /* (13, 25, 22) {real, imag} */,
  {32'hbe1a5f72, 32'hbd046b2e} /* (13, 25, 21) {real, imag} */,
  {32'h3e693226, 32'h3ea2d604} /* (13, 25, 20) {real, imag} */,
  {32'h3d51b3c8, 32'h3ee87e1b} /* (13, 25, 19) {real, imag} */,
  {32'h3da95782, 32'h3cb96acc} /* (13, 25, 18) {real, imag} */,
  {32'h3e4a45a5, 32'hbd8b3fe8} /* (13, 25, 17) {real, imag} */,
  {32'hbecd3524, 32'hbe11d20c} /* (13, 25, 16) {real, imag} */,
  {32'h3e301ccf, 32'hbeca9326} /* (13, 25, 15) {real, imag} */,
  {32'hbdb0bc38, 32'hbf07df6a} /* (13, 25, 14) {real, imag} */,
  {32'hbd9e3db2, 32'hbe75a208} /* (13, 25, 13) {real, imag} */,
  {32'h3edc767b, 32'hbc2d32a0} /* (13, 25, 12) {real, imag} */,
  {32'hbead4107, 32'h3ee4d3b6} /* (13, 25, 11) {real, imag} */,
  {32'h3d65382a, 32'hbea2babc} /* (13, 25, 10) {real, imag} */,
  {32'h3e63b5a9, 32'h3ed238b5} /* (13, 25, 9) {real, imag} */,
  {32'h3e3f1851, 32'h3d8a33e2} /* (13, 25, 8) {real, imag} */,
  {32'h3e8b5e9b, 32'hbc8895f8} /* (13, 25, 7) {real, imag} */,
  {32'hbe4e8e8b, 32'hbaa10700} /* (13, 25, 6) {real, imag} */,
  {32'hbe7eb5ac, 32'hbef34fdc} /* (13, 25, 5) {real, imag} */,
  {32'hbe88dfd9, 32'h3c1577b0} /* (13, 25, 4) {real, imag} */,
  {32'hbdc12d74, 32'h3f0d8e94} /* (13, 25, 3) {real, imag} */,
  {32'h3ea3de80, 32'h3eb004e8} /* (13, 25, 2) {real, imag} */,
  {32'h3ecd5d92, 32'h3e36d18f} /* (13, 25, 1) {real, imag} */,
  {32'hbe41bbab, 32'hbf1745c3} /* (13, 25, 0) {real, imag} */,
  {32'hbfaf2eba, 32'h3f4285bf} /* (13, 24, 31) {real, imag} */,
  {32'h3f6e168a, 32'h3f4566d0} /* (13, 24, 30) {real, imag} */,
  {32'h3f2b6674, 32'h3e05acd5} /* (13, 24, 29) {real, imag} */,
  {32'hbeff26c8, 32'h3f375150} /* (13, 24, 28) {real, imag} */,
  {32'hbd624394, 32'hbe8d3d73} /* (13, 24, 27) {real, imag} */,
  {32'h3efdf968, 32'h3d733aa4} /* (13, 24, 26) {real, imag} */,
  {32'hbe627e16, 32'h3cf43fe4} /* (13, 24, 25) {real, imag} */,
  {32'h3e3c68aa, 32'hbddec6c6} /* (13, 24, 24) {real, imag} */,
  {32'hbe833544, 32'hbe27c22e} /* (13, 24, 23) {real, imag} */,
  {32'hbedc900a, 32'h3e43f10e} /* (13, 24, 22) {real, imag} */,
  {32'h3f9db97e, 32'h3ef37893} /* (13, 24, 21) {real, imag} */,
  {32'h3eb7d65b, 32'hbe9b9e99} /* (13, 24, 20) {real, imag} */,
  {32'h3e85eec9, 32'h3e95ed24} /* (13, 24, 19) {real, imag} */,
  {32'h3e05cd18, 32'h3e814a58} /* (13, 24, 18) {real, imag} */,
  {32'h3d7288a8, 32'hbdeb9f65} /* (13, 24, 17) {real, imag} */,
  {32'h3d86819b, 32'hbf556a2c} /* (13, 24, 16) {real, imag} */,
  {32'hbe17df1d, 32'h3da52309} /* (13, 24, 15) {real, imag} */,
  {32'h3de71316, 32'hbd4fbf30} /* (13, 24, 14) {real, imag} */,
  {32'h3eb4266c, 32'hbe0cd034} /* (13, 24, 13) {real, imag} */,
  {32'hbe9b07d9, 32'h3e03730e} /* (13, 24, 12) {real, imag} */,
  {32'h3eebbe2a, 32'hbd254296} /* (13, 24, 11) {real, imag} */,
  {32'hbf4e4388, 32'hbf011a72} /* (13, 24, 10) {real, imag} */,
  {32'h3e3c2698, 32'hbe960ba1} /* (13, 24, 9) {real, imag} */,
  {32'h3f88647e, 32'h3e8d5614} /* (13, 24, 8) {real, imag} */,
  {32'h3eba8a2f, 32'h3b940f88} /* (13, 24, 7) {real, imag} */,
  {32'hbda6b85a, 32'h3e9b6cd0} /* (13, 24, 6) {real, imag} */,
  {32'h3f7c592c, 32'hbe503528} /* (13, 24, 5) {real, imag} */,
  {32'h3b08a380, 32'hbf48c3f1} /* (13, 24, 4) {real, imag} */,
  {32'h3f2eb311, 32'h3f233ae5} /* (13, 24, 3) {real, imag} */,
  {32'h3f1b81c7, 32'hbf41a334} /* (13, 24, 2) {real, imag} */,
  {32'hbfcf58c9, 32'h3f58d77e} /* (13, 24, 1) {real, imag} */,
  {32'hbf2f2008, 32'h3f04792d} /* (13, 24, 0) {real, imag} */,
  {32'hbe880924, 32'hbf34aedd} /* (13, 23, 31) {real, imag} */,
  {32'hbd04cb04, 32'h3f0cea07} /* (13, 23, 30) {real, imag} */,
  {32'hbd07f916, 32'h3ea2b074} /* (13, 23, 29) {real, imag} */,
  {32'hbe898ff6, 32'hbee895be} /* (13, 23, 28) {real, imag} */,
  {32'h3e963c95, 32'h3ebd15b0} /* (13, 23, 27) {real, imag} */,
  {32'hbedca715, 32'h3eb56770} /* (13, 23, 26) {real, imag} */,
  {32'h3e458030, 32'hbf5f3370} /* (13, 23, 25) {real, imag} */,
  {32'hbdd70b94, 32'hbe02e662} /* (13, 23, 24) {real, imag} */,
  {32'hbece9714, 32'hbefb700d} /* (13, 23, 23) {real, imag} */,
  {32'hbeafb682, 32'h3e9ac6fa} /* (13, 23, 22) {real, imag} */,
  {32'h3ec24fe6, 32'hbbfb2660} /* (13, 23, 21) {real, imag} */,
  {32'hbe297dab, 32'hbe86ea06} /* (13, 23, 20) {real, imag} */,
  {32'hbd9e5efa, 32'hbeb8f85d} /* (13, 23, 19) {real, imag} */,
  {32'h3f31bf8d, 32'h3d03d4b8} /* (13, 23, 18) {real, imag} */,
  {32'hbeaa80fb, 32'h3e81612c} /* (13, 23, 17) {real, imag} */,
  {32'hbe6abf9a, 32'hbea7d7c8} /* (13, 23, 16) {real, imag} */,
  {32'hbec002a4, 32'hbf077b3f} /* (13, 23, 15) {real, imag} */,
  {32'hbe21cd9e, 32'h3e8dddbe} /* (13, 23, 14) {real, imag} */,
  {32'h3e83ac4e, 32'hbc532780} /* (13, 23, 13) {real, imag} */,
  {32'h3df44b37, 32'h3ec1a116} /* (13, 23, 12) {real, imag} */,
  {32'hbf1c89b2, 32'h3da41e4d} /* (13, 23, 11) {real, imag} */,
  {32'hbda645ae, 32'hbe45fc3f} /* (13, 23, 10) {real, imag} */,
  {32'h3f0e1bf5, 32'hbedbe339} /* (13, 23, 9) {real, imag} */,
  {32'hbdb7ded2, 32'hbf06331b} /* (13, 23, 8) {real, imag} */,
  {32'hbe824eaf, 32'h3e12e09c} /* (13, 23, 7) {real, imag} */,
  {32'hbc8a5f70, 32'hbdb4fcf9} /* (13, 23, 6) {real, imag} */,
  {32'hbf0fadd6, 32'hbe7f303e} /* (13, 23, 5) {real, imag} */,
  {32'h3f4802d2, 32'h3e372d2a} /* (13, 23, 4) {real, imag} */,
  {32'h3ed9941a, 32'hbc3a3180} /* (13, 23, 3) {real, imag} */,
  {32'h3f218c14, 32'h3ee6f0fe} /* (13, 23, 2) {real, imag} */,
  {32'h3c759ad0, 32'hbedf00bd} /* (13, 23, 1) {real, imag} */,
  {32'hbdd3332f, 32'h3ed469e4} /* (13, 23, 0) {real, imag} */,
  {32'h3f2dc711, 32'hbdc55a7c} /* (13, 22, 31) {real, imag} */,
  {32'hbd0666a0, 32'h3f2eea29} /* (13, 22, 30) {real, imag} */,
  {32'hbe42680c, 32'h3ed82738} /* (13, 22, 29) {real, imag} */,
  {32'h3f146580, 32'hbd2180c8} /* (13, 22, 28) {real, imag} */,
  {32'h3db54b56, 32'hbe8bc7c1} /* (13, 22, 27) {real, imag} */,
  {32'hbf0819c7, 32'hbe0e4ff8} /* (13, 22, 26) {real, imag} */,
  {32'h3f3cdc03, 32'hbe4b21b2} /* (13, 22, 25) {real, imag} */,
  {32'hbf372f7e, 32'hbf113b78} /* (13, 22, 24) {real, imag} */,
  {32'h3f00c720, 32'h3e4e1d96} /* (13, 22, 23) {real, imag} */,
  {32'hbd15e1b8, 32'h3e8abcfb} /* (13, 22, 22) {real, imag} */,
  {32'h3f26130f, 32'hbe8f9e3a} /* (13, 22, 21) {real, imag} */,
  {32'hbf52cade, 32'hbdb23997} /* (13, 22, 20) {real, imag} */,
  {32'hbec0b2da, 32'h3ce77738} /* (13, 22, 19) {real, imag} */,
  {32'hbe9572b4, 32'h3f1b9d76} /* (13, 22, 18) {real, imag} */,
  {32'h3e197282, 32'hbf047c52} /* (13, 22, 17) {real, imag} */,
  {32'h3e8cbc64, 32'hbe8898c4} /* (13, 22, 16) {real, imag} */,
  {32'h3eaa81dc, 32'hbd296c30} /* (13, 22, 15) {real, imag} */,
  {32'hbe9fe6e2, 32'hbbe5d1d0} /* (13, 22, 14) {real, imag} */,
  {32'h3d020a7c, 32'hbf3469d6} /* (13, 22, 13) {real, imag} */,
  {32'hbeef42cc, 32'hbdc90442} /* (13, 22, 12) {real, imag} */,
  {32'hbea7cfd8, 32'hbd8d4ed0} /* (13, 22, 11) {real, imag} */,
  {32'h3e5484eb, 32'h3e8c8177} /* (13, 22, 10) {real, imag} */,
  {32'h3e4f7b84, 32'h3b3acf40} /* (13, 22, 9) {real, imag} */,
  {32'hbe87b5ba, 32'hbe3e29d8} /* (13, 22, 8) {real, imag} */,
  {32'hbeb5893a, 32'hbd9277a2} /* (13, 22, 7) {real, imag} */,
  {32'h3e44d813, 32'hbef11c7e} /* (13, 22, 6) {real, imag} */,
  {32'h3e5f293c, 32'hbeb21a0b} /* (13, 22, 5) {real, imag} */,
  {32'h3da94be6, 32'h3f1b0f5b} /* (13, 22, 4) {real, imag} */,
  {32'hbe27593d, 32'h3d85be93} /* (13, 22, 3) {real, imag} */,
  {32'h3ea494da, 32'h3ebe2712} /* (13, 22, 2) {real, imag} */,
  {32'hbd730f36, 32'hbf214af6} /* (13, 22, 1) {real, imag} */,
  {32'h3eb196e6, 32'hbedbb700} /* (13, 22, 0) {real, imag} */,
  {32'hbeb39b49, 32'h3ea65f06} /* (13, 21, 31) {real, imag} */,
  {32'hbf4b90c4, 32'hbe425e86} /* (13, 21, 30) {real, imag} */,
  {32'h3ea4024d, 32'h3ebc1d6d} /* (13, 21, 29) {real, imag} */,
  {32'h3d1bb8ea, 32'h3f09e496} /* (13, 21, 28) {real, imag} */,
  {32'h3e4d29f8, 32'hbdc07806} /* (13, 21, 27) {real, imag} */,
  {32'hbe4105f6, 32'hbe977122} /* (13, 21, 26) {real, imag} */,
  {32'hbe25dc36, 32'h3e9a48fa} /* (13, 21, 25) {real, imag} */,
  {32'h3f0ec45d, 32'h3dd03761} /* (13, 21, 24) {real, imag} */,
  {32'h3f01cddc, 32'h3e88e343} /* (13, 21, 23) {real, imag} */,
  {32'h3d81ff48, 32'h3f362de9} /* (13, 21, 22) {real, imag} */,
  {32'hbe4e0f58, 32'h3da4e4db} /* (13, 21, 21) {real, imag} */,
  {32'hbed3cf73, 32'h3e0dac17} /* (13, 21, 20) {real, imag} */,
  {32'h3e823aed, 32'h3e32ac36} /* (13, 21, 19) {real, imag} */,
  {32'h3e43b4ba, 32'hbe80818e} /* (13, 21, 18) {real, imag} */,
  {32'hbd269eec, 32'hbe3c3a6c} /* (13, 21, 17) {real, imag} */,
  {32'hbdab358d, 32'h3e9f04ac} /* (13, 21, 16) {real, imag} */,
  {32'h3e0754f7, 32'hbdc9a734} /* (13, 21, 15) {real, imag} */,
  {32'hbe43e76e, 32'hbe19ed15} /* (13, 21, 14) {real, imag} */,
  {32'h3d0a85a6, 32'h3e16c683} /* (13, 21, 13) {real, imag} */,
  {32'h3f1794b1, 32'hbe8f9875} /* (13, 21, 12) {real, imag} */,
  {32'hbdbfdb08, 32'hbe51e87f} /* (13, 21, 11) {real, imag} */,
  {32'hbdc98028, 32'h3ea6a11d} /* (13, 21, 10) {real, imag} */,
  {32'h3e430698, 32'h3ea324b2} /* (13, 21, 9) {real, imag} */,
  {32'hbe9680e4, 32'h3f18614e} /* (13, 21, 8) {real, imag} */,
  {32'h3e9f9d51, 32'h3f2cde1a} /* (13, 21, 7) {real, imag} */,
  {32'hbd9f3a3c, 32'h3cf27d84} /* (13, 21, 6) {real, imag} */,
  {32'h3f84d9dc, 32'hbf04f27a} /* (13, 21, 5) {real, imag} */,
  {32'hbdd79494, 32'hbe59dc14} /* (13, 21, 4) {real, imag} */,
  {32'h3ea6345a, 32'h3e79e231} /* (13, 21, 3) {real, imag} */,
  {32'hbe041063, 32'hbf151ef5} /* (13, 21, 2) {real, imag} */,
  {32'hbf0dfeed, 32'h3e22fd42} /* (13, 21, 1) {real, imag} */,
  {32'hbf23ae54, 32'h3edb33d4} /* (13, 21, 0) {real, imag} */,
  {32'h3efdd74f, 32'hbe7fc88c} /* (13, 20, 31) {real, imag} */,
  {32'hbe0a0feb, 32'hbe960ccd} /* (13, 20, 30) {real, imag} */,
  {32'h3e5a1ee7, 32'hbde9a56a} /* (13, 20, 29) {real, imag} */,
  {32'h3e192131, 32'h3e9b2403} /* (13, 20, 28) {real, imag} */,
  {32'hbe3d8fc8, 32'h3e972f61} /* (13, 20, 27) {real, imag} */,
  {32'hbcd7901c, 32'h3e8c0bc6} /* (13, 20, 26) {real, imag} */,
  {32'h3d436848, 32'hbe8e1f20} /* (13, 20, 25) {real, imag} */,
  {32'h3eb71681, 32'h3f3e037c} /* (13, 20, 24) {real, imag} */,
  {32'h3ea217ba, 32'hbda91fee} /* (13, 20, 23) {real, imag} */,
  {32'h3f13741a, 32'hbe934163} /* (13, 20, 22) {real, imag} */,
  {32'h3d12aac6, 32'hbd22a7d8} /* (13, 20, 21) {real, imag} */,
  {32'hbf1831b2, 32'h3e5cea3e} /* (13, 20, 20) {real, imag} */,
  {32'h3e4512d5, 32'h3da5ad64} /* (13, 20, 19) {real, imag} */,
  {32'hbeaabd7b, 32'hbc2cac80} /* (13, 20, 18) {real, imag} */,
  {32'h3e7d51f2, 32'hbe95e1fa} /* (13, 20, 17) {real, imag} */,
  {32'h3ec256c7, 32'hbb7a4e60} /* (13, 20, 16) {real, imag} */,
  {32'hbf07c8cd, 32'hbd33ed4e} /* (13, 20, 15) {real, imag} */,
  {32'hbdcb03c4, 32'h3f019fd7} /* (13, 20, 14) {real, imag} */,
  {32'h3d846a60, 32'h3e7352dc} /* (13, 20, 13) {real, imag} */,
  {32'hbdfc01e5, 32'hbe61b8c2} /* (13, 20, 12) {real, imag} */,
  {32'h3f09a971, 32'hbe1101f4} /* (13, 20, 11) {real, imag} */,
  {32'hbed799aa, 32'hbea25968} /* (13, 20, 10) {real, imag} */,
  {32'h3e818a04, 32'h3f19007c} /* (13, 20, 9) {real, imag} */,
  {32'h3cfe79e0, 32'h3e22e54e} /* (13, 20, 8) {real, imag} */,
  {32'h3e2d3606, 32'h3e8e89d7} /* (13, 20, 7) {real, imag} */,
  {32'hbea00f58, 32'h3ea5303a} /* (13, 20, 6) {real, imag} */,
  {32'h3d96ccbf, 32'hbee29c9c} /* (13, 20, 5) {real, imag} */,
  {32'h3dccd2bc, 32'h3da02eae} /* (13, 20, 4) {real, imag} */,
  {32'h3e1acb6b, 32'h3e27677b} /* (13, 20, 3) {real, imag} */,
  {32'h3e98bb7a, 32'hbe8f194c} /* (13, 20, 2) {real, imag} */,
  {32'hbe7714dd, 32'hbec20c3a} /* (13, 20, 1) {real, imag} */,
  {32'h3e9577c5, 32'hbe3e5094} /* (13, 20, 0) {real, imag} */,
  {32'hbcd77128, 32'hbe8e54f4} /* (13, 19, 31) {real, imag} */,
  {32'h3ecd7fca, 32'h3da27610} /* (13, 19, 30) {real, imag} */,
  {32'hbe40ccfa, 32'hbe500e12} /* (13, 19, 29) {real, imag} */,
  {32'h3e6d2ce4, 32'h3ebf26f6} /* (13, 19, 28) {real, imag} */,
  {32'h3e0bdb40, 32'hbe1f1380} /* (13, 19, 27) {real, imag} */,
  {32'hbee9dc64, 32'hbcf449ff} /* (13, 19, 26) {real, imag} */,
  {32'h3f0b46ce, 32'h3d0d89be} /* (13, 19, 25) {real, imag} */,
  {32'hbe896f89, 32'hbb8a9530} /* (13, 19, 24) {real, imag} */,
  {32'h3f1370d2, 32'hbec03763} /* (13, 19, 23) {real, imag} */,
  {32'h3d772da0, 32'hbf0ac702} /* (13, 19, 22) {real, imag} */,
  {32'h3f0f5569, 32'h3f19e6de} /* (13, 19, 21) {real, imag} */,
  {32'hbece3f00, 32'h3ed1db15} /* (13, 19, 20) {real, imag} */,
  {32'hbe5f2ce5, 32'h3e279e87} /* (13, 19, 19) {real, imag} */,
  {32'hbe996368, 32'h3e479c64} /* (13, 19, 18) {real, imag} */,
  {32'h3e8bdef0, 32'hbd5bdf38} /* (13, 19, 17) {real, imag} */,
  {32'h3d89ee53, 32'hbd84d1d2} /* (13, 19, 16) {real, imag} */,
  {32'hbe688e7a, 32'hbe49c748} /* (13, 19, 15) {real, imag} */,
  {32'hbe08c2fc, 32'hbe892e43} /* (13, 19, 14) {real, imag} */,
  {32'h3e0cf60d, 32'h3ecde788} /* (13, 19, 13) {real, imag} */,
  {32'h3e940bfc, 32'hbf1850d8} /* (13, 19, 12) {real, imag} */,
  {32'hbe644154, 32'h3b0bc040} /* (13, 19, 11) {real, imag} */,
  {32'h3e9d8683, 32'h3e002bf2} /* (13, 19, 10) {real, imag} */,
  {32'hbed9ff89, 32'h3f357e97} /* (13, 19, 9) {real, imag} */,
  {32'h3b82ff60, 32'h3e5f9bc2} /* (13, 19, 8) {real, imag} */,
  {32'hb921f800, 32'h3ecd6056} /* (13, 19, 7) {real, imag} */,
  {32'h3dfef437, 32'hbe768747} /* (13, 19, 6) {real, imag} */,
  {32'h3bdfc4e0, 32'h3df1bf63} /* (13, 19, 5) {real, imag} */,
  {32'h3bb60550, 32'hbd7866a0} /* (13, 19, 4) {real, imag} */,
  {32'hbe28e77a, 32'hbe2c6b89} /* (13, 19, 3) {real, imag} */,
  {32'h3da5c2fe, 32'h3e85f5b2} /* (13, 19, 2) {real, imag} */,
  {32'h3e8d8ba8, 32'h3d757bee} /* (13, 19, 1) {real, imag} */,
  {32'hbe3e72e7, 32'hbea01e94} /* (13, 19, 0) {real, imag} */,
  {32'hbe4c06da, 32'h3e5e18c0} /* (13, 18, 31) {real, imag} */,
  {32'hbeb42df6, 32'h3da66c61} /* (13, 18, 30) {real, imag} */,
  {32'h3ddad5c6, 32'hbeb81d8f} /* (13, 18, 29) {real, imag} */,
  {32'h3d54ab8a, 32'h3e20e2de} /* (13, 18, 28) {real, imag} */,
  {32'hbd301364, 32'h3e986912} /* (13, 18, 27) {real, imag} */,
  {32'h3e7724b4, 32'h3ec5a8c8} /* (13, 18, 26) {real, imag} */,
  {32'h3de7134b, 32'hbdc64a78} /* (13, 18, 25) {real, imag} */,
  {32'h3f18e5ce, 32'h3e7edd0b} /* (13, 18, 24) {real, imag} */,
  {32'h3e87939f, 32'hbe3edeaa} /* (13, 18, 23) {real, imag} */,
  {32'h3e49e630, 32'hbe55e684} /* (13, 18, 22) {real, imag} */,
  {32'hbdb8c0e2, 32'h3ed754be} /* (13, 18, 21) {real, imag} */,
  {32'h3ed3fc98, 32'hbe14a579} /* (13, 18, 20) {real, imag} */,
  {32'hbcca35ec, 32'h3de75ae9} /* (13, 18, 19) {real, imag} */,
  {32'hbf17d4bb, 32'hbeca884e} /* (13, 18, 18) {real, imag} */,
  {32'h3caec848, 32'h3e801454} /* (13, 18, 17) {real, imag} */,
  {32'hbe7242fe, 32'h3e92f976} /* (13, 18, 16) {real, imag} */,
  {32'hbdf678ef, 32'h3ee02056} /* (13, 18, 15) {real, imag} */,
  {32'h3ddcf84b, 32'hbe12d94d} /* (13, 18, 14) {real, imag} */,
  {32'h3da9df13, 32'h3e56e8c6} /* (13, 18, 13) {real, imag} */,
  {32'h3ee38884, 32'hbdd88530} /* (13, 18, 12) {real, imag} */,
  {32'h3e2c6de1, 32'hbefd9373} /* (13, 18, 11) {real, imag} */,
  {32'h3e78ddf3, 32'hbdffeecf} /* (13, 18, 10) {real, imag} */,
  {32'hbe3ecf51, 32'hbeb8e88d} /* (13, 18, 9) {real, imag} */,
  {32'h3e38dec9, 32'h3e2961fe} /* (13, 18, 8) {real, imag} */,
  {32'hbd7591dd, 32'h3ed24851} /* (13, 18, 7) {real, imag} */,
  {32'hbe873512, 32'hbeaf93c2} /* (13, 18, 6) {real, imag} */,
  {32'h3dfe47ed, 32'h3e75d1b9} /* (13, 18, 5) {real, imag} */,
  {32'hbd899b6d, 32'h3de8024c} /* (13, 18, 4) {real, imag} */,
  {32'hbc83d60e, 32'hbe76715a} /* (13, 18, 3) {real, imag} */,
  {32'h3d93633c, 32'hbe7e5396} /* (13, 18, 2) {real, imag} */,
  {32'hbd069910, 32'h3ea13749} /* (13, 18, 1) {real, imag} */,
  {32'h3ec368f6, 32'hbda1809a} /* (13, 18, 0) {real, imag} */,
  {32'hbd82e4c3, 32'hbe34d510} /* (13, 17, 31) {real, imag} */,
  {32'hbca0749a, 32'h3d7b6ff4} /* (13, 17, 30) {real, imag} */,
  {32'hbe2e56c0, 32'h3ce89162} /* (13, 17, 29) {real, imag} */,
  {32'hbcb36080, 32'h3e83cfdb} /* (13, 17, 28) {real, imag} */,
  {32'h3e59ea56, 32'hbe0d647c} /* (13, 17, 27) {real, imag} */,
  {32'hbdbdd78c, 32'h3e133e4c} /* (13, 17, 26) {real, imag} */,
  {32'hbbc4fa00, 32'h3d33b460} /* (13, 17, 25) {real, imag} */,
  {32'h3d8c08e7, 32'hbdac70a5} /* (13, 17, 24) {real, imag} */,
  {32'hbcba45e0, 32'h3e716a8c} /* (13, 17, 23) {real, imag} */,
  {32'hbeccbf40, 32'hbe229c18} /* (13, 17, 22) {real, imag} */,
  {32'h3de23768, 32'hbeb2a45c} /* (13, 17, 21) {real, imag} */,
  {32'h3ea84c1f, 32'hbe62201f} /* (13, 17, 20) {real, imag} */,
  {32'h3ef3e296, 32'h3ea34b35} /* (13, 17, 19) {real, imag} */,
  {32'hbd80bb80, 32'hbe631441} /* (13, 17, 18) {real, imag} */,
  {32'h3e0e47a4, 32'h3e7dc46f} /* (13, 17, 17) {real, imag} */,
  {32'h3dc98102, 32'hbee5651c} /* (13, 17, 16) {real, imag} */,
  {32'h3ef7f109, 32'h398cfd00} /* (13, 17, 15) {real, imag} */,
  {32'h3dfed566, 32'hbd001847} /* (13, 17, 14) {real, imag} */,
  {32'h3cb526e8, 32'h3e699656} /* (13, 17, 13) {real, imag} */,
  {32'hbe106268, 32'h3ba540c0} /* (13, 17, 12) {real, imag} */,
  {32'hb8df6600, 32'h3e765f3e} /* (13, 17, 11) {real, imag} */,
  {32'hbdc18bcd, 32'h3edfef96} /* (13, 17, 10) {real, imag} */,
  {32'h3e4abc93, 32'h3e24dd00} /* (13, 17, 9) {real, imag} */,
  {32'h3e4e3534, 32'hbe95c48a} /* (13, 17, 8) {real, imag} */,
  {32'h3e4084a6, 32'h3d911c80} /* (13, 17, 7) {real, imag} */,
  {32'h3c506588, 32'hbd8b80b8} /* (13, 17, 6) {real, imag} */,
  {32'hbc5064e0, 32'h3db18b88} /* (13, 17, 5) {real, imag} */,
  {32'hbdadd383, 32'hbe0732db} /* (13, 17, 4) {real, imag} */,
  {32'h3dff7780, 32'hbefe5476} /* (13, 17, 3) {real, imag} */,
  {32'hbe429cbb, 32'hbe8d56aa} /* (13, 17, 2) {real, imag} */,
  {32'hbe62ec0d, 32'hbd35c15d} /* (13, 17, 1) {real, imag} */,
  {32'hbd9ffe99, 32'hbf117b54} /* (13, 17, 0) {real, imag} */,
  {32'hbe290dca, 32'hbe09a814} /* (13, 16, 31) {real, imag} */,
  {32'hbdb4709d, 32'hbe1296ad} /* (13, 16, 30) {real, imag} */,
  {32'hbe2d5425, 32'hbebc1497} /* (13, 16, 29) {real, imag} */,
  {32'h3b8f268c, 32'hbe898ede} /* (13, 16, 28) {real, imag} */,
  {32'h3e9624b4, 32'h3e10476c} /* (13, 16, 27) {real, imag} */,
  {32'hbdd105e4, 32'h3e257725} /* (13, 16, 26) {real, imag} */,
  {32'hbeb975ce, 32'h3d30b5f2} /* (13, 16, 25) {real, imag} */,
  {32'h3baddba0, 32'hbe3ed29e} /* (13, 16, 24) {real, imag} */,
  {32'h3d80c653, 32'hbf027f50} /* (13, 16, 23) {real, imag} */,
  {32'h3e6430da, 32'hbe32d6a3} /* (13, 16, 22) {real, imag} */,
  {32'h3e29cb18, 32'hbe8bf90a} /* (13, 16, 21) {real, imag} */,
  {32'hbe690af8, 32'h3e5948a0} /* (13, 16, 20) {real, imag} */,
  {32'hbf0eb076, 32'hbe54038b} /* (13, 16, 19) {real, imag} */,
  {32'hbd99ef09, 32'hbed9b9cf} /* (13, 16, 18) {real, imag} */,
  {32'h3e7bc62e, 32'h3e012948} /* (13, 16, 17) {real, imag} */,
  {32'hbe4f80e2, 32'h00000000} /* (13, 16, 16) {real, imag} */,
  {32'h3e7bc62e, 32'hbe012948} /* (13, 16, 15) {real, imag} */,
  {32'hbd99ef09, 32'h3ed9b9cf} /* (13, 16, 14) {real, imag} */,
  {32'hbf0eb076, 32'h3e54038b} /* (13, 16, 13) {real, imag} */,
  {32'hbe690af8, 32'hbe5948a0} /* (13, 16, 12) {real, imag} */,
  {32'h3e29cb18, 32'h3e8bf90a} /* (13, 16, 11) {real, imag} */,
  {32'h3e6430da, 32'h3e32d6a3} /* (13, 16, 10) {real, imag} */,
  {32'h3d80c653, 32'h3f027f50} /* (13, 16, 9) {real, imag} */,
  {32'h3baddba0, 32'h3e3ed29e} /* (13, 16, 8) {real, imag} */,
  {32'hbeb975ce, 32'hbd30b5f2} /* (13, 16, 7) {real, imag} */,
  {32'hbdd105e4, 32'hbe257725} /* (13, 16, 6) {real, imag} */,
  {32'h3e9624b4, 32'hbe10476c} /* (13, 16, 5) {real, imag} */,
  {32'h3b8f268c, 32'h3e898ede} /* (13, 16, 4) {real, imag} */,
  {32'hbe2d5425, 32'h3ebc1497} /* (13, 16, 3) {real, imag} */,
  {32'hbdb4709d, 32'h3e1296ad} /* (13, 16, 2) {real, imag} */,
  {32'hbe290dca, 32'h3e09a814} /* (13, 16, 1) {real, imag} */,
  {32'h3e8812b7, 32'h00000000} /* (13, 16, 0) {real, imag} */,
  {32'hbe62ec0d, 32'h3d35c15d} /* (13, 15, 31) {real, imag} */,
  {32'hbe429cbb, 32'h3e8d56aa} /* (13, 15, 30) {real, imag} */,
  {32'h3dff7780, 32'h3efe5476} /* (13, 15, 29) {real, imag} */,
  {32'hbdadd383, 32'h3e0732db} /* (13, 15, 28) {real, imag} */,
  {32'hbc5064e0, 32'hbdb18b88} /* (13, 15, 27) {real, imag} */,
  {32'h3c506588, 32'h3d8b80b8} /* (13, 15, 26) {real, imag} */,
  {32'h3e4084a6, 32'hbd911c80} /* (13, 15, 25) {real, imag} */,
  {32'h3e4e3534, 32'h3e95c48a} /* (13, 15, 24) {real, imag} */,
  {32'h3e4abc93, 32'hbe24dd00} /* (13, 15, 23) {real, imag} */,
  {32'hbdc18bcd, 32'hbedfef96} /* (13, 15, 22) {real, imag} */,
  {32'hb8df6600, 32'hbe765f3e} /* (13, 15, 21) {real, imag} */,
  {32'hbe106268, 32'hbba540c0} /* (13, 15, 20) {real, imag} */,
  {32'h3cb526e8, 32'hbe699656} /* (13, 15, 19) {real, imag} */,
  {32'h3dfed566, 32'h3d001847} /* (13, 15, 18) {real, imag} */,
  {32'h3ef7f109, 32'hb98cfd00} /* (13, 15, 17) {real, imag} */,
  {32'h3dc98102, 32'h3ee5651c} /* (13, 15, 16) {real, imag} */,
  {32'h3e0e47a4, 32'hbe7dc46f} /* (13, 15, 15) {real, imag} */,
  {32'hbd80bb80, 32'h3e631441} /* (13, 15, 14) {real, imag} */,
  {32'h3ef3e296, 32'hbea34b35} /* (13, 15, 13) {real, imag} */,
  {32'h3ea84c1f, 32'h3e62201f} /* (13, 15, 12) {real, imag} */,
  {32'h3de23768, 32'h3eb2a45c} /* (13, 15, 11) {real, imag} */,
  {32'hbeccbf40, 32'h3e229c18} /* (13, 15, 10) {real, imag} */,
  {32'hbcba45e0, 32'hbe716a8c} /* (13, 15, 9) {real, imag} */,
  {32'h3d8c08e7, 32'h3dac70a5} /* (13, 15, 8) {real, imag} */,
  {32'hbbc4fa00, 32'hbd33b460} /* (13, 15, 7) {real, imag} */,
  {32'hbdbdd78c, 32'hbe133e4c} /* (13, 15, 6) {real, imag} */,
  {32'h3e59ea56, 32'h3e0d647c} /* (13, 15, 5) {real, imag} */,
  {32'hbcb36080, 32'hbe83cfdb} /* (13, 15, 4) {real, imag} */,
  {32'hbe2e56c0, 32'hbce89162} /* (13, 15, 3) {real, imag} */,
  {32'hbca0749a, 32'hbd7b6ff4} /* (13, 15, 2) {real, imag} */,
  {32'hbd82e4c3, 32'h3e34d510} /* (13, 15, 1) {real, imag} */,
  {32'hbd9ffe99, 32'h3f117b54} /* (13, 15, 0) {real, imag} */,
  {32'hbd069910, 32'hbea13749} /* (13, 14, 31) {real, imag} */,
  {32'h3d93633c, 32'h3e7e5396} /* (13, 14, 30) {real, imag} */,
  {32'hbc83d60e, 32'h3e76715a} /* (13, 14, 29) {real, imag} */,
  {32'hbd899b6d, 32'hbde8024c} /* (13, 14, 28) {real, imag} */,
  {32'h3dfe47ed, 32'hbe75d1b9} /* (13, 14, 27) {real, imag} */,
  {32'hbe873512, 32'h3eaf93c2} /* (13, 14, 26) {real, imag} */,
  {32'hbd7591dd, 32'hbed24851} /* (13, 14, 25) {real, imag} */,
  {32'h3e38dec9, 32'hbe2961fe} /* (13, 14, 24) {real, imag} */,
  {32'hbe3ecf51, 32'h3eb8e88d} /* (13, 14, 23) {real, imag} */,
  {32'h3e78ddf3, 32'h3dffeecf} /* (13, 14, 22) {real, imag} */,
  {32'h3e2c6de1, 32'h3efd9373} /* (13, 14, 21) {real, imag} */,
  {32'h3ee38884, 32'h3dd88530} /* (13, 14, 20) {real, imag} */,
  {32'h3da9df13, 32'hbe56e8c6} /* (13, 14, 19) {real, imag} */,
  {32'h3ddcf84b, 32'h3e12d94d} /* (13, 14, 18) {real, imag} */,
  {32'hbdf678ef, 32'hbee02056} /* (13, 14, 17) {real, imag} */,
  {32'hbe7242fe, 32'hbe92f976} /* (13, 14, 16) {real, imag} */,
  {32'h3caec848, 32'hbe801454} /* (13, 14, 15) {real, imag} */,
  {32'hbf17d4bb, 32'h3eca884e} /* (13, 14, 14) {real, imag} */,
  {32'hbcca35ec, 32'hbde75ae9} /* (13, 14, 13) {real, imag} */,
  {32'h3ed3fc98, 32'h3e14a579} /* (13, 14, 12) {real, imag} */,
  {32'hbdb8c0e2, 32'hbed754be} /* (13, 14, 11) {real, imag} */,
  {32'h3e49e630, 32'h3e55e684} /* (13, 14, 10) {real, imag} */,
  {32'h3e87939f, 32'h3e3edeaa} /* (13, 14, 9) {real, imag} */,
  {32'h3f18e5ce, 32'hbe7edd0b} /* (13, 14, 8) {real, imag} */,
  {32'h3de7134b, 32'h3dc64a78} /* (13, 14, 7) {real, imag} */,
  {32'h3e7724b4, 32'hbec5a8c8} /* (13, 14, 6) {real, imag} */,
  {32'hbd301364, 32'hbe986912} /* (13, 14, 5) {real, imag} */,
  {32'h3d54ab8a, 32'hbe20e2de} /* (13, 14, 4) {real, imag} */,
  {32'h3ddad5c6, 32'h3eb81d8f} /* (13, 14, 3) {real, imag} */,
  {32'hbeb42df6, 32'hbda66c61} /* (13, 14, 2) {real, imag} */,
  {32'hbe4c06da, 32'hbe5e18c0} /* (13, 14, 1) {real, imag} */,
  {32'h3ec368f6, 32'h3da1809a} /* (13, 14, 0) {real, imag} */,
  {32'h3e8d8ba8, 32'hbd757bee} /* (13, 13, 31) {real, imag} */,
  {32'h3da5c2fe, 32'hbe85f5b2} /* (13, 13, 30) {real, imag} */,
  {32'hbe28e77a, 32'h3e2c6b89} /* (13, 13, 29) {real, imag} */,
  {32'h3bb60550, 32'h3d7866a0} /* (13, 13, 28) {real, imag} */,
  {32'h3bdfc4e0, 32'hbdf1bf63} /* (13, 13, 27) {real, imag} */,
  {32'h3dfef437, 32'h3e768747} /* (13, 13, 26) {real, imag} */,
  {32'hb921f800, 32'hbecd6056} /* (13, 13, 25) {real, imag} */,
  {32'h3b82ff60, 32'hbe5f9bc2} /* (13, 13, 24) {real, imag} */,
  {32'hbed9ff89, 32'hbf357e97} /* (13, 13, 23) {real, imag} */,
  {32'h3e9d8683, 32'hbe002bf2} /* (13, 13, 22) {real, imag} */,
  {32'hbe644154, 32'hbb0bc040} /* (13, 13, 21) {real, imag} */,
  {32'h3e940bfc, 32'h3f1850d8} /* (13, 13, 20) {real, imag} */,
  {32'h3e0cf60d, 32'hbecde788} /* (13, 13, 19) {real, imag} */,
  {32'hbe08c2fc, 32'h3e892e43} /* (13, 13, 18) {real, imag} */,
  {32'hbe688e7a, 32'h3e49c748} /* (13, 13, 17) {real, imag} */,
  {32'h3d89ee53, 32'h3d84d1d2} /* (13, 13, 16) {real, imag} */,
  {32'h3e8bdef0, 32'h3d5bdf38} /* (13, 13, 15) {real, imag} */,
  {32'hbe996368, 32'hbe479c64} /* (13, 13, 14) {real, imag} */,
  {32'hbe5f2ce5, 32'hbe279e87} /* (13, 13, 13) {real, imag} */,
  {32'hbece3f00, 32'hbed1db15} /* (13, 13, 12) {real, imag} */,
  {32'h3f0f5569, 32'hbf19e6de} /* (13, 13, 11) {real, imag} */,
  {32'h3d772da0, 32'h3f0ac702} /* (13, 13, 10) {real, imag} */,
  {32'h3f1370d2, 32'h3ec03763} /* (13, 13, 9) {real, imag} */,
  {32'hbe896f89, 32'h3b8a9530} /* (13, 13, 8) {real, imag} */,
  {32'h3f0b46ce, 32'hbd0d89be} /* (13, 13, 7) {real, imag} */,
  {32'hbee9dc64, 32'h3cf449ff} /* (13, 13, 6) {real, imag} */,
  {32'h3e0bdb40, 32'h3e1f1380} /* (13, 13, 5) {real, imag} */,
  {32'h3e6d2ce4, 32'hbebf26f6} /* (13, 13, 4) {real, imag} */,
  {32'hbe40ccfa, 32'h3e500e12} /* (13, 13, 3) {real, imag} */,
  {32'h3ecd7fca, 32'hbda27610} /* (13, 13, 2) {real, imag} */,
  {32'hbcd77128, 32'h3e8e54f4} /* (13, 13, 1) {real, imag} */,
  {32'hbe3e72e7, 32'h3ea01e94} /* (13, 13, 0) {real, imag} */,
  {32'hbe7714dd, 32'h3ec20c3a} /* (13, 12, 31) {real, imag} */,
  {32'h3e98bb7a, 32'h3e8f194c} /* (13, 12, 30) {real, imag} */,
  {32'h3e1acb6b, 32'hbe27677b} /* (13, 12, 29) {real, imag} */,
  {32'h3dccd2bc, 32'hbda02eae} /* (13, 12, 28) {real, imag} */,
  {32'h3d96ccbf, 32'h3ee29c9c} /* (13, 12, 27) {real, imag} */,
  {32'hbea00f58, 32'hbea5303a} /* (13, 12, 26) {real, imag} */,
  {32'h3e2d3606, 32'hbe8e89d7} /* (13, 12, 25) {real, imag} */,
  {32'h3cfe79e0, 32'hbe22e54e} /* (13, 12, 24) {real, imag} */,
  {32'h3e818a04, 32'hbf19007c} /* (13, 12, 23) {real, imag} */,
  {32'hbed799aa, 32'h3ea25968} /* (13, 12, 22) {real, imag} */,
  {32'h3f09a971, 32'h3e1101f4} /* (13, 12, 21) {real, imag} */,
  {32'hbdfc01e5, 32'h3e61b8c2} /* (13, 12, 20) {real, imag} */,
  {32'h3d846a60, 32'hbe7352dc} /* (13, 12, 19) {real, imag} */,
  {32'hbdcb03c4, 32'hbf019fd7} /* (13, 12, 18) {real, imag} */,
  {32'hbf07c8cd, 32'h3d33ed4e} /* (13, 12, 17) {real, imag} */,
  {32'h3ec256c7, 32'h3b7a4e60} /* (13, 12, 16) {real, imag} */,
  {32'h3e7d51f2, 32'h3e95e1fa} /* (13, 12, 15) {real, imag} */,
  {32'hbeaabd7b, 32'h3c2cac80} /* (13, 12, 14) {real, imag} */,
  {32'h3e4512d5, 32'hbda5ad64} /* (13, 12, 13) {real, imag} */,
  {32'hbf1831b2, 32'hbe5cea3e} /* (13, 12, 12) {real, imag} */,
  {32'h3d12aac6, 32'h3d22a7d8} /* (13, 12, 11) {real, imag} */,
  {32'h3f13741a, 32'h3e934163} /* (13, 12, 10) {real, imag} */,
  {32'h3ea217ba, 32'h3da91fee} /* (13, 12, 9) {real, imag} */,
  {32'h3eb71681, 32'hbf3e037c} /* (13, 12, 8) {real, imag} */,
  {32'h3d436848, 32'h3e8e1f20} /* (13, 12, 7) {real, imag} */,
  {32'hbcd7901c, 32'hbe8c0bc6} /* (13, 12, 6) {real, imag} */,
  {32'hbe3d8fc8, 32'hbe972f61} /* (13, 12, 5) {real, imag} */,
  {32'h3e192131, 32'hbe9b2403} /* (13, 12, 4) {real, imag} */,
  {32'h3e5a1ee7, 32'h3de9a56a} /* (13, 12, 3) {real, imag} */,
  {32'hbe0a0feb, 32'h3e960ccd} /* (13, 12, 2) {real, imag} */,
  {32'h3efdd74f, 32'h3e7fc88c} /* (13, 12, 1) {real, imag} */,
  {32'h3e9577c5, 32'h3e3e5094} /* (13, 12, 0) {real, imag} */,
  {32'hbf0dfeed, 32'hbe22fd42} /* (13, 11, 31) {real, imag} */,
  {32'hbe041063, 32'h3f151ef5} /* (13, 11, 30) {real, imag} */,
  {32'h3ea6345a, 32'hbe79e231} /* (13, 11, 29) {real, imag} */,
  {32'hbdd79494, 32'h3e59dc14} /* (13, 11, 28) {real, imag} */,
  {32'h3f84d9dc, 32'h3f04f27a} /* (13, 11, 27) {real, imag} */,
  {32'hbd9f3a3c, 32'hbcf27d84} /* (13, 11, 26) {real, imag} */,
  {32'h3e9f9d51, 32'hbf2cde1a} /* (13, 11, 25) {real, imag} */,
  {32'hbe9680e4, 32'hbf18614e} /* (13, 11, 24) {real, imag} */,
  {32'h3e430698, 32'hbea324b2} /* (13, 11, 23) {real, imag} */,
  {32'hbdc98028, 32'hbea6a11d} /* (13, 11, 22) {real, imag} */,
  {32'hbdbfdb08, 32'h3e51e87f} /* (13, 11, 21) {real, imag} */,
  {32'h3f1794b1, 32'h3e8f9875} /* (13, 11, 20) {real, imag} */,
  {32'h3d0a85a6, 32'hbe16c683} /* (13, 11, 19) {real, imag} */,
  {32'hbe43e76e, 32'h3e19ed15} /* (13, 11, 18) {real, imag} */,
  {32'h3e0754f7, 32'h3dc9a734} /* (13, 11, 17) {real, imag} */,
  {32'hbdab358d, 32'hbe9f04ac} /* (13, 11, 16) {real, imag} */,
  {32'hbd269eec, 32'h3e3c3a6c} /* (13, 11, 15) {real, imag} */,
  {32'h3e43b4ba, 32'h3e80818e} /* (13, 11, 14) {real, imag} */,
  {32'h3e823aed, 32'hbe32ac36} /* (13, 11, 13) {real, imag} */,
  {32'hbed3cf73, 32'hbe0dac17} /* (13, 11, 12) {real, imag} */,
  {32'hbe4e0f58, 32'hbda4e4db} /* (13, 11, 11) {real, imag} */,
  {32'h3d81ff48, 32'hbf362de9} /* (13, 11, 10) {real, imag} */,
  {32'h3f01cddc, 32'hbe88e343} /* (13, 11, 9) {real, imag} */,
  {32'h3f0ec45d, 32'hbdd03761} /* (13, 11, 8) {real, imag} */,
  {32'hbe25dc36, 32'hbe9a48fa} /* (13, 11, 7) {real, imag} */,
  {32'hbe4105f6, 32'h3e977122} /* (13, 11, 6) {real, imag} */,
  {32'h3e4d29f8, 32'h3dc07806} /* (13, 11, 5) {real, imag} */,
  {32'h3d1bb8ea, 32'hbf09e496} /* (13, 11, 4) {real, imag} */,
  {32'h3ea4024d, 32'hbebc1d6d} /* (13, 11, 3) {real, imag} */,
  {32'hbf4b90c4, 32'h3e425e86} /* (13, 11, 2) {real, imag} */,
  {32'hbeb39b49, 32'hbea65f06} /* (13, 11, 1) {real, imag} */,
  {32'hbf23ae54, 32'hbedb33d4} /* (13, 11, 0) {real, imag} */,
  {32'hbd730f36, 32'h3f214af6} /* (13, 10, 31) {real, imag} */,
  {32'h3ea494da, 32'hbebe2712} /* (13, 10, 30) {real, imag} */,
  {32'hbe27593d, 32'hbd85be93} /* (13, 10, 29) {real, imag} */,
  {32'h3da94be6, 32'hbf1b0f5b} /* (13, 10, 28) {real, imag} */,
  {32'h3e5f293c, 32'h3eb21a0b} /* (13, 10, 27) {real, imag} */,
  {32'h3e44d813, 32'h3ef11c7e} /* (13, 10, 26) {real, imag} */,
  {32'hbeb5893a, 32'h3d9277a2} /* (13, 10, 25) {real, imag} */,
  {32'hbe87b5ba, 32'h3e3e29d8} /* (13, 10, 24) {real, imag} */,
  {32'h3e4f7b84, 32'hbb3acf40} /* (13, 10, 23) {real, imag} */,
  {32'h3e5484eb, 32'hbe8c8177} /* (13, 10, 22) {real, imag} */,
  {32'hbea7cfd8, 32'h3d8d4ed0} /* (13, 10, 21) {real, imag} */,
  {32'hbeef42cc, 32'h3dc90442} /* (13, 10, 20) {real, imag} */,
  {32'h3d020a7c, 32'h3f3469d6} /* (13, 10, 19) {real, imag} */,
  {32'hbe9fe6e2, 32'h3be5d1d0} /* (13, 10, 18) {real, imag} */,
  {32'h3eaa81dc, 32'h3d296c30} /* (13, 10, 17) {real, imag} */,
  {32'h3e8cbc64, 32'h3e8898c4} /* (13, 10, 16) {real, imag} */,
  {32'h3e197282, 32'h3f047c52} /* (13, 10, 15) {real, imag} */,
  {32'hbe9572b4, 32'hbf1b9d76} /* (13, 10, 14) {real, imag} */,
  {32'hbec0b2da, 32'hbce77738} /* (13, 10, 13) {real, imag} */,
  {32'hbf52cade, 32'h3db23997} /* (13, 10, 12) {real, imag} */,
  {32'h3f26130f, 32'h3e8f9e3a} /* (13, 10, 11) {real, imag} */,
  {32'hbd15e1b8, 32'hbe8abcfb} /* (13, 10, 10) {real, imag} */,
  {32'h3f00c720, 32'hbe4e1d96} /* (13, 10, 9) {real, imag} */,
  {32'hbf372f7e, 32'h3f113b78} /* (13, 10, 8) {real, imag} */,
  {32'h3f3cdc03, 32'h3e4b21b2} /* (13, 10, 7) {real, imag} */,
  {32'hbf0819c7, 32'h3e0e4ff8} /* (13, 10, 6) {real, imag} */,
  {32'h3db54b56, 32'h3e8bc7c1} /* (13, 10, 5) {real, imag} */,
  {32'h3f146580, 32'h3d2180c8} /* (13, 10, 4) {real, imag} */,
  {32'hbe42680c, 32'hbed82738} /* (13, 10, 3) {real, imag} */,
  {32'hbd0666a0, 32'hbf2eea29} /* (13, 10, 2) {real, imag} */,
  {32'h3f2dc711, 32'h3dc55a7c} /* (13, 10, 1) {real, imag} */,
  {32'h3eb196e6, 32'h3edbb700} /* (13, 10, 0) {real, imag} */,
  {32'h3c759ad0, 32'h3edf00bd} /* (13, 9, 31) {real, imag} */,
  {32'h3f218c14, 32'hbee6f0fe} /* (13, 9, 30) {real, imag} */,
  {32'h3ed9941a, 32'h3c3a3180} /* (13, 9, 29) {real, imag} */,
  {32'h3f4802d2, 32'hbe372d2a} /* (13, 9, 28) {real, imag} */,
  {32'hbf0fadd6, 32'h3e7f303e} /* (13, 9, 27) {real, imag} */,
  {32'hbc8a5f70, 32'h3db4fcf9} /* (13, 9, 26) {real, imag} */,
  {32'hbe824eaf, 32'hbe12e09c} /* (13, 9, 25) {real, imag} */,
  {32'hbdb7ded2, 32'h3f06331b} /* (13, 9, 24) {real, imag} */,
  {32'h3f0e1bf5, 32'h3edbe339} /* (13, 9, 23) {real, imag} */,
  {32'hbda645ae, 32'h3e45fc3f} /* (13, 9, 22) {real, imag} */,
  {32'hbf1c89b2, 32'hbda41e4d} /* (13, 9, 21) {real, imag} */,
  {32'h3df44b37, 32'hbec1a116} /* (13, 9, 20) {real, imag} */,
  {32'h3e83ac4e, 32'h3c532780} /* (13, 9, 19) {real, imag} */,
  {32'hbe21cd9e, 32'hbe8dddbe} /* (13, 9, 18) {real, imag} */,
  {32'hbec002a4, 32'h3f077b3f} /* (13, 9, 17) {real, imag} */,
  {32'hbe6abf9a, 32'h3ea7d7c8} /* (13, 9, 16) {real, imag} */,
  {32'hbeaa80fb, 32'hbe81612c} /* (13, 9, 15) {real, imag} */,
  {32'h3f31bf8d, 32'hbd03d4b8} /* (13, 9, 14) {real, imag} */,
  {32'hbd9e5efa, 32'h3eb8f85d} /* (13, 9, 13) {real, imag} */,
  {32'hbe297dab, 32'h3e86ea06} /* (13, 9, 12) {real, imag} */,
  {32'h3ec24fe6, 32'h3bfb2660} /* (13, 9, 11) {real, imag} */,
  {32'hbeafb682, 32'hbe9ac6fa} /* (13, 9, 10) {real, imag} */,
  {32'hbece9714, 32'h3efb700d} /* (13, 9, 9) {real, imag} */,
  {32'hbdd70b94, 32'h3e02e662} /* (13, 9, 8) {real, imag} */,
  {32'h3e458030, 32'h3f5f3370} /* (13, 9, 7) {real, imag} */,
  {32'hbedca715, 32'hbeb56770} /* (13, 9, 6) {real, imag} */,
  {32'h3e963c95, 32'hbebd15b0} /* (13, 9, 5) {real, imag} */,
  {32'hbe898ff6, 32'h3ee895be} /* (13, 9, 4) {real, imag} */,
  {32'hbd07f916, 32'hbea2b074} /* (13, 9, 3) {real, imag} */,
  {32'hbd04cb04, 32'hbf0cea07} /* (13, 9, 2) {real, imag} */,
  {32'hbe880924, 32'h3f34aedd} /* (13, 9, 1) {real, imag} */,
  {32'hbdd3332f, 32'hbed469e4} /* (13, 9, 0) {real, imag} */,
  {32'hbfcf58c9, 32'hbf58d77e} /* (13, 8, 31) {real, imag} */,
  {32'h3f1b81c7, 32'h3f41a334} /* (13, 8, 30) {real, imag} */,
  {32'h3f2eb311, 32'hbf233ae5} /* (13, 8, 29) {real, imag} */,
  {32'h3b08a380, 32'h3f48c3f1} /* (13, 8, 28) {real, imag} */,
  {32'h3f7c592c, 32'h3e503528} /* (13, 8, 27) {real, imag} */,
  {32'hbda6b85a, 32'hbe9b6cd0} /* (13, 8, 26) {real, imag} */,
  {32'h3eba8a2f, 32'hbb940f88} /* (13, 8, 25) {real, imag} */,
  {32'h3f88647e, 32'hbe8d5614} /* (13, 8, 24) {real, imag} */,
  {32'h3e3c2698, 32'h3e960ba1} /* (13, 8, 23) {real, imag} */,
  {32'hbf4e4388, 32'h3f011a72} /* (13, 8, 22) {real, imag} */,
  {32'h3eebbe2a, 32'h3d254296} /* (13, 8, 21) {real, imag} */,
  {32'hbe9b07d9, 32'hbe03730e} /* (13, 8, 20) {real, imag} */,
  {32'h3eb4266c, 32'h3e0cd034} /* (13, 8, 19) {real, imag} */,
  {32'h3de71316, 32'h3d4fbf30} /* (13, 8, 18) {real, imag} */,
  {32'hbe17df1d, 32'hbda52309} /* (13, 8, 17) {real, imag} */,
  {32'h3d86819b, 32'h3f556a2c} /* (13, 8, 16) {real, imag} */,
  {32'h3d7288a8, 32'h3deb9f65} /* (13, 8, 15) {real, imag} */,
  {32'h3e05cd18, 32'hbe814a58} /* (13, 8, 14) {real, imag} */,
  {32'h3e85eec9, 32'hbe95ed24} /* (13, 8, 13) {real, imag} */,
  {32'h3eb7d65b, 32'h3e9b9e99} /* (13, 8, 12) {real, imag} */,
  {32'h3f9db97e, 32'hbef37893} /* (13, 8, 11) {real, imag} */,
  {32'hbedc900a, 32'hbe43f10e} /* (13, 8, 10) {real, imag} */,
  {32'hbe833544, 32'h3e27c22e} /* (13, 8, 9) {real, imag} */,
  {32'h3e3c68aa, 32'h3ddec6c6} /* (13, 8, 8) {real, imag} */,
  {32'hbe627e16, 32'hbcf43fe4} /* (13, 8, 7) {real, imag} */,
  {32'h3efdf968, 32'hbd733aa4} /* (13, 8, 6) {real, imag} */,
  {32'hbd624394, 32'h3e8d3d73} /* (13, 8, 5) {real, imag} */,
  {32'hbeff26c8, 32'hbf375150} /* (13, 8, 4) {real, imag} */,
  {32'h3f2b6674, 32'hbe05acd5} /* (13, 8, 3) {real, imag} */,
  {32'h3f6e168a, 32'hbf4566d0} /* (13, 8, 2) {real, imag} */,
  {32'hbfaf2eba, 32'hbf4285bf} /* (13, 8, 1) {real, imag} */,
  {32'hbf2f2008, 32'hbf04792d} /* (13, 8, 0) {real, imag} */,
  {32'h3ecd5d92, 32'hbe36d18f} /* (13, 7, 31) {real, imag} */,
  {32'h3ea3de80, 32'hbeb004e8} /* (13, 7, 30) {real, imag} */,
  {32'hbdc12d74, 32'hbf0d8e94} /* (13, 7, 29) {real, imag} */,
  {32'hbe88dfd9, 32'hbc1577b0} /* (13, 7, 28) {real, imag} */,
  {32'hbe7eb5ac, 32'h3ef34fdc} /* (13, 7, 27) {real, imag} */,
  {32'hbe4e8e8b, 32'h3aa10700} /* (13, 7, 26) {real, imag} */,
  {32'h3e8b5e9b, 32'h3c8895f8} /* (13, 7, 25) {real, imag} */,
  {32'h3e3f1851, 32'hbd8a33e2} /* (13, 7, 24) {real, imag} */,
  {32'h3e63b5a9, 32'hbed238b5} /* (13, 7, 23) {real, imag} */,
  {32'h3d65382a, 32'h3ea2babc} /* (13, 7, 22) {real, imag} */,
  {32'hbead4107, 32'hbee4d3b6} /* (13, 7, 21) {real, imag} */,
  {32'h3edc767b, 32'h3c2d32a0} /* (13, 7, 20) {real, imag} */,
  {32'hbd9e3db2, 32'h3e75a208} /* (13, 7, 19) {real, imag} */,
  {32'hbdb0bc38, 32'h3f07df6a} /* (13, 7, 18) {real, imag} */,
  {32'h3e301ccf, 32'h3eca9326} /* (13, 7, 17) {real, imag} */,
  {32'hbecd3524, 32'h3e11d20c} /* (13, 7, 16) {real, imag} */,
  {32'h3e4a45a5, 32'h3d8b3fe8} /* (13, 7, 15) {real, imag} */,
  {32'h3da95782, 32'hbcb96acc} /* (13, 7, 14) {real, imag} */,
  {32'h3d51b3c8, 32'hbee87e1b} /* (13, 7, 13) {real, imag} */,
  {32'h3e693226, 32'hbea2d604} /* (13, 7, 12) {real, imag} */,
  {32'hbe1a5f72, 32'h3d046b2e} /* (13, 7, 11) {real, imag} */,
  {32'hbe25bddc, 32'h3eaae05d} /* (13, 7, 10) {real, imag} */,
  {32'hbe1566b0, 32'h3e8e7455} /* (13, 7, 9) {real, imag} */,
  {32'hbefe0184, 32'hbe35bd42} /* (13, 7, 8) {real, imag} */,
  {32'h3d7833a8, 32'hbda34031} /* (13, 7, 7) {real, imag} */,
  {32'h3ec50506, 32'hbd2df2d8} /* (13, 7, 6) {real, imag} */,
  {32'h3ee1087c, 32'hbd9e804a} /* (13, 7, 5) {real, imag} */,
  {32'hbf286111, 32'h3e0cb928} /* (13, 7, 4) {real, imag} */,
  {32'hbdc46cfc, 32'h3ed43637} /* (13, 7, 3) {real, imag} */,
  {32'h3ee7deae, 32'hbee6f549} /* (13, 7, 2) {real, imag} */,
  {32'h3ee9c74d, 32'h3fbf104b} /* (13, 7, 1) {real, imag} */,
  {32'hbe41bbab, 32'h3f1745c3} /* (13, 7, 0) {real, imag} */,
  {32'hbee64e1a, 32'hbe0adba3} /* (13, 6, 31) {real, imag} */,
  {32'h3fa9db9c, 32'hbf476efd} /* (13, 6, 30) {real, imag} */,
  {32'h3df57450, 32'hbf1817bb} /* (13, 6, 29) {real, imag} */,
  {32'hbe6e3792, 32'hbe957319} /* (13, 6, 28) {real, imag} */,
  {32'h3f2c914a, 32'h3d6336be} /* (13, 6, 27) {real, imag} */,
  {32'h3edbfc44, 32'h3e479ad8} /* (13, 6, 26) {real, imag} */,
  {32'h3d7944b4, 32'hbedb0ebc} /* (13, 6, 25) {real, imag} */,
  {32'h3d049590, 32'h3ccf6850} /* (13, 6, 24) {real, imag} */,
  {32'h3d8229a9, 32'hbe4e1962} /* (13, 6, 23) {real, imag} */,
  {32'h3dd5be40, 32'h3f18c41e} /* (13, 6, 22) {real, imag} */,
  {32'hbc848af8, 32'hbdaa0f5e} /* (13, 6, 21) {real, imag} */,
  {32'hbe1db331, 32'h3d919c30} /* (13, 6, 20) {real, imag} */,
  {32'h3e895335, 32'h3ebec5c2} /* (13, 6, 19) {real, imag} */,
  {32'h3e9bf044, 32'hbeb7df40} /* (13, 6, 18) {real, imag} */,
  {32'hbe1c5098, 32'h3d03a1c8} /* (13, 6, 17) {real, imag} */,
  {32'hbeb3c81d, 32'hbd24bdec} /* (13, 6, 16) {real, imag} */,
  {32'h3e38ad38, 32'hbe8f9a67} /* (13, 6, 15) {real, imag} */,
  {32'h3e83e04a, 32'hbea80c0f} /* (13, 6, 14) {real, imag} */,
  {32'h3f035f85, 32'h3ddc0136} /* (13, 6, 13) {real, imag} */,
  {32'h3df64150, 32'hbd959ac3} /* (13, 6, 12) {real, imag} */,
  {32'hbcce3ed0, 32'h3f5a7a4e} /* (13, 6, 11) {real, imag} */,
  {32'hbd91fb8b, 32'hbf22e4eb} /* (13, 6, 10) {real, imag} */,
  {32'hbeb16944, 32'h3edc55bc} /* (13, 6, 9) {real, imag} */,
  {32'h3f3aa759, 32'h3d1bdf78} /* (13, 6, 8) {real, imag} */,
  {32'hbeefb5fe, 32'h3e411700} /* (13, 6, 7) {real, imag} */,
  {32'hbed43b88, 32'hbf2f63c4} /* (13, 6, 6) {real, imag} */,
  {32'hbf2c545c, 32'hbf22170a} /* (13, 6, 5) {real, imag} */,
  {32'hbf2f4012, 32'h3e05c350} /* (13, 6, 4) {real, imag} */,
  {32'hbd739ad0, 32'h3e7469ec} /* (13, 6, 3) {real, imag} */,
  {32'h3f77b36e, 32'h3ec9b3ee} /* (13, 6, 2) {real, imag} */,
  {32'hbf4455c4, 32'hbf32da9a} /* (13, 6, 1) {real, imag} */,
  {32'h3e76795a, 32'h3f360a7b} /* (13, 6, 0) {real, imag} */,
  {32'hc0363146, 32'hbe01a5b4} /* (13, 5, 31) {real, imag} */,
  {32'h3f013790, 32'h3eb8a0b9} /* (13, 5, 30) {real, imag} */,
  {32'h3e5c56b6, 32'h3f2d358a} /* (13, 5, 29) {real, imag} */,
  {32'hbf172e40, 32'h3e86de6e} /* (13, 5, 28) {real, imag} */,
  {32'h3f83f2be, 32'h3e9c3dfb} /* (13, 5, 27) {real, imag} */,
  {32'h3ea384c4, 32'h3e81ae72} /* (13, 5, 26) {real, imag} */,
  {32'h3e61e970, 32'hbeaf145e} /* (13, 5, 25) {real, imag} */,
  {32'hbd7696ac, 32'hbf239c88} /* (13, 5, 24) {real, imag} */,
  {32'h3c489760, 32'h3f8c54eb} /* (13, 5, 23) {real, imag} */,
  {32'h3e91f752, 32'h3dc2755a} /* (13, 5, 22) {real, imag} */,
  {32'h3f078da4, 32'hbe70f856} /* (13, 5, 21) {real, imag} */,
  {32'hbee795e5, 32'h3e708931} /* (13, 5, 20) {real, imag} */,
  {32'hbebad052, 32'hbe559138} /* (13, 5, 19) {real, imag} */,
  {32'h3e2dddfe, 32'hbe68ec86} /* (13, 5, 18) {real, imag} */,
  {32'h3e4bab56, 32'h3c957c20} /* (13, 5, 17) {real, imag} */,
  {32'hbe0e8f1e, 32'hbea1450c} /* (13, 5, 16) {real, imag} */,
  {32'hbf39ec88, 32'h3e1ed446} /* (13, 5, 15) {real, imag} */,
  {32'h3d529ed2, 32'h3e1929b3} /* (13, 5, 14) {real, imag} */,
  {32'hbe967bc6, 32'hbeac0b6e} /* (13, 5, 13) {real, imag} */,
  {32'h3f29452e, 32'hbf5bfb07} /* (13, 5, 12) {real, imag} */,
  {32'h3e2cc1d8, 32'h3f00485e} /* (13, 5, 11) {real, imag} */,
  {32'hbd775528, 32'h3d81d2b2} /* (13, 5, 10) {real, imag} */,
  {32'h3ef5407a, 32'hbc8607c0} /* (13, 5, 9) {real, imag} */,
  {32'hbe5c47e2, 32'h3e4b32e7} /* (13, 5, 8) {real, imag} */,
  {32'h3e9c90d6, 32'hbedb972a} /* (13, 5, 7) {real, imag} */,
  {32'hbe36526f, 32'h3f847398} /* (13, 5, 6) {real, imag} */,
  {32'h3eaeb203, 32'hbbdf9100} /* (13, 5, 5) {real, imag} */,
  {32'h3e973b86, 32'hbec777c2} /* (13, 5, 4) {real, imag} */,
  {32'hbd944124, 32'h3ed24846} /* (13, 5, 3) {real, imag} */,
  {32'h3e65bdfc, 32'h3f962bd2} /* (13, 5, 2) {real, imag} */,
  {32'hc046f1cc, 32'hbfaf97c2} /* (13, 5, 1) {real, imag} */,
  {32'hbfef3a4c, 32'hbf92d780} /* (13, 5, 0) {real, imag} */,
  {32'h3ff63424, 32'h3ffeb9e1} /* (13, 4, 31) {real, imag} */,
  {32'hc02e7a55, 32'hc02671e1} /* (13, 4, 30) {real, imag} */,
  {32'hbf2e96af, 32'hbec08be4} /* (13, 4, 29) {real, imag} */,
  {32'h3fd8e3ca, 32'h3f7fa87d} /* (13, 4, 28) {real, imag} */,
  {32'hbf1a2cce, 32'hbe81cccb} /* (13, 4, 27) {real, imag} */,
  {32'hbe5001d2, 32'hbe48ca52} /* (13, 4, 26) {real, imag} */,
  {32'h3e360ff3, 32'h3e7eea37} /* (13, 4, 25) {real, imag} */,
  {32'h3d5d60bc, 32'hbf3f91f0} /* (13, 4, 24) {real, imag} */,
  {32'h3e0589ea, 32'hbf0d8598} /* (13, 4, 23) {real, imag} */,
  {32'h3e275a64, 32'hbb933c00} /* (13, 4, 22) {real, imag} */,
  {32'hbee2338a, 32'h3e964ae7} /* (13, 4, 21) {real, imag} */,
  {32'hbed910d7, 32'hbed22389} /* (13, 4, 20) {real, imag} */,
  {32'h3ebc092b, 32'hbecbc68e} /* (13, 4, 19) {real, imag} */,
  {32'h3e2b6e14, 32'h3eeace81} /* (13, 4, 18) {real, imag} */,
  {32'h3e97c6a2, 32'hbca10444} /* (13, 4, 17) {real, imag} */,
  {32'h3d5ec480, 32'h3e3f1d7d} /* (13, 4, 16) {real, imag} */,
  {32'h3e5e528c, 32'hbd861a46} /* (13, 4, 15) {real, imag} */,
  {32'hbd732c70, 32'hbecbbd1f} /* (13, 4, 14) {real, imag} */,
  {32'h3e8f1810, 32'hbe982688} /* (13, 4, 13) {real, imag} */,
  {32'hbdbc8419, 32'h3eb5cf08} /* (13, 4, 12) {real, imag} */,
  {32'h3ee72d82, 32'h3ddc4be5} /* (13, 4, 11) {real, imag} */,
  {32'hbef2e426, 32'h3d537064} /* (13, 4, 10) {real, imag} */,
  {32'h3eabf314, 32'h3c1fd3e0} /* (13, 4, 9) {real, imag} */,
  {32'h3c08b118, 32'hbf2796ce} /* (13, 4, 8) {real, imag} */,
  {32'hbeb8111a, 32'hbe6f40a5} /* (13, 4, 7) {real, imag} */,
  {32'hbeb4e8dc, 32'h3e95d063} /* (13, 4, 6) {real, imag} */,
  {32'hbe95d4a8, 32'hbf92b3a1} /* (13, 4, 5) {real, imag} */,
  {32'hbe95f132, 32'h3f150263} /* (13, 4, 4) {real, imag} */,
  {32'hbebd5dd2, 32'h3f466230} /* (13, 4, 3) {real, imag} */,
  {32'hbff38a88, 32'hc014fddf} /* (13, 4, 2) {real, imag} */,
  {32'h40c134bb, 32'h3f23fbe6} /* (13, 4, 1) {real, imag} */,
  {32'h3eb80e20, 32'hbeaec639} /* (13, 4, 0) {real, imag} */,
  {32'hc0a3e835, 32'h3fb61e82} /* (13, 3, 31) {real, imag} */,
  {32'h4031e709, 32'hc01ad8bc} /* (13, 3, 30) {real, imag} */,
  {32'hbec42026, 32'h3f2e3352} /* (13, 3, 29) {real, imag} */,
  {32'h3f819c62, 32'h3f610618} /* (13, 3, 28) {real, imag} */,
  {32'hbe966041, 32'h3e8d634d} /* (13, 3, 27) {real, imag} */,
  {32'hbf5ef5ef, 32'h3c8bc6b0} /* (13, 3, 26) {real, imag} */,
  {32'h3ef954ec, 32'h3e845988} /* (13, 3, 25) {real, imag} */,
  {32'h3e92f958, 32'hbf1f822c} /* (13, 3, 24) {real, imag} */,
  {32'h3ae40c80, 32'h3e68fc8d} /* (13, 3, 23) {real, imag} */,
  {32'h3dd4200c, 32'h3f1f8cf4} /* (13, 3, 22) {real, imag} */,
  {32'hbe2ea28d, 32'hbe353435} /* (13, 3, 21) {real, imag} */,
  {32'hbe8bb8bf, 32'hbec4d7fd} /* (13, 3, 20) {real, imag} */,
  {32'hbe176c15, 32'hbea2b43e} /* (13, 3, 19) {real, imag} */,
  {32'hbdd19008, 32'h3e79caa6} /* (13, 3, 18) {real, imag} */,
  {32'hbe1b4100, 32'h3eb06c75} /* (13, 3, 17) {real, imag} */,
  {32'h3e0c217f, 32'hbd97d838} /* (13, 3, 16) {real, imag} */,
  {32'h3e862dcb, 32'hbef59eb1} /* (13, 3, 15) {real, imag} */,
  {32'hbe940fbd, 32'h3e5fb95f} /* (13, 3, 14) {real, imag} */,
  {32'hbd628a90, 32'h3e5394ce} /* (13, 3, 13) {real, imag} */,
  {32'h3e8734c1, 32'hbebae193} /* (13, 3, 12) {real, imag} */,
  {32'h3f1c4002, 32'hbe2ebbca} /* (13, 3, 11) {real, imag} */,
  {32'hbeb55213, 32'h3e48641c} /* (13, 3, 10) {real, imag} */,
  {32'hbf2665ad, 32'hbf45a785} /* (13, 3, 9) {real, imag} */,
  {32'h3ed44653, 32'hbe632b28} /* (13, 3, 8) {real, imag} */,
  {32'h3f073f7e, 32'h3e545d4e} /* (13, 3, 7) {real, imag} */,
  {32'h3e1ada3e, 32'hbe5748a0} /* (13, 3, 6) {real, imag} */,
  {32'h3e12de62, 32'h3f815ec2} /* (13, 3, 5) {real, imag} */,
  {32'hbe71406c, 32'h3e9adfc1} /* (13, 3, 4) {real, imag} */,
  {32'h3d881768, 32'h3ee725fc} /* (13, 3, 3) {real, imag} */,
  {32'hbf7e4c2e, 32'hc00f0f16} /* (13, 3, 2) {real, imag} */,
  {32'h409fb372, 32'h403e16a3} /* (13, 3, 1) {real, imag} */,
  {32'h3d2660e0, 32'hbeeacc22} /* (13, 3, 0) {real, imag} */,
  {32'hc2015e68, 32'hbf818fb5} /* (13, 2, 31) {real, imag} */,
  {32'h4180fd8c, 32'hc0bc423d} /* (13, 2, 30) {real, imag} */,
  {32'h3f0ee477, 32'h3fb6c940} /* (13, 2, 29) {real, imag} */,
  {32'hbffc727d, 32'h401aa5a0} /* (13, 2, 28) {real, imag} */,
  {32'h3fd2dfd8, 32'hbfaeb7d0} /* (13, 2, 27) {real, imag} */,
  {32'h3f71b084, 32'hbf164333} /* (13, 2, 26) {real, imag} */,
  {32'hbf3f6962, 32'h3ea68bfe} /* (13, 2, 25) {real, imag} */,
  {32'h3f0a2f20, 32'hbf9cc432} /* (13, 2, 24) {real, imag} */,
  {32'hbf2a734e, 32'h3d9195c8} /* (13, 2, 23) {real, imag} */,
  {32'h3d7be8a6, 32'h3e451894} /* (13, 2, 22) {real, imag} */,
  {32'h3f45c5b7, 32'hbf165722} /* (13, 2, 21) {real, imag} */,
  {32'hbe88a3c5, 32'hbd023a6c} /* (13, 2, 20) {real, imag} */,
  {32'hbebd2edf, 32'h3ebdddff} /* (13, 2, 19) {real, imag} */,
  {32'h3e52eaa6, 32'hbe39d64a} /* (13, 2, 18) {real, imag} */,
  {32'h3e271e94, 32'hbdf1e27c} /* (13, 2, 17) {real, imag} */,
  {32'h3dc048ba, 32'hbe89ff00} /* (13, 2, 16) {real, imag} */,
  {32'hbdfa6fe6, 32'h3d80c659} /* (13, 2, 15) {real, imag} */,
  {32'h3e06d73e, 32'hbcc77020} /* (13, 2, 14) {real, imag} */,
  {32'hbdc41c38, 32'hbd727df8} /* (13, 2, 13) {real, imag} */,
  {32'h3ec4da32, 32'hbd19dd4a} /* (13, 2, 12) {real, imag} */,
  {32'h3d8a8dfa, 32'h3e8e0133} /* (13, 2, 11) {real, imag} */,
  {32'hbdf3e737, 32'h3daed053} /* (13, 2, 10) {real, imag} */,
  {32'hbea9a519, 32'hbe9a11d5} /* (13, 2, 9) {real, imag} */,
  {32'h3f320941, 32'hbe489240} /* (13, 2, 8) {real, imag} */,
  {32'hbf04c831, 32'hbec8bc52} /* (13, 2, 7) {real, imag} */,
  {32'h3e42dbcf, 32'h3f20b9a9} /* (13, 2, 6) {real, imag} */,
  {32'h3fad1202, 32'h4012c31d} /* (13, 2, 5) {real, imag} */,
  {32'hc0294460, 32'hc000e95a} /* (13, 2, 4) {real, imag} */,
  {32'h3eb0d0ee, 32'h3e976950} /* (13, 2, 3) {real, imag} */,
  {32'h411f13b5, 32'hc0325670} /* (13, 2, 2) {real, imag} */,
  {32'hc19114de, 32'h40028f76} /* (13, 2, 1) {real, imag} */,
  {32'hc180e086, 32'hc001dfa2} /* (13, 2, 0) {real, imag} */,
  {32'h422a3b02, 32'hc11bc8b7} /* (13, 1, 31) {real, imag} */,
  {32'hc13454ff, 32'hbb5bd280} /* (13, 1, 30) {real, imag} */,
  {32'h3dfb94b8, 32'h3fc90d33} /* (13, 1, 29) {real, imag} */,
  {32'h400aae68, 32'h3f0e8612} /* (13, 1, 28) {real, imag} */,
  {32'hc050536d, 32'h3f139335} /* (13, 1, 27) {real, imag} */,
  {32'h3f715cf4, 32'h3cf31240} /* (13, 1, 26) {real, imag} */,
  {32'h3e4f47b6, 32'h3e0a0662} /* (13, 1, 25) {real, imag} */,
  {32'hbf45ff5d, 32'h3f673836} /* (13, 1, 24) {real, imag} */,
  {32'hbf665271, 32'h3e9d0d82} /* (13, 1, 23) {real, imag} */,
  {32'h3ed6a2ef, 32'h3ee7e2aa} /* (13, 1, 22) {real, imag} */,
  {32'h3e77833e, 32'h3f5130c4} /* (13, 1, 21) {real, imag} */,
  {32'hbe4962ea, 32'hbe16c8ee} /* (13, 1, 20) {real, imag} */,
  {32'h3dba2386, 32'hbe880944} /* (13, 1, 19) {real, imag} */,
  {32'hbcf6c148, 32'h3e9373e6} /* (13, 1, 18) {real, imag} */,
  {32'hbe6b603b, 32'hbeb797e4} /* (13, 1, 17) {real, imag} */,
  {32'h3d1e4d7a, 32'h3deb9c43} /* (13, 1, 16) {real, imag} */,
  {32'hbe15677c, 32'hbe504219} /* (13, 1, 15) {real, imag} */,
  {32'h3e5aa498, 32'h3ec2f752} /* (13, 1, 14) {real, imag} */,
  {32'hbd891a82, 32'hbe127560} /* (13, 1, 13) {real, imag} */,
  {32'h3f032e1e, 32'hbda09c45} /* (13, 1, 12) {real, imag} */,
  {32'hbee84b84, 32'h3e587810} /* (13, 1, 11) {real, imag} */,
  {32'h3e55f99e, 32'hbe5461a2} /* (13, 1, 10) {real, imag} */,
  {32'h3dacbf30, 32'h3e23a6f9} /* (13, 1, 9) {real, imag} */,
  {32'hbe787749, 32'hbfba3654} /* (13, 1, 8) {real, imag} */,
  {32'h3f84747f, 32'h3e6777a5} /* (13, 1, 7) {real, imag} */,
  {32'hbea6abd0, 32'hbfbc441e} /* (13, 1, 6) {real, imag} */,
  {32'hbfdabc92, 32'hbf27d83a} /* (13, 1, 5) {real, imag} */,
  {32'hbf2e13db, 32'h4023767e} /* (13, 1, 4) {real, imag} */,
  {32'hc034c27d, 32'hbe5ada78} /* (13, 1, 3) {real, imag} */,
  {32'hc182e8c4, 32'hc16c369e} /* (13, 1, 2) {real, imag} */,
  {32'h4261b185, 32'h42086478} /* (13, 1, 1) {real, imag} */,
  {32'h4250d69a, 32'h4009118f} /* (13, 1, 0) {real, imag} */,
  {32'h41fa1af5, 32'hc1d98278} /* (13, 0, 31) {real, imag} */,
  {32'hc0b2fb1d, 32'h4104ef35} /* (13, 0, 30) {real, imag} */,
  {32'hbf768721, 32'hbbe20200} /* (13, 0, 29) {real, imag} */,
  {32'h3e1d109e, 32'h3f2c3145} /* (13, 0, 28) {real, imag} */,
  {32'hbfd6f2b6, 32'hbef15a62} /* (13, 0, 27) {real, imag} */,
  {32'h3da55f1a, 32'hbf5f5d9e} /* (13, 0, 26) {real, imag} */,
  {32'hbdd1d744, 32'hbf6aa92c} /* (13, 0, 25) {real, imag} */,
  {32'h3ec054a7, 32'h3f457d3e} /* (13, 0, 24) {real, imag} */,
  {32'hbeb22841, 32'h3f09bb5e} /* (13, 0, 23) {real, imag} */,
  {32'hbf26f5f7, 32'hbe5839a9} /* (13, 0, 22) {real, imag} */,
  {32'hbf076cb2, 32'hbd5b4c0c} /* (13, 0, 21) {real, imag} */,
  {32'h3d812962, 32'h3d8b0f61} /* (13, 0, 20) {real, imag} */,
  {32'h3e4141ed, 32'hbf5ab894} /* (13, 0, 19) {real, imag} */,
  {32'hbd246338, 32'h3ef81e04} /* (13, 0, 18) {real, imag} */,
  {32'h3e622d90, 32'h3eb4fbaf} /* (13, 0, 17) {real, imag} */,
  {32'hbea2e0fd, 32'h00000000} /* (13, 0, 16) {real, imag} */,
  {32'h3e622d90, 32'hbeb4fbaf} /* (13, 0, 15) {real, imag} */,
  {32'hbd246338, 32'hbef81e04} /* (13, 0, 14) {real, imag} */,
  {32'h3e4141ed, 32'h3f5ab894} /* (13, 0, 13) {real, imag} */,
  {32'h3d812962, 32'hbd8b0f61} /* (13, 0, 12) {real, imag} */,
  {32'hbf076cb2, 32'h3d5b4c0c} /* (13, 0, 11) {real, imag} */,
  {32'hbf26f5f7, 32'h3e5839a9} /* (13, 0, 10) {real, imag} */,
  {32'hbeb22841, 32'hbf09bb5e} /* (13, 0, 9) {real, imag} */,
  {32'h3ec054a7, 32'hbf457d3e} /* (13, 0, 8) {real, imag} */,
  {32'hbdd1d744, 32'h3f6aa92c} /* (13, 0, 7) {real, imag} */,
  {32'h3da55f1a, 32'h3f5f5d9e} /* (13, 0, 6) {real, imag} */,
  {32'hbfd6f2b6, 32'h3ef15a62} /* (13, 0, 5) {real, imag} */,
  {32'h3e1d109e, 32'hbf2c3145} /* (13, 0, 4) {real, imag} */,
  {32'hbf768721, 32'h3be20200} /* (13, 0, 3) {real, imag} */,
  {32'hc0b2fb1d, 32'hc104ef35} /* (13, 0, 2) {real, imag} */,
  {32'h41fa1af5, 32'h41d98278} /* (13, 0, 1) {real, imag} */,
  {32'h424de24c, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h428a1a57, 32'hc2242047} /* (12, 31, 31) {real, imag} */,
  {32'hc1978599, 32'h41840624} /* (12, 31, 30) {real, imag} */,
  {32'hbefc7a62, 32'h3c31b2c0} /* (12, 31, 29) {real, imag} */,
  {32'hbf55e5f8, 32'hc00a5466} /* (12, 31, 28) {real, imag} */,
  {32'hc017b820, 32'h3eb30fcc} /* (12, 31, 27) {real, imag} */,
  {32'hbd3dca10, 32'h3f786efc} /* (12, 31, 26) {real, imag} */,
  {32'h3f1c62ee, 32'hbe7e0faa} /* (12, 31, 25) {real, imag} */,
  {32'hbe98265b, 32'h3fad55c8} /* (12, 31, 24) {real, imag} */,
  {32'hbe018bd4, 32'h3e355bcb} /* (12, 31, 23) {real, imag} */,
  {32'hbe90a74c, 32'h3de27cf8} /* (12, 31, 22) {real, imag} */,
  {32'hbd06ff92, 32'h3f2ca6b3} /* (12, 31, 21) {real, imag} */,
  {32'h3e891fa2, 32'h3eedba92} /* (12, 31, 20) {real, imag} */,
  {32'hbda3e17f, 32'h3db5f07d} /* (12, 31, 19) {real, imag} */,
  {32'h3e4a4ffc, 32'h3dd1755e} /* (12, 31, 18) {real, imag} */,
  {32'h3e8515ae, 32'hbe53341d} /* (12, 31, 17) {real, imag} */,
  {32'h3c9d3b54, 32'hbd845edd} /* (12, 31, 16) {real, imag} */,
  {32'h3ea4ae14, 32'hbe9f5256} /* (12, 31, 15) {real, imag} */,
  {32'h3f0bc016, 32'hbe1f11d7} /* (12, 31, 14) {real, imag} */,
  {32'hbe3b366d, 32'hbebb3332} /* (12, 31, 13) {real, imag} */,
  {32'hbf34d5fa, 32'hbd948662} /* (12, 31, 12) {real, imag} */,
  {32'hbf3a5049, 32'hbf508e26} /* (12, 31, 11) {real, imag} */,
  {32'h3f595c2a, 32'hbf51dde3} /* (12, 31, 10) {real, imag} */,
  {32'hbf070fa2, 32'h3e6ff2d8} /* (12, 31, 9) {real, imag} */,
  {32'hbee3a5e7, 32'h3d453760} /* (12, 31, 8) {real, imag} */,
  {32'h3c752830, 32'h3e43bb92} /* (12, 31, 7) {real, imag} */,
  {32'h3eb7bf7e, 32'h3d43a2e8} /* (12, 31, 6) {real, imag} */,
  {32'hc082d0df, 32'h3f12267f} /* (12, 31, 5) {real, imag} */,
  {32'h4028dd31, 32'hbfc3f438} /* (12, 31, 4) {real, imag} */,
  {32'h3c4c7e60, 32'hbf514ad1} /* (12, 31, 3) {real, imag} */,
  {32'hc14996dd, 32'hbf1d7d75} /* (12, 31, 2) {real, imag} */,
  {32'h42482ad4, 32'h411e442a} /* (12, 31, 1) {real, imag} */,
  {32'h42827137, 32'hc07c5dd8} /* (12, 31, 0) {real, imag} */,
  {32'hc1a77074, 32'hc01ec049} /* (12, 30, 31) {real, imag} */,
  {32'h4133884d, 32'h408b266a} /* (12, 30, 30) {real, imag} */,
  {32'h3eead44f, 32'hbdcdec46} /* (12, 30, 29) {real, imag} */,
  {32'hc03f031d, 32'h3fe13fe7} /* (12, 30, 28) {real, imag} */,
  {32'h3f9fe174, 32'hc014b361} /* (12, 30, 27) {real, imag} */,
  {32'h3e554688, 32'hbf6dd322} /* (12, 30, 26) {real, imag} */,
  {32'hbf3aad82, 32'h3e2f3b90} /* (12, 30, 25) {real, imag} */,
  {32'h3f123302, 32'hbeeedf45} /* (12, 30, 24) {real, imag} */,
  {32'hbedda304, 32'h3d56421c} /* (12, 30, 23) {real, imag} */,
  {32'hbe1c5747, 32'h3d83ad38} /* (12, 30, 22) {real, imag} */,
  {32'h3d835d5e, 32'hbf594946} /* (12, 30, 21) {real, imag} */,
  {32'h3e49d1cf, 32'hbeff73f2} /* (12, 30, 20) {real, imag} */,
  {32'h3cd80674, 32'h3e076737} /* (12, 30, 19) {real, imag} */,
  {32'h3f1fb44e, 32'hbf352066} /* (12, 30, 18) {real, imag} */,
  {32'hbeb70633, 32'h3e1610f8} /* (12, 30, 17) {real, imag} */,
  {32'h3dafd85c, 32'hbdde13b1} /* (12, 30, 16) {real, imag} */,
  {32'hbea23768, 32'hbe9c3d1c} /* (12, 30, 15) {real, imag} */,
  {32'h3c87fa99, 32'h3f156b41} /* (12, 30, 14) {real, imag} */,
  {32'h3be4a3a0, 32'hbe407170} /* (12, 30, 13) {real, imag} */,
  {32'hbf0883d2, 32'hbda4e536} /* (12, 30, 12) {real, imag} */,
  {32'h3f182ee2, 32'h3e680d46} /* (12, 30, 11) {real, imag} */,
  {32'hbca616c0, 32'hbe9de8c6} /* (12, 30, 10) {real, imag} */,
  {32'hbed5106e, 32'hbde2f3b2} /* (12, 30, 9) {real, imag} */,
  {32'h3e1fef56, 32'h3fad5feb} /* (12, 30, 8) {real, imag} */,
  {32'hbf2564aa, 32'hbd9e9024} /* (12, 30, 7) {real, imag} */,
  {32'h3f401a4f, 32'h3d838ca4} /* (12, 30, 6) {real, imag} */,
  {32'h3f8a77f5, 32'h3ffff0ed} /* (12, 30, 5) {real, imag} */,
  {32'hbf5dc005, 32'hbfe4f300} /* (12, 30, 4) {real, imag} */,
  {32'h3ec652fa, 32'hbf59fe6a} /* (12, 30, 3) {real, imag} */,
  {32'h4190d81c, 32'h409eaae8} /* (12, 30, 2) {real, imag} */,
  {32'hc217a83c, 32'h3ef8cf0d} /* (12, 30, 1) {real, imag} */,
  {32'hc1970c5e, 32'h402e9758} /* (12, 30, 0) {real, imag} */,
  {32'h4092a3e9, 32'hc06a5577} /* (12, 29, 31) {real, imag} */,
  {32'hbea8edd3, 32'h404fd050} /* (12, 29, 30) {real, imag} */,
  {32'hbf22e696, 32'h3dbb32f8} /* (12, 29, 29) {real, imag} */,
  {32'hbf27b10e, 32'hbdc836a2} /* (12, 29, 28) {real, imag} */,
  {32'h3cefd260, 32'hbf8c5d78} /* (12, 29, 27) {real, imag} */,
  {32'h3f60d454, 32'hbf274a15} /* (12, 29, 26) {real, imag} */,
  {32'h3ec21172, 32'h3f040ec2} /* (12, 29, 25) {real, imag} */,
  {32'hbe9f6a52, 32'hbf11faf9} /* (12, 29, 24) {real, imag} */,
  {32'hbe732a41, 32'hbd21388e} /* (12, 29, 23) {real, imag} */,
  {32'h3edaeefa, 32'h3e573c36} /* (12, 29, 22) {real, imag} */,
  {32'h3b9b77f8, 32'hbd70360a} /* (12, 29, 21) {real, imag} */,
  {32'hbcf77728, 32'hbe802321} /* (12, 29, 20) {real, imag} */,
  {32'h3e60bfcd, 32'hbcc11428} /* (12, 29, 19) {real, imag} */,
  {32'h3ec0d174, 32'h3f366366} /* (12, 29, 18) {real, imag} */,
  {32'h3aa6f400, 32'h3da872c3} /* (12, 29, 17) {real, imag} */,
  {32'h3d2b2892, 32'hbe83207f} /* (12, 29, 16) {real, imag} */,
  {32'hbc7d6064, 32'hbeb0ecf8} /* (12, 29, 15) {real, imag} */,
  {32'hbeb1414e, 32'h3ecda552} /* (12, 29, 14) {real, imag} */,
  {32'hbe38b918, 32'h3e4ad76c} /* (12, 29, 13) {real, imag} */,
  {32'hbe1c74ba, 32'hbcfe70c4} /* (12, 29, 12) {real, imag} */,
  {32'hbe8648f9, 32'hbd893eac} /* (12, 29, 11) {real, imag} */,
  {32'h3d8f9476, 32'h3e7131d8} /* (12, 29, 10) {real, imag} */,
  {32'h3f40d3d6, 32'hbe09f5b6} /* (12, 29, 9) {real, imag} */,
  {32'h3f330560, 32'h3f4cfaf7} /* (12, 29, 8) {real, imag} */,
  {32'h3e679dbc, 32'hbdaaa85f} /* (12, 29, 7) {real, imag} */,
  {32'hbe2f6f4c, 32'hbefea88b} /* (12, 29, 6) {real, imag} */,
  {32'hbf26ba80, 32'hbe03b5f0} /* (12, 29, 5) {real, imag} */,
  {32'h3fc5e4f9, 32'hbfa3d5ea} /* (12, 29, 4) {real, imag} */,
  {32'hbf42fd55, 32'hbef1830f} /* (12, 29, 3) {real, imag} */,
  {32'h400bdc71, 32'h4076a746} /* (12, 29, 2) {real, imag} */,
  {32'hc0af9341, 32'hc006f384} /* (12, 29, 1) {real, imag} */,
  {32'hbe8d2149, 32'hbe47578c} /* (12, 29, 0) {real, imag} */,
  {32'h40b7d9a4, 32'hbf832bea} /* (12, 28, 31) {real, imag} */,
  {32'hc00a8819, 32'h40257cce} /* (12, 28, 30) {real, imag} */,
  {32'h3f263a80, 32'hbe8b4e3e} /* (12, 28, 29) {real, imag} */,
  {32'h3d4ab608, 32'hbedd0d77} /* (12, 28, 28) {real, imag} */,
  {32'h3f0753c1, 32'h3fc69815} /* (12, 28, 27) {real, imag} */,
  {32'hbee4fdca, 32'hbed3d029} /* (12, 28, 26) {real, imag} */,
  {32'hbd700cdf, 32'h3d7d57e8} /* (12, 28, 25) {real, imag} */,
  {32'h3d25d519, 32'h3f9f6337} /* (12, 28, 24) {real, imag} */,
  {32'hbf068d64, 32'hbd1128a8} /* (12, 28, 23) {real, imag} */,
  {32'hbd0847ca, 32'hbf329544} /* (12, 28, 22) {real, imag} */,
  {32'hbee2df5e, 32'h3e592f7f} /* (12, 28, 21) {real, imag} */,
  {32'hbee678b6, 32'h3d0de550} /* (12, 28, 20) {real, imag} */,
  {32'hbe0fada2, 32'hbe9db3ae} /* (12, 28, 19) {real, imag} */,
  {32'h3e5d89da, 32'h3e7ea952} /* (12, 28, 18) {real, imag} */,
  {32'hbdcc54b7, 32'hbddd78bf} /* (12, 28, 17) {real, imag} */,
  {32'h3d37afbe, 32'h3d3b251e} /* (12, 28, 16) {real, imag} */,
  {32'h3e02338f, 32'hbf035316} /* (12, 28, 15) {real, imag} */,
  {32'hbebff452, 32'hbdc7fd40} /* (12, 28, 14) {real, imag} */,
  {32'hbc7d0cf0, 32'h3e5cf40a} /* (12, 28, 13) {real, imag} */,
  {32'h3eacc460, 32'h3e49beae} /* (12, 28, 12) {real, imag} */,
  {32'hbeb11b24, 32'hbf3e53de} /* (12, 28, 11) {real, imag} */,
  {32'hbdc6726b, 32'h3e6b4496} /* (12, 28, 10) {real, imag} */,
  {32'hbe8eedca, 32'h3ed6346c} /* (12, 28, 9) {real, imag} */,
  {32'h3ea3a800, 32'h3ee37b8e} /* (12, 28, 8) {real, imag} */,
  {32'h3f41bb7c, 32'hbd07b904} /* (12, 28, 7) {real, imag} */,
  {32'hbd309fd0, 32'h3e61f966} /* (12, 28, 6) {real, imag} */,
  {32'hbf21bf81, 32'h3f89961c} /* (12, 28, 5) {real, imag} */,
  {32'h3f8d7230, 32'hbe587f00} /* (12, 28, 4) {real, imag} */,
  {32'h3e95a513, 32'h3e9e767e} /* (12, 28, 3) {real, imag} */,
  {32'hc05cea31, 32'h401ef263} /* (12, 28, 2) {real, imag} */,
  {32'h3f727b0d, 32'hc006c60a} /* (12, 28, 1) {real, imag} */,
  {32'h3fa3de4b, 32'h3e2d0483} /* (12, 28, 0) {real, imag} */,
  {32'hc00f1aa0, 32'h401778cd} /* (12, 27, 31) {real, imag} */,
  {32'h3f16b9ec, 32'hbfbe9b2e} /* (12, 27, 30) {real, imag} */,
  {32'h3d169efc, 32'h3ea47fc8} /* (12, 27, 29) {real, imag} */,
  {32'hbdd18a98, 32'h3f8fa1ff} /* (12, 27, 28) {real, imag} */,
  {32'h3fa2f932, 32'hbf4a88df} /* (12, 27, 27) {real, imag} */,
  {32'h3e8ef28b, 32'hbe388fac} /* (12, 27, 26) {real, imag} */,
  {32'hbed6146b, 32'h3dd49664} /* (12, 27, 25) {real, imag} */,
  {32'h3ebe32db, 32'h3d3d766c} /* (12, 27, 24) {real, imag} */,
  {32'h3f4a58fd, 32'hbf2897eb} /* (12, 27, 23) {real, imag} */,
  {32'hbe9a86c0, 32'hbecbbc92} /* (12, 27, 22) {real, imag} */,
  {32'h3e6f5cb0, 32'hbebb6d1c} /* (12, 27, 21) {real, imag} */,
  {32'h3ee46224, 32'h3d2a26f8} /* (12, 27, 20) {real, imag} */,
  {32'hbe6751e9, 32'hbe634ba0} /* (12, 27, 19) {real, imag} */,
  {32'hbf27de4e, 32'hbe52b6f0} /* (12, 27, 18) {real, imag} */,
  {32'h3d896b4e, 32'hbd323a2e} /* (12, 27, 17) {real, imag} */,
  {32'h3e7af88e, 32'hbba99bc0} /* (12, 27, 16) {real, imag} */,
  {32'h3dba5002, 32'h3e7f7cd6} /* (12, 27, 15) {real, imag} */,
  {32'hbe8e6636, 32'h3dcb7434} /* (12, 27, 14) {real, imag} */,
  {32'hbdc710e5, 32'hbf3bc358} /* (12, 27, 13) {real, imag} */,
  {32'h3e219a58, 32'h3debb680} /* (12, 27, 12) {real, imag} */,
  {32'h3f15e960, 32'h3d63c09e} /* (12, 27, 11) {real, imag} */,
  {32'h3eb6a4df, 32'h3e4e5ece} /* (12, 27, 10) {real, imag} */,
  {32'h3ebbef24, 32'h3da990b2} /* (12, 27, 9) {real, imag} */,
  {32'h3ee46d1a, 32'h3f214e6a} /* (12, 27, 8) {real, imag} */,
  {32'h3e91643e, 32'h3efbe684} /* (12, 27, 7) {real, imag} */,
  {32'hbe0a0898, 32'h3dc530d6} /* (12, 27, 6) {real, imag} */,
  {32'h3ebd4f8e, 32'hbf5b9038} /* (12, 27, 5) {real, imag} */,
  {32'hbedd801a, 32'hbf9fcc3e} /* (12, 27, 4) {real, imag} */,
  {32'hbdd46108, 32'hbbf14600} /* (12, 27, 3) {real, imag} */,
  {32'h3f20296b, 32'hbec39b3d} /* (12, 27, 2) {real, imag} */,
  {32'hc05779ce, 32'h3f01bdaa} /* (12, 27, 1) {real, imag} */,
  {32'hc0336c5a, 32'h3f51c64b} /* (12, 27, 0) {real, imag} */,
  {32'h3f40688c, 32'h3ea56c48} /* (12, 26, 31) {real, imag} */,
  {32'h3e621dd1, 32'h3e282dc7} /* (12, 26, 30) {real, imag} */,
  {32'hbd5a4105, 32'hbed058cc} /* (12, 26, 29) {real, imag} */,
  {32'h3ea76cbc, 32'h3f06d6ae} /* (12, 26, 28) {real, imag} */,
  {32'h3eec1961, 32'h3f6b224e} /* (12, 26, 27) {real, imag} */,
  {32'h3d0748fe, 32'h3f0dff78} /* (12, 26, 26) {real, imag} */,
  {32'hbea09ccd, 32'hbe43c6fc} /* (12, 26, 25) {real, imag} */,
  {32'h3e76e78d, 32'h3e9d95cf} /* (12, 26, 24) {real, imag} */,
  {32'hbf71ccb5, 32'h3da0763e} /* (12, 26, 23) {real, imag} */,
  {32'hbf14698a, 32'h3ec35a5e} /* (12, 26, 22) {real, imag} */,
  {32'hbda2c197, 32'hbc95855c} /* (12, 26, 21) {real, imag} */,
  {32'hbd579764, 32'hbe2b156b} /* (12, 26, 20) {real, imag} */,
  {32'hbe37ac2e, 32'hbe4b43c5} /* (12, 26, 19) {real, imag} */,
  {32'h3e95d21d, 32'h3ec410c2} /* (12, 26, 18) {real, imag} */,
  {32'h3da93c3f, 32'h3cce4a20} /* (12, 26, 17) {real, imag} */,
  {32'hbe78fa08, 32'hbdf247e3} /* (12, 26, 16) {real, imag} */,
  {32'h3e780efa, 32'h3e906fff} /* (12, 26, 15) {real, imag} */,
  {32'hbea77344, 32'h3d978d2d} /* (12, 26, 14) {real, imag} */,
  {32'h3ec5368a, 32'hbee748ca} /* (12, 26, 13) {real, imag} */,
  {32'h3e825b10, 32'h3d5da844} /* (12, 26, 12) {real, imag} */,
  {32'h3d759cd4, 32'h3dc98209} /* (12, 26, 11) {real, imag} */,
  {32'h3f56f712, 32'h3eb0ef90} /* (12, 26, 10) {real, imag} */,
  {32'hbcadade8, 32'h3e11acab} /* (12, 26, 9) {real, imag} */,
  {32'hbeac8ba4, 32'hbe2e2e86} /* (12, 26, 8) {real, imag} */,
  {32'h3d15db3c, 32'h3e7a869f} /* (12, 26, 7) {real, imag} */,
  {32'hbcd27f58, 32'hbe8adc55} /* (12, 26, 6) {real, imag} */,
  {32'hbdcd6dd6, 32'hbef7188a} /* (12, 26, 5) {real, imag} */,
  {32'hbe2373d8, 32'h3f0ec897} /* (12, 26, 4) {real, imag} */,
  {32'h3ef0c5af, 32'h3f0cd5b2} /* (12, 26, 3) {real, imag} */,
  {32'h3f870773, 32'h3dadedc6} /* (12, 26, 2) {real, imag} */,
  {32'h3ec8d60a, 32'h3f09383b} /* (12, 26, 1) {real, imag} */,
  {32'h3e579f30, 32'hbf092917} /* (12, 26, 0) {real, imag} */,
  {32'h3f32866c, 32'hbf1a62ae} /* (12, 25, 31) {real, imag} */,
  {32'hbeaad936, 32'h3e8de49f} /* (12, 25, 30) {real, imag} */,
  {32'hbf2baeea, 32'hbf219736} /* (12, 25, 29) {real, imag} */,
  {32'hbe89305b, 32'hbf435708} /* (12, 25, 28) {real, imag} */,
  {32'hbb904e60, 32'hbe6dab12} /* (12, 25, 27) {real, imag} */,
  {32'h3e8e4e3f, 32'h3c5027e0} /* (12, 25, 26) {real, imag} */,
  {32'hbe6e6d63, 32'hbd7c670f} /* (12, 25, 25) {real, imag} */,
  {32'h3eb73284, 32'h3dc92c72} /* (12, 25, 24) {real, imag} */,
  {32'hbea9ec26, 32'h3e902867} /* (12, 25, 23) {real, imag} */,
  {32'h3eb7f084, 32'hbe4eae74} /* (12, 25, 22) {real, imag} */,
  {32'h3f46678c, 32'h3e89de8a} /* (12, 25, 21) {real, imag} */,
  {32'h3df6e958, 32'h3d6a1e50} /* (12, 25, 20) {real, imag} */,
  {32'hbd4ee135, 32'h3f209ca0} /* (12, 25, 19) {real, imag} */,
  {32'hbe3fcbee, 32'h3d0a4222} /* (12, 25, 18) {real, imag} */,
  {32'h3e995c5a, 32'h3dda43c5} /* (12, 25, 17) {real, imag} */,
  {32'hbeba4e07, 32'hbe9ec426} /* (12, 25, 16) {real, imag} */,
  {32'hbe3aef45, 32'hbe87c313} /* (12, 25, 15) {real, imag} */,
  {32'h3cb9c740, 32'hbe503f0a} /* (12, 25, 14) {real, imag} */,
  {32'hbe5b93a7, 32'hbe540646} /* (12, 25, 13) {real, imag} */,
  {32'h3e4ba3a8, 32'hbe8a611a} /* (12, 25, 12) {real, imag} */,
  {32'h3f31bf63, 32'h3eb0db68} /* (12, 25, 11) {real, imag} */,
  {32'hbdc94967, 32'hbf1576f0} /* (12, 25, 10) {real, imag} */,
  {32'hbee8ce72, 32'h3e6cdbfa} /* (12, 25, 9) {real, imag} */,
  {32'hbe469ca6, 32'h3eeda232} /* (12, 25, 8) {real, imag} */,
  {32'h3f0e6da7, 32'hbf00ff3c} /* (12, 25, 7) {real, imag} */,
  {32'h3d58d4d9, 32'hbe94ef5a} /* (12, 25, 6) {real, imag} */,
  {32'hbd8de3ca, 32'h3ed9da9e} /* (12, 25, 5) {real, imag} */,
  {32'hbbf71ae0, 32'hbe80fbe1} /* (12, 25, 4) {real, imag} */,
  {32'hbe266d90, 32'hbd9902ab} /* (12, 25, 3) {real, imag} */,
  {32'h3d8ba543, 32'h3f283cd6} /* (12, 25, 2) {real, imag} */,
  {32'h3f0864b8, 32'h3f06813c} /* (12, 25, 1) {real, imag} */,
  {32'h3d0a5948, 32'hbe9dbf1c} /* (12, 25, 0) {real, imag} */,
  {32'hbfa71c54, 32'hbdb36e38} /* (12, 24, 31) {real, imag} */,
  {32'h3e9f72d3, 32'hbf1c418b} /* (12, 24, 30) {real, imag} */,
  {32'hbe4c5146, 32'hbe52beb6} /* (12, 24, 29) {real, imag} */,
  {32'hbf7e4fbb, 32'h3f81c3e9} /* (12, 24, 28) {real, imag} */,
  {32'h3f38f709, 32'h3e925a6d} /* (12, 24, 27) {real, imag} */,
  {32'h3ebbce2b, 32'h3eefa4ac} /* (12, 24, 26) {real, imag} */,
  {32'hbf102ce7, 32'h3d294934} /* (12, 24, 25) {real, imag} */,
  {32'h3ea96b24, 32'h3da807c6} /* (12, 24, 24) {real, imag} */,
  {32'h3df7b3d4, 32'hbd032c72} /* (12, 24, 23) {real, imag} */,
  {32'h3f18462c, 32'hbdd75580} /* (12, 24, 22) {real, imag} */,
  {32'h3e0d3d5d, 32'h3f11cd84} /* (12, 24, 21) {real, imag} */,
  {32'h3ea14265, 32'hbf70923e} /* (12, 24, 20) {real, imag} */,
  {32'hbf5fd550, 32'hbf02e46c} /* (12, 24, 19) {real, imag} */,
  {32'hbe890ca4, 32'h3ebd1332} /* (12, 24, 18) {real, imag} */,
  {32'h3df2397a, 32'hbed0a0ba} /* (12, 24, 17) {real, imag} */,
  {32'h3e0bee82, 32'h3e032daf} /* (12, 24, 16) {real, imag} */,
  {32'h3e755ed6, 32'h3e045e9e} /* (12, 24, 15) {real, imag} */,
  {32'h3f05b8f0, 32'hbd229cb2} /* (12, 24, 14) {real, imag} */,
  {32'hbee02cc6, 32'h3e8ace42} /* (12, 24, 13) {real, imag} */,
  {32'h3f043314, 32'h3e40ca62} /* (12, 24, 12) {real, imag} */,
  {32'h3f0af3dd, 32'h3b8b2610} /* (12, 24, 11) {real, imag} */,
  {32'hbecc24f9, 32'hbf0b88c2} /* (12, 24, 10) {real, imag} */,
  {32'h3d4af790, 32'h3e9e647d} /* (12, 24, 9) {real, imag} */,
  {32'h3da65bd6, 32'hbe94c569} /* (12, 24, 8) {real, imag} */,
  {32'h3d3b2a06, 32'h3eaa99d8} /* (12, 24, 7) {real, imag} */,
  {32'h3dd7b212, 32'hbe989799} /* (12, 24, 6) {real, imag} */,
  {32'h3f2c1f4b, 32'h3e9a1a5d} /* (12, 24, 5) {real, imag} */,
  {32'h3e89fe48, 32'h3f00a829} /* (12, 24, 4) {real, imag} */,
  {32'h3dbe2a16, 32'h3efd3084} /* (12, 24, 3) {real, imag} */,
  {32'h3f67b91d, 32'hbecf02ca} /* (12, 24, 2) {real, imag} */,
  {32'hbfb68768, 32'h3f43492a} /* (12, 24, 1) {real, imag} */,
  {32'hbf218586, 32'h3f659562} /* (12, 24, 0) {real, imag} */,
  {32'h3f8c88e0, 32'hbefba136} /* (12, 23, 31) {real, imag} */,
  {32'hbeb2cf29, 32'h3ec50dc2} /* (12, 23, 30) {real, imag} */,
  {32'h3f14694d, 32'h3f273b66} /* (12, 23, 29) {real, imag} */,
  {32'hbea3440a, 32'hbe8694be} /* (12, 23, 28) {real, imag} */,
  {32'hbe8e991e, 32'hbeec5cd1} /* (12, 23, 27) {real, imag} */,
  {32'hbf0d0231, 32'hbed6ed2e} /* (12, 23, 26) {real, imag} */,
  {32'h3eb47e58, 32'hbe810b1f} /* (12, 23, 25) {real, imag} */,
  {32'hbd48f9b8, 32'h3e0550f6} /* (12, 23, 24) {real, imag} */,
  {32'h3f28d9da, 32'h3e01fdc0} /* (12, 23, 23) {real, imag} */,
  {32'hbec4eb94, 32'h3e904fb8} /* (12, 23, 22) {real, imag} */,
  {32'hbefee0a2, 32'h3d647501} /* (12, 23, 21) {real, imag} */,
  {32'hbe85bdbf, 32'h3e426312} /* (12, 23, 20) {real, imag} */,
  {32'hbec508e0, 32'hbe8603a0} /* (12, 23, 19) {real, imag} */,
  {32'h3e2feba0, 32'h3e01e7d2} /* (12, 23, 18) {real, imag} */,
  {32'h3dcf1389, 32'hbb737140} /* (12, 23, 17) {real, imag} */,
  {32'hbc959970, 32'hbe48ca82} /* (12, 23, 16) {real, imag} */,
  {32'h3de2ee80, 32'hbe56a21a} /* (12, 23, 15) {real, imag} */,
  {32'h3dabe536, 32'h3e16da72} /* (12, 23, 14) {real, imag} */,
  {32'h3eeb7e76, 32'hbdd0ba5d} /* (12, 23, 13) {real, imag} */,
  {32'h3e2cd43c, 32'hbc888848} /* (12, 23, 12) {real, imag} */,
  {32'hbe54d71b, 32'hbdde34ba} /* (12, 23, 11) {real, imag} */,
  {32'h3dc731f8, 32'h3e452e51} /* (12, 23, 10) {real, imag} */,
  {32'h3de7e15b, 32'hbec4c022} /* (12, 23, 9) {real, imag} */,
  {32'hbf69029f, 32'h3df3fe1a} /* (12, 23, 8) {real, imag} */,
  {32'hbe8bfbea, 32'h3e309ac7} /* (12, 23, 7) {real, imag} */,
  {32'hbd91b4d8, 32'hbd976184} /* (12, 23, 6) {real, imag} */,
  {32'hbedfdec0, 32'hbe1180ca} /* (12, 23, 5) {real, imag} */,
  {32'h3e130aa4, 32'h3e9f0be6} /* (12, 23, 4) {real, imag} */,
  {32'h3defb2a9, 32'h3e75a3de} /* (12, 23, 3) {real, imag} */,
  {32'h3e7139b0, 32'h3e0ba34c} /* (12, 23, 2) {real, imag} */,
  {32'hbf2c26a2, 32'hbed81372} /* (12, 23, 1) {real, imag} */,
  {32'hbe5846d4, 32'h3eb62a85} /* (12, 23, 0) {real, imag} */,
  {32'h3dfe1902, 32'hbe5c5910} /* (12, 22, 31) {real, imag} */,
  {32'hbe2b7df5, 32'h3f516798} /* (12, 22, 30) {real, imag} */,
  {32'h3dd5a988, 32'h3d24b378} /* (12, 22, 29) {real, imag} */,
  {32'hbeab3b36, 32'hbf3e0441} /* (12, 22, 28) {real, imag} */,
  {32'h3f12f1d9, 32'h3f0ec082} /* (12, 22, 27) {real, imag} */,
  {32'h3da65c2a, 32'h3f002e80} /* (12, 22, 26) {real, imag} */,
  {32'h3e86ba6c, 32'hbef8915e} /* (12, 22, 25) {real, imag} */,
  {32'hbd582168, 32'h3e015e4e} /* (12, 22, 24) {real, imag} */,
  {32'h3e13d84c, 32'h3d948162} /* (12, 22, 23) {real, imag} */,
  {32'hbee3e382, 32'hbe8fcf0f} /* (12, 22, 22) {real, imag} */,
  {32'h3d7092a0, 32'h3e7888d9} /* (12, 22, 21) {real, imag} */,
  {32'hbe2d19d0, 32'h3ee55c6c} /* (12, 22, 20) {real, imag} */,
  {32'h3de6aef2, 32'h3eaf487a} /* (12, 22, 19) {real, imag} */,
  {32'h3ca27404, 32'h3d2d560c} /* (12, 22, 18) {real, imag} */,
  {32'h3e851009, 32'hbeba4702} /* (12, 22, 17) {real, imag} */,
  {32'hbeec8e7e, 32'hbdfc09dd} /* (12, 22, 16) {real, imag} */,
  {32'hbdc4ab12, 32'h3e0a335e} /* (12, 22, 15) {real, imag} */,
  {32'hbccae3b0, 32'hbe8ad5ee} /* (12, 22, 14) {real, imag} */,
  {32'h3ebb9b44, 32'h3e34e42a} /* (12, 22, 13) {real, imag} */,
  {32'h3d206ae4, 32'h3d9c2027} /* (12, 22, 12) {real, imag} */,
  {32'h3ecfaca5, 32'h3ed87aac} /* (12, 22, 11) {real, imag} */,
  {32'h3e9a7328, 32'hbcd635a8} /* (12, 22, 10) {real, imag} */,
  {32'hbf2078e2, 32'hbeef731e} /* (12, 22, 9) {real, imag} */,
  {32'h3efc55c3, 32'h3efc540c} /* (12, 22, 8) {real, imag} */,
  {32'hbf039a38, 32'hbdfccb74} /* (12, 22, 7) {real, imag} */,
  {32'h3dc1c780, 32'h3eddd260} /* (12, 22, 6) {real, imag} */,
  {32'hbedde302, 32'hbea06066} /* (12, 22, 5) {real, imag} */,
  {32'h3e07cbfa, 32'hbe0c8678} /* (12, 22, 4) {real, imag} */,
  {32'hbe626c69, 32'h3e732102} /* (12, 22, 3) {real, imag} */,
  {32'hbe08eda4, 32'hb973f800} /* (12, 22, 2) {real, imag} */,
  {32'h3dcabc3a, 32'hbefacf8d} /* (12, 22, 1) {real, imag} */,
  {32'hbd4dcbf4, 32'h3d97835a} /* (12, 22, 0) {real, imag} */,
  {32'hbf834f73, 32'h3f03b45a} /* (12, 21, 31) {real, imag} */,
  {32'hbedf6022, 32'hbe0e3276} /* (12, 21, 30) {real, imag} */,
  {32'h3f4c6d1a, 32'h3e2fa69c} /* (12, 21, 29) {real, imag} */,
  {32'h3d026e04, 32'hbcbce460} /* (12, 21, 28) {real, imag} */,
  {32'hbe5ecbde, 32'hbebb6016} /* (12, 21, 27) {real, imag} */,
  {32'hbdfd1fda, 32'h3f052fba} /* (12, 21, 26) {real, imag} */,
  {32'h3e228a16, 32'hbe5698ec} /* (12, 21, 25) {real, imag} */,
  {32'hbd0f15a0, 32'hbd021db8} /* (12, 21, 24) {real, imag} */,
  {32'hbcaf3f30, 32'h3f04f9f2} /* (12, 21, 23) {real, imag} */,
  {32'h3c0c34a0, 32'hbe53f7b6} /* (12, 21, 22) {real, imag} */,
  {32'hbcdc20a8, 32'hbee69013} /* (12, 21, 21) {real, imag} */,
  {32'hbeb219e8, 32'h3d92b9ce} /* (12, 21, 20) {real, imag} */,
  {32'h3ddeaaac, 32'h3e133988} /* (12, 21, 19) {real, imag} */,
  {32'hbdfaa75d, 32'h3ebde7ae} /* (12, 21, 18) {real, imag} */,
  {32'hbe5f6904, 32'h3e0f6480} /* (12, 21, 17) {real, imag} */,
  {32'hbed5b970, 32'h3e4bf572} /* (12, 21, 16) {real, imag} */,
  {32'h3e7092f5, 32'hbe909226} /* (12, 21, 15) {real, imag} */,
  {32'hbec86a28, 32'h3d417662} /* (12, 21, 14) {real, imag} */,
  {32'h3f4734fa, 32'hbccd33dc} /* (12, 21, 13) {real, imag} */,
  {32'hbe26ae40, 32'h3edeb3c2} /* (12, 21, 12) {real, imag} */,
  {32'h3ecbbf9e, 32'hbee7477e} /* (12, 21, 11) {real, imag} */,
  {32'h3e654954, 32'hbd67e868} /* (12, 21, 10) {real, imag} */,
  {32'h3e4a8dd2, 32'hbeae6fc1} /* (12, 21, 9) {real, imag} */,
  {32'h3ed39253, 32'hbe8fdd7c} /* (12, 21, 8) {real, imag} */,
  {32'hbf6b4003, 32'h3f1f3120} /* (12, 21, 7) {real, imag} */,
  {32'h3eaba9e8, 32'hbd7bf840} /* (12, 21, 6) {real, imag} */,
  {32'h3e6d1526, 32'h3eeb689e} /* (12, 21, 5) {real, imag} */,
  {32'hbcda4168, 32'hbcb040c0} /* (12, 21, 4) {real, imag} */,
  {32'h3d645410, 32'h3dccb406} /* (12, 21, 3) {real, imag} */,
  {32'h3e5363fc, 32'hbeabe2e8} /* (12, 21, 2) {real, imag} */,
  {32'hbebfcec4, 32'h3f167562} /* (12, 21, 1) {real, imag} */,
  {32'hbf0a8386, 32'h3e3e7d22} /* (12, 21, 0) {real, imag} */,
  {32'h3e7337c8, 32'h3c9418a0} /* (12, 20, 31) {real, imag} */,
  {32'hbea66d18, 32'hbda4d354} /* (12, 20, 30) {real, imag} */,
  {32'hbda3b7c8, 32'h3ee61765} /* (12, 20, 29) {real, imag} */,
  {32'hbdea3c6c, 32'hbedf0697} /* (12, 20, 28) {real, imag} */,
  {32'hbe9436e9, 32'hbe1e677e} /* (12, 20, 27) {real, imag} */,
  {32'hbe067068, 32'h3ddb58c5} /* (12, 20, 26) {real, imag} */,
  {32'h3cc05360, 32'hbe849ec0} /* (12, 20, 25) {real, imag} */,
  {32'h3e4d632e, 32'h3c302380} /* (12, 20, 24) {real, imag} */,
  {32'h3b610580, 32'hbf2fb08a} /* (12, 20, 23) {real, imag} */,
  {32'h3f25f23c, 32'hbf0e306e} /* (12, 20, 22) {real, imag} */,
  {32'hbd270f42, 32'hbef86d17} /* (12, 20, 21) {real, imag} */,
  {32'h3f14f2aa, 32'h3e34e7f0} /* (12, 20, 20) {real, imag} */,
  {32'h3d7d2d48, 32'h3e8ac66a} /* (12, 20, 19) {real, imag} */,
  {32'h3e81f0a9, 32'hbd7db680} /* (12, 20, 18) {real, imag} */,
  {32'hbec87338, 32'h3f345976} /* (12, 20, 17) {real, imag} */,
  {32'hbd0dc800, 32'hbe9a3c52} /* (12, 20, 16) {real, imag} */,
  {32'h3c97fe48, 32'hbdac5759} /* (12, 20, 15) {real, imag} */,
  {32'hbe6eb2ab, 32'hbf1872ae} /* (12, 20, 14) {real, imag} */,
  {32'hbdad76ca, 32'hbe07159a} /* (12, 20, 13) {real, imag} */,
  {32'h3ec3922c, 32'h3eebcc95} /* (12, 20, 12) {real, imag} */,
  {32'hbe880318, 32'h3e7ef1de} /* (12, 20, 11) {real, imag} */,
  {32'hbd9d0888, 32'h3f12ca60} /* (12, 20, 10) {real, imag} */,
  {32'h3e578f7f, 32'h3e9e9134} /* (12, 20, 9) {real, imag} */,
  {32'h3de170ae, 32'hbdc57417} /* (12, 20, 8) {real, imag} */,
  {32'h3ebf21a0, 32'hbeaeb222} /* (12, 20, 7) {real, imag} */,
  {32'hbf400daa, 32'hbe9d8693} /* (12, 20, 6) {real, imag} */,
  {32'h3e9a6eef, 32'hbe8e1ac0} /* (12, 20, 5) {real, imag} */,
  {32'hbf218d62, 32'h3e985a0e} /* (12, 20, 4) {real, imag} */,
  {32'h3e11ea00, 32'h3f2198bc} /* (12, 20, 3) {real, imag} */,
  {32'hbec1bcf4, 32'h3e5708b8} /* (12, 20, 2) {real, imag} */,
  {32'hbe3e874d, 32'hbd9329a6} /* (12, 20, 1) {real, imag} */,
  {32'h3ef2f83e, 32'hbe2d0092} /* (12, 20, 0) {real, imag} */,
  {32'h3d83ccea, 32'hbdc277a7} /* (12, 19, 31) {real, imag} */,
  {32'h3e8f0c9d, 32'h3cff1520} /* (12, 19, 30) {real, imag} */,
  {32'hbe239940, 32'h3e5401b2} /* (12, 19, 29) {real, imag} */,
  {32'h3e06036e, 32'hbf4010a4} /* (12, 19, 28) {real, imag} */,
  {32'h3eb7ee46, 32'h3e470ab4} /* (12, 19, 27) {real, imag} */,
  {32'hbe5db408, 32'h3e1b1316} /* (12, 19, 26) {real, imag} */,
  {32'h3f0cfb45, 32'h3e051d0a} /* (12, 19, 25) {real, imag} */,
  {32'hbc1b0ff0, 32'h3e79c87e} /* (12, 19, 24) {real, imag} */,
  {32'hbe63249d, 32'hbb7ebee0} /* (12, 19, 23) {real, imag} */,
  {32'hbe980126, 32'h3e829b13} /* (12, 19, 22) {real, imag} */,
  {32'hbe33bc6a, 32'h3e0834a9} /* (12, 19, 21) {real, imag} */,
  {32'h3eb44d4f, 32'h3eb251eb} /* (12, 19, 20) {real, imag} */,
  {32'h3ee1cc70, 32'hbe7f0e7c} /* (12, 19, 19) {real, imag} */,
  {32'hbdbdb11c, 32'h3e9f5429} /* (12, 19, 18) {real, imag} */,
  {32'h3e9492f8, 32'h3db4e552} /* (12, 19, 17) {real, imag} */,
  {32'hbe8062f2, 32'hbc893d2c} /* (12, 19, 16) {real, imag} */,
  {32'h3d21a1d2, 32'h3db9fbc8} /* (12, 19, 15) {real, imag} */,
  {32'h3e9ab7a6, 32'hbe47ad18} /* (12, 19, 14) {real, imag} */,
  {32'h3cdbcea4, 32'h3df1e649} /* (12, 19, 13) {real, imag} */,
  {32'hbcaec320, 32'hbc63d140} /* (12, 19, 12) {real, imag} */,
  {32'hbe3f0222, 32'hbd67d49c} /* (12, 19, 11) {real, imag} */,
  {32'h3f225326, 32'hbf2d1844} /* (12, 19, 10) {real, imag} */,
  {32'hbeb814f6, 32'h3d09dc84} /* (12, 19, 9) {real, imag} */,
  {32'h3d8cd287, 32'hbe38f510} /* (12, 19, 8) {real, imag} */,
  {32'h3eaf3170, 32'h3df731c8} /* (12, 19, 7) {real, imag} */,
  {32'h3e4ea723, 32'hbd3b1a57} /* (12, 19, 6) {real, imag} */,
  {32'hbee44dd6, 32'h3f03020a} /* (12, 19, 5) {real, imag} */,
  {32'h3e4aeecc, 32'hbdcf1528} /* (12, 19, 4) {real, imag} */,
  {32'h3c6dc580, 32'hbd254666} /* (12, 19, 3) {real, imag} */,
  {32'hbe1b5811, 32'hbe34f2dd} /* (12, 19, 2) {real, imag} */,
  {32'h3e58c7cf, 32'hbe8a5177} /* (12, 19, 1) {real, imag} */,
  {32'h3d93f162, 32'hbe209a76} /* (12, 19, 0) {real, imag} */,
  {32'hbe017e78, 32'h3d5d81ce} /* (12, 18, 31) {real, imag} */,
  {32'h3e10307c, 32'hbdfd2cdc} /* (12, 18, 30) {real, imag} */,
  {32'hbe34a66b, 32'h3e2f07a3} /* (12, 18, 29) {real, imag} */,
  {32'hbebb83d0, 32'h3d0bf2ec} /* (12, 18, 28) {real, imag} */,
  {32'hbe53b863, 32'hbf332638} /* (12, 18, 27) {real, imag} */,
  {32'hbe36f300, 32'hbd83f87c} /* (12, 18, 26) {real, imag} */,
  {32'h3db1cd35, 32'h3e8b6377} /* (12, 18, 25) {real, imag} */,
  {32'hbd834c0c, 32'h3e07dcc4} /* (12, 18, 24) {real, imag} */,
  {32'hbb13c0c0, 32'hbee2cb74} /* (12, 18, 23) {real, imag} */,
  {32'hbe256c3d, 32'h3edd488a} /* (12, 18, 22) {real, imag} */,
  {32'hbed95416, 32'hbf1ad53a} /* (12, 18, 21) {real, imag} */,
  {32'h3e393705, 32'h3e8d30c8} /* (12, 18, 20) {real, imag} */,
  {32'h3e9b8c15, 32'h3f03ba70} /* (12, 18, 19) {real, imag} */,
  {32'h3e53911a, 32'hbd73eff0} /* (12, 18, 18) {real, imag} */,
  {32'h3d8f7ed8, 32'hbecdac09} /* (12, 18, 17) {real, imag} */,
  {32'h3f0acf87, 32'h3ec5cea3} /* (12, 18, 16) {real, imag} */,
  {32'hbb91f8e0, 32'h3e610868} /* (12, 18, 15) {real, imag} */,
  {32'hbcc920b4, 32'h3dc0929f} /* (12, 18, 14) {real, imag} */,
  {32'hbe416301, 32'hbef53cf4} /* (12, 18, 13) {real, imag} */,
  {32'hbe29b85a, 32'hbe3146cd} /* (12, 18, 12) {real, imag} */,
  {32'hbe7fcd52, 32'h3e21c17b} /* (12, 18, 11) {real, imag} */,
  {32'hbd1c6788, 32'hbd25a96a} /* (12, 18, 10) {real, imag} */,
  {32'h3e9e4a18, 32'h3e4a374c} /* (12, 18, 9) {real, imag} */,
  {32'h3eb7ecc2, 32'h3e9c6160} /* (12, 18, 8) {real, imag} */,
  {32'hbbf40fc0, 32'h3dd44ca6} /* (12, 18, 7) {real, imag} */,
  {32'hbe3c2b9c, 32'h3cd9e61c} /* (12, 18, 6) {real, imag} */,
  {32'hbef2c10e, 32'hbf2b7596} /* (12, 18, 5) {real, imag} */,
  {32'hbee664b1, 32'h3e7d9d26} /* (12, 18, 4) {real, imag} */,
  {32'h3d3908a6, 32'h3d84b85e} /* (12, 18, 3) {real, imag} */,
  {32'h3d9b15e6, 32'h3dc8a5b4} /* (12, 18, 2) {real, imag} */,
  {32'hbe679179, 32'hbd578598} /* (12, 18, 1) {real, imag} */,
  {32'h3d2c0611, 32'h3e9af71e} /* (12, 18, 0) {real, imag} */,
  {32'hbdedbe28, 32'hbe2f7bf5} /* (12, 17, 31) {real, imag} */,
  {32'hbecb0194, 32'h3e397bf6} /* (12, 17, 30) {real, imag} */,
  {32'h3e1c4aaa, 32'hbc6e4ce8} /* (12, 17, 29) {real, imag} */,
  {32'hbd846534, 32'hbdd6f5f3} /* (12, 17, 28) {real, imag} */,
  {32'h3cc1e67c, 32'h3e5b53d2} /* (12, 17, 27) {real, imag} */,
  {32'h3e1853fd, 32'hbf0a42a2} /* (12, 17, 26) {real, imag} */,
  {32'h3dec32e3, 32'h3e45d243} /* (12, 17, 25) {real, imag} */,
  {32'hbee62a82, 32'hbee3aed8} /* (12, 17, 24) {real, imag} */,
  {32'hbd5f34dc, 32'h3ec28782} /* (12, 17, 23) {real, imag} */,
  {32'hbdf399a7, 32'h3d5a526e} /* (12, 17, 22) {real, imag} */,
  {32'h3ed48c87, 32'h3e0daf24} /* (12, 17, 21) {real, imag} */,
  {32'h3de1c8b7, 32'hbd842c9c} /* (12, 17, 20) {real, imag} */,
  {32'hbe27082e, 32'hbe888e34} /* (12, 17, 19) {real, imag} */,
  {32'h3e03ada6, 32'hbe14c1c4} /* (12, 17, 18) {real, imag} */,
  {32'hbde0e474, 32'hbd98584e} /* (12, 17, 17) {real, imag} */,
  {32'hbe4f8362, 32'hbe654ba5} /* (12, 17, 16) {real, imag} */,
  {32'hbe761406, 32'hbd70824c} /* (12, 17, 15) {real, imag} */,
  {32'hbebb465c, 32'h3e0719aa} /* (12, 17, 14) {real, imag} */,
  {32'hbe0d21eb, 32'hbd5a4218} /* (12, 17, 13) {real, imag} */,
  {32'hbe853d36, 32'h3c9759dc} /* (12, 17, 12) {real, imag} */,
  {32'h3dc2cd1e, 32'hbdf0813e} /* (12, 17, 11) {real, imag} */,
  {32'h3ec47398, 32'h3ece63bd} /* (12, 17, 10) {real, imag} */,
  {32'hbd0f6096, 32'hbd915f1c} /* (12, 17, 9) {real, imag} */,
  {32'hbd026fa4, 32'h3e26ae6a} /* (12, 17, 8) {real, imag} */,
  {32'hbed77d76, 32'h3e590872} /* (12, 17, 7) {real, imag} */,
  {32'hbe98b0dd, 32'h3e626087} /* (12, 17, 6) {real, imag} */,
  {32'h3da1a312, 32'hbde67816} /* (12, 17, 5) {real, imag} */,
  {32'h3eb71132, 32'h3e52f912} /* (12, 17, 4) {real, imag} */,
  {32'hbe0b4282, 32'hbc2561e0} /* (12, 17, 3) {real, imag} */,
  {32'hbe25fdf8, 32'h3d241f1e} /* (12, 17, 2) {real, imag} */,
  {32'h3e1982a7, 32'hbd9742f6} /* (12, 17, 1) {real, imag} */,
  {32'h3e81092f, 32'hbe7bc172} /* (12, 17, 0) {real, imag} */,
  {32'hbe37ab8a, 32'h3dae1d4e} /* (12, 16, 31) {real, imag} */,
  {32'hbe28b886, 32'h3e34cb12} /* (12, 16, 30) {real, imag} */,
  {32'hbdff2b97, 32'h3dc1d87e} /* (12, 16, 29) {real, imag} */,
  {32'h3e0aa74e, 32'h3ec7d54a} /* (12, 16, 28) {real, imag} */,
  {32'h3dc69758, 32'h3e0a1e37} /* (12, 16, 27) {real, imag} */,
  {32'hbdfa28e6, 32'hbe0b5b4e} /* (12, 16, 26) {real, imag} */,
  {32'h3ee167c4, 32'hbbfdfec0} /* (12, 16, 25) {real, imag} */,
  {32'h3e9e6992, 32'hbdb047ef} /* (12, 16, 24) {real, imag} */,
  {32'h3e21e68a, 32'h3ed68856} /* (12, 16, 23) {real, imag} */,
  {32'hbd324c68, 32'h3e2cc2cf} /* (12, 16, 22) {real, imag} */,
  {32'hbe827a9f, 32'h3db1efa0} /* (12, 16, 21) {real, imag} */,
  {32'hbde95eae, 32'hbdbdf524} /* (12, 16, 20) {real, imag} */,
  {32'h3ccc5ba0, 32'hbd9d366b} /* (12, 16, 19) {real, imag} */,
  {32'h3ec18d42, 32'h3d0e0240} /* (12, 16, 18) {real, imag} */,
  {32'h3ef2caaa, 32'h3dc92da0} /* (12, 16, 17) {real, imag} */,
  {32'h3e096b48, 32'h00000000} /* (12, 16, 16) {real, imag} */,
  {32'h3ef2caaa, 32'hbdc92da0} /* (12, 16, 15) {real, imag} */,
  {32'h3ec18d42, 32'hbd0e0240} /* (12, 16, 14) {real, imag} */,
  {32'h3ccc5ba0, 32'h3d9d366b} /* (12, 16, 13) {real, imag} */,
  {32'hbde95eae, 32'h3dbdf524} /* (12, 16, 12) {real, imag} */,
  {32'hbe827a9f, 32'hbdb1efa0} /* (12, 16, 11) {real, imag} */,
  {32'hbd324c68, 32'hbe2cc2cf} /* (12, 16, 10) {real, imag} */,
  {32'h3e21e68a, 32'hbed68856} /* (12, 16, 9) {real, imag} */,
  {32'h3e9e6992, 32'h3db047ef} /* (12, 16, 8) {real, imag} */,
  {32'h3ee167c4, 32'h3bfdfec0} /* (12, 16, 7) {real, imag} */,
  {32'hbdfa28e6, 32'h3e0b5b4e} /* (12, 16, 6) {real, imag} */,
  {32'h3dc69758, 32'hbe0a1e37} /* (12, 16, 5) {real, imag} */,
  {32'h3e0aa74e, 32'hbec7d54a} /* (12, 16, 4) {real, imag} */,
  {32'hbdff2b97, 32'hbdc1d87e} /* (12, 16, 3) {real, imag} */,
  {32'hbe28b886, 32'hbe34cb12} /* (12, 16, 2) {real, imag} */,
  {32'hbe37ab8a, 32'hbdae1d4e} /* (12, 16, 1) {real, imag} */,
  {32'h3e5392c0, 32'h00000000} /* (12, 16, 0) {real, imag} */,
  {32'h3e1982a7, 32'h3d9742f6} /* (12, 15, 31) {real, imag} */,
  {32'hbe25fdf8, 32'hbd241f1e} /* (12, 15, 30) {real, imag} */,
  {32'hbe0b4282, 32'h3c2561e0} /* (12, 15, 29) {real, imag} */,
  {32'h3eb71132, 32'hbe52f912} /* (12, 15, 28) {real, imag} */,
  {32'h3da1a312, 32'h3de67816} /* (12, 15, 27) {real, imag} */,
  {32'hbe98b0dd, 32'hbe626087} /* (12, 15, 26) {real, imag} */,
  {32'hbed77d76, 32'hbe590872} /* (12, 15, 25) {real, imag} */,
  {32'hbd026fa4, 32'hbe26ae6a} /* (12, 15, 24) {real, imag} */,
  {32'hbd0f6096, 32'h3d915f1c} /* (12, 15, 23) {real, imag} */,
  {32'h3ec47398, 32'hbece63bd} /* (12, 15, 22) {real, imag} */,
  {32'h3dc2cd1e, 32'h3df0813e} /* (12, 15, 21) {real, imag} */,
  {32'hbe853d36, 32'hbc9759dc} /* (12, 15, 20) {real, imag} */,
  {32'hbe0d21eb, 32'h3d5a4218} /* (12, 15, 19) {real, imag} */,
  {32'hbebb465c, 32'hbe0719aa} /* (12, 15, 18) {real, imag} */,
  {32'hbe761406, 32'h3d70824c} /* (12, 15, 17) {real, imag} */,
  {32'hbe4f8362, 32'h3e654ba5} /* (12, 15, 16) {real, imag} */,
  {32'hbde0e474, 32'h3d98584e} /* (12, 15, 15) {real, imag} */,
  {32'h3e03ada6, 32'h3e14c1c4} /* (12, 15, 14) {real, imag} */,
  {32'hbe27082e, 32'h3e888e34} /* (12, 15, 13) {real, imag} */,
  {32'h3de1c8b7, 32'h3d842c9c} /* (12, 15, 12) {real, imag} */,
  {32'h3ed48c87, 32'hbe0daf24} /* (12, 15, 11) {real, imag} */,
  {32'hbdf399a7, 32'hbd5a526e} /* (12, 15, 10) {real, imag} */,
  {32'hbd5f34dc, 32'hbec28782} /* (12, 15, 9) {real, imag} */,
  {32'hbee62a82, 32'h3ee3aed8} /* (12, 15, 8) {real, imag} */,
  {32'h3dec32e3, 32'hbe45d243} /* (12, 15, 7) {real, imag} */,
  {32'h3e1853fd, 32'h3f0a42a2} /* (12, 15, 6) {real, imag} */,
  {32'h3cc1e67c, 32'hbe5b53d2} /* (12, 15, 5) {real, imag} */,
  {32'hbd846534, 32'h3dd6f5f3} /* (12, 15, 4) {real, imag} */,
  {32'h3e1c4aaa, 32'h3c6e4ce8} /* (12, 15, 3) {real, imag} */,
  {32'hbecb0194, 32'hbe397bf6} /* (12, 15, 2) {real, imag} */,
  {32'hbdedbe28, 32'h3e2f7bf5} /* (12, 15, 1) {real, imag} */,
  {32'h3e81092f, 32'h3e7bc172} /* (12, 15, 0) {real, imag} */,
  {32'hbe679179, 32'h3d578598} /* (12, 14, 31) {real, imag} */,
  {32'h3d9b15e6, 32'hbdc8a5b4} /* (12, 14, 30) {real, imag} */,
  {32'h3d3908a6, 32'hbd84b85e} /* (12, 14, 29) {real, imag} */,
  {32'hbee664b1, 32'hbe7d9d26} /* (12, 14, 28) {real, imag} */,
  {32'hbef2c10e, 32'h3f2b7596} /* (12, 14, 27) {real, imag} */,
  {32'hbe3c2b9c, 32'hbcd9e61c} /* (12, 14, 26) {real, imag} */,
  {32'hbbf40fc0, 32'hbdd44ca6} /* (12, 14, 25) {real, imag} */,
  {32'h3eb7ecc2, 32'hbe9c6160} /* (12, 14, 24) {real, imag} */,
  {32'h3e9e4a18, 32'hbe4a374c} /* (12, 14, 23) {real, imag} */,
  {32'hbd1c6788, 32'h3d25a96a} /* (12, 14, 22) {real, imag} */,
  {32'hbe7fcd52, 32'hbe21c17b} /* (12, 14, 21) {real, imag} */,
  {32'hbe29b85a, 32'h3e3146cd} /* (12, 14, 20) {real, imag} */,
  {32'hbe416301, 32'h3ef53cf4} /* (12, 14, 19) {real, imag} */,
  {32'hbcc920b4, 32'hbdc0929f} /* (12, 14, 18) {real, imag} */,
  {32'hbb91f8e0, 32'hbe610868} /* (12, 14, 17) {real, imag} */,
  {32'h3f0acf87, 32'hbec5cea3} /* (12, 14, 16) {real, imag} */,
  {32'h3d8f7ed8, 32'h3ecdac09} /* (12, 14, 15) {real, imag} */,
  {32'h3e53911a, 32'h3d73eff0} /* (12, 14, 14) {real, imag} */,
  {32'h3e9b8c15, 32'hbf03ba70} /* (12, 14, 13) {real, imag} */,
  {32'h3e393705, 32'hbe8d30c8} /* (12, 14, 12) {real, imag} */,
  {32'hbed95416, 32'h3f1ad53a} /* (12, 14, 11) {real, imag} */,
  {32'hbe256c3d, 32'hbedd488a} /* (12, 14, 10) {real, imag} */,
  {32'hbb13c0c0, 32'h3ee2cb74} /* (12, 14, 9) {real, imag} */,
  {32'hbd834c0c, 32'hbe07dcc4} /* (12, 14, 8) {real, imag} */,
  {32'h3db1cd35, 32'hbe8b6377} /* (12, 14, 7) {real, imag} */,
  {32'hbe36f300, 32'h3d83f87c} /* (12, 14, 6) {real, imag} */,
  {32'hbe53b863, 32'h3f332638} /* (12, 14, 5) {real, imag} */,
  {32'hbebb83d0, 32'hbd0bf2ec} /* (12, 14, 4) {real, imag} */,
  {32'hbe34a66b, 32'hbe2f07a3} /* (12, 14, 3) {real, imag} */,
  {32'h3e10307c, 32'h3dfd2cdc} /* (12, 14, 2) {real, imag} */,
  {32'hbe017e78, 32'hbd5d81ce} /* (12, 14, 1) {real, imag} */,
  {32'h3d2c0611, 32'hbe9af71e} /* (12, 14, 0) {real, imag} */,
  {32'h3e58c7cf, 32'h3e8a5177} /* (12, 13, 31) {real, imag} */,
  {32'hbe1b5811, 32'h3e34f2dd} /* (12, 13, 30) {real, imag} */,
  {32'h3c6dc580, 32'h3d254666} /* (12, 13, 29) {real, imag} */,
  {32'h3e4aeecc, 32'h3dcf1528} /* (12, 13, 28) {real, imag} */,
  {32'hbee44dd6, 32'hbf03020a} /* (12, 13, 27) {real, imag} */,
  {32'h3e4ea723, 32'h3d3b1a57} /* (12, 13, 26) {real, imag} */,
  {32'h3eaf3170, 32'hbdf731c8} /* (12, 13, 25) {real, imag} */,
  {32'h3d8cd287, 32'h3e38f510} /* (12, 13, 24) {real, imag} */,
  {32'hbeb814f6, 32'hbd09dc84} /* (12, 13, 23) {real, imag} */,
  {32'h3f225326, 32'h3f2d1844} /* (12, 13, 22) {real, imag} */,
  {32'hbe3f0222, 32'h3d67d49c} /* (12, 13, 21) {real, imag} */,
  {32'hbcaec320, 32'h3c63d140} /* (12, 13, 20) {real, imag} */,
  {32'h3cdbcea4, 32'hbdf1e649} /* (12, 13, 19) {real, imag} */,
  {32'h3e9ab7a6, 32'h3e47ad18} /* (12, 13, 18) {real, imag} */,
  {32'h3d21a1d2, 32'hbdb9fbc8} /* (12, 13, 17) {real, imag} */,
  {32'hbe8062f2, 32'h3c893d2c} /* (12, 13, 16) {real, imag} */,
  {32'h3e9492f8, 32'hbdb4e552} /* (12, 13, 15) {real, imag} */,
  {32'hbdbdb11c, 32'hbe9f5429} /* (12, 13, 14) {real, imag} */,
  {32'h3ee1cc70, 32'h3e7f0e7c} /* (12, 13, 13) {real, imag} */,
  {32'h3eb44d4f, 32'hbeb251eb} /* (12, 13, 12) {real, imag} */,
  {32'hbe33bc6a, 32'hbe0834a9} /* (12, 13, 11) {real, imag} */,
  {32'hbe980126, 32'hbe829b13} /* (12, 13, 10) {real, imag} */,
  {32'hbe63249d, 32'h3b7ebee0} /* (12, 13, 9) {real, imag} */,
  {32'hbc1b0ff0, 32'hbe79c87e} /* (12, 13, 8) {real, imag} */,
  {32'h3f0cfb45, 32'hbe051d0a} /* (12, 13, 7) {real, imag} */,
  {32'hbe5db408, 32'hbe1b1316} /* (12, 13, 6) {real, imag} */,
  {32'h3eb7ee46, 32'hbe470ab4} /* (12, 13, 5) {real, imag} */,
  {32'h3e06036e, 32'h3f4010a4} /* (12, 13, 4) {real, imag} */,
  {32'hbe239940, 32'hbe5401b2} /* (12, 13, 3) {real, imag} */,
  {32'h3e8f0c9d, 32'hbcff1520} /* (12, 13, 2) {real, imag} */,
  {32'h3d83ccea, 32'h3dc277a7} /* (12, 13, 1) {real, imag} */,
  {32'h3d93f162, 32'h3e209a76} /* (12, 13, 0) {real, imag} */,
  {32'hbe3e874d, 32'h3d9329a6} /* (12, 12, 31) {real, imag} */,
  {32'hbec1bcf4, 32'hbe5708b8} /* (12, 12, 30) {real, imag} */,
  {32'h3e11ea00, 32'hbf2198bc} /* (12, 12, 29) {real, imag} */,
  {32'hbf218d62, 32'hbe985a0e} /* (12, 12, 28) {real, imag} */,
  {32'h3e9a6eef, 32'h3e8e1ac0} /* (12, 12, 27) {real, imag} */,
  {32'hbf400daa, 32'h3e9d8693} /* (12, 12, 26) {real, imag} */,
  {32'h3ebf21a0, 32'h3eaeb222} /* (12, 12, 25) {real, imag} */,
  {32'h3de170ae, 32'h3dc57417} /* (12, 12, 24) {real, imag} */,
  {32'h3e578f7f, 32'hbe9e9134} /* (12, 12, 23) {real, imag} */,
  {32'hbd9d0888, 32'hbf12ca60} /* (12, 12, 22) {real, imag} */,
  {32'hbe880318, 32'hbe7ef1de} /* (12, 12, 21) {real, imag} */,
  {32'h3ec3922c, 32'hbeebcc95} /* (12, 12, 20) {real, imag} */,
  {32'hbdad76ca, 32'h3e07159a} /* (12, 12, 19) {real, imag} */,
  {32'hbe6eb2ab, 32'h3f1872ae} /* (12, 12, 18) {real, imag} */,
  {32'h3c97fe48, 32'h3dac5759} /* (12, 12, 17) {real, imag} */,
  {32'hbd0dc800, 32'h3e9a3c52} /* (12, 12, 16) {real, imag} */,
  {32'hbec87338, 32'hbf345976} /* (12, 12, 15) {real, imag} */,
  {32'h3e81f0a9, 32'h3d7db680} /* (12, 12, 14) {real, imag} */,
  {32'h3d7d2d48, 32'hbe8ac66a} /* (12, 12, 13) {real, imag} */,
  {32'h3f14f2aa, 32'hbe34e7f0} /* (12, 12, 12) {real, imag} */,
  {32'hbd270f42, 32'h3ef86d17} /* (12, 12, 11) {real, imag} */,
  {32'h3f25f23c, 32'h3f0e306e} /* (12, 12, 10) {real, imag} */,
  {32'h3b610580, 32'h3f2fb08a} /* (12, 12, 9) {real, imag} */,
  {32'h3e4d632e, 32'hbc302380} /* (12, 12, 8) {real, imag} */,
  {32'h3cc05360, 32'h3e849ec0} /* (12, 12, 7) {real, imag} */,
  {32'hbe067068, 32'hbddb58c5} /* (12, 12, 6) {real, imag} */,
  {32'hbe9436e9, 32'h3e1e677e} /* (12, 12, 5) {real, imag} */,
  {32'hbdea3c6c, 32'h3edf0697} /* (12, 12, 4) {real, imag} */,
  {32'hbda3b7c8, 32'hbee61765} /* (12, 12, 3) {real, imag} */,
  {32'hbea66d18, 32'h3da4d354} /* (12, 12, 2) {real, imag} */,
  {32'h3e7337c8, 32'hbc9418a0} /* (12, 12, 1) {real, imag} */,
  {32'h3ef2f83e, 32'h3e2d0092} /* (12, 12, 0) {real, imag} */,
  {32'hbebfcec4, 32'hbf167562} /* (12, 11, 31) {real, imag} */,
  {32'h3e5363fc, 32'h3eabe2e8} /* (12, 11, 30) {real, imag} */,
  {32'h3d645410, 32'hbdccb406} /* (12, 11, 29) {real, imag} */,
  {32'hbcda4168, 32'h3cb040c0} /* (12, 11, 28) {real, imag} */,
  {32'h3e6d1526, 32'hbeeb689e} /* (12, 11, 27) {real, imag} */,
  {32'h3eaba9e8, 32'h3d7bf840} /* (12, 11, 26) {real, imag} */,
  {32'hbf6b4003, 32'hbf1f3120} /* (12, 11, 25) {real, imag} */,
  {32'h3ed39253, 32'h3e8fdd7c} /* (12, 11, 24) {real, imag} */,
  {32'h3e4a8dd2, 32'h3eae6fc1} /* (12, 11, 23) {real, imag} */,
  {32'h3e654954, 32'h3d67e868} /* (12, 11, 22) {real, imag} */,
  {32'h3ecbbf9e, 32'h3ee7477e} /* (12, 11, 21) {real, imag} */,
  {32'hbe26ae40, 32'hbedeb3c2} /* (12, 11, 20) {real, imag} */,
  {32'h3f4734fa, 32'h3ccd33dc} /* (12, 11, 19) {real, imag} */,
  {32'hbec86a28, 32'hbd417662} /* (12, 11, 18) {real, imag} */,
  {32'h3e7092f5, 32'h3e909226} /* (12, 11, 17) {real, imag} */,
  {32'hbed5b970, 32'hbe4bf572} /* (12, 11, 16) {real, imag} */,
  {32'hbe5f6904, 32'hbe0f6480} /* (12, 11, 15) {real, imag} */,
  {32'hbdfaa75d, 32'hbebde7ae} /* (12, 11, 14) {real, imag} */,
  {32'h3ddeaaac, 32'hbe133988} /* (12, 11, 13) {real, imag} */,
  {32'hbeb219e8, 32'hbd92b9ce} /* (12, 11, 12) {real, imag} */,
  {32'hbcdc20a8, 32'h3ee69013} /* (12, 11, 11) {real, imag} */,
  {32'h3c0c34a0, 32'h3e53f7b6} /* (12, 11, 10) {real, imag} */,
  {32'hbcaf3f30, 32'hbf04f9f2} /* (12, 11, 9) {real, imag} */,
  {32'hbd0f15a0, 32'h3d021db8} /* (12, 11, 8) {real, imag} */,
  {32'h3e228a16, 32'h3e5698ec} /* (12, 11, 7) {real, imag} */,
  {32'hbdfd1fda, 32'hbf052fba} /* (12, 11, 6) {real, imag} */,
  {32'hbe5ecbde, 32'h3ebb6016} /* (12, 11, 5) {real, imag} */,
  {32'h3d026e04, 32'h3cbce460} /* (12, 11, 4) {real, imag} */,
  {32'h3f4c6d1a, 32'hbe2fa69c} /* (12, 11, 3) {real, imag} */,
  {32'hbedf6022, 32'h3e0e3276} /* (12, 11, 2) {real, imag} */,
  {32'hbf834f73, 32'hbf03b45a} /* (12, 11, 1) {real, imag} */,
  {32'hbf0a8386, 32'hbe3e7d22} /* (12, 11, 0) {real, imag} */,
  {32'h3dcabc3a, 32'h3efacf8d} /* (12, 10, 31) {real, imag} */,
  {32'hbe08eda4, 32'h3973f800} /* (12, 10, 30) {real, imag} */,
  {32'hbe626c69, 32'hbe732102} /* (12, 10, 29) {real, imag} */,
  {32'h3e07cbfa, 32'h3e0c8678} /* (12, 10, 28) {real, imag} */,
  {32'hbedde302, 32'h3ea06066} /* (12, 10, 27) {real, imag} */,
  {32'h3dc1c780, 32'hbeddd260} /* (12, 10, 26) {real, imag} */,
  {32'hbf039a38, 32'h3dfccb74} /* (12, 10, 25) {real, imag} */,
  {32'h3efc55c3, 32'hbefc540c} /* (12, 10, 24) {real, imag} */,
  {32'hbf2078e2, 32'h3eef731e} /* (12, 10, 23) {real, imag} */,
  {32'h3e9a7328, 32'h3cd635a8} /* (12, 10, 22) {real, imag} */,
  {32'h3ecfaca5, 32'hbed87aac} /* (12, 10, 21) {real, imag} */,
  {32'h3d206ae4, 32'hbd9c2027} /* (12, 10, 20) {real, imag} */,
  {32'h3ebb9b44, 32'hbe34e42a} /* (12, 10, 19) {real, imag} */,
  {32'hbccae3b0, 32'h3e8ad5ee} /* (12, 10, 18) {real, imag} */,
  {32'hbdc4ab12, 32'hbe0a335e} /* (12, 10, 17) {real, imag} */,
  {32'hbeec8e7e, 32'h3dfc09dd} /* (12, 10, 16) {real, imag} */,
  {32'h3e851009, 32'h3eba4702} /* (12, 10, 15) {real, imag} */,
  {32'h3ca27404, 32'hbd2d560c} /* (12, 10, 14) {real, imag} */,
  {32'h3de6aef2, 32'hbeaf487a} /* (12, 10, 13) {real, imag} */,
  {32'hbe2d19d0, 32'hbee55c6c} /* (12, 10, 12) {real, imag} */,
  {32'h3d7092a0, 32'hbe7888d9} /* (12, 10, 11) {real, imag} */,
  {32'hbee3e382, 32'h3e8fcf0f} /* (12, 10, 10) {real, imag} */,
  {32'h3e13d84c, 32'hbd948162} /* (12, 10, 9) {real, imag} */,
  {32'hbd582168, 32'hbe015e4e} /* (12, 10, 8) {real, imag} */,
  {32'h3e86ba6c, 32'h3ef8915e} /* (12, 10, 7) {real, imag} */,
  {32'h3da65c2a, 32'hbf002e80} /* (12, 10, 6) {real, imag} */,
  {32'h3f12f1d9, 32'hbf0ec082} /* (12, 10, 5) {real, imag} */,
  {32'hbeab3b36, 32'h3f3e0441} /* (12, 10, 4) {real, imag} */,
  {32'h3dd5a988, 32'hbd24b378} /* (12, 10, 3) {real, imag} */,
  {32'hbe2b7df5, 32'hbf516798} /* (12, 10, 2) {real, imag} */,
  {32'h3dfe1902, 32'h3e5c5910} /* (12, 10, 1) {real, imag} */,
  {32'hbd4dcbf4, 32'hbd97835a} /* (12, 10, 0) {real, imag} */,
  {32'hbf2c26a2, 32'h3ed81372} /* (12, 9, 31) {real, imag} */,
  {32'h3e7139b0, 32'hbe0ba34c} /* (12, 9, 30) {real, imag} */,
  {32'h3defb2a9, 32'hbe75a3de} /* (12, 9, 29) {real, imag} */,
  {32'h3e130aa4, 32'hbe9f0be6} /* (12, 9, 28) {real, imag} */,
  {32'hbedfdec0, 32'h3e1180ca} /* (12, 9, 27) {real, imag} */,
  {32'hbd91b4d8, 32'h3d976184} /* (12, 9, 26) {real, imag} */,
  {32'hbe8bfbea, 32'hbe309ac7} /* (12, 9, 25) {real, imag} */,
  {32'hbf69029f, 32'hbdf3fe1a} /* (12, 9, 24) {real, imag} */,
  {32'h3de7e15b, 32'h3ec4c022} /* (12, 9, 23) {real, imag} */,
  {32'h3dc731f8, 32'hbe452e51} /* (12, 9, 22) {real, imag} */,
  {32'hbe54d71b, 32'h3dde34ba} /* (12, 9, 21) {real, imag} */,
  {32'h3e2cd43c, 32'h3c888848} /* (12, 9, 20) {real, imag} */,
  {32'h3eeb7e76, 32'h3dd0ba5d} /* (12, 9, 19) {real, imag} */,
  {32'h3dabe536, 32'hbe16da72} /* (12, 9, 18) {real, imag} */,
  {32'h3de2ee80, 32'h3e56a21a} /* (12, 9, 17) {real, imag} */,
  {32'hbc959970, 32'h3e48ca82} /* (12, 9, 16) {real, imag} */,
  {32'h3dcf1389, 32'h3b737140} /* (12, 9, 15) {real, imag} */,
  {32'h3e2feba0, 32'hbe01e7d2} /* (12, 9, 14) {real, imag} */,
  {32'hbec508e0, 32'h3e8603a0} /* (12, 9, 13) {real, imag} */,
  {32'hbe85bdbf, 32'hbe426312} /* (12, 9, 12) {real, imag} */,
  {32'hbefee0a2, 32'hbd647501} /* (12, 9, 11) {real, imag} */,
  {32'hbec4eb94, 32'hbe904fb8} /* (12, 9, 10) {real, imag} */,
  {32'h3f28d9da, 32'hbe01fdc0} /* (12, 9, 9) {real, imag} */,
  {32'hbd48f9b8, 32'hbe0550f6} /* (12, 9, 8) {real, imag} */,
  {32'h3eb47e58, 32'h3e810b1f} /* (12, 9, 7) {real, imag} */,
  {32'hbf0d0231, 32'h3ed6ed2e} /* (12, 9, 6) {real, imag} */,
  {32'hbe8e991e, 32'h3eec5cd1} /* (12, 9, 5) {real, imag} */,
  {32'hbea3440a, 32'h3e8694be} /* (12, 9, 4) {real, imag} */,
  {32'h3f14694d, 32'hbf273b66} /* (12, 9, 3) {real, imag} */,
  {32'hbeb2cf29, 32'hbec50dc2} /* (12, 9, 2) {real, imag} */,
  {32'h3f8c88e0, 32'h3efba136} /* (12, 9, 1) {real, imag} */,
  {32'hbe5846d4, 32'hbeb62a85} /* (12, 9, 0) {real, imag} */,
  {32'hbfb68768, 32'hbf43492a} /* (12, 8, 31) {real, imag} */,
  {32'h3f67b91d, 32'h3ecf02ca} /* (12, 8, 30) {real, imag} */,
  {32'h3dbe2a16, 32'hbefd3084} /* (12, 8, 29) {real, imag} */,
  {32'h3e89fe48, 32'hbf00a829} /* (12, 8, 28) {real, imag} */,
  {32'h3f2c1f4b, 32'hbe9a1a5d} /* (12, 8, 27) {real, imag} */,
  {32'h3dd7b212, 32'h3e989799} /* (12, 8, 26) {real, imag} */,
  {32'h3d3b2a06, 32'hbeaa99d8} /* (12, 8, 25) {real, imag} */,
  {32'h3da65bd6, 32'h3e94c569} /* (12, 8, 24) {real, imag} */,
  {32'h3d4af790, 32'hbe9e647d} /* (12, 8, 23) {real, imag} */,
  {32'hbecc24f9, 32'h3f0b88c2} /* (12, 8, 22) {real, imag} */,
  {32'h3f0af3dd, 32'hbb8b2610} /* (12, 8, 21) {real, imag} */,
  {32'h3f043314, 32'hbe40ca62} /* (12, 8, 20) {real, imag} */,
  {32'hbee02cc6, 32'hbe8ace42} /* (12, 8, 19) {real, imag} */,
  {32'h3f05b8f0, 32'h3d229cb2} /* (12, 8, 18) {real, imag} */,
  {32'h3e755ed6, 32'hbe045e9e} /* (12, 8, 17) {real, imag} */,
  {32'h3e0bee82, 32'hbe032daf} /* (12, 8, 16) {real, imag} */,
  {32'h3df2397a, 32'h3ed0a0ba} /* (12, 8, 15) {real, imag} */,
  {32'hbe890ca4, 32'hbebd1332} /* (12, 8, 14) {real, imag} */,
  {32'hbf5fd550, 32'h3f02e46c} /* (12, 8, 13) {real, imag} */,
  {32'h3ea14265, 32'h3f70923e} /* (12, 8, 12) {real, imag} */,
  {32'h3e0d3d5d, 32'hbf11cd84} /* (12, 8, 11) {real, imag} */,
  {32'h3f18462c, 32'h3dd75580} /* (12, 8, 10) {real, imag} */,
  {32'h3df7b3d4, 32'h3d032c72} /* (12, 8, 9) {real, imag} */,
  {32'h3ea96b24, 32'hbda807c6} /* (12, 8, 8) {real, imag} */,
  {32'hbf102ce7, 32'hbd294934} /* (12, 8, 7) {real, imag} */,
  {32'h3ebbce2b, 32'hbeefa4ac} /* (12, 8, 6) {real, imag} */,
  {32'h3f38f709, 32'hbe925a6d} /* (12, 8, 5) {real, imag} */,
  {32'hbf7e4fbb, 32'hbf81c3e9} /* (12, 8, 4) {real, imag} */,
  {32'hbe4c5146, 32'h3e52beb6} /* (12, 8, 3) {real, imag} */,
  {32'h3e9f72d3, 32'h3f1c418b} /* (12, 8, 2) {real, imag} */,
  {32'hbfa71c54, 32'h3db36e38} /* (12, 8, 1) {real, imag} */,
  {32'hbf218586, 32'hbf659562} /* (12, 8, 0) {real, imag} */,
  {32'h3f0864b8, 32'hbf06813c} /* (12, 7, 31) {real, imag} */,
  {32'h3d8ba543, 32'hbf283cd6} /* (12, 7, 30) {real, imag} */,
  {32'hbe266d90, 32'h3d9902ab} /* (12, 7, 29) {real, imag} */,
  {32'hbbf71ae0, 32'h3e80fbe1} /* (12, 7, 28) {real, imag} */,
  {32'hbd8de3ca, 32'hbed9da9e} /* (12, 7, 27) {real, imag} */,
  {32'h3d58d4d9, 32'h3e94ef5a} /* (12, 7, 26) {real, imag} */,
  {32'h3f0e6da7, 32'h3f00ff3c} /* (12, 7, 25) {real, imag} */,
  {32'hbe469ca6, 32'hbeeda232} /* (12, 7, 24) {real, imag} */,
  {32'hbee8ce72, 32'hbe6cdbfa} /* (12, 7, 23) {real, imag} */,
  {32'hbdc94967, 32'h3f1576f0} /* (12, 7, 22) {real, imag} */,
  {32'h3f31bf63, 32'hbeb0db68} /* (12, 7, 21) {real, imag} */,
  {32'h3e4ba3a8, 32'h3e8a611a} /* (12, 7, 20) {real, imag} */,
  {32'hbe5b93a7, 32'h3e540646} /* (12, 7, 19) {real, imag} */,
  {32'h3cb9c740, 32'h3e503f0a} /* (12, 7, 18) {real, imag} */,
  {32'hbe3aef45, 32'h3e87c313} /* (12, 7, 17) {real, imag} */,
  {32'hbeba4e07, 32'h3e9ec426} /* (12, 7, 16) {real, imag} */,
  {32'h3e995c5a, 32'hbdda43c5} /* (12, 7, 15) {real, imag} */,
  {32'hbe3fcbee, 32'hbd0a4222} /* (12, 7, 14) {real, imag} */,
  {32'hbd4ee135, 32'hbf209ca0} /* (12, 7, 13) {real, imag} */,
  {32'h3df6e958, 32'hbd6a1e50} /* (12, 7, 12) {real, imag} */,
  {32'h3f46678c, 32'hbe89de8a} /* (12, 7, 11) {real, imag} */,
  {32'h3eb7f084, 32'h3e4eae74} /* (12, 7, 10) {real, imag} */,
  {32'hbea9ec26, 32'hbe902867} /* (12, 7, 9) {real, imag} */,
  {32'h3eb73284, 32'hbdc92c72} /* (12, 7, 8) {real, imag} */,
  {32'hbe6e6d63, 32'h3d7c670f} /* (12, 7, 7) {real, imag} */,
  {32'h3e8e4e3f, 32'hbc5027e0} /* (12, 7, 6) {real, imag} */,
  {32'hbb904e60, 32'h3e6dab12} /* (12, 7, 5) {real, imag} */,
  {32'hbe89305b, 32'h3f435708} /* (12, 7, 4) {real, imag} */,
  {32'hbf2baeea, 32'h3f219736} /* (12, 7, 3) {real, imag} */,
  {32'hbeaad936, 32'hbe8de49f} /* (12, 7, 2) {real, imag} */,
  {32'h3f32866c, 32'h3f1a62ae} /* (12, 7, 1) {real, imag} */,
  {32'h3d0a5948, 32'h3e9dbf1c} /* (12, 7, 0) {real, imag} */,
  {32'h3ec8d60a, 32'hbf09383b} /* (12, 6, 31) {real, imag} */,
  {32'h3f870773, 32'hbdadedc6} /* (12, 6, 30) {real, imag} */,
  {32'h3ef0c5af, 32'hbf0cd5b2} /* (12, 6, 29) {real, imag} */,
  {32'hbe2373d8, 32'hbf0ec897} /* (12, 6, 28) {real, imag} */,
  {32'hbdcd6dd6, 32'h3ef7188a} /* (12, 6, 27) {real, imag} */,
  {32'hbcd27f58, 32'h3e8adc55} /* (12, 6, 26) {real, imag} */,
  {32'h3d15db3c, 32'hbe7a869f} /* (12, 6, 25) {real, imag} */,
  {32'hbeac8ba4, 32'h3e2e2e86} /* (12, 6, 24) {real, imag} */,
  {32'hbcadade8, 32'hbe11acab} /* (12, 6, 23) {real, imag} */,
  {32'h3f56f712, 32'hbeb0ef90} /* (12, 6, 22) {real, imag} */,
  {32'h3d759cd4, 32'hbdc98209} /* (12, 6, 21) {real, imag} */,
  {32'h3e825b10, 32'hbd5da844} /* (12, 6, 20) {real, imag} */,
  {32'h3ec5368a, 32'h3ee748ca} /* (12, 6, 19) {real, imag} */,
  {32'hbea77344, 32'hbd978d2d} /* (12, 6, 18) {real, imag} */,
  {32'h3e780efa, 32'hbe906fff} /* (12, 6, 17) {real, imag} */,
  {32'hbe78fa08, 32'h3df247e3} /* (12, 6, 16) {real, imag} */,
  {32'h3da93c3f, 32'hbcce4a20} /* (12, 6, 15) {real, imag} */,
  {32'h3e95d21d, 32'hbec410c2} /* (12, 6, 14) {real, imag} */,
  {32'hbe37ac2e, 32'h3e4b43c5} /* (12, 6, 13) {real, imag} */,
  {32'hbd579764, 32'h3e2b156b} /* (12, 6, 12) {real, imag} */,
  {32'hbda2c197, 32'h3c95855c} /* (12, 6, 11) {real, imag} */,
  {32'hbf14698a, 32'hbec35a5e} /* (12, 6, 10) {real, imag} */,
  {32'hbf71ccb5, 32'hbda0763e} /* (12, 6, 9) {real, imag} */,
  {32'h3e76e78d, 32'hbe9d95cf} /* (12, 6, 8) {real, imag} */,
  {32'hbea09ccd, 32'h3e43c6fc} /* (12, 6, 7) {real, imag} */,
  {32'h3d0748fe, 32'hbf0dff78} /* (12, 6, 6) {real, imag} */,
  {32'h3eec1961, 32'hbf6b224e} /* (12, 6, 5) {real, imag} */,
  {32'h3ea76cbc, 32'hbf06d6ae} /* (12, 6, 4) {real, imag} */,
  {32'hbd5a4105, 32'h3ed058cc} /* (12, 6, 3) {real, imag} */,
  {32'h3e621dd1, 32'hbe282dc7} /* (12, 6, 2) {real, imag} */,
  {32'h3f40688c, 32'hbea56c48} /* (12, 6, 1) {real, imag} */,
  {32'h3e579f30, 32'h3f092917} /* (12, 6, 0) {real, imag} */,
  {32'hc05779ce, 32'hbf01bdaa} /* (12, 5, 31) {real, imag} */,
  {32'h3f20296b, 32'h3ec39b3d} /* (12, 5, 30) {real, imag} */,
  {32'hbdd46108, 32'h3bf14600} /* (12, 5, 29) {real, imag} */,
  {32'hbedd801a, 32'h3f9fcc3e} /* (12, 5, 28) {real, imag} */,
  {32'h3ebd4f8e, 32'h3f5b9038} /* (12, 5, 27) {real, imag} */,
  {32'hbe0a0898, 32'hbdc530d6} /* (12, 5, 26) {real, imag} */,
  {32'h3e91643e, 32'hbefbe684} /* (12, 5, 25) {real, imag} */,
  {32'h3ee46d1a, 32'hbf214e6a} /* (12, 5, 24) {real, imag} */,
  {32'h3ebbef24, 32'hbda990b2} /* (12, 5, 23) {real, imag} */,
  {32'h3eb6a4df, 32'hbe4e5ece} /* (12, 5, 22) {real, imag} */,
  {32'h3f15e960, 32'hbd63c09e} /* (12, 5, 21) {real, imag} */,
  {32'h3e219a58, 32'hbdebb680} /* (12, 5, 20) {real, imag} */,
  {32'hbdc710e5, 32'h3f3bc358} /* (12, 5, 19) {real, imag} */,
  {32'hbe8e6636, 32'hbdcb7434} /* (12, 5, 18) {real, imag} */,
  {32'h3dba5002, 32'hbe7f7cd6} /* (12, 5, 17) {real, imag} */,
  {32'h3e7af88e, 32'h3ba99bc0} /* (12, 5, 16) {real, imag} */,
  {32'h3d896b4e, 32'h3d323a2e} /* (12, 5, 15) {real, imag} */,
  {32'hbf27de4e, 32'h3e52b6f0} /* (12, 5, 14) {real, imag} */,
  {32'hbe6751e9, 32'h3e634ba0} /* (12, 5, 13) {real, imag} */,
  {32'h3ee46224, 32'hbd2a26f8} /* (12, 5, 12) {real, imag} */,
  {32'h3e6f5cb0, 32'h3ebb6d1c} /* (12, 5, 11) {real, imag} */,
  {32'hbe9a86c0, 32'h3ecbbc92} /* (12, 5, 10) {real, imag} */,
  {32'h3f4a58fd, 32'h3f2897eb} /* (12, 5, 9) {real, imag} */,
  {32'h3ebe32db, 32'hbd3d766c} /* (12, 5, 8) {real, imag} */,
  {32'hbed6146b, 32'hbdd49664} /* (12, 5, 7) {real, imag} */,
  {32'h3e8ef28b, 32'h3e388fac} /* (12, 5, 6) {real, imag} */,
  {32'h3fa2f932, 32'h3f4a88df} /* (12, 5, 5) {real, imag} */,
  {32'hbdd18a98, 32'hbf8fa1ff} /* (12, 5, 4) {real, imag} */,
  {32'h3d169efc, 32'hbea47fc8} /* (12, 5, 3) {real, imag} */,
  {32'h3f16b9ec, 32'h3fbe9b2e} /* (12, 5, 2) {real, imag} */,
  {32'hc00f1aa0, 32'hc01778cd} /* (12, 5, 1) {real, imag} */,
  {32'hc0336c5a, 32'hbf51c64b} /* (12, 5, 0) {real, imag} */,
  {32'h3f727b0d, 32'h4006c60a} /* (12, 4, 31) {real, imag} */,
  {32'hc05cea31, 32'hc01ef263} /* (12, 4, 30) {real, imag} */,
  {32'h3e95a513, 32'hbe9e767e} /* (12, 4, 29) {real, imag} */,
  {32'h3f8d7230, 32'h3e587f00} /* (12, 4, 28) {real, imag} */,
  {32'hbf21bf81, 32'hbf89961c} /* (12, 4, 27) {real, imag} */,
  {32'hbd309fd0, 32'hbe61f966} /* (12, 4, 26) {real, imag} */,
  {32'h3f41bb7c, 32'h3d07b904} /* (12, 4, 25) {real, imag} */,
  {32'h3ea3a800, 32'hbee37b8e} /* (12, 4, 24) {real, imag} */,
  {32'hbe8eedca, 32'hbed6346c} /* (12, 4, 23) {real, imag} */,
  {32'hbdc6726b, 32'hbe6b4496} /* (12, 4, 22) {real, imag} */,
  {32'hbeb11b24, 32'h3f3e53de} /* (12, 4, 21) {real, imag} */,
  {32'h3eacc460, 32'hbe49beae} /* (12, 4, 20) {real, imag} */,
  {32'hbc7d0cf0, 32'hbe5cf40a} /* (12, 4, 19) {real, imag} */,
  {32'hbebff452, 32'h3dc7fd40} /* (12, 4, 18) {real, imag} */,
  {32'h3e02338f, 32'h3f035316} /* (12, 4, 17) {real, imag} */,
  {32'h3d37afbe, 32'hbd3b251e} /* (12, 4, 16) {real, imag} */,
  {32'hbdcc54b7, 32'h3ddd78bf} /* (12, 4, 15) {real, imag} */,
  {32'h3e5d89da, 32'hbe7ea952} /* (12, 4, 14) {real, imag} */,
  {32'hbe0fada2, 32'h3e9db3ae} /* (12, 4, 13) {real, imag} */,
  {32'hbee678b6, 32'hbd0de550} /* (12, 4, 12) {real, imag} */,
  {32'hbee2df5e, 32'hbe592f7f} /* (12, 4, 11) {real, imag} */,
  {32'hbd0847ca, 32'h3f329544} /* (12, 4, 10) {real, imag} */,
  {32'hbf068d64, 32'h3d1128a8} /* (12, 4, 9) {real, imag} */,
  {32'h3d25d519, 32'hbf9f6337} /* (12, 4, 8) {real, imag} */,
  {32'hbd700cdf, 32'hbd7d57e8} /* (12, 4, 7) {real, imag} */,
  {32'hbee4fdca, 32'h3ed3d029} /* (12, 4, 6) {real, imag} */,
  {32'h3f0753c1, 32'hbfc69815} /* (12, 4, 5) {real, imag} */,
  {32'h3d4ab608, 32'h3edd0d77} /* (12, 4, 4) {real, imag} */,
  {32'h3f263a80, 32'h3e8b4e3e} /* (12, 4, 3) {real, imag} */,
  {32'hc00a8819, 32'hc0257cce} /* (12, 4, 2) {real, imag} */,
  {32'h40b7d9a4, 32'h3f832bea} /* (12, 4, 1) {real, imag} */,
  {32'h3fa3de4b, 32'hbe2d0483} /* (12, 4, 0) {real, imag} */,
  {32'hc0af9341, 32'h4006f384} /* (12, 3, 31) {real, imag} */,
  {32'h400bdc71, 32'hc076a746} /* (12, 3, 30) {real, imag} */,
  {32'hbf42fd55, 32'h3ef1830f} /* (12, 3, 29) {real, imag} */,
  {32'h3fc5e4f9, 32'h3fa3d5ea} /* (12, 3, 28) {real, imag} */,
  {32'hbf26ba80, 32'h3e03b5f0} /* (12, 3, 27) {real, imag} */,
  {32'hbe2f6f4c, 32'h3efea88b} /* (12, 3, 26) {real, imag} */,
  {32'h3e679dbc, 32'h3daaa85f} /* (12, 3, 25) {real, imag} */,
  {32'h3f330560, 32'hbf4cfaf7} /* (12, 3, 24) {real, imag} */,
  {32'h3f40d3d6, 32'h3e09f5b6} /* (12, 3, 23) {real, imag} */,
  {32'h3d8f9476, 32'hbe7131d8} /* (12, 3, 22) {real, imag} */,
  {32'hbe8648f9, 32'h3d893eac} /* (12, 3, 21) {real, imag} */,
  {32'hbe1c74ba, 32'h3cfe70c4} /* (12, 3, 20) {real, imag} */,
  {32'hbe38b918, 32'hbe4ad76c} /* (12, 3, 19) {real, imag} */,
  {32'hbeb1414e, 32'hbecda552} /* (12, 3, 18) {real, imag} */,
  {32'hbc7d6064, 32'h3eb0ecf8} /* (12, 3, 17) {real, imag} */,
  {32'h3d2b2892, 32'h3e83207f} /* (12, 3, 16) {real, imag} */,
  {32'h3aa6f400, 32'hbda872c3} /* (12, 3, 15) {real, imag} */,
  {32'h3ec0d174, 32'hbf366366} /* (12, 3, 14) {real, imag} */,
  {32'h3e60bfcd, 32'h3cc11428} /* (12, 3, 13) {real, imag} */,
  {32'hbcf77728, 32'h3e802321} /* (12, 3, 12) {real, imag} */,
  {32'h3b9b77f8, 32'h3d70360a} /* (12, 3, 11) {real, imag} */,
  {32'h3edaeefa, 32'hbe573c36} /* (12, 3, 10) {real, imag} */,
  {32'hbe732a41, 32'h3d21388e} /* (12, 3, 9) {real, imag} */,
  {32'hbe9f6a52, 32'h3f11faf9} /* (12, 3, 8) {real, imag} */,
  {32'h3ec21172, 32'hbf040ec2} /* (12, 3, 7) {real, imag} */,
  {32'h3f60d454, 32'h3f274a15} /* (12, 3, 6) {real, imag} */,
  {32'h3cefd260, 32'h3f8c5d78} /* (12, 3, 5) {real, imag} */,
  {32'hbf27b10e, 32'h3dc836a2} /* (12, 3, 4) {real, imag} */,
  {32'hbf22e696, 32'hbdbb32f8} /* (12, 3, 3) {real, imag} */,
  {32'hbea8edd3, 32'hc04fd050} /* (12, 3, 2) {real, imag} */,
  {32'h4092a3e9, 32'h406a5577} /* (12, 3, 1) {real, imag} */,
  {32'hbe8d2149, 32'h3e47578c} /* (12, 3, 0) {real, imag} */,
  {32'hc217a83c, 32'hbef8cf0d} /* (12, 2, 31) {real, imag} */,
  {32'h4190d81c, 32'hc09eaae8} /* (12, 2, 30) {real, imag} */,
  {32'h3ec652fa, 32'h3f59fe6a} /* (12, 2, 29) {real, imag} */,
  {32'hbf5dc005, 32'h3fe4f300} /* (12, 2, 28) {real, imag} */,
  {32'h3f8a77f5, 32'hbffff0ed} /* (12, 2, 27) {real, imag} */,
  {32'h3f401a4f, 32'hbd838ca4} /* (12, 2, 26) {real, imag} */,
  {32'hbf2564aa, 32'h3d9e9024} /* (12, 2, 25) {real, imag} */,
  {32'h3e1fef56, 32'hbfad5feb} /* (12, 2, 24) {real, imag} */,
  {32'hbed5106e, 32'h3de2f3b2} /* (12, 2, 23) {real, imag} */,
  {32'hbca616c0, 32'h3e9de8c6} /* (12, 2, 22) {real, imag} */,
  {32'h3f182ee2, 32'hbe680d46} /* (12, 2, 21) {real, imag} */,
  {32'hbf0883d2, 32'h3da4e536} /* (12, 2, 20) {real, imag} */,
  {32'h3be4a3a0, 32'h3e407170} /* (12, 2, 19) {real, imag} */,
  {32'h3c87fa99, 32'hbf156b41} /* (12, 2, 18) {real, imag} */,
  {32'hbea23768, 32'h3e9c3d1c} /* (12, 2, 17) {real, imag} */,
  {32'h3dafd85c, 32'h3dde13b1} /* (12, 2, 16) {real, imag} */,
  {32'hbeb70633, 32'hbe1610f8} /* (12, 2, 15) {real, imag} */,
  {32'h3f1fb44e, 32'h3f352066} /* (12, 2, 14) {real, imag} */,
  {32'h3cd80674, 32'hbe076737} /* (12, 2, 13) {real, imag} */,
  {32'h3e49d1cf, 32'h3eff73f2} /* (12, 2, 12) {real, imag} */,
  {32'h3d835d5e, 32'h3f594946} /* (12, 2, 11) {real, imag} */,
  {32'hbe1c5747, 32'hbd83ad38} /* (12, 2, 10) {real, imag} */,
  {32'hbedda304, 32'hbd56421c} /* (12, 2, 9) {real, imag} */,
  {32'h3f123302, 32'h3eeedf45} /* (12, 2, 8) {real, imag} */,
  {32'hbf3aad82, 32'hbe2f3b90} /* (12, 2, 7) {real, imag} */,
  {32'h3e554688, 32'h3f6dd322} /* (12, 2, 6) {real, imag} */,
  {32'h3f9fe174, 32'h4014b361} /* (12, 2, 5) {real, imag} */,
  {32'hc03f031d, 32'hbfe13fe7} /* (12, 2, 4) {real, imag} */,
  {32'h3eead44f, 32'h3dcdec46} /* (12, 2, 3) {real, imag} */,
  {32'h4133884d, 32'hc08b266a} /* (12, 2, 2) {real, imag} */,
  {32'hc1a77074, 32'h401ec049} /* (12, 2, 1) {real, imag} */,
  {32'hc1970c5e, 32'hc02e9758} /* (12, 2, 0) {real, imag} */,
  {32'h42482ad4, 32'hc11e442a} /* (12, 1, 31) {real, imag} */,
  {32'hc14996dd, 32'h3f1d7d75} /* (12, 1, 30) {real, imag} */,
  {32'h3c4c7e60, 32'h3f514ad1} /* (12, 1, 29) {real, imag} */,
  {32'h4028dd31, 32'h3fc3f438} /* (12, 1, 28) {real, imag} */,
  {32'hc082d0df, 32'hbf12267f} /* (12, 1, 27) {real, imag} */,
  {32'h3eb7bf7e, 32'hbd43a2e8} /* (12, 1, 26) {real, imag} */,
  {32'h3c752830, 32'hbe43bb92} /* (12, 1, 25) {real, imag} */,
  {32'hbee3a5e7, 32'hbd453760} /* (12, 1, 24) {real, imag} */,
  {32'hbf070fa2, 32'hbe6ff2d8} /* (12, 1, 23) {real, imag} */,
  {32'h3f595c2a, 32'h3f51dde3} /* (12, 1, 22) {real, imag} */,
  {32'hbf3a5049, 32'h3f508e26} /* (12, 1, 21) {real, imag} */,
  {32'hbf34d5fa, 32'h3d948662} /* (12, 1, 20) {real, imag} */,
  {32'hbe3b366d, 32'h3ebb3332} /* (12, 1, 19) {real, imag} */,
  {32'h3f0bc016, 32'h3e1f11d7} /* (12, 1, 18) {real, imag} */,
  {32'h3ea4ae14, 32'h3e9f5256} /* (12, 1, 17) {real, imag} */,
  {32'h3c9d3b54, 32'h3d845edd} /* (12, 1, 16) {real, imag} */,
  {32'h3e8515ae, 32'h3e53341d} /* (12, 1, 15) {real, imag} */,
  {32'h3e4a4ffc, 32'hbdd1755e} /* (12, 1, 14) {real, imag} */,
  {32'hbda3e17f, 32'hbdb5f07d} /* (12, 1, 13) {real, imag} */,
  {32'h3e891fa2, 32'hbeedba92} /* (12, 1, 12) {real, imag} */,
  {32'hbd06ff92, 32'hbf2ca6b3} /* (12, 1, 11) {real, imag} */,
  {32'hbe90a74c, 32'hbde27cf8} /* (12, 1, 10) {real, imag} */,
  {32'hbe018bd4, 32'hbe355bcb} /* (12, 1, 9) {real, imag} */,
  {32'hbe98265b, 32'hbfad55c8} /* (12, 1, 8) {real, imag} */,
  {32'h3f1c62ee, 32'h3e7e0faa} /* (12, 1, 7) {real, imag} */,
  {32'hbd3dca10, 32'hbf786efc} /* (12, 1, 6) {real, imag} */,
  {32'hc017b820, 32'hbeb30fcc} /* (12, 1, 5) {real, imag} */,
  {32'hbf55e5f8, 32'h400a5466} /* (12, 1, 4) {real, imag} */,
  {32'hbefc7a62, 32'hbc31b2c0} /* (12, 1, 3) {real, imag} */,
  {32'hc1978599, 32'hc1840624} /* (12, 1, 2) {real, imag} */,
  {32'h428a1a57, 32'h42242047} /* (12, 1, 1) {real, imag} */,
  {32'h42827137, 32'h407c5dd8} /* (12, 1, 0) {real, imag} */,
  {32'h421cf0bc, 32'hc203701f} /* (12, 0, 31) {real, imag} */,
  {32'hc0c30253, 32'h411168d5} /* (12, 0, 30) {real, imag} */,
  {32'hbfbb3ad8, 32'h3ed4aeb0} /* (12, 0, 29) {real, imag} */,
  {32'h3d40c4de, 32'h3fb36765} /* (12, 0, 28) {real, imag} */,
  {32'hbfd42466, 32'h3e006153} /* (12, 0, 27) {real, imag} */,
  {32'hbf8cf3cc, 32'hbeb6a980} /* (12, 0, 26) {real, imag} */,
  {32'h3d42a6f6, 32'hbf796b02} /* (12, 0, 25) {real, imag} */,
  {32'hbe0e3e02, 32'h3f71e5c6} /* (12, 0, 24) {real, imag} */,
  {32'hbde688be, 32'h3f147590} /* (12, 0, 23) {real, imag} */,
  {32'hbf569249, 32'h3ed7f8e4} /* (12, 0, 22) {real, imag} */,
  {32'hbdd8c978, 32'hbe1d5898} /* (12, 0, 21) {real, imag} */,
  {32'hbe6f1c08, 32'hbd9b6488} /* (12, 0, 20) {real, imag} */,
  {32'hbc85d79c, 32'h3eb56a60} /* (12, 0, 19) {real, imag} */,
  {32'hbc629920, 32'hbee2bfce} /* (12, 0, 18) {real, imag} */,
  {32'hbd944bf5, 32'hbea1eb9c} /* (12, 0, 17) {real, imag} */,
  {32'h3dc175e4, 32'h00000000} /* (12, 0, 16) {real, imag} */,
  {32'hbd944bf5, 32'h3ea1eb9c} /* (12, 0, 15) {real, imag} */,
  {32'hbc629920, 32'h3ee2bfce} /* (12, 0, 14) {real, imag} */,
  {32'hbc85d79c, 32'hbeb56a60} /* (12, 0, 13) {real, imag} */,
  {32'hbe6f1c08, 32'h3d9b6488} /* (12, 0, 12) {real, imag} */,
  {32'hbdd8c978, 32'h3e1d5898} /* (12, 0, 11) {real, imag} */,
  {32'hbf569249, 32'hbed7f8e4} /* (12, 0, 10) {real, imag} */,
  {32'hbde688be, 32'hbf147590} /* (12, 0, 9) {real, imag} */,
  {32'hbe0e3e02, 32'hbf71e5c6} /* (12, 0, 8) {real, imag} */,
  {32'h3d42a6f6, 32'h3f796b02} /* (12, 0, 7) {real, imag} */,
  {32'hbf8cf3cc, 32'h3eb6a980} /* (12, 0, 6) {real, imag} */,
  {32'hbfd42466, 32'hbe006153} /* (12, 0, 5) {real, imag} */,
  {32'h3d40c4de, 32'hbfb36765} /* (12, 0, 4) {real, imag} */,
  {32'hbfbb3ad8, 32'hbed4aeb0} /* (12, 0, 3) {real, imag} */,
  {32'hc0c30253, 32'hc11168d5} /* (12, 0, 2) {real, imag} */,
  {32'h421cf0bc, 32'h4203701f} /* (12, 0, 1) {real, imag} */,
  {32'h427ee150, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h4299e3e7, 32'hc22fb621} /* (11, 31, 31) {real, imag} */,
  {32'hc1a3c4f9, 32'h4191f708} /* (11, 31, 30) {real, imag} */,
  {32'h3f1a8a95, 32'hbeaf0cb7} /* (11, 31, 29) {real, imag} */,
  {32'hbf090778, 32'hbf86aac5} /* (11, 31, 28) {real, imag} */,
  {32'hc04977e0, 32'h3f5b971f} /* (11, 31, 27) {real, imag} */,
  {32'hbf9ff0dc, 32'h3f1ed53d} /* (11, 31, 26) {real, imag} */,
  {32'h3ed375ce, 32'hbed247be} /* (11, 31, 25) {real, imag} */,
  {32'hbf2dc14c, 32'h3f5476fd} /* (11, 31, 24) {real, imag} */,
  {32'hbdea4a50, 32'hbec9b67f} /* (11, 31, 23) {real, imag} */,
  {32'hbd9b7a58, 32'h3f4c444a} /* (11, 31, 22) {real, imag} */,
  {32'hbe3e8105, 32'hbd8599f8} /* (11, 31, 21) {real, imag} */,
  {32'h3e810d18, 32'h3caadd90} /* (11, 31, 20) {real, imag} */,
  {32'h3e2ead9e, 32'h3e533833} /* (11, 31, 19) {real, imag} */,
  {32'h3de4843e, 32'h3ec94fd0} /* (11, 31, 18) {real, imag} */,
  {32'h3e02144c, 32'hbede22b7} /* (11, 31, 17) {real, imag} */,
  {32'h3e0d58e0, 32'hbd8b5178} /* (11, 31, 16) {real, imag} */,
  {32'h3de2abba, 32'h3db27d7b} /* (11, 31, 15) {real, imag} */,
  {32'h3ec92734, 32'hbe2cc043} /* (11, 31, 14) {real, imag} */,
  {32'hbed4bc87, 32'h3e811ae7} /* (11, 31, 13) {real, imag} */,
  {32'hbc74ff30, 32'h3e6bd418} /* (11, 31, 12) {real, imag} */,
  {32'hbf24b3b3, 32'hbf03fd85} /* (11, 31, 11) {real, imag} */,
  {32'h3f30ff67, 32'hbedd148e} /* (11, 31, 10) {real, imag} */,
  {32'hbe278aaa, 32'hbd16b98c} /* (11, 31, 9) {real, imag} */,
  {32'hbf3be2a0, 32'hbeb5c5c2} /* (11, 31, 8) {real, imag} */,
  {32'hbc9e8988, 32'h3cb8fcc0} /* (11, 31, 7) {real, imag} */,
  {32'hbebe4c19, 32'h3e979d96} /* (11, 31, 6) {real, imag} */,
  {32'hc04bfb52, 32'h3f42caa2} /* (11, 31, 5) {real, imag} */,
  {32'h4012dd6a, 32'hc019fd52} /* (11, 31, 4) {real, imag} */,
  {32'hbf860f91, 32'hbeb92c88} /* (11, 31, 3) {real, imag} */,
  {32'hc150f2a6, 32'hbfa397b6} /* (11, 31, 2) {real, imag} */,
  {32'h425828b8, 32'h4128e473} /* (11, 31, 1) {real, imag} */,
  {32'h428eea0c, 32'hc08f22b4} /* (11, 31, 0) {real, imag} */,
  {32'hc1b22ee0, 32'hc094410d} /* (11, 30, 31) {real, imag} */,
  {32'h414fd23c, 32'h4094bb92} /* (11, 30, 30) {real, imag} */,
  {32'h3f420d4e, 32'hbea83537} /* (11, 30, 29) {real, imag} */,
  {32'hc038eb7c, 32'h3fe0db92} /* (11, 30, 28) {real, imag} */,
  {32'h3f83386e, 32'hc027a44e} /* (11, 30, 27) {real, imag} */,
  {32'h3e7d25a2, 32'hbf006988} /* (11, 30, 26) {real, imag} */,
  {32'h3e7c800a, 32'h3eadf187} /* (11, 30, 25) {real, imag} */,
  {32'h3f39ea27, 32'h3e3bcba8} /* (11, 30, 24) {real, imag} */,
  {32'hbe1ec5e5, 32'hbdb048d6} /* (11, 30, 23) {real, imag} */,
  {32'hbee9774a, 32'hbedd6098} /* (11, 30, 22) {real, imag} */,
  {32'hbd9d7fdb, 32'hbeaa87b8} /* (11, 30, 21) {real, imag} */,
  {32'hbe261eab, 32'hbe9d2899} /* (11, 30, 20) {real, imag} */,
  {32'hbe0631ae, 32'hbeb72442} /* (11, 30, 19) {real, imag} */,
  {32'hbe73e864, 32'hbef43ab2} /* (11, 30, 18) {real, imag} */,
  {32'hbdd2eabc, 32'h3c8399b4} /* (11, 30, 17) {real, imag} */,
  {32'h3e8832fd, 32'hbe946250} /* (11, 30, 16) {real, imag} */,
  {32'hbdce5bdc, 32'h3c9afbc8} /* (11, 30, 15) {real, imag} */,
  {32'h3ddb82a4, 32'h3da4a3b0} /* (11, 30, 14) {real, imag} */,
  {32'h3e443f56, 32'h3e249ffc} /* (11, 30, 13) {real, imag} */,
  {32'h3dbc91c2, 32'h3e6d56de} /* (11, 30, 12) {real, imag} */,
  {32'h3e54685b, 32'h3f07d2e6} /* (11, 30, 11) {real, imag} */,
  {32'hbe3819b6, 32'hbd57072e} /* (11, 30, 10) {real, imag} */,
  {32'hbec4d794, 32'hbd5c5d61} /* (11, 30, 9) {real, imag} */,
  {32'h3f1d2549, 32'h3f28191e} /* (11, 30, 8) {real, imag} */,
  {32'h3d87a0e0, 32'hbf19f4ae} /* (11, 30, 7) {real, imag} */,
  {32'h3f2733b4, 32'hbd2e574c} /* (11, 30, 6) {real, imag} */,
  {32'h3fe5d2a9, 32'h3ff8bc99} /* (11, 30, 5) {real, imag} */,
  {32'hbf1dab10, 32'hc015816a} /* (11, 30, 4) {real, imag} */,
  {32'h3ee63a8e, 32'hbf0f9b23} /* (11, 30, 3) {real, imag} */,
  {32'h41946cf5, 32'h40a9b6b9} /* (11, 30, 2) {real, imag} */,
  {32'hc222d3e7, 32'h4025fec6} /* (11, 30, 1) {real, imag} */,
  {32'hc1b05fe6, 32'h403997dd} /* (11, 30, 0) {real, imag} */,
  {32'h407a8474, 32'hc0384752} /* (11, 29, 31) {real, imag} */,
  {32'h3e6a39a6, 32'h403f8072} /* (11, 29, 30) {real, imag} */,
  {32'hbf6791f8, 32'hbf1ded94} /* (11, 29, 29) {real, imag} */,
  {32'hbf70392a, 32'hbeaa3156} /* (11, 29, 28) {real, imag} */,
  {32'hbe5c2517, 32'hbf045129} /* (11, 29, 27) {real, imag} */,
  {32'h3eabb0d2, 32'hbef33f0e} /* (11, 29, 26) {real, imag} */,
  {32'h3dcea700, 32'h3eeaf6a7} /* (11, 29, 25) {real, imag} */,
  {32'h3c1138e0, 32'h3e70f7d0} /* (11, 29, 24) {real, imag} */,
  {32'hbdf16e68, 32'hbdc1a13a} /* (11, 29, 23) {real, imag} */,
  {32'h3d1710a0, 32'hbe6d1b36} /* (11, 29, 22) {real, imag} */,
  {32'h3e88b0bc, 32'hbb0c3880} /* (11, 29, 21) {real, imag} */,
  {32'hbe812b32, 32'hbde951ac} /* (11, 29, 20) {real, imag} */,
  {32'h3e6cedaa, 32'h3e086d88} /* (11, 29, 19) {real, imag} */,
  {32'h3ee76c87, 32'h3f251786} /* (11, 29, 18) {real, imag} */,
  {32'hbebb24df, 32'hbe8e0241} /* (11, 29, 17) {real, imag} */,
  {32'h3e3d5da3, 32'hbde1fd4c} /* (11, 29, 16) {real, imag} */,
  {32'h3e3d38b9, 32'hbf041238} /* (11, 29, 15) {real, imag} */,
  {32'h3eb4affd, 32'h3da0026a} /* (11, 29, 14) {real, imag} */,
  {32'hbf07b2e5, 32'h3e014518} /* (11, 29, 13) {real, imag} */,
  {32'h3de4c866, 32'hbdd47bf8} /* (11, 29, 12) {real, imag} */,
  {32'h3ea2f6f6, 32'hbed8ef20} /* (11, 29, 11) {real, imag} */,
  {32'hbe24b3df, 32'hbd3cf700} /* (11, 29, 10) {real, imag} */,
  {32'h3cf1a5d8, 32'h3f14ef0d} /* (11, 29, 9) {real, imag} */,
  {32'h3efb6f24, 32'h3e854884} /* (11, 29, 8) {real, imag} */,
  {32'h3ed6db18, 32'hbed4215b} /* (11, 29, 7) {real, imag} */,
  {32'h3ef68f00, 32'hbf3e8ddb} /* (11, 29, 6) {real, imag} */,
  {32'hbf9c72a8, 32'hbf2b8ddc} /* (11, 29, 5) {real, imag} */,
  {32'h3f9165ae, 32'hbfa3b7ce} /* (11, 29, 4) {real, imag} */,
  {32'hbf04aeb0, 32'hbdf15d71} /* (11, 29, 3) {real, imag} */,
  {32'h3ff5944e, 32'h4091ba98} /* (11, 29, 2) {real, imag} */,
  {32'hc08b19d8, 32'hc0269cd3} /* (11, 29, 1) {real, imag} */,
  {32'h3e5248fc, 32'hbecf0fc0} /* (11, 29, 0) {real, imag} */,
  {32'h40c08df8, 32'hbf9aa2ac} /* (11, 28, 31) {real, imag} */,
  {32'hc025b734, 32'h3feaf7c2} /* (11, 28, 30) {real, imag} */,
  {32'h3f44c972, 32'hbd0db810} /* (11, 28, 29) {real, imag} */,
  {32'h3e0864dc, 32'hbf9d08d7} /* (11, 28, 28) {real, imag} */,
  {32'h3f144aaa, 32'h3f3d6c61} /* (11, 28, 27) {real, imag} */,
  {32'hbee1ea33, 32'hbf4cde3e} /* (11, 28, 26) {real, imag} */,
  {32'h3edd8def, 32'h3ec6b910} /* (11, 28, 25) {real, imag} */,
  {32'hbf0470a1, 32'h3f1d0aa0} /* (11, 28, 24) {real, imag} */,
  {32'hbe6fe966, 32'hbea02c9a} /* (11, 28, 23) {real, imag} */,
  {32'hbf2c3ae6, 32'h3e1685fd} /* (11, 28, 22) {real, imag} */,
  {32'h3da61298, 32'h3e0a158f} /* (11, 28, 21) {real, imag} */,
  {32'h3e174fb1, 32'hbd36711f} /* (11, 28, 20) {real, imag} */,
  {32'hbdbd8d3c, 32'hbd05ca08} /* (11, 28, 19) {real, imag} */,
  {32'h3eb47fd0, 32'h3ed4a1c6} /* (11, 28, 18) {real, imag} */,
  {32'hbd54d751, 32'h3d8c8a8c} /* (11, 28, 17) {real, imag} */,
  {32'h3cde33e4, 32'hbe09c9a2} /* (11, 28, 16) {real, imag} */,
  {32'h3e220678, 32'hbe1290b5} /* (11, 28, 15) {real, imag} */,
  {32'hbe522f46, 32'h3f219aa7} /* (11, 28, 14) {real, imag} */,
  {32'h3e3f2560, 32'hbe3cba06} /* (11, 28, 13) {real, imag} */,
  {32'h3f1d46bd, 32'hbe8f87bd} /* (11, 28, 12) {real, imag} */,
  {32'hbee0655e, 32'hbe19afab} /* (11, 28, 11) {real, imag} */,
  {32'hbe7226ea, 32'h3e00b536} /* (11, 28, 10) {real, imag} */,
  {32'h3f147f2e, 32'h3e9ab064} /* (11, 28, 9) {real, imag} */,
  {32'hbd12162c, 32'h3e87a07a} /* (11, 28, 8) {real, imag} */,
  {32'h3f192fcc, 32'hbe8f1535} /* (11, 28, 7) {real, imag} */,
  {32'hbe5f84ac, 32'h3e192348} /* (11, 28, 6) {real, imag} */,
  {32'hbe172a33, 32'hbe867687} /* (11, 28, 5) {real, imag} */,
  {32'h3e2cb6dd, 32'h3d4c8da0} /* (11, 28, 4) {real, imag} */,
  {32'hbeaa0525, 32'h3ed6b3d5} /* (11, 28, 3) {real, imag} */,
  {32'hc06acd1f, 32'h402eaad3} /* (11, 28, 2) {real, imag} */,
  {32'h3f712752, 32'hc03171a3} /* (11, 28, 1) {real, imag} */,
  {32'h3fb71a2a, 32'h3c53c900} /* (11, 28, 0) {real, imag} */,
  {32'hbed2afba, 32'h401b86e8} /* (11, 27, 31) {real, imag} */,
  {32'h3f1c603c, 32'hbf62af0e} /* (11, 27, 30) {real, imag} */,
  {32'hbf61aeae, 32'h3e9ab5d8} /* (11, 27, 29) {real, imag} */,
  {32'h3e3385ed, 32'h3e8fdb2b} /* (11, 27, 28) {real, imag} */,
  {32'h3f8c3aec, 32'h3ae5d000} /* (11, 27, 27) {real, imag} */,
  {32'hbf86c45e, 32'h3ce43060} /* (11, 27, 26) {real, imag} */,
  {32'h3e457cf0, 32'hbea66bd1} /* (11, 27, 25) {real, imag} */,
  {32'h3f158817, 32'hbf3456b8} /* (11, 27, 24) {real, imag} */,
  {32'hbe5808dd, 32'h3e759015} /* (11, 27, 23) {real, imag} */,
  {32'hbeec06de, 32'hbebd5356} /* (11, 27, 22) {real, imag} */,
  {32'h3f27ecc2, 32'h3e97f42c} /* (11, 27, 21) {real, imag} */,
  {32'h3e999806, 32'hbf21c47b} /* (11, 27, 20) {real, imag} */,
  {32'h3e993244, 32'hbe55e48a} /* (11, 27, 19) {real, imag} */,
  {32'hbe568376, 32'hbe5dd840} /* (11, 27, 18) {real, imag} */,
  {32'h3e9ad574, 32'h3e469c88} /* (11, 27, 17) {real, imag} */,
  {32'hbe66084e, 32'hbdd32214} /* (11, 27, 16) {real, imag} */,
  {32'h3c5b8f30, 32'hbd8f20ed} /* (11, 27, 15) {real, imag} */,
  {32'hbe6c6be4, 32'hbe2e0a89} /* (11, 27, 14) {real, imag} */,
  {32'h3f13b0f3, 32'hbed2a230} /* (11, 27, 13) {real, imag} */,
  {32'h3e5d3ebd, 32'hbb9af880} /* (11, 27, 12) {real, imag} */,
  {32'hbe3b3320, 32'h3f0b8876} /* (11, 27, 11) {real, imag} */,
  {32'h3df2929e, 32'hbe3d5cf2} /* (11, 27, 10) {real, imag} */,
  {32'hbda6fa62, 32'h3e8064bc} /* (11, 27, 9) {real, imag} */,
  {32'h3eed21c6, 32'h3f954064} /* (11, 27, 8) {real, imag} */,
  {32'h3e287fe2, 32'h3dcd7b0d} /* (11, 27, 7) {real, imag} */,
  {32'h3ec4eb58, 32'h3e99232a} /* (11, 27, 6) {real, imag} */,
  {32'h3eb895f0, 32'hbf1b62d4} /* (11, 27, 5) {real, imag} */,
  {32'hbeff6a43, 32'hbfcc7d5a} /* (11, 27, 4) {real, imag} */,
  {32'hbf2c5d22, 32'hbe405c8f} /* (11, 27, 3) {real, imag} */,
  {32'h3eb10ea8, 32'h3c455ca0} /* (11, 27, 2) {real, imag} */,
  {32'hc05d9576, 32'h3e022142} /* (11, 27, 1) {real, imag} */,
  {32'hbfe523e2, 32'h3f33bf32} /* (11, 27, 0) {real, imag} */,
  {32'h3e496e12, 32'hbdfa914c} /* (11, 26, 31) {real, imag} */,
  {32'h3f3d3b27, 32'hbdaec9d4} /* (11, 26, 30) {real, imag} */,
  {32'h3eacf6ce, 32'hbebb53ce} /* (11, 26, 29) {real, imag} */,
  {32'h3dd7e907, 32'hbd0121ee} /* (11, 26, 28) {real, imag} */,
  {32'h3dde31f8, 32'h3e7f9437} /* (11, 26, 27) {real, imag} */,
  {32'h3ee78efc, 32'h3e916e6f} /* (11, 26, 26) {real, imag} */,
  {32'h3e30c996, 32'hbe438d3f} /* (11, 26, 25) {real, imag} */,
  {32'hbeb1b418, 32'h3f206d98} /* (11, 26, 24) {real, imag} */,
  {32'hbea1182b, 32'h3d8bfc3c} /* (11, 26, 23) {real, imag} */,
  {32'hbdbfbdf4, 32'hbe4e27d4} /* (11, 26, 22) {real, imag} */,
  {32'h3d128438, 32'h3f177d73} /* (11, 26, 21) {real, imag} */,
  {32'hbd44be28, 32'h3ebd48fb} /* (11, 26, 20) {real, imag} */,
  {32'h3cd834ba, 32'hbe739882} /* (11, 26, 19) {real, imag} */,
  {32'hbe3887f2, 32'hbe208380} /* (11, 26, 18) {real, imag} */,
  {32'hbd2420db, 32'hbd045aae} /* (11, 26, 17) {real, imag} */,
  {32'h3e1365f0, 32'hbd960636} /* (11, 26, 16) {real, imag} */,
  {32'h3e8eadfe, 32'h3ed3b2f1} /* (11, 26, 15) {real, imag} */,
  {32'hbe28c3f6, 32'hbe9c6a6e} /* (11, 26, 14) {real, imag} */,
  {32'hbe34c180, 32'hbef721e5} /* (11, 26, 13) {real, imag} */,
  {32'h3d1137b0, 32'h3e7d4931} /* (11, 26, 12) {real, imag} */,
  {32'h3e1dd059, 32'hbea02712} /* (11, 26, 11) {real, imag} */,
  {32'h3ef72a30, 32'hbea22b18} /* (11, 26, 10) {real, imag} */,
  {32'h3e64c837, 32'hbf27a0c4} /* (11, 26, 9) {real, imag} */,
  {32'hbdaf5070, 32'hbf1b8af7} /* (11, 26, 8) {real, imag} */,
  {32'hbe3778a6, 32'h3ea446f7} /* (11, 26, 7) {real, imag} */,
  {32'h3e9ccf90, 32'hbf4d0c5c} /* (11, 26, 6) {real, imag} */,
  {32'h3f271be8, 32'hbca172e0} /* (11, 26, 5) {real, imag} */,
  {32'h3ef13f90, 32'h3f83cec3} /* (11, 26, 4) {real, imag} */,
  {32'h3e11186f, 32'h3ed2a84f} /* (11, 26, 3) {real, imag} */,
  {32'h3caec7f0, 32'h3f1a41e2} /* (11, 26, 2) {real, imag} */,
  {32'h3f7382c9, 32'h3fa32261} /* (11, 26, 1) {real, imag} */,
  {32'h3df8911e, 32'hbf19aa50} /* (11, 26, 0) {real, imag} */,
  {32'hbde0d314, 32'hbe96a4fc} /* (11, 25, 31) {real, imag} */,
  {32'hbdea312c, 32'hbdf8a121} /* (11, 25, 30) {real, imag} */,
  {32'h3d8b8ac8, 32'h3dee98b8} /* (11, 25, 29) {real, imag} */,
  {32'h3f2e6631, 32'hbe33dd2e} /* (11, 25, 28) {real, imag} */,
  {32'hbf4b1748, 32'h3de69f6a} /* (11, 25, 27) {real, imag} */,
  {32'h3e91be26, 32'h3f833c4d} /* (11, 25, 26) {real, imag} */,
  {32'h3e646a5a, 32'hbf09aafa} /* (11, 25, 25) {real, imag} */,
  {32'h3ef76976, 32'h3e005d6e} /* (11, 25, 24) {real, imag} */,
  {32'hbdd3c95a, 32'h3d256820} /* (11, 25, 23) {real, imag} */,
  {32'h3ed14df9, 32'hbe529eee} /* (11, 25, 22) {real, imag} */,
  {32'h3e9414b0, 32'h3df14dfa} /* (11, 25, 21) {real, imag} */,
  {32'hbe422bf9, 32'h3dfc8c97} /* (11, 25, 20) {real, imag} */,
  {32'hbe3237b0, 32'hbe9fc0a6} /* (11, 25, 19) {real, imag} */,
  {32'hbe057f89, 32'h3d506940} /* (11, 25, 18) {real, imag} */,
  {32'hbde92234, 32'hbdc99aee} /* (11, 25, 17) {real, imag} */,
  {32'hbe8c16fe, 32'hbec322db} /* (11, 25, 16) {real, imag} */,
  {32'hbe19e815, 32'h3e9055f4} /* (11, 25, 15) {real, imag} */,
  {32'hbea36167, 32'hbcbecba8} /* (11, 25, 14) {real, imag} */,
  {32'h3f1a8ff8, 32'hbf83f69d} /* (11, 25, 13) {real, imag} */,
  {32'h3e0ee328, 32'hbd2431d7} /* (11, 25, 12) {real, imag} */,
  {32'h3e9e146e, 32'hbef2cda1} /* (11, 25, 11) {real, imag} */,
  {32'hbe168f50, 32'hbec70a82} /* (11, 25, 10) {real, imag} */,
  {32'hbedf1173, 32'hbea355d0} /* (11, 25, 9) {real, imag} */,
  {32'hbf7d756e, 32'h3eca1301} /* (11, 25, 8) {real, imag} */,
  {32'h3f1e7bb1, 32'h3bdfcf80} /* (11, 25, 7) {real, imag} */,
  {32'hbea12222, 32'h3df766e0} /* (11, 25, 6) {real, imag} */,
  {32'h3ea651bb, 32'hbea1b3fe} /* (11, 25, 5) {real, imag} */,
  {32'hbe2f5151, 32'hbe5eb02a} /* (11, 25, 4) {real, imag} */,
  {32'h3eec3f48, 32'hbead2d1a} /* (11, 25, 3) {real, imag} */,
  {32'hbe8cbe28, 32'hbd1c4440} /* (11, 25, 2) {real, imag} */,
  {32'h3f2d2a66, 32'hbe9a4ffc} /* (11, 25, 1) {real, imag} */,
  {32'h3e9efa4e, 32'hbe815e98} /* (11, 25, 0) {real, imag} */,
  {32'hbf84a9f2, 32'h3eb331fa} /* (11, 24, 31) {real, imag} */,
  {32'h3f953914, 32'hbf2dfb5d} /* (11, 24, 30) {real, imag} */,
  {32'hbdf0239e, 32'h3e7c8c1d} /* (11, 24, 29) {real, imag} */,
  {32'hbf80dcdc, 32'h3e6926af} /* (11, 24, 28) {real, imag} */,
  {32'h3d741750, 32'hbea874d9} /* (11, 24, 27) {real, imag} */,
  {32'h3e6f565e, 32'hbedbfcbf} /* (11, 24, 26) {real, imag} */,
  {32'hbf215946, 32'h3e9bf3ab} /* (11, 24, 25) {real, imag} */,
  {32'hbeddd500, 32'h3dadc656} /* (11, 24, 24) {real, imag} */,
  {32'hbed5ce7a, 32'h3f011965} /* (11, 24, 23) {real, imag} */,
  {32'h3e63c7f9, 32'hbee47665} /* (11, 24, 22) {real, imag} */,
  {32'hbe44d19c, 32'hbf02e78f} /* (11, 24, 21) {real, imag} */,
  {32'h3eb833d1, 32'h3efa3d9e} /* (11, 24, 20) {real, imag} */,
  {32'hbe4dceea, 32'h3e378920} /* (11, 24, 19) {real, imag} */,
  {32'h3ed3b056, 32'hbeb773e8} /* (11, 24, 18) {real, imag} */,
  {32'hbf0f04f8, 32'hbd94091a} /* (11, 24, 17) {real, imag} */,
  {32'hbc5ec990, 32'hbdae279a} /* (11, 24, 16) {real, imag} */,
  {32'hbdc52532, 32'hbe395ec6} /* (11, 24, 15) {real, imag} */,
  {32'h3e98ede9, 32'hbd0b25cc} /* (11, 24, 14) {real, imag} */,
  {32'hbd02f46f, 32'h3d512ee8} /* (11, 24, 13) {real, imag} */,
  {32'h3f05e238, 32'hbe09b4d3} /* (11, 24, 12) {real, imag} */,
  {32'h3e3e4f85, 32'h3e36f008} /* (11, 24, 11) {real, imag} */,
  {32'h3f212279, 32'hbda445e2} /* (11, 24, 10) {real, imag} */,
  {32'h3e01bd6e, 32'hbc886570} /* (11, 24, 9) {real, imag} */,
  {32'hbefe0448, 32'h3eae5000} /* (11, 24, 8) {real, imag} */,
  {32'h3e912d4e, 32'h3f3ef202} /* (11, 24, 7) {real, imag} */,
  {32'h3d0d93e8, 32'hbfa38c64} /* (11, 24, 6) {real, imag} */,
  {32'h3cdaabb0, 32'h3e9da75e} /* (11, 24, 5) {real, imag} */,
  {32'h3ec76264, 32'hbe9808f9} /* (11, 24, 4) {real, imag} */,
  {32'hbf89217c, 32'hbdeabc1e} /* (11, 24, 3) {real, imag} */,
  {32'h3f898232, 32'h3e677cc2} /* (11, 24, 2) {real, imag} */,
  {32'hbfda8b79, 32'h3f751222} /* (11, 24, 1) {real, imag} */,
  {32'h3d510ab4, 32'h3f1e97e1} /* (11, 24, 0) {real, imag} */,
  {32'h3e70aee9, 32'hbf1c7f16} /* (11, 23, 31) {real, imag} */,
  {32'hbdac88ba, 32'h3f4a0b98} /* (11, 23, 30) {real, imag} */,
  {32'h3eb69645, 32'h3eca50e5} /* (11, 23, 29) {real, imag} */,
  {32'hbf1b5f7a, 32'hbcc6ec5c} /* (11, 23, 28) {real, imag} */,
  {32'h3dc0ac38, 32'hbd402a8c} /* (11, 23, 27) {real, imag} */,
  {32'h3dbc9064, 32'hbdad84bc} /* (11, 23, 26) {real, imag} */,
  {32'hbdddc92d, 32'h3f1799ac} /* (11, 23, 25) {real, imag} */,
  {32'hbebe460c, 32'h3f0ec476} /* (11, 23, 24) {real, imag} */,
  {32'h3d90ead4, 32'hbf3fa93a} /* (11, 23, 23) {real, imag} */,
  {32'hbea8e8e6, 32'hbf09faa8} /* (11, 23, 22) {real, imag} */,
  {32'hbe81576e, 32'hbc5522d0} /* (11, 23, 21) {real, imag} */,
  {32'h3eb4be96, 32'h3f2f811e} /* (11, 23, 20) {real, imag} */,
  {32'hbf3ff504, 32'h3e95b854} /* (11, 23, 19) {real, imag} */,
  {32'h3c08e448, 32'hbd0f42a4} /* (11, 23, 18) {real, imag} */,
  {32'hbdcf503f, 32'hbad2cfc0} /* (11, 23, 17) {real, imag} */,
  {32'hbe09bd6c, 32'h3dead762} /* (11, 23, 16) {real, imag} */,
  {32'hbdc2613f, 32'hbe256aea} /* (11, 23, 15) {real, imag} */,
  {32'hbb897f40, 32'hbe8dbfaa} /* (11, 23, 14) {real, imag} */,
  {32'h3f86eaa8, 32'h3e865e67} /* (11, 23, 13) {real, imag} */,
  {32'h3e0282d8, 32'hbecbb1ab} /* (11, 23, 12) {real, imag} */,
  {32'hbeaad22d, 32'h3ec18e8c} /* (11, 23, 11) {real, imag} */,
  {32'hbe207753, 32'h3f44f3b6} /* (11, 23, 10) {real, imag} */,
  {32'hbe07df60, 32'hbea8f6ba} /* (11, 23, 9) {real, imag} */,
  {32'h3e607521, 32'hbef464f5} /* (11, 23, 8) {real, imag} */,
  {32'h3bde8d80, 32'hbeb241a2} /* (11, 23, 7) {real, imag} */,
  {32'h3ef86a6f, 32'h3edde02e} /* (11, 23, 6) {real, imag} */,
  {32'hbe8c7099, 32'hbd8061ee} /* (11, 23, 5) {real, imag} */,
  {32'hbe095366, 32'h3df8bf2c} /* (11, 23, 4) {real, imag} */,
  {32'h3e901d72, 32'hbd1d8090} /* (11, 23, 3) {real, imag} */,
  {32'h3ecd0668, 32'h3f1ccfe2} /* (11, 23, 2) {real, imag} */,
  {32'hbf984f52, 32'hbf04d277} /* (11, 23, 1) {real, imag} */,
  {32'h3d3538c0, 32'h3d70d664} /* (11, 23, 0) {real, imag} */,
  {32'hbe20c462, 32'hbf537303} /* (11, 22, 31) {real, imag} */,
  {32'h3e98ce9f, 32'h3edf67af} /* (11, 22, 30) {real, imag} */,
  {32'h3d22fa94, 32'hbefe02ba} /* (11, 22, 29) {real, imag} */,
  {32'h3ebdd00e, 32'hbf5dffd4} /* (11, 22, 28) {real, imag} */,
  {32'h3f53c16c, 32'h3e9bd967} /* (11, 22, 27) {real, imag} */,
  {32'h3e7a3b61, 32'h3f2e1520} /* (11, 22, 26) {real, imag} */,
  {32'hbe7268c6, 32'h3d98f59f} /* (11, 22, 25) {real, imag} */,
  {32'hbd082b3e, 32'h3e48ed3e} /* (11, 22, 24) {real, imag} */,
  {32'h3eeaf9ec, 32'hbe831f08} /* (11, 22, 23) {real, imag} */,
  {32'hbd06bd9c, 32'h3f1387fd} /* (11, 22, 22) {real, imag} */,
  {32'h3ca2d1e0, 32'h3c6a53ec} /* (11, 22, 21) {real, imag} */,
  {32'hbd0e4ae4, 32'h3d89aee4} /* (11, 22, 20) {real, imag} */,
  {32'h3db092fd, 32'hbe9dc1d2} /* (11, 22, 19) {real, imag} */,
  {32'h3e2bbcd6, 32'h39b03700} /* (11, 22, 18) {real, imag} */,
  {32'hbe53228e, 32'hbe5a562f} /* (11, 22, 17) {real, imag} */,
  {32'hbeb19682, 32'h3db6da8c} /* (11, 22, 16) {real, imag} */,
  {32'h3f0e6d35, 32'hbf0a5b19} /* (11, 22, 15) {real, imag} */,
  {32'h3b867e88, 32'h3f048862} /* (11, 22, 14) {real, imag} */,
  {32'hbdf9ffba, 32'h3e4a1133} /* (11, 22, 13) {real, imag} */,
  {32'hbda925b3, 32'hbe8c407c} /* (11, 22, 12) {real, imag} */,
  {32'h3e1afe57, 32'hbdb590ef} /* (11, 22, 11) {real, imag} */,
  {32'hbdd52da9, 32'hbe1b4a54} /* (11, 22, 10) {real, imag} */,
  {32'h3dfcda40, 32'hbeda0be4} /* (11, 22, 9) {real, imag} */,
  {32'hbe15afdb, 32'h3d9b9178} /* (11, 22, 8) {real, imag} */,
  {32'hbe6fc91f, 32'hbdf0e1aa} /* (11, 22, 7) {real, imag} */,
  {32'h3da05897, 32'h3e5150f6} /* (11, 22, 6) {real, imag} */,
  {32'hbf5c28b8, 32'h3d652cf4} /* (11, 22, 5) {real, imag} */,
  {32'h3f1455c2, 32'h3eaf83a5} /* (11, 22, 4) {real, imag} */,
  {32'hbdd5a50f, 32'h3eaa051c} /* (11, 22, 3) {real, imag} */,
  {32'hbe1f7792, 32'hbc1538c0} /* (11, 22, 2) {real, imag} */,
  {32'h3ceb9808, 32'hbf521d4a} /* (11, 22, 1) {real, imag} */,
  {32'h3e865a20, 32'h3f1f1d5c} /* (11, 22, 0) {real, imag} */,
  {32'hbd92ec86, 32'h3f1039a0} /* (11, 21, 31) {real, imag} */,
  {32'hbeb8ee30, 32'hbf9b35fa} /* (11, 21, 30) {real, imag} */,
  {32'hbe6b313e, 32'hbf3307cc} /* (11, 21, 29) {real, imag} */,
  {32'h3f23fbab, 32'h3ebd531d} /* (11, 21, 28) {real, imag} */,
  {32'h3e14d8cc, 32'hbf145781} /* (11, 21, 27) {real, imag} */,
  {32'h3e925f86, 32'h3e697029} /* (11, 21, 26) {real, imag} */,
  {32'hbee5c47d, 32'hbf289a4a} /* (11, 21, 25) {real, imag} */,
  {32'h3ea075c7, 32'hbdd4866c} /* (11, 21, 24) {real, imag} */,
  {32'h3f50c1f3, 32'h3ea84b4a} /* (11, 21, 23) {real, imag} */,
  {32'h3d5228dc, 32'h3e2c909c} /* (11, 21, 22) {real, imag} */,
  {32'hbe9e15db, 32'h3d8b6dbb} /* (11, 21, 21) {real, imag} */,
  {32'h3d9523e6, 32'h3dd734d8} /* (11, 21, 20) {real, imag} */,
  {32'hbe5389a6, 32'hbe9e0c86} /* (11, 21, 19) {real, imag} */,
  {32'h3dab0bda, 32'h3e280de6} /* (11, 21, 18) {real, imag} */,
  {32'hbda50bf2, 32'h3e5c7f05} /* (11, 21, 17) {real, imag} */,
  {32'h3de6e886, 32'hbeabbf1b} /* (11, 21, 16) {real, imag} */,
  {32'h3dcb7bc2, 32'h3c8a608c} /* (11, 21, 15) {real, imag} */,
  {32'hbe1deea0, 32'hbee7038a} /* (11, 21, 14) {real, imag} */,
  {32'hbebf1045, 32'hbeb77c16} /* (11, 21, 13) {real, imag} */,
  {32'h3eba9203, 32'hbdfffb18} /* (11, 21, 12) {real, imag} */,
  {32'h3ebffb10, 32'hbdcce78f} /* (11, 21, 11) {real, imag} */,
  {32'hbcde28d8, 32'h3e9b4528} /* (11, 21, 10) {real, imag} */,
  {32'hbef5e3d4, 32'h3ed82d8b} /* (11, 21, 9) {real, imag} */,
  {32'h3eb3a3a4, 32'h3e712c23} /* (11, 21, 8) {real, imag} */,
  {32'h3e032bbc, 32'hbf0be722} /* (11, 21, 7) {real, imag} */,
  {32'hbedc2d73, 32'h3e98c248} /* (11, 21, 6) {real, imag} */,
  {32'hbd466ff4, 32'hbe3e0c47} /* (11, 21, 5) {real, imag} */,
  {32'hbe9de1f4, 32'hbecfe524} /* (11, 21, 4) {real, imag} */,
  {32'h3e07ed19, 32'h3e4f819d} /* (11, 21, 3) {real, imag} */,
  {32'h3f79d3a5, 32'h3d14ec22} /* (11, 21, 2) {real, imag} */,
  {32'hbdb380c4, 32'h3efb3e32} /* (11, 21, 1) {real, imag} */,
  {32'hbeb5545f, 32'h3f216ea7} /* (11, 21, 0) {real, imag} */,
  {32'hbde3695b, 32'h3e15891c} /* (11, 20, 31) {real, imag} */,
  {32'h3ef2e050, 32'hbf0d7f35} /* (11, 20, 30) {real, imag} */,
  {32'h3e22d303, 32'hbe13375d} /* (11, 20, 29) {real, imag} */,
  {32'h3e738eff, 32'h3ea772a9} /* (11, 20, 28) {real, imag} */,
  {32'hbe0ffabb, 32'h3ee285c3} /* (11, 20, 27) {real, imag} */,
  {32'h3e41ffaf, 32'h3e9ab223} /* (11, 20, 26) {real, imag} */,
  {32'hbd6b6770, 32'h3f4c102a} /* (11, 20, 25) {real, imag} */,
  {32'h3e6f5be3, 32'hbe9d7268} /* (11, 20, 24) {real, imag} */,
  {32'hbf2121f3, 32'h3eca41b9} /* (11, 20, 23) {real, imag} */,
  {32'h3e452cd5, 32'h3e55974e} /* (11, 20, 22) {real, imag} */,
  {32'h3c503760, 32'hbe89f1bb} /* (11, 20, 21) {real, imag} */,
  {32'h3db20812, 32'hbeb841ec} /* (11, 20, 20) {real, imag} */,
  {32'hbe766565, 32'hbd537c0e} /* (11, 20, 19) {real, imag} */,
  {32'hbe878bea, 32'hbd03e6e8} /* (11, 20, 18) {real, imag} */,
  {32'h3d9e775d, 32'hbd23f000} /* (11, 20, 17) {real, imag} */,
  {32'hbccc20e0, 32'h3ed24812} /* (11, 20, 16) {real, imag} */,
  {32'hbe07b7b6, 32'h3b81d900} /* (11, 20, 15) {real, imag} */,
  {32'hbeb72d10, 32'h3e565268} /* (11, 20, 14) {real, imag} */,
  {32'h3ceafb29, 32'hbd9bc556} /* (11, 20, 13) {real, imag} */,
  {32'hbdeaa10f, 32'hbebfd042} /* (11, 20, 12) {real, imag} */,
  {32'hbf44d284, 32'hbda4c847} /* (11, 20, 11) {real, imag} */,
  {32'h3eac6647, 32'h3bd53848} /* (11, 20, 10) {real, imag} */,
  {32'hbe86c1d8, 32'hbec0a258} /* (11, 20, 9) {real, imag} */,
  {32'h3e958ee5, 32'h3c328be0} /* (11, 20, 8) {real, imag} */,
  {32'h3e65d586, 32'hbe3ae68b} /* (11, 20, 7) {real, imag} */,
  {32'h3e257376, 32'hbf0fdb31} /* (11, 20, 6) {real, imag} */,
  {32'hbc353f78, 32'h3ee2c80d} /* (11, 20, 5) {real, imag} */,
  {32'hbe439c81, 32'h3e5e2a18} /* (11, 20, 4) {real, imag} */,
  {32'hbe7df11e, 32'hbee46e74} /* (11, 20, 3) {real, imag} */,
  {32'hbee4309e, 32'h3e3e6c70} /* (11, 20, 2) {real, imag} */,
  {32'h3e4672de, 32'hbf04bc29} /* (11, 20, 1) {real, imag} */,
  {32'hbe61425c, 32'hbc50e4b0} /* (11, 20, 0) {real, imag} */,
  {32'h3d15c668, 32'hbd911c0a} /* (11, 19, 31) {real, imag} */,
  {32'hbe11c23a, 32'hbe1daca4} /* (11, 19, 30) {real, imag} */,
  {32'hbe24eb29, 32'h3e01f15a} /* (11, 19, 29) {real, imag} */,
  {32'hbd50df80, 32'hbeac2f2f} /* (11, 19, 28) {real, imag} */,
  {32'hbe4373d7, 32'h3e5fb4b8} /* (11, 19, 27) {real, imag} */,
  {32'hbd9a6f36, 32'h3daae0e8} /* (11, 19, 26) {real, imag} */,
  {32'h3d16e688, 32'hbe05a003} /* (11, 19, 25) {real, imag} */,
  {32'hbe621b77, 32'h3dcd0250} /* (11, 19, 24) {real, imag} */,
  {32'hbe9230ce, 32'h3d0392b0} /* (11, 19, 23) {real, imag} */,
  {32'hbe86a2ba, 32'hbe051f84} /* (11, 19, 22) {real, imag} */,
  {32'hbe817d07, 32'h3d94afd8} /* (11, 19, 21) {real, imag} */,
  {32'hbbf3b080, 32'h3ec0da66} /* (11, 19, 20) {real, imag} */,
  {32'h3dd805d4, 32'hbe8c3366} /* (11, 19, 19) {real, imag} */,
  {32'h3d90f658, 32'hbecbe1c0} /* (11, 19, 18) {real, imag} */,
  {32'hbcc1dc32, 32'h3ed2f052} /* (11, 19, 17) {real, imag} */,
  {32'hbebd39f7, 32'hbe1a6498} /* (11, 19, 16) {real, imag} */,
  {32'hbc9baa30, 32'hbcd957c0} /* (11, 19, 15) {real, imag} */,
  {32'hbe30363a, 32'h3e061102} /* (11, 19, 14) {real, imag} */,
  {32'hbd6e6358, 32'hbedb616f} /* (11, 19, 13) {real, imag} */,
  {32'hbef622fd, 32'h3f573804} /* (11, 19, 12) {real, imag} */,
  {32'h3d8ac154, 32'hbe9d95f8} /* (11, 19, 11) {real, imag} */,
  {32'hbd8c0820, 32'h3e4362a9} /* (11, 19, 10) {real, imag} */,
  {32'h3f2b6688, 32'hbe189d22} /* (11, 19, 9) {real, imag} */,
  {32'hbd4b059a, 32'h3ed6c84e} /* (11, 19, 8) {real, imag} */,
  {32'h3de94022, 32'h3f100edf} /* (11, 19, 7) {real, imag} */,
  {32'hbee889f8, 32'h3e636d4f} /* (11, 19, 6) {real, imag} */,
  {32'h3dc01413, 32'hbd590f24} /* (11, 19, 5) {real, imag} */,
  {32'h3ef6718e, 32'hbeab1a06} /* (11, 19, 4) {real, imag} */,
  {32'h3e9e3c0c, 32'hbd1fc780} /* (11, 19, 3) {real, imag} */,
  {32'hbdd42f68, 32'hbddfacf6} /* (11, 19, 2) {real, imag} */,
  {32'hbd912bbe, 32'h3f16aa90} /* (11, 19, 1) {real, imag} */,
  {32'h3e288106, 32'hbe942a72} /* (11, 19, 0) {real, imag} */,
  {32'h3d95ef78, 32'h3f36066c} /* (11, 18, 31) {real, imag} */,
  {32'h3ed46afe, 32'hbd35a16e} /* (11, 18, 30) {real, imag} */,
  {32'hbe4ee6a6, 32'h3e8d9c2b} /* (11, 18, 29) {real, imag} */,
  {32'hbec21abb, 32'h3e095554} /* (11, 18, 28) {real, imag} */,
  {32'h3dfa3fae, 32'hbe202af8} /* (11, 18, 27) {real, imag} */,
  {32'hbe578ec7, 32'hbde1b9ea} /* (11, 18, 26) {real, imag} */,
  {32'hbe5f56e1, 32'h3daa17d7} /* (11, 18, 25) {real, imag} */,
  {32'h3e0f5067, 32'hbe911576} /* (11, 18, 24) {real, imag} */,
  {32'hbdc09792, 32'hbe6391d0} /* (11, 18, 23) {real, imag} */,
  {32'h3f218260, 32'hbf62ded8} /* (11, 18, 22) {real, imag} */,
  {32'hbe2a871c, 32'hbe53b42c} /* (11, 18, 21) {real, imag} */,
  {32'hbf20be93, 32'hbd3f45f0} /* (11, 18, 20) {real, imag} */,
  {32'h3cc554ba, 32'h3d4d2a28} /* (11, 18, 19) {real, imag} */,
  {32'h3d256a10, 32'hbc2fee50} /* (11, 18, 18) {real, imag} */,
  {32'hbe0de419, 32'hbeb8bd86} /* (11, 18, 17) {real, imag} */,
  {32'hbea80a04, 32'hbdb780e8} /* (11, 18, 16) {real, imag} */,
  {32'h3e814dcc, 32'hbeb1108e} /* (11, 18, 15) {real, imag} */,
  {32'hbe4a3592, 32'h3e9d602a} /* (11, 18, 14) {real, imag} */,
  {32'h3d16892c, 32'h3ec5f1f9} /* (11, 18, 13) {real, imag} */,
  {32'hbe81937c, 32'h3e600c7e} /* (11, 18, 12) {real, imag} */,
  {32'h3ea72d1c, 32'hbe2d5542} /* (11, 18, 11) {real, imag} */,
  {32'h3d7b0e5c, 32'hbe706a8c} /* (11, 18, 10) {real, imag} */,
  {32'hbc401cf8, 32'h3d7466c6} /* (11, 18, 9) {real, imag} */,
  {32'hbc38d630, 32'hbc5c4af0} /* (11, 18, 8) {real, imag} */,
  {32'h3d93bd2e, 32'h3db662ba} /* (11, 18, 7) {real, imag} */,
  {32'hbdf88ba6, 32'h3d86c544} /* (11, 18, 6) {real, imag} */,
  {32'h3d05a945, 32'h3eeedaa0} /* (11, 18, 5) {real, imag} */,
  {32'hbebe4a8b, 32'hbed2f601} /* (11, 18, 4) {real, imag} */,
  {32'hbe89f2de, 32'hbe861db8} /* (11, 18, 3) {real, imag} */,
  {32'hbe8451c0, 32'hbede4891} /* (11, 18, 2) {real, imag} */,
  {32'hbea3e667, 32'h3e8f57ad} /* (11, 18, 1) {real, imag} */,
  {32'hbc631000, 32'h3ea6cb40} /* (11, 18, 0) {real, imag} */,
  {32'hbe67d8ea, 32'hbdef4b10} /* (11, 17, 31) {real, imag} */,
  {32'h3e9cb621, 32'h3e5bb5ce} /* (11, 17, 30) {real, imag} */,
  {32'h3ea3adf0, 32'hbcc2ec2c} /* (11, 17, 29) {real, imag} */,
  {32'hbf1a87e6, 32'h3e6e0ab2} /* (11, 17, 28) {real, imag} */,
  {32'hbd27d0a8, 32'hbe3aedf7} /* (11, 17, 27) {real, imag} */,
  {32'hbd3f304e, 32'hbd9b66c2} /* (11, 17, 26) {real, imag} */,
  {32'h3d0fa0da, 32'h3e8dbeef} /* (11, 17, 25) {real, imag} */,
  {32'h3edf3b0b, 32'hbe5da07c} /* (11, 17, 24) {real, imag} */,
  {32'hbcd46b20, 32'hbe836108} /* (11, 17, 23) {real, imag} */,
  {32'hbe9c8eea, 32'h3b97c360} /* (11, 17, 22) {real, imag} */,
  {32'hbf166a3b, 32'h3e5f9263} /* (11, 17, 21) {real, imag} */,
  {32'h3e447840, 32'h3e72808d} /* (11, 17, 20) {real, imag} */,
  {32'h3e6ac7d1, 32'hbcfd0278} /* (11, 17, 19) {real, imag} */,
  {32'h3e4a2a56, 32'h3ec9b688} /* (11, 17, 18) {real, imag} */,
  {32'h3dc467b8, 32'hbd570918} /* (11, 17, 17) {real, imag} */,
  {32'hbebac271, 32'hbe4ed706} /* (11, 17, 16) {real, imag} */,
  {32'h3cac8b08, 32'hbe11a62c} /* (11, 17, 15) {real, imag} */,
  {32'hbd9648c8, 32'h3c8cf8c0} /* (11, 17, 14) {real, imag} */,
  {32'hbed019c3, 32'h3e14c8d8} /* (11, 17, 13) {real, imag} */,
  {32'hbe333a3e, 32'h3f26a527} /* (11, 17, 12) {real, imag} */,
  {32'hbe0bbcbe, 32'h3e6e97b9} /* (11, 17, 11) {real, imag} */,
  {32'hbef3654e, 32'h3e5c453b} /* (11, 17, 10) {real, imag} */,
  {32'hbd888dfb, 32'h3998c400} /* (11, 17, 9) {real, imag} */,
  {32'hbd9f7f29, 32'hbe7ff7a0} /* (11, 17, 8) {real, imag} */,
  {32'hbedeb238, 32'hbdb6dd46} /* (11, 17, 7) {real, imag} */,
  {32'h3f155488, 32'hbda694d9} /* (11, 17, 6) {real, imag} */,
  {32'hbe7909a4, 32'hbe99c4c0} /* (11, 17, 5) {real, imag} */,
  {32'h3ebd2a3e, 32'hbe68a866} /* (11, 17, 4) {real, imag} */,
  {32'h3c8f490c, 32'h3daf6a65} /* (11, 17, 3) {real, imag} */,
  {32'h3e1e65d0, 32'hbd8f4217} /* (11, 17, 2) {real, imag} */,
  {32'hbe0aa525, 32'hbe54fd9a} /* (11, 17, 1) {real, imag} */,
  {32'h3e04a3d0, 32'hbe38b3b6} /* (11, 17, 0) {real, imag} */,
  {32'hbd16f33c, 32'h3dee0960} /* (11, 16, 31) {real, imag} */,
  {32'hbe352dba, 32'h3aa9de80} /* (11, 16, 30) {real, imag} */,
  {32'h3db54424, 32'h3eb7a8d0} /* (11, 16, 29) {real, imag} */,
  {32'h3d7f32f0, 32'h3e35080f} /* (11, 16, 28) {real, imag} */,
  {32'h3e2ace02, 32'hbe683f19} /* (11, 16, 27) {real, imag} */,
  {32'h3b55c140, 32'h3d00010a} /* (11, 16, 26) {real, imag} */,
  {32'h3c924c06, 32'hbe04cfde} /* (11, 16, 25) {real, imag} */,
  {32'h3d93e9a8, 32'hbde58e27} /* (11, 16, 24) {real, imag} */,
  {32'hbe0e808d, 32'hbdcd5fe9} /* (11, 16, 23) {real, imag} */,
  {32'h3db594ee, 32'h3ce68f1b} /* (11, 16, 22) {real, imag} */,
  {32'hbdcbd210, 32'h3c1bdff4} /* (11, 16, 21) {real, imag} */,
  {32'h3e1a6da4, 32'h3f12dd71} /* (11, 16, 20) {real, imag} */,
  {32'hbe05af36, 32'h3e41d001} /* (11, 16, 19) {real, imag} */,
  {32'h3e3264de, 32'h3e35fd6d} /* (11, 16, 18) {real, imag} */,
  {32'h3dbb9cae, 32'hbe534d36} /* (11, 16, 17) {real, imag} */,
  {32'h3e0e5488, 32'h00000000} /* (11, 16, 16) {real, imag} */,
  {32'h3dbb9cae, 32'h3e534d36} /* (11, 16, 15) {real, imag} */,
  {32'h3e3264de, 32'hbe35fd6d} /* (11, 16, 14) {real, imag} */,
  {32'hbe05af36, 32'hbe41d001} /* (11, 16, 13) {real, imag} */,
  {32'h3e1a6da4, 32'hbf12dd71} /* (11, 16, 12) {real, imag} */,
  {32'hbdcbd210, 32'hbc1bdff4} /* (11, 16, 11) {real, imag} */,
  {32'h3db594ee, 32'hbce68f1b} /* (11, 16, 10) {real, imag} */,
  {32'hbe0e808d, 32'h3dcd5fe9} /* (11, 16, 9) {real, imag} */,
  {32'h3d93e9a8, 32'h3de58e27} /* (11, 16, 8) {real, imag} */,
  {32'h3c924c06, 32'h3e04cfde} /* (11, 16, 7) {real, imag} */,
  {32'h3b55c140, 32'hbd00010a} /* (11, 16, 6) {real, imag} */,
  {32'h3e2ace02, 32'h3e683f19} /* (11, 16, 5) {real, imag} */,
  {32'h3d7f32f0, 32'hbe35080f} /* (11, 16, 4) {real, imag} */,
  {32'h3db54424, 32'hbeb7a8d0} /* (11, 16, 3) {real, imag} */,
  {32'hbe352dba, 32'hbaa9de80} /* (11, 16, 2) {real, imag} */,
  {32'hbd16f33c, 32'hbdee0960} /* (11, 16, 1) {real, imag} */,
  {32'hbded7256, 32'h00000000} /* (11, 16, 0) {real, imag} */,
  {32'hbe0aa525, 32'h3e54fd9a} /* (11, 15, 31) {real, imag} */,
  {32'h3e1e65d0, 32'h3d8f4217} /* (11, 15, 30) {real, imag} */,
  {32'h3c8f490c, 32'hbdaf6a65} /* (11, 15, 29) {real, imag} */,
  {32'h3ebd2a3e, 32'h3e68a866} /* (11, 15, 28) {real, imag} */,
  {32'hbe7909a4, 32'h3e99c4c0} /* (11, 15, 27) {real, imag} */,
  {32'h3f155488, 32'h3da694d9} /* (11, 15, 26) {real, imag} */,
  {32'hbedeb238, 32'h3db6dd46} /* (11, 15, 25) {real, imag} */,
  {32'hbd9f7f29, 32'h3e7ff7a0} /* (11, 15, 24) {real, imag} */,
  {32'hbd888dfb, 32'hb998c400} /* (11, 15, 23) {real, imag} */,
  {32'hbef3654e, 32'hbe5c453b} /* (11, 15, 22) {real, imag} */,
  {32'hbe0bbcbe, 32'hbe6e97b9} /* (11, 15, 21) {real, imag} */,
  {32'hbe333a3e, 32'hbf26a527} /* (11, 15, 20) {real, imag} */,
  {32'hbed019c3, 32'hbe14c8d8} /* (11, 15, 19) {real, imag} */,
  {32'hbd9648c8, 32'hbc8cf8c0} /* (11, 15, 18) {real, imag} */,
  {32'h3cac8b08, 32'h3e11a62c} /* (11, 15, 17) {real, imag} */,
  {32'hbebac271, 32'h3e4ed706} /* (11, 15, 16) {real, imag} */,
  {32'h3dc467b8, 32'h3d570918} /* (11, 15, 15) {real, imag} */,
  {32'h3e4a2a56, 32'hbec9b688} /* (11, 15, 14) {real, imag} */,
  {32'h3e6ac7d1, 32'h3cfd0278} /* (11, 15, 13) {real, imag} */,
  {32'h3e447840, 32'hbe72808d} /* (11, 15, 12) {real, imag} */,
  {32'hbf166a3b, 32'hbe5f9263} /* (11, 15, 11) {real, imag} */,
  {32'hbe9c8eea, 32'hbb97c360} /* (11, 15, 10) {real, imag} */,
  {32'hbcd46b20, 32'h3e836108} /* (11, 15, 9) {real, imag} */,
  {32'h3edf3b0b, 32'h3e5da07c} /* (11, 15, 8) {real, imag} */,
  {32'h3d0fa0da, 32'hbe8dbeef} /* (11, 15, 7) {real, imag} */,
  {32'hbd3f304e, 32'h3d9b66c2} /* (11, 15, 6) {real, imag} */,
  {32'hbd27d0a8, 32'h3e3aedf7} /* (11, 15, 5) {real, imag} */,
  {32'hbf1a87e6, 32'hbe6e0ab2} /* (11, 15, 4) {real, imag} */,
  {32'h3ea3adf0, 32'h3cc2ec2c} /* (11, 15, 3) {real, imag} */,
  {32'h3e9cb621, 32'hbe5bb5ce} /* (11, 15, 2) {real, imag} */,
  {32'hbe67d8ea, 32'h3def4b10} /* (11, 15, 1) {real, imag} */,
  {32'h3e04a3d0, 32'h3e38b3b6} /* (11, 15, 0) {real, imag} */,
  {32'hbea3e667, 32'hbe8f57ad} /* (11, 14, 31) {real, imag} */,
  {32'hbe8451c0, 32'h3ede4891} /* (11, 14, 30) {real, imag} */,
  {32'hbe89f2de, 32'h3e861db8} /* (11, 14, 29) {real, imag} */,
  {32'hbebe4a8b, 32'h3ed2f601} /* (11, 14, 28) {real, imag} */,
  {32'h3d05a945, 32'hbeeedaa0} /* (11, 14, 27) {real, imag} */,
  {32'hbdf88ba6, 32'hbd86c544} /* (11, 14, 26) {real, imag} */,
  {32'h3d93bd2e, 32'hbdb662ba} /* (11, 14, 25) {real, imag} */,
  {32'hbc38d630, 32'h3c5c4af0} /* (11, 14, 24) {real, imag} */,
  {32'hbc401cf8, 32'hbd7466c6} /* (11, 14, 23) {real, imag} */,
  {32'h3d7b0e5c, 32'h3e706a8c} /* (11, 14, 22) {real, imag} */,
  {32'h3ea72d1c, 32'h3e2d5542} /* (11, 14, 21) {real, imag} */,
  {32'hbe81937c, 32'hbe600c7e} /* (11, 14, 20) {real, imag} */,
  {32'h3d16892c, 32'hbec5f1f9} /* (11, 14, 19) {real, imag} */,
  {32'hbe4a3592, 32'hbe9d602a} /* (11, 14, 18) {real, imag} */,
  {32'h3e814dcc, 32'h3eb1108e} /* (11, 14, 17) {real, imag} */,
  {32'hbea80a04, 32'h3db780e8} /* (11, 14, 16) {real, imag} */,
  {32'hbe0de419, 32'h3eb8bd86} /* (11, 14, 15) {real, imag} */,
  {32'h3d256a10, 32'h3c2fee50} /* (11, 14, 14) {real, imag} */,
  {32'h3cc554ba, 32'hbd4d2a28} /* (11, 14, 13) {real, imag} */,
  {32'hbf20be93, 32'h3d3f45f0} /* (11, 14, 12) {real, imag} */,
  {32'hbe2a871c, 32'h3e53b42c} /* (11, 14, 11) {real, imag} */,
  {32'h3f218260, 32'h3f62ded8} /* (11, 14, 10) {real, imag} */,
  {32'hbdc09792, 32'h3e6391d0} /* (11, 14, 9) {real, imag} */,
  {32'h3e0f5067, 32'h3e911576} /* (11, 14, 8) {real, imag} */,
  {32'hbe5f56e1, 32'hbdaa17d7} /* (11, 14, 7) {real, imag} */,
  {32'hbe578ec7, 32'h3de1b9ea} /* (11, 14, 6) {real, imag} */,
  {32'h3dfa3fae, 32'h3e202af8} /* (11, 14, 5) {real, imag} */,
  {32'hbec21abb, 32'hbe095554} /* (11, 14, 4) {real, imag} */,
  {32'hbe4ee6a6, 32'hbe8d9c2b} /* (11, 14, 3) {real, imag} */,
  {32'h3ed46afe, 32'h3d35a16e} /* (11, 14, 2) {real, imag} */,
  {32'h3d95ef78, 32'hbf36066c} /* (11, 14, 1) {real, imag} */,
  {32'hbc631000, 32'hbea6cb40} /* (11, 14, 0) {real, imag} */,
  {32'hbd912bbe, 32'hbf16aa90} /* (11, 13, 31) {real, imag} */,
  {32'hbdd42f68, 32'h3ddfacf6} /* (11, 13, 30) {real, imag} */,
  {32'h3e9e3c0c, 32'h3d1fc780} /* (11, 13, 29) {real, imag} */,
  {32'h3ef6718e, 32'h3eab1a06} /* (11, 13, 28) {real, imag} */,
  {32'h3dc01413, 32'h3d590f24} /* (11, 13, 27) {real, imag} */,
  {32'hbee889f8, 32'hbe636d4f} /* (11, 13, 26) {real, imag} */,
  {32'h3de94022, 32'hbf100edf} /* (11, 13, 25) {real, imag} */,
  {32'hbd4b059a, 32'hbed6c84e} /* (11, 13, 24) {real, imag} */,
  {32'h3f2b6688, 32'h3e189d22} /* (11, 13, 23) {real, imag} */,
  {32'hbd8c0820, 32'hbe4362a9} /* (11, 13, 22) {real, imag} */,
  {32'h3d8ac154, 32'h3e9d95f8} /* (11, 13, 21) {real, imag} */,
  {32'hbef622fd, 32'hbf573804} /* (11, 13, 20) {real, imag} */,
  {32'hbd6e6358, 32'h3edb616f} /* (11, 13, 19) {real, imag} */,
  {32'hbe30363a, 32'hbe061102} /* (11, 13, 18) {real, imag} */,
  {32'hbc9baa30, 32'h3cd957c0} /* (11, 13, 17) {real, imag} */,
  {32'hbebd39f7, 32'h3e1a6498} /* (11, 13, 16) {real, imag} */,
  {32'hbcc1dc32, 32'hbed2f052} /* (11, 13, 15) {real, imag} */,
  {32'h3d90f658, 32'h3ecbe1c0} /* (11, 13, 14) {real, imag} */,
  {32'h3dd805d4, 32'h3e8c3366} /* (11, 13, 13) {real, imag} */,
  {32'hbbf3b080, 32'hbec0da66} /* (11, 13, 12) {real, imag} */,
  {32'hbe817d07, 32'hbd94afd8} /* (11, 13, 11) {real, imag} */,
  {32'hbe86a2ba, 32'h3e051f84} /* (11, 13, 10) {real, imag} */,
  {32'hbe9230ce, 32'hbd0392b0} /* (11, 13, 9) {real, imag} */,
  {32'hbe621b77, 32'hbdcd0250} /* (11, 13, 8) {real, imag} */,
  {32'h3d16e688, 32'h3e05a003} /* (11, 13, 7) {real, imag} */,
  {32'hbd9a6f36, 32'hbdaae0e8} /* (11, 13, 6) {real, imag} */,
  {32'hbe4373d7, 32'hbe5fb4b8} /* (11, 13, 5) {real, imag} */,
  {32'hbd50df80, 32'h3eac2f2f} /* (11, 13, 4) {real, imag} */,
  {32'hbe24eb29, 32'hbe01f15a} /* (11, 13, 3) {real, imag} */,
  {32'hbe11c23a, 32'h3e1daca4} /* (11, 13, 2) {real, imag} */,
  {32'h3d15c668, 32'h3d911c0a} /* (11, 13, 1) {real, imag} */,
  {32'h3e288106, 32'h3e942a72} /* (11, 13, 0) {real, imag} */,
  {32'h3e4672de, 32'h3f04bc29} /* (11, 12, 31) {real, imag} */,
  {32'hbee4309e, 32'hbe3e6c70} /* (11, 12, 30) {real, imag} */,
  {32'hbe7df11e, 32'h3ee46e74} /* (11, 12, 29) {real, imag} */,
  {32'hbe439c81, 32'hbe5e2a18} /* (11, 12, 28) {real, imag} */,
  {32'hbc353f78, 32'hbee2c80d} /* (11, 12, 27) {real, imag} */,
  {32'h3e257376, 32'h3f0fdb31} /* (11, 12, 26) {real, imag} */,
  {32'h3e65d586, 32'h3e3ae68b} /* (11, 12, 25) {real, imag} */,
  {32'h3e958ee5, 32'hbc328be0} /* (11, 12, 24) {real, imag} */,
  {32'hbe86c1d8, 32'h3ec0a258} /* (11, 12, 23) {real, imag} */,
  {32'h3eac6647, 32'hbbd53848} /* (11, 12, 22) {real, imag} */,
  {32'hbf44d284, 32'h3da4c847} /* (11, 12, 21) {real, imag} */,
  {32'hbdeaa10f, 32'h3ebfd042} /* (11, 12, 20) {real, imag} */,
  {32'h3ceafb29, 32'h3d9bc556} /* (11, 12, 19) {real, imag} */,
  {32'hbeb72d10, 32'hbe565268} /* (11, 12, 18) {real, imag} */,
  {32'hbe07b7b6, 32'hbb81d900} /* (11, 12, 17) {real, imag} */,
  {32'hbccc20e0, 32'hbed24812} /* (11, 12, 16) {real, imag} */,
  {32'h3d9e775d, 32'h3d23f000} /* (11, 12, 15) {real, imag} */,
  {32'hbe878bea, 32'h3d03e6e8} /* (11, 12, 14) {real, imag} */,
  {32'hbe766565, 32'h3d537c0e} /* (11, 12, 13) {real, imag} */,
  {32'h3db20812, 32'h3eb841ec} /* (11, 12, 12) {real, imag} */,
  {32'h3c503760, 32'h3e89f1bb} /* (11, 12, 11) {real, imag} */,
  {32'h3e452cd5, 32'hbe55974e} /* (11, 12, 10) {real, imag} */,
  {32'hbf2121f3, 32'hbeca41b9} /* (11, 12, 9) {real, imag} */,
  {32'h3e6f5be3, 32'h3e9d7268} /* (11, 12, 8) {real, imag} */,
  {32'hbd6b6770, 32'hbf4c102a} /* (11, 12, 7) {real, imag} */,
  {32'h3e41ffaf, 32'hbe9ab223} /* (11, 12, 6) {real, imag} */,
  {32'hbe0ffabb, 32'hbee285c3} /* (11, 12, 5) {real, imag} */,
  {32'h3e738eff, 32'hbea772a9} /* (11, 12, 4) {real, imag} */,
  {32'h3e22d303, 32'h3e13375d} /* (11, 12, 3) {real, imag} */,
  {32'h3ef2e050, 32'h3f0d7f35} /* (11, 12, 2) {real, imag} */,
  {32'hbde3695b, 32'hbe15891c} /* (11, 12, 1) {real, imag} */,
  {32'hbe61425c, 32'h3c50e4b0} /* (11, 12, 0) {real, imag} */,
  {32'hbdb380c4, 32'hbefb3e32} /* (11, 11, 31) {real, imag} */,
  {32'h3f79d3a5, 32'hbd14ec22} /* (11, 11, 30) {real, imag} */,
  {32'h3e07ed19, 32'hbe4f819d} /* (11, 11, 29) {real, imag} */,
  {32'hbe9de1f4, 32'h3ecfe524} /* (11, 11, 28) {real, imag} */,
  {32'hbd466ff4, 32'h3e3e0c47} /* (11, 11, 27) {real, imag} */,
  {32'hbedc2d73, 32'hbe98c248} /* (11, 11, 26) {real, imag} */,
  {32'h3e032bbc, 32'h3f0be722} /* (11, 11, 25) {real, imag} */,
  {32'h3eb3a3a4, 32'hbe712c23} /* (11, 11, 24) {real, imag} */,
  {32'hbef5e3d4, 32'hbed82d8b} /* (11, 11, 23) {real, imag} */,
  {32'hbcde28d8, 32'hbe9b4528} /* (11, 11, 22) {real, imag} */,
  {32'h3ebffb10, 32'h3dcce78f} /* (11, 11, 21) {real, imag} */,
  {32'h3eba9203, 32'h3dfffb18} /* (11, 11, 20) {real, imag} */,
  {32'hbebf1045, 32'h3eb77c16} /* (11, 11, 19) {real, imag} */,
  {32'hbe1deea0, 32'h3ee7038a} /* (11, 11, 18) {real, imag} */,
  {32'h3dcb7bc2, 32'hbc8a608c} /* (11, 11, 17) {real, imag} */,
  {32'h3de6e886, 32'h3eabbf1b} /* (11, 11, 16) {real, imag} */,
  {32'hbda50bf2, 32'hbe5c7f05} /* (11, 11, 15) {real, imag} */,
  {32'h3dab0bda, 32'hbe280de6} /* (11, 11, 14) {real, imag} */,
  {32'hbe5389a6, 32'h3e9e0c86} /* (11, 11, 13) {real, imag} */,
  {32'h3d9523e6, 32'hbdd734d8} /* (11, 11, 12) {real, imag} */,
  {32'hbe9e15db, 32'hbd8b6dbb} /* (11, 11, 11) {real, imag} */,
  {32'h3d5228dc, 32'hbe2c909c} /* (11, 11, 10) {real, imag} */,
  {32'h3f50c1f3, 32'hbea84b4a} /* (11, 11, 9) {real, imag} */,
  {32'h3ea075c7, 32'h3dd4866c} /* (11, 11, 8) {real, imag} */,
  {32'hbee5c47d, 32'h3f289a4a} /* (11, 11, 7) {real, imag} */,
  {32'h3e925f86, 32'hbe697029} /* (11, 11, 6) {real, imag} */,
  {32'h3e14d8cc, 32'h3f145781} /* (11, 11, 5) {real, imag} */,
  {32'h3f23fbab, 32'hbebd531d} /* (11, 11, 4) {real, imag} */,
  {32'hbe6b313e, 32'h3f3307cc} /* (11, 11, 3) {real, imag} */,
  {32'hbeb8ee30, 32'h3f9b35fa} /* (11, 11, 2) {real, imag} */,
  {32'hbd92ec86, 32'hbf1039a0} /* (11, 11, 1) {real, imag} */,
  {32'hbeb5545f, 32'hbf216ea7} /* (11, 11, 0) {real, imag} */,
  {32'h3ceb9808, 32'h3f521d4a} /* (11, 10, 31) {real, imag} */,
  {32'hbe1f7792, 32'h3c1538c0} /* (11, 10, 30) {real, imag} */,
  {32'hbdd5a50f, 32'hbeaa051c} /* (11, 10, 29) {real, imag} */,
  {32'h3f1455c2, 32'hbeaf83a5} /* (11, 10, 28) {real, imag} */,
  {32'hbf5c28b8, 32'hbd652cf4} /* (11, 10, 27) {real, imag} */,
  {32'h3da05897, 32'hbe5150f6} /* (11, 10, 26) {real, imag} */,
  {32'hbe6fc91f, 32'h3df0e1aa} /* (11, 10, 25) {real, imag} */,
  {32'hbe15afdb, 32'hbd9b9178} /* (11, 10, 24) {real, imag} */,
  {32'h3dfcda40, 32'h3eda0be4} /* (11, 10, 23) {real, imag} */,
  {32'hbdd52da9, 32'h3e1b4a54} /* (11, 10, 22) {real, imag} */,
  {32'h3e1afe57, 32'h3db590ef} /* (11, 10, 21) {real, imag} */,
  {32'hbda925b3, 32'h3e8c407c} /* (11, 10, 20) {real, imag} */,
  {32'hbdf9ffba, 32'hbe4a1133} /* (11, 10, 19) {real, imag} */,
  {32'h3b867e88, 32'hbf048862} /* (11, 10, 18) {real, imag} */,
  {32'h3f0e6d35, 32'h3f0a5b19} /* (11, 10, 17) {real, imag} */,
  {32'hbeb19682, 32'hbdb6da8c} /* (11, 10, 16) {real, imag} */,
  {32'hbe53228e, 32'h3e5a562f} /* (11, 10, 15) {real, imag} */,
  {32'h3e2bbcd6, 32'hb9b03700} /* (11, 10, 14) {real, imag} */,
  {32'h3db092fd, 32'h3e9dc1d2} /* (11, 10, 13) {real, imag} */,
  {32'hbd0e4ae4, 32'hbd89aee4} /* (11, 10, 12) {real, imag} */,
  {32'h3ca2d1e0, 32'hbc6a53ec} /* (11, 10, 11) {real, imag} */,
  {32'hbd06bd9c, 32'hbf1387fd} /* (11, 10, 10) {real, imag} */,
  {32'h3eeaf9ec, 32'h3e831f08} /* (11, 10, 9) {real, imag} */,
  {32'hbd082b3e, 32'hbe48ed3e} /* (11, 10, 8) {real, imag} */,
  {32'hbe7268c6, 32'hbd98f59f} /* (11, 10, 7) {real, imag} */,
  {32'h3e7a3b61, 32'hbf2e1520} /* (11, 10, 6) {real, imag} */,
  {32'h3f53c16c, 32'hbe9bd967} /* (11, 10, 5) {real, imag} */,
  {32'h3ebdd00e, 32'h3f5dffd4} /* (11, 10, 4) {real, imag} */,
  {32'h3d22fa94, 32'h3efe02ba} /* (11, 10, 3) {real, imag} */,
  {32'h3e98ce9f, 32'hbedf67af} /* (11, 10, 2) {real, imag} */,
  {32'hbe20c462, 32'h3f537303} /* (11, 10, 1) {real, imag} */,
  {32'h3e865a20, 32'hbf1f1d5c} /* (11, 10, 0) {real, imag} */,
  {32'hbf984f52, 32'h3f04d277} /* (11, 9, 31) {real, imag} */,
  {32'h3ecd0668, 32'hbf1ccfe2} /* (11, 9, 30) {real, imag} */,
  {32'h3e901d72, 32'h3d1d8090} /* (11, 9, 29) {real, imag} */,
  {32'hbe095366, 32'hbdf8bf2c} /* (11, 9, 28) {real, imag} */,
  {32'hbe8c7099, 32'h3d8061ee} /* (11, 9, 27) {real, imag} */,
  {32'h3ef86a6f, 32'hbedde02e} /* (11, 9, 26) {real, imag} */,
  {32'h3bde8d80, 32'h3eb241a2} /* (11, 9, 25) {real, imag} */,
  {32'h3e607521, 32'h3ef464f5} /* (11, 9, 24) {real, imag} */,
  {32'hbe07df60, 32'h3ea8f6ba} /* (11, 9, 23) {real, imag} */,
  {32'hbe207753, 32'hbf44f3b6} /* (11, 9, 22) {real, imag} */,
  {32'hbeaad22d, 32'hbec18e8c} /* (11, 9, 21) {real, imag} */,
  {32'h3e0282d8, 32'h3ecbb1ab} /* (11, 9, 20) {real, imag} */,
  {32'h3f86eaa8, 32'hbe865e67} /* (11, 9, 19) {real, imag} */,
  {32'hbb897f40, 32'h3e8dbfaa} /* (11, 9, 18) {real, imag} */,
  {32'hbdc2613f, 32'h3e256aea} /* (11, 9, 17) {real, imag} */,
  {32'hbe09bd6c, 32'hbdead762} /* (11, 9, 16) {real, imag} */,
  {32'hbdcf503f, 32'h3ad2cfc0} /* (11, 9, 15) {real, imag} */,
  {32'h3c08e448, 32'h3d0f42a4} /* (11, 9, 14) {real, imag} */,
  {32'hbf3ff504, 32'hbe95b854} /* (11, 9, 13) {real, imag} */,
  {32'h3eb4be96, 32'hbf2f811e} /* (11, 9, 12) {real, imag} */,
  {32'hbe81576e, 32'h3c5522d0} /* (11, 9, 11) {real, imag} */,
  {32'hbea8e8e6, 32'h3f09faa8} /* (11, 9, 10) {real, imag} */,
  {32'h3d90ead4, 32'h3f3fa93a} /* (11, 9, 9) {real, imag} */,
  {32'hbebe460c, 32'hbf0ec476} /* (11, 9, 8) {real, imag} */,
  {32'hbdddc92d, 32'hbf1799ac} /* (11, 9, 7) {real, imag} */,
  {32'h3dbc9064, 32'h3dad84bc} /* (11, 9, 6) {real, imag} */,
  {32'h3dc0ac38, 32'h3d402a8c} /* (11, 9, 5) {real, imag} */,
  {32'hbf1b5f7a, 32'h3cc6ec5c} /* (11, 9, 4) {real, imag} */,
  {32'h3eb69645, 32'hbeca50e5} /* (11, 9, 3) {real, imag} */,
  {32'hbdac88ba, 32'hbf4a0b98} /* (11, 9, 2) {real, imag} */,
  {32'h3e70aee9, 32'h3f1c7f16} /* (11, 9, 1) {real, imag} */,
  {32'h3d3538c0, 32'hbd70d664} /* (11, 9, 0) {real, imag} */,
  {32'hbfda8b79, 32'hbf751222} /* (11, 8, 31) {real, imag} */,
  {32'h3f898232, 32'hbe677cc2} /* (11, 8, 30) {real, imag} */,
  {32'hbf89217c, 32'h3deabc1e} /* (11, 8, 29) {real, imag} */,
  {32'h3ec76264, 32'h3e9808f9} /* (11, 8, 28) {real, imag} */,
  {32'h3cdaabb0, 32'hbe9da75e} /* (11, 8, 27) {real, imag} */,
  {32'h3d0d93e8, 32'h3fa38c64} /* (11, 8, 26) {real, imag} */,
  {32'h3e912d4e, 32'hbf3ef202} /* (11, 8, 25) {real, imag} */,
  {32'hbefe0448, 32'hbeae5000} /* (11, 8, 24) {real, imag} */,
  {32'h3e01bd6e, 32'h3c886570} /* (11, 8, 23) {real, imag} */,
  {32'h3f212279, 32'h3da445e2} /* (11, 8, 22) {real, imag} */,
  {32'h3e3e4f85, 32'hbe36f008} /* (11, 8, 21) {real, imag} */,
  {32'h3f05e238, 32'h3e09b4d3} /* (11, 8, 20) {real, imag} */,
  {32'hbd02f46f, 32'hbd512ee8} /* (11, 8, 19) {real, imag} */,
  {32'h3e98ede9, 32'h3d0b25cc} /* (11, 8, 18) {real, imag} */,
  {32'hbdc52532, 32'h3e395ec6} /* (11, 8, 17) {real, imag} */,
  {32'hbc5ec990, 32'h3dae279a} /* (11, 8, 16) {real, imag} */,
  {32'hbf0f04f8, 32'h3d94091a} /* (11, 8, 15) {real, imag} */,
  {32'h3ed3b056, 32'h3eb773e8} /* (11, 8, 14) {real, imag} */,
  {32'hbe4dceea, 32'hbe378920} /* (11, 8, 13) {real, imag} */,
  {32'h3eb833d1, 32'hbefa3d9e} /* (11, 8, 12) {real, imag} */,
  {32'hbe44d19c, 32'h3f02e78f} /* (11, 8, 11) {real, imag} */,
  {32'h3e63c7f9, 32'h3ee47665} /* (11, 8, 10) {real, imag} */,
  {32'hbed5ce7a, 32'hbf011965} /* (11, 8, 9) {real, imag} */,
  {32'hbeddd500, 32'hbdadc656} /* (11, 8, 8) {real, imag} */,
  {32'hbf215946, 32'hbe9bf3ab} /* (11, 8, 7) {real, imag} */,
  {32'h3e6f565e, 32'h3edbfcbf} /* (11, 8, 6) {real, imag} */,
  {32'h3d741750, 32'h3ea874d9} /* (11, 8, 5) {real, imag} */,
  {32'hbf80dcdc, 32'hbe6926af} /* (11, 8, 4) {real, imag} */,
  {32'hbdf0239e, 32'hbe7c8c1d} /* (11, 8, 3) {real, imag} */,
  {32'h3f953914, 32'h3f2dfb5d} /* (11, 8, 2) {real, imag} */,
  {32'hbf84a9f2, 32'hbeb331fa} /* (11, 8, 1) {real, imag} */,
  {32'h3d510ab4, 32'hbf1e97e1} /* (11, 8, 0) {real, imag} */,
  {32'h3f2d2a66, 32'h3e9a4ffc} /* (11, 7, 31) {real, imag} */,
  {32'hbe8cbe28, 32'h3d1c4440} /* (11, 7, 30) {real, imag} */,
  {32'h3eec3f48, 32'h3ead2d1a} /* (11, 7, 29) {real, imag} */,
  {32'hbe2f5151, 32'h3e5eb02a} /* (11, 7, 28) {real, imag} */,
  {32'h3ea651bb, 32'h3ea1b3fe} /* (11, 7, 27) {real, imag} */,
  {32'hbea12222, 32'hbdf766e0} /* (11, 7, 26) {real, imag} */,
  {32'h3f1e7bb1, 32'hbbdfcf80} /* (11, 7, 25) {real, imag} */,
  {32'hbf7d756e, 32'hbeca1301} /* (11, 7, 24) {real, imag} */,
  {32'hbedf1173, 32'h3ea355d0} /* (11, 7, 23) {real, imag} */,
  {32'hbe168f50, 32'h3ec70a82} /* (11, 7, 22) {real, imag} */,
  {32'h3e9e146e, 32'h3ef2cda1} /* (11, 7, 21) {real, imag} */,
  {32'h3e0ee328, 32'h3d2431d7} /* (11, 7, 20) {real, imag} */,
  {32'h3f1a8ff8, 32'h3f83f69d} /* (11, 7, 19) {real, imag} */,
  {32'hbea36167, 32'h3cbecba8} /* (11, 7, 18) {real, imag} */,
  {32'hbe19e815, 32'hbe9055f4} /* (11, 7, 17) {real, imag} */,
  {32'hbe8c16fe, 32'h3ec322db} /* (11, 7, 16) {real, imag} */,
  {32'hbde92234, 32'h3dc99aee} /* (11, 7, 15) {real, imag} */,
  {32'hbe057f89, 32'hbd506940} /* (11, 7, 14) {real, imag} */,
  {32'hbe3237b0, 32'h3e9fc0a6} /* (11, 7, 13) {real, imag} */,
  {32'hbe422bf9, 32'hbdfc8c97} /* (11, 7, 12) {real, imag} */,
  {32'h3e9414b0, 32'hbdf14dfa} /* (11, 7, 11) {real, imag} */,
  {32'h3ed14df9, 32'h3e529eee} /* (11, 7, 10) {real, imag} */,
  {32'hbdd3c95a, 32'hbd256820} /* (11, 7, 9) {real, imag} */,
  {32'h3ef76976, 32'hbe005d6e} /* (11, 7, 8) {real, imag} */,
  {32'h3e646a5a, 32'h3f09aafa} /* (11, 7, 7) {real, imag} */,
  {32'h3e91be26, 32'hbf833c4d} /* (11, 7, 6) {real, imag} */,
  {32'hbf4b1748, 32'hbde69f6a} /* (11, 7, 5) {real, imag} */,
  {32'h3f2e6631, 32'h3e33dd2e} /* (11, 7, 4) {real, imag} */,
  {32'h3d8b8ac8, 32'hbdee98b8} /* (11, 7, 3) {real, imag} */,
  {32'hbdea312c, 32'h3df8a121} /* (11, 7, 2) {real, imag} */,
  {32'hbde0d314, 32'h3e96a4fc} /* (11, 7, 1) {real, imag} */,
  {32'h3e9efa4e, 32'h3e815e98} /* (11, 7, 0) {real, imag} */,
  {32'h3f7382c9, 32'hbfa32261} /* (11, 6, 31) {real, imag} */,
  {32'h3caec7f0, 32'hbf1a41e2} /* (11, 6, 30) {real, imag} */,
  {32'h3e11186f, 32'hbed2a84f} /* (11, 6, 29) {real, imag} */,
  {32'h3ef13f90, 32'hbf83cec3} /* (11, 6, 28) {real, imag} */,
  {32'h3f271be8, 32'h3ca172e0} /* (11, 6, 27) {real, imag} */,
  {32'h3e9ccf90, 32'h3f4d0c5c} /* (11, 6, 26) {real, imag} */,
  {32'hbe3778a6, 32'hbea446f7} /* (11, 6, 25) {real, imag} */,
  {32'hbdaf5070, 32'h3f1b8af7} /* (11, 6, 24) {real, imag} */,
  {32'h3e64c837, 32'h3f27a0c4} /* (11, 6, 23) {real, imag} */,
  {32'h3ef72a30, 32'h3ea22b18} /* (11, 6, 22) {real, imag} */,
  {32'h3e1dd059, 32'h3ea02712} /* (11, 6, 21) {real, imag} */,
  {32'h3d1137b0, 32'hbe7d4931} /* (11, 6, 20) {real, imag} */,
  {32'hbe34c180, 32'h3ef721e5} /* (11, 6, 19) {real, imag} */,
  {32'hbe28c3f6, 32'h3e9c6a6e} /* (11, 6, 18) {real, imag} */,
  {32'h3e8eadfe, 32'hbed3b2f1} /* (11, 6, 17) {real, imag} */,
  {32'h3e1365f0, 32'h3d960636} /* (11, 6, 16) {real, imag} */,
  {32'hbd2420db, 32'h3d045aae} /* (11, 6, 15) {real, imag} */,
  {32'hbe3887f2, 32'h3e208380} /* (11, 6, 14) {real, imag} */,
  {32'h3cd834ba, 32'h3e739882} /* (11, 6, 13) {real, imag} */,
  {32'hbd44be28, 32'hbebd48fb} /* (11, 6, 12) {real, imag} */,
  {32'h3d128438, 32'hbf177d73} /* (11, 6, 11) {real, imag} */,
  {32'hbdbfbdf4, 32'h3e4e27d4} /* (11, 6, 10) {real, imag} */,
  {32'hbea1182b, 32'hbd8bfc3c} /* (11, 6, 9) {real, imag} */,
  {32'hbeb1b418, 32'hbf206d98} /* (11, 6, 8) {real, imag} */,
  {32'h3e30c996, 32'h3e438d3f} /* (11, 6, 7) {real, imag} */,
  {32'h3ee78efc, 32'hbe916e6f} /* (11, 6, 6) {real, imag} */,
  {32'h3dde31f8, 32'hbe7f9437} /* (11, 6, 5) {real, imag} */,
  {32'h3dd7e907, 32'h3d0121ee} /* (11, 6, 4) {real, imag} */,
  {32'h3eacf6ce, 32'h3ebb53ce} /* (11, 6, 3) {real, imag} */,
  {32'h3f3d3b27, 32'h3daec9d4} /* (11, 6, 2) {real, imag} */,
  {32'h3e496e12, 32'h3dfa914c} /* (11, 6, 1) {real, imag} */,
  {32'h3df8911e, 32'h3f19aa50} /* (11, 6, 0) {real, imag} */,
  {32'hc05d9576, 32'hbe022142} /* (11, 5, 31) {real, imag} */,
  {32'h3eb10ea8, 32'hbc455ca0} /* (11, 5, 30) {real, imag} */,
  {32'hbf2c5d22, 32'h3e405c8f} /* (11, 5, 29) {real, imag} */,
  {32'hbeff6a43, 32'h3fcc7d5a} /* (11, 5, 28) {real, imag} */,
  {32'h3eb895f0, 32'h3f1b62d4} /* (11, 5, 27) {real, imag} */,
  {32'h3ec4eb58, 32'hbe99232a} /* (11, 5, 26) {real, imag} */,
  {32'h3e287fe2, 32'hbdcd7b0d} /* (11, 5, 25) {real, imag} */,
  {32'h3eed21c6, 32'hbf954064} /* (11, 5, 24) {real, imag} */,
  {32'hbda6fa62, 32'hbe8064bc} /* (11, 5, 23) {real, imag} */,
  {32'h3df2929e, 32'h3e3d5cf2} /* (11, 5, 22) {real, imag} */,
  {32'hbe3b3320, 32'hbf0b8876} /* (11, 5, 21) {real, imag} */,
  {32'h3e5d3ebd, 32'h3b9af880} /* (11, 5, 20) {real, imag} */,
  {32'h3f13b0f3, 32'h3ed2a230} /* (11, 5, 19) {real, imag} */,
  {32'hbe6c6be4, 32'h3e2e0a89} /* (11, 5, 18) {real, imag} */,
  {32'h3c5b8f30, 32'h3d8f20ed} /* (11, 5, 17) {real, imag} */,
  {32'hbe66084e, 32'h3dd32214} /* (11, 5, 16) {real, imag} */,
  {32'h3e9ad574, 32'hbe469c88} /* (11, 5, 15) {real, imag} */,
  {32'hbe568376, 32'h3e5dd840} /* (11, 5, 14) {real, imag} */,
  {32'h3e993244, 32'h3e55e48a} /* (11, 5, 13) {real, imag} */,
  {32'h3e999806, 32'h3f21c47b} /* (11, 5, 12) {real, imag} */,
  {32'h3f27ecc2, 32'hbe97f42c} /* (11, 5, 11) {real, imag} */,
  {32'hbeec06de, 32'h3ebd5356} /* (11, 5, 10) {real, imag} */,
  {32'hbe5808dd, 32'hbe759015} /* (11, 5, 9) {real, imag} */,
  {32'h3f158817, 32'h3f3456b8} /* (11, 5, 8) {real, imag} */,
  {32'h3e457cf0, 32'h3ea66bd1} /* (11, 5, 7) {real, imag} */,
  {32'hbf86c45e, 32'hbce43060} /* (11, 5, 6) {real, imag} */,
  {32'h3f8c3aec, 32'hbae5d000} /* (11, 5, 5) {real, imag} */,
  {32'h3e3385ed, 32'hbe8fdb2b} /* (11, 5, 4) {real, imag} */,
  {32'hbf61aeae, 32'hbe9ab5d8} /* (11, 5, 3) {real, imag} */,
  {32'h3f1c603c, 32'h3f62af0e} /* (11, 5, 2) {real, imag} */,
  {32'hbed2afba, 32'hc01b86e8} /* (11, 5, 1) {real, imag} */,
  {32'hbfe523e2, 32'hbf33bf32} /* (11, 5, 0) {real, imag} */,
  {32'h3f712752, 32'h403171a3} /* (11, 4, 31) {real, imag} */,
  {32'hc06acd1f, 32'hc02eaad3} /* (11, 4, 30) {real, imag} */,
  {32'hbeaa0525, 32'hbed6b3d5} /* (11, 4, 29) {real, imag} */,
  {32'h3e2cb6dd, 32'hbd4c8da0} /* (11, 4, 28) {real, imag} */,
  {32'hbe172a33, 32'h3e867687} /* (11, 4, 27) {real, imag} */,
  {32'hbe5f84ac, 32'hbe192348} /* (11, 4, 26) {real, imag} */,
  {32'h3f192fcc, 32'h3e8f1535} /* (11, 4, 25) {real, imag} */,
  {32'hbd12162c, 32'hbe87a07a} /* (11, 4, 24) {real, imag} */,
  {32'h3f147f2e, 32'hbe9ab064} /* (11, 4, 23) {real, imag} */,
  {32'hbe7226ea, 32'hbe00b536} /* (11, 4, 22) {real, imag} */,
  {32'hbee0655e, 32'h3e19afab} /* (11, 4, 21) {real, imag} */,
  {32'h3f1d46bd, 32'h3e8f87bd} /* (11, 4, 20) {real, imag} */,
  {32'h3e3f2560, 32'h3e3cba06} /* (11, 4, 19) {real, imag} */,
  {32'hbe522f46, 32'hbf219aa7} /* (11, 4, 18) {real, imag} */,
  {32'h3e220678, 32'h3e1290b5} /* (11, 4, 17) {real, imag} */,
  {32'h3cde33e4, 32'h3e09c9a2} /* (11, 4, 16) {real, imag} */,
  {32'hbd54d751, 32'hbd8c8a8c} /* (11, 4, 15) {real, imag} */,
  {32'h3eb47fd0, 32'hbed4a1c6} /* (11, 4, 14) {real, imag} */,
  {32'hbdbd8d3c, 32'h3d05ca08} /* (11, 4, 13) {real, imag} */,
  {32'h3e174fb1, 32'h3d36711f} /* (11, 4, 12) {real, imag} */,
  {32'h3da61298, 32'hbe0a158f} /* (11, 4, 11) {real, imag} */,
  {32'hbf2c3ae6, 32'hbe1685fd} /* (11, 4, 10) {real, imag} */,
  {32'hbe6fe966, 32'h3ea02c9a} /* (11, 4, 9) {real, imag} */,
  {32'hbf0470a1, 32'hbf1d0aa0} /* (11, 4, 8) {real, imag} */,
  {32'h3edd8def, 32'hbec6b910} /* (11, 4, 7) {real, imag} */,
  {32'hbee1ea33, 32'h3f4cde3e} /* (11, 4, 6) {real, imag} */,
  {32'h3f144aaa, 32'hbf3d6c61} /* (11, 4, 5) {real, imag} */,
  {32'h3e0864dc, 32'h3f9d08d7} /* (11, 4, 4) {real, imag} */,
  {32'h3f44c972, 32'h3d0db810} /* (11, 4, 3) {real, imag} */,
  {32'hc025b734, 32'hbfeaf7c2} /* (11, 4, 2) {real, imag} */,
  {32'h40c08df8, 32'h3f9aa2ac} /* (11, 4, 1) {real, imag} */,
  {32'h3fb71a2a, 32'hbc53c900} /* (11, 4, 0) {real, imag} */,
  {32'hc08b19d8, 32'h40269cd3} /* (11, 3, 31) {real, imag} */,
  {32'h3ff5944e, 32'hc091ba98} /* (11, 3, 30) {real, imag} */,
  {32'hbf04aeb0, 32'h3df15d71} /* (11, 3, 29) {real, imag} */,
  {32'h3f9165ae, 32'h3fa3b7ce} /* (11, 3, 28) {real, imag} */,
  {32'hbf9c72a8, 32'h3f2b8ddc} /* (11, 3, 27) {real, imag} */,
  {32'h3ef68f00, 32'h3f3e8ddb} /* (11, 3, 26) {real, imag} */,
  {32'h3ed6db18, 32'h3ed4215b} /* (11, 3, 25) {real, imag} */,
  {32'h3efb6f24, 32'hbe854884} /* (11, 3, 24) {real, imag} */,
  {32'h3cf1a5d8, 32'hbf14ef0d} /* (11, 3, 23) {real, imag} */,
  {32'hbe24b3df, 32'h3d3cf700} /* (11, 3, 22) {real, imag} */,
  {32'h3ea2f6f6, 32'h3ed8ef20} /* (11, 3, 21) {real, imag} */,
  {32'h3de4c866, 32'h3dd47bf8} /* (11, 3, 20) {real, imag} */,
  {32'hbf07b2e5, 32'hbe014518} /* (11, 3, 19) {real, imag} */,
  {32'h3eb4affd, 32'hbda0026a} /* (11, 3, 18) {real, imag} */,
  {32'h3e3d38b9, 32'h3f041238} /* (11, 3, 17) {real, imag} */,
  {32'h3e3d5da3, 32'h3de1fd4c} /* (11, 3, 16) {real, imag} */,
  {32'hbebb24df, 32'h3e8e0241} /* (11, 3, 15) {real, imag} */,
  {32'h3ee76c87, 32'hbf251786} /* (11, 3, 14) {real, imag} */,
  {32'h3e6cedaa, 32'hbe086d88} /* (11, 3, 13) {real, imag} */,
  {32'hbe812b32, 32'h3de951ac} /* (11, 3, 12) {real, imag} */,
  {32'h3e88b0bc, 32'h3b0c3880} /* (11, 3, 11) {real, imag} */,
  {32'h3d1710a0, 32'h3e6d1b36} /* (11, 3, 10) {real, imag} */,
  {32'hbdf16e68, 32'h3dc1a13a} /* (11, 3, 9) {real, imag} */,
  {32'h3c1138e0, 32'hbe70f7d0} /* (11, 3, 8) {real, imag} */,
  {32'h3dcea700, 32'hbeeaf6a7} /* (11, 3, 7) {real, imag} */,
  {32'h3eabb0d2, 32'h3ef33f0e} /* (11, 3, 6) {real, imag} */,
  {32'hbe5c2517, 32'h3f045129} /* (11, 3, 5) {real, imag} */,
  {32'hbf70392a, 32'h3eaa3156} /* (11, 3, 4) {real, imag} */,
  {32'hbf6791f8, 32'h3f1ded94} /* (11, 3, 3) {real, imag} */,
  {32'h3e6a39a6, 32'hc03f8072} /* (11, 3, 2) {real, imag} */,
  {32'h407a8474, 32'h40384752} /* (11, 3, 1) {real, imag} */,
  {32'h3e5248fc, 32'h3ecf0fc0} /* (11, 3, 0) {real, imag} */,
  {32'hc222d3e7, 32'hc025fec6} /* (11, 2, 31) {real, imag} */,
  {32'h41946cf5, 32'hc0a9b6b9} /* (11, 2, 30) {real, imag} */,
  {32'h3ee63a8e, 32'h3f0f9b23} /* (11, 2, 29) {real, imag} */,
  {32'hbf1dab10, 32'h4015816a} /* (11, 2, 28) {real, imag} */,
  {32'h3fe5d2a9, 32'hbff8bc99} /* (11, 2, 27) {real, imag} */,
  {32'h3f2733b4, 32'h3d2e574c} /* (11, 2, 26) {real, imag} */,
  {32'h3d87a0e0, 32'h3f19f4ae} /* (11, 2, 25) {real, imag} */,
  {32'h3f1d2549, 32'hbf28191e} /* (11, 2, 24) {real, imag} */,
  {32'hbec4d794, 32'h3d5c5d61} /* (11, 2, 23) {real, imag} */,
  {32'hbe3819b6, 32'h3d57072e} /* (11, 2, 22) {real, imag} */,
  {32'h3e54685b, 32'hbf07d2e6} /* (11, 2, 21) {real, imag} */,
  {32'h3dbc91c2, 32'hbe6d56de} /* (11, 2, 20) {real, imag} */,
  {32'h3e443f56, 32'hbe249ffc} /* (11, 2, 19) {real, imag} */,
  {32'h3ddb82a4, 32'hbda4a3b0} /* (11, 2, 18) {real, imag} */,
  {32'hbdce5bdc, 32'hbc9afbc8} /* (11, 2, 17) {real, imag} */,
  {32'h3e8832fd, 32'h3e946250} /* (11, 2, 16) {real, imag} */,
  {32'hbdd2eabc, 32'hbc8399b4} /* (11, 2, 15) {real, imag} */,
  {32'hbe73e864, 32'h3ef43ab2} /* (11, 2, 14) {real, imag} */,
  {32'hbe0631ae, 32'h3eb72442} /* (11, 2, 13) {real, imag} */,
  {32'hbe261eab, 32'h3e9d2899} /* (11, 2, 12) {real, imag} */,
  {32'hbd9d7fdb, 32'h3eaa87b8} /* (11, 2, 11) {real, imag} */,
  {32'hbee9774a, 32'h3edd6098} /* (11, 2, 10) {real, imag} */,
  {32'hbe1ec5e5, 32'h3db048d6} /* (11, 2, 9) {real, imag} */,
  {32'h3f39ea27, 32'hbe3bcba8} /* (11, 2, 8) {real, imag} */,
  {32'h3e7c800a, 32'hbeadf187} /* (11, 2, 7) {real, imag} */,
  {32'h3e7d25a2, 32'h3f006988} /* (11, 2, 6) {real, imag} */,
  {32'h3f83386e, 32'h4027a44e} /* (11, 2, 5) {real, imag} */,
  {32'hc038eb7c, 32'hbfe0db92} /* (11, 2, 4) {real, imag} */,
  {32'h3f420d4e, 32'h3ea83537} /* (11, 2, 3) {real, imag} */,
  {32'h414fd23c, 32'hc094bb92} /* (11, 2, 2) {real, imag} */,
  {32'hc1b22ee0, 32'h4094410d} /* (11, 2, 1) {real, imag} */,
  {32'hc1b05fe6, 32'hc03997dd} /* (11, 2, 0) {real, imag} */,
  {32'h425828b8, 32'hc128e473} /* (11, 1, 31) {real, imag} */,
  {32'hc150f2a6, 32'h3fa397b6} /* (11, 1, 30) {real, imag} */,
  {32'hbf860f91, 32'h3eb92c88} /* (11, 1, 29) {real, imag} */,
  {32'h4012dd6a, 32'h4019fd52} /* (11, 1, 28) {real, imag} */,
  {32'hc04bfb52, 32'hbf42caa2} /* (11, 1, 27) {real, imag} */,
  {32'hbebe4c19, 32'hbe979d96} /* (11, 1, 26) {real, imag} */,
  {32'hbc9e8988, 32'hbcb8fcc0} /* (11, 1, 25) {real, imag} */,
  {32'hbf3be2a0, 32'h3eb5c5c2} /* (11, 1, 24) {real, imag} */,
  {32'hbe278aaa, 32'h3d16b98c} /* (11, 1, 23) {real, imag} */,
  {32'h3f30ff67, 32'h3edd148e} /* (11, 1, 22) {real, imag} */,
  {32'hbf24b3b3, 32'h3f03fd85} /* (11, 1, 21) {real, imag} */,
  {32'hbc74ff30, 32'hbe6bd418} /* (11, 1, 20) {real, imag} */,
  {32'hbed4bc87, 32'hbe811ae7} /* (11, 1, 19) {real, imag} */,
  {32'h3ec92734, 32'h3e2cc043} /* (11, 1, 18) {real, imag} */,
  {32'h3de2abba, 32'hbdb27d7b} /* (11, 1, 17) {real, imag} */,
  {32'h3e0d58e0, 32'h3d8b5178} /* (11, 1, 16) {real, imag} */,
  {32'h3e02144c, 32'h3ede22b7} /* (11, 1, 15) {real, imag} */,
  {32'h3de4843e, 32'hbec94fd0} /* (11, 1, 14) {real, imag} */,
  {32'h3e2ead9e, 32'hbe533833} /* (11, 1, 13) {real, imag} */,
  {32'h3e810d18, 32'hbcaadd90} /* (11, 1, 12) {real, imag} */,
  {32'hbe3e8105, 32'h3d8599f8} /* (11, 1, 11) {real, imag} */,
  {32'hbd9b7a58, 32'hbf4c444a} /* (11, 1, 10) {real, imag} */,
  {32'hbdea4a50, 32'h3ec9b67f} /* (11, 1, 9) {real, imag} */,
  {32'hbf2dc14c, 32'hbf5476fd} /* (11, 1, 8) {real, imag} */,
  {32'h3ed375ce, 32'h3ed247be} /* (11, 1, 7) {real, imag} */,
  {32'hbf9ff0dc, 32'hbf1ed53d} /* (11, 1, 6) {real, imag} */,
  {32'hc04977e0, 32'hbf5b971f} /* (11, 1, 5) {real, imag} */,
  {32'hbf090778, 32'h3f86aac5} /* (11, 1, 4) {real, imag} */,
  {32'h3f1a8a95, 32'h3eaf0cb7} /* (11, 1, 3) {real, imag} */,
  {32'hc1a3c4f9, 32'hc191f708} /* (11, 1, 2) {real, imag} */,
  {32'h4299e3e7, 32'h422fb621} /* (11, 1, 1) {real, imag} */,
  {32'h428eea0c, 32'h408f22b4} /* (11, 1, 0) {real, imag} */,
  {32'h422f8898, 32'hc20f875f} /* (11, 0, 31) {real, imag} */,
  {32'hc0d361cb, 32'h41193e16} /* (11, 0, 30) {real, imag} */,
  {32'hbfd27aea, 32'h3ee27042} /* (11, 0, 29) {real, imag} */,
  {32'hbeffd20c, 32'h3f87513c} /* (11, 0, 28) {real, imag} */,
  {32'hbfbd83d5, 32'h3fac4a98} /* (11, 0, 27) {real, imag} */,
  {32'hbe5424e8, 32'h3d943660} /* (11, 0, 26) {real, imag} */,
  {32'h3f38b7ee, 32'hbeb8fe24} /* (11, 0, 25) {real, imag} */,
  {32'h3ed02eed, 32'h3ec8aa2a} /* (11, 0, 24) {real, imag} */,
  {32'hbe9c6dd5, 32'h3f197224} /* (11, 0, 23) {real, imag} */,
  {32'h3ebf3bdc, 32'h3d52e7c4} /* (11, 0, 22) {real, imag} */,
  {32'hbe9176a8, 32'h3e90c282} /* (11, 0, 21) {real, imag} */,
  {32'hbe1e8999, 32'hbd48f784} /* (11, 0, 20) {real, imag} */,
  {32'hbe2231af, 32'hbe4c03cc} /* (11, 0, 19) {real, imag} */,
  {32'h3e8a32a0, 32'hbe02c9d3} /* (11, 0, 18) {real, imag} */,
  {32'hbd847984, 32'hbe7ab4f5} /* (11, 0, 17) {real, imag} */,
  {32'hbe8f5536, 32'h00000000} /* (11, 0, 16) {real, imag} */,
  {32'hbd847984, 32'h3e7ab4f5} /* (11, 0, 15) {real, imag} */,
  {32'h3e8a32a0, 32'h3e02c9d3} /* (11, 0, 14) {real, imag} */,
  {32'hbe2231af, 32'h3e4c03cc} /* (11, 0, 13) {real, imag} */,
  {32'hbe1e8999, 32'h3d48f784} /* (11, 0, 12) {real, imag} */,
  {32'hbe9176a8, 32'hbe90c282} /* (11, 0, 11) {real, imag} */,
  {32'h3ebf3bdc, 32'hbd52e7c4} /* (11, 0, 10) {real, imag} */,
  {32'hbe9c6dd5, 32'hbf197224} /* (11, 0, 9) {real, imag} */,
  {32'h3ed02eed, 32'hbec8aa2a} /* (11, 0, 8) {real, imag} */,
  {32'h3f38b7ee, 32'h3eb8fe24} /* (11, 0, 7) {real, imag} */,
  {32'hbe5424e8, 32'hbd943660} /* (11, 0, 6) {real, imag} */,
  {32'hbfbd83d5, 32'hbfac4a98} /* (11, 0, 5) {real, imag} */,
  {32'hbeffd20c, 32'hbf87513c} /* (11, 0, 4) {real, imag} */,
  {32'hbfd27aea, 32'hbee27042} /* (11, 0, 3) {real, imag} */,
  {32'hc0d361cb, 32'hc1193e16} /* (11, 0, 2) {real, imag} */,
  {32'h422f8898, 32'h420f875f} /* (11, 0, 1) {real, imag} */,
  {32'h4291a423, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h429efe91, 32'hc22ba8a3} /* (10, 31, 31) {real, imag} */,
  {32'hc1a6c6c3, 32'h419153f9} /* (10, 31, 30) {real, imag} */,
  {32'h3eba26f6, 32'hbf0fa254} /* (10, 31, 29) {real, imag} */,
  {32'h3f6e46f0, 32'hbf14ad6e} /* (10, 31, 28) {real, imag} */,
  {32'hc018ff05, 32'h3fae35bf} /* (10, 31, 27) {real, imag} */,
  {32'hbf72cde9, 32'h3ee495df} /* (10, 31, 26) {real, imag} */,
  {32'h3f4bec46, 32'hbdd85798} /* (10, 31, 25) {real, imag} */,
  {32'hbe4b65a5, 32'h3f9efba0} /* (10, 31, 24) {real, imag} */,
  {32'h3ed610f2, 32'hbed36679} /* (10, 31, 23) {real, imag} */,
  {32'hbf3840ff, 32'h3f264742} /* (10, 31, 22) {real, imag} */,
  {32'hbe0245ae, 32'h3f012527} /* (10, 31, 21) {real, imag} */,
  {32'hbe209591, 32'h3e33e00a} /* (10, 31, 20) {real, imag} */,
  {32'h3d8bff88, 32'hbddfbd1d} /* (10, 31, 19) {real, imag} */,
  {32'hbf000dfd, 32'h3e059b5b} /* (10, 31, 18) {real, imag} */,
  {32'h3dd1caf9, 32'hbdf32b67} /* (10, 31, 17) {real, imag} */,
  {32'h3e383cba, 32'hbe952a10} /* (10, 31, 16) {real, imag} */,
  {32'h3d11158e, 32'hbdcc2d37} /* (10, 31, 15) {real, imag} */,
  {32'hbe10a2dc, 32'hbf1a1f74} /* (10, 31, 14) {real, imag} */,
  {32'h3eadb4a1, 32'h3e440fd4} /* (10, 31, 13) {real, imag} */,
  {32'h3d80cd76, 32'hbf225556} /* (10, 31, 12) {real, imag} */,
  {32'hbf190ec6, 32'hbf0a5b84} /* (10, 31, 11) {real, imag} */,
  {32'h3efbaf31, 32'hbe619633} /* (10, 31, 10) {real, imag} */,
  {32'hbec5b17c, 32'h3e1df8ba} /* (10, 31, 9) {real, imag} */,
  {32'hbec17d14, 32'hbefe305e} /* (10, 31, 8) {real, imag} */,
  {32'h3f1a37d0, 32'h3e3df30c} /* (10, 31, 7) {real, imag} */,
  {32'hbe439d6c, 32'hbf22217c} /* (10, 31, 6) {real, imag} */,
  {32'hc02c58a1, 32'hbe316332} /* (10, 31, 5) {real, imag} */,
  {32'h40240b94, 32'hc048fb02} /* (10, 31, 4) {real, imag} */,
  {32'hbfbf9288, 32'h3ec0efc8} /* (10, 31, 3) {real, imag} */,
  {32'hc148ff00, 32'hc0035e8e} /* (10, 31, 2) {real, imag} */,
  {32'h425bfc61, 32'h414114bf} /* (10, 31, 1) {real, imag} */,
  {32'h4293f624, 32'hc09af701} /* (10, 31, 0) {real, imag} */,
  {32'hc1b96d1f, 32'hc0c32882} /* (10, 30, 31) {real, imag} */,
  {32'h41596382, 32'h407b0336} /* (10, 30, 30) {real, imag} */,
  {32'h3e98f22c, 32'hbf3bb3fa} /* (10, 30, 29) {real, imag} */,
  {32'hc05a8845, 32'h3fa34d5f} /* (10, 30, 28) {real, imag} */,
  {32'h3f38be07, 32'hc024d4b0} /* (10, 30, 27) {real, imag} */,
  {32'h3ea0cdd9, 32'h3ebc4cc4} /* (10, 30, 26) {real, imag} */,
  {32'hbe30361a, 32'hbe10cd6e} /* (10, 30, 25) {real, imag} */,
  {32'h3e9e3d37, 32'hbed981f6} /* (10, 30, 24) {real, imag} */,
  {32'h3e24d237, 32'hbe96ef5e} /* (10, 30, 23) {real, imag} */,
  {32'hbe85d3ce, 32'h3e9270b6} /* (10, 30, 22) {real, imag} */,
  {32'h3df65eba, 32'hbef4724e} /* (10, 30, 21) {real, imag} */,
  {32'h3c2f0bb0, 32'h3e3a3025} /* (10, 30, 20) {real, imag} */,
  {32'hbee26ec2, 32'h3d4fc3ce} /* (10, 30, 19) {real, imag} */,
  {32'hbe5e5ca0, 32'h3e47287e} /* (10, 30, 18) {real, imag} */,
  {32'h3e30702c, 32'h3dd96098} /* (10, 30, 17) {real, imag} */,
  {32'h3d4072d6, 32'h3c0ce4e4} /* (10, 30, 16) {real, imag} */,
  {32'hbe9f4e31, 32'h3e2609e4} /* (10, 30, 15) {real, imag} */,
  {32'h3edc69c6, 32'h3c7554c0} /* (10, 30, 14) {real, imag} */,
  {32'hbe9bee8f, 32'hbebb9980} /* (10, 30, 13) {real, imag} */,
  {32'hbd993ade, 32'hbee4c944} /* (10, 30, 12) {real, imag} */,
  {32'h3e825ba0, 32'h3f4d0b2e} /* (10, 30, 11) {real, imag} */,
  {32'hbf3e6041, 32'h3dee3dcc} /* (10, 30, 10) {real, imag} */,
  {32'hbed9558d, 32'hbefda11c} /* (10, 30, 9) {real, imag} */,
  {32'h3f7fbe08, 32'h3f3e5976} /* (10, 30, 8) {real, imag} */,
  {32'hbd4eed28, 32'hbe84b9c6} /* (10, 30, 7) {real, imag} */,
  {32'h3edb121c, 32'h3eb1844a} /* (10, 30, 6) {real, imag} */,
  {32'h3fecdb99, 32'h4003366a} /* (10, 30, 5) {real, imag} */,
  {32'hbf5745ae, 32'hc017b2b2} /* (10, 30, 4) {real, imag} */,
  {32'h3f9c33fc, 32'hbef9fe47} /* (10, 30, 3) {real, imag} */,
  {32'h419603b2, 32'h40b75182} /* (10, 30, 2) {real, imag} */,
  {32'hc225fe8d, 32'h401c5516} /* (10, 30, 1) {real, imag} */,
  {32'hc1ba787e, 32'h40483579} /* (10, 30, 0) {real, imag} */,
  {32'h4062072d, 32'hc02f14e8} /* (10, 29, 31) {real, imag} */,
  {32'hbe89bafa, 32'h403cc3f5} /* (10, 29, 30) {real, imag} */,
  {32'hbf62777a, 32'hbf3f6ded} /* (10, 29, 29) {real, imag} */,
  {32'hbf808b65, 32'hbec21998} /* (10, 29, 28) {real, imag} */,
  {32'hbee41416, 32'hbe23e9b0} /* (10, 29, 27) {real, imag} */,
  {32'hbe131ff0, 32'h3da8e1e6} /* (10, 29, 26) {real, imag} */,
  {32'hbf3941ad, 32'hbddb583a} /* (10, 29, 25) {real, imag} */,
  {32'hbe28a9cd, 32'hbecd286b} /* (10, 29, 24) {real, imag} */,
  {32'h3e30e5d8, 32'h3e271cfc} /* (10, 29, 23) {real, imag} */,
  {32'h3ec3d934, 32'hbf0a43c2} /* (10, 29, 22) {real, imag} */,
  {32'h3e46ee46, 32'hbe9d725a} /* (10, 29, 21) {real, imag} */,
  {32'h3e82f34d, 32'h3ef44d4e} /* (10, 29, 20) {real, imag} */,
  {32'hbdf93449, 32'h3e823aba} /* (10, 29, 19) {real, imag} */,
  {32'h3db7676e, 32'h3f03083f} /* (10, 29, 18) {real, imag} */,
  {32'h3ece35d1, 32'h3df7aef0} /* (10, 29, 17) {real, imag} */,
  {32'h3e80181d, 32'h3ea35781} /* (10, 29, 16) {real, imag} */,
  {32'h3e78e119, 32'h3ea7a2b7} /* (10, 29, 15) {real, imag} */,
  {32'h3bbf6c60, 32'h3e661e3c} /* (10, 29, 14) {real, imag} */,
  {32'hbdd0782a, 32'hbe0ed0de} /* (10, 29, 13) {real, imag} */,
  {32'hbe4069a9, 32'h3de3beb6} /* (10, 29, 12) {real, imag} */,
  {32'h3e05c79c, 32'hbecb789a} /* (10, 29, 11) {real, imag} */,
  {32'hbf4fb06f, 32'h3e81a298} /* (10, 29, 10) {real, imag} */,
  {32'hbea5ea66, 32'hbd78f1ec} /* (10, 29, 9) {real, imag} */,
  {32'h3ecfb88f, 32'hbc9aa348} /* (10, 29, 8) {real, imag} */,
  {32'hbda912a0, 32'hbecd37e6} /* (10, 29, 7) {real, imag} */,
  {32'h3e90f1bc, 32'hbeccc7d7} /* (10, 29, 6) {real, imag} */,
  {32'hbfa50c8d, 32'hbe98a6f2} /* (10, 29, 5) {real, imag} */,
  {32'h3fe266e6, 32'hbf71744a} /* (10, 29, 4) {real, imag} */,
  {32'hbf0d50d6, 32'h3eeaafbd} /* (10, 29, 3) {real, imag} */,
  {32'h400616b9, 32'h4086af0b} /* (10, 29, 2) {real, imag} */,
  {32'hc0932d8f, 32'hc0169b15} /* (10, 29, 1) {real, imag} */,
  {32'hbf0b8942, 32'hbed3d01e} /* (10, 29, 0) {real, imag} */,
  {32'h40a0d659, 32'hbf74a87c} /* (10, 28, 31) {real, imag} */,
  {32'hbff23e65, 32'h40067505} /* (10, 28, 30) {real, imag} */,
  {32'hbf3e0e15, 32'hbf48c00c} /* (10, 28, 29) {real, imag} */,
  {32'h3e83c62a, 32'hbfad6279} /* (10, 28, 28) {real, imag} */,
  {32'h3f3b4502, 32'h3f6a884e} /* (10, 28, 27) {real, imag} */,
  {32'hbe8e99b2, 32'hbe708c46} /* (10, 28, 26) {real, imag} */,
  {32'hbe0ea97a, 32'h3ef0f572} /* (10, 28, 25) {real, imag} */,
  {32'hbe7a4f8a, 32'h3f15bba6} /* (10, 28, 24) {real, imag} */,
  {32'h3ea8f3dc, 32'hbcc6fc50} /* (10, 28, 23) {real, imag} */,
  {32'h3e4785c2, 32'hbe36f94a} /* (10, 28, 22) {real, imag} */,
  {32'h3ead264f, 32'h3f24f36a} /* (10, 28, 21) {real, imag} */,
  {32'hbd55ee12, 32'hbe80befa} /* (10, 28, 20) {real, imag} */,
  {32'h3e998148, 32'h3e35d58a} /* (10, 28, 19) {real, imag} */,
  {32'h3ecb1034, 32'h3e51dd42} /* (10, 28, 18) {real, imag} */,
  {32'hbef15748, 32'hbdc2e7de} /* (10, 28, 17) {real, imag} */,
  {32'hbe412340, 32'hbe3e4c8e} /* (10, 28, 16) {real, imag} */,
  {32'hbce94099, 32'hbe9789d1} /* (10, 28, 15) {real, imag} */,
  {32'hbef985ac, 32'h3e54fb4d} /* (10, 28, 14) {real, imag} */,
  {32'hbda2d4be, 32'hbdfe574f} /* (10, 28, 13) {real, imag} */,
  {32'hbd26e504, 32'hbe22caea} /* (10, 28, 12) {real, imag} */,
  {32'h3d9a743e, 32'h3ec84bda} /* (10, 28, 11) {real, imag} */,
  {32'hbd7cab1e, 32'h3ecc7819} /* (10, 28, 10) {real, imag} */,
  {32'h3f818976, 32'hbdaa7794} /* (10, 28, 9) {real, imag} */,
  {32'h3e7a51c2, 32'h3f32c919} /* (10, 28, 8) {real, imag} */,
  {32'h3f0a8bbe, 32'h3ea248d0} /* (10, 28, 7) {real, imag} */,
  {32'hbf42a438, 32'hbf764a91} /* (10, 28, 6) {real, imag} */,
  {32'hbf3df03a, 32'h3db74726} /* (10, 28, 5) {real, imag} */,
  {32'h3f59b136, 32'h3d1431c0} /* (10, 28, 4) {real, imag} */,
  {32'hbea2bd6f, 32'h3e9e0276} /* (10, 28, 3) {real, imag} */,
  {32'hc0531cbd, 32'h3fde677d} /* (10, 28, 2) {real, imag} */,
  {32'h3fcfee04, 32'hc0431e08} /* (10, 28, 1) {real, imag} */,
  {32'h3f8e4851, 32'hbf48d2d6} /* (10, 28, 0) {real, imag} */,
  {32'hbf397270, 32'h4016f74f} /* (10, 27, 31) {real, imag} */,
  {32'h3e358d21, 32'hbfcf3922} /* (10, 27, 30) {real, imag} */,
  {32'hbd0781a6, 32'hbe67cf3e} /* (10, 27, 29) {real, imag} */,
  {32'hbec98c26, 32'h3dec0e60} /* (10, 27, 28) {real, imag} */,
  {32'h3eeb48f2, 32'hbdca52fc} /* (10, 27, 27) {real, imag} */,
  {32'hbec2a20a, 32'hbe36320f} /* (10, 27, 26) {real, imag} */,
  {32'h3e61c7d1, 32'h3eecdcec} /* (10, 27, 25) {real, imag} */,
  {32'h3e13ef7c, 32'hbf2614c8} /* (10, 27, 24) {real, imag} */,
  {32'h3e0065c7, 32'h3d4b01ae} /* (10, 27, 23) {real, imag} */,
  {32'hbdcc3ce4, 32'hbe7836f4} /* (10, 27, 22) {real, imag} */,
  {32'hbebe69ec, 32'h3dbb47d4} /* (10, 27, 21) {real, imag} */,
  {32'h3eb04136, 32'h3cd58a98} /* (10, 27, 20) {real, imag} */,
  {32'h3ef04e62, 32'hbdc5caa6} /* (10, 27, 19) {real, imag} */,
  {32'h3d50c5a8, 32'hbf0303a3} /* (10, 27, 18) {real, imag} */,
  {32'hbecc0665, 32'hbeb8def2} /* (10, 27, 17) {real, imag} */,
  {32'hbeb65de8, 32'h3bf428e0} /* (10, 27, 16) {real, imag} */,
  {32'h3d872c74, 32'h3ecef872} /* (10, 27, 15) {real, imag} */,
  {32'hbeb46b8a, 32'h3f08a1de} /* (10, 27, 14) {real, imag} */,
  {32'hbe251228, 32'h3e947946} /* (10, 27, 13) {real, imag} */,
  {32'h3ccb6310, 32'h3e089820} /* (10, 27, 12) {real, imag} */,
  {32'h3eb941ec, 32'h3f0fbac8} /* (10, 27, 11) {real, imag} */,
  {32'hbcf08d80, 32'h3f06e724} /* (10, 27, 10) {real, imag} */,
  {32'hbe7c6160, 32'hbf2be7ec} /* (10, 27, 9) {real, imag} */,
  {32'hbe7d51ed, 32'h3f4e30a1} /* (10, 27, 8) {real, imag} */,
  {32'hbe8b137d, 32'hbeaaa6b6} /* (10, 27, 7) {real, imag} */,
  {32'h3d16d8a6, 32'h3e2ccbba} /* (10, 27, 6) {real, imag} */,
  {32'hbca065c0, 32'hbf089e1a} /* (10, 27, 5) {real, imag} */,
  {32'hbf18c64c, 32'hbfa4a9bc} /* (10, 27, 4) {real, imag} */,
  {32'h3e632c50, 32'h3e2e0a9c} /* (10, 27, 3) {real, imag} */,
  {32'h3f262202, 32'hbd3336e4} /* (10, 27, 2) {real, imag} */,
  {32'hc06abc8a, 32'h3f8d0e4b} /* (10, 27, 1) {real, imag} */,
  {32'hbfffea3c, 32'h3f2f539a} /* (10, 27, 0) {real, imag} */,
  {32'h3e12ea6f, 32'hbde0ba35} /* (10, 26, 31) {real, imag} */,
  {32'h3e340756, 32'h3f653a70} /* (10, 26, 30) {real, imag} */,
  {32'hbf0660e2, 32'hbe99004f} /* (10, 26, 29) {real, imag} */,
  {32'hbef0f791, 32'hbe2dc047} /* (10, 26, 28) {real, imag} */,
  {32'h3ef51b72, 32'hbf10de38} /* (10, 26, 27) {real, imag} */,
  {32'h3e880f86, 32'hbe7865d0} /* (10, 26, 26) {real, imag} */,
  {32'h3e5b68c6, 32'hbc9a1a74} /* (10, 26, 25) {real, imag} */,
  {32'h3eb2085c, 32'h3ecd03a0} /* (10, 26, 24) {real, imag} */,
  {32'hbe575db9, 32'h3eada22c} /* (10, 26, 23) {real, imag} */,
  {32'hbea864fe, 32'h3f0a5a38} /* (10, 26, 22) {real, imag} */,
  {32'hbd415018, 32'h3dbb5f55} /* (10, 26, 21) {real, imag} */,
  {32'h3e3c5ec8, 32'hbd35c8d8} /* (10, 26, 20) {real, imag} */,
  {32'h3e575e53, 32'hbc185e58} /* (10, 26, 19) {real, imag} */,
  {32'h3e160ce0, 32'hbe18a832} /* (10, 26, 18) {real, imag} */,
  {32'hbe8d7742, 32'h3ea4c742} /* (10, 26, 17) {real, imag} */,
  {32'hbe4e252f, 32'hbe3410c8} /* (10, 26, 16) {real, imag} */,
  {32'hbe4f61ad, 32'hbeb07e25} /* (10, 26, 15) {real, imag} */,
  {32'h3edc0d4e, 32'hbe228c80} /* (10, 26, 14) {real, imag} */,
  {32'h3df485ac, 32'hbe8f34d3} /* (10, 26, 13) {real, imag} */,
  {32'h3e307835, 32'h3dacd542} /* (10, 26, 12) {real, imag} */,
  {32'h3f04eafa, 32'hbdc7a064} /* (10, 26, 11) {real, imag} */,
  {32'hbec9291f, 32'h3e9e04d6} /* (10, 26, 10) {real, imag} */,
  {32'h3f1723af, 32'hbf3aa62b} /* (10, 26, 9) {real, imag} */,
  {32'hbf0733ec, 32'h3d9e231a} /* (10, 26, 8) {real, imag} */,
  {32'h3de9f31a, 32'hbd3ea0aa} /* (10, 26, 7) {real, imag} */,
  {32'h3f0ce352, 32'h3dc80454} /* (10, 26, 6) {real, imag} */,
  {32'hbdf34e34, 32'h3f026ce0} /* (10, 26, 5) {real, imag} */,
  {32'h3f055990, 32'h3ef45ae2} /* (10, 26, 4) {real, imag} */,
  {32'h3eb775b0, 32'hbe630794} /* (10, 26, 3) {real, imag} */,
  {32'h3e33ca98, 32'h3f179fa5} /* (10, 26, 2) {real, imag} */,
  {32'h3e5830fb, 32'h3f6faceb} /* (10, 26, 1) {real, imag} */,
  {32'h3ef69ea5, 32'hbf890978} /* (10, 26, 0) {real, imag} */,
  {32'h3e91935c, 32'hbf849c11} /* (10, 25, 31) {real, imag} */,
  {32'hbf6f7fec, 32'hbe2fa876} /* (10, 25, 30) {real, imag} */,
  {32'h3e2d01ea, 32'hbc9be220} /* (10, 25, 29) {real, imag} */,
  {32'h3e899ee6, 32'h3d5119ac} /* (10, 25, 28) {real, imag} */,
  {32'hbebc49d7, 32'h3ef34e13} /* (10, 25, 27) {real, imag} */,
  {32'h3f2d079d, 32'h3ec7d92e} /* (10, 25, 26) {real, imag} */,
  {32'h3ca3ec04, 32'hbe4a5ba0} /* (10, 25, 25) {real, imag} */,
  {32'hbe6a2445, 32'h3df8ea24} /* (10, 25, 24) {real, imag} */,
  {32'h3e78411d, 32'hbe6b41af} /* (10, 25, 23) {real, imag} */,
  {32'hbe912bac, 32'h3f0bc44e} /* (10, 25, 22) {real, imag} */,
  {32'h3e847a21, 32'hbd88cd62} /* (10, 25, 21) {real, imag} */,
  {32'hbdcdaff6, 32'h3e7992ea} /* (10, 25, 20) {real, imag} */,
  {32'hbe11c783, 32'hbf0c4352} /* (10, 25, 19) {real, imag} */,
  {32'hbe2f21c1, 32'hbe37241a} /* (10, 25, 18) {real, imag} */,
  {32'hbde49754, 32'hbdc2f983} /* (10, 25, 17) {real, imag} */,
  {32'h3e2c5d66, 32'hbe1f3b01} /* (10, 25, 16) {real, imag} */,
  {32'hbe9373db, 32'hbca716b4} /* (10, 25, 15) {real, imag} */,
  {32'h3e0dbfbd, 32'hbd05f2dc} /* (10, 25, 14) {real, imag} */,
  {32'h3e94a0c8, 32'h3c7d6268} /* (10, 25, 13) {real, imag} */,
  {32'hbf04d64e, 32'h3e94327a} /* (10, 25, 12) {real, imag} */,
  {32'h3edbf115, 32'hbe5c1bf8} /* (10, 25, 11) {real, imag} */,
  {32'h3e3a942b, 32'h3d83dab0} /* (10, 25, 10) {real, imag} */,
  {32'hbf06f702, 32'h3ee9e925} /* (10, 25, 9) {real, imag} */,
  {32'hbf246fb4, 32'hbda1a142} /* (10, 25, 8) {real, imag} */,
  {32'h3e763c32, 32'h3e9856da} /* (10, 25, 7) {real, imag} */,
  {32'h3d1aec8c, 32'hbc5979c0} /* (10, 25, 6) {real, imag} */,
  {32'hbe8c15e7, 32'hbe31358c} /* (10, 25, 5) {real, imag} */,
  {32'h3d660260, 32'hbe7d965e} /* (10, 25, 4) {real, imag} */,
  {32'hbf436b20, 32'hbf7f86b0} /* (10, 25, 3) {real, imag} */,
  {32'hbecbf404, 32'h3f4c03fe} /* (10, 25, 2) {real, imag} */,
  {32'h3f345426, 32'hbf33471e} /* (10, 25, 1) {real, imag} */,
  {32'h3e1304cd, 32'h3e56311a} /* (10, 25, 0) {real, imag} */,
  {32'hbf2d2c34, 32'h3f20f196} /* (10, 24, 31) {real, imag} */,
  {32'h3f66be6d, 32'hbea10aa6} /* (10, 24, 30) {real, imag} */,
  {32'hbd69c1f0, 32'hbd844dea} /* (10, 24, 29) {real, imag} */,
  {32'hbf18bc52, 32'h3d4fee58} /* (10, 24, 28) {real, imag} */,
  {32'h3ed45845, 32'h3eb2d86a} /* (10, 24, 27) {real, imag} */,
  {32'h3ebd43ec, 32'hbe46fdc7} /* (10, 24, 26) {real, imag} */,
  {32'h3f52ab84, 32'hbe7806b1} /* (10, 24, 25) {real, imag} */,
  {32'h3e687609, 32'hbd9fe71c} /* (10, 24, 24) {real, imag} */,
  {32'hbeb8d2d8, 32'hbebc13a2} /* (10, 24, 23) {real, imag} */,
  {32'h3e3573bc, 32'hbe8ba8b5} /* (10, 24, 22) {real, imag} */,
  {32'h3e807f1a, 32'hbe3e2169} /* (10, 24, 21) {real, imag} */,
  {32'h3ef1e022, 32'hbc496a18} /* (10, 24, 20) {real, imag} */,
  {32'hbf088a74, 32'hbdca7901} /* (10, 24, 19) {real, imag} */,
  {32'h3e5f11f0, 32'h3e8ae8e6} /* (10, 24, 18) {real, imag} */,
  {32'hbe497abf, 32'h3cc3a9f2} /* (10, 24, 17) {real, imag} */,
  {32'h3e44da08, 32'hbd98bed6} /* (10, 24, 16) {real, imag} */,
  {32'h3b5a7270, 32'h3dc904d4} /* (10, 24, 15) {real, imag} */,
  {32'h3e5aee5c, 32'h3d0d43ac} /* (10, 24, 14) {real, imag} */,
  {32'h3e2f29d7, 32'h3e2352b2} /* (10, 24, 13) {real, imag} */,
  {32'hbe4eebb0, 32'hbefd0eab} /* (10, 24, 12) {real, imag} */,
  {32'hbf43b31c, 32'hbec361e6} /* (10, 24, 11) {real, imag} */,
  {32'h3ea944f4, 32'hbf022d24} /* (10, 24, 10) {real, imag} */,
  {32'h39c02e00, 32'h3e1fece4} /* (10, 24, 9) {real, imag} */,
  {32'h3e6bd6da, 32'hbdacd5d8} /* (10, 24, 8) {real, imag} */,
  {32'h3e66b0ee, 32'h3e1f6f35} /* (10, 24, 7) {real, imag} */,
  {32'hbe3aa38a, 32'hbbe81530} /* (10, 24, 6) {real, imag} */,
  {32'h3ea3aa99, 32'hbf2579c8} /* (10, 24, 5) {real, imag} */,
  {32'h3d94b4e0, 32'hbee822cc} /* (10, 24, 4) {real, imag} */,
  {32'hbf4fcd71, 32'h3eb1a35c} /* (10, 24, 3) {real, imag} */,
  {32'h3f518910, 32'h3e537ba4} /* (10, 24, 2) {real, imag} */,
  {32'hbfb24ca9, 32'h3e95a032} /* (10, 24, 1) {real, imag} */,
  {32'hbe707ef0, 32'h3d8f89fc} /* (10, 24, 0) {real, imag} */,
  {32'hbead7b7c, 32'hbe3de6b8} /* (10, 23, 31) {real, imag} */,
  {32'h3e9e96bb, 32'h3cc981d0} /* (10, 23, 30) {real, imag} */,
  {32'h3edda0d6, 32'hbe4f3848} /* (10, 23, 29) {real, imag} */,
  {32'hbf06fc80, 32'h3e29addd} /* (10, 23, 28) {real, imag} */,
  {32'hbf522072, 32'hbed7c20d} /* (10, 23, 27) {real, imag} */,
  {32'h3ee89094, 32'h3e5c2979} /* (10, 23, 26) {real, imag} */,
  {32'hbe922fa2, 32'hbecefc3d} /* (10, 23, 25) {real, imag} */,
  {32'hbeb5bec8, 32'hbe809cb6} /* (10, 23, 24) {real, imag} */,
  {32'hbcf29870, 32'h3e087d20} /* (10, 23, 23) {real, imag} */,
  {32'h3e573946, 32'h3eb1deb1} /* (10, 23, 22) {real, imag} */,
  {32'h3ec72496, 32'h3e2bf07f} /* (10, 23, 21) {real, imag} */,
  {32'hbec5b78c, 32'hbdde6720} /* (10, 23, 20) {real, imag} */,
  {32'h3de1e7b6, 32'h3e9fb2e6} /* (10, 23, 19) {real, imag} */,
  {32'hbdb635f4, 32'h3dbc833a} /* (10, 23, 18) {real, imag} */,
  {32'hbcaf4150, 32'hbeaf4e2e} /* (10, 23, 17) {real, imag} */,
  {32'h3e079d7f, 32'hbdfdba8f} /* (10, 23, 16) {real, imag} */,
  {32'hbea82b3c, 32'hbf023df6} /* (10, 23, 15) {real, imag} */,
  {32'h3d4cee5c, 32'h3eb12e48} /* (10, 23, 14) {real, imag} */,
  {32'h3deb7ec2, 32'h3e8cd24a} /* (10, 23, 13) {real, imag} */,
  {32'h3e49da7e, 32'h3e8c08d7} /* (10, 23, 12) {real, imag} */,
  {32'hbd853802, 32'h3ca36c64} /* (10, 23, 11) {real, imag} */,
  {32'hbf1427e9, 32'hbe82f0e6} /* (10, 23, 10) {real, imag} */,
  {32'h3d91e82e, 32'hbecf8337} /* (10, 23, 9) {real, imag} */,
  {32'hbd16f18c, 32'h3e360382} /* (10, 23, 8) {real, imag} */,
  {32'hbeadcd50, 32'hbf0190c1} /* (10, 23, 7) {real, imag} */,
  {32'hbcf179d0, 32'hbdd685ff} /* (10, 23, 6) {real, imag} */,
  {32'h3f0f3cf5, 32'h3ee7d96e} /* (10, 23, 5) {real, imag} */,
  {32'h3f14934c, 32'h3f029b66} /* (10, 23, 4) {real, imag} */,
  {32'h3dbfb233, 32'hbf0e6b00} /* (10, 23, 3) {real, imag} */,
  {32'h3d9dce12, 32'h3e1385a6} /* (10, 23, 2) {real, imag} */,
  {32'hbe65a079, 32'hbedb8d0e} /* (10, 23, 1) {real, imag} */,
  {32'h3e3517b8, 32'hbe56c3dc} /* (10, 23, 0) {real, imag} */,
  {32'h3e59c25e, 32'h3f108b20} /* (10, 22, 31) {real, imag} */,
  {32'h3eb895e7, 32'h3e193912} /* (10, 22, 30) {real, imag} */,
  {32'h3f0d75af, 32'hbe868f18} /* (10, 22, 29) {real, imag} */,
  {32'h3d9825ee, 32'hbc1b75d0} /* (10, 22, 28) {real, imag} */,
  {32'hbdab4a98, 32'hbe57adaa} /* (10, 22, 27) {real, imag} */,
  {32'h3da83776, 32'hbf767f42} /* (10, 22, 26) {real, imag} */,
  {32'hbe5804ea, 32'h3e3ea2dc} /* (10, 22, 25) {real, imag} */,
  {32'h3eae088a, 32'hbe4f30ef} /* (10, 22, 24) {real, imag} */,
  {32'hbc805a22, 32'hbed81694} /* (10, 22, 23) {real, imag} */,
  {32'hbf10f4c0, 32'hbe90c952} /* (10, 22, 22) {real, imag} */,
  {32'hbc63c410, 32'hbc00e9b0} /* (10, 22, 21) {real, imag} */,
  {32'h3d091e00, 32'h3dca9fc3} /* (10, 22, 20) {real, imag} */,
  {32'h3e1003ce, 32'hbe85c85e} /* (10, 22, 19) {real, imag} */,
  {32'hbe961929, 32'h3f287432} /* (10, 22, 18) {real, imag} */,
  {32'hbe194ae7, 32'h3d97c988} /* (10, 22, 17) {real, imag} */,
  {32'h3e968a7a, 32'hbcad6051} /* (10, 22, 16) {real, imag} */,
  {32'h3ddec206, 32'hbe5138ca} /* (10, 22, 15) {real, imag} */,
  {32'hbebbf96e, 32'hbef3cac3} /* (10, 22, 14) {real, imag} */,
  {32'hbf498cd9, 32'hbe11347f} /* (10, 22, 13) {real, imag} */,
  {32'hbe5bbeca, 32'h3ea46791} /* (10, 22, 12) {real, imag} */,
  {32'hbcedc230, 32'hbd932a68} /* (10, 22, 11) {real, imag} */,
  {32'h3f0e6c07, 32'hbe6dadd4} /* (10, 22, 10) {real, imag} */,
  {32'h3f9a1203, 32'h3f22080c} /* (10, 22, 9) {real, imag} */,
  {32'h3cd2c518, 32'hbed996de} /* (10, 22, 8) {real, imag} */,
  {32'hbf026acb, 32'h3e0b28e0} /* (10, 22, 7) {real, imag} */,
  {32'hbea3ff92, 32'hbdc8b41c} /* (10, 22, 6) {real, imag} */,
  {32'h3ea63e9d, 32'h3cfeaff0} /* (10, 22, 5) {real, imag} */,
  {32'hbed7ba32, 32'h3edcc7e4} /* (10, 22, 4) {real, imag} */,
  {32'hbf0609a1, 32'hbf0f223e} /* (10, 22, 3) {real, imag} */,
  {32'hbf02c7f1, 32'h3eab0303} /* (10, 22, 2) {real, imag} */,
  {32'h3edd45b6, 32'hbf3acea2} /* (10, 22, 1) {real, imag} */,
  {32'h3e613321, 32'h3ecb08e4} /* (10, 22, 0) {real, imag} */,
  {32'h3ddd58c0, 32'h3f619644} /* (10, 21, 31) {real, imag} */,
  {32'h3ecdcae8, 32'hbf6a414a} /* (10, 21, 30) {real, imag} */,
  {32'h3e893868, 32'h3ed120c0} /* (10, 21, 29) {real, imag} */,
  {32'hbe1f56df, 32'hbd4a6b50} /* (10, 21, 28) {real, imag} */,
  {32'hbe1ff534, 32'h3e280f58} /* (10, 21, 27) {real, imag} */,
  {32'hbec33582, 32'hbc19f688} /* (10, 21, 26) {real, imag} */,
  {32'h3eba55ca, 32'h3b246ec0} /* (10, 21, 25) {real, imag} */,
  {32'hbdcb67e1, 32'hbe0cbced} /* (10, 21, 24) {real, imag} */,
  {32'h3d6526d8, 32'hbdfe96a8} /* (10, 21, 23) {real, imag} */,
  {32'h3e22dfa0, 32'hbeeba651} /* (10, 21, 22) {real, imag} */,
  {32'h3d873354, 32'h3ed7ca2c} /* (10, 21, 21) {real, imag} */,
  {32'h3e67de01, 32'h3dc29630} /* (10, 21, 20) {real, imag} */,
  {32'h3e83ec10, 32'hbd9fe034} /* (10, 21, 19) {real, imag} */,
  {32'hbce94eb0, 32'hbe448978} /* (10, 21, 18) {real, imag} */,
  {32'hbd0cab43, 32'h3e0a2d41} /* (10, 21, 17) {real, imag} */,
  {32'h3d5e7fe8, 32'h3e2f9a24} /* (10, 21, 16) {real, imag} */,
  {32'hbd214410, 32'hbd8fefb8} /* (10, 21, 15) {real, imag} */,
  {32'h3d616fd0, 32'hbe551636} /* (10, 21, 14) {real, imag} */,
  {32'h3e8fb54c, 32'h3ead9d10} /* (10, 21, 13) {real, imag} */,
  {32'hbe4e49e6, 32'hbd290bbc} /* (10, 21, 12) {real, imag} */,
  {32'hbdbc2e66, 32'h3dc0431c} /* (10, 21, 11) {real, imag} */,
  {32'hbe353044, 32'h3e9066e5} /* (10, 21, 10) {real, imag} */,
  {32'hbdcbd6b4, 32'h3ec59990} /* (10, 21, 9) {real, imag} */,
  {32'h3ea2f08e, 32'h3e69b0ca} /* (10, 21, 8) {real, imag} */,
  {32'h3ceadecc, 32'h3d9e0f44} /* (10, 21, 7) {real, imag} */,
  {32'h3d7da398, 32'h3ec95140} /* (10, 21, 6) {real, imag} */,
  {32'hbe18f5cc, 32'hbf3b91f0} /* (10, 21, 5) {real, imag} */,
  {32'hbe6d3def, 32'hbe9922e0} /* (10, 21, 4) {real, imag} */,
  {32'h3e070ad0, 32'hbe482455} /* (10, 21, 3) {real, imag} */,
  {32'h3f086ff5, 32'h3ed0a396} /* (10, 21, 2) {real, imag} */,
  {32'hbf354e9f, 32'h3f56649e} /* (10, 21, 1) {real, imag} */,
  {32'hbe8117b3, 32'h3e9bf5fa} /* (10, 21, 0) {real, imag} */,
  {32'h3d363077, 32'h3eb17e1a} /* (10, 20, 31) {real, imag} */,
  {32'h3e1e5fac, 32'hbd273846} /* (10, 20, 30) {real, imag} */,
  {32'h3a80cbc0, 32'h3cfdb7b8} /* (10, 20, 29) {real, imag} */,
  {32'h3d626a58, 32'h3bef53c0} /* (10, 20, 28) {real, imag} */,
  {32'h3d358808, 32'hbe1997ae} /* (10, 20, 27) {real, imag} */,
  {32'hbe13d743, 32'hbe9b6d45} /* (10, 20, 26) {real, imag} */,
  {32'h3ddd3a60, 32'h3d35a350} /* (10, 20, 25) {real, imag} */,
  {32'h3ebdef97, 32'h3ea7fe78} /* (10, 20, 24) {real, imag} */,
  {32'hbe2f8391, 32'h3eae4d25} /* (10, 20, 23) {real, imag} */,
  {32'h3dbf504a, 32'hbf0adf40} /* (10, 20, 22) {real, imag} */,
  {32'h3eb733ec, 32'h3e91b54c} /* (10, 20, 21) {real, imag} */,
  {32'h3e75f3a3, 32'hbf6ced0c} /* (10, 20, 20) {real, imag} */,
  {32'h3e3a8f47, 32'hbda021fe} /* (10, 20, 19) {real, imag} */,
  {32'hbc9c8914, 32'hbbc75dc0} /* (10, 20, 18) {real, imag} */,
  {32'hbc8172fa, 32'hbe59c364} /* (10, 20, 17) {real, imag} */,
  {32'h3e354b75, 32'h3ee5d598} /* (10, 20, 16) {real, imag} */,
  {32'h3f1ab58a, 32'h3e296599} /* (10, 20, 15) {real, imag} */,
  {32'h3f2fb95c, 32'hbed92250} /* (10, 20, 14) {real, imag} */,
  {32'h3ecc2470, 32'hbc7779b0} /* (10, 20, 13) {real, imag} */,
  {32'h3ed2590b, 32'h3edba271} /* (10, 20, 12) {real, imag} */,
  {32'hbe325d14, 32'hbf16fb79} /* (10, 20, 11) {real, imag} */,
  {32'hbe075636, 32'hbf195dfc} /* (10, 20, 10) {real, imag} */,
  {32'hbee76069, 32'hbe2f3fc4} /* (10, 20, 9) {real, imag} */,
  {32'hbf32548e, 32'h3f10ad5c} /* (10, 20, 8) {real, imag} */,
  {32'h3acf3c00, 32'h3e8f4533} /* (10, 20, 7) {real, imag} */,
  {32'h3c90fbce, 32'hbd8159b1} /* (10, 20, 6) {real, imag} */,
  {32'hbef98fe0, 32'hbd295612} /* (10, 20, 5) {real, imag} */,
  {32'h3f18d651, 32'hbee0cd8e} /* (10, 20, 4) {real, imag} */,
  {32'hbddaf31c, 32'hbe6fe81a} /* (10, 20, 3) {real, imag} */,
  {32'hbd2ea8d4, 32'h3e2095f6} /* (10, 20, 2) {real, imag} */,
  {32'h3d8bf65c, 32'h3df497fc} /* (10, 20, 1) {real, imag} */,
  {32'h3ee8350e, 32'h3d8c8508} /* (10, 20, 0) {real, imag} */,
  {32'h3e323490, 32'hbee63914} /* (10, 19, 31) {real, imag} */,
  {32'hbc0a9490, 32'hbde5422e} /* (10, 19, 30) {real, imag} */,
  {32'hbead8fbf, 32'h3e72091a} /* (10, 19, 29) {real, imag} */,
  {32'hbeae5727, 32'hbd99a04c} /* (10, 19, 28) {real, imag} */,
  {32'h3e499f61, 32'hbd1af158} /* (10, 19, 27) {real, imag} */,
  {32'h3f1c23d8, 32'h3e4505f7} /* (10, 19, 26) {real, imag} */,
  {32'hbf2c7dc0, 32'hbcf3c0ca} /* (10, 19, 25) {real, imag} */,
  {32'hbdb40354, 32'h3e8d177e} /* (10, 19, 24) {real, imag} */,
  {32'hbf3660cc, 32'h3c9663b0} /* (10, 19, 23) {real, imag} */,
  {32'h3e5f9149, 32'hbe98da90} /* (10, 19, 22) {real, imag} */,
  {32'hbe7896e7, 32'h3d789f4c} /* (10, 19, 21) {real, imag} */,
  {32'hbe96b404, 32'hbf420a74} /* (10, 19, 20) {real, imag} */,
  {32'h3ed4107a, 32'hbead62a8} /* (10, 19, 19) {real, imag} */,
  {32'h3ee80b84, 32'hbd3aedd6} /* (10, 19, 18) {real, imag} */,
  {32'hbe0c162a, 32'hbdfa210e} /* (10, 19, 17) {real, imag} */,
  {32'h3e2f03d6, 32'h3dfc8cda} /* (10, 19, 16) {real, imag} */,
  {32'h3ddedb84, 32'h3f0ae738} /* (10, 19, 15) {real, imag} */,
  {32'hbe4c3f0a, 32'h3dd69af3} /* (10, 19, 14) {real, imag} */,
  {32'h3c4af8c0, 32'hbefc77d8} /* (10, 19, 13) {real, imag} */,
  {32'hbf169dd6, 32'h3e15e2fa} /* (10, 19, 12) {real, imag} */,
  {32'h3e9cd426, 32'h3e993716} /* (10, 19, 11) {real, imag} */,
  {32'hbe622446, 32'hbec8f396} /* (10, 19, 10) {real, imag} */,
  {32'hbd9cc818, 32'hbe54d5bc} /* (10, 19, 9) {real, imag} */,
  {32'h3f0111f8, 32'h3e8cf746} /* (10, 19, 8) {real, imag} */,
  {32'h3e9dead6, 32'hbd890416} /* (10, 19, 7) {real, imag} */,
  {32'hbe932130, 32'h3ea19e85} /* (10, 19, 6) {real, imag} */,
  {32'hbc994300, 32'h3c5e28a0} /* (10, 19, 5) {real, imag} */,
  {32'hbf2b81e9, 32'hbe2e1866} /* (10, 19, 4) {real, imag} */,
  {32'hbdbae008, 32'h3ec7b4ee} /* (10, 19, 3) {real, imag} */,
  {32'h3ea28d1b, 32'hbd94a478} /* (10, 19, 2) {real, imag} */,
  {32'h3e0747f5, 32'h3def4240} /* (10, 19, 1) {real, imag} */,
  {32'hbe87d3e4, 32'h3e061249} /* (10, 19, 0) {real, imag} */,
  {32'hbe4b93d4, 32'h3eb84052} /* (10, 18, 31) {real, imag} */,
  {32'hbee0aa65, 32'hbe92c846} /* (10, 18, 30) {real, imag} */,
  {32'h3defd0c1, 32'hbe73f306} /* (10, 18, 29) {real, imag} */,
  {32'hbe64ea3c, 32'h3dfb6aad} /* (10, 18, 28) {real, imag} */,
  {32'hbecc9a3d, 32'hbde27354} /* (10, 18, 27) {real, imag} */,
  {32'hbe8fb9c9, 32'hbee9e6c8} /* (10, 18, 26) {real, imag} */,
  {32'h3d0c5564, 32'hbe67fa78} /* (10, 18, 25) {real, imag} */,
  {32'h3d2314e8, 32'hbc2b1246} /* (10, 18, 24) {real, imag} */,
  {32'h3e1cb73e, 32'h3e670cf2} /* (10, 18, 23) {real, imag} */,
  {32'hbd5cc1ac, 32'hbe4935a2} /* (10, 18, 22) {real, imag} */,
  {32'hbe8282fd, 32'hbeb35619} /* (10, 18, 21) {real, imag} */,
  {32'hbe002586, 32'h3e1a33f8} /* (10, 18, 20) {real, imag} */,
  {32'hbd2475ec, 32'h3e619900} /* (10, 18, 19) {real, imag} */,
  {32'hbf269095, 32'hbe8886d4} /* (10, 18, 18) {real, imag} */,
  {32'hbe489a27, 32'h3e910f98} /* (10, 18, 17) {real, imag} */,
  {32'hbea29c90, 32'h3d4bee20} /* (10, 18, 16) {real, imag} */,
  {32'hbe1ebb90, 32'hbdfca7f7} /* (10, 18, 15) {real, imag} */,
  {32'hbef5dc4c, 32'hbd045bb6} /* (10, 18, 14) {real, imag} */,
  {32'hbe3f9eac, 32'hbe12f9cf} /* (10, 18, 13) {real, imag} */,
  {32'h3ec31bd0, 32'hbd2973f8} /* (10, 18, 12) {real, imag} */,
  {32'hbebc7bc3, 32'hb9e2e580} /* (10, 18, 11) {real, imag} */,
  {32'h3efa794a, 32'hbe61b230} /* (10, 18, 10) {real, imag} */,
  {32'hbeadd784, 32'h3c9d87c8} /* (10, 18, 9) {real, imag} */,
  {32'h3e0b06ce, 32'hbcd12674} /* (10, 18, 8) {real, imag} */,
  {32'h3e68882c, 32'hbc14e880} /* (10, 18, 7) {real, imag} */,
  {32'h3d503c48, 32'hbd8e8f8a} /* (10, 18, 6) {real, imag} */,
  {32'h3e0da36a, 32'hbea789a6} /* (10, 18, 5) {real, imag} */,
  {32'hbc8fafa4, 32'h3f18f33e} /* (10, 18, 4) {real, imag} */,
  {32'hbd7283b4, 32'hbec05b34} /* (10, 18, 3) {real, imag} */,
  {32'h3ea1f970, 32'hbd835f1a} /* (10, 18, 2) {real, imag} */,
  {32'hbdfc3d54, 32'h3defd73c} /* (10, 18, 1) {real, imag} */,
  {32'h3e3817ae, 32'hbabf4500} /* (10, 18, 0) {real, imag} */,
  {32'h3c3a0ab0, 32'h3d992a1e} /* (10, 17, 31) {real, imag} */,
  {32'h3eb0822e, 32'h3d38a801} /* (10, 17, 30) {real, imag} */,
  {32'h3e197e5f, 32'h3d0d814c} /* (10, 17, 29) {real, imag} */,
  {32'hbe08bbd0, 32'h3c0cf420} /* (10, 17, 28) {real, imag} */,
  {32'hbd4ea818, 32'hbe87a424} /* (10, 17, 27) {real, imag} */,
  {32'hbdd1947f, 32'hbec285c1} /* (10, 17, 26) {real, imag} */,
  {32'hbd899612, 32'hbe1bfdbb} /* (10, 17, 25) {real, imag} */,
  {32'h3dd9ede6, 32'hbddee504} /* (10, 17, 24) {real, imag} */,
  {32'h3e7444c5, 32'h3d26f574} /* (10, 17, 23) {real, imag} */,
  {32'hbe0165e2, 32'hbea44cc3} /* (10, 17, 22) {real, imag} */,
  {32'h3e90b14c, 32'hbd500dc0} /* (10, 17, 21) {real, imag} */,
  {32'hbcbee0c0, 32'h3d6653cb} /* (10, 17, 20) {real, imag} */,
  {32'h3e8e1378, 32'h3ee1c03a} /* (10, 17, 19) {real, imag} */,
  {32'h3e122540, 32'h3e22ac6c} /* (10, 17, 18) {real, imag} */,
  {32'hbd481c40, 32'h3ea3ba62} /* (10, 17, 17) {real, imag} */,
  {32'hbd4a1a4d, 32'h3dd98e40} /* (10, 17, 16) {real, imag} */,
  {32'h3d8b0468, 32'hbd0166ac} /* (10, 17, 15) {real, imag} */,
  {32'h3cbda87d, 32'hbdbea20c} /* (10, 17, 14) {real, imag} */,
  {32'h3e61be9c, 32'hbeb14358} /* (10, 17, 13) {real, imag} */,
  {32'hbd71bebc, 32'hbdc7a6fa} /* (10, 17, 12) {real, imag} */,
  {32'hbe617af8, 32'hbec422e6} /* (10, 17, 11) {real, imag} */,
  {32'hbedbcf1f, 32'hbd55be90} /* (10, 17, 10) {real, imag} */,
  {32'h3d83ee6a, 32'h3e65a8fc} /* (10, 17, 9) {real, imag} */,
  {32'hbe3f516a, 32'h3d1370ef} /* (10, 17, 8) {real, imag} */,
  {32'h3ea8045a, 32'hbe0c9e97} /* (10, 17, 7) {real, imag} */,
  {32'h3d53490d, 32'hbeba02aa} /* (10, 17, 6) {real, imag} */,
  {32'hbcf5c7f8, 32'h3d92d3fa} /* (10, 17, 5) {real, imag} */,
  {32'h3e0e4152, 32'hbe1a45a4} /* (10, 17, 4) {real, imag} */,
  {32'hbda8f10e, 32'h3ea34b36} /* (10, 17, 3) {real, imag} */,
  {32'h3c88b810, 32'h3ebd5f0c} /* (10, 17, 2) {real, imag} */,
  {32'hbe91233c, 32'hbeaee632} /* (10, 17, 1) {real, imag} */,
  {32'hbd64cf9e, 32'h3d057ca2} /* (10, 17, 0) {real, imag} */,
  {32'h3e20a4de, 32'h3e13ad0a} /* (10, 16, 31) {real, imag} */,
  {32'h3e952492, 32'h3cc8019c} /* (10, 16, 30) {real, imag} */,
  {32'hbe1cb169, 32'h3dfba4c1} /* (10, 16, 29) {real, imag} */,
  {32'hbb0e80e0, 32'h3e8b8c0c} /* (10, 16, 28) {real, imag} */,
  {32'h3d7e8f82, 32'h3dc78213} /* (10, 16, 27) {real, imag} */,
  {32'h3e27d178, 32'h3da0b31e} /* (10, 16, 26) {real, imag} */,
  {32'hbe3f5ce9, 32'h3e0a15d2} /* (10, 16, 25) {real, imag} */,
  {32'hbec58213, 32'hbd54d3cc} /* (10, 16, 24) {real, imag} */,
  {32'hbe106e0e, 32'hbe2bffa1} /* (10, 16, 23) {real, imag} */,
  {32'h3e4b6be0, 32'h3ab41c00} /* (10, 16, 22) {real, imag} */,
  {32'hbe5d8390, 32'hbee03c63} /* (10, 16, 21) {real, imag} */,
  {32'hbcfd9048, 32'hbde69390} /* (10, 16, 20) {real, imag} */,
  {32'h3df1d3a7, 32'hbe92e71c} /* (10, 16, 19) {real, imag} */,
  {32'h3e0165b9, 32'hbecfa58c} /* (10, 16, 18) {real, imag} */,
  {32'h3eb5cee0, 32'hbd473f12} /* (10, 16, 17) {real, imag} */,
  {32'hbe729103, 32'h00000000} /* (10, 16, 16) {real, imag} */,
  {32'h3eb5cee0, 32'h3d473f12} /* (10, 16, 15) {real, imag} */,
  {32'h3e0165b9, 32'h3ecfa58c} /* (10, 16, 14) {real, imag} */,
  {32'h3df1d3a7, 32'h3e92e71c} /* (10, 16, 13) {real, imag} */,
  {32'hbcfd9048, 32'h3de69390} /* (10, 16, 12) {real, imag} */,
  {32'hbe5d8390, 32'h3ee03c63} /* (10, 16, 11) {real, imag} */,
  {32'h3e4b6be0, 32'hbab41c00} /* (10, 16, 10) {real, imag} */,
  {32'hbe106e0e, 32'h3e2bffa1} /* (10, 16, 9) {real, imag} */,
  {32'hbec58213, 32'h3d54d3cc} /* (10, 16, 8) {real, imag} */,
  {32'hbe3f5ce9, 32'hbe0a15d2} /* (10, 16, 7) {real, imag} */,
  {32'h3e27d178, 32'hbda0b31e} /* (10, 16, 6) {real, imag} */,
  {32'h3d7e8f82, 32'hbdc78213} /* (10, 16, 5) {real, imag} */,
  {32'hbb0e80e0, 32'hbe8b8c0c} /* (10, 16, 4) {real, imag} */,
  {32'hbe1cb169, 32'hbdfba4c1} /* (10, 16, 3) {real, imag} */,
  {32'h3e952492, 32'hbcc8019c} /* (10, 16, 2) {real, imag} */,
  {32'h3e20a4de, 32'hbe13ad0a} /* (10, 16, 1) {real, imag} */,
  {32'hbd861760, 32'h00000000} /* (10, 16, 0) {real, imag} */,
  {32'hbe91233c, 32'h3eaee632} /* (10, 15, 31) {real, imag} */,
  {32'h3c88b810, 32'hbebd5f0c} /* (10, 15, 30) {real, imag} */,
  {32'hbda8f10e, 32'hbea34b36} /* (10, 15, 29) {real, imag} */,
  {32'h3e0e4152, 32'h3e1a45a4} /* (10, 15, 28) {real, imag} */,
  {32'hbcf5c7f8, 32'hbd92d3fa} /* (10, 15, 27) {real, imag} */,
  {32'h3d53490d, 32'h3eba02aa} /* (10, 15, 26) {real, imag} */,
  {32'h3ea8045a, 32'h3e0c9e97} /* (10, 15, 25) {real, imag} */,
  {32'hbe3f516a, 32'hbd1370ef} /* (10, 15, 24) {real, imag} */,
  {32'h3d83ee6a, 32'hbe65a8fc} /* (10, 15, 23) {real, imag} */,
  {32'hbedbcf1f, 32'h3d55be90} /* (10, 15, 22) {real, imag} */,
  {32'hbe617af8, 32'h3ec422e6} /* (10, 15, 21) {real, imag} */,
  {32'hbd71bebc, 32'h3dc7a6fa} /* (10, 15, 20) {real, imag} */,
  {32'h3e61be9c, 32'h3eb14358} /* (10, 15, 19) {real, imag} */,
  {32'h3cbda87d, 32'h3dbea20c} /* (10, 15, 18) {real, imag} */,
  {32'h3d8b0468, 32'h3d0166ac} /* (10, 15, 17) {real, imag} */,
  {32'hbd4a1a4d, 32'hbdd98e40} /* (10, 15, 16) {real, imag} */,
  {32'hbd481c40, 32'hbea3ba62} /* (10, 15, 15) {real, imag} */,
  {32'h3e122540, 32'hbe22ac6c} /* (10, 15, 14) {real, imag} */,
  {32'h3e8e1378, 32'hbee1c03a} /* (10, 15, 13) {real, imag} */,
  {32'hbcbee0c0, 32'hbd6653cb} /* (10, 15, 12) {real, imag} */,
  {32'h3e90b14c, 32'h3d500dc0} /* (10, 15, 11) {real, imag} */,
  {32'hbe0165e2, 32'h3ea44cc3} /* (10, 15, 10) {real, imag} */,
  {32'h3e7444c5, 32'hbd26f574} /* (10, 15, 9) {real, imag} */,
  {32'h3dd9ede6, 32'h3ddee504} /* (10, 15, 8) {real, imag} */,
  {32'hbd899612, 32'h3e1bfdbb} /* (10, 15, 7) {real, imag} */,
  {32'hbdd1947f, 32'h3ec285c1} /* (10, 15, 6) {real, imag} */,
  {32'hbd4ea818, 32'h3e87a424} /* (10, 15, 5) {real, imag} */,
  {32'hbe08bbd0, 32'hbc0cf420} /* (10, 15, 4) {real, imag} */,
  {32'h3e197e5f, 32'hbd0d814c} /* (10, 15, 3) {real, imag} */,
  {32'h3eb0822e, 32'hbd38a801} /* (10, 15, 2) {real, imag} */,
  {32'h3c3a0ab0, 32'hbd992a1e} /* (10, 15, 1) {real, imag} */,
  {32'hbd64cf9e, 32'hbd057ca2} /* (10, 15, 0) {real, imag} */,
  {32'hbdfc3d54, 32'hbdefd73c} /* (10, 14, 31) {real, imag} */,
  {32'h3ea1f970, 32'h3d835f1a} /* (10, 14, 30) {real, imag} */,
  {32'hbd7283b4, 32'h3ec05b34} /* (10, 14, 29) {real, imag} */,
  {32'hbc8fafa4, 32'hbf18f33e} /* (10, 14, 28) {real, imag} */,
  {32'h3e0da36a, 32'h3ea789a6} /* (10, 14, 27) {real, imag} */,
  {32'h3d503c48, 32'h3d8e8f8a} /* (10, 14, 26) {real, imag} */,
  {32'h3e68882c, 32'h3c14e880} /* (10, 14, 25) {real, imag} */,
  {32'h3e0b06ce, 32'h3cd12674} /* (10, 14, 24) {real, imag} */,
  {32'hbeadd784, 32'hbc9d87c8} /* (10, 14, 23) {real, imag} */,
  {32'h3efa794a, 32'h3e61b230} /* (10, 14, 22) {real, imag} */,
  {32'hbebc7bc3, 32'h39e2e580} /* (10, 14, 21) {real, imag} */,
  {32'h3ec31bd0, 32'h3d2973f8} /* (10, 14, 20) {real, imag} */,
  {32'hbe3f9eac, 32'h3e12f9cf} /* (10, 14, 19) {real, imag} */,
  {32'hbef5dc4c, 32'h3d045bb6} /* (10, 14, 18) {real, imag} */,
  {32'hbe1ebb90, 32'h3dfca7f7} /* (10, 14, 17) {real, imag} */,
  {32'hbea29c90, 32'hbd4bee20} /* (10, 14, 16) {real, imag} */,
  {32'hbe489a27, 32'hbe910f98} /* (10, 14, 15) {real, imag} */,
  {32'hbf269095, 32'h3e8886d4} /* (10, 14, 14) {real, imag} */,
  {32'hbd2475ec, 32'hbe619900} /* (10, 14, 13) {real, imag} */,
  {32'hbe002586, 32'hbe1a33f8} /* (10, 14, 12) {real, imag} */,
  {32'hbe8282fd, 32'h3eb35619} /* (10, 14, 11) {real, imag} */,
  {32'hbd5cc1ac, 32'h3e4935a2} /* (10, 14, 10) {real, imag} */,
  {32'h3e1cb73e, 32'hbe670cf2} /* (10, 14, 9) {real, imag} */,
  {32'h3d2314e8, 32'h3c2b1246} /* (10, 14, 8) {real, imag} */,
  {32'h3d0c5564, 32'h3e67fa78} /* (10, 14, 7) {real, imag} */,
  {32'hbe8fb9c9, 32'h3ee9e6c8} /* (10, 14, 6) {real, imag} */,
  {32'hbecc9a3d, 32'h3de27354} /* (10, 14, 5) {real, imag} */,
  {32'hbe64ea3c, 32'hbdfb6aad} /* (10, 14, 4) {real, imag} */,
  {32'h3defd0c1, 32'h3e73f306} /* (10, 14, 3) {real, imag} */,
  {32'hbee0aa65, 32'h3e92c846} /* (10, 14, 2) {real, imag} */,
  {32'hbe4b93d4, 32'hbeb84052} /* (10, 14, 1) {real, imag} */,
  {32'h3e3817ae, 32'h3abf4500} /* (10, 14, 0) {real, imag} */,
  {32'h3e0747f5, 32'hbdef4240} /* (10, 13, 31) {real, imag} */,
  {32'h3ea28d1b, 32'h3d94a478} /* (10, 13, 30) {real, imag} */,
  {32'hbdbae008, 32'hbec7b4ee} /* (10, 13, 29) {real, imag} */,
  {32'hbf2b81e9, 32'h3e2e1866} /* (10, 13, 28) {real, imag} */,
  {32'hbc994300, 32'hbc5e28a0} /* (10, 13, 27) {real, imag} */,
  {32'hbe932130, 32'hbea19e85} /* (10, 13, 26) {real, imag} */,
  {32'h3e9dead6, 32'h3d890416} /* (10, 13, 25) {real, imag} */,
  {32'h3f0111f8, 32'hbe8cf746} /* (10, 13, 24) {real, imag} */,
  {32'hbd9cc818, 32'h3e54d5bc} /* (10, 13, 23) {real, imag} */,
  {32'hbe622446, 32'h3ec8f396} /* (10, 13, 22) {real, imag} */,
  {32'h3e9cd426, 32'hbe993716} /* (10, 13, 21) {real, imag} */,
  {32'hbf169dd6, 32'hbe15e2fa} /* (10, 13, 20) {real, imag} */,
  {32'h3c4af8c0, 32'h3efc77d8} /* (10, 13, 19) {real, imag} */,
  {32'hbe4c3f0a, 32'hbdd69af3} /* (10, 13, 18) {real, imag} */,
  {32'h3ddedb84, 32'hbf0ae738} /* (10, 13, 17) {real, imag} */,
  {32'h3e2f03d6, 32'hbdfc8cda} /* (10, 13, 16) {real, imag} */,
  {32'hbe0c162a, 32'h3dfa210e} /* (10, 13, 15) {real, imag} */,
  {32'h3ee80b84, 32'h3d3aedd6} /* (10, 13, 14) {real, imag} */,
  {32'h3ed4107a, 32'h3ead62a8} /* (10, 13, 13) {real, imag} */,
  {32'hbe96b404, 32'h3f420a74} /* (10, 13, 12) {real, imag} */,
  {32'hbe7896e7, 32'hbd789f4c} /* (10, 13, 11) {real, imag} */,
  {32'h3e5f9149, 32'h3e98da90} /* (10, 13, 10) {real, imag} */,
  {32'hbf3660cc, 32'hbc9663b0} /* (10, 13, 9) {real, imag} */,
  {32'hbdb40354, 32'hbe8d177e} /* (10, 13, 8) {real, imag} */,
  {32'hbf2c7dc0, 32'h3cf3c0ca} /* (10, 13, 7) {real, imag} */,
  {32'h3f1c23d8, 32'hbe4505f7} /* (10, 13, 6) {real, imag} */,
  {32'h3e499f61, 32'h3d1af158} /* (10, 13, 5) {real, imag} */,
  {32'hbeae5727, 32'h3d99a04c} /* (10, 13, 4) {real, imag} */,
  {32'hbead8fbf, 32'hbe72091a} /* (10, 13, 3) {real, imag} */,
  {32'hbc0a9490, 32'h3de5422e} /* (10, 13, 2) {real, imag} */,
  {32'h3e323490, 32'h3ee63914} /* (10, 13, 1) {real, imag} */,
  {32'hbe87d3e4, 32'hbe061249} /* (10, 13, 0) {real, imag} */,
  {32'h3d8bf65c, 32'hbdf497fc} /* (10, 12, 31) {real, imag} */,
  {32'hbd2ea8d4, 32'hbe2095f6} /* (10, 12, 30) {real, imag} */,
  {32'hbddaf31c, 32'h3e6fe81a} /* (10, 12, 29) {real, imag} */,
  {32'h3f18d651, 32'h3ee0cd8e} /* (10, 12, 28) {real, imag} */,
  {32'hbef98fe0, 32'h3d295612} /* (10, 12, 27) {real, imag} */,
  {32'h3c90fbce, 32'h3d8159b1} /* (10, 12, 26) {real, imag} */,
  {32'h3acf3c00, 32'hbe8f4533} /* (10, 12, 25) {real, imag} */,
  {32'hbf32548e, 32'hbf10ad5c} /* (10, 12, 24) {real, imag} */,
  {32'hbee76069, 32'h3e2f3fc4} /* (10, 12, 23) {real, imag} */,
  {32'hbe075636, 32'h3f195dfc} /* (10, 12, 22) {real, imag} */,
  {32'hbe325d14, 32'h3f16fb79} /* (10, 12, 21) {real, imag} */,
  {32'h3ed2590b, 32'hbedba271} /* (10, 12, 20) {real, imag} */,
  {32'h3ecc2470, 32'h3c7779b0} /* (10, 12, 19) {real, imag} */,
  {32'h3f2fb95c, 32'h3ed92250} /* (10, 12, 18) {real, imag} */,
  {32'h3f1ab58a, 32'hbe296599} /* (10, 12, 17) {real, imag} */,
  {32'h3e354b75, 32'hbee5d598} /* (10, 12, 16) {real, imag} */,
  {32'hbc8172fa, 32'h3e59c364} /* (10, 12, 15) {real, imag} */,
  {32'hbc9c8914, 32'h3bc75dc0} /* (10, 12, 14) {real, imag} */,
  {32'h3e3a8f47, 32'h3da021fe} /* (10, 12, 13) {real, imag} */,
  {32'h3e75f3a3, 32'h3f6ced0c} /* (10, 12, 12) {real, imag} */,
  {32'h3eb733ec, 32'hbe91b54c} /* (10, 12, 11) {real, imag} */,
  {32'h3dbf504a, 32'h3f0adf40} /* (10, 12, 10) {real, imag} */,
  {32'hbe2f8391, 32'hbeae4d25} /* (10, 12, 9) {real, imag} */,
  {32'h3ebdef97, 32'hbea7fe78} /* (10, 12, 8) {real, imag} */,
  {32'h3ddd3a60, 32'hbd35a350} /* (10, 12, 7) {real, imag} */,
  {32'hbe13d743, 32'h3e9b6d45} /* (10, 12, 6) {real, imag} */,
  {32'h3d358808, 32'h3e1997ae} /* (10, 12, 5) {real, imag} */,
  {32'h3d626a58, 32'hbbef53c0} /* (10, 12, 4) {real, imag} */,
  {32'h3a80cbc0, 32'hbcfdb7b8} /* (10, 12, 3) {real, imag} */,
  {32'h3e1e5fac, 32'h3d273846} /* (10, 12, 2) {real, imag} */,
  {32'h3d363077, 32'hbeb17e1a} /* (10, 12, 1) {real, imag} */,
  {32'h3ee8350e, 32'hbd8c8508} /* (10, 12, 0) {real, imag} */,
  {32'hbf354e9f, 32'hbf56649e} /* (10, 11, 31) {real, imag} */,
  {32'h3f086ff5, 32'hbed0a396} /* (10, 11, 30) {real, imag} */,
  {32'h3e070ad0, 32'h3e482455} /* (10, 11, 29) {real, imag} */,
  {32'hbe6d3def, 32'h3e9922e0} /* (10, 11, 28) {real, imag} */,
  {32'hbe18f5cc, 32'h3f3b91f0} /* (10, 11, 27) {real, imag} */,
  {32'h3d7da398, 32'hbec95140} /* (10, 11, 26) {real, imag} */,
  {32'h3ceadecc, 32'hbd9e0f44} /* (10, 11, 25) {real, imag} */,
  {32'h3ea2f08e, 32'hbe69b0ca} /* (10, 11, 24) {real, imag} */,
  {32'hbdcbd6b4, 32'hbec59990} /* (10, 11, 23) {real, imag} */,
  {32'hbe353044, 32'hbe9066e5} /* (10, 11, 22) {real, imag} */,
  {32'hbdbc2e66, 32'hbdc0431c} /* (10, 11, 21) {real, imag} */,
  {32'hbe4e49e6, 32'h3d290bbc} /* (10, 11, 20) {real, imag} */,
  {32'h3e8fb54c, 32'hbead9d10} /* (10, 11, 19) {real, imag} */,
  {32'h3d616fd0, 32'h3e551636} /* (10, 11, 18) {real, imag} */,
  {32'hbd214410, 32'h3d8fefb8} /* (10, 11, 17) {real, imag} */,
  {32'h3d5e7fe8, 32'hbe2f9a24} /* (10, 11, 16) {real, imag} */,
  {32'hbd0cab43, 32'hbe0a2d41} /* (10, 11, 15) {real, imag} */,
  {32'hbce94eb0, 32'h3e448978} /* (10, 11, 14) {real, imag} */,
  {32'h3e83ec10, 32'h3d9fe034} /* (10, 11, 13) {real, imag} */,
  {32'h3e67de01, 32'hbdc29630} /* (10, 11, 12) {real, imag} */,
  {32'h3d873354, 32'hbed7ca2c} /* (10, 11, 11) {real, imag} */,
  {32'h3e22dfa0, 32'h3eeba651} /* (10, 11, 10) {real, imag} */,
  {32'h3d6526d8, 32'h3dfe96a8} /* (10, 11, 9) {real, imag} */,
  {32'hbdcb67e1, 32'h3e0cbced} /* (10, 11, 8) {real, imag} */,
  {32'h3eba55ca, 32'hbb246ec0} /* (10, 11, 7) {real, imag} */,
  {32'hbec33582, 32'h3c19f688} /* (10, 11, 6) {real, imag} */,
  {32'hbe1ff534, 32'hbe280f58} /* (10, 11, 5) {real, imag} */,
  {32'hbe1f56df, 32'h3d4a6b50} /* (10, 11, 4) {real, imag} */,
  {32'h3e893868, 32'hbed120c0} /* (10, 11, 3) {real, imag} */,
  {32'h3ecdcae8, 32'h3f6a414a} /* (10, 11, 2) {real, imag} */,
  {32'h3ddd58c0, 32'hbf619644} /* (10, 11, 1) {real, imag} */,
  {32'hbe8117b3, 32'hbe9bf5fa} /* (10, 11, 0) {real, imag} */,
  {32'h3edd45b6, 32'h3f3acea2} /* (10, 10, 31) {real, imag} */,
  {32'hbf02c7f1, 32'hbeab0303} /* (10, 10, 30) {real, imag} */,
  {32'hbf0609a1, 32'h3f0f223e} /* (10, 10, 29) {real, imag} */,
  {32'hbed7ba32, 32'hbedcc7e4} /* (10, 10, 28) {real, imag} */,
  {32'h3ea63e9d, 32'hbcfeaff0} /* (10, 10, 27) {real, imag} */,
  {32'hbea3ff92, 32'h3dc8b41c} /* (10, 10, 26) {real, imag} */,
  {32'hbf026acb, 32'hbe0b28e0} /* (10, 10, 25) {real, imag} */,
  {32'h3cd2c518, 32'h3ed996de} /* (10, 10, 24) {real, imag} */,
  {32'h3f9a1203, 32'hbf22080c} /* (10, 10, 23) {real, imag} */,
  {32'h3f0e6c07, 32'h3e6dadd4} /* (10, 10, 22) {real, imag} */,
  {32'hbcedc230, 32'h3d932a68} /* (10, 10, 21) {real, imag} */,
  {32'hbe5bbeca, 32'hbea46791} /* (10, 10, 20) {real, imag} */,
  {32'hbf498cd9, 32'h3e11347f} /* (10, 10, 19) {real, imag} */,
  {32'hbebbf96e, 32'h3ef3cac3} /* (10, 10, 18) {real, imag} */,
  {32'h3ddec206, 32'h3e5138ca} /* (10, 10, 17) {real, imag} */,
  {32'h3e968a7a, 32'h3cad6051} /* (10, 10, 16) {real, imag} */,
  {32'hbe194ae7, 32'hbd97c988} /* (10, 10, 15) {real, imag} */,
  {32'hbe961929, 32'hbf287432} /* (10, 10, 14) {real, imag} */,
  {32'h3e1003ce, 32'h3e85c85e} /* (10, 10, 13) {real, imag} */,
  {32'h3d091e00, 32'hbdca9fc3} /* (10, 10, 12) {real, imag} */,
  {32'hbc63c410, 32'h3c00e9b0} /* (10, 10, 11) {real, imag} */,
  {32'hbf10f4c0, 32'h3e90c952} /* (10, 10, 10) {real, imag} */,
  {32'hbc805a22, 32'h3ed81694} /* (10, 10, 9) {real, imag} */,
  {32'h3eae088a, 32'h3e4f30ef} /* (10, 10, 8) {real, imag} */,
  {32'hbe5804ea, 32'hbe3ea2dc} /* (10, 10, 7) {real, imag} */,
  {32'h3da83776, 32'h3f767f42} /* (10, 10, 6) {real, imag} */,
  {32'hbdab4a98, 32'h3e57adaa} /* (10, 10, 5) {real, imag} */,
  {32'h3d9825ee, 32'h3c1b75d0} /* (10, 10, 4) {real, imag} */,
  {32'h3f0d75af, 32'h3e868f18} /* (10, 10, 3) {real, imag} */,
  {32'h3eb895e7, 32'hbe193912} /* (10, 10, 2) {real, imag} */,
  {32'h3e59c25e, 32'hbf108b20} /* (10, 10, 1) {real, imag} */,
  {32'h3e613321, 32'hbecb08e4} /* (10, 10, 0) {real, imag} */,
  {32'hbe65a079, 32'h3edb8d0e} /* (10, 9, 31) {real, imag} */,
  {32'h3d9dce12, 32'hbe1385a6} /* (10, 9, 30) {real, imag} */,
  {32'h3dbfb233, 32'h3f0e6b00} /* (10, 9, 29) {real, imag} */,
  {32'h3f14934c, 32'hbf029b66} /* (10, 9, 28) {real, imag} */,
  {32'h3f0f3cf5, 32'hbee7d96e} /* (10, 9, 27) {real, imag} */,
  {32'hbcf179d0, 32'h3dd685ff} /* (10, 9, 26) {real, imag} */,
  {32'hbeadcd50, 32'h3f0190c1} /* (10, 9, 25) {real, imag} */,
  {32'hbd16f18c, 32'hbe360382} /* (10, 9, 24) {real, imag} */,
  {32'h3d91e82e, 32'h3ecf8337} /* (10, 9, 23) {real, imag} */,
  {32'hbf1427e9, 32'h3e82f0e6} /* (10, 9, 22) {real, imag} */,
  {32'hbd853802, 32'hbca36c64} /* (10, 9, 21) {real, imag} */,
  {32'h3e49da7e, 32'hbe8c08d7} /* (10, 9, 20) {real, imag} */,
  {32'h3deb7ec2, 32'hbe8cd24a} /* (10, 9, 19) {real, imag} */,
  {32'h3d4cee5c, 32'hbeb12e48} /* (10, 9, 18) {real, imag} */,
  {32'hbea82b3c, 32'h3f023df6} /* (10, 9, 17) {real, imag} */,
  {32'h3e079d7f, 32'h3dfdba8f} /* (10, 9, 16) {real, imag} */,
  {32'hbcaf4150, 32'h3eaf4e2e} /* (10, 9, 15) {real, imag} */,
  {32'hbdb635f4, 32'hbdbc833a} /* (10, 9, 14) {real, imag} */,
  {32'h3de1e7b6, 32'hbe9fb2e6} /* (10, 9, 13) {real, imag} */,
  {32'hbec5b78c, 32'h3dde6720} /* (10, 9, 12) {real, imag} */,
  {32'h3ec72496, 32'hbe2bf07f} /* (10, 9, 11) {real, imag} */,
  {32'h3e573946, 32'hbeb1deb1} /* (10, 9, 10) {real, imag} */,
  {32'hbcf29870, 32'hbe087d20} /* (10, 9, 9) {real, imag} */,
  {32'hbeb5bec8, 32'h3e809cb6} /* (10, 9, 8) {real, imag} */,
  {32'hbe922fa2, 32'h3ecefc3d} /* (10, 9, 7) {real, imag} */,
  {32'h3ee89094, 32'hbe5c2979} /* (10, 9, 6) {real, imag} */,
  {32'hbf522072, 32'h3ed7c20d} /* (10, 9, 5) {real, imag} */,
  {32'hbf06fc80, 32'hbe29addd} /* (10, 9, 4) {real, imag} */,
  {32'h3edda0d6, 32'h3e4f3848} /* (10, 9, 3) {real, imag} */,
  {32'h3e9e96bb, 32'hbcc981d0} /* (10, 9, 2) {real, imag} */,
  {32'hbead7b7c, 32'h3e3de6b8} /* (10, 9, 1) {real, imag} */,
  {32'h3e3517b8, 32'h3e56c3dc} /* (10, 9, 0) {real, imag} */,
  {32'hbfb24ca9, 32'hbe95a032} /* (10, 8, 31) {real, imag} */,
  {32'h3f518910, 32'hbe537ba4} /* (10, 8, 30) {real, imag} */,
  {32'hbf4fcd71, 32'hbeb1a35c} /* (10, 8, 29) {real, imag} */,
  {32'h3d94b4e0, 32'h3ee822cc} /* (10, 8, 28) {real, imag} */,
  {32'h3ea3aa99, 32'h3f2579c8} /* (10, 8, 27) {real, imag} */,
  {32'hbe3aa38a, 32'h3be81530} /* (10, 8, 26) {real, imag} */,
  {32'h3e66b0ee, 32'hbe1f6f35} /* (10, 8, 25) {real, imag} */,
  {32'h3e6bd6da, 32'h3dacd5d8} /* (10, 8, 24) {real, imag} */,
  {32'h39c02e00, 32'hbe1fece4} /* (10, 8, 23) {real, imag} */,
  {32'h3ea944f4, 32'h3f022d24} /* (10, 8, 22) {real, imag} */,
  {32'hbf43b31c, 32'h3ec361e6} /* (10, 8, 21) {real, imag} */,
  {32'hbe4eebb0, 32'h3efd0eab} /* (10, 8, 20) {real, imag} */,
  {32'h3e2f29d7, 32'hbe2352b2} /* (10, 8, 19) {real, imag} */,
  {32'h3e5aee5c, 32'hbd0d43ac} /* (10, 8, 18) {real, imag} */,
  {32'h3b5a7270, 32'hbdc904d4} /* (10, 8, 17) {real, imag} */,
  {32'h3e44da08, 32'h3d98bed6} /* (10, 8, 16) {real, imag} */,
  {32'hbe497abf, 32'hbcc3a9f2} /* (10, 8, 15) {real, imag} */,
  {32'h3e5f11f0, 32'hbe8ae8e6} /* (10, 8, 14) {real, imag} */,
  {32'hbf088a74, 32'h3dca7901} /* (10, 8, 13) {real, imag} */,
  {32'h3ef1e022, 32'h3c496a18} /* (10, 8, 12) {real, imag} */,
  {32'h3e807f1a, 32'h3e3e2169} /* (10, 8, 11) {real, imag} */,
  {32'h3e3573bc, 32'h3e8ba8b5} /* (10, 8, 10) {real, imag} */,
  {32'hbeb8d2d8, 32'h3ebc13a2} /* (10, 8, 9) {real, imag} */,
  {32'h3e687609, 32'h3d9fe71c} /* (10, 8, 8) {real, imag} */,
  {32'h3f52ab84, 32'h3e7806b1} /* (10, 8, 7) {real, imag} */,
  {32'h3ebd43ec, 32'h3e46fdc7} /* (10, 8, 6) {real, imag} */,
  {32'h3ed45845, 32'hbeb2d86a} /* (10, 8, 5) {real, imag} */,
  {32'hbf18bc52, 32'hbd4fee58} /* (10, 8, 4) {real, imag} */,
  {32'hbd69c1f0, 32'h3d844dea} /* (10, 8, 3) {real, imag} */,
  {32'h3f66be6d, 32'h3ea10aa6} /* (10, 8, 2) {real, imag} */,
  {32'hbf2d2c34, 32'hbf20f196} /* (10, 8, 1) {real, imag} */,
  {32'hbe707ef0, 32'hbd8f89fc} /* (10, 8, 0) {real, imag} */,
  {32'h3f345426, 32'h3f33471e} /* (10, 7, 31) {real, imag} */,
  {32'hbecbf404, 32'hbf4c03fe} /* (10, 7, 30) {real, imag} */,
  {32'hbf436b20, 32'h3f7f86b0} /* (10, 7, 29) {real, imag} */,
  {32'h3d660260, 32'h3e7d965e} /* (10, 7, 28) {real, imag} */,
  {32'hbe8c15e7, 32'h3e31358c} /* (10, 7, 27) {real, imag} */,
  {32'h3d1aec8c, 32'h3c5979c0} /* (10, 7, 26) {real, imag} */,
  {32'h3e763c32, 32'hbe9856da} /* (10, 7, 25) {real, imag} */,
  {32'hbf246fb4, 32'h3da1a142} /* (10, 7, 24) {real, imag} */,
  {32'hbf06f702, 32'hbee9e925} /* (10, 7, 23) {real, imag} */,
  {32'h3e3a942b, 32'hbd83dab0} /* (10, 7, 22) {real, imag} */,
  {32'h3edbf115, 32'h3e5c1bf8} /* (10, 7, 21) {real, imag} */,
  {32'hbf04d64e, 32'hbe94327a} /* (10, 7, 20) {real, imag} */,
  {32'h3e94a0c8, 32'hbc7d6268} /* (10, 7, 19) {real, imag} */,
  {32'h3e0dbfbd, 32'h3d05f2dc} /* (10, 7, 18) {real, imag} */,
  {32'hbe9373db, 32'h3ca716b4} /* (10, 7, 17) {real, imag} */,
  {32'h3e2c5d66, 32'h3e1f3b01} /* (10, 7, 16) {real, imag} */,
  {32'hbde49754, 32'h3dc2f983} /* (10, 7, 15) {real, imag} */,
  {32'hbe2f21c1, 32'h3e37241a} /* (10, 7, 14) {real, imag} */,
  {32'hbe11c783, 32'h3f0c4352} /* (10, 7, 13) {real, imag} */,
  {32'hbdcdaff6, 32'hbe7992ea} /* (10, 7, 12) {real, imag} */,
  {32'h3e847a21, 32'h3d88cd62} /* (10, 7, 11) {real, imag} */,
  {32'hbe912bac, 32'hbf0bc44e} /* (10, 7, 10) {real, imag} */,
  {32'h3e78411d, 32'h3e6b41af} /* (10, 7, 9) {real, imag} */,
  {32'hbe6a2445, 32'hbdf8ea24} /* (10, 7, 8) {real, imag} */,
  {32'h3ca3ec04, 32'h3e4a5ba0} /* (10, 7, 7) {real, imag} */,
  {32'h3f2d079d, 32'hbec7d92e} /* (10, 7, 6) {real, imag} */,
  {32'hbebc49d7, 32'hbef34e13} /* (10, 7, 5) {real, imag} */,
  {32'h3e899ee6, 32'hbd5119ac} /* (10, 7, 4) {real, imag} */,
  {32'h3e2d01ea, 32'h3c9be220} /* (10, 7, 3) {real, imag} */,
  {32'hbf6f7fec, 32'h3e2fa876} /* (10, 7, 2) {real, imag} */,
  {32'h3e91935c, 32'h3f849c11} /* (10, 7, 1) {real, imag} */,
  {32'h3e1304cd, 32'hbe56311a} /* (10, 7, 0) {real, imag} */,
  {32'h3e5830fb, 32'hbf6faceb} /* (10, 6, 31) {real, imag} */,
  {32'h3e33ca98, 32'hbf179fa5} /* (10, 6, 30) {real, imag} */,
  {32'h3eb775b0, 32'h3e630794} /* (10, 6, 29) {real, imag} */,
  {32'h3f055990, 32'hbef45ae2} /* (10, 6, 28) {real, imag} */,
  {32'hbdf34e34, 32'hbf026ce0} /* (10, 6, 27) {real, imag} */,
  {32'h3f0ce352, 32'hbdc80454} /* (10, 6, 26) {real, imag} */,
  {32'h3de9f31a, 32'h3d3ea0aa} /* (10, 6, 25) {real, imag} */,
  {32'hbf0733ec, 32'hbd9e231a} /* (10, 6, 24) {real, imag} */,
  {32'h3f1723af, 32'h3f3aa62b} /* (10, 6, 23) {real, imag} */,
  {32'hbec9291f, 32'hbe9e04d6} /* (10, 6, 22) {real, imag} */,
  {32'h3f04eafa, 32'h3dc7a064} /* (10, 6, 21) {real, imag} */,
  {32'h3e307835, 32'hbdacd542} /* (10, 6, 20) {real, imag} */,
  {32'h3df485ac, 32'h3e8f34d3} /* (10, 6, 19) {real, imag} */,
  {32'h3edc0d4e, 32'h3e228c80} /* (10, 6, 18) {real, imag} */,
  {32'hbe4f61ad, 32'h3eb07e25} /* (10, 6, 17) {real, imag} */,
  {32'hbe4e252f, 32'h3e3410c8} /* (10, 6, 16) {real, imag} */,
  {32'hbe8d7742, 32'hbea4c742} /* (10, 6, 15) {real, imag} */,
  {32'h3e160ce0, 32'h3e18a832} /* (10, 6, 14) {real, imag} */,
  {32'h3e575e53, 32'h3c185e58} /* (10, 6, 13) {real, imag} */,
  {32'h3e3c5ec8, 32'h3d35c8d8} /* (10, 6, 12) {real, imag} */,
  {32'hbd415018, 32'hbdbb5f55} /* (10, 6, 11) {real, imag} */,
  {32'hbea864fe, 32'hbf0a5a38} /* (10, 6, 10) {real, imag} */,
  {32'hbe575db9, 32'hbeada22c} /* (10, 6, 9) {real, imag} */,
  {32'h3eb2085c, 32'hbecd03a0} /* (10, 6, 8) {real, imag} */,
  {32'h3e5b68c6, 32'h3c9a1a74} /* (10, 6, 7) {real, imag} */,
  {32'h3e880f86, 32'h3e7865d0} /* (10, 6, 6) {real, imag} */,
  {32'h3ef51b72, 32'h3f10de38} /* (10, 6, 5) {real, imag} */,
  {32'hbef0f791, 32'h3e2dc047} /* (10, 6, 4) {real, imag} */,
  {32'hbf0660e2, 32'h3e99004f} /* (10, 6, 3) {real, imag} */,
  {32'h3e340756, 32'hbf653a70} /* (10, 6, 2) {real, imag} */,
  {32'h3e12ea6f, 32'h3de0ba35} /* (10, 6, 1) {real, imag} */,
  {32'h3ef69ea5, 32'h3f890978} /* (10, 6, 0) {real, imag} */,
  {32'hc06abc8a, 32'hbf8d0e4b} /* (10, 5, 31) {real, imag} */,
  {32'h3f262202, 32'h3d3336e4} /* (10, 5, 30) {real, imag} */,
  {32'h3e632c50, 32'hbe2e0a9c} /* (10, 5, 29) {real, imag} */,
  {32'hbf18c64c, 32'h3fa4a9bc} /* (10, 5, 28) {real, imag} */,
  {32'hbca065c0, 32'h3f089e1a} /* (10, 5, 27) {real, imag} */,
  {32'h3d16d8a6, 32'hbe2ccbba} /* (10, 5, 26) {real, imag} */,
  {32'hbe8b137d, 32'h3eaaa6b6} /* (10, 5, 25) {real, imag} */,
  {32'hbe7d51ed, 32'hbf4e30a1} /* (10, 5, 24) {real, imag} */,
  {32'hbe7c6160, 32'h3f2be7ec} /* (10, 5, 23) {real, imag} */,
  {32'hbcf08d80, 32'hbf06e724} /* (10, 5, 22) {real, imag} */,
  {32'h3eb941ec, 32'hbf0fbac8} /* (10, 5, 21) {real, imag} */,
  {32'h3ccb6310, 32'hbe089820} /* (10, 5, 20) {real, imag} */,
  {32'hbe251228, 32'hbe947946} /* (10, 5, 19) {real, imag} */,
  {32'hbeb46b8a, 32'hbf08a1de} /* (10, 5, 18) {real, imag} */,
  {32'h3d872c74, 32'hbecef872} /* (10, 5, 17) {real, imag} */,
  {32'hbeb65de8, 32'hbbf428e0} /* (10, 5, 16) {real, imag} */,
  {32'hbecc0665, 32'h3eb8def2} /* (10, 5, 15) {real, imag} */,
  {32'h3d50c5a8, 32'h3f0303a3} /* (10, 5, 14) {real, imag} */,
  {32'h3ef04e62, 32'h3dc5caa6} /* (10, 5, 13) {real, imag} */,
  {32'h3eb04136, 32'hbcd58a98} /* (10, 5, 12) {real, imag} */,
  {32'hbebe69ec, 32'hbdbb47d4} /* (10, 5, 11) {real, imag} */,
  {32'hbdcc3ce4, 32'h3e7836f4} /* (10, 5, 10) {real, imag} */,
  {32'h3e0065c7, 32'hbd4b01ae} /* (10, 5, 9) {real, imag} */,
  {32'h3e13ef7c, 32'h3f2614c8} /* (10, 5, 8) {real, imag} */,
  {32'h3e61c7d1, 32'hbeecdcec} /* (10, 5, 7) {real, imag} */,
  {32'hbec2a20a, 32'h3e36320f} /* (10, 5, 6) {real, imag} */,
  {32'h3eeb48f2, 32'h3dca52fc} /* (10, 5, 5) {real, imag} */,
  {32'hbec98c26, 32'hbdec0e60} /* (10, 5, 4) {real, imag} */,
  {32'hbd0781a6, 32'h3e67cf3e} /* (10, 5, 3) {real, imag} */,
  {32'h3e358d21, 32'h3fcf3922} /* (10, 5, 2) {real, imag} */,
  {32'hbf397270, 32'hc016f74f} /* (10, 5, 1) {real, imag} */,
  {32'hbfffea3c, 32'hbf2f539a} /* (10, 5, 0) {real, imag} */,
  {32'h3fcfee04, 32'h40431e08} /* (10, 4, 31) {real, imag} */,
  {32'hc0531cbd, 32'hbfde677d} /* (10, 4, 30) {real, imag} */,
  {32'hbea2bd6f, 32'hbe9e0276} /* (10, 4, 29) {real, imag} */,
  {32'h3f59b136, 32'hbd1431c0} /* (10, 4, 28) {real, imag} */,
  {32'hbf3df03a, 32'hbdb74726} /* (10, 4, 27) {real, imag} */,
  {32'hbf42a438, 32'h3f764a91} /* (10, 4, 26) {real, imag} */,
  {32'h3f0a8bbe, 32'hbea248d0} /* (10, 4, 25) {real, imag} */,
  {32'h3e7a51c2, 32'hbf32c919} /* (10, 4, 24) {real, imag} */,
  {32'h3f818976, 32'h3daa7794} /* (10, 4, 23) {real, imag} */,
  {32'hbd7cab1e, 32'hbecc7819} /* (10, 4, 22) {real, imag} */,
  {32'h3d9a743e, 32'hbec84bda} /* (10, 4, 21) {real, imag} */,
  {32'hbd26e504, 32'h3e22caea} /* (10, 4, 20) {real, imag} */,
  {32'hbda2d4be, 32'h3dfe574f} /* (10, 4, 19) {real, imag} */,
  {32'hbef985ac, 32'hbe54fb4d} /* (10, 4, 18) {real, imag} */,
  {32'hbce94099, 32'h3e9789d1} /* (10, 4, 17) {real, imag} */,
  {32'hbe412340, 32'h3e3e4c8e} /* (10, 4, 16) {real, imag} */,
  {32'hbef15748, 32'h3dc2e7de} /* (10, 4, 15) {real, imag} */,
  {32'h3ecb1034, 32'hbe51dd42} /* (10, 4, 14) {real, imag} */,
  {32'h3e998148, 32'hbe35d58a} /* (10, 4, 13) {real, imag} */,
  {32'hbd55ee12, 32'h3e80befa} /* (10, 4, 12) {real, imag} */,
  {32'h3ead264f, 32'hbf24f36a} /* (10, 4, 11) {real, imag} */,
  {32'h3e4785c2, 32'h3e36f94a} /* (10, 4, 10) {real, imag} */,
  {32'h3ea8f3dc, 32'h3cc6fc50} /* (10, 4, 9) {real, imag} */,
  {32'hbe7a4f8a, 32'hbf15bba6} /* (10, 4, 8) {real, imag} */,
  {32'hbe0ea97a, 32'hbef0f572} /* (10, 4, 7) {real, imag} */,
  {32'hbe8e99b2, 32'h3e708c46} /* (10, 4, 6) {real, imag} */,
  {32'h3f3b4502, 32'hbf6a884e} /* (10, 4, 5) {real, imag} */,
  {32'h3e83c62a, 32'h3fad6279} /* (10, 4, 4) {real, imag} */,
  {32'hbf3e0e15, 32'h3f48c00c} /* (10, 4, 3) {real, imag} */,
  {32'hbff23e65, 32'hc0067505} /* (10, 4, 2) {real, imag} */,
  {32'h40a0d659, 32'h3f74a87c} /* (10, 4, 1) {real, imag} */,
  {32'h3f8e4851, 32'h3f48d2d6} /* (10, 4, 0) {real, imag} */,
  {32'hc0932d8f, 32'h40169b15} /* (10, 3, 31) {real, imag} */,
  {32'h400616b9, 32'hc086af0b} /* (10, 3, 30) {real, imag} */,
  {32'hbf0d50d6, 32'hbeeaafbd} /* (10, 3, 29) {real, imag} */,
  {32'h3fe266e6, 32'h3f71744a} /* (10, 3, 28) {real, imag} */,
  {32'hbfa50c8d, 32'h3e98a6f2} /* (10, 3, 27) {real, imag} */,
  {32'h3e90f1bc, 32'h3eccc7d7} /* (10, 3, 26) {real, imag} */,
  {32'hbda912a0, 32'h3ecd37e6} /* (10, 3, 25) {real, imag} */,
  {32'h3ecfb88f, 32'h3c9aa348} /* (10, 3, 24) {real, imag} */,
  {32'hbea5ea66, 32'h3d78f1ec} /* (10, 3, 23) {real, imag} */,
  {32'hbf4fb06f, 32'hbe81a298} /* (10, 3, 22) {real, imag} */,
  {32'h3e05c79c, 32'h3ecb789a} /* (10, 3, 21) {real, imag} */,
  {32'hbe4069a9, 32'hbde3beb6} /* (10, 3, 20) {real, imag} */,
  {32'hbdd0782a, 32'h3e0ed0de} /* (10, 3, 19) {real, imag} */,
  {32'h3bbf6c60, 32'hbe661e3c} /* (10, 3, 18) {real, imag} */,
  {32'h3e78e119, 32'hbea7a2b7} /* (10, 3, 17) {real, imag} */,
  {32'h3e80181d, 32'hbea35781} /* (10, 3, 16) {real, imag} */,
  {32'h3ece35d1, 32'hbdf7aef0} /* (10, 3, 15) {real, imag} */,
  {32'h3db7676e, 32'hbf03083f} /* (10, 3, 14) {real, imag} */,
  {32'hbdf93449, 32'hbe823aba} /* (10, 3, 13) {real, imag} */,
  {32'h3e82f34d, 32'hbef44d4e} /* (10, 3, 12) {real, imag} */,
  {32'h3e46ee46, 32'h3e9d725a} /* (10, 3, 11) {real, imag} */,
  {32'h3ec3d934, 32'h3f0a43c2} /* (10, 3, 10) {real, imag} */,
  {32'h3e30e5d8, 32'hbe271cfc} /* (10, 3, 9) {real, imag} */,
  {32'hbe28a9cd, 32'h3ecd286b} /* (10, 3, 8) {real, imag} */,
  {32'hbf3941ad, 32'h3ddb583a} /* (10, 3, 7) {real, imag} */,
  {32'hbe131ff0, 32'hbda8e1e6} /* (10, 3, 6) {real, imag} */,
  {32'hbee41416, 32'h3e23e9b0} /* (10, 3, 5) {real, imag} */,
  {32'hbf808b65, 32'h3ec21998} /* (10, 3, 4) {real, imag} */,
  {32'hbf62777a, 32'h3f3f6ded} /* (10, 3, 3) {real, imag} */,
  {32'hbe89bafa, 32'hc03cc3f5} /* (10, 3, 2) {real, imag} */,
  {32'h4062072d, 32'h402f14e8} /* (10, 3, 1) {real, imag} */,
  {32'hbf0b8942, 32'h3ed3d01e} /* (10, 3, 0) {real, imag} */,
  {32'hc225fe8d, 32'hc01c5516} /* (10, 2, 31) {real, imag} */,
  {32'h419603b2, 32'hc0b75182} /* (10, 2, 30) {real, imag} */,
  {32'h3f9c33fc, 32'h3ef9fe47} /* (10, 2, 29) {real, imag} */,
  {32'hbf5745ae, 32'h4017b2b2} /* (10, 2, 28) {real, imag} */,
  {32'h3fecdb99, 32'hc003366a} /* (10, 2, 27) {real, imag} */,
  {32'h3edb121c, 32'hbeb1844a} /* (10, 2, 26) {real, imag} */,
  {32'hbd4eed28, 32'h3e84b9c6} /* (10, 2, 25) {real, imag} */,
  {32'h3f7fbe08, 32'hbf3e5976} /* (10, 2, 24) {real, imag} */,
  {32'hbed9558d, 32'h3efda11c} /* (10, 2, 23) {real, imag} */,
  {32'hbf3e6041, 32'hbdee3dcc} /* (10, 2, 22) {real, imag} */,
  {32'h3e825ba0, 32'hbf4d0b2e} /* (10, 2, 21) {real, imag} */,
  {32'hbd993ade, 32'h3ee4c944} /* (10, 2, 20) {real, imag} */,
  {32'hbe9bee8f, 32'h3ebb9980} /* (10, 2, 19) {real, imag} */,
  {32'h3edc69c6, 32'hbc7554c0} /* (10, 2, 18) {real, imag} */,
  {32'hbe9f4e31, 32'hbe2609e4} /* (10, 2, 17) {real, imag} */,
  {32'h3d4072d6, 32'hbc0ce4e4} /* (10, 2, 16) {real, imag} */,
  {32'h3e30702c, 32'hbdd96098} /* (10, 2, 15) {real, imag} */,
  {32'hbe5e5ca0, 32'hbe47287e} /* (10, 2, 14) {real, imag} */,
  {32'hbee26ec2, 32'hbd4fc3ce} /* (10, 2, 13) {real, imag} */,
  {32'h3c2f0bb0, 32'hbe3a3025} /* (10, 2, 12) {real, imag} */,
  {32'h3df65eba, 32'h3ef4724e} /* (10, 2, 11) {real, imag} */,
  {32'hbe85d3ce, 32'hbe9270b6} /* (10, 2, 10) {real, imag} */,
  {32'h3e24d237, 32'h3e96ef5e} /* (10, 2, 9) {real, imag} */,
  {32'h3e9e3d37, 32'h3ed981f6} /* (10, 2, 8) {real, imag} */,
  {32'hbe30361a, 32'h3e10cd6e} /* (10, 2, 7) {real, imag} */,
  {32'h3ea0cdd9, 32'hbebc4cc4} /* (10, 2, 6) {real, imag} */,
  {32'h3f38be07, 32'h4024d4b0} /* (10, 2, 5) {real, imag} */,
  {32'hc05a8845, 32'hbfa34d5f} /* (10, 2, 4) {real, imag} */,
  {32'h3e98f22c, 32'h3f3bb3fa} /* (10, 2, 3) {real, imag} */,
  {32'h41596382, 32'hc07b0336} /* (10, 2, 2) {real, imag} */,
  {32'hc1b96d1f, 32'h40c32882} /* (10, 2, 1) {real, imag} */,
  {32'hc1ba787e, 32'hc0483579} /* (10, 2, 0) {real, imag} */,
  {32'h425bfc61, 32'hc14114bf} /* (10, 1, 31) {real, imag} */,
  {32'hc148ff00, 32'h40035e8e} /* (10, 1, 30) {real, imag} */,
  {32'hbfbf9288, 32'hbec0efc8} /* (10, 1, 29) {real, imag} */,
  {32'h40240b94, 32'h4048fb02} /* (10, 1, 28) {real, imag} */,
  {32'hc02c58a1, 32'h3e316332} /* (10, 1, 27) {real, imag} */,
  {32'hbe439d6c, 32'h3f22217c} /* (10, 1, 26) {real, imag} */,
  {32'h3f1a37d0, 32'hbe3df30c} /* (10, 1, 25) {real, imag} */,
  {32'hbec17d14, 32'h3efe305e} /* (10, 1, 24) {real, imag} */,
  {32'hbec5b17c, 32'hbe1df8ba} /* (10, 1, 23) {real, imag} */,
  {32'h3efbaf31, 32'h3e619633} /* (10, 1, 22) {real, imag} */,
  {32'hbf190ec6, 32'h3f0a5b84} /* (10, 1, 21) {real, imag} */,
  {32'h3d80cd76, 32'h3f225556} /* (10, 1, 20) {real, imag} */,
  {32'h3eadb4a1, 32'hbe440fd4} /* (10, 1, 19) {real, imag} */,
  {32'hbe10a2dc, 32'h3f1a1f74} /* (10, 1, 18) {real, imag} */,
  {32'h3d11158e, 32'h3dcc2d37} /* (10, 1, 17) {real, imag} */,
  {32'h3e383cba, 32'h3e952a10} /* (10, 1, 16) {real, imag} */,
  {32'h3dd1caf9, 32'h3df32b67} /* (10, 1, 15) {real, imag} */,
  {32'hbf000dfd, 32'hbe059b5b} /* (10, 1, 14) {real, imag} */,
  {32'h3d8bff88, 32'h3ddfbd1d} /* (10, 1, 13) {real, imag} */,
  {32'hbe209591, 32'hbe33e00a} /* (10, 1, 12) {real, imag} */,
  {32'hbe0245ae, 32'hbf012527} /* (10, 1, 11) {real, imag} */,
  {32'hbf3840ff, 32'hbf264742} /* (10, 1, 10) {real, imag} */,
  {32'h3ed610f2, 32'h3ed36679} /* (10, 1, 9) {real, imag} */,
  {32'hbe4b65a5, 32'hbf9efba0} /* (10, 1, 8) {real, imag} */,
  {32'h3f4bec46, 32'h3dd85798} /* (10, 1, 7) {real, imag} */,
  {32'hbf72cde9, 32'hbee495df} /* (10, 1, 6) {real, imag} */,
  {32'hc018ff05, 32'hbfae35bf} /* (10, 1, 5) {real, imag} */,
  {32'h3f6e46f0, 32'h3f14ad6e} /* (10, 1, 4) {real, imag} */,
  {32'h3eba26f6, 32'h3f0fa254} /* (10, 1, 3) {real, imag} */,
  {32'hc1a6c6c3, 32'hc19153f9} /* (10, 1, 2) {real, imag} */,
  {32'h429efe91, 32'h422ba8a3} /* (10, 1, 1) {real, imag} */,
  {32'h4293f624, 32'h409af701} /* (10, 1, 0) {real, imag} */,
  {32'h42362b0a, 32'hc2130090} /* (10, 0, 31) {real, imag} */,
  {32'hc0ca9d4c, 32'h412fe09a} /* (10, 0, 30) {real, imag} */,
  {32'hc0017688, 32'h3f02c4d1} /* (10, 0, 29) {real, imag} */,
  {32'hbec4c8d5, 32'h3f4c18e6} /* (10, 0, 28) {real, imag} */,
  {32'hbfedba18, 32'h3f5be344} /* (10, 0, 27) {real, imag} */,
  {32'hbc787650, 32'h3e30d6e8} /* (10, 0, 26) {real, imag} */,
  {32'h3e937829, 32'hbed5b1c4} /* (10, 0, 25) {real, imag} */,
  {32'hbe02dc94, 32'h3f926efa} /* (10, 0, 24) {real, imag} */,
  {32'h3e533a04, 32'hbde3b507} /* (10, 0, 23) {real, imag} */,
  {32'h3e86aa57, 32'h3d954caa} /* (10, 0, 22) {real, imag} */,
  {32'h3d4badf6, 32'h3ec472e2} /* (10, 0, 21) {real, imag} */,
  {32'hbd0569cc, 32'hbc6e6f18} /* (10, 0, 20) {real, imag} */,
  {32'hbdf4a4ee, 32'hbf1b686a} /* (10, 0, 19) {real, imag} */,
  {32'h3dd8b5f0, 32'hbe4c7708} /* (10, 0, 18) {real, imag} */,
  {32'hbd778be0, 32'h3d1be7bc} /* (10, 0, 17) {real, imag} */,
  {32'hbeda7012, 32'h00000000} /* (10, 0, 16) {real, imag} */,
  {32'hbd778be0, 32'hbd1be7bc} /* (10, 0, 15) {real, imag} */,
  {32'h3dd8b5f0, 32'h3e4c7708} /* (10, 0, 14) {real, imag} */,
  {32'hbdf4a4ee, 32'h3f1b686a} /* (10, 0, 13) {real, imag} */,
  {32'hbd0569cc, 32'h3c6e6f18} /* (10, 0, 12) {real, imag} */,
  {32'h3d4badf6, 32'hbec472e2} /* (10, 0, 11) {real, imag} */,
  {32'h3e86aa57, 32'hbd954caa} /* (10, 0, 10) {real, imag} */,
  {32'h3e533a04, 32'h3de3b507} /* (10, 0, 9) {real, imag} */,
  {32'hbe02dc94, 32'hbf926efa} /* (10, 0, 8) {real, imag} */,
  {32'h3e937829, 32'h3ed5b1c4} /* (10, 0, 7) {real, imag} */,
  {32'hbc787650, 32'hbe30d6e8} /* (10, 0, 6) {real, imag} */,
  {32'hbfedba18, 32'hbf5be344} /* (10, 0, 5) {real, imag} */,
  {32'hbec4c8d5, 32'hbf4c18e6} /* (10, 0, 4) {real, imag} */,
  {32'hc0017688, 32'hbf02c4d1} /* (10, 0, 3) {real, imag} */,
  {32'hc0ca9d4c, 32'hc12fe09a} /* (10, 0, 2) {real, imag} */,
  {32'h42362b0a, 32'h42130090} /* (10, 0, 1) {real, imag} */,
  {32'h4299ca44, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h4299b1b4, 32'hc2209d10} /* (9, 31, 31) {real, imag} */,
  {32'hc19b750a, 32'h418b2cf5} /* (9, 31, 30) {real, imag} */,
  {32'hbef75210, 32'hbeededac} /* (9, 31, 29) {real, imag} */,
  {32'h400c7824, 32'hbea10898} /* (9, 31, 28) {real, imag} */,
  {32'hc0388f86, 32'h3f35d8cf} /* (9, 31, 27) {real, imag} */,
  {32'hbf9272ca, 32'h3edbcfb1} /* (9, 31, 26) {real, imag} */,
  {32'h3f07fa93, 32'h3e3fd081} /* (9, 31, 25) {real, imag} */,
  {32'hbe92a991, 32'h3f5873d2} /* (9, 31, 24) {real, imag} */,
  {32'h3c465ae0, 32'hbeb77dbe} /* (9, 31, 23) {real, imag} */,
  {32'hbf26cade, 32'h3ef3b006} /* (9, 31, 22) {real, imag} */,
  {32'h3dcec3a4, 32'h3f240c9a} /* (9, 31, 21) {real, imag} */,
  {32'h3e7cdd38, 32'h3f0a3c1d} /* (9, 31, 20) {real, imag} */,
  {32'h3ec8b3bf, 32'h3ce36a60} /* (9, 31, 19) {real, imag} */,
  {32'h3ddad65a, 32'h3e90be98} /* (9, 31, 18) {real, imag} */,
  {32'hbedaedf0, 32'hbe0217d0} /* (9, 31, 17) {real, imag} */,
  {32'hbd90715f, 32'hbe7c766a} /* (9, 31, 16) {real, imag} */,
  {32'h3c161ec4, 32'hbd40c49c} /* (9, 31, 15) {real, imag} */,
  {32'hbf030a4a, 32'hbf443cca} /* (9, 31, 14) {real, imag} */,
  {32'h3e098cc8, 32'h3ea3a916} /* (9, 31, 13) {real, imag} */,
  {32'h3ea4890c, 32'hbe8d52f6} /* (9, 31, 12) {real, imag} */,
  {32'hbf5d6582, 32'hbeb4f38a} /* (9, 31, 11) {real, imag} */,
  {32'hbddacc0c, 32'hbe2adedc} /* (9, 31, 10) {real, imag} */,
  {32'h3ecaca9c, 32'hbca45c50} /* (9, 31, 9) {real, imag} */,
  {32'hbf69ef22, 32'hbdf1dc1c} /* (9, 31, 8) {real, imag} */,
  {32'h3f967626, 32'h3f3868f7} /* (9, 31, 7) {real, imag} */,
  {32'hbf208e7c, 32'h3eb89bdc} /* (9, 31, 6) {real, imag} */,
  {32'hc0295a45, 32'h3f5c97f4} /* (9, 31, 5) {real, imag} */,
  {32'h401d877b, 32'hc040738a} /* (9, 31, 4) {real, imag} */,
  {32'hbfb36371, 32'h3f22051b} /* (9, 31, 3) {real, imag} */,
  {32'hc13bee4a, 32'hc00e708b} /* (9, 31, 2) {real, imag} */,
  {32'h4252283a, 32'h4153f00b} /* (9, 31, 1) {real, imag} */,
  {32'h42905eca, 32'hc0dc289a} /* (9, 31, 0) {real, imag} */,
  {32'hc1b2a101, 32'hc0c46f42} /* (9, 30, 31) {real, imag} */,
  {32'h4158527b, 32'h406c34d2} /* (9, 30, 30) {real, imag} */,
  {32'hbf0dac46, 32'hbeaf5658} /* (9, 30, 29) {real, imag} */,
  {32'hc038aad1, 32'h3fcab37a} /* (9, 30, 28) {real, imag} */,
  {32'h3fb90c3a, 32'hbfb1fd35} /* (9, 30, 27) {real, imag} */,
  {32'h3f02dcee, 32'h3eb37d9d} /* (9, 30, 26) {real, imag} */,
  {32'hbf5f366c, 32'h3d0f0c70} /* (9, 30, 25) {real, imag} */,
  {32'h3f10afbf, 32'hbe9f2e7b} /* (9, 30, 24) {real, imag} */,
  {32'h3e9d899e, 32'hbeb4fd31} /* (9, 30, 23) {real, imag} */,
  {32'hbeffd13e, 32'h3ec70152} /* (9, 30, 22) {real, imag} */,
  {32'h3e8e2894, 32'hbea7577c} /* (9, 30, 21) {real, imag} */,
  {32'h3e9d3200, 32'h3e3ca626} /* (9, 30, 20) {real, imag} */,
  {32'h3dc7ec5c, 32'h3c9b9480} /* (9, 30, 19) {real, imag} */,
  {32'hbdaec384, 32'hbe32e074} /* (9, 30, 18) {real, imag} */,
  {32'hbdba2220, 32'h3eac8000} /* (9, 30, 17) {real, imag} */,
  {32'h3e5eddd0, 32'h3e1b5aa5} /* (9, 30, 16) {real, imag} */,
  {32'hbe130a8a, 32'hbd47aecc} /* (9, 30, 15) {real, imag} */,
  {32'hbd77cdf2, 32'h3f63eb3d} /* (9, 30, 14) {real, imag} */,
  {32'h3e426e5c, 32'h3e137cb0} /* (9, 30, 13) {real, imag} */,
  {32'hbdbb6334, 32'hbe2abf42} /* (9, 30, 12) {real, imag} */,
  {32'hbe7b4764, 32'hba4078c0} /* (9, 30, 11) {real, imag} */,
  {32'h3d038d64, 32'hbde19436} /* (9, 30, 10) {real, imag} */,
  {32'h3eb5e4b7, 32'hbf10bdaf} /* (9, 30, 9) {real, imag} */,
  {32'h3f6ffc58, 32'h3f16d7ef} /* (9, 30, 8) {real, imag} */,
  {32'hbe99d8cb, 32'h3e4b52c9} /* (9, 30, 7) {real, imag} */,
  {32'h3ed40f24, 32'h3f1890a7} /* (9, 30, 6) {real, imag} */,
  {32'h402bba8f, 32'h3f8fb289} /* (9, 30, 5) {real, imag} */,
  {32'hbf06c26b, 32'hc012eebb} /* (9, 30, 4) {real, imag} */,
  {32'h3f1a4284, 32'hbfb0401d} /* (9, 30, 3) {real, imag} */,
  {32'h418f54ac, 32'h40b538f6} /* (9, 30, 2) {real, imag} */,
  {32'hc222fd64, 32'h3fc2606e} /* (9, 30, 1) {real, imag} */,
  {32'hc1aff663, 32'h4080b112} /* (9, 30, 0) {real, imag} */,
  {32'h40452f9a, 32'hc05115a2} /* (9, 29, 31) {real, imag} */,
  {32'hbcd755c0, 32'h404a9267} /* (9, 29, 30) {real, imag} */,
  {32'hbf7177e0, 32'hbe88571a} /* (9, 29, 29) {real, imag} */,
  {32'hbfa221b2, 32'hbdfff548} /* (9, 29, 28) {real, imag} */,
  {32'hbe59758c, 32'hbdf82040} /* (9, 29, 27) {real, imag} */,
  {32'hbc92e8c0, 32'hbf28b76b} /* (9, 29, 26) {real, imag} */,
  {32'hbe83746e, 32'h3e377d52} /* (9, 29, 25) {real, imag} */,
  {32'hbf4b02f4, 32'hbea48d92} /* (9, 29, 24) {real, imag} */,
  {32'hbb6c5a10, 32'hbe40f446} /* (9, 29, 23) {real, imag} */,
  {32'hbebcffc4, 32'hbed62576} /* (9, 29, 22) {real, imag} */,
  {32'hbdc5076c, 32'h3d165254} /* (9, 29, 21) {real, imag} */,
  {32'h3ee01a8e, 32'hbe50f065} /* (9, 29, 20) {real, imag} */,
  {32'hbdcb693a, 32'hbe6ca620} /* (9, 29, 19) {real, imag} */,
  {32'hbe2f22ad, 32'hbe34f981} /* (9, 29, 18) {real, imag} */,
  {32'h3e9df930, 32'hbe896487} /* (9, 29, 17) {real, imag} */,
  {32'h3dcf2860, 32'h3e4c41ff} /* (9, 29, 16) {real, imag} */,
  {32'h3e298de0, 32'h3ebcb9e8} /* (9, 29, 15) {real, imag} */,
  {32'h3e99840e, 32'hbe1a57d2} /* (9, 29, 14) {real, imag} */,
  {32'h3eaac4d1, 32'h3d868634} /* (9, 29, 13) {real, imag} */,
  {32'h3e35d577, 32'hbdbea28a} /* (9, 29, 12) {real, imag} */,
  {32'hbe1bd94e, 32'h3eb5716c} /* (9, 29, 11) {real, imag} */,
  {32'hbebfc771, 32'hbcd43014} /* (9, 29, 10) {real, imag} */,
  {32'hbe5acbc2, 32'hbe8e4e75} /* (9, 29, 9) {real, imag} */,
  {32'h3f0ce24b, 32'h3f10014e} /* (9, 29, 8) {real, imag} */,
  {32'hbf122f2b, 32'h3e42ea38} /* (9, 29, 7) {real, imag} */,
  {32'h3d14d3d8, 32'hbeda4ed6} /* (9, 29, 6) {real, imag} */,
  {32'hbfa4ce6e, 32'h3eba1917} /* (9, 29, 5) {real, imag} */,
  {32'h3f6f50c3, 32'hbe01faa6} /* (9, 29, 4) {real, imag} */,
  {32'h3d5336b4, 32'hbf6b199d} /* (9, 29, 3) {real, imag} */,
  {32'h400a0160, 32'h40aa8cc7} /* (9, 29, 2) {real, imag} */,
  {32'hc07eea4c, 32'hbfa78557} /* (9, 29, 1) {real, imag} */,
  {32'hbea0eb90, 32'h3f6257cc} /* (9, 29, 0) {real, imag} */,
  {32'h408dff05, 32'hbf894c94} /* (9, 28, 31) {real, imag} */,
  {32'hbfc694f6, 32'h40288ca7} /* (9, 28, 30) {real, imag} */,
  {32'hbf9c4e87, 32'hbfd32e9c} /* (9, 28, 29) {real, imag} */,
  {32'h3eeaa38e, 32'hbf1dab8d} /* (9, 28, 28) {real, imag} */,
  {32'hbe500e40, 32'h3f5059f2} /* (9, 28, 27) {real, imag} */,
  {32'h3f3d1858, 32'h3d9e1364} /* (9, 28, 26) {real, imag} */,
  {32'hbd5eb5e0, 32'h3effa0e4} /* (9, 28, 25) {real, imag} */,
  {32'hbe95bbe0, 32'h3e9c68a3} /* (9, 28, 24) {real, imag} */,
  {32'h3e325510, 32'h3e0f40c4} /* (9, 28, 23) {real, imag} */,
  {32'h3e9ae7a4, 32'hbe0fb2c9} /* (9, 28, 22) {real, imag} */,
  {32'h3e5a790f, 32'h3ead6fdd} /* (9, 28, 21) {real, imag} */,
  {32'hbf5897d5, 32'hbe8eb4ec} /* (9, 28, 20) {real, imag} */,
  {32'hbe0c0e3e, 32'h3e2fb75a} /* (9, 28, 19) {real, imag} */,
  {32'h3d2d2042, 32'h3e3dc6a5} /* (9, 28, 18) {real, imag} */,
  {32'h3e22a01a, 32'hbe00f911} /* (9, 28, 17) {real, imag} */,
  {32'hbe47b2e5, 32'hbd5ba0e2} /* (9, 28, 16) {real, imag} */,
  {32'h3e98a53c, 32'h3e21dc22} /* (9, 28, 15) {real, imag} */,
  {32'hbe87a3f4, 32'h3d9d2ee4} /* (9, 28, 14) {real, imag} */,
  {32'hbedf7d20, 32'h3f024abc} /* (9, 28, 13) {real, imag} */,
  {32'h3ef4b962, 32'h3d912bfa} /* (9, 28, 12) {real, imag} */,
  {32'hbda38ece, 32'hbf32aba0} /* (9, 28, 11) {real, imag} */,
  {32'hbe5f5969, 32'h3e0ba6f6} /* (9, 28, 10) {real, imag} */,
  {32'h3ee5f52a, 32'h3d8ffaf8} /* (9, 28, 9) {real, imag} */,
  {32'h3e016374, 32'h3ec259ce} /* (9, 28, 8) {real, imag} */,
  {32'h3ddb1766, 32'hbf0c45ad} /* (9, 28, 7) {real, imag} */,
  {32'hbedd4d0a, 32'hbea8cd71} /* (9, 28, 6) {real, imag} */,
  {32'hbf2f5c3e, 32'h3f3e297f} /* (9, 28, 5) {real, imag} */,
  {32'h3f83af83, 32'hbe37006e} /* (9, 28, 4) {real, imag} */,
  {32'hbed35150, 32'h3e9a7a75} /* (9, 28, 3) {real, imag} */,
  {32'hc03b769c, 32'h4018c6ae} /* (9, 28, 2) {real, imag} */,
  {32'h3f3382f6, 32'hc04c40c4} /* (9, 28, 1) {real, imag} */,
  {32'h3f94a618, 32'hbf419450} /* (9, 28, 0) {real, imag} */,
  {32'hbf8e53da, 32'h40183dde} /* (9, 27, 31) {real, imag} */,
  {32'h3f7aff09, 32'hbf9ee39a} /* (9, 27, 30) {real, imag} */,
  {32'hbf6dfd25, 32'h3ec1ee4b} /* (9, 27, 29) {real, imag} */,
  {32'hbeb0a827, 32'h3e1f1190} /* (9, 27, 28) {real, imag} */,
  {32'h3f9b9724, 32'hbebd4d47} /* (9, 27, 27) {real, imag} */,
  {32'hbe1e2312, 32'hbeab7902} /* (9, 27, 26) {real, imag} */,
  {32'hbe032666, 32'h3eec7b3a} /* (9, 27, 25) {real, imag} */,
  {32'hbb803680, 32'h3d49e728} /* (9, 27, 24) {real, imag} */,
  {32'h3e2298c5, 32'h3e441566} /* (9, 27, 23) {real, imag} */,
  {32'h3d8fa0ac, 32'hbf681e0d} /* (9, 27, 22) {real, imag} */,
  {32'hbd8cb252, 32'hbf0f4ff0} /* (9, 27, 21) {real, imag} */,
  {32'hbd1b9978, 32'hbd22a30f} /* (9, 27, 20) {real, imag} */,
  {32'hbda84551, 32'hbd754bd0} /* (9, 27, 19) {real, imag} */,
  {32'h3e9496c4, 32'h3cdce59c} /* (9, 27, 18) {real, imag} */,
  {32'h3e526ddc, 32'hbc6436b4} /* (9, 27, 17) {real, imag} */,
  {32'h3ebdd0d8, 32'hbc3d9e50} /* (9, 27, 16) {real, imag} */,
  {32'hbde7b16a, 32'hbe6ed38f} /* (9, 27, 15) {real, imag} */,
  {32'h3d59e90c, 32'h3d87e700} /* (9, 27, 14) {real, imag} */,
  {32'hbedefd1a, 32'hbea8249b} /* (9, 27, 13) {real, imag} */,
  {32'hbe9141a3, 32'h3df477c2} /* (9, 27, 12) {real, imag} */,
  {32'h3eab022b, 32'hbd8c35a6} /* (9, 27, 11) {real, imag} */,
  {32'hbf33b325, 32'h3bcd0100} /* (9, 27, 10) {real, imag} */,
  {32'h3e9501cb, 32'hbcbaa684} /* (9, 27, 9) {real, imag} */,
  {32'h3ebd15c2, 32'h3d889c91} /* (9, 27, 8) {real, imag} */,
  {32'hbe2c7bdc, 32'hbf211e4b} /* (9, 27, 7) {real, imag} */,
  {32'h3eac16aa, 32'hbf438d36} /* (9, 27, 6) {real, imag} */,
  {32'hbdfb17c8, 32'hbe909960} /* (9, 27, 5) {real, imag} */,
  {32'hbe85b0bb, 32'hbd3b7200} /* (9, 27, 4) {real, imag} */,
  {32'h3f1c6dff, 32'hbec5efd5} /* (9, 27, 3) {real, imag} */,
  {32'h3f048bb4, 32'h3e87af27} /* (9, 27, 2) {real, imag} */,
  {32'hc051ec08, 32'h3e01e296} /* (9, 27, 1) {real, imag} */,
  {32'hbfd9bfcc, 32'h3f6fe0a2} /* (9, 27, 0) {real, imag} */,
  {32'h3ea90938, 32'hbe9a57f6} /* (9, 26, 31) {real, imag} */,
  {32'hbf5ffff6, 32'h3f40c6d2} /* (9, 26, 30) {real, imag} */,
  {32'hbe607254, 32'h3e4d7805} /* (9, 26, 29) {real, imag} */,
  {32'h3eb292da, 32'h3d410dc0} /* (9, 26, 28) {real, imag} */,
  {32'h3e67392e, 32'h3bd6fd80} /* (9, 26, 27) {real, imag} */,
  {32'h3ed6bd63, 32'hbe806a9d} /* (9, 26, 26) {real, imag} */,
  {32'h3e42633a, 32'hbe302450} /* (9, 26, 25) {real, imag} */,
  {32'h3e5d23a8, 32'h3ea34e5d} /* (9, 26, 24) {real, imag} */,
  {32'hbd68a5fc, 32'hbde432de} /* (9, 26, 23) {real, imag} */,
  {32'hbdd745cc, 32'hbf296a98} /* (9, 26, 22) {real, imag} */,
  {32'h3edff534, 32'hbf31599c} /* (9, 26, 21) {real, imag} */,
  {32'hbf02cfed, 32'hbec014dc} /* (9, 26, 20) {real, imag} */,
  {32'hbc460770, 32'hbd7850f4} /* (9, 26, 19) {real, imag} */,
  {32'hbe1861d8, 32'h3e231c67} /* (9, 26, 18) {real, imag} */,
  {32'h3e9278fa, 32'hbe08cb0a} /* (9, 26, 17) {real, imag} */,
  {32'hbea97b59, 32'h3d971e7e} /* (9, 26, 16) {real, imag} */,
  {32'hbe3c3bb4, 32'hbe73f20d} /* (9, 26, 15) {real, imag} */,
  {32'h3dce8858, 32'hbea47d7c} /* (9, 26, 14) {real, imag} */,
  {32'h3e57ff22, 32'h3e8faeaa} /* (9, 26, 13) {real, imag} */,
  {32'h3cbc3738, 32'hbde2e628} /* (9, 26, 12) {real, imag} */,
  {32'h3e83c4a6, 32'hbe946f09} /* (9, 26, 11) {real, imag} */,
  {32'h3e595fcf, 32'h3ec2d8b2} /* (9, 26, 10) {real, imag} */,
  {32'h3e495adb, 32'hbebdbd84} /* (9, 26, 9) {real, imag} */,
  {32'hbe118b75, 32'hbdc1bd62} /* (9, 26, 8) {real, imag} */,
  {32'hbea1ca64, 32'hbd1de6e6} /* (9, 26, 7) {real, imag} */,
  {32'h3f31d271, 32'hbf278c22} /* (9, 26, 6) {real, imag} */,
  {32'hbe2df51d, 32'h3dff1a2c} /* (9, 26, 5) {real, imag} */,
  {32'h3f39c2ba, 32'h3f2820c9} /* (9, 26, 4) {real, imag} */,
  {32'hba710200, 32'hbedc52b8} /* (9, 26, 3) {real, imag} */,
  {32'h3e8c098d, 32'hbe25c617} /* (9, 26, 2) {real, imag} */,
  {32'h3d906338, 32'hbeec182d} /* (9, 26, 1) {real, imag} */,
  {32'h3d9f004c, 32'hbf1194ac} /* (9, 26, 0) {real, imag} */,
  {32'h3ba8d720, 32'hbf346930} /* (9, 25, 31) {real, imag} */,
  {32'hbe954f9d, 32'h3f50af36} /* (9, 25, 30) {real, imag} */,
  {32'hbd7318cc, 32'hbe24c9dc} /* (9, 25, 29) {real, imag} */,
  {32'h3da6d8df, 32'hbe980da2} /* (9, 25, 28) {real, imag} */,
  {32'h3f2e0abc, 32'hbe01ccb5} /* (9, 25, 27) {real, imag} */,
  {32'h3ce893f0, 32'h3e9cf9f4} /* (9, 25, 26) {real, imag} */,
  {32'h3e7c3dca, 32'h3eb65872} /* (9, 25, 25) {real, imag} */,
  {32'hbeb37814, 32'hbe3b3a40} /* (9, 25, 24) {real, imag} */,
  {32'h3e7d5ab0, 32'hbf0c4f5b} /* (9, 25, 23) {real, imag} */,
  {32'h3ea78658, 32'h3e651bba} /* (9, 25, 22) {real, imag} */,
  {32'h3e4e1327, 32'hbe18c76a} /* (9, 25, 21) {real, imag} */,
  {32'hbe8702ef, 32'hbd1d1b9a} /* (9, 25, 20) {real, imag} */,
  {32'h3e51304a, 32'h3f2a97e8} /* (9, 25, 19) {real, imag} */,
  {32'hbf0d5daf, 32'hbda7a090} /* (9, 25, 18) {real, imag} */,
  {32'hbec4446e, 32'hbe0ac34c} /* (9, 25, 17) {real, imag} */,
  {32'hbd90a314, 32'h3db4c2ca} /* (9, 25, 16) {real, imag} */,
  {32'h3eaeb7af, 32'hbd8ed740} /* (9, 25, 15) {real, imag} */,
  {32'h3da5c396, 32'h3e6a10f6} /* (9, 25, 14) {real, imag} */,
  {32'h3eb20fea, 32'hbea917ba} /* (9, 25, 13) {real, imag} */,
  {32'h3e6fbfe4, 32'hbeb56422} /* (9, 25, 12) {real, imag} */,
  {32'hbe8f11e6, 32'h3de9ed31} /* (9, 25, 11) {real, imag} */,
  {32'h3e0fe90a, 32'hbeb4339a} /* (9, 25, 10) {real, imag} */,
  {32'hbf3f03b2, 32'h3da4b61c} /* (9, 25, 9) {real, imag} */,
  {32'hbd203af8, 32'h3f29dd94} /* (9, 25, 8) {real, imag} */,
  {32'hbe15c019, 32'h3eda9bc7} /* (9, 25, 7) {real, imag} */,
  {32'hbd9429f6, 32'hbd8b1ec8} /* (9, 25, 6) {real, imag} */,
  {32'hbf264e32, 32'hbe9998ba} /* (9, 25, 5) {real, imag} */,
  {32'hbe85b476, 32'h3e5cacf0} /* (9, 25, 4) {real, imag} */,
  {32'hbe80d1fe, 32'hbe808979} /* (9, 25, 3) {real, imag} */,
  {32'h3cb320f0, 32'h3f456090} /* (9, 25, 2) {real, imag} */,
  {32'h3f0d0f0b, 32'hbec206ed} /* (9, 25, 1) {real, imag} */,
  {32'hbe13b8dd, 32'hbe392cb6} /* (9, 25, 0) {real, imag} */,
  {32'hbe409db9, 32'h3f0e2ef2} /* (9, 24, 31) {real, imag} */,
  {32'h3e5b9691, 32'h3ea6c05a} /* (9, 24, 30) {real, imag} */,
  {32'hbcb4bb00, 32'hbeb7909a} /* (9, 24, 29) {real, imag} */,
  {32'h3e659cee, 32'hbde04ecc} /* (9, 24, 28) {real, imag} */,
  {32'h3f21bb48, 32'h3daa1284} /* (9, 24, 27) {real, imag} */,
  {32'hbe335e82, 32'hbd1467ec} /* (9, 24, 26) {real, imag} */,
  {32'h3ee87c3a, 32'hbf87439c} /* (9, 24, 25) {real, imag} */,
  {32'hbed6b7f6, 32'hbf13374b} /* (9, 24, 24) {real, imag} */,
  {32'h3dd726ba, 32'hbeb8668b} /* (9, 24, 23) {real, imag} */,
  {32'hbe4d28c2, 32'hbded0bb8} /* (9, 24, 22) {real, imag} */,
  {32'hbe2638de, 32'h3dc91660} /* (9, 24, 21) {real, imag} */,
  {32'hbec2ac24, 32'h3d94dad1} /* (9, 24, 20) {real, imag} */,
  {32'h3d8e1b4c, 32'h3e531e45} /* (9, 24, 19) {real, imag} */,
  {32'hbe360709, 32'hbeb0e052} /* (9, 24, 18) {real, imag} */,
  {32'hbe855741, 32'hbb3de780} /* (9, 24, 17) {real, imag} */,
  {32'h3ea84177, 32'hbd88d2f0} /* (9, 24, 16) {real, imag} */,
  {32'hbe9cf51d, 32'h3f07981c} /* (9, 24, 15) {real, imag} */,
  {32'h3e343d0d, 32'hbe71d7cb} /* (9, 24, 14) {real, imag} */,
  {32'hbcd575a0, 32'hbe1d2aef} /* (9, 24, 13) {real, imag} */,
  {32'h3cf6592c, 32'h3de38db1} /* (9, 24, 12) {real, imag} */,
  {32'hbdef0b20, 32'hbeeaf8cc} /* (9, 24, 11) {real, imag} */,
  {32'hbe85869f, 32'hbe9d33b8} /* (9, 24, 10) {real, imag} */,
  {32'hbf44f950, 32'h3e2151ce} /* (9, 24, 9) {real, imag} */,
  {32'hbd901b68, 32'h3eabe38c} /* (9, 24, 8) {real, imag} */,
  {32'h3e515f48, 32'h3e02ce15} /* (9, 24, 7) {real, imag} */,
  {32'h3e1461b4, 32'h3f0e0432} /* (9, 24, 6) {real, imag} */,
  {32'h3d865b38, 32'h3c9a3428} /* (9, 24, 5) {real, imag} */,
  {32'h3e879894, 32'hbf735b23} /* (9, 24, 4) {real, imag} */,
  {32'h3d90dde7, 32'h3ee3fc8c} /* (9, 24, 3) {real, imag} */,
  {32'h3f79c2d7, 32'hbe95260e} /* (9, 24, 2) {real, imag} */,
  {32'hbfab9308, 32'h3f321bbd} /* (9, 24, 1) {real, imag} */,
  {32'hbf8b388c, 32'h3ec1f294} /* (9, 24, 0) {real, imag} */,
  {32'h3f51964f, 32'h3e87fbde} /* (9, 23, 31) {real, imag} */,
  {32'h3ee8f3cc, 32'h3ebb5eb7} /* (9, 23, 30) {real, imag} */,
  {32'h3ea90906, 32'hbebff948} /* (9, 23, 29) {real, imag} */,
  {32'hbf139144, 32'hbec81848} /* (9, 23, 28) {real, imag} */,
  {32'hbf148df5, 32'h3dbc8e90} /* (9, 23, 27) {real, imag} */,
  {32'hbe95a206, 32'hbec027aa} /* (9, 23, 26) {real, imag} */,
  {32'hbe6bc9de, 32'hbf0f8dec} /* (9, 23, 25) {real, imag} */,
  {32'h3ebfc2e9, 32'h3f0a8aa8} /* (9, 23, 24) {real, imag} */,
  {32'hbeab39a1, 32'h3dcf7b6e} /* (9, 23, 23) {real, imag} */,
  {32'h3f4839b3, 32'hbea276db} /* (9, 23, 22) {real, imag} */,
  {32'hbcf69a34, 32'h3e93a178} /* (9, 23, 21) {real, imag} */,
  {32'hbeb6e39d, 32'hbd0e6c98} /* (9, 23, 20) {real, imag} */,
  {32'hbe78d97a, 32'hbeb91768} /* (9, 23, 19) {real, imag} */,
  {32'h3d6ab22c, 32'hbd047d0a} /* (9, 23, 18) {real, imag} */,
  {32'h3de513d3, 32'h3ec68d6e} /* (9, 23, 17) {real, imag} */,
  {32'h3ead974e, 32'hbd4ffaca} /* (9, 23, 16) {real, imag} */,
  {32'hbd3aa008, 32'hbe422151} /* (9, 23, 15) {real, imag} */,
  {32'h3e5511a0, 32'hbcc0d170} /* (9, 23, 14) {real, imag} */,
  {32'hbf0e3a41, 32'hbf3287f4} /* (9, 23, 13) {real, imag} */,
  {32'hbdcdde10, 32'hbd958a28} /* (9, 23, 12) {real, imag} */,
  {32'hbebf1268, 32'h3dee6bd5} /* (9, 23, 11) {real, imag} */,
  {32'h3e263dcc, 32'h3eb4c2ee} /* (9, 23, 10) {real, imag} */,
  {32'h3dcaad82, 32'h3e4de7fe} /* (9, 23, 9) {real, imag} */,
  {32'hbebae645, 32'h3e8b0e76} /* (9, 23, 8) {real, imag} */,
  {32'h3e6a2840, 32'h3d93f88f} /* (9, 23, 7) {real, imag} */,
  {32'hbe08eafd, 32'h3d78cb20} /* (9, 23, 6) {real, imag} */,
  {32'hbdf21c05, 32'hbec97cd5} /* (9, 23, 5) {real, imag} */,
  {32'hbe0fa26c, 32'hbd8d6e22} /* (9, 23, 4) {real, imag} */,
  {32'h3eb408a2, 32'hbe6a9ccc} /* (9, 23, 3) {real, imag} */,
  {32'hbe7d5536, 32'h3f301132} /* (9, 23, 2) {real, imag} */,
  {32'hbe90f302, 32'hbf0b683c} /* (9, 23, 1) {real, imag} */,
  {32'h3e881a94, 32'h3f020bc7} /* (9, 23, 0) {real, imag} */,
  {32'h3ea33d98, 32'hbef32f6d} /* (9, 22, 31) {real, imag} */,
  {32'h3da215a1, 32'hbd15223e} /* (9, 22, 30) {real, imag} */,
  {32'h3f0c27ef, 32'h3c5b2690} /* (9, 22, 29) {real, imag} */,
  {32'hbedfd0b2, 32'hbcfc0638} /* (9, 22, 28) {real, imag} */,
  {32'hbe94ceee, 32'h3ece3614} /* (9, 22, 27) {real, imag} */,
  {32'h3df40717, 32'hbbd282e0} /* (9, 22, 26) {real, imag} */,
  {32'h3eeec109, 32'h3f0b2f41} /* (9, 22, 25) {real, imag} */,
  {32'h3e9bd2ab, 32'hbe4b51fd} /* (9, 22, 24) {real, imag} */,
  {32'h3c8a3250, 32'h3f131044} /* (9, 22, 23) {real, imag} */,
  {32'hbf4f2a5b, 32'hbc4ae300} /* (9, 22, 22) {real, imag} */,
  {32'h3e500520, 32'h3e8d35cc} /* (9, 22, 21) {real, imag} */,
  {32'hbe32f56f, 32'h3d904ae2} /* (9, 22, 20) {real, imag} */,
  {32'hbea58c60, 32'h3efed0e6} /* (9, 22, 19) {real, imag} */,
  {32'h3f3400d4, 32'hbf09e9f0} /* (9, 22, 18) {real, imag} */,
  {32'hbd86e7d6, 32'h3e1eccc1} /* (9, 22, 17) {real, imag} */,
  {32'hbe379a71, 32'h3ca849d0} /* (9, 22, 16) {real, imag} */,
  {32'h3ca8b8bc, 32'h3e779e3b} /* (9, 22, 15) {real, imag} */,
  {32'hbf0de962, 32'h3e8427ab} /* (9, 22, 14) {real, imag} */,
  {32'hbf2496b2, 32'h3e14d05a} /* (9, 22, 13) {real, imag} */,
  {32'hbce15188, 32'hbec1fef4} /* (9, 22, 12) {real, imag} */,
  {32'h3ee16c4a, 32'hbe17a936} /* (9, 22, 11) {real, imag} */,
  {32'h3e4f4308, 32'h3ea37fa5} /* (9, 22, 10) {real, imag} */,
  {32'hbce2ec48, 32'h3eb6caa0} /* (9, 22, 9) {real, imag} */,
  {32'h3e7fa908, 32'hbda4b358} /* (9, 22, 8) {real, imag} */,
  {32'hbe953db3, 32'hbdd09d0e} /* (9, 22, 7) {real, imag} */,
  {32'h3e838eeb, 32'h3dc69cf6} /* (9, 22, 6) {real, imag} */,
  {32'hbe00da64, 32'h3d170de8} /* (9, 22, 5) {real, imag} */,
  {32'hbea74539, 32'h3e351160} /* (9, 22, 4) {real, imag} */,
  {32'hbd63c370, 32'hbeb02d04} /* (9, 22, 3) {real, imag} */,
  {32'h3d36182e, 32'h3e63a9f0} /* (9, 22, 2) {real, imag} */,
  {32'h3f10603d, 32'h3ea02b35} /* (9, 22, 1) {real, imag} */,
  {32'hbf1d7a93, 32'hbe42dd4d} /* (9, 22, 0) {real, imag} */,
  {32'hbe657d9a, 32'h3ef29ca6} /* (9, 21, 31) {real, imag} */,
  {32'h3de3d485, 32'h3d2d276c} /* (9, 21, 30) {real, imag} */,
  {32'h3ea8dac4, 32'hbec34522} /* (9, 21, 29) {real, imag} */,
  {32'hbf12aa7e, 32'h3e4c5c3a} /* (9, 21, 28) {real, imag} */,
  {32'h3d5b916c, 32'hbe2c8542} /* (9, 21, 27) {real, imag} */,
  {32'h3e3d3c41, 32'h3e6499dd} /* (9, 21, 26) {real, imag} */,
  {32'hbe271438, 32'hbe02fca2} /* (9, 21, 25) {real, imag} */,
  {32'h3c60aec0, 32'hbeb6c532} /* (9, 21, 24) {real, imag} */,
  {32'hbe976cb5, 32'hbd55a670} /* (9, 21, 23) {real, imag} */,
  {32'hbe5c36e2, 32'hbdb7dd8a} /* (9, 21, 22) {real, imag} */,
  {32'hbe9f4117, 32'hbeecdde4} /* (9, 21, 21) {real, imag} */,
  {32'h3cc9d8f8, 32'h3e4ad478} /* (9, 21, 20) {real, imag} */,
  {32'h3e445724, 32'h3f05862d} /* (9, 21, 19) {real, imag} */,
  {32'h3bd86c00, 32'h3f70445d} /* (9, 21, 18) {real, imag} */,
  {32'h3ddd8ca2, 32'hbe671420} /* (9, 21, 17) {real, imag} */,
  {32'h3e4f5b26, 32'hbe983972} /* (9, 21, 16) {real, imag} */,
  {32'hbec9ee60, 32'h3d1f090b} /* (9, 21, 15) {real, imag} */,
  {32'h3cbe5aa0, 32'h3dfab20c} /* (9, 21, 14) {real, imag} */,
  {32'hbf181146, 32'hbe1d84ed} /* (9, 21, 13) {real, imag} */,
  {32'hbe8f9c8c, 32'h3eb2e161} /* (9, 21, 12) {real, imag} */,
  {32'h3eaf3a78, 32'hbef2a8d5} /* (9, 21, 11) {real, imag} */,
  {32'hbd025360, 32'hbf107dd4} /* (9, 21, 10) {real, imag} */,
  {32'h3ccb4390, 32'h3e19fbe2} /* (9, 21, 9) {real, imag} */,
  {32'h3e7c2b0e, 32'hbec49334} /* (9, 21, 8) {real, imag} */,
  {32'hbe5d9477, 32'h3e2a72a6} /* (9, 21, 7) {real, imag} */,
  {32'hbe17c05a, 32'h3d281e30} /* (9, 21, 6) {real, imag} */,
  {32'h3edc0d49, 32'hbe4795b8} /* (9, 21, 5) {real, imag} */,
  {32'h3ea1d3e2, 32'h3ef8e4d4} /* (9, 21, 4) {real, imag} */,
  {32'hbc821080, 32'hbf182141} /* (9, 21, 3) {real, imag} */,
  {32'h3dfdf1b8, 32'hbe0735ab} /* (9, 21, 2) {real, imag} */,
  {32'hbf2247c5, 32'h3ee88766} /* (9, 21, 1) {real, imag} */,
  {32'hbf3e043d, 32'h3e0cd588} /* (9, 21, 0) {real, imag} */,
  {32'h3d560cd4, 32'h3f031d6e} /* (9, 20, 31) {real, imag} */,
  {32'h3e9092e7, 32'h3e26c0a6} /* (9, 20, 30) {real, imag} */,
  {32'hbf21b6f6, 32'h3e8abe67} /* (9, 20, 29) {real, imag} */,
  {32'h3ed29958, 32'hbdfa9a4f} /* (9, 20, 28) {real, imag} */,
  {32'h3eba84b7, 32'hbecbe5c5} /* (9, 20, 27) {real, imag} */,
  {32'h3daa00a1, 32'hbe2abea6} /* (9, 20, 26) {real, imag} */,
  {32'hbf601c02, 32'h3eb5a725} /* (9, 20, 25) {real, imag} */,
  {32'hbecc63c6, 32'h3f21d086} /* (9, 20, 24) {real, imag} */,
  {32'h3de5c818, 32'hbbfcf830} /* (9, 20, 23) {real, imag} */,
  {32'hbd30a1f2, 32'h3eeb157b} /* (9, 20, 22) {real, imag} */,
  {32'h3c1b220c, 32'h3eabe35e} /* (9, 20, 21) {real, imag} */,
  {32'hbdbe7ef6, 32'h3d241738} /* (9, 20, 20) {real, imag} */,
  {32'hbe2af2cb, 32'h3ecc5bae} /* (9, 20, 19) {real, imag} */,
  {32'hbe6bbbce, 32'h3eb8770c} /* (9, 20, 18) {real, imag} */,
  {32'h3e3f0496, 32'hbea116fa} /* (9, 20, 17) {real, imag} */,
  {32'h3ccf6218, 32'hbece49be} /* (9, 20, 16) {real, imag} */,
  {32'h3c444378, 32'h3e413296} /* (9, 20, 15) {real, imag} */,
  {32'h3f24fdbe, 32'h3e900fef} /* (9, 20, 14) {real, imag} */,
  {32'hbea7c7be, 32'h3d74e84c} /* (9, 20, 13) {real, imag} */,
  {32'h3e25920b, 32'hbda99d92} /* (9, 20, 12) {real, imag} */,
  {32'h3dbcc150, 32'h3d87208a} /* (9, 20, 11) {real, imag} */,
  {32'h3e1011d6, 32'h3ebd90d3} /* (9, 20, 10) {real, imag} */,
  {32'h3e4406eb, 32'h3ecc2cac} /* (9, 20, 9) {real, imag} */,
  {32'hbf397102, 32'hbe45f8e8} /* (9, 20, 8) {real, imag} */,
  {32'h3f1ac234, 32'h3eb97f2a} /* (9, 20, 7) {real, imag} */,
  {32'hbee265ca, 32'hbdc6abaf} /* (9, 20, 6) {real, imag} */,
  {32'h3e96701f, 32'h3dfe2ba0} /* (9, 20, 5) {real, imag} */,
  {32'h3e85d2f1, 32'hbe26581b} /* (9, 20, 4) {real, imag} */,
  {32'hbe8f87ad, 32'hbe623f7c} /* (9, 20, 3) {real, imag} */,
  {32'h3e965e62, 32'h3e380b10} /* (9, 20, 2) {real, imag} */,
  {32'h3e2708ef, 32'h3e8b862d} /* (9, 20, 1) {real, imag} */,
  {32'h3d83d0ff, 32'hbea24e9a} /* (9, 20, 0) {real, imag} */,
  {32'hbc814318, 32'h3cae6ea0} /* (9, 19, 31) {real, imag} */,
  {32'h3dfce838, 32'hbc128740} /* (9, 19, 30) {real, imag} */,
  {32'hbd4e3dfe, 32'h3d512d54} /* (9, 19, 29) {real, imag} */,
  {32'h3cda5726, 32'hbe5b7154} /* (9, 19, 28) {real, imag} */,
  {32'h3e1517bb, 32'h3c8cadec} /* (9, 19, 27) {real, imag} */,
  {32'hbde5278a, 32'h3e8152e3} /* (9, 19, 26) {real, imag} */,
  {32'hbdffe130, 32'h3ec8f194} /* (9, 19, 25) {real, imag} */,
  {32'h3e09b365, 32'hbc81b7d0} /* (9, 19, 24) {real, imag} */,
  {32'hbdc385a7, 32'hbe902ba8} /* (9, 19, 23) {real, imag} */,
  {32'h3ed9abb0, 32'h3de4a862} /* (9, 19, 22) {real, imag} */,
  {32'hbeef50db, 32'h3c3c2ef8} /* (9, 19, 21) {real, imag} */,
  {32'hbe509110, 32'h3ea3fc48} /* (9, 19, 20) {real, imag} */,
  {32'h3cfc719a, 32'h3f1a9fe2} /* (9, 19, 19) {real, imag} */,
  {32'h3d2d6ea8, 32'hbd8407a4} /* (9, 19, 18) {real, imag} */,
  {32'h3e4a72ac, 32'hbeb37377} /* (9, 19, 17) {real, imag} */,
  {32'hbe9bdd34, 32'h3e23021a} /* (9, 19, 16) {real, imag} */,
  {32'h3e05e81a, 32'hbe7e6164} /* (9, 19, 15) {real, imag} */,
  {32'hbe569992, 32'hbebff6a9} /* (9, 19, 14) {real, imag} */,
  {32'h3e868832, 32'h3dbfce79} /* (9, 19, 13) {real, imag} */,
  {32'hbeb5a3f8, 32'hbe9e9e92} /* (9, 19, 12) {real, imag} */,
  {32'h3e883dcf, 32'h3ea90f2b} /* (9, 19, 11) {real, imag} */,
  {32'h3e22c20e, 32'h3d55160c} /* (9, 19, 10) {real, imag} */,
  {32'h3d01a880, 32'hbf251a62} /* (9, 19, 9) {real, imag} */,
  {32'hbd3bbcb9, 32'h3e266348} /* (9, 19, 8) {real, imag} */,
  {32'hbd385982, 32'h3e25a5ff} /* (9, 19, 7) {real, imag} */,
  {32'h3f0892e1, 32'h3e465662} /* (9, 19, 6) {real, imag} */,
  {32'h3ea3bb86, 32'h3e0c42ac} /* (9, 19, 5) {real, imag} */,
  {32'hbf09dbf3, 32'hbd087192} /* (9, 19, 4) {real, imag} */,
  {32'hbe548223, 32'hbda60bc6} /* (9, 19, 3) {real, imag} */,
  {32'h3cc11f30, 32'hbea02ff0} /* (9, 19, 2) {real, imag} */,
  {32'hbd118aa0, 32'h3df7d528} /* (9, 19, 1) {real, imag} */,
  {32'hbd961680, 32'h3ea95179} /* (9, 19, 0) {real, imag} */,
  {32'h3c185538, 32'h3ec16020} /* (9, 18, 31) {real, imag} */,
  {32'hbc895dc0, 32'h3e2ddac8} /* (9, 18, 30) {real, imag} */,
  {32'hbe50ef0a, 32'h3f175d2d} /* (9, 18, 29) {real, imag} */,
  {32'h3e141e55, 32'h3e014b97} /* (9, 18, 28) {real, imag} */,
  {32'hbe20826d, 32'h3db93c2a} /* (9, 18, 27) {real, imag} */,
  {32'hbc9fb7c8, 32'h3d020574} /* (9, 18, 26) {real, imag} */,
  {32'h3dd14bfb, 32'h3e6c2fd2} /* (9, 18, 25) {real, imag} */,
  {32'hbd724638, 32'hbde5b09e} /* (9, 18, 24) {real, imag} */,
  {32'h3c7850aa, 32'h3ebd3f9b} /* (9, 18, 23) {real, imag} */,
  {32'h3d4af9d8, 32'h3d7ea744} /* (9, 18, 22) {real, imag} */,
  {32'hbea13f18, 32'h3e841a31} /* (9, 18, 21) {real, imag} */,
  {32'h3d8b56be, 32'hbdca17d8} /* (9, 18, 20) {real, imag} */,
  {32'hbe429c40, 32'hbd705144} /* (9, 18, 19) {real, imag} */,
  {32'hbd434798, 32'h3d4d7216} /* (9, 18, 18) {real, imag} */,
  {32'h3c6c9a80, 32'hbe0a37c1} /* (9, 18, 17) {real, imag} */,
  {32'h3f1fcc36, 32'h3e425145} /* (9, 18, 16) {real, imag} */,
  {32'hbe88d54a, 32'hbdc64c2a} /* (9, 18, 15) {real, imag} */,
  {32'h3ede9881, 32'hbea29d08} /* (9, 18, 14) {real, imag} */,
  {32'hbde3dd9c, 32'hbe1b673b} /* (9, 18, 13) {real, imag} */,
  {32'hbe2397f9, 32'h3ea55073} /* (9, 18, 12) {real, imag} */,
  {32'h3ee08b89, 32'hbd91fc4a} /* (9, 18, 11) {real, imag} */,
  {32'h3e4ca8d2, 32'h3ec50ed4} /* (9, 18, 10) {real, imag} */,
  {32'hbe904790, 32'h3ea42777} /* (9, 18, 9) {real, imag} */,
  {32'h3f196520, 32'h3e446606} /* (9, 18, 8) {real, imag} */,
  {32'h3e99fd0e, 32'hbd65045d} /* (9, 18, 7) {real, imag} */,
  {32'h3d7fab80, 32'h3ec5fd48} /* (9, 18, 6) {real, imag} */,
  {32'h3e960144, 32'hbf04d019} /* (9, 18, 5) {real, imag} */,
  {32'h3e26af1d, 32'h3f0ff41c} /* (9, 18, 4) {real, imag} */,
  {32'h3da1380a, 32'hbe27399f} /* (9, 18, 3) {real, imag} */,
  {32'h3ebb4179, 32'h3e17e474} /* (9, 18, 2) {real, imag} */,
  {32'hbd0c0e90, 32'h3c3bbc60} /* (9, 18, 1) {real, imag} */,
  {32'hbde37268, 32'h3dbac67c} /* (9, 18, 0) {real, imag} */,
  {32'h3ca796b0, 32'hbe1aaf44} /* (9, 17, 31) {real, imag} */,
  {32'h3d8978fc, 32'h3e0f60da} /* (9, 17, 30) {real, imag} */,
  {32'h3e66fa50, 32'h3d8b008f} /* (9, 17, 29) {real, imag} */,
  {32'hbd9f8094, 32'hbcdbeff8} /* (9, 17, 28) {real, imag} */,
  {32'hbd7c3dba, 32'hbe6104cc} /* (9, 17, 27) {real, imag} */,
  {32'h3e365e4c, 32'hbe70c9c8} /* (9, 17, 26) {real, imag} */,
  {32'h3e8991a1, 32'hbe69294e} /* (9, 17, 25) {real, imag} */,
  {32'hbe858377, 32'hbebde941} /* (9, 17, 24) {real, imag} */,
  {32'h3e2a521a, 32'hbf0c442e} /* (9, 17, 23) {real, imag} */,
  {32'hbec8e88e, 32'h3e0fd35e} /* (9, 17, 22) {real, imag} */,
  {32'hbdd0ecc6, 32'h3eafd43e} /* (9, 17, 21) {real, imag} */,
  {32'hbcf25c58, 32'h3db47c3d} /* (9, 17, 20) {real, imag} */,
  {32'hbefff72b, 32'h3d82957f} /* (9, 17, 19) {real, imag} */,
  {32'h3e82e48d, 32'hbe8bc63e} /* (9, 17, 18) {real, imag} */,
  {32'hbea7d660, 32'h3e820f6d} /* (9, 17, 17) {real, imag} */,
  {32'hbd2522a2, 32'h3ec9e0ae} /* (9, 17, 16) {real, imag} */,
  {32'h3e194c50, 32'h3ca83448} /* (9, 17, 15) {real, imag} */,
  {32'h3e0221fb, 32'h3c57b660} /* (9, 17, 14) {real, imag} */,
  {32'h3ead267f, 32'h3e480a22} /* (9, 17, 13) {real, imag} */,
  {32'h3c3ec248, 32'h3e659767} /* (9, 17, 12) {real, imag} */,
  {32'hbe14dc14, 32'h3d1e84e4} /* (9, 17, 11) {real, imag} */,
  {32'hbe30fa66, 32'h3d05aed8} /* (9, 17, 10) {real, imag} */,
  {32'hbe2dd149, 32'hbe599b4c} /* (9, 17, 9) {real, imag} */,
  {32'h3d8b7e08, 32'hbe208d36} /* (9, 17, 8) {real, imag} */,
  {32'h3e0c981f, 32'hbd1fe508} /* (9, 17, 7) {real, imag} */,
  {32'hbe7b69c1, 32'h3ec87038} /* (9, 17, 6) {real, imag} */,
  {32'hbd2f5ea2, 32'hbd3495fa} /* (9, 17, 5) {real, imag} */,
  {32'h3da30b2b, 32'hbe0ee1e6} /* (9, 17, 4) {real, imag} */,
  {32'h3ddd3deb, 32'h3dec32e9} /* (9, 17, 3) {real, imag} */,
  {32'hbb5d3200, 32'h3ed12753} /* (9, 17, 2) {real, imag} */,
  {32'hbd41e1fc, 32'hbd729520} /* (9, 17, 1) {real, imag} */,
  {32'hbe9b1a58, 32'hbbacae00} /* (9, 17, 0) {real, imag} */,
  {32'hbdb34c11, 32'h3ea231cd} /* (9, 16, 31) {real, imag} */,
  {32'hbe90aa3c, 32'hbe776e1a} /* (9, 16, 30) {real, imag} */,
  {32'h3e29cdf6, 32'h3ddc1184} /* (9, 16, 29) {real, imag} */,
  {32'h3ddc25a0, 32'hbe8c1626} /* (9, 16, 28) {real, imag} */,
  {32'hbe7eb055, 32'hbe980731} /* (9, 16, 27) {real, imag} */,
  {32'hbdbb5791, 32'h3c438c30} /* (9, 16, 26) {real, imag} */,
  {32'h3e0105b2, 32'hbcf40510} /* (9, 16, 25) {real, imag} */,
  {32'h3d8716d4, 32'hbea15a09} /* (9, 16, 24) {real, imag} */,
  {32'hbd0f4316, 32'h3cd30130} /* (9, 16, 23) {real, imag} */,
  {32'hbe1b4fa0, 32'h3ed8dfc6} /* (9, 16, 22) {real, imag} */,
  {32'hbe1175c4, 32'hbe1faa8c} /* (9, 16, 21) {real, imag} */,
  {32'h3ecc489e, 32'hbe5b9380} /* (9, 16, 20) {real, imag} */,
  {32'h3eac45ca, 32'hbf07ed7a} /* (9, 16, 19) {real, imag} */,
  {32'hbe40f9ca, 32'hbdab1351} /* (9, 16, 18) {real, imag} */,
  {32'h3c1bd754, 32'h3ea5bc1e} /* (9, 16, 17) {real, imag} */,
  {32'h3e2d2dc8, 32'h00000000} /* (9, 16, 16) {real, imag} */,
  {32'h3c1bd754, 32'hbea5bc1e} /* (9, 16, 15) {real, imag} */,
  {32'hbe40f9ca, 32'h3dab1351} /* (9, 16, 14) {real, imag} */,
  {32'h3eac45ca, 32'h3f07ed7a} /* (9, 16, 13) {real, imag} */,
  {32'h3ecc489e, 32'h3e5b9380} /* (9, 16, 12) {real, imag} */,
  {32'hbe1175c4, 32'h3e1faa8c} /* (9, 16, 11) {real, imag} */,
  {32'hbe1b4fa0, 32'hbed8dfc6} /* (9, 16, 10) {real, imag} */,
  {32'hbd0f4316, 32'hbcd30130} /* (9, 16, 9) {real, imag} */,
  {32'h3d8716d4, 32'h3ea15a09} /* (9, 16, 8) {real, imag} */,
  {32'h3e0105b2, 32'h3cf40510} /* (9, 16, 7) {real, imag} */,
  {32'hbdbb5791, 32'hbc438c30} /* (9, 16, 6) {real, imag} */,
  {32'hbe7eb055, 32'h3e980731} /* (9, 16, 5) {real, imag} */,
  {32'h3ddc25a0, 32'h3e8c1626} /* (9, 16, 4) {real, imag} */,
  {32'h3e29cdf6, 32'hbddc1184} /* (9, 16, 3) {real, imag} */,
  {32'hbe90aa3c, 32'h3e776e1a} /* (9, 16, 2) {real, imag} */,
  {32'hbdb34c11, 32'hbea231cd} /* (9, 16, 1) {real, imag} */,
  {32'h3e1aab86, 32'h00000000} /* (9, 16, 0) {real, imag} */,
  {32'hbd41e1fc, 32'h3d729520} /* (9, 15, 31) {real, imag} */,
  {32'hbb5d3200, 32'hbed12753} /* (9, 15, 30) {real, imag} */,
  {32'h3ddd3deb, 32'hbdec32e9} /* (9, 15, 29) {real, imag} */,
  {32'h3da30b2b, 32'h3e0ee1e6} /* (9, 15, 28) {real, imag} */,
  {32'hbd2f5ea2, 32'h3d3495fa} /* (9, 15, 27) {real, imag} */,
  {32'hbe7b69c1, 32'hbec87038} /* (9, 15, 26) {real, imag} */,
  {32'h3e0c981f, 32'h3d1fe508} /* (9, 15, 25) {real, imag} */,
  {32'h3d8b7e08, 32'h3e208d36} /* (9, 15, 24) {real, imag} */,
  {32'hbe2dd149, 32'h3e599b4c} /* (9, 15, 23) {real, imag} */,
  {32'hbe30fa66, 32'hbd05aed8} /* (9, 15, 22) {real, imag} */,
  {32'hbe14dc14, 32'hbd1e84e4} /* (9, 15, 21) {real, imag} */,
  {32'h3c3ec248, 32'hbe659767} /* (9, 15, 20) {real, imag} */,
  {32'h3ead267f, 32'hbe480a22} /* (9, 15, 19) {real, imag} */,
  {32'h3e0221fb, 32'hbc57b660} /* (9, 15, 18) {real, imag} */,
  {32'h3e194c50, 32'hbca83448} /* (9, 15, 17) {real, imag} */,
  {32'hbd2522a2, 32'hbec9e0ae} /* (9, 15, 16) {real, imag} */,
  {32'hbea7d660, 32'hbe820f6d} /* (9, 15, 15) {real, imag} */,
  {32'h3e82e48d, 32'h3e8bc63e} /* (9, 15, 14) {real, imag} */,
  {32'hbefff72b, 32'hbd82957f} /* (9, 15, 13) {real, imag} */,
  {32'hbcf25c58, 32'hbdb47c3d} /* (9, 15, 12) {real, imag} */,
  {32'hbdd0ecc6, 32'hbeafd43e} /* (9, 15, 11) {real, imag} */,
  {32'hbec8e88e, 32'hbe0fd35e} /* (9, 15, 10) {real, imag} */,
  {32'h3e2a521a, 32'h3f0c442e} /* (9, 15, 9) {real, imag} */,
  {32'hbe858377, 32'h3ebde941} /* (9, 15, 8) {real, imag} */,
  {32'h3e8991a1, 32'h3e69294e} /* (9, 15, 7) {real, imag} */,
  {32'h3e365e4c, 32'h3e70c9c8} /* (9, 15, 6) {real, imag} */,
  {32'hbd7c3dba, 32'h3e6104cc} /* (9, 15, 5) {real, imag} */,
  {32'hbd9f8094, 32'h3cdbeff8} /* (9, 15, 4) {real, imag} */,
  {32'h3e66fa50, 32'hbd8b008f} /* (9, 15, 3) {real, imag} */,
  {32'h3d8978fc, 32'hbe0f60da} /* (9, 15, 2) {real, imag} */,
  {32'h3ca796b0, 32'h3e1aaf44} /* (9, 15, 1) {real, imag} */,
  {32'hbe9b1a58, 32'h3bacae00} /* (9, 15, 0) {real, imag} */,
  {32'hbd0c0e90, 32'hbc3bbc60} /* (9, 14, 31) {real, imag} */,
  {32'h3ebb4179, 32'hbe17e474} /* (9, 14, 30) {real, imag} */,
  {32'h3da1380a, 32'h3e27399f} /* (9, 14, 29) {real, imag} */,
  {32'h3e26af1d, 32'hbf0ff41c} /* (9, 14, 28) {real, imag} */,
  {32'h3e960144, 32'h3f04d019} /* (9, 14, 27) {real, imag} */,
  {32'h3d7fab80, 32'hbec5fd48} /* (9, 14, 26) {real, imag} */,
  {32'h3e99fd0e, 32'h3d65045d} /* (9, 14, 25) {real, imag} */,
  {32'h3f196520, 32'hbe446606} /* (9, 14, 24) {real, imag} */,
  {32'hbe904790, 32'hbea42777} /* (9, 14, 23) {real, imag} */,
  {32'h3e4ca8d2, 32'hbec50ed4} /* (9, 14, 22) {real, imag} */,
  {32'h3ee08b89, 32'h3d91fc4a} /* (9, 14, 21) {real, imag} */,
  {32'hbe2397f9, 32'hbea55073} /* (9, 14, 20) {real, imag} */,
  {32'hbde3dd9c, 32'h3e1b673b} /* (9, 14, 19) {real, imag} */,
  {32'h3ede9881, 32'h3ea29d08} /* (9, 14, 18) {real, imag} */,
  {32'hbe88d54a, 32'h3dc64c2a} /* (9, 14, 17) {real, imag} */,
  {32'h3f1fcc36, 32'hbe425145} /* (9, 14, 16) {real, imag} */,
  {32'h3c6c9a80, 32'h3e0a37c1} /* (9, 14, 15) {real, imag} */,
  {32'hbd434798, 32'hbd4d7216} /* (9, 14, 14) {real, imag} */,
  {32'hbe429c40, 32'h3d705144} /* (9, 14, 13) {real, imag} */,
  {32'h3d8b56be, 32'h3dca17d8} /* (9, 14, 12) {real, imag} */,
  {32'hbea13f18, 32'hbe841a31} /* (9, 14, 11) {real, imag} */,
  {32'h3d4af9d8, 32'hbd7ea744} /* (9, 14, 10) {real, imag} */,
  {32'h3c7850aa, 32'hbebd3f9b} /* (9, 14, 9) {real, imag} */,
  {32'hbd724638, 32'h3de5b09e} /* (9, 14, 8) {real, imag} */,
  {32'h3dd14bfb, 32'hbe6c2fd2} /* (9, 14, 7) {real, imag} */,
  {32'hbc9fb7c8, 32'hbd020574} /* (9, 14, 6) {real, imag} */,
  {32'hbe20826d, 32'hbdb93c2a} /* (9, 14, 5) {real, imag} */,
  {32'h3e141e55, 32'hbe014b97} /* (9, 14, 4) {real, imag} */,
  {32'hbe50ef0a, 32'hbf175d2d} /* (9, 14, 3) {real, imag} */,
  {32'hbc895dc0, 32'hbe2ddac8} /* (9, 14, 2) {real, imag} */,
  {32'h3c185538, 32'hbec16020} /* (9, 14, 1) {real, imag} */,
  {32'hbde37268, 32'hbdbac67c} /* (9, 14, 0) {real, imag} */,
  {32'hbd118aa0, 32'hbdf7d528} /* (9, 13, 31) {real, imag} */,
  {32'h3cc11f30, 32'h3ea02ff0} /* (9, 13, 30) {real, imag} */,
  {32'hbe548223, 32'h3da60bc6} /* (9, 13, 29) {real, imag} */,
  {32'hbf09dbf3, 32'h3d087192} /* (9, 13, 28) {real, imag} */,
  {32'h3ea3bb86, 32'hbe0c42ac} /* (9, 13, 27) {real, imag} */,
  {32'h3f0892e1, 32'hbe465662} /* (9, 13, 26) {real, imag} */,
  {32'hbd385982, 32'hbe25a5ff} /* (9, 13, 25) {real, imag} */,
  {32'hbd3bbcb9, 32'hbe266348} /* (9, 13, 24) {real, imag} */,
  {32'h3d01a880, 32'h3f251a62} /* (9, 13, 23) {real, imag} */,
  {32'h3e22c20e, 32'hbd55160c} /* (9, 13, 22) {real, imag} */,
  {32'h3e883dcf, 32'hbea90f2b} /* (9, 13, 21) {real, imag} */,
  {32'hbeb5a3f8, 32'h3e9e9e92} /* (9, 13, 20) {real, imag} */,
  {32'h3e868832, 32'hbdbfce79} /* (9, 13, 19) {real, imag} */,
  {32'hbe569992, 32'h3ebff6a9} /* (9, 13, 18) {real, imag} */,
  {32'h3e05e81a, 32'h3e7e6164} /* (9, 13, 17) {real, imag} */,
  {32'hbe9bdd34, 32'hbe23021a} /* (9, 13, 16) {real, imag} */,
  {32'h3e4a72ac, 32'h3eb37377} /* (9, 13, 15) {real, imag} */,
  {32'h3d2d6ea8, 32'h3d8407a4} /* (9, 13, 14) {real, imag} */,
  {32'h3cfc719a, 32'hbf1a9fe2} /* (9, 13, 13) {real, imag} */,
  {32'hbe509110, 32'hbea3fc48} /* (9, 13, 12) {real, imag} */,
  {32'hbeef50db, 32'hbc3c2ef8} /* (9, 13, 11) {real, imag} */,
  {32'h3ed9abb0, 32'hbde4a862} /* (9, 13, 10) {real, imag} */,
  {32'hbdc385a7, 32'h3e902ba8} /* (9, 13, 9) {real, imag} */,
  {32'h3e09b365, 32'h3c81b7d0} /* (9, 13, 8) {real, imag} */,
  {32'hbdffe130, 32'hbec8f194} /* (9, 13, 7) {real, imag} */,
  {32'hbde5278a, 32'hbe8152e3} /* (9, 13, 6) {real, imag} */,
  {32'h3e1517bb, 32'hbc8cadec} /* (9, 13, 5) {real, imag} */,
  {32'h3cda5726, 32'h3e5b7154} /* (9, 13, 4) {real, imag} */,
  {32'hbd4e3dfe, 32'hbd512d54} /* (9, 13, 3) {real, imag} */,
  {32'h3dfce838, 32'h3c128740} /* (9, 13, 2) {real, imag} */,
  {32'hbc814318, 32'hbcae6ea0} /* (9, 13, 1) {real, imag} */,
  {32'hbd961680, 32'hbea95179} /* (9, 13, 0) {real, imag} */,
  {32'h3e2708ef, 32'hbe8b862d} /* (9, 12, 31) {real, imag} */,
  {32'h3e965e62, 32'hbe380b10} /* (9, 12, 30) {real, imag} */,
  {32'hbe8f87ad, 32'h3e623f7c} /* (9, 12, 29) {real, imag} */,
  {32'h3e85d2f1, 32'h3e26581b} /* (9, 12, 28) {real, imag} */,
  {32'h3e96701f, 32'hbdfe2ba0} /* (9, 12, 27) {real, imag} */,
  {32'hbee265ca, 32'h3dc6abaf} /* (9, 12, 26) {real, imag} */,
  {32'h3f1ac234, 32'hbeb97f2a} /* (9, 12, 25) {real, imag} */,
  {32'hbf397102, 32'h3e45f8e8} /* (9, 12, 24) {real, imag} */,
  {32'h3e4406eb, 32'hbecc2cac} /* (9, 12, 23) {real, imag} */,
  {32'h3e1011d6, 32'hbebd90d3} /* (9, 12, 22) {real, imag} */,
  {32'h3dbcc150, 32'hbd87208a} /* (9, 12, 21) {real, imag} */,
  {32'h3e25920b, 32'h3da99d92} /* (9, 12, 20) {real, imag} */,
  {32'hbea7c7be, 32'hbd74e84c} /* (9, 12, 19) {real, imag} */,
  {32'h3f24fdbe, 32'hbe900fef} /* (9, 12, 18) {real, imag} */,
  {32'h3c444378, 32'hbe413296} /* (9, 12, 17) {real, imag} */,
  {32'h3ccf6218, 32'h3ece49be} /* (9, 12, 16) {real, imag} */,
  {32'h3e3f0496, 32'h3ea116fa} /* (9, 12, 15) {real, imag} */,
  {32'hbe6bbbce, 32'hbeb8770c} /* (9, 12, 14) {real, imag} */,
  {32'hbe2af2cb, 32'hbecc5bae} /* (9, 12, 13) {real, imag} */,
  {32'hbdbe7ef6, 32'hbd241738} /* (9, 12, 12) {real, imag} */,
  {32'h3c1b220c, 32'hbeabe35e} /* (9, 12, 11) {real, imag} */,
  {32'hbd30a1f2, 32'hbeeb157b} /* (9, 12, 10) {real, imag} */,
  {32'h3de5c818, 32'h3bfcf830} /* (9, 12, 9) {real, imag} */,
  {32'hbecc63c6, 32'hbf21d086} /* (9, 12, 8) {real, imag} */,
  {32'hbf601c02, 32'hbeb5a725} /* (9, 12, 7) {real, imag} */,
  {32'h3daa00a1, 32'h3e2abea6} /* (9, 12, 6) {real, imag} */,
  {32'h3eba84b7, 32'h3ecbe5c5} /* (9, 12, 5) {real, imag} */,
  {32'h3ed29958, 32'h3dfa9a4f} /* (9, 12, 4) {real, imag} */,
  {32'hbf21b6f6, 32'hbe8abe67} /* (9, 12, 3) {real, imag} */,
  {32'h3e9092e7, 32'hbe26c0a6} /* (9, 12, 2) {real, imag} */,
  {32'h3d560cd4, 32'hbf031d6e} /* (9, 12, 1) {real, imag} */,
  {32'h3d83d0ff, 32'h3ea24e9a} /* (9, 12, 0) {real, imag} */,
  {32'hbf2247c5, 32'hbee88766} /* (9, 11, 31) {real, imag} */,
  {32'h3dfdf1b8, 32'h3e0735ab} /* (9, 11, 30) {real, imag} */,
  {32'hbc821080, 32'h3f182141} /* (9, 11, 29) {real, imag} */,
  {32'h3ea1d3e2, 32'hbef8e4d4} /* (9, 11, 28) {real, imag} */,
  {32'h3edc0d49, 32'h3e4795b8} /* (9, 11, 27) {real, imag} */,
  {32'hbe17c05a, 32'hbd281e30} /* (9, 11, 26) {real, imag} */,
  {32'hbe5d9477, 32'hbe2a72a6} /* (9, 11, 25) {real, imag} */,
  {32'h3e7c2b0e, 32'h3ec49334} /* (9, 11, 24) {real, imag} */,
  {32'h3ccb4390, 32'hbe19fbe2} /* (9, 11, 23) {real, imag} */,
  {32'hbd025360, 32'h3f107dd4} /* (9, 11, 22) {real, imag} */,
  {32'h3eaf3a78, 32'h3ef2a8d5} /* (9, 11, 21) {real, imag} */,
  {32'hbe8f9c8c, 32'hbeb2e161} /* (9, 11, 20) {real, imag} */,
  {32'hbf181146, 32'h3e1d84ed} /* (9, 11, 19) {real, imag} */,
  {32'h3cbe5aa0, 32'hbdfab20c} /* (9, 11, 18) {real, imag} */,
  {32'hbec9ee60, 32'hbd1f090b} /* (9, 11, 17) {real, imag} */,
  {32'h3e4f5b26, 32'h3e983972} /* (9, 11, 16) {real, imag} */,
  {32'h3ddd8ca2, 32'h3e671420} /* (9, 11, 15) {real, imag} */,
  {32'h3bd86c00, 32'hbf70445d} /* (9, 11, 14) {real, imag} */,
  {32'h3e445724, 32'hbf05862d} /* (9, 11, 13) {real, imag} */,
  {32'h3cc9d8f8, 32'hbe4ad478} /* (9, 11, 12) {real, imag} */,
  {32'hbe9f4117, 32'h3eecdde4} /* (9, 11, 11) {real, imag} */,
  {32'hbe5c36e2, 32'h3db7dd8a} /* (9, 11, 10) {real, imag} */,
  {32'hbe976cb5, 32'h3d55a670} /* (9, 11, 9) {real, imag} */,
  {32'h3c60aec0, 32'h3eb6c532} /* (9, 11, 8) {real, imag} */,
  {32'hbe271438, 32'h3e02fca2} /* (9, 11, 7) {real, imag} */,
  {32'h3e3d3c41, 32'hbe6499dd} /* (9, 11, 6) {real, imag} */,
  {32'h3d5b916c, 32'h3e2c8542} /* (9, 11, 5) {real, imag} */,
  {32'hbf12aa7e, 32'hbe4c5c3a} /* (9, 11, 4) {real, imag} */,
  {32'h3ea8dac4, 32'h3ec34522} /* (9, 11, 3) {real, imag} */,
  {32'h3de3d485, 32'hbd2d276c} /* (9, 11, 2) {real, imag} */,
  {32'hbe657d9a, 32'hbef29ca6} /* (9, 11, 1) {real, imag} */,
  {32'hbf3e043d, 32'hbe0cd588} /* (9, 11, 0) {real, imag} */,
  {32'h3f10603d, 32'hbea02b35} /* (9, 10, 31) {real, imag} */,
  {32'h3d36182e, 32'hbe63a9f0} /* (9, 10, 30) {real, imag} */,
  {32'hbd63c370, 32'h3eb02d04} /* (9, 10, 29) {real, imag} */,
  {32'hbea74539, 32'hbe351160} /* (9, 10, 28) {real, imag} */,
  {32'hbe00da64, 32'hbd170de8} /* (9, 10, 27) {real, imag} */,
  {32'h3e838eeb, 32'hbdc69cf6} /* (9, 10, 26) {real, imag} */,
  {32'hbe953db3, 32'h3dd09d0e} /* (9, 10, 25) {real, imag} */,
  {32'h3e7fa908, 32'h3da4b358} /* (9, 10, 24) {real, imag} */,
  {32'hbce2ec48, 32'hbeb6caa0} /* (9, 10, 23) {real, imag} */,
  {32'h3e4f4308, 32'hbea37fa5} /* (9, 10, 22) {real, imag} */,
  {32'h3ee16c4a, 32'h3e17a936} /* (9, 10, 21) {real, imag} */,
  {32'hbce15188, 32'h3ec1fef4} /* (9, 10, 20) {real, imag} */,
  {32'hbf2496b2, 32'hbe14d05a} /* (9, 10, 19) {real, imag} */,
  {32'hbf0de962, 32'hbe8427ab} /* (9, 10, 18) {real, imag} */,
  {32'h3ca8b8bc, 32'hbe779e3b} /* (9, 10, 17) {real, imag} */,
  {32'hbe379a71, 32'hbca849d0} /* (9, 10, 16) {real, imag} */,
  {32'hbd86e7d6, 32'hbe1eccc1} /* (9, 10, 15) {real, imag} */,
  {32'h3f3400d4, 32'h3f09e9f0} /* (9, 10, 14) {real, imag} */,
  {32'hbea58c60, 32'hbefed0e6} /* (9, 10, 13) {real, imag} */,
  {32'hbe32f56f, 32'hbd904ae2} /* (9, 10, 12) {real, imag} */,
  {32'h3e500520, 32'hbe8d35cc} /* (9, 10, 11) {real, imag} */,
  {32'hbf4f2a5b, 32'h3c4ae300} /* (9, 10, 10) {real, imag} */,
  {32'h3c8a3250, 32'hbf131044} /* (9, 10, 9) {real, imag} */,
  {32'h3e9bd2ab, 32'h3e4b51fd} /* (9, 10, 8) {real, imag} */,
  {32'h3eeec109, 32'hbf0b2f41} /* (9, 10, 7) {real, imag} */,
  {32'h3df40717, 32'h3bd282e0} /* (9, 10, 6) {real, imag} */,
  {32'hbe94ceee, 32'hbece3614} /* (9, 10, 5) {real, imag} */,
  {32'hbedfd0b2, 32'h3cfc0638} /* (9, 10, 4) {real, imag} */,
  {32'h3f0c27ef, 32'hbc5b2690} /* (9, 10, 3) {real, imag} */,
  {32'h3da215a1, 32'h3d15223e} /* (9, 10, 2) {real, imag} */,
  {32'h3ea33d98, 32'h3ef32f6d} /* (9, 10, 1) {real, imag} */,
  {32'hbf1d7a93, 32'h3e42dd4d} /* (9, 10, 0) {real, imag} */,
  {32'hbe90f302, 32'h3f0b683c} /* (9, 9, 31) {real, imag} */,
  {32'hbe7d5536, 32'hbf301132} /* (9, 9, 30) {real, imag} */,
  {32'h3eb408a2, 32'h3e6a9ccc} /* (9, 9, 29) {real, imag} */,
  {32'hbe0fa26c, 32'h3d8d6e22} /* (9, 9, 28) {real, imag} */,
  {32'hbdf21c05, 32'h3ec97cd5} /* (9, 9, 27) {real, imag} */,
  {32'hbe08eafd, 32'hbd78cb20} /* (9, 9, 26) {real, imag} */,
  {32'h3e6a2840, 32'hbd93f88f} /* (9, 9, 25) {real, imag} */,
  {32'hbebae645, 32'hbe8b0e76} /* (9, 9, 24) {real, imag} */,
  {32'h3dcaad82, 32'hbe4de7fe} /* (9, 9, 23) {real, imag} */,
  {32'h3e263dcc, 32'hbeb4c2ee} /* (9, 9, 22) {real, imag} */,
  {32'hbebf1268, 32'hbdee6bd5} /* (9, 9, 21) {real, imag} */,
  {32'hbdcdde10, 32'h3d958a28} /* (9, 9, 20) {real, imag} */,
  {32'hbf0e3a41, 32'h3f3287f4} /* (9, 9, 19) {real, imag} */,
  {32'h3e5511a0, 32'h3cc0d170} /* (9, 9, 18) {real, imag} */,
  {32'hbd3aa008, 32'h3e422151} /* (9, 9, 17) {real, imag} */,
  {32'h3ead974e, 32'h3d4ffaca} /* (9, 9, 16) {real, imag} */,
  {32'h3de513d3, 32'hbec68d6e} /* (9, 9, 15) {real, imag} */,
  {32'h3d6ab22c, 32'h3d047d0a} /* (9, 9, 14) {real, imag} */,
  {32'hbe78d97a, 32'h3eb91768} /* (9, 9, 13) {real, imag} */,
  {32'hbeb6e39d, 32'h3d0e6c98} /* (9, 9, 12) {real, imag} */,
  {32'hbcf69a34, 32'hbe93a178} /* (9, 9, 11) {real, imag} */,
  {32'h3f4839b3, 32'h3ea276db} /* (9, 9, 10) {real, imag} */,
  {32'hbeab39a1, 32'hbdcf7b6e} /* (9, 9, 9) {real, imag} */,
  {32'h3ebfc2e9, 32'hbf0a8aa8} /* (9, 9, 8) {real, imag} */,
  {32'hbe6bc9de, 32'h3f0f8dec} /* (9, 9, 7) {real, imag} */,
  {32'hbe95a206, 32'h3ec027aa} /* (9, 9, 6) {real, imag} */,
  {32'hbf148df5, 32'hbdbc8e90} /* (9, 9, 5) {real, imag} */,
  {32'hbf139144, 32'h3ec81848} /* (9, 9, 4) {real, imag} */,
  {32'h3ea90906, 32'h3ebff948} /* (9, 9, 3) {real, imag} */,
  {32'h3ee8f3cc, 32'hbebb5eb7} /* (9, 9, 2) {real, imag} */,
  {32'h3f51964f, 32'hbe87fbde} /* (9, 9, 1) {real, imag} */,
  {32'h3e881a94, 32'hbf020bc7} /* (9, 9, 0) {real, imag} */,
  {32'hbfab9308, 32'hbf321bbd} /* (9, 8, 31) {real, imag} */,
  {32'h3f79c2d7, 32'h3e95260e} /* (9, 8, 30) {real, imag} */,
  {32'h3d90dde7, 32'hbee3fc8c} /* (9, 8, 29) {real, imag} */,
  {32'h3e879894, 32'h3f735b23} /* (9, 8, 28) {real, imag} */,
  {32'h3d865b38, 32'hbc9a3428} /* (9, 8, 27) {real, imag} */,
  {32'h3e1461b4, 32'hbf0e0432} /* (9, 8, 26) {real, imag} */,
  {32'h3e515f48, 32'hbe02ce15} /* (9, 8, 25) {real, imag} */,
  {32'hbd901b68, 32'hbeabe38c} /* (9, 8, 24) {real, imag} */,
  {32'hbf44f950, 32'hbe2151ce} /* (9, 8, 23) {real, imag} */,
  {32'hbe85869f, 32'h3e9d33b8} /* (9, 8, 22) {real, imag} */,
  {32'hbdef0b20, 32'h3eeaf8cc} /* (9, 8, 21) {real, imag} */,
  {32'h3cf6592c, 32'hbde38db1} /* (9, 8, 20) {real, imag} */,
  {32'hbcd575a0, 32'h3e1d2aef} /* (9, 8, 19) {real, imag} */,
  {32'h3e343d0d, 32'h3e71d7cb} /* (9, 8, 18) {real, imag} */,
  {32'hbe9cf51d, 32'hbf07981c} /* (9, 8, 17) {real, imag} */,
  {32'h3ea84177, 32'h3d88d2f0} /* (9, 8, 16) {real, imag} */,
  {32'hbe855741, 32'h3b3de780} /* (9, 8, 15) {real, imag} */,
  {32'hbe360709, 32'h3eb0e052} /* (9, 8, 14) {real, imag} */,
  {32'h3d8e1b4c, 32'hbe531e45} /* (9, 8, 13) {real, imag} */,
  {32'hbec2ac24, 32'hbd94dad1} /* (9, 8, 12) {real, imag} */,
  {32'hbe2638de, 32'hbdc91660} /* (9, 8, 11) {real, imag} */,
  {32'hbe4d28c2, 32'h3ded0bb8} /* (9, 8, 10) {real, imag} */,
  {32'h3dd726ba, 32'h3eb8668b} /* (9, 8, 9) {real, imag} */,
  {32'hbed6b7f6, 32'h3f13374b} /* (9, 8, 8) {real, imag} */,
  {32'h3ee87c3a, 32'h3f87439c} /* (9, 8, 7) {real, imag} */,
  {32'hbe335e82, 32'h3d1467ec} /* (9, 8, 6) {real, imag} */,
  {32'h3f21bb48, 32'hbdaa1284} /* (9, 8, 5) {real, imag} */,
  {32'h3e659cee, 32'h3de04ecc} /* (9, 8, 4) {real, imag} */,
  {32'hbcb4bb00, 32'h3eb7909a} /* (9, 8, 3) {real, imag} */,
  {32'h3e5b9691, 32'hbea6c05a} /* (9, 8, 2) {real, imag} */,
  {32'hbe409db9, 32'hbf0e2ef2} /* (9, 8, 1) {real, imag} */,
  {32'hbf8b388c, 32'hbec1f294} /* (9, 8, 0) {real, imag} */,
  {32'h3f0d0f0b, 32'h3ec206ed} /* (9, 7, 31) {real, imag} */,
  {32'h3cb320f0, 32'hbf456090} /* (9, 7, 30) {real, imag} */,
  {32'hbe80d1fe, 32'h3e808979} /* (9, 7, 29) {real, imag} */,
  {32'hbe85b476, 32'hbe5cacf0} /* (9, 7, 28) {real, imag} */,
  {32'hbf264e32, 32'h3e9998ba} /* (9, 7, 27) {real, imag} */,
  {32'hbd9429f6, 32'h3d8b1ec8} /* (9, 7, 26) {real, imag} */,
  {32'hbe15c019, 32'hbeda9bc7} /* (9, 7, 25) {real, imag} */,
  {32'hbd203af8, 32'hbf29dd94} /* (9, 7, 24) {real, imag} */,
  {32'hbf3f03b2, 32'hbda4b61c} /* (9, 7, 23) {real, imag} */,
  {32'h3e0fe90a, 32'h3eb4339a} /* (9, 7, 22) {real, imag} */,
  {32'hbe8f11e6, 32'hbde9ed31} /* (9, 7, 21) {real, imag} */,
  {32'h3e6fbfe4, 32'h3eb56422} /* (9, 7, 20) {real, imag} */,
  {32'h3eb20fea, 32'h3ea917ba} /* (9, 7, 19) {real, imag} */,
  {32'h3da5c396, 32'hbe6a10f6} /* (9, 7, 18) {real, imag} */,
  {32'h3eaeb7af, 32'h3d8ed740} /* (9, 7, 17) {real, imag} */,
  {32'hbd90a314, 32'hbdb4c2ca} /* (9, 7, 16) {real, imag} */,
  {32'hbec4446e, 32'h3e0ac34c} /* (9, 7, 15) {real, imag} */,
  {32'hbf0d5daf, 32'h3da7a090} /* (9, 7, 14) {real, imag} */,
  {32'h3e51304a, 32'hbf2a97e8} /* (9, 7, 13) {real, imag} */,
  {32'hbe8702ef, 32'h3d1d1b9a} /* (9, 7, 12) {real, imag} */,
  {32'h3e4e1327, 32'h3e18c76a} /* (9, 7, 11) {real, imag} */,
  {32'h3ea78658, 32'hbe651bba} /* (9, 7, 10) {real, imag} */,
  {32'h3e7d5ab0, 32'h3f0c4f5b} /* (9, 7, 9) {real, imag} */,
  {32'hbeb37814, 32'h3e3b3a40} /* (9, 7, 8) {real, imag} */,
  {32'h3e7c3dca, 32'hbeb65872} /* (9, 7, 7) {real, imag} */,
  {32'h3ce893f0, 32'hbe9cf9f4} /* (9, 7, 6) {real, imag} */,
  {32'h3f2e0abc, 32'h3e01ccb5} /* (9, 7, 5) {real, imag} */,
  {32'h3da6d8df, 32'h3e980da2} /* (9, 7, 4) {real, imag} */,
  {32'hbd7318cc, 32'h3e24c9dc} /* (9, 7, 3) {real, imag} */,
  {32'hbe954f9d, 32'hbf50af36} /* (9, 7, 2) {real, imag} */,
  {32'h3ba8d720, 32'h3f346930} /* (9, 7, 1) {real, imag} */,
  {32'hbe13b8dd, 32'h3e392cb6} /* (9, 7, 0) {real, imag} */,
  {32'h3d906338, 32'h3eec182d} /* (9, 6, 31) {real, imag} */,
  {32'h3e8c098d, 32'h3e25c617} /* (9, 6, 30) {real, imag} */,
  {32'hba710200, 32'h3edc52b8} /* (9, 6, 29) {real, imag} */,
  {32'h3f39c2ba, 32'hbf2820c9} /* (9, 6, 28) {real, imag} */,
  {32'hbe2df51d, 32'hbdff1a2c} /* (9, 6, 27) {real, imag} */,
  {32'h3f31d271, 32'h3f278c22} /* (9, 6, 26) {real, imag} */,
  {32'hbea1ca64, 32'h3d1de6e6} /* (9, 6, 25) {real, imag} */,
  {32'hbe118b75, 32'h3dc1bd62} /* (9, 6, 24) {real, imag} */,
  {32'h3e495adb, 32'h3ebdbd84} /* (9, 6, 23) {real, imag} */,
  {32'h3e595fcf, 32'hbec2d8b2} /* (9, 6, 22) {real, imag} */,
  {32'h3e83c4a6, 32'h3e946f09} /* (9, 6, 21) {real, imag} */,
  {32'h3cbc3738, 32'h3de2e628} /* (9, 6, 20) {real, imag} */,
  {32'h3e57ff22, 32'hbe8faeaa} /* (9, 6, 19) {real, imag} */,
  {32'h3dce8858, 32'h3ea47d7c} /* (9, 6, 18) {real, imag} */,
  {32'hbe3c3bb4, 32'h3e73f20d} /* (9, 6, 17) {real, imag} */,
  {32'hbea97b59, 32'hbd971e7e} /* (9, 6, 16) {real, imag} */,
  {32'h3e9278fa, 32'h3e08cb0a} /* (9, 6, 15) {real, imag} */,
  {32'hbe1861d8, 32'hbe231c67} /* (9, 6, 14) {real, imag} */,
  {32'hbc460770, 32'h3d7850f4} /* (9, 6, 13) {real, imag} */,
  {32'hbf02cfed, 32'h3ec014dc} /* (9, 6, 12) {real, imag} */,
  {32'h3edff534, 32'h3f31599c} /* (9, 6, 11) {real, imag} */,
  {32'hbdd745cc, 32'h3f296a98} /* (9, 6, 10) {real, imag} */,
  {32'hbd68a5fc, 32'h3de432de} /* (9, 6, 9) {real, imag} */,
  {32'h3e5d23a8, 32'hbea34e5d} /* (9, 6, 8) {real, imag} */,
  {32'h3e42633a, 32'h3e302450} /* (9, 6, 7) {real, imag} */,
  {32'h3ed6bd63, 32'h3e806a9d} /* (9, 6, 6) {real, imag} */,
  {32'h3e67392e, 32'hbbd6fd80} /* (9, 6, 5) {real, imag} */,
  {32'h3eb292da, 32'hbd410dc0} /* (9, 6, 4) {real, imag} */,
  {32'hbe607254, 32'hbe4d7805} /* (9, 6, 3) {real, imag} */,
  {32'hbf5ffff6, 32'hbf40c6d2} /* (9, 6, 2) {real, imag} */,
  {32'h3ea90938, 32'h3e9a57f6} /* (9, 6, 1) {real, imag} */,
  {32'h3d9f004c, 32'h3f1194ac} /* (9, 6, 0) {real, imag} */,
  {32'hc051ec08, 32'hbe01e296} /* (9, 5, 31) {real, imag} */,
  {32'h3f048bb4, 32'hbe87af27} /* (9, 5, 30) {real, imag} */,
  {32'h3f1c6dff, 32'h3ec5efd5} /* (9, 5, 29) {real, imag} */,
  {32'hbe85b0bb, 32'h3d3b7200} /* (9, 5, 28) {real, imag} */,
  {32'hbdfb17c8, 32'h3e909960} /* (9, 5, 27) {real, imag} */,
  {32'h3eac16aa, 32'h3f438d36} /* (9, 5, 26) {real, imag} */,
  {32'hbe2c7bdc, 32'h3f211e4b} /* (9, 5, 25) {real, imag} */,
  {32'h3ebd15c2, 32'hbd889c91} /* (9, 5, 24) {real, imag} */,
  {32'h3e9501cb, 32'h3cbaa684} /* (9, 5, 23) {real, imag} */,
  {32'hbf33b325, 32'hbbcd0100} /* (9, 5, 22) {real, imag} */,
  {32'h3eab022b, 32'h3d8c35a6} /* (9, 5, 21) {real, imag} */,
  {32'hbe9141a3, 32'hbdf477c2} /* (9, 5, 20) {real, imag} */,
  {32'hbedefd1a, 32'h3ea8249b} /* (9, 5, 19) {real, imag} */,
  {32'h3d59e90c, 32'hbd87e700} /* (9, 5, 18) {real, imag} */,
  {32'hbde7b16a, 32'h3e6ed38f} /* (9, 5, 17) {real, imag} */,
  {32'h3ebdd0d8, 32'h3c3d9e50} /* (9, 5, 16) {real, imag} */,
  {32'h3e526ddc, 32'h3c6436b4} /* (9, 5, 15) {real, imag} */,
  {32'h3e9496c4, 32'hbcdce59c} /* (9, 5, 14) {real, imag} */,
  {32'hbda84551, 32'h3d754bd0} /* (9, 5, 13) {real, imag} */,
  {32'hbd1b9978, 32'h3d22a30f} /* (9, 5, 12) {real, imag} */,
  {32'hbd8cb252, 32'h3f0f4ff0} /* (9, 5, 11) {real, imag} */,
  {32'h3d8fa0ac, 32'h3f681e0d} /* (9, 5, 10) {real, imag} */,
  {32'h3e2298c5, 32'hbe441566} /* (9, 5, 9) {real, imag} */,
  {32'hbb803680, 32'hbd49e728} /* (9, 5, 8) {real, imag} */,
  {32'hbe032666, 32'hbeec7b3a} /* (9, 5, 7) {real, imag} */,
  {32'hbe1e2312, 32'h3eab7902} /* (9, 5, 6) {real, imag} */,
  {32'h3f9b9724, 32'h3ebd4d47} /* (9, 5, 5) {real, imag} */,
  {32'hbeb0a827, 32'hbe1f1190} /* (9, 5, 4) {real, imag} */,
  {32'hbf6dfd25, 32'hbec1ee4b} /* (9, 5, 3) {real, imag} */,
  {32'h3f7aff09, 32'h3f9ee39a} /* (9, 5, 2) {real, imag} */,
  {32'hbf8e53da, 32'hc0183dde} /* (9, 5, 1) {real, imag} */,
  {32'hbfd9bfcc, 32'hbf6fe0a2} /* (9, 5, 0) {real, imag} */,
  {32'h3f3382f6, 32'h404c40c4} /* (9, 4, 31) {real, imag} */,
  {32'hc03b769c, 32'hc018c6ae} /* (9, 4, 30) {real, imag} */,
  {32'hbed35150, 32'hbe9a7a75} /* (9, 4, 29) {real, imag} */,
  {32'h3f83af83, 32'h3e37006e} /* (9, 4, 28) {real, imag} */,
  {32'hbf2f5c3e, 32'hbf3e297f} /* (9, 4, 27) {real, imag} */,
  {32'hbedd4d0a, 32'h3ea8cd71} /* (9, 4, 26) {real, imag} */,
  {32'h3ddb1766, 32'h3f0c45ad} /* (9, 4, 25) {real, imag} */,
  {32'h3e016374, 32'hbec259ce} /* (9, 4, 24) {real, imag} */,
  {32'h3ee5f52a, 32'hbd8ffaf8} /* (9, 4, 23) {real, imag} */,
  {32'hbe5f5969, 32'hbe0ba6f6} /* (9, 4, 22) {real, imag} */,
  {32'hbda38ece, 32'h3f32aba0} /* (9, 4, 21) {real, imag} */,
  {32'h3ef4b962, 32'hbd912bfa} /* (9, 4, 20) {real, imag} */,
  {32'hbedf7d20, 32'hbf024abc} /* (9, 4, 19) {real, imag} */,
  {32'hbe87a3f4, 32'hbd9d2ee4} /* (9, 4, 18) {real, imag} */,
  {32'h3e98a53c, 32'hbe21dc22} /* (9, 4, 17) {real, imag} */,
  {32'hbe47b2e5, 32'h3d5ba0e2} /* (9, 4, 16) {real, imag} */,
  {32'h3e22a01a, 32'h3e00f911} /* (9, 4, 15) {real, imag} */,
  {32'h3d2d2042, 32'hbe3dc6a5} /* (9, 4, 14) {real, imag} */,
  {32'hbe0c0e3e, 32'hbe2fb75a} /* (9, 4, 13) {real, imag} */,
  {32'hbf5897d5, 32'h3e8eb4ec} /* (9, 4, 12) {real, imag} */,
  {32'h3e5a790f, 32'hbead6fdd} /* (9, 4, 11) {real, imag} */,
  {32'h3e9ae7a4, 32'h3e0fb2c9} /* (9, 4, 10) {real, imag} */,
  {32'h3e325510, 32'hbe0f40c4} /* (9, 4, 9) {real, imag} */,
  {32'hbe95bbe0, 32'hbe9c68a3} /* (9, 4, 8) {real, imag} */,
  {32'hbd5eb5e0, 32'hbeffa0e4} /* (9, 4, 7) {real, imag} */,
  {32'h3f3d1858, 32'hbd9e1364} /* (9, 4, 6) {real, imag} */,
  {32'hbe500e40, 32'hbf5059f2} /* (9, 4, 5) {real, imag} */,
  {32'h3eeaa38e, 32'h3f1dab8d} /* (9, 4, 4) {real, imag} */,
  {32'hbf9c4e87, 32'h3fd32e9c} /* (9, 4, 3) {real, imag} */,
  {32'hbfc694f6, 32'hc0288ca7} /* (9, 4, 2) {real, imag} */,
  {32'h408dff05, 32'h3f894c94} /* (9, 4, 1) {real, imag} */,
  {32'h3f94a618, 32'h3f419450} /* (9, 4, 0) {real, imag} */,
  {32'hc07eea4c, 32'h3fa78557} /* (9, 3, 31) {real, imag} */,
  {32'h400a0160, 32'hc0aa8cc7} /* (9, 3, 30) {real, imag} */,
  {32'h3d5336b4, 32'h3f6b199d} /* (9, 3, 29) {real, imag} */,
  {32'h3f6f50c3, 32'h3e01faa6} /* (9, 3, 28) {real, imag} */,
  {32'hbfa4ce6e, 32'hbeba1917} /* (9, 3, 27) {real, imag} */,
  {32'h3d14d3d8, 32'h3eda4ed6} /* (9, 3, 26) {real, imag} */,
  {32'hbf122f2b, 32'hbe42ea38} /* (9, 3, 25) {real, imag} */,
  {32'h3f0ce24b, 32'hbf10014e} /* (9, 3, 24) {real, imag} */,
  {32'hbe5acbc2, 32'h3e8e4e75} /* (9, 3, 23) {real, imag} */,
  {32'hbebfc771, 32'h3cd43014} /* (9, 3, 22) {real, imag} */,
  {32'hbe1bd94e, 32'hbeb5716c} /* (9, 3, 21) {real, imag} */,
  {32'h3e35d577, 32'h3dbea28a} /* (9, 3, 20) {real, imag} */,
  {32'h3eaac4d1, 32'hbd868634} /* (9, 3, 19) {real, imag} */,
  {32'h3e99840e, 32'h3e1a57d2} /* (9, 3, 18) {real, imag} */,
  {32'h3e298de0, 32'hbebcb9e8} /* (9, 3, 17) {real, imag} */,
  {32'h3dcf2860, 32'hbe4c41ff} /* (9, 3, 16) {real, imag} */,
  {32'h3e9df930, 32'h3e896487} /* (9, 3, 15) {real, imag} */,
  {32'hbe2f22ad, 32'h3e34f981} /* (9, 3, 14) {real, imag} */,
  {32'hbdcb693a, 32'h3e6ca620} /* (9, 3, 13) {real, imag} */,
  {32'h3ee01a8e, 32'h3e50f065} /* (9, 3, 12) {real, imag} */,
  {32'hbdc5076c, 32'hbd165254} /* (9, 3, 11) {real, imag} */,
  {32'hbebcffc4, 32'h3ed62576} /* (9, 3, 10) {real, imag} */,
  {32'hbb6c5a10, 32'h3e40f446} /* (9, 3, 9) {real, imag} */,
  {32'hbf4b02f4, 32'h3ea48d92} /* (9, 3, 8) {real, imag} */,
  {32'hbe83746e, 32'hbe377d52} /* (9, 3, 7) {real, imag} */,
  {32'hbc92e8c0, 32'h3f28b76b} /* (9, 3, 6) {real, imag} */,
  {32'hbe59758c, 32'h3df82040} /* (9, 3, 5) {real, imag} */,
  {32'hbfa221b2, 32'h3dfff548} /* (9, 3, 4) {real, imag} */,
  {32'hbf7177e0, 32'h3e88571a} /* (9, 3, 3) {real, imag} */,
  {32'hbcd755c0, 32'hc04a9267} /* (9, 3, 2) {real, imag} */,
  {32'h40452f9a, 32'h405115a2} /* (9, 3, 1) {real, imag} */,
  {32'hbea0eb90, 32'hbf6257cc} /* (9, 3, 0) {real, imag} */,
  {32'hc222fd64, 32'hbfc2606e} /* (9, 2, 31) {real, imag} */,
  {32'h418f54ac, 32'hc0b538f6} /* (9, 2, 30) {real, imag} */,
  {32'h3f1a4284, 32'h3fb0401d} /* (9, 2, 29) {real, imag} */,
  {32'hbf06c26b, 32'h4012eebb} /* (9, 2, 28) {real, imag} */,
  {32'h402bba8f, 32'hbf8fb289} /* (9, 2, 27) {real, imag} */,
  {32'h3ed40f24, 32'hbf1890a7} /* (9, 2, 26) {real, imag} */,
  {32'hbe99d8cb, 32'hbe4b52c9} /* (9, 2, 25) {real, imag} */,
  {32'h3f6ffc58, 32'hbf16d7ef} /* (9, 2, 24) {real, imag} */,
  {32'h3eb5e4b7, 32'h3f10bdaf} /* (9, 2, 23) {real, imag} */,
  {32'h3d038d64, 32'h3de19436} /* (9, 2, 22) {real, imag} */,
  {32'hbe7b4764, 32'h3a4078c0} /* (9, 2, 21) {real, imag} */,
  {32'hbdbb6334, 32'h3e2abf42} /* (9, 2, 20) {real, imag} */,
  {32'h3e426e5c, 32'hbe137cb0} /* (9, 2, 19) {real, imag} */,
  {32'hbd77cdf2, 32'hbf63eb3d} /* (9, 2, 18) {real, imag} */,
  {32'hbe130a8a, 32'h3d47aecc} /* (9, 2, 17) {real, imag} */,
  {32'h3e5eddd0, 32'hbe1b5aa5} /* (9, 2, 16) {real, imag} */,
  {32'hbdba2220, 32'hbeac8000} /* (9, 2, 15) {real, imag} */,
  {32'hbdaec384, 32'h3e32e074} /* (9, 2, 14) {real, imag} */,
  {32'h3dc7ec5c, 32'hbc9b9480} /* (9, 2, 13) {real, imag} */,
  {32'h3e9d3200, 32'hbe3ca626} /* (9, 2, 12) {real, imag} */,
  {32'h3e8e2894, 32'h3ea7577c} /* (9, 2, 11) {real, imag} */,
  {32'hbeffd13e, 32'hbec70152} /* (9, 2, 10) {real, imag} */,
  {32'h3e9d899e, 32'h3eb4fd31} /* (9, 2, 9) {real, imag} */,
  {32'h3f10afbf, 32'h3e9f2e7b} /* (9, 2, 8) {real, imag} */,
  {32'hbf5f366c, 32'hbd0f0c70} /* (9, 2, 7) {real, imag} */,
  {32'h3f02dcee, 32'hbeb37d9d} /* (9, 2, 6) {real, imag} */,
  {32'h3fb90c3a, 32'h3fb1fd35} /* (9, 2, 5) {real, imag} */,
  {32'hc038aad1, 32'hbfcab37a} /* (9, 2, 4) {real, imag} */,
  {32'hbf0dac46, 32'h3eaf5658} /* (9, 2, 3) {real, imag} */,
  {32'h4158527b, 32'hc06c34d2} /* (9, 2, 2) {real, imag} */,
  {32'hc1b2a101, 32'h40c46f42} /* (9, 2, 1) {real, imag} */,
  {32'hc1aff663, 32'hc080b112} /* (9, 2, 0) {real, imag} */,
  {32'h4252283a, 32'hc153f00b} /* (9, 1, 31) {real, imag} */,
  {32'hc13bee4a, 32'h400e708b} /* (9, 1, 30) {real, imag} */,
  {32'hbfb36371, 32'hbf22051b} /* (9, 1, 29) {real, imag} */,
  {32'h401d877b, 32'h4040738a} /* (9, 1, 28) {real, imag} */,
  {32'hc0295a45, 32'hbf5c97f4} /* (9, 1, 27) {real, imag} */,
  {32'hbf208e7c, 32'hbeb89bdc} /* (9, 1, 26) {real, imag} */,
  {32'h3f967626, 32'hbf3868f7} /* (9, 1, 25) {real, imag} */,
  {32'hbf69ef22, 32'h3df1dc1c} /* (9, 1, 24) {real, imag} */,
  {32'h3ecaca9c, 32'h3ca45c50} /* (9, 1, 23) {real, imag} */,
  {32'hbddacc0c, 32'h3e2adedc} /* (9, 1, 22) {real, imag} */,
  {32'hbf5d6582, 32'h3eb4f38a} /* (9, 1, 21) {real, imag} */,
  {32'h3ea4890c, 32'h3e8d52f6} /* (9, 1, 20) {real, imag} */,
  {32'h3e098cc8, 32'hbea3a916} /* (9, 1, 19) {real, imag} */,
  {32'hbf030a4a, 32'h3f443cca} /* (9, 1, 18) {real, imag} */,
  {32'h3c161ec4, 32'h3d40c49c} /* (9, 1, 17) {real, imag} */,
  {32'hbd90715f, 32'h3e7c766a} /* (9, 1, 16) {real, imag} */,
  {32'hbedaedf0, 32'h3e0217d0} /* (9, 1, 15) {real, imag} */,
  {32'h3ddad65a, 32'hbe90be98} /* (9, 1, 14) {real, imag} */,
  {32'h3ec8b3bf, 32'hbce36a60} /* (9, 1, 13) {real, imag} */,
  {32'h3e7cdd38, 32'hbf0a3c1d} /* (9, 1, 12) {real, imag} */,
  {32'h3dcec3a4, 32'hbf240c9a} /* (9, 1, 11) {real, imag} */,
  {32'hbf26cade, 32'hbef3b006} /* (9, 1, 10) {real, imag} */,
  {32'h3c465ae0, 32'h3eb77dbe} /* (9, 1, 9) {real, imag} */,
  {32'hbe92a991, 32'hbf5873d2} /* (9, 1, 8) {real, imag} */,
  {32'h3f07fa93, 32'hbe3fd081} /* (9, 1, 7) {real, imag} */,
  {32'hbf9272ca, 32'hbedbcfb1} /* (9, 1, 6) {real, imag} */,
  {32'hc0388f86, 32'hbf35d8cf} /* (9, 1, 5) {real, imag} */,
  {32'h400c7824, 32'h3ea10898} /* (9, 1, 4) {real, imag} */,
  {32'hbef75210, 32'h3eededac} /* (9, 1, 3) {real, imag} */,
  {32'hc19b750a, 32'hc18b2cf5} /* (9, 1, 2) {real, imag} */,
  {32'h4299b1b4, 32'h42209d10} /* (9, 1, 1) {real, imag} */,
  {32'h42905eca, 32'h40dc289a} /* (9, 1, 0) {real, imag} */,
  {32'h42318a4e, 32'hc2102210} /* (9, 0, 31) {real, imag} */,
  {32'hc0bae13a, 32'h413c3442} /* (9, 0, 30) {real, imag} */,
  {32'hbfd3a414, 32'h3f5cb57c} /* (9, 0, 29) {real, imag} */,
  {32'hbe8003ec, 32'h3dcd0380} /* (9, 0, 28) {real, imag} */,
  {32'hbfeb67c0, 32'hbdfd899a} /* (9, 0, 27) {real, imag} */,
  {32'h3e8a8180, 32'hbe528827} /* (9, 0, 26) {real, imag} */,
  {32'h3eae9e63, 32'h3da1af90} /* (9, 0, 25) {real, imag} */,
  {32'h3ea21586, 32'h3fb1fbf0} /* (9, 0, 24) {real, imag} */,
  {32'hbc8879f0, 32'hbedca9bf} /* (9, 0, 23) {real, imag} */,
  {32'h3ecc5986, 32'h3f1ee578} /* (9, 0, 22) {real, imag} */,
  {32'hbee18145, 32'hbed22b5c} /* (9, 0, 21) {real, imag} */,
  {32'h3e48c07d, 32'hbdde21d0} /* (9, 0, 20) {real, imag} */,
  {32'h3e8e02ac, 32'hbeebe810} /* (9, 0, 19) {real, imag} */,
  {32'h3c86d4b4, 32'h3ed2962c} /* (9, 0, 18) {real, imag} */,
  {32'hbeca8a4a, 32'hbdf70406} /* (9, 0, 17) {real, imag} */,
  {32'h3e41a47e, 32'h00000000} /* (9, 0, 16) {real, imag} */,
  {32'hbeca8a4a, 32'h3df70406} /* (9, 0, 15) {real, imag} */,
  {32'h3c86d4b4, 32'hbed2962c} /* (9, 0, 14) {real, imag} */,
  {32'h3e8e02ac, 32'h3eebe810} /* (9, 0, 13) {real, imag} */,
  {32'h3e48c07d, 32'h3dde21d0} /* (9, 0, 12) {real, imag} */,
  {32'hbee18145, 32'h3ed22b5c} /* (9, 0, 11) {real, imag} */,
  {32'h3ecc5986, 32'hbf1ee578} /* (9, 0, 10) {real, imag} */,
  {32'hbc8879f0, 32'h3edca9bf} /* (9, 0, 9) {real, imag} */,
  {32'h3ea21586, 32'hbfb1fbf0} /* (9, 0, 8) {real, imag} */,
  {32'h3eae9e63, 32'hbda1af90} /* (9, 0, 7) {real, imag} */,
  {32'h3e8a8180, 32'h3e528827} /* (9, 0, 6) {real, imag} */,
  {32'hbfeb67c0, 32'h3dfd899a} /* (9, 0, 5) {real, imag} */,
  {32'hbe8003ec, 32'hbdcd0380} /* (9, 0, 4) {real, imag} */,
  {32'hbfd3a414, 32'hbf5cb57c} /* (9, 0, 3) {real, imag} */,
  {32'hc0bae13a, 32'hc13c3442} /* (9, 0, 2) {real, imag} */,
  {32'h42318a4e, 32'h42102210} /* (9, 0, 1) {real, imag} */,
  {32'h42966e52, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h428bb595, 32'hc20a3849} /* (8, 31, 31) {real, imag} */,
  {32'hc18af8a8, 32'h4181b2e0} /* (8, 31, 30) {real, imag} */,
  {32'hbf9060a1, 32'h3fc35b96} /* (8, 31, 29) {real, imag} */,
  {32'h3fe99c56, 32'h3f035cb3} /* (8, 31, 28) {real, imag} */,
  {32'hc01f7400, 32'h3f26fb00} /* (8, 31, 27) {real, imag} */,
  {32'hbf56180e, 32'h3de9fab4} /* (8, 31, 26) {real, imag} */,
  {32'h3eae5da6, 32'hbec9af36} /* (8, 31, 25) {real, imag} */,
  {32'hbd9f0128, 32'h3f699d99} /* (8, 31, 24) {real, imag} */,
  {32'hbe89eb2a, 32'h3f0b9a8a} /* (8, 31, 23) {real, imag} */,
  {32'hbf3db8a6, 32'h3e4da082} /* (8, 31, 22) {real, imag} */,
  {32'hbe914d2c, 32'h3f2ec71a} /* (8, 31, 21) {real, imag} */,
  {32'h3d3e162c, 32'h3f1ccdf0} /* (8, 31, 20) {real, imag} */,
  {32'h3de70ff6, 32'h3d0e4e50} /* (8, 31, 19) {real, imag} */,
  {32'h3e6556b2, 32'h3f0606e2} /* (8, 31, 18) {real, imag} */,
  {32'h3e07c8b9, 32'hbe9b5098} /* (8, 31, 17) {real, imag} */,
  {32'h3e1f1e63, 32'hbcf7e51e} /* (8, 31, 16) {real, imag} */,
  {32'hbd9f94a6, 32'hbcb1bf3c} /* (8, 31, 15) {real, imag} */,
  {32'hbeaa4c87, 32'hbf189ca2} /* (8, 31, 14) {real, imag} */,
  {32'hbdbc7b21, 32'h3e1ef37c} /* (8, 31, 13) {real, imag} */,
  {32'h3ece6234, 32'h3f220ee9} /* (8, 31, 12) {real, imag} */,
  {32'hbfae581e, 32'hbe49eff2} /* (8, 31, 11) {real, imag} */,
  {32'h3d8cc0b8, 32'hbe5bd85f} /* (8, 31, 10) {real, imag} */,
  {32'h3e133ae0, 32'hbedd209e} /* (8, 31, 9) {real, imag} */,
  {32'hbf91bc7d, 32'h3c224140} /* (8, 31, 8) {real, imag} */,
  {32'h3f15d823, 32'h3edcee22} /* (8, 31, 7) {real, imag} */,
  {32'hbf1807b8, 32'hbeaed425} /* (8, 31, 6) {real, imag} */,
  {32'hc035cc2c, 32'h3ea3a32d} /* (8, 31, 5) {real, imag} */,
  {32'h400394cd, 32'hc0207ef2} /* (8, 31, 4) {real, imag} */,
  {32'hbe80a106, 32'h3e7e2978} /* (8, 31, 3) {real, imag} */,
  {32'hc12b8065, 32'hc0169374} /* (8, 31, 2) {real, imag} */,
  {32'h4243e72d, 32'h4146ca94} /* (8, 31, 1) {real, imag} */,
  {32'h4284ce84, 32'hc0e653ae} /* (8, 31, 0) {real, imag} */,
  {32'hc1a03dbc, 32'hc0a12c7c} /* (8, 30, 31) {real, imag} */,
  {32'h414ce94e, 32'h402d8e00} /* (8, 30, 30) {real, imag} */,
  {32'hbf650215, 32'hbde02560} /* (8, 30, 29) {real, imag} */,
  {32'hc05758c2, 32'h3f43bede} /* (8, 30, 28) {real, imag} */,
  {32'h400c6076, 32'hbf5bbdea} /* (8, 30, 27) {real, imag} */,
  {32'h3d642078, 32'hbe60be35} /* (8, 30, 26) {real, imag} */,
  {32'hbf10a884, 32'h3f839adc} /* (8, 30, 25) {real, imag} */,
  {32'hbe0f4426, 32'hbd818f42} /* (8, 30, 24) {real, imag} */,
  {32'h3eec9750, 32'hbe619701} /* (8, 30, 23) {real, imag} */,
  {32'hbe3bccc2, 32'h3ce216b0} /* (8, 30, 22) {real, imag} */,
  {32'hbd5a6a86, 32'hbed848fc} /* (8, 30, 21) {real, imag} */,
  {32'h3ed3a7cb, 32'h3eb1c74c} /* (8, 30, 20) {real, imag} */,
  {32'h3e9e21f4, 32'h3e613645} /* (8, 30, 19) {real, imag} */,
  {32'hbe7ced45, 32'hbe875247} /* (8, 30, 18) {real, imag} */,
  {32'hbec8bf24, 32'hbe57b4b5} /* (8, 30, 17) {real, imag} */,
  {32'hbea1e42e, 32'hbe9acf0c} /* (8, 30, 16) {real, imag} */,
  {32'h3f0739ba, 32'hbe9d214c} /* (8, 30, 15) {real, imag} */,
  {32'hbe9a609b, 32'h3c283950} /* (8, 30, 14) {real, imag} */,
  {32'h3c8e9734, 32'h3eb0bbed} /* (8, 30, 13) {real, imag} */,
  {32'h3ef8535d, 32'h3f4f1b82} /* (8, 30, 12) {real, imag} */,
  {32'hbe87f4f8, 32'h3e7c9800} /* (8, 30, 11) {real, imag} */,
  {32'hbe952825, 32'h3deb0078} /* (8, 30, 10) {real, imag} */,
  {32'hbe8e917f, 32'h3d9d929a} /* (8, 30, 9) {real, imag} */,
  {32'h3f158887, 32'hba8cca00} /* (8, 30, 8) {real, imag} */,
  {32'h3f37d1e8, 32'hbefe53be} /* (8, 30, 7) {real, imag} */,
  {32'h3f26cd38, 32'h3ebf15dd} /* (8, 30, 6) {real, imag} */,
  {32'h402003a0, 32'h3f9caf60} /* (8, 30, 5) {real, imag} */,
  {32'hbf7f7fdc, 32'hc00ed330} /* (8, 30, 4) {real, imag} */,
  {32'hbf7b0fdb, 32'hc0120442} /* (8, 30, 3) {real, imag} */,
  {32'h418a3d64, 32'h4099eda6} /* (8, 30, 2) {real, imag} */,
  {32'hc218727c, 32'h3f7fb2f2} /* (8, 30, 1) {real, imag} */,
  {32'hc19b20e7, 32'h40958d32} /* (8, 30, 0) {real, imag} */,
  {32'h40635e97, 32'hc04fbbd8} /* (8, 29, 31) {real, imag} */,
  {32'h3e888d04, 32'h402fbae0} /* (8, 29, 30) {real, imag} */,
  {32'hbf1fe610, 32'hbe896a58} /* (8, 29, 29) {real, imag} */,
  {32'hbfda96f3, 32'hbf4322c6} /* (8, 29, 28) {real, imag} */,
  {32'h3e84af16, 32'hbf57e300} /* (8, 29, 27) {real, imag} */,
  {32'hbe6275de, 32'hbdf2ee5c} /* (8, 29, 26) {real, imag} */,
  {32'hbf4471b5, 32'hbdb48a10} /* (8, 29, 25) {real, imag} */,
  {32'h3dd39718, 32'hbed7fcbc} /* (8, 29, 24) {real, imag} */,
  {32'h3c975ec0, 32'hbe2d7edd} /* (8, 29, 23) {real, imag} */,
  {32'hbe8ab030, 32'hbc674d38} /* (8, 29, 22) {real, imag} */,
  {32'h3e4fac72, 32'h3def0eaf} /* (8, 29, 21) {real, imag} */,
  {32'h3ebe90cb, 32'h3dd27004} /* (8, 29, 20) {real, imag} */,
  {32'hbdbae50c, 32'h3dc08295} /* (8, 29, 19) {real, imag} */,
  {32'hbdf2e101, 32'h3eaa0b76} /* (8, 29, 18) {real, imag} */,
  {32'hbf0d1aa0, 32'hbdda01d8} /* (8, 29, 17) {real, imag} */,
  {32'hbeef6542, 32'hbea959d7} /* (8, 29, 16) {real, imag} */,
  {32'h3e817329, 32'h3b850ff0} /* (8, 29, 15) {real, imag} */,
  {32'hbe4bf336, 32'h3e99a022} /* (8, 29, 14) {real, imag} */,
  {32'h3ec214fb, 32'hbf075f48} /* (8, 29, 13) {real, imag} */,
  {32'h3e34b810, 32'hbd8f69e6} /* (8, 29, 12) {real, imag} */,
  {32'h3d1272ea, 32'hbe907c32} /* (8, 29, 11) {real, imag} */,
  {32'h3f3014cf, 32'hbe94608e} /* (8, 29, 10) {real, imag} */,
  {32'h3c73f120, 32'h3e920a8a} /* (8, 29, 9) {real, imag} */,
  {32'hbf419c86, 32'h3f5ee8f4} /* (8, 29, 8) {real, imag} */,
  {32'hbf45f9d7, 32'hbf33ce37} /* (8, 29, 7) {real, imag} */,
  {32'hbeb77f2f, 32'hbd34a574} /* (8, 29, 6) {real, imag} */,
  {32'hbfac0982, 32'h3e453252} /* (8, 29, 5) {real, imag} */,
  {32'h3f86a215, 32'hbe300a0c} /* (8, 29, 4) {real, imag} */,
  {32'h3e94dccb, 32'hbf8a6de0} /* (8, 29, 3) {real, imag} */,
  {32'h40094744, 32'h40990739} /* (8, 29, 2) {real, imag} */,
  {32'hc0893e46, 32'hbfb626fc} /* (8, 29, 1) {real, imag} */,
  {32'h3f0dfd16, 32'h3f884645} /* (8, 29, 0) {real, imag} */,
  {32'h409b5363, 32'hc00fdba4} /* (8, 28, 31) {real, imag} */,
  {32'hc052d024, 32'h400dc6d8} /* (8, 28, 30) {real, imag} */,
  {32'hbfbf514c, 32'hbf6f7074} /* (8, 28, 29) {real, imag} */,
  {32'h3ee00eac, 32'hbdcf0ee8} /* (8, 28, 28) {real, imag} */,
  {32'hbdf3e91d, 32'h3f9139ed} /* (8, 28, 27) {real, imag} */,
  {32'h3f762477, 32'h3de4245c} /* (8, 28, 26) {real, imag} */,
  {32'h3e12b5da, 32'h3d54d568} /* (8, 28, 25) {real, imag} */,
  {32'h3ec8bd09, 32'h3fa4d9bc} /* (8, 28, 24) {real, imag} */,
  {32'hbe50dfe5, 32'hbe11c0a3} /* (8, 28, 23) {real, imag} */,
  {32'hbe99e39d, 32'hbe1558cb} /* (8, 28, 22) {real, imag} */,
  {32'h3f14bde1, 32'hbdf2f5fa} /* (8, 28, 21) {real, imag} */,
  {32'h3d232af4, 32'hbddb2d12} /* (8, 28, 20) {real, imag} */,
  {32'hbc1c3290, 32'hbf27fdbe} /* (8, 28, 19) {real, imag} */,
  {32'h3e50ba30, 32'h3e9b4534} /* (8, 28, 18) {real, imag} */,
  {32'hbe57fe1a, 32'h3e8b5554} /* (8, 28, 17) {real, imag} */,
  {32'h3ec18759, 32'h3cec4b78} /* (8, 28, 16) {real, imag} */,
  {32'hbe896498, 32'h3c520fe0} /* (8, 28, 15) {real, imag} */,
  {32'h3cf887d8, 32'h3ec984c5} /* (8, 28, 14) {real, imag} */,
  {32'hbdcf186e, 32'hbdf59e8d} /* (8, 28, 13) {real, imag} */,
  {32'h3de4a5ae, 32'hbe0acd0c} /* (8, 28, 12) {real, imag} */,
  {32'hbd05bf0c, 32'hbee22b63} /* (8, 28, 11) {real, imag} */,
  {32'h3ebc69c6, 32'h3ee94c04} /* (8, 28, 10) {real, imag} */,
  {32'h3f34e8f0, 32'h3e03a134} /* (8, 28, 9) {real, imag} */,
  {32'hbea66fa4, 32'h3edf1371} /* (8, 28, 8) {real, imag} */,
  {32'h3e79daf2, 32'hbe5571dc} /* (8, 28, 7) {real, imag} */,
  {32'hbe82be28, 32'hbe89bfce} /* (8, 28, 6) {real, imag} */,
  {32'hbf0e30f6, 32'h3ef5b074} /* (8, 28, 5) {real, imag} */,
  {32'h3f3762c1, 32'hbf13291a} /* (8, 28, 4) {real, imag} */,
  {32'hbf3d52fa, 32'h3e21fec8} /* (8, 28, 3) {real, imag} */,
  {32'hc02c3a41, 32'h40230b6d} /* (8, 28, 2) {real, imag} */,
  {32'h3f4d1bda, 32'hc043a0d8} /* (8, 28, 1) {real, imag} */,
  {32'h3fdcba62, 32'hbf4b1984} /* (8, 28, 0) {real, imag} */,
  {32'hbf61dd3a, 32'h40003406} /* (8, 27, 31) {real, imag} */,
  {32'h3f44c139, 32'hbfb5c15c} /* (8, 27, 30) {real, imag} */,
  {32'hbeff891e, 32'h3c50c570} /* (8, 27, 29) {real, imag} */,
  {32'hbf19a4ea, 32'h3e910346} /* (8, 27, 28) {real, imag} */,
  {32'h3fc1590c, 32'hbf8f191d} /* (8, 27, 27) {real, imag} */,
  {32'hbdd0a0d8, 32'hbed5a3bd} /* (8, 27, 26) {real, imag} */,
  {32'hbeb47a94, 32'h3e9fbe62} /* (8, 27, 25) {real, imag} */,
  {32'h3f156503, 32'h3e0601c4} /* (8, 27, 24) {real, imag} */,
  {32'hbdcd9140, 32'hbe97b90d} /* (8, 27, 23) {real, imag} */,
  {32'h3e6158e9, 32'hbd82028c} /* (8, 27, 22) {real, imag} */,
  {32'h3e9b0683, 32'h3f171048} /* (8, 27, 21) {real, imag} */,
  {32'h3ea1277a, 32'h3e5823c2} /* (8, 27, 20) {real, imag} */,
  {32'hbe84c9f6, 32'hbdec48ec} /* (8, 27, 19) {real, imag} */,
  {32'hbea746a6, 32'hbf327688} /* (8, 27, 18) {real, imag} */,
  {32'h3ecca738, 32'hbd0f37a4} /* (8, 27, 17) {real, imag} */,
  {32'h3e8314b3, 32'hbda63d22} /* (8, 27, 16) {real, imag} */,
  {32'hbe21ecfa, 32'h3da0f380} /* (8, 27, 15) {real, imag} */,
  {32'hbe7480f6, 32'h3ddd50da} /* (8, 27, 14) {real, imag} */,
  {32'h3e947cb8, 32'hbe42c4a4} /* (8, 27, 13) {real, imag} */,
  {32'hbeb5eb5a, 32'h3ec210f2} /* (8, 27, 12) {real, imag} */,
  {32'h3c91f7f0, 32'h3f2f835c} /* (8, 27, 11) {real, imag} */,
  {32'h3e846867, 32'h3d5b52a8} /* (8, 27, 10) {real, imag} */,
  {32'hbcd9211c, 32'hbeaf0302} /* (8, 27, 9) {real, imag} */,
  {32'h3ee75f10, 32'h3f1b53a4} /* (8, 27, 8) {real, imag} */,
  {32'h3dc812b8, 32'hbeb77a2e} /* (8, 27, 7) {real, imag} */,
  {32'hbeffec05, 32'hbf6cd200} /* (8, 27, 6) {real, imag} */,
  {32'hbe2f85c8, 32'h3e5c86c0} /* (8, 27, 5) {real, imag} */,
  {32'h3d6c1680, 32'h3e327da9} /* (8, 27, 4) {real, imag} */,
  {32'h3f396cb6, 32'hbddccd84} /* (8, 27, 3) {real, imag} */,
  {32'h3f939c8f, 32'h3f4f5082} /* (8, 27, 2) {real, imag} */,
  {32'hc0245f32, 32'h3ea68117} /* (8, 27, 1) {real, imag} */,
  {32'hc005626f, 32'h3f2f64cd} /* (8, 27, 0) {real, imag} */,
  {32'hbec1a9e0, 32'h3ec0adb2} /* (8, 26, 31) {real, imag} */,
  {32'hbf826050, 32'h3ee3b8b4} /* (8, 26, 30) {real, imag} */,
  {32'h3e0c642c, 32'hbe2a9c49} /* (8, 26, 29) {real, imag} */,
  {32'h3ef29525, 32'h3ecf2690} /* (8, 26, 28) {real, imag} */,
  {32'h3d8b4c4c, 32'h3e12a7a7} /* (8, 26, 27) {real, imag} */,
  {32'h3ea525d6, 32'hbe902f8f} /* (8, 26, 26) {real, imag} */,
  {32'hbe878555, 32'hbf932adc} /* (8, 26, 25) {real, imag} */,
  {32'h3db17a9a, 32'hbe67cab1} /* (8, 26, 24) {real, imag} */,
  {32'hbe7e0c32, 32'hbce2edb8} /* (8, 26, 23) {real, imag} */,
  {32'h3eec69ea, 32'hbe90c792} /* (8, 26, 22) {real, imag} */,
  {32'h3ec53715, 32'h3ef3b089} /* (8, 26, 21) {real, imag} */,
  {32'h3e866f9f, 32'hbe95083d} /* (8, 26, 20) {real, imag} */,
  {32'h3eac16ae, 32'h3e01eea8} /* (8, 26, 19) {real, imag} */,
  {32'h3e83ab2e, 32'hbdabbf04} /* (8, 26, 18) {real, imag} */,
  {32'h3e1cd784, 32'h3e733dc2} /* (8, 26, 17) {real, imag} */,
  {32'hbe5fc13c, 32'h3dc6a443} /* (8, 26, 16) {real, imag} */,
  {32'h3e01d552, 32'h3e82b2b7} /* (8, 26, 15) {real, imag} */,
  {32'h3e814c70, 32'h3ea81e2f} /* (8, 26, 14) {real, imag} */,
  {32'hbe0cda54, 32'hbead1013} /* (8, 26, 13) {real, imag} */,
  {32'hbf1c9498, 32'h3f3a7193} /* (8, 26, 12) {real, imag} */,
  {32'h3eb8a24b, 32'h3ce2e78c} /* (8, 26, 11) {real, imag} */,
  {32'h3eedb58a, 32'h3dfae31e} /* (8, 26, 10) {real, imag} */,
  {32'h3f0d37be, 32'hbec6f048} /* (8, 26, 9) {real, imag} */,
  {32'h3c2c5cd8, 32'h3e322f40} /* (8, 26, 8) {real, imag} */,
  {32'h3c039ff8, 32'hbd86ad42} /* (8, 26, 7) {real, imag} */,
  {32'hbed96dca, 32'hbece255c} /* (8, 26, 6) {real, imag} */,
  {32'h3ea55606, 32'hbf027fcf} /* (8, 26, 5) {real, imag} */,
  {32'hbdab32e4, 32'h3e7af4b7} /* (8, 26, 4) {real, imag} */,
  {32'h3dc391bc, 32'hbe519c6e} /* (8, 26, 3) {real, imag} */,
  {32'hbba23fc0, 32'hbdca774a} /* (8, 26, 2) {real, imag} */,
  {32'hbe93337e, 32'h3e9d0403} /* (8, 26, 1) {real, imag} */,
  {32'hbea8f784, 32'hbeed50a2} /* (8, 26, 0) {real, imag} */,
  {32'h3ec7b797, 32'hbf4725cf} /* (8, 25, 31) {real, imag} */,
  {32'hbd3a0994, 32'h3f9b4ef0} /* (8, 25, 30) {real, imag} */,
  {32'hbf79ef90, 32'hbf4cd28a} /* (8, 25, 29) {real, imag} */,
  {32'hbec3ff04, 32'hbd24ccc9} /* (8, 25, 28) {real, imag} */,
  {32'h3e8860d2, 32'hbe12faa6} /* (8, 25, 27) {real, imag} */,
  {32'hbe94a574, 32'h3e406b47} /* (8, 25, 26) {real, imag} */,
  {32'h3e91d480, 32'h3e99ba82} /* (8, 25, 25) {real, imag} */,
  {32'h3e6466f4, 32'hbeb6c616} /* (8, 25, 24) {real, imag} */,
  {32'hbe6091b0, 32'hbef14b59} /* (8, 25, 23) {real, imag} */,
  {32'hbda04e30, 32'h3d38f2b0} /* (8, 25, 22) {real, imag} */,
  {32'h3f0371a9, 32'hbdcc8b86} /* (8, 25, 21) {real, imag} */,
  {32'hbec96cbe, 32'h3e5f5733} /* (8, 25, 20) {real, imag} */,
  {32'hbef3a30a, 32'hbd2b1194} /* (8, 25, 19) {real, imag} */,
  {32'h3ecf910f, 32'hbde10a3a} /* (8, 25, 18) {real, imag} */,
  {32'h3e578e06, 32'h3ec94efe} /* (8, 25, 17) {real, imag} */,
  {32'h3ddab75e, 32'h3c0c5a30} /* (8, 25, 16) {real, imag} */,
  {32'h3e00da92, 32'h3e412dcd} /* (8, 25, 15) {real, imag} */,
  {32'h3ec22796, 32'h3eb62cdc} /* (8, 25, 14) {real, imag} */,
  {32'h3e99e5c6, 32'h3df9f117} /* (8, 25, 13) {real, imag} */,
  {32'h3e85e7e7, 32'hbdd31ec0} /* (8, 25, 12) {real, imag} */,
  {32'hbd719858, 32'hbe1bf2a8} /* (8, 25, 11) {real, imag} */,
  {32'hbca0a856, 32'hbecea660} /* (8, 25, 10) {real, imag} */,
  {32'hbee1dde2, 32'hbdd98f37} /* (8, 25, 9) {real, imag} */,
  {32'h3dd272c6, 32'h3e54e389} /* (8, 25, 8) {real, imag} */,
  {32'hbe905f5e, 32'hbe3d15d5} /* (8, 25, 7) {real, imag} */,
  {32'h3e9c9b49, 32'h3e3fe0a8} /* (8, 25, 6) {real, imag} */,
  {32'hbe0e45ce, 32'hbbf4b720} /* (8, 25, 5) {real, imag} */,
  {32'hbe98ba23, 32'hbed3e79f} /* (8, 25, 4) {real, imag} */,
  {32'h3d8bb6b6, 32'h3e972242} /* (8, 25, 3) {real, imag} */,
  {32'h3c92f940, 32'h3ee0713a} /* (8, 25, 2) {real, imag} */,
  {32'hbe147a74, 32'h3e66c954} /* (8, 25, 1) {real, imag} */,
  {32'h3f1f600c, 32'hbe8ba742} /* (8, 25, 0) {real, imag} */,
  {32'hbf471e19, 32'h3ef5166e} /* (8, 24, 31) {real, imag} */,
  {32'h3f44b48c, 32'h3b6d9780} /* (8, 24, 30) {real, imag} */,
  {32'h3d9ebc3c, 32'hbe9e50d4} /* (8, 24, 29) {real, imag} */,
  {32'hbdefa31a, 32'h3f14aa26} /* (8, 24, 28) {real, imag} */,
  {32'h3e9cd322, 32'hbda01c7e} /* (8, 24, 27) {real, imag} */,
  {32'hbd5327c0, 32'h3f15483c} /* (8, 24, 26) {real, imag} */,
  {32'hbed2cfeb, 32'hbf40a1ed} /* (8, 24, 25) {real, imag} */,
  {32'hbe42fbc4, 32'h3ece4b69} /* (8, 24, 24) {real, imag} */,
  {32'h3b9893e0, 32'hbeb91f5d} /* (8, 24, 23) {real, imag} */,
  {32'h3f0f8dbb, 32'hbe8ea5bd} /* (8, 24, 22) {real, imag} */,
  {32'h3e5910ca, 32'hbbd9d600} /* (8, 24, 21) {real, imag} */,
  {32'h3ea00028, 32'h3c2488c8} /* (8, 24, 20) {real, imag} */,
  {32'h3dad6963, 32'h3eacf958} /* (8, 24, 19) {real, imag} */,
  {32'hbed73482, 32'hbe675785} /* (8, 24, 18) {real, imag} */,
  {32'hbc318a10, 32'hbdae8d62} /* (8, 24, 17) {real, imag} */,
  {32'h3e4ba8de, 32'hbe0ad055} /* (8, 24, 16) {real, imag} */,
  {32'h3e437693, 32'hbea8a6b2} /* (8, 24, 15) {real, imag} */,
  {32'hbe7facf9, 32'h3ebd1d44} /* (8, 24, 14) {real, imag} */,
  {32'hbe5f9239, 32'h3dde8d58} /* (8, 24, 13) {real, imag} */,
  {32'h3dd5a426, 32'hbef0035b} /* (8, 24, 12) {real, imag} */,
  {32'h3d2c2baa, 32'hbdbae2c4} /* (8, 24, 11) {real, imag} */,
  {32'hbce0ae0b, 32'h3d3fc020} /* (8, 24, 10) {real, imag} */,
  {32'h3dcd317c, 32'h3e3db690} /* (8, 24, 9) {real, imag} */,
  {32'hbcc3dca8, 32'h3ef07c13} /* (8, 24, 8) {real, imag} */,
  {32'hbdb4541c, 32'hbed54ef3} /* (8, 24, 7) {real, imag} */,
  {32'h3f0e7085, 32'h3e212d66} /* (8, 24, 6) {real, imag} */,
  {32'h3ef5b960, 32'h3e836f92} /* (8, 24, 5) {real, imag} */,
  {32'h3f601a48, 32'h3a1b8f80} /* (8, 24, 4) {real, imag} */,
  {32'h3e0d2346, 32'hbd28f49a} /* (8, 24, 3) {real, imag} */,
  {32'h3f59f388, 32'h3daf43d6} /* (8, 24, 2) {real, imag} */,
  {32'hbfab588b, 32'h3f737c8e} /* (8, 24, 1) {real, imag} */,
  {32'hbf136038, 32'hbc9c9980} /* (8, 24, 0) {real, imag} */,
  {32'h3e2e3e34, 32'hbd0722d4} /* (8, 23, 31) {real, imag} */,
  {32'hbdd7e46f, 32'h3f03bd80} /* (8, 23, 30) {real, imag} */,
  {32'hbd6fbaca, 32'h3e4fcd6b} /* (8, 23, 29) {real, imag} */,
  {32'h3d95ba23, 32'hbe1322b6} /* (8, 23, 28) {real, imag} */,
  {32'hbda27b2c, 32'h3e997c32} /* (8, 23, 27) {real, imag} */,
  {32'hbeb08120, 32'h3dc5997a} /* (8, 23, 26) {real, imag} */,
  {32'hbe490e47, 32'hbe9f85ba} /* (8, 23, 25) {real, imag} */,
  {32'hbe1b03f5, 32'h3c9a4628} /* (8, 23, 24) {real, imag} */,
  {32'hbed3f2af, 32'hbf0018ce} /* (8, 23, 23) {real, imag} */,
  {32'hbe411e19, 32'hbe663bff} /* (8, 23, 22) {real, imag} */,
  {32'h3df5311c, 32'h3d420a96} /* (8, 23, 21) {real, imag} */,
  {32'h3f28f4ea, 32'h3ec9c5c7} /* (8, 23, 20) {real, imag} */,
  {32'h3d2a1ac8, 32'h3ef65ef1} /* (8, 23, 19) {real, imag} */,
  {32'h3d3c5d70, 32'hbe85b13e} /* (8, 23, 18) {real, imag} */,
  {32'hbe72c9bc, 32'hbede0108} /* (8, 23, 17) {real, imag} */,
  {32'h3d82d384, 32'hbe3e27b1} /* (8, 23, 16) {real, imag} */,
  {32'hbd9b7c33, 32'h3e0e8632} /* (8, 23, 15) {real, imag} */,
  {32'hbe651436, 32'hbdac8e8e} /* (8, 23, 14) {real, imag} */,
  {32'hbe5363be, 32'h3e86977a} /* (8, 23, 13) {real, imag} */,
  {32'h3eec6859, 32'hbe361877} /* (8, 23, 12) {real, imag} */,
  {32'h3e3222a0, 32'hbf54de4c} /* (8, 23, 11) {real, imag} */,
  {32'h3e9cdd0c, 32'h3e69511c} /* (8, 23, 10) {real, imag} */,
  {32'hbcbd1fe0, 32'hbe7fe028} /* (8, 23, 9) {real, imag} */,
  {32'hbe293a42, 32'hbe5e5bd6} /* (8, 23, 8) {real, imag} */,
  {32'hbcf9a7f4, 32'h3f1895d0} /* (8, 23, 7) {real, imag} */,
  {32'hbdb22c92, 32'h3ee73680} /* (8, 23, 6) {real, imag} */,
  {32'hbf0ff435, 32'h3d9502f0} /* (8, 23, 5) {real, imag} */,
  {32'hbf1a9344, 32'h3cdea538} /* (8, 23, 4) {real, imag} */,
  {32'h3e440757, 32'hbca37808} /* (8, 23, 3) {real, imag} */,
  {32'h3f001be1, 32'h3f482d02} /* (8, 23, 2) {real, imag} */,
  {32'hbf375939, 32'hbf2ed1db} /* (8, 23, 1) {real, imag} */,
  {32'hbf3f00d0, 32'h3f5687ce} /* (8, 23, 0) {real, imag} */,
  {32'hbe2d8c29, 32'h3dca7a20} /* (8, 22, 31) {real, imag} */,
  {32'h3eca5af5, 32'hbe3fcc9a} /* (8, 22, 30) {real, imag} */,
  {32'hbebb5051, 32'hbcec78da} /* (8, 22, 29) {real, imag} */,
  {32'h3ebf70de, 32'hbe8ac131} /* (8, 22, 28) {real, imag} */,
  {32'hbec315e2, 32'h3dd06771} /* (8, 22, 27) {real, imag} */,
  {32'hbf27dd91, 32'h3cabeaf8} /* (8, 22, 26) {real, imag} */,
  {32'h3e4dfa1c, 32'h3e95ff91} /* (8, 22, 25) {real, imag} */,
  {32'hbcfd9608, 32'hbe6d07b5} /* (8, 22, 24) {real, imag} */,
  {32'h3f2562d9, 32'h3e4b6f1b} /* (8, 22, 23) {real, imag} */,
  {32'h3e13403a, 32'h3e75245a} /* (8, 22, 22) {real, imag} */,
  {32'h3aa40b00, 32'hbe36ad7c} /* (8, 22, 21) {real, imag} */,
  {32'h3eae1097, 32'h3e173398} /* (8, 22, 20) {real, imag} */,
  {32'h3d935819, 32'hbeb23515} /* (8, 22, 19) {real, imag} */,
  {32'hbdc84b42, 32'h3ddd3018} /* (8, 22, 18) {real, imag} */,
  {32'h3d47fd52, 32'hbe869a98} /* (8, 22, 17) {real, imag} */,
  {32'hbe69f8aa, 32'hbdd1bed6} /* (8, 22, 16) {real, imag} */,
  {32'h3e87b5ef, 32'h3ddb90a8} /* (8, 22, 15) {real, imag} */,
  {32'h3cf22020, 32'h3e00fdc8} /* (8, 22, 14) {real, imag} */,
  {32'h3eb94fca, 32'hbe85d9a4} /* (8, 22, 13) {real, imag} */,
  {32'h3e9d7941, 32'h3cbb224c} /* (8, 22, 12) {real, imag} */,
  {32'h3eaa4f8a, 32'hbe9e9dbc} /* (8, 22, 11) {real, imag} */,
  {32'hbd873572, 32'h3e2c138b} /* (8, 22, 10) {real, imag} */,
  {32'hbee86a9b, 32'h3e6e3314} /* (8, 22, 9) {real, imag} */,
  {32'hbe4067f1, 32'h3ebb7f13} /* (8, 22, 8) {real, imag} */,
  {32'hbf0ec2d2, 32'h3db72eea} /* (8, 22, 7) {real, imag} */,
  {32'hbed3bc4d, 32'hbe4d4586} /* (8, 22, 6) {real, imag} */,
  {32'h3dd2d82c, 32'hbe69bf85} /* (8, 22, 5) {real, imag} */,
  {32'h3f29b56d, 32'h3d7b3d02} /* (8, 22, 4) {real, imag} */,
  {32'hbbb5b3c0, 32'h3e1983d6} /* (8, 22, 3) {real, imag} */,
  {32'hbea0172c, 32'h3d8884f8} /* (8, 22, 2) {real, imag} */,
  {32'h3c032b70, 32'h3d617bc8} /* (8, 22, 1) {real, imag} */,
  {32'hbe7a5f81, 32'hbe9d3b3a} /* (8, 22, 0) {real, imag} */,
  {32'hbdeffe40, 32'h3eedc1f0} /* (8, 21, 31) {real, imag} */,
  {32'h3e940654, 32'hbea62ab4} /* (8, 21, 30) {real, imag} */,
  {32'hbd5b6708, 32'hbe85d7ee} /* (8, 21, 29) {real, imag} */,
  {32'h3ec05847, 32'h3da04283} /* (8, 21, 28) {real, imag} */,
  {32'hbf55675d, 32'h3dd1725d} /* (8, 21, 27) {real, imag} */,
  {32'h3def1ea0, 32'hbd3ae576} /* (8, 21, 26) {real, imag} */,
  {32'hbe65c5c7, 32'h3e11e722} /* (8, 21, 25) {real, imag} */,
  {32'hbed94768, 32'h3f023c90} /* (8, 21, 24) {real, imag} */,
  {32'h3ed3a870, 32'h3cef63f0} /* (8, 21, 23) {real, imag} */,
  {32'hbf2d1132, 32'hbf89808d} /* (8, 21, 22) {real, imag} */,
  {32'h3ddaa7eb, 32'hbe361875} /* (8, 21, 21) {real, imag} */,
  {32'hbebb9580, 32'h3e5529b4} /* (8, 21, 20) {real, imag} */,
  {32'hbf9a57ec, 32'hbe4217a2} /* (8, 21, 19) {real, imag} */,
  {32'h3df24476, 32'h3dc5c6de} /* (8, 21, 18) {real, imag} */,
  {32'h3e0c9fca, 32'h3d1e3f94} /* (8, 21, 17) {real, imag} */,
  {32'h3cdf0d10, 32'h3e61f965} /* (8, 21, 16) {real, imag} */,
  {32'h3c531500, 32'hbedb2730} /* (8, 21, 15) {real, imag} */,
  {32'hbc2e9c68, 32'h3e880698} /* (8, 21, 14) {real, imag} */,
  {32'h3d41f4f6, 32'h3e7666f6} /* (8, 21, 13) {real, imag} */,
  {32'h3eee6cb2, 32'hbea80ce9} /* (8, 21, 12) {real, imag} */,
  {32'h3e91e5b4, 32'h3ea629f5} /* (8, 21, 11) {real, imag} */,
  {32'hbea809dd, 32'h3d880f88} /* (8, 21, 10) {real, imag} */,
  {32'hbe162e51, 32'hbd1c200a} /* (8, 21, 9) {real, imag} */,
  {32'hbdf316e6, 32'h3d80e447} /* (8, 21, 8) {real, imag} */,
  {32'hbe1a6464, 32'h3deeb3aa} /* (8, 21, 7) {real, imag} */,
  {32'h3dd299e0, 32'h3e971ca4} /* (8, 21, 6) {real, imag} */,
  {32'h3f241030, 32'hbd99b1ba} /* (8, 21, 5) {real, imag} */,
  {32'h3e199a44, 32'hbeea3174} /* (8, 21, 4) {real, imag} */,
  {32'hbda49d82, 32'h3da3a120} /* (8, 21, 3) {real, imag} */,
  {32'h3dfc0f6c, 32'hbee03e2a} /* (8, 21, 2) {real, imag} */,
  {32'h3e7dfe98, 32'hbda7f2ca} /* (8, 21, 1) {real, imag} */,
  {32'hbf5e58f0, 32'h3f719ffb} /* (8, 21, 0) {real, imag} */,
  {32'h3e964e44, 32'hbe2767df} /* (8, 20, 31) {real, imag} */,
  {32'hbe4f9ebc, 32'hbf044609} /* (8, 20, 30) {real, imag} */,
  {32'h3e1690b5, 32'h3ed008e3} /* (8, 20, 29) {real, imag} */,
  {32'hbe2bb416, 32'h3dbc0d68} /* (8, 20, 28) {real, imag} */,
  {32'h3f331400, 32'hbec98edf} /* (8, 20, 27) {real, imag} */,
  {32'h3e2c6c5d, 32'h3d3ea744} /* (8, 20, 26) {real, imag} */,
  {32'hbebc7917, 32'hbd9626de} /* (8, 20, 25) {real, imag} */,
  {32'hbdeaa95c, 32'hbf3cc3af} /* (8, 20, 24) {real, imag} */,
  {32'h3f02d65b, 32'h3e9e3488} /* (8, 20, 23) {real, imag} */,
  {32'hbdbf40d0, 32'hbc68ac20} /* (8, 20, 22) {real, imag} */,
  {32'hbe0b7635, 32'h3e229e51} /* (8, 20, 21) {real, imag} */,
  {32'h3ee67d72, 32'h3e86a9d9} /* (8, 20, 20) {real, imag} */,
  {32'hbf25fd20, 32'hbcaeaa56} /* (8, 20, 19) {real, imag} */,
  {32'hbdb2a3cf, 32'hbe84ae1c} /* (8, 20, 18) {real, imag} */,
  {32'hbc0e81a0, 32'h3eb70b26} /* (8, 20, 17) {real, imag} */,
  {32'hbdc11a54, 32'h3d24a7fb} /* (8, 20, 16) {real, imag} */,
  {32'hbc056ee0, 32'hbe1df81c} /* (8, 20, 15) {real, imag} */,
  {32'hbf0f969b, 32'hbe433a74} /* (8, 20, 14) {real, imag} */,
  {32'hbe97baba, 32'hbe630d05} /* (8, 20, 13) {real, imag} */,
  {32'hbeb42018, 32'h3f2e2721} /* (8, 20, 12) {real, imag} */,
  {32'h3c9eabb0, 32'hbe9b6490} /* (8, 20, 11) {real, imag} */,
  {32'h3f254578, 32'hbec38cf4} /* (8, 20, 10) {real, imag} */,
  {32'hbeb740dd, 32'h3e57cb75} /* (8, 20, 9) {real, imag} */,
  {32'hbd547254, 32'hbe2c0f58} /* (8, 20, 8) {real, imag} */,
  {32'h3e9bdbd0, 32'hbecd104e} /* (8, 20, 7) {real, imag} */,
  {32'hbe9fa9a6, 32'h3f1922f0} /* (8, 20, 6) {real, imag} */,
  {32'hbd8cf69e, 32'h3ef71a44} /* (8, 20, 5) {real, imag} */,
  {32'hbe71c692, 32'h3e14ec5a} /* (8, 20, 4) {real, imag} */,
  {32'h3e7b81ee, 32'hbe044b1c} /* (8, 20, 3) {real, imag} */,
  {32'h3d9d0cf0, 32'h3e31f03c} /* (8, 20, 2) {real, imag} */,
  {32'h3db57610, 32'h3ea56b63} /* (8, 20, 1) {real, imag} */,
  {32'h3e4dc9ca, 32'hbf24456d} /* (8, 20, 0) {real, imag} */,
  {32'hbd560340, 32'hbf5f2a90} /* (8, 19, 31) {real, imag} */,
  {32'h3edf8476, 32'h3e06bf90} /* (8, 19, 30) {real, imag} */,
  {32'h3ec70a8a, 32'hbe460a50} /* (8, 19, 29) {real, imag} */,
  {32'hbe4b0e2a, 32'hbd24fce8} /* (8, 19, 28) {real, imag} */,
  {32'h3e318cee, 32'h3e21d524} /* (8, 19, 27) {real, imag} */,
  {32'h3ec35672, 32'hbd397b96} /* (8, 19, 26) {real, imag} */,
  {32'h3f07d2ae, 32'hbe0118e3} /* (8, 19, 25) {real, imag} */,
  {32'h3ef09d9e, 32'h3ee100cc} /* (8, 19, 24) {real, imag} */,
  {32'hbde1841e, 32'h3ef0edfd} /* (8, 19, 23) {real, imag} */,
  {32'h3f0754ba, 32'h3ddb34a1} /* (8, 19, 22) {real, imag} */,
  {32'hbda34285, 32'h3ef796d4} /* (8, 19, 21) {real, imag} */,
  {32'h3e1de766, 32'h3d2cb26e} /* (8, 19, 20) {real, imag} */,
  {32'hbd9bf15e, 32'hbed31dab} /* (8, 19, 19) {real, imag} */,
  {32'h3e702d84, 32'h3e6f9274} /* (8, 19, 18) {real, imag} */,
  {32'hbe4bd461, 32'h3f0324c6} /* (8, 19, 17) {real, imag} */,
  {32'hbe546d20, 32'hbdf051fc} /* (8, 19, 16) {real, imag} */,
  {32'hbe23d86a, 32'h3d295134} /* (8, 19, 15) {real, imag} */,
  {32'h3c7faf78, 32'h3d58aad2} /* (8, 19, 14) {real, imag} */,
  {32'h3db22354, 32'hbe2b7052} /* (8, 19, 13) {real, imag} */,
  {32'h3e620512, 32'hbe54add5} /* (8, 19, 12) {real, imag} */,
  {32'h3c738708, 32'h3eb266ea} /* (8, 19, 11) {real, imag} */,
  {32'hbf17b72e, 32'hbd0d4124} /* (8, 19, 10) {real, imag} */,
  {32'hbc03c000, 32'hbde6dccf} /* (8, 19, 9) {real, imag} */,
  {32'h3ea198f4, 32'hbdee8b9d} /* (8, 19, 8) {real, imag} */,
  {32'h3e5a69d9, 32'hbe77b405} /* (8, 19, 7) {real, imag} */,
  {32'hbd302a70, 32'hbedbd2ba} /* (8, 19, 6) {real, imag} */,
  {32'h3b27c080, 32'hbe469d80} /* (8, 19, 5) {real, imag} */,
  {32'h3ebc6651, 32'hbe698e8c} /* (8, 19, 4) {real, imag} */,
  {32'h3e3ee376, 32'hbf17228e} /* (8, 19, 3) {real, imag} */,
  {32'hbe1dd4cc, 32'hbe758c77} /* (8, 19, 2) {real, imag} */,
  {32'hbe48bcfe, 32'hbd077c8c} /* (8, 19, 1) {real, imag} */,
  {32'h3ea4106c, 32'hbd67d78c} /* (8, 19, 0) {real, imag} */,
  {32'h3ed3cbfc, 32'h3ebe0170} /* (8, 18, 31) {real, imag} */,
  {32'h3e5e92e4, 32'h3cce3590} /* (8, 18, 30) {real, imag} */,
  {32'hbd3468ae, 32'hbe422841} /* (8, 18, 29) {real, imag} */,
  {32'hbd893222, 32'hbdb19555} /* (8, 18, 28) {real, imag} */,
  {32'hbd4bf918, 32'hbe162fc3} /* (8, 18, 27) {real, imag} */,
  {32'hbe4d9866, 32'h3e3b6f6b} /* (8, 18, 26) {real, imag} */,
  {32'hbe82d1bb, 32'h3e2486a8} /* (8, 18, 25) {real, imag} */,
  {32'h3e2e1984, 32'hbdb89546} /* (8, 18, 24) {real, imag} */,
  {32'h3dad071c, 32'h3e99f14b} /* (8, 18, 23) {real, imag} */,
  {32'hbf35da82, 32'hbe9a5929} /* (8, 18, 22) {real, imag} */,
  {32'h3cacc550, 32'hbeb9f222} /* (8, 18, 21) {real, imag} */,
  {32'h3d17e292, 32'h3e1677bf} /* (8, 18, 20) {real, imag} */,
  {32'h3e859c40, 32'hbd6b6bb4} /* (8, 18, 19) {real, imag} */,
  {32'h3e9dd618, 32'hbea68fc6} /* (8, 18, 18) {real, imag} */,
  {32'h3e9217a2, 32'h3ea6007e} /* (8, 18, 17) {real, imag} */,
  {32'hbf0b1ffe, 32'h3d8c377c} /* (8, 18, 16) {real, imag} */,
  {32'hbccad3cc, 32'hbebfefff} /* (8, 18, 15) {real, imag} */,
  {32'h3e406da6, 32'hbf1681eb} /* (8, 18, 14) {real, imag} */,
  {32'h3ef8a3fa, 32'h3f2de270} /* (8, 18, 13) {real, imag} */,
  {32'hba164c80, 32'hbd6c8ea0} /* (8, 18, 12) {real, imag} */,
  {32'h3e81ae28, 32'hbe54a2f5} /* (8, 18, 11) {real, imag} */,
  {32'hbe6fcd54, 32'hbdfb8b1e} /* (8, 18, 10) {real, imag} */,
  {32'h3e45076d, 32'hbf0b0d72} /* (8, 18, 9) {real, imag} */,
  {32'h3ed291d2, 32'hbea28c56} /* (8, 18, 8) {real, imag} */,
  {32'h3e79f6af, 32'hbce6ef0a} /* (8, 18, 7) {real, imag} */,
  {32'hbf03255f, 32'hbdc48660} /* (8, 18, 6) {real, imag} */,
  {32'hbe158731, 32'h3eb8ac37} /* (8, 18, 5) {real, imag} */,
  {32'hbd0a8f68, 32'h3ee625a4} /* (8, 18, 4) {real, imag} */,
  {32'hbeadf0c4, 32'h3ef3deb8} /* (8, 18, 3) {real, imag} */,
  {32'h3ef0c486, 32'hbebc062e} /* (8, 18, 2) {real, imag} */,
  {32'hbe862702, 32'h3ea6ea14} /* (8, 18, 1) {real, imag} */,
  {32'h3c8ca660, 32'h3dabf25a} /* (8, 18, 0) {real, imag} */,
  {32'h3d0e012d, 32'hbeb3a4ea} /* (8, 17, 31) {real, imag} */,
  {32'h3e8c50c6, 32'h3e1cfc3b} /* (8, 17, 30) {real, imag} */,
  {32'hbdab26d9, 32'h3e5fb314} /* (8, 17, 29) {real, imag} */,
  {32'hbed946f0, 32'h3e07ec6e} /* (8, 17, 28) {real, imag} */,
  {32'hbe0ca3c6, 32'h3e1a15b2} /* (8, 17, 27) {real, imag} */,
  {32'h3e7ac458, 32'h3da669fc} /* (8, 17, 26) {real, imag} */,
  {32'hbe4c4750, 32'hbf096a83} /* (8, 17, 25) {real, imag} */,
  {32'hbe46a24e, 32'h3eda9349} /* (8, 17, 24) {real, imag} */,
  {32'hbeeca334, 32'h3ee68d29} /* (8, 17, 23) {real, imag} */,
  {32'hbdb38cf8, 32'h3e59e5ee} /* (8, 17, 22) {real, imag} */,
  {32'h3df06822, 32'h3d2e9684} /* (8, 17, 21) {real, imag} */,
  {32'hbe547a24, 32'h3e9bbb61} /* (8, 17, 20) {real, imag} */,
  {32'h3eb9af5d, 32'h3e457532} /* (8, 17, 19) {real, imag} */,
  {32'h3e59f8e6, 32'hbd933b6a} /* (8, 17, 18) {real, imag} */,
  {32'h3e023d30, 32'hbe3a3d87} /* (8, 17, 17) {real, imag} */,
  {32'h3d5e628a, 32'hbe71ee05} /* (8, 17, 16) {real, imag} */,
  {32'h3d894588, 32'hbe9614e8} /* (8, 17, 15) {real, imag} */,
  {32'h3e1b4bc4, 32'h3da486b5} /* (8, 17, 14) {real, imag} */,
  {32'hbd97cf07, 32'hbd18820d} /* (8, 17, 13) {real, imag} */,
  {32'h3c4ae3e8, 32'hbe37ed34} /* (8, 17, 12) {real, imag} */,
  {32'hbeb7caba, 32'h3e43dd1d} /* (8, 17, 11) {real, imag} */,
  {32'hbed5a555, 32'h3ea2f15a} /* (8, 17, 10) {real, imag} */,
  {32'h3e4c4202, 32'h3ee928ce} /* (8, 17, 9) {real, imag} */,
  {32'h3e917906, 32'h3dc245a0} /* (8, 17, 8) {real, imag} */,
  {32'hbd80e1bc, 32'h3e2641bc} /* (8, 17, 7) {real, imag} */,
  {32'h3ea4e711, 32'hbe9a6108} /* (8, 17, 6) {real, imag} */,
  {32'h3d9ccc46, 32'h38d27400} /* (8, 17, 5) {real, imag} */,
  {32'h3e996059, 32'hbd3ab5dd} /* (8, 17, 4) {real, imag} */,
  {32'hbea9a8a8, 32'hbe86613c} /* (8, 17, 3) {real, imag} */,
  {32'hbdb7b425, 32'hbe5e7c51} /* (8, 17, 2) {real, imag} */,
  {32'hbdb23438, 32'hbe0f1eba} /* (8, 17, 1) {real, imag} */,
  {32'hbdb391aa, 32'h3d8b89ec} /* (8, 17, 0) {real, imag} */,
  {32'hbdf1a164, 32'hbdbd0f4b} /* (8, 16, 31) {real, imag} */,
  {32'h3cd15d20, 32'h3e5df9d8} /* (8, 16, 30) {real, imag} */,
  {32'hbecec1f0, 32'h3e63ae31} /* (8, 16, 29) {real, imag} */,
  {32'hbdc2d52a, 32'hbce642b4} /* (8, 16, 28) {real, imag} */,
  {32'h3d2e27a4, 32'hbdbf2e16} /* (8, 16, 27) {real, imag} */,
  {32'h3cd76894, 32'h3e952469} /* (8, 16, 26) {real, imag} */,
  {32'hbdf7881e, 32'h3b95c4c0} /* (8, 16, 25) {real, imag} */,
  {32'hbe8d6653, 32'h3e011a58} /* (8, 16, 24) {real, imag} */,
  {32'hbf09dcba, 32'hbea9071c} /* (8, 16, 23) {real, imag} */,
  {32'hbdf633f4, 32'hbeb660f1} /* (8, 16, 22) {real, imag} */,
  {32'h3e845d9c, 32'hbe0bc16b} /* (8, 16, 21) {real, imag} */,
  {32'h3c361460, 32'hbdf39e24} /* (8, 16, 20) {real, imag} */,
  {32'hbd87c45e, 32'hbe01fba8} /* (8, 16, 19) {real, imag} */,
  {32'hbf146b04, 32'hbd66915f} /* (8, 16, 18) {real, imag} */,
  {32'h3dec8df0, 32'hbdcbea1b} /* (8, 16, 17) {real, imag} */,
  {32'h3ecc5874, 32'h00000000} /* (8, 16, 16) {real, imag} */,
  {32'h3dec8df0, 32'h3dcbea1b} /* (8, 16, 15) {real, imag} */,
  {32'hbf146b04, 32'h3d66915f} /* (8, 16, 14) {real, imag} */,
  {32'hbd87c45e, 32'h3e01fba8} /* (8, 16, 13) {real, imag} */,
  {32'h3c361460, 32'h3df39e24} /* (8, 16, 12) {real, imag} */,
  {32'h3e845d9c, 32'h3e0bc16b} /* (8, 16, 11) {real, imag} */,
  {32'hbdf633f4, 32'h3eb660f1} /* (8, 16, 10) {real, imag} */,
  {32'hbf09dcba, 32'h3ea9071c} /* (8, 16, 9) {real, imag} */,
  {32'hbe8d6653, 32'hbe011a58} /* (8, 16, 8) {real, imag} */,
  {32'hbdf7881e, 32'hbb95c4c0} /* (8, 16, 7) {real, imag} */,
  {32'h3cd76894, 32'hbe952469} /* (8, 16, 6) {real, imag} */,
  {32'h3d2e27a4, 32'h3dbf2e16} /* (8, 16, 5) {real, imag} */,
  {32'hbdc2d52a, 32'h3ce642b4} /* (8, 16, 4) {real, imag} */,
  {32'hbecec1f0, 32'hbe63ae31} /* (8, 16, 3) {real, imag} */,
  {32'h3cd15d20, 32'hbe5df9d8} /* (8, 16, 2) {real, imag} */,
  {32'hbdf1a164, 32'h3dbd0f4b} /* (8, 16, 1) {real, imag} */,
  {32'h3e7d9edc, 32'h00000000} /* (8, 16, 0) {real, imag} */,
  {32'hbdb23438, 32'h3e0f1eba} /* (8, 15, 31) {real, imag} */,
  {32'hbdb7b425, 32'h3e5e7c51} /* (8, 15, 30) {real, imag} */,
  {32'hbea9a8a8, 32'h3e86613c} /* (8, 15, 29) {real, imag} */,
  {32'h3e996059, 32'h3d3ab5dd} /* (8, 15, 28) {real, imag} */,
  {32'h3d9ccc46, 32'hb8d27400} /* (8, 15, 27) {real, imag} */,
  {32'h3ea4e711, 32'h3e9a6108} /* (8, 15, 26) {real, imag} */,
  {32'hbd80e1bc, 32'hbe2641bc} /* (8, 15, 25) {real, imag} */,
  {32'h3e917906, 32'hbdc245a0} /* (8, 15, 24) {real, imag} */,
  {32'h3e4c4202, 32'hbee928ce} /* (8, 15, 23) {real, imag} */,
  {32'hbed5a555, 32'hbea2f15a} /* (8, 15, 22) {real, imag} */,
  {32'hbeb7caba, 32'hbe43dd1d} /* (8, 15, 21) {real, imag} */,
  {32'h3c4ae3e8, 32'h3e37ed34} /* (8, 15, 20) {real, imag} */,
  {32'hbd97cf07, 32'h3d18820d} /* (8, 15, 19) {real, imag} */,
  {32'h3e1b4bc4, 32'hbda486b5} /* (8, 15, 18) {real, imag} */,
  {32'h3d894588, 32'h3e9614e8} /* (8, 15, 17) {real, imag} */,
  {32'h3d5e628a, 32'h3e71ee05} /* (8, 15, 16) {real, imag} */,
  {32'h3e023d30, 32'h3e3a3d87} /* (8, 15, 15) {real, imag} */,
  {32'h3e59f8e6, 32'h3d933b6a} /* (8, 15, 14) {real, imag} */,
  {32'h3eb9af5d, 32'hbe457532} /* (8, 15, 13) {real, imag} */,
  {32'hbe547a24, 32'hbe9bbb61} /* (8, 15, 12) {real, imag} */,
  {32'h3df06822, 32'hbd2e9684} /* (8, 15, 11) {real, imag} */,
  {32'hbdb38cf8, 32'hbe59e5ee} /* (8, 15, 10) {real, imag} */,
  {32'hbeeca334, 32'hbee68d29} /* (8, 15, 9) {real, imag} */,
  {32'hbe46a24e, 32'hbeda9349} /* (8, 15, 8) {real, imag} */,
  {32'hbe4c4750, 32'h3f096a83} /* (8, 15, 7) {real, imag} */,
  {32'h3e7ac458, 32'hbda669fc} /* (8, 15, 6) {real, imag} */,
  {32'hbe0ca3c6, 32'hbe1a15b2} /* (8, 15, 5) {real, imag} */,
  {32'hbed946f0, 32'hbe07ec6e} /* (8, 15, 4) {real, imag} */,
  {32'hbdab26d9, 32'hbe5fb314} /* (8, 15, 3) {real, imag} */,
  {32'h3e8c50c6, 32'hbe1cfc3b} /* (8, 15, 2) {real, imag} */,
  {32'h3d0e012d, 32'h3eb3a4ea} /* (8, 15, 1) {real, imag} */,
  {32'hbdb391aa, 32'hbd8b89ec} /* (8, 15, 0) {real, imag} */,
  {32'hbe862702, 32'hbea6ea14} /* (8, 14, 31) {real, imag} */,
  {32'h3ef0c486, 32'h3ebc062e} /* (8, 14, 30) {real, imag} */,
  {32'hbeadf0c4, 32'hbef3deb8} /* (8, 14, 29) {real, imag} */,
  {32'hbd0a8f68, 32'hbee625a4} /* (8, 14, 28) {real, imag} */,
  {32'hbe158731, 32'hbeb8ac37} /* (8, 14, 27) {real, imag} */,
  {32'hbf03255f, 32'h3dc48660} /* (8, 14, 26) {real, imag} */,
  {32'h3e79f6af, 32'h3ce6ef0a} /* (8, 14, 25) {real, imag} */,
  {32'h3ed291d2, 32'h3ea28c56} /* (8, 14, 24) {real, imag} */,
  {32'h3e45076d, 32'h3f0b0d72} /* (8, 14, 23) {real, imag} */,
  {32'hbe6fcd54, 32'h3dfb8b1e} /* (8, 14, 22) {real, imag} */,
  {32'h3e81ae28, 32'h3e54a2f5} /* (8, 14, 21) {real, imag} */,
  {32'hba164c80, 32'h3d6c8ea0} /* (8, 14, 20) {real, imag} */,
  {32'h3ef8a3fa, 32'hbf2de270} /* (8, 14, 19) {real, imag} */,
  {32'h3e406da6, 32'h3f1681eb} /* (8, 14, 18) {real, imag} */,
  {32'hbccad3cc, 32'h3ebfefff} /* (8, 14, 17) {real, imag} */,
  {32'hbf0b1ffe, 32'hbd8c377c} /* (8, 14, 16) {real, imag} */,
  {32'h3e9217a2, 32'hbea6007e} /* (8, 14, 15) {real, imag} */,
  {32'h3e9dd618, 32'h3ea68fc6} /* (8, 14, 14) {real, imag} */,
  {32'h3e859c40, 32'h3d6b6bb4} /* (8, 14, 13) {real, imag} */,
  {32'h3d17e292, 32'hbe1677bf} /* (8, 14, 12) {real, imag} */,
  {32'h3cacc550, 32'h3eb9f222} /* (8, 14, 11) {real, imag} */,
  {32'hbf35da82, 32'h3e9a5929} /* (8, 14, 10) {real, imag} */,
  {32'h3dad071c, 32'hbe99f14b} /* (8, 14, 9) {real, imag} */,
  {32'h3e2e1984, 32'h3db89546} /* (8, 14, 8) {real, imag} */,
  {32'hbe82d1bb, 32'hbe2486a8} /* (8, 14, 7) {real, imag} */,
  {32'hbe4d9866, 32'hbe3b6f6b} /* (8, 14, 6) {real, imag} */,
  {32'hbd4bf918, 32'h3e162fc3} /* (8, 14, 5) {real, imag} */,
  {32'hbd893222, 32'h3db19555} /* (8, 14, 4) {real, imag} */,
  {32'hbd3468ae, 32'h3e422841} /* (8, 14, 3) {real, imag} */,
  {32'h3e5e92e4, 32'hbcce3590} /* (8, 14, 2) {real, imag} */,
  {32'h3ed3cbfc, 32'hbebe0170} /* (8, 14, 1) {real, imag} */,
  {32'h3c8ca660, 32'hbdabf25a} /* (8, 14, 0) {real, imag} */,
  {32'hbe48bcfe, 32'h3d077c8c} /* (8, 13, 31) {real, imag} */,
  {32'hbe1dd4cc, 32'h3e758c77} /* (8, 13, 30) {real, imag} */,
  {32'h3e3ee376, 32'h3f17228e} /* (8, 13, 29) {real, imag} */,
  {32'h3ebc6651, 32'h3e698e8c} /* (8, 13, 28) {real, imag} */,
  {32'h3b27c080, 32'h3e469d80} /* (8, 13, 27) {real, imag} */,
  {32'hbd302a70, 32'h3edbd2ba} /* (8, 13, 26) {real, imag} */,
  {32'h3e5a69d9, 32'h3e77b405} /* (8, 13, 25) {real, imag} */,
  {32'h3ea198f4, 32'h3dee8b9d} /* (8, 13, 24) {real, imag} */,
  {32'hbc03c000, 32'h3de6dccf} /* (8, 13, 23) {real, imag} */,
  {32'hbf17b72e, 32'h3d0d4124} /* (8, 13, 22) {real, imag} */,
  {32'h3c738708, 32'hbeb266ea} /* (8, 13, 21) {real, imag} */,
  {32'h3e620512, 32'h3e54add5} /* (8, 13, 20) {real, imag} */,
  {32'h3db22354, 32'h3e2b7052} /* (8, 13, 19) {real, imag} */,
  {32'h3c7faf78, 32'hbd58aad2} /* (8, 13, 18) {real, imag} */,
  {32'hbe23d86a, 32'hbd295134} /* (8, 13, 17) {real, imag} */,
  {32'hbe546d20, 32'h3df051fc} /* (8, 13, 16) {real, imag} */,
  {32'hbe4bd461, 32'hbf0324c6} /* (8, 13, 15) {real, imag} */,
  {32'h3e702d84, 32'hbe6f9274} /* (8, 13, 14) {real, imag} */,
  {32'hbd9bf15e, 32'h3ed31dab} /* (8, 13, 13) {real, imag} */,
  {32'h3e1de766, 32'hbd2cb26e} /* (8, 13, 12) {real, imag} */,
  {32'hbda34285, 32'hbef796d4} /* (8, 13, 11) {real, imag} */,
  {32'h3f0754ba, 32'hbddb34a1} /* (8, 13, 10) {real, imag} */,
  {32'hbde1841e, 32'hbef0edfd} /* (8, 13, 9) {real, imag} */,
  {32'h3ef09d9e, 32'hbee100cc} /* (8, 13, 8) {real, imag} */,
  {32'h3f07d2ae, 32'h3e0118e3} /* (8, 13, 7) {real, imag} */,
  {32'h3ec35672, 32'h3d397b96} /* (8, 13, 6) {real, imag} */,
  {32'h3e318cee, 32'hbe21d524} /* (8, 13, 5) {real, imag} */,
  {32'hbe4b0e2a, 32'h3d24fce8} /* (8, 13, 4) {real, imag} */,
  {32'h3ec70a8a, 32'h3e460a50} /* (8, 13, 3) {real, imag} */,
  {32'h3edf8476, 32'hbe06bf90} /* (8, 13, 2) {real, imag} */,
  {32'hbd560340, 32'h3f5f2a90} /* (8, 13, 1) {real, imag} */,
  {32'h3ea4106c, 32'h3d67d78c} /* (8, 13, 0) {real, imag} */,
  {32'h3db57610, 32'hbea56b63} /* (8, 12, 31) {real, imag} */,
  {32'h3d9d0cf0, 32'hbe31f03c} /* (8, 12, 30) {real, imag} */,
  {32'h3e7b81ee, 32'h3e044b1c} /* (8, 12, 29) {real, imag} */,
  {32'hbe71c692, 32'hbe14ec5a} /* (8, 12, 28) {real, imag} */,
  {32'hbd8cf69e, 32'hbef71a44} /* (8, 12, 27) {real, imag} */,
  {32'hbe9fa9a6, 32'hbf1922f0} /* (8, 12, 26) {real, imag} */,
  {32'h3e9bdbd0, 32'h3ecd104e} /* (8, 12, 25) {real, imag} */,
  {32'hbd547254, 32'h3e2c0f58} /* (8, 12, 24) {real, imag} */,
  {32'hbeb740dd, 32'hbe57cb75} /* (8, 12, 23) {real, imag} */,
  {32'h3f254578, 32'h3ec38cf4} /* (8, 12, 22) {real, imag} */,
  {32'h3c9eabb0, 32'h3e9b6490} /* (8, 12, 21) {real, imag} */,
  {32'hbeb42018, 32'hbf2e2721} /* (8, 12, 20) {real, imag} */,
  {32'hbe97baba, 32'h3e630d05} /* (8, 12, 19) {real, imag} */,
  {32'hbf0f969b, 32'h3e433a74} /* (8, 12, 18) {real, imag} */,
  {32'hbc056ee0, 32'h3e1df81c} /* (8, 12, 17) {real, imag} */,
  {32'hbdc11a54, 32'hbd24a7fb} /* (8, 12, 16) {real, imag} */,
  {32'hbc0e81a0, 32'hbeb70b26} /* (8, 12, 15) {real, imag} */,
  {32'hbdb2a3cf, 32'h3e84ae1c} /* (8, 12, 14) {real, imag} */,
  {32'hbf25fd20, 32'h3caeaa56} /* (8, 12, 13) {real, imag} */,
  {32'h3ee67d72, 32'hbe86a9d9} /* (8, 12, 12) {real, imag} */,
  {32'hbe0b7635, 32'hbe229e51} /* (8, 12, 11) {real, imag} */,
  {32'hbdbf40d0, 32'h3c68ac20} /* (8, 12, 10) {real, imag} */,
  {32'h3f02d65b, 32'hbe9e3488} /* (8, 12, 9) {real, imag} */,
  {32'hbdeaa95c, 32'h3f3cc3af} /* (8, 12, 8) {real, imag} */,
  {32'hbebc7917, 32'h3d9626de} /* (8, 12, 7) {real, imag} */,
  {32'h3e2c6c5d, 32'hbd3ea744} /* (8, 12, 6) {real, imag} */,
  {32'h3f331400, 32'h3ec98edf} /* (8, 12, 5) {real, imag} */,
  {32'hbe2bb416, 32'hbdbc0d68} /* (8, 12, 4) {real, imag} */,
  {32'h3e1690b5, 32'hbed008e3} /* (8, 12, 3) {real, imag} */,
  {32'hbe4f9ebc, 32'h3f044609} /* (8, 12, 2) {real, imag} */,
  {32'h3e964e44, 32'h3e2767df} /* (8, 12, 1) {real, imag} */,
  {32'h3e4dc9ca, 32'h3f24456d} /* (8, 12, 0) {real, imag} */,
  {32'h3e7dfe98, 32'h3da7f2ca} /* (8, 11, 31) {real, imag} */,
  {32'h3dfc0f6c, 32'h3ee03e2a} /* (8, 11, 30) {real, imag} */,
  {32'hbda49d82, 32'hbda3a120} /* (8, 11, 29) {real, imag} */,
  {32'h3e199a44, 32'h3eea3174} /* (8, 11, 28) {real, imag} */,
  {32'h3f241030, 32'h3d99b1ba} /* (8, 11, 27) {real, imag} */,
  {32'h3dd299e0, 32'hbe971ca4} /* (8, 11, 26) {real, imag} */,
  {32'hbe1a6464, 32'hbdeeb3aa} /* (8, 11, 25) {real, imag} */,
  {32'hbdf316e6, 32'hbd80e447} /* (8, 11, 24) {real, imag} */,
  {32'hbe162e51, 32'h3d1c200a} /* (8, 11, 23) {real, imag} */,
  {32'hbea809dd, 32'hbd880f88} /* (8, 11, 22) {real, imag} */,
  {32'h3e91e5b4, 32'hbea629f5} /* (8, 11, 21) {real, imag} */,
  {32'h3eee6cb2, 32'h3ea80ce9} /* (8, 11, 20) {real, imag} */,
  {32'h3d41f4f6, 32'hbe7666f6} /* (8, 11, 19) {real, imag} */,
  {32'hbc2e9c68, 32'hbe880698} /* (8, 11, 18) {real, imag} */,
  {32'h3c531500, 32'h3edb2730} /* (8, 11, 17) {real, imag} */,
  {32'h3cdf0d10, 32'hbe61f965} /* (8, 11, 16) {real, imag} */,
  {32'h3e0c9fca, 32'hbd1e3f94} /* (8, 11, 15) {real, imag} */,
  {32'h3df24476, 32'hbdc5c6de} /* (8, 11, 14) {real, imag} */,
  {32'hbf9a57ec, 32'h3e4217a2} /* (8, 11, 13) {real, imag} */,
  {32'hbebb9580, 32'hbe5529b4} /* (8, 11, 12) {real, imag} */,
  {32'h3ddaa7eb, 32'h3e361875} /* (8, 11, 11) {real, imag} */,
  {32'hbf2d1132, 32'h3f89808d} /* (8, 11, 10) {real, imag} */,
  {32'h3ed3a870, 32'hbcef63f0} /* (8, 11, 9) {real, imag} */,
  {32'hbed94768, 32'hbf023c90} /* (8, 11, 8) {real, imag} */,
  {32'hbe65c5c7, 32'hbe11e722} /* (8, 11, 7) {real, imag} */,
  {32'h3def1ea0, 32'h3d3ae576} /* (8, 11, 6) {real, imag} */,
  {32'hbf55675d, 32'hbdd1725d} /* (8, 11, 5) {real, imag} */,
  {32'h3ec05847, 32'hbda04283} /* (8, 11, 4) {real, imag} */,
  {32'hbd5b6708, 32'h3e85d7ee} /* (8, 11, 3) {real, imag} */,
  {32'h3e940654, 32'h3ea62ab4} /* (8, 11, 2) {real, imag} */,
  {32'hbdeffe40, 32'hbeedc1f0} /* (8, 11, 1) {real, imag} */,
  {32'hbf5e58f0, 32'hbf719ffb} /* (8, 11, 0) {real, imag} */,
  {32'h3c032b70, 32'hbd617bc8} /* (8, 10, 31) {real, imag} */,
  {32'hbea0172c, 32'hbd8884f8} /* (8, 10, 30) {real, imag} */,
  {32'hbbb5b3c0, 32'hbe1983d6} /* (8, 10, 29) {real, imag} */,
  {32'h3f29b56d, 32'hbd7b3d02} /* (8, 10, 28) {real, imag} */,
  {32'h3dd2d82c, 32'h3e69bf85} /* (8, 10, 27) {real, imag} */,
  {32'hbed3bc4d, 32'h3e4d4586} /* (8, 10, 26) {real, imag} */,
  {32'hbf0ec2d2, 32'hbdb72eea} /* (8, 10, 25) {real, imag} */,
  {32'hbe4067f1, 32'hbebb7f13} /* (8, 10, 24) {real, imag} */,
  {32'hbee86a9b, 32'hbe6e3314} /* (8, 10, 23) {real, imag} */,
  {32'hbd873572, 32'hbe2c138b} /* (8, 10, 22) {real, imag} */,
  {32'h3eaa4f8a, 32'h3e9e9dbc} /* (8, 10, 21) {real, imag} */,
  {32'h3e9d7941, 32'hbcbb224c} /* (8, 10, 20) {real, imag} */,
  {32'h3eb94fca, 32'h3e85d9a4} /* (8, 10, 19) {real, imag} */,
  {32'h3cf22020, 32'hbe00fdc8} /* (8, 10, 18) {real, imag} */,
  {32'h3e87b5ef, 32'hbddb90a8} /* (8, 10, 17) {real, imag} */,
  {32'hbe69f8aa, 32'h3dd1bed6} /* (8, 10, 16) {real, imag} */,
  {32'h3d47fd52, 32'h3e869a98} /* (8, 10, 15) {real, imag} */,
  {32'hbdc84b42, 32'hbddd3018} /* (8, 10, 14) {real, imag} */,
  {32'h3d935819, 32'h3eb23515} /* (8, 10, 13) {real, imag} */,
  {32'h3eae1097, 32'hbe173398} /* (8, 10, 12) {real, imag} */,
  {32'h3aa40b00, 32'h3e36ad7c} /* (8, 10, 11) {real, imag} */,
  {32'h3e13403a, 32'hbe75245a} /* (8, 10, 10) {real, imag} */,
  {32'h3f2562d9, 32'hbe4b6f1b} /* (8, 10, 9) {real, imag} */,
  {32'hbcfd9608, 32'h3e6d07b5} /* (8, 10, 8) {real, imag} */,
  {32'h3e4dfa1c, 32'hbe95ff91} /* (8, 10, 7) {real, imag} */,
  {32'hbf27dd91, 32'hbcabeaf8} /* (8, 10, 6) {real, imag} */,
  {32'hbec315e2, 32'hbdd06771} /* (8, 10, 5) {real, imag} */,
  {32'h3ebf70de, 32'h3e8ac131} /* (8, 10, 4) {real, imag} */,
  {32'hbebb5051, 32'h3cec78da} /* (8, 10, 3) {real, imag} */,
  {32'h3eca5af5, 32'h3e3fcc9a} /* (8, 10, 2) {real, imag} */,
  {32'hbe2d8c29, 32'hbdca7a20} /* (8, 10, 1) {real, imag} */,
  {32'hbe7a5f81, 32'h3e9d3b3a} /* (8, 10, 0) {real, imag} */,
  {32'hbf375939, 32'h3f2ed1db} /* (8, 9, 31) {real, imag} */,
  {32'h3f001be1, 32'hbf482d02} /* (8, 9, 30) {real, imag} */,
  {32'h3e440757, 32'h3ca37808} /* (8, 9, 29) {real, imag} */,
  {32'hbf1a9344, 32'hbcdea538} /* (8, 9, 28) {real, imag} */,
  {32'hbf0ff435, 32'hbd9502f0} /* (8, 9, 27) {real, imag} */,
  {32'hbdb22c92, 32'hbee73680} /* (8, 9, 26) {real, imag} */,
  {32'hbcf9a7f4, 32'hbf1895d0} /* (8, 9, 25) {real, imag} */,
  {32'hbe293a42, 32'h3e5e5bd6} /* (8, 9, 24) {real, imag} */,
  {32'hbcbd1fe0, 32'h3e7fe028} /* (8, 9, 23) {real, imag} */,
  {32'h3e9cdd0c, 32'hbe69511c} /* (8, 9, 22) {real, imag} */,
  {32'h3e3222a0, 32'h3f54de4c} /* (8, 9, 21) {real, imag} */,
  {32'h3eec6859, 32'h3e361877} /* (8, 9, 20) {real, imag} */,
  {32'hbe5363be, 32'hbe86977a} /* (8, 9, 19) {real, imag} */,
  {32'hbe651436, 32'h3dac8e8e} /* (8, 9, 18) {real, imag} */,
  {32'hbd9b7c33, 32'hbe0e8632} /* (8, 9, 17) {real, imag} */,
  {32'h3d82d384, 32'h3e3e27b1} /* (8, 9, 16) {real, imag} */,
  {32'hbe72c9bc, 32'h3ede0108} /* (8, 9, 15) {real, imag} */,
  {32'h3d3c5d70, 32'h3e85b13e} /* (8, 9, 14) {real, imag} */,
  {32'h3d2a1ac8, 32'hbef65ef1} /* (8, 9, 13) {real, imag} */,
  {32'h3f28f4ea, 32'hbec9c5c7} /* (8, 9, 12) {real, imag} */,
  {32'h3df5311c, 32'hbd420a96} /* (8, 9, 11) {real, imag} */,
  {32'hbe411e19, 32'h3e663bff} /* (8, 9, 10) {real, imag} */,
  {32'hbed3f2af, 32'h3f0018ce} /* (8, 9, 9) {real, imag} */,
  {32'hbe1b03f5, 32'hbc9a4628} /* (8, 9, 8) {real, imag} */,
  {32'hbe490e47, 32'h3e9f85ba} /* (8, 9, 7) {real, imag} */,
  {32'hbeb08120, 32'hbdc5997a} /* (8, 9, 6) {real, imag} */,
  {32'hbda27b2c, 32'hbe997c32} /* (8, 9, 5) {real, imag} */,
  {32'h3d95ba23, 32'h3e1322b6} /* (8, 9, 4) {real, imag} */,
  {32'hbd6fbaca, 32'hbe4fcd6b} /* (8, 9, 3) {real, imag} */,
  {32'hbdd7e46f, 32'hbf03bd80} /* (8, 9, 2) {real, imag} */,
  {32'h3e2e3e34, 32'h3d0722d4} /* (8, 9, 1) {real, imag} */,
  {32'hbf3f00d0, 32'hbf5687ce} /* (8, 9, 0) {real, imag} */,
  {32'hbfab588b, 32'hbf737c8e} /* (8, 8, 31) {real, imag} */,
  {32'h3f59f388, 32'hbdaf43d6} /* (8, 8, 30) {real, imag} */,
  {32'h3e0d2346, 32'h3d28f49a} /* (8, 8, 29) {real, imag} */,
  {32'h3f601a48, 32'hba1b8f80} /* (8, 8, 28) {real, imag} */,
  {32'h3ef5b960, 32'hbe836f92} /* (8, 8, 27) {real, imag} */,
  {32'h3f0e7085, 32'hbe212d66} /* (8, 8, 26) {real, imag} */,
  {32'hbdb4541c, 32'h3ed54ef3} /* (8, 8, 25) {real, imag} */,
  {32'hbcc3dca8, 32'hbef07c13} /* (8, 8, 24) {real, imag} */,
  {32'h3dcd317c, 32'hbe3db690} /* (8, 8, 23) {real, imag} */,
  {32'hbce0ae0b, 32'hbd3fc020} /* (8, 8, 22) {real, imag} */,
  {32'h3d2c2baa, 32'h3dbae2c4} /* (8, 8, 21) {real, imag} */,
  {32'h3dd5a426, 32'h3ef0035b} /* (8, 8, 20) {real, imag} */,
  {32'hbe5f9239, 32'hbdde8d58} /* (8, 8, 19) {real, imag} */,
  {32'hbe7facf9, 32'hbebd1d44} /* (8, 8, 18) {real, imag} */,
  {32'h3e437693, 32'h3ea8a6b2} /* (8, 8, 17) {real, imag} */,
  {32'h3e4ba8de, 32'h3e0ad055} /* (8, 8, 16) {real, imag} */,
  {32'hbc318a10, 32'h3dae8d62} /* (8, 8, 15) {real, imag} */,
  {32'hbed73482, 32'h3e675785} /* (8, 8, 14) {real, imag} */,
  {32'h3dad6963, 32'hbeacf958} /* (8, 8, 13) {real, imag} */,
  {32'h3ea00028, 32'hbc2488c8} /* (8, 8, 12) {real, imag} */,
  {32'h3e5910ca, 32'h3bd9d600} /* (8, 8, 11) {real, imag} */,
  {32'h3f0f8dbb, 32'h3e8ea5bd} /* (8, 8, 10) {real, imag} */,
  {32'h3b9893e0, 32'h3eb91f5d} /* (8, 8, 9) {real, imag} */,
  {32'hbe42fbc4, 32'hbece4b69} /* (8, 8, 8) {real, imag} */,
  {32'hbed2cfeb, 32'h3f40a1ed} /* (8, 8, 7) {real, imag} */,
  {32'hbd5327c0, 32'hbf15483c} /* (8, 8, 6) {real, imag} */,
  {32'h3e9cd322, 32'h3da01c7e} /* (8, 8, 5) {real, imag} */,
  {32'hbdefa31a, 32'hbf14aa26} /* (8, 8, 4) {real, imag} */,
  {32'h3d9ebc3c, 32'h3e9e50d4} /* (8, 8, 3) {real, imag} */,
  {32'h3f44b48c, 32'hbb6d9780} /* (8, 8, 2) {real, imag} */,
  {32'hbf471e19, 32'hbef5166e} /* (8, 8, 1) {real, imag} */,
  {32'hbf136038, 32'h3c9c9980} /* (8, 8, 0) {real, imag} */,
  {32'hbe147a74, 32'hbe66c954} /* (8, 7, 31) {real, imag} */,
  {32'h3c92f940, 32'hbee0713a} /* (8, 7, 30) {real, imag} */,
  {32'h3d8bb6b6, 32'hbe972242} /* (8, 7, 29) {real, imag} */,
  {32'hbe98ba23, 32'h3ed3e79f} /* (8, 7, 28) {real, imag} */,
  {32'hbe0e45ce, 32'h3bf4b720} /* (8, 7, 27) {real, imag} */,
  {32'h3e9c9b49, 32'hbe3fe0a8} /* (8, 7, 26) {real, imag} */,
  {32'hbe905f5e, 32'h3e3d15d5} /* (8, 7, 25) {real, imag} */,
  {32'h3dd272c6, 32'hbe54e389} /* (8, 7, 24) {real, imag} */,
  {32'hbee1dde2, 32'h3dd98f37} /* (8, 7, 23) {real, imag} */,
  {32'hbca0a856, 32'h3ecea660} /* (8, 7, 22) {real, imag} */,
  {32'hbd719858, 32'h3e1bf2a8} /* (8, 7, 21) {real, imag} */,
  {32'h3e85e7e7, 32'h3dd31ec0} /* (8, 7, 20) {real, imag} */,
  {32'h3e99e5c6, 32'hbdf9f117} /* (8, 7, 19) {real, imag} */,
  {32'h3ec22796, 32'hbeb62cdc} /* (8, 7, 18) {real, imag} */,
  {32'h3e00da92, 32'hbe412dcd} /* (8, 7, 17) {real, imag} */,
  {32'h3ddab75e, 32'hbc0c5a30} /* (8, 7, 16) {real, imag} */,
  {32'h3e578e06, 32'hbec94efe} /* (8, 7, 15) {real, imag} */,
  {32'h3ecf910f, 32'h3de10a3a} /* (8, 7, 14) {real, imag} */,
  {32'hbef3a30a, 32'h3d2b1194} /* (8, 7, 13) {real, imag} */,
  {32'hbec96cbe, 32'hbe5f5733} /* (8, 7, 12) {real, imag} */,
  {32'h3f0371a9, 32'h3dcc8b86} /* (8, 7, 11) {real, imag} */,
  {32'hbda04e30, 32'hbd38f2b0} /* (8, 7, 10) {real, imag} */,
  {32'hbe6091b0, 32'h3ef14b59} /* (8, 7, 9) {real, imag} */,
  {32'h3e6466f4, 32'h3eb6c616} /* (8, 7, 8) {real, imag} */,
  {32'h3e91d480, 32'hbe99ba82} /* (8, 7, 7) {real, imag} */,
  {32'hbe94a574, 32'hbe406b47} /* (8, 7, 6) {real, imag} */,
  {32'h3e8860d2, 32'h3e12faa6} /* (8, 7, 5) {real, imag} */,
  {32'hbec3ff04, 32'h3d24ccc9} /* (8, 7, 4) {real, imag} */,
  {32'hbf79ef90, 32'h3f4cd28a} /* (8, 7, 3) {real, imag} */,
  {32'hbd3a0994, 32'hbf9b4ef0} /* (8, 7, 2) {real, imag} */,
  {32'h3ec7b797, 32'h3f4725cf} /* (8, 7, 1) {real, imag} */,
  {32'h3f1f600c, 32'h3e8ba742} /* (8, 7, 0) {real, imag} */,
  {32'hbe93337e, 32'hbe9d0403} /* (8, 6, 31) {real, imag} */,
  {32'hbba23fc0, 32'h3dca774a} /* (8, 6, 30) {real, imag} */,
  {32'h3dc391bc, 32'h3e519c6e} /* (8, 6, 29) {real, imag} */,
  {32'hbdab32e4, 32'hbe7af4b7} /* (8, 6, 28) {real, imag} */,
  {32'h3ea55606, 32'h3f027fcf} /* (8, 6, 27) {real, imag} */,
  {32'hbed96dca, 32'h3ece255c} /* (8, 6, 26) {real, imag} */,
  {32'h3c039ff8, 32'h3d86ad42} /* (8, 6, 25) {real, imag} */,
  {32'h3c2c5cd8, 32'hbe322f40} /* (8, 6, 24) {real, imag} */,
  {32'h3f0d37be, 32'h3ec6f048} /* (8, 6, 23) {real, imag} */,
  {32'h3eedb58a, 32'hbdfae31e} /* (8, 6, 22) {real, imag} */,
  {32'h3eb8a24b, 32'hbce2e78c} /* (8, 6, 21) {real, imag} */,
  {32'hbf1c9498, 32'hbf3a7193} /* (8, 6, 20) {real, imag} */,
  {32'hbe0cda54, 32'h3ead1013} /* (8, 6, 19) {real, imag} */,
  {32'h3e814c70, 32'hbea81e2f} /* (8, 6, 18) {real, imag} */,
  {32'h3e01d552, 32'hbe82b2b7} /* (8, 6, 17) {real, imag} */,
  {32'hbe5fc13c, 32'hbdc6a443} /* (8, 6, 16) {real, imag} */,
  {32'h3e1cd784, 32'hbe733dc2} /* (8, 6, 15) {real, imag} */,
  {32'h3e83ab2e, 32'h3dabbf04} /* (8, 6, 14) {real, imag} */,
  {32'h3eac16ae, 32'hbe01eea8} /* (8, 6, 13) {real, imag} */,
  {32'h3e866f9f, 32'h3e95083d} /* (8, 6, 12) {real, imag} */,
  {32'h3ec53715, 32'hbef3b089} /* (8, 6, 11) {real, imag} */,
  {32'h3eec69ea, 32'h3e90c792} /* (8, 6, 10) {real, imag} */,
  {32'hbe7e0c32, 32'h3ce2edb8} /* (8, 6, 9) {real, imag} */,
  {32'h3db17a9a, 32'h3e67cab1} /* (8, 6, 8) {real, imag} */,
  {32'hbe878555, 32'h3f932adc} /* (8, 6, 7) {real, imag} */,
  {32'h3ea525d6, 32'h3e902f8f} /* (8, 6, 6) {real, imag} */,
  {32'h3d8b4c4c, 32'hbe12a7a7} /* (8, 6, 5) {real, imag} */,
  {32'h3ef29525, 32'hbecf2690} /* (8, 6, 4) {real, imag} */,
  {32'h3e0c642c, 32'h3e2a9c49} /* (8, 6, 3) {real, imag} */,
  {32'hbf826050, 32'hbee3b8b4} /* (8, 6, 2) {real, imag} */,
  {32'hbec1a9e0, 32'hbec0adb2} /* (8, 6, 1) {real, imag} */,
  {32'hbea8f784, 32'h3eed50a2} /* (8, 6, 0) {real, imag} */,
  {32'hc0245f32, 32'hbea68117} /* (8, 5, 31) {real, imag} */,
  {32'h3f939c8f, 32'hbf4f5082} /* (8, 5, 30) {real, imag} */,
  {32'h3f396cb6, 32'h3ddccd84} /* (8, 5, 29) {real, imag} */,
  {32'h3d6c1680, 32'hbe327da9} /* (8, 5, 28) {real, imag} */,
  {32'hbe2f85c8, 32'hbe5c86c0} /* (8, 5, 27) {real, imag} */,
  {32'hbeffec05, 32'h3f6cd200} /* (8, 5, 26) {real, imag} */,
  {32'h3dc812b8, 32'h3eb77a2e} /* (8, 5, 25) {real, imag} */,
  {32'h3ee75f10, 32'hbf1b53a4} /* (8, 5, 24) {real, imag} */,
  {32'hbcd9211c, 32'h3eaf0302} /* (8, 5, 23) {real, imag} */,
  {32'h3e846867, 32'hbd5b52a8} /* (8, 5, 22) {real, imag} */,
  {32'h3c91f7f0, 32'hbf2f835c} /* (8, 5, 21) {real, imag} */,
  {32'hbeb5eb5a, 32'hbec210f2} /* (8, 5, 20) {real, imag} */,
  {32'h3e947cb8, 32'h3e42c4a4} /* (8, 5, 19) {real, imag} */,
  {32'hbe7480f6, 32'hbddd50da} /* (8, 5, 18) {real, imag} */,
  {32'hbe21ecfa, 32'hbda0f380} /* (8, 5, 17) {real, imag} */,
  {32'h3e8314b3, 32'h3da63d22} /* (8, 5, 16) {real, imag} */,
  {32'h3ecca738, 32'h3d0f37a4} /* (8, 5, 15) {real, imag} */,
  {32'hbea746a6, 32'h3f327688} /* (8, 5, 14) {real, imag} */,
  {32'hbe84c9f6, 32'h3dec48ec} /* (8, 5, 13) {real, imag} */,
  {32'h3ea1277a, 32'hbe5823c2} /* (8, 5, 12) {real, imag} */,
  {32'h3e9b0683, 32'hbf171048} /* (8, 5, 11) {real, imag} */,
  {32'h3e6158e9, 32'h3d82028c} /* (8, 5, 10) {real, imag} */,
  {32'hbdcd9140, 32'h3e97b90d} /* (8, 5, 9) {real, imag} */,
  {32'h3f156503, 32'hbe0601c4} /* (8, 5, 8) {real, imag} */,
  {32'hbeb47a94, 32'hbe9fbe62} /* (8, 5, 7) {real, imag} */,
  {32'hbdd0a0d8, 32'h3ed5a3bd} /* (8, 5, 6) {real, imag} */,
  {32'h3fc1590c, 32'h3f8f191d} /* (8, 5, 5) {real, imag} */,
  {32'hbf19a4ea, 32'hbe910346} /* (8, 5, 4) {real, imag} */,
  {32'hbeff891e, 32'hbc50c570} /* (8, 5, 3) {real, imag} */,
  {32'h3f44c139, 32'h3fb5c15c} /* (8, 5, 2) {real, imag} */,
  {32'hbf61dd3a, 32'hc0003406} /* (8, 5, 1) {real, imag} */,
  {32'hc005626f, 32'hbf2f64cd} /* (8, 5, 0) {real, imag} */,
  {32'h3f4d1bda, 32'h4043a0d8} /* (8, 4, 31) {real, imag} */,
  {32'hc02c3a41, 32'hc0230b6d} /* (8, 4, 30) {real, imag} */,
  {32'hbf3d52fa, 32'hbe21fec8} /* (8, 4, 29) {real, imag} */,
  {32'h3f3762c1, 32'h3f13291a} /* (8, 4, 28) {real, imag} */,
  {32'hbf0e30f6, 32'hbef5b074} /* (8, 4, 27) {real, imag} */,
  {32'hbe82be28, 32'h3e89bfce} /* (8, 4, 26) {real, imag} */,
  {32'h3e79daf2, 32'h3e5571dc} /* (8, 4, 25) {real, imag} */,
  {32'hbea66fa4, 32'hbedf1371} /* (8, 4, 24) {real, imag} */,
  {32'h3f34e8f0, 32'hbe03a134} /* (8, 4, 23) {real, imag} */,
  {32'h3ebc69c6, 32'hbee94c04} /* (8, 4, 22) {real, imag} */,
  {32'hbd05bf0c, 32'h3ee22b63} /* (8, 4, 21) {real, imag} */,
  {32'h3de4a5ae, 32'h3e0acd0c} /* (8, 4, 20) {real, imag} */,
  {32'hbdcf186e, 32'h3df59e8d} /* (8, 4, 19) {real, imag} */,
  {32'h3cf887d8, 32'hbec984c5} /* (8, 4, 18) {real, imag} */,
  {32'hbe896498, 32'hbc520fe0} /* (8, 4, 17) {real, imag} */,
  {32'h3ec18759, 32'hbcec4b78} /* (8, 4, 16) {real, imag} */,
  {32'hbe57fe1a, 32'hbe8b5554} /* (8, 4, 15) {real, imag} */,
  {32'h3e50ba30, 32'hbe9b4534} /* (8, 4, 14) {real, imag} */,
  {32'hbc1c3290, 32'h3f27fdbe} /* (8, 4, 13) {real, imag} */,
  {32'h3d232af4, 32'h3ddb2d12} /* (8, 4, 12) {real, imag} */,
  {32'h3f14bde1, 32'h3df2f5fa} /* (8, 4, 11) {real, imag} */,
  {32'hbe99e39d, 32'h3e1558cb} /* (8, 4, 10) {real, imag} */,
  {32'hbe50dfe5, 32'h3e11c0a3} /* (8, 4, 9) {real, imag} */,
  {32'h3ec8bd09, 32'hbfa4d9bc} /* (8, 4, 8) {real, imag} */,
  {32'h3e12b5da, 32'hbd54d568} /* (8, 4, 7) {real, imag} */,
  {32'h3f762477, 32'hbde4245c} /* (8, 4, 6) {real, imag} */,
  {32'hbdf3e91d, 32'hbf9139ed} /* (8, 4, 5) {real, imag} */,
  {32'h3ee00eac, 32'h3dcf0ee8} /* (8, 4, 4) {real, imag} */,
  {32'hbfbf514c, 32'h3f6f7074} /* (8, 4, 3) {real, imag} */,
  {32'hc052d024, 32'hc00dc6d8} /* (8, 4, 2) {real, imag} */,
  {32'h409b5363, 32'h400fdba4} /* (8, 4, 1) {real, imag} */,
  {32'h3fdcba62, 32'h3f4b1984} /* (8, 4, 0) {real, imag} */,
  {32'hc0893e46, 32'h3fb626fc} /* (8, 3, 31) {real, imag} */,
  {32'h40094744, 32'hc0990739} /* (8, 3, 30) {real, imag} */,
  {32'h3e94dccb, 32'h3f8a6de0} /* (8, 3, 29) {real, imag} */,
  {32'h3f86a215, 32'h3e300a0c} /* (8, 3, 28) {real, imag} */,
  {32'hbfac0982, 32'hbe453252} /* (8, 3, 27) {real, imag} */,
  {32'hbeb77f2f, 32'h3d34a574} /* (8, 3, 26) {real, imag} */,
  {32'hbf45f9d7, 32'h3f33ce37} /* (8, 3, 25) {real, imag} */,
  {32'hbf419c86, 32'hbf5ee8f4} /* (8, 3, 24) {real, imag} */,
  {32'h3c73f120, 32'hbe920a8a} /* (8, 3, 23) {real, imag} */,
  {32'h3f3014cf, 32'h3e94608e} /* (8, 3, 22) {real, imag} */,
  {32'h3d1272ea, 32'h3e907c32} /* (8, 3, 21) {real, imag} */,
  {32'h3e34b810, 32'h3d8f69e6} /* (8, 3, 20) {real, imag} */,
  {32'h3ec214fb, 32'h3f075f48} /* (8, 3, 19) {real, imag} */,
  {32'hbe4bf336, 32'hbe99a022} /* (8, 3, 18) {real, imag} */,
  {32'h3e817329, 32'hbb850ff0} /* (8, 3, 17) {real, imag} */,
  {32'hbeef6542, 32'h3ea959d7} /* (8, 3, 16) {real, imag} */,
  {32'hbf0d1aa0, 32'h3dda01d8} /* (8, 3, 15) {real, imag} */,
  {32'hbdf2e101, 32'hbeaa0b76} /* (8, 3, 14) {real, imag} */,
  {32'hbdbae50c, 32'hbdc08295} /* (8, 3, 13) {real, imag} */,
  {32'h3ebe90cb, 32'hbdd27004} /* (8, 3, 12) {real, imag} */,
  {32'h3e4fac72, 32'hbdef0eaf} /* (8, 3, 11) {real, imag} */,
  {32'hbe8ab030, 32'h3c674d38} /* (8, 3, 10) {real, imag} */,
  {32'h3c975ec0, 32'h3e2d7edd} /* (8, 3, 9) {real, imag} */,
  {32'h3dd39718, 32'h3ed7fcbc} /* (8, 3, 8) {real, imag} */,
  {32'hbf4471b5, 32'h3db48a10} /* (8, 3, 7) {real, imag} */,
  {32'hbe6275de, 32'h3df2ee5c} /* (8, 3, 6) {real, imag} */,
  {32'h3e84af16, 32'h3f57e300} /* (8, 3, 5) {real, imag} */,
  {32'hbfda96f3, 32'h3f4322c6} /* (8, 3, 4) {real, imag} */,
  {32'hbf1fe610, 32'h3e896a58} /* (8, 3, 3) {real, imag} */,
  {32'h3e888d04, 32'hc02fbae0} /* (8, 3, 2) {real, imag} */,
  {32'h40635e97, 32'h404fbbd8} /* (8, 3, 1) {real, imag} */,
  {32'h3f0dfd16, 32'hbf884645} /* (8, 3, 0) {real, imag} */,
  {32'hc218727c, 32'hbf7fb2f2} /* (8, 2, 31) {real, imag} */,
  {32'h418a3d64, 32'hc099eda6} /* (8, 2, 30) {real, imag} */,
  {32'hbf7b0fdb, 32'h40120442} /* (8, 2, 29) {real, imag} */,
  {32'hbf7f7fdc, 32'h400ed330} /* (8, 2, 28) {real, imag} */,
  {32'h402003a0, 32'hbf9caf60} /* (8, 2, 27) {real, imag} */,
  {32'h3f26cd38, 32'hbebf15dd} /* (8, 2, 26) {real, imag} */,
  {32'h3f37d1e8, 32'h3efe53be} /* (8, 2, 25) {real, imag} */,
  {32'h3f158887, 32'h3a8cca00} /* (8, 2, 24) {real, imag} */,
  {32'hbe8e917f, 32'hbd9d929a} /* (8, 2, 23) {real, imag} */,
  {32'hbe952825, 32'hbdeb0078} /* (8, 2, 22) {real, imag} */,
  {32'hbe87f4f8, 32'hbe7c9800} /* (8, 2, 21) {real, imag} */,
  {32'h3ef8535d, 32'hbf4f1b82} /* (8, 2, 20) {real, imag} */,
  {32'h3c8e9734, 32'hbeb0bbed} /* (8, 2, 19) {real, imag} */,
  {32'hbe9a609b, 32'hbc283950} /* (8, 2, 18) {real, imag} */,
  {32'h3f0739ba, 32'h3e9d214c} /* (8, 2, 17) {real, imag} */,
  {32'hbea1e42e, 32'h3e9acf0c} /* (8, 2, 16) {real, imag} */,
  {32'hbec8bf24, 32'h3e57b4b5} /* (8, 2, 15) {real, imag} */,
  {32'hbe7ced45, 32'h3e875247} /* (8, 2, 14) {real, imag} */,
  {32'h3e9e21f4, 32'hbe613645} /* (8, 2, 13) {real, imag} */,
  {32'h3ed3a7cb, 32'hbeb1c74c} /* (8, 2, 12) {real, imag} */,
  {32'hbd5a6a86, 32'h3ed848fc} /* (8, 2, 11) {real, imag} */,
  {32'hbe3bccc2, 32'hbce216b0} /* (8, 2, 10) {real, imag} */,
  {32'h3eec9750, 32'h3e619701} /* (8, 2, 9) {real, imag} */,
  {32'hbe0f4426, 32'h3d818f42} /* (8, 2, 8) {real, imag} */,
  {32'hbf10a884, 32'hbf839adc} /* (8, 2, 7) {real, imag} */,
  {32'h3d642078, 32'h3e60be35} /* (8, 2, 6) {real, imag} */,
  {32'h400c6076, 32'h3f5bbdea} /* (8, 2, 5) {real, imag} */,
  {32'hc05758c2, 32'hbf43bede} /* (8, 2, 4) {real, imag} */,
  {32'hbf650215, 32'h3de02560} /* (8, 2, 3) {real, imag} */,
  {32'h414ce94e, 32'hc02d8e00} /* (8, 2, 2) {real, imag} */,
  {32'hc1a03dbc, 32'h40a12c7c} /* (8, 2, 1) {real, imag} */,
  {32'hc19b20e7, 32'hc0958d32} /* (8, 2, 0) {real, imag} */,
  {32'h4243e72d, 32'hc146ca94} /* (8, 1, 31) {real, imag} */,
  {32'hc12b8065, 32'h40169374} /* (8, 1, 30) {real, imag} */,
  {32'hbe80a106, 32'hbe7e2978} /* (8, 1, 29) {real, imag} */,
  {32'h400394cd, 32'h40207ef2} /* (8, 1, 28) {real, imag} */,
  {32'hc035cc2c, 32'hbea3a32d} /* (8, 1, 27) {real, imag} */,
  {32'hbf1807b8, 32'h3eaed425} /* (8, 1, 26) {real, imag} */,
  {32'h3f15d823, 32'hbedcee22} /* (8, 1, 25) {real, imag} */,
  {32'hbf91bc7d, 32'hbc224140} /* (8, 1, 24) {real, imag} */,
  {32'h3e133ae0, 32'h3edd209e} /* (8, 1, 23) {real, imag} */,
  {32'h3d8cc0b8, 32'h3e5bd85f} /* (8, 1, 22) {real, imag} */,
  {32'hbfae581e, 32'h3e49eff2} /* (8, 1, 21) {real, imag} */,
  {32'h3ece6234, 32'hbf220ee9} /* (8, 1, 20) {real, imag} */,
  {32'hbdbc7b21, 32'hbe1ef37c} /* (8, 1, 19) {real, imag} */,
  {32'hbeaa4c87, 32'h3f189ca2} /* (8, 1, 18) {real, imag} */,
  {32'hbd9f94a6, 32'h3cb1bf3c} /* (8, 1, 17) {real, imag} */,
  {32'h3e1f1e63, 32'h3cf7e51e} /* (8, 1, 16) {real, imag} */,
  {32'h3e07c8b9, 32'h3e9b5098} /* (8, 1, 15) {real, imag} */,
  {32'h3e6556b2, 32'hbf0606e2} /* (8, 1, 14) {real, imag} */,
  {32'h3de70ff6, 32'hbd0e4e50} /* (8, 1, 13) {real, imag} */,
  {32'h3d3e162c, 32'hbf1ccdf0} /* (8, 1, 12) {real, imag} */,
  {32'hbe914d2c, 32'hbf2ec71a} /* (8, 1, 11) {real, imag} */,
  {32'hbf3db8a6, 32'hbe4da082} /* (8, 1, 10) {real, imag} */,
  {32'hbe89eb2a, 32'hbf0b9a8a} /* (8, 1, 9) {real, imag} */,
  {32'hbd9f0128, 32'hbf699d99} /* (8, 1, 8) {real, imag} */,
  {32'h3eae5da6, 32'h3ec9af36} /* (8, 1, 7) {real, imag} */,
  {32'hbf56180e, 32'hbde9fab4} /* (8, 1, 6) {real, imag} */,
  {32'hc01f7400, 32'hbf26fb00} /* (8, 1, 5) {real, imag} */,
  {32'h3fe99c56, 32'hbf035cb3} /* (8, 1, 4) {real, imag} */,
  {32'hbf9060a1, 32'hbfc35b96} /* (8, 1, 3) {real, imag} */,
  {32'hc18af8a8, 32'hc181b2e0} /* (8, 1, 2) {real, imag} */,
  {32'h428bb595, 32'h420a3849} /* (8, 1, 1) {real, imag} */,
  {32'h4284ce84, 32'h40e653ae} /* (8, 1, 0) {real, imag} */,
  {32'h42204da9, 32'hc2055672} /* (8, 0, 31) {real, imag} */,
  {32'hc0adcf1c, 32'h41232011} /* (8, 0, 30) {real, imag} */,
  {32'hbe86b557, 32'h3e1f5e94} /* (8, 0, 29) {real, imag} */,
  {32'hbe4079a0, 32'h3f589bdf} /* (8, 0, 28) {real, imag} */,
  {32'hc00e92c8, 32'h3e2aefa2} /* (8, 0, 27) {real, imag} */,
  {32'h3f7e832a, 32'hbeefa759} /* (8, 0, 26) {real, imag} */,
  {32'hbe9fa627, 32'hbf156852} /* (8, 0, 25) {real, imag} */,
  {32'h3f3dd5ec, 32'h3f5fd780} /* (8, 0, 24) {real, imag} */,
  {32'h3e818c46, 32'hbd0a9a0c} /* (8, 0, 23) {real, imag} */,
  {32'hbd15a502, 32'h3f361edd} /* (8, 0, 22) {real, imag} */,
  {32'hbf023ac5, 32'h3df8373c} /* (8, 0, 21) {real, imag} */,
  {32'hbeb4a3e7, 32'hbf447486} /* (8, 0, 20) {real, imag} */,
  {32'h3ed03e82, 32'hbde662b8} /* (8, 0, 19) {real, imag} */,
  {32'hbe1536d3, 32'h3e30edf6} /* (8, 0, 18) {real, imag} */,
  {32'hbe949894, 32'h3b6ed660} /* (8, 0, 17) {real, imag} */,
  {32'hbea70673, 32'h00000000} /* (8, 0, 16) {real, imag} */,
  {32'hbe949894, 32'hbb6ed660} /* (8, 0, 15) {real, imag} */,
  {32'hbe1536d3, 32'hbe30edf6} /* (8, 0, 14) {real, imag} */,
  {32'h3ed03e82, 32'h3de662b8} /* (8, 0, 13) {real, imag} */,
  {32'hbeb4a3e7, 32'h3f447486} /* (8, 0, 12) {real, imag} */,
  {32'hbf023ac5, 32'hbdf8373c} /* (8, 0, 11) {real, imag} */,
  {32'hbd15a502, 32'hbf361edd} /* (8, 0, 10) {real, imag} */,
  {32'h3e818c46, 32'h3d0a9a0c} /* (8, 0, 9) {real, imag} */,
  {32'h3f3dd5ec, 32'hbf5fd780} /* (8, 0, 8) {real, imag} */,
  {32'hbe9fa627, 32'h3f156852} /* (8, 0, 7) {real, imag} */,
  {32'h3f7e832a, 32'h3eefa759} /* (8, 0, 6) {real, imag} */,
  {32'hc00e92c8, 32'hbe2aefa2} /* (8, 0, 5) {real, imag} */,
  {32'hbe4079a0, 32'hbf589bdf} /* (8, 0, 4) {real, imag} */,
  {32'hbe86b557, 32'hbe1f5e94} /* (8, 0, 3) {real, imag} */,
  {32'hc0adcf1c, 32'hc1232011} /* (8, 0, 2) {real, imag} */,
  {32'h42204da9, 32'h42055672} /* (8, 0, 1) {real, imag} */,
  {32'h4289bc66, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h42646005, 32'hc1dac369} /* (7, 31, 31) {real, imag} */,
  {32'hc1686dfe, 32'h4166db87} /* (7, 31, 30) {real, imag} */,
  {32'hbfb3fe73, 32'h403ea9b8} /* (7, 31, 29) {real, imag} */,
  {32'h3fc5eefc, 32'h3ed82628} /* (7, 31, 28) {real, imag} */,
  {32'hc0147832, 32'h3f851748} /* (7, 31, 27) {real, imag} */,
  {32'hbf2184f3, 32'h3d6e1918} /* (7, 31, 26) {real, imag} */,
  {32'h3f046d3d, 32'hbf2afaa4} /* (7, 31, 25) {real, imag} */,
  {32'hbee5b8e3, 32'h3fa474f4} /* (7, 31, 24) {real, imag} */,
  {32'hbe8ef8eb, 32'hbd7e84c2} /* (7, 31, 23) {real, imag} */,
  {32'hbe231a3c, 32'hbea874cf} /* (7, 31, 22) {real, imag} */,
  {32'hbf0baf35, 32'h3ef3dd65} /* (7, 31, 21) {real, imag} */,
  {32'h3d1a5122, 32'h3e9f9a44} /* (7, 31, 20) {real, imag} */,
  {32'hbebeed78, 32'h3eac31bb} /* (7, 31, 19) {real, imag} */,
  {32'hbe9d4807, 32'hbdcd7a80} /* (7, 31, 18) {real, imag} */,
  {32'hbdd8398b, 32'hbe70c7a2} /* (7, 31, 17) {real, imag} */,
  {32'hbc730e68, 32'h3f094ed0} /* (7, 31, 16) {real, imag} */,
  {32'hbe6c9447, 32'hbc2b8dd8} /* (7, 31, 15) {real, imag} */,
  {32'h3d0eb8f4, 32'hbf294be0} /* (7, 31, 14) {real, imag} */,
  {32'h3da5fd46, 32'hbe839e28} /* (7, 31, 13) {real, imag} */,
  {32'h3c943e00, 32'hbe0934b4} /* (7, 31, 12) {real, imag} */,
  {32'hbe97b321, 32'hbf74c342} /* (7, 31, 11) {real, imag} */,
  {32'h3f1bf955, 32'h3e10a892} /* (7, 31, 10) {real, imag} */,
  {32'h3e23d984, 32'hbe770729} /* (7, 31, 9) {real, imag} */,
  {32'hbf45bb0f, 32'hbf4386b2} /* (7, 31, 8) {real, imag} */,
  {32'h3e941749, 32'h3dd14667} /* (7, 31, 7) {real, imag} */,
  {32'hbf18a781, 32'hbf66c1b7} /* (7, 31, 6) {real, imag} */,
  {32'hc03cfb34, 32'hbccd7808} /* (7, 31, 5) {real, imag} */,
  {32'h3fd2bdee, 32'hc00425f4} /* (7, 31, 4) {real, imag} */,
  {32'h3fb125cc, 32'h3f9fd7f0} /* (7, 31, 3) {real, imag} */,
  {32'hc109f35d, 32'hbf981785} /* (7, 31, 2) {real, imag} */,
  {32'h4224cfda, 32'h412909f4} /* (7, 31, 1) {real, imag} */,
  {32'h425eaf4e, 32'hc0e99daf} /* (7, 31, 0) {real, imag} */,
  {32'hc181a06e, 32'hc0400cee} /* (7, 30, 31) {real, imag} */,
  {32'h413fb028, 32'h3fd2eee3} /* (7, 30, 30) {real, imag} */,
  {32'hbf6510e5, 32'hbf86f27a} /* (7, 30, 29) {real, imag} */,
  {32'hc06d82c2, 32'h3f245c96} /* (7, 30, 28) {real, imag} */,
  {32'h3fda86e0, 32'hbf90dd2d} /* (7, 30, 27) {real, imag} */,
  {32'h3e94d677, 32'hbd1d75c8} /* (7, 30, 26) {real, imag} */,
  {32'hbe546ab6, 32'h3f2bb5e4} /* (7, 30, 25) {real, imag} */,
  {32'hbdca8438, 32'hbe66ec32} /* (7, 30, 24) {real, imag} */,
  {32'h3e7dfff3, 32'hbf2d5409} /* (7, 30, 23) {real, imag} */,
  {32'h3e9e3bfc, 32'hbc12d3a0} /* (7, 30, 22) {real, imag} */,
  {32'h3ef320d2, 32'hbec73896} /* (7, 30, 21) {real, imag} */,
  {32'hbf046e42, 32'hbeabe0dc} /* (7, 30, 20) {real, imag} */,
  {32'hbf0bbdb3, 32'h3cc94fd0} /* (7, 30, 19) {real, imag} */,
  {32'h3e8ca669, 32'h3e902aaf} /* (7, 30, 18) {real, imag} */,
  {32'h3ea490e8, 32'hbe522017} /* (7, 30, 17) {real, imag} */,
  {32'hbdd779f8, 32'hbdf4dd6a} /* (7, 30, 16) {real, imag} */,
  {32'hbb200920, 32'hbd342c24} /* (7, 30, 15) {real, imag} */,
  {32'h3da5f04c, 32'h3e7a5f60} /* (7, 30, 14) {real, imag} */,
  {32'hbe17bc02, 32'hbc8d77c0} /* (7, 30, 13) {real, imag} */,
  {32'h3f013f15, 32'h3f0553c3} /* (7, 30, 12) {real, imag} */,
  {32'h3f067f99, 32'h3e0ce1fb} /* (7, 30, 11) {real, imag} */,
  {32'h3f2d37ac, 32'hbf312e16} /* (7, 30, 10) {real, imag} */,
  {32'h3e6886ca, 32'h3e244ae9} /* (7, 30, 9) {real, imag} */,
  {32'h3f7d0b22, 32'hbe8b4666} /* (7, 30, 8) {real, imag} */,
  {32'hbf1e8dac, 32'hbdee44a0} /* (7, 30, 7) {real, imag} */,
  {32'h3f17941f, 32'h3eb919e7} /* (7, 30, 6) {real, imag} */,
  {32'h3fb5edfc, 32'h3f969f3e} /* (7, 30, 5) {real, imag} */,
  {32'hbe3c7818, 32'hbfa50f79} /* (7, 30, 4) {real, imag} */,
  {32'hbfc1ec25, 32'hbfc9bce9} /* (7, 30, 3) {real, imag} */,
  {32'h41744116, 32'h40849647} /* (7, 30, 2) {real, imag} */,
  {32'hc1fc0336, 32'hbf08d424} /* (7, 30, 1) {real, imag} */,
  {32'hc1820d36, 32'h40b5fa66} /* (7, 30, 0) {real, imag} */,
  {32'h40843c7c, 32'hc0857b78} /* (7, 29, 31) {real, imag} */,
  {32'hbf29105c, 32'h3fe1f7be} /* (7, 29, 30) {real, imag} */,
  {32'hbe2802b7, 32'h3e8ff03a} /* (7, 29, 29) {real, imag} */,
  {32'hbfc3bbb3, 32'hbf362de3} /* (7, 29, 28) {real, imag} */,
  {32'h3f7de1fa, 32'h3e1b275c} /* (7, 29, 27) {real, imag} */,
  {32'h3da4ca54, 32'h3eae0949} /* (7, 29, 26) {real, imag} */,
  {32'hbde4a047, 32'hbe1ebce2} /* (7, 29, 25) {real, imag} */,
  {32'hbe1f597f, 32'hbea916c2} /* (7, 29, 24) {real, imag} */,
  {32'h3e5684a1, 32'hbeef3847} /* (7, 29, 23) {real, imag} */,
  {32'hbd38eaf2, 32'h3d520ec0} /* (7, 29, 22) {real, imag} */,
  {32'hbe437236, 32'h3f24e890} /* (7, 29, 21) {real, imag} */,
  {32'h3cddf110, 32'h3ee98afb} /* (7, 29, 20) {real, imag} */,
  {32'hbe44cb0a, 32'h3ddc5322} /* (7, 29, 19) {real, imag} */,
  {32'h3ef04e0a, 32'hbe9f7362} /* (7, 29, 18) {real, imag} */,
  {32'h3dcc3cc8, 32'hbe0c597a} /* (7, 29, 17) {real, imag} */,
  {32'h3d1c0f3c, 32'h3eb20dcc} /* (7, 29, 16) {real, imag} */,
  {32'hbdace640, 32'hbbd2f7e0} /* (7, 29, 15) {real, imag} */,
  {32'h3c3af8d0, 32'h3e7f8842} /* (7, 29, 14) {real, imag} */,
  {32'h3f0b3650, 32'hbe3e71e4} /* (7, 29, 13) {real, imag} */,
  {32'hbeac9c55, 32'h3df810d4} /* (7, 29, 12) {real, imag} */,
  {32'h3dd3417b, 32'h3f0785b6} /* (7, 29, 11) {real, imag} */,
  {32'h3c2d01e8, 32'hbdda4ed5} /* (7, 29, 10) {real, imag} */,
  {32'h3d560968, 32'hbb4c3340} /* (7, 29, 9) {real, imag} */,
  {32'hbf37a790, 32'h3f337252} /* (7, 29, 8) {real, imag} */,
  {32'hbf40829c, 32'hbf18d497} /* (7, 29, 7) {real, imag} */,
  {32'hbf3852fa, 32'h3db55df0} /* (7, 29, 6) {real, imag} */,
  {32'hbdd8e7a2, 32'hbe8c36d4} /* (7, 29, 5) {real, imag} */,
  {32'h3fa71c10, 32'hbf4aaf40} /* (7, 29, 4) {real, imag} */,
  {32'hbee905a8, 32'h3d08cbd0} /* (7, 29, 3) {real, imag} */,
  {32'h3ff0769c, 32'h406ccdb2} /* (7, 29, 2) {real, imag} */,
  {32'hc08efc8b, 32'hbfdd5adc} /* (7, 29, 1) {real, imag} */,
  {32'h3f32150d, 32'hbe87d89d} /* (7, 29, 0) {real, imag} */,
  {32'h407063b8, 32'hc0457a32} /* (7, 28, 31) {real, imag} */,
  {32'hc0190dcb, 32'h402b1fba} /* (7, 28, 30) {real, imag} */,
  {32'hbf05c3a1, 32'h3d2f91d4} /* (7, 28, 29) {real, imag} */,
  {32'h3e6be8f6, 32'hbfa712dd} /* (7, 28, 28) {real, imag} */,
  {32'hbcdedd60, 32'h3f91f9ac} /* (7, 28, 27) {real, imag} */,
  {32'h3e830cb3, 32'hbeac2d98} /* (7, 28, 26) {real, imag} */,
  {32'hbd7fc7d0, 32'hbc8f5dc0} /* (7, 28, 25) {real, imag} */,
  {32'hbe66e362, 32'h3f168b22} /* (7, 28, 24) {real, imag} */,
  {32'h3ee88ac6, 32'h3f29b961} /* (7, 28, 23) {real, imag} */,
  {32'h3de7b9ff, 32'h3d283df4} /* (7, 28, 22) {real, imag} */,
  {32'h3e746279, 32'h3efabb78} /* (7, 28, 21) {real, imag} */,
  {32'hbe6c5af8, 32'hbe4475a4} /* (7, 28, 20) {real, imag} */,
  {32'h3ee76cc0, 32'hbde738e8} /* (7, 28, 19) {real, imag} */,
  {32'hbef5f890, 32'h3e41ae46} /* (7, 28, 18) {real, imag} */,
  {32'hbed00cd0, 32'hbe4ed7ab} /* (7, 28, 17) {real, imag} */,
  {32'h3c32f91e, 32'hbe4e1870} /* (7, 28, 16) {real, imag} */,
  {32'h3ebee65c, 32'hbbe689e0} /* (7, 28, 15) {real, imag} */,
  {32'hbe8b6e3d, 32'h3e54d238} /* (7, 28, 14) {real, imag} */,
  {32'hbd864640, 32'hbed8e026} /* (7, 28, 13) {real, imag} */,
  {32'hbe1e878a, 32'hbf2416ee} /* (7, 28, 12) {real, imag} */,
  {32'h3dabc3fe, 32'h3f260e9b} /* (7, 28, 11) {real, imag} */,
  {32'h3edb850a, 32'h3e007bca} /* (7, 28, 10) {real, imag} */,
  {32'hbea0e940, 32'h3ea4124b} /* (7, 28, 9) {real, imag} */,
  {32'hbd6feb08, 32'h3f1b9cba} /* (7, 28, 8) {real, imag} */,
  {32'h3e268ac1, 32'hbdc40a28} /* (7, 28, 7) {real, imag} */,
  {32'hbec9cb68, 32'h3dcfe96c} /* (7, 28, 6) {real, imag} */,
  {32'hbe6b7eb1, 32'h3ddc04f6} /* (7, 28, 5) {real, imag} */,
  {32'h3f93734a, 32'hbe6b6c8a} /* (7, 28, 4) {real, imag} */,
  {32'h3e957314, 32'h3f06ddf6} /* (7, 28, 3) {real, imag} */,
  {32'hc0285c1c, 32'h4006f907} /* (7, 28, 2) {real, imag} */,
  {32'h3e975e9a, 32'hc02cb87c} /* (7, 28, 1) {real, imag} */,
  {32'h3fecdcee, 32'hbde8c630} /* (7, 28, 0) {real, imag} */,
  {32'hbfa45525, 32'h3f46695a} /* (7, 27, 31) {real, imag} */,
  {32'h3fabcdc6, 32'hbf95d816} /* (7, 27, 30) {real, imag} */,
  {32'hbdaea4b0, 32'hbbd7ca00} /* (7, 27, 29) {real, imag} */,
  {32'h3cb8c840, 32'hbdbd9c08} /* (7, 27, 28) {real, imag} */,
  {32'h3f34209c, 32'hbea71331} /* (7, 27, 27) {real, imag} */,
  {32'h3f207657, 32'hbf02c462} /* (7, 27, 26) {real, imag} */,
  {32'hbea6cc80, 32'hbe2de43c} /* (7, 27, 25) {real, imag} */,
  {32'h3e135f5c, 32'h3eab7649} /* (7, 27, 24) {real, imag} */,
  {32'h3e51ea63, 32'hbc9bcab8} /* (7, 27, 23) {real, imag} */,
  {32'h3e3d048e, 32'h3ee79b66} /* (7, 27, 22) {real, imag} */,
  {32'hbf0e6e03, 32'h3e6dddd6} /* (7, 27, 21) {real, imag} */,
  {32'h3d9296a0, 32'h3eb17fe6} /* (7, 27, 20) {real, imag} */,
  {32'hbd3eb399, 32'h3e9f3793} /* (7, 27, 19) {real, imag} */,
  {32'hbf145932, 32'hbe0eedc1} /* (7, 27, 18) {real, imag} */,
  {32'hbe6a741d, 32'h3df18934} /* (7, 27, 17) {real, imag} */,
  {32'h3e132f00, 32'h3ea58512} /* (7, 27, 16) {real, imag} */,
  {32'h3df10008, 32'h3b236d90} /* (7, 27, 15) {real, imag} */,
  {32'hbe63b8c2, 32'h3ee4fb40} /* (7, 27, 14) {real, imag} */,
  {32'h3e8f3b08, 32'h3d4e455a} /* (7, 27, 13) {real, imag} */,
  {32'hbde91f84, 32'h3e0f2456} /* (7, 27, 12) {real, imag} */,
  {32'h3e9e0cba, 32'hbe61ff8f} /* (7, 27, 11) {real, imag} */,
  {32'h3e53d02f, 32'hbdb71ad8} /* (7, 27, 10) {real, imag} */,
  {32'hbe53c55e, 32'h3e8d5f4a} /* (7, 27, 9) {real, imag} */,
  {32'h3b616da0, 32'h3ec34b04} /* (7, 27, 8) {real, imag} */,
  {32'hbeea7a8e, 32'hbe430939} /* (7, 27, 7) {real, imag} */,
  {32'hbe8ab28a, 32'hbe0fe854} /* (7, 27, 6) {real, imag} */,
  {32'h3eb6d98f, 32'h3ea258a2} /* (7, 27, 5) {real, imag} */,
  {32'hbec22102, 32'hbdfd4d28} /* (7, 27, 4) {real, imag} */,
  {32'hbdfba380, 32'h3e30f9c2} /* (7, 27, 3) {real, imag} */,
  {32'h3fceb1ae, 32'h3f8b7256} /* (7, 27, 2) {real, imag} */,
  {32'hc02473b8, 32'hbde037e4} /* (7, 27, 1) {real, imag} */,
  {32'hc011524c, 32'h3f514b9c} /* (7, 27, 0) {real, imag} */,
  {32'hbf13b9d5, 32'hbe69946b} /* (7, 26, 31) {real, imag} */,
  {32'hbf5113e2, 32'h3e6c2cf0} /* (7, 26, 30) {real, imag} */,
  {32'hbeaf9bba, 32'hbf5075a5} /* (7, 26, 29) {real, imag} */,
  {32'h3d99aa8d, 32'hbd3934b0} /* (7, 26, 28) {real, imag} */,
  {32'hbdaecab3, 32'hbdb08da5} /* (7, 26, 27) {real, imag} */,
  {32'hbe3ccbb8, 32'h3d894240} /* (7, 26, 26) {real, imag} */,
  {32'h3f693bd0, 32'hbee61d14} /* (7, 26, 25) {real, imag} */,
  {32'h3ede53c4, 32'h3e109405} /* (7, 26, 24) {real, imag} */,
  {32'hbed4eb66, 32'h3e1182ce} /* (7, 26, 23) {real, imag} */,
  {32'h3da55ca0, 32'h3ea80a7c} /* (7, 26, 22) {real, imag} */,
  {32'h3ea3c58f, 32'h3e9b1729} /* (7, 26, 21) {real, imag} */,
  {32'hbe7fb441, 32'hbeeb2218} /* (7, 26, 20) {real, imag} */,
  {32'h3e23694b, 32'h3e55c90a} /* (7, 26, 19) {real, imag} */,
  {32'hbe835005, 32'hbea0de34} /* (7, 26, 18) {real, imag} */,
  {32'hbe27d23e, 32'h3c1f0050} /* (7, 26, 17) {real, imag} */,
  {32'hbebcde08, 32'h3e4460b1} /* (7, 26, 16) {real, imag} */,
  {32'hbda3ccdf, 32'hbe1dfd7f} /* (7, 26, 15) {real, imag} */,
  {32'hbe38ec60, 32'hbdc02754} /* (7, 26, 14) {real, imag} */,
  {32'hbe306ddb, 32'hbe99f858} /* (7, 26, 13) {real, imag} */,
  {32'h3d20ae34, 32'h3e422b18} /* (7, 26, 12) {real, imag} */,
  {32'hbe52eb6b, 32'h3e16b662} /* (7, 26, 11) {real, imag} */,
  {32'hbe120264, 32'hbde8ad34} /* (7, 26, 10) {real, imag} */,
  {32'h3f1449ef, 32'h3e464a8b} /* (7, 26, 9) {real, imag} */,
  {32'h3d6e5368, 32'h3e9bad3f} /* (7, 26, 8) {real, imag} */,
  {32'h3ef6317a, 32'hbc982130} /* (7, 26, 7) {real, imag} */,
  {32'hbdd01ac8, 32'h3b8b0f80} /* (7, 26, 6) {real, imag} */,
  {32'h3f15b2eb, 32'hbf0ca3a8} /* (7, 26, 5) {real, imag} */,
  {32'hbe7ac502, 32'hbedcfbeb} /* (7, 26, 4) {real, imag} */,
  {32'hbe1780cf, 32'h3ee6be86} /* (7, 26, 3) {real, imag} */,
  {32'hbdd8836c, 32'h3ecc5e3d} /* (7, 26, 2) {real, imag} */,
  {32'h3e533625, 32'hbf0933b2} /* (7, 26, 1) {real, imag} */,
  {32'hbd75e64c, 32'h3ebb646a} /* (7, 26, 0) {real, imag} */,
  {32'hbe5d6c84, 32'hbf1536a7} /* (7, 25, 31) {real, imag} */,
  {32'hbe17c106, 32'h3f917784} /* (7, 25, 30) {real, imag} */,
  {32'hbed8e1a7, 32'hbf4ae47e} /* (7, 25, 29) {real, imag} */,
  {32'h3e2eee4c, 32'hbf42c4ed} /* (7, 25, 28) {real, imag} */,
  {32'h3f96df1b, 32'h3e8c6c8e} /* (7, 25, 27) {real, imag} */,
  {32'h3f276907, 32'hbdfb301c} /* (7, 25, 26) {real, imag} */,
  {32'hbe83307d, 32'h3f2f7cd4} /* (7, 25, 25) {real, imag} */,
  {32'hbf07e855, 32'h3ea1c52c} /* (7, 25, 24) {real, imag} */,
  {32'h3edbee02, 32'hbf48148e} /* (7, 25, 23) {real, imag} */,
  {32'h3f3be576, 32'hbed6a8b7} /* (7, 25, 22) {real, imag} */,
  {32'hbed81164, 32'hbca11a40} /* (7, 25, 21) {real, imag} */,
  {32'hbe666e14, 32'h3f0a44c0} /* (7, 25, 20) {real, imag} */,
  {32'h3e12eede, 32'hbed51574} /* (7, 25, 19) {real, imag} */,
  {32'h3dded06a, 32'h3e77b616} /* (7, 25, 18) {real, imag} */,
  {32'hbc0aacd8, 32'h3e2205ee} /* (7, 25, 17) {real, imag} */,
  {32'hbe34ef65, 32'h3e037ec5} /* (7, 25, 16) {real, imag} */,
  {32'hbe7390a4, 32'hbd9b40ee} /* (7, 25, 15) {real, imag} */,
  {32'h3deeb45a, 32'h3d9364be} /* (7, 25, 14) {real, imag} */,
  {32'hbd2bb8d8, 32'hbe67849d} /* (7, 25, 13) {real, imag} */,
  {32'hbd2041be, 32'hbe017d28} /* (7, 25, 12) {real, imag} */,
  {32'h3df0ce72, 32'h3eb7e75b} /* (7, 25, 11) {real, imag} */,
  {32'hbe501160, 32'hbdafb3ab} /* (7, 25, 10) {real, imag} */,
  {32'hbe8e9fde, 32'h3e3e0516} /* (7, 25, 9) {real, imag} */,
  {32'h3e994be8, 32'h3e894afa} /* (7, 25, 8) {real, imag} */,
  {32'hbe987117, 32'hbf47916c} /* (7, 25, 7) {real, imag} */,
  {32'hbd6c870c, 32'hbef1a2a0} /* (7, 25, 6) {real, imag} */,
  {32'h3e8b9255, 32'h3e289574} /* (7, 25, 5) {real, imag} */,
  {32'hbd977096, 32'hbe2f4bf6} /* (7, 25, 4) {real, imag} */,
  {32'hbf41cbe2, 32'hbe02e6f2} /* (7, 25, 3) {real, imag} */,
  {32'h3e8b396a, 32'h3e0d12c4} /* (7, 25, 2) {real, imag} */,
  {32'hbe0097ac, 32'h3e83c292} /* (7, 25, 1) {real, imag} */,
  {32'h3edc6cf6, 32'hbe880cec} /* (7, 25, 0) {real, imag} */,
  {32'hbf05bea2, 32'h3f88ba72} /* (7, 24, 31) {real, imag} */,
  {32'h3f2bc60a, 32'hbe1a63d8} /* (7, 24, 30) {real, imag} */,
  {32'h3e271798, 32'hbe79c8ad} /* (7, 24, 29) {real, imag} */,
  {32'hbef51275, 32'h3f0353c9} /* (7, 24, 28) {real, imag} */,
  {32'hbf0a9c0a, 32'hbdc1f356} /* (7, 24, 27) {real, imag} */,
  {32'hbf039bc4, 32'hbd2ab288} /* (7, 24, 26) {real, imag} */,
  {32'hbed62194, 32'hbe42a799} /* (7, 24, 25) {real, imag} */,
  {32'hbe02bea0, 32'hbf6d49e8} /* (7, 24, 24) {real, imag} */,
  {32'hbefc6ebc, 32'h3eb580c1} /* (7, 24, 23) {real, imag} */,
  {32'h3e7224d9, 32'h3e327aeb} /* (7, 24, 22) {real, imag} */,
  {32'h3dec51f4, 32'hbf1448a2} /* (7, 24, 21) {real, imag} */,
  {32'hbd93d438, 32'h3e00b5a3} /* (7, 24, 20) {real, imag} */,
  {32'hbf2678ba, 32'hbe2b537b} /* (7, 24, 19) {real, imag} */,
  {32'h3f2bd7d9, 32'h3e9d457a} /* (7, 24, 18) {real, imag} */,
  {32'h3e0c8756, 32'h3eafee88} /* (7, 24, 17) {real, imag} */,
  {32'hbe8cce62, 32'hbe0cbf28} /* (7, 24, 16) {real, imag} */,
  {32'hbf05b17a, 32'hbe91e174} /* (7, 24, 15) {real, imag} */,
  {32'h3eae1656, 32'hbe91e712} /* (7, 24, 14) {real, imag} */,
  {32'hbe01fc1c, 32'hbd1fc260} /* (7, 24, 13) {real, imag} */,
  {32'hbe50db5c, 32'hbf0be5fb} /* (7, 24, 12) {real, imag} */,
  {32'hbe33c6bd, 32'hbed468ce} /* (7, 24, 11) {real, imag} */,
  {32'h3d17da88, 32'hbcd96878} /* (7, 24, 10) {real, imag} */,
  {32'h3e800960, 32'h3ef33d78} /* (7, 24, 9) {real, imag} */,
  {32'h3eda3f11, 32'h3f340aad} /* (7, 24, 8) {real, imag} */,
  {32'hbe8ed724, 32'h3edbc6aa} /* (7, 24, 7) {real, imag} */,
  {32'h3ea100f8, 32'h3ec3c935} /* (7, 24, 6) {real, imag} */,
  {32'h3f7b1944, 32'h3ed9517a} /* (7, 24, 5) {real, imag} */,
  {32'h3ed69b50, 32'hbdf7efea} /* (7, 24, 4) {real, imag} */,
  {32'h3e82b91c, 32'h3e8acfe4} /* (7, 24, 3) {real, imag} */,
  {32'h3f67772d, 32'hbf0daf33} /* (7, 24, 2) {real, imag} */,
  {32'hbfc45dc3, 32'h3f30f6f4} /* (7, 24, 1) {real, imag} */,
  {32'hbf559ae1, 32'h3f1d5430} /* (7, 24, 0) {real, imag} */,
  {32'hbf23e8b2, 32'hbd353f94} /* (7, 23, 31) {real, imag} */,
  {32'hbefc6eb4, 32'h3e10460c} /* (7, 23, 30) {real, imag} */,
  {32'hbd90ddc5, 32'hbeaa54ab} /* (7, 23, 29) {real, imag} */,
  {32'h3e83b555, 32'hbe7d0e40} /* (7, 23, 28) {real, imag} */,
  {32'hbe1c122e, 32'hbeb099cb} /* (7, 23, 27) {real, imag} */,
  {32'hbee34717, 32'h3e738c0e} /* (7, 23, 26) {real, imag} */,
  {32'h3d01b375, 32'hbf009196} /* (7, 23, 25) {real, imag} */,
  {32'hbdf344c6, 32'h3db57eaa} /* (7, 23, 24) {real, imag} */,
  {32'hbea5075c, 32'hbf2dd430} /* (7, 23, 23) {real, imag} */,
  {32'h3e71f827, 32'h3e50a882} /* (7, 23, 22) {real, imag} */,
  {32'h3e8f7d66, 32'hbd048a34} /* (7, 23, 21) {real, imag} */,
  {32'h3db8f8d8, 32'hbe262cc7} /* (7, 23, 20) {real, imag} */,
  {32'hbd83aa64, 32'h3ed94fea} /* (7, 23, 19) {real, imag} */,
  {32'h3e81c450, 32'hbd9c057d} /* (7, 23, 18) {real, imag} */,
  {32'h3e040bd2, 32'h3ea91a2e} /* (7, 23, 17) {real, imag} */,
  {32'h3dd9950a, 32'hbe8b14f2} /* (7, 23, 16) {real, imag} */,
  {32'h3dfef25a, 32'hbe72c3b0} /* (7, 23, 15) {real, imag} */,
  {32'hbef6a155, 32'h3e2e0d62} /* (7, 23, 14) {real, imag} */,
  {32'h3eed8db2, 32'hbeb7a2ad} /* (7, 23, 13) {real, imag} */,
  {32'h3d918b70, 32'h3dd6a280} /* (7, 23, 12) {real, imag} */,
  {32'hbcc3aa10, 32'h3e95329b} /* (7, 23, 11) {real, imag} */,
  {32'h3f293f92, 32'h3e2e5ddf} /* (7, 23, 10) {real, imag} */,
  {32'hbf0d934e, 32'h3f08890a} /* (7, 23, 9) {real, imag} */,
  {32'h3e3a57d0, 32'h3ed76f5c} /* (7, 23, 8) {real, imag} */,
  {32'hbf0c599b, 32'h3e2cb604} /* (7, 23, 7) {real, imag} */,
  {32'h3d678818, 32'h3e3594ca} /* (7, 23, 6) {real, imag} */,
  {32'hbee8ea77, 32'hbe70daf6} /* (7, 23, 5) {real, imag} */,
  {32'hbd018f2a, 32'hbc3bfb90} /* (7, 23, 4) {real, imag} */,
  {32'hbcb4d3a8, 32'h3c870108} /* (7, 23, 3) {real, imag} */,
  {32'h3edf4c0a, 32'h3f33a7da} /* (7, 23, 2) {real, imag} */,
  {32'hbec7f4f4, 32'hbf48ff99} /* (7, 23, 1) {real, imag} */,
  {32'hbe8cab70, 32'h3e2a75bb} /* (7, 23, 0) {real, imag} */,
  {32'h3f0882a9, 32'h3e15d1f6} /* (7, 22, 31) {real, imag} */,
  {32'h3d02fdbc, 32'h3ebcd440} /* (7, 22, 30) {real, imag} */,
  {32'hbe3bae5b, 32'hbf25982e} /* (7, 22, 29) {real, imag} */,
  {32'hbd687f66, 32'h3d4cdc9c} /* (7, 22, 28) {real, imag} */,
  {32'h3f23294a, 32'h3e2dd336} /* (7, 22, 27) {real, imag} */,
  {32'hbea51743, 32'hbec68402} /* (7, 22, 26) {real, imag} */,
  {32'hbe44900e, 32'h3ed2e7ee} /* (7, 22, 25) {real, imag} */,
  {32'hbe00ef45, 32'h3ddd1a5a} /* (7, 22, 24) {real, imag} */,
  {32'h3e59d1c7, 32'hbe3e809b} /* (7, 22, 23) {real, imag} */,
  {32'hbecb8a6c, 32'hbdea8332} /* (7, 22, 22) {real, imag} */,
  {32'h3e78ab78, 32'h3f29c9e2} /* (7, 22, 21) {real, imag} */,
  {32'h3e932994, 32'hbf0c2d91} /* (7, 22, 20) {real, imag} */,
  {32'h3ef1a90e, 32'h3e7572c3} /* (7, 22, 19) {real, imag} */,
  {32'hbecd89c3, 32'h3ec21b37} /* (7, 22, 18) {real, imag} */,
  {32'hbd443ac6, 32'h3e25e844} /* (7, 22, 17) {real, imag} */,
  {32'hbbfc1ca0, 32'h3e58a611} /* (7, 22, 16) {real, imag} */,
  {32'hbe894e9a, 32'h3e507b9e} /* (7, 22, 15) {real, imag} */,
  {32'hbde5f34c, 32'hbc6bb9f0} /* (7, 22, 14) {real, imag} */,
  {32'h3e7647c9, 32'hbf0f47b8} /* (7, 22, 13) {real, imag} */,
  {32'h3f48129a, 32'hbced4e20} /* (7, 22, 12) {real, imag} */,
  {32'h3f56fd4b, 32'h3c9a2da0} /* (7, 22, 11) {real, imag} */,
  {32'hbf156590, 32'h3e84fa9e} /* (7, 22, 10) {real, imag} */,
  {32'h3e51ca1c, 32'h3e6a8bae} /* (7, 22, 9) {real, imag} */,
  {32'hbed9c1e3, 32'hbe01fc71} /* (7, 22, 8) {real, imag} */,
  {32'h3dea54c2, 32'h3effd1dc} /* (7, 22, 7) {real, imag} */,
  {32'h3e968c53, 32'h3e1623a9} /* (7, 22, 6) {real, imag} */,
  {32'h3e8a3e92, 32'h3eda078d} /* (7, 22, 5) {real, imag} */,
  {32'h3cb10efc, 32'hbf05fc28} /* (7, 22, 4) {real, imag} */,
  {32'hbeb719f2, 32'h3ec0d69b} /* (7, 22, 3) {real, imag} */,
  {32'hbec630ac, 32'hbe3d22a0} /* (7, 22, 2) {real, imag} */,
  {32'hbc32af60, 32'hbe542cf5} /* (7, 22, 1) {real, imag} */,
  {32'hbdeb884c, 32'hbf52b5c6} /* (7, 22, 0) {real, imag} */,
  {32'h3d4db350, 32'h3f517db1} /* (7, 21, 31) {real, imag} */,
  {32'hbe169c6f, 32'hbf032e61} /* (7, 21, 30) {real, imag} */,
  {32'h3ee543e2, 32'h3f377cc1} /* (7, 21, 29) {real, imag} */,
  {32'h3e4c5f40, 32'h3f32c1ce} /* (7, 21, 28) {real, imag} */,
  {32'hbdbf3f74, 32'hbe89e67c} /* (7, 21, 27) {real, imag} */,
  {32'h3e9bc99a, 32'hbf2789de} /* (7, 21, 26) {real, imag} */,
  {32'h3e9dbd94, 32'hbe1d6376} /* (7, 21, 25) {real, imag} */,
  {32'hbd98252c, 32'hbe102c8e} /* (7, 21, 24) {real, imag} */,
  {32'h3ec918f2, 32'h3f1376bf} /* (7, 21, 23) {real, imag} */,
  {32'hbf0973e0, 32'hbf1d56b6} /* (7, 21, 22) {real, imag} */,
  {32'hbdf5e3b8, 32'hbeba6fa0} /* (7, 21, 21) {real, imag} */,
  {32'h3cef6e68, 32'h3ec9e075} /* (7, 21, 20) {real, imag} */,
  {32'hbd8808e4, 32'h3cabaec8} /* (7, 21, 19) {real, imag} */,
  {32'hbec4b906, 32'h3ed244d0} /* (7, 21, 18) {real, imag} */,
  {32'h3ea1e5d8, 32'hbe4cee7b} /* (7, 21, 17) {real, imag} */,
  {32'h3e9d38f0, 32'hbe0d4c9e} /* (7, 21, 16) {real, imag} */,
  {32'hbe7a9f6b, 32'h3e053ebd} /* (7, 21, 15) {real, imag} */,
  {32'h3eab4a7f, 32'hbe3352f6} /* (7, 21, 14) {real, imag} */,
  {32'h3e47a9da, 32'h3c9864c8} /* (7, 21, 13) {real, imag} */,
  {32'h3f462406, 32'hbcd89b24} /* (7, 21, 12) {real, imag} */,
  {32'h3f0962ff, 32'h3e9918f2} /* (7, 21, 11) {real, imag} */,
  {32'hbe15bd6e, 32'h3e85abdd} /* (7, 21, 10) {real, imag} */,
  {32'hbf539410, 32'hbeec07e5} /* (7, 21, 9) {real, imag} */,
  {32'hbe6b2e5a, 32'hbee1b4fe} /* (7, 21, 8) {real, imag} */,
  {32'hbf35b176, 32'h3de7affe} /* (7, 21, 7) {real, imag} */,
  {32'h3e8b401b, 32'hbe50c105} /* (7, 21, 6) {real, imag} */,
  {32'h3d661b48, 32'hbe85c4f9} /* (7, 21, 5) {real, imag} */,
  {32'hbeb28038, 32'h3e98b778} /* (7, 21, 4) {real, imag} */,
  {32'h3e9bab4c, 32'hbeb335a0} /* (7, 21, 3) {real, imag} */,
  {32'h3f32056c, 32'hbba6c680} /* (7, 21, 2) {real, imag} */,
  {32'h3c8e2b00, 32'h3e677718} /* (7, 21, 1) {real, imag} */,
  {32'hbea2e90c, 32'h3ea458d1} /* (7, 21, 0) {real, imag} */,
  {32'h3efbb391, 32'h3cf186dc} /* (7, 20, 31) {real, imag} */,
  {32'h3d02cfe8, 32'h3de9a7a4} /* (7, 20, 30) {real, imag} */,
  {32'hbf1545bc, 32'h3e5505fb} /* (7, 20, 29) {real, imag} */,
  {32'h3f10a7b4, 32'h3ec0f98f} /* (7, 20, 28) {real, imag} */,
  {32'hbf087442, 32'h3d8faf84} /* (7, 20, 27) {real, imag} */,
  {32'hbdb9d5a5, 32'hbee2a084} /* (7, 20, 26) {real, imag} */,
  {32'h3ee141d8, 32'h3e63025e} /* (7, 20, 25) {real, imag} */,
  {32'h3b3fd940, 32'hbe5a5c30} /* (7, 20, 24) {real, imag} */,
  {32'hbee444bc, 32'h3d9f49a0} /* (7, 20, 23) {real, imag} */,
  {32'h3ecb822c, 32'hbf2ebbb2} /* (7, 20, 22) {real, imag} */,
  {32'hbdc75460, 32'h3e0fcab2} /* (7, 20, 21) {real, imag} */,
  {32'h3ed99a99, 32'h3ca7eb98} /* (7, 20, 20) {real, imag} */,
  {32'hbec6d037, 32'hbeaf92d9} /* (7, 20, 19) {real, imag} */,
  {32'h3e29b576, 32'hbedad8ec} /* (7, 20, 18) {real, imag} */,
  {32'hbdde01bc, 32'hbe253c40} /* (7, 20, 17) {real, imag} */,
  {32'h3c7bdf68, 32'h3ecb2b0a} /* (7, 20, 16) {real, imag} */,
  {32'h3ec4dfd9, 32'hbcf52dd8} /* (7, 20, 15) {real, imag} */,
  {32'hbdb18f0a, 32'hbcd24c74} /* (7, 20, 14) {real, imag} */,
  {32'hbe982b34, 32'h3e9fc0a0} /* (7, 20, 13) {real, imag} */,
  {32'h3e50f5a6, 32'hbe7179f9} /* (7, 20, 12) {real, imag} */,
  {32'hbd749c70, 32'h3f0925ac} /* (7, 20, 11) {real, imag} */,
  {32'hbef37009, 32'h3d52ad0a} /* (7, 20, 10) {real, imag} */,
  {32'h3dca60c8, 32'hbee0a0d4} /* (7, 20, 9) {real, imag} */,
  {32'hbe652549, 32'hbc4e9b38} /* (7, 20, 8) {real, imag} */,
  {32'h3df383e4, 32'hbc25c390} /* (7, 20, 7) {real, imag} */,
  {32'h3e54237e, 32'hbeeb17d3} /* (7, 20, 6) {real, imag} */,
  {32'hbdb2bab4, 32'h3dace1da} /* (7, 20, 5) {real, imag} */,
  {32'hbec80d48, 32'hbee1a35a} /* (7, 20, 4) {real, imag} */,
  {32'h3d05e688, 32'hbe75f75c} /* (7, 20, 3) {real, imag} */,
  {32'hbdcd4a68, 32'h3bf120a0} /* (7, 20, 2) {real, imag} */,
  {32'h3e3bbf3f, 32'h3db8c002} /* (7, 20, 1) {real, imag} */,
  {32'h3d075290, 32'h3d4e2638} /* (7, 20, 0) {real, imag} */,
  {32'h3dbd99d8, 32'h3d8d5caf} /* (7, 19, 31) {real, imag} */,
  {32'hbde4611e, 32'h3f052dee} /* (7, 19, 30) {real, imag} */,
  {32'hbca401dc, 32'hbf053e70} /* (7, 19, 29) {real, imag} */,
  {32'hbd443800, 32'hbe3e6f38} /* (7, 19, 28) {real, imag} */,
  {32'h3e0277e3, 32'hbc49f240} /* (7, 19, 27) {real, imag} */,
  {32'hbcf6df52, 32'hbd8752b4} /* (7, 19, 26) {real, imag} */,
  {32'h3e438365, 32'hbe218244} /* (7, 19, 25) {real, imag} */,
  {32'h3ca94f20, 32'h3ea50654} /* (7, 19, 24) {real, imag} */,
  {32'hbe28f11e, 32'hbea8b7c8} /* (7, 19, 23) {real, imag} */,
  {32'hbf079be7, 32'hbdf2b803} /* (7, 19, 22) {real, imag} */,
  {32'h3e074c6a, 32'hbefd1442} /* (7, 19, 21) {real, imag} */,
  {32'h3e84509c, 32'hbf16d098} /* (7, 19, 20) {real, imag} */,
  {32'h3ec6b91e, 32'h3dcec295} /* (7, 19, 19) {real, imag} */,
  {32'hbefb6811, 32'hbdf04fe4} /* (7, 19, 18) {real, imag} */,
  {32'h3e89f7f2, 32'hbe38d96e} /* (7, 19, 17) {real, imag} */,
  {32'h3e1a3d28, 32'h3eae913f} /* (7, 19, 16) {real, imag} */,
  {32'h3d47e5c8, 32'h3e3cbe55} /* (7, 19, 15) {real, imag} */,
  {32'hbf21e2a2, 32'h3e7aaa42} /* (7, 19, 14) {real, imag} */,
  {32'h3f1c4835, 32'hbec21c1e} /* (7, 19, 13) {real, imag} */,
  {32'hbedd9231, 32'h3ea34ee2} /* (7, 19, 12) {real, imag} */,
  {32'hbeff6fb7, 32'h3d572648} /* (7, 19, 11) {real, imag} */,
  {32'hbdb81c86, 32'h3da0c01a} /* (7, 19, 10) {real, imag} */,
  {32'hbe8b3242, 32'h3c256240} /* (7, 19, 9) {real, imag} */,
  {32'hbe87782a, 32'h3ea38236} /* (7, 19, 8) {real, imag} */,
  {32'h3ed8c5ef, 32'hbd0015f7} /* (7, 19, 7) {real, imag} */,
  {32'h3ebc0425, 32'h3e5bd481} /* (7, 19, 6) {real, imag} */,
  {32'hbd56da74, 32'h3e63a6a2} /* (7, 19, 5) {real, imag} */,
  {32'h3d57359c, 32'hbd3b7c36} /* (7, 19, 4) {real, imag} */,
  {32'h3e1206f4, 32'hbedb394b} /* (7, 19, 3) {real, imag} */,
  {32'hbeb97424, 32'hbe37d039} /* (7, 19, 2) {real, imag} */,
  {32'h3dfbd264, 32'hbf05c4a3} /* (7, 19, 1) {real, imag} */,
  {32'hbf7b397e, 32'hbe91f938} /* (7, 19, 0) {real, imag} */,
  {32'h3df510c3, 32'h3e8e3876} /* (7, 18, 31) {real, imag} */,
  {32'h3d950098, 32'h3d07f502} /* (7, 18, 30) {real, imag} */,
  {32'h3cd042fc, 32'h3d31ef7a} /* (7, 18, 29) {real, imag} */,
  {32'hbd9eeefe, 32'hbe726661} /* (7, 18, 28) {real, imag} */,
  {32'hbdfbcb5c, 32'hbebd04bc} /* (7, 18, 27) {real, imag} */,
  {32'h3e0f65eb, 32'hbe737ed1} /* (7, 18, 26) {real, imag} */,
  {32'hbe8851d1, 32'hbd861c64} /* (7, 18, 25) {real, imag} */,
  {32'h3ddf5f28, 32'hbe4946fb} /* (7, 18, 24) {real, imag} */,
  {32'hbec112f2, 32'hbed49f0a} /* (7, 18, 23) {real, imag} */,
  {32'h3e37e22e, 32'h3f13b553} /* (7, 18, 22) {real, imag} */,
  {32'hbda172fc, 32'h3e203442} /* (7, 18, 21) {real, imag} */,
  {32'h3c169d7c, 32'hbe5a4ded} /* (7, 18, 20) {real, imag} */,
  {32'hbe54050a, 32'h3e86250e} /* (7, 18, 19) {real, imag} */,
  {32'hbeb6d7f9, 32'hbeb84937} /* (7, 18, 18) {real, imag} */,
  {32'hbe7baca8, 32'h3cf648d2} /* (7, 18, 17) {real, imag} */,
  {32'h3c231ee0, 32'hbe9d823d} /* (7, 18, 16) {real, imag} */,
  {32'h3e17e3bf, 32'h3da3a8a4} /* (7, 18, 15) {real, imag} */,
  {32'hbf5e5060, 32'h3eac2a5a} /* (7, 18, 14) {real, imag} */,
  {32'hbe588c8a, 32'hbd875a36} /* (7, 18, 13) {real, imag} */,
  {32'h3e8de5f9, 32'h3d8b8bb8} /* (7, 18, 12) {real, imag} */,
  {32'h3d486b98, 32'h3ef5521a} /* (7, 18, 11) {real, imag} */,
  {32'hbd6fa308, 32'hbdf20082} /* (7, 18, 10) {real, imag} */,
  {32'hbe293415, 32'hbe75f9e8} /* (7, 18, 9) {real, imag} */,
  {32'h3da27ffb, 32'h3e66fb3c} /* (7, 18, 8) {real, imag} */,
  {32'hbd382fa0, 32'h3ea9d277} /* (7, 18, 7) {real, imag} */,
  {32'h3ea49dcf, 32'h3e41649d} /* (7, 18, 6) {real, imag} */,
  {32'hbe2bad20, 32'hbe575517} /* (7, 18, 5) {real, imag} */,
  {32'hbd02c188, 32'hbe225260} /* (7, 18, 4) {real, imag} */,
  {32'h3e6ceec2, 32'h3ea331b3} /* (7, 18, 3) {real, imag} */,
  {32'h3d21eb46, 32'hbd942837} /* (7, 18, 2) {real, imag} */,
  {32'hbdd579ac, 32'h3ef52167} /* (7, 18, 1) {real, imag} */,
  {32'h3ce44210, 32'h3d436878} /* (7, 18, 0) {real, imag} */,
  {32'hbd1a5630, 32'hbeb1a1ae} /* (7, 17, 31) {real, imag} */,
  {32'hbe2b5312, 32'hbe1e506d} /* (7, 17, 30) {real, imag} */,
  {32'h3df6ce39, 32'hbe146c30} /* (7, 17, 29) {real, imag} */,
  {32'hbe4f6fb6, 32'hbef99252} /* (7, 17, 28) {real, imag} */,
  {32'h3efac091, 32'hbdad2930} /* (7, 17, 27) {real, imag} */,
  {32'hbb526ea0, 32'h3d49347b} /* (7, 17, 26) {real, imag} */,
  {32'hbf130ff1, 32'hbad46600} /* (7, 17, 25) {real, imag} */,
  {32'h3e8c8707, 32'h3d81977c} /* (7, 17, 24) {real, imag} */,
  {32'h3e8c45e0, 32'h3f34d70e} /* (7, 17, 23) {real, imag} */,
  {32'h3eb53b57, 32'hbeda02d3} /* (7, 17, 22) {real, imag} */,
  {32'h3e9ff032, 32'hbc1f1310} /* (7, 17, 21) {real, imag} */,
  {32'hbf0c5bda, 32'h3e0f4022} /* (7, 17, 20) {real, imag} */,
  {32'h3e35191c, 32'hbde18967} /* (7, 17, 19) {real, imag} */,
  {32'h3e41c9ac, 32'hbd01b52c} /* (7, 17, 18) {real, imag} */,
  {32'h3e204870, 32'hbe73cfaa} /* (7, 17, 17) {real, imag} */,
  {32'h3d28c5e8, 32'h3da6eae5} /* (7, 17, 16) {real, imag} */,
  {32'h3cfcc4a8, 32'h3d8f5cdf} /* (7, 17, 15) {real, imag} */,
  {32'hbd25383c, 32'h3d217690} /* (7, 17, 14) {real, imag} */,
  {32'hbe9ae312, 32'hbdea00f9} /* (7, 17, 13) {real, imag} */,
  {32'h3e6e959c, 32'hbea59852} /* (7, 17, 12) {real, imag} */,
  {32'hbe944dde, 32'hbe4ab9a1} /* (7, 17, 11) {real, imag} */,
  {32'hbce0b400, 32'hbe87b6c0} /* (7, 17, 10) {real, imag} */,
  {32'hbe4cc6c1, 32'h3e0b6d76} /* (7, 17, 9) {real, imag} */,
  {32'hbc89c1c4, 32'h3f24c34b} /* (7, 17, 8) {real, imag} */,
  {32'hbd78e47e, 32'hbed907a0} /* (7, 17, 7) {real, imag} */,
  {32'hbd5125e9, 32'hbebd0f10} /* (7, 17, 6) {real, imag} */,
  {32'h3d360db2, 32'hbda1e23e} /* (7, 17, 5) {real, imag} */,
  {32'h3e1abc20, 32'h3de98cd2} /* (7, 17, 4) {real, imag} */,
  {32'h3b89d3b0, 32'h3ede79de} /* (7, 17, 3) {real, imag} */,
  {32'h3ddf0dba, 32'hbdf7bbee} /* (7, 17, 2) {real, imag} */,
  {32'hbee603b6, 32'hbdffe5f6} /* (7, 17, 1) {real, imag} */,
  {32'h3e1455e5, 32'hbe0b0b16} /* (7, 17, 0) {real, imag} */,
  {32'h3df4e3b7, 32'hbd5f50e8} /* (7, 16, 31) {real, imag} */,
  {32'hbd0cdcd6, 32'h3d9c9011} /* (7, 16, 30) {real, imag} */,
  {32'h3e8040b6, 32'hbe0d0173} /* (7, 16, 29) {real, imag} */,
  {32'hbdbf8820, 32'h3e293748} /* (7, 16, 28) {real, imag} */,
  {32'hbce2850a, 32'h3dff56ba} /* (7, 16, 27) {real, imag} */,
  {32'h3da216bb, 32'h3bf253e0} /* (7, 16, 26) {real, imag} */,
  {32'h3eab43b8, 32'hbe728cc2} /* (7, 16, 25) {real, imag} */,
  {32'hbeb0e6d7, 32'h3e2ef458} /* (7, 16, 24) {real, imag} */,
  {32'h3e1c7e90, 32'h3ece4b64} /* (7, 16, 23) {real, imag} */,
  {32'h3d9ea4d6, 32'hbd301c84} /* (7, 16, 22) {real, imag} */,
  {32'h3c976c64, 32'hbf202613} /* (7, 16, 21) {real, imag} */,
  {32'hbe1eb12b, 32'h3d41250c} /* (7, 16, 20) {real, imag} */,
  {32'h3ec40c76, 32'hbc9261ac} /* (7, 16, 19) {real, imag} */,
  {32'hbd2ceb20, 32'hbb55fec8} /* (7, 16, 18) {real, imag} */,
  {32'h3e0e6c82, 32'h3e2435a2} /* (7, 16, 17) {real, imag} */,
  {32'h3e37514e, 32'h00000000} /* (7, 16, 16) {real, imag} */,
  {32'h3e0e6c82, 32'hbe2435a2} /* (7, 16, 15) {real, imag} */,
  {32'hbd2ceb20, 32'h3b55fec8} /* (7, 16, 14) {real, imag} */,
  {32'h3ec40c76, 32'h3c9261ac} /* (7, 16, 13) {real, imag} */,
  {32'hbe1eb12b, 32'hbd41250c} /* (7, 16, 12) {real, imag} */,
  {32'h3c976c64, 32'h3f202613} /* (7, 16, 11) {real, imag} */,
  {32'h3d9ea4d6, 32'h3d301c84} /* (7, 16, 10) {real, imag} */,
  {32'h3e1c7e90, 32'hbece4b64} /* (7, 16, 9) {real, imag} */,
  {32'hbeb0e6d7, 32'hbe2ef458} /* (7, 16, 8) {real, imag} */,
  {32'h3eab43b8, 32'h3e728cc2} /* (7, 16, 7) {real, imag} */,
  {32'h3da216bb, 32'hbbf253e0} /* (7, 16, 6) {real, imag} */,
  {32'hbce2850a, 32'hbdff56ba} /* (7, 16, 5) {real, imag} */,
  {32'hbdbf8820, 32'hbe293748} /* (7, 16, 4) {real, imag} */,
  {32'h3e8040b6, 32'h3e0d0173} /* (7, 16, 3) {real, imag} */,
  {32'hbd0cdcd6, 32'hbd9c9011} /* (7, 16, 2) {real, imag} */,
  {32'h3df4e3b7, 32'h3d5f50e8} /* (7, 16, 1) {real, imag} */,
  {32'hbe6296d6, 32'h00000000} /* (7, 16, 0) {real, imag} */,
  {32'hbee603b6, 32'h3dffe5f6} /* (7, 15, 31) {real, imag} */,
  {32'h3ddf0dba, 32'h3df7bbee} /* (7, 15, 30) {real, imag} */,
  {32'h3b89d3b0, 32'hbede79de} /* (7, 15, 29) {real, imag} */,
  {32'h3e1abc20, 32'hbde98cd2} /* (7, 15, 28) {real, imag} */,
  {32'h3d360db2, 32'h3da1e23e} /* (7, 15, 27) {real, imag} */,
  {32'hbd5125e9, 32'h3ebd0f10} /* (7, 15, 26) {real, imag} */,
  {32'hbd78e47e, 32'h3ed907a0} /* (7, 15, 25) {real, imag} */,
  {32'hbc89c1c4, 32'hbf24c34b} /* (7, 15, 24) {real, imag} */,
  {32'hbe4cc6c1, 32'hbe0b6d76} /* (7, 15, 23) {real, imag} */,
  {32'hbce0b400, 32'h3e87b6c0} /* (7, 15, 22) {real, imag} */,
  {32'hbe944dde, 32'h3e4ab9a1} /* (7, 15, 21) {real, imag} */,
  {32'h3e6e959c, 32'h3ea59852} /* (7, 15, 20) {real, imag} */,
  {32'hbe9ae312, 32'h3dea00f9} /* (7, 15, 19) {real, imag} */,
  {32'hbd25383c, 32'hbd217690} /* (7, 15, 18) {real, imag} */,
  {32'h3cfcc4a8, 32'hbd8f5cdf} /* (7, 15, 17) {real, imag} */,
  {32'h3d28c5e8, 32'hbda6eae5} /* (7, 15, 16) {real, imag} */,
  {32'h3e204870, 32'h3e73cfaa} /* (7, 15, 15) {real, imag} */,
  {32'h3e41c9ac, 32'h3d01b52c} /* (7, 15, 14) {real, imag} */,
  {32'h3e35191c, 32'h3de18967} /* (7, 15, 13) {real, imag} */,
  {32'hbf0c5bda, 32'hbe0f4022} /* (7, 15, 12) {real, imag} */,
  {32'h3e9ff032, 32'h3c1f1310} /* (7, 15, 11) {real, imag} */,
  {32'h3eb53b57, 32'h3eda02d3} /* (7, 15, 10) {real, imag} */,
  {32'h3e8c45e0, 32'hbf34d70e} /* (7, 15, 9) {real, imag} */,
  {32'h3e8c8707, 32'hbd81977c} /* (7, 15, 8) {real, imag} */,
  {32'hbf130ff1, 32'h3ad46600} /* (7, 15, 7) {real, imag} */,
  {32'hbb526ea0, 32'hbd49347b} /* (7, 15, 6) {real, imag} */,
  {32'h3efac091, 32'h3dad2930} /* (7, 15, 5) {real, imag} */,
  {32'hbe4f6fb6, 32'h3ef99252} /* (7, 15, 4) {real, imag} */,
  {32'h3df6ce39, 32'h3e146c30} /* (7, 15, 3) {real, imag} */,
  {32'hbe2b5312, 32'h3e1e506d} /* (7, 15, 2) {real, imag} */,
  {32'hbd1a5630, 32'h3eb1a1ae} /* (7, 15, 1) {real, imag} */,
  {32'h3e1455e5, 32'h3e0b0b16} /* (7, 15, 0) {real, imag} */,
  {32'hbdd579ac, 32'hbef52167} /* (7, 14, 31) {real, imag} */,
  {32'h3d21eb46, 32'h3d942837} /* (7, 14, 30) {real, imag} */,
  {32'h3e6ceec2, 32'hbea331b3} /* (7, 14, 29) {real, imag} */,
  {32'hbd02c188, 32'h3e225260} /* (7, 14, 28) {real, imag} */,
  {32'hbe2bad20, 32'h3e575517} /* (7, 14, 27) {real, imag} */,
  {32'h3ea49dcf, 32'hbe41649d} /* (7, 14, 26) {real, imag} */,
  {32'hbd382fa0, 32'hbea9d277} /* (7, 14, 25) {real, imag} */,
  {32'h3da27ffb, 32'hbe66fb3c} /* (7, 14, 24) {real, imag} */,
  {32'hbe293415, 32'h3e75f9e8} /* (7, 14, 23) {real, imag} */,
  {32'hbd6fa308, 32'h3df20082} /* (7, 14, 22) {real, imag} */,
  {32'h3d486b98, 32'hbef5521a} /* (7, 14, 21) {real, imag} */,
  {32'h3e8de5f9, 32'hbd8b8bb8} /* (7, 14, 20) {real, imag} */,
  {32'hbe588c8a, 32'h3d875a36} /* (7, 14, 19) {real, imag} */,
  {32'hbf5e5060, 32'hbeac2a5a} /* (7, 14, 18) {real, imag} */,
  {32'h3e17e3bf, 32'hbda3a8a4} /* (7, 14, 17) {real, imag} */,
  {32'h3c231ee0, 32'h3e9d823d} /* (7, 14, 16) {real, imag} */,
  {32'hbe7baca8, 32'hbcf648d2} /* (7, 14, 15) {real, imag} */,
  {32'hbeb6d7f9, 32'h3eb84937} /* (7, 14, 14) {real, imag} */,
  {32'hbe54050a, 32'hbe86250e} /* (7, 14, 13) {real, imag} */,
  {32'h3c169d7c, 32'h3e5a4ded} /* (7, 14, 12) {real, imag} */,
  {32'hbda172fc, 32'hbe203442} /* (7, 14, 11) {real, imag} */,
  {32'h3e37e22e, 32'hbf13b553} /* (7, 14, 10) {real, imag} */,
  {32'hbec112f2, 32'h3ed49f0a} /* (7, 14, 9) {real, imag} */,
  {32'h3ddf5f28, 32'h3e4946fb} /* (7, 14, 8) {real, imag} */,
  {32'hbe8851d1, 32'h3d861c64} /* (7, 14, 7) {real, imag} */,
  {32'h3e0f65eb, 32'h3e737ed1} /* (7, 14, 6) {real, imag} */,
  {32'hbdfbcb5c, 32'h3ebd04bc} /* (7, 14, 5) {real, imag} */,
  {32'hbd9eeefe, 32'h3e726661} /* (7, 14, 4) {real, imag} */,
  {32'h3cd042fc, 32'hbd31ef7a} /* (7, 14, 3) {real, imag} */,
  {32'h3d950098, 32'hbd07f502} /* (7, 14, 2) {real, imag} */,
  {32'h3df510c3, 32'hbe8e3876} /* (7, 14, 1) {real, imag} */,
  {32'h3ce44210, 32'hbd436878} /* (7, 14, 0) {real, imag} */,
  {32'h3dfbd264, 32'h3f05c4a3} /* (7, 13, 31) {real, imag} */,
  {32'hbeb97424, 32'h3e37d039} /* (7, 13, 30) {real, imag} */,
  {32'h3e1206f4, 32'h3edb394b} /* (7, 13, 29) {real, imag} */,
  {32'h3d57359c, 32'h3d3b7c36} /* (7, 13, 28) {real, imag} */,
  {32'hbd56da74, 32'hbe63a6a2} /* (7, 13, 27) {real, imag} */,
  {32'h3ebc0425, 32'hbe5bd481} /* (7, 13, 26) {real, imag} */,
  {32'h3ed8c5ef, 32'h3d0015f7} /* (7, 13, 25) {real, imag} */,
  {32'hbe87782a, 32'hbea38236} /* (7, 13, 24) {real, imag} */,
  {32'hbe8b3242, 32'hbc256240} /* (7, 13, 23) {real, imag} */,
  {32'hbdb81c86, 32'hbda0c01a} /* (7, 13, 22) {real, imag} */,
  {32'hbeff6fb7, 32'hbd572648} /* (7, 13, 21) {real, imag} */,
  {32'hbedd9231, 32'hbea34ee2} /* (7, 13, 20) {real, imag} */,
  {32'h3f1c4835, 32'h3ec21c1e} /* (7, 13, 19) {real, imag} */,
  {32'hbf21e2a2, 32'hbe7aaa42} /* (7, 13, 18) {real, imag} */,
  {32'h3d47e5c8, 32'hbe3cbe55} /* (7, 13, 17) {real, imag} */,
  {32'h3e1a3d28, 32'hbeae913f} /* (7, 13, 16) {real, imag} */,
  {32'h3e89f7f2, 32'h3e38d96e} /* (7, 13, 15) {real, imag} */,
  {32'hbefb6811, 32'h3df04fe4} /* (7, 13, 14) {real, imag} */,
  {32'h3ec6b91e, 32'hbdcec295} /* (7, 13, 13) {real, imag} */,
  {32'h3e84509c, 32'h3f16d098} /* (7, 13, 12) {real, imag} */,
  {32'h3e074c6a, 32'h3efd1442} /* (7, 13, 11) {real, imag} */,
  {32'hbf079be7, 32'h3df2b803} /* (7, 13, 10) {real, imag} */,
  {32'hbe28f11e, 32'h3ea8b7c8} /* (7, 13, 9) {real, imag} */,
  {32'h3ca94f20, 32'hbea50654} /* (7, 13, 8) {real, imag} */,
  {32'h3e438365, 32'h3e218244} /* (7, 13, 7) {real, imag} */,
  {32'hbcf6df52, 32'h3d8752b4} /* (7, 13, 6) {real, imag} */,
  {32'h3e0277e3, 32'h3c49f240} /* (7, 13, 5) {real, imag} */,
  {32'hbd443800, 32'h3e3e6f38} /* (7, 13, 4) {real, imag} */,
  {32'hbca401dc, 32'h3f053e70} /* (7, 13, 3) {real, imag} */,
  {32'hbde4611e, 32'hbf052dee} /* (7, 13, 2) {real, imag} */,
  {32'h3dbd99d8, 32'hbd8d5caf} /* (7, 13, 1) {real, imag} */,
  {32'hbf7b397e, 32'h3e91f938} /* (7, 13, 0) {real, imag} */,
  {32'h3e3bbf3f, 32'hbdb8c002} /* (7, 12, 31) {real, imag} */,
  {32'hbdcd4a68, 32'hbbf120a0} /* (7, 12, 30) {real, imag} */,
  {32'h3d05e688, 32'h3e75f75c} /* (7, 12, 29) {real, imag} */,
  {32'hbec80d48, 32'h3ee1a35a} /* (7, 12, 28) {real, imag} */,
  {32'hbdb2bab4, 32'hbdace1da} /* (7, 12, 27) {real, imag} */,
  {32'h3e54237e, 32'h3eeb17d3} /* (7, 12, 26) {real, imag} */,
  {32'h3df383e4, 32'h3c25c390} /* (7, 12, 25) {real, imag} */,
  {32'hbe652549, 32'h3c4e9b38} /* (7, 12, 24) {real, imag} */,
  {32'h3dca60c8, 32'h3ee0a0d4} /* (7, 12, 23) {real, imag} */,
  {32'hbef37009, 32'hbd52ad0a} /* (7, 12, 22) {real, imag} */,
  {32'hbd749c70, 32'hbf0925ac} /* (7, 12, 21) {real, imag} */,
  {32'h3e50f5a6, 32'h3e7179f9} /* (7, 12, 20) {real, imag} */,
  {32'hbe982b34, 32'hbe9fc0a0} /* (7, 12, 19) {real, imag} */,
  {32'hbdb18f0a, 32'h3cd24c74} /* (7, 12, 18) {real, imag} */,
  {32'h3ec4dfd9, 32'h3cf52dd8} /* (7, 12, 17) {real, imag} */,
  {32'h3c7bdf68, 32'hbecb2b0a} /* (7, 12, 16) {real, imag} */,
  {32'hbdde01bc, 32'h3e253c40} /* (7, 12, 15) {real, imag} */,
  {32'h3e29b576, 32'h3edad8ec} /* (7, 12, 14) {real, imag} */,
  {32'hbec6d037, 32'h3eaf92d9} /* (7, 12, 13) {real, imag} */,
  {32'h3ed99a99, 32'hbca7eb98} /* (7, 12, 12) {real, imag} */,
  {32'hbdc75460, 32'hbe0fcab2} /* (7, 12, 11) {real, imag} */,
  {32'h3ecb822c, 32'h3f2ebbb2} /* (7, 12, 10) {real, imag} */,
  {32'hbee444bc, 32'hbd9f49a0} /* (7, 12, 9) {real, imag} */,
  {32'h3b3fd940, 32'h3e5a5c30} /* (7, 12, 8) {real, imag} */,
  {32'h3ee141d8, 32'hbe63025e} /* (7, 12, 7) {real, imag} */,
  {32'hbdb9d5a5, 32'h3ee2a084} /* (7, 12, 6) {real, imag} */,
  {32'hbf087442, 32'hbd8faf84} /* (7, 12, 5) {real, imag} */,
  {32'h3f10a7b4, 32'hbec0f98f} /* (7, 12, 4) {real, imag} */,
  {32'hbf1545bc, 32'hbe5505fb} /* (7, 12, 3) {real, imag} */,
  {32'h3d02cfe8, 32'hbde9a7a4} /* (7, 12, 2) {real, imag} */,
  {32'h3efbb391, 32'hbcf186dc} /* (7, 12, 1) {real, imag} */,
  {32'h3d075290, 32'hbd4e2638} /* (7, 12, 0) {real, imag} */,
  {32'h3c8e2b00, 32'hbe677718} /* (7, 11, 31) {real, imag} */,
  {32'h3f32056c, 32'h3ba6c680} /* (7, 11, 30) {real, imag} */,
  {32'h3e9bab4c, 32'h3eb335a0} /* (7, 11, 29) {real, imag} */,
  {32'hbeb28038, 32'hbe98b778} /* (7, 11, 28) {real, imag} */,
  {32'h3d661b48, 32'h3e85c4f9} /* (7, 11, 27) {real, imag} */,
  {32'h3e8b401b, 32'h3e50c105} /* (7, 11, 26) {real, imag} */,
  {32'hbf35b176, 32'hbde7affe} /* (7, 11, 25) {real, imag} */,
  {32'hbe6b2e5a, 32'h3ee1b4fe} /* (7, 11, 24) {real, imag} */,
  {32'hbf539410, 32'h3eec07e5} /* (7, 11, 23) {real, imag} */,
  {32'hbe15bd6e, 32'hbe85abdd} /* (7, 11, 22) {real, imag} */,
  {32'h3f0962ff, 32'hbe9918f2} /* (7, 11, 21) {real, imag} */,
  {32'h3f462406, 32'h3cd89b24} /* (7, 11, 20) {real, imag} */,
  {32'h3e47a9da, 32'hbc9864c8} /* (7, 11, 19) {real, imag} */,
  {32'h3eab4a7f, 32'h3e3352f6} /* (7, 11, 18) {real, imag} */,
  {32'hbe7a9f6b, 32'hbe053ebd} /* (7, 11, 17) {real, imag} */,
  {32'h3e9d38f0, 32'h3e0d4c9e} /* (7, 11, 16) {real, imag} */,
  {32'h3ea1e5d8, 32'h3e4cee7b} /* (7, 11, 15) {real, imag} */,
  {32'hbec4b906, 32'hbed244d0} /* (7, 11, 14) {real, imag} */,
  {32'hbd8808e4, 32'hbcabaec8} /* (7, 11, 13) {real, imag} */,
  {32'h3cef6e68, 32'hbec9e075} /* (7, 11, 12) {real, imag} */,
  {32'hbdf5e3b8, 32'h3eba6fa0} /* (7, 11, 11) {real, imag} */,
  {32'hbf0973e0, 32'h3f1d56b6} /* (7, 11, 10) {real, imag} */,
  {32'h3ec918f2, 32'hbf1376bf} /* (7, 11, 9) {real, imag} */,
  {32'hbd98252c, 32'h3e102c8e} /* (7, 11, 8) {real, imag} */,
  {32'h3e9dbd94, 32'h3e1d6376} /* (7, 11, 7) {real, imag} */,
  {32'h3e9bc99a, 32'h3f2789de} /* (7, 11, 6) {real, imag} */,
  {32'hbdbf3f74, 32'h3e89e67c} /* (7, 11, 5) {real, imag} */,
  {32'h3e4c5f40, 32'hbf32c1ce} /* (7, 11, 4) {real, imag} */,
  {32'h3ee543e2, 32'hbf377cc1} /* (7, 11, 3) {real, imag} */,
  {32'hbe169c6f, 32'h3f032e61} /* (7, 11, 2) {real, imag} */,
  {32'h3d4db350, 32'hbf517db1} /* (7, 11, 1) {real, imag} */,
  {32'hbea2e90c, 32'hbea458d1} /* (7, 11, 0) {real, imag} */,
  {32'hbc32af60, 32'h3e542cf5} /* (7, 10, 31) {real, imag} */,
  {32'hbec630ac, 32'h3e3d22a0} /* (7, 10, 30) {real, imag} */,
  {32'hbeb719f2, 32'hbec0d69b} /* (7, 10, 29) {real, imag} */,
  {32'h3cb10efc, 32'h3f05fc28} /* (7, 10, 28) {real, imag} */,
  {32'h3e8a3e92, 32'hbeda078d} /* (7, 10, 27) {real, imag} */,
  {32'h3e968c53, 32'hbe1623a9} /* (7, 10, 26) {real, imag} */,
  {32'h3dea54c2, 32'hbeffd1dc} /* (7, 10, 25) {real, imag} */,
  {32'hbed9c1e3, 32'h3e01fc71} /* (7, 10, 24) {real, imag} */,
  {32'h3e51ca1c, 32'hbe6a8bae} /* (7, 10, 23) {real, imag} */,
  {32'hbf156590, 32'hbe84fa9e} /* (7, 10, 22) {real, imag} */,
  {32'h3f56fd4b, 32'hbc9a2da0} /* (7, 10, 21) {real, imag} */,
  {32'h3f48129a, 32'h3ced4e20} /* (7, 10, 20) {real, imag} */,
  {32'h3e7647c9, 32'h3f0f47b8} /* (7, 10, 19) {real, imag} */,
  {32'hbde5f34c, 32'h3c6bb9f0} /* (7, 10, 18) {real, imag} */,
  {32'hbe894e9a, 32'hbe507b9e} /* (7, 10, 17) {real, imag} */,
  {32'hbbfc1ca0, 32'hbe58a611} /* (7, 10, 16) {real, imag} */,
  {32'hbd443ac6, 32'hbe25e844} /* (7, 10, 15) {real, imag} */,
  {32'hbecd89c3, 32'hbec21b37} /* (7, 10, 14) {real, imag} */,
  {32'h3ef1a90e, 32'hbe7572c3} /* (7, 10, 13) {real, imag} */,
  {32'h3e932994, 32'h3f0c2d91} /* (7, 10, 12) {real, imag} */,
  {32'h3e78ab78, 32'hbf29c9e2} /* (7, 10, 11) {real, imag} */,
  {32'hbecb8a6c, 32'h3dea8332} /* (7, 10, 10) {real, imag} */,
  {32'h3e59d1c7, 32'h3e3e809b} /* (7, 10, 9) {real, imag} */,
  {32'hbe00ef45, 32'hbddd1a5a} /* (7, 10, 8) {real, imag} */,
  {32'hbe44900e, 32'hbed2e7ee} /* (7, 10, 7) {real, imag} */,
  {32'hbea51743, 32'h3ec68402} /* (7, 10, 6) {real, imag} */,
  {32'h3f23294a, 32'hbe2dd336} /* (7, 10, 5) {real, imag} */,
  {32'hbd687f66, 32'hbd4cdc9c} /* (7, 10, 4) {real, imag} */,
  {32'hbe3bae5b, 32'h3f25982e} /* (7, 10, 3) {real, imag} */,
  {32'h3d02fdbc, 32'hbebcd440} /* (7, 10, 2) {real, imag} */,
  {32'h3f0882a9, 32'hbe15d1f6} /* (7, 10, 1) {real, imag} */,
  {32'hbdeb884c, 32'h3f52b5c6} /* (7, 10, 0) {real, imag} */,
  {32'hbec7f4f4, 32'h3f48ff99} /* (7, 9, 31) {real, imag} */,
  {32'h3edf4c0a, 32'hbf33a7da} /* (7, 9, 30) {real, imag} */,
  {32'hbcb4d3a8, 32'hbc870108} /* (7, 9, 29) {real, imag} */,
  {32'hbd018f2a, 32'h3c3bfb90} /* (7, 9, 28) {real, imag} */,
  {32'hbee8ea77, 32'h3e70daf6} /* (7, 9, 27) {real, imag} */,
  {32'h3d678818, 32'hbe3594ca} /* (7, 9, 26) {real, imag} */,
  {32'hbf0c599b, 32'hbe2cb604} /* (7, 9, 25) {real, imag} */,
  {32'h3e3a57d0, 32'hbed76f5c} /* (7, 9, 24) {real, imag} */,
  {32'hbf0d934e, 32'hbf08890a} /* (7, 9, 23) {real, imag} */,
  {32'h3f293f92, 32'hbe2e5ddf} /* (7, 9, 22) {real, imag} */,
  {32'hbcc3aa10, 32'hbe95329b} /* (7, 9, 21) {real, imag} */,
  {32'h3d918b70, 32'hbdd6a280} /* (7, 9, 20) {real, imag} */,
  {32'h3eed8db2, 32'h3eb7a2ad} /* (7, 9, 19) {real, imag} */,
  {32'hbef6a155, 32'hbe2e0d62} /* (7, 9, 18) {real, imag} */,
  {32'h3dfef25a, 32'h3e72c3b0} /* (7, 9, 17) {real, imag} */,
  {32'h3dd9950a, 32'h3e8b14f2} /* (7, 9, 16) {real, imag} */,
  {32'h3e040bd2, 32'hbea91a2e} /* (7, 9, 15) {real, imag} */,
  {32'h3e81c450, 32'h3d9c057d} /* (7, 9, 14) {real, imag} */,
  {32'hbd83aa64, 32'hbed94fea} /* (7, 9, 13) {real, imag} */,
  {32'h3db8f8d8, 32'h3e262cc7} /* (7, 9, 12) {real, imag} */,
  {32'h3e8f7d66, 32'h3d048a34} /* (7, 9, 11) {real, imag} */,
  {32'h3e71f827, 32'hbe50a882} /* (7, 9, 10) {real, imag} */,
  {32'hbea5075c, 32'h3f2dd430} /* (7, 9, 9) {real, imag} */,
  {32'hbdf344c6, 32'hbdb57eaa} /* (7, 9, 8) {real, imag} */,
  {32'h3d01b375, 32'h3f009196} /* (7, 9, 7) {real, imag} */,
  {32'hbee34717, 32'hbe738c0e} /* (7, 9, 6) {real, imag} */,
  {32'hbe1c122e, 32'h3eb099cb} /* (7, 9, 5) {real, imag} */,
  {32'h3e83b555, 32'h3e7d0e40} /* (7, 9, 4) {real, imag} */,
  {32'hbd90ddc5, 32'h3eaa54ab} /* (7, 9, 3) {real, imag} */,
  {32'hbefc6eb4, 32'hbe10460c} /* (7, 9, 2) {real, imag} */,
  {32'hbf23e8b2, 32'h3d353f94} /* (7, 9, 1) {real, imag} */,
  {32'hbe8cab70, 32'hbe2a75bb} /* (7, 9, 0) {real, imag} */,
  {32'hbfc45dc3, 32'hbf30f6f4} /* (7, 8, 31) {real, imag} */,
  {32'h3f67772d, 32'h3f0daf33} /* (7, 8, 30) {real, imag} */,
  {32'h3e82b91c, 32'hbe8acfe4} /* (7, 8, 29) {real, imag} */,
  {32'h3ed69b50, 32'h3df7efea} /* (7, 8, 28) {real, imag} */,
  {32'h3f7b1944, 32'hbed9517a} /* (7, 8, 27) {real, imag} */,
  {32'h3ea100f8, 32'hbec3c935} /* (7, 8, 26) {real, imag} */,
  {32'hbe8ed724, 32'hbedbc6aa} /* (7, 8, 25) {real, imag} */,
  {32'h3eda3f11, 32'hbf340aad} /* (7, 8, 24) {real, imag} */,
  {32'h3e800960, 32'hbef33d78} /* (7, 8, 23) {real, imag} */,
  {32'h3d17da88, 32'h3cd96878} /* (7, 8, 22) {real, imag} */,
  {32'hbe33c6bd, 32'h3ed468ce} /* (7, 8, 21) {real, imag} */,
  {32'hbe50db5c, 32'h3f0be5fb} /* (7, 8, 20) {real, imag} */,
  {32'hbe01fc1c, 32'h3d1fc260} /* (7, 8, 19) {real, imag} */,
  {32'h3eae1656, 32'h3e91e712} /* (7, 8, 18) {real, imag} */,
  {32'hbf05b17a, 32'h3e91e174} /* (7, 8, 17) {real, imag} */,
  {32'hbe8cce62, 32'h3e0cbf28} /* (7, 8, 16) {real, imag} */,
  {32'h3e0c8756, 32'hbeafee88} /* (7, 8, 15) {real, imag} */,
  {32'h3f2bd7d9, 32'hbe9d457a} /* (7, 8, 14) {real, imag} */,
  {32'hbf2678ba, 32'h3e2b537b} /* (7, 8, 13) {real, imag} */,
  {32'hbd93d438, 32'hbe00b5a3} /* (7, 8, 12) {real, imag} */,
  {32'h3dec51f4, 32'h3f1448a2} /* (7, 8, 11) {real, imag} */,
  {32'h3e7224d9, 32'hbe327aeb} /* (7, 8, 10) {real, imag} */,
  {32'hbefc6ebc, 32'hbeb580c1} /* (7, 8, 9) {real, imag} */,
  {32'hbe02bea0, 32'h3f6d49e8} /* (7, 8, 8) {real, imag} */,
  {32'hbed62194, 32'h3e42a799} /* (7, 8, 7) {real, imag} */,
  {32'hbf039bc4, 32'h3d2ab288} /* (7, 8, 6) {real, imag} */,
  {32'hbf0a9c0a, 32'h3dc1f356} /* (7, 8, 5) {real, imag} */,
  {32'hbef51275, 32'hbf0353c9} /* (7, 8, 4) {real, imag} */,
  {32'h3e271798, 32'h3e79c8ad} /* (7, 8, 3) {real, imag} */,
  {32'h3f2bc60a, 32'h3e1a63d8} /* (7, 8, 2) {real, imag} */,
  {32'hbf05bea2, 32'hbf88ba72} /* (7, 8, 1) {real, imag} */,
  {32'hbf559ae1, 32'hbf1d5430} /* (7, 8, 0) {real, imag} */,
  {32'hbe0097ac, 32'hbe83c292} /* (7, 7, 31) {real, imag} */,
  {32'h3e8b396a, 32'hbe0d12c4} /* (7, 7, 30) {real, imag} */,
  {32'hbf41cbe2, 32'h3e02e6f2} /* (7, 7, 29) {real, imag} */,
  {32'hbd977096, 32'h3e2f4bf6} /* (7, 7, 28) {real, imag} */,
  {32'h3e8b9255, 32'hbe289574} /* (7, 7, 27) {real, imag} */,
  {32'hbd6c870c, 32'h3ef1a2a0} /* (7, 7, 26) {real, imag} */,
  {32'hbe987117, 32'h3f47916c} /* (7, 7, 25) {real, imag} */,
  {32'h3e994be8, 32'hbe894afa} /* (7, 7, 24) {real, imag} */,
  {32'hbe8e9fde, 32'hbe3e0516} /* (7, 7, 23) {real, imag} */,
  {32'hbe501160, 32'h3dafb3ab} /* (7, 7, 22) {real, imag} */,
  {32'h3df0ce72, 32'hbeb7e75b} /* (7, 7, 21) {real, imag} */,
  {32'hbd2041be, 32'h3e017d28} /* (7, 7, 20) {real, imag} */,
  {32'hbd2bb8d8, 32'h3e67849d} /* (7, 7, 19) {real, imag} */,
  {32'h3deeb45a, 32'hbd9364be} /* (7, 7, 18) {real, imag} */,
  {32'hbe7390a4, 32'h3d9b40ee} /* (7, 7, 17) {real, imag} */,
  {32'hbe34ef65, 32'hbe037ec5} /* (7, 7, 16) {real, imag} */,
  {32'hbc0aacd8, 32'hbe2205ee} /* (7, 7, 15) {real, imag} */,
  {32'h3dded06a, 32'hbe77b616} /* (7, 7, 14) {real, imag} */,
  {32'h3e12eede, 32'h3ed51574} /* (7, 7, 13) {real, imag} */,
  {32'hbe666e14, 32'hbf0a44c0} /* (7, 7, 12) {real, imag} */,
  {32'hbed81164, 32'h3ca11a40} /* (7, 7, 11) {real, imag} */,
  {32'h3f3be576, 32'h3ed6a8b7} /* (7, 7, 10) {real, imag} */,
  {32'h3edbee02, 32'h3f48148e} /* (7, 7, 9) {real, imag} */,
  {32'hbf07e855, 32'hbea1c52c} /* (7, 7, 8) {real, imag} */,
  {32'hbe83307d, 32'hbf2f7cd4} /* (7, 7, 7) {real, imag} */,
  {32'h3f276907, 32'h3dfb301c} /* (7, 7, 6) {real, imag} */,
  {32'h3f96df1b, 32'hbe8c6c8e} /* (7, 7, 5) {real, imag} */,
  {32'h3e2eee4c, 32'h3f42c4ed} /* (7, 7, 4) {real, imag} */,
  {32'hbed8e1a7, 32'h3f4ae47e} /* (7, 7, 3) {real, imag} */,
  {32'hbe17c106, 32'hbf917784} /* (7, 7, 2) {real, imag} */,
  {32'hbe5d6c84, 32'h3f1536a7} /* (7, 7, 1) {real, imag} */,
  {32'h3edc6cf6, 32'h3e880cec} /* (7, 7, 0) {real, imag} */,
  {32'h3e533625, 32'h3f0933b2} /* (7, 6, 31) {real, imag} */,
  {32'hbdd8836c, 32'hbecc5e3d} /* (7, 6, 30) {real, imag} */,
  {32'hbe1780cf, 32'hbee6be86} /* (7, 6, 29) {real, imag} */,
  {32'hbe7ac502, 32'h3edcfbeb} /* (7, 6, 28) {real, imag} */,
  {32'h3f15b2eb, 32'h3f0ca3a8} /* (7, 6, 27) {real, imag} */,
  {32'hbdd01ac8, 32'hbb8b0f80} /* (7, 6, 26) {real, imag} */,
  {32'h3ef6317a, 32'h3c982130} /* (7, 6, 25) {real, imag} */,
  {32'h3d6e5368, 32'hbe9bad3f} /* (7, 6, 24) {real, imag} */,
  {32'h3f1449ef, 32'hbe464a8b} /* (7, 6, 23) {real, imag} */,
  {32'hbe120264, 32'h3de8ad34} /* (7, 6, 22) {real, imag} */,
  {32'hbe52eb6b, 32'hbe16b662} /* (7, 6, 21) {real, imag} */,
  {32'h3d20ae34, 32'hbe422b18} /* (7, 6, 20) {real, imag} */,
  {32'hbe306ddb, 32'h3e99f858} /* (7, 6, 19) {real, imag} */,
  {32'hbe38ec60, 32'h3dc02754} /* (7, 6, 18) {real, imag} */,
  {32'hbda3ccdf, 32'h3e1dfd7f} /* (7, 6, 17) {real, imag} */,
  {32'hbebcde08, 32'hbe4460b1} /* (7, 6, 16) {real, imag} */,
  {32'hbe27d23e, 32'hbc1f0050} /* (7, 6, 15) {real, imag} */,
  {32'hbe835005, 32'h3ea0de34} /* (7, 6, 14) {real, imag} */,
  {32'h3e23694b, 32'hbe55c90a} /* (7, 6, 13) {real, imag} */,
  {32'hbe7fb441, 32'h3eeb2218} /* (7, 6, 12) {real, imag} */,
  {32'h3ea3c58f, 32'hbe9b1729} /* (7, 6, 11) {real, imag} */,
  {32'h3da55ca0, 32'hbea80a7c} /* (7, 6, 10) {real, imag} */,
  {32'hbed4eb66, 32'hbe1182ce} /* (7, 6, 9) {real, imag} */,
  {32'h3ede53c4, 32'hbe109405} /* (7, 6, 8) {real, imag} */,
  {32'h3f693bd0, 32'h3ee61d14} /* (7, 6, 7) {real, imag} */,
  {32'hbe3ccbb8, 32'hbd894240} /* (7, 6, 6) {real, imag} */,
  {32'hbdaecab3, 32'h3db08da5} /* (7, 6, 5) {real, imag} */,
  {32'h3d99aa8d, 32'h3d3934b0} /* (7, 6, 4) {real, imag} */,
  {32'hbeaf9bba, 32'h3f5075a5} /* (7, 6, 3) {real, imag} */,
  {32'hbf5113e2, 32'hbe6c2cf0} /* (7, 6, 2) {real, imag} */,
  {32'hbf13b9d5, 32'h3e69946b} /* (7, 6, 1) {real, imag} */,
  {32'hbd75e64c, 32'hbebb646a} /* (7, 6, 0) {real, imag} */,
  {32'hc02473b8, 32'h3de037e4} /* (7, 5, 31) {real, imag} */,
  {32'h3fceb1ae, 32'hbf8b7256} /* (7, 5, 30) {real, imag} */,
  {32'hbdfba380, 32'hbe30f9c2} /* (7, 5, 29) {real, imag} */,
  {32'hbec22102, 32'h3dfd4d28} /* (7, 5, 28) {real, imag} */,
  {32'h3eb6d98f, 32'hbea258a2} /* (7, 5, 27) {real, imag} */,
  {32'hbe8ab28a, 32'h3e0fe854} /* (7, 5, 26) {real, imag} */,
  {32'hbeea7a8e, 32'h3e430939} /* (7, 5, 25) {real, imag} */,
  {32'h3b616da0, 32'hbec34b04} /* (7, 5, 24) {real, imag} */,
  {32'hbe53c55e, 32'hbe8d5f4a} /* (7, 5, 23) {real, imag} */,
  {32'h3e53d02f, 32'h3db71ad8} /* (7, 5, 22) {real, imag} */,
  {32'h3e9e0cba, 32'h3e61ff8f} /* (7, 5, 21) {real, imag} */,
  {32'hbde91f84, 32'hbe0f2456} /* (7, 5, 20) {real, imag} */,
  {32'h3e8f3b08, 32'hbd4e455a} /* (7, 5, 19) {real, imag} */,
  {32'hbe63b8c2, 32'hbee4fb40} /* (7, 5, 18) {real, imag} */,
  {32'h3df10008, 32'hbb236d90} /* (7, 5, 17) {real, imag} */,
  {32'h3e132f00, 32'hbea58512} /* (7, 5, 16) {real, imag} */,
  {32'hbe6a741d, 32'hbdf18934} /* (7, 5, 15) {real, imag} */,
  {32'hbf145932, 32'h3e0eedc1} /* (7, 5, 14) {real, imag} */,
  {32'hbd3eb399, 32'hbe9f3793} /* (7, 5, 13) {real, imag} */,
  {32'h3d9296a0, 32'hbeb17fe6} /* (7, 5, 12) {real, imag} */,
  {32'hbf0e6e03, 32'hbe6dddd6} /* (7, 5, 11) {real, imag} */,
  {32'h3e3d048e, 32'hbee79b66} /* (7, 5, 10) {real, imag} */,
  {32'h3e51ea63, 32'h3c9bcab8} /* (7, 5, 9) {real, imag} */,
  {32'h3e135f5c, 32'hbeab7649} /* (7, 5, 8) {real, imag} */,
  {32'hbea6cc80, 32'h3e2de43c} /* (7, 5, 7) {real, imag} */,
  {32'h3f207657, 32'h3f02c462} /* (7, 5, 6) {real, imag} */,
  {32'h3f34209c, 32'h3ea71331} /* (7, 5, 5) {real, imag} */,
  {32'h3cb8c840, 32'h3dbd9c08} /* (7, 5, 4) {real, imag} */,
  {32'hbdaea4b0, 32'h3bd7ca00} /* (7, 5, 3) {real, imag} */,
  {32'h3fabcdc6, 32'h3f95d816} /* (7, 5, 2) {real, imag} */,
  {32'hbfa45525, 32'hbf46695a} /* (7, 5, 1) {real, imag} */,
  {32'hc011524c, 32'hbf514b9c} /* (7, 5, 0) {real, imag} */,
  {32'h3e975e9a, 32'h402cb87c} /* (7, 4, 31) {real, imag} */,
  {32'hc0285c1c, 32'hc006f907} /* (7, 4, 30) {real, imag} */,
  {32'h3e957314, 32'hbf06ddf6} /* (7, 4, 29) {real, imag} */,
  {32'h3f93734a, 32'h3e6b6c8a} /* (7, 4, 28) {real, imag} */,
  {32'hbe6b7eb1, 32'hbddc04f6} /* (7, 4, 27) {real, imag} */,
  {32'hbec9cb68, 32'hbdcfe96c} /* (7, 4, 26) {real, imag} */,
  {32'h3e268ac1, 32'h3dc40a28} /* (7, 4, 25) {real, imag} */,
  {32'hbd6feb08, 32'hbf1b9cba} /* (7, 4, 24) {real, imag} */,
  {32'hbea0e940, 32'hbea4124b} /* (7, 4, 23) {real, imag} */,
  {32'h3edb850a, 32'hbe007bca} /* (7, 4, 22) {real, imag} */,
  {32'h3dabc3fe, 32'hbf260e9b} /* (7, 4, 21) {real, imag} */,
  {32'hbe1e878a, 32'h3f2416ee} /* (7, 4, 20) {real, imag} */,
  {32'hbd864640, 32'h3ed8e026} /* (7, 4, 19) {real, imag} */,
  {32'hbe8b6e3d, 32'hbe54d238} /* (7, 4, 18) {real, imag} */,
  {32'h3ebee65c, 32'h3be689e0} /* (7, 4, 17) {real, imag} */,
  {32'h3c32f91e, 32'h3e4e1870} /* (7, 4, 16) {real, imag} */,
  {32'hbed00cd0, 32'h3e4ed7ab} /* (7, 4, 15) {real, imag} */,
  {32'hbef5f890, 32'hbe41ae46} /* (7, 4, 14) {real, imag} */,
  {32'h3ee76cc0, 32'h3de738e8} /* (7, 4, 13) {real, imag} */,
  {32'hbe6c5af8, 32'h3e4475a4} /* (7, 4, 12) {real, imag} */,
  {32'h3e746279, 32'hbefabb78} /* (7, 4, 11) {real, imag} */,
  {32'h3de7b9ff, 32'hbd283df4} /* (7, 4, 10) {real, imag} */,
  {32'h3ee88ac6, 32'hbf29b961} /* (7, 4, 9) {real, imag} */,
  {32'hbe66e362, 32'hbf168b22} /* (7, 4, 8) {real, imag} */,
  {32'hbd7fc7d0, 32'h3c8f5dc0} /* (7, 4, 7) {real, imag} */,
  {32'h3e830cb3, 32'h3eac2d98} /* (7, 4, 6) {real, imag} */,
  {32'hbcdedd60, 32'hbf91f9ac} /* (7, 4, 5) {real, imag} */,
  {32'h3e6be8f6, 32'h3fa712dd} /* (7, 4, 4) {real, imag} */,
  {32'hbf05c3a1, 32'hbd2f91d4} /* (7, 4, 3) {real, imag} */,
  {32'hc0190dcb, 32'hc02b1fba} /* (7, 4, 2) {real, imag} */,
  {32'h407063b8, 32'h40457a32} /* (7, 4, 1) {real, imag} */,
  {32'h3fecdcee, 32'h3de8c630} /* (7, 4, 0) {real, imag} */,
  {32'hc08efc8b, 32'h3fdd5adc} /* (7, 3, 31) {real, imag} */,
  {32'h3ff0769c, 32'hc06ccdb2} /* (7, 3, 30) {real, imag} */,
  {32'hbee905a8, 32'hbd08cbd0} /* (7, 3, 29) {real, imag} */,
  {32'h3fa71c10, 32'h3f4aaf40} /* (7, 3, 28) {real, imag} */,
  {32'hbdd8e7a2, 32'h3e8c36d4} /* (7, 3, 27) {real, imag} */,
  {32'hbf3852fa, 32'hbdb55df0} /* (7, 3, 26) {real, imag} */,
  {32'hbf40829c, 32'h3f18d497} /* (7, 3, 25) {real, imag} */,
  {32'hbf37a790, 32'hbf337252} /* (7, 3, 24) {real, imag} */,
  {32'h3d560968, 32'h3b4c3340} /* (7, 3, 23) {real, imag} */,
  {32'h3c2d01e8, 32'h3dda4ed5} /* (7, 3, 22) {real, imag} */,
  {32'h3dd3417b, 32'hbf0785b6} /* (7, 3, 21) {real, imag} */,
  {32'hbeac9c55, 32'hbdf810d4} /* (7, 3, 20) {real, imag} */,
  {32'h3f0b3650, 32'h3e3e71e4} /* (7, 3, 19) {real, imag} */,
  {32'h3c3af8d0, 32'hbe7f8842} /* (7, 3, 18) {real, imag} */,
  {32'hbdace640, 32'h3bd2f7e0} /* (7, 3, 17) {real, imag} */,
  {32'h3d1c0f3c, 32'hbeb20dcc} /* (7, 3, 16) {real, imag} */,
  {32'h3dcc3cc8, 32'h3e0c597a} /* (7, 3, 15) {real, imag} */,
  {32'h3ef04e0a, 32'h3e9f7362} /* (7, 3, 14) {real, imag} */,
  {32'hbe44cb0a, 32'hbddc5322} /* (7, 3, 13) {real, imag} */,
  {32'h3cddf110, 32'hbee98afb} /* (7, 3, 12) {real, imag} */,
  {32'hbe437236, 32'hbf24e890} /* (7, 3, 11) {real, imag} */,
  {32'hbd38eaf2, 32'hbd520ec0} /* (7, 3, 10) {real, imag} */,
  {32'h3e5684a1, 32'h3eef3847} /* (7, 3, 9) {real, imag} */,
  {32'hbe1f597f, 32'h3ea916c2} /* (7, 3, 8) {real, imag} */,
  {32'hbde4a047, 32'h3e1ebce2} /* (7, 3, 7) {real, imag} */,
  {32'h3da4ca54, 32'hbeae0949} /* (7, 3, 6) {real, imag} */,
  {32'h3f7de1fa, 32'hbe1b275c} /* (7, 3, 5) {real, imag} */,
  {32'hbfc3bbb3, 32'h3f362de3} /* (7, 3, 4) {real, imag} */,
  {32'hbe2802b7, 32'hbe8ff03a} /* (7, 3, 3) {real, imag} */,
  {32'hbf29105c, 32'hbfe1f7be} /* (7, 3, 2) {real, imag} */,
  {32'h40843c7c, 32'h40857b78} /* (7, 3, 1) {real, imag} */,
  {32'h3f32150d, 32'h3e87d89d} /* (7, 3, 0) {real, imag} */,
  {32'hc1fc0336, 32'h3f08d424} /* (7, 2, 31) {real, imag} */,
  {32'h41744116, 32'hc0849647} /* (7, 2, 30) {real, imag} */,
  {32'hbfc1ec25, 32'h3fc9bce9} /* (7, 2, 29) {real, imag} */,
  {32'hbe3c7818, 32'h3fa50f79} /* (7, 2, 28) {real, imag} */,
  {32'h3fb5edfc, 32'hbf969f3e} /* (7, 2, 27) {real, imag} */,
  {32'h3f17941f, 32'hbeb919e7} /* (7, 2, 26) {real, imag} */,
  {32'hbf1e8dac, 32'h3dee44a0} /* (7, 2, 25) {real, imag} */,
  {32'h3f7d0b22, 32'h3e8b4666} /* (7, 2, 24) {real, imag} */,
  {32'h3e6886ca, 32'hbe244ae9} /* (7, 2, 23) {real, imag} */,
  {32'h3f2d37ac, 32'h3f312e16} /* (7, 2, 22) {real, imag} */,
  {32'h3f067f99, 32'hbe0ce1fb} /* (7, 2, 21) {real, imag} */,
  {32'h3f013f15, 32'hbf0553c3} /* (7, 2, 20) {real, imag} */,
  {32'hbe17bc02, 32'h3c8d77c0} /* (7, 2, 19) {real, imag} */,
  {32'h3da5f04c, 32'hbe7a5f60} /* (7, 2, 18) {real, imag} */,
  {32'hbb200920, 32'h3d342c24} /* (7, 2, 17) {real, imag} */,
  {32'hbdd779f8, 32'h3df4dd6a} /* (7, 2, 16) {real, imag} */,
  {32'h3ea490e8, 32'h3e522017} /* (7, 2, 15) {real, imag} */,
  {32'h3e8ca669, 32'hbe902aaf} /* (7, 2, 14) {real, imag} */,
  {32'hbf0bbdb3, 32'hbcc94fd0} /* (7, 2, 13) {real, imag} */,
  {32'hbf046e42, 32'h3eabe0dc} /* (7, 2, 12) {real, imag} */,
  {32'h3ef320d2, 32'h3ec73896} /* (7, 2, 11) {real, imag} */,
  {32'h3e9e3bfc, 32'h3c12d3a0} /* (7, 2, 10) {real, imag} */,
  {32'h3e7dfff3, 32'h3f2d5409} /* (7, 2, 9) {real, imag} */,
  {32'hbdca8438, 32'h3e66ec32} /* (7, 2, 8) {real, imag} */,
  {32'hbe546ab6, 32'hbf2bb5e4} /* (7, 2, 7) {real, imag} */,
  {32'h3e94d677, 32'h3d1d75c8} /* (7, 2, 6) {real, imag} */,
  {32'h3fda86e0, 32'h3f90dd2d} /* (7, 2, 5) {real, imag} */,
  {32'hc06d82c2, 32'hbf245c96} /* (7, 2, 4) {real, imag} */,
  {32'hbf6510e5, 32'h3f86f27a} /* (7, 2, 3) {real, imag} */,
  {32'h413fb028, 32'hbfd2eee3} /* (7, 2, 2) {real, imag} */,
  {32'hc181a06e, 32'h40400cee} /* (7, 2, 1) {real, imag} */,
  {32'hc1820d36, 32'hc0b5fa66} /* (7, 2, 0) {real, imag} */,
  {32'h4224cfda, 32'hc12909f4} /* (7, 1, 31) {real, imag} */,
  {32'hc109f35d, 32'h3f981785} /* (7, 1, 30) {real, imag} */,
  {32'h3fb125cc, 32'hbf9fd7f0} /* (7, 1, 29) {real, imag} */,
  {32'h3fd2bdee, 32'h400425f4} /* (7, 1, 28) {real, imag} */,
  {32'hc03cfb34, 32'h3ccd7808} /* (7, 1, 27) {real, imag} */,
  {32'hbf18a781, 32'h3f66c1b7} /* (7, 1, 26) {real, imag} */,
  {32'h3e941749, 32'hbdd14667} /* (7, 1, 25) {real, imag} */,
  {32'hbf45bb0f, 32'h3f4386b2} /* (7, 1, 24) {real, imag} */,
  {32'h3e23d984, 32'h3e770729} /* (7, 1, 23) {real, imag} */,
  {32'h3f1bf955, 32'hbe10a892} /* (7, 1, 22) {real, imag} */,
  {32'hbe97b321, 32'h3f74c342} /* (7, 1, 21) {real, imag} */,
  {32'h3c943e00, 32'h3e0934b4} /* (7, 1, 20) {real, imag} */,
  {32'h3da5fd46, 32'h3e839e28} /* (7, 1, 19) {real, imag} */,
  {32'h3d0eb8f4, 32'h3f294be0} /* (7, 1, 18) {real, imag} */,
  {32'hbe6c9447, 32'h3c2b8dd8} /* (7, 1, 17) {real, imag} */,
  {32'hbc730e68, 32'hbf094ed0} /* (7, 1, 16) {real, imag} */,
  {32'hbdd8398b, 32'h3e70c7a2} /* (7, 1, 15) {real, imag} */,
  {32'hbe9d4807, 32'h3dcd7a80} /* (7, 1, 14) {real, imag} */,
  {32'hbebeed78, 32'hbeac31bb} /* (7, 1, 13) {real, imag} */,
  {32'h3d1a5122, 32'hbe9f9a44} /* (7, 1, 12) {real, imag} */,
  {32'hbf0baf35, 32'hbef3dd65} /* (7, 1, 11) {real, imag} */,
  {32'hbe231a3c, 32'h3ea874cf} /* (7, 1, 10) {real, imag} */,
  {32'hbe8ef8eb, 32'h3d7e84c2} /* (7, 1, 9) {real, imag} */,
  {32'hbee5b8e3, 32'hbfa474f4} /* (7, 1, 8) {real, imag} */,
  {32'h3f046d3d, 32'h3f2afaa4} /* (7, 1, 7) {real, imag} */,
  {32'hbf2184f3, 32'hbd6e1918} /* (7, 1, 6) {real, imag} */,
  {32'hc0147832, 32'hbf851748} /* (7, 1, 5) {real, imag} */,
  {32'h3fc5eefc, 32'hbed82628} /* (7, 1, 4) {real, imag} */,
  {32'hbfb3fe73, 32'hc03ea9b8} /* (7, 1, 3) {real, imag} */,
  {32'hc1686dfe, 32'hc166db87} /* (7, 1, 2) {real, imag} */,
  {32'h42646005, 32'h41dac369} /* (7, 1, 1) {real, imag} */,
  {32'h425eaf4e, 32'h40e99daf} /* (7, 1, 0) {real, imag} */,
  {32'h42046afa, 32'hc1db6a80} /* (7, 0, 31) {real, imag} */,
  {32'hc04eac6a, 32'h410336f2} /* (7, 0, 30) {real, imag} */,
  {32'hbe0e4fcc, 32'hbf33fe6b} /* (7, 0, 29) {real, imag} */,
  {32'h3ee35448, 32'h3dfd0fa0} /* (7, 0, 28) {real, imag} */,
  {32'hbfff0831, 32'h3f516c1a} /* (7, 0, 27) {real, imag} */,
  {32'h3dbf935e, 32'h3ec30877} /* (7, 0, 26) {real, imag} */,
  {32'h3eef6a72, 32'hbfb195fa} /* (7, 0, 25) {real, imag} */,
  {32'hbf0874d8, 32'h3d760830} /* (7, 0, 24) {real, imag} */,
  {32'h3eab376c, 32'hbdd520a8} /* (7, 0, 23) {real, imag} */,
  {32'hbed145dc, 32'h3dc0b683} /* (7, 0, 22) {real, imag} */,
  {32'hbeaf2eea, 32'h3eab4290} /* (7, 0, 21) {real, imag} */,
  {32'h3d4057d8, 32'hbf19f9a7} /* (7, 0, 20) {real, imag} */,
  {32'h3da45ecc, 32'hbc947a5c} /* (7, 0, 19) {real, imag} */,
  {32'h3e36ba40, 32'h3f01ca2b} /* (7, 0, 18) {real, imag} */,
  {32'h3e0432d0, 32'hbe529cc9} /* (7, 0, 17) {real, imag} */,
  {32'hbe207d94, 32'h00000000} /* (7, 0, 16) {real, imag} */,
  {32'h3e0432d0, 32'h3e529cc9} /* (7, 0, 15) {real, imag} */,
  {32'h3e36ba40, 32'hbf01ca2b} /* (7, 0, 14) {real, imag} */,
  {32'h3da45ecc, 32'h3c947a5c} /* (7, 0, 13) {real, imag} */,
  {32'h3d4057d8, 32'h3f19f9a7} /* (7, 0, 12) {real, imag} */,
  {32'hbeaf2eea, 32'hbeab4290} /* (7, 0, 11) {real, imag} */,
  {32'hbed145dc, 32'hbdc0b683} /* (7, 0, 10) {real, imag} */,
  {32'h3eab376c, 32'h3dd520a8} /* (7, 0, 9) {real, imag} */,
  {32'hbf0874d8, 32'hbd760830} /* (7, 0, 8) {real, imag} */,
  {32'h3eef6a72, 32'h3fb195fa} /* (7, 0, 7) {real, imag} */,
  {32'h3dbf935e, 32'hbec30877} /* (7, 0, 6) {real, imag} */,
  {32'hbfff0831, 32'hbf516c1a} /* (7, 0, 5) {real, imag} */,
  {32'h3ee35448, 32'hbdfd0fa0} /* (7, 0, 4) {real, imag} */,
  {32'hbe0e4fcc, 32'h3f33fe6b} /* (7, 0, 3) {real, imag} */,
  {32'hc04eac6a, 32'hc10336f2} /* (7, 0, 2) {real, imag} */,
  {32'h42046afa, 32'h41db6a80} /* (7, 0, 1) {real, imag} */,
  {32'h42718902, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h421cbd4a, 32'hc1881355} /* (6, 31, 31) {real, imag} */,
  {32'hc124e64a, 32'h411b9bf8} /* (6, 31, 30) {real, imag} */,
  {32'hbf2575ee, 32'h4007893d} /* (6, 31, 29) {real, imag} */,
  {32'h3fc182cd, 32'h3f5536de} /* (6, 31, 28) {real, imag} */,
  {32'hbff02b8e, 32'h3e98e236} /* (6, 31, 27) {real, imag} */,
  {32'hbef51b62, 32'h3d1dba94} /* (6, 31, 26) {real, imag} */,
  {32'h3f430ac0, 32'hbe626ffa} /* (6, 31, 25) {real, imag} */,
  {32'hbea4d526, 32'h3f86c0c2} /* (6, 31, 24) {real, imag} */,
  {32'h3eae01e9, 32'h3b8a9480} /* (6, 31, 23) {real, imag} */,
  {32'hbe9af5bc, 32'h3d8c86b1} /* (6, 31, 22) {real, imag} */,
  {32'hbf1db160, 32'h3f3e8369} /* (6, 31, 21) {real, imag} */,
  {32'hbd90ba32, 32'hbd48daac} /* (6, 31, 20) {real, imag} */,
  {32'h3c2fa580, 32'hbd3ad3db} /* (6, 31, 19) {real, imag} */,
  {32'h3e8d0e80, 32'h3f007478} /* (6, 31, 18) {real, imag} */,
  {32'hbea13968, 32'hbda5f118} /* (6, 31, 17) {real, imag} */,
  {32'hbe6b0cce, 32'hbdde0e18} /* (6, 31, 16) {real, imag} */,
  {32'h3dcb5712, 32'hbde78f7a} /* (6, 31, 15) {real, imag} */,
  {32'hbef69b04, 32'hbe055a8b} /* (6, 31, 14) {real, imag} */,
  {32'h3d9c0e6e, 32'h3e826814} /* (6, 31, 13) {real, imag} */,
  {32'h3eebc1d6, 32'hbe3de156} /* (6, 31, 12) {real, imag} */,
  {32'hbf2b8a8c, 32'hbf80b772} /* (6, 31, 11) {real, imag} */,
  {32'h3eaf1eac, 32'h3e73cda2} /* (6, 31, 10) {real, imag} */,
  {32'h3d492f8c, 32'h3ee4a539} /* (6, 31, 9) {real, imag} */,
  {32'hbf2f5090, 32'hbe2bc1d1} /* (6, 31, 8) {real, imag} */,
  {32'hbf093dee, 32'h3d326728} /* (6, 31, 7) {real, imag} */,
  {32'h3ec17d26, 32'hbddfc2fa} /* (6, 31, 6) {real, imag} */,
  {32'hc0374f0c, 32'h3ee28e0a} /* (6, 31, 5) {real, imag} */,
  {32'h3fbed70e, 32'hbfc619ab} /* (6, 31, 4) {real, imag} */,
  {32'h40049d73, 32'h3f05217f} /* (6, 31, 3) {real, imag} */,
  {32'hc0b93089, 32'h3c345180} /* (6, 31, 2) {real, imag} */,
  {32'h41de82cb, 32'h40f286c0} /* (6, 31, 1) {real, imag} */,
  {32'h421fd30a, 32'hc0eb3175} /* (6, 31, 0) {real, imag} */,
  {32'hc11ecffa, 32'hc027fa80} /* (6, 30, 31) {real, imag} */,
  {32'h40d87e37, 32'h3d4528c0} /* (6, 30, 30) {real, imag} */,
  {32'hbee67c55, 32'hbfa03d1e} /* (6, 30, 29) {real, imag} */,
  {32'hc02e24a7, 32'h3da2a7b0} /* (6, 30, 28) {real, imag} */,
  {32'h3fb40b32, 32'hbe96e888} /* (6, 30, 27) {real, imag} */,
  {32'h3e28c640, 32'hbf094c50} /* (6, 30, 26) {real, imag} */,
  {32'hbe16b2b2, 32'h3f031a6c} /* (6, 30, 25) {real, imag} */,
  {32'h3f586070, 32'hbe1d26fc} /* (6, 30, 24) {real, imag} */,
  {32'h3ec30072, 32'hbef2c842} /* (6, 30, 23) {real, imag} */,
  {32'h3e47f755, 32'h3d57fb10} /* (6, 30, 22) {real, imag} */,
  {32'h3eae24dc, 32'hbf3dc8dc} /* (6, 30, 21) {real, imag} */,
  {32'hbebc19f0, 32'h3db15e10} /* (6, 30, 20) {real, imag} */,
  {32'h3d981f1e, 32'h3cffed15} /* (6, 30, 19) {real, imag} */,
  {32'h3e38db14, 32'hbdb5f704} /* (6, 30, 18) {real, imag} */,
  {32'h3dbf3712, 32'h3e86dd8c} /* (6, 30, 17) {real, imag} */,
  {32'hbb96e840, 32'h3ce291a8} /* (6, 30, 16) {real, imag} */,
  {32'hbdd0d590, 32'hbdd68cb6} /* (6, 30, 15) {real, imag} */,
  {32'hbeb67104, 32'h3ec8d701} /* (6, 30, 14) {real, imag} */,
  {32'h3e7990fa, 32'hbe9849d3} /* (6, 30, 13) {real, imag} */,
  {32'h3d44a074, 32'hbeca98a3} /* (6, 30, 12) {real, imag} */,
  {32'h3dc58a1d, 32'h3f03d576} /* (6, 30, 11) {real, imag} */,
  {32'h3c32a800, 32'h3d928536} /* (6, 30, 10) {real, imag} */,
  {32'hbef8c1be, 32'hbcf957e0} /* (6, 30, 9) {real, imag} */,
  {32'h3fad6493, 32'hbea87c6b} /* (6, 30, 8) {real, imag} */,
  {32'hbdcaef3c, 32'h3e96ee08} /* (6, 30, 7) {real, imag} */,
  {32'h3e81b47c, 32'hbd055b60} /* (6, 30, 6) {real, imag} */,
  {32'h3f308e0d, 32'h3f7c1d8b} /* (6, 30, 5) {real, imag} */,
  {32'h3e894bd4, 32'hbf76120d} /* (6, 30, 4) {real, imag} */,
  {32'hbfc88758, 32'hbf9287ec} /* (6, 30, 3) {real, imag} */,
  {32'h41307012, 32'h402c400d} /* (6, 30, 2) {real, imag} */,
  {32'hc19ffd87, 32'h3d449930} /* (6, 30, 1) {real, imag} */,
  {32'hc12ed24a, 32'h40925213} /* (6, 30, 0) {real, imag} */,
  {32'h40345df8, 32'hc06d5064} /* (6, 29, 31) {real, imag} */,
  {32'h3e3c4c3c, 32'h3eb546da} /* (6, 29, 30) {real, imag} */,
  {32'hbf4c68e0, 32'h3ebcb546} /* (6, 29, 29) {real, imag} */,
  {32'hbf51e1ba, 32'hbe8b9f11} /* (6, 29, 28) {real, imag} */,
  {32'h3f75f994, 32'h3f549451} /* (6, 29, 27) {real, imag} */,
  {32'h3dafb600, 32'h3f8e3130} /* (6, 29, 26) {real, imag} */,
  {32'hbea18e82, 32'hbd9f6da6} /* (6, 29, 25) {real, imag} */,
  {32'hbefbed88, 32'h3f199556} /* (6, 29, 24) {real, imag} */,
  {32'h3f148835, 32'hbd2958d0} /* (6, 29, 23) {real, imag} */,
  {32'hbf150e76, 32'hbe4fa509} /* (6, 29, 22) {real, imag} */,
  {32'h3efea02c, 32'hbccfda6c} /* (6, 29, 21) {real, imag} */,
  {32'hbdb9026c, 32'h3eea9420} /* (6, 29, 20) {real, imag} */,
  {32'h3d86d394, 32'h3ea7f34b} /* (6, 29, 19) {real, imag} */,
  {32'h3f4bcf8a, 32'hbe3ae89a} /* (6, 29, 18) {real, imag} */,
  {32'hbed1dd8e, 32'hbe8c2277} /* (6, 29, 17) {real, imag} */,
  {32'hbccab9f4, 32'hbd64e2ca} /* (6, 29, 16) {real, imag} */,
  {32'h3eb11e3c, 32'hbe484078} /* (6, 29, 15) {real, imag} */,
  {32'hbd26261c, 32'h3e1f8920} /* (6, 29, 14) {real, imag} */,
  {32'h3f23faa6, 32'hbeb90170} /* (6, 29, 13) {real, imag} */,
  {32'hbdb5145c, 32'hbea5aad0} /* (6, 29, 12) {real, imag} */,
  {32'hbe9cd648, 32'hbef3e68d} /* (6, 29, 11) {real, imag} */,
  {32'h3c507750, 32'h3e1d62cf} /* (6, 29, 10) {real, imag} */,
  {32'h3e8eb618, 32'h3da4a6cc} /* (6, 29, 9) {real, imag} */,
  {32'h3e8637ef, 32'h3f32ed8c} /* (6, 29, 8) {real, imag} */,
  {32'hbcebe0a0, 32'h3e95739a} /* (6, 29, 7) {real, imag} */,
  {32'hbf912008, 32'hbe665e23} /* (6, 29, 6) {real, imag} */,
  {32'h3e1591c0, 32'h3e3fc9e7} /* (6, 29, 5) {real, imag} */,
  {32'h3f4e4a34, 32'hbf54a4a1} /* (6, 29, 4) {real, imag} */,
  {32'h3e575f26, 32'h3c230910} /* (6, 29, 3) {real, imag} */,
  {32'h3f1eac7a, 32'h407caf3a} /* (6, 29, 2) {real, imag} */,
  {32'hc03b06ef, 32'hbf75c638} /* (6, 29, 1) {real, imag} */,
  {32'h3f45c137, 32'hc001562d} /* (6, 29, 0) {real, imag} */,
  {32'h3fe94d46, 32'hc0122f85} /* (6, 28, 31) {real, imag} */,
  {32'hbfdb88d7, 32'h3fc63d81} /* (6, 28, 30) {real, imag} */,
  {32'hbe8cc302, 32'hbe2bf7cc} /* (6, 28, 29) {real, imag} */,
  {32'h3e8935ba, 32'hbf1139ee} /* (6, 28, 28) {real, imag} */,
  {32'hbf0b23d4, 32'h3edf882c} /* (6, 28, 27) {real, imag} */,
  {32'hbefad5f8, 32'hbf705d98} /* (6, 28, 26) {real, imag} */,
  {32'h3dbeec46, 32'hbd832086} /* (6, 28, 25) {real, imag} */,
  {32'hbf3a7c42, 32'hbeb384fd} /* (6, 28, 24) {real, imag} */,
  {32'h3ef00d3c, 32'h3ed13acf} /* (6, 28, 23) {real, imag} */,
  {32'hbea01d00, 32'hbd84a154} /* (6, 28, 22) {real, imag} */,
  {32'h3d3fa660, 32'h3df82686} /* (6, 28, 21) {real, imag} */,
  {32'hbc915ad0, 32'hbf427f36} /* (6, 28, 20) {real, imag} */,
  {32'h3ed482d6, 32'h3f145c59} /* (6, 28, 19) {real, imag} */,
  {32'h3ce36570, 32'h3ed94274} /* (6, 28, 18) {real, imag} */,
  {32'hbe40b34d, 32'hbe99a613} /* (6, 28, 17) {real, imag} */,
  {32'hbdbba422, 32'hbe478412} /* (6, 28, 16) {real, imag} */,
  {32'h3e6d938a, 32'h3ddd3a06} /* (6, 28, 15) {real, imag} */,
  {32'h3edc3030, 32'h3ec33461} /* (6, 28, 14) {real, imag} */,
  {32'hbd7049ac, 32'h3def67c2} /* (6, 28, 13) {real, imag} */,
  {32'h3ef6841e, 32'h3c71e348} /* (6, 28, 12) {real, imag} */,
  {32'h3ea4f472, 32'hbd7dfa78} /* (6, 28, 11) {real, imag} */,
  {32'hbf1a3ab7, 32'h3d414a5a} /* (6, 28, 10) {real, imag} */,
  {32'hbe796c39, 32'h3e09e54c} /* (6, 28, 9) {real, imag} */,
  {32'hbf2270ce, 32'h3e69add8} /* (6, 28, 8) {real, imag} */,
  {32'hbdb25355, 32'hbe84d2ef} /* (6, 28, 7) {real, imag} */,
  {32'h3d8a21b4, 32'h3f1ae96e} /* (6, 28, 6) {real, imag} */,
  {32'h3d700f0a, 32'hbec44c9e} /* (6, 28, 5) {real, imag} */,
  {32'h3eb9a3ff, 32'h3ed341c9} /* (6, 28, 4) {real, imag} */,
  {32'h3e8e828e, 32'hbec496fe} /* (6, 28, 3) {real, imag} */,
  {32'hbfb6af96, 32'h3fd036cd} /* (6, 28, 2) {real, imag} */,
  {32'h3e971e0e, 32'hbfde02ae} /* (6, 28, 1) {real, imag} */,
  {32'h3fbff7ff, 32'h3e6215a8} /* (6, 28, 0) {real, imag} */,
  {32'hbf08b77c, 32'h3fd01214} /* (6, 27, 31) {real, imag} */,
  {32'h3f6b0e63, 32'hbf9b3060} /* (6, 27, 30) {real, imag} */,
  {32'hbb4ec240, 32'hbecff8c1} /* (6, 27, 29) {real, imag} */,
  {32'hbe37f7a2, 32'h3eabd8e5} /* (6, 27, 28) {real, imag} */,
  {32'h3d833d94, 32'hbe727dc0} /* (6, 27, 27) {real, imag} */,
  {32'h3ec310f8, 32'hbe8564d2} /* (6, 27, 26) {real, imag} */,
  {32'hbe8bff0d, 32'h3df9e8f8} /* (6, 27, 25) {real, imag} */,
  {32'h3dd63eac, 32'h3ecbdfd9} /* (6, 27, 24) {real, imag} */,
  {32'hbe98c2e6, 32'h3e891009} /* (6, 27, 23) {real, imag} */,
  {32'hbe242274, 32'hbe9dfa80} /* (6, 27, 22) {real, imag} */,
  {32'h3eb0dca6, 32'hbeb7c138} /* (6, 27, 21) {real, imag} */,
  {32'hbe6fae90, 32'h3f3e7872} /* (6, 27, 20) {real, imag} */,
  {32'h3e57544c, 32'hbeab5fde} /* (6, 27, 19) {real, imag} */,
  {32'h3d16ab78, 32'hbd8f2bf4} /* (6, 27, 18) {real, imag} */,
  {32'h3d49d02c, 32'h3a0529c0} /* (6, 27, 17) {real, imag} */,
  {32'h3b26b440, 32'h3e5d36f9} /* (6, 27, 16) {real, imag} */,
  {32'hbe7662e1, 32'hbd0164ac} /* (6, 27, 15) {real, imag} */,
  {32'hbb075d60, 32'h3d7046f4} /* (6, 27, 14) {real, imag} */,
  {32'hbde26f96, 32'h3eb253e6} /* (6, 27, 13) {real, imag} */,
  {32'h3ea41177, 32'h3ed80c18} /* (6, 27, 12) {real, imag} */,
  {32'h3e6ea60b, 32'h3f5a0ec7} /* (6, 27, 11) {real, imag} */,
  {32'hbef62ffc, 32'hbf3ef540} /* (6, 27, 10) {real, imag} */,
  {32'h3d8ebfca, 32'h3e0d85e3} /* (6, 27, 9) {real, imag} */,
  {32'hbe704bf9, 32'hbe7a7c4f} /* (6, 27, 8) {real, imag} */,
  {32'hbe1b52d6, 32'hbe4b9210} /* (6, 27, 7) {real, imag} */,
  {32'h3e23f8b1, 32'h3d7b6f42} /* (6, 27, 6) {real, imag} */,
  {32'h3f840590, 32'hbed45966} /* (6, 27, 5) {real, imag} */,
  {32'hbf9219f4, 32'h3e2db710} /* (6, 27, 4) {real, imag} */,
  {32'hbf1598a2, 32'hbde25794} /* (6, 27, 3) {real, imag} */,
  {32'h3fc61b96, 32'hbf259a98} /* (6, 27, 2) {real, imag} */,
  {32'hbfe929f8, 32'hbfb528e2} /* (6, 27, 1) {real, imag} */,
  {32'hbfdde6d8, 32'h3f602773} /* (6, 27, 0) {real, imag} */,
  {32'hbf725449, 32'hbf3a5230} /* (6, 26, 31) {real, imag} */,
  {32'hbfb23dbd, 32'hbeb87a7e} /* (6, 26, 30) {real, imag} */,
  {32'hbf3a26b1, 32'h3f1fc4f8} /* (6, 26, 29) {real, imag} */,
  {32'h3e9b2dc6, 32'hbe1521bc} /* (6, 26, 28) {real, imag} */,
  {32'hbe752a8c, 32'hbed241eb} /* (6, 26, 27) {real, imag} */,
  {32'hba791200, 32'hbea9fe2c} /* (6, 26, 26) {real, imag} */,
  {32'h3f4354a0, 32'h3ec22846} /* (6, 26, 25) {real, imag} */,
  {32'h3cc6d490, 32'hbe815a9a} /* (6, 26, 24) {real, imag} */,
  {32'h3dccd7a8, 32'hbf42697a} /* (6, 26, 23) {real, imag} */,
  {32'h3e47178b, 32'hbe5809a2} /* (6, 26, 22) {real, imag} */,
  {32'h3ed5870c, 32'h3ca19fd0} /* (6, 26, 21) {real, imag} */,
  {32'hbe09dd10, 32'h3e049a1f} /* (6, 26, 20) {real, imag} */,
  {32'hbdf8291c, 32'h3e6cdc0a} /* (6, 26, 19) {real, imag} */,
  {32'hbd27852a, 32'h3df1f654} /* (6, 26, 18) {real, imag} */,
  {32'h3a236900, 32'hbe89df2c} /* (6, 26, 17) {real, imag} */,
  {32'hbd32243c, 32'hbd8431d0} /* (6, 26, 16) {real, imag} */,
  {32'hbf22b1f6, 32'h3ef07c04} /* (6, 26, 15) {real, imag} */,
  {32'h3e0ed292, 32'hbea61958} /* (6, 26, 14) {real, imag} */,
  {32'hbe85bcb2, 32'h3f2c5708} /* (6, 26, 13) {real, imag} */,
  {32'h3d0cbbc6, 32'hbda87c12} /* (6, 26, 12) {real, imag} */,
  {32'hbede5b16, 32'h3e88b3ef} /* (6, 26, 11) {real, imag} */,
  {32'h3e13aefc, 32'hbdcc3652} /* (6, 26, 10) {real, imag} */,
  {32'hbd8b0936, 32'h3f0a3c23} /* (6, 26, 9) {real, imag} */,
  {32'hbd021c32, 32'h3d200d60} /* (6, 26, 8) {real, imag} */,
  {32'h3e8cc555, 32'hbf058720} /* (6, 26, 7) {real, imag} */,
  {32'h3f053e5a, 32'h3ea2980e} /* (6, 26, 6) {real, imag} */,
  {32'hbd36bffc, 32'hbe77c3e6} /* (6, 26, 5) {real, imag} */,
  {32'h3e747737, 32'h3e7202ba} /* (6, 26, 4) {real, imag} */,
  {32'hbe98f380, 32'hbddae2c4} /* (6, 26, 3) {real, imag} */,
  {32'hbeda9cf6, 32'h3f1195f0} /* (6, 26, 2) {real, imag} */,
  {32'h3ec7d0d2, 32'hbf3dc1ec} /* (6, 26, 1) {real, imag} */,
  {32'h3cf6d520, 32'h3f391890} /* (6, 26, 0) {real, imag} */,
  {32'hbe25e802, 32'hbf2a930f} /* (6, 25, 31) {real, imag} */,
  {32'h3e2e506c, 32'h3f25af8c} /* (6, 25, 30) {real, imag} */,
  {32'h3d3921c8, 32'hbea8c78a} /* (6, 25, 29) {real, imag} */,
  {32'h3f196716, 32'hbedf5b22} /* (6, 25, 28) {real, imag} */,
  {32'h3ed30722, 32'h3df5e6c2} /* (6, 25, 27) {real, imag} */,
  {32'h3f43ecb4, 32'hbe32e572} /* (6, 25, 26) {real, imag} */,
  {32'hbd2c60c8, 32'hbe331cb9} /* (6, 25, 25) {real, imag} */,
  {32'hbdfde2d2, 32'hbe70d761} /* (6, 25, 24) {real, imag} */,
  {32'h3f180028, 32'hbd6a490c} /* (6, 25, 23) {real, imag} */,
  {32'h3ce27ac0, 32'h3e1385b9} /* (6, 25, 22) {real, imag} */,
  {32'hbe16216c, 32'h3de5748e} /* (6, 25, 21) {real, imag} */,
  {32'hbcc11de0, 32'h3e07f729} /* (6, 25, 20) {real, imag} */,
  {32'h3e8b6d3c, 32'hbd8215d1} /* (6, 25, 19) {real, imag} */,
  {32'h3e848564, 32'h3d562005} /* (6, 25, 18) {real, imag} */,
  {32'hbeccd932, 32'hbe5119ce} /* (6, 25, 17) {real, imag} */,
  {32'hbef72f22, 32'h3d8f89d1} /* (6, 25, 16) {real, imag} */,
  {32'hbc94f88a, 32'h3e5173dc} /* (6, 25, 15) {real, imag} */,
  {32'h3d834462, 32'h3f0c8496} /* (6, 25, 14) {real, imag} */,
  {32'hbee8c74a, 32'hbebda0e6} /* (6, 25, 13) {real, imag} */,
  {32'hbe03e732, 32'h3ea979fe} /* (6, 25, 12) {real, imag} */,
  {32'h3e7eebc2, 32'hbd692808} /* (6, 25, 11) {real, imag} */,
  {32'hbe6106c7, 32'hbf4cfa39} /* (6, 25, 10) {real, imag} */,
  {32'hbedc88d2, 32'hbde44d00} /* (6, 25, 9) {real, imag} */,
  {32'h3e2a2e4a, 32'h3d4c0168} /* (6, 25, 8) {real, imag} */,
  {32'h3ea9dc72, 32'h3f2e2f00} /* (6, 25, 7) {real, imag} */,
  {32'hbf223f48, 32'h3c7113c0} /* (6, 25, 6) {real, imag} */,
  {32'hbd83be64, 32'hbf12afb1} /* (6, 25, 5) {real, imag} */,
  {32'hbf56b4e8, 32'h3e01b000} /* (6, 25, 4) {real, imag} */,
  {32'hbef274f6, 32'hbee590e5} /* (6, 25, 3) {real, imag} */,
  {32'hbd9232a4, 32'hbefade4b} /* (6, 25, 2) {real, imag} */,
  {32'h3f08278e, 32'hbf1b5262} /* (6, 25, 1) {real, imag} */,
  {32'h3e7f5802, 32'h3df08bed} /* (6, 25, 0) {real, imag} */,
  {32'hbf694d0c, 32'h3f480658} /* (6, 24, 31) {real, imag} */,
  {32'h3f6dbb79, 32'hbea4b57d} /* (6, 24, 30) {real, imag} */,
  {32'h3d528dc0, 32'hbe577852} /* (6, 24, 29) {real, imag} */,
  {32'hbed68347, 32'h3efc68f3} /* (6, 24, 28) {real, imag} */,
  {32'hbf070efe, 32'hbe43ea96} /* (6, 24, 27) {real, imag} */,
  {32'hbf42933c, 32'hbdb61ffd} /* (6, 24, 26) {real, imag} */,
  {32'h3e1c97c8, 32'hbdc3b98c} /* (6, 24, 25) {real, imag} */,
  {32'hbd8591a4, 32'hbf0a90ec} /* (6, 24, 24) {real, imag} */,
  {32'hbf028819, 32'hbf08bd20} /* (6, 24, 23) {real, imag} */,
  {32'hbe2ef400, 32'h3b1cf000} /* (6, 24, 22) {real, imag} */,
  {32'h3e9a4d44, 32'hbe70dc23} /* (6, 24, 21) {real, imag} */,
  {32'h3cb8a91e, 32'hbebeaca8} /* (6, 24, 20) {real, imag} */,
  {32'h3e29b190, 32'h3d37515a} /* (6, 24, 19) {real, imag} */,
  {32'h3e15d88f, 32'h3eb24ddb} /* (6, 24, 18) {real, imag} */,
  {32'h3ea793e2, 32'hbe9f2b87} /* (6, 24, 17) {real, imag} */,
  {32'h3e6cc261, 32'hbe8837df} /* (6, 24, 16) {real, imag} */,
  {32'hbe7f0707, 32'hbc1366a0} /* (6, 24, 15) {real, imag} */,
  {32'hbd8644c8, 32'h3db0405b} /* (6, 24, 14) {real, imag} */,
  {32'h3e23beff, 32'hbdf827ee} /* (6, 24, 13) {real, imag} */,
  {32'hbe84844e, 32'h3dc8abd2} /* (6, 24, 12) {real, imag} */,
  {32'h3ed2de4a, 32'hbe376523} /* (6, 24, 11) {real, imag} */,
  {32'hbdfd1440, 32'hbe5a7b1a} /* (6, 24, 10) {real, imag} */,
  {32'h3e937530, 32'hbd8adae6} /* (6, 24, 9) {real, imag} */,
  {32'h3eb2582e, 32'h3e9dcacc} /* (6, 24, 8) {real, imag} */,
  {32'hbbcbe340, 32'h3eb63465} /* (6, 24, 7) {real, imag} */,
  {32'h3d57a6c8, 32'h3e0c094a} /* (6, 24, 6) {real, imag} */,
  {32'h3f39e2a0, 32'h3eeb7a88} /* (6, 24, 5) {real, imag} */,
  {32'hbf2c51df, 32'hbf11b442} /* (6, 24, 4) {real, imag} */,
  {32'h3ed0e104, 32'hbf2c9af2} /* (6, 24, 3) {real, imag} */,
  {32'h3f19af10, 32'hbdf0a2e7} /* (6, 24, 2) {real, imag} */,
  {32'hbf70afaa, 32'h3f22f0a1} /* (6, 24, 1) {real, imag} */,
  {32'hbf72cf56, 32'h3f87d76e} /* (6, 24, 0) {real, imag} */,
  {32'h3cce5bf4, 32'hbe1c9553} /* (6, 23, 31) {real, imag} */,
  {32'hbdf7f940, 32'h3f1459c4} /* (6, 23, 30) {real, imag} */,
  {32'h3f5c493b, 32'hbe88a96e} /* (6, 23, 29) {real, imag} */,
  {32'hbe1a39c2, 32'h3f081570} /* (6, 23, 28) {real, imag} */,
  {32'h3ec08947, 32'h3cf5cf70} /* (6, 23, 27) {real, imag} */,
  {32'h3e8a79d8, 32'hbe50e5e9} /* (6, 23, 26) {real, imag} */,
  {32'h3f00addf, 32'h3d3a01c8} /* (6, 23, 25) {real, imag} */,
  {32'h3e54b958, 32'hbd1a0578} /* (6, 23, 24) {real, imag} */,
  {32'h3e8a5192, 32'hbf109d0d} /* (6, 23, 23) {real, imag} */,
  {32'hbda39f27, 32'h3fb35d9a} /* (6, 23, 22) {real, imag} */,
  {32'hbe352fd7, 32'h3d431454} /* (6, 23, 21) {real, imag} */,
  {32'hbccb9760, 32'hbe8be03e} /* (6, 23, 20) {real, imag} */,
  {32'hbc6e6230, 32'hbe62c92f} /* (6, 23, 19) {real, imag} */,
  {32'hbd2013cc, 32'hbd153b81} /* (6, 23, 18) {real, imag} */,
  {32'hbee71edd, 32'hbe5a9202} /* (6, 23, 17) {real, imag} */,
  {32'hbd61fe60, 32'hbded0371} /* (6, 23, 16) {real, imag} */,
  {32'hbe27da75, 32'hbf00523f} /* (6, 23, 15) {real, imag} */,
  {32'h3e8fcd0c, 32'h3cf701e0} /* (6, 23, 14) {real, imag} */,
  {32'hbf6ed2e7, 32'hbf052710} /* (6, 23, 13) {real, imag} */,
  {32'h3ee6138f, 32'hbf4ecede} /* (6, 23, 12) {real, imag} */,
  {32'h3de46ef2, 32'h3ecb4c3a} /* (6, 23, 11) {real, imag} */,
  {32'hbe11229d, 32'h3e9b054f} /* (6, 23, 10) {real, imag} */,
  {32'h3d6528c9, 32'hbdc538a4} /* (6, 23, 9) {real, imag} */,
  {32'hbe05a6f4, 32'hbeee75a0} /* (6, 23, 8) {real, imag} */,
  {32'hbcc02e40, 32'hbe956fd3} /* (6, 23, 7) {real, imag} */,
  {32'hbddb1b77, 32'h3efa202d} /* (6, 23, 6) {real, imag} */,
  {32'hbd4946c6, 32'hbe78137a} /* (6, 23, 5) {real, imag} */,
  {32'hbdd3a2d6, 32'hbf0db652} /* (6, 23, 4) {real, imag} */,
  {32'hbec487f8, 32'h3ee68f96} /* (6, 23, 3) {real, imag} */,
  {32'h3be3eb40, 32'hbe5eb6b6} /* (6, 23, 2) {real, imag} */,
  {32'hbda91446, 32'hbf560dc0} /* (6, 23, 1) {real, imag} */,
  {32'hbec10ec0, 32'hbf12713c} /* (6, 23, 0) {real, imag} */,
  {32'h3f0ff111, 32'h3e51efee} /* (6, 22, 31) {real, imag} */,
  {32'hbed515e8, 32'h3f4d9bfa} /* (6, 22, 30) {real, imag} */,
  {32'hbf00027c, 32'hbdb07a14} /* (6, 22, 29) {real, imag} */,
  {32'hbd156669, 32'hbe0e48ca} /* (6, 22, 28) {real, imag} */,
  {32'h3e4ab31c, 32'h3e95d26b} /* (6, 22, 27) {real, imag} */,
  {32'h3c85f5f0, 32'hbebe755f} /* (6, 22, 26) {real, imag} */,
  {32'h3ed8df24, 32'hbe30fc8a} /* (6, 22, 25) {real, imag} */,
  {32'h3eb1462a, 32'h3ef306be} /* (6, 22, 24) {real, imag} */,
  {32'hbefc7dad, 32'h3f2cf84a} /* (6, 22, 23) {real, imag} */,
  {32'hbf2d4f58, 32'hbf463174} /* (6, 22, 22) {real, imag} */,
  {32'h3ef500b2, 32'h3eb33171} /* (6, 22, 21) {real, imag} */,
  {32'hbe1ec6ba, 32'hbe61c4a4} /* (6, 22, 20) {real, imag} */,
  {32'hbf0d9cce, 32'hbe8925aa} /* (6, 22, 19) {real, imag} */,
  {32'h3ea6951e, 32'hbf2780e8} /* (6, 22, 18) {real, imag} */,
  {32'hbd7339b6, 32'hbe549d4b} /* (6, 22, 17) {real, imag} */,
  {32'hbe444769, 32'h3e700cda} /* (6, 22, 16) {real, imag} */,
  {32'h3e91f71c, 32'hba557e40} /* (6, 22, 15) {real, imag} */,
  {32'hbe7dd2f2, 32'hbcbbf0f0} /* (6, 22, 14) {real, imag} */,
  {32'hbe839fa8, 32'hbe224a5a} /* (6, 22, 13) {real, imag} */,
  {32'hbe02e346, 32'h3e2e9ec9} /* (6, 22, 12) {real, imag} */,
  {32'hbe424b6a, 32'h3ecadcae} /* (6, 22, 11) {real, imag} */,
  {32'h3d6eeaf8, 32'hbf3229a6} /* (6, 22, 10) {real, imag} */,
  {32'h3dc9d454, 32'h3d45b920} /* (6, 22, 9) {real, imag} */,
  {32'h3e4cce45, 32'h3ed72acc} /* (6, 22, 8) {real, imag} */,
  {32'h3d8ca2ac, 32'hbdd5916a} /* (6, 22, 7) {real, imag} */,
  {32'h3ee7e346, 32'h3ef31b00} /* (6, 22, 6) {real, imag} */,
  {32'h3d465e04, 32'hbd374894} /* (6, 22, 5) {real, imag} */,
  {32'h3ecbc55e, 32'hbc0f17b4} /* (6, 22, 4) {real, imag} */,
  {32'hbe2f7e17, 32'h3f269520} /* (6, 22, 3) {real, imag} */,
  {32'hbe645c46, 32'h3f7184d0} /* (6, 22, 2) {real, imag} */,
  {32'hbf1044d4, 32'hbe65fece} /* (6, 22, 1) {real, imag} */,
  {32'hbea071da, 32'hbf86e6e9} /* (6, 22, 0) {real, imag} */,
  {32'hbd37f768, 32'h3f6db7e6} /* (6, 21, 31) {real, imag} */,
  {32'hbdd9996d, 32'hbf5beb42} /* (6, 21, 30) {real, imag} */,
  {32'hbe7f92cc, 32'hbeb646dc} /* (6, 21, 29) {real, imag} */,
  {32'hbe9fdb73, 32'hbf1a6a70} /* (6, 21, 28) {real, imag} */,
  {32'h3e52859e, 32'h3c947108} /* (6, 21, 27) {real, imag} */,
  {32'hbe11a11d, 32'h3e8557e7} /* (6, 21, 26) {real, imag} */,
  {32'hbec8d70a, 32'h3e9404d3} /* (6, 21, 25) {real, imag} */,
  {32'hbe35955e, 32'hbede14a7} /* (6, 21, 24) {real, imag} */,
  {32'hbd17ae9e, 32'h3f17bedd} /* (6, 21, 23) {real, imag} */,
  {32'hbe1024b4, 32'h3f03142c} /* (6, 21, 22) {real, imag} */,
  {32'hbe9b0f5c, 32'hbc576300} /* (6, 21, 21) {real, imag} */,
  {32'h3f082813, 32'hbda67abe} /* (6, 21, 20) {real, imag} */,
  {32'h3e4fae3a, 32'hbed2e5a7} /* (6, 21, 19) {real, imag} */,
  {32'hbe22462e, 32'hbdb9feb3} /* (6, 21, 18) {real, imag} */,
  {32'hba19d200, 32'hbed45cfa} /* (6, 21, 17) {real, imag} */,
  {32'hbda44595, 32'hbd0ce07c} /* (6, 21, 16) {real, imag} */,
  {32'hbe4458a1, 32'h3cb9c6b0} /* (6, 21, 15) {real, imag} */,
  {32'hbe07e2a4, 32'h3d99176c} /* (6, 21, 14) {real, imag} */,
  {32'h3ea33bdf, 32'h3f2d7946} /* (6, 21, 13) {real, imag} */,
  {32'hbe3e7283, 32'hbdc5ff8a} /* (6, 21, 12) {real, imag} */,
  {32'hbe8fefee, 32'hbf2fe4c0} /* (6, 21, 11) {real, imag} */,
  {32'hbe738ee1, 32'hbecb77a8} /* (6, 21, 10) {real, imag} */,
  {32'h3ec0c697, 32'hbe50aa52} /* (6, 21, 9) {real, imag} */,
  {32'h3ec8ac3c, 32'hbe0fe6e7} /* (6, 21, 8) {real, imag} */,
  {32'h3e9fa7ec, 32'h3eab5800} /* (6, 21, 7) {real, imag} */,
  {32'h3e9140fd, 32'h3e948570} /* (6, 21, 6) {real, imag} */,
  {32'hbdeda93c, 32'hbdb3c00e} /* (6, 21, 5) {real, imag} */,
  {32'hbdb2f47c, 32'h3e2e7080} /* (6, 21, 4) {real, imag} */,
  {32'hbdb6736e, 32'hbdc8e4e8} /* (6, 21, 3) {real, imag} */,
  {32'h3e24a528, 32'hbe6b88ba} /* (6, 21, 2) {real, imag} */,
  {32'hbeb4a1f9, 32'h3f1a9502} /* (6, 21, 1) {real, imag} */,
  {32'h3ec7da22, 32'h3ea1e9e4} /* (6, 21, 0) {real, imag} */,
  {32'hbe4ed62d, 32'h3edaa48c} /* (6, 20, 31) {real, imag} */,
  {32'hbd0fc158, 32'hbe1d2c56} /* (6, 20, 30) {real, imag} */,
  {32'hbf03f567, 32'hbda882c2} /* (6, 20, 29) {real, imag} */,
  {32'h3e7f155f, 32'hbdb1dc27} /* (6, 20, 28) {real, imag} */,
  {32'h3c8d16a8, 32'hbe230e64} /* (6, 20, 27) {real, imag} */,
  {32'hbe2be016, 32'hbe6c3316} /* (6, 20, 26) {real, imag} */,
  {32'h3eca39c4, 32'h3d988ce8} /* (6, 20, 25) {real, imag} */,
  {32'h3e567a64, 32'hbeed9831} /* (6, 20, 24) {real, imag} */,
  {32'h3e8747b1, 32'hbea769fc} /* (6, 20, 23) {real, imag} */,
  {32'hbefec0df, 32'hbd0e52d4} /* (6, 20, 22) {real, imag} */,
  {32'hbe5cd7bf, 32'hbca734b8} /* (6, 20, 21) {real, imag} */,
  {32'h3d955a42, 32'h3ef43535} /* (6, 20, 20) {real, imag} */,
  {32'h3e5a52e5, 32'h3ecb18c0} /* (6, 20, 19) {real, imag} */,
  {32'hbeb97bd8, 32'hbd12bcd6} /* (6, 20, 18) {real, imag} */,
  {32'h3e0d8432, 32'hbf0a4295} /* (6, 20, 17) {real, imag} */,
  {32'hbd0ddca4, 32'hbe57546a} /* (6, 20, 16) {real, imag} */,
  {32'h3e99cc85, 32'h3e73e896} /* (6, 20, 15) {real, imag} */,
  {32'h3e194d21, 32'h3d75cf3a} /* (6, 20, 14) {real, imag} */,
  {32'h3e41eb62, 32'hbed16cb2} /* (6, 20, 13) {real, imag} */,
  {32'hbd65cd34, 32'h3ee53052} /* (6, 20, 12) {real, imag} */,
  {32'h3eb44244, 32'hbe211ca6} /* (6, 20, 11) {real, imag} */,
  {32'h3e294351, 32'hbe0f4ea8} /* (6, 20, 10) {real, imag} */,
  {32'h3e3121b8, 32'h3e5c1c5f} /* (6, 20, 9) {real, imag} */,
  {32'hbe784860, 32'h3e10cdfb} /* (6, 20, 8) {real, imag} */,
  {32'hbedf9120, 32'hbe969f67} /* (6, 20, 7) {real, imag} */,
  {32'h3e4481cd, 32'hbe8256d8} /* (6, 20, 6) {real, imag} */,
  {32'h3eabe18c, 32'hbd2fa3a8} /* (6, 20, 5) {real, imag} */,
  {32'h3e3ae797, 32'h3eab363d} /* (6, 20, 4) {real, imag} */,
  {32'hbb5b9980, 32'h3d2447c0} /* (6, 20, 3) {real, imag} */,
  {32'hbdd5bb68, 32'h3e15d054} /* (6, 20, 2) {real, imag} */,
  {32'h3e965b8e, 32'h3e92a665} /* (6, 20, 1) {real, imag} */,
  {32'hbe382c6d, 32'hbeaff3fb} /* (6, 20, 0) {real, imag} */,
  {32'h3e8dbce0, 32'hbee36ef1} /* (6, 19, 31) {real, imag} */,
  {32'h3e6e07ef, 32'h3edb1e67} /* (6, 19, 30) {real, imag} */,
  {32'hbc57e720, 32'h3d0de098} /* (6, 19, 29) {real, imag} */,
  {32'hbc1da860, 32'hbe462b30} /* (6, 19, 28) {real, imag} */,
  {32'h3e6b2508, 32'h3bce38c0} /* (6, 19, 27) {real, imag} */,
  {32'h3f05fd17, 32'h3e165e2c} /* (6, 19, 26) {real, imag} */,
  {32'hbea5e8ff, 32'hbe873b4c} /* (6, 19, 25) {real, imag} */,
  {32'h3e753082, 32'hbeef2f3c} /* (6, 19, 24) {real, imag} */,
  {32'hbf091b2a, 32'h3d9233cc} /* (6, 19, 23) {real, imag} */,
  {32'hbe0332c3, 32'h3e32fdd0} /* (6, 19, 22) {real, imag} */,
  {32'hbd831afc, 32'hbe9b34a4} /* (6, 19, 21) {real, imag} */,
  {32'h3e4fd7c7, 32'h3dbf0d94} /* (6, 19, 20) {real, imag} */,
  {32'hbed5dff2, 32'hbea54b22} /* (6, 19, 19) {real, imag} */,
  {32'h3dbf30cc, 32'hbd8aa9ac} /* (6, 19, 18) {real, imag} */,
  {32'hbdb2cf15, 32'h3edacb83} /* (6, 19, 17) {real, imag} */,
  {32'h3d423c69, 32'hbe0b07aa} /* (6, 19, 16) {real, imag} */,
  {32'h3dca2956, 32'hbb74d020} /* (6, 19, 15) {real, imag} */,
  {32'hbe10d9d0, 32'hbe359d22} /* (6, 19, 14) {real, imag} */,
  {32'h3e5b5c0c, 32'h3ed388e0} /* (6, 19, 13) {real, imag} */,
  {32'hbee00398, 32'h3e1adec6} /* (6, 19, 12) {real, imag} */,
  {32'hbe145755, 32'hbe3824ad} /* (6, 19, 11) {real, imag} */,
  {32'h3eaf4f85, 32'h3e947e7c} /* (6, 19, 10) {real, imag} */,
  {32'h3dc007ec, 32'h3e83fdcd} /* (6, 19, 9) {real, imag} */,
  {32'h3d74bdd2, 32'hbe44d71c} /* (6, 19, 8) {real, imag} */,
  {32'h3eacc9fc, 32'hbd9f30b1} /* (6, 19, 7) {real, imag} */,
  {32'hbca71a80, 32'hbb647d20} /* (6, 19, 6) {real, imag} */,
  {32'hbee83e9e, 32'h3d60d5c8} /* (6, 19, 5) {real, imag} */,
  {32'hbd9f39d6, 32'h3e160674} /* (6, 19, 4) {real, imag} */,
  {32'h3e8a05fc, 32'hbe577f42} /* (6, 19, 3) {real, imag} */,
  {32'hbe55c405, 32'hbae76e00} /* (6, 19, 2) {real, imag} */,
  {32'hbd48976c, 32'h3f124165} /* (6, 19, 1) {real, imag} */,
  {32'h3e3a8ad4, 32'hbef70261} /* (6, 19, 0) {real, imag} */,
  {32'hbe82f185, 32'h3c40a250} /* (6, 18, 31) {real, imag} */,
  {32'h3ecac3cd, 32'hbe25643b} /* (6, 18, 30) {real, imag} */,
  {32'h3e8e9177, 32'hbd86d5e0} /* (6, 18, 29) {real, imag} */,
  {32'hbe9108cd, 32'h3d1482fe} /* (6, 18, 28) {real, imag} */,
  {32'hbd0f22ca, 32'hbed2e9de} /* (6, 18, 27) {real, imag} */,
  {32'hbdf251f1, 32'hbedc36ab} /* (6, 18, 26) {real, imag} */,
  {32'hbea2c903, 32'hbe86e040} /* (6, 18, 25) {real, imag} */,
  {32'hbe841503, 32'h3c278f8c} /* (6, 18, 24) {real, imag} */,
  {32'h3e1bb96e, 32'h3dc30c34} /* (6, 18, 23) {real, imag} */,
  {32'h3ef25a54, 32'hbe23eecb} /* (6, 18, 22) {real, imag} */,
  {32'hbf71a9d2, 32'hb9c59c00} /* (6, 18, 21) {real, imag} */,
  {32'hbd0fee60, 32'hbd2d7970} /* (6, 18, 20) {real, imag} */,
  {32'h3e54d026, 32'h3e21ca1a} /* (6, 18, 19) {real, imag} */,
  {32'h3df21caa, 32'hbe84c775} /* (6, 18, 18) {real, imag} */,
  {32'h3e924ea5, 32'hbe8982cb} /* (6, 18, 17) {real, imag} */,
  {32'hbe6ba45d, 32'hbde6018d} /* (6, 18, 16) {real, imag} */,
  {32'hbe875ab4, 32'hbe483d84} /* (6, 18, 15) {real, imag} */,
  {32'h3eaf5613, 32'h3e7a4688} /* (6, 18, 14) {real, imag} */,
  {32'hbe44d74e, 32'h3eb5534a} /* (6, 18, 13) {real, imag} */,
  {32'h3e25dc33, 32'hbf335d1c} /* (6, 18, 12) {real, imag} */,
  {32'h3e81cbd8, 32'h3c7f4a1c} /* (6, 18, 11) {real, imag} */,
  {32'hbf134589, 32'h3ee066d4} /* (6, 18, 10) {real, imag} */,
  {32'hbea37c36, 32'h3edae775} /* (6, 18, 9) {real, imag} */,
  {32'hbede746a, 32'h3f24235c} /* (6, 18, 8) {real, imag} */,
  {32'hbee78cb6, 32'h3d18e298} /* (6, 18, 7) {real, imag} */,
  {32'hbb319e80, 32'hbe13b5b0} /* (6, 18, 6) {real, imag} */,
  {32'h3d87038a, 32'hbe55fa26} /* (6, 18, 5) {real, imag} */,
  {32'h3d2e7a76, 32'hbe830567} /* (6, 18, 4) {real, imag} */,
  {32'h3e098c6c, 32'hbed3724e} /* (6, 18, 3) {real, imag} */,
  {32'hbe26fa77, 32'hbe8f1400} /* (6, 18, 2) {real, imag} */,
  {32'h3ec5b862, 32'h3f6842cb} /* (6, 18, 1) {real, imag} */,
  {32'hbd54305a, 32'h3e33f654} /* (6, 18, 0) {real, imag} */,
  {32'h3f1afcd5, 32'hbdd87615} /* (6, 17, 31) {real, imag} */,
  {32'hbbf3d8ac, 32'h3e83ae97} /* (6, 17, 30) {real, imag} */,
  {32'hbd028770, 32'hbe1f5162} /* (6, 17, 29) {real, imag} */,
  {32'hbdd3b349, 32'h3eb4afaa} /* (6, 17, 28) {real, imag} */,
  {32'hbe232944, 32'hbe76c924} /* (6, 17, 27) {real, imag} */,
  {32'h3d0e4ec7, 32'h3e1f85e6} /* (6, 17, 26) {real, imag} */,
  {32'h3d52125a, 32'hbe689ea9} /* (6, 17, 25) {real, imag} */,
  {32'h3df092c6, 32'hbd7b747f} /* (6, 17, 24) {real, imag} */,
  {32'hbe60568a, 32'hbdd488be} /* (6, 17, 23) {real, imag} */,
  {32'h3e0bcedd, 32'h3e45db8e} /* (6, 17, 22) {real, imag} */,
  {32'h3c201520, 32'hbe0c7cb5} /* (6, 17, 21) {real, imag} */,
  {32'h3f5bac1c, 32'hbe3f0a02} /* (6, 17, 20) {real, imag} */,
  {32'hbd4e231a, 32'h3ce105f4} /* (6, 17, 19) {real, imag} */,
  {32'hbe3d0bb8, 32'hbace8880} /* (6, 17, 18) {real, imag} */,
  {32'h3dcc515f, 32'hbd8277d0} /* (6, 17, 17) {real, imag} */,
  {32'h3d8f7799, 32'hbe672008} /* (6, 17, 16) {real, imag} */,
  {32'hbdf3b8c2, 32'h3e138784} /* (6, 17, 15) {real, imag} */,
  {32'h3dab3009, 32'h3ec146c8} /* (6, 17, 14) {real, imag} */,
  {32'h3e7b13e4, 32'hbce47030} /* (6, 17, 13) {real, imag} */,
  {32'hbe0f6dd6, 32'h3e4bf2c2} /* (6, 17, 12) {real, imag} */,
  {32'hbeafa412, 32'h3c44f178} /* (6, 17, 11) {real, imag} */,
  {32'hbea1d247, 32'hbd8cf674} /* (6, 17, 10) {real, imag} */,
  {32'hbe89a6a4, 32'hbee3382c} /* (6, 17, 9) {real, imag} */,
  {32'hbe801617, 32'hbd83cee5} /* (6, 17, 8) {real, imag} */,
  {32'hbec1223e, 32'h3eb34b8d} /* (6, 17, 7) {real, imag} */,
  {32'hbc4ce680, 32'hbdd7daca} /* (6, 17, 6) {real, imag} */,
  {32'hbe2e1419, 32'hbe1b375b} /* (6, 17, 5) {real, imag} */,
  {32'hbe464bdc, 32'hbe5ec928} /* (6, 17, 4) {real, imag} */,
  {32'h3e900784, 32'h3dd1e196} /* (6, 17, 3) {real, imag} */,
  {32'h3d59a640, 32'hbdbaa65e} /* (6, 17, 2) {real, imag} */,
  {32'hbdcc4072, 32'hbe7ea9b8} /* (6, 17, 1) {real, imag} */,
  {32'h3e3c5de9, 32'hbf05407f} /* (6, 17, 0) {real, imag} */,
  {32'h3e8eb71d, 32'h3e8e33a8} /* (6, 16, 31) {real, imag} */,
  {32'hbe17d354, 32'h3de395a8} /* (6, 16, 30) {real, imag} */,
  {32'hbdf90023, 32'h3d9a2dfe} /* (6, 16, 29) {real, imag} */,
  {32'hbeb17221, 32'h3e129320} /* (6, 16, 28) {real, imag} */,
  {32'hbeac5cc6, 32'h3e17071e} /* (6, 16, 27) {real, imag} */,
  {32'h3e3c0cbc, 32'h3d024932} /* (6, 16, 26) {real, imag} */,
  {32'h3e85dc86, 32'h3e367cea} /* (6, 16, 25) {real, imag} */,
  {32'h3c181170, 32'h3f04b9bd} /* (6, 16, 24) {real, imag} */,
  {32'hbe538b17, 32'hbe918f54} /* (6, 16, 23) {real, imag} */,
  {32'h3e81e50c, 32'hbe714794} /* (6, 16, 22) {real, imag} */,
  {32'hbc7aad38, 32'h3e869a4b} /* (6, 16, 21) {real, imag} */,
  {32'h3e18b88b, 32'h3e1505bc} /* (6, 16, 20) {real, imag} */,
  {32'h3e5c9502, 32'hbe80211a} /* (6, 16, 19) {real, imag} */,
  {32'h3ed3fafc, 32'hbeaa6044} /* (6, 16, 18) {real, imag} */,
  {32'hbdbd87f6, 32'h3ede7e4a} /* (6, 16, 17) {real, imag} */,
  {32'hbe83e90f, 32'h00000000} /* (6, 16, 16) {real, imag} */,
  {32'hbdbd87f6, 32'hbede7e4a} /* (6, 16, 15) {real, imag} */,
  {32'h3ed3fafc, 32'h3eaa6044} /* (6, 16, 14) {real, imag} */,
  {32'h3e5c9502, 32'h3e80211a} /* (6, 16, 13) {real, imag} */,
  {32'h3e18b88b, 32'hbe1505bc} /* (6, 16, 12) {real, imag} */,
  {32'hbc7aad38, 32'hbe869a4b} /* (6, 16, 11) {real, imag} */,
  {32'h3e81e50c, 32'h3e714794} /* (6, 16, 10) {real, imag} */,
  {32'hbe538b17, 32'h3e918f54} /* (6, 16, 9) {real, imag} */,
  {32'h3c181170, 32'hbf04b9bd} /* (6, 16, 8) {real, imag} */,
  {32'h3e85dc86, 32'hbe367cea} /* (6, 16, 7) {real, imag} */,
  {32'h3e3c0cbc, 32'hbd024932} /* (6, 16, 6) {real, imag} */,
  {32'hbeac5cc6, 32'hbe17071e} /* (6, 16, 5) {real, imag} */,
  {32'hbeb17221, 32'hbe129320} /* (6, 16, 4) {real, imag} */,
  {32'hbdf90023, 32'hbd9a2dfe} /* (6, 16, 3) {real, imag} */,
  {32'hbe17d354, 32'hbde395a8} /* (6, 16, 2) {real, imag} */,
  {32'h3e8eb71d, 32'hbe8e33a8} /* (6, 16, 1) {real, imag} */,
  {32'h3ebe759d, 32'h00000000} /* (6, 16, 0) {real, imag} */,
  {32'hbdcc4072, 32'h3e7ea9b8} /* (6, 15, 31) {real, imag} */,
  {32'h3d59a640, 32'h3dbaa65e} /* (6, 15, 30) {real, imag} */,
  {32'h3e900784, 32'hbdd1e196} /* (6, 15, 29) {real, imag} */,
  {32'hbe464bdc, 32'h3e5ec928} /* (6, 15, 28) {real, imag} */,
  {32'hbe2e1419, 32'h3e1b375b} /* (6, 15, 27) {real, imag} */,
  {32'hbc4ce680, 32'h3dd7daca} /* (6, 15, 26) {real, imag} */,
  {32'hbec1223e, 32'hbeb34b8d} /* (6, 15, 25) {real, imag} */,
  {32'hbe801617, 32'h3d83cee5} /* (6, 15, 24) {real, imag} */,
  {32'hbe89a6a4, 32'h3ee3382c} /* (6, 15, 23) {real, imag} */,
  {32'hbea1d247, 32'h3d8cf674} /* (6, 15, 22) {real, imag} */,
  {32'hbeafa412, 32'hbc44f178} /* (6, 15, 21) {real, imag} */,
  {32'hbe0f6dd6, 32'hbe4bf2c2} /* (6, 15, 20) {real, imag} */,
  {32'h3e7b13e4, 32'h3ce47030} /* (6, 15, 19) {real, imag} */,
  {32'h3dab3009, 32'hbec146c8} /* (6, 15, 18) {real, imag} */,
  {32'hbdf3b8c2, 32'hbe138784} /* (6, 15, 17) {real, imag} */,
  {32'h3d8f7799, 32'h3e672008} /* (6, 15, 16) {real, imag} */,
  {32'h3dcc515f, 32'h3d8277d0} /* (6, 15, 15) {real, imag} */,
  {32'hbe3d0bb8, 32'h3ace8880} /* (6, 15, 14) {real, imag} */,
  {32'hbd4e231a, 32'hbce105f4} /* (6, 15, 13) {real, imag} */,
  {32'h3f5bac1c, 32'h3e3f0a02} /* (6, 15, 12) {real, imag} */,
  {32'h3c201520, 32'h3e0c7cb5} /* (6, 15, 11) {real, imag} */,
  {32'h3e0bcedd, 32'hbe45db8e} /* (6, 15, 10) {real, imag} */,
  {32'hbe60568a, 32'h3dd488be} /* (6, 15, 9) {real, imag} */,
  {32'h3df092c6, 32'h3d7b747f} /* (6, 15, 8) {real, imag} */,
  {32'h3d52125a, 32'h3e689ea9} /* (6, 15, 7) {real, imag} */,
  {32'h3d0e4ec7, 32'hbe1f85e6} /* (6, 15, 6) {real, imag} */,
  {32'hbe232944, 32'h3e76c924} /* (6, 15, 5) {real, imag} */,
  {32'hbdd3b349, 32'hbeb4afaa} /* (6, 15, 4) {real, imag} */,
  {32'hbd028770, 32'h3e1f5162} /* (6, 15, 3) {real, imag} */,
  {32'hbbf3d8ac, 32'hbe83ae97} /* (6, 15, 2) {real, imag} */,
  {32'h3f1afcd5, 32'h3dd87615} /* (6, 15, 1) {real, imag} */,
  {32'h3e3c5de9, 32'h3f05407f} /* (6, 15, 0) {real, imag} */,
  {32'h3ec5b862, 32'hbf6842cb} /* (6, 14, 31) {real, imag} */,
  {32'hbe26fa77, 32'h3e8f1400} /* (6, 14, 30) {real, imag} */,
  {32'h3e098c6c, 32'h3ed3724e} /* (6, 14, 29) {real, imag} */,
  {32'h3d2e7a76, 32'h3e830567} /* (6, 14, 28) {real, imag} */,
  {32'h3d87038a, 32'h3e55fa26} /* (6, 14, 27) {real, imag} */,
  {32'hbb319e80, 32'h3e13b5b0} /* (6, 14, 26) {real, imag} */,
  {32'hbee78cb6, 32'hbd18e298} /* (6, 14, 25) {real, imag} */,
  {32'hbede746a, 32'hbf24235c} /* (6, 14, 24) {real, imag} */,
  {32'hbea37c36, 32'hbedae775} /* (6, 14, 23) {real, imag} */,
  {32'hbf134589, 32'hbee066d4} /* (6, 14, 22) {real, imag} */,
  {32'h3e81cbd8, 32'hbc7f4a1c} /* (6, 14, 21) {real, imag} */,
  {32'h3e25dc33, 32'h3f335d1c} /* (6, 14, 20) {real, imag} */,
  {32'hbe44d74e, 32'hbeb5534a} /* (6, 14, 19) {real, imag} */,
  {32'h3eaf5613, 32'hbe7a4688} /* (6, 14, 18) {real, imag} */,
  {32'hbe875ab4, 32'h3e483d84} /* (6, 14, 17) {real, imag} */,
  {32'hbe6ba45d, 32'h3de6018d} /* (6, 14, 16) {real, imag} */,
  {32'h3e924ea5, 32'h3e8982cb} /* (6, 14, 15) {real, imag} */,
  {32'h3df21caa, 32'h3e84c775} /* (6, 14, 14) {real, imag} */,
  {32'h3e54d026, 32'hbe21ca1a} /* (6, 14, 13) {real, imag} */,
  {32'hbd0fee60, 32'h3d2d7970} /* (6, 14, 12) {real, imag} */,
  {32'hbf71a9d2, 32'h39c59c00} /* (6, 14, 11) {real, imag} */,
  {32'h3ef25a54, 32'h3e23eecb} /* (6, 14, 10) {real, imag} */,
  {32'h3e1bb96e, 32'hbdc30c34} /* (6, 14, 9) {real, imag} */,
  {32'hbe841503, 32'hbc278f8c} /* (6, 14, 8) {real, imag} */,
  {32'hbea2c903, 32'h3e86e040} /* (6, 14, 7) {real, imag} */,
  {32'hbdf251f1, 32'h3edc36ab} /* (6, 14, 6) {real, imag} */,
  {32'hbd0f22ca, 32'h3ed2e9de} /* (6, 14, 5) {real, imag} */,
  {32'hbe9108cd, 32'hbd1482fe} /* (6, 14, 4) {real, imag} */,
  {32'h3e8e9177, 32'h3d86d5e0} /* (6, 14, 3) {real, imag} */,
  {32'h3ecac3cd, 32'h3e25643b} /* (6, 14, 2) {real, imag} */,
  {32'hbe82f185, 32'hbc40a250} /* (6, 14, 1) {real, imag} */,
  {32'hbd54305a, 32'hbe33f654} /* (6, 14, 0) {real, imag} */,
  {32'hbd48976c, 32'hbf124165} /* (6, 13, 31) {real, imag} */,
  {32'hbe55c405, 32'h3ae76e00} /* (6, 13, 30) {real, imag} */,
  {32'h3e8a05fc, 32'h3e577f42} /* (6, 13, 29) {real, imag} */,
  {32'hbd9f39d6, 32'hbe160674} /* (6, 13, 28) {real, imag} */,
  {32'hbee83e9e, 32'hbd60d5c8} /* (6, 13, 27) {real, imag} */,
  {32'hbca71a80, 32'h3b647d20} /* (6, 13, 26) {real, imag} */,
  {32'h3eacc9fc, 32'h3d9f30b1} /* (6, 13, 25) {real, imag} */,
  {32'h3d74bdd2, 32'h3e44d71c} /* (6, 13, 24) {real, imag} */,
  {32'h3dc007ec, 32'hbe83fdcd} /* (6, 13, 23) {real, imag} */,
  {32'h3eaf4f85, 32'hbe947e7c} /* (6, 13, 22) {real, imag} */,
  {32'hbe145755, 32'h3e3824ad} /* (6, 13, 21) {real, imag} */,
  {32'hbee00398, 32'hbe1adec6} /* (6, 13, 20) {real, imag} */,
  {32'h3e5b5c0c, 32'hbed388e0} /* (6, 13, 19) {real, imag} */,
  {32'hbe10d9d0, 32'h3e359d22} /* (6, 13, 18) {real, imag} */,
  {32'h3dca2956, 32'h3b74d020} /* (6, 13, 17) {real, imag} */,
  {32'h3d423c69, 32'h3e0b07aa} /* (6, 13, 16) {real, imag} */,
  {32'hbdb2cf15, 32'hbedacb83} /* (6, 13, 15) {real, imag} */,
  {32'h3dbf30cc, 32'h3d8aa9ac} /* (6, 13, 14) {real, imag} */,
  {32'hbed5dff2, 32'h3ea54b22} /* (6, 13, 13) {real, imag} */,
  {32'h3e4fd7c7, 32'hbdbf0d94} /* (6, 13, 12) {real, imag} */,
  {32'hbd831afc, 32'h3e9b34a4} /* (6, 13, 11) {real, imag} */,
  {32'hbe0332c3, 32'hbe32fdd0} /* (6, 13, 10) {real, imag} */,
  {32'hbf091b2a, 32'hbd9233cc} /* (6, 13, 9) {real, imag} */,
  {32'h3e753082, 32'h3eef2f3c} /* (6, 13, 8) {real, imag} */,
  {32'hbea5e8ff, 32'h3e873b4c} /* (6, 13, 7) {real, imag} */,
  {32'h3f05fd17, 32'hbe165e2c} /* (6, 13, 6) {real, imag} */,
  {32'h3e6b2508, 32'hbbce38c0} /* (6, 13, 5) {real, imag} */,
  {32'hbc1da860, 32'h3e462b30} /* (6, 13, 4) {real, imag} */,
  {32'hbc57e720, 32'hbd0de098} /* (6, 13, 3) {real, imag} */,
  {32'h3e6e07ef, 32'hbedb1e67} /* (6, 13, 2) {real, imag} */,
  {32'h3e8dbce0, 32'h3ee36ef1} /* (6, 13, 1) {real, imag} */,
  {32'h3e3a8ad4, 32'h3ef70261} /* (6, 13, 0) {real, imag} */,
  {32'h3e965b8e, 32'hbe92a665} /* (6, 12, 31) {real, imag} */,
  {32'hbdd5bb68, 32'hbe15d054} /* (6, 12, 30) {real, imag} */,
  {32'hbb5b9980, 32'hbd2447c0} /* (6, 12, 29) {real, imag} */,
  {32'h3e3ae797, 32'hbeab363d} /* (6, 12, 28) {real, imag} */,
  {32'h3eabe18c, 32'h3d2fa3a8} /* (6, 12, 27) {real, imag} */,
  {32'h3e4481cd, 32'h3e8256d8} /* (6, 12, 26) {real, imag} */,
  {32'hbedf9120, 32'h3e969f67} /* (6, 12, 25) {real, imag} */,
  {32'hbe784860, 32'hbe10cdfb} /* (6, 12, 24) {real, imag} */,
  {32'h3e3121b8, 32'hbe5c1c5f} /* (6, 12, 23) {real, imag} */,
  {32'h3e294351, 32'h3e0f4ea8} /* (6, 12, 22) {real, imag} */,
  {32'h3eb44244, 32'h3e211ca6} /* (6, 12, 21) {real, imag} */,
  {32'hbd65cd34, 32'hbee53052} /* (6, 12, 20) {real, imag} */,
  {32'h3e41eb62, 32'h3ed16cb2} /* (6, 12, 19) {real, imag} */,
  {32'h3e194d21, 32'hbd75cf3a} /* (6, 12, 18) {real, imag} */,
  {32'h3e99cc85, 32'hbe73e896} /* (6, 12, 17) {real, imag} */,
  {32'hbd0ddca4, 32'h3e57546a} /* (6, 12, 16) {real, imag} */,
  {32'h3e0d8432, 32'h3f0a4295} /* (6, 12, 15) {real, imag} */,
  {32'hbeb97bd8, 32'h3d12bcd6} /* (6, 12, 14) {real, imag} */,
  {32'h3e5a52e5, 32'hbecb18c0} /* (6, 12, 13) {real, imag} */,
  {32'h3d955a42, 32'hbef43535} /* (6, 12, 12) {real, imag} */,
  {32'hbe5cd7bf, 32'h3ca734b8} /* (6, 12, 11) {real, imag} */,
  {32'hbefec0df, 32'h3d0e52d4} /* (6, 12, 10) {real, imag} */,
  {32'h3e8747b1, 32'h3ea769fc} /* (6, 12, 9) {real, imag} */,
  {32'h3e567a64, 32'h3eed9831} /* (6, 12, 8) {real, imag} */,
  {32'h3eca39c4, 32'hbd988ce8} /* (6, 12, 7) {real, imag} */,
  {32'hbe2be016, 32'h3e6c3316} /* (6, 12, 6) {real, imag} */,
  {32'h3c8d16a8, 32'h3e230e64} /* (6, 12, 5) {real, imag} */,
  {32'h3e7f155f, 32'h3db1dc27} /* (6, 12, 4) {real, imag} */,
  {32'hbf03f567, 32'h3da882c2} /* (6, 12, 3) {real, imag} */,
  {32'hbd0fc158, 32'h3e1d2c56} /* (6, 12, 2) {real, imag} */,
  {32'hbe4ed62d, 32'hbedaa48c} /* (6, 12, 1) {real, imag} */,
  {32'hbe382c6d, 32'h3eaff3fb} /* (6, 12, 0) {real, imag} */,
  {32'hbeb4a1f9, 32'hbf1a9502} /* (6, 11, 31) {real, imag} */,
  {32'h3e24a528, 32'h3e6b88ba} /* (6, 11, 30) {real, imag} */,
  {32'hbdb6736e, 32'h3dc8e4e8} /* (6, 11, 29) {real, imag} */,
  {32'hbdb2f47c, 32'hbe2e7080} /* (6, 11, 28) {real, imag} */,
  {32'hbdeda93c, 32'h3db3c00e} /* (6, 11, 27) {real, imag} */,
  {32'h3e9140fd, 32'hbe948570} /* (6, 11, 26) {real, imag} */,
  {32'h3e9fa7ec, 32'hbeab5800} /* (6, 11, 25) {real, imag} */,
  {32'h3ec8ac3c, 32'h3e0fe6e7} /* (6, 11, 24) {real, imag} */,
  {32'h3ec0c697, 32'h3e50aa52} /* (6, 11, 23) {real, imag} */,
  {32'hbe738ee1, 32'h3ecb77a8} /* (6, 11, 22) {real, imag} */,
  {32'hbe8fefee, 32'h3f2fe4c0} /* (6, 11, 21) {real, imag} */,
  {32'hbe3e7283, 32'h3dc5ff8a} /* (6, 11, 20) {real, imag} */,
  {32'h3ea33bdf, 32'hbf2d7946} /* (6, 11, 19) {real, imag} */,
  {32'hbe07e2a4, 32'hbd99176c} /* (6, 11, 18) {real, imag} */,
  {32'hbe4458a1, 32'hbcb9c6b0} /* (6, 11, 17) {real, imag} */,
  {32'hbda44595, 32'h3d0ce07c} /* (6, 11, 16) {real, imag} */,
  {32'hba19d200, 32'h3ed45cfa} /* (6, 11, 15) {real, imag} */,
  {32'hbe22462e, 32'h3db9feb3} /* (6, 11, 14) {real, imag} */,
  {32'h3e4fae3a, 32'h3ed2e5a7} /* (6, 11, 13) {real, imag} */,
  {32'h3f082813, 32'h3da67abe} /* (6, 11, 12) {real, imag} */,
  {32'hbe9b0f5c, 32'h3c576300} /* (6, 11, 11) {real, imag} */,
  {32'hbe1024b4, 32'hbf03142c} /* (6, 11, 10) {real, imag} */,
  {32'hbd17ae9e, 32'hbf17bedd} /* (6, 11, 9) {real, imag} */,
  {32'hbe35955e, 32'h3ede14a7} /* (6, 11, 8) {real, imag} */,
  {32'hbec8d70a, 32'hbe9404d3} /* (6, 11, 7) {real, imag} */,
  {32'hbe11a11d, 32'hbe8557e7} /* (6, 11, 6) {real, imag} */,
  {32'h3e52859e, 32'hbc947108} /* (6, 11, 5) {real, imag} */,
  {32'hbe9fdb73, 32'h3f1a6a70} /* (6, 11, 4) {real, imag} */,
  {32'hbe7f92cc, 32'h3eb646dc} /* (6, 11, 3) {real, imag} */,
  {32'hbdd9996d, 32'h3f5beb42} /* (6, 11, 2) {real, imag} */,
  {32'hbd37f768, 32'hbf6db7e6} /* (6, 11, 1) {real, imag} */,
  {32'h3ec7da22, 32'hbea1e9e4} /* (6, 11, 0) {real, imag} */,
  {32'hbf1044d4, 32'h3e65fece} /* (6, 10, 31) {real, imag} */,
  {32'hbe645c46, 32'hbf7184d0} /* (6, 10, 30) {real, imag} */,
  {32'hbe2f7e17, 32'hbf269520} /* (6, 10, 29) {real, imag} */,
  {32'h3ecbc55e, 32'h3c0f17b4} /* (6, 10, 28) {real, imag} */,
  {32'h3d465e04, 32'h3d374894} /* (6, 10, 27) {real, imag} */,
  {32'h3ee7e346, 32'hbef31b00} /* (6, 10, 26) {real, imag} */,
  {32'h3d8ca2ac, 32'h3dd5916a} /* (6, 10, 25) {real, imag} */,
  {32'h3e4cce45, 32'hbed72acc} /* (6, 10, 24) {real, imag} */,
  {32'h3dc9d454, 32'hbd45b920} /* (6, 10, 23) {real, imag} */,
  {32'h3d6eeaf8, 32'h3f3229a6} /* (6, 10, 22) {real, imag} */,
  {32'hbe424b6a, 32'hbecadcae} /* (6, 10, 21) {real, imag} */,
  {32'hbe02e346, 32'hbe2e9ec9} /* (6, 10, 20) {real, imag} */,
  {32'hbe839fa8, 32'h3e224a5a} /* (6, 10, 19) {real, imag} */,
  {32'hbe7dd2f2, 32'h3cbbf0f0} /* (6, 10, 18) {real, imag} */,
  {32'h3e91f71c, 32'h3a557e40} /* (6, 10, 17) {real, imag} */,
  {32'hbe444769, 32'hbe700cda} /* (6, 10, 16) {real, imag} */,
  {32'hbd7339b6, 32'h3e549d4b} /* (6, 10, 15) {real, imag} */,
  {32'h3ea6951e, 32'h3f2780e8} /* (6, 10, 14) {real, imag} */,
  {32'hbf0d9cce, 32'h3e8925aa} /* (6, 10, 13) {real, imag} */,
  {32'hbe1ec6ba, 32'h3e61c4a4} /* (6, 10, 12) {real, imag} */,
  {32'h3ef500b2, 32'hbeb33171} /* (6, 10, 11) {real, imag} */,
  {32'hbf2d4f58, 32'h3f463174} /* (6, 10, 10) {real, imag} */,
  {32'hbefc7dad, 32'hbf2cf84a} /* (6, 10, 9) {real, imag} */,
  {32'h3eb1462a, 32'hbef306be} /* (6, 10, 8) {real, imag} */,
  {32'h3ed8df24, 32'h3e30fc8a} /* (6, 10, 7) {real, imag} */,
  {32'h3c85f5f0, 32'h3ebe755f} /* (6, 10, 6) {real, imag} */,
  {32'h3e4ab31c, 32'hbe95d26b} /* (6, 10, 5) {real, imag} */,
  {32'hbd156669, 32'h3e0e48ca} /* (6, 10, 4) {real, imag} */,
  {32'hbf00027c, 32'h3db07a14} /* (6, 10, 3) {real, imag} */,
  {32'hbed515e8, 32'hbf4d9bfa} /* (6, 10, 2) {real, imag} */,
  {32'h3f0ff111, 32'hbe51efee} /* (6, 10, 1) {real, imag} */,
  {32'hbea071da, 32'h3f86e6e9} /* (6, 10, 0) {real, imag} */,
  {32'hbda91446, 32'h3f560dc0} /* (6, 9, 31) {real, imag} */,
  {32'h3be3eb40, 32'h3e5eb6b6} /* (6, 9, 30) {real, imag} */,
  {32'hbec487f8, 32'hbee68f96} /* (6, 9, 29) {real, imag} */,
  {32'hbdd3a2d6, 32'h3f0db652} /* (6, 9, 28) {real, imag} */,
  {32'hbd4946c6, 32'h3e78137a} /* (6, 9, 27) {real, imag} */,
  {32'hbddb1b77, 32'hbefa202d} /* (6, 9, 26) {real, imag} */,
  {32'hbcc02e40, 32'h3e956fd3} /* (6, 9, 25) {real, imag} */,
  {32'hbe05a6f4, 32'h3eee75a0} /* (6, 9, 24) {real, imag} */,
  {32'h3d6528c9, 32'h3dc538a4} /* (6, 9, 23) {real, imag} */,
  {32'hbe11229d, 32'hbe9b054f} /* (6, 9, 22) {real, imag} */,
  {32'h3de46ef2, 32'hbecb4c3a} /* (6, 9, 21) {real, imag} */,
  {32'h3ee6138f, 32'h3f4ecede} /* (6, 9, 20) {real, imag} */,
  {32'hbf6ed2e7, 32'h3f052710} /* (6, 9, 19) {real, imag} */,
  {32'h3e8fcd0c, 32'hbcf701e0} /* (6, 9, 18) {real, imag} */,
  {32'hbe27da75, 32'h3f00523f} /* (6, 9, 17) {real, imag} */,
  {32'hbd61fe60, 32'h3ded0371} /* (6, 9, 16) {real, imag} */,
  {32'hbee71edd, 32'h3e5a9202} /* (6, 9, 15) {real, imag} */,
  {32'hbd2013cc, 32'h3d153b81} /* (6, 9, 14) {real, imag} */,
  {32'hbc6e6230, 32'h3e62c92f} /* (6, 9, 13) {real, imag} */,
  {32'hbccb9760, 32'h3e8be03e} /* (6, 9, 12) {real, imag} */,
  {32'hbe352fd7, 32'hbd431454} /* (6, 9, 11) {real, imag} */,
  {32'hbda39f27, 32'hbfb35d9a} /* (6, 9, 10) {real, imag} */,
  {32'h3e8a5192, 32'h3f109d0d} /* (6, 9, 9) {real, imag} */,
  {32'h3e54b958, 32'h3d1a0578} /* (6, 9, 8) {real, imag} */,
  {32'h3f00addf, 32'hbd3a01c8} /* (6, 9, 7) {real, imag} */,
  {32'h3e8a79d8, 32'h3e50e5e9} /* (6, 9, 6) {real, imag} */,
  {32'h3ec08947, 32'hbcf5cf70} /* (6, 9, 5) {real, imag} */,
  {32'hbe1a39c2, 32'hbf081570} /* (6, 9, 4) {real, imag} */,
  {32'h3f5c493b, 32'h3e88a96e} /* (6, 9, 3) {real, imag} */,
  {32'hbdf7f940, 32'hbf1459c4} /* (6, 9, 2) {real, imag} */,
  {32'h3cce5bf4, 32'h3e1c9553} /* (6, 9, 1) {real, imag} */,
  {32'hbec10ec0, 32'h3f12713c} /* (6, 9, 0) {real, imag} */,
  {32'hbf70afaa, 32'hbf22f0a1} /* (6, 8, 31) {real, imag} */,
  {32'h3f19af10, 32'h3df0a2e7} /* (6, 8, 30) {real, imag} */,
  {32'h3ed0e104, 32'h3f2c9af2} /* (6, 8, 29) {real, imag} */,
  {32'hbf2c51df, 32'h3f11b442} /* (6, 8, 28) {real, imag} */,
  {32'h3f39e2a0, 32'hbeeb7a88} /* (6, 8, 27) {real, imag} */,
  {32'h3d57a6c8, 32'hbe0c094a} /* (6, 8, 26) {real, imag} */,
  {32'hbbcbe340, 32'hbeb63465} /* (6, 8, 25) {real, imag} */,
  {32'h3eb2582e, 32'hbe9dcacc} /* (6, 8, 24) {real, imag} */,
  {32'h3e937530, 32'h3d8adae6} /* (6, 8, 23) {real, imag} */,
  {32'hbdfd1440, 32'h3e5a7b1a} /* (6, 8, 22) {real, imag} */,
  {32'h3ed2de4a, 32'h3e376523} /* (6, 8, 21) {real, imag} */,
  {32'hbe84844e, 32'hbdc8abd2} /* (6, 8, 20) {real, imag} */,
  {32'h3e23beff, 32'h3df827ee} /* (6, 8, 19) {real, imag} */,
  {32'hbd8644c8, 32'hbdb0405b} /* (6, 8, 18) {real, imag} */,
  {32'hbe7f0707, 32'h3c1366a0} /* (6, 8, 17) {real, imag} */,
  {32'h3e6cc261, 32'h3e8837df} /* (6, 8, 16) {real, imag} */,
  {32'h3ea793e2, 32'h3e9f2b87} /* (6, 8, 15) {real, imag} */,
  {32'h3e15d88f, 32'hbeb24ddb} /* (6, 8, 14) {real, imag} */,
  {32'h3e29b190, 32'hbd37515a} /* (6, 8, 13) {real, imag} */,
  {32'h3cb8a91e, 32'h3ebeaca8} /* (6, 8, 12) {real, imag} */,
  {32'h3e9a4d44, 32'h3e70dc23} /* (6, 8, 11) {real, imag} */,
  {32'hbe2ef400, 32'hbb1cf000} /* (6, 8, 10) {real, imag} */,
  {32'hbf028819, 32'h3f08bd20} /* (6, 8, 9) {real, imag} */,
  {32'hbd8591a4, 32'h3f0a90ec} /* (6, 8, 8) {real, imag} */,
  {32'h3e1c97c8, 32'h3dc3b98c} /* (6, 8, 7) {real, imag} */,
  {32'hbf42933c, 32'h3db61ffd} /* (6, 8, 6) {real, imag} */,
  {32'hbf070efe, 32'h3e43ea96} /* (6, 8, 5) {real, imag} */,
  {32'hbed68347, 32'hbefc68f3} /* (6, 8, 4) {real, imag} */,
  {32'h3d528dc0, 32'h3e577852} /* (6, 8, 3) {real, imag} */,
  {32'h3f6dbb79, 32'h3ea4b57d} /* (6, 8, 2) {real, imag} */,
  {32'hbf694d0c, 32'hbf480658} /* (6, 8, 1) {real, imag} */,
  {32'hbf72cf56, 32'hbf87d76e} /* (6, 8, 0) {real, imag} */,
  {32'h3f08278e, 32'h3f1b5262} /* (6, 7, 31) {real, imag} */,
  {32'hbd9232a4, 32'h3efade4b} /* (6, 7, 30) {real, imag} */,
  {32'hbef274f6, 32'h3ee590e5} /* (6, 7, 29) {real, imag} */,
  {32'hbf56b4e8, 32'hbe01b000} /* (6, 7, 28) {real, imag} */,
  {32'hbd83be64, 32'h3f12afb1} /* (6, 7, 27) {real, imag} */,
  {32'hbf223f48, 32'hbc7113c0} /* (6, 7, 26) {real, imag} */,
  {32'h3ea9dc72, 32'hbf2e2f00} /* (6, 7, 25) {real, imag} */,
  {32'h3e2a2e4a, 32'hbd4c0168} /* (6, 7, 24) {real, imag} */,
  {32'hbedc88d2, 32'h3de44d00} /* (6, 7, 23) {real, imag} */,
  {32'hbe6106c7, 32'h3f4cfa39} /* (6, 7, 22) {real, imag} */,
  {32'h3e7eebc2, 32'h3d692808} /* (6, 7, 21) {real, imag} */,
  {32'hbe03e732, 32'hbea979fe} /* (6, 7, 20) {real, imag} */,
  {32'hbee8c74a, 32'h3ebda0e6} /* (6, 7, 19) {real, imag} */,
  {32'h3d834462, 32'hbf0c8496} /* (6, 7, 18) {real, imag} */,
  {32'hbc94f88a, 32'hbe5173dc} /* (6, 7, 17) {real, imag} */,
  {32'hbef72f22, 32'hbd8f89d1} /* (6, 7, 16) {real, imag} */,
  {32'hbeccd932, 32'h3e5119ce} /* (6, 7, 15) {real, imag} */,
  {32'h3e848564, 32'hbd562005} /* (6, 7, 14) {real, imag} */,
  {32'h3e8b6d3c, 32'h3d8215d1} /* (6, 7, 13) {real, imag} */,
  {32'hbcc11de0, 32'hbe07f729} /* (6, 7, 12) {real, imag} */,
  {32'hbe16216c, 32'hbde5748e} /* (6, 7, 11) {real, imag} */,
  {32'h3ce27ac0, 32'hbe1385b9} /* (6, 7, 10) {real, imag} */,
  {32'h3f180028, 32'h3d6a490c} /* (6, 7, 9) {real, imag} */,
  {32'hbdfde2d2, 32'h3e70d761} /* (6, 7, 8) {real, imag} */,
  {32'hbd2c60c8, 32'h3e331cb9} /* (6, 7, 7) {real, imag} */,
  {32'h3f43ecb4, 32'h3e32e572} /* (6, 7, 6) {real, imag} */,
  {32'h3ed30722, 32'hbdf5e6c2} /* (6, 7, 5) {real, imag} */,
  {32'h3f196716, 32'h3edf5b22} /* (6, 7, 4) {real, imag} */,
  {32'h3d3921c8, 32'h3ea8c78a} /* (6, 7, 3) {real, imag} */,
  {32'h3e2e506c, 32'hbf25af8c} /* (6, 7, 2) {real, imag} */,
  {32'hbe25e802, 32'h3f2a930f} /* (6, 7, 1) {real, imag} */,
  {32'h3e7f5802, 32'hbdf08bed} /* (6, 7, 0) {real, imag} */,
  {32'h3ec7d0d2, 32'h3f3dc1ec} /* (6, 6, 31) {real, imag} */,
  {32'hbeda9cf6, 32'hbf1195f0} /* (6, 6, 30) {real, imag} */,
  {32'hbe98f380, 32'h3ddae2c4} /* (6, 6, 29) {real, imag} */,
  {32'h3e747737, 32'hbe7202ba} /* (6, 6, 28) {real, imag} */,
  {32'hbd36bffc, 32'h3e77c3e6} /* (6, 6, 27) {real, imag} */,
  {32'h3f053e5a, 32'hbea2980e} /* (6, 6, 26) {real, imag} */,
  {32'h3e8cc555, 32'h3f058720} /* (6, 6, 25) {real, imag} */,
  {32'hbd021c32, 32'hbd200d60} /* (6, 6, 24) {real, imag} */,
  {32'hbd8b0936, 32'hbf0a3c23} /* (6, 6, 23) {real, imag} */,
  {32'h3e13aefc, 32'h3dcc3652} /* (6, 6, 22) {real, imag} */,
  {32'hbede5b16, 32'hbe88b3ef} /* (6, 6, 21) {real, imag} */,
  {32'h3d0cbbc6, 32'h3da87c12} /* (6, 6, 20) {real, imag} */,
  {32'hbe85bcb2, 32'hbf2c5708} /* (6, 6, 19) {real, imag} */,
  {32'h3e0ed292, 32'h3ea61958} /* (6, 6, 18) {real, imag} */,
  {32'hbf22b1f6, 32'hbef07c04} /* (6, 6, 17) {real, imag} */,
  {32'hbd32243c, 32'h3d8431d0} /* (6, 6, 16) {real, imag} */,
  {32'h3a236900, 32'h3e89df2c} /* (6, 6, 15) {real, imag} */,
  {32'hbd27852a, 32'hbdf1f654} /* (6, 6, 14) {real, imag} */,
  {32'hbdf8291c, 32'hbe6cdc0a} /* (6, 6, 13) {real, imag} */,
  {32'hbe09dd10, 32'hbe049a1f} /* (6, 6, 12) {real, imag} */,
  {32'h3ed5870c, 32'hbca19fd0} /* (6, 6, 11) {real, imag} */,
  {32'h3e47178b, 32'h3e5809a2} /* (6, 6, 10) {real, imag} */,
  {32'h3dccd7a8, 32'h3f42697a} /* (6, 6, 9) {real, imag} */,
  {32'h3cc6d490, 32'h3e815a9a} /* (6, 6, 8) {real, imag} */,
  {32'h3f4354a0, 32'hbec22846} /* (6, 6, 7) {real, imag} */,
  {32'hba791200, 32'h3ea9fe2c} /* (6, 6, 6) {real, imag} */,
  {32'hbe752a8c, 32'h3ed241eb} /* (6, 6, 5) {real, imag} */,
  {32'h3e9b2dc6, 32'h3e1521bc} /* (6, 6, 4) {real, imag} */,
  {32'hbf3a26b1, 32'hbf1fc4f8} /* (6, 6, 3) {real, imag} */,
  {32'hbfb23dbd, 32'h3eb87a7e} /* (6, 6, 2) {real, imag} */,
  {32'hbf725449, 32'h3f3a5230} /* (6, 6, 1) {real, imag} */,
  {32'h3cf6d520, 32'hbf391890} /* (6, 6, 0) {real, imag} */,
  {32'hbfe929f8, 32'h3fb528e2} /* (6, 5, 31) {real, imag} */,
  {32'h3fc61b96, 32'h3f259a98} /* (6, 5, 30) {real, imag} */,
  {32'hbf1598a2, 32'h3de25794} /* (6, 5, 29) {real, imag} */,
  {32'hbf9219f4, 32'hbe2db710} /* (6, 5, 28) {real, imag} */,
  {32'h3f840590, 32'h3ed45966} /* (6, 5, 27) {real, imag} */,
  {32'h3e23f8b1, 32'hbd7b6f42} /* (6, 5, 26) {real, imag} */,
  {32'hbe1b52d6, 32'h3e4b9210} /* (6, 5, 25) {real, imag} */,
  {32'hbe704bf9, 32'h3e7a7c4f} /* (6, 5, 24) {real, imag} */,
  {32'h3d8ebfca, 32'hbe0d85e3} /* (6, 5, 23) {real, imag} */,
  {32'hbef62ffc, 32'h3f3ef540} /* (6, 5, 22) {real, imag} */,
  {32'h3e6ea60b, 32'hbf5a0ec7} /* (6, 5, 21) {real, imag} */,
  {32'h3ea41177, 32'hbed80c18} /* (6, 5, 20) {real, imag} */,
  {32'hbde26f96, 32'hbeb253e6} /* (6, 5, 19) {real, imag} */,
  {32'hbb075d60, 32'hbd7046f4} /* (6, 5, 18) {real, imag} */,
  {32'hbe7662e1, 32'h3d0164ac} /* (6, 5, 17) {real, imag} */,
  {32'h3b26b440, 32'hbe5d36f9} /* (6, 5, 16) {real, imag} */,
  {32'h3d49d02c, 32'hba0529c0} /* (6, 5, 15) {real, imag} */,
  {32'h3d16ab78, 32'h3d8f2bf4} /* (6, 5, 14) {real, imag} */,
  {32'h3e57544c, 32'h3eab5fde} /* (6, 5, 13) {real, imag} */,
  {32'hbe6fae90, 32'hbf3e7872} /* (6, 5, 12) {real, imag} */,
  {32'h3eb0dca6, 32'h3eb7c138} /* (6, 5, 11) {real, imag} */,
  {32'hbe242274, 32'h3e9dfa80} /* (6, 5, 10) {real, imag} */,
  {32'hbe98c2e6, 32'hbe891009} /* (6, 5, 9) {real, imag} */,
  {32'h3dd63eac, 32'hbecbdfd9} /* (6, 5, 8) {real, imag} */,
  {32'hbe8bff0d, 32'hbdf9e8f8} /* (6, 5, 7) {real, imag} */,
  {32'h3ec310f8, 32'h3e8564d2} /* (6, 5, 6) {real, imag} */,
  {32'h3d833d94, 32'h3e727dc0} /* (6, 5, 5) {real, imag} */,
  {32'hbe37f7a2, 32'hbeabd8e5} /* (6, 5, 4) {real, imag} */,
  {32'hbb4ec240, 32'h3ecff8c1} /* (6, 5, 3) {real, imag} */,
  {32'h3f6b0e63, 32'h3f9b3060} /* (6, 5, 2) {real, imag} */,
  {32'hbf08b77c, 32'hbfd01214} /* (6, 5, 1) {real, imag} */,
  {32'hbfdde6d8, 32'hbf602773} /* (6, 5, 0) {real, imag} */,
  {32'h3e971e0e, 32'h3fde02ae} /* (6, 4, 31) {real, imag} */,
  {32'hbfb6af96, 32'hbfd036cd} /* (6, 4, 30) {real, imag} */,
  {32'h3e8e828e, 32'h3ec496fe} /* (6, 4, 29) {real, imag} */,
  {32'h3eb9a3ff, 32'hbed341c9} /* (6, 4, 28) {real, imag} */,
  {32'h3d700f0a, 32'h3ec44c9e} /* (6, 4, 27) {real, imag} */,
  {32'h3d8a21b4, 32'hbf1ae96e} /* (6, 4, 26) {real, imag} */,
  {32'hbdb25355, 32'h3e84d2ef} /* (6, 4, 25) {real, imag} */,
  {32'hbf2270ce, 32'hbe69add8} /* (6, 4, 24) {real, imag} */,
  {32'hbe796c39, 32'hbe09e54c} /* (6, 4, 23) {real, imag} */,
  {32'hbf1a3ab7, 32'hbd414a5a} /* (6, 4, 22) {real, imag} */,
  {32'h3ea4f472, 32'h3d7dfa78} /* (6, 4, 21) {real, imag} */,
  {32'h3ef6841e, 32'hbc71e348} /* (6, 4, 20) {real, imag} */,
  {32'hbd7049ac, 32'hbdef67c2} /* (6, 4, 19) {real, imag} */,
  {32'h3edc3030, 32'hbec33461} /* (6, 4, 18) {real, imag} */,
  {32'h3e6d938a, 32'hbddd3a06} /* (6, 4, 17) {real, imag} */,
  {32'hbdbba422, 32'h3e478412} /* (6, 4, 16) {real, imag} */,
  {32'hbe40b34d, 32'h3e99a613} /* (6, 4, 15) {real, imag} */,
  {32'h3ce36570, 32'hbed94274} /* (6, 4, 14) {real, imag} */,
  {32'h3ed482d6, 32'hbf145c59} /* (6, 4, 13) {real, imag} */,
  {32'hbc915ad0, 32'h3f427f36} /* (6, 4, 12) {real, imag} */,
  {32'h3d3fa660, 32'hbdf82686} /* (6, 4, 11) {real, imag} */,
  {32'hbea01d00, 32'h3d84a154} /* (6, 4, 10) {real, imag} */,
  {32'h3ef00d3c, 32'hbed13acf} /* (6, 4, 9) {real, imag} */,
  {32'hbf3a7c42, 32'h3eb384fd} /* (6, 4, 8) {real, imag} */,
  {32'h3dbeec46, 32'h3d832086} /* (6, 4, 7) {real, imag} */,
  {32'hbefad5f8, 32'h3f705d98} /* (6, 4, 6) {real, imag} */,
  {32'hbf0b23d4, 32'hbedf882c} /* (6, 4, 5) {real, imag} */,
  {32'h3e8935ba, 32'h3f1139ee} /* (6, 4, 4) {real, imag} */,
  {32'hbe8cc302, 32'h3e2bf7cc} /* (6, 4, 3) {real, imag} */,
  {32'hbfdb88d7, 32'hbfc63d81} /* (6, 4, 2) {real, imag} */,
  {32'h3fe94d46, 32'h40122f85} /* (6, 4, 1) {real, imag} */,
  {32'h3fbff7ff, 32'hbe6215a8} /* (6, 4, 0) {real, imag} */,
  {32'hc03b06ef, 32'h3f75c638} /* (6, 3, 31) {real, imag} */,
  {32'h3f1eac7a, 32'hc07caf3a} /* (6, 3, 30) {real, imag} */,
  {32'h3e575f26, 32'hbc230910} /* (6, 3, 29) {real, imag} */,
  {32'h3f4e4a34, 32'h3f54a4a1} /* (6, 3, 28) {real, imag} */,
  {32'h3e1591c0, 32'hbe3fc9e7} /* (6, 3, 27) {real, imag} */,
  {32'hbf912008, 32'h3e665e23} /* (6, 3, 26) {real, imag} */,
  {32'hbcebe0a0, 32'hbe95739a} /* (6, 3, 25) {real, imag} */,
  {32'h3e8637ef, 32'hbf32ed8c} /* (6, 3, 24) {real, imag} */,
  {32'h3e8eb618, 32'hbda4a6cc} /* (6, 3, 23) {real, imag} */,
  {32'h3c507750, 32'hbe1d62cf} /* (6, 3, 22) {real, imag} */,
  {32'hbe9cd648, 32'h3ef3e68d} /* (6, 3, 21) {real, imag} */,
  {32'hbdb5145c, 32'h3ea5aad0} /* (6, 3, 20) {real, imag} */,
  {32'h3f23faa6, 32'h3eb90170} /* (6, 3, 19) {real, imag} */,
  {32'hbd26261c, 32'hbe1f8920} /* (6, 3, 18) {real, imag} */,
  {32'h3eb11e3c, 32'h3e484078} /* (6, 3, 17) {real, imag} */,
  {32'hbccab9f4, 32'h3d64e2ca} /* (6, 3, 16) {real, imag} */,
  {32'hbed1dd8e, 32'h3e8c2277} /* (6, 3, 15) {real, imag} */,
  {32'h3f4bcf8a, 32'h3e3ae89a} /* (6, 3, 14) {real, imag} */,
  {32'h3d86d394, 32'hbea7f34b} /* (6, 3, 13) {real, imag} */,
  {32'hbdb9026c, 32'hbeea9420} /* (6, 3, 12) {real, imag} */,
  {32'h3efea02c, 32'h3ccfda6c} /* (6, 3, 11) {real, imag} */,
  {32'hbf150e76, 32'h3e4fa509} /* (6, 3, 10) {real, imag} */,
  {32'h3f148835, 32'h3d2958d0} /* (6, 3, 9) {real, imag} */,
  {32'hbefbed88, 32'hbf199556} /* (6, 3, 8) {real, imag} */,
  {32'hbea18e82, 32'h3d9f6da6} /* (6, 3, 7) {real, imag} */,
  {32'h3dafb600, 32'hbf8e3130} /* (6, 3, 6) {real, imag} */,
  {32'h3f75f994, 32'hbf549451} /* (6, 3, 5) {real, imag} */,
  {32'hbf51e1ba, 32'h3e8b9f11} /* (6, 3, 4) {real, imag} */,
  {32'hbf4c68e0, 32'hbebcb546} /* (6, 3, 3) {real, imag} */,
  {32'h3e3c4c3c, 32'hbeb546da} /* (6, 3, 2) {real, imag} */,
  {32'h40345df8, 32'h406d5064} /* (6, 3, 1) {real, imag} */,
  {32'h3f45c137, 32'h4001562d} /* (6, 3, 0) {real, imag} */,
  {32'hc19ffd87, 32'hbd449930} /* (6, 2, 31) {real, imag} */,
  {32'h41307012, 32'hc02c400d} /* (6, 2, 30) {real, imag} */,
  {32'hbfc88758, 32'h3f9287ec} /* (6, 2, 29) {real, imag} */,
  {32'h3e894bd4, 32'h3f76120d} /* (6, 2, 28) {real, imag} */,
  {32'h3f308e0d, 32'hbf7c1d8b} /* (6, 2, 27) {real, imag} */,
  {32'h3e81b47c, 32'h3d055b60} /* (6, 2, 26) {real, imag} */,
  {32'hbdcaef3c, 32'hbe96ee08} /* (6, 2, 25) {real, imag} */,
  {32'h3fad6493, 32'h3ea87c6b} /* (6, 2, 24) {real, imag} */,
  {32'hbef8c1be, 32'h3cf957e0} /* (6, 2, 23) {real, imag} */,
  {32'h3c32a800, 32'hbd928536} /* (6, 2, 22) {real, imag} */,
  {32'h3dc58a1d, 32'hbf03d576} /* (6, 2, 21) {real, imag} */,
  {32'h3d44a074, 32'h3eca98a3} /* (6, 2, 20) {real, imag} */,
  {32'h3e7990fa, 32'h3e9849d3} /* (6, 2, 19) {real, imag} */,
  {32'hbeb67104, 32'hbec8d701} /* (6, 2, 18) {real, imag} */,
  {32'hbdd0d590, 32'h3dd68cb6} /* (6, 2, 17) {real, imag} */,
  {32'hbb96e840, 32'hbce291a8} /* (6, 2, 16) {real, imag} */,
  {32'h3dbf3712, 32'hbe86dd8c} /* (6, 2, 15) {real, imag} */,
  {32'h3e38db14, 32'h3db5f704} /* (6, 2, 14) {real, imag} */,
  {32'h3d981f1e, 32'hbcffed15} /* (6, 2, 13) {real, imag} */,
  {32'hbebc19f0, 32'hbdb15e10} /* (6, 2, 12) {real, imag} */,
  {32'h3eae24dc, 32'h3f3dc8dc} /* (6, 2, 11) {real, imag} */,
  {32'h3e47f755, 32'hbd57fb10} /* (6, 2, 10) {real, imag} */,
  {32'h3ec30072, 32'h3ef2c842} /* (6, 2, 9) {real, imag} */,
  {32'h3f586070, 32'h3e1d26fc} /* (6, 2, 8) {real, imag} */,
  {32'hbe16b2b2, 32'hbf031a6c} /* (6, 2, 7) {real, imag} */,
  {32'h3e28c640, 32'h3f094c50} /* (6, 2, 6) {real, imag} */,
  {32'h3fb40b32, 32'h3e96e888} /* (6, 2, 5) {real, imag} */,
  {32'hc02e24a7, 32'hbda2a7b0} /* (6, 2, 4) {real, imag} */,
  {32'hbee67c55, 32'h3fa03d1e} /* (6, 2, 3) {real, imag} */,
  {32'h40d87e37, 32'hbd4528c0} /* (6, 2, 2) {real, imag} */,
  {32'hc11ecffa, 32'h4027fa80} /* (6, 2, 1) {real, imag} */,
  {32'hc12ed24a, 32'hc0925213} /* (6, 2, 0) {real, imag} */,
  {32'h41de82cb, 32'hc0f286c0} /* (6, 1, 31) {real, imag} */,
  {32'hc0b93089, 32'hbc345180} /* (6, 1, 30) {real, imag} */,
  {32'h40049d73, 32'hbf05217f} /* (6, 1, 29) {real, imag} */,
  {32'h3fbed70e, 32'h3fc619ab} /* (6, 1, 28) {real, imag} */,
  {32'hc0374f0c, 32'hbee28e0a} /* (6, 1, 27) {real, imag} */,
  {32'h3ec17d26, 32'h3ddfc2fa} /* (6, 1, 26) {real, imag} */,
  {32'hbf093dee, 32'hbd326728} /* (6, 1, 25) {real, imag} */,
  {32'hbf2f5090, 32'h3e2bc1d1} /* (6, 1, 24) {real, imag} */,
  {32'h3d492f8c, 32'hbee4a539} /* (6, 1, 23) {real, imag} */,
  {32'h3eaf1eac, 32'hbe73cda2} /* (6, 1, 22) {real, imag} */,
  {32'hbf2b8a8c, 32'h3f80b772} /* (6, 1, 21) {real, imag} */,
  {32'h3eebc1d6, 32'h3e3de156} /* (6, 1, 20) {real, imag} */,
  {32'h3d9c0e6e, 32'hbe826814} /* (6, 1, 19) {real, imag} */,
  {32'hbef69b04, 32'h3e055a8b} /* (6, 1, 18) {real, imag} */,
  {32'h3dcb5712, 32'h3de78f7a} /* (6, 1, 17) {real, imag} */,
  {32'hbe6b0cce, 32'h3dde0e18} /* (6, 1, 16) {real, imag} */,
  {32'hbea13968, 32'h3da5f118} /* (6, 1, 15) {real, imag} */,
  {32'h3e8d0e80, 32'hbf007478} /* (6, 1, 14) {real, imag} */,
  {32'h3c2fa580, 32'h3d3ad3db} /* (6, 1, 13) {real, imag} */,
  {32'hbd90ba32, 32'h3d48daac} /* (6, 1, 12) {real, imag} */,
  {32'hbf1db160, 32'hbf3e8369} /* (6, 1, 11) {real, imag} */,
  {32'hbe9af5bc, 32'hbd8c86b1} /* (6, 1, 10) {real, imag} */,
  {32'h3eae01e9, 32'hbb8a9480} /* (6, 1, 9) {real, imag} */,
  {32'hbea4d526, 32'hbf86c0c2} /* (6, 1, 8) {real, imag} */,
  {32'h3f430ac0, 32'h3e626ffa} /* (6, 1, 7) {real, imag} */,
  {32'hbef51b62, 32'hbd1dba94} /* (6, 1, 6) {real, imag} */,
  {32'hbff02b8e, 32'hbe98e236} /* (6, 1, 5) {real, imag} */,
  {32'h3fc182cd, 32'hbf5536de} /* (6, 1, 4) {real, imag} */,
  {32'hbf2575ee, 32'hc007893d} /* (6, 1, 3) {real, imag} */,
  {32'hc124e64a, 32'hc11b9bf8} /* (6, 1, 2) {real, imag} */,
  {32'h421cbd4a, 32'h41881355} /* (6, 1, 1) {real, imag} */,
  {32'h421fd30a, 32'h40eb3175} /* (6, 1, 0) {real, imag} */,
  {32'h41b4b0b3, 32'hc19ddcf1} /* (6, 0, 31) {real, imag} */,
  {32'hbfa79c50, 32'h40a7e5d8} /* (6, 0, 30) {real, imag} */,
  {32'h3f12fde1, 32'hbfac198c} /* (6, 0, 29) {real, imag} */,
  {32'h3da06320, 32'hbfaaa057} /* (6, 0, 28) {real, imag} */,
  {32'hbf9de18c, 32'h3f0d89e8} /* (6, 0, 27) {real, imag} */,
  {32'h3f50e4d7, 32'h3e57dbc4} /* (6, 0, 26) {real, imag} */,
  {32'h3f48a551, 32'hbf9805d5} /* (6, 0, 25) {real, imag} */,
  {32'hbe2ad428, 32'h3e8bf166} /* (6, 0, 24) {real, imag} */,
  {32'hbf1e1595, 32'h3e1ada58} /* (6, 0, 23) {real, imag} */,
  {32'hbdea688c, 32'hbe798d73} /* (6, 0, 22) {real, imag} */,
  {32'hbf009f9b, 32'h3f1a9d37} /* (6, 0, 21) {real, imag} */,
  {32'h3e842066, 32'hbe545dd4} /* (6, 0, 20) {real, imag} */,
  {32'h3eb47180, 32'h3efacb18} /* (6, 0, 19) {real, imag} */,
  {32'hbe4c7530, 32'h3ee84676} /* (6, 0, 18) {real, imag} */,
  {32'hbd984504, 32'h3cfd14f2} /* (6, 0, 17) {real, imag} */,
  {32'h3eb6c008, 32'h00000000} /* (6, 0, 16) {real, imag} */,
  {32'hbd984504, 32'hbcfd14f2} /* (6, 0, 15) {real, imag} */,
  {32'hbe4c7530, 32'hbee84676} /* (6, 0, 14) {real, imag} */,
  {32'h3eb47180, 32'hbefacb18} /* (6, 0, 13) {real, imag} */,
  {32'h3e842066, 32'h3e545dd4} /* (6, 0, 12) {real, imag} */,
  {32'hbf009f9b, 32'hbf1a9d37} /* (6, 0, 11) {real, imag} */,
  {32'hbdea688c, 32'h3e798d73} /* (6, 0, 10) {real, imag} */,
  {32'hbf1e1595, 32'hbe1ada58} /* (6, 0, 9) {real, imag} */,
  {32'hbe2ad428, 32'hbe8bf166} /* (6, 0, 8) {real, imag} */,
  {32'h3f48a551, 32'h3f9805d5} /* (6, 0, 7) {real, imag} */,
  {32'h3f50e4d7, 32'hbe57dbc4} /* (6, 0, 6) {real, imag} */,
  {32'hbf9de18c, 32'hbf0d89e8} /* (6, 0, 5) {real, imag} */,
  {32'h3da06320, 32'h3faaa057} /* (6, 0, 4) {real, imag} */,
  {32'h3f12fde1, 32'h3fac198c} /* (6, 0, 3) {real, imag} */,
  {32'hbfa79c50, 32'hc0a7e5d8} /* (6, 0, 2) {real, imag} */,
  {32'h41b4b0b3, 32'h419ddcf1} /* (6, 0, 1) {real, imag} */,
  {32'h42434370, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'h413db712, 32'hbfee91b4} /* (5, 31, 31) {real, imag} */,
  {32'hbe5733e0, 32'h3ee0f640} /* (5, 31, 30) {real, imag} */,
  {32'hbe8d3652, 32'h3fdc2658} /* (5, 31, 29) {real, imag} */,
  {32'h3f4ad6a5, 32'h3f8f0810} /* (5, 31, 28) {real, imag} */,
  {32'hbeae5fb8, 32'hbf38a617} /* (5, 31, 27) {real, imag} */,
  {32'hbf2ee3e4, 32'h3ece317d} /* (5, 31, 26) {real, imag} */,
  {32'hbe25dcbc, 32'hbf058868} /* (5, 31, 25) {real, imag} */,
  {32'h3f5a4d77, 32'hbe683474} /* (5, 31, 24) {real, imag} */,
  {32'hbf09c200, 32'hbedb87cb} /* (5, 31, 23) {real, imag} */,
  {32'hbe8c54b5, 32'h3ea38f9a} /* (5, 31, 22) {real, imag} */,
  {32'h3ed92f8f, 32'h3ec2139a} /* (5, 31, 21) {real, imag} */,
  {32'h3e4e8303, 32'h3d9a8872} /* (5, 31, 20) {real, imag} */,
  {32'h3ea3cbba, 32'hbe174527} /* (5, 31, 19) {real, imag} */,
  {32'h3e977e17, 32'h3ea9c5c3} /* (5, 31, 18) {real, imag} */,
  {32'h3e0d8ff3, 32'hbe2f6c15} /* (5, 31, 17) {real, imag} */,
  {32'h3d804ef8, 32'h3e329433} /* (5, 31, 16) {real, imag} */,
  {32'h3dc76a4a, 32'h3c5a9ad0} /* (5, 31, 15) {real, imag} */,
  {32'hbe0f312c, 32'h3eb0c575} /* (5, 31, 14) {real, imag} */,
  {32'h3d83e909, 32'h3e8817c7} /* (5, 31, 13) {real, imag} */,
  {32'h3e323de7, 32'h3ec0ed13} /* (5, 31, 12) {real, imag} */,
  {32'hbe8faa5a, 32'hbb5df380} /* (5, 31, 11) {real, imag} */,
  {32'hbdf2237e, 32'h3dbcf99a} /* (5, 31, 10) {real, imag} */,
  {32'h3ed8dd67, 32'h3e8f8268} /* (5, 31, 9) {real, imag} */,
  {32'h3df48864, 32'h3e945451} /* (5, 31, 8) {real, imag} */,
  {32'hbfabb13e, 32'h3deb6a01} /* (5, 31, 7) {real, imag} */,
  {32'h3e962453, 32'h3ebb854e} /* (5, 31, 6) {real, imag} */,
  {32'h3f0af44c, 32'hbedf17a4} /* (5, 31, 5) {real, imag} */,
  {32'h3e2bdf6e, 32'h3f3f581d} /* (5, 31, 4) {real, imag} */,
  {32'h3fe71a97, 32'h3ee16697} /* (5, 31, 3) {real, imag} */,
  {32'h3f36ace0, 32'h3d28e240} /* (5, 31, 2) {real, imag} */,
  {32'h40e4b078, 32'h4056416a} /* (5, 31, 1) {real, imag} */,
  {32'h418da16e, 32'hc09b2d54} /* (5, 31, 0) {real, imag} */,
  {32'h3f37f910, 32'hbf9e8910} /* (5, 30, 31) {real, imag} */,
  {32'hbfe434ce, 32'hc0233f10} /* (5, 30, 30) {real, imag} */,
  {32'hbc8c5e20, 32'hbe53845a} /* (5, 30, 29) {real, imag} */,
  {32'h3e69d564, 32'hbf37755f} /* (5, 30, 28) {real, imag} */,
  {32'h3f57b7b1, 32'h3f8572b9} /* (5, 30, 27) {real, imag} */,
  {32'h3de43a27, 32'hbf0aa4ce} /* (5, 30, 26) {real, imag} */,
  {32'hbe0e2d9e, 32'h3edad9da} /* (5, 30, 25) {real, imag} */,
  {32'h3d3c7780, 32'h3df81028} /* (5, 30, 24) {real, imag} */,
  {32'h3e0d99a5, 32'hbf72d973} /* (5, 30, 23) {real, imag} */,
  {32'hbebba530, 32'hbe2734c4} /* (5, 30, 22) {real, imag} */,
  {32'hbe050fc0, 32'h3e85ed4b} /* (5, 30, 21) {real, imag} */,
  {32'h3d093194, 32'h3df2a765} /* (5, 30, 20) {real, imag} */,
  {32'hbcf721f6, 32'hba16c400} /* (5, 30, 19) {real, imag} */,
  {32'h3a183500, 32'h3e7a9fd2} /* (5, 30, 18) {real, imag} */,
  {32'hbe69b948, 32'hbe3aa6bc} /* (5, 30, 17) {real, imag} */,
  {32'h3e2d36a2, 32'h3df7a9c0} /* (5, 30, 16) {real, imag} */,
  {32'h3e489513, 32'h3e66a7aa} /* (5, 30, 15) {real, imag} */,
  {32'hbd44fca8, 32'h3de3166a} /* (5, 30, 14) {real, imag} */,
  {32'hbe0a04a7, 32'h3ee593ee} /* (5, 30, 13) {real, imag} */,
  {32'h3edc5e12, 32'hbdbbf454} /* (5, 30, 12) {real, imag} */,
  {32'hbe3ca46b, 32'hbe8931f6} /* (5, 30, 11) {real, imag} */,
  {32'h3db22634, 32'h3e5d055c} /* (5, 30, 10) {real, imag} */,
  {32'hbd122184, 32'h3db564d5} /* (5, 30, 9) {real, imag} */,
  {32'h3e8a1216, 32'hbf97f9fd} /* (5, 30, 8) {real, imag} */,
  {32'h3ed844fa, 32'h3e99bcf4} /* (5, 30, 7) {real, imag} */,
  {32'hbf5dc0ea, 32'hbf279de6} /* (5, 30, 6) {real, imag} */,
  {32'hbf7bb23d, 32'hbe1478f8} /* (5, 30, 5) {real, imag} */,
  {32'h3ec8cbb6, 32'h3f203f07} /* (5, 30, 4) {real, imag} */,
  {32'h3c68f2a0, 32'hbf4aec4b} /* (5, 30, 3) {real, imag} */,
  {32'h3f4c8e18, 32'h3ea0cfc0} /* (5, 30, 2) {real, imag} */,
  {32'hbeb3b740, 32'hbd213220} /* (5, 30, 1) {real, imag} */,
  {32'hc014f34e, 32'h3fe141c1} /* (5, 30, 0) {real, imag} */,
  {32'h3ecdc5ec, 32'hbfc72d42} /* (5, 29, 31) {real, imag} */,
  {32'h3f8ccf79, 32'hc00f49d4} /* (5, 29, 30) {real, imag} */,
  {32'hbe9be700, 32'hbeb04cda} /* (5, 29, 29) {real, imag} */,
  {32'h3e99a51e, 32'hbe72991e} /* (5, 29, 28) {real, imag} */,
  {32'hbeb9ce16, 32'h3ea959d8} /* (5, 29, 27) {real, imag} */,
  {32'h3d1133d8, 32'h3f09c1ca} /* (5, 29, 26) {real, imag} */,
  {32'hbea4e860, 32'h3f588e82} /* (5, 29, 25) {real, imag} */,
  {32'hbde75284, 32'hbee8f030} /* (5, 29, 24) {real, imag} */,
  {32'h3c204300, 32'h3e4ade51} /* (5, 29, 23) {real, imag} */,
  {32'h3e38ed07, 32'h3e835e4b} /* (5, 29, 22) {real, imag} */,
  {32'hbee4a6f0, 32'h3f04311a} /* (5, 29, 21) {real, imag} */,
  {32'hbe4aedd3, 32'h3de3fdbc} /* (5, 29, 20) {real, imag} */,
  {32'h3ec5e166, 32'hbe0737b9} /* (5, 29, 19) {real, imag} */,
  {32'h3e727b56, 32'h3ebbdd81} /* (5, 29, 18) {real, imag} */,
  {32'h3ebe8ced, 32'h3dd02368} /* (5, 29, 17) {real, imag} */,
  {32'hbe63e7d6, 32'h3daf8c2e} /* (5, 29, 16) {real, imag} */,
  {32'hbd8b5172, 32'hbe1722b0} /* (5, 29, 15) {real, imag} */,
  {32'hbdcaf1af, 32'h3db22665} /* (5, 29, 14) {real, imag} */,
  {32'h3d4381a2, 32'hbeb2229f} /* (5, 29, 13) {real, imag} */,
  {32'h3f425ffc, 32'h3c24ff00} /* (5, 29, 12) {real, imag} */,
  {32'hbde46820, 32'hbe87ea03} /* (5, 29, 11) {real, imag} */,
  {32'hbdbab9b4, 32'h3e7d48bf} /* (5, 29, 10) {real, imag} */,
  {32'h3eff16f8, 32'h3de6b7cc} /* (5, 29, 9) {real, imag} */,
  {32'h3f32f2b8, 32'h3e00b4a0} /* (5, 29, 8) {real, imag} */,
  {32'hbec8c62a, 32'hbf0575b2} /* (5, 29, 7) {real, imag} */,
  {32'hbf56869f, 32'h3e31d670} /* (5, 29, 6) {real, imag} */,
  {32'hbea280e9, 32'h3f29ae8a} /* (5, 29, 5) {real, imag} */,
  {32'hbec7d1a5, 32'hbde85338} /* (5, 29, 4) {real, imag} */,
  {32'h3d80ca96, 32'hbee5ae72} /* (5, 29, 3) {real, imag} */,
  {32'hbea8df48, 32'h3fa72ee2} /* (5, 29, 2) {real, imag} */,
  {32'h3e666eb8, 32'h3fb21549} /* (5, 29, 1) {real, imag} */,
  {32'h3f00fbc1, 32'hbfd02bfb} /* (5, 29, 0) {real, imag} */,
  {32'hc01bb8b4, 32'hbefeec40} /* (5, 28, 31) {real, imag} */,
  {32'h3f495216, 32'h3ecf0d84} /* (5, 28, 30) {real, imag} */,
  {32'hbf40fcdb, 32'hbf555504} /* (5, 28, 29) {real, imag} */,
  {32'h3f2c6584, 32'h3dd7dc70} /* (5, 28, 28) {real, imag} */,
  {32'h3ea869ff, 32'hbdf8d2e8} /* (5, 28, 27) {real, imag} */,
  {32'hbd7564a8, 32'hbd8440a2} /* (5, 28, 26) {real, imag} */,
  {32'hbf2154e8, 32'h3d9cf48c} /* (5, 28, 25) {real, imag} */,
  {32'h3e4286f5, 32'hbedbdea7} /* (5, 28, 24) {real, imag} */,
  {32'hbf06559a, 32'h3dab3a16} /* (5, 28, 23) {real, imag} */,
  {32'h3e34f5f8, 32'h3f412023} /* (5, 28, 22) {real, imag} */,
  {32'h3eec92c8, 32'hbeb8d52b} /* (5, 28, 21) {real, imag} */,
  {32'hbe77a766, 32'hbedd9f64} /* (5, 28, 20) {real, imag} */,
  {32'hbeffb710, 32'h3e345d8e} /* (5, 28, 19) {real, imag} */,
  {32'h3e9636c0, 32'hbef555e4} /* (5, 28, 18) {real, imag} */,
  {32'hbd122ef4, 32'h3d85d776} /* (5, 28, 17) {real, imag} */,
  {32'hbe35a500, 32'hbe40947a} /* (5, 28, 16) {real, imag} */,
  {32'h3e5093aa, 32'hbd8f0679} /* (5, 28, 15) {real, imag} */,
  {32'hbec59a7d, 32'hbe6c0dc0} /* (5, 28, 14) {real, imag} */,
  {32'hbe8757a0, 32'hbe5a7be6} /* (5, 28, 13) {real, imag} */,
  {32'h3e9c0740, 32'hbf30f3f4} /* (5, 28, 12) {real, imag} */,
  {32'h3e9d3956, 32'h3ec1769a} /* (5, 28, 11) {real, imag} */,
  {32'h3e7c4804, 32'hbde13fb9} /* (5, 28, 10) {real, imag} */,
  {32'h3e1053ae, 32'hbda8cc36} /* (5, 28, 9) {real, imag} */,
  {32'h3f0513a0, 32'h3ebf80f6} /* (5, 28, 8) {real, imag} */,
  {32'h3e033a1c, 32'hbf0ca0ee} /* (5, 28, 7) {real, imag} */,
  {32'hbf33df08, 32'h3ea3a6f8} /* (5, 28, 6) {real, imag} */,
  {32'h3ea3e4e8, 32'h3f39a4fa} /* (5, 28, 5) {real, imag} */,
  {32'h3dcaacb2, 32'hbf038016} /* (5, 28, 4) {real, imag} */,
  {32'h3de3e05d, 32'hbc5388e0} /* (5, 28, 3) {real, imag} */,
  {32'h3e163ce8, 32'hbf4fc354} /* (5, 28, 2) {real, imag} */,
  {32'hbf3dc213, 32'h3f5a51e3} /* (5, 28, 1) {real, imag} */,
  {32'h3eecc939, 32'h3f1148c0} /* (5, 28, 0) {real, imag} */,
  {32'h3f30f85b, 32'hbe42a416} /* (5, 27, 31) {real, imag} */,
  {32'hbdb35e44, 32'hbf28c87a} /* (5, 27, 30) {real, imag} */,
  {32'h3f121aa2, 32'hbd95bdc8} /* (5, 27, 29) {real, imag} */,
  {32'hbf2c5ab0, 32'hbe75a5a7} /* (5, 27, 28) {real, imag} */,
  {32'hbf25ea98, 32'hbe313d60} /* (5, 27, 27) {real, imag} */,
  {32'h3e99459e, 32'h3e76ff96} /* (5, 27, 26) {real, imag} */,
  {32'hbe900a19, 32'h3e1db134} /* (5, 27, 25) {real, imag} */,
  {32'h3e0314cb, 32'hbcb04f04} /* (5, 27, 24) {real, imag} */,
  {32'hbebc02c4, 32'hbdebb5b2} /* (5, 27, 23) {real, imag} */,
  {32'h3d8bf216, 32'hbf0b22d7} /* (5, 27, 22) {real, imag} */,
  {32'h3ea9aed5, 32'h3e643aae} /* (5, 27, 21) {real, imag} */,
  {32'h3de5d141, 32'hbd052890} /* (5, 27, 20) {real, imag} */,
  {32'h3ec3b0f5, 32'hbef2e301} /* (5, 27, 19) {real, imag} */,
  {32'h3e90f440, 32'hbd279ab0} /* (5, 27, 18) {real, imag} */,
  {32'hbe437a24, 32'hbcce99d0} /* (5, 27, 17) {real, imag} */,
  {32'h3dbc5b44, 32'hbd8bc834} /* (5, 27, 16) {real, imag} */,
  {32'hbcf23f26, 32'h3e58b7c0} /* (5, 27, 15) {real, imag} */,
  {32'hbea9bb6a, 32'hbd5c5dd0} /* (5, 27, 14) {real, imag} */,
  {32'hbf17544b, 32'hbea4f7b0} /* (5, 27, 13) {real, imag} */,
  {32'hbe79b317, 32'h3ea42bfc} /* (5, 27, 12) {real, imag} */,
  {32'hbe151511, 32'h3eb50d00} /* (5, 27, 11) {real, imag} */,
  {32'hbf094323, 32'h3f247f57} /* (5, 27, 10) {real, imag} */,
  {32'hbe648fd3, 32'hbef1ab4c} /* (5, 27, 9) {real, imag} */,
  {32'hbf86198c, 32'hbe713ff4} /* (5, 27, 8) {real, imag} */,
  {32'h3e0c633e, 32'hbe3357cb} /* (5, 27, 7) {real, imag} */,
  {32'h3e843aba, 32'hbf1c612a} /* (5, 27, 6) {real, imag} */,
  {32'hbf0e1474, 32'hbf0cc338} /* (5, 27, 5) {real, imag} */,
  {32'hbea55a2d, 32'h3e1cb3a8} /* (5, 27, 4) {real, imag} */,
  {32'hbf2a7356, 32'h3f0ffdd3} /* (5, 27, 3) {real, imag} */,
  {32'hbe97236a, 32'h3e96ccb4} /* (5, 27, 2) {real, imag} */,
  {32'h3f53eb6e, 32'hbfcbbef5} /* (5, 27, 1) {real, imag} */,
  {32'h3ec555c0, 32'hbebd4a1d} /* (5, 27, 0) {real, imag} */,
  {32'hbe47c574, 32'hbe91f4fc} /* (5, 26, 31) {real, imag} */,
  {32'hbf27baa6, 32'h3e947dc7} /* (5, 26, 30) {real, imag} */,
  {32'hbf10c6c7, 32'h3f518a6a} /* (5, 26, 29) {real, imag} */,
  {32'hbdf6ee08, 32'hbe6df240} /* (5, 26, 28) {real, imag} */,
  {32'hbe02b7ec, 32'hbeb3b206} /* (5, 26, 27) {real, imag} */,
  {32'hbee65fb4, 32'hbed859f0} /* (5, 26, 26) {real, imag} */,
  {32'h3f30b280, 32'hbecb180e} /* (5, 26, 25) {real, imag} */,
  {32'hbee656ca, 32'h3e9d9254} /* (5, 26, 24) {real, imag} */,
  {32'h3dbe11b5, 32'h3edb7dc6} /* (5, 26, 23) {real, imag} */,
  {32'h3ef1ac8c, 32'hbdb35291} /* (5, 26, 22) {real, imag} */,
  {32'hbe34b2c8, 32'hbf4a9f41} /* (5, 26, 21) {real, imag} */,
  {32'h3ef76cf8, 32'h3e9fda51} /* (5, 26, 20) {real, imag} */,
  {32'hbceebc44, 32'hbda115cc} /* (5, 26, 19) {real, imag} */,
  {32'h3e9e5949, 32'hbe90a921} /* (5, 26, 18) {real, imag} */,
  {32'hbe35093c, 32'h3c9d8fb0} /* (5, 26, 17) {real, imag} */,
  {32'h3e9d9664, 32'h3e1e84f9} /* (5, 26, 16) {real, imag} */,
  {32'hbec1dec0, 32'h3e673c00} /* (5, 26, 15) {real, imag} */,
  {32'h3e5a7398, 32'hbe3755c4} /* (5, 26, 14) {real, imag} */,
  {32'h3e841f64, 32'hbe6c22ca} /* (5, 26, 13) {real, imag} */,
  {32'hbe351ba0, 32'h3d838da6} /* (5, 26, 12) {real, imag} */,
  {32'hbe928324, 32'h3d122710} /* (5, 26, 11) {real, imag} */,
  {32'hbe410445, 32'hbe9a4a3e} /* (5, 26, 10) {real, imag} */,
  {32'hbeb20f12, 32'hbd83fec0} /* (5, 26, 9) {real, imag} */,
  {32'hbe1a1248, 32'h3e8a33c2} /* (5, 26, 8) {real, imag} */,
  {32'h3d3e8ef0, 32'hbf3f54c4} /* (5, 26, 7) {real, imag} */,
  {32'hbe543026, 32'h3ea28410} /* (5, 26, 6) {real, imag} */,
  {32'h3e9fd09a, 32'hbe9117ca} /* (5, 26, 5) {real, imag} */,
  {32'h3e246f0c, 32'hbdc8b702} /* (5, 26, 4) {real, imag} */,
  {32'h3ed9d75c, 32'h3df818f2} /* (5, 26, 3) {real, imag} */,
  {32'hbed13f72, 32'h3e5dfb50} /* (5, 26, 2) {real, imag} */,
  {32'h3e998fc4, 32'hbf0085d1} /* (5, 26, 1) {real, imag} */,
  {32'h3f5fb55f, 32'hbd99fc88} /* (5, 26, 0) {real, imag} */,
  {32'hbe404a2c, 32'h3e412c74} /* (5, 25, 31) {real, imag} */,
  {32'hbdb6ac94, 32'hbf284746} /* (5, 25, 30) {real, imag} */,
  {32'hbedcdeb8, 32'h3e8c5c02} /* (5, 25, 29) {real, imag} */,
  {32'h3e1e4d49, 32'hbdf467e9} /* (5, 25, 28) {real, imag} */,
  {32'h3e739498, 32'hbf553d65} /* (5, 25, 27) {real, imag} */,
  {32'h3ef19e32, 32'hbe8074f6} /* (5, 25, 26) {real, imag} */,
  {32'hba674b00, 32'h3e471e1a} /* (5, 25, 25) {real, imag} */,
  {32'h3e6ecada, 32'h3e8f0c44} /* (5, 25, 24) {real, imag} */,
  {32'h3eb93cf0, 32'hbe235dd0} /* (5, 25, 23) {real, imag} */,
  {32'h3ee1f372, 32'hbf252934} /* (5, 25, 22) {real, imag} */,
  {32'hbde91222, 32'hbcf65400} /* (5, 25, 21) {real, imag} */,
  {32'hbddb13d8, 32'h3dc6b91b} /* (5, 25, 20) {real, imag} */,
  {32'hbed7c307, 32'hbe289e3a} /* (5, 25, 19) {real, imag} */,
  {32'hbf120707, 32'h3e53b173} /* (5, 25, 18) {real, imag} */,
  {32'hbe88002e, 32'hbeaa0ed7} /* (5, 25, 17) {real, imag} */,
  {32'hb98ca000, 32'h3e7862e6} /* (5, 25, 16) {real, imag} */,
  {32'h3e61d406, 32'hbd4c68ca} /* (5, 25, 15) {real, imag} */,
  {32'h3e46bf23, 32'hbdea803c} /* (5, 25, 14) {real, imag} */,
  {32'hbed5d0e7, 32'hbcfdc1bc} /* (5, 25, 13) {real, imag} */,
  {32'h3f23d00a, 32'h3eb57b93} /* (5, 25, 12) {real, imag} */,
  {32'h3e331f54, 32'hbf24a22c} /* (5, 25, 11) {real, imag} */,
  {32'h3f0c4dce, 32'hbb94a840} /* (5, 25, 10) {real, imag} */,
  {32'hbeb261c1, 32'hbea7cffe} /* (5, 25, 9) {real, imag} */,
  {32'hbeb20a57, 32'hbc8d35c0} /* (5, 25, 8) {real, imag} */,
  {32'h3ed88aaa, 32'h3e9614e8} /* (5, 25, 7) {real, imag} */,
  {32'hbc9f5088, 32'h3d6e2380} /* (5, 25, 6) {real, imag} */,
  {32'hbf14175a, 32'h3db2148b} /* (5, 25, 5) {real, imag} */,
  {32'hbf387f12, 32'h3f29df0d} /* (5, 25, 4) {real, imag} */,
  {32'hbe68f533, 32'h3e0af9b9} /* (5, 25, 3) {real, imag} */,
  {32'hbefd8e0f, 32'h3e9ecef2} /* (5, 25, 2) {real, imag} */,
  {32'h3d4581c8, 32'hbdf0a808} /* (5, 25, 1) {real, imag} */,
  {32'hbf4d6622, 32'h3ebf51a2} /* (5, 25, 0) {real, imag} */,
  {32'hbe912e80, 32'h3e753e30} /* (5, 24, 31) {real, imag} */,
  {32'h3e713ecb, 32'h3e6f1504} /* (5, 24, 30) {real, imag} */,
  {32'hbe344206, 32'h3e1a4529} /* (5, 24, 29) {real, imag} */,
  {32'h3e66258a, 32'h3dcb7efa} /* (5, 24, 28) {real, imag} */,
  {32'hbf35eea0, 32'hbec09eed} /* (5, 24, 27) {real, imag} */,
  {32'h3ed6a992, 32'h3d834150} /* (5, 24, 26) {real, imag} */,
  {32'h3c1451a0, 32'h3f457def} /* (5, 24, 25) {real, imag} */,
  {32'h3f22d6f9, 32'h3f1d4ef0} /* (5, 24, 24) {real, imag} */,
  {32'h3ecb9567, 32'hbf6a13d1} /* (5, 24, 23) {real, imag} */,
  {32'h3e229406, 32'h3d16a530} /* (5, 24, 22) {real, imag} */,
  {32'hbe006a5d, 32'h3dea46d8} /* (5, 24, 21) {real, imag} */,
  {32'hbde032ec, 32'h3e976986} /* (5, 24, 20) {real, imag} */,
  {32'h3e88043d, 32'h3d945a0c} /* (5, 24, 19) {real, imag} */,
  {32'hbf246d56, 32'h3cc38f70} /* (5, 24, 18) {real, imag} */,
  {32'h3e0404e8, 32'hbed579f0} /* (5, 24, 17) {real, imag} */,
  {32'h3d550078, 32'hbb159f00} /* (5, 24, 16) {real, imag} */,
  {32'hbd228ffe, 32'h3e7f0ae5} /* (5, 24, 15) {real, imag} */,
  {32'h3e018228, 32'hbe88c96f} /* (5, 24, 14) {real, imag} */,
  {32'hbdaa7c90, 32'h3c8f4f8c} /* (5, 24, 13) {real, imag} */,
  {32'hbdfd75ec, 32'h3f2ae442} /* (5, 24, 12) {real, imag} */,
  {32'hbe8895d0, 32'h3d3520fc} /* (5, 24, 11) {real, imag} */,
  {32'hbebb29f2, 32'hbd883ea6} /* (5, 24, 10) {real, imag} */,
  {32'h3deed3b4, 32'h3f49870d} /* (5, 24, 9) {real, imag} */,
  {32'hbea19344, 32'hbe8adec8} /* (5, 24, 8) {real, imag} */,
  {32'h3e997b30, 32'hbefcb568} /* (5, 24, 7) {real, imag} */,
  {32'h3ecd5601, 32'hbeb262ae} /* (5, 24, 6) {real, imag} */,
  {32'hbcc70b30, 32'h3e2e78c8} /* (5, 24, 5) {real, imag} */,
  {32'hbef708f6, 32'h3c9ab9f8} /* (5, 24, 4) {real, imag} */,
  {32'h3f9cdcc2, 32'hbf3ae395} /* (5, 24, 3) {real, imag} */,
  {32'hbf04ca1b, 32'hbe7c7f3c} /* (5, 24, 2) {real, imag} */,
  {32'h3f48c834, 32'hbdb78f20} /* (5, 24, 1) {real, imag} */,
  {32'h3f008bc4, 32'h3afda380} /* (5, 24, 0) {real, imag} */,
  {32'hbbe20460, 32'h3dc2bd24} /* (5, 23, 31) {real, imag} */,
  {32'h3dd0b726, 32'h3f4f311e} /* (5, 23, 30) {real, imag} */,
  {32'h3eab8df4, 32'hbf05d461} /* (5, 23, 29) {real, imag} */,
  {32'hbd7f1fc9, 32'h3f06e5ad} /* (5, 23, 28) {real, imag} */,
  {32'hbdef98d2, 32'hbd33b218} /* (5, 23, 27) {real, imag} */,
  {32'hbe7d489a, 32'hbdbb11f4} /* (5, 23, 26) {real, imag} */,
  {32'h3eb9749e, 32'h3e2621b5} /* (5, 23, 25) {real, imag} */,
  {32'h3efd1c13, 32'hbde0c50e} /* (5, 23, 24) {real, imag} */,
  {32'h3e209265, 32'h3c5ebbe0} /* (5, 23, 23) {real, imag} */,
  {32'hbcc5e3f0, 32'hbe56f1f7} /* (5, 23, 22) {real, imag} */,
  {32'hbd040fa8, 32'hbd935475} /* (5, 23, 21) {real, imag} */,
  {32'hbd64dd5a, 32'h3cc7e6b4} /* (5, 23, 20) {real, imag} */,
  {32'h3ed69261, 32'hbea596f1} /* (5, 23, 19) {real, imag} */,
  {32'hbda6930c, 32'h3d842717} /* (5, 23, 18) {real, imag} */,
  {32'hbed15fac, 32'hbd9f29bd} /* (5, 23, 17) {real, imag} */,
  {32'h3eb4b578, 32'hbd3bcba4} /* (5, 23, 16) {real, imag} */,
  {32'hbeba543b, 32'hbef82337} /* (5, 23, 15) {real, imag} */,
  {32'hbe0a96b0, 32'hbcc13bb0} /* (5, 23, 14) {real, imag} */,
  {32'hbd88a902, 32'hbdff1d1e} /* (5, 23, 13) {real, imag} */,
  {32'hbe9d05cb, 32'hbf2c9d6f} /* (5, 23, 12) {real, imag} */,
  {32'h3e75fd1e, 32'h3f4b0d00} /* (5, 23, 11) {real, imag} */,
  {32'h3ee0129a, 32'hbf303b75} /* (5, 23, 10) {real, imag} */,
  {32'hbe9510a3, 32'hbea0a68c} /* (5, 23, 9) {real, imag} */,
  {32'h3ea00395, 32'h3f15590e} /* (5, 23, 8) {real, imag} */,
  {32'h3e83f7d9, 32'h3d0a971e} /* (5, 23, 7) {real, imag} */,
  {32'h3e8ca1db, 32'hbe4be539} /* (5, 23, 6) {real, imag} */,
  {32'h3ea1adaa, 32'hbdc6052e} /* (5, 23, 5) {real, imag} */,
  {32'hbc8d0ef0, 32'hbd8a337b} /* (5, 23, 4) {real, imag} */,
  {32'hbe4f04b8, 32'hbdda12e7} /* (5, 23, 3) {real, imag} */,
  {32'h3eecaea1, 32'hbdbb0e50} /* (5, 23, 2) {real, imag} */,
  {32'h3c7e92c0, 32'h3ecba3d6} /* (5, 23, 1) {real, imag} */,
  {32'hbf4b01aa, 32'hbe699c2b} /* (5, 23, 0) {real, imag} */,
  {32'hbe0dabc1, 32'hbdd74f13} /* (5, 22, 31) {real, imag} */,
  {32'hbd3fcfc0, 32'h3ba808c0} /* (5, 22, 30) {real, imag} */,
  {32'hbe40d714, 32'h3ee7400a} /* (5, 22, 29) {real, imag} */,
  {32'h3e76b8ec, 32'h3ed12cfb} /* (5, 22, 28) {real, imag} */,
  {32'hbe94e008, 32'hbd53c355} /* (5, 22, 27) {real, imag} */,
  {32'hbe38f7ae, 32'hbe54b468} /* (5, 22, 26) {real, imag} */,
  {32'h3efa40ef, 32'hbf6912dc} /* (5, 22, 25) {real, imag} */,
  {32'h3ea0c52b, 32'h3db5ad86} /* (5, 22, 24) {real, imag} */,
  {32'hbeb58b81, 32'hbe51b6d8} /* (5, 22, 23) {real, imag} */,
  {32'hbe73928f, 32'hbe2b51c0} /* (5, 22, 22) {real, imag} */,
  {32'hbea71ce0, 32'hbe7cc2e8} /* (5, 22, 21) {real, imag} */,
  {32'hbe29ffeb, 32'h3f030938} /* (5, 22, 20) {real, imag} */,
  {32'h3e8bdff8, 32'h3d064b18} /* (5, 22, 19) {real, imag} */,
  {32'hbddf35bf, 32'h3ea103e9} /* (5, 22, 18) {real, imag} */,
  {32'h3ef5f945, 32'hbd810e84} /* (5, 22, 17) {real, imag} */,
  {32'h3df3b228, 32'h3ee704f8} /* (5, 22, 16) {real, imag} */,
  {32'h3e4c5d40, 32'h3df6f8e0} /* (5, 22, 15) {real, imag} */,
  {32'h3ec9bc5b, 32'h3cf7b5a0} /* (5, 22, 14) {real, imag} */,
  {32'h3eb24e00, 32'h3e95c321} /* (5, 22, 13) {real, imag} */,
  {32'hbe05de3c, 32'hbd0b5d20} /* (5, 22, 12) {real, imag} */,
  {32'hbef37412, 32'h3ef363c6} /* (5, 22, 11) {real, imag} */,
  {32'h3ea216bb, 32'hbd2e9bd0} /* (5, 22, 10) {real, imag} */,
  {32'h3b82ad60, 32'hbdcb63d0} /* (5, 22, 9) {real, imag} */,
  {32'hbef940ab, 32'h3dc93e24} /* (5, 22, 8) {real, imag} */,
  {32'h3ef63b46, 32'hbced8c98} /* (5, 22, 7) {real, imag} */,
  {32'hbd6a1660, 32'hbf40d422} /* (5, 22, 6) {real, imag} */,
  {32'h3f245438, 32'hbed35840} /* (5, 22, 5) {real, imag} */,
  {32'hbe665807, 32'h3ef34f98} /* (5, 22, 4) {real, imag} */,
  {32'hbf08572e, 32'h3c8c3ef0} /* (5, 22, 3) {real, imag} */,
  {32'hbd8228fa, 32'h3ecf340e} /* (5, 22, 2) {real, imag} */,
  {32'h3bc85d00, 32'h3f204356} /* (5, 22, 1) {real, imag} */,
  {32'hbd981a96, 32'h3dfa0e62} /* (5, 22, 0) {real, imag} */,
  {32'h3cf3e850, 32'h3dd2a51c} /* (5, 21, 31) {real, imag} */,
  {32'h3df263ba, 32'h3de5f150} /* (5, 21, 30) {real, imag} */,
  {32'h3eb85ce4, 32'h3ece1650} /* (5, 21, 29) {real, imag} */,
  {32'h3df15e5c, 32'hbe25fda6} /* (5, 21, 28) {real, imag} */,
  {32'hbdeb6e30, 32'hbba03940} /* (5, 21, 27) {real, imag} */,
  {32'hbf1d2e01, 32'hbec4937d} /* (5, 21, 26) {real, imag} */,
  {32'hbf0ab3bc, 32'hbe3726a1} /* (5, 21, 25) {real, imag} */,
  {32'h3e913596, 32'h3f19388d} /* (5, 21, 24) {real, imag} */,
  {32'h3e993f90, 32'hbe7cb2aa} /* (5, 21, 23) {real, imag} */,
  {32'hbf419235, 32'h3ece4880} /* (5, 21, 22) {real, imag} */,
  {32'h3f8669de, 32'h3e891faf} /* (5, 21, 21) {real, imag} */,
  {32'hbc98dfa8, 32'h3e5b7208} /* (5, 21, 20) {real, imag} */,
  {32'hbd2fb4f0, 32'hbd51925c} /* (5, 21, 19) {real, imag} */,
  {32'h3e792761, 32'h3d3b1e6e} /* (5, 21, 18) {real, imag} */,
  {32'hbea8055f, 32'h3ec1d208} /* (5, 21, 17) {real, imag} */,
  {32'h3e41cf64, 32'hbef80adc} /* (5, 21, 16) {real, imag} */,
  {32'h3dcdca04, 32'h3e970c31} /* (5, 21, 15) {real, imag} */,
  {32'h3d2fe550, 32'hbe4281dc} /* (5, 21, 14) {real, imag} */,
  {32'h3e855f9e, 32'hbf3682dc} /* (5, 21, 13) {real, imag} */,
  {32'h3d09294c, 32'hbed68298} /* (5, 21, 12) {real, imag} */,
  {32'hbf2391b8, 32'hbe36cba8} /* (5, 21, 11) {real, imag} */,
  {32'h3d9ea37f, 32'h3f3e2b62} /* (5, 21, 10) {real, imag} */,
  {32'h3e8ddaa7, 32'h3b80a580} /* (5, 21, 9) {real, imag} */,
  {32'h3d3649ec, 32'hbc5250f4} /* (5, 21, 8) {real, imag} */,
  {32'hbe2f601e, 32'hbe5ae229} /* (5, 21, 7) {real, imag} */,
  {32'h3d3a3cbe, 32'h3dbb1007} /* (5, 21, 6) {real, imag} */,
  {32'h3d35225d, 32'hbe707d85} /* (5, 21, 5) {real, imag} */,
  {32'h3ea660cc, 32'hbe93e792} /* (5, 21, 4) {real, imag} */,
  {32'hbebd9c4a, 32'hbe0808ea} /* (5, 21, 3) {real, imag} */,
  {32'h3e83f4c8, 32'hbe80b28b} /* (5, 21, 2) {real, imag} */,
  {32'h3e8452f9, 32'hbd34856c} /* (5, 21, 1) {real, imag} */,
  {32'h3ec28fa2, 32'hbe02283a} /* (5, 21, 0) {real, imag} */,
  {32'hbe3c0c8a, 32'hbf0dc2fd} /* (5, 20, 31) {real, imag} */,
  {32'hbd2e3164, 32'hbdcbf450} /* (5, 20, 30) {real, imag} */,
  {32'h3e24241b, 32'h3e73a5c4} /* (5, 20, 29) {real, imag} */,
  {32'hbed0da8d, 32'hbdd081b4} /* (5, 20, 28) {real, imag} */,
  {32'h3ea23ef4, 32'h3db76ea4} /* (5, 20, 27) {real, imag} */,
  {32'hbe04ab83, 32'h3e37d11e} /* (5, 20, 26) {real, imag} */,
  {32'hbe1055fc, 32'hbea36c39} /* (5, 20, 25) {real, imag} */,
  {32'hbf0c6683, 32'h3d02331a} /* (5, 20, 24) {real, imag} */,
  {32'h3f21872b, 32'h3eb57864} /* (5, 20, 23) {real, imag} */,
  {32'hbeb1f893, 32'h3efd427d} /* (5, 20, 22) {real, imag} */,
  {32'hbec6574e, 32'hbe310006} /* (5, 20, 21) {real, imag} */,
  {32'hbdd093c2, 32'hbdbc14c6} /* (5, 20, 20) {real, imag} */,
  {32'hbe625e4f, 32'h3b22cae0} /* (5, 20, 19) {real, imag} */,
  {32'h3e348476, 32'h3f7b357e} /* (5, 20, 18) {real, imag} */,
  {32'h3edc9a3b, 32'h3e401e7c} /* (5, 20, 17) {real, imag} */,
  {32'hbba02378, 32'hbd0ee302} /* (5, 20, 16) {real, imag} */,
  {32'hbe169107, 32'hbe3abffc} /* (5, 20, 15) {real, imag} */,
  {32'hbf26a305, 32'h3e8552b2} /* (5, 20, 14) {real, imag} */,
  {32'h3da180c9, 32'h3ca5d5e8} /* (5, 20, 13) {real, imag} */,
  {32'h3f00e988, 32'hbeb16ad8} /* (5, 20, 12) {real, imag} */,
  {32'h3d86d1f0, 32'h3c9fd600} /* (5, 20, 11) {real, imag} */,
  {32'h3d87c3dc, 32'hbd1b2e48} /* (5, 20, 10) {real, imag} */,
  {32'h3dd04df8, 32'hbb865ec0} /* (5, 20, 9) {real, imag} */,
  {32'h3de3e5ac, 32'h3e6a61aa} /* (5, 20, 8) {real, imag} */,
  {32'h3f143038, 32'h3ea9a46f} /* (5, 20, 7) {real, imag} */,
  {32'hbefa2a50, 32'h3eef3b9b} /* (5, 20, 6) {real, imag} */,
  {32'h3e29bbd0, 32'hbe8f5b2e} /* (5, 20, 5) {real, imag} */,
  {32'h3dc40aae, 32'h3e83d723} /* (5, 20, 4) {real, imag} */,
  {32'h3eb0e622, 32'h3e269f62} /* (5, 20, 3) {real, imag} */,
  {32'hbeba82db, 32'hbdd01010} /* (5, 20, 2) {real, imag} */,
  {32'h3e810ec2, 32'hbdd5e8ff} /* (5, 20, 1) {real, imag} */,
  {32'hbdb6b83b, 32'h3e0de54f} /* (5, 20, 0) {real, imag} */,
  {32'h3eb9855c, 32'hbdf9b093} /* (5, 19, 31) {real, imag} */,
  {32'h3f18f6e2, 32'h3dca2038} /* (5, 19, 30) {real, imag} */,
  {32'hbcc78968, 32'hbe15b681} /* (5, 19, 29) {real, imag} */,
  {32'hbda865aa, 32'h3dc5e060} /* (5, 19, 28) {real, imag} */,
  {32'hbd542d0c, 32'hbda37863} /* (5, 19, 27) {real, imag} */,
  {32'h3e7d2ebd, 32'hbcb1f160} /* (5, 19, 26) {real, imag} */,
  {32'hbf81b858, 32'h3e4288e3} /* (5, 19, 25) {real, imag} */,
  {32'hbe0e4869, 32'hbe131f24} /* (5, 19, 24) {real, imag} */,
  {32'hbe8deca8, 32'h3f373d28} /* (5, 19, 23) {real, imag} */,
  {32'hbe78ace0, 32'hbd85cb6f} /* (5, 19, 22) {real, imag} */,
  {32'h3e0a3995, 32'hbdd72415} /* (5, 19, 21) {real, imag} */,
  {32'h3d01dcf0, 32'hbe68e627} /* (5, 19, 20) {real, imag} */,
  {32'h3f1b2ba8, 32'h3c0d2b00} /* (5, 19, 19) {real, imag} */,
  {32'hbe88b50a, 32'hbe2e82b3} /* (5, 19, 18) {real, imag} */,
  {32'hbc3fba30, 32'hba8361c0} /* (5, 19, 17) {real, imag} */,
  {32'hbf07f109, 32'hbe3a3a99} /* (5, 19, 16) {real, imag} */,
  {32'hbf100920, 32'hbda7b89e} /* (5, 19, 15) {real, imag} */,
  {32'h3d2a9c4c, 32'hbeb164bf} /* (5, 19, 14) {real, imag} */,
  {32'hbe80feaf, 32'h3e952e21} /* (5, 19, 13) {real, imag} */,
  {32'h3f0084d0, 32'h3e451996} /* (5, 19, 12) {real, imag} */,
  {32'h3e7c8d94, 32'h3ee07f4a} /* (5, 19, 11) {real, imag} */,
  {32'h3eb3c7ad, 32'hbedab884} /* (5, 19, 10) {real, imag} */,
  {32'hbf19aeab, 32'h3e8a5c4e} /* (5, 19, 9) {real, imag} */,
  {32'h3e7316e3, 32'h3e6bebea} /* (5, 19, 8) {real, imag} */,
  {32'hbd29b7ac, 32'h3eed1c26} /* (5, 19, 7) {real, imag} */,
  {32'hbe80aafb, 32'h3deafedf} /* (5, 19, 6) {real, imag} */,
  {32'hbe6bf916, 32'hbd2e7a75} /* (5, 19, 5) {real, imag} */,
  {32'hbe3553f5, 32'hbe702624} /* (5, 19, 4) {real, imag} */,
  {32'hbe25f7a8, 32'h3d7eb500} /* (5, 19, 3) {real, imag} */,
  {32'h3ecfebe8, 32'hbec3690e} /* (5, 19, 2) {real, imag} */,
  {32'hbecc137a, 32'h3e2495e0} /* (5, 19, 1) {real, imag} */,
  {32'hbdef7c10, 32'h3e8885ee} /* (5, 19, 0) {real, imag} */,
  {32'hbe45f160, 32'hbce0ee68} /* (5, 18, 31) {real, imag} */,
  {32'h3ecac6fb, 32'h3d89f858} /* (5, 18, 30) {real, imag} */,
  {32'hbe827a36, 32'h3e3aa91e} /* (5, 18, 29) {real, imag} */,
  {32'hbf0953d5, 32'hbe2ca796} /* (5, 18, 28) {real, imag} */,
  {32'h3e33dbc6, 32'hbeab6ecb} /* (5, 18, 27) {real, imag} */,
  {32'h3d34f0e2, 32'hbea25b9a} /* (5, 18, 26) {real, imag} */,
  {32'hbd027480, 32'hbe99c425} /* (5, 18, 25) {real, imag} */,
  {32'h3ef56960, 32'h3eb92c5e} /* (5, 18, 24) {real, imag} */,
  {32'h3de26e82, 32'hbdf5728e} /* (5, 18, 23) {real, imag} */,
  {32'hbe8ff64f, 32'hbe8ee591} /* (5, 18, 22) {real, imag} */,
  {32'h3e9322d0, 32'h3ddf69ed} /* (5, 18, 21) {real, imag} */,
  {32'hbe307fd2, 32'hbe5718bc} /* (5, 18, 20) {real, imag} */,
  {32'h3edcf6aa, 32'h3dde1e5b} /* (5, 18, 19) {real, imag} */,
  {32'hbdd5a78c, 32'h3d26bde0} /* (5, 18, 18) {real, imag} */,
  {32'h3e9d2856, 32'hbc792c80} /* (5, 18, 17) {real, imag} */,
  {32'h3d597eb6, 32'h3e6931e8} /* (5, 18, 16) {real, imag} */,
  {32'hbe8e125b, 32'hbda242f0} /* (5, 18, 15) {real, imag} */,
  {32'h3d1f72a0, 32'hbd04ba49} /* (5, 18, 14) {real, imag} */,
  {32'h3e142203, 32'h3e0c05ea} /* (5, 18, 13) {real, imag} */,
  {32'hbf4014d6, 32'h3f0917a9} /* (5, 18, 12) {real, imag} */,
  {32'h3ed794c4, 32'h3e9a96ee} /* (5, 18, 11) {real, imag} */,
  {32'h3df8a6e0, 32'h3dd893e8} /* (5, 18, 10) {real, imag} */,
  {32'h3e131115, 32'h3be75f60} /* (5, 18, 9) {real, imag} */,
  {32'hbeaab1bd, 32'h3d84f46e} /* (5, 18, 8) {real, imag} */,
  {32'hbe3ba65c, 32'h3eb9c137} /* (5, 18, 7) {real, imag} */,
  {32'hbe2b839e, 32'hbf437dd4} /* (5, 18, 6) {real, imag} */,
  {32'hbcbf6192, 32'hbe5d055b} /* (5, 18, 5) {real, imag} */,
  {32'hbd57b380, 32'h3d00d494} /* (5, 18, 4) {real, imag} */,
  {32'h3d612bb2, 32'hbe34571c} /* (5, 18, 3) {real, imag} */,
  {32'hbbf5afc0, 32'h3eb3d49e} /* (5, 18, 2) {real, imag} */,
  {32'hbde9ea98, 32'hbd3b6d14} /* (5, 18, 1) {real, imag} */,
  {32'h3e78027d, 32'hbdf89667} /* (5, 18, 0) {real, imag} */,
  {32'h3e60fedc, 32'hbdcfbb1a} /* (5, 17, 31) {real, imag} */,
  {32'hbd209aec, 32'hbdbb95c4} /* (5, 17, 30) {real, imag} */,
  {32'h3e2740f3, 32'h3e72522c} /* (5, 17, 29) {real, imag} */,
  {32'h3b5cd830, 32'h3dfec538} /* (5, 17, 28) {real, imag} */,
  {32'hbe75fa7e, 32'h3d8d809e} /* (5, 17, 27) {real, imag} */,
  {32'h3d2ccb6a, 32'h3e9a91b3} /* (5, 17, 26) {real, imag} */,
  {32'hbe6359f1, 32'hbdda3ab8} /* (5, 17, 25) {real, imag} */,
  {32'hbe80b9b4, 32'h3d8c1a7f} /* (5, 17, 24) {real, imag} */,
  {32'hbeeafb42, 32'hbd401b70} /* (5, 17, 23) {real, imag} */,
  {32'h3ce9b578, 32'h3e07e303} /* (5, 17, 22) {real, imag} */,
  {32'hbeee822e, 32'hbda8a9a0} /* (5, 17, 21) {real, imag} */,
  {32'h3e7e2638, 32'hbcf1a7bc} /* (5, 17, 20) {real, imag} */,
  {32'hbeb00d40, 32'hbeb65ca3} /* (5, 17, 19) {real, imag} */,
  {32'h3e4ff076, 32'h3da10e90} /* (5, 17, 18) {real, imag} */,
  {32'hbe1de6c6, 32'hbc6cb940} /* (5, 17, 17) {real, imag} */,
  {32'h3ed395fc, 32'h3e017a56} /* (5, 17, 16) {real, imag} */,
  {32'h3b5e14e0, 32'hbea0a528} /* (5, 17, 15) {real, imag} */,
  {32'hbdbc3826, 32'h3e1e534a} /* (5, 17, 14) {real, imag} */,
  {32'hbdd90254, 32'h3ecc16ee} /* (5, 17, 13) {real, imag} */,
  {32'hbe93ce23, 32'hbf205cec} /* (5, 17, 12) {real, imag} */,
  {32'h3eb9af98, 32'hbe5d49a3} /* (5, 17, 11) {real, imag} */,
  {32'hbd76f309, 32'h3e3f0b98} /* (5, 17, 10) {real, imag} */,
  {32'hbe40ded7, 32'h3eb3d3ce} /* (5, 17, 9) {real, imag} */,
  {32'hbd835b20, 32'hbdaf2b16} /* (5, 17, 8) {real, imag} */,
  {32'hbe1a46af, 32'hbc5d8c3c} /* (5, 17, 7) {real, imag} */,
  {32'h3e2624ff, 32'h3eaf5ee6} /* (5, 17, 6) {real, imag} */,
  {32'hbe66afe8, 32'hbca4b638} /* (5, 17, 5) {real, imag} */,
  {32'h3e55378b, 32'hbea122ec} /* (5, 17, 4) {real, imag} */,
  {32'h3db52118, 32'hbe13a120} /* (5, 17, 3) {real, imag} */,
  {32'h3dc17a50, 32'hbdb62afa} /* (5, 17, 2) {real, imag} */,
  {32'hbe169fa5, 32'h3f46d50c} /* (5, 17, 1) {real, imag} */,
  {32'h3e2a6297, 32'h3ea828a1} /* (5, 17, 0) {real, imag} */,
  {32'h3db41599, 32'hbc207780} /* (5, 16, 31) {real, imag} */,
  {32'h3c80112c, 32'h3e172c8e} /* (5, 16, 30) {real, imag} */,
  {32'h3e1829ee, 32'h3e25ef6e} /* (5, 16, 29) {real, imag} */,
  {32'hbe7a71f0, 32'h3c73ffa0} /* (5, 16, 28) {real, imag} */,
  {32'h3df1b6f1, 32'hbe981466} /* (5, 16, 27) {real, imag} */,
  {32'hbec4b57c, 32'h3dbee64f} /* (5, 16, 26) {real, imag} */,
  {32'hbd99108e, 32'hbd767f28} /* (5, 16, 25) {real, imag} */,
  {32'hbde375d6, 32'hbc395448} /* (5, 16, 24) {real, imag} */,
  {32'hbcb23e72, 32'hbe6505a2} /* (5, 16, 23) {real, imag} */,
  {32'hbe52b9ea, 32'h3d502c79} /* (5, 16, 22) {real, imag} */,
  {32'h3e579aea, 32'h3e82946c} /* (5, 16, 21) {real, imag} */,
  {32'h3ea38c95, 32'hbd729e50} /* (5, 16, 20) {real, imag} */,
  {32'h3e9bc8a7, 32'h3ee9cb23} /* (5, 16, 19) {real, imag} */,
  {32'hbe04d942, 32'hbd667c24} /* (5, 16, 18) {real, imag} */,
  {32'h3b296dc0, 32'hbe3d5427} /* (5, 16, 17) {real, imag} */,
  {32'hbdd62ad7, 32'h00000000} /* (5, 16, 16) {real, imag} */,
  {32'h3b296dc0, 32'h3e3d5427} /* (5, 16, 15) {real, imag} */,
  {32'hbe04d942, 32'h3d667c24} /* (5, 16, 14) {real, imag} */,
  {32'h3e9bc8a7, 32'hbee9cb23} /* (5, 16, 13) {real, imag} */,
  {32'h3ea38c95, 32'h3d729e50} /* (5, 16, 12) {real, imag} */,
  {32'h3e579aea, 32'hbe82946c} /* (5, 16, 11) {real, imag} */,
  {32'hbe52b9ea, 32'hbd502c79} /* (5, 16, 10) {real, imag} */,
  {32'hbcb23e72, 32'h3e6505a2} /* (5, 16, 9) {real, imag} */,
  {32'hbde375d6, 32'h3c395448} /* (5, 16, 8) {real, imag} */,
  {32'hbd99108e, 32'h3d767f28} /* (5, 16, 7) {real, imag} */,
  {32'hbec4b57c, 32'hbdbee64f} /* (5, 16, 6) {real, imag} */,
  {32'h3df1b6f1, 32'h3e981466} /* (5, 16, 5) {real, imag} */,
  {32'hbe7a71f0, 32'hbc73ffa0} /* (5, 16, 4) {real, imag} */,
  {32'h3e1829ee, 32'hbe25ef6e} /* (5, 16, 3) {real, imag} */,
  {32'h3c80112c, 32'hbe172c8e} /* (5, 16, 2) {real, imag} */,
  {32'h3db41599, 32'h3c207780} /* (5, 16, 1) {real, imag} */,
  {32'h3ec8d2a7, 32'h00000000} /* (5, 16, 0) {real, imag} */,
  {32'hbe169fa5, 32'hbf46d50c} /* (5, 15, 31) {real, imag} */,
  {32'h3dc17a50, 32'h3db62afa} /* (5, 15, 30) {real, imag} */,
  {32'h3db52118, 32'h3e13a120} /* (5, 15, 29) {real, imag} */,
  {32'h3e55378b, 32'h3ea122ec} /* (5, 15, 28) {real, imag} */,
  {32'hbe66afe8, 32'h3ca4b638} /* (5, 15, 27) {real, imag} */,
  {32'h3e2624ff, 32'hbeaf5ee6} /* (5, 15, 26) {real, imag} */,
  {32'hbe1a46af, 32'h3c5d8c3c} /* (5, 15, 25) {real, imag} */,
  {32'hbd835b20, 32'h3daf2b16} /* (5, 15, 24) {real, imag} */,
  {32'hbe40ded7, 32'hbeb3d3ce} /* (5, 15, 23) {real, imag} */,
  {32'hbd76f309, 32'hbe3f0b98} /* (5, 15, 22) {real, imag} */,
  {32'h3eb9af98, 32'h3e5d49a3} /* (5, 15, 21) {real, imag} */,
  {32'hbe93ce23, 32'h3f205cec} /* (5, 15, 20) {real, imag} */,
  {32'hbdd90254, 32'hbecc16ee} /* (5, 15, 19) {real, imag} */,
  {32'hbdbc3826, 32'hbe1e534a} /* (5, 15, 18) {real, imag} */,
  {32'h3b5e14e0, 32'h3ea0a528} /* (5, 15, 17) {real, imag} */,
  {32'h3ed395fc, 32'hbe017a56} /* (5, 15, 16) {real, imag} */,
  {32'hbe1de6c6, 32'h3c6cb940} /* (5, 15, 15) {real, imag} */,
  {32'h3e4ff076, 32'hbda10e90} /* (5, 15, 14) {real, imag} */,
  {32'hbeb00d40, 32'h3eb65ca3} /* (5, 15, 13) {real, imag} */,
  {32'h3e7e2638, 32'h3cf1a7bc} /* (5, 15, 12) {real, imag} */,
  {32'hbeee822e, 32'h3da8a9a0} /* (5, 15, 11) {real, imag} */,
  {32'h3ce9b578, 32'hbe07e303} /* (5, 15, 10) {real, imag} */,
  {32'hbeeafb42, 32'h3d401b70} /* (5, 15, 9) {real, imag} */,
  {32'hbe80b9b4, 32'hbd8c1a7f} /* (5, 15, 8) {real, imag} */,
  {32'hbe6359f1, 32'h3dda3ab8} /* (5, 15, 7) {real, imag} */,
  {32'h3d2ccb6a, 32'hbe9a91b3} /* (5, 15, 6) {real, imag} */,
  {32'hbe75fa7e, 32'hbd8d809e} /* (5, 15, 5) {real, imag} */,
  {32'h3b5cd830, 32'hbdfec538} /* (5, 15, 4) {real, imag} */,
  {32'h3e2740f3, 32'hbe72522c} /* (5, 15, 3) {real, imag} */,
  {32'hbd209aec, 32'h3dbb95c4} /* (5, 15, 2) {real, imag} */,
  {32'h3e60fedc, 32'h3dcfbb1a} /* (5, 15, 1) {real, imag} */,
  {32'h3e2a6297, 32'hbea828a1} /* (5, 15, 0) {real, imag} */,
  {32'hbde9ea98, 32'h3d3b6d14} /* (5, 14, 31) {real, imag} */,
  {32'hbbf5afc0, 32'hbeb3d49e} /* (5, 14, 30) {real, imag} */,
  {32'h3d612bb2, 32'h3e34571c} /* (5, 14, 29) {real, imag} */,
  {32'hbd57b380, 32'hbd00d494} /* (5, 14, 28) {real, imag} */,
  {32'hbcbf6192, 32'h3e5d055b} /* (5, 14, 27) {real, imag} */,
  {32'hbe2b839e, 32'h3f437dd4} /* (5, 14, 26) {real, imag} */,
  {32'hbe3ba65c, 32'hbeb9c137} /* (5, 14, 25) {real, imag} */,
  {32'hbeaab1bd, 32'hbd84f46e} /* (5, 14, 24) {real, imag} */,
  {32'h3e131115, 32'hbbe75f60} /* (5, 14, 23) {real, imag} */,
  {32'h3df8a6e0, 32'hbdd893e8} /* (5, 14, 22) {real, imag} */,
  {32'h3ed794c4, 32'hbe9a96ee} /* (5, 14, 21) {real, imag} */,
  {32'hbf4014d6, 32'hbf0917a9} /* (5, 14, 20) {real, imag} */,
  {32'h3e142203, 32'hbe0c05ea} /* (5, 14, 19) {real, imag} */,
  {32'h3d1f72a0, 32'h3d04ba49} /* (5, 14, 18) {real, imag} */,
  {32'hbe8e125b, 32'h3da242f0} /* (5, 14, 17) {real, imag} */,
  {32'h3d597eb6, 32'hbe6931e8} /* (5, 14, 16) {real, imag} */,
  {32'h3e9d2856, 32'h3c792c80} /* (5, 14, 15) {real, imag} */,
  {32'hbdd5a78c, 32'hbd26bde0} /* (5, 14, 14) {real, imag} */,
  {32'h3edcf6aa, 32'hbdde1e5b} /* (5, 14, 13) {real, imag} */,
  {32'hbe307fd2, 32'h3e5718bc} /* (5, 14, 12) {real, imag} */,
  {32'h3e9322d0, 32'hbddf69ed} /* (5, 14, 11) {real, imag} */,
  {32'hbe8ff64f, 32'h3e8ee591} /* (5, 14, 10) {real, imag} */,
  {32'h3de26e82, 32'h3df5728e} /* (5, 14, 9) {real, imag} */,
  {32'h3ef56960, 32'hbeb92c5e} /* (5, 14, 8) {real, imag} */,
  {32'hbd027480, 32'h3e99c425} /* (5, 14, 7) {real, imag} */,
  {32'h3d34f0e2, 32'h3ea25b9a} /* (5, 14, 6) {real, imag} */,
  {32'h3e33dbc6, 32'h3eab6ecb} /* (5, 14, 5) {real, imag} */,
  {32'hbf0953d5, 32'h3e2ca796} /* (5, 14, 4) {real, imag} */,
  {32'hbe827a36, 32'hbe3aa91e} /* (5, 14, 3) {real, imag} */,
  {32'h3ecac6fb, 32'hbd89f858} /* (5, 14, 2) {real, imag} */,
  {32'hbe45f160, 32'h3ce0ee68} /* (5, 14, 1) {real, imag} */,
  {32'h3e78027d, 32'h3df89667} /* (5, 14, 0) {real, imag} */,
  {32'hbecc137a, 32'hbe2495e0} /* (5, 13, 31) {real, imag} */,
  {32'h3ecfebe8, 32'h3ec3690e} /* (5, 13, 30) {real, imag} */,
  {32'hbe25f7a8, 32'hbd7eb500} /* (5, 13, 29) {real, imag} */,
  {32'hbe3553f5, 32'h3e702624} /* (5, 13, 28) {real, imag} */,
  {32'hbe6bf916, 32'h3d2e7a75} /* (5, 13, 27) {real, imag} */,
  {32'hbe80aafb, 32'hbdeafedf} /* (5, 13, 26) {real, imag} */,
  {32'hbd29b7ac, 32'hbeed1c26} /* (5, 13, 25) {real, imag} */,
  {32'h3e7316e3, 32'hbe6bebea} /* (5, 13, 24) {real, imag} */,
  {32'hbf19aeab, 32'hbe8a5c4e} /* (5, 13, 23) {real, imag} */,
  {32'h3eb3c7ad, 32'h3edab884} /* (5, 13, 22) {real, imag} */,
  {32'h3e7c8d94, 32'hbee07f4a} /* (5, 13, 21) {real, imag} */,
  {32'h3f0084d0, 32'hbe451996} /* (5, 13, 20) {real, imag} */,
  {32'hbe80feaf, 32'hbe952e21} /* (5, 13, 19) {real, imag} */,
  {32'h3d2a9c4c, 32'h3eb164bf} /* (5, 13, 18) {real, imag} */,
  {32'hbf100920, 32'h3da7b89e} /* (5, 13, 17) {real, imag} */,
  {32'hbf07f109, 32'h3e3a3a99} /* (5, 13, 16) {real, imag} */,
  {32'hbc3fba30, 32'h3a8361c0} /* (5, 13, 15) {real, imag} */,
  {32'hbe88b50a, 32'h3e2e82b3} /* (5, 13, 14) {real, imag} */,
  {32'h3f1b2ba8, 32'hbc0d2b00} /* (5, 13, 13) {real, imag} */,
  {32'h3d01dcf0, 32'h3e68e627} /* (5, 13, 12) {real, imag} */,
  {32'h3e0a3995, 32'h3dd72415} /* (5, 13, 11) {real, imag} */,
  {32'hbe78ace0, 32'h3d85cb6f} /* (5, 13, 10) {real, imag} */,
  {32'hbe8deca8, 32'hbf373d28} /* (5, 13, 9) {real, imag} */,
  {32'hbe0e4869, 32'h3e131f24} /* (5, 13, 8) {real, imag} */,
  {32'hbf81b858, 32'hbe4288e3} /* (5, 13, 7) {real, imag} */,
  {32'h3e7d2ebd, 32'h3cb1f160} /* (5, 13, 6) {real, imag} */,
  {32'hbd542d0c, 32'h3da37863} /* (5, 13, 5) {real, imag} */,
  {32'hbda865aa, 32'hbdc5e060} /* (5, 13, 4) {real, imag} */,
  {32'hbcc78968, 32'h3e15b681} /* (5, 13, 3) {real, imag} */,
  {32'h3f18f6e2, 32'hbdca2038} /* (5, 13, 2) {real, imag} */,
  {32'h3eb9855c, 32'h3df9b093} /* (5, 13, 1) {real, imag} */,
  {32'hbdef7c10, 32'hbe8885ee} /* (5, 13, 0) {real, imag} */,
  {32'h3e810ec2, 32'h3dd5e8ff} /* (5, 12, 31) {real, imag} */,
  {32'hbeba82db, 32'h3dd01010} /* (5, 12, 30) {real, imag} */,
  {32'h3eb0e622, 32'hbe269f62} /* (5, 12, 29) {real, imag} */,
  {32'h3dc40aae, 32'hbe83d723} /* (5, 12, 28) {real, imag} */,
  {32'h3e29bbd0, 32'h3e8f5b2e} /* (5, 12, 27) {real, imag} */,
  {32'hbefa2a50, 32'hbeef3b9b} /* (5, 12, 26) {real, imag} */,
  {32'h3f143038, 32'hbea9a46f} /* (5, 12, 25) {real, imag} */,
  {32'h3de3e5ac, 32'hbe6a61aa} /* (5, 12, 24) {real, imag} */,
  {32'h3dd04df8, 32'h3b865ec0} /* (5, 12, 23) {real, imag} */,
  {32'h3d87c3dc, 32'h3d1b2e48} /* (5, 12, 22) {real, imag} */,
  {32'h3d86d1f0, 32'hbc9fd600} /* (5, 12, 21) {real, imag} */,
  {32'h3f00e988, 32'h3eb16ad8} /* (5, 12, 20) {real, imag} */,
  {32'h3da180c9, 32'hbca5d5e8} /* (5, 12, 19) {real, imag} */,
  {32'hbf26a305, 32'hbe8552b2} /* (5, 12, 18) {real, imag} */,
  {32'hbe169107, 32'h3e3abffc} /* (5, 12, 17) {real, imag} */,
  {32'hbba02378, 32'h3d0ee302} /* (5, 12, 16) {real, imag} */,
  {32'h3edc9a3b, 32'hbe401e7c} /* (5, 12, 15) {real, imag} */,
  {32'h3e348476, 32'hbf7b357e} /* (5, 12, 14) {real, imag} */,
  {32'hbe625e4f, 32'hbb22cae0} /* (5, 12, 13) {real, imag} */,
  {32'hbdd093c2, 32'h3dbc14c6} /* (5, 12, 12) {real, imag} */,
  {32'hbec6574e, 32'h3e310006} /* (5, 12, 11) {real, imag} */,
  {32'hbeb1f893, 32'hbefd427d} /* (5, 12, 10) {real, imag} */,
  {32'h3f21872b, 32'hbeb57864} /* (5, 12, 9) {real, imag} */,
  {32'hbf0c6683, 32'hbd02331a} /* (5, 12, 8) {real, imag} */,
  {32'hbe1055fc, 32'h3ea36c39} /* (5, 12, 7) {real, imag} */,
  {32'hbe04ab83, 32'hbe37d11e} /* (5, 12, 6) {real, imag} */,
  {32'h3ea23ef4, 32'hbdb76ea4} /* (5, 12, 5) {real, imag} */,
  {32'hbed0da8d, 32'h3dd081b4} /* (5, 12, 4) {real, imag} */,
  {32'h3e24241b, 32'hbe73a5c4} /* (5, 12, 3) {real, imag} */,
  {32'hbd2e3164, 32'h3dcbf450} /* (5, 12, 2) {real, imag} */,
  {32'hbe3c0c8a, 32'h3f0dc2fd} /* (5, 12, 1) {real, imag} */,
  {32'hbdb6b83b, 32'hbe0de54f} /* (5, 12, 0) {real, imag} */,
  {32'h3e8452f9, 32'h3d34856c} /* (5, 11, 31) {real, imag} */,
  {32'h3e83f4c8, 32'h3e80b28b} /* (5, 11, 30) {real, imag} */,
  {32'hbebd9c4a, 32'h3e0808ea} /* (5, 11, 29) {real, imag} */,
  {32'h3ea660cc, 32'h3e93e792} /* (5, 11, 28) {real, imag} */,
  {32'h3d35225d, 32'h3e707d85} /* (5, 11, 27) {real, imag} */,
  {32'h3d3a3cbe, 32'hbdbb1007} /* (5, 11, 26) {real, imag} */,
  {32'hbe2f601e, 32'h3e5ae229} /* (5, 11, 25) {real, imag} */,
  {32'h3d3649ec, 32'h3c5250f4} /* (5, 11, 24) {real, imag} */,
  {32'h3e8ddaa7, 32'hbb80a580} /* (5, 11, 23) {real, imag} */,
  {32'h3d9ea37f, 32'hbf3e2b62} /* (5, 11, 22) {real, imag} */,
  {32'hbf2391b8, 32'h3e36cba8} /* (5, 11, 21) {real, imag} */,
  {32'h3d09294c, 32'h3ed68298} /* (5, 11, 20) {real, imag} */,
  {32'h3e855f9e, 32'h3f3682dc} /* (5, 11, 19) {real, imag} */,
  {32'h3d2fe550, 32'h3e4281dc} /* (5, 11, 18) {real, imag} */,
  {32'h3dcdca04, 32'hbe970c31} /* (5, 11, 17) {real, imag} */,
  {32'h3e41cf64, 32'h3ef80adc} /* (5, 11, 16) {real, imag} */,
  {32'hbea8055f, 32'hbec1d208} /* (5, 11, 15) {real, imag} */,
  {32'h3e792761, 32'hbd3b1e6e} /* (5, 11, 14) {real, imag} */,
  {32'hbd2fb4f0, 32'h3d51925c} /* (5, 11, 13) {real, imag} */,
  {32'hbc98dfa8, 32'hbe5b7208} /* (5, 11, 12) {real, imag} */,
  {32'h3f8669de, 32'hbe891faf} /* (5, 11, 11) {real, imag} */,
  {32'hbf419235, 32'hbece4880} /* (5, 11, 10) {real, imag} */,
  {32'h3e993f90, 32'h3e7cb2aa} /* (5, 11, 9) {real, imag} */,
  {32'h3e913596, 32'hbf19388d} /* (5, 11, 8) {real, imag} */,
  {32'hbf0ab3bc, 32'h3e3726a1} /* (5, 11, 7) {real, imag} */,
  {32'hbf1d2e01, 32'h3ec4937d} /* (5, 11, 6) {real, imag} */,
  {32'hbdeb6e30, 32'h3ba03940} /* (5, 11, 5) {real, imag} */,
  {32'h3df15e5c, 32'h3e25fda6} /* (5, 11, 4) {real, imag} */,
  {32'h3eb85ce4, 32'hbece1650} /* (5, 11, 3) {real, imag} */,
  {32'h3df263ba, 32'hbde5f150} /* (5, 11, 2) {real, imag} */,
  {32'h3cf3e850, 32'hbdd2a51c} /* (5, 11, 1) {real, imag} */,
  {32'h3ec28fa2, 32'h3e02283a} /* (5, 11, 0) {real, imag} */,
  {32'h3bc85d00, 32'hbf204356} /* (5, 10, 31) {real, imag} */,
  {32'hbd8228fa, 32'hbecf340e} /* (5, 10, 30) {real, imag} */,
  {32'hbf08572e, 32'hbc8c3ef0} /* (5, 10, 29) {real, imag} */,
  {32'hbe665807, 32'hbef34f98} /* (5, 10, 28) {real, imag} */,
  {32'h3f245438, 32'h3ed35840} /* (5, 10, 27) {real, imag} */,
  {32'hbd6a1660, 32'h3f40d422} /* (5, 10, 26) {real, imag} */,
  {32'h3ef63b46, 32'h3ced8c98} /* (5, 10, 25) {real, imag} */,
  {32'hbef940ab, 32'hbdc93e24} /* (5, 10, 24) {real, imag} */,
  {32'h3b82ad60, 32'h3dcb63d0} /* (5, 10, 23) {real, imag} */,
  {32'h3ea216bb, 32'h3d2e9bd0} /* (5, 10, 22) {real, imag} */,
  {32'hbef37412, 32'hbef363c6} /* (5, 10, 21) {real, imag} */,
  {32'hbe05de3c, 32'h3d0b5d20} /* (5, 10, 20) {real, imag} */,
  {32'h3eb24e00, 32'hbe95c321} /* (5, 10, 19) {real, imag} */,
  {32'h3ec9bc5b, 32'hbcf7b5a0} /* (5, 10, 18) {real, imag} */,
  {32'h3e4c5d40, 32'hbdf6f8e0} /* (5, 10, 17) {real, imag} */,
  {32'h3df3b228, 32'hbee704f8} /* (5, 10, 16) {real, imag} */,
  {32'h3ef5f945, 32'h3d810e84} /* (5, 10, 15) {real, imag} */,
  {32'hbddf35bf, 32'hbea103e9} /* (5, 10, 14) {real, imag} */,
  {32'h3e8bdff8, 32'hbd064b18} /* (5, 10, 13) {real, imag} */,
  {32'hbe29ffeb, 32'hbf030938} /* (5, 10, 12) {real, imag} */,
  {32'hbea71ce0, 32'h3e7cc2e8} /* (5, 10, 11) {real, imag} */,
  {32'hbe73928f, 32'h3e2b51c0} /* (5, 10, 10) {real, imag} */,
  {32'hbeb58b81, 32'h3e51b6d8} /* (5, 10, 9) {real, imag} */,
  {32'h3ea0c52b, 32'hbdb5ad86} /* (5, 10, 8) {real, imag} */,
  {32'h3efa40ef, 32'h3f6912dc} /* (5, 10, 7) {real, imag} */,
  {32'hbe38f7ae, 32'h3e54b468} /* (5, 10, 6) {real, imag} */,
  {32'hbe94e008, 32'h3d53c355} /* (5, 10, 5) {real, imag} */,
  {32'h3e76b8ec, 32'hbed12cfb} /* (5, 10, 4) {real, imag} */,
  {32'hbe40d714, 32'hbee7400a} /* (5, 10, 3) {real, imag} */,
  {32'hbd3fcfc0, 32'hbba808c0} /* (5, 10, 2) {real, imag} */,
  {32'hbe0dabc1, 32'h3dd74f13} /* (5, 10, 1) {real, imag} */,
  {32'hbd981a96, 32'hbdfa0e62} /* (5, 10, 0) {real, imag} */,
  {32'h3c7e92c0, 32'hbecba3d6} /* (5, 9, 31) {real, imag} */,
  {32'h3eecaea1, 32'h3dbb0e50} /* (5, 9, 30) {real, imag} */,
  {32'hbe4f04b8, 32'h3dda12e7} /* (5, 9, 29) {real, imag} */,
  {32'hbc8d0ef0, 32'h3d8a337b} /* (5, 9, 28) {real, imag} */,
  {32'h3ea1adaa, 32'h3dc6052e} /* (5, 9, 27) {real, imag} */,
  {32'h3e8ca1db, 32'h3e4be539} /* (5, 9, 26) {real, imag} */,
  {32'h3e83f7d9, 32'hbd0a971e} /* (5, 9, 25) {real, imag} */,
  {32'h3ea00395, 32'hbf15590e} /* (5, 9, 24) {real, imag} */,
  {32'hbe9510a3, 32'h3ea0a68c} /* (5, 9, 23) {real, imag} */,
  {32'h3ee0129a, 32'h3f303b75} /* (5, 9, 22) {real, imag} */,
  {32'h3e75fd1e, 32'hbf4b0d00} /* (5, 9, 21) {real, imag} */,
  {32'hbe9d05cb, 32'h3f2c9d6f} /* (5, 9, 20) {real, imag} */,
  {32'hbd88a902, 32'h3dff1d1e} /* (5, 9, 19) {real, imag} */,
  {32'hbe0a96b0, 32'h3cc13bb0} /* (5, 9, 18) {real, imag} */,
  {32'hbeba543b, 32'h3ef82337} /* (5, 9, 17) {real, imag} */,
  {32'h3eb4b578, 32'h3d3bcba4} /* (5, 9, 16) {real, imag} */,
  {32'hbed15fac, 32'h3d9f29bd} /* (5, 9, 15) {real, imag} */,
  {32'hbda6930c, 32'hbd842717} /* (5, 9, 14) {real, imag} */,
  {32'h3ed69261, 32'h3ea596f1} /* (5, 9, 13) {real, imag} */,
  {32'hbd64dd5a, 32'hbcc7e6b4} /* (5, 9, 12) {real, imag} */,
  {32'hbd040fa8, 32'h3d935475} /* (5, 9, 11) {real, imag} */,
  {32'hbcc5e3f0, 32'h3e56f1f7} /* (5, 9, 10) {real, imag} */,
  {32'h3e209265, 32'hbc5ebbe0} /* (5, 9, 9) {real, imag} */,
  {32'h3efd1c13, 32'h3de0c50e} /* (5, 9, 8) {real, imag} */,
  {32'h3eb9749e, 32'hbe2621b5} /* (5, 9, 7) {real, imag} */,
  {32'hbe7d489a, 32'h3dbb11f4} /* (5, 9, 6) {real, imag} */,
  {32'hbdef98d2, 32'h3d33b218} /* (5, 9, 5) {real, imag} */,
  {32'hbd7f1fc9, 32'hbf06e5ad} /* (5, 9, 4) {real, imag} */,
  {32'h3eab8df4, 32'h3f05d461} /* (5, 9, 3) {real, imag} */,
  {32'h3dd0b726, 32'hbf4f311e} /* (5, 9, 2) {real, imag} */,
  {32'hbbe20460, 32'hbdc2bd24} /* (5, 9, 1) {real, imag} */,
  {32'hbf4b01aa, 32'h3e699c2b} /* (5, 9, 0) {real, imag} */,
  {32'h3f48c834, 32'h3db78f20} /* (5, 8, 31) {real, imag} */,
  {32'hbf04ca1b, 32'h3e7c7f3c} /* (5, 8, 30) {real, imag} */,
  {32'h3f9cdcc2, 32'h3f3ae395} /* (5, 8, 29) {real, imag} */,
  {32'hbef708f6, 32'hbc9ab9f8} /* (5, 8, 28) {real, imag} */,
  {32'hbcc70b30, 32'hbe2e78c8} /* (5, 8, 27) {real, imag} */,
  {32'h3ecd5601, 32'h3eb262ae} /* (5, 8, 26) {real, imag} */,
  {32'h3e997b30, 32'h3efcb568} /* (5, 8, 25) {real, imag} */,
  {32'hbea19344, 32'h3e8adec8} /* (5, 8, 24) {real, imag} */,
  {32'h3deed3b4, 32'hbf49870d} /* (5, 8, 23) {real, imag} */,
  {32'hbebb29f2, 32'h3d883ea6} /* (5, 8, 22) {real, imag} */,
  {32'hbe8895d0, 32'hbd3520fc} /* (5, 8, 21) {real, imag} */,
  {32'hbdfd75ec, 32'hbf2ae442} /* (5, 8, 20) {real, imag} */,
  {32'hbdaa7c90, 32'hbc8f4f8c} /* (5, 8, 19) {real, imag} */,
  {32'h3e018228, 32'h3e88c96f} /* (5, 8, 18) {real, imag} */,
  {32'hbd228ffe, 32'hbe7f0ae5} /* (5, 8, 17) {real, imag} */,
  {32'h3d550078, 32'h3b159f00} /* (5, 8, 16) {real, imag} */,
  {32'h3e0404e8, 32'h3ed579f0} /* (5, 8, 15) {real, imag} */,
  {32'hbf246d56, 32'hbcc38f70} /* (5, 8, 14) {real, imag} */,
  {32'h3e88043d, 32'hbd945a0c} /* (5, 8, 13) {real, imag} */,
  {32'hbde032ec, 32'hbe976986} /* (5, 8, 12) {real, imag} */,
  {32'hbe006a5d, 32'hbdea46d8} /* (5, 8, 11) {real, imag} */,
  {32'h3e229406, 32'hbd16a530} /* (5, 8, 10) {real, imag} */,
  {32'h3ecb9567, 32'h3f6a13d1} /* (5, 8, 9) {real, imag} */,
  {32'h3f22d6f9, 32'hbf1d4ef0} /* (5, 8, 8) {real, imag} */,
  {32'h3c1451a0, 32'hbf457def} /* (5, 8, 7) {real, imag} */,
  {32'h3ed6a992, 32'hbd834150} /* (5, 8, 6) {real, imag} */,
  {32'hbf35eea0, 32'h3ec09eed} /* (5, 8, 5) {real, imag} */,
  {32'h3e66258a, 32'hbdcb7efa} /* (5, 8, 4) {real, imag} */,
  {32'hbe344206, 32'hbe1a4529} /* (5, 8, 3) {real, imag} */,
  {32'h3e713ecb, 32'hbe6f1504} /* (5, 8, 2) {real, imag} */,
  {32'hbe912e80, 32'hbe753e30} /* (5, 8, 1) {real, imag} */,
  {32'h3f008bc4, 32'hbafda380} /* (5, 8, 0) {real, imag} */,
  {32'h3d4581c8, 32'h3df0a808} /* (5, 7, 31) {real, imag} */,
  {32'hbefd8e0f, 32'hbe9ecef2} /* (5, 7, 30) {real, imag} */,
  {32'hbe68f533, 32'hbe0af9b9} /* (5, 7, 29) {real, imag} */,
  {32'hbf387f12, 32'hbf29df0d} /* (5, 7, 28) {real, imag} */,
  {32'hbf14175a, 32'hbdb2148b} /* (5, 7, 27) {real, imag} */,
  {32'hbc9f5088, 32'hbd6e2380} /* (5, 7, 26) {real, imag} */,
  {32'h3ed88aaa, 32'hbe9614e8} /* (5, 7, 25) {real, imag} */,
  {32'hbeb20a57, 32'h3c8d35c0} /* (5, 7, 24) {real, imag} */,
  {32'hbeb261c1, 32'h3ea7cffe} /* (5, 7, 23) {real, imag} */,
  {32'h3f0c4dce, 32'h3b94a840} /* (5, 7, 22) {real, imag} */,
  {32'h3e331f54, 32'h3f24a22c} /* (5, 7, 21) {real, imag} */,
  {32'h3f23d00a, 32'hbeb57b93} /* (5, 7, 20) {real, imag} */,
  {32'hbed5d0e7, 32'h3cfdc1bc} /* (5, 7, 19) {real, imag} */,
  {32'h3e46bf23, 32'h3dea803c} /* (5, 7, 18) {real, imag} */,
  {32'h3e61d406, 32'h3d4c68ca} /* (5, 7, 17) {real, imag} */,
  {32'hb98ca000, 32'hbe7862e6} /* (5, 7, 16) {real, imag} */,
  {32'hbe88002e, 32'h3eaa0ed7} /* (5, 7, 15) {real, imag} */,
  {32'hbf120707, 32'hbe53b173} /* (5, 7, 14) {real, imag} */,
  {32'hbed7c307, 32'h3e289e3a} /* (5, 7, 13) {real, imag} */,
  {32'hbddb13d8, 32'hbdc6b91b} /* (5, 7, 12) {real, imag} */,
  {32'hbde91222, 32'h3cf65400} /* (5, 7, 11) {real, imag} */,
  {32'h3ee1f372, 32'h3f252934} /* (5, 7, 10) {real, imag} */,
  {32'h3eb93cf0, 32'h3e235dd0} /* (5, 7, 9) {real, imag} */,
  {32'h3e6ecada, 32'hbe8f0c44} /* (5, 7, 8) {real, imag} */,
  {32'hba674b00, 32'hbe471e1a} /* (5, 7, 7) {real, imag} */,
  {32'h3ef19e32, 32'h3e8074f6} /* (5, 7, 6) {real, imag} */,
  {32'h3e739498, 32'h3f553d65} /* (5, 7, 5) {real, imag} */,
  {32'h3e1e4d49, 32'h3df467e9} /* (5, 7, 4) {real, imag} */,
  {32'hbedcdeb8, 32'hbe8c5c02} /* (5, 7, 3) {real, imag} */,
  {32'hbdb6ac94, 32'h3f284746} /* (5, 7, 2) {real, imag} */,
  {32'hbe404a2c, 32'hbe412c74} /* (5, 7, 1) {real, imag} */,
  {32'hbf4d6622, 32'hbebf51a2} /* (5, 7, 0) {real, imag} */,
  {32'h3e998fc4, 32'h3f0085d1} /* (5, 6, 31) {real, imag} */,
  {32'hbed13f72, 32'hbe5dfb50} /* (5, 6, 30) {real, imag} */,
  {32'h3ed9d75c, 32'hbdf818f2} /* (5, 6, 29) {real, imag} */,
  {32'h3e246f0c, 32'h3dc8b702} /* (5, 6, 28) {real, imag} */,
  {32'h3e9fd09a, 32'h3e9117ca} /* (5, 6, 27) {real, imag} */,
  {32'hbe543026, 32'hbea28410} /* (5, 6, 26) {real, imag} */,
  {32'h3d3e8ef0, 32'h3f3f54c4} /* (5, 6, 25) {real, imag} */,
  {32'hbe1a1248, 32'hbe8a33c2} /* (5, 6, 24) {real, imag} */,
  {32'hbeb20f12, 32'h3d83fec0} /* (5, 6, 23) {real, imag} */,
  {32'hbe410445, 32'h3e9a4a3e} /* (5, 6, 22) {real, imag} */,
  {32'hbe928324, 32'hbd122710} /* (5, 6, 21) {real, imag} */,
  {32'hbe351ba0, 32'hbd838da6} /* (5, 6, 20) {real, imag} */,
  {32'h3e841f64, 32'h3e6c22ca} /* (5, 6, 19) {real, imag} */,
  {32'h3e5a7398, 32'h3e3755c4} /* (5, 6, 18) {real, imag} */,
  {32'hbec1dec0, 32'hbe673c00} /* (5, 6, 17) {real, imag} */,
  {32'h3e9d9664, 32'hbe1e84f9} /* (5, 6, 16) {real, imag} */,
  {32'hbe35093c, 32'hbc9d8fb0} /* (5, 6, 15) {real, imag} */,
  {32'h3e9e5949, 32'h3e90a921} /* (5, 6, 14) {real, imag} */,
  {32'hbceebc44, 32'h3da115cc} /* (5, 6, 13) {real, imag} */,
  {32'h3ef76cf8, 32'hbe9fda51} /* (5, 6, 12) {real, imag} */,
  {32'hbe34b2c8, 32'h3f4a9f41} /* (5, 6, 11) {real, imag} */,
  {32'h3ef1ac8c, 32'h3db35291} /* (5, 6, 10) {real, imag} */,
  {32'h3dbe11b5, 32'hbedb7dc6} /* (5, 6, 9) {real, imag} */,
  {32'hbee656ca, 32'hbe9d9254} /* (5, 6, 8) {real, imag} */,
  {32'h3f30b280, 32'h3ecb180e} /* (5, 6, 7) {real, imag} */,
  {32'hbee65fb4, 32'h3ed859f0} /* (5, 6, 6) {real, imag} */,
  {32'hbe02b7ec, 32'h3eb3b206} /* (5, 6, 5) {real, imag} */,
  {32'hbdf6ee08, 32'h3e6df240} /* (5, 6, 4) {real, imag} */,
  {32'hbf10c6c7, 32'hbf518a6a} /* (5, 6, 3) {real, imag} */,
  {32'hbf27baa6, 32'hbe947dc7} /* (5, 6, 2) {real, imag} */,
  {32'hbe47c574, 32'h3e91f4fc} /* (5, 6, 1) {real, imag} */,
  {32'h3f5fb55f, 32'h3d99fc88} /* (5, 6, 0) {real, imag} */,
  {32'h3f53eb6e, 32'h3fcbbef5} /* (5, 5, 31) {real, imag} */,
  {32'hbe97236a, 32'hbe96ccb4} /* (5, 5, 30) {real, imag} */,
  {32'hbf2a7356, 32'hbf0ffdd3} /* (5, 5, 29) {real, imag} */,
  {32'hbea55a2d, 32'hbe1cb3a8} /* (5, 5, 28) {real, imag} */,
  {32'hbf0e1474, 32'h3f0cc338} /* (5, 5, 27) {real, imag} */,
  {32'h3e843aba, 32'h3f1c612a} /* (5, 5, 26) {real, imag} */,
  {32'h3e0c633e, 32'h3e3357cb} /* (5, 5, 25) {real, imag} */,
  {32'hbf86198c, 32'h3e713ff4} /* (5, 5, 24) {real, imag} */,
  {32'hbe648fd3, 32'h3ef1ab4c} /* (5, 5, 23) {real, imag} */,
  {32'hbf094323, 32'hbf247f57} /* (5, 5, 22) {real, imag} */,
  {32'hbe151511, 32'hbeb50d00} /* (5, 5, 21) {real, imag} */,
  {32'hbe79b317, 32'hbea42bfc} /* (5, 5, 20) {real, imag} */,
  {32'hbf17544b, 32'h3ea4f7b0} /* (5, 5, 19) {real, imag} */,
  {32'hbea9bb6a, 32'h3d5c5dd0} /* (5, 5, 18) {real, imag} */,
  {32'hbcf23f26, 32'hbe58b7c0} /* (5, 5, 17) {real, imag} */,
  {32'h3dbc5b44, 32'h3d8bc834} /* (5, 5, 16) {real, imag} */,
  {32'hbe437a24, 32'h3cce99d0} /* (5, 5, 15) {real, imag} */,
  {32'h3e90f440, 32'h3d279ab0} /* (5, 5, 14) {real, imag} */,
  {32'h3ec3b0f5, 32'h3ef2e301} /* (5, 5, 13) {real, imag} */,
  {32'h3de5d141, 32'h3d052890} /* (5, 5, 12) {real, imag} */,
  {32'h3ea9aed5, 32'hbe643aae} /* (5, 5, 11) {real, imag} */,
  {32'h3d8bf216, 32'h3f0b22d7} /* (5, 5, 10) {real, imag} */,
  {32'hbebc02c4, 32'h3debb5b2} /* (5, 5, 9) {real, imag} */,
  {32'h3e0314cb, 32'h3cb04f04} /* (5, 5, 8) {real, imag} */,
  {32'hbe900a19, 32'hbe1db134} /* (5, 5, 7) {real, imag} */,
  {32'h3e99459e, 32'hbe76ff96} /* (5, 5, 6) {real, imag} */,
  {32'hbf25ea98, 32'h3e313d60} /* (5, 5, 5) {real, imag} */,
  {32'hbf2c5ab0, 32'h3e75a5a7} /* (5, 5, 4) {real, imag} */,
  {32'h3f121aa2, 32'h3d95bdc8} /* (5, 5, 3) {real, imag} */,
  {32'hbdb35e44, 32'h3f28c87a} /* (5, 5, 2) {real, imag} */,
  {32'h3f30f85b, 32'h3e42a416} /* (5, 5, 1) {real, imag} */,
  {32'h3ec555c0, 32'h3ebd4a1d} /* (5, 5, 0) {real, imag} */,
  {32'hbf3dc213, 32'hbf5a51e3} /* (5, 4, 31) {real, imag} */,
  {32'h3e163ce8, 32'h3f4fc354} /* (5, 4, 30) {real, imag} */,
  {32'h3de3e05d, 32'h3c5388e0} /* (5, 4, 29) {real, imag} */,
  {32'h3dcaacb2, 32'h3f038016} /* (5, 4, 28) {real, imag} */,
  {32'h3ea3e4e8, 32'hbf39a4fa} /* (5, 4, 27) {real, imag} */,
  {32'hbf33df08, 32'hbea3a6f8} /* (5, 4, 26) {real, imag} */,
  {32'h3e033a1c, 32'h3f0ca0ee} /* (5, 4, 25) {real, imag} */,
  {32'h3f0513a0, 32'hbebf80f6} /* (5, 4, 24) {real, imag} */,
  {32'h3e1053ae, 32'h3da8cc36} /* (5, 4, 23) {real, imag} */,
  {32'h3e7c4804, 32'h3de13fb9} /* (5, 4, 22) {real, imag} */,
  {32'h3e9d3956, 32'hbec1769a} /* (5, 4, 21) {real, imag} */,
  {32'h3e9c0740, 32'h3f30f3f4} /* (5, 4, 20) {real, imag} */,
  {32'hbe8757a0, 32'h3e5a7be6} /* (5, 4, 19) {real, imag} */,
  {32'hbec59a7d, 32'h3e6c0dc0} /* (5, 4, 18) {real, imag} */,
  {32'h3e5093aa, 32'h3d8f0679} /* (5, 4, 17) {real, imag} */,
  {32'hbe35a500, 32'h3e40947a} /* (5, 4, 16) {real, imag} */,
  {32'hbd122ef4, 32'hbd85d776} /* (5, 4, 15) {real, imag} */,
  {32'h3e9636c0, 32'h3ef555e4} /* (5, 4, 14) {real, imag} */,
  {32'hbeffb710, 32'hbe345d8e} /* (5, 4, 13) {real, imag} */,
  {32'hbe77a766, 32'h3edd9f64} /* (5, 4, 12) {real, imag} */,
  {32'h3eec92c8, 32'h3eb8d52b} /* (5, 4, 11) {real, imag} */,
  {32'h3e34f5f8, 32'hbf412023} /* (5, 4, 10) {real, imag} */,
  {32'hbf06559a, 32'hbdab3a16} /* (5, 4, 9) {real, imag} */,
  {32'h3e4286f5, 32'h3edbdea7} /* (5, 4, 8) {real, imag} */,
  {32'hbf2154e8, 32'hbd9cf48c} /* (5, 4, 7) {real, imag} */,
  {32'hbd7564a8, 32'h3d8440a2} /* (5, 4, 6) {real, imag} */,
  {32'h3ea869ff, 32'h3df8d2e8} /* (5, 4, 5) {real, imag} */,
  {32'h3f2c6584, 32'hbdd7dc70} /* (5, 4, 4) {real, imag} */,
  {32'hbf40fcdb, 32'h3f555504} /* (5, 4, 3) {real, imag} */,
  {32'h3f495216, 32'hbecf0d84} /* (5, 4, 2) {real, imag} */,
  {32'hc01bb8b4, 32'h3efeec40} /* (5, 4, 1) {real, imag} */,
  {32'h3eecc939, 32'hbf1148c0} /* (5, 4, 0) {real, imag} */,
  {32'h3e666eb8, 32'hbfb21549} /* (5, 3, 31) {real, imag} */,
  {32'hbea8df48, 32'hbfa72ee2} /* (5, 3, 30) {real, imag} */,
  {32'h3d80ca96, 32'h3ee5ae72} /* (5, 3, 29) {real, imag} */,
  {32'hbec7d1a5, 32'h3de85338} /* (5, 3, 28) {real, imag} */,
  {32'hbea280e9, 32'hbf29ae8a} /* (5, 3, 27) {real, imag} */,
  {32'hbf56869f, 32'hbe31d670} /* (5, 3, 26) {real, imag} */,
  {32'hbec8c62a, 32'h3f0575b2} /* (5, 3, 25) {real, imag} */,
  {32'h3f32f2b8, 32'hbe00b4a0} /* (5, 3, 24) {real, imag} */,
  {32'h3eff16f8, 32'hbde6b7cc} /* (5, 3, 23) {real, imag} */,
  {32'hbdbab9b4, 32'hbe7d48bf} /* (5, 3, 22) {real, imag} */,
  {32'hbde46820, 32'h3e87ea03} /* (5, 3, 21) {real, imag} */,
  {32'h3f425ffc, 32'hbc24ff00} /* (5, 3, 20) {real, imag} */,
  {32'h3d4381a2, 32'h3eb2229f} /* (5, 3, 19) {real, imag} */,
  {32'hbdcaf1af, 32'hbdb22665} /* (5, 3, 18) {real, imag} */,
  {32'hbd8b5172, 32'h3e1722b0} /* (5, 3, 17) {real, imag} */,
  {32'hbe63e7d6, 32'hbdaf8c2e} /* (5, 3, 16) {real, imag} */,
  {32'h3ebe8ced, 32'hbdd02368} /* (5, 3, 15) {real, imag} */,
  {32'h3e727b56, 32'hbebbdd81} /* (5, 3, 14) {real, imag} */,
  {32'h3ec5e166, 32'h3e0737b9} /* (5, 3, 13) {real, imag} */,
  {32'hbe4aedd3, 32'hbde3fdbc} /* (5, 3, 12) {real, imag} */,
  {32'hbee4a6f0, 32'hbf04311a} /* (5, 3, 11) {real, imag} */,
  {32'h3e38ed07, 32'hbe835e4b} /* (5, 3, 10) {real, imag} */,
  {32'h3c204300, 32'hbe4ade51} /* (5, 3, 9) {real, imag} */,
  {32'hbde75284, 32'h3ee8f030} /* (5, 3, 8) {real, imag} */,
  {32'hbea4e860, 32'hbf588e82} /* (5, 3, 7) {real, imag} */,
  {32'h3d1133d8, 32'hbf09c1ca} /* (5, 3, 6) {real, imag} */,
  {32'hbeb9ce16, 32'hbea959d8} /* (5, 3, 5) {real, imag} */,
  {32'h3e99a51e, 32'h3e72991e} /* (5, 3, 4) {real, imag} */,
  {32'hbe9be700, 32'h3eb04cda} /* (5, 3, 3) {real, imag} */,
  {32'h3f8ccf79, 32'h400f49d4} /* (5, 3, 2) {real, imag} */,
  {32'h3ecdc5ec, 32'h3fc72d42} /* (5, 3, 1) {real, imag} */,
  {32'h3f00fbc1, 32'h3fd02bfb} /* (5, 3, 0) {real, imag} */,
  {32'hbeb3b740, 32'h3d213220} /* (5, 2, 31) {real, imag} */,
  {32'h3f4c8e18, 32'hbea0cfc0} /* (5, 2, 30) {real, imag} */,
  {32'h3c68f2a0, 32'h3f4aec4b} /* (5, 2, 29) {real, imag} */,
  {32'h3ec8cbb6, 32'hbf203f07} /* (5, 2, 28) {real, imag} */,
  {32'hbf7bb23d, 32'h3e1478f8} /* (5, 2, 27) {real, imag} */,
  {32'hbf5dc0ea, 32'h3f279de6} /* (5, 2, 26) {real, imag} */,
  {32'h3ed844fa, 32'hbe99bcf4} /* (5, 2, 25) {real, imag} */,
  {32'h3e8a1216, 32'h3f97f9fd} /* (5, 2, 24) {real, imag} */,
  {32'hbd122184, 32'hbdb564d5} /* (5, 2, 23) {real, imag} */,
  {32'h3db22634, 32'hbe5d055c} /* (5, 2, 22) {real, imag} */,
  {32'hbe3ca46b, 32'h3e8931f6} /* (5, 2, 21) {real, imag} */,
  {32'h3edc5e12, 32'h3dbbf454} /* (5, 2, 20) {real, imag} */,
  {32'hbe0a04a7, 32'hbee593ee} /* (5, 2, 19) {real, imag} */,
  {32'hbd44fca8, 32'hbde3166a} /* (5, 2, 18) {real, imag} */,
  {32'h3e489513, 32'hbe66a7aa} /* (5, 2, 17) {real, imag} */,
  {32'h3e2d36a2, 32'hbdf7a9c0} /* (5, 2, 16) {real, imag} */,
  {32'hbe69b948, 32'h3e3aa6bc} /* (5, 2, 15) {real, imag} */,
  {32'h3a183500, 32'hbe7a9fd2} /* (5, 2, 14) {real, imag} */,
  {32'hbcf721f6, 32'h3a16c400} /* (5, 2, 13) {real, imag} */,
  {32'h3d093194, 32'hbdf2a765} /* (5, 2, 12) {real, imag} */,
  {32'hbe050fc0, 32'hbe85ed4b} /* (5, 2, 11) {real, imag} */,
  {32'hbebba530, 32'h3e2734c4} /* (5, 2, 10) {real, imag} */,
  {32'h3e0d99a5, 32'h3f72d973} /* (5, 2, 9) {real, imag} */,
  {32'h3d3c7780, 32'hbdf81028} /* (5, 2, 8) {real, imag} */,
  {32'hbe0e2d9e, 32'hbedad9da} /* (5, 2, 7) {real, imag} */,
  {32'h3de43a27, 32'h3f0aa4ce} /* (5, 2, 6) {real, imag} */,
  {32'h3f57b7b1, 32'hbf8572b9} /* (5, 2, 5) {real, imag} */,
  {32'h3e69d564, 32'h3f37755f} /* (5, 2, 4) {real, imag} */,
  {32'hbc8c5e20, 32'h3e53845a} /* (5, 2, 3) {real, imag} */,
  {32'hbfe434ce, 32'h40233f10} /* (5, 2, 2) {real, imag} */,
  {32'h3f37f910, 32'h3f9e8910} /* (5, 2, 1) {real, imag} */,
  {32'hc014f34e, 32'hbfe141c1} /* (5, 2, 0) {real, imag} */,
  {32'h40e4b078, 32'hc056416a} /* (5, 1, 31) {real, imag} */,
  {32'h3f36ace0, 32'hbd28e240} /* (5, 1, 30) {real, imag} */,
  {32'h3fe71a97, 32'hbee16697} /* (5, 1, 29) {real, imag} */,
  {32'h3e2bdf6e, 32'hbf3f581d} /* (5, 1, 28) {real, imag} */,
  {32'h3f0af44c, 32'h3edf17a4} /* (5, 1, 27) {real, imag} */,
  {32'h3e962453, 32'hbebb854e} /* (5, 1, 26) {real, imag} */,
  {32'hbfabb13e, 32'hbdeb6a01} /* (5, 1, 25) {real, imag} */,
  {32'h3df48864, 32'hbe945451} /* (5, 1, 24) {real, imag} */,
  {32'h3ed8dd67, 32'hbe8f8268} /* (5, 1, 23) {real, imag} */,
  {32'hbdf2237e, 32'hbdbcf99a} /* (5, 1, 22) {real, imag} */,
  {32'hbe8faa5a, 32'h3b5df380} /* (5, 1, 21) {real, imag} */,
  {32'h3e323de7, 32'hbec0ed13} /* (5, 1, 20) {real, imag} */,
  {32'h3d83e909, 32'hbe8817c7} /* (5, 1, 19) {real, imag} */,
  {32'hbe0f312c, 32'hbeb0c575} /* (5, 1, 18) {real, imag} */,
  {32'h3dc76a4a, 32'hbc5a9ad0} /* (5, 1, 17) {real, imag} */,
  {32'h3d804ef8, 32'hbe329433} /* (5, 1, 16) {real, imag} */,
  {32'h3e0d8ff3, 32'h3e2f6c15} /* (5, 1, 15) {real, imag} */,
  {32'h3e977e17, 32'hbea9c5c3} /* (5, 1, 14) {real, imag} */,
  {32'h3ea3cbba, 32'h3e174527} /* (5, 1, 13) {real, imag} */,
  {32'h3e4e8303, 32'hbd9a8872} /* (5, 1, 12) {real, imag} */,
  {32'h3ed92f8f, 32'hbec2139a} /* (5, 1, 11) {real, imag} */,
  {32'hbe8c54b5, 32'hbea38f9a} /* (5, 1, 10) {real, imag} */,
  {32'hbf09c200, 32'h3edb87cb} /* (5, 1, 9) {real, imag} */,
  {32'h3f5a4d77, 32'h3e683474} /* (5, 1, 8) {real, imag} */,
  {32'hbe25dcbc, 32'h3f058868} /* (5, 1, 7) {real, imag} */,
  {32'hbf2ee3e4, 32'hbece317d} /* (5, 1, 6) {real, imag} */,
  {32'hbeae5fb8, 32'h3f38a617} /* (5, 1, 5) {real, imag} */,
  {32'h3f4ad6a5, 32'hbf8f0810} /* (5, 1, 4) {real, imag} */,
  {32'hbe8d3652, 32'hbfdc2658} /* (5, 1, 3) {real, imag} */,
  {32'hbe5733e0, 32'hbee0f640} /* (5, 1, 2) {real, imag} */,
  {32'h413db712, 32'h3fee91b4} /* (5, 1, 1) {real, imag} */,
  {32'h418da16e, 32'h409b2d54} /* (5, 1, 0) {real, imag} */,
  {32'h410356ac, 32'hc0f93bbd} /* (5, 0, 31) {real, imag} */,
  {32'h3f43ad50, 32'h3fbc8958} /* (5, 0, 30) {real, imag} */,
  {32'h402dd7ae, 32'hbff1b01a} /* (5, 0, 29) {real, imag} */,
  {32'hbe371328, 32'hbf87e979} /* (5, 0, 28) {real, imag} */,
  {32'hbe1187dc, 32'h3ec67ab6} /* (5, 0, 27) {real, imag} */,
  {32'h3f9dceac, 32'h3e216244} /* (5, 0, 26) {real, imag} */,
  {32'h3d7a7ad0, 32'h3e9f5024} /* (5, 0, 25) {real, imag} */,
  {32'h3bab5990, 32'hbf552410} /* (5, 0, 24) {real, imag} */,
  {32'hbd375518, 32'h3f667ff8} /* (5, 0, 23) {real, imag} */,
  {32'hbf1fab31, 32'h3f0ff853} /* (5, 0, 22) {real, imag} */,
  {32'hbeb81530, 32'h3e0008e0} /* (5, 0, 21) {real, imag} */,
  {32'hbf22b0b6, 32'h3c0047b0} /* (5, 0, 20) {real, imag} */,
  {32'hbe3f891d, 32'h3e884f85} /* (5, 0, 19) {real, imag} */,
  {32'hbcd53c18, 32'h3ea7789c} /* (5, 0, 18) {real, imag} */,
  {32'hbeafc400, 32'h3e380350} /* (5, 0, 17) {real, imag} */,
  {32'hbeb96b34, 32'h00000000} /* (5, 0, 16) {real, imag} */,
  {32'hbeafc400, 32'hbe380350} /* (5, 0, 15) {real, imag} */,
  {32'hbcd53c18, 32'hbea7789c} /* (5, 0, 14) {real, imag} */,
  {32'hbe3f891d, 32'hbe884f85} /* (5, 0, 13) {real, imag} */,
  {32'hbf22b0b6, 32'hbc0047b0} /* (5, 0, 12) {real, imag} */,
  {32'hbeb81530, 32'hbe0008e0} /* (5, 0, 11) {real, imag} */,
  {32'hbf1fab31, 32'hbf0ff853} /* (5, 0, 10) {real, imag} */,
  {32'hbd375518, 32'hbf667ff8} /* (5, 0, 9) {real, imag} */,
  {32'h3bab5990, 32'h3f552410} /* (5, 0, 8) {real, imag} */,
  {32'h3d7a7ad0, 32'hbe9f5024} /* (5, 0, 7) {real, imag} */,
  {32'h3f9dceac, 32'hbe216244} /* (5, 0, 6) {real, imag} */,
  {32'hbe1187dc, 32'hbec67ab6} /* (5, 0, 5) {real, imag} */,
  {32'hbe371328, 32'h3f87e979} /* (5, 0, 4) {real, imag} */,
  {32'h402dd7ae, 32'h3ff1b01a} /* (5, 0, 3) {real, imag} */,
  {32'h3f43ad50, 32'hbfbc8958} /* (5, 0, 2) {real, imag} */,
  {32'h410356ac, 32'h40f93bbd} /* (5, 0, 1) {real, imag} */,
  {32'h41f6a686, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hc13b4b8d, 32'h412d18d3} /* (4, 31, 31) {real, imag} */,
  {32'h40e356ee, 32'hc0bbd49a} /* (4, 31, 30) {real, imag} */,
  {32'h3ecbffd6, 32'h3fcb2118} /* (4, 31, 29) {real, imag} */,
  {32'h3e1f04c4, 32'h3fa3ec2c} /* (4, 31, 28) {real, imag} */,
  {32'h3ff8e9ef, 32'hbf53ca10} /* (4, 31, 27) {real, imag} */,
  {32'hbf311f6b, 32'h3f4bc0dd} /* (4, 31, 26) {real, imag} */,
  {32'hbeeb9284, 32'h3db51bf0} /* (4, 31, 25) {real, imag} */,
  {32'h3d074130, 32'hbf964f38} /* (4, 31, 24) {real, imag} */,
  {32'hbf2ba055, 32'hbf05b886} /* (4, 31, 23) {real, imag} */,
  {32'h3e80b80e, 32'hbdf1e4ad} /* (4, 31, 22) {real, imag} */,
  {32'hbe3badc9, 32'hbf0922e1} /* (4, 31, 21) {real, imag} */,
  {32'hbdee09ec, 32'h3e2d394b} /* (4, 31, 20) {real, imag} */,
  {32'h3e373c2e, 32'h3ddaeacf} /* (4, 31, 19) {real, imag} */,
  {32'hbf463230, 32'hbf11c066} /* (4, 31, 18) {real, imag} */,
  {32'h3eb9a562, 32'hbd9c5e2a} /* (4, 31, 17) {real, imag} */,
  {32'hbed63d96, 32'h3e87be28} /* (4, 31, 16) {real, imag} */,
  {32'h3e9b17d8, 32'hbea7b11e} /* (4, 31, 15) {real, imag} */,
  {32'h3e16341b, 32'h3f0e4304} /* (4, 31, 14) {real, imag} */,
  {32'h3e340592, 32'h3e4212ce} /* (4, 31, 13) {real, imag} */,
  {32'h3de14bda, 32'hbdd941ec} /* (4, 31, 12) {real, imag} */,
  {32'h3f3f87c2, 32'h3e8fe028} /* (4, 31, 11) {real, imag} */,
  {32'hbe2d9324, 32'h3f0bf683} /* (4, 31, 10) {real, imag} */,
  {32'hbe08855e, 32'hbd9f0d88} /* (4, 31, 9) {real, imag} */,
  {32'h3f3acac0, 32'h3ecb082a} /* (4, 31, 8) {real, imag} */,
  {32'hbf41b6c6, 32'h3dfe6a5a} /* (4, 31, 7) {real, imag} */,
  {32'h3ef6b5ca, 32'h3f0101b6} /* (4, 31, 6) {real, imag} */,
  {32'h404b796e, 32'hbe290a2e} /* (4, 31, 5) {real, imag} */,
  {32'hbfdeee70, 32'h400f469a} /* (4, 31, 4) {real, imag} */,
  {32'h3fc82ec2, 32'h3fa0f71e} /* (4, 31, 3) {real, imag} */,
  {32'h40a68dc8, 32'hbf7c72eb} /* (4, 31, 2) {real, imag} */,
  {32'hc1131668, 32'hbf1a93d0} /* (4, 31, 1) {real, imag} */,
  {32'hbf22e928, 32'hbfdfb30c} /* (4, 31, 0) {real, imag} */,
  {32'h4109ad3f, 32'hbd665600} /* (4, 30, 31) {real, imag} */,
  {32'hc0e31e4d, 32'hc0792c8a} /* (4, 30, 30) {real, imag} */,
  {32'hbefa7a2c, 32'hbe94b956} /* (4, 30, 29) {real, imag} */,
  {32'h4035abc9, 32'hbe2026fe} /* (4, 30, 28) {real, imag} */,
  {32'hbf271aba, 32'h3ff13038} /* (4, 30, 27) {real, imag} */,
  {32'h3eb8a4d6, 32'hbf0b1eda} /* (4, 30, 26) {real, imag} */,
  {32'h3f31302c, 32'h3e613a6d} /* (4, 30, 25) {real, imag} */,
  {32'hbf7238c7, 32'h3ec6e651} /* (4, 30, 24) {real, imag} */,
  {32'h3e3c9e98, 32'hbe1f63ce} /* (4, 30, 23) {real, imag} */,
  {32'h3e8ce546, 32'hbf2d22cf} /* (4, 30, 22) {real, imag} */,
  {32'hbe9bf068, 32'h3eac79e1} /* (4, 30, 21) {real, imag} */,
  {32'h3eb47e97, 32'hbe9c15f8} /* (4, 30, 20) {real, imag} */,
  {32'hbe3d1688, 32'h3e0bf04b} /* (4, 30, 19) {real, imag} */,
  {32'hbe18bb90, 32'h3f1c22a7} /* (4, 30, 18) {real, imag} */,
  {32'h3e1adc31, 32'hbebaa487} /* (4, 30, 17) {real, imag} */,
  {32'h3e66aef0, 32'h3e52a889} /* (4, 30, 16) {real, imag} */,
  {32'hbd236e56, 32'h3f0d98d2} /* (4, 30, 15) {real, imag} */,
  {32'h3e1776e0, 32'hbde90e34} /* (4, 30, 14) {real, imag} */,
  {32'hbde67f96, 32'h3e8bb15a} /* (4, 30, 13) {real, imag} */,
  {32'h3ea518f8, 32'h3de16509} /* (4, 30, 12) {real, imag} */,
  {32'hbea76fd4, 32'hbf2028fa} /* (4, 30, 11) {real, imag} */,
  {32'h3c80fd80, 32'hbea4ad02} /* (4, 30, 10) {real, imag} */,
  {32'hbea2c4dc, 32'hbe227409} /* (4, 30, 9) {real, imag} */,
  {32'hbea1c3ec, 32'hbffee26a} /* (4, 30, 8) {real, imag} */,
  {32'h3e8819cc, 32'h3f8ac40f} /* (4, 30, 7) {real, imag} */,
  {32'hbf5336de, 32'hbf7f7bee} /* (4, 30, 6) {real, imag} */,
  {32'hbfc77ed0, 32'hbf27ce8e} /* (4, 30, 5) {real, imag} */,
  {32'h3e9b3a96, 32'h400ba956} /* (4, 30, 4) {real, imag} */,
  {32'h3cf6fe20, 32'hbf74cdb0} /* (4, 30, 3) {real, imag} */,
  {32'hc0ed9e45, 32'hbfcbfea8} /* (4, 30, 2) {real, imag} */,
  {32'h416ccb8f, 32'hbf609371} /* (4, 30, 1) {real, imag} */,
  {32'h40af23e6, 32'hbe8f84c4} /* (4, 30, 0) {real, imag} */,
  {32'hc0178967, 32'hbea990d8} /* (4, 29, 31) {real, imag} */,
  {32'h3edb17d7, 32'hc0613b1e} /* (4, 29, 30) {real, imag} */,
  {32'hbe8f8a99, 32'h3f0e8801} /* (4, 29, 29) {real, imag} */,
  {32'h3f550140, 32'h3f3e00e3} /* (4, 29, 28) {real, imag} */,
  {32'hbf5aba0f, 32'h3e9c7bec} /* (4, 29, 27) {real, imag} */,
  {32'h3be85580, 32'h3ea6a326} /* (4, 29, 26) {real, imag} */,
  {32'hbe11466c, 32'h3f78531c} /* (4, 29, 25) {real, imag} */,
  {32'h3cd52ca8, 32'hbee70325} /* (4, 29, 24) {real, imag} */,
  {32'hbe2a23b5, 32'h3dd2ad2c} /* (4, 29, 23) {real, imag} */,
  {32'h3d145574, 32'h3e0afe0c} /* (4, 29, 22) {real, imag} */,
  {32'hbef04451, 32'h3e04d772} /* (4, 29, 21) {real, imag} */,
  {32'h3e9e4222, 32'h3e9d30db} /* (4, 29, 20) {real, imag} */,
  {32'h3e9d5c2e, 32'hbdccbda8} /* (4, 29, 19) {real, imag} */,
  {32'hbd358f34, 32'hbed2fef7} /* (4, 29, 18) {real, imag} */,
  {32'h3e16a47c, 32'hbc0ec6a8} /* (4, 29, 17) {real, imag} */,
  {32'h3e9a36fe, 32'h3ea8093b} /* (4, 29, 16) {real, imag} */,
  {32'h3e9d0c24, 32'hbdb7d1b9} /* (4, 29, 15) {real, imag} */,
  {32'hbf16f64a, 32'h3de31ac6} /* (4, 29, 14) {real, imag} */,
  {32'hbe79d999, 32'h3e517123} /* (4, 29, 13) {real, imag} */,
  {32'h3d4ae430, 32'h3bc9e8f4} /* (4, 29, 12) {real, imag} */,
  {32'hbea73458, 32'h3e7a333c} /* (4, 29, 11) {real, imag} */,
  {32'h3eb01c06, 32'h3efbac9d} /* (4, 29, 10) {real, imag} */,
  {32'hbe20fa2c, 32'h3f179d86} /* (4, 29, 9) {real, imag} */,
  {32'h3df8f89e, 32'hbf32c1a8} /* (4, 29, 8) {real, imag} */,
  {32'hbe79a733, 32'hbed1590e} /* (4, 29, 7) {real, imag} */,
  {32'hbe7d5344, 32'h3eebf55c} /* (4, 29, 6) {real, imag} */,
  {32'h3f817646, 32'h3f449091} /* (4, 29, 5) {real, imag} */,
  {32'hbf4b52c6, 32'h3eb8f8bd} /* (4, 29, 4) {real, imag} */,
  {32'hbc756a00, 32'hbe8f23ed} /* (4, 29, 3) {real, imag} */,
  {32'hbfbae113, 32'hbf8d1e00} /* (4, 29, 2) {real, imag} */,
  {32'h40289fe7, 32'h3fd97180} /* (4, 29, 1) {real, imag} */,
  {32'h3ed3a6a1, 32'hbf4cb1aa} /* (4, 29, 0) {real, imag} */,
  {32'hc098991c, 32'h3fc626ac} /* (4, 28, 31) {real, imag} */,
  {32'h40321df1, 32'hbfc393a6} /* (4, 28, 30) {real, imag} */,
  {32'hbf1e1673, 32'hbf659480} /* (4, 28, 29) {real, imag} */,
  {32'h3f3820bc, 32'h3f075424} /* (4, 28, 28) {real, imag} */,
  {32'h3f274907, 32'h3e3dd40c} /* (4, 28, 27) {real, imag} */,
  {32'h3ddecf00, 32'h3eac1a5e} /* (4, 28, 26) {real, imag} */,
  {32'hbf256632, 32'hbe51664a} /* (4, 28, 25) {real, imag} */,
  {32'h3db48c1a, 32'hbe8dd106} /* (4, 28, 24) {real, imag} */,
  {32'hbc7ef2d0, 32'hbed6adb8} /* (4, 28, 23) {real, imag} */,
  {32'h3ec4f75c, 32'h3ed9ae4a} /* (4, 28, 22) {real, imag} */,
  {32'hbc5fd01c, 32'h3ea8f18f} /* (4, 28, 21) {real, imag} */,
  {32'hbca8b274, 32'h3c6ca9c0} /* (4, 28, 20) {real, imag} */,
  {32'hbe0385e5, 32'h3d9add16} /* (4, 28, 19) {real, imag} */,
  {32'hbdc79f21, 32'hbed15276} /* (4, 28, 18) {real, imag} */,
  {32'hbe7b58e8, 32'h3d274958} /* (4, 28, 17) {real, imag} */,
  {32'hbe4f493b, 32'h3e7d1e16} /* (4, 28, 16) {real, imag} */,
  {32'hbdbe688e, 32'hbebb3a58} /* (4, 28, 15) {real, imag} */,
  {32'h3b0bd940, 32'hbe54eab6} /* (4, 28, 14) {real, imag} */,
  {32'h3e57c127, 32'h3e2afcbc} /* (4, 28, 13) {real, imag} */,
  {32'hbe11bdc4, 32'hbe09679a} /* (4, 28, 12) {real, imag} */,
  {32'h3f72c0ca, 32'h3e7dac7d} /* (4, 28, 11) {real, imag} */,
  {32'h3eadcdbb, 32'h3dd7924f} /* (4, 28, 10) {real, imag} */,
  {32'h3d2460c8, 32'hbdfec0db} /* (4, 28, 9) {real, imag} */,
  {32'h3e96f687, 32'h3c375778} /* (4, 28, 8) {real, imag} */,
  {32'h3e93b0b0, 32'hbb89ec20} /* (4, 28, 7) {real, imag} */,
  {32'hbfa3cb80, 32'h3eb98b2c} /* (4, 28, 6) {real, imag} */,
  {32'h3d2a71c2, 32'h3eec7ef0} /* (4, 28, 5) {real, imag} */,
  {32'hbf0fc2ba, 32'hbe73c6e3} /* (4, 28, 4) {real, imag} */,
  {32'hbe483d1a, 32'hbe72d4fc} /* (4, 28, 3) {real, imag} */,
  {32'h3fa91cb5, 32'hc039daec} /* (4, 28, 2) {real, imag} */,
  {32'hbfa23b39, 32'h4024f48e} /* (4, 28, 1) {real, imag} */,
  {32'hbfb7cfd6, 32'h3ea04cc8} /* (4, 28, 0) {real, imag} */,
  {32'h40247c5e, 32'hbfa17a40} /* (4, 27, 31) {real, imag} */,
  {32'h3e79080c, 32'hbf462afb} /* (4, 27, 30) {real, imag} */,
  {32'h3f28b277, 32'hbde41184} /* (4, 27, 29) {real, imag} */,
  {32'h3f0ac180, 32'h3e732361} /* (4, 27, 28) {real, imag} */,
  {32'hbf4d0fde, 32'h3f75e207} /* (4, 27, 27) {real, imag} */,
  {32'hbeaa11f4, 32'h3edaaea5} /* (4, 27, 26) {real, imag} */,
  {32'hbd14a736, 32'hbe1b60f2} /* (4, 27, 25) {real, imag} */,
  {32'h3dcc4244, 32'h3dc8e5ae} /* (4, 27, 24) {real, imag} */,
  {32'hbc57a1f0, 32'hbd33ff90} /* (4, 27, 23) {real, imag} */,
  {32'h3e5bab23, 32'hbf0dbbd8} /* (4, 27, 22) {real, imag} */,
  {32'hbdd5cc9e, 32'h3f522e0e} /* (4, 27, 21) {real, imag} */,
  {32'hbe184681, 32'hbdcbee1c} /* (4, 27, 20) {real, imag} */,
  {32'hbdd0a042, 32'h3eaa4d8f} /* (4, 27, 19) {real, imag} */,
  {32'h3eaa229e, 32'h3e5f34f4} /* (4, 27, 18) {real, imag} */,
  {32'h3e691b94, 32'h3e248f20} /* (4, 27, 17) {real, imag} */,
  {32'hbd87ff72, 32'hbe824680} /* (4, 27, 16) {real, imag} */,
  {32'hbe61e64c, 32'hbe74062e} /* (4, 27, 15) {real, imag} */,
  {32'h3eafd40e, 32'hbe60cafe} /* (4, 27, 14) {real, imag} */,
  {32'hbeba10a6, 32'hbd254dc0} /* (4, 27, 13) {real, imag} */,
  {32'hbe6de98c, 32'hbe0eaf0e} /* (4, 27, 12) {real, imag} */,
  {32'hbe8a65c0, 32'hbf6962b4} /* (4, 27, 11) {real, imag} */,
  {32'hbd876fa0, 32'hbc95ce48} /* (4, 27, 10) {real, imag} */,
  {32'h3e35de95, 32'h3ee10bf2} /* (4, 27, 9) {real, imag} */,
  {32'hbe8a68f8, 32'h3d4bb67e} /* (4, 27, 8) {real, imag} */,
  {32'h3f445c7e, 32'hbea7cbc8} /* (4, 27, 7) {real, imag} */,
  {32'hbe9a5dea, 32'hbea95625} /* (4, 27, 6) {real, imag} */,
  {32'hbf2819a3, 32'h3e199575} /* (4, 27, 5) {real, imag} */,
  {32'h3f3a9428, 32'h3f2f9882} /* (4, 27, 4) {real, imag} */,
  {32'hbdbb7eaa, 32'h3ebb7e25} /* (4, 27, 3) {real, imag} */,
  {32'hbfafeab3, 32'h3ecd9c0a} /* (4, 27, 2) {real, imag} */,
  {32'h3fda6421, 32'hbf324c80} /* (4, 27, 1) {real, imag} */,
  {32'h4023bf55, 32'h3e32cd1c} /* (4, 27, 0) {real, imag} */,
  {32'h3f08b211, 32'hbec4fc49} /* (4, 26, 31) {real, imag} */,
  {32'hbf2e8ad9, 32'h3e091fca} /* (4, 26, 30) {real, imag} */,
  {32'hbeb4a0be, 32'hbe4159b7} /* (4, 26, 29) {real, imag} */,
  {32'hbe39af60, 32'h3e9a5db0} /* (4, 26, 28) {real, imag} */,
  {32'hbe1d9fa9, 32'hbe41d63a} /* (4, 26, 27) {real, imag} */,
  {32'hbf22dcb0, 32'h3e9ad7a4} /* (4, 26, 26) {real, imag} */,
  {32'h3ea255d4, 32'hbeb40a5b} /* (4, 26, 25) {real, imag} */,
  {32'hbf2af1fe, 32'h3cc8a370} /* (4, 26, 24) {real, imag} */,
  {32'h3e4f6151, 32'h3cb19528} /* (4, 26, 23) {real, imag} */,
  {32'h3cbc4608, 32'h3dc93292} /* (4, 26, 22) {real, imag} */,
  {32'hbecd18c7, 32'hbe54a510} /* (4, 26, 21) {real, imag} */,
  {32'h3e6cc65e, 32'hbde58426} /* (4, 26, 20) {real, imag} */,
  {32'h3f00fb91, 32'h3dfe01a6} /* (4, 26, 19) {real, imag} */,
  {32'hbd4d22e8, 32'h3ec5f147} /* (4, 26, 18) {real, imag} */,
  {32'hbc5222a8, 32'hbd87ce34} /* (4, 26, 17) {real, imag} */,
  {32'h3d8cfa67, 32'h3e15ce90} /* (4, 26, 16) {real, imag} */,
  {32'h3e72f80c, 32'h3da8b098} /* (4, 26, 15) {real, imag} */,
  {32'h3df843ba, 32'hbcb136bc} /* (4, 26, 14) {real, imag} */,
  {32'hbe469ca9, 32'h3e112fe4} /* (4, 26, 13) {real, imag} */,
  {32'hbf29831d, 32'hbe513631} /* (4, 26, 12) {real, imag} */,
  {32'hbe76a4e3, 32'h3f20ff26} /* (4, 26, 11) {real, imag} */,
  {32'hbe068bab, 32'hbf036a8e} /* (4, 26, 10) {real, imag} */,
  {32'hbeeb0d7a, 32'h3e18251d} /* (4, 26, 9) {real, imag} */,
  {32'hbe892ce3, 32'hbec74fc6} /* (4, 26, 8) {real, imag} */,
  {32'hbcc943f4, 32'h3e925770} /* (4, 26, 7) {real, imag} */,
  {32'hbd5e71a8, 32'h3e6cfeaa} /* (4, 26, 6) {real, imag} */,
  {32'h3d300010, 32'hbf1e2a76} /* (4, 26, 5) {real, imag} */,
  {32'h3d8c20e0, 32'h3d083090} /* (4, 26, 4) {real, imag} */,
  {32'h3f32089d, 32'hbcb828b0} /* (4, 26, 3) {real, imag} */,
  {32'h3edb9333, 32'hbc4951e0} /* (4, 26, 2) {real, imag} */,
  {32'h3f0566bc, 32'hbf271802} /* (4, 26, 1) {real, imag} */,
  {32'h3ed1757b, 32'h3f126d0f} /* (4, 26, 0) {real, imag} */,
  {32'h3ba29c00, 32'h3f5e5ed0} /* (4, 25, 31) {real, imag} */,
  {32'h3f16639d, 32'hbea53c32} /* (4, 25, 30) {real, imag} */,
  {32'hbbf6f0c0, 32'hbe867624} /* (4, 25, 29) {real, imag} */,
  {32'hbeedb3c9, 32'h3ec112b2} /* (4, 25, 28) {real, imag} */,
  {32'h3f89f01a, 32'hbf463306} /* (4, 25, 27) {real, imag} */,
  {32'h3e9e4c54, 32'hbdacc3eb} /* (4, 25, 26) {real, imag} */,
  {32'hbf188057, 32'hbe9e5b11} /* (4, 25, 25) {real, imag} */,
  {32'h3e2e003e, 32'h3cf75d50} /* (4, 25, 24) {real, imag} */,
  {32'h3eab1276, 32'hbdbbbd5c} /* (4, 25, 23) {real, imag} */,
  {32'h3e270dfa, 32'h3e4a626a} /* (4, 25, 22) {real, imag} */,
  {32'hbe2e9a42, 32'hbeb57e0f} /* (4, 25, 21) {real, imag} */,
  {32'hbf2de3e2, 32'hbda93420} /* (4, 25, 20) {real, imag} */,
  {32'hbf1e20eb, 32'hbeb0b5a8} /* (4, 25, 19) {real, imag} */,
  {32'hbef14e8a, 32'h3ccad230} /* (4, 25, 18) {real, imag} */,
  {32'hbee01659, 32'h3f0135a8} /* (4, 25, 17) {real, imag} */,
  {32'h3ed9987f, 32'h3dea32b2} /* (4, 25, 16) {real, imag} */,
  {32'hbce03174, 32'hbea19cce} /* (4, 25, 15) {real, imag} */,
  {32'h3efa3896, 32'h3e55b06f} /* (4, 25, 14) {real, imag} */,
  {32'hbe506284, 32'hbef64ad2} /* (4, 25, 13) {real, imag} */,
  {32'h3e9cd558, 32'h3e234132} /* (4, 25, 12) {real, imag} */,
  {32'hbe22fec1, 32'hbf007f1a} /* (4, 25, 11) {real, imag} */,
  {32'hbd6918f8, 32'h3ea5e41c} /* (4, 25, 10) {real, imag} */,
  {32'hbd3d584e, 32'hbed32650} /* (4, 25, 9) {real, imag} */,
  {32'hbed37006, 32'h3f11a78a} /* (4, 25, 8) {real, imag} */,
  {32'h3df8483a, 32'h3e3d772a} /* (4, 25, 7) {real, imag} */,
  {32'h3eae43f3, 32'h3e6014c9} /* (4, 25, 6) {real, imag} */,
  {32'h3f2061da, 32'hbe5c7b8c} /* (4, 25, 5) {real, imag} */,
  {32'hbf0f8df0, 32'h3f3938dc} /* (4, 25, 4) {real, imag} */,
  {32'hbe950396, 32'h3eb57b46} /* (4, 25, 3) {real, imag} */,
  {32'hbe18814a, 32'hbf5ac3cc} /* (4, 25, 2) {real, imag} */,
  {32'hbf5c7086, 32'h3cb7d3cc} /* (4, 25, 1) {real, imag} */,
  {32'hbf46088a, 32'h3e9a5c4a} /* (4, 25, 0) {real, imag} */,
  {32'hbd71f918, 32'hbee5830c} /* (4, 24, 31) {real, imag} */,
  {32'hbf286cd2, 32'h3f10e353} /* (4, 24, 30) {real, imag} */,
  {32'hbd431862, 32'hbd446f18} /* (4, 24, 29) {real, imag} */,
  {32'hbe065ddb, 32'h3d06cc7c} /* (4, 24, 28) {real, imag} */,
  {32'hbc0eb100, 32'h3f0d97ea} /* (4, 24, 27) {real, imag} */,
  {32'hbe48d5a6, 32'hbec9d87e} /* (4, 24, 26) {real, imag} */,
  {32'hbe340eec, 32'hbda7aa38} /* (4, 24, 25) {real, imag} */,
  {32'hbe8a4634, 32'hbe6baaee} /* (4, 24, 24) {real, imag} */,
  {32'h3eccecfc, 32'hbf1ba022} /* (4, 24, 23) {real, imag} */,
  {32'h3f0e1ac9, 32'h3d60d3f0} /* (4, 24, 22) {real, imag} */,
  {32'hbe84945a, 32'h39f0ea00} /* (4, 24, 21) {real, imag} */,
  {32'hbddcd5b1, 32'hbe0f38d0} /* (4, 24, 20) {real, imag} */,
  {32'h3e35ac29, 32'h3edccfc0} /* (4, 24, 19) {real, imag} */,
  {32'h3e885a50, 32'hbf09a7e1} /* (4, 24, 18) {real, imag} */,
  {32'hbd5e8f66, 32'h3c5d7da8} /* (4, 24, 17) {real, imag} */,
  {32'h3b99a478, 32'h3e8f44ca} /* (4, 24, 16) {real, imag} */,
  {32'h3e99801e, 32'hbdcfb8c2} /* (4, 24, 15) {real, imag} */,
  {32'h3dc06782, 32'hbd98b7ca} /* (4, 24, 14) {real, imag} */,
  {32'hbea4bbd2, 32'hbe97fa5e} /* (4, 24, 13) {real, imag} */,
  {32'h3ebf15fd, 32'h3ef5e13e} /* (4, 24, 12) {real, imag} */,
  {32'h3cfa9ac8, 32'hbed6ecc7} /* (4, 24, 11) {real, imag} */,
  {32'hbed1cd81, 32'hbea06be6} /* (4, 24, 10) {real, imag} */,
  {32'hbf24db44, 32'h3e880e71} /* (4, 24, 9) {real, imag} */,
  {32'hbf1d6e1d, 32'h3e2ba6a3} /* (4, 24, 8) {real, imag} */,
  {32'hbeb77614, 32'hbe2ac088} /* (4, 24, 7) {real, imag} */,
  {32'h3e56a198, 32'h3e9450e8} /* (4, 24, 6) {real, imag} */,
  {32'h3e5a4f68, 32'h3ecaa07c} /* (4, 24, 5) {real, imag} */,
  {32'h3edcc0f6, 32'h3db013d6} /* (4, 24, 4) {real, imag} */,
  {32'h3e1e0f20, 32'hbe5504e2} /* (4, 24, 3) {real, imag} */,
  {32'hbf8c18a4, 32'h3ec378a6} /* (4, 24, 2) {real, imag} */,
  {32'h3fbe96a6, 32'hbe8b7fcf} /* (4, 24, 1) {real, imag} */,
  {32'h3f2f95a3, 32'hbf892d0c} /* (4, 24, 0) {real, imag} */,
  {32'hbeea0e35, 32'h3e4d133a} /* (4, 23, 31) {real, imag} */,
  {32'h3d2c7528, 32'hbdbcf69b} /* (4, 23, 30) {real, imag} */,
  {32'h3eb8de7e, 32'hbf3dc7bc} /* (4, 23, 29) {real, imag} */,
  {32'h3d9deec0, 32'h3eebca74} /* (4, 23, 28) {real, imag} */,
  {32'hbdf974ac, 32'h3e9b95cb} /* (4, 23, 27) {real, imag} */,
  {32'hbd7954a6, 32'hbe834225} /* (4, 23, 26) {real, imag} */,
  {32'h3dd05204, 32'hbe14f5f6} /* (4, 23, 25) {real, imag} */,
  {32'hbd969ac7, 32'h3b8840c0} /* (4, 23, 24) {real, imag} */,
  {32'hbe745db9, 32'hbe12ba80} /* (4, 23, 23) {real, imag} */,
  {32'h3ee0bf4a, 32'h3ef882b2} /* (4, 23, 22) {real, imag} */,
  {32'hbee3b1f2, 32'h3e9cfedb} /* (4, 23, 21) {real, imag} */,
  {32'hbdaf059b, 32'h3eef5fd4} /* (4, 23, 20) {real, imag} */,
  {32'hbde8e66c, 32'hbbe52670} /* (4, 23, 19) {real, imag} */,
  {32'hbe1cbca8, 32'h3d6bb618} /* (4, 23, 18) {real, imag} */,
  {32'hbd81b6be, 32'h3e0684ca} /* (4, 23, 17) {real, imag} */,
  {32'hbebb66d0, 32'h3f062175} /* (4, 23, 16) {real, imag} */,
  {32'h3e0d9339, 32'hbe6942b7} /* (4, 23, 15) {real, imag} */,
  {32'hbe0b90d4, 32'hbe7c0f7f} /* (4, 23, 14) {real, imag} */,
  {32'hbf1d4502, 32'hbd5d1250} /* (4, 23, 13) {real, imag} */,
  {32'h3e6ca350, 32'hbf12c51f} /* (4, 23, 12) {real, imag} */,
  {32'hbe0a4ea4, 32'h3ebc2587} /* (4, 23, 11) {real, imag} */,
  {32'hbe3c7260, 32'h3ef998b5} /* (4, 23, 10) {real, imag} */,
  {32'hbee0d8c3, 32'h3f3468e2} /* (4, 23, 9) {real, imag} */,
  {32'hbe00a85d, 32'hbe0702c8} /* (4, 23, 8) {real, imag} */,
  {32'hbe55a559, 32'hbedf8cf1} /* (4, 23, 7) {real, imag} */,
  {32'h3f28c2ad, 32'hbd81ea50} /* (4, 23, 6) {real, imag} */,
  {32'h3f31bbc6, 32'hbf01be5f} /* (4, 23, 5) {real, imag} */,
  {32'h3e02b1e6, 32'h3e6508a4} /* (4, 23, 4) {real, imag} */,
  {32'hbdf576c4, 32'h3ed560b5} /* (4, 23, 3) {real, imag} */,
  {32'h3dc8b4a4, 32'h3d5a6310} /* (4, 23, 2) {real, imag} */,
  {32'h3e8b6442, 32'h3cf435d0} /* (4, 23, 1) {real, imag} */,
  {32'hbe2ce468, 32'hbef4ddbd} /* (4, 23, 0) {real, imag} */,
  {32'hbed97c3b, 32'h3d288c3e} /* (4, 22, 31) {real, imag} */,
  {32'h3f1c9715, 32'hbe9a3eb5} /* (4, 22, 30) {real, imag} */,
  {32'hbe599177, 32'h3e70a243} /* (4, 22, 29) {real, imag} */,
  {32'hbd10d1b0, 32'h3e6468db} /* (4, 22, 28) {real, imag} */,
  {32'h3e8ae95b, 32'h3f164c3e} /* (4, 22, 27) {real, imag} */,
  {32'h3f0101bf, 32'hbeba6e1c} /* (4, 22, 26) {real, imag} */,
  {32'hbeacfcfa, 32'hbe8abef6} /* (4, 22, 25) {real, imag} */,
  {32'hbe8be33c, 32'hbe834964} /* (4, 22, 24) {real, imag} */,
  {32'hbc29cb40, 32'hbeefd94e} /* (4, 22, 23) {real, imag} */,
  {32'h3e9c961c, 32'h3e91d848} /* (4, 22, 22) {real, imag} */,
  {32'h3f24c715, 32'hbe75e8d0} /* (4, 22, 21) {real, imag} */,
  {32'h3f18d087, 32'h3e541000} /* (4, 22, 20) {real, imag} */,
  {32'hbd7d0e64, 32'hbe4a823c} /* (4, 22, 19) {real, imag} */,
  {32'hbe2b5cd8, 32'hbe6eacd3} /* (4, 22, 18) {real, imag} */,
  {32'h3e0e69dd, 32'h3e0bf8c9} /* (4, 22, 17) {real, imag} */,
  {32'h3d950843, 32'hbecd3674} /* (4, 22, 16) {real, imag} */,
  {32'h3d34f966, 32'hbe429718} /* (4, 22, 15) {real, imag} */,
  {32'hbd98bdc8, 32'hbe143618} /* (4, 22, 14) {real, imag} */,
  {32'hbd42e5b0, 32'hbd81ef3a} /* (4, 22, 13) {real, imag} */,
  {32'h3ee3d019, 32'hbe38ee5a} /* (4, 22, 12) {real, imag} */,
  {32'hbe50fc34, 32'h3ece4c9a} /* (4, 22, 11) {real, imag} */,
  {32'hbe90e90c, 32'hbec90885} /* (4, 22, 10) {real, imag} */,
  {32'h3dcda5a8, 32'h3d35c26f} /* (4, 22, 9) {real, imag} */,
  {32'hbe94c565, 32'hbf36e4c9} /* (4, 22, 8) {real, imag} */,
  {32'hbe26dc0e, 32'h3e258dfe} /* (4, 22, 7) {real, imag} */,
  {32'h3e9f318c, 32'h3e4dbfd4} /* (4, 22, 6) {real, imag} */,
  {32'h3f42bee3, 32'hbedf7075} /* (4, 22, 5) {real, imag} */,
  {32'hbdc9591a, 32'hbd6b2b8c} /* (4, 22, 4) {real, imag} */,
  {32'hbf189a9f, 32'hbf223602} /* (4, 22, 3) {real, imag} */,
  {32'h3d21578a, 32'h3ea9f866} /* (4, 22, 2) {real, imag} */,
  {32'h3ef6bb58, 32'h3eb9fcc1} /* (4, 22, 1) {real, imag} */,
  {32'hbf03c667, 32'h3f292d22} /* (4, 22, 0) {real, imag} */,
  {32'hbd80a81a, 32'hbf9cb290} /* (4, 21, 31) {real, imag} */,
  {32'hbde18118, 32'h3edd7304} /* (4, 21, 30) {real, imag} */,
  {32'hbf35d760, 32'h3e37a610} /* (4, 21, 29) {real, imag} */,
  {32'hbd4eb084, 32'h3e98016b} /* (4, 21, 28) {real, imag} */,
  {32'hbec0be68, 32'hbdfc301c} /* (4, 21, 27) {real, imag} */,
  {32'h3f250f17, 32'hbe6324a2} /* (4, 21, 26) {real, imag} */,
  {32'h3eefe189, 32'hbbcdcc80} /* (4, 21, 25) {real, imag} */,
  {32'hbe86a89a, 32'h3dd365a8} /* (4, 21, 24) {real, imag} */,
  {32'hbeb61251, 32'hbe5591b2} /* (4, 21, 23) {real, imag} */,
  {32'hbea8364b, 32'hbdfd36ed} /* (4, 21, 22) {real, imag} */,
  {32'hbe9466bd, 32'h3ebf53b6} /* (4, 21, 21) {real, imag} */,
  {32'hbeddd17f, 32'h3e98d912} /* (4, 21, 20) {real, imag} */,
  {32'hbdf6f52d, 32'h3ea551cf} /* (4, 21, 19) {real, imag} */,
  {32'h3f21c805, 32'h3e141a42} /* (4, 21, 18) {real, imag} */,
  {32'hbc2ccc60, 32'hbe71afcc} /* (4, 21, 17) {real, imag} */,
  {32'h3e6cb998, 32'hbd9648f4} /* (4, 21, 16) {real, imag} */,
  {32'hbe286992, 32'h3ee7172c} /* (4, 21, 15) {real, imag} */,
  {32'hbed95252, 32'hbe7de3e4} /* (4, 21, 14) {real, imag} */,
  {32'hbda16326, 32'hbd80c008} /* (4, 21, 13) {real, imag} */,
  {32'h3e86405e, 32'h3de4a1c0} /* (4, 21, 12) {real, imag} */,
  {32'hbea8abac, 32'h3cf83dd8} /* (4, 21, 11) {real, imag} */,
  {32'hbe8a2ce6, 32'hbe9dcb7a} /* (4, 21, 10) {real, imag} */,
  {32'h3c8a7eac, 32'h3e9a53f4} /* (4, 21, 9) {real, imag} */,
  {32'hbe20a292, 32'hbe3e1d1a} /* (4, 21, 8) {real, imag} */,
  {32'h3e97809e, 32'hbd805c28} /* (4, 21, 7) {real, imag} */,
  {32'hbe41eb7a, 32'hbdfc5a1c} /* (4, 21, 6) {real, imag} */,
  {32'hbe0294f9, 32'h3ee8d502} /* (4, 21, 5) {real, imag} */,
  {32'h3e53e39a, 32'hbd7e3264} /* (4, 21, 4) {real, imag} */,
  {32'hbeef962b, 32'hbdfcf4a6} /* (4, 21, 3) {real, imag} */,
  {32'hbee50f46, 32'h3e904dd9} /* (4, 21, 2) {real, imag} */,
  {32'h3e7be16f, 32'hbf142e25} /* (4, 21, 1) {real, imag} */,
  {32'h3f8660cc, 32'hbe762072} /* (4, 21, 0) {real, imag} */,
  {32'h3dd9867b, 32'h3e577070} /* (4, 20, 31) {real, imag} */,
  {32'h3da535a3, 32'hbe345999} /* (4, 20, 30) {real, imag} */,
  {32'hbea6fb48, 32'h3e50cad7} /* (4, 20, 29) {real, imag} */,
  {32'hbe8eb760, 32'hbed9936b} /* (4, 20, 28) {real, imag} */,
  {32'h3e7cbcdc, 32'h3f36f8ff} /* (4, 20, 27) {real, imag} */,
  {32'h3e52346c, 32'hbe0a482a} /* (4, 20, 26) {real, imag} */,
  {32'h3e28c94b, 32'h3d031de0} /* (4, 20, 25) {real, imag} */,
  {32'h3edb36f0, 32'hbef6469d} /* (4, 20, 24) {real, imag} */,
  {32'h3ea34800, 32'hbdf32792} /* (4, 20, 23) {real, imag} */,
  {32'hbf160b06, 32'h3e2f4732} /* (4, 20, 22) {real, imag} */,
  {32'h3e0b461e, 32'h3db3efdf} /* (4, 20, 21) {real, imag} */,
  {32'h3ee8d0a4, 32'hbe95f91b} /* (4, 20, 20) {real, imag} */,
  {32'hbe331ccc, 32'hbe92a0fc} /* (4, 20, 19) {real, imag} */,
  {32'h3eb9f0cf, 32'hbdbb215c} /* (4, 20, 18) {real, imag} */,
  {32'hbf0d3e21, 32'hbddfc7d6} /* (4, 20, 17) {real, imag} */,
  {32'hbb46f680, 32'h3cebf288} /* (4, 20, 16) {real, imag} */,
  {32'h3ed59e90, 32'hbe18a8d2} /* (4, 20, 15) {real, imag} */,
  {32'h3e6cb76b, 32'hbe2bb938} /* (4, 20, 14) {real, imag} */,
  {32'h3f1c222a, 32'h3db256e8} /* (4, 20, 13) {real, imag} */,
  {32'hbe9566e1, 32'h3d3e69f4} /* (4, 20, 12) {real, imag} */,
  {32'h39016000, 32'hbf08e4d9} /* (4, 20, 11) {real, imag} */,
  {32'h3ef58f7e, 32'h3f3e8e2a} /* (4, 20, 10) {real, imag} */,
  {32'hbe9ddc40, 32'h3c8bfca0} /* (4, 20, 9) {real, imag} */,
  {32'h3e68b00e, 32'h3d3359f4} /* (4, 20, 8) {real, imag} */,
  {32'hbdc72cac, 32'h3f254263} /* (4, 20, 7) {real, imag} */,
  {32'hbef66a56, 32'h3e0d9a7e} /* (4, 20, 6) {real, imag} */,
  {32'h3e94ae47, 32'h3e2ffd42} /* (4, 20, 5) {real, imag} */,
  {32'h3e869960, 32'hbd8170a0} /* (4, 20, 4) {real, imag} */,
  {32'hbebf797f, 32'hbe366946} /* (4, 20, 3) {real, imag} */,
  {32'hbe8c0730, 32'hbeeb5854} /* (4, 20, 2) {real, imag} */,
  {32'hbe12be58, 32'hbde1b2b9} /* (4, 20, 1) {real, imag} */,
  {32'hbe80a0d0, 32'hbc03ff10} /* (4, 20, 0) {real, imag} */,
  {32'h3e91592d, 32'h3e9b3ebe} /* (4, 19, 31) {real, imag} */,
  {32'h3e45f5c0, 32'hbe9386b2} /* (4, 19, 30) {real, imag} */,
  {32'hbd8b7f01, 32'h3e572df0} /* (4, 19, 29) {real, imag} */,
  {32'hbe87b390, 32'h3e2b80d3} /* (4, 19, 28) {real, imag} */,
  {32'hbeb83d48, 32'hbe35f46f} /* (4, 19, 27) {real, imag} */,
  {32'hbe9a9d6b, 32'h3eed9c43} /* (4, 19, 26) {real, imag} */,
  {32'hbf0f7b47, 32'h3ed0524d} /* (4, 19, 25) {real, imag} */,
  {32'hbe005535, 32'hbf28e5b8} /* (4, 19, 24) {real, imag} */,
  {32'h3e94b8cc, 32'hbac65fc0} /* (4, 19, 23) {real, imag} */,
  {32'hbee302b2, 32'hbdd0da09} /* (4, 19, 22) {real, imag} */,
  {32'h3e31df36, 32'h3e20080a} /* (4, 19, 21) {real, imag} */,
  {32'h3e3d52d2, 32'hbe03ca20} /* (4, 19, 20) {real, imag} */,
  {32'hbe7dda77, 32'hbf1649ec} /* (4, 19, 19) {real, imag} */,
  {32'hbe443ee4, 32'hbd7aeee6} /* (4, 19, 18) {real, imag} */,
  {32'h3e9e907c, 32'h3f1a865a} /* (4, 19, 17) {real, imag} */,
  {32'h3dc0963c, 32'h3dc8b7de} /* (4, 19, 16) {real, imag} */,
  {32'hbe4b41bc, 32'h3e87c172} /* (4, 19, 15) {real, imag} */,
  {32'h3d23191c, 32'h3ead724b} /* (4, 19, 14) {real, imag} */,
  {32'hbeaf2e17, 32'h3d99b804} /* (4, 19, 13) {real, imag} */,
  {32'hbed8cec0, 32'h3e94864b} /* (4, 19, 12) {real, imag} */,
  {32'h3f20011e, 32'hbe260d2a} /* (4, 19, 11) {real, imag} */,
  {32'h3d0d87ea, 32'h3e91e0fb} /* (4, 19, 10) {real, imag} */,
  {32'hbed2ef3e, 32'hbf00729b} /* (4, 19, 9) {real, imag} */,
  {32'h3eb89654, 32'h3d2bfe5a} /* (4, 19, 8) {real, imag} */,
  {32'h3e209502, 32'hbeef0977} /* (4, 19, 7) {real, imag} */,
  {32'hbe8c9da8, 32'h3e3eee28} /* (4, 19, 6) {real, imag} */,
  {32'hbe2f39b6, 32'h3e8a70b6} /* (4, 19, 5) {real, imag} */,
  {32'h3c856927, 32'h3c9bd0c4} /* (4, 19, 4) {real, imag} */,
  {32'h3d8be66a, 32'h3ef76306} /* (4, 19, 3) {real, imag} */,
  {32'h3dfcea61, 32'hbcb68af6} /* (4, 19, 2) {real, imag} */,
  {32'hbee0b363, 32'h3e37e0a3} /* (4, 19, 1) {real, imag} */,
  {32'hbe433b5f, 32'hbe1027fc} /* (4, 19, 0) {real, imag} */,
  {32'hbf0a05a3, 32'h3e60aee1} /* (4, 18, 31) {real, imag} */,
  {32'hbdaaf6bd, 32'h3c0213c0} /* (4, 18, 30) {real, imag} */,
  {32'h3db8bb9c, 32'h3d68c250} /* (4, 18, 29) {real, imag} */,
  {32'h3e84afd4, 32'hbea5e6fa} /* (4, 18, 28) {real, imag} */,
  {32'h3dc71f62, 32'h3e1e4bd3} /* (4, 18, 27) {real, imag} */,
  {32'h3d578dca, 32'hbd02e044} /* (4, 18, 26) {real, imag} */,
  {32'hbe1d71e9, 32'h3ec6baf8} /* (4, 18, 25) {real, imag} */,
  {32'hbda6c327, 32'h3e6a7a70} /* (4, 18, 24) {real, imag} */,
  {32'h3f1e105c, 32'h3e8493b0} /* (4, 18, 23) {real, imag} */,
  {32'hbdfbd376, 32'h3de50202} /* (4, 18, 22) {real, imag} */,
  {32'h3d3a54bc, 32'hbed90d88} /* (4, 18, 21) {real, imag} */,
  {32'hbe157404, 32'h3e1ec32d} /* (4, 18, 20) {real, imag} */,
  {32'hbe4e4b89, 32'hbd2dfac0} /* (4, 18, 19) {real, imag} */,
  {32'hbd254628, 32'hbdd53c6d} /* (4, 18, 18) {real, imag} */,
  {32'hbeae5476, 32'h3d0adf76} /* (4, 18, 17) {real, imag} */,
  {32'hbd60d194, 32'h3dbe6cdf} /* (4, 18, 16) {real, imag} */,
  {32'h3dc4b6a1, 32'h3d908d10} /* (4, 18, 15) {real, imag} */,
  {32'h3d9ec598, 32'h3f0b9cac} /* (4, 18, 14) {real, imag} */,
  {32'hbeb4b0c8, 32'hbd84bc37} /* (4, 18, 13) {real, imag} */,
  {32'h3d733c53, 32'h3d0ab9f6} /* (4, 18, 12) {real, imag} */,
  {32'h3e6a2bc0, 32'hbee08db6} /* (4, 18, 11) {real, imag} */,
  {32'h3d448ec6, 32'hbcc29cbc} /* (4, 18, 10) {real, imag} */,
  {32'h3d735d00, 32'h3eb6083b} /* (4, 18, 9) {real, imag} */,
  {32'h3e82b6af, 32'hbe37f8ff} /* (4, 18, 8) {real, imag} */,
  {32'h3e0baa91, 32'hbb8d7200} /* (4, 18, 7) {real, imag} */,
  {32'hbe28bfca, 32'hbe981029} /* (4, 18, 6) {real, imag} */,
  {32'h3e20ec51, 32'h3ecb2452} /* (4, 18, 5) {real, imag} */,
  {32'hbe6a904e, 32'hbd20bdac} /* (4, 18, 4) {real, imag} */,
  {32'h3e520597, 32'h3eefc10b} /* (4, 18, 3) {real, imag} */,
  {32'hbe13a2fb, 32'h3c8aa980} /* (4, 18, 2) {real, imag} */,
  {32'h3ebde1f4, 32'hbed57bf3} /* (4, 18, 1) {real, imag} */,
  {32'h3ca9b15e, 32'hbe5edb95} /* (4, 18, 0) {real, imag} */,
  {32'hbe4e915e, 32'h3eaad585} /* (4, 17, 31) {real, imag} */,
  {32'hbe1e7fbf, 32'hbeb20965} /* (4, 17, 30) {real, imag} */,
  {32'h3e8b052b, 32'h3e8388e3} /* (4, 17, 29) {real, imag} */,
  {32'h3e55bcfd, 32'h3d3ce4e8} /* (4, 17, 28) {real, imag} */,
  {32'hbf10df56, 32'hbbad5d40} /* (4, 17, 27) {real, imag} */,
  {32'h3e4202ed, 32'h3d6b4678} /* (4, 17, 26) {real, imag} */,
  {32'h3c03eda0, 32'hbc8a4d10} /* (4, 17, 25) {real, imag} */,
  {32'hbdced95c, 32'hbdafb7ec} /* (4, 17, 24) {real, imag} */,
  {32'h3ec5e632, 32'h3e9853f9} /* (4, 17, 23) {real, imag} */,
  {32'hbccc1b28, 32'hbca54784} /* (4, 17, 22) {real, imag} */,
  {32'hbdcd0397, 32'h3e92d95f} /* (4, 17, 21) {real, imag} */,
  {32'h3e4216bc, 32'hbc2571e8} /* (4, 17, 20) {real, imag} */,
  {32'h3eba046b, 32'h3df0409d} /* (4, 17, 19) {real, imag} */,
  {32'hbe73638c, 32'h3ea6615b} /* (4, 17, 18) {real, imag} */,
  {32'h3d65a899, 32'hbeaee702} /* (4, 17, 17) {real, imag} */,
  {32'h3e5385fb, 32'h3d76b002} /* (4, 17, 16) {real, imag} */,
  {32'hbe70028f, 32'hbd878ec2} /* (4, 17, 15) {real, imag} */,
  {32'h3ea29559, 32'hbe2cea4b} /* (4, 17, 14) {real, imag} */,
  {32'h3ee2ad1a, 32'hbead88ec} /* (4, 17, 13) {real, imag} */,
  {32'h3eb81c9f, 32'hbe096874} /* (4, 17, 12) {real, imag} */,
  {32'hbe175db5, 32'hbe87388f} /* (4, 17, 11) {real, imag} */,
  {32'hbea76710, 32'h3e64d1de} /* (4, 17, 10) {real, imag} */,
  {32'hbe1b4556, 32'h3e858ba0} /* (4, 17, 9) {real, imag} */,
  {32'hbe476142, 32'h3c70f058} /* (4, 17, 8) {real, imag} */,
  {32'h3d80417a, 32'h3e9a65e8} /* (4, 17, 7) {real, imag} */,
  {32'h3eb4265a, 32'h3e4de41e} /* (4, 17, 6) {real, imag} */,
  {32'h3e0f970e, 32'h3deffe47} /* (4, 17, 5) {real, imag} */,
  {32'hbe0b4a0f, 32'hbcdf786a} /* (4, 17, 4) {real, imag} */,
  {32'hbe2da9ab, 32'hbe6b0174} /* (4, 17, 3) {real, imag} */,
  {32'hbde232dc, 32'hbdaafca2} /* (4, 17, 2) {real, imag} */,
  {32'h3ded84ea, 32'h3ef30ca4} /* (4, 17, 1) {real, imag} */,
  {32'hbe009e79, 32'h3f22b519} /* (4, 17, 0) {real, imag} */,
  {32'hbe5b38cf, 32'hbe761d66} /* (4, 16, 31) {real, imag} */,
  {32'hbe423126, 32'hbd6881d1} /* (4, 16, 30) {real, imag} */,
  {32'hbe2f5818, 32'hbcd2d4c8} /* (4, 16, 29) {real, imag} */,
  {32'h3e496e2b, 32'hbe967279} /* (4, 16, 28) {real, imag} */,
  {32'h3e6262ac, 32'hbe8d45fb} /* (4, 16, 27) {real, imag} */,
  {32'h3d4fb3e2, 32'h3c4603a0} /* (4, 16, 26) {real, imag} */,
  {32'hbde635f8, 32'hbed0ec38} /* (4, 16, 25) {real, imag} */,
  {32'h3ddb328b, 32'hbe1227fa} /* (4, 16, 24) {real, imag} */,
  {32'hbcfe2158, 32'h3d88556e} /* (4, 16, 23) {real, imag} */,
  {32'hbea95421, 32'hbebf21c7} /* (4, 16, 22) {real, imag} */,
  {32'hbe81bf54, 32'hbd805d54} /* (4, 16, 21) {real, imag} */,
  {32'h3dc5a84b, 32'hbdf1e326} /* (4, 16, 20) {real, imag} */,
  {32'h3e016963, 32'hbe4eb01b} /* (4, 16, 19) {real, imag} */,
  {32'hbe6cf7f7, 32'hbd3073a4} /* (4, 16, 18) {real, imag} */,
  {32'hb8e8f000, 32'hbd68c78a} /* (4, 16, 17) {real, imag} */,
  {32'hbdc0580e, 32'h00000000} /* (4, 16, 16) {real, imag} */,
  {32'hb8e8f000, 32'h3d68c78a} /* (4, 16, 15) {real, imag} */,
  {32'hbe6cf7f7, 32'h3d3073a4} /* (4, 16, 14) {real, imag} */,
  {32'h3e016963, 32'h3e4eb01b} /* (4, 16, 13) {real, imag} */,
  {32'h3dc5a84b, 32'h3df1e326} /* (4, 16, 12) {real, imag} */,
  {32'hbe81bf54, 32'h3d805d54} /* (4, 16, 11) {real, imag} */,
  {32'hbea95421, 32'h3ebf21c7} /* (4, 16, 10) {real, imag} */,
  {32'hbcfe2158, 32'hbd88556e} /* (4, 16, 9) {real, imag} */,
  {32'h3ddb328b, 32'h3e1227fa} /* (4, 16, 8) {real, imag} */,
  {32'hbde635f8, 32'h3ed0ec38} /* (4, 16, 7) {real, imag} */,
  {32'h3d4fb3e2, 32'hbc4603a0} /* (4, 16, 6) {real, imag} */,
  {32'h3e6262ac, 32'h3e8d45fb} /* (4, 16, 5) {real, imag} */,
  {32'h3e496e2b, 32'h3e967279} /* (4, 16, 4) {real, imag} */,
  {32'hbe2f5818, 32'h3cd2d4c8} /* (4, 16, 3) {real, imag} */,
  {32'hbe423126, 32'h3d6881d1} /* (4, 16, 2) {real, imag} */,
  {32'hbe5b38cf, 32'h3e761d66} /* (4, 16, 1) {real, imag} */,
  {32'h3d9871fc, 32'h00000000} /* (4, 16, 0) {real, imag} */,
  {32'h3ded84ea, 32'hbef30ca4} /* (4, 15, 31) {real, imag} */,
  {32'hbde232dc, 32'h3daafca2} /* (4, 15, 30) {real, imag} */,
  {32'hbe2da9ab, 32'h3e6b0174} /* (4, 15, 29) {real, imag} */,
  {32'hbe0b4a0f, 32'h3cdf786a} /* (4, 15, 28) {real, imag} */,
  {32'h3e0f970e, 32'hbdeffe47} /* (4, 15, 27) {real, imag} */,
  {32'h3eb4265a, 32'hbe4de41e} /* (4, 15, 26) {real, imag} */,
  {32'h3d80417a, 32'hbe9a65e8} /* (4, 15, 25) {real, imag} */,
  {32'hbe476142, 32'hbc70f058} /* (4, 15, 24) {real, imag} */,
  {32'hbe1b4556, 32'hbe858ba0} /* (4, 15, 23) {real, imag} */,
  {32'hbea76710, 32'hbe64d1de} /* (4, 15, 22) {real, imag} */,
  {32'hbe175db5, 32'h3e87388f} /* (4, 15, 21) {real, imag} */,
  {32'h3eb81c9f, 32'h3e096874} /* (4, 15, 20) {real, imag} */,
  {32'h3ee2ad1a, 32'h3ead88ec} /* (4, 15, 19) {real, imag} */,
  {32'h3ea29559, 32'h3e2cea4b} /* (4, 15, 18) {real, imag} */,
  {32'hbe70028f, 32'h3d878ec2} /* (4, 15, 17) {real, imag} */,
  {32'h3e5385fb, 32'hbd76b002} /* (4, 15, 16) {real, imag} */,
  {32'h3d65a899, 32'h3eaee702} /* (4, 15, 15) {real, imag} */,
  {32'hbe73638c, 32'hbea6615b} /* (4, 15, 14) {real, imag} */,
  {32'h3eba046b, 32'hbdf0409d} /* (4, 15, 13) {real, imag} */,
  {32'h3e4216bc, 32'h3c2571e8} /* (4, 15, 12) {real, imag} */,
  {32'hbdcd0397, 32'hbe92d95f} /* (4, 15, 11) {real, imag} */,
  {32'hbccc1b28, 32'h3ca54784} /* (4, 15, 10) {real, imag} */,
  {32'h3ec5e632, 32'hbe9853f9} /* (4, 15, 9) {real, imag} */,
  {32'hbdced95c, 32'h3dafb7ec} /* (4, 15, 8) {real, imag} */,
  {32'h3c03eda0, 32'h3c8a4d10} /* (4, 15, 7) {real, imag} */,
  {32'h3e4202ed, 32'hbd6b4678} /* (4, 15, 6) {real, imag} */,
  {32'hbf10df56, 32'h3bad5d40} /* (4, 15, 5) {real, imag} */,
  {32'h3e55bcfd, 32'hbd3ce4e8} /* (4, 15, 4) {real, imag} */,
  {32'h3e8b052b, 32'hbe8388e3} /* (4, 15, 3) {real, imag} */,
  {32'hbe1e7fbf, 32'h3eb20965} /* (4, 15, 2) {real, imag} */,
  {32'hbe4e915e, 32'hbeaad585} /* (4, 15, 1) {real, imag} */,
  {32'hbe009e79, 32'hbf22b519} /* (4, 15, 0) {real, imag} */,
  {32'h3ebde1f4, 32'h3ed57bf3} /* (4, 14, 31) {real, imag} */,
  {32'hbe13a2fb, 32'hbc8aa980} /* (4, 14, 30) {real, imag} */,
  {32'h3e520597, 32'hbeefc10b} /* (4, 14, 29) {real, imag} */,
  {32'hbe6a904e, 32'h3d20bdac} /* (4, 14, 28) {real, imag} */,
  {32'h3e20ec51, 32'hbecb2452} /* (4, 14, 27) {real, imag} */,
  {32'hbe28bfca, 32'h3e981029} /* (4, 14, 26) {real, imag} */,
  {32'h3e0baa91, 32'h3b8d7200} /* (4, 14, 25) {real, imag} */,
  {32'h3e82b6af, 32'h3e37f8ff} /* (4, 14, 24) {real, imag} */,
  {32'h3d735d00, 32'hbeb6083b} /* (4, 14, 23) {real, imag} */,
  {32'h3d448ec6, 32'h3cc29cbc} /* (4, 14, 22) {real, imag} */,
  {32'h3e6a2bc0, 32'h3ee08db6} /* (4, 14, 21) {real, imag} */,
  {32'h3d733c53, 32'hbd0ab9f6} /* (4, 14, 20) {real, imag} */,
  {32'hbeb4b0c8, 32'h3d84bc37} /* (4, 14, 19) {real, imag} */,
  {32'h3d9ec598, 32'hbf0b9cac} /* (4, 14, 18) {real, imag} */,
  {32'h3dc4b6a1, 32'hbd908d10} /* (4, 14, 17) {real, imag} */,
  {32'hbd60d194, 32'hbdbe6cdf} /* (4, 14, 16) {real, imag} */,
  {32'hbeae5476, 32'hbd0adf76} /* (4, 14, 15) {real, imag} */,
  {32'hbd254628, 32'h3dd53c6d} /* (4, 14, 14) {real, imag} */,
  {32'hbe4e4b89, 32'h3d2dfac0} /* (4, 14, 13) {real, imag} */,
  {32'hbe157404, 32'hbe1ec32d} /* (4, 14, 12) {real, imag} */,
  {32'h3d3a54bc, 32'h3ed90d88} /* (4, 14, 11) {real, imag} */,
  {32'hbdfbd376, 32'hbde50202} /* (4, 14, 10) {real, imag} */,
  {32'h3f1e105c, 32'hbe8493b0} /* (4, 14, 9) {real, imag} */,
  {32'hbda6c327, 32'hbe6a7a70} /* (4, 14, 8) {real, imag} */,
  {32'hbe1d71e9, 32'hbec6baf8} /* (4, 14, 7) {real, imag} */,
  {32'h3d578dca, 32'h3d02e044} /* (4, 14, 6) {real, imag} */,
  {32'h3dc71f62, 32'hbe1e4bd3} /* (4, 14, 5) {real, imag} */,
  {32'h3e84afd4, 32'h3ea5e6fa} /* (4, 14, 4) {real, imag} */,
  {32'h3db8bb9c, 32'hbd68c250} /* (4, 14, 3) {real, imag} */,
  {32'hbdaaf6bd, 32'hbc0213c0} /* (4, 14, 2) {real, imag} */,
  {32'hbf0a05a3, 32'hbe60aee1} /* (4, 14, 1) {real, imag} */,
  {32'h3ca9b15e, 32'h3e5edb95} /* (4, 14, 0) {real, imag} */,
  {32'hbee0b363, 32'hbe37e0a3} /* (4, 13, 31) {real, imag} */,
  {32'h3dfcea61, 32'h3cb68af6} /* (4, 13, 30) {real, imag} */,
  {32'h3d8be66a, 32'hbef76306} /* (4, 13, 29) {real, imag} */,
  {32'h3c856927, 32'hbc9bd0c4} /* (4, 13, 28) {real, imag} */,
  {32'hbe2f39b6, 32'hbe8a70b6} /* (4, 13, 27) {real, imag} */,
  {32'hbe8c9da8, 32'hbe3eee28} /* (4, 13, 26) {real, imag} */,
  {32'h3e209502, 32'h3eef0977} /* (4, 13, 25) {real, imag} */,
  {32'h3eb89654, 32'hbd2bfe5a} /* (4, 13, 24) {real, imag} */,
  {32'hbed2ef3e, 32'h3f00729b} /* (4, 13, 23) {real, imag} */,
  {32'h3d0d87ea, 32'hbe91e0fb} /* (4, 13, 22) {real, imag} */,
  {32'h3f20011e, 32'h3e260d2a} /* (4, 13, 21) {real, imag} */,
  {32'hbed8cec0, 32'hbe94864b} /* (4, 13, 20) {real, imag} */,
  {32'hbeaf2e17, 32'hbd99b804} /* (4, 13, 19) {real, imag} */,
  {32'h3d23191c, 32'hbead724b} /* (4, 13, 18) {real, imag} */,
  {32'hbe4b41bc, 32'hbe87c172} /* (4, 13, 17) {real, imag} */,
  {32'h3dc0963c, 32'hbdc8b7de} /* (4, 13, 16) {real, imag} */,
  {32'h3e9e907c, 32'hbf1a865a} /* (4, 13, 15) {real, imag} */,
  {32'hbe443ee4, 32'h3d7aeee6} /* (4, 13, 14) {real, imag} */,
  {32'hbe7dda77, 32'h3f1649ec} /* (4, 13, 13) {real, imag} */,
  {32'h3e3d52d2, 32'h3e03ca20} /* (4, 13, 12) {real, imag} */,
  {32'h3e31df36, 32'hbe20080a} /* (4, 13, 11) {real, imag} */,
  {32'hbee302b2, 32'h3dd0da09} /* (4, 13, 10) {real, imag} */,
  {32'h3e94b8cc, 32'h3ac65fc0} /* (4, 13, 9) {real, imag} */,
  {32'hbe005535, 32'h3f28e5b8} /* (4, 13, 8) {real, imag} */,
  {32'hbf0f7b47, 32'hbed0524d} /* (4, 13, 7) {real, imag} */,
  {32'hbe9a9d6b, 32'hbeed9c43} /* (4, 13, 6) {real, imag} */,
  {32'hbeb83d48, 32'h3e35f46f} /* (4, 13, 5) {real, imag} */,
  {32'hbe87b390, 32'hbe2b80d3} /* (4, 13, 4) {real, imag} */,
  {32'hbd8b7f01, 32'hbe572df0} /* (4, 13, 3) {real, imag} */,
  {32'h3e45f5c0, 32'h3e9386b2} /* (4, 13, 2) {real, imag} */,
  {32'h3e91592d, 32'hbe9b3ebe} /* (4, 13, 1) {real, imag} */,
  {32'hbe433b5f, 32'h3e1027fc} /* (4, 13, 0) {real, imag} */,
  {32'hbe12be58, 32'h3de1b2b9} /* (4, 12, 31) {real, imag} */,
  {32'hbe8c0730, 32'h3eeb5854} /* (4, 12, 30) {real, imag} */,
  {32'hbebf797f, 32'h3e366946} /* (4, 12, 29) {real, imag} */,
  {32'h3e869960, 32'h3d8170a0} /* (4, 12, 28) {real, imag} */,
  {32'h3e94ae47, 32'hbe2ffd42} /* (4, 12, 27) {real, imag} */,
  {32'hbef66a56, 32'hbe0d9a7e} /* (4, 12, 26) {real, imag} */,
  {32'hbdc72cac, 32'hbf254263} /* (4, 12, 25) {real, imag} */,
  {32'h3e68b00e, 32'hbd3359f4} /* (4, 12, 24) {real, imag} */,
  {32'hbe9ddc40, 32'hbc8bfca0} /* (4, 12, 23) {real, imag} */,
  {32'h3ef58f7e, 32'hbf3e8e2a} /* (4, 12, 22) {real, imag} */,
  {32'h39016000, 32'h3f08e4d9} /* (4, 12, 21) {real, imag} */,
  {32'hbe9566e1, 32'hbd3e69f4} /* (4, 12, 20) {real, imag} */,
  {32'h3f1c222a, 32'hbdb256e8} /* (4, 12, 19) {real, imag} */,
  {32'h3e6cb76b, 32'h3e2bb938} /* (4, 12, 18) {real, imag} */,
  {32'h3ed59e90, 32'h3e18a8d2} /* (4, 12, 17) {real, imag} */,
  {32'hbb46f680, 32'hbcebf288} /* (4, 12, 16) {real, imag} */,
  {32'hbf0d3e21, 32'h3ddfc7d6} /* (4, 12, 15) {real, imag} */,
  {32'h3eb9f0cf, 32'h3dbb215c} /* (4, 12, 14) {real, imag} */,
  {32'hbe331ccc, 32'h3e92a0fc} /* (4, 12, 13) {real, imag} */,
  {32'h3ee8d0a4, 32'h3e95f91b} /* (4, 12, 12) {real, imag} */,
  {32'h3e0b461e, 32'hbdb3efdf} /* (4, 12, 11) {real, imag} */,
  {32'hbf160b06, 32'hbe2f4732} /* (4, 12, 10) {real, imag} */,
  {32'h3ea34800, 32'h3df32792} /* (4, 12, 9) {real, imag} */,
  {32'h3edb36f0, 32'h3ef6469d} /* (4, 12, 8) {real, imag} */,
  {32'h3e28c94b, 32'hbd031de0} /* (4, 12, 7) {real, imag} */,
  {32'h3e52346c, 32'h3e0a482a} /* (4, 12, 6) {real, imag} */,
  {32'h3e7cbcdc, 32'hbf36f8ff} /* (4, 12, 5) {real, imag} */,
  {32'hbe8eb760, 32'h3ed9936b} /* (4, 12, 4) {real, imag} */,
  {32'hbea6fb48, 32'hbe50cad7} /* (4, 12, 3) {real, imag} */,
  {32'h3da535a3, 32'h3e345999} /* (4, 12, 2) {real, imag} */,
  {32'h3dd9867b, 32'hbe577070} /* (4, 12, 1) {real, imag} */,
  {32'hbe80a0d0, 32'h3c03ff10} /* (4, 12, 0) {real, imag} */,
  {32'h3e7be16f, 32'h3f142e25} /* (4, 11, 31) {real, imag} */,
  {32'hbee50f46, 32'hbe904dd9} /* (4, 11, 30) {real, imag} */,
  {32'hbeef962b, 32'h3dfcf4a6} /* (4, 11, 29) {real, imag} */,
  {32'h3e53e39a, 32'h3d7e3264} /* (4, 11, 28) {real, imag} */,
  {32'hbe0294f9, 32'hbee8d502} /* (4, 11, 27) {real, imag} */,
  {32'hbe41eb7a, 32'h3dfc5a1c} /* (4, 11, 26) {real, imag} */,
  {32'h3e97809e, 32'h3d805c28} /* (4, 11, 25) {real, imag} */,
  {32'hbe20a292, 32'h3e3e1d1a} /* (4, 11, 24) {real, imag} */,
  {32'h3c8a7eac, 32'hbe9a53f4} /* (4, 11, 23) {real, imag} */,
  {32'hbe8a2ce6, 32'h3e9dcb7a} /* (4, 11, 22) {real, imag} */,
  {32'hbea8abac, 32'hbcf83dd8} /* (4, 11, 21) {real, imag} */,
  {32'h3e86405e, 32'hbde4a1c0} /* (4, 11, 20) {real, imag} */,
  {32'hbda16326, 32'h3d80c008} /* (4, 11, 19) {real, imag} */,
  {32'hbed95252, 32'h3e7de3e4} /* (4, 11, 18) {real, imag} */,
  {32'hbe286992, 32'hbee7172c} /* (4, 11, 17) {real, imag} */,
  {32'h3e6cb998, 32'h3d9648f4} /* (4, 11, 16) {real, imag} */,
  {32'hbc2ccc60, 32'h3e71afcc} /* (4, 11, 15) {real, imag} */,
  {32'h3f21c805, 32'hbe141a42} /* (4, 11, 14) {real, imag} */,
  {32'hbdf6f52d, 32'hbea551cf} /* (4, 11, 13) {real, imag} */,
  {32'hbeddd17f, 32'hbe98d912} /* (4, 11, 12) {real, imag} */,
  {32'hbe9466bd, 32'hbebf53b6} /* (4, 11, 11) {real, imag} */,
  {32'hbea8364b, 32'h3dfd36ed} /* (4, 11, 10) {real, imag} */,
  {32'hbeb61251, 32'h3e5591b2} /* (4, 11, 9) {real, imag} */,
  {32'hbe86a89a, 32'hbdd365a8} /* (4, 11, 8) {real, imag} */,
  {32'h3eefe189, 32'h3bcdcc80} /* (4, 11, 7) {real, imag} */,
  {32'h3f250f17, 32'h3e6324a2} /* (4, 11, 6) {real, imag} */,
  {32'hbec0be68, 32'h3dfc301c} /* (4, 11, 5) {real, imag} */,
  {32'hbd4eb084, 32'hbe98016b} /* (4, 11, 4) {real, imag} */,
  {32'hbf35d760, 32'hbe37a610} /* (4, 11, 3) {real, imag} */,
  {32'hbde18118, 32'hbedd7304} /* (4, 11, 2) {real, imag} */,
  {32'hbd80a81a, 32'h3f9cb290} /* (4, 11, 1) {real, imag} */,
  {32'h3f8660cc, 32'h3e762072} /* (4, 11, 0) {real, imag} */,
  {32'h3ef6bb58, 32'hbeb9fcc1} /* (4, 10, 31) {real, imag} */,
  {32'h3d21578a, 32'hbea9f866} /* (4, 10, 30) {real, imag} */,
  {32'hbf189a9f, 32'h3f223602} /* (4, 10, 29) {real, imag} */,
  {32'hbdc9591a, 32'h3d6b2b8c} /* (4, 10, 28) {real, imag} */,
  {32'h3f42bee3, 32'h3edf7075} /* (4, 10, 27) {real, imag} */,
  {32'h3e9f318c, 32'hbe4dbfd4} /* (4, 10, 26) {real, imag} */,
  {32'hbe26dc0e, 32'hbe258dfe} /* (4, 10, 25) {real, imag} */,
  {32'hbe94c565, 32'h3f36e4c9} /* (4, 10, 24) {real, imag} */,
  {32'h3dcda5a8, 32'hbd35c26f} /* (4, 10, 23) {real, imag} */,
  {32'hbe90e90c, 32'h3ec90885} /* (4, 10, 22) {real, imag} */,
  {32'hbe50fc34, 32'hbece4c9a} /* (4, 10, 21) {real, imag} */,
  {32'h3ee3d019, 32'h3e38ee5a} /* (4, 10, 20) {real, imag} */,
  {32'hbd42e5b0, 32'h3d81ef3a} /* (4, 10, 19) {real, imag} */,
  {32'hbd98bdc8, 32'h3e143618} /* (4, 10, 18) {real, imag} */,
  {32'h3d34f966, 32'h3e429718} /* (4, 10, 17) {real, imag} */,
  {32'h3d950843, 32'h3ecd3674} /* (4, 10, 16) {real, imag} */,
  {32'h3e0e69dd, 32'hbe0bf8c9} /* (4, 10, 15) {real, imag} */,
  {32'hbe2b5cd8, 32'h3e6eacd3} /* (4, 10, 14) {real, imag} */,
  {32'hbd7d0e64, 32'h3e4a823c} /* (4, 10, 13) {real, imag} */,
  {32'h3f18d087, 32'hbe541000} /* (4, 10, 12) {real, imag} */,
  {32'h3f24c715, 32'h3e75e8d0} /* (4, 10, 11) {real, imag} */,
  {32'h3e9c961c, 32'hbe91d848} /* (4, 10, 10) {real, imag} */,
  {32'hbc29cb40, 32'h3eefd94e} /* (4, 10, 9) {real, imag} */,
  {32'hbe8be33c, 32'h3e834964} /* (4, 10, 8) {real, imag} */,
  {32'hbeacfcfa, 32'h3e8abef6} /* (4, 10, 7) {real, imag} */,
  {32'h3f0101bf, 32'h3eba6e1c} /* (4, 10, 6) {real, imag} */,
  {32'h3e8ae95b, 32'hbf164c3e} /* (4, 10, 5) {real, imag} */,
  {32'hbd10d1b0, 32'hbe6468db} /* (4, 10, 4) {real, imag} */,
  {32'hbe599177, 32'hbe70a243} /* (4, 10, 3) {real, imag} */,
  {32'h3f1c9715, 32'h3e9a3eb5} /* (4, 10, 2) {real, imag} */,
  {32'hbed97c3b, 32'hbd288c3e} /* (4, 10, 1) {real, imag} */,
  {32'hbf03c667, 32'hbf292d22} /* (4, 10, 0) {real, imag} */,
  {32'h3e8b6442, 32'hbcf435d0} /* (4, 9, 31) {real, imag} */,
  {32'h3dc8b4a4, 32'hbd5a6310} /* (4, 9, 30) {real, imag} */,
  {32'hbdf576c4, 32'hbed560b5} /* (4, 9, 29) {real, imag} */,
  {32'h3e02b1e6, 32'hbe6508a4} /* (4, 9, 28) {real, imag} */,
  {32'h3f31bbc6, 32'h3f01be5f} /* (4, 9, 27) {real, imag} */,
  {32'h3f28c2ad, 32'h3d81ea50} /* (4, 9, 26) {real, imag} */,
  {32'hbe55a559, 32'h3edf8cf1} /* (4, 9, 25) {real, imag} */,
  {32'hbe00a85d, 32'h3e0702c8} /* (4, 9, 24) {real, imag} */,
  {32'hbee0d8c3, 32'hbf3468e2} /* (4, 9, 23) {real, imag} */,
  {32'hbe3c7260, 32'hbef998b5} /* (4, 9, 22) {real, imag} */,
  {32'hbe0a4ea4, 32'hbebc2587} /* (4, 9, 21) {real, imag} */,
  {32'h3e6ca350, 32'h3f12c51f} /* (4, 9, 20) {real, imag} */,
  {32'hbf1d4502, 32'h3d5d1250} /* (4, 9, 19) {real, imag} */,
  {32'hbe0b90d4, 32'h3e7c0f7f} /* (4, 9, 18) {real, imag} */,
  {32'h3e0d9339, 32'h3e6942b7} /* (4, 9, 17) {real, imag} */,
  {32'hbebb66d0, 32'hbf062175} /* (4, 9, 16) {real, imag} */,
  {32'hbd81b6be, 32'hbe0684ca} /* (4, 9, 15) {real, imag} */,
  {32'hbe1cbca8, 32'hbd6bb618} /* (4, 9, 14) {real, imag} */,
  {32'hbde8e66c, 32'h3be52670} /* (4, 9, 13) {real, imag} */,
  {32'hbdaf059b, 32'hbeef5fd4} /* (4, 9, 12) {real, imag} */,
  {32'hbee3b1f2, 32'hbe9cfedb} /* (4, 9, 11) {real, imag} */,
  {32'h3ee0bf4a, 32'hbef882b2} /* (4, 9, 10) {real, imag} */,
  {32'hbe745db9, 32'h3e12ba80} /* (4, 9, 9) {real, imag} */,
  {32'hbd969ac7, 32'hbb8840c0} /* (4, 9, 8) {real, imag} */,
  {32'h3dd05204, 32'h3e14f5f6} /* (4, 9, 7) {real, imag} */,
  {32'hbd7954a6, 32'h3e834225} /* (4, 9, 6) {real, imag} */,
  {32'hbdf974ac, 32'hbe9b95cb} /* (4, 9, 5) {real, imag} */,
  {32'h3d9deec0, 32'hbeebca74} /* (4, 9, 4) {real, imag} */,
  {32'h3eb8de7e, 32'h3f3dc7bc} /* (4, 9, 3) {real, imag} */,
  {32'h3d2c7528, 32'h3dbcf69b} /* (4, 9, 2) {real, imag} */,
  {32'hbeea0e35, 32'hbe4d133a} /* (4, 9, 1) {real, imag} */,
  {32'hbe2ce468, 32'h3ef4ddbd} /* (4, 9, 0) {real, imag} */,
  {32'h3fbe96a6, 32'h3e8b7fcf} /* (4, 8, 31) {real, imag} */,
  {32'hbf8c18a4, 32'hbec378a6} /* (4, 8, 30) {real, imag} */,
  {32'h3e1e0f20, 32'h3e5504e2} /* (4, 8, 29) {real, imag} */,
  {32'h3edcc0f6, 32'hbdb013d6} /* (4, 8, 28) {real, imag} */,
  {32'h3e5a4f68, 32'hbecaa07c} /* (4, 8, 27) {real, imag} */,
  {32'h3e56a198, 32'hbe9450e8} /* (4, 8, 26) {real, imag} */,
  {32'hbeb77614, 32'h3e2ac088} /* (4, 8, 25) {real, imag} */,
  {32'hbf1d6e1d, 32'hbe2ba6a3} /* (4, 8, 24) {real, imag} */,
  {32'hbf24db44, 32'hbe880e71} /* (4, 8, 23) {real, imag} */,
  {32'hbed1cd81, 32'h3ea06be6} /* (4, 8, 22) {real, imag} */,
  {32'h3cfa9ac8, 32'h3ed6ecc7} /* (4, 8, 21) {real, imag} */,
  {32'h3ebf15fd, 32'hbef5e13e} /* (4, 8, 20) {real, imag} */,
  {32'hbea4bbd2, 32'h3e97fa5e} /* (4, 8, 19) {real, imag} */,
  {32'h3dc06782, 32'h3d98b7ca} /* (4, 8, 18) {real, imag} */,
  {32'h3e99801e, 32'h3dcfb8c2} /* (4, 8, 17) {real, imag} */,
  {32'h3b99a478, 32'hbe8f44ca} /* (4, 8, 16) {real, imag} */,
  {32'hbd5e8f66, 32'hbc5d7da8} /* (4, 8, 15) {real, imag} */,
  {32'h3e885a50, 32'h3f09a7e1} /* (4, 8, 14) {real, imag} */,
  {32'h3e35ac29, 32'hbedccfc0} /* (4, 8, 13) {real, imag} */,
  {32'hbddcd5b1, 32'h3e0f38d0} /* (4, 8, 12) {real, imag} */,
  {32'hbe84945a, 32'hb9f0ea00} /* (4, 8, 11) {real, imag} */,
  {32'h3f0e1ac9, 32'hbd60d3f0} /* (4, 8, 10) {real, imag} */,
  {32'h3eccecfc, 32'h3f1ba022} /* (4, 8, 9) {real, imag} */,
  {32'hbe8a4634, 32'h3e6baaee} /* (4, 8, 8) {real, imag} */,
  {32'hbe340eec, 32'h3da7aa38} /* (4, 8, 7) {real, imag} */,
  {32'hbe48d5a6, 32'h3ec9d87e} /* (4, 8, 6) {real, imag} */,
  {32'hbc0eb100, 32'hbf0d97ea} /* (4, 8, 5) {real, imag} */,
  {32'hbe065ddb, 32'hbd06cc7c} /* (4, 8, 4) {real, imag} */,
  {32'hbd431862, 32'h3d446f18} /* (4, 8, 3) {real, imag} */,
  {32'hbf286cd2, 32'hbf10e353} /* (4, 8, 2) {real, imag} */,
  {32'hbd71f918, 32'h3ee5830c} /* (4, 8, 1) {real, imag} */,
  {32'h3f2f95a3, 32'h3f892d0c} /* (4, 8, 0) {real, imag} */,
  {32'hbf5c7086, 32'hbcb7d3cc} /* (4, 7, 31) {real, imag} */,
  {32'hbe18814a, 32'h3f5ac3cc} /* (4, 7, 30) {real, imag} */,
  {32'hbe950396, 32'hbeb57b46} /* (4, 7, 29) {real, imag} */,
  {32'hbf0f8df0, 32'hbf3938dc} /* (4, 7, 28) {real, imag} */,
  {32'h3f2061da, 32'h3e5c7b8c} /* (4, 7, 27) {real, imag} */,
  {32'h3eae43f3, 32'hbe6014c9} /* (4, 7, 26) {real, imag} */,
  {32'h3df8483a, 32'hbe3d772a} /* (4, 7, 25) {real, imag} */,
  {32'hbed37006, 32'hbf11a78a} /* (4, 7, 24) {real, imag} */,
  {32'hbd3d584e, 32'h3ed32650} /* (4, 7, 23) {real, imag} */,
  {32'hbd6918f8, 32'hbea5e41c} /* (4, 7, 22) {real, imag} */,
  {32'hbe22fec1, 32'h3f007f1a} /* (4, 7, 21) {real, imag} */,
  {32'h3e9cd558, 32'hbe234132} /* (4, 7, 20) {real, imag} */,
  {32'hbe506284, 32'h3ef64ad2} /* (4, 7, 19) {real, imag} */,
  {32'h3efa3896, 32'hbe55b06f} /* (4, 7, 18) {real, imag} */,
  {32'hbce03174, 32'h3ea19cce} /* (4, 7, 17) {real, imag} */,
  {32'h3ed9987f, 32'hbdea32b2} /* (4, 7, 16) {real, imag} */,
  {32'hbee01659, 32'hbf0135a8} /* (4, 7, 15) {real, imag} */,
  {32'hbef14e8a, 32'hbccad230} /* (4, 7, 14) {real, imag} */,
  {32'hbf1e20eb, 32'h3eb0b5a8} /* (4, 7, 13) {real, imag} */,
  {32'hbf2de3e2, 32'h3da93420} /* (4, 7, 12) {real, imag} */,
  {32'hbe2e9a42, 32'h3eb57e0f} /* (4, 7, 11) {real, imag} */,
  {32'h3e270dfa, 32'hbe4a626a} /* (4, 7, 10) {real, imag} */,
  {32'h3eab1276, 32'h3dbbbd5c} /* (4, 7, 9) {real, imag} */,
  {32'h3e2e003e, 32'hbcf75d50} /* (4, 7, 8) {real, imag} */,
  {32'hbf188057, 32'h3e9e5b11} /* (4, 7, 7) {real, imag} */,
  {32'h3e9e4c54, 32'h3dacc3eb} /* (4, 7, 6) {real, imag} */,
  {32'h3f89f01a, 32'h3f463306} /* (4, 7, 5) {real, imag} */,
  {32'hbeedb3c9, 32'hbec112b2} /* (4, 7, 4) {real, imag} */,
  {32'hbbf6f0c0, 32'h3e867624} /* (4, 7, 3) {real, imag} */,
  {32'h3f16639d, 32'h3ea53c32} /* (4, 7, 2) {real, imag} */,
  {32'h3ba29c00, 32'hbf5e5ed0} /* (4, 7, 1) {real, imag} */,
  {32'hbf46088a, 32'hbe9a5c4a} /* (4, 7, 0) {real, imag} */,
  {32'h3f0566bc, 32'h3f271802} /* (4, 6, 31) {real, imag} */,
  {32'h3edb9333, 32'h3c4951e0} /* (4, 6, 30) {real, imag} */,
  {32'h3f32089d, 32'h3cb828b0} /* (4, 6, 29) {real, imag} */,
  {32'h3d8c20e0, 32'hbd083090} /* (4, 6, 28) {real, imag} */,
  {32'h3d300010, 32'h3f1e2a76} /* (4, 6, 27) {real, imag} */,
  {32'hbd5e71a8, 32'hbe6cfeaa} /* (4, 6, 26) {real, imag} */,
  {32'hbcc943f4, 32'hbe925770} /* (4, 6, 25) {real, imag} */,
  {32'hbe892ce3, 32'h3ec74fc6} /* (4, 6, 24) {real, imag} */,
  {32'hbeeb0d7a, 32'hbe18251d} /* (4, 6, 23) {real, imag} */,
  {32'hbe068bab, 32'h3f036a8e} /* (4, 6, 22) {real, imag} */,
  {32'hbe76a4e3, 32'hbf20ff26} /* (4, 6, 21) {real, imag} */,
  {32'hbf29831d, 32'h3e513631} /* (4, 6, 20) {real, imag} */,
  {32'hbe469ca9, 32'hbe112fe4} /* (4, 6, 19) {real, imag} */,
  {32'h3df843ba, 32'h3cb136bc} /* (4, 6, 18) {real, imag} */,
  {32'h3e72f80c, 32'hbda8b098} /* (4, 6, 17) {real, imag} */,
  {32'h3d8cfa67, 32'hbe15ce90} /* (4, 6, 16) {real, imag} */,
  {32'hbc5222a8, 32'h3d87ce34} /* (4, 6, 15) {real, imag} */,
  {32'hbd4d22e8, 32'hbec5f147} /* (4, 6, 14) {real, imag} */,
  {32'h3f00fb91, 32'hbdfe01a6} /* (4, 6, 13) {real, imag} */,
  {32'h3e6cc65e, 32'h3de58426} /* (4, 6, 12) {real, imag} */,
  {32'hbecd18c7, 32'h3e54a510} /* (4, 6, 11) {real, imag} */,
  {32'h3cbc4608, 32'hbdc93292} /* (4, 6, 10) {real, imag} */,
  {32'h3e4f6151, 32'hbcb19528} /* (4, 6, 9) {real, imag} */,
  {32'hbf2af1fe, 32'hbcc8a370} /* (4, 6, 8) {real, imag} */,
  {32'h3ea255d4, 32'h3eb40a5b} /* (4, 6, 7) {real, imag} */,
  {32'hbf22dcb0, 32'hbe9ad7a4} /* (4, 6, 6) {real, imag} */,
  {32'hbe1d9fa9, 32'h3e41d63a} /* (4, 6, 5) {real, imag} */,
  {32'hbe39af60, 32'hbe9a5db0} /* (4, 6, 4) {real, imag} */,
  {32'hbeb4a0be, 32'h3e4159b7} /* (4, 6, 3) {real, imag} */,
  {32'hbf2e8ad9, 32'hbe091fca} /* (4, 6, 2) {real, imag} */,
  {32'h3f08b211, 32'h3ec4fc49} /* (4, 6, 1) {real, imag} */,
  {32'h3ed1757b, 32'hbf126d0f} /* (4, 6, 0) {real, imag} */,
  {32'h3fda6421, 32'h3f324c80} /* (4, 5, 31) {real, imag} */,
  {32'hbfafeab3, 32'hbecd9c0a} /* (4, 5, 30) {real, imag} */,
  {32'hbdbb7eaa, 32'hbebb7e25} /* (4, 5, 29) {real, imag} */,
  {32'h3f3a9428, 32'hbf2f9882} /* (4, 5, 28) {real, imag} */,
  {32'hbf2819a3, 32'hbe199575} /* (4, 5, 27) {real, imag} */,
  {32'hbe9a5dea, 32'h3ea95625} /* (4, 5, 26) {real, imag} */,
  {32'h3f445c7e, 32'h3ea7cbc8} /* (4, 5, 25) {real, imag} */,
  {32'hbe8a68f8, 32'hbd4bb67e} /* (4, 5, 24) {real, imag} */,
  {32'h3e35de95, 32'hbee10bf2} /* (4, 5, 23) {real, imag} */,
  {32'hbd876fa0, 32'h3c95ce48} /* (4, 5, 22) {real, imag} */,
  {32'hbe8a65c0, 32'h3f6962b4} /* (4, 5, 21) {real, imag} */,
  {32'hbe6de98c, 32'h3e0eaf0e} /* (4, 5, 20) {real, imag} */,
  {32'hbeba10a6, 32'h3d254dc0} /* (4, 5, 19) {real, imag} */,
  {32'h3eafd40e, 32'h3e60cafe} /* (4, 5, 18) {real, imag} */,
  {32'hbe61e64c, 32'h3e74062e} /* (4, 5, 17) {real, imag} */,
  {32'hbd87ff72, 32'h3e824680} /* (4, 5, 16) {real, imag} */,
  {32'h3e691b94, 32'hbe248f20} /* (4, 5, 15) {real, imag} */,
  {32'h3eaa229e, 32'hbe5f34f4} /* (4, 5, 14) {real, imag} */,
  {32'hbdd0a042, 32'hbeaa4d8f} /* (4, 5, 13) {real, imag} */,
  {32'hbe184681, 32'h3dcbee1c} /* (4, 5, 12) {real, imag} */,
  {32'hbdd5cc9e, 32'hbf522e0e} /* (4, 5, 11) {real, imag} */,
  {32'h3e5bab23, 32'h3f0dbbd8} /* (4, 5, 10) {real, imag} */,
  {32'hbc57a1f0, 32'h3d33ff90} /* (4, 5, 9) {real, imag} */,
  {32'h3dcc4244, 32'hbdc8e5ae} /* (4, 5, 8) {real, imag} */,
  {32'hbd14a736, 32'h3e1b60f2} /* (4, 5, 7) {real, imag} */,
  {32'hbeaa11f4, 32'hbedaaea5} /* (4, 5, 6) {real, imag} */,
  {32'hbf4d0fde, 32'hbf75e207} /* (4, 5, 5) {real, imag} */,
  {32'h3f0ac180, 32'hbe732361} /* (4, 5, 4) {real, imag} */,
  {32'h3f28b277, 32'h3de41184} /* (4, 5, 3) {real, imag} */,
  {32'h3e79080c, 32'h3f462afb} /* (4, 5, 2) {real, imag} */,
  {32'h40247c5e, 32'h3fa17a40} /* (4, 5, 1) {real, imag} */,
  {32'h4023bf55, 32'hbe32cd1c} /* (4, 5, 0) {real, imag} */,
  {32'hbfa23b39, 32'hc024f48e} /* (4, 4, 31) {real, imag} */,
  {32'h3fa91cb5, 32'h4039daec} /* (4, 4, 30) {real, imag} */,
  {32'hbe483d1a, 32'h3e72d4fc} /* (4, 4, 29) {real, imag} */,
  {32'hbf0fc2ba, 32'h3e73c6e3} /* (4, 4, 28) {real, imag} */,
  {32'h3d2a71c2, 32'hbeec7ef0} /* (4, 4, 27) {real, imag} */,
  {32'hbfa3cb80, 32'hbeb98b2c} /* (4, 4, 26) {real, imag} */,
  {32'h3e93b0b0, 32'h3b89ec20} /* (4, 4, 25) {real, imag} */,
  {32'h3e96f687, 32'hbc375778} /* (4, 4, 24) {real, imag} */,
  {32'h3d2460c8, 32'h3dfec0db} /* (4, 4, 23) {real, imag} */,
  {32'h3eadcdbb, 32'hbdd7924f} /* (4, 4, 22) {real, imag} */,
  {32'h3f72c0ca, 32'hbe7dac7d} /* (4, 4, 21) {real, imag} */,
  {32'hbe11bdc4, 32'h3e09679a} /* (4, 4, 20) {real, imag} */,
  {32'h3e57c127, 32'hbe2afcbc} /* (4, 4, 19) {real, imag} */,
  {32'h3b0bd940, 32'h3e54eab6} /* (4, 4, 18) {real, imag} */,
  {32'hbdbe688e, 32'h3ebb3a58} /* (4, 4, 17) {real, imag} */,
  {32'hbe4f493b, 32'hbe7d1e16} /* (4, 4, 16) {real, imag} */,
  {32'hbe7b58e8, 32'hbd274958} /* (4, 4, 15) {real, imag} */,
  {32'hbdc79f21, 32'h3ed15276} /* (4, 4, 14) {real, imag} */,
  {32'hbe0385e5, 32'hbd9add16} /* (4, 4, 13) {real, imag} */,
  {32'hbca8b274, 32'hbc6ca9c0} /* (4, 4, 12) {real, imag} */,
  {32'hbc5fd01c, 32'hbea8f18f} /* (4, 4, 11) {real, imag} */,
  {32'h3ec4f75c, 32'hbed9ae4a} /* (4, 4, 10) {real, imag} */,
  {32'hbc7ef2d0, 32'h3ed6adb8} /* (4, 4, 9) {real, imag} */,
  {32'h3db48c1a, 32'h3e8dd106} /* (4, 4, 8) {real, imag} */,
  {32'hbf256632, 32'h3e51664a} /* (4, 4, 7) {real, imag} */,
  {32'h3ddecf00, 32'hbeac1a5e} /* (4, 4, 6) {real, imag} */,
  {32'h3f274907, 32'hbe3dd40c} /* (4, 4, 5) {real, imag} */,
  {32'h3f3820bc, 32'hbf075424} /* (4, 4, 4) {real, imag} */,
  {32'hbf1e1673, 32'h3f659480} /* (4, 4, 3) {real, imag} */,
  {32'h40321df1, 32'h3fc393a6} /* (4, 4, 2) {real, imag} */,
  {32'hc098991c, 32'hbfc626ac} /* (4, 4, 1) {real, imag} */,
  {32'hbfb7cfd6, 32'hbea04cc8} /* (4, 4, 0) {real, imag} */,
  {32'h40289fe7, 32'hbfd97180} /* (4, 3, 31) {real, imag} */,
  {32'hbfbae113, 32'h3f8d1e00} /* (4, 3, 30) {real, imag} */,
  {32'hbc756a00, 32'h3e8f23ed} /* (4, 3, 29) {real, imag} */,
  {32'hbf4b52c6, 32'hbeb8f8bd} /* (4, 3, 28) {real, imag} */,
  {32'h3f817646, 32'hbf449091} /* (4, 3, 27) {real, imag} */,
  {32'hbe7d5344, 32'hbeebf55c} /* (4, 3, 26) {real, imag} */,
  {32'hbe79a733, 32'h3ed1590e} /* (4, 3, 25) {real, imag} */,
  {32'h3df8f89e, 32'h3f32c1a8} /* (4, 3, 24) {real, imag} */,
  {32'hbe20fa2c, 32'hbf179d86} /* (4, 3, 23) {real, imag} */,
  {32'h3eb01c06, 32'hbefbac9d} /* (4, 3, 22) {real, imag} */,
  {32'hbea73458, 32'hbe7a333c} /* (4, 3, 21) {real, imag} */,
  {32'h3d4ae430, 32'hbbc9e8f4} /* (4, 3, 20) {real, imag} */,
  {32'hbe79d999, 32'hbe517123} /* (4, 3, 19) {real, imag} */,
  {32'hbf16f64a, 32'hbde31ac6} /* (4, 3, 18) {real, imag} */,
  {32'h3e9d0c24, 32'h3db7d1b9} /* (4, 3, 17) {real, imag} */,
  {32'h3e9a36fe, 32'hbea8093b} /* (4, 3, 16) {real, imag} */,
  {32'h3e16a47c, 32'h3c0ec6a8} /* (4, 3, 15) {real, imag} */,
  {32'hbd358f34, 32'h3ed2fef7} /* (4, 3, 14) {real, imag} */,
  {32'h3e9d5c2e, 32'h3dccbda8} /* (4, 3, 13) {real, imag} */,
  {32'h3e9e4222, 32'hbe9d30db} /* (4, 3, 12) {real, imag} */,
  {32'hbef04451, 32'hbe04d772} /* (4, 3, 11) {real, imag} */,
  {32'h3d145574, 32'hbe0afe0c} /* (4, 3, 10) {real, imag} */,
  {32'hbe2a23b5, 32'hbdd2ad2c} /* (4, 3, 9) {real, imag} */,
  {32'h3cd52ca8, 32'h3ee70325} /* (4, 3, 8) {real, imag} */,
  {32'hbe11466c, 32'hbf78531c} /* (4, 3, 7) {real, imag} */,
  {32'h3be85580, 32'hbea6a326} /* (4, 3, 6) {real, imag} */,
  {32'hbf5aba0f, 32'hbe9c7bec} /* (4, 3, 5) {real, imag} */,
  {32'h3f550140, 32'hbf3e00e3} /* (4, 3, 4) {real, imag} */,
  {32'hbe8f8a99, 32'hbf0e8801} /* (4, 3, 3) {real, imag} */,
  {32'h3edb17d7, 32'h40613b1e} /* (4, 3, 2) {real, imag} */,
  {32'hc0178967, 32'h3ea990d8} /* (4, 3, 1) {real, imag} */,
  {32'h3ed3a6a1, 32'h3f4cb1aa} /* (4, 3, 0) {real, imag} */,
  {32'h416ccb8f, 32'h3f609371} /* (4, 2, 31) {real, imag} */,
  {32'hc0ed9e45, 32'h3fcbfea8} /* (4, 2, 30) {real, imag} */,
  {32'h3cf6fe20, 32'h3f74cdb0} /* (4, 2, 29) {real, imag} */,
  {32'h3e9b3a96, 32'hc00ba956} /* (4, 2, 28) {real, imag} */,
  {32'hbfc77ed0, 32'h3f27ce8e} /* (4, 2, 27) {real, imag} */,
  {32'hbf5336de, 32'h3f7f7bee} /* (4, 2, 26) {real, imag} */,
  {32'h3e8819cc, 32'hbf8ac40f} /* (4, 2, 25) {real, imag} */,
  {32'hbea1c3ec, 32'h3ffee26a} /* (4, 2, 24) {real, imag} */,
  {32'hbea2c4dc, 32'h3e227409} /* (4, 2, 23) {real, imag} */,
  {32'h3c80fd80, 32'h3ea4ad02} /* (4, 2, 22) {real, imag} */,
  {32'hbea76fd4, 32'h3f2028fa} /* (4, 2, 21) {real, imag} */,
  {32'h3ea518f8, 32'hbde16509} /* (4, 2, 20) {real, imag} */,
  {32'hbde67f96, 32'hbe8bb15a} /* (4, 2, 19) {real, imag} */,
  {32'h3e1776e0, 32'h3de90e34} /* (4, 2, 18) {real, imag} */,
  {32'hbd236e56, 32'hbf0d98d2} /* (4, 2, 17) {real, imag} */,
  {32'h3e66aef0, 32'hbe52a889} /* (4, 2, 16) {real, imag} */,
  {32'h3e1adc31, 32'h3ebaa487} /* (4, 2, 15) {real, imag} */,
  {32'hbe18bb90, 32'hbf1c22a7} /* (4, 2, 14) {real, imag} */,
  {32'hbe3d1688, 32'hbe0bf04b} /* (4, 2, 13) {real, imag} */,
  {32'h3eb47e97, 32'h3e9c15f8} /* (4, 2, 12) {real, imag} */,
  {32'hbe9bf068, 32'hbeac79e1} /* (4, 2, 11) {real, imag} */,
  {32'h3e8ce546, 32'h3f2d22cf} /* (4, 2, 10) {real, imag} */,
  {32'h3e3c9e98, 32'h3e1f63ce} /* (4, 2, 9) {real, imag} */,
  {32'hbf7238c7, 32'hbec6e651} /* (4, 2, 8) {real, imag} */,
  {32'h3f31302c, 32'hbe613a6d} /* (4, 2, 7) {real, imag} */,
  {32'h3eb8a4d6, 32'h3f0b1eda} /* (4, 2, 6) {real, imag} */,
  {32'hbf271aba, 32'hbff13038} /* (4, 2, 5) {real, imag} */,
  {32'h4035abc9, 32'h3e2026fe} /* (4, 2, 4) {real, imag} */,
  {32'hbefa7a2c, 32'h3e94b956} /* (4, 2, 3) {real, imag} */,
  {32'hc0e31e4d, 32'h40792c8a} /* (4, 2, 2) {real, imag} */,
  {32'h4109ad3f, 32'h3d665600} /* (4, 2, 1) {real, imag} */,
  {32'h40af23e6, 32'h3e8f84c4} /* (4, 2, 0) {real, imag} */,
  {32'hc1131668, 32'h3f1a93d0} /* (4, 1, 31) {real, imag} */,
  {32'h40a68dc8, 32'h3f7c72eb} /* (4, 1, 30) {real, imag} */,
  {32'h3fc82ec2, 32'hbfa0f71e} /* (4, 1, 29) {real, imag} */,
  {32'hbfdeee70, 32'hc00f469a} /* (4, 1, 28) {real, imag} */,
  {32'h404b796e, 32'h3e290a2e} /* (4, 1, 27) {real, imag} */,
  {32'h3ef6b5ca, 32'hbf0101b6} /* (4, 1, 26) {real, imag} */,
  {32'hbf41b6c6, 32'hbdfe6a5a} /* (4, 1, 25) {real, imag} */,
  {32'h3f3acac0, 32'hbecb082a} /* (4, 1, 24) {real, imag} */,
  {32'hbe08855e, 32'h3d9f0d88} /* (4, 1, 23) {real, imag} */,
  {32'hbe2d9324, 32'hbf0bf683} /* (4, 1, 22) {real, imag} */,
  {32'h3f3f87c2, 32'hbe8fe028} /* (4, 1, 21) {real, imag} */,
  {32'h3de14bda, 32'h3dd941ec} /* (4, 1, 20) {real, imag} */,
  {32'h3e340592, 32'hbe4212ce} /* (4, 1, 19) {real, imag} */,
  {32'h3e16341b, 32'hbf0e4304} /* (4, 1, 18) {real, imag} */,
  {32'h3e9b17d8, 32'h3ea7b11e} /* (4, 1, 17) {real, imag} */,
  {32'hbed63d96, 32'hbe87be28} /* (4, 1, 16) {real, imag} */,
  {32'h3eb9a562, 32'h3d9c5e2a} /* (4, 1, 15) {real, imag} */,
  {32'hbf463230, 32'h3f11c066} /* (4, 1, 14) {real, imag} */,
  {32'h3e373c2e, 32'hbddaeacf} /* (4, 1, 13) {real, imag} */,
  {32'hbdee09ec, 32'hbe2d394b} /* (4, 1, 12) {real, imag} */,
  {32'hbe3badc9, 32'h3f0922e1} /* (4, 1, 11) {real, imag} */,
  {32'h3e80b80e, 32'h3df1e4ad} /* (4, 1, 10) {real, imag} */,
  {32'hbf2ba055, 32'h3f05b886} /* (4, 1, 9) {real, imag} */,
  {32'h3d074130, 32'h3f964f38} /* (4, 1, 8) {real, imag} */,
  {32'hbeeb9284, 32'hbdb51bf0} /* (4, 1, 7) {real, imag} */,
  {32'hbf311f6b, 32'hbf4bc0dd} /* (4, 1, 6) {real, imag} */,
  {32'h3ff8e9ef, 32'h3f53ca10} /* (4, 1, 5) {real, imag} */,
  {32'h3e1f04c4, 32'hbfa3ec2c} /* (4, 1, 4) {real, imag} */,
  {32'h3ecbffd6, 32'hbfcb2118} /* (4, 1, 3) {real, imag} */,
  {32'h40e356ee, 32'h40bbd49a} /* (4, 1, 2) {real, imag} */,
  {32'hc13b4b8d, 32'hc12d18d3} /* (4, 1, 1) {real, imag} */,
  {32'hbf22e928, 32'h3fdfb30c} /* (4, 1, 0) {real, imag} */,
  {32'hc0802b48, 32'h400b010e} /* (4, 0, 31) {real, imag} */,
  {32'h403178a0, 32'hbf8606a2} /* (4, 0, 30) {real, imag} */,
  {32'h402be6c6, 32'hbfc1d192} /* (4, 0, 29) {real, imag} */,
  {32'hbedb2781, 32'hc012e12e} /* (4, 0, 28) {real, imag} */,
  {32'h3fb5b418, 32'hbdc69068} /* (4, 0, 27) {real, imag} */,
  {32'h3f927170, 32'h3e991dd9} /* (4, 0, 26) {real, imag} */,
  {32'hbdc77c15, 32'h3e957b5c} /* (4, 0, 25) {real, imag} */,
  {32'hbf32e364, 32'hbf2d7932} /* (4, 0, 24) {real, imag} */,
  {32'h3db1fdf6, 32'hbe90a344} /* (4, 0, 23) {real, imag} */,
  {32'hbec1cffa, 32'hbeac7ff3} /* (4, 0, 22) {real, imag} */,
  {32'hbea3e3a0, 32'hbb4f8200} /* (4, 0, 21) {real, imag} */,
  {32'hbec9125f, 32'h3e2d5d7f} /* (4, 0, 20) {real, imag} */,
  {32'h3ee31407, 32'hbd2b79c4} /* (4, 0, 19) {real, imag} */,
  {32'h3e8c9958, 32'hbe3a2333} /* (4, 0, 18) {real, imag} */,
  {32'h3c8a8574, 32'h3e60d6f9} /* (4, 0, 17) {real, imag} */,
  {32'hbe304bee, 32'h00000000} /* (4, 0, 16) {real, imag} */,
  {32'h3c8a8574, 32'hbe60d6f9} /* (4, 0, 15) {real, imag} */,
  {32'h3e8c9958, 32'h3e3a2333} /* (4, 0, 14) {real, imag} */,
  {32'h3ee31407, 32'h3d2b79c4} /* (4, 0, 13) {real, imag} */,
  {32'hbec9125f, 32'hbe2d5d7f} /* (4, 0, 12) {real, imag} */,
  {32'hbea3e3a0, 32'h3b4f8200} /* (4, 0, 11) {real, imag} */,
  {32'hbec1cffa, 32'h3eac7ff3} /* (4, 0, 10) {real, imag} */,
  {32'h3db1fdf6, 32'h3e90a344} /* (4, 0, 9) {real, imag} */,
  {32'hbf32e364, 32'h3f2d7932} /* (4, 0, 8) {real, imag} */,
  {32'hbdc77c15, 32'hbe957b5c} /* (4, 0, 7) {real, imag} */,
  {32'h3f927170, 32'hbe991dd9} /* (4, 0, 6) {real, imag} */,
  {32'h3fb5b418, 32'h3dc69068} /* (4, 0, 5) {real, imag} */,
  {32'hbedb2781, 32'h4012e12e} /* (4, 0, 4) {real, imag} */,
  {32'h402be6c6, 32'h3fc1d192} /* (4, 0, 3) {real, imag} */,
  {32'h403178a0, 32'h3f8606a2} /* (4, 0, 2) {real, imag} */,
  {32'hc0802b48, 32'hc00b010e} /* (4, 0, 1) {real, imag} */,
  {32'h417d0662, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hc1c44884, 32'h418832a4} /* (3, 31, 31) {real, imag} */,
  {32'h411a0f1a, 32'hc10021d2} /* (3, 31, 30) {real, imag} */,
  {32'h3f9b1624, 32'h3f3d9cc4} /* (3, 31, 29) {real, imag} */,
  {32'hbf83f346, 32'h3f747e24} /* (3, 31, 28) {real, imag} */,
  {32'h3fff9bfe, 32'hbff6da63} /* (3, 31, 27) {real, imag} */,
  {32'hbdefcfec, 32'h3e5ba976} /* (3, 31, 26) {real, imag} */,
  {32'hbe5d5c60, 32'h3f0e732e} /* (3, 31, 25) {real, imag} */,
  {32'h3edd3728, 32'hbfaee7e5} /* (3, 31, 24) {real, imag} */,
  {32'hbec2dda8, 32'hbdf4d03e} /* (3, 31, 23) {real, imag} */,
  {32'h3e88b990, 32'hbecf17c0} /* (3, 31, 22) {real, imag} */,
  {32'h3ef17016, 32'hbf27e156} /* (3, 31, 21) {real, imag} */,
  {32'hbe8f4d6d, 32'hbdaa845d} /* (3, 31, 20) {real, imag} */,
  {32'hbd6c08e1, 32'h3e954215} /* (3, 31, 19) {real, imag} */,
  {32'hbe1c4f4c, 32'hbe1673d0} /* (3, 31, 18) {real, imag} */,
  {32'h3ea0b3ae, 32'hbe32bac3} /* (3, 31, 17) {real, imag} */,
  {32'h3e9d0f66, 32'hbc5563e0} /* (3, 31, 16) {real, imag} */,
  {32'h3e764116, 32'hbd6efffc} /* (3, 31, 15) {real, imag} */,
  {32'hbe76c315, 32'h3ee605fe} /* (3, 31, 14) {real, imag} */,
  {32'h3d7c7ecc, 32'h3d7e7eaa} /* (3, 31, 13) {real, imag} */,
  {32'hbd984bf1, 32'hbe0f84c3} /* (3, 31, 12) {real, imag} */,
  {32'h3f73d926, 32'h3f20416a} /* (3, 31, 11) {real, imag} */,
  {32'hbe75bda2, 32'hbdf06ba6} /* (3, 31, 10) {real, imag} */,
  {32'hbe788bdc, 32'h3d6695f0} /* (3, 31, 9) {real, imag} */,
  {32'h3f2b861f, 32'h3f44082b} /* (3, 31, 8) {real, imag} */,
  {32'hbf23b710, 32'hbe869f60} /* (3, 31, 7) {real, imag} */,
  {32'h3f95c0bb, 32'h3ec80d04} /* (3, 31, 6) {real, imag} */,
  {32'h407bad4c, 32'h3e45e14c} /* (3, 31, 5) {real, imag} */,
  {32'hc0354e47, 32'h3fccad5a} /* (3, 31, 4) {real, imag} */,
  {32'h3fdce602, 32'h3fa27adc} /* (3, 31, 3) {real, imag} */,
  {32'h40fb0f50, 32'hbfaefbf8} /* (3, 31, 2) {real, imag} */,
  {32'hc1910235, 32'hc03fa448} /* (3, 31, 1) {real, imag} */,
  {32'hc12818e4, 32'hbf85d494} /* (3, 31, 0) {real, imag} */,
  {32'h4143a854, 32'h3ed85dc0} /* (3, 30, 31) {real, imag} */,
  {32'hc10d518a, 32'hc08a34a9} /* (3, 30, 30) {real, imag} */,
  {32'hbf969306, 32'hbe0134c8} /* (3, 30, 29) {real, imag} */,
  {32'h4048385c, 32'h3e5b6714} /* (3, 30, 28) {real, imag} */,
  {32'hbfbca142, 32'h3f96aa0b} /* (3, 30, 27) {real, imag} */,
  {32'h3eac336c, 32'hbcb89968} /* (3, 30, 26) {real, imag} */,
  {32'h3f8a966e, 32'h3eaa65c0} /* (3, 30, 25) {real, imag} */,
  {32'hbf6a1dc3, 32'hbc9eed90} /* (3, 30, 24) {real, imag} */,
  {32'h3e5b206a, 32'h3ec81ca8} /* (3, 30, 23) {real, imag} */,
  {32'h3ef132e3, 32'hbb47f600} /* (3, 30, 22) {real, imag} */,
  {32'hbecd68e3, 32'hbed40cdc} /* (3, 30, 21) {real, imag} */,
  {32'h3f2e555e, 32'h3d5d6fe0} /* (3, 30, 20) {real, imag} */,
  {32'hbdeb1114, 32'h3dc5d86c} /* (3, 30, 19) {real, imag} */,
  {32'h3d99eede, 32'h3ed01514} /* (3, 30, 18) {real, imag} */,
  {32'h3f1017f2, 32'h3ebd9e46} /* (3, 30, 17) {real, imag} */,
  {32'h3d9a680a, 32'h3d151ce0} /* (3, 30, 16) {real, imag} */,
  {32'h3d98a610, 32'hbe8d610e} /* (3, 30, 15) {real, imag} */,
  {32'hbde30920, 32'hbf070199} /* (3, 30, 14) {real, imag} */,
  {32'hbd7a1530, 32'hbea4b86a} /* (3, 30, 13) {real, imag} */,
  {32'h3d8c8370, 32'h3ea1a997} /* (3, 30, 12) {real, imag} */,
  {32'hbeb0dc3a, 32'hbf6aa619} /* (3, 30, 11) {real, imag} */,
  {32'h3f0021a0, 32'h3f1acde5} /* (3, 30, 10) {real, imag} */,
  {32'hbf61a859, 32'h3e9e5474} /* (3, 30, 9) {real, imag} */,
  {32'hbf8256fc, 32'hbf1dd252} /* (3, 30, 8) {real, imag} */,
  {32'h3f4076aa, 32'h3f278db5} /* (3, 30, 7) {real, imag} */,
  {32'hbf09978d, 32'hbd15b70c} /* (3, 30, 6) {real, imag} */,
  {32'hbfc6582c, 32'hbfb746a4} /* (3, 30, 5) {real, imag} */,
  {32'h3f7495c3, 32'h4005928a} /* (3, 30, 4) {real, imag} */,
  {32'h3f41b4d3, 32'hbfb49180} /* (3, 30, 3) {real, imag} */,
  {32'hc127120c, 32'hc03dd0ef} /* (3, 30, 2) {real, imag} */,
  {32'h41a76ee7, 32'hbfc6afd1} /* (3, 30, 1) {real, imag} */,
  {32'h410ead27, 32'hc0203054} /* (3, 30, 0) {real, imag} */,
  {32'hc0574aea, 32'h3f4def58} /* (3, 29, 31) {real, imag} */,
  {32'hbed396bb, 32'hc08631b4} /* (3, 29, 30) {real, imag} */,
  {32'hbfa39ca2, 32'h3fb61e24} /* (3, 29, 29) {real, imag} */,
  {32'h3fa999f5, 32'hbe0b924e} /* (3, 29, 28) {real, imag} */,
  {32'hbf9c85a2, 32'hbf3b0683} /* (3, 29, 27) {real, imag} */,
  {32'h3d03ae38, 32'h3f7179c1} /* (3, 29, 26) {real, imag} */,
  {32'h3e7b7fe4, 32'h3f7dbab3} /* (3, 29, 25) {real, imag} */,
  {32'hbe0270ca, 32'hbef89a55} /* (3, 29, 24) {real, imag} */,
  {32'h3f528e27, 32'hbe275646} /* (3, 29, 23) {real, imag} */,
  {32'hbc5f8084, 32'h3e8457ae} /* (3, 29, 22) {real, imag} */,
  {32'hbf3133de, 32'h3f153ff2} /* (3, 29, 21) {real, imag} */,
  {32'hbe0284ce, 32'hbe7cf968} /* (3, 29, 20) {real, imag} */,
  {32'hbf26515f, 32'h3c8dd438} /* (3, 29, 19) {real, imag} */,
  {32'h3dc7d21b, 32'hbf352ec5} /* (3, 29, 18) {real, imag} */,
  {32'hbe7a3db0, 32'h3ccef150} /* (3, 29, 17) {real, imag} */,
  {32'hbe5f8e05, 32'h3e1e2474} /* (3, 29, 16) {real, imag} */,
  {32'hbe6490de, 32'hbd71d8f6} /* (3, 29, 15) {real, imag} */,
  {32'hbe015074, 32'h3d352572} /* (3, 29, 14) {real, imag} */,
  {32'h3e99d8fd, 32'hbcd00d48} /* (3, 29, 13) {real, imag} */,
  {32'hbcbe50f8, 32'hbe7f4ea1} /* (3, 29, 12) {real, imag} */,
  {32'h3dbf9ba4, 32'h3f13fba6} /* (3, 29, 11) {real, imag} */,
  {32'h3e5a1afa, 32'hbe9d646e} /* (3, 29, 10) {real, imag} */,
  {32'hbeec682b, 32'h3f12afbf} /* (3, 29, 9) {real, imag} */,
  {32'hbd8a957c, 32'hbf84ae04} /* (3, 29, 8) {real, imag} */,
  {32'hbe1dcb9f, 32'hbdc04326} /* (3, 29, 7) {real, imag} */,
  {32'hbdbe99dc, 32'hbe598268} /* (3, 29, 6) {real, imag} */,
  {32'h3f940c60, 32'h3d8b7768} /* (3, 29, 5) {real, imag} */,
  {32'hbec6ea7d, 32'h3e9f9c17} /* (3, 29, 4) {real, imag} */,
  {32'hbe5d3dea, 32'h3f541960} /* (3, 29, 3) {real, imag} */,
  {32'hbff9392a, 32'hbfbe9b4f} /* (3, 29, 2) {real, imag} */,
  {32'h408d693c, 32'h3fc3905a} /* (3, 29, 1) {real, imag} */,
  {32'h3f2f1a47, 32'h3f246520} /* (3, 29, 0) {real, imag} */,
  {32'hc0a90769, 32'h3ff63bdb} /* (3, 28, 31) {real, imag} */,
  {32'h403d88de, 32'hc01a7d25} /* (3, 28, 30) {real, imag} */,
  {32'h3e6e9915, 32'hbf964ecb} /* (3, 28, 29) {real, imag} */,
  {32'hbf6b9e66, 32'h3ecda3b2} /* (3, 28, 28) {real, imag} */,
  {32'h3ddc91a7, 32'hbf2f52e0} /* (3, 28, 27) {real, imag} */,
  {32'h3ec2633a, 32'hbeb13475} /* (3, 28, 26) {real, imag} */,
  {32'hbd24c26c, 32'hbed12b39} /* (3, 28, 25) {real, imag} */,
  {32'h3e599c9a, 32'hbed528f3} /* (3, 28, 24) {real, imag} */,
  {32'h3ef50e6d, 32'h3a458e00} /* (3, 28, 23) {real, imag} */,
  {32'hbcd33949, 32'h3e8df6e2} /* (3, 28, 22) {real, imag} */,
  {32'hbde75d09, 32'hbe05063c} /* (3, 28, 21) {real, imag} */,
  {32'hbd456ce4, 32'h3d989268} /* (3, 28, 20) {real, imag} */,
  {32'h3dfd4172, 32'hbef852bc} /* (3, 28, 19) {real, imag} */,
  {32'h3e0a91ea, 32'hbe4b3f46} /* (3, 28, 18) {real, imag} */,
  {32'h3c474160, 32'hbdb09dfa} /* (3, 28, 17) {real, imag} */,
  {32'h3e1c84eb, 32'h3cdfb802} /* (3, 28, 16) {real, imag} */,
  {32'hbde6faed, 32'h3debf3dc} /* (3, 28, 15) {real, imag} */,
  {32'h3f096b6d, 32'h3e8d1e38} /* (3, 28, 14) {real, imag} */,
  {32'hbddb2d97, 32'h3ec28c36} /* (3, 28, 13) {real, imag} */,
  {32'hbeb82a31, 32'hbef951d0} /* (3, 28, 12) {real, imag} */,
  {32'h3f6f032a, 32'h3d9e9408} /* (3, 28, 11) {real, imag} */,
  {32'hbf379946, 32'h3dd549cf} /* (3, 28, 10) {real, imag} */,
  {32'hbf222e48, 32'hbe2b3b33} /* (3, 28, 9) {real, imag} */,
  {32'hbeaf5aba, 32'h3eee86c6} /* (3, 28, 8) {real, imag} */,
  {32'h3da4a93c, 32'h3ee6029e} /* (3, 28, 7) {real, imag} */,
  {32'hbea4f123, 32'h3ea41377} /* (3, 28, 6) {real, imag} */,
  {32'h3f5cb5ec, 32'h3ddb6954} /* (3, 28, 5) {real, imag} */,
  {32'hbe48bb24, 32'h3f0ce2e6} /* (3, 28, 4) {real, imag} */,
  {32'hbeff6766, 32'hbf8d0e7c} /* (3, 28, 3) {real, imag} */,
  {32'h3f4fcfdd, 32'hc03c406b} /* (3, 28, 2) {real, imag} */,
  {32'hbfbf4fee, 32'h40359c6e} /* (3, 28, 1) {real, imag} */,
  {32'hc014b735, 32'h3f1912a0} /* (3, 28, 0) {real, imag} */,
  {32'h402d387a, 32'hc0213378} /* (3, 27, 31) {real, imag} */,
  {32'hbebbd2b8, 32'h3ece01e2} /* (3, 27, 30) {real, imag} */,
  {32'hbf0d44cc, 32'hbec15a4a} /* (3, 27, 29) {real, imag} */,
  {32'h3f098b80, 32'hbdeafea3} /* (3, 27, 28) {real, imag} */,
  {32'hbee268c2, 32'h3f5169f8} /* (3, 27, 27) {real, imag} */,
  {32'hbf46d7da, 32'h3c914be0} /* (3, 27, 26) {real, imag} */,
  {32'hbdefafa2, 32'h3c936170} /* (3, 27, 25) {real, imag} */,
  {32'hbe26f0f7, 32'hbe840b32} /* (3, 27, 24) {real, imag} */,
  {32'h3f292b9c, 32'hbe5e24e6} /* (3, 27, 23) {real, imag} */,
  {32'h3e801ca2, 32'h3e3adf63} /* (3, 27, 22) {real, imag} */,
  {32'hbe3d1e5c, 32'h3ec81b5c} /* (3, 27, 21) {real, imag} */,
  {32'hbdf7577a, 32'hbdc62f58} /* (3, 27, 20) {real, imag} */,
  {32'h3e06db1a, 32'h3ef70352} /* (3, 27, 19) {real, imag} */,
  {32'h3d10a7da, 32'h3dbcb9af} /* (3, 27, 18) {real, imag} */,
  {32'hbd75f7d0, 32'h3f208712} /* (3, 27, 17) {real, imag} */,
  {32'hbeb116d6, 32'hbdb16ca3} /* (3, 27, 16) {real, imag} */,
  {32'hbc858400, 32'h3db7161f} /* (3, 27, 15) {real, imag} */,
  {32'hbedc369e, 32'h3e4a5b06} /* (3, 27, 14) {real, imag} */,
  {32'hbbc7bff0, 32'hbc262428} /* (3, 27, 13) {real, imag} */,
  {32'h3d93a400, 32'hbe88234e} /* (3, 27, 12) {real, imag} */,
  {32'hbf3fe3c3, 32'hbe66d764} /* (3, 27, 11) {real, imag} */,
  {32'hbeeb317b, 32'hbe8f51a2} /* (3, 27, 10) {real, imag} */,
  {32'hbd3c3498, 32'h3d8fd190} /* (3, 27, 9) {real, imag} */,
  {32'hbed1bd33, 32'hbdb87ddf} /* (3, 27, 8) {real, imag} */,
  {32'h3eb2d7c6, 32'hbeaab2f3} /* (3, 27, 7) {real, imag} */,
  {32'h3ddb8fba, 32'h3e3f3041} /* (3, 27, 6) {real, imag} */,
  {32'hbf52a943, 32'h3b906940} /* (3, 27, 5) {real, imag} */,
  {32'h3ec839a4, 32'h3f53533c} /* (3, 27, 4) {real, imag} */,
  {32'hbf101288, 32'h3e9af5fe} /* (3, 27, 3) {real, imag} */,
  {32'hbf98ac70, 32'hbdf8793c} /* (3, 27, 2) {real, imag} */,
  {32'h40158132, 32'h3e9695ba} /* (3, 27, 1) {real, imag} */,
  {32'h402529fb, 32'hbe347bcc} /* (3, 27, 0) {real, imag} */,
  {32'h3f399064, 32'h3ee206e8} /* (3, 26, 31) {real, imag} */,
  {32'hbf39221e, 32'hbecae763} /* (3, 26, 30) {real, imag} */,
  {32'hbdf85086, 32'hbe8f9a78} /* (3, 26, 29) {real, imag} */,
  {32'h3e46cade, 32'h3e2d7ddf} /* (3, 26, 28) {real, imag} */,
  {32'hbe8cb9d0, 32'h3ea7a7ed} /* (3, 26, 27) {real, imag} */,
  {32'hbf0b1ac1, 32'hbf268040} /* (3, 26, 26) {real, imag} */,
  {32'h3c904cc0, 32'hbecb2459} /* (3, 26, 25) {real, imag} */,
  {32'hbe0237e0, 32'h3eddae3d} /* (3, 26, 24) {real, imag} */,
  {32'hbe3d4ef4, 32'hbf760b21} /* (3, 26, 23) {real, imag} */,
  {32'h3e86224c, 32'h3ee6339f} /* (3, 26, 22) {real, imag} */,
  {32'hbe3a49c6, 32'h3ef25f8d} /* (3, 26, 21) {real, imag} */,
  {32'hbea505c2, 32'h3da85200} /* (3, 26, 20) {real, imag} */,
  {32'h3da80080, 32'hbe2fcbaf} /* (3, 26, 19) {real, imag} */,
  {32'h3e1d5838, 32'hbf3da12e} /* (3, 26, 18) {real, imag} */,
  {32'h3df45eb3, 32'h3e82141e} /* (3, 26, 17) {real, imag} */,
  {32'hbdf7445e, 32'h3ed2bf78} /* (3, 26, 16) {real, imag} */,
  {32'h3e1d6b26, 32'h3e250f48} /* (3, 26, 15) {real, imag} */,
  {32'h3e4f3657, 32'hbd986a4f} /* (3, 26, 14) {real, imag} */,
  {32'hbe2cd20b, 32'hbf441508} /* (3, 26, 13) {real, imag} */,
  {32'h3e694d1f, 32'hbeb9d0e8} /* (3, 26, 12) {real, imag} */,
  {32'hbe546c24, 32'h3e8d787e} /* (3, 26, 11) {real, imag} */,
  {32'h3ec55666, 32'hbe32c313} /* (3, 26, 10) {real, imag} */,
  {32'h3ea2ae8b, 32'h3eaa042e} /* (3, 26, 9) {real, imag} */,
  {32'hbd9bb2cb, 32'h3dda1d24} /* (3, 26, 8) {real, imag} */,
  {32'h3d903a40, 32'h3f0ba4ee} /* (3, 26, 7) {real, imag} */,
  {32'h3e5357d8, 32'h3cc0b7dc} /* (3, 26, 6) {real, imag} */,
  {32'hbea7f426, 32'h3dfca9d5} /* (3, 26, 5) {real, imag} */,
  {32'hbede31f8, 32'h3f09fed7} /* (3, 26, 4) {real, imag} */,
  {32'h3db755d5, 32'h3f1f923e} /* (3, 26, 3) {real, imag} */,
  {32'hbe759d0a, 32'hbe00d8a4} /* (3, 26, 2) {real, imag} */,
  {32'h3f0875dc, 32'hbe597d12} /* (3, 26, 1) {real, imag} */,
  {32'h3e3fa0c0, 32'hbf121be8} /* (3, 26, 0) {real, imag} */,
  {32'hbf452674, 32'h3f2095c4} /* (3, 25, 31) {real, imag} */,
  {32'hbf339dd0, 32'hbf2ef548} /* (3, 25, 30) {real, imag} */,
  {32'h3dd5ab94, 32'hbe291b0c} /* (3, 25, 29) {real, imag} */,
  {32'hbed666ca, 32'h3edf1892} /* (3, 25, 28) {real, imag} */,
  {32'h3e8961e6, 32'hbe6e6ddc} /* (3, 25, 27) {real, imag} */,
  {32'h3d2db710, 32'h3ebeaf2e} /* (3, 25, 26) {real, imag} */,
  {32'h3e39ddc6, 32'hbe570a64} /* (3, 25, 25) {real, imag} */,
  {32'h3f0ac668, 32'hbdd2764f} /* (3, 25, 24) {real, imag} */,
  {32'hbdf6bb98, 32'hbe7452f5} /* (3, 25, 23) {real, imag} */,
  {32'hbea09473, 32'hbdac2a0b} /* (3, 25, 22) {real, imag} */,
  {32'h3d804150, 32'hbb8b8cc0} /* (3, 25, 21) {real, imag} */,
  {32'h3e1939c2, 32'hbe7bc9f3} /* (3, 25, 20) {real, imag} */,
  {32'hbd905cd0, 32'h3b6d7910} /* (3, 25, 19) {real, imag} */,
  {32'h3dbdb9ae, 32'h3eaccbce} /* (3, 25, 18) {real, imag} */,
  {32'h3e3acb01, 32'hbef99858} /* (3, 25, 17) {real, imag} */,
  {32'h3e1f9ba1, 32'hbe9d8b2c} /* (3, 25, 16) {real, imag} */,
  {32'h3e0ca606, 32'hbeb97b27} /* (3, 25, 15) {real, imag} */,
  {32'h3d6c73e0, 32'h3e8a1bdf} /* (3, 25, 14) {real, imag} */,
  {32'hbf40079e, 32'h3d2adafa} /* (3, 25, 13) {real, imag} */,
  {32'hbdbae56e, 32'h3f155723} /* (3, 25, 12) {real, imag} */,
  {32'hbf0273e0, 32'h3da4f8c4} /* (3, 25, 11) {real, imag} */,
  {32'h3f08a7ee, 32'h3dc88598} /* (3, 25, 10) {real, imag} */,
  {32'hbe8fae3d, 32'hbecca355} /* (3, 25, 9) {real, imag} */,
  {32'hbde1e0da, 32'hbeb689b2} /* (3, 25, 8) {real, imag} */,
  {32'h3ec3d47f, 32'h3e877fdc} /* (3, 25, 7) {real, imag} */,
  {32'h3c1838b8, 32'h3eee68dd} /* (3, 25, 6) {real, imag} */,
  {32'h3dff5c90, 32'hbf9a7570} /* (3, 25, 5) {real, imag} */,
  {32'h3e445caa, 32'h3ed8006a} /* (3, 25, 4) {real, imag} */,
  {32'hbeb6d1c1, 32'hbeb3ad58} /* (3, 25, 3) {real, imag} */,
  {32'hbf238152, 32'hbe911ebe} /* (3, 25, 2) {real, imag} */,
  {32'hbe6a2697, 32'hbe39e3f5} /* (3, 25, 1) {real, imag} */,
  {32'h3d001530, 32'h3f42fbc8} /* (3, 25, 0) {real, imag} */,
  {32'h3f568b2c, 32'hbeff3716} /* (3, 24, 31) {real, imag} */,
  {32'hbe7c8e74, 32'h3ee69e65} /* (3, 24, 30) {real, imag} */,
  {32'hbc39f5a0, 32'h3e4613e7} /* (3, 24, 29) {real, imag} */,
  {32'hbdbe2faa, 32'hbe7b362b} /* (3, 24, 28) {real, imag} */,
  {32'h3f05b43c, 32'hbec3507d} /* (3, 24, 27) {real, imag} */,
  {32'hbf1b7d94, 32'h3ee4ab5c} /* (3, 24, 26) {real, imag} */,
  {32'hbf2b1071, 32'h3d90b513} /* (3, 24, 25) {real, imag} */,
  {32'h3dfa66d0, 32'h3e0ae26a} /* (3, 24, 24) {real, imag} */,
  {32'hbf217df1, 32'h3ebeaa35} /* (3, 24, 23) {real, imag} */,
  {32'h3e47d849, 32'h3e6548f9} /* (3, 24, 22) {real, imag} */,
  {32'h3dd01dbe, 32'h3f2045ca} /* (3, 24, 21) {real, imag} */,
  {32'h3df2b496, 32'hbed4dd65} /* (3, 24, 20) {real, imag} */,
  {32'h3e6da44c, 32'hbec4359d} /* (3, 24, 19) {real, imag} */,
  {32'hbea46025, 32'hbeab1fb1} /* (3, 24, 18) {real, imag} */,
  {32'hbdc18874, 32'hbec77203} /* (3, 24, 17) {real, imag} */,
  {32'hbd924c6c, 32'h3e180376} /* (3, 24, 16) {real, imag} */,
  {32'hbe330534, 32'hbe2ee2ed} /* (3, 24, 15) {real, imag} */,
  {32'h3ef57653, 32'hbd384b90} /* (3, 24, 14) {real, imag} */,
  {32'h3eb8a4a5, 32'h3f12a83c} /* (3, 24, 13) {real, imag} */,
  {32'hbf1c18fc, 32'hbe39d0db} /* (3, 24, 12) {real, imag} */,
  {32'hbc1addd0, 32'hbe5a8a6c} /* (3, 24, 11) {real, imag} */,
  {32'hbf05e9a2, 32'h3ee119ce} /* (3, 24, 10) {real, imag} */,
  {32'h3dddffc0, 32'h3d23e08a} /* (3, 24, 9) {real, imag} */,
  {32'hbf0bd345, 32'hbdd3873a} /* (3, 24, 8) {real, imag} */,
  {32'hbda835a4, 32'hbf3efe2a} /* (3, 24, 7) {real, imag} */,
  {32'h3ea80922, 32'hbd9857fe} /* (3, 24, 6) {real, imag} */,
  {32'h3d653d38, 32'h3ebdca90} /* (3, 24, 5) {real, imag} */,
  {32'h3ec6c75a, 32'hbe7c48c6} /* (3, 24, 4) {real, imag} */,
  {32'hbebd730f, 32'hbd462678} /* (3, 24, 3) {real, imag} */,
  {32'hbf2f06e6, 32'h3e6b2454} /* (3, 24, 2) {real, imag} */,
  {32'h3f8a98e4, 32'hbf1fbb66} /* (3, 24, 1) {real, imag} */,
  {32'h3f7f2c6b, 32'h3d60d17c} /* (3, 24, 0) {real, imag} */,
  {32'hbf0a2e3a, 32'h3ebd4c96} /* (3, 23, 31) {real, imag} */,
  {32'hbf0768a5, 32'h3f05182e} /* (3, 23, 30) {real, imag} */,
  {32'hbe077ff0, 32'h3ddec512} /* (3, 23, 29) {real, imag} */,
  {32'h3e7902c4, 32'hbdd2e12c} /* (3, 23, 28) {real, imag} */,
  {32'hbe5d6d98, 32'h3ea4125c} /* (3, 23, 27) {real, imag} */,
  {32'hbdc90815, 32'hbe25dadb} /* (3, 23, 26) {real, imag} */,
  {32'hbec0ffb4, 32'hbe8b4001} /* (3, 23, 25) {real, imag} */,
  {32'h3e1b48cc, 32'h3ea5f5d1} /* (3, 23, 24) {real, imag} */,
  {32'hbee975fe, 32'hbe9809f4} /* (3, 23, 23) {real, imag} */,
  {32'h3edf4076, 32'h3e37cd06} /* (3, 23, 22) {real, imag} */,
  {32'hbe1ccdee, 32'hbe462345} /* (3, 23, 21) {real, imag} */,
  {32'h3df374ea, 32'h3e42124e} /* (3, 23, 20) {real, imag} */,
  {32'hbed5af34, 32'h3ef2dd10} /* (3, 23, 19) {real, imag} */,
  {32'hbeb393e2, 32'hbe822eb7} /* (3, 23, 18) {real, imag} */,
  {32'h3db444b7, 32'hbe7b7945} /* (3, 23, 17) {real, imag} */,
  {32'h3f0696a6, 32'h3dd04efe} /* (3, 23, 16) {real, imag} */,
  {32'h3debd1ce, 32'h3ef02bec} /* (3, 23, 15) {real, imag} */,
  {32'hbebbd9a7, 32'h3b9c6780} /* (3, 23, 14) {real, imag} */,
  {32'h3eab68ae, 32'h3ef1a71d} /* (3, 23, 13) {real, imag} */,
  {32'h3eb99065, 32'h3cfce810} /* (3, 23, 12) {real, imag} */,
  {32'h3f037697, 32'h3def8a92} /* (3, 23, 11) {real, imag} */,
  {32'hbe8ff34e, 32'h3e792fe1} /* (3, 23, 10) {real, imag} */,
  {32'hbf0533b4, 32'h3e62feb2} /* (3, 23, 9) {real, imag} */,
  {32'h3bcb6a20, 32'hbdfe1c7a} /* (3, 23, 8) {real, imag} */,
  {32'hbdf8b6cf, 32'h3ed8016a} /* (3, 23, 7) {real, imag} */,
  {32'h3eedaa92, 32'hbd203998} /* (3, 23, 6) {real, imag} */,
  {32'hbd87aff2, 32'hbeb06dee} /* (3, 23, 5) {real, imag} */,
  {32'h3ec195fe, 32'h3e937224} /* (3, 23, 4) {real, imag} */,
  {32'hbdcf9f44, 32'h3ef40dad} /* (3, 23, 3) {real, imag} */,
  {32'h3e7e2ed4, 32'hbf69e4d9} /* (3, 23, 2) {real, imag} */,
  {32'hbdd90cb8, 32'h3c9092f0} /* (3, 23, 1) {real, imag} */,
  {32'h3ccbb360, 32'h3ea76479} /* (3, 23, 0) {real, imag} */,
  {32'hbf200e12, 32'h3eee733d} /* (3, 22, 31) {real, imag} */,
  {32'h3e3e55c4, 32'hbe99704c} /* (3, 22, 30) {real, imag} */,
  {32'h3eebea81, 32'hbe308406} /* (3, 22, 29) {real, imag} */,
  {32'h3eda2cd6, 32'h3da1855c} /* (3, 22, 28) {real, imag} */,
  {32'h3e31154a, 32'h3b4fb480} /* (3, 22, 27) {real, imag} */,
  {32'hbe373321, 32'h3e2950ee} /* (3, 22, 26) {real, imag} */,
  {32'h3bb87920, 32'h3e6b6fb7} /* (3, 22, 25) {real, imag} */,
  {32'h3ba39060, 32'h3dbd7c9c} /* (3, 22, 24) {real, imag} */,
  {32'h3c97cc60, 32'hbd7ca512} /* (3, 22, 23) {real, imag} */,
  {32'hbe5ea870, 32'hbe8dac7f} /* (3, 22, 22) {real, imag} */,
  {32'hbdba28c2, 32'hbe5f49b6} /* (3, 22, 21) {real, imag} */,
  {32'hbeb81f01, 32'h3c3aef40} /* (3, 22, 20) {real, imag} */,
  {32'hbe73d368, 32'h3f41df08} /* (3, 22, 19) {real, imag} */,
  {32'h3f0268fe, 32'hbd6726d4} /* (3, 22, 18) {real, imag} */,
  {32'h3dc9b26c, 32'hbc8ceb3c} /* (3, 22, 17) {real, imag} */,
  {32'h3c6b55b0, 32'h3dcd061e} /* (3, 22, 16) {real, imag} */,
  {32'hbd5fd0fe, 32'h3f16e3be} /* (3, 22, 15) {real, imag} */,
  {32'hbedb6ddf, 32'h3eaf0b16} /* (3, 22, 14) {real, imag} */,
  {32'h3e9de6d0, 32'hbeaf7530} /* (3, 22, 13) {real, imag} */,
  {32'hbf4731b5, 32'hbecd33c6} /* (3, 22, 12) {real, imag} */,
  {32'hbd814bd8, 32'h3e94751e} /* (3, 22, 11) {real, imag} */,
  {32'h3dcf12ca, 32'hbe8a3227} /* (3, 22, 10) {real, imag} */,
  {32'h3ca421a8, 32'hbdd5a9bd} /* (3, 22, 9) {real, imag} */,
  {32'h3ec889e6, 32'hbe49cba8} /* (3, 22, 8) {real, imag} */,
  {32'hbd1fbf50, 32'hbe1f18fb} /* (3, 22, 7) {real, imag} */,
  {32'h3e8ce39a, 32'h3e257569} /* (3, 22, 6) {real, imag} */,
  {32'h3e10f64a, 32'h3da28e2c} /* (3, 22, 5) {real, imag} */,
  {32'hbe0f5abd, 32'hbf1291a7} /* (3, 22, 4) {real, imag} */,
  {32'h3bf74a40, 32'hbb97a280} /* (3, 22, 3) {real, imag} */,
  {32'hbd8a837a, 32'hbea0931d} /* (3, 22, 2) {real, imag} */,
  {32'h3de968bc, 32'h3e5c94ea} /* (3, 22, 1) {real, imag} */,
  {32'hbd2e8794, 32'h3eea89a4} /* (3, 22, 0) {real, imag} */,
  {32'hbe026c8d, 32'hbf117748} /* (3, 21, 31) {real, imag} */,
  {32'hbee8f55e, 32'h3e04d13a} /* (3, 21, 30) {real, imag} */,
  {32'h3b282cc0, 32'hbe751122} /* (3, 21, 29) {real, imag} */,
  {32'hbed3f8e0, 32'h3ee016bd} /* (3, 21, 28) {real, imag} */,
  {32'h3e9b4267, 32'h3f124668} /* (3, 21, 27) {real, imag} */,
  {32'hbd84b2d8, 32'h3c0ad390} /* (3, 21, 26) {real, imag} */,
  {32'hbdfa530d, 32'hbee73cd8} /* (3, 21, 25) {real, imag} */,
  {32'h3e71db52, 32'h3cfb5f10} /* (3, 21, 24) {real, imag} */,
  {32'hbeea7a37, 32'h3e337583} /* (3, 21, 23) {real, imag} */,
  {32'hbd0b2d10, 32'hbc76a790} /* (3, 21, 22) {real, imag} */,
  {32'h3e8ddda0, 32'hbe8c12f2} /* (3, 21, 21) {real, imag} */,
  {32'h3e318217, 32'h3e9a70ce} /* (3, 21, 20) {real, imag} */,
  {32'h3d13e7f0, 32'hbe83ec52} /* (3, 21, 19) {real, imag} */,
  {32'hbdcc2d51, 32'h3dd16b6c} /* (3, 21, 18) {real, imag} */,
  {32'h3e3a1630, 32'h3d964d2f} /* (3, 21, 17) {real, imag} */,
  {32'hbe34f2b6, 32'h3cf06112} /* (3, 21, 16) {real, imag} */,
  {32'h3f2bdfb8, 32'hbea05288} /* (3, 21, 15) {real, imag} */,
  {32'hbeec0ee8, 32'hbdf40bba} /* (3, 21, 14) {real, imag} */,
  {32'hbe238bd1, 32'h3f27837d} /* (3, 21, 13) {real, imag} */,
  {32'hbcfc7180, 32'h3f2cc6a0} /* (3, 21, 12) {real, imag} */,
  {32'h3de1972c, 32'hbe8a92a0} /* (3, 21, 11) {real, imag} */,
  {32'hbde347e0, 32'hbd3c25a0} /* (3, 21, 10) {real, imag} */,
  {32'hbdf967b4, 32'hbe0606eb} /* (3, 21, 9) {real, imag} */,
  {32'h3eb6aafc, 32'h3f42862e} /* (3, 21, 8) {real, imag} */,
  {32'h3ea4a3a4, 32'hbe47cd29} /* (3, 21, 7) {real, imag} */,
  {32'h3f0d698a, 32'hbef77fef} /* (3, 21, 6) {real, imag} */,
  {32'h3d47ecf0, 32'h3e2d23c4} /* (3, 21, 5) {real, imag} */,
  {32'hbea4719a, 32'h3e432178} /* (3, 21, 4) {real, imag} */,
  {32'hbef58f6c, 32'hbd51f008} /* (3, 21, 3) {real, imag} */,
  {32'hbeac15c8, 32'h3eed1399} /* (3, 21, 2) {real, imag} */,
  {32'h3e5d762a, 32'hbe3e8fb5} /* (3, 21, 1) {real, imag} */,
  {32'h3f26dd2d, 32'hbebaa684} /* (3, 21, 0) {real, imag} */,
  {32'h3e672c3d, 32'hbdcc8274} /* (3, 20, 31) {real, imag} */,
  {32'h3e6b3f40, 32'hbeab2879} /* (3, 20, 30) {real, imag} */,
  {32'hbd6df798, 32'hbe03d550} /* (3, 20, 29) {real, imag} */,
  {32'hbe2133c4, 32'hbd622198} /* (3, 20, 28) {real, imag} */,
  {32'h3e43ed76, 32'h3f32b0c6} /* (3, 20, 27) {real, imag} */,
  {32'h3de76a85, 32'hbdb5bac1} /* (3, 20, 26) {real, imag} */,
  {32'h3f418ee1, 32'hbcb43d30} /* (3, 20, 25) {real, imag} */,
  {32'hb9eb5400, 32'h3eb3360e} /* (3, 20, 24) {real, imag} */,
  {32'h3e9c4dce, 32'h3eee7aa6} /* (3, 20, 23) {real, imag} */,
  {32'hbe900bc9, 32'hbeac7909} /* (3, 20, 22) {real, imag} */,
  {32'h3e7e8c02, 32'h3e9a32da} /* (3, 20, 21) {real, imag} */,
  {32'hbe1226d4, 32'hbdc09794} /* (3, 20, 20) {real, imag} */,
  {32'h3ddab282, 32'h3edda2c4} /* (3, 20, 19) {real, imag} */,
  {32'h3e0eacf4, 32'hbe84159c} /* (3, 20, 18) {real, imag} */,
  {32'h3dd31b00, 32'h3f01cc01} /* (3, 20, 17) {real, imag} */,
  {32'h3c3e6c78, 32'hbe3a2447} /* (3, 20, 16) {real, imag} */,
  {32'hbe312852, 32'h3ded8388} /* (3, 20, 15) {real, imag} */,
  {32'h3c7a6198, 32'hbdc10f46} /* (3, 20, 14) {real, imag} */,
  {32'h3ccc4f93, 32'h3f296897} /* (3, 20, 13) {real, imag} */,
  {32'h3e5f4d6e, 32'h3e705337} /* (3, 20, 12) {real, imag} */,
  {32'hbe3f8e5c, 32'hbc5c39f0} /* (3, 20, 11) {real, imag} */,
  {32'hbec77fd7, 32'h3dce40b8} /* (3, 20, 10) {real, imag} */,
  {32'hbe3b21ac, 32'h3d62d5aa} /* (3, 20, 9) {real, imag} */,
  {32'hbdc6a1d0, 32'h3eacc927} /* (3, 20, 8) {real, imag} */,
  {32'hbe4b1d44, 32'h3f213274} /* (3, 20, 7) {real, imag} */,
  {32'hbea67c12, 32'hbe369909} /* (3, 20, 6) {real, imag} */,
  {32'hbe9420e1, 32'hbee72536} /* (3, 20, 5) {real, imag} */,
  {32'hbebd42d1, 32'hbe035657} /* (3, 20, 4) {real, imag} */,
  {32'h3f0d5465, 32'h3e5909fd} /* (3, 20, 3) {real, imag} */,
  {32'hbea4de64, 32'hbe1953b4} /* (3, 20, 2) {real, imag} */,
  {32'h3f189506, 32'hbdd33bcc} /* (3, 20, 1) {real, imag} */,
  {32'hbee5ed97, 32'hbe258766} /* (3, 20, 0) {real, imag} */,
  {32'h3da20d60, 32'h3dfb8b53} /* (3, 19, 31) {real, imag} */,
  {32'hbcd0e952, 32'hbdc6ecd6} /* (3, 19, 30) {real, imag} */,
  {32'h3e4a58db, 32'hbcd5ed54} /* (3, 19, 29) {real, imag} */,
  {32'h3e1364ce, 32'h3e82ab26} /* (3, 19, 28) {real, imag} */,
  {32'h3eccc968, 32'hbe9e8ad1} /* (3, 19, 27) {real, imag} */,
  {32'h3ecd4ec6, 32'h3d9f9374} /* (3, 19, 26) {real, imag} */,
  {32'h3e1b7cc4, 32'hbe2e12a2} /* (3, 19, 25) {real, imag} */,
  {32'h3c91b174, 32'h3cd13f20} /* (3, 19, 24) {real, imag} */,
  {32'hbef9c696, 32'h3d9f2d5e} /* (3, 19, 23) {real, imag} */,
  {32'h3e975b80, 32'hbe27ad02} /* (3, 19, 22) {real, imag} */,
  {32'hbe829d16, 32'hbe9c4ecd} /* (3, 19, 21) {real, imag} */,
  {32'h3f272f9d, 32'hbde0c1b2} /* (3, 19, 20) {real, imag} */,
  {32'hbe7ff44b, 32'h3e05812d} /* (3, 19, 19) {real, imag} */,
  {32'h3d8a2d0c, 32'h3db7e304} /* (3, 19, 18) {real, imag} */,
  {32'hbe22f203, 32'hbe059f36} /* (3, 19, 17) {real, imag} */,
  {32'hbeec9b28, 32'hbdaf9e58} /* (3, 19, 16) {real, imag} */,
  {32'h3e83c2ce, 32'h3ec36130} /* (3, 19, 15) {real, imag} */,
  {32'h3cae3de8, 32'h3ee93b55} /* (3, 19, 14) {real, imag} */,
  {32'h3f55f08d, 32'hbed070a7} /* (3, 19, 13) {real, imag} */,
  {32'hbedef586, 32'hbeab5ada} /* (3, 19, 12) {real, imag} */,
  {32'hbef13456, 32'hbe416c70} /* (3, 19, 11) {real, imag} */,
  {32'hbda468d6, 32'h3eb99afa} /* (3, 19, 10) {real, imag} */,
  {32'hbc8b7f00, 32'hbde78680} /* (3, 19, 9) {real, imag} */,
  {32'hbe8d8d51, 32'h3d18c112} /* (3, 19, 8) {real, imag} */,
  {32'h3edde473, 32'hbdeaba22} /* (3, 19, 7) {real, imag} */,
  {32'hbdb6bb0c, 32'hbf1814e9} /* (3, 19, 6) {real, imag} */,
  {32'hbdaaa1f5, 32'h3d8018ef} /* (3, 19, 5) {real, imag} */,
  {32'hbec6581c, 32'hbd8b62e6} /* (3, 19, 4) {real, imag} */,
  {32'hbd847644, 32'hbdcdd59c} /* (3, 19, 3) {real, imag} */,
  {32'h3c135290, 32'hbe2e7bbe} /* (3, 19, 2) {real, imag} */,
  {32'hbed5ed5b, 32'h3f03d542} /* (3, 19, 1) {real, imag} */,
  {32'hbdbd253c, 32'hbe58081f} /* (3, 19, 0) {real, imag} */,
  {32'h3e2ce9e7, 32'hbd29722c} /* (3, 18, 31) {real, imag} */,
  {32'h3cc785b0, 32'h3e02e060} /* (3, 18, 30) {real, imag} */,
  {32'h3eb17464, 32'h3e0d9fce} /* (3, 18, 29) {real, imag} */,
  {32'h3eed7627, 32'hbe88927c} /* (3, 18, 28) {real, imag} */,
  {32'h3e6cbd49, 32'h3eca0f1b} /* (3, 18, 27) {real, imag} */,
  {32'hbe351a2a, 32'h3eca6ea9} /* (3, 18, 26) {real, imag} */,
  {32'hbe66829c, 32'h3e98d21e} /* (3, 18, 25) {real, imag} */,
  {32'h3e582e92, 32'h3ea8e378} /* (3, 18, 24) {real, imag} */,
  {32'hbed35f4e, 32'h3c601300} /* (3, 18, 23) {real, imag} */,
  {32'hbed75152, 32'h3ed9f1fa} /* (3, 18, 22) {real, imag} */,
  {32'h3cd10c34, 32'hbe7bad0c} /* (3, 18, 21) {real, imag} */,
  {32'h3cd1e0e0, 32'hbd88a746} /* (3, 18, 20) {real, imag} */,
  {32'hbda4af24, 32'h3da28e50} /* (3, 18, 19) {real, imag} */,
  {32'h3e7157c9, 32'h3d0b86b6} /* (3, 18, 18) {real, imag} */,
  {32'h3eec00a6, 32'hbecc3e6e} /* (3, 18, 17) {real, imag} */,
  {32'h3e247b0c, 32'h3e13cb4f} /* (3, 18, 16) {real, imag} */,
  {32'hbe87bef5, 32'h3e14d477} /* (3, 18, 15) {real, imag} */,
  {32'h3e23a33c, 32'hbed62ba5} /* (3, 18, 14) {real, imag} */,
  {32'h3d4185ae, 32'h3e1884ea} /* (3, 18, 13) {real, imag} */,
  {32'h3f276336, 32'hbf477922} /* (3, 18, 12) {real, imag} */,
  {32'h3d101b8f, 32'hbe981124} /* (3, 18, 11) {real, imag} */,
  {32'h3d76e6ac, 32'h3e0bfcbe} /* (3, 18, 10) {real, imag} */,
  {32'hbd8068a2, 32'hbde08108} /* (3, 18, 9) {real, imag} */,
  {32'h3e47ef51, 32'hbf0742ab} /* (3, 18, 8) {real, imag} */,
  {32'hbda2908c, 32'hbdb44f16} /* (3, 18, 7) {real, imag} */,
  {32'hbd78c904, 32'h3d0ab0b0} /* (3, 18, 6) {real, imag} */,
  {32'hbdf78222, 32'h3dcaad2a} /* (3, 18, 5) {real, imag} */,
  {32'h3ef4c9a7, 32'hbd9d9d0c} /* (3, 18, 4) {real, imag} */,
  {32'h3dab9bd0, 32'h3e3b6606} /* (3, 18, 3) {real, imag} */,
  {32'hbec5518f, 32'h3ebca2c9} /* (3, 18, 2) {real, imag} */,
  {32'h3eda6b83, 32'hbea37c83} /* (3, 18, 1) {real, imag} */,
  {32'h3dcb75d9, 32'hbe8a9760} /* (3, 18, 0) {real, imag} */,
  {32'hbd82bef5, 32'h3db49e4c} /* (3, 17, 31) {real, imag} */,
  {32'h3d6fadc3, 32'hbeb4bf0e} /* (3, 17, 30) {real, imag} */,
  {32'hbed137ce, 32'h3e651844} /* (3, 17, 29) {real, imag} */,
  {32'h3e53fe81, 32'h3d6e4a48} /* (3, 17, 28) {real, imag} */,
  {32'hbdefb324, 32'hbdaeea3c} /* (3, 17, 27) {real, imag} */,
  {32'h3e5c1b06, 32'hbd425ea8} /* (3, 17, 26) {real, imag} */,
  {32'h3e62e9ca, 32'hbc152eb0} /* (3, 17, 25) {real, imag} */,
  {32'h3d992db4, 32'h3c1855c0} /* (3, 17, 24) {real, imag} */,
  {32'h3ea332ea, 32'h3c10d488} /* (3, 17, 23) {real, imag} */,
  {32'hbdef1fb4, 32'h3e21da3c} /* (3, 17, 22) {real, imag} */,
  {32'h3e032e79, 32'h3e5e422c} /* (3, 17, 21) {real, imag} */,
  {32'hbdeaae78, 32'hbe34fc42} /* (3, 17, 20) {real, imag} */,
  {32'h3d56a0ec, 32'h3ee3d199} /* (3, 17, 19) {real, imag} */,
  {32'h3d457dee, 32'hbf0fa455} /* (3, 17, 18) {real, imag} */,
  {32'hbc6e2838, 32'h3d4a274b} /* (3, 17, 17) {real, imag} */,
  {32'hbdd6c23e, 32'h3e3581cf} /* (3, 17, 16) {real, imag} */,
  {32'hbedece11, 32'hbedb097a} /* (3, 17, 15) {real, imag} */,
  {32'h3e651ebe, 32'h3e14fab6} /* (3, 17, 14) {real, imag} */,
  {32'hbdb6e076, 32'h3ba512b0} /* (3, 17, 13) {real, imag} */,
  {32'hbec4edd5, 32'h3dcd9698} /* (3, 17, 12) {real, imag} */,
  {32'hbd9921ea, 32'hbe7531c2} /* (3, 17, 11) {real, imag} */,
  {32'h3e9ffe01, 32'hbb013ec0} /* (3, 17, 10) {real, imag} */,
  {32'hbebf4e4a, 32'hbe711b7e} /* (3, 17, 9) {real, imag} */,
  {32'h3dbe3356, 32'hbedfb927} /* (3, 17, 8) {real, imag} */,
  {32'hbe5e7f50, 32'h3d75ffb2} /* (3, 17, 7) {real, imag} */,
  {32'h3d9b0ce0, 32'h3ee56b6a} /* (3, 17, 6) {real, imag} */,
  {32'hbd5c9790, 32'hbe2f4da0} /* (3, 17, 5) {real, imag} */,
  {32'h3e921fb2, 32'h3e345898} /* (3, 17, 4) {real, imag} */,
  {32'hbcd0c874, 32'hbea8899a} /* (3, 17, 3) {real, imag} */,
  {32'h3de1ce5c, 32'hbd28500f} /* (3, 17, 2) {real, imag} */,
  {32'h3dee6316, 32'h3e330d33} /* (3, 17, 1) {real, imag} */,
  {32'h3e9d0d19, 32'h3cbb022c} /* (3, 17, 0) {real, imag} */,
  {32'h3e696a10, 32'hbd0e7800} /* (3, 16, 31) {real, imag} */,
  {32'hbddf4384, 32'h3ebfe7be} /* (3, 16, 30) {real, imag} */,
  {32'hbcbbdfc6, 32'h3e6c09b6} /* (3, 16, 29) {real, imag} */,
  {32'h3dd361a9, 32'hbde01d82} /* (3, 16, 28) {real, imag} */,
  {32'hbe4e3961, 32'h3ee2aa68} /* (3, 16, 27) {real, imag} */,
  {32'h3e10e393, 32'hbeb53092} /* (3, 16, 26) {real, imag} */,
  {32'h3cbf0402, 32'h3dba76aa} /* (3, 16, 25) {real, imag} */,
  {32'h3dc66056, 32'h3c5ad700} /* (3, 16, 24) {real, imag} */,
  {32'h3e25d198, 32'h3dafe2c4} /* (3, 16, 23) {real, imag} */,
  {32'hbcaf0f28, 32'hbdb2d9fc} /* (3, 16, 22) {real, imag} */,
  {32'h3e8c88d6, 32'h3e46ed7c} /* (3, 16, 21) {real, imag} */,
  {32'h3dcb9e76, 32'h3eda6a7e} /* (3, 16, 20) {real, imag} */,
  {32'hbee9f72c, 32'h3d3227dd} /* (3, 16, 19) {real, imag} */,
  {32'hbe64fda0, 32'h3da0cc7e} /* (3, 16, 18) {real, imag} */,
  {32'hbe5f95d6, 32'h3e1c711d} /* (3, 16, 17) {real, imag} */,
  {32'hbdecc3a2, 32'h00000000} /* (3, 16, 16) {real, imag} */,
  {32'hbe5f95d6, 32'hbe1c711d} /* (3, 16, 15) {real, imag} */,
  {32'hbe64fda0, 32'hbda0cc7e} /* (3, 16, 14) {real, imag} */,
  {32'hbee9f72c, 32'hbd3227dd} /* (3, 16, 13) {real, imag} */,
  {32'h3dcb9e76, 32'hbeda6a7e} /* (3, 16, 12) {real, imag} */,
  {32'h3e8c88d6, 32'hbe46ed7c} /* (3, 16, 11) {real, imag} */,
  {32'hbcaf0f28, 32'h3db2d9fc} /* (3, 16, 10) {real, imag} */,
  {32'h3e25d198, 32'hbdafe2c4} /* (3, 16, 9) {real, imag} */,
  {32'h3dc66056, 32'hbc5ad700} /* (3, 16, 8) {real, imag} */,
  {32'h3cbf0402, 32'hbdba76aa} /* (3, 16, 7) {real, imag} */,
  {32'h3e10e393, 32'h3eb53092} /* (3, 16, 6) {real, imag} */,
  {32'hbe4e3961, 32'hbee2aa68} /* (3, 16, 5) {real, imag} */,
  {32'h3dd361a9, 32'h3de01d82} /* (3, 16, 4) {real, imag} */,
  {32'hbcbbdfc6, 32'hbe6c09b6} /* (3, 16, 3) {real, imag} */,
  {32'hbddf4384, 32'hbebfe7be} /* (3, 16, 2) {real, imag} */,
  {32'h3e696a10, 32'h3d0e7800} /* (3, 16, 1) {real, imag} */,
  {32'hbdd26ab0, 32'h00000000} /* (3, 16, 0) {real, imag} */,
  {32'h3dee6316, 32'hbe330d33} /* (3, 15, 31) {real, imag} */,
  {32'h3de1ce5c, 32'h3d28500f} /* (3, 15, 30) {real, imag} */,
  {32'hbcd0c874, 32'h3ea8899a} /* (3, 15, 29) {real, imag} */,
  {32'h3e921fb2, 32'hbe345898} /* (3, 15, 28) {real, imag} */,
  {32'hbd5c9790, 32'h3e2f4da0} /* (3, 15, 27) {real, imag} */,
  {32'h3d9b0ce0, 32'hbee56b6a} /* (3, 15, 26) {real, imag} */,
  {32'hbe5e7f50, 32'hbd75ffb2} /* (3, 15, 25) {real, imag} */,
  {32'h3dbe3356, 32'h3edfb927} /* (3, 15, 24) {real, imag} */,
  {32'hbebf4e4a, 32'h3e711b7e} /* (3, 15, 23) {real, imag} */,
  {32'h3e9ffe01, 32'h3b013ec0} /* (3, 15, 22) {real, imag} */,
  {32'hbd9921ea, 32'h3e7531c2} /* (3, 15, 21) {real, imag} */,
  {32'hbec4edd5, 32'hbdcd9698} /* (3, 15, 20) {real, imag} */,
  {32'hbdb6e076, 32'hbba512b0} /* (3, 15, 19) {real, imag} */,
  {32'h3e651ebe, 32'hbe14fab6} /* (3, 15, 18) {real, imag} */,
  {32'hbedece11, 32'h3edb097a} /* (3, 15, 17) {real, imag} */,
  {32'hbdd6c23e, 32'hbe3581cf} /* (3, 15, 16) {real, imag} */,
  {32'hbc6e2838, 32'hbd4a274b} /* (3, 15, 15) {real, imag} */,
  {32'h3d457dee, 32'h3f0fa455} /* (3, 15, 14) {real, imag} */,
  {32'h3d56a0ec, 32'hbee3d199} /* (3, 15, 13) {real, imag} */,
  {32'hbdeaae78, 32'h3e34fc42} /* (3, 15, 12) {real, imag} */,
  {32'h3e032e79, 32'hbe5e422c} /* (3, 15, 11) {real, imag} */,
  {32'hbdef1fb4, 32'hbe21da3c} /* (3, 15, 10) {real, imag} */,
  {32'h3ea332ea, 32'hbc10d488} /* (3, 15, 9) {real, imag} */,
  {32'h3d992db4, 32'hbc1855c0} /* (3, 15, 8) {real, imag} */,
  {32'h3e62e9ca, 32'h3c152eb0} /* (3, 15, 7) {real, imag} */,
  {32'h3e5c1b06, 32'h3d425ea8} /* (3, 15, 6) {real, imag} */,
  {32'hbdefb324, 32'h3daeea3c} /* (3, 15, 5) {real, imag} */,
  {32'h3e53fe81, 32'hbd6e4a48} /* (3, 15, 4) {real, imag} */,
  {32'hbed137ce, 32'hbe651844} /* (3, 15, 3) {real, imag} */,
  {32'h3d6fadc3, 32'h3eb4bf0e} /* (3, 15, 2) {real, imag} */,
  {32'hbd82bef5, 32'hbdb49e4c} /* (3, 15, 1) {real, imag} */,
  {32'h3e9d0d19, 32'hbcbb022c} /* (3, 15, 0) {real, imag} */,
  {32'h3eda6b83, 32'h3ea37c83} /* (3, 14, 31) {real, imag} */,
  {32'hbec5518f, 32'hbebca2c9} /* (3, 14, 30) {real, imag} */,
  {32'h3dab9bd0, 32'hbe3b6606} /* (3, 14, 29) {real, imag} */,
  {32'h3ef4c9a7, 32'h3d9d9d0c} /* (3, 14, 28) {real, imag} */,
  {32'hbdf78222, 32'hbdcaad2a} /* (3, 14, 27) {real, imag} */,
  {32'hbd78c904, 32'hbd0ab0b0} /* (3, 14, 26) {real, imag} */,
  {32'hbda2908c, 32'h3db44f16} /* (3, 14, 25) {real, imag} */,
  {32'h3e47ef51, 32'h3f0742ab} /* (3, 14, 24) {real, imag} */,
  {32'hbd8068a2, 32'h3de08108} /* (3, 14, 23) {real, imag} */,
  {32'h3d76e6ac, 32'hbe0bfcbe} /* (3, 14, 22) {real, imag} */,
  {32'h3d101b8f, 32'h3e981124} /* (3, 14, 21) {real, imag} */,
  {32'h3f276336, 32'h3f477922} /* (3, 14, 20) {real, imag} */,
  {32'h3d4185ae, 32'hbe1884ea} /* (3, 14, 19) {real, imag} */,
  {32'h3e23a33c, 32'h3ed62ba5} /* (3, 14, 18) {real, imag} */,
  {32'hbe87bef5, 32'hbe14d477} /* (3, 14, 17) {real, imag} */,
  {32'h3e247b0c, 32'hbe13cb4f} /* (3, 14, 16) {real, imag} */,
  {32'h3eec00a6, 32'h3ecc3e6e} /* (3, 14, 15) {real, imag} */,
  {32'h3e7157c9, 32'hbd0b86b6} /* (3, 14, 14) {real, imag} */,
  {32'hbda4af24, 32'hbda28e50} /* (3, 14, 13) {real, imag} */,
  {32'h3cd1e0e0, 32'h3d88a746} /* (3, 14, 12) {real, imag} */,
  {32'h3cd10c34, 32'h3e7bad0c} /* (3, 14, 11) {real, imag} */,
  {32'hbed75152, 32'hbed9f1fa} /* (3, 14, 10) {real, imag} */,
  {32'hbed35f4e, 32'hbc601300} /* (3, 14, 9) {real, imag} */,
  {32'h3e582e92, 32'hbea8e378} /* (3, 14, 8) {real, imag} */,
  {32'hbe66829c, 32'hbe98d21e} /* (3, 14, 7) {real, imag} */,
  {32'hbe351a2a, 32'hbeca6ea9} /* (3, 14, 6) {real, imag} */,
  {32'h3e6cbd49, 32'hbeca0f1b} /* (3, 14, 5) {real, imag} */,
  {32'h3eed7627, 32'h3e88927c} /* (3, 14, 4) {real, imag} */,
  {32'h3eb17464, 32'hbe0d9fce} /* (3, 14, 3) {real, imag} */,
  {32'h3cc785b0, 32'hbe02e060} /* (3, 14, 2) {real, imag} */,
  {32'h3e2ce9e7, 32'h3d29722c} /* (3, 14, 1) {real, imag} */,
  {32'h3dcb75d9, 32'h3e8a9760} /* (3, 14, 0) {real, imag} */,
  {32'hbed5ed5b, 32'hbf03d542} /* (3, 13, 31) {real, imag} */,
  {32'h3c135290, 32'h3e2e7bbe} /* (3, 13, 30) {real, imag} */,
  {32'hbd847644, 32'h3dcdd59c} /* (3, 13, 29) {real, imag} */,
  {32'hbec6581c, 32'h3d8b62e6} /* (3, 13, 28) {real, imag} */,
  {32'hbdaaa1f5, 32'hbd8018ef} /* (3, 13, 27) {real, imag} */,
  {32'hbdb6bb0c, 32'h3f1814e9} /* (3, 13, 26) {real, imag} */,
  {32'h3edde473, 32'h3deaba22} /* (3, 13, 25) {real, imag} */,
  {32'hbe8d8d51, 32'hbd18c112} /* (3, 13, 24) {real, imag} */,
  {32'hbc8b7f00, 32'h3de78680} /* (3, 13, 23) {real, imag} */,
  {32'hbda468d6, 32'hbeb99afa} /* (3, 13, 22) {real, imag} */,
  {32'hbef13456, 32'h3e416c70} /* (3, 13, 21) {real, imag} */,
  {32'hbedef586, 32'h3eab5ada} /* (3, 13, 20) {real, imag} */,
  {32'h3f55f08d, 32'h3ed070a7} /* (3, 13, 19) {real, imag} */,
  {32'h3cae3de8, 32'hbee93b55} /* (3, 13, 18) {real, imag} */,
  {32'h3e83c2ce, 32'hbec36130} /* (3, 13, 17) {real, imag} */,
  {32'hbeec9b28, 32'h3daf9e58} /* (3, 13, 16) {real, imag} */,
  {32'hbe22f203, 32'h3e059f36} /* (3, 13, 15) {real, imag} */,
  {32'h3d8a2d0c, 32'hbdb7e304} /* (3, 13, 14) {real, imag} */,
  {32'hbe7ff44b, 32'hbe05812d} /* (3, 13, 13) {real, imag} */,
  {32'h3f272f9d, 32'h3de0c1b2} /* (3, 13, 12) {real, imag} */,
  {32'hbe829d16, 32'h3e9c4ecd} /* (3, 13, 11) {real, imag} */,
  {32'h3e975b80, 32'h3e27ad02} /* (3, 13, 10) {real, imag} */,
  {32'hbef9c696, 32'hbd9f2d5e} /* (3, 13, 9) {real, imag} */,
  {32'h3c91b174, 32'hbcd13f20} /* (3, 13, 8) {real, imag} */,
  {32'h3e1b7cc4, 32'h3e2e12a2} /* (3, 13, 7) {real, imag} */,
  {32'h3ecd4ec6, 32'hbd9f9374} /* (3, 13, 6) {real, imag} */,
  {32'h3eccc968, 32'h3e9e8ad1} /* (3, 13, 5) {real, imag} */,
  {32'h3e1364ce, 32'hbe82ab26} /* (3, 13, 4) {real, imag} */,
  {32'h3e4a58db, 32'h3cd5ed54} /* (3, 13, 3) {real, imag} */,
  {32'hbcd0e952, 32'h3dc6ecd6} /* (3, 13, 2) {real, imag} */,
  {32'h3da20d60, 32'hbdfb8b53} /* (3, 13, 1) {real, imag} */,
  {32'hbdbd253c, 32'h3e58081f} /* (3, 13, 0) {real, imag} */,
  {32'h3f189506, 32'h3dd33bcc} /* (3, 12, 31) {real, imag} */,
  {32'hbea4de64, 32'h3e1953b4} /* (3, 12, 30) {real, imag} */,
  {32'h3f0d5465, 32'hbe5909fd} /* (3, 12, 29) {real, imag} */,
  {32'hbebd42d1, 32'h3e035657} /* (3, 12, 28) {real, imag} */,
  {32'hbe9420e1, 32'h3ee72536} /* (3, 12, 27) {real, imag} */,
  {32'hbea67c12, 32'h3e369909} /* (3, 12, 26) {real, imag} */,
  {32'hbe4b1d44, 32'hbf213274} /* (3, 12, 25) {real, imag} */,
  {32'hbdc6a1d0, 32'hbeacc927} /* (3, 12, 24) {real, imag} */,
  {32'hbe3b21ac, 32'hbd62d5aa} /* (3, 12, 23) {real, imag} */,
  {32'hbec77fd7, 32'hbdce40b8} /* (3, 12, 22) {real, imag} */,
  {32'hbe3f8e5c, 32'h3c5c39f0} /* (3, 12, 21) {real, imag} */,
  {32'h3e5f4d6e, 32'hbe705337} /* (3, 12, 20) {real, imag} */,
  {32'h3ccc4f93, 32'hbf296897} /* (3, 12, 19) {real, imag} */,
  {32'h3c7a6198, 32'h3dc10f46} /* (3, 12, 18) {real, imag} */,
  {32'hbe312852, 32'hbded8388} /* (3, 12, 17) {real, imag} */,
  {32'h3c3e6c78, 32'h3e3a2447} /* (3, 12, 16) {real, imag} */,
  {32'h3dd31b00, 32'hbf01cc01} /* (3, 12, 15) {real, imag} */,
  {32'h3e0eacf4, 32'h3e84159c} /* (3, 12, 14) {real, imag} */,
  {32'h3ddab282, 32'hbedda2c4} /* (3, 12, 13) {real, imag} */,
  {32'hbe1226d4, 32'h3dc09794} /* (3, 12, 12) {real, imag} */,
  {32'h3e7e8c02, 32'hbe9a32da} /* (3, 12, 11) {real, imag} */,
  {32'hbe900bc9, 32'h3eac7909} /* (3, 12, 10) {real, imag} */,
  {32'h3e9c4dce, 32'hbeee7aa6} /* (3, 12, 9) {real, imag} */,
  {32'hb9eb5400, 32'hbeb3360e} /* (3, 12, 8) {real, imag} */,
  {32'h3f418ee1, 32'h3cb43d30} /* (3, 12, 7) {real, imag} */,
  {32'h3de76a85, 32'h3db5bac1} /* (3, 12, 6) {real, imag} */,
  {32'h3e43ed76, 32'hbf32b0c6} /* (3, 12, 5) {real, imag} */,
  {32'hbe2133c4, 32'h3d622198} /* (3, 12, 4) {real, imag} */,
  {32'hbd6df798, 32'h3e03d550} /* (3, 12, 3) {real, imag} */,
  {32'h3e6b3f40, 32'h3eab2879} /* (3, 12, 2) {real, imag} */,
  {32'h3e672c3d, 32'h3dcc8274} /* (3, 12, 1) {real, imag} */,
  {32'hbee5ed97, 32'h3e258766} /* (3, 12, 0) {real, imag} */,
  {32'h3e5d762a, 32'h3e3e8fb5} /* (3, 11, 31) {real, imag} */,
  {32'hbeac15c8, 32'hbeed1399} /* (3, 11, 30) {real, imag} */,
  {32'hbef58f6c, 32'h3d51f008} /* (3, 11, 29) {real, imag} */,
  {32'hbea4719a, 32'hbe432178} /* (3, 11, 28) {real, imag} */,
  {32'h3d47ecf0, 32'hbe2d23c4} /* (3, 11, 27) {real, imag} */,
  {32'h3f0d698a, 32'h3ef77fef} /* (3, 11, 26) {real, imag} */,
  {32'h3ea4a3a4, 32'h3e47cd29} /* (3, 11, 25) {real, imag} */,
  {32'h3eb6aafc, 32'hbf42862e} /* (3, 11, 24) {real, imag} */,
  {32'hbdf967b4, 32'h3e0606eb} /* (3, 11, 23) {real, imag} */,
  {32'hbde347e0, 32'h3d3c25a0} /* (3, 11, 22) {real, imag} */,
  {32'h3de1972c, 32'h3e8a92a0} /* (3, 11, 21) {real, imag} */,
  {32'hbcfc7180, 32'hbf2cc6a0} /* (3, 11, 20) {real, imag} */,
  {32'hbe238bd1, 32'hbf27837d} /* (3, 11, 19) {real, imag} */,
  {32'hbeec0ee8, 32'h3df40bba} /* (3, 11, 18) {real, imag} */,
  {32'h3f2bdfb8, 32'h3ea05288} /* (3, 11, 17) {real, imag} */,
  {32'hbe34f2b6, 32'hbcf06112} /* (3, 11, 16) {real, imag} */,
  {32'h3e3a1630, 32'hbd964d2f} /* (3, 11, 15) {real, imag} */,
  {32'hbdcc2d51, 32'hbdd16b6c} /* (3, 11, 14) {real, imag} */,
  {32'h3d13e7f0, 32'h3e83ec52} /* (3, 11, 13) {real, imag} */,
  {32'h3e318217, 32'hbe9a70ce} /* (3, 11, 12) {real, imag} */,
  {32'h3e8ddda0, 32'h3e8c12f2} /* (3, 11, 11) {real, imag} */,
  {32'hbd0b2d10, 32'h3c76a790} /* (3, 11, 10) {real, imag} */,
  {32'hbeea7a37, 32'hbe337583} /* (3, 11, 9) {real, imag} */,
  {32'h3e71db52, 32'hbcfb5f10} /* (3, 11, 8) {real, imag} */,
  {32'hbdfa530d, 32'h3ee73cd8} /* (3, 11, 7) {real, imag} */,
  {32'hbd84b2d8, 32'hbc0ad390} /* (3, 11, 6) {real, imag} */,
  {32'h3e9b4267, 32'hbf124668} /* (3, 11, 5) {real, imag} */,
  {32'hbed3f8e0, 32'hbee016bd} /* (3, 11, 4) {real, imag} */,
  {32'h3b282cc0, 32'h3e751122} /* (3, 11, 3) {real, imag} */,
  {32'hbee8f55e, 32'hbe04d13a} /* (3, 11, 2) {real, imag} */,
  {32'hbe026c8d, 32'h3f117748} /* (3, 11, 1) {real, imag} */,
  {32'h3f26dd2d, 32'h3ebaa684} /* (3, 11, 0) {real, imag} */,
  {32'h3de968bc, 32'hbe5c94ea} /* (3, 10, 31) {real, imag} */,
  {32'hbd8a837a, 32'h3ea0931d} /* (3, 10, 30) {real, imag} */,
  {32'h3bf74a40, 32'h3b97a280} /* (3, 10, 29) {real, imag} */,
  {32'hbe0f5abd, 32'h3f1291a7} /* (3, 10, 28) {real, imag} */,
  {32'h3e10f64a, 32'hbda28e2c} /* (3, 10, 27) {real, imag} */,
  {32'h3e8ce39a, 32'hbe257569} /* (3, 10, 26) {real, imag} */,
  {32'hbd1fbf50, 32'h3e1f18fb} /* (3, 10, 25) {real, imag} */,
  {32'h3ec889e6, 32'h3e49cba8} /* (3, 10, 24) {real, imag} */,
  {32'h3ca421a8, 32'h3dd5a9bd} /* (3, 10, 23) {real, imag} */,
  {32'h3dcf12ca, 32'h3e8a3227} /* (3, 10, 22) {real, imag} */,
  {32'hbd814bd8, 32'hbe94751e} /* (3, 10, 21) {real, imag} */,
  {32'hbf4731b5, 32'h3ecd33c6} /* (3, 10, 20) {real, imag} */,
  {32'h3e9de6d0, 32'h3eaf7530} /* (3, 10, 19) {real, imag} */,
  {32'hbedb6ddf, 32'hbeaf0b16} /* (3, 10, 18) {real, imag} */,
  {32'hbd5fd0fe, 32'hbf16e3be} /* (3, 10, 17) {real, imag} */,
  {32'h3c6b55b0, 32'hbdcd061e} /* (3, 10, 16) {real, imag} */,
  {32'h3dc9b26c, 32'h3c8ceb3c} /* (3, 10, 15) {real, imag} */,
  {32'h3f0268fe, 32'h3d6726d4} /* (3, 10, 14) {real, imag} */,
  {32'hbe73d368, 32'hbf41df08} /* (3, 10, 13) {real, imag} */,
  {32'hbeb81f01, 32'hbc3aef40} /* (3, 10, 12) {real, imag} */,
  {32'hbdba28c2, 32'h3e5f49b6} /* (3, 10, 11) {real, imag} */,
  {32'hbe5ea870, 32'h3e8dac7f} /* (3, 10, 10) {real, imag} */,
  {32'h3c97cc60, 32'h3d7ca512} /* (3, 10, 9) {real, imag} */,
  {32'h3ba39060, 32'hbdbd7c9c} /* (3, 10, 8) {real, imag} */,
  {32'h3bb87920, 32'hbe6b6fb7} /* (3, 10, 7) {real, imag} */,
  {32'hbe373321, 32'hbe2950ee} /* (3, 10, 6) {real, imag} */,
  {32'h3e31154a, 32'hbb4fb480} /* (3, 10, 5) {real, imag} */,
  {32'h3eda2cd6, 32'hbda1855c} /* (3, 10, 4) {real, imag} */,
  {32'h3eebea81, 32'h3e308406} /* (3, 10, 3) {real, imag} */,
  {32'h3e3e55c4, 32'h3e99704c} /* (3, 10, 2) {real, imag} */,
  {32'hbf200e12, 32'hbeee733d} /* (3, 10, 1) {real, imag} */,
  {32'hbd2e8794, 32'hbeea89a4} /* (3, 10, 0) {real, imag} */,
  {32'hbdd90cb8, 32'hbc9092f0} /* (3, 9, 31) {real, imag} */,
  {32'h3e7e2ed4, 32'h3f69e4d9} /* (3, 9, 30) {real, imag} */,
  {32'hbdcf9f44, 32'hbef40dad} /* (3, 9, 29) {real, imag} */,
  {32'h3ec195fe, 32'hbe937224} /* (3, 9, 28) {real, imag} */,
  {32'hbd87aff2, 32'h3eb06dee} /* (3, 9, 27) {real, imag} */,
  {32'h3eedaa92, 32'h3d203998} /* (3, 9, 26) {real, imag} */,
  {32'hbdf8b6cf, 32'hbed8016a} /* (3, 9, 25) {real, imag} */,
  {32'h3bcb6a20, 32'h3dfe1c7a} /* (3, 9, 24) {real, imag} */,
  {32'hbf0533b4, 32'hbe62feb2} /* (3, 9, 23) {real, imag} */,
  {32'hbe8ff34e, 32'hbe792fe1} /* (3, 9, 22) {real, imag} */,
  {32'h3f037697, 32'hbdef8a92} /* (3, 9, 21) {real, imag} */,
  {32'h3eb99065, 32'hbcfce810} /* (3, 9, 20) {real, imag} */,
  {32'h3eab68ae, 32'hbef1a71d} /* (3, 9, 19) {real, imag} */,
  {32'hbebbd9a7, 32'hbb9c6780} /* (3, 9, 18) {real, imag} */,
  {32'h3debd1ce, 32'hbef02bec} /* (3, 9, 17) {real, imag} */,
  {32'h3f0696a6, 32'hbdd04efe} /* (3, 9, 16) {real, imag} */,
  {32'h3db444b7, 32'h3e7b7945} /* (3, 9, 15) {real, imag} */,
  {32'hbeb393e2, 32'h3e822eb7} /* (3, 9, 14) {real, imag} */,
  {32'hbed5af34, 32'hbef2dd10} /* (3, 9, 13) {real, imag} */,
  {32'h3df374ea, 32'hbe42124e} /* (3, 9, 12) {real, imag} */,
  {32'hbe1ccdee, 32'h3e462345} /* (3, 9, 11) {real, imag} */,
  {32'h3edf4076, 32'hbe37cd06} /* (3, 9, 10) {real, imag} */,
  {32'hbee975fe, 32'h3e9809f4} /* (3, 9, 9) {real, imag} */,
  {32'h3e1b48cc, 32'hbea5f5d1} /* (3, 9, 8) {real, imag} */,
  {32'hbec0ffb4, 32'h3e8b4001} /* (3, 9, 7) {real, imag} */,
  {32'hbdc90815, 32'h3e25dadb} /* (3, 9, 6) {real, imag} */,
  {32'hbe5d6d98, 32'hbea4125c} /* (3, 9, 5) {real, imag} */,
  {32'h3e7902c4, 32'h3dd2e12c} /* (3, 9, 4) {real, imag} */,
  {32'hbe077ff0, 32'hbddec512} /* (3, 9, 3) {real, imag} */,
  {32'hbf0768a5, 32'hbf05182e} /* (3, 9, 2) {real, imag} */,
  {32'hbf0a2e3a, 32'hbebd4c96} /* (3, 9, 1) {real, imag} */,
  {32'h3ccbb360, 32'hbea76479} /* (3, 9, 0) {real, imag} */,
  {32'h3f8a98e4, 32'h3f1fbb66} /* (3, 8, 31) {real, imag} */,
  {32'hbf2f06e6, 32'hbe6b2454} /* (3, 8, 30) {real, imag} */,
  {32'hbebd730f, 32'h3d462678} /* (3, 8, 29) {real, imag} */,
  {32'h3ec6c75a, 32'h3e7c48c6} /* (3, 8, 28) {real, imag} */,
  {32'h3d653d38, 32'hbebdca90} /* (3, 8, 27) {real, imag} */,
  {32'h3ea80922, 32'h3d9857fe} /* (3, 8, 26) {real, imag} */,
  {32'hbda835a4, 32'h3f3efe2a} /* (3, 8, 25) {real, imag} */,
  {32'hbf0bd345, 32'h3dd3873a} /* (3, 8, 24) {real, imag} */,
  {32'h3dddffc0, 32'hbd23e08a} /* (3, 8, 23) {real, imag} */,
  {32'hbf05e9a2, 32'hbee119ce} /* (3, 8, 22) {real, imag} */,
  {32'hbc1addd0, 32'h3e5a8a6c} /* (3, 8, 21) {real, imag} */,
  {32'hbf1c18fc, 32'h3e39d0db} /* (3, 8, 20) {real, imag} */,
  {32'h3eb8a4a5, 32'hbf12a83c} /* (3, 8, 19) {real, imag} */,
  {32'h3ef57653, 32'h3d384b90} /* (3, 8, 18) {real, imag} */,
  {32'hbe330534, 32'h3e2ee2ed} /* (3, 8, 17) {real, imag} */,
  {32'hbd924c6c, 32'hbe180376} /* (3, 8, 16) {real, imag} */,
  {32'hbdc18874, 32'h3ec77203} /* (3, 8, 15) {real, imag} */,
  {32'hbea46025, 32'h3eab1fb1} /* (3, 8, 14) {real, imag} */,
  {32'h3e6da44c, 32'h3ec4359d} /* (3, 8, 13) {real, imag} */,
  {32'h3df2b496, 32'h3ed4dd65} /* (3, 8, 12) {real, imag} */,
  {32'h3dd01dbe, 32'hbf2045ca} /* (3, 8, 11) {real, imag} */,
  {32'h3e47d849, 32'hbe6548f9} /* (3, 8, 10) {real, imag} */,
  {32'hbf217df1, 32'hbebeaa35} /* (3, 8, 9) {real, imag} */,
  {32'h3dfa66d0, 32'hbe0ae26a} /* (3, 8, 8) {real, imag} */,
  {32'hbf2b1071, 32'hbd90b513} /* (3, 8, 7) {real, imag} */,
  {32'hbf1b7d94, 32'hbee4ab5c} /* (3, 8, 6) {real, imag} */,
  {32'h3f05b43c, 32'h3ec3507d} /* (3, 8, 5) {real, imag} */,
  {32'hbdbe2faa, 32'h3e7b362b} /* (3, 8, 4) {real, imag} */,
  {32'hbc39f5a0, 32'hbe4613e7} /* (3, 8, 3) {real, imag} */,
  {32'hbe7c8e74, 32'hbee69e65} /* (3, 8, 2) {real, imag} */,
  {32'h3f568b2c, 32'h3eff3716} /* (3, 8, 1) {real, imag} */,
  {32'h3f7f2c6b, 32'hbd60d17c} /* (3, 8, 0) {real, imag} */,
  {32'hbe6a2697, 32'h3e39e3f5} /* (3, 7, 31) {real, imag} */,
  {32'hbf238152, 32'h3e911ebe} /* (3, 7, 30) {real, imag} */,
  {32'hbeb6d1c1, 32'h3eb3ad58} /* (3, 7, 29) {real, imag} */,
  {32'h3e445caa, 32'hbed8006a} /* (3, 7, 28) {real, imag} */,
  {32'h3dff5c90, 32'h3f9a7570} /* (3, 7, 27) {real, imag} */,
  {32'h3c1838b8, 32'hbeee68dd} /* (3, 7, 26) {real, imag} */,
  {32'h3ec3d47f, 32'hbe877fdc} /* (3, 7, 25) {real, imag} */,
  {32'hbde1e0da, 32'h3eb689b2} /* (3, 7, 24) {real, imag} */,
  {32'hbe8fae3d, 32'h3ecca355} /* (3, 7, 23) {real, imag} */,
  {32'h3f08a7ee, 32'hbdc88598} /* (3, 7, 22) {real, imag} */,
  {32'hbf0273e0, 32'hbda4f8c4} /* (3, 7, 21) {real, imag} */,
  {32'hbdbae56e, 32'hbf155723} /* (3, 7, 20) {real, imag} */,
  {32'hbf40079e, 32'hbd2adafa} /* (3, 7, 19) {real, imag} */,
  {32'h3d6c73e0, 32'hbe8a1bdf} /* (3, 7, 18) {real, imag} */,
  {32'h3e0ca606, 32'h3eb97b27} /* (3, 7, 17) {real, imag} */,
  {32'h3e1f9ba1, 32'h3e9d8b2c} /* (3, 7, 16) {real, imag} */,
  {32'h3e3acb01, 32'h3ef99858} /* (3, 7, 15) {real, imag} */,
  {32'h3dbdb9ae, 32'hbeaccbce} /* (3, 7, 14) {real, imag} */,
  {32'hbd905cd0, 32'hbb6d7910} /* (3, 7, 13) {real, imag} */,
  {32'h3e1939c2, 32'h3e7bc9f3} /* (3, 7, 12) {real, imag} */,
  {32'h3d804150, 32'h3b8b8cc0} /* (3, 7, 11) {real, imag} */,
  {32'hbea09473, 32'h3dac2a0b} /* (3, 7, 10) {real, imag} */,
  {32'hbdf6bb98, 32'h3e7452f5} /* (3, 7, 9) {real, imag} */,
  {32'h3f0ac668, 32'h3dd2764f} /* (3, 7, 8) {real, imag} */,
  {32'h3e39ddc6, 32'h3e570a64} /* (3, 7, 7) {real, imag} */,
  {32'h3d2db710, 32'hbebeaf2e} /* (3, 7, 6) {real, imag} */,
  {32'h3e8961e6, 32'h3e6e6ddc} /* (3, 7, 5) {real, imag} */,
  {32'hbed666ca, 32'hbedf1892} /* (3, 7, 4) {real, imag} */,
  {32'h3dd5ab94, 32'h3e291b0c} /* (3, 7, 3) {real, imag} */,
  {32'hbf339dd0, 32'h3f2ef548} /* (3, 7, 2) {real, imag} */,
  {32'hbf452674, 32'hbf2095c4} /* (3, 7, 1) {real, imag} */,
  {32'h3d001530, 32'hbf42fbc8} /* (3, 7, 0) {real, imag} */,
  {32'h3f0875dc, 32'h3e597d12} /* (3, 6, 31) {real, imag} */,
  {32'hbe759d0a, 32'h3e00d8a4} /* (3, 6, 30) {real, imag} */,
  {32'h3db755d5, 32'hbf1f923e} /* (3, 6, 29) {real, imag} */,
  {32'hbede31f8, 32'hbf09fed7} /* (3, 6, 28) {real, imag} */,
  {32'hbea7f426, 32'hbdfca9d5} /* (3, 6, 27) {real, imag} */,
  {32'h3e5357d8, 32'hbcc0b7dc} /* (3, 6, 26) {real, imag} */,
  {32'h3d903a40, 32'hbf0ba4ee} /* (3, 6, 25) {real, imag} */,
  {32'hbd9bb2cb, 32'hbdda1d24} /* (3, 6, 24) {real, imag} */,
  {32'h3ea2ae8b, 32'hbeaa042e} /* (3, 6, 23) {real, imag} */,
  {32'h3ec55666, 32'h3e32c313} /* (3, 6, 22) {real, imag} */,
  {32'hbe546c24, 32'hbe8d787e} /* (3, 6, 21) {real, imag} */,
  {32'h3e694d1f, 32'h3eb9d0e8} /* (3, 6, 20) {real, imag} */,
  {32'hbe2cd20b, 32'h3f441508} /* (3, 6, 19) {real, imag} */,
  {32'h3e4f3657, 32'h3d986a4f} /* (3, 6, 18) {real, imag} */,
  {32'h3e1d6b26, 32'hbe250f48} /* (3, 6, 17) {real, imag} */,
  {32'hbdf7445e, 32'hbed2bf78} /* (3, 6, 16) {real, imag} */,
  {32'h3df45eb3, 32'hbe82141e} /* (3, 6, 15) {real, imag} */,
  {32'h3e1d5838, 32'h3f3da12e} /* (3, 6, 14) {real, imag} */,
  {32'h3da80080, 32'h3e2fcbaf} /* (3, 6, 13) {real, imag} */,
  {32'hbea505c2, 32'hbda85200} /* (3, 6, 12) {real, imag} */,
  {32'hbe3a49c6, 32'hbef25f8d} /* (3, 6, 11) {real, imag} */,
  {32'h3e86224c, 32'hbee6339f} /* (3, 6, 10) {real, imag} */,
  {32'hbe3d4ef4, 32'h3f760b21} /* (3, 6, 9) {real, imag} */,
  {32'hbe0237e0, 32'hbeddae3d} /* (3, 6, 8) {real, imag} */,
  {32'h3c904cc0, 32'h3ecb2459} /* (3, 6, 7) {real, imag} */,
  {32'hbf0b1ac1, 32'h3f268040} /* (3, 6, 6) {real, imag} */,
  {32'hbe8cb9d0, 32'hbea7a7ed} /* (3, 6, 5) {real, imag} */,
  {32'h3e46cade, 32'hbe2d7ddf} /* (3, 6, 4) {real, imag} */,
  {32'hbdf85086, 32'h3e8f9a78} /* (3, 6, 3) {real, imag} */,
  {32'hbf39221e, 32'h3ecae763} /* (3, 6, 2) {real, imag} */,
  {32'h3f399064, 32'hbee206e8} /* (3, 6, 1) {real, imag} */,
  {32'h3e3fa0c0, 32'h3f121be8} /* (3, 6, 0) {real, imag} */,
  {32'h40158132, 32'hbe9695ba} /* (3, 5, 31) {real, imag} */,
  {32'hbf98ac70, 32'h3df8793c} /* (3, 5, 30) {real, imag} */,
  {32'hbf101288, 32'hbe9af5fe} /* (3, 5, 29) {real, imag} */,
  {32'h3ec839a4, 32'hbf53533c} /* (3, 5, 28) {real, imag} */,
  {32'hbf52a943, 32'hbb906940} /* (3, 5, 27) {real, imag} */,
  {32'h3ddb8fba, 32'hbe3f3041} /* (3, 5, 26) {real, imag} */,
  {32'h3eb2d7c6, 32'h3eaab2f3} /* (3, 5, 25) {real, imag} */,
  {32'hbed1bd33, 32'h3db87ddf} /* (3, 5, 24) {real, imag} */,
  {32'hbd3c3498, 32'hbd8fd190} /* (3, 5, 23) {real, imag} */,
  {32'hbeeb317b, 32'h3e8f51a2} /* (3, 5, 22) {real, imag} */,
  {32'hbf3fe3c3, 32'h3e66d764} /* (3, 5, 21) {real, imag} */,
  {32'h3d93a400, 32'h3e88234e} /* (3, 5, 20) {real, imag} */,
  {32'hbbc7bff0, 32'h3c262428} /* (3, 5, 19) {real, imag} */,
  {32'hbedc369e, 32'hbe4a5b06} /* (3, 5, 18) {real, imag} */,
  {32'hbc858400, 32'hbdb7161f} /* (3, 5, 17) {real, imag} */,
  {32'hbeb116d6, 32'h3db16ca3} /* (3, 5, 16) {real, imag} */,
  {32'hbd75f7d0, 32'hbf208712} /* (3, 5, 15) {real, imag} */,
  {32'h3d10a7da, 32'hbdbcb9af} /* (3, 5, 14) {real, imag} */,
  {32'h3e06db1a, 32'hbef70352} /* (3, 5, 13) {real, imag} */,
  {32'hbdf7577a, 32'h3dc62f58} /* (3, 5, 12) {real, imag} */,
  {32'hbe3d1e5c, 32'hbec81b5c} /* (3, 5, 11) {real, imag} */,
  {32'h3e801ca2, 32'hbe3adf63} /* (3, 5, 10) {real, imag} */,
  {32'h3f292b9c, 32'h3e5e24e6} /* (3, 5, 9) {real, imag} */,
  {32'hbe26f0f7, 32'h3e840b32} /* (3, 5, 8) {real, imag} */,
  {32'hbdefafa2, 32'hbc936170} /* (3, 5, 7) {real, imag} */,
  {32'hbf46d7da, 32'hbc914be0} /* (3, 5, 6) {real, imag} */,
  {32'hbee268c2, 32'hbf5169f8} /* (3, 5, 5) {real, imag} */,
  {32'h3f098b80, 32'h3deafea3} /* (3, 5, 4) {real, imag} */,
  {32'hbf0d44cc, 32'h3ec15a4a} /* (3, 5, 3) {real, imag} */,
  {32'hbebbd2b8, 32'hbece01e2} /* (3, 5, 2) {real, imag} */,
  {32'h402d387a, 32'h40213378} /* (3, 5, 1) {real, imag} */,
  {32'h402529fb, 32'h3e347bcc} /* (3, 5, 0) {real, imag} */,
  {32'hbfbf4fee, 32'hc0359c6e} /* (3, 4, 31) {real, imag} */,
  {32'h3f4fcfdd, 32'h403c406b} /* (3, 4, 30) {real, imag} */,
  {32'hbeff6766, 32'h3f8d0e7c} /* (3, 4, 29) {real, imag} */,
  {32'hbe48bb24, 32'hbf0ce2e6} /* (3, 4, 28) {real, imag} */,
  {32'h3f5cb5ec, 32'hbddb6954} /* (3, 4, 27) {real, imag} */,
  {32'hbea4f123, 32'hbea41377} /* (3, 4, 26) {real, imag} */,
  {32'h3da4a93c, 32'hbee6029e} /* (3, 4, 25) {real, imag} */,
  {32'hbeaf5aba, 32'hbeee86c6} /* (3, 4, 24) {real, imag} */,
  {32'hbf222e48, 32'h3e2b3b33} /* (3, 4, 23) {real, imag} */,
  {32'hbf379946, 32'hbdd549cf} /* (3, 4, 22) {real, imag} */,
  {32'h3f6f032a, 32'hbd9e9408} /* (3, 4, 21) {real, imag} */,
  {32'hbeb82a31, 32'h3ef951d0} /* (3, 4, 20) {real, imag} */,
  {32'hbddb2d97, 32'hbec28c36} /* (3, 4, 19) {real, imag} */,
  {32'h3f096b6d, 32'hbe8d1e38} /* (3, 4, 18) {real, imag} */,
  {32'hbde6faed, 32'hbdebf3dc} /* (3, 4, 17) {real, imag} */,
  {32'h3e1c84eb, 32'hbcdfb802} /* (3, 4, 16) {real, imag} */,
  {32'h3c474160, 32'h3db09dfa} /* (3, 4, 15) {real, imag} */,
  {32'h3e0a91ea, 32'h3e4b3f46} /* (3, 4, 14) {real, imag} */,
  {32'h3dfd4172, 32'h3ef852bc} /* (3, 4, 13) {real, imag} */,
  {32'hbd456ce4, 32'hbd989268} /* (3, 4, 12) {real, imag} */,
  {32'hbde75d09, 32'h3e05063c} /* (3, 4, 11) {real, imag} */,
  {32'hbcd33949, 32'hbe8df6e2} /* (3, 4, 10) {real, imag} */,
  {32'h3ef50e6d, 32'hba458e00} /* (3, 4, 9) {real, imag} */,
  {32'h3e599c9a, 32'h3ed528f3} /* (3, 4, 8) {real, imag} */,
  {32'hbd24c26c, 32'h3ed12b39} /* (3, 4, 7) {real, imag} */,
  {32'h3ec2633a, 32'h3eb13475} /* (3, 4, 6) {real, imag} */,
  {32'h3ddc91a7, 32'h3f2f52e0} /* (3, 4, 5) {real, imag} */,
  {32'hbf6b9e66, 32'hbecda3b2} /* (3, 4, 4) {real, imag} */,
  {32'h3e6e9915, 32'h3f964ecb} /* (3, 4, 3) {real, imag} */,
  {32'h403d88de, 32'h401a7d25} /* (3, 4, 2) {real, imag} */,
  {32'hc0a90769, 32'hbff63bdb} /* (3, 4, 1) {real, imag} */,
  {32'hc014b735, 32'hbf1912a0} /* (3, 4, 0) {real, imag} */,
  {32'h408d693c, 32'hbfc3905a} /* (3, 3, 31) {real, imag} */,
  {32'hbff9392a, 32'h3fbe9b4f} /* (3, 3, 30) {real, imag} */,
  {32'hbe5d3dea, 32'hbf541960} /* (3, 3, 29) {real, imag} */,
  {32'hbec6ea7d, 32'hbe9f9c17} /* (3, 3, 28) {real, imag} */,
  {32'h3f940c60, 32'hbd8b7768} /* (3, 3, 27) {real, imag} */,
  {32'hbdbe99dc, 32'h3e598268} /* (3, 3, 26) {real, imag} */,
  {32'hbe1dcb9f, 32'h3dc04326} /* (3, 3, 25) {real, imag} */,
  {32'hbd8a957c, 32'h3f84ae04} /* (3, 3, 24) {real, imag} */,
  {32'hbeec682b, 32'hbf12afbf} /* (3, 3, 23) {real, imag} */,
  {32'h3e5a1afa, 32'h3e9d646e} /* (3, 3, 22) {real, imag} */,
  {32'h3dbf9ba4, 32'hbf13fba6} /* (3, 3, 21) {real, imag} */,
  {32'hbcbe50f8, 32'h3e7f4ea1} /* (3, 3, 20) {real, imag} */,
  {32'h3e99d8fd, 32'h3cd00d48} /* (3, 3, 19) {real, imag} */,
  {32'hbe015074, 32'hbd352572} /* (3, 3, 18) {real, imag} */,
  {32'hbe6490de, 32'h3d71d8f6} /* (3, 3, 17) {real, imag} */,
  {32'hbe5f8e05, 32'hbe1e2474} /* (3, 3, 16) {real, imag} */,
  {32'hbe7a3db0, 32'hbccef150} /* (3, 3, 15) {real, imag} */,
  {32'h3dc7d21b, 32'h3f352ec5} /* (3, 3, 14) {real, imag} */,
  {32'hbf26515f, 32'hbc8dd438} /* (3, 3, 13) {real, imag} */,
  {32'hbe0284ce, 32'h3e7cf968} /* (3, 3, 12) {real, imag} */,
  {32'hbf3133de, 32'hbf153ff2} /* (3, 3, 11) {real, imag} */,
  {32'hbc5f8084, 32'hbe8457ae} /* (3, 3, 10) {real, imag} */,
  {32'h3f528e27, 32'h3e275646} /* (3, 3, 9) {real, imag} */,
  {32'hbe0270ca, 32'h3ef89a55} /* (3, 3, 8) {real, imag} */,
  {32'h3e7b7fe4, 32'hbf7dbab3} /* (3, 3, 7) {real, imag} */,
  {32'h3d03ae38, 32'hbf7179c1} /* (3, 3, 6) {real, imag} */,
  {32'hbf9c85a2, 32'h3f3b0683} /* (3, 3, 5) {real, imag} */,
  {32'h3fa999f5, 32'h3e0b924e} /* (3, 3, 4) {real, imag} */,
  {32'hbfa39ca2, 32'hbfb61e24} /* (3, 3, 3) {real, imag} */,
  {32'hbed396bb, 32'h408631b4} /* (3, 3, 2) {real, imag} */,
  {32'hc0574aea, 32'hbf4def58} /* (3, 3, 1) {real, imag} */,
  {32'h3f2f1a47, 32'hbf246520} /* (3, 3, 0) {real, imag} */,
  {32'h41a76ee7, 32'h3fc6afd1} /* (3, 2, 31) {real, imag} */,
  {32'hc127120c, 32'h403dd0ef} /* (3, 2, 30) {real, imag} */,
  {32'h3f41b4d3, 32'h3fb49180} /* (3, 2, 29) {real, imag} */,
  {32'h3f7495c3, 32'hc005928a} /* (3, 2, 28) {real, imag} */,
  {32'hbfc6582c, 32'h3fb746a4} /* (3, 2, 27) {real, imag} */,
  {32'hbf09978d, 32'h3d15b70c} /* (3, 2, 26) {real, imag} */,
  {32'h3f4076aa, 32'hbf278db5} /* (3, 2, 25) {real, imag} */,
  {32'hbf8256fc, 32'h3f1dd252} /* (3, 2, 24) {real, imag} */,
  {32'hbf61a859, 32'hbe9e5474} /* (3, 2, 23) {real, imag} */,
  {32'h3f0021a0, 32'hbf1acde5} /* (3, 2, 22) {real, imag} */,
  {32'hbeb0dc3a, 32'h3f6aa619} /* (3, 2, 21) {real, imag} */,
  {32'h3d8c8370, 32'hbea1a997} /* (3, 2, 20) {real, imag} */,
  {32'hbd7a1530, 32'h3ea4b86a} /* (3, 2, 19) {real, imag} */,
  {32'hbde30920, 32'h3f070199} /* (3, 2, 18) {real, imag} */,
  {32'h3d98a610, 32'h3e8d610e} /* (3, 2, 17) {real, imag} */,
  {32'h3d9a680a, 32'hbd151ce0} /* (3, 2, 16) {real, imag} */,
  {32'h3f1017f2, 32'hbebd9e46} /* (3, 2, 15) {real, imag} */,
  {32'h3d99eede, 32'hbed01514} /* (3, 2, 14) {real, imag} */,
  {32'hbdeb1114, 32'hbdc5d86c} /* (3, 2, 13) {real, imag} */,
  {32'h3f2e555e, 32'hbd5d6fe0} /* (3, 2, 12) {real, imag} */,
  {32'hbecd68e3, 32'h3ed40cdc} /* (3, 2, 11) {real, imag} */,
  {32'h3ef132e3, 32'h3b47f600} /* (3, 2, 10) {real, imag} */,
  {32'h3e5b206a, 32'hbec81ca8} /* (3, 2, 9) {real, imag} */,
  {32'hbf6a1dc3, 32'h3c9eed90} /* (3, 2, 8) {real, imag} */,
  {32'h3f8a966e, 32'hbeaa65c0} /* (3, 2, 7) {real, imag} */,
  {32'h3eac336c, 32'h3cb89968} /* (3, 2, 6) {real, imag} */,
  {32'hbfbca142, 32'hbf96aa0b} /* (3, 2, 5) {real, imag} */,
  {32'h4048385c, 32'hbe5b6714} /* (3, 2, 4) {real, imag} */,
  {32'hbf969306, 32'h3e0134c8} /* (3, 2, 3) {real, imag} */,
  {32'hc10d518a, 32'h408a34a9} /* (3, 2, 2) {real, imag} */,
  {32'h4143a854, 32'hbed85dc0} /* (3, 2, 1) {real, imag} */,
  {32'h410ead27, 32'h40203054} /* (3, 2, 0) {real, imag} */,
  {32'hc1910235, 32'h403fa448} /* (3, 1, 31) {real, imag} */,
  {32'h40fb0f50, 32'h3faefbf8} /* (3, 1, 30) {real, imag} */,
  {32'h3fdce602, 32'hbfa27adc} /* (3, 1, 29) {real, imag} */,
  {32'hc0354e47, 32'hbfccad5a} /* (3, 1, 28) {real, imag} */,
  {32'h407bad4c, 32'hbe45e14c} /* (3, 1, 27) {real, imag} */,
  {32'h3f95c0bb, 32'hbec80d04} /* (3, 1, 26) {real, imag} */,
  {32'hbf23b710, 32'h3e869f60} /* (3, 1, 25) {real, imag} */,
  {32'h3f2b861f, 32'hbf44082b} /* (3, 1, 24) {real, imag} */,
  {32'hbe788bdc, 32'hbd6695f0} /* (3, 1, 23) {real, imag} */,
  {32'hbe75bda2, 32'h3df06ba6} /* (3, 1, 22) {real, imag} */,
  {32'h3f73d926, 32'hbf20416a} /* (3, 1, 21) {real, imag} */,
  {32'hbd984bf1, 32'h3e0f84c3} /* (3, 1, 20) {real, imag} */,
  {32'h3d7c7ecc, 32'hbd7e7eaa} /* (3, 1, 19) {real, imag} */,
  {32'hbe76c315, 32'hbee605fe} /* (3, 1, 18) {real, imag} */,
  {32'h3e764116, 32'h3d6efffc} /* (3, 1, 17) {real, imag} */,
  {32'h3e9d0f66, 32'h3c5563e0} /* (3, 1, 16) {real, imag} */,
  {32'h3ea0b3ae, 32'h3e32bac3} /* (3, 1, 15) {real, imag} */,
  {32'hbe1c4f4c, 32'h3e1673d0} /* (3, 1, 14) {real, imag} */,
  {32'hbd6c08e1, 32'hbe954215} /* (3, 1, 13) {real, imag} */,
  {32'hbe8f4d6d, 32'h3daa845d} /* (3, 1, 12) {real, imag} */,
  {32'h3ef17016, 32'h3f27e156} /* (3, 1, 11) {real, imag} */,
  {32'h3e88b990, 32'h3ecf17c0} /* (3, 1, 10) {real, imag} */,
  {32'hbec2dda8, 32'h3df4d03e} /* (3, 1, 9) {real, imag} */,
  {32'h3edd3728, 32'h3faee7e5} /* (3, 1, 8) {real, imag} */,
  {32'hbe5d5c60, 32'hbf0e732e} /* (3, 1, 7) {real, imag} */,
  {32'hbdefcfec, 32'hbe5ba976} /* (3, 1, 6) {real, imag} */,
  {32'h3fff9bfe, 32'h3ff6da63} /* (3, 1, 5) {real, imag} */,
  {32'hbf83f346, 32'hbf747e24} /* (3, 1, 4) {real, imag} */,
  {32'h3f9b1624, 32'hbf3d9cc4} /* (3, 1, 3) {real, imag} */,
  {32'h411a0f1a, 32'h410021d2} /* (3, 1, 2) {real, imag} */,
  {32'hc1c44884, 32'hc18832a4} /* (3, 1, 1) {real, imag} */,
  {32'hc12818e4, 32'h3f85d494} /* (3, 1, 0) {real, imag} */,
  {32'hc1292762, 32'h40f47352} /* (3, 0, 31) {real, imag} */,
  {32'h4019d169, 32'hc024c5ca} /* (3, 0, 30) {real, imag} */,
  {32'h4030fd5c, 32'hbf6a1274} /* (3, 0, 29) {real, imag} */,
  {32'h3e247e74, 32'hc02ad320} /* (3, 0, 28) {real, imag} */,
  {32'h4008722f, 32'hbf8cffe2} /* (3, 0, 27) {real, imag} */,
  {32'h3ecb2ff0, 32'h3ecb0d58} /* (3, 0, 26) {real, imag} */,
  {32'hbe3f1e92, 32'h3edf3371} /* (3, 0, 25) {real, imag} */,
  {32'hbd79635e, 32'hbe19c28b} /* (3, 0, 24) {real, imag} */,
  {32'h3f85765f, 32'h3e400726} /* (3, 0, 23) {real, imag} */,
  {32'hbdb10cea, 32'hbe14ebd2} /* (3, 0, 22) {real, imag} */,
  {32'hbe561730, 32'h3dcd512e} /* (3, 0, 21) {real, imag} */,
  {32'hbe1e658d, 32'h3e0c61b5} /* (3, 0, 20) {real, imag} */,
  {32'hbd620dfb, 32'hbf3a82a8} /* (3, 0, 19) {real, imag} */,
  {32'h3e187b08, 32'h3f15e7b8} /* (3, 0, 18) {real, imag} */,
  {32'h3d72f5fb, 32'hbeb85c4e} /* (3, 0, 17) {real, imag} */,
  {32'h3c3a3178, 32'h00000000} /* (3, 0, 16) {real, imag} */,
  {32'h3d72f5fb, 32'h3eb85c4e} /* (3, 0, 15) {real, imag} */,
  {32'h3e187b08, 32'hbf15e7b8} /* (3, 0, 14) {real, imag} */,
  {32'hbd620dfb, 32'h3f3a82a8} /* (3, 0, 13) {real, imag} */,
  {32'hbe1e658d, 32'hbe0c61b5} /* (3, 0, 12) {real, imag} */,
  {32'hbe561730, 32'hbdcd512e} /* (3, 0, 11) {real, imag} */,
  {32'hbdb10cea, 32'h3e14ebd2} /* (3, 0, 10) {real, imag} */,
  {32'h3f85765f, 32'hbe400726} /* (3, 0, 9) {real, imag} */,
  {32'hbd79635e, 32'h3e19c28b} /* (3, 0, 8) {real, imag} */,
  {32'hbe3f1e92, 32'hbedf3371} /* (3, 0, 7) {real, imag} */,
  {32'h3ecb2ff0, 32'hbecb0d58} /* (3, 0, 6) {real, imag} */,
  {32'h4008722f, 32'h3f8cffe2} /* (3, 0, 5) {real, imag} */,
  {32'h3e247e74, 32'h402ad320} /* (3, 0, 4) {real, imag} */,
  {32'h4030fd5c, 32'h3f6a1274} /* (3, 0, 3) {real, imag} */,
  {32'h4019d169, 32'h4024c5ca} /* (3, 0, 2) {real, imag} */,
  {32'hc1292762, 32'hc0f47352} /* (3, 0, 1) {real, imag} */,
  {32'h408d095b, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc1e907cd, 32'h4193725e} /* (2, 31, 31) {real, imag} */,
  {32'h4123d54f, 32'hc108fcd8} /* (2, 31, 30) {real, imag} */,
  {32'h3fdfb448, 32'h3f2572b7} /* (2, 31, 29) {real, imag} */,
  {32'hbec22e86, 32'h3f7c6dd4} /* (2, 31, 28) {real, imag} */,
  {32'h3fd29f59, 32'hbfdbb22c} /* (2, 31, 27) {real, imag} */,
  {32'hbd84efc0, 32'hbc28db40} /* (2, 31, 26) {real, imag} */,
  {32'hbe58990b, 32'h3f3c837d} /* (2, 31, 25) {real, imag} */,
  {32'h3f334014, 32'hbf684d50} /* (2, 31, 24) {real, imag} */,
  {32'hbdc21ad4, 32'h3dd26afe} /* (2, 31, 23) {real, imag} */,
  {32'h3eda6014, 32'h3e0ffaf9} /* (2, 31, 22) {real, imag} */,
  {32'h3ef4ad1b, 32'hbecc2a32} /* (2, 31, 21) {real, imag} */,
  {32'h3efb333c, 32'h3d6dfbac} /* (2, 31, 20) {real, imag} */,
  {32'hbd9c7f60, 32'h3ef8d327} /* (2, 31, 19) {real, imag} */,
  {32'hbd52ac05, 32'hbe87a08e} /* (2, 31, 18) {real, imag} */,
  {32'h3da1b65a, 32'h3e17137f} /* (2, 31, 17) {real, imag} */,
  {32'hbe923ff8, 32'hbdf6a105} /* (2, 31, 16) {real, imag} */,
  {32'hbdcc8e17, 32'h3ecbe896} /* (2, 31, 15) {real, imag} */,
  {32'hbe5a80d5, 32'h3e1335a7} /* (2, 31, 14) {real, imag} */,
  {32'hbec0ea95, 32'h3ea28405} /* (2, 31, 13) {real, imag} */,
  {32'hbde56644, 32'hbf00bf32} /* (2, 31, 12) {real, imag} */,
  {32'h3f98df18, 32'h3ef2fb38} /* (2, 31, 11) {real, imag} */,
  {32'hbec762d8, 32'hbe9302f3} /* (2, 31, 10) {real, imag} */,
  {32'h3e4952ea, 32'h3e1471c9} /* (2, 31, 9) {real, imag} */,
  {32'h3f65e12a, 32'h3e4913ce} /* (2, 31, 8) {real, imag} */,
  {32'hbd98bdc8, 32'hbe39249a} /* (2, 31, 7) {real, imag} */,
  {32'h3f97b59e, 32'h3efa58a0} /* (2, 31, 6) {real, imag} */,
  {32'h4084ef9c, 32'h3ddfabef} /* (2, 31, 5) {real, imag} */,
  {32'hc03afd8c, 32'h3fb203bd} /* (2, 31, 4) {real, imag} */,
  {32'h3fc721b1, 32'h3fa2b064} /* (2, 31, 3) {real, imag} */,
  {32'h40f6d04c, 32'hbf80fcee} /* (2, 31, 2) {real, imag} */,
  {32'hc19f114e, 32'hc058475e} /* (2, 31, 1) {real, imag} */,
  {32'hc17f6ad2, 32'hbfe409e0} /* (2, 31, 0) {real, imag} */,
  {32'h41344612, 32'h3e3d3590} /* (2, 30, 31) {real, imag} */,
  {32'hc0ff12ef, 32'hc0988f98} /* (2, 30, 30) {real, imag} */,
  {32'hbf8ddc1e, 32'h3f73b55d} /* (2, 30, 29) {real, imag} */,
  {32'h404dc345, 32'hbf535bdc} /* (2, 30, 28) {real, imag} */,
  {32'hbfc5dc90, 32'h3fba7fcf} /* (2, 30, 27) {real, imag} */,
  {32'hbf23c7fa, 32'h3eedf2fa} /* (2, 30, 26) {real, imag} */,
  {32'hbb4a1c60, 32'hbe319e9c} /* (2, 30, 25) {real, imag} */,
  {32'hbf6abcf3, 32'hbec75f89} /* (2, 30, 24) {real, imag} */,
  {32'h3d8c895c, 32'hbe3a4594} /* (2, 30, 23) {real, imag} */,
  {32'h3f62c600, 32'hbf551546} /* (2, 30, 22) {real, imag} */,
  {32'hbcf416b0, 32'h3e9a876e} /* (2, 30, 21) {real, imag} */,
  {32'h3e6155bc, 32'hbf0125af} /* (2, 30, 20) {real, imag} */,
  {32'h3e5f7c14, 32'h3c37d33c} /* (2, 30, 19) {real, imag} */,
  {32'hbce1e188, 32'h3eee348c} /* (2, 30, 18) {real, imag} */,
  {32'hbdde694b, 32'h3ea9fd95} /* (2, 30, 17) {real, imag} */,
  {32'hbd9b6993, 32'h3ebe64ba} /* (2, 30, 16) {real, imag} */,
  {32'h3df66859, 32'h3e999c0a} /* (2, 30, 15) {real, imag} */,
  {32'hbe9f2aeb, 32'hbd087d60} /* (2, 30, 14) {real, imag} */,
  {32'hbe56a184, 32'hbdbb0f18} /* (2, 30, 13) {real, imag} */,
  {32'h3e7e08b0, 32'hbdee65f0} /* (2, 30, 12) {real, imag} */,
  {32'hbe46ffd5, 32'hbf455133} /* (2, 30, 11) {real, imag} */,
  {32'hbe89b59e, 32'h3f23d72c} /* (2, 30, 10) {real, imag} */,
  {32'hbea2e60a, 32'h3e801244} /* (2, 30, 9) {real, imag} */,
  {32'hbfa6c5cf, 32'hbf7a9ce7} /* (2, 30, 8) {real, imag} */,
  {32'h3e3a5829, 32'h3ea17e15} /* (2, 30, 7) {real, imag} */,
  {32'h3e0bec05, 32'h3ebcc014} /* (2, 30, 6) {real, imag} */,
  {32'hbf86e118, 32'hbfdcccc6} /* (2, 30, 5) {real, imag} */,
  {32'h3fceb7cb, 32'h3fbcfc89} /* (2, 30, 4) {real, imag} */,
  {32'h3fcee380, 32'hbf53104c} /* (2, 30, 3) {real, imag} */,
  {32'hc13249c6, 32'hc01af864} /* (2, 30, 2) {real, imag} */,
  {32'h41b4eca6, 32'hc00fcaa9} /* (2, 30, 1) {real, imag} */,
  {32'h4122e7b4, 32'hc05a7243} /* (2, 30, 0) {real, imag} */,
  {32'hc0382e10, 32'h3f87d672} /* (2, 29, 31) {real, imag} */,
  {32'hbf0db9a5, 32'hc0961d4e} /* (2, 29, 30) {real, imag} */,
  {32'hbfcc7612, 32'h3f8b7d8f} /* (2, 29, 29) {real, imag} */,
  {32'h3f642d9d, 32'hbec7f2b6} /* (2, 29, 28) {real, imag} */,
  {32'hbf5bc29f, 32'hbf952930} /* (2, 29, 27) {real, imag} */,
  {32'hbf38addb, 32'hbdd97af5} /* (2, 29, 26) {real, imag} */,
  {32'h3f035836, 32'h3ef16260} /* (2, 29, 25) {real, imag} */,
  {32'hbda3ce2b, 32'hbefaed6a} /* (2, 29, 24) {real, imag} */,
  {32'h3d84f7df, 32'h3b559fc0} /* (2, 29, 23) {real, imag} */,
  {32'h3f1c9116, 32'hbec80c61} /* (2, 29, 22) {real, imag} */,
  {32'hbdb4dfe4, 32'h3edf0747} /* (2, 29, 21) {real, imag} */,
  {32'h3f10bf80, 32'h3e2be3f5} /* (2, 29, 20) {real, imag} */,
  {32'h3a919280, 32'hbe64f9c9} /* (2, 29, 19) {real, imag} */,
  {32'h3e7bec9c, 32'hbf223d2e} /* (2, 29, 18) {real, imag} */,
  {32'h3e25ce7a, 32'h3ecbbb35} /* (2, 29, 17) {real, imag} */,
  {32'hbe2ea740, 32'h3e4d155c} /* (2, 29, 16) {real, imag} */,
  {32'h3ead34a8, 32'h3e8ebe38} /* (2, 29, 15) {real, imag} */,
  {32'h3dc5b7aa, 32'h3ce7d948} /* (2, 29, 14) {real, imag} */,
  {32'hbd728ede, 32'hbe60d55c} /* (2, 29, 13) {real, imag} */,
  {32'hbe6a4bf8, 32'hbf11a97e} /* (2, 29, 12) {real, imag} */,
  {32'hbd04c948, 32'h3e5d0195} /* (2, 29, 11) {real, imag} */,
  {32'hbc9c84b2, 32'hbe3cbd52} /* (2, 29, 10) {real, imag} */,
  {32'hbeb04b02, 32'h3f87833b} /* (2, 29, 9) {real, imag} */,
  {32'hbe716765, 32'hbf3aff6c} /* (2, 29, 8) {real, imag} */,
  {32'hbe901cc3, 32'hbe6f7cab} /* (2, 29, 7) {real, imag} */,
  {32'h3e43fa4c, 32'hbedda79e} /* (2, 29, 6) {real, imag} */,
  {32'h3dbd9806, 32'hbe6c0c68} /* (2, 29, 5) {real, imag} */,
  {32'hbdd3c17c, 32'h3eaf335c} /* (2, 29, 4) {real, imag} */,
  {32'hbfa7278c, 32'h3f5b0308} /* (2, 29, 3) {real, imag} */,
  {32'hc0173cba, 32'hc00ef77f} /* (2, 29, 2) {real, imag} */,
  {32'h409f3a08, 32'h40344ce4} /* (2, 29, 1) {real, imag} */,
  {32'h3f8173f0, 32'h3f7a2460} /* (2, 29, 0) {real, imag} */,
  {32'hc0b43598, 32'h3fcadba7} /* (2, 28, 31) {real, imag} */,
  {32'h404fc2b9, 32'hc064f8c0} /* (2, 28, 30) {real, imag} */,
  {32'h3cb979d8, 32'hbf0945fd} /* (2, 28, 29) {real, imag} */,
  {32'hbd776008, 32'h3df663f8} /* (2, 28, 28) {real, imag} */,
  {32'hbe7d19a4, 32'hbdb4b3c8} /* (2, 28, 27) {real, imag} */,
  {32'h3e8d8a5e, 32'hbe99e61c} /* (2, 28, 26) {real, imag} */,
  {32'hbf1b42ef, 32'hbe2b6100} /* (2, 28, 25) {real, imag} */,
  {32'hbe6594d2, 32'hbf1eab97} /* (2, 28, 24) {real, imag} */,
  {32'h3e8ee724, 32'h3dfdff68} /* (2, 28, 23) {real, imag} */,
  {32'hbdf81cf6, 32'h3cd35630} /* (2, 28, 22) {real, imag} */,
  {32'hbe235982, 32'hbe5e1908} /* (2, 28, 21) {real, imag} */,
  {32'h3e66bf48, 32'hbe077e5e} /* (2, 28, 20) {real, imag} */,
  {32'h3eea7e04, 32'hbea0ecc4} /* (2, 28, 19) {real, imag} */,
  {32'h3ec32590, 32'hbce3aff8} /* (2, 28, 18) {real, imag} */,
  {32'h3e1db033, 32'h3dddb040} /* (2, 28, 17) {real, imag} */,
  {32'h3e35f934, 32'hbe0b0111} /* (2, 28, 16) {real, imag} */,
  {32'hbdb70de8, 32'h3e6665e8} /* (2, 28, 15) {real, imag} */,
  {32'hbec61abe, 32'h3ea18f56} /* (2, 28, 14) {real, imag} */,
  {32'hbf07d80d, 32'h3bfef6f0} /* (2, 28, 13) {real, imag} */,
  {32'h3ddd6d09, 32'h3eaa590e} /* (2, 28, 12) {real, imag} */,
  {32'h3f4e5102, 32'h3e6da2c0} /* (2, 28, 11) {real, imag} */,
  {32'hbe742a00, 32'hbeb98fe1} /* (2, 28, 10) {real, imag} */,
  {32'hbeacb2fe, 32'h3e923672} /* (2, 28, 9) {real, imag} */,
  {32'h3de39b4b, 32'h3f03ca5a} /* (2, 28, 8) {real, imag} */,
  {32'hbe8b6d49, 32'h3f1ae8d8} /* (2, 28, 7) {real, imag} */,
  {32'h3ec98ca3, 32'h3f23b74d} /* (2, 28, 6) {real, imag} */,
  {32'h3f621601, 32'hbeea027e} /* (2, 28, 5) {real, imag} */,
  {32'hbf7ad8bc, 32'h3f5225da} /* (2, 28, 4) {real, imag} */,
  {32'hbee2ad07, 32'hbe440cc0} /* (2, 28, 3) {real, imag} */,
  {32'h3f095e18, 32'hc02dbd78} /* (2, 28, 2) {real, imag} */,
  {32'hc0041c49, 32'h400e6902} /* (2, 28, 1) {real, imag} */,
  {32'hc00863b4, 32'h3f268f73} /* (2, 28, 0) {real, imag} */,
  {32'h4011edd5, 32'hc04a7164} /* (2, 27, 31) {real, imag} */,
  {32'h3d236350, 32'h3ef6ef05} /* (2, 27, 30) {real, imag} */,
  {32'hbdb30576, 32'h3e8a9a44} /* (2, 27, 29) {real, imag} */,
  {32'hbe4cd964, 32'h3e51a49e} /* (2, 27, 28) {real, imag} */,
  {32'hbf1e7668, 32'h3f32d0ee} /* (2, 27, 27) {real, imag} */,
  {32'h3dabcdac, 32'h3e40f16b} /* (2, 27, 26) {real, imag} */,
  {32'hbf651ffa, 32'hbe7d9fb2} /* (2, 27, 25) {real, imag} */,
  {32'hbd162258, 32'h3e96aa06} /* (2, 27, 24) {real, imag} */,
  {32'hbe82b1ad, 32'hbe9ed95f} /* (2, 27, 23) {real, imag} */,
  {32'h3e4af08c, 32'h3d580a00} /* (2, 27, 22) {real, imag} */,
  {32'hbdd27d98, 32'hbe18d8da} /* (2, 27, 21) {real, imag} */,
  {32'hbdc72d94, 32'h3dcae2e4} /* (2, 27, 20) {real, imag} */,
  {32'h3e8012bd, 32'hbeb48675} /* (2, 27, 19) {real, imag} */,
  {32'hbcdf6284, 32'h3eb53fc7} /* (2, 27, 18) {real, imag} */,
  {32'hbe886afb, 32'hbe47f49f} /* (2, 27, 17) {real, imag} */,
  {32'h3e91e5e0, 32'h3e56248c} /* (2, 27, 16) {real, imag} */,
  {32'hbdd1213a, 32'hbe011b00} /* (2, 27, 15) {real, imag} */,
  {32'hbf0e74c7, 32'hbde30a50} /* (2, 27, 14) {real, imag} */,
  {32'h3dae8e9a, 32'hbc4b9d50} /* (2, 27, 13) {real, imag} */,
  {32'hbe7c73f5, 32'h3d73d980} /* (2, 27, 12) {real, imag} */,
  {32'hbe74f15c, 32'hbe724d09} /* (2, 27, 11) {real, imag} */,
  {32'hbe47007e, 32'h3df92480} /* (2, 27, 10) {real, imag} */,
  {32'hbe78e73d, 32'hbec5bba7} /* (2, 27, 9) {real, imag} */,
  {32'h3d44bdd4, 32'hbf524eee} /* (2, 27, 8) {real, imag} */,
  {32'hbe2a7ce8, 32'hbd950796} /* (2, 27, 7) {real, imag} */,
  {32'h3eaddb16, 32'h3ef89de1} /* (2, 27, 6) {real, imag} */,
  {32'hbf7852a9, 32'hbe072b6d} /* (2, 27, 5) {real, imag} */,
  {32'h3e935a02, 32'h3eb2de17} /* (2, 27, 4) {real, imag} */,
  {32'hbe1d0e2e, 32'hbec35bb5} /* (2, 27, 3) {real, imag} */,
  {32'hbfcd1080, 32'h3f3cd08a} /* (2, 27, 2) {real, imag} */,
  {32'h404374f4, 32'hbe62deb0} /* (2, 27, 1) {real, imag} */,
  {32'h4031a711, 32'hbf3409b8} /* (2, 27, 0) {real, imag} */,
  {32'h3e5e2112, 32'h3eba4cd4} /* (2, 26, 31) {real, imag} */,
  {32'hbe74f1c0, 32'h3f3ae389} /* (2, 26, 30) {real, imag} */,
  {32'hb7c04000, 32'h3d28bd04} /* (2, 26, 29) {real, imag} */,
  {32'h3e26ed69, 32'h3e08ef7d} /* (2, 26, 28) {real, imag} */,
  {32'h3ddca074, 32'h3c5403c0} /* (2, 26, 27) {real, imag} */,
  {32'hbe8756ac, 32'hbe193721} /* (2, 26, 26) {real, imag} */,
  {32'hbe1e0792, 32'hbf042dd0} /* (2, 26, 25) {real, imag} */,
  {32'hbe8830ee, 32'h3e392f8c} /* (2, 26, 24) {real, imag} */,
  {32'hbb84da00, 32'hbf2a2bf2} /* (2, 26, 23) {real, imag} */,
  {32'h3f1efe4b, 32'h3dadf6e0} /* (2, 26, 22) {real, imag} */,
  {32'h3ec9d4e2, 32'h3e1715d6} /* (2, 26, 21) {real, imag} */,
  {32'hbf067ea1, 32'h3ed555f3} /* (2, 26, 20) {real, imag} */,
  {32'hbe874c1c, 32'hbe7d7acb} /* (2, 26, 19) {real, imag} */,
  {32'hbd78361a, 32'h3ebd399a} /* (2, 26, 18) {real, imag} */,
  {32'h3d55a3c0, 32'h3dc0acfd} /* (2, 26, 17) {real, imag} */,
  {32'h3c2766e0, 32'h3e9d811d} /* (2, 26, 16) {real, imag} */,
  {32'hbe6dd045, 32'hbdca342e} /* (2, 26, 15) {real, imag} */,
  {32'hbdfb883a, 32'h3e9c2f56} /* (2, 26, 14) {real, imag} */,
  {32'h3e75d092, 32'hb955fc00} /* (2, 26, 13) {real, imag} */,
  {32'h3e9db68c, 32'hbeab7e73} /* (2, 26, 12) {real, imag} */,
  {32'hbd3a5e68, 32'hbe20e058} /* (2, 26, 11) {real, imag} */,
  {32'h3eec288f, 32'h3eb4ecea} /* (2, 26, 10) {real, imag} */,
  {32'hbeca77ae, 32'hbe06a392} /* (2, 26, 9) {real, imag} */,
  {32'hbe383389, 32'hbf1d6487} /* (2, 26, 8) {real, imag} */,
  {32'hbe9718a6, 32'h3dcfb7dc} /* (2, 26, 7) {real, imag} */,
  {32'h3e23e206, 32'h3e98681d} /* (2, 26, 6) {real, imag} */,
  {32'h3d4f3b7e, 32'h3f648fdc} /* (2, 26, 5) {real, imag} */,
  {32'hbf44d0d5, 32'h3f40d341} /* (2, 26, 4) {real, imag} */,
  {32'h3eaa4c3a, 32'hbe92bf4c} /* (2, 26, 3) {real, imag} */,
  {32'hbd146e00, 32'h3e7da365} /* (2, 26, 2) {real, imag} */,
  {32'hbea15b1a, 32'hbf0164d5} /* (2, 26, 1) {real, imag} */,
  {32'h3f07d9f9, 32'hbe9d8f51} /* (2, 26, 0) {real, imag} */,
  {32'hbf025b20, 32'h3eb25113} /* (2, 25, 31) {real, imag} */,
  {32'hbec20da0, 32'hbee273dc} /* (2, 25, 30) {real, imag} */,
  {32'h3ed40ffa, 32'hbddf7ff5} /* (2, 25, 29) {real, imag} */,
  {32'hbe6aa11a, 32'h3ee703ce} /* (2, 25, 28) {real, imag} */,
  {32'hbc38ad50, 32'hbeed54a2} /* (2, 25, 27) {real, imag} */,
  {32'hbe4600fe, 32'h3e2677f6} /* (2, 25, 26) {real, imag} */,
  {32'h3e2cf734, 32'hbdd9a068} /* (2, 25, 25) {real, imag} */,
  {32'hbe12352e, 32'h3ea3e63d} /* (2, 25, 24) {real, imag} */,
  {32'h3eb6064f, 32'hbeef7157} /* (2, 25, 23) {real, imag} */,
  {32'h3ec4f5cb, 32'hbf567524} /* (2, 25, 22) {real, imag} */,
  {32'hbed772f4, 32'h3e90dfd7} /* (2, 25, 21) {real, imag} */,
  {32'h3d5d95f0, 32'h3dabb37a} /* (2, 25, 20) {real, imag} */,
  {32'h3de53529, 32'hbe85883c} /* (2, 25, 19) {real, imag} */,
  {32'hbee6df53, 32'h3ed91c12} /* (2, 25, 18) {real, imag} */,
  {32'h3ec19d14, 32'h3d535672} /* (2, 25, 17) {real, imag} */,
  {32'hbe37e982, 32'hbe0d246c} /* (2, 25, 16) {real, imag} */,
  {32'h3e706de8, 32'h3e69b89e} /* (2, 25, 15) {real, imag} */,
  {32'hbeb51c5b, 32'hbdae3b68} /* (2, 25, 14) {real, imag} */,
  {32'h3ed15753, 32'h3e34edfa} /* (2, 25, 13) {real, imag} */,
  {32'h3cd7bca0, 32'h3dc2dc70} /* (2, 25, 12) {real, imag} */,
  {32'h3e5f7bbe, 32'hbe337c92} /* (2, 25, 11) {real, imag} */,
  {32'hbefd8217, 32'hbebaff4a} /* (2, 25, 10) {real, imag} */,
  {32'hbf3c1c48, 32'hbe62cba6} /* (2, 25, 9) {real, imag} */,
  {32'h3d9ac684, 32'hbd44d5a2} /* (2, 25, 8) {real, imag} */,
  {32'hbee43679, 32'hbf307d50} /* (2, 25, 7) {real, imag} */,
  {32'hbd3aaf78, 32'hbe8a8f43} /* (2, 25, 6) {real, imag} */,
  {32'h3d0119c0, 32'hbed95507} /* (2, 25, 5) {real, imag} */,
  {32'hbf01c744, 32'hbdc42776} /* (2, 25, 4) {real, imag} */,
  {32'hbf2cc2b0, 32'h3ec5907c} /* (2, 25, 3) {real, imag} */,
  {32'hbd269134, 32'h3e6a0951} /* (2, 25, 2) {real, imag} */,
  {32'hbe426dd5, 32'hbdc963f4} /* (2, 25, 1) {real, imag} */,
  {32'h3d16af50, 32'h3ed53c41} /* (2, 25, 0) {real, imag} */,
  {32'h3ee902b0, 32'hbf750973} /* (2, 24, 31) {real, imag} */,
  {32'h3e2734a7, 32'h3f454375} /* (2, 24, 30) {real, imag} */,
  {32'hbdcdde4a, 32'h3cd2aa68} /* (2, 24, 29) {real, imag} */,
  {32'h3d8c1e7c, 32'hbd8461c4} /* (2, 24, 28) {real, imag} */,
  {32'h3d8b8650, 32'h3ddba5de} /* (2, 24, 27) {real, imag} */,
  {32'hbebaf802, 32'h3f70b3d3} /* (2, 24, 26) {real, imag} */,
  {32'hbf29fc84, 32'h3ed41de4} /* (2, 24, 25) {real, imag} */,
  {32'hbde98978, 32'h3b918130} /* (2, 24, 24) {real, imag} */,
  {32'hbee676e3, 32'hbf407b0d} /* (2, 24, 23) {real, imag} */,
  {32'hbc47f550, 32'hbeaa5696} /* (2, 24, 22) {real, imag} */,
  {32'hbe927c2a, 32'h3f4461f6} /* (2, 24, 21) {real, imag} */,
  {32'h3f12fbcb, 32'h3dbda9a6} /* (2, 24, 20) {real, imag} */,
  {32'hbe24a334, 32'h3eb60167} /* (2, 24, 19) {real, imag} */,
  {32'hbd5336d8, 32'h3e9dd96e} /* (2, 24, 18) {real, imag} */,
  {32'h3e11d26a, 32'hbedb532d} /* (2, 24, 17) {real, imag} */,
  {32'h3d949860, 32'hbf0a1288} /* (2, 24, 16) {real, imag} */,
  {32'h3e468b38, 32'h3e497ef6} /* (2, 24, 15) {real, imag} */,
  {32'h3b63d300, 32'h3e27d313} /* (2, 24, 14) {real, imag} */,
  {32'hbd99d4fa, 32'hbf1023ba} /* (2, 24, 13) {real, imag} */,
  {32'h3eb3342d, 32'h3e68bfe0} /* (2, 24, 12) {real, imag} */,
  {32'h3e02e90b, 32'h3ed33d32} /* (2, 24, 11) {real, imag} */,
  {32'hbd8cda56, 32'h3f6a78f4} /* (2, 24, 10) {real, imag} */,
  {32'h3f3f32c0, 32'hbe7bc8dc} /* (2, 24, 9) {real, imag} */,
  {32'h3e101ce9, 32'hbf2225b7} /* (2, 24, 8) {real, imag} */,
  {32'h3f0faff6, 32'hbf4dd8e2} /* (2, 24, 7) {real, imag} */,
  {32'h3ebd1d6f, 32'hbeef7384} /* (2, 24, 6) {real, imag} */,
  {32'hbd06ab10, 32'h3e1bc73a} /* (2, 24, 5) {real, imag} */,
  {32'h3d3b2d59, 32'hbf49c9f2} /* (2, 24, 4) {real, imag} */,
  {32'hbf1fb35e, 32'h3f0e88a5} /* (2, 24, 3) {real, imag} */,
  {32'hbf8cfa02, 32'hbf6694d0} /* (2, 24, 2) {real, imag} */,
  {32'h3fbfe59d, 32'hbf1a4594} /* (2, 24, 1) {real, imag} */,
  {32'h3e7aa4c2, 32'hbd8992f0} /* (2, 24, 0) {real, imag} */,
  {32'hbf1094c7, 32'h3f5e04b6} /* (2, 23, 31) {real, imag} */,
  {32'h3e12d7fa, 32'h3ec7a555} /* (2, 23, 30) {real, imag} */,
  {32'hbf3ba9c5, 32'hbefc9595} /* (2, 23, 29) {real, imag} */,
  {32'hbea039f0, 32'h3ed57300} /* (2, 23, 28) {real, imag} */,
  {32'hbea2f81e, 32'h3f2e8e61} /* (2, 23, 27) {real, imag} */,
  {32'hbd9f40ed, 32'hbf37eaa1} /* (2, 23, 26) {real, imag} */,
  {32'hbd2aa3ec, 32'h3e32d79c} /* (2, 23, 25) {real, imag} */,
  {32'hbecd9aeb, 32'h3d03aaf6} /* (2, 23, 24) {real, imag} */,
  {32'h3eb26b84, 32'hbe24bb01} /* (2, 23, 23) {real, imag} */,
  {32'hbe987cda, 32'h3cd01440} /* (2, 23, 22) {real, imag} */,
  {32'hbe2a84de, 32'hbf060715} /* (2, 23, 21) {real, imag} */,
  {32'hbf2bb034, 32'hbe8a4675} /* (2, 23, 20) {real, imag} */,
  {32'h3eabaef6, 32'h3db07e73} /* (2, 23, 19) {real, imag} */,
  {32'hbed47af4, 32'hbea99f77} /* (2, 23, 18) {real, imag} */,
  {32'hbed5590c, 32'hbebe7896} /* (2, 23, 17) {real, imag} */,
  {32'h3e23887c, 32'hbe94810c} /* (2, 23, 16) {real, imag} */,
  {32'hbe8a31cd, 32'h3e5ac8f3} /* (2, 23, 15) {real, imag} */,
  {32'h3f5158db, 32'h3d82c7c2} /* (2, 23, 14) {real, imag} */,
  {32'hbe981f7c, 32'hbdf661ab} /* (2, 23, 13) {real, imag} */,
  {32'hbf0f57a3, 32'h3e2e70ea} /* (2, 23, 12) {real, imag} */,
  {32'hbe5e5bd8, 32'hbf09042c} /* (2, 23, 11) {real, imag} */,
  {32'h3d3e1a2a, 32'hbcfb5d38} /* (2, 23, 10) {real, imag} */,
  {32'h3d8433e4, 32'h3d8d001e} /* (2, 23, 9) {real, imag} */,
  {32'hbec3e457, 32'hbdc5fdf8} /* (2, 23, 8) {real, imag} */,
  {32'hbddafe68, 32'h3d438a10} /* (2, 23, 7) {real, imag} */,
  {32'h3ea0bcd6, 32'h3d85d455} /* (2, 23, 6) {real, imag} */,
  {32'h3f1f648f, 32'hbe9d3858} /* (2, 23, 5) {real, imag} */,
  {32'h3e2edf54, 32'hbdbee195} /* (2, 23, 4) {real, imag} */,
  {32'hbc887320, 32'h3e7e949e} /* (2, 23, 3) {real, imag} */,
  {32'h3ede5689, 32'hbf55a3cb} /* (2, 23, 2) {real, imag} */,
  {32'h3ee18f6c, 32'hbe236b1b} /* (2, 23, 1) {real, imag} */,
  {32'hbedba0ba, 32'h3f0a62da} /* (2, 23, 0) {real, imag} */,
  {32'hbf235a44, 32'h3ebe38d8} /* (2, 22, 31) {real, imag} */,
  {32'hbeea6a0a, 32'hbf18ed13} /* (2, 22, 30) {real, imag} */,
  {32'h3f51fe31, 32'hbd9f0d0e} /* (2, 22, 29) {real, imag} */,
  {32'h3c7972a8, 32'hbea0fe8f} /* (2, 22, 28) {real, imag} */,
  {32'h3b9514e0, 32'hbed1916e} /* (2, 22, 27) {real, imag} */,
  {32'h3ef4b908, 32'h3e43f601} /* (2, 22, 26) {real, imag} */,
  {32'h3ea4ffbc, 32'hbd953900} /* (2, 22, 25) {real, imag} */,
  {32'hbeda52f2, 32'hbe2761d4} /* (2, 22, 24) {real, imag} */,
  {32'h3e7d4cbf, 32'hbf0818b2} /* (2, 22, 23) {real, imag} */,
  {32'h3f0e1da1, 32'hbde0f4ee} /* (2, 22, 22) {real, imag} */,
  {32'hbe6962f4, 32'h3f16297a} /* (2, 22, 21) {real, imag} */,
  {32'hbed48b1e, 32'h3dae6715} /* (2, 22, 20) {real, imag} */,
  {32'h3e00f4e8, 32'h3f094c5c} /* (2, 22, 19) {real, imag} */,
  {32'h3ddb1868, 32'h3d640ea8} /* (2, 22, 18) {real, imag} */,
  {32'h3c3d2228, 32'h3e5d7372} /* (2, 22, 17) {real, imag} */,
  {32'h3e95e3f7, 32'hbe3b5cc8} /* (2, 22, 16) {real, imag} */,
  {32'hbec3f2f8, 32'h3c4ecd68} /* (2, 22, 15) {real, imag} */,
  {32'h3df2225e, 32'hbebd9596} /* (2, 22, 14) {real, imag} */,
  {32'h3eae2f0a, 32'h3f27b408} /* (2, 22, 13) {real, imag} */,
  {32'hbdd4028c, 32'hbdf47258} /* (2, 22, 12) {real, imag} */,
  {32'hbdad610c, 32'h3f25b692} /* (2, 22, 11) {real, imag} */,
  {32'hbeeca7f2, 32'h3c7cc3e0} /* (2, 22, 10) {real, imag} */,
  {32'hbe36b027, 32'h3e9d074b} /* (2, 22, 9) {real, imag} */,
  {32'hbee505a2, 32'h3e37af91} /* (2, 22, 8) {real, imag} */,
  {32'hbe2ab2c3, 32'h3e0dad3a} /* (2, 22, 7) {real, imag} */,
  {32'h3e6af2d5, 32'h3e3bca7f} /* (2, 22, 6) {real, imag} */,
  {32'h3e0272f6, 32'h3d2c3246} /* (2, 22, 5) {real, imag} */,
  {32'hbf21e576, 32'h3dab89c0} /* (2, 22, 4) {real, imag} */,
  {32'hbf167067, 32'hbe6d43c3} /* (2, 22, 3) {real, imag} */,
  {32'h3eb4688d, 32'hbf452bea} /* (2, 22, 2) {real, imag} */,
  {32'h3d640ef4, 32'h3e140576} /* (2, 22, 1) {real, imag} */,
  {32'h3efee158, 32'h3ea28b36} /* (2, 22, 0) {real, imag} */,
  {32'h3e950630, 32'hbf242e12} /* (2, 21, 31) {real, imag} */,
  {32'hbcc124f0, 32'h3f0fba86} /* (2, 21, 30) {real, imag} */,
  {32'h3d9c9bb6, 32'hbed340b8} /* (2, 21, 29) {real, imag} */,
  {32'h3e7e8260, 32'h3e951a90} /* (2, 21, 28) {real, imag} */,
  {32'h3ea38fa2, 32'hbd3ccc18} /* (2, 21, 27) {real, imag} */,
  {32'hbc36be80, 32'h3c8b53d0} /* (2, 21, 26) {real, imag} */,
  {32'hbe39bb5b, 32'h3cdd1108} /* (2, 21, 25) {real, imag} */,
  {32'h3efa817c, 32'h3f00c014} /* (2, 21, 24) {real, imag} */,
  {32'h3eaa1890, 32'h3e56139b} /* (2, 21, 23) {real, imag} */,
  {32'h3d70c590, 32'h3df58f2a} /* (2, 21, 22) {real, imag} */,
  {32'h3e43509c, 32'h3ea2aa90} /* (2, 21, 21) {real, imag} */,
  {32'h3d9f56b1, 32'h3d3609f4} /* (2, 21, 20) {real, imag} */,
  {32'hbe9a8fa0, 32'h3dc2fc27} /* (2, 21, 19) {real, imag} */,
  {32'h3e57970c, 32'hbe5f68fe} /* (2, 21, 18) {real, imag} */,
  {32'hbd6ab7b8, 32'hbdf6ca36} /* (2, 21, 17) {real, imag} */,
  {32'hbd5b6788, 32'hbeb19e82} /* (2, 21, 16) {real, imag} */,
  {32'hbe0f21e6, 32'h3df487d9} /* (2, 21, 15) {real, imag} */,
  {32'h3e993444, 32'h3d4771e8} /* (2, 21, 14) {real, imag} */,
  {32'h3a429e00, 32'hbe5a7cd4} /* (2, 21, 13) {real, imag} */,
  {32'h3e3b2d34, 32'hbcdbb608} /* (2, 21, 12) {real, imag} */,
  {32'hbe2e3806, 32'hbedeedac} /* (2, 21, 11) {real, imag} */,
  {32'h3eed52aa, 32'hbc96f6d4} /* (2, 21, 10) {real, imag} */,
  {32'hbd9560a0, 32'hbea5ad45} /* (2, 21, 9) {real, imag} */,
  {32'h3ea47580, 32'h3de19368} /* (2, 21, 8) {real, imag} */,
  {32'hbe6fdc5e, 32'h3e079e98} /* (2, 21, 7) {real, imag} */,
  {32'h3d7498f4, 32'hbe90fb77} /* (2, 21, 6) {real, imag} */,
  {32'h3e9dc6fe, 32'hbe38c42c} /* (2, 21, 5) {real, imag} */,
  {32'hbe6dcd6c, 32'hbcc849c8} /* (2, 21, 4) {real, imag} */,
  {32'hbdae3c38, 32'h3ea20466} /* (2, 21, 3) {real, imag} */,
  {32'hbf2b3811, 32'hbe019c74} /* (2, 21, 2) {real, imag} */,
  {32'h3f16ef36, 32'hbf922388} /* (2, 21, 1) {real, imag} */,
  {32'h3eb469dc, 32'hbea93396} /* (2, 21, 0) {real, imag} */,
  {32'hbdbc6b0b, 32'h3de0ab28} /* (2, 20, 31) {real, imag} */,
  {32'hbe9f8386, 32'hbd0f6bde} /* (2, 20, 30) {real, imag} */,
  {32'hbd9da997, 32'h3d8f896a} /* (2, 20, 29) {real, imag} */,
  {32'h3d4cda0e, 32'hbc5e1908} /* (2, 20, 28) {real, imag} */,
  {32'hbd5c7068, 32'hbcad4e88} /* (2, 20, 27) {real, imag} */,
  {32'hbdc79020, 32'h3e7131ba} /* (2, 20, 26) {real, imag} */,
  {32'hbf25acc6, 32'hbe68b30e} /* (2, 20, 25) {real, imag} */,
  {32'h3e149283, 32'h3ec53686} /* (2, 20, 24) {real, imag} */,
  {32'h3dd14877, 32'h3e8f5550} /* (2, 20, 23) {real, imag} */,
  {32'h3ef59b44, 32'h3ed7f1b0} /* (2, 20, 22) {real, imag} */,
  {32'hbec41ed2, 32'h3eee752c} /* (2, 20, 21) {real, imag} */,
  {32'hbdf55008, 32'hbd40e9b6} /* (2, 20, 20) {real, imag} */,
  {32'hbebc8b41, 32'hbf399c3b} /* (2, 20, 19) {real, imag} */,
  {32'hbe90827b, 32'h3d6d0518} /* (2, 20, 18) {real, imag} */,
  {32'hbd308ad7, 32'hbf068468} /* (2, 20, 17) {real, imag} */,
  {32'h3d7ec3eb, 32'hbee2345c} /* (2, 20, 16) {real, imag} */,
  {32'hbe981faa, 32'hbefa7d9a} /* (2, 20, 15) {real, imag} */,
  {32'hbe95a57c, 32'hbf1794f4} /* (2, 20, 14) {real, imag} */,
  {32'hbedbbd3a, 32'hbea9b239} /* (2, 20, 13) {real, imag} */,
  {32'h3f0eb4a7, 32'hbe3c2441} /* (2, 20, 12) {real, imag} */,
  {32'h3eb23823, 32'h3e1c4437} /* (2, 20, 11) {real, imag} */,
  {32'h3da6977c, 32'h3e7338b4} /* (2, 20, 10) {real, imag} */,
  {32'h3e6e8af4, 32'h3d1d3ac2} /* (2, 20, 9) {real, imag} */,
  {32'hbde658fb, 32'hbe67bbda} /* (2, 20, 8) {real, imag} */,
  {32'h3ea4e712, 32'h3eb265a9} /* (2, 20, 7) {real, imag} */,
  {32'h3e1bc772, 32'hbeb81e78} /* (2, 20, 6) {real, imag} */,
  {32'h3ecb292f, 32'h3e9180f5} /* (2, 20, 5) {real, imag} */,
  {32'h3e4bb529, 32'hbe1215a5} /* (2, 20, 4) {real, imag} */,
  {32'h3ee40260, 32'h3ecde44a} /* (2, 20, 3) {real, imag} */,
  {32'h3ddc449c, 32'hbbcd1c00} /* (2, 20, 2) {real, imag} */,
  {32'h3ef0e490, 32'h3edbdf4a} /* (2, 20, 1) {real, imag} */,
  {32'h3e716628, 32'h3e94c54f} /* (2, 20, 0) {real, imag} */,
  {32'h3e6f7810, 32'hbebbfd7e} /* (2, 19, 31) {real, imag} */,
  {32'h3d019a4c, 32'hbe428f84} /* (2, 19, 30) {real, imag} */,
  {32'hbd52f394, 32'hbeb8a80e} /* (2, 19, 29) {real, imag} */,
  {32'hbf2a6816, 32'hbec58ec1} /* (2, 19, 28) {real, imag} */,
  {32'h3ee84603, 32'h3e4aa200} /* (2, 19, 27) {real, imag} */,
  {32'hbdc38270, 32'h3eaf16e2} /* (2, 19, 26) {real, imag} */,
  {32'hbe9ff6e7, 32'hbe04d333} /* (2, 19, 25) {real, imag} */,
  {32'hbeee1339, 32'hbebf2640} /* (2, 19, 24) {real, imag} */,
  {32'h3e56e36a, 32'h3f114560} /* (2, 19, 23) {real, imag} */,
  {32'hbee5cde0, 32'hbe2d3300} /* (2, 19, 22) {real, imag} */,
  {32'hbe5edf98, 32'h3f051b42} /* (2, 19, 21) {real, imag} */,
  {32'hbe7b67b8, 32'h3e8393ec} /* (2, 19, 20) {real, imag} */,
  {32'hbd421e2c, 32'h3d53e811} /* (2, 19, 19) {real, imag} */,
  {32'hbea73eb3, 32'hbf25edd2} /* (2, 19, 18) {real, imag} */,
  {32'h3d8bc480, 32'h3d7f4fa8} /* (2, 19, 17) {real, imag} */,
  {32'hbe9b85b5, 32'h3d98817a} /* (2, 19, 16) {real, imag} */,
  {32'hbd0f46cc, 32'hbec9d364} /* (2, 19, 15) {real, imag} */,
  {32'h3ec0b11e, 32'h3e99b99c} /* (2, 19, 14) {real, imag} */,
  {32'hbf1a3f60, 32'hbe8a7fa4} /* (2, 19, 13) {real, imag} */,
  {32'hbd3beefe, 32'h3dff0648} /* (2, 19, 12) {real, imag} */,
  {32'hbd0fe33e, 32'hbdd703f4} /* (2, 19, 11) {real, imag} */,
  {32'hbd7f01e4, 32'h3e8ec673} /* (2, 19, 10) {real, imag} */,
  {32'hbe851097, 32'h3dfe5f90} /* (2, 19, 9) {real, imag} */,
  {32'h3eb198b7, 32'h3b247140} /* (2, 19, 8) {real, imag} */,
  {32'h3e6872aa, 32'hbe9c3797} /* (2, 19, 7) {real, imag} */,
  {32'hbd672312, 32'h3c297e40} /* (2, 19, 6) {real, imag} */,
  {32'hbe250985, 32'h3cbdd89c} /* (2, 19, 5) {real, imag} */,
  {32'hbe2a4ce2, 32'h3d706b86} /* (2, 19, 4) {real, imag} */,
  {32'hbdad0beb, 32'hbe1f769b} /* (2, 19, 3) {real, imag} */,
  {32'h3dfccfd0, 32'h3e8f5806} /* (2, 19, 2) {real, imag} */,
  {32'hbedf89ee, 32'h3ed1069c} /* (2, 19, 1) {real, imag} */,
  {32'hbe981e2c, 32'h3eeda6e7} /* (2, 19, 0) {real, imag} */,
  {32'h3ebb3896, 32'hbe253f58} /* (2, 18, 31) {real, imag} */,
  {32'hbe83baef, 32'hbd8d0212} /* (2, 18, 30) {real, imag} */,
  {32'hbe5e521f, 32'hbd31053c} /* (2, 18, 29) {real, imag} */,
  {32'h3dd679a6, 32'hbd6802a4} /* (2, 18, 28) {real, imag} */,
  {32'hbd7436f4, 32'h3ec5ea9a} /* (2, 18, 27) {real, imag} */,
  {32'h3da2065c, 32'hbe5d0cd6} /* (2, 18, 26) {real, imag} */,
  {32'hbe981398, 32'hbf3688f7} /* (2, 18, 25) {real, imag} */,
  {32'hbec75721, 32'hbe1cf1c8} /* (2, 18, 24) {real, imag} */,
  {32'h3f1832ab, 32'hbf1ad2be} /* (2, 18, 23) {real, imag} */,
  {32'hbec82816, 32'hbdfe589a} /* (2, 18, 22) {real, imag} */,
  {32'h3f033589, 32'h3ed1827f} /* (2, 18, 21) {real, imag} */,
  {32'h3dfba27e, 32'h3eecef91} /* (2, 18, 20) {real, imag} */,
  {32'h3df0356a, 32'h3f2b96d4} /* (2, 18, 19) {real, imag} */,
  {32'hbdd4b400, 32'h3de8e0a8} /* (2, 18, 18) {real, imag} */,
  {32'h3eab93a1, 32'hbdde86b9} /* (2, 18, 17) {real, imag} */,
  {32'hbea1e99a, 32'h3e2a8c38} /* (2, 18, 16) {real, imag} */,
  {32'h3e2d576a, 32'hbe550b62} /* (2, 18, 15) {real, imag} */,
  {32'hbe8f9e87, 32'hbe5ac9da} /* (2, 18, 14) {real, imag} */,
  {32'hbcda2604, 32'hbd40c930} /* (2, 18, 13) {real, imag} */,
  {32'hbe78bda5, 32'h3f21dab2} /* (2, 18, 12) {real, imag} */,
  {32'hbdccdf7a, 32'h3f212ffd} /* (2, 18, 11) {real, imag} */,
  {32'h3e3485ba, 32'hbef8ba26} /* (2, 18, 10) {real, imag} */,
  {32'hbf54a70c, 32'h3d98bfa4} /* (2, 18, 9) {real, imag} */,
  {32'hbe5fdadc, 32'hbdeb5801} /* (2, 18, 8) {real, imag} */,
  {32'hb9886000, 32'hbe9f29b1} /* (2, 18, 7) {real, imag} */,
  {32'h3deaf564, 32'h3e8d6366} /* (2, 18, 6) {real, imag} */,
  {32'hbe27f9c1, 32'hbd4f33ac} /* (2, 18, 5) {real, imag} */,
  {32'h3f010098, 32'hbeb7ddf6} /* (2, 18, 4) {real, imag} */,
  {32'h3e87526f, 32'h3e99e75c} /* (2, 18, 3) {real, imag} */,
  {32'hbdd69866, 32'h3e9bee80} /* (2, 18, 2) {real, imag} */,
  {32'h3d16bee4, 32'hbf36e4a8} /* (2, 18, 1) {real, imag} */,
  {32'hbda335c2, 32'h3dbc2b16} /* (2, 18, 0) {real, imag} */,
  {32'h3e050424, 32'h3ee7f44e} /* (2, 17, 31) {real, imag} */,
  {32'hbe59381c, 32'hbe362eac} /* (2, 17, 30) {real, imag} */,
  {32'h3dff4cd4, 32'hbe1550e2} /* (2, 17, 29) {real, imag} */,
  {32'h3e979a10, 32'hbe42257c} /* (2, 17, 28) {real, imag} */,
  {32'hbe37ea58, 32'h3e1850a3} /* (2, 17, 27) {real, imag} */,
  {32'h3e49ae36, 32'hbe895caf} /* (2, 17, 26) {real, imag} */,
  {32'h3e2a3227, 32'h3dad37dd} /* (2, 17, 25) {real, imag} */,
  {32'hbe75700a, 32'hbdd851be} /* (2, 17, 24) {real, imag} */,
  {32'hbeddcc0b, 32'hbe262cb2} /* (2, 17, 23) {real, imag} */,
  {32'h3ec07082, 32'hbda0d6bb} /* (2, 17, 22) {real, imag} */,
  {32'hbe11caf8, 32'h3effb04e} /* (2, 17, 21) {real, imag} */,
  {32'h3e2dbdbd, 32'hbe0bb1b2} /* (2, 17, 20) {real, imag} */,
  {32'hbe8a0bab, 32'hbe2027f4} /* (2, 17, 19) {real, imag} */,
  {32'hbe73958f, 32'h3d6deb6c} /* (2, 17, 18) {real, imag} */,
  {32'hbe0fb784, 32'h3d8774a4} /* (2, 17, 17) {real, imag} */,
  {32'h3e723a0f, 32'h3e84618b} /* (2, 17, 16) {real, imag} */,
  {32'hbe2eac21, 32'h3d407d54} /* (2, 17, 15) {real, imag} */,
  {32'hbe3c6c8e, 32'hbe13338e} /* (2, 17, 14) {real, imag} */,
  {32'h3c6c7c80, 32'h3f25c8b3} /* (2, 17, 13) {real, imag} */,
  {32'h3dc109e3, 32'hbee8077a} /* (2, 17, 12) {real, imag} */,
  {32'h3ef49654, 32'hbb2dd580} /* (2, 17, 11) {real, imag} */,
  {32'h3ddcafee, 32'hbe4aae3e} /* (2, 17, 10) {real, imag} */,
  {32'h3e85bd25, 32'hbeb39f98} /* (2, 17, 9) {real, imag} */,
  {32'h3f06f1f6, 32'h3ea681b7} /* (2, 17, 8) {real, imag} */,
  {32'hbe32404f, 32'hbefc9060} /* (2, 17, 7) {real, imag} */,
  {32'h3e0485f8, 32'hbd8991a5} /* (2, 17, 6) {real, imag} */,
  {32'h3f017b3a, 32'h3ecab793} /* (2, 17, 5) {real, imag} */,
  {32'hbdc9e498, 32'h3e2b07c4} /* (2, 17, 4) {real, imag} */,
  {32'hbe262469, 32'h3dab9b77} /* (2, 17, 3) {real, imag} */,
  {32'hbe548bf0, 32'hbd1184a0} /* (2, 17, 2) {real, imag} */,
  {32'hbe4a0338, 32'h3e82f1aa} /* (2, 17, 1) {real, imag} */,
  {32'hbe68dfd4, 32'h3c655a88} /* (2, 17, 0) {real, imag} */,
  {32'h3daeef54, 32'h3df3060d} /* (2, 16, 31) {real, imag} */,
  {32'h3e18ae3f, 32'h3e338c2c} /* (2, 16, 30) {real, imag} */,
  {32'hbeb7959d, 32'h3f1dd25c} /* (2, 16, 29) {real, imag} */,
  {32'h3e1d9bd3, 32'h3e871093} /* (2, 16, 28) {real, imag} */,
  {32'h3e1497b6, 32'hbdfd1a38} /* (2, 16, 27) {real, imag} */,
  {32'h3d6885fa, 32'h3e55665a} /* (2, 16, 26) {real, imag} */,
  {32'hbdba188e, 32'hbd51fd80} /* (2, 16, 25) {real, imag} */,
  {32'hbe835dc0, 32'h3ec7dd90} /* (2, 16, 24) {real, imag} */,
  {32'hbe8b892e, 32'hbe7a6985} /* (2, 16, 23) {real, imag} */,
  {32'h3d112fa4, 32'hbe8ec5ce} /* (2, 16, 22) {real, imag} */,
  {32'hbe14e864, 32'h3e6d4942} /* (2, 16, 21) {real, imag} */,
  {32'h3e8123b7, 32'hbcff4288} /* (2, 16, 20) {real, imag} */,
  {32'h3e3df236, 32'hbebd7a9a} /* (2, 16, 19) {real, imag} */,
  {32'h3e60ddd1, 32'hbbb29d00} /* (2, 16, 18) {real, imag} */,
  {32'hbe4b72b6, 32'hbe6cb332} /* (2, 16, 17) {real, imag} */,
  {32'hbcb147a8, 32'h00000000} /* (2, 16, 16) {real, imag} */,
  {32'hbe4b72b6, 32'h3e6cb332} /* (2, 16, 15) {real, imag} */,
  {32'h3e60ddd1, 32'h3bb29d00} /* (2, 16, 14) {real, imag} */,
  {32'h3e3df236, 32'h3ebd7a9a} /* (2, 16, 13) {real, imag} */,
  {32'h3e8123b7, 32'h3cff4288} /* (2, 16, 12) {real, imag} */,
  {32'hbe14e864, 32'hbe6d4942} /* (2, 16, 11) {real, imag} */,
  {32'h3d112fa4, 32'h3e8ec5ce} /* (2, 16, 10) {real, imag} */,
  {32'hbe8b892e, 32'h3e7a6985} /* (2, 16, 9) {real, imag} */,
  {32'hbe835dc0, 32'hbec7dd90} /* (2, 16, 8) {real, imag} */,
  {32'hbdba188e, 32'h3d51fd80} /* (2, 16, 7) {real, imag} */,
  {32'h3d6885fa, 32'hbe55665a} /* (2, 16, 6) {real, imag} */,
  {32'h3e1497b6, 32'h3dfd1a38} /* (2, 16, 5) {real, imag} */,
  {32'h3e1d9bd3, 32'hbe871093} /* (2, 16, 4) {real, imag} */,
  {32'hbeb7959d, 32'hbf1dd25c} /* (2, 16, 3) {real, imag} */,
  {32'h3e18ae3f, 32'hbe338c2c} /* (2, 16, 2) {real, imag} */,
  {32'h3daeef54, 32'hbdf3060d} /* (2, 16, 1) {real, imag} */,
  {32'hbe24dba6, 32'h00000000} /* (2, 16, 0) {real, imag} */,
  {32'hbe4a0338, 32'hbe82f1aa} /* (2, 15, 31) {real, imag} */,
  {32'hbe548bf0, 32'h3d1184a0} /* (2, 15, 30) {real, imag} */,
  {32'hbe262469, 32'hbdab9b77} /* (2, 15, 29) {real, imag} */,
  {32'hbdc9e498, 32'hbe2b07c4} /* (2, 15, 28) {real, imag} */,
  {32'h3f017b3a, 32'hbecab793} /* (2, 15, 27) {real, imag} */,
  {32'h3e0485f8, 32'h3d8991a5} /* (2, 15, 26) {real, imag} */,
  {32'hbe32404f, 32'h3efc9060} /* (2, 15, 25) {real, imag} */,
  {32'h3f06f1f6, 32'hbea681b7} /* (2, 15, 24) {real, imag} */,
  {32'h3e85bd25, 32'h3eb39f98} /* (2, 15, 23) {real, imag} */,
  {32'h3ddcafee, 32'h3e4aae3e} /* (2, 15, 22) {real, imag} */,
  {32'h3ef49654, 32'h3b2dd580} /* (2, 15, 21) {real, imag} */,
  {32'h3dc109e3, 32'h3ee8077a} /* (2, 15, 20) {real, imag} */,
  {32'h3c6c7c80, 32'hbf25c8b3} /* (2, 15, 19) {real, imag} */,
  {32'hbe3c6c8e, 32'h3e13338e} /* (2, 15, 18) {real, imag} */,
  {32'hbe2eac21, 32'hbd407d54} /* (2, 15, 17) {real, imag} */,
  {32'h3e723a0f, 32'hbe84618b} /* (2, 15, 16) {real, imag} */,
  {32'hbe0fb784, 32'hbd8774a4} /* (2, 15, 15) {real, imag} */,
  {32'hbe73958f, 32'hbd6deb6c} /* (2, 15, 14) {real, imag} */,
  {32'hbe8a0bab, 32'h3e2027f4} /* (2, 15, 13) {real, imag} */,
  {32'h3e2dbdbd, 32'h3e0bb1b2} /* (2, 15, 12) {real, imag} */,
  {32'hbe11caf8, 32'hbeffb04e} /* (2, 15, 11) {real, imag} */,
  {32'h3ec07082, 32'h3da0d6bb} /* (2, 15, 10) {real, imag} */,
  {32'hbeddcc0b, 32'h3e262cb2} /* (2, 15, 9) {real, imag} */,
  {32'hbe75700a, 32'h3dd851be} /* (2, 15, 8) {real, imag} */,
  {32'h3e2a3227, 32'hbdad37dd} /* (2, 15, 7) {real, imag} */,
  {32'h3e49ae36, 32'h3e895caf} /* (2, 15, 6) {real, imag} */,
  {32'hbe37ea58, 32'hbe1850a3} /* (2, 15, 5) {real, imag} */,
  {32'h3e979a10, 32'h3e42257c} /* (2, 15, 4) {real, imag} */,
  {32'h3dff4cd4, 32'h3e1550e2} /* (2, 15, 3) {real, imag} */,
  {32'hbe59381c, 32'h3e362eac} /* (2, 15, 2) {real, imag} */,
  {32'h3e050424, 32'hbee7f44e} /* (2, 15, 1) {real, imag} */,
  {32'hbe68dfd4, 32'hbc655a88} /* (2, 15, 0) {real, imag} */,
  {32'h3d16bee4, 32'h3f36e4a8} /* (2, 14, 31) {real, imag} */,
  {32'hbdd69866, 32'hbe9bee80} /* (2, 14, 30) {real, imag} */,
  {32'h3e87526f, 32'hbe99e75c} /* (2, 14, 29) {real, imag} */,
  {32'h3f010098, 32'h3eb7ddf6} /* (2, 14, 28) {real, imag} */,
  {32'hbe27f9c1, 32'h3d4f33ac} /* (2, 14, 27) {real, imag} */,
  {32'h3deaf564, 32'hbe8d6366} /* (2, 14, 26) {real, imag} */,
  {32'hb9886000, 32'h3e9f29b1} /* (2, 14, 25) {real, imag} */,
  {32'hbe5fdadc, 32'h3deb5801} /* (2, 14, 24) {real, imag} */,
  {32'hbf54a70c, 32'hbd98bfa4} /* (2, 14, 23) {real, imag} */,
  {32'h3e3485ba, 32'h3ef8ba26} /* (2, 14, 22) {real, imag} */,
  {32'hbdccdf7a, 32'hbf212ffd} /* (2, 14, 21) {real, imag} */,
  {32'hbe78bda5, 32'hbf21dab2} /* (2, 14, 20) {real, imag} */,
  {32'hbcda2604, 32'h3d40c930} /* (2, 14, 19) {real, imag} */,
  {32'hbe8f9e87, 32'h3e5ac9da} /* (2, 14, 18) {real, imag} */,
  {32'h3e2d576a, 32'h3e550b62} /* (2, 14, 17) {real, imag} */,
  {32'hbea1e99a, 32'hbe2a8c38} /* (2, 14, 16) {real, imag} */,
  {32'h3eab93a1, 32'h3dde86b9} /* (2, 14, 15) {real, imag} */,
  {32'hbdd4b400, 32'hbde8e0a8} /* (2, 14, 14) {real, imag} */,
  {32'h3df0356a, 32'hbf2b96d4} /* (2, 14, 13) {real, imag} */,
  {32'h3dfba27e, 32'hbeecef91} /* (2, 14, 12) {real, imag} */,
  {32'h3f033589, 32'hbed1827f} /* (2, 14, 11) {real, imag} */,
  {32'hbec82816, 32'h3dfe589a} /* (2, 14, 10) {real, imag} */,
  {32'h3f1832ab, 32'h3f1ad2be} /* (2, 14, 9) {real, imag} */,
  {32'hbec75721, 32'h3e1cf1c8} /* (2, 14, 8) {real, imag} */,
  {32'hbe981398, 32'h3f3688f7} /* (2, 14, 7) {real, imag} */,
  {32'h3da2065c, 32'h3e5d0cd6} /* (2, 14, 6) {real, imag} */,
  {32'hbd7436f4, 32'hbec5ea9a} /* (2, 14, 5) {real, imag} */,
  {32'h3dd679a6, 32'h3d6802a4} /* (2, 14, 4) {real, imag} */,
  {32'hbe5e521f, 32'h3d31053c} /* (2, 14, 3) {real, imag} */,
  {32'hbe83baef, 32'h3d8d0212} /* (2, 14, 2) {real, imag} */,
  {32'h3ebb3896, 32'h3e253f58} /* (2, 14, 1) {real, imag} */,
  {32'hbda335c2, 32'hbdbc2b16} /* (2, 14, 0) {real, imag} */,
  {32'hbedf89ee, 32'hbed1069c} /* (2, 13, 31) {real, imag} */,
  {32'h3dfccfd0, 32'hbe8f5806} /* (2, 13, 30) {real, imag} */,
  {32'hbdad0beb, 32'h3e1f769b} /* (2, 13, 29) {real, imag} */,
  {32'hbe2a4ce2, 32'hbd706b86} /* (2, 13, 28) {real, imag} */,
  {32'hbe250985, 32'hbcbdd89c} /* (2, 13, 27) {real, imag} */,
  {32'hbd672312, 32'hbc297e40} /* (2, 13, 26) {real, imag} */,
  {32'h3e6872aa, 32'h3e9c3797} /* (2, 13, 25) {real, imag} */,
  {32'h3eb198b7, 32'hbb247140} /* (2, 13, 24) {real, imag} */,
  {32'hbe851097, 32'hbdfe5f90} /* (2, 13, 23) {real, imag} */,
  {32'hbd7f01e4, 32'hbe8ec673} /* (2, 13, 22) {real, imag} */,
  {32'hbd0fe33e, 32'h3dd703f4} /* (2, 13, 21) {real, imag} */,
  {32'hbd3beefe, 32'hbdff0648} /* (2, 13, 20) {real, imag} */,
  {32'hbf1a3f60, 32'h3e8a7fa4} /* (2, 13, 19) {real, imag} */,
  {32'h3ec0b11e, 32'hbe99b99c} /* (2, 13, 18) {real, imag} */,
  {32'hbd0f46cc, 32'h3ec9d364} /* (2, 13, 17) {real, imag} */,
  {32'hbe9b85b5, 32'hbd98817a} /* (2, 13, 16) {real, imag} */,
  {32'h3d8bc480, 32'hbd7f4fa8} /* (2, 13, 15) {real, imag} */,
  {32'hbea73eb3, 32'h3f25edd2} /* (2, 13, 14) {real, imag} */,
  {32'hbd421e2c, 32'hbd53e811} /* (2, 13, 13) {real, imag} */,
  {32'hbe7b67b8, 32'hbe8393ec} /* (2, 13, 12) {real, imag} */,
  {32'hbe5edf98, 32'hbf051b42} /* (2, 13, 11) {real, imag} */,
  {32'hbee5cde0, 32'h3e2d3300} /* (2, 13, 10) {real, imag} */,
  {32'h3e56e36a, 32'hbf114560} /* (2, 13, 9) {real, imag} */,
  {32'hbeee1339, 32'h3ebf2640} /* (2, 13, 8) {real, imag} */,
  {32'hbe9ff6e7, 32'h3e04d333} /* (2, 13, 7) {real, imag} */,
  {32'hbdc38270, 32'hbeaf16e2} /* (2, 13, 6) {real, imag} */,
  {32'h3ee84603, 32'hbe4aa200} /* (2, 13, 5) {real, imag} */,
  {32'hbf2a6816, 32'h3ec58ec1} /* (2, 13, 4) {real, imag} */,
  {32'hbd52f394, 32'h3eb8a80e} /* (2, 13, 3) {real, imag} */,
  {32'h3d019a4c, 32'h3e428f84} /* (2, 13, 2) {real, imag} */,
  {32'h3e6f7810, 32'h3ebbfd7e} /* (2, 13, 1) {real, imag} */,
  {32'hbe981e2c, 32'hbeeda6e7} /* (2, 13, 0) {real, imag} */,
  {32'h3ef0e490, 32'hbedbdf4a} /* (2, 12, 31) {real, imag} */,
  {32'h3ddc449c, 32'h3bcd1c00} /* (2, 12, 30) {real, imag} */,
  {32'h3ee40260, 32'hbecde44a} /* (2, 12, 29) {real, imag} */,
  {32'h3e4bb529, 32'h3e1215a5} /* (2, 12, 28) {real, imag} */,
  {32'h3ecb292f, 32'hbe9180f5} /* (2, 12, 27) {real, imag} */,
  {32'h3e1bc772, 32'h3eb81e78} /* (2, 12, 26) {real, imag} */,
  {32'h3ea4e712, 32'hbeb265a9} /* (2, 12, 25) {real, imag} */,
  {32'hbde658fb, 32'h3e67bbda} /* (2, 12, 24) {real, imag} */,
  {32'h3e6e8af4, 32'hbd1d3ac2} /* (2, 12, 23) {real, imag} */,
  {32'h3da6977c, 32'hbe7338b4} /* (2, 12, 22) {real, imag} */,
  {32'h3eb23823, 32'hbe1c4437} /* (2, 12, 21) {real, imag} */,
  {32'h3f0eb4a7, 32'h3e3c2441} /* (2, 12, 20) {real, imag} */,
  {32'hbedbbd3a, 32'h3ea9b239} /* (2, 12, 19) {real, imag} */,
  {32'hbe95a57c, 32'h3f1794f4} /* (2, 12, 18) {real, imag} */,
  {32'hbe981faa, 32'h3efa7d9a} /* (2, 12, 17) {real, imag} */,
  {32'h3d7ec3eb, 32'h3ee2345c} /* (2, 12, 16) {real, imag} */,
  {32'hbd308ad7, 32'h3f068468} /* (2, 12, 15) {real, imag} */,
  {32'hbe90827b, 32'hbd6d0518} /* (2, 12, 14) {real, imag} */,
  {32'hbebc8b41, 32'h3f399c3b} /* (2, 12, 13) {real, imag} */,
  {32'hbdf55008, 32'h3d40e9b6} /* (2, 12, 12) {real, imag} */,
  {32'hbec41ed2, 32'hbeee752c} /* (2, 12, 11) {real, imag} */,
  {32'h3ef59b44, 32'hbed7f1b0} /* (2, 12, 10) {real, imag} */,
  {32'h3dd14877, 32'hbe8f5550} /* (2, 12, 9) {real, imag} */,
  {32'h3e149283, 32'hbec53686} /* (2, 12, 8) {real, imag} */,
  {32'hbf25acc6, 32'h3e68b30e} /* (2, 12, 7) {real, imag} */,
  {32'hbdc79020, 32'hbe7131ba} /* (2, 12, 6) {real, imag} */,
  {32'hbd5c7068, 32'h3cad4e88} /* (2, 12, 5) {real, imag} */,
  {32'h3d4cda0e, 32'h3c5e1908} /* (2, 12, 4) {real, imag} */,
  {32'hbd9da997, 32'hbd8f896a} /* (2, 12, 3) {real, imag} */,
  {32'hbe9f8386, 32'h3d0f6bde} /* (2, 12, 2) {real, imag} */,
  {32'hbdbc6b0b, 32'hbde0ab28} /* (2, 12, 1) {real, imag} */,
  {32'h3e716628, 32'hbe94c54f} /* (2, 12, 0) {real, imag} */,
  {32'h3f16ef36, 32'h3f922388} /* (2, 11, 31) {real, imag} */,
  {32'hbf2b3811, 32'h3e019c74} /* (2, 11, 30) {real, imag} */,
  {32'hbdae3c38, 32'hbea20466} /* (2, 11, 29) {real, imag} */,
  {32'hbe6dcd6c, 32'h3cc849c8} /* (2, 11, 28) {real, imag} */,
  {32'h3e9dc6fe, 32'h3e38c42c} /* (2, 11, 27) {real, imag} */,
  {32'h3d7498f4, 32'h3e90fb77} /* (2, 11, 26) {real, imag} */,
  {32'hbe6fdc5e, 32'hbe079e98} /* (2, 11, 25) {real, imag} */,
  {32'h3ea47580, 32'hbde19368} /* (2, 11, 24) {real, imag} */,
  {32'hbd9560a0, 32'h3ea5ad45} /* (2, 11, 23) {real, imag} */,
  {32'h3eed52aa, 32'h3c96f6d4} /* (2, 11, 22) {real, imag} */,
  {32'hbe2e3806, 32'h3edeedac} /* (2, 11, 21) {real, imag} */,
  {32'h3e3b2d34, 32'h3cdbb608} /* (2, 11, 20) {real, imag} */,
  {32'h3a429e00, 32'h3e5a7cd4} /* (2, 11, 19) {real, imag} */,
  {32'h3e993444, 32'hbd4771e8} /* (2, 11, 18) {real, imag} */,
  {32'hbe0f21e6, 32'hbdf487d9} /* (2, 11, 17) {real, imag} */,
  {32'hbd5b6788, 32'h3eb19e82} /* (2, 11, 16) {real, imag} */,
  {32'hbd6ab7b8, 32'h3df6ca36} /* (2, 11, 15) {real, imag} */,
  {32'h3e57970c, 32'h3e5f68fe} /* (2, 11, 14) {real, imag} */,
  {32'hbe9a8fa0, 32'hbdc2fc27} /* (2, 11, 13) {real, imag} */,
  {32'h3d9f56b1, 32'hbd3609f4} /* (2, 11, 12) {real, imag} */,
  {32'h3e43509c, 32'hbea2aa90} /* (2, 11, 11) {real, imag} */,
  {32'h3d70c590, 32'hbdf58f2a} /* (2, 11, 10) {real, imag} */,
  {32'h3eaa1890, 32'hbe56139b} /* (2, 11, 9) {real, imag} */,
  {32'h3efa817c, 32'hbf00c014} /* (2, 11, 8) {real, imag} */,
  {32'hbe39bb5b, 32'hbcdd1108} /* (2, 11, 7) {real, imag} */,
  {32'hbc36be80, 32'hbc8b53d0} /* (2, 11, 6) {real, imag} */,
  {32'h3ea38fa2, 32'h3d3ccc18} /* (2, 11, 5) {real, imag} */,
  {32'h3e7e8260, 32'hbe951a90} /* (2, 11, 4) {real, imag} */,
  {32'h3d9c9bb6, 32'h3ed340b8} /* (2, 11, 3) {real, imag} */,
  {32'hbcc124f0, 32'hbf0fba86} /* (2, 11, 2) {real, imag} */,
  {32'h3e950630, 32'h3f242e12} /* (2, 11, 1) {real, imag} */,
  {32'h3eb469dc, 32'h3ea93396} /* (2, 11, 0) {real, imag} */,
  {32'h3d640ef4, 32'hbe140576} /* (2, 10, 31) {real, imag} */,
  {32'h3eb4688d, 32'h3f452bea} /* (2, 10, 30) {real, imag} */,
  {32'hbf167067, 32'h3e6d43c3} /* (2, 10, 29) {real, imag} */,
  {32'hbf21e576, 32'hbdab89c0} /* (2, 10, 28) {real, imag} */,
  {32'h3e0272f6, 32'hbd2c3246} /* (2, 10, 27) {real, imag} */,
  {32'h3e6af2d5, 32'hbe3bca7f} /* (2, 10, 26) {real, imag} */,
  {32'hbe2ab2c3, 32'hbe0dad3a} /* (2, 10, 25) {real, imag} */,
  {32'hbee505a2, 32'hbe37af91} /* (2, 10, 24) {real, imag} */,
  {32'hbe36b027, 32'hbe9d074b} /* (2, 10, 23) {real, imag} */,
  {32'hbeeca7f2, 32'hbc7cc3e0} /* (2, 10, 22) {real, imag} */,
  {32'hbdad610c, 32'hbf25b692} /* (2, 10, 21) {real, imag} */,
  {32'hbdd4028c, 32'h3df47258} /* (2, 10, 20) {real, imag} */,
  {32'h3eae2f0a, 32'hbf27b408} /* (2, 10, 19) {real, imag} */,
  {32'h3df2225e, 32'h3ebd9596} /* (2, 10, 18) {real, imag} */,
  {32'hbec3f2f8, 32'hbc4ecd68} /* (2, 10, 17) {real, imag} */,
  {32'h3e95e3f7, 32'h3e3b5cc8} /* (2, 10, 16) {real, imag} */,
  {32'h3c3d2228, 32'hbe5d7372} /* (2, 10, 15) {real, imag} */,
  {32'h3ddb1868, 32'hbd640ea8} /* (2, 10, 14) {real, imag} */,
  {32'h3e00f4e8, 32'hbf094c5c} /* (2, 10, 13) {real, imag} */,
  {32'hbed48b1e, 32'hbdae6715} /* (2, 10, 12) {real, imag} */,
  {32'hbe6962f4, 32'hbf16297a} /* (2, 10, 11) {real, imag} */,
  {32'h3f0e1da1, 32'h3de0f4ee} /* (2, 10, 10) {real, imag} */,
  {32'h3e7d4cbf, 32'h3f0818b2} /* (2, 10, 9) {real, imag} */,
  {32'hbeda52f2, 32'h3e2761d4} /* (2, 10, 8) {real, imag} */,
  {32'h3ea4ffbc, 32'h3d953900} /* (2, 10, 7) {real, imag} */,
  {32'h3ef4b908, 32'hbe43f601} /* (2, 10, 6) {real, imag} */,
  {32'h3b9514e0, 32'h3ed1916e} /* (2, 10, 5) {real, imag} */,
  {32'h3c7972a8, 32'h3ea0fe8f} /* (2, 10, 4) {real, imag} */,
  {32'h3f51fe31, 32'h3d9f0d0e} /* (2, 10, 3) {real, imag} */,
  {32'hbeea6a0a, 32'h3f18ed13} /* (2, 10, 2) {real, imag} */,
  {32'hbf235a44, 32'hbebe38d8} /* (2, 10, 1) {real, imag} */,
  {32'h3efee158, 32'hbea28b36} /* (2, 10, 0) {real, imag} */,
  {32'h3ee18f6c, 32'h3e236b1b} /* (2, 9, 31) {real, imag} */,
  {32'h3ede5689, 32'h3f55a3cb} /* (2, 9, 30) {real, imag} */,
  {32'hbc887320, 32'hbe7e949e} /* (2, 9, 29) {real, imag} */,
  {32'h3e2edf54, 32'h3dbee195} /* (2, 9, 28) {real, imag} */,
  {32'h3f1f648f, 32'h3e9d3858} /* (2, 9, 27) {real, imag} */,
  {32'h3ea0bcd6, 32'hbd85d455} /* (2, 9, 26) {real, imag} */,
  {32'hbddafe68, 32'hbd438a10} /* (2, 9, 25) {real, imag} */,
  {32'hbec3e457, 32'h3dc5fdf8} /* (2, 9, 24) {real, imag} */,
  {32'h3d8433e4, 32'hbd8d001e} /* (2, 9, 23) {real, imag} */,
  {32'h3d3e1a2a, 32'h3cfb5d38} /* (2, 9, 22) {real, imag} */,
  {32'hbe5e5bd8, 32'h3f09042c} /* (2, 9, 21) {real, imag} */,
  {32'hbf0f57a3, 32'hbe2e70ea} /* (2, 9, 20) {real, imag} */,
  {32'hbe981f7c, 32'h3df661ab} /* (2, 9, 19) {real, imag} */,
  {32'h3f5158db, 32'hbd82c7c2} /* (2, 9, 18) {real, imag} */,
  {32'hbe8a31cd, 32'hbe5ac8f3} /* (2, 9, 17) {real, imag} */,
  {32'h3e23887c, 32'h3e94810c} /* (2, 9, 16) {real, imag} */,
  {32'hbed5590c, 32'h3ebe7896} /* (2, 9, 15) {real, imag} */,
  {32'hbed47af4, 32'h3ea99f77} /* (2, 9, 14) {real, imag} */,
  {32'h3eabaef6, 32'hbdb07e73} /* (2, 9, 13) {real, imag} */,
  {32'hbf2bb034, 32'h3e8a4675} /* (2, 9, 12) {real, imag} */,
  {32'hbe2a84de, 32'h3f060715} /* (2, 9, 11) {real, imag} */,
  {32'hbe987cda, 32'hbcd01440} /* (2, 9, 10) {real, imag} */,
  {32'h3eb26b84, 32'h3e24bb01} /* (2, 9, 9) {real, imag} */,
  {32'hbecd9aeb, 32'hbd03aaf6} /* (2, 9, 8) {real, imag} */,
  {32'hbd2aa3ec, 32'hbe32d79c} /* (2, 9, 7) {real, imag} */,
  {32'hbd9f40ed, 32'h3f37eaa1} /* (2, 9, 6) {real, imag} */,
  {32'hbea2f81e, 32'hbf2e8e61} /* (2, 9, 5) {real, imag} */,
  {32'hbea039f0, 32'hbed57300} /* (2, 9, 4) {real, imag} */,
  {32'hbf3ba9c5, 32'h3efc9595} /* (2, 9, 3) {real, imag} */,
  {32'h3e12d7fa, 32'hbec7a555} /* (2, 9, 2) {real, imag} */,
  {32'hbf1094c7, 32'hbf5e04b6} /* (2, 9, 1) {real, imag} */,
  {32'hbedba0ba, 32'hbf0a62da} /* (2, 9, 0) {real, imag} */,
  {32'h3fbfe59d, 32'h3f1a4594} /* (2, 8, 31) {real, imag} */,
  {32'hbf8cfa02, 32'h3f6694d0} /* (2, 8, 30) {real, imag} */,
  {32'hbf1fb35e, 32'hbf0e88a5} /* (2, 8, 29) {real, imag} */,
  {32'h3d3b2d59, 32'h3f49c9f2} /* (2, 8, 28) {real, imag} */,
  {32'hbd06ab10, 32'hbe1bc73a} /* (2, 8, 27) {real, imag} */,
  {32'h3ebd1d6f, 32'h3eef7384} /* (2, 8, 26) {real, imag} */,
  {32'h3f0faff6, 32'h3f4dd8e2} /* (2, 8, 25) {real, imag} */,
  {32'h3e101ce9, 32'h3f2225b7} /* (2, 8, 24) {real, imag} */,
  {32'h3f3f32c0, 32'h3e7bc8dc} /* (2, 8, 23) {real, imag} */,
  {32'hbd8cda56, 32'hbf6a78f4} /* (2, 8, 22) {real, imag} */,
  {32'h3e02e90b, 32'hbed33d32} /* (2, 8, 21) {real, imag} */,
  {32'h3eb3342d, 32'hbe68bfe0} /* (2, 8, 20) {real, imag} */,
  {32'hbd99d4fa, 32'h3f1023ba} /* (2, 8, 19) {real, imag} */,
  {32'h3b63d300, 32'hbe27d313} /* (2, 8, 18) {real, imag} */,
  {32'h3e468b38, 32'hbe497ef6} /* (2, 8, 17) {real, imag} */,
  {32'h3d949860, 32'h3f0a1288} /* (2, 8, 16) {real, imag} */,
  {32'h3e11d26a, 32'h3edb532d} /* (2, 8, 15) {real, imag} */,
  {32'hbd5336d8, 32'hbe9dd96e} /* (2, 8, 14) {real, imag} */,
  {32'hbe24a334, 32'hbeb60167} /* (2, 8, 13) {real, imag} */,
  {32'h3f12fbcb, 32'hbdbda9a6} /* (2, 8, 12) {real, imag} */,
  {32'hbe927c2a, 32'hbf4461f6} /* (2, 8, 11) {real, imag} */,
  {32'hbc47f550, 32'h3eaa5696} /* (2, 8, 10) {real, imag} */,
  {32'hbee676e3, 32'h3f407b0d} /* (2, 8, 9) {real, imag} */,
  {32'hbde98978, 32'hbb918130} /* (2, 8, 8) {real, imag} */,
  {32'hbf29fc84, 32'hbed41de4} /* (2, 8, 7) {real, imag} */,
  {32'hbebaf802, 32'hbf70b3d3} /* (2, 8, 6) {real, imag} */,
  {32'h3d8b8650, 32'hbddba5de} /* (2, 8, 5) {real, imag} */,
  {32'h3d8c1e7c, 32'h3d8461c4} /* (2, 8, 4) {real, imag} */,
  {32'hbdcdde4a, 32'hbcd2aa68} /* (2, 8, 3) {real, imag} */,
  {32'h3e2734a7, 32'hbf454375} /* (2, 8, 2) {real, imag} */,
  {32'h3ee902b0, 32'h3f750973} /* (2, 8, 1) {real, imag} */,
  {32'h3e7aa4c2, 32'h3d8992f0} /* (2, 8, 0) {real, imag} */,
  {32'hbe426dd5, 32'h3dc963f4} /* (2, 7, 31) {real, imag} */,
  {32'hbd269134, 32'hbe6a0951} /* (2, 7, 30) {real, imag} */,
  {32'hbf2cc2b0, 32'hbec5907c} /* (2, 7, 29) {real, imag} */,
  {32'hbf01c744, 32'h3dc42776} /* (2, 7, 28) {real, imag} */,
  {32'h3d0119c0, 32'h3ed95507} /* (2, 7, 27) {real, imag} */,
  {32'hbd3aaf78, 32'h3e8a8f43} /* (2, 7, 26) {real, imag} */,
  {32'hbee43679, 32'h3f307d50} /* (2, 7, 25) {real, imag} */,
  {32'h3d9ac684, 32'h3d44d5a2} /* (2, 7, 24) {real, imag} */,
  {32'hbf3c1c48, 32'h3e62cba6} /* (2, 7, 23) {real, imag} */,
  {32'hbefd8217, 32'h3ebaff4a} /* (2, 7, 22) {real, imag} */,
  {32'h3e5f7bbe, 32'h3e337c92} /* (2, 7, 21) {real, imag} */,
  {32'h3cd7bca0, 32'hbdc2dc70} /* (2, 7, 20) {real, imag} */,
  {32'h3ed15753, 32'hbe34edfa} /* (2, 7, 19) {real, imag} */,
  {32'hbeb51c5b, 32'h3dae3b68} /* (2, 7, 18) {real, imag} */,
  {32'h3e706de8, 32'hbe69b89e} /* (2, 7, 17) {real, imag} */,
  {32'hbe37e982, 32'h3e0d246c} /* (2, 7, 16) {real, imag} */,
  {32'h3ec19d14, 32'hbd535672} /* (2, 7, 15) {real, imag} */,
  {32'hbee6df53, 32'hbed91c12} /* (2, 7, 14) {real, imag} */,
  {32'h3de53529, 32'h3e85883c} /* (2, 7, 13) {real, imag} */,
  {32'h3d5d95f0, 32'hbdabb37a} /* (2, 7, 12) {real, imag} */,
  {32'hbed772f4, 32'hbe90dfd7} /* (2, 7, 11) {real, imag} */,
  {32'h3ec4f5cb, 32'h3f567524} /* (2, 7, 10) {real, imag} */,
  {32'h3eb6064f, 32'h3eef7157} /* (2, 7, 9) {real, imag} */,
  {32'hbe12352e, 32'hbea3e63d} /* (2, 7, 8) {real, imag} */,
  {32'h3e2cf734, 32'h3dd9a068} /* (2, 7, 7) {real, imag} */,
  {32'hbe4600fe, 32'hbe2677f6} /* (2, 7, 6) {real, imag} */,
  {32'hbc38ad50, 32'h3eed54a2} /* (2, 7, 5) {real, imag} */,
  {32'hbe6aa11a, 32'hbee703ce} /* (2, 7, 4) {real, imag} */,
  {32'h3ed40ffa, 32'h3ddf7ff5} /* (2, 7, 3) {real, imag} */,
  {32'hbec20da0, 32'h3ee273dc} /* (2, 7, 2) {real, imag} */,
  {32'hbf025b20, 32'hbeb25113} /* (2, 7, 1) {real, imag} */,
  {32'h3d16af50, 32'hbed53c41} /* (2, 7, 0) {real, imag} */,
  {32'hbea15b1a, 32'h3f0164d5} /* (2, 6, 31) {real, imag} */,
  {32'hbd146e00, 32'hbe7da365} /* (2, 6, 30) {real, imag} */,
  {32'h3eaa4c3a, 32'h3e92bf4c} /* (2, 6, 29) {real, imag} */,
  {32'hbf44d0d5, 32'hbf40d341} /* (2, 6, 28) {real, imag} */,
  {32'h3d4f3b7e, 32'hbf648fdc} /* (2, 6, 27) {real, imag} */,
  {32'h3e23e206, 32'hbe98681d} /* (2, 6, 26) {real, imag} */,
  {32'hbe9718a6, 32'hbdcfb7dc} /* (2, 6, 25) {real, imag} */,
  {32'hbe383389, 32'h3f1d6487} /* (2, 6, 24) {real, imag} */,
  {32'hbeca77ae, 32'h3e06a392} /* (2, 6, 23) {real, imag} */,
  {32'h3eec288f, 32'hbeb4ecea} /* (2, 6, 22) {real, imag} */,
  {32'hbd3a5e68, 32'h3e20e058} /* (2, 6, 21) {real, imag} */,
  {32'h3e9db68c, 32'h3eab7e73} /* (2, 6, 20) {real, imag} */,
  {32'h3e75d092, 32'h3955fc00} /* (2, 6, 19) {real, imag} */,
  {32'hbdfb883a, 32'hbe9c2f56} /* (2, 6, 18) {real, imag} */,
  {32'hbe6dd045, 32'h3dca342e} /* (2, 6, 17) {real, imag} */,
  {32'h3c2766e0, 32'hbe9d811d} /* (2, 6, 16) {real, imag} */,
  {32'h3d55a3c0, 32'hbdc0acfd} /* (2, 6, 15) {real, imag} */,
  {32'hbd78361a, 32'hbebd399a} /* (2, 6, 14) {real, imag} */,
  {32'hbe874c1c, 32'h3e7d7acb} /* (2, 6, 13) {real, imag} */,
  {32'hbf067ea1, 32'hbed555f3} /* (2, 6, 12) {real, imag} */,
  {32'h3ec9d4e2, 32'hbe1715d6} /* (2, 6, 11) {real, imag} */,
  {32'h3f1efe4b, 32'hbdadf6e0} /* (2, 6, 10) {real, imag} */,
  {32'hbb84da00, 32'h3f2a2bf2} /* (2, 6, 9) {real, imag} */,
  {32'hbe8830ee, 32'hbe392f8c} /* (2, 6, 8) {real, imag} */,
  {32'hbe1e0792, 32'h3f042dd0} /* (2, 6, 7) {real, imag} */,
  {32'hbe8756ac, 32'h3e193721} /* (2, 6, 6) {real, imag} */,
  {32'h3ddca074, 32'hbc5403c0} /* (2, 6, 5) {real, imag} */,
  {32'h3e26ed69, 32'hbe08ef7d} /* (2, 6, 4) {real, imag} */,
  {32'hb7c04000, 32'hbd28bd04} /* (2, 6, 3) {real, imag} */,
  {32'hbe74f1c0, 32'hbf3ae389} /* (2, 6, 2) {real, imag} */,
  {32'h3e5e2112, 32'hbeba4cd4} /* (2, 6, 1) {real, imag} */,
  {32'h3f07d9f9, 32'h3e9d8f51} /* (2, 6, 0) {real, imag} */,
  {32'h404374f4, 32'h3e62deb0} /* (2, 5, 31) {real, imag} */,
  {32'hbfcd1080, 32'hbf3cd08a} /* (2, 5, 30) {real, imag} */,
  {32'hbe1d0e2e, 32'h3ec35bb5} /* (2, 5, 29) {real, imag} */,
  {32'h3e935a02, 32'hbeb2de17} /* (2, 5, 28) {real, imag} */,
  {32'hbf7852a9, 32'h3e072b6d} /* (2, 5, 27) {real, imag} */,
  {32'h3eaddb16, 32'hbef89de1} /* (2, 5, 26) {real, imag} */,
  {32'hbe2a7ce8, 32'h3d950796} /* (2, 5, 25) {real, imag} */,
  {32'h3d44bdd4, 32'h3f524eee} /* (2, 5, 24) {real, imag} */,
  {32'hbe78e73d, 32'h3ec5bba7} /* (2, 5, 23) {real, imag} */,
  {32'hbe47007e, 32'hbdf92480} /* (2, 5, 22) {real, imag} */,
  {32'hbe74f15c, 32'h3e724d09} /* (2, 5, 21) {real, imag} */,
  {32'hbe7c73f5, 32'hbd73d980} /* (2, 5, 20) {real, imag} */,
  {32'h3dae8e9a, 32'h3c4b9d50} /* (2, 5, 19) {real, imag} */,
  {32'hbf0e74c7, 32'h3de30a50} /* (2, 5, 18) {real, imag} */,
  {32'hbdd1213a, 32'h3e011b00} /* (2, 5, 17) {real, imag} */,
  {32'h3e91e5e0, 32'hbe56248c} /* (2, 5, 16) {real, imag} */,
  {32'hbe886afb, 32'h3e47f49f} /* (2, 5, 15) {real, imag} */,
  {32'hbcdf6284, 32'hbeb53fc7} /* (2, 5, 14) {real, imag} */,
  {32'h3e8012bd, 32'h3eb48675} /* (2, 5, 13) {real, imag} */,
  {32'hbdc72d94, 32'hbdcae2e4} /* (2, 5, 12) {real, imag} */,
  {32'hbdd27d98, 32'h3e18d8da} /* (2, 5, 11) {real, imag} */,
  {32'h3e4af08c, 32'hbd580a00} /* (2, 5, 10) {real, imag} */,
  {32'hbe82b1ad, 32'h3e9ed95f} /* (2, 5, 9) {real, imag} */,
  {32'hbd162258, 32'hbe96aa06} /* (2, 5, 8) {real, imag} */,
  {32'hbf651ffa, 32'h3e7d9fb2} /* (2, 5, 7) {real, imag} */,
  {32'h3dabcdac, 32'hbe40f16b} /* (2, 5, 6) {real, imag} */,
  {32'hbf1e7668, 32'hbf32d0ee} /* (2, 5, 5) {real, imag} */,
  {32'hbe4cd964, 32'hbe51a49e} /* (2, 5, 4) {real, imag} */,
  {32'hbdb30576, 32'hbe8a9a44} /* (2, 5, 3) {real, imag} */,
  {32'h3d236350, 32'hbef6ef05} /* (2, 5, 2) {real, imag} */,
  {32'h4011edd5, 32'h404a7164} /* (2, 5, 1) {real, imag} */,
  {32'h4031a711, 32'h3f3409b8} /* (2, 5, 0) {real, imag} */,
  {32'hc0041c49, 32'hc00e6902} /* (2, 4, 31) {real, imag} */,
  {32'h3f095e18, 32'h402dbd78} /* (2, 4, 30) {real, imag} */,
  {32'hbee2ad07, 32'h3e440cc0} /* (2, 4, 29) {real, imag} */,
  {32'hbf7ad8bc, 32'hbf5225da} /* (2, 4, 28) {real, imag} */,
  {32'h3f621601, 32'h3eea027e} /* (2, 4, 27) {real, imag} */,
  {32'h3ec98ca3, 32'hbf23b74d} /* (2, 4, 26) {real, imag} */,
  {32'hbe8b6d49, 32'hbf1ae8d8} /* (2, 4, 25) {real, imag} */,
  {32'h3de39b4b, 32'hbf03ca5a} /* (2, 4, 24) {real, imag} */,
  {32'hbeacb2fe, 32'hbe923672} /* (2, 4, 23) {real, imag} */,
  {32'hbe742a00, 32'h3eb98fe1} /* (2, 4, 22) {real, imag} */,
  {32'h3f4e5102, 32'hbe6da2c0} /* (2, 4, 21) {real, imag} */,
  {32'h3ddd6d09, 32'hbeaa590e} /* (2, 4, 20) {real, imag} */,
  {32'hbf07d80d, 32'hbbfef6f0} /* (2, 4, 19) {real, imag} */,
  {32'hbec61abe, 32'hbea18f56} /* (2, 4, 18) {real, imag} */,
  {32'hbdb70de8, 32'hbe6665e8} /* (2, 4, 17) {real, imag} */,
  {32'h3e35f934, 32'h3e0b0111} /* (2, 4, 16) {real, imag} */,
  {32'h3e1db033, 32'hbdddb040} /* (2, 4, 15) {real, imag} */,
  {32'h3ec32590, 32'h3ce3aff8} /* (2, 4, 14) {real, imag} */,
  {32'h3eea7e04, 32'h3ea0ecc4} /* (2, 4, 13) {real, imag} */,
  {32'h3e66bf48, 32'h3e077e5e} /* (2, 4, 12) {real, imag} */,
  {32'hbe235982, 32'h3e5e1908} /* (2, 4, 11) {real, imag} */,
  {32'hbdf81cf6, 32'hbcd35630} /* (2, 4, 10) {real, imag} */,
  {32'h3e8ee724, 32'hbdfdff68} /* (2, 4, 9) {real, imag} */,
  {32'hbe6594d2, 32'h3f1eab97} /* (2, 4, 8) {real, imag} */,
  {32'hbf1b42ef, 32'h3e2b6100} /* (2, 4, 7) {real, imag} */,
  {32'h3e8d8a5e, 32'h3e99e61c} /* (2, 4, 6) {real, imag} */,
  {32'hbe7d19a4, 32'h3db4b3c8} /* (2, 4, 5) {real, imag} */,
  {32'hbd776008, 32'hbdf663f8} /* (2, 4, 4) {real, imag} */,
  {32'h3cb979d8, 32'h3f0945fd} /* (2, 4, 3) {real, imag} */,
  {32'h404fc2b9, 32'h4064f8c0} /* (2, 4, 2) {real, imag} */,
  {32'hc0b43598, 32'hbfcadba7} /* (2, 4, 1) {real, imag} */,
  {32'hc00863b4, 32'hbf268f73} /* (2, 4, 0) {real, imag} */,
  {32'h409f3a08, 32'hc0344ce4} /* (2, 3, 31) {real, imag} */,
  {32'hc0173cba, 32'h400ef77f} /* (2, 3, 30) {real, imag} */,
  {32'hbfa7278c, 32'hbf5b0308} /* (2, 3, 29) {real, imag} */,
  {32'hbdd3c17c, 32'hbeaf335c} /* (2, 3, 28) {real, imag} */,
  {32'h3dbd9806, 32'h3e6c0c68} /* (2, 3, 27) {real, imag} */,
  {32'h3e43fa4c, 32'h3edda79e} /* (2, 3, 26) {real, imag} */,
  {32'hbe901cc3, 32'h3e6f7cab} /* (2, 3, 25) {real, imag} */,
  {32'hbe716765, 32'h3f3aff6c} /* (2, 3, 24) {real, imag} */,
  {32'hbeb04b02, 32'hbf87833b} /* (2, 3, 23) {real, imag} */,
  {32'hbc9c84b2, 32'h3e3cbd52} /* (2, 3, 22) {real, imag} */,
  {32'hbd04c948, 32'hbe5d0195} /* (2, 3, 21) {real, imag} */,
  {32'hbe6a4bf8, 32'h3f11a97e} /* (2, 3, 20) {real, imag} */,
  {32'hbd728ede, 32'h3e60d55c} /* (2, 3, 19) {real, imag} */,
  {32'h3dc5b7aa, 32'hbce7d948} /* (2, 3, 18) {real, imag} */,
  {32'h3ead34a8, 32'hbe8ebe38} /* (2, 3, 17) {real, imag} */,
  {32'hbe2ea740, 32'hbe4d155c} /* (2, 3, 16) {real, imag} */,
  {32'h3e25ce7a, 32'hbecbbb35} /* (2, 3, 15) {real, imag} */,
  {32'h3e7bec9c, 32'h3f223d2e} /* (2, 3, 14) {real, imag} */,
  {32'h3a919280, 32'h3e64f9c9} /* (2, 3, 13) {real, imag} */,
  {32'h3f10bf80, 32'hbe2be3f5} /* (2, 3, 12) {real, imag} */,
  {32'hbdb4dfe4, 32'hbedf0747} /* (2, 3, 11) {real, imag} */,
  {32'h3f1c9116, 32'h3ec80c61} /* (2, 3, 10) {real, imag} */,
  {32'h3d84f7df, 32'hbb559fc0} /* (2, 3, 9) {real, imag} */,
  {32'hbda3ce2b, 32'h3efaed6a} /* (2, 3, 8) {real, imag} */,
  {32'h3f035836, 32'hbef16260} /* (2, 3, 7) {real, imag} */,
  {32'hbf38addb, 32'h3dd97af5} /* (2, 3, 6) {real, imag} */,
  {32'hbf5bc29f, 32'h3f952930} /* (2, 3, 5) {real, imag} */,
  {32'h3f642d9d, 32'h3ec7f2b6} /* (2, 3, 4) {real, imag} */,
  {32'hbfcc7612, 32'hbf8b7d8f} /* (2, 3, 3) {real, imag} */,
  {32'hbf0db9a5, 32'h40961d4e} /* (2, 3, 2) {real, imag} */,
  {32'hc0382e10, 32'hbf87d672} /* (2, 3, 1) {real, imag} */,
  {32'h3f8173f0, 32'hbf7a2460} /* (2, 3, 0) {real, imag} */,
  {32'h41b4eca6, 32'h400fcaa9} /* (2, 2, 31) {real, imag} */,
  {32'hc13249c6, 32'h401af864} /* (2, 2, 30) {real, imag} */,
  {32'h3fcee380, 32'h3f53104c} /* (2, 2, 29) {real, imag} */,
  {32'h3fceb7cb, 32'hbfbcfc89} /* (2, 2, 28) {real, imag} */,
  {32'hbf86e118, 32'h3fdcccc6} /* (2, 2, 27) {real, imag} */,
  {32'h3e0bec05, 32'hbebcc014} /* (2, 2, 26) {real, imag} */,
  {32'h3e3a5829, 32'hbea17e15} /* (2, 2, 25) {real, imag} */,
  {32'hbfa6c5cf, 32'h3f7a9ce7} /* (2, 2, 24) {real, imag} */,
  {32'hbea2e60a, 32'hbe801244} /* (2, 2, 23) {real, imag} */,
  {32'hbe89b59e, 32'hbf23d72c} /* (2, 2, 22) {real, imag} */,
  {32'hbe46ffd5, 32'h3f455133} /* (2, 2, 21) {real, imag} */,
  {32'h3e7e08b0, 32'h3dee65f0} /* (2, 2, 20) {real, imag} */,
  {32'hbe56a184, 32'h3dbb0f18} /* (2, 2, 19) {real, imag} */,
  {32'hbe9f2aeb, 32'h3d087d60} /* (2, 2, 18) {real, imag} */,
  {32'h3df66859, 32'hbe999c0a} /* (2, 2, 17) {real, imag} */,
  {32'hbd9b6993, 32'hbebe64ba} /* (2, 2, 16) {real, imag} */,
  {32'hbdde694b, 32'hbea9fd95} /* (2, 2, 15) {real, imag} */,
  {32'hbce1e188, 32'hbeee348c} /* (2, 2, 14) {real, imag} */,
  {32'h3e5f7c14, 32'hbc37d33c} /* (2, 2, 13) {real, imag} */,
  {32'h3e6155bc, 32'h3f0125af} /* (2, 2, 12) {real, imag} */,
  {32'hbcf416b0, 32'hbe9a876e} /* (2, 2, 11) {real, imag} */,
  {32'h3f62c600, 32'h3f551546} /* (2, 2, 10) {real, imag} */,
  {32'h3d8c895c, 32'h3e3a4594} /* (2, 2, 9) {real, imag} */,
  {32'hbf6abcf3, 32'h3ec75f89} /* (2, 2, 8) {real, imag} */,
  {32'hbb4a1c60, 32'h3e319e9c} /* (2, 2, 7) {real, imag} */,
  {32'hbf23c7fa, 32'hbeedf2fa} /* (2, 2, 6) {real, imag} */,
  {32'hbfc5dc90, 32'hbfba7fcf} /* (2, 2, 5) {real, imag} */,
  {32'h404dc345, 32'h3f535bdc} /* (2, 2, 4) {real, imag} */,
  {32'hbf8ddc1e, 32'hbf73b55d} /* (2, 2, 3) {real, imag} */,
  {32'hc0ff12ef, 32'h40988f98} /* (2, 2, 2) {real, imag} */,
  {32'h41344612, 32'hbe3d3590} /* (2, 2, 1) {real, imag} */,
  {32'h4122e7b4, 32'h405a7243} /* (2, 2, 0) {real, imag} */,
  {32'hc19f114e, 32'h4058475e} /* (2, 1, 31) {real, imag} */,
  {32'h40f6d04c, 32'h3f80fcee} /* (2, 1, 30) {real, imag} */,
  {32'h3fc721b1, 32'hbfa2b064} /* (2, 1, 29) {real, imag} */,
  {32'hc03afd8c, 32'hbfb203bd} /* (2, 1, 28) {real, imag} */,
  {32'h4084ef9c, 32'hbddfabef} /* (2, 1, 27) {real, imag} */,
  {32'h3f97b59e, 32'hbefa58a0} /* (2, 1, 26) {real, imag} */,
  {32'hbd98bdc8, 32'h3e39249a} /* (2, 1, 25) {real, imag} */,
  {32'h3f65e12a, 32'hbe4913ce} /* (2, 1, 24) {real, imag} */,
  {32'h3e4952ea, 32'hbe1471c9} /* (2, 1, 23) {real, imag} */,
  {32'hbec762d8, 32'h3e9302f3} /* (2, 1, 22) {real, imag} */,
  {32'h3f98df18, 32'hbef2fb38} /* (2, 1, 21) {real, imag} */,
  {32'hbde56644, 32'h3f00bf32} /* (2, 1, 20) {real, imag} */,
  {32'hbec0ea95, 32'hbea28405} /* (2, 1, 19) {real, imag} */,
  {32'hbe5a80d5, 32'hbe1335a7} /* (2, 1, 18) {real, imag} */,
  {32'hbdcc8e17, 32'hbecbe896} /* (2, 1, 17) {real, imag} */,
  {32'hbe923ff8, 32'h3df6a105} /* (2, 1, 16) {real, imag} */,
  {32'h3da1b65a, 32'hbe17137f} /* (2, 1, 15) {real, imag} */,
  {32'hbd52ac05, 32'h3e87a08e} /* (2, 1, 14) {real, imag} */,
  {32'hbd9c7f60, 32'hbef8d327} /* (2, 1, 13) {real, imag} */,
  {32'h3efb333c, 32'hbd6dfbac} /* (2, 1, 12) {real, imag} */,
  {32'h3ef4ad1b, 32'h3ecc2a32} /* (2, 1, 11) {real, imag} */,
  {32'h3eda6014, 32'hbe0ffaf9} /* (2, 1, 10) {real, imag} */,
  {32'hbdc21ad4, 32'hbdd26afe} /* (2, 1, 9) {real, imag} */,
  {32'h3f334014, 32'h3f684d50} /* (2, 1, 8) {real, imag} */,
  {32'hbe58990b, 32'hbf3c837d} /* (2, 1, 7) {real, imag} */,
  {32'hbd84efc0, 32'h3c28db40} /* (2, 1, 6) {real, imag} */,
  {32'h3fd29f59, 32'h3fdbb22c} /* (2, 1, 5) {real, imag} */,
  {32'hbec22e86, 32'hbf7c6dd4} /* (2, 1, 4) {real, imag} */,
  {32'h3fdfb448, 32'hbf2572b7} /* (2, 1, 3) {real, imag} */,
  {32'h4123d54f, 32'h4108fcd8} /* (2, 1, 2) {real, imag} */,
  {32'hc1e907cd, 32'hc193725e} /* (2, 1, 1) {real, imag} */,
  {32'hc17f6ad2, 32'h3fe409e0} /* (2, 1, 0) {real, imag} */,
  {32'hc15cc43f, 32'h410dbc6d} /* (2, 0, 31) {real, imag} */,
  {32'h3fc4186a, 32'hc059a97f} /* (2, 0, 30) {real, imag} */,
  {32'h3fde9dc8, 32'hbfbf6985} /* (2, 0, 29) {real, imag} */,
  {32'hbf431f38, 32'hc02140fc} /* (2, 0, 28) {real, imag} */,
  {32'h3fc95d5a, 32'hbef539ec} /* (2, 0, 27) {real, imag} */,
  {32'hbe2d891a, 32'h3f22a445} /* (2, 0, 26) {real, imag} */,
  {32'hbd0dd2e0, 32'h3f815abd} /* (2, 0, 25) {real, imag} */,
  {32'h3f3504e8, 32'hbf18807d} /* (2, 0, 24) {real, imag} */,
  {32'h3e47f683, 32'hbe144859} /* (2, 0, 23) {real, imag} */,
  {32'h3f02a5e5, 32'hbeecd5ec} /* (2, 0, 22) {real, imag} */,
  {32'h3e94ceee, 32'hbf1d0e7c} /* (2, 0, 21) {real, imag} */,
  {32'hbda36602, 32'h3d4e0100} /* (2, 0, 20) {real, imag} */,
  {32'h3e06c8c0, 32'h3e817cc7} /* (2, 0, 19) {real, imag} */,
  {32'hbe59c974, 32'hbdb6fda0} /* (2, 0, 18) {real, imag} */,
  {32'h3e84ae48, 32'hbe3609ac} /* (2, 0, 17) {real, imag} */,
  {32'hbd0dcba4, 32'h00000000} /* (2, 0, 16) {real, imag} */,
  {32'h3e84ae48, 32'h3e3609ac} /* (2, 0, 15) {real, imag} */,
  {32'hbe59c974, 32'h3db6fda0} /* (2, 0, 14) {real, imag} */,
  {32'h3e06c8c0, 32'hbe817cc7} /* (2, 0, 13) {real, imag} */,
  {32'hbda36602, 32'hbd4e0100} /* (2, 0, 12) {real, imag} */,
  {32'h3e94ceee, 32'h3f1d0e7c} /* (2, 0, 11) {real, imag} */,
  {32'h3f02a5e5, 32'h3eecd5ec} /* (2, 0, 10) {real, imag} */,
  {32'h3e47f683, 32'h3e144859} /* (2, 0, 9) {real, imag} */,
  {32'h3f3504e8, 32'h3f18807d} /* (2, 0, 8) {real, imag} */,
  {32'hbd0dd2e0, 32'hbf815abd} /* (2, 0, 7) {real, imag} */,
  {32'hbe2d891a, 32'hbf22a445} /* (2, 0, 6) {real, imag} */,
  {32'h3fc95d5a, 32'h3ef539ec} /* (2, 0, 5) {real, imag} */,
  {32'hbf431f38, 32'h402140fc} /* (2, 0, 4) {real, imag} */,
  {32'h3fde9dc8, 32'h3fbf6985} /* (2, 0, 3) {real, imag} */,
  {32'h3fc4186a, 32'h4059a97f} /* (2, 0, 2) {real, imag} */,
  {32'hc15cc43f, 32'hc10dbc6d} /* (2, 0, 1) {real, imag} */,
  {32'hc06389c6, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc1c06709, 32'h417a5546} /* (1, 31, 31) {real, imag} */,
  {32'h410ca72a, 32'hc0e7a1a0} /* (1, 31, 30) {real, imag} */,
  {32'h3ff2a66d, 32'hbe36f578} /* (1, 31, 29) {real, imag} */,
  {32'h3ebed3af, 32'h3fa88e11} /* (1, 31, 28) {real, imag} */,
  {32'h3ff1ea94, 32'hbf93293c} /* (1, 31, 27) {real, imag} */,
  {32'h3eb2f384, 32'hbecff0a1} /* (1, 31, 26) {real, imag} */,
  {32'hbee6e3e4, 32'h3f816cbe} /* (1, 31, 25) {real, imag} */,
  {32'h3ee78477, 32'hbee9f1c1} /* (1, 31, 24) {real, imag} */,
  {32'hbe6e5500, 32'hbf42b294} /* (1, 31, 23) {real, imag} */,
  {32'hbe7a3e6b, 32'h3ecd8960} /* (1, 31, 22) {real, imag} */,
  {32'hbe8a07af, 32'hbdf5b93a} /* (1, 31, 21) {real, imag} */,
  {32'h3e99a388, 32'h3e185f5d} /* (1, 31, 20) {real, imag} */,
  {32'hbeb885de, 32'hbd5a0810} /* (1, 31, 19) {real, imag} */,
  {32'hbe4cf26a, 32'hbec8672d} /* (1, 31, 18) {real, imag} */,
  {32'h3e7bf15b, 32'h3dfbf001} /* (1, 31, 17) {real, imag} */,
  {32'hbb465be0, 32'hbd1acad8} /* (1, 31, 16) {real, imag} */,
  {32'hbda598f4, 32'hbe0488f5} /* (1, 31, 15) {real, imag} */,
  {32'hbcc04404, 32'h3d029cc4} /* (1, 31, 14) {real, imag} */,
  {32'h3db06312, 32'hbb88d180} /* (1, 31, 13) {real, imag} */,
  {32'hbda15bc4, 32'h3e155167} /* (1, 31, 12) {real, imag} */,
  {32'h3f0e4ef0, 32'h3f076ade} /* (1, 31, 11) {real, imag} */,
  {32'hbebc61bc, 32'h3d6ceea2} /* (1, 31, 10) {real, imag} */,
  {32'hbe09ee3c, 32'h3f2f7294} /* (1, 31, 9) {real, imag} */,
  {32'h3f8fce5a, 32'h3f4885b3} /* (1, 31, 8) {real, imag} */,
  {32'hbf2bf0db, 32'h3dbb6654} /* (1, 31, 7) {real, imag} */,
  {32'h3e9ffd6c, 32'h3e825ed4} /* (1, 31, 6) {real, imag} */,
  {32'h406dde0b, 32'h3dfa27d4} /* (1, 31, 5) {real, imag} */,
  {32'hc029ed83, 32'h3f157882} /* (1, 31, 4) {real, imag} */,
  {32'h3f5b8bbf, 32'h3f148293} /* (1, 31, 3) {real, imag} */,
  {32'h40b0976e, 32'h3ef7ed99} /* (1, 31, 2) {real, imag} */,
  {32'hc183a91f, 32'hbfec4749} /* (1, 31, 1) {real, imag} */,
  {32'hc17707f3, 32'hc0052fc4} /* (1, 31, 0) {real, imag} */,
  {32'h41020a3a, 32'hbdcc3680} /* (1, 30, 31) {real, imag} */,
  {32'hc0dea3d9, 32'hc0601cae} /* (1, 30, 30) {real, imag} */,
  {32'hbd314b08, 32'h3fa1752f} /* (1, 30, 29) {real, imag} */,
  {32'h4059c255, 32'hbf014f84} /* (1, 30, 28) {real, imag} */,
  {32'hbfb43e4e, 32'h3f96daa0} /* (1, 30, 27) {real, imag} */,
  {32'hbdc4de90, 32'hbe54c3b8} /* (1, 30, 26) {real, imag} */,
  {32'h3e7c76e6, 32'hbf489424} /* (1, 30, 25) {real, imag} */,
  {32'hbfb0dda9, 32'h3f50ae8d} /* (1, 30, 24) {real, imag} */,
  {32'h3e0f55cc, 32'h3e3d88ce} /* (1, 30, 23) {real, imag} */,
  {32'hbd3afe7c, 32'h3dabc9de} /* (1, 30, 22) {real, imag} */,
  {32'hbe858d7c, 32'h3f0e832c} /* (1, 30, 21) {real, imag} */,
  {32'hbe3e1710, 32'hbe6d7e51} /* (1, 30, 20) {real, imag} */,
  {32'h3c03dd34, 32'h3c9152d4} /* (1, 30, 19) {real, imag} */,
  {32'h3e929baf, 32'h3e25698b} /* (1, 30, 18) {real, imag} */,
  {32'hbc9697ac, 32'hbdb2f798} /* (1, 30, 17) {real, imag} */,
  {32'hbdcf1f28, 32'hbe163c10} /* (1, 30, 16) {real, imag} */,
  {32'h3c4c8e70, 32'h3e080d63} /* (1, 30, 15) {real, imag} */,
  {32'hbe72bc28, 32'h3e1c15e1} /* (1, 30, 14) {real, imag} */,
  {32'hbe0ebab4, 32'h3f0e5fca} /* (1, 30, 13) {real, imag} */,
  {32'h3ddab3fc, 32'hbd0af4f2} /* (1, 30, 12) {real, imag} */,
  {32'hbe558bcb, 32'hbe9e36ee} /* (1, 30, 11) {real, imag} */,
  {32'hbd9d6ec2, 32'h3f2495f4} /* (1, 30, 10) {real, imag} */,
  {32'hbe9d502c, 32'hbcbfbcd8} /* (1, 30, 9) {real, imag} */,
  {32'hbf84197a, 32'hbf8f10a5} /* (1, 30, 8) {real, imag} */,
  {32'hbb077180, 32'h3e9fc5a6} /* (1, 30, 7) {real, imag} */,
  {32'h3e5584f0, 32'h3d05f77c} /* (1, 30, 6) {real, imag} */,
  {32'hbf8dfeb2, 32'hbfd8bd12} /* (1, 30, 5) {real, imag} */,
  {32'h3faede74, 32'h3f10ddc8} /* (1, 30, 4) {real, imag} */,
  {32'h3f6ac239, 32'h3f3057f4} /* (1, 30, 3) {real, imag} */,
  {32'hc1141f88, 32'hbf2755ad} /* (1, 30, 2) {real, imag} */,
  {32'h418f74bf, 32'hbffa5ecc} /* (1, 30, 1) {real, imag} */,
  {32'h40fe832c, 32'hc0109d07} /* (1, 30, 0) {real, imag} */,
  {32'hbfe040ab, 32'h3fb0f71b} /* (1, 29, 31) {real, imag} */,
  {32'hbeed933c, 32'hc0810ee2} /* (1, 29, 30) {real, imag} */,
  {32'hbc8ea8a0, 32'h3fd76169} /* (1, 29, 29) {real, imag} */,
  {32'h3f4f4536, 32'hbf76624c} /* (1, 29, 28) {real, imag} */,
  {32'hbf8aa5ba, 32'hbf4c3352} /* (1, 29, 27) {real, imag} */,
  {32'hbf6c64a1, 32'h3e643823} /* (1, 29, 26) {real, imag} */,
  {32'hbeb7f387, 32'h3e896234} /* (1, 29, 25) {real, imag} */,
  {32'hbf480f7f, 32'hbe6ac2d3} /* (1, 29, 24) {real, imag} */,
  {32'h3eaf9e06, 32'h3e6396cd} /* (1, 29, 23) {real, imag} */,
  {32'h3ef1946d, 32'h3e0d1c7c} /* (1, 29, 22) {real, imag} */,
  {32'h3cb590bc, 32'hbe03afda} /* (1, 29, 21) {real, imag} */,
  {32'h3f83e9a2, 32'hbe86bbfa} /* (1, 29, 20) {real, imag} */,
  {32'hbd4c04a8, 32'h3d039dfa} /* (1, 29, 19) {real, imag} */,
  {32'h3e517a24, 32'hbc200a20} /* (1, 29, 18) {real, imag} */,
  {32'hbdf62f1f, 32'h3e25abd8} /* (1, 29, 17) {real, imag} */,
  {32'hbe28feef, 32'h3e23aef1} /* (1, 29, 16) {real, imag} */,
  {32'h3e2b0b36, 32'h3e5f740f} /* (1, 29, 15) {real, imag} */,
  {32'hbe8159bf, 32'h3e3b8e81} /* (1, 29, 14) {real, imag} */,
  {32'hbe9d04f2, 32'h3ab47c80} /* (1, 29, 13) {real, imag} */,
  {32'hbdd8362d, 32'h3e67449f} /* (1, 29, 12) {real, imag} */,
  {32'h3e138120, 32'hbd6ea84c} /* (1, 29, 11) {real, imag} */,
  {32'h3dac2f60, 32'hbe4cea51} /* (1, 29, 10) {real, imag} */,
  {32'hbd84dfec, 32'h3dc41726} /* (1, 29, 9) {real, imag} */,
  {32'h3e256d94, 32'hbf56d76b} /* (1, 29, 8) {real, imag} */,
  {32'hbe610c0c, 32'h3d5f7c08} /* (1, 29, 7) {real, imag} */,
  {32'hbeed045e, 32'h3e381de8} /* (1, 29, 6) {real, imag} */,
  {32'h3f0a60e2, 32'hbe48ee59} /* (1, 29, 5) {real, imag} */,
  {32'hbf3d8d26, 32'h3e61d365} /* (1, 29, 4) {real, imag} */,
  {32'h3dfeba0c, 32'hbe625ee6} /* (1, 29, 3) {real, imag} */,
  {32'hbfbd3fcd, 32'hc01f93e2} /* (1, 29, 2) {real, imag} */,
  {32'h4071bf5d, 32'h3fe6f6e8} /* (1, 29, 1) {real, imag} */,
  {32'h3f83a094, 32'h3e019160} /* (1, 29, 0) {real, imag} */,
  {32'hc08950b2, 32'h3f08f442} /* (1, 28, 31) {real, imag} */,
  {32'h3ff95d7a, 32'hc04ce668} /* (1, 28, 30) {real, imag} */,
  {32'hbe1bed98, 32'hbf60093c} /* (1, 28, 29) {real, imag} */,
  {32'hbe437dfe, 32'h3dfeace4} /* (1, 28, 28) {real, imag} */,
  {32'h3ede9a6a, 32'h3e6fd804} /* (1, 28, 27) {real, imag} */,
  {32'h3ea2613e, 32'h3e8287ca} /* (1, 28, 26) {real, imag} */,
  {32'hbdc7fb76, 32'h3f41493c} /* (1, 28, 25) {real, imag} */,
  {32'h3e9a62b5, 32'hbeced2bc} /* (1, 28, 24) {real, imag} */,
  {32'h3f157666, 32'h3dc939f8} /* (1, 28, 23) {real, imag} */,
  {32'h3f0bf991, 32'h3ebd8b50} /* (1, 28, 22) {real, imag} */,
  {32'h3ec2196a, 32'hbf41e220} /* (1, 28, 21) {real, imag} */,
  {32'h3c93d7b0, 32'h3efc6572} /* (1, 28, 20) {real, imag} */,
  {32'hbdac4d18, 32'hbdbd7285} /* (1, 28, 19) {real, imag} */,
  {32'hbebf8ab7, 32'hbe848f24} /* (1, 28, 18) {real, imag} */,
  {32'h3e419fd7, 32'h3e6b5ae4} /* (1, 28, 17) {real, imag} */,
  {32'hbd17e2d1, 32'hbd8ae2d4} /* (1, 28, 16) {real, imag} */,
  {32'hbd724d82, 32'h3e8b8125} /* (1, 28, 15) {real, imag} */,
  {32'h3de64002, 32'hbe3a67af} /* (1, 28, 14) {real, imag} */,
  {32'hbe060f2a, 32'hbeb8a946} /* (1, 28, 13) {real, imag} */,
  {32'h3bbb6dc0, 32'hbee3625f} /* (1, 28, 12) {real, imag} */,
  {32'h3e4aad7f, 32'hbc98db48} /* (1, 28, 11) {real, imag} */,
  {32'hbe71c418, 32'h3e4049ac} /* (1, 28, 10) {real, imag} */,
  {32'hbea8a5ea, 32'h3d1d3c5e} /* (1, 28, 9) {real, imag} */,
  {32'hbe30c3f8, 32'hbe519bf0} /* (1, 28, 8) {real, imag} */,
  {32'hbeda273c, 32'h3e693c79} /* (1, 28, 7) {real, imag} */,
  {32'h3ebffdc7, 32'h3ee4533c} /* (1, 28, 6) {real, imag} */,
  {32'h3f06b53a, 32'h3e8bf7db} /* (1, 28, 5) {real, imag} */,
  {32'hbf479f2d, 32'h3e90a672} /* (1, 28, 4) {real, imag} */,
  {32'hbf20dca4, 32'h3f657670} /* (1, 28, 3) {real, imag} */,
  {32'h3fb6463c, 32'hc02a9da4} /* (1, 28, 2) {real, imag} */,
  {32'hc0015b13, 32'h3f83face} /* (1, 28, 1) {real, imag} */,
  {32'hbe736c28, 32'h3eec282c} /* (1, 28, 0) {real, imag} */,
  {32'h3f94f23c, 32'hc0198b9e} /* (1, 27, 31) {real, imag} */,
  {32'h3ed07e1a, 32'h3f1984ec} /* (1, 27, 30) {real, imag} */,
  {32'hbea82c4a, 32'h3eb3fcdf} /* (1, 27, 29) {real, imag} */,
  {32'hbdba54a4, 32'hbe73e479} /* (1, 27, 28) {real, imag} */,
  {32'hbf2f9810, 32'h3f5ca75e} /* (1, 27, 27) {real, imag} */,
  {32'hbdc50b38, 32'h3d3aa5f8} /* (1, 27, 26) {real, imag} */,
  {32'h3e83a914, 32'hbf228b1a} /* (1, 27, 25) {real, imag} */,
  {32'hbea3b4e2, 32'hbe0c542b} /* (1, 27, 24) {real, imag} */,
  {32'h3e397122, 32'hbe86fcf1} /* (1, 27, 23) {real, imag} */,
  {32'hbde429e1, 32'h3e420fee} /* (1, 27, 22) {real, imag} */,
  {32'hbddcc620, 32'h3dc7cae0} /* (1, 27, 21) {real, imag} */,
  {32'hbe2ce988, 32'hbe1df586} /* (1, 27, 20) {real, imag} */,
  {32'h3f546830, 32'hbe95de7e} /* (1, 27, 19) {real, imag} */,
  {32'hbd93eb5b, 32'hbdaba0ec} /* (1, 27, 18) {real, imag} */,
  {32'hbe191f49, 32'h3ddd1643} /* (1, 27, 17) {real, imag} */,
  {32'hbe57aec0, 32'hbe4d419e} /* (1, 27, 16) {real, imag} */,
  {32'hbe7e8df4, 32'h3cbb0b80} /* (1, 27, 15) {real, imag} */,
  {32'h3e2c25ed, 32'hbf29d7fd} /* (1, 27, 14) {real, imag} */,
  {32'h3ea58f90, 32'hbd8d1d31} /* (1, 27, 13) {real, imag} */,
  {32'h3ed9a23e, 32'h3f2dbab0} /* (1, 27, 12) {real, imag} */,
  {32'hbd74e636, 32'h3e2f373e} /* (1, 27, 11) {real, imag} */,
  {32'hbeef3ca9, 32'h3ddb2a3c} /* (1, 27, 10) {real, imag} */,
  {32'h3de67237, 32'h3e4235e6} /* (1, 27, 9) {real, imag} */,
  {32'h3ee0eb45, 32'h3e2859c1} /* (1, 27, 8) {real, imag} */,
  {32'hbeca9a49, 32'hbdcac330} /* (1, 27, 7) {real, imag} */,
  {32'hbe89540c, 32'h3e0659a0} /* (1, 27, 6) {real, imag} */,
  {32'h3e14e870, 32'hbe708b84} /* (1, 27, 5) {real, imag} */,
  {32'h3e500b12, 32'hbdf7c8c4} /* (1, 27, 4) {real, imag} */,
  {32'hbf1c3c64, 32'hbefe0336} /* (1, 27, 3) {real, imag} */,
  {32'hbfd200b2, 32'h3e5a0a54} /* (1, 27, 2) {real, imag} */,
  {32'h403a7a75, 32'hbe263c01} /* (1, 27, 1) {real, imag} */,
  {32'h3fe9f865, 32'hbf62d3fc} /* (1, 27, 0) {real, imag} */,
  {32'hbe6b1d73, 32'hbef8f41f} /* (1, 26, 31) {real, imag} */,
  {32'hbd13083a, 32'h3edae54e} /* (1, 26, 30) {real, imag} */,
  {32'hbe12ce66, 32'h3e0a7b99} /* (1, 26, 29) {real, imag} */,
  {32'h3ebb8db3, 32'h3e3f7a34} /* (1, 26, 28) {real, imag} */,
  {32'hbe6cd2ec, 32'hbe050018} /* (1, 26, 27) {real, imag} */,
  {32'hbeaf52bc, 32'h3eaeacde} /* (1, 26, 26) {real, imag} */,
  {32'h3f0ed710, 32'h3ee9b823} /* (1, 26, 25) {real, imag} */,
  {32'h3e4fa023, 32'h3e1d5f82} /* (1, 26, 24) {real, imag} */,
  {32'h3eb633a2, 32'hbf37881c} /* (1, 26, 23) {real, imag} */,
  {32'h3e556ef7, 32'h3e1f2bea} /* (1, 26, 22) {real, imag} */,
  {32'hbe710ea5, 32'h3f171586} /* (1, 26, 21) {real, imag} */,
  {32'h3d704aa6, 32'hbc0ce738} /* (1, 26, 20) {real, imag} */,
  {32'hbec98a73, 32'h3e5e144f} /* (1, 26, 19) {real, imag} */,
  {32'hbd4c8d94, 32'hbde8828c} /* (1, 26, 18) {real, imag} */,
  {32'hbe872f8b, 32'h3ddf33f3} /* (1, 26, 17) {real, imag} */,
  {32'h3d872552, 32'h3d54d534} /* (1, 26, 16) {real, imag} */,
  {32'h3e285ce6, 32'h3e494e18} /* (1, 26, 15) {real, imag} */,
  {32'h39760f00, 32'h3c5447c0} /* (1, 26, 14) {real, imag} */,
  {32'h3d4664c8, 32'h3ead85a8} /* (1, 26, 13) {real, imag} */,
  {32'h3d8c5642, 32'h3d2782f4} /* (1, 26, 12) {real, imag} */,
  {32'hbed40b4a, 32'h3d0ce6bc} /* (1, 26, 11) {real, imag} */,
  {32'h3e03d81e, 32'h3e0a2866} /* (1, 26, 10) {real, imag} */,
  {32'hbf0ffe2d, 32'hbf014d38} /* (1, 26, 9) {real, imag} */,
  {32'h3d6e86fe, 32'hbdf2c71c} /* (1, 26, 8) {real, imag} */,
  {32'h3e43a154, 32'h3d421e1b} /* (1, 26, 7) {real, imag} */,
  {32'h3ecbbdc4, 32'hbec9a774} /* (1, 26, 6) {real, imag} */,
  {32'h3f34d0f1, 32'h3f72a08a} /* (1, 26, 5) {real, imag} */,
  {32'hbeefda0e, 32'h3e61da77} /* (1, 26, 4) {real, imag} */,
  {32'h3eb0fbe8, 32'h3e9f8ea8} /* (1, 26, 3) {real, imag} */,
  {32'hbf4789eb, 32'hbea017b4} /* (1, 26, 2) {real, imag} */,
  {32'hbec4f184, 32'hbf9b40b0} /* (1, 26, 1) {real, imag} */,
  {32'h3f0e5d0a, 32'h3f636aa2} /* (1, 26, 0) {real, imag} */,
  {32'h3f51151a, 32'h3f277e1e} /* (1, 25, 31) {real, imag} */,
  {32'hbf098137, 32'h3ed01e73} /* (1, 25, 30) {real, imag} */,
  {32'hbd8dc441, 32'hbd85942c} /* (1, 25, 29) {real, imag} */,
  {32'hbda17e03, 32'h3e0ebd06} /* (1, 25, 28) {real, imag} */,
  {32'hbc8f3640, 32'hbe9815ef} /* (1, 25, 27) {real, imag} */,
  {32'hbf139ba1, 32'hbf14fb68} /* (1, 25, 26) {real, imag} */,
  {32'hbec0ddf4, 32'hbe99bf2a} /* (1, 25, 25) {real, imag} */,
  {32'h3e1f2ec5, 32'hbde935d6} /* (1, 25, 24) {real, imag} */,
  {32'h3f22f6a7, 32'hbe0d7394} /* (1, 25, 23) {real, imag} */,
  {32'h3c101f30, 32'hbefc68e1} /* (1, 25, 22) {real, imag} */,
  {32'h3d22fd10, 32'hbeb0e3ca} /* (1, 25, 21) {real, imag} */,
  {32'hbe1b811c, 32'h3f16de2e} /* (1, 25, 20) {real, imag} */,
  {32'h3d0da13a, 32'hbea7c5aa} /* (1, 25, 19) {real, imag} */,
  {32'h3e9d5ff9, 32'hbdc141d7} /* (1, 25, 18) {real, imag} */,
  {32'h3e13ccde, 32'h3e49dbf3} /* (1, 25, 17) {real, imag} */,
  {32'h3d43da76, 32'hbe907443} /* (1, 25, 16) {real, imag} */,
  {32'h3d791e88, 32'hbeaf13bb} /* (1, 25, 15) {real, imag} */,
  {32'hbe3a4bcd, 32'hbd06f212} /* (1, 25, 14) {real, imag} */,
  {32'h3c799620, 32'h3e1bcc8e} /* (1, 25, 13) {real, imag} */,
  {32'h3daa86cc, 32'hbed1c43b} /* (1, 25, 12) {real, imag} */,
  {32'hbe8bd851, 32'hbea4799c} /* (1, 25, 11) {real, imag} */,
  {32'hbe2d12c5, 32'hbda14859} /* (1, 25, 10) {real, imag} */,
  {32'hbe7f30e0, 32'hbf058c34} /* (1, 25, 9) {real, imag} */,
  {32'h3f0c6722, 32'h3f104206} /* (1, 25, 8) {real, imag} */,
  {32'h3ed27864, 32'hbe2e0394} /* (1, 25, 7) {real, imag} */,
  {32'h3ef3035a, 32'hbe218678} /* (1, 25, 6) {real, imag} */,
  {32'h3e2cac73, 32'h3eca0fa9} /* (1, 25, 5) {real, imag} */,
  {32'hbf18e080, 32'hbf71ff0b} /* (1, 25, 4) {real, imag} */,
  {32'hbd84dc1e, 32'h3e850fda} /* (1, 25, 3) {real, imag} */,
  {32'h3ea01c43, 32'h3e006194} /* (1, 25, 2) {real, imag} */,
  {32'hbec03e15, 32'hbeac4c32} /* (1, 25, 1) {real, imag} */,
  {32'h3e024878, 32'h3ec38335} /* (1, 25, 0) {real, imag} */,
  {32'h3f1cd2fe, 32'hbf401539} /* (1, 24, 31) {real, imag} */,
  {32'h3e613ea0, 32'hbd68a410} /* (1, 24, 30) {real, imag} */,
  {32'hbd517810, 32'hbe700332} /* (1, 24, 29) {real, imag} */,
  {32'hbedb42a8, 32'hbef91a5c} /* (1, 24, 28) {real, imag} */,
  {32'hba003180, 32'h3f99c8b8} /* (1, 24, 27) {real, imag} */,
  {32'hbe86b9b5, 32'h3e113d61} /* (1, 24, 26) {real, imag} */,
  {32'h3d3b497f, 32'hbead7771} /* (1, 24, 25) {real, imag} */,
  {32'h3e16c6ec, 32'h3f0f1c30} /* (1, 24, 24) {real, imag} */,
  {32'h3f0db74a, 32'hbebae5c8} /* (1, 24, 23) {real, imag} */,
  {32'h3b716b40, 32'hbf4d9fa6} /* (1, 24, 22) {real, imag} */,
  {32'h3f1fb2e6, 32'h3e8c34c1} /* (1, 24, 21) {real, imag} */,
  {32'hbe1d7f00, 32'h3f0003a6} /* (1, 24, 20) {real, imag} */,
  {32'hbec76b29, 32'h3eff3d72} /* (1, 24, 19) {real, imag} */,
  {32'h3e3cf9d0, 32'h3e3dc29b} /* (1, 24, 18) {real, imag} */,
  {32'h3e960138, 32'hbd13f65a} /* (1, 24, 17) {real, imag} */,
  {32'hbeac6ca6, 32'hbc416e00} /* (1, 24, 16) {real, imag} */,
  {32'h3e1d2dd6, 32'hbd424678} /* (1, 24, 15) {real, imag} */,
  {32'h3e0cc3fa, 32'hbe20d0de} /* (1, 24, 14) {real, imag} */,
  {32'hbe6085cb, 32'h3f17b956} /* (1, 24, 13) {real, imag} */,
  {32'hbede279d, 32'hbeb590d4} /* (1, 24, 12) {real, imag} */,
  {32'hbd768dac, 32'hbdf1b8b4} /* (1, 24, 11) {real, imag} */,
  {32'hbf06bce8, 32'h3ec06f47} /* (1, 24, 10) {real, imag} */,
  {32'h3f4b5f18, 32'hbe1d946a} /* (1, 24, 9) {real, imag} */,
  {32'hbe3b3142, 32'hbf2aee09} /* (1, 24, 8) {real, imag} */,
  {32'h3f8aba94, 32'hbdfd6eb3} /* (1, 24, 7) {real, imag} */,
  {32'hbdad3904, 32'hbed929c0} /* (1, 24, 6) {real, imag} */,
  {32'hbd4df8dc, 32'hbe8ff2a9} /* (1, 24, 5) {real, imag} */,
  {32'hbe086cff, 32'hbe45847c} /* (1, 24, 4) {real, imag} */,
  {32'hbdc4f1d9, 32'h3e1179f8} /* (1, 24, 3) {real, imag} */,
  {32'hbfd29dcf, 32'hbe4b78a6} /* (1, 24, 2) {real, imag} */,
  {32'h3f711a69, 32'hbee74c57} /* (1, 24, 1) {real, imag} */,
  {32'h3ebd11e8, 32'hbf603a32} /* (1, 24, 0) {real, imag} */,
  {32'hbe8e552b, 32'h3db52514} /* (1, 23, 31) {real, imag} */,
  {32'h3ec125ce, 32'hbed3bd05} /* (1, 23, 30) {real, imag} */,
  {32'hbebb5cc7, 32'hbed64c92} /* (1, 23, 29) {real, imag} */,
  {32'h3ed68702, 32'h3ec87c8b} /* (1, 23, 28) {real, imag} */,
  {32'hbcf27446, 32'hbd02ba00} /* (1, 23, 27) {real, imag} */,
  {32'hbe6ab588, 32'h3eaf42f8} /* (1, 23, 26) {real, imag} */,
  {32'hbde6a554, 32'hbdb3650c} /* (1, 23, 25) {real, imag} */,
  {32'hbdebf525, 32'hbd6850dc} /* (1, 23, 24) {real, imag} */,
  {32'h3ea3a31c, 32'h3c9b3600} /* (1, 23, 23) {real, imag} */,
  {32'hbe725d7b, 32'h3c3173b0} /* (1, 23, 22) {real, imag} */,
  {32'hbf08f3f8, 32'h3e5abfc4} /* (1, 23, 21) {real, imag} */,
  {32'h3e277d6e, 32'h3e39f892} /* (1, 23, 20) {real, imag} */,
  {32'h3e8361fd, 32'hbeb7fa8a} /* (1, 23, 19) {real, imag} */,
  {32'hbe871240, 32'h3f54cd14} /* (1, 23, 18) {real, imag} */,
  {32'hbe3abfc1, 32'h3dc43745} /* (1, 23, 17) {real, imag} */,
  {32'h3eb7ba78, 32'hbefe5414} /* (1, 23, 16) {real, imag} */,
  {32'h3ea02ca9, 32'h3e4af2c9} /* (1, 23, 15) {real, imag} */,
  {32'h3f3e3707, 32'hbe75d65e} /* (1, 23, 14) {real, imag} */,
  {32'hbe5e9e70, 32'hbdeec3e7} /* (1, 23, 13) {real, imag} */,
  {32'h3dbbc618, 32'h3f3530d8} /* (1, 23, 12) {real, imag} */,
  {32'h3e059c0c, 32'h3bd5aaf0} /* (1, 23, 11) {real, imag} */,
  {32'h3cf499f0, 32'hbea83ca4} /* (1, 23, 10) {real, imag} */,
  {32'h3e16b32a, 32'h3e727178} /* (1, 23, 9) {real, imag} */,
  {32'hbd69bc28, 32'h3e9b5c50} /* (1, 23, 8) {real, imag} */,
  {32'hbea9d2a1, 32'hbdb3779c} /* (1, 23, 7) {real, imag} */,
  {32'h3eb5482e, 32'h3ee84416} /* (1, 23, 6) {real, imag} */,
  {32'hbe88f268, 32'h3d6878b4} /* (1, 23, 5) {real, imag} */,
  {32'hbe0fa4fa, 32'h3edb21b0} /* (1, 23, 4) {real, imag} */,
  {32'hbf1aaf46, 32'h3ee3bcd9} /* (1, 23, 3) {real, imag} */,
  {32'h3ea44570, 32'hbf3205d8} /* (1, 23, 2) {real, imag} */,
  {32'h3de2b852, 32'h3d913358} /* (1, 23, 1) {real, imag} */,
  {32'hbf0a8538, 32'h3e12a964} /* (1, 23, 0) {real, imag} */,
  {32'h3ea4812f, 32'h3e220dbf} /* (1, 22, 31) {real, imag} */,
  {32'h3f05fbdb, 32'hbf409c35} /* (1, 22, 30) {real, imag} */,
  {32'h3f2beed9, 32'h3df4c832} /* (1, 22, 29) {real, imag} */,
  {32'h3eb88261, 32'hbd9e7290} /* (1, 22, 28) {real, imag} */,
  {32'hbeb70d5d, 32'h3e3b5a28} /* (1, 22, 27) {real, imag} */,
  {32'hbd4c6432, 32'h3eacfd34} /* (1, 22, 26) {real, imag} */,
  {32'h3e9007c5, 32'hbd577bb0} /* (1, 22, 25) {real, imag} */,
  {32'hbe86cf96, 32'h3de35627} /* (1, 22, 24) {real, imag} */,
  {32'h3f5539bd, 32'hbd419654} /* (1, 22, 23) {real, imag} */,
  {32'h3e66bda4, 32'h3cb19d40} /* (1, 22, 22) {real, imag} */,
  {32'hbd974a9a, 32'hbe92cf26} /* (1, 22, 21) {real, imag} */,
  {32'hbef039fe, 32'h3d673fb8} /* (1, 22, 20) {real, imag} */,
  {32'h3e47dd2e, 32'hbe2fccbd} /* (1, 22, 19) {real, imag} */,
  {32'hbe8a1818, 32'h3eb61ec6} /* (1, 22, 18) {real, imag} */,
  {32'hbd6fd5d6, 32'hbe569edb} /* (1, 22, 17) {real, imag} */,
  {32'h3c739c9c, 32'hbbe57490} /* (1, 22, 16) {real, imag} */,
  {32'h3e41586e, 32'h3d2b7cf1} /* (1, 22, 15) {real, imag} */,
  {32'h3bc0de80, 32'h3bd88c80} /* (1, 22, 14) {real, imag} */,
  {32'h3e94d66d, 32'hbe5c6843} /* (1, 22, 13) {real, imag} */,
  {32'hbded2d71, 32'h3e92f8aa} /* (1, 22, 12) {real, imag} */,
  {32'hbf2299eb, 32'hbd6abe00} /* (1, 22, 11) {real, imag} */,
  {32'h3db7e58a, 32'hbe870906} /* (1, 22, 10) {real, imag} */,
  {32'h3e319b6c, 32'h3e8c05bb} /* (1, 22, 9) {real, imag} */,
  {32'h3f138efc, 32'hbef740eb} /* (1, 22, 8) {real, imag} */,
  {32'hbee56ea3, 32'hbbf80170} /* (1, 22, 7) {real, imag} */,
  {32'hbdec8cce, 32'hbdecba56} /* (1, 22, 6) {real, imag} */,
  {32'hbe5a165a, 32'hbe301014} /* (1, 22, 5) {real, imag} */,
  {32'hbe18bc94, 32'h3f3ffd7a} /* (1, 22, 4) {real, imag} */,
  {32'hbec099ad, 32'h3d0339dc} /* (1, 22, 3) {real, imag} */,
  {32'hbe442deb, 32'hbf0f3aab} /* (1, 22, 2) {real, imag} */,
  {32'hbe216149, 32'h3f0bf583} /* (1, 22, 1) {real, imag} */,
  {32'hbe16715b, 32'h3df40b1b} /* (1, 22, 0) {real, imag} */,
  {32'h3e96c5a9, 32'hbf4648ba} /* (1, 21, 31) {real, imag} */,
  {32'h3c238630, 32'h3e87bf42} /* (1, 21, 30) {real, imag} */,
  {32'hbe7573c7, 32'h3e654a0e} /* (1, 21, 29) {real, imag} */,
  {32'h3e2159ee, 32'h3ead5863} /* (1, 21, 28) {real, imag} */,
  {32'hbf04e76e, 32'h3dd4e9f2} /* (1, 21, 27) {real, imag} */,
  {32'h3eb61936, 32'h3e4d924a} /* (1, 21, 26) {real, imag} */,
  {32'hbdb74810, 32'h3ed55ec7} /* (1, 21, 25) {real, imag} */,
  {32'hbe125c6d, 32'hbe5715ce} /* (1, 21, 24) {real, imag} */,
  {32'hbe3ab9c7, 32'h3e992834} /* (1, 21, 23) {real, imag} */,
  {32'hbf21cfdc, 32'h3e25002c} /* (1, 21, 22) {real, imag} */,
  {32'hbf55a5ba, 32'h3ed70f54} /* (1, 21, 21) {real, imag} */,
  {32'hbe089dd6, 32'hbdadd05c} /* (1, 21, 20) {real, imag} */,
  {32'h3e369232, 32'h3dff284b} /* (1, 21, 19) {real, imag} */,
  {32'hbe1e9db6, 32'hbe3ef119} /* (1, 21, 18) {real, imag} */,
  {32'hbe082d6a, 32'hbd3e56e0} /* (1, 21, 17) {real, imag} */,
  {32'h3e89c370, 32'hbda20bdc} /* (1, 21, 16) {real, imag} */,
  {32'h3ea69198, 32'hbd5c752e} /* (1, 21, 15) {real, imag} */,
  {32'hbdf1b51a, 32'hbd439730} /* (1, 21, 14) {real, imag} */,
  {32'hbe11bad0, 32'h3eefd6a0} /* (1, 21, 13) {real, imag} */,
  {32'hbf3f550b, 32'hbf1f608a} /* (1, 21, 12) {real, imag} */,
  {32'h3e3f6a4e, 32'h3d9f6de8} /* (1, 21, 11) {real, imag} */,
  {32'h3df4b7d0, 32'hbecb9166} /* (1, 21, 10) {real, imag} */,
  {32'h3f20f686, 32'h3f64d2bc} /* (1, 21, 9) {real, imag} */,
  {32'h3d9c4ec0, 32'h3d4a48ec} /* (1, 21, 8) {real, imag} */,
  {32'hbe594781, 32'hbe2d65be} /* (1, 21, 7) {real, imag} */,
  {32'h3ee688b1, 32'hbe3b41a2} /* (1, 21, 6) {real, imag} */,
  {32'h3d20cf58, 32'h3ea62851} /* (1, 21, 5) {real, imag} */,
  {32'h3deb047d, 32'hbdceeba6} /* (1, 21, 4) {real, imag} */,
  {32'hbea9e59b, 32'hbdbd3033} /* (1, 21, 3) {real, imag} */,
  {32'h3d891694, 32'h3f82ebab} /* (1, 21, 2) {real, imag} */,
  {32'h3efd130a, 32'hbee8a13c} /* (1, 21, 1) {real, imag} */,
  {32'h3e86cab6, 32'hbbc904c0} /* (1, 21, 0) {real, imag} */,
  {32'h3edafe84, 32'h3d278650} /* (1, 20, 31) {real, imag} */,
  {32'h3da84aac, 32'h3e340a9f} /* (1, 20, 30) {real, imag} */,
  {32'hbe5596ab, 32'h3de06392} /* (1, 20, 29) {real, imag} */,
  {32'h3ea7c00e, 32'h3e9d6d54} /* (1, 20, 28) {real, imag} */,
  {32'h3ed4e110, 32'h3abb1200} /* (1, 20, 27) {real, imag} */,
  {32'h3e9ea700, 32'hbd259c4c} /* (1, 20, 26) {real, imag} */,
  {32'hbf05950c, 32'hbeb5006d} /* (1, 20, 25) {real, imag} */,
  {32'h3ee6a2ab, 32'h3e2997a6} /* (1, 20, 24) {real, imag} */,
  {32'hbd5d60de, 32'hbf007a08} /* (1, 20, 23) {real, imag} */,
  {32'hbe8c87b4, 32'h3f0a885e} /* (1, 20, 22) {real, imag} */,
  {32'h3da01b1c, 32'hbe59f333} /* (1, 20, 21) {real, imag} */,
  {32'hbeb4c4c5, 32'hbe28c624} /* (1, 20, 20) {real, imag} */,
  {32'hbe26bb34, 32'hbd7504d3} /* (1, 20, 19) {real, imag} */,
  {32'h3dbc29ca, 32'hbeb17393} /* (1, 20, 18) {real, imag} */,
  {32'h3dcc12c5, 32'hbdf38f18} /* (1, 20, 17) {real, imag} */,
  {32'hbe7647b9, 32'h3ec6b940} /* (1, 20, 16) {real, imag} */,
  {32'hbe5c62fa, 32'hbe7995c8} /* (1, 20, 15) {real, imag} */,
  {32'h3d0aa540, 32'hbe1df7e2} /* (1, 20, 14) {real, imag} */,
  {32'h3e231b11, 32'hbe3d6a6e} /* (1, 20, 13) {real, imag} */,
  {32'h3eb542f0, 32'hbf035dbf} /* (1, 20, 12) {real, imag} */,
  {32'hbe98bac0, 32'hbf298280} /* (1, 20, 11) {real, imag} */,
  {32'h3ec28a1a, 32'hbf2a89dc} /* (1, 20, 10) {real, imag} */,
  {32'h3e953e57, 32'hbef73b13} /* (1, 20, 9) {real, imag} */,
  {32'hbb8c2fb0, 32'hbd7305ec} /* (1, 20, 8) {real, imag} */,
  {32'h3d780acc, 32'hbcc45540} /* (1, 20, 7) {real, imag} */,
  {32'hbd5d55ae, 32'h3f0abd73} /* (1, 20, 6) {real, imag} */,
  {32'h3e86f25d, 32'hbf0b4dc0} /* (1, 20, 5) {real, imag} */,
  {32'hbe62cd9b, 32'hbe40ab02} /* (1, 20, 4) {real, imag} */,
  {32'hbdf79448, 32'h3ec215a5} /* (1, 20, 3) {real, imag} */,
  {32'h3eb45048, 32'h3e8616d7} /* (1, 20, 2) {real, imag} */,
  {32'h3d92b59a, 32'h3e94729c} /* (1, 20, 1) {real, imag} */,
  {32'hbcf62a40, 32'h3ecad71e} /* (1, 20, 0) {real, imag} */,
  {32'hbda56825, 32'h3ec57fcc} /* (1, 19, 31) {real, imag} */,
  {32'h3e3ecfec, 32'h3d8ac2fe} /* (1, 19, 30) {real, imag} */,
  {32'h3d635e22, 32'h3e30e12a} /* (1, 19, 29) {real, imag} */,
  {32'hbf052c0b, 32'hbd591d9e} /* (1, 19, 28) {real, imag} */,
  {32'hbe6af962, 32'hbebe858a} /* (1, 19, 27) {real, imag} */,
  {32'hbec4c908, 32'hbe90ede7} /* (1, 19, 26) {real, imag} */,
  {32'hbde18e2d, 32'hbe1dbc97} /* (1, 19, 25) {real, imag} */,
  {32'h3c32db10, 32'h3f0073a7} /* (1, 19, 24) {real, imag} */,
  {32'h3daae28d, 32'hbee20a86} /* (1, 19, 23) {real, imag} */,
  {32'hbe28e52d, 32'h3c09a218} /* (1, 19, 22) {real, imag} */,
  {32'h3ec1f3f6, 32'hbee3ccfa} /* (1, 19, 21) {real, imag} */,
  {32'h3c17a974, 32'hbd552c1f} /* (1, 19, 20) {real, imag} */,
  {32'h3e2bd1b6, 32'h3e5b6b62} /* (1, 19, 19) {real, imag} */,
  {32'hbd95c139, 32'h3df400e2} /* (1, 19, 18) {real, imag} */,
  {32'hbe9ac91c, 32'h3e81b6fa} /* (1, 19, 17) {real, imag} */,
  {32'h3ebecef7, 32'h3e54aed0} /* (1, 19, 16) {real, imag} */,
  {32'h3deb8420, 32'h3dfba3c8} /* (1, 19, 15) {real, imag} */,
  {32'hbe8aedc6, 32'h3e1f5051} /* (1, 19, 14) {real, imag} */,
  {32'hbdfc8c1a, 32'h3ec20d1a} /* (1, 19, 13) {real, imag} */,
  {32'hbeb6a9cb, 32'hbd7b5eb0} /* (1, 19, 12) {real, imag} */,
  {32'hbe904d76, 32'hbec74363} /* (1, 19, 11) {real, imag} */,
  {32'hbddcff03, 32'hbebd1363} /* (1, 19, 10) {real, imag} */,
  {32'h3d9c4b86, 32'h3e9dd876} /* (1, 19, 9) {real, imag} */,
  {32'h3e7b1dbe, 32'hbeabd69a} /* (1, 19, 8) {real, imag} */,
  {32'hbdb2b49e, 32'hbebfe009} /* (1, 19, 7) {real, imag} */,
  {32'hbd2948a0, 32'h3f0028ad} /* (1, 19, 6) {real, imag} */,
  {32'h3d5bf183, 32'h3b9e4700} /* (1, 19, 5) {real, imag} */,
  {32'h3ef6cac0, 32'hbdbae56e} /* (1, 19, 4) {real, imag} */,
  {32'h3e227013, 32'hbd8257f2} /* (1, 19, 3) {real, imag} */,
  {32'hbe67591d, 32'hbe015fc4} /* (1, 19, 2) {real, imag} */,
  {32'h3e86d454, 32'h3f0d5f76} /* (1, 19, 1) {real, imag} */,
  {32'h3ea99211, 32'h3e150007} /* (1, 19, 0) {real, imag} */,
  {32'hbf0f97df, 32'h3e667e3d} /* (1, 18, 31) {real, imag} */,
  {32'hbee690a8, 32'h3e2e223c} /* (1, 18, 30) {real, imag} */,
  {32'h3b472880, 32'hbccb7c58} /* (1, 18, 29) {real, imag} */,
  {32'hbe1df35c, 32'h3e28c910} /* (1, 18, 28) {real, imag} */,
  {32'hbdf86e2a, 32'hbedb119c} /* (1, 18, 27) {real, imag} */,
  {32'h3e65c6d6, 32'hbe52d583} /* (1, 18, 26) {real, imag} */,
  {32'hbdb5ac44, 32'h3e9ee528} /* (1, 18, 25) {real, imag} */,
  {32'h3d70232d, 32'h3da566aa} /* (1, 18, 24) {real, imag} */,
  {32'hbe58c643, 32'h3e10ac9e} /* (1, 18, 23) {real, imag} */,
  {32'h3d20aed8, 32'hbe2b6368} /* (1, 18, 22) {real, imag} */,
  {32'hbd219912, 32'h3ea4a12c} /* (1, 18, 21) {real, imag} */,
  {32'h3e300b71, 32'hbed25cce} /* (1, 18, 20) {real, imag} */,
  {32'hbe944026, 32'hbec31138} /* (1, 18, 19) {real, imag} */,
  {32'hbdf65832, 32'hbdb9e6c6} /* (1, 18, 18) {real, imag} */,
  {32'h3e14daf7, 32'hbdbbc36c} /* (1, 18, 17) {real, imag} */,
  {32'h3dba4766, 32'hbea0ffc0} /* (1, 18, 16) {real, imag} */,
  {32'hbb8951c0, 32'hbeadf99c} /* (1, 18, 15) {real, imag} */,
  {32'h3e2a6b18, 32'h3e12061e} /* (1, 18, 14) {real, imag} */,
  {32'h3f1f58e6, 32'h3d4ba22c} /* (1, 18, 13) {real, imag} */,
  {32'h3ef32082, 32'h3e72a4eb} /* (1, 18, 12) {real, imag} */,
  {32'h3e16d8f8, 32'hbf1a86a9} /* (1, 18, 11) {real, imag} */,
  {32'hbcf54428, 32'h3ecbf014} /* (1, 18, 10) {real, imag} */,
  {32'h3d155c7a, 32'h3e10c694} /* (1, 18, 9) {real, imag} */,
  {32'h3e1ac114, 32'h3ed3aa40} /* (1, 18, 8) {real, imag} */,
  {32'h3bc006b8, 32'hbc147c20} /* (1, 18, 7) {real, imag} */,
  {32'h3e32eef9, 32'h3eb5b28e} /* (1, 18, 6) {real, imag} */,
  {32'hbecb91d7, 32'hbda5fd93} /* (1, 18, 5) {real, imag} */,
  {32'hbd4ecebc, 32'hbe916f43} /* (1, 18, 4) {real, imag} */,
  {32'h3eb18c83, 32'h3dd98260} /* (1, 18, 3) {real, imag} */,
  {32'hbef8c550, 32'h3dab7dfa} /* (1, 18, 2) {real, imag} */,
  {32'hbe0c637c, 32'hbc936354} /* (1, 18, 1) {real, imag} */,
  {32'hbe9e9437, 32'hbd859c86} /* (1, 18, 0) {real, imag} */,
  {32'h3dc129f3, 32'h3e09e56e} /* (1, 17, 31) {real, imag} */,
  {32'h3dfb83ca, 32'h3e2d8ce6} /* (1, 17, 30) {real, imag} */,
  {32'hbe5283ff, 32'hbe269da9} /* (1, 17, 29) {real, imag} */,
  {32'hbda634c0, 32'hbe07a5ed} /* (1, 17, 28) {real, imag} */,
  {32'hbea27820, 32'hbe0823f7} /* (1, 17, 27) {real, imag} */,
  {32'hbe5db638, 32'hbe8bf850} /* (1, 17, 26) {real, imag} */,
  {32'h3e70b512, 32'hbe2ba8cb} /* (1, 17, 25) {real, imag} */,
  {32'hbec9de7b, 32'h3f01a7f1} /* (1, 17, 24) {real, imag} */,
  {32'h3d87361d, 32'h3e9afada} /* (1, 17, 23) {real, imag} */,
  {32'hbece02ef, 32'hbd016590} /* (1, 17, 22) {real, imag} */,
  {32'h3db17e18, 32'hbe2044e7} /* (1, 17, 21) {real, imag} */,
  {32'hbdd81d0c, 32'hbe73f267} /* (1, 17, 20) {real, imag} */,
  {32'h3e24b0fe, 32'h3ddede74} /* (1, 17, 19) {real, imag} */,
  {32'hbe6cbc98, 32'hbe06c5cd} /* (1, 17, 18) {real, imag} */,
  {32'h3e98434c, 32'hbea2723f} /* (1, 17, 17) {real, imag} */,
  {32'hbe5df71c, 32'hbe9930ad} /* (1, 17, 16) {real, imag} */,
  {32'hbd1440e4, 32'h3e00c11c} /* (1, 17, 15) {real, imag} */,
  {32'hbec5c9b6, 32'h3dfa9cce} /* (1, 17, 14) {real, imag} */,
  {32'hbeb06334, 32'h3d8f6439} /* (1, 17, 13) {real, imag} */,
  {32'h3e0308a0, 32'h3d8c5857} /* (1, 17, 12) {real, imag} */,
  {32'hbcd30078, 32'hbe0231cf} /* (1, 17, 11) {real, imag} */,
  {32'hbdbec784, 32'hbe99aece} /* (1, 17, 10) {real, imag} */,
  {32'h3d8d98cc, 32'h3d4e759c} /* (1, 17, 9) {real, imag} */,
  {32'h3e085084, 32'h3e98e121} /* (1, 17, 8) {real, imag} */,
  {32'h3e87e19e, 32'hbe80fbdb} /* (1, 17, 7) {real, imag} */,
  {32'hbcab1038, 32'h3bc2db98} /* (1, 17, 6) {real, imag} */,
  {32'hbd952254, 32'h3e976b9a} /* (1, 17, 5) {real, imag} */,
  {32'hbcae7550, 32'h3e685883} /* (1, 17, 4) {real, imag} */,
  {32'hbef4daee, 32'h3c0dada0} /* (1, 17, 3) {real, imag} */,
  {32'hbea56c5c, 32'hbe04fd1c} /* (1, 17, 2) {real, imag} */,
  {32'h3e4666a1, 32'h3e14f99a} /* (1, 17, 1) {real, imag} */,
  {32'hbd4f956a, 32'hbea610be} /* (1, 17, 0) {real, imag} */,
  {32'h3df4f4c2, 32'hbd5ca2f2} /* (1, 16, 31) {real, imag} */,
  {32'hbe465f0b, 32'h3e249a73} /* (1, 16, 30) {real, imag} */,
  {32'h3d85a698, 32'hbdb3b368} /* (1, 16, 29) {real, imag} */,
  {32'hbba5c220, 32'hbe908f80} /* (1, 16, 28) {real, imag} */,
  {32'hbed7f5c4, 32'hbedd6793} /* (1, 16, 27) {real, imag} */,
  {32'hbd54d36c, 32'h3e1957e2} /* (1, 16, 26) {real, imag} */,
  {32'hbe93012e, 32'hbdfb8668} /* (1, 16, 25) {real, imag} */,
  {32'h3e6ca209, 32'h3dd1bad0} /* (1, 16, 24) {real, imag} */,
  {32'hbed2891f, 32'hbd5ef902} /* (1, 16, 23) {real, imag} */,
  {32'h3dfbf7f8, 32'h3ed1d192} /* (1, 16, 22) {real, imag} */,
  {32'hbea19b42, 32'hbd8f6abe} /* (1, 16, 21) {real, imag} */,
  {32'hbe3b12d1, 32'h3d828016} /* (1, 16, 20) {real, imag} */,
  {32'hbd58a67a, 32'hbd8fd57f} /* (1, 16, 19) {real, imag} */,
  {32'h3e8d3d59, 32'h3de69eae} /* (1, 16, 18) {real, imag} */,
  {32'hbdca72b2, 32'h3d897635} /* (1, 16, 17) {real, imag} */,
  {32'h3f182cc1, 32'h00000000} /* (1, 16, 16) {real, imag} */,
  {32'hbdca72b2, 32'hbd897635} /* (1, 16, 15) {real, imag} */,
  {32'h3e8d3d59, 32'hbde69eae} /* (1, 16, 14) {real, imag} */,
  {32'hbd58a67a, 32'h3d8fd57f} /* (1, 16, 13) {real, imag} */,
  {32'hbe3b12d1, 32'hbd828016} /* (1, 16, 12) {real, imag} */,
  {32'hbea19b42, 32'h3d8f6abe} /* (1, 16, 11) {real, imag} */,
  {32'h3dfbf7f8, 32'hbed1d192} /* (1, 16, 10) {real, imag} */,
  {32'hbed2891f, 32'h3d5ef902} /* (1, 16, 9) {real, imag} */,
  {32'h3e6ca209, 32'hbdd1bad0} /* (1, 16, 8) {real, imag} */,
  {32'hbe93012e, 32'h3dfb8668} /* (1, 16, 7) {real, imag} */,
  {32'hbd54d36c, 32'hbe1957e2} /* (1, 16, 6) {real, imag} */,
  {32'hbed7f5c4, 32'h3edd6793} /* (1, 16, 5) {real, imag} */,
  {32'hbba5c220, 32'h3e908f80} /* (1, 16, 4) {real, imag} */,
  {32'h3d85a698, 32'h3db3b368} /* (1, 16, 3) {real, imag} */,
  {32'hbe465f0b, 32'hbe249a73} /* (1, 16, 2) {real, imag} */,
  {32'h3df4f4c2, 32'h3d5ca2f2} /* (1, 16, 1) {real, imag} */,
  {32'h3da0d4a0, 32'h00000000} /* (1, 16, 0) {real, imag} */,
  {32'h3e4666a1, 32'hbe14f99a} /* (1, 15, 31) {real, imag} */,
  {32'hbea56c5c, 32'h3e04fd1c} /* (1, 15, 30) {real, imag} */,
  {32'hbef4daee, 32'hbc0dada0} /* (1, 15, 29) {real, imag} */,
  {32'hbcae7550, 32'hbe685883} /* (1, 15, 28) {real, imag} */,
  {32'hbd952254, 32'hbe976b9a} /* (1, 15, 27) {real, imag} */,
  {32'hbcab1038, 32'hbbc2db98} /* (1, 15, 26) {real, imag} */,
  {32'h3e87e19e, 32'h3e80fbdb} /* (1, 15, 25) {real, imag} */,
  {32'h3e085084, 32'hbe98e121} /* (1, 15, 24) {real, imag} */,
  {32'h3d8d98cc, 32'hbd4e759c} /* (1, 15, 23) {real, imag} */,
  {32'hbdbec784, 32'h3e99aece} /* (1, 15, 22) {real, imag} */,
  {32'hbcd30078, 32'h3e0231cf} /* (1, 15, 21) {real, imag} */,
  {32'h3e0308a0, 32'hbd8c5857} /* (1, 15, 20) {real, imag} */,
  {32'hbeb06334, 32'hbd8f6439} /* (1, 15, 19) {real, imag} */,
  {32'hbec5c9b6, 32'hbdfa9cce} /* (1, 15, 18) {real, imag} */,
  {32'hbd1440e4, 32'hbe00c11c} /* (1, 15, 17) {real, imag} */,
  {32'hbe5df71c, 32'h3e9930ad} /* (1, 15, 16) {real, imag} */,
  {32'h3e98434c, 32'h3ea2723f} /* (1, 15, 15) {real, imag} */,
  {32'hbe6cbc98, 32'h3e06c5cd} /* (1, 15, 14) {real, imag} */,
  {32'h3e24b0fe, 32'hbddede74} /* (1, 15, 13) {real, imag} */,
  {32'hbdd81d0c, 32'h3e73f267} /* (1, 15, 12) {real, imag} */,
  {32'h3db17e18, 32'h3e2044e7} /* (1, 15, 11) {real, imag} */,
  {32'hbece02ef, 32'h3d016590} /* (1, 15, 10) {real, imag} */,
  {32'h3d87361d, 32'hbe9afada} /* (1, 15, 9) {real, imag} */,
  {32'hbec9de7b, 32'hbf01a7f1} /* (1, 15, 8) {real, imag} */,
  {32'h3e70b512, 32'h3e2ba8cb} /* (1, 15, 7) {real, imag} */,
  {32'hbe5db638, 32'h3e8bf850} /* (1, 15, 6) {real, imag} */,
  {32'hbea27820, 32'h3e0823f7} /* (1, 15, 5) {real, imag} */,
  {32'hbda634c0, 32'h3e07a5ed} /* (1, 15, 4) {real, imag} */,
  {32'hbe5283ff, 32'h3e269da9} /* (1, 15, 3) {real, imag} */,
  {32'h3dfb83ca, 32'hbe2d8ce6} /* (1, 15, 2) {real, imag} */,
  {32'h3dc129f3, 32'hbe09e56e} /* (1, 15, 1) {real, imag} */,
  {32'hbd4f956a, 32'h3ea610be} /* (1, 15, 0) {real, imag} */,
  {32'hbe0c637c, 32'h3c936354} /* (1, 14, 31) {real, imag} */,
  {32'hbef8c550, 32'hbdab7dfa} /* (1, 14, 30) {real, imag} */,
  {32'h3eb18c83, 32'hbdd98260} /* (1, 14, 29) {real, imag} */,
  {32'hbd4ecebc, 32'h3e916f43} /* (1, 14, 28) {real, imag} */,
  {32'hbecb91d7, 32'h3da5fd93} /* (1, 14, 27) {real, imag} */,
  {32'h3e32eef9, 32'hbeb5b28e} /* (1, 14, 26) {real, imag} */,
  {32'h3bc006b8, 32'h3c147c20} /* (1, 14, 25) {real, imag} */,
  {32'h3e1ac114, 32'hbed3aa40} /* (1, 14, 24) {real, imag} */,
  {32'h3d155c7a, 32'hbe10c694} /* (1, 14, 23) {real, imag} */,
  {32'hbcf54428, 32'hbecbf014} /* (1, 14, 22) {real, imag} */,
  {32'h3e16d8f8, 32'h3f1a86a9} /* (1, 14, 21) {real, imag} */,
  {32'h3ef32082, 32'hbe72a4eb} /* (1, 14, 20) {real, imag} */,
  {32'h3f1f58e6, 32'hbd4ba22c} /* (1, 14, 19) {real, imag} */,
  {32'h3e2a6b18, 32'hbe12061e} /* (1, 14, 18) {real, imag} */,
  {32'hbb8951c0, 32'h3eadf99c} /* (1, 14, 17) {real, imag} */,
  {32'h3dba4766, 32'h3ea0ffc0} /* (1, 14, 16) {real, imag} */,
  {32'h3e14daf7, 32'h3dbbc36c} /* (1, 14, 15) {real, imag} */,
  {32'hbdf65832, 32'h3db9e6c6} /* (1, 14, 14) {real, imag} */,
  {32'hbe944026, 32'h3ec31138} /* (1, 14, 13) {real, imag} */,
  {32'h3e300b71, 32'h3ed25cce} /* (1, 14, 12) {real, imag} */,
  {32'hbd219912, 32'hbea4a12c} /* (1, 14, 11) {real, imag} */,
  {32'h3d20aed8, 32'h3e2b6368} /* (1, 14, 10) {real, imag} */,
  {32'hbe58c643, 32'hbe10ac9e} /* (1, 14, 9) {real, imag} */,
  {32'h3d70232d, 32'hbda566aa} /* (1, 14, 8) {real, imag} */,
  {32'hbdb5ac44, 32'hbe9ee528} /* (1, 14, 7) {real, imag} */,
  {32'h3e65c6d6, 32'h3e52d583} /* (1, 14, 6) {real, imag} */,
  {32'hbdf86e2a, 32'h3edb119c} /* (1, 14, 5) {real, imag} */,
  {32'hbe1df35c, 32'hbe28c910} /* (1, 14, 4) {real, imag} */,
  {32'h3b472880, 32'h3ccb7c58} /* (1, 14, 3) {real, imag} */,
  {32'hbee690a8, 32'hbe2e223c} /* (1, 14, 2) {real, imag} */,
  {32'hbf0f97df, 32'hbe667e3d} /* (1, 14, 1) {real, imag} */,
  {32'hbe9e9437, 32'h3d859c86} /* (1, 14, 0) {real, imag} */,
  {32'h3e86d454, 32'hbf0d5f76} /* (1, 13, 31) {real, imag} */,
  {32'hbe67591d, 32'h3e015fc4} /* (1, 13, 30) {real, imag} */,
  {32'h3e227013, 32'h3d8257f2} /* (1, 13, 29) {real, imag} */,
  {32'h3ef6cac0, 32'h3dbae56e} /* (1, 13, 28) {real, imag} */,
  {32'h3d5bf183, 32'hbb9e4700} /* (1, 13, 27) {real, imag} */,
  {32'hbd2948a0, 32'hbf0028ad} /* (1, 13, 26) {real, imag} */,
  {32'hbdb2b49e, 32'h3ebfe009} /* (1, 13, 25) {real, imag} */,
  {32'h3e7b1dbe, 32'h3eabd69a} /* (1, 13, 24) {real, imag} */,
  {32'h3d9c4b86, 32'hbe9dd876} /* (1, 13, 23) {real, imag} */,
  {32'hbddcff03, 32'h3ebd1363} /* (1, 13, 22) {real, imag} */,
  {32'hbe904d76, 32'h3ec74363} /* (1, 13, 21) {real, imag} */,
  {32'hbeb6a9cb, 32'h3d7b5eb0} /* (1, 13, 20) {real, imag} */,
  {32'hbdfc8c1a, 32'hbec20d1a} /* (1, 13, 19) {real, imag} */,
  {32'hbe8aedc6, 32'hbe1f5051} /* (1, 13, 18) {real, imag} */,
  {32'h3deb8420, 32'hbdfba3c8} /* (1, 13, 17) {real, imag} */,
  {32'h3ebecef7, 32'hbe54aed0} /* (1, 13, 16) {real, imag} */,
  {32'hbe9ac91c, 32'hbe81b6fa} /* (1, 13, 15) {real, imag} */,
  {32'hbd95c139, 32'hbdf400e2} /* (1, 13, 14) {real, imag} */,
  {32'h3e2bd1b6, 32'hbe5b6b62} /* (1, 13, 13) {real, imag} */,
  {32'h3c17a974, 32'h3d552c1f} /* (1, 13, 12) {real, imag} */,
  {32'h3ec1f3f6, 32'h3ee3ccfa} /* (1, 13, 11) {real, imag} */,
  {32'hbe28e52d, 32'hbc09a218} /* (1, 13, 10) {real, imag} */,
  {32'h3daae28d, 32'h3ee20a86} /* (1, 13, 9) {real, imag} */,
  {32'h3c32db10, 32'hbf0073a7} /* (1, 13, 8) {real, imag} */,
  {32'hbde18e2d, 32'h3e1dbc97} /* (1, 13, 7) {real, imag} */,
  {32'hbec4c908, 32'h3e90ede7} /* (1, 13, 6) {real, imag} */,
  {32'hbe6af962, 32'h3ebe858a} /* (1, 13, 5) {real, imag} */,
  {32'hbf052c0b, 32'h3d591d9e} /* (1, 13, 4) {real, imag} */,
  {32'h3d635e22, 32'hbe30e12a} /* (1, 13, 3) {real, imag} */,
  {32'h3e3ecfec, 32'hbd8ac2fe} /* (1, 13, 2) {real, imag} */,
  {32'hbda56825, 32'hbec57fcc} /* (1, 13, 1) {real, imag} */,
  {32'h3ea99211, 32'hbe150007} /* (1, 13, 0) {real, imag} */,
  {32'h3d92b59a, 32'hbe94729c} /* (1, 12, 31) {real, imag} */,
  {32'h3eb45048, 32'hbe8616d7} /* (1, 12, 30) {real, imag} */,
  {32'hbdf79448, 32'hbec215a5} /* (1, 12, 29) {real, imag} */,
  {32'hbe62cd9b, 32'h3e40ab02} /* (1, 12, 28) {real, imag} */,
  {32'h3e86f25d, 32'h3f0b4dc0} /* (1, 12, 27) {real, imag} */,
  {32'hbd5d55ae, 32'hbf0abd73} /* (1, 12, 26) {real, imag} */,
  {32'h3d780acc, 32'h3cc45540} /* (1, 12, 25) {real, imag} */,
  {32'hbb8c2fb0, 32'h3d7305ec} /* (1, 12, 24) {real, imag} */,
  {32'h3e953e57, 32'h3ef73b13} /* (1, 12, 23) {real, imag} */,
  {32'h3ec28a1a, 32'h3f2a89dc} /* (1, 12, 22) {real, imag} */,
  {32'hbe98bac0, 32'h3f298280} /* (1, 12, 21) {real, imag} */,
  {32'h3eb542f0, 32'h3f035dbf} /* (1, 12, 20) {real, imag} */,
  {32'h3e231b11, 32'h3e3d6a6e} /* (1, 12, 19) {real, imag} */,
  {32'h3d0aa540, 32'h3e1df7e2} /* (1, 12, 18) {real, imag} */,
  {32'hbe5c62fa, 32'h3e7995c8} /* (1, 12, 17) {real, imag} */,
  {32'hbe7647b9, 32'hbec6b940} /* (1, 12, 16) {real, imag} */,
  {32'h3dcc12c5, 32'h3df38f18} /* (1, 12, 15) {real, imag} */,
  {32'h3dbc29ca, 32'h3eb17393} /* (1, 12, 14) {real, imag} */,
  {32'hbe26bb34, 32'h3d7504d3} /* (1, 12, 13) {real, imag} */,
  {32'hbeb4c4c5, 32'h3e28c624} /* (1, 12, 12) {real, imag} */,
  {32'h3da01b1c, 32'h3e59f333} /* (1, 12, 11) {real, imag} */,
  {32'hbe8c87b4, 32'hbf0a885e} /* (1, 12, 10) {real, imag} */,
  {32'hbd5d60de, 32'h3f007a08} /* (1, 12, 9) {real, imag} */,
  {32'h3ee6a2ab, 32'hbe2997a6} /* (1, 12, 8) {real, imag} */,
  {32'hbf05950c, 32'h3eb5006d} /* (1, 12, 7) {real, imag} */,
  {32'h3e9ea700, 32'h3d259c4c} /* (1, 12, 6) {real, imag} */,
  {32'h3ed4e110, 32'hbabb1200} /* (1, 12, 5) {real, imag} */,
  {32'h3ea7c00e, 32'hbe9d6d54} /* (1, 12, 4) {real, imag} */,
  {32'hbe5596ab, 32'hbde06392} /* (1, 12, 3) {real, imag} */,
  {32'h3da84aac, 32'hbe340a9f} /* (1, 12, 2) {real, imag} */,
  {32'h3edafe84, 32'hbd278650} /* (1, 12, 1) {real, imag} */,
  {32'hbcf62a40, 32'hbecad71e} /* (1, 12, 0) {real, imag} */,
  {32'h3efd130a, 32'h3ee8a13c} /* (1, 11, 31) {real, imag} */,
  {32'h3d891694, 32'hbf82ebab} /* (1, 11, 30) {real, imag} */,
  {32'hbea9e59b, 32'h3dbd3033} /* (1, 11, 29) {real, imag} */,
  {32'h3deb047d, 32'h3dceeba6} /* (1, 11, 28) {real, imag} */,
  {32'h3d20cf58, 32'hbea62851} /* (1, 11, 27) {real, imag} */,
  {32'h3ee688b1, 32'h3e3b41a2} /* (1, 11, 26) {real, imag} */,
  {32'hbe594781, 32'h3e2d65be} /* (1, 11, 25) {real, imag} */,
  {32'h3d9c4ec0, 32'hbd4a48ec} /* (1, 11, 24) {real, imag} */,
  {32'h3f20f686, 32'hbf64d2bc} /* (1, 11, 23) {real, imag} */,
  {32'h3df4b7d0, 32'h3ecb9166} /* (1, 11, 22) {real, imag} */,
  {32'h3e3f6a4e, 32'hbd9f6de8} /* (1, 11, 21) {real, imag} */,
  {32'hbf3f550b, 32'h3f1f608a} /* (1, 11, 20) {real, imag} */,
  {32'hbe11bad0, 32'hbeefd6a0} /* (1, 11, 19) {real, imag} */,
  {32'hbdf1b51a, 32'h3d439730} /* (1, 11, 18) {real, imag} */,
  {32'h3ea69198, 32'h3d5c752e} /* (1, 11, 17) {real, imag} */,
  {32'h3e89c370, 32'h3da20bdc} /* (1, 11, 16) {real, imag} */,
  {32'hbe082d6a, 32'h3d3e56e0} /* (1, 11, 15) {real, imag} */,
  {32'hbe1e9db6, 32'h3e3ef119} /* (1, 11, 14) {real, imag} */,
  {32'h3e369232, 32'hbdff284b} /* (1, 11, 13) {real, imag} */,
  {32'hbe089dd6, 32'h3dadd05c} /* (1, 11, 12) {real, imag} */,
  {32'hbf55a5ba, 32'hbed70f54} /* (1, 11, 11) {real, imag} */,
  {32'hbf21cfdc, 32'hbe25002c} /* (1, 11, 10) {real, imag} */,
  {32'hbe3ab9c7, 32'hbe992834} /* (1, 11, 9) {real, imag} */,
  {32'hbe125c6d, 32'h3e5715ce} /* (1, 11, 8) {real, imag} */,
  {32'hbdb74810, 32'hbed55ec7} /* (1, 11, 7) {real, imag} */,
  {32'h3eb61936, 32'hbe4d924a} /* (1, 11, 6) {real, imag} */,
  {32'hbf04e76e, 32'hbdd4e9f2} /* (1, 11, 5) {real, imag} */,
  {32'h3e2159ee, 32'hbead5863} /* (1, 11, 4) {real, imag} */,
  {32'hbe7573c7, 32'hbe654a0e} /* (1, 11, 3) {real, imag} */,
  {32'h3c238630, 32'hbe87bf42} /* (1, 11, 2) {real, imag} */,
  {32'h3e96c5a9, 32'h3f4648ba} /* (1, 11, 1) {real, imag} */,
  {32'h3e86cab6, 32'h3bc904c0} /* (1, 11, 0) {real, imag} */,
  {32'hbe216149, 32'hbf0bf583} /* (1, 10, 31) {real, imag} */,
  {32'hbe442deb, 32'h3f0f3aab} /* (1, 10, 30) {real, imag} */,
  {32'hbec099ad, 32'hbd0339dc} /* (1, 10, 29) {real, imag} */,
  {32'hbe18bc94, 32'hbf3ffd7a} /* (1, 10, 28) {real, imag} */,
  {32'hbe5a165a, 32'h3e301014} /* (1, 10, 27) {real, imag} */,
  {32'hbdec8cce, 32'h3decba56} /* (1, 10, 26) {real, imag} */,
  {32'hbee56ea3, 32'h3bf80170} /* (1, 10, 25) {real, imag} */,
  {32'h3f138efc, 32'h3ef740eb} /* (1, 10, 24) {real, imag} */,
  {32'h3e319b6c, 32'hbe8c05bb} /* (1, 10, 23) {real, imag} */,
  {32'h3db7e58a, 32'h3e870906} /* (1, 10, 22) {real, imag} */,
  {32'hbf2299eb, 32'h3d6abe00} /* (1, 10, 21) {real, imag} */,
  {32'hbded2d71, 32'hbe92f8aa} /* (1, 10, 20) {real, imag} */,
  {32'h3e94d66d, 32'h3e5c6843} /* (1, 10, 19) {real, imag} */,
  {32'h3bc0de80, 32'hbbd88c80} /* (1, 10, 18) {real, imag} */,
  {32'h3e41586e, 32'hbd2b7cf1} /* (1, 10, 17) {real, imag} */,
  {32'h3c739c9c, 32'h3be57490} /* (1, 10, 16) {real, imag} */,
  {32'hbd6fd5d6, 32'h3e569edb} /* (1, 10, 15) {real, imag} */,
  {32'hbe8a1818, 32'hbeb61ec6} /* (1, 10, 14) {real, imag} */,
  {32'h3e47dd2e, 32'h3e2fccbd} /* (1, 10, 13) {real, imag} */,
  {32'hbef039fe, 32'hbd673fb8} /* (1, 10, 12) {real, imag} */,
  {32'hbd974a9a, 32'h3e92cf26} /* (1, 10, 11) {real, imag} */,
  {32'h3e66bda4, 32'hbcb19d40} /* (1, 10, 10) {real, imag} */,
  {32'h3f5539bd, 32'h3d419654} /* (1, 10, 9) {real, imag} */,
  {32'hbe86cf96, 32'hbde35627} /* (1, 10, 8) {real, imag} */,
  {32'h3e9007c5, 32'h3d577bb0} /* (1, 10, 7) {real, imag} */,
  {32'hbd4c6432, 32'hbeacfd34} /* (1, 10, 6) {real, imag} */,
  {32'hbeb70d5d, 32'hbe3b5a28} /* (1, 10, 5) {real, imag} */,
  {32'h3eb88261, 32'h3d9e7290} /* (1, 10, 4) {real, imag} */,
  {32'h3f2beed9, 32'hbdf4c832} /* (1, 10, 3) {real, imag} */,
  {32'h3f05fbdb, 32'h3f409c35} /* (1, 10, 2) {real, imag} */,
  {32'h3ea4812f, 32'hbe220dbf} /* (1, 10, 1) {real, imag} */,
  {32'hbe16715b, 32'hbdf40b1b} /* (1, 10, 0) {real, imag} */,
  {32'h3de2b852, 32'hbd913358} /* (1, 9, 31) {real, imag} */,
  {32'h3ea44570, 32'h3f3205d8} /* (1, 9, 30) {real, imag} */,
  {32'hbf1aaf46, 32'hbee3bcd9} /* (1, 9, 29) {real, imag} */,
  {32'hbe0fa4fa, 32'hbedb21b0} /* (1, 9, 28) {real, imag} */,
  {32'hbe88f268, 32'hbd6878b4} /* (1, 9, 27) {real, imag} */,
  {32'h3eb5482e, 32'hbee84416} /* (1, 9, 26) {real, imag} */,
  {32'hbea9d2a1, 32'h3db3779c} /* (1, 9, 25) {real, imag} */,
  {32'hbd69bc28, 32'hbe9b5c50} /* (1, 9, 24) {real, imag} */,
  {32'h3e16b32a, 32'hbe727178} /* (1, 9, 23) {real, imag} */,
  {32'h3cf499f0, 32'h3ea83ca4} /* (1, 9, 22) {real, imag} */,
  {32'h3e059c0c, 32'hbbd5aaf0} /* (1, 9, 21) {real, imag} */,
  {32'h3dbbc618, 32'hbf3530d8} /* (1, 9, 20) {real, imag} */,
  {32'hbe5e9e70, 32'h3deec3e7} /* (1, 9, 19) {real, imag} */,
  {32'h3f3e3707, 32'h3e75d65e} /* (1, 9, 18) {real, imag} */,
  {32'h3ea02ca9, 32'hbe4af2c9} /* (1, 9, 17) {real, imag} */,
  {32'h3eb7ba78, 32'h3efe5414} /* (1, 9, 16) {real, imag} */,
  {32'hbe3abfc1, 32'hbdc43745} /* (1, 9, 15) {real, imag} */,
  {32'hbe871240, 32'hbf54cd14} /* (1, 9, 14) {real, imag} */,
  {32'h3e8361fd, 32'h3eb7fa8a} /* (1, 9, 13) {real, imag} */,
  {32'h3e277d6e, 32'hbe39f892} /* (1, 9, 12) {real, imag} */,
  {32'hbf08f3f8, 32'hbe5abfc4} /* (1, 9, 11) {real, imag} */,
  {32'hbe725d7b, 32'hbc3173b0} /* (1, 9, 10) {real, imag} */,
  {32'h3ea3a31c, 32'hbc9b3600} /* (1, 9, 9) {real, imag} */,
  {32'hbdebf525, 32'h3d6850dc} /* (1, 9, 8) {real, imag} */,
  {32'hbde6a554, 32'h3db3650c} /* (1, 9, 7) {real, imag} */,
  {32'hbe6ab588, 32'hbeaf42f8} /* (1, 9, 6) {real, imag} */,
  {32'hbcf27446, 32'h3d02ba00} /* (1, 9, 5) {real, imag} */,
  {32'h3ed68702, 32'hbec87c8b} /* (1, 9, 4) {real, imag} */,
  {32'hbebb5cc7, 32'h3ed64c92} /* (1, 9, 3) {real, imag} */,
  {32'h3ec125ce, 32'h3ed3bd05} /* (1, 9, 2) {real, imag} */,
  {32'hbe8e552b, 32'hbdb52514} /* (1, 9, 1) {real, imag} */,
  {32'hbf0a8538, 32'hbe12a964} /* (1, 9, 0) {real, imag} */,
  {32'h3f711a69, 32'h3ee74c57} /* (1, 8, 31) {real, imag} */,
  {32'hbfd29dcf, 32'h3e4b78a6} /* (1, 8, 30) {real, imag} */,
  {32'hbdc4f1d9, 32'hbe1179f8} /* (1, 8, 29) {real, imag} */,
  {32'hbe086cff, 32'h3e45847c} /* (1, 8, 28) {real, imag} */,
  {32'hbd4df8dc, 32'h3e8ff2a9} /* (1, 8, 27) {real, imag} */,
  {32'hbdad3904, 32'h3ed929c0} /* (1, 8, 26) {real, imag} */,
  {32'h3f8aba94, 32'h3dfd6eb3} /* (1, 8, 25) {real, imag} */,
  {32'hbe3b3142, 32'h3f2aee09} /* (1, 8, 24) {real, imag} */,
  {32'h3f4b5f18, 32'h3e1d946a} /* (1, 8, 23) {real, imag} */,
  {32'hbf06bce8, 32'hbec06f47} /* (1, 8, 22) {real, imag} */,
  {32'hbd768dac, 32'h3df1b8b4} /* (1, 8, 21) {real, imag} */,
  {32'hbede279d, 32'h3eb590d4} /* (1, 8, 20) {real, imag} */,
  {32'hbe6085cb, 32'hbf17b956} /* (1, 8, 19) {real, imag} */,
  {32'h3e0cc3fa, 32'h3e20d0de} /* (1, 8, 18) {real, imag} */,
  {32'h3e1d2dd6, 32'h3d424678} /* (1, 8, 17) {real, imag} */,
  {32'hbeac6ca6, 32'h3c416e00} /* (1, 8, 16) {real, imag} */,
  {32'h3e960138, 32'h3d13f65a} /* (1, 8, 15) {real, imag} */,
  {32'h3e3cf9d0, 32'hbe3dc29b} /* (1, 8, 14) {real, imag} */,
  {32'hbec76b29, 32'hbeff3d72} /* (1, 8, 13) {real, imag} */,
  {32'hbe1d7f00, 32'hbf0003a6} /* (1, 8, 12) {real, imag} */,
  {32'h3f1fb2e6, 32'hbe8c34c1} /* (1, 8, 11) {real, imag} */,
  {32'h3b716b40, 32'h3f4d9fa6} /* (1, 8, 10) {real, imag} */,
  {32'h3f0db74a, 32'h3ebae5c8} /* (1, 8, 9) {real, imag} */,
  {32'h3e16c6ec, 32'hbf0f1c30} /* (1, 8, 8) {real, imag} */,
  {32'h3d3b497f, 32'h3ead7771} /* (1, 8, 7) {real, imag} */,
  {32'hbe86b9b5, 32'hbe113d61} /* (1, 8, 6) {real, imag} */,
  {32'hba003180, 32'hbf99c8b8} /* (1, 8, 5) {real, imag} */,
  {32'hbedb42a8, 32'h3ef91a5c} /* (1, 8, 4) {real, imag} */,
  {32'hbd517810, 32'h3e700332} /* (1, 8, 3) {real, imag} */,
  {32'h3e613ea0, 32'h3d68a410} /* (1, 8, 2) {real, imag} */,
  {32'h3f1cd2fe, 32'h3f401539} /* (1, 8, 1) {real, imag} */,
  {32'h3ebd11e8, 32'h3f603a32} /* (1, 8, 0) {real, imag} */,
  {32'hbec03e15, 32'h3eac4c32} /* (1, 7, 31) {real, imag} */,
  {32'h3ea01c43, 32'hbe006194} /* (1, 7, 30) {real, imag} */,
  {32'hbd84dc1e, 32'hbe850fda} /* (1, 7, 29) {real, imag} */,
  {32'hbf18e080, 32'h3f71ff0b} /* (1, 7, 28) {real, imag} */,
  {32'h3e2cac73, 32'hbeca0fa9} /* (1, 7, 27) {real, imag} */,
  {32'h3ef3035a, 32'h3e218678} /* (1, 7, 26) {real, imag} */,
  {32'h3ed27864, 32'h3e2e0394} /* (1, 7, 25) {real, imag} */,
  {32'h3f0c6722, 32'hbf104206} /* (1, 7, 24) {real, imag} */,
  {32'hbe7f30e0, 32'h3f058c34} /* (1, 7, 23) {real, imag} */,
  {32'hbe2d12c5, 32'h3da14859} /* (1, 7, 22) {real, imag} */,
  {32'hbe8bd851, 32'h3ea4799c} /* (1, 7, 21) {real, imag} */,
  {32'h3daa86cc, 32'h3ed1c43b} /* (1, 7, 20) {real, imag} */,
  {32'h3c799620, 32'hbe1bcc8e} /* (1, 7, 19) {real, imag} */,
  {32'hbe3a4bcd, 32'h3d06f212} /* (1, 7, 18) {real, imag} */,
  {32'h3d791e88, 32'h3eaf13bb} /* (1, 7, 17) {real, imag} */,
  {32'h3d43da76, 32'h3e907443} /* (1, 7, 16) {real, imag} */,
  {32'h3e13ccde, 32'hbe49dbf3} /* (1, 7, 15) {real, imag} */,
  {32'h3e9d5ff9, 32'h3dc141d7} /* (1, 7, 14) {real, imag} */,
  {32'h3d0da13a, 32'h3ea7c5aa} /* (1, 7, 13) {real, imag} */,
  {32'hbe1b811c, 32'hbf16de2e} /* (1, 7, 12) {real, imag} */,
  {32'h3d22fd10, 32'h3eb0e3ca} /* (1, 7, 11) {real, imag} */,
  {32'h3c101f30, 32'h3efc68e1} /* (1, 7, 10) {real, imag} */,
  {32'h3f22f6a7, 32'h3e0d7394} /* (1, 7, 9) {real, imag} */,
  {32'h3e1f2ec5, 32'h3de935d6} /* (1, 7, 8) {real, imag} */,
  {32'hbec0ddf4, 32'h3e99bf2a} /* (1, 7, 7) {real, imag} */,
  {32'hbf139ba1, 32'h3f14fb68} /* (1, 7, 6) {real, imag} */,
  {32'hbc8f3640, 32'h3e9815ef} /* (1, 7, 5) {real, imag} */,
  {32'hbda17e03, 32'hbe0ebd06} /* (1, 7, 4) {real, imag} */,
  {32'hbd8dc441, 32'h3d85942c} /* (1, 7, 3) {real, imag} */,
  {32'hbf098137, 32'hbed01e73} /* (1, 7, 2) {real, imag} */,
  {32'h3f51151a, 32'hbf277e1e} /* (1, 7, 1) {real, imag} */,
  {32'h3e024878, 32'hbec38335} /* (1, 7, 0) {real, imag} */,
  {32'hbec4f184, 32'h3f9b40b0} /* (1, 6, 31) {real, imag} */,
  {32'hbf4789eb, 32'h3ea017b4} /* (1, 6, 30) {real, imag} */,
  {32'h3eb0fbe8, 32'hbe9f8ea8} /* (1, 6, 29) {real, imag} */,
  {32'hbeefda0e, 32'hbe61da77} /* (1, 6, 28) {real, imag} */,
  {32'h3f34d0f1, 32'hbf72a08a} /* (1, 6, 27) {real, imag} */,
  {32'h3ecbbdc4, 32'h3ec9a774} /* (1, 6, 26) {real, imag} */,
  {32'h3e43a154, 32'hbd421e1b} /* (1, 6, 25) {real, imag} */,
  {32'h3d6e86fe, 32'h3df2c71c} /* (1, 6, 24) {real, imag} */,
  {32'hbf0ffe2d, 32'h3f014d38} /* (1, 6, 23) {real, imag} */,
  {32'h3e03d81e, 32'hbe0a2866} /* (1, 6, 22) {real, imag} */,
  {32'hbed40b4a, 32'hbd0ce6bc} /* (1, 6, 21) {real, imag} */,
  {32'h3d8c5642, 32'hbd2782f4} /* (1, 6, 20) {real, imag} */,
  {32'h3d4664c8, 32'hbead85a8} /* (1, 6, 19) {real, imag} */,
  {32'h39760f00, 32'hbc5447c0} /* (1, 6, 18) {real, imag} */,
  {32'h3e285ce6, 32'hbe494e18} /* (1, 6, 17) {real, imag} */,
  {32'h3d872552, 32'hbd54d534} /* (1, 6, 16) {real, imag} */,
  {32'hbe872f8b, 32'hbddf33f3} /* (1, 6, 15) {real, imag} */,
  {32'hbd4c8d94, 32'h3de8828c} /* (1, 6, 14) {real, imag} */,
  {32'hbec98a73, 32'hbe5e144f} /* (1, 6, 13) {real, imag} */,
  {32'h3d704aa6, 32'h3c0ce738} /* (1, 6, 12) {real, imag} */,
  {32'hbe710ea5, 32'hbf171586} /* (1, 6, 11) {real, imag} */,
  {32'h3e556ef7, 32'hbe1f2bea} /* (1, 6, 10) {real, imag} */,
  {32'h3eb633a2, 32'h3f37881c} /* (1, 6, 9) {real, imag} */,
  {32'h3e4fa023, 32'hbe1d5f82} /* (1, 6, 8) {real, imag} */,
  {32'h3f0ed710, 32'hbee9b823} /* (1, 6, 7) {real, imag} */,
  {32'hbeaf52bc, 32'hbeaeacde} /* (1, 6, 6) {real, imag} */,
  {32'hbe6cd2ec, 32'h3e050018} /* (1, 6, 5) {real, imag} */,
  {32'h3ebb8db3, 32'hbe3f7a34} /* (1, 6, 4) {real, imag} */,
  {32'hbe12ce66, 32'hbe0a7b99} /* (1, 6, 3) {real, imag} */,
  {32'hbd13083a, 32'hbedae54e} /* (1, 6, 2) {real, imag} */,
  {32'hbe6b1d73, 32'h3ef8f41f} /* (1, 6, 1) {real, imag} */,
  {32'h3f0e5d0a, 32'hbf636aa2} /* (1, 6, 0) {real, imag} */,
  {32'h403a7a75, 32'h3e263c01} /* (1, 5, 31) {real, imag} */,
  {32'hbfd200b2, 32'hbe5a0a54} /* (1, 5, 30) {real, imag} */,
  {32'hbf1c3c64, 32'h3efe0336} /* (1, 5, 29) {real, imag} */,
  {32'h3e500b12, 32'h3df7c8c4} /* (1, 5, 28) {real, imag} */,
  {32'h3e14e870, 32'h3e708b84} /* (1, 5, 27) {real, imag} */,
  {32'hbe89540c, 32'hbe0659a0} /* (1, 5, 26) {real, imag} */,
  {32'hbeca9a49, 32'h3dcac330} /* (1, 5, 25) {real, imag} */,
  {32'h3ee0eb45, 32'hbe2859c1} /* (1, 5, 24) {real, imag} */,
  {32'h3de67237, 32'hbe4235e6} /* (1, 5, 23) {real, imag} */,
  {32'hbeef3ca9, 32'hbddb2a3c} /* (1, 5, 22) {real, imag} */,
  {32'hbd74e636, 32'hbe2f373e} /* (1, 5, 21) {real, imag} */,
  {32'h3ed9a23e, 32'hbf2dbab0} /* (1, 5, 20) {real, imag} */,
  {32'h3ea58f90, 32'h3d8d1d31} /* (1, 5, 19) {real, imag} */,
  {32'h3e2c25ed, 32'h3f29d7fd} /* (1, 5, 18) {real, imag} */,
  {32'hbe7e8df4, 32'hbcbb0b80} /* (1, 5, 17) {real, imag} */,
  {32'hbe57aec0, 32'h3e4d419e} /* (1, 5, 16) {real, imag} */,
  {32'hbe191f49, 32'hbddd1643} /* (1, 5, 15) {real, imag} */,
  {32'hbd93eb5b, 32'h3daba0ec} /* (1, 5, 14) {real, imag} */,
  {32'h3f546830, 32'h3e95de7e} /* (1, 5, 13) {real, imag} */,
  {32'hbe2ce988, 32'h3e1df586} /* (1, 5, 12) {real, imag} */,
  {32'hbddcc620, 32'hbdc7cae0} /* (1, 5, 11) {real, imag} */,
  {32'hbde429e1, 32'hbe420fee} /* (1, 5, 10) {real, imag} */,
  {32'h3e397122, 32'h3e86fcf1} /* (1, 5, 9) {real, imag} */,
  {32'hbea3b4e2, 32'h3e0c542b} /* (1, 5, 8) {real, imag} */,
  {32'h3e83a914, 32'h3f228b1a} /* (1, 5, 7) {real, imag} */,
  {32'hbdc50b38, 32'hbd3aa5f8} /* (1, 5, 6) {real, imag} */,
  {32'hbf2f9810, 32'hbf5ca75e} /* (1, 5, 5) {real, imag} */,
  {32'hbdba54a4, 32'h3e73e479} /* (1, 5, 4) {real, imag} */,
  {32'hbea82c4a, 32'hbeb3fcdf} /* (1, 5, 3) {real, imag} */,
  {32'h3ed07e1a, 32'hbf1984ec} /* (1, 5, 2) {real, imag} */,
  {32'h3f94f23c, 32'h40198b9e} /* (1, 5, 1) {real, imag} */,
  {32'h3fe9f865, 32'h3f62d3fc} /* (1, 5, 0) {real, imag} */,
  {32'hc0015b13, 32'hbf83face} /* (1, 4, 31) {real, imag} */,
  {32'h3fb6463c, 32'h402a9da4} /* (1, 4, 30) {real, imag} */,
  {32'hbf20dca4, 32'hbf657670} /* (1, 4, 29) {real, imag} */,
  {32'hbf479f2d, 32'hbe90a672} /* (1, 4, 28) {real, imag} */,
  {32'h3f06b53a, 32'hbe8bf7db} /* (1, 4, 27) {real, imag} */,
  {32'h3ebffdc7, 32'hbee4533c} /* (1, 4, 26) {real, imag} */,
  {32'hbeda273c, 32'hbe693c79} /* (1, 4, 25) {real, imag} */,
  {32'hbe30c3f8, 32'h3e519bf0} /* (1, 4, 24) {real, imag} */,
  {32'hbea8a5ea, 32'hbd1d3c5e} /* (1, 4, 23) {real, imag} */,
  {32'hbe71c418, 32'hbe4049ac} /* (1, 4, 22) {real, imag} */,
  {32'h3e4aad7f, 32'h3c98db48} /* (1, 4, 21) {real, imag} */,
  {32'h3bbb6dc0, 32'h3ee3625f} /* (1, 4, 20) {real, imag} */,
  {32'hbe060f2a, 32'h3eb8a946} /* (1, 4, 19) {real, imag} */,
  {32'h3de64002, 32'h3e3a67af} /* (1, 4, 18) {real, imag} */,
  {32'hbd724d82, 32'hbe8b8125} /* (1, 4, 17) {real, imag} */,
  {32'hbd17e2d1, 32'h3d8ae2d4} /* (1, 4, 16) {real, imag} */,
  {32'h3e419fd7, 32'hbe6b5ae4} /* (1, 4, 15) {real, imag} */,
  {32'hbebf8ab7, 32'h3e848f24} /* (1, 4, 14) {real, imag} */,
  {32'hbdac4d18, 32'h3dbd7285} /* (1, 4, 13) {real, imag} */,
  {32'h3c93d7b0, 32'hbefc6572} /* (1, 4, 12) {real, imag} */,
  {32'h3ec2196a, 32'h3f41e220} /* (1, 4, 11) {real, imag} */,
  {32'h3f0bf991, 32'hbebd8b50} /* (1, 4, 10) {real, imag} */,
  {32'h3f157666, 32'hbdc939f8} /* (1, 4, 9) {real, imag} */,
  {32'h3e9a62b5, 32'h3eced2bc} /* (1, 4, 8) {real, imag} */,
  {32'hbdc7fb76, 32'hbf41493c} /* (1, 4, 7) {real, imag} */,
  {32'h3ea2613e, 32'hbe8287ca} /* (1, 4, 6) {real, imag} */,
  {32'h3ede9a6a, 32'hbe6fd804} /* (1, 4, 5) {real, imag} */,
  {32'hbe437dfe, 32'hbdfeace4} /* (1, 4, 4) {real, imag} */,
  {32'hbe1bed98, 32'h3f60093c} /* (1, 4, 3) {real, imag} */,
  {32'h3ff95d7a, 32'h404ce668} /* (1, 4, 2) {real, imag} */,
  {32'hc08950b2, 32'hbf08f442} /* (1, 4, 1) {real, imag} */,
  {32'hbe736c28, 32'hbeec282c} /* (1, 4, 0) {real, imag} */,
  {32'h4071bf5d, 32'hbfe6f6e8} /* (1, 3, 31) {real, imag} */,
  {32'hbfbd3fcd, 32'h401f93e2} /* (1, 3, 30) {real, imag} */,
  {32'h3dfeba0c, 32'h3e625ee6} /* (1, 3, 29) {real, imag} */,
  {32'hbf3d8d26, 32'hbe61d365} /* (1, 3, 28) {real, imag} */,
  {32'h3f0a60e2, 32'h3e48ee59} /* (1, 3, 27) {real, imag} */,
  {32'hbeed045e, 32'hbe381de8} /* (1, 3, 26) {real, imag} */,
  {32'hbe610c0c, 32'hbd5f7c08} /* (1, 3, 25) {real, imag} */,
  {32'h3e256d94, 32'h3f56d76b} /* (1, 3, 24) {real, imag} */,
  {32'hbd84dfec, 32'hbdc41726} /* (1, 3, 23) {real, imag} */,
  {32'h3dac2f60, 32'h3e4cea51} /* (1, 3, 22) {real, imag} */,
  {32'h3e138120, 32'h3d6ea84c} /* (1, 3, 21) {real, imag} */,
  {32'hbdd8362d, 32'hbe67449f} /* (1, 3, 20) {real, imag} */,
  {32'hbe9d04f2, 32'hbab47c80} /* (1, 3, 19) {real, imag} */,
  {32'hbe8159bf, 32'hbe3b8e81} /* (1, 3, 18) {real, imag} */,
  {32'h3e2b0b36, 32'hbe5f740f} /* (1, 3, 17) {real, imag} */,
  {32'hbe28feef, 32'hbe23aef1} /* (1, 3, 16) {real, imag} */,
  {32'hbdf62f1f, 32'hbe25abd8} /* (1, 3, 15) {real, imag} */,
  {32'h3e517a24, 32'h3c200a20} /* (1, 3, 14) {real, imag} */,
  {32'hbd4c04a8, 32'hbd039dfa} /* (1, 3, 13) {real, imag} */,
  {32'h3f83e9a2, 32'h3e86bbfa} /* (1, 3, 12) {real, imag} */,
  {32'h3cb590bc, 32'h3e03afda} /* (1, 3, 11) {real, imag} */,
  {32'h3ef1946d, 32'hbe0d1c7c} /* (1, 3, 10) {real, imag} */,
  {32'h3eaf9e06, 32'hbe6396cd} /* (1, 3, 9) {real, imag} */,
  {32'hbf480f7f, 32'h3e6ac2d3} /* (1, 3, 8) {real, imag} */,
  {32'hbeb7f387, 32'hbe896234} /* (1, 3, 7) {real, imag} */,
  {32'hbf6c64a1, 32'hbe643823} /* (1, 3, 6) {real, imag} */,
  {32'hbf8aa5ba, 32'h3f4c3352} /* (1, 3, 5) {real, imag} */,
  {32'h3f4f4536, 32'h3f76624c} /* (1, 3, 4) {real, imag} */,
  {32'hbc8ea8a0, 32'hbfd76169} /* (1, 3, 3) {real, imag} */,
  {32'hbeed933c, 32'h40810ee2} /* (1, 3, 2) {real, imag} */,
  {32'hbfe040ab, 32'hbfb0f71b} /* (1, 3, 1) {real, imag} */,
  {32'h3f83a094, 32'hbe019160} /* (1, 3, 0) {real, imag} */,
  {32'h418f74bf, 32'h3ffa5ecc} /* (1, 2, 31) {real, imag} */,
  {32'hc1141f88, 32'h3f2755ad} /* (1, 2, 30) {real, imag} */,
  {32'h3f6ac239, 32'hbf3057f4} /* (1, 2, 29) {real, imag} */,
  {32'h3faede74, 32'hbf10ddc8} /* (1, 2, 28) {real, imag} */,
  {32'hbf8dfeb2, 32'h3fd8bd12} /* (1, 2, 27) {real, imag} */,
  {32'h3e5584f0, 32'hbd05f77c} /* (1, 2, 26) {real, imag} */,
  {32'hbb077180, 32'hbe9fc5a6} /* (1, 2, 25) {real, imag} */,
  {32'hbf84197a, 32'h3f8f10a5} /* (1, 2, 24) {real, imag} */,
  {32'hbe9d502c, 32'h3cbfbcd8} /* (1, 2, 23) {real, imag} */,
  {32'hbd9d6ec2, 32'hbf2495f4} /* (1, 2, 22) {real, imag} */,
  {32'hbe558bcb, 32'h3e9e36ee} /* (1, 2, 21) {real, imag} */,
  {32'h3ddab3fc, 32'h3d0af4f2} /* (1, 2, 20) {real, imag} */,
  {32'hbe0ebab4, 32'hbf0e5fca} /* (1, 2, 19) {real, imag} */,
  {32'hbe72bc28, 32'hbe1c15e1} /* (1, 2, 18) {real, imag} */,
  {32'h3c4c8e70, 32'hbe080d63} /* (1, 2, 17) {real, imag} */,
  {32'hbdcf1f28, 32'h3e163c10} /* (1, 2, 16) {real, imag} */,
  {32'hbc9697ac, 32'h3db2f798} /* (1, 2, 15) {real, imag} */,
  {32'h3e929baf, 32'hbe25698b} /* (1, 2, 14) {real, imag} */,
  {32'h3c03dd34, 32'hbc9152d4} /* (1, 2, 13) {real, imag} */,
  {32'hbe3e1710, 32'h3e6d7e51} /* (1, 2, 12) {real, imag} */,
  {32'hbe858d7c, 32'hbf0e832c} /* (1, 2, 11) {real, imag} */,
  {32'hbd3afe7c, 32'hbdabc9de} /* (1, 2, 10) {real, imag} */,
  {32'h3e0f55cc, 32'hbe3d88ce} /* (1, 2, 9) {real, imag} */,
  {32'hbfb0dda9, 32'hbf50ae8d} /* (1, 2, 8) {real, imag} */,
  {32'h3e7c76e6, 32'h3f489424} /* (1, 2, 7) {real, imag} */,
  {32'hbdc4de90, 32'h3e54c3b8} /* (1, 2, 6) {real, imag} */,
  {32'hbfb43e4e, 32'hbf96daa0} /* (1, 2, 5) {real, imag} */,
  {32'h4059c255, 32'h3f014f84} /* (1, 2, 4) {real, imag} */,
  {32'hbd314b08, 32'hbfa1752f} /* (1, 2, 3) {real, imag} */,
  {32'hc0dea3d9, 32'h40601cae} /* (1, 2, 2) {real, imag} */,
  {32'h41020a3a, 32'h3dcc3680} /* (1, 2, 1) {real, imag} */,
  {32'h40fe832c, 32'h40109d07} /* (1, 2, 0) {real, imag} */,
  {32'hc183a91f, 32'h3fec4749} /* (1, 1, 31) {real, imag} */,
  {32'h40b0976e, 32'hbef7ed99} /* (1, 1, 30) {real, imag} */,
  {32'h3f5b8bbf, 32'hbf148293} /* (1, 1, 29) {real, imag} */,
  {32'hc029ed83, 32'hbf157882} /* (1, 1, 28) {real, imag} */,
  {32'h406dde0b, 32'hbdfa27d4} /* (1, 1, 27) {real, imag} */,
  {32'h3e9ffd6c, 32'hbe825ed4} /* (1, 1, 26) {real, imag} */,
  {32'hbf2bf0db, 32'hbdbb6654} /* (1, 1, 25) {real, imag} */,
  {32'h3f8fce5a, 32'hbf4885b3} /* (1, 1, 24) {real, imag} */,
  {32'hbe09ee3c, 32'hbf2f7294} /* (1, 1, 23) {real, imag} */,
  {32'hbebc61bc, 32'hbd6ceea2} /* (1, 1, 22) {real, imag} */,
  {32'h3f0e4ef0, 32'hbf076ade} /* (1, 1, 21) {real, imag} */,
  {32'hbda15bc4, 32'hbe155167} /* (1, 1, 20) {real, imag} */,
  {32'h3db06312, 32'h3b88d180} /* (1, 1, 19) {real, imag} */,
  {32'hbcc04404, 32'hbd029cc4} /* (1, 1, 18) {real, imag} */,
  {32'hbda598f4, 32'h3e0488f5} /* (1, 1, 17) {real, imag} */,
  {32'hbb465be0, 32'h3d1acad8} /* (1, 1, 16) {real, imag} */,
  {32'h3e7bf15b, 32'hbdfbf001} /* (1, 1, 15) {real, imag} */,
  {32'hbe4cf26a, 32'h3ec8672d} /* (1, 1, 14) {real, imag} */,
  {32'hbeb885de, 32'h3d5a0810} /* (1, 1, 13) {real, imag} */,
  {32'h3e99a388, 32'hbe185f5d} /* (1, 1, 12) {real, imag} */,
  {32'hbe8a07af, 32'h3df5b93a} /* (1, 1, 11) {real, imag} */,
  {32'hbe7a3e6b, 32'hbecd8960} /* (1, 1, 10) {real, imag} */,
  {32'hbe6e5500, 32'h3f42b294} /* (1, 1, 9) {real, imag} */,
  {32'h3ee78477, 32'h3ee9f1c1} /* (1, 1, 8) {real, imag} */,
  {32'hbee6e3e4, 32'hbf816cbe} /* (1, 1, 7) {real, imag} */,
  {32'h3eb2f384, 32'h3ecff0a1} /* (1, 1, 6) {real, imag} */,
  {32'h3ff1ea94, 32'h3f93293c} /* (1, 1, 5) {real, imag} */,
  {32'h3ebed3af, 32'hbfa88e11} /* (1, 1, 4) {real, imag} */,
  {32'h3ff2a66d, 32'h3e36f578} /* (1, 1, 3) {real, imag} */,
  {32'h410ca72a, 32'h40e7a1a0} /* (1, 1, 2) {real, imag} */,
  {32'hc1c06709, 32'hc17a5546} /* (1, 1, 1) {real, imag} */,
  {32'hc17707f3, 32'h40052fc4} /* (1, 1, 0) {real, imag} */,
  {32'hc1320afc, 32'h40db72e7} /* (1, 0, 31) {real, imag} */,
  {32'h3eaf7d10, 32'hc00f4804} /* (1, 0, 30) {real, imag} */,
  {32'h3fb6ff0d, 32'hbf3f489c} /* (1, 0, 29) {real, imag} */,
  {32'hbf5bd2bf, 32'hc00369d2} /* (1, 0, 28) {real, imag} */,
  {32'h400f374c, 32'h3f0e43d0} /* (1, 0, 27) {real, imag} */,
  {32'h3e92bbc5, 32'hbe1a78e3} /* (1, 0, 26) {real, imag} */,
  {32'hbf100e2b, 32'h3f8e648c} /* (1, 0, 25) {real, imag} */,
  {32'hbd369cb0, 32'hbf751311} /* (1, 0, 24) {real, imag} */,
  {32'hbddb412c, 32'hbef24727} /* (1, 0, 23) {real, imag} */,
  {32'h3eb5bd18, 32'h3e980ece} /* (1, 0, 22) {real, imag} */,
  {32'h3f068c37, 32'hbdfb6c40} /* (1, 0, 21) {real, imag} */,
  {32'h3ea95788, 32'h3eca5be8} /* (1, 0, 20) {real, imag} */,
  {32'h3ea19658, 32'h3eb72024} /* (1, 0, 19) {real, imag} */,
  {32'hbdd5fe0a, 32'hbf2da58a} /* (1, 0, 18) {real, imag} */,
  {32'hbeb4423a, 32'h3dbbb1e4} /* (1, 0, 17) {real, imag} */,
  {32'h3e0ba361, 32'h00000000} /* (1, 0, 16) {real, imag} */,
  {32'hbeb4423a, 32'hbdbbb1e4} /* (1, 0, 15) {real, imag} */,
  {32'hbdd5fe0a, 32'h3f2da58a} /* (1, 0, 14) {real, imag} */,
  {32'h3ea19658, 32'hbeb72024} /* (1, 0, 13) {real, imag} */,
  {32'h3ea95788, 32'hbeca5be8} /* (1, 0, 12) {real, imag} */,
  {32'h3f068c37, 32'h3dfb6c40} /* (1, 0, 11) {real, imag} */,
  {32'h3eb5bd18, 32'hbe980ece} /* (1, 0, 10) {real, imag} */,
  {32'hbddb412c, 32'h3ef24727} /* (1, 0, 9) {real, imag} */,
  {32'hbd369cb0, 32'h3f751311} /* (1, 0, 8) {real, imag} */,
  {32'hbf100e2b, 32'hbf8e648c} /* (1, 0, 7) {real, imag} */,
  {32'h3e92bbc5, 32'h3e1a78e3} /* (1, 0, 6) {real, imag} */,
  {32'h400f374c, 32'hbf0e43d0} /* (1, 0, 5) {real, imag} */,
  {32'hbf5bd2bf, 32'h400369d2} /* (1, 0, 4) {real, imag} */,
  {32'h3fb6ff0d, 32'h3f3f489c} /* (1, 0, 3) {real, imag} */,
  {32'h3eaf7d10, 32'h400f4804} /* (1, 0, 2) {real, imag} */,
  {32'hc1320afc, 32'hc0db72e7} /* (1, 0, 1) {real, imag} */,
  {32'hc0c89817, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hc1210d46, 32'h4103b8de} /* (0, 31, 31) {real, imag} */,
  {32'h4032ad2b, 32'hbfd8411c} /* (0, 31, 30) {real, imag} */,
  {32'h3fcebd20, 32'h3da9676e} /* (0, 31, 29) {real, imag} */,
  {32'h3effe53b, 32'h3f02d502} /* (0, 31, 28) {real, imag} */,
  {32'h3f1b3910, 32'hbed2d494} /* (0, 31, 27) {real, imag} */,
  {32'h3efe81df, 32'hbe68c852} /* (0, 31, 26) {real, imag} */,
  {32'hbe492e41, 32'h3e613823} /* (0, 31, 25) {real, imag} */,
  {32'hbdc95710, 32'hbf0ae0d9} /* (0, 31, 24) {real, imag} */,
  {32'hbdb5966f, 32'h3e1c186a} /* (0, 31, 23) {real, imag} */,
  {32'hbe3aef38, 32'h3e68e6e2} /* (0, 31, 22) {real, imag} */,
  {32'h3efd81e2, 32'h3d4a66d0} /* (0, 31, 21) {real, imag} */,
  {32'hbd91da41, 32'h3e0e09c6} /* (0, 31, 20) {real, imag} */,
  {32'h3e6b60be, 32'h3e565758} /* (0, 31, 19) {real, imag} */,
  {32'hbe1b913e, 32'h3d810da8} /* (0, 31, 18) {real, imag} */,
  {32'h3e51671a, 32'hbce35cb4} /* (0, 31, 17) {real, imag} */,
  {32'h3d964b88, 32'h3dc5bb2c} /* (0, 31, 16) {real, imag} */,
  {32'h3d53c3fc, 32'h3e656e7c} /* (0, 31, 15) {real, imag} */,
  {32'h3e3ec258, 32'h3d584e8a} /* (0, 31, 14) {real, imag} */,
  {32'h3c8f7db8, 32'h3e145df1} /* (0, 31, 13) {real, imag} */,
  {32'hbd31340a, 32'hbeda5d96} /* (0, 31, 12) {real, imag} */,
  {32'h3e9387d7, 32'h3f01534a} /* (0, 31, 11) {real, imag} */,
  {32'hbe826137, 32'hbeadc5ba} /* (0, 31, 10) {real, imag} */,
  {32'h3ee52414, 32'h3f02562b} /* (0, 31, 9) {real, imag} */,
  {32'h3e0c6d49, 32'h3ec55d3b} /* (0, 31, 8) {real, imag} */,
  {32'hbe134e91, 32'h3e6ace5c} /* (0, 31, 7) {real, imag} */,
  {32'hbc981580, 32'hbe2ac079} /* (0, 31, 6) {real, imag} */,
  {32'h3ffc6b5a, 32'hbed2b368} /* (0, 31, 5) {real, imag} */,
  {32'hbf8ab738, 32'h3d6f9e20} /* (0, 31, 4) {real, imag} */,
  {32'h3f6e39b6, 32'hbc65b580} /* (0, 31, 3) {real, imag} */,
  {32'h3ffd3b82, 32'h3ed2b7fe} /* (0, 31, 2) {real, imag} */,
  {32'hc0c0868e, 32'h3e54e948} /* (0, 31, 1) {real, imag} */,
  {32'hc0da7e04, 32'hc023a2bb} /* (0, 31, 0) {real, imag} */,
  {32'h40205470, 32'hbf21e13a} /* (0, 30, 31) {real, imag} */,
  {32'hc03a574a, 32'hbfdc7406} /* (0, 30, 30) {real, imag} */,
  {32'hbe81ae78, 32'h3f32e1fd} /* (0, 30, 29) {real, imag} */,
  {32'h3feb503f, 32'hbeab9a7c} /* (0, 30, 28) {real, imag} */,
  {32'hbf414726, 32'h3f7d7cca} /* (0, 30, 27) {real, imag} */,
  {32'h3f065b1a, 32'hbebc831f} /* (0, 30, 26) {real, imag} */,
  {32'h3eb53c14, 32'hbd8fd624} /* (0, 30, 25) {real, imag} */,
  {32'hbf578e4e, 32'h3ea76c4c} /* (0, 30, 24) {real, imag} */,
  {32'hbe57c989, 32'h3e17beb0} /* (0, 30, 23) {real, imag} */,
  {32'hbe1f318b, 32'h3e733898} /* (0, 30, 22) {real, imag} */,
  {32'hbda9148e, 32'h3f1a7ce4} /* (0, 30, 21) {real, imag} */,
  {32'h3e140a1a, 32'h3ed4c76c} /* (0, 30, 20) {real, imag} */,
  {32'hbeac2314, 32'h3b5147c0} /* (0, 30, 19) {real, imag} */,
  {32'hbd64927c, 32'h3e422bf2} /* (0, 30, 18) {real, imag} */,
  {32'h3eb94f7b, 32'h3d88a388} /* (0, 30, 17) {real, imag} */,
  {32'h3d866a5d, 32'hbc42bb98} /* (0, 30, 16) {real, imag} */,
  {32'h3d2166da, 32'hbde5dc8d} /* (0, 30, 15) {real, imag} */,
  {32'h3d18607a, 32'h3c150cc8} /* (0, 30, 14) {real, imag} */,
  {32'hbd8fdfd8, 32'hbc2b661c} /* (0, 30, 13) {real, imag} */,
  {32'hbe8dc2ff, 32'hbd95b914} /* (0, 30, 12) {real, imag} */,
  {32'hbe25812b, 32'h3e2b840c} /* (0, 30, 11) {real, imag} */,
  {32'h3d7fac9e, 32'hbd518d80} /* (0, 30, 10) {real, imag} */,
  {32'h3c2a9ca0, 32'hbd7d2270} /* (0, 30, 9) {real, imag} */,
  {32'hbeac923b, 32'hbee8ff5c} /* (0, 30, 8) {real, imag} */,
  {32'hbd259288, 32'hbe8f07cc} /* (0, 30, 7) {real, imag} */,
  {32'hbe2b37a6, 32'hbec75e7f} /* (0, 30, 6) {real, imag} */,
  {32'hbf1ec512, 32'hbf8ea3fe} /* (0, 30, 5) {real, imag} */,
  {32'h3ed61c24, 32'h3e4e82a8} /* (0, 30, 4) {real, imag} */,
  {32'h3ee5c05c, 32'h3f5defee} /* (0, 30, 3) {real, imag} */,
  {32'hc07bb0a2, 32'hbe0d3768} /* (0, 30, 2) {real, imag} */,
  {32'h40f44033, 32'hbe862dad} /* (0, 30, 1) {real, imag} */,
  {32'h402d914c, 32'hbf3351a6} /* (0, 30, 0) {real, imag} */,
  {32'hbf02c6cb, 32'h3f9ab240} /* (0, 29, 31) {real, imag} */,
  {32'hbf370cdb, 32'hbfdbd312} /* (0, 29, 30) {real, imag} */,
  {32'h3eaf456d, 32'h3f5b544e} /* (0, 29, 29) {real, imag} */,
  {32'h3f16c8c0, 32'hbf7f74dc} /* (0, 29, 28) {real, imag} */,
  {32'hbe8dcb31, 32'hbeac67e3} /* (0, 29, 27) {real, imag} */,
  {32'hbeb37fe9, 32'h3ef4799d} /* (0, 29, 26) {real, imag} */,
  {32'hbf457eec, 32'h3da5fdee} /* (0, 29, 25) {real, imag} */,
  {32'h3e8c4836, 32'hbcc3eca8} /* (0, 29, 24) {real, imag} */,
  {32'h3d17a1b0, 32'h3e9885db} /* (0, 29, 23) {real, imag} */,
  {32'h3dffded0, 32'hbd0f6e84} /* (0, 29, 22) {real, imag} */,
  {32'h3e486d54, 32'hbe1ab7b3} /* (0, 29, 21) {real, imag} */,
  {32'h3ec52218, 32'hbd5b2794} /* (0, 29, 20) {real, imag} */,
  {32'hbddd2074, 32'h3e456582} /* (0, 29, 19) {real, imag} */,
  {32'hbea03e7d, 32'h3bd1d0b0} /* (0, 29, 18) {real, imag} */,
  {32'h3dda3198, 32'h3cd62a30} /* (0, 29, 17) {real, imag} */,
  {32'h3b585e60, 32'hbe764c0b} /* (0, 29, 16) {real, imag} */,
  {32'h3df7e26c, 32'h3dc6c0ce} /* (0, 29, 15) {real, imag} */,
  {32'hbea9fc0a, 32'hbdcf693f} /* (0, 29, 14) {real, imag} */,
  {32'h3ba7c4c0, 32'hbe746267} /* (0, 29, 13) {real, imag} */,
  {32'hbe88847e, 32'hbe0f7f18} /* (0, 29, 12) {real, imag} */,
  {32'hbe30606e, 32'hbe074786} /* (0, 29, 11) {real, imag} */,
  {32'hbe65b4d7, 32'h3e0f8d13} /* (0, 29, 10) {real, imag} */,
  {32'hbe274892, 32'hba7d0b40} /* (0, 29, 9) {real, imag} */,
  {32'h3e6592e6, 32'hbec32a4e} /* (0, 29, 8) {real, imag} */,
  {32'hbd3e1d08, 32'h3eb338ee} /* (0, 29, 7) {real, imag} */,
  {32'h3ce8ed32, 32'hbe0d7896} /* (0, 29, 6) {real, imag} */,
  {32'h3ef66c44, 32'h3f00d3a8} /* (0, 29, 5) {real, imag} */,
  {32'hbec4cc1f, 32'h3e108fb3} /* (0, 29, 4) {real, imag} */,
  {32'h3f233db4, 32'hbecf82f2} /* (0, 29, 3) {real, imag} */,
  {32'hbf1e0af6, 32'hbf06614a} /* (0, 29, 2) {real, imag} */,
  {32'h3fb3a764, 32'h3e63c504} /* (0, 29, 1) {real, imag} */,
  {32'h3f5e95d2, 32'hbed052ca} /* (0, 29, 0) {real, imag} */,
  {32'hbfb201f0, 32'hbec2a4a8} /* (0, 28, 31) {real, imag} */,
  {32'h3f28f9f0, 32'hbf79347e} /* (0, 28, 30) {real, imag} */,
  {32'h3e7011c4, 32'hbf805571} /* (0, 28, 29) {real, imag} */,
  {32'h3bef90c0, 32'hbcee57e0} /* (0, 28, 28) {real, imag} */,
  {32'h3e9ecd13, 32'h3c908ab8} /* (0, 28, 27) {real, imag} */,
  {32'hbde01044, 32'hbdc2bed8} /* (0, 28, 26) {real, imag} */,
  {32'hbea48d1c, 32'h3f074adc} /* (0, 28, 25) {real, imag} */,
  {32'h3ea8080e, 32'hbc8e2758} /* (0, 28, 24) {real, imag} */,
  {32'h3e3a30ce, 32'hbe64d338} /* (0, 28, 23) {real, imag} */,
  {32'h3ee62196, 32'hbe3933a0} /* (0, 28, 22) {real, imag} */,
  {32'hbe0d3248, 32'hbeb7699d} /* (0, 28, 21) {real, imag} */,
  {32'h3dc4ab8b, 32'h3d963b42} /* (0, 28, 20) {real, imag} */,
  {32'h3d6cef18, 32'hbca8af5c} /* (0, 28, 19) {real, imag} */,
  {32'hbdda7a3a, 32'hbe6efe3a} /* (0, 28, 18) {real, imag} */,
  {32'hbcef2788, 32'h3d08e8af} /* (0, 28, 17) {real, imag} */,
  {32'h3e27c95a, 32'h3e1e68fa} /* (0, 28, 16) {real, imag} */,
  {32'hbdaba366, 32'h3dc064af} /* (0, 28, 15) {real, imag} */,
  {32'h3d651bad, 32'hbeb03466} /* (0, 28, 14) {real, imag} */,
  {32'hbeaa9756, 32'hbe4a0ea1} /* (0, 28, 13) {real, imag} */,
  {32'hbe6c5250, 32'hbe66bfde} /* (0, 28, 12) {real, imag} */,
  {32'h3dc64a1a, 32'h3d87eb44} /* (0, 28, 11) {real, imag} */,
  {32'hbe050e62, 32'hbd0eb1b6} /* (0, 28, 10) {real, imag} */,
  {32'hbf11d060, 32'h3eef9dcf} /* (0, 28, 9) {real, imag} */,
  {32'hbdaf0890, 32'h3f0a6271} /* (0, 28, 8) {real, imag} */,
  {32'h3f4cb336, 32'hbf0bce38} /* (0, 28, 7) {real, imag} */,
  {32'h3d566aa0, 32'h3e9ad78c} /* (0, 28, 6) {real, imag} */,
  {32'hbd481890, 32'h3e61c18b} /* (0, 28, 5) {real, imag} */,
  {32'hbe249ea4, 32'hbe84c117} /* (0, 28, 4) {real, imag} */,
  {32'hbeb63d48, 32'h3e83d145} /* (0, 28, 3) {real, imag} */,
  {32'hbe0e65d8, 32'hbfa8d210} /* (0, 28, 2) {real, imag} */,
  {32'hbf5afaea, 32'h3f081c40} /* (0, 28, 1) {real, imag} */,
  {32'h3f344f1b, 32'h3ebf2c90} /* (0, 28, 0) {real, imag} */,
  {32'hbe998fdb, 32'hbf57dc4d} /* (0, 27, 31) {real, imag} */,
  {32'h3ebddea6, 32'h3edcdc75} /* (0, 27, 30) {real, imag} */,
  {32'hbeaff2a9, 32'h3e9e4730} /* (0, 27, 29) {real, imag} */,
  {32'hbe3ca84a, 32'hbeedb3a4} /* (0, 27, 28) {real, imag} */,
  {32'h3e33d0be, 32'hbe3f2f64} /* (0, 27, 27) {real, imag} */,
  {32'hbed97cb2, 32'hbe382e02} /* (0, 27, 26) {real, imag} */,
  {32'h3eb99b89, 32'hbdaf1e4e} /* (0, 27, 25) {real, imag} */,
  {32'h3c1bd958, 32'hbb4c4700} /* (0, 27, 24) {real, imag} */,
  {32'h3e1e367b, 32'h3db7d278} /* (0, 27, 23) {real, imag} */,
  {32'hbe4517f8, 32'hbe2691d6} /* (0, 27, 22) {real, imag} */,
  {32'hbb9c2280, 32'h3eae8819} /* (0, 27, 21) {real, imag} */,
  {32'hbe487ffa, 32'hbd4c1718} /* (0, 27, 20) {real, imag} */,
  {32'h3e1ef95f, 32'hbe5f9f68} /* (0, 27, 19) {real, imag} */,
  {32'h3e5c2cb4, 32'h3ded3b7d} /* (0, 27, 18) {real, imag} */,
  {32'h3e3b2a26, 32'h3e215a44} /* (0, 27, 17) {real, imag} */,
  {32'hbd572b74, 32'hbe3f6484} /* (0, 27, 16) {real, imag} */,
  {32'hbd32b73a, 32'h3e060916} /* (0, 27, 15) {real, imag} */,
  {32'hbe673106, 32'hbe9b38c9} /* (0, 27, 14) {real, imag} */,
  {32'h3e29dc56, 32'hbd1396f8} /* (0, 27, 13) {real, imag} */,
  {32'hbe593810, 32'h3e384952} /* (0, 27, 12) {real, imag} */,
  {32'hbef21631, 32'h3e1a8403} /* (0, 27, 11) {real, imag} */,
  {32'hbeca591c, 32'hbe884caf} /* (0, 27, 10) {real, imag} */,
  {32'h3e0373c4, 32'hbd682520} /* (0, 27, 9) {real, imag} */,
  {32'hbdbe4454, 32'h3ed63453} /* (0, 27, 8) {real, imag} */,
  {32'hbe36de07, 32'hbb8e9f00} /* (0, 27, 7) {real, imag} */,
  {32'h3eabec51, 32'hbe0adcee} /* (0, 27, 6) {real, imag} */,
  {32'h3e18191d, 32'hbe88a1b4} /* (0, 27, 5) {real, imag} */,
  {32'h3ec23f02, 32'hbd1bbcb8} /* (0, 27, 4) {real, imag} */,
  {32'hbf0b99ef, 32'hbecb6c8e} /* (0, 27, 3) {real, imag} */,
  {32'hbf2d3a30, 32'hbe617768} /* (0, 27, 2) {real, imag} */,
  {32'h3f8ebaf4, 32'h3ebe497d} /* (0, 27, 1) {real, imag} */,
  {32'h3f6f0010, 32'h3dbbaf20} /* (0, 27, 0) {real, imag} */,
  {32'hbe6b36e7, 32'h3e30d796} /* (0, 26, 31) {real, imag} */,
  {32'hbddc1a98, 32'h3e6eb2bc} /* (0, 26, 30) {real, imag} */,
  {32'h3ed50ada, 32'hbdb45c6d} /* (0, 26, 29) {real, imag} */,
  {32'h3f0716b4, 32'h3e8eb088} /* (0, 26, 28) {real, imag} */,
  {32'hbe4ce642, 32'h3da64dfd} /* (0, 26, 27) {real, imag} */,
  {32'hbec5b992, 32'hbe091e86} /* (0, 26, 26) {real, imag} */,
  {32'h3dd53024, 32'hbe1c772a} /* (0, 26, 25) {real, imag} */,
  {32'h3d01fe79, 32'h3e8c96dc} /* (0, 26, 24) {real, imag} */,
  {32'h3e8145e6, 32'h3e0af1ed} /* (0, 26, 23) {real, imag} */,
  {32'hbe715624, 32'hbee03869} /* (0, 26, 22) {real, imag} */,
  {32'hbd8182cc, 32'hbe83ac96} /* (0, 26, 21) {real, imag} */,
  {32'hbc47f460, 32'hbe8c3284} /* (0, 26, 20) {real, imag} */,
  {32'h3cdb65c0, 32'h3e4133c4} /* (0, 26, 19) {real, imag} */,
  {32'hbeb99698, 32'hbec5a30d} /* (0, 26, 18) {real, imag} */,
  {32'hbdcf2eee, 32'h3ddbb8f9} /* (0, 26, 17) {real, imag} */,
  {32'h3d3f7191, 32'hbe3c1f6a} /* (0, 26, 16) {real, imag} */,
  {32'h3e417bbd, 32'hbb8a4338} /* (0, 26, 15) {real, imag} */,
  {32'h3d586e88, 32'hbcc56300} /* (0, 26, 14) {real, imag} */,
  {32'h3e42233c, 32'h3e037bce} /* (0, 26, 13) {real, imag} */,
  {32'h3e3ae08d, 32'hbc632920} /* (0, 26, 12) {real, imag} */,
  {32'h3e827bd2, 32'h3c6a96f8} /* (0, 26, 11) {real, imag} */,
  {32'hbdc18b20, 32'h3e119bd7} /* (0, 26, 10) {real, imag} */,
  {32'h3e7d5bbc, 32'h3da83170} /* (0, 26, 9) {real, imag} */,
  {32'hbcfa254c, 32'h3e29e5ad} /* (0, 26, 8) {real, imag} */,
  {32'h3eaa21b2, 32'hbdea7ee0} /* (0, 26, 7) {real, imag} */,
  {32'h3d795568, 32'hbe25c11a} /* (0, 26, 6) {real, imag} */,
  {32'h3f038458, 32'h3e65e4a5} /* (0, 26, 5) {real, imag} */,
  {32'hbe296ee3, 32'hbedcf7c7} /* (0, 26, 4) {real, imag} */,
  {32'h3e8488b7, 32'h3f638a55} /* (0, 26, 3) {real, imag} */,
  {32'hbf4e89bd, 32'hbf1e2916} /* (0, 26, 2) {real, imag} */,
  {32'hbd822fbc, 32'hbf019710} /* (0, 26, 1) {real, imag} */,
  {32'hbda6a99e, 32'h3f7c7d9c} /* (0, 26, 0) {real, imag} */,
  {32'h3f596da6, 32'h3f487663} /* (0, 25, 31) {real, imag} */,
  {32'hbef4a89c, 32'h3eae7ef2} /* (0, 25, 30) {real, imag} */,
  {32'h3e45e34e, 32'h3e11ed56} /* (0, 25, 29) {real, imag} */,
  {32'h3e3bdf66, 32'hbcf69778} /* (0, 25, 28) {real, imag} */,
  {32'h3e92a3c2, 32'hbea9f5e2} /* (0, 25, 27) {real, imag} */,
  {32'hbee17a78, 32'hbe90177a} /* (0, 25, 26) {real, imag} */,
  {32'hbe9da280, 32'h3d84d830} /* (0, 25, 25) {real, imag} */,
  {32'hbd9e525e, 32'h3e560bf1} /* (0, 25, 24) {real, imag} */,
  {32'h3e518d0e, 32'hbe354ca8} /* (0, 25, 23) {real, imag} */,
  {32'hbe3b40a9, 32'h3e54bbe8} /* (0, 25, 22) {real, imag} */,
  {32'h3e5143f1, 32'hbdb41e54} /* (0, 25, 21) {real, imag} */,
  {32'hbe32a501, 32'hbe92f19e} /* (0, 25, 20) {real, imag} */,
  {32'hbb095340, 32'hbe961296} /* (0, 25, 19) {real, imag} */,
  {32'h3e53a96e, 32'h3e01df98} /* (0, 25, 18) {real, imag} */,
  {32'hbb753800, 32'hbdf80a80} /* (0, 25, 17) {real, imag} */,
  {32'hbdc39498, 32'h3e8d5fe4} /* (0, 25, 16) {real, imag} */,
  {32'hbe2ec7b8, 32'hbdb4d5c0} /* (0, 25, 15) {real, imag} */,
  {32'hbe8ec66e, 32'h3d505e94} /* (0, 25, 14) {real, imag} */,
  {32'hbc2127e0, 32'hbe55de2a} /* (0, 25, 13) {real, imag} */,
  {32'h39a3a800, 32'h3d50d9da} /* (0, 25, 12) {real, imag} */,
  {32'h3e40076c, 32'h3caf30f0} /* (0, 25, 11) {real, imag} */,
  {32'h3ddc391c, 32'h3e38618f} /* (0, 25, 10) {real, imag} */,
  {32'hbd6621b4, 32'h3c8ceee0} /* (0, 25, 9) {real, imag} */,
  {32'h3e08ba00, 32'h3e15ea24} /* (0, 25, 8) {real, imag} */,
  {32'h3dc9718e, 32'h3c858ea8} /* (0, 25, 7) {real, imag} */,
  {32'hbe2d4f6c, 32'hbcddc930} /* (0, 25, 6) {real, imag} */,
  {32'hbe252ca6, 32'h3dc39573} /* (0, 25, 5) {real, imag} */,
  {32'h3e95bab6, 32'hbed9c31b} /* (0, 25, 4) {real, imag} */,
  {32'hbe77c858, 32'hbf08692d} /* (0, 25, 3) {real, imag} */,
  {32'h3eb5eefe, 32'hb9fe4400} /* (0, 25, 2) {real, imag} */,
  {32'hbe228002, 32'hbe9cad96} /* (0, 25, 1) {real, imag} */,
  {32'hbdd7ffec, 32'h3ea0a24c} /* (0, 25, 0) {real, imag} */,
  {32'h3d1c3980, 32'hbf215289} /* (0, 24, 31) {real, imag} */,
  {32'hbf095349, 32'hbe099336} /* (0, 24, 30) {real, imag} */,
  {32'hbf01de38, 32'hbe047694} /* (0, 24, 29) {real, imag} */,
  {32'h3d9dca6a, 32'hbd93c4b8} /* (0, 24, 28) {real, imag} */,
  {32'h3e7d9973, 32'h3e5d3c6a} /* (0, 24, 27) {real, imag} */,
  {32'hbea76a7e, 32'h3e849026} /* (0, 24, 26) {real, imag} */,
  {32'h3e68aebc, 32'hbebc7027} /* (0, 24, 25) {real, imag} */,
  {32'h3de2c7ba, 32'h3cd03f30} /* (0, 24, 24) {real, imag} */,
  {32'hbd8960bc, 32'h3d019d68} /* (0, 24, 23) {real, imag} */,
  {32'hbeb63392, 32'hbdb29500} /* (0, 24, 22) {real, imag} */,
  {32'h3e90954c, 32'h3e4322b9} /* (0, 24, 21) {real, imag} */,
  {32'hbe35ab09, 32'h3e2b1723} /* (0, 24, 20) {real, imag} */,
  {32'hbdc350fc, 32'hbe8e22ae} /* (0, 24, 19) {real, imag} */,
  {32'h3e5c36e6, 32'hbed2eba7} /* (0, 24, 18) {real, imag} */,
  {32'h3dd755f0, 32'hbccc52b0} /* (0, 24, 17) {real, imag} */,
  {32'hbcb1fc00, 32'h3eb5419e} /* (0, 24, 16) {real, imag} */,
  {32'hbdc98d65, 32'h3d947032} /* (0, 24, 15) {real, imag} */,
  {32'h3ead80d0, 32'h3e0ca485} /* (0, 24, 14) {real, imag} */,
  {32'h3e687837, 32'hbe21c36d} /* (0, 24, 13) {real, imag} */,
  {32'hbe3f7d6b, 32'h3d3ea540} /* (0, 24, 12) {real, imag} */,
  {32'hbe29e3f4, 32'hbeba7491} /* (0, 24, 11) {real, imag} */,
  {32'hbe7ce8e5, 32'h3ee69015} /* (0, 24, 10) {real, imag} */,
  {32'h3ebc6d8b, 32'h3e0b0487} /* (0, 24, 9) {real, imag} */,
  {32'hbefcc5e2, 32'hbe3510ec} /* (0, 24, 8) {real, imag} */,
  {32'h3e8b3d56, 32'h3eb9ac7d} /* (0, 24, 7) {real, imag} */,
  {32'h3e2eaff6, 32'hbd9deacc} /* (0, 24, 6) {real, imag} */,
  {32'hbe00034a, 32'h3e2e6ea0} /* (0, 24, 5) {real, imag} */,
  {32'h3ef610dc, 32'h3e16e9e6} /* (0, 24, 4) {real, imag} */,
  {32'hbcbcf3d8, 32'h3e1037e1} /* (0, 24, 3) {real, imag} */,
  {32'hbf864771, 32'h3e869517} /* (0, 24, 2) {real, imag} */,
  {32'h3e4c7b92, 32'hbf0850e1} /* (0, 24, 1) {real, imag} */,
  {32'h3f31299e, 32'hbf15be20} /* (0, 24, 0) {real, imag} */,
  {32'hbf1d2422, 32'hbe07ce90} /* (0, 23, 31) {real, imag} */,
  {32'h3d3e5a24, 32'hbccc68c0} /* (0, 23, 30) {real, imag} */,
  {32'hbd62ccbc, 32'h3eb84dc6} /* (0, 23, 29) {real, imag} */,
  {32'hbd991e32, 32'hbe82cb4f} /* (0, 23, 28) {real, imag} */,
  {32'hbcd8159a, 32'hbd8fc468} /* (0, 23, 27) {real, imag} */,
  {32'h3ea15090, 32'hbd2aa520} /* (0, 23, 26) {real, imag} */,
  {32'h3dd6d538, 32'hbd41c0f2} /* (0, 23, 25) {real, imag} */,
  {32'hbd5ff710, 32'hbec85cc8} /* (0, 23, 24) {real, imag} */,
  {32'hbe5bfd9e, 32'h3d863f86} /* (0, 23, 23) {real, imag} */,
  {32'h3e7b4aa0, 32'hbe94dc92} /* (0, 23, 22) {real, imag} */,
  {32'hbeece180, 32'hbbe24fc0} /* (0, 23, 21) {real, imag} */,
  {32'h3e9a2ed5, 32'hbe887a14} /* (0, 23, 20) {real, imag} */,
  {32'hbd737254, 32'hbc54f2a8} /* (0, 23, 19) {real, imag} */,
  {32'hbe87b8ca, 32'hbb2b0560} /* (0, 23, 18) {real, imag} */,
  {32'h3d4d0d20, 32'h3d9ec486} /* (0, 23, 17) {real, imag} */,
  {32'h3e18bb41, 32'h3c008c40} /* (0, 23, 16) {real, imag} */,
  {32'hbde5454f, 32'h3e4a01d3} /* (0, 23, 15) {real, imag} */,
  {32'hbe426d7d, 32'hbdd1c736} /* (0, 23, 14) {real, imag} */,
  {32'h3e45325c, 32'hbc242578} /* (0, 23, 13) {real, imag} */,
  {32'h3ce7ee98, 32'h3e445ea4} /* (0, 23, 12) {real, imag} */,
  {32'hbc961320, 32'hbcf1d198} /* (0, 23, 11) {real, imag} */,
  {32'hbb284880, 32'hbea560ce} /* (0, 23, 10) {real, imag} */,
  {32'h3d491348, 32'hbdd6c3f6} /* (0, 23, 9) {real, imag} */,
  {32'h3e2f73ce, 32'h3ea8cbb5} /* (0, 23, 8) {real, imag} */,
  {32'h3e9bcfd6, 32'h3c94dd58} /* (0, 23, 7) {real, imag} */,
  {32'hbcf691a0, 32'h3e5ec45f} /* (0, 23, 6) {real, imag} */,
  {32'h3e6cf843, 32'h3ca73028} /* (0, 23, 5) {real, imag} */,
  {32'hbecee360, 32'h3f0cf41b} /* (0, 23, 4) {real, imag} */,
  {32'hbf2dc512, 32'hbec1766c} /* (0, 23, 3) {real, imag} */,
  {32'h3f1e3a69, 32'hbf02174f} /* (0, 23, 2) {real, imag} */,
  {32'h3c5c3c28, 32'h3e0d45cf} /* (0, 23, 1) {real, imag} */,
  {32'hbecf06c5, 32'h3e08554c} /* (0, 23, 0) {real, imag} */,
  {32'hbf1a8a3c, 32'h3c27da90} /* (0, 22, 31) {real, imag} */,
  {32'h3f17403c, 32'hbf3ef3a2} /* (0, 22, 30) {real, imag} */,
  {32'hbd48e058, 32'hbda6387b} /* (0, 22, 29) {real, imag} */,
  {32'h3e085a68, 32'h3e8568ba} /* (0, 22, 28) {real, imag} */,
  {32'hbdd6b508, 32'h3c334c28} /* (0, 22, 27) {real, imag} */,
  {32'hbd746e2c, 32'h3ce63958} /* (0, 22, 26) {real, imag} */,
  {32'h3e0d32b6, 32'h3db87fa8} /* (0, 22, 25) {real, imag} */,
  {32'h3e18f172, 32'h3dcffbb4} /* (0, 22, 24) {real, imag} */,
  {32'h3d5080fa, 32'h3eeaf5ae} /* (0, 22, 23) {real, imag} */,
  {32'h3e865f62, 32'h3dfea096} /* (0, 22, 22) {real, imag} */,
  {32'h3e2645f5, 32'h3daf4698} /* (0, 22, 21) {real, imag} */,
  {32'hbedc6ba2, 32'h3ee8ca45} /* (0, 22, 20) {real, imag} */,
  {32'h3eb29ef4, 32'h3d8b6914} /* (0, 22, 19) {real, imag} */,
  {32'h3e30295c, 32'h3e0f237e} /* (0, 22, 18) {real, imag} */,
  {32'hbdfcda8c, 32'hbde25f92} /* (0, 22, 17) {real, imag} */,
  {32'h3d80c70a, 32'h3e2d92bc} /* (0, 22, 16) {real, imag} */,
  {32'h3ccd43ec, 32'hbb0fbd00} /* (0, 22, 15) {real, imag} */,
  {32'hbe312066, 32'h3d6eb666} /* (0, 22, 14) {real, imag} */,
  {32'h3e1af9f8, 32'hbca74830} /* (0, 22, 13) {real, imag} */,
  {32'h3dcd83c4, 32'hbe74f3b2} /* (0, 22, 12) {real, imag} */,
  {32'h3dcfbbfc, 32'h3e603e80} /* (0, 22, 11) {real, imag} */,
  {32'hbe10570f, 32'h3e4502aa} /* (0, 22, 10) {real, imag} */,
  {32'h3e588486, 32'h3ebb5b48} /* (0, 22, 9) {real, imag} */,
  {32'h3ee739a8, 32'h3e8964e2} /* (0, 22, 8) {real, imag} */,
  {32'h3c97c970, 32'h3dea99db} /* (0, 22, 7) {real, imag} */,
  {32'hbd1dd44c, 32'hbeae7ede} /* (0, 22, 6) {real, imag} */,
  {32'h3ef420ec, 32'hbe216d08} /* (0, 22, 5) {real, imag} */,
  {32'hbe997e51, 32'h3e94e99f} /* (0, 22, 4) {real, imag} */,
  {32'hbe09faa3, 32'h3dd393fd} /* (0, 22, 3) {real, imag} */,
  {32'hbcde3410, 32'hbe882b57} /* (0, 22, 2) {real, imag} */,
  {32'hbd083304, 32'h3da16f7e} /* (0, 22, 1) {real, imag} */,
  {32'h3ded1ed8, 32'h3d92ae52} /* (0, 22, 0) {real, imag} */,
  {32'h3e06507f, 32'h3e027d23} /* (0, 21, 31) {real, imag} */,
  {32'h3dd5c0b4, 32'h3ec0fcdd} /* (0, 21, 30) {real, imag} */,
  {32'h3e539569, 32'h3da46088} /* (0, 21, 29) {real, imag} */,
  {32'hbde18ee6, 32'h3eab2984} /* (0, 21, 28) {real, imag} */,
  {32'hbebc1c0e, 32'hbe5ca805} /* (0, 21, 27) {real, imag} */,
  {32'h3dd2335c, 32'h3dbf15e8} /* (0, 21, 26) {real, imag} */,
  {32'h3e04aa46, 32'h3d0404ad} /* (0, 21, 25) {real, imag} */,
  {32'hbd94bec8, 32'hbe6c6655} /* (0, 21, 24) {real, imag} */,
  {32'h3dec915e, 32'hbda091b0} /* (0, 21, 23) {real, imag} */,
  {32'hbf5bcabc, 32'h3e27c818} /* (0, 21, 22) {real, imag} */,
  {32'h3e93d3dd, 32'h3df88aaf} /* (0, 21, 21) {real, imag} */,
  {32'hbe3f1264, 32'hbf1e6e4c} /* (0, 21, 20) {real, imag} */,
  {32'hbd1ed97c, 32'h3db2b870} /* (0, 21, 19) {real, imag} */,
  {32'h3ed922de, 32'h3defb1ae} /* (0, 21, 18) {real, imag} */,
  {32'hbdde2b16, 32'hbd966295} /* (0, 21, 17) {real, imag} */,
  {32'hbdc536e2, 32'hbe0cdd56} /* (0, 21, 16) {real, imag} */,
  {32'hbd16fbdc, 32'h3e60963b} /* (0, 21, 15) {real, imag} */,
  {32'hbe01069c, 32'hbe9ac822} /* (0, 21, 14) {real, imag} */,
  {32'hbddd6290, 32'hbe697720} /* (0, 21, 13) {real, imag} */,
  {32'h3e5997b7, 32'hbe0c1200} /* (0, 21, 12) {real, imag} */,
  {32'hbe10e220, 32'h3f4bfbb0} /* (0, 21, 11) {real, imag} */,
  {32'h3d5891e0, 32'hbd04e3e0} /* (0, 21, 10) {real, imag} */,
  {32'hbd8379f0, 32'h3dba598a} /* (0, 21, 9) {real, imag} */,
  {32'h3e4d3e85, 32'hbeab0f0e} /* (0, 21, 8) {real, imag} */,
  {32'hbdb3ea35, 32'hbdadfd22} /* (0, 21, 7) {real, imag} */,
  {32'h3ead1b80, 32'hbe903f66} /* (0, 21, 6) {real, imag} */,
  {32'hbdaca0d0, 32'h3c2dc5e0} /* (0, 21, 5) {real, imag} */,
  {32'hbe7d3084, 32'h3e3e8708} /* (0, 21, 4) {real, imag} */,
  {32'hbe8cd5c8, 32'hbeab2fb0} /* (0, 21, 3) {real, imag} */,
  {32'h3e99aab3, 32'h3e0ab698} /* (0, 21, 2) {real, imag} */,
  {32'h3eb178fe, 32'hbcc35440} /* (0, 21, 1) {real, imag} */,
  {32'hbdba6690, 32'hbd01b194} /* (0, 21, 0) {real, imag} */,
  {32'h3e8eb132, 32'h3e541659} /* (0, 20, 31) {real, imag} */,
  {32'h3ea95892, 32'hbe3ea2dc} /* (0, 20, 30) {real, imag} */,
  {32'h3be04d40, 32'h3c5aa400} /* (0, 20, 29) {real, imag} */,
  {32'hbe090d53, 32'hbe92c8ac} /* (0, 20, 28) {real, imag} */,
  {32'hbe1a7e45, 32'h3ead2906} /* (0, 20, 27) {real, imag} */,
  {32'hbe4af0b4, 32'h3e14d2d4} /* (0, 20, 26) {real, imag} */,
  {32'h3e43e9cb, 32'hbeb11fae} /* (0, 20, 25) {real, imag} */,
  {32'h3c16a380, 32'h3ea39878} /* (0, 20, 24) {real, imag} */,
  {32'h3da2b5da, 32'h3d274ca4} /* (0, 20, 23) {real, imag} */,
  {32'h3e32803a, 32'h3e2946ec} /* (0, 20, 22) {real, imag} */,
  {32'hbee376d2, 32'hbd36d37d} /* (0, 20, 21) {real, imag} */,
  {32'h3e01db02, 32'hbe764178} /* (0, 20, 20) {real, imag} */,
  {32'h3e1d30c5, 32'h3e6c944c} /* (0, 20, 19) {real, imag} */,
  {32'hbe37dc10, 32'h3e9b09ea} /* (0, 20, 18) {real, imag} */,
  {32'h3d387988, 32'h3e7e05e2} /* (0, 20, 17) {real, imag} */,
  {32'hbdb6decc, 32'hbde7f565} /* (0, 20, 16) {real, imag} */,
  {32'hbde4950b, 32'hbe666601} /* (0, 20, 15) {real, imag} */,
  {32'h3e590713, 32'h3d89e298} /* (0, 20, 14) {real, imag} */,
  {32'h3ee955fa, 32'hbe1a2e1f} /* (0, 20, 13) {real, imag} */,
  {32'h3c40d330, 32'hbd638e80} /* (0, 20, 12) {real, imag} */,
  {32'h3e2ee37a, 32'h3dd03379} /* (0, 20, 11) {real, imag} */,
  {32'h3d5792e7, 32'h3c87b970} /* (0, 20, 10) {real, imag} */,
  {32'hbd42d440, 32'hbef317e6} /* (0, 20, 9) {real, imag} */,
  {32'hbe329a89, 32'hbe6e6bc2} /* (0, 20, 8) {real, imag} */,
  {32'h3e17d8c8, 32'h3e045798} /* (0, 20, 7) {real, imag} */,
  {32'hbdcd6beb, 32'h3e6afc59} /* (0, 20, 6) {real, imag} */,
  {32'hbe8cc4ce, 32'hbcff5c10} /* (0, 20, 5) {real, imag} */,
  {32'hbe7f7558, 32'h3d181770} /* (0, 20, 4) {real, imag} */,
  {32'hbdbf5527, 32'h3eaea198} /* (0, 20, 3) {real, imag} */,
  {32'hbdf76348, 32'h3e891bc9} /* (0, 20, 2) {real, imag} */,
  {32'h3e17eaae, 32'hbeefd661} /* (0, 20, 1) {real, imag} */,
  {32'h3cd6b808, 32'h3e95a892} /* (0, 20, 0) {real, imag} */,
  {32'h3e78e841, 32'hbd8f6b7a} /* (0, 19, 31) {real, imag} */,
  {32'h3ca7aac8, 32'h3e3d4474} /* (0, 19, 30) {real, imag} */,
  {32'h3da1bf94, 32'hbe08b5f2} /* (0, 19, 29) {real, imag} */,
  {32'h3cd4a6f0, 32'h3e894a27} /* (0, 19, 28) {real, imag} */,
  {32'h3d0ac577, 32'hbd201be2} /* (0, 19, 27) {real, imag} */,
  {32'h3d935c45, 32'h3e230dc8} /* (0, 19, 26) {real, imag} */,
  {32'hbeb15e52, 32'hbdff6773} /* (0, 19, 25) {real, imag} */,
  {32'h3ed633b8, 32'h3eaaf2ad} /* (0, 19, 24) {real, imag} */,
  {32'hbe032715, 32'hbed9868e} /* (0, 19, 23) {real, imag} */,
  {32'h3eeeaa25, 32'hbd070090} /* (0, 19, 22) {real, imag} */,
  {32'hbe674fca, 32'hbda4fbe2} /* (0, 19, 21) {real, imag} */,
  {32'hbcba666c, 32'hbd0ab2bc} /* (0, 19, 20) {real, imag} */,
  {32'h3e2ae4e4, 32'h3ddd25f4} /* (0, 19, 19) {real, imag} */,
  {32'hbe715950, 32'h3e51732c} /* (0, 19, 18) {real, imag} */,
  {32'h3e8931e8, 32'hbd053820} /* (0, 19, 17) {real, imag} */,
  {32'h3e29d8cc, 32'h3d73633e} /* (0, 19, 16) {real, imag} */,
  {32'hbdf82996, 32'hbe86075f} /* (0, 19, 15) {real, imag} */,
  {32'hbea299ff, 32'hbec431a4} /* (0, 19, 14) {real, imag} */,
  {32'hbe64ee0b, 32'hbd7a5cfc} /* (0, 19, 13) {real, imag} */,
  {32'hbd8d2450, 32'h3d5198c6} /* (0, 19, 12) {real, imag} */,
  {32'hbe58370b, 32'h3e4e7ddc} /* (0, 19, 11) {real, imag} */,
  {32'h3e6d362e, 32'h3e3c0318} /* (0, 19, 10) {real, imag} */,
  {32'h3d23fc20, 32'hbd204528} /* (0, 19, 9) {real, imag} */,
  {32'hbcfc21a8, 32'hbe55211e} /* (0, 19, 8) {real, imag} */,
  {32'h3e544ec2, 32'hbe51b25e} /* (0, 19, 7) {real, imag} */,
  {32'h3e5547a3, 32'h3e2184ae} /* (0, 19, 6) {real, imag} */,
  {32'hba052a00, 32'h3e2495a1} /* (0, 19, 5) {real, imag} */,
  {32'hbd9f4ee0, 32'h3ea9aa18} /* (0, 19, 4) {real, imag} */,
  {32'hbebb4432, 32'hbe6b22b4} /* (0, 19, 3) {real, imag} */,
  {32'h3f132189, 32'hbe6a3c26} /* (0, 19, 2) {real, imag} */,
  {32'hbdec0cf6, 32'h3ea4aa5b} /* (0, 19, 1) {real, imag} */,
  {32'hbed0aa9e, 32'hbe920454} /* (0, 19, 0) {real, imag} */,
  {32'hbeadba82, 32'hbeb069c2} /* (0, 18, 31) {real, imag} */,
  {32'hbe2f8be0, 32'h3e6bd1c5} /* (0, 18, 30) {real, imag} */,
  {32'h3e5fe07b, 32'h3e31b8f0} /* (0, 18, 29) {real, imag} */,
  {32'h3d491ffe, 32'hbe4211f3} /* (0, 18, 28) {real, imag} */,
  {32'hbdeaed0e, 32'h3eab82a8} /* (0, 18, 27) {real, imag} */,
  {32'h3e096dd9, 32'hbd215c56} /* (0, 18, 26) {real, imag} */,
  {32'h3e89e1c8, 32'h3e39f2ac} /* (0, 18, 25) {real, imag} */,
  {32'h3d91924d, 32'h3e96d925} /* (0, 18, 24) {real, imag} */,
  {32'hbe9cd7b3, 32'h3e56e5a6} /* (0, 18, 23) {real, imag} */,
  {32'hbe5480df, 32'hbe4a639c} /* (0, 18, 22) {real, imag} */,
  {32'h3eb951a8, 32'hbdca1988} /* (0, 18, 21) {real, imag} */,
  {32'h3ea77c65, 32'hbdc319b0} /* (0, 18, 20) {real, imag} */,
  {32'h3e39f2cb, 32'h3e103641} /* (0, 18, 19) {real, imag} */,
  {32'h3dc1fdda, 32'hbbc9b6a0} /* (0, 18, 18) {real, imag} */,
  {32'hbd87ce5a, 32'h3e3e04d2} /* (0, 18, 17) {real, imag} */,
  {32'h3ceacbd0, 32'h3e8dfeda} /* (0, 18, 16) {real, imag} */,
  {32'hbde0cec8, 32'h3e014057} /* (0, 18, 15) {real, imag} */,
  {32'h3e37c2e0, 32'hbe8ec21c} /* (0, 18, 14) {real, imag} */,
  {32'hbd110ed8, 32'h3d45e6d1} /* (0, 18, 13) {real, imag} */,
  {32'h3e6677ec, 32'hbd4a7e48} /* (0, 18, 12) {real, imag} */,
  {32'h3de850ce, 32'hbdd5941a} /* (0, 18, 11) {real, imag} */,
  {32'hbdc903ba, 32'h3f23fa4c} /* (0, 18, 10) {real, imag} */,
  {32'h3e97543b, 32'hbe472560} /* (0, 18, 9) {real, imag} */,
  {32'h3d2bb6bc, 32'h3e1baf7f} /* (0, 18, 8) {real, imag} */,
  {32'hbda873ea, 32'h3e8dfeb8} /* (0, 18, 7) {real, imag} */,
  {32'hbe0fd1b0, 32'hbde7df2a} /* (0, 18, 6) {real, imag} */,
  {32'h3d8d82e9, 32'h3e90bf2f} /* (0, 18, 5) {real, imag} */,
  {32'h3e6568f4, 32'hbe664bd6} /* (0, 18, 4) {real, imag} */,
  {32'hbdfe843b, 32'hbd899d90} /* (0, 18, 3) {real, imag} */,
  {32'hbecf2ede, 32'h3a7a4140} /* (0, 18, 2) {real, imag} */,
  {32'hbd5dee9d, 32'hbaece880} /* (0, 18, 1) {real, imag} */,
  {32'hbd173234, 32'hbe282256} /* (0, 18, 0) {real, imag} */,
  {32'hbe01b70a, 32'h3e0854c5} /* (0, 17, 31) {real, imag} */,
  {32'h3ea2d3ac, 32'hbe9a5886} /* (0, 17, 30) {real, imag} */,
  {32'hbd9f4d2c, 32'h3d70c0e0} /* (0, 17, 29) {real, imag} */,
  {32'h3d200d95, 32'h3c535ac8} /* (0, 17, 28) {real, imag} */,
  {32'h3cc64c90, 32'h3c6e2a94} /* (0, 17, 27) {real, imag} */,
  {32'hbe4c0428, 32'hbdad6152} /* (0, 17, 26) {real, imag} */,
  {32'h3e3a15dd, 32'h3dfbe8f0} /* (0, 17, 25) {real, imag} */,
  {32'hbd902eea, 32'h3e603b9c} /* (0, 17, 24) {real, imag} */,
  {32'hbe2f5d75, 32'h3d9eb344} /* (0, 17, 23) {real, imag} */,
  {32'h3e98ebc2, 32'h3d952545} /* (0, 17, 22) {real, imag} */,
  {32'hbe0598f7, 32'hbd317698} /* (0, 17, 21) {real, imag} */,
  {32'hbe1926db, 32'h3ea9051f} /* (0, 17, 20) {real, imag} */,
  {32'h3e767076, 32'hbe4127a4} /* (0, 17, 19) {real, imag} */,
  {32'hbcd18498, 32'h3dc0b6e1} /* (0, 17, 18) {real, imag} */,
  {32'hbdff0f10, 32'h3c52ef60} /* (0, 17, 17) {real, imag} */,
  {32'hbe3881d8, 32'h3d18aabf} /* (0, 17, 16) {real, imag} */,
  {32'h3e617661, 32'h3c4b38f0} /* (0, 17, 15) {real, imag} */,
  {32'h3e3e0e12, 32'h3e41f5f7} /* (0, 17, 14) {real, imag} */,
  {32'hbe5bcc14, 32'hbe6fb84e} /* (0, 17, 13) {real, imag} */,
  {32'hbdee8ea6, 32'h3e8d7cc4} /* (0, 17, 12) {real, imag} */,
  {32'hbe0b652e, 32'hbe86a54a} /* (0, 17, 11) {real, imag} */,
  {32'hbd82f204, 32'h3cee853c} /* (0, 17, 10) {real, imag} */,
  {32'h3e5813b7, 32'h3e64c010} /* (0, 17, 9) {real, imag} */,
  {32'hbda9cbb0, 32'hbd5e1f86} /* (0, 17, 8) {real, imag} */,
  {32'h3c4e0710, 32'hbbad8780} /* (0, 17, 7) {real, imag} */,
  {32'h3d49092c, 32'hbe12264a} /* (0, 17, 6) {real, imag} */,
  {32'h3dbdcdc2, 32'hbdb78610} /* (0, 17, 5) {real, imag} */,
  {32'hbe0848c6, 32'hbd8b5424} /* (0, 17, 4) {real, imag} */,
  {32'h3d9f3e45, 32'h3c0ec9d0} /* (0, 17, 3) {real, imag} */,
  {32'hbd224610, 32'hbed6b678} /* (0, 17, 2) {real, imag} */,
  {32'h3dc7ee00, 32'h3ea95790} /* (0, 17, 1) {real, imag} */,
  {32'hbbdcd958, 32'hbda991a8} /* (0, 17, 0) {real, imag} */,
  {32'hbd4c849f, 32'h3cbc5e48} /* (0, 16, 31) {real, imag} */,
  {32'h3dad4e08, 32'h3daf5ef0} /* (0, 16, 30) {real, imag} */,
  {32'hbdddcefa, 32'hbc9ff684} /* (0, 16, 29) {real, imag} */,
  {32'h3b943478, 32'h3d568590} /* (0, 16, 28) {real, imag} */,
  {32'hbd0c2900, 32'hba0d8e00} /* (0, 16, 27) {real, imag} */,
  {32'hbd9444f2, 32'h3ce9e3c8} /* (0, 16, 26) {real, imag} */,
  {32'hbc2c0010, 32'h3eaec518} /* (0, 16, 25) {real, imag} */,
  {32'h3df2689c, 32'hbd4a4df4} /* (0, 16, 24) {real, imag} */,
  {32'h3ea58d3c, 32'hbd071eba} /* (0, 16, 23) {real, imag} */,
  {32'hbdab123b, 32'h3de2eccd} /* (0, 16, 22) {real, imag} */,
  {32'h3cba52fa, 32'h3dc05df8} /* (0, 16, 21) {real, imag} */,
  {32'hbe91ef80, 32'h3dfb6fd8} /* (0, 16, 20) {real, imag} */,
  {32'hbc81d956, 32'h3ee00c18} /* (0, 16, 19) {real, imag} */,
  {32'hbda57574, 32'h3d925b1d} /* (0, 16, 18) {real, imag} */,
  {32'hbce1921a, 32'h3e0ac1e1} /* (0, 16, 17) {real, imag} */,
  {32'hbba186f8, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hbce1921a, 32'hbe0ac1e1} /* (0, 16, 15) {real, imag} */,
  {32'hbda57574, 32'hbd925b1d} /* (0, 16, 14) {real, imag} */,
  {32'hbc81d956, 32'hbee00c18} /* (0, 16, 13) {real, imag} */,
  {32'hbe91ef80, 32'hbdfb6fd8} /* (0, 16, 12) {real, imag} */,
  {32'h3cba52fa, 32'hbdc05df8} /* (0, 16, 11) {real, imag} */,
  {32'hbdab123b, 32'hbde2eccd} /* (0, 16, 10) {real, imag} */,
  {32'h3ea58d3c, 32'h3d071eba} /* (0, 16, 9) {real, imag} */,
  {32'h3df2689c, 32'h3d4a4df4} /* (0, 16, 8) {real, imag} */,
  {32'hbc2c0010, 32'hbeaec518} /* (0, 16, 7) {real, imag} */,
  {32'hbd9444f2, 32'hbce9e3c8} /* (0, 16, 6) {real, imag} */,
  {32'hbd0c2900, 32'h3a0d8e00} /* (0, 16, 5) {real, imag} */,
  {32'h3b943478, 32'hbd568590} /* (0, 16, 4) {real, imag} */,
  {32'hbdddcefa, 32'h3c9ff684} /* (0, 16, 3) {real, imag} */,
  {32'h3dad4e08, 32'hbdaf5ef0} /* (0, 16, 2) {real, imag} */,
  {32'hbd4c849f, 32'hbcbc5e48} /* (0, 16, 1) {real, imag} */,
  {32'h3ef765c6, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h3dc7ee00, 32'hbea95790} /* (0, 15, 31) {real, imag} */,
  {32'hbd224610, 32'h3ed6b678} /* (0, 15, 30) {real, imag} */,
  {32'h3d9f3e45, 32'hbc0ec9d0} /* (0, 15, 29) {real, imag} */,
  {32'hbe0848c6, 32'h3d8b5424} /* (0, 15, 28) {real, imag} */,
  {32'h3dbdcdc2, 32'h3db78610} /* (0, 15, 27) {real, imag} */,
  {32'h3d49092c, 32'h3e12264a} /* (0, 15, 26) {real, imag} */,
  {32'h3c4e0710, 32'h3bad8780} /* (0, 15, 25) {real, imag} */,
  {32'hbda9cbb0, 32'h3d5e1f86} /* (0, 15, 24) {real, imag} */,
  {32'h3e5813b7, 32'hbe64c010} /* (0, 15, 23) {real, imag} */,
  {32'hbd82f204, 32'hbcee853c} /* (0, 15, 22) {real, imag} */,
  {32'hbe0b652e, 32'h3e86a54a} /* (0, 15, 21) {real, imag} */,
  {32'hbdee8ea6, 32'hbe8d7cc4} /* (0, 15, 20) {real, imag} */,
  {32'hbe5bcc14, 32'h3e6fb84e} /* (0, 15, 19) {real, imag} */,
  {32'h3e3e0e12, 32'hbe41f5f7} /* (0, 15, 18) {real, imag} */,
  {32'h3e617661, 32'hbc4b38f0} /* (0, 15, 17) {real, imag} */,
  {32'hbe3881d8, 32'hbd18aabf} /* (0, 15, 16) {real, imag} */,
  {32'hbdff0f10, 32'hbc52ef60} /* (0, 15, 15) {real, imag} */,
  {32'hbcd18498, 32'hbdc0b6e1} /* (0, 15, 14) {real, imag} */,
  {32'h3e767076, 32'h3e4127a4} /* (0, 15, 13) {real, imag} */,
  {32'hbe1926db, 32'hbea9051f} /* (0, 15, 12) {real, imag} */,
  {32'hbe0598f7, 32'h3d317698} /* (0, 15, 11) {real, imag} */,
  {32'h3e98ebc2, 32'hbd952545} /* (0, 15, 10) {real, imag} */,
  {32'hbe2f5d75, 32'hbd9eb344} /* (0, 15, 9) {real, imag} */,
  {32'hbd902eea, 32'hbe603b9c} /* (0, 15, 8) {real, imag} */,
  {32'h3e3a15dd, 32'hbdfbe8f0} /* (0, 15, 7) {real, imag} */,
  {32'hbe4c0428, 32'h3dad6152} /* (0, 15, 6) {real, imag} */,
  {32'h3cc64c90, 32'hbc6e2a94} /* (0, 15, 5) {real, imag} */,
  {32'h3d200d95, 32'hbc535ac8} /* (0, 15, 4) {real, imag} */,
  {32'hbd9f4d2c, 32'hbd70c0e0} /* (0, 15, 3) {real, imag} */,
  {32'h3ea2d3ac, 32'h3e9a5886} /* (0, 15, 2) {real, imag} */,
  {32'hbe01b70a, 32'hbe0854c5} /* (0, 15, 1) {real, imag} */,
  {32'hbbdcd958, 32'h3da991a8} /* (0, 15, 0) {real, imag} */,
  {32'hbd5dee9d, 32'h3aece880} /* (0, 14, 31) {real, imag} */,
  {32'hbecf2ede, 32'hba7a4140} /* (0, 14, 30) {real, imag} */,
  {32'hbdfe843b, 32'h3d899d90} /* (0, 14, 29) {real, imag} */,
  {32'h3e6568f4, 32'h3e664bd6} /* (0, 14, 28) {real, imag} */,
  {32'h3d8d82e9, 32'hbe90bf2f} /* (0, 14, 27) {real, imag} */,
  {32'hbe0fd1b0, 32'h3de7df2a} /* (0, 14, 26) {real, imag} */,
  {32'hbda873ea, 32'hbe8dfeb8} /* (0, 14, 25) {real, imag} */,
  {32'h3d2bb6bc, 32'hbe1baf7f} /* (0, 14, 24) {real, imag} */,
  {32'h3e97543b, 32'h3e472560} /* (0, 14, 23) {real, imag} */,
  {32'hbdc903ba, 32'hbf23fa4c} /* (0, 14, 22) {real, imag} */,
  {32'h3de850ce, 32'h3dd5941a} /* (0, 14, 21) {real, imag} */,
  {32'h3e6677ec, 32'h3d4a7e48} /* (0, 14, 20) {real, imag} */,
  {32'hbd110ed8, 32'hbd45e6d1} /* (0, 14, 19) {real, imag} */,
  {32'h3e37c2e0, 32'h3e8ec21c} /* (0, 14, 18) {real, imag} */,
  {32'hbde0cec8, 32'hbe014057} /* (0, 14, 17) {real, imag} */,
  {32'h3ceacbd0, 32'hbe8dfeda} /* (0, 14, 16) {real, imag} */,
  {32'hbd87ce5a, 32'hbe3e04d2} /* (0, 14, 15) {real, imag} */,
  {32'h3dc1fdda, 32'h3bc9b6a0} /* (0, 14, 14) {real, imag} */,
  {32'h3e39f2cb, 32'hbe103641} /* (0, 14, 13) {real, imag} */,
  {32'h3ea77c65, 32'h3dc319b0} /* (0, 14, 12) {real, imag} */,
  {32'h3eb951a8, 32'h3dca1988} /* (0, 14, 11) {real, imag} */,
  {32'hbe5480df, 32'h3e4a639c} /* (0, 14, 10) {real, imag} */,
  {32'hbe9cd7b3, 32'hbe56e5a6} /* (0, 14, 9) {real, imag} */,
  {32'h3d91924d, 32'hbe96d925} /* (0, 14, 8) {real, imag} */,
  {32'h3e89e1c8, 32'hbe39f2ac} /* (0, 14, 7) {real, imag} */,
  {32'h3e096dd9, 32'h3d215c56} /* (0, 14, 6) {real, imag} */,
  {32'hbdeaed0e, 32'hbeab82a8} /* (0, 14, 5) {real, imag} */,
  {32'h3d491ffe, 32'h3e4211f3} /* (0, 14, 4) {real, imag} */,
  {32'h3e5fe07b, 32'hbe31b8f0} /* (0, 14, 3) {real, imag} */,
  {32'hbe2f8be0, 32'hbe6bd1c5} /* (0, 14, 2) {real, imag} */,
  {32'hbeadba82, 32'h3eb069c2} /* (0, 14, 1) {real, imag} */,
  {32'hbd173234, 32'h3e282256} /* (0, 14, 0) {real, imag} */,
  {32'hbdec0cf6, 32'hbea4aa5b} /* (0, 13, 31) {real, imag} */,
  {32'h3f132189, 32'h3e6a3c26} /* (0, 13, 30) {real, imag} */,
  {32'hbebb4432, 32'h3e6b22b4} /* (0, 13, 29) {real, imag} */,
  {32'hbd9f4ee0, 32'hbea9aa18} /* (0, 13, 28) {real, imag} */,
  {32'hba052a00, 32'hbe2495a1} /* (0, 13, 27) {real, imag} */,
  {32'h3e5547a3, 32'hbe2184ae} /* (0, 13, 26) {real, imag} */,
  {32'h3e544ec2, 32'h3e51b25e} /* (0, 13, 25) {real, imag} */,
  {32'hbcfc21a8, 32'h3e55211e} /* (0, 13, 24) {real, imag} */,
  {32'h3d23fc20, 32'h3d204528} /* (0, 13, 23) {real, imag} */,
  {32'h3e6d362e, 32'hbe3c0318} /* (0, 13, 22) {real, imag} */,
  {32'hbe58370b, 32'hbe4e7ddc} /* (0, 13, 21) {real, imag} */,
  {32'hbd8d2450, 32'hbd5198c6} /* (0, 13, 20) {real, imag} */,
  {32'hbe64ee0b, 32'h3d7a5cfc} /* (0, 13, 19) {real, imag} */,
  {32'hbea299ff, 32'h3ec431a4} /* (0, 13, 18) {real, imag} */,
  {32'hbdf82996, 32'h3e86075f} /* (0, 13, 17) {real, imag} */,
  {32'h3e29d8cc, 32'hbd73633e} /* (0, 13, 16) {real, imag} */,
  {32'h3e8931e8, 32'h3d053820} /* (0, 13, 15) {real, imag} */,
  {32'hbe715950, 32'hbe51732c} /* (0, 13, 14) {real, imag} */,
  {32'h3e2ae4e4, 32'hbddd25f4} /* (0, 13, 13) {real, imag} */,
  {32'hbcba666c, 32'h3d0ab2bc} /* (0, 13, 12) {real, imag} */,
  {32'hbe674fca, 32'h3da4fbe2} /* (0, 13, 11) {real, imag} */,
  {32'h3eeeaa25, 32'h3d070090} /* (0, 13, 10) {real, imag} */,
  {32'hbe032715, 32'h3ed9868e} /* (0, 13, 9) {real, imag} */,
  {32'h3ed633b8, 32'hbeaaf2ad} /* (0, 13, 8) {real, imag} */,
  {32'hbeb15e52, 32'h3dff6773} /* (0, 13, 7) {real, imag} */,
  {32'h3d935c45, 32'hbe230dc8} /* (0, 13, 6) {real, imag} */,
  {32'h3d0ac577, 32'h3d201be2} /* (0, 13, 5) {real, imag} */,
  {32'h3cd4a6f0, 32'hbe894a27} /* (0, 13, 4) {real, imag} */,
  {32'h3da1bf94, 32'h3e08b5f2} /* (0, 13, 3) {real, imag} */,
  {32'h3ca7aac8, 32'hbe3d4474} /* (0, 13, 2) {real, imag} */,
  {32'h3e78e841, 32'h3d8f6b7a} /* (0, 13, 1) {real, imag} */,
  {32'hbed0aa9e, 32'h3e920454} /* (0, 13, 0) {real, imag} */,
  {32'h3e17eaae, 32'h3eefd661} /* (0, 12, 31) {real, imag} */,
  {32'hbdf76348, 32'hbe891bc9} /* (0, 12, 30) {real, imag} */,
  {32'hbdbf5527, 32'hbeaea198} /* (0, 12, 29) {real, imag} */,
  {32'hbe7f7558, 32'hbd181770} /* (0, 12, 28) {real, imag} */,
  {32'hbe8cc4ce, 32'h3cff5c10} /* (0, 12, 27) {real, imag} */,
  {32'hbdcd6beb, 32'hbe6afc59} /* (0, 12, 26) {real, imag} */,
  {32'h3e17d8c8, 32'hbe045798} /* (0, 12, 25) {real, imag} */,
  {32'hbe329a89, 32'h3e6e6bc2} /* (0, 12, 24) {real, imag} */,
  {32'hbd42d440, 32'h3ef317e6} /* (0, 12, 23) {real, imag} */,
  {32'h3d5792e7, 32'hbc87b970} /* (0, 12, 22) {real, imag} */,
  {32'h3e2ee37a, 32'hbdd03379} /* (0, 12, 21) {real, imag} */,
  {32'h3c40d330, 32'h3d638e80} /* (0, 12, 20) {real, imag} */,
  {32'h3ee955fa, 32'h3e1a2e1f} /* (0, 12, 19) {real, imag} */,
  {32'h3e590713, 32'hbd89e298} /* (0, 12, 18) {real, imag} */,
  {32'hbde4950b, 32'h3e666601} /* (0, 12, 17) {real, imag} */,
  {32'hbdb6decc, 32'h3de7f565} /* (0, 12, 16) {real, imag} */,
  {32'h3d387988, 32'hbe7e05e2} /* (0, 12, 15) {real, imag} */,
  {32'hbe37dc10, 32'hbe9b09ea} /* (0, 12, 14) {real, imag} */,
  {32'h3e1d30c5, 32'hbe6c944c} /* (0, 12, 13) {real, imag} */,
  {32'h3e01db02, 32'h3e764178} /* (0, 12, 12) {real, imag} */,
  {32'hbee376d2, 32'h3d36d37d} /* (0, 12, 11) {real, imag} */,
  {32'h3e32803a, 32'hbe2946ec} /* (0, 12, 10) {real, imag} */,
  {32'h3da2b5da, 32'hbd274ca4} /* (0, 12, 9) {real, imag} */,
  {32'h3c16a380, 32'hbea39878} /* (0, 12, 8) {real, imag} */,
  {32'h3e43e9cb, 32'h3eb11fae} /* (0, 12, 7) {real, imag} */,
  {32'hbe4af0b4, 32'hbe14d2d4} /* (0, 12, 6) {real, imag} */,
  {32'hbe1a7e45, 32'hbead2906} /* (0, 12, 5) {real, imag} */,
  {32'hbe090d53, 32'h3e92c8ac} /* (0, 12, 4) {real, imag} */,
  {32'h3be04d40, 32'hbc5aa400} /* (0, 12, 3) {real, imag} */,
  {32'h3ea95892, 32'h3e3ea2dc} /* (0, 12, 2) {real, imag} */,
  {32'h3e8eb132, 32'hbe541659} /* (0, 12, 1) {real, imag} */,
  {32'h3cd6b808, 32'hbe95a892} /* (0, 12, 0) {real, imag} */,
  {32'h3eb178fe, 32'h3cc35440} /* (0, 11, 31) {real, imag} */,
  {32'h3e99aab3, 32'hbe0ab698} /* (0, 11, 30) {real, imag} */,
  {32'hbe8cd5c8, 32'h3eab2fb0} /* (0, 11, 29) {real, imag} */,
  {32'hbe7d3084, 32'hbe3e8708} /* (0, 11, 28) {real, imag} */,
  {32'hbdaca0d0, 32'hbc2dc5e0} /* (0, 11, 27) {real, imag} */,
  {32'h3ead1b80, 32'h3e903f66} /* (0, 11, 26) {real, imag} */,
  {32'hbdb3ea35, 32'h3dadfd22} /* (0, 11, 25) {real, imag} */,
  {32'h3e4d3e85, 32'h3eab0f0e} /* (0, 11, 24) {real, imag} */,
  {32'hbd8379f0, 32'hbdba598a} /* (0, 11, 23) {real, imag} */,
  {32'h3d5891e0, 32'h3d04e3e0} /* (0, 11, 22) {real, imag} */,
  {32'hbe10e220, 32'hbf4bfbb0} /* (0, 11, 21) {real, imag} */,
  {32'h3e5997b7, 32'h3e0c1200} /* (0, 11, 20) {real, imag} */,
  {32'hbddd6290, 32'h3e697720} /* (0, 11, 19) {real, imag} */,
  {32'hbe01069c, 32'h3e9ac822} /* (0, 11, 18) {real, imag} */,
  {32'hbd16fbdc, 32'hbe60963b} /* (0, 11, 17) {real, imag} */,
  {32'hbdc536e2, 32'h3e0cdd56} /* (0, 11, 16) {real, imag} */,
  {32'hbdde2b16, 32'h3d966295} /* (0, 11, 15) {real, imag} */,
  {32'h3ed922de, 32'hbdefb1ae} /* (0, 11, 14) {real, imag} */,
  {32'hbd1ed97c, 32'hbdb2b870} /* (0, 11, 13) {real, imag} */,
  {32'hbe3f1264, 32'h3f1e6e4c} /* (0, 11, 12) {real, imag} */,
  {32'h3e93d3dd, 32'hbdf88aaf} /* (0, 11, 11) {real, imag} */,
  {32'hbf5bcabc, 32'hbe27c818} /* (0, 11, 10) {real, imag} */,
  {32'h3dec915e, 32'h3da091b0} /* (0, 11, 9) {real, imag} */,
  {32'hbd94bec8, 32'h3e6c6655} /* (0, 11, 8) {real, imag} */,
  {32'h3e04aa46, 32'hbd0404ad} /* (0, 11, 7) {real, imag} */,
  {32'h3dd2335c, 32'hbdbf15e8} /* (0, 11, 6) {real, imag} */,
  {32'hbebc1c0e, 32'h3e5ca805} /* (0, 11, 5) {real, imag} */,
  {32'hbde18ee6, 32'hbeab2984} /* (0, 11, 4) {real, imag} */,
  {32'h3e539569, 32'hbda46088} /* (0, 11, 3) {real, imag} */,
  {32'h3dd5c0b4, 32'hbec0fcdd} /* (0, 11, 2) {real, imag} */,
  {32'h3e06507f, 32'hbe027d23} /* (0, 11, 1) {real, imag} */,
  {32'hbdba6690, 32'h3d01b194} /* (0, 11, 0) {real, imag} */,
  {32'hbd083304, 32'hbda16f7e} /* (0, 10, 31) {real, imag} */,
  {32'hbcde3410, 32'h3e882b57} /* (0, 10, 30) {real, imag} */,
  {32'hbe09faa3, 32'hbdd393fd} /* (0, 10, 29) {real, imag} */,
  {32'hbe997e51, 32'hbe94e99f} /* (0, 10, 28) {real, imag} */,
  {32'h3ef420ec, 32'h3e216d08} /* (0, 10, 27) {real, imag} */,
  {32'hbd1dd44c, 32'h3eae7ede} /* (0, 10, 26) {real, imag} */,
  {32'h3c97c970, 32'hbdea99db} /* (0, 10, 25) {real, imag} */,
  {32'h3ee739a8, 32'hbe8964e2} /* (0, 10, 24) {real, imag} */,
  {32'h3e588486, 32'hbebb5b48} /* (0, 10, 23) {real, imag} */,
  {32'hbe10570f, 32'hbe4502aa} /* (0, 10, 22) {real, imag} */,
  {32'h3dcfbbfc, 32'hbe603e80} /* (0, 10, 21) {real, imag} */,
  {32'h3dcd83c4, 32'h3e74f3b2} /* (0, 10, 20) {real, imag} */,
  {32'h3e1af9f8, 32'h3ca74830} /* (0, 10, 19) {real, imag} */,
  {32'hbe312066, 32'hbd6eb666} /* (0, 10, 18) {real, imag} */,
  {32'h3ccd43ec, 32'h3b0fbd00} /* (0, 10, 17) {real, imag} */,
  {32'h3d80c70a, 32'hbe2d92bc} /* (0, 10, 16) {real, imag} */,
  {32'hbdfcda8c, 32'h3de25f92} /* (0, 10, 15) {real, imag} */,
  {32'h3e30295c, 32'hbe0f237e} /* (0, 10, 14) {real, imag} */,
  {32'h3eb29ef4, 32'hbd8b6914} /* (0, 10, 13) {real, imag} */,
  {32'hbedc6ba2, 32'hbee8ca45} /* (0, 10, 12) {real, imag} */,
  {32'h3e2645f5, 32'hbdaf4698} /* (0, 10, 11) {real, imag} */,
  {32'h3e865f62, 32'hbdfea096} /* (0, 10, 10) {real, imag} */,
  {32'h3d5080fa, 32'hbeeaf5ae} /* (0, 10, 9) {real, imag} */,
  {32'h3e18f172, 32'hbdcffbb4} /* (0, 10, 8) {real, imag} */,
  {32'h3e0d32b6, 32'hbdb87fa8} /* (0, 10, 7) {real, imag} */,
  {32'hbd746e2c, 32'hbce63958} /* (0, 10, 6) {real, imag} */,
  {32'hbdd6b508, 32'hbc334c28} /* (0, 10, 5) {real, imag} */,
  {32'h3e085a68, 32'hbe8568ba} /* (0, 10, 4) {real, imag} */,
  {32'hbd48e058, 32'h3da6387b} /* (0, 10, 3) {real, imag} */,
  {32'h3f17403c, 32'h3f3ef3a2} /* (0, 10, 2) {real, imag} */,
  {32'hbf1a8a3c, 32'hbc27da90} /* (0, 10, 1) {real, imag} */,
  {32'h3ded1ed8, 32'hbd92ae52} /* (0, 10, 0) {real, imag} */,
  {32'h3c5c3c28, 32'hbe0d45cf} /* (0, 9, 31) {real, imag} */,
  {32'h3f1e3a69, 32'h3f02174f} /* (0, 9, 30) {real, imag} */,
  {32'hbf2dc512, 32'h3ec1766c} /* (0, 9, 29) {real, imag} */,
  {32'hbecee360, 32'hbf0cf41b} /* (0, 9, 28) {real, imag} */,
  {32'h3e6cf843, 32'hbca73028} /* (0, 9, 27) {real, imag} */,
  {32'hbcf691a0, 32'hbe5ec45f} /* (0, 9, 26) {real, imag} */,
  {32'h3e9bcfd6, 32'hbc94dd58} /* (0, 9, 25) {real, imag} */,
  {32'h3e2f73ce, 32'hbea8cbb5} /* (0, 9, 24) {real, imag} */,
  {32'h3d491348, 32'h3dd6c3f6} /* (0, 9, 23) {real, imag} */,
  {32'hbb284880, 32'h3ea560ce} /* (0, 9, 22) {real, imag} */,
  {32'hbc961320, 32'h3cf1d198} /* (0, 9, 21) {real, imag} */,
  {32'h3ce7ee98, 32'hbe445ea4} /* (0, 9, 20) {real, imag} */,
  {32'h3e45325c, 32'h3c242578} /* (0, 9, 19) {real, imag} */,
  {32'hbe426d7d, 32'h3dd1c736} /* (0, 9, 18) {real, imag} */,
  {32'hbde5454f, 32'hbe4a01d3} /* (0, 9, 17) {real, imag} */,
  {32'h3e18bb41, 32'hbc008c40} /* (0, 9, 16) {real, imag} */,
  {32'h3d4d0d20, 32'hbd9ec486} /* (0, 9, 15) {real, imag} */,
  {32'hbe87b8ca, 32'h3b2b0560} /* (0, 9, 14) {real, imag} */,
  {32'hbd737254, 32'h3c54f2a8} /* (0, 9, 13) {real, imag} */,
  {32'h3e9a2ed5, 32'h3e887a14} /* (0, 9, 12) {real, imag} */,
  {32'hbeece180, 32'h3be24fc0} /* (0, 9, 11) {real, imag} */,
  {32'h3e7b4aa0, 32'h3e94dc92} /* (0, 9, 10) {real, imag} */,
  {32'hbe5bfd9e, 32'hbd863f86} /* (0, 9, 9) {real, imag} */,
  {32'hbd5ff710, 32'h3ec85cc8} /* (0, 9, 8) {real, imag} */,
  {32'h3dd6d538, 32'h3d41c0f2} /* (0, 9, 7) {real, imag} */,
  {32'h3ea15090, 32'h3d2aa520} /* (0, 9, 6) {real, imag} */,
  {32'hbcd8159a, 32'h3d8fc468} /* (0, 9, 5) {real, imag} */,
  {32'hbd991e32, 32'h3e82cb4f} /* (0, 9, 4) {real, imag} */,
  {32'hbd62ccbc, 32'hbeb84dc6} /* (0, 9, 3) {real, imag} */,
  {32'h3d3e5a24, 32'h3ccc68c0} /* (0, 9, 2) {real, imag} */,
  {32'hbf1d2422, 32'h3e07ce90} /* (0, 9, 1) {real, imag} */,
  {32'hbecf06c5, 32'hbe08554c} /* (0, 9, 0) {real, imag} */,
  {32'h3e4c7b92, 32'h3f0850e1} /* (0, 8, 31) {real, imag} */,
  {32'hbf864771, 32'hbe869517} /* (0, 8, 30) {real, imag} */,
  {32'hbcbcf3d8, 32'hbe1037e1} /* (0, 8, 29) {real, imag} */,
  {32'h3ef610dc, 32'hbe16e9e6} /* (0, 8, 28) {real, imag} */,
  {32'hbe00034a, 32'hbe2e6ea0} /* (0, 8, 27) {real, imag} */,
  {32'h3e2eaff6, 32'h3d9deacc} /* (0, 8, 26) {real, imag} */,
  {32'h3e8b3d56, 32'hbeb9ac7d} /* (0, 8, 25) {real, imag} */,
  {32'hbefcc5e2, 32'h3e3510ec} /* (0, 8, 24) {real, imag} */,
  {32'h3ebc6d8b, 32'hbe0b0487} /* (0, 8, 23) {real, imag} */,
  {32'hbe7ce8e5, 32'hbee69015} /* (0, 8, 22) {real, imag} */,
  {32'hbe29e3f4, 32'h3eba7491} /* (0, 8, 21) {real, imag} */,
  {32'hbe3f7d6b, 32'hbd3ea540} /* (0, 8, 20) {real, imag} */,
  {32'h3e687837, 32'h3e21c36d} /* (0, 8, 19) {real, imag} */,
  {32'h3ead80d0, 32'hbe0ca485} /* (0, 8, 18) {real, imag} */,
  {32'hbdc98d65, 32'hbd947032} /* (0, 8, 17) {real, imag} */,
  {32'hbcb1fc00, 32'hbeb5419e} /* (0, 8, 16) {real, imag} */,
  {32'h3dd755f0, 32'h3ccc52b0} /* (0, 8, 15) {real, imag} */,
  {32'h3e5c36e6, 32'h3ed2eba7} /* (0, 8, 14) {real, imag} */,
  {32'hbdc350fc, 32'h3e8e22ae} /* (0, 8, 13) {real, imag} */,
  {32'hbe35ab09, 32'hbe2b1723} /* (0, 8, 12) {real, imag} */,
  {32'h3e90954c, 32'hbe4322b9} /* (0, 8, 11) {real, imag} */,
  {32'hbeb63392, 32'h3db29500} /* (0, 8, 10) {real, imag} */,
  {32'hbd8960bc, 32'hbd019d68} /* (0, 8, 9) {real, imag} */,
  {32'h3de2c7ba, 32'hbcd03f30} /* (0, 8, 8) {real, imag} */,
  {32'h3e68aebc, 32'h3ebc7027} /* (0, 8, 7) {real, imag} */,
  {32'hbea76a7e, 32'hbe849026} /* (0, 8, 6) {real, imag} */,
  {32'h3e7d9973, 32'hbe5d3c6a} /* (0, 8, 5) {real, imag} */,
  {32'h3d9dca6a, 32'h3d93c4b8} /* (0, 8, 4) {real, imag} */,
  {32'hbf01de38, 32'h3e047694} /* (0, 8, 3) {real, imag} */,
  {32'hbf095349, 32'h3e099336} /* (0, 8, 2) {real, imag} */,
  {32'h3d1c3980, 32'h3f215289} /* (0, 8, 1) {real, imag} */,
  {32'h3f31299e, 32'h3f15be20} /* (0, 8, 0) {real, imag} */,
  {32'hbe228002, 32'h3e9cad96} /* (0, 7, 31) {real, imag} */,
  {32'h3eb5eefe, 32'h39fe4400} /* (0, 7, 30) {real, imag} */,
  {32'hbe77c858, 32'h3f08692d} /* (0, 7, 29) {real, imag} */,
  {32'h3e95bab6, 32'h3ed9c31b} /* (0, 7, 28) {real, imag} */,
  {32'hbe252ca6, 32'hbdc39573} /* (0, 7, 27) {real, imag} */,
  {32'hbe2d4f6c, 32'h3cddc930} /* (0, 7, 26) {real, imag} */,
  {32'h3dc9718e, 32'hbc858ea8} /* (0, 7, 25) {real, imag} */,
  {32'h3e08ba00, 32'hbe15ea24} /* (0, 7, 24) {real, imag} */,
  {32'hbd6621b4, 32'hbc8ceee0} /* (0, 7, 23) {real, imag} */,
  {32'h3ddc391c, 32'hbe38618f} /* (0, 7, 22) {real, imag} */,
  {32'h3e40076c, 32'hbcaf30f0} /* (0, 7, 21) {real, imag} */,
  {32'h39a3a800, 32'hbd50d9da} /* (0, 7, 20) {real, imag} */,
  {32'hbc2127e0, 32'h3e55de2a} /* (0, 7, 19) {real, imag} */,
  {32'hbe8ec66e, 32'hbd505e94} /* (0, 7, 18) {real, imag} */,
  {32'hbe2ec7b8, 32'h3db4d5c0} /* (0, 7, 17) {real, imag} */,
  {32'hbdc39498, 32'hbe8d5fe4} /* (0, 7, 16) {real, imag} */,
  {32'hbb753800, 32'h3df80a80} /* (0, 7, 15) {real, imag} */,
  {32'h3e53a96e, 32'hbe01df98} /* (0, 7, 14) {real, imag} */,
  {32'hbb095340, 32'h3e961296} /* (0, 7, 13) {real, imag} */,
  {32'hbe32a501, 32'h3e92f19e} /* (0, 7, 12) {real, imag} */,
  {32'h3e5143f1, 32'h3db41e54} /* (0, 7, 11) {real, imag} */,
  {32'hbe3b40a9, 32'hbe54bbe8} /* (0, 7, 10) {real, imag} */,
  {32'h3e518d0e, 32'h3e354ca8} /* (0, 7, 9) {real, imag} */,
  {32'hbd9e525e, 32'hbe560bf1} /* (0, 7, 8) {real, imag} */,
  {32'hbe9da280, 32'hbd84d830} /* (0, 7, 7) {real, imag} */,
  {32'hbee17a78, 32'h3e90177a} /* (0, 7, 6) {real, imag} */,
  {32'h3e92a3c2, 32'h3ea9f5e2} /* (0, 7, 5) {real, imag} */,
  {32'h3e3bdf66, 32'h3cf69778} /* (0, 7, 4) {real, imag} */,
  {32'h3e45e34e, 32'hbe11ed56} /* (0, 7, 3) {real, imag} */,
  {32'hbef4a89c, 32'hbeae7ef2} /* (0, 7, 2) {real, imag} */,
  {32'h3f596da6, 32'hbf487663} /* (0, 7, 1) {real, imag} */,
  {32'hbdd7ffec, 32'hbea0a24c} /* (0, 7, 0) {real, imag} */,
  {32'hbd822fbc, 32'h3f019710} /* (0, 6, 31) {real, imag} */,
  {32'hbf4e89bd, 32'h3f1e2916} /* (0, 6, 30) {real, imag} */,
  {32'h3e8488b7, 32'hbf638a55} /* (0, 6, 29) {real, imag} */,
  {32'hbe296ee3, 32'h3edcf7c7} /* (0, 6, 28) {real, imag} */,
  {32'h3f038458, 32'hbe65e4a5} /* (0, 6, 27) {real, imag} */,
  {32'h3d795568, 32'h3e25c11a} /* (0, 6, 26) {real, imag} */,
  {32'h3eaa21b2, 32'h3dea7ee0} /* (0, 6, 25) {real, imag} */,
  {32'hbcfa254c, 32'hbe29e5ad} /* (0, 6, 24) {real, imag} */,
  {32'h3e7d5bbc, 32'hbda83170} /* (0, 6, 23) {real, imag} */,
  {32'hbdc18b20, 32'hbe119bd7} /* (0, 6, 22) {real, imag} */,
  {32'h3e827bd2, 32'hbc6a96f8} /* (0, 6, 21) {real, imag} */,
  {32'h3e3ae08d, 32'h3c632920} /* (0, 6, 20) {real, imag} */,
  {32'h3e42233c, 32'hbe037bce} /* (0, 6, 19) {real, imag} */,
  {32'h3d586e88, 32'h3cc56300} /* (0, 6, 18) {real, imag} */,
  {32'h3e417bbd, 32'h3b8a4338} /* (0, 6, 17) {real, imag} */,
  {32'h3d3f7191, 32'h3e3c1f6a} /* (0, 6, 16) {real, imag} */,
  {32'hbdcf2eee, 32'hbddbb8f9} /* (0, 6, 15) {real, imag} */,
  {32'hbeb99698, 32'h3ec5a30d} /* (0, 6, 14) {real, imag} */,
  {32'h3cdb65c0, 32'hbe4133c4} /* (0, 6, 13) {real, imag} */,
  {32'hbc47f460, 32'h3e8c3284} /* (0, 6, 12) {real, imag} */,
  {32'hbd8182cc, 32'h3e83ac96} /* (0, 6, 11) {real, imag} */,
  {32'hbe715624, 32'h3ee03869} /* (0, 6, 10) {real, imag} */,
  {32'h3e8145e6, 32'hbe0af1ed} /* (0, 6, 9) {real, imag} */,
  {32'h3d01fe79, 32'hbe8c96dc} /* (0, 6, 8) {real, imag} */,
  {32'h3dd53024, 32'h3e1c772a} /* (0, 6, 7) {real, imag} */,
  {32'hbec5b992, 32'h3e091e86} /* (0, 6, 6) {real, imag} */,
  {32'hbe4ce642, 32'hbda64dfd} /* (0, 6, 5) {real, imag} */,
  {32'h3f0716b4, 32'hbe8eb088} /* (0, 6, 4) {real, imag} */,
  {32'h3ed50ada, 32'h3db45c6d} /* (0, 6, 3) {real, imag} */,
  {32'hbddc1a98, 32'hbe6eb2bc} /* (0, 6, 2) {real, imag} */,
  {32'hbe6b36e7, 32'hbe30d796} /* (0, 6, 1) {real, imag} */,
  {32'hbda6a99e, 32'hbf7c7d9c} /* (0, 6, 0) {real, imag} */,
  {32'h3f8ebaf4, 32'hbebe497d} /* (0, 5, 31) {real, imag} */,
  {32'hbf2d3a30, 32'h3e617768} /* (0, 5, 30) {real, imag} */,
  {32'hbf0b99ef, 32'h3ecb6c8e} /* (0, 5, 29) {real, imag} */,
  {32'h3ec23f02, 32'h3d1bbcb8} /* (0, 5, 28) {real, imag} */,
  {32'h3e18191d, 32'h3e88a1b4} /* (0, 5, 27) {real, imag} */,
  {32'h3eabec51, 32'h3e0adcee} /* (0, 5, 26) {real, imag} */,
  {32'hbe36de07, 32'h3b8e9f00} /* (0, 5, 25) {real, imag} */,
  {32'hbdbe4454, 32'hbed63453} /* (0, 5, 24) {real, imag} */,
  {32'h3e0373c4, 32'h3d682520} /* (0, 5, 23) {real, imag} */,
  {32'hbeca591c, 32'h3e884caf} /* (0, 5, 22) {real, imag} */,
  {32'hbef21631, 32'hbe1a8403} /* (0, 5, 21) {real, imag} */,
  {32'hbe593810, 32'hbe384952} /* (0, 5, 20) {real, imag} */,
  {32'h3e29dc56, 32'h3d1396f8} /* (0, 5, 19) {real, imag} */,
  {32'hbe673106, 32'h3e9b38c9} /* (0, 5, 18) {real, imag} */,
  {32'hbd32b73a, 32'hbe060916} /* (0, 5, 17) {real, imag} */,
  {32'hbd572b74, 32'h3e3f6484} /* (0, 5, 16) {real, imag} */,
  {32'h3e3b2a26, 32'hbe215a44} /* (0, 5, 15) {real, imag} */,
  {32'h3e5c2cb4, 32'hbded3b7d} /* (0, 5, 14) {real, imag} */,
  {32'h3e1ef95f, 32'h3e5f9f68} /* (0, 5, 13) {real, imag} */,
  {32'hbe487ffa, 32'h3d4c1718} /* (0, 5, 12) {real, imag} */,
  {32'hbb9c2280, 32'hbeae8819} /* (0, 5, 11) {real, imag} */,
  {32'hbe4517f8, 32'h3e2691d6} /* (0, 5, 10) {real, imag} */,
  {32'h3e1e367b, 32'hbdb7d278} /* (0, 5, 9) {real, imag} */,
  {32'h3c1bd958, 32'h3b4c4700} /* (0, 5, 8) {real, imag} */,
  {32'h3eb99b89, 32'h3daf1e4e} /* (0, 5, 7) {real, imag} */,
  {32'hbed97cb2, 32'h3e382e02} /* (0, 5, 6) {real, imag} */,
  {32'h3e33d0be, 32'h3e3f2f64} /* (0, 5, 5) {real, imag} */,
  {32'hbe3ca84a, 32'h3eedb3a4} /* (0, 5, 4) {real, imag} */,
  {32'hbeaff2a9, 32'hbe9e4730} /* (0, 5, 3) {real, imag} */,
  {32'h3ebddea6, 32'hbedcdc75} /* (0, 5, 2) {real, imag} */,
  {32'hbe998fdb, 32'h3f57dc4d} /* (0, 5, 1) {real, imag} */,
  {32'h3f6f0010, 32'hbdbbaf20} /* (0, 5, 0) {real, imag} */,
  {32'hbf5afaea, 32'hbf081c40} /* (0, 4, 31) {real, imag} */,
  {32'hbe0e65d8, 32'h3fa8d210} /* (0, 4, 30) {real, imag} */,
  {32'hbeb63d48, 32'hbe83d145} /* (0, 4, 29) {real, imag} */,
  {32'hbe249ea4, 32'h3e84c117} /* (0, 4, 28) {real, imag} */,
  {32'hbd481890, 32'hbe61c18b} /* (0, 4, 27) {real, imag} */,
  {32'h3d566aa0, 32'hbe9ad78c} /* (0, 4, 26) {real, imag} */,
  {32'h3f4cb336, 32'h3f0bce38} /* (0, 4, 25) {real, imag} */,
  {32'hbdaf0890, 32'hbf0a6271} /* (0, 4, 24) {real, imag} */,
  {32'hbf11d060, 32'hbeef9dcf} /* (0, 4, 23) {real, imag} */,
  {32'hbe050e62, 32'h3d0eb1b6} /* (0, 4, 22) {real, imag} */,
  {32'h3dc64a1a, 32'hbd87eb44} /* (0, 4, 21) {real, imag} */,
  {32'hbe6c5250, 32'h3e66bfde} /* (0, 4, 20) {real, imag} */,
  {32'hbeaa9756, 32'h3e4a0ea1} /* (0, 4, 19) {real, imag} */,
  {32'h3d651bad, 32'h3eb03466} /* (0, 4, 18) {real, imag} */,
  {32'hbdaba366, 32'hbdc064af} /* (0, 4, 17) {real, imag} */,
  {32'h3e27c95a, 32'hbe1e68fa} /* (0, 4, 16) {real, imag} */,
  {32'hbcef2788, 32'hbd08e8af} /* (0, 4, 15) {real, imag} */,
  {32'hbdda7a3a, 32'h3e6efe3a} /* (0, 4, 14) {real, imag} */,
  {32'h3d6cef18, 32'h3ca8af5c} /* (0, 4, 13) {real, imag} */,
  {32'h3dc4ab8b, 32'hbd963b42} /* (0, 4, 12) {real, imag} */,
  {32'hbe0d3248, 32'h3eb7699d} /* (0, 4, 11) {real, imag} */,
  {32'h3ee62196, 32'h3e3933a0} /* (0, 4, 10) {real, imag} */,
  {32'h3e3a30ce, 32'h3e64d338} /* (0, 4, 9) {real, imag} */,
  {32'h3ea8080e, 32'h3c8e2758} /* (0, 4, 8) {real, imag} */,
  {32'hbea48d1c, 32'hbf074adc} /* (0, 4, 7) {real, imag} */,
  {32'hbde01044, 32'h3dc2bed8} /* (0, 4, 6) {real, imag} */,
  {32'h3e9ecd13, 32'hbc908ab8} /* (0, 4, 5) {real, imag} */,
  {32'h3bef90c0, 32'h3cee57e0} /* (0, 4, 4) {real, imag} */,
  {32'h3e7011c4, 32'h3f805571} /* (0, 4, 3) {real, imag} */,
  {32'h3f28f9f0, 32'h3f79347e} /* (0, 4, 2) {real, imag} */,
  {32'hbfb201f0, 32'h3ec2a4a8} /* (0, 4, 1) {real, imag} */,
  {32'h3f344f1b, 32'hbebf2c90} /* (0, 4, 0) {real, imag} */,
  {32'h3fb3a764, 32'hbe63c504} /* (0, 3, 31) {real, imag} */,
  {32'hbf1e0af6, 32'h3f06614a} /* (0, 3, 30) {real, imag} */,
  {32'h3f233db4, 32'h3ecf82f2} /* (0, 3, 29) {real, imag} */,
  {32'hbec4cc1f, 32'hbe108fb3} /* (0, 3, 28) {real, imag} */,
  {32'h3ef66c44, 32'hbf00d3a8} /* (0, 3, 27) {real, imag} */,
  {32'h3ce8ed32, 32'h3e0d7896} /* (0, 3, 26) {real, imag} */,
  {32'hbd3e1d08, 32'hbeb338ee} /* (0, 3, 25) {real, imag} */,
  {32'h3e6592e6, 32'h3ec32a4e} /* (0, 3, 24) {real, imag} */,
  {32'hbe274892, 32'h3a7d0b40} /* (0, 3, 23) {real, imag} */,
  {32'hbe65b4d7, 32'hbe0f8d13} /* (0, 3, 22) {real, imag} */,
  {32'hbe30606e, 32'h3e074786} /* (0, 3, 21) {real, imag} */,
  {32'hbe88847e, 32'h3e0f7f18} /* (0, 3, 20) {real, imag} */,
  {32'h3ba7c4c0, 32'h3e746267} /* (0, 3, 19) {real, imag} */,
  {32'hbea9fc0a, 32'h3dcf693f} /* (0, 3, 18) {real, imag} */,
  {32'h3df7e26c, 32'hbdc6c0ce} /* (0, 3, 17) {real, imag} */,
  {32'h3b585e60, 32'h3e764c0b} /* (0, 3, 16) {real, imag} */,
  {32'h3dda3198, 32'hbcd62a30} /* (0, 3, 15) {real, imag} */,
  {32'hbea03e7d, 32'hbbd1d0b0} /* (0, 3, 14) {real, imag} */,
  {32'hbddd2074, 32'hbe456582} /* (0, 3, 13) {real, imag} */,
  {32'h3ec52218, 32'h3d5b2794} /* (0, 3, 12) {real, imag} */,
  {32'h3e486d54, 32'h3e1ab7b3} /* (0, 3, 11) {real, imag} */,
  {32'h3dffded0, 32'h3d0f6e84} /* (0, 3, 10) {real, imag} */,
  {32'h3d17a1b0, 32'hbe9885db} /* (0, 3, 9) {real, imag} */,
  {32'h3e8c4836, 32'h3cc3eca8} /* (0, 3, 8) {real, imag} */,
  {32'hbf457eec, 32'hbda5fdee} /* (0, 3, 7) {real, imag} */,
  {32'hbeb37fe9, 32'hbef4799d} /* (0, 3, 6) {real, imag} */,
  {32'hbe8dcb31, 32'h3eac67e3} /* (0, 3, 5) {real, imag} */,
  {32'h3f16c8c0, 32'h3f7f74dc} /* (0, 3, 4) {real, imag} */,
  {32'h3eaf456d, 32'hbf5b544e} /* (0, 3, 3) {real, imag} */,
  {32'hbf370cdb, 32'h3fdbd312} /* (0, 3, 2) {real, imag} */,
  {32'hbf02c6cb, 32'hbf9ab240} /* (0, 3, 1) {real, imag} */,
  {32'h3f5e95d2, 32'h3ed052ca} /* (0, 3, 0) {real, imag} */,
  {32'h40f44033, 32'h3e862dad} /* (0, 2, 31) {real, imag} */,
  {32'hc07bb0a2, 32'h3e0d3768} /* (0, 2, 30) {real, imag} */,
  {32'h3ee5c05c, 32'hbf5defee} /* (0, 2, 29) {real, imag} */,
  {32'h3ed61c24, 32'hbe4e82a8} /* (0, 2, 28) {real, imag} */,
  {32'hbf1ec512, 32'h3f8ea3fe} /* (0, 2, 27) {real, imag} */,
  {32'hbe2b37a6, 32'h3ec75e7f} /* (0, 2, 26) {real, imag} */,
  {32'hbd259288, 32'h3e8f07cc} /* (0, 2, 25) {real, imag} */,
  {32'hbeac923b, 32'h3ee8ff5c} /* (0, 2, 24) {real, imag} */,
  {32'h3c2a9ca0, 32'h3d7d2270} /* (0, 2, 23) {real, imag} */,
  {32'h3d7fac9e, 32'h3d518d80} /* (0, 2, 22) {real, imag} */,
  {32'hbe25812b, 32'hbe2b840c} /* (0, 2, 21) {real, imag} */,
  {32'hbe8dc2ff, 32'h3d95b914} /* (0, 2, 20) {real, imag} */,
  {32'hbd8fdfd8, 32'h3c2b661c} /* (0, 2, 19) {real, imag} */,
  {32'h3d18607a, 32'hbc150cc8} /* (0, 2, 18) {real, imag} */,
  {32'h3d2166da, 32'h3de5dc8d} /* (0, 2, 17) {real, imag} */,
  {32'h3d866a5d, 32'h3c42bb98} /* (0, 2, 16) {real, imag} */,
  {32'h3eb94f7b, 32'hbd88a388} /* (0, 2, 15) {real, imag} */,
  {32'hbd64927c, 32'hbe422bf2} /* (0, 2, 14) {real, imag} */,
  {32'hbeac2314, 32'hbb5147c0} /* (0, 2, 13) {real, imag} */,
  {32'h3e140a1a, 32'hbed4c76c} /* (0, 2, 12) {real, imag} */,
  {32'hbda9148e, 32'hbf1a7ce4} /* (0, 2, 11) {real, imag} */,
  {32'hbe1f318b, 32'hbe733898} /* (0, 2, 10) {real, imag} */,
  {32'hbe57c989, 32'hbe17beb0} /* (0, 2, 9) {real, imag} */,
  {32'hbf578e4e, 32'hbea76c4c} /* (0, 2, 8) {real, imag} */,
  {32'h3eb53c14, 32'h3d8fd624} /* (0, 2, 7) {real, imag} */,
  {32'h3f065b1a, 32'h3ebc831f} /* (0, 2, 6) {real, imag} */,
  {32'hbf414726, 32'hbf7d7cca} /* (0, 2, 5) {real, imag} */,
  {32'h3feb503f, 32'h3eab9a7c} /* (0, 2, 4) {real, imag} */,
  {32'hbe81ae78, 32'hbf32e1fd} /* (0, 2, 3) {real, imag} */,
  {32'hc03a574a, 32'h3fdc7406} /* (0, 2, 2) {real, imag} */,
  {32'h40205470, 32'h3f21e13a} /* (0, 2, 1) {real, imag} */,
  {32'h402d914c, 32'h3f3351a6} /* (0, 2, 0) {real, imag} */,
  {32'hc0c0868e, 32'hbe54e948} /* (0, 1, 31) {real, imag} */,
  {32'h3ffd3b82, 32'hbed2b7fe} /* (0, 1, 30) {real, imag} */,
  {32'h3f6e39b6, 32'h3c65b580} /* (0, 1, 29) {real, imag} */,
  {32'hbf8ab738, 32'hbd6f9e20} /* (0, 1, 28) {real, imag} */,
  {32'h3ffc6b5a, 32'h3ed2b368} /* (0, 1, 27) {real, imag} */,
  {32'hbc981580, 32'h3e2ac079} /* (0, 1, 26) {real, imag} */,
  {32'hbe134e91, 32'hbe6ace5c} /* (0, 1, 25) {real, imag} */,
  {32'h3e0c6d49, 32'hbec55d3b} /* (0, 1, 24) {real, imag} */,
  {32'h3ee52414, 32'hbf02562b} /* (0, 1, 23) {real, imag} */,
  {32'hbe826137, 32'h3eadc5ba} /* (0, 1, 22) {real, imag} */,
  {32'h3e9387d7, 32'hbf01534a} /* (0, 1, 21) {real, imag} */,
  {32'hbd31340a, 32'h3eda5d96} /* (0, 1, 20) {real, imag} */,
  {32'h3c8f7db8, 32'hbe145df1} /* (0, 1, 19) {real, imag} */,
  {32'h3e3ec258, 32'hbd584e8a} /* (0, 1, 18) {real, imag} */,
  {32'h3d53c3fc, 32'hbe656e7c} /* (0, 1, 17) {real, imag} */,
  {32'h3d964b88, 32'hbdc5bb2c} /* (0, 1, 16) {real, imag} */,
  {32'h3e51671a, 32'h3ce35cb4} /* (0, 1, 15) {real, imag} */,
  {32'hbe1b913e, 32'hbd810da8} /* (0, 1, 14) {real, imag} */,
  {32'h3e6b60be, 32'hbe565758} /* (0, 1, 13) {real, imag} */,
  {32'hbd91da41, 32'hbe0e09c6} /* (0, 1, 12) {real, imag} */,
  {32'h3efd81e2, 32'hbd4a66d0} /* (0, 1, 11) {real, imag} */,
  {32'hbe3aef38, 32'hbe68e6e2} /* (0, 1, 10) {real, imag} */,
  {32'hbdb5966f, 32'hbe1c186a} /* (0, 1, 9) {real, imag} */,
  {32'hbdc95710, 32'h3f0ae0d9} /* (0, 1, 8) {real, imag} */,
  {32'hbe492e41, 32'hbe613823} /* (0, 1, 7) {real, imag} */,
  {32'h3efe81df, 32'h3e68c852} /* (0, 1, 6) {real, imag} */,
  {32'h3f1b3910, 32'h3ed2d494} /* (0, 1, 5) {real, imag} */,
  {32'h3effe53b, 32'hbf02d502} /* (0, 1, 4) {real, imag} */,
  {32'h3fcebd20, 32'hbda9676e} /* (0, 1, 3) {real, imag} */,
  {32'h4032ad2b, 32'h3fd8411c} /* (0, 1, 2) {real, imag} */,
  {32'hc1210d46, 32'hc103b8de} /* (0, 1, 1) {real, imag} */,
  {32'hc0da7e04, 32'h4023a2bb} /* (0, 1, 0) {real, imag} */,
  {32'hc09d55bc, 32'h403b5f38} /* (0, 0, 31) {real, imag} */,
  {32'hbf320c7b, 32'h3f42d454} /* (0, 0, 30) {real, imag} */,
  {32'h3f01198f, 32'h3e3d7522} /* (0, 0, 29) {real, imag} */,
  {32'hbf162c74, 32'hbf64475a} /* (0, 0, 28) {real, imag} */,
  {32'h3fdde962, 32'h3e1430e4} /* (0, 0, 27) {real, imag} */,
  {32'hbe2c66be, 32'hbef7e7cb} /* (0, 0, 26) {real, imag} */,
  {32'hbf1c3a57, 32'h3ef7d1f7} /* (0, 0, 25) {real, imag} */,
  {32'hbb8e3780, 32'hbece46c3} /* (0, 0, 24) {real, imag} */,
  {32'h3ea1b702, 32'h3dc5463f} /* (0, 0, 23) {real, imag} */,
  {32'hbe1c0618, 32'h3ea24160} /* (0, 0, 22) {real, imag} */,
  {32'h3dd0d97c, 32'h3de48f5e} /* (0, 0, 21) {real, imag} */,
  {32'h3e74146c, 32'h3ec35b98} /* (0, 0, 20) {real, imag} */,
  {32'hbe7409a4, 32'hbd48477d} /* (0, 0, 19) {real, imag} */,
  {32'h3e829ec4, 32'hbea56217} /* (0, 0, 18) {real, imag} */,
  {32'hbe5f606a, 32'hbdcad3e3} /* (0, 0, 17) {real, imag} */,
  {32'hbd59867a, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'hbe5f606a, 32'h3dcad3e3} /* (0, 0, 15) {real, imag} */,
  {32'h3e829ec4, 32'h3ea56217} /* (0, 0, 14) {real, imag} */,
  {32'hbe7409a4, 32'h3d48477d} /* (0, 0, 13) {real, imag} */,
  {32'h3e74146c, 32'hbec35b98} /* (0, 0, 12) {real, imag} */,
  {32'h3dd0d97c, 32'hbde48f5e} /* (0, 0, 11) {real, imag} */,
  {32'hbe1c0618, 32'hbea24160} /* (0, 0, 10) {real, imag} */,
  {32'h3ea1b702, 32'hbdc5463f} /* (0, 0, 9) {real, imag} */,
  {32'hbb8e3780, 32'h3ece46c3} /* (0, 0, 8) {real, imag} */,
  {32'hbf1c3a57, 32'hbef7d1f7} /* (0, 0, 7) {real, imag} */,
  {32'hbe2c66be, 32'h3ef7e7cb} /* (0, 0, 6) {real, imag} */,
  {32'h3fdde962, 32'hbe1430e4} /* (0, 0, 5) {real, imag} */,
  {32'hbf162c74, 32'h3f64475a} /* (0, 0, 4) {real, imag} */,
  {32'h3f01198f, 32'hbe3d7522} /* (0, 0, 3) {real, imag} */,
  {32'hbf320c7b, 32'hbf42d454} /* (0, 0, 2) {real, imag} */,
  {32'hc09d55bc, 32'hc03b5f38} /* (0, 0, 1) {real, imag} */,
  {32'hc0885967, 32'h00000000} /* (0, 0, 0) {real, imag} */};
