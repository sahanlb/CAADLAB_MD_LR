-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
RgC9CO9Dwkz4EvAURdFi3LlD5FVBz/QbS3Skste+tKRVe+ikaKMUsP739GrAWwNw
gt0xBw7Q8tgDiyoliPF9sgwiIDpZaLakshiDu6FJtOvbYvVXk6iT+NOOCHgF+yU8
TE3iXuUKV7LW0pm6Ty4/gdJtXKEEDKWviOT1Tj0cj1s=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5683)

`protect DATA_BLOCK
+W5miNn07Q6PCgYG23iSHSulFer4qr1Ixy8lojoT+FgZS6W65YmF7bbelz/iTHjf
rprm6rTINOC3EhmrzMeG1l9iNbxEyQp9FUR+weeKgzsQEbqEl91/haT0OvT8Nd5K
kc548C3HlQ/Jjw4uyNoudBmrbRH1TE1iSTiMdrthhf75dZM8hemGuJB3l051LlMT
LhCNpdbD3M6MC/36Prcj4RksYunzNpKGNoQfk27S7kMcfen7wUicPs22/4+QQLtC
dIn0nXwNOAne0cHdmyeBIGdteQfoCo+YODNpnmTzXSfD3lNGLQYZy9vYBgswylmf
HWCalDQxUrjDgb8ZY35+KUPH5XFk8dbS2iuXAV6v5Kr590SAipweFN4ErVrboGWO
hRVb0IiDOLQA3tOTOa+ICRdZjgC5WHRCnqw+YVgEkd18t1keYap0b28peBuTHDD0
Wlg2CrjEMlDmpZ7IR8dJLQAxzo5EhZo551f4f+iN34SoyTf1yd5j5BQ/POOn8Eip
VR6nOcbA9Ct4wFAHpG8r/pwt2zO/yB+VuFuJWtJyVK9VA94IOVV3DEodYAiWA86v
svzhnNqs/jxXhG7op0QJmi2UiQedH8d3iuzuRJI3qiiUa61qjLID95waIBZn6KZr
72L4MtLoUx8WRVnqpSrQfDo8KK3env/Se2aQRC8cXNnR+/x72YnYO3HQ5J2uofDi
vUg9ZNrDqBD5hqsoBF7Q8sSjgQubCC+l+4mpq0TunMrxbz2OuzNTJlCYks/yv2eH
F/f1JCIHA1UuA9C9t0cE+y9AsmHIaC8eGikFibLbquLp5ncYkQ2wk0hWma1UKeAX
8RMKkhUBQEmw7/Pj6gzHiXx/bktVhLAOGS7kqvBfP2W0zYU1HEC+Nx+JLiXZSIsD
q2bUnKk8+FEBBD4YqBG6aRdC9Pu+tjD9WQ6WyUqUhQRQeWdXLwAV3ORDI90CwjeR
w0Ah1wi9wQrEVUyNXcLX+6scJkFOPQhdIlL5b8W+5tNR4uZfll8LAMGM6Q7b3qZ8
aJPeaqJZrMd/Zr599KhN7AzhTz9+wDsTyMx7PaAWAPgUYcmgrRpFtXLRR27eDxeM
WtmTaI2IZtHWO+F0KW8uU23Xdbs8xAE2qMoP7ryzs/gm+F9WIQj922XivNmC0Tge
fgNnutj7AIQWl2xdWUw6pB/BMOvju+QyIDDBLmH/KfZbHL3Jwj0tRyZ4HTzE10QV
uThmPTZp3dsA6T76tnN2hdS8EdQXzm3PRzFx8DERNKLKtCYRrCj2704MDS7xWgEj
eTwXG67bKLhThaUYLj/8ExEh5I/Vau1CeE/9PL0u6iloMpdLiNvAutYjg5DYAZCh
v6MUj+NObS0JDgwLxOoxh3Od6ziqaOLv/dciu/m/S+zIDIqsULByyN7l8UVzdl59
PwovGkmGz0Pk2wA7MJmfs3y1gDAZbc73mxmwjbH1EQLkOqdQzXGsi1NnrrZw4uNi
sXV9KJ4eeZjC3C1BKBQEqrcC32zBwDRhfFnlDeqNGST4VzNgVc1DVZGJvV80eFsB
ZcNDbB5jUXKmajNiL9+elow6GTNeYnKazPYKMy9GNJ3QPOqL550Isfv3ujtSY78P
IiR9Oi44HcAD3++0qlW9pgq7kbgsMB5r3lh6Avx5dYMNgrLUa/Abq8rtcXn4lkC9
A6MY09y9ADPz8EcvpNVMaUkQC3sarlXDmFnI7sRzd/qXFGfPRL5++NXXDvaRmWx7
SUARX7g7RJnaebpiA+rOAicENBdmROjIyNWHiQx8FX7Zz8doZSjLO3DnfhQn4ntO
mBPMmqn0i1E3zgKK0mPn5Wqu/iBhvk22+Kwhd67HiWTY1pfqiBnOhvloDoW2yfhs
R3Y97+qMiSw1LhkY30yaXkxk86+UEYxpPiTDLnjpBbqPYSwG1DAmxnSseT96JlzW
5nYewNI9hWh3W062/HgCwP3o/D0DYnLejIivEstWe2kTK6xMfHlJB6XMtsJIfJr7
obFTCznTswvUWuU77a/x1DZWy6EnNN9iYEtNEn3Qw/zrUenfuBoX3iOtNjiBgWcO
omGvcQ7OM85ggKQU9tRwsz8eH0YIp+klMpjGn5KXLwN8ansINziUpCx4i7MqU/Po
y//TZGh+BAuZ/xvPzXxQurdMsbSMkpyx0L5AA55c6k8oYZvisGiUua78yFfzpeda
gvKVXYl1APbF0APPjlO/dGCmx07kCkXs/VjMAIQP+bpzzt5JH38VHTBDadh0UyON
zZIISMz9vOx3zmQElmFn9gibthXd90aYWY/E12Wxt1mOa94FEYfGq+3Iws9c63YU
/3MQTZir2gfK9srz5X2cTlalMPaaAM0MORhbqZCXgQM83QeW1vvbPrtBw59/iz7e
qJPFYnC5ypZ30QataExWYc+/9GaiCXf7HFKPYop81wygX2+TyaPlAcQAJ0uPIGSy
yAstL+d2dBQbHBfhW0gWUxDETpVipsJa68Eatu0XB26r6iVPb+59OVu6rCLycHR2
RWUlGAVFXtyf0SjPPTcyMezSxxeOp+9lXwaDWr3noR/Re3JVKsPguanIVqkENtHY
LXiwGq4RCgeQ+rt7kDNYNiFTAId5DueU4OAMZ8SU73Ix7C00Y1ZKa/eWQ47r6k4X
U7G/cC+MuXA96Eqmo/CywUhAQCWb0I73GdPlULdlGakPLSnFJ//7CN1L/Rsza30u
4pi6Vki+Wuc5G44CZ70HUrwSUoN2a9C3vjVZPcKCD5+MNucedfwwu3X/tjB4adpd
B1O7t2s7SsChosuaWDs1cFoNP2tC8YZ/bj/tSFa7bTnCN0BD4rx/ubVuZouxsPfL
u5fe8Tn9m9tEKNYW2CWFvHwu9RyJNi4vhFm29UJQAOYLDEhRmgoLAR2c1ZEnkEHY
B5SYyVuV10URsNYn+O74xUwfSKfRp6UuwurNTX2Qc8rmBLDkWnZZqG5qKyyLaWTO
HEYjwd3OwblKBqvIYTcXqy6lqmau1n+iCbMg91h+GXw88u0ZXiefellv7qPbJZZV
ryu7vAvE6ua5owlSN9wuZa/gOkyzh3XhGjCuasJOt3sXBZQNcF/JkXLGffO0Ml4M
Y1XZtI7yLy9PphULnUbWe8DIUxrII75dTFNVNaO0mHsjgn6qLp9qpvRxpeNc06n5
woB6u10ov8uB2tWTbWfcR9xdgBOA2mcZvP++n2l7RO4k8pFmVJQ534/3fSd/D8Re
8Loc4514M520X0waNgk2jKxqXfALcICxzN1CWJV8y0rbR+QjBu5wIOKWEERlHnGr
H6PL4luQR3WBxyuwIaAU+9VELi5zo8pxJ8ygmonB/RhgXBrv/pBAIgBJ5wIBk84i
Nq9LL9VO2dUS8OI02wF33rVqvI/vL7UpwJSmxqwmE3GZDqgGbATAvb4vnk3wzO9n
nmtqE1PPqZGVm3iJYS6SWp1x3sLBecsSgN304m46jYd1sKOnEL/pQmAZx/ZgOJcL
dDe6ERtt0H9CJXa67fcJhhujQpMqANpDjSyzJaL6sX8VjRWuhfP7LjVA4yLPu9KU
3/5piSpAPx+/6aCBDXeEc2z9U34nPNBAGT/LQXWwPTgLyqwrHIPCJ/TcFBdydmeq
UFAKXHoVR004TnpXCkyPQIjnEftXXxQpMpY9lYOIL06Q+ssf/gCxRJsYZHaQICmT
xDKA4u4BYi4Sng0f5bbaTuID+RfMACpOl2E2DYlxdHCPiTqi9TaN5F2hAXh6BlZJ
KQUPSUzit6q3nNl330ffRVuoR7YCyqpATMjVmYfn3LaomjoUTOadV8dn/voH5S+0
Vf7Y8fqdz5CThXsCEwTCezJvNH8Hgq0O7P4gNm7Hf2j7jkam2RU43QYhF7ZgIKjQ
sE84fyojeQiPlB0a3ych1P6x3KAEduktmj89V+dkvlQGq1dZOpybQLz8ecmpp40h
FCPh6WBcmP4cS4wUAPVqAYgCn16jq7P5x7GOGpwvRhQi3RbK4ugpiCGAXzrL2Jgn
QiReM6/F8kuYmqqPTmSQ20nCLfCzb0x5bTblm3wtj2E/YKGVCApCAlMiUx08k6DH
Oq3TiZH3FAkbHIo4d93sfhQki62Ru60niQ3CTB0VGAsldxwRGpu8hWxAm+5X+juJ
sK/7Wcg67FGRZR0v0WACGBTskZ5vzsM0oTjVYJLB1ENIq3FB9YWVQDkl9iGaC+kJ
1sVk1alZtuZ04q/+A3XzkB7lo+4XDG8R1x4egDZ1wy8GCt73udd6wlT1jr84u/tk
b2PL89eN/Oc4FKYauR3Qm24m1rAHZ1UqdpZ/DOfrhu88ALsAQ5waOQyIS/7MgS3B
MpXI6mytRq0xhPjZlUKBEl9poDB4uxaECrojipItdtRH/xT3dcSZEKydCKTAzWXL
JfALkdTE4VV5pb/lh5Oa1cgGBBcfV10Zuemhp3eX6Y0tFHvM0QyYXda7zIHfTBBa
DMf0OUvBsEmu5TR+rbaYlGrVVAfXWduLff3l2otVDJfZbeC3ryVaN3i+m8jV20G8
DnTRmJFhiqfi25gMKo7cAbiJAcS26VtEWq9Fg6eoEYWw01c1zIjes+kOMxWTwfw3
DQthjWLao1bFMaYqbf/Ze63XYLfuyKsB0TZhjkzuMaFdoDUicH7dcX8TGGYnoTEQ
XEWM7Q07pKUVBAH6pBBqnnhFJo05SKiQMPRWjC2v6xGL+ALnP4svEJ/cn1RpSEBl
xhGgTuwD8FyKqJ9f9ME99JvEobv886V8yo9s7sE4H4QQ2HeIawPe00jmeHnpEtMn
9M0PKM0Id01/q2ASXplNBfwYg1vVPf3bGO1s0JE+BtrtZjrT6WfR8Bp8wE+wkuXn
uZVXQPOkhIuI5qthP+ESQ/ROAKKnsln/lsx3rJc8uAAh9Db4qaZC+RaIDUHQ+FvR
kv0M5S9glIctI0RUFoYhR9CyKTdqRrarRDVP7ZsxGtnIw/QmomWMveF2FRH/DlOT
ySQpeD7uOE1HBbJIybXgY2O4F6P5gntaxFIMUmu/pnEh2wQkc9gJxjj3CVWGbpzJ
TlKqoKoiTSKJ8SqCwCNp5qoqwLUQjI1DOIO1oYH7a5lVVFi96wYVbYtr4Yq9sRnk
f/hbw8iSxDnLm/2gBsxH4ifAdBl96MktTIdwJII1faoeaImpKO40GTC8Uty0U4YW
/6+nFAWoZCP6zhd43EtNP0SGmG0H87okTzFScfOKPsVgILK5sEoU9Wk3qKSqB2de
QfRzhdZewM9uGGraOdQbDqnoRne5G4XhdJ3tq0ocn8igVmkhN6bS0LAfzVQwIoxd
aaz981u8Afpzvu8jqgzhhfvz8HtMsb9lG2UTEZ0qAEoxGY1mWC7G0nKdayts6ZAO
NqxFUtWWf/h0FMtGmXMyKzaotfpFQzYQVInlyChzNIsjXFEnYQw6bpn5uF5UtWi8
NnMg4PZJjhS3aZ8aX/JmPYJLO+SBjJTAu7PkldtYDHwqyapjy1Crh/8ocvnoJCZL
Pg77F1mMiQ25Otd6JvPlTlLWl42Yo3B2WaUotzXot1J5JS30i3PyUHYm0jFTyl2K
9Qip8G1+CQMSjoveIcuyzmhGQCKFpgIeH9omkNykvti17JcYurm2E0oPcVBAZEzT
prY4tKH2/gWFgG9QmNeOpuebT0DLav0RfGvS3TUIPGGIZtZmyk1tS8LVNA3h5YVF
9OznTNawal2eKs+IbU6dI3Ppjc9MBeM6my+lRu1XY3HzvLKNzjML1QvXlKjxYbxk
yx8GdQf0MqeE5RG+h4gE7FIF4ce8N/BWQ/v7j3uqPoZZOpfwxN7zUpkJzNQzxE8Q
74a7LY13oCl/tev4rE1B/nMyOdqakxlZUcERjMm7s0vS7QXwL5B8GNAMG1/cf4jU
G20l4socfFerzlQplcWv2VTpifmO1m4ppJdVALv21K5HnWpF95MQ2l6y51LbzUWT
0cxGSe4at06XGZDdWfy4LOk4vD+jzmKcKtc0GfQTxDQX++q9e8sDNH0MIaMPtFfl
BVzy+QgMjuRcRWoDdizSDwev0wcZOQCG72FMkZOn8CuPeSxR1slFj7KUYHG52RXk
Owj3soZGrdmQA5IXVMz+rU5zgN+rMQbF1APrLKb5jD841KNnBXlSTYs1f7O92wW0
eTl2hNuR5SSq5QH25GYIedfThVtAT1rj4RAfd1oudg4p7J26SHHn56w7KiogGngv
cyHJa8PXgRlMVvEuFulGEjfNLe+E01pvNa/qL87fVU13L0VdIq3jtm1IKknuTZxh
S7kfp8CBbjIlMHddUYPtXACeiqF4jLCrUZtLg05U+aDDcyJfZRDPT4Y01nN1HIXB
Q0CK8KvFQWMPVW5/E8CI/S18GIHl1dxIPNNn1ftnJKBVvym7JqLY0Ovzqyze52Fu
5klQMkDG6aMeEV86V7sr3obnpUlFPcMO9Eyiwf3LYFyU1uUvoEVBJIdIGLIOqr8i
4zL0nU83wuUPAYlu7uGds3YO/T39W9BXIaIEN30qYqZbTAaQEWU/pFv5Lto0BqJc
RKh2qwtTLOKJdnAb2zN4g2i7NyNdaOkDpgSmhAmXr2royBSGy89kaDpEzMhOzjjR
acfrIeMWcdjDNq2JjYRNjN4S1axshvnPuOS6Q+3QCqHdHEwuW/fE69whf646ZmNs
JKlEmTW0xxJLxhy5Q34v/70COd4nyIfMTcUiu3mdk9ssT5j/TR2zA+Z3YEr05PYh
DX8GAR71zI9/ut7monszhHfsnYfuG9uLG18KqAPiboysbFWusjUo0JGzSR4cl4Vz
IjVUhGZmrNbdM9KeFC+aN/uPnGTcw0YpcZxlb8d6fbHWdfiY8pBIzx/6H7IEau3V
N6oPiPW0sAbX/DkCJCsOeBqfPTqhjsUm410aiKpchHvr6xiPfCc87Auz3vNQNiCi
SG6DbzW9xkmy0dZv6pMS6yHJCuwo6XXPNL30U2JIYU2zYk1aNlZYHLigqzHitoF8
s87N3y2p1yxuWQSpuPzA430a16fc1YWFdDqrdgPwPfBxfSIwCj36XwU9vgPOznSs
7GsA7q5JYLcRws7H0+14hP7vJXwnxFlTQENxq5GLFDi3IZzA/NJwS0wqcyNAkbSH
XbNq0yN22xZkdplqLR2lMrjctTwMR3QHKLZ4BqLy2JYvuz/rhqO8j7C82vsV6hJP
nuPy2Csp1G6t40l9VlSgw1KcJVy3PiBIhkyfmPUFNYEyuX5MaxeUHcGo6wVQ+q4y
JE5Q7Pn/ac0/nAQhL3EiyqwJdkwD7bPxHmzXUHXGA9mdnv7whdYkdooDxWNCshW1
KKsphVuCh4mXFOuglA4UxtPfIhIX1x8sbj0/X06Ywuq5ennj5lXx9DUYqw5dNcdw
6UUW/Gx3J4DvGGORdfhdpAJmK5bU7bKa+JMDvu+o6SPsMDOjkG2E0fI1rKEMvW7H
4Sz+jgAvQimeHpW1abW9QAkbBmVxZ8ckJOZM2O+j5AJ/HqBXePW9dysCBiU4Wyjn
bqtKBpoyzhpN7gPb8rN1V2uPk4uIBwVP7UtFWoCUdmvgPJHUbOt6IQfoQT/ur3IL
/9ujaRgGMpG6f2lZXBc8T1tmSbsjC7JYOUqku7D9L900aR5RObllpfYJAtMpuch4
1p8w90qy2NMRqMxw3GN//RGPhh9Da76OMxJfa1kLwYZM5xIRos93MviDbThf17aQ
`protect END_PROTECTED