-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Q44A81PR0gIQRJjsakQWpnUGtq9cJFXI9uOw1jf49hgQBitsUOyHi5ybhEsJPqH4
Kf67oJHCZUIRK5fKxVtYPYt+kBEW88j8tDbXSSP1hKoNASvxxiXfEGmN/CDnDTSM
8mK1Xsr/a9R8ZgMKM/+kxCCWk9J5M0DOYIwpaxCsXOq5wRaiiV1q5Q==
--pragma protect end_key_block
--pragma protect digest_block
OskUbLpDQ5ros+otF7/wRO6oViI=
--pragma protect end_digest_block
--pragma protect data_block
JlywjQmMvir6KxsVh2Zq6a8Jk1rEyTNOg1vH7tnPAYHFDk1vLYUeBqH+wgeZHPR3
V6EAiYZjTkkutygJqJTlDjXTKe5O4LyICLH74FEJ1dXo+unnO6pQ/rdpxM7KngE6
6WEuEJMa6dEBxTg4MZVliR0WROyBPWaRM5MGPzLHuiwg7f8ro81Joiz0CFRLY/XS
tORnWWSzuwYGQuw9vK57HbaPlmgLlHF1/uTVK/hGz63SJArem/v19iu2PD9iG5N5
bJs0UdqRT0zLAyt8qGc6ov1LZZDf9Hb/fVxMle2AGxvrzZ/Gj2MeM3qdjWlZgnxt
ZeXR571/6aRn1imjvSLtPtgxHHb055JlKiULnBIYpcTKermXjvD/U8A9C1st10PH
PCDOPV9NjvAczwbZphj9RVq5+QmBrU6O/wE8HGcAcFLPVbnn0enC8l1UFe5jhToF
Ir3zvY/YwKWXFLt4kVtHChb876279cdXALppO8dJhAn9DC9GKeocsR1PbH/4fysw
U2ZiQnchprT15Xk3UjHrd07ja12zy2lxMwPJyDleBfzQOzIi+nvViUeEKC7mnAn4
AuYItJ3asWDFIwYseVjTJ9OfHlldQvY7XM/YAU3ZdtruGdFvbdw/J2+hao1Omi5u
YOU15FJlmGn72tpFp/yTYRNm1ZYI5ksWvrrwsIvKx9FZ+a3VmNPTn1/V1EtxNkj0
xzRuHsV1C0kLpx176Lv85aik1qAOXAhdCLai7LIY293jwUT/dDp5UDm00vsH0o2I
UnMWIR8hREjlEH3yOm4j3EdshA6je1/mvH4XTRuJ0cUIezUW96QQnwvStpq+UszH
+0SoRXeI9Of3I/dDZqaozJoRI9Keowbk2MSj1zXj1wTF8TxQKmwiUaa9/dBHYG79
sz1JMElNjKDvS/fckEH1h4/YzqzUAbYSoIv+/3cRedG6+zoaGjZ5lFyumWFjAzAM
5G3jQdZwaqhWoSO4/UF6s0XUHszpHo75vFCxhSv3EzIqr8xUdGjo98A3fmFCy2J5
Sm0Y4uu6FA78blRtHW8sUtvn4RrLCUoSA6LvwG7yQ1npSRLLJC4farsXSsujR//V
G5R/FxUXOfa6qhryzd4vhQ7BwTExwfXvdxsrsXi2Hy+rdXORIHikHDX9q8IpE/lU
47TEScLyXw0XcyQdZEdfbIbf2bIDLSNXOfFtqQHkuJTsKtbs/uRfSETotSm3Lq/v
OHt3YDoEWpUvKH5IWQWR/BOdwq9fosy8lMQkbuWAo/NG0m5sK9EteTPsQjRuJEM0
10faBIDmI5GLQz95vvsWpIyF5vLmWUWYck58qka+V2nASL4yiSx8DjR8YJDr1o2d
VaIbL6og7O//NoevSukP6guZUA9p35nNYUtlypgE6WRPLzA/2TXQZVNMTYwYYCZy
BxNgPqeyiqyjyRxkY0xMeSeoMeqjkZ7Y6IVc2kB1YXQ4Fu9po64rjVX6oC/1eKml
OXyZLuZGfF7byNu63HJNe8s7bz1aj6IMP7xCRXpcuQXsy+yQIboNTaOCK6ssh5+B
q5AJAI51Y0KIiw3/4yrmXbnQSaoMvd9WFpNofQto0SgyTldZw25h5VcnXWBGs0ZL
HaD903cVcXXArmUtdSDGUnFqVEUWxyh4jttvzkcXQs1lNOIzdmNORvOKNBQcde8e
uHKLm06PNXNwu/vB7THl/4C+IPmfVVSCGWT6Su4HR2xwNLHtesFosD5a6L0aw3Ne
UdIKylZPUA0j9P1egV1IHuHQUw4WX5NphZKNiJIsZPfIg3Xl1CE+RPLs2YI1oxRy
OqrzcrZBZO2M3fEqnXaT+5CxrH5nYEM9c3VNaG9so82kxwjiBVKXI+9Dd9jWJqkq
A/3S6kIcICKva437AiH4YRBfhj3hRzoeLZPsmMcPglI0TCj3MMSgbI0kupolfS8H
02icG6HLWsEAbHvha+wUhJDSZrtzQsJ3l4tSLuYxzlqHV/3pyJNEtX/jlqO2KJl8
ZWhvirzj2VkSybDoQoTb1tANf02NwkgJBZ82wYUTPd1wlAacfr8jVwG9iQidu10n
W1xzI3F5m8kcOhIOKXrjSmVN14Ck35ZZGyB81AVn7aR6CH1EDFvH5qR4G6J87rml
rs4B+wx6f9d7FWIxRop4Ta3PCiPZvhb0TaoZ+rDcoqxOJLKdSwgTTQMToawre14T
mJaO0YnzwgYEeC2m1TVdGawAJj+xIPreWGvMhMEirWx5FFtxphaDJBgJwDg52C6W
d+4YfEIfWt/hMs6/5EItM9dgFbnTqZ+U2iEVZFzF64/SHD9ERCHs+ZG4Iy7+3ooY
b9RoZgk2TczYuywQ94EsUvclNHi2/YwD8r1RP2XDCIKGPdd3B3F0AN51CIJ90Lbc
hSnaT/otj27GBtz3EaBHMPA1wbpGcsiDEmmRZiYk7gErNvLgp+zSVzgMYghKCLTX
IsPkQcFlus8vMFIR2/VpeCD33tOEpldK5WHPwPKXlH+7U3HODb6jG5mqS3TUP9Zi
GbLXHseIDtG8qmSYePLKjLU3XYz37E7glB4kXzqqb3+MDCLJTrLyrlNs9k6EdyYZ
YQD1kfS/7x0gBsFyZdVmzHT5rvE6CrYYMLutlozo+3sAJP5T36tgZHD6XfIPWG/J
bJE495OzajCoD/X8GJxF3syOtTu8rtTP4ZVeGrziL0H2jZ4l3GUwKtdu4rhC2ty7
LwtbA01HRhyqVk+mPKvtzuFAnPch/qDz4u67wNlV28dkM9d0oLoPIrB+0ZnLO9/l
YYNJ93cYU9FNWfqx+WWSXvcazn4C+T9Gz+4zpk/hX4XopZVXmnyqR846LYJF+S3A
eB2qMxDUm8WAf1tsnr/AOpbIdf2x/ylsk5aZQLfpjXESkGTVPMI3sDfghg/9WwL6
LsJTYz8orW96H2k2FvHdV64+xxaU4UneA/hDuTN8hwMBgbhgaW8HCMkYC8UMwMt0
KRNh6/QIu/k2SQ0hoMGOUeXA4FFv2brNXtlj4JUOVE8dyfp0MCwr1/M9iT1tjyKk
15u2dBCI1G5nd0Zy2JOqfIWrGrM0P9MP4ppHgZd6DQd20aaHCcM/9GeUodFhq9zz
rsYNTYVheXxvG1ZUG8rYzVOqD5F5Jgruzcy6NFYLzWd3MbTaZy1p7GtHgH/JblD1
gO0zXfUapYgfB7A0HQsai1ud5HLUU6mDC32ICjEGYowxQp1xJb6b2KdqNmAxV/W5
f78bN6rG0X6+WuYd7V+LZ0hGsMXMjqrhdiZN7+RgYU/NJEl1qQEU38DZwpgO42sW
dTRiF3bZ/1uO2nA9fvsUR6m9i0Dp4QsWPLHEdfy2QzPGP8cxw2dIS/18mY/PRd7a
6dCnPqNSnrX0WkrIdfTH4vMSaYiqOeGI+wA6VoVsEMnv/IxsVGeEDdPY/g9OkHmL
uf9jBNmYlKhnCXwJtdOYs7O1B4GzgB/T9xj0MgT9eNcN3GM5JHfL5iXlGQrZ4EVU
Smpz6zwG4NX/sbxrG6WB12Vpn5ykBgd4IjZrcPU+nNcgwXaLESi6lbyA0u1uZfTN
INa/gwngU70Ix9QGhzn0BWSCCRG5fHwOZSZVkonclhuORaf3wCG0GCh2ZOsxe0GB
Vk3+J4spaaD9t7ItGedYitqCj7eIuJ1dbdvKvAr5lW/LMUsXwV8Gc1+p43VVlRlI
Dl4dnkD0Y3ilF+KvoQE/BsTEWyuGhiF/Ym+G+BAzhggrQ8dmtY5v9MFdXJxOJ/sI
Ca781ZZnEzSo1/kdl3YbcGa4KlxIV7DIgutpBsgv8f07ZRGV68TJ7y90Q5QSd6ky
VB+pymtQZZKtkQDIuQoIlenKU5YwcSun65RQ3ZEsXyGFh7RMa50QDPrskAwUPO4G
H07Qtls0WUe7UKnht3JnsSUgUPIs57BOwmIFEV8ZN5kgE10hc3P+OHYRSP5QjDf/
+aMUphtBFCFKAdQGW05k3tBEvijdgejrkVwLOeb1Fg3yF+BHOMwQaD8aT7I6HRyD
BrxoTqIaVD+DYTgOFN8QA4VcSZ1n0Hpb4gZwPoezxZGxOmAoZe4N2thTxTGXawfz
r01nQRp70V/mTfBvH+xn+JbKrgMqg7tmYqM3/TUWxiamESPOIIFPoxmcSUu/ZBU9
z2NejWuFkTqLM3VoEMl+C6hJbknjFskOtlUK+T+iHkuol7AQl2sQkeDHzWD0V1il
d2SPthxxCeSeEKAOF8QExqohT9Qmafj0ZtmQl3jy4xEpOc8GongfaNT69SLwGSU3
aHyCCv0vmqHkR/B4kc1sBUu9cHry9kgZNYr376zLPZ0tqcwseITyTMOHrxi9Ujz+
24d2vJj54/HvVB2W3aDqT7WDEKsskP3aBLh0rwB4NZ0zcESqaJAG+m4K+3MHS2wJ
mY8mSxe4Fimc3Fl92QQkYP1umPvtfTcADjbANPs1eq38K9t/DHI8A67cQXjrE8s4
KoNblcVMYI1A+nXXPOJbzm480YGsXYOLnsw7xv37yBJSR7kxl1r1/+tsXqWUjLkA
S8W1xL42Sh3Us0Zxc7unCzu5w0lPqoV3SCM2/C8pLmzC9TzVeduT/KJb2Ngmt4tS
fiqfLkMhpZFsklxWj2V8vlfeYX4nctnUxLHcYTbSWpzsfWH2doX8plJ71xDXSZsz
5JgG9rF3lGZAxDuT6tiGt9Ku3e4jdhNdh64FwVLy31+KTz4R3sS2eLZF2b59nMAo
NZ0OVv/6LDFSiFVJgC8mP+YbG1XIX93+iqH26cbkbDnEbBpUPd/KkBsdMRl9iLyH
LKYpUEVUBeaXlfErgqlxxT/gBYNplsC6lh+4Ga3nlRAZMp5BlGNzXgg1kkZIV0q6
OhzG2mJKE4aTk1laNHsjThuxtBS41+s7mFYquAO28ENeXTYP9E/x+bt0GdFOC7Mi
dKjniUQFq77RAuacnOkQMXe/KJKiFxWz9b2wmpZZL1DIHa2FVmDVEfxjS9V+7lF3
dvzy94Y0a67SnPEb5VK/SVQo7IgfkWj2f0NSmFzubymOfCaI1uPMZ70bMJPFSrBI
KI3lxdaNXQ+ud6KseE5INRiXwmlFMDikbbAAk6orWJEnnGVUpCSieT7zz3vLyyXI
qEY6fMQnIqzz04LHCcnpAaMX4thLIgG772Nt4vuKyGJfwNtio22Mbe+91jhYh1qJ
zs2GkBYwcskUc+EY1kn5JmhNxtsNEfYSJiq6bCEFRUep0rO2bt44XP1dLaC2uJXc
SZ9x96PUYnKzu2H3LpF2zuMuyJjxonHrCsSZVF86+EVucJWtC0Vg97pCPx2U6tki
xw80Yo3zt7Gh/nDrypkuFrxCUitc1YPxon/o7lZjeE2i6bvDw35H5sFAIsDP0iso
8yXdeQBoi/JJFis1gxo+B9Nz92crWwTK5jhFR91JsEMUydInUwqUmb+r6hDxi+C5
WeeqdJO1cVEb5YEeCxF+eOhWlVmKl342a4R8A2mPEUFzHg+QCko4F9VnAfLux/eF
1+aWswuOa6/3ByGncr5uYIfEOSs7LnlZ6Trk4KNkrTkIXmg0KBMXAdVTQtLQuaMk
aNvSxXsv3I+zrFf4sQbOuzlZ+0cSGTk0qc96f3g0Mm1DJVTiiSOwN1fkNXf16lMg
zcIgos2mh7Wk5+bmrpIPYZZIbzN7Wq4EfkysWxZEAQCWmUZ/2pbofoudQikmOnn4
qVg7bryzbvgBqE1/ygxsUsmqgbafngilsrqptS9MTIbB97yMp49PPLf0/Z+UUEix
/jCfCkUxkr/VgLhhZWRMSpa4ix8PYGoowI4XF6FoYPiDa2iCFetIyqemfXhta9t6
hmcTYOWcTS1MiCgZ0JO/SSwcEo90iyJaB3tIA7mk6FiDgNcgrjQEFe9lsO/Xq/8E
S9mzxd+coVudG9vGHgTJ/Yu+UBemSSyH6HHTzKibDAbWPTv+NJnoyONwikVSuAb6
8I9MKDjL8ryzhsxl7esTl5Jdky8S2GhFE44IvofLjV1nZQzASt/lrCDMb64Dtjnw
rlsCXRfQ9OhVDiaBngxdrFahSvwpenbWnvQMwWNK+XDMR/HM7r9dPBDUecvgr7xg
Ril9gh88NhXCa5rIgX6/T0MfUF+ihtPkgGTxqBnFY7hr3vdcrtrdudmfD7iEzDGi
mgpwkGUXFkxPe3i2cR8ft+kGM9gnRS7dwdW0kqvkkpEeepUJT637GJOzbS6avi9Y
IwQ6dMhN//zGkfbLCEFTuKhn9iwTkR4aKH993h9lkteaChaJPF/EldUQTiuO44be
+8dZfSAUE+Jp313yW3rxlKACSYbYzTfWfbLxW+bvS8mAXlN+ALjnAo+l4wIR3Bm4
A4kp8aHLJhtFzhvnMHyHczj6yOXCkTePz0MLuldyZ40nQe1ogYtvQJbMl/mZNPI4
4xIbRPo5uk3/X6lW7JgjQdHO6SnMPc6EpVfazgXl94PVPAm6d9Boev4aEtCdX4FQ
oSWby2Z4VYRi+7dTSQmafQeitVO1ww+KyrW/dZOVW4+9qf7lxKAgjoNBn3NLbdY/
5OXlXZTl9RnAjGC/kyJwEDze4OiakcKCrZ0R6JH6+t4xhZDOuayKHxtuKYxTTtuB
lFeaMvCz027F0G+IVCb9pZFWNduWQeS8MtwdC3nCjTUue3pHLKlfyNeD4gGo4o9N
8rPVE+5jug8cWOCzsYwOA3OSkrOwL4dg7U9gjrwXHJ25yEk0RJiZuq3TKhydcQ3T
jEzj5IsPjFj7ePBe/dt/He9TO4dKlNGepOjvPuzJcXLmMXOBbZMqIuOdXdiGJfq5
krZyeyN8WRTMKwbA83cUOuN/hLpOXW3ax4RlQNasQOw=
--pragma protect end_data_block
--pragma protect digest_block
d4thxYif4pwdjQ4fQvUclazGPrM=
--pragma protect end_digest_block
--pragma protect end_protected
