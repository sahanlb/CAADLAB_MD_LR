localparam [0:4095][0:2][31:0] P_FORCE = {
  {32'hc41ca24e, 32'h435160db, 32'h42832ab9},
  {32'h44268986, 32'h42f65070, 32'h441cae5f},
  {32'hc31e4319, 32'h43e12906, 32'hc3f2b95f},
  {32'hc31fa70a, 32'h441e929a, 32'hc3b24c50},
  {32'hc2f3838e, 32'h4390b2b3, 32'h4386a8a8},
  {32'hc389368d, 32'h4393c268, 32'h43854b1b},
  {32'hc31a674f, 32'hc3171daf, 32'hc3180c3e},
  {32'h423548fb, 32'hc3d0ebd3, 32'h43de1d2e},
  {32'hc4113e72, 32'h4276e571, 32'h43e12c6c},
  {32'hc33d1421, 32'h437db54c, 32'h420a6d4d},
  {32'hc1666ba0, 32'h436e4ceb, 32'hc2ed99d7},
  {32'hc1c317f0, 32'h43ac294b, 32'h43a33cc3},
  {32'h438b6f44, 32'hc3211758, 32'h43b34ee5},
  {32'h42ce4787, 32'h4275cdb6, 32'hc3d2fc2e},
  {32'h4315792d, 32'hc3c386e5, 32'hc0586719},
  {32'h44039fdf, 32'h434780e8, 32'hc3d3400a},
  {32'h41f4b676, 32'hc32bea54, 32'hc327aeb3},
  {32'hc1a41c18, 32'hc2d0541b, 32'hc385314a},
  {32'h42930ecc, 32'h43c25b50, 32'hc302acc8},
  {32'hc3831d54, 32'h4300232d, 32'h43478830},
  {32'h43ab5744, 32'h43ace7de, 32'hc3841b18},
  {32'hc3fb0ebc, 32'hc36fe305, 32'h4396db16},
  {32'h42341c82, 32'h43100782, 32'h441d3c83},
  {32'hc35fe150, 32'hc3470b47, 32'hc26f47ed},
  {32'hc3e740e2, 32'h439b785d, 32'h4421888c},
  {32'h43d27c8a, 32'h430f5d9d, 32'hc262de92},
  {32'hc1b52c3c, 32'hc2a9dbc1, 32'h4225e64e},
  {32'h42d308f1, 32'h43413fc7, 32'hc35e5603},
  {32'h4385a1ef, 32'hc228107b, 32'h443442a5},
  {32'hc2ef3e4c, 32'hc387cef6, 32'h439ac31f},
  {32'hc315467d, 32'hc3fbbfce, 32'h42545ecd},
  {32'h4292fd8c, 32'hc2f71331, 32'h4412697a},
  {32'hc2a28a5b, 32'h4316df2f, 32'hc39e64e0},
  {32'hc29f615a, 32'hc2cfbd8e, 32'hc32c5007},
  {32'hc33c43b9, 32'hc3b677a6, 32'hc3949a68},
  {32'hc401eeba, 32'hc31fd0c8, 32'hc36c25b2},
  {32'h431f3ddb, 32'h43e46995, 32'hc39e1a05},
  {32'hc340c646, 32'h42c34957, 32'hc2bc11f2},
  {32'hc2f1a1aa, 32'hc2622041, 32'hc3060e47},
  {32'h4321daf7, 32'h43a6b770, 32'h43fac69f},
  {32'hc362c8fe, 32'h4392965c, 32'hc1818dae},
  {32'h42d0a190, 32'hc3b9a70f, 32'h42362897},
  {32'h435ff349, 32'hc30aae3c, 32'h42fc32b5},
  {32'h4354e9f5, 32'h4291d084, 32'h420fa857},
  {32'h43d1c08f, 32'h42c7c722, 32'h43467790},
  {32'hc31d0b8b, 32'hc3822528, 32'hc38c975c},
  {32'hc2df9276, 32'hc394b79a, 32'hc31d7b1d},
  {32'h43ceeba2, 32'hc2f1b64b, 32'hc3644a76},
  {32'h43a3a8e8, 32'h40afd8d4, 32'h429ab18f},
  {32'hc16836d4, 32'h43d96a21, 32'hc16390da},
  {32'h433317f9, 32'hc2178a7b, 32'h42b218a9},
  {32'hc34e0631, 32'h427d5983, 32'hc29eb618},
  {32'h436d9960, 32'h43167bbd, 32'hc239dc81},
  {32'hc2dfae0a, 32'h4386517f, 32'h430f49ee},
  {32'hc2f29bf8, 32'h43a011cb, 32'h435faa7a},
  {32'h4380c0cb, 32'hc3d4e760, 32'h4363aa67},
  {32'hc18aa6b0, 32'h43c6b8d2, 32'h41bf309d},
  {32'hc40dfff7, 32'hc3998033, 32'hc40f9d70},
  {32'hc332ab18, 32'h42b3a545, 32'hc1f266e4},
  {32'h4333f497, 32'hc2bf7c10, 32'h41e2f754},
  {32'h43c749b6, 32'h431438cf, 32'h43815c49},
  {32'h4188883f, 32'hc41e3e51, 32'h4272121d},
  {32'hc338beef, 32'hc3744043, 32'hc314e15e},
  {32'h43384a10, 32'h43b24462, 32'hc2b2a265},
  {32'h439b89ad, 32'hc3165370, 32'h43ab1e93},
  {32'h439e895f, 32'h413df954, 32'hc3de2a36},
  {32'h43aed9d4, 32'hc2a86065, 32'h4286df2e},
  {32'hc2b26624, 32'h4363989c, 32'hc2ec84c6},
  {32'h43310595, 32'hc3aac707, 32'h40b118b6},
  {32'hc31bc1b3, 32'hc2c392f5, 32'h436e2473},
  {32'h4387acc2, 32'h4306bf26, 32'hc36e229a},
  {32'hc213a2bc, 32'h43887415, 32'hc36df70b},
  {32'h42b6abca, 32'hc26c98c7, 32'hc342369d},
  {32'h436e1caf, 32'hc3fd6698, 32'h42592724},
  {32'h43040bab, 32'hc350d654, 32'hc3438fe3},
  {32'hc16b9fea, 32'h413ac65e, 32'h41d0ae7e},
  {32'h43abebe7, 32'hc3e779c7, 32'hc3f387bc},
  {32'h4255ee66, 32'h4234ea48, 32'hc382ec34},
  {32'hc391b550, 32'hc3c1d006, 32'h4404f08c},
  {32'hc20f7bf7, 32'h4367ae0f, 32'h43ab6407},
  {32'hc12c6d9e, 32'h43267185, 32'hc3051133},
  {32'h43cf85d9, 32'hc3d8091d, 32'h43e829fc},
  {32'h4350209b, 32'hc31727a3, 32'hc2be98da},
  {32'hc4430c6e, 32'h43cd3630, 32'hc221e8c9},
  {32'h431f8ecc, 32'hc40a9a29, 32'h413370dd},
  {32'h4305aef1, 32'h4360c28b, 32'hc27f9ec7},
  {32'h42834eda, 32'h4348cc01, 32'h42db3ae7},
  {32'hc37a9e29, 32'h43078520, 32'hc304320e},
  {32'h438c217b, 32'hc2a745d5, 32'h438c2e71},
  {32'hc241d2c0, 32'hc31b574d, 32'h43c87f24},
  {32'h421c1439, 32'h4246e4f2, 32'hc1413c09},
  {32'h43ee5874, 32'h42985f35, 32'hc3ca7d9f},
  {32'h428677c3, 32'h43562d97, 32'hc3ae05e4},
  {32'h43a46e19, 32'hc1221fb0, 32'h42de3b00},
  {32'h420d4a90, 32'h44175377, 32'h4370ec0e},
  {32'h42ce3646, 32'hc2fb11d2, 32'hc383638d},
  {32'h40ecf436, 32'h42ff201d, 32'hc3a3a4b8},
  {32'h4306c874, 32'h4101dd97, 32'h42abed22},
  {32'hc3987b57, 32'h42f063d0, 32'hc2f3116d},
  {32'hc2c791f7, 32'hc353aaa0, 32'hc36a9ead},
  {32'hc302396c, 32'h4380f856, 32'h42c5f59f},
  {32'hc2c52b21, 32'hc204569f, 32'hc2d0e563},
  {32'hc21943cd, 32'h443b751a, 32'h437afdf9},
  {32'h43aca284, 32'hc30ae4d3, 32'hc34260f8},
  {32'hc2360236, 32'hc1591be3, 32'h42e73af6},
  {32'h43274b90, 32'hc3813cb6, 32'hc3754a8a},
  {32'hc1faaa91, 32'h4388d87a, 32'hc13d1453},
  {32'hc2de3883, 32'hc343d12a, 32'hc36d8012},
  {32'h4371e611, 32'hc305d318, 32'hc2199180},
  {32'h42e668d6, 32'hc35b5db7, 32'h43995281},
  {32'hc36e8eaf, 32'h4387d6f9, 32'h4357b753},
  {32'hc402728e, 32'h438ac07b, 32'hc2bce23a},
  {32'h43921a3c, 32'h43086ed1, 32'h4398421a},
  {32'h43ad6295, 32'h4289c4d5, 32'hc388cf17},
  {32'hc3dad64d, 32'hc3b09d7f, 32'h4286fed4},
  {32'h43ab7870, 32'h43372385, 32'h440280ce},
  {32'hc359edc7, 32'h42e06190, 32'h41a1da1b},
  {32'hc201ea5f, 32'h4123a384, 32'h42af6c94},
  {32'h41b0996d, 32'h4312aca7, 32'h42f9710a},
  {32'hc4383d83, 32'h43eb35c3, 32'h43bb025c},
  {32'hc2f809ca, 32'h4387906b, 32'h431875c0},
  {32'hc320c1df, 32'h43436d46, 32'h43668f38},
  {32'h42698740, 32'hc3ca076f, 32'h4328411e},
  {32'hc10ef43a, 32'hc2c572dd, 32'hc223129c},
  {32'h43bd7c7c, 32'hc3bf8d92, 32'hc2407bb9},
  {32'hc3025bae, 32'h422759e4, 32'hc303353d},
  {32'h42a09250, 32'hc2d00eaa, 32'hc3ca3c2f},
  {32'hc0cdda9c, 32'hc35f2b68, 32'hc3ac3a49},
  {32'h42cb3414, 32'h43137deb, 32'hc2e7a519},
  {32'hc39a4066, 32'h43e5c98d, 32'h4413584d},
  {32'h43ceaeb7, 32'h43a41cfa, 32'hc2c6216a},
  {32'h433bca26, 32'hc2de03a7, 32'h42936200},
  {32'h430336f0, 32'hc3956be3, 32'h4380b83d},
  {32'h423c877a, 32'h42cc4f3f, 32'h43fedf21},
  {32'h42ae9cf6, 32'h43d6ee05, 32'h418b69ac},
  {32'h4382d25e, 32'hc39bd342, 32'hc2531655},
  {32'h43422ccc, 32'h41ce0d67, 32'h43bcc7b4},
  {32'h42da1ff3, 32'h40f308ff, 32'hc380faf8},
  {32'hc2ac5661, 32'hc263c11c, 32'h4294fa2d},
  {32'h42c25f95, 32'h43b5ba00, 32'h4386303c},
  {32'h42d4b8c3, 32'hc386760d, 32'h435c895f},
  {32'h42d30e1a, 32'hc39ac121, 32'hc35bfefe},
  {32'h41ccb20c, 32'h4323d558, 32'h43605d4f},
  {32'hc30c1060, 32'hc2c04faa, 32'h431be46c},
  {32'hc345a10e, 32'h421a24d5, 32'h43ed6b13},
  {32'hc3916f41, 32'hc3c5c809, 32'hc2e56f17},
  {32'hc35c8e8a, 32'h432c7662, 32'h43225ce4},
  {32'h438fa5ee, 32'hc31b038b, 32'h4303ef61},
  {32'hc2fa8538, 32'h433361a7, 32'h43304df1},
  {32'h403c29a0, 32'h4357209d, 32'hc28312c0},
  {32'hc3164a52, 32'hc313209b, 32'h42e2b462},
  {32'hc05275a0, 32'hc39bd96a, 32'hc1ed6995},
  {32'hc437893c, 32'hc382687a, 32'hc23bf330},
  {32'hc2fa2c83, 32'hc380d1aa, 32'hc3aea0cd},
  {32'hc2ede284, 32'hc3a801ff, 32'hc24f44fe},
  {32'h433ad501, 32'hc3c9cc62, 32'hc28b6263},
  {32'hc38bb613, 32'hc2e49459, 32'h43077ec6},
  {32'h4476c2c3, 32'h43cdb07e, 32'hc337c653},
  {32'hc38e1c50, 32'hc335eff3, 32'hc3839a90},
  {32'hc414cac4, 32'h42befda8, 32'hc19a42e8},
  {32'h4331fc47, 32'h4314b1ab, 32'hc39ebddb},
  {32'hc2be1ce7, 32'hc3e73dba, 32'h43149471},
  {32'hc31f685c, 32'hc2a1f0bc, 32'hc2a940a5},
  {32'h439839e6, 32'h4272e380, 32'h425dc102},
  {32'h42ba0cec, 32'h41e22c00, 32'hc30e178b},
  {32'hc44d6a36, 32'h4341f87d, 32'hc3d1606a},
  {32'h43a04fdb, 32'h4289d6c3, 32'hc2adb908},
  {32'h438001f8, 32'h43834b1e, 32'h439f65a1},
  {32'hc1f40b88, 32'hc37b01ed, 32'h42d2666c},
  {32'h43318393, 32'hc2c67ba6, 32'h43cd2cb4},
  {32'hc2f4da17, 32'hc32ae7d6, 32'h4385901b},
  {32'h434e9409, 32'h427fce45, 32'h4073ebb4},
  {32'hc28e5fc8, 32'h41d5bfff, 32'h4382e51e},
  {32'h4268d4ae, 32'h43186e54, 32'hc311df2c},
  {32'hc3014634, 32'h42cba548, 32'h431e14d1},
  {32'hc2b792a6, 32'h4376b4d9, 32'hc3c38cde},
  {32'h41a5e840, 32'hc3f5dfff, 32'hc1c3ebd7},
  {32'h43462a43, 32'hc1b194e2, 32'h43a36582},
  {32'h43c3a59a, 32'hc2bbf4d3, 32'hc3dd1535},
  {32'h40ae66d2, 32'hc2d17100, 32'h42b03c4f},
  {32'hc2d6a20f, 32'h429ee39d, 32'h4368eb05},
  {32'hc341fb64, 32'h4384d55b, 32'h437bf90a},
  {32'h43e6ffad, 32'h439d9fe1, 32'h4385fa9e},
  {32'hc3cc3550, 32'h42e0707d, 32'h4310b999},
  {32'h43c33198, 32'h422cf70a, 32'hc3a8fd8a},
  {32'hc38265b5, 32'h43dc610f, 32'hc4032943},
  {32'hc3602e84, 32'hc2c83638, 32'hc06f51db},
  {32'h43b9cf44, 32'hc27ba4cb, 32'h42c72550},
  {32'h42854f0e, 32'hc2edddfe, 32'h42ca8bd0},
  {32'hc30aafb9, 32'h3e8ad6e0, 32'hc3648105},
  {32'h44012ac4, 32'h3f81e0dc, 32'h4418be39},
  {32'h430df7b7, 32'h41c64a0c, 32'h4383ae42},
  {32'h43c01625, 32'hc281c7d8, 32'h430bac3e},
  {32'h43793b88, 32'h4383ee9e, 32'hc3786086},
  {32'hc3b92116, 32'hc3875a1f, 32'h429e0201},
  {32'hc31ad738, 32'hc36a4211, 32'hc3f7db68},
  {32'h431a12f3, 32'hc33d7783, 32'h43955e72},
  {32'h4376b5aa, 32'hc35210e9, 32'h4395ebb7},
  {32'hc2286d80, 32'h43959ca7, 32'hc310e82a},
  {32'h431b324b, 32'h4324e0ff, 32'h40bf1162},
  {32'hc3863fe1, 32'hc192c595, 32'hc400abc5},
  {32'h430e8f4c, 32'h4237ec36, 32'hc2d0ac7e},
  {32'h4384dcde, 32'h43b2d6b2, 32'hc397953f},
  {32'hc440a6f2, 32'h43eec89a, 32'hc3af6bcb},
  {32'h423fd1b6, 32'h426a53b5, 32'hc20cda1a},
  {32'h43f8efb9, 32'h425d170b, 32'hc3c63c25},
  {32'h42489db0, 32'hc2d728d0, 32'hc1913f6c},
  {32'hc213345b, 32'hc3959276, 32'hc1918596},
  {32'h431235eb, 32'hc2f188ed, 32'hc39b81e7},
  {32'h4422a05b, 32'h439b5f5d, 32'h430bc461},
  {32'h43975a61, 32'h43e480da, 32'h42e5f74a},
  {32'hc39d9e72, 32'h4326427b, 32'h436a7372},
  {32'h431096b6, 32'h4395396d, 32'h4282aabe},
  {32'h42bc08cb, 32'h426c31dd, 32'h44065db6},
  {32'h41be0f0a, 32'h41ac1d73, 32'h4348dda2},
  {32'hc37fe386, 32'h4216d557, 32'hc20e8566},
  {32'hc30ca624, 32'hc1fe4872, 32'hc39be034},
  {32'h42392fb6, 32'hc309044a, 32'h43c4d0a9},
  {32'hc3719261, 32'h439a95b6, 32'hc302cb9e},
  {32'h43e75048, 32'h4304fc19, 32'hc2866f52},
  {32'hc1eb60c0, 32'h43fa667f, 32'hc356577a},
  {32'hc380ced2, 32'hc3887b3e, 32'h43031151},
  {32'h4314bb12, 32'hc2da0b3c, 32'h42576bb7},
  {32'hc2b0af6c, 32'hc3c0fd10, 32'hc34653f0},
  {32'hc31c5d93, 32'hc3746eac, 32'hc2cc1288},
  {32'h421cd17c, 32'h420bc960, 32'h43e73b16},
  {32'h42fbffbe, 32'hc2d9de1e, 32'h42a7a1b3},
  {32'h42bbb16e, 32'h42ea49b4, 32'hc2d108b8},
  {32'hc2883ae6, 32'h42be1eff, 32'hc3a56477},
  {32'hc3a01bdf, 32'h434b0ca4, 32'h3fbb7ec0},
  {32'h4232ed35, 32'h4385b21b, 32'hc2c50ab1},
  {32'hc25253cb, 32'hc3a9626b, 32'hc39ae684},
  {32'h43007824, 32'hbe5f4300, 32'h434d4530},
  {32'h429bf80f, 32'hc286cb59, 32'hc2c8c068},
  {32'hc2f7ff40, 32'hc307fb32, 32'hc366bebe},
  {32'hc3501d8e, 32'h428d7363, 32'h43769282},
  {32'h43632b9f, 32'h418f5b99, 32'hc38dac3b},
  {32'hc3ee98f6, 32'h432b088b, 32'h43b9eb86},
  {32'h42a1dcc8, 32'hc37e4c0f, 32'hc394e6e5},
  {32'hc3413746, 32'h440075f1, 32'h42be2f05},
  {32'h43212679, 32'hc2e8e396, 32'hc2cb96d5},
  {32'h41ad641b, 32'hc37cc90f, 32'h43885ccf},
  {32'hc2ff8388, 32'hc3c259c5, 32'h43a34544},
  {32'hc305f06a, 32'h4301bc43, 32'hc2ecbd4e},
  {32'hc187cb40, 32'h43619e80, 32'h43146b68},
  {32'hc1914d83, 32'h43229a71, 32'hc303310b},
  {32'hc3bc3d18, 32'hc204241b, 32'hc374ef13},
  {32'h43e9aeae, 32'h440bde00, 32'hc1cb50e6},
  {32'h41e2974c, 32'hc1476c5c, 32'hc3c25620},
  {32'h417ed2a0, 32'hc38ed3bb, 32'hc31d8ba6},
  {32'h42f3218b, 32'hc39abc64, 32'h4415a907},
  {32'hc2b06530, 32'hc30ccf78, 32'hc2a5b49d},
  {32'h42e9e797, 32'h431b8ed0, 32'h431a1195},
  {32'h43cde9ed, 32'hc18ec912, 32'h40af51c5},
  {32'h43771b05, 32'hc19b7342, 32'h4425aaca},
  {32'hc25614e9, 32'hc327fde9, 32'hc2d241a5},
  {32'h43306a21, 32'h43590e36, 32'hc342ae45},
  {32'h409e390b, 32'h43a8e4e3, 32'h436c6123},
  {32'hc362c0ff, 32'hc114e735, 32'h434cac5f},
  {32'h441bdec2, 32'h435c1fff, 32'hc38f2134},
  {32'h3f824d70, 32'hc33b0039, 32'hbfe7ea14},
  {32'h429699c9, 32'hc203d7a4, 32'h431fca31},
  {32'h43141a9e, 32'hc3985968, 32'hc3d24544},
  {32'hc3d5d573, 32'h4313c7be, 32'hc2e762f3},
  {32'hc3ab1f5c, 32'h437ac33c, 32'h4418b854},
  {32'hc304258f, 32'hc25ffbf9, 32'h437c0ddb},
  {32'h428f2079, 32'h43cbe02b, 32'hc3898c4d},
  {32'hc2bd1236, 32'hc308111c, 32'h43b2b7ba},
  {32'h43197a65, 32'hc2b6700e, 32'hc3994cd1},
  {32'h422c86da, 32'h42d735d8, 32'h439ada71},
  {32'hc30a7f1c, 32'h41c42e30, 32'h43a63c35},
  {32'hc0c473e0, 32'hc321555b, 32'h442ef7e4},
  {32'hc4015abb, 32'h438437dd, 32'hc4345f02},
  {32'h4393a606, 32'h432b1e08, 32'h40820860},
  {32'h43496a01, 32'hc2914c89, 32'hc318373c},
  {32'h4341e9d9, 32'hc3301e0f, 32'hc3290169},
  {32'hc3ae5845, 32'hc2af397d, 32'hc34e1d0b},
  {32'h4250861c, 32'hc3ba4383, 32'h41d6cb53},
  {32'hc30ffc79, 32'h42160a1c, 32'hc3476868},
  {32'hc3ba6cf5, 32'h433cf833, 32'h4338ed53},
  {32'h43aa5137, 32'hc36105c5, 32'hc38835a6},
  {32'h439ca8c0, 32'h439e5209, 32'hc3c7aec7},
  {32'h42cdbb2d, 32'hc1e62aa1, 32'hc295e8b3},
  {32'h42e45d62, 32'hc28373d7, 32'hc349d8b6},
  {32'hc32ad948, 32'hc3eb2022, 32'h43250984},
  {32'hc2f37a24, 32'h43e4a8ce, 32'h432cbcac},
  {32'hc31095b0, 32'h42019aeb, 32'h41e85252},
  {32'hc2fab065, 32'h42a0bd30, 32'hc2d39557},
  {32'hc376ff2a, 32'h430a565e, 32'hc3b8d5fa},
  {32'hc2888de8, 32'h4321d8f9, 32'h43a37378},
  {32'h438b51f3, 32'hc38b798f, 32'h4249f629},
  {32'hc3431a28, 32'hc1ab6068, 32'h4390e47b},
  {32'hc31df47b, 32'hc34b63cf, 32'hc2a255a4},
  {32'hc19977b2, 32'h4394ef9f, 32'hc3383ae4},
  {32'h435c29e5, 32'hc390ab83, 32'h42f702d4},
  {32'h42dd055d, 32'hc2e569d0, 32'hc419aa52},
  {32'h438b1b47, 32'hc1564b87, 32'hc3827d6f},
  {32'h430e3eb4, 32'h429cdda4, 32'hbeb2c700},
  {32'h431f918f, 32'h430e56fe, 32'h421d456a},
  {32'hc36bbb40, 32'h4398eafd, 32'hc38137bf},
  {32'h42315024, 32'h432cc0b1, 32'h4338522c},
  {32'h441cbb07, 32'hc32c8afb, 32'h4417c741},
  {32'hc24cce76, 32'h4385345b, 32'h42d7f2b4},
  {32'h42e87072, 32'hc18e235d, 32'h43c569c4},
  {32'h43941ae4, 32'hc353b288, 32'hc3695c3b},
  {32'h43458bc1, 32'hc204b2ba, 32'h4400b414},
  {32'h438b502a, 32'hc28254b0, 32'h436f2d06},
  {32'h4369e26e, 32'h42a80d76, 32'hc3efb0ca},
  {32'hc3e67eac, 32'h431ae63d, 32'h43fe53b8},
  {32'h430dc289, 32'hc1ff9b71, 32'h42ae737e},
  {32'h4371c2ab, 32'hc34e21dc, 32'hc3e24f5f},
  {32'hc3ce1d6e, 32'hc3f0ae42, 32'hc23b9c45},
  {32'h43356321, 32'hc40e7532, 32'h434230b2},
  {32'hc18f43a4, 32'h43a6e6e6, 32'h42f48e93},
  {32'hc3749d46, 32'h434b1df2, 32'h42b8cbbb},
  {32'hc359ca16, 32'h43b3d717, 32'hc3baf854},
  {32'hc2ae74ef, 32'h439e4843, 32'h430625bf},
  {32'h438a0066, 32'hc386614d, 32'hc2bba76e},
  {32'hc3a85a3c, 32'h42e8f36d, 32'h43da31fa},
  {32'h4429d27f, 32'hc1810675, 32'hc3e15dc7},
  {32'hc2cf0fce, 32'h43bbbbaa, 32'hc33546da},
  {32'hc3071f5e, 32'h42166a96, 32'h42f550bb},
  {32'h4228600b, 32'hc25da4ad, 32'hc3059c74},
  {32'hc3b7ee32, 32'hc2e1e629, 32'h430b4ec9},
  {32'hc402395c, 32'h438c4a67, 32'hc308b487},
  {32'hc1c23c4c, 32'hc3d6ff66, 32'hc2ac2782},
  {32'hc360554b, 32'h4380c186, 32'hc2c067a7},
  {32'hc30c839a, 32'h44175a54, 32'hc3d4e9b6},
  {32'h438d9c13, 32'h440ed683, 32'h4371089a},
  {32'hc18e6aee, 32'hc20891f5, 32'hc3a6a398},
  {32'hc2bc3db5, 32'h42f5aec6, 32'hc3bb4f22},
  {32'h443b095e, 32'hc08ccb40, 32'hc340170f},
  {32'h40ecc122, 32'h42a2507c, 32'h429b1457},
  {32'hc2e2789d, 32'hc34d61dc, 32'h42f2304a},
  {32'h439208a1, 32'hc3baf7f6, 32'hc3c68fb9},
  {32'hc3825181, 32'hc321784c, 32'h43e7f84d},
  {32'hc35af75e, 32'hc255c0e6, 32'hc32e5d7d},
  {32'h412f02d0, 32'hc2f0cb6a, 32'hc39cd0fb},
  {32'hc27b6253, 32'h442ac59e, 32'h444ebac9},
  {32'h412d60ca, 32'h40158077, 32'hc30f4486},
  {32'hc21fdb1a, 32'hc2bcfd00, 32'h4289227a},
  {32'hc394e7b5, 32'hc4092a48, 32'hc3c0540a},
  {32'hc3663906, 32'h4406a435, 32'h4396f7ad},
  {32'hc1e92884, 32'hc26c53a3, 32'hc33b0f7f},
  {32'h440b2089, 32'h42e4339d, 32'hc1b1007e},
  {32'hc2c50956, 32'hc2ae4c4a, 32'hc2a94c3b},
  {32'hc2fdd959, 32'h43cb713e, 32'h42dc4a8b},
  {32'hc1e157f3, 32'h43d826e3, 32'h439beb97},
  {32'hc3b27314, 32'hc30a433a, 32'h4313b471},
  {32'h4378224f, 32'hc34c818d, 32'h43959c01},
  {32'h425c7afe, 32'hc319e681, 32'hc3622b79},
  {32'hc29389cb, 32'hc2d4225b, 32'h41e9aa66},
  {32'h4351b88b, 32'hc3c18326, 32'h43bcc3e3},
  {32'hc33ce734, 32'hc32821a7, 32'hc1e307c1},
  {32'h4288ea9c, 32'h43abb80f, 32'h43983d85},
  {32'h43028159, 32'hc2fc1913, 32'h4382358c},
  {32'hc39c8bef, 32'hc32cb994, 32'hc3657c56},
  {32'h42591cd7, 32'hc3bb11be, 32'h43ca3b4c},
  {32'hc3830d46, 32'hc3549a84, 32'hc2db7446},
  {32'hc2c0e519, 32'h42b5045b, 32'hc35c83aa},
  {32'hc28fff59, 32'h4207bcc2, 32'h428f3cde},
  {32'hc212c36d, 32'h40f96f35, 32'hc38f5277},
  {32'h42ac81ea, 32'h43600e47, 32'h4348c29a},
  {32'hc35dd3d3, 32'h4384badb, 32'hc33989ef},
  {32'hc2de0b10, 32'h4382ee6d, 32'h428a6489},
  {32'h4342e1d9, 32'hc4276671, 32'h43ddc693},
  {32'h42dcb032, 32'h4333cf1d, 32'h43640e56},
  {32'h439ba371, 32'h426cbbb5, 32'hc3a23140},
  {32'hc32b3327, 32'hc35e03f6, 32'h43b84c4a},
  {32'hc3912785, 32'h43ba1a03, 32'h438a5598},
  {32'hc2cefa38, 32'h440f20ca, 32'h43d7abe8},
  {32'hc387875b, 32'hc384c91e, 32'hc3909754},
  {32'hc37a85a2, 32'hc2b4355a, 32'hc35697e8},
  {32'h42969328, 32'h4389d2f1, 32'h42b5172e},
  {32'hc38679e8, 32'h431a9484, 32'hc24617b8},
  {32'h41aa9104, 32'h4286a8d2, 32'h43b22ac6},
  {32'h42a2a234, 32'hc3dd06be, 32'h423c09fb},
  {32'h43e5fd2a, 32'hbff7ea8d, 32'hc2be58f3},
  {32'h43af52a8, 32'hc1dbfb08, 32'hc3d349e3},
  {32'h42725334, 32'hc3622c42, 32'hc3909ca7},
  {32'hc385d480, 32'h43a11b06, 32'hc209c961},
  {32'hc21c75f8, 32'h4369bb00, 32'h43818363},
  {32'h42cb2cc8, 32'hc2ff7410, 32'hc380f55d},
  {32'h42ce16a0, 32'hc34a4802, 32'hc3419389},
  {32'h4345cc98, 32'h43111cc1, 32'h420b0d36},
  {32'h43d2bfc2, 32'hc3bbdfcd, 32'h41155f74},
  {32'hc416a8ac, 32'hc3b946cc, 32'hc3cdfc11},
  {32'hc2698324, 32'hc2f2462b, 32'h43ca7fbd},
  {32'h4339afd6, 32'h41f8f25e, 32'hc3bfe14f},
  {32'hc3cc0203, 32'h433f9e11, 32'hc3d911bd},
  {32'h4386516e, 32'h43ed5ac6, 32'hc3297aac},
  {32'h433dfccb, 32'h4405490a, 32'hc3c62ee3},
  {32'h4110fa40, 32'h433697ed, 32'h42a27ede},
  {32'h42e87014, 32'h43279b46, 32'hc372ffb4},
  {32'h44028637, 32'hc2935aee, 32'hc35694f1},
  {32'hc39c39fe, 32'hc3ca1239, 32'h434e9300},
  {32'hc300eab6, 32'h41012781, 32'hc36b9912},
  {32'h41e928cf, 32'h4039e3d9, 32'hc3bb59a5},
  {32'h42a022fa, 32'hc377dfb4, 32'hc2948d67},
  {32'hc36fc65b, 32'h43a8a80d, 32'h42edc836},
  {32'h43a74d89, 32'hc36f23d7, 32'h426b770b},
  {32'h4212035f, 32'hc3ab1b25, 32'hc1813c82},
  {32'hc3571154, 32'hc319715a, 32'hc330d645},
  {32'h439fbf44, 32'h43203884, 32'h431fb194},
  {32'hc38da05a, 32'hc21e476d, 32'h409ebbbd},
  {32'hc388e9ad, 32'h43da4656, 32'h41b6bdce},
  {32'h43f6c08d, 32'hc30b3406, 32'h43bc8a41},
  {32'hc4062fd6, 32'hc395ad17, 32'hc0dbe75c},
  {32'hc3fa1eea, 32'h42a3469b, 32'hc413c641},
  {32'hc3e5f9e2, 32'h439e40a7, 32'hc26dcf40},
  {32'h432e5420, 32'h43b75920, 32'h427960f1},
  {32'hc19065cb, 32'hc320863e, 32'h41713baf},
  {32'h431b7cb8, 32'hc28e537b, 32'h41f76736},
  {32'hc2dfffd2, 32'h435a2870, 32'hc3b6fbaa},
  {32'hc399a423, 32'hc326bbfe, 32'h421cd1df},
  {32'h432034cd, 32'hc30fe1e6, 32'hc40c0781},
  {32'hc29bde8f, 32'hc3841677, 32'h43895036},
  {32'h43a79446, 32'h4318502f, 32'h43a4b66e},
  {32'h4404b353, 32'h43b9bfb1, 32'hc2783a1a},
  {32'h41fc9df4, 32'hc3d17cf8, 32'hc269e496},
  {32'hc2daf6cd, 32'hc2bbd028, 32'hc34f6331},
  {32'h41b33988, 32'hc110f2a7, 32'h423a189c},
  {32'h422274e3, 32'h42c70532, 32'h42463a8b},
  {32'h426bc2f2, 32'h435f9917, 32'h42466a88},
  {32'hc3570c3c, 32'hc2ea79a4, 32'h4269a471},
  {32'hc3d29103, 32'h4318bcb8, 32'h43d2682c},
  {32'hc3ee7f24, 32'h420f86d2, 32'hc375fd7f},
  {32'h42f7fc69, 32'h439b8117, 32'hc32916b7},
  {32'h43c82b27, 32'hc3464087, 32'h402f0424},
  {32'hc3ad4650, 32'hc2e8b6bd, 32'h437a9aae},
  {32'h4410e31c, 32'hc3c5a6d5, 32'hc31dfc6b},
  {32'hc2c2efba, 32'hc37e578e, 32'h42a6068c},
  {32'h430abdec, 32'h42acd29f, 32'hc3a4d7fc},
  {32'h4366f733, 32'h433d6242, 32'hc24810ce},
  {32'hc4009d21, 32'h422dd8f0, 32'hc294e63c},
  {32'h42ec217a, 32'h41cbbb46, 32'hc2e6dd62},
  {32'h4382d88f, 32'h435deecd, 32'hc34c33a8},
  {32'hc1b32076, 32'h433589d2, 32'hc3c1a11c},
  {32'h41b689c4, 32'hc2a31d72, 32'h42f232b2},
  {32'h433e8baa, 32'h43b1383a, 32'hc3005469},
  {32'hc391ec9f, 32'hc2cdfecc, 32'hc386e92e},
  {32'hc28fea57, 32'hc0badb3a, 32'hc0cf37a4},
  {32'hc3eb55aa, 32'h42fec651, 32'h43900589},
  {32'h42e5f802, 32'hc379c74b, 32'hc23d3915},
  {32'h40eaee4a, 32'h43169665, 32'h43bdea90},
  {32'h4277e1c7, 32'h44042fc2, 32'hc4230670},
  {32'hc3b39ba4, 32'hc352ac76, 32'h4281b7f1},
  {32'h433a5929, 32'hc1ac5b2a, 32'hc31b7f57},
  {32'hc246aac4, 32'hc3e97ecd, 32'h430eb603},
  {32'hc39b1b3b, 32'h4384cabc, 32'hc3b15e21},
  {32'hc3af25ac, 32'h4307c8b0, 32'hc2cd50ba},
  {32'h43095ce8, 32'h431db15b, 32'h43e5db9d},
  {32'h436112e2, 32'h4325b178, 32'h439d2000},
  {32'hc2506256, 32'hc39468a5, 32'h437e5bfc},
  {32'h442d5112, 32'h4380cf8c, 32'hc308c6e0},
  {32'hc3057d7a, 32'hc3c643d5, 32'hc24a1414},
  {32'hc3a2b8e7, 32'h435ccb7a, 32'h43a23ff4},
  {32'hc3659c6d, 32'h435b3935, 32'h423ff650},
  {32'h42efc787, 32'h43160365, 32'h437000a3},
  {32'hc3a38422, 32'hc38453c9, 32'h4282519c},
  {32'h440e2636, 32'hc3692828, 32'h4371b018},
  {32'hc3b87aca, 32'hc3f5f8cf, 32'h4163276a},
  {32'hc32a52bc, 32'h444585e3, 32'hc3c8c031},
  {32'hc2b54339, 32'h441d52f5, 32'hc34d15cc},
  {32'hc275ef77, 32'h441443aa, 32'h419b731b},
  {32'h42e00985, 32'hc3a36355, 32'h435a06ef},
  {32'hc2662458, 32'hc3bab98a, 32'hc3459e1b},
  {32'hc402ac2a, 32'hc31a37c5, 32'hc3328321},
  {32'h4296250f, 32'h422ce4a1, 32'h42d44885},
  {32'h4258aa8c, 32'h432eeddf, 32'hc415efc3},
  {32'hc4361621, 32'h43a58a87, 32'h43b4fb2b},
  {32'h43c23fba, 32'h42427721, 32'hc26723c0},
  {32'h4334910a, 32'hc3db03b2, 32'hc2d61fb9},
  {32'h42cc4859, 32'h43be1882, 32'hc2b38d6c},
  {32'hc25e8392, 32'h42e7c112, 32'hc3a6cbe4},
  {32'h43ae04d6, 32'hc377afa4, 32'hc2192c18},
  {32'hc3e88826, 32'hc3f3aefa, 32'hc3f7daa2},
  {32'h4354fe37, 32'hc2cce9be, 32'hc3982a82},
  {32'hc399f428, 32'h4419a2ea, 32'hc30e454f},
  {32'hc384af77, 32'h43518f9e, 32'hc36153be},
  {32'hc3903904, 32'h43a3f0a5, 32'h440c2820},
  {32'h4374f1f2, 32'hc37809ec, 32'hc41f085b},
  {32'hc31f50b8, 32'hc3cdc4ff, 32'hc3ea05b5},
  {32'h42b08b0f, 32'hc331a0d3, 32'h42b56f74},
  {32'hc24cb19c, 32'hc2a36d06, 32'hc35e3776},
  {32'hc2f35f5f, 32'hc3ddd27a, 32'hc3a8d40c},
  {32'h436f31b0, 32'hc39d422d, 32'hc263c28a},
  {32'h43941901, 32'hc3815b94, 32'h442a682c},
  {32'hc3c49f1e, 32'h43cc8e13, 32'hc3bf4800},
  {32'hc4018364, 32'hc3496871, 32'hc3890669},
  {32'hc22626da, 32'h43c37d74, 32'h4373983d},
  {32'hc23d90d1, 32'hc26a0a06, 32'hc250c9e4},
  {32'h428b719d, 32'hc2b7aaf4, 32'hc35e8508},
  {32'h434511aa, 32'hc2dc0d41, 32'hc294ffe6},
  {32'hc309395e, 32'h433bf6bf, 32'h43992ab0},
  {32'hc357b658, 32'hc266d806, 32'hc2f616d5},
  {32'h439e0923, 32'h42519ce3, 32'hc3132557},
  {32'h443b0994, 32'h4387d2e2, 32'hc2a14372},
  {32'h43303389, 32'hc356ca1b, 32'h4332c983},
  {32'h4324033b, 32'h42859582, 32'hc2f38bd0},
  {32'hc3d628d6, 32'h430b2f82, 32'h42f79bd2},
  {32'h43d47377, 32'hc34d4072, 32'h438b391c},
  {32'h43f150d6, 32'h4389d6cf, 32'h42ab5ff8},
  {32'h432959ff, 32'hc3df2955, 32'hc3cfe060},
  {32'hc3a79e1a, 32'h4318dd47, 32'hc322f0d0},
  {32'h42a87bb0, 32'hc174ad61, 32'h42c5e409},
  {32'hc19de6e9, 32'h42314c3b, 32'h42f7afda},
  {32'h43bd1804, 32'h43436878, 32'h41872313},
  {32'hc31bcd17, 32'h42e89f2e, 32'hc38a72eb},
  {32'hc39182dd, 32'hc390c8ab, 32'hc2ffec84},
  {32'hc36f1a9b, 32'h40a14234, 32'h41e9538e},
  {32'h43897d93, 32'hc2df2760, 32'hc34db1a5},
  {32'hc3c4ab4d, 32'hc334da0d, 32'h43818e55},
  {32'hc40068f4, 32'h43a063c4, 32'hc2fca0c8},
  {32'h43af08f7, 32'hc3c0d0d3, 32'h41fdff3f},
  {32'hc3e20c37, 32'hc3920f70, 32'hc3863dfa},
  {32'hc37f5658, 32'h434635bc, 32'h43763a42},
  {32'hc35e4014, 32'h4388e63b, 32'h4319a480},
  {32'hc38005b7, 32'hc34210bc, 32'h4150324a},
  {32'h4333171b, 32'h4247d737, 32'hc2a37810},
  {32'h434434e9, 32'hc387c2ab, 32'h4383e50e},
  {32'h41b1d346, 32'hc3af445c, 32'h43435326},
  {32'hc219087e, 32'h431e3954, 32'hc29645b3},
  {32'h4332a042, 32'hc2d38653, 32'hc3ca9a13},
  {32'hc32e4c65, 32'hc14c1de1, 32'hc2edd746},
  {32'hc349735d, 32'h41b757d3, 32'h417638ea},
  {32'hc3f8e552, 32'hc3080ab9, 32'hc27b59c6},
  {32'h42d756a5, 32'hc3b8e043, 32'hc26aaf25},
  {32'h42d35784, 32'h43020119, 32'hc3544a0d},
  {32'h4333a73a, 32'hc33ef914, 32'hc416133f},
  {32'hc44a4aac, 32'hc2c6309b, 32'hc27cc914},
  {32'hc33308c3, 32'hc2b39b92, 32'hc21901da},
  {32'h433b380a, 32'h43434a32, 32'hc3ca0e2d},
  {32'hc2d86368, 32'h42d5a1df, 32'hc2063a83},
  {32'hc3379c92, 32'h43cd2fec, 32'h43cba233},
  {32'h43c9a79c, 32'hc1b83e81, 32'h43ad2e30},
  {32'hc27c75a4, 32'h42d85b71, 32'hc41d5df8},
  {32'hc3cebdc7, 32'h43ebf675, 32'h42071b1e},
  {32'h43b00f72, 32'hc2069175, 32'hc38f90e4},
  {32'hc38dc29e, 32'h431300f3, 32'hc388b219},
  {32'hc3a524ab, 32'h43809200, 32'hc2acb20c},
  {32'h41b39090, 32'hc105374f, 32'h43936f11},
  {32'hc3ab156b, 32'h439e5a4a, 32'hc381b947},
  {32'hc3d5fd02, 32'hc1a730a4, 32'h43db285c},
  {32'hc24b9058, 32'h420c7f39, 32'h41618e7c},
  {32'hc39872b6, 32'h43bd3db1, 32'h43366c88},
  {32'h41bf4b51, 32'h42b9db1e, 32'h42c4b827},
  {32'h43827e8a, 32'hc2e89e9d, 32'hc120b8e9},
  {32'h434f85ea, 32'hc3135083, 32'hc2a233a3},
  {32'h4381d77a, 32'hc31897f8, 32'hc384b40d},
  {32'h43974f8c, 32'h43038414, 32'hc37ddaa6},
  {32'h437a4896, 32'h42c41a20, 32'h440e18a4},
  {32'h43efefce, 32'h43694d47, 32'h438a74f2},
  {32'hc13dcabd, 32'h424f1374, 32'hc30ae9cb},
  {32'hc360103e, 32'h43a6c587, 32'h43209480},
  {32'hc3b4c57f, 32'hc1d253cd, 32'h42eda5a9},
  {32'h436ac9e0, 32'hc39f1680, 32'hc3cd26cf},
  {32'hc3bf6903, 32'h42de4add, 32'h42992855},
  {32'hc39c676c, 32'h43a4fb6e, 32'hc38ddf1a},
  {32'h42bd95cd, 32'h4389478b, 32'hc3ccd86e},
  {32'h43887106, 32'h4301630c, 32'hc2c8f830},
  {32'h424587dc, 32'hc2fa275e, 32'h42ee17c2},
  {32'hc2a3f409, 32'hc3fc383b, 32'h435e389d},
  {32'hc4199567, 32'h43e9b721, 32'hc309f9a3},
  {32'hc41c0393, 32'hc071658e, 32'hc264d45f},
  {32'h434c17ce, 32'h4211b2b8, 32'h43b9d699},
  {32'hc32e5c27, 32'hc3a4093a, 32'h4390c79f},
  {32'hc30b207c, 32'hc30357a3, 32'hc1ffd9e9},
  {32'h44086244, 32'hc2c55471, 32'h440d51a6},
  {32'hc2d0fdef, 32'h41ebad98, 32'hc1681411},
  {32'h44030308, 32'h42099b71, 32'h43aa20da},
  {32'h438713ba, 32'h437b0aa7, 32'h43982a53},
  {32'hc3954169, 32'hc26a6081, 32'h4308cbfc},
  {32'hc3a71132, 32'hc398ece7, 32'hc1da41ae},
  {32'h43428ca3, 32'hc391b9bf, 32'hc2df4224},
  {32'hc2bc7f6b, 32'hc3a47e81, 32'h43a3914f},
  {32'h428a6ddf, 32'hc2c958af, 32'h4371ffb0},
  {32'hc20e7fe1, 32'hc3e331d1, 32'hc3298b41},
  {32'hc375b947, 32'h4300897a, 32'h43bbaa3b},
  {32'hc28b49e7, 32'hc35946fd, 32'h433c676a},
  {32'h43b8fc49, 32'h42d0aa10, 32'h42ce3a6d},
  {32'h43604a22, 32'hc2be15b1, 32'h42ed1efa},
  {32'h43c629fb, 32'h40b164b7, 32'hc380347b},
  {32'h43ddb42a, 32'h41f3c517, 32'hc406ccad},
  {32'h41206e89, 32'h429c1517, 32'hc3445212},
  {32'hc265775a, 32'h430b35c5, 32'h43653062},
  {32'hc23ab136, 32'hc34979e3, 32'hc2cb0e91},
  {32'h423c3c42, 32'h433e913a, 32'h42b2787d},
  {32'hc372609c, 32'hc30b9a5b, 32'h4358712b},
  {32'h42cb6172, 32'hc255532a, 32'h442194a3},
  {32'hc3676f7e, 32'h43d4180f, 32'hc3a1276c},
  {32'hbe76e184, 32'h43b53fdd, 32'hc3ada0a6},
  {32'h4395347e, 32'hc28c66a4, 32'h437ae1a7},
  {32'h42e94e5a, 32'hc347177a, 32'h433ba26a},
  {32'hc2a9359c, 32'h4275815e, 32'h4304127f},
  {32'h4441af1e, 32'hc25af9b8, 32'h447cb871},
  {32'hc3ad28b4, 32'h43682ec4, 32'hc2fff832},
  {32'h43131efb, 32'h436fe1d2, 32'hc2e805c4},
  {32'h439208a4, 32'hc2821374, 32'h438ed95f},
  {32'h42d7d3bc, 32'h43736641, 32'h42bffb6e},
  {32'h42b165b0, 32'hc33cad3b, 32'h436ec4c1},
  {32'hc12f422a, 32'h43912c54, 32'hc341b52a},
  {32'hc2f9fbb4, 32'hc2a52c76, 32'hc362354d},
  {32'hc39bc2a5, 32'hbfb05fa2, 32'hc3482069},
  {32'h42c166dc, 32'h438f76bc, 32'hc3176372},
  {32'hc3356890, 32'hc2ca7076, 32'h436ddb63},
  {32'hc2a23e77, 32'hc32eeea0, 32'h411f8e41},
  {32'hc2d45f46, 32'h429051ae, 32'hc340bc0d},
  {32'hc3487958, 32'hc3808e93, 32'h430b91f6},
  {32'hc2afb891, 32'hc2ef31c7, 32'hc42ca226},
  {32'h4386f906, 32'hc3d15f55, 32'hc3e5c232},
  {32'hc3d11248, 32'hc353838d, 32'hc1d924a7},
  {32'hc2a768c4, 32'h432013c1, 32'hc3a303db},
  {32'h42974b32, 32'h4367aa65, 32'hc380fbc8},
  {32'h434ed015, 32'hc1b4fa00, 32'h43acf847},
  {32'hc3010330, 32'h43187255, 32'h42efd6a5},
  {32'h4354c2e1, 32'hc29057c7, 32'hc2111485},
  {32'h438e5f29, 32'h42f2bae1, 32'h40f7d11a},
  {32'h43ab2606, 32'hc3430d98, 32'hc375f259},
  {32'h4351a922, 32'h421ac75d, 32'h42ae4610},
  {32'hc3d53ae0, 32'hc26f61e4, 32'h43aae79d},
  {32'h42c8d7ab, 32'h440d6342, 32'hc3177876},
  {32'h438be2a8, 32'hc397f78a, 32'hc35cf180},
  {32'hc3944870, 32'h433a2abe, 32'h424287ca},
  {32'h40a2c9b2, 32'h43581c90, 32'h43cbbdc4},
  {32'h4347756b, 32'h43b7f7fc, 32'hc308616d},
  {32'hc27f3929, 32'h4319b2a2, 32'hc29c79ee},
  {32'hc356af4b, 32'hc398b10a, 32'hc2dbf5a0},
  {32'h439a42e0, 32'hc25646d3, 32'h43bd9003},
  {32'h42a52a03, 32'hc374d468, 32'h43974bd0},
  {32'hc320cdd7, 32'hc429e33a, 32'h4246a3e1},
  {32'h4327c5d3, 32'h435d5a40, 32'hc0a15204},
  {32'hc342fe6e, 32'h42ed9b56, 32'hc2b8b7ab},
  {32'h43957366, 32'hc1564f79, 32'h43a1e844},
  {32'h42a8d94e, 32'hc28d711c, 32'h3faa0efd},
  {32'hc3d3a400, 32'h440d5111, 32'h43308e22},
  {32'h42db6dd4, 32'hc0bddd60, 32'hc3c13953},
  {32'h43e3bb8b, 32'hc307daac, 32'hc303bd8e},
  {32'hc2892334, 32'hc2c8ff72, 32'h43b80d4c},
  {32'h4387e43a, 32'h419b9e0b, 32'hc3857000},
  {32'hc39603c2, 32'h43c51f6a, 32'hc3774ccc},
  {32'hc3bdb5b8, 32'h42a356ea, 32'hc305e980},
  {32'h42ab161a, 32'h42e62a20, 32'hc2661505},
  {32'hc2f2abd7, 32'hc2b8655e, 32'hc16ed0c6},
  {32'hc3842c8d, 32'hc3963f1e, 32'hc385067b},
  {32'hc3dea519, 32'h42f0294e, 32'h4407425b},
  {32'h431e0105, 32'h4159045e, 32'h41f21982},
  {32'hc34e1dd0, 32'hc2454a86, 32'h42832e6f},
  {32'hc39ab3a0, 32'h429a6a3e, 32'hc37ea854},
  {32'hc1fd0f30, 32'hc2345d2c, 32'h439837e6},
  {32'hc29c4e30, 32'h4407bde5, 32'hc4085e6a},
  {32'h41479c90, 32'h431fc37f, 32'h43ea7442},
  {32'hc31c03cc, 32'h43d8407d, 32'h42c928f6},
  {32'hc3a31ffc, 32'hc2fe7c89, 32'hc206d7d5},
  {32'hc3e14503, 32'hc3c01ab6, 32'h432b16ce},
  {32'h43a06b1a, 32'hc33f31a9, 32'hc32bae9d},
  {32'hc2b7cfee, 32'hc3d21417, 32'h4291d2a7},
  {32'hc39f50a9, 32'hc32a6bf8, 32'h425af09a},
  {32'hc29f2781, 32'h43a3ec82, 32'hc344c716},
  {32'hc37647f7, 32'h41dcf969, 32'h42efab0b},
  {32'h436b8f82, 32'h437737a3, 32'h43ec4b1e},
  {32'hc2e5c74e, 32'h419f6226, 32'h42faf840},
  {32'hc430293c, 32'h44046d83, 32'hc3976bcf},
  {32'h41bfcef8, 32'h4377945a, 32'hc4249cd1},
  {32'h43b07a84, 32'hc373db7a, 32'hc37514ec},
  {32'hc33d599f, 32'hc4074274, 32'h432cf933},
  {32'hc2cb7dd8, 32'hc26a3db3, 32'hc3058083},
  {32'h42a04444, 32'h4231a710, 32'h43accaec},
  {32'hc2d2a4c2, 32'h43a52f68, 32'hc355396a},
  {32'hc3165b17, 32'hc2ed9130, 32'hc3602730},
  {32'h44692914, 32'h43ec6e48, 32'hc3470d24},
  {32'h431c5ecb, 32'h43a2dbd0, 32'hc2293d56},
  {32'hc31b9238, 32'hc2d806f2, 32'h43981386},
  {32'h43551974, 32'hc20869e4, 32'hc385af3e},
  {32'h43716a39, 32'hc2ab423e, 32'h42b33ecc},
  {32'hc4146316, 32'h42b253d3, 32'hc432271c},
  {32'h4405912c, 32'hc2c070fc, 32'h443a9749},
  {32'h431921bf, 32'hc120b90a, 32'hc3ba1c42},
  {32'hc3a8ac86, 32'h429a448d, 32'h4340fd5d},
  {32'hc1ae03e0, 32'h4360d9d6, 32'h42243006},
  {32'h4328ac93, 32'hc2a99de8, 32'hc2ffeebf},
  {32'h436c9c4e, 32'hc383ea33, 32'h42df4a37},
  {32'h425e0c7c, 32'hc3d0c53d, 32'h431052a7},
  {32'hc42d422e, 32'hc3be3b1a, 32'hc332af40},
  {32'h42731630, 32'hc22449b2, 32'hc14b28af},
  {32'hc2ad3cf2, 32'h4301a9bd, 32'h43535667},
  {32'h438a3279, 32'h43a01a5b, 32'hc3a6aba4},
  {32'h43103967, 32'hc2688479, 32'h421e981b},
  {32'hc3369200, 32'hc39caade, 32'h43a3443f},
  {32'h43cdd403, 32'h43724be9, 32'hc2240d22},
  {32'h438b7c50, 32'hc2acc785, 32'h4288fefc},
  {32'h433d5011, 32'h42826f77, 32'hc401befa},
  {32'hc31ca357, 32'hc2b7c175, 32'hc300929e},
  {32'hc3a06894, 32'hc3f679e4, 32'hc2cd01e7},
  {32'h43b92820, 32'hc318eecb, 32'hc36bf98b},
  {32'h4287d6ad, 32'hc25ab369, 32'h4389b9da},
  {32'hc3ca7683, 32'h42ead07b, 32'h43603bda},
  {32'h431dd18f, 32'h426593cc, 32'hc35f0b65},
  {32'hc22d226b, 32'h42f85c9b, 32'h4392cb54},
  {32'hc353c1aa, 32'h42dbd15f, 32'hc2d6404c},
  {32'h431bd967, 32'h433f38b8, 32'h43b1bc72},
  {32'h432536df, 32'h4389e0cc, 32'h3fd9d850},
  {32'h416f6aa0, 32'hc23b8d38, 32'hc230d9f0},
  {32'h42f3a546, 32'h432d3735, 32'h43b4f9db},
  {32'hc38b0878, 32'h433a44f3, 32'h429e208a},
  {32'hc3074ce6, 32'h420991f1, 32'hc3160f6c},
  {32'h442796d6, 32'h44432623, 32'hc38b7577},
  {32'hc469e60f, 32'h43e1d035, 32'hc26fd94e},
  {32'hc227df81, 32'hc3e8f01e, 32'h44280cfb},
  {32'hc2bce917, 32'h43fb250a, 32'hc374a67f},
  {32'h4320d23c, 32'hc1dabfe6, 32'hc3874c4d},
  {32'h42d5111f, 32'hc2bee68b, 32'h42ff7b61},
  {32'hc3a93a12, 32'hc2ce1c14, 32'hc3186fd1},
  {32'h43429f40, 32'h43e92ad6, 32'h43b85fc7},
  {32'h425b750c, 32'h442bb473, 32'hc3a12fae},
  {32'hc2a4e4ec, 32'h4324dbbd, 32'h434927be},
  {32'hc38d429e, 32'h4317f7cb, 32'hc2b91291},
  {32'h42f74d83, 32'hc3ad7302, 32'hc2a9bea0},
  {32'h434e05a2, 32'hc2085a8b, 32'h42ff5755},
  {32'hc3c5bb63, 32'hc17a0149, 32'h430c12a5},
  {32'hc1f7319c, 32'h43db4254, 32'h4396283a},
  {32'hc29c408a, 32'h43d7345b, 32'h4212d7b8},
  {32'h43a1d752, 32'hc3cf2a27, 32'hc3bc4854},
  {32'h431f493c, 32'hc24d3897, 32'h43a47401},
  {32'h43b17134, 32'hc2fe3dc5, 32'h434d5e4e},
  {32'hc33e52d9, 32'hc2c6f8c6, 32'h4387590c},
  {32'hc3984156, 32'h43022bb5, 32'hc3ef00bb},
  {32'hc326b07b, 32'hc3644349, 32'h42b6d0d8},
  {32'h430192df, 32'hc3c363d3, 32'h4397bfec},
  {32'hc393fb78, 32'h43273361, 32'hc2c36cdf},
  {32'h442db9f8, 32'h42ca8c8c, 32'h442fc750},
  {32'h43646480, 32'hc3433e04, 32'hc282c6c2},
  {32'hc304eab6, 32'h43ee41d3, 32'hc40fe45f},
  {32'h436e5e6d, 32'h4283d018, 32'h41bb50de},
  {32'h431c8a03, 32'h43033dd7, 32'h42bbcce0},
  {32'h41b04a63, 32'h438b8e3e, 32'hc346d0ac},
  {32'h43733aa0, 32'hc2efb969, 32'hc322fe69},
  {32'hc2d42870, 32'hc3755156, 32'hc2e6c0fc},
  {32'hc394addc, 32'h4326b678, 32'h4284cb7d},
  {32'h43bbb344, 32'hc21cbf86, 32'h42313626},
  {32'h423d30e3, 32'h439298cd, 32'hc3b6b2e8},
  {32'h42ab351d, 32'h43021172, 32'hc3a060a8},
  {32'h43be2823, 32'h43b1bc13, 32'hc3c314e6},
  {32'hc3bea547, 32'hc3427223, 32'h42e13b1e},
  {32'hc3b7cda0, 32'hc1c1fa95, 32'hc2d1c710},
  {32'h4216cc54, 32'hc35968a6, 32'hc3082aa0},
  {32'h43165b52, 32'hc263277c, 32'hc2ae7dac},
  {32'hc31661b0, 32'hc2e6f86e, 32'h4216c0f8},
  {32'hc25a5912, 32'hc2019a4a, 32'hc3172fde},
  {32'h43c5b660, 32'h44066ec1, 32'h42e61fd5},
  {32'hc2715eec, 32'h438cba8d, 32'hc2e88d9a},
  {32'h43c490bf, 32'h4311f799, 32'hc2804280},
  {32'hc3b03d27, 32'h4403d169, 32'h42d6d32d},
  {32'hc349fcfd, 32'h42223903, 32'h436b0e1c},
  {32'h433082b4, 32'hc2b5e798, 32'h43980ca8},
  {32'hc450e0ad, 32'hc33fecbd, 32'h43524b84},
  {32'hc32dc092, 32'hc19c535f, 32'hc3083258},
  {32'hc2ac3980, 32'h430fef2e, 32'h4359a828},
  {32'hc3939b78, 32'hc316a68d, 32'hc28190c5},
  {32'h414ac54d, 32'hc34e150e, 32'hc37b873b},
  {32'hc34e36ae, 32'h43cd96eb, 32'h42bab388},
  {32'h42e72f1f, 32'hc35c0e2b, 32'hc2332f35},
  {32'hc20eccae, 32'hc2cf5216, 32'hc35daee8},
  {32'hc3675b87, 32'h43868b77, 32'h4385d172},
  {32'h42e8259a, 32'hc403e3f2, 32'hc2821d29},
  {32'h434e5a71, 32'h41b5dbb4, 32'h440fce32},
  {32'hc319c487, 32'h436d745f, 32'h42bcf08c},
  {32'hc43f2c31, 32'hc3cec8f0, 32'hc33c966f},
  {32'h433e2c86, 32'hc2a5bb96, 32'hc1918726},
  {32'hc2932e0e, 32'h42efdf66, 32'h43697cf2},
  {32'h44076685, 32'h43b78de8, 32'hc3b2f083},
  {32'h4286e63e, 32'hc2ae683b, 32'h417e6f58},
  {32'h43c41b01, 32'hc398e1f1, 32'hc3209f23},
  {32'hc31e37b3, 32'hc3060d6c, 32'hc3b4b4cf},
  {32'hc1d8ffb9, 32'h426fd3ca, 32'h430eb3dd},
  {32'h435f0301, 32'hc36d526c, 32'hc2e947a9},
  {32'h43464850, 32'hc3082598, 32'h433a5902},
  {32'hc3b4e212, 32'hc2bf8c28, 32'hc1495bd6},
  {32'h43e3f6ef, 32'h4288b7b3, 32'h42ce397a},
  {32'h438af09b, 32'h42579471, 32'hc3b36dd4},
  {32'hc30c4fb2, 32'hc438cd9c, 32'hc3d75940},
  {32'h43639eba, 32'h4315da28, 32'hc3c2e554},
  {32'h425c9f92, 32'hc3c405ee, 32'h4340823f},
  {32'h43e6efd2, 32'h42ace2a9, 32'h42e91aae},
  {32'h41c7164d, 32'hc3909d9e, 32'hc31770cc},
  {32'hc3d9d6ac, 32'hc31098d5, 32'hc307725c},
  {32'hc425da3e, 32'h41bc971f, 32'hc334cc4b},
  {32'hc2d17308, 32'h43df6464, 32'h43b02266},
  {32'hc3116156, 32'h42ce563a, 32'h42ecde9b},
  {32'h4235b688, 32'h431d281d, 32'h434c79d5},
  {32'h43a4f9a6, 32'hc3b5c77b, 32'h43823b19},
  {32'hc38f93ea, 32'h42d90f0c, 32'h4292ba94},
  {32'hc3366ab0, 32'h41c5e8e9, 32'h42ce1dd8},
  {32'h43c3220c, 32'hc387a6a8, 32'h42ca54fc},
  {32'hc3fe088c, 32'h4228bb0e, 32'h43f19ffe},
  {32'h423ea710, 32'hc2e364eb, 32'hc2707b80},
  {32'h429c22dc, 32'hc220a6e7, 32'h43272d2a},
  {32'h44117498, 32'hc33bfae2, 32'h40b1d368},
  {32'h434307bc, 32'h43eba28a, 32'hc2e455d6},
  {32'h439f63ca, 32'hc22bfb8f, 32'h438038c5},
  {32'hc2dafc84, 32'h43a7a56a, 32'hc34c7856},
  {32'hc3a86e4a, 32'h439619a0, 32'h4281f96e},
  {32'hc32aff2b, 32'h42855ba3, 32'hc3c30c8e},
  {32'hc2cd336b, 32'h429183df, 32'h42ec6f98},
  {32'h4362d8e4, 32'hc34c4875, 32'h4352601b},
  {32'h43ed2be4, 32'h43965e2e, 32'h43841f72},
  {32'hc412f7b9, 32'h430241d2, 32'h42fb6261},
  {32'hc3801452, 32'hc29c2fff, 32'hc224bad7},
  {32'h43bb209c, 32'hc1e45b51, 32'h432a6836},
  {32'hc326345a, 32'h4305b345, 32'h43925f92},
  {32'hc24b18f6, 32'h43d91a49, 32'h42807e4a},
  {32'h441aff38, 32'h430f1fb0, 32'h44848c53},
  {32'hc2c4a9d4, 32'hc331f6d7, 32'hc3228526},
  {32'h42890d4e, 32'h440b54ee, 32'hc3de6be7},
  {32'h42ac9e8b, 32'h43a8d24c, 32'h43809a84},
  {32'hc396d4b5, 32'hc31ae319, 32'hc1afb60f},
  {32'h43460064, 32'hc2b74a4f, 32'h4384a7b0},
  {32'hc2bf9938, 32'hc34917b5, 32'hc27efd7a},
  {32'h4301fae8, 32'hc397eb05, 32'h42028432},
  {32'hc2a3747d, 32'h437bd868, 32'hc3004609},
  {32'hc4077a32, 32'h428e3efd, 32'hc22dc51a},
  {32'h42ca0dd0, 32'h432d3edd, 32'hc3a0fa54},
  {32'hc39d9033, 32'hc178fa9d, 32'hc1509d88},
  {32'h432ddf87, 32'hc384e395, 32'hc32b0525},
  {32'hbf370a00, 32'h40760a40, 32'hc30f178d},
  {32'hc2e0b3a5, 32'hc37fdd29, 32'h426ce4f3},
  {32'h43af4de6, 32'hc2d3406a, 32'hc2908274},
  {32'hc0ef7a1a, 32'hc240908a, 32'hc3e80604},
  {32'hc1e3f7fc, 32'hc396800f, 32'hc2a02e96},
  {32'h4298851a, 32'h425f8c01, 32'h43368a2b},
  {32'h434a10b1, 32'h40c6cac9, 32'h43b9263a},
  {32'h41cef2d6, 32'h431ec793, 32'h439fa438},
  {32'h433d3f76, 32'h4339c826, 32'h4412bfec},
  {32'hc38f8a59, 32'hc2adcc63, 32'h42a33973},
  {32'hc23f3ed4, 32'h42e03506, 32'h43e6fac9},
  {32'h43fefdf8, 32'hbfd06a56, 32'hc2e8122e},
  {32'h43b7cc6a, 32'h42229d81, 32'hc3526dc0},
  {32'hc300a5b1, 32'hc31bb712, 32'hc23ffdf4},
  {32'h4414b9c3, 32'hc0e50cc8, 32'h44112b1a},
  {32'hc3be8e91, 32'h43ec588d, 32'hc3983aec},
  {32'hc37a1c32, 32'h43bf6e67, 32'hc406198a},
  {32'h430a576c, 32'h42582d58, 32'hc31e8bb0},
  {32'hc1991169, 32'hc2b1b78b, 32'hc3d1f79a},
  {32'h43c29df6, 32'h434b1023, 32'hc10edba8},
  {32'h43435a5e, 32'hc2fe992b, 32'h4356d965},
  {32'hc3e9fe51, 32'h43428ead, 32'hc38a3a63},
  {32'h43c45e0f, 32'h4412ff0c, 32'h42a2e54c},
  {32'hc2d8f244, 32'h419788f9, 32'hc24506f7},
  {32'hc3b27bb3, 32'hc213b125, 32'hc373d918},
  {32'h43b022d1, 32'h440faac6, 32'h43785a83},
  {32'hc4068abb, 32'h4363a4c4, 32'h44137016},
  {32'hc321320c, 32'hc361653b, 32'h439182e4},
  {32'hc11522c0, 32'hc38b159e, 32'hc399e9a6},
  {32'hc2acf95b, 32'hc341debe, 32'hc190dd8b},
  {32'hc336b390, 32'h426165f0, 32'h42945c2e},
  {32'hc1b6cbc0, 32'hc2c2ebee, 32'hc404f475},
  {32'h435aaeda, 32'hc35acbfd, 32'hc3b22692},
  {32'h42e05ade, 32'hc395cb21, 32'h437d6492},
  {32'hc3106886, 32'h43d874b4, 32'h43f1429b},
  {32'hc268b92c, 32'hc37c9802, 32'hc30906b6},
  {32'hc2e0c72a, 32'h43a41429, 32'h433ad1f2},
  {32'hc40f7c14, 32'h43af171d, 32'h4401638e},
  {32'h439ef850, 32'h43aa9e17, 32'h43ff50d9},
  {32'hc273a281, 32'hc4246d64, 32'h43cbe83a},
  {32'h437eb004, 32'hc394da18, 32'h44183ffb},
  {32'hc1df8c3c, 32'hc297501f, 32'hc37292c8},
  {32'hc40e6b84, 32'hc3aaae97, 32'h42846749},
  {32'h42910f19, 32'h4214520a, 32'hc321f2c8},
  {32'h430e3e54, 32'h43d05aba, 32'h425fcd98},
  {32'hc37b7169, 32'hc4459782, 32'h437cff0d},
  {32'h40d6d2bc, 32'hc252abbe, 32'h4376589d},
  {32'h43898da9, 32'hc3919f39, 32'h43596972},
  {32'hc3e5d482, 32'hc310a345, 32'hc266849f},
  {32'h3f8cad80, 32'hc331bba4, 32'hc0a81193},
  {32'h438af0ac, 32'h432fab39, 32'hc2df0163},
  {32'hc3556258, 32'hc381176f, 32'hc3245423},
  {32'h42bc5b83, 32'h43800c96, 32'h440bf206},
  {32'h42b258e9, 32'h42d0dd4d, 32'hc33f99ea},
  {32'hc30717d5, 32'h44327c4d, 32'h43c53a76},
  {32'h4107fc27, 32'h43a59165, 32'h43a23ea7},
  {32'h43c0d616, 32'hc355e711, 32'hc360bd95},
  {32'hc3fc5978, 32'hc401f38a, 32'hc31d5c76},
  {32'hc2ac96f9, 32'h42d16cfd, 32'h438c988b},
  {32'h435677e7, 32'hc390ee59, 32'h431ee3eb},
  {32'h4190df96, 32'h43f20f04, 32'h42bbe0c8},
  {32'h43b4dd93, 32'h42de4bd5, 32'h422763e9},
  {32'h42345088, 32'h4383b2c5, 32'h4384f227},
  {32'h43a7d5f2, 32'h435bbc57, 32'hc3a980fb},
  {32'hc33ccbb0, 32'hc3010227, 32'hc4072af8},
  {32'h43859a56, 32'h42cdec20, 32'h439f1cb2},
  {32'h43332204, 32'h4431454e, 32'hc30f1a5d},
  {32'hc38ed1c0, 32'hc42b9fcf, 32'hc3931288},
  {32'hc102e19c, 32'h4374167c, 32'hc1e26978},
  {32'hc38b9392, 32'h4157696a, 32'h42f56ed8},
  {32'h43d4eed1, 32'h4399994f, 32'h43dc484d},
  {32'h415d80a8, 32'h43c6f58d, 32'hc27a7d84},
  {32'hc32af1af, 32'h42bf0227, 32'hc399bb43},
  {32'h4361490c, 32'hc38bb5d6, 32'h4342b3f4},
  {32'h42954dc0, 32'h4388219b, 32'h42583a0c},
  {32'hc44a3ab4, 32'hc2addb4a, 32'h42fc15dc},
  {32'hc317c03d, 32'h43353144, 32'hc319b6ea},
  {32'hc3a1c983, 32'hc0c73602, 32'hc22ee08f},
  {32'hc3149249, 32'hc2fc78bd, 32'hc2dc470e},
  {32'h434e0185, 32'h43643e48, 32'h41eac0a4},
  {32'h42505cbd, 32'h43b8f7e4, 32'hc31b1bc2},
  {32'h42ed89c5, 32'h433d0f03, 32'hc2bb181e},
  {32'hc3e7ba36, 32'hc3b5b422, 32'h412260c9},
  {32'h43d52f27, 32'h42ab7a96, 32'hc3a50b25},
  {32'hc3e00226, 32'h42974f27, 32'h4107ffa7},
  {32'hc25cbb72, 32'h4325e99a, 32'hc1c61448},
  {32'hc3b28a4d, 32'h43490e6c, 32'h42883110},
  {32'h439dd275, 32'h4372ed39, 32'h44344670},
  {32'hc3a5fc3c, 32'h435e122d, 32'hc1c7d1f5},
  {32'h444fbcc0, 32'h43578400, 32'hc20c6453},
  {32'h41fe2b3a, 32'hc3437643, 32'h42e22e67},
  {32'hc3a6a3d0, 32'h433d65dd, 32'h439a5509},
  {32'h43964066, 32'h436fd0e8, 32'h432c2b83},
  {32'h432164a7, 32'h433bb638, 32'hc1859359},
  {32'h420dfe50, 32'hc38a14c7, 32'hc36d9c1d},
  {32'h43fa1b4f, 32'h430a4b3e, 32'h44208d0f},
  {32'hc3be64a5, 32'hc2ddead5, 32'hc2704cbd},
  {32'h42180702, 32'h42b4c93c, 32'hc347e10a},
  {32'hc22aed18, 32'h4412335e, 32'h41479c2e},
  {32'h43082f34, 32'h4363fe03, 32'h41334e6d},
  {32'hc3ada6df, 32'h425fa1c5, 32'hc30c324e},
  {32'h42aa7f24, 32'hc3fcc458, 32'h43eb72ac},
  {32'hc3f0945e, 32'h43a4df3e, 32'hc3259f21},
  {32'hc0942c0b, 32'h4311ccaf, 32'h430e1e7f},
  {32'h433c07b8, 32'h428b16af, 32'hc38bd302},
  {32'h43fa3db4, 32'hc34be0db, 32'hc2991f0d},
  {32'hc39dcedb, 32'hc3fb4d81, 32'hc3374332},
  {32'h43b8144b, 32'h43aa976c, 32'hc384be92},
  {32'hc399d04f, 32'hc3337034, 32'h43dfca26},
  {32'hc1303fd6, 32'h428a4b8f, 32'hc402419b},
  {32'h43566b5e, 32'hc3773ed0, 32'h43cd81a9},
  {32'h42dc02e7, 32'hc40416d4, 32'hc23bb0c5},
  {32'hc245dd2c, 32'h43968591, 32'hc31ccec8},
  {32'h43452edc, 32'hc392e461, 32'hc39c53e1},
  {32'hc2f7845a, 32'hc3abe778, 32'h417566c5},
  {32'hc3b24a07, 32'hc2f39022, 32'h43518467},
  {32'h4425659a, 32'hc1283f2d, 32'hc282b0f2},
  {32'hc391e718, 32'hc2b97859, 32'hc2669fb2},
  {32'h415b228e, 32'hc27ba0db, 32'hc3ddae13},
  {32'h439386e1, 32'hc355c95c, 32'hc3f72b1b},
  {32'hc3fd99c7, 32'h438b5e7f, 32'h4213572f},
  {32'h41065b96, 32'h43f020e9, 32'h42f74a9a},
  {32'h432461d6, 32'h42f03314, 32'h43db5195},
  {32'hc3182051, 32'h4372bb0e, 32'hc3937dfe},
  {32'h439f7d01, 32'h440a3a60, 32'hc3c4106d},
  {32'h4372798f, 32'h4362fa90, 32'hc2be6fec},
  {32'hc3ea9b38, 32'h43d47409, 32'hc3467555},
  {32'h42da2f87, 32'hc285dba2, 32'h43790c1c},
  {32'hc282ff44, 32'hc40eef39, 32'h432ca58c},
  {32'hc3d1e195, 32'hc3216b06, 32'hc1aa311f},
  {32'hc32485ab, 32'h40a8c918, 32'hc2881865},
  {32'h43ae027e, 32'hc348c90e, 32'h422eddb6},
  {32'hc29aadf5, 32'hc2ae49d0, 32'hc37483e6},
  {32'hc2d4325c, 32'h42ede738, 32'h43525d3e},
  {32'hc409b1a9, 32'hc39bb66a, 32'h428a917e},
  {32'h43a7790e, 32'h43bbdb90, 32'hc2d81d0a},
  {32'hc37eb2bd, 32'hc2032bd2, 32'hc26daafe},
  {32'h44091cbb, 32'hc35decab, 32'hc3202ffd},
  {32'hc41c80dc, 32'h42b64b21, 32'h4364816c},
  {32'hc3a96c20, 32'hc36896cb, 32'h41e26868},
  {32'h42f36c24, 32'hc38d6ee3, 32'hc40b7520},
  {32'h42ce5db4, 32'h439f305c, 32'h439414f0},
  {32'hc3c2766c, 32'h42aff035, 32'h44106787},
  {32'h43bab72b, 32'hc2c3e0aa, 32'hc32b005c},
  {32'h431cda2e, 32'h43031b74, 32'hc3a6836a},
  {32'h42869e6c, 32'hc29b727f, 32'hc38b9a25},
  {32'h43a085f2, 32'h43b0f22e, 32'hc3de4fd5},
  {32'hc3b394c6, 32'h425f3644, 32'hc397e400},
  {32'hc14dcb8a, 32'h427af379, 32'hc2d033f3},
  {32'h4321ce8c, 32'hc30ce6f1, 32'hc30ba47e},
  {32'hc3be7c74, 32'hc363cbef, 32'hc2726cc6},
  {32'hc40b75a4, 32'hc21cb902, 32'hc3e1da09},
  {32'h4304a7ca, 32'h4398ab7e, 32'hc30db08e},
  {32'hc353f176, 32'h44848cce, 32'hc37ae77c},
  {32'h43344b5e, 32'hc29ae06a, 32'h42c38a72},
  {32'hc35d71d1, 32'h43803f9a, 32'h42d87a75},
  {32'hc3f65e15, 32'h4132d1b8, 32'hc352cbcb},
  {32'h4280be60, 32'h41a79ef6, 32'hc1f40cdb},
  {32'h4347c6ba, 32'h43b169e5, 32'hc391fc26},
  {32'h4338e2c4, 32'h430a6a14, 32'h43a3157e},
  {32'hc3cdfe7a, 32'hc38c737d, 32'h43af7755},
  {32'hc2c0514f, 32'h4380b2e3, 32'hc358bbd5},
  {32'hc3ff67f6, 32'h4300b1aa, 32'hc33f7422},
  {32'hc3263036, 32'hc382d854, 32'hc2ec17ea},
  {32'h43d978c6, 32'hc28a85a3, 32'hc3b51985},
  {32'h433e047f, 32'h424cc121, 32'h41d21da0},
  {32'h43353893, 32'hc3f570ba, 32'hc421002c},
  {32'h42b07b76, 32'hc222c230, 32'h43a48fcd},
  {32'hc38a79b0, 32'h4333fb1d, 32'hc3395f44},
  {32'h439d5c01, 32'h41dc2006, 32'hc405db15},
  {32'h43e70670, 32'hc2d7ea76, 32'hc39b82c1},
  {32'hc32ed857, 32'h41be8a66, 32'hc35300ee},
  {32'h4170d11b, 32'h43ae613f, 32'hc3a01bc8},
  {32'h42f6e110, 32'hc2f20663, 32'hc33bb796},
  {32'h41bb0bf8, 32'hc388f23a, 32'h43430a44},
  {32'hc268ee0a, 32'h41dd5751, 32'hc32a2857},
  {32'h44188e17, 32'h42a0d1be, 32'h44442b97},
  {32'hc2e6b573, 32'hc3f9b090, 32'h42f27307},
  {32'hc258621c, 32'h4348b7d9, 32'hc310f5ca},
  {32'hc378ea00, 32'hc04565aa, 32'hc27877fa},
  {32'h4353f5f1, 32'h4284fe48, 32'hc27f4d21},
  {32'hc3065a49, 32'hc3b02560, 32'hc3c4bcad},
  {32'h438af84d, 32'h42ee70c0, 32'h43f94603},
  {32'hc4211a1a, 32'h438d844d, 32'h4359712c},
  {32'hc2f9139e, 32'hc28c191f, 32'h4364871b},
  {32'hc3151806, 32'hc26815c8, 32'h416eaff5},
  {32'hc281d98c, 32'h43985767, 32'h43ac9662},
  {32'h433eb52f, 32'hc3376080, 32'h42638e41},
  {32'h43179b24, 32'h42669506, 32'hc1b8b9d3},
  {32'hc2db7b25, 32'hc301bb5e, 32'h41da944e},
  {32'h4204367c, 32'hc39590cf, 32'h430fcdd1},
  {32'h439f0c75, 32'hc384e0b8, 32'hc31e1cf2},
  {32'hc283dad5, 32'hc2f2e400, 32'h428a9bfd},
  {32'hc4024a44, 32'h4347fa62, 32'h438e4cde},
  {32'hc3402df7, 32'h431b43bf, 32'hc34b5a86},
  {32'h4362df00, 32'h4364b196, 32'h42a7843f},
  {32'hc3fe0781, 32'h436a2062, 32'hc31148d9},
  {32'h44256531, 32'h432b862e, 32'h42deb657},
  {32'hc3d2f6d6, 32'hc22e2767, 32'hc29a0763},
  {32'hc3b86480, 32'h43141814, 32'h42a68c45},
  {32'h4200bd8d, 32'h437a56ba, 32'h42dee27b},
  {32'h411bcb70, 32'h41f6e76d, 32'hc30f3e36},
  {32'hc3567902, 32'hc3bb8176, 32'hc35dc0d5},
  {32'h43d476b2, 32'hc2f07004, 32'h43710f56},
  {32'hc31b597d, 32'h4384a2f2, 32'hc2de3cab},
  {32'h42d167ba, 32'hc3e60264, 32'h3fb4ee98},
  {32'h43af0391, 32'h4397df22, 32'hc2bc20c0},
  {32'h439159c2, 32'hc29c8fe1, 32'h42f032bd},
  {32'hc32cfd65, 32'hc320f3c6, 32'h42d15eed},
  {32'h44041fdc, 32'hc3f8457a, 32'h43bf2cc5},
  {32'hc42f94d7, 32'hc3ead344, 32'hc338566e},
  {32'hc28f4150, 32'h4202ad14, 32'hc0893200},
  {32'hbfd81c78, 32'hc277167c, 32'h429906b9},
  {32'hc3a74147, 32'h439021b8, 32'h42d05d26},
  {32'h437e232c, 32'h43869450, 32'hc37a3926},
  {32'h434bd62f, 32'hc3a1be1c, 32'hc34d7d9b},
  {32'h430d4887, 32'hc3c37e8f, 32'hc3a69a99},
  {32'h429abbf0, 32'h43307bba, 32'h41a2a4ca},
  {32'hc31f37fd, 32'hc2b54a50, 32'h4236511d},
  {32'hc32f41f8, 32'h422a4b04, 32'hc2728b7b},
  {32'hc38ba805, 32'hc354a9ac, 32'h426c7537},
  {32'hc3853161, 32'h438b850f, 32'h4250fad2},
  {32'hc2908000, 32'h421866d3, 32'hc3281f90},
  {32'h430f4fdc, 32'hc2642c37, 32'h430f6fab},
  {32'hc362f096, 32'hc3646915, 32'h42e257cc},
  {32'hc263418a, 32'hc30f7055, 32'hc34604e4},
  {32'hc307f00a, 32'hc3ad68e7, 32'hc3985658},
  {32'hc096d430, 32'h40d25253, 32'h43baf5cc},
  {32'hc2cea978, 32'h434996b0, 32'hc38ae0fd},
  {32'hc3e07a86, 32'hc3c9d8d7, 32'hc3b1dcd9},
  {32'h43e1f857, 32'h414bb666, 32'h440217b8},
  {32'hc2723355, 32'h42a6631a, 32'h42ab4940},
  {32'hc2bdfd7c, 32'h42e7f8e3, 32'h4349d853},
  {32'h42e6fedd, 32'h434ee892, 32'h43197988},
  {32'hc3894c40, 32'hc38dae4c, 32'hc35fc921},
  {32'hc252d980, 32'hc40bfeb3, 32'hc382ab4c},
  {32'hc30eafbf, 32'hc40c5a42, 32'h43906a1a},
  {32'h42fc8ad0, 32'hc386f470, 32'hc3881c1f},
  {32'hc33bb95c, 32'h4259f809, 32'hc0c8de94},
  {32'hc33e85ae, 32'hc3a19f14, 32'hc3a46da8},
  {32'hc3ba226f, 32'hc1f53f96, 32'h42f93088},
  {32'hc1671f10, 32'hc396182d, 32'hc2f754cb},
  {32'h440c1ceb, 32'hc33497d8, 32'hc3c3c1ce},
  {32'h430eb817, 32'h4391332d, 32'hc4597694},
  {32'hc3d3e267, 32'h437bb362, 32'h43f8ad1e},
  {32'h42ce7b41, 32'hc2535715, 32'hc22ef4c4},
  {32'hc3e3e800, 32'hc2b95c81, 32'hc32c33fb},
  {32'hc102e087, 32'hc34c2680, 32'hc33cd308},
  {32'hc398c6d6, 32'hc3a930a4, 32'hc382ad78},
  {32'hc3c36b3e, 32'hc30bd506, 32'h43573caa},
  {32'hc38079d8, 32'hc354ffd0, 32'h4372dc1e},
  {32'h43baa989, 32'hc38d6854, 32'hc11269b5},
  {32'hc390de89, 32'h43198268, 32'hc31dfd1c},
  {32'hc29aa2c8, 32'h42047375, 32'hc2aeebed},
  {32'hc26e5301, 32'hc2fafd5a, 32'h439d7932},
  {32'hc33a0150, 32'hc2e74ff2, 32'h43a03e5c},
  {32'hc2d3abfb, 32'hc3da56fb, 32'hc3c4460e},
  {32'h433e41c4, 32'hc3f9802e, 32'hc360ebc0},
  {32'hc3ac8e56, 32'hbffb0cb2, 32'h4369cb89},
  {32'hc3b18526, 32'hc3dfd350, 32'hc30d251e},
  {32'h4323f7db, 32'h43c7ed4e, 32'hc2068da6},
  {32'hc385b3bc, 32'h43a2eeb7, 32'hc395af2a},
  {32'hc39b4040, 32'h42e59462, 32'hc2d74bd5},
  {32'h4345da6d, 32'hc31182de, 32'h4470b16f},
  {32'hc141aa8c, 32'hc1aa5efc, 32'hc359adbc},
  {32'hc2bda551, 32'h434638fd, 32'h42abea73},
  {32'hc353c0b7, 32'h42e2bb35, 32'hc32e07db},
  {32'h4331160c, 32'h435c8cca, 32'h431d120d},
  {32'hc231fa99, 32'hc289b495, 32'h42dc6ec2},
  {32'h4166268a, 32'h41b1f62f, 32'hc38bdc43},
  {32'hc1a16c4c, 32'h42ad03e5, 32'hc395daf5},
  {32'hc1b6cfb7, 32'h4319bc3b, 32'hc3a24cf6},
  {32'hc206af53, 32'h424005d2, 32'hc3a1d191},
  {32'hc384185a, 32'h40a45bb9, 32'hc332d91e},
  {32'hc310ad65, 32'hc2da3918, 32'hc38893cd},
  {32'h43351dab, 32'hc3aa8de1, 32'h434d0615},
  {32'hc16a68c4, 32'h43961a16, 32'h445d5bb0},
  {32'hc23c5e62, 32'h43a7319c, 32'h4358ee90},
  {32'h43cf3ffd, 32'h4261178a, 32'hc39b3f32},
  {32'h42bf8c9f, 32'h4326d4fa, 32'h42907720},
  {32'hc4051c98, 32'hc3a2eb43, 32'h42985363},
  {32'h4345e150, 32'hc2a3c75a, 32'h439406c0},
  {32'hc30bb228, 32'hc30b95ad, 32'h42ee2a02},
  {32'h41deb050, 32'h429fe4b4, 32'hc2883e20},
  {32'h439e1716, 32'hc281e2bd, 32'h43d059a8},
  {32'hc2c78fa4, 32'h414976e8, 32'hc3c2bebc},
  {32'h438ebc95, 32'h43dae180, 32'hc34006ef},
  {32'h43b080aa, 32'h44087caa, 32'hc3546ee1},
  {32'h43849764, 32'hc291355d, 32'hc28267dd},
  {32'h426bb6b9, 32'hc31c658f, 32'h4379eaba},
  {32'h42343677, 32'hc4011059, 32'h426ed132},
  {32'hc3f397f8, 32'h424da996, 32'hc275381c},
  {32'hc3314028, 32'hc20bcd30, 32'hc30c385d},
  {32'hc321d5a1, 32'hc3dcb9d4, 32'hc334aa91},
  {32'hc4013fa1, 32'h434ca8c7, 32'h4422e1d2},
  {32'hc382aa9a, 32'hc2b84f53, 32'h438c2fd4},
  {32'h42a54ea9, 32'h42ce9cf4, 32'hc31ccbd1},
  {32'h41d777a0, 32'hc378b959, 32'hc2d0a8a9},
  {32'hc2d1d135, 32'hc39200e6, 32'hc3de0f26},
  {32'h44098c93, 32'hc1baf0a8, 32'hc34286e9},
  {32'hc3a4a061, 32'hc39303f5, 32'hbfefc668},
  {32'hc225514f, 32'hc35cbb9a, 32'h4371f124},
  {32'hc3ad8a56, 32'h41d43c4d, 32'h43851806},
  {32'hc3ad68d6, 32'h439729bc, 32'hc36d1c73},
  {32'hc3eda32d, 32'h415c9b5c, 32'h43d785cf},
  {32'h442733bb, 32'h436bfcab, 32'hc3977879},
  {32'hc266d901, 32'hc39d2664, 32'hc2b9e10b},
  {32'hc23fe8c7, 32'hc38d7eb1, 32'hc25064b5},
  {32'h43fcd906, 32'hc1a8df5c, 32'h42c78777},
  {32'hc1fc488a, 32'hc3500150, 32'h434be931},
  {32'h41837030, 32'h43cba27c, 32'hc39f01ff},
  {32'h43a8896a, 32'hc39bc963, 32'h4379b886},
  {32'hc3de94c5, 32'h43cfafdc, 32'hc3cf41f7},
  {32'h42f83a03, 32'h440504db, 32'hc34868a8},
  {32'h43884681, 32'h4431d94c, 32'hc33d6020},
  {32'hc36aa19c, 32'h440b8e51, 32'hc2e7a987},
  {32'h419c0fa1, 32'hc3c0a818, 32'hc2354640},
  {32'h432106c0, 32'hc3f194ec, 32'h4428f0f0},
  {32'hc38740c8, 32'hc34396d7, 32'hc2c17b0c},
  {32'hc2784d1a, 32'hc1d8fd8e, 32'h443dee3d},
  {32'h43b4fc51, 32'hc3006d15, 32'hc22753e3},
  {32'hc31d5fdd, 32'h439dea27, 32'h4396b691},
  {32'h433ccfb9, 32'h4155fcd4, 32'hc35e5c22},
  {32'h438087b0, 32'hc337568d, 32'h431ea744},
  {32'hc42e496c, 32'h42b3316c, 32'h43199f79},
  {32'hc1bd1e0a, 32'h42b211a7, 32'h4380a591},
  {32'h40b91dc8, 32'hc2aaa194, 32'hc34b473b},
  {32'h4309bdc8, 32'hc40c3d2e, 32'hc302bd03},
  {32'hc3bd7ab5, 32'hc385409c, 32'hc3801104},
  {32'h42a4986c, 32'h438511eb, 32'h43de1349},
  {32'hc339e4a8, 32'h436b376f, 32'hc091fc0f},
  {32'h43b19654, 32'h42b3e87b, 32'h437c70be},
  {32'hc3d80df4, 32'hc3826f03, 32'h436084ff},
  {32'h4313f8a2, 32'hc29d296f, 32'hc3af4117},
  {32'hc2e29c2e, 32'h4306debc, 32'hc376fda4},
  {32'h4420a2c3, 32'h43940868, 32'h442174ad},
  {32'hc2f52cb7, 32'h4435abe6, 32'h43c2740d},
  {32'hc21368c2, 32'h43bc953a, 32'h43e5e086},
  {32'h43857f90, 32'h439ee984, 32'h4310d160},
  {32'hc40ae8e1, 32'h438598be, 32'hc3f42326},
  {32'h428c0c28, 32'hc35c349d, 32'hc30161e4},
  {32'h419d1e1f, 32'hc3cfd217, 32'h443621f1},
  {32'hc2c63eea, 32'h42cbaf1e, 32'hc3a22c9b},
  {32'hc1ac9bf2, 32'hc341c3f0, 32'hc34be440},
  {32'hc32e9730, 32'h429da129, 32'h3f32b230},
  {32'hc390d41a, 32'h42dfd6e5, 32'hc3801ba4},
  {32'h42d5241d, 32'hc200c30c, 32'h441b1c6f},
  {32'h43088ffa, 32'h432d420b, 32'hc32f6535},
  {32'hc41bf47c, 32'h43834855, 32'h4402225e},
  {32'hc354e2a4, 32'hc24ffeb9, 32'h4362b201},
  {32'hc339eb37, 32'h40fd0e95, 32'hc2ca2b58},
  {32'hc3ba0d80, 32'h44080741, 32'hc197b11f},
  {32'hc38d960a, 32'hc2ac870d, 32'hc3b46a8c},
  {32'h43fc4323, 32'h42b09b65, 32'hc30d8f19},
  {32'hc38c3a19, 32'hc403bfa7, 32'hc3ab7ad6},
  {32'hc2f5fa25, 32'hc30c65d7, 32'hc38223dc},
  {32'hc3aa2547, 32'h44506a89, 32'h433a97c8},
  {32'hc3d43107, 32'h43b06664, 32'hc345993d},
  {32'hc40ce183, 32'h4383f9da, 32'hc406cc63},
  {32'h441806a5, 32'h42bd5e1c, 32'hc1b4a061},
  {32'h414f264e, 32'h4212c641, 32'h41d966ea},
  {32'hc3879d6a, 32'hc34cbd34, 32'hc3966628},
  {32'h43328080, 32'hc346cf2e, 32'hc1b97588},
  {32'hc41f0117, 32'hc14fbb80, 32'h43db5ecf},
  {32'h41b8d7a2, 32'h432f6110, 32'hc3a88c22},
  {32'h43dde683, 32'h43a5cc88, 32'hc32e8192},
  {32'h4434976f, 32'h42850053, 32'hc30546f8},
  {32'h435fd9c3, 32'h431db3a4, 32'hc253060c},
  {32'h439a0864, 32'h42aa0668, 32'h4380935f},
  {32'hc2a27739, 32'hc3c8e7a7, 32'h432978b9},
  {32'hc34bf976, 32'h42ec8208, 32'h43ed2c36},
  {32'h428a8889, 32'hc311f2e3, 32'h436924e9},
  {32'h42a0d62c, 32'hc38ee94c, 32'hc3a4d988},
  {32'h4178e2b2, 32'h431a4900, 32'h4328e1c4},
  {32'h43b1e391, 32'hc38a3253, 32'hc33e2c78},
  {32'hc3899a3e, 32'h434effc8, 32'h434a2351},
  {32'hc361e57f, 32'h438e5731, 32'hc13db17c},
  {32'hc33f615e, 32'h441457e2, 32'h4442065d},
  {32'hc3815d08, 32'hc3797714, 32'h4398d01a},
  {32'hc30c9044, 32'hc3a891a5, 32'hc3a9bb87},
  {32'h42ca7ffc, 32'hc23071b9, 32'hc3fed361},
  {32'hc4122b09, 32'hc39ad10c, 32'hc2a50b1c},
  {32'h4301a039, 32'hc23005f3, 32'hc3774259},
  {32'h43913daf, 32'hc2b9a80d, 32'h4364b77c},
  {32'h430edd3c, 32'hc2fc1787, 32'hc19c465a},
  {32'hc3d52963, 32'h4409eda6, 32'hc37cbb10},
  {32'hc3111b4a, 32'hc3818d5b, 32'h42063248},
  {32'h4323ac0d, 32'h43ecc41e, 32'h432e377a},
  {32'h41dcf9e3, 32'h40ba99ac, 32'h41af0434},
  {32'hc2c23010, 32'h4328b70b, 32'h42ce48c4},
  {32'h43101545, 32'h4318f53b, 32'hc3a06364},
  {32'h434157bc, 32'hc3b43c64, 32'h433de4dc},
  {32'h442d3ae5, 32'h4385623a, 32'h442a88de},
  {32'hc31de286, 32'h429b7a0b, 32'h4304935b},
  {32'hc2ef5fb5, 32'h439a64ed, 32'hc41434d2},
  {32'h42a5ff18, 32'h43c98601, 32'hc309206a},
  {32'h438727ad, 32'hc31737ef, 32'hc330c049},
  {32'hc2292074, 32'hc290679d, 32'h4282421c},
  {32'h43a77f00, 32'h43a56508, 32'hc279c4a1},
  {32'hc3fa81b5, 32'h43266840, 32'h4305e10e},
  {32'hc2ef3316, 32'h42b0b69d, 32'hc289c8c6},
  {32'hc3207032, 32'h432d662a, 32'hc41f82e4},
  {32'hc42235c7, 32'h43bba394, 32'h43bdeb4e},
  {32'h429e2ae4, 32'hc365f2a0, 32'hc2792c2a},
  {32'hc30869ee, 32'h42f3e9cf, 32'hc330ed5a},
  {32'hc3228ebb, 32'hc3ecc5a9, 32'h437c494b},
  {32'h426e4f8a, 32'h43683a22, 32'hc078ae30},
  {32'h42af61eb, 32'h420c881d, 32'hc3269a38},
  {32'hc2d040ae, 32'hc2709a2b, 32'h4301d4df},
  {32'hc36ee3a8, 32'h43aa6597, 32'h4396f939},
  {32'hc31de452, 32'h429e4643, 32'h42cfc943},
  {32'h43535bcb, 32'h4090768d, 32'hc3bdf0a4},
  {32'hc4021cf8, 32'h43b0a9ed, 32'h431c2756},
  {32'h44298ca0, 32'h41e25ae6, 32'hc2c8aa99},
  {32'hc3247c47, 32'hc40606a2, 32'hc3128013},
  {32'hc37d98e6, 32'hc33a0659, 32'h43dd6e26},
  {32'h4408d4b9, 32'hc26edb99, 32'hc4137cc2},
  {32'h43351518, 32'hc3e54381, 32'h4372f276},
  {32'hc3878736, 32'hc3dbbc8d, 32'hc24e53b4},
  {32'h429f64b2, 32'hc293ef81, 32'hc23c199d},
  {32'h430e9234, 32'h411ed25a, 32'h429ce3c1},
  {32'h433cd6ec, 32'h41e9086c, 32'h431424c8},
  {32'h42b89fec, 32'h435261ad, 32'h436be210},
  {32'hc3997446, 32'hc305f4d1, 32'hc2dd86e4},
  {32'h43b0565d, 32'h4295fb8b, 32'h4337b182},
  {32'hc301060e, 32'h43f20983, 32'hc385d62e},
  {32'h438f8aa1, 32'hc26d9400, 32'hc373bfc0},
  {32'h428de987, 32'h430e6cd2, 32'h41a89655},
  {32'h4356fc08, 32'h43925f4c, 32'hc397dcf8},
  {32'h41bd6d12, 32'hc30c0b86, 32'h440f6cba},
  {32'h426acc99, 32'hc3453380, 32'h43a58437},
  {32'h42bf78a1, 32'hc36484c2, 32'hc368a43b},
  {32'hc1c71868, 32'hc365adfe, 32'hc21d3efc},
  {32'hc1ad71b6, 32'h40c9bdcc, 32'hc3f596af},
  {32'h43a806d8, 32'h42e0cbef, 32'hc3fd5853},
  {32'hc1fed98f, 32'hc30790cf, 32'h41ecddb8},
  {32'hc3e9cb1f, 32'h4316224c, 32'h42ab1589},
  {32'hc3c99aa0, 32'h4170c164, 32'h43a375da},
  {32'hc2eb6332, 32'hc33c6ba6, 32'h4364b0b3},
  {32'h41ed2860, 32'h439308ee, 32'h43006610},
  {32'hc2314043, 32'hc386943d, 32'h419f2dec},
  {32'hc2f63865, 32'hc30f7df6, 32'hc2fc767d},
  {32'hc2d68e5c, 32'h41eddb48, 32'hc1df98be},
  {32'h43d09fbf, 32'hc31b6da1, 32'hc27d00c6},
  {32'h425292e4, 32'hc288bed8, 32'h426bf2fa},
  {32'hc2d65dd2, 32'h4313e1c0, 32'h43ee42c2},
  {32'h43cd1018, 32'hc39a109f, 32'h4390fe51},
  {32'hc3969982, 32'h4300fccf, 32'hc2ba08c0},
  {32'hc2106ecc, 32'hc3003ff8, 32'hc3a236b4},
  {32'h43958b87, 32'h43ed490a, 32'hc3f7181f},
  {32'h431a193e, 32'h43765dd6, 32'hc3bd89ce},
  {32'h42a7b56c, 32'hc236dbd5, 32'h423f1480},
  {32'hc341fc3a, 32'h42e2471d, 32'hc26d17d1},
  {32'hc3dd2e08, 32'h43f3da19, 32'hc28097ae},
  {32'hc21e53de, 32'h437de4e3, 32'h4401dc20},
  {32'h43189458, 32'hc3a1b986, 32'hc4277d75},
  {32'h42918f94, 32'h43b479b7, 32'hc336fd6d},
  {32'hc2b46862, 32'h420f712b, 32'h43506f05},
  {32'h4353e479, 32'h4413f454, 32'hc3db2c68},
  {32'hc39e61d4, 32'h439250c6, 32'hc2769d87},
  {32'h43873c0e, 32'h43bab1f1, 32'hc405525f},
  {32'h42e21fd1, 32'h41911430, 32'hc31fe164},
  {32'hc431e488, 32'hc217ddc9, 32'hc2526800},
  {32'h43bc7453, 32'hc35f0d2c, 32'h4212b52d},
  {32'hc39242e6, 32'hc362956c, 32'hc3b55a73},
  {32'hc2cd3ec1, 32'h3f3437ac, 32'h40fe90c4},
  {32'hc2f79c07, 32'h43653ff4, 32'hc2823d23},
  {32'hc34b3a52, 32'hc3d480ea, 32'h43ed80bb},
  {32'hc2e57d48, 32'h43223ce3, 32'h42fc35f1},
  {32'hc40b9afa, 32'hc378ceb1, 32'h42875119},
  {32'h42b84295, 32'h430cd714, 32'h42081b9c},
  {32'hc3b64552, 32'hc2e74649, 32'h4348b8e0},
  {32'hc3d8a307, 32'hc2b5d277, 32'hc3869d9f},
  {32'hc101d100, 32'hc30ebba5, 32'hc2fbbe4e},
  {32'hc4074308, 32'h4335dba4, 32'h4017954e},
  {32'hc3c017cf, 32'h43225324, 32'h43ea3381},
  {32'hc37c853b, 32'h43c3f51b, 32'h3f60b0c4},
  {32'hc36e6235, 32'h43d9bd13, 32'hc3aa1115},
  {32'hc2c194d8, 32'hc22c98a5, 32'hc1f25547},
  {32'h42261bf4, 32'hc3980349, 32'hc2e1ed20},
  {32'hc3905ccb, 32'h436388fd, 32'h4309b9e8},
  {32'hc3b9edfc, 32'h436b181c, 32'h43c71c35},
  {32'hc3a109fb, 32'h4337e25c, 32'h421a5eb4},
  {32'hc1234416, 32'h4336dfd0, 32'h4305dd9f},
  {32'hc3042a9f, 32'hc3a2d5a5, 32'h42071008},
  {32'h4299ecb4, 32'h4204037a, 32'hc3d7f26f},
  {32'hc2073aa6, 32'hc3883b72, 32'h439549b7},
  {32'hc2a1647e, 32'h43c3e124, 32'hc2885604},
  {32'h41761d62, 32'hc34690f4, 32'hc3ddfb30},
  {32'hc2159172, 32'hc226a006, 32'hc254b297},
  {32'hc3861192, 32'hc217af4d, 32'hc2a73e60},
  {32'h4292029d, 32'hc3386662, 32'hc31bec40},
  {32'h44111f3a, 32'hc329787b, 32'hc3136cf2},
  {32'h4421c49f, 32'hc28d79e3, 32'h4354eff6},
  {32'h426757e8, 32'h43e4256f, 32'hc4385773},
  {32'hc28fbbca, 32'hc2553ecf, 32'h43011d2f},
  {32'hc2e9e614, 32'h429b19af, 32'hc3a8581e},
  {32'h44394e90, 32'hc30c33a7, 32'hc286b6a4},
  {32'hc3fee4c3, 32'h438d4e02, 32'hc217eeb8},
  {32'hc3443cfe, 32'h41eeb518, 32'hc31d644f},
  {32'h43806d5c, 32'hc2fd9552, 32'h42eba0eb},
  {32'hc3bbe254, 32'hc407d864, 32'hc2937572},
  {32'h4380cccb, 32'hc0962fb0, 32'hc38968cd},
  {32'hc2cac090, 32'h43fd622f, 32'h4324eab7},
  {32'hc2928fbc, 32'hc3dd8de7, 32'h42cbe2e4},
  {32'h429afc84, 32'hc1d4a136, 32'hc3923743},
  {32'hc2f98283, 32'hc2399f45, 32'hc2064743},
  {32'hc399c48e, 32'h42717b0a, 32'h43ef4777},
  {32'hc338e143, 32'hc2df1672, 32'hc14cc97f},
  {32'h432963b1, 32'hc282736c, 32'hc3feea08},
  {32'hc39d8feb, 32'h4282fffe, 32'h431974f7},
  {32'h43315b62, 32'hc3a9602a, 32'hc325a478},
  {32'hc364f738, 32'h42d7aa29, 32'hc1e1d461},
  {32'hc383c1e8, 32'h41d8b785, 32'h41928a60},
  {32'hc3852c72, 32'hc365db8c, 32'h403b615a},
  {32'h4309844e, 32'hc3b815d0, 32'hc40b527f},
  {32'h3f97dac0, 32'hc3259c3e, 32'hc3fc411a},
  {32'hc32ac253, 32'h437dfec6, 32'h43d842a1},
  {32'h4366ddd2, 32'hc23f58cc, 32'h43a2f3ea},
  {32'hc3fd3f24, 32'h437eec8d, 32'hc2faa055},
  {32'h43c484ea, 32'h42cc70af, 32'h4389cabf},
  {32'h41df810c, 32'h43633391, 32'h4373d58e},
  {32'hc3d0a7a3, 32'h42dbb695, 32'hc3f625da},
  {32'h413506ce, 32'h429bd029, 32'h4344ef9a},
  {32'h43d17bb2, 32'h42afd158, 32'h43d5bebb},
  {32'hc39e8c28, 32'hc375c964, 32'h427172d5},
  {32'h4253bd04, 32'hc3321533, 32'hc159f1d2},
  {32'h430bf325, 32'hc38b352b, 32'h4393a72b},
  {32'hc30f8c6b, 32'h43995107, 32'hc3a885ec},
  {32'hc425a6ee, 32'hc28c6dfc, 32'hc3f6a657},
  {32'h42f6d50f, 32'hc2d7f9c3, 32'h43d14fe7},
  {32'h4393bd63, 32'h4138131a, 32'h42a89415},
  {32'hc36c4bd1, 32'h42ed6c64, 32'h43f31ccf},
  {32'h43283ec3, 32'h42e83711, 32'h43507c5a},
  {32'h43eaf12d, 32'h42bccf21, 32'h43ed66fe},
  {32'hc34af720, 32'hc3a08c4b, 32'h42e1c993},
  {32'h42de2fff, 32'h430e1fc0, 32'hc3852052},
  {32'hc22ac45a, 32'h433d39b1, 32'h439f7cc6},
  {32'hc3be3fbb, 32'hc2df2e01, 32'hc31e145d},
  {32'h42f653c7, 32'h432cb318, 32'h433107af},
  {32'h42a06c08, 32'h435959bd, 32'hc2abb0ff},
  {32'h4360ff2a, 32'hc3f5e765, 32'h4386a4d0},
  {32'hc3149ae7, 32'hc3f6ac9f, 32'hc160eda7},
  {32'hc3d60c17, 32'h4350c485, 32'hc2887681},
  {32'h42e1eaea, 32'h42e909b6, 32'hc41982c9},
  {32'hc30d2327, 32'h43ee28e7, 32'h4318adc7},
  {32'h426acdcb, 32'h433d198d, 32'h43f254ce},
  {32'hc380c609, 32'h436cb62a, 32'h430250f9},
  {32'h43d188c8, 32'h4201744e, 32'h42e2e359},
  {32'hc3de363a, 32'hbf1aff10, 32'h43eb7aa8},
  {32'hc3318556, 32'h4267149d, 32'hc1c7431e},
  {32'h4392f53d, 32'h432fb10d, 32'hc3e4e0ce},
  {32'hc3648617, 32'h43999efd, 32'hc203c173},
  {32'hc37d67f9, 32'h4330b2c2, 32'hc38f01e9},
  {32'h436de746, 32'h433d9a24, 32'h4370495b},
  {32'hc3177774, 32'h43da3003, 32'hc3fcf6ae},
  {32'hc3688ed4, 32'h42a24599, 32'hc1954ec9},
  {32'hc3215422, 32'h43ac5366, 32'h431cb823},
  {32'hc38fcee3, 32'h42df60fa, 32'h43aae5f8},
  {32'h43be2916, 32'hc36fdf80, 32'hc2f1b283},
  {32'h42aaf42f, 32'hc3a7b3af, 32'h439685bc},
  {32'h43797295, 32'hc4082838, 32'hc39ce0f6},
  {32'h41259c8e, 32'h43e74313, 32'h434eec1d},
  {32'h4378c7b7, 32'hc2229b3a, 32'hc3e16d15},
  {32'hc18c3686, 32'hc31c411c, 32'h430e9b0b},
  {32'hc22e401a, 32'hc1c89a90, 32'h43de6c1f},
  {32'hc389036e, 32'h4390932f, 32'h4260e9c8},
  {32'hc3484ce2, 32'hc2b832b8, 32'h43c456a2},
  {32'hc213964e, 32'hc3d95f47, 32'h40d04d48},
  {32'h433d2fa6, 32'h41bbfcde, 32'hc2b241ea},
  {32'h42d51f22, 32'hc0fdecca, 32'h42625df1},
  {32'h41ae7c5b, 32'h42f3c436, 32'hc3248237},
  {32'h433bf6b7, 32'h42e51128, 32'h436164c3},
  {32'hc4013fd4, 32'hc308a31a, 32'h43101cb5},
  {32'h43a2e029, 32'h438e9fc8, 32'hc337ea95},
  {32'hc226d72a, 32'h417c511c, 32'h42e8caa0},
  {32'hc3ce19a7, 32'h43260258, 32'hc4242bf0},
  {32'h43f1dd74, 32'h434c5958, 32'h427add0d},
  {32'h43b0030f, 32'hc2880d23, 32'h4351799e},
  {32'hc420ab3e, 32'h42cf8be6, 32'h4398a029},
  {32'hc40e45c1, 32'hc39ea763, 32'hc316a52e},
  {32'h43f2c323, 32'hc3ea0916, 32'h43910f96},
  {32'hc37e8df2, 32'h42a1070b, 32'hc2172086},
  {32'hc2822e6e, 32'h42ae2d3f, 32'hc2ec8640},
  {32'h42ca9bbc, 32'h43657812, 32'h4389494b},
  {32'hc310c534, 32'hc334730b, 32'hc2232727},
  {32'h428a19e8, 32'h43007486, 32'hc387b7a0},
  {32'hc1f2e7cc, 32'hc3738bd9, 32'h441a967b},
  {32'hc306f48d, 32'h413dd1ea, 32'h41e4d0fa},
  {32'hc36e44af, 32'h438fd8ba, 32'hc1d0658f},
  {32'h42a5b586, 32'hc331eb0a, 32'hc2d456dc},
  {32'h43b9d39c, 32'h43a84266, 32'hc379879b},
  {32'h43682f72, 32'hc1a86901, 32'hc2de3a30},
  {32'h437234c8, 32'h40e785f0, 32'hc31f0689},
  {32'hc2530cc0, 32'h43335867, 32'hc34c82df},
  {32'hc3cc3982, 32'hc36494c8, 32'h431595e2},
  {32'h438cdef6, 32'h4364a446, 32'h42bbc431},
  {32'hc37d6b5e, 32'h427dc3cf, 32'h4264ddde},
  {32'hc2a79816, 32'hc323ab3f, 32'hc1c6d37b},
  {32'h43192391, 32'hc31cebd1, 32'h41953002},
  {32'hc3764fe9, 32'h437d53fa, 32'hc3944a94},
  {32'hc3dbc848, 32'hc3c5eace, 32'h438b8f49},
  {32'h43add612, 32'h440d0579, 32'hc3fe0b45},
  {32'h4301ccfa, 32'h43a5b254, 32'h40cc281d},
  {32'hc39d2b35, 32'hc3252a45, 32'h437ce096},
  {32'h4314d3f2, 32'h442365db, 32'h433c4ccc},
  {32'hc4149232, 32'h40db12c8, 32'h3fdd524a},
  {32'hc18d5af4, 32'h4304f923, 32'hc2c84d6a},
  {32'h440181be, 32'h42a3181d, 32'hc320d922},
  {32'h4118c110, 32'h436ea721, 32'hc3cbdd9e},
  {32'hc3419c9b, 32'hc2920c3b, 32'h438ca2f0},
  {32'h43649b70, 32'h41a6e206, 32'h42aeed50},
  {32'hc2a1c4d5, 32'hc29c2034, 32'hc3812c26},
  {32'hc3051861, 32'hc3a4218f, 32'hc393407a},
  {32'h43938d30, 32'hc32bbae0, 32'h44474064},
  {32'hc33eb4aa, 32'hc314ab57, 32'h42cbda6b},
  {32'hc022f3d0, 32'hc1d65a61, 32'hc2a291f5},
  {32'hc21717a0, 32'h424cb860, 32'hc1645fbe},
  {32'h42944cce, 32'hc3ec70c9, 32'h4316ccef},
  {32'hc33077ce, 32'hc28b488f, 32'h42b1f9bd},
  {32'h43eeb776, 32'h43153106, 32'hc39ad287},
  {32'hc284016e, 32'h43a37f38, 32'hc40b5f23},
  {32'hc3046b6b, 32'hc2c2daed, 32'hc3087d15},
  {32'h43cbab81, 32'h43bb4a8e, 32'h42dff620},
  {32'hc3ae1062, 32'h411bd4f8, 32'h4308e4f5},
  {32'hc3a2e539, 32'h435b676c, 32'hc2d7ee6b},
  {32'h438c51b0, 32'h433d988c, 32'hc3fa1cb7},
  {32'hc2f6b71b, 32'h43b4d2e8, 32'h44356b49},
  {32'hc3d5b7a1, 32'hc3e80d0c, 32'h431e8b0a},
  {32'hc324809a, 32'h418cea89, 32'h42a549b3},
  {32'hc395bfd1, 32'hc3ee1ead, 32'hc2a65c0e},
  {32'h43b350b7, 32'hc3ec11a3, 32'hc2de5241},
  {32'h44290e79, 32'h4381c94a, 32'hc3318ce9},
  {32'hc35362bd, 32'hc3cb28ec, 32'hc2a5753a},
  {32'h43114d9c, 32'hc41052f3, 32'hc2980720},
  {32'h43731bab, 32'hc3c21c4d, 32'h43a3595e},
  {32'hc3c3fd3f, 32'hc3c12e50, 32'hc3a16bb7},
  {32'hc3d7cdf6, 32'hc3128d11, 32'hc39dc509},
  {32'hc23ef09e, 32'h42afe5eb, 32'hc349b17c},
  {32'hc2efc12b, 32'hc337f567, 32'h43370959},
  {32'hc39e2edf, 32'h436847ee, 32'hc2e75f9c},
  {32'h42b121c2, 32'hc2c27d8d, 32'h424880c0},
  {32'hc3dda443, 32'h434f796c, 32'hc3275484},
  {32'hc3059878, 32'hc3389b65, 32'h428d063f},
  {32'h43394136, 32'hc34ed6a8, 32'h41ceb8c4},
  {32'hc378579c, 32'h433c76e5, 32'hc2d5935a},
  {32'hc1af5504, 32'h4397e92e, 32'h4267f4c8},
  {32'h43083eb3, 32'hc29e7197, 32'hc3453273},
  {32'hc3a742f0, 32'hc3977236, 32'hc3837bec},
  {32'h43d379dd, 32'h4418c1ac, 32'hc3af6cf3},
  {32'hc31423f8, 32'hc2bad817, 32'hc3dd5dbb},
  {32'hc27ddda7, 32'h433fc67d, 32'hc4033206},
  {32'hc3183ac5, 32'hc3719afd, 32'hc36b3d73},
  {32'hc315c89a, 32'h43868e7f, 32'h4398c2f1},
  {32'h421d4bcd, 32'hc1a2ef91, 32'h4397b137},
  {32'hc330abdf, 32'h42504b3e, 32'h44101d19},
  {32'hc1cf22f1, 32'h41ef52ad, 32'h4424744a},
  {32'h41f905a8, 32'h4385a428, 32'hc3806990},
  {32'hc37763f0, 32'hc3484e0c, 32'hc1117d76},
  {32'h42ac5fbf, 32'h43145d26, 32'h435ec22f},
  {32'h430fcabf, 32'hc3647ebc, 32'h40c3ae84},
  {32'hc2257270, 32'hc3fc9972, 32'hc3aa459d},
  {32'h43dace17, 32'hc168ef9a, 32'h43eb262a},
  {32'h42630282, 32'hc34aad7f, 32'h43792789},
  {32'hc2134320, 32'hc2a9ce0f, 32'hc2ad04c0},
  {32'h435a98f4, 32'h438155ee, 32'hc28704d5},
  {32'h43e14dca, 32'hc2df158d, 32'h43d6a73a},
  {32'hc219c098, 32'hc37e305a, 32'h43a3e278},
  {32'h43a30396, 32'hc21e810d, 32'h430edacb},
  {32'h43931853, 32'hc28611ef, 32'hc3db2951},
  {32'h42facd51, 32'h433087c4, 32'h4329cf27},
  {32'h43e0e740, 32'h43d39b0c, 32'h43767791},
  {32'hc302cd09, 32'hc29cfd17, 32'hc25397a9},
  {32'hc350b17f, 32'hc36c8f24, 32'hc398184c},
  {32'hc409d08b, 32'h41d417d9, 32'hc2893d45},
  {32'hc3bfa42c, 32'h43afa98d, 32'hc24c3340},
  {32'h4307f300, 32'h4329c41d, 32'hc3f4b108},
  {32'h439223cf, 32'hc276aaec, 32'hc25912db},
  {32'hc340fa99, 32'hc2f41fd6, 32'hc3eb4f0d},
  {32'hc32f0206, 32'h429097b2, 32'h42e71cba},
  {32'h412d2438, 32'hc3ccf512, 32'hc2613406},
  {32'hc41193fe, 32'hc42653cd, 32'hc35bc6f3},
  {32'h4303cabd, 32'h41e0f7ce, 32'h432e35fe},
  {32'h43eb63f5, 32'h429c558e, 32'h42eb9d3b},
  {32'h40da4c65, 32'hc23ce59c, 32'hc2c3e3de},
  {32'hc3bf7893, 32'hc38876b4, 32'hc39f35a6},
  {32'h4335b162, 32'h41d603d6, 32'hc2da891f},
  {32'h4264954b, 32'hc3ab9f81, 32'hc332bfea},
  {32'h42af7d66, 32'h414648de, 32'h4319dcc0},
  {32'h441bc2dc, 32'hc2dcfc53, 32'h444d9b5d},
  {32'hc36b86c5, 32'hc3a0145b, 32'h43f8c8eb},
  {32'hc37c1bb1, 32'h4316ed85, 32'hc397f531},
  {32'h43325f3e, 32'hc3e30f6e, 32'h43bdd114},
  {32'hc29b742d, 32'h421bf80a, 32'hc1090c1a},
  {32'h41b592dd, 32'hc3062041, 32'h43e40e5d},
  {32'h4304591b, 32'hc3cc91a7, 32'hc143edab},
  {32'hc3d4d645, 32'hc3a9f497, 32'hc35d7214},
  {32'h42d79fe7, 32'h43878a8f, 32'h43921fc5},
  {32'hc33edc11, 32'hc35e2d2b, 32'h411f6801},
  {32'hc3b6dc02, 32'h439c5c43, 32'h43b2e6ca},
  {32'h42eae381, 32'hc3a84891, 32'h438e33c2},
  {32'h413af2d2, 32'hc334a962, 32'hc30cd302},
  {32'hc3108db6, 32'h4390bd2e, 32'h43f21357},
  {32'hc308f1ae, 32'hc39b8352, 32'hc3f040b4},
  {32'hc300b9d9, 32'h42c20e3a, 32'h43a9d43e},
  {32'hc3ff94d0, 32'hc30170d4, 32'h40d2b6fc},
  {32'hc41a94dd, 32'h4357e7b6, 32'h438c8d47},
  {32'hc3d2bdd3, 32'h43e3bcf7, 32'hc3141d87},
  {32'hc3fe033f, 32'h4342418b, 32'hc31356ab},
  {32'hc3f55c4e, 32'h43e760ae, 32'h4300cf83},
  {32'h4340f50e, 32'h413e7414, 32'h42fbb544},
  {32'h4337fecb, 32'h41c50a65, 32'hc361ecaf},
  {32'hc304f1cd, 32'h43393b7e, 32'h42072eab},
  {32'h43789e26, 32'hc3b3b1aa, 32'hc402403a},
  {32'h42d8cea3, 32'hc3896962, 32'hc356743a},
  {32'hc1c12ac0, 32'hc1c7f48e, 32'hc312c38f},
  {32'hc1b72228, 32'hc33c8e90, 32'hc1ab5260},
  {32'h41a806b6, 32'hc385a59f, 32'hc1781d29},
  {32'hc3937566, 32'hc2881818, 32'hc3d82ae6},
  {32'hc2a7a54e, 32'h43480971, 32'h42840442},
  {32'h43df1cde, 32'hc34e67ee, 32'h43852f7c},
  {32'hc2a4d2d7, 32'h439963d4, 32'h43a4dfc8},
  {32'h43a16b79, 32'hc3327be2, 32'h440e4b3e},
  {32'hc2fa7722, 32'h43756e9d, 32'h43c1e2f0},
  {32'h42ba17bb, 32'h4125033a, 32'h41e5c106},
  {32'h4226e8b1, 32'hc312f146, 32'hc3feaadf},
  {32'hc407a644, 32'h438e0129, 32'h43f88bb8},
  {32'hc34cc503, 32'h42a45c20, 32'hc4120bae},
  {32'hc1ca05e8, 32'hc34328fa, 32'hc3694909},
  {32'hc416353e, 32'h43c909b4, 32'hc193853d},
  {32'h42564515, 32'h4343b68f, 32'hc40cf4e2},
  {32'h434eeed2, 32'h435211d9, 32'hc353a106},
  {32'hc343c710, 32'hc3529a7c, 32'h4385f1ed},
  {32'hc2a0b967, 32'h430cfd94, 32'h438949fe},
  {32'h40c255c0, 32'hc2b2d296, 32'h43adb02a},
  {32'hc387f6de, 32'h43469fa4, 32'h41a8d6bd},
  {32'hc391eb14, 32'h430e9b78, 32'hc2ce95b3},
  {32'hc3e59c36, 32'h43117049, 32'h43cce0c6},
  {32'hc402006b, 32'hc2a63534, 32'hc2003f9e},
  {32'hc4177891, 32'hc259a4d4, 32'hc317149d},
  {32'h442ccd9f, 32'hc2960967, 32'hc391414d},
  {32'h419bd48c, 32'hc32651bf, 32'h436ef639},
  {32'hc3b88214, 32'hc33865ed, 32'hc30daa18},
  {32'h435575c4, 32'hc384aa34, 32'hc24aecc5},
  {32'hc389e425, 32'h4303c3b9, 32'hc2597381},
  {32'hc2d9a87c, 32'hc2265a83, 32'hc3e10071},
  {32'h43a9471f, 32'hc3334bbe, 32'hc2dc23c3},
  {32'h420813ac, 32'h4336c1a1, 32'h422eff42},
  {32'h43782109, 32'hc389a195, 32'h43a7143e},
  {32'h43328194, 32'h4337a4e4, 32'hc284e0c8},
  {32'hc19f2502, 32'hc334de1e, 32'hc2871293},
  {32'hc2f523e1, 32'hc19e899b, 32'h435ed0fa},
  {32'h433a7caf, 32'hc33b291c, 32'hc2d3301e},
  {32'hc4338617, 32'h439652c7, 32'h44033e5a},
  {32'h420353a3, 32'hc2f032a9, 32'h427f4c30},
  {32'h436442a2, 32'h42b5aba3, 32'h4302bdfe},
  {32'hc1ee712b, 32'hc3f90c1f, 32'h42bef176},
  {32'h43830d34, 32'h43a8457c, 32'hc318519b},
  {32'h4380bd18, 32'hc3bd7812, 32'hc1c64eee},
  {32'hc34a9a75, 32'h4184ba2b, 32'h4267ce7c},
  {32'hc34db6b0, 32'hc19601a6, 32'h436ddf3f},
  {32'hc2b75985, 32'hc2e69839, 32'h41430960},
  {32'h4326cd84, 32'h437802d0, 32'h43ce6d3a},
  {32'hc3513ffd, 32'h42bcb8bf, 32'h42d6e60c},
  {32'hc3bde00d, 32'h4335246e, 32'h43d39330},
  {32'hc3681f74, 32'h43c4bb17, 32'hc34fc028},
  {32'h41b5fb2f, 32'hc38ac975, 32'hc3839254},
  {32'hc28b404d, 32'hc3cf4623, 32'hc2038d83},
  {32'hc305640c, 32'hc3ceea5d, 32'hc162630a},
  {32'hc35f89f1, 32'h434735f3, 32'hc3d0acfb},
  {32'h4339c559, 32'h438de68a, 32'h436e4131},
  {32'hc117a72e, 32'hc29d0a81, 32'h43555fc3},
  {32'h438c236b, 32'h42cb1150, 32'h42f7d067},
  {32'hc1faff5b, 32'h43c1da90, 32'h42204ca3},
  {32'hc3d8bf58, 32'h43a5858f, 32'h43461379},
  {32'h42fc3217, 32'hc12bdffc, 32'hc399138e},
  {32'h435a9fa5, 32'hc33888c2, 32'h439599a0},
  {32'hc41a56ad, 32'hc32350b2, 32'hc3212868},
  {32'hc28b9127, 32'h4396f524, 32'hc32e6ff9},
  {32'hc3e5a7af, 32'hc3694218, 32'hc3290a7e},
  {32'h423797fa, 32'hc3b416ba, 32'h43a86b6f},
  {32'h43c4223e, 32'hc27d67e6, 32'h43147656},
  {32'h42edb540, 32'h4114a66a, 32'h4322a9ad},
  {32'h4419a47e, 32'hc3b247a4, 32'hc228a3df},
  {32'h442320b7, 32'h4394b74e, 32'hc295bc79},
  {32'h434c41b4, 32'hc3962d8f, 32'h4237ec9d},
  {32'hc405dcfe, 32'hc3870d68, 32'h4298f79a},
  {32'h42555359, 32'h42d7b753, 32'h432d70b5},
  {32'h43b89a22, 32'hc20397b4, 32'hc300861d},
  {32'h440e32a6, 32'hc3bd0364, 32'h43423d5a},
  {32'hc3c9a471, 32'h432e7855, 32'h421aadca},
  {32'hc2fe74d9, 32'h4144b28d, 32'h44313a96},
  {32'hc307fa04, 32'h421bab3c, 32'hc3a53e65},
  {32'h415a7c08, 32'hc2de2b2b, 32'h437978cb},
  {32'hc229c2da, 32'h43919759, 32'hc18433e0},
  {32'h41d05fa8, 32'h42e9202f, 32'h4247ce5d},
  {32'hc2869a2e, 32'h43ab1dbc, 32'hc1c633d1},
  {32'h42cd7897, 32'h43d71363, 32'h425a385d},
  {32'hc3a6636b, 32'h43b5e541, 32'hc1997598},
  {32'h42861f99, 32'h4384f850, 32'hc390f55e},
  {32'hc136c048, 32'h43b3a88a, 32'h4350b9aa},
  {32'hc2d0099c, 32'hc2705b66, 32'h43814412},
  {32'h41b2da0d, 32'hc3a20042, 32'h439a7a8b},
  {32'hc2a515a5, 32'hc3fca03c, 32'hc33dca4b},
  {32'h42b60e9b, 32'h415c2a58, 32'h438230b6},
  {32'h42c445f7, 32'h43384135, 32'hc2d7fa78},
  {32'h42591ddb, 32'h42daf04f, 32'hc40eb5ea},
  {32'hc3d397e3, 32'h417ae764, 32'h4334f027},
  {32'h4216ad98, 32'hc3509dca, 32'h431223f2},
  {32'h423d6d8f, 32'hc3c64e9d, 32'h425e29c0},
  {32'h4349e2b8, 32'hc3ce1fa6, 32'hc2bf2025},
  {32'hc3398e68, 32'hc24a9f9b, 32'h43860b47},
  {32'h40c983dc, 32'h4252e08a, 32'hc3234ffa},
  {32'hc3b05f3e, 32'hc331e4a2, 32'h4347b189},
  {32'h431ab79f, 32'hc30b59cf, 32'h411f8687},
  {32'h40b2a08d, 32'h43519258, 32'hc3533bba},
  {32'hc32f15cc, 32'h43a7b2cc, 32'hc286e820},
  {32'h435fe2b4, 32'h4265da74, 32'h42888471},
  {32'h43272638, 32'hc2edf35e, 32'h43f4ca9e},
  {32'hc3b75380, 32'hc2f21188, 32'hc3ef59ec},
  {32'hc4366b28, 32'h4342faf0, 32'hc17924f7},
  {32'h44142e24, 32'hc3381242, 32'hc29a1d31},
  {32'hc1888868, 32'hc225ad96, 32'hc0c17cbb},
  {32'h439db79f, 32'hc2d7adb9, 32'hc336f57a},
  {32'hc34e76a0, 32'h42e8f148, 32'h43578e00},
  {32'hc2a0680b, 32'h4380e168, 32'h42f9fa6d},
  {32'hc30dbdb6, 32'h435d11fc, 32'h439a037e},
  {32'h43b3e745, 32'h43b64c91, 32'hc3698be7},
  {32'h431ddeba, 32'hc383dad5, 32'h43883bcd},
  {32'hc1c7bf59, 32'hc38fbdf9, 32'hc0c6c4d1},
  {32'h42632fc0, 32'hc18f445a, 32'hc36a5020},
  {32'hc3cf4ba3, 32'h434600cd, 32'hc1218f91},
  {32'hc335612a, 32'hc3892143, 32'h432b3faa},
  {32'hc3d4c6cb, 32'h43807fb7, 32'hc2ce6ede},
  {32'hc23b839f, 32'hc2ee8583, 32'h4428d26c},
  {32'hc275cd6d, 32'h43c47260, 32'h42bb87f4},
  {32'h42bd5c12, 32'hc30eaf39, 32'hc3e0c805},
  {32'hc3e1c233, 32'h419ccfbc, 32'h421bf842},
  {32'hc3203f3d, 32'hc332a5eb, 32'h428d2302},
  {32'hc387e610, 32'h42bb9bbd, 32'hc3990c50},
  {32'hc40e7bdd, 32'hc36adba1, 32'hc199777d},
  {32'h42e51163, 32'hc2d60287, 32'hc4137261},
  {32'h4341d219, 32'h43be51c8, 32'hc4126b97},
  {32'h4326dfd2, 32'hc3b53636, 32'h438efa1e},
  {32'hc38bc0fa, 32'h429f29cc, 32'h439d20ff},
  {32'h42a060f5, 32'hc380b2ff, 32'hc2e63bc3},
  {32'hc32d4cc5, 32'hc3b307ce, 32'hc254476a},
  {32'hc38c0a35, 32'hc36fc6d7, 32'h42aa0f33},
  {32'h4399d565, 32'hc313e178, 32'h437c8746},
  {32'h43e94a7d, 32'hc2c312a0, 32'hc39a6f1f},
  {32'h4349f8ba, 32'h435d7850, 32'hc3f34073},
  {32'h432b5924, 32'hc29947d1, 32'hc18e26c0},
  {32'hc38603fb, 32'h431c6e6c, 32'h42263f72},
  {32'hc3d54dd7, 32'hc2e4ca73, 32'hc4167c2c},
  {32'hc38d4238, 32'h440fe83d, 32'hc3995f59},
  {32'hc105cdad, 32'h439c97bc, 32'hc2ba00c3},
  {32'hc37d2cd6, 32'h434d899f, 32'h424c7863},
  {32'h433c0097, 32'hc32ca8b0, 32'hc2eb2f24},
  {32'hc2f5e5e1, 32'hc2f6a1f8, 32'h429f9e5f},
  {32'hc227a09a, 32'hc36e092c, 32'h44514f8c},
  {32'hc30cf4fb, 32'h42ce4983, 32'hc34dd73e},
  {32'h44118aea, 32'h43a423d0, 32'hc39b9a78},
  {32'h430eb68c, 32'h3f7f020a, 32'h42dc166f},
  {32'h4364736f, 32'hc35ff6eb, 32'hc2af486c},
  {32'hc3ef7b38, 32'h4379afa7, 32'h41d0d320},
  {32'h4385cbc1, 32'hc312b46f, 32'h43a40ca5},
  {32'h42b5e03e, 32'hc30a9ebc, 32'hc353eb41},
  {32'h4283cfb1, 32'hc3154b79, 32'hc23af833},
  {32'hc2929770, 32'h42bcc114, 32'h437d03b5},
  {32'h43d0088f, 32'hc3165f77, 32'h43499927},
  {32'hc39b28ea, 32'h431d9b64, 32'h4389cb65},
  {32'hc3c1c5c4, 32'h429d27f0, 32'hc2a69210},
  {32'h4272d718, 32'h42c93c6f, 32'h43f5d500},
  {32'hc38697a3, 32'hc23b364c, 32'hc13effea},
  {32'hc3bc094f, 32'h438dde0e, 32'hc2074976},
  {32'h4196d7c0, 32'hc34d933b, 32'h43c6b7bb},
  {32'hc405d9b3, 32'h413cd654, 32'h439a1781},
  {32'hc3103095, 32'h41cdad08, 32'h4357504c},
  {32'hbe84a380, 32'hc261de1c, 32'hc0209320},
  {32'hc2908d43, 32'h439cb685, 32'hc41130b0},
  {32'h4320a2a9, 32'h43853011, 32'h43594e04},
  {32'h430242fe, 32'hc39f0742, 32'h41f9ca98},
  {32'hc36ad4a2, 32'hc3b78a06, 32'hc38153b7},
  {32'hc383d75c, 32'hc414ce55, 32'hc1b92c12},
  {32'h4368c792, 32'hc1d56029, 32'hc136e4b0},
  {32'hc35c129b, 32'hc3c068da, 32'h42884376},
  {32'hc363f575, 32'hc31bed77, 32'hc207ac4c},
  {32'h42632a3e, 32'h4351293c, 32'hc3be2a63},
  {32'hc2aa87d8, 32'h422281eb, 32'h413f2251},
  {32'hc38f2b18, 32'hc34d973d, 32'hc19d97a6},
  {32'hc42469f3, 32'hc3322159, 32'hc210c08a},
  {32'h433f8d40, 32'hc3814da8, 32'h427663ac},
  {32'hc344a685, 32'hc358c6d7, 32'h4391b37e},
  {32'h43964cca, 32'h42ce6bc5, 32'hc36059fa},
  {32'h43af69f5, 32'hc39f277f, 32'h4285f582},
  {32'hc33669c3, 32'h432903e8, 32'h4225f5cf},
  {32'hc3a89cae, 32'h43431c97, 32'h4388601b},
  {32'h440cea50, 32'h42c74d55, 32'h421bcfec},
  {32'h430d3e08, 32'hc2db9958, 32'h4317399c},
  {32'hc3c05be3, 32'hc2620df5, 32'h43acea3b},
  {32'h40359b60, 32'h431512a6, 32'hc38c5474},
  {32'hc459b09e, 32'hc31e49c3, 32'h43071386},
  {32'h406663b8, 32'hc3849b1a, 32'h426cd2f4},
  {32'h43360558, 32'hc338163a, 32'h4222157a},
  {32'hc2ab0656, 32'hc3a0f63c, 32'h43ab058d},
  {32'h44325340, 32'hc3171263, 32'h44152b48},
  {32'hc3be5e7a, 32'h42e2f22e, 32'hc2a36555},
  {32'h416a30f8, 32'h438d1f33, 32'hc36c3ed0},
  {32'h43a7366d, 32'h440d13bd, 32'hc3431f5a},
  {32'hc3b55fbf, 32'h43686d40, 32'hc3b39843},
  {32'hc3b6f2f2, 32'hc318945d, 32'h42c0a8db},
  {32'h4365fc92, 32'hc416f16f, 32'h43be70be},
  {32'h419896dc, 32'hc3850906, 32'h438c6b16},
  {32'hc2519b2e, 32'h41792da5, 32'h4337f50a},
  {32'h4265d038, 32'hc30c98d7, 32'hc319b84c},
  {32'hc3a47c90, 32'hc36897c6, 32'h441da4e8},
  {32'hc130184c, 32'h42078848, 32'h424e9235},
  {32'h43afc2fa, 32'hc2e60c28, 32'hc2b6e103},
  {32'h4351eb5f, 32'hc3ab9501, 32'h43966887},
  {32'hc38c42d2, 32'h42c6eb6f, 32'hc2c61c86},
  {32'h4440430e, 32'h4335bd80, 32'hc320c25f},
  {32'h4300ae7f, 32'hc36a16ac, 32'h42ec0a34},
  {32'hc35e9a88, 32'hc3b82850, 32'hc346efa4},
  {32'hc30c1643, 32'h43a03d88, 32'h433a6b08},
  {32'hc2b3bfbc, 32'h43f256e7, 32'h435073f4},
  {32'h43001053, 32'h4330b968, 32'hc29f2f6a},
  {32'hc3ba17a7, 32'hc3a6f3ef, 32'h436822bd},
  {32'hc2fe3128, 32'h434092f5, 32'hbf8923b9},
  {32'h41fef8b4, 32'hc3202e8c, 32'hc3a40b07},
  {32'h43696250, 32'hc3823280, 32'h414c8f2a},
  {32'hbfd1af00, 32'h4330de7a, 32'h439045e9},
  {32'hc22cbb48, 32'h42338d4f, 32'hc3ea6518},
  {32'h42bccb4b, 32'hc1ad8393, 32'h41df8fb6},
  {32'hc388bb7c, 32'h43ca018c, 32'hc3d2091d},
  {32'h415e3960, 32'hc38eb9ef, 32'hc36ade34},
  {32'h43e4444c, 32'h4399e6f0, 32'hc2818606},
  {32'h4355925e, 32'h432d58ce, 32'hc370a951},
  {32'hc304f10c, 32'hc31502b7, 32'hc266ca5b},
  {32'h42e90cd2, 32'hc3777b41, 32'h43a47ca0},
  {32'hc4182a2f, 32'hc3297ed1, 32'hc3b9d9cf},
  {32'hc01f68e0, 32'h426846b6, 32'h43eb7b31},
  {32'hc2c67de1, 32'hc1d73b5f, 32'hc34866de},
  {32'h4348e147, 32'h43907bcc, 32'h41af2d4f},
  {32'h43642f0a, 32'h439e2d79, 32'h43c5e9cc},
  {32'hc01e5de0, 32'h43e85c72, 32'hc4526f35},
  {32'h431ae362, 32'hc2f69ebb, 32'hc39185e3},
  {32'hc4178aca, 32'hc3b05ad7, 32'hc2e00633},
  {32'h439d37c8, 32'hc3a8dae9, 32'h41b90ce2},
  {32'hc43e467e, 32'hc39b2bdb, 32'h42f8df20},
  {32'hc39c3fcd, 32'h4291768f, 32'h4380b330},
  {32'h42bc2704, 32'hc2c69404, 32'h42bc84e9},
  {32'h443fbb7b, 32'h42f1b716, 32'hc3da4a9e},
  {32'hc43b82d4, 32'hc293f9d4, 32'h41f349b7},
  {32'hc2086301, 32'h42bfe12b, 32'h438e132d},
  {32'hc24d667c, 32'hc3573015, 32'hc2a3cdd1},
  {32'hc36c09c7, 32'hc3186bd8, 32'hc1592a28},
  {32'h42cbe73d, 32'h42dea527, 32'hc261b26a},
  {32'hc37f7738, 32'hc223485e, 32'h42cf6372},
  {32'hc1f78b39, 32'hc37b8af7, 32'h4238bd89},
  {32'h439755d5, 32'h433e594b, 32'h42ea65be},
  {32'h421ce61c, 32'hc18c003e, 32'h43549263},
  {32'hc2be2855, 32'hc3fdd43f, 32'h43007454},
  {32'hc3aa7741, 32'hc2471018, 32'hc32ad9d5},
  {32'hc204325f, 32'h421b1df5, 32'hc1c97b91},
  {32'h439a2a45, 32'hc3922982, 32'h429ca8de},
  {32'hc36decbb, 32'h41f4f94d, 32'h43b04014},
  {32'hc36c5601, 32'h439351b1, 32'h429b48f3},
  {32'h4330a290, 32'h42acabaa, 32'h43840f54},
  {32'h4115a4d8, 32'hc38cb705, 32'hc19bcd5b},
  {32'hc27d9d96, 32'h4253a357, 32'hc3787204},
  {32'h42d55761, 32'hc1a27947, 32'hc2d94796},
  {32'h4323243b, 32'h43635878, 32'hc31e046c},
  {32'hc283c751, 32'h423ae006, 32'h43f8e8de},
  {32'h434f172b, 32'h428625db, 32'hc3127aea},
  {32'h4348152c, 32'hc2949ab1, 32'hc3cd9c7d},
  {32'hc3bac0b6, 32'hc36ee85c, 32'h4363d1a7},
  {32'hc2b69ade, 32'hc37465cf, 32'hc3b0c86e},
  {32'h42b0b219, 32'hc371a9bb, 32'hc42159b6},
  {32'hc37b7f2f, 32'h4119c871, 32'h43ab603e},
  {32'hc3de7bd3, 32'h42f6584d, 32'h42c1f88d},
  {32'h42d782ef, 32'hc3fbd873, 32'h43ce62f7},
  {32'hc419969c, 32'h43db9a17, 32'h42cec2a9},
  {32'hc187316c, 32'hc3bac50e, 32'h43a9b1db},
  {32'h42b1ba54, 32'h42a10724, 32'h4383f5b3},
  {32'h429bc576, 32'hc2d7269e, 32'h42e7d0e8},
  {32'h42f40739, 32'hc409b0c4, 32'h42c52015},
  {32'h43199a3c, 32'h4299ce3b, 32'h43b281b2},
  {32'hc3a7b948, 32'h437a293e, 32'hc3b19c61},
  {32'h438724d4, 32'hc3b62f9b, 32'h42dfa03b},
  {32'h4365cf9c, 32'h43c020cb, 32'h4363df62},
  {32'hc28ad25b, 32'h4418a64c, 32'hc1787030},
  {32'hc347d815, 32'hc2c692b4, 32'hc39f9731},
  {32'h43967f1f, 32'hc3e2ad18, 32'hc318f7cb},
  {32'h43665a24, 32'hc26149ac, 32'h41b30119},
  {32'hc3961d14, 32'h438aae75, 32'h4345e6f2},
  {32'h427c54c7, 32'hc31d6088, 32'hc39b965d},
  {32'hc2d804c2, 32'hc238acf4, 32'hc2269515},
  {32'hc29f4b4b, 32'hc30f8d2c, 32'h41c95855},
  {32'h42f46260, 32'h43c7fcff, 32'hc2c2e174},
  {32'hc3335f22, 32'hc384143e, 32'h42b7f59f},
  {32'hc385a349, 32'hc1a693c2, 32'hc408eb43},
  {32'h43752576, 32'hc29ba6be, 32'hc1f5c556},
  {32'hc27ad168, 32'h429fa052, 32'h425cfa30},
  {32'hc42144d7, 32'hc2a1e48c, 32'hc2874e6f},
  {32'hc37b77c9, 32'h43eb0a24, 32'h41343714},
  {32'h4417ce30, 32'h41ee7806, 32'hc4152575},
  {32'hc1f544f8, 32'h4294aedb, 32'hc07cd83f},
  {32'hc2ff6b62, 32'hc33f0e91, 32'h43e19bf5},
  {32'hc4078286, 32'h43a2c606, 32'hc3b77114},
  {32'hc3f1659c, 32'hc3e4f9d2, 32'hc3af1490},
  {32'h433fba08, 32'hc32b5943, 32'h42fdd1fe},
  {32'hc3103e45, 32'h430f8bd2, 32'hc2671bbc},
  {32'h43276aea, 32'h42855ac6, 32'hc3c00207},
  {32'h42132d8c, 32'h4388f911, 32'h43c69199},
  {32'h43159177, 32'hc33dcb64, 32'hc34595e4},
  {32'hc3f0def8, 32'h43cd8497, 32'h436198a3},
  {32'h43883736, 32'h423d1235, 32'h43b095dc},
  {32'hc2ddbffd, 32'hc2189871, 32'h4390709a},
  {32'hc1212f34, 32'hc307b4dc, 32'h3ea01800},
  {32'h438e3013, 32'hc3438149, 32'h442a328c},
  {32'h427070db, 32'hc3660af1, 32'hc31a5ceb},
  {32'hc2b6c27c, 32'hc2deb632, 32'h43652217},
  {32'hc31921e4, 32'hc34329c6, 32'hc3d7478b},
  {32'h43aad8e2, 32'h42b4a018, 32'hc203320f},
  {32'h42093417, 32'h4387792e, 32'hc32b1b9c},
  {32'h4243dbe8, 32'h433205f2, 32'hc2d60249},
  {32'hc3467f24, 32'hc3af83f1, 32'hc1873f73},
  {32'hc31972eb, 32'hc382a1bc, 32'hc371edfb},
  {32'h43c1951c, 32'hc3e5e863, 32'hc1a14ff8},
  {32'h42096649, 32'hc229de31, 32'hc16b6ccc},
  {32'hc2877d40, 32'hc393f74d, 32'hc39dbc0b},
  {32'hc39680c7, 32'h4433e961, 32'h41f18e74},
  {32'h4320abfe, 32'hc2f3b9de, 32'hc30097b5},
  {32'h4236bba8, 32'hc2b56179, 32'hc30c4379},
  {32'h43e56aac, 32'hc2864b59, 32'hc316c6c0},
  {32'hc2cf7bc7, 32'h4360584c, 32'hc294bd43},
  {32'hc3c84b5a, 32'h40a32820, 32'hc2abea84},
  {32'h43d41988, 32'hc34ddbcf, 32'hc24d2916},
  {32'hc31d469e, 32'hc309d78f, 32'hc3854349},
  {32'h42444330, 32'h41ccd1a2, 32'hc3480c7e},
  {32'h430bd1f0, 32'hc3c88a09, 32'hc3a9221a},
  {32'h419539bc, 32'h433b8586, 32'hc33c7cd4},
  {32'h43e29fd6, 32'h43aad034, 32'h435e31a1},
  {32'h435a96db, 32'h4363e1d7, 32'h439688b3},
  {32'hc38b31a6, 32'h4358504a, 32'h4388fd47},
  {32'h42a3e206, 32'hc2f76623, 32'h42df651a},
  {32'h423d2cfa, 32'h43aa331b, 32'h4264ed90},
  {32'h4241fcd2, 32'hc3d6cec6, 32'h431e146d},
  {32'h435f3ad4, 32'hc3c7ee2f, 32'h4314c762},
  {32'h43a71458, 32'hc35a41e5, 32'h42ab5428},
  {32'hc3f15c47, 32'hc3ac2458, 32'h42483760},
  {32'h44098e58, 32'hc26ae72c, 32'h443bb712},
  {32'hc444a9b0, 32'h4239f261, 32'h42cd699f},
  {32'h43807231, 32'h433b1ddb, 32'hc381a05f},
  {32'hc1238774, 32'hc32150c0, 32'hc31c352a},
  {32'h43c3b9b6, 32'hc3995e40, 32'h43368120},
  {32'hc39de2ed, 32'hc396e4d7, 32'hc307c997},
  {32'hc2cb4cfb, 32'h42fde337, 32'h4202b760},
  {32'h4347f286, 32'hc372ff78, 32'hc245da5e},
  {32'hc3378739, 32'h42e34fd0, 32'h4273e602},
  {32'h427d97b0, 32'h42e7116a, 32'hc393d5d3},
  {32'hc1a5ecd8, 32'h43284336, 32'h44164b71},
  {32'h425a8787, 32'h439e791a, 32'hc32f41c0},
  {32'hc38ba0a5, 32'hc2ff4d4a, 32'h43a7280a},
  {32'h434d580c, 32'hc1c5b5ff, 32'hc32aef96},
  {32'hc3a5c26e, 32'h42e2f9f8, 32'hc2debfcf},
  {32'hc334b1a2, 32'hc31a4edc, 32'hc06893f6},
  {32'h4425ea4f, 32'hc398629d, 32'h43b56b55},
  {32'hc3b8ad34, 32'h43e42ff9, 32'hc3dd76ed},
  {32'hc2a210cf, 32'h43a437ba, 32'hc3fd40c1},
  {32'hc3bfa55c, 32'hc3620feb, 32'hc35df502},
  {32'h42670ce4, 32'hc2f13739, 32'hc2a1a1a1},
  {32'hc3d42326, 32'h42f4fa86, 32'h4315af9e},
  {32'h43f3beda, 32'hc327404c, 32'hc3661680},
  {32'hc247d015, 32'hc310a00d, 32'hc3080d4f},
  {32'h439e568e, 32'h437b7d17, 32'h415f05cc},
  {32'hc1659402, 32'h43ea9448, 32'hc207c3c0},
  {32'h4290554d, 32'h43a20392, 32'hc3c1838f},
  {32'hc0ec35dd, 32'hc3926d23, 32'hc19f15db},
  {32'h43e93b42, 32'hc3b156c7, 32'hc3a44768},
  {32'hc38115e6, 32'h436802e2, 32'h432289da},
  {32'hc2a8c0ce, 32'h42d707e4, 32'hc1e36bc9},
  {32'h43ad7ddd, 32'h42cf63f5, 32'h43376aa0},
  {32'hc395c036, 32'hc3c60043, 32'hc381b958},
  {32'hc3c599be, 32'hc35763e6, 32'hc41ce3a9},
  {32'hc3a57eee, 32'h42d8f76e, 32'h43436440},
  {32'hc339eba7, 32'hc29f8488, 32'hc2f6599b},
  {32'hc314a51e, 32'h4341516e, 32'hc3ad5e3a},
  {32'h4300288a, 32'h418bb2c9, 32'h42d41bdb},
  {32'h4374f0f6, 32'hc323aa7c, 32'hc36545d8},
  {32'hc27656f4, 32'hc31791f4, 32'h42049ddf},
  {32'h43840944, 32'h41b6b6d6, 32'h433cdae5},
  {32'hc410ac21, 32'hc3603dc7, 32'h4368987b},
  {32'h4338f010, 32'h42461330, 32'h439127a6},
  {32'h410e5b80, 32'h42e39561, 32'h43ff279e},
  {32'hc3c84bfe, 32'h437d8a27, 32'hc3a2286f},
  {32'h419a4408, 32'h42bc1c6e, 32'h40f71f5c},
  {32'h432b6230, 32'h439bb781, 32'h42d4de9a},
  {32'hc1f9d4fc, 32'h432d13cf, 32'h41bbecef},
  {32'hc2390cea, 32'hc282b86c, 32'h43ea6315},
  {32'hc257e4c2, 32'h4386f1d4, 32'hc2c3b007},
  {32'hc2a49b9b, 32'h434c0924, 32'hc389d450},
  {32'hc3030e92, 32'hc2372234, 32'h43b3d3c2},
  {32'h41382bb4, 32'h4371762f, 32'hc3d7d006},
  {32'hc08372e2, 32'h4351243c, 32'h43a0fe0a},
  {32'h4392df88, 32'hc34ad81f, 32'h439cdb8e},
  {32'h438fa9b8, 32'hc23f2e3b, 32'hc2600209},
  {32'h43295c8b, 32'h42a84957, 32'h420201a6},
  {32'h43a0e677, 32'h42eb9658, 32'hc2fb647f},
  {32'h43c42b52, 32'hc2d5a337, 32'hc3c5740c},
  {32'hc39cf202, 32'h4237c13e, 32'hc3651f94},
  {32'hc2ddb303, 32'hc3d3f8fe, 32'hc225f5ab},
  {32'h426110c4, 32'h43c9cc78, 32'h42af7da6},
  {32'h43a1f191, 32'hc384011c, 32'hc311b5e1},
  {32'h421b46fd, 32'h42917375, 32'h42e91b5c},
  {32'hc3d9a8ca, 32'h422ba9e6, 32'h43ba1336},
  {32'hc3137086, 32'h43a92e15, 32'hc3c82733},
  {32'h42a82b37, 32'hc39f5ec1, 32'h43657806},
  {32'hc31f0849, 32'hc367dd64, 32'h43246075},
  {32'hc4032b58, 32'h433325e1, 32'h43865156},
  {32'h43fb0efc, 32'h42f91549, 32'h432ae027},
  {32'h43a86def, 32'h43b424af, 32'h429f6aa8},
  {32'hc2bcff4a, 32'h40b9f4ca, 32'h43a469b7},
  {32'h4302f074, 32'h429b80e4, 32'hc306982e},
  {32'hc2d1978d, 32'h41297500, 32'h4175f17f},
  {32'h42b7af73, 32'h4316d0ee, 32'h438eabaf},
  {32'h4383ddfc, 32'hc387eece, 32'h433b4d1c},
  {32'h4051e400, 32'hc38962df, 32'h436232b0},
  {32'h423fb31f, 32'hc2709547, 32'h421c4912},
  {32'h43d53fc9, 32'hc396cd15, 32'hc2c04b26},
  {32'h42dda252, 32'hc342bbc3, 32'hc3b95f53},
  {32'hc2ccaa80, 32'h4405ad48, 32'hc292404b},
  {32'h429266c1, 32'hc291795a, 32'hc1b6daff},
  {32'hc3364147, 32'h4282ee5d, 32'hc1c68d6f},
  {32'hc2d01ef4, 32'hc293dfff, 32'h43005cdb},
  {32'hc3ce1c5a, 32'hc1c6363a, 32'h40d05b3e},
  {32'h43c4624e, 32'hc2f2d87b, 32'hc37c8efe},
  {32'h432d61e9, 32'hc3309f85, 32'hc3b83183},
  {32'hc3b768ff, 32'hc3a3bb41, 32'hc416b0a2},
  {32'h43632fad, 32'hc3b48359, 32'hc251b751},
  {32'h430ccbf3, 32'hc354f27a, 32'hc304f96d},
  {32'hc39a2c77, 32'hc25b6ef4, 32'hc2500ade},
  {32'hc2a54d9e, 32'h4291e81f, 32'h43a3974a},
  {32'hc2909e88, 32'h43a92ebb, 32'hc36775b1},
  {32'hc38d7786, 32'h439a2f72, 32'h43de3f38},
  {32'hc28b2059, 32'hc368db95, 32'h433a3ba5},
  {32'h4345c115, 32'hc261f37d, 32'hc2d15df0},
  {32'hc34e907e, 32'h43aa3776, 32'hc397c60e},
  {32'h43697726, 32'hc320b1e1, 32'hc3b1b1e6},
  {32'hc3658d18, 32'h42e7f6e3, 32'hc3a525ea},
  {32'h4122ea24, 32'hc341a49a, 32'hc38641b4},
  {32'h435527fa, 32'h43bbece4, 32'h425b5bf6},
  {32'hc3201c1e, 32'h4319385d, 32'hc3992514},
  {32'hc26ee967, 32'hc2f5b5fb, 32'hc397b8f5},
  {32'h43fd16f3, 32'hc37900e1, 32'h43a38803},
  {32'hc32425f6, 32'hc22342c8, 32'h421d6209},
  {32'h4341e1c9, 32'h42a5d8d0, 32'hc2119b7a},
  {32'hc1646118, 32'h43027c7f, 32'hc37c8e80},
  {32'h42b0c5ee, 32'hc2b76554, 32'hc2e22bfe},
  {32'h439baed4, 32'h44035059, 32'h435286de},
  {32'hc387d638, 32'h41d84b87, 32'hc37119a6},
  {32'hc386f3c6, 32'h438ed93a, 32'hc2e7dc33},
  {32'hc2993455, 32'hc33926b6, 32'h43273ae1},
  {32'hc289cf4c, 32'hc3886504, 32'hc3101964},
  {32'hc218b914, 32'hc34cb233, 32'h43881060},
  {32'hc317a17f, 32'hc2cc3bbf, 32'h42ecd0c5},
  {32'hc225c7d5, 32'h439278a1, 32'hc2aec2ce},
  {32'h4424c06a, 32'hc3b802df, 32'hc32600b1},
  {32'hc4339c38, 32'hc2d688fe, 32'h42ce4991},
  {32'hc23f042f, 32'hc35279b4, 32'h43fc955a},
  {32'h4384c203, 32'h436a7254, 32'hc3240161},
  {32'h43c10e33, 32'hc38cfd60, 32'h426ab76e},
  {32'h4438c7e0, 32'h426706eb, 32'h3ff85d90},
  {32'hc379b66b, 32'h438231b7, 32'hc2d09db1},
  {32'h422b0a30, 32'hc314e0d9, 32'h42a7c6cd},
  {32'h3f507d00, 32'h428d5301, 32'h43e110a3},
  {32'hc35374c0, 32'hc3c17a72, 32'h42edbe26},
  {32'h43f330fb, 32'h43873bf6, 32'h43e85413},
  {32'hc2884126, 32'h43e8a81d, 32'h42e6000f},
  {32'h421d9d50, 32'h42ad6c84, 32'hc3c75902},
  {32'hc2fef942, 32'hc31afe00, 32'hc3564760},
  {32'h4335855b, 32'hc3df18d8, 32'h43d4e3f1},
  {32'hc2f728ca, 32'hc38bea80, 32'h400a514e},
  {32'h427b69d8, 32'h42bdd300, 32'h4367f191},
  {32'h431bedb2, 32'hc395409e, 32'hc380e495},
  {32'hc4335441, 32'h436c9630, 32'h44087bad},
  {32'h437afcdf, 32'h428c4149, 32'h43807696},
  {32'hc2843cd1, 32'h439e6230, 32'hc2e3546e},
  {32'hc31573fb, 32'hc2d1bb3b, 32'h435c71cb},
  {32'h430f652d, 32'h43f5080a, 32'hc3abdf64},
  {32'h43e6448a, 32'hc415cd95, 32'hc3861634},
  {32'hc2c917ff, 32'hc316a263, 32'hc10d40fc},
  {32'h44096b85, 32'h42a5bdb2, 32'hc2cc2dab},
  {32'h43b3de92, 32'hc30d59d6, 32'h43ae1a98},
  {32'hc3e66d50, 32'h43b81647, 32'hc371f78a},
  {32'h437e4b95, 32'h434a7495, 32'hc2da2e28},
  {32'h43c7aeed, 32'h415f5cb3, 32'h43ba2e8c},
  {32'h426cb8d0, 32'hc3a6ee18, 32'h42e886a3},
  {32'hc384f873, 32'hc38094f7, 32'hc3436503},
  {32'h42fe476c, 32'hc330221d, 32'h432f8ce2},
  {32'h43fdfd3c, 32'hc1cae18a, 32'hc36fb589},
  {32'hc2c3f8ac, 32'hc3299ada, 32'hc3510a44},
  {32'h44016184, 32'hc3924ba4, 32'h433afa45},
  {32'hc30ae6c5, 32'h4409d15b, 32'h43e73052},
  {32'hc405cd05, 32'h425e0d43, 32'hc3b3ac98},
  {32'h431770df, 32'h4402a025, 32'hc342c36f},
  {32'hc385c5ad, 32'hc3855e05, 32'h431f9116},
  {32'h433e2abf, 32'hc21d4d03, 32'h4335839c},
  {32'h43a1a0eb, 32'hc2b2b198, 32'h437b13c2},
  {32'h42e1bfa2, 32'hc21ee970, 32'hc3e7bb0a},
  {32'hc2a9bc96, 32'hc3ced621, 32'h4455bb77},
  {32'hc1c37730, 32'h4409f4e7, 32'h433d187d},
  {32'h430461a3, 32'h439b6bbd, 32'hc4178d58},
  {32'h4284602e, 32'hbf0e3085, 32'h43fd1332},
  {32'h43f2b9a4, 32'hc25883fc, 32'hc2eb8b69},
  {32'h43942d79, 32'h42a2817b, 32'hc3415b04},
  {32'hc24b4504, 32'h4381a174, 32'h41bf00fe},
  {32'h406e3300, 32'h42856559, 32'h427234ec},
  {32'hc3d86b95, 32'hc3d49d1d, 32'h42554374},
  {32'hc30921c3, 32'h42888eb0, 32'h43d2239c},
  {32'h42800275, 32'hc31c1bea, 32'h43c0133f},
  {32'h43655bc4, 32'hc252ce55, 32'hc35ccbc7},
  {32'hc33b2566, 32'h43a52029, 32'hc356e869},
  {32'h433782b2, 32'hc2d9838e, 32'hc30adb3d},
  {32'hc267e88d, 32'h4278c744, 32'hc1c8b74f},
  {32'hc3d48ed4, 32'h4347653c, 32'h43ce6c78},
  {32'h43950af6, 32'hc38d6f71, 32'h408a8ce2},
  {32'hc33abfd0, 32'h42ebd550, 32'hc27802bf},
  {32'hc2f824ae, 32'h43016f80, 32'h414634dc},
  {32'h441fa32a, 32'h43d5c19b, 32'h444b446f},
  {32'h432ba327, 32'h43141645, 32'hc3449de1},
  {32'h43ae9d19, 32'h42ef5e26, 32'hc3dee3d4},
  {32'h43d5d54b, 32'h4405aa6b, 32'hc3bf5281},
  {32'hc3b6048c, 32'h41169efb, 32'h3f97979d},
  {32'hc095eea4, 32'hc33b553e, 32'hc29723fc},
  {32'hc2520fd6, 32'hc2eece63, 32'hc25a0edb},
  {32'hc3e9cf99, 32'hc3ad19ed, 32'hc33ab87a},
  {32'hc2b3e5be, 32'h42f4a491, 32'hc2e05f45},
  {32'h438f65f3, 32'hc3ed1009, 32'hc3a5286d},
  {32'hc3d7b2c3, 32'h439dd96f, 32'h43a22ab8},
  {32'h43072500, 32'hc2a99cbe, 32'h43ecfb5e},
  {32'h43ad6898, 32'hc40cfc62, 32'hc2026752},
  {32'hc32a29ae, 32'hc2a88ae9, 32'h430ce925},
  {32'h43cc99fd, 32'h436ca5be, 32'hc2d8dc76},
  {32'hc3711d7b, 32'hc34ba3e5, 32'h428ea93a},
  {32'hc38a7b8a, 32'hc32f0920, 32'h43455c75},
  {32'h43a3c286, 32'hc30d8c7e, 32'h4218319f},
  {32'hc3790708, 32'h4354ce3c, 32'hbfbe005a},
  {32'hc27f70ca, 32'h41983946, 32'hc3ab6a46},
  {32'hc3df1b0c, 32'hc224479d, 32'h43b264a2},
  {32'h42599368, 32'hc3391c99, 32'hc3af6d45},
  {32'h41eabab7, 32'hc23fd4ca, 32'hc38f9356},
  {32'hc2ba9dc3, 32'h436354a1, 32'h438cb221},
  {32'h438a2ce5, 32'h43a3f101, 32'h403020f4},
  {32'hc3147664, 32'h438b1c7f, 32'h42c96a61},
  {32'hc38f040e, 32'h4322fea3, 32'hc390c954},
  {32'h433843c8, 32'hc35cf484, 32'h43285792},
  {32'hc3c50632, 32'h435205f0, 32'h400a0e77},
  {32'hc373bb3e, 32'hc1ba842c, 32'hc295cee1},
  {32'h43b35d5c, 32'h43f36547, 32'h43063fe8},
  {32'hc348d61a, 32'h438d1c91, 32'hc3373377},
  {32'hc3e09f12, 32'h43569354, 32'h42108e96},
  {32'h4380fdba, 32'hc38566df, 32'hc3ebc48a},
  {32'h428d6508, 32'hc387c684, 32'hc3763e49},
  {32'hc1c7dea5, 32'hc10008fc, 32'h435c12bb},
  {32'hc2d3b133, 32'h4268c54d, 32'hc457ed94},
  {32'hc39ef6cf, 32'h4329d9e2, 32'h42e6d7c3},
  {32'h4320e96f, 32'h430c2971, 32'hc33cd2c2},
  {32'hc24f30d0, 32'h43456657, 32'h42f79f93},
  {32'hc30759b0, 32'hc108b25b, 32'h43aa8379},
  {32'hc28be9c6, 32'hc2027f7a, 32'hc3590b7a},
  {32'h43372619, 32'hc4058808, 32'hc303e694},
  {32'hc3c0178d, 32'hc35f740f, 32'h4351e211},
  {32'h4418dca2, 32'hc2e87669, 32'h42851fa4},
  {32'h431d46db, 32'h4351959a, 32'h4234d14b},
  {32'h43c168ea, 32'hc28816a1, 32'hc35e2402},
  {32'h4193bc44, 32'h438ddc0d, 32'hc16418a3},
  {32'h434d0d14, 32'h422277ab, 32'h42e1cb01},
  {32'h42bedbfc, 32'hc18183db, 32'h41c3fd08},
  {32'hc3b049ea, 32'hc3d70cf1, 32'h4320e376},
  {32'h436c9668, 32'hc318f77a, 32'h41adea87},
  {32'h440d7224, 32'h40830daf, 32'hc2ec4064},
  {32'hc40b7f4b, 32'h42ab2fab, 32'hc443053e},
  {32'h431741b6, 32'hc31961c0, 32'hc34a70cc},
  {32'hc3955fb8, 32'h4218c41a, 32'hc3c1f8ac},
  {32'h41a59960, 32'h43325203, 32'h41b2dd2a},
  {32'h432a1f93, 32'h43af7c9b, 32'hc2e47f0c},
  {32'hc30c76b0, 32'hc2016b1c, 32'hc40fdcc7},
  {32'h435bb603, 32'hc3982ae2, 32'h41fd923e},
  {32'h41b96e3d, 32'hc39edf39, 32'h42f3e117},
  {32'hc329617a, 32'hc3afc426, 32'h43173b0c},
  {32'hc399a61f, 32'h40c3726a, 32'h41dbe80b},
  {32'hc367c438, 32'h41e6fe58, 32'hc3de9727},
  {32'h4364010c, 32'h43538370, 32'hc3186719},
  {32'h426fd3ee, 32'h4300d586, 32'hc284277b},
  {32'h418350af, 32'h4336d732, 32'hc3d3354b},
  {32'hc2cbfd0a, 32'hc3f96cb5, 32'h4400481a},
  {32'hc2c48667, 32'h431ff10b, 32'hc384b07e},
  {32'h43be4979, 32'hc334d73e, 32'hc365a1ee},
  {32'hc31bbe0c, 32'hc32a71ba, 32'h437b81cc},
  {32'hc302bdd2, 32'h43eb4022, 32'h437dcf82},
  {32'hc3619d0d, 32'h4374337a, 32'h43858070},
  {32'h434b0b04, 32'hc3057a60, 32'hc38e8cee},
  {32'hc36d1eac, 32'h4400d9e7, 32'hc3b0cfdf},
  {32'h41bd5dc5, 32'h438272df, 32'hc4409e44},
  {32'h42402398, 32'h43811538, 32'hc31e22f2},
  {32'hc302beda, 32'hc2f6c262, 32'h42d95d1e},
  {32'h43461fa7, 32'hc2ce7528, 32'h42bfa7c8},
  {32'h43139714, 32'hc3450f0f, 32'h432940a2},
  {32'h4441461d, 32'hc40b0b72, 32'h43e111da},
  {32'h4345936e, 32'h42c2ae9a, 32'h4326d6d2},
  {32'hc2bae212, 32'h438b07ac, 32'hc2f717ca},
  {32'hc3535836, 32'h43b12b9c, 32'hc37c2a69},
  {32'h43551ab2, 32'h43beddcc, 32'h436957b0},
  {32'hc38e98f7, 32'h4390bbfe, 32'hc3fce868},
  {32'hc3f109f3, 32'hc3a70ec0, 32'h43839860},
  {32'hc30d1cb8, 32'hc35f595b, 32'hc16fb81a},
  {32'hc2a443ba, 32'hc31b28dc, 32'hc3bcd412},
  {32'h438c9152, 32'hc41e44be, 32'h43eed5e8},
  {32'h43047427, 32'h428e7bd3, 32'hc39088e9},
  {32'h431f1a56, 32'hc3c3fa40, 32'h43ab27d3},
  {32'hc2a8bfb6, 32'hc2041a99, 32'hc37ca170},
  {32'hc3836e09, 32'hc30cfaea, 32'h41d866b6},
  {32'hc2ae928d, 32'hc30e3cce, 32'h42dc323c},
  {32'hc32782e4, 32'h437b446b, 32'hc3f08774},
  {32'h431e252c, 32'hc314f46d, 32'hc392b387},
  {32'h4091b007, 32'hc40350d8, 32'hc294b028},
  {32'hc2e5aa58, 32'hc20eaceb, 32'h4108e6e3},
  {32'hc196232a, 32'hc34869f0, 32'h429cd7c4},
  {32'h4367a7f2, 32'hc373faf0, 32'h427e679f},
  {32'hc3eebca5, 32'h4273419c, 32'h4267c915},
  {32'hc24c7618, 32'h4369bd4a, 32'h43c4c68a},
  {32'h413aade7, 32'h43e40123, 32'hc34014e9},
  {32'hc454b739, 32'h412cb958, 32'h43e252e0},
  {32'h43a15080, 32'h432171d2, 32'h432728de},
  {32'h43abb51f, 32'hc2be6ac1, 32'hc22be550},
  {32'hc38c5788, 32'hc1949dca, 32'hc39a1238},
  {32'h43038d4a, 32'hc3b009bd, 32'hc305aba1},
  {32'hc445f692, 32'hc3663a84, 32'hc29f6a7d},
  {32'hc1c1ea05, 32'hc3e468fd, 32'hc35d82e0},
  {32'hc3331390, 32'h43efeac2, 32'hc3b675df},
  {32'hc35025ce, 32'h42fde4b6, 32'hc39ae4b9},
  {32'h42f078a0, 32'hc2a8a74f, 32'hc359862c},
  {32'h43b2e4bc, 32'h43b1f1e4, 32'hc3261dc5},
  {32'h433bf583, 32'h42c03dc7, 32'h42afddb5},
  {32'hc213a7c1, 32'hc1b6edba, 32'hc24572c6},
  {32'h43e5e5c9, 32'hc3abd4ce, 32'h43255078},
  {32'hc15c66c0, 32'h433f8bbb, 32'hc2a38d9b},
  {32'hc29b088f, 32'hc35e41bd, 32'hc31681a0},
  {32'h41ceb9f8, 32'hc3d014fa, 32'hc3e9c258},
  {32'hc29d1989, 32'hc3c7996a, 32'h439d66b1},
  {32'h3f4a0c80, 32'h438219cc, 32'h425e68ad},
  {32'h43953937, 32'hc329abdf, 32'hc414620e},
  {32'hc34a3528, 32'hc404ec61, 32'hc423e072},
  {32'hc3859501, 32'h435bcccd, 32'h43da3703},
  {32'h4342fda0, 32'h439de3c6, 32'hc3503fe2},
  {32'h441ea794, 32'h4250b0e6, 32'h42dca83e},
  {32'hc3ebae80, 32'h4303e275, 32'h43ce06ae},
  {32'h43cf4083, 32'h43556a62, 32'h42ee5c71},
  {32'hc3b543c9, 32'hc269a188, 32'hc4107f72},
  {32'hc42bede0, 32'h43882c9b, 32'hc2bd5408},
  {32'h43cbe1ea, 32'h42c2c7d5, 32'hc3513110},
  {32'hc2f7a4de, 32'hc408055a, 32'h439842c0},
  {32'h42db6c12, 32'hc2b8136e, 32'hc37cbc23},
  {32'h42dcecdc, 32'hc1d5296c, 32'h443881b7},
  {32'h430f7214, 32'hc231a219, 32'h42870456},
  {32'hc30fb597, 32'h42b0118a, 32'hc4012f9d},
  {32'h42aacd22, 32'h427febb0, 32'hc32a1b14},
  {32'hc397b48e, 32'hc3f0531a, 32'hc32d3201},
  {32'h42953f88, 32'hc31828ae, 32'h429f6d34},
  {32'h4366af94, 32'hc3ae8939, 32'h423632d5},
  {32'hc3698bc2, 32'hc3a94d8e, 32'hc252f8f4},
  {32'hc11ee1cc, 32'hc36d165b, 32'h43291461},
  {32'hc36ed788, 32'hc06051a8, 32'h41d498ae},
  {32'h42d1d788, 32'hc3c6a4fd, 32'h438e0b87},
  {32'h433f3a53, 32'h429a69ec, 32'h42fba90d},
  {32'h432c8b51, 32'h440a1ded, 32'hc2d93746},
  {32'hc3f079e7, 32'h4372b570, 32'hc27d36ea},
  {32'hc18272b8, 32'hc3916cc2, 32'hc32d0956},
  {32'hc396abac, 32'h41b12b02, 32'hc38696c4},
  {32'hc4042e5a, 32'hc1c95e5b, 32'h4300e379},
  {32'hc3195e58, 32'h432320fc, 32'h43478ad4},
  {32'h438719bd, 32'h43516d84, 32'h43e72250},
  {32'hc2a9bb2c, 32'h43b14aa9, 32'h40417cb0},
  {32'h436a78e1, 32'h43ef5319, 32'h43ba714b},
  {32'h41bd760c, 32'hc35ab1c1, 32'h4380837a},
  {32'hc370a00a, 32'hc393fe92, 32'h43e87a7f},
  {32'hc21278ba, 32'h424726f4, 32'h42cdcd4c},
  {32'h43d99aac, 32'hc3159a57, 32'hc2e9aa8a},
  {32'h42aacaa9, 32'h4232b33b, 32'h402f28af},
  {32'hc38e0549, 32'hc1a13be2, 32'hc3900ab8},
  {32'hc3a543d1, 32'h439d7b38, 32'h42be1aa1},
  {32'h443e1cad, 32'h431bca8c, 32'hc33dc3e9},
  {32'h439d3912, 32'h440d8dfb, 32'hc36b5066},
  {32'hc1c00615, 32'hc2b03a9a, 32'hc098512e},
  {32'hc2bfa396, 32'hc310b854, 32'h42136a58},
  {32'h4211a312, 32'hc33aeb1e, 32'hc2a28add},
  {32'hc260d300, 32'hc3440bdd, 32'hc158ced1},
  {32'hc3f183f8, 32'hc3098765, 32'h4164c9ba},
  {32'h436c6a16, 32'hc2f22a95, 32'hc31f4316},
  {32'h43a99740, 32'hc3b47085, 32'hc3a0f679},
  {32'hc36b1462, 32'hc2c071e0, 32'h4161338a},
  {32'hc3af5630, 32'hc35e90ed, 32'h4360230d},
  {32'h4348e2c1, 32'h43bcd8ad, 32'hc3869ee2},
  {32'hc40e3b93, 32'h419f1fc2, 32'h43b2e979},
  {32'hc2b62bb7, 32'h427366f4, 32'hc3d2e996},
  {32'h439d95cf, 32'h434c3203, 32'h43a85ae8},
  {32'hc412ae1d, 32'h43a14638, 32'hc248ef35},
  {32'hc3d578b4, 32'h434a142b, 32'h425057c4},
  {32'hc3f73663, 32'h436fb165, 32'h4378b0dd},
  {32'hc2b4fe43, 32'hc2520235, 32'hc2d765e6},
  {32'hc40b5f13, 32'h43a2c791, 32'h43238811},
  {32'hc3295127, 32'hc395f6c4, 32'hc319b4d2},
  {32'hc389134e, 32'h4399eb61, 32'hc29e6908},
  {32'hc328e58e, 32'hc239094e, 32'h43c51028},
  {32'h4300ca34, 32'h430e3ccf, 32'h43fdc1e2},
  {32'h41a99f4a, 32'hc38c6373, 32'h436aaac7},
  {32'hc2b8613e, 32'hc31ee214, 32'h4269e076},
  {32'h42f57b12, 32'hc36abaca, 32'h4400e491},
  {32'h42e99e30, 32'h4303ef24, 32'h4380fb5b},
  {32'h4393119b, 32'h4396d57c, 32'hc0587b10},
  {32'hc1861fa2, 32'hc2f8d27c, 32'h438ab86a},
  {32'hc34601db, 32'hc3a57985, 32'hc3262d9f},
  {32'hc3c05f8c, 32'hc40fa511, 32'h43a06d16},
  {32'h42a23089, 32'h41441e22, 32'hc3387742},
  {32'h423c6a93, 32'hc3da07cb, 32'hc40ba7eb},
  {32'hc300b2ed, 32'hc22b9e9e, 32'h439fce47},
  {32'hc263d75d, 32'h42eda4a0, 32'h43a14738},
  {32'h4409e9ec, 32'hc39d1102, 32'h438ddbd1},
  {32'h433eb45a, 32'h42693040, 32'hc151b2cc},
  {32'hc3180b4c, 32'hc2b6df9e, 32'h430b5f91},
  {32'h424ab282, 32'hc2224066, 32'h4345aa91},
  {32'h40fb1300, 32'h436a9b2a, 32'hc3370680},
  {32'h4209fb0a, 32'hc3c527cf, 32'h437d7927},
  {32'h4359a95d, 32'hc192b1de, 32'h4183eeae},
  {32'hc3b54070, 32'h412ad05e, 32'hc3e5a6ba},
  {32'hc250429a, 32'h43a0c1db, 32'h41a0e2fd},
  {32'hc347a4dc, 32'h438f853b, 32'h4302172a},
  {32'hc3e762b1, 32'hc3124a58, 32'hc2a770b3},
  {32'h435bbe88, 32'hc3bb7206, 32'h430d9b50},
  {32'hc40889b2, 32'hc33dfe06, 32'hc37aed02},
  {32'hc37faea6, 32'h431e47f5, 32'hc2459c92},
  {32'h4422d129, 32'h438e9f02, 32'h44160236},
  {32'h4256949e, 32'hc30ad732, 32'hc2ad71b6},
  {32'h432f1f41, 32'hc128bd41, 32'hc3798646},
  {32'h42a37858, 32'h42d3f7f7, 32'h43e88716},
  {32'hc3b91d9f, 32'hc3ed52f9, 32'hc317e85e},
  {32'h3fb71640, 32'h436df802, 32'hc346e6c9},
  {32'h42606b68, 32'h433865e1, 32'h42bd988d},
  {32'h435d3689, 32'h4317a0b0, 32'hc395ab5b},
  {32'hc344339f, 32'hc027adbc, 32'h4281091e},
  {32'h439abb26, 32'hc3c128b5, 32'h428b0f0c},
  {32'hc3c50512, 32'hc31cb4c3, 32'hc3003496},
  {32'hc396c6b6, 32'h438b7a26, 32'h43ca30cc},
  {32'h4362132e, 32'hc3247434, 32'hc32ba18f},
  {32'h42a98396, 32'h42fedd63, 32'h43ad600f},
  {32'hc31662c3, 32'h42a04ed7, 32'hc1e5f0f0},
  {32'h425e7e14, 32'h439ad60b, 32'h43959996},
  {32'hc40098a2, 32'hc38cc42a, 32'h432cc3ea},
  {32'h429e8b0e, 32'hc3b60759, 32'hc1b7c6d4},
  {32'h43f4ed20, 32'h422441b1, 32'h421b67bc},
  {32'hc2f6510d, 32'hc31df7f3, 32'h42ca7c57},
  {32'hc264adaa, 32'h436f5e23, 32'hc3914aa3},
  {32'hc2272ae5, 32'h42999641, 32'hc12a4768},
  {32'hc289ea5c, 32'hc2448056, 32'hc2a9bb78},
  {32'hc15b2ae0, 32'hc3f64725, 32'hc32f7597},
  {32'h446131d1, 32'h439d3f18, 32'hc38538df},
  {32'h4232bffd, 32'hc4181ed1, 32'hc306b7ee},
  {32'hc2ac7da0, 32'h4383db51, 32'hc32966aa},
  {32'h4380e0eb, 32'h444370a8, 32'h42f1b62a},
  {32'hc3beb5db, 32'hc3dc7fe4, 32'h43acf184},
  {32'hc31d1fac, 32'hc3e37545, 32'h42beceb4},
  {32'h43b5a832, 32'h434ea45a, 32'h4439aab7},
  {32'hc21dbb7f, 32'hc2f2f24f, 32'hc35e2b88},
  {32'hc438b7b3, 32'h43226bda, 32'hc1bf95e0},
  {32'h426e6065, 32'h4411d50d, 32'h4397255b},
  {32'hc2c25a9a, 32'hc3b9cbfc, 32'hc32381ac},
  {32'hc1f3a39a, 32'h42a57bc5, 32'h43a9a374},
  {32'h4325c131, 32'hc3ca49ef, 32'h43d514ce},
  {32'hc41f2448, 32'h433e28f8, 32'h4032c7aa},
  {32'hc21acd62, 32'hc33cff01, 32'hc2dbcfac},
  {32'h4234e86c, 32'hc2fc8fb7, 32'hc2b83745},
  {32'hc3e90c00, 32'hc18f94d6, 32'h4394368a},
  {32'h439f95cc, 32'h42d447bd, 32'h434fb459},
  {32'hc2e82947, 32'h4322bb02, 32'hc379daff},
  {32'hc0e5e820, 32'h42b03765, 32'hc39dcfba},
  {32'h432a0f20, 32'hc3e515af, 32'h4381e814},
  {32'h42409d71, 32'hc36b0b3f, 32'h42a4a862},
  {32'hc32b2ffd, 32'hc30ade15, 32'h43502ac7},
  {32'hc32369f7, 32'h42b9a812, 32'hc3b00d57},
  {32'hc1e3225e, 32'hc29b3339, 32'hc2e5490f},
  {32'h431eb13c, 32'hc3fdaf4b, 32'h43c09cdf},
  {32'hc40538ec, 32'h43f80e78, 32'hc29c0047},
  {32'hc28ffa80, 32'h433befcd, 32'h431e537e},
  {32'h43775192, 32'h4382a2b9, 32'hc3609ce9},
  {32'h43f0b862, 32'hc26fbc47, 32'hc303ec04},
  {32'h434d473c, 32'h43258298, 32'hc34f8225},
  {32'h40fdcc3c, 32'h43281e99, 32'h431a20db},
  {32'hc3ef931e, 32'hc22cdf10, 32'h4236d4c3},
  {32'h44010519, 32'hc4534e20, 32'h4395f4de},
  {32'hc3a78ce2, 32'h4345d958, 32'hc38f07dd},
  {32'hc3dd5408, 32'h43808a52, 32'h43a80f9c},
  {32'h43ab8155, 32'h43329f6e, 32'h43e1e6d5},
  {32'hc29c2308, 32'hc3ca06de, 32'hc31b7658},
  {32'hc321248f, 32'hc2a25f38, 32'h42d6ea7c},
  {32'h42b147cc, 32'h427f24a6, 32'hc2ef3572},
  {32'hc31e2fe6, 32'hc2e7c459, 32'hc337238b},
  {32'hbce14400, 32'hc241d2f9, 32'hc17e00ab},
  {32'h4353af47, 32'h418cc252, 32'h43752b87},
  {32'h41d98806, 32'h433547ce, 32'hc39c8885},
  {32'h42e4261e, 32'h423766c0, 32'h42ad2a56},
  {32'h434c68f7, 32'h4326db6a, 32'h420cd839},
  {32'h438a9692, 32'h4323a535, 32'h43b38ce3},
  {32'hc29a0454, 32'hc33d0d27, 32'h41b1d6a7},
  {32'hc273fad8, 32'hc39bb78a, 32'hc3ef1f10},
  {32'hc23af58c, 32'hc38f5914, 32'h431eaf66},
  {32'hc3c1cebb, 32'h42bcd9c5, 32'hc28f531f},
  {32'h42862bc3, 32'hc34dc95f, 32'h42d44c9a},
  {32'hc3f02751, 32'h42f6b3c7, 32'hc355269e},
  {32'hc2f248b8, 32'hc3636331, 32'h43158e6e},
  {32'hc3258d70, 32'h4325eecd, 32'h43822c3c},
  {32'hc296e3fa, 32'hc2520687, 32'hc4024d7c},
  {32'hc2cf97a3, 32'h42baa5c6, 32'h428d9585},
  {32'h43a8cfcd, 32'h431ab9ae, 32'h4371cf01},
  {32'hc3380734, 32'hc3a98a8f, 32'hc30081d3},
  {32'hc3000e8f, 32'hc3a163b9, 32'hc2ddbbfd},
  {32'h42f9c5bd, 32'hc3df9d1b, 32'h43c472e0},
  {32'hc3f47a49, 32'h437f17e7, 32'hc23181cf},
  {32'h4367ad60, 32'h440a4a40, 32'hc31d766b},
  {32'h4381f62a, 32'h42ef563e, 32'h420fb168},
  {32'h418109d0, 32'hc3a58c0f, 32'h438e95e9},
  {32'hc32a7242, 32'h4319930d, 32'h43fa89c3},
  {32'hc10f20b0, 32'hc4084b12, 32'h438ace4c},
  {32'h42c6b954, 32'hc2a17136, 32'hc27637de},
  {32'hc35865b4, 32'hc3b9d9ff, 32'h4343fa33},
  {32'hc0787100, 32'hc306bfc1, 32'hc38eb75b},
  {32'hc3cf0d2a, 32'h42cdae50, 32'h438cfb7e},
  {32'h4367162a, 32'hc3adeaec, 32'hc23ca1e3},
  {32'hc2f598ef, 32'h42bf930f, 32'hc3a4261c},
  {32'h42996c43, 32'hc3724fb5, 32'h43403690},
  {32'hbf4e0bce, 32'h429531c0, 32'h42030be6},
  {32'h43aac494, 32'hc21ff7da, 32'h42192fb1},
  {32'h4367333b, 32'hc3d4f63d, 32'hc408fc1f},
  {32'hc3945009, 32'h411a2b35, 32'h439b3efa},
  {32'h4302dc57, 32'hc241821d, 32'h42ddf8ba},
  {32'h42ce67cb, 32'h430745e4, 32'hc3b27c33},
  {32'hc34073f3, 32'h424d8586, 32'hc1f323a2},
  {32'h4275e67c, 32'hc36b9111, 32'h432eaad4},
  {32'h43455351, 32'hc167cd9c, 32'hc327de5a},
  {32'hc130f9fc, 32'hc4072a2b, 32'hc3287392},
  {32'h42a3413e, 32'h4326d4ef, 32'h4398a31f},
  {32'hc3ab0456, 32'hc4047d42, 32'hc2387d51},
  {32'h43412c55, 32'h43de78e5, 32'h4300c262},
  {32'h43b2f00b, 32'hc3b0c728, 32'h42856168},
  {32'hc3251e9c, 32'h437d35f4, 32'h43650660},
  {32'h42b9c325, 32'h41daff03, 32'hc394b68a},
  {32'h411775b2, 32'h4303eb38, 32'h432c2e2f},
  {32'hc312000f, 32'hc2d3a10f, 32'h4295dfd5},
  {32'hc2c5ceb6, 32'hc3ded122, 32'hc2ea7932},
  {32'h41d4ffb1, 32'hc360925d, 32'hc2f2a203},
  {32'hc3dd1e0e, 32'h439c68ac, 32'h431c101b},
  {32'h3f9e29d8, 32'h434161e9, 32'hc37352cc},
  {32'h42e80b52, 32'hc2b44918, 32'hc3f69552},
  {32'hc418d1f2, 32'h4386b181, 32'h441ad015},
  {32'h432ccdb1, 32'hc3a79e37, 32'hc377e583},
  {32'h44165613, 32'h4309cee2, 32'hc36a183c},
  {32'hc1a9ada8, 32'hc34663e8, 32'h42ee722d},
  {32'h4379448a, 32'h43f36b9f, 32'hc2c35305},
  {32'hc35fc97e, 32'hc2d0e308, 32'h432f23b5},
  {32'h41019eac, 32'hc27f4bf1, 32'h42f3e2be},
  {32'hc3218ca1, 32'hc3d922ad, 32'hc39194d2},
  {32'hc3e8a25d, 32'h43f98ca9, 32'hc36cc4ff},
  {32'hc310699b, 32'h43c3e56a, 32'h440ca99c},
  {32'hc3fb60ad, 32'h422c5788, 32'h420263c9},
  {32'h43633456, 32'hc341b2fa, 32'hc3d35463},
  {32'hc4421b21, 32'h438b8aa2, 32'h43699e99},
  {32'hc26aa1c6, 32'hc414545e, 32'hc3b030fb},
  {32'h430210c6, 32'hc154b2a6, 32'hc2a6cf6e},
  {32'hc2ccca09, 32'hc20e5346, 32'h439b45e2},
  {32'h433d4d57, 32'hc3b906c2, 32'h43ea2551},
  {32'hc3d30006, 32'h43284457, 32'hc31ac804},
  {32'hc3662cd4, 32'h430b105a, 32'hc288c078},
  {32'h435c4319, 32'h42d281a4, 32'h40244198},
  {32'h42c75a2c, 32'h42c852a8, 32'hc3b4876c},
  {32'hc28587bb, 32'hc32d867f, 32'hc30a5cfa},
  {32'h4339aa49, 32'hc391edc5, 32'h4393650a},
  {32'h430ab574, 32'hc38dd557, 32'hc34dab82},
  {32'hc3b3381c, 32'h43ac7783, 32'h421588ca},
  {32'hc381574a, 32'h437279d7, 32'h43b1f303},
  {32'h43880c6f, 32'hc1883ea2, 32'hc328c670},
  {32'h425cf374, 32'hc2f93ff8, 32'h43120789},
  {32'h408b51a9, 32'h4257797b, 32'h43011492},
  {32'hc30fcdb2, 32'hc282e50f, 32'hc3fa5eb6},
  {32'hc3fbdb0c, 32'hc20b894f, 32'h4361dbe8},
  {32'h428016bc, 32'hc382e708, 32'hc39f3861},
  {32'h43612b40, 32'hc1721929, 32'h419a38e2},
  {32'hc3fa5469, 32'h43830fcd, 32'hc3377c03},
  {32'hc322d534, 32'hc2bc71fa, 32'hc3a10c28},
  {32'hc372abb0, 32'hc2705ff3, 32'hc21f62d1},
  {32'hc3af5c66, 32'hc35e5499, 32'hc388fb5c},
  {32'hc38731d7, 32'hc31218d0, 32'h40dd6c81},
  {32'h43b90bdf, 32'hc373efbb, 32'h43e2f3bc},
  {32'h433aa7bc, 32'h432011ad, 32'hc3d07bc6},
  {32'hc397b6bb, 32'h4378392f, 32'hc3d7453b},
  {32'h430a9c29, 32'h43b94ee3, 32'hc36e26f0},
  {32'hc36dd7df, 32'h438d6c11, 32'h43c07bbb},
  {32'hc32b69f4, 32'hc3260327, 32'h42e47071},
  {32'h42689f06, 32'hc1d555f6, 32'h43cf1ad6},
  {32'hc382b3e1, 32'h43656a66, 32'h423718a1},
  {32'hc3064f84, 32'h42bd3617, 32'hc393b027},
  {32'h4312dc89, 32'h439dbeaf, 32'hc27b75ed},
  {32'hc3314226, 32'hc31c03c1, 32'hc3448969},
  {32'h423765fa, 32'h4338552c, 32'h42b72aba},
  {32'h43a1d392, 32'h4346da93, 32'hc0d7f0fa},
  {32'hc3e3ad5f, 32'hc19745a0, 32'hc2b6fa88},
  {32'h4136de10, 32'h42109c8a, 32'h4272b510},
  {32'h4319de7b, 32'h43d6728f, 32'hc3a574b2},
  {32'h43e15622, 32'h43c8f91e, 32'hc0eae278},
  {32'h42e2b6d0, 32'hc383d035, 32'hc15bd14a},
  {32'hc388f9db, 32'h439b0740, 32'h40178ff6},
  {32'hc35b2958, 32'h442be60e, 32'hc2d7c741},
  {32'hc383a2c7, 32'h415f410b, 32'hc2b799be},
  {32'h440ab657, 32'hc1cb9bb8, 32'h425e9284},
  {32'h42a29cc5, 32'hc258d263, 32'hc2b4cc9c},
  {32'hc42dde5c, 32'h431658b8, 32'h436e0a36},
  {32'hc21506bd, 32'hc37fcc8f, 32'hc3a7675f},
  {32'h43e4c93a, 32'h43537e29, 32'hc26a2bc5},
  {32'hc337a6be, 32'hc33bb69a, 32'h436abfe1},
  {32'h44069e3a, 32'h425a7cad, 32'hc35b2656},
  {32'hc43350fc, 32'h4257913d, 32'hc3f417da},
  {32'hc36f69c4, 32'hc2e3f03e, 32'hc346356c},
  {32'hc1f2f694, 32'h43e594f6, 32'hc2ea1c71},
  {32'hc3ab1d2d, 32'hc3fff3b5, 32'hc28ea488},
  {32'h43526086, 32'h43a945d1, 32'hc3b67061},
  {32'h43dd24e8, 32'h432dc62f, 32'h44024adc},
  {32'hc2b845a2, 32'hc34bd801, 32'hc3266810},
  {32'hc3824226, 32'h4411f68d, 32'h42ca5ba6},
  {32'h41ade560, 32'h41db5a6d, 32'hc39c6019},
  {32'hc2ebf411, 32'h4277c3ab, 32'hc33f7d2f},
  {32'h43b09532, 32'h434365c6, 32'h423d3e8b},
  {32'h4345d83c, 32'hc1a9fe4c, 32'hc12c1f6c},
  {32'hc2cc6e0e, 32'h41a79023, 32'h42960756},
  {32'h42c339b8, 32'h43d6c3e2, 32'h43d55c6c},
  {32'h41f07354, 32'h4260bb10, 32'hc327683a},
  {32'h4300a497, 32'h4324cd5c, 32'hc3bb2607},
  {32'h43bae4da, 32'h43489094, 32'hc3667ab7},
  {32'h43063b3f, 32'hc1feccf3, 32'hc3205c35},
  {32'hc3c204bc, 32'h42c638d8, 32'h43a85b7f},
  {32'hc1af487d, 32'hc2f7e526, 32'h41045d20},
  {32'h426c25aa, 32'h43204957, 32'hc3d614d0},
  {32'hc386e182, 32'hc30092c9, 32'h436f17fc},
  {32'h424e8b64, 32'h430cb56a, 32'h438ee913},
  {32'hc3cbd06c, 32'hc2ab64e7, 32'h43be930c},
  {32'hc3bb02f9, 32'h4398ac24, 32'hc32db79b},
  {32'hc4049eb6, 32'h42baf93b, 32'h42455665},
  {32'h43a8e9de, 32'h4327fe29, 32'h430da0e1},
  {32'h43959135, 32'h438b0d61, 32'hc3687766},
  {32'hc3db7f2a, 32'h430547dc, 32'h425118ed},
  {32'hc3387062, 32'hc3832c47, 32'hc24bb18e},
  {32'hc42f8565, 32'hc38dced6, 32'h439fd127},
  {32'hc30eab18, 32'hc3e719a8, 32'hc38f483d},
  {32'h439592ff, 32'hc30b0d9e, 32'h43d68b23},
  {32'h43cc5d9d, 32'h439d0d80, 32'hc2553a13},
  {32'hc33755c4, 32'h44305acd, 32'hc319e6b8},
  {32'h439ef70f, 32'hc186934a, 32'h43d27397},
  {32'hc3856f73, 32'hc290b3f5, 32'hc2c274f1},
  {32'h43890d6a, 32'hc306c7b8, 32'h42fee6b0},
  {32'h43af624e, 32'hc34a744f, 32'h4303beed},
  {32'hc22cb834, 32'h42bbc3a0, 32'hc396dbbd},
  {32'hc3883a67, 32'h40cd5c06, 32'h4386bd3c},
  {32'hc32a1412, 32'hc39ca837, 32'hc3ecc1c4},
  {32'hc137b33e, 32'h44014510, 32'hc3d3f641},
  {32'h43e145c0, 32'h439fd080, 32'h432603d9},
  {32'h437b542c, 32'hbf9f53e0, 32'h43113834},
  {32'hc3e7421e, 32'h438e93f3, 32'hc36ddcc2},
  {32'h434e0f3b, 32'hc1f0b49a, 32'hc36f23c0},
  {32'hc36141b8, 32'hc3f0071f, 32'h410afb61},
  {32'hc3411168, 32'h42d096b2, 32'hc3937a38},
  {32'hc31846ca, 32'h4325d459, 32'h41a5c9bd},
  {32'h4323937d, 32'h432480a9, 32'hc423f6f3},
  {32'h4313d442, 32'h4042e3b0, 32'hc3a72e1a},
  {32'hc2f53045, 32'h438bc9d2, 32'h440dedc6},
  {32'h42dcac4c, 32'hc3ea8fde, 32'h42e065ef},
  {32'hc3b08e1f, 32'hc3a3ac58, 32'hc3101604},
  {32'hc433883a, 32'h43a7e004, 32'hc390daa2},
  {32'h4388ca8f, 32'h439c64ef, 32'hc3ddd54a},
  {32'hc34bb3ca, 32'hc368ebd3, 32'hc34a31d2},
  {32'h433cc412, 32'hc4027a10, 32'hc29dd108},
  {32'h433c05a6, 32'h40114a70, 32'hc34e9e05},
  {32'h3ffd28b8, 32'h43047460, 32'hc32b0e0e},
  {32'hc335a24c, 32'hc3a4f187, 32'hc2a89943},
  {32'hc3026a60, 32'h43a718f4, 32'h43a45511},
  {32'hc33fd60e, 32'h43042e7a, 32'hc3abffb1},
  {32'h431e4e33, 32'hc28514f6, 32'h4294761c},
  {32'h428efa83, 32'h42ec1f8f, 32'hc3963c82},
  {32'hc33216c2, 32'hc23e8b86, 32'h43570df0},
  {32'h42918b88, 32'h43664ada, 32'h4323d7ce},
  {32'hc36a3acb, 32'h42f5b307, 32'hc3b4c782},
  {32'h422fb645, 32'hc3b034df, 32'h43acd5bf},
  {32'h42eb4c61, 32'hc24b11b4, 32'hc2ceda30},
  {32'h4354a6de, 32'h42bfbfdd, 32'hc3714b38},
  {32'hc3903c6e, 32'hc3695472, 32'h439f8276},
  {32'hc1fc3580, 32'h4312b16b, 32'hc2e13f20},
  {32'hc1c1f9b1, 32'hc2fc91af, 32'hc35ead9f},
  {32'hc1409812, 32'h439d86dd, 32'hc34b9458},
  {32'hc2e12bb5, 32'h4312ff8a, 32'hc426c628},
  {32'hc2dfc552, 32'h42cc1407, 32'hc2e9b49c},
  {32'h42b1689d, 32'h42ca952c, 32'hc30dda13},
  {32'h4416e6e9, 32'h4273b1ef, 32'h43a9e66f},
  {32'h43ae4634, 32'hc2743ad6, 32'hc3e5c11d},
  {32'hc38d548a, 32'hc2082e19, 32'hc3648b94},
  {32'h42d1cab4, 32'hc39207bc, 32'h430ecd65},
  {32'h4339bdac, 32'h43294e59, 32'h43dc3bb1},
  {32'hc40032fe, 32'hc15cb940, 32'h43fdd234},
  {32'hc2ff50ae, 32'hc32037e9, 32'hc3362ac4},
  {32'hc2037be6, 32'hc3f5de1e, 32'h436d0998},
  {32'h42eff4cb, 32'hc3627a04, 32'h42312502},
  {32'hc40f9dcc, 32'h43e3d4c6, 32'h43ac766c},
  {32'hc38015e3, 32'h42ca433f, 32'hc37c35db},
  {32'h42b60519, 32'hc32bc868, 32'h42d52d86},
  {32'h4314c66b, 32'h3e638fd0, 32'hc263c335},
  {32'h43a2e1ca, 32'hc326edce, 32'h431e218d},
  {32'hc2448012, 32'h4394649f, 32'hc37e7078},
  {32'hc29d5621, 32'hc24f74c9, 32'h431cb975},
  {32'h435fd401, 32'hc30b2ddc, 32'hc1a9f020},
  {32'hc3ce8a8e, 32'h43c0b18a, 32'h439cf58e},
  {32'h43b2fa9b, 32'h43c95cf9, 32'h442eb714},
  {32'hc21dbb45, 32'h433defde, 32'hc38e1fdf},
  {32'h431f1080, 32'h43856969, 32'hc2a3397a},
  {32'hc37eb5e8, 32'h428542cf, 32'hc4060d2d},
  {32'h43e4eb24, 32'hc3ac5a95, 32'h42e578fc},
  {32'hc362a541, 32'h428526a0, 32'h42693c26},
  {32'h42854fe8, 32'hc30b159e, 32'hc416c772},
  {32'h436f5193, 32'h42b7cbeb, 32'hc31eb46d},
  {32'hc3bb48dd, 32'hc40271e5, 32'hc187f147},
  {32'hc3efb63d, 32'h42a47f73, 32'hc1bf36fa},
  {32'h43a28f66, 32'hc3d8b3a2, 32'h4338b471},
  {32'hc318a042, 32'hc34255ba, 32'h433b6f04},
  {32'h43fe1509, 32'hc2435e48, 32'h4348c8bc},
  {32'h441dcce8, 32'h437568b4, 32'h433d9731},
  {32'h43cc997e, 32'hc311c804, 32'h440a8ec9},
  {32'h4289b250, 32'h43a015b3, 32'hc380b573},
  {32'h42c89534, 32'hc360d0b1, 32'hc2dceee2},
  {32'h425b3706, 32'h40cb483a, 32'h422900a3},
  {32'hc40e4b5f, 32'h43b9b399, 32'h43e5bd2f},
  {32'h435afa31, 32'h4349073e, 32'hc2e62511},
  {32'h42d34a8a, 32'hc2c38867, 32'hc2116996},
  {32'h43429a6d, 32'h42af9190, 32'h427f0d30},
  {32'h43856a70, 32'hc3cdc356, 32'h43d45268},
  {32'h420f1639, 32'h436fab22, 32'hc3c1a4b4},
  {32'hc2048f96, 32'hc3887a75, 32'h4403817d},
  {32'hc29bee75, 32'h4211e5bc, 32'hc25c5e77},
  {32'hc20f8232, 32'hc245174a, 32'h4336e492},
  {32'h432b93d2, 32'hc2539bb8, 32'h43a1435c},
  {32'h437468af, 32'hc3795f1d, 32'hc4075d44},
  {32'hc3d8507c, 32'hc3825383, 32'h439fba5a},
  {32'h42b799ad, 32'h43d93efe, 32'h42bb62be},
  {32'h429f3252, 32'h4405bbd9, 32'hc4661757},
  {32'hc3959f2d, 32'h43a6ce21, 32'hc345f727},
  {32'hc36ddec9, 32'h433c71da, 32'hc3e3991a},
  {32'h42287d50, 32'h43089fda, 32'h41329b58},
  {32'h442bbb79, 32'h41e99cee, 32'hc32f0b4e},
  {32'h419c4e34, 32'h438071ee, 32'h4337cacd},
  {32'h43c6ca18, 32'hc2ef6a42, 32'h4366dc01},
  {32'h4195c9b0, 32'hc3aed2b3, 32'h433b2ff5},
  {32'hc30efb51, 32'h426b043e, 32'h43dab9ce},
  {32'h440a8b34, 32'hc1cce505, 32'hc4119023},
  {32'hc36cf843, 32'hc420ee4a, 32'hc3309e36},
  {32'h43d65b76, 32'hc419910b, 32'h440a6a20},
  {32'h43b12c77, 32'hbf9b2620, 32'h441ce5fb},
  {32'hc2fb2ce1, 32'h41c5359d, 32'h4338948d},
  {32'h43e9912b, 32'hc23f72e9, 32'h43d2436c},
  {32'h429a43c4, 32'h4347c6d9, 32'hc1b299e5},
  {32'h4313e3dd, 32'h429a9e03, 32'hc20c1ecc},
  {32'hc34b2590, 32'hc390d956, 32'hc368995c},
  {32'h42645b7c, 32'h43b99824, 32'h432d83a4},
  {32'hc3cbdb43, 32'h43a0284d, 32'hc36dee60},
  {32'hc2ceddc8, 32'hc288cdd5, 32'h4381854e},
  {32'hc348ad94, 32'h4339dff5, 32'hc335d57a},
  {32'hc3890fb8, 32'h43556154, 32'h43af059a},
  {32'h4372c7dc, 32'h43016991, 32'hc3231f80},
  {32'h4233d41c, 32'hc3233eea, 32'hc30600bc},
  {32'h421d7f14, 32'hc377227f, 32'h42dfc2ef},
  {32'hc3887dc9, 32'h434986d1, 32'hc3ba5b6c},
  {32'h437514a7, 32'h40f53dcb, 32'hc3841e08},
  {32'hc1b3726c, 32'hc3321290, 32'hc2610155},
  {32'hc3629ffe, 32'hc3840631, 32'hc3700a2b},
  {32'h4387b032, 32'hc36afd9a, 32'h43b7d6a5},
  {32'h437f203d, 32'hc1bc9b4d, 32'hc385ba3a},
  {32'h413804c0, 32'hc3a9b54a, 32'hc228b612},
  {32'h443b199b, 32'h433a97c2, 32'hc21557bd},
  {32'h42d25b15, 32'hc16c374a, 32'h42ef153a},
  {32'hc3243e47, 32'hc20c3e02, 32'h4284053e},
  {32'h42d6f828, 32'h4410ca6c, 32'h4355c600},
  {32'hc39ab0c8, 32'hc416ae1e, 32'hc344ca0a},
  {32'hc303fe34, 32'h43a04a7a, 32'hc2f10dc2},
  {32'h4390762d, 32'hc3a62377, 32'h42b0bd5b},
  {32'hc2709e13, 32'hc342a5a7, 32'hc33cd1c4},
  {32'h43cc3fd4, 32'h4338d77a, 32'h43ed3588},
  {32'h43be9e52, 32'hc3e7d415, 32'h43935689},
  {32'h439fc4a7, 32'hc1927a1b, 32'h4217fbea},
  {32'h416fba6e, 32'hc1a99b21, 32'hc3022945},
  {32'h432ab2a2, 32'hc1cc645b, 32'hc20a7711},
  {32'hc3c76946, 32'h4271c4ad, 32'h43a27ddf},
  {32'hc384e37c, 32'hc169c117, 32'h432b88a6},
  {32'h4368320f, 32'hc26843f8, 32'hc2f56289},
  {32'h4302b164, 32'h43f12128, 32'hc361fbf3},
  {32'h43987926, 32'hc2aafee5, 32'h4235b448},
  {32'hc2926a07, 32'hc1abe6d1, 32'h41020e96},
  {32'hc1ff3cd6, 32'hc416ad39, 32'h4391a622},
  {32'hc3533336, 32'h4227af74, 32'hc3599d8d},
  {32'h43edf108, 32'h42e154a9, 32'hc30b6282},
  {32'h438053bf, 32'h427398f5, 32'hc2ab58de},
  {32'hc381fc9a, 32'h420f7e2e, 32'hc36e37b7},
  {32'h41b65bb0, 32'hc16567fc, 32'h4264c8df},
  {32'hc377577a, 32'h4384bb66, 32'h43ab7cc1},
  {32'hc4034ded, 32'h408afcb5, 32'h42a46240},
  {32'h42d13f05, 32'h43d1bf4b, 32'hc460a9c9},
  {32'h42ad3df4, 32'h4403d869, 32'h4300ef8a},
  {32'h40c9074c, 32'hc344834e, 32'hc390a52c},
  {32'h438d5b47, 32'h4328f555, 32'h43654c92},
  {32'h42874edc, 32'hc2b39c35, 32'hc28b2482},
  {32'hc3d231e7, 32'hc229a27e, 32'hc2fc4153},
  {32'hc37d70a3, 32'hc3135f76, 32'h43fd2588},
  {32'h42ec4c5c, 32'h426fe066, 32'h42c324df},
  {32'h433e4b45, 32'hc3288a1d, 32'hc2d1f4ef},
  {32'hc067b17a, 32'h41745826, 32'hc3bc8cc9},
  {32'h439f1b38, 32'hc17528c3, 32'hc1a5bbdc},
  {32'h43663310, 32'hc39c2c55, 32'h437a717a},
  {32'h431a3c62, 32'hc3935a01, 32'h41d3bfc7},
  {32'h423a44ec, 32'h418e7dda, 32'hc36a161a},
  {32'hc39c0b3b, 32'h433769e2, 32'h441ad6ac},
  {32'hc31de878, 32'h41cdfba6, 32'hc2a66e86},
  {32'h42d4668d, 32'hc37200ea, 32'h4396363b},
  {32'hc2fe6c82, 32'hc3a12595, 32'h43afff43},
  {32'hc2a24991, 32'h42d48a94, 32'h4243cf12},
  {32'hc37b6435, 32'hc40782fa, 32'h41e62b9e},
  {32'h43b05596, 32'h435d28c4, 32'hc393b08d},
  {32'hc0fa8cd0, 32'hc3171e08, 32'hc3d98835},
  {32'hc40c164f, 32'h423ca2e2, 32'hc3f9c6b4},
  {32'h4289c8b4, 32'hc3851f11, 32'hc415f0c3},
  {32'hc3e64281, 32'hc24bc01f, 32'hc35defad},
  {32'h42d16e9b, 32'h4308283e, 32'h438f2896},
  {32'hc41b1d81, 32'hc3cd7c70, 32'h439fddd6},
  {32'h431fdf68, 32'h4354945d, 32'h4397105a},
  {32'hc3cf3fe6, 32'h4399f322, 32'hc311cc47},
  {32'hc3dc8d0d, 32'h4133d07b, 32'h43eec71c},
  {32'h43b64d6d, 32'hc0f33a64, 32'h433241a9},
  {32'h42dbe1d2, 32'h419a8b92, 32'h42d41859},
  {32'h4380f152, 32'hc2d07e08, 32'hc11ebf6a},
  {32'h4415277d, 32'hc32fc5c2, 32'h438475f6},
  {32'hc3d547a4, 32'hc29cfc3e, 32'hc1a39e92},
  {32'hc32f1aac, 32'hc317083c, 32'h43361bcd},
  {32'hc31ee5f0, 32'hc3cd80bd, 32'h431af23a},
  {32'h428ac518, 32'h4216eb9d, 32'hc35d0466},
  {32'hc3b1d155, 32'hc3394b7f, 32'hc25d93dc},
  {32'h42532874, 32'hc38e54b6, 32'hc312126b},
  {32'h432971ed, 32'hc2cadc18, 32'hc30a5018},
  {32'h40e612d4, 32'h438e5839, 32'hc26532f4},
  {32'hc37f508b, 32'hc2a80849, 32'h436a31e8},
  {32'hc35806fe, 32'hc38e6511, 32'h3ed2c243},
  {32'hc333ae4c, 32'h439e7ac0, 32'h4353304e},
  {32'h42b3d807, 32'hc3107487, 32'hc34e01eb},
  {32'hc3021404, 32'hc35c3576, 32'h438a5e1c},
  {32'hc2a5f0d6, 32'h433c8a16, 32'hc3429900},
  {32'h438966c3, 32'hc30ef9cc, 32'h42ee527f},
  {32'hc31bdbc6, 32'hc37d25d9, 32'hc3195629},
  {32'hc2238917, 32'hc3579880, 32'hc40e943a},
  {32'h43825283, 32'h425a3800, 32'hc3dcd5cb},
  {32'h410d2704, 32'h4385eca2, 32'h440e0aeb},
  {32'h43c0170d, 32'h428cf1e7, 32'hc31d486e},
  {32'hc26e75e0, 32'h434f8581, 32'h441700f3},
  {32'h43470398, 32'h440cb2a0, 32'h42dda4e0},
  {32'hc3152611, 32'hc3957b79, 32'hc3f20fa9},
  {32'hc3417ad6, 32'hc1275588, 32'h432e3434},
  {32'hc34cb9d4, 32'h4165e5c3, 32'hc374f5cc},
  {32'h4380f090, 32'hc38366f8, 32'h43d5a09d},
  {32'h43acade2, 32'hc33203c2, 32'h43e7c7af},
  {32'hc385403b, 32'h42aed8a0, 32'h41849bce},
  {32'hc1a6f9d4, 32'h434e2b38, 32'hc341275b},
  {32'h44097f71, 32'h4412c5c6, 32'hc2d3b1a3},
  {32'hc30bc73f, 32'h43cf0a4a, 32'hc36fdf9f},
  {32'hc3302934, 32'hc3c84bcf, 32'hc25e2f9b},
  {32'h438f3b9b, 32'hc35a772f, 32'h433616a5},
  {32'h43ccdab0, 32'hc331f8f5, 32'h429f3462},
  {32'h43322004, 32'h421a444c, 32'h42a3fd1e},
  {32'hc1a56c20, 32'hc30f9e5c, 32'hc279b2aa},
  {32'hc39f0fa3, 32'hc21febd7, 32'hc386f56b},
  {32'hc22c21b4, 32'hc364412b, 32'h441857f1},
  {32'h43ac175d, 32'hc36232b7, 32'hc32c6cf5},
  {32'h43a8a3fb, 32'h43671ada, 32'hc41aaa45},
  {32'hc3a6a4ce, 32'hc30dbb3b, 32'hc2df2dc8},
  {32'h4347f1b3, 32'h427c7e4c, 32'hc411817e},
  {32'hc3bec577, 32'hc373cefc, 32'h439087c8},
  {32'hc390c1f9, 32'h43404a94, 32'hc2c24dbc},
  {32'h43a3d24a, 32'hc39737b0, 32'h4389c9a2},
  {32'hc332106d, 32'hc2ecf76a, 32'h43035a78},
  {32'h4173eeac, 32'h43d0e0b2, 32'h440ff1c0},
  {32'hc3615fb8, 32'hc38972f8, 32'h43b0d203},
  {32'h42648e82, 32'hc38f1113, 32'h439dfe37},
  {32'hc44dbafe, 32'hc349cb2e, 32'h4362d147},
  {32'hc3465652, 32'h435bb52a, 32'h43119dd2},
  {32'hc3c8199c, 32'hc2db5e61, 32'hc303fcf8},
  {32'h421da339, 32'hc3cc61d0, 32'h4382fee2},
  {32'h4298162e, 32'hc34acbef, 32'h43cafe56},
  {32'hc3856e40, 32'h43874b5c, 32'hc348dcc2},
  {32'hc3932bd2, 32'h431769d0, 32'hc30630a1},
  {32'h43008c5d, 32'hc295a8c3, 32'hc36e9add},
  {32'h430997dd, 32'hc402c0b7, 32'hc353400e},
  {32'hc1f6b47c, 32'hc3ba5480, 32'hc335cfc3},
  {32'h437c8321, 32'hc21c5d36, 32'h41c3603b},
  {32'hc3e19b51, 32'h438afc3b, 32'hc295cebd},
  {32'h436be8bb, 32'h435d26b3, 32'h4338dd47},
  {32'h43709c9b, 32'hc37d31ed, 32'hc3a6584a},
  {32'h43ae3ea3, 32'h43b13a60, 32'h43a0f49d},
  {32'hc3a19e4c, 32'h428521d9, 32'h437419ad},
  {32'h4350453c, 32'h432b121c, 32'hc3c9f1f8},
  {32'hc32196c2, 32'hc3731b25, 32'hc1abf46b},
  {32'h4291f1ee, 32'hc24d815d, 32'hc3605669},
  {32'h43b36c70, 32'h43cfc3c7, 32'h42a08a48},
  {32'h4359f12b, 32'hc384c96c, 32'hc27869e2},
  {32'hc3903d99, 32'h438de378, 32'hc3fad481},
  {32'h4280db10, 32'hc3e9aa2f, 32'hc3d02e8e},
  {32'hc3a7f787, 32'h4391fc39, 32'h4262ea7e},
  {32'hc34e8284, 32'hc366f32a, 32'h41c0a200},
  {32'h42ae38f4, 32'h4305d456, 32'hc30d9d0a},
  {32'h43a5f9db, 32'h418238fe, 32'hc399a2a4},
  {32'h43a47ef5, 32'hc33bbf0a, 32'hc2d3044b},
  {32'h43ee5040, 32'h42f47948, 32'hc2a98d9b},
  {32'h43c9e2d7, 32'h41f63e85, 32'hc30764a4},
  {32'h4395e7c1, 32'hc42258b2, 32'h438ad17c},
  {32'h433c20be, 32'h43122786, 32'hc36ac1db},
  {32'hc3883d80, 32'hc171e73f, 32'hc3990c13},
  {32'h43f8f915, 32'h434db1d2, 32'h438ebeea},
  {32'h42c589c7, 32'hc38c048d, 32'h44185977},
  {32'h420f8b0e, 32'h43575e5f, 32'h42177c2b},
  {32'h42e9f541, 32'hc307770f, 32'h4319be83},
  {32'h42f13c81, 32'hc348c046, 32'hc39bc3b0},
  {32'h423af87c, 32'hc2bc0c3f, 32'hc28bd8e1},
  {32'hc2af8014, 32'h43339bda, 32'h4408b0d6},
  {32'h434de5fe, 32'h435c1bbd, 32'hc31d2027},
  {32'hc37987b5, 32'h41976e3e, 32'hc3f800c7},
  {32'hc30acb84, 32'h41a0adbb, 32'h4239512b},
  {32'h436343bb, 32'hc22ef0e2, 32'h42dc55eb},
  {32'hc2589748, 32'h41b03c0a, 32'h436808cc},
  {32'h402b8160, 32'hc2db7300, 32'hc31df7f0},
  {32'h42753179, 32'hc2b08f95, 32'h42958ad3},
  {32'hc4424da6, 32'hc3815600, 32'hc3ca1177},
  {32'hc3b53f71, 32'h40b463f4, 32'hc3ef9110},
  {32'hc33938ce, 32'hc319f3ee, 32'hc1f6e328},
  {32'hc3b0ca57, 32'hc318ceef, 32'hc2b4f154},
  {32'hc344880b, 32'h43a58500, 32'hc3c4fd7b},
  {32'h442e5b32, 32'hc2e14c91, 32'h4293d8c0},
  {32'h43b3daf8, 32'h42f82f80, 32'hc363222c},
  {32'h436cc086, 32'hc2c8ebbb, 32'h43fd1961},
  {32'h4346f300, 32'hc36bdb91, 32'hc3b49ce3},
  {32'hc33452fc, 32'h42266acf, 32'h4390e5a3},
  {32'hc0bb413a, 32'hc39a7d43, 32'hc2688cd4},
  {32'h42a7499a, 32'hc2de6538, 32'hc3a1921e},
  {32'hc2b8b43e, 32'h439384de, 32'h3ea92b00},
  {32'hc3bd7e24, 32'h424571da, 32'hc28d3d77},
  {32'hc40ab6b4, 32'h43abf0db, 32'h41e86573},
  {32'hc3eae0c3, 32'hc30cd4d1, 32'h4329da5f},
  {32'hc2d854cd, 32'hc2af3f84, 32'hc2c1b732},
  {32'hc3125372, 32'hc3680f9e, 32'hc2b08ccf},
  {32'h435e3faf, 32'hc31c8b03, 32'hc3f5a563},
  {32'hc3724868, 32'hc2ff3699, 32'h440253c4},
  {32'hc404a022, 32'h4178dbd0, 32'h420b5f68},
  {32'hc38f64ad, 32'h42ce375d, 32'hc2997fdd},
  {32'h436457dd, 32'hc30a8f8a, 32'hc3942108},
  {32'hc199ca20, 32'h43b272f3, 32'h438d41a0},
  {32'hc1624784, 32'h42326e45, 32'hc2eacfdb},
  {32'hc319b31b, 32'h430d0525, 32'h43318986},
  {32'h439d7e34, 32'h436f26d9, 32'hc2bbdecb},
  {32'hc39b338a, 32'hc2c9c8a0, 32'h42da04a5},
  {32'h438c9ccf, 32'hc3857c80, 32'hc4357fb8},
  {32'hc30b9f74, 32'hc36ff197, 32'hc31752cf},
  {32'h43fff37c, 32'hc341bcce, 32'h43e434c0},
  {32'hc3befedc, 32'hc37234e0, 32'h43f7f91b},
  {32'hc0fcc410, 32'h430f90a5, 32'hc41d217a},
  {32'hc2d24514, 32'h43ed234d, 32'h43a0b7dc},
  {32'hc1d938fc, 32'hc40a7873, 32'hc1eeb57d},
  {32'hc26fb572, 32'h426556f3, 32'h42985c6a},
  {32'hc2a6f216, 32'hc325a415, 32'hc29976d4},
  {32'hc40a2176, 32'hc04301d4, 32'h4017b834},
  {32'h42905aed, 32'h4286add2, 32'h43d5f88f},
  {32'hc22dbb75, 32'h4366a2cd, 32'hc2c93723},
  {32'h43ac1526, 32'hc241d58d, 32'h425573f5},
  {32'hc37c4f04, 32'h43e524d3, 32'hc2857fed},
  {32'h4344e0bc, 32'h43cf40b5, 32'hc34dd618},
  {32'hc2f1c013, 32'hc360361d, 32'hc399b971},
  {32'hc2ad0c6d, 32'hc32ed6a7, 32'h3ffd9940},
  {32'hc2aa7e70, 32'hc30b43e8, 32'h41a5d9d6},
  {32'h421ca02a, 32'hc33d4522, 32'h43f62fc9},
  {32'h43a1ff9f, 32'h43430548, 32'hc4003b33},
  {32'h42a47001, 32'hc38066bd, 32'hc2a031d2},
  {32'h4251703d, 32'h41910a8a, 32'hc32b6385},
  {32'h42449224, 32'h43716218, 32'hc242c9f4},
  {32'h42c350fe, 32'hc404d345, 32'h43d05e0f},
  {32'hc2a448ef, 32'hc39a8679, 32'hc3b96c16},
  {32'h4251a163, 32'h4368891d, 32'hc2cdf7be},
  {32'hc3e69aec, 32'hc362656e, 32'h43207cda},
  {32'hc36ec4bc, 32'hc376a435, 32'h421252e2},
  {32'h43339a76, 32'hc3951b2d, 32'h431ec1d1},
  {32'hc24d0759, 32'h42af00bf, 32'hc2520322},
  {32'h4317987a, 32'hc399290d, 32'hc29e406d},
  {32'h44458062, 32'h43a468ed, 32'hc31697a3},
  {32'hc292ae5e, 32'hc26d9ea3, 32'hc3a00098},
  {32'hc3770eba, 32'hc29f3c9d, 32'h434c21f9},
  {32'h437d7c24, 32'hc291e346, 32'hc2d741b7},
  {32'hc33042ae, 32'h40c93288, 32'h43dd9625},
  {32'hc39f0d70, 32'h4305fc62, 32'hc337d6f3},
  {32'hc0e9b950, 32'h436782bc, 32'hc3a0cec6},
  {32'hc3864118, 32'h43bd1bf9, 32'hc3a88e7f},
  {32'hc3016cd7, 32'h434b1a16, 32'h439ddd09},
  {32'h43c861de, 32'h442c7406, 32'hc2a5e0f6},
  {32'h4212005c, 32'hc44bf1b1, 32'h42f9dc11},
  {32'hc349e7aa, 32'hc354850d, 32'h439bd71a},
  {32'hc1fb98ac, 32'h43a43350, 32'h433f4dc9},
  {32'hc3d57ebf, 32'h434fb8d7, 32'hc33362fb},
  {32'h419b5353, 32'h4232db8f, 32'hc36d59e0},
  {32'hc26a2644, 32'hc231b89a, 32'hc3c7e919},
  {32'h430b4588, 32'h437ba854, 32'h4294548f},
  {32'hc2d9eb42, 32'h4284c1e5, 32'hc3ded09b},
  {32'hc2ac720b, 32'h42f4e5cd, 32'hc2f1d5be},
  {32'hc3156201, 32'hc39cc956, 32'hc2051700},
  {32'h43019588, 32'h43839c7a, 32'h4214c87c},
  {32'h438c8718, 32'h4376301d, 32'h422311ca},
  {32'hc371647b, 32'hc3e169dd, 32'hc440d739},
  {32'hc38f1586, 32'hc348e9e6, 32'hc335d738},
  {32'h4185b2e3, 32'hc2db776a, 32'hc39c09ff},
  {32'hc29b0452, 32'h4341391f, 32'hc2184440},
  {32'h42820cbc, 32'hc30dc559, 32'hc40f9be1},
  {32'hc2faeb70, 32'hc373c277, 32'h436a28e4},
  {32'hc320156c, 32'h43def79a, 32'hc3d0f5fc},
  {32'hc37004a1, 32'h42d11366, 32'h43d52a52},
  {32'h43a126d8, 32'h437fc68b, 32'h41fcab5d},
  {32'h428bf417, 32'h4299cba0, 32'h428028d0},
  {32'h42340af1, 32'h421f4f27, 32'hc3b88895},
  {32'hc285c03e, 32'hc2ed2418, 32'h443285cc},
  {32'hc376591f, 32'h43948f7b, 32'hc2b216c0},
  {32'hc3343d1d, 32'hc20ff3b2, 32'h4199ebc5},
  {32'hc2c867aa, 32'h42d42209, 32'hc2e2bebe},
  {32'hc3d1d8e8, 32'h4223b217, 32'hc355a93c},
  {32'hc2de3c67, 32'hc3c5b608, 32'hc1b2beab},
  {32'hc2605ec2, 32'h43b22634, 32'h43194f98},
  {32'hc38d324f, 32'h430b2012, 32'h414dfbc8},
  {32'h4105b033, 32'hc1381819, 32'h4269d5b9},
  {32'hc337b5ac, 32'h44115447, 32'h436b9ede},
  {32'h430df4d6, 32'h4237616d, 32'h4286de6a},
  {32'h438a8ade, 32'h42c12b12, 32'h426979f0},
  {32'hc3888d80, 32'h43667f51, 32'hc246f00a},
  {32'hc3814343, 32'hc418d32b, 32'hc02d0227},
  {32'hc33f24de, 32'h439eef72, 32'hc35b3ff7},
  {32'h438041b6, 32'h420c83c8, 32'h4268040e},
  {32'hc3fe4e8c, 32'hc2be4cca, 32'h42da66ce},
  {32'hc392690f, 32'hc318b199, 32'hc32e69c5},
  {32'h42876dd8, 32'h43f4bf6a, 32'h43619b5f},
  {32'hc0d3cb08, 32'h43db674d, 32'h442d884a},
  {32'h42118117, 32'h43a60970, 32'hc324b78f},
  {32'h43b27384, 32'h432df313, 32'hc3d02400},
  {32'hc3860a06, 32'h42f781c0, 32'hc39d858a},
  {32'hc3c5df80, 32'hc29202f9, 32'hc2063af1},
  {32'h41f40a30, 32'h4198a058, 32'h43a53372},
  {32'hc3c6a674, 32'hc299a03d, 32'hc3423f58},
  {32'hc3b50310, 32'hc31915ab, 32'hc2859a8e},
  {32'h44372bdd, 32'h42aa441e, 32'h3fd74a66},
  {32'hc3088fbd, 32'h43f8d6e0, 32'hc3d3a520},
  {32'h423b66c4, 32'h43382420, 32'hc2fcece0},
  {32'h42693626, 32'h437b0974, 32'hc3237c45},
  {32'hc2fa7479, 32'hc26366ff, 32'hc33594b3},
  {32'h427c18ed, 32'hc2afaa7e, 32'hc3380eb7},
  {32'hc3b86826, 32'h4333a1b9, 32'h42da9678},
  {32'hc295330a, 32'hc30eb2df, 32'h4296ac7e},
  {32'h426e3dc1, 32'hc381a46f, 32'h43af483c},
  {32'h43acff2b, 32'h43a25f50, 32'h42c30eef},
  {32'hc3f95da6, 32'h43738a7f, 32'h43f1037e},
  {32'h42b88ef2, 32'hc23f525f, 32'h4329317d},
  {32'hc38d1674, 32'h437101a2, 32'h43835a12},
  {32'h41b01807, 32'h441a549f, 32'h4425e74a},
  {32'h422bf0bc, 32'hc2e0e379, 32'h43c9aa0d},
  {32'hc333661c, 32'hc3dbef9a, 32'hc3dfa8da},
  {32'hc328fac6, 32'h4414d4ae, 32'h40ef8c1c},
  {32'h42c22429, 32'hc3de6a1c, 32'hc3484ca8},
  {32'hc2d13461, 32'h42e74912, 32'h4336a16c},
  {32'h4392e62f, 32'h4364db6b, 32'hc2e956b0},
  {32'hc401bf1b, 32'hc133c06d, 32'h4390bf67},
  {32'h43981f6a, 32'hc31577e1, 32'h4337c49a},
  {32'hc3b889ea, 32'h436ec928, 32'hc34a6ede},
  {32'hc412913c, 32'h43132efb, 32'h43dc09f3},
  {32'h441be7e3, 32'h4388a91f, 32'h4429a106},
  {32'hc2fd9edf, 32'hc4042bcf, 32'hc2b885c8},
  {32'hc2d94324, 32'hc1b7c0c6, 32'hc2e7dbad},
  {32'h43c5d080, 32'h4395c79a, 32'h4458b8b2},
  {32'h4377d21a, 32'hc31fd798, 32'hc347f93e},
  {32'h43e575a4, 32'h4124ff36, 32'hc2aacab3},
  {32'h433062e6, 32'h428561eb, 32'h43f28a90},
  {32'h42b39c76, 32'h4354eb20, 32'h430f9bd5},
  {32'hc2aec879, 32'hc35c7822, 32'h43628bc5},
  {32'h42492e30, 32'h42e35ec7, 32'hc2fef555},
  {32'hc41b1de3, 32'h4370d272, 32'h4362acbb},
  {32'hc2529488, 32'hc3588088, 32'h4364f73f},
  {32'h435773be, 32'hc1b37c39, 32'hc3e5c37c},
  {32'h4295fa17, 32'h4386a631, 32'hc39dd3aa},
  {32'h43637852, 32'h43929eba, 32'h43e62580},
  {32'hc13d36d7, 32'h43054d7f, 32'hc35e8601},
  {32'h42915a5f, 32'hc3cc55e8, 32'h43447b75},
  {32'hc2f78e16, 32'h431e7cf9, 32'hc397ae7d},
  {32'h4186ef7b, 32'h4152ce12, 32'hc353c964},
  {32'h43699ee5, 32'h4290df74, 32'h429a6d31},
  {32'hc3bbb9c9, 32'h42fb8efe, 32'h437fc743},
  {32'hc2bd0766, 32'h43f22360, 32'hc2e26335},
  {32'hc245b5a4, 32'hc2d64e13, 32'hc39eea98},
  {32'hc42b203e, 32'h439c89fe, 32'hc39ba570},
  {32'h4406d234, 32'h3fcd8f6e, 32'hc30158f9},
  {32'hc3822db0, 32'hc3450d30, 32'hc3725f25},
  {32'hc38b344f, 32'h42ed9f67, 32'h433eaeb1},
  {32'h43b0d67f, 32'hc2b9c31b, 32'h437ddc00},
  {32'hc3e34284, 32'hc166d462, 32'h43c0e802},
  {32'hc2b0c5a0, 32'h43c7008e, 32'hc34b586e},
  {32'hc1ba8612, 32'h4261cfec, 32'hc3d2da4e},
  {32'hc4051da6, 32'hc3c18905, 32'hc360e52c},
  {32'hc398b9e3, 32'hc2a4228c, 32'hc3b5d9b4},
  {32'h42bac9fb, 32'hc1a8dfc8, 32'hc3a4c0cf},
  {32'h43033837, 32'hc33d8478, 32'hc2e178b5},
  {32'hc327a1ea, 32'hc3cdaab4, 32'hc3b361dc},
  {32'h413c7510, 32'hc3c6b896, 32'h43196d27},
  {32'h42c66e68, 32'hc19d5807, 32'hc30c88a6},
  {32'hc200a4dc, 32'hc3022d28, 32'h433b4325},
  {32'hc3fda9e1, 32'hc36525a6, 32'h4300322d},
  {32'h4206f945, 32'h4348bd56, 32'hc37ec06e},
  {32'h439cf82f, 32'h43c417e8, 32'h43a2e78f},
  {32'hc275b9c4, 32'h4397c57d, 32'h42c9d6fe},
  {32'hc30c4276, 32'h42ac3cc7, 32'h42f414ba},
  {32'hc1547ab6, 32'hc3080d49, 32'hc3c7a776},
  {32'h43a34854, 32'h43353b31, 32'hc1c3034a},
  {32'hc38a93cc, 32'h435a77ba, 32'hc2fa5d5c},
  {32'hc396c2f4, 32'hc35ee3bf, 32'hc3bb585a},
  {32'hc1d7b00c, 32'hc30aad69, 32'h430b25f5},
  {32'hc30b930d, 32'h43b7833a, 32'h42a0252e},
  {32'h421219f8, 32'hc3fada10, 32'hc321701e},
  {32'h44000917, 32'h440ce5d6, 32'hc3b3d6d4},
  {32'hc393fc3e, 32'h43a1a5be, 32'h43779b40},
  {32'hc38ecd93, 32'hc4010044, 32'hc3dd851e},
  {32'h41c60de8, 32'hc2470d73, 32'h43a6533f},
  {32'hc38abc0b, 32'hc36a5624, 32'hc34e5787},
  {32'hc2dd4db0, 32'hc36e6f38, 32'hc2d7b4a7},
  {32'h43468ec9, 32'h437db184, 32'hc20b54af},
  {32'hc1f101bd, 32'h436b3ea3, 32'hc381ff9e},
  {32'hc3b5d45c, 32'h42fdcac7, 32'h42956fcf},
  {32'h435e9083, 32'h428668a2, 32'hc2b51631},
  {32'h431581d3, 32'h438c0e15, 32'hc3285dad},
  {32'h4263941a, 32'hc2fc3e6f, 32'h42b33979},
  {32'h42af4362, 32'hc2e96bf7, 32'h431bacb6},
  {32'hc3bc9294, 32'h41b5a788, 32'h430a87c7},
  {32'hc382a663, 32'hc3a1a9c4, 32'h43ec1d91},
  {32'h434af48d, 32'h404ee870, 32'hc3d8c299},
  {32'hc2f7dffb, 32'h437b6371, 32'h432f4be4},
  {32'h437f934a, 32'h428d0494, 32'h42e356a4},
  {32'h41b6eeb8, 32'h4391f838, 32'hc29c703b},
  {32'h433f4abb, 32'hc41aceed, 32'h43d3b088},
  {32'hc3105e98, 32'hc2e427d1, 32'hc3e79bb3},
  {32'h421cc39a, 32'h44001863, 32'hc467da0c},
  {32'hc41e108b, 32'hc3731530, 32'h42a5eab4},
  {32'hc31e04c0, 32'h434a9ff6, 32'h433481fa},
  {32'h437eccca, 32'h433cd906, 32'h43c5cb33},
  {32'hc3f14f4e, 32'h43a736ad, 32'hc32f0643},
  {32'h431612d9, 32'h420b1481, 32'h42c98b0f},
  {32'hc31cbb57, 32'h4292b01d, 32'h4379d5aa},
  {32'hc2866627, 32'hc1a4d5f7, 32'hc33aeca6},
  {32'hc3dfe46e, 32'h433851c7, 32'h43dd5389},
  {32'h4266a842, 32'h430ceb54, 32'h42e1c728},
  {32'hc2a82f61, 32'h43b7dcbb, 32'h42461f9c},
  {32'hc3357bfa, 32'h42b422d9, 32'h42b601f1},
  {32'hc1555d99, 32'h43a7029e, 32'hc33a8c9b},
  {32'hc35569fd, 32'hc3697417, 32'hc2fdacc6},
  {32'hc3ae25b4, 32'h4299cff4, 32'hc3ca5a8c},
  {32'hc3807ab7, 32'h424203e0, 32'hc30e15c2},
  {32'hc2351aa1, 32'h4310ebf9, 32'hc2557b88},
  {32'h42a5fe7a, 32'h42fa7010, 32'h4317a829},
  {32'h427c5828, 32'hc30bdde1, 32'h4228e92c},
  {32'hc3e66be6, 32'h425aa7ff, 32'h430992ac},
  {32'hc391f33a, 32'h430f182a, 32'h43e90517},
  {32'hc2c978b5, 32'hc3969cb8, 32'h438c531f},
  {32'hc35c1bbb, 32'hc1ac0fc5, 32'h430c0787},
  {32'h42ebb856, 32'hc0ea8b8c, 32'hc30a40c3},
  {32'h42b34904, 32'h43e52f92, 32'hc326b396},
  {32'hc3410ae2, 32'hc3c14fc7, 32'h4305efe2},
  {32'h424064d9, 32'h42a39f06, 32'h4339d89e},
  {32'h43d563cd, 32'hc1c58e13, 32'hc33965b1},
  {32'hc2a5773e, 32'hc3535e3f, 32'hc3ca5c91},
  {32'hc3eb4276, 32'hc341ba72, 32'hc406ee2c},
  {32'hc3a3e77f, 32'h438c1d28, 32'h434a8644},
  {32'h43614390, 32'hc36851c2, 32'h43006772},
  {32'hc40307cb, 32'h43f4b4ca, 32'hc289cf06},
  {32'hc30c5bc8, 32'hc2479ca3, 32'hc24d2a21},
  {32'h435888dd, 32'h4327e9e3, 32'h430263a2},
  {32'h42a233ba, 32'hc309e96a, 32'hc3ab164e},
  {32'h42ca1b45, 32'h431be09e, 32'h435e9d42},
  {32'hc301f42e, 32'hc2ffa453, 32'h4396c0a5},
  {32'hc2cbdfb5, 32'hc1964d4e, 32'hc33f5814},
  {32'h4425cf30, 32'h43958df4, 32'h43ebc368},
  {32'hc3fdaaa8, 32'hc39c756d, 32'hc3269b6d},
  {32'hc3abdc84, 32'h422c0bd4, 32'h41751d5c},
  {32'hc2d03ef8, 32'h43d6f287, 32'hc237f804},
  {32'hc3a94a4d, 32'h42c6e849, 32'hc292d7f5},
  {32'h42436a71, 32'hc389971f, 32'h429c990c},
  {32'hc2956e14, 32'hc36f2b72, 32'h43708533},
  {32'hc164084e, 32'hc2a6cb18, 32'hc2c7ce57},
  {32'h42cf9704, 32'h436a8940, 32'h429d7aa6},
  {32'h42cee258, 32'h435e7f2c, 32'hc379c83d},
  {32'hc455eb56, 32'hc3b79469, 32'hc14f5afc},
  {32'h42e904f0, 32'h42b293e8, 32'hc20b3ba5},
  {32'h40799640, 32'h42cf73ba, 32'h42fdd927},
  {32'h420a1954, 32'hc2ca8178, 32'hc0fc0fd1},
  {32'h42621d9f, 32'h429973b2, 32'hc1bd2715},
  {32'h4397328c, 32'hc3b7c3f0, 32'hc40a35af},
  {32'hc3b188e0, 32'hc3ea6b74, 32'hc05bd44b},
  {32'hc351cd33, 32'h43583342, 32'hc3759529},
  {32'h439ef52e, 32'hc3c5d1c9, 32'h423cf177},
  {32'h438f4661, 32'h429e2f05, 32'hc3219493},
  {32'hc3c27f8c, 32'hc3b69e36, 32'hc243f323},
  {32'h440e15ed, 32'h438405da, 32'hc28a97d4},
  {32'h42ec8fbe, 32'hc12b3c06, 32'h434abe69},
  {32'hc423471d, 32'hc323f818, 32'h43163b1a},
  {32'h42e77603, 32'hc3165fe5, 32'hc38682b3},
  {32'hc3160a51, 32'hc2c933e9, 32'h429c55b7},
  {32'hc289ce7f, 32'hc3f592e9, 32'hc3c2e097},
  {32'h43e5572e, 32'hc332e13c, 32'h43e05fd9},
  {32'h42bc0c7e, 32'hc318f664, 32'hc2000dbf},
  {32'hc2d09b8c, 32'h438944a5, 32'h43e39bfd},
  {32'hc38d6778, 32'h42f690d4, 32'h4189cf22},
  {32'hc14547c0, 32'h4319e76d, 32'h43c47975},
  {32'h42da5aae, 32'hc2275dbb, 32'hc2aca143},
  {32'h43431b38, 32'hc39ebf3c, 32'h432cfd09},
  {32'h42ba9667, 32'hc291918c, 32'h42e2b414},
  {32'hc39819a4, 32'h420a5c1f, 32'hc35c5e8b},
  {32'hc39b5b9f, 32'hc38275c3, 32'hc39d95e2},
  {32'hc3ab35c2, 32'h42deea57, 32'h43c7fd2d},
  {32'hc37b4a2d, 32'h42d4cf9d, 32'h41fbeac4},
  {32'h437e07cb, 32'hc2ae5d6e, 32'hc399a438},
  {32'h418cb71d, 32'hc3d8d969, 32'h430ac24c},
  {32'hc3549299, 32'hc3b80e6c, 32'hc3bdf4ec},
  {32'hc2b6bc3e, 32'h43d36d1c, 32'hc2391b3c},
  {32'h41966349, 32'hc3b89045, 32'hc0d45d08},
  {32'hc37e918a, 32'hc3263b06, 32'hc3e6c889},
  {32'h431cda73, 32'hc3f62171, 32'hc3d658b8},
  {32'h4306b1ee, 32'h43701910, 32'hc352e271},
  {32'h40822a60, 32'h439d93ce, 32'h423be291},
  {32'h4403ba83, 32'h4379c6a6, 32'hc37ad932},
  {32'hc2f510f0, 32'hc2956128, 32'h4340ff0a},
  {32'hc3e6c844, 32'hc38d6492, 32'hc30f2fcc},
  {32'h43759cfc, 32'hc1940acb, 32'hc2b7928b},
  {32'hc398f490, 32'hc406feb1, 32'h4386829a},
  {32'hc3035644, 32'hc2c475a7, 32'hc006d9b3},
  {32'h44287b23, 32'hc3323462, 32'h43c41d14},
  {32'hc22f38ed, 32'h4391cd78, 32'hc3f04265},
  {32'hc28f7254, 32'h43b7892d, 32'h43b5e7f2},
  {32'hc30ffd50, 32'h43df5ee3, 32'hc222ee6f},
  {32'hc39dc411, 32'hc38ea49b, 32'hc33b617c},
  {32'hc29c474f, 32'hc3d2771c, 32'h432bc797},
  {32'h41c121ac, 32'hc38ccdb9, 32'h43188d29},
  {32'hc3c5270c, 32'hc292d553, 32'h435c7e43},
  {32'h4201a612, 32'h42ec2eac, 32'h41d93afa},
  {32'hc201d360, 32'h42d044b0, 32'h43b064d5},
  {32'hc40e1b25, 32'h43b8e7ad, 32'h43adff9d},
  {32'h41cef3b2, 32'hc3a3001e, 32'hc246095c},
  {32'hc2d288d2, 32'hc37b0902, 32'h434a4b73},
  {32'hc3626df5, 32'h43ca804c, 32'h43047660},
  {32'hc2ecfcc9, 32'hc354bfe5, 32'h42964182},
  {32'hc321ee0a, 32'h42fe126c, 32'hc353739e},
  {32'hc2c02767, 32'hc3aa4a71, 32'hc366b24c},
  {32'hc3056731, 32'h43a2757f, 32'h430cdf16},
  {32'h4306f4d8, 32'hc37700be, 32'hc38c6827},
  {32'hc3cbdbd0, 32'hc36131da, 32'h430dd329},
  {32'h430eac1a, 32'hc30bfd92, 32'hc1d5ea24},
  {32'h43342964, 32'hc30ccd92, 32'h4377f390},
  {32'h422f27e7, 32'h43bcf54a, 32'hc38f17f4},
  {32'hc434c759, 32'hc33abf58, 32'hc1b94705},
  {32'h43f21363, 32'h42dc129b, 32'h434b50a2},
  {32'hc38f09aa, 32'hc404028a, 32'hc281c36c},
  {32'hc3354db5, 32'h43cd6d07, 32'h43906035},
  {32'hc0971ba0, 32'h439da657, 32'h42392b88},
  {32'hc27a9599, 32'hc2efaffe, 32'hc29349ab},
  {32'h42fc5a2a, 32'h43ba8b1a, 32'hc391a243},
  {32'h424edb36, 32'h431f5b51, 32'h435356bb},
  {32'hc2d98fc6, 32'hc2ae51b3, 32'h43917550},
  {32'hc3155856, 32'h438436e1, 32'h42bca834},
  {32'h43a005cb, 32'h4338b53c, 32'h426a8474},
  {32'hc329ec80, 32'hc392a52e, 32'hc38dfc2c},
  {32'hc3dd202c, 32'h43c1472f, 32'h43b1cd57},
  {32'h43b08a34, 32'h43913771, 32'hc375e19b},
  {32'hc2aa4d3a, 32'h430ef55b, 32'h442b9dcf},
  {32'hc1aa1147, 32'h43af4e41, 32'hc3dc1876},
  {32'hc2ed78f3, 32'h43a97604, 32'h42183ec0},
  {32'hc3656cd7, 32'hc1c5b76f, 32'hc2fd256f},
  {32'hc2a6f628, 32'hc3ad5e31, 32'hc38ab196},
  {32'h428ef6b0, 32'hc3ccbd3d, 32'hc41b7434},
  {32'h4284f65d, 32'hc2d0db29, 32'hc31a1524},
  {32'h419449d4, 32'hc383289f, 32'hc3a83a92},
  {32'h4372a83b, 32'h4342e6e1, 32'hc4179207},
  {32'h4389562f, 32'h429a671e, 32'hc3957372},
  {32'hc3b54137, 32'h4299bafc, 32'h443147c7},
  {32'h4356837f, 32'hc339e067, 32'hc35050a3},
  {32'hc3410c75, 32'hc1b20a18, 32'h42f26d6e},
  {32'hc259191a, 32'hc3b21764, 32'h4294b6b5},
  {32'h43c782ae, 32'h438f84e8, 32'hc30d7c20},
  {32'hc3d38a57, 32'hc3a5962d, 32'h4341d6b4},
  {32'h42fe6de8, 32'h4292503a, 32'hc2de5604},
  {32'h43ed14d2, 32'h42f389f6, 32'h4329f8c2},
  {32'hc3c5f102, 32'h438fdc50, 32'hc316479e},
  {32'h423673cd, 32'hc3504337, 32'hc2b9a8e9},
  {32'hc3b09c16, 32'h44144208, 32'h42ac58c5},
  {32'hc378e67c, 32'h4411529c, 32'hc3600e5d},
  {32'hc3633e0b, 32'hc2b57b54, 32'hc3d0b599},
  {32'h43945f5d, 32'hc427e1d7, 32'hc2d973f5},
  {32'hc3a43016, 32'hc29d46c7, 32'h43981bac},
  {32'h42cfe258, 32'h43731682, 32'h404788e0},
  {32'hc3956f67, 32'hc2e0de89, 32'hc2bb0ba8},
  {32'hc43360c4, 32'h43c168ee, 32'h44039c09},
  {32'h42c34314, 32'h442bcb0d, 32'hc3b945d7},
  {32'hc33b421a, 32'h43ab4132, 32'hc203d525},
  {32'h432fadcd, 32'h433fae52, 32'hc21b268a},
  {32'hc28f88b7, 32'h43542aaf, 32'h436f990e},
  {32'h43a17e2d, 32'h428c6116, 32'hc32fccaf},
  {32'hc3c00628, 32'hc2f3ab15, 32'hc31f1c6b},
  {32'h412d1756, 32'hc388de46, 32'hc425034d},
  {32'h40126fc8, 32'h43cfe982, 32'hc2cbca35},
  {32'h42ef0479, 32'h4304a0d2, 32'hc31023a3},
  {32'h4264a424, 32'h435e5717, 32'h424a0bfc},
  {32'hc35044fb, 32'h41411550, 32'h443e4320},
  {32'hc2c24f0e, 32'h43d5ebac, 32'h43036e33},
  {32'h4394e365, 32'hc31ad730, 32'h43a84e55},
  {32'h429f1c9e, 32'h435de071, 32'hc2bf3aef},
  {32'hc2d5fb65, 32'h433019cd, 32'hc2922161},
  {32'h43b33ef2, 32'hc30464ae, 32'h42a0a1ed},
  {32'h4381fbba, 32'h4345c382, 32'h4284fd98},
  {32'h43209b51, 32'h415b05fc, 32'h412332b1},
  {32'h42be2be9, 32'hc374f8e8, 32'hc150f19c},
  {32'h4013b779, 32'h43c75112, 32'h43b00efe},
  {32'hc380fb27, 32'hc3ac69b9, 32'hc2ae903a},
  {32'h43a85369, 32'h42b2d3af, 32'h4299b4d7},
  {32'h42a9df06, 32'hc30a786d, 32'hc3d13ef8},
  {32'h44058cf8, 32'hc3d61a32, 32'h43cc7a67},
  {32'h420a5dca, 32'h4303cfbe, 32'h42aa13d4},
  {32'h432d55b8, 32'hc3b99193, 32'hc3c94157},
  {32'h43223968, 32'h43454da4, 32'hc3388a19},
  {32'hc30ab738, 32'hc32069ec, 32'hc20dfaaa},
  {32'hc3373c94, 32'h4314476b, 32'hc38f45d1},
  {32'h43908adf, 32'h41d90358, 32'hc2553693},
  {32'hc3629070, 32'h43c7b1ce, 32'hc3776572},
  {32'hc2a2d776, 32'h4255738c, 32'h43749529},
  {32'h4230eebe, 32'h4325c507, 32'hc39fd576},
  {32'hc37c892d, 32'h4304c92f, 32'h42e3d037},
  {32'hc2fb63fc, 32'hc32c37d9, 32'h43269e12},
  {32'h441ac51f, 32'hc20e747d, 32'hc2dc6022},
  {32'hc3845015, 32'hc326f8bd, 32'h432eb827},
  {32'h43a36a34, 32'hc321fe45, 32'h434b73a3},
  {32'hc23708da, 32'h4347d97e, 32'hc351f9dd},
  {32'h426e643c, 32'hc3c88a2d, 32'h437f7956},
  {32'h4309b527, 32'hc34d09ac, 32'hc3164201},
  {32'h423a60aa, 32'hc3b780e6, 32'hc2384e7c},
  {32'hc3613e00, 32'h428ebc6a, 32'hc2a061bc},
  {32'h43eb55d0, 32'hc2d159af, 32'h439d26e4},
  {32'h42938a11, 32'h42bfb83c, 32'hc27d5f27},
  {32'hc37f3ec7, 32'h43e6927c, 32'hc3ca727f},
  {32'h41b04660, 32'h42baf5c8, 32'h435d64c4},
  {32'hc328b268, 32'hc360e59e, 32'h42317745},
  {32'hc30885f5, 32'hc214a93d, 32'hc2a01138},
  {32'h42214fb5, 32'hc3c5f182, 32'h4387c17d},
  {32'h3f7fc400, 32'hc2d46bed, 32'h429e7552},
  {32'h4386afdc, 32'hc40ee408, 32'h43a7d2ae},
  {32'h420d983d, 32'hc32181ad, 32'hc28cdcc5},
  {32'h440bdf98, 32'hc3b8c950, 32'h438710cf},
  {32'h41c3c4bc, 32'h43871454, 32'h42d3670e},
  {32'h4319ee63, 32'hc3dceb0a, 32'h401cf19e},
  {32'hc1dcb59e, 32'hc396a1c2, 32'h43bfdac2},
  {32'hc346e5e7, 32'h41329e61, 32'hc40303b6},
  {32'h43f720b0, 32'h4283dfb3, 32'hc262f75b},
  {32'hc403e671, 32'hc3974c0f, 32'h42008cbd},
  {32'hc3e79b8a, 32'hc0dbacec, 32'h42ba572e},
  {32'h43cfba59, 32'h42bb5463, 32'hc30e8b73},
  {32'h4433507c, 32'h423698cd, 32'hc3be4ce5},
  {32'hc388bdb2, 32'hc3c66aab, 32'h434e060c},
  {32'hc2f7afed, 32'hc3d8aa32, 32'hc37d655f},
  {32'h435be93a, 32'h439fb8f4, 32'hc3b5d915},
  {32'h44045fdb, 32'h41b2dba9, 32'h42ba394f},
  {32'h41ad5e8b, 32'hc2f59bd7, 32'h439b0f7e},
  {32'h42ec5028, 32'h4385075a, 32'hc24a537c},
  {32'hc31ff2f4, 32'h42c8b4e3, 32'h42c817e8},
  {32'hc3016b53, 32'h4356ffe0, 32'hc2b7b700},
  {32'hc39a847e, 32'h43ac812c, 32'hc2cd51a5},
  {32'hc2b9a04e, 32'h43ff0ef3, 32'hc3f7f818},
  {32'h43805e33, 32'h4411ad19, 32'h42479d4a},
  {32'hc3f8d614, 32'h431429c0, 32'hc38cca25},
  {32'h439a0f9d, 32'hc37782a1, 32'h43087668},
  {32'h4305de46, 32'hc3a7d424, 32'h41dd5a62},
  {32'h4248fbbd, 32'hc2e17ac9, 32'h42959ba4},
  {32'h43a5552d, 32'hc33faf6f, 32'hc2db6ae3},
  {32'hc2b2a3d6, 32'h43699fb0, 32'hc355fe61},
  {32'hc2dd2b8b, 32'hc2ae9f46, 32'hc356d4cb},
  {32'h429ab7de, 32'h43408d33, 32'h442d6434},
  {32'hc2cf5b43, 32'h4386f4cb, 32'hc335151a},
  {32'hc3c8eb4d, 32'h43143c5f, 32'h43036fed},
  {32'hc3bb2f10, 32'h432a839b, 32'h4368806b},
  {32'h441596a0, 32'hc2f33d1a, 32'h428768d6},
  {32'h43133c66, 32'hc3aa7e31, 32'h43147e58},
  {32'hc39a4695, 32'h433d4aca, 32'h4349940d},
  {32'h43791af3, 32'hc33755bc, 32'h43dcc1df},
  {32'hc3cf67a8, 32'hc44a48f9, 32'hc3e8c7e4},
  {32'h4261c85e, 32'h41d3c9f8, 32'hc2e5a60b},
  {32'h43c767b9, 32'h42f1ec2b, 32'h42f4368a},
  {32'h4323982c, 32'h43001bbf, 32'h41afd0a8},
  {32'hc2b82328, 32'h435a9560, 32'hc3d93a6c},
  {32'hc31db968, 32'hc28c2757, 32'hc3533cc0},
  {32'h42cee2f6, 32'hc330c0e9, 32'h42b70701},
  {32'hc3dbfa84, 32'h419af013, 32'hc29ce916},
  {32'h438f3034, 32'h4264c5c6, 32'h43ba58e7},
  {32'hc3c1f13a, 32'hc3cbe095, 32'hc365c291},
  {32'h4233594f, 32'hc39680a0, 32'h4311980c},
  {32'h43540587, 32'h43961a6b, 32'h43afba69},
  {32'hc22f748a, 32'hc2f606ec, 32'h438ab3da},
  {32'hc300adac, 32'hc2bf68d8, 32'hc34f05e1},
  {32'h4382b3d0, 32'hc3d6baa0, 32'h43b5c8cc},
  {32'hc2d20834, 32'hc2619c85, 32'hc3d26fbe},
  {32'h42086ba0, 32'hc277c898, 32'h438187c6},
  {32'hc3443d01, 32'hc37b4c90, 32'hc42e4518},
  {32'hc196ae35, 32'h438168a6, 32'h429955ed},
  {32'hc2b05c4d, 32'h43e32c12, 32'h43398220},
  {32'h433fa4e3, 32'h42f5eb52, 32'hc39d8126},
  {32'h415dcd4e, 32'h42fa5eff, 32'h43990d95},
  {32'hc1d3b514, 32'h43112c10, 32'hc33c6e01},
  {32'h43dd7381, 32'hc3071697, 32'hc30da276},
  {32'hc3ed8124, 32'h42aaa67d, 32'hc208f83c},
  {32'h42e4b550, 32'h429ca65d, 32'h43b4e008},
  {32'h43da7fff, 32'hc33cde54, 32'h42cf609a},
  {32'h43815ce3, 32'hc334cf5f, 32'hc2fc643c},
  {32'hc33143c8, 32'hc397a30b, 32'h43af12f9},
  {32'h433ff217, 32'h430fb20a, 32'h43fdb845},
  {32'hc3a58838, 32'h42d1cb44, 32'hc3c1d933},
  {32'hc29f8c6e, 32'hc3556693, 32'h43382d1f},
  {32'h439c325b, 32'h43524c7e, 32'h43310ec5},
  {32'hc343a5d0, 32'hc3a47b7b, 32'hc13c9204},
  {32'hc399baa5, 32'h4387b951, 32'hc3147eb9},
  {32'h440bac04, 32'hc34b1cc6, 32'h43c74e3d},
  {32'hc21b25c5, 32'h438b5198, 32'hc3a6aa47},
  {32'h43c8685f, 32'hc299919b, 32'h429785de},
  {32'h423512f8, 32'h41c8ab69, 32'hc3983bf4},
  {32'hc334a3a1, 32'h4381bba4, 32'hc385fd62},
  {32'hc0ee48cc, 32'hc3b2bdfd, 32'h442bcf4d},
  {32'h42d01d9c, 32'hc3d538be, 32'hc40bfd91},
  {32'h42be719e, 32'hc3816630, 32'hc2d67c1a},
  {32'h431f024d, 32'h42535abd, 32'h41f4e6c9},
  {32'hc3a7e975, 32'h4354e8bd, 32'h42d6067a},
  {32'hc31f3c3f, 32'hc1d3b7e5, 32'h42baa317},
  {32'h4376afd0, 32'h4307d297, 32'h432dd270},
  {32'h43e37d27, 32'hc316dfce, 32'hc3dff5b1},
  {32'hc3bb45c4, 32'hc308f962, 32'hc02e8a41},
  {32'hc3394e2e, 32'hc3693085, 32'hc32146cb},
  {32'hc1e03f5f, 32'hc2bb169d, 32'hc30d0c63},
  {32'h43b5a7a5, 32'h42e84faa, 32'h436c9322},
  {32'hc3b1b220, 32'h434f0bd1, 32'h43615e97},
  {32'h43143bcb, 32'hc39ef5c3, 32'h437fd756},
  {32'h4392b4a5, 32'hc2cd90bd, 32'h42f2c4cd},
  {32'h408097e0, 32'h42bb1aa6, 32'hc2fb8c55},
  {32'h4386f1d4, 32'h3e3df900, 32'hc3a5ee65},
  {32'hc21a789e, 32'h4379212c, 32'hc3952552},
  {32'hc3002240, 32'hc3378c38, 32'hc3190bff},
  {32'h438ed75a, 32'h42005272, 32'hc3995a17},
  {32'hc36bef3a, 32'h43af1c8b, 32'hc2bd8642},
  {32'h43259a93, 32'hc34bd08f, 32'h438cec0e},
  {32'hc2a78676, 32'h431969ef, 32'h43724c4a},
  {32'hc3c7c288, 32'h43899c81, 32'h421dcca3},
  {32'hc2aa27dc, 32'hc3c27ca1, 32'hc34442fc},
  {32'h43621f61, 32'hc3048771, 32'h441d8f52},
  {32'hc34ebb8e, 32'h42451138, 32'hc155d1dc},
  {32'hc3f8f7cd, 32'hc41405cd, 32'h4214c3ab},
  {32'h43b52922, 32'hc3dabe04, 32'h438daa89},
  {32'hc42fa9a5, 32'h430a985e, 32'h4291562b},
  {32'h42129ac0, 32'hc2eea0c3, 32'hc3468c03},
  {32'hc368ba06, 32'hc312a946, 32'h4206b9a5},
  {32'h43347d10, 32'h437d3604, 32'hc393b603},
  {32'h42e9c5dd, 32'hc3346097, 32'hc3193760},
  {32'h42928d20, 32'hc354513e, 32'h435693eb},
  {32'hc3bfac5b, 32'hc3b85275, 32'h4208c398},
  {32'hc2ee6f38, 32'hc2ee4f1e, 32'hc3d529b9},
  {32'hc1de0520, 32'hc3c43ea6, 32'h4357b342},
  {32'h4397d5af, 32'hc2c98652, 32'h436fa19c},
  {32'h410d2673, 32'hc38780ab, 32'hc3ae1b82},
  {32'hc346e90f, 32'h4342e7eb, 32'h4332c504},
  {32'hc26dcf4d, 32'h42972898, 32'hc33ee38d},
  {32'hc3734133, 32'h43f0a149, 32'h43d88c7c},
  {32'hc3805482, 32'h4336dd7d, 32'h43e23b40},
  {32'h425e4893, 32'h43fdf995, 32'hc16af022},
  {32'hc250e2ba, 32'hc2e05148, 32'h4359e713},
  {32'h43c50fb6, 32'hc2b0416a, 32'hc3d04da3},
  {32'hc37fb17d, 32'hc235e1ad, 32'h43d10336},
  {32'hc1cf6150, 32'h42fe6730, 32'h43011969},
  {32'h43ad9e84, 32'h42fa8e68, 32'hc3cba2b0},
  {32'hc3b15c6e, 32'h43462449, 32'hc232a59e},
  {32'h42f33033, 32'hc3b8f524, 32'h41a493d3},
  {32'h43ab5cb8, 32'hc349e5fa, 32'h43bb21b9},
  {32'hc2ad5eee, 32'hc0574395, 32'hc41439de},
  {32'hc2c208fe, 32'hc2f865e7, 32'hc30959bc},
  {32'h44134af8, 32'hc3ae81ee, 32'h44292bd9},
  {32'hc25d02d6, 32'hc38bab52, 32'h42b1bdf7},
  {32'h4228acd6, 32'h4090f5d0, 32'h426af519},
  {32'h435b70b3, 32'hc308a3c0, 32'h4315dcc3},
  {32'hc419671f, 32'h426cf366, 32'h4340893a},
  {32'hc3328f16, 32'hc2e9efb1, 32'h4379b9e5},
  {32'h4302a638, 32'h4380100f, 32'hc3a11800},
  {32'hc3d9f64d, 32'hc399b197, 32'h41de2cf9},
  {32'h435dbf92, 32'h4384e91a, 32'hc2440401},
  {32'h43f4bd88, 32'hc3989030, 32'hc337b4c7},
  {32'hc32a5998, 32'hc1e839f8, 32'h42b7843f},
  {32'hc3aecd47, 32'h438f1bc0, 32'h4358231f},
  {32'hc2f61d89, 32'h43a1cce5, 32'h437db04a},
  {32'hc3355af0, 32'h43757fec, 32'hc13a9738},
  {32'hc3baaa00, 32'h41485558, 32'hc3f1d3a5},
  {32'h42709ae1, 32'h4301c19e, 32'hc2c33a1e},
  {32'hc1994d64, 32'h4411f84e, 32'hc2ca071d},
  {32'hc4292d5e, 32'hc390393a, 32'hc2fcd323},
  {32'h43041e84, 32'h3fccd994, 32'h4387e46e},
  {32'hc3b6ba5e, 32'hc32a06ef, 32'h439ca79e},
  {32'hc37391d5, 32'hc3bad7be, 32'hc292266f},
  {32'h42e52395, 32'hc2c32122, 32'h41f69e01},
  {32'h416cc77e, 32'hc2fc8c59, 32'hc3b0d6b2},
  {32'hc3efeac3, 32'hc290fe47, 32'hc38688a3},
  {32'h4309ecab, 32'hc35b0ba8, 32'h4427faa2},
  {32'h42eacbe0, 32'h433b2a7a, 32'hc15e5122},
  {32'hc39aef45, 32'h41cdbf65, 32'hc304e9d7},
  {32'hc13b8458, 32'hc31ed2fa, 32'hc306694c},
  {32'hc37b2bb6, 32'hc2dcba21, 32'hc382bf60},
  {32'h419196b0, 32'hc205115d, 32'h439a95e3},
  {32'h430e8ac2, 32'hc3645dc3, 32'h42b13c04},
  {32'hc2841892, 32'hc2570bf0, 32'hc3fd60b9},
  {32'h439184d0, 32'h4267583f, 32'h434b46ee},
  {32'h433b9332, 32'hc278d1f7, 32'hc1d8e606},
  {32'h43143c20, 32'h4367d7b7, 32'h4347880b},
  {32'h42b20929, 32'hc305ac15, 32'hc3c0a9cc},
  {32'hbf9bab80, 32'h4400394a, 32'h42c891df},
  {32'hc28fd935, 32'hc3b1df7b, 32'hc3adeee6},
  {32'hc241a7ac, 32'h4315eb15, 32'h43a7de40},
  {32'h4348588f, 32'h42ba3130, 32'hc40d48b9},
  {32'h43553cf1, 32'hc33398a8, 32'hc1c0eef9},
  {32'hc21f66c6, 32'h404eb838, 32'h43b8c0a4},
  {32'h4351d345, 32'h43006920, 32'hc2ff9143},
  {32'hc36524dc, 32'h42f050b6, 32'h42d3d16d},
  {32'hc3579011, 32'h42d6636a, 32'hc19195c2},
  {32'h43549ea8, 32'hc23d6027, 32'hc3c95fdb},
  {32'hc1cd2aca, 32'h431e2b76, 32'hc22da227},
  {32'hc3d28c3c, 32'hc38397e7, 32'hc2c93f7c},
  {32'h429581f0, 32'hc3995698, 32'hc32400e4},
  {32'hc401fbe4, 32'hc4002e74, 32'h4221619c},
  {32'hc406ff92, 32'h41e5d88e, 32'hc426722c},
  {32'h43006e2d, 32'h43ed3f04, 32'hc1a8f72d},
  {32'hc390258c, 32'hc400c0f9, 32'hc26ae59e},
  {32'hc3467d8e, 32'hc391fd43, 32'hc20e0607},
  {32'h4334de94, 32'hc3ec559c, 32'h440b2cdb},
  {32'hc377029c, 32'hc380b348, 32'hc32adef9},
  {32'hc325f216, 32'h4234acad, 32'h43301155},
  {32'h4383bc16, 32'h43177fac, 32'hc3be45af},
  {32'hc3f3a828, 32'h43b856f6, 32'h439dc9ac},
  {32'h43a8886c, 32'h4302d7a4, 32'h43b8fe4f},
  {32'h421bdbfd, 32'hc3456bb8, 32'hc34467a0},
  {32'hc34442a2, 32'hc40dc804, 32'h42b28dd9},
  {32'hc372a71c, 32'hc0620900, 32'hc31a3b99},
  {32'h42a7ec81, 32'hc3fd26d7, 32'hc2f2525a},
  {32'h435ab272, 32'hc3c7c8f2, 32'h435fa7af},
  {32'h42a77cc2, 32'h422b2602, 32'hc32d3220},
  {32'hc302090b, 32'h42cb53c0, 32'hc1e5af43},
  {32'h433c4628, 32'h434bd6c9, 32'h43f1a626},
  {32'h42092ecb, 32'h428d321a, 32'h43c05f4c},
  {32'hc2cfb0c9, 32'h4354fb3a, 32'h43991c2c},
  {32'h430b1fad, 32'h43c2d429, 32'h43a49adf},
  {32'hc343fe64, 32'h42abfbd3, 32'hc2ae0b9b},
  {32'h43b8de11, 32'h42625f3c, 32'hc31016b9},
  {32'hc3036886, 32'h42dc081b, 32'h432a6682},
  {32'hc258ca78, 32'hc26a37c6, 32'h4277a395},
  {32'hc2b53e0e, 32'hc11e8696, 32'hc3ddc1aa},
  {32'hc3bf408f, 32'hc3cb05c4, 32'hc34a7bd1},
  {32'h42312eb8, 32'h434ce346, 32'h43488d2c},
  {32'h42b43fbf, 32'h43044bd3, 32'h42eb3a85},
  {32'h42a157c6, 32'h440d6354, 32'h41df4518},
  {32'h43a4b16e, 32'hc3304296, 32'h41d91a71},
  {32'h4343733e, 32'hc3892a25, 32'hc33539bb},
  {32'hc3a7cf69, 32'h4354fcc2, 32'h4310c54f},
  {32'h432e959c, 32'h40cd6780, 32'h42f71d88},
  {32'h42887c0e, 32'hc37d41a7, 32'h42c5c6c8},
  {32'h43b4da05, 32'h43a13b6f, 32'hc3b19c96},
  {32'hc32cad94, 32'hc2b16971, 32'h423dc775},
  {32'hc2b56130, 32'h43b2c2d6, 32'hc42a06c7},
  {32'h41ade24a, 32'h42f51269, 32'h439667fc},
  {32'hc21c05c6, 32'h417803db, 32'hc3da47b8},
  {32'hc1dcdec0, 32'hc34ea53c, 32'h431489e6},
  {32'hc3d5bd54, 32'h4355b473, 32'hc36d9f4a},
  {32'hc3911ae4, 32'h42f5cbaa, 32'h43540000},
  {32'hc33f7104, 32'h42688580, 32'h4334b6e3},
  {32'h440e54b7, 32'h426f8d8d, 32'h43023922},
  {32'hc3680b5b, 32'h43bd4858, 32'h441f8aa8},
  {32'h4364b0be, 32'h4364491a, 32'h425cb6c4},
  {32'h42146dd7, 32'h439bbf51, 32'hc2ec9f27},
  {32'hc3125f9a, 32'hc30d22c8, 32'h43317f19},
  {32'h42eb57f0, 32'hc2515887, 32'h427178eb},
  {32'hc3a6b142, 32'h432fad8a, 32'hc36fadfe},
  {32'hc422a071, 32'h430def9d, 32'hc3be0a57},
  {32'h42787477, 32'h4392e3b4, 32'h4395930d},
  {32'hc3d8df07, 32'h41b95884, 32'hc347d773},
  {32'hc36ef798, 32'h44385df6, 32'h42c71491},
  {32'hc3caf5d5, 32'hc35f7552, 32'hc31448a1},
  {32'h4314c985, 32'h4349fb7c, 32'hc1a41369},
  {32'hc3635839, 32'hc29eb268, 32'hc3ab4bd6},
  {32'h4384f21a, 32'hc26d3cee, 32'hc339c187},
  {32'hc2ae5e6c, 32'h4282ebb7, 32'h43b3cdfc},
  {32'hc392b18c, 32'h422023d3, 32'h44502b1f},
  {32'h431076dc, 32'hc279f458, 32'hc35a0e7c},
  {32'hc3a0caf6, 32'h43bf0510, 32'h4264ebe8},
  {32'hc406d757, 32'hc23b6b7e, 32'h43a418a6},
  {32'h42071ba4, 32'h42c36a73, 32'h4376542f},
  {32'h4398cc29, 32'h3fc270e0, 32'hc2e2f02d},
  {32'hc22a3310, 32'hc3028d4d, 32'h41e36673},
  {32'h43980146, 32'h42591cca, 32'h4391e2a7},
  {32'hc3189e93, 32'hc3648fd6, 32'h43a468cb},
  {32'hc31cc0e5, 32'hc02212a5, 32'hc2f8279f},
  {32'h438ca025, 32'hc31aeee5, 32'h43291d88},
  {32'h42679c90, 32'h424c456d, 32'hc1ecab9b},
  {32'h42d4ab6e, 32'hc342d807, 32'hc1c7f46d},
  {32'hc39de853, 32'hc2289c3e, 32'h433a664a},
  {32'hc145f3b0, 32'hc3d24c8e, 32'h41f65bca},
  {32'hc3149bee, 32'hc3c7134f, 32'h43bda4b0},
  {32'h431534da, 32'h42d1f72a, 32'hc38317f6},
  {32'h4365502f, 32'h40e150b8, 32'hc374b625},
  {32'h42e69556, 32'hc436ba39, 32'hc2a6b9bc},
  {32'h43e96d20, 32'h43a487ff, 32'h440463df},
  {32'hc323b165, 32'hc2d74385, 32'h42caeefc},
  {32'hc37d07f4, 32'h4399ae5e, 32'h431223de},
  {32'h42c51a38, 32'h4309d24e, 32'h42517940},
  {32'h42500c1d, 32'hc36ce904, 32'h42009c0a},
  {32'h42bfa2e9, 32'hc3b0dfdb, 32'hc351a042},
  {32'hc2ac8a5a, 32'hc3c159fa, 32'hc35913ca},
  {32'hc1373cd8, 32'h425be10d, 32'hc39f0e94},
  {32'h43a3a532, 32'h43f97738, 32'h42d29d54},
  {32'h42ea9f41, 32'hc3aacb82, 32'hc42136b4},
  {32'hc412ac3d, 32'h43bf6fc2, 32'h43a3f895},
  {32'h43448da9, 32'h4305b292, 32'hc0760049},
  {32'hc3203424, 32'hc286c8fa, 32'hc38ec60a},
  {32'hc3270b9c, 32'h438ad2c5, 32'hc29debf6},
  {32'h42f5e078, 32'hc2706a84, 32'hc30204ff},
  {32'hc2e385fd, 32'hc23ac688, 32'hc1b41b92},
  {32'h4318de0f, 32'h42275a33, 32'h42e241d1},
  {32'h4061f4c0, 32'hc2a6e5ca, 32'h42412652},
  {32'h439b6a8f, 32'hc3659def, 32'h41bd2050},
  {32'h43dd5512, 32'hc31ef39a, 32'hc2c1bc2f},
  {32'hc42c6bcc, 32'hc1b865ad, 32'h4092b9dc},
  {32'h4343aa4f, 32'h439b6d97, 32'hc2baa5c1},
  {32'h429bd938, 32'h43f5b5ea, 32'hc38feac0},
  {32'h40d231fc, 32'hc3a3874b, 32'h430b93c0},
  {32'h43f0a5aa, 32'h42aa228e, 32'h428128ec},
  {32'hc39a9016, 32'hc341f5ea, 32'h43b10499},
  {32'h43470992, 32'h4393fe43, 32'h4009bae0},
  {32'h430783d7, 32'hc417051a, 32'hc3619fdb},
  {32'hc353c619, 32'h3fcae488, 32'h4221dc47},
  {32'hc4279751, 32'h4399e421, 32'h436ccc32},
  {32'hc3425ec2, 32'h4412011f, 32'h432a9c27},
  {32'h42c11d34, 32'h42ca4246, 32'hc304145b},
  {32'h43c7df36, 32'h414343b6, 32'h4358c6bb},
  {32'h435bda1a, 32'hc29033cf, 32'h43e34ffc},
  {32'h418d6083, 32'hc2849303, 32'h42906c4e},
  {32'hc1b2d196, 32'h42c8aa18, 32'h43265e5d},
  {32'h43399334, 32'hc3eadba2, 32'hc3ae1bb1},
  {32'h4371c325, 32'h4295d0ba, 32'hc34800c4},
  {32'hc28acf72, 32'h428165c1, 32'hc26ea580},
  {32'h439e19fd, 32'hc2d4fd10, 32'hc19b9480},
  {32'h43b769cd, 32'h41d90264, 32'h42c7f7ef},
  {32'hc28f85ee, 32'hc2ec984a, 32'hc410691c},
  {32'h435b3ac0, 32'hc3c5201a, 32'h420aad69},
  {32'h42a3ce84, 32'hc43681d8, 32'hc331f97a},
  {32'h430c1426, 32'h429a8acd, 32'h419b0cef},
  {32'h42dc3341, 32'hc3c490e9, 32'h41a5501b},
  {32'h43908309, 32'h43949a2c, 32'hc3cc711d},
  {32'h43facbc7, 32'h42833733, 32'h4383f7b4},
  {32'h430e98bc, 32'h4403e5d8, 32'hc414940f},
  {32'hc4007fa8, 32'hc394dbb0, 32'h4077da59},
  {32'hc313ba8e, 32'hc326c327, 32'h42dfce9c},
  {32'h42f41ca0, 32'hc251831a, 32'hc31a9a96},
  {32'hc32f43a5, 32'hc329cfd7, 32'h432873b4},
  {32'hc3474426, 32'h41aa55dd, 32'hc38504e5},
  {32'hc30cb179, 32'h4238ecf2, 32'hc1a17b83},
  {32'hc422d558, 32'h43ad0bf7, 32'hc2c21b2a},
  {32'hc3f3dec4, 32'hc2ff6275, 32'hc42a7e6a},
  {32'h43a6ab30, 32'h439458a6, 32'hc375f7e1},
  {32'h41c47b28, 32'hc2499b1c, 32'hc2b5c6aa},
  {32'h436babcd, 32'hc3b0939d, 32'h422c46f6},
  {32'hc2e9fc18, 32'hc30399cb, 32'hc2b1e11f},
  {32'h436867a6, 32'hc2da055d, 32'h43eb8e3a},
  {32'hc35cd34c, 32'hc2f10b68, 32'h4420bad3},
  {32'h42ec4539, 32'h4174e640, 32'hc33f2346},
  {32'hc3c11d24, 32'h43418e00, 32'h4309fa06},
  {32'h43f20541, 32'h421f6786, 32'h442029a1},
  {32'hc3a8950b, 32'h42c8a36d, 32'h43e0adcc},
  {32'h43b73bd9, 32'h42d20fc4, 32'hc3b21276},
  {32'hc21a9f38, 32'hc38eb6e9, 32'hc2324e0b},
  {32'h4374181c, 32'h43bfab78, 32'h41b018c0},
  {32'h434b06cb, 32'h42e1cb57, 32'h42b12d47},
  {32'hc030d440, 32'hc233f70c, 32'hc3423ae3},
  {32'hc21f46e4, 32'h423deab8, 32'hc36f7c2f},
  {32'h43a78837, 32'hc20a53b5, 32'hc2d0778f},
  {32'hc29e6346, 32'hc00319cb, 32'h43a2c27c},
  {32'h4408f382, 32'hc19d532a, 32'hc3b7ea00},
  {32'hc274e696, 32'hc367b51e, 32'h43a72bc3},
  {32'hc40b008d, 32'hc37220e8, 32'h43f36e3f},
  {32'h44059a79, 32'h4350ef9a, 32'hc33e0182},
  {32'h435319d0, 32'hc3b03ff2, 32'h43f6532b},
  {32'hc02aaf00, 32'hc3c6492e, 32'h43808ee7},
  {32'h4439e091, 32'hc2e63e5d, 32'h4449b067},
  {32'h42a27f90, 32'h437a924e, 32'hc31fe2a2},
  {32'h42dbafc4, 32'h42e1570e, 32'h432add22},
  {32'hc1855e3a, 32'hc35dbfb5, 32'hc2682ee8},
  {32'hc20ae6ed, 32'h434bb8b5, 32'h42ebd59a},
  {32'h3f97c9d8, 32'h42af33b3, 32'hc305dc73},
  {32'hc33af392, 32'hc3d07194, 32'hbfb761f0},
  {32'h41bcac02, 32'hc214f906, 32'hc32e98aa},
  {32'hc38917ad, 32'h4204796c, 32'hc2fa46c4},
  {32'h41cf5d2b, 32'hc19c8b03, 32'hc1d84bcb},
  {32'hc3a32042, 32'h43a2b48f, 32'h43e0adcd},
  {32'hc39d4470, 32'hc27188b8, 32'h432ef7c4},
  {32'h42f30cdc, 32'hc33bd45f, 32'h43b7ac8d},
  {32'h4194f722, 32'hc24ecc5f, 32'h41faddde},
  {32'hc3307f64, 32'h422b537f, 32'hc364c538},
  {32'h438edbf7, 32'hc3228dea, 32'h4391ad62},
  {32'hc3448866, 32'h431e5a4e, 32'hc41b4733},
  {32'hc2df4e31, 32'hc22281dc, 32'h430b88a2},
  {32'h43384b8e, 32'h4080981e, 32'h43d8834b},
  {32'hc2b44e0e, 32'h4117af81, 32'h4422baf6},
  {32'h4037e14c, 32'hc3b6b341, 32'h433f1ef2},
  {32'hc2e943b0, 32'hc33acc78, 32'hc23bca90},
  {32'hc450abf0, 32'h42227994, 32'hc30615aa},
  {32'hc3052821, 32'h434e99fe, 32'hc258100c},
  {32'hc2a2231b, 32'h43b626e1, 32'h438d0935},
  {32'h42eb4948, 32'h43fc2208, 32'hc30a3fe3},
  {32'h4116ae08, 32'hc2f01739, 32'h432a0b12},
  {32'h42c7efdc, 32'hc1537645, 32'hc1ddf560},
  {32'h436f68d8, 32'h4352dbac, 32'hc39c5d08},
  {32'hc3b3f728, 32'h44111dda, 32'h4325fce0},
  {32'h44224680, 32'h441a7383, 32'h4339c493},
  {32'hc2a0e263, 32'hc137ff94, 32'hc395d7a9},
  {32'hc23371dc, 32'hc39ca2e7, 32'h43a242bb},
  {32'hc313a86d, 32'h3fcfe4e8, 32'hc2205a89},
  {32'h426a3104, 32'h42eb50bd, 32'hc25625a5},
  {32'hc23acc25, 32'hc0519693, 32'h42a31ea9},
  {32'hc2929d9c, 32'h4305af66, 32'hc3c03694},
  {32'h4384daf3, 32'h42177196, 32'h44358e45},
  {32'h43b1606d, 32'h43e4d1b8, 32'h42852886},
  {32'h41e86d99, 32'hc34b7ae8, 32'h42a88b26},
  {32'hc3542f6b, 32'h4190f416, 32'hc2719239},
  {32'h432097dd, 32'hc361a01e, 32'hc2f2e930},
  {32'hc28a7fb9, 32'hc382b161, 32'hc386d0a8},
  {32'hc323105b, 32'h438e42d8, 32'hc42af2cf},
  {32'hc3aa35df, 32'h4307bd69, 32'hc235d0d9},
  {32'h42d68fe9, 32'hc284a442, 32'hc26c4b3f},
  {32'hc3c0da31, 32'h423ae16c, 32'hc294ac35},
  {32'hc3d15515, 32'h435561b1, 32'hc2faf0c0},
  {32'h435fc65d, 32'h43829427, 32'hc4083971},
  {32'h440570be, 32'hc2896182, 32'hc2e73af7},
  {32'h435b1384, 32'hc36e8607, 32'hc2fb8bd4},
  {32'h431091f1, 32'h42f50f25, 32'hc17cbc9a},
  {32'hc29f37bb, 32'h41f87f90, 32'hc32d748d},
  {32'hc4041dd6, 32'hc2b9bd66, 32'hc2c0d642},
  {32'h43ac54c5, 32'h409596f3, 32'h4396fa7c},
  {32'hc323d511, 32'h42afa6bd, 32'hc34c150a},
  {32'h42ec9633, 32'h428d54b6, 32'h42a48278},
  {32'h42eb77e3, 32'h43981ba8, 32'h42cb1443},
  {32'h43068fa5, 32'hc349f99e, 32'hc24972fd},
  {32'hc382adcc, 32'hc3a3039c, 32'hc36d4dbb},
  {32'h430a7160, 32'hc3d12b6c, 32'hc2503c9c},
  {32'hc42a98ba, 32'hc2f9d2f3, 32'hc328a7fc},
  {32'h42849b12, 32'h412c9480, 32'h401b61b0},
  {32'h43744e30, 32'hc3104ca7, 32'hc31ac24a},
  {32'h4105f6bf, 32'h4421136e, 32'hc38d66a4},
  {32'h437e3e00, 32'hc3786d7b, 32'hc31d8ede},
  {32'h41c1c0f2, 32'h43740644, 32'hc396e5ae},
  {32'h434f7cff, 32'hc365e5f3, 32'h4343c6db},
  {32'hc192ccd5, 32'hc3935a2e, 32'hc345ff83},
  {32'h43a366a2, 32'hc408483a, 32'hc3ca7283},
  {32'hc2ceaed8, 32'h4341794e, 32'hc38d2c63},
  {32'hc15a8098, 32'hc10a5f1a, 32'h4316b509},
  {32'h42367e71, 32'h42b992c4, 32'h43dbfabe},
  {32'h42fac96e, 32'h43383ea3, 32'h414bc6c2},
  {32'hc32702d0, 32'hc2345af8, 32'hc2270cd8},
  {32'h442cf9dc, 32'hc2e2f4c4, 32'hc1ab1ef5},
  {32'h4310d031, 32'h425c83ce, 32'hc39cb800},
  {32'hc3286f2c, 32'hc30e36bc, 32'hc3bc801a},
  {32'h42929794, 32'h440f24b7, 32'h4353a88c},
  {32'hc3405bd1, 32'h41534f18, 32'h43a3f0cf},
  {32'h42d6661a, 32'h43597b24, 32'h43b1e839},
  {32'h421e216c, 32'h4234a404, 32'h43c1cda3},
  {32'h434a5708, 32'hc29bb8f9, 32'hc347b384},
  {32'hc3ae4322, 32'hc385fff1, 32'hc401182b},
  {32'hc2865cd0, 32'h43b7e870, 32'h4309e41d},
  {32'hc43678fb, 32'hc38e7bc2, 32'h438c02bb},
  {32'hc3910595, 32'hc36c6904, 32'hc3f9f1b8},
  {32'hc2b2217b, 32'h43b9f83e, 32'h420634e8},
  {32'hc0e6954d, 32'hc3844b92, 32'hc25a8eef},
  {32'hc3d51131, 32'h429672ac, 32'hc33d48f0},
  {32'hc36df7fa, 32'h43855279, 32'hc2823a1f},
  {32'hc1c6e780, 32'h4381bd5c, 32'h4276189e},
  {32'h434bdf27, 32'hc1d820c1, 32'h434038e8},
  {32'h4258b4b4, 32'h4323fd0e, 32'hc2a0286f},
  {32'hc380af29, 32'h42d492c2, 32'h43cd4893},
  {32'hc215920d, 32'h42bf10f5, 32'h4252c5d2},
  {32'hc222747e, 32'hc240f037, 32'hc321704f},
  {32'h43b2df39, 32'hc3192a59, 32'h4202f281},
  {32'hc3f90c45, 32'h43987edd, 32'h43896093},
  {32'hc196fea0, 32'hc39abb99, 32'h43ad82f7},
  {32'h43ae8511, 32'hc1c0875e, 32'hc330a5d0},
  {32'hc3b20859, 32'hc3da925a, 32'h439c6284},
  {32'h434e18ed, 32'h420d0da6, 32'hc298c254},
  {32'hc2d6a9ea, 32'h43e73865, 32'hc32fee85},
  {32'hc4114208, 32'hc32e36f9, 32'hc3786707},
  {32'h4422125a, 32'h43daa0fe, 32'hc3a125ea},
  {32'hc32d839a, 32'hc22ef804, 32'h4067b000},
  {32'h43047da8, 32'h42634d2d, 32'h428f007a},
  {32'h43e12d8e, 32'hc305dff5, 32'h4428775a},
  {32'h422941a0, 32'h4293b0a9, 32'h426147c4},
  {32'hc32e4527, 32'h440f8e8d, 32'h42ead0ab},
  {32'hc3c9ab68, 32'hc2a2989d, 32'hc27d31e6},
  {32'hc2c5b460, 32'hc3d9e5b3, 32'h41afba37},
  {32'h440e5b24, 32'hc33162db, 32'h4248c834},
  {32'h42f22b4c, 32'h4028ac46, 32'hc2ad238d},
  {32'hc3b87d1f, 32'hc2a1dddc, 32'hc2d06c02},
  {32'hc3b5b4fc, 32'h438b692d, 32'h439012e1},
  {32'h431e685b, 32'h410812ef, 32'hc3a4463b},
  {32'h4347f638, 32'h41be2da1, 32'hc367cfc7},
  {32'h4286b53d, 32'h415c8544, 32'hc362d2ef},
  {32'h43fe8d13, 32'h43bb73ad, 32'hc3c93da2},
  {32'hc2e6d062, 32'hc40e3c37, 32'hc21ffba2},
  {32'hc36c031c, 32'hc26d293e, 32'h4315a8b2},
  {32'h420fc0d0, 32'hc3c22aba, 32'hc2ebfda9},
  {32'h42a2eec1, 32'hc3b31d71, 32'hc302a604},
  {32'hc3063401, 32'h41cd7190, 32'hc3fdddc5},
  {32'h43546332, 32'h411ef770, 32'h42f6c470},
  {32'h43acc94e, 32'h42b7412c, 32'hc3b83986},
  {32'h40c123e0, 32'hc2e6702d, 32'h434dcb2f},
  {32'hc3adff65, 32'h43544b33, 32'h4395abc2},
  {32'hc325dab9, 32'hc3320b09, 32'hc1a0035a},
  {32'hc21adbd0, 32'hc33ff0a1, 32'hc3930847},
  {32'h4419d8c4, 32'h43d4f6b7, 32'hc3d2e99b},
  {32'hc308b82d, 32'hc2d20a92, 32'h42d93e6f},
  {32'h43409322, 32'hc339dd90, 32'h4218f325},
  {32'h441c5dd3, 32'h433f0398, 32'h4408e9b4},
  {32'hc30172c1, 32'h4399b6e2, 32'hc425084d},
  {32'hc28f668a, 32'hc347fe3c, 32'hc32c9208},
  {32'hc3353ce1, 32'h440dcdf0, 32'h431b75dc},
  {32'hc2e5ae49, 32'hc32b2373, 32'hc3184f2d},
  {32'hc21fe1d2, 32'hc373411a, 32'hc3f136da},
  {32'h4376f092, 32'h4219ef98, 32'hc3247d01},
  {32'hc2c92bb6, 32'hc32e0656, 32'h4203ecc3},
  {32'h41dfa3b8, 32'hc23166da, 32'hc27f5464},
  {32'h42b28a4a, 32'h4257c92f, 32'hc4016009},
  {32'hc384ffeb, 32'h43c1928f, 32'h43938fc3},
  {32'h426ff265, 32'hc28a25be, 32'hc2a754dc},
  {32'h43a9665e, 32'hc3211121, 32'hc2a8cec5},
  {32'hc36946e4, 32'h42c0726d, 32'hc2ba2877},
  {32'hc4462b1a, 32'hc3fae4a7, 32'hc285d2ce},
  {32'h42e83e64, 32'hc408c2a4, 32'hc419da77},
  {32'hc20d3d26, 32'hc2f9403e, 32'h4295fda4},
  {32'hc2955e58, 32'h4364e916, 32'hc2d7a283},
  {32'hc32dc219, 32'hc4075c1a, 32'hc36d3cbd},
  {32'h434b86b0, 32'hc32e469a, 32'h437bfebd},
  {32'hc34f91e2, 32'h42b1effc, 32'h439a7e75},
  {32'h44260230, 32'h4369e695, 32'hc38beb36},
  {32'hc3106cdd, 32'h4391871f, 32'h42f376bc},
  {32'h3e44ac00, 32'hc30a666a, 32'h4385769a},
  {32'h43219fd5, 32'hc1aad76b, 32'h43576b58},
  {32'hc3ea04b8, 32'hc3ba239a, 32'h4329d706},
  {32'hc1b6dc00, 32'hc3c30a31, 32'hc3eab1b3},
  {32'h43b6f818, 32'h427c7b99, 32'hc2eff526},
  {32'hc30a8dac, 32'h425744b8, 32'hc27d38a9},
  {32'hc3914a98, 32'h4213526d, 32'hc4638e75},
  {32'h442763be, 32'h4321ed0b, 32'h43446b9c},
  {32'hc355408c, 32'h42aa1f4b, 32'h41bb378b},
  {32'hc379ba67, 32'h41ced22c, 32'h423047bd},
  {32'h40f83d40, 32'hc3a58e8c, 32'h43044d2b},
  {32'h43426f4b, 32'h42b3f7ad, 32'hc1700bd0},
  {32'hc2c61930, 32'hc36871b8, 32'h43940d4f},
  {32'h4398e03c, 32'h438e198f, 32'hc3ba35d5},
  {32'h4311c0f8, 32'h43516018, 32'h43fbaea2},
  {32'h429f56be, 32'hc36de9be, 32'h432b9b7c},
  {32'h4389dbde, 32'h42036137, 32'h430ea159},
  {32'h4384a2c5, 32'h431ece05, 32'hc34b49e6},
  {32'hc3ab5566, 32'h42b64cc2, 32'hc35b1478},
  {32'h429085f6, 32'hc2cf363a, 32'hc29284f0},
  {32'h43379b64, 32'hc1f6d090, 32'h42da01a4},
  {32'hc0efe5f2, 32'h4358eda4, 32'hc34f1838},
  {32'h436f055d, 32'hc3a08408, 32'h41b12b3a},
  {32'hc2db05a4, 32'hc33a6c28, 32'h425dc1a9},
  {32'h42b2bd0e, 32'hc21cabfc, 32'hc45e8aa1},
  {32'h42bd818e, 32'h437e4670, 32'h42ef5ec3},
  {32'h40f01fa4, 32'h437638ae, 32'hc2b5e395},
  {32'hc3cb3cdc, 32'hc38b58a2, 32'h438704b2},
  {32'h42df94b6, 32'h423a4bf1, 32'h4341e4f6},
  {32'hc2a81cff, 32'hc30bd503, 32'h42a062ff},
  {32'hc29eccb8, 32'hc3a38dca, 32'hc3634a5c},
  {32'h44020570, 32'h431b06f8, 32'hc34a5c86},
  {32'hc3eac16c, 32'h4357e4f6, 32'hc376e637},
  {32'h43341789, 32'hc3b5365f, 32'h42861ff2},
  {32'h41b6eb66, 32'h43bed45c, 32'h43b87865},
  {32'hc284a21c, 32'hc3876e01, 32'hc3263c4f},
  {32'h424f3b50, 32'hc362aeb0, 32'hc29dd858},
  {32'h4325d39f, 32'hc1954cf6, 32'h42845f96},
  {32'h433f602a, 32'h42ec7b8d, 32'hc31b4d42},
  {32'h43a81103, 32'hc392b6bf, 32'h41b2a3e8},
  {32'h42e04669, 32'h420ec734, 32'hc375e1c9},
  {32'hc2ff2332, 32'hc17ca92a, 32'h43782331},
  {32'hc38d465b, 32'hc35142b1, 32'hc352cf93},
  {32'h41c56140, 32'hc1f503e8, 32'hc300d5e1},
  {32'h4398b454, 32'h4378c85e, 32'hc424a221},
  {32'hc3068786, 32'hc2d01703, 32'hc2bda6b0},
  {32'h43a6a45c, 32'hc291440c, 32'h41abf3f7},
  {32'hc3a2fae0, 32'h4331f777, 32'hc28c2cb3},
  {32'h4030dfcc, 32'hc3308433, 32'hc39f3ca6},
  {32'hc32ec262, 32'hc31b7300, 32'hc3a9354f},
  {32'hc3e708ae, 32'h42f8d056, 32'hc2c610c4},
  {32'hc3aa573e, 32'hc30eca20, 32'h433b61c7},
  {32'h440059e7, 32'h43693d68, 32'h41644d11},
  {32'hc357d1fe, 32'h4337dc8e, 32'hc40c4785},
  {32'h429bde88, 32'h42a94765, 32'hc3484bc0},
  {32'hc1db0e6e, 32'hc31b2ef7, 32'hc35c97d3},
  {32'hc4146f72, 32'hc27c4d0c, 32'h4413d775},
  {32'h42d81bc2, 32'hc3d5c7cc, 32'h440823e1},
  {32'h4349e3ea, 32'hc34307ee, 32'h43227dae},
  {32'hc366357a, 32'h4343b32b, 32'hc3945591},
  {32'hc397728f, 32'h424f1522, 32'hc2c92b18},
  {32'h42d813c2, 32'h433a2572, 32'h43907e0e},
  {32'hc3be5689, 32'h4412279c, 32'hc3721232},
  {32'h43cac1a4, 32'hc26f4358, 32'h43766d33},
  {32'h42aded86, 32'hc2eb585e, 32'hc390c36b},
  {32'hc42eecf3, 32'hc3ff8df6, 32'hc337da1f},
  {32'hc34c895e, 32'h43bdbba3, 32'hc31a7adc},
  {32'hc1fb59e8, 32'h4388d2d6, 32'hc3863499},
  {32'h434ad76a, 32'h43e18468, 32'hc3420936},
  {32'hc34f9c13, 32'hc34e9c1f, 32'h42c9b9d3},
  {32'h42733a12, 32'hc30c2e3a, 32'hc3221419},
  {32'h4332cdea, 32'hc296108c, 32'h42e351fc},
  {32'h4415f208, 32'h441052bb, 32'hc3e1b37c},
  {32'h4327d7d6, 32'hc16e2dfc, 32'h4348ea02},
  {32'hc3a1fe87, 32'h4299bc2b, 32'hc39a8672},
  {32'hc3820c48, 32'hc15cecd8, 32'h432c1e57},
  {32'hc281559f, 32'hc3d3fbbd, 32'h421b741f},
  {32'hc2fbed94, 32'hc25a13b3, 32'h433bbc12},
  {32'h40e9d780, 32'hc3647cdb, 32'h43aca6e4},
  {32'h4398c4b7, 32'hc29f2635, 32'hc3959f79},
  {32'hc312c70e, 32'hc3462af1, 32'h432a63e5},
  {32'h42511162, 32'h427678ad, 32'h4416a6ce},
  {32'h422c2273, 32'h43610094, 32'h42ab4a5f},
  {32'hc40ccab0, 32'hc3b3996c, 32'h425ed43b},
  {32'h42e70fca, 32'h4420ad4e, 32'hc20609bb},
  {32'hc1e9af00, 32'hc38a4ff3, 32'hc2ef6d40},
  {32'h4310b6c7, 32'h42f631cc, 32'h43847823},
  {32'hc3fe2c86, 32'hc36c824b, 32'hc38a071b},
  {32'h4292e654, 32'h4173721c, 32'hc04a95dd},
  {32'hc3014b98, 32'h41dc3cb3, 32'hc314484c},
  {32'hc2d4a71e, 32'hc2866024, 32'hc371ad19},
  {32'h44319858, 32'hc31b7f1f, 32'hc3853820},
  {32'h439a6888, 32'hc3a1b0bd, 32'hc3fceec5},
  {32'h43036245, 32'h42946508, 32'h41b6a8df},
  {32'h4248b85d, 32'h42f786b3, 32'h40d97fa8},
  {32'hc3948ebe, 32'h438d09e0, 32'hc2f53246},
  {32'h43c3deb4, 32'hc20e5515, 32'hc3186feb},
  {32'h43919f65, 32'h439b01fa, 32'h42d5618b},
  {32'h428fe95e, 32'hc35fbca9, 32'hc0eccba8},
  {32'h413e5ce0, 32'h4372b6b4, 32'hc2cccdd8},
  {32'hc280cc22, 32'h425428e0, 32'h41ab08f1},
  {32'hc3459c45, 32'h438a1102, 32'hc4459a7a},
  {32'hc297c022, 32'h43827420, 32'h42e27c61},
  {32'hc395fa99, 32'hc38168c2, 32'hc3723702},
  {32'h4399149d, 32'h42a0464f, 32'h437d44a6},
  {32'hc3d6e084, 32'h43ec32fb, 32'hc2982627},
  {32'h43b2dab6, 32'hc33fe3cf, 32'h419a1a97},
  {32'hc2a478e6, 32'hc303962e, 32'hc2d43808},
  {32'hc2eeeef4, 32'hc302122c, 32'h41ab7512},
  {32'h43a3ca0e, 32'h42986331, 32'h42cb6b85},
  {32'h43e415ea, 32'h429b76b6, 32'hc1d19864},
  {32'h438305dc, 32'hc233679b, 32'h43d40fd4},
  {32'h42cde55f, 32'hc37e9442, 32'h439c074f},
  {32'h43d7dc73, 32'h43907b2b, 32'hc3a966a4},
  {32'h41505b40, 32'h42a2afdd, 32'hc39012fb},
  {32'h4383b433, 32'h441e210f, 32'h42036b00},
  {32'hc21307d1, 32'h4277266f, 32'h420bb66e},
  {32'hc117b4d0, 32'hc25f38ea, 32'hc319efb7},
  {32'h436c2997, 32'hc20ea1dd, 32'hc1982c88},
  {32'hc35b6a1e, 32'hc32b759e, 32'hc2c33d10},
  {32'hc163b9cf, 32'h42a384ca, 32'h439fb526},
  {32'hc214d3dc, 32'h4185544b, 32'hc314736a},
  {32'h41be227c, 32'h4395d147, 32'hc3dadaa3},
  {32'h411ba040, 32'hc29012d4, 32'h440fad6b},
  {32'h43dba786, 32'h4391b61d, 32'hc3481d44},
  {32'h42d7c302, 32'hc427c095, 32'h43b34711},
  {32'hc15dfe34, 32'h42f44caa, 32'h430c4ab5},
  {32'h43a798ae, 32'hc35ed08f, 32'hc3b9f458},
  {32'hc3fa8c66, 32'hc313e47b, 32'h42d09dd4},
  {32'hc417bb0e, 32'hc2f56a19, 32'hc425f1a5},
  {32'hc3c3a853, 32'hc3e311be, 32'hc3f4ed9a},
  {32'h405ebc42, 32'hc34383e1, 32'h4356461a},
  {32'h42736bae, 32'hc32ae90c, 32'h439f98ba},
  {32'h42cda587, 32'h4323c3c7, 32'hc336f7d5},
  {32'h42a17f3a, 32'h43250991, 32'h4228dde6},
  {32'h43e3ea36, 32'hc3006c14, 32'h427a367b},
  {32'hc2d71afd, 32'hc3445553, 32'h43284ff7},
  {32'hc389e9a5, 32'hc3c715a8, 32'h438a64c5},
  {32'hc0186940, 32'h438789a6, 32'h43406a75},
  {32'hc340b622, 32'h4310ad10, 32'h427901c0},
  {32'hc33bdafe, 32'h4328c7eb, 32'h432f5987},
  {32'hc2f5abb9, 32'h43e8c2fa, 32'hc2c05183},
  {32'h43af50b6, 32'hc38d2923, 32'h43cc9d07},
  {32'hc3ee2d17, 32'h42db4e67, 32'hc3a80d24},
  {32'h438b6578, 32'hc319a08d, 32'h41af88f3},
  {32'h43ba3211, 32'hc323027d, 32'h43bb8f9f},
  {32'hc4222454, 32'hc3187192, 32'hc3f61bb3},
  {32'hc26cf18e, 32'hc37797d7, 32'h43715b4c},
  {32'hc3ca5e7e, 32'hc238337e, 32'h41bb05f6},
  {32'hc1f234d4, 32'h43337685, 32'h42ac8412},
  {32'hc1f45ce7, 32'hc2df7c0c, 32'hc336b98c},
  {32'h4382a937, 32'h4283cd22, 32'hc0a94ebc},
  {32'hc2ed86a6, 32'h4309f041, 32'h43e91487},
  {32'h41e8fcea, 32'hc414d612, 32'h435b09bf},
  {32'h442867de, 32'hc315d77d, 32'hc2dbb0e4},
  {32'hc3954760, 32'h4367f1b3, 32'hc306bf60},
  {32'h42bb43b5, 32'hc323940e, 32'hc3a1eee5},
  {32'h43aecced, 32'hc2c49b11, 32'hc2feda3b},
  {32'h43b8f048, 32'hc39655a9, 32'h41e3b91a},
  {32'hc2814278, 32'hbe98ed80, 32'h43dc3486},
  {32'h430a3f7b, 32'h4296bed6, 32'h43a3370b},
  {32'hc29b4040, 32'h440e91c4, 32'h4292696f},
  {32'hc4091be6, 32'hc2f2778a, 32'h4377d42c},
  {32'h43c577dd, 32'h42e9f491, 32'h43008fe6},
  {32'hc36aecad, 32'h4327705e, 32'hc3b53f39},
  {32'hc2ef3c30, 32'h4348ca61, 32'hc325f704},
  {32'h42deedae, 32'hc0cf0b14, 32'h42ad6388},
  {32'hc3d6e7d7, 32'h4388c34f, 32'hc380ba12},
  {32'hc3a43158, 32'hc2d7e7fb, 32'hc3f22666},
  {32'h43c8bea8, 32'h4417bf79, 32'hc2fa1fe8},
  {32'hc3371508, 32'hc3ec3880, 32'hc20afb96},
  {32'hc2cffe7e, 32'hc32f355c, 32'h42a195a7},
  {32'h43961b38, 32'hc370771f, 32'hc2bf1355},
  {32'hc3c8eb86, 32'hc133b530, 32'hc339a01b},
  {32'hc37f1534, 32'hc2a869b9, 32'h4357f85f},
  {32'h4354517f, 32'h439cb9fe, 32'hc349f536},
  {32'hc3af0cee, 32'h43db42ef, 32'h43c17269},
  {32'h430a14fb, 32'h4215b1f8, 32'h42f7cd0d},
  {32'hc34a357f, 32'h4353973f, 32'hc30f7185},
  {32'hc2aa53c8, 32'hc4245094, 32'h43526bfd},
  {32'h43286382, 32'hc32b88c0, 32'hc2a635a3},
  {32'hc142cfb0, 32'hc3159580, 32'h41d47b92},
  {32'hc3873b78, 32'h43a561fa, 32'hc25a06fa},
  {32'h418603f6, 32'hc39a4e32, 32'hc4198396},
  {32'hc3026534, 32'h4083c788, 32'hc2174c3a},
  {32'h41f46d2b, 32'h41953842, 32'hc396768b},
  {32'h4316350c, 32'h433c3072, 32'hc4158560},
  {32'h4405d44a, 32'hc25ce1b4, 32'h4283a39c},
  {32'h4348b0c7, 32'h426017c0, 32'hc313c3f4},
  {32'hc3b9f67b, 32'hc33119bd, 32'hc37e72d2},
  {32'h440aa094, 32'h43932fe9, 32'hc1625581},
  {32'hc3a722ce, 32'hc2330cc5, 32'h43417aa4},
  {32'hc15188a8, 32'h419b29d3, 32'h42921886},
  {32'h42a61068, 32'hc3a303e1, 32'h42d556ac},
  {32'h40dbcc60, 32'h440c9851, 32'hc38c6263},
  {32'hc23762e0, 32'hc29d4b60, 32'hc3367e9a},
  {32'h42619bb0, 32'hc32daad6, 32'h43921a28},
  {32'hc0c32a20, 32'hc3a6c2c0, 32'h41fd8bf5},
  {32'h434cd214, 32'h432a85d5, 32'hc2deb12d},
  {32'hc2044364, 32'hc40888cf, 32'hc33b8d59},
  {32'hc410a4ec, 32'hc32e2111, 32'hc2c0444a},
  {32'hc32a95b7, 32'h422ebecb, 32'h4342e686},
  {32'hc1ea7a6e, 32'hc0c0c9fc, 32'h4247ee56},
  {32'h4365c019, 32'hc3afdebb, 32'hc1052aed},
  {32'h410e760a, 32'h426e8b06, 32'h42d10bc5},
  {32'hc2e390a8, 32'h42ac6d0b, 32'hc33398a5},
  {32'h4369c1b8, 32'h4377a0c7, 32'hc41af7ac},
  {32'h43ae018d, 32'hc2c419d6, 32'hc2e5cfa7},
  {32'h441791ee, 32'hc30967a4, 32'h42d4b14e},
  {32'hc3a3928f, 32'h41a25c90, 32'hc2bba31e},
  {32'hc3bfba16, 32'h43e165db, 32'h430fb41c},
  {32'hc22b4148, 32'hc214b502, 32'h42b1652b},
  {32'h44417cea, 32'hc19da5d4, 32'hc352b4ba},
  {32'hc3d9ffdf, 32'h437188f5, 32'h43cf8fb3},
  {32'h444f69c3, 32'h42ea0c7a, 32'hc3dddfc5},
  {32'hc40e1b8d, 32'hc337d813, 32'h432589f7},
  {32'hc2b7ade8, 32'hc43e5e08, 32'hc40d22bc},
  {32'h4388062d, 32'h42fab38c, 32'h424c8b9d},
  {32'hc2bdc234, 32'h41ace806, 32'h42e44116},
  {32'hc35ff31a, 32'hc3a2d8f6, 32'h43139fb1},
  {32'h44131468, 32'h43537605, 32'hc27a5110},
  {32'hc394792b, 32'hc369dbd6, 32'h42c8a54b},
  {32'h439fd2f9, 32'h43ea68e8, 32'h436cf481},
  {32'hc1297acc, 32'h4403857e, 32'h41c28607},
  {32'hc2762e3f, 32'h4396e187, 32'h43a552d0},
  {32'h42e85498, 32'h41ccd1e4, 32'h429d9b10},
  {32'h41b6b95d, 32'hc37ad4ad, 32'hc2e85494},
  {32'hc1dfe084, 32'h42a66340, 32'h4353f2a6},
  {32'hc221c7d6, 32'h42e5cb79, 32'h42235882},
  {32'h423b7c2d, 32'h421e6ef6, 32'hc38b4b0a},
  {32'h41aca052, 32'hc4302c31, 32'hc211f8a5},
  {32'h423039fe, 32'hc2a69e76, 32'hc2e3db0c},
  {32'h43d620a3, 32'hc3c0047f, 32'hc3a780fd},
  {32'h41fcf1e8, 32'h4146c45f, 32'h439bc578},
  {32'hc32fc9a4, 32'h43aefb3c, 32'hc400cb6b},
  {32'hc30dc704, 32'hc3956cb6, 32'hc3707a5d},
  {32'hc305ac48, 32'hc340c4b6, 32'hc2483d1d},
  {32'hc368f9d2, 32'h4068ccc0, 32'h43927283},
  {32'h42708735, 32'h4269402f, 32'hc389fefd},
  {32'hc1aef7f1, 32'hc2cf7314, 32'h43835a98},
  {32'hc3d3a630, 32'h42ca5548, 32'hc4121a0e},
  {32'hc382c70d, 32'h431410d9, 32'h42fa1730},
  {32'hc353e008, 32'h41bb6b8c, 32'hc2aa0659},
  {32'hc3c2c44c, 32'h4363e3ca, 32'h4406c5f2},
  {32'h43431965, 32'hc1e95a7e, 32'h42aa2604},
  {32'hc2fd2a99, 32'h43816575, 32'h440b67c3},
  {32'h43cec1f6, 32'hc391bad6, 32'h43d51c8e},
  {32'h40a7d4b0, 32'hc31a569d, 32'h43640833},
  {32'hc38d9db6, 32'h43a9e63a, 32'hc30ccd6b},
  {32'hc2917d46, 32'hc37522fa, 32'h42e6d3b3},
  {32'h43a4d44a, 32'h436397f9, 32'hc25fa628},
  {32'hc2befb36, 32'hc2445220, 32'h43c56ce3},
  {32'hc1e38e60, 32'h42a45ea4, 32'hc338ede3},
  {32'h42efb87d, 32'hc3d41f55, 32'h4426667e},
  {32'hc3e135b0, 32'hc2f973ae, 32'h42c7ca53},
  {32'hc1c372e0, 32'hc3d14203, 32'hc3b3ec1d},
  {32'hc33ffee3, 32'h42f6d52f, 32'hbff22ddc},
  {32'h41c63a78, 32'hc325f7ca, 32'h433ccdb8},
  {32'hc2d8424e, 32'hc311b9f9, 32'hc1e6658d},
  {32'h43557243, 32'h442cf4ec, 32'hc3adef19},
  {32'hc3af0ade, 32'h42daf8b0, 32'hc3ada28e},
  {32'hc31771de, 32'hc3d6a012, 32'hc39d7d52},
  {32'h43e73282, 32'h4243a2d3, 32'hc2c49807},
  {32'h427b7f87, 32'hc1a86612, 32'h42d32caf},
  {32'h428ea552, 32'hc3256d88, 32'hc4131c3a},
  {32'h432a2e03, 32'h43c93334, 32'hc3d52645},
  {32'h435ae831, 32'hc1a74ea9, 32'h4209d53d},
  {32'hc3079590, 32'h43627e21, 32'hc326194f},
  {32'hc2074d9c, 32'h432aea94, 32'h43caae84},
  {32'hc3dbc0e0, 32'h42c421e0, 32'hc3868d52},
  {32'hc3a4cfee, 32'hc0844f04, 32'h42f59584},
  {32'h437a4551, 32'h3ef30f60, 32'h42c5afab},
  {32'hc3954454, 32'hc3a4bfbd, 32'hc296c043},
  {32'h3f4fe380, 32'h43266bf2, 32'h43678f25},
  {32'h43a3bd88, 32'h4376a4c9, 32'h430d0389},
  {32'hc3045d6b, 32'h42ef608f, 32'hc3a8308b},
  {32'h4361c646, 32'h43d1622a, 32'hc3afe134},
  {32'h438aaf90, 32'h4401edb2, 32'h436d0ce9},
  {32'hc3a21436, 32'h423f39a4, 32'hc37a5265},
  {32'hc29b9aca, 32'h41b8e6c5, 32'hc2e3d29b},
  {32'h43716ad3, 32'h423bfb06, 32'h4423b2d9},
  {32'hc404005e, 32'hc3193e26, 32'h43bb3e3c},
  {32'hc25592ba, 32'h42b41e59, 32'hc31b5290},
  {32'hc35219e2, 32'hc32564ed, 32'hc331f84e},
  {32'hc3c49a7a, 32'h3ff61780, 32'hc35e211d},
  {32'hc3ecfbdb, 32'hc3aa1632, 32'h41e48b60},
  {32'h432696c4, 32'h4391ee93, 32'hc3ac0b39},
  {32'hc3b44338, 32'hc33c24da, 32'h43569f0e},
  {32'h43b3dd36, 32'hc37b5d20, 32'hc35b5ab2},
  {32'h422c8794, 32'h43f4d86c, 32'hc4530e25},
  {32'hc31dcf11, 32'hc2016e3f, 32'h42615ad9},
  {32'h431e850e, 32'hc34e9f93, 32'h42e30b9b},
  {32'h4314991d, 32'hc3e28a40, 32'hc32ee3c1},
  {32'h43aa0507, 32'hc3d0d4a7, 32'hc3224167},
  {32'h43c15355, 32'h4296ba14, 32'h42ded943},
  {32'hc04ec4ec, 32'h42e21699, 32'h4420fa2d},
  {32'hc38a657a, 32'h441b2757, 32'hc1c70a7e},
  {32'hc2439fe2, 32'h4323aabf, 32'hc36b185d},
  {32'h43e93f4d, 32'hc3161abd, 32'h431966e8},
  {32'hc2e73358, 32'hc277c982, 32'hc31f8cf3},
  {32'h43611c9d, 32'hc39120b8, 32'h44006510},
  {32'h44020522, 32'h433bb37d, 32'h43cb3021},
  {32'hc403587a, 32'h42024885, 32'hc279df31},
  {32'hc30a99da, 32'h44080ee8, 32'h430d1043},
  {32'h41d1ab64, 32'h439f6d23, 32'hc3d7e809},
  {32'h4255fe58, 32'h437ae1d0, 32'h43364650},
  {32'h4236c62c, 32'hc30f1599, 32'hc2ac6ee6},
  {32'hc3d1a383, 32'h431cc6d0, 32'h42404544},
  {32'h42c18af5, 32'h4384db56, 32'h409647e8},
  {32'h43d8bc73, 32'h4334fd1c, 32'h435d771d},
  {32'hc3835e4d, 32'hc3b67cf5, 32'h43d7a6aa},
  {32'hc25883a8, 32'h425b2980, 32'hc218aa85},
  {32'h43c08e72, 32'hc30207ae, 32'hc381e2ad},
  {32'hc3b43ee0, 32'h43e747ba, 32'h44069101},
  {32'hc0cf6646, 32'h422a8aea, 32'hc3b4579a},
  {32'h437c0fa8, 32'h43c9156c, 32'h431afafa},
  {32'hc3338d20, 32'hc38cfa4f, 32'hc3a3d6e8},
  {32'hc409d04c, 32'h4363aebd, 32'h438672ca},
  {32'h420f366e, 32'h435ad541, 32'h43c4f7c3},
  {32'h421713ce, 32'hc39c7712, 32'hc1e2f655},
  {32'hc208f376, 32'h4321d6a4, 32'hc3ccbcaa},
  {32'h4451c0ff, 32'h43897af4, 32'hc1d81a86},
  {32'hc2793766, 32'hc32cf6d0, 32'hc34911f4},
  {32'hc2908c19, 32'hc1eb23ef, 32'h42c65157},
  {32'h437b2517, 32'h433e5c22, 32'h4366f45f},
  {32'hc0983f4c, 32'h43573c90, 32'hc30aca0c},
  {32'hc33a1820, 32'h4338b4e0, 32'h426db4fe},
  {32'h43b32a61, 32'hc35b37e6, 32'h44119620},
  {32'hc33b24ae, 32'h418eb1c6, 32'hc37b0198},
  {32'h42c6700f, 32'h438be23b, 32'hc3576d26},
  {32'h412f5364, 32'h4335fd91, 32'hc29944b2},
  {32'h435de276, 32'h43449700, 32'h4380dd64},
  {32'h410eb2b0, 32'h42f2b788, 32'h43e5ea06},
  {32'h41600a18, 32'h43edab94, 32'h43473d59},
  {32'h4295373e, 32'hc2bec2ca, 32'hc2370d18},
  {32'hc307d744, 32'h4337cb4d, 32'h42d47307},
  {32'hc1a03312, 32'h4383763a, 32'hc302a81e},
  {32'hc3bfc7e5, 32'hc3682dee, 32'h42accb60},
  {32'hc383167d, 32'hc382c69a, 32'h4358d6e8},
  {32'h440bb4a2, 32'h4354f493, 32'hc3d1f505},
  {32'hc3225b8e, 32'hc2d5dce3, 32'hc3a0046a},
  {32'hc2d1fffe, 32'hc2f21f5c, 32'hc36f4221},
  {32'hc38f28c9, 32'hc1d71d6b, 32'h42106f02},
  {32'hc37c4b97, 32'h42bc4c92, 32'hc2ff8aba},
  {32'h4215a635, 32'h41cd862b, 32'hc2bb7ec0},
  {32'h4352b99e, 32'h442ea676, 32'hc34e59d3},
  {32'h43827725, 32'hc2ea1cb2, 32'h4413795d},
  {32'h43704b22, 32'h439df614, 32'hc35b7cec},
  {32'hc398f57e, 32'hc2c84dbc, 32'hc39338ad},
  {32'h42b878f6, 32'h41f14e92, 32'hc175eaf0},
  {32'hc22e3027, 32'h42afa5ae, 32'h42fa8bec},
  {32'hc1c80b50, 32'h41cfe247, 32'hc3526b7a},
  {32'h43dbeeb3, 32'hc3cd5222, 32'h43a68234},
  {32'hc34e1cf1, 32'h43211d78, 32'hc2e8288d},
  {32'h4407a300, 32'h438cf895, 32'h43983429},
  {32'hc38311e6, 32'h427ad20d, 32'hc3b322cd},
  {32'hc2e521d0, 32'hc3cb20fa, 32'hc2dc39d8},
  {32'hc13479ea, 32'hc3aeb2de, 32'hc375c1dd},
  {32'hc1ae0060, 32'hc21815e2, 32'h42dd982d},
  {32'h42271248, 32'hc2a3e859, 32'hc406f235},
  {32'h44072b20, 32'h418596b1, 32'h44021106},
  {32'h43ccf765, 32'hc226a706, 32'hc38cecd1},
  {32'hc338931d, 32'h43614daa, 32'h42908d7d},
  {32'hc32b6726, 32'h41e11d20, 32'h42902c0a},
  {32'hc273bbb5, 32'h42799480, 32'hc4143034},
  {32'h43e331c4, 32'hc2c1fd28, 32'hc3b7bbce},
  {32'hc33491b5, 32'h4107016c, 32'hc31adc55},
  {32'hc3e2d81a, 32'hc3abc70a, 32'hc422d449},
  {32'hc388268e, 32'h42fe0e66, 32'hc35dbeb1},
  {32'h4255ae50, 32'h41e256b1, 32'h42b5959d},
  {32'hc3eae506, 32'h4433b0e9, 32'hc3709b06},
  {32'h442f9efb, 32'h436004c2, 32'hc336ca55},
  {32'hc385a32e, 32'hc359865e, 32'hc37db621},
  {32'hc35a7cef, 32'hc2e74dd6, 32'h42ea6364},
  {32'h43e7e5cc, 32'hc2b49c20, 32'h42c610e6},
  {32'hc32a9b2e, 32'h4305b6b9, 32'hc3becd58},
  {32'hc3b9cfed, 32'hc3596749, 32'hc2917332},
  {32'h436e1750, 32'h42ded5df, 32'h433ca058},
  {32'h43f3ec9e, 32'h431c7d22, 32'hc3477857},
  {32'h43e4dbc1, 32'h437c4410, 32'h43ebfcd2},
  {32'h3faa1ec0, 32'h4260574e, 32'hc358626a},
  {32'hc33ceded, 32'h43036f0b, 32'h41eb3911},
  {32'h431bfa4e, 32'hc304d009, 32'hc2a658b4},
  {32'hc3b56115, 32'h435912b6, 32'hc304bde4},
  {32'hc1f526a8, 32'h435bca9e, 32'hc300ba83},
  {32'h429c22b0, 32'h439ea67e, 32'hc3a9791f},
  {32'hc3cd847b, 32'hc214caa2, 32'h430315c6},
  {32'hc2bf0c9d, 32'hc38ec8e1, 32'h4385f16d},
  {32'hc26a96a3, 32'hc104480e, 32'hc3c1f234},
  {32'hc2ba4b3e, 32'h42e95bed, 32'h439b50a6},
  {32'hc42e822c, 32'h4317af2a, 32'hc1a99e4b},
  {32'hc188c98a, 32'hc33edc0e, 32'hc3b152fb},
  {32'hc3b2f8a7, 32'h42291892, 32'hc3215ed1},
  {32'hc3dc3bee, 32'hc3361138, 32'hc3577691},
  {32'hc2ed5f46, 32'hc38e9220, 32'h43d48cf7},
  {32'h43e1598d, 32'hc182c856, 32'hc3c83edc},
  {32'h4212d0a0, 32'h4322cba6, 32'hc39249c7},
  {32'hc3a1b582, 32'hc245c61a, 32'hbe63ebe0},
  {32'hc0424948, 32'h431ec967, 32'h42b638e2},
  {32'h4400d3fe, 32'h41802849, 32'hc2fbbec9}};
