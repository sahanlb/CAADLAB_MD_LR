-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HMN0rSkqrdUmGbRI/KQDaJBxxnz6RNykBkOtmPJeD35FKFVXdlNiPBueayMMLwQxHGGSjkliU8E7
r75oAfgYqUfcAWpfnj5PE3em+s3uJbyqdIRqhmYXLP4mlHpBzBJeRQ1bf8JCVCglvA1rdErJh0P5
1zSeehK6ZZGEu9y3/cx/aG9VO0zrlZNb3dBYuwn3PY6U8Nd3LWsMFd6+QdkQJMkX3qIEDNpfFUOG
HlkezcREwFcFVZfFEFr4rF3oUx91qOEcN5EXJyc3hj9RieznrHsighJ6+ldYTNkl8jsN7c70mes1
JWUqgIR9VPnuo3z3lHvQ2rLfmp7CrRB+QRazAA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20112)
`protect data_block
/RBnXek7dJknoEcVEKF/vWQwbLxxVp6jjnPK/hJVOtvPAGTZjDqw0LqLcB+hvnvoNSKEC/97UdLm
dq67+UUNOcK3q9CZqJHYPX8OLZrDj6AIa8vbvDp+RVPkL20WbIGRHfHz0H2XhQ9AsqtC9HU0wWfh
/WZC4n5YvNEyIDs8Fw7LxU+0rt62n9AHFWvTiGElJmZoShVm4vEO2/eoRlMgJMi40kWEqxH7v/h9
NIGYCZf+fOje0jpL6nShqpSVhCOxzLqTVUhnaz6ORb4jqapUDZRhMOh3HpKsZwmMTJqM41u5IbJY
12xUdQWvEnlIUgAmlxlM2CKZ0ck5WbQ0Ti/nk+IAsSLKks1mGYCMZHsh98Sy1OWlPfOqa2hsFa6T
z5ZpMgZJHZHt/2n8DCJEPHReZht24kojsEAEnMh31l9PGvJfK0tbbdSvbzK5nR2KFVAXZjnli7ok
R7uyC86kJ3lkyF5tnlab/momyZZQIeRjld1p661z1BV8e+Oj5xHa2ln9xqJgmXDx1CBE8Xcn0Jj/
Bav3unQrBOlcgOFZB04bbJtRLM89a/ipU03YffY7DWAUwVU0t/9T3jea96NhDHxJwAzkICI9eo2m
JnIdae3d+LDHwf5l8XOYsqwiyh+KVOKLXXRUU+/LXDQ4gPfeTsnyVeEN7GdFLbm//ELpvDCyhiSr
qjPMzGj54oBAug1mNzwUyLh4GzVRQ1srbaqRYVpTA73/dWM5N50RlSaUu9AxfoODxX0LIslCDCLO
B9eRstZT9aYyHsLYLRptJGN8xiTMDqZzi8PKgzVMyw+SGFoum66gd1+u/kE4H5RwsfqjtuMHpRa4
YpJJFDE6xTKzXFH872VXUV48FxFzAw+S8d8Ma+2IvwHRRudfOUhLUc0UmTvv4/dvC6xFwVCNRO9V
+HW24T+ibdjTsWxaOVQLozbh4jw0mYaZ7BaRF29bta7AAyCb2io6pmz805ODjaBOCOqUoVv27j9/
aW9GvAErVE/bRiAdMQOmyWDWDM0Y/08LJJSXsZC4cQ4epP+LFpb5CMJTOpwUUblmqdshpB1nq3kC
0+Bgbd9X5I902+9ESOL+9rC6exvm0zfxYXyMCC6iH+aLLy/SpGnkfHmd1Xvu8olvkSq7Ee2SIl4w
0FQ+LFh7VI6w7dtZgCTPpE9y6eRZvkdF2tTUXgOweCLTz1o6ttncleDgr1nlg+PeEj0DXahfZuGd
rJzH1Z4oRmjj1JzUwCFqupJ71Duj1CtC3nMwFH2jtSgEXobOJAACCOE6jnc6oE2QSDXyN31GeFVn
lTAO73gh84NVgtcUsRIRrw+6iM1Rd7Vns2re22hnvjgSmicHj3+MUS1YtgFsYU7HR8G/ZOFAL5fc
cZbC79Zz3KQUsEwBmeZ3++dG4t0WeFa5lm5VTgFibLFSFn76tgremXMLh6UoAjhBPrypHYBnL2og
NwQuAGkg3jiVNTfJEnjJcmXT8BuqlT0WEWTNMQxYDtL+zphg2Po8hwkJePn0zky9jXc2OJJ535pv
G9kbSnymuPU1//wpXq3Vj1nhlDNcqO4jEGNu4SL6u0svP5JzrRXpY0QvZXzS0Chg/jfDMRw6J7rO
iqAlTnNI66MFiMfuMdf6/kSB5kokrm9SobJT22yc+KE4qP0zn2LxOkFHhJZMw8XoVLrilduMVvXa
Rr0y9T3d89iRWHmzK70xJ3wuztdIFPaQ5z9QPzy5IuOozA7tC216DClt6lcK/civHMfFuD0cV9bJ
T8lXc+ubLCiGoRP4T50cJR2vsE9/MJ7VdyRVbSYEG6KEP4Q4l2x8IVBxyLAOKJwPFL6MD4ddC2p+
AzKn6uw3C/gRHKCa7cLDbk9MMGW4Egd9yNmy+uYvK3VIL5I0mUa7DqwqiKJoPZY+qbpqB+CZzL2k
umUv4bDtgQ+i2aTiHw80trg5JL8mTzSlc97zBhB41cfJbLu/LqZ2nTzz2xKk7JQLjfeOqlAGFkbx
AXVGo01PbHrURr5SACOjvbgk0lY5gpirT66RGRhs8Oqf7kViqRRji8LGHj3yyS+I2ku3en6sQkbS
AGQ7VpUcTKDbtf3na0cQspJNzGIk563TjjenagTKOA9Cevhe2j9TFLEcqHmaSNeiCOgTXd6Hi3GY
tMmrTpBX74fS3nunf5kGx6zvIBvdLBntqNziz8AMEr+RDdBO5XMJM/Z2RJ79t4m+oaFMbFku4w0t
4dG4Vcmj+c1okoDBTANwlZlcUT8/V0dJGQJaI+rKM6Cbv5zTcQZ/KnUGBnith8zZOltFlOi4mDib
pKa5kyx3SrmhBLK9lBNCAVpcfIohRwCyCVaVjbSsnlqv5kXMIoC3LLvg5hW/uPwV57owVAi5olJS
bD8YybDrPXTbkf/cziSkAW3qv1PKpDxGn7AylLYVruE2b/15oZxNskZoXpJknw3KFEDDJAyIQi0/
bm+zminrU2iQ4B2FaWOa3rw+DWKrB9I0Kmfn/s2pXgQgSho1qe3HcN6zNZEUR574vvwbMjsZQEao
Yw8t3txPI2AihlYCuIBj9hBEeVqBI5xgRodpy+m90+aPrxZ9qagWr/bxFgAtwIjY1Jr0kl1DjT+v
GqegVjnctR+YfbeCZFphHr7ozuS3mf6kyz9WfxUUJEUA4IIqU0c+Y4t1JlZ/Eq6QRdPhbDnrJ+VC
uj8H62up2Vl5IRRE1MSv7m1IvhnQsPVVoMZK9cRZzn3xSC+nUXbtlKgtj1l0UwB48V7nVS8LSkaN
l5YpTQLKYCipfJEiaf6UHaLEc7+23sanGMD+wXRLVHiZ9NCBtnEPNBKPKjRXYmQAfpGP02VbjQkG
YWdnMWj1lunMpUaPoXF0IuwoPucIlL5wpAl1CjhK7h2GAnw+hHgAWDPfgxHbuMRVAuWhZhxC6GO4
sn1iLnCaKACVzCquPonpuc7qZukPyMHWHudbSDwUqRrBB8V3DEXiOK5y3YkhUkg1zz+JzVaARBRM
HGyQpht4WbWKMZa3h7q+ebJbxWoSvGeWm2U4eDoYC5tTKeKp7tdKGSubnapYvVC1vUXVVKRKj1lg
7pns5x2z5dw2cnNVNSlWJLozPNtinctnAKeN/OeXczC7jakPVqrsoJ/LgrK3jjVqBLR7O5g7s/zq
V2WcyWhSUfQmJL/g7Z/Cnes4YD8NDFdA24RsVJG0N+v6elXc2qFpORPpfYCikiWRjcrdMdySFQOD
zSAuQjRoRug+1nX6ZtbkTtr7pX3ksAl+yGh/jw/n3WjdX7rUjrrBqVW2GKWswfWf8RFjvFgys1vR
MMXXg4AFGO3hNigYlgpJ5IXIozsYKYIwaKcfs0pv0yvQh9wPhyVPcHfzgCaXHyoEamRhiCz5Kfmy
DSUrzmO7D1/93Itbxxf8DwMWU/q6Yati194d1RoD95RrcW8bgfX+jHNy3v2Sa6eiVDfZ7VJ8+WAw
91MwSc4bcN+TkHXIVA9x/xboQfvH8CsnxRzhC9olR4LBp4JadDRJiEmVIsju82M+JVOfo7c21tNN
gKrDOBCdWDNAeXUWYuy1Rc3A2Wr1Lw9xw79wBGGiDpyGCWOhZbSrSgVq1KjK6GvLeC43ktf/PvCN
pQLasNKrfd3o8kSDxFuU/FnSVquykICidFQKzgFzUhnbP8SxkKvTR4Y9sen8WE3pOc1v3ZARY+At
fkDy9E57+6Z47U4CjQ/ShRvl8ZDH/8KblCyKgGLs8+/NhxUCmyuA1DIXM8yUCss1eDIORu4fIgNX
Xhg/0zBhJHzDcD6vGA64583dJazTciLNWoZA/gVHyHILWs4sV0yzakGhhiWLUzotn1oUPaOpWmrs
1Ddh2/vCj+jHxE/JgwBBm/oKR4vBmucVH2HiZD7rZNw1s7BeVRd7OZxuyUtdxLqyo+51NT5XqJk2
12Ulm30dX8E3YTNBs0uNE/+xkPpk6Zs5amD1oSwJDZRX+yvt25PBVbIiScJbHSHn9JrAfSY982Ou
A6GtK9rJf6/G3vw6NbEczhsLiKT3LUZ2wUQzqVFYgFB8vsbhugku+HO/f8PJa5qRN/ZuFU3k7PQZ
VFJcm50S3sUeDboA0rn/ABykVa8f8xmv/Ldabo9Gq2y9CTRDOSyReUOzHgX8njS0Ub/Iwxy/mZ+8
4s5uMg3ABx1R2As2EWYTXlgEutuZ3TsFi1l5Db1zMUyIzuRWMDRm0PHzzrgALDKLQKybXyKuwS3n
e1DKxUfOkZ3dQ5dbZZzFtUuW48MnVK8iTd6ej8qHgV/mfDlTKs7Jy9Q97p4DPyhxESKXbZieN7/y
O9VJom0IGOlXQ2Pzc8gQvnwdxFLBaw3eG0zpvspxw4O6Nx7fgwlQubClQwmCQmPsxs+WvfHbHLRY
YZ2i9G6fe/ixEUgvsBuKQnykoV9oljCvk5Umr4FF763q6/aNi+NZ4Ck+IN4RBOup+B9VpVZjZa8u
Lc0/yL3Y336db+R9+s+eNndHKJ8zZmV6MTsmGDMshAJ5PsA0F3wWGBXy8TwMNFviY29mhh4uMyTs
f8eTnL6MqyUtT/o6fvmMz51pvXyqj2hBAXs9o92rO3F+jJ6Thh3yAgI+UcpCSQTn8/f7+hcf7tgB
qBnTu/dlfDlx22my6Y+En0r96AW+veik8z6aP1cxm5o9VR7nfYDxyT/SghTXMjXOGDxAZZe2itwY
mK7BIR0QqIrve20RTxsWsizWLnHswAQd0bynWaqUJyq16IKQtsS64+3JcjE7OFt8BDNigrHksv8J
hQFzYwoK6Yvb4FZbw74tQeLlA7AwCv/8D3SpRsiO3NHoyWG/9QK7mtaLCf4ogUMLeToCjbI41SDM
75rDSmCiQj3S+cIM4UXsKWKv9Qs02FYJePHGVlWGIM4lNxdjON9r3a1ACrJN88WqEY+KakayKuTK
e9coh/Po8XlAzrxrMdNcFKBYdDdwdClXHMacjiFxPbxz3WRSw992z7vYPH/wvfV1lFtGg2DJNlC3
aWjmfQblFVWbcDNt83TWbpMoqSkXHe0VMdEyQhc4LRtkOy/VSg5m7yD3KPlx3s5LjnvNiNMjplOr
XoOFdgi2nQDOZ6NbIe3tq+56WD01js0syYjgnvB6LAqk58zUfcI6GnOfh1iso+GWj9oAeo7+Gbk7
Tqxc7bbv8PGN8WmY6Q/5jkWCMi0w6s2+LHhoEMHfDDPrdproRGVID+w84e6FGP+goBFsioKANl/m
+74w8v8gMgEv5WDdVklo6g1rYzbXbP4SMBj3CYVPAZQdcAxATfHX7q6n853rTyAqe3Rz+CBUOCNa
2nbBrHqwB3safSsX1sDtkcU7qELxzdtQWhz9d9+azfZavFjsw4UH2uqlTkjmZLQCDaVswaKxS9tL
e1vOq7dQU0HgRI2yBr2H1lguPP+t2swVsUZec7IG88848c/ZnSqgYO8gRDtzjwLAiboqZU4GYit4
UT8pUEjT3M8j/qPm8ygg080FVOsDVlpmnn4vgXjxJVVeV0bvC5mgjykJqe/N2EHCceeQbBf/q4RL
56UlnS8mA4f+e7Ck2OJVXlvDp/e42V6r/tDWKmDihgncRWnD2mcUE5ghKeyTdfSftMkfiAImtl+w
velWiF7xLeI8OqDzzpSbBQ83mo26ztYYAszueAbd9GOPWgk49a6GZhIrf1oZ6HEJRVLxP/iHdeEQ
/mjueE5MiVAbcnZMffkC88yPyz93pImpbvDAU4SahubW9jQocMRQ+ccW2FKbKqhXf/eNIT0tYSE4
BdAIUHw6bIkBkkl7xb0mL1P/QQvVgcc/th04X/vYS993ScwLnSm+WXvRJZLAC49+fR/JyE5sI+WW
D3P6VG/FOrFGCAEty50IdWbg1/EdMJybM5sp9oe9gZO0IXxGo/aqtt+N1NL4VHC0dAEIvzLbg0cB
6dHUBXanJ16IMWtzNsGXAZfEDnhzdDwCgWTe+W/rUBpvs6VSxT6sKol+0/F69J98BuQ8iyKq7hNL
4ASokGJtZkVVQh7pNuHUOdjy8J8ZqaBphBGWJGKEdiXuaVX3KdO1jihFaMxIzmJJTjoQ/AKe4ZgQ
bHQpINjePUOzUZxDQLbEEbv8Y80Kjaybv16LS09wquu8I7ueB6fJb76ZjxTtD48Sb7CnR9jJGrGo
4U3qoDrcfy4ZXV51kNHymQZEU2BIjM+nY+VzRPXFhf9IdfYYIgXTOh9E3JT6UIJEpAErsriVdfyL
Ffbe4OP8xxRFaaHmPuwjWCbaS1r1MoEx2jZJjHd7Dz1M+E0TTl4cE9zGtuV8zfNvUTswfsxRR/hO
YMeTM0U0npX0/gLXZB5Bc7nqBSxVQfizTKVszQ9a5zMTsgo7YLDh5MXADs4YZAtal7RukAZjngm0
nJhZd61KsSILDVcXrTtY4cDY0FkJRPIsI6XX4oALKEQYQYA8WC8iSKtiALgBEtJgfXEt9619/ssE
KRnBzPN15U4WXGRQtQfEyElTaCuYm8Ckmoly3rL/zdUqBJ9aC1bd/ECxInWWdK/QVs4fqYAUxUD/
qH2C4s3wn0c/HEDR86E7oCGdXTwdItoosSLPqKmkjC1TmEUBaMj2jcqCdGNp6miKS2o1d6O6THsl
BvWE/daPRHf7ODSKPMuttUJdoVMG9Nni8nQJl02I5cYtWJTRoKLhlby/gOn+6qaO70n1/U4p1qXN
DYApmIIdFkeVNaZUVXSpzvEeUUcloC777UCqdlt4xlArz3qp577OLl9tru74Gop/5+QtKpIWBI33
b0ZoOj4L/6SS8xjz/2JvYdVX6L/WerAsoxWfILJNgFOXcFGmfRNObJZBXiqG7C7swlT4LdnFOHHj
C9f3yG4ebBm+k/I59kfeuo9l0RG/xsAjMjfW9oUeY59eJIljOqo8MjlwVqFY5+7DzdwUPsU9S3f2
O4T3YNzy0VsvmgrFNMYdUd7a73KpYxWkpJzT6l/+xC7eyA9SM8xcJpYmMeO2I7oh0TIUpmVE2bWK
uJ7EhDhStA21V6dNXeceN/ASl28fCAjlX+3fgxEYgk8SEZwTjmbmHc4wO5+TDnNie1KbriyZyV8u
I12AMCPmDmQOu0yxJUyqF+nKvEKqWsarE2Mzn+1jvtoTivXyywOf5Hw4ku9Jge0JCAvkeMeWvNXY
niiuEDdePgmTHfjooectCNqVe+u8XB/OUNv4hHKgJxrnglIV+aryflP3UB7BjUaeikCwCawZVl3F
Yh+bQOmlApqdV+hNcgil5NdP+Qc9OTKc1fFpqJqKIyFJYYDXL3AnlysuuGBi/XALoucz6rlYfJNq
YqUV6GdbzLS+RBHM83NCN5joNd0lWmTAwEn2PLtVJjjxmhP2e1xbmsrOz+mYmookakOvMkm+TIj/
pzlxtH2I7LfYB8tk+amYMG4jofVvBveQxLwD/gtDT9YuoXqM8ekxhYSicd4tWd/v6SskTv3Gm1xr
PiHH1ogaD62amr3MGASXOHrzAigcOjVovwQF0d7LH994OipmSj5rSOeBqQaAzaYf49TrOGzvxZA6
tzalB6OzPw9UNO8QJGlvxu2XdBoCSkybFAHJ+1SjCzBFtsnohaq4B7F0/LAY6hYYuZDhNCo3NnOo
EOqOdUzYpgutUjOXFFBTYcUE49Zb1C5RzwWeW4hFkYcNljjZT/Q+rv9wO/MUaGd9UfGWLF7HzBw7
6bHOOCVfydNJkcv5MRo4TP9F0mPlbWUB8JG2Y9Rj0zwIBNuNNIykTpYWbZE/8vFuRDX0vzf3QQU0
Q+7GY7rW3HCkoL3KY0v+GDRCFySZcc0p+ehjTOdfF01QA6MI9hto7f1XsU8XBnEBcQ6rxqxCQ7p/
E3wp161P0DzqYVB/5IBaQNImpiedmXenVuc72SdRiHaqAnFQJbGC+usHvi7/11nxBXZuHPJqDnfK
XvKSOwesowZvKCYZt+ZKGFO2OSdoRiIrCbBPUrq0yVJEHJ1I4KwsN9/ee1ktA3hqtXkvLpqiA/1b
Kiku/DzrSYVpUb6XTqQHxZ8H26UxepxNehx3o3Gvxz97orxxd4aKryAGTlVjkaEUJXrvJub59fX7
rHY67yqOlYNlcBw6gJFSOfjM3VTdnw/6RCNuMXEcPZpueBFq1kZFFGjbGpQ9e85JwCz4nsNQ208L
GYuPqlY3BEVCtj7CjaYOaCyr/qoE7FmHJEZwQeTSjzdb8WwZkxVJSFJgVjreK+kiOqIFpTh1RicV
7TZ0qz2FE8rwkFoJrTjwO9aWspkJzuPR69MFJnG19vbXgE2fT2n0zrZ1gbytSf/Ze3MlD553aMY2
ZaiPhhokIu2Dp1CXvPlXesD0BayGFByTM0JI1kduUyWtivFo+jZ3PLEuEAyGOGJWBJPW/bQILbc6
oYfqY/hZKwWIiCGMnsEganz4n7+/1llPKIUGP8l7Hdk3Kp5m8eyJjfyyS2JhthZGgsdYUH29fywp
RK1WEGxF0xUEenU5Fin11LWXlc4hkcZ/NDms2lR/nS9RXCcXGT+5IGXPncxdxxvjSVvYg7C7JssB
1uB0UjfWIJM3fSYRUs9ruf847wEeKo4CGrbjQGdvqhR4IcTXAGpEUrVwpxWIzizEvGEn+61sVChm
+lsD3gpNhF+gO145vBzkUnFxCM3y8Kdz6DOP+RaOSn9NxXGcQ5V16oOiuSvlwh8hrm3ueDTxfh64
vUsVU4WFkTg/dLIhdUCXmplaScIKKhXSkOppaFnKkgjIlR7bqEowtscsylL42qgvgB0ko3VT0Tth
ikVQQHpgPBgaZoFNfPgQnmepHoAbn3WAH9Yxjl8yhl7Xfr3JAAOCm7L4rEXRwQXD3z54LrWKbtxM
4QBeoBxn3TTwlZvohqS8zp/RJh/kMAyQqqmkXxZWpSA1WjOYNS1cKlqojKJHriSyB6S+eRxImGFX
UNz0pBwLMeIOsuIF0HrLzfpYaPS8pgfAaIt/HinPs+cPJ9q/Lvi+BVT9QDuRlq1s6XHabRe2bPIP
RN4o1bA0Pcb7wnaNz5aLmL7x6D6iSXJyMFzVoCGpjBFJu0zvXPkJn3nlVhw67ZZeXsanqFIXe3DH
1u53ArSbAt1r4DmcQIWEIGBrMVndjlIWjvEp3aPhmtsu6Iqzh5WUDrNARZDhffBUJV0RNFfD60nc
816hCr5TKkbQqpqc6qQepQpuY7n4C6nhpXQlCK4s6XtEEDg52C6A1xpLNPzja7iPYNC8XHhMQHMK
ODIpO1yKbHx9wny8xJ7cbGZRr0+jYpwasgMqALL6TfnIuRVuNV2eWNtvbbEIQptljfLFP7Og5/Nk
9+sfDAYlvf0rpbS5l9bVQJzVVGjZv9AuPc3vSx7axSWYfTXf4+d5Oup9yd89oV2dP4NtGO0vBfr5
LBpsQe2aE3LQPt/+UcALCJ+Nm4J/1oApUGOs96qc7m4UVGRjAZ3OtpFKJPSFm/gZ0rq3mHNgsAzZ
/mD8aSrvneiR30Z4FktxBZXxksa0pPGm5559MXhEYYaOLMoLRx7xZw/yrr0qOboCOsGc0zzEHHVi
4iXd40isi8iwRGBWEaYx1KFdcKvPBw+6Pyzb97A4SM1cfFZU8I8MI7k0d0QhrbneFOHeis/SxgBZ
YfCuT0WdyeRQ9MLjPdtQfZj/EXN8elc9xNwEUwpwYFtYFl2NfslUrXFsz0cH5E4ccv6W0eXD3LH/
bvM3aS7/8ylk8rER1mHT055tywMxhkAjdqb43+QGpVlXAnI0O9r1q2Qkv4nsyt77nx/OeB5uo20t
Wmmx+zdDkp6Hqk7wNNQq7sf2/Dd4CzbvA1k1QswDZAJoaIF7C2MOIgAjjkXTSmOdSUm4DXdJ/e0W
4Nd1lIBeSBqo/h5lf3Xv1Gm0ni3Wx2k1+Jt2vHoEiqQRr9yLOmJQnMPklpzxNznk1XQ/xVZJB+eu
q6WdDNqqJIZ8At6XU0Nkkh3aKEnLVQJr0xHrKCHOU0RUzUnG/k3mBuAmIELGuAZp7hMepPGoReVB
S3nNH0ynklMDyLCJp1wpm58Sz/TEOR5Exq4lAzm5uIIBtQbSr9OeXgeKiiCjc4KyqnxgeomL4Wxs
e5wnyGvFOQkjIdhHxOwlcDrnMB8phyT+34Bmdh/rmosRRXdOmWhYl3w84M770DR4IMtqzGFMBORu
qbXd3B3cI/oXDFsLba89rjnOS2yVyrx280Ka2ctN7ZiPQRUeDaTC/IFfAPVouqu4zyPZV+2XfiQr
Ssewh/ZhY0j61orIMXYLM63k1Ufb805ZhO2HksF0Wwjp4BpzunNFd9KhE6XIkOpadtJigZFeTdwl
/PGPZgXinHqxPEn15yYJiC1hXkX6s5FkF/RHPRFFLuIS/olSJHrYD9q/t1ujnqwpf/qnuCdA7Ytg
3Xp9Vbwpe1Xrd28i7Wqyyp88TZCiTRe3yF2EpvQYhT7SN0YIOChzKnsPJmUl7LHwtTny85SUXMoD
/Br2Vw0I+dTQo8YUf0ES2ohk61XYHcpDkqdRlnSfP02sp/vYZUJQNNhxrDYVs4V9/Q9gDaXqDvEJ
vAr3kcfKdqhDQACXJv4DADJMb/dGF1SJDtWK2zFc6b2Rh3VagLqV0J313dktONMAd5OkTt04Hqo7
hTDmHGENl3w/gKxa6QzcpptWKZ+5Uw5zuoXttCv0BERhKPFgNyVQea5kmVcQX3/9R4E1jZ9CQ53E
SD4CKOZP5frMkQu4IzSBp26auepjxw3qWOYx5GszF3MqOhsIkUhiDyJmswBXWZi6jWh7jRg2ceZk
lur7Ybci+axk9pPKkWgGnZis6aRm7tUfLiVGWunJlFyJ9P7JL1l+iZZHSC5sZsw40j4ZJKGwyut4
nBRoKrAQW8maAUvD5h0Te8HDtJrg/6Od7xDu59EppRSfdIoC9dkVDtLx+ZRijXbSQXn5d3Pr7/7E
6yLZARfptP0lC5yQ5xgGIuhaQTrMK+/y6vf3uZUBtV7pIdbTuHHNoTqL9rNOH/4K6i5HYYWL4wz/
y9u2ccfZYbWLiR/JKxjEJPSvjOHbJY/sEKYpSHmjCgJQRX5fPPKExml3JcUtX4SRv/ey/+V31QYJ
Gcj3hgUlpA9OUWrNj4SXpzW4ras+AyuYK2noSXx0A+i1ndyScTbICiYCRdA7dxwJ/fnaI5HJq4nS
73j0bwAW7ZCU+eZgE+I/JyQ0xiuSTLAQbZHvtKkOE2q0W+Iiq491eTwMEZIUHhzyYS2wK+jMQPIO
kaxqI3VaPwKH6rNWpsS/AFKb/gONz2RAjpB7IDviMtvT67nZsplu1QqPiL+ciVItBytV7QLeHiTR
+3NBUekvCrMuHCcJZu4XMYEWEQ74wGPm9+o+oFVs95H48/204gsEpDBlY8rsV0UnnLVHX47PYNyh
/aA60HCH91fFxbUTGV99rU69EZKOjDi351sX3X0fo5PfYwoufF31a9piiBJCYm609hDlDkrbYt0V
l0V9V8Agy1eLgIggZTye/zMdEwkpng4A3jddxOb71X1PfEf41dvRgF8t/yx8l/R7fLQWyz5v+HS8
se0Dip4N5+xN+95aKvFPPCDW7gxvLykdPfCW9nHhL9MiepnqAILSfzuzNFSvGUhyljr9WIKMZ0C4
YH4GW82vTdIvgG+5mSYUU+r78TL2j7nxJYrFkewmGlrkeZBIJPDKARejqe6Zd8c9hciiMt/FVSIe
HdyHtJC2adBtOVCkk9UAWf3/b6Tf5oBE+h3C6x5jatk+XUcwnvywV+hgMMOj7uMA7ws4gY0xP3CT
fL7ulPdTEBxEV36183njnpmK8Gf7puC2o+41NyFXEAFBgX3bsH/jZpNH7SddoMJDofs3E910dOW1
yKWqkIt48ciiDsuhftVM4k8FewmyYUNYWdyH/GbmxETf8CE3HIWDIzZcfoQhjMEup3SAiXzx+E+P
UDPdWwRqxAYQwT/lgSt0ZyTX8iglLbw3Hy/LxuH1iAGmreXOP9wnhviE926VrZMes3LL1lD+TWMn
dQMDXA1cSsTKMA/4Wl5tGfmt537TQkHdkyo3VxPlEbRScOb8F9b0Tm6v9k10y9yBskbuA1GbxuJS
z1KKjI3+z0sb8cydiL8IoWwo51KYEPGmsWPQnR5vSlm2g+aHckJGee4FJ3iHVRpM0WQ0j+hSuRZ4
fMGoPB6kCf2VlrHmXLKNCblil2F+RAqPmS2M6QqOIIiMHoNVSAvxIp5RPpC/TvsHvjoqsHMx8b9M
ki31r7x7PjHdPuWSUZtvrvrsxt0YMny/tlCvJ2zEh8Fz68HTlUQszl3OurK95AXMC7LzyQKKHbcX
9MAQIbnhTuKdzjzC1r2VYbFuljvq9JMIP52DEqjpqDQH+VvkudOUw5ekFbZmD1nqD4RspjoH71H+
kH0xZCT1V/m+EOeTILVUpzWnqn/U/nEZz/c1WV0dswJHdEoCRVn45PkTn0LL4loIvPL6UMVKpSim
wuYlDAgrtDXHDapq1tth2al6e1yBh0etjpm9XhmQzNjv7pu22tKPvCfF/OXDTLZSesyvXrMgBSof
8KeAEXs9LyQYqhTH53QEI+cVmt9to99V8HaM3fGGskBe96xaR5S/OAUkp7iItmr0MXFCBKkPveDS
+3NRhR3gBi5GorHWzsWeSV1mnn4fyyCtro/VGizfYPjUwLRyGZb9Jg/MlWuBm6unlF/giaUFikEG
1xgOybO6nAsfcx1uiuJzxbESCKa09u8QiEdWQHkMYfggA8g29hDl58Q8WBsO8ShcYQiohfeHKCQ0
f+Bot/A/MLr4im+kScQ+ueaEXBwuAI7l612IbTw+WWByq4PmsbqiQOFFkOhpzKpkifUUY2Tx+/hQ
PXSxn+DXBTWSXiyDWLrRvJqucqAUgr07CfZ90enQGeeZJV5PCMmd2bSv89DSMq3JpalYgHt4Ya6T
uulqjVoTSo8KCOAJtzPd3xyZQiAX9PsQX1QoIPYztR18XpcjS0RQEpODZWYgOUXup3CPaSXhvCo2
cmRIGVfIam19D3aMclDDKhgcZDm6PJhMhLc15M9YdU/7x82OOlaF5KVBmejnFdh61IVzh3b86c9v
NNg5+60KImSQdzNrQx84J3OoMZc0TTfa3L4yxB+tzVBnZP18SepiJsDH/D5xHAriQlXXBt9T+cI/
btAAG0p+/pWpHF1clouiCET+g3pwd40sEKadahO6ugXKggTtI0AXKeOgyzA7+HZpMf+bGwu8u9B1
k9JvTBXWeMhaGEWac3yEjy0uK19ZWYhAgQrrtBDQ8xKelCtl3POuSglB0UlqmogXLNmJtP8V8FB5
lVxcafoW+jpymYOu0w0kbHzfFJ+FfCXRBeiQtTFrpDRLQXfrPc+eWHD++Bo56IXGdDvWTssxjEq4
TqD0uSFR47FWRPbrWaXMVhg4g23DlSdL5ZWuOGWYK8LNmhgW2QRlDc/fSE4UbIgbl4cS/P09nCvv
EkodmYcVbYxtJEwbuKJF9k/OON/15UOi5ituhZfftRracGL/doKnz2T40NLpdcbyln4T250Z0Sxu
jRN31Rh90amiK0S76b1EIjY5o4jDnuANalL+QQ56SPBV+54GvN6BuSzjlZXJthpGLsGBE1CmZzLw
eVjWRAqLCLmJnwaha/vPJjx5TCx2LJnMjuTX1ywKX47EYg/2/fwjxNY47Ky1h5Xoi4GtHAqo0ZcH
dpany+umBRhgGyERZkISBHQNRND0nzyoe6f3wL7xgJGG/VGHDtqeSDfLj3fTyC+dvsFfSa7zDgXi
PXXFvAJlORcoh+8Ow3YCSdPAkpn2NrF91aHQVfaGwjH+xYtHnFb9c1dX9IxrWmGS/wTRfZBYFS+z
L+d7qI7yufApQ8n5vDKJyvo2e7tmLUo8d20tHjds7kKWODNSc2KGIewdf4xthroJxvnkxXmLMNle
77iDQL8GWyVuEQSchsTVzyBK7ahzcv0pvkAvawuWN4DhCBzjkdcBpwfDMtRhyUL64Rh8xZTPLf2g
NfUt4bHhiNpfSmklQ9UqC8i4GKBA2zzIgTqV8gTDlZLvB8JSRQgI9zLPB4N/fEs68DIGuMmqg9IQ
BGB2cJzLhKUPT2UBU/q9dlzi2Z8amo3WBPSl7eFZWvqGEpH4RI6t4se9AK2I8UCdokYlvwFYfn44
QqWD9meTI7B/yBPzgmxptTW/1uIIZ/tzzhguUVsURwYpFAyP8+YHX6n6oMZA/i4KMz1hx2kPyQHi
sYd0/zO/w+PxFdWLfIemqMbW6NovFb+scuFm2HVldpDSLfiMEXZRSUSoAAwpcTppdoEZS9Afy2ne
FNho7sX3eI8djcBPzChq2eajLdOSXXzhU35fLd857pXc9TsAnGPWdgp5zDrKltMfiwn0ckFIC2vN
z7J6G7gpTBuPgnQ3G/361bZk2nLdscA+1mmmZBI1ElFvYQ76TtJo+yNf+QGou+NWr5iKP6TQ0x6r
RdiwFnX6N3buAHU/I0b3Y6sJde74fa2qMuu3lxLQUfBY8ypA8Sn7aRigyVaJBFgR1epu5px6j2kv
xdgx5WTvSrLPknxwP2ADF83Zeiv4JwPMPKHVFh0k9bEUIgNY7r26YyS3zTlmF45SfC5Vp23GnepZ
9Ja90KoFH3pqgYtaZKw4jl3g25M+Zn1APXXUSP/qc3J7AV6a7EXfxK6NxQbcR3relriZ5uYGb0XA
/ZQlnrC1dGh9K8Q0xw/s+3SAXHinvK6XPrGRupHrEwdju+l9VvvWSsBkQRPFFNDlQ8gscbOErr0J
YA1P7EGnKriNfhcaQGOJoGvtRzBtfTe1OWmnbwqVY6kBnvz2hU/1KcLRQEzfqHMYd0WctyhVycJT
89RAcxAC2I15bEwswJTIzp07alpgHldOOdVj/gAc2Go1aWxbf13cCdgKL1dQS9g10CzYuo8TLGMT
hQJTGV9HTxRqd1zf/eLr8k7nG/QxmVA9/MPud5nijzBgcVtsnZXZSyQ/Y/wW+omjYWp7aSvOWi/A
4XP0XRqX8CxevzRHu6plsZWhr0WM1h3CBAuF1aO6VXNtYcIUZjHTOjJjq8FWd75EU8+cEAS6CuE2
xC2lioj7/6i3tBvvi1VFs4I3uCzshyauxOCfXk06aRZ8IZTd0UzSySjNtXIzF0GTjHNob9oxSq8x
pXIqSdKz4Idh8LLLu4EoyVWOjOZi5NLMdHcmCIWQz8svxijl09CsBL81gcx4JnTKIzQNSVtIM3VE
/ifNDd9TRWZrwsdqkbTZ7lhNiZjcoQ6zwAVnTw3nANQPmwG/AOhWIY5wRFzZFzZpPipRO5mXXIsC
nGcqkiSWQHfTBuhd3+DX5KJtY0CledGdT6Xe3EmOyQV1rZ72L5P4Ommw+Y6Y/8f8UUdQFMWuoeS3
4+JwFajCBKDsaqM70z5QNwmmE2R93hOyQvmaMHmARgb12Dh2ZN6/CYULXt6iuHHoavN2srH0I5qQ
67mnbtqdm+u3Zjzwp8KSy5gwTmpUDCbwc6w4FkKTWrCfL1br5a4j7npqxJ17vjYx0I3OQPWj6tcc
V2Uw4RlDZyeyi6kLyANBsqHlR1sN4x7lzs7EzeO6LcS89jECHcScu3BxIwru0SKBzJ7kOAyHg9A2
IgBqlyv2j/fy37+pB2MZmKQ9rJ7KGu02EuFdiVyo8Ma4eRAX2ZPlDR57+NpEddKkwJX4gTxtYvs2
DwYbgOvinXL2buXY+h83I0GgjuvbLeQ7pNN/LnBOGHCkNO3/++DNL2gC2x8OmH3Gj8vn9JGCxDsu
lnG4ahBwUhheupmOTI3MMWE7CT4XdueBq2WW9VeB0+pr9sj9uJecQPfON82qyjJZ7NhhlQmxIncU
hdVyChWbxXWUIojnzO8S7LxYh3CqNdg17JUDM/X6Tr7Mt9jyvjqbWMAoPprR1kSvUCZcN9tYPDZ/
KvIPJxp5zijnQL+DAW3HFmE91GpmyTHrHBZR+g674kdSzvecVqOrta9bNKVACH1I/SIyLXa7oBL8
BvmBYfuhYTZsI3c9OgEtrHYVQ0cTHSSxWDRscQfF3pgdJ5D8NrPL4601VWCBTFmfSulbpmW92XNC
23uVSQL0msp0gdIoH1/0atJ3CvsVMEflhw0xEYDhHscIpDbVCkmUvRrAZrzfK8UUmlt/qoWcTtcp
DTZ6zK1CrY572hBmZjvk60SA2ZaT85ijKRpwZvzGEAuQPFxggRO/s86RRXWGOhLlg4tzgZoQbNhJ
s03uJi1mHG7Egfzb4XnwK22XblgtLUnHKDW8MwKohfSYT9UgcjWpQo+alGBs/HLUEXPF8ZuYhaXc
aSCw5PeR8Gm3CDP8Yn/Js9pCLjWUR+d6Wud7SVHveqYLMRSDln+trRyc3mViylFhjvqG/usShN6r
UDvJ3KUxiBKhGcjJw8RhvfaDQIjsjcu/IHscQyKTKGLV2e6X0K+acc2Ld7lC+tHegH3gESPWAVNi
EtstxmpIzkQgo9Q9I/IOxeOL2/0uieU2tv8iFlGvdyLqy402m8RihRG3YVr7LDD2vbJ7fZUQutLO
GYzAfkCChXgHYh4DA2G0tY8+F1/04v6vOW/gD+p9Xohpim83gxGwutTnWLFB2c3BhCeLqRcrXuw5
b0KR6FoA9Awu11KFSJ8CjaHJ1gArL4ssfJ+g2gFhQ659ezK6QeYDEHsMCQOTJhsTG19fcuUrxK06
3zbU9P0pP5iakfRBS3mrnjxBBzgrFeSMVS/KtwG4h+tz4IG/dL1r/hMngy3gYfvWqp2+VFSr56Q/
tkCneFE2HzA951ILGFSsaWHDPZU5h7Yv5tk2ibd1IW8yvusvtydk2YAD6NVqEwwkafEFwQc6eGE3
9mhJZaZtl7+97RDvSK4j0xrx/90dEBjOkSdj9m7JUoKClvSHJ1unrFo5PdLwWp7lgJt8R8z6FG4I
066yzeJyPNDq36qeBk1fdAqTX1ryq7rnNgWMVLmme0TSF5awQlbJu7+kEp2Pt+S0R4cQx43+pVKH
VjCNZ0MEV4nEkzGmYptIiaNypMO0pVpoYMX9VCkyeC2E9vBGt7puxidVc177/EZ6UJY0/OGj+T5c
SMUeB272fOU9dj7Gi+IVWX8kyRwvGZRSmXCyaSE2YDOjqGRiqgELY9QNLNBKfMQkQymcuSST2Ac8
7vltTZR5GaEAJ6xfu/cp/TrV6OIz8wqqJEW2y2O8EwMgOMNtnFgnMeJm2SPVLLMV28B8EXTFm5jn
NpcMDRe3/ggcpWN9ONA8zvRKfgBFb+sEehFDm1EeCyVALLdmOOXGtjLHJMZ68MciQymx/BggqKPk
rIiSs1YdJPUQYSgDL/bL+oKZEx42/K9KwnydNU5MgKqGnaj+PCZ6+zgVdQ6InO53d9lbiQbvl5yE
DJZF0ArdOSwUSByYOoI8jOv5tqdB7kOMd0SuLTvpEWJiIeLI8MrcCPX78tqTqqAR6twFTv49oywD
dIhv214d+rKOvt5JA5PwhYrXm7TlONAm+tb7TXKR5blOEj1d39wOB0AuQpdYr+qHamZvKnztAhYW
e/EVzCJu9meBN91ju5wXZbxbh+ZztYF6RmHrtkVC2T9FYWl2vP2lAO/6yD+bFugaipUNE5hs4LA2
0MAdrBz9bv+jEm82ulwoGM5mMT4uHFtrg5DHwp1VsTVoUhuTfIbpN06Pi5x2FtfxuTyK861UXHYW
w+TTT+l3rjkh21SVeP5eh4l2Tk51BHAUr5YQdmBXOhLxoCZV5PO0ozQ3qGiDEk9MthE3uX0qvIBt
Wnrh6J9H3W6DvycokR8K50NidcwITGCvgcox+jKmMjkdu7mYNLImmiYnIWZ74LChRWRt1FIVqt5v
8x4y5RCzTONHHeNU+p6PCmbfi19GGofSiK7Fww7WNNZfm2+YCfJCBmfHC2VWjjGMnzizT5iv9+xD
LnUymwmgvz6Bm+rH3SaEHbtHpF3V8wunObbhZzN12KY4p9wkRAi6O9jrCOJBIbsg2/Z+hufnmUoc
IqzPT5pfCvERGfOeojLMv4kyfDUY7WBQbEOaq+hMnGASFm1D731nlQNhvYyjhAzxL0RDTpuYfhyy
AuzSJdhQxUFBDXSOtUjARLTxxYooEnbimrhIeat+g/F8smSgAO+2RsoRMTfDDKi7TM4KKXxMLpuv
7krOslhfPw5zpN99Pr4C0w4dPvi2gaMpI8LsGiOKe6JBAwFTTaUy4qxyTW7XAaaGWbCtu/54ucLb
SevhgQpKapfzmWEOl/P5Whvd55hLdHPMKLnLBA49EPGjah9eiqIWQfnU1/pD18Gxw/rOh5qMkIKk
j7Fc+KVVvIfK/aRb1fZkLvrAh5J/T7kqCpDPSM+uqEK/r+K1aXtYlNoF4VfFZPfaUPRk+o4CZdyP
RBhchQTmLZi1h1M3DvV5FoL/kg8pGvmk9MKMfyDrJdzczI9emQCewboZFbK1xiXT+G+g2ZEOfg92
gnkOXpDCIwdcvNnJex/jHoDLSJKokmJgVTBmXRLjqEiQ+8JBF2K7Hj2fNisq5FSVjuNUAza8dOmU
C2Y3RSLGhxpn5hJYe/nITj2SQj0/GKkdNOdF97hdJWaKvAIX3zX2UnQTPfIiq4OaON0dLArF4Hgb
bT+59y74dF73UFka3Oa3gcKQzqtv0hce+Z3kNsH/3ZYCYYKb8zX/CMhy+IlOA1F0NgaIqQCXux13
lrrDB78kFpRpshnKgUYUntMExMTNZn7R4izNnN0yWvifPBwVGkh+rOySj+iW+62GDFUe24jbPC7F
iHuycsLWgZMd6OizEgspY09HgI4NxO/U3AiVGHKibBh/PqNcXQNMkTy1mN7npqx+Wj+JuXyGE4gw
Ag7I2/LtIZUOSI/tOofyLisdRynGwrTD1rQ7LeZOTre4sux39fzBWGpXLNBOY0rDUZkb4ttBqqr7
7yl0fkff5vk4hm7t/9figw92+BjG5pU/Zk7icC498P8c9WV7ciV4uEdMzGP38rwjKEv0PCfV+db+
rdq+M4CqP+YAeEo8MiF3rSeR+ndvT0mJrSxTBpR83P5XHRNU0UESgKFn14I/dQoRb3my6e2iRsTW
cuJPlNXWxqk05+741DhvDCQk8nsZmJH1Ilzc5GR4OvoyU7PbbfOd3QXxzmpTEcM/U/2nhQsGFeET
hNaUmakqO74PcFaW9v6lCoUprCMwg1EUHsiV3hcdVfkhm/Mp0bsMYK/n9wWAIddSfVR9H+Rtyt72
5VerStZs4JOQU8uz+l0pd358ddBNOr3ZGp039PcFR0SCrAMHx0x1izEDGB3rsO4yslO3sihVuu8O
lVtD3AbVTEfpnPKLv2JdY5iqX97NZIMTLEiIVav+70Glrrc8wnyq3RH2akRqYPWMyVYsEbYrTIop
ZzzIqt+RfPd0dluGFBB1746SJIwHv3ptzPJBOxj0hMK6RWUJfkCv/UsOgbxOlxR5QPZT48koHkLR
UvfkFQHcYlHqiqE5aQiW2pSp5ME7iz1wSJ/E0pCy7AZ+ytxLlHPXvucZl+ioTdfkM+u+kdBQvDnZ
0M8WJbk1OssCvddxevUsWrzXDNtKlxnsOkzyuaUUt1AJEaRksdQGphIChc8wCU/oGAgbpMaRn/9p
smqKscouazxuaqSUIWQyHh3cc2STBPki0Ukh+84Qe34DlVue3TvfmY3BoaEE+GrzAE9Ic6ALVdzv
hxcAWxXW3Tn6R9eP2KIGrHWH25X+dxg+zdBxi2vctEc7D6DSX0fwbZTR+rhWXj5BxDB94IQPD4MJ
XA3y4W3mNS388jCQ3/mD9O40ZKlfp3jH1w3DxXj6Ku9nZ231RHWR9WNmQsR16T6zg7mL6F0zrUJX
31kt6xsz47JJUbDUyHdLvC1VKGOg7XXB8CKw5On9z5dvZ+8WJrUDOzOSSDY3EOnoDdRZRBzVHxEu
BCNw01OWcNozYN0d8bNFDPyOZkN0C7kg8NL39YFLKekdtThMTtmCm9mT20SyXa7iDYm1vXo5rknp
Tlqq/QkuWCyzp75VPJlxUUlOsoWuKYIiw8wUkBfPtuRrd84czI9VLxcVFePMBiRnbVbLRly4Y83t
ii1+krOnXZXcysA7BMX5xWyW7jKo5kuHMAQLOOY3gTm4H+PxqN0CVPiDENizXjgK/w5wApfk8UpW
vC+LA9WL414Py2f8sk3asS59EF77q4+wDwTVPZydUD5Yz1CRtYrJFJTYwbuDlco2x6YpDM0IP8m9
6LwrRenibdGTnK2Z4ITfVeJP1k4c+fwODdmJ8U/WOioi+vXGK61ONn9IBDelYxyy2pzKKXqLJ0++
9095hZVudnpnKHb2LWNA6L3Zseuin25DetoQej1jDqoUV/1ifKVzsof+VPMm7a/7G8oc4n/b7gUo
9Siv06o1H01j4iS8VFyLG4VMvisAVjLiYfjiSkjSfzFFq3xi1JJKqj+wNcxFrJhPDnpNFlhyXLSa
EjPP7ylB/R1j9/10OV9Ca69HnJlJZzZZEOsnZTjkde4mXL3/UpRXgVpUffqgtnLKYbDSEFNUOp7Q
gpKMn79Qf7jFpl0A35r0uZQ0DVWs9oJohL0Km4atfHRIGlDM9V3KNiVibt0Nf1fu5ujp6pcXrwL6
40slsnPxi2Hbn45IyNz9qKcK64EevbnXmCNbrY6AdrlpjZzBmmIN7mDnvmKGCi8+KwNK6YZ2N+p4
W8Z6iTq12Iq1Ir+5OX25ydBQxGuE9by4LiSmuWo3/+d7w50uzeT4B++LwMaD/FGhouf54bXMFwcP
CEeXVnWDKjDNieW8/oELJ+ZBpqBScAF2FhyG+VANgftNPGj3Ganzvzzf+b3r9eyURhI4nXEFp1OA
hI6dY2ShnDhZ83bUk27rHWtrn/NCePsJycC0HT/Xdl2IKXkOLkpz29U0rh6KjmffYJwZB4h0Uukk
x1UzOr98LLqNyaTszagyJUKoEMrWYcIBXTDCXWk4zGrauaRauX0rnWBfM1aA2pvqdJ391ccPdMFy
x5VXLr4OGemTK8nt1CzdRx7wfE4yKS04RR1NE8+SdBku+jgPj7sVlEgJz4OU3baJ/U3J4Vgq3Y/W
HN6ykCiHCw1LzhE8Ha6ZksRWI815ZBKzOXWGtWRroNxWgPQIb61qf4G9wAtFOmqYycU7UanIohzu
4MwKZ9B9kbAYqZVj0vqlMYaEIOEBRoNSEbD2/TrVGlSpZuqRWk23167F2hYmYf0Pk+6u+zQ1+s26
7knN6k+A62rxsQJHL2copZxt/pvdZOqvkakQArXeukB7RH419Wk9t600RhVJSOW5YtODCoUsGa+4
3regHwpjadyDScPffE5LbcsJW1bPVNlpnWY9gsWzF5G7mjEj7EELeP4WmuWSsx8tEtIDRHMA3nZT
hodMjdUX1ygPSU6ATx9g6z5htujax6ZfsMGJXa9dpw9Yb4tgw3hh6mL6/N3S4bexorQT7pNwaehc
ZXVpxtTyfRMF2Z53xa18u4xrQ4yKLEWVIE5RJ64hCh6zmHnedmrWosfKH8q+YMViGpC6Uq1HKtJQ
/L8XMm/Wmgt5ZFxQSGoSWLbmFo/aLSJVWsE0rVB7hTudisHF+6AzovGZM4qtKeAB6ZimEzCLmd9w
7ljw917c61jBHu82BceonOGmYSwK93yldOtq/swV0xRQlKPcqdry7gvxzZeqs58NfUWTgSu0KKie
D2YEdpz7qwiubBQ9Egjo9FLPuxkRoPHSjIOmBkV41Bg6r2AiUFTqhf9/holpOv3fEQM443QVnHh/
SS4ipWA3BGUY9ONXVrBm83VwVkV0OrogzekqHI6T89Aj95olttRMN7fRHgSMe3JZNpRaB/OdWGsa
xsG6FCCeG9unxRyaalyVWfFl8wVhwy8igu96Rq1eNeiUAC4SoPJsYeH97nfVIquGutzt60mf2Cuy
N90TfMASDyyzZwZrQXOwIn7szQ/4AfdAn9USkaXYChpVpbZ5C32EJnfvUIiZUXpU5dnKfr/L8DeN
b4cCtb/FKOCPWAajYl4hXdaDVZ6UoSD6kEcDEE9Kkk8tV45SkeWpHm9SeGSLwlNE5BYMhs+zK6+M
yZNPoKDZ87+8QAQo6ZrTdoDvffXgApzrMKMT1qfCZ/45iK3Iwt99y+EVksZz5xrd0mSN8568JPcu
sVUB13FUxnpQHHYyqAnkn48TAMlvvSJ4ja9ODvqEq4bekFec+KyDmpi+/nSK6S4MHW12M8JnjJ+y
217YbUeq0zSSLO1nJgjXKKbTcllZDIuc1NtgBgQqfoCveIZgWxbjXpnYtnBh2QfLvbgxtYCiY7C6
kJKbTORlR+LMH41yaQOMEH/Y78jyBOr3BsM7CYBeSncpSZaheGqt99VEf3i6CfFeNQvntUk6x+44
UOLG9XBAkCIY4me/MuFgRXuNqY0dBAKfc2EK1+OyU1+qo0P8fpWnu7THyPWOjXubAwv5nsaD+3R9
tZAURZTBdS3wFN4x7kweVKx46Wa+7LveGmOEvt+U9C9DRAirgb0BQdN2tlIezffPvgPZf435u8Yi
KNRE8fRRp2x2oSF5iEUnWeVipvZWgpUdNaJ/nAIcI9XgNq2cNOIi4HW4NLlDsAH9SR43h1xe46wR
Jb3Hpcgbe83NgIsJq9VcrsoDes+u+2WgJIBGv+puzxhSNf3BY+AXPJQ46SDitebCxlS4vJUdm1T+
XlBmkYHpqTk5mC6fK3bBcokr8dBb4xpaijArteDf/Xo0GMoGo7m2YvpOgTXi5juh+cueqgX62dNS
JUijlz4KWhyZ9KoSv+0al8wKafbd4LjPtURMaMLbeIenQMn5o+82FoD7Tk2tfmVWnUum9Tcisfs6
/tZxEiME7WuKfLOhXi0PVv0t1rG/mrFGIRzlbZDi+Lv74Cg5AdeeC0A6bj8Xf55HqY2+nUQL3nOv
5qNOv5JPnVuNFprufZ2hnwuzQ/gMWUM5TwSfgvr7ij+qiVuFAnpOmrNywYgQIMNjRqdHEDaHztTs
k90uJhuhQE+cQU7tcT10HQStDs8Ns1mRanV2o0+QBIB/jbMzaduy8etLoaK31yffF6pYuTRaKJKd
8FvY4EVwaWSHlRnnFl23961kATwGBmAGmg8x97MaHYYohYQTYEDSSRKVemOIfgjj4zHX/4lfbz5x
jDdcg8CVKsYCySmXoyJFNyU9aFdl2PtfiR1z1iwikzkJ+lbfQA31fqgTgBUYfg/iYyUefIJPfQ6E
XJoQT4G0mffWmyx8PjN+yXrl+FrwGPyYV9oqW+6OptiXOf9oVoJ0iNss28kE6I6shvPNJGvXGYsX
EsaU53KFFTCbPE1Po+IUU7QffSLQDvJwtYni7FAtC3N+H2esUfN7b8w85uDWtsDU8AEhrQjzx4jQ
YKijl1Igy+iJSCTN1yyGHwzCZjtQYalTjCL47Ieijj8e2BwIoVvwW3GLvmoZkz7dY7unJ+w1APFI
rOSzkwpYm+R4iPEaTDmRq583gnAH2EZ4y2pP1ZQDAx/iapwC1DHQYUljHR/ANd6/P9ueIT5Ci2PK
aBMu7c8JccA9BetoE5/K0YW0MwiC+tWymHcN9Yyxp+gTRc0FreS9p3nGITUp/U3V+lvmlD+jKSNV
VzO9c333fSAjdM+ZwXyaO5Ql0H28D6WWzwFk+beSy6ymFDQyypviKKWXbEF3mtm/Yt8PflvhY5eZ
81mBD6/6T44kls5Iq0zXgZToQ5SgU1v26TAoeMbkPsvCVhSY4v3lkClCzSluQvbniwwd11dz9Vlj
tzqR2LwQRXG1QG/GdxbvfCvY6KkNUHQzWqxFxfiulMJrpNQYS3oAieUhhRyKClspQMcloRhsur3r
2GjmSl3nTTzIQmi1ePqS5AEiK6fsQ26Zu8VquKc1Ja/H8q3vkZG79H+aB0dsgl40GP4hp+8arOE+
aRNffqVDDA2wK9yqaPqVGuvJeX/xkDvudavJfMGma0uaxGixGaBzOGYcbDt8zZHsJU77ZmKS67kV
WZabg+Zzk9E9B58oWvbHvKn5vc/tIQbXLqsU5/XQ+T04WdkRv54zxiqZml+8wO1/+6ItLxJqzl4E
9/SNQK+5fKR1jQztCrwk1HqZTKVpjhuUeyeb4TOF1XGfiilb4OqQMY3iJA+RQIyIGaDfjyn1YPvN
RMnJxStY71haCPC5UAmAxb6kDOlBTJz/sqJYtIj9V7l1SPHAUVALNgDbL00oTM+wbU8scBV0B0/z
G+ukL20Oz+5nCus6EUiIsFCDYYcOTM0C2r/+qgEcFIMBtJW+MNBPZXNpxfl4pCdNWWtXjGgZq/aY
hC+Yz3sa/UUgB1290v14Ri7ZJoEJS1WJaYMXyuK3pZx80tI+3bh3B5hnsGNjRAhBmN7H0FQa9oUf
jBUeDYPWZnFMk0lxbO6YashWSlp0OICFANn/I4lnKlhqqTVZxJzRqFJ0HQTNgPeFAGgaEYlCh0bX
n+leEeJ+2W2HLeITAVmDvMZnI8987cBuKyQRIaGoDVvm9HaOxk8PEsS+IW7e4CTgQ2C+e27Nlg0W
9DuFr3J7tfijM33+44hNDzrwbHSICPPJU1ir6prGqKIpkqH06jR/aClyRzop3ewABOeQU1GzWILT
1B+TRWafn6W+mQu4ZYNOvQxRrvfBBe8AoEt24PV8HNCUaKjPTUJbicnlAjoEKgDiq/OC3bKmmTpX
ehIDNOjrCQ3OYMebZ7q5gbhQ55/CPnPSULBL5ycOWw5kNQasVoFHm4U+ETNI/UP+EOPhNyeG+4Fn
sU/81VgxKtmiJXFMBjqEtya1eP7p9IiAJNM67V3u7IfVlrySq9nE/1VgrNYgLzSW8eZL/Ca8sQxB
w2mL0QPDIidAky5kKLoaXxblYwZdlOXWwD91SfBqR1Hiy0JjJJ8OYmgulcLhbAoAd8JSk51U/75n
0+SuZVkpIerruE8ELjAJoo0ve3TRUdufesqWoN4BbR2NFmKyqxx08jaRWLtKob6+SP4cFUajqfk3
1Ro0h1ZNBji99+4ARw+ZWBnDs0VnbBKr8kVklSrklIQlDSLRH1T3A6+I8gJzgg1Gw6EHNp7aB3bE
xhiOLsO5Uy94KeBZg6D/y1PBQDLV+9eMk4XySGPWvghaFY6ndADLik76jqNd+T5I9LooJCESD0Bs
VxIHpoFgmdA07xBV7RL/TGFtnrHHI7X7coOe3R85Gvr/3eDMZtfNCwc0HYmlscivmQlqFfM1a38b
aBhrZbgOY9qGX+ruI8wO5biH6DnkQ7BzCLBnAtirrGnIwbLyNonJRP36Aj573eWuRP/CJrYQzcoZ
1a3n283UtIJAW2DK4Q5KEBpMyZcR4YW9FCMImI3eyvgJtx9ks/RJL0dX7jjt1kuETfF51sGQKMgA
ULeqEc6LWdiGpJeCitk65ULTVntCF46tb74tKFp0TleL0sZxtdeXBMxUD4SDJszXavwxOMkEkVxH
1wO9lTUcH+/daeGEFsf7vyoq3v/7d7i4ccCBuUxeI1l7vUiwzkgKpWzVcZN/VRE++wyvNFxjtcwD
Htkgi+4H0UsSLOCMCOyeCAYrsHk1zTeWEYHLbpUDMs845hUFucQ8ddMd4jVD29xvTwtCNxdU+GIm
cTo8ONAqTwEtvTUhrFKHYxCwrVGhdonmwnAAvpXpAGaNDd4b0zv3QaXPxkvJlkRFMYrCiKrvjeq3
MkpQ/ei6GLhNmXbMyRwuyKtsIVacGAzhV3ptSfSFQPmBbl8rLhVphLOs8hk9SH+pLJ1C4Mpevolx
DP8v650HQGeXqsQZKLDWBF0/Sktk7WmJbmeW55lfg4BNFIwXZWqO0QDsQUOfG1FxBVkpYDWdukkm
AoUOv8DAkQSHbXktm5WwG3LpBoUN1d2fGruQHQLapJcP0P5iBOT6DGw7uI11Jj+FIhzbZs13J1mn
10GB0FozFzcsO9CWXDYsmjDFYAJL5ndky2ePq0D+ODaz5tvUeH5mLTN2rySzTYfqYWNBaeptPgQc
kA+NdXOH4NRfX6nO53o3E1pIu8uoUaqHmVyXvPqZeg+1NJTi5gqQ2te+vZEqOiij24HZuS0cKW4e
YUn7J+lmQeyfSBdksGdB3fUbQ/jVBY01HzoMWaWcriabSGhjnky74s6AY5s1zZvg/Te0glVUcLEn
1g6F0BpL4k12NrnNSEE2UqqcS16377cwB48xXHAfTKctTojiqfEJ6Y0q6qmnWD8d8slL5WQ6c+lB
/39hB/QzyYUFcYCaRMdYdQ0Om6pFVN0W31drUq+bywilBcS0VWIg7v333xceP7vzKPjC8LRQVdz7
s9uL1OcO+sC0GSExkmERdRBCL+CF4NSm742bXgd0q1g9yueXBDVib6LFeksPDOEv9+gFqkgRdK43
2xl6Be1IeVilsEILe2O33jBU7Q5ASSiws/2T+kqNDb5kMyUcZMURV4mFNxvGLKfjQedG9kuZVmuu
qcFr4NOGDUSgjXnqkJVHQnsu2+xj/6GgvvOaEFT5JxaOmZBE0w9dahPn/fZXv7dA8S9YUIRdqrIN
8ffDT828x66zq+CEZ637ChasDOJJBSso5c2E8OSfuaPu38M3J6RQEhntGoGny9KOBwYcxN2W/9C1
poBjLysadbmy1aNxsAzB3572AHgGrHLqyA4xrUUdn8OIutvTwfy3OfaozT6bpHRpmHegYUodfTC2
5L+gmjn0Ta8QWFZoYBI249mQl+7AOvbZI6ckNHPVY4DqbF+cPNahOIdkWwEpU++6btT+OvPo2ND8
mB5RNa5OpG6q7WB/dWNtljmbXZxYzZqWWZU3/Q6QXRaGj7NEQPxGQ2eDWt5ibtEoXuzFOotap91j
7mpeKM/IW9WrMOjTRb8jA4F8ECMELp3LxSq3veD8u67brlJLvUvjK0LLvExgGyPR+b8Rz8oyiaBB
L/trtXx/q8QUGvCO92DSd/DCm4y4+nJyy2DojNnr8Thn1cx4ctdbqhkHrVzBynA5KLo/zKmrp4+B
b8B/PFHn1N8cLoqu1Z1ENWcobsF/pwyzidg+d7fqr5gr1goI5MKB0gDbozCSVfuP4ICUexnIoogA
5BVdY/D7bQqn2oD5WTdGLT7j2Rz5tj86Sp9X7lTALsZIgp+ne+YLJ9Jnx/y60aem
`protect end_protected
