localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTY_CHK = {
  {32'h4022ddbb, 32'hc15a51ce} /* (15, 15, 15) {real, imag} */,
  {32'hbfed6999, 32'hc098c435} /* (15, 15, 14) {real, imag} */,
  {32'h4072d7e0, 32'h3e0cab98} /* (15, 15, 13) {real, imag} */,
  {32'h4078a7bc, 32'h408c66ed} /* (15, 15, 12) {real, imag} */,
  {32'hc0a9172d, 32'h40b4d249} /* (15, 15, 11) {real, imag} */,
  {32'hc1117fc8, 32'h40b596d4} /* (15, 15, 10) {real, imag} */,
  {32'hc06b997b, 32'h40ef9a80} /* (15, 15, 9) {real, imag} */,
  {32'h41061487, 32'h40f77d56} /* (15, 15, 8) {real, imag} */,
  {32'h405664e7, 32'h40b318a6} /* (15, 15, 7) {real, imag} */,
  {32'hbdb3e790, 32'hc0f0005c} /* (15, 15, 6) {real, imag} */,
  {32'hc0036953, 32'hc12184c4} /* (15, 15, 5) {real, imag} */,
  {32'hc053c8ab, 32'hc1112ef0} /* (15, 15, 4) {real, imag} */,
  {32'h412721d9, 32'h3ff13a06} /* (15, 15, 3) {real, imag} */,
  {32'h41252939, 32'h4134ce67} /* (15, 15, 2) {real, imag} */,
  {32'hbfe300aa, 32'h40b2345d} /* (15, 15, 1) {real, imag} */,
  {32'hc04ffc67, 32'hc0140e00} /* (15, 15, 0) {real, imag} */,
  {32'hbfc665b9, 32'h40a2bbc8} /* (15, 14, 15) {real, imag} */,
  {32'hc054ea5b, 32'h4144090e} /* (15, 14, 14) {real, imag} */,
  {32'hc09fd2e0, 32'h4112f1bc} /* (15, 14, 13) {real, imag} */,
  {32'hc03e690f, 32'h40db615d} /* (15, 14, 12) {real, imag} */,
  {32'hc016f80c, 32'hc07d4d9a} /* (15, 14, 11) {real, imag} */,
  {32'h3f4d550e, 32'h3f1cf0d6} /* (15, 14, 10) {real, imag} */,
  {32'h4008a175, 32'h40ee0f39} /* (15, 14, 9) {real, imag} */,
  {32'h40b968f9, 32'hbfe0ef3e} /* (15, 14, 8) {real, imag} */,
  {32'h3ea712fc, 32'h3f124818} /* (15, 14, 7) {real, imag} */,
  {32'h3f482a70, 32'h40fd331d} /* (15, 14, 6) {real, imag} */,
  {32'hc0a1c2e2, 32'h40dff288} /* (15, 14, 5) {real, imag} */,
  {32'hc0086946, 32'hbfc1d89c} /* (15, 14, 4) {real, imag} */,
  {32'hc028a500, 32'hbfc70f04} /* (15, 14, 3) {real, imag} */,
  {32'hc05eed10, 32'hc0b15d74} /* (15, 14, 2) {real, imag} */,
  {32'h3f99f580, 32'hc09f8541} /* (15, 14, 1) {real, imag} */,
  {32'h4082ce30, 32'h3ff4c59f} /* (15, 14, 0) {real, imag} */,
  {32'hc0a18550, 32'hc0088712} /* (15, 13, 15) {real, imag} */,
  {32'hc04a1150, 32'h3fe4405a} /* (15, 13, 14) {real, imag} */,
  {32'hbfd6114e, 32'h40fd07bc} /* (15, 13, 13) {real, imag} */,
  {32'h4036d7d4, 32'h3e30d400} /* (15, 13, 12) {real, imag} */,
  {32'h411dafab, 32'hc07e9736} /* (15, 13, 11) {real, imag} */,
  {32'h4105e3c8, 32'hc0c138be} /* (15, 13, 10) {real, imag} */,
  {32'h40e34e38, 32'hc0236ee2} /* (15, 13, 9) {real, imag} */,
  {32'h40d8b3e1, 32'hc05165ca} /* (15, 13, 8) {real, imag} */,
  {32'hbf9b85cc, 32'hc119150a} /* (15, 13, 7) {real, imag} */,
  {32'hbff8c8ee, 32'hc00ea7e1} /* (15, 13, 6) {real, imag} */,
  {32'hc00b10fd, 32'h40949f88} /* (15, 13, 5) {real, imag} */,
  {32'hc12837a2, 32'hbfd8d9ea} /* (15, 13, 4) {real, imag} */,
  {32'hc16001bd, 32'hc07ec468} /* (15, 13, 3) {real, imag} */,
  {32'hc0bf0fee, 32'hc0061128} /* (15, 13, 2) {real, imag} */,
  {32'h40a21c7f, 32'h409df68a} /* (15, 13, 1) {real, imag} */,
  {32'hc0415242, 32'hbe9df210} /* (15, 13, 0) {real, imag} */,
  {32'h3fee11af, 32'h40378732} /* (15, 12, 15) {real, imag} */,
  {32'h40ba0014, 32'h40728696} /* (15, 12, 14) {real, imag} */,
  {32'h3feab27c, 32'h405cbb86} /* (15, 12, 13) {real, imag} */,
  {32'hc0c6f970, 32'h3fe6d0d2} /* (15, 12, 12) {real, imag} */,
  {32'hc0b7e1b6, 32'h3f485190} /* (15, 12, 11) {real, imag} */,
  {32'hbfcd25b4, 32'h405c19ff} /* (15, 12, 10) {real, imag} */,
  {32'hbfb6f250, 32'hc03b9d61} /* (15, 12, 9) {real, imag} */,
  {32'hc0c9b726, 32'hc0d36d04} /* (15, 12, 8) {real, imag} */,
  {32'hc1028096, 32'h4095903a} /* (15, 12, 7) {real, imag} */,
  {32'hc0488df4, 32'h40ebe22b} /* (15, 12, 6) {real, imag} */,
  {32'h40880707, 32'h40cfca54} /* (15, 12, 5) {real, imag} */,
  {32'h3f0fe1a8, 32'hc0a34855} /* (15, 12, 4) {real, imag} */,
  {32'h3e93cec0, 32'h402b8902} /* (15, 12, 3) {real, imag} */,
  {32'h41085e34, 32'h40ae6f62} /* (15, 12, 2) {real, imag} */,
  {32'h40ae89ff, 32'h3f3abf84} /* (15, 12, 1) {real, imag} */,
  {32'hbf8b3d4b, 32'h3e6f6ca0} /* (15, 12, 0) {real, imag} */,
  {32'h3f0f2c22, 32'hbf9b9697} /* (15, 11, 15) {real, imag} */,
  {32'h3fb734cd, 32'hc0c66555} /* (15, 11, 14) {real, imag} */,
  {32'h3f9ae81e, 32'hc0b18da4} /* (15, 11, 13) {real, imag} */,
  {32'hc00315a0, 32'hc0d17ac7} /* (15, 11, 12) {real, imag} */,
  {32'hc02c6458, 32'h402bd80a} /* (15, 11, 11) {real, imag} */,
  {32'hc0a16374, 32'h3f900df4} /* (15, 11, 10) {real, imag} */,
  {32'hc02f92cc, 32'hbf7b7890} /* (15, 11, 9) {real, imag} */,
  {32'h3f3c6388, 32'h3f3a74c8} /* (15, 11, 8) {real, imag} */,
  {32'h40adf6dc, 32'hc0c8e8f2} /* (15, 11, 7) {real, imag} */,
  {32'h408b5d72, 32'hc111ed84} /* (15, 11, 6) {real, imag} */,
  {32'hbf21392c, 32'hc0d534e3} /* (15, 11, 5) {real, imag} */,
  {32'hbfb4843a, 32'hc0cbbbe7} /* (15, 11, 4) {real, imag} */,
  {32'hbf9ae63c, 32'hc0e55006} /* (15, 11, 3) {real, imag} */,
  {32'hc07c9163, 32'h3f402c5a} /* (15, 11, 2) {real, imag} */,
  {32'hc0205409, 32'h403524e7} /* (15, 11, 1) {real, imag} */,
  {32'hbfc0bca6, 32'hc030f520} /* (15, 11, 0) {real, imag} */,
  {32'hbf8a2858, 32'h3f519eb0} /* (15, 10, 15) {real, imag} */,
  {32'hbf010630, 32'hc08154f2} /* (15, 10, 14) {real, imag} */,
  {32'h4043476b, 32'hc0a9fedb} /* (15, 10, 13) {real, imag} */,
  {32'h40a8ec3b, 32'h406e8a3f} /* (15, 10, 12) {real, imag} */,
  {32'h4052e8a6, 32'h3f22716c} /* (15, 10, 11) {real, imag} */,
  {32'hbe7a3df4, 32'hbfbfc4cc} /* (15, 10, 10) {real, imag} */,
  {32'h405d8756, 32'hc065f75c} /* (15, 10, 9) {real, imag} */,
  {32'h40536c28, 32'hc00b021a} /* (15, 10, 8) {real, imag} */,
  {32'h3f4ac536, 32'h401c6fd8} /* (15, 10, 7) {real, imag} */,
  {32'hbef265d8, 32'h4069776d} /* (15, 10, 6) {real, imag} */,
  {32'hc02cbb53, 32'hbf8a00fe} /* (15, 10, 5) {real, imag} */,
  {32'h4088b2b3, 32'h3f40b354} /* (15, 10, 4) {real, imag} */,
  {32'h409cb9ae, 32'h4022d9f0} /* (15, 10, 3) {real, imag} */,
  {32'hbec7b7d0, 32'h3f9188f5} /* (15, 10, 2) {real, imag} */,
  {32'hc0699be6, 32'hbf4adb8e} /* (15, 10, 1) {real, imag} */,
  {32'hba11c000, 32'h3f99f883} /* (15, 10, 0) {real, imag} */,
  {32'h3e9fc232, 32'hbff1b38c} /* (15, 9, 15) {real, imag} */,
  {32'hbea5f56c, 32'h3f285bb6} /* (15, 9, 14) {real, imag} */,
  {32'hbe007788, 32'h40063dd5} /* (15, 9, 13) {real, imag} */,
  {32'h3f90025e, 32'hc00b0f46} /* (15, 9, 12) {real, imag} */,
  {32'hbf2d3a73, 32'hbffc3a3f} /* (15, 9, 11) {real, imag} */,
  {32'hbf41a620, 32'hc01306c9} /* (15, 9, 10) {real, imag} */,
  {32'hbd5c4a80, 32'h3fe09638} /* (15, 9, 9) {real, imag} */,
  {32'h3ed4a2fc, 32'hbebbc380} /* (15, 9, 8) {real, imag} */,
  {32'h3d9faa98, 32'hc0230b72} /* (15, 9, 7) {real, imag} */,
  {32'h3f9f2baa, 32'hbe814f6a} /* (15, 9, 6) {real, imag} */,
  {32'h401d0ceb, 32'hbf347f5a} /* (15, 9, 5) {real, imag} */,
  {32'h40665e9a, 32'h3e8a15c8} /* (15, 9, 4) {real, imag} */,
  {32'h3fa15db0, 32'hbf4f9f92} /* (15, 9, 3) {real, imag} */,
  {32'hbf1fed2c, 32'h3f59289c} /* (15, 9, 2) {real, imag} */,
  {32'h4003f557, 32'h404cca58} /* (15, 9, 1) {real, imag} */,
  {32'h3eeea5d0, 32'h3ef3cbf0} /* (15, 9, 0) {real, imag} */,
  {32'hbe912a88, 32'h3e7383a0} /* (15, 8, 15) {real, imag} */,
  {32'h3ff1b44a, 32'h3dff4e80} /* (15, 8, 14) {real, imag} */,
  {32'hbfc52204, 32'hc00c29c3} /* (15, 8, 13) {real, imag} */,
  {32'h3e33af00, 32'hbf7495f4} /* (15, 8, 12) {real, imag} */,
  {32'h3efa4f38, 32'h3ff412ee} /* (15, 8, 11) {real, imag} */,
  {32'h400a2426, 32'hbd9d4cf0} /* (15, 8, 10) {real, imag} */,
  {32'hbefe2a68, 32'hbfc138f1} /* (15, 8, 9) {real, imag} */,
  {32'hc04dad22, 32'hbff15a9a} /* (15, 8, 8) {real, imag} */,
  {32'h3d32ec60, 32'hc04be960} /* (15, 8, 7) {real, imag} */,
  {32'hbd665d00, 32'h3f9744d1} /* (15, 8, 6) {real, imag} */,
  {32'hbf738500, 32'h4050d6fe} /* (15, 8, 5) {real, imag} */,
  {32'h3e3c9c80, 32'h4032b2b4} /* (15, 8, 4) {real, imag} */,
  {32'h3d2863e0, 32'h3dc6dd80} /* (15, 8, 3) {real, imag} */,
  {32'hbf9c2a26, 32'h3f82a31a} /* (15, 8, 2) {real, imag} */,
  {32'hc00a7ee6, 32'h3f5c7a94} /* (15, 8, 1) {real, imag} */,
  {32'hc01c9c11, 32'h3f1ed806} /* (15, 8, 0) {real, imag} */,
  {32'hbf812fb0, 32'hbf260418} /* (15, 7, 15) {real, imag} */,
  {32'h3ff32a0f, 32'h3f34994e} /* (15, 7, 14) {real, imag} */,
  {32'h406907f4, 32'h40318187} /* (15, 7, 13) {real, imag} */,
  {32'h3e33802c, 32'hbe5f8964} /* (15, 7, 12) {real, imag} */,
  {32'h3f01f8ad, 32'hbfee83e1} /* (15, 7, 11) {real, imag} */,
  {32'h3f05f7f0, 32'hbfc32ed2} /* (15, 7, 10) {real, imag} */,
  {32'hbd1e8200, 32'h3ffedf6c} /* (15, 7, 9) {real, imag} */,
  {32'h3f1519f2, 32'h40b8e6ee} /* (15, 7, 8) {real, imag} */,
  {32'hbefdf1d2, 32'h408f6a19} /* (15, 7, 7) {real, imag} */,
  {32'hbef353d2, 32'hbf8fc3a2} /* (15, 7, 6) {real, imag} */,
  {32'hbf25f2f4, 32'h3f57f936} /* (15, 7, 5) {real, imag} */,
  {32'h3f5e7b20, 32'h3f029d4c} /* (15, 7, 4) {real, imag} */,
  {32'hbf1d5f70, 32'hbfa1910b} /* (15, 7, 3) {real, imag} */,
  {32'h40141013, 32'hbfff36ce} /* (15, 7, 2) {real, imag} */,
  {32'h4089f9f4, 32'hbf89f9c3} /* (15, 7, 1) {real, imag} */,
  {32'h400b4622, 32'h3f98b69c} /* (15, 7, 0) {real, imag} */,
  {32'h401e6c25, 32'h40a60dda} /* (15, 6, 15) {real, imag} */,
  {32'h4093da05, 32'h40504429} /* (15, 6, 14) {real, imag} */,
  {32'hbee8ad48, 32'hc0a4b6cb} /* (15, 6, 13) {real, imag} */,
  {32'hbfad2f4f, 32'hbf81d1f6} /* (15, 6, 12) {real, imag} */,
  {32'h3f96619c, 32'h4022dccb} /* (15, 6, 11) {real, imag} */,
  {32'hbfa714b8, 32'hc0274d58} /* (15, 6, 10) {real, imag} */,
  {32'hbfb1a319, 32'hc0a773d6} /* (15, 6, 9) {real, imag} */,
  {32'hbfae7fcb, 32'hbfce2330} /* (15, 6, 8) {real, imag} */,
  {32'hc0479cb2, 32'hbf9e450b} /* (15, 6, 7) {real, imag} */,
  {32'hbf838596, 32'hbec1c598} /* (15, 6, 6) {real, imag} */,
  {32'hbfeda80e, 32'hbf137c8b} /* (15, 6, 5) {real, imag} */,
  {32'h40c452e5, 32'h3da59920} /* (15, 6, 4) {real, imag} */,
  {32'h406b1bd8, 32'h3f9b2bb5} /* (15, 6, 3) {real, imag} */,
  {32'h3fe6ec88, 32'hbf8be511} /* (15, 6, 2) {real, imag} */,
  {32'h40210af4, 32'h400e3e34} /* (15, 6, 1) {real, imag} */,
  {32'h3f8be298, 32'h408c614c} /* (15, 6, 0) {real, imag} */,
  {32'h408f18bb, 32'h4072591a} /* (15, 5, 15) {real, imag} */,
  {32'hbe8c4fe4, 32'h40870d43} /* (15, 5, 14) {real, imag} */,
  {32'hc09274ce, 32'h40854222} /* (15, 5, 13) {real, imag} */,
  {32'h3fc54b10, 32'h3feeb67c} /* (15, 5, 12) {real, imag} */,
  {32'hbeabb9a0, 32'hc0416ff4} /* (15, 5, 11) {real, imag} */,
  {32'h3f4bdf94, 32'h3f877154} /* (15, 5, 10) {real, imag} */,
  {32'hc05458bc, 32'hbed0a8e0} /* (15, 5, 9) {real, imag} */,
  {32'hc114e906, 32'hc0d655e1} /* (15, 5, 8) {real, imag} */,
  {32'hc09edaaa, 32'hc056452c} /* (15, 5, 7) {real, imag} */,
  {32'hbf0bd8a0, 32'hc03c9b47} /* (15, 5, 6) {real, imag} */,
  {32'h3fc0dd7e, 32'hbc12f800} /* (15, 5, 5) {real, imag} */,
  {32'hbe017030, 32'h3fc35d14} /* (15, 5, 4) {real, imag} */,
  {32'h3dea6340, 32'h3fbf6fe6} /* (15, 5, 3) {real, imag} */,
  {32'hc0a7115a, 32'h3f2f970c} /* (15, 5, 2) {real, imag} */,
  {32'hc0577399, 32'hbfbf4762} /* (15, 5, 1) {real, imag} */,
  {32'h40ac9b24, 32'hc0019e50} /* (15, 5, 0) {real, imag} */,
  {32'hc0baa896, 32'hbffe7b1d} /* (15, 4, 15) {real, imag} */,
  {32'hc11d1882, 32'h40bd4b31} /* (15, 4, 14) {real, imag} */,
  {32'hc084e747, 32'h412df8aa} /* (15, 4, 13) {real, imag} */,
  {32'h402c26e8, 32'h4012f92b} /* (15, 4, 12) {real, imag} */,
  {32'hc081fc6a, 32'h3d2c3f80} /* (15, 4, 11) {real, imag} */,
  {32'hc0bf1001, 32'h3f9b46f2} /* (15, 4, 10) {real, imag} */,
  {32'hc0d5be20, 32'h40e70662} /* (15, 4, 9) {real, imag} */,
  {32'hbf2b8e50, 32'h4067bd0d} /* (15, 4, 8) {real, imag} */,
  {32'hc0495f08, 32'h41066386} /* (15, 4, 7) {real, imag} */,
  {32'h4087040e, 32'h40b9f0db} /* (15, 4, 6) {real, imag} */,
  {32'h40e33929, 32'h40e465ca} /* (15, 4, 5) {real, imag} */,
  {32'h40575db2, 32'h40c3a763} /* (15, 4, 4) {real, imag} */,
  {32'h410ee522, 32'hbf9a3c97} /* (15, 4, 3) {real, imag} */,
  {32'h4116d3b4, 32'hc01fcf5b} /* (15, 4, 2) {real, imag} */,
  {32'h4086c73b, 32'hc0d6957e} /* (15, 4, 1) {real, imag} */,
  {32'hc08cd836, 32'hc083fb8c} /* (15, 4, 0) {real, imag} */,
  {32'hbec61428, 32'hbfaeaef1} /* (15, 3, 15) {real, imag} */,
  {32'h40454f34, 32'hc0a42db6} /* (15, 3, 14) {real, imag} */,
  {32'h40dad4ce, 32'hc08b3cfe} /* (15, 3, 13) {real, imag} */,
  {32'h40e68e6a, 32'hc02d5360} /* (15, 3, 12) {real, imag} */,
  {32'hc09d4644, 32'h3f0a4452} /* (15, 3, 11) {real, imag} */,
  {32'hc1821158, 32'h40abc744} /* (15, 3, 10) {real, imag} */,
  {32'hc170e040, 32'hc1142b72} /* (15, 3, 9) {real, imag} */,
  {32'hc0caef89, 32'hc001812e} /* (15, 3, 8) {real, imag} */,
  {32'h3fbe561a, 32'hc0221096} /* (15, 3, 7) {real, imag} */,
  {32'h40b0b626, 32'h3f0d2744} /* (15, 3, 6) {real, imag} */,
  {32'hbfc37fce, 32'hc11a1638} /* (15, 3, 5) {real, imag} */,
  {32'hc13c623e, 32'hbdecfe80} /* (15, 3, 4) {real, imag} */,
  {32'hbf838c70, 32'hbe97ff90} /* (15, 3, 3) {real, imag} */,
  {32'h4069ae23, 32'hc03e13fe} /* (15, 3, 2) {real, imag} */,
  {32'h4078e706, 32'hc08f9950} /* (15, 3, 1) {real, imag} */,
  {32'hc016fc74, 32'hc0de8a57} /* (15, 3, 0) {real, imag} */,
  {32'hbff07d3b, 32'h404c3c93} /* (15, 2, 15) {real, imag} */,
  {32'h40ccde6a, 32'hc030d138} /* (15, 2, 14) {real, imag} */,
  {32'h400b4224, 32'hc137ed30} /* (15, 2, 13) {real, imag} */,
  {32'hc01f21e9, 32'hc1542abc} /* (15, 2, 12) {real, imag} */,
  {32'h3fa9609f, 32'hc12c8186} /* (15, 2, 11) {real, imag} */,
  {32'hc0879099, 32'hbedd1040} /* (15, 2, 10) {real, imag} */,
  {32'h40db19bc, 32'h40e97613} /* (15, 2, 9) {real, imag} */,
  {32'hc139f26a, 32'h410664aa} /* (15, 2, 8) {real, imag} */,
  {32'hc0545a14, 32'h411b29b0} /* (15, 2, 7) {real, imag} */,
  {32'h4127bb8b, 32'h40d10e4b} /* (15, 2, 6) {real, imag} */,
  {32'h41946c88, 32'h40473d50} /* (15, 2, 5) {real, imag} */,
  {32'h4135a7fe, 32'h4166f47a} /* (15, 2, 4) {real, imag} */,
  {32'h3f9adfe0, 32'h4150fc08} /* (15, 2, 3) {real, imag} */,
  {32'h3eb4e110, 32'h405d9740} /* (15, 2, 2) {real, imag} */,
  {32'hc1519fee, 32'h4105896b} /* (15, 2, 1) {real, imag} */,
  {32'hc0e6bdfa, 32'h403438f6} /* (15, 2, 0) {real, imag} */,
  {32'hbf90ed9a, 32'hc0fb6273} /* (15, 1, 15) {real, imag} */,
  {32'h400032fe, 32'h3e2d60a0} /* (15, 1, 14) {real, imag} */,
  {32'h3f40c410, 32'h3ea217dc} /* (15, 1, 13) {real, imag} */,
  {32'hc06e2d08, 32'h40b42c75} /* (15, 1, 12) {real, imag} */,
  {32'h4095859b, 32'h40f1fac7} /* (15, 1, 11) {real, imag} */,
  {32'hc00eac82, 32'hc11d97cc} /* (15, 1, 10) {real, imag} */,
  {32'h40bfcb0a, 32'hc0d7a734} /* (15, 1, 9) {real, imag} */,
  {32'h404c61b0, 32'hbfd17280} /* (15, 1, 8) {real, imag} */,
  {32'hbf643104, 32'hc050775c} /* (15, 1, 7) {real, imag} */,
  {32'hc035aac4, 32'h40f5e216} /* (15, 1, 6) {real, imag} */,
  {32'hbfd53d36, 32'h4130994c} /* (15, 1, 5) {real, imag} */,
  {32'hc0e243fa, 32'hbf22b428} /* (15, 1, 4) {real, imag} */,
  {32'hc15f7deb, 32'hc0b0ee74} /* (15, 1, 3) {real, imag} */,
  {32'hbff9aed8, 32'hbfa69438} /* (15, 1, 2) {real, imag} */,
  {32'h4039c151, 32'hc0e2680b} /* (15, 1, 1) {real, imag} */,
  {32'hc0920942, 32'hc0c13ada} /* (15, 1, 0) {real, imag} */,
  {32'hbfbaaf54, 32'hc0de9a29} /* (15, 0, 15) {real, imag} */,
  {32'hc1193de5, 32'hc10fbf6b} /* (15, 0, 14) {real, imag} */,
  {32'h406fe0e2, 32'h3fe6aada} /* (15, 0, 13) {real, imag} */,
  {32'h41585c6c, 32'hc0a5e49e} /* (15, 0, 12) {real, imag} */,
  {32'h40df48fe, 32'hc0ed6e02} /* (15, 0, 11) {real, imag} */,
  {32'h41476c78, 32'h400acd20} /* (15, 0, 10) {real, imag} */,
  {32'hc103f713, 32'hc098eaa1} /* (15, 0, 9) {real, imag} */,
  {32'h404fe66a, 32'h3e0f4270} /* (15, 0, 8) {real, imag} */,
  {32'hbfb3c773, 32'hc11e1d8d} /* (15, 0, 7) {real, imag} */,
  {32'hc1929d0a, 32'h4091f8ca} /* (15, 0, 6) {real, imag} */,
  {32'hc1a86718, 32'h41853068} /* (15, 0, 5) {real, imag} */,
  {32'hc11a16ae, 32'hc0c68c86} /* (15, 0, 4) {real, imag} */,
  {32'h3f27f4aa, 32'hc12985ad} /* (15, 0, 3) {real, imag} */,
  {32'hbf93a9fe, 32'hc10ee227} /* (15, 0, 2) {real, imag} */,
  {32'h401330fa, 32'hc09681c2} /* (15, 0, 1) {real, imag} */,
  {32'h40fef530, 32'h3f2deb12} /* (15, 0, 0) {real, imag} */,
  {32'h40012f0d, 32'hc0a083a3} /* (14, 15, 15) {real, imag} */,
  {32'h40ebd6e4, 32'hc16111e8} /* (14, 15, 14) {real, imag} */,
  {32'hbfdc2700, 32'hc12db6fe} /* (14, 15, 13) {real, imag} */,
  {32'h4053dff2, 32'hbffccc40} /* (14, 15, 12) {real, imag} */,
  {32'h407b98a6, 32'h4127d691} /* (14, 15, 11) {real, imag} */,
  {32'h41041e67, 32'h408f3b26} /* (14, 15, 10) {real, imag} */,
  {32'h415cbc82, 32'hc174d5c2} /* (14, 15, 9) {real, imag} */,
  {32'h40748956, 32'hc0e5a755} /* (14, 15, 8) {real, imag} */,
  {32'h40db76a5, 32'h40aa330a} /* (14, 15, 7) {real, imag} */,
  {32'h410129a4, 32'h40dce82c} /* (14, 15, 6) {real, imag} */,
  {32'h410b98c6, 32'h40e8fcd6} /* (14, 15, 5) {real, imag} */,
  {32'hc017026e, 32'h4129cb49} /* (14, 15, 4) {real, imag} */,
  {32'hc137e89a, 32'h3fad55b8} /* (14, 15, 3) {real, imag} */,
  {32'hc095e15f, 32'hbfa8eac4} /* (14, 15, 2) {real, imag} */,
  {32'hc05bf431, 32'h4036163d} /* (14, 15, 1) {real, imag} */,
  {32'hc091ee38, 32'hbf21b1b4} /* (14, 15, 0) {real, imag} */,
  {32'h40c86fb7, 32'h4085f157} /* (14, 14, 15) {real, imag} */,
  {32'h3ff69560, 32'h4154cf00} /* (14, 14, 14) {real, imag} */,
  {32'h40ff0268, 32'hc02be188} /* (14, 14, 13) {real, imag} */,
  {32'h41a614cb, 32'hc1425ddb} /* (14, 14, 12) {real, imag} */,
  {32'h40167198, 32'hc09651ae} /* (14, 14, 11) {real, imag} */,
  {32'hc0f420b6, 32'hbedd49a0} /* (14, 14, 10) {real, imag} */,
  {32'hc112e76d, 32'h40b39a38} /* (14, 14, 9) {real, imag} */,
  {32'hc059956a, 32'hbe26e6a0} /* (14, 14, 8) {real, imag} */,
  {32'h3fa99f34, 32'h4107bc72} /* (14, 14, 7) {real, imag} */,
  {32'hbffaa2a0, 32'h409b100c} /* (14, 14, 6) {real, imag} */,
  {32'h40b16fc4, 32'hc09c3c0e} /* (14, 14, 5) {real, imag} */,
  {32'h3f2f03e6, 32'h40c655f2} /* (14, 14, 4) {real, imag} */,
  {32'h4081af97, 32'h410fc3a4} /* (14, 14, 3) {real, imag} */,
  {32'hc0be89c6, 32'hc017c15a} /* (14, 14, 2) {real, imag} */,
  {32'hc0eb90d3, 32'hc1079d9a} /* (14, 14, 1) {real, imag} */,
  {32'hc016eee0, 32'hc098d7be} /* (14, 14, 0) {real, imag} */,
  {32'h407b3e59, 32'h3f257dca} /* (14, 13, 15) {real, imag} */,
  {32'h40939506, 32'hc1230f42} /* (14, 13, 14) {real, imag} */,
  {32'hbf760f13, 32'hc000f572} /* (14, 13, 13) {real, imag} */,
  {32'hc10e8358, 32'h40f84a0d} /* (14, 13, 12) {real, imag} */,
  {32'hc0f4df02, 32'h3f72436f} /* (14, 13, 11) {real, imag} */,
  {32'h3f69f23c, 32'h3fff7294} /* (14, 13, 10) {real, imag} */,
  {32'h400e699e, 32'hbfb501de} /* (14, 13, 9) {real, imag} */,
  {32'hc0550052, 32'hc0dbf4ec} /* (14, 13, 8) {real, imag} */,
  {32'hc0b175fe, 32'hc028f5eb} /* (14, 13, 7) {real, imag} */,
  {32'hc0d06a93, 32'hbf534870} /* (14, 13, 6) {real, imag} */,
  {32'hc120e63d, 32'hbff4ddaf} /* (14, 13, 5) {real, imag} */,
  {32'hc0b40c22, 32'h40126e76} /* (14, 13, 4) {real, imag} */,
  {32'hc011dc38, 32'hbfbc2148} /* (14, 13, 3) {real, imag} */,
  {32'h3fc974a4, 32'h40092706} /* (14, 13, 2) {real, imag} */,
  {32'h3fdaa885, 32'h40a7ed8c} /* (14, 13, 1) {real, imag} */,
  {32'hc0f79c5d, 32'h40da488c} /* (14, 13, 0) {real, imag} */,
  {32'hc0c150e1, 32'hc0a0226a} /* (14, 12, 15) {real, imag} */,
  {32'hc0d2a300, 32'hc1169f12} /* (14, 12, 14) {real, imag} */,
  {32'h3e94ae24, 32'hc0ca276e} /* (14, 12, 13) {real, imag} */,
  {32'h3f713aa0, 32'h3f880a04} /* (14, 12, 12) {real, imag} */,
  {32'hc0171099, 32'h40ad1c21} /* (14, 12, 11) {real, imag} */,
  {32'hc04f69e0, 32'hc05141f2} /* (14, 12, 10) {real, imag} */,
  {32'hbf2cd3f0, 32'hc0154cf8} /* (14, 12, 9) {real, imag} */,
  {32'hc09f0fc1, 32'hbfd7052c} /* (14, 12, 8) {real, imag} */,
  {32'hbf1f3ad8, 32'hbfb61376} /* (14, 12, 7) {real, imag} */,
  {32'hc091595a, 32'h407c870c} /* (14, 12, 6) {real, imag} */,
  {32'hc0c64c3a, 32'h408dd898} /* (14, 12, 5) {real, imag} */,
  {32'hbeb826b2, 32'h407a0fda} /* (14, 12, 4) {real, imag} */,
  {32'h407f276e, 32'h40e8cf12} /* (14, 12, 3) {real, imag} */,
  {32'h40a4276a, 32'h40802794} /* (14, 12, 2) {real, imag} */,
  {32'hc0ce8a97, 32'h40aa20e2} /* (14, 12, 1) {real, imag} */,
  {32'hc0862a0a, 32'h4080211d} /* (14, 12, 0) {real, imag} */,
  {32'hbfc2eae0, 32'h3e6ce860} /* (14, 11, 15) {real, imag} */,
  {32'hc0871b10, 32'h3f62ff34} /* (14, 11, 14) {real, imag} */,
  {32'hc0c5e813, 32'h40040c22} /* (14, 11, 13) {real, imag} */,
  {32'hbfa2d20e, 32'h40783345} /* (14, 11, 12) {real, imag} */,
  {32'hc05f4d92, 32'hc0ce8286} /* (14, 11, 11) {real, imag} */,
  {32'hc0558982, 32'hc0fdf62a} /* (14, 11, 10) {real, imag} */,
  {32'h40c6fed8, 32'hc017936a} /* (14, 11, 9) {real, imag} */,
  {32'h3f8823e1, 32'hc01c18ba} /* (14, 11, 8) {real, imag} */,
  {32'h3ecf8610, 32'h3fc710fa} /* (14, 11, 7) {real, imag} */,
  {32'h4083322e, 32'hc090544b} /* (14, 11, 6) {real, imag} */,
  {32'hc01f37c8, 32'hc0f4ad26} /* (14, 11, 5) {real, imag} */,
  {32'h3eb1a868, 32'hbde30960} /* (14, 11, 4) {real, imag} */,
  {32'hc062bcfb, 32'h40442ecc} /* (14, 11, 3) {real, imag} */,
  {32'hbffb7734, 32'hbf8886d8} /* (14, 11, 2) {real, imag} */,
  {32'h404408b6, 32'hc03d72d6} /* (14, 11, 1) {real, imag} */,
  {32'hbf0f1874, 32'hbff45587} /* (14, 11, 0) {real, imag} */,
  {32'h3ee48046, 32'h3eb13bbc} /* (14, 10, 15) {real, imag} */,
  {32'h4017a474, 32'h3f943035} /* (14, 10, 14) {real, imag} */,
  {32'hbf8f5b64, 32'h3da0d1e0} /* (14, 10, 13) {real, imag} */,
  {32'h405fa6af, 32'h3f67cef7} /* (14, 10, 12) {real, imag} */,
  {32'h406bdb12, 32'hc053f92e} /* (14, 10, 11) {real, imag} */,
  {32'h400f2cbe, 32'hbf30e1ca} /* (14, 10, 10) {real, imag} */,
  {32'hbf1217f4, 32'h4043003c} /* (14, 10, 9) {real, imag} */,
  {32'h40029168, 32'hbfc010b3} /* (14, 10, 8) {real, imag} */,
  {32'hbfc37bc2, 32'hc0483106} /* (14, 10, 7) {real, imag} */,
  {32'hc08f3c0a, 32'h3e1f91b8} /* (14, 10, 6) {real, imag} */,
  {32'h3ea36108, 32'hbea23baa} /* (14, 10, 5) {real, imag} */,
  {32'hc09c4de6, 32'h3fe1e8d7} /* (14, 10, 4) {real, imag} */,
  {32'hc0c72654, 32'hc01a9cb3} /* (14, 10, 3) {real, imag} */,
  {32'hbf6d3c96, 32'hc04d9fac} /* (14, 10, 2) {real, imag} */,
  {32'hbe4d59fc, 32'h3fa366d5} /* (14, 10, 1) {real, imag} */,
  {32'hbf7bf162, 32'hbff59053} /* (14, 10, 0) {real, imag} */,
  {32'hbf179efc, 32'hbd1c3580} /* (14, 9, 15) {real, imag} */,
  {32'h3f38e769, 32'h3f6f674c} /* (14, 9, 14) {real, imag} */,
  {32'h4078f63e, 32'h3f5524ff} /* (14, 9, 13) {real, imag} */,
  {32'h3eb75fdc, 32'h3eea0e9c} /* (14, 9, 12) {real, imag} */,
  {32'h3fdfd17a, 32'h3f32019b} /* (14, 9, 11) {real, imag} */,
  {32'h402bda6d, 32'h3f80a2c0} /* (14, 9, 10) {real, imag} */,
  {32'hbfd31d4c, 32'h3f34f018} /* (14, 9, 9) {real, imag} */,
  {32'hbfe14746, 32'h3f7feb5c} /* (14, 9, 8) {real, imag} */,
  {32'hbf295f62, 32'h3f7e540a} /* (14, 9, 7) {real, imag} */,
  {32'h3f5ac99c, 32'hc04599da} /* (14, 9, 6) {real, imag} */,
  {32'h4025244a, 32'hc025fc80} /* (14, 9, 5) {real, imag} */,
  {32'h3efc1524, 32'hc00926e9} /* (14, 9, 4) {real, imag} */,
  {32'h3fe41b06, 32'h3fb3e725} /* (14, 9, 3) {real, imag} */,
  {32'hbf2d58a0, 32'h403f9822} /* (14, 9, 2) {real, imag} */,
  {32'hc02ce289, 32'hbf0edda4} /* (14, 9, 1) {real, imag} */,
  {32'h3f8d76cd, 32'h3e102518} /* (14, 9, 0) {real, imag} */,
  {32'hbfbb733f, 32'h3fe206cf} /* (14, 8, 15) {real, imag} */,
  {32'h3f1fc818, 32'h40074eb0} /* (14, 8, 14) {real, imag} */,
  {32'h3faa8556, 32'h3f282808} /* (14, 8, 13) {real, imag} */,
  {32'h3ec0b7c0, 32'h3fa8024c} /* (14, 8, 12) {real, imag} */,
  {32'h3f4d305a, 32'h3ed76880} /* (14, 8, 11) {real, imag} */,
  {32'h3f74bc2c, 32'h3ed36784} /* (14, 8, 10) {real, imag} */,
  {32'h3daa9ed0, 32'hbff31df2} /* (14, 8, 9) {real, imag} */,
  {32'hbf2ca090, 32'hc0485a06} /* (14, 8, 8) {real, imag} */,
  {32'hbf2d6a48, 32'hc01e0390} /* (14, 8, 7) {real, imag} */,
  {32'hbfe37036, 32'h3fd55f00} /* (14, 8, 6) {real, imag} */,
  {32'hc00d41f4, 32'h3eebeae0} /* (14, 8, 5) {real, imag} */,
  {32'hbf8edd7e, 32'hc07c35b4} /* (14, 8, 4) {real, imag} */,
  {32'h40564d5b, 32'hc05d981e} /* (14, 8, 3) {real, imag} */,
  {32'h406b5331, 32'hbfcf16c6} /* (14, 8, 2) {real, imag} */,
  {32'hbf17ab58, 32'hc0570cd8} /* (14, 8, 1) {real, imag} */,
  {32'hc0085853, 32'hc02cf0b7} /* (14, 8, 0) {real, imag} */,
  {32'h40503180, 32'hbf927568} /* (14, 7, 15) {real, imag} */,
  {32'h3f7947a1, 32'h3f096fb4} /* (14, 7, 14) {real, imag} */,
  {32'hc01fc530, 32'h3fb51530} /* (14, 7, 13) {real, imag} */,
  {32'h3f68ab5e, 32'hbf2c8bd6} /* (14, 7, 12) {real, imag} */,
  {32'h3f626838, 32'hbf81d11e} /* (14, 7, 11) {real, imag} */,
  {32'h3fd3ac0e, 32'h4003c448} /* (14, 7, 10) {real, imag} */,
  {32'h3f0df650, 32'h3fa27b84} /* (14, 7, 9) {real, imag} */,
  {32'hbda16cc8, 32'hbea99c60} /* (14, 7, 8) {real, imag} */,
  {32'h3f6626ea, 32'hbfa90439} /* (14, 7, 7) {real, imag} */,
  {32'h4026136f, 32'hbf20a98a} /* (14, 7, 6) {real, imag} */,
  {32'h401e8b96, 32'h3fc5d5a5} /* (14, 7, 5) {real, imag} */,
  {32'h3fc0939f, 32'h4026a0c5} /* (14, 7, 4) {real, imag} */,
  {32'hbfeb2bf2, 32'hbe10f538} /* (14, 7, 3) {real, imag} */,
  {32'hbf817f0c, 32'hbfb2eff4} /* (14, 7, 2) {real, imag} */,
  {32'hc01a1ab5, 32'h3f7bb244} /* (14, 7, 1) {real, imag} */,
  {32'hbf8cf6c5, 32'h3ff717b3} /* (14, 7, 0) {real, imag} */,
  {32'hbf0f93c5, 32'h3fb188d9} /* (14, 6, 15) {real, imag} */,
  {32'h3f01d7f8, 32'h3ff5f5eb} /* (14, 6, 14) {real, imag} */,
  {32'h4049400e, 32'h3fb6df2e} /* (14, 6, 13) {real, imag} */,
  {32'h3fc17236, 32'hbef087b2} /* (14, 6, 12) {real, imag} */,
  {32'hbf55aed0, 32'hbffa1840} /* (14, 6, 11) {real, imag} */,
  {32'h3f815899, 32'h3fb6edd9} /* (14, 6, 10) {real, imag} */,
  {32'h3f8a5afe, 32'h4041bd02} /* (14, 6, 9) {real, imag} */,
  {32'hc020a6a0, 32'h3ed57c74} /* (14, 6, 8) {real, imag} */,
  {32'hc0429831, 32'hbfb70730} /* (14, 6, 7) {real, imag} */,
  {32'h3fff1e40, 32'hbf909a45} /* (14, 6, 6) {real, imag} */,
  {32'h409cf436, 32'h3f6c09bd} /* (14, 6, 5) {real, imag} */,
  {32'h4013ffbc, 32'hbf843569} /* (14, 6, 4) {real, imag} */,
  {32'h3fcc0130, 32'hc0680fab} /* (14, 6, 3) {real, imag} */,
  {32'h3f77e352, 32'hbfe6dec0} /* (14, 6, 2) {real, imag} */,
  {32'h3fb49a70, 32'hc081908a} /* (14, 6, 1) {real, imag} */,
  {32'hbf41402a, 32'hbf8aefe9} /* (14, 6, 0) {real, imag} */,
  {32'h3e61005c, 32'h40073579} /* (14, 5, 15) {real, imag} */,
  {32'h40b00d8e, 32'hc04ec903} /* (14, 5, 14) {real, imag} */,
  {32'h40d82e51, 32'hc0d0768b} /* (14, 5, 13) {real, imag} */,
  {32'h402ca191, 32'hc00e0793} /* (14, 5, 12) {real, imag} */,
  {32'h40a40a93, 32'hc0221c74} /* (14, 5, 11) {real, imag} */,
  {32'hc0959e7f, 32'hc0916bea} /* (14, 5, 10) {real, imag} */,
  {32'hc06a1fb7, 32'hc095e5bc} /* (14, 5, 9) {real, imag} */,
  {32'hbe633e28, 32'hc0273858} /* (14, 5, 8) {real, imag} */,
  {32'hbed07670, 32'hc04c1f7d} /* (14, 5, 7) {real, imag} */,
  {32'h3f2996b0, 32'hc0ae805f} /* (14, 5, 6) {real, imag} */,
  {32'hbcc29300, 32'hc09865ba} /* (14, 5, 5) {real, imag} */,
  {32'hbf7c9f4c, 32'h3fee0eb2} /* (14, 5, 4) {real, imag} */,
  {32'hbfe1fa7a, 32'h4008509a} /* (14, 5, 3) {real, imag} */,
  {32'h3f438178, 32'h406ab50a} /* (14, 5, 2) {real, imag} */,
  {32'hbed6bc9c, 32'h403945ca} /* (14, 5, 1) {real, imag} */,
  {32'h401d261f, 32'h3fac3619} /* (14, 5, 0) {real, imag} */,
  {32'hc0949e63, 32'h3fe379c9} /* (14, 4, 15) {real, imag} */,
  {32'hc100af50, 32'h40d9ea35} /* (14, 4, 14) {real, imag} */,
  {32'hbfdf78f7, 32'h40bb19a2} /* (14, 4, 13) {real, imag} */,
  {32'h408b517e, 32'hc0f15c8b} /* (14, 4, 12) {real, imag} */,
  {32'h401c88a7, 32'hc0878291} /* (14, 4, 11) {real, imag} */,
  {32'hc0c476be, 32'h400e9804} /* (14, 4, 10) {real, imag} */,
  {32'hc11a034f, 32'hc0625c76} /* (14, 4, 9) {real, imag} */,
  {32'hc09024f5, 32'hc07b823e} /* (14, 4, 8) {real, imag} */,
  {32'h41326866, 32'h40865480} /* (14, 4, 7) {real, imag} */,
  {32'h40c2378a, 32'hc0932802} /* (14, 4, 6) {real, imag} */,
  {32'hbfdd92c0, 32'hc1275d9a} /* (14, 4, 5) {real, imag} */,
  {32'hbefb5432, 32'hc02fe0f2} /* (14, 4, 4) {real, imag} */,
  {32'h40ee8c85, 32'h4038b114} /* (14, 4, 3) {real, imag} */,
  {32'h3f901178, 32'h3ff15644} /* (14, 4, 2) {real, imag} */,
  {32'h40a9673f, 32'hbf499ea0} /* (14, 4, 1) {real, imag} */,
  {32'h40b56bec, 32'h3ed54c20} /* (14, 4, 0) {real, imag} */,
  {32'h4003d5e3, 32'hc07ded5a} /* (14, 3, 15) {real, imag} */,
  {32'hc0357920, 32'hc07eb460} /* (14, 3, 14) {real, imag} */,
  {32'hbf51ec4b, 32'h40fe02a7} /* (14, 3, 13) {real, imag} */,
  {32'h4090278f, 32'h4047a296} /* (14, 3, 12) {real, imag} */,
  {32'h40f61dca, 32'h40133d76} /* (14, 3, 11) {real, imag} */,
  {32'hc00964e5, 32'h40af92c8} /* (14, 3, 10) {real, imag} */,
  {32'hc056e7e2, 32'h406a1a29} /* (14, 3, 9) {real, imag} */,
  {32'h3eed36ac, 32'hbfa63568} /* (14, 3, 8) {real, imag} */,
  {32'h3f8d1688, 32'hbfd8172a} /* (14, 3, 7) {real, imag} */,
  {32'hbf533828, 32'h410a22e2} /* (14, 3, 6) {real, imag} */,
  {32'hc08568da, 32'h3ffe3b3b} /* (14, 3, 5) {real, imag} */,
  {32'hbfac649e, 32'hc0e5ad0b} /* (14, 3, 4) {real, imag} */,
  {32'hc0912418, 32'hc0982a7b} /* (14, 3, 3) {real, imag} */,
  {32'hc1118e04, 32'h403fb474} /* (14, 3, 2) {real, imag} */,
  {32'h3fb5d257, 32'hbfa6df1f} /* (14, 3, 1) {real, imag} */,
  {32'h40a7aaa1, 32'hc0b0fbb0} /* (14, 3, 0) {real, imag} */,
  {32'hc0c68d29, 32'h40c6ddfd} /* (14, 2, 15) {real, imag} */,
  {32'hc17eb554, 32'h41425ce8} /* (14, 2, 14) {real, imag} */,
  {32'hc1933e7e, 32'h41473472} /* (14, 2, 13) {real, imag} */,
  {32'hc0d76bec, 32'h41592b99} /* (14, 2, 12) {real, imag} */,
  {32'h40811a01, 32'h413301ad} /* (14, 2, 11) {real, imag} */,
  {32'h40a5e47e, 32'h4025e8c3} /* (14, 2, 10) {real, imag} */,
  {32'hbfd8a368, 32'hc0c808a8} /* (14, 2, 9) {real, imag} */,
  {32'h3fd0e345, 32'hc0a708b3} /* (14, 2, 8) {real, imag} */,
  {32'h410c53e4, 32'hbfad9ca2} /* (14, 2, 7) {real, imag} */,
  {32'h40fe5e1e, 32'hc0598318} /* (14, 2, 6) {real, imag} */,
  {32'h3e58d1b0, 32'hc1066d77} /* (14, 2, 5) {real, imag} */,
  {32'hc0506546, 32'hc140b301} /* (14, 2, 4) {real, imag} */,
  {32'h3fd80113, 32'hc15458da} /* (14, 2, 3) {real, imag} */,
  {32'h3fa6ef1a, 32'hc0929c43} /* (14, 2, 2) {real, imag} */,
  {32'h405bec6e, 32'h4078d2b7} /* (14, 2, 1) {real, imag} */,
  {32'h3fe87f29, 32'h40214fb7} /* (14, 2, 0) {real, imag} */,
  {32'h3f843748, 32'hc046e772} /* (14, 1, 15) {real, imag} */,
  {32'hc0e5b0f8, 32'hc0f4556f} /* (14, 1, 14) {real, imag} */,
  {32'hc1724658, 32'hc123f6e6} /* (14, 1, 13) {real, imag} */,
  {32'hc1307b8c, 32'hc0d32c28} /* (14, 1, 12) {real, imag} */,
  {32'hbf91930b, 32'h40df3dfa} /* (14, 1, 11) {real, imag} */,
  {32'hc01f5d9c, 32'h41658447} /* (14, 1, 10) {real, imag} */,
  {32'hc0567d28, 32'h400a90f8} /* (14, 1, 9) {real, imag} */,
  {32'hbf3d5a6e, 32'h3f9ce4e4} /* (14, 1, 8) {real, imag} */,
  {32'h3fcb7adc, 32'h3fd5a735} /* (14, 1, 7) {real, imag} */,
  {32'hbfcad94a, 32'h40ce5bfe} /* (14, 1, 6) {real, imag} */,
  {32'hc115883a, 32'h3f09143c} /* (14, 1, 5) {real, imag} */,
  {32'hc0e5a97f, 32'hc0c03896} /* (14, 1, 4) {real, imag} */,
  {32'hc00685f2, 32'h400fd24d} /* (14, 1, 3) {real, imag} */,
  {32'hc08dcf69, 32'h40cd03ed} /* (14, 1, 2) {real, imag} */,
  {32'hc0a713bc, 32'h408b4efc} /* (14, 1, 1) {real, imag} */,
  {32'hc06430d4, 32'hc0a12668} /* (14, 1, 0) {real, imag} */,
  {32'h3eb685bc, 32'h3fb2c287} /* (14, 0, 15) {real, imag} */,
  {32'h4107f024, 32'h402f72b8} /* (14, 0, 14) {real, imag} */,
  {32'h407bcc25, 32'h41132d04} /* (14, 0, 13) {real, imag} */,
  {32'h40c43a5c, 32'h41450e62} /* (14, 0, 12) {real, imag} */,
  {32'h406c2714, 32'h41398d4a} /* (14, 0, 11) {real, imag} */,
  {32'h402a14f1, 32'h3fdd0063} /* (14, 0, 10) {real, imag} */,
  {32'h4040303c, 32'hc00c3619} /* (14, 0, 9) {real, imag} */,
  {32'hbf52b970, 32'h4059e926} /* (14, 0, 8) {real, imag} */,
  {32'hc0e3d55d, 32'h4189d7fa} /* (14, 0, 7) {real, imag} */,
  {32'h40960446, 32'h408f0c89} /* (14, 0, 6) {real, imag} */,
  {32'h401a5a8a, 32'h401ed3c6} /* (14, 0, 5) {real, imag} */,
  {32'h4062034d, 32'h41115963} /* (14, 0, 4) {real, imag} */,
  {32'hc003d271, 32'h3ebe0998} /* (14, 0, 3) {real, imag} */,
  {32'h40b453d8, 32'hbe3c5230} /* (14, 0, 2) {real, imag} */,
  {32'h40dcfb57, 32'h414c6ad0} /* (14, 0, 1) {real, imag} */,
  {32'h3ffdef8a, 32'h41263e29} /* (14, 0, 0) {real, imag} */,
  {32'h3f851744, 32'h40708b8c} /* (13, 15, 15) {real, imag} */,
  {32'h4007af3a, 32'h3c655000} /* (13, 15, 14) {real, imag} */,
  {32'hc00430b8, 32'hc007d16e} /* (13, 15, 13) {real, imag} */,
  {32'hbe936ebd, 32'hc16c3a87} /* (13, 15, 12) {real, imag} */,
  {32'h40b7b798, 32'hc12abfdc} /* (13, 15, 11) {real, imag} */,
  {32'h4066b7a7, 32'hc0f704e4} /* (13, 15, 10) {real, imag} */,
  {32'h401ad572, 32'h3eac7700} /* (13, 15, 9) {real, imag} */,
  {32'hbf90b43a, 32'h3f920188} /* (13, 15, 8) {real, imag} */,
  {32'hc11aaf28, 32'hbf80705e} /* (13, 15, 7) {real, imag} */,
  {32'hbfd9ab86, 32'h3fb65448} /* (13, 15, 6) {real, imag} */,
  {32'hbfaf29b2, 32'h40e6fe2a} /* (13, 15, 5) {real, imag} */,
  {32'hbc191400, 32'h40288d2a} /* (13, 15, 4) {real, imag} */,
  {32'hbfa31090, 32'hc071555f} /* (13, 15, 3) {real, imag} */,
  {32'hc138642a, 32'hc081054b} /* (13, 15, 2) {real, imag} */,
  {32'hc0be56a6, 32'hc111ab18} /* (13, 15, 1) {real, imag} */,
  {32'hc08918b8, 32'hc001e309} /* (13, 15, 0) {real, imag} */,
  {32'hc04822b8, 32'hc01475df} /* (13, 14, 15) {real, imag} */,
  {32'hc1180530, 32'hc0eff4e2} /* (13, 14, 14) {real, imag} */,
  {32'hc14e5079, 32'hc116dfe2} /* (13, 14, 13) {real, imag} */,
  {32'hc14059c2, 32'h3f67bffb} /* (13, 14, 12) {real, imag} */,
  {32'hc0bf5e92, 32'h40a36e58} /* (13, 14, 11) {real, imag} */,
  {32'h3d7dff80, 32'h3e8aa6ac} /* (13, 14, 10) {real, imag} */,
  {32'h401ef9c4, 32'h401b6a30} /* (13, 14, 9) {real, imag} */,
  {32'h408937d2, 32'h3fce95a2} /* (13, 14, 8) {real, imag} */,
  {32'hbef84f58, 32'h404d0604} /* (13, 14, 7) {real, imag} */,
  {32'hc11cc0e5, 32'h410ce28e} /* (13, 14, 6) {real, imag} */,
  {32'hc0f2994e, 32'h4103442c} /* (13, 14, 5) {real, imag} */,
  {32'h406ca0a0, 32'h3f5ee624} /* (13, 14, 4) {real, imag} */,
  {32'h3fd1a3a8, 32'hbf5e5d11} /* (13, 14, 3) {real, imag} */,
  {32'hbc411600, 32'h3fe35a6c} /* (13, 14, 2) {real, imag} */,
  {32'h40d408ef, 32'h3fa22e48} /* (13, 14, 1) {real, imag} */,
  {32'h40f67578, 32'hc03e03cb} /* (13, 14, 0) {real, imag} */,
  {32'h40909bc0, 32'hc0ca2f34} /* (13, 13, 15) {real, imag} */,
  {32'h4092036c, 32'hc0a68358} /* (13, 13, 14) {real, imag} */,
  {32'hbfd54192, 32'h3df57e20} /* (13, 13, 13) {real, imag} */,
  {32'h40861ea3, 32'hbfdef296} /* (13, 13, 12) {real, imag} */,
  {32'hc0623bf1, 32'hbe182e90} /* (13, 13, 11) {real, imag} */,
  {32'hc090a77c, 32'hc037598f} /* (13, 13, 10) {real, imag} */,
  {32'h3f3c93e8, 32'hc1023446} /* (13, 13, 9) {real, imag} */,
  {32'h40bf22b4, 32'h3f35582a} /* (13, 13, 8) {real, imag} */,
  {32'h40651ff0, 32'h4032dd9a} /* (13, 13, 7) {real, imag} */,
  {32'h4117ce8e, 32'hc0ab5920} /* (13, 13, 6) {real, imag} */,
  {32'h40c3c09c, 32'hbf0e403a} /* (13, 13, 5) {real, imag} */,
  {32'hbd765ff0, 32'h3fc28c06} /* (13, 13, 4) {real, imag} */,
  {32'hc00ca082, 32'h3ffbb364} /* (13, 13, 3) {real, imag} */,
  {32'hbfecabc0, 32'hbf9b8f16} /* (13, 13, 2) {real, imag} */,
  {32'hbe2b2fe0, 32'h406f3756} /* (13, 13, 1) {real, imag} */,
  {32'hbf85f555, 32'h40e3926a} /* (13, 13, 0) {real, imag} */,
  {32'h404e34fb, 32'hc03817b8} /* (13, 12, 15) {real, imag} */,
  {32'h4027b99b, 32'hbde7a8f0} /* (13, 12, 14) {real, imag} */,
  {32'hc034d7ca, 32'h40b27098} /* (13, 12, 13) {real, imag} */,
  {32'hc0345eb6, 32'h40b827c4} /* (13, 12, 12) {real, imag} */,
  {32'h4002f943, 32'h4061cecd} /* (13, 12, 11) {real, imag} */,
  {32'hbf86fee3, 32'h406b6c76} /* (13, 12, 10) {real, imag} */,
  {32'hc10cd18c, 32'h40df6170} /* (13, 12, 9) {real, imag} */,
  {32'hc00ca583, 32'h40f0aa6f} /* (13, 12, 8) {real, imag} */,
  {32'hc03757c8, 32'h402bed9c} /* (13, 12, 7) {real, imag} */,
  {32'hc0fc6172, 32'hc0dd96df} /* (13, 12, 6) {real, imag} */,
  {32'hc12af485, 32'hbfc67e2a} /* (13, 12, 5) {real, imag} */,
  {32'hc11043b9, 32'h3fc5db19} /* (13, 12, 4) {real, imag} */,
  {32'h3ef5b258, 32'hbf812b48} /* (13, 12, 3) {real, imag} */,
  {32'h40918854, 32'h3e897bcc} /* (13, 12, 2) {real, imag} */,
  {32'h3ff68b42, 32'h3eca84c0} /* (13, 12, 1) {real, imag} */,
  {32'h402c1f50, 32'hbec36994} /* (13, 12, 0) {real, imag} */,
  {32'h4061a39a, 32'h4002c462} /* (13, 11, 15) {real, imag} */,
  {32'h410d5328, 32'h401ff13e} /* (13, 11, 14) {real, imag} */,
  {32'h3fd8f499, 32'hbf0aaa1c} /* (13, 11, 13) {real, imag} */,
  {32'hc0496f6e, 32'h3f9803c1} /* (13, 11, 12) {real, imag} */,
  {32'h3f3bcbd0, 32'h3fb3e21e} /* (13, 11, 11) {real, imag} */,
  {32'h4041ac86, 32'h40dd15f2} /* (13, 11, 10) {real, imag} */,
  {32'hbf92608c, 32'h400620c5} /* (13, 11, 9) {real, imag} */,
  {32'hc03ad1e1, 32'hc04122f1} /* (13, 11, 8) {real, imag} */,
  {32'hbfaa337e, 32'hbfbe0a85} /* (13, 11, 7) {real, imag} */,
  {32'hc08209ee, 32'h40801241} /* (13, 11, 6) {real, imag} */,
  {32'hc090ff58, 32'h41118e30} /* (13, 11, 5) {real, imag} */,
  {32'hbf811530, 32'h4075e924} /* (13, 11, 4) {real, imag} */,
  {32'h3f6dd3a6, 32'hbf91d8c5} /* (13, 11, 3) {real, imag} */,
  {32'h3e910617, 32'h40744e9e} /* (13, 11, 2) {real, imag} */,
  {32'hbff09708, 32'h40d09002} /* (13, 11, 1) {real, imag} */,
  {32'hc00c49d8, 32'h3fa7f5b8} /* (13, 11, 0) {real, imag} */,
  {32'hbe97507c, 32'h3f8351bb} /* (13, 10, 15) {real, imag} */,
  {32'hbf5f5688, 32'h3fd4f2ce} /* (13, 10, 14) {real, imag} */,
  {32'hbfb67e58, 32'h40215065} /* (13, 10, 13) {real, imag} */,
  {32'hbeb8597c, 32'h3e4f0517} /* (13, 10, 12) {real, imag} */,
  {32'h3faf6ab2, 32'hbdbeb0e0} /* (13, 10, 11) {real, imag} */,
  {32'h3fc5caf1, 32'h4021c351} /* (13, 10, 10) {real, imag} */,
  {32'h3f5c66c0, 32'h3fbe5b0f} /* (13, 10, 9) {real, imag} */,
  {32'hbfe96942, 32'hbea3e9c0} /* (13, 10, 8) {real, imag} */,
  {32'h3e528470, 32'hbf88c548} /* (13, 10, 7) {real, imag} */,
  {32'hbf01b3a0, 32'h3f859d32} /* (13, 10, 6) {real, imag} */,
  {32'hc09f4267, 32'hc01812c6} /* (13, 10, 5) {real, imag} */,
  {32'hc0a441ff, 32'hbfe606f8} /* (13, 10, 4) {real, imag} */,
  {32'hbf76f9d8, 32'hc03da87a} /* (13, 10, 3) {real, imag} */,
  {32'hc0566884, 32'hbf851b10} /* (13, 10, 2) {real, imag} */,
  {32'hc09b71a3, 32'hbd4729c0} /* (13, 10, 1) {real, imag} */,
  {32'hbfcbdb2f, 32'h3f011c08} /* (13, 10, 0) {real, imag} */,
  {32'hbf6b1f84, 32'h3dbaff30} /* (13, 9, 15) {real, imag} */,
  {32'hc00113ed, 32'hbf91aee7} /* (13, 9, 14) {real, imag} */,
  {32'hbf92a9e1, 32'hbfb12103} /* (13, 9, 13) {real, imag} */,
  {32'h3eeddbf2, 32'hbebef9f8} /* (13, 9, 12) {real, imag} */,
  {32'h3fb6becb, 32'h3fdd4205} /* (13, 9, 11) {real, imag} */,
  {32'hbede6a2a, 32'hbf4ff264} /* (13, 9, 10) {real, imag} */,
  {32'h3faa19af, 32'hbfca78b5} /* (13, 9, 9) {real, imag} */,
  {32'h3f8cf930, 32'hbfb45090} /* (13, 9, 8) {real, imag} */,
  {32'h40160a1b, 32'hc00e643e} /* (13, 9, 7) {real, imag} */,
  {32'h3fbe6456, 32'hbf34257c} /* (13, 9, 6) {real, imag} */,
  {32'h3e33dcb4, 32'hbf92ee07} /* (13, 9, 5) {real, imag} */,
  {32'hc041123e, 32'h3fb2b5bc} /* (13, 9, 4) {real, imag} */,
  {32'hc02c9e96, 32'h400daf91} /* (13, 9, 3) {real, imag} */,
  {32'hbf17e2ce, 32'h3fb27352} /* (13, 9, 2) {real, imag} */,
  {32'h3fcf7d10, 32'h3ff499f5} /* (13, 9, 1) {real, imag} */,
  {32'h3f7ac783, 32'h3f8c031f} /* (13, 9, 0) {real, imag} */,
  {32'h3f05e647, 32'h3d997560} /* (13, 8, 15) {real, imag} */,
  {32'hbfd3ec9e, 32'h3f6c4c57} /* (13, 8, 14) {real, imag} */,
  {32'hbf8cd3f8, 32'hbf397728} /* (13, 8, 13) {real, imag} */,
  {32'hbf0fcb10, 32'hbf65e948} /* (13, 8, 12) {real, imag} */,
  {32'h3f87e420, 32'hbfcbe974} /* (13, 8, 11) {real, imag} */,
  {32'hbf72957c, 32'hbf606a80} /* (13, 8, 10) {real, imag} */,
  {32'h3f0f9488, 32'h40082bd0} /* (13, 8, 9) {real, imag} */,
  {32'hbe451610, 32'h3f90f1f8} /* (13, 8, 8) {real, imag} */,
  {32'hbf0192d8, 32'h3f71e660} /* (13, 8, 7) {real, imag} */,
  {32'hbf99436b, 32'h3f5cce50} /* (13, 8, 6) {real, imag} */,
  {32'h3faad803, 32'hbe9ddec8} /* (13, 8, 5) {real, imag} */,
  {32'h400df912, 32'hbe9469b0} /* (13, 8, 4) {real, imag} */,
  {32'h3f5a6f44, 32'h403d1e45} /* (13, 8, 3) {real, imag} */,
  {32'h3fa77f32, 32'h3fb70aca} /* (13, 8, 2) {real, imag} */,
  {32'hbf032764, 32'hbf9d4978} /* (13, 8, 1) {real, imag} */,
  {32'h3f2b435c, 32'h3e3df508} /* (13, 8, 0) {real, imag} */,
  {32'hbf2fcbd4, 32'hbebd80f4} /* (13, 7, 15) {real, imag} */,
  {32'hc079322d, 32'hc02c30d0} /* (13, 7, 14) {real, imag} */,
  {32'hbfe49d59, 32'hbfdaaced} /* (13, 7, 13) {real, imag} */,
  {32'hbfd079da, 32'h400e52f1} /* (13, 7, 12) {real, imag} */,
  {32'hbe177ef8, 32'h3fd131ab} /* (13, 7, 11) {real, imag} */,
  {32'hbfa85cea, 32'h3f11a304} /* (13, 7, 10) {real, imag} */,
  {32'hc00cf5a2, 32'h3fb0033d} /* (13, 7, 9) {real, imag} */,
  {32'hbff4a280, 32'hbf8fb188} /* (13, 7, 8) {real, imag} */,
  {32'hbe8621c8, 32'h3e713098} /* (13, 7, 7) {real, imag} */,
  {32'h3ee56c88, 32'h3f587c5c} /* (13, 7, 6) {real, imag} */,
  {32'hbfcfca6a, 32'hbeb06fec} /* (13, 7, 5) {real, imag} */,
  {32'hbf1c6da0, 32'hbfab1b8a} /* (13, 7, 4) {real, imag} */,
  {32'h3fe15f2c, 32'hbf117b73} /* (13, 7, 3) {real, imag} */,
  {32'h402958fc, 32'h3fb7d89c} /* (13, 7, 2) {real, imag} */,
  {32'hbd9d43d8, 32'h3fdffd3d} /* (13, 7, 1) {real, imag} */,
  {32'h3e4acb64, 32'hbd0f2020} /* (13, 7, 0) {real, imag} */,
  {32'h3fe8d0d7, 32'hbf8f1abb} /* (13, 6, 15) {real, imag} */,
  {32'h40547842, 32'h400743f3} /* (13, 6, 14) {real, imag} */,
  {32'h3fa1256c, 32'h3ffc1a32} /* (13, 6, 13) {real, imag} */,
  {32'h3f049282, 32'h3cde4878} /* (13, 6, 12) {real, imag} */,
  {32'h3d0737c0, 32'hbf97bffe} /* (13, 6, 11) {real, imag} */,
  {32'h3f14424a, 32'hc03ee4df} /* (13, 6, 10) {real, imag} */,
  {32'hbd471c40, 32'hbf7e1e2a} /* (13, 6, 9) {real, imag} */,
  {32'h3f96fd82, 32'h4061893e} /* (13, 6, 8) {real, imag} */,
  {32'h40249c38, 32'h3f9511dc} /* (13, 6, 7) {real, imag} */,
  {32'h3f699dd0, 32'hc08a75ac} /* (13, 6, 6) {real, imag} */,
  {32'h3f8bab8f, 32'hbf32590a} /* (13, 6, 5) {real, imag} */,
  {32'hc06f9e4a, 32'h3e83c9c0} /* (13, 6, 4) {real, imag} */,
  {32'hc047a560, 32'h3f93e848} /* (13, 6, 3) {real, imag} */,
  {32'hbfd3f569, 32'h3f98e360} /* (13, 6, 2) {real, imag} */,
  {32'hc021628e, 32'hc074890f} /* (13, 6, 1) {real, imag} */,
  {32'hbfd93b67, 32'hc027ea38} /* (13, 6, 0) {real, imag} */,
  {32'hbe8805f0, 32'hc08dec8c} /* (13, 5, 15) {real, imag} */,
  {32'h40477286, 32'hc0b66cb9} /* (13, 5, 14) {real, imag} */,
  {32'hbf05469e, 32'h4044d386} /* (13, 5, 13) {real, imag} */,
  {32'hc0a1128d, 32'h408e4acd} /* (13, 5, 12) {real, imag} */,
  {32'hc03ae89c, 32'h40ee8838} /* (13, 5, 11) {real, imag} */,
  {32'h3f262550, 32'h409aa3f2} /* (13, 5, 10) {real, imag} */,
  {32'hc04766a2, 32'h401eae43} /* (13, 5, 9) {real, imag} */,
  {32'h3f475114, 32'h4016f107} /* (13, 5, 8) {real, imag} */,
  {32'h40141cce, 32'hbf73386a} /* (13, 5, 7) {real, imag} */,
  {32'hc0146840, 32'hbf99d72b} /* (13, 5, 6) {real, imag} */,
  {32'hc0815834, 32'hc03871ee} /* (13, 5, 5) {real, imag} */,
  {32'hc0acf4bb, 32'hc0147862} /* (13, 5, 4) {real, imag} */,
  {32'hbf134b46, 32'hbfef7705} /* (13, 5, 3) {real, imag} */,
  {32'h3eccd631, 32'hbf792ac0} /* (13, 5, 2) {real, imag} */,
  {32'h3f976b6c, 32'hc098e34a} /* (13, 5, 1) {real, imag} */,
  {32'h3b743400, 32'hbff8e82c} /* (13, 5, 0) {real, imag} */,
  {32'h40b43022, 32'h3fc8a6d0} /* (13, 4, 15) {real, imag} */,
  {32'hc0168ae1, 32'h401c3134} /* (13, 4, 14) {real, imag} */,
  {32'hc1137d74, 32'hbec1b7e0} /* (13, 4, 13) {real, imag} */,
  {32'hc060215e, 32'h4007287d} /* (13, 4, 12) {real, imag} */,
  {32'hc04e1039, 32'hc0c0ae6e} /* (13, 4, 11) {real, imag} */,
  {32'hbfc0f7d1, 32'hc00b612a} /* (13, 4, 10) {real, imag} */,
  {32'h3f189108, 32'hbf88d152} /* (13, 4, 9) {real, imag} */,
  {32'hc108d1f7, 32'hc0c70d3d} /* (13, 4, 8) {real, imag} */,
  {32'hc06a0ce8, 32'hc0b3cca4} /* (13, 4, 7) {real, imag} */,
  {32'h4051b3d4, 32'h3e5b2580} /* (13, 4, 6) {real, imag} */,
  {32'h40b1f11e, 32'h401f2ea3} /* (13, 4, 5) {real, imag} */,
  {32'h3ff4d5c8, 32'h3febe58f} /* (13, 4, 4) {real, imag} */,
  {32'hbf9e837e, 32'h3f25e388} /* (13, 4, 3) {real, imag} */,
  {32'h40b56b54, 32'h3f4a6442} /* (13, 4, 2) {real, imag} */,
  {32'h4015faff, 32'h40285ee6} /* (13, 4, 1) {real, imag} */,
  {32'h3f9191a7, 32'h4012cbe8} /* (13, 4, 0) {real, imag} */,
  {32'hc0994dc0, 32'hbee99b38} /* (13, 3, 15) {real, imag} */,
  {32'hc0f4d63e, 32'hc085bc62} /* (13, 3, 14) {real, imag} */,
  {32'hc0548dbb, 32'h401ff014} /* (13, 3, 13) {real, imag} */,
  {32'h40dd8fe9, 32'h40a8a9fa} /* (13, 3, 12) {real, imag} */,
  {32'h3ff94a5e, 32'hc03b1f57} /* (13, 3, 11) {real, imag} */,
  {32'hc0cea2f8, 32'h400f38e5} /* (13, 3, 10) {real, imag} */,
  {32'hc1331a6c, 32'h40d5e709} /* (13, 3, 9) {real, imag} */,
  {32'hc00f59c8, 32'h3fd80d4f} /* (13, 3, 8) {real, imag} */,
  {32'hbfb85479, 32'hbfc98c11} /* (13, 3, 7) {real, imag} */,
  {32'h3fcbe87c, 32'hbf7424b0} /* (13, 3, 6) {real, imag} */,
  {32'h403edadf, 32'hbf848f7d} /* (13, 3, 5) {real, imag} */,
  {32'h3f39f0c7, 32'hc0c54b78} /* (13, 3, 4) {real, imag} */,
  {32'hbf04a34a, 32'hc10062e8} /* (13, 3, 3) {real, imag} */,
  {32'hc0073209, 32'h3f1bb38d} /* (13, 3, 2) {real, imag} */,
  {32'hc0b0cdd2, 32'h407632d2} /* (13, 3, 1) {real, imag} */,
  {32'h408c20df, 32'h3feeff8a} /* (13, 3, 0) {real, imag} */,
  {32'h40ad3dac, 32'h3fe8561a} /* (13, 2, 15) {real, imag} */,
  {32'h402ec3a4, 32'h4061473c} /* (13, 2, 14) {real, imag} */,
  {32'h4092be36, 32'hc0bc18e8} /* (13, 2, 13) {real, imag} */,
  {32'h40eef218, 32'hbfbab0f6} /* (13, 2, 12) {real, imag} */,
  {32'hbfb3044e, 32'hc02f3f8c} /* (13, 2, 11) {real, imag} */,
  {32'h40a6c569, 32'hc01e1a48} /* (13, 2, 10) {real, imag} */,
  {32'h40ac97c2, 32'hc0488ebe} /* (13, 2, 9) {real, imag} */,
  {32'hc0423772, 32'hc08e05d2} /* (13, 2, 8) {real, imag} */,
  {32'hc059efd0, 32'hbf5d1088} /* (13, 2, 7) {real, imag} */,
  {32'hbfc742d0, 32'h406ec3b1} /* (13, 2, 6) {real, imag} */,
  {32'h408a8c76, 32'hbed60c50} /* (13, 2, 5) {real, imag} */,
  {32'h40d56008, 32'hc00f7d01} /* (13, 2, 4) {real, imag} */,
  {32'h4017285e, 32'h3fa47788} /* (13, 2, 3) {real, imag} */,
  {32'hc0a67351, 32'h3fc18114} /* (13, 2, 2) {real, imag} */,
  {32'hbf9ae904, 32'h3f923988} /* (13, 2, 1) {real, imag} */,
  {32'hc00da770, 32'h404ab8db} /* (13, 2, 0) {real, imag} */,
  {32'hc1562156, 32'h3ffed4d0} /* (13, 1, 15) {real, imag} */,
  {32'hc0394340, 32'h408a58ea} /* (13, 1, 14) {real, imag} */,
  {32'h414675bf, 32'hc066ef62} /* (13, 1, 13) {real, imag} */,
  {32'h3eb3d899, 32'hbf7722b0} /* (13, 1, 12) {real, imag} */,
  {32'h3fcccf26, 32'hc07cc1a8} /* (13, 1, 11) {real, imag} */,
  {32'h3e559230, 32'hc0c4beec} /* (13, 1, 10) {real, imag} */,
  {32'hc0bedf5b, 32'hc0885cd2} /* (13, 1, 9) {real, imag} */,
  {32'h3ee99467, 32'hc0bfc9d0} /* (13, 1, 8) {real, imag} */,
  {32'h410446b0, 32'h40d4f368} /* (13, 1, 7) {real, imag} */,
  {32'h40b460cc, 32'h4129747d} /* (13, 1, 6) {real, imag} */,
  {32'h40c41600, 32'h3f9c7b72} /* (13, 1, 5) {real, imag} */,
  {32'h4112c66d, 32'h3f0fde82} /* (13, 1, 4) {real, imag} */,
  {32'hbf103cb8, 32'h40532bf3} /* (13, 1, 3) {real, imag} */,
  {32'hc0df82c0, 32'h400ba57e} /* (13, 1, 2) {real, imag} */,
  {32'h40275de3, 32'h40b08ebb} /* (13, 1, 1) {real, imag} */,
  {32'hbfde9226, 32'hc004624b} /* (13, 1, 0) {real, imag} */,
  {32'h401f79f8, 32'h3e033b68} /* (13, 0, 15) {real, imag} */,
  {32'h40c83d92, 32'hc033d667} /* (13, 0, 14) {real, imag} */,
  {32'hc10e5195, 32'h4091bf7d} /* (13, 0, 13) {real, imag} */,
  {32'hc198f436, 32'h4101bc4e} /* (13, 0, 12) {real, imag} */,
  {32'hbe323c60, 32'h413f7f12} /* (13, 0, 11) {real, imag} */,
  {32'h40d8c476, 32'h4060d794} /* (13, 0, 10) {real, imag} */,
  {32'hc048d1a0, 32'h40906081} /* (13, 0, 9) {real, imag} */,
  {32'hc01e1339, 32'h403eaf82} /* (13, 0, 8) {real, imag} */,
  {32'h41500a76, 32'h40de48c2} /* (13, 0, 7) {real, imag} */,
  {32'h3f072472, 32'hbf479a08} /* (13, 0, 6) {real, imag} */,
  {32'hbe345e38, 32'hc097bab6} /* (13, 0, 5) {real, imag} */,
  {32'h41122348, 32'h408ba01f} /* (13, 0, 4) {real, imag} */,
  {32'h40b185b2, 32'h41080d6d} /* (13, 0, 3) {real, imag} */,
  {32'h40bda81a, 32'h406fe571} /* (13, 0, 2) {real, imag} */,
  {32'h40e433d0, 32'h4011f49a} /* (13, 0, 1) {real, imag} */,
  {32'h4084b746, 32'h3ec7d8c4} /* (13, 0, 0) {real, imag} */,
  {32'h4028d9fe, 32'hbf6655b8} /* (12, 15, 15) {real, imag} */,
  {32'h3f0c1dc8, 32'hbdad1020} /* (12, 15, 14) {real, imag} */,
  {32'hc0e6e292, 32'hc039b8b2} /* (12, 15, 13) {real, imag} */,
  {32'hc0d86470, 32'h3f84ed48} /* (12, 15, 12) {real, imag} */,
  {32'hbfa330e7, 32'hbf1b93dc} /* (12, 15, 11) {real, imag} */,
  {32'hc0645fd2, 32'hc034f680} /* (12, 15, 10) {real, imag} */,
  {32'h40954079, 32'h4016425c} /* (12, 15, 9) {real, imag} */,
  {32'h409289e1, 32'h409cb435} /* (12, 15, 8) {real, imag} */,
  {32'hbff29420, 32'h40f1b7db} /* (12, 15, 7) {real, imag} */,
  {32'hc045582c, 32'h40e20c0a} /* (12, 15, 6) {real, imag} */,
  {32'h3fb8322e, 32'h40cd1586} /* (12, 15, 5) {real, imag} */,
  {32'h40a3ac42, 32'h409cb276} /* (12, 15, 4) {real, imag} */,
  {32'h40abd252, 32'hc01fa9c0} /* (12, 15, 3) {real, imag} */,
  {32'hc031cc5c, 32'hc1027b90} /* (12, 15, 2) {real, imag} */,
  {32'hc0bfe546, 32'hc08369c3} /* (12, 15, 1) {real, imag} */,
  {32'hc08d1234, 32'hc096afa2} /* (12, 15, 0) {real, imag} */,
  {32'hc088d882, 32'h3ee7c252} /* (12, 14, 15) {real, imag} */,
  {32'hc0941867, 32'hbf95fb8e} /* (12, 14, 14) {real, imag} */,
  {32'hbf1be394, 32'h3f04cc72} /* (12, 14, 13) {real, imag} */,
  {32'hc00b0e50, 32'hbdc024e0} /* (12, 14, 12) {real, imag} */,
  {32'hc09ff407, 32'hbffa8ff0} /* (12, 14, 11) {real, imag} */,
  {32'hbf6c9300, 32'h3ff481cc} /* (12, 14, 10) {real, imag} */,
  {32'hc11832be, 32'h4032b426} /* (12, 14, 9) {real, imag} */,
  {32'hc0aafae1, 32'h40d243d2} /* (12, 14, 8) {real, imag} */,
  {32'hc08651ec, 32'h411d610d} /* (12, 14, 7) {real, imag} */,
  {32'h40006190, 32'h402a7d6d} /* (12, 14, 6) {real, imag} */,
  {32'h403689df, 32'h400a64c6} /* (12, 14, 5) {real, imag} */,
  {32'hc039bdd6, 32'hbe5216c0} /* (12, 14, 4) {real, imag} */,
  {32'hc102bda5, 32'hc0621b6a} /* (12, 14, 3) {real, imag} */,
  {32'hc02e1644, 32'hbf99e220} /* (12, 14, 2) {real, imag} */,
  {32'h40578dfe, 32'h403b3cbc} /* (12, 14, 1) {real, imag} */,
  {32'h40a08914, 32'h3ff74a9e} /* (12, 14, 0) {real, imag} */,
  {32'h3f39600f, 32'hbec9349c} /* (12, 13, 15) {real, imag} */,
  {32'h3fd50078, 32'hbf101700} /* (12, 13, 14) {real, imag} */,
  {32'h407f0cce, 32'hbff974ac} /* (12, 13, 13) {real, imag} */,
  {32'hc02f2c97, 32'h3f586210} /* (12, 13, 12) {real, imag} */,
  {32'hbdb46900, 32'h40049d4c} /* (12, 13, 11) {real, imag} */,
  {32'h40a6c27d, 32'h40219922} /* (12, 13, 10) {real, imag} */,
  {32'h3fe4c40c, 32'h3fb04842} /* (12, 13, 9) {real, imag} */,
  {32'h400dc3e3, 32'h40247197} /* (12, 13, 8) {real, imag} */,
  {32'h408faf76, 32'hc064034f} /* (12, 13, 7) {real, imag} */,
  {32'h40a71e42, 32'h3f37c434} /* (12, 13, 6) {real, imag} */,
  {32'hbfd28df9, 32'h40b06f97} /* (12, 13, 5) {real, imag} */,
  {32'hc08e611b, 32'hbff698b1} /* (12, 13, 4) {real, imag} */,
  {32'h3fd48dc1, 32'hc08c7007} /* (12, 13, 3) {real, imag} */,
  {32'h3fa0043d, 32'hc08566d4} /* (12, 13, 2) {real, imag} */,
  {32'hc0d7b8b6, 32'hbfc730a2} /* (12, 13, 1) {real, imag} */,
  {32'h3f4286dc, 32'hbffea9dc} /* (12, 13, 0) {real, imag} */,
  {32'h3e4d3468, 32'hbfac174a} /* (12, 12, 15) {real, imag} */,
  {32'h4035d777, 32'hc04fa21a} /* (12, 12, 14) {real, imag} */,
  {32'h4088cbd0, 32'h3fb17094} /* (12, 12, 13) {real, imag} */,
  {32'h40db9117, 32'hbf3de27f} /* (12, 12, 12) {real, imag} */,
  {32'hc013339a, 32'hbf0b6667} /* (12, 12, 11) {real, imag} */,
  {32'hc0003390, 32'h3e0f0708} /* (12, 12, 10) {real, imag} */,
  {32'hbfccbdcf, 32'hc0503ea3} /* (12, 12, 9) {real, imag} */,
  {32'hbf9f4ba4, 32'h3dd121e8} /* (12, 12, 8) {real, imag} */,
  {32'h3fe1b439, 32'hc015dd33} /* (12, 12, 7) {real, imag} */,
  {32'hc0262673, 32'hbfa76200} /* (12, 12, 6) {real, imag} */,
  {32'hc0846a53, 32'h4008e6ad} /* (12, 12, 5) {real, imag} */,
  {32'hbefc5cdc, 32'hbd5736a0} /* (12, 12, 4) {real, imag} */,
  {32'h3f9b8e63, 32'h401fc226} /* (12, 12, 3) {real, imag} */,
  {32'h400d53dd, 32'h40ab86c1} /* (12, 12, 2) {real, imag} */,
  {32'h40c16b74, 32'hbfd9bf43} /* (12, 12, 1) {real, imag} */,
  {32'h407e89d7, 32'hc0599dd6} /* (12, 12, 0) {real, imag} */,
  {32'h3dbe78f0, 32'h3e9c4f62} /* (12, 11, 15) {real, imag} */,
  {32'h40008749, 32'hbfd17def} /* (12, 11, 14) {real, imag} */,
  {32'hbf0a45bc, 32'h402786d6} /* (12, 11, 13) {real, imag} */,
  {32'hc0106354, 32'h4033dfc0} /* (12, 11, 12) {real, imag} */,
  {32'hbe1126f0, 32'hbdaffcf0} /* (12, 11, 11) {real, imag} */,
  {32'h400c1ae2, 32'hbdc79d30} /* (12, 11, 10) {real, imag} */,
  {32'h404b23ac, 32'h405ae024} /* (12, 11, 9) {real, imag} */,
  {32'h40979169, 32'h4075650e} /* (12, 11, 8) {real, imag} */,
  {32'h403b9631, 32'h4017a914} /* (12, 11, 7) {real, imag} */,
  {32'hc0836d3d, 32'h3efb5920} /* (12, 11, 6) {real, imag} */,
  {32'hbf469fa8, 32'hc06fd8d2} /* (12, 11, 5) {real, imag} */,
  {32'h40957875, 32'hc10245d6} /* (12, 11, 4) {real, imag} */,
  {32'h3fcbc4f2, 32'hc0431aea} /* (12, 11, 3) {real, imag} */,
  {32'hbff95b24, 32'hbf675e65} /* (12, 11, 2) {real, imag} */,
  {32'hc0fcd0c5, 32'hc028055f} /* (12, 11, 1) {real, imag} */,
  {32'hc0793a9c, 32'hbecab364} /* (12, 11, 0) {real, imag} */,
  {32'hbf2d5406, 32'h3f399609} /* (12, 10, 15) {real, imag} */,
  {32'hc06275de, 32'hbf8162a0} /* (12, 10, 14) {real, imag} */,
  {32'hc0a0f6be, 32'hc086ce39} /* (12, 10, 13) {real, imag} */,
  {32'hc08712a2, 32'hc06173e6} /* (12, 10, 12) {real, imag} */,
  {32'hc0317948, 32'hbe278c60} /* (12, 10, 11) {real, imag} */,
  {32'hc0878d29, 32'hbfd95fd4} /* (12, 10, 10) {real, imag} */,
  {32'hc06f5a09, 32'hc0548625} /* (12, 10, 9) {real, imag} */,
  {32'h400a2bfe, 32'hc01868da} /* (12, 10, 8) {real, imag} */,
  {32'h40344219, 32'h402b4208} /* (12, 10, 7) {real, imag} */,
  {32'h4039ad94, 32'h3f80e10e} /* (12, 10, 6) {real, imag} */,
  {32'hbf0f1132, 32'hc0063ad8} /* (12, 10, 5) {real, imag} */,
  {32'hbe105d68, 32'hc0829c46} /* (12, 10, 4) {real, imag} */,
  {32'h4012acf8, 32'hc0682e68} /* (12, 10, 3) {real, imag} */,
  {32'h4056eb1a, 32'hc028e7ca} /* (12, 10, 2) {real, imag} */,
  {32'hbf2a9962, 32'hc0648162} /* (12, 10, 1) {real, imag} */,
  {32'hbf1b7aa2, 32'hbfe023c8} /* (12, 10, 0) {real, imag} */,
  {32'h3eef46dc, 32'h3ff40c98} /* (12, 9, 15) {real, imag} */,
  {32'h3d1b23e0, 32'h4023b415} /* (12, 9, 14) {real, imag} */,
  {32'hbfde1b6f, 32'h3fc259b9} /* (12, 9, 13) {real, imag} */,
  {32'hc02b4fde, 32'h4026e207} /* (12, 9, 12) {real, imag} */,
  {32'hbfced358, 32'h3fc93893} /* (12, 9, 11) {real, imag} */,
  {32'h3fa321eb, 32'hbea335b0} /* (12, 9, 10) {real, imag} */,
  {32'hbe8119e8, 32'hbf534b86} /* (12, 9, 9) {real, imag} */,
  {32'hbfe2e01e, 32'h3f37ec64} /* (12, 9, 8) {real, imag} */,
  {32'h3fb6cfaa, 32'h4006599d} /* (12, 9, 7) {real, imag} */,
  {32'h3fae8bcd, 32'h404c8bf4} /* (12, 9, 6) {real, imag} */,
  {32'h3f78411c, 32'h3f2628ec} /* (12, 9, 5) {real, imag} */,
  {32'h3fe73389, 32'hbe24c2d8} /* (12, 9, 4) {real, imag} */,
  {32'h3fcd9a56, 32'h4016de76} /* (12, 9, 3) {real, imag} */,
  {32'h40244cdc, 32'hbdf832b0} /* (12, 9, 2) {real, imag} */,
  {32'h3ec755dc, 32'hbf1d1161} /* (12, 9, 1) {real, imag} */,
  {32'hbead2bae, 32'hbe39f9d4} /* (12, 9, 0) {real, imag} */,
  {32'hbf58fca8, 32'h3f5fae44} /* (12, 8, 15) {real, imag} */,
  {32'h3f2a9250, 32'h3f8f1a6e} /* (12, 8, 14) {real, imag} */,
  {32'h3ec578b4, 32'hbf565024} /* (12, 8, 13) {real, imag} */,
  {32'hc03de178, 32'hbfa57ec0} /* (12, 8, 12) {real, imag} */,
  {32'hbf4d4430, 32'hbf8c7ad0} /* (12, 8, 11) {real, imag} */,
  {32'hbfacb43f, 32'hbf54d854} /* (12, 8, 10) {real, imag} */,
  {32'hbfd7193d, 32'hbf3931aa} /* (12, 8, 9) {real, imag} */,
  {32'hbf72a1e8, 32'hbf4e1450} /* (12, 8, 8) {real, imag} */,
  {32'hc05e7bc6, 32'h3ff9870a} /* (12, 8, 7) {real, imag} */,
  {32'hc04c084d, 32'h3f86d1cc} /* (12, 8, 6) {real, imag} */,
  {32'hbe828948, 32'hbf1dd4fc} /* (12, 8, 5) {real, imag} */,
  {32'hbf2c6ee4, 32'hbd76d6e0} /* (12, 8, 4) {real, imag} */,
  {32'hbe8c34a4, 32'h3d84a1e0} /* (12, 8, 3) {real, imag} */,
  {32'h3ee36306, 32'hbea389e2} /* (12, 8, 2) {real, imag} */,
  {32'h3f9bf544, 32'hbe0c1ca0} /* (12, 8, 1) {real, imag} */,
  {32'h3f11f3cc, 32'hbf2226e2} /* (12, 8, 0) {real, imag} */,
  {32'hbfee302b, 32'hbe9e9710} /* (12, 7, 15) {real, imag} */,
  {32'hbf03faf2, 32'hbef5cc38} /* (12, 7, 14) {real, imag} */,
  {32'hbe4ca238, 32'hbf268d7e} /* (12, 7, 13) {real, imag} */,
  {32'h3f595e5f, 32'hc022e9d5} /* (12, 7, 12) {real, imag} */,
  {32'h3f84bba2, 32'hbfe5bda5} /* (12, 7, 11) {real, imag} */,
  {32'h3f0ec402, 32'hbef93308} /* (12, 7, 10) {real, imag} */,
  {32'h4020dcb8, 32'hbf19f552} /* (12, 7, 9) {real, imag} */,
  {32'h3fd18f7a, 32'hbca55780} /* (12, 7, 8) {real, imag} */,
  {32'hbed4a620, 32'h3f91aa0e} /* (12, 7, 7) {real, imag} */,
  {32'h3edfa554, 32'h3fd03e78} /* (12, 7, 6) {real, imag} */,
  {32'hbfd5f27e, 32'h406170e3} /* (12, 7, 5) {real, imag} */,
  {32'hbf8e4b41, 32'h4017f332} /* (12, 7, 4) {real, imag} */,
  {32'h3ef09e78, 32'h3f36617c} /* (12, 7, 3) {real, imag} */,
  {32'hbf0ad050, 32'h3e31b738} /* (12, 7, 2) {real, imag} */,
  {32'hbe46d528, 32'h3f1ace3f} /* (12, 7, 1) {real, imag} */,
  {32'hbf72737b, 32'hbe072c94} /* (12, 7, 0) {real, imag} */,
  {32'h3f97ae6d, 32'h3f31afa7} /* (12, 6, 15) {real, imag} */,
  {32'h3e8aa528, 32'hbf077870} /* (12, 6, 14) {real, imag} */,
  {32'hbf160f6c, 32'h3fa3b3f4} /* (12, 6, 13) {real, imag} */,
  {32'hc00698fe, 32'h4095313f} /* (12, 6, 12) {real, imag} */,
  {32'hc02f7012, 32'h4076a04a} /* (12, 6, 11) {real, imag} */,
  {32'h3f862d18, 32'h4082e8e5} /* (12, 6, 10) {real, imag} */,
  {32'h3fcf9096, 32'h401178f1} /* (12, 6, 9) {real, imag} */,
  {32'h3eb4c954, 32'h3e935d10} /* (12, 6, 8) {real, imag} */,
  {32'h404ffca3, 32'hc00ae632} /* (12, 6, 7) {real, imag} */,
  {32'h4017ca3e, 32'hc002f8c9} /* (12, 6, 6) {real, imag} */,
  {32'h3f0a6b92, 32'hc002b4d0} /* (12, 6, 5) {real, imag} */,
  {32'hbfbae697, 32'hbf9ff8fa} /* (12, 6, 4) {real, imag} */,
  {32'hc0c1fa62, 32'h3f5dd31a} /* (12, 6, 3) {real, imag} */,
  {32'hc08d8dc4, 32'h3bc80800} /* (12, 6, 2) {real, imag} */,
  {32'h3f61c2aa, 32'hc03b68c4} /* (12, 6, 1) {real, imag} */,
  {32'h3f961065, 32'hbf7ae5e5} /* (12, 6, 0) {real, imag} */,
  {32'hc0524d8a, 32'h400685bb} /* (12, 5, 15) {real, imag} */,
  {32'hc0031905, 32'h40221874} /* (12, 5, 14) {real, imag} */,
  {32'h3fe84a6c, 32'h3f224d6e} /* (12, 5, 13) {real, imag} */,
  {32'h402ce082, 32'hc0272f42} /* (12, 5, 12) {real, imag} */,
  {32'hc01c98c3, 32'hbfdb9b2e} /* (12, 5, 11) {real, imag} */,
  {32'hbff27934, 32'hbffe4019} /* (12, 5, 10) {real, imag} */,
  {32'h4066ebb0, 32'hbdebecc0} /* (12, 5, 9) {real, imag} */,
  {32'h409c3deb, 32'hc04108e2} /* (12, 5, 8) {real, imag} */,
  {32'h400a020d, 32'hc06d2686} /* (12, 5, 7) {real, imag} */,
  {32'h402240f4, 32'hc02794c0} /* (12, 5, 6) {real, imag} */,
  {32'hbf19984c, 32'hc0530756} /* (12, 5, 5) {real, imag} */,
  {32'hc0208808, 32'hc00eef14} /* (12, 5, 4) {real, imag} */,
  {32'hc0b020d0, 32'hbfabf5cb} /* (12, 5, 3) {real, imag} */,
  {32'hc0dc703d, 32'hc026b0d8} /* (12, 5, 2) {real, imag} */,
  {32'hc08db547, 32'hbfb030b2} /* (12, 5, 1) {real, imag} */,
  {32'hc09572c0, 32'hbf03534a} /* (12, 5, 0) {real, imag} */,
  {32'h3ff79f6d, 32'h3fc5aa56} /* (12, 4, 15) {real, imag} */,
  {32'h40b36eac, 32'hbfbb1244} /* (12, 4, 14) {real, imag} */,
  {32'h404d18b2, 32'hc049f7e6} /* (12, 4, 13) {real, imag} */,
  {32'h3f8050cc, 32'hbce398e0} /* (12, 4, 12) {real, imag} */,
  {32'hbf34bdc2, 32'h3fc53990} /* (12, 4, 11) {real, imag} */,
  {32'h401faef2, 32'h40291e70} /* (12, 4, 10) {real, imag} */,
  {32'hc086ee2e, 32'hbf0167e4} /* (12, 4, 9) {real, imag} */,
  {32'hc0c75278, 32'h3f6f6bb3} /* (12, 4, 8) {real, imag} */,
  {32'hc032d70a, 32'h401660b9} /* (12, 4, 7) {real, imag} */,
  {32'h40103705, 32'hc076b700} /* (12, 4, 6) {real, imag} */,
  {32'h403a5876, 32'hc08db666} /* (12, 4, 5) {real, imag} */,
  {32'hc02220e6, 32'hc042d660} /* (12, 4, 4) {real, imag} */,
  {32'hbe9fbe5c, 32'h3eaf3444} /* (12, 4, 3) {real, imag} */,
  {32'hbfea6116, 32'h3d81acc0} /* (12, 4, 2) {real, imag} */,
  {32'hc0c469c2, 32'hc067a7c6} /* (12, 4, 1) {real, imag} */,
  {32'hbe3d6fd0, 32'hc049bdba} /* (12, 4, 0) {real, imag} */,
  {32'hc0188a8d, 32'h4052b0b8} /* (12, 3, 15) {real, imag} */,
  {32'hbf957a54, 32'h3f4b8494} /* (12, 3, 14) {real, imag} */,
  {32'h3fb6bb0b, 32'h3f91face} /* (12, 3, 13) {real, imag} */,
  {32'hc094b5ea, 32'h3fb68304} /* (12, 3, 12) {real, imag} */,
  {32'h3e9f7c1c, 32'h3f7d97c7} /* (12, 3, 11) {real, imag} */,
  {32'h40b65077, 32'hbfe1caec} /* (12, 3, 10) {real, imag} */,
  {32'h3fd607c6, 32'hc06e211d} /* (12, 3, 9) {real, imag} */,
  {32'h40823f74, 32'hc04e6491} /* (12, 3, 8) {real, imag} */,
  {32'h4029a52f, 32'hc07ff065} /* (12, 3, 7) {real, imag} */,
  {32'hbff5fd9d, 32'h40a2cbd4} /* (12, 3, 6) {real, imag} */,
  {32'h403e48c0, 32'hbfb22e8c} /* (12, 3, 5) {real, imag} */,
  {32'h402cf490, 32'h3fa8d429} /* (12, 3, 4) {real, imag} */,
  {32'h400e29d2, 32'h40860d51} /* (12, 3, 3) {real, imag} */,
  {32'hbf0fe6ca, 32'hc06761c3} /* (12, 3, 2) {real, imag} */,
  {32'h3ef0e9a0, 32'hc043f353} /* (12, 3, 1) {real, imag} */,
  {32'hc03b696b, 32'hbfd53ce6} /* (12, 3, 0) {real, imag} */,
  {32'hc042d9ac, 32'h3f461807} /* (12, 2, 15) {real, imag} */,
  {32'hc01f9162, 32'h407c46c9} /* (12, 2, 14) {real, imag} */,
  {32'hc04657f0, 32'hbf812c51} /* (12, 2, 13) {real, imag} */,
  {32'hc0da5acc, 32'h401739b9} /* (12, 2, 12) {real, imag} */,
  {32'hc003dd30, 32'hc000bf1c} /* (12, 2, 11) {real, imag} */,
  {32'hc0926be5, 32'hc0d22297} /* (12, 2, 10) {real, imag} */,
  {32'h405b75b5, 32'hbfac76d0} /* (12, 2, 9) {real, imag} */,
  {32'h41010fbc, 32'h40a2266a} /* (12, 2, 8) {real, imag} */,
  {32'hbfa50717, 32'h40063403} /* (12, 2, 7) {real, imag} */,
  {32'h3f492936, 32'h4050c349} /* (12, 2, 6) {real, imag} */,
  {32'hc0801fe0, 32'h411b77de} /* (12, 2, 5) {real, imag} */,
  {32'hc0bc0209, 32'h41354a57} /* (12, 2, 4) {real, imag} */,
  {32'hc059ce30, 32'h4121b2c6} /* (12, 2, 3) {real, imag} */,
  {32'hbefd95d0, 32'h4113be08} /* (12, 2, 2) {real, imag} */,
  {32'h40b422d9, 32'h40a97ec6} /* (12, 2, 1) {real, imag} */,
  {32'hbf87bfae, 32'h4041d2fd} /* (12, 2, 0) {real, imag} */,
  {32'h40ca34fd, 32'hc0c17528} /* (12, 1, 15) {real, imag} */,
  {32'h40a3e66b, 32'hc0e540c2} /* (12, 1, 14) {real, imag} */,
  {32'h40182438, 32'h3f83e4a5} /* (12, 1, 13) {real, imag} */,
  {32'h40a12c60, 32'hc030770c} /* (12, 1, 12) {real, imag} */,
  {32'h408d4cac, 32'h3fd1d80a} /* (12, 1, 11) {real, imag} */,
  {32'hc027dd24, 32'hbf022b64} /* (12, 1, 10) {real, imag} */,
  {32'hbfe8a013, 32'hbe332578} /* (12, 1, 9) {real, imag} */,
  {32'h408c3f9b, 32'hc03c25e6} /* (12, 1, 8) {real, imag} */,
  {32'h40d4e06c, 32'hc1041038} /* (12, 1, 7) {real, imag} */,
  {32'hbb295a00, 32'hc0fdb4da} /* (12, 1, 6) {real, imag} */,
  {32'h40fae020, 32'hc103fa25} /* (12, 1, 5) {real, imag} */,
  {32'h41250b9c, 32'hc0bdc92e} /* (12, 1, 4) {real, imag} */,
  {32'h41211621, 32'hc0118ffc} /* (12, 1, 3) {real, imag} */,
  {32'h410f4637, 32'hbf8a5be4} /* (12, 1, 2) {real, imag} */,
  {32'h40c42e3a, 32'h405c1a22} /* (12, 1, 1) {real, imag} */,
  {32'h40733727, 32'h3faf5268} /* (12, 1, 0) {real, imag} */,
  {32'hc10168da, 32'hbf377a04} /* (12, 0, 15) {real, imag} */,
  {32'hc114c731, 32'h40d873ae} /* (12, 0, 14) {real, imag} */,
  {32'hbf7d5d12, 32'h40da243c} /* (12, 0, 13) {real, imag} */,
  {32'h40e13e3c, 32'h4087e1ee} /* (12, 0, 12) {real, imag} */,
  {32'hbfb9f728, 32'hc0184136} /* (12, 0, 11) {real, imag} */,
  {32'hc053c0e0, 32'hc08c80fa} /* (12, 0, 10) {real, imag} */,
  {32'h3f59a95e, 32'hc0070462} /* (12, 0, 9) {real, imag} */,
  {32'hc0b37fea, 32'hbe81c2b0} /* (12, 0, 8) {real, imag} */,
  {32'hbef149dc, 32'hbfa6f086} /* (12, 0, 7) {real, imag} */,
  {32'h410acf61, 32'hc0b00471} /* (12, 0, 6) {real, imag} */,
  {32'h40cbf716, 32'hbfe2ecf6} /* (12, 0, 5) {real, imag} */,
  {32'hc06b15df, 32'hc07400d6} /* (12, 0, 4) {real, imag} */,
  {32'hc05cc092, 32'hc09d2620} /* (12, 0, 3) {real, imag} */,
  {32'h3f88d412, 32'hbfc84b9e} /* (12, 0, 2) {real, imag} */,
  {32'hbfe5f2a2, 32'h408eb61d} /* (12, 0, 1) {real, imag} */,
  {32'hc0a0edde, 32'h40729e2c} /* (12, 0, 0) {real, imag} */,
  {32'hbf6a227e, 32'h3ee8abf0} /* (11, 15, 15) {real, imag} */,
  {32'h4053399f, 32'hc00363a7} /* (11, 15, 14) {real, imag} */,
  {32'h410917a2, 32'h3ff0b9eb} /* (11, 15, 13) {real, imag} */,
  {32'h406380a4, 32'hc04694d5} /* (11, 15, 12) {real, imag} */,
  {32'hbfe3f067, 32'hc08bf833} /* (11, 15, 11) {real, imag} */,
  {32'hc0a84c45, 32'hc0649778} /* (11, 15, 10) {real, imag} */,
  {32'hc122850a, 32'hc0ce837c} /* (11, 15, 9) {real, imag} */,
  {32'hbff51234, 32'hc0a899f5} /* (11, 15, 8) {real, imag} */,
  {32'h40264e02, 32'h3fb093ff} /* (11, 15, 7) {real, imag} */,
  {32'h4014f022, 32'h40c8892c} /* (11, 15, 6) {real, imag} */,
  {32'h40edd002, 32'h3ffb2c87} /* (11, 15, 5) {real, imag} */,
  {32'h405590c0, 32'hc01436e8} /* (11, 15, 4) {real, imag} */,
  {32'hbfc25008, 32'hc09e01e8} /* (11, 15, 3) {real, imag} */,
  {32'h3c29afc0, 32'hc07b6e31} /* (11, 15, 2) {real, imag} */,
  {32'h40b4f9f7, 32'hc054733a} /* (11, 15, 1) {real, imag} */,
  {32'h3ffd3f16, 32'hbf90e820} /* (11, 15, 0) {real, imag} */,
  {32'h40915eba, 32'h409033d9} /* (11, 14, 15) {real, imag} */,
  {32'h3ff7da14, 32'h40a241b8} /* (11, 14, 14) {real, imag} */,
  {32'hc0bcd78b, 32'h401f7e8f} /* (11, 14, 13) {real, imag} */,
  {32'hc0af812e, 32'h3d235398} /* (11, 14, 12) {real, imag} */,
  {32'h3f6754ac, 32'hc01d5dd2} /* (11, 14, 11) {real, imag} */,
  {32'hbff15626, 32'h3e9fc4a0} /* (11, 14, 10) {real, imag} */,
  {32'hc06e6e7a, 32'h3ea0b4a0} /* (11, 14, 9) {real, imag} */,
  {32'hc06d0050, 32'h400234ad} /* (11, 14, 8) {real, imag} */,
  {32'hbf7afbdc, 32'h3f2ccda4} /* (11, 14, 7) {real, imag} */,
  {32'hbea55044, 32'hc09283e4} /* (11, 14, 6) {real, imag} */,
  {32'hc0c2affa, 32'h406feaf4} /* (11, 14, 5) {real, imag} */,
  {32'h3e8d4ffc, 32'h408662be} /* (11, 14, 4) {real, imag} */,
  {32'h40adc114, 32'hc0691e09} /* (11, 14, 3) {real, imag} */,
  {32'h40f2d487, 32'hc0af0d1f} /* (11, 14, 2) {real, imag} */,
  {32'h4110b9ee, 32'hc08c0fca} /* (11, 14, 1) {real, imag} */,
  {32'h406df29a, 32'hbe368740} /* (11, 14, 0) {real, imag} */,
  {32'hbd162b58, 32'hc07fd71d} /* (11, 13, 15) {real, imag} */,
  {32'hbeb4aa00, 32'hbeaf0dca} /* (11, 13, 14) {real, imag} */,
  {32'hbec79298, 32'h402ec823} /* (11, 13, 13) {real, imag} */,
  {32'hc09619a0, 32'hc05bd93a} /* (11, 13, 12) {real, imag} */,
  {32'h3f8d0f84, 32'hc035d95e} /* (11, 13, 11) {real, imag} */,
  {32'h408045be, 32'h3fc22990} /* (11, 13, 10) {real, imag} */,
  {32'hbfee1b0a, 32'h40152776} /* (11, 13, 9) {real, imag} */,
  {32'hbf487980, 32'h3eab9e50} /* (11, 13, 8) {real, imag} */,
  {32'hbe47410c, 32'h3f2cd4f8} /* (11, 13, 7) {real, imag} */,
  {32'h3fbc620a, 32'h3fee3d98} /* (11, 13, 6) {real, imag} */,
  {32'h406adaca, 32'h4008caa8} /* (11, 13, 5) {real, imag} */,
  {32'h40529257, 32'h407641a6} /* (11, 13, 4) {real, imag} */,
  {32'h3f03442b, 32'h4037489c} /* (11, 13, 3) {real, imag} */,
  {32'hc08fb51a, 32'hbe9e9b28} /* (11, 13, 2) {real, imag} */,
  {32'h3ecadcc0, 32'h40428d12} /* (11, 13, 1) {real, imag} */,
  {32'h40868ee0, 32'hbfa0c09d} /* (11, 13, 0) {real, imag} */,
  {32'hbff11d1c, 32'h3f21c0e6} /* (11, 12, 15) {real, imag} */,
  {32'h3f462d62, 32'hbfe30f07} /* (11, 12, 14) {real, imag} */,
  {32'h4026580e, 32'hbff80cfd} /* (11, 12, 13) {real, imag} */,
  {32'h3ef32a4c, 32'hbefaf8e0} /* (11, 12, 12) {real, imag} */,
  {32'h401775e0, 32'hbf4bd04e} /* (11, 12, 11) {real, imag} */,
  {32'h3efb1f22, 32'hbfc724a4} /* (11, 12, 10) {real, imag} */,
  {32'h3f7cbdaf, 32'hbf8443b9} /* (11, 12, 9) {real, imag} */,
  {32'hbf500046, 32'hc0aa05c6} /* (11, 12, 8) {real, imag} */,
  {32'hbfb04fe2, 32'hc0b21380} /* (11, 12, 7) {real, imag} */,
  {32'h3fd6632c, 32'h3fa8b501} /* (11, 12, 6) {real, imag} */,
  {32'h3fa2a92e, 32'h3d1cd8e0} /* (11, 12, 5) {real, imag} */,
  {32'hbfda22b6, 32'hbe966e61} /* (11, 12, 4) {real, imag} */,
  {32'hc0237f2b, 32'h3fe26aad} /* (11, 12, 3) {real, imag} */,
  {32'hc01897c0, 32'h404933ae} /* (11, 12, 2) {real, imag} */,
  {32'hc08bb4f4, 32'h40ad10e8} /* (11, 12, 1) {real, imag} */,
  {32'hc01708f6, 32'h405dffbb} /* (11, 12, 0) {real, imag} */,
  {32'hbf4f813e, 32'hbf26097d} /* (11, 11, 15) {real, imag} */,
  {32'hbfcc4d62, 32'h3fdf1741} /* (11, 11, 14) {real, imag} */,
  {32'h40034004, 32'h40181658} /* (11, 11, 13) {real, imag} */,
  {32'h4029a1ec, 32'h406ce8e0} /* (11, 11, 12) {real, imag} */,
  {32'h3f01e3fc, 32'h3f8848fa} /* (11, 11, 11) {real, imag} */,
  {32'h3eb6ba6c, 32'hbf3ebaf8} /* (11, 11, 10) {real, imag} */,
  {32'hbc47fd80, 32'h3eb4176c} /* (11, 11, 9) {real, imag} */,
  {32'hc02c623e, 32'h3f960bca} /* (11, 11, 8) {real, imag} */,
  {32'hc088c94c, 32'hbfc93326} /* (11, 11, 7) {real, imag} */,
  {32'hc082c0ac, 32'hc049a00a} /* (11, 11, 6) {real, imag} */,
  {32'hc082dd79, 32'hc0799b3b} /* (11, 11, 5) {real, imag} */,
  {32'hbf892d80, 32'hbea34930} /* (11, 11, 4) {real, imag} */,
  {32'h3f001a3d, 32'h40688d86} /* (11, 11, 3) {real, imag} */,
  {32'h3fa81ad0, 32'hbe859ad0} /* (11, 11, 2) {real, imag} */,
  {32'h3f19b33c, 32'hc0247d40} /* (11, 11, 1) {real, imag} */,
  {32'hbece5fce, 32'hbd53df18} /* (11, 11, 0) {real, imag} */,
  {32'hbf8ee4b2, 32'h3ed14cc4} /* (11, 10, 15) {real, imag} */,
  {32'h3e0a0a44, 32'h3f5e5ca6} /* (11, 10, 14) {real, imag} */,
  {32'h3f6abf99, 32'hbf10d370} /* (11, 10, 13) {real, imag} */,
  {32'h3ffc7c98, 32'hbf87d278} /* (11, 10, 12) {real, imag} */,
  {32'h3fdee455, 32'hbecf42ec} /* (11, 10, 11) {real, imag} */,
  {32'h401afffe, 32'hbfaae22a} /* (11, 10, 10) {real, imag} */,
  {32'h400b1510, 32'hbe84db60} /* (11, 10, 9) {real, imag} */,
  {32'h3fe38da2, 32'h402b906f} /* (11, 10, 8) {real, imag} */,
  {32'h3f9299f1, 32'h3f50a5a5} /* (11, 10, 7) {real, imag} */,
  {32'h3eff8772, 32'h3f70a450} /* (11, 10, 6) {real, imag} */,
  {32'h403d3e6e, 32'h400af6a8} /* (11, 10, 5) {real, imag} */,
  {32'h40547f78, 32'h4066bfa7} /* (11, 10, 4) {real, imag} */,
  {32'h3d85b740, 32'hbeb31d58} /* (11, 10, 3) {real, imag} */,
  {32'hbf86187a, 32'hc003a0ac} /* (11, 10, 2) {real, imag} */,
  {32'hbf9f87b1, 32'hbf550a20} /* (11, 10, 1) {real, imag} */,
  {32'hc02f97f0, 32'h3e4c3f88} /* (11, 10, 0) {real, imag} */,
  {32'hbe62cd18, 32'hbed560cc} /* (11, 9, 15) {real, imag} */,
  {32'h3e991892, 32'hbf7d2d66} /* (11, 9, 14) {real, imag} */,
  {32'hbe8a36e8, 32'hbf1e65ef} /* (11, 9, 13) {real, imag} */,
  {32'h3e7add84, 32'hbe8eafae} /* (11, 9, 12) {real, imag} */,
  {32'h3f4e802c, 32'h3f6b1ebd} /* (11, 9, 11) {real, imag} */,
  {32'h3fb4849a, 32'hbf85cc37} /* (11, 9, 10) {real, imag} */,
  {32'h3fe2a704, 32'hbf876fb6} /* (11, 9, 9) {real, imag} */,
  {32'hbe294818, 32'hbd346ae0} /* (11, 9, 8) {real, imag} */,
  {32'hbf095a35, 32'h3e9ce86c} /* (11, 9, 7) {real, imag} */,
  {32'h3f0d77f8, 32'hbd96f278} /* (11, 9, 6) {real, imag} */,
  {32'h3ec9ae70, 32'h3f027e46} /* (11, 9, 5) {real, imag} */,
  {32'h3f847da0, 32'h3fa6ad16} /* (11, 9, 4) {real, imag} */,
  {32'hbffe0d2e, 32'hbea5cfac} /* (11, 9, 3) {real, imag} */,
  {32'hc01005f2, 32'hbfeca782} /* (11, 9, 2) {real, imag} */,
  {32'hbeb039fa, 32'hbfd5f102} /* (11, 9, 1) {real, imag} */,
  {32'h3e917dfa, 32'hbf33f134} /* (11, 9, 0) {real, imag} */,
  {32'hbd9b7290, 32'hbfa07de5} /* (11, 8, 15) {real, imag} */,
  {32'hbf3fa2f8, 32'hbf568ac6} /* (11, 8, 14) {real, imag} */,
  {32'h3ee4757c, 32'h3f8a7af8} /* (11, 8, 13) {real, imag} */,
  {32'h3ff43268, 32'hbf329b88} /* (11, 8, 12) {real, imag} */,
  {32'h3f4f6332, 32'hbf2f1012} /* (11, 8, 11) {real, imag} */,
  {32'h3f6909b2, 32'hbd173480} /* (11, 8, 10) {real, imag} */,
  {32'hbe42b550, 32'h3eb9c534} /* (11, 8, 9) {real, imag} */,
  {32'hbfba86ec, 32'hbd346c60} /* (11, 8, 8) {real, imag} */,
  {32'hbf85d611, 32'hbf72a968} /* (11, 8, 7) {real, imag} */,
  {32'hbf897f10, 32'hbfc74176} /* (11, 8, 6) {real, imag} */,
  {32'hbf5bfbc0, 32'hbfd86277} /* (11, 8, 5) {real, imag} */,
  {32'hbfa18bfc, 32'hbf26245e} /* (11, 8, 4) {real, imag} */,
  {32'hbfdea800, 32'hbf1c8a5a} /* (11, 8, 3) {real, imag} */,
  {32'hbfe83312, 32'h3d717650} /* (11, 8, 2) {real, imag} */,
  {32'hbe0b9614, 32'h3f79f6dc} /* (11, 8, 1) {real, imag} */,
  {32'h3f429d2c, 32'h3def1f40} /* (11, 8, 0) {real, imag} */,
  {32'h3f294bca, 32'hbf04d71c} /* (11, 7, 15) {real, imag} */,
  {32'h3f4c6a23, 32'h3e91a29c} /* (11, 7, 14) {real, imag} */,
  {32'h3f7b6d3c, 32'hbf9317aa} /* (11, 7, 13) {real, imag} */,
  {32'hbf377083, 32'hbe8705fe} /* (11, 7, 12) {real, imag} */,
  {32'hbf052568, 32'h3f54037d} /* (11, 7, 11) {real, imag} */,
  {32'hbe9b7010, 32'h3fa87fb5} /* (11, 7, 10) {real, imag} */,
  {32'hbfa92d64, 32'hbfb516e4} /* (11, 7, 9) {real, imag} */,
  {32'hbf76e042, 32'hc003b004} /* (11, 7, 8) {real, imag} */,
  {32'hbf7a341b, 32'hbfd89419} /* (11, 7, 7) {real, imag} */,
  {32'hbf14cbe4, 32'hbf9dc70c} /* (11, 7, 6) {real, imag} */,
  {32'h3fbe6bd0, 32'hbfb03f9f} /* (11, 7, 5) {real, imag} */,
  {32'h3f65692d, 32'hbfdecbca} /* (11, 7, 4) {real, imag} */,
  {32'hbcf12120, 32'hbf0d9032} /* (11, 7, 3) {real, imag} */,
  {32'h3f009916, 32'h3f5e4acd} /* (11, 7, 2) {real, imag} */,
  {32'h3f10ba55, 32'h3ec2c732} /* (11, 7, 1) {real, imag} */,
  {32'hbc363940, 32'h3e7248b6} /* (11, 7, 0) {real, imag} */,
  {32'hbfca40ee, 32'hbfd9c989} /* (11, 6, 15) {real, imag} */,
  {32'hbf8fe888, 32'h3e45a608} /* (11, 6, 14) {real, imag} */,
  {32'h3dc5b4c8, 32'h3fd24b46} /* (11, 6, 13) {real, imag} */,
  {32'hbf8b04fe, 32'h3fe2ebfc} /* (11, 6, 12) {real, imag} */,
  {32'hbf4a580e, 32'h3fe90511} /* (11, 6, 11) {real, imag} */,
  {32'h3fdf02db, 32'h3f2c2b3d} /* (11, 6, 10) {real, imag} */,
  {32'h3f29497e, 32'h3fcd9396} /* (11, 6, 9) {real, imag} */,
  {32'hbef26ea8, 32'h3faddffe} /* (11, 6, 8) {real, imag} */,
  {32'hbe700488, 32'h4010c005} /* (11, 6, 7) {real, imag} */,
  {32'hbf9e9ace, 32'h3f45c210} /* (11, 6, 6) {real, imag} */,
  {32'hbfbfa1b8, 32'hbf5a5490} /* (11, 6, 5) {real, imag} */,
  {32'hbf4596ca, 32'h3f83c07e} /* (11, 6, 4) {real, imag} */,
  {32'hc014ed20, 32'h3fffc8ba} /* (11, 6, 3) {real, imag} */,
  {32'hc02cda24, 32'hbee1ae44} /* (11, 6, 2) {real, imag} */,
  {32'h3d6c6660, 32'hc018fb3c} /* (11, 6, 1) {real, imag} */,
  {32'h3e2642f8, 32'hc02469ee} /* (11, 6, 0) {real, imag} */,
  {32'hbe789478, 32'h3fdfface} /* (11, 5, 15) {real, imag} */,
  {32'h3f262dc0, 32'h40216010} /* (11, 5, 14) {real, imag} */,
  {32'h3fa5c9ea, 32'hc0075620} /* (11, 5, 13) {real, imag} */,
  {32'h3f21b588, 32'hc016dc72} /* (11, 5, 12) {real, imag} */,
  {32'h3fa0abce, 32'hbfd987c4} /* (11, 5, 11) {real, imag} */,
  {32'h4020470c, 32'h3daca700} /* (11, 5, 10) {real, imag} */,
  {32'h3fa226d0, 32'h40853fc2} /* (11, 5, 9) {real, imag} */,
  {32'hbfe1c284, 32'h407291ed} /* (11, 5, 8) {real, imag} */,
  {32'hbef68240, 32'h406f7695} /* (11, 5, 7) {real, imag} */,
  {32'hbf822620, 32'h4012ed76} /* (11, 5, 6) {real, imag} */,
  {32'h3e862c94, 32'hbff047ae} /* (11, 5, 5) {real, imag} */,
  {32'h401cf9de, 32'hc0668990} /* (11, 5, 4) {real, imag} */,
  {32'h3ff3b652, 32'hbf4f0b78} /* (11, 5, 3) {real, imag} */,
  {32'h3f3b04b3, 32'h3f87183c} /* (11, 5, 2) {real, imag} */,
  {32'h3faf7676, 32'hbeb28e14} /* (11, 5, 1) {real, imag} */,
  {32'hbeac3c42, 32'h3f657380} /* (11, 5, 0) {real, imag} */,
  {32'h3fa06ba8, 32'hc0427a2e} /* (11, 4, 15) {real, imag} */,
  {32'h3f7e0992, 32'hc05531d0} /* (11, 4, 14) {real, imag} */,
  {32'hbf47d7ba, 32'hbf92df93} /* (11, 4, 13) {real, imag} */,
  {32'h4027136a, 32'hc026a70d} /* (11, 4, 12) {real, imag} */,
  {32'h3f804f5d, 32'hbfa29067} /* (11, 4, 11) {real, imag} */,
  {32'hbf8a09d2, 32'h3e418968} /* (11, 4, 10) {real, imag} */,
  {32'h3f83dc78, 32'h40213b12} /* (11, 4, 9) {real, imag} */,
  {32'h403d7564, 32'h3f939702} /* (11, 4, 8) {real, imag} */,
  {32'hc0086f7f, 32'hbfabded0} /* (11, 4, 7) {real, imag} */,
  {32'h405c69c6, 32'hc09c5a0d} /* (11, 4, 6) {real, imag} */,
  {32'h4044bdc9, 32'hbffd1731} /* (11, 4, 5) {real, imag} */,
  {32'hbf662ee5, 32'h3d595478} /* (11, 4, 4) {real, imag} */,
  {32'h3f4c6fed, 32'h3f965ed9} /* (11, 4, 3) {real, imag} */,
  {32'hbf93185c, 32'h4048958a} /* (11, 4, 2) {real, imag} */,
  {32'h3f65a61c, 32'h405abdf0} /* (11, 4, 1) {real, imag} */,
  {32'h3f3260ba, 32'hbee56d98} /* (11, 4, 0) {real, imag} */,
  {32'h3f77664a, 32'h3f26f084} /* (11, 3, 15) {real, imag} */,
  {32'hc03705ab, 32'h3e8f1b2a} /* (11, 3, 14) {real, imag} */,
  {32'hc0330ab4, 32'hbfee4091} /* (11, 3, 13) {real, imag} */,
  {32'hbfca1bf6, 32'hc01d509c} /* (11, 3, 12) {real, imag} */,
  {32'hc02d6792, 32'hc04dc9de} /* (11, 3, 11) {real, imag} */,
  {32'h404e3a60, 32'hc0939e20} /* (11, 3, 10) {real, imag} */,
  {32'h40221577, 32'h3e439f28} /* (11, 3, 9) {real, imag} */,
  {32'hc045f1b8, 32'h40b19c9a} /* (11, 3, 8) {real, imag} */,
  {32'hbfeb6742, 32'h4048e5f4} /* (11, 3, 7) {real, imag} */,
  {32'hbfd115ca, 32'h3fad91aa} /* (11, 3, 6) {real, imag} */,
  {32'hbf24d416, 32'h40076be6} /* (11, 3, 5) {real, imag} */,
  {32'h40089b01, 32'h3e85d660} /* (11, 3, 4) {real, imag} */,
  {32'h3f98255e, 32'hc059aa60} /* (11, 3, 3) {real, imag} */,
  {32'hbf53acec, 32'hc07ffd75} /* (11, 3, 2) {real, imag} */,
  {32'hbe30bb90, 32'h3f992fe0} /* (11, 3, 1) {real, imag} */,
  {32'h3ff9c060, 32'h3fe8f4c3} /* (11, 3, 0) {real, imag} */,
  {32'h3e874c68, 32'h40991a5d} /* (11, 2, 15) {real, imag} */,
  {32'h40849c74, 32'h3e5d6a90} /* (11, 2, 14) {real, imag} */,
  {32'h4092e323, 32'hbfec20bb} /* (11, 2, 13) {real, imag} */,
  {32'h408965ea, 32'h3ef52427} /* (11, 2, 12) {real, imag} */,
  {32'hc0aad736, 32'hbe657918} /* (11, 2, 11) {real, imag} */,
  {32'hc01d4285, 32'h4047ff72} /* (11, 2, 10) {real, imag} */,
  {32'hc0145afe, 32'hc0cc5fc4} /* (11, 2, 9) {real, imag} */,
  {32'hbf18bb28, 32'hc0b7f65c} /* (11, 2, 8) {real, imag} */,
  {32'h3f6be5d4, 32'hc06dd27f} /* (11, 2, 7) {real, imag} */,
  {32'hbfddd363, 32'h3f8c1c22} /* (11, 2, 6) {real, imag} */,
  {32'h3f8c993c, 32'h40a51194} /* (11, 2, 5) {real, imag} */,
  {32'hc003b42a, 32'hc0a56c98} /* (11, 2, 4) {real, imag} */,
  {32'h3f4aa968, 32'hc0d68bd0} /* (11, 2, 3) {real, imag} */,
  {32'h3edc0790, 32'h3f5f6188} /* (11, 2, 2) {real, imag} */,
  {32'hc0758cba, 32'h3f20bb54} /* (11, 2, 1) {real, imag} */,
  {32'h3e1f0248, 32'hbf68bc20} /* (11, 2, 0) {real, imag} */,
  {32'h40523aa4, 32'h40790e4e} /* (11, 1, 15) {real, imag} */,
  {32'h403ec375, 32'h4050c411} /* (11, 1, 14) {real, imag} */,
  {32'h3f7691c8, 32'hbfc6fa45} /* (11, 1, 13) {real, imag} */,
  {32'hbe467cb8, 32'h4024358d} /* (11, 1, 12) {real, imag} */,
  {32'h40b0a71a, 32'h401b0d2c} /* (11, 1, 11) {real, imag} */,
  {32'hbfa169fb, 32'hc02b9220} /* (11, 1, 10) {real, imag} */,
  {32'hc082e0bb, 32'hbfb820e0} /* (11, 1, 9) {real, imag} */,
  {32'h405affba, 32'hbfd2b4ed} /* (11, 1, 8) {real, imag} */,
  {32'h3fb73058, 32'hbe645fb8} /* (11, 1, 7) {real, imag} */,
  {32'hc0a4e56b, 32'h40ca6844} /* (11, 1, 6) {real, imag} */,
  {32'hbfd807d8, 32'h3d866b10} /* (11, 1, 5) {real, imag} */,
  {32'hbf06d226, 32'hc0720f52} /* (11, 1, 4) {real, imag} */,
  {32'hbfd3b9c2, 32'h3d89f360} /* (11, 1, 3) {real, imag} */,
  {32'h3f6b82ca, 32'hbf84ee26} /* (11, 1, 2) {real, imag} */,
  {32'h402e257a, 32'hbd223b60} /* (11, 1, 1) {real, imag} */,
  {32'h40b9a2e4, 32'h3ffb1ecc} /* (11, 1, 0) {real, imag} */,
  {32'hbf88b629, 32'hbf051832} /* (11, 0, 15) {real, imag} */,
  {32'hc047d1f5, 32'h3e4adc68} /* (11, 0, 14) {real, imag} */,
  {32'h407e3a6a, 32'h40a2fe00} /* (11, 0, 13) {real, imag} */,
  {32'h40dea0a0, 32'h40bc220f} /* (11, 0, 12) {real, imag} */,
  {32'h3f4b5162, 32'h4050bcda} /* (11, 0, 11) {real, imag} */,
  {32'hc081909a, 32'h406af976} /* (11, 0, 10) {real, imag} */,
  {32'h404a8ebd, 32'h40569bc0} /* (11, 0, 9) {real, imag} */,
  {32'h4065b244, 32'h4077219a} /* (11, 0, 8) {real, imag} */,
  {32'hbff308f3, 32'h40514d46} /* (11, 0, 7) {real, imag} */,
  {32'h4030def6, 32'hbf0e354f} /* (11, 0, 6) {real, imag} */,
  {32'h40b455c8, 32'h403cd912} /* (11, 0, 5) {real, imag} */,
  {32'h4037cade, 32'h400e6324} /* (11, 0, 4) {real, imag} */,
  {32'h40942433, 32'h4024531c} /* (11, 0, 3) {real, imag} */,
  {32'h40b1eb58, 32'hbfd82a54} /* (11, 0, 2) {real, imag} */,
  {32'h3f3f12d5, 32'hbeb1d448} /* (11, 0, 1) {real, imag} */,
  {32'hbf94f5f6, 32'h40c36efb} /* (11, 0, 0) {real, imag} */,
  {32'hbf844675, 32'h3fe3a66f} /* (10, 15, 15) {real, imag} */,
  {32'hbf0817c6, 32'h40d294fa} /* (10, 15, 14) {real, imag} */,
  {32'h40a79e64, 32'h40c97118} /* (10, 15, 13) {real, imag} */,
  {32'h406af226, 32'h3f2c3ab4} /* (10, 15, 12) {real, imag} */,
  {32'hbe80fd8c, 32'hc08d4990} /* (10, 15, 11) {real, imag} */,
  {32'h3ece8988, 32'h3ec560b6} /* (10, 15, 10) {real, imag} */,
  {32'h402f54ad, 32'h3ff06d46} /* (10, 15, 9) {real, imag} */,
  {32'h400636da, 32'h40810710} /* (10, 15, 8) {real, imag} */,
  {32'hbf7e1bba, 32'hbf2881e8} /* (10, 15, 7) {real, imag} */,
  {32'hbe0a6f58, 32'hc000db76} /* (10, 15, 6) {real, imag} */,
  {32'h40eae60c, 32'h3f9a7a4d} /* (10, 15, 5) {real, imag} */,
  {32'h40cea718, 32'hbf9feb22} /* (10, 15, 4) {real, imag} */,
  {32'h4087885e, 32'hbe89acc6} /* (10, 15, 3) {real, imag} */,
  {32'h400898e4, 32'h4041d103} /* (10, 15, 2) {real, imag} */,
  {32'h3e3e12d2, 32'hc0550cf7} /* (10, 15, 1) {real, imag} */,
  {32'h3f486384, 32'hc0b55152} /* (10, 15, 0) {real, imag} */,
  {32'hc0131ac1, 32'hc02befbb} /* (10, 14, 15) {real, imag} */,
  {32'hbf37fa38, 32'hc0b6b888} /* (10, 14, 14) {real, imag} */,
  {32'h40565e8c, 32'hc0a2aca6} /* (10, 14, 13) {real, imag} */,
  {32'h406e693b, 32'hc09dd05b} /* (10, 14, 12) {real, imag} */,
  {32'h3fd8bbc2, 32'hc09caa21} /* (10, 14, 11) {real, imag} */,
  {32'h403b9b5a, 32'hc0cab301} /* (10, 14, 10) {real, imag} */,
  {32'h405fb9ce, 32'hbef6785b} /* (10, 14, 9) {real, imag} */,
  {32'hbf1f3dae, 32'h3fc992ec} /* (10, 14, 8) {real, imag} */,
  {32'hbf128fcd, 32'hbf088bd2} /* (10, 14, 7) {real, imag} */,
  {32'h40c72056, 32'h4085c70d} /* (10, 14, 6) {real, imag} */,
  {32'h40ffd4aa, 32'h40c25867} /* (10, 14, 5) {real, imag} */,
  {32'h40282f9c, 32'h4039c91d} /* (10, 14, 4) {real, imag} */,
  {32'hbf94da12, 32'h3f5412c5} /* (10, 14, 3) {real, imag} */,
  {32'h3f1f21ce, 32'hbed665ec} /* (10, 14, 2) {real, imag} */,
  {32'h3f06dd17, 32'hc026d153} /* (10, 14, 1) {real, imag} */,
  {32'hbd264db8, 32'hc0395a40} /* (10, 14, 0) {real, imag} */,
  {32'hbf01f94a, 32'h3f4336b2} /* (10, 13, 15) {real, imag} */,
  {32'hbfc0f2cc, 32'h4037a6b3} /* (10, 13, 14) {real, imag} */,
  {32'hbe2e51e0, 32'h40a265fe} /* (10, 13, 13) {real, imag} */,
  {32'h3ffb75ce, 32'h403e031a} /* (10, 13, 12) {real, imag} */,
  {32'hbf851e23, 32'h3f58f50a} /* (10, 13, 11) {real, imag} */,
  {32'hc02e5870, 32'hbf85b8d8} /* (10, 13, 10) {real, imag} */,
  {32'h3eb2acb6, 32'hbf24e147} /* (10, 13, 9) {real, imag} */,
  {32'h3faa74f2, 32'h3e7efca8} /* (10, 13, 8) {real, imag} */,
  {32'h400ca872, 32'h3f420d78} /* (10, 13, 7) {real, imag} */,
  {32'h3f75d247, 32'h3f870327} /* (10, 13, 6) {real, imag} */,
  {32'hbb6b6600, 32'hbfa80404} /* (10, 13, 5) {real, imag} */,
  {32'h3f3bf784, 32'h3e6e60f0} /* (10, 13, 4) {real, imag} */,
  {32'h3d1d03a4, 32'h404268b9} /* (10, 13, 3) {real, imag} */,
  {32'hbf9231dc, 32'h40741208} /* (10, 13, 2) {real, imag} */,
  {32'hbf15aaf0, 32'h401ac7f8} /* (10, 13, 1) {real, imag} */,
  {32'hbb941100, 32'hbfa47e00} /* (10, 13, 0) {real, imag} */,
  {32'h3fa192eb, 32'hbf38d151} /* (10, 12, 15) {real, imag} */,
  {32'h402c9c3e, 32'h3fb8224f} /* (10, 12, 14) {real, imag} */,
  {32'h40025ff9, 32'h402090c0} /* (10, 12, 13) {real, imag} */,
  {32'h3e0aa746, 32'h3feea880} /* (10, 12, 12) {real, imag} */,
  {32'hbf81c1b2, 32'hc0682378} /* (10, 12, 11) {real, imag} */,
  {32'hbfa88216, 32'hbffd68a4} /* (10, 12, 10) {real, imag} */,
  {32'hc024fcf4, 32'hc0116d06} /* (10, 12, 9) {real, imag} */,
  {32'hc0211907, 32'hc0378f80} /* (10, 12, 8) {real, imag} */,
  {32'hbfdf75c4, 32'hbff33d52} /* (10, 12, 7) {real, imag} */,
  {32'hbfa57a0a, 32'h3f81972d} /* (10, 12, 6) {real, imag} */,
  {32'hc026de41, 32'h40549ba2} /* (10, 12, 5) {real, imag} */,
  {32'hc02c02be, 32'h3f710aa8} /* (10, 12, 4) {real, imag} */,
  {32'hbfd2d634, 32'hc03e6403} /* (10, 12, 3) {real, imag} */,
  {32'h3f29a9ef, 32'hbf317379} /* (10, 12, 2) {real, imag} */,
  {32'h3f65ffae, 32'hbfe97053} /* (10, 12, 1) {real, imag} */,
  {32'hbee34280, 32'hbe49a1a4} /* (10, 12, 0) {real, imag} */,
  {32'h3fa5a416, 32'h3ec82e12} /* (10, 11, 15) {real, imag} */,
  {32'hbf77803a, 32'h3faf7ec2} /* (10, 11, 14) {real, imag} */,
  {32'hbecb3eb8, 32'hbfea0b3c} /* (10, 11, 13) {real, imag} */,
  {32'h3ffbf0fa, 32'hbfe760bb} /* (10, 11, 12) {real, imag} */,
  {32'h3fc46a6a, 32'hbfc64eeb} /* (10, 11, 11) {real, imag} */,
  {32'h3e8da59a, 32'hbfd2b27b} /* (10, 11, 10) {real, imag} */,
  {32'hc00b8900, 32'h40248dd2} /* (10, 11, 9) {real, imag} */,
  {32'hbffb90ce, 32'h3fcffd0f} /* (10, 11, 8) {real, imag} */,
  {32'h3f2d6106, 32'hbef7d882} /* (10, 11, 7) {real, imag} */,
  {32'h3fd64de6, 32'hc062334a} /* (10, 11, 6) {real, imag} */,
  {32'hbf7b2672, 32'hc00d6e77} /* (10, 11, 5) {real, imag} */,
  {32'hc0318e01, 32'hc0013846} /* (10, 11, 4) {real, imag} */,
  {32'h3f8512f1, 32'hc021ecfc} /* (10, 11, 3) {real, imag} */,
  {32'h4027dd6b, 32'hbfcc211c} /* (10, 11, 2) {real, imag} */,
  {32'h4014c91f, 32'h3df89ea0} /* (10, 11, 1) {real, imag} */,
  {32'h3f0f5f4f, 32'h3d99bc18} /* (10, 11, 0) {real, imag} */,
  {32'hbfc7143a, 32'h4003d72c} /* (10, 10, 15) {real, imag} */,
  {32'hbf97e032, 32'h403b914f} /* (10, 10, 14) {real, imag} */,
  {32'hbf2b74e1, 32'h3fb70252} /* (10, 10, 13) {real, imag} */,
  {32'hbf9d03d2, 32'hbe181998} /* (10, 10, 12) {real, imag} */,
  {32'hbf25bbf4, 32'hbf151252} /* (10, 10, 11) {real, imag} */,
  {32'h3e8f0104, 32'h3e2fce78} /* (10, 10, 10) {real, imag} */,
  {32'hbe9b5026, 32'h3d81e5e8} /* (10, 10, 9) {real, imag} */,
  {32'h3d9eca24, 32'hbf355723} /* (10, 10, 8) {real, imag} */,
  {32'hbf56ecca, 32'hbeee03d4} /* (10, 10, 7) {real, imag} */,
  {32'hc0166320, 32'h3ee7fd34} /* (10, 10, 6) {real, imag} */,
  {32'hbfa12597, 32'h3f689dde} /* (10, 10, 5) {real, imag} */,
  {32'hbf8131e6, 32'hbfd9e561} /* (10, 10, 4) {real, imag} */,
  {32'hbee3f13c, 32'hbfa4a15a} /* (10, 10, 3) {real, imag} */,
  {32'hbee222ef, 32'h3ec953e2} /* (10, 10, 2) {real, imag} */,
  {32'hbf586c87, 32'h3f162d49} /* (10, 10, 1) {real, imag} */,
  {32'hbda5147c, 32'h3eaafd0a} /* (10, 10, 0) {real, imag} */,
  {32'h3e8eef96, 32'hbf6492d8} /* (10, 9, 15) {real, imag} */,
  {32'h3f995a75, 32'hbfd7ff61} /* (10, 9, 14) {real, imag} */,
  {32'h3f2ba0de, 32'hbd9216a0} /* (10, 9, 13) {real, imag} */,
  {32'hbeae2eb4, 32'h3f8085ba} /* (10, 9, 12) {real, imag} */,
  {32'h3f53ebd2, 32'h3edef67c} /* (10, 9, 11) {real, imag} */,
  {32'h3fcd1bdf, 32'h3ebadd8e} /* (10, 9, 10) {real, imag} */,
  {32'hbd8e9ba8, 32'hbf70be04} /* (10, 9, 9) {real, imag} */,
  {32'h3e7986d0, 32'hbf776dd3} /* (10, 9, 8) {real, imag} */,
  {32'h3f366be6, 32'h3ea6bd60} /* (10, 9, 7) {real, imag} */,
  {32'h3f6cdf56, 32'h3f9ad172} /* (10, 9, 6) {real, imag} */,
  {32'h3eb4bb6c, 32'h3efcea7f} /* (10, 9, 5) {real, imag} */,
  {32'h3feb1127, 32'h3e439f58} /* (10, 9, 4) {real, imag} */,
  {32'h3e83b3e8, 32'hbf011add} /* (10, 9, 3) {real, imag} */,
  {32'hbf6475e1, 32'h3f59ee04} /* (10, 9, 2) {real, imag} */,
  {32'hbf350d0e, 32'h3fa30698} /* (10, 9, 1) {real, imag} */,
  {32'hbe1d8e57, 32'h3f691191} /* (10, 9, 0) {real, imag} */,
  {32'h3d675080, 32'hbf4fb580} /* (10, 8, 15) {real, imag} */,
  {32'h3ee55084, 32'hbefa9b6c} /* (10, 8, 14) {real, imag} */,
  {32'h3f80c102, 32'h3f4ebd70} /* (10, 8, 13) {real, imag} */,
  {32'h3ef0946e, 32'h3f196eaa} /* (10, 8, 12) {real, imag} */,
  {32'h3f058902, 32'h3f938d00} /* (10, 8, 11) {real, imag} */,
  {32'hbe5a9488, 32'h3faec572} /* (10, 8, 10) {real, imag} */,
  {32'hbf916d57, 32'hbf526de9} /* (10, 8, 9) {real, imag} */,
  {32'h3db55ea0, 32'hbf90ac16} /* (10, 8, 8) {real, imag} */,
  {32'h3f7a5c36, 32'hbf17f72a} /* (10, 8, 7) {real, imag} */,
  {32'h3dcc7200, 32'hbf3b7140} /* (10, 8, 6) {real, imag} */,
  {32'hbbd4f100, 32'hbf89b55a} /* (10, 8, 5) {real, imag} */,
  {32'hbecd0b6c, 32'hbe23fac8} /* (10, 8, 4) {real, imag} */,
  {32'h3e582ea0, 32'hbee941e0} /* (10, 8, 3) {real, imag} */,
  {32'h3eaf8df8, 32'hbf365888} /* (10, 8, 2) {real, imag} */,
  {32'hbdf98084, 32'hbf0a89fc} /* (10, 8, 1) {real, imag} */,
  {32'h3ee9c314, 32'hbf046df4} /* (10, 8, 0) {real, imag} */,
  {32'h3f179c2b, 32'h3e84c5ef} /* (10, 7, 15) {real, imag} */,
  {32'h3ef17fe3, 32'h3d9fa2d0} /* (10, 7, 14) {real, imag} */,
  {32'hbec079ec, 32'hbf9d65ee} /* (10, 7, 13) {real, imag} */,
  {32'h3e286e68, 32'hbf8419e0} /* (10, 7, 12) {real, imag} */,
  {32'h3f8d73c5, 32'h3e9ffbec} /* (10, 7, 11) {real, imag} */,
  {32'h3f62e3e6, 32'h3fd2a39e} /* (10, 7, 10) {real, imag} */,
  {32'h3f84ac32, 32'h3f8a3282} /* (10, 7, 9) {real, imag} */,
  {32'h3f80f110, 32'hbde0c6d8} /* (10, 7, 8) {real, imag} */,
  {32'hbe19eb1c, 32'hbe9f2510} /* (10, 7, 7) {real, imag} */,
  {32'hbef49353, 32'hbda1e4b8} /* (10, 7, 6) {real, imag} */,
  {32'hbf1bac32, 32'hbf568ed6} /* (10, 7, 5) {real, imag} */,
  {32'h3f7de196, 32'hbf318420} /* (10, 7, 4) {real, imag} */,
  {32'h3ff313aa, 32'hbfe390b2} /* (10, 7, 3) {real, imag} */,
  {32'h3d0826f0, 32'hbf817ae1} /* (10, 7, 2) {real, imag} */,
  {32'hbf774ff6, 32'h3e65869c} /* (10, 7, 1) {real, imag} */,
  {32'hbe93abfc, 32'h3b912780} /* (10, 7, 0) {real, imag} */,
  {32'hbf82f66a, 32'hbea401f4} /* (10, 6, 15) {real, imag} */,
  {32'hbfd3e86a, 32'h3eff7408} /* (10, 6, 14) {real, imag} */,
  {32'h3f470da3, 32'hbcacbe80} /* (10, 6, 13) {real, imag} */,
  {32'h3fdbe5d6, 32'hc0117f3a} /* (10, 6, 12) {real, imag} */,
  {32'h401fae78, 32'hbfcf6277} /* (10, 6, 11) {real, imag} */,
  {32'hbffed3f7, 32'hbf2d31ea} /* (10, 6, 10) {real, imag} */,
  {32'hbff15324, 32'h3fcce56c} /* (10, 6, 9) {real, imag} */,
  {32'h3ef30db1, 32'hbec7b0ee} /* (10, 6, 8) {real, imag} */,
  {32'hbed63910, 32'hbcf2d0a0} /* (10, 6, 7) {real, imag} */,
  {32'hbf8c793b, 32'h3f91f559} /* (10, 6, 6) {real, imag} */,
  {32'h3f8f8b03, 32'h3fe246c1} /* (10, 6, 5) {real, imag} */,
  {32'h3f796e9c, 32'h3fea8fdd} /* (10, 6, 4) {real, imag} */,
  {32'h3e26fcc0, 32'hbf39533f} /* (10, 6, 3) {real, imag} */,
  {32'h3ee05059, 32'h3de43598} /* (10, 6, 2) {real, imag} */,
  {32'hbf6d3e99, 32'h3fb2152c} /* (10, 6, 1) {real, imag} */,
  {32'hbf448f38, 32'h3e24ccb4} /* (10, 6, 0) {real, imag} */,
  {32'hbf9ba958, 32'hbf8379de} /* (10, 5, 15) {real, imag} */,
  {32'h3d92c050, 32'hbe6d8b9c} /* (10, 5, 14) {real, imag} */,
  {32'h401c983d, 32'h3e7ec800} /* (10, 5, 13) {real, imag} */,
  {32'h3f9bb01c, 32'h3df791b0} /* (10, 5, 12) {real, imag} */,
  {32'hc04078fb, 32'h3dfa5b30} /* (10, 5, 11) {real, imag} */,
  {32'hbf5a492f, 32'hc031de44} /* (10, 5, 10) {real, imag} */,
  {32'h3f546f4e, 32'hbfc4e3bb} /* (10, 5, 9) {real, imag} */,
  {32'h3f3542f4, 32'hbefafa7c} /* (10, 5, 8) {real, imag} */,
  {32'h3fb6fe0b, 32'h3f951bc6} /* (10, 5, 7) {real, imag} */,
  {32'h3e098bcc, 32'hbffa3e7b} /* (10, 5, 6) {real, imag} */,
  {32'h400c93b2, 32'hbf3432ad} /* (10, 5, 5) {real, imag} */,
  {32'h3fb4878a, 32'h3f59b677} /* (10, 5, 4) {real, imag} */,
  {32'h3f9eece5, 32'hbedc26dc} /* (10, 5, 3) {real, imag} */,
  {32'h40052279, 32'h3f03a1ab} /* (10, 5, 2) {real, imag} */,
  {32'h3fb4dcba, 32'hbe849d20} /* (10, 5, 1) {real, imag} */,
  {32'hbf911ad2, 32'hbf804d2e} /* (10, 5, 0) {real, imag} */,
  {32'hc0158808, 32'hbf34eb6b} /* (10, 4, 15) {real, imag} */,
  {32'h3f8d0ce2, 32'hc046b992} /* (10, 4, 14) {real, imag} */,
  {32'h406357fd, 32'hc029d438} /* (10, 4, 13) {real, imag} */,
  {32'h3f1c2a98, 32'hbcfe3a20} /* (10, 4, 12) {real, imag} */,
  {32'hbfcb9238, 32'hbe9630cc} /* (10, 4, 11) {real, imag} */,
  {32'h3f46e9eb, 32'hc0555f88} /* (10, 4, 10) {real, imag} */,
  {32'h3f6d2aa6, 32'hc0d792c1} /* (10, 4, 9) {real, imag} */,
  {32'h409c51f2, 32'hbf89ad08} /* (10, 4, 8) {real, imag} */,
  {32'h4094b581, 32'hbfb1c38c} /* (10, 4, 7) {real, imag} */,
  {32'hbdf24998, 32'hc000c920} /* (10, 4, 6) {real, imag} */,
  {32'hbfc8ff72, 32'h3fa1b93f} /* (10, 4, 5) {real, imag} */,
  {32'h3fd8a530, 32'h3fae2138} /* (10, 4, 4) {real, imag} */,
  {32'h3d50fd90, 32'h3e5008b0} /* (10, 4, 3) {real, imag} */,
  {32'hbf1b82c3, 32'hbf2ce2cf} /* (10, 4, 2) {real, imag} */,
  {32'hbf9df56f, 32'h3f84501b} /* (10, 4, 1) {real, imag} */,
  {32'hbfe85f40, 32'h3fa7e216} /* (10, 4, 0) {real, imag} */,
  {32'hc01fecf8, 32'h40185a3a} /* (10, 3, 15) {real, imag} */,
  {32'hbf9a9c74, 32'h408abc55} /* (10, 3, 14) {real, imag} */,
  {32'h3fc9f8e5, 32'h405b9654} /* (10, 3, 13) {real, imag} */,
  {32'hbfc1975c, 32'hbf68c676} /* (10, 3, 12) {real, imag} */,
  {32'hc031c844, 32'hbff91a45} /* (10, 3, 11) {real, imag} */,
  {32'h3e5ea308, 32'hbfa6fc00} /* (10, 3, 10) {real, imag} */,
  {32'hbf87e5b2, 32'hbf5c51e5} /* (10, 3, 9) {real, imag} */,
  {32'hc07640cb, 32'h407fc688} /* (10, 3, 8) {real, imag} */,
  {32'hc0838eeb, 32'h40220182} /* (10, 3, 7) {real, imag} */,
  {32'hc01a6174, 32'hbf5987a2} /* (10, 3, 6) {real, imag} */,
  {32'hc06db010, 32'h3f3be70d} /* (10, 3, 5) {real, imag} */,
  {32'hc068c8ad, 32'h40413be7} /* (10, 3, 4) {real, imag} */,
  {32'hbe99d37c, 32'h404cdcc7} /* (10, 3, 3) {real, imag} */,
  {32'h3f9c86d4, 32'hbf382840} /* (10, 3, 2) {real, imag} */,
  {32'h4089c815, 32'h3f1e180a} /* (10, 3, 1) {real, imag} */,
  {32'h402ec1ac, 32'h3fdea1a4} /* (10, 3, 0) {real, imag} */,
  {32'h3f82baca, 32'h3fe84ee2} /* (10, 2, 15) {real, imag} */,
  {32'h403ca726, 32'h3ec30fc8} /* (10, 2, 14) {real, imag} */,
  {32'h3eb08f04, 32'hbfe7803a} /* (10, 2, 13) {real, imag} */,
  {32'h40260565, 32'h3e9fd630} /* (10, 2, 12) {real, imag} */,
  {32'hbfeda528, 32'h3f446248} /* (10, 2, 11) {real, imag} */,
  {32'hc0273c10, 32'h3fe9067c} /* (10, 2, 10) {real, imag} */,
  {32'hbf2d85f6, 32'h3e498002} /* (10, 2, 9) {real, imag} */,
  {32'h3f855a19, 32'h40166b60} /* (10, 2, 8) {real, imag} */,
  {32'hc0133575, 32'hbf19c8ba} /* (10, 2, 7) {real, imag} */,
  {32'h3fab64f6, 32'hbf9a4ff9} /* (10, 2, 6) {real, imag} */,
  {32'h40631aec, 32'hbe0d9c20} /* (10, 2, 5) {real, imag} */,
  {32'h4058bbd2, 32'hc0734bc3} /* (10, 2, 4) {real, imag} */,
  {32'hc01992d9, 32'hc0297e8d} /* (10, 2, 3) {real, imag} */,
  {32'hc013976c, 32'hc03477dc} /* (10, 2, 2) {real, imag} */,
  {32'h3f96d78a, 32'hc0259b27} /* (10, 2, 1) {real, imag} */,
  {32'h3ed3b273, 32'h3e9ca41c} /* (10, 2, 0) {real, imag} */,
  {32'hc003b74c, 32'hc008b047} /* (10, 1, 15) {real, imag} */,
  {32'hbee40baa, 32'hbcfef680} /* (10, 1, 14) {real, imag} */,
  {32'hbde4fda0, 32'h40423440} /* (10, 1, 13) {real, imag} */,
  {32'hc02ebff6, 32'h40248996} /* (10, 1, 12) {real, imag} */,
  {32'hc05a1b96, 32'h403612fa} /* (10, 1, 11) {real, imag} */,
  {32'hc0b91eea, 32'h3f98a174} /* (10, 1, 10) {real, imag} */,
  {32'hbfb22d1a, 32'hbf3f1fec} /* (10, 1, 9) {real, imag} */,
  {32'hc037defa, 32'hc07d65a5} /* (10, 1, 8) {real, imag} */,
  {32'h3e09e4d6, 32'hc0bb418a} /* (10, 1, 7) {real, imag} */,
  {32'hbf9d603b, 32'hc0a479a5} /* (10, 1, 6) {real, imag} */,
  {32'hc0910808, 32'hc0230114} /* (10, 1, 5) {real, imag} */,
  {32'hc0c69464, 32'h400f0439} /* (10, 1, 4) {real, imag} */,
  {32'hc04261dc, 32'hbdc33ff8} /* (10, 1, 3) {real, imag} */,
  {32'h3ffc26a5, 32'hbe98abd8} /* (10, 1, 2) {real, imag} */,
  {32'hbf4498a8, 32'hc09703e4} /* (10, 1, 1) {real, imag} */,
  {32'h3f16f80c, 32'hc04a54bc} /* (10, 1, 0) {real, imag} */,
  {32'h4010587e, 32'hbed53338} /* (10, 0, 15) {real, imag} */,
  {32'h3fe5a165, 32'hc05689dc} /* (10, 0, 14) {real, imag} */,
  {32'hbfabb546, 32'hc0bffb68} /* (10, 0, 13) {real, imag} */,
  {32'hbfdc17bc, 32'hbf397662} /* (10, 0, 12) {real, imag} */,
  {32'h4003b11c, 32'h4022b245} /* (10, 0, 11) {real, imag} */,
  {32'h3fba2a88, 32'h3fbe872a} /* (10, 0, 10) {real, imag} */,
  {32'h3eeea20c, 32'hbe57c73c} /* (10, 0, 9) {real, imag} */,
  {32'h3f8439de, 32'hbf9bd93a} /* (10, 0, 8) {real, imag} */,
  {32'hbfbfb753, 32'hc05d12fe} /* (10, 0, 7) {real, imag} */,
  {32'hc086a728, 32'hc07a2bb6} /* (10, 0, 6) {real, imag} */,
  {32'hc001a514, 32'hc09a3002} /* (10, 0, 5) {real, imag} */,
  {32'hbd8e5fce, 32'h3eacc868} /* (10, 0, 4) {real, imag} */,
  {32'h4024aaca, 32'h4050a070} /* (10, 0, 3) {real, imag} */,
  {32'h402ab9b1, 32'h40239db8} /* (10, 0, 2) {real, imag} */,
  {32'h3f090148, 32'h40869a8e} /* (10, 0, 1) {real, imag} */,
  {32'hbfbe46b4, 32'h4030c9e7} /* (10, 0, 0) {real, imag} */,
  {32'h4024cb65, 32'h404e41a6} /* (9, 15, 15) {real, imag} */,
  {32'h3fcdc566, 32'h3fda6c6f} /* (9, 15, 14) {real, imag} */,
  {32'h3f6bae73, 32'h3f1845c5} /* (9, 15, 13) {real, imag} */,
  {32'h4011a9c2, 32'h40652e3a} /* (9, 15, 12) {real, imag} */,
  {32'hbf7d8ac4, 32'h406e1e8a} /* (9, 15, 11) {real, imag} */,
  {32'hc00b8778, 32'h3f3e3e28} /* (9, 15, 10) {real, imag} */,
  {32'hbf6f5db2, 32'h401b9c62} /* (9, 15, 9) {real, imag} */,
  {32'hbeb240f8, 32'h3f6c0a2c} /* (9, 15, 8) {real, imag} */,
  {32'h3e8ddf3c, 32'hbfa7aeb0} /* (9, 15, 7) {real, imag} */,
  {32'hbfa3b2a6, 32'h3fd81d77} /* (9, 15, 6) {real, imag} */,
  {32'hc09b7350, 32'hbf065a5e} /* (9, 15, 5) {real, imag} */,
  {32'hc0029a93, 32'hc035f223} /* (9, 15, 4) {real, imag} */,
  {32'h400b2e22, 32'hbdd9c610} /* (9, 15, 3) {real, imag} */,
  {32'h4037780b, 32'h3e66e150} /* (9, 15, 2) {real, imag} */,
  {32'hbf7f0b2d, 32'hbeafafbc} /* (9, 15, 1) {real, imag} */,
  {32'hbf1444c0, 32'hbfcdcd9b} /* (9, 15, 0) {real, imag} */,
  {32'hbf5eefe0, 32'hc013f678} /* (9, 14, 15) {real, imag} */,
  {32'h3e7e2428, 32'hc012d856} /* (9, 14, 14) {real, imag} */,
  {32'hbf71a474, 32'h3f79c6e4} /* (9, 14, 13) {real, imag} */,
  {32'hbfe25038, 32'h3f5ac1d6} /* (9, 14, 12) {real, imag} */,
  {32'hbf0943ea, 32'h4021989c} /* (9, 14, 11) {real, imag} */,
  {32'hbfc8c712, 32'h3ffaebce} /* (9, 14, 10) {real, imag} */,
  {32'hc030a9f0, 32'hc015b16b} /* (9, 14, 9) {real, imag} */,
  {32'hbf5ede62, 32'hbec4e848} /* (9, 14, 8) {real, imag} */,
  {32'hbf95be27, 32'hbf4b8029} /* (9, 14, 7) {real, imag} */,
  {32'h3f428da1, 32'hc03362f4} /* (9, 14, 6) {real, imag} */,
  {32'h3fff8d05, 32'hc00aa3ae} /* (9, 14, 5) {real, imag} */,
  {32'h3fd802d4, 32'h3f9c9586} /* (9, 14, 4) {real, imag} */,
  {32'h40052f91, 32'hbeb97316} /* (9, 14, 3) {real, imag} */,
  {32'hbf19ebc2, 32'hbe814f18} /* (9, 14, 2) {real, imag} */,
  {32'hbfaca183, 32'h3fb105b9} /* (9, 14, 1) {real, imag} */,
  {32'hbd1ce38c, 32'h3f9ace24} /* (9, 14, 0) {real, imag} */,
  {32'hbf825468, 32'hbeeb30b4} /* (9, 13, 15) {real, imag} */,
  {32'hc03d75ee, 32'hbf7d20fb} /* (9, 13, 14) {real, imag} */,
  {32'hc01b91aa, 32'h3e155188} /* (9, 13, 13) {real, imag} */,
  {32'h3f26bc74, 32'h401ef07e} /* (9, 13, 12) {real, imag} */,
  {32'h3f89c6f4, 32'h3fe3f676} /* (9, 13, 11) {real, imag} */,
  {32'hbef7c688, 32'hbcf81800} /* (9, 13, 10) {real, imag} */,
  {32'hbe5a60b4, 32'hbf85b907} /* (9, 13, 9) {real, imag} */,
  {32'hbf2b097d, 32'hbf7f8fd4} /* (9, 13, 8) {real, imag} */,
  {32'h3fa54be8, 32'hbf86490c} /* (9, 13, 7) {real, imag} */,
  {32'h3e5fd120, 32'hc07b4800} /* (9, 13, 6) {real, imag} */,
  {32'hc007952a, 32'hc0762267} /* (9, 13, 5) {real, imag} */,
  {32'hbdba3562, 32'hbf8d9e26} /* (9, 13, 4) {real, imag} */,
  {32'hbfc4dee6, 32'hbf26c3ac} /* (9, 13, 3) {real, imag} */,
  {32'hbe113408, 32'hbf88c6c8} /* (9, 13, 2) {real, imag} */,
  {32'h3e51d2f4, 32'hbfc1bbb0} /* (9, 13, 1) {real, imag} */,
  {32'hbf226abb, 32'hbe0ae334} /* (9, 13, 0) {real, imag} */,
  {32'hbf0de03e, 32'h3e112c32} /* (9, 12, 15) {real, imag} */,
  {32'hbfc02f27, 32'h40060cb0} /* (9, 12, 14) {real, imag} */,
  {32'hc02d9a80, 32'h3fb3a36a} /* (9, 12, 13) {real, imag} */,
  {32'hbfcb902c, 32'h3d7bc520} /* (9, 12, 12) {real, imag} */,
  {32'hbe8da824, 32'hbede6087} /* (9, 12, 11) {real, imag} */,
  {32'h3f10dcad, 32'hbd2e7ba0} /* (9, 12, 10) {real, imag} */,
  {32'h3f998bae, 32'hbdaedc40} /* (9, 12, 9) {real, imag} */,
  {32'h402df69e, 32'h3e364794} /* (9, 12, 8) {real, imag} */,
  {32'h402e0efc, 32'h3f542d0b} /* (9, 12, 7) {real, imag} */,
  {32'h40065f58, 32'hbf114b1d} /* (9, 12, 6) {real, imag} */,
  {32'h3fbc32ad, 32'hc05417c1} /* (9, 12, 5) {real, imag} */,
  {32'h3fe5d8f0, 32'hbfdc0bec} /* (9, 12, 4) {real, imag} */,
  {32'h3f927f6e, 32'h3eacccd3} /* (9, 12, 3) {real, imag} */,
  {32'h3e092fd4, 32'h3e8b3bd0} /* (9, 12, 2) {real, imag} */,
  {32'hbfacedf6, 32'h3f882df1} /* (9, 12, 1) {real, imag} */,
  {32'hbfb226c8, 32'h3fa4ce18} /* (9, 12, 0) {real, imag} */,
  {32'hbf130d5f, 32'h3f96336f} /* (9, 11, 15) {real, imag} */,
  {32'h3f2a9792, 32'h3f6e4bb7} /* (9, 11, 14) {real, imag} */,
  {32'h3fb56eb3, 32'h3e8e7008} /* (9, 11, 13) {real, imag} */,
  {32'h3cc23380, 32'hbf146e60} /* (9, 11, 12) {real, imag} */,
  {32'hc002e026, 32'h3f884766} /* (9, 11, 11) {real, imag} */,
  {32'hc01b1321, 32'h3fcd08c8} /* (9, 11, 10) {real, imag} */,
  {32'hbeb4b670, 32'h3efb7ec4} /* (9, 11, 9) {real, imag} */,
  {32'hbff84c8b, 32'hbf8a0749} /* (9, 11, 8) {real, imag} */,
  {32'hbfcdc48e, 32'hbfabfec2} /* (9, 11, 7) {real, imag} */,
  {32'hbf49b6f6, 32'h3ef58312} /* (9, 11, 6) {real, imag} */,
  {32'hbf8b0bd5, 32'h3f2e11b4} /* (9, 11, 5) {real, imag} */,
  {32'hbf9eb9a0, 32'h3da6f5ba} /* (9, 11, 4) {real, imag} */,
  {32'hbf813078, 32'hbf42140e} /* (9, 11, 3) {real, imag} */,
  {32'hbfbe420a, 32'hbf28234c} /* (9, 11, 2) {real, imag} */,
  {32'hbf9588d4, 32'h3eb3f338} /* (9, 11, 1) {real, imag} */,
  {32'hb9e6f800, 32'h3ea66392} /* (9, 11, 0) {real, imag} */,
  {32'hbd42f718, 32'h3ee2a8fa} /* (9, 10, 15) {real, imag} */,
  {32'hbc152600, 32'h3f2f8609} /* (9, 10, 14) {real, imag} */,
  {32'h3de7b630, 32'h3e90f100} /* (9, 10, 13) {real, imag} */,
  {32'hbfeec062, 32'h3f63123a} /* (9, 10, 12) {real, imag} */,
  {32'hbfe1bbba, 32'h3fee0f3f} /* (9, 10, 11) {real, imag} */,
  {32'h3f45ce3a, 32'h3e52728c} /* (9, 10, 10) {real, imag} */,
  {32'h3f998613, 32'h3efd5e56} /* (9, 10, 9) {real, imag} */,
  {32'h3f501c92, 32'h3e86ab1e} /* (9, 10, 8) {real, imag} */,
  {32'h3e31f7d2, 32'hbec47dec} /* (9, 10, 7) {real, imag} */,
  {32'hbec95786, 32'h3ec409c1} /* (9, 10, 6) {real, imag} */,
  {32'hbf129f02, 32'h3e301192} /* (9, 10, 5) {real, imag} */,
  {32'hbf0473a9, 32'h3eaf9ce8} /* (9, 10, 4) {real, imag} */,
  {32'h3f7ddae3, 32'h3fa69e8e} /* (9, 10, 3) {real, imag} */,
  {32'h40088ac6, 32'hbee0eae9} /* (9, 10, 2) {real, imag} */,
  {32'h3f070217, 32'h3f83eaec} /* (9, 10, 1) {real, imag} */,
  {32'hbd9f22c4, 32'h3fb33eae} /* (9, 10, 0) {real, imag} */,
  {32'hbf0aa12b, 32'h3e3b4eec} /* (9, 9, 15) {real, imag} */,
  {32'hbfe59330, 32'h3f67f0b8} /* (9, 9, 14) {real, imag} */,
  {32'hbf15ebb0, 32'h3ec42be8} /* (9, 9, 13) {real, imag} */,
  {32'h3f6bb75a, 32'hbf4bc32c} /* (9, 9, 12) {real, imag} */,
  {32'h3fd35190, 32'hbedd10f8} /* (9, 9, 11) {real, imag} */,
  {32'h3f822e25, 32'h3eb02c1a} /* (9, 9, 10) {real, imag} */,
  {32'h3f121c28, 32'h3d811310} /* (9, 9, 9) {real, imag} */,
  {32'h3f402337, 32'hbf89c6e2} /* (9, 9, 8) {real, imag} */,
  {32'hbf7834a0, 32'h3c9e9220} /* (9, 9, 7) {real, imag} */,
  {32'hbe677846, 32'hbeac8969} /* (9, 9, 6) {real, imag} */,
  {32'h3fb714bc, 32'hbe09a252} /* (9, 9, 5) {real, imag} */,
  {32'h3f5dd9a6, 32'hbec37be0} /* (9, 9, 4) {real, imag} */,
  {32'h3f3fdab5, 32'hbf3cd797} /* (9, 9, 3) {real, imag} */,
  {32'h3f12a42e, 32'hbedc406c} /* (9, 9, 2) {real, imag} */,
  {32'hbd9bdc78, 32'hbf0bcde4} /* (9, 9, 1) {real, imag} */,
  {32'hbdee7a11, 32'h3e038169} /* (9, 9, 0) {real, imag} */,
  {32'h3f23e2d0, 32'hbe061658} /* (9, 8, 15) {real, imag} */,
  {32'h3c9ff340, 32'h3e3574d4} /* (9, 8, 14) {real, imag} */,
  {32'hbe8111d4, 32'h3e0f1e68} /* (9, 8, 13) {real, imag} */,
  {32'h3e86a750, 32'hbe7f3bf8} /* (9, 8, 12) {real, imag} */,
  {32'hbe0d6288, 32'hbf10f956} /* (9, 8, 11) {real, imag} */,
  {32'h3e532750, 32'hbf2f7550} /* (9, 8, 10) {real, imag} */,
  {32'h3e8817fe, 32'hbe552196} /* (9, 8, 9) {real, imag} */,
  {32'h3d93a010, 32'h3f8129f2} /* (9, 8, 8) {real, imag} */,
  {32'hbe02f75b, 32'h3ecbd900} /* (9, 8, 7) {real, imag} */,
  {32'hbf184d44, 32'hbf2e2536} /* (9, 8, 6) {real, imag} */,
  {32'hbe9e0408, 32'h3ed5debe} /* (9, 8, 5) {real, imag} */,
  {32'hbe2719f4, 32'h3fb1dea2} /* (9, 8, 4) {real, imag} */,
  {32'hbd2257e8, 32'h3ebc314c} /* (9, 8, 3) {real, imag} */,
  {32'h3dad1708, 32'h3e5bbcb0} /* (9, 8, 2) {real, imag} */,
  {32'h3f46ffac, 32'h3e011270} /* (9, 8, 1) {real, imag} */,
  {32'h3f62b75a, 32'h3c48dc80} /* (9, 8, 0) {real, imag} */,
  {32'h3f0f2def, 32'h3ec4f856} /* (9, 7, 15) {real, imag} */,
  {32'h3eae4998, 32'h3f21ecba} /* (9, 7, 14) {real, imag} */,
  {32'hbeec9c1c, 32'h3f472820} /* (9, 7, 13) {real, imag} */,
  {32'hbf39a926, 32'h3e8aacb0} /* (9, 7, 12) {real, imag} */,
  {32'hbef7f408, 32'hbea65fe8} /* (9, 7, 11) {real, imag} */,
  {32'hbdd085d0, 32'hbf315a13} /* (9, 7, 10) {real, imag} */,
  {32'hbf175854, 32'hbea3d5fc} /* (9, 7, 9) {real, imag} */,
  {32'hbebc1e4a, 32'hbee028a2} /* (9, 7, 8) {real, imag} */,
  {32'hbebfeca7, 32'hbf2427df} /* (9, 7, 7) {real, imag} */,
  {32'hbe00da22, 32'hbe586dde} /* (9, 7, 6) {real, imag} */,
  {32'hbf2abb95, 32'hbd8d5764} /* (9, 7, 5) {real, imag} */,
  {32'hbfd1b82f, 32'hbe504c60} /* (9, 7, 4) {real, imag} */,
  {32'hbf39dccb, 32'hbf0b7a03} /* (9, 7, 3) {real, imag} */,
  {32'h3f332a8e, 32'hbe2cfa78} /* (9, 7, 2) {real, imag} */,
  {32'h3f806ea0, 32'h3e5cece0} /* (9, 7, 1) {real, imag} */,
  {32'h3e968884, 32'hbd86ddee} /* (9, 7, 0) {real, imag} */,
  {32'hbe920b21, 32'h3e332b5d} /* (9, 6, 15) {real, imag} */,
  {32'h3d824460, 32'h3f309217} /* (9, 6, 14) {real, imag} */,
  {32'hbf0dc7c6, 32'h3eacaa72} /* (9, 6, 13) {real, imag} */,
  {32'h3eb11900, 32'h3f48b992} /* (9, 6, 12) {real, imag} */,
  {32'h3f62253c, 32'h3f5bece2} /* (9, 6, 11) {real, imag} */,
  {32'h3d5e3640, 32'h3f6448af} /* (9, 6, 10) {real, imag} */,
  {32'hbf40a1ce, 32'h3fae68ca} /* (9, 6, 9) {real, imag} */,
  {32'hbdab1d74, 32'h3fe083de} /* (9, 6, 8) {real, imag} */,
  {32'h3e0466a2, 32'h3d807ec2} /* (9, 6, 7) {real, imag} */,
  {32'hbf29afa9, 32'hbe693026} /* (9, 6, 6) {real, imag} */,
  {32'hbf5387d2, 32'hbee034bf} /* (9, 6, 5) {real, imag} */,
  {32'h3e9cf016, 32'h3f9e94d2} /* (9, 6, 4) {real, imag} */,
  {32'h3f1bca55, 32'h3ee04622} /* (9, 6, 3) {real, imag} */,
  {32'h3f8bb0fe, 32'hbee2e8bf} /* (9, 6, 2) {real, imag} */,
  {32'h3fc73f58, 32'h3ee5f33e} /* (9, 6, 1) {real, imag} */,
  {32'h3f5fd03a, 32'hbea57296} /* (9, 6, 0) {real, imag} */,
  {32'hbfc74586, 32'h3f6b6fbe} /* (9, 5, 15) {real, imag} */,
  {32'hbfe99a71, 32'h3fdae71c} /* (9, 5, 14) {real, imag} */,
  {32'h3eae6370, 32'h3fda0068} /* (9, 5, 13) {real, imag} */,
  {32'h3f843590, 32'h3f97a258} /* (9, 5, 12) {real, imag} */,
  {32'h3face730, 32'h3e349ad0} /* (9, 5, 11) {real, imag} */,
  {32'h3ee4ec3a, 32'hbe503000} /* (9, 5, 10) {real, imag} */,
  {32'h3fe8289c, 32'hbfd7e2c1} /* (9, 5, 9) {real, imag} */,
  {32'h4019d62d, 32'hbfd8da3b} /* (9, 5, 8) {real, imag} */,
  {32'h3ec97028, 32'hbff9ae90} /* (9, 5, 7) {real, imag} */,
  {32'hbef1535b, 32'hbf49e2a5} /* (9, 5, 6) {real, imag} */,
  {32'hbf27ad16, 32'h3f11c5cc} /* (9, 5, 5) {real, imag} */,
  {32'hbee8cb26, 32'hbcb26558} /* (9, 5, 4) {real, imag} */,
  {32'hbf1f05a6, 32'hbcabfe30} /* (9, 5, 3) {real, imag} */,
  {32'hbeb43766, 32'h3ea15504} /* (9, 5, 2) {real, imag} */,
  {32'hbf2bf545, 32'h401f7605} /* (9, 5, 1) {real, imag} */,
  {32'hbf9ba75e, 32'h3f7acd11} /* (9, 5, 0) {real, imag} */,
  {32'h3f0a89b6, 32'h3f3defdc} /* (9, 4, 15) {real, imag} */,
  {32'hbef18bb4, 32'h3f3b741a} /* (9, 4, 14) {real, imag} */,
  {32'hbf721a40, 32'h3f81b6b6} /* (9, 4, 13) {real, imag} */,
  {32'h3fbe5876, 32'h3e525dd8} /* (9, 4, 12) {real, imag} */,
  {32'h4007a2f2, 32'hbf5b20b8} /* (9, 4, 11) {real, imag} */,
  {32'hbf465c47, 32'hc043a6e8} /* (9, 4, 10) {real, imag} */,
  {32'hbfa54bae, 32'hc0658e12} /* (9, 4, 9) {real, imag} */,
  {32'hbff7243c, 32'hbfe3040a} /* (9, 4, 8) {real, imag} */,
  {32'hc00727a8, 32'hbe6b686c} /* (9, 4, 7) {real, imag} */,
  {32'hbf8b815c, 32'h3e806842} /* (9, 4, 6) {real, imag} */,
  {32'hc00d7b3c, 32'h3d785b40} /* (9, 4, 5) {real, imag} */,
  {32'hbfa065dc, 32'hbfa5afcc} /* (9, 4, 4) {real, imag} */,
  {32'h3fdb840c, 32'h3f4fce16} /* (9, 4, 3) {real, imag} */,
  {32'h3fcd71da, 32'h40241046} /* (9, 4, 2) {real, imag} */,
  {32'h3f699e63, 32'h3f8a0fc3} /* (9, 4, 1) {real, imag} */,
  {32'h40117979, 32'h3eec887e} /* (9, 4, 0) {real, imag} */,
  {32'hbf61add5, 32'hbfc84bfd} /* (9, 3, 15) {real, imag} */,
  {32'hc0164560, 32'hbffb73a2} /* (9, 3, 14) {real, imag} */,
  {32'hbfd7f350, 32'hbff2e4d1} /* (9, 3, 13) {real, imag} */,
  {32'hbf062050, 32'h3fa65811} /* (9, 3, 12) {real, imag} */,
  {32'hbd5fccb0, 32'h3fba9862} /* (9, 3, 11) {real, imag} */,
  {32'h3f23d072, 32'hc0325c10} /* (9, 3, 10) {real, imag} */,
  {32'h3e88a4ca, 32'hbff0a2f5} /* (9, 3, 9) {real, imag} */,
  {32'h3eedf672, 32'hbf90120e} /* (9, 3, 8) {real, imag} */,
  {32'hbd320210, 32'hbf693403} /* (9, 3, 7) {real, imag} */,
  {32'hbf1a27fd, 32'hbe252980} /* (9, 3, 6) {real, imag} */,
  {32'hc008905a, 32'h3fc592ba} /* (9, 3, 5) {real, imag} */,
  {32'hba568b00, 32'h3f32d565} /* (9, 3, 4) {real, imag} */,
  {32'h3f4bb5fb, 32'h3f997e88} /* (9, 3, 3) {real, imag} */,
  {32'h3e869fc4, 32'h3ed2c2a4} /* (9, 3, 2) {real, imag} */,
  {32'hbf91e974, 32'hbffb3c74} /* (9, 3, 1) {real, imag} */,
  {32'hbed7d5e2, 32'hbf83d5ea} /* (9, 3, 0) {real, imag} */,
  {32'hbfbd69bc, 32'hbfc3efde} /* (9, 2, 15) {real, imag} */,
  {32'hc01dd31e, 32'hc07fa064} /* (9, 2, 14) {real, imag} */,
  {32'hbfb980a4, 32'hbe8cf577} /* (9, 2, 13) {real, imag} */,
  {32'h3f9ec25e, 32'h3f4d3e7e} /* (9, 2, 12) {real, imag} */,
  {32'h3fd9ba87, 32'hbf286b43} /* (9, 2, 11) {real, imag} */,
  {32'h400f54e7, 32'h3f75d0d5} /* (9, 2, 10) {real, imag} */,
  {32'h3fe70780, 32'h409172a6} /* (9, 2, 9) {real, imag} */,
  {32'h3f9cf76b, 32'h40a26a6a} /* (9, 2, 8) {real, imag} */,
  {32'h3ffb1c51, 32'h3e13cac4} /* (9, 2, 7) {real, imag} */,
  {32'h3ffbc2f6, 32'h3f2e94c8} /* (9, 2, 6) {real, imag} */,
  {32'hc02525f8, 32'hbd735160} /* (9, 2, 5) {real, imag} */,
  {32'hbf944250, 32'hbf4da564} /* (9, 2, 4) {real, imag} */,
  {32'h4024a473, 32'hbefe04b8} /* (9, 2, 3) {real, imag} */,
  {32'h405ebc5c, 32'h3f4b9e20} /* (9, 2, 2) {real, imag} */,
  {32'hbcc94c00, 32'h3f8be0b5} /* (9, 2, 1) {real, imag} */,
  {32'hbe5d2517, 32'hbdad5cc8} /* (9, 2, 0) {real, imag} */,
  {32'h3f53121f, 32'hbf4a7330} /* (9, 1, 15) {real, imag} */,
  {32'h3fa0cc40, 32'h3f82e401} /* (9, 1, 14) {real, imag} */,
  {32'h3f915d4f, 32'h3dfc1e88} /* (9, 1, 13) {real, imag} */,
  {32'h3f76fb5e, 32'hbd6bcfc0} /* (9, 1, 12) {real, imag} */,
  {32'hbf8b8db0, 32'hbe229660} /* (9, 1, 11) {real, imag} */,
  {32'h3e301688, 32'hc07b8d0a} /* (9, 1, 10) {real, imag} */,
  {32'hc07e1ed0, 32'hc0bf3557} /* (9, 1, 9) {real, imag} */,
  {32'hbff2a62e, 32'hc01b292d} /* (9, 1, 8) {real, imag} */,
  {32'h4002f6d2, 32'h4002a096} /* (9, 1, 7) {real, imag} */,
  {32'h3ebea9a6, 32'h400ef8a6} /* (9, 1, 6) {real, imag} */,
  {32'h405643f3, 32'h40277320} /* (9, 1, 5) {real, imag} */,
  {32'h402f0d29, 32'h3f8336d6} /* (9, 1, 4) {real, imag} */,
  {32'hbf7a6579, 32'h400beaf8} /* (9, 1, 3) {real, imag} */,
  {32'hc0303c75, 32'h40b32b58} /* (9, 1, 2) {real, imag} */,
  {32'hbeaa278a, 32'h4010da18} /* (9, 1, 1) {real, imag} */,
  {32'h3ec5e118, 32'h3f874781} /* (9, 1, 0) {real, imag} */,
  {32'h3f627bc8, 32'hc03143d4} /* (9, 0, 15) {real, imag} */,
  {32'h403e19c2, 32'hbf77da87} /* (9, 0, 14) {real, imag} */,
  {32'hbea57b0c, 32'hbfaa8875} /* (9, 0, 13) {real, imag} */,
  {32'hc0178427, 32'hbfe29bcd} /* (9, 0, 12) {real, imag} */,
  {32'h3fbf4b11, 32'h405f6944} /* (9, 0, 11) {real, imag} */,
  {32'hbf102a08, 32'h4094925c} /* (9, 0, 10) {real, imag} */,
  {32'h3ed9c042, 32'h3f08fdd6} /* (9, 0, 9) {real, imag} */,
  {32'hbfd5e124, 32'h3df64118} /* (9, 0, 8) {real, imag} */,
  {32'hbed2bdc4, 32'hc085ca5c} /* (9, 0, 7) {real, imag} */,
  {32'h3e0401f8, 32'hc038ba4c} /* (9, 0, 6) {real, imag} */,
  {32'h404a136d, 32'hbec4325a} /* (9, 0, 5) {real, imag} */,
  {32'h3fdfc706, 32'hbf57c6f5} /* (9, 0, 4) {real, imag} */,
  {32'hbf04face, 32'hc05e7b80} /* (9, 0, 3) {real, imag} */,
  {32'hbfee4b68, 32'hc063accb} /* (9, 0, 2) {real, imag} */,
  {32'h3f59f37e, 32'hc0759c31} /* (9, 0, 1) {real, imag} */,
  {32'h3f0f64dc, 32'hc00a9870} /* (9, 0, 0) {real, imag} */,
  {32'hbf45d614, 32'hc0141257} /* (8, 15, 15) {real, imag} */,
  {32'hbfcb3abb, 32'hbf3ba5ff} /* (8, 15, 14) {real, imag} */,
  {32'hbfcff98c, 32'h3e17fabe} /* (8, 15, 13) {real, imag} */,
  {32'hbe858f19, 32'h3f7b9c23} /* (8, 15, 12) {real, imag} */,
  {32'hbfbd7010, 32'h4027f912} /* (8, 15, 11) {real, imag} */,
  {32'h3f90b0a8, 32'h403763c1} /* (8, 15, 10) {real, imag} */,
  {32'h3f8da351, 32'h40280d80} /* (8, 15, 9) {real, imag} */,
  {32'hc00e4f72, 32'hbee01bab} /* (8, 15, 8) {real, imag} */,
  {32'hbf4b5bea, 32'hbfe83028} /* (8, 15, 7) {real, imag} */,
  {32'h3ee87c9e, 32'hbc35ed00} /* (8, 15, 6) {real, imag} */,
  {32'h3f8fdfc6, 32'h3f7b4314} /* (8, 15, 5) {real, imag} */,
  {32'h3fe10908, 32'h3fda50c8} /* (8, 15, 4) {real, imag} */,
  {32'h40073ca5, 32'hbfa11f8b} /* (8, 15, 3) {real, imag} */,
  {32'h3f58250e, 32'hbf017e38} /* (8, 15, 2) {real, imag} */,
  {32'hbf460598, 32'hbedbfa5a} /* (8, 15, 1) {real, imag} */,
  {32'hbff982cd, 32'hbfa13a3c} /* (8, 15, 0) {real, imag} */,
  {32'h3e08e782, 32'hbff67b43} /* (8, 14, 15) {real, imag} */,
  {32'hbe0cdedd, 32'hbee962f2} /* (8, 14, 14) {real, imag} */,
  {32'h3f78d899, 32'h3dddeb0c} /* (8, 14, 13) {real, imag} */,
  {32'h3fb31d9c, 32'hbd168f50} /* (8, 14, 12) {real, imag} */,
  {32'h4033b1d6, 32'hc016f10e} /* (8, 14, 11) {real, imag} */,
  {32'h3f08ead6, 32'h4012f125} /* (8, 14, 10) {real, imag} */,
  {32'h3f225027, 32'h408fa2d1} /* (8, 14, 9) {real, imag} */,
  {32'h3f811c33, 32'h4028f300} /* (8, 14, 8) {real, imag} */,
  {32'h3e16556e, 32'h4041c32c} /* (8, 14, 7) {real, imag} */,
  {32'hc034d77a, 32'h402eebaa} /* (8, 14, 6) {real, imag} */,
  {32'hc056d557, 32'hbe74dd8d} /* (8, 14, 5) {real, imag} */,
  {32'hbfa0b2e9, 32'hbee66144} /* (8, 14, 4) {real, imag} */,
  {32'h3ec23232, 32'h3e766dd4} /* (8, 14, 3) {real, imag} */,
  {32'hbdec1b09, 32'hbeb28a33} /* (8, 14, 2) {real, imag} */,
  {32'hc02c616a, 32'h3dd80ed1} /* (8, 14, 1) {real, imag} */,
  {32'hbea3c2ab, 32'h3f894096} /* (8, 14, 0) {real, imag} */,
  {32'hbfd6e7dd, 32'hbf0541fd} /* (8, 13, 15) {real, imag} */,
  {32'h3e4ac6d4, 32'hbd86e2a8} /* (8, 13, 14) {real, imag} */,
  {32'hbf85203b, 32'hbf673dfa} /* (8, 13, 13) {real, imag} */,
  {32'hbfab38f5, 32'hc025a44e} /* (8, 13, 12) {real, imag} */,
  {32'hbface369, 32'hbf5c69ab} /* (8, 13, 11) {real, imag} */,
  {32'hc02bb0ee, 32'h3e8c85e6} /* (8, 13, 10) {real, imag} */,
  {32'h3fa82bd6, 32'h3ff29408} /* (8, 13, 9) {real, imag} */,
  {32'h3faba187, 32'hbd2f2bb8} /* (8, 13, 8) {real, imag} */,
  {32'hbf7af9f8, 32'h3f630aaa} /* (8, 13, 7) {real, imag} */,
  {32'hbe703fc8, 32'h3e412ce8} /* (8, 13, 6) {real, imag} */,
  {32'h3ff6a051, 32'h3f44490a} /* (8, 13, 5) {real, imag} */,
  {32'h3f6013b7, 32'h40082474} /* (8, 13, 4) {real, imag} */,
  {32'h3ed357cd, 32'h3fb22346} /* (8, 13, 3) {real, imag} */,
  {32'hbf5f85d1, 32'hbe8ffdae} /* (8, 13, 2) {real, imag} */,
  {32'hbf81174e, 32'hbf48821c} /* (8, 13, 1) {real, imag} */,
  {32'hbfb7cde2, 32'h3e9b77ce} /* (8, 13, 0) {real, imag} */,
  {32'hbf2ea370, 32'hbf3129df} /* (8, 12, 15) {real, imag} */,
  {32'h3e7ad61c, 32'hbfc7f9db} /* (8, 12, 14) {real, imag} */,
  {32'h3fb1dd73, 32'hbfc8d3ae} /* (8, 12, 13) {real, imag} */,
  {32'h3f8e3a67, 32'h3d030608} /* (8, 12, 12) {real, imag} */,
  {32'h3e5a8ece, 32'h3f01f4bb} /* (8, 12, 11) {real, imag} */,
  {32'h3fbf410c, 32'h3e9778a7} /* (8, 12, 10) {real, imag} */,
  {32'h403faae1, 32'hbfa761d1} /* (8, 12, 9) {real, imag} */,
  {32'h3fd8cb06, 32'hc026c692} /* (8, 12, 8) {real, imag} */,
  {32'h3fcd66e0, 32'hbfebd216} /* (8, 12, 7) {real, imag} */,
  {32'h3d4711e0, 32'hbf897823} /* (8, 12, 6) {real, imag} */,
  {32'h3db6a3e0, 32'hbf12afc5} /* (8, 12, 5) {real, imag} */,
  {32'hc01c78de, 32'hbf2a2fa1} /* (8, 12, 4) {real, imag} */,
  {32'hc007c743, 32'hbe2c04b4} /* (8, 12, 3) {real, imag} */,
  {32'hbfd83bc3, 32'hbf19e3f4} /* (8, 12, 2) {real, imag} */,
  {32'h3d2b1450, 32'h3f08c5c7} /* (8, 12, 1) {real, imag} */,
  {32'h3e3fd43c, 32'hbe99cec0} /* (8, 12, 0) {real, imag} */,
  {32'h3ec38484, 32'h3f15fe67} /* (8, 11, 15) {real, imag} */,
  {32'hbf70a77b, 32'h3f54a06b} /* (8, 11, 14) {real, imag} */,
  {32'hbd8bb86c, 32'h3eb9da55} /* (8, 11, 13) {real, imag} */,
  {32'h3f809173, 32'hbf5df2de} /* (8, 11, 12) {real, imag} */,
  {32'h3f7b9f82, 32'hbefa559a} /* (8, 11, 11) {real, imag} */,
  {32'h3efd8970, 32'hbefc86fe} /* (8, 11, 10) {real, imag} */,
  {32'hbedd01e6, 32'h3f026484} /* (8, 11, 9) {real, imag} */,
  {32'hbf34ec72, 32'h3ef15117} /* (8, 11, 8) {real, imag} */,
  {32'hbf6078ec, 32'hbe8d0308} /* (8, 11, 7) {real, imag} */,
  {32'h3f8ff46b, 32'hc00ed658} /* (8, 11, 6) {real, imag} */,
  {32'h400266c2, 32'hc00a672e} /* (8, 11, 5) {real, imag} */,
  {32'h3ff5862c, 32'hbf92bbfa} /* (8, 11, 4) {real, imag} */,
  {32'h3ee07cbf, 32'hbf09b8d5} /* (8, 11, 3) {real, imag} */,
  {32'hbea2fb26, 32'hbf055ac9} /* (8, 11, 2) {real, imag} */,
  {32'hbe8967c8, 32'h3ec759cc} /* (8, 11, 1) {real, imag} */,
  {32'h3f98dc0e, 32'h3f9095f0} /* (8, 11, 0) {real, imag} */,
  {32'h3e8a9373, 32'hbf459e9e} /* (8, 10, 15) {real, imag} */,
  {32'h3e53a661, 32'hbf284d9d} /* (8, 10, 14) {real, imag} */,
  {32'h3eac4d9e, 32'hbe338d5a} /* (8, 10, 13) {real, imag} */,
  {32'h3f3dada8, 32'h3ea4b73e} /* (8, 10, 12) {real, imag} */,
  {32'hbe60af58, 32'hbe19b488} /* (8, 10, 11) {real, imag} */,
  {32'hbf079090, 32'hbf3ef568} /* (8, 10, 10) {real, imag} */,
  {32'hbfac28c0, 32'h3ee3a7f0} /* (8, 10, 9) {real, imag} */,
  {32'hbf017f4e, 32'h3ec67cf4} /* (8, 10, 8) {real, imag} */,
  {32'h3e8625a7, 32'h3daaf1e0} /* (8, 10, 7) {real, imag} */,
  {32'hbeb18cbc, 32'h3f207e1a} /* (8, 10, 6) {real, imag} */,
  {32'hbe1d3280, 32'h3eed665a} /* (8, 10, 5) {real, imag} */,
  {32'h3f130328, 32'h3f3c054c} /* (8, 10, 4) {real, imag} */,
  {32'h3e68b804, 32'h3f9f342e} /* (8, 10, 3) {real, imag} */,
  {32'hbea00108, 32'h3faa9a67} /* (8, 10, 2) {real, imag} */,
  {32'hbf26ea72, 32'hbd9a97bf} /* (8, 10, 1) {real, imag} */,
  {32'hbf0cca11, 32'hbee3f7e7} /* (8, 10, 0) {real, imag} */,
  {32'hbf026dfc, 32'hbe7f00e0} /* (8, 9, 15) {real, imag} */,
  {32'hbe888338, 32'hbe5a0cc4} /* (8, 9, 14) {real, imag} */,
  {32'h3aee1000, 32'hbe5130fa} /* (8, 9, 13) {real, imag} */,
  {32'h3e256dce, 32'hbf5f301d} /* (8, 9, 12) {real, imag} */,
  {32'h3f0db294, 32'hbf25b487} /* (8, 9, 11) {real, imag} */,
  {32'h3f3a57b8, 32'hbf21de5c} /* (8, 9, 10) {real, imag} */,
  {32'h3ea6e0a7, 32'hbf610a5a} /* (8, 9, 9) {real, imag} */,
  {32'h3e916508, 32'hbf093781} /* (8, 9, 8) {real, imag} */,
  {32'h3f53b540, 32'hbe864076} /* (8, 9, 7) {real, imag} */,
  {32'hbe5d018b, 32'h3f74dca0} /* (8, 9, 6) {real, imag} */,
  {32'hbf4c0d61, 32'h3e9e57f8} /* (8, 9, 5) {real, imag} */,
  {32'hbf0923b0, 32'hbe6cee0c} /* (8, 9, 4) {real, imag} */,
  {32'h3f08524d, 32'hbe949584} /* (8, 9, 3) {real, imag} */,
  {32'h3ecb9b9c, 32'hbefd4118} /* (8, 9, 2) {real, imag} */,
  {32'h3eeda6ad, 32'h3ae79a00} /* (8, 9, 1) {real, imag} */,
  {32'h3e6e5078, 32'h3d607130} /* (8, 9, 0) {real, imag} */,
  {32'h3f34a683, 32'h00000000} /* (8, 8, 15) {real, imag} */,
  {32'h3f13412a, 32'h00000000} /* (8, 8, 14) {real, imag} */,
  {32'h3bcbbf80, 32'h00000000} /* (8, 8, 13) {real, imag} */,
  {32'hbc86b710, 32'h00000000} /* (8, 8, 12) {real, imag} */,
  {32'hbddae1fc, 32'h00000000} /* (8, 8, 11) {real, imag} */,
  {32'hbf2f5d1a, 32'h00000000} /* (8, 8, 10) {real, imag} */,
  {32'hbfcc2ac7, 32'h00000000} /* (8, 8, 9) {real, imag} */,
  {32'hbeab31ba, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'hbf41bd79, 32'h00000000} /* (8, 8, 7) {real, imag} */,
  {32'hbe4cb820, 32'h00000000} /* (8, 8, 6) {real, imag} */,
  {32'hbea2131e, 32'h00000000} /* (8, 8, 5) {real, imag} */,
  {32'hbedc8420, 32'h00000000} /* (8, 8, 4) {real, imag} */,
  {32'h3f10d20e, 32'h00000000} /* (8, 8, 3) {real, imag} */,
  {32'h3f60c130, 32'h00000000} /* (8, 8, 2) {real, imag} */,
  {32'h3f6b7377, 32'h00000000} /* (8, 8, 1) {real, imag} */,
  {32'h3ea75156, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'hbf026dfc, 32'h3e7f00e0} /* (8, 7, 15) {real, imag} */,
  {32'hbe888338, 32'h3e5a0cc4} /* (8, 7, 14) {real, imag} */,
  {32'h3aee1000, 32'h3e5130fa} /* (8, 7, 13) {real, imag} */,
  {32'h3e256dce, 32'h3f5f301d} /* (8, 7, 12) {real, imag} */,
  {32'h3f0db294, 32'h3f25b487} /* (8, 7, 11) {real, imag} */,
  {32'h3f3a57b8, 32'h3f21de5c} /* (8, 7, 10) {real, imag} */,
  {32'h3ea6e0a7, 32'h3f610a5a} /* (8, 7, 9) {real, imag} */,
  {32'h3e916508, 32'h3f093781} /* (8, 7, 8) {real, imag} */,
  {32'h3f53b540, 32'h3e864076} /* (8, 7, 7) {real, imag} */,
  {32'hbe5d018b, 32'hbf74dca0} /* (8, 7, 6) {real, imag} */,
  {32'hbf4c0d61, 32'hbe9e57f8} /* (8, 7, 5) {real, imag} */,
  {32'hbf0923b0, 32'h3e6cee0c} /* (8, 7, 4) {real, imag} */,
  {32'h3f08524d, 32'h3e949584} /* (8, 7, 3) {real, imag} */,
  {32'h3ecb9b9c, 32'h3efd4118} /* (8, 7, 2) {real, imag} */,
  {32'h3eeda6ad, 32'hbae79a00} /* (8, 7, 1) {real, imag} */,
  {32'h3e6e5078, 32'hbd607130} /* (8, 7, 0) {real, imag} */,
  {32'h3e8a9373, 32'h3f459e9e} /* (8, 6, 15) {real, imag} */,
  {32'h3e53a661, 32'h3f284d9d} /* (8, 6, 14) {real, imag} */,
  {32'h3eac4d9e, 32'h3e338d5a} /* (8, 6, 13) {real, imag} */,
  {32'h3f3dada8, 32'hbea4b73e} /* (8, 6, 12) {real, imag} */,
  {32'hbe60af58, 32'h3e19b488} /* (8, 6, 11) {real, imag} */,
  {32'hbf079090, 32'h3f3ef568} /* (8, 6, 10) {real, imag} */,
  {32'hbfac28c0, 32'hbee3a7f0} /* (8, 6, 9) {real, imag} */,
  {32'hbf017f4e, 32'hbec67cf4} /* (8, 6, 8) {real, imag} */,
  {32'h3e8625a7, 32'hbdaaf1e0} /* (8, 6, 7) {real, imag} */,
  {32'hbeb18cbc, 32'hbf207e1a} /* (8, 6, 6) {real, imag} */,
  {32'hbe1d3280, 32'hbeed665a} /* (8, 6, 5) {real, imag} */,
  {32'h3f130328, 32'hbf3c054c} /* (8, 6, 4) {real, imag} */,
  {32'h3e68b804, 32'hbf9f342e} /* (8, 6, 3) {real, imag} */,
  {32'hbea00108, 32'hbfaa9a67} /* (8, 6, 2) {real, imag} */,
  {32'hbf26ea72, 32'h3d9a97bf} /* (8, 6, 1) {real, imag} */,
  {32'hbf0cca11, 32'h3ee3f7e7} /* (8, 6, 0) {real, imag} */,
  {32'h3ec38484, 32'hbf15fe67} /* (8, 5, 15) {real, imag} */,
  {32'hbf70a77b, 32'hbf54a06b} /* (8, 5, 14) {real, imag} */,
  {32'hbd8bb86c, 32'hbeb9da55} /* (8, 5, 13) {real, imag} */,
  {32'h3f809173, 32'h3f5df2de} /* (8, 5, 12) {real, imag} */,
  {32'h3f7b9f82, 32'h3efa559a} /* (8, 5, 11) {real, imag} */,
  {32'h3efd8970, 32'h3efc86fe} /* (8, 5, 10) {real, imag} */,
  {32'hbedd01e6, 32'hbf026484} /* (8, 5, 9) {real, imag} */,
  {32'hbf34ec72, 32'hbef15117} /* (8, 5, 8) {real, imag} */,
  {32'hbf6078ec, 32'h3e8d0308} /* (8, 5, 7) {real, imag} */,
  {32'h3f8ff46b, 32'h400ed658} /* (8, 5, 6) {real, imag} */,
  {32'h400266c2, 32'h400a672e} /* (8, 5, 5) {real, imag} */,
  {32'h3ff5862c, 32'h3f92bbfa} /* (8, 5, 4) {real, imag} */,
  {32'h3ee07cbf, 32'h3f09b8d5} /* (8, 5, 3) {real, imag} */,
  {32'hbea2fb26, 32'h3f055ac9} /* (8, 5, 2) {real, imag} */,
  {32'hbe8967c8, 32'hbec759cc} /* (8, 5, 1) {real, imag} */,
  {32'h3f98dc0e, 32'hbf9095f0} /* (8, 5, 0) {real, imag} */,
  {32'hbf2ea370, 32'h3f3129df} /* (8, 4, 15) {real, imag} */,
  {32'h3e7ad61c, 32'h3fc7f9db} /* (8, 4, 14) {real, imag} */,
  {32'h3fb1dd73, 32'h3fc8d3ae} /* (8, 4, 13) {real, imag} */,
  {32'h3f8e3a67, 32'hbd030608} /* (8, 4, 12) {real, imag} */,
  {32'h3e5a8ece, 32'hbf01f4bb} /* (8, 4, 11) {real, imag} */,
  {32'h3fbf410c, 32'hbe9778a7} /* (8, 4, 10) {real, imag} */,
  {32'h403faae1, 32'h3fa761d1} /* (8, 4, 9) {real, imag} */,
  {32'h3fd8cb06, 32'h4026c692} /* (8, 4, 8) {real, imag} */,
  {32'h3fcd66e0, 32'h3febd216} /* (8, 4, 7) {real, imag} */,
  {32'h3d4711e0, 32'h3f897823} /* (8, 4, 6) {real, imag} */,
  {32'h3db6a3e0, 32'h3f12afc5} /* (8, 4, 5) {real, imag} */,
  {32'hc01c78de, 32'h3f2a2fa1} /* (8, 4, 4) {real, imag} */,
  {32'hc007c743, 32'h3e2c04b4} /* (8, 4, 3) {real, imag} */,
  {32'hbfd83bc3, 32'h3f19e3f4} /* (8, 4, 2) {real, imag} */,
  {32'h3d2b1450, 32'hbf08c5c7} /* (8, 4, 1) {real, imag} */,
  {32'h3e3fd43c, 32'h3e99cec0} /* (8, 4, 0) {real, imag} */,
  {32'hbfd6e7dd, 32'h3f0541fd} /* (8, 3, 15) {real, imag} */,
  {32'h3e4ac6d4, 32'h3d86e2a8} /* (8, 3, 14) {real, imag} */,
  {32'hbf85203b, 32'h3f673dfa} /* (8, 3, 13) {real, imag} */,
  {32'hbfab38f5, 32'h4025a44e} /* (8, 3, 12) {real, imag} */,
  {32'hbface369, 32'h3f5c69ab} /* (8, 3, 11) {real, imag} */,
  {32'hc02bb0ee, 32'hbe8c85e6} /* (8, 3, 10) {real, imag} */,
  {32'h3fa82bd6, 32'hbff29408} /* (8, 3, 9) {real, imag} */,
  {32'h3faba187, 32'h3d2f2bb8} /* (8, 3, 8) {real, imag} */,
  {32'hbf7af9f8, 32'hbf630aaa} /* (8, 3, 7) {real, imag} */,
  {32'hbe703fc8, 32'hbe412ce8} /* (8, 3, 6) {real, imag} */,
  {32'h3ff6a051, 32'hbf44490a} /* (8, 3, 5) {real, imag} */,
  {32'h3f6013b7, 32'hc0082474} /* (8, 3, 4) {real, imag} */,
  {32'h3ed357cd, 32'hbfb22346} /* (8, 3, 3) {real, imag} */,
  {32'hbf5f85d1, 32'h3e8ffdae} /* (8, 3, 2) {real, imag} */,
  {32'hbf81174e, 32'h3f48821c} /* (8, 3, 1) {real, imag} */,
  {32'hbfb7cde2, 32'hbe9b77ce} /* (8, 3, 0) {real, imag} */,
  {32'h3e08e782, 32'h3ff67b43} /* (8, 2, 15) {real, imag} */,
  {32'hbe0cdedd, 32'h3ee962f2} /* (8, 2, 14) {real, imag} */,
  {32'h3f78d899, 32'hbdddeb0c} /* (8, 2, 13) {real, imag} */,
  {32'h3fb31d9c, 32'h3d168f50} /* (8, 2, 12) {real, imag} */,
  {32'h4033b1d6, 32'h4016f10e} /* (8, 2, 11) {real, imag} */,
  {32'h3f08ead6, 32'hc012f125} /* (8, 2, 10) {real, imag} */,
  {32'h3f225027, 32'hc08fa2d1} /* (8, 2, 9) {real, imag} */,
  {32'h3f811c33, 32'hc028f300} /* (8, 2, 8) {real, imag} */,
  {32'h3e16556e, 32'hc041c32c} /* (8, 2, 7) {real, imag} */,
  {32'hc034d77a, 32'hc02eebaa} /* (8, 2, 6) {real, imag} */,
  {32'hc056d557, 32'h3e74dd8d} /* (8, 2, 5) {real, imag} */,
  {32'hbfa0b2e9, 32'h3ee66144} /* (8, 2, 4) {real, imag} */,
  {32'h3ec23232, 32'hbe766dd4} /* (8, 2, 3) {real, imag} */,
  {32'hbdec1b09, 32'h3eb28a33} /* (8, 2, 2) {real, imag} */,
  {32'hc02c616a, 32'hbdd80ed1} /* (8, 2, 1) {real, imag} */,
  {32'hbea3c2ab, 32'hbf894096} /* (8, 2, 0) {real, imag} */,
  {32'hbf45d614, 32'h40141257} /* (8, 1, 15) {real, imag} */,
  {32'hbfcb3abb, 32'h3f3ba5ff} /* (8, 1, 14) {real, imag} */,
  {32'hbfcff98c, 32'hbe17fabe} /* (8, 1, 13) {real, imag} */,
  {32'hbe858f19, 32'hbf7b9c23} /* (8, 1, 12) {real, imag} */,
  {32'hbfbd7010, 32'hc027f912} /* (8, 1, 11) {real, imag} */,
  {32'h3f90b0a8, 32'hc03763c1} /* (8, 1, 10) {real, imag} */,
  {32'h3f8da351, 32'hc0280d80} /* (8, 1, 9) {real, imag} */,
  {32'hc00e4f72, 32'h3ee01bab} /* (8, 1, 8) {real, imag} */,
  {32'hbf4b5bea, 32'h3fe83028} /* (8, 1, 7) {real, imag} */,
  {32'h3ee87c9e, 32'h3c35ed00} /* (8, 1, 6) {real, imag} */,
  {32'h3f8fdfc6, 32'hbf7b4314} /* (8, 1, 5) {real, imag} */,
  {32'h3fe10908, 32'hbfda50c8} /* (8, 1, 4) {real, imag} */,
  {32'h40073ca5, 32'h3fa11f8b} /* (8, 1, 3) {real, imag} */,
  {32'h3f58250e, 32'h3f017e38} /* (8, 1, 2) {real, imag} */,
  {32'hbf460598, 32'h3edbfa5a} /* (8, 1, 1) {real, imag} */,
  {32'hbff982cd, 32'h3fa13a3c} /* (8, 1, 0) {real, imag} */,
  {32'h401b19ed, 32'h00000000} /* (8, 0, 15) {real, imag} */,
  {32'h3fbed77b, 32'h00000000} /* (8, 0, 14) {real, imag} */,
  {32'hbc593cc0, 32'h00000000} /* (8, 0, 13) {real, imag} */,
  {32'hbed1a0b7, 32'h00000000} /* (8, 0, 12) {real, imag} */,
  {32'h3f73d21e, 32'h00000000} /* (8, 0, 11) {real, imag} */,
  {32'h3f6e3822, 32'h00000000} /* (8, 0, 10) {real, imag} */,
  {32'hbf1c7a4a, 32'h00000000} /* (8, 0, 9) {real, imag} */,
  {32'hbdfd28c8, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'hbfba83f0, 32'h00000000} /* (8, 0, 7) {real, imag} */,
  {32'h3f9e1b82, 32'h00000000} /* (8, 0, 6) {real, imag} */,
  {32'hbf693091, 32'h00000000} /* (8, 0, 5) {real, imag} */,
  {32'hbf35b25e, 32'h00000000} /* (8, 0, 4) {real, imag} */,
  {32'hbec81eac, 32'h00000000} /* (8, 0, 3) {real, imag} */,
  {32'h3e9f6fe9, 32'h00000000} /* (8, 0, 2) {real, imag} */,
  {32'h3e7d007c, 32'h00000000} /* (8, 0, 1) {real, imag} */,
  {32'h3f965602, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h3f53121f, 32'h3f4a7330} /* (7, 15, 15) {real, imag} */,
  {32'h3fa0cc40, 32'hbf82e401} /* (7, 15, 14) {real, imag} */,
  {32'h3f915d4f, 32'hbdfc1e88} /* (7, 15, 13) {real, imag} */,
  {32'h3f76fb5e, 32'h3d6bcfc0} /* (7, 15, 12) {real, imag} */,
  {32'hbf8b8db0, 32'h3e229660} /* (7, 15, 11) {real, imag} */,
  {32'h3e301688, 32'h407b8d0a} /* (7, 15, 10) {real, imag} */,
  {32'hc07e1ed0, 32'h40bf3557} /* (7, 15, 9) {real, imag} */,
  {32'hbff2a62e, 32'h401b292d} /* (7, 15, 8) {real, imag} */,
  {32'h4002f6d2, 32'hc002a096} /* (7, 15, 7) {real, imag} */,
  {32'h3ebea9a6, 32'hc00ef8a6} /* (7, 15, 6) {real, imag} */,
  {32'h405643f3, 32'hc0277320} /* (7, 15, 5) {real, imag} */,
  {32'h402f0d29, 32'hbf8336d6} /* (7, 15, 4) {real, imag} */,
  {32'hbf7a6579, 32'hc00beaf8} /* (7, 15, 3) {real, imag} */,
  {32'hc0303c75, 32'hc0b32b58} /* (7, 15, 2) {real, imag} */,
  {32'hbeaa278a, 32'hc010da18} /* (7, 15, 1) {real, imag} */,
  {32'h3ec5e118, 32'hbf874781} /* (7, 15, 0) {real, imag} */,
  {32'hbfbd69bc, 32'h3fc3efde} /* (7, 14, 15) {real, imag} */,
  {32'hc01dd31e, 32'h407fa064} /* (7, 14, 14) {real, imag} */,
  {32'hbfb980a4, 32'h3e8cf577} /* (7, 14, 13) {real, imag} */,
  {32'h3f9ec25e, 32'hbf4d3e7e} /* (7, 14, 12) {real, imag} */,
  {32'h3fd9ba87, 32'h3f286b43} /* (7, 14, 11) {real, imag} */,
  {32'h400f54e7, 32'hbf75d0d5} /* (7, 14, 10) {real, imag} */,
  {32'h3fe70780, 32'hc09172a6} /* (7, 14, 9) {real, imag} */,
  {32'h3f9cf76b, 32'hc0a26a6a} /* (7, 14, 8) {real, imag} */,
  {32'h3ffb1c51, 32'hbe13cac4} /* (7, 14, 7) {real, imag} */,
  {32'h3ffbc2f6, 32'hbf2e94c8} /* (7, 14, 6) {real, imag} */,
  {32'hc02525f8, 32'h3d735160} /* (7, 14, 5) {real, imag} */,
  {32'hbf944250, 32'h3f4da564} /* (7, 14, 4) {real, imag} */,
  {32'h4024a473, 32'h3efe04b8} /* (7, 14, 3) {real, imag} */,
  {32'h405ebc5c, 32'hbf4b9e20} /* (7, 14, 2) {real, imag} */,
  {32'hbcc94c00, 32'hbf8be0b5} /* (7, 14, 1) {real, imag} */,
  {32'hbe5d2517, 32'h3dad5cc8} /* (7, 14, 0) {real, imag} */,
  {32'hbf61add5, 32'h3fc84bfd} /* (7, 13, 15) {real, imag} */,
  {32'hc0164560, 32'h3ffb73a2} /* (7, 13, 14) {real, imag} */,
  {32'hbfd7f350, 32'h3ff2e4d1} /* (7, 13, 13) {real, imag} */,
  {32'hbf062050, 32'hbfa65811} /* (7, 13, 12) {real, imag} */,
  {32'hbd5fccb0, 32'hbfba9862} /* (7, 13, 11) {real, imag} */,
  {32'h3f23d072, 32'h40325c10} /* (7, 13, 10) {real, imag} */,
  {32'h3e88a4ca, 32'h3ff0a2f5} /* (7, 13, 9) {real, imag} */,
  {32'h3eedf672, 32'h3f90120e} /* (7, 13, 8) {real, imag} */,
  {32'hbd320210, 32'h3f693403} /* (7, 13, 7) {real, imag} */,
  {32'hbf1a27fd, 32'h3e252980} /* (7, 13, 6) {real, imag} */,
  {32'hc008905a, 32'hbfc592ba} /* (7, 13, 5) {real, imag} */,
  {32'hba568b00, 32'hbf32d565} /* (7, 13, 4) {real, imag} */,
  {32'h3f4bb5fb, 32'hbf997e88} /* (7, 13, 3) {real, imag} */,
  {32'h3e869fc4, 32'hbed2c2a4} /* (7, 13, 2) {real, imag} */,
  {32'hbf91e974, 32'h3ffb3c74} /* (7, 13, 1) {real, imag} */,
  {32'hbed7d5e2, 32'h3f83d5ea} /* (7, 13, 0) {real, imag} */,
  {32'h3f0a89b6, 32'hbf3defdc} /* (7, 12, 15) {real, imag} */,
  {32'hbef18bb4, 32'hbf3b741a} /* (7, 12, 14) {real, imag} */,
  {32'hbf721a40, 32'hbf81b6b6} /* (7, 12, 13) {real, imag} */,
  {32'h3fbe5876, 32'hbe525dd8} /* (7, 12, 12) {real, imag} */,
  {32'h4007a2f2, 32'h3f5b20b8} /* (7, 12, 11) {real, imag} */,
  {32'hbf465c47, 32'h4043a6e8} /* (7, 12, 10) {real, imag} */,
  {32'hbfa54bae, 32'h40658e12} /* (7, 12, 9) {real, imag} */,
  {32'hbff7243c, 32'h3fe3040a} /* (7, 12, 8) {real, imag} */,
  {32'hc00727a8, 32'h3e6b686c} /* (7, 12, 7) {real, imag} */,
  {32'hbf8b815c, 32'hbe806842} /* (7, 12, 6) {real, imag} */,
  {32'hc00d7b3c, 32'hbd785b40} /* (7, 12, 5) {real, imag} */,
  {32'hbfa065dc, 32'h3fa5afcc} /* (7, 12, 4) {real, imag} */,
  {32'h3fdb840c, 32'hbf4fce16} /* (7, 12, 3) {real, imag} */,
  {32'h3fcd71da, 32'hc0241046} /* (7, 12, 2) {real, imag} */,
  {32'h3f699e63, 32'hbf8a0fc3} /* (7, 12, 1) {real, imag} */,
  {32'h40117979, 32'hbeec887e} /* (7, 12, 0) {real, imag} */,
  {32'hbfc74586, 32'hbf6b6fbe} /* (7, 11, 15) {real, imag} */,
  {32'hbfe99a71, 32'hbfdae71c} /* (7, 11, 14) {real, imag} */,
  {32'h3eae6370, 32'hbfda0068} /* (7, 11, 13) {real, imag} */,
  {32'h3f843590, 32'hbf97a258} /* (7, 11, 12) {real, imag} */,
  {32'h3face730, 32'hbe349ad0} /* (7, 11, 11) {real, imag} */,
  {32'h3ee4ec3a, 32'h3e503000} /* (7, 11, 10) {real, imag} */,
  {32'h3fe8289c, 32'h3fd7e2c1} /* (7, 11, 9) {real, imag} */,
  {32'h4019d62d, 32'h3fd8da3b} /* (7, 11, 8) {real, imag} */,
  {32'h3ec97028, 32'h3ff9ae90} /* (7, 11, 7) {real, imag} */,
  {32'hbef1535b, 32'h3f49e2a5} /* (7, 11, 6) {real, imag} */,
  {32'hbf27ad16, 32'hbf11c5cc} /* (7, 11, 5) {real, imag} */,
  {32'hbee8cb26, 32'h3cb26558} /* (7, 11, 4) {real, imag} */,
  {32'hbf1f05a6, 32'h3cabfe30} /* (7, 11, 3) {real, imag} */,
  {32'hbeb43766, 32'hbea15504} /* (7, 11, 2) {real, imag} */,
  {32'hbf2bf545, 32'hc01f7605} /* (7, 11, 1) {real, imag} */,
  {32'hbf9ba75e, 32'hbf7acd11} /* (7, 11, 0) {real, imag} */,
  {32'hbe920b21, 32'hbe332b5d} /* (7, 10, 15) {real, imag} */,
  {32'h3d824460, 32'hbf309217} /* (7, 10, 14) {real, imag} */,
  {32'hbf0dc7c6, 32'hbeacaa72} /* (7, 10, 13) {real, imag} */,
  {32'h3eb11900, 32'hbf48b992} /* (7, 10, 12) {real, imag} */,
  {32'h3f62253c, 32'hbf5bece2} /* (7, 10, 11) {real, imag} */,
  {32'h3d5e3640, 32'hbf6448af} /* (7, 10, 10) {real, imag} */,
  {32'hbf40a1ce, 32'hbfae68ca} /* (7, 10, 9) {real, imag} */,
  {32'hbdab1d74, 32'hbfe083de} /* (7, 10, 8) {real, imag} */,
  {32'h3e0466a2, 32'hbd807ec2} /* (7, 10, 7) {real, imag} */,
  {32'hbf29afa9, 32'h3e693026} /* (7, 10, 6) {real, imag} */,
  {32'hbf5387d2, 32'h3ee034bf} /* (7, 10, 5) {real, imag} */,
  {32'h3e9cf016, 32'hbf9e94d2} /* (7, 10, 4) {real, imag} */,
  {32'h3f1bca55, 32'hbee04622} /* (7, 10, 3) {real, imag} */,
  {32'h3f8bb0fe, 32'h3ee2e8bf} /* (7, 10, 2) {real, imag} */,
  {32'h3fc73f58, 32'hbee5f33e} /* (7, 10, 1) {real, imag} */,
  {32'h3f5fd03a, 32'h3ea57296} /* (7, 10, 0) {real, imag} */,
  {32'h3f0f2def, 32'hbec4f856} /* (7, 9, 15) {real, imag} */,
  {32'h3eae4998, 32'hbf21ecba} /* (7, 9, 14) {real, imag} */,
  {32'hbeec9c1c, 32'hbf472820} /* (7, 9, 13) {real, imag} */,
  {32'hbf39a926, 32'hbe8aacb0} /* (7, 9, 12) {real, imag} */,
  {32'hbef7f408, 32'h3ea65fe8} /* (7, 9, 11) {real, imag} */,
  {32'hbdd085d0, 32'h3f315a13} /* (7, 9, 10) {real, imag} */,
  {32'hbf175854, 32'h3ea3d5fc} /* (7, 9, 9) {real, imag} */,
  {32'hbebc1e4a, 32'h3ee028a2} /* (7, 9, 8) {real, imag} */,
  {32'hbebfeca7, 32'h3f2427df} /* (7, 9, 7) {real, imag} */,
  {32'hbe00da22, 32'h3e586dde} /* (7, 9, 6) {real, imag} */,
  {32'hbf2abb95, 32'h3d8d5764} /* (7, 9, 5) {real, imag} */,
  {32'hbfd1b82f, 32'h3e504c60} /* (7, 9, 4) {real, imag} */,
  {32'hbf39dccb, 32'h3f0b7a03} /* (7, 9, 3) {real, imag} */,
  {32'h3f332a8e, 32'h3e2cfa78} /* (7, 9, 2) {real, imag} */,
  {32'h3f806ea0, 32'hbe5cece0} /* (7, 9, 1) {real, imag} */,
  {32'h3e968884, 32'h3d86ddee} /* (7, 9, 0) {real, imag} */,
  {32'h3f23e2d0, 32'h3e061658} /* (7, 8, 15) {real, imag} */,
  {32'h3c9ff340, 32'hbe3574d4} /* (7, 8, 14) {real, imag} */,
  {32'hbe8111d4, 32'hbe0f1e68} /* (7, 8, 13) {real, imag} */,
  {32'h3e86a750, 32'h3e7f3bf8} /* (7, 8, 12) {real, imag} */,
  {32'hbe0d6288, 32'h3f10f956} /* (7, 8, 11) {real, imag} */,
  {32'h3e532750, 32'h3f2f7550} /* (7, 8, 10) {real, imag} */,
  {32'h3e8817fe, 32'h3e552196} /* (7, 8, 9) {real, imag} */,
  {32'h3d93a010, 32'hbf8129f2} /* (7, 8, 8) {real, imag} */,
  {32'hbe02f75b, 32'hbecbd900} /* (7, 8, 7) {real, imag} */,
  {32'hbf184d44, 32'h3f2e2536} /* (7, 8, 6) {real, imag} */,
  {32'hbe9e0408, 32'hbed5debe} /* (7, 8, 5) {real, imag} */,
  {32'hbe2719f4, 32'hbfb1dea2} /* (7, 8, 4) {real, imag} */,
  {32'hbd2257e8, 32'hbebc314c} /* (7, 8, 3) {real, imag} */,
  {32'h3dad1708, 32'hbe5bbcb0} /* (7, 8, 2) {real, imag} */,
  {32'h3f46ffac, 32'hbe011270} /* (7, 8, 1) {real, imag} */,
  {32'h3f62b75a, 32'hbc48dc80} /* (7, 8, 0) {real, imag} */,
  {32'hbf0aa12b, 32'hbe3b4eec} /* (7, 7, 15) {real, imag} */,
  {32'hbfe59330, 32'hbf67f0b8} /* (7, 7, 14) {real, imag} */,
  {32'hbf15ebb0, 32'hbec42be8} /* (7, 7, 13) {real, imag} */,
  {32'h3f6bb75a, 32'h3f4bc32c} /* (7, 7, 12) {real, imag} */,
  {32'h3fd35190, 32'h3edd10f8} /* (7, 7, 11) {real, imag} */,
  {32'h3f822e25, 32'hbeb02c1a} /* (7, 7, 10) {real, imag} */,
  {32'h3f121c28, 32'hbd811310} /* (7, 7, 9) {real, imag} */,
  {32'h3f402337, 32'h3f89c6e2} /* (7, 7, 8) {real, imag} */,
  {32'hbf7834a0, 32'hbc9e9220} /* (7, 7, 7) {real, imag} */,
  {32'hbe677846, 32'h3eac8969} /* (7, 7, 6) {real, imag} */,
  {32'h3fb714bc, 32'h3e09a252} /* (7, 7, 5) {real, imag} */,
  {32'h3f5dd9a6, 32'h3ec37be0} /* (7, 7, 4) {real, imag} */,
  {32'h3f3fdab5, 32'h3f3cd797} /* (7, 7, 3) {real, imag} */,
  {32'h3f12a42e, 32'h3edc406c} /* (7, 7, 2) {real, imag} */,
  {32'hbd9bdc78, 32'h3f0bcde4} /* (7, 7, 1) {real, imag} */,
  {32'hbdee7a11, 32'hbe038169} /* (7, 7, 0) {real, imag} */,
  {32'hbd42f718, 32'hbee2a8fa} /* (7, 6, 15) {real, imag} */,
  {32'hbc152600, 32'hbf2f8609} /* (7, 6, 14) {real, imag} */,
  {32'h3de7b630, 32'hbe90f100} /* (7, 6, 13) {real, imag} */,
  {32'hbfeec062, 32'hbf63123a} /* (7, 6, 12) {real, imag} */,
  {32'hbfe1bbba, 32'hbfee0f3f} /* (7, 6, 11) {real, imag} */,
  {32'h3f45ce3a, 32'hbe52728c} /* (7, 6, 10) {real, imag} */,
  {32'h3f998613, 32'hbefd5e56} /* (7, 6, 9) {real, imag} */,
  {32'h3f501c92, 32'hbe86ab1e} /* (7, 6, 8) {real, imag} */,
  {32'h3e31f7d2, 32'h3ec47dec} /* (7, 6, 7) {real, imag} */,
  {32'hbec95786, 32'hbec409c1} /* (7, 6, 6) {real, imag} */,
  {32'hbf129f02, 32'hbe301192} /* (7, 6, 5) {real, imag} */,
  {32'hbf0473a9, 32'hbeaf9ce8} /* (7, 6, 4) {real, imag} */,
  {32'h3f7ddae3, 32'hbfa69e8e} /* (7, 6, 3) {real, imag} */,
  {32'h40088ac6, 32'h3ee0eae9} /* (7, 6, 2) {real, imag} */,
  {32'h3f070217, 32'hbf83eaec} /* (7, 6, 1) {real, imag} */,
  {32'hbd9f22c4, 32'hbfb33eae} /* (7, 6, 0) {real, imag} */,
  {32'hbf130d5f, 32'hbf96336f} /* (7, 5, 15) {real, imag} */,
  {32'h3f2a9792, 32'hbf6e4bb7} /* (7, 5, 14) {real, imag} */,
  {32'h3fb56eb3, 32'hbe8e7008} /* (7, 5, 13) {real, imag} */,
  {32'h3cc23380, 32'h3f146e60} /* (7, 5, 12) {real, imag} */,
  {32'hc002e026, 32'hbf884766} /* (7, 5, 11) {real, imag} */,
  {32'hc01b1321, 32'hbfcd08c8} /* (7, 5, 10) {real, imag} */,
  {32'hbeb4b670, 32'hbefb7ec4} /* (7, 5, 9) {real, imag} */,
  {32'hbff84c8b, 32'h3f8a0749} /* (7, 5, 8) {real, imag} */,
  {32'hbfcdc48e, 32'h3fabfec2} /* (7, 5, 7) {real, imag} */,
  {32'hbf49b6f6, 32'hbef58312} /* (7, 5, 6) {real, imag} */,
  {32'hbf8b0bd5, 32'hbf2e11b4} /* (7, 5, 5) {real, imag} */,
  {32'hbf9eb9a0, 32'hbda6f5ba} /* (7, 5, 4) {real, imag} */,
  {32'hbf813078, 32'h3f42140e} /* (7, 5, 3) {real, imag} */,
  {32'hbfbe420a, 32'h3f28234c} /* (7, 5, 2) {real, imag} */,
  {32'hbf9588d4, 32'hbeb3f338} /* (7, 5, 1) {real, imag} */,
  {32'hb9e6f800, 32'hbea66392} /* (7, 5, 0) {real, imag} */,
  {32'hbf0de03e, 32'hbe112c32} /* (7, 4, 15) {real, imag} */,
  {32'hbfc02f27, 32'hc0060cb0} /* (7, 4, 14) {real, imag} */,
  {32'hc02d9a80, 32'hbfb3a36a} /* (7, 4, 13) {real, imag} */,
  {32'hbfcb902c, 32'hbd7bc520} /* (7, 4, 12) {real, imag} */,
  {32'hbe8da824, 32'h3ede6087} /* (7, 4, 11) {real, imag} */,
  {32'h3f10dcad, 32'h3d2e7ba0} /* (7, 4, 10) {real, imag} */,
  {32'h3f998bae, 32'h3daedc40} /* (7, 4, 9) {real, imag} */,
  {32'h402df69e, 32'hbe364794} /* (7, 4, 8) {real, imag} */,
  {32'h402e0efc, 32'hbf542d0b} /* (7, 4, 7) {real, imag} */,
  {32'h40065f58, 32'h3f114b1d} /* (7, 4, 6) {real, imag} */,
  {32'h3fbc32ad, 32'h405417c1} /* (7, 4, 5) {real, imag} */,
  {32'h3fe5d8f0, 32'h3fdc0bec} /* (7, 4, 4) {real, imag} */,
  {32'h3f927f6e, 32'hbeacccd3} /* (7, 4, 3) {real, imag} */,
  {32'h3e092fd4, 32'hbe8b3bd0} /* (7, 4, 2) {real, imag} */,
  {32'hbfacedf6, 32'hbf882df1} /* (7, 4, 1) {real, imag} */,
  {32'hbfb226c8, 32'hbfa4ce18} /* (7, 4, 0) {real, imag} */,
  {32'hbf825468, 32'h3eeb30b4} /* (7, 3, 15) {real, imag} */,
  {32'hc03d75ee, 32'h3f7d20fb} /* (7, 3, 14) {real, imag} */,
  {32'hc01b91aa, 32'hbe155188} /* (7, 3, 13) {real, imag} */,
  {32'h3f26bc74, 32'hc01ef07e} /* (7, 3, 12) {real, imag} */,
  {32'h3f89c6f4, 32'hbfe3f676} /* (7, 3, 11) {real, imag} */,
  {32'hbef7c688, 32'h3cf81800} /* (7, 3, 10) {real, imag} */,
  {32'hbe5a60b4, 32'h3f85b907} /* (7, 3, 9) {real, imag} */,
  {32'hbf2b097d, 32'h3f7f8fd4} /* (7, 3, 8) {real, imag} */,
  {32'h3fa54be8, 32'h3f86490c} /* (7, 3, 7) {real, imag} */,
  {32'h3e5fd120, 32'h407b4800} /* (7, 3, 6) {real, imag} */,
  {32'hc007952a, 32'h40762267} /* (7, 3, 5) {real, imag} */,
  {32'hbdba3562, 32'h3f8d9e26} /* (7, 3, 4) {real, imag} */,
  {32'hbfc4dee6, 32'h3f26c3ac} /* (7, 3, 3) {real, imag} */,
  {32'hbe113408, 32'h3f88c6c8} /* (7, 3, 2) {real, imag} */,
  {32'h3e51d2f4, 32'h3fc1bbb0} /* (7, 3, 1) {real, imag} */,
  {32'hbf226abb, 32'h3e0ae334} /* (7, 3, 0) {real, imag} */,
  {32'hbf5eefe0, 32'h4013f678} /* (7, 2, 15) {real, imag} */,
  {32'h3e7e2428, 32'h4012d856} /* (7, 2, 14) {real, imag} */,
  {32'hbf71a474, 32'hbf79c6e4} /* (7, 2, 13) {real, imag} */,
  {32'hbfe25038, 32'hbf5ac1d6} /* (7, 2, 12) {real, imag} */,
  {32'hbf0943ea, 32'hc021989c} /* (7, 2, 11) {real, imag} */,
  {32'hbfc8c712, 32'hbffaebce} /* (7, 2, 10) {real, imag} */,
  {32'hc030a9f0, 32'h4015b16b} /* (7, 2, 9) {real, imag} */,
  {32'hbf5ede62, 32'h3ec4e848} /* (7, 2, 8) {real, imag} */,
  {32'hbf95be27, 32'h3f4b8029} /* (7, 2, 7) {real, imag} */,
  {32'h3f428da1, 32'h403362f4} /* (7, 2, 6) {real, imag} */,
  {32'h3fff8d05, 32'h400aa3ae} /* (7, 2, 5) {real, imag} */,
  {32'h3fd802d4, 32'hbf9c9586} /* (7, 2, 4) {real, imag} */,
  {32'h40052f91, 32'h3eb97316} /* (7, 2, 3) {real, imag} */,
  {32'hbf19ebc2, 32'h3e814f18} /* (7, 2, 2) {real, imag} */,
  {32'hbfaca183, 32'hbfb105b9} /* (7, 2, 1) {real, imag} */,
  {32'hbd1ce38c, 32'hbf9ace24} /* (7, 2, 0) {real, imag} */,
  {32'h4024cb65, 32'hc04e41a6} /* (7, 1, 15) {real, imag} */,
  {32'h3fcdc566, 32'hbfda6c6f} /* (7, 1, 14) {real, imag} */,
  {32'h3f6bae73, 32'hbf1845c5} /* (7, 1, 13) {real, imag} */,
  {32'h4011a9c2, 32'hc0652e3a} /* (7, 1, 12) {real, imag} */,
  {32'hbf7d8ac4, 32'hc06e1e8a} /* (7, 1, 11) {real, imag} */,
  {32'hc00b8778, 32'hbf3e3e28} /* (7, 1, 10) {real, imag} */,
  {32'hbf6f5db2, 32'hc01b9c62} /* (7, 1, 9) {real, imag} */,
  {32'hbeb240f8, 32'hbf6c0a2c} /* (7, 1, 8) {real, imag} */,
  {32'h3e8ddf3c, 32'h3fa7aeb0} /* (7, 1, 7) {real, imag} */,
  {32'hbfa3b2a6, 32'hbfd81d77} /* (7, 1, 6) {real, imag} */,
  {32'hc09b7350, 32'h3f065a5e} /* (7, 1, 5) {real, imag} */,
  {32'hc0029a93, 32'h4035f223} /* (7, 1, 4) {real, imag} */,
  {32'h400b2e22, 32'h3dd9c610} /* (7, 1, 3) {real, imag} */,
  {32'h4037780b, 32'hbe66e150} /* (7, 1, 2) {real, imag} */,
  {32'hbf7f0b2d, 32'h3eafafbc} /* (7, 1, 1) {real, imag} */,
  {32'hbf1444c0, 32'h3fcdcd9b} /* (7, 1, 0) {real, imag} */,
  {32'h3f627bc8, 32'h403143d4} /* (7, 0, 15) {real, imag} */,
  {32'h403e19c2, 32'h3f77da87} /* (7, 0, 14) {real, imag} */,
  {32'hbea57b0c, 32'h3faa8875} /* (7, 0, 13) {real, imag} */,
  {32'hc0178427, 32'h3fe29bcd} /* (7, 0, 12) {real, imag} */,
  {32'h3fbf4b11, 32'hc05f6944} /* (7, 0, 11) {real, imag} */,
  {32'hbf102a08, 32'hc094925c} /* (7, 0, 10) {real, imag} */,
  {32'h3ed9c042, 32'hbf08fdd6} /* (7, 0, 9) {real, imag} */,
  {32'hbfd5e124, 32'hbdf64118} /* (7, 0, 8) {real, imag} */,
  {32'hbed2bdc4, 32'h4085ca5c} /* (7, 0, 7) {real, imag} */,
  {32'h3e0401f8, 32'h4038ba4c} /* (7, 0, 6) {real, imag} */,
  {32'h404a136d, 32'h3ec4325a} /* (7, 0, 5) {real, imag} */,
  {32'h3fdfc706, 32'h3f57c6f5} /* (7, 0, 4) {real, imag} */,
  {32'hbf04face, 32'h405e7b80} /* (7, 0, 3) {real, imag} */,
  {32'hbfee4b68, 32'h4063accb} /* (7, 0, 2) {real, imag} */,
  {32'h3f59f37e, 32'h40759c31} /* (7, 0, 1) {real, imag} */,
  {32'h3f0f64dc, 32'h400a9870} /* (7, 0, 0) {real, imag} */,
  {32'hc003b74c, 32'h4008b047} /* (6, 15, 15) {real, imag} */,
  {32'hbee40baa, 32'h3cfef680} /* (6, 15, 14) {real, imag} */,
  {32'hbde4fda0, 32'hc0423440} /* (6, 15, 13) {real, imag} */,
  {32'hc02ebff6, 32'hc0248996} /* (6, 15, 12) {real, imag} */,
  {32'hc05a1b96, 32'hc03612fa} /* (6, 15, 11) {real, imag} */,
  {32'hc0b91eea, 32'hbf98a174} /* (6, 15, 10) {real, imag} */,
  {32'hbfb22d1a, 32'h3f3f1fec} /* (6, 15, 9) {real, imag} */,
  {32'hc037defa, 32'h407d65a5} /* (6, 15, 8) {real, imag} */,
  {32'h3e09e4d6, 32'h40bb418a} /* (6, 15, 7) {real, imag} */,
  {32'hbf9d603b, 32'h40a479a5} /* (6, 15, 6) {real, imag} */,
  {32'hc0910808, 32'h40230114} /* (6, 15, 5) {real, imag} */,
  {32'hc0c69464, 32'hc00f0439} /* (6, 15, 4) {real, imag} */,
  {32'hc04261dc, 32'h3dc33ff8} /* (6, 15, 3) {real, imag} */,
  {32'h3ffc26a5, 32'h3e98abd8} /* (6, 15, 2) {real, imag} */,
  {32'hbf4498a8, 32'h409703e4} /* (6, 15, 1) {real, imag} */,
  {32'h3f16f80c, 32'h404a54bc} /* (6, 15, 0) {real, imag} */,
  {32'h3f82baca, 32'hbfe84ee2} /* (6, 14, 15) {real, imag} */,
  {32'h403ca726, 32'hbec30fc8} /* (6, 14, 14) {real, imag} */,
  {32'h3eb08f04, 32'h3fe7803a} /* (6, 14, 13) {real, imag} */,
  {32'h40260565, 32'hbe9fd630} /* (6, 14, 12) {real, imag} */,
  {32'hbfeda528, 32'hbf446248} /* (6, 14, 11) {real, imag} */,
  {32'hc0273c10, 32'hbfe9067c} /* (6, 14, 10) {real, imag} */,
  {32'hbf2d85f6, 32'hbe498002} /* (6, 14, 9) {real, imag} */,
  {32'h3f855a19, 32'hc0166b60} /* (6, 14, 8) {real, imag} */,
  {32'hc0133575, 32'h3f19c8ba} /* (6, 14, 7) {real, imag} */,
  {32'h3fab64f6, 32'h3f9a4ff9} /* (6, 14, 6) {real, imag} */,
  {32'h40631aec, 32'h3e0d9c20} /* (6, 14, 5) {real, imag} */,
  {32'h4058bbd2, 32'h40734bc3} /* (6, 14, 4) {real, imag} */,
  {32'hc01992d9, 32'h40297e8d} /* (6, 14, 3) {real, imag} */,
  {32'hc013976c, 32'h403477dc} /* (6, 14, 2) {real, imag} */,
  {32'h3f96d78a, 32'h40259b27} /* (6, 14, 1) {real, imag} */,
  {32'h3ed3b273, 32'hbe9ca41c} /* (6, 14, 0) {real, imag} */,
  {32'hc01fecf8, 32'hc0185a3a} /* (6, 13, 15) {real, imag} */,
  {32'hbf9a9c74, 32'hc08abc55} /* (6, 13, 14) {real, imag} */,
  {32'h3fc9f8e5, 32'hc05b9654} /* (6, 13, 13) {real, imag} */,
  {32'hbfc1975c, 32'h3f68c676} /* (6, 13, 12) {real, imag} */,
  {32'hc031c844, 32'h3ff91a45} /* (6, 13, 11) {real, imag} */,
  {32'h3e5ea308, 32'h3fa6fc00} /* (6, 13, 10) {real, imag} */,
  {32'hbf87e5b2, 32'h3f5c51e5} /* (6, 13, 9) {real, imag} */,
  {32'hc07640cb, 32'hc07fc688} /* (6, 13, 8) {real, imag} */,
  {32'hc0838eeb, 32'hc0220182} /* (6, 13, 7) {real, imag} */,
  {32'hc01a6174, 32'h3f5987a2} /* (6, 13, 6) {real, imag} */,
  {32'hc06db010, 32'hbf3be70d} /* (6, 13, 5) {real, imag} */,
  {32'hc068c8ad, 32'hc0413be7} /* (6, 13, 4) {real, imag} */,
  {32'hbe99d37c, 32'hc04cdcc7} /* (6, 13, 3) {real, imag} */,
  {32'h3f9c86d4, 32'h3f382840} /* (6, 13, 2) {real, imag} */,
  {32'h4089c815, 32'hbf1e180a} /* (6, 13, 1) {real, imag} */,
  {32'h402ec1ac, 32'hbfdea1a4} /* (6, 13, 0) {real, imag} */,
  {32'hc0158808, 32'h3f34eb6b} /* (6, 12, 15) {real, imag} */,
  {32'h3f8d0ce2, 32'h4046b992} /* (6, 12, 14) {real, imag} */,
  {32'h406357fd, 32'h4029d438} /* (6, 12, 13) {real, imag} */,
  {32'h3f1c2a98, 32'h3cfe3a20} /* (6, 12, 12) {real, imag} */,
  {32'hbfcb9238, 32'h3e9630cc} /* (6, 12, 11) {real, imag} */,
  {32'h3f46e9eb, 32'h40555f88} /* (6, 12, 10) {real, imag} */,
  {32'h3f6d2aa6, 32'h40d792c1} /* (6, 12, 9) {real, imag} */,
  {32'h409c51f2, 32'h3f89ad08} /* (6, 12, 8) {real, imag} */,
  {32'h4094b581, 32'h3fb1c38c} /* (6, 12, 7) {real, imag} */,
  {32'hbdf24998, 32'h4000c920} /* (6, 12, 6) {real, imag} */,
  {32'hbfc8ff72, 32'hbfa1b93f} /* (6, 12, 5) {real, imag} */,
  {32'h3fd8a530, 32'hbfae2138} /* (6, 12, 4) {real, imag} */,
  {32'h3d50fd90, 32'hbe5008b0} /* (6, 12, 3) {real, imag} */,
  {32'hbf1b82c3, 32'h3f2ce2cf} /* (6, 12, 2) {real, imag} */,
  {32'hbf9df56f, 32'hbf84501b} /* (6, 12, 1) {real, imag} */,
  {32'hbfe85f40, 32'hbfa7e216} /* (6, 12, 0) {real, imag} */,
  {32'hbf9ba958, 32'h3f8379de} /* (6, 11, 15) {real, imag} */,
  {32'h3d92c050, 32'h3e6d8b9c} /* (6, 11, 14) {real, imag} */,
  {32'h401c983d, 32'hbe7ec800} /* (6, 11, 13) {real, imag} */,
  {32'h3f9bb01c, 32'hbdf791b0} /* (6, 11, 12) {real, imag} */,
  {32'hc04078fb, 32'hbdfa5b30} /* (6, 11, 11) {real, imag} */,
  {32'hbf5a492f, 32'h4031de44} /* (6, 11, 10) {real, imag} */,
  {32'h3f546f4e, 32'h3fc4e3bb} /* (6, 11, 9) {real, imag} */,
  {32'h3f3542f4, 32'h3efafa7c} /* (6, 11, 8) {real, imag} */,
  {32'h3fb6fe0b, 32'hbf951bc6} /* (6, 11, 7) {real, imag} */,
  {32'h3e098bcc, 32'h3ffa3e7b} /* (6, 11, 6) {real, imag} */,
  {32'h400c93b2, 32'h3f3432ad} /* (6, 11, 5) {real, imag} */,
  {32'h3fb4878a, 32'hbf59b677} /* (6, 11, 4) {real, imag} */,
  {32'h3f9eece5, 32'h3edc26dc} /* (6, 11, 3) {real, imag} */,
  {32'h40052279, 32'hbf03a1ab} /* (6, 11, 2) {real, imag} */,
  {32'h3fb4dcba, 32'h3e849d20} /* (6, 11, 1) {real, imag} */,
  {32'hbf911ad2, 32'h3f804d2e} /* (6, 11, 0) {real, imag} */,
  {32'hbf82f66a, 32'h3ea401f4} /* (6, 10, 15) {real, imag} */,
  {32'hbfd3e86a, 32'hbeff7408} /* (6, 10, 14) {real, imag} */,
  {32'h3f470da3, 32'h3cacbe80} /* (6, 10, 13) {real, imag} */,
  {32'h3fdbe5d6, 32'h40117f3a} /* (6, 10, 12) {real, imag} */,
  {32'h401fae78, 32'h3fcf6277} /* (6, 10, 11) {real, imag} */,
  {32'hbffed3f7, 32'h3f2d31ea} /* (6, 10, 10) {real, imag} */,
  {32'hbff15324, 32'hbfcce56c} /* (6, 10, 9) {real, imag} */,
  {32'h3ef30db1, 32'h3ec7b0ee} /* (6, 10, 8) {real, imag} */,
  {32'hbed63910, 32'h3cf2d0a0} /* (6, 10, 7) {real, imag} */,
  {32'hbf8c793b, 32'hbf91f559} /* (6, 10, 6) {real, imag} */,
  {32'h3f8f8b03, 32'hbfe246c1} /* (6, 10, 5) {real, imag} */,
  {32'h3f796e9c, 32'hbfea8fdd} /* (6, 10, 4) {real, imag} */,
  {32'h3e26fcc0, 32'h3f39533f} /* (6, 10, 3) {real, imag} */,
  {32'h3ee05059, 32'hbde43598} /* (6, 10, 2) {real, imag} */,
  {32'hbf6d3e99, 32'hbfb2152c} /* (6, 10, 1) {real, imag} */,
  {32'hbf448f38, 32'hbe24ccb4} /* (6, 10, 0) {real, imag} */,
  {32'h3f179c2b, 32'hbe84c5ef} /* (6, 9, 15) {real, imag} */,
  {32'h3ef17fe3, 32'hbd9fa2d0} /* (6, 9, 14) {real, imag} */,
  {32'hbec079ec, 32'h3f9d65ee} /* (6, 9, 13) {real, imag} */,
  {32'h3e286e68, 32'h3f8419e0} /* (6, 9, 12) {real, imag} */,
  {32'h3f8d73c5, 32'hbe9ffbec} /* (6, 9, 11) {real, imag} */,
  {32'h3f62e3e6, 32'hbfd2a39e} /* (6, 9, 10) {real, imag} */,
  {32'h3f84ac32, 32'hbf8a3282} /* (6, 9, 9) {real, imag} */,
  {32'h3f80f110, 32'h3de0c6d8} /* (6, 9, 8) {real, imag} */,
  {32'hbe19eb1c, 32'h3e9f2510} /* (6, 9, 7) {real, imag} */,
  {32'hbef49353, 32'h3da1e4b8} /* (6, 9, 6) {real, imag} */,
  {32'hbf1bac32, 32'h3f568ed6} /* (6, 9, 5) {real, imag} */,
  {32'h3f7de196, 32'h3f318420} /* (6, 9, 4) {real, imag} */,
  {32'h3ff313aa, 32'h3fe390b2} /* (6, 9, 3) {real, imag} */,
  {32'h3d0826f0, 32'h3f817ae1} /* (6, 9, 2) {real, imag} */,
  {32'hbf774ff6, 32'hbe65869c} /* (6, 9, 1) {real, imag} */,
  {32'hbe93abfc, 32'hbb912780} /* (6, 9, 0) {real, imag} */,
  {32'h3d675080, 32'h3f4fb580} /* (6, 8, 15) {real, imag} */,
  {32'h3ee55084, 32'h3efa9b6c} /* (6, 8, 14) {real, imag} */,
  {32'h3f80c102, 32'hbf4ebd70} /* (6, 8, 13) {real, imag} */,
  {32'h3ef0946e, 32'hbf196eaa} /* (6, 8, 12) {real, imag} */,
  {32'h3f058902, 32'hbf938d00} /* (6, 8, 11) {real, imag} */,
  {32'hbe5a9488, 32'hbfaec572} /* (6, 8, 10) {real, imag} */,
  {32'hbf916d57, 32'h3f526de9} /* (6, 8, 9) {real, imag} */,
  {32'h3db55ea0, 32'h3f90ac16} /* (6, 8, 8) {real, imag} */,
  {32'h3f7a5c36, 32'h3f17f72a} /* (6, 8, 7) {real, imag} */,
  {32'h3dcc7200, 32'h3f3b7140} /* (6, 8, 6) {real, imag} */,
  {32'hbbd4f100, 32'h3f89b55a} /* (6, 8, 5) {real, imag} */,
  {32'hbecd0b6c, 32'h3e23fac8} /* (6, 8, 4) {real, imag} */,
  {32'h3e582ea0, 32'h3ee941e0} /* (6, 8, 3) {real, imag} */,
  {32'h3eaf8df8, 32'h3f365888} /* (6, 8, 2) {real, imag} */,
  {32'hbdf98084, 32'h3f0a89fc} /* (6, 8, 1) {real, imag} */,
  {32'h3ee9c314, 32'h3f046df4} /* (6, 8, 0) {real, imag} */,
  {32'h3e8eef96, 32'h3f6492d8} /* (6, 7, 15) {real, imag} */,
  {32'h3f995a75, 32'h3fd7ff61} /* (6, 7, 14) {real, imag} */,
  {32'h3f2ba0de, 32'h3d9216a0} /* (6, 7, 13) {real, imag} */,
  {32'hbeae2eb4, 32'hbf8085ba} /* (6, 7, 12) {real, imag} */,
  {32'h3f53ebd2, 32'hbedef67c} /* (6, 7, 11) {real, imag} */,
  {32'h3fcd1bdf, 32'hbebadd8e} /* (6, 7, 10) {real, imag} */,
  {32'hbd8e9ba8, 32'h3f70be04} /* (6, 7, 9) {real, imag} */,
  {32'h3e7986d0, 32'h3f776dd3} /* (6, 7, 8) {real, imag} */,
  {32'h3f366be6, 32'hbea6bd60} /* (6, 7, 7) {real, imag} */,
  {32'h3f6cdf56, 32'hbf9ad172} /* (6, 7, 6) {real, imag} */,
  {32'h3eb4bb6c, 32'hbefcea7f} /* (6, 7, 5) {real, imag} */,
  {32'h3feb1127, 32'hbe439f58} /* (6, 7, 4) {real, imag} */,
  {32'h3e83b3e8, 32'h3f011add} /* (6, 7, 3) {real, imag} */,
  {32'hbf6475e1, 32'hbf59ee04} /* (6, 7, 2) {real, imag} */,
  {32'hbf350d0e, 32'hbfa30698} /* (6, 7, 1) {real, imag} */,
  {32'hbe1d8e57, 32'hbf691191} /* (6, 7, 0) {real, imag} */,
  {32'hbfc7143a, 32'hc003d72c} /* (6, 6, 15) {real, imag} */,
  {32'hbf97e032, 32'hc03b914f} /* (6, 6, 14) {real, imag} */,
  {32'hbf2b74e1, 32'hbfb70252} /* (6, 6, 13) {real, imag} */,
  {32'hbf9d03d2, 32'h3e181998} /* (6, 6, 12) {real, imag} */,
  {32'hbf25bbf4, 32'h3f151252} /* (6, 6, 11) {real, imag} */,
  {32'h3e8f0104, 32'hbe2fce78} /* (6, 6, 10) {real, imag} */,
  {32'hbe9b5026, 32'hbd81e5e8} /* (6, 6, 9) {real, imag} */,
  {32'h3d9eca24, 32'h3f355723} /* (6, 6, 8) {real, imag} */,
  {32'hbf56ecca, 32'h3eee03d4} /* (6, 6, 7) {real, imag} */,
  {32'hc0166320, 32'hbee7fd34} /* (6, 6, 6) {real, imag} */,
  {32'hbfa12597, 32'hbf689dde} /* (6, 6, 5) {real, imag} */,
  {32'hbf8131e6, 32'h3fd9e561} /* (6, 6, 4) {real, imag} */,
  {32'hbee3f13c, 32'h3fa4a15a} /* (6, 6, 3) {real, imag} */,
  {32'hbee222ef, 32'hbec953e2} /* (6, 6, 2) {real, imag} */,
  {32'hbf586c87, 32'hbf162d49} /* (6, 6, 1) {real, imag} */,
  {32'hbda5147c, 32'hbeaafd0a} /* (6, 6, 0) {real, imag} */,
  {32'h3fa5a416, 32'hbec82e12} /* (6, 5, 15) {real, imag} */,
  {32'hbf77803a, 32'hbfaf7ec2} /* (6, 5, 14) {real, imag} */,
  {32'hbecb3eb8, 32'h3fea0b3c} /* (6, 5, 13) {real, imag} */,
  {32'h3ffbf0fa, 32'h3fe760bb} /* (6, 5, 12) {real, imag} */,
  {32'h3fc46a6a, 32'h3fc64eeb} /* (6, 5, 11) {real, imag} */,
  {32'h3e8da59a, 32'h3fd2b27b} /* (6, 5, 10) {real, imag} */,
  {32'hc00b8900, 32'hc0248dd2} /* (6, 5, 9) {real, imag} */,
  {32'hbffb90ce, 32'hbfcffd0f} /* (6, 5, 8) {real, imag} */,
  {32'h3f2d6106, 32'h3ef7d882} /* (6, 5, 7) {real, imag} */,
  {32'h3fd64de6, 32'h4062334a} /* (6, 5, 6) {real, imag} */,
  {32'hbf7b2672, 32'h400d6e77} /* (6, 5, 5) {real, imag} */,
  {32'hc0318e01, 32'h40013846} /* (6, 5, 4) {real, imag} */,
  {32'h3f8512f1, 32'h4021ecfc} /* (6, 5, 3) {real, imag} */,
  {32'h4027dd6b, 32'h3fcc211c} /* (6, 5, 2) {real, imag} */,
  {32'h4014c91f, 32'hbdf89ea0} /* (6, 5, 1) {real, imag} */,
  {32'h3f0f5f4f, 32'hbd99bc18} /* (6, 5, 0) {real, imag} */,
  {32'h3fa192eb, 32'h3f38d151} /* (6, 4, 15) {real, imag} */,
  {32'h402c9c3e, 32'hbfb8224f} /* (6, 4, 14) {real, imag} */,
  {32'h40025ff9, 32'hc02090c0} /* (6, 4, 13) {real, imag} */,
  {32'h3e0aa746, 32'hbfeea880} /* (6, 4, 12) {real, imag} */,
  {32'hbf81c1b2, 32'h40682378} /* (6, 4, 11) {real, imag} */,
  {32'hbfa88216, 32'h3ffd68a4} /* (6, 4, 10) {real, imag} */,
  {32'hc024fcf4, 32'h40116d06} /* (6, 4, 9) {real, imag} */,
  {32'hc0211907, 32'h40378f80} /* (6, 4, 8) {real, imag} */,
  {32'hbfdf75c4, 32'h3ff33d52} /* (6, 4, 7) {real, imag} */,
  {32'hbfa57a0a, 32'hbf81972d} /* (6, 4, 6) {real, imag} */,
  {32'hc026de41, 32'hc0549ba2} /* (6, 4, 5) {real, imag} */,
  {32'hc02c02be, 32'hbf710aa8} /* (6, 4, 4) {real, imag} */,
  {32'hbfd2d634, 32'h403e6403} /* (6, 4, 3) {real, imag} */,
  {32'h3f29a9ef, 32'h3f317379} /* (6, 4, 2) {real, imag} */,
  {32'h3f65ffae, 32'h3fe97053} /* (6, 4, 1) {real, imag} */,
  {32'hbee34280, 32'h3e49a1a4} /* (6, 4, 0) {real, imag} */,
  {32'hbf01f94a, 32'hbf4336b2} /* (6, 3, 15) {real, imag} */,
  {32'hbfc0f2cc, 32'hc037a6b3} /* (6, 3, 14) {real, imag} */,
  {32'hbe2e51e0, 32'hc0a265fe} /* (6, 3, 13) {real, imag} */,
  {32'h3ffb75ce, 32'hc03e031a} /* (6, 3, 12) {real, imag} */,
  {32'hbf851e23, 32'hbf58f50a} /* (6, 3, 11) {real, imag} */,
  {32'hc02e5870, 32'h3f85b8d8} /* (6, 3, 10) {real, imag} */,
  {32'h3eb2acb6, 32'h3f24e147} /* (6, 3, 9) {real, imag} */,
  {32'h3faa74f2, 32'hbe7efca8} /* (6, 3, 8) {real, imag} */,
  {32'h400ca872, 32'hbf420d78} /* (6, 3, 7) {real, imag} */,
  {32'h3f75d247, 32'hbf870327} /* (6, 3, 6) {real, imag} */,
  {32'hbb6b6600, 32'h3fa80404} /* (6, 3, 5) {real, imag} */,
  {32'h3f3bf784, 32'hbe6e60f0} /* (6, 3, 4) {real, imag} */,
  {32'h3d1d03a4, 32'hc04268b9} /* (6, 3, 3) {real, imag} */,
  {32'hbf9231dc, 32'hc0741208} /* (6, 3, 2) {real, imag} */,
  {32'hbf15aaf0, 32'hc01ac7f8} /* (6, 3, 1) {real, imag} */,
  {32'hbb941100, 32'h3fa47e00} /* (6, 3, 0) {real, imag} */,
  {32'hc0131ac1, 32'h402befbb} /* (6, 2, 15) {real, imag} */,
  {32'hbf37fa38, 32'h40b6b888} /* (6, 2, 14) {real, imag} */,
  {32'h40565e8c, 32'h40a2aca6} /* (6, 2, 13) {real, imag} */,
  {32'h406e693b, 32'h409dd05b} /* (6, 2, 12) {real, imag} */,
  {32'h3fd8bbc2, 32'h409caa21} /* (6, 2, 11) {real, imag} */,
  {32'h403b9b5a, 32'h40cab301} /* (6, 2, 10) {real, imag} */,
  {32'h405fb9ce, 32'h3ef6785b} /* (6, 2, 9) {real, imag} */,
  {32'hbf1f3dae, 32'hbfc992ec} /* (6, 2, 8) {real, imag} */,
  {32'hbf128fcd, 32'h3f088bd2} /* (6, 2, 7) {real, imag} */,
  {32'h40c72056, 32'hc085c70d} /* (6, 2, 6) {real, imag} */,
  {32'h40ffd4aa, 32'hc0c25867} /* (6, 2, 5) {real, imag} */,
  {32'h40282f9c, 32'hc039c91d} /* (6, 2, 4) {real, imag} */,
  {32'hbf94da12, 32'hbf5412c5} /* (6, 2, 3) {real, imag} */,
  {32'h3f1f21ce, 32'h3ed665ec} /* (6, 2, 2) {real, imag} */,
  {32'h3f06dd17, 32'h4026d153} /* (6, 2, 1) {real, imag} */,
  {32'hbd264db8, 32'h40395a40} /* (6, 2, 0) {real, imag} */,
  {32'hbf844675, 32'hbfe3a66f} /* (6, 1, 15) {real, imag} */,
  {32'hbf0817c6, 32'hc0d294fa} /* (6, 1, 14) {real, imag} */,
  {32'h40a79e64, 32'hc0c97118} /* (6, 1, 13) {real, imag} */,
  {32'h406af226, 32'hbf2c3ab4} /* (6, 1, 12) {real, imag} */,
  {32'hbe80fd8c, 32'h408d4990} /* (6, 1, 11) {real, imag} */,
  {32'h3ece8988, 32'hbec560b6} /* (6, 1, 10) {real, imag} */,
  {32'h402f54ad, 32'hbff06d46} /* (6, 1, 9) {real, imag} */,
  {32'h400636da, 32'hc0810710} /* (6, 1, 8) {real, imag} */,
  {32'hbf7e1bba, 32'h3f2881e8} /* (6, 1, 7) {real, imag} */,
  {32'hbe0a6f58, 32'h4000db76} /* (6, 1, 6) {real, imag} */,
  {32'h40eae60c, 32'hbf9a7a4d} /* (6, 1, 5) {real, imag} */,
  {32'h40cea718, 32'h3f9feb22} /* (6, 1, 4) {real, imag} */,
  {32'h4087885e, 32'h3e89acc6} /* (6, 1, 3) {real, imag} */,
  {32'h400898e4, 32'hc041d103} /* (6, 1, 2) {real, imag} */,
  {32'h3e3e12d2, 32'h40550cf7} /* (6, 1, 1) {real, imag} */,
  {32'h3f486384, 32'h40b55152} /* (6, 1, 0) {real, imag} */,
  {32'h4010587e, 32'h3ed53338} /* (6, 0, 15) {real, imag} */,
  {32'h3fe5a165, 32'h405689dc} /* (6, 0, 14) {real, imag} */,
  {32'hbfabb546, 32'h40bffb68} /* (6, 0, 13) {real, imag} */,
  {32'hbfdc17bc, 32'h3f397662} /* (6, 0, 12) {real, imag} */,
  {32'h4003b11c, 32'hc022b245} /* (6, 0, 11) {real, imag} */,
  {32'h3fba2a88, 32'hbfbe872a} /* (6, 0, 10) {real, imag} */,
  {32'h3eeea20c, 32'h3e57c73c} /* (6, 0, 9) {real, imag} */,
  {32'h3f8439de, 32'h3f9bd93a} /* (6, 0, 8) {real, imag} */,
  {32'hbfbfb753, 32'h405d12fe} /* (6, 0, 7) {real, imag} */,
  {32'hc086a728, 32'h407a2bb6} /* (6, 0, 6) {real, imag} */,
  {32'hc001a514, 32'h409a3002} /* (6, 0, 5) {real, imag} */,
  {32'hbd8e5fce, 32'hbeacc868} /* (6, 0, 4) {real, imag} */,
  {32'h4024aaca, 32'hc050a070} /* (6, 0, 3) {real, imag} */,
  {32'h402ab9b1, 32'hc0239db8} /* (6, 0, 2) {real, imag} */,
  {32'h3f090148, 32'hc0869a8e} /* (6, 0, 1) {real, imag} */,
  {32'hbfbe46b4, 32'hc030c9e7} /* (6, 0, 0) {real, imag} */,
  {32'h40523aa4, 32'hc0790e4e} /* (5, 15, 15) {real, imag} */,
  {32'h403ec375, 32'hc050c411} /* (5, 15, 14) {real, imag} */,
  {32'h3f7691c8, 32'h3fc6fa45} /* (5, 15, 13) {real, imag} */,
  {32'hbe467cb8, 32'hc024358d} /* (5, 15, 12) {real, imag} */,
  {32'h40b0a71a, 32'hc01b0d2c} /* (5, 15, 11) {real, imag} */,
  {32'hbfa169fb, 32'h402b9220} /* (5, 15, 10) {real, imag} */,
  {32'hc082e0bb, 32'h3fb820e0} /* (5, 15, 9) {real, imag} */,
  {32'h405affba, 32'h3fd2b4ed} /* (5, 15, 8) {real, imag} */,
  {32'h3fb73058, 32'h3e645fb8} /* (5, 15, 7) {real, imag} */,
  {32'hc0a4e56b, 32'hc0ca6844} /* (5, 15, 6) {real, imag} */,
  {32'hbfd807d8, 32'hbd866b10} /* (5, 15, 5) {real, imag} */,
  {32'hbf06d226, 32'h40720f52} /* (5, 15, 4) {real, imag} */,
  {32'hbfd3b9c2, 32'hbd89f360} /* (5, 15, 3) {real, imag} */,
  {32'h3f6b82ca, 32'h3f84ee26} /* (5, 15, 2) {real, imag} */,
  {32'h402e257a, 32'h3d223b60} /* (5, 15, 1) {real, imag} */,
  {32'h40b9a2e4, 32'hbffb1ecc} /* (5, 15, 0) {real, imag} */,
  {32'h3e874c68, 32'hc0991a5d} /* (5, 14, 15) {real, imag} */,
  {32'h40849c74, 32'hbe5d6a90} /* (5, 14, 14) {real, imag} */,
  {32'h4092e323, 32'h3fec20bb} /* (5, 14, 13) {real, imag} */,
  {32'h408965ea, 32'hbef52427} /* (5, 14, 12) {real, imag} */,
  {32'hc0aad736, 32'h3e657918} /* (5, 14, 11) {real, imag} */,
  {32'hc01d4285, 32'hc047ff72} /* (5, 14, 10) {real, imag} */,
  {32'hc0145afe, 32'h40cc5fc4} /* (5, 14, 9) {real, imag} */,
  {32'hbf18bb28, 32'h40b7f65c} /* (5, 14, 8) {real, imag} */,
  {32'h3f6be5d4, 32'h406dd27f} /* (5, 14, 7) {real, imag} */,
  {32'hbfddd363, 32'hbf8c1c22} /* (5, 14, 6) {real, imag} */,
  {32'h3f8c993c, 32'hc0a51194} /* (5, 14, 5) {real, imag} */,
  {32'hc003b42a, 32'h40a56c98} /* (5, 14, 4) {real, imag} */,
  {32'h3f4aa968, 32'h40d68bd0} /* (5, 14, 3) {real, imag} */,
  {32'h3edc0790, 32'hbf5f6188} /* (5, 14, 2) {real, imag} */,
  {32'hc0758cba, 32'hbf20bb54} /* (5, 14, 1) {real, imag} */,
  {32'h3e1f0248, 32'h3f68bc20} /* (5, 14, 0) {real, imag} */,
  {32'h3f77664a, 32'hbf26f084} /* (5, 13, 15) {real, imag} */,
  {32'hc03705ab, 32'hbe8f1b2a} /* (5, 13, 14) {real, imag} */,
  {32'hc0330ab4, 32'h3fee4091} /* (5, 13, 13) {real, imag} */,
  {32'hbfca1bf6, 32'h401d509c} /* (5, 13, 12) {real, imag} */,
  {32'hc02d6792, 32'h404dc9de} /* (5, 13, 11) {real, imag} */,
  {32'h404e3a60, 32'h40939e20} /* (5, 13, 10) {real, imag} */,
  {32'h40221577, 32'hbe439f28} /* (5, 13, 9) {real, imag} */,
  {32'hc045f1b8, 32'hc0b19c9a} /* (5, 13, 8) {real, imag} */,
  {32'hbfeb6742, 32'hc048e5f4} /* (5, 13, 7) {real, imag} */,
  {32'hbfd115ca, 32'hbfad91aa} /* (5, 13, 6) {real, imag} */,
  {32'hbf24d416, 32'hc0076be6} /* (5, 13, 5) {real, imag} */,
  {32'h40089b01, 32'hbe85d660} /* (5, 13, 4) {real, imag} */,
  {32'h3f98255e, 32'h4059aa60} /* (5, 13, 3) {real, imag} */,
  {32'hbf53acec, 32'h407ffd75} /* (5, 13, 2) {real, imag} */,
  {32'hbe30bb90, 32'hbf992fe0} /* (5, 13, 1) {real, imag} */,
  {32'h3ff9c060, 32'hbfe8f4c3} /* (5, 13, 0) {real, imag} */,
  {32'h3fa06ba8, 32'h40427a2e} /* (5, 12, 15) {real, imag} */,
  {32'h3f7e0992, 32'h405531d0} /* (5, 12, 14) {real, imag} */,
  {32'hbf47d7ba, 32'h3f92df93} /* (5, 12, 13) {real, imag} */,
  {32'h4027136a, 32'h4026a70d} /* (5, 12, 12) {real, imag} */,
  {32'h3f804f5d, 32'h3fa29067} /* (5, 12, 11) {real, imag} */,
  {32'hbf8a09d2, 32'hbe418968} /* (5, 12, 10) {real, imag} */,
  {32'h3f83dc78, 32'hc0213b12} /* (5, 12, 9) {real, imag} */,
  {32'h403d7564, 32'hbf939702} /* (5, 12, 8) {real, imag} */,
  {32'hc0086f7f, 32'h3fabded0} /* (5, 12, 7) {real, imag} */,
  {32'h405c69c6, 32'h409c5a0d} /* (5, 12, 6) {real, imag} */,
  {32'h4044bdc9, 32'h3ffd1731} /* (5, 12, 5) {real, imag} */,
  {32'hbf662ee5, 32'hbd595478} /* (5, 12, 4) {real, imag} */,
  {32'h3f4c6fed, 32'hbf965ed9} /* (5, 12, 3) {real, imag} */,
  {32'hbf93185c, 32'hc048958a} /* (5, 12, 2) {real, imag} */,
  {32'h3f65a61c, 32'hc05abdf0} /* (5, 12, 1) {real, imag} */,
  {32'h3f3260ba, 32'h3ee56d98} /* (5, 12, 0) {real, imag} */,
  {32'hbe789478, 32'hbfdfface} /* (5, 11, 15) {real, imag} */,
  {32'h3f262dc0, 32'hc0216010} /* (5, 11, 14) {real, imag} */,
  {32'h3fa5c9ea, 32'h40075620} /* (5, 11, 13) {real, imag} */,
  {32'h3f21b588, 32'h4016dc72} /* (5, 11, 12) {real, imag} */,
  {32'h3fa0abce, 32'h3fd987c4} /* (5, 11, 11) {real, imag} */,
  {32'h4020470c, 32'hbdaca700} /* (5, 11, 10) {real, imag} */,
  {32'h3fa226d0, 32'hc0853fc2} /* (5, 11, 9) {real, imag} */,
  {32'hbfe1c284, 32'hc07291ed} /* (5, 11, 8) {real, imag} */,
  {32'hbef68240, 32'hc06f7695} /* (5, 11, 7) {real, imag} */,
  {32'hbf822620, 32'hc012ed76} /* (5, 11, 6) {real, imag} */,
  {32'h3e862c94, 32'h3ff047ae} /* (5, 11, 5) {real, imag} */,
  {32'h401cf9de, 32'h40668990} /* (5, 11, 4) {real, imag} */,
  {32'h3ff3b652, 32'h3f4f0b78} /* (5, 11, 3) {real, imag} */,
  {32'h3f3b04b3, 32'hbf87183c} /* (5, 11, 2) {real, imag} */,
  {32'h3faf7676, 32'h3eb28e14} /* (5, 11, 1) {real, imag} */,
  {32'hbeac3c42, 32'hbf657380} /* (5, 11, 0) {real, imag} */,
  {32'hbfca40ee, 32'h3fd9c989} /* (5, 10, 15) {real, imag} */,
  {32'hbf8fe888, 32'hbe45a608} /* (5, 10, 14) {real, imag} */,
  {32'h3dc5b4c8, 32'hbfd24b46} /* (5, 10, 13) {real, imag} */,
  {32'hbf8b04fe, 32'hbfe2ebfc} /* (5, 10, 12) {real, imag} */,
  {32'hbf4a580e, 32'hbfe90511} /* (5, 10, 11) {real, imag} */,
  {32'h3fdf02db, 32'hbf2c2b3d} /* (5, 10, 10) {real, imag} */,
  {32'h3f29497e, 32'hbfcd9396} /* (5, 10, 9) {real, imag} */,
  {32'hbef26ea8, 32'hbfaddffe} /* (5, 10, 8) {real, imag} */,
  {32'hbe700488, 32'hc010c005} /* (5, 10, 7) {real, imag} */,
  {32'hbf9e9ace, 32'hbf45c210} /* (5, 10, 6) {real, imag} */,
  {32'hbfbfa1b8, 32'h3f5a5490} /* (5, 10, 5) {real, imag} */,
  {32'hbf4596ca, 32'hbf83c07e} /* (5, 10, 4) {real, imag} */,
  {32'hc014ed20, 32'hbfffc8ba} /* (5, 10, 3) {real, imag} */,
  {32'hc02cda24, 32'h3ee1ae44} /* (5, 10, 2) {real, imag} */,
  {32'h3d6c6660, 32'h4018fb3c} /* (5, 10, 1) {real, imag} */,
  {32'h3e2642f8, 32'h402469ee} /* (5, 10, 0) {real, imag} */,
  {32'h3f294bca, 32'h3f04d71c} /* (5, 9, 15) {real, imag} */,
  {32'h3f4c6a23, 32'hbe91a29c} /* (5, 9, 14) {real, imag} */,
  {32'h3f7b6d3c, 32'h3f9317aa} /* (5, 9, 13) {real, imag} */,
  {32'hbf377083, 32'h3e8705fe} /* (5, 9, 12) {real, imag} */,
  {32'hbf052568, 32'hbf54037d} /* (5, 9, 11) {real, imag} */,
  {32'hbe9b7010, 32'hbfa87fb5} /* (5, 9, 10) {real, imag} */,
  {32'hbfa92d64, 32'h3fb516e4} /* (5, 9, 9) {real, imag} */,
  {32'hbf76e042, 32'h4003b004} /* (5, 9, 8) {real, imag} */,
  {32'hbf7a341b, 32'h3fd89419} /* (5, 9, 7) {real, imag} */,
  {32'hbf14cbe4, 32'h3f9dc70c} /* (5, 9, 6) {real, imag} */,
  {32'h3fbe6bd0, 32'h3fb03f9f} /* (5, 9, 5) {real, imag} */,
  {32'h3f65692d, 32'h3fdecbca} /* (5, 9, 4) {real, imag} */,
  {32'hbcf12120, 32'h3f0d9032} /* (5, 9, 3) {real, imag} */,
  {32'h3f009916, 32'hbf5e4acd} /* (5, 9, 2) {real, imag} */,
  {32'h3f10ba55, 32'hbec2c732} /* (5, 9, 1) {real, imag} */,
  {32'hbc363940, 32'hbe7248b6} /* (5, 9, 0) {real, imag} */,
  {32'hbd9b7290, 32'h3fa07de5} /* (5, 8, 15) {real, imag} */,
  {32'hbf3fa2f8, 32'h3f568ac6} /* (5, 8, 14) {real, imag} */,
  {32'h3ee4757c, 32'hbf8a7af8} /* (5, 8, 13) {real, imag} */,
  {32'h3ff43268, 32'h3f329b88} /* (5, 8, 12) {real, imag} */,
  {32'h3f4f6332, 32'h3f2f1012} /* (5, 8, 11) {real, imag} */,
  {32'h3f6909b2, 32'h3d173480} /* (5, 8, 10) {real, imag} */,
  {32'hbe42b550, 32'hbeb9c534} /* (5, 8, 9) {real, imag} */,
  {32'hbfba86ec, 32'h3d346c60} /* (5, 8, 8) {real, imag} */,
  {32'hbf85d611, 32'h3f72a968} /* (5, 8, 7) {real, imag} */,
  {32'hbf897f10, 32'h3fc74176} /* (5, 8, 6) {real, imag} */,
  {32'hbf5bfbc0, 32'h3fd86277} /* (5, 8, 5) {real, imag} */,
  {32'hbfa18bfc, 32'h3f26245e} /* (5, 8, 4) {real, imag} */,
  {32'hbfdea800, 32'h3f1c8a5a} /* (5, 8, 3) {real, imag} */,
  {32'hbfe83312, 32'hbd717650} /* (5, 8, 2) {real, imag} */,
  {32'hbe0b9614, 32'hbf79f6dc} /* (5, 8, 1) {real, imag} */,
  {32'h3f429d2c, 32'hbdef1f40} /* (5, 8, 0) {real, imag} */,
  {32'hbe62cd18, 32'h3ed560cc} /* (5, 7, 15) {real, imag} */,
  {32'h3e991892, 32'h3f7d2d66} /* (5, 7, 14) {real, imag} */,
  {32'hbe8a36e8, 32'h3f1e65ef} /* (5, 7, 13) {real, imag} */,
  {32'h3e7add84, 32'h3e8eafae} /* (5, 7, 12) {real, imag} */,
  {32'h3f4e802c, 32'hbf6b1ebd} /* (5, 7, 11) {real, imag} */,
  {32'h3fb4849a, 32'h3f85cc37} /* (5, 7, 10) {real, imag} */,
  {32'h3fe2a704, 32'h3f876fb6} /* (5, 7, 9) {real, imag} */,
  {32'hbe294818, 32'h3d346ae0} /* (5, 7, 8) {real, imag} */,
  {32'hbf095a35, 32'hbe9ce86c} /* (5, 7, 7) {real, imag} */,
  {32'h3f0d77f8, 32'h3d96f278} /* (5, 7, 6) {real, imag} */,
  {32'h3ec9ae70, 32'hbf027e46} /* (5, 7, 5) {real, imag} */,
  {32'h3f847da0, 32'hbfa6ad16} /* (5, 7, 4) {real, imag} */,
  {32'hbffe0d2e, 32'h3ea5cfac} /* (5, 7, 3) {real, imag} */,
  {32'hc01005f2, 32'h3feca782} /* (5, 7, 2) {real, imag} */,
  {32'hbeb039fa, 32'h3fd5f102} /* (5, 7, 1) {real, imag} */,
  {32'h3e917dfa, 32'h3f33f134} /* (5, 7, 0) {real, imag} */,
  {32'hbf8ee4b2, 32'hbed14cc4} /* (5, 6, 15) {real, imag} */,
  {32'h3e0a0a44, 32'hbf5e5ca6} /* (5, 6, 14) {real, imag} */,
  {32'h3f6abf99, 32'h3f10d370} /* (5, 6, 13) {real, imag} */,
  {32'h3ffc7c98, 32'h3f87d278} /* (5, 6, 12) {real, imag} */,
  {32'h3fdee455, 32'h3ecf42ec} /* (5, 6, 11) {real, imag} */,
  {32'h401afffe, 32'h3faae22a} /* (5, 6, 10) {real, imag} */,
  {32'h400b1510, 32'h3e84db60} /* (5, 6, 9) {real, imag} */,
  {32'h3fe38da2, 32'hc02b906f} /* (5, 6, 8) {real, imag} */,
  {32'h3f9299f1, 32'hbf50a5a5} /* (5, 6, 7) {real, imag} */,
  {32'h3eff8772, 32'hbf70a450} /* (5, 6, 6) {real, imag} */,
  {32'h403d3e6e, 32'hc00af6a8} /* (5, 6, 5) {real, imag} */,
  {32'h40547f78, 32'hc066bfa7} /* (5, 6, 4) {real, imag} */,
  {32'h3d85b740, 32'h3eb31d58} /* (5, 6, 3) {real, imag} */,
  {32'hbf86187a, 32'h4003a0ac} /* (5, 6, 2) {real, imag} */,
  {32'hbf9f87b1, 32'h3f550a20} /* (5, 6, 1) {real, imag} */,
  {32'hc02f97f0, 32'hbe4c3f88} /* (5, 6, 0) {real, imag} */,
  {32'hbf4f813e, 32'h3f26097d} /* (5, 5, 15) {real, imag} */,
  {32'hbfcc4d62, 32'hbfdf1741} /* (5, 5, 14) {real, imag} */,
  {32'h40034004, 32'hc0181658} /* (5, 5, 13) {real, imag} */,
  {32'h4029a1ec, 32'hc06ce8e0} /* (5, 5, 12) {real, imag} */,
  {32'h3f01e3fc, 32'hbf8848fa} /* (5, 5, 11) {real, imag} */,
  {32'h3eb6ba6c, 32'h3f3ebaf8} /* (5, 5, 10) {real, imag} */,
  {32'hbc47fd80, 32'hbeb4176c} /* (5, 5, 9) {real, imag} */,
  {32'hc02c623e, 32'hbf960bca} /* (5, 5, 8) {real, imag} */,
  {32'hc088c94c, 32'h3fc93326} /* (5, 5, 7) {real, imag} */,
  {32'hc082c0ac, 32'h4049a00a} /* (5, 5, 6) {real, imag} */,
  {32'hc082dd79, 32'h40799b3b} /* (5, 5, 5) {real, imag} */,
  {32'hbf892d80, 32'h3ea34930} /* (5, 5, 4) {real, imag} */,
  {32'h3f001a3d, 32'hc0688d86} /* (5, 5, 3) {real, imag} */,
  {32'h3fa81ad0, 32'h3e859ad0} /* (5, 5, 2) {real, imag} */,
  {32'h3f19b33c, 32'h40247d40} /* (5, 5, 1) {real, imag} */,
  {32'hbece5fce, 32'h3d53df18} /* (5, 5, 0) {real, imag} */,
  {32'hbff11d1c, 32'hbf21c0e6} /* (5, 4, 15) {real, imag} */,
  {32'h3f462d62, 32'h3fe30f07} /* (5, 4, 14) {real, imag} */,
  {32'h4026580e, 32'h3ff80cfd} /* (5, 4, 13) {real, imag} */,
  {32'h3ef32a4c, 32'h3efaf8e0} /* (5, 4, 12) {real, imag} */,
  {32'h401775e0, 32'h3f4bd04e} /* (5, 4, 11) {real, imag} */,
  {32'h3efb1f22, 32'h3fc724a4} /* (5, 4, 10) {real, imag} */,
  {32'h3f7cbdaf, 32'h3f8443b9} /* (5, 4, 9) {real, imag} */,
  {32'hbf500046, 32'h40aa05c6} /* (5, 4, 8) {real, imag} */,
  {32'hbfb04fe2, 32'h40b21380} /* (5, 4, 7) {real, imag} */,
  {32'h3fd6632c, 32'hbfa8b501} /* (5, 4, 6) {real, imag} */,
  {32'h3fa2a92e, 32'hbd1cd8e0} /* (5, 4, 5) {real, imag} */,
  {32'hbfda22b6, 32'h3e966e61} /* (5, 4, 4) {real, imag} */,
  {32'hc0237f2b, 32'hbfe26aad} /* (5, 4, 3) {real, imag} */,
  {32'hc01897c0, 32'hc04933ae} /* (5, 4, 2) {real, imag} */,
  {32'hc08bb4f4, 32'hc0ad10e8} /* (5, 4, 1) {real, imag} */,
  {32'hc01708f6, 32'hc05dffbb} /* (5, 4, 0) {real, imag} */,
  {32'hbd162b58, 32'h407fd71d} /* (5, 3, 15) {real, imag} */,
  {32'hbeb4aa00, 32'h3eaf0dca} /* (5, 3, 14) {real, imag} */,
  {32'hbec79298, 32'hc02ec823} /* (5, 3, 13) {real, imag} */,
  {32'hc09619a0, 32'h405bd93a} /* (5, 3, 12) {real, imag} */,
  {32'h3f8d0f84, 32'h4035d95e} /* (5, 3, 11) {real, imag} */,
  {32'h408045be, 32'hbfc22990} /* (5, 3, 10) {real, imag} */,
  {32'hbfee1b0a, 32'hc0152776} /* (5, 3, 9) {real, imag} */,
  {32'hbf487980, 32'hbeab9e50} /* (5, 3, 8) {real, imag} */,
  {32'hbe47410c, 32'hbf2cd4f8} /* (5, 3, 7) {real, imag} */,
  {32'h3fbc620a, 32'hbfee3d98} /* (5, 3, 6) {real, imag} */,
  {32'h406adaca, 32'hc008caa8} /* (5, 3, 5) {real, imag} */,
  {32'h40529257, 32'hc07641a6} /* (5, 3, 4) {real, imag} */,
  {32'h3f03442b, 32'hc037489c} /* (5, 3, 3) {real, imag} */,
  {32'hc08fb51a, 32'h3e9e9b28} /* (5, 3, 2) {real, imag} */,
  {32'h3ecadcc0, 32'hc0428d12} /* (5, 3, 1) {real, imag} */,
  {32'h40868ee0, 32'h3fa0c09d} /* (5, 3, 0) {real, imag} */,
  {32'h40915eba, 32'hc09033d9} /* (5, 2, 15) {real, imag} */,
  {32'h3ff7da14, 32'hc0a241b8} /* (5, 2, 14) {real, imag} */,
  {32'hc0bcd78b, 32'hc01f7e8f} /* (5, 2, 13) {real, imag} */,
  {32'hc0af812e, 32'hbd235398} /* (5, 2, 12) {real, imag} */,
  {32'h3f6754ac, 32'h401d5dd2} /* (5, 2, 11) {real, imag} */,
  {32'hbff15626, 32'hbe9fc4a0} /* (5, 2, 10) {real, imag} */,
  {32'hc06e6e7a, 32'hbea0b4a0} /* (5, 2, 9) {real, imag} */,
  {32'hc06d0050, 32'hc00234ad} /* (5, 2, 8) {real, imag} */,
  {32'hbf7afbdc, 32'hbf2ccda4} /* (5, 2, 7) {real, imag} */,
  {32'hbea55044, 32'h409283e4} /* (5, 2, 6) {real, imag} */,
  {32'hc0c2affa, 32'hc06feaf4} /* (5, 2, 5) {real, imag} */,
  {32'h3e8d4ffc, 32'hc08662be} /* (5, 2, 4) {real, imag} */,
  {32'h40adc114, 32'h40691e09} /* (5, 2, 3) {real, imag} */,
  {32'h40f2d487, 32'h40af0d1f} /* (5, 2, 2) {real, imag} */,
  {32'h4110b9ee, 32'h408c0fca} /* (5, 2, 1) {real, imag} */,
  {32'h406df29a, 32'h3e368740} /* (5, 2, 0) {real, imag} */,
  {32'hbf6a227e, 32'hbee8abf0} /* (5, 1, 15) {real, imag} */,
  {32'h4053399f, 32'h400363a7} /* (5, 1, 14) {real, imag} */,
  {32'h410917a2, 32'hbff0b9eb} /* (5, 1, 13) {real, imag} */,
  {32'h406380a4, 32'h404694d5} /* (5, 1, 12) {real, imag} */,
  {32'hbfe3f067, 32'h408bf833} /* (5, 1, 11) {real, imag} */,
  {32'hc0a84c45, 32'h40649778} /* (5, 1, 10) {real, imag} */,
  {32'hc122850a, 32'h40ce837c} /* (5, 1, 9) {real, imag} */,
  {32'hbff51234, 32'h40a899f5} /* (5, 1, 8) {real, imag} */,
  {32'h40264e02, 32'hbfb093ff} /* (5, 1, 7) {real, imag} */,
  {32'h4014f022, 32'hc0c8892c} /* (5, 1, 6) {real, imag} */,
  {32'h40edd002, 32'hbffb2c87} /* (5, 1, 5) {real, imag} */,
  {32'h405590c0, 32'h401436e8} /* (5, 1, 4) {real, imag} */,
  {32'hbfc25008, 32'h409e01e8} /* (5, 1, 3) {real, imag} */,
  {32'h3c29afc0, 32'h407b6e31} /* (5, 1, 2) {real, imag} */,
  {32'h40b4f9f7, 32'h4054733a} /* (5, 1, 1) {real, imag} */,
  {32'h3ffd3f16, 32'h3f90e820} /* (5, 1, 0) {real, imag} */,
  {32'hbf88b629, 32'h3f051832} /* (5, 0, 15) {real, imag} */,
  {32'hc047d1f5, 32'hbe4adc68} /* (5, 0, 14) {real, imag} */,
  {32'h407e3a6a, 32'hc0a2fe00} /* (5, 0, 13) {real, imag} */,
  {32'h40dea0a0, 32'hc0bc220f} /* (5, 0, 12) {real, imag} */,
  {32'h3f4b5162, 32'hc050bcda} /* (5, 0, 11) {real, imag} */,
  {32'hc081909a, 32'hc06af976} /* (5, 0, 10) {real, imag} */,
  {32'h404a8ebd, 32'hc0569bc0} /* (5, 0, 9) {real, imag} */,
  {32'h4065b244, 32'hc077219a} /* (5, 0, 8) {real, imag} */,
  {32'hbff308f3, 32'hc0514d46} /* (5, 0, 7) {real, imag} */,
  {32'h4030def6, 32'h3f0e354f} /* (5, 0, 6) {real, imag} */,
  {32'h40b455c8, 32'hc03cd912} /* (5, 0, 5) {real, imag} */,
  {32'h4037cade, 32'hc00e6324} /* (5, 0, 4) {real, imag} */,
  {32'h40942433, 32'hc024531c} /* (5, 0, 3) {real, imag} */,
  {32'h40b1eb58, 32'h3fd82a54} /* (5, 0, 2) {real, imag} */,
  {32'h3f3f12d5, 32'h3eb1d448} /* (5, 0, 1) {real, imag} */,
  {32'hbf94f5f6, 32'hc0c36efb} /* (5, 0, 0) {real, imag} */,
  {32'h40ca34fd, 32'h40c17528} /* (4, 15, 15) {real, imag} */,
  {32'h40a3e66b, 32'h40e540c2} /* (4, 15, 14) {real, imag} */,
  {32'h40182438, 32'hbf83e4a5} /* (4, 15, 13) {real, imag} */,
  {32'h40a12c60, 32'h4030770c} /* (4, 15, 12) {real, imag} */,
  {32'h408d4cac, 32'hbfd1d80a} /* (4, 15, 11) {real, imag} */,
  {32'hc027dd24, 32'h3f022b64} /* (4, 15, 10) {real, imag} */,
  {32'hbfe8a013, 32'h3e332578} /* (4, 15, 9) {real, imag} */,
  {32'h408c3f9b, 32'h403c25e6} /* (4, 15, 8) {real, imag} */,
  {32'h40d4e06c, 32'h41041038} /* (4, 15, 7) {real, imag} */,
  {32'hbb295a00, 32'h40fdb4da} /* (4, 15, 6) {real, imag} */,
  {32'h40fae020, 32'h4103fa25} /* (4, 15, 5) {real, imag} */,
  {32'h41250b9c, 32'h40bdc92e} /* (4, 15, 4) {real, imag} */,
  {32'h41211621, 32'h40118ffc} /* (4, 15, 3) {real, imag} */,
  {32'h410f4637, 32'h3f8a5be4} /* (4, 15, 2) {real, imag} */,
  {32'h40c42e3a, 32'hc05c1a22} /* (4, 15, 1) {real, imag} */,
  {32'h40733727, 32'hbfaf5268} /* (4, 15, 0) {real, imag} */,
  {32'hc042d9ac, 32'hbf461807} /* (4, 14, 15) {real, imag} */,
  {32'hc01f9162, 32'hc07c46c9} /* (4, 14, 14) {real, imag} */,
  {32'hc04657f0, 32'h3f812c51} /* (4, 14, 13) {real, imag} */,
  {32'hc0da5acc, 32'hc01739b9} /* (4, 14, 12) {real, imag} */,
  {32'hc003dd30, 32'h4000bf1c} /* (4, 14, 11) {real, imag} */,
  {32'hc0926be5, 32'h40d22297} /* (4, 14, 10) {real, imag} */,
  {32'h405b75b5, 32'h3fac76d0} /* (4, 14, 9) {real, imag} */,
  {32'h41010fbc, 32'hc0a2266a} /* (4, 14, 8) {real, imag} */,
  {32'hbfa50717, 32'hc0063403} /* (4, 14, 7) {real, imag} */,
  {32'h3f492936, 32'hc050c349} /* (4, 14, 6) {real, imag} */,
  {32'hc0801fe0, 32'hc11b77de} /* (4, 14, 5) {real, imag} */,
  {32'hc0bc0209, 32'hc1354a57} /* (4, 14, 4) {real, imag} */,
  {32'hc059ce30, 32'hc121b2c6} /* (4, 14, 3) {real, imag} */,
  {32'hbefd95d0, 32'hc113be08} /* (4, 14, 2) {real, imag} */,
  {32'h40b422d9, 32'hc0a97ec6} /* (4, 14, 1) {real, imag} */,
  {32'hbf87bfae, 32'hc041d2fd} /* (4, 14, 0) {real, imag} */,
  {32'hc0188a8d, 32'hc052b0b8} /* (4, 13, 15) {real, imag} */,
  {32'hbf957a54, 32'hbf4b8494} /* (4, 13, 14) {real, imag} */,
  {32'h3fb6bb0b, 32'hbf91face} /* (4, 13, 13) {real, imag} */,
  {32'hc094b5ea, 32'hbfb68304} /* (4, 13, 12) {real, imag} */,
  {32'h3e9f7c1c, 32'hbf7d97c7} /* (4, 13, 11) {real, imag} */,
  {32'h40b65077, 32'h3fe1caec} /* (4, 13, 10) {real, imag} */,
  {32'h3fd607c6, 32'h406e211d} /* (4, 13, 9) {real, imag} */,
  {32'h40823f74, 32'h404e6491} /* (4, 13, 8) {real, imag} */,
  {32'h4029a52f, 32'h407ff065} /* (4, 13, 7) {real, imag} */,
  {32'hbff5fd9d, 32'hc0a2cbd4} /* (4, 13, 6) {real, imag} */,
  {32'h403e48c0, 32'h3fb22e8c} /* (4, 13, 5) {real, imag} */,
  {32'h402cf490, 32'hbfa8d429} /* (4, 13, 4) {real, imag} */,
  {32'h400e29d2, 32'hc0860d51} /* (4, 13, 3) {real, imag} */,
  {32'hbf0fe6ca, 32'h406761c3} /* (4, 13, 2) {real, imag} */,
  {32'h3ef0e9a0, 32'h4043f353} /* (4, 13, 1) {real, imag} */,
  {32'hc03b696b, 32'h3fd53ce6} /* (4, 13, 0) {real, imag} */,
  {32'h3ff79f6d, 32'hbfc5aa56} /* (4, 12, 15) {real, imag} */,
  {32'h40b36eac, 32'h3fbb1244} /* (4, 12, 14) {real, imag} */,
  {32'h404d18b2, 32'h4049f7e6} /* (4, 12, 13) {real, imag} */,
  {32'h3f8050cc, 32'h3ce398e0} /* (4, 12, 12) {real, imag} */,
  {32'hbf34bdc2, 32'hbfc53990} /* (4, 12, 11) {real, imag} */,
  {32'h401faef2, 32'hc0291e70} /* (4, 12, 10) {real, imag} */,
  {32'hc086ee2e, 32'h3f0167e4} /* (4, 12, 9) {real, imag} */,
  {32'hc0c75278, 32'hbf6f6bb3} /* (4, 12, 8) {real, imag} */,
  {32'hc032d70a, 32'hc01660b9} /* (4, 12, 7) {real, imag} */,
  {32'h40103705, 32'h4076b700} /* (4, 12, 6) {real, imag} */,
  {32'h403a5876, 32'h408db666} /* (4, 12, 5) {real, imag} */,
  {32'hc02220e6, 32'h4042d660} /* (4, 12, 4) {real, imag} */,
  {32'hbe9fbe5c, 32'hbeaf3444} /* (4, 12, 3) {real, imag} */,
  {32'hbfea6116, 32'hbd81acc0} /* (4, 12, 2) {real, imag} */,
  {32'hc0c469c2, 32'h4067a7c6} /* (4, 12, 1) {real, imag} */,
  {32'hbe3d6fd0, 32'h4049bdba} /* (4, 12, 0) {real, imag} */,
  {32'hc0524d8a, 32'hc00685bb} /* (4, 11, 15) {real, imag} */,
  {32'hc0031905, 32'hc0221874} /* (4, 11, 14) {real, imag} */,
  {32'h3fe84a6c, 32'hbf224d6e} /* (4, 11, 13) {real, imag} */,
  {32'h402ce082, 32'h40272f42} /* (4, 11, 12) {real, imag} */,
  {32'hc01c98c3, 32'h3fdb9b2e} /* (4, 11, 11) {real, imag} */,
  {32'hbff27934, 32'h3ffe4019} /* (4, 11, 10) {real, imag} */,
  {32'h4066ebb0, 32'h3debecc0} /* (4, 11, 9) {real, imag} */,
  {32'h409c3deb, 32'h404108e2} /* (4, 11, 8) {real, imag} */,
  {32'h400a020d, 32'h406d2686} /* (4, 11, 7) {real, imag} */,
  {32'h402240f4, 32'h402794c0} /* (4, 11, 6) {real, imag} */,
  {32'hbf19984c, 32'h40530756} /* (4, 11, 5) {real, imag} */,
  {32'hc0208808, 32'h400eef14} /* (4, 11, 4) {real, imag} */,
  {32'hc0b020d0, 32'h3fabf5cb} /* (4, 11, 3) {real, imag} */,
  {32'hc0dc703d, 32'h4026b0d8} /* (4, 11, 2) {real, imag} */,
  {32'hc08db547, 32'h3fb030b2} /* (4, 11, 1) {real, imag} */,
  {32'hc09572c0, 32'h3f03534a} /* (4, 11, 0) {real, imag} */,
  {32'h3f97ae6d, 32'hbf31afa7} /* (4, 10, 15) {real, imag} */,
  {32'h3e8aa528, 32'h3f077870} /* (4, 10, 14) {real, imag} */,
  {32'hbf160f6c, 32'hbfa3b3f4} /* (4, 10, 13) {real, imag} */,
  {32'hc00698fe, 32'hc095313f} /* (4, 10, 12) {real, imag} */,
  {32'hc02f7012, 32'hc076a04a} /* (4, 10, 11) {real, imag} */,
  {32'h3f862d18, 32'hc082e8e5} /* (4, 10, 10) {real, imag} */,
  {32'h3fcf9096, 32'hc01178f1} /* (4, 10, 9) {real, imag} */,
  {32'h3eb4c954, 32'hbe935d10} /* (4, 10, 8) {real, imag} */,
  {32'h404ffca3, 32'h400ae632} /* (4, 10, 7) {real, imag} */,
  {32'h4017ca3e, 32'h4002f8c9} /* (4, 10, 6) {real, imag} */,
  {32'h3f0a6b92, 32'h4002b4d0} /* (4, 10, 5) {real, imag} */,
  {32'hbfbae697, 32'h3f9ff8fa} /* (4, 10, 4) {real, imag} */,
  {32'hc0c1fa62, 32'hbf5dd31a} /* (4, 10, 3) {real, imag} */,
  {32'hc08d8dc4, 32'hbbc80800} /* (4, 10, 2) {real, imag} */,
  {32'h3f61c2aa, 32'h403b68c4} /* (4, 10, 1) {real, imag} */,
  {32'h3f961065, 32'h3f7ae5e5} /* (4, 10, 0) {real, imag} */,
  {32'hbfee302b, 32'h3e9e9710} /* (4, 9, 15) {real, imag} */,
  {32'hbf03faf2, 32'h3ef5cc38} /* (4, 9, 14) {real, imag} */,
  {32'hbe4ca238, 32'h3f268d7e} /* (4, 9, 13) {real, imag} */,
  {32'h3f595e5f, 32'h4022e9d5} /* (4, 9, 12) {real, imag} */,
  {32'h3f84bba2, 32'h3fe5bda5} /* (4, 9, 11) {real, imag} */,
  {32'h3f0ec402, 32'h3ef93308} /* (4, 9, 10) {real, imag} */,
  {32'h4020dcb8, 32'h3f19f552} /* (4, 9, 9) {real, imag} */,
  {32'h3fd18f7a, 32'h3ca55780} /* (4, 9, 8) {real, imag} */,
  {32'hbed4a620, 32'hbf91aa0e} /* (4, 9, 7) {real, imag} */,
  {32'h3edfa554, 32'hbfd03e78} /* (4, 9, 6) {real, imag} */,
  {32'hbfd5f27e, 32'hc06170e3} /* (4, 9, 5) {real, imag} */,
  {32'hbf8e4b41, 32'hc017f332} /* (4, 9, 4) {real, imag} */,
  {32'h3ef09e78, 32'hbf36617c} /* (4, 9, 3) {real, imag} */,
  {32'hbf0ad050, 32'hbe31b738} /* (4, 9, 2) {real, imag} */,
  {32'hbe46d528, 32'hbf1ace3f} /* (4, 9, 1) {real, imag} */,
  {32'hbf72737b, 32'h3e072c94} /* (4, 9, 0) {real, imag} */,
  {32'hbf58fca8, 32'hbf5fae44} /* (4, 8, 15) {real, imag} */,
  {32'h3f2a9250, 32'hbf8f1a6e} /* (4, 8, 14) {real, imag} */,
  {32'h3ec578b4, 32'h3f565024} /* (4, 8, 13) {real, imag} */,
  {32'hc03de178, 32'h3fa57ec0} /* (4, 8, 12) {real, imag} */,
  {32'hbf4d4430, 32'h3f8c7ad0} /* (4, 8, 11) {real, imag} */,
  {32'hbfacb43f, 32'h3f54d854} /* (4, 8, 10) {real, imag} */,
  {32'hbfd7193d, 32'h3f3931aa} /* (4, 8, 9) {real, imag} */,
  {32'hbf72a1e8, 32'h3f4e1450} /* (4, 8, 8) {real, imag} */,
  {32'hc05e7bc6, 32'hbff9870a} /* (4, 8, 7) {real, imag} */,
  {32'hc04c084d, 32'hbf86d1cc} /* (4, 8, 6) {real, imag} */,
  {32'hbe828948, 32'h3f1dd4fc} /* (4, 8, 5) {real, imag} */,
  {32'hbf2c6ee4, 32'h3d76d6e0} /* (4, 8, 4) {real, imag} */,
  {32'hbe8c34a4, 32'hbd84a1e0} /* (4, 8, 3) {real, imag} */,
  {32'h3ee36306, 32'h3ea389e2} /* (4, 8, 2) {real, imag} */,
  {32'h3f9bf544, 32'h3e0c1ca0} /* (4, 8, 1) {real, imag} */,
  {32'h3f11f3cc, 32'h3f2226e2} /* (4, 8, 0) {real, imag} */,
  {32'h3eef46dc, 32'hbff40c98} /* (4, 7, 15) {real, imag} */,
  {32'h3d1b23e0, 32'hc023b415} /* (4, 7, 14) {real, imag} */,
  {32'hbfde1b6f, 32'hbfc259b9} /* (4, 7, 13) {real, imag} */,
  {32'hc02b4fde, 32'hc026e207} /* (4, 7, 12) {real, imag} */,
  {32'hbfced358, 32'hbfc93893} /* (4, 7, 11) {real, imag} */,
  {32'h3fa321eb, 32'h3ea335b0} /* (4, 7, 10) {real, imag} */,
  {32'hbe8119e8, 32'h3f534b86} /* (4, 7, 9) {real, imag} */,
  {32'hbfe2e01e, 32'hbf37ec64} /* (4, 7, 8) {real, imag} */,
  {32'h3fb6cfaa, 32'hc006599d} /* (4, 7, 7) {real, imag} */,
  {32'h3fae8bcd, 32'hc04c8bf4} /* (4, 7, 6) {real, imag} */,
  {32'h3f78411c, 32'hbf2628ec} /* (4, 7, 5) {real, imag} */,
  {32'h3fe73389, 32'h3e24c2d8} /* (4, 7, 4) {real, imag} */,
  {32'h3fcd9a56, 32'hc016de76} /* (4, 7, 3) {real, imag} */,
  {32'h40244cdc, 32'h3df832b0} /* (4, 7, 2) {real, imag} */,
  {32'h3ec755dc, 32'h3f1d1161} /* (4, 7, 1) {real, imag} */,
  {32'hbead2bae, 32'h3e39f9d4} /* (4, 7, 0) {real, imag} */,
  {32'hbf2d5406, 32'hbf399609} /* (4, 6, 15) {real, imag} */,
  {32'hc06275de, 32'h3f8162a0} /* (4, 6, 14) {real, imag} */,
  {32'hc0a0f6be, 32'h4086ce39} /* (4, 6, 13) {real, imag} */,
  {32'hc08712a2, 32'h406173e6} /* (4, 6, 12) {real, imag} */,
  {32'hc0317948, 32'h3e278c60} /* (4, 6, 11) {real, imag} */,
  {32'hc0878d29, 32'h3fd95fd4} /* (4, 6, 10) {real, imag} */,
  {32'hc06f5a09, 32'h40548625} /* (4, 6, 9) {real, imag} */,
  {32'h400a2bfe, 32'h401868da} /* (4, 6, 8) {real, imag} */,
  {32'h40344219, 32'hc02b4208} /* (4, 6, 7) {real, imag} */,
  {32'h4039ad94, 32'hbf80e10e} /* (4, 6, 6) {real, imag} */,
  {32'hbf0f1132, 32'h40063ad8} /* (4, 6, 5) {real, imag} */,
  {32'hbe105d68, 32'h40829c46} /* (4, 6, 4) {real, imag} */,
  {32'h4012acf8, 32'h40682e68} /* (4, 6, 3) {real, imag} */,
  {32'h4056eb1a, 32'h4028e7ca} /* (4, 6, 2) {real, imag} */,
  {32'hbf2a9962, 32'h40648162} /* (4, 6, 1) {real, imag} */,
  {32'hbf1b7aa2, 32'h3fe023c8} /* (4, 6, 0) {real, imag} */,
  {32'h3dbe78f0, 32'hbe9c4f62} /* (4, 5, 15) {real, imag} */,
  {32'h40008749, 32'h3fd17def} /* (4, 5, 14) {real, imag} */,
  {32'hbf0a45bc, 32'hc02786d6} /* (4, 5, 13) {real, imag} */,
  {32'hc0106354, 32'hc033dfc0} /* (4, 5, 12) {real, imag} */,
  {32'hbe1126f0, 32'h3daffcf0} /* (4, 5, 11) {real, imag} */,
  {32'h400c1ae2, 32'h3dc79d30} /* (4, 5, 10) {real, imag} */,
  {32'h404b23ac, 32'hc05ae024} /* (4, 5, 9) {real, imag} */,
  {32'h40979169, 32'hc075650e} /* (4, 5, 8) {real, imag} */,
  {32'h403b9631, 32'hc017a914} /* (4, 5, 7) {real, imag} */,
  {32'hc0836d3d, 32'hbefb5920} /* (4, 5, 6) {real, imag} */,
  {32'hbf469fa8, 32'h406fd8d2} /* (4, 5, 5) {real, imag} */,
  {32'h40957875, 32'h410245d6} /* (4, 5, 4) {real, imag} */,
  {32'h3fcbc4f2, 32'h40431aea} /* (4, 5, 3) {real, imag} */,
  {32'hbff95b24, 32'h3f675e65} /* (4, 5, 2) {real, imag} */,
  {32'hc0fcd0c5, 32'h4028055f} /* (4, 5, 1) {real, imag} */,
  {32'hc0793a9c, 32'h3ecab364} /* (4, 5, 0) {real, imag} */,
  {32'h3e4d3468, 32'h3fac174a} /* (4, 4, 15) {real, imag} */,
  {32'h4035d777, 32'h404fa21a} /* (4, 4, 14) {real, imag} */,
  {32'h4088cbd0, 32'hbfb17094} /* (4, 4, 13) {real, imag} */,
  {32'h40db9117, 32'h3f3de27f} /* (4, 4, 12) {real, imag} */,
  {32'hc013339a, 32'h3f0b6667} /* (4, 4, 11) {real, imag} */,
  {32'hc0003390, 32'hbe0f0708} /* (4, 4, 10) {real, imag} */,
  {32'hbfccbdcf, 32'h40503ea3} /* (4, 4, 9) {real, imag} */,
  {32'hbf9f4ba4, 32'hbdd121e8} /* (4, 4, 8) {real, imag} */,
  {32'h3fe1b439, 32'h4015dd33} /* (4, 4, 7) {real, imag} */,
  {32'hc0262673, 32'h3fa76200} /* (4, 4, 6) {real, imag} */,
  {32'hc0846a53, 32'hc008e6ad} /* (4, 4, 5) {real, imag} */,
  {32'hbefc5cdc, 32'h3d5736a0} /* (4, 4, 4) {real, imag} */,
  {32'h3f9b8e63, 32'hc01fc226} /* (4, 4, 3) {real, imag} */,
  {32'h400d53dd, 32'hc0ab86c1} /* (4, 4, 2) {real, imag} */,
  {32'h40c16b74, 32'h3fd9bf43} /* (4, 4, 1) {real, imag} */,
  {32'h407e89d7, 32'h40599dd6} /* (4, 4, 0) {real, imag} */,
  {32'h3f39600f, 32'h3ec9349c} /* (4, 3, 15) {real, imag} */,
  {32'h3fd50078, 32'h3f101700} /* (4, 3, 14) {real, imag} */,
  {32'h407f0cce, 32'h3ff974ac} /* (4, 3, 13) {real, imag} */,
  {32'hc02f2c97, 32'hbf586210} /* (4, 3, 12) {real, imag} */,
  {32'hbdb46900, 32'hc0049d4c} /* (4, 3, 11) {real, imag} */,
  {32'h40a6c27d, 32'hc0219922} /* (4, 3, 10) {real, imag} */,
  {32'h3fe4c40c, 32'hbfb04842} /* (4, 3, 9) {real, imag} */,
  {32'h400dc3e3, 32'hc0247197} /* (4, 3, 8) {real, imag} */,
  {32'h408faf76, 32'h4064034f} /* (4, 3, 7) {real, imag} */,
  {32'h40a71e42, 32'hbf37c434} /* (4, 3, 6) {real, imag} */,
  {32'hbfd28df9, 32'hc0b06f97} /* (4, 3, 5) {real, imag} */,
  {32'hc08e611b, 32'h3ff698b1} /* (4, 3, 4) {real, imag} */,
  {32'h3fd48dc1, 32'h408c7007} /* (4, 3, 3) {real, imag} */,
  {32'h3fa0043d, 32'h408566d4} /* (4, 3, 2) {real, imag} */,
  {32'hc0d7b8b6, 32'h3fc730a2} /* (4, 3, 1) {real, imag} */,
  {32'h3f4286dc, 32'h3ffea9dc} /* (4, 3, 0) {real, imag} */,
  {32'hc088d882, 32'hbee7c252} /* (4, 2, 15) {real, imag} */,
  {32'hc0941867, 32'h3f95fb8e} /* (4, 2, 14) {real, imag} */,
  {32'hbf1be394, 32'hbf04cc72} /* (4, 2, 13) {real, imag} */,
  {32'hc00b0e50, 32'h3dc024e0} /* (4, 2, 12) {real, imag} */,
  {32'hc09ff407, 32'h3ffa8ff0} /* (4, 2, 11) {real, imag} */,
  {32'hbf6c9300, 32'hbff481cc} /* (4, 2, 10) {real, imag} */,
  {32'hc11832be, 32'hc032b426} /* (4, 2, 9) {real, imag} */,
  {32'hc0aafae1, 32'hc0d243d2} /* (4, 2, 8) {real, imag} */,
  {32'hc08651ec, 32'hc11d610d} /* (4, 2, 7) {real, imag} */,
  {32'h40006190, 32'hc02a7d6d} /* (4, 2, 6) {real, imag} */,
  {32'h403689df, 32'hc00a64c6} /* (4, 2, 5) {real, imag} */,
  {32'hc039bdd6, 32'h3e5216c0} /* (4, 2, 4) {real, imag} */,
  {32'hc102bda5, 32'h40621b6a} /* (4, 2, 3) {real, imag} */,
  {32'hc02e1644, 32'h3f99e220} /* (4, 2, 2) {real, imag} */,
  {32'h40578dfe, 32'hc03b3cbc} /* (4, 2, 1) {real, imag} */,
  {32'h40a08914, 32'hbff74a9e} /* (4, 2, 0) {real, imag} */,
  {32'h4028d9fe, 32'h3f6655b8} /* (4, 1, 15) {real, imag} */,
  {32'h3f0c1dc8, 32'h3dad1020} /* (4, 1, 14) {real, imag} */,
  {32'hc0e6e292, 32'h4039b8b2} /* (4, 1, 13) {real, imag} */,
  {32'hc0d86470, 32'hbf84ed48} /* (4, 1, 12) {real, imag} */,
  {32'hbfa330e7, 32'h3f1b93dc} /* (4, 1, 11) {real, imag} */,
  {32'hc0645fd2, 32'h4034f680} /* (4, 1, 10) {real, imag} */,
  {32'h40954079, 32'hc016425c} /* (4, 1, 9) {real, imag} */,
  {32'h409289e1, 32'hc09cb435} /* (4, 1, 8) {real, imag} */,
  {32'hbff29420, 32'hc0f1b7db} /* (4, 1, 7) {real, imag} */,
  {32'hc045582c, 32'hc0e20c0a} /* (4, 1, 6) {real, imag} */,
  {32'h3fb8322e, 32'hc0cd1586} /* (4, 1, 5) {real, imag} */,
  {32'h40a3ac42, 32'hc09cb276} /* (4, 1, 4) {real, imag} */,
  {32'h40abd252, 32'h401fa9c0} /* (4, 1, 3) {real, imag} */,
  {32'hc031cc5c, 32'h41027b90} /* (4, 1, 2) {real, imag} */,
  {32'hc0bfe546, 32'h408369c3} /* (4, 1, 1) {real, imag} */,
  {32'hc08d1234, 32'h4096afa2} /* (4, 1, 0) {real, imag} */,
  {32'hc10168da, 32'h3f377a04} /* (4, 0, 15) {real, imag} */,
  {32'hc114c731, 32'hc0d873ae} /* (4, 0, 14) {real, imag} */,
  {32'hbf7d5d12, 32'hc0da243c} /* (4, 0, 13) {real, imag} */,
  {32'h40e13e3c, 32'hc087e1ee} /* (4, 0, 12) {real, imag} */,
  {32'hbfb9f728, 32'h40184136} /* (4, 0, 11) {real, imag} */,
  {32'hc053c0e0, 32'h408c80fa} /* (4, 0, 10) {real, imag} */,
  {32'h3f59a95e, 32'h40070462} /* (4, 0, 9) {real, imag} */,
  {32'hc0b37fea, 32'h3e81c2b0} /* (4, 0, 8) {real, imag} */,
  {32'hbef149dc, 32'h3fa6f086} /* (4, 0, 7) {real, imag} */,
  {32'h410acf61, 32'h40b00471} /* (4, 0, 6) {real, imag} */,
  {32'h40cbf716, 32'h3fe2ecf6} /* (4, 0, 5) {real, imag} */,
  {32'hc06b15df, 32'h407400d6} /* (4, 0, 4) {real, imag} */,
  {32'hc05cc092, 32'h409d2620} /* (4, 0, 3) {real, imag} */,
  {32'h3f88d412, 32'h3fc84b9e} /* (4, 0, 2) {real, imag} */,
  {32'hbfe5f2a2, 32'hc08eb61d} /* (4, 0, 1) {real, imag} */,
  {32'hc0a0edde, 32'hc0729e2c} /* (4, 0, 0) {real, imag} */,
  {32'hc1562156, 32'hbffed4d0} /* (3, 15, 15) {real, imag} */,
  {32'hc0394340, 32'hc08a58ea} /* (3, 15, 14) {real, imag} */,
  {32'h414675bf, 32'h4066ef62} /* (3, 15, 13) {real, imag} */,
  {32'h3eb3d899, 32'h3f7722b0} /* (3, 15, 12) {real, imag} */,
  {32'h3fcccf26, 32'h407cc1a8} /* (3, 15, 11) {real, imag} */,
  {32'h3e559230, 32'h40c4beec} /* (3, 15, 10) {real, imag} */,
  {32'hc0bedf5b, 32'h40885cd2} /* (3, 15, 9) {real, imag} */,
  {32'h3ee99467, 32'h40bfc9d0} /* (3, 15, 8) {real, imag} */,
  {32'h410446b0, 32'hc0d4f368} /* (3, 15, 7) {real, imag} */,
  {32'h40b460cc, 32'hc129747d} /* (3, 15, 6) {real, imag} */,
  {32'h40c41600, 32'hbf9c7b72} /* (3, 15, 5) {real, imag} */,
  {32'h4112c66d, 32'hbf0fde82} /* (3, 15, 4) {real, imag} */,
  {32'hbf103cb8, 32'hc0532bf3} /* (3, 15, 3) {real, imag} */,
  {32'hc0df82c0, 32'hc00ba57e} /* (3, 15, 2) {real, imag} */,
  {32'h40275de3, 32'hc0b08ebb} /* (3, 15, 1) {real, imag} */,
  {32'hbfde9226, 32'h4004624b} /* (3, 15, 0) {real, imag} */,
  {32'h40ad3dac, 32'hbfe8561a} /* (3, 14, 15) {real, imag} */,
  {32'h402ec3a4, 32'hc061473c} /* (3, 14, 14) {real, imag} */,
  {32'h4092be36, 32'h40bc18e8} /* (3, 14, 13) {real, imag} */,
  {32'h40eef218, 32'h3fbab0f6} /* (3, 14, 12) {real, imag} */,
  {32'hbfb3044e, 32'h402f3f8c} /* (3, 14, 11) {real, imag} */,
  {32'h40a6c569, 32'h401e1a48} /* (3, 14, 10) {real, imag} */,
  {32'h40ac97c2, 32'h40488ebe} /* (3, 14, 9) {real, imag} */,
  {32'hc0423772, 32'h408e05d2} /* (3, 14, 8) {real, imag} */,
  {32'hc059efd0, 32'h3f5d1088} /* (3, 14, 7) {real, imag} */,
  {32'hbfc742d0, 32'hc06ec3b1} /* (3, 14, 6) {real, imag} */,
  {32'h408a8c76, 32'h3ed60c50} /* (3, 14, 5) {real, imag} */,
  {32'h40d56008, 32'h400f7d01} /* (3, 14, 4) {real, imag} */,
  {32'h4017285e, 32'hbfa47788} /* (3, 14, 3) {real, imag} */,
  {32'hc0a67351, 32'hbfc18114} /* (3, 14, 2) {real, imag} */,
  {32'hbf9ae904, 32'hbf923988} /* (3, 14, 1) {real, imag} */,
  {32'hc00da770, 32'hc04ab8db} /* (3, 14, 0) {real, imag} */,
  {32'hc0994dc0, 32'h3ee99b38} /* (3, 13, 15) {real, imag} */,
  {32'hc0f4d63e, 32'h4085bc62} /* (3, 13, 14) {real, imag} */,
  {32'hc0548dbb, 32'hc01ff014} /* (3, 13, 13) {real, imag} */,
  {32'h40dd8fe9, 32'hc0a8a9fa} /* (3, 13, 12) {real, imag} */,
  {32'h3ff94a5e, 32'h403b1f57} /* (3, 13, 11) {real, imag} */,
  {32'hc0cea2f8, 32'hc00f38e5} /* (3, 13, 10) {real, imag} */,
  {32'hc1331a6c, 32'hc0d5e709} /* (3, 13, 9) {real, imag} */,
  {32'hc00f59c8, 32'hbfd80d4f} /* (3, 13, 8) {real, imag} */,
  {32'hbfb85479, 32'h3fc98c11} /* (3, 13, 7) {real, imag} */,
  {32'h3fcbe87c, 32'h3f7424b0} /* (3, 13, 6) {real, imag} */,
  {32'h403edadf, 32'h3f848f7d} /* (3, 13, 5) {real, imag} */,
  {32'h3f39f0c7, 32'h40c54b78} /* (3, 13, 4) {real, imag} */,
  {32'hbf04a34a, 32'h410062e8} /* (3, 13, 3) {real, imag} */,
  {32'hc0073209, 32'hbf1bb38d} /* (3, 13, 2) {real, imag} */,
  {32'hc0b0cdd2, 32'hc07632d2} /* (3, 13, 1) {real, imag} */,
  {32'h408c20df, 32'hbfeeff8a} /* (3, 13, 0) {real, imag} */,
  {32'h40b43022, 32'hbfc8a6d0} /* (3, 12, 15) {real, imag} */,
  {32'hc0168ae1, 32'hc01c3134} /* (3, 12, 14) {real, imag} */,
  {32'hc1137d74, 32'h3ec1b7e0} /* (3, 12, 13) {real, imag} */,
  {32'hc060215e, 32'hc007287d} /* (3, 12, 12) {real, imag} */,
  {32'hc04e1039, 32'h40c0ae6e} /* (3, 12, 11) {real, imag} */,
  {32'hbfc0f7d1, 32'h400b612a} /* (3, 12, 10) {real, imag} */,
  {32'h3f189108, 32'h3f88d152} /* (3, 12, 9) {real, imag} */,
  {32'hc108d1f7, 32'h40c70d3d} /* (3, 12, 8) {real, imag} */,
  {32'hc06a0ce8, 32'h40b3cca4} /* (3, 12, 7) {real, imag} */,
  {32'h4051b3d4, 32'hbe5b2580} /* (3, 12, 6) {real, imag} */,
  {32'h40b1f11e, 32'hc01f2ea3} /* (3, 12, 5) {real, imag} */,
  {32'h3ff4d5c8, 32'hbfebe58f} /* (3, 12, 4) {real, imag} */,
  {32'hbf9e837e, 32'hbf25e388} /* (3, 12, 3) {real, imag} */,
  {32'h40b56b54, 32'hbf4a6442} /* (3, 12, 2) {real, imag} */,
  {32'h4015faff, 32'hc0285ee6} /* (3, 12, 1) {real, imag} */,
  {32'h3f9191a7, 32'hc012cbe8} /* (3, 12, 0) {real, imag} */,
  {32'hbe8805f0, 32'h408dec8c} /* (3, 11, 15) {real, imag} */,
  {32'h40477286, 32'h40b66cb9} /* (3, 11, 14) {real, imag} */,
  {32'hbf05469e, 32'hc044d386} /* (3, 11, 13) {real, imag} */,
  {32'hc0a1128d, 32'hc08e4acd} /* (3, 11, 12) {real, imag} */,
  {32'hc03ae89c, 32'hc0ee8838} /* (3, 11, 11) {real, imag} */,
  {32'h3f262550, 32'hc09aa3f2} /* (3, 11, 10) {real, imag} */,
  {32'hc04766a2, 32'hc01eae43} /* (3, 11, 9) {real, imag} */,
  {32'h3f475114, 32'hc016f107} /* (3, 11, 8) {real, imag} */,
  {32'h40141cce, 32'h3f73386a} /* (3, 11, 7) {real, imag} */,
  {32'hc0146840, 32'h3f99d72b} /* (3, 11, 6) {real, imag} */,
  {32'hc0815834, 32'h403871ee} /* (3, 11, 5) {real, imag} */,
  {32'hc0acf4bb, 32'h40147862} /* (3, 11, 4) {real, imag} */,
  {32'hbf134b46, 32'h3fef7705} /* (3, 11, 3) {real, imag} */,
  {32'h3eccd631, 32'h3f792ac0} /* (3, 11, 2) {real, imag} */,
  {32'h3f976b6c, 32'h4098e34a} /* (3, 11, 1) {real, imag} */,
  {32'h3b743400, 32'h3ff8e82c} /* (3, 11, 0) {real, imag} */,
  {32'h3fe8d0d7, 32'h3f8f1abb} /* (3, 10, 15) {real, imag} */,
  {32'h40547842, 32'hc00743f3} /* (3, 10, 14) {real, imag} */,
  {32'h3fa1256c, 32'hbffc1a32} /* (3, 10, 13) {real, imag} */,
  {32'h3f049282, 32'hbcde4878} /* (3, 10, 12) {real, imag} */,
  {32'h3d0737c0, 32'h3f97bffe} /* (3, 10, 11) {real, imag} */,
  {32'h3f14424a, 32'h403ee4df} /* (3, 10, 10) {real, imag} */,
  {32'hbd471c40, 32'h3f7e1e2a} /* (3, 10, 9) {real, imag} */,
  {32'h3f96fd82, 32'hc061893e} /* (3, 10, 8) {real, imag} */,
  {32'h40249c38, 32'hbf9511dc} /* (3, 10, 7) {real, imag} */,
  {32'h3f699dd0, 32'h408a75ac} /* (3, 10, 6) {real, imag} */,
  {32'h3f8bab8f, 32'h3f32590a} /* (3, 10, 5) {real, imag} */,
  {32'hc06f9e4a, 32'hbe83c9c0} /* (3, 10, 4) {real, imag} */,
  {32'hc047a560, 32'hbf93e848} /* (3, 10, 3) {real, imag} */,
  {32'hbfd3f569, 32'hbf98e360} /* (3, 10, 2) {real, imag} */,
  {32'hc021628e, 32'h4074890f} /* (3, 10, 1) {real, imag} */,
  {32'hbfd93b67, 32'h4027ea38} /* (3, 10, 0) {real, imag} */,
  {32'hbf2fcbd4, 32'h3ebd80f4} /* (3, 9, 15) {real, imag} */,
  {32'hc079322d, 32'h402c30d0} /* (3, 9, 14) {real, imag} */,
  {32'hbfe49d59, 32'h3fdaaced} /* (3, 9, 13) {real, imag} */,
  {32'hbfd079da, 32'hc00e52f1} /* (3, 9, 12) {real, imag} */,
  {32'hbe177ef8, 32'hbfd131ab} /* (3, 9, 11) {real, imag} */,
  {32'hbfa85cea, 32'hbf11a304} /* (3, 9, 10) {real, imag} */,
  {32'hc00cf5a2, 32'hbfb0033d} /* (3, 9, 9) {real, imag} */,
  {32'hbff4a280, 32'h3f8fb188} /* (3, 9, 8) {real, imag} */,
  {32'hbe8621c8, 32'hbe713098} /* (3, 9, 7) {real, imag} */,
  {32'h3ee56c88, 32'hbf587c5c} /* (3, 9, 6) {real, imag} */,
  {32'hbfcfca6a, 32'h3eb06fec} /* (3, 9, 5) {real, imag} */,
  {32'hbf1c6da0, 32'h3fab1b8a} /* (3, 9, 4) {real, imag} */,
  {32'h3fe15f2c, 32'h3f117b73} /* (3, 9, 3) {real, imag} */,
  {32'h402958fc, 32'hbfb7d89c} /* (3, 9, 2) {real, imag} */,
  {32'hbd9d43d8, 32'hbfdffd3d} /* (3, 9, 1) {real, imag} */,
  {32'h3e4acb64, 32'h3d0f2020} /* (3, 9, 0) {real, imag} */,
  {32'h3f05e647, 32'hbd997560} /* (3, 8, 15) {real, imag} */,
  {32'hbfd3ec9e, 32'hbf6c4c57} /* (3, 8, 14) {real, imag} */,
  {32'hbf8cd3f8, 32'h3f397728} /* (3, 8, 13) {real, imag} */,
  {32'hbf0fcb10, 32'h3f65e948} /* (3, 8, 12) {real, imag} */,
  {32'h3f87e420, 32'h3fcbe974} /* (3, 8, 11) {real, imag} */,
  {32'hbf72957c, 32'h3f606a80} /* (3, 8, 10) {real, imag} */,
  {32'h3f0f9488, 32'hc0082bd0} /* (3, 8, 9) {real, imag} */,
  {32'hbe451610, 32'hbf90f1f8} /* (3, 8, 8) {real, imag} */,
  {32'hbf0192d8, 32'hbf71e660} /* (3, 8, 7) {real, imag} */,
  {32'hbf99436b, 32'hbf5cce50} /* (3, 8, 6) {real, imag} */,
  {32'h3faad803, 32'h3e9ddec8} /* (3, 8, 5) {real, imag} */,
  {32'h400df912, 32'h3e9469b0} /* (3, 8, 4) {real, imag} */,
  {32'h3f5a6f44, 32'hc03d1e45} /* (3, 8, 3) {real, imag} */,
  {32'h3fa77f32, 32'hbfb70aca} /* (3, 8, 2) {real, imag} */,
  {32'hbf032764, 32'h3f9d4978} /* (3, 8, 1) {real, imag} */,
  {32'h3f2b435c, 32'hbe3df508} /* (3, 8, 0) {real, imag} */,
  {32'hbf6b1f84, 32'hbdbaff30} /* (3, 7, 15) {real, imag} */,
  {32'hc00113ed, 32'h3f91aee7} /* (3, 7, 14) {real, imag} */,
  {32'hbf92a9e1, 32'h3fb12103} /* (3, 7, 13) {real, imag} */,
  {32'h3eeddbf2, 32'h3ebef9f8} /* (3, 7, 12) {real, imag} */,
  {32'h3fb6becb, 32'hbfdd4205} /* (3, 7, 11) {real, imag} */,
  {32'hbede6a2a, 32'h3f4ff264} /* (3, 7, 10) {real, imag} */,
  {32'h3faa19af, 32'h3fca78b5} /* (3, 7, 9) {real, imag} */,
  {32'h3f8cf930, 32'h3fb45090} /* (3, 7, 8) {real, imag} */,
  {32'h40160a1b, 32'h400e643e} /* (3, 7, 7) {real, imag} */,
  {32'h3fbe6456, 32'h3f34257c} /* (3, 7, 6) {real, imag} */,
  {32'h3e33dcb4, 32'h3f92ee07} /* (3, 7, 5) {real, imag} */,
  {32'hc041123e, 32'hbfb2b5bc} /* (3, 7, 4) {real, imag} */,
  {32'hc02c9e96, 32'hc00daf91} /* (3, 7, 3) {real, imag} */,
  {32'hbf17e2ce, 32'hbfb27352} /* (3, 7, 2) {real, imag} */,
  {32'h3fcf7d10, 32'hbff499f5} /* (3, 7, 1) {real, imag} */,
  {32'h3f7ac783, 32'hbf8c031f} /* (3, 7, 0) {real, imag} */,
  {32'hbe97507c, 32'hbf8351bb} /* (3, 6, 15) {real, imag} */,
  {32'hbf5f5688, 32'hbfd4f2ce} /* (3, 6, 14) {real, imag} */,
  {32'hbfb67e58, 32'hc0215065} /* (3, 6, 13) {real, imag} */,
  {32'hbeb8597c, 32'hbe4f0517} /* (3, 6, 12) {real, imag} */,
  {32'h3faf6ab2, 32'h3dbeb0e0} /* (3, 6, 11) {real, imag} */,
  {32'h3fc5caf1, 32'hc021c351} /* (3, 6, 10) {real, imag} */,
  {32'h3f5c66c0, 32'hbfbe5b0f} /* (3, 6, 9) {real, imag} */,
  {32'hbfe96942, 32'h3ea3e9c0} /* (3, 6, 8) {real, imag} */,
  {32'h3e528470, 32'h3f88c548} /* (3, 6, 7) {real, imag} */,
  {32'hbf01b3a0, 32'hbf859d32} /* (3, 6, 6) {real, imag} */,
  {32'hc09f4267, 32'h401812c6} /* (3, 6, 5) {real, imag} */,
  {32'hc0a441ff, 32'h3fe606f8} /* (3, 6, 4) {real, imag} */,
  {32'hbf76f9d8, 32'h403da87a} /* (3, 6, 3) {real, imag} */,
  {32'hc0566884, 32'h3f851b10} /* (3, 6, 2) {real, imag} */,
  {32'hc09b71a3, 32'h3d4729c0} /* (3, 6, 1) {real, imag} */,
  {32'hbfcbdb2f, 32'hbf011c08} /* (3, 6, 0) {real, imag} */,
  {32'h4061a39a, 32'hc002c462} /* (3, 5, 15) {real, imag} */,
  {32'h410d5328, 32'hc01ff13e} /* (3, 5, 14) {real, imag} */,
  {32'h3fd8f499, 32'h3f0aaa1c} /* (3, 5, 13) {real, imag} */,
  {32'hc0496f6e, 32'hbf9803c1} /* (3, 5, 12) {real, imag} */,
  {32'h3f3bcbd0, 32'hbfb3e21e} /* (3, 5, 11) {real, imag} */,
  {32'h4041ac86, 32'hc0dd15f2} /* (3, 5, 10) {real, imag} */,
  {32'hbf92608c, 32'hc00620c5} /* (3, 5, 9) {real, imag} */,
  {32'hc03ad1e1, 32'h404122f1} /* (3, 5, 8) {real, imag} */,
  {32'hbfaa337e, 32'h3fbe0a85} /* (3, 5, 7) {real, imag} */,
  {32'hc08209ee, 32'hc0801241} /* (3, 5, 6) {real, imag} */,
  {32'hc090ff58, 32'hc1118e30} /* (3, 5, 5) {real, imag} */,
  {32'hbf811530, 32'hc075e924} /* (3, 5, 4) {real, imag} */,
  {32'h3f6dd3a6, 32'h3f91d8c5} /* (3, 5, 3) {real, imag} */,
  {32'h3e910617, 32'hc0744e9e} /* (3, 5, 2) {real, imag} */,
  {32'hbff09708, 32'hc0d09002} /* (3, 5, 1) {real, imag} */,
  {32'hc00c49d8, 32'hbfa7f5b8} /* (3, 5, 0) {real, imag} */,
  {32'h404e34fb, 32'h403817b8} /* (3, 4, 15) {real, imag} */,
  {32'h4027b99b, 32'h3de7a8f0} /* (3, 4, 14) {real, imag} */,
  {32'hc034d7ca, 32'hc0b27098} /* (3, 4, 13) {real, imag} */,
  {32'hc0345eb6, 32'hc0b827c4} /* (3, 4, 12) {real, imag} */,
  {32'h4002f943, 32'hc061cecd} /* (3, 4, 11) {real, imag} */,
  {32'hbf86fee3, 32'hc06b6c76} /* (3, 4, 10) {real, imag} */,
  {32'hc10cd18c, 32'hc0df6170} /* (3, 4, 9) {real, imag} */,
  {32'hc00ca583, 32'hc0f0aa6f} /* (3, 4, 8) {real, imag} */,
  {32'hc03757c8, 32'hc02bed9c} /* (3, 4, 7) {real, imag} */,
  {32'hc0fc6172, 32'h40dd96df} /* (3, 4, 6) {real, imag} */,
  {32'hc12af485, 32'h3fc67e2a} /* (3, 4, 5) {real, imag} */,
  {32'hc11043b9, 32'hbfc5db19} /* (3, 4, 4) {real, imag} */,
  {32'h3ef5b258, 32'h3f812b48} /* (3, 4, 3) {real, imag} */,
  {32'h40918854, 32'hbe897bcc} /* (3, 4, 2) {real, imag} */,
  {32'h3ff68b42, 32'hbeca84c0} /* (3, 4, 1) {real, imag} */,
  {32'h402c1f50, 32'h3ec36994} /* (3, 4, 0) {real, imag} */,
  {32'h40909bc0, 32'h40ca2f34} /* (3, 3, 15) {real, imag} */,
  {32'h4092036c, 32'h40a68358} /* (3, 3, 14) {real, imag} */,
  {32'hbfd54192, 32'hbdf57e20} /* (3, 3, 13) {real, imag} */,
  {32'h40861ea3, 32'h3fdef296} /* (3, 3, 12) {real, imag} */,
  {32'hc0623bf1, 32'h3e182e90} /* (3, 3, 11) {real, imag} */,
  {32'hc090a77c, 32'h4037598f} /* (3, 3, 10) {real, imag} */,
  {32'h3f3c93e8, 32'h41023446} /* (3, 3, 9) {real, imag} */,
  {32'h40bf22b4, 32'hbf35582a} /* (3, 3, 8) {real, imag} */,
  {32'h40651ff0, 32'hc032dd9a} /* (3, 3, 7) {real, imag} */,
  {32'h4117ce8e, 32'h40ab5920} /* (3, 3, 6) {real, imag} */,
  {32'h40c3c09c, 32'h3f0e403a} /* (3, 3, 5) {real, imag} */,
  {32'hbd765ff0, 32'hbfc28c06} /* (3, 3, 4) {real, imag} */,
  {32'hc00ca082, 32'hbffbb364} /* (3, 3, 3) {real, imag} */,
  {32'hbfecabc0, 32'h3f9b8f16} /* (3, 3, 2) {real, imag} */,
  {32'hbe2b2fe0, 32'hc06f3756} /* (3, 3, 1) {real, imag} */,
  {32'hbf85f555, 32'hc0e3926a} /* (3, 3, 0) {real, imag} */,
  {32'hc04822b8, 32'h401475df} /* (3, 2, 15) {real, imag} */,
  {32'hc1180530, 32'h40eff4e2} /* (3, 2, 14) {real, imag} */,
  {32'hc14e5079, 32'h4116dfe2} /* (3, 2, 13) {real, imag} */,
  {32'hc14059c2, 32'hbf67bffb} /* (3, 2, 12) {real, imag} */,
  {32'hc0bf5e92, 32'hc0a36e58} /* (3, 2, 11) {real, imag} */,
  {32'h3d7dff80, 32'hbe8aa6ac} /* (3, 2, 10) {real, imag} */,
  {32'h401ef9c4, 32'hc01b6a30} /* (3, 2, 9) {real, imag} */,
  {32'h408937d2, 32'hbfce95a2} /* (3, 2, 8) {real, imag} */,
  {32'hbef84f58, 32'hc04d0604} /* (3, 2, 7) {real, imag} */,
  {32'hc11cc0e5, 32'hc10ce28e} /* (3, 2, 6) {real, imag} */,
  {32'hc0f2994e, 32'hc103442c} /* (3, 2, 5) {real, imag} */,
  {32'h406ca0a0, 32'hbf5ee624} /* (3, 2, 4) {real, imag} */,
  {32'h3fd1a3a8, 32'h3f5e5d11} /* (3, 2, 3) {real, imag} */,
  {32'hbc411600, 32'hbfe35a6c} /* (3, 2, 2) {real, imag} */,
  {32'h40d408ef, 32'hbfa22e48} /* (3, 2, 1) {real, imag} */,
  {32'h40f67578, 32'h403e03cb} /* (3, 2, 0) {real, imag} */,
  {32'h3f851744, 32'hc0708b8c} /* (3, 1, 15) {real, imag} */,
  {32'h4007af3a, 32'hbc655000} /* (3, 1, 14) {real, imag} */,
  {32'hc00430b8, 32'h4007d16e} /* (3, 1, 13) {real, imag} */,
  {32'hbe936ebd, 32'h416c3a87} /* (3, 1, 12) {real, imag} */,
  {32'h40b7b798, 32'h412abfdc} /* (3, 1, 11) {real, imag} */,
  {32'h4066b7a7, 32'h40f704e4} /* (3, 1, 10) {real, imag} */,
  {32'h401ad572, 32'hbeac7700} /* (3, 1, 9) {real, imag} */,
  {32'hbf90b43a, 32'hbf920188} /* (3, 1, 8) {real, imag} */,
  {32'hc11aaf28, 32'h3f80705e} /* (3, 1, 7) {real, imag} */,
  {32'hbfd9ab86, 32'hbfb65448} /* (3, 1, 6) {real, imag} */,
  {32'hbfaf29b2, 32'hc0e6fe2a} /* (3, 1, 5) {real, imag} */,
  {32'hbc191400, 32'hc0288d2a} /* (3, 1, 4) {real, imag} */,
  {32'hbfa31090, 32'h4071555f} /* (3, 1, 3) {real, imag} */,
  {32'hc138642a, 32'h4081054b} /* (3, 1, 2) {real, imag} */,
  {32'hc0be56a6, 32'h4111ab18} /* (3, 1, 1) {real, imag} */,
  {32'hc08918b8, 32'h4001e309} /* (3, 1, 0) {real, imag} */,
  {32'h401f79f8, 32'hbe033b68} /* (3, 0, 15) {real, imag} */,
  {32'h40c83d92, 32'h4033d667} /* (3, 0, 14) {real, imag} */,
  {32'hc10e5195, 32'hc091bf7d} /* (3, 0, 13) {real, imag} */,
  {32'hc198f436, 32'hc101bc4e} /* (3, 0, 12) {real, imag} */,
  {32'hbe323c60, 32'hc13f7f12} /* (3, 0, 11) {real, imag} */,
  {32'h40d8c476, 32'hc060d794} /* (3, 0, 10) {real, imag} */,
  {32'hc048d1a0, 32'hc0906081} /* (3, 0, 9) {real, imag} */,
  {32'hc01e1339, 32'hc03eaf82} /* (3, 0, 8) {real, imag} */,
  {32'h41500a76, 32'hc0de48c2} /* (3, 0, 7) {real, imag} */,
  {32'h3f072472, 32'h3f479a08} /* (3, 0, 6) {real, imag} */,
  {32'hbe345e38, 32'h4097bab6} /* (3, 0, 5) {real, imag} */,
  {32'h41122348, 32'hc08ba01f} /* (3, 0, 4) {real, imag} */,
  {32'h40b185b2, 32'hc1080d6d} /* (3, 0, 3) {real, imag} */,
  {32'h40bda81a, 32'hc06fe571} /* (3, 0, 2) {real, imag} */,
  {32'h40e433d0, 32'hc011f49a} /* (3, 0, 1) {real, imag} */,
  {32'h4084b746, 32'hbec7d8c4} /* (3, 0, 0) {real, imag} */,
  {32'h3f843748, 32'h4046e772} /* (2, 15, 15) {real, imag} */,
  {32'hc0e5b0f8, 32'h40f4556f} /* (2, 15, 14) {real, imag} */,
  {32'hc1724658, 32'h4123f6e6} /* (2, 15, 13) {real, imag} */,
  {32'hc1307b8c, 32'h40d32c28} /* (2, 15, 12) {real, imag} */,
  {32'hbf91930b, 32'hc0df3dfa} /* (2, 15, 11) {real, imag} */,
  {32'hc01f5d9c, 32'hc1658447} /* (2, 15, 10) {real, imag} */,
  {32'hc0567d28, 32'hc00a90f8} /* (2, 15, 9) {real, imag} */,
  {32'hbf3d5a6e, 32'hbf9ce4e4} /* (2, 15, 8) {real, imag} */,
  {32'h3fcb7adc, 32'hbfd5a735} /* (2, 15, 7) {real, imag} */,
  {32'hbfcad94a, 32'hc0ce5bfe} /* (2, 15, 6) {real, imag} */,
  {32'hc115883a, 32'hbf09143c} /* (2, 15, 5) {real, imag} */,
  {32'hc0e5a97f, 32'h40c03896} /* (2, 15, 4) {real, imag} */,
  {32'hc00685f2, 32'hc00fd24d} /* (2, 15, 3) {real, imag} */,
  {32'hc08dcf69, 32'hc0cd03ed} /* (2, 15, 2) {real, imag} */,
  {32'hc0a713bc, 32'hc08b4efc} /* (2, 15, 1) {real, imag} */,
  {32'hc06430d4, 32'h40a12668} /* (2, 15, 0) {real, imag} */,
  {32'hc0c68d29, 32'hc0c6ddfd} /* (2, 14, 15) {real, imag} */,
  {32'hc17eb554, 32'hc1425ce8} /* (2, 14, 14) {real, imag} */,
  {32'hc1933e7e, 32'hc1473472} /* (2, 14, 13) {real, imag} */,
  {32'hc0d76bec, 32'hc1592b99} /* (2, 14, 12) {real, imag} */,
  {32'h40811a01, 32'hc13301ad} /* (2, 14, 11) {real, imag} */,
  {32'h40a5e47e, 32'hc025e8c3} /* (2, 14, 10) {real, imag} */,
  {32'hbfd8a368, 32'h40c808a8} /* (2, 14, 9) {real, imag} */,
  {32'h3fd0e345, 32'h40a708b3} /* (2, 14, 8) {real, imag} */,
  {32'h410c53e4, 32'h3fad9ca2} /* (2, 14, 7) {real, imag} */,
  {32'h40fe5e1e, 32'h40598318} /* (2, 14, 6) {real, imag} */,
  {32'h3e58d1b0, 32'h41066d77} /* (2, 14, 5) {real, imag} */,
  {32'hc0506546, 32'h4140b301} /* (2, 14, 4) {real, imag} */,
  {32'h3fd80113, 32'h415458da} /* (2, 14, 3) {real, imag} */,
  {32'h3fa6ef1a, 32'h40929c43} /* (2, 14, 2) {real, imag} */,
  {32'h405bec6e, 32'hc078d2b7} /* (2, 14, 1) {real, imag} */,
  {32'h3fe87f29, 32'hc0214fb7} /* (2, 14, 0) {real, imag} */,
  {32'h4003d5e3, 32'h407ded5a} /* (2, 13, 15) {real, imag} */,
  {32'hc0357920, 32'h407eb460} /* (2, 13, 14) {real, imag} */,
  {32'hbf51ec4b, 32'hc0fe02a7} /* (2, 13, 13) {real, imag} */,
  {32'h4090278f, 32'hc047a296} /* (2, 13, 12) {real, imag} */,
  {32'h40f61dca, 32'hc0133d76} /* (2, 13, 11) {real, imag} */,
  {32'hc00964e5, 32'hc0af92c8} /* (2, 13, 10) {real, imag} */,
  {32'hc056e7e2, 32'hc06a1a29} /* (2, 13, 9) {real, imag} */,
  {32'h3eed36ac, 32'h3fa63568} /* (2, 13, 8) {real, imag} */,
  {32'h3f8d1688, 32'h3fd8172a} /* (2, 13, 7) {real, imag} */,
  {32'hbf533828, 32'hc10a22e2} /* (2, 13, 6) {real, imag} */,
  {32'hc08568da, 32'hbffe3b3b} /* (2, 13, 5) {real, imag} */,
  {32'hbfac649e, 32'h40e5ad0b} /* (2, 13, 4) {real, imag} */,
  {32'hc0912418, 32'h40982a7b} /* (2, 13, 3) {real, imag} */,
  {32'hc1118e04, 32'hc03fb474} /* (2, 13, 2) {real, imag} */,
  {32'h3fb5d257, 32'h3fa6df1f} /* (2, 13, 1) {real, imag} */,
  {32'h40a7aaa1, 32'h40b0fbb0} /* (2, 13, 0) {real, imag} */,
  {32'hc0949e63, 32'hbfe379c9} /* (2, 12, 15) {real, imag} */,
  {32'hc100af50, 32'hc0d9ea35} /* (2, 12, 14) {real, imag} */,
  {32'hbfdf78f7, 32'hc0bb19a2} /* (2, 12, 13) {real, imag} */,
  {32'h408b517e, 32'h40f15c8b} /* (2, 12, 12) {real, imag} */,
  {32'h401c88a7, 32'h40878291} /* (2, 12, 11) {real, imag} */,
  {32'hc0c476be, 32'hc00e9804} /* (2, 12, 10) {real, imag} */,
  {32'hc11a034f, 32'h40625c76} /* (2, 12, 9) {real, imag} */,
  {32'hc09024f5, 32'h407b823e} /* (2, 12, 8) {real, imag} */,
  {32'h41326866, 32'hc0865480} /* (2, 12, 7) {real, imag} */,
  {32'h40c2378a, 32'h40932802} /* (2, 12, 6) {real, imag} */,
  {32'hbfdd92c0, 32'h41275d9a} /* (2, 12, 5) {real, imag} */,
  {32'hbefb5432, 32'h402fe0f2} /* (2, 12, 4) {real, imag} */,
  {32'h40ee8c85, 32'hc038b114} /* (2, 12, 3) {real, imag} */,
  {32'h3f901178, 32'hbff15644} /* (2, 12, 2) {real, imag} */,
  {32'h40a9673f, 32'h3f499ea0} /* (2, 12, 1) {real, imag} */,
  {32'h40b56bec, 32'hbed54c20} /* (2, 12, 0) {real, imag} */,
  {32'h3e61005c, 32'hc0073579} /* (2, 11, 15) {real, imag} */,
  {32'h40b00d8e, 32'h404ec903} /* (2, 11, 14) {real, imag} */,
  {32'h40d82e51, 32'h40d0768b} /* (2, 11, 13) {real, imag} */,
  {32'h402ca191, 32'h400e0793} /* (2, 11, 12) {real, imag} */,
  {32'h40a40a93, 32'h40221c74} /* (2, 11, 11) {real, imag} */,
  {32'hc0959e7f, 32'h40916bea} /* (2, 11, 10) {real, imag} */,
  {32'hc06a1fb7, 32'h4095e5bc} /* (2, 11, 9) {real, imag} */,
  {32'hbe633e28, 32'h40273858} /* (2, 11, 8) {real, imag} */,
  {32'hbed07670, 32'h404c1f7d} /* (2, 11, 7) {real, imag} */,
  {32'h3f2996b0, 32'h40ae805f} /* (2, 11, 6) {real, imag} */,
  {32'hbcc29300, 32'h409865ba} /* (2, 11, 5) {real, imag} */,
  {32'hbf7c9f4c, 32'hbfee0eb2} /* (2, 11, 4) {real, imag} */,
  {32'hbfe1fa7a, 32'hc008509a} /* (2, 11, 3) {real, imag} */,
  {32'h3f438178, 32'hc06ab50a} /* (2, 11, 2) {real, imag} */,
  {32'hbed6bc9c, 32'hc03945ca} /* (2, 11, 1) {real, imag} */,
  {32'h401d261f, 32'hbfac3619} /* (2, 11, 0) {real, imag} */,
  {32'hbf0f93c5, 32'hbfb188d9} /* (2, 10, 15) {real, imag} */,
  {32'h3f01d7f8, 32'hbff5f5eb} /* (2, 10, 14) {real, imag} */,
  {32'h4049400e, 32'hbfb6df2e} /* (2, 10, 13) {real, imag} */,
  {32'h3fc17236, 32'h3ef087b2} /* (2, 10, 12) {real, imag} */,
  {32'hbf55aed0, 32'h3ffa1840} /* (2, 10, 11) {real, imag} */,
  {32'h3f815899, 32'hbfb6edd9} /* (2, 10, 10) {real, imag} */,
  {32'h3f8a5afe, 32'hc041bd02} /* (2, 10, 9) {real, imag} */,
  {32'hc020a6a0, 32'hbed57c74} /* (2, 10, 8) {real, imag} */,
  {32'hc0429831, 32'h3fb70730} /* (2, 10, 7) {real, imag} */,
  {32'h3fff1e40, 32'h3f909a45} /* (2, 10, 6) {real, imag} */,
  {32'h409cf436, 32'hbf6c09bd} /* (2, 10, 5) {real, imag} */,
  {32'h4013ffbc, 32'h3f843569} /* (2, 10, 4) {real, imag} */,
  {32'h3fcc0130, 32'h40680fab} /* (2, 10, 3) {real, imag} */,
  {32'h3f77e352, 32'h3fe6dec0} /* (2, 10, 2) {real, imag} */,
  {32'h3fb49a70, 32'h4081908a} /* (2, 10, 1) {real, imag} */,
  {32'hbf41402a, 32'h3f8aefe9} /* (2, 10, 0) {real, imag} */,
  {32'h40503180, 32'h3f927568} /* (2, 9, 15) {real, imag} */,
  {32'h3f7947a1, 32'hbf096fb4} /* (2, 9, 14) {real, imag} */,
  {32'hc01fc530, 32'hbfb51530} /* (2, 9, 13) {real, imag} */,
  {32'h3f68ab5e, 32'h3f2c8bd6} /* (2, 9, 12) {real, imag} */,
  {32'h3f626838, 32'h3f81d11e} /* (2, 9, 11) {real, imag} */,
  {32'h3fd3ac0e, 32'hc003c448} /* (2, 9, 10) {real, imag} */,
  {32'h3f0df650, 32'hbfa27b84} /* (2, 9, 9) {real, imag} */,
  {32'hbda16cc8, 32'h3ea99c60} /* (2, 9, 8) {real, imag} */,
  {32'h3f6626ea, 32'h3fa90439} /* (2, 9, 7) {real, imag} */,
  {32'h4026136f, 32'h3f20a98a} /* (2, 9, 6) {real, imag} */,
  {32'h401e8b96, 32'hbfc5d5a5} /* (2, 9, 5) {real, imag} */,
  {32'h3fc0939f, 32'hc026a0c5} /* (2, 9, 4) {real, imag} */,
  {32'hbfeb2bf2, 32'h3e10f538} /* (2, 9, 3) {real, imag} */,
  {32'hbf817f0c, 32'h3fb2eff4} /* (2, 9, 2) {real, imag} */,
  {32'hc01a1ab5, 32'hbf7bb244} /* (2, 9, 1) {real, imag} */,
  {32'hbf8cf6c5, 32'hbff717b3} /* (2, 9, 0) {real, imag} */,
  {32'hbfbb733f, 32'hbfe206cf} /* (2, 8, 15) {real, imag} */,
  {32'h3f1fc818, 32'hc0074eb0} /* (2, 8, 14) {real, imag} */,
  {32'h3faa8556, 32'hbf282808} /* (2, 8, 13) {real, imag} */,
  {32'h3ec0b7c0, 32'hbfa8024c} /* (2, 8, 12) {real, imag} */,
  {32'h3f4d305a, 32'hbed76880} /* (2, 8, 11) {real, imag} */,
  {32'h3f74bc2c, 32'hbed36784} /* (2, 8, 10) {real, imag} */,
  {32'h3daa9ed0, 32'h3ff31df2} /* (2, 8, 9) {real, imag} */,
  {32'hbf2ca090, 32'h40485a06} /* (2, 8, 8) {real, imag} */,
  {32'hbf2d6a48, 32'h401e0390} /* (2, 8, 7) {real, imag} */,
  {32'hbfe37036, 32'hbfd55f00} /* (2, 8, 6) {real, imag} */,
  {32'hc00d41f4, 32'hbeebeae0} /* (2, 8, 5) {real, imag} */,
  {32'hbf8edd7e, 32'h407c35b4} /* (2, 8, 4) {real, imag} */,
  {32'h40564d5b, 32'h405d981e} /* (2, 8, 3) {real, imag} */,
  {32'h406b5331, 32'h3fcf16c6} /* (2, 8, 2) {real, imag} */,
  {32'hbf17ab58, 32'h40570cd8} /* (2, 8, 1) {real, imag} */,
  {32'hc0085853, 32'h402cf0b7} /* (2, 8, 0) {real, imag} */,
  {32'hbf179efc, 32'h3d1c3580} /* (2, 7, 15) {real, imag} */,
  {32'h3f38e769, 32'hbf6f674c} /* (2, 7, 14) {real, imag} */,
  {32'h4078f63e, 32'hbf5524ff} /* (2, 7, 13) {real, imag} */,
  {32'h3eb75fdc, 32'hbeea0e9c} /* (2, 7, 12) {real, imag} */,
  {32'h3fdfd17a, 32'hbf32019b} /* (2, 7, 11) {real, imag} */,
  {32'h402bda6d, 32'hbf80a2c0} /* (2, 7, 10) {real, imag} */,
  {32'hbfd31d4c, 32'hbf34f018} /* (2, 7, 9) {real, imag} */,
  {32'hbfe14746, 32'hbf7feb5c} /* (2, 7, 8) {real, imag} */,
  {32'hbf295f62, 32'hbf7e540a} /* (2, 7, 7) {real, imag} */,
  {32'h3f5ac99c, 32'h404599da} /* (2, 7, 6) {real, imag} */,
  {32'h4025244a, 32'h4025fc80} /* (2, 7, 5) {real, imag} */,
  {32'h3efc1524, 32'h400926e9} /* (2, 7, 4) {real, imag} */,
  {32'h3fe41b06, 32'hbfb3e725} /* (2, 7, 3) {real, imag} */,
  {32'hbf2d58a0, 32'hc03f9822} /* (2, 7, 2) {real, imag} */,
  {32'hc02ce289, 32'h3f0edda4} /* (2, 7, 1) {real, imag} */,
  {32'h3f8d76cd, 32'hbe102518} /* (2, 7, 0) {real, imag} */,
  {32'h3ee48046, 32'hbeb13bbc} /* (2, 6, 15) {real, imag} */,
  {32'h4017a474, 32'hbf943035} /* (2, 6, 14) {real, imag} */,
  {32'hbf8f5b64, 32'hbda0d1e0} /* (2, 6, 13) {real, imag} */,
  {32'h405fa6af, 32'hbf67cef7} /* (2, 6, 12) {real, imag} */,
  {32'h406bdb12, 32'h4053f92e} /* (2, 6, 11) {real, imag} */,
  {32'h400f2cbe, 32'h3f30e1ca} /* (2, 6, 10) {real, imag} */,
  {32'hbf1217f4, 32'hc043003c} /* (2, 6, 9) {real, imag} */,
  {32'h40029168, 32'h3fc010b3} /* (2, 6, 8) {real, imag} */,
  {32'hbfc37bc2, 32'h40483106} /* (2, 6, 7) {real, imag} */,
  {32'hc08f3c0a, 32'hbe1f91b8} /* (2, 6, 6) {real, imag} */,
  {32'h3ea36108, 32'h3ea23baa} /* (2, 6, 5) {real, imag} */,
  {32'hc09c4de6, 32'hbfe1e8d7} /* (2, 6, 4) {real, imag} */,
  {32'hc0c72654, 32'h401a9cb3} /* (2, 6, 3) {real, imag} */,
  {32'hbf6d3c96, 32'h404d9fac} /* (2, 6, 2) {real, imag} */,
  {32'hbe4d59fc, 32'hbfa366d5} /* (2, 6, 1) {real, imag} */,
  {32'hbf7bf162, 32'h3ff59053} /* (2, 6, 0) {real, imag} */,
  {32'hbfc2eae0, 32'hbe6ce860} /* (2, 5, 15) {real, imag} */,
  {32'hc0871b10, 32'hbf62ff34} /* (2, 5, 14) {real, imag} */,
  {32'hc0c5e813, 32'hc0040c22} /* (2, 5, 13) {real, imag} */,
  {32'hbfa2d20e, 32'hc0783345} /* (2, 5, 12) {real, imag} */,
  {32'hc05f4d92, 32'h40ce8286} /* (2, 5, 11) {real, imag} */,
  {32'hc0558982, 32'h40fdf62a} /* (2, 5, 10) {real, imag} */,
  {32'h40c6fed8, 32'h4017936a} /* (2, 5, 9) {real, imag} */,
  {32'h3f8823e1, 32'h401c18ba} /* (2, 5, 8) {real, imag} */,
  {32'h3ecf8610, 32'hbfc710fa} /* (2, 5, 7) {real, imag} */,
  {32'h4083322e, 32'h4090544b} /* (2, 5, 6) {real, imag} */,
  {32'hc01f37c8, 32'h40f4ad26} /* (2, 5, 5) {real, imag} */,
  {32'h3eb1a868, 32'h3de30960} /* (2, 5, 4) {real, imag} */,
  {32'hc062bcfb, 32'hc0442ecc} /* (2, 5, 3) {real, imag} */,
  {32'hbffb7734, 32'h3f8886d8} /* (2, 5, 2) {real, imag} */,
  {32'h404408b6, 32'h403d72d6} /* (2, 5, 1) {real, imag} */,
  {32'hbf0f1874, 32'h3ff45587} /* (2, 5, 0) {real, imag} */,
  {32'hc0c150e1, 32'h40a0226a} /* (2, 4, 15) {real, imag} */,
  {32'hc0d2a300, 32'h41169f12} /* (2, 4, 14) {real, imag} */,
  {32'h3e94ae24, 32'h40ca276e} /* (2, 4, 13) {real, imag} */,
  {32'h3f713aa0, 32'hbf880a04} /* (2, 4, 12) {real, imag} */,
  {32'hc0171099, 32'hc0ad1c21} /* (2, 4, 11) {real, imag} */,
  {32'hc04f69e0, 32'h405141f2} /* (2, 4, 10) {real, imag} */,
  {32'hbf2cd3f0, 32'h40154cf8} /* (2, 4, 9) {real, imag} */,
  {32'hc09f0fc1, 32'h3fd7052c} /* (2, 4, 8) {real, imag} */,
  {32'hbf1f3ad8, 32'h3fb61376} /* (2, 4, 7) {real, imag} */,
  {32'hc091595a, 32'hc07c870c} /* (2, 4, 6) {real, imag} */,
  {32'hc0c64c3a, 32'hc08dd898} /* (2, 4, 5) {real, imag} */,
  {32'hbeb826b2, 32'hc07a0fda} /* (2, 4, 4) {real, imag} */,
  {32'h407f276e, 32'hc0e8cf12} /* (2, 4, 3) {real, imag} */,
  {32'h40a4276a, 32'hc0802794} /* (2, 4, 2) {real, imag} */,
  {32'hc0ce8a97, 32'hc0aa20e2} /* (2, 4, 1) {real, imag} */,
  {32'hc0862a0a, 32'hc080211d} /* (2, 4, 0) {real, imag} */,
  {32'h407b3e59, 32'hbf257dca} /* (2, 3, 15) {real, imag} */,
  {32'h40939506, 32'h41230f42} /* (2, 3, 14) {real, imag} */,
  {32'hbf760f13, 32'h4000f572} /* (2, 3, 13) {real, imag} */,
  {32'hc10e8358, 32'hc0f84a0d} /* (2, 3, 12) {real, imag} */,
  {32'hc0f4df02, 32'hbf72436f} /* (2, 3, 11) {real, imag} */,
  {32'h3f69f23c, 32'hbfff7294} /* (2, 3, 10) {real, imag} */,
  {32'h400e699e, 32'h3fb501de} /* (2, 3, 9) {real, imag} */,
  {32'hc0550052, 32'h40dbf4ec} /* (2, 3, 8) {real, imag} */,
  {32'hc0b175fe, 32'h4028f5eb} /* (2, 3, 7) {real, imag} */,
  {32'hc0d06a93, 32'h3f534870} /* (2, 3, 6) {real, imag} */,
  {32'hc120e63d, 32'h3ff4ddaf} /* (2, 3, 5) {real, imag} */,
  {32'hc0b40c22, 32'hc0126e76} /* (2, 3, 4) {real, imag} */,
  {32'hc011dc38, 32'h3fbc2148} /* (2, 3, 3) {real, imag} */,
  {32'h3fc974a4, 32'hc0092706} /* (2, 3, 2) {real, imag} */,
  {32'h3fdaa885, 32'hc0a7ed8c} /* (2, 3, 1) {real, imag} */,
  {32'hc0f79c5d, 32'hc0da488c} /* (2, 3, 0) {real, imag} */,
  {32'h40c86fb7, 32'hc085f157} /* (2, 2, 15) {real, imag} */,
  {32'h3ff69560, 32'hc154cf00} /* (2, 2, 14) {real, imag} */,
  {32'h40ff0268, 32'h402be188} /* (2, 2, 13) {real, imag} */,
  {32'h41a614cb, 32'h41425ddb} /* (2, 2, 12) {real, imag} */,
  {32'h40167198, 32'h409651ae} /* (2, 2, 11) {real, imag} */,
  {32'hc0f420b6, 32'h3edd49a0} /* (2, 2, 10) {real, imag} */,
  {32'hc112e76d, 32'hc0b39a38} /* (2, 2, 9) {real, imag} */,
  {32'hc059956a, 32'h3e26e6a0} /* (2, 2, 8) {real, imag} */,
  {32'h3fa99f34, 32'hc107bc72} /* (2, 2, 7) {real, imag} */,
  {32'hbffaa2a0, 32'hc09b100c} /* (2, 2, 6) {real, imag} */,
  {32'h40b16fc4, 32'h409c3c0e} /* (2, 2, 5) {real, imag} */,
  {32'h3f2f03e6, 32'hc0c655f2} /* (2, 2, 4) {real, imag} */,
  {32'h4081af97, 32'hc10fc3a4} /* (2, 2, 3) {real, imag} */,
  {32'hc0be89c6, 32'h4017c15a} /* (2, 2, 2) {real, imag} */,
  {32'hc0eb90d3, 32'h41079d9a} /* (2, 2, 1) {real, imag} */,
  {32'hc016eee0, 32'h4098d7be} /* (2, 2, 0) {real, imag} */,
  {32'h40012f0d, 32'h40a083a3} /* (2, 1, 15) {real, imag} */,
  {32'h40ebd6e4, 32'h416111e8} /* (2, 1, 14) {real, imag} */,
  {32'hbfdc2700, 32'h412db6fe} /* (2, 1, 13) {real, imag} */,
  {32'h4053dff2, 32'h3ffccc40} /* (2, 1, 12) {real, imag} */,
  {32'h407b98a6, 32'hc127d691} /* (2, 1, 11) {real, imag} */,
  {32'h41041e67, 32'hc08f3b26} /* (2, 1, 10) {real, imag} */,
  {32'h415cbc82, 32'h4174d5c2} /* (2, 1, 9) {real, imag} */,
  {32'h40748956, 32'h40e5a755} /* (2, 1, 8) {real, imag} */,
  {32'h40db76a5, 32'hc0aa330a} /* (2, 1, 7) {real, imag} */,
  {32'h410129a4, 32'hc0dce82c} /* (2, 1, 6) {real, imag} */,
  {32'h410b98c6, 32'hc0e8fcd6} /* (2, 1, 5) {real, imag} */,
  {32'hc017026e, 32'hc129cb49} /* (2, 1, 4) {real, imag} */,
  {32'hc137e89a, 32'hbfad55b8} /* (2, 1, 3) {real, imag} */,
  {32'hc095e15f, 32'h3fa8eac4} /* (2, 1, 2) {real, imag} */,
  {32'hc05bf431, 32'hc036163d} /* (2, 1, 1) {real, imag} */,
  {32'hc091ee38, 32'h3f21b1b4} /* (2, 1, 0) {real, imag} */,
  {32'h3eb685bc, 32'hbfb2c287} /* (2, 0, 15) {real, imag} */,
  {32'h4107f024, 32'hc02f72b8} /* (2, 0, 14) {real, imag} */,
  {32'h407bcc25, 32'hc1132d04} /* (2, 0, 13) {real, imag} */,
  {32'h40c43a5c, 32'hc1450e62} /* (2, 0, 12) {real, imag} */,
  {32'h406c2714, 32'hc1398d4a} /* (2, 0, 11) {real, imag} */,
  {32'h402a14f1, 32'hbfdd0063} /* (2, 0, 10) {real, imag} */,
  {32'h4040303c, 32'h400c3619} /* (2, 0, 9) {real, imag} */,
  {32'hbf52b970, 32'hc059e926} /* (2, 0, 8) {real, imag} */,
  {32'hc0e3d55d, 32'hc189d7fa} /* (2, 0, 7) {real, imag} */,
  {32'h40960446, 32'hc08f0c89} /* (2, 0, 6) {real, imag} */,
  {32'h401a5a8a, 32'hc01ed3c6} /* (2, 0, 5) {real, imag} */,
  {32'h4062034d, 32'hc1115963} /* (2, 0, 4) {real, imag} */,
  {32'hc003d271, 32'hbebe0998} /* (2, 0, 3) {real, imag} */,
  {32'h40b453d8, 32'h3e3c5230} /* (2, 0, 2) {real, imag} */,
  {32'h40dcfb57, 32'hc14c6ad0} /* (2, 0, 1) {real, imag} */,
  {32'h3ffdef8a, 32'hc1263e29} /* (2, 0, 0) {real, imag} */,
  {32'hbf90ed9a, 32'h40fb6273} /* (1, 15, 15) {real, imag} */,
  {32'h400032fe, 32'hbe2d60a0} /* (1, 15, 14) {real, imag} */,
  {32'h3f40c410, 32'hbea217dc} /* (1, 15, 13) {real, imag} */,
  {32'hc06e2d08, 32'hc0b42c75} /* (1, 15, 12) {real, imag} */,
  {32'h4095859b, 32'hc0f1fac7} /* (1, 15, 11) {real, imag} */,
  {32'hc00eac82, 32'h411d97cc} /* (1, 15, 10) {real, imag} */,
  {32'h40bfcb0a, 32'h40d7a734} /* (1, 15, 9) {real, imag} */,
  {32'h404c61b0, 32'h3fd17280} /* (1, 15, 8) {real, imag} */,
  {32'hbf643104, 32'h4050775c} /* (1, 15, 7) {real, imag} */,
  {32'hc035aac4, 32'hc0f5e216} /* (1, 15, 6) {real, imag} */,
  {32'hbfd53d36, 32'hc130994c} /* (1, 15, 5) {real, imag} */,
  {32'hc0e243fa, 32'h3f22b428} /* (1, 15, 4) {real, imag} */,
  {32'hc15f7deb, 32'h40b0ee74} /* (1, 15, 3) {real, imag} */,
  {32'hbff9aed8, 32'h3fa69438} /* (1, 15, 2) {real, imag} */,
  {32'h4039c151, 32'h40e2680b} /* (1, 15, 1) {real, imag} */,
  {32'hc0920942, 32'h40c13ada} /* (1, 15, 0) {real, imag} */,
  {32'hbff07d3b, 32'hc04c3c93} /* (1, 14, 15) {real, imag} */,
  {32'h40ccde6a, 32'h4030d138} /* (1, 14, 14) {real, imag} */,
  {32'h400b4224, 32'h4137ed30} /* (1, 14, 13) {real, imag} */,
  {32'hc01f21e9, 32'h41542abc} /* (1, 14, 12) {real, imag} */,
  {32'h3fa9609f, 32'h412c8186} /* (1, 14, 11) {real, imag} */,
  {32'hc0879099, 32'h3edd1040} /* (1, 14, 10) {real, imag} */,
  {32'h40db19bc, 32'hc0e97613} /* (1, 14, 9) {real, imag} */,
  {32'hc139f26a, 32'hc10664aa} /* (1, 14, 8) {real, imag} */,
  {32'hc0545a14, 32'hc11b29b0} /* (1, 14, 7) {real, imag} */,
  {32'h4127bb8b, 32'hc0d10e4b} /* (1, 14, 6) {real, imag} */,
  {32'h41946c88, 32'hc0473d50} /* (1, 14, 5) {real, imag} */,
  {32'h4135a7fe, 32'hc166f47a} /* (1, 14, 4) {real, imag} */,
  {32'h3f9adfe0, 32'hc150fc08} /* (1, 14, 3) {real, imag} */,
  {32'h3eb4e110, 32'hc05d9740} /* (1, 14, 2) {real, imag} */,
  {32'hc1519fee, 32'hc105896b} /* (1, 14, 1) {real, imag} */,
  {32'hc0e6bdfa, 32'hc03438f6} /* (1, 14, 0) {real, imag} */,
  {32'hbec61428, 32'h3faeaef1} /* (1, 13, 15) {real, imag} */,
  {32'h40454f34, 32'h40a42db6} /* (1, 13, 14) {real, imag} */,
  {32'h40dad4ce, 32'h408b3cfe} /* (1, 13, 13) {real, imag} */,
  {32'h40e68e6a, 32'h402d5360} /* (1, 13, 12) {real, imag} */,
  {32'hc09d4644, 32'hbf0a4452} /* (1, 13, 11) {real, imag} */,
  {32'hc1821158, 32'hc0abc744} /* (1, 13, 10) {real, imag} */,
  {32'hc170e040, 32'h41142b72} /* (1, 13, 9) {real, imag} */,
  {32'hc0caef89, 32'h4001812e} /* (1, 13, 8) {real, imag} */,
  {32'h3fbe561a, 32'h40221096} /* (1, 13, 7) {real, imag} */,
  {32'h40b0b626, 32'hbf0d2744} /* (1, 13, 6) {real, imag} */,
  {32'hbfc37fce, 32'h411a1638} /* (1, 13, 5) {real, imag} */,
  {32'hc13c623e, 32'h3decfe80} /* (1, 13, 4) {real, imag} */,
  {32'hbf838c70, 32'h3e97ff90} /* (1, 13, 3) {real, imag} */,
  {32'h4069ae23, 32'h403e13fe} /* (1, 13, 2) {real, imag} */,
  {32'h4078e706, 32'h408f9950} /* (1, 13, 1) {real, imag} */,
  {32'hc016fc74, 32'h40de8a57} /* (1, 13, 0) {real, imag} */,
  {32'hc0baa896, 32'h3ffe7b1d} /* (1, 12, 15) {real, imag} */,
  {32'hc11d1882, 32'hc0bd4b31} /* (1, 12, 14) {real, imag} */,
  {32'hc084e747, 32'hc12df8aa} /* (1, 12, 13) {real, imag} */,
  {32'h402c26e8, 32'hc012f92b} /* (1, 12, 12) {real, imag} */,
  {32'hc081fc6a, 32'hbd2c3f80} /* (1, 12, 11) {real, imag} */,
  {32'hc0bf1001, 32'hbf9b46f2} /* (1, 12, 10) {real, imag} */,
  {32'hc0d5be20, 32'hc0e70662} /* (1, 12, 9) {real, imag} */,
  {32'hbf2b8e50, 32'hc067bd0d} /* (1, 12, 8) {real, imag} */,
  {32'hc0495f08, 32'hc1066386} /* (1, 12, 7) {real, imag} */,
  {32'h4087040e, 32'hc0b9f0db} /* (1, 12, 6) {real, imag} */,
  {32'h40e33929, 32'hc0e465ca} /* (1, 12, 5) {real, imag} */,
  {32'h40575db2, 32'hc0c3a763} /* (1, 12, 4) {real, imag} */,
  {32'h410ee522, 32'h3f9a3c97} /* (1, 12, 3) {real, imag} */,
  {32'h4116d3b4, 32'h401fcf5b} /* (1, 12, 2) {real, imag} */,
  {32'h4086c73b, 32'h40d6957e} /* (1, 12, 1) {real, imag} */,
  {32'hc08cd836, 32'h4083fb8c} /* (1, 12, 0) {real, imag} */,
  {32'h408f18bb, 32'hc072591a} /* (1, 11, 15) {real, imag} */,
  {32'hbe8c4fe4, 32'hc0870d43} /* (1, 11, 14) {real, imag} */,
  {32'hc09274ce, 32'hc0854222} /* (1, 11, 13) {real, imag} */,
  {32'h3fc54b10, 32'hbfeeb67c} /* (1, 11, 12) {real, imag} */,
  {32'hbeabb9a0, 32'h40416ff4} /* (1, 11, 11) {real, imag} */,
  {32'h3f4bdf94, 32'hbf877154} /* (1, 11, 10) {real, imag} */,
  {32'hc05458bc, 32'h3ed0a8e0} /* (1, 11, 9) {real, imag} */,
  {32'hc114e906, 32'h40d655e1} /* (1, 11, 8) {real, imag} */,
  {32'hc09edaaa, 32'h4056452c} /* (1, 11, 7) {real, imag} */,
  {32'hbf0bd8a0, 32'h403c9b47} /* (1, 11, 6) {real, imag} */,
  {32'h3fc0dd7e, 32'h3c12f800} /* (1, 11, 5) {real, imag} */,
  {32'hbe017030, 32'hbfc35d14} /* (1, 11, 4) {real, imag} */,
  {32'h3dea6340, 32'hbfbf6fe6} /* (1, 11, 3) {real, imag} */,
  {32'hc0a7115a, 32'hbf2f970c} /* (1, 11, 2) {real, imag} */,
  {32'hc0577399, 32'h3fbf4762} /* (1, 11, 1) {real, imag} */,
  {32'h40ac9b24, 32'h40019e50} /* (1, 11, 0) {real, imag} */,
  {32'h401e6c25, 32'hc0a60dda} /* (1, 10, 15) {real, imag} */,
  {32'h4093da05, 32'hc0504429} /* (1, 10, 14) {real, imag} */,
  {32'hbee8ad48, 32'h40a4b6cb} /* (1, 10, 13) {real, imag} */,
  {32'hbfad2f4f, 32'h3f81d1f6} /* (1, 10, 12) {real, imag} */,
  {32'h3f96619c, 32'hc022dccb} /* (1, 10, 11) {real, imag} */,
  {32'hbfa714b8, 32'h40274d58} /* (1, 10, 10) {real, imag} */,
  {32'hbfb1a319, 32'h40a773d6} /* (1, 10, 9) {real, imag} */,
  {32'hbfae7fcb, 32'h3fce2330} /* (1, 10, 8) {real, imag} */,
  {32'hc0479cb2, 32'h3f9e450b} /* (1, 10, 7) {real, imag} */,
  {32'hbf838596, 32'h3ec1c598} /* (1, 10, 6) {real, imag} */,
  {32'hbfeda80e, 32'h3f137c8b} /* (1, 10, 5) {real, imag} */,
  {32'h40c452e5, 32'hbda59920} /* (1, 10, 4) {real, imag} */,
  {32'h406b1bd8, 32'hbf9b2bb5} /* (1, 10, 3) {real, imag} */,
  {32'h3fe6ec88, 32'h3f8be511} /* (1, 10, 2) {real, imag} */,
  {32'h40210af4, 32'hc00e3e34} /* (1, 10, 1) {real, imag} */,
  {32'h3f8be298, 32'hc08c614c} /* (1, 10, 0) {real, imag} */,
  {32'hbf812fb0, 32'h3f260418} /* (1, 9, 15) {real, imag} */,
  {32'h3ff32a0f, 32'hbf34994e} /* (1, 9, 14) {real, imag} */,
  {32'h406907f4, 32'hc0318187} /* (1, 9, 13) {real, imag} */,
  {32'h3e33802c, 32'h3e5f8964} /* (1, 9, 12) {real, imag} */,
  {32'h3f01f8ad, 32'h3fee83e1} /* (1, 9, 11) {real, imag} */,
  {32'h3f05f7f0, 32'h3fc32ed2} /* (1, 9, 10) {real, imag} */,
  {32'hbd1e8200, 32'hbffedf6c} /* (1, 9, 9) {real, imag} */,
  {32'h3f1519f2, 32'hc0b8e6ee} /* (1, 9, 8) {real, imag} */,
  {32'hbefdf1d2, 32'hc08f6a19} /* (1, 9, 7) {real, imag} */,
  {32'hbef353d2, 32'h3f8fc3a2} /* (1, 9, 6) {real, imag} */,
  {32'hbf25f2f4, 32'hbf57f936} /* (1, 9, 5) {real, imag} */,
  {32'h3f5e7b20, 32'hbf029d4c} /* (1, 9, 4) {real, imag} */,
  {32'hbf1d5f70, 32'h3fa1910b} /* (1, 9, 3) {real, imag} */,
  {32'h40141013, 32'h3fff36ce} /* (1, 9, 2) {real, imag} */,
  {32'h4089f9f4, 32'h3f89f9c3} /* (1, 9, 1) {real, imag} */,
  {32'h400b4622, 32'hbf98b69c} /* (1, 9, 0) {real, imag} */,
  {32'hbe912a88, 32'hbe7383a0} /* (1, 8, 15) {real, imag} */,
  {32'h3ff1b44a, 32'hbdff4e80} /* (1, 8, 14) {real, imag} */,
  {32'hbfc52204, 32'h400c29c3} /* (1, 8, 13) {real, imag} */,
  {32'h3e33af00, 32'h3f7495f4} /* (1, 8, 12) {real, imag} */,
  {32'h3efa4f38, 32'hbff412ee} /* (1, 8, 11) {real, imag} */,
  {32'h400a2426, 32'h3d9d4cf0} /* (1, 8, 10) {real, imag} */,
  {32'hbefe2a68, 32'h3fc138f1} /* (1, 8, 9) {real, imag} */,
  {32'hc04dad22, 32'h3ff15a9a} /* (1, 8, 8) {real, imag} */,
  {32'h3d32ec60, 32'h404be960} /* (1, 8, 7) {real, imag} */,
  {32'hbd665d00, 32'hbf9744d1} /* (1, 8, 6) {real, imag} */,
  {32'hbf738500, 32'hc050d6fe} /* (1, 8, 5) {real, imag} */,
  {32'h3e3c9c80, 32'hc032b2b4} /* (1, 8, 4) {real, imag} */,
  {32'h3d2863e0, 32'hbdc6dd80} /* (1, 8, 3) {real, imag} */,
  {32'hbf9c2a26, 32'hbf82a31a} /* (1, 8, 2) {real, imag} */,
  {32'hc00a7ee6, 32'hbf5c7a94} /* (1, 8, 1) {real, imag} */,
  {32'hc01c9c11, 32'hbf1ed806} /* (1, 8, 0) {real, imag} */,
  {32'h3e9fc232, 32'h3ff1b38c} /* (1, 7, 15) {real, imag} */,
  {32'hbea5f56c, 32'hbf285bb6} /* (1, 7, 14) {real, imag} */,
  {32'hbe007788, 32'hc0063dd5} /* (1, 7, 13) {real, imag} */,
  {32'h3f90025e, 32'h400b0f46} /* (1, 7, 12) {real, imag} */,
  {32'hbf2d3a73, 32'h3ffc3a3f} /* (1, 7, 11) {real, imag} */,
  {32'hbf41a620, 32'h401306c9} /* (1, 7, 10) {real, imag} */,
  {32'hbd5c4a80, 32'hbfe09638} /* (1, 7, 9) {real, imag} */,
  {32'h3ed4a2fc, 32'h3ebbc380} /* (1, 7, 8) {real, imag} */,
  {32'h3d9faa98, 32'h40230b72} /* (1, 7, 7) {real, imag} */,
  {32'h3f9f2baa, 32'h3e814f6a} /* (1, 7, 6) {real, imag} */,
  {32'h401d0ceb, 32'h3f347f5a} /* (1, 7, 5) {real, imag} */,
  {32'h40665e9a, 32'hbe8a15c8} /* (1, 7, 4) {real, imag} */,
  {32'h3fa15db0, 32'h3f4f9f92} /* (1, 7, 3) {real, imag} */,
  {32'hbf1fed2c, 32'hbf59289c} /* (1, 7, 2) {real, imag} */,
  {32'h4003f557, 32'hc04cca58} /* (1, 7, 1) {real, imag} */,
  {32'h3eeea5d0, 32'hbef3cbf0} /* (1, 7, 0) {real, imag} */,
  {32'hbf8a2858, 32'hbf519eb0} /* (1, 6, 15) {real, imag} */,
  {32'hbf010630, 32'h408154f2} /* (1, 6, 14) {real, imag} */,
  {32'h4043476b, 32'h40a9fedb} /* (1, 6, 13) {real, imag} */,
  {32'h40a8ec3b, 32'hc06e8a3f} /* (1, 6, 12) {real, imag} */,
  {32'h4052e8a6, 32'hbf22716c} /* (1, 6, 11) {real, imag} */,
  {32'hbe7a3df4, 32'h3fbfc4cc} /* (1, 6, 10) {real, imag} */,
  {32'h405d8756, 32'h4065f75c} /* (1, 6, 9) {real, imag} */,
  {32'h40536c28, 32'h400b021a} /* (1, 6, 8) {real, imag} */,
  {32'h3f4ac536, 32'hc01c6fd8} /* (1, 6, 7) {real, imag} */,
  {32'hbef265d8, 32'hc069776d} /* (1, 6, 6) {real, imag} */,
  {32'hc02cbb53, 32'h3f8a00fe} /* (1, 6, 5) {real, imag} */,
  {32'h4088b2b3, 32'hbf40b354} /* (1, 6, 4) {real, imag} */,
  {32'h409cb9ae, 32'hc022d9f0} /* (1, 6, 3) {real, imag} */,
  {32'hbec7b7d0, 32'hbf9188f5} /* (1, 6, 2) {real, imag} */,
  {32'hc0699be6, 32'h3f4adb8e} /* (1, 6, 1) {real, imag} */,
  {32'hba11c000, 32'hbf99f883} /* (1, 6, 0) {real, imag} */,
  {32'h3f0f2c22, 32'h3f9b9697} /* (1, 5, 15) {real, imag} */,
  {32'h3fb734cd, 32'h40c66555} /* (1, 5, 14) {real, imag} */,
  {32'h3f9ae81e, 32'h40b18da4} /* (1, 5, 13) {real, imag} */,
  {32'hc00315a0, 32'h40d17ac7} /* (1, 5, 12) {real, imag} */,
  {32'hc02c6458, 32'hc02bd80a} /* (1, 5, 11) {real, imag} */,
  {32'hc0a16374, 32'hbf900df4} /* (1, 5, 10) {real, imag} */,
  {32'hc02f92cc, 32'h3f7b7890} /* (1, 5, 9) {real, imag} */,
  {32'h3f3c6388, 32'hbf3a74c8} /* (1, 5, 8) {real, imag} */,
  {32'h40adf6dc, 32'h40c8e8f2} /* (1, 5, 7) {real, imag} */,
  {32'h408b5d72, 32'h4111ed84} /* (1, 5, 6) {real, imag} */,
  {32'hbf21392c, 32'h40d534e3} /* (1, 5, 5) {real, imag} */,
  {32'hbfb4843a, 32'h40cbbbe7} /* (1, 5, 4) {real, imag} */,
  {32'hbf9ae63c, 32'h40e55006} /* (1, 5, 3) {real, imag} */,
  {32'hc07c9163, 32'hbf402c5a} /* (1, 5, 2) {real, imag} */,
  {32'hc0205409, 32'hc03524e7} /* (1, 5, 1) {real, imag} */,
  {32'hbfc0bca6, 32'h4030f520} /* (1, 5, 0) {real, imag} */,
  {32'h3fee11af, 32'hc0378732} /* (1, 4, 15) {real, imag} */,
  {32'h40ba0014, 32'hc0728696} /* (1, 4, 14) {real, imag} */,
  {32'h3feab27c, 32'hc05cbb86} /* (1, 4, 13) {real, imag} */,
  {32'hc0c6f970, 32'hbfe6d0d2} /* (1, 4, 12) {real, imag} */,
  {32'hc0b7e1b6, 32'hbf485190} /* (1, 4, 11) {real, imag} */,
  {32'hbfcd25b4, 32'hc05c19ff} /* (1, 4, 10) {real, imag} */,
  {32'hbfb6f250, 32'h403b9d61} /* (1, 4, 9) {real, imag} */,
  {32'hc0c9b726, 32'h40d36d04} /* (1, 4, 8) {real, imag} */,
  {32'hc1028096, 32'hc095903a} /* (1, 4, 7) {real, imag} */,
  {32'hc0488df4, 32'hc0ebe22b} /* (1, 4, 6) {real, imag} */,
  {32'h40880707, 32'hc0cfca54} /* (1, 4, 5) {real, imag} */,
  {32'h3f0fe1a8, 32'h40a34855} /* (1, 4, 4) {real, imag} */,
  {32'h3e93cec0, 32'hc02b8902} /* (1, 4, 3) {real, imag} */,
  {32'h41085e34, 32'hc0ae6f62} /* (1, 4, 2) {real, imag} */,
  {32'h40ae89ff, 32'hbf3abf84} /* (1, 4, 1) {real, imag} */,
  {32'hbf8b3d4b, 32'hbe6f6ca0} /* (1, 4, 0) {real, imag} */,
  {32'hc0a18550, 32'h40088712} /* (1, 3, 15) {real, imag} */,
  {32'hc04a1150, 32'hbfe4405a} /* (1, 3, 14) {real, imag} */,
  {32'hbfd6114e, 32'hc0fd07bc} /* (1, 3, 13) {real, imag} */,
  {32'h4036d7d4, 32'hbe30d400} /* (1, 3, 12) {real, imag} */,
  {32'h411dafab, 32'h407e9736} /* (1, 3, 11) {real, imag} */,
  {32'h4105e3c8, 32'h40c138be} /* (1, 3, 10) {real, imag} */,
  {32'h40e34e38, 32'h40236ee2} /* (1, 3, 9) {real, imag} */,
  {32'h40d8b3e1, 32'h405165ca} /* (1, 3, 8) {real, imag} */,
  {32'hbf9b85cc, 32'h4119150a} /* (1, 3, 7) {real, imag} */,
  {32'hbff8c8ee, 32'h400ea7e1} /* (1, 3, 6) {real, imag} */,
  {32'hc00b10fd, 32'hc0949f88} /* (1, 3, 5) {real, imag} */,
  {32'hc12837a2, 32'h3fd8d9ea} /* (1, 3, 4) {real, imag} */,
  {32'hc16001bd, 32'h407ec468} /* (1, 3, 3) {real, imag} */,
  {32'hc0bf0fee, 32'h40061128} /* (1, 3, 2) {real, imag} */,
  {32'h40a21c7f, 32'hc09df68a} /* (1, 3, 1) {real, imag} */,
  {32'hc0415242, 32'h3e9df210} /* (1, 3, 0) {real, imag} */,
  {32'hbfc665b9, 32'hc0a2bbc8} /* (1, 2, 15) {real, imag} */,
  {32'hc054ea5b, 32'hc144090e} /* (1, 2, 14) {real, imag} */,
  {32'hc09fd2e0, 32'hc112f1bc} /* (1, 2, 13) {real, imag} */,
  {32'hc03e690f, 32'hc0db615d} /* (1, 2, 12) {real, imag} */,
  {32'hc016f80c, 32'h407d4d9a} /* (1, 2, 11) {real, imag} */,
  {32'h3f4d550e, 32'hbf1cf0d6} /* (1, 2, 10) {real, imag} */,
  {32'h4008a175, 32'hc0ee0f39} /* (1, 2, 9) {real, imag} */,
  {32'h40b968f9, 32'h3fe0ef3e} /* (1, 2, 8) {real, imag} */,
  {32'h3ea712fc, 32'hbf124818} /* (1, 2, 7) {real, imag} */,
  {32'h3f482a70, 32'hc0fd331d} /* (1, 2, 6) {real, imag} */,
  {32'hc0a1c2e2, 32'hc0dff288} /* (1, 2, 5) {real, imag} */,
  {32'hc0086946, 32'h3fc1d89c} /* (1, 2, 4) {real, imag} */,
  {32'hc028a500, 32'h3fc70f04} /* (1, 2, 3) {real, imag} */,
  {32'hc05eed10, 32'h40b15d74} /* (1, 2, 2) {real, imag} */,
  {32'h3f99f580, 32'h409f8541} /* (1, 2, 1) {real, imag} */,
  {32'h4082ce30, 32'hbff4c59f} /* (1, 2, 0) {real, imag} */,
  {32'h4022ddbb, 32'h415a51ce} /* (1, 1, 15) {real, imag} */,
  {32'hbfed6999, 32'h4098c435} /* (1, 1, 14) {real, imag} */,
  {32'h4072d7e0, 32'hbe0cab98} /* (1, 1, 13) {real, imag} */,
  {32'h4078a7bc, 32'hc08c66ed} /* (1, 1, 12) {real, imag} */,
  {32'hc0a9172d, 32'hc0b4d249} /* (1, 1, 11) {real, imag} */,
  {32'hc1117fc8, 32'hc0b596d4} /* (1, 1, 10) {real, imag} */,
  {32'hc06b997b, 32'hc0ef9a80} /* (1, 1, 9) {real, imag} */,
  {32'h41061487, 32'hc0f77d56} /* (1, 1, 8) {real, imag} */,
  {32'h405664e7, 32'hc0b318a6} /* (1, 1, 7) {real, imag} */,
  {32'hbdb3e790, 32'h40f0005c} /* (1, 1, 6) {real, imag} */,
  {32'hc0036953, 32'h412184c4} /* (1, 1, 5) {real, imag} */,
  {32'hc053c8ab, 32'h41112ef0} /* (1, 1, 4) {real, imag} */,
  {32'h412721d9, 32'hbff13a06} /* (1, 1, 3) {real, imag} */,
  {32'h41252939, 32'hc134ce67} /* (1, 1, 2) {real, imag} */,
  {32'hbfe300aa, 32'hc0b2345d} /* (1, 1, 1) {real, imag} */,
  {32'hc04ffc67, 32'h40140e00} /* (1, 1, 0) {real, imag} */,
  {32'hbfbaaf54, 32'h40de9a29} /* (1, 0, 15) {real, imag} */,
  {32'hc1193de5, 32'h410fbf6b} /* (1, 0, 14) {real, imag} */,
  {32'h406fe0e2, 32'hbfe6aada} /* (1, 0, 13) {real, imag} */,
  {32'h41585c6c, 32'h40a5e49e} /* (1, 0, 12) {real, imag} */,
  {32'h40df48fe, 32'h40ed6e02} /* (1, 0, 11) {real, imag} */,
  {32'h41476c78, 32'hc00acd20} /* (1, 0, 10) {real, imag} */,
  {32'hc103f713, 32'h4098eaa1} /* (1, 0, 9) {real, imag} */,
  {32'h404fe66a, 32'hbe0f4270} /* (1, 0, 8) {real, imag} */,
  {32'hbfb3c773, 32'h411e1d8d} /* (1, 0, 7) {real, imag} */,
  {32'hc1929d0a, 32'hc091f8ca} /* (1, 0, 6) {real, imag} */,
  {32'hc1a86718, 32'hc1853068} /* (1, 0, 5) {real, imag} */,
  {32'hc11a16ae, 32'h40c68c86} /* (1, 0, 4) {real, imag} */,
  {32'h3f27f4aa, 32'h412985ad} /* (1, 0, 3) {real, imag} */,
  {32'hbf93a9fe, 32'h410ee227} /* (1, 0, 2) {real, imag} */,
  {32'h401330fa, 32'h409681c2} /* (1, 0, 1) {real, imag} */,
  {32'h40fef530, 32'hbf2deb12} /* (1, 0, 0) {real, imag} */,
  {32'hc1179cce, 32'hc1192ea6} /* (0, 15, 15) {real, imag} */,
  {32'hc10525d1, 32'hc007e0cc} /* (0, 15, 14) {real, imag} */,
  {32'h4114de86, 32'h404f3fae} /* (0, 15, 13) {real, imag} */,
  {32'h4135b108, 32'h404b8542} /* (0, 15, 12) {real, imag} */,
  {32'h40441b1e, 32'h3f7f82d0} /* (0, 15, 11) {real, imag} */,
  {32'hc0ef881b, 32'h3fd55420} /* (0, 15, 10) {real, imag} */,
  {32'hc119c0cc, 32'h40503ba2} /* (0, 15, 9) {real, imag} */,
  {32'h3faa63d3, 32'h3f44b196} /* (0, 15, 8) {real, imag} */,
  {32'hc074c589, 32'h40656154} /* (0, 15, 7) {real, imag} */,
  {32'h406556ec, 32'h3cfae680} /* (0, 15, 6) {real, imag} */,
  {32'h3fa74678, 32'hc12f0ba2} /* (0, 15, 5) {real, imag} */,
  {32'hc05324c0, 32'hc0976cf7} /* (0, 15, 4) {real, imag} */,
  {32'hc06c9129, 32'h3f21ffb0} /* (0, 15, 3) {real, imag} */,
  {32'hc0604eb8, 32'hc00cdd05} /* (0, 15, 2) {real, imag} */,
  {32'hc105f002, 32'hc12e8e28} /* (0, 15, 1) {real, imag} */,
  {32'hbfe827fc, 32'hbf9358e6} /* (0, 15, 0) {real, imag} */,
  {32'h40caf222, 32'hc07ac38a} /* (0, 14, 15) {real, imag} */,
  {32'h3f24454e, 32'h3fcb4933} /* (0, 14, 14) {real, imag} */,
  {32'hbf754160, 32'h4148e68c} /* (0, 14, 13) {real, imag} */,
  {32'hbea25e3c, 32'h410160f0} /* (0, 14, 12) {real, imag} */,
  {32'h40852f00, 32'h40723f55} /* (0, 14, 11) {real, imag} */,
  {32'h40f85ce5, 32'h40b1400a} /* (0, 14, 10) {real, imag} */,
  {32'hc00062d5, 32'h4046397a} /* (0, 14, 9) {real, imag} */,
  {32'hc0679195, 32'h40a7d6fa} /* (0, 14, 8) {real, imag} */,
  {32'h3fc5ed6e, 32'hbfeb82c6} /* (0, 14, 7) {real, imag} */,
  {32'hc1087f7c, 32'hc15183c0} /* (0, 14, 6) {real, imag} */,
  {32'hc08d1551, 32'hc081b5a7} /* (0, 14, 5) {real, imag} */,
  {32'hbfa13dbb, 32'h40cc7a2a} /* (0, 14, 4) {real, imag} */,
  {32'hbfa92ce6, 32'h4113ebdc} /* (0, 14, 3) {real, imag} */,
  {32'h40301323, 32'h4123ff6c} /* (0, 14, 2) {real, imag} */,
  {32'hc04a6654, 32'h406e976a} /* (0, 14, 1) {real, imag} */,
  {32'hc011bcdd, 32'hc048b1f2} /* (0, 14, 0) {real, imag} */,
  {32'hc03f2a0e, 32'hc0ac4b1f} /* (0, 13, 15) {real, imag} */,
  {32'hbfb616db, 32'hc0e137aa} /* (0, 13, 14) {real, imag} */,
  {32'h40395ab0, 32'h407693ca} /* (0, 13, 13) {real, imag} */,
  {32'h408029a8, 32'h3f7ef4f7} /* (0, 13, 12) {real, imag} */,
  {32'hc1131358, 32'hc1375593} /* (0, 13, 11) {real, imag} */,
  {32'hbfcb762e, 32'hbfb1a563} /* (0, 13, 10) {real, imag} */,
  {32'h4149db08, 32'h41166e48} /* (0, 13, 9) {real, imag} */,
  {32'h406a4f8a, 32'h4028f29a} /* (0, 13, 8) {real, imag} */,
  {32'hc03a146c, 32'hc08fa502} /* (0, 13, 7) {real, imag} */,
  {32'h40847dd1, 32'hc066f01e} /* (0, 13, 6) {real, imag} */,
  {32'h410c470b, 32'hc021a26f} /* (0, 13, 5) {real, imag} */,
  {32'h4191be20, 32'hc029b599} /* (0, 13, 4) {real, imag} */,
  {32'h40d3030d, 32'hc05d8fa2} /* (0, 13, 3) {real, imag} */,
  {32'h40384162, 32'hc12c3c58} /* (0, 13, 2) {real, imag} */,
  {32'h3fa9db5c, 32'hc14a2c0e} /* (0, 13, 1) {real, imag} */,
  {32'hc02170ac, 32'hc0583e5a} /* (0, 13, 0) {real, imag} */,
  {32'h3e2814d8, 32'h3e56696e} /* (0, 12, 15) {real, imag} */,
  {32'h40f7a888, 32'hc069c41f} /* (0, 12, 14) {real, imag} */,
  {32'h41046632, 32'hc085b8c8} /* (0, 12, 13) {real, imag} */,
  {32'hbfcc3dba, 32'hbe7cbaa8} /* (0, 12, 12) {real, imag} */,
  {32'hc10e2f1e, 32'hc0481fdc} /* (0, 12, 11) {real, imag} */,
  {32'h401984a8, 32'h4076436c} /* (0, 12, 10) {real, imag} */,
  {32'h404da213, 32'h40715eae} /* (0, 12, 9) {real, imag} */,
  {32'h3fc9e304, 32'h3f9e8504} /* (0, 12, 8) {real, imag} */,
  {32'hc1040d3f, 32'h409f88b5} /* (0, 12, 7) {real, imag} */,
  {32'hc10f63b6, 32'h4117bb64} /* (0, 12, 6) {real, imag} */,
  {32'h404a9b76, 32'h40b62dc5} /* (0, 12, 5) {real, imag} */,
  {32'h40282a73, 32'h41148010} /* (0, 12, 4) {real, imag} */,
  {32'h403eaa2b, 32'hbfd15d4f} /* (0, 12, 3) {real, imag} */,
  {32'h412cc449, 32'hc0184ad4} /* (0, 12, 2) {real, imag} */,
  {32'h410f639e, 32'h40aa2431} /* (0, 12, 1) {real, imag} */,
  {32'hbf852964, 32'h405e91e2} /* (0, 12, 0) {real, imag} */,
  {32'hc0829223, 32'h3fc2f4d4} /* (0, 11, 15) {real, imag} */,
  {32'hc02b77e2, 32'h407d28b7} /* (0, 11, 14) {real, imag} */,
  {32'hbe8d7bc4, 32'hbdcbc010} /* (0, 11, 13) {real, imag} */,
  {32'h407f5485, 32'hbf31621f} /* (0, 11, 12) {real, imag} */,
  {32'h404af058, 32'hc07b06b3} /* (0, 11, 11) {real, imag} */,
  {32'h40a4700c, 32'hc00c4068} /* (0, 11, 10) {real, imag} */,
  {32'h40896b8c, 32'h40856786} /* (0, 11, 9) {real, imag} */,
  {32'h40afdacd, 32'h40b3afe7} /* (0, 11, 8) {real, imag} */,
  {32'hbfb195f8, 32'hbfb75209} /* (0, 11, 7) {real, imag} */,
  {32'hbfbbcded, 32'h4055ce06} /* (0, 11, 6) {real, imag} */,
  {32'hc0757cbd, 32'h405f533d} /* (0, 11, 5) {real, imag} */,
  {32'hc0480b00, 32'h40cc0f96} /* (0, 11, 4) {real, imag} */,
  {32'h40a2a443, 32'h408a5065} /* (0, 11, 3) {real, imag} */,
  {32'h40da5c33, 32'h40439358} /* (0, 11, 2) {real, imag} */,
  {32'h408d1c63, 32'hc0253cca} /* (0, 11, 1) {real, imag} */,
  {32'h4082c02b, 32'hc012089a} /* (0, 11, 0) {real, imag} */,
  {32'h4000fa34, 32'h3fa465bc} /* (0, 10, 15) {real, imag} */,
  {32'h4053fcdc, 32'h3f13530e} /* (0, 10, 14) {real, imag} */,
  {32'h3eaffe90, 32'h40732c86} /* (0, 10, 13) {real, imag} */,
  {32'hc0087a8e, 32'h403132f4} /* (0, 10, 12) {real, imag} */,
  {32'h3f941408, 32'h407b0e17} /* (0, 10, 11) {real, imag} */,
  {32'hbfe5d0cc, 32'h3f255d50} /* (0, 10, 10) {real, imag} */,
  {32'h3f9af3dc, 32'h4010ae94} /* (0, 10, 9) {real, imag} */,
  {32'h4088a8c1, 32'hbda88da0} /* (0, 10, 8) {real, imag} */,
  {32'h406d6be9, 32'hc04df157} /* (0, 10, 7) {real, imag} */,
  {32'h40767bd5, 32'hc04fc058} /* (0, 10, 6) {real, imag} */,
  {32'h405efdf1, 32'h403d5027} /* (0, 10, 5) {real, imag} */,
  {32'h3f93ae9b, 32'hbfebbbe8} /* (0, 10, 4) {real, imag} */,
  {32'hbfc8edc6, 32'hc087295c} /* (0, 10, 3) {real, imag} */,
  {32'h3f721429, 32'hc0df3f77} /* (0, 10, 2) {real, imag} */,
  {32'h3f2753d0, 32'hbefd5ac0} /* (0, 10, 1) {real, imag} */,
  {32'h3fbd8c3c, 32'h40439446} /* (0, 10, 0) {real, imag} */,
  {32'h3ec93ee0, 32'hbec7a7f0} /* (0, 9, 15) {real, imag} */,
  {32'h3dea4e80, 32'h3db93010} /* (0, 9, 14) {real, imag} */,
  {32'hbee76b10, 32'h3f81014c} /* (0, 9, 13) {real, imag} */,
  {32'hbf8edf14, 32'h3f5e9c98} /* (0, 9, 12) {real, imag} */,
  {32'hbeac7350, 32'h3ec86970} /* (0, 9, 11) {real, imag} */,
  {32'hc056af4a, 32'hbfba0006} /* (0, 9, 10) {real, imag} */,
  {32'hc09ffee5, 32'h3f2af71a} /* (0, 9, 9) {real, imag} */,
  {32'h3ec6214c, 32'hbe54624a} /* (0, 9, 8) {real, imag} */,
  {32'h3f7fa84c, 32'hbf7c0938} /* (0, 9, 7) {real, imag} */,
  {32'hbfc28e07, 32'hbf9d9e28} /* (0, 9, 6) {real, imag} */,
  {32'hbf28ecf7, 32'hbff47c40} /* (0, 9, 5) {real, imag} */,
  {32'h3f5f7740, 32'hbfcd2284} /* (0, 9, 4) {real, imag} */,
  {32'h408223ca, 32'h3f9a0662} /* (0, 9, 3) {real, imag} */,
  {32'h409b2164, 32'h407367c9} /* (0, 9, 2) {real, imag} */,
  {32'h402a554e, 32'h3fc7732c} /* (0, 9, 1) {real, imag} */,
  {32'h3fdc4516, 32'h3df52020} /* (0, 9, 0) {real, imag} */,
  {32'h401011bf, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'h3e039b50, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'hbf8a3b60, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'hbf89e5ae, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'hc04a6cfe, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'hc065bb68, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hc056fd17, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'hbfe84126, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hbfbf8998, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hbf4f5ca8, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'h3f830bac, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'h3fa255e6, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'hc060158c, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'hc0f59916, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'hc06f7b34, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'h3e587f80, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h3ec93ee0, 32'h3ec7a7f0} /* (0, 7, 15) {real, imag} */,
  {32'h3dea4e80, 32'hbdb93010} /* (0, 7, 14) {real, imag} */,
  {32'hbee76b10, 32'hbf81014c} /* (0, 7, 13) {real, imag} */,
  {32'hbf8edf14, 32'hbf5e9c98} /* (0, 7, 12) {real, imag} */,
  {32'hbeac7350, 32'hbec86970} /* (0, 7, 11) {real, imag} */,
  {32'hc056af4a, 32'h3fba0006} /* (0, 7, 10) {real, imag} */,
  {32'hc09ffee5, 32'hbf2af71a} /* (0, 7, 9) {real, imag} */,
  {32'h3ec6214c, 32'h3e54624a} /* (0, 7, 8) {real, imag} */,
  {32'h3f7fa84c, 32'h3f7c0938} /* (0, 7, 7) {real, imag} */,
  {32'hbfc28e07, 32'h3f9d9e28} /* (0, 7, 6) {real, imag} */,
  {32'hbf28ecf7, 32'h3ff47c40} /* (0, 7, 5) {real, imag} */,
  {32'h3f5f7740, 32'h3fcd2284} /* (0, 7, 4) {real, imag} */,
  {32'h408223ca, 32'hbf9a0662} /* (0, 7, 3) {real, imag} */,
  {32'h409b2164, 32'hc07367c9} /* (0, 7, 2) {real, imag} */,
  {32'h402a554e, 32'hbfc7732c} /* (0, 7, 1) {real, imag} */,
  {32'h3fdc4516, 32'hbdf52020} /* (0, 7, 0) {real, imag} */,
  {32'h4000fa34, 32'hbfa465bc} /* (0, 6, 15) {real, imag} */,
  {32'h4053fcdc, 32'hbf13530e} /* (0, 6, 14) {real, imag} */,
  {32'h3eaffe90, 32'hc0732c86} /* (0, 6, 13) {real, imag} */,
  {32'hc0087a8e, 32'hc03132f4} /* (0, 6, 12) {real, imag} */,
  {32'h3f941408, 32'hc07b0e17} /* (0, 6, 11) {real, imag} */,
  {32'hbfe5d0cc, 32'hbf255d50} /* (0, 6, 10) {real, imag} */,
  {32'h3f9af3dc, 32'hc010ae94} /* (0, 6, 9) {real, imag} */,
  {32'h4088a8c1, 32'h3da88da0} /* (0, 6, 8) {real, imag} */,
  {32'h406d6be9, 32'h404df157} /* (0, 6, 7) {real, imag} */,
  {32'h40767bd5, 32'h404fc058} /* (0, 6, 6) {real, imag} */,
  {32'h405efdf1, 32'hc03d5027} /* (0, 6, 5) {real, imag} */,
  {32'h3f93ae9b, 32'h3febbbe8} /* (0, 6, 4) {real, imag} */,
  {32'hbfc8edc6, 32'h4087295c} /* (0, 6, 3) {real, imag} */,
  {32'h3f721429, 32'h40df3f77} /* (0, 6, 2) {real, imag} */,
  {32'h3f2753d0, 32'h3efd5ac0} /* (0, 6, 1) {real, imag} */,
  {32'h3fbd8c3c, 32'hc0439446} /* (0, 6, 0) {real, imag} */,
  {32'hc0829223, 32'hbfc2f4d4} /* (0, 5, 15) {real, imag} */,
  {32'hc02b77e2, 32'hc07d28b7} /* (0, 5, 14) {real, imag} */,
  {32'hbe8d7bc4, 32'h3dcbc010} /* (0, 5, 13) {real, imag} */,
  {32'h407f5485, 32'h3f31621f} /* (0, 5, 12) {real, imag} */,
  {32'h404af058, 32'h407b06b3} /* (0, 5, 11) {real, imag} */,
  {32'h40a4700c, 32'h400c4068} /* (0, 5, 10) {real, imag} */,
  {32'h40896b8c, 32'hc0856786} /* (0, 5, 9) {real, imag} */,
  {32'h40afdacd, 32'hc0b3afe7} /* (0, 5, 8) {real, imag} */,
  {32'hbfb195f8, 32'h3fb75209} /* (0, 5, 7) {real, imag} */,
  {32'hbfbbcded, 32'hc055ce06} /* (0, 5, 6) {real, imag} */,
  {32'hc0757cbd, 32'hc05f533d} /* (0, 5, 5) {real, imag} */,
  {32'hc0480b00, 32'hc0cc0f96} /* (0, 5, 4) {real, imag} */,
  {32'h40a2a443, 32'hc08a5065} /* (0, 5, 3) {real, imag} */,
  {32'h40da5c33, 32'hc0439358} /* (0, 5, 2) {real, imag} */,
  {32'h408d1c63, 32'h40253cca} /* (0, 5, 1) {real, imag} */,
  {32'h4082c02b, 32'h4012089a} /* (0, 5, 0) {real, imag} */,
  {32'h3e2814d8, 32'hbe56696e} /* (0, 4, 15) {real, imag} */,
  {32'h40f7a888, 32'h4069c41f} /* (0, 4, 14) {real, imag} */,
  {32'h41046632, 32'h4085b8c8} /* (0, 4, 13) {real, imag} */,
  {32'hbfcc3dba, 32'h3e7cbaa8} /* (0, 4, 12) {real, imag} */,
  {32'hc10e2f1e, 32'h40481fdc} /* (0, 4, 11) {real, imag} */,
  {32'h401984a8, 32'hc076436c} /* (0, 4, 10) {real, imag} */,
  {32'h404da213, 32'hc0715eae} /* (0, 4, 9) {real, imag} */,
  {32'h3fc9e304, 32'hbf9e8504} /* (0, 4, 8) {real, imag} */,
  {32'hc1040d3f, 32'hc09f88b5} /* (0, 4, 7) {real, imag} */,
  {32'hc10f63b6, 32'hc117bb64} /* (0, 4, 6) {real, imag} */,
  {32'h404a9b76, 32'hc0b62dc5} /* (0, 4, 5) {real, imag} */,
  {32'h40282a73, 32'hc1148010} /* (0, 4, 4) {real, imag} */,
  {32'h403eaa2b, 32'h3fd15d4f} /* (0, 4, 3) {real, imag} */,
  {32'h412cc449, 32'h40184ad4} /* (0, 4, 2) {real, imag} */,
  {32'h410f639e, 32'hc0aa2431} /* (0, 4, 1) {real, imag} */,
  {32'hbf852964, 32'hc05e91e2} /* (0, 4, 0) {real, imag} */,
  {32'hc03f2a0e, 32'h40ac4b1f} /* (0, 3, 15) {real, imag} */,
  {32'hbfb616db, 32'h40e137aa} /* (0, 3, 14) {real, imag} */,
  {32'h40395ab0, 32'hc07693ca} /* (0, 3, 13) {real, imag} */,
  {32'h408029a8, 32'hbf7ef4f7} /* (0, 3, 12) {real, imag} */,
  {32'hc1131358, 32'h41375593} /* (0, 3, 11) {real, imag} */,
  {32'hbfcb762e, 32'h3fb1a563} /* (0, 3, 10) {real, imag} */,
  {32'h4149db08, 32'hc1166e48} /* (0, 3, 9) {real, imag} */,
  {32'h406a4f8a, 32'hc028f29a} /* (0, 3, 8) {real, imag} */,
  {32'hc03a146c, 32'h408fa502} /* (0, 3, 7) {real, imag} */,
  {32'h40847dd1, 32'h4066f01e} /* (0, 3, 6) {real, imag} */,
  {32'h410c470b, 32'h4021a26f} /* (0, 3, 5) {real, imag} */,
  {32'h4191be20, 32'h4029b599} /* (0, 3, 4) {real, imag} */,
  {32'h40d3030d, 32'h405d8fa2} /* (0, 3, 3) {real, imag} */,
  {32'h40384162, 32'h412c3c58} /* (0, 3, 2) {real, imag} */,
  {32'h3fa9db5c, 32'h414a2c0e} /* (0, 3, 1) {real, imag} */,
  {32'hc02170ac, 32'h40583e5a} /* (0, 3, 0) {real, imag} */,
  {32'h40caf222, 32'h407ac38a} /* (0, 2, 15) {real, imag} */,
  {32'h3f24454e, 32'hbfcb4933} /* (0, 2, 14) {real, imag} */,
  {32'hbf754160, 32'hc148e68c} /* (0, 2, 13) {real, imag} */,
  {32'hbea25e3c, 32'hc10160f0} /* (0, 2, 12) {real, imag} */,
  {32'h40852f00, 32'hc0723f55} /* (0, 2, 11) {real, imag} */,
  {32'h40f85ce5, 32'hc0b1400a} /* (0, 2, 10) {real, imag} */,
  {32'hc00062d5, 32'hc046397a} /* (0, 2, 9) {real, imag} */,
  {32'hc0679195, 32'hc0a7d6fa} /* (0, 2, 8) {real, imag} */,
  {32'h3fc5ed6e, 32'h3feb82c6} /* (0, 2, 7) {real, imag} */,
  {32'hc1087f7c, 32'h415183c0} /* (0, 2, 6) {real, imag} */,
  {32'hc08d1551, 32'h4081b5a7} /* (0, 2, 5) {real, imag} */,
  {32'hbfa13dbb, 32'hc0cc7a2a} /* (0, 2, 4) {real, imag} */,
  {32'hbfa92ce6, 32'hc113ebdc} /* (0, 2, 3) {real, imag} */,
  {32'h40301323, 32'hc123ff6c} /* (0, 2, 2) {real, imag} */,
  {32'hc04a6654, 32'hc06e976a} /* (0, 2, 1) {real, imag} */,
  {32'hc011bcdd, 32'h4048b1f2} /* (0, 2, 0) {real, imag} */,
  {32'hc1179cce, 32'h41192ea6} /* (0, 1, 15) {real, imag} */,
  {32'hc10525d1, 32'h4007e0cc} /* (0, 1, 14) {real, imag} */,
  {32'h4114de86, 32'hc04f3fae} /* (0, 1, 13) {real, imag} */,
  {32'h4135b108, 32'hc04b8542} /* (0, 1, 12) {real, imag} */,
  {32'h40441b1e, 32'hbf7f82d0} /* (0, 1, 11) {real, imag} */,
  {32'hc0ef881b, 32'hbfd55420} /* (0, 1, 10) {real, imag} */,
  {32'hc119c0cc, 32'hc0503ba2} /* (0, 1, 9) {real, imag} */,
  {32'h3faa63d3, 32'hbf44b196} /* (0, 1, 8) {real, imag} */,
  {32'hc074c589, 32'hc0656154} /* (0, 1, 7) {real, imag} */,
  {32'h406556ec, 32'hbcfae680} /* (0, 1, 6) {real, imag} */,
  {32'h3fa74678, 32'h412f0ba2} /* (0, 1, 5) {real, imag} */,
  {32'hc05324c0, 32'h40976cf7} /* (0, 1, 4) {real, imag} */,
  {32'hc06c9129, 32'hbf21ffb0} /* (0, 1, 3) {real, imag} */,
  {32'hc0604eb8, 32'h400cdd05} /* (0, 1, 2) {real, imag} */,
  {32'hc105f002, 32'h412e8e28} /* (0, 1, 1) {real, imag} */,
  {32'hbfe827fc, 32'h3f9358e6} /* (0, 1, 0) {real, imag} */,
  {32'h3fad0629, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'hc092d18a, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'hc04a7da6, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h40931666, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'h4108b856, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'hc167249e, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'h400b9649, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'hc0dfdf64, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h41326934, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'h4124180e, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'h3f2bcaa8, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'h40c342f4, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'hc0c3fa42, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'hc1ef7a2e, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'h3faba088, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'h4198784f, 32'h00000000} /* (0, 0, 0) {real, imag} */};
