-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vGNLFLmrb94otyc1HO/RvyHSPgzu7D3JcsCXqiyoy085MIwiuJjNmg1n24/AY7aM
MbavSF1M+7ivRcC9s7GOIDbwmV2sd4OgIlFaTimHlKZ21U6yYfZTKMz87CgDBCN6
s8dKMt8b2h+Zgba0L9q/jB9jbdNUG+8g2gI0L49UU0BSUMHws0bh6w==
--pragma protect end_key_block
--pragma protect digest_block
JyDNiqGvzZ6nHx//b5U08e7Zs94=
--pragma protect end_digest_block
--pragma protect data_block
P/KJOxFa5hVdJeWzg91ivcYiHMCd6AJWVBjdav09d6S+L6MTgXS18Jg7hBzyDtO9
Dlw8J5i8vqPzvbSV4QmIDODVNbg4DKI2ygd37Ik7+7TKM1ltzFZ+Q9iXQQdXD681
z9FFyhIuVx0gk9F8pLn+fWogFGBHb8Kpi6hnb4LE6chl2BYMKOB0bNuazbYWX78Y
df1E6IBoNec/QNo+ew8EMTWdqicOAwHUqtNGdDl+6N8x1pCEH+Dwn7KMhtWhzFDj
V6NZJjtPb3Os0rL+7hTLWWQ/zbXLoLROTeObfG3w4yVeCgS52Ly6umhLSX++xWiM
92vh9l8mV2Lwevfhyq7T4cgBE+FkDeVB9K0LDT1GvKYrEx2yHl4VgNhkBdqdxirf
NQgTS6YRPkOGBtbCuuPNzDQoCABmI44MDmA6nbsbrAIIqv4kgfg684zWeqWjAqJy
e17K/BecZLQ9dRIsNhn74GUViaOXeOHT36C60+R1CwweZModQVRbvT9n5/BNwcGE
NFJzFXydLEhNOlFf7dfMU85KChIovdRvBEOoiU82HnO5lFaimeRE4Fh1mJh3aLZM
0spgoxCnPHoN0kTKFoSDIHdu8rDfNHz+e08v1haFlofz2Yiv0DQvse9Gc/tTEwBY
9cCyKrpFqpGnzizgKsWXpI3QKx4fhwxyPSpnHe0I5cy1msdqjYHLoYDJh3rxw1oh
A9nqFwr6tQZfof7LjQYnUH9JQz0K+ToIc33zXQCq9TCSaRuT02Cgq4T+blxHJqQ4
9JbTzfsjlgX0R5GHsQ8hj+P+XxQq30UlYqfcdIcL010YTQ6RoQxxSG1srn2uPnAv
tkzHgbAE93JhfDDZOPdCgjTL9jWkp7qADJzeY+Hu1k5DjFJxGgKmcVYGzo4sd3Jn
ilzx2uCRrsUvefhk0fhrNVhL3OAFlMGAoDDhk+JmtjtrfKQCp/KkM+q2MnmeLmoM
Q/K6Uij6UhAj7Ei5MCkF68f9PklgukwwC/++umTrJjtsGlzhalGiicfsv5CU8mSd
D9kHEmTA5qjv/6XRDrLUOXbi3NA8keCsYrOI6m1MM/Z2lbCAqSghzBssQJNXLr8p
hGUQMoVtzmCSImtewIDsSCokCCrc9OGd5pH1gR1DO9qgOSq2xeYr/B2VHcTqiTp7
qK9sPI8iG0MkaVQaCI3kIlPz0TrY58+WS8fP12AqHlgVovwGMU9IrPNs3BpMmsnp
Eyn6h2h1YNFF564DdcwFW36O9UR4mvRHMRYrHSTr9kfiV5PEa5J+lePJNsoB/94h
86NAzFD5c2MEXPn8FyAVQYxeVd0rT5YY6OaagthQSiNYSyf7ip9IlLtGzm7aWL2k
T8Nmn5IJhBNDbJVdEswxw2y3yTUU7qF6qiAAg2boOPpFch9OFUWAWGeCtCxIgAvM
PvT7ep2iHNK7+QJ6SMkVpYe5D+45SZ+FcRyd2rD3fGwGWETfFbdMgJXcwqD602LT
0ApAoi5zLD5bvHLJ6dAmbiblflTAEZBobPQbS+fA+mDo3d9UnHliBcKPn1oKcycG
sMOo776d7tvh6/3fJ2Ywa+O+5IlKvtmlTrUoNjoFkig55nSzty5mlOA8UwdY4PMj
oue5/KL+ZW5Sl+sI/nWgmBSPtnIHc1HsF7oWpHtSgCTNTonQ+UiiFgEOyPBI19XA
Q7IJ6SsCfDGCWAb+B1auXRShWxGhGjbVhNtjsz8T4JQnIWFJ3+5YgARazwUbfCas
iNrK1m5olXH2RGh5WpbTIXn8aALyxeqJFFAw6gp00wcIr7S1JiCR/jit1wvWCmvl
stLR7wRkFWAxTPwo90TsvKu3zCOurHVDYU6O85Kq3GgPv7YN10C+OLIE138z2xWV
IsYY7JbVX9W7WB31Z4iMmEBinWYdlTsT23O5US7QuFpBczauPW1HOcZZnYQXXjxP
79slQHpJJBcvX07vlnJGzt0YGq8xUQmDBcVNwTP8MvQbLggHYQ8OODZcbC8vwc4x
vKktlwsHYL9sxuGFjmkS9uVnYtP3JeeCztyBkEOWn6Mr5DMRC0hCsKX39m8tE4cr
dpNoiQ7pwtvsUBYNBfXk2LPz3XbgsHIpK5VMOPxkwmyACMNYyHg9HZ8BZ4tmTjyW
a352WMBIuckF1X6da/UQeqtS9GdhAJ9TWbbM8u/xU5nbgC6H/efiK8vArcKA24bq
rMnWddmGM58kUOz4gBdq5u830nRYQ8kjiLBuDGPE2OwcPPH0Hhji5R2cEeyosO2x
ZbKSk40TKSXV2iHPOU+YQWkYvWWOZe5opD4KFlVhvn1m8bv6CCpUB7520zJjvqmE
McGVLp0aMp9iReoHP22MxGwOKnFQyMVhRgkMdRrr4gG1SupWBb/zfQ+MGazLHaEr
E7F/O+9mjIjn3MleOogq8WW++88WAL8Gn/Vv2aM2sX01bJurN7/atEA0M3+qMK2b
sZvcglAY1783ZAx7LLJ1dY5wxUz4GsP3s1AtZ/jx8fgPgebT+WNOXn7ycs3/jo0e
6oGFH/l8+FIdUQeVNtXrd4IMtXl0RgfjJawaGda5wQuS+pqTdXyPZFecwsyxg5fI
Qys2o7uEC17Y00MuQ13ZrytY28lIyhyF3GQm4x1wwEgwtZOwNc/NaGhWK6OtcHoH
JTfybcmsvR383FbW80vzQndUGDC29jv+bwidikNnTKsEh4IkC8xHTOfVZ31Vy6kE
MaRnNZq5BoQ5ATgG6zYovkCzQTY0B/d6vi9jYsDZb8Hq9EtxrbIf6oxtlRstsZ/t
7g8eMFEsIb0zO/if9ymBE98Hi+MpZOIXePw0THqEO/xJ8Q+mrRCBD/kUgLPNpgtp
RFSw2l6Nkd4M+UXXZ5QKL7ceLopDRP9V7T8F+ifZ+cMHSMSIh9PpXXPKr4zea8Z/
HDwdKlrHwGYlOxturXD1nAWrhO8QWKZ+2MCH1Y/pmD23gIkkp7C6kxs3yTT1uclY
/8CbRGgZxl2X3NOVhX68gwJstwt3Nr6t6PZBpWamyGDn4kNrZpoZWUPR/Igw6ToE
sQuxI/cHlboNBqbppjSa7MPjj5mdNBPAI1jK2FJ2W0y0WkzGvvGIl4TR29qsjrW3
yvFNcIU2iWlph83NhzMVFaDRERl6QjLSD0MugqXrAxbgqMXnLpY9O0l1+X1FPCEd
hANFIM8O863zV7AypSgKvWaxb9vhbjLWXv2SjNbmJcQWTb4J7tdC1GMt4oTifRQm
+7PFwg22M0cyt+ZopTu/7HdAS0nG/2+OcFtq2HyPlWQ2oVt+jon5ZTLEdADJ2mKx
SBvPvPxJ09tcu+nH63Emuql6ntzal1v43YUvdU614Py62rgGsxyw+MLzIWqA1T6y
Lv41vKbo7naG7jzE0WsWYJwHHKfI6OSCOXc5CZ58RDbb0jNhpNRL0ILP/oEmt5o8
6zZIRKWh3h5SudcV+1z8T82jQFPcq9kx6xW911IXniKrOh5j+dkFataa5Y4Lzcqg
c/9km5y0ZvkQDV4JDuPSE6vnWNhTYHNj/pQ3+Q4Eb2nI69JkAy1YOPsGfcG+s43N
NICRbTifGBxdFiHz+7s1Wwo1UF2eWiey6uy8JLjM3auxBNXtxfSG5GQT43n68H+z
DPhnFGzCh5EE01jpg7lZnQ5Qa+7yrEfndWwT2WN+dyrIRGZM4gdjbXaTJwW1OjeB
gYyoHzOs5joPoUYVlhES53w+SbFcfhkXtxUCjYjnEIiP3M0f/HbEaGqFOr5nAYFB
Un+hCJ6nnPVcFpzrGjrO//NU8zTO6/CPONia7cGiVPs2bEimP1CjRb0Xji5IiTrr
grhzkBeDVBjauUgbiRBTrvoCWz+IozRfFRVu6u6lRwyYnktAXSdUISbCk+X71ewT
FmJtVaZvgEaYj2DgqygTkRWq0AesqxBSG76VoT4VFUNxrJ8AWJSA/6psMr9sj7S7
ioiuZ8bi0xy7icnZxcxdsqUEjENVjlAfOyZWZs/KsCDINoHkDZWFmC4PAy9XhrdM
jWHsVougjr3sLNcO0WtMv+/j2/MAaDruvqaRluLSp1wiuGccHF7YJ+D3bTDCd7Ka
JuuS1C86VkFAA34+AVYKZKtT0sAAqUCB08DU7T0cHnBlMV+UgwWf9BfPLAM+bZI4
iDtfGgtR6Ij553QWg+RKC9YInfc4E9c0a4a0sz57vfi5Zofvd9Z9eMiuoXxMoFOh
CgZJYQKpFvwco0APolSKKquhTm9Co32zvDVwZQ7PqEhFnBPa+EmIrAtvUgd5SdzO
0bre9oqeZ6HD1QauR6Hoaeo8JWhoMA6iYKkrYGChpY4J4dVBkrTee4AS5vIgrVOF
ZckcOEAOfGdODj2oedwdgQL1NromNfp79SNPj/EG9gk9+EivvPw0V6YQ9SXgc2ix
VzB0aWOfydsScvf0PleVY77nTOL0ar31vPJArwTcqPhxbsPHmCdCAS8eAod6Z2A5
YeMbjRdw06wYcFYvEt+/0gyE3LWT3EIyOzYdvLQn3qyef8cpvDW3z3xdNT7+Zzsd
VVjkhU3vnjhfiauI2RfVK+g4J03fD0RIJQCKUwDGHfEUhNucGoFd2ooldHuYGOy5
Rm73+JamHceGpNor4ht1xhOGzmMNCuFawT/Udc9zLndJ3hPYRnawjkRh0oObMBI6
K1Ub2vFdy6NFriOMwzK8hJ6qG/dDfsMjSvIXcoTIPbtTTqVFzjUzVQWeRl9lryRY
FuHZs87XCbg13ePtmbSKQ2TGzbBbb1E/p0VhIPNDLM2cWVvIbHNMyLjufZVcZSKa
uFvXHakXGSdO2JbqLijOXTyMZuw4NppaE4rkLcLVVpXY98lAOVJpR0IipPd3wbY7
hBkURrzFLeabFWX5ZTN+As1LOescVScMshkMZmsAPq2FHP4aC/Mhc/L0DC8Csc/C
q8wXSzBuu0z+N5AGBgNDPvhGAWlEUJjPDwwAa/KWqyp9nUPLdYzM8xCqNGdi4BhQ
9I4DRXk6wv7IO0cXivSPiqrGDBJzluDjzxJV51GtgoOfHVT2Yr/vbY/F2970C1PZ
dCkCc244N7KPOzVFFpGe9MTfQ/rJfghGxLFiX8E3v/+3ogcREEuHRoypJ7HZe4Y+
qvp8m/GuL4ywzJnEl0wJso/gtblocxQrSnDufZEpepfTBOKQWud4UvoyYRx4TseU
+jGeS8huCDsO896LYHo17dEwKThmahpjyhpdejmbtQMPZom74NEfcoA0HxNlMRUj
q2YKKsrJ3JVkxHK4qYJ3uBFzcLBK+ihMugQAKa+VDia7sUfON7k2sCoBHhzhEJ5v
/0Rpu9CBBJVKepfBGJAsUxdX775u4UpFzqQ8ft2HngI8E/RKrYgbuIubkN0N+ENy
dKnhNnJwayyF9zlW0JQj0Z2vJWaNp7GIaEOIRbWTThnMaxT2fU7CnhNS5I14Z/81
HeojfUJU2FJBtoALuaJiMoOp0g5vTvnUpqmuK+tQQ4J1iV5PNjL3/XOc/V8iXNzH
VuSFN/sZEdwa7cX2kcWg0vzuf3szt7BCcRamOSUrLglKqABsEtl1jTnvbHqRFdEK
Z2IfUfdQWvYPOTDZAvDQnY6KFYb020Q58YW2Qv0xTaib2xaQQaC++4I3qCn9zVQU
/c4sqtaSV8kWTu1E5GTUWOff2oKb4nKSyAx8XQQHIZAebJQC0N/394eJViMSwRHW
TXm97iT/u5ZIJysP+7LscntC3XMbyhj61iXNhm5nMAc+2T8tFqK734sHpx1pR2+2
vrurqwKL6e9DkifAZ76poWVBo+U51Yz92KpHzT+VDJnB+82rhvbp/ix+DQlil10s
+M1Blu3QmOncMfY7IMKAJwZvcJuMWbPL1xND5E+5nor/ayqNBHTNj9YiqLBDf1bL
0+AcEoCrZ+NavGhVoRNRNVPlxnGbjKpogyb+qcqTsPBg7nTn9AuYxqxwowyMst8x
uy++aShFkO6xT8m7Lf5qznz0xIOuF1whe6L4ldRoH1EPMYRQzDo+R2gh6eABWssq
YQNOLX31HCm8hcY2spYFLRofJBnW9uadaH4Of1AM5WlDojf2Ak8OJKmGKx3eQV+J
La1ZQlXFymA5J9dZkVzHc1JzeWcpvtGjCqFQ/ZuTtyaIZYCTg9Aq1uFF5XJEzhQp
WvP+fcckIPZCypkIuinSZBLSmu0SBQM4Ai192uei8ZRTihvoRIGZKj/Gh9DRGn/i
bRT2LtaUzOPxg5kL3rdQyfscgItTkac1QfxA7jMbzfsXvkRY6EUpi2YespbBlofU
V6tcOhv9LVc1tWDuTEvYYMTgg4JUKSw8hRCCRcGbkU4dGqVDt146H3DbRv7169mS
RWdq57//1zSVSeLKnLtBwWVvhMtwtoMWS0gDnED1Zt5o19n8Gaw6TCKlJypjsvsb
0j2lFzbB1EYvCvu0hTQoz+w7Fg1ANjh7yAGX1Ik+OaF57dphjAp9DreKPuDtvH+w
7mygsQkUqFUZUa75XWBMudORYaBacRieKbH5sBxxwDPzeOxxYkMxzA4SoiB4WLXx
bB6HKkbqy6WUhz0fDZvXPIW9XFpdXHs9HsKszGK6trBSPx4Txh5ZIlkzLazXRV61
XeKCgEbCLjfQ3zJTPb8SI2OCRZpQWbCNOMgqUwSJ/us5NuwgBbGQKM+DbNdZ1mlS
WG7uNvB3dpGiyYd7k3BlGxquvqRDinTq5kJZgxghmaJklEz0E0zdxz9s0nT4v9zG
2RK5afqFToi0y5qTrzPU4vzH+IISwdHKnMTFA+HA14ykkaZ8C2aaSsPyUBmO3NRf
0pVbPjZB4PRyDSs+q8/SoXKZttxiYJA5PReoepoXs2thqdSHKyXkvxUJJW28lA19
u18RFbvtii8ko6f69GWJONQ8Lfa2qnK2uXBXKHbH5RVQZKGQE4Tms39UJJoLcaRi
KdGvlfJ7MlO83tbo7WsNgf9PhAJI/BThjLUzlXbafwC8eRxLh8aeJz0NaEvtDfhK
XhxDsk7e7Q9WTmnykTMtyN4BH+z8INRRBsNO1BKL3E8W7gFJGR2CuQn9/q92W5x8
MjueeMGcNAFtvL/S5WHw0PSXt+su7pXX+M+dugamaJZyQL8hlMw+B8RmDIRKksU7
cM+GNlvb9I/+0fRnvnnyjBN/6oCdIZPYuW1prndcUUsf7B1ADMZ+AMmM/+prDEae
nqQIosXevM9yf5u/h5GZchlDrV5wzHFd4On83zrtr/YO6w+pVLmUoJn8DzTlJfMT
ailQhQ9AN0dpUouTau/uze1FmSz87Vcs/cfFs8RAv0t19zfrKmjaZnuxQzaITvnx
yFntP19h+Uw/nHAycaueM6g57800DwEj17nED/k2xEwNN1iCdJYvnlMBJpILnaUz
CPDlQLOXaYnKQacrVswMNe0Y7biWwXsEGhK9cFozrUD6H+tEd43EhkQ5CEgJFzGI
bwz7CkqcnHMEdVXad/BIXS6d3DOe03MlpWzBjx5hYh8geP3GppFvcpq6pSgJ8sCl
Y3mjpuU43FKGL5JBxNSIpg0juL2bh6xs1MgnMM4WaEoKTyk1nl6HlbZr3d8gMFJb
iDQ2hnbnH49AT7T0Qblk/klqMHm+71h98fidfrM9tMhQ3Yrkdqx7XRrUBHuZSZDJ
H3VPrCarDFJ84SzQMlkiX+GZ/6F95hK2X/r5CNoyBvlHR9Q+FqBloB+Nef/teFKt
zvAJiEJwoc5QHu9JhNglf1wftTYz7haqc4BcXiqf+3BMsfZKT833bg/DDD+gdFgH
tKO5M99mNcSPF5TxA5bu+OaL3n1MZHK6zBBYaUAHc5RQknf7zrhX7N33UmNVU9UN
rJtYeivvWLmEec2yydewldK64g2Aihl3Cd2OVGyW045PpTlQgtZGqYdhXvdAMpwD
meY+83/xhM/EqLUEwhAVpeBki00rztEwDIvBMTLBv1LK9v/yF00iD8i58PN4BNgc
v7w70qsrkYrdcFb40EeahgCJDe4uTdHNj2DcyrnrHD08hPJt0VDXC1fDfAeKg0UB
8ABdXvaaxQAP9SxAIqRiPNKpxXN6KK/2Mg9yWn3hRzLe7nHe+4lbRpDIJuTaKam+
lEWQhIX82Pr1uuVQQ70GIufUqIl5jJshH9FWpkf847kZBI+Zz1PhLnouHGqmA2xi
c5kcCxkpK7IhxCaATOtpEdy/06JvXrZUAyWGZS/3qBg1+zK9yhtdyZikrW7FWPvs
pyWNdwo5+roTWxF3KGHjVwUjfhANp3/Q21CUrrIEuzVEuxCvpWuhqgPdepeQ6cxv
aDsj+4+TXfwKA5MPYULyDeRg0didZuk/TnIojMwLEnyc60t6yS2x53OeII1TLx+3
Et2oQ5rqYBxkuSQ0T/2jxGst2zbZYCsyixnWTO1s+6ZYQ16TuXnHP/wa9H3mm3GH
PjjjVADpfTTviU4ueLV14CoT5y2mVXSUHlKIe9sWLG+l1O2b2tR14djEv3MJC1U1
fZmfX6SbMj1WSvWwXWaBafgCvzNB690Cv/qd5NeyXOU0meOIHH+I9HI6rWmGIeqw
dlnRBgLAU/375d5Vw6Y3lB9UduJr54DJnLzPfZ6F6UfZD4vf7RYVZRfAfRHAUCk4
CXpTosPnMosU0ZmOktJFNiSv5bBjSaB7z7L+NRD3ipRh1S9sDpk3qoKJXCR9lC45
f2mvUJ1Fj/E9IXde4Cwa7+vJvetgM8ndaoxxRELiX6mam12i5VEzjBXQG3NpFx7d
ypAbp1WyI18PFzdzAuhRabDEYcT3s6iT9pSWi5d8sieEr2ARIzjXSsAG4QtQI14G
moCtXMQE0buCIh8yBUmGCodlwRzFN42hQ8RkprPUz6wZf8NhZnJamY39bvSyM1RX
NcbCdgkfM8reCnMxiJd+pC4Kblo5ybyER3Y730ZC9xwaMD8AaDHkNYCX5zkQw30v
z2nvj65naM4pB9jRxcBB1F/NgS09xDlMEZeMFhpiLBArQr7hY01pKGfx8cPgk7/J
izfFdLOAYrJdhE1k8lSzcQi6jPSCijxXZLUjGTJ1jnY0EyCflN4YymLVRRp31Vbm
7T1sMAkD5OmqnrCUyJHZXD2CaoyefuuOaho8vCcjOleSSQ27lwayNtZC6ipTo1PC
qh0YVkxXNGsW95HfE4mwW0m7E1Dz6NoSP8NwtmziLqiogtavR6YtxIeZu/6IysIM
H1PpEp14xPn1ZNVk0GjSPmmyPyRZxlCRMMwI4ccmriTJB0SL1Wd/EXn1q/B73D6u
gIA/C/CVUGL7KWu9Mto7xi6vJMU9TrXosQPsfX+aSEO3Yf1I0lLRPTf4a57daefR
dy0fqLSJS3yt3FEVNaOlvnu5pVXSYs7ujDFOF89n1u9RYZ+CCj4fpX4qPnfPyDB9
EiR22W96NfEntzK8UANg9GRw5GiI4zP1m1Os7quVuGFb67lEF16/an2BYCgIi3dp
BkS2CnK22ZLdTA5iDzJpAg6CmoWWKyydzUsEJCFPjc8pXS8nlDqcIC5HshDyzcgn
QRvqfi4xuRSDgaNfzMlliVGHeO/vmrdl88qg7ny9u35Oin93X0vs5GXQ3Wwr8ip0
aDPPzb4TS7LRoTi2vjsi2qWIZm3owlcM3IopwAsZKqRbkOdU/It+oHR8BmNBstPa
krIkYlH7xv5e0WGXCC/ndeGH2yqtWxDpM6EInzUepEdDUgwwPU04aX0ur7wT3zik
vH5OMGCulP+O9VV5aqHM+wKzwe1b7SjerHbi007bktNzLRVeVL7QXCvAOsI8EHQt
Mycs1MJnsnLDJprZyArl2YN7pGtVil+0fRbdARLayeiUb2fgGS3fE+2/NjGCYwGh
lb7DJLsYKsW6kfxP8aPN0ofKLARDJ65IXzGwP6C29dHqWwbyq++ZJ53PIRws+hv+
kNMbprNHPTHYotwnYTdce9uAty2w1513/dvJ1Np6xsJ5l78US2GUxi5ynCyuKz5S
E6230UtntZWLOK7mJD/19lpMekNxLpsYVfb1jN1oPu+79LuwE5RJtt2GCbqU9yxA
3FyWVyx/elHV6w1od+xf7K2Y+qeqyYy2MlK9KgGQiAk3eKsEmR/ymXw4pU5qsxDY
pDo2eEl+GcPP0OZDc95uS5zWFk+b4gPdfh69jA+vd09RCuQmI6EkrE20fclPRFYf
iYE2PgSJOuC4uUMhtpQZ+0oWYRTeG1RfKO2AXJP+SJS3AEaqTrjGzFo397tkwTW4
z4eEpi5gy1cE+Dud4Nz8vWnkxzOr5g3TRZw5UqT4fCxXHWKuvHCq1UQijudPGQSn
NMEZ1wxdGowSW+nbmP6gt4DR0ZJ0d7XD3gIgPtZGE0BTw9FICmOQkJgZgKHaKblk
Qeh4rTSi+S34fj/AoAYYQlaT2rY1bhCYjnxn1HOdSkEb8lu4Jem6LMP9W3v+wX98
bWG06h227p8+sQhisb/fuTWD5RZFxWVX1KQCJTnbFXvD/JgH9Kli5fwWraKkCPYL
9nI2KJLixACpXnAV5gNVdBfrlA8dYvkvaTkgVYm2nOUn++6iXVMsS59LPOvhVcmG

--pragma protect end_data_block
--pragma protect digest_block
iV/PgH8db6AcG+Jk1yvqzbU0Rvc=
--pragma protect end_digest_block
--pragma protect end_protected
