-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
3bXzxxqHnPQQxf7dfo3P15R+63UnMBL1EjaCgBO7DIGoJzIf/kmvQNd89M/pvbPX
0A82sUZw7AtyoDDeOUKYS+GlnZpYriCRpJEvREnQxBIrpQ2l7/MlceajnBtPJUAP
dYhpM3WPrmt5RIzPkk1D1e+S24JWYTfLLIL8s4f9dec=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 23312)
`protect data_block
uODwHsxafe2cuiHMgo6QwT/0ma1XWc61LOQhqc2vTn5fDuPLiF99IDfYa76YDsm+
u2jAlVB6B32QtNJJwu1/ZZU9uqWCYr4k2zYApzaH+MDGDQQU43ZlngRWIDR09e9L
ea8WuULhJoTX3HZ5Die3Q8pTMv3MA8RdmheaVm/kenlHNT1K4RjeokXPUfr++1E2
fz1t8o9GoTywMOVKNWfuhwf6wkZoNkYGqjQV/us9Ka4b8RhOr7vTfhZV2Ulc4iUX
W4mwM4XMflosVxFmvFc8Ci7yBgblUiLzV8RTmmMacPQm0uN78ODJbmB0Dj08mww1
pXN4fvviJnY3KWUcGCeXyiERrwV11Y/TzeoayMhW/4f+mwNhRKoC59mkml87BwAi
m+sJCn8Zbbfx0Hv/ITSBnF0TivjdZFLhO0UmPqkiKsR5b3CYYMWDZQBa6FJ+fL9B
Kv7ZwhH9gcGzFxuF6xdMb4Wo0kvl9ApkdY/zFGb91QEMn5qh9dflgvd0oN19axho
vkJrtg6pXbH38Gx1Uj7N5tCH3UKEz3KaRXuc7Tr1lFsGILMU6V4Rj8u3nywEuhmc
Lqa1yPjXy4AJoGTNS191152fhRuP69htJMo/xiGg26QgQeptsSUUfuvjPA+Vq1fm
fHruxgYVov96P/fnnZdmuZJjR35EBEU8wHFno72Zrn/+5V8INgAM2KD87GuSL2QU
ZXNecdb9XiaU5SiJndwTEF3MYNDovXHoyxMVClmtbqaawZXa1dwfGCOSiymQY/E+
Oc41JFv6KpqZSP3PXYqRBiZz+7WQhytryvUkfPQnZHA018CITWMYwhjfP9XJUcLP
akfz0YtsZU1kmVpaUUG+7juVNtJBtikEgOk8kZf9MVei8Q9pXOS2JGL8DIfqJB6B
dkE605/HUtUUuOmQWjFjSzlUfvDzoB+V8rxNPio4439iVeYKmJxoexU91hr2U2Ax
zDV2+nCtBTl4Bty4yAdUY+X44VtoMKgP7WINDn+LdfJr/YfCOfguLI7DkGNLOSI9
UccCtJxywenh4alnN7U9Toh/YwdTAyGXBb6QRvBN1ADwQB4BXH+8GvE6TBAU1eib
lDwIPLeBzq0JpBNTK2on/DNQZRwVxz+tf5gfJms7ixeTQuWTCPKgz+SkGS4Hv/tk
ZyfLXoKwihf2pumWHBiEpvYitRLzRJJifhiS/X+EMFs+JypOFUVj0irRxDmPlQJ8
tzZWcbk2s8q3LdMgq5UN/I8Ln1FOUglcq6N0CHBqCYQv39KK/wDha+M4DSkRViQE
WAjI/jtDQOhLRkJf0RHcPkmhZvCztOCnOwY14J5PKXckONwgSgGKpHuQ8YqiVMLB
FnfEGr4XN+tBZkMH+IqVrBfB40rbGdL54DR+oVjCv+4ujFltBdHqzRhlJonkgJO+
CiivGnyu1JnlIBPxLq4Me7ixE6Bki/HXCny4HMwzS7eTaylxJFXD7//ToFPnqFUV
xFttjNjTxgjP59zE0MWbJa8KyHX1rX/MA5og8wkYzcdkyauQYf3x9ntCCIAwLzwn
tgjn3LY7lXWlrPie+7TsufCAdgdBrIo619F5f/ZiCpnG9UMq3IW8KO0MtnED3SpT
95ytJb1j3tfkkan3KCYTu07sByI4M5KUWZAYT9Rl7SQJcirgvnvAf9/Oac71SiCt
40eoAWxeD/3VWQRJbocROTPk/siWmY7MmM3HyiKXX9wLakHVA48yDsxBk12F3607
NlXC8T/kTRnWo/8g8iI+P6cE8FiA0d0WJrfrp86/PO/6nbtUF/Z/NFd732lyHgBq
8CkvjhIwAtY+XVvkW6zk2VU8oREXg7RuBpADmXYeqEvWzORddDgubftjWr4e3vMi
1QFUCB2ccHyXPN3KR/vPew8hXZf5LMkUIts2YRbN9ovtEoCrzPeZn4mh0g8Lm+Ns
fk74TFnBZnNqtgAq3nIfbk0Xq5fRV31mAeMLYvzv+8Bfpp9UitCh2O5iGmz1xSTI
6lHy3EnFkH0CbiCMeXKVt10X/MUGjlfPOcv6ufOwC9JzFIY4MihgMs61fGhm0AMa
+uubYSfdAVnb/TkMCBUxqId4kSae2rtt6UUaO1F4LEt5bHZ/9JfgDP0CIyu6VFyc
WesNJ4bKtELra7cKyI0X1doCQgr2iF7yfxFJvA4bC55J2z49W2CxQ1hIOt+W2qmh
QREmbAaaLyXQINr2aZ7fz7FmtbjTNVkV7xOM27OVy6KvrfYLWswhXGsVPhp+lw2H
uVrUtbusendkTpQhNKkWKSOhfvsvVMqF02ClR7u8kFtvHLpYpQsubIr8++BYQBC5
W44oiyfNfUmdI6Yha1j/jsQ5WEIRUkVX484g26ZR+lTOCOVJew/661dI8iA0lPZA
8xVDzIyDMTmCPrWmc+aPDCgDbxNGm7hm/iVkbjvtBCp5fvTbB4toM1tdcih7XJSD
iqJQWp0j6slbo4Y4c00a4v2g78GM63t9mPMdfD40agZnn9IccqFmegNT0Z2dt1kb
lscdOoijM02TjeDueDx2YDbiJ38kERf1rB5mYriAsf95snFr5SFLGhLqq2+cA1cv
JLerDshvDVvIlFmfiFrLgNfPecEyzAYNe4QrJK0s5yfsBg7+pq7O8XL8qXkSt6k2
ZeHfoIaMpa49BDY4I0j4vZs9oCUjbQQU3lE1GPZP2WcEgXSs1JMHLiGNfkDfrWoZ
thd/tD5wP9yo3ee4fxVpxqS9cy36yvmxvCrbd00RKp6Wa53GlkvMjzkUQ51pp0mB
ekIKQUTi0VuGJXVaMw8XwdSwTT2lpqjlB3zHaOWpXsS3Y8+bZe1QsazZz0Lymn6C
ggwUjAo/U6+r9QpaOpQjCxGEFbR9iUV8QzXUOBxwsPaPgKJ6WED4dxB1rAASVcR/
9gLryC7olY+lV2bWdSZfBfysB281jihNx2pXAvVNgl/L2cbQvYW6JHpIoOLf5jSh
etLK2uM85dKBKAXmQgfiSYhH8bNIDujFafvQ6WpekXPy+GwQZAIhMdJGF8eItbC/
jot5+spSTcqGA+6fXLjyVRQb7nvbiURnwEaEKIv8/jbvvJPrXzPY7pfkZF5ng97w
5dfu8RPs6b9zoY6Y//tK13ANJAUhDIe99Bji+pBPD1k7VFDgJzUSaypdkW1ZXaze
NKmfQLirz9Be4d1O4wGfzNHppTtcx+9v43xPb1XcAo48FBWaxwlwfCd9cKqeonTX
oBk2w59+eLSi0nT5EWM3bLLkDj/U17uDDnLqY4lL79x7OnM6cLQmuyxscd9pz1NY
wiQGtxxoq7YghO8a/IwbwGWtIKwcC6Bsv+mejd1Jaiwms9VvDzmKnSrA9+ssFrHb
BFdpimzX0n4bD2Tejw/8YyxvZ7S+Nab/YlSQsPCxrypSJxPEvfxJNKrImkl9cQD+
GSdB8zNlncF+vyFGTAkYYw7pyMzus48YOvk5VtleTcK8TBhPbQapPw/mcE/rqP1o
Tpr5CPD1n9GLLsZwOfWvFWQJsepbtQjedN9tJMXHLGCYmfHdyawTehh5QLi3pG2O
ijUgjtwrif9dBvs/HBNtDPwrw5wmZ1phFgrhAV91oiRqdiK647HadfODY41nr3p0
Hw7Nw5+bNUN7d07KYS5iPgPtQo5tp3YTBoBjmRy3hd8vLmz22C8fTBYbamfWerWv
RS+iE8Tjai5LFXE8ZCbky6hXe9fBc3CoK1Plp3x866dWoj4g3SORTngksRtXhxNC
7/NBVwJfrveuwqv8ej1w6SxCCEWjMierjjN6uZNXdJ3dwt1ACxvxkuHyXkcoqQTT
D9+zf2joVbSmxznTsuJkkjLbv/PUsDOcoejRCeI97pTgvjrdDmVzib501mU0+HFS
byU1Fr5/Tm/b8qM25cjkGuckBKRAfYz0dwpwsHetThA+NkUa1Lf/IwUdhCua8tt6
ULmKksUW53Bxc6V2sgrZRJUkkf3IhM14W2usi++LzWN+/jXT6C9L0afDSX/JQsV6
tDHeaW1lA1ePe8FU867D0RReZpEiVLBr7wbMXGovNnVt8ztA54T/RD1/GhXT4UCv
PMr1iBHR+qKR5vH7jDphuktEBhrs0XqwHLf3zXPQrPtatIdTkflbpCAbu1XEoq2Q
669TQ13ZitXuRJPvITlBkCumles4KFwR2qi1k4qMw1A9hw8A6f8AF5bYRzZQnMpo
T1LA0YImN3fpPQ/vEpWaYWJ36VqiIDiRzMIj72rJh1PxBxHn7/1p/GEDHVBNpk3+
9tnOjjw/ajpjhT9aROs74LSRrMGJYajLl/CLm/giutnTzZW8wln/ueE2wP24B0nM
ghmi7yNkl3pHcbkx1EdMgLfN9TkVH+XT+eV+ZB1/3DOuhs5ZHhL+j0sU9zw5k3Rw
3OGFQ+w95NGAqDs4E51WnthPGmHkO9dxvvR0MKekNOE8yF7prqGliiDoC9PeXE/n
lVeOXAIqud47B3InccpRS3vXKuF5nAKdd4OfB9q+6hj/BFFEbnjac9zlAdUif6Sx
6+/IVex9dsEa/JRmdTrt5hDuj5deGI05qxIz0sXVvZokj7RJLk5d9vHPOTZTJcbV
PwibeW0ELCBvGv1I3HCveKup0XtrCrnIxzLzHHX1lpwnHOxlFTBWiFgVzvV+veqm
QdTiH9ooV56ZS3tnSf7iJ0IQMj77Yj/TPEaIkF/OX/P1xM+4ZREf/jsrh/zBg14d
rf4wUdIQuCOsObrNeMRaD+IRQhKwxW61P2kc1yGRIoy7jziMvQUBhywoOHbRgI5I
4mYyXzgMbaQ97QNL1zNPWzv1bi73ny4kbm9bl9USsKli3/BwmrY5LQijjNZjyK32
D1yzBlguviFWDp287+3uf4EECjvRyNxnQrMfAY5qGPYzf+l8yplrJMk017h92J4F
ojBzE6+nN5FszUkyjXmbpqRkgjCO0bKCpDcVUyVECatGm6kuOdfjBnzQe6DZhRoc
U6bQn5587iMEBLJ8MAeiB93J+Cpw5I2tGbCky7JjV5qewEkWLgzVD3VSCipIk74s
re8Mj1HlSI/3HWx52tylf+mXaFx8EQbQ+8xbXkmar4kezbS6JDGjFu0XUGOhTNqg
7VHV1ylN/ynLVkjjz3CYJAZuHQR2qvRLaZ3kU9UWB//ZxI14DhUiwPzrIDepZqEr
JtGhQjknr1BqcmMUegJnNCUKUKJFjpWGRam+MWNqqQlXN+JRA1Aki9ea2OieQLZ6
UbP44w5aD54XCs9dZuAISd6dpGP5/AaLWLNgEh47Gh5sYyGdeS5yrQppGzk0Rxlo
fezj7yqP4Ril0papDiUuD/5zZSm+AoEqg1XVxFsgonQ3Ls8qG9a8R/TORy2GmGIF
1lJXzpo9aVAfkenbEglLTfem851Jq2F2VwZ2Vmyu+rZ+AXTDQT4AcajLjHFuGxM/
v7v3VnqZnuFv5GLHJMDr3FbuvlWc0lPyD/zMZtBwTXn8YYzXjn/5E0aD2Pkch11i
MdVqGZ8pdHUe2E29MaRNtbS8NIgAJZdVARUb70PaY/TM5ndLdeoVfl2Jt52vBYyk
L7OvPl3OQnUsqlrkO8hBg7gB+dXy/EmVDsP1R2cQoFtJq2htjGuu0KUJFq+Itose
j4vYoiBQMWNXtjEINu8xwBscp/d5GehtBxrdutb9bWUzRAi/2lKqzcolSp+fm7qJ
kBoZOkFrciFFIf5C/CZopBucqS92VhbvHTzT2A2iCgnxV/sGYGfpsBwf64Q+QkS9
9W6sW/5HEhdEAqbsSR0SEKO/mbo/MNMvkr6xgoF0Vdv7v2bhIDp+EbyKhPHyMP0H
t3rc1Rb+g6+dQ8spYc1CJ/cdoARWTUF+LnyHrtq8KS8BHAvn1hoGQftOBaaYvJhb
p23o16GF4QZ3JPERfGXQG4y2m0IEkP/8mjju9/A78SHYVeEi1njFN7Ia4UfLyE+T
qINUi1kCNUdbYBK2T5q8iFms2Oe8Nn3l3mNp2UqlLiLoBzzHRE48vqiOdZ6RcxRe
BhIuRAniDKSSiWbmouOjdCMKldWKSVJtD4/7f3YSCftMGouXswl/90BGDFaEymir
v4Jzc9J0TIO31IId82oWn7koBxLNdG9acjRTtC/yscY7OWnCdZmH+opMCOQjHstR
khyivS/tN2alC+M0aLJY+KqpnTnASIS1LGTJpMKKT6hhOaHRYlc7yge5Q16T5jxv
C3Q6NjOOxNC+tx/Stf4DWOCeGzXF3ukMjB1r5sLbbsRitowU5p6OdwFmB5CacvFt
6Vba3hXTKa0lx/MFvDJyF9iojswe2Su0EZkR4hjYYAYL0Bb7WjTi4oFIggtGd6pt
340KLiTmiPcV7PmZEzVzeEIsXdjCmBUDYiXlAhTS4J3Wahiu+dmep56zVaR06dzA
p3RFwtX5THGtJAyn4sOrTaSSD29qaMCjFbVBcDLCggwrsOfF4Dj9vlGDPiRCFtQm
YxuFJZBNkJVeKMJQafqAuKvq45rKvQfCZZnPsSpba/YYQmMknqHeLkdj53UNMa8E
1bF7wgWLaki9R01iXbMH/53r33vfli9QInRWQUY1gAZzzS9ThrKTFQzFpJWhwX18
9lJ01JZsFLL6pvr+Mu3PoGWMwbXCrCO6fiPKKm9bCvOZ9VgHNhbFperewoCsuY9I
bYqWpn46JNI+ZX3DhHKWx65VTZmedUwEYbVttQVSXbox0LunOtMf5/G9mQ9CDpNi
AboEWGd2nPqkWpxfwFVggd6Z/30migkrRCVlljx6wBWy6p79Brihs4jL1bJpxktg
E3zx6Y4aV1PsKEr8pT/m9iFXTXwUQguiA6YlF9LD0JIH+iArsBY1gNn0o3VF/cSH
MyQtjPcuX3OmTdB+aBK2YV5TAvd6KCCqjxd9uRgOKruIKw3sM9eQYyt2rBW7IqRx
1gMftPvoPZkVGwxW+JWs9OfBFCAyxy2und7hcPbLVBwmxaYXP6aY3fQn4d3HVfxi
zoM2NpEwvxXeyKXqZ+TxYLZ4+qTa/OzO8YLd0HZb7o9nfj7uPflpGrbh4xCdNfar
3tGkFlSUACKVcqoOZ4KR1nE5p/uwv6ooHGhnPwrCTWEJvUnq8IW2UEi4nCQ0MN36
BSpcaw5ebwnyV9Uc+HmquYZr7xuxBxZwXhVNrnxUwFwWCDLSGwk8qYaQH9kdWrJ6
EDLJNp3Jui8AhH5SQofylK1HtyLcq3nXLt87VYHSN23k1CbfmAwNMEzgBnWil8ZJ
zXA2F1kGctJ5aVLQPyATMlhK3iD/4rZ+PDEWoE2oTEtEHyxTKa5BicTkvqsnklWH
No8VKHLc3MimcTAYciXmuOe48yX4LFDL3qVp/hfrSc/Xihf618uwB6qqNtrNBeoo
mIXgAWtBXgB4ykxR1V4McMM3JwHopxZHr1EyO/68NjXI9UIAHEeMe6WHTfewWdvj
c3K0DnRRdH4Es8bF+fQLSkpkTfBKBSnpqUnHmzcxU1hExSe0CNRIP4zKg8GTNm3r
XCMpiYM5CVrf3OplTkqYrxXR/Er/crBSgWbb869lxL78BiPg2QofGcWBDjU2fS63
h7sd/RHWCDcBFNmwhxW9Pen1g/9P+RqTQ1sgow3RzgAtxWQruockXjC41In+ekUx
UNJuadQR6jz0GM8AShARMm1BON0WdOQBuoSR7O4o5SyNy9v2dDQkhAib1D7S/Q4e
/hmHFTZYEr90HFc3KqyL4RvYapP1ai5Gidfp728wmYLwSQd/paNE87/2ZB7GizSm
tC37dWWVLhWIugnMzzmcJnJr1MTBRFegD9SRlOupn2Db1JOIJCvsIGIlj3u2cAaT
nGdz0ccXm/ySTf1CDvIEVWA3rmU2LYbS8jG5kixQUMoDGRRcUOF4Ng9O1FpLf4i9
y4rWMThA0TZPgT/2DF0NPyeVi73Hb0XjPS59In0AbdVAliExAmvjAfXLZ+wX5xll
3x1XHMeJZGUbS5Dh/lC3QG1mRVxncDXsdqWweMLblBzmtyon6Q/b7mOCe3M6N9pM
/IgvgtUaSqMXdXbgGSyY/EH351oXwTLN6Zgd/5USBtG3jwcfzzM7VzB4wwP8U9Hk
Agl+lrZ77C2UktWBGuD3ZT4wc9wbUP2/+DJIBz7o5MokhXun4ZVxfqUHSw0wNmTs
Jk+mLRK/J7ZHsK/Qf2h5PtTdw9El9wfyZK0HKCftpkHa/riGJiLQo9liC7r7Y0vb
LCzLt16w8BJkEIxX6C2veFqi+HGfmFliK+U/eBtcjTYbotdunSWBJjEVn32rfqlQ
u9SzIqIk9cKQE4d+DpetKMA1iRvD35N+b2YmvjMsN2p15TOzy9w8Q1lsOgt9qjxV
LppZxJ0mfgvHsX8XMAVJBoTB9HtsNGyTfZqf5g/oFo+fvdEXuNmfTYFCpy4UY5yo
/3e0ydEcaTpeIt3ap6VrOkBnpFp/pqVwm5nGZPmKvf1y1EK68OaCoXjTa0nr11UP
lIWGXI6EYgPTU47L+l1V3H+sOy/q1QhDPHNaOI/vB+F7+x+eQfjSj34AaRSyq/q4
JwpckQQAVUxNQVYH9xvmIYGLzBVplObWMNJEjWf6ZK7ELgnAGUWNG0bAUN//TQ8w
A1o3wsUFJaTO+mXMTYyyJGA04aP15MLNqY+4Wp4G0GP0RSwO+gNHH7Z2WO/r31YW
o5PoUiiEokkuWqWB2YyjVWMhe+XTFq5+K2e4aMkt9TS/+PuNoSTb9t5qAJdkSceX
xd327DWGEMEYJ9j9oG9fyG+wE9AmgX58TirXJ4RwEIzdp4OtIwwa7dUCUPeWfQa9
LeuD3dbKULVFkrMfvg+vh+xKCydrLRJy2zFBlVRNAQP1XiHFXJbhEJOvjHvuGjyw
9AwF1WxkLbhPtT3UeoZRmckoJN+Gl58zfvSpkFwXRCjI69hMOTM17RwKOdlsu2Pa
nKAQ6Es3JztebeWZAF1VhMRcpiXEbCvibki1Q5oqhT4GiuW0y1dcqxUhCf2Upch+
RXSxBsT1CpAovFd6QjvKDkqt1cXnme+VC46zlbecl4tuATgEVvSA7u8/ng4+QHCO
bckjPvhuaAkDQMAyc8kajiq2cJsB4q5myNJr6jGfybSF1kk39DtYXBiVU6f3qsS5
tM2XvNDpACPabfccSsOEBcall430CHLmQQwXNoQGseklgSr/u4O6mFQOCBr5WYHW
27soQLE6bdhPGSJaidviQGKGV/E+TGvuNoUlQOy6okPjL1Qs81JpbtpoGtCfDz+5
Ja2EqakzL5QUn0ALK0IpmwFz0FldQY5y649rKwxyNOjscYnk6EfdAYApuwyEujlG
1qTfPPNZuUIxbDrbLJfW90UJU0BTBfrcdEM/eV1CzD6AnJ4+etGzr1U+04VZC3+Q
Kijbtz9lSDb43ye2GH1QtQBsX42WEFsRicYa50j6M+0hg/mjUTxYGfMlySv6baim
K7l/Fk36Nod/OxpNU/x8X0P5nDCE5O4dFUQ+HidhI2EUeTyl+vzLzaWGN1K7zDlI
ds92w+1dkerCXUbeN8xemhIwTmWwEBucKRvOCeBm3ogixR/ywdaIJj4abzw/30ZK
FCfdjViN2AHkcLIYHJfQUvu4avcW5Clz7WXl/CmmiM0PszIoEFJ1rYhSn0eDJTSX
opIr1EaV3haorOMiZTuuP+q/RxsrwpZrgbk9Pho1qp1DDw7anI9/pb77ts5NUSUp
bE/FAgySwTrkZt8NatXtPoSGpPn5iURb59NfXILFYgLqlwZhHCjSYGna36bzBcgM
IILS3wC/2KRhWtS/XeOnTYzOXpMT7nbYN4t4erOiJqEIf+wBKAvL3tPDZ2HjQIV0
Q91bqmPxIH662wplx2WWm8GQdJGTFLf/AU7V9RoqyK/nz4mErrNu2diCiLdwUj04
MWS0FEwDwd8HOLG23LgH0eV3+HXYlm0BmCc0r4/5UCxiB/yX7782ywl8htLj3qCq
eFf7etJNGqLFgeUpT3Zb/siSlUKbqdSX8Nl6lT5lik/UPm8bkBTYsbYi7L9Pt1BQ
uhzbWdqr4T3SDdYNLwBfmuMic1560PifgJEi88LUfLGsMFcxMLOFKC6BDuC/bNEl
MT9opuiaiq0ZX2hwx/eFLipW9YGnZYW8YbENGg/DVfZRUSVboMtP+m2iArKeC58r
1pYOVg06PjFOOLYYVEcUR0C3/14XEaFPOOrwf6IlLpikzmR5o1wx0IUDuu3+Ap9H
mIT1P/1WAT/O6OzCwRzB0/ulBqrbCqUNh6a7IeXVhDHVsMiwdTO37HDW7VB486dF
JxF2k4DQuAsagqAx44bTM287xiQQpF0SmD0gcE0qxk00spha19iAC5UwLnvVLN7Z
zpQAY68SZD1MmNU1T9lzBJQKMbmI4pCsWw2HL+eeE+ovp8AZFn7B37R75g+amHoe
Kn/4DdFI8P/xnrvhufDf3b9UxEF8Ej210QLQZF2CwH1gc29fpEkqBXQ6c2FwO0Hi
JHRjyNplVJ4sFFs0q3Caj/mNQOK/Ly++u58Z82ONvP+YbwU5ShH+XMsrvs20v31d
NOgdwn0kQVzBmvp/HlSzyLSMlS0CX/Up44DtGy7OOIOklf6b7pwJdNC9cV3Lnyqe
cHDGkeMGwW87t4+zROOENDgwoA+7UVSceSp4CTZfdYLAbc9HYHffV/ohGkXu17VJ
EBKsI0PBlUIaQNv4oEIinNC0ZxbIbCmhe7T9ZzbBdF5ct+bmQ4OkzsnXZfLAweVl
cbVm7QDDDe6j+uYslIXrFO+rCg3RYY4qdHJlZp/P49QhY0fpf+sMI+OPRM5H/3vh
zuieO1x+Vb4LqH5hjb37qj5PgKxTVqDDpuUxwA7tJFqmLkRTL+8aU8k/zyYn2Jvp
LI2WkCapV0n5J08LJfqPE5EJITBI7l55600tcD2Jg+QC+YaKOHroIooAkLn5oAy6
zxayjT1fMwxtoGbBc/0niKkOQmrCtnjvEf5G0rAyusxArgdibmd+uCrSRNrViRWD
uZ9p9/0ZdpS1XTmYHE+b9H1AN2c+lI6UpEhBz2FbQ4NjgG7PCVncUWhPpHnfCOqq
ik3s6DbZXMXplrklbD7qJ1OVK3TEcnOo5sRjMSA/ZR6OntV/MvQECE6haQIPE4ui
Y39mwJBgMj+EOFCi16iHaRzSSNbc7aH+Toje/5YP5UjMx5C/OP81nI0rVdu3Qckv
LHio5+DCKv+N8gFv5aBbxUYXryMDqA/5ZaTp/6DgGUxcTWGqfFugaKdVdPtFT5x4
/cPlasJpP1ql8Hgi1gSCecUDEapJkeAv0AX1llVY6RgAb27S+3Gny5taz1xSZNqU
xNz22rGEPZ+R7wrNQ7A7Wd1LwivQRsjcLTOe/GsiZ0Dg3GEKuzRlvmMhQPI1mftS
y6P48FTBxq91POTB7/rRkqtcoMHEFJCURPuxFpWUE95++JRgxwaLpAKF1tcJBy2Q
vv8IwRfKWNLxk+KWBqZP5wXXCeHcDk7r4K4IRqDFm5qqmk52CnKPgoKlVZgpmAvR
XdHTkwWLszNuToSaBhxb/nI665CxwaiZ5do8TgeRbLKwP1vWoT3zf4HwZJXqy1FH
xkjPNBv0lWruON98bcNUEAu5+FUyGqIE6PM4KIJPFKjCt48pIttRJq4K0+6/dzt9
1QeD0WFeLrdTBvexY8S4GoEyafsqekdFpQc8jf+gGT/A0cJq9wckw0EhlRqOWwXu
FxTW0dy0+wHcppCYjFkwvjbZAgBwqY5d+YL1IMPR6WecanqXej0B4fywLwfUISJq
DAek1tUva5xYcGGZSJ7y14VUd0DNjAxknzTxIV6pdz3E+vjNoC68r6gRRGxYcpaE
+WLjMC8mM1aIYy8y2YfUgUxA1PMqcvnUXHCk3rmqDv8NJ/MNPLkXCsj8kI4ONtcq
Tzi420q1eefefYY20hDMPN0sUBWJRy2rnc6acAtKeGKaJJF58Z3hkZnHzPhzMJ3c
UVbBsPqOPunMzNvo4SaejOYtQI5itwv3L+vnk6bkl5GWVmc11kSUdm4sLkPl2zEu
HsHue8+Scnj4Ger5/n0zQliL2/vL0KVxqhFQmAH+ILj9Decuhhzf/4jbrIHjDgk2
K9A10W4HfrxlDyiVFmPcDS+4SXPK/0UwoWKSGqvLFGdxV6mEndJBZIaSc2sOEDj+
wjKMGCH45J6armnkgCTLmxpblAnkWA7+TXaRGibp8m4sm/yhq2R5BQug4V2qFmg5
mMwS9y3xXz1X/h01Ow8n1YcbDspzluHUrSk7v7WVdcQM2nXo/ZBxNMLYaqjHdwv7
+0CdnlOEB00M8AesQNEG8IvX5IVwwMK0BE9Ug2ZeOEOAQnauIiXZu2mGrlqtexne
DgvXbPkZlCiUcQiMnl0UmUh87LcmlKEs6TzWe3H+JVYWJETC3DZLRineA8Sf6Eqd
nDqXtlqD6MbEVX7gxmCDurtflBCUykLPUwUGWpi9cW19ESNpuCjnFw24oxwPcq9o
qE21id/aHxcPUkUy/x129iZVx2L5qo/Dlpo1A/rMTrbHU4/wmLY3GlIklHdnWwzB
fM4aj4+Q613Fa/pOKgTjNxTAg1sJ2FM619V5RrddCIZbJSGYzogG7s0uJSV1sKGZ
ZrlrbDqu1RmabcjuzDSR0XoJFhxvUUDKM2sKxeb8xxilUZpOsjBto9Zc9Wuf6Yjt
5DrcalJMGKZg1kztb+Gx2wpxtDFitSpT8Mt+IRWRkRXZfe1bdhFUnSF0aSsJFvg8
tv62SDnoA60oed24h3tDgwDGgBESafGzYmYNqkswEIqtWlNEuEuhLtPGMOfLtFKu
ama0qn6kct23pX/vZ6TVoy8K38Y+pKQ01xAZcgAyh1JELJ6f9p/1pA/fWsK2gmBs
/EM6MWGCc7qWIN2Xgiw/Ja/czved2LFOYkpmLfIv5upE/FvpvY/t76RXQZDZk/lk
9DhPjZrLVT3j2hweX7uyTrrwSWIjOlSfqCyTX0r5rVw0qMB1JdKOD0jVtRhdGC4+
OJtj1rQ+fvwhZEHIa4KP+QPREc9l8hUBdq6EMxiEv1TBJLaTwlPpI6tPN12RQzxK
xx7UyjBBFZ99hQ2vLQ/C0tPqVJG+yVhfXk/mtPVKVHxniBmV4DxOXxy7jG/i2ePn
7VJhGk699oUpVUTRbEQ+1pj6kpJoKB8qHcSJUyxN+dTWrPC5McxspCm77F/DwMtn
ck9syiYw7Cy/BolE4VEAtwfKPAdb3kcCODa84ISeIq+R888C4dfBNuieqHyFP2am
0nkOYBGshDpg0XG1+U8Wkjo7K5LqNv3vwoKxGeL3vmpwfuzr+Jy1IxM+1RSa89rv
3u2R3EglcupweUZdpdEkDtt0mG7SkhDCQdMompIU6wFxCZtXM7sCGE3YjXLFIF+3
rMYBHRLDJUD3+geA0/AGVGJTtyO3G5zFgzyYHvYZDEbPCmNRUGhoqf+jM8oNISfO
8M9FMMIlYVWAcJyzdZzDrziF94KV4t4LAeHOvUUgA6cSmGqT93AaLBAUdW40degm
YgsQGeEdkxFbsZpSjjqykCUMeSC6EI4S3YSYXl9dO81gkL3gDnFF714ULLcZRXfz
RrnlJ3vdgfLBhPWZVQrURNKjQE2hUNgZIcjdt01bLkfV1FYKeWSBn4f1BgAfdEMi
zdL3m5Jn7oAnvpB9qriRyNgaA+TPAUt8H3d58UizNtF1LN6QQMoA0Ff+j8idHTW+
pH494hgdnPEC2x8HBek5UUuwq/R4SiKAVmpGaAbeKbEp91o7Y6cevhtULnWZ78Db
FJ7EH0n2xOtiog4Ga00QHMrVErdbyARv9IlV9tFJyA95EPMm009wEoqatCh2alcu
oaVQwWGf5n7pe0EvDSTFJe4ny9elpwmSUXjfuYW2I0nY9OfVea/GDqNdUzKq2QYX
Rzxbt/HBYCZibQd+2F58qdO/LBH36whKIqRTTvXafkNlwQ4lxh9TRbs1+mm8fjk5
yCM5xLQ6oTEcOJm2zJ2R/77WvvPeDdOaD4M0Ryo18IapKMIcn+RLO7JIsQMxdCbq
ACWIp85I0RHAWTD+xXRglpwecHdypxHX4dKjG1a1eGuOOXC/NnXb3hu5MCUKpKwT
LUUNNUcC/Aun4s0uRjNHV9UebjES37swzqtAdFK4DCf8LuBgYyDRCO2wY56ic1LT
6RExYHrOVvKR2Ge7C5+e3JKfYOP9rVMTiACQaWAxGP1WkYNbWJJeAHafzCbkUg6C
SXiJ/jYbWEP2yD5IevI/FPkbnX95C46RFU+xfrhGDkORWzar8fr96/IPzdCUMIGw
h7pOWlA5wTmhZIC2w58JnnJrvPa02o86Q5qNKUAKR3NoLAzI5puyQxeQJLMKUw4X
Fj9bwVmYsX5i7CIy9LaBq/Db7mu144v/nPp3EqtnAIbO9BK8z5veAzwpehXssQGw
fO0G1NnHtyy8d34eaEKTbcWLsYCHapBE7lt6118j83/A6T58fwGlT9H+5qHbZfy0
bPY/mOSLRV14NQaIAGTQ3nRsEublr65Bfh2iDYN0wZKwwQX+KFWvoJwEqwIzXQM/
UeVn7CGy0QxKreIPJxJXObWjt0ofjbAeTqr6J6jcU+BD+RglNY1s3qMRkJiJD+2s
xklVkAkY80DYQO1nZkMGuxHpKCrtPQDKrNOwQh1s+KILpvl0iUakVUetFBLhDXRE
AbTCAp3YbE8jAAYaoq+f1mcxpBx/XWu52TcLyccx9ZEVBz2Y4QABAiPgxib1ulCl
XfhofRBptdiWhxj/2wkAgFKeM4//3PllKWQVb7z9yvt+kRznEswTJp3GeZHYCZIg
v0r+lYtVHz80aaOGSJInYjg+J2F/nm2lmMJFdTTTUASpILo8eqe+bvLNa5ax3hfd
w1RJNxl0tdqgm1o9ewhroOo4V+e9j6o15Xzpz6blZN+4xiqlQF29z9Q3+cTzVj2L
WBYL9XqrGgIB4SFzBXD1rsYz6NNQPdY1ixwXQQUb/flLm79cvfZ2Ps6aXDP25R49
miltyhsN4lGrkqn85cShdnufhDsj83+CWJfKCxBnAFCCehelweioO5znZeckpwDa
R1MU2K+c1oxblIXd9Epv1sFGOeD3v0vS20OMD1cqcRoD3PwYtgO3vzse9OjtKcHx
P85P9/RlSkgumXFyb62RWRdI0T22fXg/Q6Mt+Ntza0MZXFOIlsio/WSF8waizB1j
JVr3jywW9LViQww5U93/APE8uDZfc+iOJQm29siDvI91pMEygkQm2REW9EC4weBF
sPI0AyuNDuj98zSaxrIgkGZqRQ4en2Xz3dRBloU12besZttX/toTI0XJwynEYYt7
vk/ETf8+vBayoiCzIdYNlxuzH6p4dEXXBrLL4G3lh0RbwMw3U3wKDdGDvcahx/rq
S6l2gPWlBsEjBmW1/9U2ySofggcGRFGgqBx7MFp/G9VBmvixoVSnGmK0bIXRuaDN
zxk3M2RiJYH5B07royr2HrT6+q5WmWeoqvXRGA66y8Wo3AZEnN/v+mJRJKvCCeqZ
50etyeA8JN+RLgTWgMSzR7TgffNcL6LySib9opHQVPK5nSgFTNqyA3gDsRjmTMvP
8BwgWEkgZnXKWxO4fm2Ke03ajLwQCrqjkzXh0CycaIrU9jGGR9HJdsKOJTDIWUw3
A1LSmJABObcmzV0qoJ4ApzVS9Jc520UdPoI3z3llmLmpzIT2pyIi4EjAr3l4H7Gd
VzaYqOMKTUszUKDunvHdddnSpekT6QN3L8d9991adY3T+le1PogkU4zr7vMJsv9X
Vq2zwb135Z3/zknhsFdUMaJV54kT3S/tDjy20d0LtMVNsA6d7eWhrcGW8LuxoBql
/l/pBuw+naCcaPxZprEKoi0LXipoD7u3w6ZkWActFUwExnsljkyY3DeI3rxpNdX+
VgyE2flKTNjjFRsQjjY2a6WkzO/zpgL6F6wR544x81V4+WIrb3s+oly7brv0IDnS
n5AeWRhJ5y6pjjBPpMVm3o8kapE8Dx+djb+dzDqL1SXsuI6YXk9/DtZIVVfk8MTl
eicU66Cb7bHJFBcawIGnHRF017yzlSgIghdR7uf5U5FWlAXc0xtiTKPGlCj+8VjC
kuayhxvLfv0M6Dr6SMJ/EF00mpzthkKV35R+DUU1RakVPwXPiuc8f60VQlkgwPVu
WhZVdrmVai6bXSVNjgJmhz4trELQwzS08aRCpABHRTlXhI+P+xZpAojE2bSrZww8
LkAWW4PaphCAdUbEumh7oFlIkn9jKOq+XEG2Mup7FuyVRGB+4hdZI0a45wzM7bfD
eyNLdLLGviyo9XSCSqVdk7BEnAlI8sFJeAstcc/DCrupOoD3fhOmT7EzwY9LHJ/5
nSklCJkCxDr09n20SmP6oQs5amXNfmJY5X//7EJ/rmv0c+gowZkIc3FAeMleTM4l
Q5MQm1vhjh5YzOsXkmTmU0MrBrz2Trt7v+BFwTd65DJ6QPrL/VabjF6PW6g98EfC
nfJgcAsAcOrshum3jmT7Yjky7hJQ2zAr6NZnHuPcothehMHWdMnL7vAgjPOT77Jc
/d4u13JKtibFPsbunqhWPWf6IwnVjttKfpbwcZxfwB98wDdulRrHkHNiCrab3YIv
pmdxGCqXfhST61qEUUvwj/HuVFXBvM5kmy6oIn3DH3enxNKyyBB1B9S14Z6RxP/3
c/KGRAVzGabrC0FeAS/CDnqH0wRzEtf6EsPwbjtFRtDsycGguZu+HgEd1g3s/Jm4
HAonsA4hPlxDv1XF6Tl6Py7AEd4kkk3LcR4zw6TPCIDoP3OASTWGWbz4lAZpwVTy
En4fHZIJ2vWKsHT2xnR+jUbFZQIYsdxm/2HuCQ8xEi34ahkzPH/+qzOeWIRIBmIB
Jd+iXhC4eZRoqQm+6VUZ2XgHnPi4RYyzrwukL6VS34+j5D8+IRwdt9VqObVgp9kq
I8KZvrkIEfutjmLJ+HVG/lnHmBunr3c8bzJsdfB1wVuCTlIBEILzZw0Djf/NtfuL
lvYGKZC2vm2+ZEEeBK/9p+L5wTRPuCKXstpjXt8O72ez2SVZflMZm9l9GwW8BoQo
KUOZbI8b4/cSXVF+9n2GSR3dYH49f/PG1H2hxvuLUJG30kO0v0rCSLfeYpfsMeHW
HgeMsrOjqhxuSDHhlmk19QYgelOy+Vfb7fs8idh4jm1gGFNHS2T8z/zACPJdZH1v
Zrm8Bd2RfAq4W3oaU3/yfpWxe2nIHE6jO/9UTNaB3oxZBbryJ9AMRT3PtuRGjeYx
bozHu16JYOIX7GUAB6h+hht+aStvAFYbRj4nQx+rVs4KhriOty9O4FmFdZCu5td6
NkMGJ8nxCSNONsFqClmjXdYop7CCwJcFytjlHwvjz0oBGV899kzvVsnPJaZ4ON0C
/BZlBF9j5G7C40u7v6nEaKVS6onM3tTMc8LZzD3jdbEXmPzk0/USi2Jv6Jj8Wfkh
VCai0DWnMsi4UG0MxMW95h7wJm+Jzn8Cj7I2IUO6c2L8hFDpJkbQ7+ozOCOv9WPC
LX56Ggx6j6ya6yYtRIVZZRQTGgwGH4yTCWtoMx3m889greibYO0n4Nm8iea/81pk
ZN/UY84UA+pVY3RGvIbCA0c5uzJg5kGdI66JXQZCfcdp7UvPvr4Yvnj2Y7RHju+5
GKuoU0IZ/aa89aH4fpcVvEZfg/+ifTgRcOC8oWDoriqgAy2FjxJWXFrU8VrjIDfQ
c0W05xmoiw46G6pm4h5jWacX85NsJnLG86xiPuFlOyXVjpfoUoG9PblyU4gu+Jd0
FJH6DzpI0IaW5enWc8P/z04vG8FuCpKY1cXP43KzC2CFocernw0uBkQ8yT7Gr3ZQ
EASi31bbxM0kEx0EEkjnFDRJ1Nx2Z8ZZp7HKr6WbIoE3Djo8WXNk3lNwTf9Gbbm7
dU5n/LR5QEmnRfaI7/JeLCMcDyo22ClZa3+TRGDLTKHp3NOMwl1wG+whQRaF4Dma
z+kPgyEerBGPpPhFNEwvL3TnChMdQLTGKpAej3YnIDVhCmK9Qm3aqjRYCjD+lBxt
mHFLDoA6Td+G8buh2vy3naqjMM+MN/BsurCuPotVIutoZ4tEiq8+98HbNfC6Zqmz
VLnXkqTOLODJa9MT2v/+pmMSbWUBlx1QEWNHUNUnx9r7eOCFMSI9nOnyP8aKngwg
tMCFJZ8+t6T3EMLj+Wsdvly9R46bLcYc5nDkEX/SnMFwNARrxVio8HwvJpT++WII
Ne+cdXYMrgpCTsenwAiy13N2Mf+U02RdJUasrJK9bniMzMDcVU2caVa0K3pSPqaj
xx8k/7ynkkzTnUnjGf4/cQgyP7DYqRSSC5n66GUVj/AEtmbtcAu0ZeiLQ3aw2XBe
MaQEF2qYoZAYnUBr9+SC9BGfJWNdfWt6aChk+BIY5HLClW8rIivQZBjCAsCj7fRf
SrN0LrUg+dnwBtV8rGeD+s9E0XMAk3CuDO15hrKRbWRwt0rcU0s1RsY+J+yijVNT
1vtpEDc+t0VgWeF1TqQLD0L0mbBcQW8igYfTXxJ2NA8ByKhmhEK/3Ve1BqvSCNUb
leRmaCn48TJQu9pr+N5Z5hvI2Y/ob0i/6jMlmYiPIlTRzm0aEEGGHDyxgnd5FADj
DJ6O9HJ7Z7q6+lWS0LSpljiXBAWIMGtxowRk6ZJe59FiP+B7p+TVgGRYdLDvuaRh
RZJnmp9VIeVwA3jqeG9hBK9yQpo1LYOCPvg2Hj/WrINEFSuVua8lXDx5CojrqeSq
2v4IdwVH5vXzCMb5o/5MHZLo2ksQeZDgavPH4nCM8vDlZmpMhhc8axMh0ZciuV5w
TRTVosUY3Kne/y4ZYdOqoD3VgYQ/mRws8i3I47MV3+CQHMJBRygQvN457PieuqDf
dIw2dqjc2PDfnAPpBNewsfTEQWnkflKEQFVHgPiHBi7Mnh5IvBXeOKVpja4cJs/H
YRKdkTrtuUUhd7DZqawcskZXVMgz4c3KuztNF9dcFrKY9NVxx80yFRem9EIKj2Z+
bl3ui/G/YstTQrRRG/uylKxwXF2Pq+gQ7XMp6/4stQQzjUmTnzi5IadOtyOq9k/H
ClER9SrRjGLaWqFSGkF3dvmnWqcXmNElgXWe46zbAYVytNy+KYdt3DXu3r602CcG
TVo1Zx8gCQGgcrkATL5aRfJRlxrRzJx2ATSmoRJWfQf4V+/OPKcWzSPKg1MagQfC
HI+n+gXAiD4kT12juGYot3BZjRU/qulEJhnJC6iOecwlM7xZobfHLDdvXm9366uP
UOiInZcm/Wkd38Dqnd3RT8D1Z7heb7LvBXuHyn2ZuK+ap+eBxgFI0bc9N5MAJ1fc
ZjXZtIF83zl1Wt75qt+QDMZh+zr+RQyU/QnyL5uRDkZ5nCrty1DCWygrxrkYGtnX
fpIxyV8ez8ku5mkX91KZbk32jZq9rvww+moxT5DZ/4tsJWzrAMrbE2kSjBnLWbbU
erlB+OmBusz2CysJ00JDT0xJXHlPwUDJjSqYkCxIwLrvVfueEOC+2fMVqjZNku1s
caGy5oQSOtaDf4oE+QpP7gtuHogaStE14ULYlyaj14KSXQm5cky9q4HtF+/OIOZZ
h1OmQ+I2i2XbPOa12oSIUttXgI2p6faSB9KxjcXLaCYQ9SgZPqlSsIfxlHHV3FVf
Pf3hK6XQhrRSogvMpTR2rseTLOb2B58gWEjysZGVwi/pbhOGpZgzOwn5nA1yCBVI
/awtj84RzZXVp4sAkA0KP6Za9PglltCb9CaJtf3vRf+6EaD1FVb9zRMzJxWUnHeR
qbQuzcvCJTzS3tV4dXItu3263BYlXVCJVTnZqlHRtf86lHpXEvB/EtnNX4P7G47h
22LODWw0eFBSbdi7DVSK4Sr/BDHlRinIkGfxWMBD9Z7JS0hhcctARIebXB7WbQhd
wTUHZ1Y8k8sp8X0wSBiE1EubH8hNQW/rPQlO3+js+Fd4a9hdFYk+L4Qk2FkV+FM6
UjpZc+jSRVRH9qQn/WgUYiCwdmMG821ZyDNhDEK8JS/HBO9PfB4iLV1Kf6EJt5IF
yalI4PrNTmkOZJFOv8nIP4XiSyzQsOjn4CeOgwX23k/HjCledtjXpU0tTDPE8moZ
H+fYpX7hHLfQF6C2x95CiyliP7OeMWXnmqvD0oEtF2g69SwmpNc86oXL2fktC9WY
YWvBKn5F8auwYDPIa29LHDiQxoFU+8j58xzoyUAKJ6Bp+q+Noe5sc5qdNAcHOEs3
90XGOEabYPAM7VzZCDQqV6FwV91UBgXP9xeP4hYJP/uiWyw6UWP1wovlJQpZC/LA
mnYGdvs3UitoPgZ7Vn1xObJwQUxOeWUgyKaVVZLkDf1tzYRLxgxyBdAqoVwqQd4e
JkSjOmI1K4J/qW0Nj8niYAkkxYuJizHyQ1bes+U0sqRiZVGsX1xkApr4CsO7sMhp
cQI4ltX5QIMjfE519U+ZhcPyE6e+tWanKqU2nQiwkMcxPRPuRIO2IOgCNcHbpUJC
GYeH9aVHM8WyXPMebt7ycR5GT7fBcJ+kf3xHcxE8q0T4hH62s7GfEJvkY6gf3fqM
FTW2o2J8JHiJcC79Ci3MpgsVxVmkp729nnds05FbZAFMrFqEdTjX59qXcytzHqZS
Y9IotwE10j2Ygz2dUvne8/8loV/OioHToWgbHHOUBMj28rXEBuGsb3u/sSCVpyK5
mMjQGayFXviosItB61XI5V/KPcBSyHvnybIPO1WjlKZ3DddUZ7s07EuusI/zarkr
qIQm+yogJGi47ArpZqwJ7NiEYTvxzIsY8xfnr8R5ILKVVOxRuD4ghnL5IBdMVVxn
PJ1PV8Bd5+0MetDpE64jNiom2HouRPmwloqmX78Sg6SJx7c0Wwzw3x8z7W9FO0Pp
LGXmc34xqNxmNoiy3XlUQmAz6CjdT/Nx0oZlsVJskEbIOWJx/HPGhkHKThtGT8a3
zC4PSaWWCdEiFWc0Aa6kU+IArlKtoGpXs38IS7qkkbv5UtemctZZ7NvT3AFHNP3U
D3bKsF1ui18yLcjk5kyF9uOs8HJVXmw+PtZQDZzvi8Ksiltbtg9F30WGslE1/Eu6
J0OPLLIe2e9szpW33gs/WVkYcxMgAcCdzFOrS5kHzO8CSQYO90TCe9p+MZ8jff4R
4F2sWE2sKJoAQBeApJ4foLZev8+xHeaPwLpo+g57xmOnWvXgFeTnwmNC/3s8GqCv
qLWydjgzhDaDdpGWebogRC8qE/HCFIJiEKTmhsmBKuEOsMFlJbgAl/IGpPMc4VuT
4uOVeBuh7QwC3+yz0OXFOekpHvwZ/a5oz0tmd7f2E4OzadswjY6snr9XlklsQjTX
Q3Ur5Qohyn5rlgVVXTVNwys8Y4Ft1y9bz6oBroZO1LnNvZ9OoRNDFTcaV+Qfi7at
Xkz7E5Ud9cfEBZWaJ6+G5hoGCv1gLOrU1Jm2m3a4EGTkqcobxOIDASmxLs+ac7Og
8rb40Ozwd1bugRU2C2irMXjT7QENF0YJ9+oorMIUKu2ep0Zu0rBsrogukFj5PXwA
A5R+CmRqYiwgojnw5EZelaCizjTA+9xjYCGznW68O1Z1Rs3KP8OdlXW4S3TQM5v/
tenAU/OibYp1VeId3WgyH99NqW8GRjudOd/ORQlKLcmI+bdWfwUlegR36HoO4nPW
m9ynfFNJ13YytAbGuODTVoVqgeJcOQ5nQz1zf+acwzQJe7Dje4sjdSOxiS3OtPzw
cE6pwBdvI3w1sNX9uGGX5t3iAdLhWDFbNDJTDcIro+MUe/IVlpsc1XTu9/itdt9J
8S2m0pMBDbKNRJvIjnMeDKr2qyfKoZcaivYAehX8plHcfk/Ccu7y4Yi5Ane6ToEX
qih942Y1hxvvV6ZY6O3CvoTWzLjKczuNGl9UeqCAEmPwz1+OKbgq+FkEwPVupaNf
0V5/beWWMS0ccsM6iKCzwJmpkeJW+ZKD2NaL+z06mMtMjm9EbzWL6xeYCuKTDrgQ
o7D8RnGO9YmBGAGWnr7Xjuwv6oqM1KcDE8jEoVx7e4OKT5FP6IzTlYYMsKykDLtf
saN7w8qmKFv2+TJU5sytaLtKd/QDP4kZCAMzesewQgVOtYRaWs7fcYGS1IBLmjTg
+KIwyz73fRkR21R9UQdurUhahlCvC10f17gcXjIm4D9Q2x4ckSSHKNv3DsOb3sob
TdmtCW7/Agi+tlv9Kf5ALWNBak4CM6cC8ef18XAMSLMhNmNh2e+Wc6dFteuKPsp4
fx/QPdbe34RIbfRBrj9CxNnHnmAMPBZGn6GXskDS9MyOIv6JSjZL3FWz0dwLkTO2
W4uHa4bN6Zf00mf+iWASOnRMQnYFNIY9DYjMUAzgL2iwW3hL3HW5AHf3w3wk5efa
b6Jzu5Y6CIN82c0Ro3STRT+YQ84v5CYNJR3TWS/YAzYWw3NelCCXnsOkluna8zn3
xFwMVSXipbhxXrKd8lRVYduN+285r5JJSbIR244jJwKFBsVYC2puitwRTmjuAaDb
rcG2URK2OARXXCKaM+pXYsHRVNvGRZzD/Iuyxo0hZDi5uuyJahmK3ZIaFMA7GZOX
61vwmeg2aZNyUaNSZmc1NNUm06NqcYt9yEmRy9hlLNCZeWa+CSvxZhEBFF2rn54Y
vFosCKobpms7402YaHQRYiC64ijELz/TXi/EvovvFXcpATTpO3g2l91lM1uXb9EG
4rlv+rYcNJLnq9pp3i9h37uZLa8R1kSRGEv52HcNlCyvt08/stizaDWCn6PauM32
NJgUHqhrDMkgKt2p/U6sRbNL3pPgBNd+Aew0ccyID/TMHz+9LOObZBIfUDBlowg5
6j80lopyZwY8Qn3OiciWYnc88wpj9aj5qrCDkn+vLacwEEh/hMqm//TQSilzd9uy
E7SiYe9APZbdJ3P/Ajb6E1ShgEx42PT44u3n8nfkU4t83oto79v5bPBA5Ci6Rcc1
I4/9+Utj3NMgZfbi0kX2fID729R36nPrXXRMjL+G7HrcdnzDkas3/zaI4gmnmQQm
LGKzruNxrJEkv1yk6RQ1VCY/4P7Z5tLUa6GO8Alv65DMWEW64vTIMXFQszAIz6SG
4OiVfZo4N6mTvQuyjHdkDkBojZv8CmfvOyK8tx0awSbMYMQ8pgNwVNZ9Bmwdj4wQ
QJUs+VtZXE/Tm5NOrdqzNwUKzApIQvCLlMFKD3Z2zT7LvKzbP72MRjTQ+DjRrsbG
3R/Uymj6phhe3QpiiKMFdBO9rwSPu7mINJq2DDFnlCkaiEYqtBkbXvm9BRZmeJyR
T0RKsCwqnolZEeThXxysuOdV/NUaIpxgFONtQHOxYutsk8KBZMQUPSIjBQECVx6w
drNI4d4kSa8lGrEI3hrvnCZdgBkKbb7fx4vOM6UPUOX5dxx2/YSE7XHtN5rOp/5D
1hD/2FpAUah2tAyjx00yvQchMJHhkAGcDNiH24nZUqOzB7RI+f9vANCztqinCK/y
gwRPBW7zJ06c12YrK7urclZIJ45jXSj1ITYniz/bYA71pV5dfBNTbYDxNc0I5gLP
ySsdHZ0ORnVO2fC2BLHM/tRQ52eZcjh5YcPEiNX265VcqFxI9cmZUjpH+gRc2vPi
C5fu2uAzA/UiIBzTYGQDXuRm0BSjhMLOqYAGZj9QShigcoZjvUItA8QX6R6UQi+t
gIbUcfMZ4k7X/+ns7GmUVey+jXtfbjl5M3Oo2fTCv2rUBNBop0uP3wkGHLYsMeWT
9tdEwZK8AdBiwWjIkL6hHkg4uUTj9hv7UUsoD/wVvjLqm48wVTNAqS6+3WW+wK0l
iKcMpG3N56C1hG4UnPj0vDss9RTCZmIAmzzKSnBsn/l+M6CTYNadPqa6go1FDk17
WvqjCeRzSDn22MeAt4XKoDr/u8vSLO5/E/QfweiBrcu3aSymUVN7BsRFZwGP0KPs
uW6ETTcF+IMBkW1Kc/utmrG444MVP9gNCTMC5w/+tGs6IIrKzEOU9mHmtqVIjcRm
bh6kzIr3d6vvlW/gnDGnfN8n9KL1KUvA/P1v/jlpFXyd0RIA9viaqvggZh51Meuz
iEyzx/8m1gjECXf1IUGlb3IWYd4YAqVEewQyzKM++qh57rX1e9QB03QJKs4RdX0D
UR/7R4/BQhMbNXjKihCPqAyCdvIa2NK80TjG9MoZCsiPGNZQt6ivxzBK5ClQ2U2i
NDKWfesPMNc0UbFPK9wSlfN+R64EOEMsRUBmjhufIFcsE0EJ2oj9E3gyGM18750F
JRPeIURap8qSnFFK0FudrE1B+gQWdwrcYFoYvbLElO9jsHA71dwDNPCzOB6eyiBP
+QQF/OiIfdkhi5AoWOtaBrNiqfniKogcErW5RcxAwSrNFuOT/eQHAeHAxn2Cvwmr
b4OhyGYKhf3PHtXnzG45ASl5zBI93dpf+tlpcsHP3I+QN6HCUTgSbm7QsTTlNsyZ
c5iCA86TVY+aQIYH6w9ptg8FZHVxlj2tRPX+c+YbWJ6bjzqA4KDYe06cHA77ADFP
iNqOebs3IkeiGoosONrITEvlS0Xkuts4JIsO0vH1HVw0AhQGmXrfW9o+YiEOhqXN
F6kGtHSlBb0gjkZSIHeVDsVL0RRVQ5QQFWV/csndggy1O+r07687Oes1ELfhbbVd
42V857Ms6bNXMHJl8ViNT1rOjXWOrtwtaEVxdmyJByc2Ll+vHfGXG5O4Pb/2qhWk
os2D1skoEKCG472O6pA11mo5IBmlIP1kdHIxXPpDOgWyitP7/Bpaiq+3Yy1JXSfR
lUb+njWGw4Nwn7rzbukSyKV3xYFVIgrVD7VsDv1C/9E1k9WozVqegNND1QmP9olk
BDXW+DOuMGlWewasnMwooC5lbGcZCZgMCl8SeW8BRZO0+62DBH505kUeKkF7ivd0
PitAG9GjQki99JFe81IyzuiLz3NS3Zzj/dZTMrWX91mx4mQ1uwbcNcIIypF/6TVc
qOcdOPiBXpXf0qXtwInn7T5DmSSzsD5hGK+2HKHYnXwEHM9ZT7mz7+MzW2w6UJDF
k0lj/3GxaSVvEMwk3Pa1chAZiBPW2y0Buy0ectU5NWj86/skZIMtSoawcarUfFs3
GuyqAJtVItvTXsqU/Mpm2/luKn44OWQayb3bPGyUzDPUWHYcDmN42noLBSMiQuaw
2uqa9wsqT+SPGPgFQBgRZepU6XMgbf4Ovg5ctuJONvMhp56EltSYMqLCFn7vmZ/3
QXjFpSrsl4APgsh4xfy4DnpVjJdPzQD0zyN7GLB0mD9OVc9wibANBPlrsYm9aMfo
01EIpO/GobV/ZIiApR6uiArjhIDeqMVqersXwKJd1wHXyLiHO4nQXDIkD4QVgxky
1fm62RpIQsDa5TWdc1XcUkf0mCr/jgZRGO6wcO/wVg21jcJabyL60OpYqpWX7txj
ttgActer5GN1a0ULF5Vhzt1PFcDJBpG/dAMVoG7GE3/ukUn3kD/D59B7/2xC+mxI
8aBsOMu4Yw84ygZNNMrDP420l7GqPEjkRrYh88GlkQYylw8L0bV9gBSJxiQXmN3g
9s6JFDZD80DDv35oG6JsUK5AC+KtCk0VZDKFdL0czIQh/LX/zv8yuCzHD3qe7j4J
GAKpZuBmZsSWy4z5vCUm4VDAl2ZJRDs37YfpIcf7ORUOwPwJqoCVp8o2sa/9vEQH
2DSqAZx0qhPcxBKEt8e5SBtgHYXGvkJP5YKFpeNvo7Oy0zmw53VZalHOBywnWKaD
/FlzfRpORfmu+6BH2Nl6PAL4KfYf/LqA5ZHPAOtqdCzI5OWto40jmbXYykSFEn9Z
OvLmU1ldqP1RSOt3msQQLU+oaLakvVxIkjqCNRAxYPowv6KN3VKZdVIF9N0sRveP
SgQ5u1dpoaeJt03txo0EMXxUiD13i3e+Hm/3eOtOjKgfQQcN0tOuW6/HLX0+ZFDW
XTbibh9sqNwo5q0W4pMTaI0K8zYtOFA8a5Fu3aZjYIWezKdQXR9imQE/Pb9oJ8s7
ISFcy+V8j4cHDn7Sr+FPIsLyE7oXOLHgMnnyGhuEy/dJvbni2DdsLOngiB/WunsH
qFrILnVUr+dW7i83tqr05CLoxefHIzhEqnn2SNj0LVdK0NbpvjukR9J3Tm9xD/Fu
xs5QnBbDLYxYrGtW+lstu1iY3QCZK3F7jsMUbsJZz14R927jQrlbKgrxhOnbXvPt
mEVLpFrXpbLn59aIDYJ+bGpFhXgKepuhh4hhu3jbur6n8FR1ZUfSHv29P4Rg+HfI
absdxb9oQHPpaP4rUlfrro3BbbVLFESkWKCLX9T0T5H6POXoUCfs93wpAxF2HYQL
07dUA3par6cQywcwKADxh1wBkujfEPLtdxDMesKXjA34mIe3lkQFrmXZT8+q03bo
lLecKd6EkDfez5qlYKfQceAGpvgxMpgzYsdLWUAJGQz9Da2Pdg8pduYsYmDiWToX
G9LTvxeWbbwR7FbrTx1peZrgvGHnaynKfEry5Wqa0FUFNrEyzDZ4IbcViyoksuO4
ElGgcrd5jFnLrcvKhUaxv02gXdVyrDMLU9jjBJCHSX8t3xLdIk209Telsn+iLd27
yPPr1dNga2d9fY9FMmgvKmrBgg9z4tcXHtqbzD0vwSgA8gSErqeqQSDYRh1ODVdt
RwzuE6fnjS9PlKFE9pWSHHbu6UjrnWp+y0E0CKHdsN4bcV7zJSU+hAjUEc3q/Apz
78Z4Au49jH5VXx+t3nHcPvsRCsDUP3yUx30vLGQk94t+cd9ik8VEckmVdWBvB9L4
wHsdsKWcVoLFlV+vACKE7tmr1uRjqKzL5noZ6evY7EbzJAOvtw1797C1mUYfHI8P
1BDky3ZP5eolOddKPbz68+8EN+xocJ8FhukJDKUcz+JHjLZzpj8HN7964ImeuSrW
apxe9Q9Cmrf8xMxgN+Ljc0hanKoVB7JhjS3fqUSn8unlUxnmHhQTDz3hg6z2AQH7
CrZnjpIa499ddhFtoGq+8FKFaTS4cGd/gIlxMRU1jVRrhHln9Xipeo3Hc2O4aHiK
LM7Xf+L5+nrX9u1qU3bzPxzaqgOHKdNe0TPML3BVzX5Y165YtKN8NfY9BYWS8llL
+yDKq+AOvoBiEIJ12mOAwSsyLUarRewQat122wc+MGJrOKJ8Beb3skzEVKS6CoJ9
dLv6RN5OTacgfi0O6a1ca6lcuFSuaxcYsI9h5ekmPfrnIZK8du97EXhxVWDyTI36
+el5dS4GW/QOUYziDV62GMNSjnMgTuU+z9RQWcfo9ozNM/5XB1gkpQr8CY4nw3NP
rJD6YvHNQUO2wrWquL67RNWpr2gijVU6AN3UTOu25hD5w63yCUz5uq99jmraO0Bi
aG7BTAmfR5g347+j/K4AQ0Pu2GGLSWCI8+oqWqu6MPHswe2SVpqJPog9qjhNvjOi
vZZKiID6TpuaqP/MpPWZTLu9h3/ifS+jMV4XNX/3Zbh21+4UkQvcpYzsDmr02Wlu
GsFUVJRb/YAcw0JJv2i6JHq7VT0FDSVwBWV17r4I+pa84PJUqjJiwDWVrtT8E6M0
V6/w9Jxi24lSnD9iVMH1PgobaTiAdbCaMzm7BOx9LUmKlmKwDLSW8yxprusfBVmG
FsKkBwyyMgsbgXMJYkfNeb4XgbzP8f6Oz62sHHbctdkaBQgP/z43Ml7LoneXJ49b
Jqt7nDpwKszO8mWWpbSjNOU31yKOwUFoPUyGPl/6xtA36jradRrbiND5hws8RNcj
a9TM1a8ybm1tqbBmuikBIMbPuMT42FTdtQ2sxI2fRNEHxwthEoNcRkO+wyuqWZ7b
nZW+P/hGyl7N0svrAwdkds0dD8Bcm9KT2ZTXeYl6X2E7OOzpduOC5OMRcCU1djgA
xH4LoYufd5zmLhmGZ3zK0w8zMERhxqMQk2swAa/Op+j+kSMofNuax+tP8J9NEel9
AlH8mi6R1hu5g6+lglX6fyuceC63Q2Fh2xqF9yA1XBZTQTTVi12SxU3C5YhFeK0q
7ItI/YWm9oQkIbcVMS7mdQOKhSQLcPJaYHbwBUahiczO/pqkoQKimsZLjB+X8CG2
43o7Y2TYVfSHs/Lak+/ncDIyufQe4+K5g63E5wUdMisSxzAnDyIopqlqsjicZNiF
hhA52ik1KUmx4LDVicNUxF5GW0yoKRIlFQ0UKKrxuBbQJqOz7Oqa+H39Y609aSrM
SQ/mg5+CcUTZ8xjZ6SYZH8ux4JKT441pDOxcBw836N6OSdW7jnu9PsqB7DnaLjRd
jBHJNv4DHNF1BldrJ0xdA19dd/JByOj+kdH1NAsZHgpiwUDSDLN5d0X3ouj2Ht0G
5dp15NJlIAQz21QQtHMGmqNZepQLjwsUmPJpiIsHzZyIlsQcm+7zbW13so802UN5
J/M5StjRm4MitAYpV9DIop4g5RWD9Tua5m6yhT1J0x989LaDuvR0qef80LGdBIfo
1dBU/cC/TIjbywyZBBAfS5+hg58MklCTIUBBx0zYIiY7uOPB6O/nvfcBCeKUi4S+
my/U3v24/9sUv7YFC2k0dBVJZeDt691qCjfEkYYFgp9vVmqhu38R1ByhOfklAxvl
uPKrrqE3FkUt741W5mSg1GB+fOPH2Z15vKt/qQLenxihxvOAReAz9aUG1+9D1Y+c
lRKXnPAWU88/ClRDakrj4F2nXRNzLyh4FfgveVibK78KgTOOKpMsr5NeoE+LdYvd
H1+/09pr3eDwxfmnkqveClUyCFtoenyHTqHD+LWo0jCPttBH3jN7TCHMrApBTM3J
gFMUn9zxs6yujqwVQuVt3s0uiNEGMFG+l39CM8M9nP3MCgjI7QdkEbdNZ0YVi9LV
XS7eVN+WBm4FSsDr50pQegt4NDw/iedGwcHKjoG6Ec2K2Qi5I+6zR+sdKYDQnPmG
uX0MkdVvhWAAInFY3jwLxL1whtMaEndB/N+54ogfiZV4ZHPqJsrTYrlNLzaUw9iK
FhUiiqxZSShZyRBwFCfKWGdAH0YAlIDNGEHChX4Tm/C9kyN0RVmVVAQXJvHyLv4a
9kWf+YZX5N9YpmigY7VJFMPW0S5h2DOzF5J2LgGOGlhACXlFBtEGh/NCiqafFjPr
HWCoSzfJGtepIqUwWpQoBO2muJOueXdxvXte8ACyo5/pg/kLvQ70vaS2jK7WRHo4
5AQ8FWcGnHGB+0TFSE53OWFOHZwMuWS+iL1H5Fm5mR8FZ3e6QDhyS7yaYcTBw4Ti
db7U2v6KM8bktIxzy5Y2FxR+Q4IfQ7ay0O6lhAvoqAcT6JARnbS1fEDQ53fIIczN
Jld2PtitXsP/411YfU6g7M3UUxYh0q5xXKc0t7xjW5DbGaQf4j9IrjIudflJoP8J
o0QAdsIG7Eg9DN2T43+oOGNS9DqW0O9buaPkiZBTrq1Ov0FgZTVV7yRcWKxmMyFa
LdkQd6OKcTy4L7LH2hbsAkAmaq9H1JQCD+Q59/4hd8oR2cqiiEmPWGt/wqpV0Yg0
5C8pkHGgF/yCaxyKT8LvrDxQ+AaMA0+QrL4LwC5MyK1cFW/bysvndBhy2k6lEKEo
KggfQsuFfPhaNJmO5a/2bAYHOGCyFm0XfrI14oYxlzBVTShMXsMQBdRZCdrZFLZ8
VVc75PB+de+kN/PNLwQJvpk9L/dFh5f3a8n7epxl7UP8eihWB7+tQcKzK/wkMDtQ
CLs339tcQNbLcEp2wgF/EO7wJBYucDmOz5LGPcxlw9rVN73o7U5lcsbfQWDgOVLU
I8sBbbQJxU1yekUg6moCsbrU8v+Qv6e8zhzZ2L5W3eH9fr3FKFNXvOWHKobd/5qO
8QraqXgg9HCO0SOBNTROPCJnFG65VvEKDojDzbqVAARa4nCEdq27yghd46iK8+jK
/d/SjDsUQwvO8YJY16FNrhAsvf7Y4PKbOTXYsvQrsoU/XLi6ctJifdsbaDtqomoc
kYR2lXueRUE4LDazBrKihM4LK4+O8MiTMAWB6Ub4yNgVO3Tth3Nc4o3bJoG2Tg3V
b20H11+ItRGp62Fc4XQYYEPTMls4VsSXc3vHg9G2g/D6cfyu2vS9hY7v7dra9ZuK
JzdXlDCAGP1gSMqLqS8iIQzwTgR+16scPDlREpq7QAk6BzAh7LHn6cbK9e8W2xpc
8m6caDSOfFCWRbbhbL+CN2vPWD0FAMogUZqheRAons1TD+14754ukLr3sjVOqq4I
TIvdHYrNWmex9FSHvqBf3uU2tP+8Q4i+3exnMNevJnl0KeEqhKC5xxVRYPSFFIaC
dYoh7H3qQioPGdmS//KE3WC2HArBGVXi2+7npvcB4XBp703eGi2WUznXGCgGt4y0
2n8rAnFi5hgv7u5HOSMx0768+tUPw03scOy68cywByjIl+MSijTI/G3XOuj9zr25
1AP2vtUb2b94fzP7d2u+csePLxnPkPfeADCY9RavUPt0TFibdz1wApb/1CIiSWQ4
aJTlYK0bK1NJujm5w/WG55yP45QXCXCbn8RMjwacwWCN8sAcBk4C1IXWw/p70Nk3
ZqT3L5pvH9LMUSJG2ePptRQfjtXx3K++hX3hFGgCA9GcJfvWVFaNzdYsX19p6WC1
JXI2nsXFoxtEjp3DIthZDVpB6uB6vmpXZwCA6obkDlEJ24h4RThroaChLW7roHBG
2PWesjiV3SGlBWUUxjKxiixEcQfe/ENR58qdiqG7jUJNlZ6qyYdDXpWpA7R0ZGYo
EudKn7ZYMJEQaa3vHSXBX3u7m0BNyWGSPpQ/8Ch59JrXqV2n3/TtrOJNh51OxuVs
MKs9xVZJDlIrXUxEW/35h2iCME+fop0YT6/N++5FMNBRPslmf7OrZLppUr/MdRgi
1VlxbhEaXOPbcgLyZA5pyOoDlU3AQygkJUHTuGiuaWdrLbZTivmbeQtpMKStD7Yu
2vQzQO8od0bQhPrBDxItYr2i2iQFBY+RIDJ9Gx0Lh/shB3XlLJMHL+12GH7IlhjL
UstnsbZxN5IaGPFLeW05yr0cJ6foNvGfZdEj8ngVB5TAjmhLwdWK95+Obem/segl
SmQY/hdP1DLmgpSSiCOhw9Hnz2PZJxFbK6WI6Dnbid9oqqVwjwzJ5Bjgp0cydLpV
jsOTdclQLA65Ogr1E7Q9l3r+/rwSs8VDWPwpmqr7ksJRvq3IDeNrxPy/bMAA5IJE
T6wTeXl5aF+kCOQOoMzMlpKdjANmmVYETesHb4SGlA4jBnTqSEAri8l4feZhkAbJ
QQ1myXNEud14tiSHxZCyght//mQ4vCPzLJ8ovK9vGtVcd5uREn6MkYwfR8+lcNEJ
zefDEJqXI4n/gTHtgxz8S9a2qI3XGiqd/BGhnZwqL9mkNzP9MNeQ4+KCOpJlqrNz
BtPEHO3M6ZjibiysDohaDmr3qwhkAQstCRxXDTpb+vQ=
`protect end_protected
