-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
jOufMMz2S/O8ueRD5psUgC5SnfcliOWXaDVy7gy0azPZBK9g2kRlFDVCOAfjSvLF
R/iTzgznSz2u3MzI2xSXW5A5UR762gyaOEOH98OoHqLxqq8h00JojXdzgkJUhj4b
2+VP2Jx3RpNjEnqLGZM1+X/ElJd3I4kxnj5CVcRlT+8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 36336)
`protect data_block
l3ZgHa5gmiKwyeGJPc+cJu6kfqZkQUVMBqAKdexhB/Bv62A2qN6iq+oJ0uq9/JEP
0fCSm/ZzNGfM890n8gNtGO/QCLBsuzY/EZqcEYDzIYnBWtrFWUYFItyydan8/VTS
oigsHj2/DmYPf2cA6qKS8BU+EbV/IbJakExatWyoQ1G5ZBmmbnYL2fMGiGa1wibr
4nUReciCs17L9vZ45AihSweVvJVm/RU4byj/fJ50Ugb0hOHclK3OZs8Gs13czpt+
GTPgic2EQC9HhFhHG50b7r0gKy+f7UuTag/MdhoVjaRMPg+l4xvbihUz7KllRzxe
K+hGVLmAzvY+gbGchLzENNKfPgyx7+j2gXZ+GPVTunCei7YEKdcZph42LgXrN+nP
SFrEem8JkaOhRMKGdJkgIUniEOuEJ2WlMRAiVizH4JI7rgVaqUqFwJYT48oYhiQX
WGWBUc0PWRszEoWNypws/8K46YEdng0omuuWwTToPcVxRj+9XtTLs3Vdv8McjvWH
mPwH8egwH9ADdaZ85jrpSd5Yg+IDoI9XkfyYmbElcxXBVVSsRKHkpuIATBi6QLqs
qLQM2lSo6XDzZ2NiEqBb4aCOsRxyyBzlpIio9wyVujwVguRaoGJIq8Cad+zWKnqw
YgcCdwWUGyLuv8wVL6Nd+7oUzvwGho+RPwHkbUPSVeEmEb/mvbCnv6dkg6Xwh6kA
8dq9Hnr7HlydqC0ASqhkjSzXDy3yF9q2+RIdRY1t5Gek766/xwZ6U5cxk7tp2qxH
ICecFX5QDcQKW1AOHjdJA/F6qt+hDWNFfwN7Zi3766f63ErrcXGciEXjTetGtZtm
ZgyNe9OxaPYyhMhbatU3vlTQ690w0Z6+AQ7lGv2Vwd81uxJdFJI+M3Tt8vLfLNkg
ylQkth45soHN/YR73RGSm9IfumvfCCr1HTgysZ2n31wug3MXSfegrjFGZ78h8ywP
CurtWKYkpYOdFvQgT9ZUQJlyAygfXhEHOr0H6su/KzDuhCEHamvigvPWdocazETY
qcxhtKXz9dud1uVAjCOc4Bb+35YY9fdsy7BtvuNlWC/BbEZaLzbf2MgRx76jgxc8
pbMnFSFN17U4yDZGNfXdEGTNTwQKAzDSxb6a1IVB02+tF9U1X4IaCowPRAnOyiMr
/bnCwW2j8CnyWoQ/UCfE1syfp4jdeCNOEgo9PvSDjHDXnkEmEXO0qfy/K7jHatdi
eb/k+0zCTjKkJgiMpWCMUTVvULB2o91X5SeDUKbf2dgFCxBSGQ3Aw6L+ksIQFPJz
GRaVXULDLWRpx1Rtb0Hah89EX9g30Au72ZckDIDvpqgEkdyXaNOMWN1uXh5UHqAB
Fpg7BhrhBN6h6Tw4HPRQw9YsQTa5V/GxxJAJHK0uYoy1Z/Cp71bo2Bup+RrC+McW
pWHUZNFytIOtBPbaHeVJTQpebCclwHJA4ByDZEoY0jDurFQWXCRthkcVKK0px53G
vWBwReIVxyTdB0gQ+5qPhdQqJkzrqkj1pb1fo+UZfNSWRtRelzFFibCDeUqZmWSh
AOjg9cg3EqU5r7aAbuktJX+ogxMchLATeuWViDvZglQhD0upc9QpNjxsMoG0JgeL
Z5t/npLMWH+5k0ac6D38QGGCO2X5rkbG4vf2RvAA2NlI5pXWRqzt3yEiBG8Dpg8n
1mFFXSK7MkT+yZe/UXZ1lTXmHDqGfGo78IUN666u0bkqbt0uvLVnn/1K2r1VW4QA
UpwjbkQzcbMOMrkhxsIQHyUB2UGAiPz85DhfKF72U6F+UfB5PTXfUjxIY71cpsHo
4OQEwCp1qBg9v5U7ZWloZjdlbHOBj64huezr40cLEVcNcbqP/2eIixJKjYjedKgQ
aEWcMM0dY47Ss6TpVFmf9QMPR+awuRk7fRNfVMdEJZs/chcoeNdtRe29WuEx/bTb
h7VrUcLctHdSjgY7g0H10iZJA2na9jFMrZGrz9bwnNlrgraz/3hNozx3HeEoKpbb
gJ48mj+7rIigW+dEzKCy4Zxwa3thMs/Ryom+YMcg80oKX6pXfvCk/exIKm9b9Xd7
VveuK1wRrkw8WaL7/TwtwI4WE1tW3wkynPwB+6tYIKSrUVqUaWdKtd7cyaR6JVP/
rY2wa8R6DtLKySDlutuOOkATtxp77Et1t8LmvyCZoVunzVCZfZCTVufFJ5SAvJQO
64AbUhkI1pWpAXakwOEMXia2aoup1A8po8NZLK0T3JDcJSZT4PpXqZeKio2sMC7/
HvHZ96BTQxAWfXeMh92hvsPPFOlce1DILgiyXPbiMkdLDIBEzVhrocY4JZAmAYNX
MWcSRqUx34VHBOgkmOwmCVh4fzLQS/XYN+2PZLuoYEyR8Fh322GBCbNDx7eTqiFw
A974AHRdeUO/LF+kyg3d55KGSwZcsHzggerqVvxvsBnuptp8u6Ug4aQ8s/xpEi5r
Bf9AMcE8GqR4hbA6TgLyw4zn3HszXo5TA3SzVq1Dvo/PDEIaWyCV2DB16YYhX9n4
R5qnLtYwixTBRC2xZjENpq8Z9/ZErQh1ILNZ8IE7v1QE/87dIZHGG+c8ApZ3QigD
eVl31NjRpCXwIkzZiw6GtomZMIo7RLigRR6uwbULOQrpQN/XmQxxNvuACS1xGu37
XZrDhuy+GuqzfBvIui9CyT7P3KlBbMi7kcQ4L7K+Ya+Bs3y00jF8X2OZ337dl4ML
mojrx1Zhc777nfx/RvP0Qlcac9p7Str5MlkvglkQVSaZdLpRYJYL8SPcl88pmZuE
NyN2jp/MbEc3wn/5WE+6VV77svA7xGHS6PipfK6iDD75sUqXxp5b6o2zGAjU7GP+
zdFYm7yo3zMVf+EJRUjVnz1knIgeRPobk/tGG4/Kj4pp4uQA6ry4AjovHKAffDCy
+qzBBouwXemLXkvdKVk3pjbhbD8mAn2c3VEzey6MSxp40usQY97ajo3q6ZiAmuOI
mHG2zfvSulP0MKm5TPGTLBydAEQoxFRRMx9BNrPtdM7vDylUuBgTnNFIHuJ5ibCt
/lj0PmuvEV2I1eCF9tQy6p1uqwhuSt+LvJv63ou4u+hmu+sp8yv+jOSnouQuqFxw
0Yf2mm2Af9BEtAOEkJit5wdHCh77+OwUQMkdLdiBth7t0aklTteQ4iW3JaAvj8En
H2S6ZXXZCUtjG+VvVNS0MFwcxPwHfa174l1fOYUk+vvinBWtUgZTjvHRrmC1/AOX
HDDx9kLm4s3f5S4kAmkqzwmpxW/1PZ0ryF/zIWQ6xcQ9uS/i2VV1tToo+k9l/BkH
1LBUmd/RDVZOZKVKYJIDu2wFl673Mf2P+SDVyyR4enBdmK+RsSp//bKQT1F5z4Qf
/oM+VPM6/4hYErgC+h4CWcltC7X8DcvX0JFqgCTX0PRytd943wCckzRN0QTNtbih
XlKfrCoUi3A/mm9TTo0PILhVpFAoXAOhWLb7jEUEMExB7ThAVrBakTfnE8YAxeOw
azyAUjWV2RiRPWDYV6fHS060PPS1RdhRB5Br9IqpKQw5i48ZaikJlcmExBVFWlkK
itfWAWen/JGq7re0Vz87opblTK7llR4pmfl60HB+Pm1g0tdFylyRVvHr29yNoftA
Usq0urnWt7ZBa+PoWrBWz239jFshfm76BIkaz7s7G8kbKd9n2I8wElqCoGkY5iV+
9nyIAl2kdrin348SmPb5/WGuHyNO3WhXTi/lGkbGKRU/HssAhH7vDdR7v9RjfvV0
CbDN0mpJZMzaM8+Ghig8Ka0zDoUH5PAxBHxABfGiPcV9HGCmDqYjAw4Kf2dd9h/M
Tfi7tv1UTTd5xU+nLX1TfYUM4ZLMx6UfBhWf1BqLFdqCejzbado6A5s4T9oKJV45
4jaofYuRM6aFt4LGQtfLKX5jhuaPKRoAGjvghXslCC9KvjGGcyML1G9RdWe+I0wZ
ngaG1b8frTrsVwksQwqNCeJ06fyIlvJVMrA3Z3nnskR0G3A9sBcrQs7I0+xX4aBX
XVFfDZnOym5wJXTbL3CXVy4sEndpWjlI2y33eYGrXiNp6H70/lWMY617st0YTKH3
QjH3qHvtxg044IzTXBo6y28hiz4HJDLiVAyM1w6GF4HnoH/lf/mMNdJ2Dnwoy/sq
u0jKimWVfwDvvtLY3C3fUe3UyEEIQgVWFF8hFlymWRylYa866q20HLbWFISD1ftm
uc2g589UKGM6LZZWNaIFqWY2/TEpgQSmgXheF8x+ClOj58ZG9/minbIXLKGFpKkx
7ewcujvQC963kx0+TO7f/KyhrqHAwQRj7wyFLvKd40VAtfTykc7LJqPBvqm251y6
JT0mdP7OoNNQK0zmXeXC6VwXEnaprmQctKgKP/dF9kIpalCMRD98y4Sx1OXrUxCu
+ogYmwuQbC7/PWJ7muAIsjttu1wheG1XZ3cLqn7t804oSmRF9d1ZIIOrKXwu9K2y
Nmgyg/jakbMsfrG1D+XlzVS3xzNWbl3MYC2bCKqWf3brOIteCipcKb17w72p0Sll
OMO+JF7UgIrPRX7MQ8kj/H75C02DR924GAzg1OfjupwfUhGtHKrlViFKdcS0oUiI
4Kh7I5Ivl8VsB7WmF6fkRQPN68vBAV9bjSNy/W1HfmRxTu9uiUbBCZ5KY1JBLFx8
jtiIW94uHM9UtCb2YYWVNfbYfzz4gEvqyesVKzc8Gb0Pe1ct1Q2tZKB3whZMwCzE
bNL1bY/CLXJ+gN3+4mIQXPMoTZzK6EGR1LU5fHAX/WRaxGotGVuQbKjjcYeW1c9q
OfuAojZCbH7ETf6YaltUvQ/VwaUOFrnjOS8K59rCbuvIamQCejAOgVaS1f38Nxwt
alrnxHD1iEyl6atfA/84Dd3y36EClMdx3OEVhl7YwwwWk1BXX5jwRoRgCWniB/h9
608u+48BAOOm5FwYO7CQ+0AcGyjq3moYTOUu7Y491s/RE5udtcICR2lgW6gL4dLl
qmqHkZN3/NsnjJJMJN2g9WM8C6aiGzOyT/TW5bS2Wf3cQEwo4nyU4/EEOem8oErQ
ajMrpUyey1A3RxqO+h92q8epVxoxqj6WHjkFLZOkzeUs3dMo3yJhclJ6ICIJkHMK
8gKVVog8QbQ2NSBmAfc+HvXrmu4iyidB0o5FTF4ZHGPGUOiN4svVQSKjX1iaKkR9
h4wzSqzIosd3pea9KKfAMyOsojgfhMl9WugnHvmH/3EQ5bC1btR91pKXMFMnFiTB
1Ff0qGtKHMCqDdo0OHlmKW5Kz2Dt7P75r5D/Vxk/X4uj/Eb/rw63+VVv2DQ6sl3F
QBg0FBltuU/ld7XuaDaI2PRI9mjBevw4o1iC+VBkYBN3YPeaQj5/HkjxAhuTkQ9Y
LVKDwwW1wLFtpRhJKxNE/TQas5xO8gv2Cd1vLnw8X+MAktOc1US2AMfDbFRL23Uc
XFdjNt4U3syzPMxXe2HkDPQi5+9j+QycAj/vvMcJSN9sU4olWPLj2QWSEzGZmzjF
P0O2DLfgAqd4SILJRfn0t4h45LJGK76TGDiCj7wR/T702hsG6erhwtboIpo0U87f
oWnZbvfVRy8ZSjVvV43J5M7zhzb0+CTn8LLZWX3pdHDILVFyTLaG3fkbrcyAmeaH
ghR62QCeXdUatTxkKfY1P+0N83+Nf8rQIXfN+ZN1L3l0VumCW13ywEN24dR/re1w
pUNgsPpfgSycKENXiEUh16Za7fJP4iA58eOtChTCh+DRiP8ezJFqyMUlyWtCKOYa
CnkNegOLJyds4WngD/IM3CeWtVdFdyzv9i3ym92EhziBjkC/Z2EKC7wuaqV76ChO
qtekWOU9gmws7L3O2NpH5HULTdff2tbxc7I88N+XyRD8gbkZbiiCEVeoZxoaDEIw
xLy/a+SXrK+cUx9PfV99ATqJjC+yC5aqJI6PIcCsy023zVmY7fpPLAQ9suzAoFuh
cUYXRAMI1s55rz9/pKfd3Ppp0dRiq8y1FZ2PdET+c/ewHbDpgZYMZyov+aSst4w1
i2h3Q3U8vAIMbnrJLyG53s8CePCfObqIwoqAa4nMREAMY490gbGHpiokw9th7L8a
2M/Ve47P3YinPYBAMJ3SnbXiFiM9KMXqsPre0Ocac3u1h9It7WRqvbPkie8RgNPc
4MGw4fUxJWV6IztA6je1tU7jiTd8mcLhZbmk8O+iZGyRCSzbyT18KNcvfvjIYSKR
cYbBxA3fPf3jbGlhj56YvffZw3xHn5o51AYyvXg5ORIIQNdDwPo6scxpjs+2UpG5
GMSh6QuGfCL+0JIEnTskHjyXnKf857KYbhfEB3n3M1T8MrNNZ0yNCEY2EitbikKu
DG5x5rTNAgE759olAhh7QNTKQwmm5SXqRJY70Sdfp3uvU6tPQZ54ig4avs3r4Lmb
VxgBw+GVV/kT2fNmzKpSWFL5nTgS82U0Zx4x1X/HttHojRM/EGBE+1pR8BOXpg1b
Ae0srmntKH0oKXyCsQzFwK5prjNHT5Cy0grbk9MjFb2zFAcD6pjEX3I33a7yK0Wm
cJPpmuCQNFGOWf1gF6YOGakFAmXmqT+SjYQyfjwuQjpO4qMBs8FugHUBxzU95Zk7
iwHcV+rjfPLIJ9K9I4QYko3BXQjHEIIggvQXVP1vcDBDywL96L/DJ2PVCtd5cRVW
CfLguqvW7BvvXGvbehJbMwdIx8D5s/X0MUHojoLRTmU6UmpgGOKLe4xiCzTcpvKg
ldZ/VzIa6/j8kDrs0zM2YMTelqL5IxoVmsEtLoHmq8KnGKqHq+c3Wi3CG8NQgUfI
MRwtpk6IvgY/DZDxSJox8zgWWt0zl7cfW2puYZIg54JnEEKp0lTfiOUk1Ja6rZEK
05IC1/d1KkyYwFQCS/Bd7RfElZy4rbr+t0TSnabTjsnp+Yk16D/Fgc5rCUScfBTw
iX8SPi5xmoxf1TyeWjzvinQfb7dAT4iKe0iqpm+pBOXx/oYnFZtlUFaXAgIgNUEv
IN7SqagvZ1w51tbPC0X/wC5r8IRTWg1FPf29vO9MQb5JVnU+PzU7YRgERgno26If
c/X0pubW4jXXRkCfY79DF+pGSpqRnOFaXsx7b9OFQRLuQe3CVoj5YHm+lXT6wynU
jxeHa0/QtOEZ+gfF4F7swLUmOn8KwlT/5AJaQCQbDcGZXuy2vd0f4j0OxJEonoZU
cANYP3wucvcb4Uqm/8RBTPEA8JEQuZiEhXA5dHL7GtnET4U63dKjF0rkvZ9dzZVT
FCnsw/bZoQYyGYgNocxaP4zwdUm5ENTD+p/shCjbdqydVRwSo/nVSmXwJTt+v2WP
DrBffH53T6s+VKsNt9tonTvTFoom0rrzReKkD7BU6jSpY7AcTNcaNYC/xzMEhQxj
JDkP/CuhcsFRvtEBJwNEMEAdBRDzZm0Cy3VVZT15tE1eNqXK0QAUv9Bhc0Fyr/xj
1UM7YC0j1Fnj/Zr+pDsSy2FBIPX4KNaMmOKABrQsddWMljg0goiqrLx9EnAZ8ha7
LuP+zmR242VS9jKe6Hi+n82txLhGsaySVZmbhgOARo8U0E5SHB5KtKki8KLfDOOJ
9oXEtef/xl/Xpry6rpe5n7fCLmdvt8JcTFAa7/SV40L9RY2uJq8CPTAio4AwzYRv
jScWkYLdnrTsyTKLVTCis0dI+jfX1md+803j6g2/xJPW8OOxiS/Vb5ygOYcPn7BR
e6jS2cWTH3ElP+bAB26Z6F2CXkMj2/O37kyh4RKbzJ6CP74GnWc6U0NB6yjxmEQa
oZ/cBsh//DVwtDt1UF1DEN5O3FPcBD0rhX8Eq+AzW+5/YUf0Odw08vUX2xoP/OPe
WMQ3ocsUYgy9V/VP89fnI/NOect8ySZcYBjS7T9yiL0p57TRX61cloitVNwVvfLF
ElFCbwa06NPy+c+pxaUuE78CZzW5sMhWionkwoeJH5dSDHpqcR5sV7PGWPH2OZFm
B1YtugAfsXNvXS4/8NLZ4qpykl04a1/UfJL/r6h9QIcUpUIV/5w7jWcjzUHvvVsM
AcC+aZpOGeJkdWHT0y+W2RMl2F3Oeh6q8z0afpQI7Z0sGv9hD4gkqUeNXCXUpDK6
WmeKV8ZvBqEIMB1aUU719SetwajCkOnvsduZwnObMiZ5jx2E68kBYPGrtklSyeHq
vB2LiBFjyHyTR8lJPfT/00FZ+N0itZ7orHUDVcNPgaPUw/pm4BYltqT2Bbd3G+Gl
+9K9Ewu84NA3E2SDbdH5Y61y0knRdhFOeIy0wvnJt2JPw9mBKvPu4jc+G+nYbOWy
gVurG4YSG13PZbvVkGEgW/co8K/bb0mN1E+Yu3fIK2+3vghvmW1mgkSIV5K4WSES
DVn87LpfQXiwtBaDZPdpjC00jFvoRfNNi/F0eW9yYw9d8Ut8ALNc/nhzeWCarazb
BSvJWaZrKAwKavNjtyZ+wDTr5e1l+k0pYugGrRn9+SdF/ROJ68gOmklwwTtJ2RV+
CI37qVyGK3cKEs3+3kh14/hgo/QGJR0/qR7PBrwtr3GYvgWFhWhqmpTsc9IawTru
/+WcMPPiBotGR+Pq1xoBUQVTBstwqLqm7BdNe92HMfyH3Qa/lZ2JpTw/YNdUugRY
fz48MwZBr8c4Et1SyGIvOqOYYveRHh6b15r5jp3ZiR1dwdE3KQdIPYSt6XPl+NOP
qnkvEL44orHZ5nxQs7B9p3vP6Rq/7EJYi1jqqTxFZEoc7XKNlraOV2TxGQwsPR5R
7UDsLsSXMULmk+yNBCVoEKvcms4RE8oZNYDisGp6ORpMov6IJy9Tg0D+gUC1giKq
CB6xnBnZXy56HGpH135uN0TemH9T7nXNTWOtrhm4EdiX7vklzKqqEfdstuWVCEHA
dwbAOaSIBbAKkTnSeeD87KXeXNuHs5ANEdwzis1R7zbtPFr4gaF144+q728YOlQ7
XjWzzFFKOVCm+R7XbGj23xCr2XGxVQ8bWZRaKAPGxtmYnTjTXyy2mRhZdXaP5fCd
sx5hPwFrIcILvSGHwQihjsJBJX0Fq1/9jPopO4x8i5HhID8cgaNdUxSr6zImZLES
lXUROirCFPsdqVW5BA4XONbZW0mQRwgEkwXW2HroHcf9VKYgl8Z3qe2HNbWEd4T/
rnbASdli94mXFoqscgxHjvL+oeqAVG2ZVEpurohTeevn8SEjGVGr4e61PzyMUHTm
HtJA5jHjlOzmcWQZSVEjJv2+r1mBiJBGaodKDinteH20xWJSUiPJp+YP1Rrsoudl
maEJw9azF60wXsvdNTHWlYhT4PYetyX1Pvfe2JI0FRK2v54pGRT2wDJoBP+nLVRF
o6ZPOn1wVLxQ55vVOrgiivqCsggMbWWlC6qHtsDnfrR0o5tB4jp9fnRIyOlcP1Rq
UdVCKIYusflZ18i650qj6wPzaOlXnF7m+IaR9IzVgufWFT7EAJgIxzz15ZGzm7lX
NVVgVi3GYHMBbzoumsRl4ViKOWJO382Hk2gFPUHLQaj5e8K8ySbg8iZhGUYnVi6H
ao/N2p0Lxnjnuod2T5hqjbGt47d6E+Vq9r+eV5PsO4TIJnWB03Ey+9xnOlQdYAf/
Teaw28e46L7xcSCORScyF8QoMuGDV2nVz7y5zybibho2rFmjkcD2beCym9k1m9i3
Dnj1+DvLiY2rVKPSb9Zx/SkCqFDyCuc2pQWC1GSIUL+1M/mm1kkEtsJn4FrXmdY/
W6SshMc5DtSqKmB4xOl2a9BuzKjSFSnmHOssMtdifZgt0qOawDJVGYVoY7gI76IP
p99kQi1+izSVTJqZG7Cj9K2i5we3o3zGXtDaGPb9Ucc9o/b/4OWqyrFz4ZGzzSOB
9MiQePkZjzLHbl8V0EikkCEG05nfu5x6rFdXihknZhktLB+QBKXi5AbmTv+/VaW3
rmCaalDMlCl4MAkvomvyycNVLEjungj9ZR3GqgQ8KPdZ3inGRgroY5YVqLvuqTVj
kVA0XjeJk/Rj3wuvQt3yM8ZGEkVO6/Stov59w7ej8LMCTf0QqZETQbEnyglbbrEO
Q/ls6CIQxqv+v636Go6B90mMQ3/faCQY8SGGYemyms2nhhI2akOYBk5js/TZn4F9
mdyaQ3A8hCJVJwGKn0z9eK/eGYeFDfKeeDwGm9pd2y1SPP8E6mloL8/NxEFZ3VWy
8yOhTbDeu1Go3h2/5KvNIWs7Xv/IUzunnflVYoE4wSI7JabZR8B5XIF3hkar7tmP
UD8a6vN7Wf8qSnUPcnojSgcaTw+LMkV/5eiy/H2iCMbAH+dulUN/nrqYRa4CADVB
cTj2XcP34cyVldp5DK7WD4obigX4MAhSxi4XbOIeq/VL5KYo/SH9QmBZXGmmwp86
cK4FVwsYrCSF8859nwqFCvMMBVDLkTs22yV/AcKsSJg+LkOULkaxnd/yoH/gkZUK
yfNbB/HGljHqYJfSxpbU6nwAqlIaStyLCSohUldaQo8fxAAuq4dfgnOhUSGBYnLj
TnSZjUeWV+sDG2EpAgmGqkOxcgaBFZbmD5GRn7Mj7hyk0JFApV/GfrmXtL3+b5d6
UcrLuSJjI6BYXX6p8LF1WV6zQUWUhryRCwfgU2KTwbKvZiuiZHkDaJRwxJm7vfso
UdjJYqoIxYOOoq0K3Fo4X7+LI+Dh9JgRsgFbSm8sOdunIt2tCtZsri/dzUVl1Ufe
gjVJ31mgJXKBijk1+nh8otEpf3wBA5nidjOVJnVCVbsacCJH7vn3RIb/BU8eVpmy
MGZAUPpoaxUN4vKVubjabgvfBSBiSaBsv+0OJL5Nj/Zs6EsP/YbeiplT06HuklOU
zc71M3R8TuERNYOGx/YLAA9clveQT4sGeTxPyBB2uae+7whIOFyAzXnU/6w/6nLV
Ej/eNwN4gtRvV1mVmi0dFE/c7UuYzYpKXnepVeNIC5GbwfRBbiEWulbJpXfQp51Q
IjPtGuJqg5JUsZeusUTjgoe6rRqDMGDmaOC6jWd05L0bFR1MlGSirN/ldbY425jd
SCFIcvjgzu9VxQTZrjGZL/QwW50eWuxlgg6g1WmT6HCqrLnsxDZ3fnD9dPloOp8l
LcNnjovVN+6T9Tw96n/8Dvs9ULNI2DzzHPZc0OJphP7Q9Q0KphE8aqh8M3FMMvmq
g0l2TmLKTl35ez6Q6HR/6hc3MKG0xTR/7dEHZPLERVe0kRr7JzfDoWwkTf0ohl+g
SvA0gaOk2m5vUYWdK4luCX81UF2vvO1HOUzbgUzrSTAfKxao8nuWlarYU4YpxBPg
i0b2jFYzf/fYYhmneIb2vFbLQYACTf6o7Pqa/WKph1q+4nUTM22fHSgnaB/d735s
xcSJi9jKlSycKHRrmvQRBMUlpQ4aM+fCsIRYmJ4nMYLCQOmBbahuVBHD/aMH+DNZ
v8ZI1l0CgQurgYU8QjnLGbTY4zFuFW10F15/B8B963Ti84rZO1MtQuQmwENsbfwe
ZWX3qinmnG1o6hgFEevdVeqXprHIufC7ODhO5mX160JMzfLxn9auor64WKG/8kRR
zsvWKMhLr2gPHhp6NkCich0ylTh8A6EHEf98z+RCH0USPhOjAB6stZpROyZvBt6V
gg2gcnzZAVVM84Nco5R9+3Tcvyfk9Hx62eEdECieRN2zKkykYPERLJTvV/gXLa8C
/YutrhMpnf5q47rNlOZ8TW8O3YRP7pGJ8hW1C6TjdmaHWuM6epqXbxj6CKIecol4
36ipMnQw+J/8cDEJH51zyh5gRgokGYofRnzG23G3F9KaC0yyTMIH6JgoNwM6DynE
KgdzDBFO8b4NSNDXsEPc+sVTqGUo0xqvKOLzyDOlgW+U0OtwaB3/CvFWkloOnZHB
4ShwCgxIExYsp59Jv24kF3RKwp7+9V0ducGSraNJ18iMOX+5ySdCVWdJ2BwilH0A
X/gSemUj85d2lG0u1wOvAzwY0NerApzd7iiysPTra+RQft0038uj9J+56qIfrj1L
Efm5rqowVFlG1fcjr3CB5phT7CsDQvB5lhbMdpBAKKHvK+RnGAWtJCGII4oSEB+F
6uZqS4BN2Pu2H9fHx9L2kZRYedizTde/OpR4LyhmCFcZEIGRbL6SI5hjeWolWCxQ
gZ/fB8GZhUjQLm2XzINaT1O5RYMVwqAWJCI++4p+Y5hHbK1umCFYXxSDgSgBULJV
+Pk5VN7JuTsCrGY2YGMPo/gcCBcW4TTsirX4UPzJHAtAwpV1u7GGv4wUH0Pj/euu
aUZwfR96scQyn4u+yPKpIQ0wDKpMq0yZ/nYFBURJ3zIVFDzb9PAYgAoNB7pb3BN/
tTTWaCiVVTaJuOVP6RsJLoKEosHaKUaKov6sFJNXWSHV8NqF9qtzQNsxVqOLxxEf
fedfkI+7HGlJbo6yDW2SFhyb19xYj/l+UjNcAwDC9rG/cQ1tz7zjzb1clGLa8p0G
dI9BfRKf4iRqVvqQQRB7YxP9BcJQ3tCP3ADYWcPSKmTwI9GG/6WifAm3SUy198XY
GOoOjtsCGBQOUVLdJy5ehSs8iCVQ7WBe6um6HTBTGB6UWvusoFyf2xPg+HkvK+FH
3uI+V/CbA0fyoFi3kWU3r6tVSNFDQOvMfETq23W3xSSOqKKrpdIde2y1ysm9WTaX
CORUgTEc3jSSnbI6EpUHO2k7mCDOATXbbRJHXDUhgsy9ZxgayyZU4g4rutllLN8s
mQGwKZ+/ABPWfp37slQ8AKPUoCfsVNh8ytBuoQ+xhdtg4E6vy1T4mEkPtoeF6B8g
aarhWGxDC7bhpJLomAYqLwAHAE6Teyykidv11MKG9w20GHNQ9YvEzSu/07qr2wse
GfZFk9in/aXS3km6OfuC6GsAFkwv48ok5J8GH64RzSgpyUeWcM/3l5iso+rXVKed
N/VLz6N+GUXbtO2Hv3mEnZSTBx4kd5wDVq/2Kvd9l/skAZeMR3LHlMu9A+cVH5N2
FRNRcvLzqA3tiW065+Yaoa1zMLPvJX1GyPTB2ttvM+PSQjUgtcbG326CrGh7bBRq
3Lw46p9YGVr7DMTbQbmDmIpmTeFGNY9FBNBEt+ZGhr1iVcv0r5Bg3vhZAqZoDi/e
mkPIt5uZ6i15XzvtrHgpmG26OWIveYe1yzAQFGd3gs8O+k2fIUvnAn6F4gJBcwSJ
Jw4vf5tW1JdLhbVIJuLsqQ/jkoqGYyOIDgC9ja7CKoNqNVil8ZeT01UvAYdfiGf3
tTN/BGmUVWgAs7fiLoUWSv9ubAPvT6txF1G0UlpO/aAnFSRNZn1QLLYW/uMe9qyw
kfxzaUR5X+8So4Gk3Bu3AFCFuM9xkbqpFMJVisgk5EWacs+OQn0n9rlhrNjq5hf9
WbwQivylKkpaNTyTe5eVyMoYo4wqezDke2le2MEnGnQK2zuDjBRl4GvFv1ukmp9r
JxuGQijEOt4l4Dg0NGAZyzVmwvLMgd07QNPdv3gnIbz8ina5X4cdy+mK8rr+8qK9
1VQpvDMiLuqJVMgSDClh4PgwB/HQ4nXSTpBCTG9zGcGEkzhNvCidAjI6Thx0+82w
NFkLVw8RoexxGetVGHPT9SYAz2A0xoTUTQxQVpwtdSnH4obUnrHRJkFRPRfo3q+u
j6lJrM/itpMj8PCAiw+mLX0sXh1DxGL5rztBpSonsBhEvlSwtHT58qZ+kTaHQ6/U
IbpnlyXyrNTPGcw3LEi01aQEe/800fmLohn2Ibe4p6Y4c4xqCmkPSTBkPGh4FV2u
KqLd6dOks+3RIrgE7HMxgwNga/6t34jM5dy9m18IwuoxxOLeg8ioEYJUOawDVZax
yU2FjYZ0UAqDtJmXbJwWwPs0g3bYLx53NebqDlKGkMnJwxEOCamX2af8VpjXb/6Y
lEB5NbgZxhKfo86t4FfYJ1vexNDc5Z+1xTqeG8eaRhzKSdGnsLXD+tzLuTOdJuu8
vhSBFJ4oBsFganpo/ux6Nem/ttwNlI7L9We2u+1wqb3DCp0XWKXU34TWbM5CTGKv
Vo0LxLFpMHnH/XWBhF9cd/96c29ORbo6XXBRl8wRtCAEROliWMQ3UuXIHFIupHIM
lx/HzV9A6nJtgfeqRlduhouZa1NKnYdMM0bhORpMqMOLt9v0TpEIdunud+9xRJTu
YatsACm8ZewHfWcVjZDsA24J1ZM9T8/5sh/t4B3ZNlJFsBFAltZOIb2Hvavrd7zB
bSIbIjjVhi40sXtwP/TuV240wv1W5Slfqlaf8KijISoaicLbJiWSDP9TcZd+YNhy
kDZQDybSDSE8/JcTNHRcIcTJ8ea33hBAJR/bsTZFDIKHanYyQOlbz2kX5Pw7asTp
reZ1TC3DXDibbanjJc6Agf+FD0N7Td3cizekQeql96az/HNifBfGYhaX9KxcaEDB
Xg+pg5gG7iBXrTYY0gr171YCvS9Qr00i66T72WrMlHhye+mVFR33uQ+DXuOtaQuC
OogdVlh3xjLjPUPvH5gqItQR8EWf/XiAiV1dWS2GAx2PDYZ11oOw7zaFJUjsblLm
4oTcL/Bz8Lkwv/11+S/05J6DU6mxUbuEtO+SofrQw3NPBRoeILjUhBQi7lL5BuLC
nDyuyq+jClrko8nZL6h1q7aQ6wS5AxoZe46shQt4bm3dDcRebQ+E1JFDA7UZk6W0
uOj8LecFyXSIxawk88FA3FoX7bkss9kCXdSLrFw+IkjpmhPjNvbLZB+NUwBpgIba
KC1KoXU2rcYYEYiz7CRIgNSSBw3aDq3q1+x1IC2bi53v0w7Bc3RFty4NzjlOsLUy
KGV+PDU9pQdPf/zYIubwrzaeKWfxqjUS1iaYODGwe7JbjWu7I0dWIjto/eAHoAo7
it5ElapyZLiOEROP266F6pTkjT0+5wW9nNHTED21tIY2njCimMdmO5AFyG1M8RL9
Kq/kQMv50XV+ruRRn+pi+D2GcDUNO7nsxA76fcG8Avlg4IWy22tQ6zH3BdCB/7q3
tqtrXFPIg0aGheeHdD9pNpzcoeczY+BEEydQ+dBUxOhcZoQTIvzRGtjmj64DG2+k
B2lm9YysBodIcHawA0z/4f1YCy5HJ70OQHHvuBY9u02rKFFNgxFGR3Ki8fie5ot2
2Wr9cGr9eiHXZMFthd4o8sgRQeniJVrFzQznNhFsjs815S4sobFtu6Ef9RLZfnHu
mGSdLqUYj9zAHjbUrUVHWiL7PR1YAw1LYkFlQIsWJMEzqjuEoP3QVsKhkiGquBBX
ftm3RYCFXh9T8KLInsh4MDwJZudFZqAXj2IPFNGomaAGwL4fK6LR7Wd5B7fCeLKL
sOyrmMa8FuNn1HK0JgFvkSNi/k9tUiG9/W/Py5GH3kdyNggVYkakJ7BIiJYyMb4c
1wLGSV9TfsQ1080mp++p+xVLA/kexxFJ1d77GyX8dxZe2CD/uWm+dSHcjfMG1+ad
fWdSCbH8ouqWYsEFpfbqR/XuRbbgYOaHSeFIvKHzawPTVu0VfTMjxn7Urn0J7OYG
QhFGrSk8/Ae0wHW5J6SZ4iB2PhGZ+arkFM/ssDOidCKQmvfm/5+jTcan3UP+R/4C
OI54tO1Ce0LBRAqNBX29HL6Jcz+nEnBFhSDryHjNu2X2Vr04P0x4Rv0vh3tUXBMy
f9AABPSzmENVuCsVvvCsjZOdnA0k/Rf42JGL75EU6sWR8H8E+rgq4R+MwPZNnni6
aO3quedSAb6yQbLyNlmu2uzCiKsrp6fhIxclL1Z1wXNVdQWoy7X3NIkbNh/LflfX
ho/GjLiezGJL9kIzVnLCE5dST/o4fa/3QJSFG6I/9DZCNvMMWLl2cbW255yEoj+U
n55drHiOlHup++/ji3B8FoH9cGFdg21iFSTRPAAKxgXysmDaEDi2d9s5ML8lmLKg
KUHZhJF1ImI1u++V6r/trbEorFy4n/NgnYQ4ToLzremCAWUyF8Hax8jUu1i2j9iN
56kDIigF79O+MO/+Y2yI78aaM7rHkXpFdsAXAGY+zRpkqfSiKLD1hMVrcdwb1K0M
t5aWMo1xN4wwl4jAs57mh+SNIOuXkO1X+u5wMUnx/qF4VcPfSI4dbKzA/erL/M+F
inQJomGycKnbAuR1aJ7NvmZs8l0aPWJj5227cctg6t4cKwNLOeVU+vyGQR7RTwou
CmRy6LD4Wu2wR6P8TsNAYzWj18ac2W2Hc1D4uVgD9kcbhXZ7uvucn22TO9Hd4kFm
XUNUP7mMLBBSrpyvUDwdg7de3V24IKOVGDLFHqGCUEgIW9m2ImMSZ5ciuVvFOWCZ
JT6+n0ALIsmPDJEhWMIvZ2JM/g+YpmKs2eR6rvd8eddzu3eU1sKDvD5AgWkpuSMO
R4LCb7J4RK9JAZDphwpsixTINI+asYYBUjVQZwdxtNYQrpwkxblLVhfrlb1V4sHu
4ZozsSaoLjFV/IkroKsXRWurlTvRGgSNW5bInYnM0ot4yE3b275J1RouBybYkukX
7XgwiI0EpNo1uJB8+HNZzTH8FCbPEJn4DuJYwrbvuOOJC776+f/UJXPXGhuGrb+Y
xePtesEWwznJ5VyWYsw8O6folTpXtzLP4YQsLyiAyHtknzRYrvvERadWvHqalcMj
IQjUTPeASfuOJDe+tor+FsMwhtc2RvMweTU6qfDqkigOVDUBvMXPmpVOz5yLyfV7
70eabfJbd1asXjtevZEGw/LVMRTj37gF33HTihuvigc9p0ylKZ59DAfT9cw0r+08
R+ab04PBiEejNQLcB1oCCYa0ZORi9yMOHs4bnR7aaQyvfvUlsdLbJ4YevluKUW3P
1KCrScz3lzQdtZrZJCu6pJ44tfiftT3LJPmyj2JHzFgGCVlaBb56nxJHmoYVpnsZ
IJ3NQ0RUEY0w4kg+BzAKYuC8Oh5RtUgDuT/aPVP2ykh27ctSrhYUB54ayfY8irDv
AX25upqlxproNeqp/QRGVjyhGDVBLmAldpjkFAZMc6LYkxU9qZqgo1+I+eRTrRnb
Nch0TjhMw8bMcNgJUUCq9t8KcjmcoDA+GwEy3fHfO1JtEFoRooGikJEZH1C/hlFT
MRLrG4akeq/enCFcZ8tiZnc/bDFXDeFv6S+ziKXT6dfGfgAHpzk+35t6Yf8VcXDh
bfvIsvm0f02HQUerI+yLXX6qGXIMG3pLbPqnUEck0wEQdYiutoS3muMrTTWobRtH
Sc85d/vbwdTX/jgXsK8/+D8rM6MIafurTi4g5UXBfHvnFGyX/QRYMDjtDtneKFpp
yafswaFKsjxJ6s0AHPGBsvtKqOqBkvf6PqIobUSf/mlyUTmFnMuVQneWzDE1G8C5
k3Y7cjtCgRzm2/UZigezcNL4oUH3wq0/1nwiOKC/BDyxV2BCG/KHsykFYDj1Jujt
M9ej2go323BSKB4XJNyuqMyovoGd+a1Pma2vRsaS3+Yb07VwZ4cESHc/6AaOy0s6
cIrGsIGaVdwiIy6VjOmomTeqqMGvs+qNZcaNFSTvMLGfZG994tCul4H41HLKf0GS
kxzi1c2gHCUlOekJeKoOqyDSFS2D+emoa8TWNlqDuc3Z0b5s4yIIIGhXT2k8dzbl
j3H+DMIWKTzvUYD790oltIfRJtEQ3jZV8Lf4KPa+818UPwvdjJKxQQ4b/LRQHSc/
CxOJjOYRWcIBq0kG5ckJubqih9UtJwC+v3V3VeFQlTf47Byy0H+u1OuPeBiYfQku
q4DEQ/CZeCPlHZjSxalXpxz292Abae36uBFbCTTXFGAENirbcE4B8ZQ2ZLJqMsfk
o3JNLSufydYU2OiR4yAD/XM5oTFMJNxHQUQeM7UwhTHIj1afga+STUWcKde0xyvl
PP6lh75vuDjEddXcTYeGyQvebAwdDGvqQQ9oo8pswW1nJuoY/x3kb2VCoQQjtok5
mJmpHcLRyvmYSj0D4gzoL82MgCN/vmWBMJUNk+ksHivetqOzc0Z17BQN0n+EjxZp
rO4lCw5Txy+q4thBYheN9T5XBHv2vvU8HXLmc9SFpI4bg51a/lhNLIP844inB0jQ
8HDrJqIU8NfVQ2BpciMuuNCwptKD+srtbWJwbW8o+H04rg4qqB/94yCwDXx718nm
u0PyQFq4MuOB/ldgnkueOgw6oQWSenmPcM/xBhOHmDCMOgHuf74h1yCU4uLdJvqf
HuBwMK9089t0J4QNmvQTaLtB9/Le5196vP1pDB6649Gy0AzSTqTrsI//M/MJrCEw
Z+8Vg65a28pXxIIZhsB60slO7Z5noVrmtx344S83ttl38kWk9qMzIuX/rLvLPzW7
z7aA2w+qVMySTpiDn6+flTZMAVMTmDpzzX4YOgA4GjCTm7GAQmb14K2vnXPS+Tvz
X4NjhQqbQxw5zl8eCkSgyC4NKmV1Vt5cXt6IUC5g9vGJ+56ENltdlKDiKL1j1yko
ZdQEl+Wl5XuufhLJfTn2qPFvz76x0A+eSmrHgDlOQConHyJa7wkffYPCexIhCFmU
+Kg4kva95EOJ2fydXxnFHlQ4A0WlFi/krEvQ6R8Tn3co4S5Az0fjqVLHEdmcTl7r
DBofJZ6dNGPY/cDQfH0WXELFMLG/aB0FA9QiIz05o4cmCJV4E+DAbUa6nGdpGNKl
B1ZYK54SH3hJCIFk6tPYRms0/h8FnJZv4z5rMG6OU5kWF/bpapKem2+bZvKgolyj
xw6eAJLap4nZ2xuat6gQjLZo4lZf32Vmt4HG9H0DMAdLtcEN3NDGiYnlk8LCups+
k5PSmQiMToldzrwfcXTfpqFJRHZW3mFXbyP3/7tvsPaCLbGCMsxsebjX2JFG+cJX
INznVTbDbnV652MdTz2QI2ZFEfhK+ex21hcWyZxs9TG7LO19G/3T3FJtPecl04bV
Tj+rks/XdQnZoOWe5QtF9A6DRUY1CF7Q7b3shnCaavFIYO1ZzFNs9+gAPmT2LY1z
vTzVhxfIiMJX1wWebaY1teDB+IwNnq1TLa6RXAJ3A6izjw5/v+VXuDvPrAGHKE5d
1en8fsmUPPPqXMQXfMMBsFBp+Xzol7HCkmZOX16nwXRum81ZYzERPspaxa3yzojq
cobzgAlc/vemOjVFk9QMjMXZG+a4zzU95UeuELATAkoPw9bGRPh73k5LoPz2v8HX
evWB2a1bMPCgF1bwhGu9rlZpGNEYpfNDDopZFpNpxNib5jUcSMv90JaL3JXTqSke
QJqi/HTdq5JEie5d8XOoNvENldM48QSlymh1pztJ9A+ClmbWGSMZnWUwcoGoLBN5
ABDteBi835PibBuuYbBxvgspIp2M9nRrmEcLS32FZLKHYMkU0pyab3FL4IosTLIN
GmSPG+lOx+ONO9g33M2FsDOZRoJdV6dMmbEdnsT6pTF0KxMFe3Fa+OfgebnUKQVv
vcQeDVt8GIsutwTji3kP3STmi4SYJURoXxtTHqWnZTyiaHCd4TYbijWkY1rB4OJI
QBbIZy8aMdexe5UP+uNdqNo3qwLQyKFtafjXZFp4WIkQxRZFweMZj/05m36eePd8
d0cJWBSA8p2DSProOg16OTqUjsHsQzJurlYoEDmUBTjdFU+8vZsZY19VGxvmu5co
NFq0QD1sLvj28ltHhu5grzRS8uRYwVR5Ox78C/PcwvWP01rfDr5F8OoKtpc+DIl4
IkOdlVm4YDhLwjKC83qx1LXO8DF/fCKot56rtq1x4yNXsiCyZyndXv+OdcLZrrTI
4y1IlsvABRhUnS6c4v63xSUPOx1H8tdhyE8hWXnMvSYHiZdYsIZDV/5arSmNgy8R
KtcpJnQRw0M0Dg2eDcJKzdcfQbF3BPdGaQ/141Jw7Xe2n9nWcVUCg28orMCo8dp1
oPW9KirhjjQrhStQ3W1xoVGq7k7CySfoOj+4OjzFeExQfTxcLeR7yhJ9YI/w2wAI
eoXgtwQE4OVcP49/sZ5uX4BmAWx5UlSWZjjCjr2hcRmjjlLQS07ZZahvF70i9bNK
3m2rx9gY3lJJ8+zm4MMq+3uQY2TzbW51KgLdWPsWNzhmdwjpMBbyutkXaNKJsdwj
xBP5BkuhER08bsSMOy6rg+s/d/I8BNlzdzQBZmbElbXchDlXv2OctiJsfSVb6e4e
loSmq4D8T7QsBTUhbSUY4TU5p9dzRVIOoY/X0bYeStTPAwp2eVXmY4LuBqIOXJfE
h8IsOEJXwgLtcj8IjsISai2DUtXhbIrnnzdIflbQbgmpMlA1G7uOdQPwXrnVjsBf
8FnazMZDRm3YRMKh+aiVFHlPtA8qGGQ49QgMX2N9X5l6b6NHu28vsjlLgHi7Mzko
hodtD7dwxUdTxGXU0pa8BtkRJFR3kEzMONCntJZghuHVdSyqQnh9/l2j753WhQqE
GqMhGLE9u7qR2TnDz2ibmBYb+citCOtNqMrOgNZ/A+S+os9jpEcHxoKs/qMRMs+Y
HAbpW7/yj/smSpyp5UxXT9rvO5ZqEuBGgPcOEqRGzajpRk8L1+w9iT39BGUZF87m
rFBBwg4frOQ2+/UHEknOfq0jQK1VrGAVYJ+Iqps8gkUIE8cU+fS7yL2G/7ec1gTl
ewxg5+btipv3kzRJXypU+DZXCLvYDtJ/y2IvBnwyIyYBpT8gQ6YDxApzc7vK/wE4
qnS3hUmdt+ccYZHgECZWA2LNiTbD5whGUTkUO+9teX8+m5v/6KRZl4DakHYdZOLq
pImk2A3quiA9WJyoSkiER1Ks8JtCkPXrDVzFUxv7W/53FIgGYQ6eltuBb4J3DXmy
aLI//sfyerkekq31kbH1Av9p8Q/sG/lroiIvpwk3BeRLbXGMtRia6C59TurjosOt
cLWUksUHjSFKoZ67jEQVmLk1jQdsYOA+zx+LdfY5a8yK2DEc/o4OGrP9y1b6ajNa
jUwp7HyWQA0BgMAWWhcXtl999Jed+WUoRvUxdiW/mcNCq+EwliaD4kAAOadT/G5y
JhTnMdsdxFoW2nz/H82sHXG+Q9GEt0QyXkvoMJBj8N+KRfPVnbbcbV+tIDAJoLfH
1PQEFXFzp2jwjGTQvz+9C8NfYuMk5P8qUiAB8ctFaXa/CmoA1AfmJ9x6vjR6Ntsc
0suuDpdwMH3FLdiSR7kNE4qATQjcO2iC74gCY90fj7vj+VQ48oqxHt/rNvKYyzuz
PdVW4DOJyiUrs72HbQdIe/f2XUpryfzHxa8b3OZvFbsBcpdRu7c+J+FmhpW9l6o0
qQcFb5Y5trK9erzwxpNRAFyMvhcLs8rTOLa/BfSqtl8fF0zhsCdZ04Y4iOhDZoch
5EQZaEnU1dFGfNqiFYJocT5BbKW8Sg93bJdIdkZmCjU5dzn/j9TlfAot7Lp02WoX
SjluZvjkdOrMPjPiHKgU4H1vf9JwF+Ikw+XZxon9t0svG9MNvdp9LDRz9t0BsgQx
HZRsgfAHaQ6GdvUTTg3Sne0XDnJrfyqrXYMY31aW8PA9XokqFxWAOsxwZRADeYg2
dXXO3y1xCy0MpVaH2vXMEF7EE1FS/2Z4FlJOAMNoMBKh6zYrhkc0ihnBYyIYQq5t
jeGVkAVgXdw5L+D4vsCWjdxa5Yvrw7dDk2sZShomVVuMT+kRcBdJ40hQXzB9brDO
Dp1nfMiQdou0lrcIu3FR7u1mGbM/FuPMHpepxVNj07VkQGdVodZGy3E9CN9/TNVk
xphy5E8BAxaB6ltIOeI7h3linVteTe+1Xko/eEtHjgcVa6OdoIgMyFRQeHeqZMX8
TlBuDCPfOI7opfrM59qYClgiwiUC2xiRxD7u/8evZoHJIT4F9sm9bO3Wx9i7pscc
nVnq5ZKgPTIcFQPLvPbXXmsuvnmx+DICLWWnn8ME7Z4037OjAVwuzzMQW2U9GtLI
MkUvSh8KsRrn3UxB1HSrfjFkIwdWpyzFynt0J94tOeQxIYkvDJ35UmyNNbjndXjw
/0rhWYNw7Ms5ULWbGUD7/5RV9SpDqV4A34VjWHoctfo2aG39qGCWL0mrmWtyctq1
bdrU+MqHdZLo/nJbRaU3woR94vKYrzcYAgOtZR8coTSDfAVFMsb8DwhbeZhMnyXo
WRgib32GtgeYXyR7CwXsNH2ti6jTYzjp81i1QU9rZVrvBVxo5ZWJAg+rjo5rvpBL
4eHs41c1rd30aczRAaXpnllabdSaHk/NwLQnL5Zg7kdoc6/pzd6F3B2ZywFIdMVx
0EICuOZcbVxI3ooqxK4EBYO/Q6Q2K1d+T8BOF46D7wP3iKdqwfz0fWNkqZF4utRk
gkrAcd47yYmKBfQlCZ/wlcLPlSKEajQvc3IV76YUJsXG8v6YibhnB7sJpAnxbXVx
mDLQ02mH0e+zz2q7OCfZ9xC5UmmdSFEUAnKuAxlkXv+WrlsAxXo0LH9DMBHXGhEv
29KkhJwJPf/XwmaHkKgJpuwfbznr3WirVXVayrv8sEQtT9061++ZPTvRlKScc7UK
J1l5jWf/K8NNClAh1p6tGAioLdeGRZ02YCu3Iy8G5hSLrUERUNc0aXsSI/5Xugac
lYSnFCcQNz74rDqab+pne56XO++aTUjJBdLVhD6VmWI6I+MTvXsLyyE4euy6T5rG
Aacb/aOLb7B8ZQ1cbR33fBXX+9zB/Nk8Vipx29GGMQER77jJfHjHUSInBt82bIcQ
0yHmNSr7Il79mJPdqxHiRBUFG26NcEtoT0cKdLBfpKK81B4Whp+q/Mb/LKTZYDPr
z0dz2VOPd6PM9TQ/TusX0OrpancfpBeUcnqoMnnkEBazdsiTXJvmJ8AJQOWgVHpN
AvrfWOEn9SKd0TGMVZfker98uEGpTtR2dL0KL7HDtNsr7QfW+au8YLMTsTTSWgdT
dlwwop8YLvGEU/YVSquvam3O4ieajNr5CYIksoaoKQ7NF+TU9eni/oVtZcQgMVH5
B49LbglpTIkTS1hHIBYb6Q8d1uDugoPdjMtmRxIfFKMuDqH+thlyqKY9Z1JtovvQ
jFwCY984EDxtJMsqimOQDrHw5WhfQ4o33jBcT8DHGXEV4jWF6T0sqlP/k3JMRTU3
YwCxbsIlaKk7wwQ2/w+CgxCG1Y1Pbn6ltKsVi/+1TM+agZpcOtrPOZJS+ajxoknP
V2NShcOV/ZIzEE1v4noGytISSIp0YlBYBtl0pbn84YyLuQEKlC4g67Q6KZKfAx9L
z62gBq6mNf+KkRFGgcZC8m5Zy6V3g5qiVRxg7w219N22abqn9czHuQpjPknk5/kT
AofmsHhmwVw/rcPXthsFBJGiOkgdXbKYOK4P2L/jO7DSPB4DQJO7O9UDC2BcpR3w
6qWx6148fyC300FyOSN9W9qg/WpPiSMaPV8CaQsoGNcI+03+j0mcsySNravfZpbx
BFXsupe2B7y8f+2OCrdCh5+Dd2mFdY3y5NW7O6zcQCn6ZBUkqosZq+jDBSVl/Z69
s+LdV03EShwCgLb3izSHla6RydVtD8BM5EIw/j3WlVwktOrJDhktL3RuTWRXMqqv
vbX/mWYuviDvnLBisMzNU5+CG6MCtK8QtEnEAzjILGU+RT4qXrNTgB0UB1gADsAo
1qYrLj33pInUcL51xP+DFDOTLYPfJDcVcJv9o9ruRve8bxPIvqC67RYzYIVav8Gd
yrwt/w/ia7UGOnKkJ9tixkk6LZHSbTvXWH1zmjJjWbgGpX+W6HN/lHwLx8USlWT8
Ic9D7/ciCGBLwEFj7Wh57aXOvSIFedWIXxLeNfplCbODSWfrc+h3YTh9zXhkWnHi
14YKzNH8FJ2Pl4EyHpl/jLyy7CO9quiISbdXC6eX9jSxPAQv7yzjW9JrwriyZVMl
JR2m51oqA+8fKIQj4ATlzTHxxuvss91wTB1eJ+cLQSpQ1IH0qJYU1F0UWAbWlGoz
PxH0ULr5UX7OFgaXtqGLNskKprUnVbc7AsBR5xVgIZA43GYlqKZ3LmRCObpVatw5
QsyiKdnLpPQNJvd0akIa/SMtNDeQMeQEKwpGMFmJjC8jc42IoCMzxu13HEaGc7Pg
wUafs3OFLZkn+sSfUxLHIVs06lnBjimWo6N2Ahd9fKuxmNfimtKwhJ8jlfYynGf8
MenKalqSNlulDmpVk3Z2FLIrFblAS2T9JkmB0+OMNoP67dRdpQ737zw+RObYKSXp
4d+QDqLZojbPymMjuo4ZeryY+2xBf4SlBgCTrtXL1gbgISP7vf0lY0FMpxjnVcXU
1/HaMAo88wdfME2Y0Sgb0Ti+NJv4gSebEsptpkzxrZQqwAUuDII1fk7Dspgp77qa
iMSH3321uknERacil5kdwmFE5NZ+kmhZE2XlmzXBgHoKWXVbDg0l4PrCA/dbN28R
EsJgabeqh4SD7gmBjeL9xHKXpafj1a6jnYbgK2kbd+m25hwzgX34J61Q8anVrVRk
DzcKPw+3Nw+T949AH6+FX3cJcPN41SJtPh2go/p2MGv6NG6xbv9bz0Bb7m3TGuqS
BzqLoCgnvmcuHDL4/x39c+wJMvKmROSxXleH1rTVDpevSjxgDDCla+I4J+TKLRoO
L1K4a0FsDY5JWrIKgajnqjB1zRFdRFItD+wLTa5JJANI1mqZP78w9fZyjRkqB0js
wX8kLf7Bz/Yhn2Z1vt6X/t3P8TCl8fhOJp98/lH2oHpDPzZEvm9EWe1t1rNoi7KE
LvDqmFuNFYzHJgaFuu1SmDpaBsIYjsmUFz6yL6dOLUiypZ5sn088qIyqdLNjkX97
kRPsHQPCWm1P+vvrM9go8IoFX3SBGSUjhdSukb4tAoXgpjcLDBm+DcWceQ9ldqBg
MswVcdpJ0942ZGa70GEOIyuqV94dnAFOAxqCzHSmBUKKklBh8Gl7sxfkUT80GDRK
SdhmRfBbwsh6qOEm+Fe7qqb3kImKwjBgfWEoeyngWO87V+oDUHdzEJfS3CrGV/ou
G3Wmm8FJL/TnmqtWD8uu+MRqwewRtib8x9ScxSZ30GtzczF6teoF0MglLDDkR7QA
mWBtm9IBUZwDgrN5LrHmEf7jQkVy2eqe2GZBnvIN2JN4uy/6N81DoYPjljh+PZ2P
Jl/yWdEDOfV3xI9ika6CAZ0+J81gS8fAwGv4dTM5RWEFGU2J+xuTjga+Syv9CqEj
0ZCQoEgZEjjs8NKe9YMldyuUXLXY6pXmUSe0jk5dQv4S7t+8bwN7+yIxY5vtpDyq
Q9TXQGegqgWCwhH5gOrOEK1zQMWA7yTF9MMB4AOeqSDAnkUwnF5j/VtEjSVf7tpl
uBXlgfdLtrWFFkkpC+Vh1MLBEL/xoiA1BEhI7t6pzrFgrm3ydAq5c278N05L7Df6
v6Tv4YsjZYqiISs9xecTMR2mMBINGqtSeFKRZq5GwqEkC21HpA9f6fzBbJgrCcgU
i6Xd/Bxv6T8gC5TrpmHAa0mOrIUBxKRMUXU771YKf4/uUQDsLBHaNlO04j0KBlZO
VU9xHZIc/4wLAtuhCrlRuNIewR3hFMWCsdn17fEEHiLwgvPrREHwekPSgxfGDzhL
V+3TRplvm3VKa7d7y2BOcq+npIi6UTVayrYsRxHFoSt6vW67arUs2e13UDysGyHG
TnYjr8mVy886tkmo3Oom/tl8Avu9oYwPj5yEZvPknz3DrNucqKxU62QxqNNDhDQz
Z5j5HABUuIy1U/aYPmPixSJHM+AHnyE+NsShOv9lPkdI/h8kb1MiFuO5bRO7I9GS
N0omuDWJtvbALT6FeZLz506cQC+IbCvRMb4PkhdRq6ac6S/D4Y3wPLIg2RSAm2p7
rJytXXQdxHGcjqjUZ2hP9rxWoXETp9kSnKTv/w3hIwxlEYBiCVwu6tKa/yEgx54U
kzVyex2eihiN/7bZ+Re8sCzhH+U616G2Fe6An0uqvzN4pm7SRIw3y/wfQLtERB5q
8cLiNRHtHy2BLwIqRCjBhslx2E1dQNguy6p7RclX3FGolm45EduudMqtPtC/3Ddg
D83o2G8s2rek4EGNUo7zzZC4Fn/aGxkWOlgrrbPhS62uOs5U7MfSRMSYoUkFFFOs
hRi07arW1aUBrahvgb5W3y9V9evtpnnh2AJalHhKXioKDvh6syqZG35mg94bhUYi
865aqLwe2Qtfx+JNYwhmM6sK5lHkrafQBS3syfy4TZvfzCs5EAJ0uIqXJVLclogV
Vm1kiKkQO4GrstFu19xcS7SBIhwOz731FK+Hkvj9QootQHXUoPHwLCSDYjyjNjWz
0I1/hbmOZOO+LAEL/3SVwS+GyAq2luRvBf8wx1QXqBZv4WaoXcqJbnijX906hJgL
jeScJQzYYdD9x+lYstlqu0CftN2jJOipxBJ0ODRArTVThW4rDe7cHG5cDz0wJsRB
wvQTBIjtl090tUY/wQLYvzPFbhvDxUKnbPu4MPuDwopiFBV1jylw5zcMBgfqMNx9
beqcWiSiDavn72jmnIKKDOZmo2PZ1GHQ/2b9vgBRaB0t+iyet1WaAawt0rsDKgxR
iVKDDQaaxMunmeZ1aZJtEBDMbY/qdD48IkIX/I+J2qBCw0fTXoiChHEzVGGws9q+
+VPH7AbbIh+sLY/sI53Akc22hbrShX5nR+9IBOvFNHn+3bLyOo421he1JJQjcdsO
CbzREY18AIOfUHKD8NfirmrzCf5TwRs2Pqu+FvfmQ4saFPq+WN/sBMyvzqpv65Vb
aRmTi2zV3D3+LNC8899CbdQxqJmwD4I7PkLG5mjVKd+RXP7WeGQF5T82MPc5TGf2
+IhIVjZIt+aMQimr63J5WOt6mKMTe15Y3HeLPwroJ5SIqk1hNxTyJkoSmucro2qz
mfnG0aKpzyKEEHBKLod+1/NJkbXDv2HWdn15fjEK6VxLVzah5PQfRFgjpqQYISxV
g6+bud32md76xy5WIP2NWVpprsGPhHyv/ORVzeYWBoXnshmZwpeZ4Ox3Fjql43Ws
xqO9mfvHlj206k7Px7VycscH3kDP3DNjJMDvX9Yv4R7FmqyTuGMbPDlO+FmLIsGa
eDebmqwzmyzsq3Voj6JEDKWYTKWnTsZeK1g1JiUvYgd+AOR1KQ2+conxPt0NJ1+b
aQpNjR2uIWD0fyGH6EaeOeF9Ce/N7JvJiWECtSKSJ18d0T+Sy2Lv4wkuksGzhUZ5
po8zhs+IQR5gAD0wqd2SUFg/b0B00IhnfxsN7gn+LQR+rLGNols6xy66fiwxs9Ma
5l/soy3PE2AjiqvRf6rvupFzbU6TXcxh920ssV8lAa3xdBxC8ehNQWBA62vkQJNh
18vAnV3dYHzdv6gY+lXNVTIorUOEh8jg34rFHKLD/NNsEdL7mbK9dq3IWIS3yjXY
ZzxFSYcHYcrQ8MHJwWsT+pplj5jwZUXjtULnavQgg538YXiIUtvEtNCaM3ZsKnsg
6pwCfPWgLMWVBgP9cmjrhY81I+dz+NkB+MP+yTfeO5XhnpDX45bPjgieMaxpQOdl
eBODc/WAk+Pa5vYhhS1vjCu9Yuq7J+kT0qpRicRj8aWTGBh7Fim6Xg1lSoYFneEH
9FgnndnAZgcpsg1hZ8xSX+//oOp06/iIccKjCJDqu1QxVNu7fV8Q5g8jIL9v324S
8m/gHKrKqzItB7CzJshhx2+05Dkc8gbRhOSVkKZPVHhYQysINccWqA6bCUS2G1bf
C2AiofJvb7mpYb/qYmkWnATaUCUsZHIyiQPTfojQe+T00EJjPOEgecPvqLmXas+3
UrmQRtDikVmmrnmwpEwfDTAEwtJKE2seS3jpM5DBnyawte496erxmkm7hV8Y/IbB
HOEdEeCbZ8Sw4xT53VRljWMmNqQgfHlgm8Pdb56nWghO6q7zbFsLEIpvMcZsIU8Q
+kajb8sEDCqS9O5LrtmFZvQ/tZ4yUbSVrLp+s+x5aNTQGOPo9QIBAZng5Uu10MPl
fCzAxCKQutI7js3OfmSNnL5R9tC3My/zqaV2mun5nR/t9MVrK93oAKe3xNqa3bZw
TEVWgT02UNsy/ZDDF/uHq8CwUZFwkyWr3Ak8CPB+iCM6ElyeFmvfS3PYSWcLjxyV
fWpWNgs0CVQ6uO1+ONhfPb+4bOAG0jcz7L4kVGVQ71KAjlTlYTen7e7FBHAtHqZj
r+RZIwNBPBIt43EkuRK3e1z2zQNwOz+xSemi3nz3qKkNZaSOLCS5XIzQvr/Xazhm
BahiKLaNJkk+zGeTVGq/zk//zBVjeD8SbrLICFi0pK4QGCh4M7yjt+vnmujAFskH
5KT7ixutuNBMwf28KxxYzLsGH8lW8lKV6fnMLXmXSL/dgrds4/qv3zKxIOqh5EW1
joNq1J7Qf2c+h4UD04xANGdQvwD27sCY3P1yXUsBPcEUcCTMkqWEEPum1ErwEjdt
JzIMts8XXTw6q64GcNYsgLyrS+rsVwMdtBtakT0UsiSjtBU3/4p49hdXnajtba6E
xq55o4hSxMu0bFR/4OSNCphTfQSFtB40Ayq7w5u6gc9qUmFsmcGzED9mrq5JVWI3
OPTEzev2NEh5Q+DHC4IKVWzjIwGB24g4Zb3yoJ0PHizxwmuMBHJmkrktDnhHDxws
Rs83RJFga+6l+krJgaj8ZmnFmwQd3TYEW+zIJuDv5grCAstKJCBm/bauo0NaepWQ
6rmOXcGJBOHT9g7FzO+IV8SqaBG/tvA8SI6Fb11DjrRbZzPDIy7lnmP9V7ATnQ9p
BVcTyqDnXcNKWErkszyPZ4QwMCe40BNF7aTmMqYJRAtX9gagblYQaXftJDgGMgRW
1WCX6wiL9jSBQoKDkIKlFCB4mu5/9MLSplbeJkFA5N6Z5wIRvBzMSi85wa8MkrgO
tlEHYGjiQiY1HDYiY+Q3IIV/rqgIuPmokoDUQgKPRHleM0hpJTiXbNIrPtdHXwdD
C9brF0VGPb9LT3hCeXU91xsWROu1xtIVQobp8yjlkayggHEvWpg3SFnSRWWU1GnF
R7S/59l3gu0NsMSznp5+ozxFcZ+A9aJarAlHtCShf/2js6iN0o+qCVkRunAlYzDd
P8ICUMZ0bcS9PgX8UkuXwNI+t2TxjPpYyfOEEzTBXn3hPjhUesM1Qx9bB7xNnCCM
VJfMEzf7AdsbzEKzMzPhPioe3AFrV39jLd+d0ztOPVMhQlhpJghHr+KRcCaVGXN1
NSW40rG/f+VcCWiCCCnXovenAA2AgOvbzHP+LSKfoX35cv29IW+hlZbZdU4NEdsU
RL10JRNgtASTZjPyg3AdTNgE2/MEIbAR4rqHsEoqYMYLkYavtEQnBCM5em9qvaZ0
jVvPRVuJ0XMAsA3WScZf1r45LpIV7E7UAEktjaV/q3w6NHraY8RS/XNqLKSwGYC9
Yq+qtV/g6cLD/A2tAHEKbdnmzijRG3qZk1ubMNghwiMdCigkEIFqDdc7CwbUUBHS
Dli2mPuCcqSXHSTL4sesvj4QlHRjmqk7zW08p/W5jnBlODo3qjnipY4ixA40U1Zt
rFqxWXFIQCG4PpvTWcfZ0GsoSgtCqjk3e7+Hl941xG31U9iJHxeHG80Byr4l1JBF
WeCuWdyaDvlYLwDUqdc/WBC31EzzVDn60qsiVk0b/wZPYNNAGgL6n8ZDLEIV2/Se
PtNpl6RPHV9TPcWN5ty82oyojBK7738WXzQUn0vzWOdr5NEhenUwBFXcn4TfH48m
aESvweFQp4VnUWznbq0Unf2ssXiZFUcQO+L9XX+TXUOT/V5RTHF6OjduwJVNNevm
KG47Cjb/OH7dmiamjZoAMyIuhHBcoXwPPLS/cjwkd3ORIJq+pZ+YFErbECes+w+v
6LREkr+HVMvaYZiJzuMLsO007ARY2UtH9EcajgRXS/3ufJDWPQJslIqehFc6GHVm
V46cLmJhPxjOlHnhfFSQjbCcp2RAipocBid4CqbiizUAye9ubYdTHb+87ZeZbZI7
v5QnRq8LgkR0Hl65Z+wlJ4EsIUcgkcnp/KtKkUYo5qNUMBP2oc5V1AYE7jw+2nG3
kd1zCeUX59wnxKWoGY+BGrx3ur7Cqnsl7SwTwkrI5O6DVkQ130VIE/qOd6pZDihW
iT9aun7cJiD9PZHlqtcw1m8b3iSuejSpjdkdXspium5Vs14IhDCRnLXgUM6jaFWn
Uhbcz30qU39pzeNn1MbPRpAtUCh8iE1oeej8CeYD6QIrnLEMScoj3WVimimrZuSd
7cDabkjGPmWwL0ez1YHuznN5xWVTPEwCtmr/1PoxmNBZLY6YkvyRlURLT7bWZ+wB
2i8VWi3EAtdQP0mJgurPHxhosMEMyiNvtiVEQQ7eDnCeFGMZS1lC94ODFG3QkWe8
lNW1awP576o8NPFk/hIT3DitZaF3T6Q63clk1IP4LrA4eDtl/nURBNvYZ3xAbuIj
Q+kIknb8rclVjGaXuJFcCY3bGj7hbu8w/08401D/Bu34vo0n+DAsZW6+C69Vnyrf
lQ5sNuqOXQHf74nkbT0rtoOI2BRNTEOL9PvxfA/jdh8XFPE3VF1ZNLh1W9SdM3lO
voUJz/PrgGjrgZcj2GwMcKWnkncqHa3dZHPDNh8yuOHcbZbNlPkmOQgOcKcMzV3g
vXb2K1D7pf8sN8MM3aXy0nnsaC2fTiinxmhnc5xvota+K03pxGHCJtaRHCz62MtI
NxWT0C7bTA/NmbvXFeJOZfiYYE1CdN6V5bWBhs7tYL9Q+BDb/oh+C0kaqo8g1/Lj
qh6mP54Bt3Y/3/LZ+xNwCWHOVo+wUMg5GVpMpZvIozWNWW8z9iIFpDpiq1sCRkwG
BZ1drowmjHg5TCL3iWxXzBOSoej2QThNkFMK6jBsOWnc4LzLbbRdmz5bWuGbS/Pg
Y+1bL4MUXDNRgf85OSnr+B8oi1494q4NoMwbl4WhSmSy8FAlufkANx7dBys9uK5X
DtnJDM6sxUZg9NFfNCcxbjDtSWc/zP1t3D9JHtbnK2efYQRFUoK3jXMaxcEVH7oy
mV7q7mMF2u4ercnainGDx0ZRBg/S7njR16C1haozGCWyDlrYzRyN3mmQYg6bQQzg
CSAIjKmcVKczfsv9akdjV9qoqy1+yHBhNuhbRJc3fKZ9vr05kRul0N9jlAXrJL6y
ypAncJ3F9Br5CG5LSpcsqYYGgtApamPYedtiHDI0DnLOM3sK/aMPbD5/iXaetNsy
fnMxamInagN/3T33KEwA9JZogn+b8eClYMtRvYE8WmUywuiuGaOS2DY2/JSDx/jx
0fj6OsjeB/ZqmGocGHRIVPNyJkYTu/Vnh+7rTU89M8fSikyCVbiXmlUj2+kfOjXm
1BHu+CcAuRNEKwr0Ri23fjOfGL/WzcMyODPQJrI4mn12xhsOZ589/5yVxep4e7O5
twT0aA++hGjH0xJAogE3JX4iTTFN636vcZZFWkOhHO0VXiBKtLNufioheUTGJK13
jyL8Z/khd4wkTN6uRZfQKnDFn6Xt8BUBlSkUvwTvghN4E6R1zAiUjpTU1BKoC2xc
WULT2+mJH6pfX/mZd9WfB+CG8m8HhqACzZ97qXdu6sY7LVR/9yBNTCz8A7dcoCaw
SdZmDk4iCyYPOSJyw6JONsnFtavVjsUTdcTaIj+eDXXzMsROc/uVWTcV4qhMacaa
L6UHelkPBdtYUCaB3fU8W6ymBPnBtJQmvOKl5tsTws77GnSrK28mkh/BDQJRhUtk
jnR18zMrYTJCcCsOUQhCKS/oZ1hLwEZDvE1E+Wc38SvWr5pYJddR7gJEubp95gRu
M+iK9WNR1MqjJwQWGQKgS39jNuPyy6ZlgMiEkUsLIEdY9EDxlbiTujlk//EvCCRW
saiZanKsu4AsK/CRdfAHnB9RQ2VLtof/71SrXiLf5rE7w09naqVaFwItTqesZpGj
8h90nALmcthLCMq8egCr8xg79P39xgbFgGxgCjy+/JSylkBOhP/NPw6iMAw4Uv7/
rk6xr/GLfaPC2O/aYTkIb4DWL+VJXqXetaZWq675KoELB1sAFr5uP49k8AJb8CjC
bb/FgJdGBL1Mg4NpPK1ypKa3faVZ3buwoevKH1h5Hj4RkdPZcfpYm+tO1whOqY2L
cPYcPWZkZ5WiVK/KFoiZUSgYWMgm97yr8FRvAIbJax07ePq5WzYhns82jqEUkS6n
phwgp1piG1v62zGbn2ibTmRVEqND8oZ+Wyk2OxucIEFzmdlek/G8/3eqjhey62xd
PJNsLdTBRlSF3UxCx1ZGmJ5ZRYodC2rgJrfPbjHNn7Y06OCG4DE9WCQ7Y312vhWb
gWm6XvI+p5hnUQUAchsScaWbu4x/6o/cm/9/q5Txz6EdHgakD0yi3DiQ3tCzvf1z
/MOYNCht1SaqmwpfL7pUMan4vh/vHnzmY3sy6dJdnzLfO1q6PnLRMJELrY7M7Sdk
oE8ayz1hGd1d8Gv8BFFvLewwIwAedpwO4Fp5jj4Vs1tVjN+Saoj7s6UqOm6xspeo
+kiaFT9xOIWN5Zpsj4jnT037AnXyy5Y1Rj0IcBjiAcC1HmQePZt5YonIGoH7NkUu
dlCSfK+otCVPBV9tXa91AIL4XQjnPLm8yMi+ItsPQRd4NMd/wmg8SVgHQAJrtyb1
CrsyaaxvGY7Hltrzb7QlHSyAIB+jTOVMVUrlTlrrWRLoLKiQG7D4A6qf/x+VHtdD
0q9G3m0IL8OxnFTrDhH/Nf5SYlZ2+eu1rRdhq2AmlFCkZTduMpxfu/1ancBu9/+q
nqeJyJOziNufQ49cYdG6hunCmMP1SFYvb5iVnm3EtcnsCPS4L1ywX9jyzAaw4z4f
Gcpt9p8EC5VPz6dZlRo8kZetbNTuj8O51/20VUsGLjHpj2bVb6fhbZe3R9b4umyf
o6sp7JUMccd8/v4vbRU91az/TdIWOAIRaT1LzRTZQqkxDkzNf4u9+b11a5HM384A
ue6ENmLvOCwloGeIMyMNWGaODdgBxibewm1uoVuyTpyYUwbcC3C2E62DxO+9anoN
y4ErnZzI+SPxRlGsx7Z669Blnw/a5ybmnyKx5qD+76lJCL5eEcIU3cOTTksMSNr+
yTBPR5rEEHwvndimBecsrF4I8QAqBKkT5ay75F3DRv1HrK7NN0/tKxa7i7x4Z7X2
ALrJPxJArclaluw9bxG3rPs2tBP96PThejyQvi5eMaX8wWtHYVRkE5OY2voQY9X6
1xrUdBBAvkAJIJnvjuf1sZmn8RSBVHbCJ0w+LBPlmzACkT+X4dJxDHey/QAgmgGh
05B5Y5V2XlnEsMEFEiISVMG8SWQO4atmYll/6WaOiiAGAYGWzD6CXwjuTcUZvt0P
pfv0rbeb0C684I4Mk9c713p+BrRsEvmkumPRVHsA4n2mXtmR9eLNU5gD2rBNsvMH
O4EeZ8WSsDWrwmN/LOvQfDwcK7K5ddPRVkqhV+fNz65sPE0mn7cQJzG4G1LBrbr6
SOs8937QSIB5kpn0WGM97miB+OJhdzoOPEcoBnHgMEZCXKbo5wChTcWR69lMwb7w
GWaLSSZ1lqTo9g/DSCn0UrZuGZQZdUfoiqViAfb40Xk6iOCCNX6pG5DxaCnV7QxE
VI51I3BY6a36+vccjry2wZO1dHrionK1B7zWBZOJGfchhzdYSFPpzMzzXZdktZ0+
ZjcrfaJFzqN9G25ylbBPG4RgEEy8xk843wkq+MRWrK7aJ9FOPPa79mn8uYY/7Jcm
daGGm3fMc+EgJDtFH+N4OeS8r3f4uJkSG/KFurFIYJUtv2goSq+flxmldrwFkqdf
o5lb3IG7Vv+nHwIv5ERMTS4+wd05SGWhfaPzUgGO3Jq8rqpU7ow3YNLbVf18aZnG
lT+fr+4k5UdIM/begr/+ZCLof/PLZs24VXRpYLD/dCqdvZxAcuVr4y9kxUdODP0L
B6ITmsamoVBCC0Cx0QSj0P0Wqllbsw345ja5A78eM2kh19FMaViG9eONOF7kaygH
rvSz0ordwvC/mEihv2XFaBgf1rZnUT1wGtwainD19yc+o9SNuxZXgMaxQ6bk6AZv
uc1ILnwM23Xn0NqzRAdmHgwq27RK3hkGejnRt5hMfwhuqX9NKW3XSoYozcgCupgp
siJV+moqKO14bXLlAyorNJQVCXd6BNPM5DYkFua6E83qPzJezyhw6hWm6TWYQ9rQ
8cpSZN8DPzdhGOjY5bFA3NIsvE0Vub8/QgMGvQJOyABAFybvN0yzJkTwDvzRKOv9
fk68lWgY6MlYb53sU1XMEzsNmK0OyxEdFCb7/SSby5gy2azA9s+W8XoIXvnxAMl1
Ri2KVHa1cPGKhdyfqBb6lah9DGTsfoQw9I5+LdzeQ6uhSYRNe8fQpo6m48hT7nbB
U62guE72E99ba0vofz7ThxzKVE8mu8gP/z7bT+l3MuGXRmLMqvSO3AC4AyOdovKk
0W8N20fGGFQao+e8Q8kfpHCXEPyEAW12712/ZrzQClgQ45TGmd2Wt3t2TBssh8nQ
8lgq26u1XWB4zVw5aK+caPcLQN41jSjVg8WmaFIYPpCMFEjl5yaUJ3s1mEyh7s+F
mmGUPDpOooviw2dwpGHgotDn4PL4rR49LVr30HzEFF4PJmCNpGu6UJJNJmfRwV8b
4Y7jbWlbaI9V5J9D1aqS74hGcEfBI63CaUAf8cU11iSEbN9MvSF5fbPGcmAimcUg
T2ExLB96FuW/niX9M3X7xoJ8FiIeF8GEpurkBWJJ+rSbvQmJouxh/7hMWr7oXJBr
IN0u8Z6xykpMufg0NK/Ru3wUbKTAfR4CwUltUI8HP4mNeBF2oR0Cl5tylgTU6XdA
L0cTeZzavyLQ1qXA7ZXVTpauPUBs+k0HR4qkXy07Anblwp8kgVuk719bQ+qVA4GD
b6CJUFHPeJP7UnBQlnmulCFSkeAhiepeUP7qnGwMf+thcy4g0FPwEP3SVhEGgOWc
78FJTIkHItcBtm5vNOiG/gylPOUl2epGQXyWbuoV5CBnQcXdvdpgZzw2kenbbFLG
OKx5JqS456nftys7kGqUJJn742Ol1tO9F8U1DBRdfgw99uxG2S8WnTb3rqNMhsYY
VNE5eum849s2jy7ZGXhztcNFnS/tE+D6VnwGEglMvp4MjSQVXDZgRo6x5zUqy3zE
g7rZmjzzk+kz2bLa3qlKce5vdbsu0lx9yJInqzYf4yCwfw/ijj4k/ooVKDs6fx3Q
T07fnEFZQJyNRnw6R9zF5qmixgjcrOuWBHbT7Oq9bO0/yJ8Q/yvImFC0HxRjdUgi
gsnYG8AyrLuyr1yf4tHy0r8FYhWu8cnRpc9HRkQX5VDcV1aUodCkhKAgpSoYSSTx
MEYkHlvPGqVpUIqkUhr1eZLa8TlEqmSRRKw7qye718zfai8DhlQMgxgXnHgQkSLM
bpoMRd5j+J2Xbeg0YU61XszVOv/m8z//KTRC+5KjTwJFS9CUYQQzaZop+bH0X1fP
juv3IQp9+PeSyzSrwUWiD4H/d8LP+7+hU9+pchibRJwcADVsUFJFFueaU2Q7a3QU
jsU+jRAUT76nQu3XOqVV0bRDstzTenL759KkrHZuMm357T2eSFBvKSP42oQKaGxw
/i1FTApc0e2/l7sjkbN1OSL5m88r8KqaslXCYHM/TRdHYE8AZhnzwF8rF/4/emIK
hZL2BBV4Bgi4beK7YDIeMwxjOKKr/F3h4YhQERsk74rY9iftEne0/IOOGG0q+UV9
pNbnZcpimLip6p61392KVSWV+ZLARErgxWF/PeQ+XtKVfUC4Wiv5ZN3NhyLK0jcU
rYCbGoK3026UUN8Dfbv7zCCTqAyWcV+2/t9PJ5IqIHZNZDq6UAFLtyYgSQIHxtxl
7BCXR+KfuzLKJ+Ddboxg8x4RBldgnUsKs1n4FkEDvuQXiQFAT2N9L8AGXFBpY4f4
zCTxB5coO5A3uFebFA/w2Q4Uk5Wyc2AIkGPcAFQAnItsvHSGZwWLG2AI8nyX1Jt3
P4+Z5MTojiivcNs1eCOmEWc14I1iegIfyWqZZA768bRfhCznxJdOsZjO9pgN7/LY
UOcjj3o/jCnoWK7XzirF8xU0tA8EZ4vWiO6tLd8JORZA52Lkn2QHhZTJFmuFWSXB
KsRdjnSe/vhtDtuWAGiYvYjGapcw6CRcwLYX7Ds4eItvWJD8tWrm5oLOy6Ft8HSS
F4URoRFBS0PCHeM1tQHJrqKxlfLncsGWQk7F3PyI6hTJ4yHEm9MpxKO7VmG6FrBi
Nn4kcm/kBdGYk0TP3+ilHT/UDkzOnHkA3ntGHZK+uk0S4G9xegomFmvgww64fWcm
6rRbbCIO5KeFk5hiKb4t7bQ9V3ujNjEZepu+Vji6gPWE70yem6tQA865lQWtKQmU
3yQqzETtkNbJgxsozUxx3DJWFEI/SIYhoFDeTtZ+PyCL8PlmmCAgX5v8l4dl4s/v
hBS9e47l2PzeSCRgZLjQyzMSqthOCOy64nE7qa9txs9gBIQRiqtHcHzKEf3bHyMU
jA15n3Cfex+An73D21dyLsXqlP8ySbs/6GoKdY6+De10M9oslOGeDNDnvqzSMOxu
1SYx0jjJ1Qdb0jel681ETchIvGuPG/dfKYs4M5UnWB7Z3Tt+WtTjznVTZeug6nx3
5lHNdtRa8ETs2TFZkPfZK7wp9xrtXHGg5LQ1jpQ0BpyRngU6myDv9hJxPiiG6Pq7
oqsT+5OAuGL39quJX/HuYFwPrVp2poyq6R8qw7QUIRUCg4Ei7mN/Kxuk8aiYPtjl
sgTP6w2UCl0HJsOJyVnJsF+RuG4Qt9cml1C1P6BvVK8YbaHKcyZzcWb9dDydpqyq
o1XjHUPdLVmqCR/emCOgKLTltETZTaSNKKFl1WUjZqteKSxXdXmVispghjhY4sQn
rvYcGD/rIDdIaLncXPlaEV8kk8WwWnimmmFSTbOyplUT2fSM2hPEmEPlirttE7wq
2tcrMaKsxtG/tbni2329C006hdDnj3J6tRuyA/QFTSVkA8mtq7+IK/0VXO2C2GtN
3eoffE3bnou3dY45PYoZxr4CQOwZUpINJuAUYdXQmmb8LlG/X5AqpRkr60W5nnvh
c+HvKURlba2DLLPJllJAo/vTfiMoCVwUee8Dn7CPqP1gDUCywgWglyTg76ThcFKB
Q+5CXa9hlvuMyI2h9GSMvVA4L3gNFnNr9J/xIFgywsMX2hTGlrL992WIY/s2pi/P
96X740YjT1l0QpkYB9S0Qv733/5dibLiKqLHT+znsHuTJVgpLA4Jc/Kzo/aWPVNW
pQTh96w0XLjDzoKSrTnJT8ACTlwO8X5w89aRDt7Jufnt6ojDsplVFQBSLmGLQAKk
bZtF/29ik9OK0AGCsh+TUlbjrd7H1GTYE7mIPUYg7gizcSkj8spK/pvpuy+OgVk6
QBG5vT/8otWnIklsEBaV9aifOukvfioy+2UyMwhoXLff0ecx+V36DgQwVA3Jc/8S
ThLGsyKC0bwLkzrd/D6SZ3MwhQIaA1/v49zMjBEFvD0gywvtJfXhnql6rR94Wo8N
4Z/R/dC07Ml94t8FopseHuIBSwa3mzyDhxdWyW593Qu8Qh7jDPhFPc4dHs0B2i/9
3BGOHZLpQCV26rUXKMXjIPSbEUp0fPlE0pcnfdJMB9deB9EaFRCPS8u/bsGjbIeF
E6pDY8h850JQ806NV6Q7Ea6SvKUgXqyKGKJBFVL6pS3GPzyIfUncm6yDU3aJjn67
xiChzm5hNupxntzqGjXQGPHFtpKWRr1OqlOW3/x0/NblbuLG0IoCE5E22PO7qs0n
5FBZTaRoBHMa1e4Zyn6Wux9PBAgI+FqKWnp4gUhfBl41y/bFwScrBtBKHSP+FHgu
jbOTwsUFMTKitjhyOsuhc3hup3Qk5nfYo5Dj+UVn62Akuxs+s1bqDbHvYsS/yW0Z
swrSjzpLPvb2pKgVMcqF0h3MtQzBXgyTQUeo+pMjFkT91qPSesQ2jjVw27X+gxrr
HnbEQEg0i0D9Bva1WpXehJw8prYVHHRZ7oOObEpEC0rSENS57YQJ5u4UnB31ATxm
ON3NBj33wrQtQoQODrsPstdq30zYfITS+AJJPy3WGv690i+Zjblp2NXqqIPNxBzN
2rNULGV+H0gd39Wivdh8wJxa9B5jAyLJRQyBGrFghu0XRO96XoLj0Qz6fsB8mJ7P
10LeWL22aKMBiBK9xW0K6fnUGYaDX3GmDjvISnjTbv9aNrf8oj8qUb4j1tLLBVam
KU9OYd1oHNeEeEH5JlgFaIVdMxk9CjjL8OgmgByuP4X1t/Th/N+Sank3vWnMH8iU
TnbHokKo0O3sKiw+bNStXgWu5Es7u7ex6l5jX/5ITktVUL09KgCEtWmO9B64lSpb
M6dcSer+J3o1BVxaFvWzoZOhYV/g27k8z1E1JGuzWXOLZbNg+EpOXPASO/wQmwRs
9O4HHS/AvpCWwdI+0Ijq3zoJtErgCBsl4+E2/qT2gtVi8x6pCz8anZ7MfbtCDX44
ttyb+fWVQuNKo6N4gIyvm71YRxtyZoXtsfRQMMfZGt/TBYZuU/mESvGDWdYEiRt2
KNgg0s1PvGXPNNAg+EaRVM95bz8CF2X0IuLjWVJQIHpjCv4nV8b/LtRUEj+X8ddN
i9KGc1rnf8cnWf5SO/jhsXvnMlMc0zdNXnkFuj9LeZEnaJ4WqzjU7v7SggfKtTf4
CwTPf9XQCkzkt9OgOWwoJQFU/kgeJAMuKEeIKAM4M8vPmzJQkKuSwhAdE516wM7a
ru8a5O+/wydURK5RhUo+WSNVd96h/iMfq8fYacZrFgumswP3YfbdymBishjf6TiI
ugPIda7MFvJLIo8fOL5g6EJsj55MrPWm8PsvLk8L0tfUBkU47FLaGHviVWuN9oVv
l3H6gHtJTG8mZVcQWZmKNcJfCZ78dWzU3bomf68CE8RZlbYidOOTpKXcE/Cmgruf
4rpvnZ/4R1ups3TNYWiq19ZdME2KpHF68cQEh92zf/YAODQ5nORhofKn5MkTrBuv
Bqsb6UmwHxKW5EdK1xP8LE/qAhMPpeY7QK3/yPNeHqNQTf+cCQy32iuRWTCTz/hO
3JGjyQT2XAuTcRby2M4Ig46tfxCAJrEWbUron4L1Xt6bY2KdVi0mg0rm/Jwy/wzk
1Oa8BV+ldA0QVJsJKjJNktxNxye7c+c6HW4VmWrB+HG5InumnMPzzHqU/G4x669X
GhERPKTuV29/cx60onIPgKMmmpEiCB4o7w7gjEtjGhHFuUddwcKJOneLmThfy0SC
WmNjTXevxiG8C0IhlIKPW2vpLMEHF3993UMqVMceu1ozePrVYTD8zwNmNgS9btjw
blfXFe/haerEg4hyHem2QMIx0gb3H3TFo5hCMqtec2boPSqM2gO3fnLQIzMT0j/W
6/eQL4ikE13N19DDgCFeKXdQhAJPGC7ia7AUfMz8kzGn2GmlL7a2mpb06syx2rSS
36GfJC10V74jO6HO2HlThldzZrNOd96Mirwam6mMrU0uiuv3layLQ0CFojByg7n0
1/buFoviCAVM7T21SsbzjbWcf5kMN3XbyXW+Xzg8KNS8W7xlliRJV/RgqUrZ1IOd
+slTT5xGRwjYR3t5rq/NJ89zNRHAdFnJjBRdl5vphm23nMgDkI3ZY0QLPo6U62Nv
Eas9FESqK4fGJuMIaI0O1uYinVo3UFjkIsWQL7BZ+8f55Kt1JfkBRIBZC3b/YGxw
SrmC6b99MMl5pXwsbHSm7bN/zK9J2Sv3BIX000JKU31xCqFl3MW5D9EYtjpcd72F
SuKlFYwh+24YB2BDDygXAsqD6OpARwEuhXJYGpdmwdnBIB0Tu6kPg2C+aEygEb9j
IRMxOzwP/0B3n50rGn5/NltZIUBig1EvcfskopSU5iLuHodlO1bpSG1CBoGobbyd
jjGF+NnXoMA2HdNLFUe1HZXQ5Z/99BUGMDWcbk87RVbqumprd+s6ljeGkyvjCQNi
G8sSrkqNIaYRH7Zy0kmcTPE/bqPXi6zKV9TbyemAGEqG0RPuaFMIdPzpcgwINF4/
JEgHmIwJnZkS/ZgCcktW5n/UAUKq7dQZbkib+PydwD3uNGQ3Y0tlqHCVBqyQPHip
du+tAY3eAfOcsWGKPe+ceM6i2MF8WKmgfl4vj3Mjyp7MaETqNts4Wcj9//uyUdl/
wW5m7FjDjZWvp7uSuDlRNj2L2uAFjMZPgwCttX2sDFsKtksFlh1xRaOy5LPCFfXS
VyounQZLk35U0wuPj2Q/vy6WtoW15vYWctYMhsOCznB/5I6EFyy0dqorZMkwUamn
sFmyUmIpJ7BW7EALbzdCfzRX4v4SEKjFNMxTlUslkCWsdAFqBhtdq4GvJY6a6Xkd
nXUaNhoVHqHzzu4nfEq2eyRiLZNIc2bvO3fj1mVcZfJUOKcgHCGQicloYBI9BGLh
2t9+JudGZn9KeNes2vgWN8xadpQ7x+DwPk9fGXPfOx+AI7qefHtR4xNG+McYjTss
eQKwv+3btkvY6cdtPOPakpRBPwWz8YTpb/w511qcRlGvQMTURbIV2PaSLUA1q5Jb
uBfwOwmQ5XXB2VeSOcmbaaV8mgRlRv3ydZsrQmwMJtaT5kfC1cDXxKRAxQ3Co2QF
6MrwVl2w3Zr46t4YNfZVwLvA26kIomcQbUQQGTUsCWXFvSKTTfruedDCSnangBpB
LIULklQG5r59P9fjWVUO1fuFfzKJkRZ9/Qk6epfHL8k9IDFUgLuojqgWtN1F+lXP
3vAXe2+q9jO+O/rDhGnEjRuKUw+94/gz9ydOHkNMjiYJpHeZLXok11QlwiAx//+E
iiA2G+VDOotafNxluf1Up6Fo+qXqbYWr465CSTxjN8ziZ+7s0pLjaSYP2qr2kCVg
MoyqADWNhqKAf84F2kZY9EgZ48ae5vLVr7fGzUx8U8ZIgCHvFjh7cFV/WeD5Twip
NOc6XL3SVTZccP1S6gb4NNgIJDj218BJCQxwZTbgGyI0YBbyfWExybHiore9TWwA
Eexo3iUklzssv7a0M6kOI70O3O9DYoDKFIqnz/g7RAzC/ZPO1otxS1jR4lh1acuN
RL8+l8hOCUSGqx+cFOIy6ULrXji5rU36by5v00/EyujSJho3j/13gJSSE4llFY/j
CbAMEJpbdFUaOHvrCFNCi64lFxvO32z6bDIgS9eaDfoXN5gCLUNz+Ra7vQEXn3lv
m4CxXJuzCKith3UhvK6VoOJFpNi8Z/i77FXNMrp8bsk1pixP2rjbgswb3rNzDYoQ
15ntaMwAkyEWTtk/GWEvwv1IlF616aroZDMJISB95dcvhEqQXFGdmHNchrg1RSvG
c1C3X13J37obYVJXXA7uLgYlpDIZsp2a8oy0C7VDS8STITw4Ot3snwR3JgRHNByC
1K9zSACQ6G7b7xKGYPnQqVh6+7xSi7CsH6b1c6ex3UvwTyoIHSThBNpFW3Y1oQuH
NN2VwtAROHnpzXVVEVZJbqxJaeAq77JDeO5Vx3NaJeD9J3oXWkPG69gpQ7svsEFh
ehRaN2RarBSBbm+YObj4UzsFOb830oG0ecFgYAQslB3ZHWoxKHWwJx0rWQo+ixVY
QxXMh4OfjMD8IjQxAxQqfLnd9NVEeG4QNO38t7nFlOC9Ry51KeyGdckLQfUY1xKW
4YyEH26+WzQ59VhN1XWPdID7GSsx72W1PflzZ7w7wCXr94mxu7k5lU/NVxS1ob18
1NhFL1LPyq8CU5nXLazt2LKUsfUVc4f/dvXyZ9X93Oxt9IuPh/fkkeYqstpxWXNv
o0uzWpB2xtfw1uhs5pIJ9AkuP41uA0ETWDXzrHhbmQFjp1wx8ncYz3rs7JUdAa6w
O8zvUiuV2vgS2wrcgTh8lRBS9kiTckDElLB8Gg0twjU6zkTKtjHDKhn5LI0nDZ38
vb+MHOUHsPML3snF+xFnzsRbOkYMUl1ATWLu//53aBsLY09is1ipKj4W+Ip+9XEa
I/Aplq1WL4HmY+13irjxe56C9W6MOcxIs1RS8tDLDbFdayJF0R1suqH+9QnaizbD
lbmPXTGOWaffqDBoM6t5xN8X6kUv9RZptikMdqdqDhtf8NnDVsZQXASAJHTUiQrg
4ep1NQbpT8I/pW6QM4unTZ2JfDqGcJS32K0s8aC3rjyfqmrUA9RYO6P5npzfwoOV
AbEukJpyCVZbiP4DIQF6JaZIubsPzd9Cq8Jq2G/0BZFq/pr35mh6EFuc6EsRJ0LZ
RVjFy8C27X439uzeKz2lc8EEGWHzbn9dS2ze+6ut++71j1Dz8CGucov/5tci4GcK
jfcYlKzaz8em523KtunHdv78X01cukg9GrSPEOoL6FPhvtGITOOkNF4+RZBucysL
YbRL3xju3J8CCts/s03bE4aiwkct9wsrttgN9/+cD01eHUDzMmdeBwrNjSPcDSBj
Fdqs/6PcyK3qxF9ol9rIPgmfls4Ga4n6sYP7U/kNg/Eh4ILy14/0VZ7LWWSMu42Q
74QaiVfm8TuSQduZ1x9IRmSgL82nJLfVf6/wcC8X+9EfwNiu/QmeJo0uOEst758u
a569BkH3aetQqibKgfMSvuqg0l4QuEKbCWmZLKSaMrPrafTiSh3P8n7cTXR4MgUQ
iZJdKoxSnTf0UY2OJ3GGTHV0kVh3sOot8K3KGNR/QITY28PQu9CWFhG4C8HfXrCi
Nr7OrNH9pW0U8wg1Y8YWoqVGAb5RdeQnwsuKJ+XNzKVCw78kryVqlD+79D4q3EME
+y0Lfjyf5tgSKl1sS1D0IIHnm0mORE5CBWs4Qh8obxWcjrl7gGnfESkb8TxPjWyQ
21FEuDbU8yRWOmZOW5o/exyX3Q/Ip0xlNGyoKX8TcxkmQEeDQyDx8nXes8Dyd8mJ
4JZcBhzICM6nqQ4dlxjhp4CCitQVizBAwneRvVkvH3K70AlsnvoRaIk7Fyv+bSrF
GPSGcyHCObg0LRh6pebFruqkCWbTeobcQ06Fg+nOXyJCOYNfcSeGqZCMV9qont2C
hxFzsHX3+lUWawSeFEkZIRtUflQEQ6M5BAIb6oamBtgoQ9iwgkukejKCxtDyoO/y
EYReiJeS53HRCJmgxnlfjtvh8lGd/H9lAg+PSiu2etCGewCAhL7vloKsLKTSggNV
fbpotvTMlrZWhlhX9GjSlezfFs+rn0uSrlpX4DdNWBKdEyGmJEeTqJV+7Lwk0ovh
RvqbEqLy4tr1iCepa2vLSAVIaIOw1VWFK4YVtRRRWHQGi7xm4aRpzMbwXxX1qBgN
pLQ4TJ2BYq6gBxS4RHDd0WGhfiNCc0jJugz9C2X74hOOTRF0g5vTzg8/+qmu87dp
CL/GcHou6C81uISFbuYEp9AWz9SRiOtqhkHaPS8vmKBr7SQooLw9kYKm/DnirBON
KQpW0tb/dH9NdveZUCN9zPmfOvjHYId5eHrrWeqBoXVMokNJz74ZIVx0koj7vvAj
zg8PasfjYuYSQI19jTI3/HlSTpkywFg8lbhaJFZQkB8I2MD6LPgVOlmjL1qH8q0A
FaqDKiphgxgLN/pvH7WWIwE2W+11aJ/udO9B/hkE0+Ad+fv62NhglMfcnBWqKMSl
nIT1juPEKFplQMIPMOuLOj2w5V60JjcOIB5b5ynms/7WXtVhifShAEODx5O8wP4v
44ZI4uwTf5pOQVvycrZ/V89QI5qsV14GYRFmMq6IQRZgXTEJhDLSzRae/YIecJRO
HD55CgMGjF70qgSs66SUiXvoD6EhNpRqikK1VdT379+duNt+z+2rdujmAHSI3aSQ
hePrMaf4YOy3jOn/fwzkRLJia3RS4s6fZEoiL2XqQKvaW0nid/K2J9d7Z6ulass+
YG9pysUmbhOcBp/EHMmgExet7IYkQqDKHMjGdz1S3Kb4atOKwEDZe2yuGVTZNB1D
2bPh32EH8TxLX7bbJTar3r3KFu31d2MYjhnR4I8w17/Vl5b2csD6GdKVxLUO2fk/
4uQoyACiLlwh2AZkvCWso0MHJPl1WQ9DPw+AWmTibjpmdH8s75hi0C+ykt4virnj
KgwpHDdr5ml2VjLom2LpbY+nizDVw/mrPrDPQzFuUpBVf3QCx1+FlNYeNTibF9tW
j6oA+4PM7lKVyzRJA7HWehIkOBJcYN7zedh0s4l9+jO576iUP4Fudblv+sisoRM7
aWJ+W4W3tBvTCAITrhjEW5c/KHWQZVuSHvROgkVqT4M94BG7TGJtGE/dp7JEXE0w
A2tmlj2bK9AtkcrEzQLTpYZ3Vbgn4N1lz1tbe05TmIjch7P6FQMW+xbXbiCYFYlP
2fMWoIOOfWaIXU2L91YHajn8Qgy+14htmM26P/EF3X1MH6Vvs+Oz1BO/HCuElmTb
HgVqKCiDZ/hu5HrCIKOWaXBSxJjneTPZM0Fg1m9XNbmlCrHpMWGqA1peinz8WRJi
xR+jlcFjS7ogZPhty+rZGS9TjHWwTNDZ17USBVQjTQR151fLfX9yjebrsNVjBJz7
V1gWLUJu39eM6ctdFXywYi45zHIbd0+50rRz9jChht7P4t0BM9HIoxoMjhUlSmtp
6z/ALPtprcOyRjKmVk+sBf17RzuYymUskVLXcXHhy79nQ3ULW4zzXOHEIh0lKdkk
jVhhvBHRdzmxXmflV6ueHZUS9LvAfOlpQPgdIonosFrl4/Y/KOw98/evq7xfBkrY
Ooexq3V5Vr2Qf7ZvvELiVIjDH0WlCwh03QYC1oMUrWZIyF7Ap1UlawUQam6b1Sfa
sy5uSAFdjewP4ZeSSOzvAxtT3ElEGpfLh2wbXmUjEedel2eKQWs9CtKHdulnldHC
10T93376coHouEn4iciY+8riMwL5cwN1cLQ70j2bmDGD51CvHSNo4CryMvTtu1yd
KzjfbYcLqSAGl8QfGoMfm0gmsAqzP5Pv4Fw0zffgxWe9c5fEPkacRntFUxy3ZMqx
e3G6ymubS6VKUpGPFrcJ0JNuqP89AVJUefU7jPUwljmiH0ClbjsxStMjV7cAzhNC
ydt/x1CLBEp2nbNeYqnmbJl8vjAvY/qR0apjCXXp+eH8LYrnnnSusxHlM4a4PCfz
AnDrfvoIRqzuHTzx9HDPb1J7cc8JW0wx00zv+NUFwBF7gm4djnIZ3Iga2cTAKJWb
lGld+bHqFG4AsMJA//fB+3ypX0hUwIx1HWSkHb28FvqDWQuIsuK6+L0e37GGvyfJ
5uX7g7LN7aDFeOTPqCJVa5Hfgkcvi1L3UXdwUcJglUFmHSOVsLmtKyG/41oGDzO7
yCBBR+f1q8qHSL34f8KO7xhnjqEZ7pqoB2vO2bIMABfjCJx3jkVN3jhToVvW09UX
xXjMAomwzU4u7yd6mZA8vVNuCOoIkR+uQ57sHVhl/Au+3A27UsZX7cn4zbYKT9DH
TP8Cpub8OVIZ1xChZ+bKiK/6tUZM4CWiAKrnVfhPUJGu4f4y8dM6J6tktGaE9e62
B21nIUnjXZzzL1xQA3Ye36W/8vI0ZalCZvdc1AJLyBqvgMt5gHo82IcZ4U+bgkzF
k5YJ0zwgQy831ps3fHZ0j0Y+WqGlKF+1xtSuZxzKaXvB48FyBKxifzTpL4+zsZz0
BtXQWG7Jza+ROimdmUIuOG8irYMiqjfxElHbnyzrO+wQcRzaf1kma2TbeDKfqMRr
qb0J509Vurjsu2SvDXW24YRnCcHCCHrvT2PfshvcxG+5y8cs7tAsL11cZaFk0y+8
9PGib1yIt+0nG+4ZwoC0jlEJmXfQFz0KY5ERTmQ5NJFsn7fCO4qea5gGhOM50EBT
HxEfN+5dKC7kKNce4ZXi2Lvn2K17o429A2csCbWRVNawqP0ctKjyGEEbRJms3IB4
iEGnOJdi5hhuJnUXH/TQmSfOBtIBdEO9X6B5bIEsw2/NCK6SjsTwl9gCrvYlW1ai
V6rriDr+v+Ca1j3yriehCUYOsPH6XZ7sVYx1sD2eFnr+6qhFvF00NmDg9xYGaJ7h
AwQS5oW/FmPBZtn0iJ07/Jey4u9UJiGX1sCAtftQis9wY3EDuC8/1uTpFf0a4aeN
D5bsYLsRn/s4qPrU3jthV9Mv3/Y1Qwkg5HO7+m0Gs5fpv7VO/pMD6i0wkAVMfXZJ
KTLGmAmtB0rxLvnewLuM65YXE26RwtWBTygoyfAUZeXnp58Z+WGXHe/GeO2Xk9/e
25E6/chsQJuhojNpZkfNC6SZ3pyXUETIK9sP88SZfQPkfhfCO5UbUpWY8Xbizgu7
jZSuk9ZDpJehcRoGUgYDqHwLwUdIJzlyJWqrKSe2JlVLUoQI+/nTxfcnOwmIdeVH
RGeJb9RjbLw/3bEzc1aMYfjTbjTpv2b0V+0z7f27tgTDU1DpHv5eflcswbUFI8bO
5uCwn/CkyiIcu4NgLxyTO9rZcD4/LoS+JuaokfuATLcYxQDKMZcmwZZyIO33dkRt
+rV0rl8nra/7OQ0wtC/aGd/5nnVDkNZ48Ikvum4w7jrudtQwFlQJHWTaRQ0xcEF4
B+PtC6lHWmICgejfQzZYDJ8XzKqT2lAYs3zgNaciue0fNE1u4QJgcktGgmmJehBI
u+/obr4l4IunqXMtZIWVJLH/xF0DvhzG7uW1oN2h8dTCtP1+UQAF2zV30e4nLVVw
abnOBeOLM+Vh4BIgYn/p/FwCX7usm/liT/aXBYV6mTF8T7tkCkdKoRwgccNwTvX6
/gNJrPx0tJDNvnTKVqHhexQNKfqvE2Iyrr3noll4O2dqWt6WaoW7+FcZIzOyXnBo
bcgzw1wRHrI5ughw56IC9J24JmUYzfrc7CXT/R2mMDi1NUdUOD5WXmGjma7JV9dC
JVCAqGUzc1u9pQZ11OAsjCHHf1vf+R4WNmCW4bV8p6ANxInDJZB+RmWEYCu/QFS/
dMPvNBP8+NufjXVfAl8PZ5bUZGk0bOin/WBtcQrSkgHWWALQdeTPVGZbh+I2zE+Z
zuVmGbom43/rBfZj9+uACVFMwvgWb/Dtxym8qv7rmCG0YPtTiPOzCOXIskc37iDq
I1OHMV8jyEbhCitUt9tIiJ7pFVsp/bH5pYF39m6KMX8vJtkI7gUuHParcNJb5rXK
D8sUQHD5i5Sw8oiF0vpEWM97truoHwwZrGWTEJzHN9EyS/uCSdoaOsWXwJHdknIl
6BsHVZ9l2ybOT1M3YEkQkftBbty7W1jsCw8fbVXvjHMM4IPGYYhJzF5u23UDxam6
FR9ZpZ6OUaH6RfUfJJxkffCHMyE60BZMTH2KPswIPaEywpfGFAo2lrsG2M5kwudL
MdszKxA16hPZuTU5kDluvFtTwebG19k8SeF7WFPQfffKfr8i/XTzsKmhEdLAbsEF
Ln2NUzfzNw2SJgHq2pAgtJPuIZmPyzlHArPbFulqmkR2DxnGqfrhfEUTeMN4lTST
YlOPTrwNkI7RjC96+5W4mOBJh9LXDtb+giF+4m8r82ZLkqaN2RTpmTPWQxJvLRHO
Qqs56yhn4c8Y0IMBbEWCzdfmvHlTLz8VDNmCg1YGsajXsDvAwwrjY/vx7Fe0K4Dg
J1b1mMcdYTDiRU+5nLJnipwRdOYhDh6JQiT8NUm8cgbj039bhhD+a9IumtVDzzeD
FLYudb9ump+Ym5WeaCv4CjwbMzN5pEl6juIZh9AIxe0CJzHwL1ClPwyX5bX0yhq2
Ion5swTeNScZRh2PN5DjlnVbON+6pSHyz0+fTg0sXlAPhOJhIR2eE3WBV9hLR2W6
YJTFDCdCaeaMwS8i/oRxia70t4GnUEVIyemmv5R8fIzt/Ki9IhMhhq7mvoUGa2cn
Gy9hk8TACfU/5Qi1XZ/ZjXb1/yo7/dDnZU2xkhK/9hrTBBigvf5bJdM4e5TExb9u
IenSGOfxPwKxywMZuX/aOO+VZJYRKhDeiusyDCiGD4GRgW2jzeIUCI9rhUW6YOUO
PFN6elWXESreRZNQN2uyB85SthQF6MTjUouZv2Udlf483wV/o7eduV4c3cc/dZ7J
lZlIHxS0AVkTQ8C5HEip96xfYKeeKrnQyJ5yf66ZbiRa3ecaDKU7tt9vCEhjDtHD
D434Ip5G1s8LF05NU24cw6tueVN4AoLAFkBDgpOd+7Itpline9M60YNlqaDwEsvp
Ze6PlS8iK8+Dopd2dgn3eMXdOyul3q8vO7IUAmBr/7e3sktaOdHipuHlQvQIv28v
GDUhAyJ/bI3d8+e2IM+etiatYdYGn7H052s0MQmfBqScrCPfS+MVj3GDMfUVqFQX
UGmJM6+6wph8wdbnJmA0zQsrqVnjaMoXIKfet/itQxCr12OZUjUb/D5SLMqy3Z7b
BR4bf6EBtzwypDB4jMjYsf1+rDu9K1VIn5v1jf75ix6xnKTtLxpIJXy1KGHA9mo4
RtGVcaf0rrz7kXwmuloojKMhtSkEKFSBv59AWiMIFRfnh0brcyzZJeCXIuiEbN3o
EGkhNj0cVpbjlX5a0zusHhftU3fVObPlebNyCrsOVVy6awRHs0KwFZomy/ulLzzA
Ujv2tCrlbeNkn0ejBTpfnAdGCjIOQYdnachDVxk3E4OfnCayywxx7GswbVnnqn0k
fphpiMVAgWUNKdSWfKRWbhZvr1d+5l/EzXYDxA9dnD76Bm7js/VqlPjRhnZxjI7F
w97Cd6MAbWfEyf6H7SZC42nip1laEhv3VP6LsF7Cn+pD9qa3GXQqkho7sppUxsqo
wLgcHjK3YQk19nSfxGFZ59tvDP96mhrTea8n5x6jbobcWM+fRgLmr5mKLIM5ABHb
Pzl3G0YayKAtc54kQswKZFLUmhMkHfGPSDGiDE4ogtierU3GAykXoPZsHQri3Hdp
XsMCCrV4x0oVvTFWGV/4I6kcRjqNXG2a7iENPCPDypbA3GBDdKjlTv+KpbCGhmqY
OB3tZb+re1SCh0zsKzyPjx/YTRAxXvpGBYVBi/xlUBTN8UrJo9HwVymqMyEJr0ar
S+TbepPPPn3fURQIbc6RM7hJUcLmLD+1tPGL6ZoE3xwncvFdF+7FV8Nr5ExOnBgI
y4Kk9snLpaM0s252Zaz1gFdH60ZQwuuTMUM70CIZS8zY5MxZRcS5lVNLzoMUPxS+
`protect end_protected
