-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
U0TFm2zYo+EIh+q5e3OktaL3cL686o6O4+OuDn8vVOGKg+0GKD02hFBg9hAUsNNTc7hg8fVd1+gF
5YX6eeS8aIAqd/GCd7NwmtedOj7h1yVvFg+cLNzkgZGpHrUJnsdONUaz6iztRdDmqp4HKYJ+o40b
O9uJNiLTsBOXL6yWqx10xp/EsGGZp++Me2bBLkYAnU0tZM9X3e8dVoRtqgYYC20tsPiL0G34qLGu
lu4X+U9uLdRPGBPFK5kD4ajkyrkhQ7c9RymwgSnjsr8bOD6lB4X+GvZz2M5Ezwtf+WC1VfjTjlfh
6VPaivbNX/hBLwJOFQnmwNI8IiIvlix5AnIpqQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4544)
`protect data_block
MuRdLka4zLdqxQqYFg9EI2QmtGY8BLVFn16UNMW/lEK9BqMHN4SXx6JhBnVhMXLk2gS43yTX0e08
Ymb6ZoSYVPMu/a5a+7jLivjD2a0rUhkfuNT0tSHm7g3b4N2d4J+/F8444Y/NHUlOMuRYNaX3AE91
Tx7HniwZNwbcXf4zXgIrO5uxAnIGs8CsOxi8emy+h7rjrmJQZ1JKxuf115TjgSRg0hEozo00CXI0
wyGE/a9BtGcDh0B/UZ1XfBdlGmO3kwG/PBDN+qhd8a3uVvrUgWlYAzWlco1bm7bQcISkTV5EzqKr
VFSHukX44qrAnzn2ca5R+FMwtHxXnSjT5viMM6pNT56bQvYq0J2RO9xdodpJ86RhoqfnC50G0txv
2tXEW0gBDOMkguT00NcAKL3PUJhxexUgdKGQVpu6LSMduXgIMt/DF0UW60jt4PMQ4IR19b0vusPf
QbsPAhowUfFMjHicQOYV58BBchqQcaJeCyVAM8Jcjocwd0rMd1tYJ3P4sfWYGqCTEOZtcYWmVzbr
Vzygr/ohDQkp0Znh0p/G3LMydnE2ON8c6mXjm8o5Rkt/TDWt9LPkWEuJPzblqUJRUAv1ccCTKrvt
OYHy5jMJbyS4TC4tmn35OGQ3jFfXwFcIOmO6dKahukI1PQvLJw/cJcnNOIKXuO7LD/nVc+ak2fpw
/PN8gUe5cZq6pOyOf/7/n234C41MOca7gSKqvoS4VOKQ0bIshEjXnAepFKTk0qa+UvKoJ+4I1QaS
TO7ZAqSMvWXMeUvQiCWnjxXfjWOg24E+lhm1MTQkljRWAJ5+pkaevYUnxmKKWDuHkQlpNS5YsHxt
npQehXKbGOkXpRciep4IpmTemJSEZxQ8w1voT/6IplY342x2kHlH0obopUB1laYQ9BZpvhmF0HP5
fZfW2xIx39AIqVRVfLJN5PT3CI6PrDM2GJKc4P9/oEfRlifVmXWUCArrmVSACNKdE63k97u1y/6c
IaokW0Wqf4WtoPctimRLw0kZhnTYv3MH/DAucPJaR5HfKCJ+1Bsn8z3JL64I+pMlS4Wb4NRpwtgl
vSlWxam1psBuubZGCp/UY2VAahQqkIOF+MY+lsc6Zb61ciVgT7HMFsXm7KE2gTWGX0QDegZPtHyz
Zh2miOTJ09helrUJ69qxxtA+Xs1wdHrJiYwLcfREa70is+84D4qdEpqGOlUe9RWihWWij0IXFv9t
hufYs8fsmn2q8HHK2+MBWi/wtaGIb+P1Ay/vnRJB8jaMcv+f3YsXKw6NyQULamVC8xvG7GIXo2qi
a0DJz1oB3rnB9wWCI9iUIiSKPTVvBJWDfW3QetPcIJQB+sIIUQAgycjFDJCnOB+JD06AXkAVKSmg
dqLbuqeAG6biBX684PgKMbBUccuAoKYQyRdXfx+aAbtyNujApr7qx/3C5DNXCWGuCVRogWDN9/EX
Qz1nVoPXyJHn35a1eqA8kWwK8tRlhE1oSLYcfir3aFilStipLniG5sT5KngD9zqmRh/eqKneMzeW
ndz0ry+AgDZgL7e1HtBF+8BhwRZpVMG3syBlE5Qq7429fQVIIpYGbpGc0uI1KanuR6aG0SNMre6j
I/cUy2jDuLxzYNuv9IMfSKKGtXN18fbb6fJK23BILNcp6QS/rTGOoVqoI1Mo5nHCUYezIquoJyYH
h1TmIvJLuOBghWgGeWqKnvsYKhdoIYOTjNOJAAv7rOFvZpZUisClJYP4eghi3gEaVVVgHpVeCOMP
2CLLLqU357mrevJXc/RhiK4ZBMAuYMhC9+h+R7Vct2i8Ab3V0p5HNcyRcSS8q3EuJxe3f4XwJvtb
MRdS8PNaj4o9POK+qL/VnpUlUrMqZqRGUuW0ZgOtIwW4F+4oF9mzy0/tb8E5v65+awmiQ/96q1vZ
Fxo4WOu5OiDCcT84KKsKa591x3/bLnZwlbc6PvmRxkoo2ayTbNX/Gd1ie3QLssrOzWb6esnjI8H+
jgs1wVXyRxgj4z6EQgUln3LCSGWJF6QE/EBuYAl+wcBP5Soq9g1LmPCaWbnSofv6zG3O5v/dQ070
iBaWQurz++ShbZRfI959k60/dZg6SaJNK/KfkI9Mt953hxiiy2SvQkh7O15SC/mr1Y0dHYsC2ZF4
SNZ6sZynMSD8JXTLWn0O1WVtqh5liAO5nJB/WZWz9zxEnFGDKxBfEhSBMyrP4p2oKx8u3d8qJphr
VsnIkYNbEoBs2cxjV2H6Y4mvcR1lPL9A0tjbp96fK6jUm8r6permDxoIHwqDb4OETtmrMPtKShwd
cZpS5k3XqAQBUSWqPqQClpq3aigo9pwU5eG+Tpq1xUnYvWFgDOKf1iE0gwBY0+FUCc+xzmGCEtZ2
QmxKyuo6m9bSOq9XgcsgaEiuy1LGRgi7qpUN/u3WXlOhzRdAyl9EH2RRwK+8aLRmSHDUB75sRGQo
3oBUEIj+Gmu27ko1yyqKOcAnsKWeNRjUloyjG12m+zeKEocPHiAlskuRCHyq7uuJSwIw3ggzY/Di
lZq7w5DRsUjDAPx/IARAlR7byJKFb11ZThDV7FWeBDXBLfh/dlbWTYb50pMcyOm083R21e5eRXli
WtQatV8YGMyHPbNlNAROPu4v+yW+e52FNHLxfLWEFoKExUxO/nnJ9Yvoe3iKfStNGPuEYp+hXyLv
qvFINmatWPVb3DJ2cNl7tpAaMc0fgE5eTdTd2wke6qWc6CtdzLu+KlNEyYINKKtO39X3mIy4480c
TKMt94v+DravJwDHY89meRHuC3L+zfc0Tb72d7UjS+/urlP8T3vgOKSjK0N6h0z0UhLqcXRcX0fS
hSvtBUCn8mzqB0YSNB26hPfMAb1uBXPxkWajlPHwOU9MU6zpzQ2eIy+e5Z89V9XobvB1KxFpXIgS
ANhFzenh4EJL+xfG+fvRXkGkEXqWGkaSerNq0t9iRouAUjOR2SqdEWAymBrHIFMEtvWrGr34lgMO
VC7DpmGLKXyP9eEnusj/Kx+w7CJjYRFh8FMutBWLKlc8NK1AjP2xzGTNeZ/KjX5xqljLXyPjR/ZC
fmRmem4N/IgjuK6Cr3PRR7ch6TZpdznwPfHlu8rK9s0S2irxRnRaTRIpbOE7xc93LAvjnUgAOFYw
uArIj+dc1qs4eaaO2yECWZDaGbOZl1I4k6VZphbbWSJ7LSmrH7hakPyUZqQJE7v8ImpHGZnxFK1r
W7ME6Y959f5p0L51ujoSO63uD8jpfZ1EpOq8YKrgCkFpNGXh831Dxyene7Vhdq0CyJ/jJbC26P0x
ofeBXQA/3YtO+w5Phpt1ZfxGETepsrjkIhv1BIWwRMq7d5wH8qJxJCJljU3r9UAbMffST4xURCNK
gdVTcnPfPlyWmqg5eZ2sf8p44jwGw1Sp8XSgfCNycO6gVCarpGnBKTp9F69YlVGEPxOLzwpz/xcs
neAXvaOIJZvCpyWO6UoBGqZQFXpfVEZbNtAHfC1RGzjoRJ63NC5GCP0IglLcbaD+58aDybcK7nBr
qSMzDJQbtGXcZMmqJE8u9KnS+Jz3+YP7uL6c2Q4Y5xuh+X08Q5RKKRnWLum+1FfRbBpgogAp8SRl
O3nsH1A0U7pJXTx+EMLSLb7HgLggTpJpF7SGWGCKX4pZ8tpkIzHTawjIxEHVSFeAjVQpRjvvMROR
yCe/dZAp+XMO5Lbq2xSQFGZJ+BlQz+XT+I+FxeasMs2Huc0OWRA93aMhaIHH+/mVvVRsDjQbwZFe
HC9aldE1RCk9DZSSz2cXagZab3qo5U2MoiGjtuFFtuLF5aIT/xKgPSgN4BR3O1Dpb4TGJpkFB2EZ
0s7vjR7RPiqiQNsPN8FgMH4qfye9oKBw8HpS+Y7PjReEIwtRvYRHtO4DiAaZeFCmK33W82GJ0QZt
mEUeWkS24h4VexU7GVkt6IBVnflFMrFrQEKyTODmvg3bNKxwobsOqkEh3xSkuhA4EdR5Wq/VT4q4
9iU7WGR9dHBY/CQmYQPQTvWMlQdYcDrGNKv5qo723W4ccBhMVjpubcnKyujvBzyhfTzN3j8xAvlc
Qb7spjEg7p+mvpKLgqZZFQvGuyeshmqtLdHUFOnhCUWPECCgUTnY9BWz/dnI2kZjPCY2/DAaqcp+
O6g5bsQkYPN5zwH5jFh7DZp3MgAZoo8bG6GARBh/lcEvaMWXqNgED/r5aEdUjNQJokJk4mXLhtcJ
6RtRJKtfgNkylxls9ZVAabjBRZal/hpfJxnBkEMxHtI8lBzFBiqf0f7ytCF9ZmAdWjmfRxXGZYON
DBmz1gTME0crLUFrMTDwrTNlKBV13zYt42T7ihf7jVjevdrOcJpUnl5w3fjtPT3adFz/Oe+IpN0Y
d+lI6f7YuNAjW/fUyhe4MrinvHVkTCqDk/mZBHZYNU7k077BoNDBv0g6FETVI2kfw9ZoO9Fkb38X
SI9K1dUO+q9oYU1uDrP67EQougVWEF9pnkl/CUu71OgajdUnWRYm+b7avEMc1p1zmqrM9wKzdffa
6eEy7bCoVQcu6S74wT9d4zZadPJPNSAFYcEOf0Cplzo6ucTYNoU7/1JF1+7wQyB/lmzCJUQe7oxm
3NGai9Sztw8anwaG77po2YwrcB8jXciSe11nH/YBbbgc2DEt0P9jC8V5s4oT173VfcXUyP37/TL5
i0UDYp1JkxjylWtqRP7tZMkXU3J0B3ysAFXfJmGeuSQBSs5Q2FpNdkRghuGPjPM8ewB6TgGLYheX
5ZEVu0onJRsRc9PfPMCXButEnds3vn1B14PvRv1Akj5l16cZV3ldQ9+Iyt52M2bq35mjuWjkwBy0
nu6TSrZ7cmyXthkqgg2X8MQz73GxEzvfV1hQhL+1Il4MR6F/iQ0Ws/HFhoZInkWunOubGeJlzkLQ
xqn6ebg9N22ySPuCYUVjAyF8610BbP6yUN+2eJnFN6QVkAA616PECo05reUaqTrZR1cO1l+h7FtT
yo9KeDe+JliEMSRgzhUZJ+yBtAKoLkCsOlTfGekW1MEJFeCtatJSX8dAsMFTv8mrT6BYc+UfXXZh
WXwIdZKnuZO8wa39pJk+vE6jpWx0jlSBuG8mXx3Dnc2VlVfPMZwOFZlIjAzbNdh9/QOvTBQ6c5lG
LTh+/mM/Mjx/xRZi4trlMWTKbUCyoOKjcxZF2tF49WMRLlWz/mRRZpBVc2njrfdDmu32Kdgg0bPz
l7hZ2at4QY6Yn4Vyi6DBPpUi6KIg8dfJ98/qq/BAZGY0J1/BjHMArYKweNFXwk3yAcX7VSo4oaMm
SyLI7diFfo5QMHQqGShqlhQy6JTqvYTltEmWCWV92VMBdnLuc5O5ZEPv82m9A6jXjmJJV72jQi3B
pE1jCxKUkzgY5xmQtOWYjuBvuhUI5QNQ9y8ryqxP9D4hna3ebVrCr5LtvuXSrvLfeLSsOGZTcckH
+fCPG5MMoMecV3YkpRIdepMYSojkyIh/UxJhURWh/B1Ho6nrrl4rAqTwWI/HX4LItBYCpDJsGjeO
hINSAtPihh4Vk4a1zlKa1BHIFDtVYjmUTztsjcoiSwKFP8VrlBbOXwgvQ/J8AIhWKPWQmY1rz5/R
Uog/tFKVbmLMiejDgufaOxYTUGrEnBMQllieTu52HaYrWgmVNbfN6u23Q4bXiy7E8xiiSXQ/aamq
dXDnF3UOKzGBeevB9fHVotKJ6hd/XZn5SVQndrVkDzDO78bGENFQNhjKhmJjpycFqsZLfdA7QlMY
C6pI0HDYMKYcLrnl0kuIgNAbM+crbmUiARMzNUd9F/3TuAvAn2Es2pCbwRBDuFwICMfGp092pzzw
Nw0mPZTTYYfybqYEWeUagWmFqIh5h4uzVmJ9Rv53yrA45ZMd2nqPhRg+RoKXmBr4B3DTQKlRX+RB
UFVgnd5aY5LyYXlj2DKgZWxKdVE8bCZTl99PG2Zp07+8YJ73XN9tK/cpNUtxPciTQJW2laH2Yshz
mtMF0kPl75ETNolk1AHkMD4nACkbv0LozX4tjjMW7Wt3bwsezv0yXFfldBfZzYFPPwkfnh6jpjYt
VTz8lEp7AnoPrnb8jBmSLRDoXeq2mlEeOogMHhy8Vv0B8lFfNGoNJEs=
`protect end_protected
