localparam [0:32767][0:2][31:0] P_FORCE = {
  {32'hc48b4428, 32'h43a80f60, 32'h4320680e},
  {32'hc4fa86f6, 32'hc2cb200d, 32'hc43d1f57},
  {32'h44a42e11, 32'h438b376c, 32'h44f8063f},
  {32'h43d16b8a, 32'h447cab02, 32'hc3288819},
  {32'h437e66f0, 32'hc504f6d8, 32'hc384035a},
  {32'hc491abb5, 32'h43eaebfd, 32'h43795204},
  {32'hc3f4874e, 32'hc3c6091f, 32'h438f6623},
  {32'hc39fc4b4, 32'h4510e8c3, 32'hc3b45452},
  {32'h44dfff6b, 32'hc3ca0878, 32'h43145b27},
  {32'hc4ad95d4, 32'h431a2914, 32'h43f7abad},
  {32'h44374305, 32'hc438a29c, 32'hc3b2caa2},
  {32'hc4e462f0, 32'h4393a1b3, 32'hc398ded3},
  {32'hc27b4deb, 32'hc49153bd, 32'h4134197f},
  {32'hc42b3fdf, 32'hc335ae3f, 32'h44c88b0d},
  {32'hc30e26d8, 32'hc4eb4ddd, 32'hc4204e46},
  {32'h44f533ad, 32'hc35931bc, 32'h42aeb745},
  {32'h44e63f14, 32'hc3de9fb5, 32'hc31ba902},
  {32'hc4b88912, 32'h43428afe, 32'h4495f0ce},
  {32'hc48afa78, 32'h42a2d2ad, 32'hc3c9ec8a},
  {32'hc581bc4d, 32'h4314bad7, 32'h42c33a75},
  {32'h44fe3abb, 32'h43f39a99, 32'hc36709e6},
  {32'h44696686, 32'hc2e0e0ef, 32'h443afcc3},
  {32'h4433f04d, 32'hc444bfd3, 32'hc4bbe57e},
  {32'h424caa38, 32'h45091af9, 32'h43c57ace},
  {32'hc4cf29b0, 32'hc196a5eb, 32'hc330d220},
  {32'hc47ee262, 32'h44f70841, 32'h4434a0b2},
  {32'h4334fb6a, 32'hc4979fb5, 32'hc4c7344c},
  {32'h43c91c07, 32'hc300b0b3, 32'hc4bf7d9c},
  {32'hc4932558, 32'h4281fa70, 32'h437360c7},
  {32'hc4a4db04, 32'h42813d6f, 32'hc3a13b43},
  {32'hc4ae1f29, 32'hc4094546, 32'h4386dbbd},
  {32'h4508cc4f, 32'h4408026e, 32'hc3395b7b},
  {32'hc46aad38, 32'hc39fc414, 32'h42d4f1c4},
  {32'h453979f3, 32'h43ff1b82, 32'h432e5953},
  {32'hc520cb08, 32'hc478359f, 32'hc2fc0c28},
  {32'h43e31687, 32'h450bf2f4, 32'h42a38f6f},
  {32'hc447c287, 32'hc3490832, 32'h4480a5df},
  {32'h454b68c5, 32'hc391badc, 32'h41400d78},
  {32'hc4ab67a1, 32'h43252855, 32'h4287213c},
  {32'h43c52197, 32'h45265e1c, 32'h44054eed},
  {32'hc46866df, 32'hc50f32c8, 32'hc3ae6260},
  {32'hc4c29f32, 32'h43dab2c5, 32'h441289c3},
  {32'hc4f13da1, 32'hc32e3185, 32'h43290866},
  {32'h4524ccec, 32'h440a2de6, 32'h438d1260},
  {32'h4374799a, 32'hc4759fbf, 32'h431f9c28},
  {32'h453075d6, 32'h4452c172, 32'h4301a0ff},
  {32'hc51c1737, 32'hc393d06d, 32'hc40ec8b9},
  {32'hc4a5e728, 32'h437bf08e, 32'hc2900fbf},
  {32'hc2fe342f, 32'hc4bf1c23, 32'hc455def7},
  {32'hc3d450a3, 32'h445bec64, 32'h4415b778},
  {32'h439270dc, 32'h42cf0da0, 32'hc488cdb4},
  {32'h4426540a, 32'h44c99ea6, 32'h44824251},
  {32'hc458afd1, 32'hc449f09a, 32'hc5132364},
  {32'h42ea2d08, 32'h44ed0052, 32'h438846fd},
  {32'h45106bc0, 32'hc43ae518, 32'hc2a54a8e},
  {32'hc42d9224, 32'hc4975014, 32'hc41874b3},
  {32'h4496da21, 32'h43fa6cf6, 32'h446a6da5},
  {32'hc4c8b103, 32'hc38b9ba7, 32'h41bf64c8},
  {32'hc33d082e, 32'h455cd9da, 32'hc2af1706},
  {32'hc3e9057f, 32'hc514db02, 32'h43a4b5c8},
  {32'h44749e2d, 32'h4360bcea, 32'hc3fa3323},
  {32'hc5185832, 32'hc47c4920, 32'hc4426660},
  {32'h452c2e4e, 32'h43b5ef73, 32'h43f3158f},
  {32'hc3a3051a, 32'hc3cc108b, 32'hc3f2db41},
  {32'h4353de04, 32'hc3a69931, 32'h446380f9},
  {32'hc3e24701, 32'hc4ad20ec, 32'hc2acb53a},
  {32'h44a0f9d3, 32'h441387e8, 32'hc41f360c},
  {32'hc2d8a712, 32'hc50d664b, 32'h43294818},
  {32'h44a93c19, 32'h443565f6, 32'hc43bf51d},
  {32'h44feb92e, 32'hc20cd7f2, 32'h433ac7ea},
  {32'h42f09e40, 32'h4434f2bc, 32'h43e4331e},
  {32'hc40b98a4, 32'h42f3007a, 32'h43e3723a},
  {32'h4465fa2d, 32'h431b5227, 32'hc4508356},
  {32'hc4cee6c5, 32'hc4e47195, 32'h43cfaf85},
  {32'h40e1c91c, 32'h442d7353, 32'hc488f819},
  {32'h44463ba8, 32'hc4cca2ec, 32'h4102909e},
  {32'h4501754d, 32'h441a74b6, 32'hc4016c53},
  {32'hc4f0c6e7, 32'h433806ae, 32'hc1c02230},
  {32'h43705a91, 32'h44203667, 32'hc30260b2},
  {32'hc50618d9, 32'h428b6fb6, 32'h449ebf22},
  {32'h428c134f, 32'hc3d5a86a, 32'hc5808e0f},
  {32'h44dcae6a, 32'hc45d38c1, 32'hc3cb37b7},
  {32'hc4c92170, 32'h44acdb72, 32'h43cac377},
  {32'h4422f136, 32'h438096d1, 32'h440c79ac},
  {32'hc3b149c0, 32'h44a95bd2, 32'hc3bff582},
  {32'h44f38f4b, 32'hc478169f, 32'hc3baca0b},
  {32'hc3f403d0, 32'h448af173, 32'hc3c4c7c0},
  {32'h45130d10, 32'h432f8a94, 32'hc428d3cd},
  {32'hc588ae02, 32'h43008dff, 32'h4419d416},
  {32'h44361158, 32'hc27033cd, 32'h435530d7},
  {32'hc305e3a2, 32'h4484950e, 32'hc4996e5d},
  {32'h41e14d0e, 32'hc53168cd, 32'hc4199d70},
  {32'h43ce8fa8, 32'h43d431a2, 32'h415db042},
  {32'h436b1a00, 32'hc33c341c, 32'h4528970e},
  {32'hc537a138, 32'h430361ef, 32'hc38d60c8},
  {32'h44b554a6, 32'h4362b89b, 32'h424f675d},
  {32'hc42bc8b0, 32'hc36fcdad, 32'hc3a6215b},
  {32'h43ed0c00, 32'h4400fa52, 32'hc4307c61},
  {32'h43f9a239, 32'hc3cc649c, 32'hc490aa0d},
  {32'h450ba546, 32'hc42d4f6a, 32'hc283bb85},
  {32'h40b8f770, 32'h452abeb0, 32'hc416c15e},
  {32'hc46c7e34, 32'hc40a5f7b, 32'h3fb7c5d9},
  {32'hc3d2c940, 32'h4477eef4, 32'hc4bc1328},
  {32'h435666f0, 32'hc26c4cc1, 32'h44fdb8d0},
  {32'h441a23a9, 32'h43f75e76, 32'h42c1f466},
  {32'h44728393, 32'h43f0668c, 32'h450cce38},
  {32'hc54b26d9, 32'hc329a43b, 32'hc44e780d},
  {32'h450c8298, 32'hc325be2c, 32'hc399456b},
  {32'h43298f11, 32'hc4feb5da, 32'hc5115fb9},
  {32'hc28c4ef5, 32'h4461c4a6, 32'h449340d9},
  {32'hc3962211, 32'h4358b5b6, 32'h4408668a},
  {32'hc429a666, 32'h433307bd, 32'h4356e94e},
  {32'hc2e1a420, 32'hc521a612, 32'h4382f488},
  {32'h42ece2e4, 32'hc34ff6cc, 32'hc5286ac4},
  {32'h4357b09c, 32'hc3406bd7, 32'h43baacfd},
  {32'hc3b9a882, 32'h448a1890, 32'hc4eb9a4a},
  {32'h448d603c, 32'hc4f72d83, 32'h43c712b9},
  {32'h450af122, 32'h43ffda3c, 32'h4441c154},
  {32'hc39a40ea, 32'hc483ed76, 32'hc4270fd0},
  {32'h44a5220c, 32'hc4097a36, 32'h4284a793},
  {32'hc4af4802, 32'h421de168, 32'h41f73b42},
  {32'hc486a276, 32'h43f6edbe, 32'h43d7bb5e},
  {32'h432e17ed, 32'hc4a8f95f, 32'hc420c9a6},
  {32'h441e0a43, 32'h44e12d6e, 32'hc2f46372},
  {32'h43d37a64, 32'hc4ddbc78, 32'hc2b28a7e},
  {32'hc4e8d1b6, 32'h43242fc1, 32'hc43ee75a},
  {32'hc492136c, 32'h43c821bd, 32'h4388646e},
  {32'hc588c288, 32'h43a7f9e0, 32'hc2ed4267},
  {32'h43eb57a0, 32'hc4120781, 32'h44829717},
  {32'h4313f48b, 32'h44c3bd82, 32'h43ec7dd3},
  {32'hc2c18578, 32'hc54aecab, 32'h432ea91c},
  {32'hc490a376, 32'h448e32e3, 32'hc2ae1169},
  {32'h44ef0cbe, 32'hc3a804a0, 32'h4205338a},
  {32'hc390f090, 32'h45877c70, 32'hc3a735a7},
  {32'h44c03890, 32'hc49a4c83, 32'hc347db47},
  {32'hc3c0b6cc, 32'hc494df47, 32'hc2e60688},
  {32'h448e1d17, 32'h4296e6c5, 32'h41d86ea2},
  {32'hc3cc2abe, 32'hc3bd414d, 32'h450f39e5},
  {32'hc48b1dca, 32'hc420470d, 32'h440a6d9c},
  {32'h43dcbd39, 32'h44d9c8c8, 32'hc2338f82},
  {32'hc4a68553, 32'hc2cd4e48, 32'h442ddefc},
  {32'h44599658, 32'h43ae9bda, 32'hc2c4fa55},
  {32'hc4d99e8c, 32'hc313df80, 32'h442f4be8},
  {32'h4366cbaa, 32'h43ea02d4, 32'hc3f9f135},
  {32'h43118004, 32'h442cf8d4, 32'hc3ffba36},
  {32'h431871b3, 32'hc287514b, 32'h44af086e},
  {32'h44169846, 32'hc4845d1a, 32'hc485d49a},
  {32'h43930ea5, 32'h43f816fe, 32'hc422c3d8},
  {32'hc400df21, 32'hc4cd30b1, 32'h444c0916},
  {32'h4505fef3, 32'h41eee0aa, 32'h4398c7d1},
  {32'hc4941c9e, 32'hc48e5dba, 32'h43d6f0b9},
  {32'h443fc217, 32'h42aeacbf, 32'hc4f5a221},
  {32'h443c7d25, 32'hc3a03bd4, 32'h44af518e},
  {32'h455331f2, 32'h425e3a70, 32'hc35370a9},
  {32'hc4ba8dd8, 32'hc2e0c63e, 32'h427d8132},
  {32'hc3ec9b9b, 32'hc239d08f, 32'hc31995ad},
  {32'hc5234170, 32'hc422b426, 32'h43873897},
  {32'h454ae81d, 32'hc374ad06, 32'hc1f15358},
  {32'hc52d1339, 32'h42f21a67, 32'h43a36327},
  {32'hc467e332, 32'h45510d50, 32'h43314ec2},
  {32'hc41061fb, 32'hc4a5fc6a, 32'h43d72e8c},
  {32'h44013129, 32'h44bde1d8, 32'h43825485},
  {32'hc3d34cf2, 32'h431d4062, 32'h4386a97e},
  {32'hc39c3edd, 32'h42efe02c, 32'hc499512c},
  {32'hc3bf0a43, 32'hc4626307, 32'h4502ee6a},
  {32'hc4fcf15a, 32'h42237ba9, 32'h3f87b9a0},
  {32'hc2e43143, 32'h425dc11f, 32'h44dcdf97},
  {32'h42d38890, 32'hc5264137, 32'hc38eadcd},
  {32'h438ca567, 32'h440353a2, 32'hc16ea3fe},
  {32'hc2ce3270, 32'hc4d351ae, 32'hc4df90cc},
  {32'h434b63fe, 32'h4444a677, 32'h4512d72b},
  {32'h427cc271, 32'h44b1859c, 32'hc3d7048a},
  {32'h430d7756, 32'h4433f9a4, 32'h4480c4ba},
  {32'hc3de0c3c, 32'hc38a5154, 32'hc4ab122a},
  {32'h44f97003, 32'h435963ac, 32'h431b0d6a},
  {32'hc4493406, 32'hc39c30ed, 32'hc3d55185},
  {32'h4209fcdc, 32'h43e75e2b, 32'h44a04e74},
  {32'h42780d84, 32'hc34a5e98, 32'hc50c2d28},
  {32'hc3bab78e, 32'h44b54b49, 32'h451f132c},
  {32'hc4431ae9, 32'hc4adbadb, 32'hc5021a0a},
  {32'h426e5b7c, 32'h3fb30056, 32'h442df89e},
  {32'hc39d7680, 32'hc5294c16, 32'hc44f5979},
  {32'h4549343a, 32'h447ff209, 32'hc10da8d0},
  {32'h411eb628, 32'hc46849f6, 32'h41f8ca94},
  {32'h4507bde2, 32'h43cbf1e2, 32'hc3ba0d84},
  {32'hc5349802, 32'hc3f6839d, 32'hc15335bf},
  {32'h455839e4, 32'h435b3d69, 32'h43a5eccf},
  {32'hc4534001, 32'hc35b65b5, 32'hc1663c2e},
  {32'h456c5613, 32'hc399399f, 32'h43617b70},
  {32'h43d4fc76, 32'hc4232b7c, 32'hc43b8b3f},
  {32'hc39a5955, 32'h43497546, 32'h442ca56c},
  {32'h450788e3, 32'h441395d9, 32'hc3962014},
  {32'hc4a17107, 32'h43a7d38c, 32'h44563196},
  {32'h4439ffdc, 32'hc49051b2, 32'hc49fe9b8},
  {32'hc4474d1d, 32'h4432f339, 32'h43b19838},
  {32'hc38aed70, 32'hc46ac717, 32'hc5108543},
  {32'hc53610d6, 32'h43af7444, 32'h445599b6},
  {32'h42a436d0, 32'h43e9fc2c, 32'hc4c7a1eb},
  {32'hc48c3d71, 32'hc30408e2, 32'h448d4f9e},
  {32'h4440e38c, 32'h4367f88e, 32'hc409ab6f},
  {32'hc336cabe, 32'hc326ac70, 32'h44ca58c6},
  {32'h43903dcd, 32'h431aa745, 32'hc4b2ef67},
  {32'hc52a9a15, 32'h42fb3650, 32'h43d0c224},
  {32'hc4bb91a7, 32'h43864b39, 32'hc381276f},
  {32'hc4d84d68, 32'h4468771c, 32'h44047d11},
  {32'h43d972f8, 32'hc358b28d, 32'hc497e984},
  {32'h436ecbea, 32'h440d6304, 32'h4436c673},
  {32'h4429ece0, 32'hc4c4e2e3, 32'hc3b83f79},
  {32'hc4a4cf9b, 32'h44c22003, 32'hc3518b7b},
  {32'hc4a08a42, 32'h439e4da7, 32'h4225e55b},
  {32'hc33c7dba, 32'h44bb654e, 32'hc4081ac9},
  {32'h44db6625, 32'hc45c5319, 32'h43380ed3},
  {32'hc47e0165, 32'h444925c3, 32'h422e0608},
  {32'h44e9a5ce, 32'h43dfd9c0, 32'hc343006b},
  {32'hc593bc42, 32'h434b2d41, 32'h4282bcb2},
  {32'hc506ed8e, 32'h437a4174, 32'h42b2ae38},
  {32'h44711a3f, 32'h4192bc51, 32'h44e147f4},
  {32'hc4c6b311, 32'h428884ca, 32'hc46f902d},
  {32'h44560c50, 32'hc42a9a59, 32'h43abc1ca},
  {32'h437b3534, 32'h4395614c, 32'h42fd833f},
  {32'h4508fb60, 32'hc3abe48b, 32'h4339fe7e},
  {32'hc4c53f87, 32'h412bff08, 32'hc2ec28af},
  {32'h44a3da51, 32'hc2bdab72, 32'hc2b811bc},
  {32'hc49be189, 32'h44beeb85, 32'hc3c78e45},
  {32'h440f58cc, 32'hc510a6ca, 32'hc3788ff4},
  {32'h43800f99, 32'h441ebb2d, 32'hc2914035},
  {32'h4357abf0, 32'h438d9094, 32'h44eda34e},
  {32'hc50769e2, 32'h444376af, 32'h4306c15e},
  {32'h42918b34, 32'hc418a344, 32'hc3b501eb},
  {32'hc4a64960, 32'h42839639, 32'h4408fd88},
  {32'h448dbda6, 32'hc40ff336, 32'hc3fb8b26},
  {32'hc478d7a8, 32'h43403970, 32'h43cc8e0f},
  {32'hc2c13e70, 32'h436c6491, 32'hc4eed2ca},
  {32'hc50e2c2d, 32'hc126a3bc, 32'h40a9de8a},
  {32'h44825c26, 32'h42d02c88, 32'hc409b958},
  {32'hc511c3e4, 32'hc24b000f, 32'h43adc5d8},
  {32'h440f71c8, 32'h43d0ac4a, 32'hc49500cc},
  {32'h44342ca2, 32'h44a1d77f, 32'h4299a402},
  {32'h44815b25, 32'hc444f8b8, 32'hc43cceb4},
  {32'hc30d1be7, 32'h4481b188, 32'h44838de5},
  {32'h442e2dce, 32'h43a6d2ae, 32'hc3a846e9},
  {32'hc42681a0, 32'h448bbf5f, 32'h43c571bd},
  {32'hc1aaa508, 32'hc480868d, 32'hc3d77600},
  {32'hc250ef88, 32'h4490e03e, 32'hc5076594},
  {32'hc53479a1, 32'hc348ec86, 32'h43576d99},
  {32'h44cb9c40, 32'h43e9d802, 32'hc231b2fe},
  {32'hc3d4698e, 32'hc543a79b, 32'h42a5f79a},
  {32'h4409f01c, 32'h44c93f0c, 32'h43e3b6c5},
  {32'hc50aae5f, 32'hc2686f77, 32'hbedbe83c},
  {32'h43c4df5a, 32'h44ed1cda, 32'h41da6081},
  {32'hc3901ec6, 32'hc4af4575, 32'h43ac8aa2},
  {32'h4525633b, 32'hc44ca047, 32'h4392aaa4},
  {32'hc50f8c58, 32'h4318fc06, 32'hc42c0c23},
  {32'h445c62b8, 32'h44141a95, 32'hc3bffaf2},
  {32'h4493cb27, 32'hc282488e, 32'h439907e0},
  {32'h42df7947, 32'h44dcfa76, 32'h443aaa71},
  {32'hc422be76, 32'hc456bbfd, 32'hc527bb85},
  {32'h43fcc269, 32'h445e6812, 32'h42cc244a},
  {32'hc2ed5ce9, 32'hc46e9898, 32'hc4477f8e},
  {32'h433f3232, 32'h43a8ddc9, 32'h4540f95f},
  {32'hc3bf7374, 32'hc43a6932, 32'hc3ba4bc4},
  {32'h43ba0c8d, 32'hc40e16ab, 32'h44883456},
  {32'hc4e27a03, 32'h4352d6f2, 32'hc33bf5ca},
  {32'hc4142ddc, 32'h440879cb, 32'h4358c4bf},
  {32'hc4a86d8d, 32'h42056c7f, 32'hc48e47a5},
  {32'h44711557, 32'h44c2b233, 32'h43b91642},
  {32'h438084e0, 32'h432f914d, 32'hc4bdb4ec},
  {32'h45627b0c, 32'h4333fd12, 32'h44180375},
  {32'hc525ae0e, 32'hc35c6da8, 32'h420a1d0d},
  {32'hc271caeb, 32'h450dc179, 32'hc347cd21},
  {32'h4416e7ba, 32'h4424d113, 32'h43d8bbd5},
  {32'h41d32a1b, 32'hc570cb77, 32'h43587a38},
  {32'hc2a6cb58, 32'h453439bb, 32'h43958635},
  {32'h44a0fb4b, 32'hc3112ef0, 32'h43da3c9e},
  {32'h438bb9d8, 32'h44200ec5, 32'h42f518ac},
  {32'h432f90c7, 32'hc55a5283, 32'hc1eb417d},
  {32'hc44faa9c, 32'hc28713ec, 32'h43f21f9a},
  {32'hc577dbd7, 32'hc3c428e7, 32'h42b551d1},
  {32'h44b9add2, 32'h42dba33d, 32'h4437f809},
  {32'hc4ae023b, 32'h41e41c79, 32'h4387840b},
  {32'h4462af13, 32'h4406912f, 32'hc3fa547c},
  {32'hc3be4d6a, 32'hc4183f93, 32'h446d9d69},
  {32'hc395a966, 32'h42d1c8e4, 32'hc37fbde7},
  {32'hc416b4e2, 32'hc505f61f, 32'h44294963},
  {32'h44879c34, 32'h428db147, 32'hc4211a11},
  {32'hc3b9cc42, 32'h41f0f794, 32'h4466b166},
  {32'hc3c0ca0f, 32'hc331459b, 32'hc55d5203},
  {32'hc4ac9a74, 32'h43b13bf4, 32'hc2929f13},
  {32'h446c1c00, 32'h445bbc25, 32'hc424f050},
  {32'hc43211e7, 32'hc5351fbd, 32'h43eda60b},
  {32'h4527a56d, 32'h43acb721, 32'hc4811669},
  {32'h4420f5d1, 32'hc206a7d2, 32'h4361a224},
  {32'h43e46592, 32'h4534a06d, 32'h41e9f83c},
  {32'hc3220fe0, 32'hc507fcce, 32'h42fabe67},
  {32'h45502a5a, 32'h4308e1b5, 32'hc2d65b7b},
  {32'hc4c6da7f, 32'h43333b45, 32'h43ccfb33},
  {32'h4548d9fa, 32'h43990c9a, 32'hc39f31c4},
  {32'h451a5bd7, 32'hc4473edd, 32'hc3cafc64},
  {32'hc43a78f0, 32'h43a628d1, 32'h447d63e0},
  {32'h451ea47c, 32'h43991e0b, 32'h439e37de},
  {32'hc4912f94, 32'h447fad19, 32'hc3e67064},
  {32'h42886244, 32'hc53378db, 32'hc3a402a2},
  {32'hc2da6755, 32'h4502459c, 32'h435e23c3},
  {32'hc2f9a040, 32'h440b7e44, 32'hc34766fb},
  {32'hc4ac91aa, 32'h4443e41f, 32'h4485cda0},
  {32'h444387c1, 32'hc3b68608, 32'h43a024ce},
  {32'hc52ecf98, 32'h43d20510, 32'h4430c08c},
  {32'h438e96cc, 32'hc4334de6, 32'hc3a46ed3},
  {32'h43b6432c, 32'h44817eec, 32'hc2c71bbf},
  {32'h42bc1030, 32'h437ee295, 32'h454fa4a4},
  {32'h422060fd, 32'hc379e6b4, 32'hc4ff2667},
  {32'h43616a2c, 32'hc2c713ef, 32'h446029c3},
  {32'hc4eab105, 32'h4282a6cf, 32'hc417999a},
  {32'h448fd5c1, 32'h417f0af8, 32'h43ee7255},
  {32'hc2ed42f4, 32'hc36cecf0, 32'hc499b05b},
  {32'h441ffc99, 32'hc51d7669, 32'h4317d869},
  {32'hc41c93b6, 32'h44d100fc, 32'hc46ecfe2},
  {32'h44ba79cc, 32'hc3ce1522, 32'h440ba9d6},
  {32'hc3ac6547, 32'h4526a124, 32'hc3f6ee08},
  {32'h44a31186, 32'h429736c6, 32'h448f82d7},
  {32'hc346d7ee, 32'h446cb574, 32'h4401124a},
  {32'h444d9e15, 32'h439ebd8e, 32'h44b91044},
  {32'hc50507f0, 32'h4425b02b, 32'hc4779e59},
  {32'hc41a94a6, 32'h43137090, 32'h43834286},
  {32'hc467e56b, 32'h43937061, 32'hc4771b9d},
  {32'hc467b81d, 32'h42ce2308, 32'h4494043a},
  {32'hc3c2f3f8, 32'h43cc6314, 32'hc32c389e},
  {32'h43caebee, 32'h44597879, 32'hc3565f22},
  {32'h44573014, 32'hc32e2adf, 32'hc3508ae5},
  {32'hc32a310c, 32'hc2758f6f, 32'hc550d976},
  {32'h442c13da, 32'hc3589919, 32'hc2c5e67f},
  {32'h42d4e619, 32'h44ddc238, 32'hc4b7f3ff},
  {32'h448f80da, 32'hc4913897, 32'h4353bc6a},
  {32'h42c3607e, 32'hc4d1fee7, 32'h45298235},
  {32'h43b3a1bc, 32'h431b49f4, 32'hc4e4bcfe},
  {32'hc4288273, 32'h441bd180, 32'h438aa40c},
  {32'hc49b343f, 32'h439db313, 32'h441ad00c},
  {32'hc35583f0, 32'h448929ca, 32'hc460aa9d},
  {32'h4330c518, 32'hc541a912, 32'hc3a00c02},
  {32'h44e1cd71, 32'h40e297dc, 32'h4377a7e4},
  {32'h44011b3d, 32'h43e5da1b, 32'h45549133},
  {32'hc2e4d6e0, 32'h4482348f, 32'hc4309abc},
  {32'h44031d06, 32'h44298599, 32'h42ea728b},
  {32'hc55b8270, 32'h434277c5, 32'h4366d65f},
  {32'h44730b2e, 32'h43d05853, 32'h43b42357},
  {32'hc4c31246, 32'hc2def44d, 32'hc382f34c},
  {32'h44b1337d, 32'hc470c9ff, 32'hc3cef5c2},
  {32'hc3d8d300, 32'h454c24b2, 32'hc328a267},
  {32'h43a3ca40, 32'hc4f34f63, 32'h4282259b},
  {32'hc3fc705b, 32'h44c68ad9, 32'hc4354abf},
  {32'hc2b96488, 32'hc4c41a7c, 32'h4390d90d},
  {32'h443e4896, 32'hc4a3947b, 32'h44571297},
  {32'h44afa00c, 32'hc3ec2d88, 32'hc3960b4f},
  {32'h4210aa20, 32'hc44f4f32, 32'h442349ba},
  {32'hc39d03f0, 32'hc45a14fc, 32'h43c09e32},
  {32'hc3b2511f, 32'h42c442b4, 32'hc51f9645},
  {32'hc43ac14c, 32'hc3e2a6b5, 32'h42bc0ce3},
  {32'h42c22988, 32'h454e4d35, 32'h425d040c},
  {32'hc431cb89, 32'hc515457c, 32'h4312f3dd},
  {32'hc42619a9, 32'h440fb0f3, 32'h4357edea},
  {32'hc402f0ea, 32'h417bd2ed, 32'h4220436e},
  {32'hc3a58450, 32'h43b64309, 32'h44e374bd},
  {32'h44e66814, 32'h4471c396, 32'hc49d3a14},
  {32'hc080ae2c, 32'hc3bb48a0, 32'hc532ef64},
  {32'hc3e87ea7, 32'hc4e6fad0, 32'hc39b8413},
  {32'hc3f1c741, 32'hc3a329dc, 32'hc3c80616},
  {32'hc4a006da, 32'hc462afdb, 32'h44406e2b},
  {32'h437bf5d4, 32'h44168f3c, 32'hc4a8228a},
  {32'hc3727313, 32'hc4a4b9a5, 32'hc215d0d6},
  {32'h45239c27, 32'hc417ae2d, 32'hc1c50775},
  {32'hc5945f55, 32'hc31f4d64, 32'hc3caacfa},
  {32'h441aee50, 32'hbfe8b308, 32'hc235735d},
  {32'hc3bec876, 32'hc5166b70, 32'h4343fa7d},
  {32'h4411d220, 32'h45269e4d, 32'h431a1cfb},
  {32'h44e6c926, 32'h41c167c4, 32'h434f2bde},
  {32'h44df932e, 32'h44306b0a, 32'h438c8c3a},
  {32'hc4766ef3, 32'hc4871d36, 32'h4302d3f3},
  {32'hc3b45439, 32'h4197ac5f, 32'hc413b2a4},
  {32'h4380f70c, 32'h44a4028f, 32'hc3c0b8cf},
  {32'hc482d1a4, 32'h44a883c0, 32'hc456fad6},
  {32'hc26f5580, 32'hc4f74ab8, 32'h450f599d},
  {32'h42410398, 32'hc2c2f5ae, 32'hc4424357},
  {32'h447a4ab3, 32'h444bf70f, 32'h449f0368},
  {32'hc51ec574, 32'h445bd0e7, 32'hc3e31ee9},
  {32'h4504a1b4, 32'h43b580e4, 32'hc22bf9d1},
  {32'hc4d88153, 32'hc3eb58a5, 32'hc4b15f86},
  {32'h448aa61c, 32'h43b8cdb5, 32'h449c2c93},
  {32'h42e43150, 32'h44406b34, 32'h42cbcc39},
  {32'h441a9090, 32'hc2a3940c, 32'h442257dc},
  {32'hc30bcf61, 32'h439334b7, 32'hc503c9a5},
  {32'hc3af1105, 32'h42742e0b, 32'h44b55d7b},
  {32'hc4f8aaca, 32'hc281c017, 32'hc42daab5},
  {32'h44415ce0, 32'h4381f49d, 32'h44b7647e},
  {32'h4399eca7, 32'hc3f541f5, 32'hc4e591a5},
  {32'hc38afba3, 32'h44ca55dd, 32'h44fdbc63},
  {32'hc3a76e28, 32'hc31b13bb, 32'hc4472583},
  {32'h44b33e93, 32'h431c0e01, 32'h43cccd8a},
  {32'hc532a2bf, 32'hc29c7f63, 32'h43a526f6},
  {32'h450230ad, 32'h446746c2, 32'hc2ee273d},
  {32'hc482db98, 32'hc39ad33e, 32'hc39aafd6},
  {32'h44d4075c, 32'h43a518b4, 32'hc3245f34},
  {32'hc42163c6, 32'hc489ea3c, 32'hc3448364},
  {32'hc4c23ddc, 32'h42cc743e, 32'hc3df008d},
  {32'hc452b49b, 32'hc392d1ca, 32'h4312adf0},
  {32'h4546b4f0, 32'hc106b5bc, 32'h43373d7b},
  {32'h409ced40, 32'hc4e1b569, 32'hc412dcf1},
  {32'h42253a70, 32'h4267a116, 32'h448b1969},
  {32'hc29881c0, 32'hc34880d6, 32'hc3e930d0},
  {32'h4405a26e, 32'h44a04403, 32'h44e81008},
  {32'h42d8d438, 32'hc4c6e401, 32'hc476afb9},
  {32'h4476f8d5, 32'h442d43d0, 32'h442b424a},
  {32'hc3a5c899, 32'h4297b02e, 32'hc4f241d6},
  {32'h436892f0, 32'h44cbf0ed, 32'h4511e46c},
  {32'h44446170, 32'hc491fb49, 32'hc3017076},
  {32'h434ec0c0, 32'hc4ae1218, 32'h45036964},
  {32'h43dd8758, 32'hc4c1bdb1, 32'hc43586c7},
  {32'h40033bd6, 32'hc4c17e93, 32'h449b79f8},
  {32'h45151fdb, 32'hc1d0ec1c, 32'hc32227ce},
  {32'hc468b7ec, 32'h44254865, 32'h44484b18},
  {32'h441fb01c, 32'hc420fa6c, 32'hc377dd9c},
  {32'hc3ada765, 32'h43e066e8, 32'h44e5d060},
  {32'h42bf43fc, 32'hc42ebf30, 32'hc4f7ee0f},
  {32'h4406bd92, 32'h434d9afe, 32'h44ebbb01},
  {32'h443324a1, 32'hc4835788, 32'h4283591c},
  {32'hc42ac0db, 32'h452b2a34, 32'h433ab760},
  {32'h454ec224, 32'h4429a272, 32'hc3b9ff0d},
  {32'hc50cdf73, 32'h442ab899, 32'hc2b1dd9b},
  {32'h4475a0c4, 32'hc5253f28, 32'h44009940},
  {32'hc41d9fac, 32'h443891aa, 32'h43586104},
  {32'h4419a803, 32'hc390c32c, 32'hc39c631a},
  {32'hc54920e2, 32'hc3dbf385, 32'hc3ccc7dc},
  {32'hc441c2e9, 32'h42c6f76d, 32'hc3c2e4bd},
  {32'h4526cddb, 32'hc3dbc77d, 32'hc36b493c},
  {32'hc41392b6, 32'h42e870d9, 32'hc3e5717f},
  {32'h441385dc, 32'h441083e9, 32'h43c41dfb},
  {32'h44583d62, 32'h43702df7, 32'hc3644300},
  {32'h44051488, 32'hc4a58faa, 32'h430fa642},
  {32'hc50f2a91, 32'h43e78871, 32'h42d7c413},
  {32'hc4da9d7b, 32'hc3e252fc, 32'h434073cf},
  {32'hc528360d, 32'h445cc0f0, 32'h439a25b8},
  {32'h44c579d3, 32'hc4c329d3, 32'hc1fe8330},
  {32'hc5022392, 32'h42db4395, 32'hc4100b9d},
  {32'h4430e151, 32'h44286ddf, 32'hc4819cce},
  {32'hc48127cc, 32'hc227f20a, 32'hc4670b75},
  {32'hc41f1eb9, 32'hc369cd5c, 32'hc3a35c55},
  {32'hc24ee132, 32'h444f5a79, 32'h44f7d738},
  {32'hc395055e, 32'hc4bf8c84, 32'hc4def9cd},
  {32'h43546bdc, 32'h44be854a, 32'h43cd833a},
  {32'hc42e8cfa, 32'hc33a7994, 32'hc500cf41},
  {32'hc45ac85c, 32'h4418f9a0, 32'h43f4c53b},
  {32'hc470b27a, 32'hc404cd66, 32'h420d64de},
  {32'hc536348c, 32'hc37b03bc, 32'h4342bb35},
  {32'h40311a90, 32'hc2e42522, 32'hc483bae8},
  {32'h44d18721, 32'hc282d6ad, 32'h42a474c6},
  {32'h43bd60b0, 32'hc45fcc21, 32'hc4db5830},
  {32'hc4b531d5, 32'hc2af3343, 32'h44d96cdf},
  {32'h43493d66, 32'hc3c86814, 32'hc404d9c4},
  {32'hc3eb43c4, 32'h44d97770, 32'h447434f9},
  {32'h432bde98, 32'hc493c3f9, 32'hc4a92983},
  {32'h4491a64a, 32'hc26ec7a3, 32'hc50d3b3a},
  {32'hc4d94f02, 32'h3e85a2c0, 32'h42e0d6f8},
  {32'h452019c5, 32'h43adb2dc, 32'h43a8dc15},
  {32'hc4c2aefd, 32'hc3d08f63, 32'hc48281d0},
  {32'h4480b278, 32'h421f1576, 32'h44269546},
  {32'h440a405d, 32'hc4a27f9a, 32'h423a4e9d},
  {32'h4543f195, 32'h44421fcf, 32'h42c38ed6},
  {32'hc5274189, 32'hc47d645e, 32'hc46708fe},
  {32'hc4cd97c6, 32'h4314ff59, 32'hc14c5ac0},
  {32'hc50ba972, 32'hc1cd3bd4, 32'h438d4408},
  {32'h452cd71e, 32'h42c5144c, 32'hc36aa74e},
  {32'hc4bf7733, 32'h42b04790, 32'hc2e9fb4e},
  {32'h43cb8095, 32'h43cf3bd3, 32'h44cda3b4},
  {32'hc5107198, 32'hc401d931, 32'hc40452c3},
  {32'h43079154, 32'h43ecd195, 32'h444e9266},
  {32'hc44a8f9d, 32'hc4b331ce, 32'hc2a7781f},
  {32'h44bba032, 32'h43bd0d0c, 32'hc3799f66},
  {32'h450af5e4, 32'h41bc071d, 32'hc35e99aa},
  {32'h4499587e, 32'h42b68d8c, 32'h43a7cb6a},
  {32'hc40a111c, 32'hc3f1820c, 32'hc4109507},
  {32'h44087e31, 32'h42ac9761, 32'hc34a01a5},
  {32'h3e4d0000, 32'hc407eedd, 32'hc444604b},
  {32'h43896be4, 32'h448ff881, 32'h4424de9b},
  {32'hc4129d56, 32'hc3e69c64, 32'h439942f6},
  {32'hc2247420, 32'h44d37b7f, 32'h447ae08d},
  {32'h40c35a80, 32'hc53409b0, 32'hc38564a5},
  {32'hc44ce79c, 32'h4452c1d2, 32'h4371dc2d},
  {32'hc49b9269, 32'h43fd91fe, 32'hc0d3ddf7},
  {32'hc3ef6866, 32'hc4dd4d01, 32'hc422b736},
  {32'h432c7e92, 32'h4423bab8, 32'h4408eb43},
  {32'h440bd78c, 32'hc3082720, 32'h42ff3797},
  {32'h4493b8de, 32'h448cc7f2, 32'hc1e6d912},
  {32'hc410ecbb, 32'hc3d9b430, 32'hc4324808},
  {32'h442faf6e, 32'hc2a21f48, 32'hc41add8d},
  {32'hc5875385, 32'h42af0c18, 32'h43d33ed6},
  {32'h44c986f5, 32'h44302df0, 32'h4440aa54},
  {32'hc465e4dc, 32'hc4293d87, 32'h43572ad5},
  {32'h43618e6a, 32'h44551504, 32'hc2353025},
  {32'hc442c20e, 32'hc46b4957, 32'hc3bda718},
  {32'h44f581ef, 32'h4329dec1, 32'hc2641764},
  {32'hc3557c0e, 32'hc517b752, 32'h436b83ba},
  {32'h44a5c77b, 32'h44149a11, 32'hc30dbcc1},
  {32'h4499d3a7, 32'hc28df32f, 32'h439de977},
  {32'h4487c490, 32'hc29cc052, 32'hc49c2acc},
  {32'hc447e420, 32'hc406e818, 32'h43026bb6},
  {32'h437d0348, 32'h4445ff71, 32'hc413e8e2},
  {32'hc495401b, 32'hc4ae193a, 32'h452b3526},
  {32'hc2d51459, 32'h44a90931, 32'hc4b39e1f},
  {32'hc3f7c45c, 32'h42d0c014, 32'h43814289},
  {32'h448cb86f, 32'h43999897, 32'hc406a612},
  {32'hc326bf30, 32'h422b0080, 32'h455d2118},
  {32'h44c8a39a, 32'h43c94350, 32'hc20faf74},
  {32'hc58a4c47, 32'h439364ac, 32'h41f12af0},
  {32'h444b8107, 32'hc3672335, 32'hc489da51},
  {32'h431d4610, 32'hc4bdfbdb, 32'h43a42c8b},
  {32'hc4359065, 32'h45335838, 32'h43672a12},
  {32'hc43580d0, 32'hc1b7ff5e, 32'h4409a451},
  {32'hc492645e, 32'h4494629f, 32'hc3418538},
  {32'h44d5070a, 32'hc3d3f552, 32'hc3aa2210},
  {32'h44c1b5d2, 32'hc35e154b, 32'hc39737be},
  {32'h44d6ca38, 32'hc32b8c5e, 32'hc46e39b0},
  {32'hc47c5ce4, 32'hc315172b, 32'h43e1a60f},
  {32'h44c38fbc, 32'hc453ceb2, 32'h4325f9cf},
  {32'hc438c415, 32'h44532dad, 32'hc514a8ba},
  {32'h442f2264, 32'hc1c14d6c, 32'hc3fd8885},
  {32'hc397c811, 32'h4458e477, 32'h423fa076},
  {32'h43d6fe8c, 32'hc35a5df8, 32'h4424a0cd},
  {32'hc42c151a, 32'h44180b8a, 32'hc4603301},
  {32'h44ac8816, 32'hc28702be, 32'h433d3ffc},
  {32'hc4a083fd, 32'h442d6824, 32'h43c1bf8e},
  {32'h444d47c5, 32'h442738fe, 32'h44ec96c4},
  {32'hc38f1f5b, 32'hc36df03b, 32'hc4be14ee},
  {32'h4106ee34, 32'hc4cb34f2, 32'h43937b89},
  {32'hc42308de, 32'h44930cba, 32'hc468d1bd},
  {32'hc4483a8a, 32'h431edc68, 32'hc25d57f4},
  {32'h4173a020, 32'h4441e8cc, 32'hc46ddbde},
  {32'h4420ac98, 32'hc4ac381f, 32'h44a934b0},
  {32'hc425d666, 32'hc3720902, 32'hc4513c09},
  {32'h436f9094, 32'h4389a2ad, 32'h451f8c1d},
  {32'hc486dac2, 32'hc2814098, 32'hc517eb20},
  {32'h440b0c19, 32'h42d7b828, 32'h44261814},
  {32'h43719a0d, 32'h44db2d82, 32'hc471da5a},
  {32'hc2aeba65, 32'h44de4b3b, 32'h44e6cd51},
  {32'h42b5ccd9, 32'h4482dad4, 32'hc4aa573a},
  {32'h43f9ee80, 32'h44b1ef22, 32'hc37d3f6a},
  {32'h446d7788, 32'hc4d8a0e8, 32'hc2afb6f9},
  {32'hc415353c, 32'hc3992182, 32'hc44e50c0},
  {32'hc409365b, 32'hc234c4e3, 32'h438f99bf},
  {32'hc31ad4b1, 32'h45149af9, 32'hc3eff0bd},
  {32'h44db257d, 32'hc39a4918, 32'h4417c18a},
  {32'h4386d575, 32'hc33740b7, 32'h44d61ec8},
  {32'h423f2fb4, 32'h44bf2adf, 32'hc50c5007},
  {32'hc4b2a91e, 32'hc17e7a50, 32'h4404bea0},
  {32'h44f5a2d8, 32'h43bdb750, 32'h431bfac1},
  {32'hc41a3eab, 32'h4500c7ac, 32'hc31203b8},
  {32'h44abd56a, 32'hc27ecd75, 32'hc3c8f5fa},
  {32'h438c708c, 32'h4448b6b2, 32'h43969e68},
  {32'h44908e7a, 32'hc4b1d5b7, 32'hc241f311},
  {32'hc48e6277, 32'h41bf0cf6, 32'hc3e54692},
  {32'hc4f8ca9c, 32'hc3d0596c, 32'h418a2662},
  {32'hc587bb4a, 32'h4389bfb2, 32'hc2cbcaa9},
  {32'h457b1ebf, 32'h4362e5bb, 32'h43807584},
  {32'h44c950fa, 32'h434268ea, 32'hc349c5ba},
  {32'h42cfd640, 32'hc5157a9c, 32'hc324e645},
  {32'hc4f1e9b8, 32'h43dcb8f8, 32'hc298ca92},
  {32'hc41d4470, 32'hc4254d23, 32'hc2778828},
  {32'hc53d0a6e, 32'h43ea2b6b, 32'hc3b283dd},
  {32'h455be682, 32'hc44cec42, 32'hc3972dc6},
  {32'h442714a9, 32'hc46745f9, 32'h43c61b7a},
  {32'h43b73aa7, 32'h4443174f, 32'hc452a55b},
  {32'h4351686b, 32'hc4b1b574, 32'h4505c645},
  {32'hc30aba37, 32'hc52a5835, 32'h43508ce9},
  {32'h43b1812b, 32'h439ad27e, 32'hc3a0b7af},
  {32'h444e73af, 32'h43ac9160, 32'h4391004e},
  {32'h442b910c, 32'h44e60b04, 32'h4215a003},
  {32'hc4ad168b, 32'hc201f437, 32'h448b38b3},
  {32'h451d7013, 32'h43402c7e, 32'h444cec0c},
  {32'h4420224f, 32'hc4297c9e, 32'hc392ba71},
  {32'hc540627b, 32'h429cd040, 32'hc290a2da},
  {32'h44982674, 32'hc4abec14, 32'hc45bbfe0},
  {32'h44272707, 32'h44717c07, 32'hc301ec92},
  {32'hc4df52a9, 32'hc40fb8de, 32'h43141a07},
  {32'h44e2447f, 32'h4350dc12, 32'h4393ba0e},
  {32'hc46706eb, 32'hc4b53aba, 32'h423eb2b6},
  {32'h435967d2, 32'hc417e9d4, 32'hc522dbd3},
  {32'hc42156ec, 32'hc45a8b43, 32'hc2aa812c},
  {32'hc39a433e, 32'hc3bebebe, 32'hc09899b4},
  {32'hc4bfad1c, 32'h433d819f, 32'hc2556593},
  {32'h44c04636, 32'h4010b48b, 32'hc3684a34},
  {32'hc49bc664, 32'hc4cbbf79, 32'h43170082},
  {32'h450c1f55, 32'h42bd7961, 32'h44257b53},
  {32'h439c1680, 32'hc432562e, 32'h43910dc5},
  {32'h421c9d00, 32'h45525fd5, 32'hc368a1c5},
  {32'hc4a27e40, 32'h42a17040, 32'h43199f37},
  {32'h44d62843, 32'hc395b97e, 32'hc407ddfa},
  {32'h43f049bb, 32'hc432cc03, 32'h43b97fbd},
  {32'hc410955f, 32'h4412c01e, 32'hc46111f7},
  {32'h435fd48f, 32'h449f7be0, 32'h445fb139},
  {32'h432caa94, 32'hc495d6c8, 32'h41e67882},
  {32'h455efece, 32'hc39fa08f, 32'h4317439d},
  {32'h42dff99c, 32'h417df046, 32'hc4d1d929},
  {32'h451aba4b, 32'hc368e423, 32'h42bb387c},
  {32'hc55c6a93, 32'hc353a851, 32'hc2b2e361},
  {32'hc387d028, 32'h43ba4965, 32'h44eaaff5},
  {32'h436eb976, 32'h4381ff36, 32'hc4a8f707},
  {32'h44fba3b7, 32'h42ddf26a, 32'h430bbbbf},
  {32'hc352a851, 32'hc4687280, 32'hc489eafa},
  {32'h43a491dc, 32'h44f5e816, 32'h42efbc42},
  {32'hc40125d7, 32'hc4c7c08a, 32'hc03de9cb},
  {32'h4402dfb2, 32'h44c1b435, 32'h448da80f},
  {32'hc45028ba, 32'hc3826277, 32'hc2e89bc9},
  {32'h44703556, 32'h445eb065, 32'h432900da},
  {32'hc4bf69ab, 32'hc30f427b, 32'hc4aed6c2},
  {32'h4483e761, 32'h43b0ce34, 32'h43979ca8},
  {32'hc3cb8c7c, 32'hc4e3721c, 32'hc461e8c2},
  {32'h45436748, 32'h443ff12e, 32'h43cd8e0a},
  {32'hc52c749f, 32'hc1c67294, 32'hc36e3aac},
  {32'h44ab5620, 32'h44cd91e5, 32'h432deba6},
  {32'hc4b9bf7b, 32'hc43be19d, 32'h4366d849},
  {32'h442b82b1, 32'h44252bc3, 32'hc27e8022},
  {32'hc54239cc, 32'hc1ad8318, 32'hc44ceede},
  {32'h449c1fca, 32'h42bb9729, 32'hc2c22857},
  {32'hc3341478, 32'hc0bc34df, 32'hc4fbefec},
  {32'hc4217169, 32'h44698d57, 32'h4457eef6},
  {32'hc0cf9500, 32'h43a80866, 32'hc34f129b},
  {32'h42829304, 32'h453a67d2, 32'h4396f1fd},
  {32'h44f7584d, 32'hc4631dab, 32'h43076b48},
  {32'hc42c3386, 32'h40dc2798, 32'hc202725c},
  {32'h442dfe0a, 32'h433c95e2, 32'hc4b735fd},
  {32'hc40b6f62, 32'h4437b25e, 32'h4514b566},
  {32'h43f11c90, 32'hc48d51f6, 32'hc42f1728},
  {32'hc30ef75c, 32'hc4435410, 32'h448a377d},
  {32'hc3a34e1f, 32'h4456e08b, 32'hc3a3ca3f},
  {32'h43f73548, 32'hc384679c, 32'h43dc8d04},
  {32'hc3e2ef83, 32'hc29e19f0, 32'hc53266ae},
  {32'hc4c031e4, 32'h4444b558, 32'h42e5292c},
  {32'hc352c2a0, 32'hc3f4da26, 32'hc415a21d},
  {32'h444ab862, 32'h44f6dc7b, 32'h44e43cf7},
  {32'h43ac7f1a, 32'hc4246aab, 32'hc3f620f8},
  {32'h449e9c05, 32'h42b93cb1, 32'h43507148},
  {32'hc24ee440, 32'hc5208750, 32'hc3e15ede},
  {32'hc3f9841c, 32'h44d79bd7, 32'h44485e5f},
  {32'hc4a5c7c4, 32'hc2cbaad0, 32'hc33b9475},
  {32'hc44d6074, 32'h452e27d8, 32'h42f867f6},
  {32'h452f6799, 32'hc4139a12, 32'hc1106b69},
  {32'hc510c79d, 32'h43405fee, 32'h44269fb0},
  {32'h445c4fa0, 32'hc31adf79, 32'h4380e9d4},
  {32'hc566cbe8, 32'h4383273b, 32'h44222a84},
  {32'hc42d6abf, 32'h42cfdff2, 32'hc415f4e7},
  {32'h44613578, 32'hc24e9852, 32'h43028e8f},
  {32'hc5443734, 32'h440d5bc2, 32'hc3fedb00},
  {32'h43edd014, 32'h440a881f, 32'h42601af1},
  {32'hc502b786, 32'hc459c34f, 32'hc09edc68},
  {32'h439d2029, 32'hc3dba70d, 32'h439ae645},
  {32'hc4611155, 32'h44c07f81, 32'h43131e16},
  {32'h43875fb6, 32'hc4607360, 32'h43713286},
  {32'hc3f72bbc, 32'h4402cf20, 32'hc357d705},
  {32'h44946074, 32'hc4596112, 32'h42029054},
  {32'h44c59154, 32'h439f05a7, 32'hc35aa877},
  {32'h44fb2149, 32'hc3a0bc2f, 32'hc3830c96},
  {32'hc440cea4, 32'h4445cf3c, 32'hc2daf921},
  {32'h43be8287, 32'hc4933e57, 32'hc3b33279},
  {32'hc361820a, 32'h44261739, 32'h4406283a},
  {32'h44a69fd0, 32'hc3749866, 32'hc2d2aed6},
  {32'hc2c572ff, 32'hc19e0c43, 32'h4492b9f9},
  {32'hc3b8519c, 32'hc4209071, 32'hc49a53ee},
  {32'hc4341b32, 32'h435fbaba, 32'h4428e5af},
  {32'h44982c50, 32'h43af5dcf, 32'h4321dd74},
  {32'hc3f6d87e, 32'h442c72c2, 32'h4499d009},
  {32'h4460d6ac, 32'h43312f19, 32'hc4870241},
  {32'hc37dd9c5, 32'hc048be70, 32'h44e92d79},
  {32'h44cd5715, 32'hc36dd095, 32'hc4040b8d},
  {32'hc521bc64, 32'hc0a1a456, 32'h4398edb7},
  {32'hc41aff28, 32'hc2fc75ad, 32'hc3f7b60a},
  {32'h4123d300, 32'h447c8c59, 32'h452464c5},
  {32'h4432be74, 32'hc38207b1, 32'hc5566fe8},
  {32'h454061a2, 32'h43077214, 32'hc445700a},
  {32'hc4a10552, 32'h43bec7ca, 32'h44e2e9be},
  {32'hc1bb0808, 32'h44199114, 32'h42ff1e0e},
  {32'hc3934a62, 32'hc51dd965, 32'hc2a47e3c},
  {32'h420b84c0, 32'h4559495a, 32'h43481a8d},
  {32'h44293c9e, 32'hc4c51ed6, 32'h43d771a4},
  {32'hc2947468, 32'h44ef73cf, 32'hc26cdefe},
  {32'hc4692db1, 32'hc511695d, 32'h431debfd},
  {32'hc4a78849, 32'h43ff8941, 32'hc14dcda3},
  {32'hc495cbaa, 32'hc2f95ac6, 32'h44df7d64},
  {32'h44d8c7ab, 32'h43ce1fb1, 32'hc48091de},
  {32'hc3bf0d48, 32'hc3c34e90, 32'h4470e6ca},
  {32'h438abef0, 32'h440d4e8e, 32'h43e7ca10},
  {32'hc3cd0cd0, 32'h41b958eb, 32'hc55dcbec},
  {32'hc349c91c, 32'h411437da, 32'h4501415c},
  {32'hc49f66c3, 32'hc48d9e21, 32'h4272dec6},
  {32'h439d38be, 32'h4489035e, 32'h43ac43ac},
  {32'h443ef438, 32'hc2d14536, 32'hc46a4756},
  {32'h44c028e2, 32'hc4054ce6, 32'h43d0484e},
  {32'hc543e1df, 32'h43a88a9c, 32'hc3f3c149},
  {32'hc35a4884, 32'h43a3af4b, 32'hc2c40965},
  {32'hc39d26cc, 32'hc4246266, 32'hc4c4aa5b},
  {32'hc3d48f61, 32'hc2d6675b, 32'h4545d044},
  {32'hc34ae238, 32'hc36db453, 32'hc49af807},
  {32'hc3897dcd, 32'h44e03076, 32'h4435cca8},
  {32'hc2c47513, 32'hc3e7646e, 32'hc4340c78},
  {32'h4485c18a, 32'h44248684, 32'h43c49e02},
  {32'h451cad4d, 32'hc2d7692e, 32'hc33c9529},
  {32'hc4172b7f, 32'hc483d92f, 32'hc23e033e},
  {32'h451afb60, 32'h444f7c40, 32'hc19dc8b3},
  {32'hc51f8389, 32'h42fd509a, 32'h3fe7b929},
  {32'h44835ce3, 32'h44be34fe, 32'hc13435e0},
  {32'hc4bfbfcd, 32'hc4caad2b, 32'h42ad395b},
  {32'hc495d312, 32'h431c3ae2, 32'h408a6e7c},
  {32'hc55ea7e6, 32'h43bda62c, 32'hc1c74800},
  {32'h4566059f, 32'h42f64958, 32'h42ef49c0},
  {32'hc4157052, 32'hc441e086, 32'h4453602f},
  {32'h43a130b0, 32'h44d2c684, 32'hc214d011},
  {32'hc43df709, 32'hc3e8a7ca, 32'h438da170},
  {32'h4395e22e, 32'h440aa2df, 32'hc4993340},
  {32'hc427b2cc, 32'hc432766d, 32'h4130cd64},
  {32'h448fa111, 32'h440690cc, 32'hc48dfcc6},
  {32'hc4bc1410, 32'hc3226bad, 32'h442e8181},
  {32'h4520477d, 32'h417432ee, 32'hc407fed1},
  {32'hc49360a2, 32'hc437d270, 32'hc382228a},
  {32'hc3979268, 32'h43ff4038, 32'hc2ea344e},
  {32'hc48d11d3, 32'hc5057b98, 32'h4361e7aa},
  {32'h44f542ec, 32'hc223d656, 32'hc3d7821e},
  {32'hc38eabee, 32'hc4c9164c, 32'h43b7112b},
  {32'h440152de, 32'h4467287b, 32'hc42209e4},
  {32'hc30c935b, 32'hc40e64de, 32'h4476f8cc},
  {32'h4374126b, 32'hc31b54b2, 32'hc4962e97},
  {32'hc55ae122, 32'h4364300d, 32'hc28b9182},
  {32'h451d7eac, 32'hc2942ae8, 32'hc4953bd8},
  {32'hc2c79020, 32'hc4b3ad54, 32'hc2c8f884},
  {32'hc20bb8e7, 32'h4529afad, 32'h43301679},
  {32'hc42f6a57, 32'h43a846cc, 32'hc38b0302},
  {32'h42468891, 32'h440665ce, 32'hc45ba8ff},
  {32'h42b2c24a, 32'hc51df05a, 32'hc38218ab},
  {32'h421c8726, 32'h4510f4e4, 32'hc2f0006b},
  {32'h450f6dcf, 32'h43c8c2cc, 32'hc2b56e2d},
  {32'hc4b2eabd, 32'h42e5a6e1, 32'h43a5381d},
  {32'h44ba2832, 32'hc3865ba4, 32'h447f3da7},
  {32'hc50f10fa, 32'h435c46cd, 32'hc450a9f8},
  {32'hc2fb77c3, 32'hc48dde95, 32'h4458f2bc},
  {32'hc33b30b7, 32'h44e7999c, 32'hc3264698},
  {32'h4505dbb4, 32'h43db9bff, 32'h43f921b9},
  {32'hc4cf382f, 32'h43913253, 32'hc3e5876b},
  {32'h43997d8f, 32'h43bb0ce1, 32'h44c3618b},
  {32'hc4d8235e, 32'h42675b3b, 32'hc47b2af6},
  {32'h43c8d5f4, 32'h43850a28, 32'h45154230},
  {32'h439cd327, 32'h4291b5f3, 32'h44442856},
  {32'hc2590130, 32'hc56dd042, 32'h428c602b},
  {32'hc4bdc105, 32'h44594152, 32'hc3150f16},
  {32'h4400c8c7, 32'hc46a347b, 32'hc3ad6b40},
  {32'hc35a7400, 32'h410c1040, 32'hc518e6ed},
  {32'h43e1c22e, 32'hc39c07bd, 32'h449cc7a2},
  {32'hc522003c, 32'hc35a4a80, 32'h41a7801e},
  {32'h44041b3c, 32'h43f26d86, 32'h4543d368},
  {32'hc4c3111e, 32'hc473e048, 32'hc4965833},
  {32'hc0261c80, 32'hc399df51, 32'h450a3268},
  {32'h42a751a0, 32'hc30cdd54, 32'hc49026c8},
  {32'hc1f461c0, 32'h44a0c87a, 32'h44d89e32},
  {32'h44c4cd4e, 32'hc3a18a1e, 32'hc3788339},
  {32'hc42a9ddc, 32'h4483541b, 32'h41a23886},
  {32'h440603b3, 32'hc406ea26, 32'h450b16f0},
  {32'hc4e64d10, 32'hc2a79d3d, 32'hc3fcd704},
  {32'hc3c6f928, 32'h43a6b5a0, 32'h44b9e38d},
  {32'hc39763b8, 32'h42fdbbca, 32'hc5152161},
  {32'h4133e400, 32'hc2f67b88, 32'h44ce166d},
  {32'h43fa9d22, 32'h44b00d77, 32'h44b505ba},
  {32'hc44ea9aa, 32'hc422cc7d, 32'hc3b67439},
  {32'hc3fa38fc, 32'h439260c1, 32'h45056c68},
  {32'h443809a5, 32'h431fcc84, 32'h441b29c7},
  {32'hc3dbb948, 32'h42935682, 32'hc4ac9a24},
  {32'hc2cdef9c, 32'hc53a503d, 32'hc3b21671},
  {32'hc45d4955, 32'hc3859581, 32'hc42072b6},
  {32'hc287c01f, 32'hc4370ea4, 32'hc1276096},
  {32'hc492fd0c, 32'h43979cc7, 32'hc1d24722},
  {32'h4559c7c0, 32'hc349df9e, 32'h431c1782},
  {32'hc4924468, 32'h43bc8ca6, 32'hc3cac5d8},
  {32'h4505b6cd, 32'h439303f8, 32'hc39d17bf},
  {32'hc482d98c, 32'h43974e33, 32'hc36252ce},
  {32'h44946c56, 32'hc4bb714d, 32'hc44d2bc6},
  {32'hc54599fb, 32'h43a4a263, 32'hc3a2fe53},
  {32'hc489313f, 32'hc3937738, 32'h4267d44f},
  {32'hc461e0f4, 32'h44b9ef83, 32'hc3a6fa09},
  {32'hc3ae67e0, 32'hc506c67a, 32'hc4005377},
  {32'h44435681, 32'h4143e02d, 32'h44070d9c},
  {32'h4308f950, 32'hc3956233, 32'hc55bfe7f},
  {32'hc4a77854, 32'h422c6d05, 32'h439a08fe},
  {32'hc3d190cc, 32'h423aa227, 32'h44b618b8},
  {32'h4346a996, 32'h44cb7d13, 32'hc415593c},
  {32'h43de547f, 32'hc3be3569, 32'h44b2b75c},
  {32'h4511ea67, 32'h43f4a025, 32'hc40ad5be},
  {32'h440bd1d1, 32'hc4a96ec4, 32'h44861ca9},
  {32'hc38c1e49, 32'h443de716, 32'h439b3758},
  {32'h44bd1069, 32'h43a68c08, 32'h43fc3fbf},
  {32'h42a24588, 32'h444c2f81, 32'h451e7c74},
  {32'h4387c6a3, 32'h4370b5a0, 32'hc39b138e},
  {32'h4542b015, 32'h4421bf30, 32'hc403ed73},
  {32'hc480c40f, 32'hc44007a5, 32'h44344254},
  {32'h440943b9, 32'h44280bae, 32'h433676c2},
  {32'hc3f0cc52, 32'h41d03af2, 32'h4519df64},
  {32'h424557b8, 32'h44264534, 32'hc4f51ae9},
  {32'hc40bdd10, 32'hc49cfd47, 32'hc1093230},
  {32'h4436a538, 32'h4358849e, 32'h42f94ef8},
  {32'hc49f718a, 32'h4451242d, 32'h443867c5},
  {32'h4548bc99, 32'h4353410a, 32'h438a17f7},
  {32'hc3ab7399, 32'hc4968d47, 32'h43e91940},
  {32'h44831ea6, 32'h44be7b89, 32'hc405cc45},
  {32'h44a1e441, 32'h414479ec, 32'hc3c9378e},
  {32'h453cce6a, 32'h43b1f8b9, 32'hc38eb170},
  {32'hc44a135d, 32'hc4d2e763, 32'h43200779},
  {32'h43a3bb07, 32'hc36e63ca, 32'h433d7fdd},
  {32'h4288ad53, 32'hc4a8d838, 32'h43896890},
  {32'hc4792dce, 32'h4471836e, 32'hc44057aa},
  {32'h448dd5ab, 32'h42f7417d, 32'h43db5e5c},
  {32'h43c86e90, 32'hc3ced61d, 32'hc35c410a},
  {32'h4537168a, 32'h43107462, 32'h44160e86},
  {32'hc519199b, 32'hc45ffcb0, 32'h434e930d},
  {32'h44b05847, 32'hc348888c, 32'hc2fb8804},
  {32'hc4978b14, 32'hc46768f5, 32'hc45b65e3},
  {32'h4540265c, 32'hc17d7ff1, 32'h43b117f5},
  {32'h442d40c8, 32'hc3aa9f44, 32'h40418000},
  {32'h448998f1, 32'h43715337, 32'h440cea35},
  {32'hc4035f4b, 32'h449fea5f, 32'hc518c8a6},
  {32'h44726de8, 32'h42fe86db, 32'h444824bb},
  {32'hc49155b0, 32'hc2f70b31, 32'hc4a088b0},
  {32'h4355dacc, 32'h447c2bca, 32'h44c97e7f},
  {32'h43e1137e, 32'hc41ab2e2, 32'h4311f3d8},
  {32'h451ffeb3, 32'h42ee60da, 32'h43e3ae83},
  {32'hc4711e93, 32'hc2c6b51b, 32'hc424b973},
  {32'hc4320b36, 32'h441d4c5e, 32'h43d808dd},
  {32'hc322703e, 32'hc51d597e, 32'hc3617571},
  {32'h43a49700, 32'h45490888, 32'hc1a2398b},
  {32'hc486c8d6, 32'h430baad0, 32'hc2ea5786},
  {32'h43dc5920, 32'h442027cf, 32'h4428d8cc},
  {32'hc4937358, 32'hc4e60d6f, 32'hc29cead8},
  {32'h4561ac77, 32'h438d2732, 32'h43e7d25e},
  {32'hc58aecee, 32'hc325b20b, 32'hc3e7a97b},
  {32'h450af375, 32'h41290145, 32'h422fbaf3},
  {32'hc30b51ad, 32'hc21a545b, 32'hc484945d},
  {32'h42a5f9d8, 32'hc3e21e0e, 32'h44b88791},
  {32'h43817bdb, 32'h449c10ee, 32'hc411d744},
  {32'h42f720b6, 32'h450187f6, 32'h44647cbb},
  {32'h441ecde4, 32'hc49e31f2, 32'hc42919c8},
  {32'hc536b86b, 32'hc385dea3, 32'h4403c98c},
  {32'h450c2d07, 32'hc39fcf98, 32'hc45f8485},
  {32'hc3e87896, 32'h4433aa60, 32'h44aa344a},
  {32'h44f69b6d, 32'hc3f8a752, 32'h42cdbf39},
  {32'hc47a75f9, 32'hc35228fb, 32'h4453ce02},
  {32'hc25fb7f0, 32'hc2c015c0, 32'hc48daaa5},
  {32'h42e92012, 32'hc29ec860, 32'h4413a719},
  {32'h4395a156, 32'hc5202bd0, 32'hc3a47852},
  {32'hc438aaa4, 32'h434df2ee, 32'h4451d2c0},
  {32'h45246884, 32'h43c82031, 32'hc339eadd},
  {32'hc4126471, 32'h44866e3f, 32'h4481fbfb},
  {32'hc37ded1e, 32'hc500be48, 32'hc4bdc469},
  {32'h44345742, 32'h4373256e, 32'h43fb9eab},
  {32'h45783506, 32'hc40c1aa4, 32'h43406d03},
  {32'hc373b588, 32'h45188667, 32'hc2fc3a71},
  {32'h455a1c89, 32'h429dbb81, 32'h4376b871},
  {32'hc4e0328b, 32'h44ab1fca, 32'h433a46e4},
  {32'h449325e1, 32'hc39a4a02, 32'hc1c4b1d4},
  {32'hc49c1708, 32'h43fbb885, 32'h41571376},
  {32'h44a6b30f, 32'h42562a27, 32'h4383210f},
  {32'hc533a92c, 32'hc434d705, 32'h43147275},
  {32'h44e7211c, 32'hc3dd7ef7, 32'hc3c1ea94},
  {32'h447fc6ff, 32'h42ceda70, 32'hc263f500},
  {32'hc582f144, 32'hc410983a, 32'h438e92e7},
  {32'h45107bee, 32'h435d75e2, 32'h43ae6351},
  {32'hc4feb862, 32'hc4081573, 32'hc3d1653e},
  {32'h44fa276b, 32'hc47df6a0, 32'hc3900ae5},
  {32'hc515f8ac, 32'h43e1c877, 32'h43089678},
  {32'h4420b60d, 32'hc48efc40, 32'hc30e9bc6},
  {32'hc3d8ca8a, 32'h45006332, 32'hc3332e47},
  {32'h4512250a, 32'hc4080466, 32'h438db822},
  {32'hc460f568, 32'h42870585, 32'hc3f471be},
  {32'h4513485d, 32'hc38c6f46, 32'h4364a65b},
  {32'hc3d9f0ad, 32'h4402b3e7, 32'h4454873f},
  {32'h42c4d529, 32'hc208c94e, 32'hc4716372},
  {32'h431f43e4, 32'h44ad6e8d, 32'h441ad99c},
  {32'h4485a21f, 32'hc3089423, 32'hc3e4dabc},
  {32'hc4f78ec9, 32'h43922119, 32'h430ad54c},
  {32'h44463f72, 32'h440c38f8, 32'hc43d725f},
  {32'h4345fac6, 32'h446e4481, 32'h44778b51},
  {32'h44b6b4c5, 32'hc4052ba9, 32'hc386f6a1},
  {32'hc562c97c, 32'h43a64ce8, 32'hc225bbac},
  {32'h441ecb34, 32'hc4913d2b, 32'hc4e9c67e},
  {32'h44917d09, 32'hc35134a7, 32'h438e54eb},
  {32'h439faf7e, 32'hc52a9ee1, 32'hc30f5587},
  {32'hc4ab40f1, 32'h43c9ea32, 32'hc289ac69},
  {32'h42fea1bf, 32'hc1a2560c, 32'hc4fc1be7},
  {32'hc4721f5c, 32'h44403dcc, 32'h4499be2c},
  {32'h44062807, 32'hc476fc0a, 32'hc4a1d6e0},
  {32'h452702b2, 32'hc191e6cb, 32'hc2281b7d},
  {32'hc56d574a, 32'hc2c62fc0, 32'h3faaf700},
  {32'h45275395, 32'h43d1ecea, 32'h43074a96},
  {32'hc3e7bfc4, 32'hc5157b91, 32'hc37cbfd0},
  {32'hc33258db, 32'h4577ba7d, 32'h4388eb99},
  {32'h44e79f80, 32'hc3326138, 32'hc38d01ee},
  {32'h442bc460, 32'h44a1cb4c, 32'h421f8635},
  {32'hc46258dc, 32'hc5212fc9, 32'h43b4d701},
  {32'h43dd606c, 32'h441d230b, 32'h431dc2d9},
  {32'hc2f3dfac, 32'hc3654dd4, 32'h452250e5},
  {32'h44936a8a, 32'h4390d640, 32'hc4be4235},
  {32'hc5126e2e, 32'hc3c387cb, 32'h4181b15b},
  {32'h4412aff8, 32'h445fd6f8, 32'h437617ad},
  {32'hc51306d2, 32'hc2b3fbcb, 32'hc2674f3a},
  {32'hc5051629, 32'h438b9c04, 32'h435f5926},
  {32'hc19689c0, 32'h423f12ac, 32'hc513f0b6},
  {32'h44003fbe, 32'h44477980, 32'h44e657e2},
  {32'hc4f2b7ab, 32'hc321bf99, 32'hc2fbe554},
  {32'h43a7ab80, 32'h409b3c98, 32'h44986cd7},
  {32'hc507d4de, 32'h4401736b, 32'hc3d2c4c8},
  {32'h44260c18, 32'hc407b518, 32'h43fd9024},
  {32'hc46d240b, 32'hc49380ed, 32'hc408d7a0},
  {32'h43c2f65f, 32'h4169c700, 32'h44c61f0e},
  {32'hc520cfc9, 32'hc32e206e, 32'h43bd4486},
  {32'h4326fb28, 32'h4528344d, 32'h43a80144},
  {32'hc4be98da, 32'hc4d3202b, 32'hc2bd2513},
  {32'h4434930a, 32'h42f38d3f, 32'h4434b023},
  {32'h4529b71c, 32'hc3ce5762, 32'hc413b217},
  {32'hc52c793e, 32'h429c5cd2, 32'hc33e27e6},
  {32'hc285e2e0, 32'h44f85a0f, 32'hc3b00166},
  {32'h4400f94b, 32'hc3e0f641, 32'h42a5a856},
  {32'h43ba066e, 32'h45098eb5, 32'hc2c4fdfe},
  {32'hc4505aee, 32'hc495691a, 32'hc377c502},
  {32'h45119fc2, 32'h42aaa110, 32'hc3d434f6},
  {32'hc51757dd, 32'hc31cb1fc, 32'hc3c8ea8c},
  {32'h451ba406, 32'hc3fdb809, 32'hc2959fd6},
  {32'hc4fa3ee9, 32'hc34928cb, 32'h435d7b32},
  {32'h44738e96, 32'h448c425b, 32'hc30b361f},
  {32'hc4fa785f, 32'hc2f9d227, 32'hc3145543},
  {32'hc488ba10, 32'h43ca4dbd, 32'hc2e5007c},
  {32'h43479fb2, 32'hc4b1a9a6, 32'h442fce81},
  {32'h442532db, 32'h4227a5c8, 32'hc508e156},
  {32'hc522b0b2, 32'hc25d89d0, 32'hc26f287c},
  {32'h44430fa6, 32'h42f91686, 32'hc46c7892},
  {32'hc3b32230, 32'hc4045ac2, 32'hc3d54b5a},
  {32'h433fdcbe, 32'h440b9177, 32'hc420e540},
  {32'hc308b854, 32'hc4c81790, 32'h43757557},
  {32'h451c5129, 32'h434b8f04, 32'hc46f0bc4},
  {32'hc24c8186, 32'hc2cbf8e4, 32'h44fab77b},
  {32'h4534d480, 32'h4424f48a, 32'hc39840c8},
  {32'hc2b61120, 32'h4361642b, 32'h45540dc3},
  {32'hc4103a90, 32'h41b212ba, 32'hc3256a8b},
  {32'h41ad3100, 32'h44a8d54c, 32'h451a28b5},
  {32'h44c4bf01, 32'hc3e17332, 32'hc4ab0c24},
  {32'h4413a4ec, 32'hc4979a1f, 32'hc343d3a9},
  {32'hc3e1b328, 32'h4532c87f, 32'hc39dbb02},
  {32'h44d38c76, 32'h43a388b7, 32'h43db12ee},
  {32'hc4e43cc4, 32'h4426ffbe, 32'h4436de9e},
  {32'h43e48490, 32'hc4bba651, 32'h430760ba},
  {32'h449c4dd9, 32'h43b5196f, 32'h43126db4},
  {32'h4531453c, 32'h4440b7bb, 32'h428c971e},
  {32'hc5356d09, 32'h43b9d1ad, 32'h43dd3ae3},
  {32'hc41aae7a, 32'hc44094fc, 32'h43a1d5ce},
  {32'h423234f8, 32'h44dbc82d, 32'h4395af43},
  {32'hc2226400, 32'hc47c348f, 32'h443d0b50},
  {32'h43e1871e, 32'h43d88376, 32'hc46e0fda},
  {32'h43a96351, 32'hc361d766, 32'h44fdbf62},
  {32'hc3cfc588, 32'h4435bad1, 32'hc473b25d},
  {32'h4419f3e0, 32'h432f3125, 32'hc31b849a},
  {32'hc3a737dd, 32'hc3ca0b31, 32'hc4db85f2},
  {32'h43cbfb38, 32'hc44ebc9c, 32'h43fc5243},
  {32'h440ecf23, 32'hc3b67098, 32'hc46af327},
  {32'h444da0cb, 32'hc4b0ebb0, 32'h452818e0},
  {32'hc5344353, 32'h43c578e5, 32'hc38b8e3c},
  {32'h44faef87, 32'h44288de8, 32'hc387aa63},
  {32'hc3edd898, 32'h45143871, 32'hc3e50bc9},
  {32'hc36b992e, 32'hc51153f8, 32'h442c182a},
  {32'h447c9a8e, 32'hc36a4c36, 32'hc49f89c3},
  {32'h42804c40, 32'h44201ba8, 32'h451b86bb},
  {32'hc4d74884, 32'h43c4a1f4, 32'hc4d64858},
  {32'h45224972, 32'hc2627b78, 32'hc1e6303a},
  {32'hc44a8c32, 32'hc41926dc, 32'hc4964966},
  {32'h42a1efb4, 32'hc43cba4e, 32'h44768c69},
  {32'h43373847, 32'h4485eccf, 32'hc4479b35},
  {32'hc51bcebe, 32'hc2bd15ee, 32'h4314c2aa},
  {32'h43aa1e30, 32'hc45c5c6b, 32'h44bf4717},
  {32'hc348971c, 32'h43e0e673, 32'hc50051fa},
  {32'h44e1edfe, 32'h41ebac35, 32'hc3d4609c},
  {32'hc33b3c0c, 32'h455b765d, 32'h42fa6dfe},
  {32'hc31c6cf8, 32'hc0750490, 32'h45841f0f},
  {32'h44742848, 32'hc12865da, 32'h44a00163},
  {32'hc34c5910, 32'hc4d57cec, 32'hc49b3d2a},
  {32'hc49ffcf0, 32'hc294acb6, 32'h43fe30fd},
  {32'h417e64c2, 32'hc4c9e1f9, 32'h42a3c7f2},
  {32'hc482f4a2, 32'h4382f673, 32'hc3ffd759},
  {32'hc2234da0, 32'hc4cc1b73, 32'h41168a20},
  {32'h4425996b, 32'h442be679, 32'h4396df6d},
  {32'hc1c9879c, 32'hc55cd790, 32'hc26088ae},
  {32'h4294cce8, 32'h4485994b, 32'hc4907c42},
  {32'h45252009, 32'hc3f115a5, 32'hc1a7d6a3},
  {32'hc4fec999, 32'h433b6776, 32'hc42d90c5},
  {32'h450d88e2, 32'h4362a4a0, 32'hc40e6190},
  {32'hc32182d7, 32'h4464c2eb, 32'hc43f69ec},
  {32'h44e4cd5b, 32'hc49b54bd, 32'h42ec6ce7},
  {32'hc467eca4, 32'h4411d536, 32'h434a6f82},
  {32'h43166abe, 32'hc474c918, 32'h43605345},
  {32'hc4647dc9, 32'h44b01199, 32'h43142025},
  {32'h4432c5f0, 32'hc4c2fba5, 32'hc23eda18},
  {32'h44184ecb, 32'hc4c94c3e, 32'h43a55d8b},
  {32'h44f378f9, 32'hc30de0e1, 32'hc33d5519},
  {32'hc30d4d84, 32'hc4fc1ed7, 32'h450f40f4},
  {32'hc4aff43c, 32'h440484fd, 32'h4488e92e},
  {32'h44b662ba, 32'h43b23f4c, 32'hc311f8e9},
  {32'hc496fc8e, 32'hc39c4c1d, 32'hc2f5a0d4},
  {32'h436e6c98, 32'h4469be34, 32'hc44615fc},
  {32'hc3a87524, 32'h41f91970, 32'h4581105d},
  {32'hc3930ddf, 32'h443c4c9d, 32'h4395e398},
  {32'hc361ba66, 32'h43f77797, 32'hc4523982},
  {32'hc49c468e, 32'h43c9ff00, 32'h448ae3aa},
  {32'h4382b5d8, 32'hc257614f, 32'hc4d848b5},
  {32'h43cb1fcb, 32'h43c18717, 32'hc4e96011},
  {32'hc4e89f05, 32'hc3702e6d, 32'hc29747f4},
  {32'hc49e93e4, 32'h43420769, 32'hc348e9e8},
  {32'hc49dc856, 32'hc28b11de, 32'h44e7b99e},
  {32'hc400cafd, 32'h454f1365, 32'hc2803638},
  {32'hc4fe96e7, 32'hc3a126f1, 32'h434a148d},
  {32'h44cb0ff4, 32'hc4139aec, 32'hc41b89c4},
  {32'hc4971933, 32'hc37322b1, 32'h42af5f61},
  {32'h450bed0d, 32'h43a8776e, 32'h43ad23cc},
  {32'hc560fd75, 32'hc40c032d, 32'hc27a2eac},
  {32'h43db866a, 32'h456ac5e7, 32'h42b794bd},
  {32'hc4fe4608, 32'hc34850ae, 32'h3cd92d00},
  {32'h45089740, 32'h44827639, 32'h438029d6},
  {32'h40cfae00, 32'hc5108278, 32'hc3ae5e32},
  {32'hc36d247f, 32'h44ce6cb5, 32'h43adca6b},
  {32'h4482d578, 32'hc39db32e, 32'h40a4f468},
  {32'hc4a24989, 32'h44262ce6, 32'hc34d286a},
  {32'h4346ef91, 32'h44f060f4, 32'h440ec70d},
  {32'h4505a695, 32'hc314dfe6, 32'hc16f98f6},
  {32'hc1e521f4, 32'h455c5f7d, 32'h437c523f},
  {32'hc406c1f8, 32'hc4ee5a70, 32'hbdddbc80},
  {32'hc347646c, 32'h44446714, 32'h44848785},
  {32'hc4d59258, 32'hc4ecf7fd, 32'hc4b54689},
  {32'h44bd4f9d, 32'hc22d7b38, 32'h44b13634},
  {32'hc28cee25, 32'h44196372, 32'h430ef9de},
  {32'h44be33b8, 32'h44186d24, 32'hc3834a19},
  {32'h4404f43c, 32'h44767524, 32'hc4b745f4},
  {32'h44068b5c, 32'h439af5eb, 32'h442d3fdf},
  {32'hc50de7eb, 32'hc33d3c92, 32'h42e0628e},
  {32'h44ff5c4e, 32'h43c83ba8, 32'h4303f1bb},
  {32'h441db948, 32'hc346ae20, 32'hc1b6fc2c},
  {32'h4455ac3e, 32'h4434517d, 32'h448c4b2c},
  {32'hc39e8956, 32'hc35e405e, 32'hc48ab719},
  {32'hc39e7d15, 32'h444bbfa3, 32'h41c90b3d},
  {32'hc513e482, 32'hc43adcc2, 32'h43c7f2a6},
  {32'h433d82a4, 32'h44e902d6, 32'h4354bc8c},
  {32'hc41fc4a1, 32'hc3ca6677, 32'hc3ccc2f0},
  {32'h44a9798e, 32'h441a4308, 32'h443fa719},
  {32'hc42e8015, 32'hc52e1d9e, 32'h40ac23ce},
  {32'h44092bce, 32'h43b1ced5, 32'h4242e46c},
  {32'hc3407658, 32'h42beb777, 32'h43a44c4d},
  {32'h44b34d10, 32'hc3cab734, 32'h43ebea59},
  {32'h42d911cc, 32'h4347e488, 32'hc519b8a2},
  {32'h42309bbc, 32'hc48a7b8a, 32'h446d7166},
  {32'h436649d7, 32'h436a0be0, 32'hc3600685},
  {32'h436a2c68, 32'h446eb487, 32'h44eb4eac},
  {32'hc40d5b74, 32'hc3e70067, 32'hc5493727},
  {32'h44d8a14c, 32'hc2b300c2, 32'h42823a46},
  {32'hc3cd7861, 32'hc3e3ac06, 32'hc4cb5d08},
  {32'hc304514e, 32'h449242fc, 32'h44f3d593},
  {32'h4511a09e, 32'hc2cec91f, 32'h43ed66d2},
  {32'h43a7105d, 32'hc490f13e, 32'h4517208b},
  {32'hc3a8a6f8, 32'h43eb70e9, 32'hc4b20e44},
  {32'hc4d3108a, 32'hc3b65a6f, 32'hc3864b21},
  {32'h450ff46c, 32'h4301893e, 32'hc361e3be},
  {32'hc4848d88, 32'h44d058be, 32'h431553d6},
  {32'h45004d87, 32'h436765f4, 32'h42a546f0},
  {32'hc51e2434, 32'hc30f704f, 32'h4432d814},
  {32'h4466c2aa, 32'hc4c5b10f, 32'hc4636fcd},
  {32'h43677be8, 32'hc3f112d2, 32'h44902dc3},
  {32'h45413b99, 32'hc47191ef, 32'hc2aa18f0},
  {32'hc51215b4, 32'h4426e483, 32'hc3665cd5},
  {32'h441b982a, 32'hc31f95b0, 32'hc2d7acf4},
  {32'hc4cb123f, 32'h4415e788, 32'hc33ac043},
  {32'h448c720e, 32'hc5602e45, 32'hc315f9ca},
  {32'h44981d5b, 32'h440a0e54, 32'hc3c10af1},
  {32'h441aa9f5, 32'h43b039ad, 32'hc418964c},
  {32'hc4357ce8, 32'hc40fbd02, 32'h43b3c743},
  {32'h448f8612, 32'h4325f36c, 32'hc2860383},
  {32'h44c06efe, 32'h42ffcbb6, 32'hc34ec309},
  {32'hc4c3e30f, 32'h437f232b, 32'hc4fa2f5f},
  {32'hc36d5b90, 32'h43e0aa06, 32'h4396be88},
  {32'hc493236d, 32'h43baf757, 32'h42b483e8},
  {32'h44f631bc, 32'hc479c91b, 32'h4326363b},
  {32'hc3748ecd, 32'h45436837, 32'h439e1b05},
  {32'h45217de0, 32'h43e2a132, 32'hc3a1c249},
  {32'hc5445f18, 32'h443bf424, 32'h434d08e9},
  {32'h4310b770, 32'hc4c6ac1d, 32'hc414e199},
  {32'hc4911a0d, 32'hc3e8ed6c, 32'h43ff028f},
  {32'hc2a6c7f2, 32'h43ac5bfe, 32'h4537d909},
  {32'hc4b6be8a, 32'h43e0d97f, 32'hc49a080f},
  {32'h44c03152, 32'hc2b528f5, 32'hc263cd86},
  {32'h42acb2d8, 32'h4502c9b5, 32'h43513929},
  {32'h4511ba43, 32'hc2ba1d0b, 32'hc30ab1c6},
  {32'hc4eb9c31, 32'hc0eaca59, 32'hc4022a1c},
  {32'h44416c77, 32'hc4e88621, 32'hc3b27c08},
  {32'hc415209a, 32'h44c34da1, 32'hc34d66d0},
  {32'h447a6617, 32'hc40e23f6, 32'hc3022de2},
  {32'hc4a58964, 32'hc42e7301, 32'h4422a131},
  {32'h455cbc0a, 32'hc3a0a0d4, 32'hc3f10814},
  {32'hc318bb57, 32'h44837476, 32'hc30cc907},
  {32'h42d139e3, 32'hc3065486, 32'hc53554d9},
  {32'h438d0fb7, 32'h453eba78, 32'h42be930f},
  {32'h445eeb96, 32'hc40cfd34, 32'hc4173fc3},
  {32'hc3dce6ac, 32'h433f184c, 32'h432350a2},
  {32'h45034737, 32'hc42b4bcf, 32'hc4a4a005},
  {32'h44c4e6b0, 32'hc09cdf3c, 32'hc2be84ac},
  {32'hc4b8acd0, 32'hc311c9fd, 32'h43a4f1ac},
  {32'h45413a1e, 32'h43c5f056, 32'h43e7bb16},
  {32'hc4ea50b2, 32'hc38d4694, 32'h43f5a663},
  {32'h44c97ffc, 32'hc2d3864e, 32'hc2b52df1},
  {32'h449621c8, 32'hc3b149fe, 32'hc3f757b8},
  {32'h4513fb04, 32'h4499e6cf, 32'hc25c59d8},
  {32'hc4b4cc5e, 32'hc4d260db, 32'hc3e9e129},
  {32'h43ee5856, 32'h45294018, 32'hc135085a},
  {32'hc4d5cd01, 32'hc3b6cc3f, 32'hc3ed4124},
  {32'h44355658, 32'h43740c42, 32'hc39abeef},
  {32'h44d1a2d6, 32'hc169334e, 32'h4308d372},
  {32'hc305b67a, 32'h44d106ab, 32'h442ae643},
  {32'hc4a0351b, 32'h430dc1c5, 32'hc43b4a59},
  {32'h43a957cd, 32'h44075148, 32'hc21e4f2b},
  {32'hc3e6e15a, 32'hc49a92ad, 32'hc4847f4c},
  {32'h445110e5, 32'h44e5a242, 32'h443c4eaf},
  {32'hc5093a8e, 32'hc40e287a, 32'h43ec1ada},
  {32'hc30eea40, 32'hc4ac9ee7, 32'h44f6c27f},
  {32'hc50b11ee, 32'hc3cf96de, 32'hc42d8b88},
  {32'h45057be4, 32'hc3958131, 32'hc3a70506},
  {32'hc50f2f11, 32'hc3e10690, 32'hc3902b09},
  {32'h43e4c98f, 32'h44587ba5, 32'h439e883d},
  {32'h42c03710, 32'hc489c0cc, 32'hc43b3af2},
  {32'h434af0e8, 32'h452c9a27, 32'h43b30845},
  {32'hc4553eee, 32'hc3c1bf17, 32'hc52a384a},
  {32'hc003a920, 32'hc247b979, 32'h44cea705},
  {32'hc48ecf8e, 32'h44042584, 32'h43824aac},
  {32'hc4cbdf28, 32'hc43ee1d6, 32'hc3a09880},
  {32'h42184bc9, 32'h4555626b, 32'hc2c43cd2},
  {32'h43a87ecb, 32'hc4ae2465, 32'hc399cf9d},
  {32'h44d858a6, 32'h4487e5bc, 32'hc39b0115},
  {32'hc40f139f, 32'hc4febe41, 32'hc2412f02},
  {32'hc46904ff, 32'h44233b6f, 32'h43a35225},
  {32'hc466eed2, 32'hc4984a58, 32'hc4a6b68c},
  {32'h44a59d1c, 32'h447b0473, 32'h4457bd5a},
  {32'hc413f178, 32'hc4351b77, 32'h4448fc1a},
  {32'h448e1912, 32'h43f984d5, 32'hc2e6eb8a},
  {32'hc2f51d48, 32'hc3a5d472, 32'h4501d44e},
  {32'h448cd33c, 32'h434f0343, 32'hc45c0e95},
  {32'hc4a30356, 32'hc33fa156, 32'h44147170},
  {32'h435f5217, 32'h42c1aca0, 32'hc53fa558},
  {32'hc494b751, 32'hc2bf33c1, 32'hc335ce91},
  {32'h441984fe, 32'hc39c0a62, 32'hc4c858bb},
  {32'hc445da37, 32'h4384d9c7, 32'h44f2577c},
  {32'h4532e7b9, 32'hc29e6e90, 32'hc47eb72f},
  {32'hc4b3a118, 32'hc4a0ea29, 32'h43ffd408},
  {32'h4496e41c, 32'h44847e52, 32'hc4113df0},
  {32'h42abf778, 32'hc50da5ef, 32'hc438389c},
  {32'h42b510e8, 32'h42de8e46, 32'hc520ade4},
  {32'hc434d230, 32'hc4114d1e, 32'h44b24518},
  {32'h430d3cda, 32'hc2141c6c, 32'hc3c55177},
  {32'hc5084784, 32'h42fa08de, 32'h43a72e3e},
  {32'h4520eb48, 32'hc377a34d, 32'hc494fbe6},
  {32'h44af499e, 32'hc4942f94, 32'hc457772f},
  {32'hc5038a97, 32'h44450b75, 32'h431246ed},
  {32'h427ec273, 32'hc4ea47f6, 32'hc2a2b7a5},
  {32'hc4d7e4fd, 32'h4430ac90, 32'h437a673a},
  {32'h4494290f, 32'hc42c2409, 32'h433f6d76},
  {32'hc40c0328, 32'hc391bd40, 32'hc35ffa45},
  {32'h44d956e4, 32'h43c7d69c, 32'h41158671},
  {32'hc428b876, 32'h43c1f2d0, 32'h43c78563},
  {32'h454d515e, 32'h4301c0fd, 32'h429d936f},
  {32'hc4996165, 32'h43a8766d, 32'hc38aa500},
  {32'hc36f07b4, 32'hc4d17be7, 32'h434b3b49},
  {32'hc44e338c, 32'hc2478994, 32'hc40e82d1},
  {32'hc345420c, 32'hc4abd563, 32'h445f9a3f},
  {32'hc3511456, 32'h448bf077, 32'hc41ee899},
  {32'h4464b88f, 32'hc2155f5b, 32'h4402e23b},
  {32'hc3a358e6, 32'hc398df86, 32'hc51e95e7},
  {32'h438a14c0, 32'hc2342b88, 32'h44e06b6c},
  {32'hc31255f0, 32'h433c31e2, 32'hc4d61244},
  {32'h43aac9e8, 32'hc4c71578, 32'h44c7848c},
  {32'hc55afd78, 32'h43ca8f1d, 32'hc206e8fd},
  {32'h4512c175, 32'h43912fdb, 32'hc3981bed},
  {32'hc3880466, 32'hc369686d, 32'hc498e92b},
  {32'h44bce940, 32'hc4a14ce2, 32'hc3c817da},
  {32'hc4d48d48, 32'h43be0291, 32'h437f8cd9},
  {32'hc36e5ec2, 32'h4393066d, 32'h44be8c97},
  {32'hc52e1b95, 32'h43cc0ed6, 32'hc48443cd},
  {32'h44b8a88c, 32'hc329c083, 32'h4370ae1f},
  {32'hc48db0ba, 32'hc4a20627, 32'hc48d953c},
  {32'h448ae4cc, 32'hc450c662, 32'h444426d0},
  {32'hc4c200c0, 32'h44272b0f, 32'hc3a31c82},
  {32'h434a6d98, 32'h43a7dc89, 32'h417622c2},
  {32'h44b20faa, 32'hc461d787, 32'hc36de4a3},
  {32'h42a2aefc, 32'h448f8201, 32'hc3f2de38},
  {32'hc4614dfa, 32'hc2f5c642, 32'h440211d6},
  {32'hc4850e94, 32'h430faa5e, 32'hc50efde6},
  {32'h433cafa0, 32'hc461b6bd, 32'h4480415d},
  {32'hc373d8e0, 32'hc38c3a4d, 32'h4509bbc4},
  {32'hc56a6881, 32'h41da36fc, 32'h42d76c6e},
  {32'h4432043c, 32'h445c9ab9, 32'h420f5645},
  {32'h43f9d24f, 32'hc31d9ea9, 32'h446c8c11},
  {32'h4221e6a4, 32'hc38a6ad3, 32'h439381fb},
  {32'hc3f56fc2, 32'h43bb3cc4, 32'h45018522},
  {32'h4408d3a2, 32'h440fbcad, 32'hc496427f},
  {32'h43857aaa, 32'hc35ab6d9, 32'h45295f61},
  {32'h4373a6ae, 32'h45078cfe, 32'hc39ebdc4},
  {32'h44376f9b, 32'hc425c0fc, 32'hc361a5e5},
  {32'hc5278c84, 32'hc3aa088e, 32'hc3abe64e},
  {32'h42016440, 32'h44569dcb, 32'h43721b1c},
  {32'hc54bb2f0, 32'hc242d7cb, 32'hc2c1fb49},
  {32'h440f2319, 32'hc5314b27, 32'h43feed11},
  {32'hc39cb2a2, 32'h450fa638, 32'h43ded2b3},
  {32'h4426dc97, 32'hc40d60cb, 32'h43cc977f},
  {32'hc50bfdc0, 32'h43d0a00b, 32'hc3f505a7},
  {32'hc3c624a5, 32'hc58a2a85, 32'h4311f4b4},
  {32'h444759ca, 32'h434e0e32, 32'h43f1a02f},
  {32'hc20ec4a0, 32'h4448374c, 32'hc497e7af},
  {32'h42f489a8, 32'h44a80311, 32'h44f0fefe},
  {32'hc494e47f, 32'hc43cdb17, 32'h42d3ca3a},
  {32'h44cba12c, 32'h43049c86, 32'hc342e6b3},
  {32'hc4a7f447, 32'h41c2d520, 32'h440a6ba4},
  {32'h449ead07, 32'h4417b97e, 32'hc3c95fbc},
  {32'hc1c57140, 32'hc42f17d6, 32'h4511fff8},
  {32'h44e34ccc, 32'hc29eb00c, 32'h434469ec},
  {32'hc3178970, 32'hc30b64c9, 32'h43ba7f26},
  {32'hc42dcae0, 32'hc4ec3e3e, 32'h44fb0c18},
  {32'h44dc5d70, 32'h444a8b6c, 32'hc44b6d38},
  {32'h44a7da60, 32'h44221883, 32'hc3b72f9a},
  {32'hc51eed2c, 32'hc3009ae2, 32'hc3a43e59},
  {32'h4409cf87, 32'h41141e3c, 32'hc4bb6e8f},
  {32'hc3a453fd, 32'h42aa8ada, 32'h452ae5ab},
  {32'hc2ad0180, 32'h4462ca82, 32'hc49fb29f},
  {32'h428176ef, 32'hc335456f, 32'h44b3c002},
  {32'h455a42d9, 32'hc418f2cc, 32'h4303ea19},
  {32'hc564fc2a, 32'hc405c000, 32'hc2d0690f},
  {32'h44db5b9c, 32'h43cf629d, 32'h437d861f},
  {32'hc491ee00, 32'hc4f71ff6, 32'h430a3ba6},
  {32'h440defeb, 32'h4504bed2, 32'h43be8d50},
  {32'hc306d06f, 32'hc3d97a82, 32'hc387a072},
  {32'h44378f2a, 32'h44148b98, 32'h43935853},
  {32'hc5308bb6, 32'hc3a548c3, 32'h43a59fda},
  {32'hc486a705, 32'h443ebd20, 32'hc228a307},
  {32'h43d6eba4, 32'h42ff8f30, 32'h44c61e36},
  {32'hc40ad593, 32'hc5458ecf, 32'hc35bcf44},
  {32'h44003a3c, 32'h45377f44, 32'h43e2a4bc},
  {32'h450dcf36, 32'h43cabb87, 32'hc2d74e9b},
  {32'h455670a5, 32'h43559dce, 32'h42e0dc57},
  {32'h42495530, 32'hc37300ed, 32'hc492f0d1},
  {32'h4416fb47, 32'hc30a9aa2, 32'h44835b03},
  {32'hc3bba3f7, 32'hc4f86ebb, 32'hc4aec217},
  {32'hc3b12cd6, 32'h442247a8, 32'h456e9f48},
  {32'hc50c5c38, 32'h4360d8fa, 32'h4409c9aa},
  {32'hc10da9a0, 32'hc40ff7ae, 32'h44a83ce6},
  {32'h429d9313, 32'hc3e60f53, 32'hc48bb669},
  {32'h44d4ec4c, 32'h431128f4, 32'h426738ba},
  {32'hc4e70a7e, 32'hc2e7d74d, 32'hc45277e3},
  {32'hc27ed0c8, 32'h44b991cb, 32'h43ea8206},
  {32'h43e54732, 32'hc3475e14, 32'hc4c4833b},
  {32'h43888b60, 32'h4490e393, 32'h44821041},
  {32'hc4b0f1d8, 32'hc39013ad, 32'hc43bd49d},
  {32'hc1b28e62, 32'h44e78d99, 32'hc328580f},
  {32'hc36eea2d, 32'hc4ed9298, 32'hc3e86316},
  {32'h44bf7d6a, 32'h449832f2, 32'h4409ec16},
  {32'hc4a9c0ee, 32'hc348b0fb, 32'hc39db67d},
  {32'h43a1a25e, 32'h44f8240d, 32'hc2b8554f},
  {32'h432018f1, 32'hc5282896, 32'hc3e7b06e},
  {32'hc4442c48, 32'h43f3ed99, 32'h441d61ce},
  {32'hc517296c, 32'hc360caa0, 32'hc40edb40},
  {32'h450125f5, 32'h43a6bf89, 32'hc3df5b55},
  {32'h43c5c5c8, 32'hc3efecd2, 32'hc40b52e7},
  {32'h4390ac34, 32'hc4043ad5, 32'h44ea57af},
  {32'hc42c6f60, 32'hc424b18e, 32'h429d4616},
  {32'hc4464c90, 32'h449fe5d5, 32'h4412034e},
  {32'h40aee1ea, 32'hc41a48aa, 32'hc508817e},
  {32'hc4a572d5, 32'h430af5dc, 32'h43a7c2af},
  {32'hc26880b2, 32'hc44d574d, 32'hc4bbff23},
  {32'hc3f25ab0, 32'h44876bea, 32'h44dc697e},
  {32'h43ae0006, 32'hc4568f4c, 32'hc4a1d8b0},
  {32'h43da958d, 32'h44f35465, 32'h4327ecc5},
  {32'hc3273dbc, 32'h439e0f1a, 32'hc5011cda},
  {32'hc3cc345e, 32'h4428708b, 32'h43d7b8dc},
  {32'h44f643f2, 32'hc385feff, 32'hc3c63cb6},
  {32'hc5071a9d, 32'hc1d01494, 32'h440df2cd},
  {32'hc465a60f, 32'h4392ab05, 32'hc3903bcb},
  {32'h445620aa, 32'h441cb5ac, 32'h456df144},
  {32'h43cd3bbe, 32'hc480a90e, 32'hc4179829},
  {32'hc32f4298, 32'h42f23ec3, 32'h42005055},
  {32'h43f1152c, 32'hc55ea74f, 32'h439e11da},
  {32'hc4200d0c, 32'h44f98f06, 32'h4339d5e3},
  {32'h447515d6, 32'h433c807b, 32'hc346bbaf},
  {32'hc4549b5a, 32'h450a9ddd, 32'hc39cf2f7},
  {32'h43878aba, 32'hc3ef60c0, 32'h4315f513},
  {32'hc408bf36, 32'h447c5bd9, 32'h43419f62},
  {32'h450ee645, 32'hc3dbc812, 32'hc3f64d8f},
  {32'hc4ef953c, 32'hc3d89539, 32'h434f8e7f},
  {32'hc3f26afc, 32'hc2aca429, 32'h3f4d769f},
  {32'h440ed4a6, 32'h42b27591, 32'h4380461e},
  {32'hc14046f5, 32'hc1fcab1f, 32'hc55995c1},
  {32'h448e65b4, 32'hc2a80837, 32'h4504a58d},
  {32'h4440b393, 32'hc3ada9e9, 32'h40246822},
  {32'h451f8f31, 32'hc27b50be, 32'h42720966},
  {32'hc3176892, 32'h452e2cff, 32'h439c0071},
  {32'hc4901261, 32'hc3a799f4, 32'h433ffbe7},
  {32'hc40f1f20, 32'h4531a9dc, 32'hc3a1ba09},
  {32'h4418847e, 32'hc4efe386, 32'hc382157d},
  {32'h43fb5ac0, 32'h427afc6a, 32'hc436546c},
  {32'h446016b2, 32'h441d9075, 32'h451366ca},
  {32'hc42938a4, 32'h449424b6, 32'h445c7998},
  {32'hc3c672fb, 32'hc319966b, 32'h442fe6bc},
  {32'hc50dc0d7, 32'h43f231ba, 32'h435cd3cd},
  {32'h431e121d, 32'hc4946c9c, 32'hc515b137},
  {32'hc1bde155, 32'h44183219, 32'h441f9fed},
  {32'hc1fe1cca, 32'hc316dc13, 32'hc39bf6fa},
  {32'hc3c96918, 32'h44b157a5, 32'h4467856c},
  {32'h45555233, 32'hc40d6e08, 32'h43c3a21f},
  {32'hc58db325, 32'hc31b39dd, 32'hc31ba60f},
  {32'h43c52948, 32'h445cb1ad, 32'hc4ce3e06},
  {32'hc3a6754f, 32'h42b05b22, 32'h41bbf48a},
  {32'hc447dca3, 32'hc4f01ef2, 32'hc3d49b0e},
  {32'h436b4ed2, 32'h453e8940, 32'h4415eb93},
  {32'h4551becb, 32'h43ab5a4a, 32'h43f4d80e},
  {32'hc4086344, 32'h43944260, 32'h44b36e6d},
  {32'h43e3d944, 32'hc4aff95e, 32'hc3d75d3d},
  {32'hc329a6e4, 32'hc3c25988, 32'hc4be39bf},
  {32'hc44ace38, 32'hc25ef6d1, 32'h451b43b1},
  {32'h4526c8b4, 32'h4379c6f0, 32'h43af21cb},
  {32'hc3dbe13a, 32'h4318727c, 32'hc3f38b85},
  {32'h4481cd6f, 32'h4413dc66, 32'h43bcbce9},
  {32'hc4a3b3b6, 32'hc39b619d, 32'hc1012aca},
  {32'h451fc20b, 32'h444ac3d9, 32'h4358064a},
  {32'hc5632342, 32'hc403a1c6, 32'h4414020a},
  {32'h44e957a5, 32'h4374c2f6, 32'h4426cd0f},
  {32'hc2c1c444, 32'hc49b0d67, 32'hc47f0936},
  {32'h450b0787, 32'h439864f5, 32'hc3f9134a},
  {32'h44f7dfde, 32'h435fa314, 32'h43ae106f},
  {32'h4391cab8, 32'h4496cc18, 32'h441fcbb9},
  {32'h434b4ceb, 32'hc4ec69c0, 32'hc45124e9},
  {32'h449bffe7, 32'h41507306, 32'h42963d48},
  {32'hc1b376b3, 32'hc36654fc, 32'hc553f317},
  {32'h450b4203, 32'h43711c8d, 32'hc2ce979c},
  {32'hc4bcf1d9, 32'hc415e4f9, 32'hc48ba04f},
  {32'h4531b5f0, 32'h438cb207, 32'h44186d45},
  {32'hc53d2edb, 32'h4357152b, 32'hc31c2466},
  {32'hc4173d46, 32'hc3526e3b, 32'hc20d904d},
  {32'hc47e40cc, 32'hc451f96f, 32'hc4616066},
  {32'h42379c99, 32'h451b8b78, 32'hc32ac463},
  {32'h421ae2f8, 32'hc47e27fb, 32'h4378b533},
  {32'h44ce0e91, 32'h43a6445b, 32'h4489365e},
  {32'hc4459a68, 32'hc4c9dec3, 32'h42df19f7},
  {32'h4383591e, 32'hc35e3ca9, 32'h4401eeff},
  {32'hc34f75c0, 32'hc3aa9c18, 32'h438396d9},
  {32'hc445dbc7, 32'hc493364a, 32'hc3e68dae},
  {32'h4511c6bb, 32'h43d99c77, 32'h4393ce58},
  {32'hc51675b9, 32'h43512144, 32'h4337d809},
  {32'h451e23b4, 32'hc365f431, 32'h4376b240},
  {32'hc44c9aa5, 32'hc4aabe35, 32'h42d4b8a3},
  {32'h438511fc, 32'h445a6535, 32'h435a03e0},
  {32'hc4821023, 32'hc45a657a, 32'hc45a4628},
  {32'h45049773, 32'h43d6f88a, 32'h43b444ba},
  {32'h42f47656, 32'hc3bd1bd8, 32'h444ef42a},
  {32'h4430e5b9, 32'h44db306f, 32'h43565db2},
  {32'hc4ef55e5, 32'hc1f39378, 32'hc3913cff},
  {32'hc3d86758, 32'h43366ca6, 32'hc4a991cc},
  {32'hc51bbf2f, 32'hc3f6e7ee, 32'hc1af3c7e},
  {32'h43e3dcef, 32'h44102f3b, 32'hc39b0cdb},
  {32'hc52f5c4f, 32'hc2a8b58a, 32'h43b87a2e},
  {32'h448822ee, 32'h445a09c6, 32'h44024a61},
  {32'hc488c550, 32'h4384ad0f, 32'h43335a1b},
  {32'h44899ff8, 32'h43c87f8a, 32'hc262a2e8},
  {32'hc48e8a4a, 32'hc49a1b65, 32'hc489dd99},
  {32'h4387c8cb, 32'h45347341, 32'hc39d98ef},
  {32'h44725b71, 32'h43823ea3, 32'h43795703},
  {32'h43d767af, 32'h448fdca5, 32'hc2c644a3},
  {32'hc2c23ed4, 32'hc3b254ea, 32'h44b78c53},
  {32'h4481ab97, 32'h4402eae6, 32'hc3b7b637},
  {32'hc4b37d08, 32'h434d905a, 32'h4515f38d},
  {32'h44b67d58, 32'hc390ea3a, 32'hc4afb831},
  {32'h42ccc2d0, 32'hc51aa444, 32'h40c79a9e},
  {32'hc3d47bc2, 32'h441f371c, 32'h4454bfa3},
  {32'h4457e644, 32'h43827217, 32'h41f5952e},
  {32'hc50f1795, 32'h43a4362e, 32'hc1856c49},
  {32'h44bc4122, 32'hc424c947, 32'hc2dbdb20},
  {32'hc500ebc1, 32'hc3c24187, 32'hc3b09e1b},
  {32'h45001c0e, 32'h4249c1e1, 32'hc31e05e4},
  {32'hc512679c, 32'h441f7f30, 32'h42634690},
  {32'hc37aa380, 32'h435a0f1b, 32'h43608c4d},
  {32'hc3abb8cc, 32'hc3b530b2, 32'h426d8708},
  {32'h43b21a2c, 32'hc5163db9, 32'hc288b715},
  {32'hc3d69b5e, 32'h4449e05b, 32'h42b0edbf},
  {32'h44a1a8ae, 32'h422de733, 32'h41f4d4b3},
  {32'hc51a29ce, 32'h432f96d1, 32'hc29fbfc0},
  {32'hc4876336, 32'hc3eb81b0, 32'hc39e9423},
  {32'hc2493da4, 32'hc3b44c64, 32'hc550d61f},
  {32'h44b348d8, 32'h42eb3a22, 32'hc34dc8df},
  {32'hc4f07880, 32'h435f1f52, 32'hc3d6b1d0},
  {32'hc332da50, 32'hc4fd4f2f, 32'h43645516},
  {32'hc54f26db, 32'hc2dff2b5, 32'hc3ac2705},
  {32'hc32c3d26, 32'hc38a8b38, 32'h42f9f722},
  {32'hc27767ba, 32'h453cf1b0, 32'h430303a7},
  {32'h43ddbcfb, 32'hc430c938, 32'h44df3860},
  {32'hc4fb7a9c, 32'h43cb7ed8, 32'hc10440dc},
  {32'h41146300, 32'h3f8effa0, 32'h44d3fbee},
  {32'hc365d143, 32'hc341f33e, 32'hc5416a67},
  {32'h432a0931, 32'hc1930f2c, 32'h443af9ad},
  {32'hc401a4ab, 32'h44490672, 32'hc48f62f3},
  {32'h43cf7de8, 32'hc300b47f, 32'h421f6e18},
  {32'h4474a343, 32'hc43c2f54, 32'hc2d1b73d},
  {32'hc53b3013, 32'h434f8efe, 32'h42e70a45},
  {32'hc2231380, 32'hc41b07d1, 32'h441bd205},
  {32'hc2951ab8, 32'hc1be496f, 32'hc4e2dab4},
  {32'hc4efab07, 32'hc4298bfa, 32'h412adabe},
  {32'hc4898bb6, 32'h44a208cf, 32'hc1a9aa0d},
  {32'h44963b4b, 32'hc3a195d4, 32'h4414f5af},
  {32'h4383c3cc, 32'h44f51fff, 32'h44a80bb1},
  {32'hc1ce2ce0, 32'h442f7c2b, 32'hc4e9da90},
  {32'h433b76c6, 32'h441db10e, 32'h43b80dfd},
  {32'hc49f1c72, 32'hc42c5036, 32'hc2b66045},
  {32'hc40d17a2, 32'hc36815a1, 32'hc4e37f73},
  {32'h44a6a001, 32'h43477d52, 32'h43d243d2},
  {32'h44796f12, 32'hc3f760d5, 32'hc40369a2},
  {32'h43f56842, 32'hc2a5c36e, 32'h429bf48f},
  {32'h43351a08, 32'h44dc11bf, 32'hc3e3c460},
  {32'h450e488a, 32'hc41a7a1e, 32'hc34a647b},
  {32'hc5102c98, 32'hc4836e15, 32'hc3f38c70},
  {32'h4421a148, 32'hc402c53c, 32'h44721f86},
  {32'hc4e6175f, 32'h433731e4, 32'h439505bf},
  {32'h43dc7458, 32'hc4ca14bb, 32'hc4125a88},
  {32'hc52af6e3, 32'h433a44a8, 32'hc2e8375b},
  {32'h450c93e6, 32'h439565d1, 32'h43792551},
  {32'hc3c80db3, 32'h4473cc6f, 32'h426a8be2},
  {32'h4496e1fd, 32'hc4b106c9, 32'h43271247},
  {32'h43ab1996, 32'h41a48719, 32'h44b3853a},
  {32'h450a3582, 32'h43e8ce8b, 32'hc3256fb6},
  {32'h42c294c9, 32'hc499e5f9, 32'h454a92e8},
  {32'h43971652, 32'hc52e8776, 32'h41f8709c},
  {32'h44fc0267, 32'h41ce0470, 32'hc2da3cdb},
  {32'hc332e30c, 32'hc1e14882, 32'h44e98345},
  {32'h450c2de1, 32'h43ab98b9, 32'hc3cb25de},
  {32'hc3bf684f, 32'hc30d4ba2, 32'h44daf92a},
  {32'h43b826fd, 32'h43eb1207, 32'hc499ad61},
  {32'h4338bc97, 32'h44327f32, 32'hc49706dc},
  {32'h432af678, 32'h4412ef7f, 32'h450f5871},
  {32'h4487ae1d, 32'h43318b5a, 32'hc4169e55},
  {32'h44f571be, 32'h442e449f, 32'hc2d78bd1},
  {32'hc3e9f529, 32'hc3d43ecb, 32'h44f9b3a1},
  {32'hc2588adc, 32'h44b4ed9c, 32'hc232dbda},
  {32'h431035ba, 32'hc53000b4, 32'h3f87afc0},
  {32'h452a1c2a, 32'hc1841bfe, 32'hc331f1b7},
  {32'hc4a97285, 32'hc3a4dbff, 32'hc2ba50df},
  {32'h44166a48, 32'hc3d7a722, 32'hc31d14c0},
  {32'hc43a5b68, 32'h43aeed97, 32'h42e84889},
  {32'h44aae76e, 32'h42881872, 32'hc39cce54},
  {32'hc5102531, 32'hc3e839b0, 32'h42e596d2},
  {32'h44c43324, 32'h442a7377, 32'hc3906993},
  {32'h431be0dd, 32'hc4fea48e, 32'h42e2c7e0},
  {32'h452830de, 32'h44203c72, 32'hc3baebf6},
  {32'h41f48fe0, 32'hc575dcde, 32'hc2ad9ec2},
  {32'h44714df4, 32'hc3865788, 32'hc30de1f4},
  {32'hc3a154f2, 32'h44e7de27, 32'h43768fca},
  {32'hc33aa2f0, 32'h441797e0, 32'hc4cf72f6},
  {32'h40c583a0, 32'h44e966a9, 32'h44472d03},
  {32'h44d349ad, 32'h42c2f178, 32'hc39a2068},
  {32'h44af6219, 32'h433390f8, 32'h41dd30fb},
  {32'hc4cbe402, 32'hc4246c02, 32'hc40c053d},
  {32'h4533c3a4, 32'h43d726a6, 32'hc39f8a53},
  {32'hc42cc19c, 32'hc4375509, 32'hc50a8a5c},
  {32'h42a8b0c0, 32'h446f85a3, 32'h45135651},
  {32'h4444f129, 32'hc3dd0be6, 32'hc3f32be1},
  {32'h43f410a8, 32'hc4105eb2, 32'h430bd5db},
  {32'hc3bfb5e0, 32'hc4a90ee3, 32'hc43f7e37},
  {32'hc352d0b3, 32'hc301421e, 32'h44d2f16d},
  {32'hc3e26f3f, 32'h42e21aed, 32'hc511cf16},
  {32'h424d4803, 32'h44103ce8, 32'h44127b94},
  {32'h44a67f7a, 32'hc444e015, 32'hc2ac7c70},
  {32'hc317cbb2, 32'h45110986, 32'h44c151f2},
  {32'hc4ec126e, 32'hc3a2b95a, 32'hc39174a4},
  {32'h44f59722, 32'hc3138da8, 32'h4395f387},
  {32'hc45d1883, 32'hc4fd3a68, 32'hc4146d8f},
  {32'h4393ea20, 32'h44cfeca0, 32'hc120cfa8},
  {32'h44c0111d, 32'hc3614f28, 32'hc1c820ec},
  {32'h4536fae1, 32'hc3c3ded5, 32'hc30db1b9},
  {32'hc4d952b5, 32'hc30ab3fc, 32'h43c3921d},
  {32'h454c1cb2, 32'hc28349a7, 32'h43947fa5},
  {32'hc4faf984, 32'hc29b498d, 32'h41b48153},
  {32'h4507cb9b, 32'hc2e820c5, 32'h42b0bf52},
  {32'h44e30296, 32'hc3c9937b, 32'h43b83098},
  {32'h4394b768, 32'h452840ac, 32'h42d2b6d6},
  {32'hc3781514, 32'hc422479c, 32'hc49b5ff7},
  {32'hc5483b84, 32'h44462baf, 32'h427c1ebd},
  {32'h4547966d, 32'hc2ebd809, 32'h441b661e},
  {32'hc44193e6, 32'h43d484de, 32'h4432b9be},
  {32'h44b17d16, 32'hc38d7bbe, 32'hc428cfaf},
  {32'h433d1d50, 32'h449878c4, 32'h44bffd28},
  {32'hc4e936d2, 32'hc3146401, 32'hc3863d36},
  {32'h44845c41, 32'hc4bd13f6, 32'h452bd009},
  {32'h4317978c, 32'h450d2755, 32'hc4c807df},
  {32'hc3aa37b7, 32'h4452a15f, 32'h430b20e2},
  {32'h444a97fc, 32'hc3d5b7d2, 32'hc3ca1745},
  {32'h436cbfd4, 32'h445abedc, 32'h44bbd98e},
  {32'hc336f36b, 32'h43862851, 32'hc45cf469},
  {32'hc41b0ae0, 32'h44c61b9d, 32'h445e746d},
  {32'h44c6d4be, 32'hc426afd3, 32'hc41cd459},
  {32'hc419f178, 32'h440385fe, 32'h43bc5e27},
  {32'h45180280, 32'hc462d6ff, 32'hc3b88e25},
  {32'hc4594274, 32'h452962b4, 32'h418df76c},
  {32'hc48d19b0, 32'hc31747f0, 32'hc25ef5fa},
  {32'hc3567c90, 32'h44a5d1ed, 32'h43ff0610},
  {32'h44ade3b5, 32'hc51da51c, 32'hc36c2ead},
  {32'hc51dd496, 32'hc2d202d1, 32'h42a482f9},
  {32'h42c06a16, 32'h4481c03f, 32'h43b23df3},
  {32'hc4b98f84, 32'hc1872b7e, 32'h43b17eb4},
  {32'h45026664, 32'h42d77091, 32'hc08542e7},
  {32'h4312193e, 32'h4345d62c, 32'hc27492f0},
  {32'hc500bee9, 32'hc38e582e, 32'hc47845ff},
  {32'h4508ccc9, 32'h43b5f7bc, 32'h4448ec1b},
  {32'h44ab2165, 32'h42a7f206, 32'h43496902},
  {32'h450ad528, 32'hc47d4d3b, 32'hc31583fa},
  {32'hc3e392a2, 32'h44867d2e, 32'h42d392f8},
  {32'h449f0d0a, 32'hc398f812, 32'h434528e8},
  {32'hc305ac46, 32'h45711087, 32'hc366c886},
  {32'h44f0729b, 32'hc4d656d6, 32'h43b23c3e},
  {32'hc4a2e515, 32'h428cb162, 32'hc4124a23},
  {32'h4438edfb, 32'hc44948bc, 32'hc3a99857},
  {32'hc4625afc, 32'h43aa93df, 32'hc5004680},
  {32'h444fe8e0, 32'hc2075b0c, 32'hc3213fe3},
  {32'hc24f43b0, 32'h45063e9d, 32'h4378069a},
  {32'h440f9ea0, 32'hc43247a0, 32'hc416bf4b},
  {32'hc4017928, 32'h44a73e47, 32'h442d7a03},
  {32'h446cebda, 32'hc4c08aa9, 32'hc40b6ab3},
  {32'hc3bef2bb, 32'h4413da1d, 32'h45043e27},
  {32'h44320cd6, 32'hc3abe422, 32'h43a126fa},
  {32'hc472ba6a, 32'h4439e7a8, 32'h43826a94},
  {32'h44922aca, 32'hc24d34a7, 32'hc3e0c932},
  {32'h449d6560, 32'hc2e5f4bb, 32'h44312555},
  {32'h449c3a5a, 32'hc421fe61, 32'hc4124658},
  {32'hc4f531c8, 32'h43f651ec, 32'h43743b03},
  {32'h44a9a257, 32'hc2913a54, 32'hc44f14b4},
  {32'hc4a23744, 32'h443ace27, 32'h43efaf73},
  {32'h450c6f22, 32'hc333732b, 32'hc43ee255},
  {32'hc39b31c0, 32'h4396e6fa, 32'hc2992acd},
  {32'hc4b86b90, 32'hc408bbd2, 32'h44de0a1f},
  {32'hc4891c17, 32'h43b27184, 32'hc2a2deb1},
  {32'hc507b577, 32'hc4797802, 32'hc3e3ae9e},
  {32'h4359b1be, 32'h455abd0b, 32'h4348038a},
  {32'hc522f927, 32'hc39e9e79, 32'hc24e6e9f},
  {32'hc39fb3f0, 32'h454edbc6, 32'hc398e9a3},
  {32'hc33afd4a, 32'hc4da567a, 32'h437d610f},
  {32'h4492c23a, 32'h440ee10d, 32'h436c4ff3},
  {32'hc5217345, 32'hc27578c6, 32'hc34c3a9a},
  {32'h451bc463, 32'h43c5a882, 32'h416a614a},
  {32'hc49649ee, 32'h4295ce15, 32'h421e4929},
  {32'h44a9407e, 32'h442a63d1, 32'h43f958a4},
  {32'hc2b937e4, 32'hc43ac280, 32'hc3de993a},
  {32'h42c0e868, 32'h44248349, 32'hc34927ee},
  {32'hc3f94c83, 32'hc3c22ab8, 32'hc49e26d5},
  {32'h43cb601e, 32'h44181d7c, 32'h45104b37},
  {32'hc2c10db2, 32'hc17c1aa1, 32'hc4152746},
  {32'h43dc33ac, 32'h4371d829, 32'h449003f7},
  {32'hc4a72036, 32'hc42f6f3f, 32'hc46be200},
  {32'h448884f4, 32'h438860ad, 32'hc36e8ba7},
  {32'hc4186ded, 32'hc376c91b, 32'h438a37c1},
  {32'hc391a567, 32'hc273992d, 32'h452b7ebb},
  {32'hc4f449f0, 32'hc31c8d30, 32'h424177fa},
  {32'h44104c90, 32'h44c551fe, 32'h441cf807},
  {32'hc42bf309, 32'hc4a29034, 32'hc4cca2c1},
  {32'h434f5f48, 32'h4411d6fd, 32'h445c5d94},
  {32'hc3d9a518, 32'h44a89109, 32'hc328a896},
  {32'hc509c60e, 32'hc3abba41, 32'hc3ac7eb9},
  {32'h434b0863, 32'h4513e6f1, 32'h4479535f},
  {32'h4339c6da, 32'hc4c05e0f, 32'h42883ad9},
  {32'h42a16d98, 32'h451691bd, 32'hc38bde8d},
  {32'hc469310d, 32'hc5041f32, 32'h42758499},
  {32'hc4613709, 32'h439f16df, 32'hc3b6bfcb},
  {32'hc589e186, 32'h43753489, 32'hc367f209},
  {32'hc3abde30, 32'hc2afd300, 32'hbfd45c78},
  {32'hc528d304, 32'h43aa5506, 32'h442cb247},
  {32'h44bc090c, 32'h428c390c, 32'h4416be04},
  {32'hc50a7fdd, 32'hc3a250d3, 32'h42dccf2c},
  {32'h4502e8a4, 32'h431cffde, 32'h424540bf},
  {32'h42954474, 32'hc243a305, 32'h4563febf},
  {32'h447bdb72, 32'h45215a47, 32'h415ca288},
  {32'hc4c4cd12, 32'hc28e23e6, 32'h423a315a},
  {32'h443c3b5a, 32'hc40e0a0e, 32'hc4c17c3a},
  {32'hc5383626, 32'hc2daf81e, 32'h43d013ca},
  {32'h452fbb3c, 32'hc40c272a, 32'hc35012cd},
  {32'hc3b6c7f4, 32'hc4a9483a, 32'h440c21b5},
  {32'h4409a7f6, 32'h45371108, 32'h4052faee},
  {32'h440516d5, 32'h43415e1b, 32'h438d27f4},
  {32'h43875575, 32'h4412156f, 32'hc41d36b0},
  {32'hc4bc61e2, 32'hc4104459, 32'hc41c7d9a},
  {32'h444e9d9b, 32'h3f5fdc60, 32'hc4792a66},
  {32'hc4afa829, 32'hc293a6ff, 32'h4504e580},
  {32'h45455c00, 32'hc343c5d8, 32'hc485a62b},
  {32'hc37220f4, 32'hc4ed7665, 32'h438dcffd},
  {32'hc533d035, 32'h43bc40cd, 32'h43e86919},
  {32'hc4b13ae1, 32'hc31e7e61, 32'hc2869fed},
  {32'hc3fa2ca0, 32'h452318ae, 32'h43c4af70},
  {32'h44e718d6, 32'hc48f968f, 32'h428eae5c},
  {32'h44b8b2a3, 32'h44290adc, 32'h43d9b07b},
  {32'h450fb2cf, 32'h42b1e8be, 32'hc3a0b1cf},
  {32'hc53905af, 32'h440ac845, 32'hc3962178},
  {32'h44293358, 32'hc45822e2, 32'h43362b10},
  {32'hc3115f17, 32'h44a1b82f, 32'hc452e7ee},
  {32'h44061b57, 32'hc4533005, 32'h450870fa},
  {32'hc4b5721e, 32'hc3a5bbfc, 32'hc3772dde},
  {32'h453cda40, 32'h43c271cc, 32'h43200734},
  {32'hc42feaf6, 32'h42f94201, 32'hc557cdc3},
  {32'hc46743c4, 32'h4409d4d3, 32'h4480063a},
  {32'hc517b9b6, 32'h4351650c, 32'hc459105f},
  {32'hc232e1e0, 32'h4276431f, 32'h4504d2d1},
  {32'hc5041c8f, 32'hc35f3a64, 32'hc2a0c74e},
  {32'hc314fd38, 32'hc4b18720, 32'h44f5db6d},
  {32'hc40ccd5e, 32'h44d3e8f8, 32'hc41be8eb},
  {32'hc43497d2, 32'hc338ac2b, 32'h4397a61c},
  {32'hc49e37d8, 32'h4484316d, 32'h428fc88a},
  {32'h447640db, 32'hc501d762, 32'hc3c69d75},
  {32'hc2d004d8, 32'h44bdb33e, 32'h43bd680b},
  {32'h44b84101, 32'h43ae6b43, 32'h43e92b9a},
  {32'hc3a26531, 32'h4348a4e5, 32'hc4c23b80},
  {32'h4429c980, 32'hc33aeda8, 32'h440293bf},
  {32'h43856aec, 32'hc492a8f5, 32'hc53c5772},
  {32'h438e8150, 32'h42b902d3, 32'h43ecd456},
  {32'hc4d62959, 32'h4424befc, 32'h428240cb},
  {32'h4454b9e6, 32'h441deb1f, 32'hc3ee885b},
  {32'hc2f08ee0, 32'hc51791fe, 32'h43af228e},
  {32'hc504e2ad, 32'h43ca5726, 32'hc30999fb},
  {32'h4500f70e, 32'h4347ab57, 32'h4297755e},
  {32'hc453d557, 32'h44595f04, 32'hc490fa82},
  {32'h44d40c42, 32'hc40beec8, 32'h4422cbea},
  {32'h4213c378, 32'h42d4bb80, 32'h442e337c},
  {32'h433b457f, 32'h438090e3, 32'hc534b465},
  {32'h4376c94c, 32'h43c9e16b, 32'h418dec07},
  {32'h445cd68a, 32'h437ca382, 32'h43d233d5},
  {32'hc4d5b8a0, 32'h441298d8, 32'h429c122d},
  {32'hc42f0672, 32'hc4db69da, 32'h440db9aa},
  {32'hc4a8d629, 32'hc37a010a, 32'hc31a1d7c},
  {32'h44d3f062, 32'h42ff0e32, 32'h440bcbed},
  {32'hc369cbca, 32'hc361651c, 32'hc52c281c},
  {32'hc39d692c, 32'hc43fe956, 32'hc28511fa},
  {32'hc59f5098, 32'hc3559788, 32'hc2cdd6bc},
  {32'h4551ef39, 32'h43e6c689, 32'hc44e5d5f},
  {32'hc42c9e87, 32'h445d4d0b, 32'hc38cc9aa},
  {32'h438a0773, 32'hc3f9094c, 32'hc36651ca},
  {32'hc538bcad, 32'h41c86b0b, 32'h43f80a20},
  {32'hc44ccd56, 32'hc33632d6, 32'h4352a0bc},
  {32'hc46352b6, 32'h451517aa, 32'h42eeca52},
  {32'h421fb1f8, 32'hc55aee9e, 32'h43093b8b},
  {32'h41a6cc68, 32'h4396ff36, 32'h437fa7cc},
  {32'h4436e198, 32'hc48792f6, 32'hc41e5bd1},
  {32'hc3505c8b, 32'hc4d5768a, 32'h44d56b32},
  {32'hc4fdfd1a, 32'h422c57e7, 32'h42ab3118},
  {32'h438ccfc6, 32'h45267ed8, 32'h410cd3e3},
  {32'h448e1575, 32'hc44c4a15, 32'hc349080e},
  {32'h44b9670a, 32'h441bc006, 32'hc4933fbc},
  {32'hc4486291, 32'hc5183f4a, 32'hc183bfb4},
  {32'h453206c1, 32'hc347d453, 32'h44732607},
  {32'h45118fa4, 32'hc2cdef4a, 32'h43e2b2ff},
  {32'hc49786dc, 32'hc4f1823f, 32'h44d8823e},
  {32'h43c8d7b8, 32'hc49b065e, 32'hc4873ddc},
  {32'h4441d149, 32'h422a8cfa, 32'hc31c4ba1},
  {32'hc2ee5d50, 32'hc5197bd6, 32'h423eac67},
  {32'h43909c4a, 32'h422e33f6, 32'hc48c088d},
  {32'hc4b1ac3e, 32'hc40eff9b, 32'h441a375c},
  {32'h43c5cf5e, 32'h449918bb, 32'h420358eb},
  {32'hc4e15afb, 32'hc32aee7a, 32'hc1ffb1cd},
  {32'h4545ece7, 32'hc3be5aaf, 32'h4339525b},
  {32'hc525548f, 32'hc20bd2ab, 32'h4411d214},
  {32'h440e5023, 32'hc199f66d, 32'hc4171ca6},
  {32'hc40ff704, 32'hc5168f26, 32'h43e4de10},
  {32'h43f1416c, 32'h44833bca, 32'hc0dff70c},
  {32'hc4e1fbe5, 32'hc15a3663, 32'hc1ffc038},
  {32'h432ead76, 32'h450b8a93, 32'hc3ff99a8},
  {32'h439471bc, 32'hc56149a2, 32'hc3acbdc2},
  {32'h44b04e42, 32'hc3565e95, 32'hc3340cc4},
  {32'h44946094, 32'hc461b9a9, 32'h42487651},
  {32'hc4884a14, 32'h44108920, 32'hc3f59bd2},
  {32'h44f94f94, 32'h43c359e0, 32'h44088064},
  {32'h4486d347, 32'hc417d87d, 32'hc31780fd},
  {32'h44a471ac, 32'h4384f97f, 32'h4492a410},
  {32'hc4fd4553, 32'hc403466c, 32'h438587db},
  {32'h4504697b, 32'hbf00a5c0, 32'h4380a337},
  {32'hc533eea3, 32'hc30a4c9e, 32'hc1374b1e},
  {32'h44ac2316, 32'h43f2b7a8, 32'h44522893},
  {32'hc332dae4, 32'hc44d0832, 32'h42d33762},
  {32'hc2387e20, 32'hc32dfd1c, 32'h44c3da73},
  {32'hc4846f2e, 32'hc3f9a137, 32'hc3e5c097},
  {32'h4341d422, 32'h44f71740, 32'hc1b0225e},
  {32'h428c3e60, 32'hc4814b22, 32'hc4953bb1},
  {32'h4423961b, 32'h43b90b4e, 32'h44f62f6f},
  {32'h440522f8, 32'h41b663d0, 32'hc453a8c7},
  {32'hc467bae9, 32'h4403d70c, 32'h45417fd4},
  {32'hc32efd10, 32'hc46ef7a3, 32'hc4754856},
  {32'h4380b9c3, 32'h4495ae5e, 32'h43b4af9c},
  {32'hc506dd4c, 32'hc3faef96, 32'hc285f404},
  {32'h43af9694, 32'h4505df67, 32'h41d33918},
  {32'h44fd84c5, 32'hc3800144, 32'hc3c6ad74},
  {32'h453a92b2, 32'h43ad68af, 32'h43eb3534},
  {32'hc525e991, 32'hc18a8bfb, 32'h42cea0d3},
  {32'h44ec9198, 32'h43b248f4, 32'h4406b152},
  {32'hc3a36b44, 32'hc2ce0fbc, 32'h432bbf35},
  {32'h44aef360, 32'hc446505d, 32'h40e0be8a},
  {32'hc3788dc2, 32'h44a4cfd5, 32'hc5159050},
  {32'hc2b11d53, 32'h450c7948, 32'h438386de},
  {32'h448863c0, 32'h43d1d999, 32'h4369525a},
  {32'hc492977d, 32'h43782116, 32'h4427743c},
  {32'hc3a3d5eb, 32'hc41aa3da, 32'hc49c560d},
  {32'h44900d08, 32'hc1677c67, 32'hc360e5e3},
  {32'h4352ae90, 32'hc4692dff, 32'hc4cf2822},
  {32'hc405afae, 32'h44bfa41c, 32'h44ac5011},
  {32'hc4d09181, 32'hc3862203, 32'hc35119de},
  {32'hc3a2317f, 32'hc4890314, 32'h4506092d},
  {32'h44c2c654, 32'h43c957f8, 32'hc3e4b162},
  {32'h442b1cbc, 32'hc3f3c417, 32'h43982611},
  {32'h45063d84, 32'hc2dfc4ae, 32'hc3aaf577},
  {32'hc4992442, 32'h43dcc5c8, 32'h442e6f06},
  {32'h44a68997, 32'h438e67f5, 32'hc386d4d4},
  {32'hc3107ca8, 32'h43347096, 32'h4570f903},
  {32'h439775f8, 32'h41b92770, 32'hc4de25e3},
  {32'hc45ad6f0, 32'h43cf844d, 32'h42ad74e6},
  {32'h45537e56, 32'hc44691ea, 32'hc38af0c8},
  {32'hc52d10e5, 32'h449e83e9, 32'h42b7cdba},
  {32'h447e107a, 32'hc143f1bc, 32'hc2aa8cad},
  {32'hc4c66907, 32'h44a54395, 32'h445bce0d},
  {32'h44af16ae, 32'hc5074473, 32'hc14a6358},
  {32'h449b267d, 32'h439caa34, 32'hc2afb6ef},
  {32'hc3ae1d68, 32'hc3aceb25, 32'hc3ee23e6},
  {32'hc5891ec8, 32'h436d7ad1, 32'h42df265a},
  {32'h452e7eb2, 32'h42b43038, 32'hc312126e},
  {32'h44d6ffcc, 32'h42b2a1f0, 32'h43cf85c1},
  {32'hc4d92081, 32'h42cf2f73, 32'hc3da3449},
  {32'hc1447f00, 32'hc3cd644f, 32'h4529202c},
  {32'hc259249e, 32'h450c3807, 32'hc3fbceea},
  {32'h42659f10, 32'hc2f0aeac, 32'h443379d4},
  {32'hc3d9e625, 32'h454797a2, 32'h43b8a928},
  {32'hc4ac4751, 32'hc3f64ee0, 32'h434243de},
  {32'hc421bc2a, 32'h4498041a, 32'h44293b69},
  {32'h4432133c, 32'hc5182f37, 32'h42c93328},
  {32'hc49aa111, 32'hc31c8cf6, 32'h428e78e1},
  {32'h4521f0da, 32'hc370ddcf, 32'hc2ac2934},
  {32'hc5384ae8, 32'h4396f2b2, 32'h43a85df7},
  {32'h45060056, 32'h434d0122, 32'h440b8352},
  {32'hc025f500, 32'h445086c6, 32'h451e807d},
  {32'h43feb736, 32'hc4c52be0, 32'hc40e915a},
  {32'hc43c4bc0, 32'h4445f3b4, 32'h441e856a},
  {32'hc290cbf6, 32'hc3d4fb7f, 32'hc4f4908f},
  {32'hc414a3bf, 32'h442aa493, 32'h44ba2042},
  {32'h453f1b3e, 32'h41925f88, 32'hc27eac2c},
  {32'hc4d91e9c, 32'h428a916e, 32'h44919106},
  {32'h431c0d57, 32'hc4812708, 32'hc4e2f074},
  {32'hc5294f16, 32'hc335d090, 32'hc3224503},
  {32'h450ffeda, 32'hc41a9ab4, 32'hc3fa79bd},
  {32'h430ca5fa, 32'h43a6c1af, 32'h4509edb4},
  {32'hc4156f1c, 32'hc42d6938, 32'hc400e1a3},
  {32'hc44c38f8, 32'h442d1742, 32'h44788e59},
  {32'h44c2b428, 32'hc465db05, 32'hc3c67ff4},
  {32'h451e1864, 32'h433ace95, 32'hc433271f},
  {32'hc56d1d0e, 32'h42d4d6e7, 32'h43399c9b},
  {32'hc3c31816, 32'h43bd9d67, 32'h43093639},
  {32'h42ac96c8, 32'hc510c249, 32'hc412b675},
  {32'h4475db48, 32'h449f6d07, 32'h43d24eee},
  {32'h45049e4e, 32'hc39d86d0, 32'hc2a850a9},
  {32'h4514486e, 32'h448ad36d, 32'hc3431eca},
  {32'hc35feda4, 32'hc57a4a18, 32'h43b56e95},
  {32'h425271bc, 32'h438ecba5, 32'hc2733fce},
  {32'hc4e0632e, 32'hc304a88d, 32'hc1f92331},
  {32'h43f02208, 32'h423668e4, 32'h439a6175},
  {32'hc4090d0f, 32'h43ace7d4, 32'h44307d1e},
  {32'h448f87ca, 32'h4400a66a, 32'h44986439},
  {32'hc3d70bf2, 32'hc42d0942, 32'hc45988d7},
  {32'hc482c16f, 32'hc27af9e0, 32'h438ba48d},
  {32'hc4f36331, 32'hc2ed441e, 32'hc46b08d3},
  {32'h43e4c44c, 32'h44202e88, 32'h44e23119},
  {32'hc485e4b4, 32'hc48ffeb1, 32'hc3d70193},
  {32'h4318b8e4, 32'hc42c19cb, 32'h446cd472},
  {32'hc540cb4b, 32'hc3b802e6, 32'hc3fbff48},
  {32'h45540c14, 32'h41a8afde, 32'hc3dbfdc7},
  {32'hc3f9c0da, 32'h40f612ee, 32'hc4d601a7},
  {32'h44de4982, 32'h43a6801a, 32'hc271e94c},
  {32'hc2dc6610, 32'hc387d5ac, 32'hc44e6f98},
  {32'h443623a8, 32'h44af722d, 32'h413a7e4e},
  {32'hc408a1e4, 32'hc48c3428, 32'hc4f62736},
  {32'h42883658, 32'hc3aa9477, 32'h4299bdad},
  {32'hc4c6f8b0, 32'hc36bf760, 32'h430f29f8},
  {32'h41d77380, 32'hc5312c32, 32'hc3972030},
  {32'h44825428, 32'h4471826c, 32'h4370f12e},
  {32'hc3b4b307, 32'hc35b06cd, 32'hc1e72b4c},
  {32'h444a1d7d, 32'h44f20fd9, 32'hc3965407},
  {32'hc4678a49, 32'hc5022d31, 32'h433e3d85},
  {32'h45468a80, 32'hc3a0f35e, 32'hc3d95e53},
  {32'hc4f0e39c, 32'h438290e9, 32'hc35b5be0},
  {32'h44e5bd84, 32'h43afbb02, 32'h44913929},
  {32'hc4a492d0, 32'hc2c65746, 32'hc384cee3},
  {32'h43e06d72, 32'h44b09c8a, 32'hc2bc2346},
  {32'hc448e57a, 32'hc400ff98, 32'hbea5c2d8},
  {32'hc384d105, 32'h446ba4cb, 32'hc42c9a1c},
  {32'hc514c7dd, 32'hc3d45712, 32'h43938704},
  {32'hc3873308, 32'h41d13538, 32'hc512f42c},
  {32'h436bcd06, 32'hc39fb793, 32'h44e9f5d8},
  {32'h451f967b, 32'hc3113fff, 32'h4302d8ce},
  {32'hc43f79ae, 32'h429f72f2, 32'h44fe1b3e},
  {32'hc4f10e7e, 32'h440e1b00, 32'h4281a32c},
  {32'hc403878c, 32'hc53c4cee, 32'h4400c817},
  {32'h441ae683, 32'h43c2f977, 32'hc469dbcb},
  {32'h444cf1e9, 32'hc4239c07, 32'h43870b53},
  {32'h44eed00c, 32'h43899b5b, 32'hc3101475},
  {32'hc3e7d0ab, 32'hc51af7ab, 32'hc4182009},
  {32'h43979ac8, 32'hc3853fae, 32'hc51bbb96},
  {32'hc49427a5, 32'hc29d7f67, 32'h449d3f29},
  {32'h456a43ba, 32'h425557de, 32'hc432f19c},
  {32'h44fc5383, 32'hc4444a2f, 32'hc28d3c15},
  {32'hc5834027, 32'h41818a93, 32'hc25e8b02},
  {32'h450b234c, 32'h429bc2e8, 32'hc1d749f0},
  {32'h43a69c68, 32'h44aea5c5, 32'hc3a925d4},
  {32'h451b7e78, 32'hc3bfde60, 32'hc3a44f04},
  {32'h434824ce, 32'h45260451, 32'h433bdd1d},
  {32'h4527c61d, 32'h4448bc46, 32'h4323b65a},
  {32'hc5247f55, 32'h43f76cd0, 32'h439bc8bb},
  {32'hc45a8fae, 32'hc30a6abe, 32'h42eaf2d0},
  {32'h427cb300, 32'h4530d5f7, 32'h43749fc4},
  {32'h445096db, 32'hc4acd3f0, 32'h44a48d00},
  {32'hc38916b2, 32'h44d0f516, 32'h4232b8a5},
  {32'h44180db0, 32'hc4ab2fc9, 32'hc191297c},
  {32'hc4235b81, 32'hc29d5740, 32'hc4f7bff4},
  {32'hc46be23b, 32'h43eedab8, 32'h446343ec},
  {32'hc4759c3c, 32'h4324f9c8, 32'h438a16ab},
  {32'h43bf715c, 32'h42f76470, 32'h4310158c},
  {32'h450ce652, 32'hc3ca2fca, 32'hc39ea59b},
  {32'h4411c86e, 32'hc4d350fd, 32'h41836eb6},
  {32'hc4b5f243, 32'h449523b3, 32'hc46f68be},
  {32'h44204d6c, 32'hc3e8b5c3, 32'hc2034eea},
  {32'hc3ba8ed0, 32'h44c17673, 32'hc3ae69ec},
  {32'h451f4c41, 32'h43b38cb7, 32'hc3b65154},
  {32'h4484aa85, 32'hc24b3970, 32'h4357cebc},
  {32'h44b6a998, 32'h41ce97ef, 32'h445b6e3a},
  {32'hc4fa6269, 32'hc3d3cf83, 32'hc4ab87b4},
  {32'h448c7954, 32'hc2f52485, 32'hc3188903},
  {32'h435ba838, 32'hc443e989, 32'hc56a250e},
  {32'hc35d3d38, 32'hc43921ad, 32'h4543b169},
  {32'hc4a472fd, 32'h4378daae, 32'hc3be2560},
  {32'hc4d5e4b9, 32'h43bcf1cd, 32'hc30e0b64},
  {32'h443fbe90, 32'hc52d8aac, 32'hc3ea2db9},
  {32'h4257c540, 32'h4352f6ba, 32'hc457cb5d},
  {32'h43a5ef34, 32'hc3ffcc28, 32'h446c33e6},
  {32'hc4669f39, 32'h44f07eb8, 32'hc3be6c4b},
  {32'h415f20c0, 32'hc319e4ff, 32'h451016dd},
  {32'hc381e24c, 32'hc4ee3f26, 32'h45113e71},
  {32'hc487d41c, 32'h44b19a8c, 32'hc47a241c},
  {32'h44a4980d, 32'h437929fa, 32'hc3a68253},
  {32'hc3030308, 32'h435ad299, 32'h43fcaac6},
  {32'hc3b85c9e, 32'h4350bad9, 32'hc4439312},
  {32'h44c7b054, 32'hc42e1f7a, 32'h42c69abb},
  {32'h450cd23e, 32'h435840af, 32'hc321c95c},
  {32'h433011b8, 32'hc50330fa, 32'hc2f7ebec},
  {32'h441d7498, 32'h450ad6d1, 32'hc30d0023},
  {32'h443f2872, 32'h430d5b03, 32'h43b2a4a9},
  {32'hc496400d, 32'h43c071e1, 32'hc436624c},
  {32'h450782eb, 32'hc3a1e695, 32'h44741821},
  {32'hc28bab5a, 32'h44f4a782, 32'h43213594},
  {32'h4519f6b4, 32'hc43b25e8, 32'h43dca2fd},
  {32'hc51319f9, 32'h445bbab2, 32'h42c9fb0a},
  {32'hc4122ff5, 32'hc4097a85, 32'hc31fcec8},
  {32'h434a8578, 32'h452816fc, 32'hc37da80c},
  {32'h44da3d26, 32'hc4bcb515, 32'hc2a7cec0},
  {32'hc44c9dbf, 32'h446702e0, 32'hc218de87},
  {32'hc3afc1b1, 32'hc494b847, 32'hc48b0307},
  {32'h4445a053, 32'hc3a2fd6b, 32'h45217a11},
  {32'hc2fe7726, 32'hc56823d2, 32'hc331e71b},
  {32'h445b2640, 32'h44b6b70b, 32'h430644bd},
  {32'hc1b35580, 32'hc461fe5a, 32'hc2954143},
  {32'h4462c744, 32'h41ea1ff2, 32'hc46dfc0c},
  {32'hc20d9f54, 32'hc4c1c2c5, 32'h4319c160},
  {32'h450eabfc, 32'hc18293b6, 32'hc3abdf92},
  {32'h44397d35, 32'h44180c06, 32'hc4ddc57f},
  {32'hc3301dd0, 32'h45080516, 32'h44d27b70},
  {32'h448d4d5a, 32'hc425f8d5, 32'hc4ac7788},
  {32'h438a3d16, 32'hc260acbd, 32'hc4d79824},
  {32'hc42b0e77, 32'hc442eb9b, 32'h43de12eb},
  {32'hc40e4793, 32'h44838f3a, 32'hc3a5b996},
  {32'hc44e8e00, 32'hc40a96b3, 32'h44f07314},
  {32'h42e32fca, 32'h44605615, 32'hc4dcd0a5},
  {32'hc3092db0, 32'hc3801966, 32'h448bb688},
  {32'h45366f25, 32'hc2b1dd3b, 32'hc3084cf7},
  {32'hc51dc176, 32'hc3aee2a4, 32'hc1e416a1},
  {32'h450624e7, 32'h43e5917e, 32'h4265db20},
  {32'hc41f5524, 32'hc4ce876f, 32'h432aaf63},
  {32'h43559c7c, 32'h43d8e457, 32'h43ad6e08},
  {32'hc39a926c, 32'hc3a17d13, 32'h43d2771c},
  {32'h4505a23c, 32'h44169ea3, 32'hc39fcca4},
  {32'h421cad42, 32'hc54c0139, 32'h433e2e19},
  {32'h42cec600, 32'h4482a52d, 32'h4377b4cc},
  {32'h439a6ecf, 32'hc48e3575, 32'h43d69d42},
  {32'hc437ed7f, 32'h4520cd38, 32'hc4b73d53},
  {32'hc315f0ab, 32'hc40c10c7, 32'h45031d51},
  {32'hc461c903, 32'h43cbf919, 32'h42a10dc9},
  {32'h4534f230, 32'h424c1a61, 32'h444e7ccb},
  {32'hc361d538, 32'hc4f3612d, 32'hc389283a},
  {32'hc3b00ee5, 32'h43d94ec9, 32'h43be0943},
  {32'hc382496e, 32'hc2dd032d, 32'hc5458eaf},
  {32'h43e7bb27, 32'h4456b523, 32'h4518816c},
  {32'hc4a6d91e, 32'hc416b120, 32'h43816523},
  {32'h43726d2e, 32'h45248d56, 32'h443fbda3},
  {32'h431b653b, 32'h40e2dc90, 32'hc4567a24},
  {32'h43f942ff, 32'h400e2585, 32'h44e07fd8},
  {32'hc33138a4, 32'hc4923121, 32'hc47e4a51},
  {32'h4490179c, 32'h444bfbae, 32'h443f97d7},
  {32'h44932acc, 32'h428f0600, 32'h430c06cd},
  {32'h4434a9f4, 32'h44b952ef, 32'h4434c236},
  {32'hc4fbff6f, 32'hc3b0715d, 32'hc42f7347},
  {32'h4441dbb1, 32'h43aaa799, 32'h43c64fcd},
  {32'hc2d09308, 32'hc5173446, 32'hc311364d},
  {32'h42b15132, 32'h452d1e28, 32'h44428eca},
  {32'hc4f1d0da, 32'h4241c9fd, 32'hc39151ac},
  {32'hc439be0a, 32'h4575d815, 32'h41ae1eea},
  {32'hc4571249, 32'hc41d0e23, 32'hc2794480},
  {32'h4516224c, 32'h43935d34, 32'h44275c54},
  {32'hc444bb2f, 32'h44843d57, 32'h43ebc968},
  {32'h44b3140a, 32'hc37ad0cc, 32'h43c6d26f},
  {32'h42c33acc, 32'h45051e6d, 32'hc4953248},
  {32'h4295ae7c, 32'hc4a3e191, 32'h44e51eb7},
  {32'h439916a4, 32'hc4df9a0b, 32'hc2389b37},
  {32'hc4aae7b0, 32'h44b7579d, 32'h439e3abb},
  {32'hc330f854, 32'hc415b61a, 32'hc44333af},
  {32'h4431e527, 32'h44cb34de, 32'hc3778f20},
  {32'h43a8a01a, 32'hc51c7660, 32'hc4f238d4},
  {32'hc307f250, 32'h40915108, 32'h44dd755c},
  {32'h4418015a, 32'hc47b25a3, 32'hc30847de},
  {32'h43a49562, 32'h44c711f1, 32'h43c3fcad},
  {32'h43d5cf2a, 32'hc468fb4e, 32'hc448e4f3},
  {32'h43b916ec, 32'h4512f9a4, 32'hc34a4d98},
  {32'h43e07a40, 32'hc4077783, 32'hc3ace2fe},
  {32'hc4b71f67, 32'h44942ecd, 32'hc04ef035},
  {32'hc3a9ad99, 32'hc40b4584, 32'hc4543689},
  {32'hc411ff16, 32'h44111d63, 32'h44fbb907},
  {32'h4445ca9c, 32'hc460b5a8, 32'hc3d313c4},
  {32'hc50b5574, 32'h428636a1, 32'h4141164c},
  {32'hc3808257, 32'hc497314f, 32'hc3f69459},
  {32'hc4b27851, 32'h4461c524, 32'h434b62a5},
  {32'hc49c6f80, 32'h42ad1775, 32'h408dd196},
  {32'hc55174ce, 32'h431c73ad, 32'hc34b0634},
  {32'h438f9308, 32'hc4fa5121, 32'h43bbd88f},
  {32'h4508dda6, 32'hc2aa4cbb, 32'hc386bb8a},
  {32'h42b867ea, 32'h44478179, 32'hc35a8f51},
  {32'hc5797ba5, 32'h433666be, 32'hc41651cc},
  {32'hc414d357, 32'hc3c917a2, 32'h4168d6fc},
  {32'h44eb9f3c, 32'hc3439849, 32'hc40fae65},
  {32'hc475a83c, 32'h434737f2, 32'hc50efcb7},
  {32'h4525e50f, 32'h4377c6af, 32'h42ae9858},
  {32'h44a84a94, 32'h438b1770, 32'h43131ff0},
  {32'h44cc4e74, 32'hc3b50c8f, 32'h43104929},
  {32'hc4c73ff6, 32'h43b7822c, 32'hc2c51e99},
  {32'hc34298f4, 32'h43f16d81, 32'hc3e7fbf5},
  {32'hc545e0b1, 32'h4312d782, 32'h434f5b06},
  {32'h44cdb282, 32'hc45666c4, 32'h4464576d},
  {32'h42f34fe4, 32'hc36801e9, 32'hc489bd13},
  {32'h443c7009, 32'h447fad18, 32'h44e03a1e},
  {32'hc3d1d499, 32'h437d7caa, 32'h438fd4ad},
  {32'h440508b7, 32'hc22658f1, 32'hc4326d13},
  {32'h43cc7284, 32'hc2055d12, 32'h45180b97},
  {32'h44650179, 32'hc316b158, 32'hc41140a9},
  {32'hc39d86cf, 32'h42c20856, 32'h4427ca25},
  {32'h42f16f17, 32'hc519a45d, 32'h42932e48},
  {32'hc4dbc8f0, 32'h437c66a5, 32'hc37d7dac},
  {32'h454d2f39, 32'hc2f0a348, 32'hc0ba706c},
  {32'hc4db2a16, 32'hc4427c64, 32'h441c74a3},
  {32'h44a22b9a, 32'h438a7ca0, 32'hc4a08f08},
  {32'hc3bc3be6, 32'h42b027e7, 32'hc222e832},
  {32'h44ad4c6f, 32'hc40a23c8, 32'hc3e2d8aa},
  {32'hc34d85a5, 32'h4395ed9c, 32'h441eac16},
  {32'h43e6b206, 32'h42ee060f, 32'hc2f28c9a},
  {32'hc41a4844, 32'h450dd65a, 32'h4409d5d5},
  {32'h42e9c9c0, 32'hc51c7523, 32'hc4184101},
  {32'h450ecb5b, 32'h43b66274, 32'hc3dc44f8},
  {32'hc50abdde, 32'h42fc33dc, 32'h448b8e26},
  {32'h453505fb, 32'hc358334b, 32'h43de10a0},
  {32'hc4def596, 32'hc413de75, 32'hc47bc1b8},
  {32'hc3966611, 32'h453e06ee, 32'hc30512de},
  {32'h43e76228, 32'h41c6717e, 32'h418ad44a},
  {32'h44dc0350, 32'h44a37a66, 32'hc3289222},
  {32'hc5529ef9, 32'hc35478b9, 32'h43ac17e3},
  {32'hc4de6ebd, 32'h424b89fc, 32'h43a9cfa3},
  {32'h42e09410, 32'hc157347f, 32'h446fc050},
  {32'h43e36778, 32'hc40efda1, 32'hc4dd406c},
  {32'hc408e0e3, 32'hc28b9301, 32'h43abe3f8},
  {32'h445bd0da, 32'hc2807ba8, 32'h44ea74f6},
  {32'hc3854934, 32'h42e97d9c, 32'hc5125f84},
  {32'hc476b7ce, 32'h4286828a, 32'h43cffea2},
  {32'hc545b030, 32'hc3583428, 32'hc290ef79},
  {32'h43242106, 32'h44801176, 32'h441c6544},
  {32'h4337cc0a, 32'hc307d9c4, 32'hc4bbbb84},
  {32'h4583e14f, 32'hc418264b, 32'h43f62d57},
  {32'hc432e780, 32'h43c59c2d, 32'hc4704030},
  {32'hc42c4078, 32'hc1f5a3ec, 32'hc39a2767},
  {32'hc26ba0c0, 32'hc47cba07, 32'hc4ccb1a5},
  {32'h44b0004d, 32'h3d986bb0, 32'h4419c1b3},
  {32'h44791d62, 32'h435cf612, 32'hc42f9f35},
  {32'hc39e067b, 32'h43073e88, 32'h4503d050},
  {32'hc408b110, 32'hc1ae536c, 32'hc4f37513},
  {32'h448036aa, 32'hc2d83690, 32'h449e10d7},
  {32'h44e24c23, 32'hc2db0011, 32'hc3937bf0},
  {32'hc55ad922, 32'hc3743a95, 32'h43032511},
  {32'h44de28b2, 32'h447a29f4, 32'hc36a8804},
  {32'h44e671c3, 32'hc28a2e54, 32'h4305d469},
  {32'h45169189, 32'hc33d3684, 32'hc3d9f7ab},
  {32'hc524ba13, 32'hc416a5aa, 32'h43b7b04f},
  {32'h44df8895, 32'h43fc7578, 32'hc38c7a91},
  {32'hc4f2bab1, 32'hc41853ad, 32'hc4139329},
  {32'h4543bda4, 32'hc376be7a, 32'h43232da5},
  {32'hc459ad66, 32'hc2b6e866, 32'h4352d2d8},
  {32'h44a6ecb5, 32'h4401b6e8, 32'hc4bdcfc2},
  {32'hc4a34511, 32'hc46ee20e, 32'h440e426c},
  {32'h421fafe0, 32'h42df762d, 32'hc3b5d6e5},
  {32'hc5294656, 32'h44013013, 32'hc247b621},
  {32'h4405a2c1, 32'h45016e2d, 32'hc2e2fbe9},
  {32'h439aad3c, 32'hc3265cdd, 32'hc2b2e2fc},
  {32'h433954c0, 32'h43294378, 32'hc5023c09},
  {32'hc3f5594c, 32'h43bdf5a1, 32'h4502390e},
  {32'h43cdf53b, 32'hc2e42af4, 32'hc4be565b},
  {32'hc55e4ff0, 32'h432efe01, 32'h42ca5c69},
  {32'h441f4714, 32'h452834c6, 32'hc25439f4},
  {32'h44ac0e16, 32'hc32a9214, 32'hc2c0156e},
  {32'h44047c8a, 32'h43d1487d, 32'hc4d57552},
  {32'hc4e4853d, 32'hc392c51b, 32'h4473423d},
  {32'hc43fa381, 32'h4031ab90, 32'hc4850e29},
  {32'hc4ccc433, 32'h4322ffff, 32'h4525c412},
  {32'h439f5f29, 32'hc40c64ca, 32'hc538cc76},
  {32'h4493c866, 32'hc4a00d68, 32'hc3063836},
  {32'hc4eb4c1e, 32'h432da1d9, 32'hc2f9793f},
  {32'h442e9c2e, 32'hc3c9e6c9, 32'hc3cb759f},
  {32'hc2e34120, 32'h45119788, 32'h43a3330f},
  {32'h4422121b, 32'h43c67f65, 32'h43c12d87},
  {32'h43e3bc53, 32'h44addd2a, 32'h42f5eb9d},
  {32'h45758583, 32'hc4003393, 32'hc4000fde},
  {32'hc4ffb068, 32'h43a96215, 32'h439da1b2},
  {32'h4477ed6e, 32'hc47265d3, 32'hc401c784},
  {32'hc3a784f6, 32'h4465a0ff, 32'hc517db19},
  {32'h44b20100, 32'hc40247a1, 32'h43b0d308},
  {32'hc3a65d86, 32'h436b7921, 32'hc4ab95c1},
  {32'h4388683e, 32'hc42f3260, 32'hc2e99dc1},
  {32'hc42a9eba, 32'h437a931e, 32'hc4a1a608},
  {32'h4502a5fc, 32'h4338fd3f, 32'h433be25d},
  {32'hc36aa2c8, 32'h42c7aad8, 32'hc46c291b},
  {32'hc3b452d7, 32'h444ad1e2, 32'h457e004f},
  {32'h44e59b3d, 32'h43e65cf7, 32'hc3f51d01},
  {32'h4519c4ab, 32'hc2a209f0, 32'h435162da},
  {32'hc53c2932, 32'hc22a2804, 32'h43da4f5d},
  {32'hc3b83a71, 32'hc46927cd, 32'hc30cdb7f},
  {32'hc332b428, 32'h44829592, 32'hc3a6913b},
  {32'h44571a9d, 32'hc3fedbb4, 32'h44322b93},
  {32'hc50b322b, 32'h437958db, 32'hc2fcc233},
  {32'h455216b6, 32'h432c8d6d, 32'h44014b81},
  {32'hc414b620, 32'h43c3b7c1, 32'hc422be6d},
  {32'h44143cf9, 32'hc3d452ac, 32'h44ea03de},
  {32'hc3aa4bcc, 32'hc38b3e90, 32'hc5042c10},
  {32'hc2cd8669, 32'h43fce986, 32'h44736f3b},
  {32'hc2e6fb2c, 32'h43ae5635, 32'hc48aa708},
  {32'hc4843cbc, 32'h429710c0, 32'h43891964},
  {32'h44c18669, 32'hc351cff3, 32'h44be2820},
  {32'hc53190c5, 32'h40b6902f, 32'hc39a317f},
  {32'h44c79603, 32'h43ce645e, 32'h43d4ecf0},
  {32'hc44a21ed, 32'h443cdd77, 32'hc503c056},
  {32'h444230a5, 32'hc493056b, 32'h4424c1fc},
  {32'h43267df0, 32'h44c3c2ff, 32'h44a70d70},
  {32'hc05d4dc0, 32'h4419d07e, 32'hc4e269c3},
  {32'h43a51576, 32'h44644171, 32'h41801279},
  {32'hc4e725ac, 32'hc38d5f0f, 32'hc435ea5a},
  {32'hc46c6808, 32'h4401edb7, 32'hc2938b3b},
  {32'hc3f7a2c7, 32'hc39dbb78, 32'h44a4fefd},
  {32'hc53715e4, 32'hc3610885, 32'h43a6bf80},
  {32'h4498bff5, 32'hc4556a15, 32'h443f80e0},
  {32'hc3d61944, 32'h443a100c, 32'hc4cb7dd8},
  {32'hc46d18bd, 32'hc4172412, 32'hc38f81b1},
  {32'hc47045c0, 32'h40335ed0, 32'h436ec649},
  {32'h44b0ffbe, 32'hc323eeed, 32'h436bdd75},
  {32'h44f9757e, 32'hc1acf805, 32'hc387fbb5},
  {32'h45345dbc, 32'h43ce7b26, 32'h431c2abb},
  {32'hc49955ce, 32'h43d43f08, 32'h42d3934d},
  {32'h44af378d, 32'h421b1bd8, 32'h43c4300d},
  {32'hc4367066, 32'h45139009, 32'hc43c3c02},
  {32'h4497df6e, 32'hc4988864, 32'h430d8260},
  {32'hc34be938, 32'h440f5b98, 32'hc27a8417},
  {32'hc449d6a6, 32'hc4ddc302, 32'hc50f38d9},
  {32'hc429985a, 32'hc49c4006, 32'h44b33cc5},
  {32'hc2ecf920, 32'h4310d577, 32'h451b016d},
  {32'h43a08652, 32'hc2c9dfcb, 32'hc48c6465},
  {32'h44937c4e, 32'hc2805008, 32'h4463182f},
  {32'h442787af, 32'h44a5eba7, 32'hc42a0a55},
  {32'hc4621a3b, 32'h438fd329, 32'h4501c2ea},
  {32'hc2d7773f, 32'h4498706b, 32'hc321b8d6},
  {32'hc2c299ec, 32'hc38a925e, 32'hc2a2b5ea},
  {32'hc3e44088, 32'hc49d2109, 32'h44ee867a},
  {32'h423887ce, 32'h44560d84, 32'hc50d1caa},
  {32'h4404c9b9, 32'h43e827da, 32'hc1d07a55},
  {32'hc29426f1, 32'hc3b38b86, 32'h4540ecb2},
  {32'hc3ebbe7f, 32'h44d29c69, 32'h4391874b},
  {32'hc51e6ae5, 32'hc3ed91e0, 32'h442202db},
  {32'h44d8a6cc, 32'h42483929, 32'h43903fb5},
  {32'h44a09ed5, 32'h4339fc64, 32'h441ea455},
  {32'h441954a0, 32'h4408bdea, 32'h435a5767},
  {32'hc506ac57, 32'h4438d8ec, 32'hc3c318b1},
  {32'h42e1ca7d, 32'h43c2d17d, 32'hc2e743c9},
  {32'hc382f7d4, 32'hc54f14df, 32'h44165378},
  {32'h440546bf, 32'h43c70874, 32'hc1eb0112},
  {32'hc4869ea0, 32'hc3ba04fd, 32'h432a91a2},
  {32'h4517165b, 32'h44451a04, 32'h43035c2f},
  {32'h43155f3f, 32'hc53fad7c, 32'hc1812c0e},
  {32'h4302d618, 32'h443a832c, 32'hc20b9e8c},
  {32'hc33b3d3e, 32'h4475ee8e, 32'hc33efd48},
  {32'hc3d5010c, 32'hc50b3446, 32'h424054e1},
  {32'h42ea6e90, 32'h44e6515e, 32'h446e4345},
  {32'h4395bcd2, 32'h424bd2e1, 32'h422d8a6a},
  {32'h421d787c, 32'h43456bc3, 32'h453d0c43},
  {32'hc4430e0b, 32'hc4977bc6, 32'hc3d75619},
  {32'h45022d76, 32'hc30189ef, 32'h43450883},
  {32'hc531a401, 32'hc42749c2, 32'hc459b898},
  {32'hc16cb340, 32'h450398a6, 32'h44f6c5e2},
  {32'h442cde61, 32'h42b5ae5a, 32'h42b9e805},
  {32'hc49e09b5, 32'hc5016650, 32'h44f4f9f4},
  {32'hc48864f0, 32'h440c4afe, 32'hc41a6929},
  {32'h43b3be17, 32'hc20fca65, 32'h44baf8f1},
  {32'hc483ac9e, 32'hc42d777f, 32'hc41b2423},
  {32'h4424525a, 32'h4486e0b9, 32'h43ef944b},
  {32'hc1cc9998, 32'h41a935d4, 32'hc425eabc},
  {32'hc46a7802, 32'h44bc1daa, 32'h45058c8b},
  {32'h4232e63c, 32'hc3f62440, 32'hc4bd4619},
  {32'h4320dbfd, 32'h44ee84eb, 32'hc2967ec1},
  {32'hc48b5e3c, 32'hc493e6b6, 32'hc436f986},
  {32'hc2c3df00, 32'h44f3b184, 32'hc3a1c5b7},
  {32'hc4f9fa56, 32'hc3a9a07d, 32'h435df19a},
  {32'h43dee3f8, 32'h452b8b73, 32'h44047b4e},
  {32'hc50d50a0, 32'hc3a22887, 32'hc2c5da8d},
  {32'h45258cca, 32'h42378e8a, 32'h43ead8f8},
  {32'hc3723b20, 32'h449ff5f1, 32'hc2586cfe},
  {32'h44e7d036, 32'hc31b36ec, 32'h442c81dc},
  {32'h44425a5e, 32'h42cab445, 32'hc47bc2cf},
  {32'hc3b898f8, 32'hc496af64, 32'h44e77214},
  {32'hc448cef6, 32'hc31f19fc, 32'hc49d0d64},
  {32'h4231a06e, 32'h45618cf2, 32'hc370b262},
  {32'hc408de98, 32'hc3c44184, 32'hc5334467},
  {32'h44c9c760, 32'h432dbd00, 32'h43d0806c},
  {32'h448fcdd9, 32'hc4a00658, 32'hc4907830},
  {32'hc3c57000, 32'h443880d3, 32'h44df3202},
  {32'hc4a97c6d, 32'hc386820d, 32'hc3a073ae},
  {32'h439291d6, 32'hc4ac6b9f, 32'h446fa932},
  {32'h440f60b8, 32'hc4b3cc78, 32'hc433821b},
  {32'h44092a75, 32'h4498788f, 32'hc3df3d10},
  {32'h44b20769, 32'hc383bf53, 32'hc406ea9e},
  {32'hc3de69f8, 32'h4450c2e2, 32'h44a49a7a},
  {32'hc464b5cd, 32'hc41480fe, 32'hc3ab642e},
  {32'hc4bf7643, 32'h43b7ddec, 32'h43d2c9b7},
  {32'h4465789e, 32'hc4ce7fce, 32'hc45dbd97},
  {32'h44ac65b0, 32'hc1f93b14, 32'h437123f4},
  {32'h433f2410, 32'hc562b0f7, 32'hc34fb554},
  {32'hc53ce4bf, 32'h4393ecfd, 32'hc3873d81},
  {32'hc42382a8, 32'hc432abac, 32'h42e417ee},
  {32'hc52e0505, 32'h441e6590, 32'hc3275b15},
  {32'h42d5e410, 32'hc50a2566, 32'hc3832f7b},
  {32'h43bcea01, 32'h4455566b, 32'hc29c445c},
  {32'h44a53422, 32'h43c6b879, 32'h43de4b51},
  {32'hc3b8d74c, 32'hc30a43d6, 32'h43998560},
  {32'h44aba718, 32'hc262e4f6, 32'hc3dd4e3c},
  {32'h454f1325, 32'hc3507b86, 32'hc3918024},
  {32'hc5184338, 32'h437ec729, 32'hc391e209},
  {32'h4519476e, 32'h419a2673, 32'h433b856b},
  {32'hc48406ae, 32'h430bdbec, 32'hc33f1f48},
  {32'h440e20ed, 32'hc5297e8f, 32'hc3446dcc},
  {32'hc48883bc, 32'h4452cd1a, 32'hc286c36a},
  {32'h44039674, 32'hc4695d44, 32'h438c6876},
  {32'hc4fde46f, 32'h43dab8d6, 32'hc181c25b},
  {32'h43e74185, 32'hc4b0efb0, 32'h4369e27c},
  {32'h44448ea4, 32'hc315df92, 32'hc3ef71c1},
  {32'h44a74e96, 32'hc3c9667d, 32'h447999df},
  {32'hc2ef6bb0, 32'h442e6444, 32'h4435a2f6},
  {32'hc3b422c6, 32'hc21bf71a, 32'hc1323418},
  {32'hc4676e55, 32'h43a1ff8a, 32'h44612801},
  {32'hc36977ca, 32'h423dac9d, 32'hc53f9a8e},
  {32'hc3cfbe57, 32'hc1cc5fe7, 32'h443473d7},
  {32'h427da840, 32'hc4a58229, 32'hc3c97b42},
  {32'h42da8534, 32'h44fb54f7, 32'h431e6486},
  {32'hc30e2c18, 32'hc33b551b, 32'hc3e38e57},
  {32'hc50d517c, 32'h4432da4c, 32'h44a4ec94},
  {32'h455e0055, 32'hc38b93d6, 32'hc340f9ef},
  {32'hc4b6a823, 32'h43530d0f, 32'hc329bab9},
  {32'h44eb2582, 32'hc3b1a956, 32'hc28c85eb},
  {32'hc2c621e4, 32'h4445ac07, 32'h43bc6d4c},
  {32'h4421868a, 32'h43b566c2, 32'h42654bc1},
  {32'hc3bec6ba, 32'h4536e1f7, 32'h4329205e},
  {32'h453af26a, 32'hc3e4d5e2, 32'hc409e35a},
  {32'h44424e25, 32'hc344a4c6, 32'hc52e6822},
  {32'hc53aa724, 32'h420e2807, 32'h441ab0f7},
  {32'h441c0401, 32'h4450b992, 32'hc3317e5a},
  {32'hc3a68958, 32'hc5098d49, 32'h41ab448d},
  {32'h443ed0ab, 32'h44753bb6, 32'h441924e1},
  {32'h440d735e, 32'hc3948f16, 32'h43843382},
  {32'h43cfa1ac, 32'h445020d3, 32'h42a4d925},
  {32'hc4483abf, 32'hc50a840c, 32'hc26b272e},
  {32'h43c7d38f, 32'h44c41d3e, 32'h4337a7d2},
  {32'hc50ce02e, 32'hc3b20adf, 32'hc351828b},
  {32'h440258e4, 32'h4407bbb2, 32'h43f61d96},
  {32'hc4ed5887, 32'h429c4785, 32'h43180e7f},
  {32'h4466d402, 32'h4430fcad, 32'h43e8c347},
  {32'hc390e660, 32'hc440094d, 32'hc4cf3b7c},
  {32'hc4527a6b, 32'h440928b6, 32'h43a62f49},
  {32'h43327abd, 32'hc46a2e11, 32'hc4428316},
  {32'h4479084c, 32'h447db2c6, 32'h439d3084},
  {32'hc26cafa2, 32'hc3fbc584, 32'hc35a819f},
  {32'h4540a8d2, 32'hc3ca6ae1, 32'h43530b73},
  {32'hc5145723, 32'hc3473b04, 32'hc3c526ca},
  {32'hc4220cec, 32'hc2a5b0ec, 32'hc3e5ac74},
  {32'hc4de48b6, 32'hc31dfdbd, 32'hc41138ec},
  {32'h43a1d918, 32'h44aa5d73, 32'h43c533ea},
  {32'hc4aaed66, 32'hc224438c, 32'hc3c3f3b1},
  {32'h44d9c500, 32'h43a75368, 32'h4475d107},
  {32'hc4860d8a, 32'hc381f86a, 32'hc4ffe422},
  {32'h4458e8cb, 32'h43f79480, 32'h443ee527},
  {32'hc46c0b38, 32'h441fc6eb, 32'h436eb2fb},
  {32'hc48a5bf8, 32'hc474b9d0, 32'hc309b711},
  {32'h452e3eaf, 32'h446f89db, 32'h43878df8},
  {32'h43333d8c, 32'hc4905b95, 32'h4351731b},
  {32'h44300e6f, 32'h450885f2, 32'h438c147f},
  {32'hc49187f6, 32'hc436aa39, 32'hc3cf8f27},
  {32'h45390d94, 32'h437e72c2, 32'hc364acd4},
  {32'hc45f2d38, 32'h431ab04e, 32'hc37e48c4},
  {32'h4523234e, 32'hc38ac400, 32'hc2694b23},
  {32'hc427bcb8, 32'hc420e67c, 32'hc3ad3c44},
  {32'hc1f7c9c0, 32'h44a42038, 32'hc3938148},
  {32'hc4dc184e, 32'hc30fdc4f, 32'hc389e98c},
  {32'hc4661028, 32'h441edd3e, 32'hc32475f4},
  {32'hc471825e, 32'hc30fcd30, 32'h44212339},
  {32'h44e9fdec, 32'h431a38a3, 32'hc3beb378},
  {32'hc47ece81, 32'hc40c9d9b, 32'h43be814e},
  {32'h4521bef3, 32'h44017fd3, 32'hc35d7ac6},
  {32'hc48dd5fa, 32'hbf902030, 32'h44c2d4bd},
  {32'hc492d08a, 32'h43b606ca, 32'hc3930d56},
  {32'hc4b1efb5, 32'hc50436e9, 32'h43431c0d},
  {32'h44fa86aa, 32'h449a55f7, 32'hc42cedf0},
  {32'hc3e941f4, 32'hc3d6039e, 32'h446856b8},
  {32'h416a5a00, 32'h447a5bad, 32'hc4916b59},
  {32'hc4aab120, 32'hc4797bc1, 32'h42b659a2},
  {32'hc48e85e3, 32'hc2c7c4e2, 32'hc3ff301f},
  {32'hc58bad2e, 32'h43444392, 32'h42794469},
  {32'h430dd940, 32'h432729ca, 32'hc35c5b99},
  {32'h450df03b, 32'h4194497e, 32'hc3c5884c},
  {32'hc4b72aa8, 32'h444f93ae, 32'h4458d892},
  {32'hc4d404cc, 32'h43666b85, 32'h43a07ce4},
  {32'hc4431858, 32'hc317c5ea, 32'hc404fa1c},
  {32'h44e0e2ee, 32'hc3da869d, 32'h433bb532},
  {32'h40f38680, 32'h44f3c33b, 32'h4323078a},
  {32'h45400ac9, 32'hc3d436a8, 32'hc4269b0a},
  {32'hc5204dfa, 32'h43d2d7a0, 32'h42b9988c},
  {32'h45298199, 32'h43170871, 32'h4383592f},
  {32'hc3fcd6a8, 32'h43a91674, 32'hc4339e33},
  {32'h43a4c7d0, 32'hc4ac2c3c, 32'h43460305},
  {32'h4214995e, 32'h44600343, 32'hc24e8387},
  {32'h44a91f11, 32'hc35ad5a2, 32'h4487532f},
  {32'hc5021d54, 32'h42f3c515, 32'hc344e0cf},
  {32'h42f0e9de, 32'h4291da67, 32'h44984ede},
  {32'h4094f9b0, 32'hc347be99, 32'hc4e405a3},
  {32'h4427f758, 32'h44284614, 32'hc3912512},
  {32'h44c1f230, 32'h43fbfb7e, 32'h438bc1bc},
  {32'h41ada280, 32'hc5098fb6, 32'h439a40c4},
  {32'hc4245cc3, 32'h44418e57, 32'hc49ec708},
  {32'hc4c84cd0, 32'h430267b3, 32'h425db84d},
  {32'hc3dbea2c, 32'h455d7c83, 32'h4142cf71},
  {32'h442a1c01, 32'hc5071324, 32'h43ff762b},
  {32'h43ab7bf0, 32'h44de1e22, 32'h439bc454},
  {32'h440da2f7, 32'h42055789, 32'h443fa3bb},
  {32'hc4c48fdc, 32'hc423a174, 32'hc5139cf4},
  {32'hc491a88b, 32'h42dbf823, 32'hc4000ed4},
  {32'hc37dea83, 32'h43b76e97, 32'hc4c1d377},
  {32'h44cc44d6, 32'hc3de1115, 32'h439f361f},
  {32'hc3499256, 32'h43674ec1, 32'hc40bffe9},
  {32'h43e387a4, 32'hc2c896b5, 32'hc48251f1},
  {32'h44a2876e, 32'hc37f44ac, 32'hc3336d8f},
  {32'hc492271c, 32'h4223bb3a, 32'hc40e1353},
  {32'h44113d24, 32'hc2f19250, 32'h447b56a5},
  {32'hc49dbd11, 32'h430ca402, 32'hc50074e3},
  {32'h438e9300, 32'hc537b023, 32'h431cb097},
  {32'hc37a4b70, 32'hc2c129a3, 32'h43e86647},
  {32'h41d0599b, 32'hc4dfff0f, 32'hc4f055ee},
  {32'hc39ecb27, 32'hc40dea0e, 32'h44a6ad16},
  {32'h43be9572, 32'hc4dc2fd9, 32'h43be4693},
  {32'hc444e0ce, 32'h433b1d7b, 32'hc28168b5},
  {32'h443fceb5, 32'hc2be5d65, 32'h439c1d52},
  {32'h43a0843c, 32'hc3309356, 32'hc2d17685},
  {32'h45099f1f, 32'hc3000806, 32'h4426be00},
  {32'hc419105d, 32'h44df9ee9, 32'hc4221a9e},
  {32'h451e793c, 32'hc3d8fc2b, 32'h42f999f9},
  {32'hc59b680c, 32'h432812c4, 32'hc1ad2b66},
  {32'h425243e0, 32'hc3ac5b91, 32'hc1ffa465},
  {32'h44cef176, 32'h428bcae4, 32'hc40eea61},
  {32'hc358cc28, 32'hc56f21b4, 32'hc322ea14},
  {32'hc3fa552a, 32'h4428c2b2, 32'h4358be58},
  {32'hc3f4b1d0, 32'hc422f5ee, 32'hc30354e8},
  {32'hc4168ce5, 32'h453d2dd3, 32'h4301bf39},
  {32'h44c99f3a, 32'hc48849b7, 32'h4343ae84},
  {32'h445b8b26, 32'h44237779, 32'h44b2dace},
  {32'hc3ae4150, 32'hc1f9562b, 32'hc5693062},
  {32'hc383a55e, 32'h44415467, 32'h45109893},
  {32'hc52f8d3e, 32'hc3242ff8, 32'h4426092e},
  {32'h44606091, 32'h43b07861, 32'hc477de9e},
  {32'h439a07df, 32'hc437ef39, 32'h446d62bf},
  {32'h44a18181, 32'h445aad52, 32'hc3f430b1},
  {32'hc538d0dc, 32'hc2434a84, 32'hc35c33f0},
  {32'h44b98e41, 32'hc3a2dd76, 32'hc2df8831},
  {32'h449c49a1, 32'hc338a80f, 32'h43b9e38a},
  {32'hc3375384, 32'h44b4e58e, 32'h45051757},
  {32'h449725c8, 32'hc4922fa3, 32'hc4a0a219},
  {32'h44aa328d, 32'h43f23ddf, 32'hc3ab9beb},
  {32'hc449e1d0, 32'hc4138603, 32'h43b6b37e},
  {32'h450d9bf6, 32'h430aa3f0, 32'h432a4f2d},
  {32'hc406935a, 32'h4378b8ad, 32'h453ba30b},
  {32'h43bac786, 32'h432b1010, 32'hc4de3205},
  {32'h43c4b4ce, 32'hc378f8c0, 32'h431f6b52},
  {32'h44f68fa2, 32'hc31031fe, 32'hc2a41a64},
  {32'hc4b15583, 32'hc1c6590b, 32'h444094b6},
  {32'hc486600f, 32'h439d6ef7, 32'hc39576bc},
  {32'h42d60d92, 32'hc4d1e98a, 32'hc3c2f75e},
  {32'h448d5796, 32'h443095d9, 32'hc354d209},
  {32'h450bc5fe, 32'hc213f47a, 32'hc381912c},
  {32'h450a29fd, 32'h446033b9, 32'hc3ef803e},
  {32'h437bec00, 32'hc53537b6, 32'hc38f0ec0},
  {32'h448c62ee, 32'h444eb279, 32'hc301fd5e},
  {32'hc41b8ba8, 32'hc414b172, 32'h4330bb91},
  {32'h43daab3f, 32'h449b1035, 32'hc3e43dcb},
  {32'h4210e000, 32'hc4e8c6fb, 32'h44f40194},
  {32'h43d65b70, 32'hc46de03a, 32'hc389a3a8},
  {32'h44972808, 32'h431499eb, 32'h44f8b7e4},
  {32'hc47d376b, 32'hc498298c, 32'hc346f84d},
  {32'h4435afcf, 32'h44118d62, 32'h4383faba},
  {32'hc479f19e, 32'h43883625, 32'hc457a99b},
  {32'hc305592e, 32'h44a7ee37, 32'h44ec9d3a},
  {32'h44e0e704, 32'h43902b1c, 32'hc3d4aabc},
  {32'h44150fda, 32'h43d77368, 32'hc387386a},
  {32'hc2078940, 32'h422f7b6c, 32'hc44ba1b1},
  {32'h44a8f914, 32'hc272d773, 32'h4434a8fc},
  {32'hc44b989e, 32'hc4b99e85, 32'h4233d9b9},
  {32'h43fd5bf5, 32'h44bf7e97, 32'h44824827},
  {32'hc43d78d6, 32'hc33bd62a, 32'hc303c921},
  {32'h453c7ac5, 32'h44194e1c, 32'h43c5a819},
  {32'hc33dec37, 32'hc465a9d1, 32'hc48b1790},
  {32'h453bba86, 32'hc3b439de, 32'hc10a6918},
  {32'hc47a876c, 32'hc42332cd, 32'hc2b5e627},
  {32'hc32f8c30, 32'h44ec162e, 32'h42c608e2},
  {32'hc4f3620e, 32'h4458ef58, 32'h4237d305},
  {32'h42a94de0, 32'h44e7541d, 32'h430bf9ef},
  {32'hc48adcd4, 32'hc455c7b7, 32'h43af2c08},
  {32'hc4f76dc5, 32'h42176241, 32'hc409b9d2},
  {32'hc58e609d, 32'h4368b167, 32'hc27612cd},
  {32'h45758058, 32'h431cb2a9, 32'hc3eda869},
  {32'hc3620308, 32'hc4d52e92, 32'hc43de944},
  {32'h432de967, 32'h4514f8bc, 32'hc2d4d6c4},
  {32'hc3b7d368, 32'hc3b7d2b4, 32'hc3e8414c},
  {32'h434bb34a, 32'h44d2fb42, 32'h4474946e},
  {32'hc2b88ac0, 32'hc56ea890, 32'h40284fd4},
  {32'h436c033c, 32'hc300d036, 32'h42ff47fd},
  {32'h44102e88, 32'h42f8d0af, 32'hc40d88d9},
  {32'h4345760c, 32'h43741f5e, 32'h449aadd1},
  {32'h434d43d5, 32'hc4006a8d, 32'hc4ae8312},
  {32'h43cc997e, 32'hc44debee, 32'h451b04d1},
  {32'h43523d44, 32'h44887aec, 32'hc4c15d31},
  {32'hc4487c8f, 32'h440155ef, 32'h423bc4f2},
  {32'h43e6d6dc, 32'hc4b36d38, 32'hc42be5db},
  {32'hc38c85cf, 32'h453e1583, 32'hc3585016},
  {32'h43fec526, 32'hc42011a9, 32'hc4217eff},
  {32'hc2a9bf30, 32'h44ca8406, 32'h44bcb64b},
  {32'h443329ae, 32'h44223df3, 32'hc41fadf8},
  {32'h4417cba4, 32'h429ff9ab, 32'h4472a207},
  {32'h4414f8fb, 32'hc45fb0b2, 32'hc4482e14},
  {32'hc520edb0, 32'h448555f2, 32'h43be2ba6},
  {32'h44ae550d, 32'h43017356, 32'hc1cd19e6},
  {32'hc4040edc, 32'h446a4c46, 32'hc2afc886},
  {32'h43b2a772, 32'hc409b79b, 32'hc3895b43},
  {32'hc4ab2b54, 32'h443e96fe, 32'h422735c4},
  {32'h44fb9c42, 32'h44002eb1, 32'h41e87af7},
  {32'hc4e96daf, 32'hc3f89c70, 32'h430d14e3},
  {32'h450a6cf9, 32'hc431aa08, 32'hc34d6502},
  {32'h447713ed, 32'h438f2e84, 32'h448ad0cf},
  {32'hc4d552f5, 32'hc3165961, 32'hc427d3e4},
  {32'h43a44a7f, 32'hc30de56e, 32'h455af237},
  {32'h4504f918, 32'hc37792ae, 32'hc116d37b},
  {32'h44ef39a0, 32'hc385ae0f, 32'h438cb71b},
  {32'hc3c02a20, 32'h451b2938, 32'h433e9b37},
  {32'h4426d6fa, 32'h4322e277, 32'h439200c9},
  {32'hc4d0229b, 32'h4445f194, 32'hc201f38a},
  {32'hc3a34c43, 32'hc56cf70c, 32'hc2ebc73c},
  {32'hc49a8a97, 32'hc2293e84, 32'hc4292128},
  {32'h44a6c5cc, 32'hc35ccd5d, 32'h43b05391},
  {32'hc49eaa41, 32'h435c9722, 32'hc3c8d077},
  {32'h42a9e340, 32'h42099e53, 32'hc4e83045},
  {32'hc36df79c, 32'h445c14cb, 32'hc31664d4},
  {32'h4385b3e4, 32'hc41eaa1b, 32'hc32707d8},
  {32'h446cf1fe, 32'h42f5cf26, 32'h43af6b78},
  {32'h43d1abd4, 32'hc413bee3, 32'hc4bc592e},
  {32'hc4e9b092, 32'hc37599be, 32'h443ca271},
  {32'h45220bc1, 32'hc3f3b77f, 32'h4234e0d6},
  {32'hc50d9b18, 32'h44125e72, 32'h448ad3b5},
  {32'hc35b8d59, 32'h43d8b832, 32'hc3dfb61f},
  {32'h449ce094, 32'hc2c73cca, 32'h43a8bb61},
  {32'h4422bcbc, 32'hc4edef71, 32'h41b027f6},
  {32'hc4cdcc3f, 32'hc31a5269, 32'h447e6ac3},
  {32'h432f22b5, 32'hc395332b, 32'hc3851ce1},
  {32'hc52b8b2a, 32'h441e8aae, 32'h4337c801},
  {32'h42df74ea, 32'hc527e1f6, 32'hc3a2f6b0},
  {32'h448b59ec, 32'hc3af07e0, 32'hc544648c},
  {32'hc3b7afd8, 32'hc399fd19, 32'h4467ed16},
  {32'h4305a5c0, 32'h44650a42, 32'hc47bafd6},
  {32'hc427da6e, 32'hc44f433e, 32'hc189247a},
  {32'h45398662, 32'hc2f47de0, 32'hc3141ec7},
  {32'hc415f8c4, 32'hc4381074, 32'h43a9285d},
  {32'h44dae36d, 32'h448777cc, 32'h428e6e3e},
  {32'hc4bb5ef3, 32'hc4f21d56, 32'h43a3ce48},
  {32'h454261b2, 32'h3e78e980, 32'h440174b6},
  {32'hc3ce7e48, 32'h441593e0, 32'hc4a14076},
  {32'h450a4182, 32'hc31eb54c, 32'hc30ef1fc},
  {32'hc5124827, 32'hc3cbed36, 32'hc30623aa},
  {32'h44795a1a, 32'hc378dca0, 32'h447d9daa},
  {32'hc43b500c, 32'hc49c7387, 32'hc4cc8124},
  {32'hc3f347c3, 32'h441f97ed, 32'h43c602fa},
  {32'hc3c1b60e, 32'hc38e2f0d, 32'hc4de7fb1},
  {32'h451f4ca4, 32'h43fd6a5e, 32'h429f37bf},
  {32'hc13f2c10, 32'h433f252b, 32'hc3cb113d},
  {32'h43e06270, 32'h445fd466, 32'h44b7f199},
  {32'hc4ebe526, 32'hc31383da, 32'hc499a432},
  {32'h453723e5, 32'h43285395, 32'hc45dad4c},
  {32'hc32aab6f, 32'hc53efaf4, 32'hc4080e2b},
  {32'h44566164, 32'hc1843a98, 32'h44c16a5a},
  {32'hc5127e9d, 32'h42a942c0, 32'h43157e0d},
  {32'h4499ccf2, 32'h44ae5a5d, 32'h4422c8d5},
  {32'hc2cef390, 32'hc48971e7, 32'hc3c671b8},
  {32'h440397ab, 32'h4395f224, 32'h4458f3b6},
  {32'h44e2f95c, 32'hc2d54283, 32'hc3cf8ed3},
  {32'hc5421a97, 32'h431729b6, 32'hc28337a4},
  {32'h4340b9f8, 32'h453896d8, 32'h44507cc4},
  {32'h447c3442, 32'hc3df8c20, 32'h43391758},
  {32'h4444821b, 32'h433ac537, 32'h428f1872},
  {32'hc4905f28, 32'hc3e35a13, 32'hc2ee157b},
  {32'hc3bd4d00, 32'h433c6561, 32'hc11cd088},
  {32'hc4865c82, 32'hc184a0a0, 32'hc48b90a4},
  {32'h45547ec1, 32'h433bdcf7, 32'h4238f26f},
  {32'h43dfaea4, 32'hc331b032, 32'hc42337ef},
  {32'h4503fea3, 32'hc0702670, 32'h443c61d9},
  {32'hc48b2043, 32'hc49edfef, 32'hc2b85169},
  {32'h4513d2c1, 32'h41330048, 32'hc324443f},
  {32'hc431480e, 32'hc51e134f, 32'h433aa7a0},
  {32'h44ac272a, 32'h44bd23f1, 32'hc29992f9},
  {32'hc4f3b4b2, 32'h431a764a, 32'hc3849739},
  {32'h43ab7f39, 32'h432b5a38, 32'hc3d00356},
  {32'hc30b2438, 32'h44245403, 32'h4487baed},
  {32'hc416f843, 32'h4479c0e0, 32'hc29215f6},
  {32'hc42280d3, 32'hc4ae190c, 32'h44df7e78},
  {32'h44d14076, 32'h43dc18fa, 32'hc445887d},
  {32'h43a96e66, 32'hc34f9d66, 32'h44982961},
  {32'h455b3fbd, 32'h442fdbb1, 32'hc360cf2b},
  {32'hc2f472d0, 32'hc550a0d9, 32'hc2d66a37},
  {32'h45149398, 32'h42f6caba, 32'hc30e8f6b},
  {32'hc5780304, 32'hc342dd2f, 32'h43120108},
  {32'hc3d2c688, 32'hc4149026, 32'hc5531846},
  {32'h443b79a6, 32'hc492dbd7, 32'hc36824f6},
  {32'hc5602df5, 32'h43a04fd9, 32'h4124edf8},
  {32'h44779ece, 32'hc4a0366e, 32'h43ba3417},
  {32'hc3dab1b6, 32'h4525b280, 32'h4316a123},
  {32'h44c8f081, 32'hc40de4a3, 32'hc394fbeb},
  {32'hc282a1c0, 32'hc292a9e0, 32'h4262aec4},
  {32'h44d04170, 32'hc4659e22, 32'hc3dbfcfc},
  {32'hc4fd955a, 32'h4347f1e8, 32'h4051516c},
  {32'h451d92ca, 32'hc2c5b84d, 32'h4415f17d},
  {32'hc30f1518, 32'h45074caf, 32'hc3b85674},
  {32'hc2c9ad3c, 32'hc4821882, 32'hc4504484},
  {32'hc3a06fc4, 32'h40133640, 32'hc483e7d0},
  {32'h430e7bcc, 32'h43ed5bf9, 32'h445a62a9},
  {32'hc44a8abc, 32'h44bb9bc8, 32'h4201ceb8},
  {32'h4394a346, 32'h438cb6a7, 32'h4442fd4d},
  {32'hc3e18272, 32'hc39f9e83, 32'hc50eb946},
  {32'h452d76cc, 32'hc4498867, 32'h4315c11e},
  {32'h442fa07e, 32'hc3485d87, 32'hc447331a},
  {32'h428f7840, 32'hc4bdedbe, 32'h44ff2b9c},
  {32'hc24f75c0, 32'h44c6798c, 32'hc47788f1},
  {32'hc4119909, 32'hc3bffa10, 32'h4329f868},
  {32'hc466f5bc, 32'h4355a82b, 32'hc5084dbe},
  {32'h44cb32c5, 32'hc27d4cb7, 32'h44679424},
  {32'hc4d9673a, 32'h4419155d, 32'hc3bb5343},
  {32'h44ab9473, 32'hc1729524, 32'h44c32e8c},
  {32'hc590562a, 32'h43904c19, 32'h436b31d9},
  {32'hc3a1e7c5, 32'h42b0f9a2, 32'h440460c8},
  {32'hc467d7d7, 32'h438f3c8b, 32'hc4483bcd},
  {32'hc33b3e9c, 32'h44b0b9a2, 32'h452b37ab},
  {32'h4490a6f8, 32'h43010c0a, 32'hc406704c},
  {32'h439c08db, 32'h43917199, 32'h41e43f88},
  {32'h45466a1c, 32'hc3ab89b6, 32'hc37c7c9c},
  {32'hc4827c71, 32'h43c1cb92, 32'hc41cd3e1},
  {32'h449f64ad, 32'h437d571b, 32'h43cce343},
  {32'h431e430b, 32'hc3635b80, 32'hc4e7c585},
  {32'h44dc1405, 32'hc3dbff37, 32'h44101f84},
  {32'h449476c6, 32'hc453a284, 32'h44553020},
  {32'hc416ce8f, 32'hc2905c16, 32'hc48bac7e},
  {32'h4427e927, 32'hc4cc6cf9, 32'h441d7825},
  {32'h44de3cbc, 32'hc3867f59, 32'hc3528a50},
  {32'hc4968ae2, 32'h42acdf9a, 32'hc4792ce3},
  {32'h442bcde7, 32'hc36f3e09, 32'h44596052},
  {32'hc520e25c, 32'hc3166355, 32'h4386070a},
  {32'h44ef4f32, 32'hc3a38927, 32'h4338d10c},
  {32'hc4d7e5d6, 32'h44030860, 32'hc269544e},
  {32'h4553e783, 32'hc146d1b1, 32'hc1c0c03b},
  {32'hc53acd47, 32'hc41417ba, 32'h43ae61c6},
  {32'h44b9a4d3, 32'hc30052ee, 32'h44303d6a},
  {32'h44167eba, 32'h44809492, 32'hc32fd7a3},
  {32'h43cd11d2, 32'hc500ca15, 32'h44213841},
  {32'h440042de, 32'h4566cdc5, 32'hc24571a2},
  {32'h44ad7db8, 32'hc3afa724, 32'h43ba405c},
  {32'hc5334d10, 32'h43d50382, 32'h441458f2},
  {32'h44849086, 32'hc4e0dde1, 32'h439c64b7},
  {32'h441541d8, 32'h448d2e22, 32'h44b9ed66},
  {32'h43acea0a, 32'hc4189900, 32'hc43a3f0d},
  {32'h42ac3984, 32'h44b8eb1d, 32'h451a1018},
  {32'hc52501d2, 32'h4317bd9e, 32'h4262182c},
  {32'h43f9cf2c, 32'h448da70a, 32'hc17c39d4},
  {32'hc480f24e, 32'hc3ed030c, 32'hc0801c64},
  {32'h4506c4c8, 32'h439d16d7, 32'h41c36105},
  {32'hc2cc228d, 32'hc18ace49, 32'h44d7caa5},
  {32'h44fefb37, 32'h439ed1f5, 32'hc28591e3},
  {32'h43c7409c, 32'h43833fee, 32'hc493f7a9},
  {32'hc4f9dfda, 32'hc3f5a6a8, 32'h43d38cf9},
  {32'hc26c58d0, 32'h44f42e9c, 32'hc5013e28},
  {32'h444b5d4a, 32'h440c3148, 32'hc4cdf91f},
  {32'hc3b09dea, 32'hc38c86af, 32'h44b4ffd6},
  {32'h43b0cb58, 32'h450adbe0, 32'h41793b29},
  {32'hc39a0dfb, 32'h43a08b10, 32'h44636eed},
  {32'h42883eec, 32'h43c7a9b6, 32'hc4315add},
  {32'hc436af84, 32'hc39e1bcc, 32'h430e8779},
  {32'h45239ac4, 32'hc28918a3, 32'hc3ce81a4},
  {32'hc54ec7b1, 32'h42622a4c, 32'h43862db7},
  {32'h4552fb51, 32'h439b3693, 32'hc3170c85},
  {32'hc501585f, 32'hc483f368, 32'hc2a1f31c},
  {32'h44bc83aa, 32'h440ba82b, 32'hc3e47126},
  {32'h4445ef99, 32'hc47f2ebb, 32'h427830b2},
  {32'h44e7144e, 32'h44230775, 32'hc20d28ad},
  {32'hc43f67ff, 32'hc4d0224e, 32'hc34399e3},
  {32'hc456f7c9, 32'h436e95dd, 32'h43c2c44a},
  {32'hc3477109, 32'h4368663b, 32'h43bf6f3b},
  {32'hc5108dba, 32'h4372877d, 32'hc3befbd0},
  {32'hc303cabc, 32'h4539548d, 32'h4428f32f},
  {32'h4488805e, 32'hc40ffbde, 32'hc41ae711},
  {32'h44df684a, 32'h447d0a70, 32'h4113ee3c},
  {32'hc2eba6f1, 32'hc55fe023, 32'hc3894926},
  {32'h44af4a66, 32'hc3f4b3fb, 32'h43896898},
  {32'h407e6c32, 32'hc423e292, 32'hc5342cfe},
  {32'hc31a2ec6, 32'hc1ef8e8b, 32'h44e34c6b},
  {32'hc082d4d0, 32'hc471a0e9, 32'hc1b77d70},
  {32'h43f1961c, 32'hc410def6, 32'h42f1d2d4},
  {32'hc3da8fb5, 32'hc21a7866, 32'hc4e4eb1c},
  {32'hc40f4b9e, 32'h438b8818, 32'h448d89cb},
  {32'h4149e546, 32'h4230fd2e, 32'hc4c0e274},
  {32'h445a739e, 32'h44da7c27, 32'h44058f33},
  {32'hc4e03630, 32'hc3e25f0d, 32'h436a6e89},
  {32'h4310a664, 32'h44d2b470, 32'h449ce42f},
  {32'hc536524b, 32'h423ce434, 32'hc41a1d36},
  {32'hc3c468a6, 32'h439a7d44, 32'h4318db86},
  {32'h435e105c, 32'hc52c57cd, 32'hc380dab1},
  {32'h4456f92d, 32'h44967ffb, 32'h440f0349},
  {32'h44848e46, 32'hc4b49cfd, 32'h43849c4b},
  {32'hc407e03d, 32'h45865129, 32'hc3dd0f55},
  {32'hc4abf320, 32'hc4c0ee1b, 32'h42e00b9e},
  {32'hc4380946, 32'h43a1be33, 32'h41942acb},
  {32'hc480f000, 32'hc3a400ff, 32'hc3ad7fb7},
  {32'h44f68ba4, 32'h42992092, 32'hc29c1027},
  {32'hc1c9f09f, 32'h43918581, 32'hc50a73a2},
  {32'h431a763a, 32'hc4812490, 32'h44ea930d},
  {32'hc0d8beeb, 32'h432ccfa4, 32'h43735bd2},
  {32'hc3644e4c, 32'h43c668c6, 32'h45537b29},
  {32'hc35283c8, 32'hc44a509d, 32'hc47a8646},
  {32'hc427d6e0, 32'h443de5a3, 32'h43a81995},
  {32'h439dd778, 32'hc394c8ec, 32'hc54019f8},
  {32'hc45a0288, 32'h44d96e17, 32'h44954b7d},
  {32'h44366022, 32'hc43d34a9, 32'hc43f755d},
  {32'hc3fa2710, 32'hc4c670d1, 32'h44cec0a2},
  {32'h448bbc7d, 32'h4435dc1a, 32'hc44c4bc8},
  {32'h441ea60d, 32'hc4135d04, 32'h433dd246},
  {32'hc397df89, 32'hc4b865a3, 32'hc4226005},
  {32'hc4a282b1, 32'h43c97500, 32'h4430eb14},
  {32'hc2374abf, 32'hc4a9bdd6, 32'h42fe2c90},
  {32'hc531f240, 32'h41817abe, 32'h4245d7f9},
  {32'hc36cbc02, 32'hc3d5a286, 32'hc55b92cb},
  {32'hc527ec35, 32'hc28cd54f, 32'hc38c4cb8},
  {32'h44eceeea, 32'hc4aa4598, 32'h438244c7},
  {32'hc544bf22, 32'h43e5c473, 32'hc4037298},
  {32'hc3c5417c, 32'hc4c4a555, 32'h41766de0},
  {32'hc4978997, 32'h442af013, 32'hc3e727b3},
  {32'h442812ba, 32'hc553f3b4, 32'h4311b23c},
  {32'hc5187b4a, 32'hc30098ad, 32'h43449baf},
  {32'hc3df454a, 32'hc31408b7, 32'h42902b6f},
  {32'hc5924147, 32'hc2830587, 32'hc3b27db6},
  {32'h4513e7d3, 32'hc242b5ff, 32'hc3b0ef56},
  {32'h451196a4, 32'hc2a672ea, 32'hc3e885c6},
  {32'hc4d4763c, 32'hc2418fae, 32'hc4080ee1},
  {32'h4401af38, 32'h44158977, 32'h44ad8ebc},
  {32'hc48d41d9, 32'h43d393e5, 32'hc24e03f5},
  {32'h423b76fa, 32'hc5503fdb, 32'hc2c262a3},
  {32'h43a33c48, 32'h43b11cb3, 32'h442089a7},
  {32'hc4141dae, 32'hc33d7028, 32'hc427519d},
  {32'hc55677c7, 32'h43cdd96a, 32'h41145d86},
  {32'h446b479c, 32'hc48bfa4a, 32'hc279b203},
  {32'h43e4e9f9, 32'hc1a467cc, 32'hc4624783},
  {32'h446db2a9, 32'h42ef1e3f, 32'h445e2369},
  {32'hc3a85b64, 32'h41e5da91, 32'h42f1c0d8},
  {32'hc4461616, 32'h435a3019, 32'hc45457f3},
  {32'hc434ba98, 32'h42172ccc, 32'h44162868},
  {32'h43113b7c, 32'hc4c120dd, 32'hc3f1f92e},
  {32'hc4d4f822, 32'hc10c58ff, 32'hc231a4ac},
  {32'hc408c042, 32'hc4ffd638, 32'hc42cf835},
  {32'hc4ce4786, 32'hc19c8f5e, 32'hc1ed02d1},
  {32'h40d3a680, 32'hc3640457, 32'h4218f87f},
  {32'hc4420b44, 32'hc44a7ad7, 32'h44b0bea9},
  {32'h45717f4c, 32'h442bcff8, 32'hc2d9a9a1},
  {32'hc3da4cfc, 32'hc387dfb9, 32'h429232da},
  {32'h44f4ee60, 32'hc3f722ad, 32'hc364d434},
  {32'hc3f2bef0, 32'h4413bd8c, 32'h44c10530},
  {32'hc462d5c6, 32'hc42dad37, 32'hc40638be},
  {32'hc3dc3690, 32'h450d7929, 32'hc2f5c3bf},
  {32'h429e6c48, 32'hc540e7c5, 32'h42e8f37f},
  {32'h45199296, 32'hc0861fa0, 32'hc4526e8e},
  {32'hc486c8ed, 32'hc3edd1ef, 32'h44b25613},
  {32'hc363e3aa, 32'h442635f0, 32'h432147af},
  {32'hc41ea2bd, 32'hc4c584d1, 32'hc4059bc7},
  {32'h455daf6f, 32'hc31e3dcc, 32'hc372740b},
  {32'hc5306c5e, 32'hc2d56b6b, 32'hc1b96db7},
  {32'h44bf9274, 32'h44c160b8, 32'h435ffed4},
  {32'hc53a60c5, 32'hc39fe426, 32'h43abe05a},
  {32'hc454155d, 32'h441a78c2, 32'h43b8f902},
  {32'hc52fbbf0, 32'hc40b58c5, 32'hc28cc274},
  {32'hc2711b50, 32'h43aaaaf5, 32'h441a3504},
  {32'h44d5de5f, 32'hc2ffa490, 32'h43028ebe},
  {32'h41972cf4, 32'h4420d3d5, 32'h44c2d55b},
  {32'hc536d8e6, 32'hc35dac7e, 32'hc37df857},
  {32'h43ad315c, 32'hc2497b62, 32'h4409c6f0},
  {32'hc4d9dc28, 32'hc21734c6, 32'hc48e7eef},
  {32'h4431a96e, 32'h445138fa, 32'h449abb4f},
  {32'h4441168c, 32'hc43604f6, 32'hc37b850f},
  {32'h45002c7c, 32'h4347d425, 32'h4400f811},
  {32'hc53555d1, 32'hc2c84916, 32'hc3baba8b},
  {32'h44d351d8, 32'h440b6ed2, 32'h41a3809e},
  {32'hc4d6a692, 32'hc49d0056, 32'hc382bb44},
  {32'h44807f26, 32'h439348ac, 32'h43d9cc73},
  {32'h44c42015, 32'h42a62f62, 32'h4368f62b},
  {32'h41b7aec0, 32'h4454392c, 32'h440c818a},
  {32'h43ac0f2c, 32'hc4e99951, 32'hc49ddeea},
  {32'h44d19861, 32'h43a22456, 32'hc32bd41d},
  {32'hc4a5c0db, 32'h435600ef, 32'h414497ba},
  {32'hc383fc88, 32'hc4c3a9cb, 32'hc15ccaa2},
  {32'h44dfe43d, 32'h44323532, 32'h440049ae},
  {32'h44bcf350, 32'h439dea7e, 32'h4211c6ad},
  {32'h4440b896, 32'h44cd062d, 32'h4335ec31},
  {32'hc48802a6, 32'hc4ae8261, 32'hc2d9f1a3},
  {32'h450a0ae4, 32'hc20776c4, 32'h422350a5},
  {32'hc54b5519, 32'hc3cd5739, 32'h43374f83},
  {32'h4504c8b9, 32'h43f7d332, 32'h4239e17b},
  {32'h42dbd5f0, 32'h4103ce9c, 32'h446796c3},
  {32'h44ac5638, 32'h43d6f770, 32'hc39cca79},
  {32'hc41dc8f7, 32'hc430f449, 32'hc3a79157},
  {32'h426a3d0f, 32'hc1b70b6e, 32'hc4c38f9b},
  {32'hc39a1954, 32'hc34fc1fb, 32'h43dbb85e},
  {32'h4411778c, 32'h4493500a, 32'hc3e292ae},
  {32'hc4b6f506, 32'hc2dfb6b8, 32'h43ac4301},
  {32'h451cef9a, 32'h43988814, 32'h42e7db80},
  {32'hc38dc31b, 32'h4259438b, 32'h451e5ebd},
  {32'h44c9f149, 32'h42a4a171, 32'hc3f09275},
  {32'hc35ff1e4, 32'hc519e47f, 32'h433c32cf},
  {32'h43ffcfb0, 32'h451ff2ad, 32'hc395445b},
  {32'h434ecef7, 32'hc3bdd4b2, 32'h44d2a577},
  {32'h42171207, 32'h441c4fed, 32'hc4938aeb},
  {32'hc43b5464, 32'hc4748df8, 32'h43bc3baa},
  {32'h44490e76, 32'h4372ed70, 32'hc40f99e1},
  {32'hc4c6c5a6, 32'h410300dc, 32'h4467666d},
  {32'h44d32046, 32'hbef48260, 32'hc4bcb10a},
  {32'h432ee8c8, 32'hc4d080aa, 32'hc418c13e},
  {32'hc51bf3f8, 32'h44160ab1, 32'h437821e0},
  {32'hc40d359b, 32'hc4a88dcb, 32'h42bfd4a2},
  {32'hc42ebf28, 32'h450e44ee, 32'hc4036e93},
  {32'h449b9818, 32'hc4869589, 32'hc2e7ee06},
  {32'h43e8c7fd, 32'h44256fb5, 32'hc2bd6286},
  {32'hc3f1b984, 32'hc3785d93, 32'hc49e0cea},
  {32'hc5110795, 32'h447edbca, 32'h441c22a0},
  {32'hc40c122a, 32'h41d5e33a, 32'h432702f3},
  {32'hc3ce3dde, 32'h442d3bf6, 32'hc4b7962a},
  {32'h4515c84a, 32'hc17faac0, 32'h43557cd8},
  {32'hc513782a, 32'hc392de69, 32'hc3551bfe},
  {32'h44eebcba, 32'hc486b1f2, 32'h43286d07},
  {32'hc42f052f, 32'h448cd8d9, 32'hc33f0847},
  {32'h438970f2, 32'hc2afe14d, 32'h43a7483d},
  {32'hc490906a, 32'h43c4a6e6, 32'hc3df085b},
  {32'h4428601a, 32'hc478259b, 32'h430b2700},
  {32'hc4aedbe7, 32'hc2d5c641, 32'hc30b2910},
  {32'h44488658, 32'hc4661072, 32'h44c7324e},
  {32'hc42c852c, 32'h4401a797, 32'hc51c2b31},
  {32'hc423ae0b, 32'hc45b6b56, 32'h4487c2dd},
  {32'hc4cbeca9, 32'h4491340b, 32'hc404ed5c},
  {32'h442f7d22, 32'hc4804bc9, 32'h43bcf35d},
  {32'h417442b2, 32'h43f42c7c, 32'h4210a624},
  {32'h43514783, 32'hc38c3bb7, 32'h446190cd},
  {32'hc5704180, 32'h422f2fc4, 32'hc309e9d2},
  {32'h4346e2d8, 32'hc2ea9dbc, 32'hc3cacb7e},
  {32'h441541b4, 32'h44a0e936, 32'hc4fada79},
  {32'h446ea960, 32'hc42a89c6, 32'h44246338},
  {32'hc212c680, 32'hc4c77bd2, 32'hc4156e08},
  {32'h448b760e, 32'h4329d417, 32'hc47ece3b},
  {32'h44657a0e, 32'hc3007c86, 32'h44828ccf},
  {32'hc3d1de0c, 32'hc405c78a, 32'hc5240803},
  {32'hc4a02569, 32'hc36768cc, 32'hc2d6e3f3},
  {32'hc49706da, 32'h44ca8b37, 32'hc39c5c6b},
  {32'h4482f198, 32'hc484040b, 32'h43d9ca7f},
  {32'h43fdde7e, 32'hc46e03aa, 32'h4473c50b},
  {32'hc3df656d, 32'h43ca7788, 32'hc4adb37d},
  {32'h44cd8766, 32'h43315e42, 32'hc297b4a5},
  {32'h431c2289, 32'hc243ade2, 32'h44b113bd},
  {32'hc41d774f, 32'h440ac07d, 32'hc281924b},
  {32'h43792b90, 32'hc304a020, 32'h410590be},
  {32'h438409c6, 32'h4428e38e, 32'hc4249c5f},
  {32'h4486ca12, 32'hc40cbaa2, 32'h4389f5ba},
  {32'hc3a32de3, 32'h43ccd470, 32'hc24f0b1b},
  {32'h45888e00, 32'hc3df471c, 32'h429c28bc},
  {32'hc524b336, 32'hc308a188, 32'hc3bf8e92},
  {32'h4568fc6e, 32'hc3b56cac, 32'h43c29e38},
  {32'h41be1e30, 32'h43d996db, 32'hc4402308},
  {32'h448a00aa, 32'hc4d2a1c5, 32'hc40848b2},
  {32'hc4f3dcad, 32'h43d4ab68, 32'hc20bd86a},
  {32'hc396d022, 32'hc4884a06, 32'h436f0b76},
  {32'hc4080bfe, 32'h44c8636a, 32'h4325b524},
  {32'hc382b4c2, 32'hc549a1c8, 32'hc3c0ce53},
  {32'hc4d4aa23, 32'hc26b29c6, 32'hc30b988b},
  {32'h4231f3d0, 32'h4412374b, 32'hc49481b6},
  {32'hc4794bbb, 32'h43d68ce9, 32'h4427691b},
  {32'hc4655c2a, 32'hc4510a57, 32'h448f1cd1},
  {32'h4535da14, 32'hc3858cde, 32'hc3bac699},
  {32'h44bed5b3, 32'h426472ea, 32'h4394fe67},
  {32'h441352a6, 32'h41e1d5ef, 32'hc5200f7d},
  {32'hc4509fb0, 32'hc4dcf471, 32'h43ae8cc9},
  {32'hc4fdb496, 32'h42806f7b, 32'hc28e84a4},
  {32'h443f311b, 32'h4457a0c0, 32'hc4a32f83},
  {32'hc48a60d9, 32'hc388eb65, 32'h44dff719},
  {32'hc3130b19, 32'h44ef5cac, 32'hc4cf5116},
  {32'h45122fdf, 32'h43b78be2, 32'hc39f28d6},
  {32'hc4bda304, 32'hc40aba16, 32'h438bc55d},
  {32'h434afc7e, 32'h450155b4, 32'h42707545},
  {32'hc3ccfe90, 32'hc3e3c559, 32'hc3219c2b},
  {32'h446f987a, 32'h4440cd9d, 32'hc4737172},
  {32'h44837a2b, 32'hc35baaca, 32'h43fff555},
  {32'h4544a1f8, 32'hc32fcc38, 32'h427287b8},
  {32'hc4ac5331, 32'h437b3a8c, 32'h4390021f},
  {32'h44c8e43b, 32'h42323914, 32'hc41255c3},
  {32'hc232c738, 32'hc57f1bea, 32'hc1ece864},
  {32'h44df26ce, 32'h443359c1, 32'hc291ce37},
  {32'hc45ed02b, 32'hc402eee0, 32'h438910ec},
  {32'h43cb53bb, 32'h44f18855, 32'hc3872a39},
  {32'hc4ff7ab3, 32'hc4424f66, 32'h440d72fe},
  {32'hc2774a9c, 32'h4472805e, 32'h436a7cd2},
  {32'hc458faf0, 32'hc3bc49ae, 32'h4372a409},
  {32'hc3ce70b0, 32'h44b8d49a, 32'hc4ccd442},
  {32'hc3244ade, 32'hc5080498, 32'h44a729ed},
  {32'h432dd70d, 32'hc4f00396, 32'hc2986490},
  {32'h43fe50ae, 32'h44a51cd3, 32'h44245dd1},
  {32'hc47ae1e5, 32'hc1f7074d, 32'hc498be1a},
  {32'h4435fc35, 32'h44ac32fe, 32'h42be8bea},
  {32'hc41d31ea, 32'hc3e61b57, 32'hc54672e1},
  {32'h44aec3a7, 32'hc2cbe1f2, 32'h44a63fbe},
  {32'h444a32b4, 32'h434ac060, 32'hc3a7b1be},
  {32'hc2462a5a, 32'h451cd73b, 32'h43a3ff52},
  {32'hc34cc41e, 32'hc361e3e2, 32'hc4ba2bae},
  {32'h442acf92, 32'h441e8eff, 32'h4485a0f7},
  {32'hc444e077, 32'hc3a56e3e, 32'hc412ff14},
  {32'h42ec33dc, 32'h43f19843, 32'hc212ab0e},
  {32'hc4b6e70e, 32'h43126cd5, 32'hc378146e},
  {32'h4301e110, 32'h44650cdb, 32'h442f72c5},
  {32'hc3bae18d, 32'hc4844968, 32'hc55780d0},
  {32'h449d4534, 32'h43d28a28, 32'h4407aa43},
  {32'hc3b2c686, 32'hc5654e8a, 32'h43ae767d},
  {32'h44343684, 32'h44ab3a15, 32'h443cb659},
  {32'hc528bb06, 32'h4414635b, 32'hc19bb973},
  {32'h45042676, 32'h44983c19, 32'hc29aa230},
  {32'hc3b27e38, 32'hc3b16b78, 32'hc3f60155},
  {32'h4525417d, 32'h430f44d4, 32'h436ec3d4},
  {32'hc49bcf8a, 32'h43f51000, 32'hc44cf3b1},
  {32'h453784e8, 32'hc41eb79f, 32'h440e700e},
  {32'h441437f8, 32'h4493b453, 32'hc42aed9b},
  {32'hc4567482, 32'h4433aa35, 32'h449610ef},
  {32'h44feda43, 32'h4340fb20, 32'h4388aac3},
  {32'hc37eeb92, 32'h42b4186b, 32'h454189db},
  {32'h450ba668, 32'hc391bdd0, 32'hc1009f42},
  {32'h450091e3, 32'h43df2213, 32'h426ec50e},
  {32'h453ea076, 32'h43967d47, 32'hc323c0d8},
  {32'hc3e5d375, 32'h43cbb34a, 32'h452f9ee2},
  {32'h4529e306, 32'h3fbfb000, 32'hc1c5aa20},
  {32'h444b0ccf, 32'hc42c5d0c, 32'h44e57e28},
  {32'hc3461a09, 32'hc46283ec, 32'hc4847df0},
  {32'h43c5a64d, 32'hc4f13d2d, 32'h4432f9d0},
  {32'h4528906c, 32'h42e3ef01, 32'hc4174f98},
  {32'hc512c5a6, 32'h4330332b, 32'h43ecd7f5},
  {32'hc4729267, 32'hc43fd59c, 32'hc10d3374},
  {32'hc3bf1172, 32'h44ae9ab6, 32'h44a918f3},
  {32'h43b6cf83, 32'hc398ea7e, 32'hc4b45d26},
  {32'hc34db9b4, 32'hc40b213e, 32'h44b19c63},
  {32'h43a3d1b4, 32'hc5518ab7, 32'h433437d8},
  {32'hc50ddbb2, 32'h441afad9, 32'h43b0d8c1},
  {32'h430a185c, 32'hc2dfdd77, 32'hc3621f95},
  {32'hc53ee72e, 32'hc39557f2, 32'h4189b65b},
  {32'h44619ab2, 32'hc44af7e8, 32'h43cbe651},
  {32'h44a47efa, 32'hc26b1e74, 32'h43bac39a},
  {32'h44d62f9e, 32'h4445489c, 32'hc2ddcd43},
  {32'hc52bb6b3, 32'hc2b85256, 32'hc3654552},
  {32'hc3aa387e, 32'h4337a3d6, 32'h4401218d},
  {32'h444c5a13, 32'hc2df3da1, 32'h42589903},
  {32'hc4b60bf2, 32'hc338bdd3, 32'hc4c83211},
  {32'h4507cb7e, 32'h4226c55b, 32'h432b0301},
  {32'h4365e963, 32'h44cd4287, 32'hc3c243ec},
  {32'hc28a1830, 32'hc55e2239, 32'hc26874af},
  {32'hc4b3776c, 32'h433f2627, 32'h42900458},
  {32'h43d73b6c, 32'hc4a62f5a, 32'hc2cca50a},
  {32'hc4908718, 32'h44328547, 32'h42babc2f},
  {32'h44fcce98, 32'hc475caae, 32'hc3947a53},
  {32'h443cf7b8, 32'h44482e6b, 32'h43b14d09},
  {32'h453351f0, 32'hc2bf0472, 32'h432246a2},
  {32'hc2cfaf00, 32'h44352d7f, 32'h444930be},
  {32'hc4b5d4fc, 32'hc2a00f5c, 32'hc36b4acd},
  {32'h43c20688, 32'h44814b29, 32'h43e66b82},
  {32'hc304dd46, 32'hc1a56822, 32'hc43e9982},
  {32'h43be1efa, 32'h43aa44fd, 32'h437505e3},
  {32'hc33aeea8, 32'hc52f9f49, 32'hc2b6993b},
  {32'hc2cce412, 32'h452323ea, 32'hc2333e16},
  {32'h44e19e95, 32'hbfb4a468, 32'h438b9b97},
  {32'hc49dd1e2, 32'hc43dc724, 32'h4433e54d},
  {32'h44b4b39e, 32'hc38ec884, 32'hc47ac3ca},
  {32'h4401c97c, 32'h43128b3e, 32'h4455226d},
  {32'h45004100, 32'hc3798559, 32'hc3834f28},
  {32'h426cf0d7, 32'h44073624, 32'h44e764e3},
  {32'h454cabf8, 32'h41d2c0d3, 32'h42c52aee},
  {32'hc32c6798, 32'h440090d9, 32'h4519ff2d},
  {32'h45012384, 32'hc4575688, 32'hc442bf03},
  {32'h4459f3fa, 32'h43a6d287, 32'hc32eac30},
  {32'hc55cd9a0, 32'hc364e635, 32'h414a72df},
  {32'h44bb21e0, 32'h44026e89, 32'h436f8387},
  {32'hc392ff10, 32'hc4ebfb4a, 32'h43a6f92d},
  {32'h44a58098, 32'h41528716, 32'hc3840380},
  {32'hc48bea64, 32'hc3523c17, 32'h42d30a59},
  {32'h44f57760, 32'h446dbc5c, 32'hc18e35ff},
  {32'hc4e2b7da, 32'hc4d91dfa, 32'h42da4b99},
  {32'h453a1094, 32'h43453456, 32'h43aea573},
  {32'hc31e1a1a, 32'h42ae7809, 32'h4551242d},
  {32'h44a49885, 32'h440d62e6, 32'h438f8f53},
  {32'hc32aaf26, 32'h42afb805, 32'h443d2e6f},
  {32'h445f44fe, 32'h44b30575, 32'h425cf922},
  {32'h43090f48, 32'hc3fff0f5, 32'hc462b148},
  {32'h4457acce, 32'h42ff67cf, 32'h43182560},
  {32'hc4658454, 32'hc471ce42, 32'hc3965670},
  {32'h44e13ab6, 32'h42acfd8f, 32'h441add67},
  {32'hc2cf92c6, 32'hc4193861, 32'hc40f7ebf},
  {32'h44e1f4df, 32'hc3801d60, 32'h44385c2e},
  {32'hc55b112d, 32'hc24ef476, 32'hc0c28edc},
  {32'h44a2d52e, 32'hc3a667ce, 32'hc3949de3},
  {32'hc41c0f14, 32'hc487d79b, 32'hc4ba3a53},
  {32'h448a5dcb, 32'h4246b7fe, 32'hc33be401},
  {32'hc39b237c, 32'hc1f698c1, 32'hc4c15c6f},
  {32'h43a24fff, 32'h43c2ec96, 32'h44b4bed8},
  {32'hc47e4a63, 32'hc509c471, 32'hc332c740},
  {32'hc4bcc6bb, 32'h40c6b13f, 32'h42ce20da},
  {32'hc34c5553, 32'h43be6f10, 32'hc3cb9409},
  {32'hc2a8e148, 32'hc519409d, 32'hc3821c15},
  {32'h445679bf, 32'h44a98bb9, 32'hc381725e},
  {32'h4425e246, 32'hc42cad8d, 32'hc2abd1be},
  {32'h43abf570, 32'h44f73ef0, 32'h42173dab},
  {32'hc506960a, 32'hc40572af, 32'hc30cb01e},
  {32'h44f7c7ea, 32'h41665d23, 32'hc351f8e6},
  {32'hc50b554d, 32'h436b5a4b, 32'hc305afdc},
  {32'h45686681, 32'h43963bcc, 32'h43c303ec},
  {32'hc41fc144, 32'h40f769e0, 32'h442e8902},
  {32'h43c784fc, 32'h4370e36c, 32'hc28907ed},
  {32'hc4f0daa5, 32'hc4059094, 32'hc0385375},
  {32'h43c7001e, 32'hc3cac289, 32'hc3587b0a},
  {32'hc4205d78, 32'hc29d24d2, 32'h44b9964a},
  {32'h44b39953, 32'h435557c0, 32'hc4956176},
  {32'h434243d3, 32'h43cb22b7, 32'h44ae3724},
  {32'h4519cee3, 32'hc3d6fa5b, 32'hc35be5fa},
  {32'hc514559e, 32'h4352b14a, 32'h43c3d381},
  {32'h45616e56, 32'hc38686a0, 32'hc1f73d7b},
  {32'hc47a5702, 32'hc4ef5470, 32'h449723a8},
  {32'h44d5ec7a, 32'h441ef63f, 32'hc3ba12e9},
  {32'hc2b41740, 32'hc2866d5f, 32'h4419e99a},
  {32'hc2846552, 32'h442333e2, 32'hc4e407bd},
  {32'hc53e081d, 32'hc32e3da2, 32'h43bb4670},
  {32'h454e411a, 32'hc2168ba8, 32'h43e93ebd},
  {32'hc3a54203, 32'h43e84a95, 32'h4550d977},
  {32'h457d0018, 32'h437f59ca, 32'hc3bebcfd},
  {32'h44309149, 32'hc4a19e96, 32'hc3b12566},
  {32'hc48a9886, 32'hc425b6b4, 32'h44b2c918},
  {32'hc4571bd3, 32'hc3dc4b11, 32'hc3910ae6},
  {32'hc5023d74, 32'h448016ba, 32'hc3d6f605},
  {32'h43861ff6, 32'hc2e64332, 32'hc3edeba5},
  {32'hc49002a2, 32'h436e98c8, 32'hc300a649},
  {32'h4437e4a9, 32'hc40b55b8, 32'hc49c9cbf},
  {32'hc3452bd8, 32'hbf8bfb96, 32'h440cdc5c},
  {32'h44814c86, 32'hc1be56b0, 32'h44269e2a},
  {32'hc2b341b6, 32'h4521a57d, 32'h43854976},
  {32'h430ff9c0, 32'hc55a1248, 32'h438f005a},
  {32'hc4ec6b42, 32'h42092b9c, 32'h418f7d31},
  {32'hc2cc41d8, 32'hc445067d, 32'h45001353},
  {32'hc3ebbd10, 32'h4516ac76, 32'hc3b3ff75},
  {32'h442347f8, 32'hc259de53, 32'h4262e964},
  {32'hc23fe948, 32'hc312d7ca, 32'hc55894d2},
  {32'h4389d500, 32'hc2f48519, 32'h44f4e7ec},
  {32'hc2d35204, 32'hc4320510, 32'hc4eb9e72},
  {32'h44c25262, 32'hc435310f, 32'h43b81ddf},
  {32'hc48667f2, 32'h44c85c55, 32'hc3baa32f},
  {32'h45342b57, 32'h43eb4401, 32'hc413b5b3},
  {32'hc551248a, 32'h437a32ec, 32'h42132d88},
  {32'h43c6851a, 32'hc4e204c2, 32'h4421f616},
  {32'hc4ffa345, 32'h43263145, 32'h42cc8740},
  {32'h45508e1c, 32'h439b7a8c, 32'h4395b52b},
  {32'hc41d832c, 32'hc461f17c, 32'hc5541fc8},
  {32'h44ad8181, 32'h43c1a368, 32'h42fd9024},
  {32'h436d12f6, 32'hc4521bb9, 32'hc53cffc7},
  {32'hc3889e20, 32'hc4edddc2, 32'h44d953a6},
  {32'h436469c0, 32'h448a2755, 32'hc4c71e68},
  {32'h44c270e9, 32'h4324dc28, 32'h42655b41},
  {32'h440071c9, 32'hc50412ac, 32'h43f98514},
  {32'hc4a4f1e0, 32'hc1d12ef0, 32'hc459652c},
  {32'h44461ad1, 32'hc4851fe7, 32'hc343034c},
  {32'hc47262c9, 32'h44efbd29, 32'hc378ea73},
  {32'h43a28df5, 32'hc402406d, 32'h44cd3875},
  {32'hc393248c, 32'hc47bfff9, 32'h4531711e},
  {32'hc497996c, 32'h4396461c, 32'hc4713967},
  {32'hc3a7abeb, 32'hc4c6a17c, 32'h444a6818},
  {32'h435f9e69, 32'hc4997f05, 32'hc380399d},
  {32'h4273ab58, 32'hc3a1a5c7, 32'hc51727bd},
  {32'h44006cb1, 32'h415d4825, 32'h449e0218},
  {32'h43fd25fb, 32'h43ce40af, 32'hc44ef1e1},
  {32'h447e0f58, 32'hc3bde19e, 32'h44af4a1f},
  {32'h43c70728, 32'h454e7006, 32'h427499ad},
  {32'hc3a0bb7a, 32'hc39e5426, 32'h4421d1d7},
  {32'hc53a959e, 32'hc3dfd88b, 32'h43da4557},
  {32'h44d75cfd, 32'h445fc338, 32'h441f7d26},
  {32'h450e700e, 32'h42db6085, 32'h41d56edf},
  {32'h4183f840, 32'hc522755d, 32'hc4412217},
  {32'hc4276ab5, 32'h448291a3, 32'h42f3e03c},
  {32'h437fdec6, 32'hc50bf19b, 32'h43386719},
  {32'hc4993e94, 32'h44d984c7, 32'h439bd464},
  {32'h44ab0ce8, 32'hc481be1d, 32'h4445e9e0},
  {32'hc3d9b45a, 32'h43f6ff99, 32'h44838a02},
  {32'h42e32f9c, 32'hc475d920, 32'hc48a2f19},
  {32'hc38a5a92, 32'h448f32b5, 32'h448d7492},
  {32'hc3691570, 32'hc457e7cd, 32'h448780b2},
  {32'h44f7f469, 32'hc3d3d4b0, 32'h4337b36f},
  {32'h4368a9f7, 32'hc1e7bda7, 32'h44aa7f99},
  {32'h44c898bc, 32'h442880ee, 32'hc3d77804},
  {32'hc4005687, 32'hc40574e0, 32'h4476d092},
  {32'h449418b6, 32'h41f6bf46, 32'h42c950c2},
  {32'h42bff656, 32'h4454b492, 32'hc3a3c592},
  {32'hc3a95e4c, 32'h43a97a96, 32'h4508fc49},
  {32'hc34940f3, 32'h445756e4, 32'hc50306b1},
  {32'h44afbfe3, 32'h43e266b8, 32'hc38fd23e},
  {32'hc3b468f6, 32'hc4cf2b8e, 32'hc3604c94},
  {32'h41322ad4, 32'h44c250e5, 32'h425793f6},
  {32'hc51e4ec8, 32'hc4172887, 32'h43a10fe0},
  {32'hc38d1536, 32'h43d50a94, 32'hc49c360f},
  {32'hc3620f3b, 32'hc3ccc56f, 32'hc36ee4ab},
  {32'h442dc142, 32'h430f546d, 32'hc4271b4b},
  {32'hc4a65225, 32'h438e40e4, 32'h42fc729d},
  {32'h4322ec46, 32'hc2460cdb, 32'h43127c80},
  {32'hc51bff36, 32'hc42e219d, 32'hc2b6fa83},
  {32'h4518572c, 32'h43c66373, 32'hc3b3c694},
  {32'hc3d8ff20, 32'hc41bff21, 32'h4361e86d},
  {32'h44a0a77e, 32'h44b470e0, 32'h4275f5a6},
  {32'hc3ae6618, 32'hc504b69a, 32'hc3044c65},
  {32'hc4db0c1b, 32'hc1efd4fc, 32'hc30a4002},
  {32'hc41da0f8, 32'h44982b2c, 32'h431eaf5e},
  {32'h43b0cac4, 32'h441861c5, 32'hc464e369},
  {32'h429de488, 32'hc2225678, 32'h44bc0462},
  {32'hc3f5da40, 32'hc4986b30, 32'hc2059c64},
  {32'h439539b4, 32'h451c001e, 32'h43db084e},
  {32'hc397edf1, 32'hc458481f, 32'hc5083ffe},
  {32'h445d6d45, 32'h43c5e321, 32'h43cf9938},
  {32'hc5678128, 32'h43003cef, 32'hc3f9dd86},
  {32'h43d4c464, 32'h44df99d3, 32'h44c5599b},
  {32'h43660654, 32'h44952632, 32'hc3f73275},
  {32'h43d1bcbb, 32'hc1edb3ec, 32'h44586251},
  {32'h43d98ba0, 32'hc4a6660e, 32'hc3fa53a7},
  {32'hc3b0f91a, 32'h44a5dace, 32'h433c585e},
  {32'hc52b2234, 32'hc352551a, 32'hc3d29f28},
  {32'h43bef51b, 32'h44bc1320, 32'h4444f965},
  {32'hc2485530, 32'hc3951a7c, 32'hc2c71d79},
  {32'h4522a477, 32'hc41973d6, 32'h432b7d4a},
  {32'hc3921440, 32'hc2f14cf0, 32'hc4c1a0bf},
  {32'h44c19750, 32'hc34283dc, 32'hc2355892},
  {32'hc48d6363, 32'hc4b6d062, 32'h435696ed},
  {32'h44fe39ef, 32'h44559874, 32'h4446c11d},
  {32'hc407fc9f, 32'hc393aabe, 32'hc38a85a8},
  {32'h43cf4596, 32'h44e599ce, 32'h429a2b3a},
  {32'hc5206999, 32'hc3cb835b, 32'hc349b691},
  {32'h4546c716, 32'h4359bffc, 32'h43f3aa66},
  {32'hc560e93e, 32'h42b0acb7, 32'hc2c69ed3},
  {32'h43e2ded0, 32'h432def6e, 32'h439058d4},
  {32'h446d996d, 32'hc3bb8a68, 32'hc4449120},
  {32'hc526eea6, 32'h43d66513, 32'h443d4088},
  {32'h43129408, 32'hc43ad2c8, 32'hc3eb0f53},
  {32'hc518652c, 32'h44121827, 32'h4457a16e},
  {32'hc3a47a16, 32'hc4253393, 32'hc4e1f857},
  {32'hc455d341, 32'h43d3edf2, 32'h44449630},
  {32'h43cb0d2e, 32'hc0061270, 32'hc4eb5ed2},
  {32'hc421fbbd, 32'h44dd2436, 32'h44e3906a},
  {32'h438a6030, 32'hc443799d, 32'hc3ea716d},
  {32'hc2be9004, 32'h450b5aaf, 32'h44015fe9},
  {32'h445bc6d4, 32'h4492581b, 32'hc4905499},
  {32'hc4c4da4d, 32'h43ae840c, 32'h41e74b28},
  {32'hc404cb2b, 32'hc38c2075, 32'hc5447743},
  {32'hc3d4e2b6, 32'h454f6ae1, 32'hc404a98f},
  {32'hc4140735, 32'h42f81519, 32'hc44ca2db},
  {32'hc4126ffc, 32'h44320d37, 32'h44e55486},
  {32'h44ec5f98, 32'h43376ee3, 32'h42df2836},
  {32'hc524c391, 32'h441e0210, 32'hc30b278a},
  {32'hc35b0131, 32'hc457be3d, 32'hc37f02ee},
  {32'hc55f2a94, 32'h4430df26, 32'hc3be5ea8},
  {32'h43bf1c3c, 32'hc490bd04, 32'h438b2674},
  {32'h42635282, 32'h455b4c63, 32'h43928663},
  {32'h4335665c, 32'hc437e17f, 32'hc3a6dc37},
  {32'hc4dbe2b8, 32'hc2c3bdd3, 32'h42bf0a73},
  {32'h42f75ebe, 32'hc2943c69, 32'hc3c768f0},
  {32'hc40df12a, 32'h430e8ec3, 32'hc36f9559},
  {32'hc41086f8, 32'hc20a275e, 32'hc361e760},
  {32'hc4133521, 32'h439ba6b0, 32'hc36139e4},
  {32'hc501b7c8, 32'h41944727, 32'hc40b813d},
  {32'h4499bd28, 32'hc3396439, 32'h44e874f6},
  {32'hc484697e, 32'h4327d81b, 32'hc3b923dd},
  {32'h44457fd5, 32'hc4c1e3c5, 32'hc2e98155},
  {32'h43368d34, 32'h45287b24, 32'h4468dcfb},
  {32'hc36f07fd, 32'hc452cf69, 32'h43d0ce93},
  {32'hc3c5f97c, 32'h452cfde9, 32'h4421daa5},
  {32'h43920e33, 32'hc53405c1, 32'h4364bd58},
  {32'h440e14f3, 32'hc432c064, 32'hc3dbd68c},
  {32'h4464d89c, 32'h42ae3b54, 32'h43f4af8e},
  {32'hc46c4c78, 32'hc437e529, 32'h4481e24d},
  {32'h43d26a06, 32'hc310d33e, 32'hc495af0b},
  {32'hc2c9b060, 32'h42d003c2, 32'h43c6e262},
  {32'h44000a92, 32'hc44ac2b7, 32'hc40cfdc0},
  {32'hc35cb6cd, 32'h436348e8, 32'h4346b385},
  {32'h44c62a78, 32'h43ed2ec6, 32'hc4c19595},
  {32'hc4703ebf, 32'hc43c16fd, 32'h43ff4c8f},
  {32'h44ea22b5, 32'h415ead4a, 32'h4344e660},
  {32'hc5873ebf, 32'hc26f621e, 32'hc2cc5a77},
  {32'hc20d7e00, 32'h4408eb1b, 32'hc477e519},
  {32'hc23a0b10, 32'h43e12e0e, 32'h43efc73f},
  {32'h44486cf5, 32'hc43e6168, 32'hc119ab90},
  {32'h43a059b9, 32'h44a0e3fd, 32'h449d9a26},
  {32'h453ae23b, 32'h43d4d6e5, 32'h43e90c01},
  {32'h432d9d30, 32'h44fa4ecd, 32'h44737253},
  {32'h447bcb9a, 32'hc3dbdee2, 32'hc4ebf85b},
  {32'h443474e0, 32'hc3983970, 32'hc437c4ce},
  {32'h42fb4198, 32'hc381625a, 32'h455188a4},
  {32'h44686aa1, 32'h441dda6c, 32'hc3d5be0f},
  {32'hc3ab371a, 32'hc54c80e7, 32'hc1b96253},
  {32'h4414237a, 32'h4472e8d3, 32'h43ab7026},
  {32'h4368d374, 32'hc313d7d5, 32'hc139a2ba},
  {32'h4392770a, 32'h452444c0, 32'h4406de31},
  {32'h4330c22c, 32'hc57b1513, 32'h43a4c0b8},
  {32'hc47dbdcd, 32'h4310f46c, 32'h4316eb36},
  {32'hc37c1890, 32'hc4832860, 32'h45114840},
  {32'h44057c70, 32'h4422624e, 32'h43ddac96},
  {32'h44417075, 32'h442c7f26, 32'hc3fbf2e0},
  {32'h431e1469, 32'h445432a0, 32'h4512a6cc},
  {32'hc3cc8479, 32'hc538d01d, 32'hc32040b0},
  {32'h42d71180, 32'h43c8246e, 32'h42d044a4},
  {32'hc43f690b, 32'hc2a7dc48, 32'hc3a33bf5},
  {32'h44752e45, 32'h44053373, 32'h44073f8d},
  {32'hc39bfe38, 32'h42e1d43e, 32'hc376a701},
  {32'h4411f778, 32'hc3e1f9df, 32'h43f02217},
  {32'hc4a1c6b5, 32'h437eceb4, 32'hc4a9f334},
  {32'h44daad0f, 32'h43a8273d, 32'hc3e94be4},
  {32'h43a25a64, 32'hc4f4fc0a, 32'hc3ebad83},
  {32'hc33fcdeb, 32'h4337767d, 32'h44ddf85d},
  {32'h43bfe0c7, 32'hc485e455, 32'h4275ccd6},
  {32'h42d26084, 32'h437a131d, 32'h44fcde03},
  {32'hc484d208, 32'hc48f86a5, 32'hc49a0ba4},
  {32'h4475e9be, 32'hc2eb25c6, 32'h44b43a70},
  {32'hc4be4c8a, 32'h4279d9ff, 32'hc192e692},
  {32'hc4331884, 32'hc3ef8dc8, 32'hc447056f},
  {32'hc2b77be0, 32'h449bd956, 32'h444bf4eb},
  {32'hc41a94f8, 32'hc32ca252, 32'hc2c648f0},
  {32'h442efa84, 32'h43706e0a, 32'hc40c63e9},
  {32'hc5020457, 32'hc438a943, 32'hbd60d400},
  {32'h44a13fc2, 32'hc1cde172, 32'h433a2781},
  {32'hc4fd2bcc, 32'hc2ea4db1, 32'h43a6cd5b},
  {32'h446a7843, 32'hc3d07b65, 32'h440332ab},
  {32'h43fa830f, 32'hc1899cb2, 32'h44275eec},
  {32'h4481418b, 32'h424ac0fb, 32'h44819d07},
  {32'hc4d889ff, 32'hc43e8ea8, 32'h42d3ab03},
  {32'h44177738, 32'hc17badea, 32'hc4cad69c},
  {32'h40fc8900, 32'hc4a29bba, 32'h44474e5a},
  {32'h44883f25, 32'h43df2510, 32'h42bc0a55},
  {32'hc45deacd, 32'hc38de818, 32'h4319b8dc},
  {32'hc2aad092, 32'hc344fe18, 32'hc52a215e},
  {32'hc38d1ae8, 32'h43a292d7, 32'h45522378},
  {32'h44690f48, 32'hc4423c5f, 32'hc3f46c74},
  {32'hc4222634, 32'hc476a95e, 32'h44af85f9},
  {32'hc3c5f1f0, 32'h44c11fcd, 32'hc5097eae},
  {32'h4486d00f, 32'hc362789c, 32'h4265acbe},
  {32'h443d8ee8, 32'h44a35064, 32'hc44b4223},
  {32'hc3af593d, 32'h42c5c330, 32'h45046e3c},
  {32'h43b0aad4, 32'h434bdcba, 32'hc222a958},
  {32'hc51a39a4, 32'h43be942a, 32'h441bb6b1},
  {32'h446b7d75, 32'hc40c18e7, 32'hc4cded65},
  {32'h4494ee9b, 32'hc4a92f4e, 32'hc3b2cdd9},
  {32'hc4553bd5, 32'h45375175, 32'hc2b49a24},
  {32'h44cfa260, 32'h431f1b69, 32'h43b0b3d8},
  {32'hc48c4ab6, 32'h44ea5099, 32'h43fa6102},
  {32'h442ccc20, 32'hc50db455, 32'hc38ed67a},
  {32'h4421e3f6, 32'h451c5932, 32'h42c50ca4},
  {32'h455c60a5, 32'hc41f1fce, 32'hc420a2f9},
  {32'hc5919af6, 32'h43bc2688, 32'hc405e2e3},
  {32'hc4613b2a, 32'hc2123c9c, 32'h43bf75a8},
  {32'h43109ce2, 32'hc4041d37, 32'h446ef79f},
  {32'h451b5576, 32'hc1a3710e, 32'h4395e372},
  {32'hc2e4d6fc, 32'h44e45b2f, 32'h423fd8d6},
  {32'hc1817b58, 32'hc44d4a3b, 32'h4411e0bb},
  {32'hc5252272, 32'h431663cc, 32'hc40d6ab7},
  {32'hc3f4ea82, 32'h42ef8355, 32'h4431ca07},
  {32'hc40f4dd6, 32'h42d86598, 32'hc44bbb18},
  {32'h447cedd0, 32'hc42f6b09, 32'hc34d3bad},
  {32'h448e660a, 32'h442de00f, 32'hc35ff24f},
  {32'h43b44643, 32'hc56124a9, 32'hc2f10de7},
  {32'hc4f1969e, 32'h43db11ba, 32'hc2b5652c},
  {32'h448851bb, 32'hc2c8dad7, 32'hc3bff7e7},
  {32'hc3ac51c6, 32'h44f6e595, 32'hc464be57},
  {32'h42e5e1b2, 32'hc511ea97, 32'h441a0115},
  {32'h4415f802, 32'h44b6d50a, 32'hc410ed05},
  {32'h447140bb, 32'h43ca3b92, 32'h44d42a38},
  {32'hc4b18dc6, 32'hc2feac39, 32'hc4d03e8b},
  {32'h448543fc, 32'hc2c9cb5c, 32'hc31765ca},
  {32'h43da729c, 32'hc4e92caa, 32'hc4d081ee},
  {32'hc4faf538, 32'hc3d127ad, 32'h449437e0},
  {32'hc1832f44, 32'hc3e41e81, 32'hc3665248},
  {32'hc5295c4e, 32'h42f78c01, 32'h432fd55e},
  {32'h4417986a, 32'hc46549df, 32'h42446b81},
  {32'hc433ef9b, 32'h44185811, 32'hc454bd60},
  {32'h44be6df2, 32'h42c0c9f5, 32'hc2861add},
  {32'hc54a3cc8, 32'h43dc2164, 32'hc2c48ff9},
  {32'h442edb85, 32'h43c015ab, 32'h43fcbf6a},
  {32'h45226575, 32'hc22b5299, 32'h4409ee15},
  {32'h432e6760, 32'hc4de87d3, 32'hc4d87fd6},
  {32'hc359112d, 32'h44aa3963, 32'h4443242e},
  {32'h43441c76, 32'h43842cbe, 32'hc3559457},
  {32'h43565af6, 32'hc3a7a2d7, 32'hc52c0586},
  {32'h4432fff8, 32'hc482314b, 32'hc3560764},
  {32'h4413032f, 32'h43f87794, 32'hc47155b3},
  {32'h4491fef8, 32'h42f4d5f5, 32'h44a59fb2},
  {32'hc46f5b78, 32'h437b01fe, 32'hc477146c},
  {32'h453c0f46, 32'hc42242ee, 32'h43383148},
  {32'hc4b71ea6, 32'hc29bb41a, 32'hc459cf7b},
  {32'h44035178, 32'h44182b1a, 32'hc3c53b78},
  {32'hc50e9ec6, 32'h437647b6, 32'h43ef52b4},
  {32'h44a3dec5, 32'hc453a8be, 32'hc306e795},
  {32'h43ee2282, 32'h4581daa0, 32'hc2e62465},
  {32'h4410a957, 32'hc4d0de9e, 32'h42bb43ef},
  {32'hc46471c8, 32'h44f6b17d, 32'h4348e680},
  {32'h444de2bc, 32'hc50c2fff, 32'h4354feb6},
  {32'hc3b80808, 32'hc2bc5315, 32'h43af5372},
  {32'hc421bbd3, 32'h43a361e3, 32'hc49effc7},
  {32'hc4a18979, 32'hc3256d68, 32'h4437a90d},
  {32'h42edf75e, 32'hc5208fc3, 32'h43b395fb},
  {32'h44196f5f, 32'h447c92b5, 32'h4312bad1},
  {32'h4505f351, 32'h40223b60, 32'h42d1b0db},
  {32'hc3bf086a, 32'h42dd19f1, 32'hc46fbf45},
  {32'hc4f895da, 32'hc3646416, 32'hc23fb523},
  {32'h450c6f30, 32'h43480504, 32'h442f1ae8},
  {32'h440627e3, 32'h4373b9b3, 32'hc32883b1},
  {32'h420ed2d1, 32'hc4f73180, 32'h451e3252},
  {32'h450a1016, 32'hc34ac0ee, 32'hc403b9c8},
  {32'h42b9bdf7, 32'hc354c0cb, 32'hc521950c},
  {32'hc552592f, 32'hc3fde98c, 32'h43ad302a},
  {32'h442c791d, 32'h42e41c5d, 32'hc4ba7174},
  {32'hc3dcec5c, 32'hc490bb1a, 32'h4290f1f7},
  {32'h4434424b, 32'hc2d2011f, 32'hc30e719f},
  {32'h4411c62e, 32'h43b3d857, 32'h44931484},
  {32'hbe280000, 32'h440255fb, 32'h44159d86},
  {32'hc54b4586, 32'hc32e3c4b, 32'hc20d8f5f},
  {32'h4567206a, 32'h43495960, 32'hc226a735},
  {32'hc53295fe, 32'hc47b537a, 32'h430c0c6a},
  {32'h45612fe2, 32'hc26e9b96, 32'h43516aba},
  {32'h44d75147, 32'hc2a7b650, 32'hc3a7844c},
  {32'h44f2f28b, 32'h44290a00, 32'h43a8b4af},
  {32'hc4b061b8, 32'hc48be986, 32'hc2856b8b},
  {32'hc4b96472, 32'h4332ddd2, 32'h43734133},
  {32'h43cb3c19, 32'hc4c44e9e, 32'h442ddfc7},
  {32'h43df98e1, 32'h445bf106, 32'hc4c55c18},
  {32'hc346e222, 32'hc380506c, 32'h44eb2454},
  {32'hc474909c, 32'h4377bf1b, 32'hc3bd6145},
  {32'hc32fe5d8, 32'h440c0212, 32'h44b5caa0},
  {32'hc456aaaf, 32'hc4f39b1e, 32'hc31b32c7},
  {32'hc4967684, 32'h43e24489, 32'h432ed817},
  {32'hc357dc18, 32'hc4173b9f, 32'hc5001b8a},
  {32'h44f7e06f, 32'h42f5cce8, 32'h4419979d},
  {32'hc4243c6b, 32'hc471f189, 32'h413a7eb0},
  {32'h409ab2d8, 32'h42036010, 32'h443601ba},
  {32'hc3a6d13e, 32'h442776a7, 32'hc4ce435d},
  {32'h44b93a98, 32'h4386ae23, 32'h42b0cea7},
  {32'hc3968f34, 32'hc3e7093f, 32'hc496ff83},
  {32'h4445d60a, 32'h4535c977, 32'hc305396f},
  {32'hc425e4c9, 32'h42f5beeb, 32'h43dd7d9d},
  {32'h43db38f0, 32'h4458e2b5, 32'h45044ce8},
  {32'hc4153740, 32'hc328ce0e, 32'hc4fc7f9d},
  {32'hc413d12a, 32'h4479c46c, 32'hc13432a8},
  {32'hc3fc1820, 32'hc4a3ecc7, 32'h42ed01af},
  {32'h4298c88c, 32'h458405b2, 32'h4380b8ed},
  {32'h44ab24ed, 32'hc430f19d, 32'hc34f7055},
  {32'h4407a919, 32'h44e8c247, 32'h442b3747},
  {32'hc486d34f, 32'hc4e3598e, 32'hc0fe0fce},
  {32'hc48549ad, 32'h428f22ff, 32'h438fa19b},
  {32'hc51fb855, 32'hc3a41afd, 32'h4178b32f},
  {32'h45484e91, 32'h431a7f49, 32'h43864653},
  {32'hc3135b3b, 32'hc4a4c6fe, 32'hc4197374},
  {32'h4398ebe1, 32'hc43faeec, 32'h450fe768},
  {32'hc0d51fa3, 32'h430bef98, 32'hc48e21ff},
  {32'hc436cd18, 32'h44ce6bb3, 32'h4379ebe5},
  {32'h441f8512, 32'hc4ba12c9, 32'hc34ef77c},
  {32'hc3d09a07, 32'h44b30d25, 32'h442fa324},
  {32'h4539e0df, 32'hc3a8dd12, 32'hc3c08598},
  {32'hc4cffa43, 32'h4365e6d7, 32'h44869bc3},
  {32'hc4b48317, 32'hc35af49c, 32'h423e3c6c},
  {32'hc4a3867a, 32'h440cbec3, 32'h43717ec6},
  {32'h44cc14c9, 32'h4411ec3d, 32'hc39f0c44},
  {32'h4394221b, 32'h42e58186, 32'h4409750e},
  {32'hc36ba0d1, 32'hc40b83ad, 32'h44139851},
  {32'hc3cdfc70, 32'h441da790, 32'h430a5568},
  {32'h44b5048a, 32'hc2cedae5, 32'hc431a3d0},
  {32'hc3ffa154, 32'h4498b929, 32'h4480c4f7},
  {32'h44a38f15, 32'hc4ad7bad, 32'hc482b21f},
  {32'hc51d71ba, 32'h43dcb7d9, 32'h435b6394},
  {32'h447e817e, 32'hc51af6f1, 32'h422c7504},
  {32'hc51632c2, 32'h43f2a36b, 32'h44283219},
  {32'h4361eab6, 32'hc4d7fc0c, 32'h421fe86d},
  {32'hc44cf293, 32'h450c2a27, 32'h4392aa16},
  {32'hc3531d4e, 32'hc5704d9d, 32'hc3980b79},
  {32'h44cb3c0c, 32'h433be4ec, 32'h42d46b40},
  {32'h445ef3e4, 32'h4322d3c3, 32'h436117d6},
  {32'hc4821c54, 32'h423ac087, 32'hc335100e},
  {32'h44bfbd54, 32'hc4552579, 32'hc3d37384},
  {32'h43941749, 32'h435cda53, 32'h44e3b0e0},
  {32'hc4e3e8d2, 32'h42eda9ed, 32'hc4734cca},
  {32'h44dd92d0, 32'h4382ceae, 32'h4442e068},
  {32'hc4c0dad4, 32'hc388b177, 32'h43206d9d},
  {32'h446a64c6, 32'hc50c6a14, 32'hc252ef38},
  {32'hc49bb397, 32'h4495e1ef, 32'h42fa7ad5},
  {32'hc3a69372, 32'h431a617f, 32'hc36fcaf7},
  {32'hc45e6797, 32'h45182370, 32'h4405edce},
  {32'hc3bc10d5, 32'hc578dfe0, 32'hc2d622e4},
  {32'h4402a5c1, 32'hc32e87e6, 32'hc4679dad},
  {32'h43b84af8, 32'hc2894f89, 32'hc42aefea},
  {32'hc4838a0a, 32'h44346261, 32'hc386a8c6},
  {32'hc296002b, 32'hc3fc163e, 32'hc47f4d02},
  {32'h43e3800c, 32'h449cc747, 32'h43e03ad0},
  {32'hc39dd445, 32'hc3af4d2b, 32'hc55b6935},
  {32'h42c1d37a, 32'h44463e0a, 32'h44011e6d},
  {32'h44e87eaf, 32'h43ee629f, 32'hc4a04ed6},
  {32'hc4107b7d, 32'h43c8707c, 32'h4544e422},
  {32'hc33e43a1, 32'hc3828b51, 32'hc29e8c20},
  {32'hc50d312a, 32'h444345a7, 32'h44a78d1a},
  {32'h44ac735e, 32'hc436ff90, 32'hc4995d2f},
  {32'h4480a556, 32'h43fd83f9, 32'hc34065d4},
  {32'hc3a7d7ac, 32'hc5074a5b, 32'hc27aab1a},
  {32'hc4527e71, 32'h4476ba48, 32'h41ab1627},
  {32'h44265116, 32'hc238e1f6, 32'hc4333d7f},
  {32'hc425f1a0, 32'h44c7552f, 32'hc2563338},
  {32'h4433c1bf, 32'hc345ce27, 32'hc51e3050},
  {32'h444738e6, 32'h42b88312, 32'hc3b19318},
  {32'hc3be8f89, 32'hc37c4d54, 32'h4512f152},
  {32'h448c1a04, 32'h4262b00e, 32'h4430f596},
  {32'hc5017f04, 32'hc468b4c7, 32'h4345d3ef},
  {32'h44922a00, 32'h43caeada, 32'h43cfc371},
  {32'hc3e8b376, 32'hc4883314, 32'hc2bd5831},
  {32'h432db4e0, 32'h4589f6e2, 32'h43d9bb39},
  {32'hc532b005, 32'hc3ef0310, 32'hc385842f},
  {32'hc4f4139a, 32'hc3178481, 32'h439af2e3},
  {32'hc509515d, 32'h41ceb793, 32'h43cd1a77},
  {32'h44e5d149, 32'hc35f1319, 32'hc3ca0eb8},
  {32'h450faa07, 32'hc392995f, 32'hc11fec1e},
  {32'h442fa143, 32'h440bbca7, 32'h44c5c73f},
  {32'hc44166be, 32'hc4580ff1, 32'hc5145794},
  {32'hc3e47f4a, 32'hc3483af9, 32'h44a4f912},
  {32'hc34e3f81, 32'hc2d68eb6, 32'hc524af70},
  {32'h44b34bd6, 32'h4402646b, 32'h43887de6},
  {32'h410a8200, 32'h41bcf922, 32'hc4e6917b},
  {32'hc2daee00, 32'hc42ee08e, 32'h43c7b64b},
  {32'hc564ca6f, 32'h415f22fa, 32'h43035d2e},
  {32'h4492da44, 32'hc335f72f, 32'hc3acd60f},
  {32'hc35a5ef8, 32'hc381024f, 32'hc4c9eebb},
  {32'h450efd8f, 32'h44101d88, 32'h4383e9e4},
  {32'h44ec70c2, 32'hc3ac4c0e, 32'hc1f1f444},
  {32'hc296e0cf, 32'h43f506c4, 32'h448a0bfb},
  {32'hc485e8fc, 32'hc3c80401, 32'hc46ddd59},
  {32'hc4aeb84c, 32'h432ebd58, 32'hc1c8b5ae},
  {32'hc425e505, 32'h43b91a49, 32'hc3622ab6},
  {32'hc4748344, 32'hc4937d65, 32'hc2909a8a},
  {32'h4468bfaa, 32'h44c7dec1, 32'h43d2786a},
  {32'hc51e3ad8, 32'h41e92144, 32'h43911b09},
  {32'h42f4ba9a, 32'h44e8354b, 32'hc369bfca},
  {32'hc3f75e98, 32'hc47cd5eb, 32'h43dc65b6},
  {32'h4439db07, 32'h4326a15c, 32'h433a9b8c},
  {32'hc57595b4, 32'h43ef3956, 32'h431f5047},
  {32'h44a5b270, 32'h4420c371, 32'h4209a25b},
  {32'hc4a23f81, 32'hc29b9f6b, 32'h431a9834},
  {32'h4422eda2, 32'h44956980, 32'h44059f36},
  {32'hc481e4ff, 32'hc276b048, 32'h44479bdc},
  {32'h42f2f094, 32'h4081feda, 32'hc4fee994},
  {32'h40c85141, 32'hc50a548b, 32'h42be9a56},
  {32'h43e9f677, 32'h43f5538c, 32'h4243f95c},
  {32'hc3660b3c, 32'h43d0c12f, 32'h443552a8},
  {32'h450cf70a, 32'h436ac568, 32'hc33cca94},
  {32'hc505f54d, 32'h42ac9020, 32'h44115665},
  {32'h44f92aec, 32'hc40215ba, 32'hc238b5fc},
  {32'hc48b6750, 32'hc50d1bb1, 32'h443c9119},
  {32'h44f20873, 32'h44a0e47a, 32'hc3c73715},
  {32'h43af37d4, 32'hc4cd51a8, 32'h433f3e29},
  {32'h41654a6a, 32'h43d52547, 32'hc50ee007},
  {32'hc3aba5a2, 32'h43906145, 32'h45248421},
  {32'h43532300, 32'hc390afa0, 32'hc502cea8},
  {32'hc3404fe0, 32'h43b7d558, 32'h4454b5aa},
  {32'h450e71d7, 32'hc22bed11, 32'hc43dee07},
  {32'h4436dcc6, 32'hc50da498, 32'hc3a0c330},
  {32'hc4250908, 32'h446ac041, 32'h443eca6d},
  {32'h44fcdaac, 32'h427b1b44, 32'h43f75193},
  {32'hc47da912, 32'h44882cb5, 32'hc35f9655},
  {32'h430a14e8, 32'hc539f91d, 32'hc37c6966},
  {32'h4470c539, 32'h443c620a, 32'h42392446},
  {32'h455a175a, 32'h43061660, 32'hc28b82f2},
  {32'hc48230a0, 32'hc395cc68, 32'h416ab8a0},
  {32'h44de7e69, 32'hc267de90, 32'h4400fd4f},
  {32'h4392685a, 32'h44ea9161, 32'hc346d6cc},
  {32'h43a1082d, 32'hc43cc3c3, 32'h44a7f9f4},
  {32'h4438d744, 32'h447999bf, 32'h43019ea6},
  {32'hc210ddb0, 32'hc395e84e, 32'h44fb8d1d},
  {32'hc30d7d38, 32'h438380bb, 32'hc4e6b5a6},
  {32'h44096c81, 32'hc33557d4, 32'h44060cd5},
  {32'hc2bd6c20, 32'h42c563bc, 32'hc3992f89},
  {32'h450b858a, 32'hc43ce15b, 32'h431faba6},
  {32'h43ad24ae, 32'h4299c95e, 32'hc49b0584},
  {32'h451e45c2, 32'hc3b7cc22, 32'h43a74eab},
  {32'hc4862142, 32'h448f7ef1, 32'hc32f2e67},
  {32'hc3b6f9bd, 32'hc4df25ad, 32'h4147067d},
  {32'hc259d6a0, 32'h44d3b969, 32'hc4483a1b},
  {32'h4473a68b, 32'hc5044bac, 32'hc3eff9e0},
  {32'hc2fbe1ae, 32'h44b6b179, 32'hc39ae5c2},
  {32'h43a8a00a, 32'h43d48408, 32'h443b30a5},
  {32'hc31125ca, 32'h4397103b, 32'hc4d8430d},
  {32'h4516fc88, 32'hc3a1e880, 32'hc3224fbf},
  {32'hc32955e0, 32'hc3878bb8, 32'hc4e7994a},
  {32'h44f9c222, 32'h43874acf, 32'h4370b773},
  {32'h42f75ed7, 32'h44897c2b, 32'hc44a1b84},
  {32'hc4e2746a, 32'h439d7c0c, 32'hc2084287},
  {32'h436e0421, 32'hc42d4248, 32'h44a383db},
  {32'h42aa62b2, 32'h45130a0a, 32'h43804fb7},
  {32'h44b21078, 32'h432e69f5, 32'hc16b2d1a},
  {32'hc50b8f1e, 32'h432ceade, 32'hc3df330d},
  {32'h451a580d, 32'hc3bbaf98, 32'h43c26fdc},
  {32'h4421d902, 32'h44427184, 32'h4489f124},
  {32'hc381bf90, 32'h442442cc, 32'hc4bdcf16},
  {32'hc40a68cd, 32'h44795284, 32'h431f5925},
  {32'hc323f13c, 32'hc4a2615b, 32'h4226570e},
  {32'hc4ec24a6, 32'h441037d2, 32'h433530cc},
  {32'hc274d71a, 32'hc537b8e6, 32'hc3ee98ea},
  {32'h431c0065, 32'h44e59bbd, 32'hc28726dd},
  {32'hc34bf787, 32'hc55516b3, 32'hc3c11637},
  {32'hc3f697e7, 32'h44521204, 32'hc3782921},
  {32'h4477f058, 32'hc40a3f98, 32'h42b341fc},
  {32'hc5110d1c, 32'hc3aab6a6, 32'hc34a77ea},
  {32'hc1fc6058, 32'hc3bcd532, 32'hc23c7098},
  {32'hc24867a2, 32'hc300274b, 32'hc3a429d8},
  {32'h44836866, 32'hc4b33337, 32'hc2a17db1},
  {32'hc2967c00, 32'h4418bf9c, 32'hc41ed70f},
  {32'h4354d85f, 32'hc4f8498b, 32'hc38fac76},
  {32'hc44edbb4, 32'h451bdc30, 32'h431da914},
  {32'hc3821adb, 32'hc55ce8df, 32'hc292869c},
  {32'h4473b398, 32'hc3d83511, 32'h440d184d},
  {32'h446e5a46, 32'h4476a8ef, 32'hc3eb1c42},
  {32'hc3202108, 32'h43bbb3f4, 32'h4479d1f2},
  {32'hc3daf29a, 32'hc45b10cd, 32'hc33e12f8},
  {32'h449e8ee3, 32'h4393d895, 32'hc3a84d89},
  {32'hc3da1fc6, 32'hc24d494b, 32'h447af55d},
  {32'h44138c17, 32'h4504b2e0, 32'h42ffbb82},
  {32'hc49e9f35, 32'hc3237a27, 32'hc2f047c6},
  {32'h4464d668, 32'h449555aa, 32'h43a8b72b},
  {32'h4527af78, 32'h41d989f0, 32'h43fce91a},
  {32'hc3704bb8, 32'hc4e13d3d, 32'h44f265a8},
  {32'hc40a0a59, 32'h449257a1, 32'hc51f572c},
  {32'hc1fbb8d8, 32'h447532e8, 32'hc48058ec},
  {32'hc2af34f8, 32'hc4e35539, 32'hc2e23da6},
  {32'h43e4243c, 32'hc28900ed, 32'hc4097137},
  {32'hc4466396, 32'hc480ac0b, 32'h446a1976},
  {32'hc3f866c2, 32'hc421a033, 32'hc5517c01},
  {32'hc405a93e, 32'hc3088d40, 32'h4408a056},
  {32'h45222988, 32'hc32834ef, 32'hc378ccf2},
  {32'hc5823518, 32'hc3be21a3, 32'h4450dcd7},
  {32'h44ed8c28, 32'h437e51b1, 32'hc39ec4a8},
  {32'h439dfe6b, 32'hc56218e7, 32'hc299237c},
  {32'h44eb30f4, 32'h4388818a, 32'h4258f933},
  {32'hc525d576, 32'hc379329a, 32'hc36b04af},
  {32'h450bc855, 32'h4456a81d, 32'hc38e9aa3},
  {32'hc53b349e, 32'hc354bbdc, 32'h43447cd9},
  {32'h44ce5819, 32'hc3358019, 32'hc0c0ad0c},
  {32'h44ce7336, 32'hc42e4723, 32'hc32a1188},
  {32'hc40802ea, 32'h44ed628f, 32'hc4c1805c},
  {32'hc25fe0c4, 32'hc44a0fc9, 32'h44a1ade9},
  {32'hc39abbd3, 32'hbebb12a0, 32'hc48af7ac},
  {32'h44d14f9a, 32'h441d36a4, 32'h43331574},
  {32'hc41e6b25, 32'hc3938300, 32'hc51c354d},
  {32'h447cd56b, 32'h44178ff0, 32'h43b277b6},
  {32'hc4c12c8d, 32'hc3b3a731, 32'hc46099f8},
  {32'h451983b3, 32'h43a8f8e2, 32'h43ff8ada},
  {32'h43007a29, 32'hc2bb1f14, 32'hc42b0ff1},
  {32'h437437a4, 32'hc3b8251f, 32'h44aaba96},
  {32'h4407cd56, 32'hc461e234, 32'h41880206},
  {32'hc4a25261, 32'h43d96f18, 32'hc360eebc},
  {32'h425177b0, 32'hc4942026, 32'hc48ead5e},
  {32'h4495eb88, 32'h445a821d, 32'h4242d224},
  {32'h44288706, 32'hc3d6b070, 32'hc2d4c958},
  {32'h442a031f, 32'h44817e07, 32'h44833c31},
  {32'hc4335962, 32'hc3a084c7, 32'hc45f621a},
  {32'h449a1450, 32'h4440bf26, 32'h4350b667},
  {32'hc44d5aac, 32'hc4ace6f0, 32'hc41c5f5a},
  {32'h43e6a1dc, 32'h453c60cd, 32'h430ff3f9},
  {32'hc2559bda, 32'h423e0dd1, 32'hc1c01ab8},
  {32'h44926b76, 32'h449e37fb, 32'h41e668a8},
  {32'h431a58a4, 32'hc54baed6, 32'hc3a7e596},
  {32'h450e2cd2, 32'h422f4c11, 32'h442d057b},
  {32'hc51b83b5, 32'hc25ab545, 32'h4198810e},
  {32'hc3518c6c, 32'hc3fb90dd, 32'hc4629547},
  {32'hc392426a, 32'hc4e2634c, 32'hc3658f2e},
  {32'hc3d9c80e, 32'h43abe17d, 32'h43d0180a},
  {32'hc4439e57, 32'h44143789, 32'hc4375001},
  {32'hc3e85c0c, 32'h45332f8b, 32'h42726fa0},
  {32'h4302d4ad, 32'hc4909b09, 32'hc3082394},
  {32'h4495465c, 32'h440661a6, 32'hc29ec94d},
  {32'h42c2d8e8, 32'hc4157fde, 32'hc55f34ae},
  {32'hc5681d22, 32'hc0c33c10, 32'h43434895},
  {32'h447081bf, 32'hc403a465, 32'h42c3fac1},
  {32'h43b32652, 32'hc509f9df, 32'h44f0138c},
  {32'hc366dd33, 32'hc558cba9, 32'hc3e3c12b},
  {32'h443adcdd, 32'h435068f6, 32'h43198fde},
  {32'hc3c06043, 32'hc52ca921, 32'hc3bc6172},
  {32'hc40a7a96, 32'h43f07d1a, 32'h43063d7d},
  {32'hc256f218, 32'hc054ece8, 32'hc44c1dce},
  {32'h42d7a240, 32'h44618bec, 32'h44b93c1e},
  {32'h42a4e7e0, 32'h42916fcd, 32'hc458ca9e},
  {32'h43bd071c, 32'h43d583e6, 32'h4449eb91},
  {32'h4414fc53, 32'hc557af40, 32'hc238f97c},
  {32'h430c54a4, 32'h4585f9ed, 32'h42f0189e},
  {32'h44b629c9, 32'h42699ecd, 32'hc31f3848},
  {32'h40942e10, 32'h44db7d6e, 32'h43125893},
  {32'h454ee9c8, 32'hc3ae111a, 32'h418a8a20},
  {32'hc5474091, 32'h41e3128c, 32'h423aa50d},
  {32'h4566be07, 32'h43ae960f, 32'h43c31460},
  {32'hc58a470b, 32'hc393c0c5, 32'hc369d95c},
  {32'h44193b50, 32'hc42c8c90, 32'hc3ebc8c9},
  {32'h42353358, 32'hc3b354d7, 32'hc3178a6f},
  {32'hc54e220e, 32'h43a23f70, 32'h431b9c8f},
  {32'h439ebac1, 32'h4382bc1a, 32'h451c9a75},
  {32'h431a4b78, 32'h449c55cc, 32'h424fa2de},
  {32'h4501df30, 32'hc4709719, 32'h438ad131},
  {32'hc338c611, 32'h44f67081, 32'hc282f69c},
  {32'hc4e3a0ec, 32'hc3e5ff7f, 32'h4351134b},
  {32'hc4f02666, 32'h44b77d01, 32'h430d6cfa},
  {32'h451c1250, 32'hc3dd3d0b, 32'hc2ca3c96},
  {32'h45031ac5, 32'h41a8c2c8, 32'h42b0d5a0},
  {32'h44e6ac7c, 32'hc147c77a, 32'h4403b7fb},
  {32'hc4a880f5, 32'h445350a0, 32'h443b8b0e},
  {32'h44cdac4e, 32'h42cbb2ef, 32'hc2d273fc},
  {32'hc38d4139, 32'h4304d425, 32'h44a3e35f},
  {32'hc3795b4b, 32'hc3a3907a, 32'hc50be0ab},
  {32'hc42504a7, 32'h4471d2e2, 32'h423f5817},
  {32'hc328c1ca, 32'hc4e224d3, 32'h4324b5b3},
  {32'hc5092264, 32'hbe40dd00, 32'hc398849b},
  {32'h457643ba, 32'hc3f9dd3e, 32'h433af04c},
  {32'hc514b1f0, 32'h444c60f9, 32'h42b37fca},
  {32'h4558bd8d, 32'hc3ceba4b, 32'hc3e9aca6},
  {32'h446c27a8, 32'h4439e3ee, 32'hc1f29e18},
  {32'h438afcb0, 32'hc37957ec, 32'hc5429892},
  {32'h42bd05d0, 32'h443ab97f, 32'h4506c56b},
  {32'h4281e558, 32'hc40560e7, 32'h4344049d},
  {32'hc4fd493b, 32'h437bffa5, 32'h4332093b},
  {32'h43630588, 32'hc515dc61, 32'hc4260ca1},
  {32'h450b1343, 32'h42cbe92e, 32'hc41bf044},
  {32'hc51204fe, 32'hc32d8e2d, 32'h4406ab45},
  {32'h43b93a66, 32'h443506b7, 32'hc48bed0f},
  {32'hc4afa0e0, 32'hc4d9de34, 32'hc421a809},
  {32'h4388f8a9, 32'h44f489d4, 32'h4422b41e},
  {32'hc4ea96ea, 32'hc27aa816, 32'hc3b18fe0},
  {32'h4409bc44, 32'h4566aa69, 32'hc3404b34},
  {32'hc4d276cc, 32'hc48c6dd2, 32'hc3e0cd35},
  {32'h44fa0ab4, 32'hc38eb397, 32'h43b148a6},
  {32'hc4c32090, 32'hc2ec4227, 32'hc20f59ec},
  {32'h443a064b, 32'h430a0ff6, 32'h440f5e16},
  {32'hc4e41094, 32'h4321c734, 32'h43dc3bc4},
  {32'h44f8448e, 32'hc329e9d4, 32'h430ed538},
  {32'hc5457b80, 32'hc3f88442, 32'hc3b8ced7},
  {32'hc4003ce5, 32'hc171a58a, 32'h443cc2cd},
  {32'hc3a10254, 32'h4213c70a, 32'hc53924ac},
  {32'h449a40a6, 32'h441b99d9, 32'h42d0fd47},
  {32'hc5440bb2, 32'hc411d117, 32'hc2e8f35c},
  {32'h448180fc, 32'hc3aa0438, 32'h41df4a49},
  {32'hc5855996, 32'h4354f385, 32'hc3066c12},
  {32'hc241d920, 32'h43ef6804, 32'hc36612bf},
  {32'h427fa578, 32'hc55323e2, 32'hc34e63a1},
  {32'h43c16764, 32'h4350e934, 32'h44c7dbed},
  {32'h437220dc, 32'hc4081a89, 32'hc42f013d},
  {32'hc3a71e95, 32'h42cc341e, 32'h44b6ca23},
  {32'hc509eba0, 32'hc42f6e14, 32'hc4694192},
  {32'h43cbd710, 32'hc39ceb38, 32'h4489e868},
  {32'h45093a8b, 32'hc392cd84, 32'hc3ef6b95},
  {32'hc468222e, 32'hc48f53cc, 32'hc3af5dac},
  {32'h452e88d6, 32'h4251bfc1, 32'h44231d80},
  {32'h44596159, 32'h43028b03, 32'h42f10dfc},
  {32'h449ce709, 32'h449524cb, 32'h42e52800},
  {32'hc3455c2c, 32'hc50911a2, 32'hc2008475},
  {32'hc4e6d8c6, 32'hc1cbde74, 32'hc3437d91},
  {32'hc5327a62, 32'hc3a58ab3, 32'hc3926df1},
  {32'h42bd5723, 32'h443906ef, 32'h4454f54e},
  {32'h41cc5101, 32'hc4db3b22, 32'hc2b9021a},
  {32'h438f34fd, 32'h43f01155, 32'h43bb775e},
  {32'hc4baeae6, 32'hc2ebbd06, 32'hc31e9666},
  {32'h451ec33a, 32'h430a1d42, 32'h44153f34},
  {32'hc46fa796, 32'hc438de79, 32'h43f8d0be},
  {32'h44cbca89, 32'h4464ce82, 32'hc3f4d9e0},
  {32'h44c82279, 32'hc395728a, 32'h434d2756},
  {32'h440e9581, 32'h42da0d0b, 32'hc4ccd955},
  {32'hc44e6c8d, 32'h439fd054, 32'h42ff69f3},
  {32'h4403fb77, 32'h443136ab, 32'h428f645a},
  {32'hc4dc9adc, 32'hc4cac8ca, 32'h42bd1b82},
  {32'h45594ea0, 32'h440d20ac, 32'hc37bba17},
  {32'h43abeae8, 32'h421d9b16, 32'h42cca059},
  {32'h433cf37c, 32'h4344c0a9, 32'hc4665446},
  {32'hc463a7ea, 32'hc3324c39, 32'h44444b74},
  {32'h4244d43f, 32'hc38f6f91, 32'hc5012f75},
  {32'hc5621169, 32'h42a04b3b, 32'h412ef4fb},
  {32'h43c0d70f, 32'hc4761282, 32'hc511a79e},
  {32'h44c50d30, 32'hc408ebc4, 32'hc4130c9d},
  {32'hc563995f, 32'h43910a80, 32'h42a67f8f},
  {32'h436ee632, 32'hc4f4b780, 32'hc3107015},
  {32'hc3fce048, 32'h433086fc, 32'hc303590c},
  {32'h449f3bae, 32'hc459937d, 32'hc356c49e},
  {32'h44ba3f7e, 32'h43b5f2d5, 32'hc3b7d4a4},
  {32'h44cf499c, 32'hc2dc1e6b, 32'hc4a0e2a2},
  {32'hc52c6166, 32'h4426b908, 32'h43f1da76},
  {32'h443a9123, 32'hc2dd36f6, 32'h443ea0b2},
  {32'hc48c4cda, 32'h44c3e029, 32'hc38b408f},
  {32'h43dab7d7, 32'hc43e77b7, 32'h448a4ec7},
  {32'hc31808a2, 32'h44cfff3d, 32'h4201c829},
  {32'h443932d2, 32'hc4ef3fcb, 32'h41585032},
  {32'hc4adf200, 32'hc2d3a02f, 32'hc3a62008},
  {32'hc23666a0, 32'hc34cc8d9, 32'hc2e36b24},
  {32'hc28b0dec, 32'hc3611507, 32'hc557342e},
  {32'h450dedfb, 32'h437339fb, 32'h4226387a},
  {32'h44ca5b26, 32'hc2be0022, 32'hc407b858},
  {32'h444f33ee, 32'hc41edd5d, 32'h44fdcf7e},
  {32'hc51885c0, 32'hc350b31d, 32'hc3626fa4},
  {32'h44335edf, 32'hc4890c7b, 32'h44756f06},
  {32'hc36f73ed, 32'h45188751, 32'hc2b4a4ba},
  {32'h45460bac, 32'h4433360a, 32'h427a9a1a},
  {32'hc42b4cc6, 32'h445f4121, 32'hc49639c0},
  {32'h44b9fc1a, 32'h43f0d7f8, 32'h444cfcdb},
  {32'hc4942db4, 32'h43bd75e5, 32'hc4d516d5},
  {32'h441def1e, 32'h432239a9, 32'hc34d5e08},
  {32'hc13966b0, 32'h4398df50, 32'hc509dd4d},
  {32'h4300c234, 32'hc417b7ae, 32'h44a78034},
  {32'h448d032b, 32'hc36bfca6, 32'hc3c3191a},
  {32'hc4e93034, 32'h4221bbb6, 32'h423b443d},
  {32'h44653656, 32'h3e384200, 32'h44c51efc},
  {32'hc40805d0, 32'h43928e97, 32'hc3987b33},
  {32'h43e1c499, 32'hc361edce, 32'h42934c01},
  {32'hc53f1aef, 32'h4306a138, 32'hc3f26420},
  {32'h4459a1a8, 32'hc4d962de, 32'h43ad4e2d},
  {32'h448b82ea, 32'hc494d510, 32'h448043e7},
  {32'hc400a810, 32'h4392d91e, 32'hc3a99f6b},
  {32'h44a0d630, 32'hc434fd7e, 32'h44220cff},
  {32'h44be0577, 32'h42ed762a, 32'hc383d646},
  {32'hc4c40ab0, 32'h42f32e02, 32'hc3ead27e},
  {32'hc38897a0, 32'hc4cf422d, 32'h44131636},
  {32'hc43351ec, 32'hc35eaf98, 32'h439d3ff5},
  {32'h4411539e, 32'h426a6229, 32'h44edb988},
  {32'hc353c874, 32'h43977539, 32'hc4d8f4c2},
  {32'hc47661a0, 32'hc2950eb1, 32'h435ac9fe},
  {32'hc59610f7, 32'hc3dc214c, 32'hc3026f6e},
  {32'h44cd4fac, 32'hc2bad3f6, 32'hc41dae27},
  {32'hc438858c, 32'h44541a8b, 32'hc2b9e00c},
  {32'h4365b548, 32'hc519544c, 32'hc2d1c8ab},
  {32'hc4d498e8, 32'h442c5a8a, 32'h43e8bfdf},
  {32'h4430c6cf, 32'h439c49ad, 32'h4299025c},
  {32'hc46c8e90, 32'h44f9b60f, 32'h43f084fb},
  {32'h44f17e8b, 32'hc4a6c96f, 32'hc31ed932},
  {32'hc3050394, 32'hc433f988, 32'h417dfeb8},
  {32'h43c8993e, 32'hc34218a3, 32'hc46df3b0},
  {32'hc3743662, 32'hc3a61cd2, 32'h4490e120},
  {32'h427c5ed5, 32'hc4f8f6cb, 32'h4317d849},
  {32'hc3b3960b, 32'hc24fa883, 32'hc53b6917},
  {32'hc4b9b69e, 32'hc30d156d, 32'hc40cb048},
  {32'hc3d2c78b, 32'h453a1565, 32'hc23cf95c},
  {32'hc32979bd, 32'hc4829aae, 32'h44a5f9a2},
  {32'h436424c6, 32'h44390d5d, 32'hc4673b96},
  {32'h43c1f526, 32'h440e21b7, 32'hc1db4f9d},
  {32'hc30ed100, 32'h44996ee8, 32'h44b6b2a1},
  {32'h420e1fa2, 32'hc4e42c62, 32'hc4fd7005},
  {32'h4489db6a, 32'h43b72d73, 32'hc41429fe},
  {32'hc4f29624, 32'hc3d229dc, 32'h4239344e},
  {32'h430fb004, 32'h4300b985, 32'h4400410c},
  {32'hc3f1c0fc, 32'hc465d376, 32'h440b9872},
  {32'h44f984fd, 32'h43eadefc, 32'hc2a16b15},
  {32'h44368b0b, 32'hbfbde838, 32'h4448001e},
  {32'h45209bcb, 32'h43b36d57, 32'hc3257145},
  {32'hc594a8c4, 32'hc3908400, 32'h42ecbeb0},
  {32'h451023cb, 32'h4400f2fb, 32'h4346adf0},
  {32'hc49867e6, 32'hc4008517, 32'hc364fb54},
  {32'h42ff0e5a, 32'h450bf0f1, 32'hc397eca1},
  {32'hc3d00b24, 32'hc31c985a, 32'h42764485},
  {32'hc289e6f4, 32'h44a9ca0c, 32'h42c0469b},
  {32'h43b40c3a, 32'hc5596a11, 32'h42f6dc1c},
  {32'hc465413e, 32'hc238d21f, 32'hc413752f},
  {32'h42a22b66, 32'hc42103e2, 32'h448517ec},
  {32'hc491f860, 32'hc438b73e, 32'hc4643c00},
  {32'hc3851a23, 32'hc4f6c724, 32'h44cc0d75},
  {32'h4463ad9c, 32'h429ea1ac, 32'hc496d477},
  {32'h4414d611, 32'h43fbd3e7, 32'h451c3917},
  {32'hc2c9acca, 32'hc51b229b, 32'hc42db3c0},
  {32'h451840aa, 32'hc089b4db, 32'h42a80252},
  {32'hc34770c8, 32'hc45fde52, 32'hc4be4fab},
  {32'h44211e91, 32'h44aea1b0, 32'h44862372},
  {32'h438340f2, 32'hc498fcad, 32'h442b8708},
  {32'hc3609f6b, 32'h447301f5, 32'h443b47c5},
  {32'hc3c77e44, 32'hc4ae7e13, 32'hc44cdb9c},
  {32'hc3f5ed06, 32'h4458314e, 32'h429b20f7},
  {32'h4293ff00, 32'hc3f8a76a, 32'hc4fcd0aa},
  {32'h43d5c823, 32'h45503562, 32'hc3a726c9},
  {32'h445e3e18, 32'hc20fbc57, 32'h42d4ae3f},
  {32'h425d6c68, 32'h4441624e, 32'h450b1dfc},
  {32'hc421d27a, 32'hc4a2c1e1, 32'hc4f06772},
  {32'h44613337, 32'h42198793, 32'h443e6ec4},
  {32'hc29aaf20, 32'hc55f7519, 32'hc3987eba},
  {32'h43709418, 32'h45370568, 32'h43fce855},
  {32'h44ca021a, 32'hc359bc75, 32'hc39680fb},
  {32'h440c7a3b, 32'h4503046b, 32'hc2525109},
  {32'hc2b4c550, 32'hc5460482, 32'h42ad7cb1},
  {32'h44c78fc0, 32'h426247a4, 32'h4407b9cf},
  {32'hc4230280, 32'hc3c1a0f2, 32'h41c11885},
  {32'h45298322, 32'h42896135, 32'hc21a1fb1},
  {32'h43ac8b52, 32'h44910106, 32'hc4d5d5a9},
  {32'hc34bb8e8, 32'h44ceb16d, 32'h437f624c},
  {32'h44437034, 32'h43dc0182, 32'h43b44c24},
  {32'hc2593130, 32'h4396a91e, 32'h4500f0c9},
  {32'hc31df19c, 32'hc3c40239, 32'hc3cfb726},
  {32'hc40a778c, 32'h4354625c, 32'h448b2e06},
  {32'h43d6e022, 32'hc509baae, 32'hc4ef9cec},
  {32'hc55b8c78, 32'hc3367558, 32'h4389455c},
  {32'hc3c851e2, 32'hc432c496, 32'hc382ac38},
  {32'h43bebfa6, 32'hc4808dda, 32'h44f793d3},
  {32'h4405627a, 32'hc49b8716, 32'hc3b85e57},
  {32'hc300d85c, 32'hc4875281, 32'h43fc11a7},
  {32'hc31b8573, 32'hc4df7777, 32'hc3f9a579},
  {32'h43a99746, 32'h42afbfe2, 32'h4514f9a3},
  {32'h4498d307, 32'hc40ae6d4, 32'hc29f2507},
  {32'hc510f757, 32'h4219a8c2, 32'h43f6da7f},
  {32'hc2ba8e27, 32'h435ede05, 32'hc52272ba},
  {32'h448c1b6a, 32'h430965a6, 32'h43ddd2a6},
  {32'h450d8f28, 32'hc42b26e9, 32'hc210b4cf},
  {32'hc5914589, 32'hc357ec64, 32'hc3c7ace3},
  {32'h4521a2dc, 32'h44227a71, 32'h43b273e8},
  {32'hc46fcc58, 32'h4521b640, 32'hc3b82721},
  {32'h444634da, 32'hc4317c49, 32'h439a4e09},
  {32'hc52ce734, 32'hc3839b89, 32'hc3087823},
  {32'h4524e51d, 32'h4369dfd5, 32'h42ed1815},
  {32'hc4ce6580, 32'hc2f5048f, 32'h43adbc9a},
  {32'h4476741f, 32'hc3221ea8, 32'hc3876fa8},
  {32'h44888952, 32'hc2f10026, 32'hc085e3a2},
  {32'hc50d691e, 32'hc1ff63e7, 32'hc38fc33e},
  {32'h452d2791, 32'hc1ca708b, 32'h435fa8ac},
  {32'h44d76380, 32'h432ce02d, 32'hc2b847f8},
  {32'h3f705400, 32'hc5245bca, 32'hc353b850},
  {32'hc454da5d, 32'h44d77e79, 32'h4427f99f},
  {32'hc3099750, 32'hc3cf4152, 32'h42e0739a},
  {32'hc58d4c0b, 32'hc38fdcb4, 32'hc29f15c5},
  {32'h45142ef5, 32'hc3dc0cd1, 32'h44544c5c},
  {32'hc3858180, 32'h42cca196, 32'h438d32be},
  {32'h41f7aa80, 32'h41dd5be1, 32'h450dddb0},
  {32'hc4d68516, 32'h43c57c7e, 32'h43c31709},
  {32'hc24279a0, 32'h408c8744, 32'hc48b851d},
  {32'h4416fe94, 32'h44b3f10b, 32'h44809e4f},
  {32'h44082f78, 32'hc451efe4, 32'hc3e6d00f},
  {32'hc4432de5, 32'hc2cda05b, 32'hc336ca39},
  {32'h445e6e42, 32'hc48b3642, 32'h4222601e},
  {32'hc4bd63e7, 32'h442fe2a7, 32'hc23c285d},
  {32'h450c4fd9, 32'hc3a1a723, 32'hc3a204b5},
  {32'hc567bbc5, 32'h4408da7a, 32'h435b3494},
  {32'h44b88e18, 32'hc3d2f8b7, 32'hc45066c6},
  {32'hc2a577e5, 32'h42e8ed3d, 32'h44ea6a25},
  {32'hc2bc9dd0, 32'hc3f1f2ae, 32'hc511ab0c},
  {32'hc311ae2a, 32'h43f8651b, 32'h444c2cdb},
  {32'h43de2188, 32'hc3d37bb0, 32'hc4bf277d},
  {32'hc4e7a07b, 32'h43873c99, 32'h423d9e3b},
  {32'hc375754c, 32'hc561a9cf, 32'h42383b2c},
  {32'h431f6e70, 32'hc2857d94, 32'hc4a0ceb5},
  {32'hc4fdffeb, 32'h43805a23, 32'h44bd2ca9},
  {32'h4549e0a6, 32'h419379fd, 32'h43d25a9c},
  {32'hc448c3b6, 32'hc4ee1284, 32'hc2757928},
  {32'h441433a0, 32'h44821a4e, 32'h43d433a4},
  {32'h446e2b0c, 32'hc415508d, 32'hc38ba9f3},
  {32'h44038d34, 32'h44fae6e3, 32'hc39b947c},
  {32'hc395d03e, 32'hc556b81a, 32'h44033b88},
  {32'h43c24f86, 32'h45016152, 32'h42cd28aa},
  {32'hc4524ebe, 32'hc489c998, 32'hc46e9f12},
  {32'h44444e48, 32'h44253da4, 32'h442fbdde},
  {32'hc419316a, 32'h41b4aa2a, 32'h44dfec82},
  {32'h438b5ff2, 32'h438a8548, 32'h45165017},
  {32'hc3af776d, 32'hc48b91cf, 32'hc5038aae},
  {32'hc2b8d800, 32'h43a9d5a4, 32'h45084105},
  {32'hc4d9efc0, 32'hc37026b8, 32'hc4473191},
  {32'h42a14210, 32'h44acdd77, 32'h4437ea5e},
  {32'hc4eb670e, 32'hc4317623, 32'hc2e85170},
  {32'h45099055, 32'hc21d359e, 32'h4468ad56},
  {32'hc49efe60, 32'h4434a745, 32'hc4101b6a},
  {32'h44e89269, 32'h44455e71, 32'hc3d6fe42},
  {32'hc39a57bd, 32'hc4b6825e, 32'hc4adec49},
  {32'h44bc5bb7, 32'h44815972, 32'h444fbd9b},
  {32'hc4e14e93, 32'hc3d1ac01, 32'h42f0ab7c},
  {32'hc2552e10, 32'h44d582ce, 32'h44305fd5},
  {32'hc3e698b6, 32'hc312af2f, 32'hc54fb6fd},
  {32'h44adb6fe, 32'hc379b402, 32'hc3a5642e},
  {32'h441c213a, 32'hc3d1d230, 32'h44097412},
  {32'hc426e57d, 32'hc49d006d, 32'hc2968d9b},
  {32'h43249551, 32'h44411fcc, 32'h42a76b9b},
  {32'hc4a48a5b, 32'hc2dcb8bd, 32'h432857f0},
  {32'h450a90a0, 32'h442214d3, 32'h430f0069},
  {32'hc4284881, 32'hc4e4c927, 32'h4315457b},
  {32'h43924554, 32'h432305e8, 32'hc3507e4a},
  {32'hc46ff7a0, 32'h4326ad6e, 32'hc01c3e2a},
  {32'h437bbb2c, 32'h43fce5df, 32'hc344bf9f},
  {32'hc0902bc0, 32'h44022703, 32'hc409c033},
  {32'h43b5b19b, 32'h4424b207, 32'hc4e3157c},
  {32'hc403bc6a, 32'hc3bf277b, 32'h44e1f4a5},
  {32'hc39357fa, 32'h4496d242, 32'h427b0c1f},
  {32'hc33fa8a6, 32'hc3a3d832, 32'h44963ccd},
  {32'h4447c01e, 32'h44a4cad2, 32'hc39cdc04},
  {32'hc3c5882c, 32'hc044ce62, 32'hc3d51ffe},
  {32'h429ca5bf, 32'hc2a846bb, 32'hc51f01d5},
  {32'hc4a0dea6, 32'hc31708be, 32'h441923b5},
  {32'h447f6bb2, 32'hc2432f02, 32'hc38ac882},
  {32'hc4e0bdf7, 32'hc3d35b4b, 32'h44b511ef},
  {32'h42501b40, 32'h445479c8, 32'hc4f1b594},
  {32'hc4c53912, 32'hc3c8fc7f, 32'hc3db95d3},
  {32'h41597a80, 32'h452ccbd0, 32'h422bbabb},
  {32'hc5259cc8, 32'h42f8b4e0, 32'h41eee8c0},
  {32'h45163ffe, 32'hc254b06e, 32'hc3902392},
  {32'hc3cdb288, 32'h440239e2, 32'h4539b503},
  {32'h4536cc75, 32'hc1350131, 32'hc46b296b},
  {32'h4410a4df, 32'hc4d3add3, 32'hc3cea13b},
  {32'hc4e68bd6, 32'h437a08f5, 32'h440162d1},
  {32'hc4d1ee83, 32'h437de1b5, 32'hc35faa5e},
  {32'hc373fb26, 32'h445c73b0, 32'h4382aae7},
  {32'h433fea60, 32'hc51c1ee4, 32'h423d30de},
  {32'hc4e2bb76, 32'hc36ba800, 32'hc388c941},
  {32'h4560ec12, 32'h44066b58, 32'h42c5afd6},
  {32'hc59b94b8, 32'hc2db5a5c, 32'h43ad9fb3},
  {32'h44eb9742, 32'h436db09b, 32'h442459f9},
  {32'h440a0542, 32'h45499ce2, 32'h4308aa5b},
  {32'h41ebf102, 32'hc4b7437b, 32'h42897160},
  {32'hc41d5a53, 32'h445540ab, 32'h4299bd60},
  {32'h43cbf8ec, 32'hc39d1703, 32'h44c1e7d3},
  {32'hc2a410e6, 32'h451313f6, 32'h42f1768a},
  {32'hc3a46687, 32'h4433aab0, 32'h450c4374},
  {32'hc436600b, 32'h449002a0, 32'h4454ae69},
  {32'h4484426f, 32'h4392c827, 32'h44be5782},
  {32'hc5141fa4, 32'h4323cbab, 32'h43e45dec},
  {32'h43ae9d50, 32'hc546c5f8, 32'hc336d13e},
  {32'hc56457e1, 32'h432e4539, 32'h41628adc},
  {32'h438f734d, 32'hc32e26ee, 32'hc18038ef},
  {32'hc515775a, 32'hc292bbf8, 32'hc49d5f92},
  {32'h43e62dc7, 32'hc43ea938, 32'h44d6c868},
  {32'hc4e439ca, 32'h416b4e70, 32'hc3d71ccc},
  {32'h43cb98f2, 32'h442913a6, 32'h45026a76},
  {32'hc4ac2a20, 32'hc42a34aa, 32'hc503787d},
  {32'h441b69b5, 32'h43c8fad2, 32'h44d67577},
  {32'hc480296e, 32'h43e09aec, 32'hc4286f60},
  {32'h43ec90a8, 32'hc4bd5523, 32'h44b8defe},
  {32'h4453955d, 32'hc40cf2f2, 32'hc39f1fc9},
  {32'h4397c1a0, 32'h4386428f, 32'hc41a6e9b},
  {32'h4336dc98, 32'hc356d4d6, 32'h44bb555b},
  {32'hc5069216, 32'h4467b0ae, 32'h43aa8fe6},
  {32'h450c1933, 32'h4318d99e, 32'h42dd5a5f},
  {32'hc44bf568, 32'h4402a0b3, 32'hc4e1bc11},
  {32'h43c0ef4a, 32'hc51f0bc4, 32'h43dbb9a0},
  {32'h43034a98, 32'hc4b47adb, 32'h44f39c85},
  {32'hc3150080, 32'h440ccec3, 32'hc362fd02},
  {32'hc37c7e1d, 32'hc353be4d, 32'h448d1d9a},
  {32'h44386c60, 32'hc373b2bb, 32'h448f857c},
  {32'hc529bd1c, 32'h43041d27, 32'hc4227112},
  {32'hc386de31, 32'hc3e71241, 32'h4547736a},
  {32'h43f1c8fc, 32'hc31fb0bb, 32'hc3f87e29},
  {32'hc208d39a, 32'hc3cbe37d, 32'h44a673b1},
  {32'h4365a26d, 32'h4527907e, 32'hc2b0a1be},
  {32'h44871a0d, 32'hc3bb3112, 32'hc280888e},
  {32'hc5943310, 32'hc369c25c, 32'h433a2bbb},
  {32'h450ec5d7, 32'h42271e99, 32'hc386403c},
  {32'hc1be737c, 32'h44bd1bfc, 32'hc2999367},
  {32'hc22e06e8, 32'hc5170a81, 32'hc39f12c0},
  {32'hc53188be, 32'h432d34bd, 32'h428408b9},
  {32'h448999a5, 32'hc4b825a5, 32'h42950de5},
  {32'hc54a39f7, 32'h44652c81, 32'h4429d740},
  {32'h4509f562, 32'hc4a260c6, 32'hc3972a7f},
  {32'h447887c0, 32'hc49a04c6, 32'h43ae91ff},
  {32'h43c5f8aa, 32'hc48db448, 32'hc444c900},
  {32'hc3cf21cf, 32'hc4cb6cd8, 32'h449bc956},
  {32'hc4699bee, 32'hc3da81a1, 32'h446ecf4f},
  {32'h45198227, 32'hc3677856, 32'hc392076e},
  {32'h420ec48c, 32'hc3363f40, 32'h44962aa3},
  {32'h437db630, 32'h43bf1cf1, 32'hc4e000af},
  {32'hc50d945c, 32'hc3b66f6e, 32'h43a70b74},
  {32'h449fb32f, 32'h44466efa, 32'hc3b604bb},
  {32'hc3fbc9ae, 32'h43a1616e, 32'hc38c1232},
  {32'hc327ecd0, 32'hc38d7fcf, 32'h44dacb60},
  {32'h43d7f530, 32'h414666de, 32'hc4d633b5},
  {32'h4411a254, 32'h448e5e3e, 32'hc3a7292e},
  {32'hc42a36d2, 32'hc38b82b3, 32'h4508fb35},
  {32'hc4945609, 32'h436b2a0c, 32'hc3d16c9e},
  {32'hc451ea90, 32'hc1aa1988, 32'h44a35a5c},
  {32'h43563d02, 32'h4501e075, 32'hc40066ad},
  {32'hc46e2d03, 32'hc2a9254f, 32'hc32bde1a},
  {32'h4549a062, 32'hc3896f32, 32'h429a20ea},
  {32'hc4b189cc, 32'h43fddec4, 32'hc26a38a0},
  {32'h452405f6, 32'h42b217f6, 32'hc33fd4fc},
  {32'h42f3ad9c, 32'hc51be9c2, 32'h43674e46},
  {32'hc1c31770, 32'h4552cd3d, 32'h43a520ca},
  {32'h443b7b1a, 32'hc4ffe362, 32'hc368ccc8},
  {32'hc3437d0c, 32'h44dd0472, 32'hc3c9bc38},
  {32'hc420b6f6, 32'h434e508a, 32'h42469e2e},
  {32'hc4ca356e, 32'hc22efe78, 32'h42d2dd72},
  {32'hc1ed2943, 32'h43119b46, 32'h447769b7},
  {32'h43a7e607, 32'hc4907439, 32'hc39c36c6},
  {32'hc37f3c7c, 32'hc3b9c866, 32'h450b2078},
  {32'hc3eac226, 32'h434b6324, 32'hc40419e9},
  {32'h440e4e77, 32'h43aea5b9, 32'h446ddfeb},
  {32'hc4edbdb8, 32'hc2c70518, 32'hc34d0d03},
  {32'h43b386ea, 32'h42d6138d, 32'h44ef28d3},
  {32'hc536bbdf, 32'hc3ff0396, 32'hc2a4dc67},
  {32'h451956fd, 32'h43280a5e, 32'h43e420e6},
  {32'hc41eee56, 32'hc3e9b6a2, 32'hc374f100},
  {32'h4400a02a, 32'hc50df2d1, 32'h45020553},
  {32'hc4472af0, 32'h43318523, 32'hc436a404},
  {32'h439c8dd8, 32'h43e9a52c, 32'h443acc10},
  {32'hc4a4cedb, 32'hc4298799, 32'hc3de3fab},
  {32'h421853ea, 32'h43bceb5b, 32'h44dbe410},
  {32'h43d33838, 32'hc32b518b, 32'hc4dd00a8},
  {32'hc2960770, 32'h449c578a, 32'h449a8f02},
  {32'hc42dcfd1, 32'hc48e06fa, 32'hc48f3055},
  {32'h442b85ef, 32'h41861620, 32'h426bc639},
  {32'hc5498409, 32'hc302f965, 32'h4232c8df},
  {32'h44961432, 32'h44f2481a, 32'hc2ebfee6},
  {32'hc4738b0b, 32'h431f7330, 32'h41c2d8da},
  {32'hc3e10da2, 32'h4532b638, 32'hc35eceac},
  {32'hc55767da, 32'h42dab642, 32'hc31f3814},
  {32'h4513bdb1, 32'h429bff82, 32'h4390068f},
  {32'hc5879707, 32'hc2886492, 32'hc3a1f25e},
  {32'h44522aba, 32'h439165b9, 32'h441f8861},
  {32'hc3491131, 32'h446c97f0, 32'hc50207d5},
  {32'h40c632a8, 32'hc3901ea4, 32'h44a89f77},
  {32'h430b654c, 32'hc2bf608a, 32'h433ce9a3},
  {32'hc3d27e02, 32'h454742b8, 32'hc134fb16},
  {32'h42e3fc40, 32'hc48d9a33, 32'hc4b6b691},
  {32'hc398f9f9, 32'h43dfd7cb, 32'h44ce976d},
  {32'hc3c99871, 32'hc40a1ea7, 32'hc53c74f2},
  {32'hc41714b2, 32'h43f24b9a, 32'h451f97d4},
  {32'h44e1f5bd, 32'hc2d5730c, 32'h42974b4f},
  {32'h43bff52a, 32'h43fae92d, 32'h441d01b8},
  {32'h42a02dc5, 32'hc2e5c0fe, 32'hc3ac6620},
  {32'hc319d899, 32'hc326cb17, 32'h4441c187},
  {32'h4523e72a, 32'h41d2be74, 32'hc409c013},
  {32'hc44aed1a, 32'hc1c43be5, 32'h45010e4d},
  {32'h451f466a, 32'hc38573a6, 32'hc3de8ab3},
  {32'hc48a998b, 32'h43c6a46b, 32'h44b41822},
  {32'hc2b69c6b, 32'h43025629, 32'hc56545be},
  {32'h433a6ca7, 32'hc31c1bcc, 32'h44a1b8da},
  {32'h44d474ba, 32'hc48470a6, 32'h42a571c3},
  {32'hc50de19d, 32'h4431cf62, 32'hc3e125a6},
  {32'h44d30f0f, 32'h4426ec33, 32'h4305e9c4},
  {32'hc50ae45f, 32'h44ba618e, 32'hc40502e0},
  {32'hc35ce630, 32'hc4190cf7, 32'h42c3a2c6},
  {32'h44b8469b, 32'hc3b891d4, 32'hc2c2bbf6},
  {32'h449b6bc4, 32'h4352993f, 32'h44161e5e},
  {32'hc4a7ca60, 32'h43ccea26, 32'hc43652d9},
  {32'h45874f49, 32'hc3423097, 32'hc2b66ca3},
  {32'h439bb2c2, 32'hc447c3d8, 32'h44857067},
  {32'hc2f77806, 32'hc15881ca, 32'hc56a5a82},
  {32'h44160513, 32'h433e2d85, 32'h44cab972},
  {32'hc4f37613, 32'hc3a6e817, 32'hc431d4f0},
  {32'h448d25cb, 32'hc4d79bcc, 32'h4339f00a},
  {32'hc321acc8, 32'h45268355, 32'h439ea75b},
  {32'hc4859f53, 32'hc3ecc0b3, 32'h430d5613},
  {32'hc31c361e, 32'h455fd206, 32'hc31402dc},
  {32'h4497ac60, 32'hc4dc0250, 32'hc322d8ca},
  {32'hc4352000, 32'hc387ed91, 32'hc4801fb8},
  {32'h43cb1333, 32'hc35925a5, 32'h452a82ea},
  {32'hc42b6a43, 32'hc1053b88, 32'hc4673b8e},
  {32'hc42f39e0, 32'hc3c5f233, 32'h421ba9ba},
  {32'hc4081194, 32'h447bc5f6, 32'h441d9164},
  {32'h440e80b7, 32'hc436661e, 32'hc4d24ac9},
  {32'hc537000c, 32'hc2aae0a5, 32'h40ddc79a},
  {32'h44271910, 32'h43190ca9, 32'hc4edb967},
  {32'hc4c6678a, 32'h4244ce89, 32'hc22facd4},
  {32'h44d6e3a3, 32'hc2910647, 32'h4218d65f},
  {32'hc587ebe0, 32'h418cc27f, 32'h436b0e1b},
  {32'h44b3c214, 32'h437201d0, 32'hc4a5f0a9},
  {32'h44b3ca8f, 32'h4217df90, 32'h4316ca13},
  {32'h4471fcc4, 32'hc3820a4c, 32'hc426d851},
  {32'hc4da235f, 32'h435882ec, 32'h4495507a},
  {32'hc3f74b7a, 32'hc3996c54, 32'hc38d5cbe},
  {32'hc42434f1, 32'h447c0293, 32'h43a35d5f},
  {32'h442c8a40, 32'hc1889025, 32'hc50088fb},
  {32'h44e945c7, 32'hc3e74c27, 32'hc47be42e},
  {32'hc389987a, 32'hc37f0b54, 32'h451b6b33},
  {32'h44f93eab, 32'hc1753c88, 32'h42c1f661},
  {32'hc2707aa8, 32'hc4305fd9, 32'hbf1fe360},
  {32'h43ee1876, 32'h44caae35, 32'h4253797e},
  {32'hc287ac28, 32'hc4b845ce, 32'h432dda67},
  {32'h4558a1fd, 32'h438e4ad7, 32'h43286188},
  {32'hc4b6b7d2, 32'hc4013f7e, 32'h43e64660},
  {32'h43adc550, 32'hc3476a12, 32'h4384f9be},
  {32'hc49c41bc, 32'h434d4a48, 32'hc416634a},
  {32'h44b04bdc, 32'hc3080f23, 32'h43cc8a4c},
  {32'hc4b0e370, 32'h42f1cdb0, 32'h440ce968},
  {32'h44c639ef, 32'h4381d82d, 32'h44affd21},
  {32'hc4b5123c, 32'hc4aa5977, 32'hc412856a},
  {32'hc401afb8, 32'h43b0a8e1, 32'h4489e59e},
  {32'hc4710510, 32'hc48099de, 32'hc3514e4d},
  {32'h4360f03d, 32'h442acdf2, 32'h44ee80a7},
  {32'h444c268b, 32'hc3f40d64, 32'hc456b7ee},
  {32'h44cb0860, 32'hc425212c, 32'h441ef2e2},
  {32'hc4ccb52f, 32'h4439d1c8, 32'hc499e4a9},
  {32'h43a7bf0a, 32'hc07492a0, 32'hc33cda58},
  {32'hc48c5425, 32'hc50a7918, 32'hc3ae9940},
  {32'h44474994, 32'h44d18ef6, 32'h4390b9c6},
  {32'h44304026, 32'hc455ef98, 32'h43962fdb},
  {32'hc32528d4, 32'h4535c68e, 32'hc1d5e743},
  {32'hc2647f78, 32'hc4aa37b0, 32'hc4888431},
  {32'hc455fdf7, 32'hc2d71fca, 32'hc2fc6d1e},
  {32'hc322ab90, 32'hc2f09bd3, 32'hc34a884b},
  {32'hc0ae3f50, 32'hc5556910, 32'hc2b51579},
  {32'h44fb2e01, 32'h44528920, 32'h432a1e9c},
  {32'hc4c120b5, 32'h44344ecb, 32'hc35ffa21},
  {32'h45187a45, 32'h418c36b4, 32'hc31cb632},
  {32'hc3f67904, 32'hc3b37616, 32'hc2b4df56},
  {32'hc369798a, 32'hc2c0e691, 32'h438241bf},
  {32'hc4b1cbae, 32'hc3a406eb, 32'hc407bcfc},
  {32'hc22ccd80, 32'hc3424695, 32'hc2d3b511},
  {32'hc39cb684, 32'hc4679916, 32'h43d6717c},
  {32'h4351bf16, 32'h44e4e7be, 32'h424ed201},
  {32'hc4e187a5, 32'hc3c0494e, 32'hc385167f},
  {32'hc48131fb, 32'h43430e88, 32'hc3997b82},
  {32'hc4f72cae, 32'hc2ef843e, 32'h4384d0a2},
  {32'h45016476, 32'h440a80e2, 32'h43675b68},
  {32'h44c4d7d5, 32'hc16af372, 32'hc2086c96},
  {32'h44bed339, 32'h43a53bbb, 32'hc445e10f},
  {32'hc3f9e246, 32'h43d020d2, 32'h45309ff6},
  {32'h454bc26b, 32'hc3abe4ce, 32'hc40f6dbb},
  {32'hc444e3a8, 32'hc48090a3, 32'h44442193},
  {32'h44337596, 32'h44d8b3cf, 32'h41cdeaee},
  {32'hc2866cd8, 32'hc4bf0f1b, 32'hc3b94741},
  {32'h4316ba14, 32'h44cb3c1e, 32'hc35af815},
  {32'hc45cfd41, 32'h435fcabc, 32'h44d26d95},
  {32'hc3cf6cbe, 32'hc2cff816, 32'hc487ecfe},
  {32'hc5578125, 32'hc2affab5, 32'h4410e291},
  {32'h44833993, 32'hc302f7b5, 32'hc514cbc6},
  {32'h44c07317, 32'hc4650661, 32'hc415edc9},
  {32'hc3e3f378, 32'h445a2083, 32'h448f513e},
  {32'h44a5bf4d, 32'hc3bdea2a, 32'h434f1386},
  {32'hc313a3f2, 32'h4553b1bb, 32'h42e2676e},
  {32'h444db10c, 32'hc51b4e38, 32'h440135ae},
  {32'hc46ab05a, 32'hc3560a3f, 32'hc3712cbd},
  {32'hc3dbb52c, 32'hc41c55a0, 32'hc40630e5},
  {32'hc547063a, 32'h4433e08c, 32'h439666a2},
  {32'hc39afee0, 32'hc37c3592, 32'hc2b075bf},
  {32'h43de292c, 32'h4540bf55, 32'h43673c6d},
  {32'h44490582, 32'hc4c0433d, 32'h449c0dac},
  {32'h429e00cd, 32'h445a6e61, 32'h437b2a97},
  {32'hc34da159, 32'hc490387f, 32'hc35ff5ac},
  {32'hc2804980, 32'h45164dcd, 32'h4345ee1c},
  {32'h441e925c, 32'hc3b03d5b, 32'h4423f936},
  {32'hc2dcb814, 32'hc3dfacd0, 32'hc52cf8fd},
  {32'h426d5cd0, 32'h43ffb15b, 32'h451202ab},
  {32'hc4361cee, 32'h444be084, 32'h4418fe84},
  {32'h44369be8, 32'hc47c0af1, 32'h41f7d16e},
  {32'hc4a457ab, 32'h448e7746, 32'h43267d15},
  {32'hc1d01bf4, 32'hc4b8a5d7, 32'h43c597f6},
  {32'hc4c4ca56, 32'h44d2b107, 32'hc2a1ba68},
  {32'h4533a7de, 32'hc3bdcad1, 32'hc27e43b4},
  {32'h445ab475, 32'hc3856501, 32'hc46c1bc0},
  {32'h44b6ab20, 32'h43e39b81, 32'h44be5d85},
  {32'hc5761db9, 32'hc3347c26, 32'hc28a2b7a},
  {32'h4489687e, 32'hc3c0cc6b, 32'h44651784},
  {32'hc32a6518, 32'h425b375c, 32'hc46544ec},
  {32'hc4d93bd1, 32'hc42066e5, 32'h44a85753},
  {32'h44912aff, 32'hc438680f, 32'hc2fdb667},
  {32'h430091e5, 32'hc2d7bd59, 32'hc505b12c},
  {32'h44d89734, 32'hc40562d4, 32'h43e805b8},
  {32'h438a0c30, 32'h449d1eac, 32'h41c3639e},
  {32'hc49b398e, 32'hc3027c66, 32'h445cca06},
  {32'hc492ae92, 32'h43b112ce, 32'hc3a2534d},
  {32'h44d214f5, 32'hc3a8324f, 32'h443568b9},
  {32'h4424aadd, 32'h4327f603, 32'h44af4c9e},
  {32'hc2d38724, 32'hc4ce043c, 32'hc502c70c},
  {32'h45123b74, 32'hc35dafe6, 32'hc487d6f2},
  {32'h4333da82, 32'hc3d5b8cf, 32'h43f3298a},
  {32'hc3d53c55, 32'h450ea88c, 32'hc42ba429},
  {32'h44178395, 32'hc355c295, 32'h44a709f8},
  {32'h44351291, 32'h44412280, 32'hc3294992},
  {32'h451f1ae1, 32'hc31ff70a, 32'h4319c536},
  {32'hc1d9bb00, 32'h45325d1d, 32'hc3cc659e},
  {32'hc47ee4fa, 32'h42d22a6f, 32'h43ab4a4d},
  {32'hc494bb40, 32'hc3e01959, 32'hc478e674},
  {32'hc384d4c8, 32'hc2e69cca, 32'h4486327c},
  {32'h44725902, 32'h416e5f3d, 32'h42fd8f52},
  {32'h44c6b433, 32'hc3c096f0, 32'hc2a6581a},
  {32'hc41546fc, 32'h4473c8a8, 32'hc43aa944},
  {32'h42c312ae, 32'hc446ce90, 32'h4338b29e},
  {32'hc3c449d3, 32'h44f99564, 32'h43ad8224},
  {32'h43a609cb, 32'hc533bae0, 32'hc25c948e},
  {32'h44c281f2, 32'h435222d4, 32'h4361c669},
  {32'h44df9298, 32'h445c6298, 32'hc40f2862},
  {32'hc2fbc31d, 32'hc44d61ae, 32'h44b28ba4},
  {32'h43d8ac0a, 32'hc2e340ec, 32'h4509af6e},
  {32'h43199f0e, 32'hc21771af, 32'hc515b0b4},
  {32'hc3b7f773, 32'h43a03b58, 32'h4498c1b2},
  {32'h41a3944e, 32'h44a1a51f, 32'hc3ceb4e8},
  {32'hc522cf71, 32'hc2094094, 32'h42feca94},
  {32'h44e482c2, 32'h43dbc0c6, 32'h42fbd793},
  {32'h444a94b6, 32'hc3f5b519, 32'hc36b1b9a},
  {32'h424d77f0, 32'h4470ea14, 32'h4489e167},
  {32'h43870802, 32'hc4ea3ce1, 32'hc4b3ebc6},
  {32'h43784b14, 32'hc2cf6d41, 32'hc4d0165a},
  {32'hc4881784, 32'hc4a4dd94, 32'hc3854fa0},
  {32'h439da49c, 32'hc34eee3e, 32'h43477b32},
  {32'hc4457f91, 32'h43033611, 32'h438dea3b},
  {32'h4386f488, 32'h4432e46a, 32'hc4df172e},
  {32'hc3087889, 32'hc3832f2c, 32'h448792ef},
  {32'h4535fd28, 32'hc2b5ad9a, 32'hc36a81eb},
  {32'hc3fc8844, 32'h43f4fac4, 32'h43e51c59},
  {32'h42c23cc0, 32'h41e1cee3, 32'h42b4c234},
  {32'hc543ea02, 32'hc3b629da, 32'h431576f8},
  {32'h45243a8f, 32'h43e17b08, 32'hc41154d2},
  {32'hc44eb1be, 32'hc32a18f1, 32'h434ae27f},
  {32'h44947050, 32'h44770a2e, 32'hc2450023},
  {32'hc5280d7a, 32'hc3ca9f02, 32'hc38d2020},
  {32'h455aa0d1, 32'hc3b51227, 32'hc13eaf4d},
  {32'h44210287, 32'hc3525812, 32'h43c73059},
  {32'h41e08133, 32'hc4a5ce3f, 32'hc391c4be},
  {32'h44714ff3, 32'hc3cf7dc2, 32'h445f54c3},
  {32'h45044b2a, 32'hc3c54c3e, 32'h42b37a6e},
  {32'h4450d81f, 32'hc3783fe5, 32'h45230093},
  {32'hc4ad58e7, 32'hc433c4fd, 32'hc3cd95b3},
  {32'h43714fbb, 32'hc3197df1, 32'h44e0a04a},
  {32'hc38015b8, 32'hc4bd2800, 32'hc4d73ab5},
  {32'h41541620, 32'h45013ac9, 32'h44bb1d7e},
  {32'h44257ade, 32'hc37350dc, 32'hc3b4c26f},
  {32'hc42b7680, 32'hc3624168, 32'h42c2a723},
  {32'h3ff76380, 32'h44c3248d, 32'hc4bdb156},
  {32'h447033a2, 32'h442c65e7, 32'h43a8934f},
  {32'hc426ba6b, 32'hc4fdc7ad, 32'hc2f15d8f},
  {32'h436a1bc0, 32'h43e24b6d, 32'h4520f02c},
  {32'hc493870e, 32'h4365d658, 32'hc354e7af},
  {32'hc3a0a988, 32'h44a25002, 32'h4534223d},
  {32'hc4518fbb, 32'hc47bc045, 32'hc387642d},
  {32'hc3600d23, 32'h446bb131, 32'h43e6b202},
  {32'hc4d5774e, 32'hc48db8f7, 32'hc38f33d0},
  {32'h454b7356, 32'h448e3418, 32'h4414c065},
  {32'h44d16731, 32'hc4044dbd, 32'hc38fd813},
  {32'hc35abab6, 32'h4573b45f, 32'h434c21dc},
  {32'hc4c8d82a, 32'hc4b8c498, 32'h4138457e},
  {32'h43d4ae36, 32'hc36a06f8, 32'h432cd95a},
  {32'hc55853e7, 32'h43fca34c, 32'hc261d6c6},
  {32'h4491f4c4, 32'h4393e278, 32'h4443e66d},
  {32'h440eeaa2, 32'hc4c49891, 32'hc44b78a2},
  {32'hc258d5f8, 32'hc49cae97, 32'h44c20ced},
  {32'hc2c66e60, 32'h42457d37, 32'hc3f5cbac},
  {32'hc404aa1a, 32'h43a092e9, 32'h44c465e4},
  {32'hc27c58f0, 32'hc2008cfd, 32'hc519324b},
  {32'h44dfec57, 32'hc33651c6, 32'h42fa0ba4},
  {32'h4545a487, 32'hc441c485, 32'hc427b466},
  {32'h42af425a, 32'h448f4f72, 32'h4506b6a7},
  {32'hc3fcd242, 32'hc43c4605, 32'hc4a1b9e0},
  {32'h422ed46c, 32'hc27277be, 32'h44e233b8},
  {32'hc3655928, 32'hc1a27252, 32'hc4a5e07a},
  {32'h443fea1b, 32'h4329bb8a, 32'h439a6f14},
  {32'h44d9939b, 32'h4295c3f4, 32'hc44f8066},
  {32'hc3bf2a88, 32'h45154bd0, 32'h41c6f043},
  {32'h450060f7, 32'h43bd2eaa, 32'h42ad60fc},
  {32'hc537c6bb, 32'hc2429c63, 32'h43af13a2},
  {32'h421c6aa6, 32'hc293df32, 32'hc527e1b7},
  {32'h4451edd8, 32'h428ab96a, 32'h43fe9277},
  {32'h43cfc09c, 32'hc46780be, 32'hc3ccb3fa},
  {32'hc580edaa, 32'h438f34f0, 32'h435ba244},
  {32'h452dc2ce, 32'h42b74d74, 32'hc3e0ec5f},
  {32'h442f5ec1, 32'h447e61aa, 32'h43c3f5f6},
  {32'h453746a5, 32'hc3aaf040, 32'h43966b03},
  {32'h439d35bf, 32'h43906d6f, 32'h4399ff57},
  {32'h44ba2d3f, 32'h42a9e1c1, 32'h431273dd},
  {32'hc40f8e0c, 32'hc456d33e, 32'h441b9aa7},
  {32'h4544a148, 32'hc31141fc, 32'h43a36756},
  {32'h44f36e72, 32'h40d9020f, 32'hc383c46d},
  {32'hc57c9b82, 32'h41ce4fbd, 32'h4435ac5d},
  {32'h44ad2419, 32'h43fc3949, 32'h44446791},
  {32'h43808f2b, 32'h449c904b, 32'hc3b19301},
  {32'h44ab1e0a, 32'hc4beeada, 32'h42668cae},
  {32'hc54ddc2a, 32'hc2b1ae2d, 32'hc30ef489},
  {32'hc3966973, 32'hc403b11e, 32'h43a5c86e},
  {32'hc49a77fa, 32'h44508274, 32'hc3183afc},
  {32'h4438215e, 32'hc500345d, 32'h43a7f9c0},
  {32'hc3da4477, 32'hc395bc71, 32'hc4b36a9d},
  {32'h44bf8301, 32'hc13b6716, 32'h43d48f57},
  {32'hc3b6a7b8, 32'h44245697, 32'hc515206e},
  {32'h42f8e1bd, 32'hc2c9f3e7, 32'hc39fb2b2},
  {32'h43c4a5a1, 32'h440e92b9, 32'h44fbb586},
  {32'hc36624be, 32'hc4ac9b46, 32'hc41d74e9},
  {32'hc2ba8b10, 32'h44d5ecd2, 32'hc3886ac9},
  {32'hc2c91b2e, 32'hc3abec97, 32'hc4c407fa},
  {32'h422f03e8, 32'h43a9ace4, 32'h4552cefc},
  {32'h446f20e3, 32'hc433e411, 32'hc37b4d9e},
  {32'hc41d6d08, 32'hc48b3c62, 32'h444a9cc5},
  {32'h4463b034, 32'h444dca76, 32'hc4138224},
  {32'h4399d40e, 32'h4409cb4b, 32'h44824ddf},
  {32'h454c6a38, 32'hc3cb3824, 32'hc2dbde06},
  {32'hc48d3df5, 32'h434b185c, 32'h44c335c5},
  {32'h44d1ac65, 32'hc06ddde8, 32'hc4326b96},
  {32'h43ae0608, 32'h44b5aa2a, 32'h44a1a6dc},
  {32'h45310930, 32'hc417e1ab, 32'hc350d733},
  {32'h454d1bc8, 32'hc1c445c8, 32'hc3ec972d},
  {32'hc3fd0b08, 32'hc3be8ac9, 32'h453acb13},
  {32'h43bed1b0, 32'h4341ea83, 32'h42ea7fae},
  {32'hc37da6f9, 32'hc523f5b4, 32'hc22c4a1b},
  {32'h45287a49, 32'hc3f62476, 32'h43f6082a},
  {32'h4494eaf6, 32'hc45614f5, 32'hc2979bdb},
  {32'h449c9a96, 32'h4502fdd6, 32'h43337fb2},
  {32'hc502b8cc, 32'hc3eaa060, 32'hc44f0d4a},
  {32'h44884661, 32'h412a1500, 32'h4369ed28},
  {32'hc3236100, 32'hc296c598, 32'h448ecfe7},
  {32'h4521a0ce, 32'h44039e5e, 32'hc37621d6},
  {32'h4307ca30, 32'hc3974309, 32'hc276ea4e},
  {32'h430d9a00, 32'hc2e8dcc6, 32'h454d7d5a},
  {32'hc49d0c0f, 32'hc46b47f5, 32'hc4ba41a3},
  {32'h44917fa7, 32'h43fa9859, 32'h42dc5776},
  {32'hc345547e, 32'hc531413a, 32'hc3235937},
  {32'h44f056fc, 32'h420618a9, 32'h41801864},
  {32'h43f6898e, 32'hc3a83456, 32'hc48ae636},
  {32'h44a32e50, 32'hc3f1c4c5, 32'h44b854af},
  {32'hc46fc79b, 32'hc48f4cb8, 32'hc462756d},
  {32'h45109d4e, 32'hc3419ad5, 32'h41b6bf94},
  {32'hc2fa1600, 32'hc4c10406, 32'hc44c9e4f},
  {32'hc33c5d81, 32'h42693345, 32'h452fe979},
  {32'hc496f6f4, 32'hc3b9d335, 32'h43217996},
  {32'h44270bd8, 32'h449a4dd7, 32'h44a0152b},
  {32'hc51a62ab, 32'hc3a46bc9, 32'hc2c0b510},
  {32'h453af668, 32'hc3a990b4, 32'hc41ab566},
  {32'h436712d0, 32'h42166dd5, 32'h44061759},
  {32'hc4ca1c64, 32'hc4278031, 32'hc32cce78},
  {32'h44c4016a, 32'h43d89634, 32'h440bc125},
  {32'hc4ba819a, 32'h4398fe6a, 32'h441f7f85},
  {32'h43495274, 32'h458126ce, 32'hc25adf20},
  {32'h42fdae65, 32'hc4ba5c06, 32'hc34eb041},
  {32'h4462c70f, 32'h4442f5e4, 32'h43ab81bd},
  {32'hc5463d3a, 32'hc3a6bc7b, 32'h40dd01df},
  {32'h456a1db3, 32'h44254121, 32'h4439a0b6},
  {32'hc4c582fa, 32'h42ed35b3, 32'h42da38f8},
  {32'h43c42a08, 32'h4516c20a, 32'h4370989b},
  {32'hc3c7c0bf, 32'hc455d012, 32'h4483be6a},
  {32'hc4f144ad, 32'h43a21e51, 32'hc1a293c1},
  {32'h438873c0, 32'hc2d83c5a, 32'h451ee668},
  {32'h44d26b20, 32'h434085a8, 32'h429b1467},
  {32'h44393f88, 32'hc2873d20, 32'h42bb3add},
  {32'h43a882e0, 32'h44475c41, 32'hc2ef86e1},
  {32'hc39e57fa, 32'hc3547842, 32'h445a931d},
  {32'h4473248b, 32'h43043e94, 32'h429f2fc1},
  {32'hc49a27c5, 32'hc3943f72, 32'hc3f1cd74},
  {32'h44a05268, 32'h44d3f463, 32'hc449ee37},
  {32'h42af885e, 32'h437464f8, 32'h438fcf8c},
  {32'h431940b0, 32'hbedcac40, 32'hc44228a9},
  {32'h436d9ebe, 32'hc4945341, 32'h449eedcd},
  {32'h456ca860, 32'h44329ac4, 32'hc31dcbd2},
  {32'hc5372bc8, 32'h43aa9b1b, 32'h44743d71},
  {32'h455eeba6, 32'hc41d4c9c, 32'hc46bb64c},
  {32'h44306639, 32'hc4c56a6c, 32'h42f434bc},
  {32'hc477de92, 32'h4505939e, 32'h43ac12af},
  {32'hc42f1652, 32'hc433995a, 32'h42acffb1},
  {32'hc4a8a43e, 32'h43bb41eb, 32'h4445f9a2},
  {32'h44677428, 32'hc3e346b4, 32'h43b8c830},
  {32'hc4da17b9, 32'hc32c5142, 32'hc138aa02},
  {32'h456275b7, 32'h42b9b6dd, 32'hc32a785e},
  {32'hc42d11c4, 32'h43451a36, 32'h43d16e35},
  {32'h4516b3a3, 32'hc312db75, 32'h433113ed},
  {32'hc4906916, 32'h44033c0b, 32'hc4cf5d0d},
  {32'h44a15bf7, 32'h41c26f2a, 32'h436c634b},
  {32'hc4d85c42, 32'h427e6891, 32'hc2fb9563},
  {32'h441365c6, 32'hc2c72ace, 32'h444014f8},
  {32'hc3c417db, 32'h429db895, 32'hc3857302},
  {32'h432ca13e, 32'hc3b41cf5, 32'hc285298d},
  {32'hc4830351, 32'hc4327832, 32'hc4880313},
  {32'h4315ab25, 32'hc387674f, 32'h43d4d8ac},
  {32'hc4eacb5c, 32'hc2ed6e2a, 32'hc3375d78},
  {32'h449b193a, 32'hc4016d83, 32'h44e1ad69},
  {32'hc566f955, 32'h430f9a0c, 32'h4207adba},
  {32'h440d235a, 32'hc38cec35, 32'hc2afb08a},
  {32'hc3c2aba2, 32'h4521f188, 32'h4350cce9},
  {32'h436898e0, 32'hc51d0a34, 32'h43f51213},
  {32'h44c4e130, 32'h44549aef, 32'hc397f05e},
  {32'hc2830b0c, 32'h439b7688, 32'h45678400},
  {32'hc4fd4455, 32'hc3cb02e9, 32'hc4dba7e4},
  {32'hc4f1680c, 32'hc384bfd1, 32'hc32c7673},
  {32'hc43e1f64, 32'h448e5b89, 32'hc42415c7},
  {32'hc2f82e22, 32'h43b85898, 32'h45407d6a},
  {32'hc2dffd2c, 32'h419b844f, 32'hc3c7d62e},
  {32'hc48a84aa, 32'hc137d191, 32'hc44614d0},
  {32'h44a266a7, 32'hc4dea302, 32'hc3ecc08f},
  {32'hc380719c, 32'h45080d4f, 32'h4309bf45},
  {32'h44584296, 32'h43a31bea, 32'h448386f4},
  {32'hc488a9e5, 32'h443884de, 32'hc48a6374},
  {32'h4409bd0c, 32'hc2e589d2, 32'h45110368},
  {32'h44772418, 32'hc4115044, 32'h44b0e950},
  {32'h43cfdaf2, 32'h448ce562, 32'hc5233d70},
  {32'hc397083a, 32'h44a3c1f4, 32'h433d37b0},
  {32'hc1ad39bb, 32'h41dacce6, 32'h439a5c2f},
  {32'hc41c2dd6, 32'h440b5221, 32'h439b7f01},
  {32'h4477fc5c, 32'hc3ab8f52, 32'h44295cfe},
  {32'h44d659e5, 32'hc3192f03, 32'h4318e40b},
  {32'h42f8816d, 32'hc4317c9a, 32'hc2d3b2ee},
  {32'hc34bb4c8, 32'h44b5089c, 32'hc31fb644},
  {32'h44c4ea18, 32'h42adbdc1, 32'h443905b0},
  {32'hc5833ef5, 32'hc36b1061, 32'hc3c0324d},
  {32'h450deda1, 32'hc2d2fb28, 32'h43cefda0},
  {32'hc414d064, 32'h4034ccf8, 32'hc3b09636},
  {32'hc238a4a0, 32'hc55d632a, 32'hc3849cda},
  {32'hc3441ba8, 32'h456520b6, 32'hc19dd46a},
  {32'h43a4d6ae, 32'h3fd6dc65, 32'h41c14cba},
  {32'hc528515e, 32'h4450bfac, 32'hc40c6a2d},
  {32'h43875520, 32'hc4eb0c11, 32'hc1c56246},
  {32'hc48db67c, 32'hc35c265d, 32'h4392f9f2},
  {32'hc4692c42, 32'h4375cd04, 32'hc51e1f15},
  {32'hc26d1e52, 32'h441d4e6f, 32'h4498a17e},
  {32'hc38565f4, 32'hc426bbc1, 32'h44899dff},
  {32'hc30350c0, 32'h44b44eab, 32'hc42d69e9},
  {32'hc3b89d85, 32'hc50566a8, 32'hc3053099},
  {32'hc33fc550, 32'h44141e99, 32'hc542e316},
  {32'hc3ddc782, 32'hc398770f, 32'h44238a8a},
  {32'h4511c3c2, 32'hc355436e, 32'h4404399e},
  {32'h44bebd7f, 32'hc338d1d3, 32'h44159e55},
  {32'hc3fb5035, 32'h450d416f, 32'h44c90954},
  {32'h44ac0bbc, 32'hc308e353, 32'hc48f90cb},
  {32'h435ce2f0, 32'h4486bdbe, 32'h41b20186},
  {32'hc4c4a526, 32'hc20dc611, 32'h4324f0a5},
  {32'h43f129ca, 32'h4507d5aa, 32'hc3867277},
  {32'hc4efcc31, 32'hc3c9eb80, 32'h43728783},
  {32'h4412222b, 32'h4441664b, 32'hc48479e4},
  {32'h4415a199, 32'hc385bdc9, 32'h44146409},
  {32'h450696a9, 32'hc3fef3a5, 32'hc381e7ea},
  {32'hc4d6f698, 32'h43ef77de, 32'hc3263096},
  {32'h44d2bc3a, 32'h441990ba, 32'hc34d8b38},
  {32'hc3dff086, 32'hc3d472b0, 32'hc415678e},
  {32'h43b2cf82, 32'h4524d2eb, 32'h43eaf695},
  {32'hc4e17bbf, 32'h41f4de70, 32'h42ccd5d6},
  {32'h453767c3, 32'h4453723a, 32'h40d48fde},
  {32'hc52b17d7, 32'hc40d3961, 32'h4224c4ca},
  {32'h432aad6c, 32'h4431481e, 32'hc14ea3cc},
  {32'hc3795e68, 32'h42c5df3c, 32'h4359ecad},
  {32'h445dddf9, 32'h436bc0c4, 32'hc4a9a79b},
  {32'h44d75233, 32'h42b62c74, 32'h4447bb10},
  {32'hc3b8679d, 32'hc461d2ad, 32'hc42527aa},
  {32'h42f17ce0, 32'h44f50c3e, 32'h44479953},
  {32'hc23c7100, 32'hc48122d1, 32'hc4ad18bf},
  {32'hc472dad4, 32'h4218e070, 32'h43bc2a9c},
  {32'hc432ee34, 32'hc413ffe0, 32'hc47ab954},
  {32'h4424d7d6, 32'h44800835, 32'h44a310df},
  {32'h43999500, 32'hc2baa0f0, 32'hc4c997b3},
  {32'h44059a7d, 32'hc2f00065, 32'h415585d3},
  {32'hc1a29468, 32'hc2c2b319, 32'hc4b9335c},
  {32'hc4c74682, 32'hc2bde67b, 32'h43e51144},
  {32'h4312c3de, 32'hc527d1cc, 32'hc3adb71a},
  {32'h44533cf2, 32'h44d61700, 32'hc3185c9e},
  {32'h4292cf68, 32'hc2f83dc0, 32'h4248227b},
  {32'h43766f5c, 32'h44b64a0d, 32'h44ae71d4},
  {32'hc484e012, 32'hc41d5a5b, 32'hc4988bae},
  {32'h455b7bdf, 32'hc3bd453c, 32'hc38a36d5},
  {32'hc502cef0, 32'hc479bc21, 32'h42c86fcb},
  {32'h44d939b7, 32'h449f8e26, 32'h4337c010},
  {32'h4498b78e, 32'hc4467df3, 32'hc2ea7c46},
  {32'h44d2b138, 32'h43c0eeb0, 32'hc2dae32e},
  {32'hc50c0e15, 32'hc3de6208, 32'h43d24a16},
  {32'hc219da48, 32'h440ee99a, 32'hc2d45111},
  {32'hc4cf4b06, 32'h43ea25f4, 32'hc4999138},
  {32'h4475e861, 32'h427b1cd3, 32'h43b9c4e3},
  {32'hc39ef421, 32'h44add6cb, 32'hc41b631f},
  {32'h42c994ee, 32'hc50aedba, 32'h44adb309},
  {32'hc2873918, 32'hc3cb9fde, 32'hc3bcd230},
  {32'hc4510e69, 32'h442f36ad, 32'h443256f8},
  {32'hc3e6062b, 32'hc1c3c75d, 32'hc548a2d1},
  {32'hc44bc2a6, 32'h4388920e, 32'h44932a44},
  {32'h44966028, 32'hc485bbe6, 32'hc46b3ccc},
  {32'hc561c595, 32'hc29b5c6d, 32'h435ba3fe},
  {32'h4390aeb5, 32'hc47ec268, 32'hc48de04a},
  {32'h43d359bf, 32'h454629a1, 32'h4409bf6e},
  {32'hc2c6aff0, 32'hc4a08f67, 32'hc46e2a2a},
  {32'hc3a56340, 32'hc498e417, 32'h4435ab44},
  {32'h4418bad0, 32'hc2f0cd4b, 32'hc4943198},
  {32'hc3e00624, 32'hc343518f, 32'h43a6d593},
  {32'hc2c82e10, 32'hc3d88c5e, 32'hc41225d5},
  {32'hc3146aa8, 32'h43bcfb90, 32'h45241502},
  {32'h44d46e96, 32'h43252dbe, 32'hc3c8663e},
  {32'hc4b58c32, 32'hc3cbe362, 32'h438fea57},
  {32'h456e470e, 32'hc44313bc, 32'hc1c08970},
  {32'hc45a5be3, 32'h450a8b2e, 32'h43c5f8c5},
  {32'h445cfcff, 32'hc3255be7, 32'hc31ac73a},
  {32'hc524e691, 32'h43c04319, 32'hc3391aa3},
  {32'h452b7814, 32'hc3e20fea, 32'hc3100c17},
  {32'hc4ba578a, 32'h43da8235, 32'h42e4d683},
  {32'h45236bc3, 32'h439b71aa, 32'hc281063b},
  {32'hc4cd77a4, 32'h440bf809, 32'hc40f82a2},
  {32'hc3171b7a, 32'hc3e2b552, 32'hc3490483},
  {32'h424e396c, 32'hc40c0862, 32'h447cf573},
  {32'hc49e6e9b, 32'hc1d130aa, 32'hc5106043},
  {32'h44aff532, 32'hc42fc8c6, 32'h44ab4278},
  {32'hc3b3923d, 32'h446b0441, 32'hc37df0a4},
  {32'h42952ed4, 32'hc5374659, 32'hc31c80e0},
  {32'hc36f6c3b, 32'h455b03db, 32'hc1963963},
  {32'hc501c0d9, 32'hc270281e, 32'h438e05d7},
  {32'hc407fc00, 32'h442fb927, 32'hc33da998},
  {32'h428d5333, 32'hc5006aa4, 32'h43e594cc},
  {32'hc4e41578, 32'hc3c32007, 32'hc1c124e7},
  {32'h45062712, 32'h41bb0bbd, 32'hc2f0a123},
  {32'hc38e553e, 32'hc38f4256, 32'hc51d8ec8},
  {32'hc45f31b9, 32'h43b2827e, 32'h42eb9259},
  {32'hc529aba0, 32'hc3ba9de6, 32'hc24945cc},
  {32'h43c7063c, 32'hc320a267, 32'hc50a5d59},
  {32'hc487485b, 32'h4212648b, 32'h437901b1},
  {32'h451158d8, 32'h43974831, 32'h428ce782},
  {32'hc462475c, 32'h440c8a9e, 32'h43f9cbf0},
  {32'h4550b9fc, 32'hc37d5bd7, 32'hc2f50627},
  {32'hc4a568a4, 32'h438fd50e, 32'h44a35362},
  {32'h430c7120, 32'hc38c6fe8, 32'hc4d66016},
  {32'hc4c4149c, 32'h43e2abbc, 32'hc3d69098},
  {32'h4520aacb, 32'hc3fe860e, 32'hc4853918},
  {32'hc30313f6, 32'h452a0ef3, 32'h449c5ff7},
  {32'h42db5fbc, 32'hc3ea4c91, 32'hc410ce76},
  {32'hc54fd02e, 32'h441bac30, 32'h4396fe6d},
  {32'h44d31cbb, 32'hc4221335, 32'hc4db4b49},
  {32'h43e9e168, 32'h43a95fb2, 32'hc439da60},
  {32'hc459fa69, 32'h435b4f9a, 32'h44967ec8},
  {32'h44b32e0a, 32'h4401ed71, 32'hc10a36b1},
  {32'hc3e6f2a7, 32'hc514972c, 32'hc36b032e},
  {32'h441762c8, 32'h44e460a4, 32'hc1e0fa90},
  {32'h446b0ed4, 32'hc4d83ddc, 32'hc3cd3714},
  {32'h44ca3b0c, 32'h44a6fb04, 32'h43b5fa10},
  {32'hc4885d32, 32'hc3b59ada, 32'hc36f640f},
  {32'hc4f1232a, 32'h42538494, 32'h440d1d33},
  {32'hc4c4c5fc, 32'hc293ed8b, 32'hc42e80e2},
  {32'h45193784, 32'h43092cc1, 32'h419ab2e4},
  {32'h43ca8924, 32'hc47d2c3d, 32'hc41ffea5},
  {32'h42a48b80, 32'h45248846, 32'h4358da16},
  {32'hc4908b63, 32'hc3c8dd92, 32'hc400c637},
  {32'hc4758b59, 32'h42644152, 32'h446725ec},
  {32'hc4289677, 32'hc331035c, 32'hc4a75aad},
  {32'h42ed44a5, 32'h43b4109e, 32'h4557897c},
  {32'hc3e2e028, 32'h40f7ac9c, 32'hc463aa38},
  {32'h4555d6bb, 32'h42ed9115, 32'h43214fe0},
  {32'hc4f3adca, 32'h4393d102, 32'hc381c998},
  {32'h453bb3ac, 32'h43f9a762, 32'h43029ffe},
  {32'hc3e16344, 32'hc4a3315b, 32'hc45a5667},
  {32'hc4498306, 32'h451de6e2, 32'hc38ffa76},
  {32'hc4acf301, 32'hc2d9a99d, 32'h42142280},
  {32'h4474d148, 32'h44ae270c, 32'h44aca3c7},
  {32'hc51a01a3, 32'h43156622, 32'hc44b05d2},
  {32'h44ccf5df, 32'hc3ae2e4d, 32'hc2757c0e},
  {32'h432f52b3, 32'h44ad2e4e, 32'h433d4920},
  {32'hc4c97564, 32'hc443af51, 32'h4376cb29},
  {32'h453a315e, 32'h4398c84d, 32'h4410e3cf},
  {32'hc53e4663, 32'h43b4a04d, 32'h43c3d20d},
  {32'h44c3e122, 32'h44246357, 32'hc235fff7},
  {32'hc48aff03, 32'hc4719015, 32'h418e816c},
  {32'h4458a909, 32'h4410bcbb, 32'hc41cb90e},
  {32'hc49913ce, 32'hc2c4ab65, 32'hc3c6e074},
  {32'h44dfe99e, 32'hc3929bfa, 32'hc33ae1dd},
  {32'hc497bbd1, 32'hc34f51a1, 32'hc321ede4},
  {32'h45058b6f, 32'h43a662ab, 32'h435e0bac},
  {32'hc4540e7b, 32'hc4887d76, 32'h4309ac9f},
  {32'hc4a76b27, 32'h4324f77e, 32'hc3b5cbf5},
  {32'hc3849983, 32'hc315207b, 32'h44f023f4},
  {32'h4506d8b8, 32'h43ec5918, 32'h43b19506},
  {32'hc4a56216, 32'hc3a8e367, 32'h4179c5a0},
  {32'hc13475e6, 32'hc3bf44c6, 32'hc41f15fe},
  {32'hc525761a, 32'h43414719, 32'h4335d602},
  {32'h43fdddd7, 32'h43ea4a82, 32'hc47fe91e},
  {32'hc419e358, 32'hc450801c, 32'h43c171ad},
  {32'h43025b48, 32'h44804d7d, 32'hc3c0d90b},
  {32'h442bac5c, 32'h43534a27, 32'h44a36dc3},
  {32'h43df7e08, 32'h443c60f0, 32'hc4d5d0bd},
  {32'h438ee6fd, 32'hc2810267, 32'h45138bf2},
  {32'hc48976da, 32'h43533ec8, 32'hc1a9b978},
  {32'hc4ce5b5d, 32'h43cfbe86, 32'h4520c890},
  {32'h44822169, 32'hc3791126, 32'hc4d55609},
  {32'hc2c81d60, 32'hc5376e39, 32'h432304b6},
  {32'hc435567c, 32'h44296ee3, 32'h4439a26c},
  {32'hc387f5ac, 32'hc3999428, 32'hc3fae104},
  {32'h439257c8, 32'h44c2d544, 32'hc3ad1f5e},
  {32'h43fcac52, 32'hc4e35dfb, 32'hc3c97258},
  {32'hc464bbfa, 32'h42b322d8, 32'hc3aa03a6},
  {32'hc3a4cb7e, 32'hc39732a4, 32'h429e71e3},
  {32'hc44ff9ca, 32'hc3d528f1, 32'h43a925fd},
  {32'h44e8f70e, 32'hc2f7e36c, 32'h432e7ffa},
  {32'hc4d0df8d, 32'hc1424b7f, 32'h440c577d},
  {32'h4402d054, 32'hc3dc78ac, 32'h43663910},
  {32'h43a74670, 32'h4496f4b0, 32'hc3688dab},
  {32'h44911004, 32'hc404f518, 32'h4489d9da},
  {32'hc3f847f4, 32'hc2da534f, 32'hc516cb01},
  {32'h4393e761, 32'hc4b57f92, 32'h43701a12},
  {32'hc49f3c82, 32'h44410e26, 32'hc2c4cbe1},
  {32'h4440944c, 32'h43a37b48, 32'h436c4650},
  {32'h43e0c414, 32'hc33ad776, 32'hc4ac3b87},
  {32'h44a4231c, 32'hc4961e16, 32'h433dbb5d},
  {32'hc41a23d4, 32'h44721359, 32'hc4a5c8ca},
  {32'h44a6227b, 32'h41daaaf0, 32'hc2869f40},
  {32'hc42586d5, 32'h44054dd7, 32'hc40f8077},
  {32'h445ce292, 32'hc3a39b02, 32'h43e160f8},
  {32'hc531353c, 32'hc3a4e7a8, 32'hc1b76883},
  {32'h4532600a, 32'hc156a1d6, 32'h443126ec},
  {32'hc3fafd70, 32'h42620d75, 32'hc3fb7aaa},
  {32'hc41229c6, 32'h439babd0, 32'h43b0387a},
  {32'hc4d78357, 32'h43547a60, 32'hc44ea24a},
  {32'hc4523bc2, 32'h445da13b, 32'h44d710a2},
  {32'hc4882275, 32'hc398ba46, 32'h43041c1e},
  {32'hc3c36326, 32'h4354fd80, 32'hc2f209ba},
  {32'h4431254c, 32'hc4a6b08c, 32'h426d2bc2},
  {32'hc4aa1f41, 32'h4254e848, 32'hc340eeb0},
  {32'h4361c554, 32'hc435fd21, 32'h441c778c},
  {32'hc35dcd20, 32'h43edf5b0, 32'hc4f7f4f5},
  {32'h42e9ccf8, 32'hc52af826, 32'h43b2075f},
  {32'h450753db, 32'hc487a866, 32'h44698760},
  {32'hc4e4f998, 32'h44a3cc34, 32'hc48cb217},
  {32'hc30306fd, 32'hc4a42999, 32'h4487662b},
  {32'hc43a0c2d, 32'h43a20ef2, 32'h4455ba91},
  {32'hc4946c2c, 32'h4361f7c3, 32'hc44b223e},
  {32'h42b52d61, 32'hc45f7ceb, 32'h44945bb8},
  {32'h450cd9b0, 32'h42aad780, 32'h42e292d7},
  {32'h450e67ab, 32'hc3f9c2de, 32'hc113167c},
  {32'hc46ad1f4, 32'h4470e698, 32'hc38b83c1},
  {32'h453181be, 32'h423eca8a, 32'hc3418b36},
  {32'hc599dd3f, 32'hc38d0e0f, 32'hc2d43274},
  {32'h455483e8, 32'h4214a6e4, 32'h4413c86c},
  {32'h442cd856, 32'h44ce3777, 32'hc1a77509},
  {32'h4339aae8, 32'h437d3999, 32'h43bb1c07},
  {32'h42218040, 32'h4486310e, 32'h412bb673},
  {32'h44c55911, 32'h426fee30, 32'h4307af2a},
  {32'hc50df17a, 32'h445dfee1, 32'h44347147},
  {32'h4554d586, 32'hc42d6ae1, 32'h42b9c28e},
  {32'hc3ea66e7, 32'h44a298f8, 32'h436493a9},
  {32'hc41a03a8, 32'hc4150019, 32'hc42a5629},
  {32'hc3122d26, 32'hc4f8a26e, 32'h4508084b},
  {32'h438c354e, 32'hc402976e, 32'h44e9f687},
  {32'h450e4ee6, 32'h4265472d, 32'hc21fe056},
  {32'hc45ebbba, 32'hc41f25c3, 32'hc3011100},
  {32'hc336a78d, 32'h442cc82d, 32'hc5343469},
  {32'hc3a94722, 32'h41d8eb99, 32'h44c8171a},
  {32'h43998926, 32'h44e3b67d, 32'hc2579003},
  {32'h44a3bc3a, 32'hc4211124, 32'h42d6b85f},
  {32'hc3be0d6e, 32'hc425f15b, 32'h4508033a},
  {32'hc38fe610, 32'hc4cc673a, 32'hc5038519},
  {32'h41d91bd0, 32'hc29bf574, 32'hc531dd7c},
  {32'hc3daab56, 32'hc5031698, 32'hc20f942f},
  {32'hc2d971ee, 32'h443baf02, 32'h43707d12},
  {32'hc3e1045e, 32'hc4d00937, 32'h42d5dcf1},
  {32'h44b92d2f, 32'h42e8f67e, 32'hc2879c97},
  {32'h4446b6d0, 32'h4138b608, 32'h4400784a},
  {32'h44ecdfca, 32'hc3e57a5d, 32'hc4116eb3},
  {32'hc559b125, 32'h430a158f, 32'h42fb52c5},
  {32'hc46b5b4d, 32'h42550897, 32'hc3be2693},
  {32'hc402196d, 32'hc547a36e, 32'h43436d58},
  {32'h4461e26b, 32'h44d719c2, 32'h43d3f4e7},
  {32'hc407507c, 32'hc3bec17e, 32'h4384c6fd},
  {32'hc2427dc0, 32'h457859f0, 32'h43651feb},
  {32'hc50d7012, 32'hc455d71a, 32'h4322a428},
  {32'hc3e03d4f, 32'h44377c8f, 32'h435550b0},
  {32'h41714cf8, 32'hc336382c, 32'h420cf34d},
  {32'h431a96ba, 32'hc40a603c, 32'hc34af88e},
  {32'h4413a82b, 32'h451efc16, 32'h43c52293},
  {32'h445f8762, 32'h42bb1ad5, 32'h43a412c5},
  {32'h44ce151c, 32'h43918df1, 32'h443adb4e},
  {32'hc4026426, 32'hc4539d60, 32'hc4267e5d},
  {32'h43b63566, 32'h42eb0018, 32'h40ef00df},
  {32'hc503acea, 32'hc39cad3e, 32'hc465a3dd},
  {32'h4323c7ad, 32'h44ac5bb7, 32'h44dff443},
  {32'h4445399a, 32'hc3be1915, 32'h437c0f5e},
  {32'h41401838, 32'hc48e6c26, 32'h44ea9e97},
  {32'h43fe9705, 32'h44cb5aa3, 32'hc4a7d85f},
  {32'hc4c0acbe, 32'h438550e3, 32'h43428bd3},
  {32'h43239847, 32'hc12fb8b0, 32'hc4bcac19},
  {32'h4416a09a, 32'h454ca848, 32'h42d0862a},
  {32'h44e58fcb, 32'h3fcc6a70, 32'hc365f593},
  {32'h4491a136, 32'hc1c1753e, 32'h4464bb32},
  {32'hc4e00103, 32'hc419efe0, 32'hc49d1166},
  {32'h44fa6ddd, 32'h42fad8cf, 32'h43970317},
  {32'hc49cad92, 32'hc4b1ab0b, 32'hc456905e},
  {32'h4403b318, 32'h4502ab11, 32'hc3269a11},
  {32'hc3ac4fec, 32'h43ace908, 32'hc34155ce},
  {32'h441348ef, 32'h4507d167, 32'h439291e0},
  {32'hc38102aa, 32'hc503f660, 32'h438e32b8},
  {32'h45601258, 32'h43e8c40f, 32'h43fce7cf},
  {32'hc40a9938, 32'hc3d9b28c, 32'hc414f591},
  {32'h455105bf, 32'hc3b8fe50, 32'hc35a4b57},
  {32'h4337b6f4, 32'hc40f25dd, 32'hc4b2ec60},
  {32'hc400ddd8, 32'h446a830e, 32'h4489b334},
  {32'h43492dc2, 32'h44a507ad, 32'hc4440741},
  {32'hc4a3b22f, 32'h43a8b44f, 32'h44567429},
  {32'hc24cc958, 32'hc48cd7f2, 32'hc4dbc3a6},
  {32'hc50d9350, 32'hc30d7e80, 32'h428297ab},
  {32'h428bb657, 32'hc3de16d8, 32'hc501adbf},
  {32'hc51b2d3c, 32'h438736b0, 32'h442a0619},
  {32'h44872d55, 32'hc3078361, 32'hc33f2988},
  {32'h42b204de, 32'h441536a7, 32'h4370bb8b},
  {32'hc349fffc, 32'hc406c926, 32'hc3c3e03b},
  {32'h43cde71a, 32'h4315d994, 32'hc2e83738},
  {32'h44358019, 32'hc3933f11, 32'hc44d45c4},
  {32'hc3cf9a00, 32'h451901c5, 32'h4206e54f},
  {32'h442f04d1, 32'h42e6d9b5, 32'hc443aa94},
  {32'hc4ddafbc, 32'h43b59b27, 32'h43d706b4},
  {32'hc4189a14, 32'h436eeed1, 32'hc5656978},
  {32'hc4089812, 32'h43433f82, 32'h437a2857},
  {32'h446caa24, 32'hc4dae9d0, 32'hc26fbcb4},
  {32'hc4612724, 32'h44663998, 32'h4412ae52},
  {32'h45065e3e, 32'h4400384c, 32'h428e3738},
  {32'hc4ade623, 32'h44d087d8, 32'h4198fbb9},
  {32'h445ff26c, 32'hc5371062, 32'hc390c8c8},
  {32'hc47d8780, 32'h434cf4f2, 32'h4305db31},
  {32'h44892f08, 32'h437396c6, 32'h42d4702e},
  {32'hc376d950, 32'hc3d8f5f7, 32'h43d0ad87},
  {32'hc4618550, 32'hc3c42230, 32'hc44dc7c4},
  {32'h44ced8ba, 32'h42b77b61, 32'h4400dfdc},
  {32'hc56df9ac, 32'hc38cad77, 32'h421dc38c},
  {32'h43a6dd8a, 32'hc31a6285, 32'h4517bc94},
  {32'hc53eff41, 32'hc1e50cdb, 32'hc3b1bdc6},
  {32'h44fc56a2, 32'hc308dfed, 32'h4143162c},
  {32'hc470f9c6, 32'h43be0591, 32'h42aaf9e2},
  {32'h4465202c, 32'h43426868, 32'hc397fb8e},
  {32'hc4c5c5dc, 32'h44b5f54a, 32'h421a9f4b},
  {32'h4514f56c, 32'hc42cd92a, 32'hc36b68df},
  {32'h44676db4, 32'h43f0f00d, 32'h42d61401},
  {32'h44072e04, 32'h4202d7d7, 32'h44dede53},
  {32'hc5255067, 32'h43de42bd, 32'hc3d66f3d},
  {32'h44335dc7, 32'hc43cdc7d, 32'h43504ea2},
  {32'hc3f2d3ec, 32'h44abb501, 32'h444d65cf},
  {32'h3f84c56c, 32'hc3b9e4c2, 32'hc4b28d0f},
  {32'hc4cfb324, 32'h43abb368, 32'h4407cc78},
  {32'hc28822e0, 32'h43f04130, 32'hc481b301},
  {32'hc3de4a94, 32'h438bfc9a, 32'h44694ed6},
  {32'h455b3284, 32'h4241b17a, 32'hc391c11f},
  {32'hc4832d1d, 32'h445b16f2, 32'h44138d7e},
  {32'h449b2d43, 32'hc12568c6, 32'hc3ff95f7},
  {32'hc4d1bd3b, 32'hc376f8a3, 32'hc3d6b612},
  {32'h430f7b25, 32'hc4141b0b, 32'hc49ac6d2},
  {32'h41a757b0, 32'h44f2da59, 32'h442ba19a},
  {32'hc3ecf5fd, 32'hc3274c4d, 32'hc489f602},
  {32'hc519bda8, 32'h442de886, 32'h444eb38a},
  {32'hc274272a, 32'hc4775967, 32'hc4dc46f6},
  {32'h4523cc9d, 32'hc1ca3bed, 32'hc3c2b188},
  {32'hc56ae044, 32'hc40f34be, 32'hc0e32d50},
  {32'hc486865d, 32'h4321b5be, 32'h4393943f},
  {32'hc3b4c679, 32'hc534a8cc, 32'hc3087134},
  {32'h42021c00, 32'h43927aa5, 32'h431a375c},
  {32'h4336e9da, 32'hc52edc24, 32'h432d2400},
  {32'h44619d8c, 32'h45210e13, 32'h441207ea},
  {32'hc4a97b90, 32'hc4d55a01, 32'h42d148d9},
  {32'h44e43a48, 32'hc3c9f47d, 32'h434cbd00},
  {32'hc493865f, 32'hc3c7a0fc, 32'h43937807},
  {32'h440418a9, 32'h43dda3fc, 32'h43be0095},
  {32'hc4b48106, 32'hc282a58d, 32'h43ea38f5},
  {32'h445f5520, 32'h4524597d, 32'h437aa397},
  {32'hc2d0923b, 32'hc4926446, 32'hc5024e7f},
  {32'h43984e16, 32'h4336f02a, 32'hc23ba0e9},
  {32'hc242b6d0, 32'hc3bcbc4a, 32'hc4d1e5a2},
  {32'h446063bc, 32'h44bab518, 32'h44057430},
  {32'hc3b6278a, 32'hc3ce4f4b, 32'h42fd9c3f},
  {32'h44bd2830, 32'hc4484cf5, 32'h441c4b22},
  {32'hc3729440, 32'h4462ab87, 32'hc4d04223},
  {32'h440148f3, 32'h4382b084, 32'h43642638},
  {32'hc3350f9c, 32'hc55445c1, 32'hc412125b},
  {32'h44a3608c, 32'h449cef99, 32'h43ed7772},
  {32'h44bc7aef, 32'h42af97ee, 32'h4399588c},
  {32'h4443edf6, 32'h43cb21ad, 32'h4492ab95},
  {32'hc487768a, 32'hc3a27f2e, 32'hc5395a2e},
  {32'h44d2744a, 32'hc2aa7e37, 32'h428390e0},
  {32'h437eeae4, 32'h44a95a71, 32'hc35465c2},
  {32'hc43f1ce0, 32'hc4cca3d3, 32'h4363e98f},
  {32'hc293e560, 32'h44d8ec9c, 32'h43648e04},
  {32'hc4a90dc2, 32'hc421441d, 32'h4402f719},
  {32'h44196012, 32'h44812fdb, 32'hc2d21006},
  {32'hc4fb1448, 32'hc4389f48, 32'hc31aa43b},
  {32'h4440493f, 32'h43c65735, 32'h421d385d},
  {32'hc58a1941, 32'hc31edd7e, 32'hc370f292},
  {32'h45371f21, 32'hc3a845a2, 32'h437d51be},
  {32'hc40e73cf, 32'hc28baa2f, 32'h43e2cb0e},
  {32'h44994ef4, 32'h44476434, 32'h43f563b0},
  {32'hc520a92a, 32'hc37eb838, 32'hc1a2e980},
  {32'hc2ea78a0, 32'h432c00c3, 32'hc4d69916},
  {32'hc3a03eb1, 32'hc3b6f39b, 32'h44cc95ff},
  {32'h452bf719, 32'h43c235de, 32'h43c40169},
  {32'hc3065385, 32'h43861fb3, 32'h44a7baf5},
  {32'h43b33030, 32'hc3350d17, 32'hc4d3a920},
  {32'hc156b44c, 32'h43fec907, 32'h455e54d3},
  {32'h44936c61, 32'h42e7f58f, 32'hc32ac3ad},
  {32'hc4288d67, 32'hc4bc74ac, 32'h44bc88c7},
  {32'h44bf232f, 32'h445f0b05, 32'hc412d103},
  {32'h44c5e40a, 32'h43199418, 32'h42a9b56e},
  {32'h432d450a, 32'hc34105a7, 32'hc281569b},
  {32'hc3c984e2, 32'hc4958436, 32'h436639d1},
  {32'hc47bc52a, 32'h42436c6b, 32'hc2ed7bd3},
  {32'hc44b18ba, 32'h440f4b97, 32'h454a0582},
  {32'h4570f8cc, 32'hc3911d7c, 32'hc4628d6b},
  {32'hc3a21c23, 32'hc49acf10, 32'h43962219},
  {32'hc4f17698, 32'h420dcd82, 32'h448a22f7},
  {32'h43c021ee, 32'hc5037f4d, 32'hc2ff7b33},
  {32'hc42536cc, 32'h414202cb, 32'h440e7a17},
  {32'h44dc4030, 32'hc43aba3c, 32'h43a2e768},
  {32'hc42725bc, 32'h447ab2b6, 32'hc39751da},
  {32'h45498d70, 32'hc3d34413, 32'hc42a384e},
  {32'hc558558c, 32'hc2c2ae6d, 32'hc40047f7},
  {32'hc36b7a74, 32'hc3657025, 32'h440324fc},
  {32'h42daf774, 32'h4532a625, 32'h3f0ef270},
  {32'h4446f1e4, 32'hc3ec01dc, 32'h45001166},
  {32'hc43edf76, 32'h43417a4c, 32'hc4070bc7},
  {32'h43a8da32, 32'hc522b551, 32'hc1b98c86},
  {32'hc43c3d8a, 32'h4211994a, 32'hc49319df},
  {32'h449cacc0, 32'h431d7e50, 32'h438dab29},
  {32'hc4099c93, 32'hc3889e15, 32'hc5216e28},
  {32'h44ac1c2a, 32'hc30fff31, 32'h443352e0},
  {32'h44c79514, 32'h43d97421, 32'h43ba966d},
  {32'h4508471c, 32'hc493e53d, 32'hc4006de5},
  {32'hc5385bff, 32'h44a0216d, 32'hc4375224},
  {32'hc3a1c6eb, 32'hc3bd20a3, 32'h44d3d32a},
  {32'hc4a3af1c, 32'h4405025f, 32'hc457c8bc},
  {32'h44424134, 32'hc46c9edf, 32'h4402abad},
  {32'h442c3bc7, 32'hc338f359, 32'hc124aa8c},
  {32'h44da618a, 32'h435cf761, 32'h447d297c},
  {32'hc54cfdc2, 32'h43426fd2, 32'h433cb059},
  {32'h444925fb, 32'h432504ef, 32'h449df32a},
  {32'hc4899fd2, 32'hc349b3a6, 32'hc49c68a2},
  {32'h43c3aee4, 32'hc478d94b, 32'h446a1903},
  {32'h4334145a, 32'h44956e0f, 32'hc42d1b63},
  {32'h43989a73, 32'h437b89e3, 32'hc4949758},
  {32'h446f431e, 32'hc3f9aaa5, 32'h43ee821c},
  {32'hc41a8150, 32'h431c7b16, 32'hc4d250c9},
  {32'hc4b700c6, 32'h42cb46ad, 32'hc3d8f58a},
  {32'hc44a27d0, 32'h442537f9, 32'hc4ba26fe},
  {32'h4384b7ef, 32'hc3fe596b, 32'h4523e935},
  {32'hc38c7802, 32'hc457222b, 32'h452d0734},
  {32'hc4566a05, 32'h44dc70c6, 32'hc4b83853},
  {32'hc3a6bd48, 32'hc48f3870, 32'h44ac7ec2},
  {32'h43a89255, 32'hc3085442, 32'h434bb273},
  {32'hc540713a, 32'h435ebbb2, 32'hc29a17db},
  {32'h44480a13, 32'h42ab644b, 32'h449e9859},
  {32'hc51a984a, 32'hc3e6c0e0, 32'h43bf82ef},
  {32'h4485bdf6, 32'hc43217c5, 32'h447d66b4},
  {32'hc2ff6b1c, 32'hc2ef3176, 32'hc4cf9915},
  {32'h43809942, 32'hc3fc1fa5, 32'h42f6e0d6},
  {32'hc444232b, 32'hc43948a2, 32'hc46f8944},
  {32'h4495c440, 32'h443f760b, 32'h43372604},
  {32'h44cfe9df, 32'h4240cd20, 32'hc3a54032},
  {32'h430a9760, 32'hc3e59e78, 32'hc1e2efa8},
  {32'hc4dda68c, 32'h42d1e556, 32'h430f2ffa},
  {32'h4348d986, 32'hc4b25e38, 32'hc3b3eb69},
  {32'hc575d9b0, 32'h43f9b877, 32'h4353654e},
  {32'hc31e8790, 32'hc56baa3f, 32'hc401ab44},
  {32'hc3411760, 32'h4495931f, 32'h43a3ae2e},
  {32'hc38fdc82, 32'h4475f278, 32'hc51e70ff},
  {32'h43ad3474, 32'hc499d3a4, 32'h448e210f},
  {32'hc32645e4, 32'hc0ff52c8, 32'h4521b6a6},
  {32'h450a18ea, 32'h43537dde, 32'h4314bcdd},
  {32'hc45bd990, 32'h4346820b, 32'h4493b163},
  {32'h44393102, 32'h42c5a344, 32'hc4eb871e},
  {32'hc392ae9c, 32'h4319f677, 32'h4538c725},
  {32'h4550422d, 32'hc3a25dd8, 32'h43b8805f},
  {32'h43854c1f, 32'hc4ab5d8b, 32'hc33c4d4b},
  {32'hc4aa4806, 32'h4248342b, 32'h44138343},
  {32'h450dc2f5, 32'hc43be70a, 32'hc441c2b6},
  {32'h44376dc6, 32'h4496c7a1, 32'hc34f297d},
  {32'hc461a18c, 32'hc3d2cf29, 32'h4498a675},
  {32'hc34d3c71, 32'h4381cbdc, 32'hc4c12a79},
  {32'hc41dad03, 32'h430e86d1, 32'h454657c2},
  {32'hc40623f4, 32'h439f77f6, 32'hc54c7379},
  {32'h448017d8, 32'h42673e26, 32'h4357416f},
  {32'h44feecbc, 32'h43c1ecb3, 32'h432b46d8},
  {32'hc578a0be, 32'h41b21024, 32'h4315d0a8},
  {32'hc42a6573, 32'h439134b8, 32'hc3d80732},
  {32'hc539a1c2, 32'hc421cf7f, 32'hc3ddcefb},
  {32'h438b4258, 32'h450e31e6, 32'hc3912cb9},
  {32'hc45ee0a8, 32'hc3b0b208, 32'h43c1ad84},
  {32'h4488eab3, 32'h44cc5a05, 32'h43ebf641},
  {32'hc569c245, 32'hc38a1532, 32'h429971cb},
  {32'h42c60569, 32'h44238222, 32'hc2ccb30b},
  {32'h44c93286, 32'hc39f3cfb, 32'hc1982d24},
  {32'hc3a7e322, 32'hc39fac75, 32'hc4ae3342},
  {32'hc372facd, 32'hc46bc6c7, 32'h450e1c07},
  {32'hc1f1476f, 32'h42219a80, 32'hc4ad8e79},
  {32'h452eb44f, 32'hc314213e, 32'h4393d798},
  {32'hc4a76996, 32'hc474187f, 32'h41a55170},
  {32'h43c947d0, 32'h431af5e6, 32'h435a96f3},
  {32'hc32c7409, 32'hc14e66c8, 32'h4334ba94},
  {32'h44ab61cf, 32'h442eac4e, 32'h43c54b51},
  {32'hc4de4a92, 32'hc395167b, 32'h43e3a077},
  {32'hc47f81ee, 32'hc40729bc, 32'h44984ea0},
  {32'hc39547dc, 32'h442564f1, 32'hc4d8ac6e},
  {32'h44059c20, 32'h40c3e084, 32'h44a5baf9},
  {32'hc409c07a, 32'hc26170bd, 32'hc2ed1341},
  {32'hc34a365b, 32'h438d9ea1, 32'h45040d13},
  {32'h43827de4, 32'hc2be612c, 32'h43ec3d54},
  {32'h42b98d08, 32'h441df11c, 32'h4541fe4c},
  {32'h4349ab44, 32'hc49c5974, 32'hc54b55d9},
  {32'hc3445a2a, 32'h449b6573, 32'hc3e0d1d4},
  {32'hc3bf4426, 32'hc5791544, 32'hc32b6498},
  {32'h44fb1af6, 32'h4476e969, 32'h440749d6},
  {32'h44fcef5f, 32'hc38ed320, 32'hc2565357},
  {32'h44d7a2b9, 32'h44a30b42, 32'hc2f6de00},
  {32'hc396f11e, 32'hc57580cf, 32'hc3a88915},
  {32'h4570aa30, 32'h4402e9f1, 32'h43d0d3cb},
  {32'hc59057e8, 32'h419336f1, 32'hc3c53bcc},
  {32'h44293018, 32'hc44a5f47, 32'hc43f4198},
  {32'h4423b336, 32'h419dced3, 32'hc433c094},
  {32'h43da9ebd, 32'h4468a8a7, 32'h44ac7517},
  {32'hc1a11a0c, 32'h442505ac, 32'hc48316f8},
  {32'hc44215aa, 32'h442155d9, 32'h440be4e5},
  {32'hc3aa55bd, 32'hc4479a83, 32'hc4cc7f50},
  {32'hc4c08eb4, 32'h441e0c5c, 32'h43fd0e56},
  {32'h44551469, 32'hc4e040b6, 32'hc4a87df5},
  {32'hc4bf581e, 32'h430bbe3e, 32'h44a17186},
  {32'hc459ee63, 32'hc3bd1ec1, 32'h42810089},
  {32'hc4896b95, 32'hc4141136, 32'h4489f744},
  {32'hc3426e7c, 32'h444d017f, 32'hc50f486b},
  {32'h44111f4e, 32'h42981b5f, 32'h434fd5ab},
  {32'h4427b4e4, 32'h426ce47e, 32'hc40d27f1},
  {32'hc41402de, 32'h43b625bf, 32'h44c5f4f2},
  {32'h4395b4ea, 32'hc1750104, 32'hc48fd274},
  {32'hc4b24236, 32'h428ae8d9, 32'h445775e0},
  {32'h44ca81f6, 32'h4334cf4a, 32'hc375b572},
  {32'hc41d0546, 32'hc3ef139f, 32'h43861ed1},
  {32'h44a0f957, 32'hc50d7ab0, 32'hc21e4b92},
  {32'hc4b63801, 32'h448c7a06, 32'h430f58a4},
  {32'hc2e9b3f0, 32'hc32f95bb, 32'hc2826d58},
  {32'hc4207b10, 32'hc3405896, 32'hc3b9e042},
  {32'h446a7614, 32'hc4b5beb1, 32'hc34641d8},
  {32'h44f77079, 32'h42e1dbed, 32'hc218daf1},
  {32'h45362b10, 32'h43f71978, 32'hc2cac091},
  {32'hc45206b6, 32'h4212ad0c, 32'h43a67ade},
  {32'h4583b2ac, 32'hc3861a52, 32'h440fd5c0},
  {32'hc497efe6, 32'h435904db, 32'h443fa601},
  {32'hc54140c0, 32'h4302eb85, 32'hc41a9161},
  {32'h44caa490, 32'h43692a3c, 32'h43a7876c},
  {32'h42430d20, 32'h4396be15, 32'hc3ae91aa},
  {32'h440962cf, 32'hc51defe6, 32'hc2e95360},
  {32'hc3f7d75a, 32'h43b27bec, 32'h439f0ba3},
  {32'h44b339d0, 32'hc34712a1, 32'hc3a48e9f},
  {32'h43a08ffd, 32'h45434964, 32'h43ee3e29},
  {32'h44a41cfd, 32'hc43eb9e2, 32'h43c1af5d},
  {32'h45044738, 32'hc403f0ce, 32'hc3c57877},
  {32'h442242ea, 32'hc3d57907, 32'h44c257ee},
  {32'hc489ffee, 32'h43009f1c, 32'hc4995c7e},
  {32'h445480ea, 32'hc3bbe9b5, 32'h411cbb6c},
  {32'h42c3fd72, 32'h45320a5b, 32'h43d093a0},
  {32'h43fb78ad, 32'hc31d9c09, 32'hc4cfa15e},
  {32'hc43a010c, 32'h436931c2, 32'h43c358ea},
  {32'h44d236b0, 32'hc4858b9b, 32'h4286d8d0},
  {32'hc4cf1013, 32'h42a3b4f3, 32'h448d3804},
  {32'hc3433ad0, 32'h42445eca, 32'hc41497ee},
  {32'hc579e060, 32'h4382c3f6, 32'h43892e54},
  {32'h45095d14, 32'h41c9e7b2, 32'hc44b9214},
  {32'hc3b19283, 32'h43251c9a, 32'h4492705b},
  {32'h44fe81ab, 32'hc4070f42, 32'h4288d3aa},
  {32'hc38b2940, 32'h44cdadd8, 32'h44cf8956},
  {32'h440f64fc, 32'hc35c6450, 32'hc4a869a8},
  {32'hc2e9e155, 32'h45261cd0, 32'hc340ae8f},
  {32'h42376140, 32'hc4dae46b, 32'hc4049232},
  {32'h44b782c4, 32'hc381b07d, 32'hc4dd42d5},
  {32'hc51cc849, 32'h43260db2, 32'hc2c73802},
  {32'hc3ae98c2, 32'h43bf5268, 32'h43ec2b72},
  {32'hc50027ec, 32'hc3d25e29, 32'hc3533851},
  {32'h44a9fa31, 32'h4411dd0f, 32'hc3d3f5fa},
  {32'hc44ba0ca, 32'hc4a21283, 32'h43bae261},
  {32'h449525da, 32'h44acd4f6, 32'h43bcb5e8},
  {32'hc43adff6, 32'hc458df44, 32'h43904880},
  {32'h44223bcc, 32'h448519e0, 32'h43e3b951},
  {32'hc4227820, 32'hc40448bb, 32'hc3f42306},
  {32'hc266e2a0, 32'h4387d88f, 32'hc28813bf},
  {32'hc50d6281, 32'h4196334e, 32'h43abccf8},
  {32'h43ea9852, 32'h44b7588e, 32'h442dc3ce},
  {32'h4121e028, 32'hc524a24e, 32'hc41b6be0},
  {32'hc3a0ce46, 32'h4487a6c5, 32'h440d78f1},
  {32'hc372d79d, 32'hc4aa9209, 32'h42d0a56c},
  {32'h443a8ce0, 32'h44d5d6c1, 32'h446514dc},
  {32'h449ad4d6, 32'hc40ce8b0, 32'hc30a87d1},
  {32'h44d894d6, 32'hc40e80d6, 32'h43ca76f5},
  {32'hc40845e2, 32'hc494c929, 32'hc4eb0c4d},
  {32'h4522170e, 32'h430d4a0b, 32'hc3ff79dc},
  {32'hc3c313e4, 32'hc4510cdd, 32'hc4b8d9f1},
  {32'h438e901f, 32'h44999d0b, 32'hc1cf32ca},
  {32'hc3888dd6, 32'hc451300e, 32'hc3d6fcaa},
  {32'hc3adbb9b, 32'h44ba3389, 32'h4376b7b9},
  {32'hc43637d4, 32'hc3fc8f74, 32'hc53c78f3},
  {32'h451a42ce, 32'hc2ce6ef8, 32'hc2b2e27d},
  {32'h44b6bb98, 32'h43253aca, 32'hc3089fbd},
  {32'hc42435b4, 32'hc5040080, 32'hc3b00aca},
  {32'hc35a3902, 32'h454c6685, 32'hc311fd05},
  {32'h44d5d6d3, 32'h432832b7, 32'h4234be82},
  {32'h45055d30, 32'h439bfdea, 32'hc3d31016},
  {32'hc4800fc0, 32'hc4ae4afa, 32'hc39569bd},
  {32'h453c70d8, 32'h43f32357, 32'hc3047664},
  {32'hc51d39a0, 32'hc462a7cf, 32'hc3ea5762},
  {32'h45072ca7, 32'h441934cf, 32'h438b9409},
  {32'hc480cf2b, 32'hc3f2f46b, 32'h43e78b1b},
  {32'h435bcbd0, 32'h44ebe47c, 32'hc36a65df},
  {32'hc4043924, 32'hc4a07dcb, 32'hc312209e},
  {32'h44cc0824, 32'h43b0d855, 32'hc113572e},
  {32'hc5304156, 32'hc369cc58, 32'h43853fe6},
  {32'h443abb13, 32'h44bd8728, 32'hc408bb5d},
  {32'h421279ec, 32'hc3d1e992, 32'h42cf64f5},
  {32'h44fef762, 32'hc422cfeb, 32'hc437a34d},
  {32'hc507c99c, 32'hc3b79913, 32'hc38c71ad},
  {32'h44a5d84a, 32'hc30ceb40, 32'hc4213f2c},
  {32'hc4cc034a, 32'hc4550066, 32'h43e2e5d7},
  {32'h44b4f092, 32'h44463bbf, 32'hc4c72c4c},
  {32'hc528f286, 32'hc2c94c56, 32'h42abe2a2},
  {32'h442e0b6e, 32'h447d4407, 32'hc4002aff},
  {32'h43878c35, 32'h43be332f, 32'h452279a3},
  {32'hc414eabb, 32'hc34158f7, 32'hc486bf53},
  {32'hc4c2abd9, 32'h4446f56d, 32'h45060f9a},
  {32'h448256a4, 32'hc3db275b, 32'hc53c0981},
  {32'h4400afaa, 32'hc4ab8a91, 32'hc3f96f7f},
  {32'hc368cd19, 32'h451ebc1c, 32'h4359e86a},
  {32'h44716166, 32'hc3e3619f, 32'h431680d8},
  {32'hc5029e68, 32'h44afdd61, 32'h43a0e827},
  {32'hc22f6318, 32'hc4d98c8e, 32'hc2ef4c8c},
  {32'h431f6408, 32'h43f3a59b, 32'h4185a834},
  {32'hc2ef4d00, 32'hc45708f9, 32'hc41ca20e},
  {32'hc5861e78, 32'hc39918b4, 32'h43a3abd7},
  {32'h4417693e, 32'hc2f4a258, 32'h431845f7},
  {32'hc515b5d9, 32'h43a17b9b, 32'hc44c69ee},
  {32'h450899be, 32'hc2b3f545, 32'hc2b671c8},
  {32'h4422be00, 32'h442006e5, 32'hc2bf8c9d},
  {32'h43934e20, 32'hc4d0281e, 32'h43bd2996},
  {32'hc4fc5b64, 32'hc42dbc71, 32'hc439be2b},
  {32'h438110cd, 32'hc33a4947, 32'h444510a1},
  {32'hc49e44e9, 32'hc3a1103a, 32'hc4a72909},
  {32'h44005d90, 32'h43823893, 32'h451c50eb},
  {32'hc452b54a, 32'hc2bc6797, 32'hc3c85c26},
  {32'h4449d452, 32'hc4fc0310, 32'hc2812a64},
  {32'hc28c9798, 32'h44cbbec3, 32'hc42792d8},
  {32'h4442a3bc, 32'hc397d643, 32'hc176877c},
  {32'hc3b5d630, 32'h4509daa4, 32'hc41f3735},
  {32'hc3c264b7, 32'hc41f8b1e, 32'h44e2f32a},
  {32'h4316251e, 32'h442d68f3, 32'hc03ffb98},
  {32'h4541e040, 32'h428cba30, 32'h436e8a4c},
  {32'hc53cb0e0, 32'hc2c4b45e, 32'hc3f6d1d8},
  {32'h455c0fa1, 32'h42a1c13a, 32'hc3d98f2f},
  {32'hc4920781, 32'hc34e4f3d, 32'hc3b3d43b},
  {32'h44216a84, 32'hc4658ba7, 32'h447d31c0},
  {32'h44059d45, 32'h4434cb44, 32'hc415de95},
  {32'h44e70317, 32'h432d01b7, 32'hc417c9fe},
  {32'h446771b1, 32'hc50e46e7, 32'hc3890137},
  {32'hc48a7aca, 32'h43a9e36a, 32'hc3b54c7e},
  {32'h44ad7805, 32'hc3964cbb, 32'h43b1b468},
  {32'hc418d059, 32'h452cb2a2, 32'hc29880c6},
  {32'h450a81cd, 32'hc3b75dbf, 32'h444bdabb},
  {32'h43f2ee18, 32'h43dfe820, 32'h44dc6027},
  {32'h41be960e, 32'hc4261f09, 32'hc4abd565},
  {32'h442e396c, 32'hc41f2d40, 32'h43203b2e},
  {32'h43c171aa, 32'hc455f446, 32'h43de5b0d},
  {32'hc50852af, 32'h42365de6, 32'hc408cd9a},
  {32'h447e0245, 32'h43334994, 32'h44a0300b},
  {32'hc48a3cf2, 32'h43616155, 32'h42b670c6},
  {32'h43452f30, 32'hc4832fc2, 32'h44ea010f},
  {32'hc1cd9780, 32'h44bbbd03, 32'hc36c7c8b},
  {32'h441de2fc, 32'hc2c39765, 32'h425e8560},
  {32'hc54ad3e7, 32'h43cb2f9e, 32'hc3c6a3ea},
  {32'hc35c55ac, 32'h4439ab3b, 32'h43896d5a},
  {32'h44bc4c7b, 32'h446a1feb, 32'h431a8451},
  {32'h4541b3a0, 32'h4426e785, 32'h423e9da7},
  {32'hc4472291, 32'h451c9709, 32'hc2569d21},
  {32'hc3efdbe2, 32'hc3f0d9a4, 32'hc383f348},
  {32'hc467c85c, 32'h44ee62d6, 32'h42612290},
  {32'h427285c0, 32'hc518d0e2, 32'h43b00405},
  {32'h4475502c, 32'hc35eec34, 32'h43fc7612},
  {32'hc3883ac8, 32'hc517784e, 32'hc4f7fc82},
  {32'hc488e70c, 32'hc3d286b0, 32'h442fdf53},
  {32'hc3c334a5, 32'hc49e05b2, 32'h43703f9c},
  {32'h45275cdf, 32'hc35269fe, 32'h43c4683e},
  {32'hc39a35f1, 32'hc4c5c467, 32'h43422546},
  {32'h43f35822, 32'h44ff51d4, 32'hc23f0330},
  {32'hc5074933, 32'h4332a1f1, 32'h43cea733},
  {32'hc384713c, 32'hc25094ce, 32'h428c7aba},
  {32'h44f959bb, 32'h439405e5, 32'h438ab618},
  {32'hc47e7eea, 32'hc43c67ae, 32'h449d693a},
  {32'h4411d73e, 32'h44e7c00a, 32'hc4d89557},
  {32'h4323b4d1, 32'h45136803, 32'h42accb71},
  {32'hc2e26318, 32'hc4730111, 32'h4383f8b9},
  {32'hc353f842, 32'h42c51110, 32'hc4faa6df},
  {32'hc4c3714c, 32'hc36b08ab, 32'h448f4797},
  {32'h43e29380, 32'h43fb6fd0, 32'hc3ea79b4},
  {32'h448e04ce, 32'hc269752c, 32'h4474cdb8},
  {32'h442a1656, 32'hc334e887, 32'hc3e90a5e},
  {32'hc4922552, 32'hc34f1622, 32'h4429bd13},
  {32'h44f1fb72, 32'h441eb7d7, 32'hc2b39f98},
  {32'hc3fc42f3, 32'hc5126848, 32'h42d54118},
  {32'h4527d081, 32'hc29aad33, 32'hc3060325},
  {32'h44169419, 32'hc4518c6c, 32'h4336204f},
  {32'h44a96a1b, 32'h44c33d14, 32'h42fe0e1f},
  {32'hc534a3e8, 32'h43618cb0, 32'h42822c08},
  {32'h44e78c0a, 32'h44057ba3, 32'hc34ece3f},
  {32'h4428e819, 32'hc3d6b827, 32'h42ef944a},
  {32'hc1c00d61, 32'hc3d88b6c, 32'hc4640f69},
  {32'hc36ef3fd, 32'h430f9c9c, 32'h44b6835a},
  {32'h42cef139, 32'hc44c9717, 32'hc3596da7},
  {32'h44075413, 32'h44e47fd2, 32'h43eb5717},
  {32'hc1a0d424, 32'hc404a44b, 32'hc54422c4},
  {32'h451ae9b1, 32'hc20b82ef, 32'h43f2419d},
  {32'hc2ec4520, 32'hc4247bf2, 32'hc50ad6fa},
  {32'h4462f228, 32'h446b0169, 32'h44ccb292},
  {32'hc42513ab, 32'h44ae8d0e, 32'hc29e4c33},
  {32'h433de964, 32'hc47cdbe4, 32'h444d4a25},
  {32'hc2dae0a5, 32'h444b77cd, 32'hc4aed6a5},
  {32'h443613b2, 32'h447ee129, 32'hc2f63e8c},
  {32'hc5334a6a, 32'hc379ab82, 32'h42d40982},
  {32'h42efd558, 32'h44214cb1, 32'h41815637},
  {32'h43f96acc, 32'hc35429de, 32'hc35a0604},
  {32'h44dc1c9e, 32'h434a4318, 32'h448191a6},
  {32'hc53c9ca0, 32'hc22a1aba, 32'hc3826e8f},
  {32'h4329f2b3, 32'hc24d4e78, 32'h438c1926},
  {32'hc472cd1d, 32'hc51a0904, 32'h427a6241},
  {32'h453a3bb6, 32'h4414e322, 32'hc36cef67},
  {32'hc255f9d0, 32'hc3e46640, 32'hc3f936ba},
  {32'h44d273fb, 32'h4462fd26, 32'h43527e7a},
  {32'hc50df1a7, 32'hc381eb69, 32'hc30db07c},
  {32'h4388ff7b, 32'h43988d87, 32'h43ffc10c},
  {32'hc41431ae, 32'h4306a048, 32'h431dd032},
  {32'h432afe5a, 32'h4250cd93, 32'h431a73f8},
  {32'h44868548, 32'hc26eab5c, 32'hc41c2f0c},
  {32'hc4a6e1c1, 32'hc3a05ad4, 32'h444e7405},
  {32'h41285760, 32'h44221ee8, 32'hc4ced598},
  {32'hc3326b70, 32'h44efa8c8, 32'h43dd2516},
  {32'h44b760d4, 32'hc4026316, 32'hc32e96c5},
  {32'h43eb730c, 32'h4387ad02, 32'h447bd1d2},
  {32'h43fa40b9, 32'hc3d0a783, 32'hc4cdcf3d},
  {32'hc2a3fb32, 32'h451389d1, 32'h44f4992d},
  {32'h451fd0c7, 32'h43a6837c, 32'h4318e493},
  {32'hc44ed8a6, 32'h44899242, 32'h44279236},
  {32'hc33a591d, 32'hc4b05e4e, 32'hc3742e94},
  {32'h43571d88, 32'hc381d462, 32'h42d16816},
  {32'h4396c2b0, 32'hc3564395, 32'hc4f946c6},
  {32'hc3422520, 32'h42f1285d, 32'h452ea87e},
  {32'h44dcbcbd, 32'hc0ca573b, 32'hc32ad5ac},
  {32'hc4a4a448, 32'h43a7346b, 32'h44445d5a},
  {32'h441963fb, 32'hc41e94dd, 32'hc3bcf343},
  {32'hc46473f8, 32'h436c0a00, 32'h42db18bf},
  {32'h447db8ca, 32'hc4b52fe9, 32'hc3a11483},
  {32'hc4f160a8, 32'h44658d64, 32'h4262a870},
  {32'h455b7c21, 32'h42e22d4e, 32'h421d4104},
  {32'hc45a83e4, 32'h44e443b4, 32'hc38ddad1},
  {32'h4413e958, 32'hc44f181b, 32'h43dfb299},
  {32'h44b25aa1, 32'h43474b6a, 32'hc16ef32d},
  {32'h44f4ce02, 32'hc1af0772, 32'h419fa47d},
  {32'hc56af9bf, 32'hc2a4227a, 32'h4384a4f1},
  {32'hc4eee2aa, 32'hc3aa70b1, 32'hc3915d37},
  {32'hc2c60020, 32'hc3a81504, 32'h43e47973},
  {32'hc3f6c120, 32'h43281e75, 32'hc49110e2},
  {32'h452af202, 32'h43a190cc, 32'h4420a66f},
  {32'h43e9dd17, 32'h44ca9966, 32'h43644811},
  {32'h44c3b32a, 32'hc46629e3, 32'h43f27ae4},
  {32'hc3c44bd5, 32'h44f7dde9, 32'hc2e251d3},
  {32'hc374a668, 32'hc40c9d43, 32'h42812719},
  {32'hc3ce47eb, 32'h45747889, 32'h439e3f95},
  {32'h43f24cbc, 32'hc53e9200, 32'h4026a150},
  {32'hc3ff017c, 32'hc27613d2, 32'hc45eb8b4},
  {32'h443c65f8, 32'hc0788870, 32'h440c805e},
  {32'hc2d02d00, 32'h435256c0, 32'h43ae5f55},
  {32'h433b3e12, 32'h420f5046, 32'hc5018b4b},
  {32'hc4586db4, 32'hc2812f82, 32'h4401e2c1},
  {32'h442d55c2, 32'hc4078b00, 32'hc4acd0df},
  {32'hc4932452, 32'h42df9583, 32'h43c712b9},
  {32'hc3971732, 32'hc39decd7, 32'hc4d61f13},
  {32'hc38f971c, 32'h44e45601, 32'h4398d31e},
  {32'h451832f4, 32'hc428725a, 32'h43868351},
  {32'hc567f031, 32'h43befa77, 32'h438101bd},
  {32'hc28b89d0, 32'h4496e1cb, 32'hc482cfc4},
  {32'hc4c3d739, 32'hc313427d, 32'hc356277e},
  {32'hc3c74724, 32'hc22a7988, 32'hc5568f33},
  {32'hc3cf54e6, 32'h4386943a, 32'h44b21db2},
  {32'h443eb04d, 32'hc3d71387, 32'hc4926838},
  {32'hc3245688, 32'h43983f7e, 32'h45197bcb},
  {32'hc38db988, 32'hc4b55a8f, 32'hc4563aca},
  {32'h4515d37f, 32'h4158fe7f, 32'hc472ec08},
  {32'hc4c496be, 32'h4248b764, 32'h449c1f75},
  {32'h442d0323, 32'h4453bab6, 32'hc47f6b7d},
  {32'hc4c5b73e, 32'hc4a0fdd2, 32'hc30db1a2},
  {32'h44f7692d, 32'h43abfddd, 32'h43becb12},
  {32'hc4391126, 32'hc311fe20, 32'hc40809cd},
  {32'h4434b860, 32'h4453c68a, 32'hc2bc1baa},
  {32'hc48e54d8, 32'hc4706919, 32'h43debd59},
  {32'h44bb8964, 32'hc32af4da, 32'h43a903a4},
  {32'hc5030782, 32'hc24f4852, 32'h43f0a91a},
  {32'h4492e976, 32'h442807db, 32'h43d5ed1b},
  {32'hc4a26d22, 32'hc242ae5d, 32'h4393615a},
  {32'h44390f67, 32'h4489fc6b, 32'h445602b0},
  {32'hc49270c3, 32'hc4ea80ef, 32'hc48201be},
  {32'hc4ac560c, 32'h43ace635, 32'h43512530},
  {32'hc2d189e6, 32'hc51ec756, 32'hc3769501},
  {32'h43770f7a, 32'h44dde9dc, 32'h43c5f78b},
  {32'h44d9578c, 32'h43a9ca82, 32'hc3cb7a1b},
  {32'h45278662, 32'hc38bb4be, 32'h4471c21a},
  {32'hc5163606, 32'hc43b41c0, 32'hc4889388},
  {32'h44c1c265, 32'h43185fc3, 32'hc374463b},
  {32'hc47cd692, 32'hc47f0466, 32'hc4995bc6},
  {32'h43fe15e9, 32'h44353e07, 32'h44039265},
  {32'hc3f0452a, 32'h42e291af, 32'hc412e352},
  {32'h451baabe, 32'h441f06cc, 32'h43b41253},
  {32'hc311c770, 32'hc5014287, 32'h425a1b35},
  {32'h4331a37e, 32'h44b4e8df, 32'hc3118ab2},
  {32'hc47f3720, 32'h435a5afb, 32'hc3829007},
  {32'hc522fa7c, 32'hc3805dd2, 32'h440e5bfa},
  {32'h4490adf1, 32'h44ee9ae1, 32'h419c5ff0},
  {32'hc4051292, 32'hc3ed5638, 32'hc31794d9},
  {32'h432b7ecf, 32'h4523aedc, 32'hc38c5cd8},
  {32'hc4facc99, 32'hc48bdddf, 32'hc3aef648},
  {32'hc3c0c8dc, 32'h43256791, 32'hc2b4ea98},
  {32'hc4cde349, 32'hc420e30a, 32'h4156b2d0},
  {32'h44f3bbcb, 32'hc392f2f7, 32'h4474ff49},
  {32'hc38c4b5c, 32'hc49b2d41, 32'h4344f7f4},
  {32'h4461573b, 32'h44d83d8d, 32'hc2f6a67f},
  {32'hc3fc3fe0, 32'hc47b18e0, 32'h44aa0731},
  {32'hc386f3a5, 32'h448998a4, 32'hc4196701},
  {32'hc399de1a, 32'hc2a11ed8, 32'h44cdcfec},
  {32'h44830bef, 32'h451bf135, 32'hc32709fd},
  {32'h43b4ecea, 32'hc45494c6, 32'hc3facecd},
  {32'h43b484d8, 32'hc41560b2, 32'hc4da3cec},
  {32'hc4eed56c, 32'h427b710a, 32'h43e3249f},
  {32'hc3e4bbf0, 32'h43b09820, 32'hc4a102e8},
  {32'hc519e1f8, 32'hc35efe4b, 32'hc2ee395a},
  {32'h4319d1b0, 32'h44579191, 32'hc4b958e0},
  {32'hc3091aa8, 32'hc29048fd, 32'h4469a90b},
  {32'h4514da95, 32'h43cdf68a, 32'hc2f3c28e},
  {32'hc3df03b1, 32'hc3b5ffb1, 32'h4520753b},
  {32'h44709f7e, 32'h4231333e, 32'hc35daeea},
  {32'hc49985b7, 32'h43feeeb4, 32'h44d162d2},
  {32'h4514f2fc, 32'h432cd8db, 32'hc48e4cee},
  {32'h44817b8c, 32'hc4324d95, 32'hc485491c},
  {32'hc47f0f08, 32'h443338b8, 32'h40d0a860},
  {32'hc4ec5183, 32'hc35ce753, 32'h43be9a00},
  {32'hc5547c2b, 32'h44491480, 32'h431ad57e},
  {32'h44881bee, 32'hc4248bae, 32'h434d9a02},
  {32'h44deca70, 32'h43e6747f, 32'h4204ed31},
  {32'hc1515890, 32'hc3647d9e, 32'h434596a9},
  {32'hc58f08cc, 32'hc2cc5d67, 32'hc3bbff90},
  {32'h45292faa, 32'h434da49c, 32'h43dcbca5},
  {32'hc30f246a, 32'h44c520ba, 32'h43722e69},
  {32'h437d36cc, 32'hc457800d, 32'h44c40e4c},
  {32'h4444c76d, 32'hc30038a4, 32'h43672dd6},
  {32'h433dc158, 32'hc480c3db, 32'h44ad8ed5},
  {32'hc42243b4, 32'hc2eeb43f, 32'hc5511d45},
  {32'hbe60d300, 32'hc4c11265, 32'hc297af05},
  {32'hc3cd6184, 32'hc3b163f7, 32'hc53c4250},
  {32'h43c93d58, 32'h442092b8, 32'h45124c96},
  {32'h44f277b2, 32'h41978cc5, 32'h43391ad3},
  {32'h43cbbe05, 32'hc4b16ebe, 32'h447073f4},
  {32'hc529b372, 32'h442a1c59, 32'hc4051092},
  {32'h440a4067, 32'hc2e082e2, 32'h448be0b8},
  {32'hc3b6c144, 32'h444d3bef, 32'hc4c9c502},
  {32'h440780ff, 32'hc4ec5fce, 32'h440276ab},
  {32'h4321b3cf, 32'h4412e4de, 32'hc3917623},
  {32'h44f5a526, 32'h440ed1c0, 32'h4462ba9f},
  {32'hc582a7ca, 32'hc22583a9, 32'h430e939d},
  {32'h44c6f67a, 32'h43477e81, 32'h42ecd672},
  {32'h44258ad0, 32'hc32db150, 32'hc54060ee},
  {32'h443b1394, 32'hc42cf54a, 32'h44050ade},
  {32'hc4c6b29c, 32'h444784b2, 32'hc36caa91},
  {32'hc459b99d, 32'h433f9d93, 32'hc3910012},
  {32'h44f7597b, 32'hc3ba1bc0, 32'h4305517a},
  {32'hc32eb4b6, 32'h44ddd6d4, 32'hc3aa949c},
  {32'hc3ed1844, 32'hc3bdd004, 32'h43bbeeaf},
  {32'hc30234b7, 32'h4484a58f, 32'hc4ea34da},
  {32'h44beb99d, 32'hc285f7b3, 32'h4429b232},
  {32'h45258fd2, 32'hc3b9c956, 32'h4418b8ac},
  {32'h423d1db4, 32'h4496e6b3, 32'hc4ebad1d},
  {32'hc3b5061c, 32'h406048f0, 32'h436c2812},
  {32'h4284a648, 32'hc340d74f, 32'h448baaeb},
  {32'hc502a4d2, 32'hc042fd44, 32'hc34b2923},
  {32'h44642e9c, 32'hc0decb30, 32'h43f0a0e0},
  {32'hc4031962, 32'h43169837, 32'hc3a881ae},
  {32'h42a0c80f, 32'hc4b6b65b, 32'h4380a794},
  {32'h438fb8d7, 32'hc383c558, 32'hc566fb08},
  {32'h4486949b, 32'hc40fddd4, 32'hc26e67c6},
  {32'hc53ae83a, 32'hc3e29e17, 32'h43c5b863},
  {32'h456d3c93, 32'hc346722f, 32'hc4111af5},
  {32'hc463b341, 32'h424fae61, 32'hc31e4d59},
  {32'h4522558a, 32'hc33ed490, 32'h441c6622},
  {32'hc4310468, 32'h448a2d70, 32'h4374a4d6},
  {32'h44b3864e, 32'h43e47a0a, 32'h43400918},
  {32'hbf88e000, 32'h450d14a1, 32'hc3aea16e},
  {32'h44f2b26c, 32'hc3b741f2, 32'h44198c9e},
  {32'hc4b01d9e, 32'h43cf3971, 32'hc32ec575},
  {32'hc2c9bad2, 32'hc211703c, 32'hc4f5a7b4},
  {32'hc51387b5, 32'hc2e3ff0b, 32'h43dc4be3},
  {32'h41c9f310, 32'hc2e1bd17, 32'h44aecd8a},
  {32'h42011c00, 32'h43b67235, 32'hc497f54e},
  {32'hc4a0f618, 32'hc322e506, 32'h439e6cbc},
  {32'h448901d8, 32'h44ab0722, 32'h430d4d58},
  {32'hc4a23653, 32'hc432d38d, 32'h42cfdcbc},
  {32'h42a6cce8, 32'h44b14436, 32'h44078d87},
  {32'h43b47633, 32'hc30db51d, 32'hc41e53b3},
  {32'hc35a299f, 32'hc33fb611, 32'h4498d20f},
  {32'hc3c9f5c8, 32'h439fb9ee, 32'hc4ec31e7},
  {32'h4481069c, 32'h44869219, 32'hc3fd0e16},
  {32'hc432278a, 32'h4379f497, 32'h42edbddd},
  {32'h44864d6f, 32'h44399986, 32'h436a49ad},
  {32'hc36c6190, 32'hc52ea532, 32'hc3d3f865},
  {32'h4553456a, 32'h4289f4ab, 32'h405976a0},
  {32'hc248d790, 32'hc483f2e3, 32'h43c39365},
  {32'h444900b4, 32'hc43da84a, 32'hc43c6df6},
  {32'hc507fb4c, 32'h42cab02a, 32'h429edd62},
  {32'h45017d68, 32'h43d9869f, 32'h42bb794a},
  {32'hc4915c30, 32'hc49c02e9, 32'h42e6082a},
  {32'hc304dfe3, 32'h4554cb27, 32'hc292e3e4},
  {32'h43cd1f33, 32'hc50f3f56, 32'h42701c2c},
  {32'h450a06b8, 32'h43fc4c79, 32'hc3cfc02c},
  {32'hc5090f65, 32'hc46d8eaa, 32'hc2957c59},
  {32'hc483cfa0, 32'h4270d718, 32'hc18b525a},
  {32'hc3c32f4e, 32'hc226912f, 32'h42456130},
  {32'hc4b9f467, 32'hc451e46c, 32'hc02cfe7e},
  {32'hc0ed3140, 32'hc4b115bc, 32'h44a50323},
  {32'h4490f972, 32'hc4007c87, 32'h43ec7e63},
  {32'h453be9bf, 32'h4258b24b, 32'h43ff231b},
  {32'h437767f0, 32'hc2af46ff, 32'hc5073efa},
  {32'hc46d2a8b, 32'hc37946a1, 32'h43e4a178},
  {32'hc5889a97, 32'hc38dd44c, 32'hc33cdd74},
  {32'h44d69f5a, 32'h440bb64a, 32'h445cda8d},
  {32'h43d291d4, 32'h4499f96d, 32'hc319f287},
  {32'hc398ef3e, 32'hc4e76f8c, 32'h44fe4803},
  {32'hc3b72809, 32'hc4b84ee4, 32'hc42c9d64},
  {32'hc3ccda06, 32'hc08174ff, 32'h45023aee},
  {32'hc4a0d0f6, 32'hc4410a82, 32'hc3dd8568},
  {32'h444b31eb, 32'h451981ad, 32'h425031e0},
  {32'h44ed06e1, 32'hc3df9b87, 32'hc38bd9b6},
  {32'h43e39d04, 32'h431e7812, 32'h44aca0b9},
  {32'hc25b3a18, 32'hc37222ed, 32'hc56a401f},
  {32'h4511a4d4, 32'hc31ef1f8, 32'h4461163d},
  {32'hc56dae87, 32'h43781592, 32'h42a76ff6},
  {32'h44d8fcae, 32'h4484b599, 32'h43021cba},
  {32'hc3026068, 32'hc504e611, 32'h40f52764},
  {32'h44aa9c80, 32'h449b46d0, 32'hc34139d4},
  {32'hc3363698, 32'hc5335232, 32'hc3b858f0},
  {32'h443e3ddd, 32'h44026e90, 32'h43f3a863},
  {32'hc564eaec, 32'hc21185af, 32'hc3059111},
  {32'h4503cfb6, 32'h42c50969, 32'hc3595e63},
  {32'h44fdf7ae, 32'hc3d6064f, 32'h42575134},
  {32'hbfe40500, 32'hc3c136cf, 32'h450002e1},
  {32'h43262f41, 32'hc32f1609, 32'hc4054ff9},
  {32'hc4d943a8, 32'h44b79ca8, 32'h43e1d128},
  {32'h42c42472, 32'hc4259e6c, 32'hc470cfca},
  {32'hc4456403, 32'h43e03b43, 32'h441bbaa9},
  {32'h43287366, 32'hc50f83b9, 32'hc4d33dd3},
  {32'hc4b892e9, 32'h43831dbb, 32'h44c24fe3},
  {32'hc4cc64b2, 32'hc3d0d139, 32'h43a2a81b},
  {32'h448a2d21, 32'hc4a81ece, 32'h44b38011},
  {32'hc3dbca48, 32'hc4b4c36f, 32'hc4433a9c},
  {32'h42d88326, 32'hc4c0e2cd, 32'h43cdcb5e},
  {32'h44def43c, 32'h42ce708d, 32'hc3f21032},
  {32'hc516e26c, 32'h44488cf1, 32'h43213ad1},
  {32'hc4e3540b, 32'h42b461bb, 32'hc22b8d70},
  {32'hc5373b3c, 32'h424ba198, 32'h42c80226},
  {32'hc34eb2d2, 32'hc4c36255, 32'hc53abc21},
  {32'hc31a48e8, 32'hc322a5bc, 32'hc3b19a15},
  {32'h44b60f6d, 32'hc48ac7cc, 32'hc313d0f5},
  {32'hc55c40da, 32'h4364a729, 32'h41b3ca86},
  {32'h444c57ca, 32'h4336ef44, 32'hc364a587},
  {32'hc2bf8e14, 32'h45822e29, 32'hc198bacb},
  {32'h44e375e8, 32'hc4891494, 32'h434da44e},
  {32'hc51078ed, 32'h4381d298, 32'h433caf3f},
  {32'h456fef25, 32'h43b7830d, 32'h439ab832},
  {32'hc58dc548, 32'hc33256f8, 32'hc3b63cb1},
  {32'hc493cd4c, 32'hc38f8163, 32'hc2eec517},
  {32'h44580dc4, 32'h430050bb, 32'h44c1ddc2},
  {32'hc4a7fa43, 32'h426682c4, 32'hc488de23},
  {32'h45071275, 32'h4359557e, 32'h43009a1d},
  {32'h42901658, 32'h43dc3bc3, 32'hc3cb0301},
  {32'h453bb74a, 32'hc42fe5be, 32'h42bab6ab},
  {32'hc40c5fb8, 32'h449bfd08, 32'h43d4100e},
  {32'hc4c45a1c, 32'hc3b804df, 32'h4392ece7},
  {32'hc4f7e6b7, 32'h442f36cc, 32'hc388da66},
  {32'h43f67787, 32'hc4fa8059, 32'h433db0c2},
  {32'h450382a5, 32'hc3c9c86b, 32'h425e63ca},
  {32'h435c07ae, 32'hc3e73d01, 32'h4508185d},
  {32'hc3f87eb0, 32'hc183a108, 32'hbf93aee8},
  {32'h431d7019, 32'hc3c6e407, 32'hc426ba7e},
  {32'h43a54122, 32'h43da6d57, 32'h45336161},
  {32'hc04a7380, 32'hc52d00b6, 32'hc303bd42},
  {32'hc3ba823e, 32'h43d5b59d, 32'h44a6c477},
  {32'hc31a4700, 32'hc4f95b34, 32'hc2744444},
  {32'hc41a23b0, 32'h42e20361, 32'h43335a88},
  {32'hc480605a, 32'hc41ef7e6, 32'hc32dc41e},
  {32'hc480bb8e, 32'h4421211b, 32'h428cf92e},
  {32'h4511794f, 32'hc392d95f, 32'hc4531e51},
  {32'hc4c3b22f, 32'h42a2e76e, 32'hc3c06b75},
  {32'h43ff3376, 32'hc38c9715, 32'hc4eae346},
  {32'hc36af340, 32'h438f480f, 32'h4489d3cc},
  {32'h4315acae, 32'hc4903faf, 32'hc2827a55},
  {32'h43c5996f, 32'h44afec4e, 32'h44956f2c},
  {32'h45230950, 32'hc40793c0, 32'hc4664a7d},
  {32'h43880cc0, 32'h42360dd0, 32'hc491a4d8},
  {32'hc44793a9, 32'h4315fc61, 32'h44d21b1d},
  {32'hc28be138, 32'h44160a98, 32'h4036abe4},
  {32'hc3b1342c, 32'hc54727f2, 32'h429e9784},
  {32'h4420e11f, 32'h4447f295, 32'h43948069},
  {32'hc3b1421a, 32'hc304e2e6, 32'hc3d1ce14},
  {32'h45238ab3, 32'h440ecc98, 32'hc2b5a4f8},
  {32'hc49bbeae, 32'hc4d5802d, 32'hc3d21959},
  {32'h42c0e626, 32'h446b17c5, 32'hc252ca0f},
  {32'hc2b7ebb0, 32'h43c24ad1, 32'h44946ee8},
  {32'h42bed2c8, 32'hc0aaa0ad, 32'h441f198b},
  {32'hc428a0a6, 32'hc2c23f0c, 32'h43242e22},
  {32'h4466d33f, 32'h448a7baa, 32'h4401e335},
  {32'h4396ee7f, 32'hc4aefa48, 32'h43818a7a},
  {32'hc463013a, 32'h4447c1ab, 32'h4269cd29},
  {32'h42da5910, 32'hc469637e, 32'hc4503540},
  {32'h44bc6914, 32'h443b153d, 32'h445085f1},
  {32'h4451485a, 32'hc45c488e, 32'hc416eeaf},
  {32'h456a5a0e, 32'h41d1e1d6, 32'h415a8568},
  {32'hc48131c0, 32'h4466ecaa, 32'hc495e2f9},
  {32'h44aea322, 32'h44507d9f, 32'hc41a98ca},
  {32'hc3f8bb38, 32'hc4a122c1, 32'hc4188bbc},
  {32'h421f1f28, 32'hc2c6626a, 32'h4379eeac},
  {32'hc395c2bb, 32'hc4636d08, 32'hc3e6071f},
  {32'h437cddc8, 32'h443eedad, 32'h4484c808},
  {32'hc4668270, 32'hc410cba8, 32'hc439ffba},
  {32'h451d1d92, 32'hc38d4a0b, 32'hc4034516},
  {32'hc3f12252, 32'h43032de2, 32'h435b28a3},
  {32'h43ee589c, 32'hc5108a35, 32'hc397228b},
  {32'h44d1ec96, 32'h439cde72, 32'h44289da4},
  {32'hc52078b8, 32'h4427aa71, 32'h436a8727},
  {32'h43d343b0, 32'h45251416, 32'hc16286a0},
  {32'hc4ae9cd8, 32'hc40db49c, 32'hc247fca6},
  {32'h454d9f00, 32'hc319a165, 32'hc39b0c24},
  {32'hc53fefc8, 32'hc364158f, 32'hc2b9bc32},
  {32'h45180b1b, 32'h44100743, 32'hc20a484f},
  {32'h44a5b6aa, 32'h414cecb9, 32'hc38dd08d},
  {32'h44c82069, 32'h43654a96, 32'hc2d5e5c6},
  {32'hc507bb26, 32'hc36d2f9e, 32'hc3b7c824},
  {32'h43bde3f0, 32'h4414bd24, 32'hc3808b43},
  {32'h430fea58, 32'h42ab43db, 32'h4553d082},
  {32'h43da33b0, 32'h440a30b7, 32'hc3e2c763},
  {32'hc4c1368b, 32'h420466ec, 32'h43c90a0e},
  {32'h44bbe98f, 32'h43faf7c7, 32'h4386976b},
  {32'hc3ebb3c8, 32'hc3c84ad3, 32'h43916275},
  {32'h43f5df2a, 32'h43ab611d, 32'hc41bdee1},
  {32'hc3df14d0, 32'hc5316c23, 32'h42da9d48},
  {32'h45018861, 32'h448cba84, 32'hc446afe6},
  {32'hc3482118, 32'hc3d45ea4, 32'h44503607},
  {32'h4243587a, 32'h437d4276, 32'hc4f6e035},
  {32'hc2fa3bb2, 32'hc501fbe2, 32'hc1ee6e08},
  {32'h453d4a9a, 32'h417c0290, 32'hc1b9f1e4},
  {32'hc4eaa72e, 32'h43c2f647, 32'h44691485},
  {32'h449f9532, 32'hc3d3d8a0, 32'hc3c4ba65},
  {32'h45341bfc, 32'hc38150a7, 32'hc1b8d296},
  {32'hc4019c36, 32'h454499d1, 32'h438bbe8a},
  {32'h44af52ca, 32'hc3a60934, 32'h424d33ba},
  {32'h42b98b60, 32'h451051e0, 32'hc136b7d4},
  {32'hc37b6192, 32'hc4ef107f, 32'h43cb9297},
  {32'hc4a811be, 32'h43ca91f6, 32'hc3377c72},
  {32'h438b3fc0, 32'hc49c8b15, 32'hc4264e70},
  {32'hc5435ff2, 32'h43a152d5, 32'h435d32bc},
  {32'h44fb2cac, 32'hc36c3942, 32'h43f48773},
  {32'hc31bfbb1, 32'h44cb5a00, 32'h438e4d93},
  {32'h45235506, 32'h42b0be2c, 32'h43fce42b},
  {32'hc441677e, 32'h442fe7c8, 32'hc35925f6},
  {32'hc338b722, 32'hc5564825, 32'h43c7ed0f},
  {32'hc3c8014f, 32'h438f58f0, 32'hc536eb81},
  {32'hc4cd2d15, 32'h43857fdb, 32'h43989a1a},
  {32'hc2ec10ac, 32'hc3ca86ca, 32'hc569f8f3},
  {32'h45022a14, 32'hc303502f, 32'h437fa03d},
  {32'hc498eba4, 32'h431ccb0d, 32'hc4551f7c},
  {32'h44c478e5, 32'hc496d7a6, 32'h4086739f},
  {32'hc4d737c6, 32'h44809a9b, 32'hc355c7f6},
  {32'hc3e96036, 32'hc4840529, 32'h43a40516},
  {32'hc30e8060, 32'h44ca253b, 32'hc489df4c},
  {32'h43d058e9, 32'hc42e15a4, 32'h4442fa7e},
  {32'h4401ff5e, 32'h44046a6a, 32'hc42a2d1d},
  {32'h42bb47e8, 32'h4489b8ae, 32'h45437f4d},
  {32'hc5171175, 32'hc411789c, 32'h41171055},
  {32'h45599417, 32'hc3123071, 32'hc40a9440},
  {32'hc497e3b0, 32'h43f9fab9, 32'hc46d86be},
  {32'h42b90e1c, 32'h43f6dfa7, 32'h44a54a4d},
  {32'h4431001c, 32'hc3a3ab26, 32'hc40a5fb6},
  {32'h441c6b8a, 32'h4295e24f, 32'hc3a62561},
  {32'h44ee503c, 32'hc20dac06, 32'h4407e0b2},
  {32'hc517f4de, 32'hc258811a, 32'hc3f681e8},
  {32'h44d87993, 32'h4206fd2b, 32'h43b110fe},
  {32'hc3ae51f2, 32'h446b6157, 32'hc418228f},
  {32'h44956643, 32'hc43e0e43, 32'h4480a9ca},
  {32'h44b7c0de, 32'h44ab241a, 32'h4499c42b},
  {32'hc48a12e4, 32'h4279c944, 32'hc50e08b5},
  {32'hc388968b, 32'hc383bd32, 32'h44c864b5},
  {32'hc2c99bb4, 32'h42cc12b2, 32'h447f1314},
  {32'h43f3e5a4, 32'h4482ed74, 32'h4395c79a},
  {32'h452cfade, 32'h43885471, 32'hc321622c},
  {32'h41c91d80, 32'h43218441, 32'hc4ebb035},
  {32'h4466f9e6, 32'hc3f348aa, 32'h44affce5},
  {32'hc4c653c2, 32'h4348a9ce, 32'hc419d125},
  {32'h4355df2b, 32'hc3f8b0fa, 32'h42ba9a76},
  {32'hc53bdd5a, 32'h42d13a8e, 32'hc22e3ad5},
  {32'h4250ed40, 32'hc3309b35, 32'hc38512ba},
  {32'h44f53c12, 32'hc13ce51d, 32'hc26db461},
  {32'h455a8fb3, 32'h42bc0283, 32'h433e575e},
  {32'hc4889414, 32'h4382ddeb, 32'hc3a949c9},
  {32'h44fc6386, 32'h43a9ea1a, 32'h43ecc87a},
  {32'hc4c47044, 32'h449def48, 32'h436ba51c},
  {32'h43950aba, 32'hc4975936, 32'h43ad8477},
  {32'h4391e208, 32'hc3c5a106, 32'h4463d7b9},
  {32'hc4601345, 32'hc29a7bd0, 32'hc494611b},
  {32'h43fb1fc3, 32'hc4acf6a2, 32'h44c221aa},
  {32'hc3da6f89, 32'h43bda9c1, 32'h44fc033e},
  {32'h424e9200, 32'h454072b2, 32'h43965843},
  {32'hc33ad683, 32'h4351f881, 32'h4496d69d},
  {32'h450604b8, 32'h43b77309, 32'hc3fa543b},
  {32'hc49a9bdc, 32'hc4587981, 32'hbed0684e},
  {32'h44a90b8f, 32'hc3ac2f01, 32'hc41bce33},
  {32'h4478d25b, 32'h420c03dc, 32'hc30b6824},
  {32'h44134f2f, 32'hc45ebc01, 32'h451ac74a},
  {32'hc3393c0d, 32'hc48fda41, 32'hc4e76a14},
  {32'h43c66ca2, 32'h43142bdf, 32'hc4c79ef6},
  {32'hc4846800, 32'hc3bdd91f, 32'h448eb5a5},
  {32'h442e995c, 32'h4493dc4b, 32'hc38668ff},
  {32'hc48fefa6, 32'hc3c75c84, 32'h4471bd82},
  {32'h439087cc, 32'h44a0f964, 32'hc40091b1},
  {32'hc3ee597f, 32'hc420551d, 32'h43f1f99f},
  {32'h45218878, 32'hc3923fbd, 32'hc120b689},
  {32'hc53bfbc2, 32'h4380d377, 32'hc332fe0f},
  {32'h4552f647, 32'h43d1689a, 32'hc2e31d18},
  {32'hc518f513, 32'hc45ff0cd, 32'h421028b2},
  {32'h4465b9a0, 32'h43cd4ea1, 32'h431bd244},
  {32'hc52b4641, 32'h4363b0ca, 32'hc2bc05a9},
  {32'hc2eae680, 32'h4535e93f, 32'h433ff3dc},
  {32'hc520571a, 32'hc41e8db3, 32'h43584e39},
  {32'hc4b93e04, 32'h43b69679, 32'h43b65db6},
  {32'hc46d20b6, 32'h4227d61d, 32'h421f9f1b},
  {32'h441cca74, 32'h45055583, 32'hc492ef9d},
  {32'hc35add40, 32'hc44e512a, 32'h44a81422},
  {32'hc4c4243e, 32'hc2191fe5, 32'hc3357b88},
  {32'h43aabda8, 32'h4240569a, 32'h4518d257},
  {32'hc50c0bd6, 32'hc3bc7df7, 32'hc438a932},
  {32'hc42612d2, 32'hc35d5b71, 32'h439e34da},
  {32'hc44d595e, 32'hc3b15da2, 32'hc50ce124},
  {32'h43aa2b0c, 32'h446e70e1, 32'h44923d82},
  {32'h434074b8, 32'h430f364a, 32'hc39a7dce},
  {32'hc33b0ff0, 32'hc317213a, 32'h4497400e},
  {32'hc397b4fd, 32'h44291d0a, 32'hc4a05fcb},
  {32'hc475bf6c, 32'hc20b065a, 32'h440342e7},
  {32'hc2a18b98, 32'hc51a3313, 32'hc451cfd7},
  {32'h44221408, 32'h44900ec5, 32'h4303a293},
  {32'h412ca120, 32'hc282cf0e, 32'hc4b06ab2},
  {32'h45601a13, 32'h43830b79, 32'hc388c531},
  {32'hc338dd28, 32'hc472fad2, 32'hc537f7d8},
  {32'h4406f2dc, 32'hc32a6b83, 32'h4391a3b2},
  {32'hc53e57c7, 32'h42bb2c30, 32'hc32095e3},
  {32'hc36f9560, 32'h44ed7d60, 32'h446a6f17},
  {32'hc495a787, 32'h432f4715, 32'hc4498dc2},
  {32'h433e1310, 32'h451a0abc, 32'hc3337911},
  {32'hc3a3cc14, 32'hc57baacf, 32'h4264e5da},
  {32'hc42ffad2, 32'h437a7894, 32'hc229a11b},
  {32'hc3f37a26, 32'hc39a3650, 32'h437df7ad},
  {32'h45488177, 32'hc0d41467, 32'hc0980634},
  {32'hc4a73076, 32'h4451dc10, 32'hc4f9a063},
  {32'hc3eaaad6, 32'h43049a2a, 32'h44a6b0d5},
  {32'h42df7d74, 32'hc3fda759, 32'h4272a1b2},
  {32'hc49230d6, 32'h439ec3a9, 32'h44b00d67},
  {32'hc418e07f, 32'hc530514b, 32'hc3aed6e6},
  {32'hc44d298c, 32'h440cda44, 32'h43ea657e},
  {32'h4478f1aa, 32'hc37bf95b, 32'hc48bd5c9},
  {32'hc4a5bead, 32'h430ca42f, 32'h44cbbec0},
  {32'hc466b91b, 32'hc3960de5, 32'hc44855a6},
  {32'h439d0ebc, 32'h44581cc6, 32'h449db9ca},
  {32'hc4313616, 32'h44c83b6c, 32'hc506ef48},
  {32'h437dafa3, 32'h44a34661, 32'h42bec236},
  {32'hc3e144ed, 32'hc3f7d8de, 32'hc5256198},
  {32'hc3fd59ad, 32'h4499064d, 32'h435a9466},
  {32'hc4c5ec48, 32'hc20422f0, 32'h418109b8},
  {32'hc3e70c60, 32'h448c5c14, 32'h44b662e1},
  {32'h43805b8e, 32'hc4a74707, 32'hc522be3e},
  {32'h43ceb158, 32'h447ea072, 32'h44d9ba3f},
  {32'h449c9338, 32'hc5098637, 32'hc2bb1478},
  {32'hc0f7967a, 32'h45556009, 32'hc31f20a5},
  {32'hc48972b4, 32'hc2e7afe7, 32'hc34c9e23},
  {32'hc256ab50, 32'h45290f5f, 32'hc312e724},
  {32'h43351390, 32'hc2d66c7e, 32'h4301d4eb},
  {32'h44c10c23, 32'h43e74feb, 32'hc367471c},
  {32'h44c3293e, 32'h439daef4, 32'h416882de},
  {32'hc4bd99e3, 32'hc44e63f9, 32'h43dd3f9c},
  {32'hc2dda570, 32'hc39880f3, 32'hc2b5f29e},
  {32'h44eb1bc7, 32'hc389ba02, 32'hc3874d1b},
  {32'hc4124bcd, 32'h4423e579, 32'hc4e25946},
  {32'h45094d9b, 32'h42c18e07, 32'h4422bf06},
  {32'hc4b60c03, 32'h4330fb39, 32'hc3e1e7af},
  {32'h4525747f, 32'hc4024d41, 32'h4307b0cc},
  {32'h4291dd90, 32'h4555f509, 32'hc1c7cba0},
  {32'h44a0c96e, 32'hc29290b4, 32'hc195c22f},
  {32'hc4e7f1c9, 32'h44072b84, 32'hc32ab2fc},
  {32'h44419464, 32'hc4e6c686, 32'hc31a07e4},
  {32'hc3d11912, 32'hc3271238, 32'hc31c0977},
  {32'h443d8287, 32'h41502061, 32'h44c06f7e},
  {32'hc41c7e9c, 32'h445fa038, 32'h43ac30f9},
  {32'h451cf886, 32'h43a1faff, 32'h43adc92a},
  {32'hc41413dd, 32'h4331e04d, 32'h43be931c},
  {32'h442484ad, 32'hc4204d96, 32'hc4023122},
  {32'h44705e90, 32'h43fe319b, 32'h4206814f},
  {32'h43d46bba, 32'hc47d8661, 32'hc472f005},
  {32'hc538d2b7, 32'hc3e2240b, 32'h418515b3},
  {32'hc4209098, 32'h4333e150, 32'hc4056561},
  {32'hc4ea3710, 32'hc44250db, 32'hc28f7a8c},
  {32'h4508b404, 32'hc407360b, 32'hc47e82fc},
  {32'hc49ae680, 32'h3fc0bf7c, 32'hc2cecbd1},
  {32'h43c0f548, 32'hc469ac09, 32'hc4a61ebf},
  {32'hc41068e5, 32'h4507ad27, 32'h43306a1f},
  {32'h41213580, 32'hc2f8b8e9, 32'hc497dc43},
  {32'hc4f8391b, 32'h43d2131e, 32'h441493ec},
  {32'h438d803c, 32'hc511ca75, 32'hc3bfdfe5},
  {32'h41839780, 32'hc35a20e2, 32'hc4aab678},
  {32'hc537e7ea, 32'h43413c95, 32'h443cdeba},
  {32'hc47e807e, 32'h440cdc7c, 32'h43a400ed},
  {32'hc4b5c3d4, 32'hc460c0d7, 32'hc376afbf},
  {32'h44fd0c40, 32'h43a0b922, 32'h433f8457},
  {32'h4447e7a9, 32'hc49e1c28, 32'hc3de3999},
  {32'hc3090030, 32'h44e172fa, 32'hc37671f2},
  {32'hc4eec6ba, 32'hc48c81b0, 32'hc40c0379},
  {32'hc4c47711, 32'hc36e7582, 32'h4404cca6},
  {32'hc32e33eb, 32'h43e8e9cd, 32'hc4b7cb64},
  {32'h43d39fc2, 32'hc4182e20, 32'h442b1fab},
  {32'h43f023ea, 32'h42ad9e5f, 32'h44654cae},
  {32'h436cda00, 32'h44a8e331, 32'h4484bcf8},
  {32'hc51ddf3e, 32'hc32fbb22, 32'h42191f7d},
  {32'h44dced37, 32'hc40d119f, 32'hc2f8abf5},
  {32'hc3a908bd, 32'hc1711864, 32'hc5507de3},
  {32'hc3447f9a, 32'h44d268f0, 32'h438db356},
  {32'h448deff1, 32'hc3ad1dd0, 32'hc42934de},
  {32'h430f518c, 32'h4418164c, 32'h44b54997},
  {32'hc33a7cdc, 32'h442cd570, 32'hc4a1d7c9},
  {32'h437a2600, 32'hc3beb727, 32'hc32f8c27},
  {32'h4392dc33, 32'hc55a5fdf, 32'hc41811eb},
  {32'h439f202c, 32'h4483b6a4, 32'h44168941},
  {32'hc3c40f2a, 32'hc3840dbd, 32'hc4a211e8},
  {32'hc3b2825c, 32'h4324200c, 32'h452bceb8},
  {32'hc4a65bbc, 32'hc44c7dad, 32'hc42443a9},
  {32'h44e0c963, 32'hc3b86d80, 32'hc33e4ed6},
  {32'hc332c07e, 32'h44d68908, 32'h44022cee},
  {32'hc49ba15c, 32'hc40cd21e, 32'hc446bc0c},
  {32'hc2a171c0, 32'h44647cd9, 32'h44610c4a},
  {32'hc4d17b28, 32'hc38d3e8c, 32'h43761095},
  {32'h44c4a90e, 32'h449d4a3b, 32'hc3510876},
  {32'hc3f9e261, 32'hc55367e0, 32'h43d0b2cb},
  {32'hc4aacaca, 32'h43f34646, 32'h436ce0ab},
  {32'hc54bfb9b, 32'hc24038dc, 32'hc1ba4685},
  {32'h44eac5a5, 32'hc206af83, 32'h446e9e8f},
  {32'hc50cba0e, 32'h43ea0062, 32'h43e33996},
  {32'h4354a61e, 32'h43191042, 32'hc3f5db81},
  {32'hc1db5140, 32'hc4fbe33c, 32'h4299577a},
  {32'h43ee43d2, 32'h44bac68f, 32'h4392dfb9},
  {32'hc46e0b37, 32'h42ac114e, 32'h447fb2b6},
  {32'h43e697ac, 32'h440d7d6a, 32'hc4805add},
  {32'hc506b17e, 32'h437094cc, 32'h43d18ecd},
  {32'h4525887a, 32'h43996180, 32'hc3b06309},
  {32'hc40c7f8d, 32'hc3539b2f, 32'h4443833c},
  {32'h43654e8a, 32'h43b8d0da, 32'hc410ffe1},
  {32'hc569a292, 32'hc2e276a7, 32'hc208e480},
  {32'h446fb474, 32'h44554293, 32'hc47f5ab0},
  {32'hc38e59e4, 32'hc1a48b08, 32'h441b17bd},
  {32'hc1e84000, 32'h449befd3, 32'hc40012dc},
  {32'h4381e482, 32'hc53f6a22, 32'h427a185b},
  {32'hc42ff06a, 32'hc36a0d43, 32'hc43943b0},
  {32'hc545e718, 32'hc3c17e6b, 32'h438d079e},
  {32'h44997cb6, 32'h436a90de, 32'hc4e72a16},
  {32'h44c4db69, 32'hc4eee1b0, 32'hc3a2d26f},
  {32'h427f4ec0, 32'h4529a638, 32'h4161b43c},
  {32'h452f1992, 32'h44217ed2, 32'h433aa364},
  {32'h43182dc9, 32'h453459b5, 32'hc3dff0ec},
  {32'h440d916d, 32'hc50f5932, 32'h425b96d0},
  {32'h44c46a02, 32'h42d85d71, 32'h424e2417},
  {32'h44e971dc, 32'h434daf0f, 32'h4380bc0f},
  {32'hc57f9a7c, 32'h4428dae3, 32'hc3c179c1},
  {32'h451ebb90, 32'hc3743db6, 32'h4408a76f},
  {32'hc45aa690, 32'h43c125c5, 32'hc472f95a},
  {32'h44b7b92c, 32'h438576c4, 32'hc38f127a},
  {32'h42f11580, 32'h4443e3ec, 32'h43a41360},
  {32'h441a2ca4, 32'hc35929b6, 32'h4450708b},
  {32'hc3eeb900, 32'h444adac6, 32'hc4857f70},
  {32'h436c3be2, 32'hc4bfae7a, 32'hc08c0e10},
  {32'hc51a5702, 32'h4414c4ec, 32'hc324c36f},
  {32'h442d9336, 32'h438a5004, 32'h44cbf82b},
  {32'h449bf89f, 32'hc3e2fba1, 32'hc46bf435},
  {32'h44aa58bf, 32'hc4db7373, 32'hc3805120},
  {32'hc4dd5436, 32'h446684d9, 32'hc446ef6f},
  {32'h43c96139, 32'hc336d155, 32'h42cc82d9},
  {32'hc3b569a2, 32'h441d872e, 32'hc5023154},
  {32'h4488aca8, 32'hc3183758, 32'h44a91070},
  {32'h43b381b4, 32'hc38eeafa, 32'hc485f775},
  {32'h440fee67, 32'h43eb112f, 32'h4519f78b},
  {32'hc563ab12, 32'hc3843508, 32'hc395c794},
  {32'hc405d0c4, 32'h44018f42, 32'h4483b522},
  {32'hc424f291, 32'h44896523, 32'hc4bf274f},
  {32'h447ef1b9, 32'h4428932e, 32'h448472be},
  {32'h43214d3e, 32'hc3ff2a94, 32'hc4b3fcc4},
  {32'hc37e7288, 32'h3ef95e00, 32'hc4840620},
  {32'h43457350, 32'hc4aca945, 32'h447e8687},
  {32'h43a1f448, 32'hc3b226df, 32'hc536eaa4},
  {32'hc2355439, 32'hc1a05e45, 32'h44c2a13b},
  {32'h42ffeef6, 32'h432ad961, 32'hc4cf2cdf},
  {32'h433fcfc4, 32'hc49bbe72, 32'hc22fd852},
  {32'h4300e9b0, 32'hc42887e6, 32'h4514b2e1},
  {32'h41b559e8, 32'hc3438663, 32'hc50a1078},
  {32'h4276afc0, 32'h447f7aca, 32'h4425b0ec},
  {32'hc3038b60, 32'hc2a56a6a, 32'h4318c6fe},
  {32'h420daed0, 32'h45233094, 32'hc3510172},
  {32'h44d04a0b, 32'hc40c938c, 32'h43d43f2e},
  {32'h43ad5b08, 32'h43a6352e, 32'h43809ae7},
  {32'h43da60fd, 32'hc4dfe8d3, 32'h430bc5ce},
  {32'hc428736e, 32'h431a2122, 32'hc4047215},
  {32'h4563f4b4, 32'hc3af9d86, 32'h441e63ec},
  {32'hc5358003, 32'hc39e416c, 32'hc4092134},
  {32'h44169785, 32'h442f5df9, 32'h4487117e},
  {32'hc437ea68, 32'hc1ab6dad, 32'h43401059},
  {32'h417acf7c, 32'hc4a59670, 32'h44389477},
  {32'hc4af8cd7, 32'h44319168, 32'hc34a63b4},
  {32'h4553bf50, 32'h43643a19, 32'h439d84af},
  {32'hc2e655af, 32'h457b7461, 32'h42aa9fc7},
  {32'h448920b3, 32'hc50903e7, 32'hc2af2492},
  {32'hc2888a28, 32'h44af7ed4, 32'hc29ed2a5},
  {32'h44064211, 32'h43c879fe, 32'hc46b795a},
  {32'hc37e3890, 32'h4487e1ac, 32'h44831d7b},
  {32'hc431b736, 32'hc4545fd3, 32'h438c9f3e},
  {32'h44744026, 32'h43f02b64, 32'hc3aa33b8},
  {32'h4479f951, 32'hc3f9b54d, 32'h43d53c1d},
  {32'h42f9d7ae, 32'h44a043ab, 32'hc4976c35},
  {32'hc4b24683, 32'hc440fb3b, 32'hc22ad967},
  {32'hc3186eb8, 32'h4499ed91, 32'hc3f33ddb},
  {32'hc39f3546, 32'hc45a4b7c, 32'hc322a12c},
  {32'h41262f80, 32'h4430503b, 32'h449548f0},
  {32'h42aa0f25, 32'hc3bda689, 32'hc4e1e96f},
  {32'h44959386, 32'h445b5145, 32'hc406c3f5},
  {32'hc3df557d, 32'hc3ade199, 32'h4535f3ec},
  {32'h4355a6b2, 32'h428bb14b, 32'hc49e7595},
  {32'hc43235fa, 32'hc2e17ef4, 32'h449d24e4},
  {32'hc34d448f, 32'hc2fa7b38, 32'hc54b23a5},
  {32'h44ff3ea6, 32'hc32f8856, 32'hc2995aa1},
  {32'h4572922e, 32'hc32dc1b2, 32'h441a7bef},
  {32'hc4f6e186, 32'h43db1230, 32'hc39331f5},
  {32'h43a998ce, 32'hc1a7824c, 32'h43047ec2},
  {32'hc28f1577, 32'hc4d12ed4, 32'hc3600a30},
  {32'h446a7984, 32'h44c10dce, 32'hc325ba04},
  {32'h4419af28, 32'hc4070bab, 32'hc1e7f7b9},
  {32'hc2e9964e, 32'h453985e2, 32'h4284c4d5},
  {32'hc58ab949, 32'hc30ea83a, 32'hc3591ce8},
  {32'hc367141e, 32'h44850b39, 32'hc40ff83d},
  {32'hc2a65bc8, 32'hc3cc2176, 32'hbfe454ac},
  {32'hc4334f02, 32'hc338e6d4, 32'hc41025fc},
  {32'hc22b3200, 32'h429ba8a5, 32'h43c54c48},
  {32'h447edf2c, 32'h42cbb730, 32'hc44cc85f},
  {32'h430cec5b, 32'h448e0f98, 32'h43fe8796},
  {32'hc3a34cfc, 32'hc5190060, 32'hc4028a80},
  {32'h4505add5, 32'hc3091696, 32'hc30ddf53},
  {32'hc50b756c, 32'hc4a2da7c, 32'hc47f80ba},
  {32'h438e506c, 32'h447b35cd, 32'h44b3a7e4},
  {32'h43be088b, 32'hc38c7d76, 32'hc461d355},
  {32'h4396895f, 32'h4531c805, 32'h4206f6cd},
  {32'h439487a4, 32'h439b5920, 32'hc3a62561},
  {32'h434620f4, 32'h4491c053, 32'h42d11928},
  {32'hc4056e4a, 32'hc31832d4, 32'hc47c6e85},
  {32'h441a8850, 32'h4531e0eb, 32'h424009e7},
  {32'hc4030454, 32'hc41f5764, 32'h437c8f25},
  {32'h43f943c8, 32'hc3174e50, 32'h44b788b9},
  {32'hc511f3d0, 32'hc2c1e9f9, 32'hc3bac809},
  {32'hc3a44eac, 32'h41c72360, 32'h43f00899},
  {32'hc4a86192, 32'hc4c926a4, 32'hc3218f30},
  {32'h43b53091, 32'h451a8d35, 32'hc275e978},
  {32'h43aa245c, 32'hc4c9e203, 32'hc3bf8762},
  {32'h43b58e38, 32'hc3164fd2, 32'hc232dd23},
  {32'hc4e0ce92, 32'hc3512709, 32'h427a83b9},
  {32'hc4208cf1, 32'h43150eae, 32'h4325ec25},
  {32'hc505923d, 32'h44148372, 32'h4405ed9d},
  {32'h45067b9a, 32'hc41d9055, 32'h443483ba},
  {32'hc1bfd9aa, 32'hc51a8c4f, 32'hc3edea2e},
  {32'hc484c01c, 32'h43bd31cc, 32'hc3946fb3},
  {32'hc3c57cf4, 32'h43393ad2, 32'hc3996655},
  {32'hc3f0c8c7, 32'h44a67b6f, 32'h42faff2e},
  {32'hc34644bd, 32'hc481d577, 32'hc4ae2f25},
  {32'h4385722d, 32'h4511d1e5, 32'h43913475},
  {32'hc1aba960, 32'hc433afc7, 32'hc5222901},
  {32'hc45a1c01, 32'h442927da, 32'h44ac447b},
  {32'hc44003f6, 32'h42d511c1, 32'hc4ba13f5},
  {32'hc48bdb88, 32'hc2ed9251, 32'h444e623d},
  {32'h4451f99e, 32'h4486d080, 32'hc459ea26},
  {32'h439b2d86, 32'h430a3c2a, 32'h443304e7},
  {32'h447682ff, 32'hc3702aad, 32'hc422248e},
  {32'hc48388b9, 32'h45086413, 32'h42757bae},
  {32'h4342ead3, 32'hc39b5952, 32'hc4c0d734},
  {32'hc37db83a, 32'h45005f90, 32'h44d3c69f},
  {32'h4400b7f4, 32'hc44d4822, 32'hc444a31f},
  {32'h43e1e5b6, 32'hc31aa492, 32'h442e95bf},
  {32'h44b3968d, 32'hc463193d, 32'hc2357c82},
  {32'hc4956bc0, 32'h4464bd9a, 32'h43ce2206},
  {32'hc459efe3, 32'hc394a666, 32'h411fe646},
  {32'hc33bd4d0, 32'h455a4b34, 32'hc15c6dd8},
  {32'h44b679c5, 32'hc45d9a3f, 32'h42c1a68f},
  {32'h44b21055, 32'h436b1f92, 32'h42c8e2d5},
  {32'h456ddb3c, 32'h42f133d9, 32'h428dada2},
  {32'hc58c4c1b, 32'hc30397c5, 32'hc36bfe3a},
  {32'hc31eb1f2, 32'hc3f5537c, 32'h43d633bb},
  {32'h445e43a1, 32'hc3a33b8f, 32'h449e59d1},
  {32'hc4df3472, 32'h44490031, 32'hc4517ead},
  {32'h44a6d5ef, 32'hc1a9f694, 32'h44e08ea5},
  {32'h4420849b, 32'h44b2df91, 32'h42b8a3bd},
  {32'h43e0bd30, 32'hc3c6c5a2, 32'hc4089a3b},
  {32'hc3d9c6c7, 32'h44906bec, 32'hc3ad948e},
  {32'hc3d6136e, 32'h418b6141, 32'hc1936c26},
  {32'hc4f0212e, 32'h43f4a37b, 32'hc33027d3},
  {32'h442098e2, 32'hc49ce19b, 32'hc312c906},
  {32'h43dd89f8, 32'h4327bd40, 32'hc48c1ebe},
  {32'h45060d97, 32'h428ee503, 32'h43948296},
  {32'h41ed767c, 32'h4367b165, 32'hc4484d36},
  {32'h4401ed0f, 32'hc28be806, 32'hc4bcb03e},
  {32'h435a7b78, 32'hc1fc84a8, 32'h4516df81},
  {32'h4450a1f0, 32'hc444dab2, 32'hc3ff368e},
  {32'hc49e97fe, 32'h442e7b50, 32'hc109fe33},
  {32'h449e0411, 32'h438f5927, 32'hc4aed9b7},
  {32'h429659c2, 32'h451a1c59, 32'hc394dd75},
  {32'h454e8d74, 32'h43cf7013, 32'h43ef482f},
  {32'hc5450e96, 32'hc468fad7, 32'h441f700b},
  {32'h4540f87b, 32'h42b66fb4, 32'hc3ec5cef},
  {32'hc4b20a72, 32'h434f7c58, 32'hc38721d2},
  {32'hc405b522, 32'h43832d8e, 32'hc535f208},
  {32'hc2c8ea40, 32'h42b21fbd, 32'h43f13552},
  {32'h43a2bd38, 32'hc4d1ef2d, 32'hc1941bad},
  {32'hc37bc26b, 32'h452476b1, 32'hc312d2f2},
  {32'hc35d6486, 32'hc541c1f9, 32'h4319f1f9},
  {32'h43976ec0, 32'hc42a78a3, 32'h425fe86a},
  {32'hc428ff5a, 32'hc2dd5cfe, 32'h450d8853},
  {32'hc4490baf, 32'h4364557b, 32'h43ef1a27},
  {32'hc3b082b8, 32'hc520c99e, 32'hc42e9e7f},
  {32'h42d28a2e, 32'h44f217a3, 32'h444818c3},
  {32'h4496d796, 32'hc43d8783, 32'hc36e31a4},
  {32'h44e59a9a, 32'h44be09de, 32'h4171e60a},
  {32'hc4706948, 32'hc4a84ca5, 32'h43d70fbf},
  {32'h44692bf0, 32'hc31b6a26, 32'h44116407},
  {32'hc48b2bc8, 32'h4384dd99, 32'hc48c64c8},
  {32'h4426c3e2, 32'hc41e2666, 32'hc4fd1ea4},
  {32'hc469d2dc, 32'hc40305f1, 32'hc41d09b7},
  {32'h42e5e0a0, 32'hc33ffc43, 32'h4552d688},
  {32'hc4065df3, 32'hc4164fc4, 32'hc4221c39},
  {32'h4451e026, 32'h43409375, 32'h440ea381},
  {32'h4309d17a, 32'hc4fe778d, 32'h430da654},
  {32'h44d0846d, 32'h438b6d05, 32'h42492c75},
  {32'hc3665c60, 32'hc4ac3b78, 32'hc3d082c2},
  {32'hc38ed5b2, 32'hc3532617, 32'h43a804b7},
  {32'hc4bc7e16, 32'hc447f3e9, 32'hc39c3be2},
  {32'h44353a7c, 32'h44153e70, 32'hc3e60247},
  {32'hc4a5e935, 32'hc44750a7, 32'hc43b6e35},
  {32'h44432a96, 32'h44333254, 32'h439331f7},
  {32'h43a30a0a, 32'hc4816f26, 32'hc16d66ed},
  {32'hc2cf37e1, 32'h453572f6, 32'h40bcf860},
  {32'hc4b64d9b, 32'hc49b24fc, 32'hc48940a0},
  {32'hc372d42d, 32'hc3377000, 32'h4461be63},
  {32'hc4b8c4d6, 32'hc1fc1630, 32'h43346479},
  {32'hc4d5ca25, 32'hc24cf577, 32'h439e1b52},
  {32'h43a09640, 32'h44f5e838, 32'hc2aa0524},
  {32'h42fd26f8, 32'hc43a4652, 32'h43f932bb},
  {32'h44b71671, 32'h448ef640, 32'hc2b209fa},
  {32'hc4351c04, 32'hc42e5805, 32'hc304c2b8},
  {32'hc4d7e2c4, 32'hc2be8908, 32'h42663fb5},
  {32'hc5122c92, 32'hc45ff9a2, 32'hc43efbdd},
  {32'h4480ac64, 32'h4448ee72, 32'h443211e1},
  {32'h43b82481, 32'hc4953d97, 32'hc1b5decc},
  {32'h44bdbd9d, 32'hc34be6a0, 32'h4442ffb4},
  {32'hc48c3fdf, 32'hc3bf8b6a, 32'h42fe384e},
  {32'hc486116a, 32'h43846182, 32'hc3559940},
  {32'hc4609e27, 32'hc470999e, 32'h42272789},
  {32'h43627d22, 32'hc3dd731c, 32'h421b34c8},
  {32'hc12ac428, 32'h42ae57f4, 32'h448404be},
  {32'h4303cbc8, 32'h41d44025, 32'hc4f62ae0},
  {32'hc5108d5d, 32'h425e3284, 32'hc36a0ee9},
  {32'h453c031c, 32'hc446e578, 32'hc2e4d7e8},
  {32'hc46db27e, 32'hc48c04d9, 32'h426ba5a1},
  {32'h4309484a, 32'h4526e1b3, 32'hc3c14780},
  {32'hc4ed8fb4, 32'hc3093414, 32'hc3ebc671},
  {32'hc3bd1377, 32'h43c565b0, 32'hc448e37e},
  {32'hc4a7e3ef, 32'h43467b48, 32'h4427f2e0},
  {32'hc09d648c, 32'hc39d1abc, 32'hc4d5c398},
  {32'hc3156108, 32'h43f4bd00, 32'h45263295},
  {32'h43907328, 32'hc3bf2fa6, 32'hc52fc235},
  {32'h445fdb78, 32'h4386b686, 32'hc488bf7e},
  {32'hc4c25440, 32'h4463e123, 32'hc18af417},
  {32'h43ee0812, 32'hc45f8c57, 32'h433a2e3b},
  {32'hc500eb5e, 32'h446bc677, 32'h43fb528c},
  {32'h454c3caa, 32'hc329a8b9, 32'hc3d5d218},
  {32'hc43a3f2e, 32'hc3845848, 32'hc2d3e382},
  {32'h45346c7c, 32'hc44a978b, 32'hc41f7beb},
  {32'hc5873d8f, 32'h43d6a4a8, 32'h43d72bf7},
  {32'h456e3e06, 32'h42d0306b, 32'h4334d312},
  {32'h438e351c, 32'h443b24a3, 32'hc41950e4},
  {32'h43bb128b, 32'hc41a7460, 32'h45138a39},
  {32'hc4ed4b9a, 32'h42691aeb, 32'hc346eb5e},
  {32'h44ae9485, 32'hc3fd5c1b, 32'h43ca6ba1},
  {32'hc5030494, 32'h4338488d, 32'hc331ea7c},
  {32'h4266502c, 32'hbe45e5c0, 32'h44da942a},
  {32'hc40ce8b8, 32'h44097450, 32'h445d844b},
  {32'h424a9453, 32'h436f697e, 32'h45437786},
  {32'hc48dd90e, 32'h4366726a, 32'hc3d3997d},
  {32'h455ddc68, 32'hc442b515, 32'h43a9c512},
  {32'hc28fdca8, 32'h4493f63d, 32'hc48daab0},
  {32'hc324b2ee, 32'hc448490b, 32'h43fc422a},
  {32'hc4d544f2, 32'h440f1ac9, 32'hc21c27e6},
  {32'hc3027141, 32'hc5152080, 32'h442e2149},
  {32'h440df5e3, 32'h44f32a5e, 32'hc3722621},
  {32'hc3d34b0d, 32'h441329d9, 32'h44b5048c},
  {32'hc51556a6, 32'h43016d99, 32'hc480183e},
  {32'h44c8f93c, 32'h4221d169, 32'hc3fadc58},
  {32'h4362326e, 32'h44a3ea34, 32'hc51ae57d},
  {32'hc2b4037e, 32'hc4a8be21, 32'h453cd2e2},
  {32'h441dceee, 32'hc34ec8bb, 32'hc3ddc1ee},
  {32'h4441a285, 32'h434a3798, 32'hc2fd4bdc},
  {32'h442c7699, 32'hc31b38b0, 32'h44a2a2f7},
  {32'hc3fe0855, 32'hc38e86fb, 32'hc50517ed},
  {32'h43198917, 32'h436b58aa, 32'h44e6359d},
  {32'hc40375c1, 32'h4268d5f4, 32'hc54d23f2},
  {32'h44f43c72, 32'hc3bb04e7, 32'h44078fcc},
  {32'hc293c446, 32'h449210b7, 32'h450d860a},
  {32'h43f5830a, 32'h44c124a5, 32'hc512563f},
  {32'hc4199c69, 32'hc438850f, 32'h444bfeee},
  {32'h43cda4d5, 32'hc3c78384, 32'h44b2aecd},
  {32'hc374ade2, 32'h450d7b11, 32'h43fa3634},
  {32'hc4289a22, 32'hc4ac6bda, 32'h43a66712},
  {32'h43b66838, 32'h449e5aaa, 32'h41ac5073},
  {32'h448a028b, 32'hc3777fb3, 32'h43b49b75},
  {32'hc3a7f190, 32'hc330a911, 32'hc4d0e05d},
  {32'hc49054f7, 32'hc2ef7ab4, 32'hc2a1c82b},
  {32'hc48e7bda, 32'hc42a7db6, 32'hc4942272},
  {32'h43416420, 32'h44300f91, 32'h43957add},
  {32'hc477ed9a, 32'h424c2970, 32'h43940f53},
  {32'hc415345f, 32'hc546a2eb, 32'h426d10fb},
  {32'hc31815c9, 32'h450adf73, 32'hc2a4ccc9},
  {32'h42270a98, 32'hc4940345, 32'h43283100},
  {32'h415a1800, 32'h4575fcd8, 32'hc3a8a582},
  {32'h45169211, 32'hc47a5f93, 32'h43f52e83},
  {32'hc297a09c, 32'hc449dcd7, 32'h4419e750},
  {32'hc36fd26b, 32'h44336998, 32'hc38981ea},
  {32'hc24867c0, 32'h42e3e053, 32'h449ab685},
  {32'hc49eb576, 32'hc416f8ee, 32'h4440db5b},
  {32'hc3de692a, 32'h41b7e9e5, 32'hc50975a4},
  {32'hc4cbf7e1, 32'h434e23de, 32'hc178841c},
  {32'h43e23d65, 32'h44e1a4b2, 32'hc3d5e812},
  {32'hc2b73360, 32'hc312e700, 32'h451e67ab},
  {32'h43a6874c, 32'h420c1677, 32'hc3858c18},
  {32'hc46c9a5d, 32'hc25eb184, 32'hc369fdc6},
  {32'hc36b7a38, 32'hc41adaa7, 32'h44d5960f},
  {32'h4517ecfc, 32'hc39fa25c, 32'hc4480360},
  {32'h44354a78, 32'h448922eb, 32'hc40aba2a},
  {32'hc49fe6c9, 32'hc36ca452, 32'h4202c1e2},
  {32'h4375bfc8, 32'h443a1c0a, 32'h423e8d39},
  {32'hc49f1687, 32'hc3e5aa38, 32'h448a6b63},
  {32'h43951df0, 32'h3fc63a50, 32'hc4ddd4f1},
  {32'hc491b23c, 32'h4292bf76, 32'hc3bb6e86},
  {32'h44ad9687, 32'hc33ee99b, 32'hc4206d3a},
  {32'hc4dbf33b, 32'hc35919b3, 32'h4374b803},
  {32'h45726736, 32'h42bb7093, 32'h43fa2d21},
  {32'hc4d13232, 32'hc4851fcd, 32'hc33e48eb},
  {32'h448570f2, 32'h44519c83, 32'h43e39653},
  {32'hc3f42535, 32'hc2943ba6, 32'hc32533cb},
  {32'h43ae4228, 32'h44b10a63, 32'hc3e92756},
  {32'hc55302de, 32'hc346955d, 32'h432fa4b4},
  {32'h44a55e7d, 32'hc38fba30, 32'hc281befc},
  {32'hc36f2afc, 32'hc3ba5183, 32'h4394680e},
  {32'hc4153637, 32'hc481da88, 32'hc42e2d9e},
  {32'h434823bc, 32'h44b3969f, 32'h4430171c},
  {32'h44bb77ad, 32'hc3f998ce, 32'hc3b1303a},
  {32'h43ec2d00, 32'h448d390c, 32'h43b7d7e1},
  {32'hc33814f6, 32'hc554c3b3, 32'hc39a400d},
  {32'h44f186c9, 32'hc3db6c51, 32'h4330e998},
  {32'hc4ced53d, 32'hc3613826, 32'hc44b3508},
  {32'h444c13cc, 32'hc3b4322f, 32'h445f325c},
  {32'h43e64188, 32'hc4957a45, 32'hc3a574a8},
  {32'h4476fb48, 32'hc40b58ec, 32'h443a11ab},
  {32'hc3b04538, 32'hc4ce83a4, 32'hc3cd6294},
  {32'h4333bd0c, 32'h4407bcae, 32'hc38f60e6},
  {32'hc52ed984, 32'hc29a0303, 32'h41325eb1},
  {32'h432ecb18, 32'h43c041ad, 32'h453ed0f8},
  {32'h433d5910, 32'hc4bb995b, 32'hc3765ee2},
  {32'h446f9ac0, 32'h444d0e5c, 32'h447449d6},
  {32'h420c3330, 32'hc3c72ed2, 32'hc4c901b3},
  {32'hc326f2a8, 32'h4488c3b7, 32'h437ee50e},
  {32'hc3157a1c, 32'hc535c11e, 32'hc313a66f},
  {32'h42f0ff94, 32'h44eb7d45, 32'h43f2e906},
  {32'h445086dd, 32'hc4183c4e, 32'hc400d4f4},
  {32'h44cfa4bf, 32'h4400ded5, 32'h42c50260},
  {32'hc507ddba, 32'hc3fd204b, 32'h43514186},
  {32'h443c731f, 32'h43c58ae5, 32'h43ee81fd},
  {32'hc43f063c, 32'h42fc70f2, 32'h43392149},
  {32'h453c8360, 32'hc2f4c36e, 32'h44693cc9},
  {32'h449a5489, 32'hc452d3ae, 32'hc48e0e2e},
  {32'hc338a46a, 32'hc312e55f, 32'h44a6b734},
  {32'h430e035a, 32'hc3fac285, 32'h425e64e4},
  {32'hc3e4059e, 32'h43953193, 32'h44b64d5b},
  {32'h44453ef8, 32'hc400cdcf, 32'hc37dc6b3},
  {32'hc165bee8, 32'h44766602, 32'h4452fd06},
  {32'hc37cab33, 32'hc4a55274, 32'hc4d65450},
  {32'hc3eed99d, 32'h4429c6f1, 32'h452730e6},
  {32'h45470b17, 32'h43b43e76, 32'h43be3a94},
  {32'h430bbc24, 32'hc30423f4, 32'h44c23418},
  {32'hc31aa0d5, 32'hc35f5292, 32'hc3e89d36},
  {32'h43e2d7d8, 32'hc4912e3f, 32'h44cbdbb7},
  {32'h44da72e7, 32'hc44f1176, 32'hc1a2aee9},
  {32'hc3b04802, 32'hc21dc15c, 32'h44fa0369},
  {32'h44769b62, 32'h42c8d78c, 32'hc3f74634},
  {32'hc4025717, 32'h44943808, 32'h44476b92},
  {32'h447ca2a4, 32'hc49f3489, 32'hc476a50c},
  {32'hc4e92b7d, 32'hc41da7c5, 32'h43a7fca8},
  {32'h451c6f59, 32'hc4b0017e, 32'h439146e9},
  {32'h40553000, 32'h44fe10a4, 32'h430d7750},
  {32'hc33f9183, 32'hc4fb31e1, 32'h43986193},
  {32'hc46b6c19, 32'h4522b56f, 32'h424202ae},
  {32'h4523948e, 32'h435f0c46, 32'hc3f9e0a7},
  {32'hc419a632, 32'h441b715b, 32'h426bb812},
  {32'h455a84a7, 32'h434ce523, 32'h4360c7bd},
  {32'hc4e70496, 32'hc4153d8e, 32'h436ad138},
  {32'hc4e50b30, 32'hc1926a46, 32'hc3a85622},
  {32'h43a21344, 32'h439c37c6, 32'hc2fbf52f},
  {32'hc55f6d76, 32'h441e5388, 32'hc3b50a21},
  {32'h43ee4b30, 32'h44273231, 32'h43f91017},
  {32'hc4318680, 32'h42d24204, 32'hc2f1fecb},
  {32'h43e44b50, 32'hc4b9bcb0, 32'h41d58934},
  {32'hc53fe7e6, 32'hc37c3acc, 32'h436794e1},
  {32'h45050724, 32'h43209503, 32'hc39d7e2c},
  {32'hc5089bfd, 32'h44291266, 32'hc224e2ee},
  {32'h44aa57be, 32'hc4b5d461, 32'h428b34e8},
  {32'h44874200, 32'hc37f3be2, 32'hc41a400f},
  {32'h43d9fdfc, 32'h42576547, 32'h44d1bf38},
  {32'hc48e593e, 32'hc3ff3398, 32'h440a3301},
  {32'h43d96347, 32'hc4190144, 32'hc3fa040c},
  {32'hc469c807, 32'h40909afc, 32'h440da226},
  {32'h447cfd30, 32'hc40a6ca4, 32'hc378e434},
  {32'hc3ef6ae7, 32'h429c0b20, 32'hc14d00a0},
  {32'h43813bf0, 32'hc45a206b, 32'hc474b170},
  {32'hc45e2f9b, 32'h4466ea4d, 32'hc141e4d4},
  {32'h440a51f2, 32'hc3fb7bd5, 32'h426f2581},
  {32'hc58476ca, 32'hc38f2eeb, 32'h4256211b},
  {32'h4529e772, 32'hc3902943, 32'hc48288a0},
  {32'h43431ac6, 32'hc281c48c, 32'h426b0364},
  {32'hc4023b39, 32'hc3c59c01, 32'hc4f86345},
  {32'hc4a84c40, 32'h43f4000e, 32'h441d186c},
  {32'hc394981c, 32'hc1fde29b, 32'hc3932afe},
  {32'hc36e647c, 32'h448c797e, 32'h44c0f49b},
  {32'h43ff49b4, 32'hc400e18e, 32'hc50f5e9a},
  {32'h444e67b4, 32'hc31bc51a, 32'hc525e87c},
  {32'h4294bfe6, 32'hc388d473, 32'h45521df1},
  {32'h44b5acda, 32'h43b0d51b, 32'hc38c0141},
  {32'hc49210a8, 32'hc3ccf6e8, 32'h442ad54f},
  {32'h41b7a400, 32'h4535ec86, 32'h42886695},
  {32'h44c7442b, 32'hc401d298, 32'hc363ced0},
  {32'h45137c28, 32'h446ae1e7, 32'h4213743c},
  {32'hc55d411e, 32'hc3bc521c, 32'h43aa6dca},
  {32'h437f91b9, 32'h448faa3f, 32'h428df9f2},
  {32'h432ddc20, 32'hc3144a33, 32'h43fae5b5},
  {32'h43d320c0, 32'h444afd10, 32'h441c5414},
  {32'h44024609, 32'hc27c0a2a, 32'h43800d0d},
  {32'h43d4ae0d, 32'h43d21de2, 32'h44d55d12},
  {32'h43b78ac6, 32'hc4221e0f, 32'hc446c7e0},
  {32'hc36230c1, 32'h431c4f4d, 32'h44ca7674},
  {32'h41d211c1, 32'hc46a1e41, 32'hc487b7f9},
  {32'h440cb7c8, 32'h4443b797, 32'h44c4c44f},
  {32'hc367eec0, 32'hc43e72f8, 32'hc3f71415},
  {32'h4580e5b3, 32'h414634f8, 32'h419c2494},
  {32'hc5792768, 32'h43ce0852, 32'hc393f05b},
  {32'hc4e65c44, 32'hc2a70fe9, 32'hc3105c37},
  {32'hc340ec8c, 32'hc4defd24, 32'hc4a02a6c},
  {32'hc304e27c, 32'h44a51d73, 32'h4486e4e3},
  {32'h414b8eb0, 32'h42a6c3a8, 32'hc4ced263},
  {32'h44cb0b8b, 32'h44598b31, 32'h4443695a},
  {32'hc4d312da, 32'h4385e659, 32'hc4c2a602},
  {32'hc0ae0368, 32'hc31d2cb6, 32'h44b82a90},
  {32'h44279216, 32'hc31db7ac, 32'hc2cb2dd4},
  {32'hc20009b8, 32'hc517864b, 32'hc27fb00e},
  {32'h44b8ac4b, 32'h4498b041, 32'h43f69426},
  {32'h44329bdc, 32'hc48bcd88, 32'h4183a900},
  {32'h43ee44a8, 32'h45130cda, 32'h43184939},
  {32'hc4479758, 32'hc4f282fc, 32'hc2843141},
  {32'h44ab6f5e, 32'h439f448e, 32'hc4053a40},
  {32'hc4b383e1, 32'hc344d0c3, 32'hc3d15445},
  {32'h4534502a, 32'h4390616a, 32'h44490fa7},
  {32'hc5050689, 32'h42e28db9, 32'h43c97dbf},
  {32'h44b3bc8a, 32'h444fe780, 32'h42ca83e8},
  {32'hc39eaedd, 32'hc4630452, 32'h443a5867},
  {32'hc20be10d, 32'h44e8560c, 32'hc2b45510},
  {32'hc3802c1c, 32'hc2de89c6, 32'h450408a4},
  {32'h43133af1, 32'h43a64dc9, 32'hc4d5ec60},
  {32'h4481acbc, 32'hc0be9ea7, 32'h4481e30f},
  {32'h43cccffc, 32'hc3906827, 32'hc4c5d5c4},
  {32'hc489a344, 32'h41a7cb88, 32'h44466c53},
  {32'h43abfba4, 32'h43abc7e6, 32'hc4bc8c02},
  {32'hc50a4cc6, 32'hc46a5437, 32'h433b700d},
  {32'h44065d90, 32'h450df247, 32'h422b2613},
  {32'hc40052c9, 32'hc208bbe5, 32'hc3a1766f},
  {32'h444ca537, 32'h44103952, 32'hc4abcc20},
  {32'hc3c8284c, 32'hc53c1e74, 32'h43028397},
  {32'h4434b699, 32'h438aa7bd, 32'hc41257ea},
  {32'hc3f87a10, 32'h4398fd25, 32'h449b5886},
  {32'h44e53aa4, 32'hc3c691f0, 32'hc4b4e80c},
  {32'h44c8873d, 32'hc4c7b680, 32'hc3b7ded4},
  {32'hc5099f9c, 32'h44994849, 32'hc3a9608c},
  {32'h43f78c18, 32'hc49a0244, 32'hc3335648},
  {32'hc3ffaad7, 32'h451213eb, 32'h414649ac},
  {32'h41d8500c, 32'hc53baa4f, 32'hc2503e4f},
  {32'h44b573cd, 32'h42d06648, 32'hc2dde637},
  {32'h440ddc44, 32'h44502786, 32'h43660e13},
  {32'hc50ec91e, 32'h4427c5e7, 32'h441e129f},
  {32'h453d9347, 32'hc3e3613f, 32'h43f683b0},
  {32'hc32ac1a2, 32'h4485412a, 32'h438aa9cb},
  {32'h443b1d65, 32'hc439d732, 32'h44186d10},
  {32'hc429ed8e, 32'h444a83c5, 32'hc2e98e24},
  {32'h4426b89a, 32'hc47698f3, 32'hc2420674},
  {32'hc495b372, 32'h43f735a0, 32'hc42e386e},
  {32'h43e21bb3, 32'h4393f589, 32'h4368358b},
  {32'hc506f641, 32'hc3182231, 32'hc4269ee1},
  {32'h437a0539, 32'h43370cff, 32'h45152cf4},
  {32'hc447cf72, 32'hc31ee60c, 32'hc3f32789},
  {32'h44145748, 32'hc4c05bd2, 32'h43eb2874},
  {32'hc360201b, 32'h451acf2d, 32'hc37f7418},
  {32'h4547c3da, 32'h43d93479, 32'h428af718},
  {32'hc490e3dc, 32'hc31733e1, 32'hc4b2cd84},
  {32'h4386e14f, 32'hc411f6dc, 32'hc29d5bd5},
  {32'hc2cf15fb, 32'h42405443, 32'hc374a56e},
  {32'h43326f30, 32'h4431339d, 32'h44ea332c},
  {32'hc535bc8a, 32'h43b4f8d1, 32'hc403c6c8},
  {32'h434b8de6, 32'h435ed564, 32'h431f10d9},
  {32'hc4bb78df, 32'h4323dc96, 32'hc3de8fa3},
  {32'h44806a90, 32'h43ecafc7, 32'h449fdf46},
  {32'h431238f7, 32'h44aac9aa, 32'hc410a4f6},
  {32'hc4b46d30, 32'hc36b53e7, 32'h4217e75f},
  {32'h4498daa3, 32'hc4948744, 32'h44082db6},
  {32'hc49db519, 32'h44bd957f, 32'h442d9199},
  {32'hc4a18a0e, 32'h4371a575, 32'hc3df200e},
  {32'hc4b49f33, 32'h442c5c00, 32'hc4164d83},
  {32'h42978e5a, 32'hc524bfcf, 32'h43f2541c},
  {32'h4341f110, 32'h44f41aa4, 32'h44bb0ed8},
  {32'hc47473ea, 32'hc402adf9, 32'hc3776526},
  {32'hc40275d8, 32'h4326fb77, 32'h438c9086},
  {32'h43bd5d64, 32'hc2b10c06, 32'h44de0034},
  {32'hc3331b3a, 32'h4462053e, 32'hc328ca30},
  {32'h43c979aa, 32'hc4259c53, 32'h4487c9c2},
  {32'h4304cf9c, 32'h441c65f8, 32'hc4675f7e},
  {32'h43b89021, 32'hc4ee4d90, 32'h432be78f},
  {32'hc2e37a2e, 32'h444c79b5, 32'hc4b76397},
  {32'hc353954c, 32'hc3d917dc, 32'h4449dbe7},
  {32'hc545ef72, 32'hc3cc9265, 32'hc37c70d3},
  {32'hc42778d0, 32'h43fa46b4, 32'h439f9115},
  {32'h44a3a57b, 32'h43b339b0, 32'hc3a6238a},
  {32'h451521ac, 32'hc4770839, 32'hc3beb9e8},
  {32'hc499f7da, 32'h43849bdc, 32'h41824606},
  {32'hc2fee674, 32'hc3ea65e9, 32'h434e605a},
  {32'hc589b927, 32'hc32ffafd, 32'hc2c87a48},
  {32'h43e375a9, 32'hc4fb0cdd, 32'h4370c7a4},
  {32'h43c880b0, 32'h41d650d6, 32'h4489b3a2},
  {32'hc48afe63, 32'h44288973, 32'hc40c16cd},
  {32'hc4948400, 32'hc346dbd0, 32'h43eb4f4a},
  {32'hc428d428, 32'hc41187e0, 32'h44856f16},
  {32'hc3290810, 32'h429c9424, 32'hc4890216},
  {32'h432de9e4, 32'hc4a37333, 32'h420ed48f},
  {32'h44df1c3a, 32'h42c46ba2, 32'hc43033e8},
  {32'hc4a73098, 32'hc4498e9a, 32'h43abd6c5},
  {32'h44eaa731, 32'h43b8cddf, 32'h4320b907},
  {32'h44674f4b, 32'hc3f585cf, 32'h42947715},
  {32'hc4ba3a12, 32'hc3111566, 32'h44e1c50c},
  {32'h439c2ebc, 32'hc391e8a2, 32'hc465a3be},
  {32'h440950ee, 32'h4281000a, 32'hc4b13cac},
  {32'hc3dd7cfa, 32'hc4a2fc50, 32'h43c60e8d},
  {32'h4397f857, 32'h451144a2, 32'h4018adf5},
  {32'hc5485d66, 32'hc3354854, 32'h42bdf9da},
  {32'hc37e6bc0, 32'h45465211, 32'hc2ecaace},
  {32'hc214c980, 32'hc4585a60, 32'h42c5bb1c},
  {32'h44a5d856, 32'hc42d9d42, 32'hc3e92087},
  {32'hc5275182, 32'hc2b440f8, 32'h43c3d622},
  {32'h4484d257, 32'hc28b996c, 32'h42eaae97},
  {32'hc40111bb, 32'hc50b8821, 32'h43e929c3},
  {32'h42d54100, 32'h4525d125, 32'h4348c0e7},
  {32'h449f224d, 32'hc22184e9, 32'h4384a830},
  {32'h44c9749a, 32'h447be49c, 32'hc324adae},
  {32'hc49518c6, 32'hc4c4db16, 32'h43afd3e0},
  {32'hc4909738, 32'h43e6d39f, 32'hc3ded89a},
  {32'hc34f071c, 32'h445620ee, 32'hc2a78804},
  {32'hc4c5b8d3, 32'hc1ed21fb, 32'hc4029f04},
  {32'h44759c93, 32'h44158719, 32'h43ce3462},
  {32'hc338b679, 32'hc390ed07, 32'h438e44f9},
  {32'h442095d4, 32'h442cbd7b, 32'h44db7ec8},
  {32'hc41512ee, 32'hc40e04a4, 32'hc42ccf27},
  {32'hc406f5dc, 32'h44222706, 32'h440b2440},
  {32'hc551a387, 32'hc37ecec6, 32'hc18ff456},
  {32'hc3154200, 32'h44a7f8e7, 32'h451383f8},
  {32'h44155bcc, 32'hc46f3013, 32'hc1cd62fe},
  {32'hc3f804c4, 32'h44155f72, 32'h4438e4f7},
  {32'hc2076bd0, 32'h43ede990, 32'hc489f2ea},
  {32'h450946c9, 32'h42c80534, 32'hc306158b},
  {32'hc458a4a3, 32'hc49eb32e, 32'hc3a3a41b},
  {32'h43d1afdd, 32'h44f4a16d, 32'hc3786776},
  {32'h444894b0, 32'hc152a1f2, 32'hc3aa836b},
  {32'h44a28528, 32'h43b182bc, 32'h44115308},
  {32'hc49475e2, 32'hc40149f4, 32'hc4d2c618},
  {32'hc4ab1632, 32'h444717c6, 32'h4393f64c},
  {32'hc451ad92, 32'hc51f907a, 32'h438ce392},
  {32'h4519ea3d, 32'h449744cb, 32'hc40c4c2e},
  {32'h411c0294, 32'hc40ecf4a, 32'hc3c15f39},
  {32'h450b151e, 32'h4404d4fd, 32'h4348c69a},
  {32'hc522f96c, 32'hc3ee7478, 32'h438fc7e2},
  {32'h44aa8d23, 32'h440d721b, 32'h4361efd2},
  {32'hc5140b12, 32'h42d988ae, 32'hc31a311a},
  {32'h44781cfe, 32'h42d3fab4, 32'h442c713c},
  {32'h43a975fe, 32'hc400006c, 32'hc4cd6f50},
  {32'hc48eb5d6, 32'h446b94c5, 32'h447a2d87},
  {32'h43143794, 32'hc44087ea, 32'hc37b57f7},
  {32'h41e85ac0, 32'h440b4b5f, 32'h44d531e6},
  {32'hc307eb58, 32'hc49f021b, 32'hc500413b},
  {32'h4461746b, 32'h449a3b13, 32'h43977b0d},
  {32'hc306ae58, 32'hc432fe52, 32'hc5050adb},
  {32'hc3bd2606, 32'h4460bb8a, 32'h44b66fd1},
  {32'h4473d4fa, 32'hc310e82a, 32'hc4927a98},
  {32'hc38ca8ea, 32'hc3f13f2f, 32'h449b560f},
  {32'h43308a0e, 32'h44ed80c6, 32'hc4c0aece},
  {32'h43b584b7, 32'h44058581, 32'h42ba711b},
  {32'hc2f78423, 32'hc55430de, 32'hc37416ed},
  {32'hc4150e7a, 32'h44c57092, 32'h441cf585},
  {32'h44964d9d, 32'hc37134e4, 32'hc3b35fa9},
  {32'hc4a0c346, 32'hc2c3c6ac, 32'h44916c19},
  {32'h44f52de9, 32'h42a9ed1b, 32'hc3557150},
  {32'hc4fd1f92, 32'hc32a5b48, 32'h439f231e},
  {32'h44c596ff, 32'hc4ced296, 32'hc16d35a3},
  {32'hc537d24d, 32'h424d4edc, 32'h43d600a0},
  {32'h44b40291, 32'h4321b7a1, 32'hc2a663b6},
  {32'hc47cae4e, 32'h451af29f, 32'hc2ff26b1},
  {32'h4451b8ae, 32'hc2810e54, 32'hc20bdb2a},
  {32'hc41e083a, 32'hc2902a8a, 32'h4280eadb},
  {32'h4538c12d, 32'h43167f46, 32'h43800d06},
  {32'hc56834a9, 32'hc33ebcac, 32'hc3dad591},
  {32'hc4f0ab1c, 32'hc3e52d04, 32'h41107c73},
  {32'h44a53933, 32'hc3284b34, 32'hc2337b50},
  {32'hc3dad01a, 32'h438405e8, 32'hc53e5e18},
  {32'h43ea9940, 32'hc402450e, 32'h4530f776},
  {32'hc50bc9c2, 32'hc420f248, 32'hc3d2a748},
  {32'h450bc6d4, 32'hc455ecb9, 32'hc1d533f0},
  {32'hc45f3376, 32'h441d72c6, 32'h420cc148},
  {32'hc4003d55, 32'hc355c54d, 32'h4355c3cf},
  {32'hc489454f, 32'h44f1eeaa, 32'h4129d982},
  {32'h4367e7f0, 32'hc51e7d3b, 32'hc3e2c634},
  {32'hc403ade1, 32'hc397fcd9, 32'hc377069f},
  {32'h4528c4a4, 32'h4351a40c, 32'h436c8822},
  {32'h42d48e40, 32'h4388d362, 32'hc2886d41},
  {32'h42bb06e0, 32'h42891607, 32'hc4e51b76},
  {32'h430b7f30, 32'h43b87f49, 32'h4495b7f3},
  {32'h43a984b1, 32'hc433f4db, 32'hc4e8dd81},
  {32'h4400af18, 32'h4435ba35, 32'hc3120f93},
  {32'h44ac631e, 32'hc31d94bb, 32'hc3d66904},
  {32'hc49d15a6, 32'hc2e0b6ab, 32'h43785b85},
  {32'h4561b5ae, 32'hc448e89c, 32'h43d76990},
  {32'hc51667b4, 32'hc4030af1, 32'h435c26c2},
  {32'h451d4688, 32'hc2bd1eb2, 32'hc4697de1},
  {32'h43c3aae4, 32'h41090104, 32'h42cf4c0c},
  {32'h43f178e6, 32'hc4be56ea, 32'hc407d41c},
  {32'hc51adbac, 32'h43b06b57, 32'h43c9ec1a},
  {32'h4482d9cd, 32'hc40ec35f, 32'hc4034c31},
  {32'hc448e57a, 32'h44a7b6b4, 32'h44da0be2},
  {32'hc32d944e, 32'hc2f5eee4, 32'hc4457e36},
  {32'h43d749b0, 32'h43c05135, 32'hc52be5cb},
  {32'hc4b766b3, 32'hc3843294, 32'h449fca3a},
  {32'hc43fc18a, 32'hc33d2fc2, 32'hc3fc168c},
  {32'hc5009fef, 32'hc452b31f, 32'hc2d8a12b},
  {32'h43a52e34, 32'h4439f0c8, 32'h437e7834},
  {32'h448eb07c, 32'hc2aa3326, 32'hc39972d8},
  {32'h450ac2ab, 32'h44031db2, 32'hc38997ef},
  {32'hc28d42a0, 32'hc4c66b26, 32'hc30e75a3},
  {32'hc44da7e6, 32'h4249295e, 32'h438925ce},
  {32'hc41ab89e, 32'hc3d4ea13, 32'h44f141d1},
  {32'h44871203, 32'h430a1f4c, 32'hc490e088},
  {32'h43dfd2c0, 32'hc26c5df3, 32'h4476a9ad},
  {32'h439c3e2c, 32'h453539a7, 32'h43c92574},
  {32'hc4f42149, 32'hc4254ca8, 32'hc40d27f8},
  {32'h4529b4da, 32'h43934387, 32'hc29a98ad},
  {32'hc4bf826e, 32'hc46634b4, 32'hc3ad722a},
  {32'hc3c0ee08, 32'hc2088d3c, 32'h436e7bbb},
  {32'h428ba572, 32'hc27fe022, 32'hc4b6a591},
  {32'h44a49060, 32'h43176f79, 32'h4445ef61},
  {32'hc447b3a1, 32'h43052401, 32'hc497facf},
  {32'h44bea327, 32'h43183631, 32'hc3203941},
  {32'hc49d7452, 32'hc42bff2d, 32'hc429fdf8},
  {32'h43e58196, 32'h4544444f, 32'hc2ff54f8},
  {32'hc2605481, 32'hc3aebf89, 32'hc46216f8},
  {32'hc362cc2a, 32'h43fae05f, 32'h45004a3e},
  {32'hc319cdbc, 32'hc52f5c84, 32'hc4012168},
  {32'h43b14c00, 32'h41cbfcde, 32'h436645e6},
  {32'hc3cdda02, 32'h43ff3acd, 32'h42a205a3},
  {32'hc22fce22, 32'hc5445694, 32'hc2f40f94},
  {32'hc3086ec8, 32'h455328d8, 32'h42ee6aee},
  {32'hc402d561, 32'hc45e1629, 32'h4409c2e8},
  {32'h440a1de3, 32'h441333ce, 32'h43433a5f},
  {32'hc40afa76, 32'hc503ba78, 32'h4313d3d1},
  {32'hc45e2f86, 32'h436b4985, 32'hc394becd},
  {32'hc43f82d0, 32'h43d4b6b1, 32'h435658c2},
  {32'h44e3b338, 32'h441e4633, 32'h4404e7a8},
  {32'h44820a38, 32'hc422d42e, 32'h42ccb81c},
  {32'h4364af10, 32'h446feced, 32'hc2965d4a},
  {32'hc2010038, 32'hc4a03e90, 32'h443dcdd1},
  {32'hc3310685, 32'h44ca144e, 32'h428b1af4},
  {32'hc47a83d0, 32'hc38b2d03, 32'h4414b7cd},
  {32'h447920b7, 32'h450aa2c4, 32'hc3dd738e},
  {32'hc39af6ef, 32'hc3c4865b, 32'h4306eb9e},
  {32'h44793599, 32'h43b2b4be, 32'hc468253b},
  {32'hc4787826, 32'hc41cd170, 32'hc2d269ba},
  {32'h43684588, 32'h43f1f3c2, 32'h439cb0aa},
  {32'hc542c3f8, 32'hc3873264, 32'h439c50da},
  {32'h44952e23, 32'h4466390a, 32'hc4b3441e},
  {32'hc4845bde, 32'h438b5fbe, 32'h43fb324b},
  {32'h4404c2c1, 32'h44b35205, 32'hc3fed49f},
  {32'hc40b3828, 32'hc3dceef4, 32'h43ad8fe1},
  {32'h44aad171, 32'h43eaf17b, 32'hc2c17227},
  {32'hc412cde9, 32'h430abbe0, 32'h451ddf63},
  {32'h448cb13e, 32'hc3423701, 32'hc302e996},
  {32'h45112462, 32'hc48926ed, 32'hc41d65fe},
  {32'hc42b0850, 32'hc40e77d1, 32'h44f9a5ca},
  {32'hc31a9511, 32'hc4bb248e, 32'h43cb35df},
  {32'hc483fad9, 32'h4501ef33, 32'h43e2d431},
  {32'hc310b057, 32'hc5736561, 32'h42aa3a9f},
  {32'h4390ccbf, 32'h448ed2d7, 32'hc3f2e3ae},
  {32'h4400ff2f, 32'hc457d86c, 32'hc4834832},
  {32'hc57efa5d, 32'h41b4cd42, 32'hc40d7bca},
  {32'h451027ff, 32'hc4081fd3, 32'h439d663f},
  {32'hc350c08c, 32'h44650bc5, 32'hc47827b8},
  {32'h43a586a2, 32'hc455c217, 32'h4438fd08},
  {32'h43b7276c, 32'h442d357e, 32'hc48247cc},
  {32'h42b7c5ea, 32'hc22aead1, 32'h44433096},
  {32'hc478c167, 32'h443aa458, 32'hc40cb4b7},
  {32'hc4a79d82, 32'hc30a74e5, 32'hc3416da0},
  {32'hc5221333, 32'h42d02af3, 32'hc47d29ee},
  {32'h43c0a7d8, 32'hc3562b1e, 32'h441ea8f3},
  {32'hc4fc47c7, 32'h43c2162c, 32'h43fc7409},
  {32'h44df0f73, 32'hc48fd994, 32'hc2903184},
  {32'hc3a86f54, 32'h454636aa, 32'h42f21c48},
  {32'h449bba27, 32'hc3879f93, 32'h438d3e6f},
  {32'hc34b9dae, 32'hc388c5ff, 32'hc4d89514},
  {32'h44a9e5ee, 32'hc47b6483, 32'h40cf2994},
  {32'hc2d940ce, 32'h4359a896, 32'hc3c83d97},
  {32'h452ae484, 32'h4344fd83, 32'h441a130f},
  {32'hc50e4f59, 32'hc3aabd1b, 32'hc3f54eaf},
  {32'hc3b64182, 32'hc2c8639d, 32'h43bb4eeb},
  {32'h4352874e, 32'hc4d69727, 32'hc49e8351},
  {32'h4386f023, 32'hc43cbcaf, 32'h44177430},
  {32'h440ea841, 32'h441c1a93, 32'hc47192e0},
  {32'hc4a7e465, 32'h439f3c75, 32'hc364d06c},
  {32'h43d9bbb2, 32'hc4ac2caf, 32'h43d767c3},
  {32'hc418db7c, 32'h44522b13, 32'hc304a5c8},
  {32'hc23888a0, 32'hc38fc24d, 32'h43dc13a1},
  {32'h43246b9a, 32'h45385482, 32'h439a3302},
  {32'h422813e0, 32'hc44245bc, 32'h4516220f},
  {32'h44afb94b, 32'hc4ad5e06, 32'h449d60bf},
  {32'h439c9694, 32'hc51a5fa8, 32'hc4f89c50},
  {32'h44972fcb, 32'hc3977d6c, 32'hc300b136},
  {32'hc4b6505b, 32'hc2083160, 32'h430fcc3e},
  {32'hc3c34950, 32'h43180e18, 32'hc4b65919},
  {32'h4379be35, 32'hc3d61b90, 32'h44e39b8e},
  {32'hc44b600e, 32'hc342bf41, 32'hc388ebad},
  {32'h4465270e, 32'hc4874872, 32'h4433e892},
  {32'hc52d3ac5, 32'h426c8ba7, 32'hc343c68c},
  {32'h42fe7ba0, 32'hc3d2c91e, 32'h43c2624e},
  {32'hc5953cb8, 32'h423cdbce, 32'h43380a3b},
  {32'h44c703c8, 32'hc280c8f6, 32'h42060473},
  {32'hc51729bb, 32'hc29f9f9c, 32'h4418dc9a},
  {32'h444a94e9, 32'hc497c65d, 32'h4193ad1c},
  {32'hc305e158, 32'h4525bc57, 32'hc32fd343},
  {32'h44a06dcb, 32'h4402294e, 32'h4400b0c7},
  {32'hc542747d, 32'h44163213, 32'h429b99da},
  {32'h4419f857, 32'hc50ac257, 32'hc38d2cfb},
  {32'hc3cd8456, 32'hc437861f, 32'hc3570147},
  {32'hc473c5b1, 32'h441c09d7, 32'hc5045ac9},
  {32'hc386c53a, 32'hc26f36ac, 32'h451751d6},
  {32'hc518d482, 32'hc3ae3fd5, 32'h43212eab},
  {32'h443a8bfe, 32'h44ac14e3, 32'hc39f3991},
  {32'h44e55a71, 32'hc3d42965, 32'h4272988e},
  {32'h4382cb7a, 32'h44e5f805, 32'hc37a9666},
  {32'hc4c6caf0, 32'h42e8d18a, 32'h444ee928},
  {32'h43bc3c38, 32'hc35e0063, 32'hc3f0b10d},
  {32'h4505eec5, 32'hc32f59d5, 32'h436da397},
  {32'h44079223, 32'h443bdff2, 32'h452f19d0},
  {32'h442023fb, 32'hc415d777, 32'hc4c765e6},
  {32'h440e03ce, 32'h4523c360, 32'hc306b6c7},
  {32'hc4d3adc1, 32'hc44a9ffe, 32'h43d99089},
  {32'h432676f4, 32'h43efbc19, 32'hc3462607},
  {32'hc481aaee, 32'hc3c964f4, 32'h44b6411b},
  {32'h445e7216, 32'h43a94add, 32'hc392550a},
  {32'hc4936612, 32'hc3dfc529, 32'h42bb4fa0},
  {32'h451174d0, 32'hc40fcfc3, 32'h423f9168},
  {32'hc4e98d0c, 32'hc38fd067, 32'hc334b1c9},
  {32'h44c6eaba, 32'h446ef107, 32'h427c34b2},
  {32'hc425ac8e, 32'hc4b90aea, 32'hc379ab23},
  {32'h42fdef10, 32'h43e661ee, 32'h43a631fa},
  {32'hc4ae4e55, 32'hc2fa188d, 32'hc1e0f547},
  {32'hc34ed7d8, 32'h44e257c1, 32'hc3cb65e3},
  {32'hc4989d7c, 32'hc4d439b9, 32'h436e3738},
  {32'h4514b165, 32'h427e4ffd, 32'hc3a2b1fa},
  {32'h42c8f6aa, 32'h43939ddb, 32'h4341dd47},
  {32'h432124eb, 32'h4311983f, 32'hc4e08b96},
  {32'h44d24e3e, 32'h4396541d, 32'h4429e677},
  {32'hc44d3c1a, 32'hc3c26dc7, 32'hc361b5af},
  {32'h434a35c8, 32'h41cf3cb8, 32'h447deb7f},
  {32'hc3c3163a, 32'hc50125b4, 32'hc34842be},
  {32'h44b587ad, 32'hc31c6c7e, 32'hc32d7881},
  {32'hc4bb09da, 32'hc4120b7e, 32'hc4b1c232},
  {32'h43b80994, 32'h44f09537, 32'h44693627},
  {32'h4281e1fa, 32'hc40952ce, 32'hc249f208},
  {32'h433adcfe, 32'hc451a183, 32'h44a38a3f},
  {32'hc31fc700, 32'hc3787fb8, 32'hc4988e05},
  {32'hc327be4c, 32'h44708d71, 32'hc3704480},
  {32'hc448e26a, 32'h4124c633, 32'hc4d1af96},
  {32'hc25ccbd2, 32'h44803e9e, 32'h452395f8},
  {32'hc52b506d, 32'h42ee4740, 32'h4356fd80},
  {32'h4508407e, 32'h439d585c, 32'h43351f4c},
  {32'hc39c8376, 32'h430cd95c, 32'hc4dba0f8},
  {32'h433ab42a, 32'h4447c39f, 32'h43395303},
  {32'hc51e8ac7, 32'hc435bf0a, 32'h4320e8d5},
  {32'h4380b2b5, 32'h455cebbc, 32'hc301cdfb},
  {32'h431ea5e6, 32'hc5106844, 32'h431f7313},
  {32'h444acb32, 32'h44a4e890, 32'hc39fc25e},
  {32'hc46b1263, 32'hc4fdc30c, 32'h42b97c85},
  {32'hc49a5c9c, 32'h43177f5d, 32'h44000ccf},
  {32'hc58ff3ee, 32'h4201fa1a, 32'hc38b4a83},
  {32'h45773497, 32'h437440a0, 32'hc33596af},
  {32'h4458daf3, 32'hc41d54c3, 32'hc42d249c},
  {32'hc35c0334, 32'h449a1f0a, 32'h43ff5563},
  {32'hc19b6062, 32'hc43e7823, 32'hc3f23751},
  {32'hc480a6ff, 32'h43dbc7de, 32'h44643a28},
  {32'hc1b58a1e, 32'hc4cacf7c, 32'hc3a99b64},
  {32'hc3f42a58, 32'h43ac50b2, 32'h44ff9876},
  {32'h454a21b9, 32'hc39c9817, 32'hc43d98d2},
  {32'h4365c6f0, 32'h44b3fd0f, 32'h44c37de3},
  {32'hc37fe04f, 32'hc468c446, 32'hc4a4d96c},
  {32'hc3d727e4, 32'hc372aa92, 32'h44a43c70},
  {32'hc4af8c08, 32'h44c19c88, 32'hc4919b9c},
  {32'hc407ec87, 32'hc3abc2c7, 32'h43f10fe9},
  {32'h451ea5fb, 32'hc3b5ebcc, 32'hc25873a0},
  {32'hc4487d7c, 32'h43d82218, 32'h44934aa9},
  {32'hc30868e8, 32'hc487b7fd, 32'hc329136e},
  {32'h443c5dc0, 32'h443efd42, 32'h455264fb},
  {32'hc1ec7860, 32'hc4d4c1f7, 32'hc4ada032},
  {32'hc420721a, 32'hc2505774, 32'h432f3783},
  {32'h432c48b8, 32'hc569757d, 32'hc427c4b3},
  {32'hc50aedc7, 32'h450184fc, 32'h436edef6},
  {32'hc2fd0b78, 32'h424a4350, 32'hc3577aa3},
  {32'hc47d6dae, 32'hc38238ab, 32'hc385e7e6},
  {32'h445fbafc, 32'hc5158fff, 32'hc32504b5},
  {32'hc53f294f, 32'hc329c5b1, 32'h43657cae},
  {32'h44f2f7d9, 32'hc3235a71, 32'hc3d07735},
  {32'hc59112d6, 32'h41125590, 32'h41876619},
  {32'h449e7748, 32'hc35cee76, 32'hc3aad813},
  {32'h4488d81e, 32'hc1de336c, 32'h42f20e46},
  {32'hc54e605e, 32'h42be0823, 32'hc39be5af},
  {32'hc2c41b90, 32'hc1b34424, 32'h4549ac8b},
  {32'h44ba80f0, 32'hc3d3049a, 32'hc364ab33},
  {32'h436fc8fc, 32'hc4d4f7f7, 32'h42a504c6},
  {32'hc4d427ef, 32'h443da8bf, 32'h43b11be0},
  {32'hc3833105, 32'hc489ff54, 32'hc18fa818},
  {32'hc5088e30, 32'h443f6b3f, 32'h42a89df2},
  {32'h439c63d6, 32'hc55d8e7f, 32'h41a63bfb},
  {32'hc3540032, 32'hc466c712, 32'h43b1b76a},
  {32'h4477498e, 32'hc4144abe, 32'hc3bc4df2},
  {32'hc49dd555, 32'h440d8260, 32'hc4d46f8b},
  {32'h4388af61, 32'hc4704c8c, 32'hc3a612c4},
  {32'hc403539f, 32'h4502403a, 32'h430e019e},
  {32'h42f73db0, 32'hc4b4324a, 32'hc2d2dc4a},
  {32'h44832c60, 32'h44057f1f, 32'hc382fd22},
  {32'h44463624, 32'hc3c7fb3f, 32'hc4dafad7},
  {32'h43b13fe6, 32'h45082fed, 32'h43f92f83},
  {32'h43d4e0a8, 32'hc41429d9, 32'hc2fa215e},
  {32'hc47e1434, 32'h442d6c3d, 32'h44e15699},
  {32'hc42ff588, 32'hc3878816, 32'hc4297d14},
  {32'h44ac13ec, 32'h4407afd7, 32'hc33ded7c},
  {32'h43b791b4, 32'hc415972c, 32'hc489ef0a},
  {32'hc4b30870, 32'hc1a6afb5, 32'h43e5c762},
  {32'h448d2cea, 32'hc3979915, 32'h3e47a668},
  {32'hc47fd23f, 32'h4431a638, 32'h44ac1231},
  {32'h44c394fd, 32'hc44664cd, 32'hc4abc73a},
  {32'h44786c21, 32'h441d6f2e, 32'hc4bbef21},
  {32'hc50aa21f, 32'h43b41b4f, 32'h401d1dd7},
  {32'hc4302cba, 32'h4404ee10, 32'hc41bff58},
  {32'hc4cc02bc, 32'hc3a15730, 32'hc3d042ff},
  {32'hc39b4987, 32'h452d14c2, 32'h44266803},
  {32'h4484b710, 32'hc40238f7, 32'hc32da4f8},
  {32'h449c1f88, 32'h4507f2fe, 32'h42a45ac1},
  {32'hc4e95c75, 32'hc4d50b67, 32'h4353dfe9},
  {32'h44d09f71, 32'hc3f88964, 32'hc2a66c52},
  {32'hc48ca904, 32'hc38731ca, 32'h43a32311},
  {32'h43ab5720, 32'hc36c447f, 32'hc2919e6b},
  {32'hc3d78c82, 32'h43810f2a, 32'h43216de8},
  {32'h43bbfa00, 32'h43c13681, 32'h4492322c},
  {32'hc40fac10, 32'hc30d84ee, 32'hc52c7aec},
  {32'h449e7a5e, 32'h42cc7d8a, 32'hc39855a9},
  {32'hc35c1a28, 32'hc5143ac9, 32'hc4078ab1},
  {32'h437b5bde, 32'h43df204c, 32'h45218d08},
  {32'hc1bf38ab, 32'hc310753f, 32'hc47ec9cf},
  {32'h4545d4ee, 32'hc2dbc43f, 32'h44220ca9},
  {32'hc46cac98, 32'h445e4b0e, 32'hc3ca2a7e},
  {32'h43f83c98, 32'h442ef15e, 32'hc36f13c5},
  {32'hc4ec5918, 32'hc37d66e3, 32'hc458ed67},
  {32'h44ec77d4, 32'h44096826, 32'hc15a179d},
  {32'hc4f94545, 32'hc400552d, 32'hc381479f},
  {32'h44a0feb4, 32'h4443081e, 32'h4411eebf},
  {32'hc4d6d134, 32'hc47ebca3, 32'hc34fec43},
  {32'hc43ee5ed, 32'h443eadd1, 32'h424be184},
  {32'hc4d61ab8, 32'hc38adbb0, 32'h4253e9f3},
  {32'hc3ab0b3c, 32'hc4c0a511, 32'hc3cd29d5},
  {32'h44fdb320, 32'h4415bf2a, 32'h4449d514},
  {32'hc292c6db, 32'hc4138f7f, 32'h43d7d2bc},
  {32'h455a82e1, 32'h42f412e6, 32'h4347a05c},
  {32'hc211d2e0, 32'hc51ac61a, 32'hc3407b85},
  {32'h44a206e7, 32'h43812534, 32'hc30f6427},
  {32'hc59e9339, 32'hc31e3d16, 32'h43b5b8b8},
  {32'h453ef06d, 32'h429ca26a, 32'hc10747b7},
  {32'h444905bb, 32'h438640ca, 32'hc343e2fc},
  {32'h4528606e, 32'hc184089d, 32'h43b59471},
  {32'hc45807c9, 32'hc479b9f7, 32'h44465345},
  {32'h439ee649, 32'h44624ca1, 32'hc407f13e},
  {32'hc42b3010, 32'hc3f2d25e, 32'h445a67dc},
  {32'h44066e36, 32'h45327bd6, 32'hc40ad0c2},
  {32'h442bf0c4, 32'h437a35b6, 32'h4502c3d7},
  {32'h44de0000, 32'h43cb419e, 32'hc4138e9d},
  {32'hc4d7f6ef, 32'h430207ec, 32'h44211b21},
  {32'h4348eec3, 32'h43b57bb7, 32'hc3accd48},
  {32'hc4c4410c, 32'hc49e3741, 32'h43f8bd3c},
  {32'h45010706, 32'h443adc4d, 32'hc3811e95},
  {32'hc3a38080, 32'hc35ee978, 32'h44bdedaa},
  {32'h44529e4a, 32'h44466395, 32'hc387f4ac},
  {32'hc46a45df, 32'h42e57712, 32'h44744132},
  {32'h4484585b, 32'h420b1df9, 32'hc4a63c2f},
  {32'hc4407c93, 32'h44052349, 32'h452026f6},
  {32'h43a9ed08, 32'hc362de6a, 32'hc52a2f77},
  {32'h4409d8e0, 32'hc51a9392, 32'hc3c7c9a0},
  {32'hc4eab228, 32'h440e305f, 32'hc33c8f8c},
  {32'h441d3dd5, 32'hc4191239, 32'h434a2be6},
  {32'hc53ae7e2, 32'h43eeaa74, 32'h440bc3eb},
  {32'hc3ce8e8f, 32'hc52baa28, 32'h4390602a},
  {32'hc462e684, 32'h432038f1, 32'hc401b4ec},
  {32'h440b8c0a, 32'h4294e249, 32'h430bdbdb},
  {32'hc40d4510, 32'hc40e6341, 32'hc3ac5143},
  {32'h451335d6, 32'hc356be2d, 32'h4385f2b1},
  {32'hc39695e1, 32'h43628654, 32'h43095ad4},
  {32'hc4214e7b, 32'hc52b8f5b, 32'h431ec30a},
  {32'hc34e0b80, 32'h44a40455, 32'hc340217e},
  {32'hc2dc9e05, 32'h41ce66ae, 32'h4503c1ec},
  {32'hc4f4ee03, 32'h436308c6, 32'hc2a06705},
  {32'h452632c0, 32'h43ad6934, 32'h43f1c203},
  {32'hc52fef75, 32'hc2c5526b, 32'h43247b72},
  {32'h44b22b04, 32'h4445c1a0, 32'h4281ea41},
  {32'hc3cd2ae9, 32'hc27c60ca, 32'hc449fb49},
  {32'h45327fd4, 32'hc40509d8, 32'h42293fe0},
  {32'hc44b8b2c, 32'h451fbbe7, 32'hc430c9bd},
  {32'hc3a616f3, 32'hc3d9dded, 32'h44aaafda},
  {32'hc3f34dc2, 32'hc33d5d27, 32'hc53f0cfc},
  {32'h44d2e021, 32'hc41d8fa3, 32'hc2a78338},
  {32'h449a0adf, 32'h44497819, 32'hc3d6c508},
  {32'h4485e40a, 32'h44912e2c, 32'h43bbd59a},
  {32'hc509a0a1, 32'h437470be, 32'hc4deb6e5},
  {32'h43e6fcd0, 32'h4109f071, 32'h44029643},
  {32'hc40a0682, 32'h44d578df, 32'hc4b2a486},
  {32'hc30f5b2e, 32'hc4acf9d1, 32'h453e5aea},
  {32'h43753f28, 32'hc39c51a2, 32'hc45f1ee7},
  {32'hc3da7d9e, 32'h43f90c72, 32'hc41e1c7c},
  {32'h44737b14, 32'h43be61d6, 32'h4487c549},
  {32'h41916e70, 32'hc3245ce9, 32'hc513be75},
  {32'h40014f00, 32'hc308a88e, 32'h44ae7315},
  {32'hc471870c, 32'h44b59304, 32'hc44020b4},
  {32'h44bf8a6f, 32'hc3910542, 32'h443348ff},
  {32'hc37d8238, 32'hc31b2c1b, 32'h4516780f},
  {32'hc236cac8, 32'hc4878bfa, 32'hc4e4bdc3},
  {32'hc28c2c70, 32'h4404def1, 32'h44412e55},
  {32'h439cfb82, 32'hc22ab52f, 32'h4478e611},
  {32'hc3a861dc, 32'h4512b4b1, 32'h441542e9},
  {32'h4515b8f2, 32'hc388485b, 32'h433f63eb},
  {32'hc22349a4, 32'h43e83bee, 32'hc4f86e0a},
  {32'h4436a91e, 32'hc4c44910, 32'h43fec7c2},
  {32'hc4800407, 32'h433882a3, 32'hc439a911},
  {32'hc4a4c38c, 32'hc3a0376a, 32'h434a5db2},
  {32'hc53f8c48, 32'hc2319394, 32'hc3d1eb32},
  {32'h44808ca5, 32'h441c0638, 32'h43868d8e},
  {32'h40717940, 32'h44bdeb5a, 32'hc36f40ea},
  {32'h3f116000, 32'hc4919eab, 32'h428f5722},
  {32'hc4f06008, 32'h445b9a41, 32'h43b218dd},
  {32'h44b220ba, 32'hc2c7315f, 32'h43a56979},
  {32'hc535bff7, 32'h43ecb3b6, 32'hc414c14b},
  {32'h442401aa, 32'hc5014906, 32'h43e6c43a},
  {32'hc4870aec, 32'hc16fde05, 32'h428773f3},
  {32'h445a4943, 32'hc39ec0f5, 32'hc413c949},
  {32'h41edb108, 32'hc506ff58, 32'h450bbab0},
  {32'hc39698ae, 32'hc2360afb, 32'h448f0b73},
  {32'h43e35cd4, 32'h42a411a5, 32'hc511fe02},
  {32'hc4c9978c, 32'hc3b6a888, 32'h435e3cc5},
  {32'h42693a98, 32'h4434adc2, 32'hc506b263},
  {32'hc4b6a5ca, 32'hc347137a, 32'h44d46861},
  {32'h44513962, 32'h41f17500, 32'h43cb40f8},
  {32'h44a57dc9, 32'h43c46e4b, 32'h43a315fc},
  {32'hc492b2ff, 32'hc4b3bec5, 32'h444a8680},
  {32'h44692f8d, 32'hc3929cf5, 32'hc462343d},
  {32'h440f5b6c, 32'h4313da3c, 32'hc494ad94},
  {32'hc43655fe, 32'hc4681b52, 32'h43eb7bbd},
  {32'h452e6d41, 32'hc19ab47a, 32'h43722db3},
  {32'hc2e1ef50, 32'hc4c5380a, 32'h448cc976},
  {32'hc31488e8, 32'hc2925259, 32'hc539d4be},
  {32'hc4aba62b, 32'hc40d95a9, 32'hc2c0041c},
  {32'h44d17412, 32'h438af6f5, 32'hc3d0fbce},
  {32'hc59aedec, 32'hc303fdbf, 32'h4344bdf4},
  {32'h456f437b, 32'hc1c80558, 32'hc40e37cb},
  {32'hc4f191d2, 32'h42cff74a, 32'hc358c410},
  {32'hc34b87c5, 32'h4583b4d4, 32'h4314318e},
  {32'hc41d589c, 32'hc3ab224a, 32'hc29b3f34},
  {32'h43264c6e, 32'h44b8d8e9, 32'h44049647},
  {32'hc539d4d0, 32'hc3763474, 32'h4387448c},
  {32'h430640d8, 32'h44b3b4fa, 32'hc26f1b6b},
  {32'hc372f8df, 32'h44b7f672, 32'h43a0fe5c},
  {32'h43cb2e27, 32'hc48ac5cf, 32'hc3809638},
  {32'hc364df04, 32'hc3e41c65, 32'h44850994},
  {32'h41e0c4f9, 32'hc2f91b14, 32'hc4b55da2},
  {32'h43a49d05, 32'h4252e5db, 32'h452e499f},
  {32'hc3f6b708, 32'hc29df4e3, 32'hc4e3a8e6},
  {32'h44843fd3, 32'h41a259d0, 32'h42acf725},
  {32'hc3cdcb40, 32'hc368638a, 32'hc4f3c69c},
  {32'h450d542c, 32'h42eebdc3, 32'h4430e301},
  {32'h438019c2, 32'h4489545d, 32'h4252f98a},
  {32'h44cc5ba3, 32'h42facd40, 32'h43f0f002},
  {32'hc3d3ae2a, 32'hc4ef4a56, 32'hc3d09f43},
  {32'h438305f1, 32'h447cb4f7, 32'h4415d1a8},
  {32'hc3d4a67c, 32'h417493a4, 32'hc4cf081e},
  {32'h438a599a, 32'h452ee39a, 32'h44029868},
  {32'hc4961c00, 32'hc3565f7c, 32'hc3966ab3},
  {32'hc32b9930, 32'h446d0c10, 32'h44898b14},
  {32'hc4ac92f2, 32'h4264c3a0, 32'hc3008c4c},
  {32'h456413ee, 32'hc41b6009, 32'h429a8d7b},
  {32'hc576ad3c, 32'hc38bbae6, 32'h43159e85},
  {32'h4491b54d, 32'h44d7bd70, 32'h439940d9},
  {32'hc4cd71c0, 32'h440cf2ac, 32'hc4345f88},
  {32'h44ae5cb9, 32'h44259380, 32'hc3f8fd16},
  {32'hc54d59a5, 32'hc3ad0cdb, 32'h433713fb},
  {32'h42aefe5c, 32'h43f78c6e, 32'hc14535f8},
  {32'hc5315fb4, 32'hc2e66026, 32'hc254ce89},
  {32'h44d251be, 32'h430dca06, 32'h43823db1},
  {32'h44c803bc, 32'hc39d50cc, 32'h41d94a54},
  {32'h43d8cbd0, 32'h451aec59, 32'h4093de93},
  {32'hc4713584, 32'h4449989b, 32'hc2b92297},
  {32'hc46f9658, 32'h444befb0, 32'h434cde6b},
  {32'hc3ab8a6c, 32'hc397ec63, 32'hc504ec05},
  {32'hc447c2dd, 32'h436096b4, 32'h440a81c8},
  {32'h43f4c060, 32'hc4717b77, 32'hc4afdcd0},
  {32'hc4adfab5, 32'h444ec76a, 32'h443a1306},
  {32'hc3d2e9b3, 32'hc3c4b9bc, 32'hc429aa18},
  {32'h42f7053f, 32'hc1e82674, 32'h43c00fae},
  {32'h443e97ad, 32'hc49bfbca, 32'hc3f83cba},
  {32'h42c20f72, 32'h442f6c21, 32'h435b1c8b},
  {32'h43aad8d0, 32'hc4919149, 32'hc2e77a58},
  {32'hc55dd1d4, 32'hc2c4e22c, 32'h434ac700},
  {32'hc237fe40, 32'h43979447, 32'hc4d8bbef},
  {32'hc2ddde12, 32'hc3b01652, 32'h45221e46},
  {32'h44589674, 32'hc41aad48, 32'hc4bbd6de},
  {32'h43d7e6c0, 32'h4296916c, 32'h44c9ce89},
  {32'h450bae5b, 32'hc4b4347c, 32'hc358fef5},
  {32'hc513b2c4, 32'h443bd16c, 32'hc33a51cd},
  {32'h4435773e, 32'h4384eb86, 32'hc32228a2},
  {32'hc38b3af1, 32'h452b07b1, 32'hc369b985},
  {32'h4542e480, 32'h43de6187, 32'h4349fe9d},
  {32'h421c4f28, 32'h44a7c5a9, 32'h415d97d5},
  {32'h43b9b3d0, 32'h3f570bb0, 32'hc1547a60},
  {32'hc58dd3f4, 32'h44367e31, 32'hc27b0e37},
  {32'h450ace8e, 32'hc1deeece, 32'h41bf26b4},
  {32'hc46c0b7c, 32'h44247f44, 32'h441e75e5},
  {32'hc52b9aec, 32'hc3d24d42, 32'hc41b9b36},
  {32'h4546528d, 32'h438bb428, 32'h4346c4c2},
  {32'hc44bc24e, 32'hc372858c, 32'h431a1b35},
  {32'h44086024, 32'hc3b4bf09, 32'h441c69a5},
  {32'hc3bded54, 32'h451eb99b, 32'h43ef6150},
  {32'hc426726c, 32'hc37f64f3, 32'h3f847ee5},
  {32'hc50c3416, 32'h444b120f, 32'hc38d4ef2},
  {32'h4429f9cb, 32'hc4c82993, 32'hc38fdbff},
  {32'h44dde8c2, 32'hc3e9bd7d, 32'hc303276e},
  {32'h44bfa4cc, 32'h437c97e5, 32'h4351377d},
  {32'hc4566c40, 32'h43e23c26, 32'hc42d7b0c},
  {32'h443c8d80, 32'hc37880d9, 32'hc39b767c},
  {32'hc3b8ce8c, 32'h44972be6, 32'h4485e432},
  {32'h443ff448, 32'hc413790a, 32'hc4056bf2},
  {32'h41cf7c02, 32'hc3024887, 32'h42dde82e},
  {32'hc2d894dd, 32'h43b72490, 32'hc5404345},
  {32'hc1249ff0, 32'h42aaaf47, 32'h44e657d2},
  {32'hc4c383bf, 32'hc305f22a, 32'hc3d43c42},
  {32'hc5939905, 32'h3f0d6048, 32'h429cd7b8},
  {32'h4381c004, 32'hc2d1ff51, 32'hc4af8d11},
  {32'hc468a71c, 32'hc3c5467e, 32'h441ec4e5},
  {32'h45073a23, 32'hc2c1f739, 32'hc40e138e},
  {32'hc44700c4, 32'h44e44240, 32'hc32a32aa},
  {32'hc31b92b0, 32'h44051909, 32'hc4a42ce0},
  {32'hc48fabe5, 32'h44d55310, 32'h44692f25},
  {32'h42118b9a, 32'hc52809d2, 32'hc412d741},
  {32'h4455c680, 32'h41c52a61, 32'h42cfc25b},
  {32'hc4b574a0, 32'hc19a02e2, 32'h43d4eb22},
  {32'h445235af, 32'h441eaef9, 32'hc447c55c},
  {32'hc4c698cf, 32'hc4a598b4, 32'hc15f2843},
  {32'h44236fb1, 32'h427dea08, 32'h4401f630},
  {32'hc4ef50b7, 32'h42198c2a, 32'h4322df5a},
  {32'h43ec1658, 32'h457f51d8, 32'h429034d6},
  {32'hc5794d44, 32'hc3e3c5a4, 32'h44031038},
  {32'h43beb604, 32'h44c8b7ad, 32'hc329af17},
  {32'hc42c7d4c, 32'hc40040ba, 32'h433a99a0},
  {32'h441ee35a, 32'h4409227a, 32'h432d127d},
  {32'hc4c2ad48, 32'h421bad05, 32'hc21f674f},
  {32'h45369832, 32'hc2dc075d, 32'h440da8f3},
  {32'hc201371c, 32'hc54f38d0, 32'h436702a4},
  {32'hc32cc08c, 32'h44c47b21, 32'h43fa2436},
  {32'h43275bc2, 32'h428c4d7a, 32'hc5213e34},
  {32'h450e1f44, 32'hc2c4e992, 32'h42388aa9},
  {32'hc380d356, 32'hc4005802, 32'hc2903e7f},
  {32'h454988ae, 32'hc2ef6c35, 32'h43cefad9},
  {32'hc54f0024, 32'hc3221074, 32'hc2c9880c},
  {32'h452c3c6c, 32'h430531b1, 32'hc41f0f0e},
  {32'hc3c190a6, 32'hc416f779, 32'hc4f0b847},
  {32'h450c0c9f, 32'h43819023, 32'hc33045b8},
  {32'hc49a62aa, 32'hc412a8da, 32'hc3601556},
  {32'h44ee71ed, 32'h438cf7af, 32'h43d7a909},
  {32'hc4d55801, 32'hc3c38047, 32'hc398f15e},
  {32'hc4b71816, 32'h43d7c6ec, 32'hc30fca19},
  {32'h4511e2ae, 32'hc441eb6d, 32'hc2ab7af8},
  {32'hc49718ca, 32'hc4584289, 32'hc34ba524},
  {32'h44e031f8, 32'h449b888d, 32'h43e30ee1},
  {32'hc53f54e8, 32'h4408d896, 32'h43999404},
  {32'h44334fa2, 32'h450ddea0, 32'h43b52111},
  {32'hc452571b, 32'hc40a05a4, 32'h42b1cdc9},
  {32'hc4222708, 32'hc3643d2f, 32'h4259a38c},
  {32'hc57a3d0a, 32'hc33c337c, 32'h43294793},
  {32'hc3803962, 32'h42df4af7, 32'h4400a504},
  {32'h435bc6df, 32'hc49a9e63, 32'h44cc1f44},
  {32'h45154410, 32'h4350e337, 32'h43ce67fa},
  {32'hc2dec470, 32'hc48ce161, 32'h44252524},
  {32'hc2b8205e, 32'h44e34d66, 32'h435f3acd},
  {32'hc4ae874f, 32'hc409a837, 32'h440d7206},
  {32'h425f1550, 32'h4255db40, 32'hc4c8891f},
  {32'h432b19c6, 32'h4298ec0f, 32'h435ee70d},
  {32'h444adfb0, 32'hc3d52a8c, 32'hc4845408},
  {32'hc50c180e, 32'h4243fa32, 32'h43d2f039},
  {32'hc319f2fc, 32'h446b943c, 32'h40e755b8},
  {32'hc4dc9096, 32'hc42b4690, 32'h44bb30a4},
  {32'h4561f792, 32'h43cb7093, 32'hc35ceb3f},
  {32'h44d076ee, 32'h439314ff, 32'h436a86c8},
  {32'hc38c6bad, 32'hc4048e64, 32'hc5117965},
  {32'h4398a2c6, 32'hc34954df, 32'h4502bd0c},
  {32'hc497f187, 32'h4396c666, 32'hc3a4d073},
  {32'hc57548e7, 32'h43bfc406, 32'h433badc2},
  {32'h42d991c0, 32'hc43a346f, 32'hc533715c},
  {32'h4416f02c, 32'hc51c0378, 32'hc37cb5fe},
  {32'hc3e45eec, 32'h44c7a2e5, 32'h443c2b6b},
  {32'h40202600, 32'hc301ff17, 32'hc32f8883},
  {32'hc42281de, 32'h44d5918c, 32'hc3cab143},
  {32'h443af044, 32'hc4b2c583, 32'h42ce2635},
  {32'h445dd070, 32'h42d8bd44, 32'hc39a499a},
  {32'h44d2a761, 32'h4440f99e, 32'hc2444c66},
  {32'hc411df45, 32'h43d6800b, 32'h42740205},
  {32'hc4a6da67, 32'hc3b894ae, 32'h43a946ef},
  {32'hc4c2a8a3, 32'h441c37bf, 32'hc414ba9f},
  {32'h44585fd4, 32'h44173fe0, 32'hc36b0b62},
  {32'hc480d63c, 32'h43f97827, 32'hc39736cc},
  {32'h42a1c7ac, 32'h4178184b, 32'h45451746},
  {32'hc41660a8, 32'h445f8080, 32'hc44f18d9},
  {32'h4446f99c, 32'hc3df75c3, 32'h43bebeb3},
  {32'hc468c04a, 32'h43aec421, 32'hc3a9b959},
  {32'h45137896, 32'hc3e8c92b, 32'hc23a25ba},
  {32'hc5324516, 32'hc394a744, 32'hc38a3351},
  {32'h450a0aad, 32'hc43b5131, 32'hc12a724a},
  {32'hc3d94d9c, 32'h451afb2f, 32'hc44d57b8},
  {32'hc30e868e, 32'hc3c85b2e, 32'h44493384},
  {32'hc4be88de, 32'h44d751f3, 32'hc29791b8},
  {32'h447f5b48, 32'hc400e828, 32'h448022b8},
  {32'h42e04568, 32'hc2b5cfbd, 32'hc4cce948},
  {32'h457768fa, 32'h44076ced, 32'h43c9c193},
  {32'hc41f23ed, 32'h4390786e, 32'hc493cfa0},
  {32'h44b6cf07, 32'h43247b94, 32'h41af6271},
  {32'h43fd7a3d, 32'h44a0b21a, 32'hc4cfb134},
  {32'h43f61fd0, 32'h436a3ba2, 32'h44b0902a},
  {32'hc4e24383, 32'hc3ca78fe, 32'h4276bd0c},
  {32'h44f48e2f, 32'hc2afb5c6, 32'h434c76ea},
  {32'h44c59044, 32'hc3796d82, 32'h44a981b6},
  {32'hc513030a, 32'h4340e1df, 32'hc3bfdf92},
  {32'hc3f2bf74, 32'h43e1240c, 32'h44b9a396},
  {32'hc4d0536d, 32'h4482ca5f, 32'hc3168f0e},
  {32'h43513c58, 32'hc4b53565, 32'h4401a2f3},
  {32'h4485a022, 32'h44b34150, 32'h447388ac},
  {32'hc3875082, 32'hc47e129d, 32'hc427dc40},
  {32'hc3d795ff, 32'hc49b74bb, 32'h4445d291},
  {32'h43affd53, 32'hc3953e8f, 32'h45005696},
  {32'hc54f6ab2, 32'hc3bf2c54, 32'hc20a1981},
  {32'h4065e180, 32'hc491a416, 32'h43614fa5},
  {32'h44842f3e, 32'hc2f7913f, 32'h43146bee},
  {32'h4413c18e, 32'hc4f1cfd7, 32'h42ee5701},
  {32'h42f3c994, 32'h44bbddc9, 32'hc41d4a70},
  {32'h44a8d613, 32'hc363e560, 32'h44135f6f},
  {32'hc58dd6f8, 32'hc2ead08d, 32'hc2481484},
  {32'h44f14b8b, 32'h44745bc1, 32'hc34e5cce},
  {32'h449c5c2c, 32'h44140830, 32'h438a499d},
  {32'h45287710, 32'hc3c752bc, 32'hc398d3d1},
  {32'hc3cdf33c, 32'h45030266, 32'hc3067461},
  {32'h452f9dec, 32'h4387857e, 32'h4364b150},
  {32'hc43ca43c, 32'h454567ba, 32'h43e9e1e6},
  {32'h44c06cf7, 32'hc44b57d4, 32'hc2b7d05e},
  {32'h445b2c90, 32'h4419f03d, 32'h43472187},
  {32'h43ad0f39, 32'h44f9d439, 32'hc4894baa},
  {32'hc4321712, 32'hc47e5390, 32'h44992482},
  {32'hc38337ce, 32'hc43e66c7, 32'h44479316},
  {32'h44d4a384, 32'h436af88f, 32'hc227369a},
  {32'h4499fc20, 32'hc40b1f82, 32'h435ec55c},
  {32'hc30ba0cc, 32'h450b3a57, 32'h42cc5d28},
  {32'h4374ed46, 32'hc347b12a, 32'h4537dd86},
  {32'h439f149f, 32'h4468053e, 32'h418c5c8c},
  {32'h436b5b53, 32'h438ff002, 32'hc3d7a8eb},
  {32'hc4f79f2e, 32'h445f09e4, 32'h4423b001},
  {32'h43eaa1fc, 32'hbf2c3ab0, 32'hc4bf3841},
  {32'h446db34e, 32'h43ebb787, 32'hc43ccda3},
  {32'hc51f2682, 32'hc39e80e0, 32'h42a7671c},
  {32'hc4ce9f82, 32'h43a0a315, 32'hc34313e4},
  {32'hc424abc1, 32'hc410135d, 32'h44daa806},
  {32'hc41c39d3, 32'hc3f8e75a, 32'hc525ed63},
  {32'hc3de9192, 32'hc4a471d2, 32'h43fcffb0},
  {32'h45336a5d, 32'hc3e64bf8, 32'h43574d2b},
  {32'hc5829496, 32'hc21e190d, 32'h42ed8b4a},
  {32'h4518c6e8, 32'h44203073, 32'hc3726376},
  {32'hc3194620, 32'hc3b4907c, 32'h4431fc89},
  {32'h450eaea6, 32'h4219a336, 32'h427ecb66},
  {32'hc549e5c8, 32'h432708c2, 32'h43a97223},
  {32'h444eff9c, 32'h448aa4fe, 32'hc3957274},
  {32'hc585af98, 32'hc347e98b, 32'hc397701f},
  {32'h42862f6d, 32'h44607a74, 32'h4352cfa6},
  {32'hc3f21c70, 32'h43a1808a, 32'h4459b32f},
  {32'hc40ee2d3, 32'h442fe79f, 32'hc46d3204},
  {32'h435c88c5, 32'h445c9a1b, 32'h448a56fe},
  {32'h44ec9d27, 32'hc2d3a5d1, 32'hc3c63d1a},
  {32'h440c7b7b, 32'h448f6a5e, 32'h441df8f1},
  {32'h43198a40, 32'hc493a9e4, 32'hc436a7a7},
  {32'h446605b5, 32'hc3570a7b, 32'h434afb8c},
  {32'hc4f091db, 32'hc40b5366, 32'hc47b83ef},
  {32'h44f30416, 32'h4398d6bd, 32'h44327263},
  {32'hc48ffe54, 32'hc32b37d3, 32'h4282f692},
  {32'hc3485754, 32'hc38c3771, 32'h43f31ade},
  {32'hc4892ca8, 32'h44064baa, 32'hc4c0316f},
  {32'hc4aee80a, 32'h43a1134e, 32'h42908e58},
  {32'h432ef674, 32'hc44eba3b, 32'hc4c6e601},
  {32'h44effc82, 32'h439058b3, 32'hc2b44f74},
  {32'h44d4c6e6, 32'hc4083ac5, 32'hc38d6df5},
  {32'hbedb36a0, 32'h4415b312, 32'h455412dc},
  {32'hc4c2d581, 32'h429afd58, 32'h4021a1fc},
  {32'hc419bd0e, 32'h440ed0b6, 32'hc2975aaa},
  {32'hc3aa74fa, 32'hc545420f, 32'hc41cbf50},
  {32'hc2aa0c80, 32'h4497a2fa, 32'h42f88d3a},
  {32'h4435d6e4, 32'h426eff15, 32'h42e36149},
  {32'h44500844, 32'h44922d2e, 32'hc4296bc9},
  {32'hc49dfc0c, 32'hc4910848, 32'hc2fb7369},
  {32'hc4cf24f3, 32'h42e1c7c3, 32'h41e8dd0c},
  {32'hc4523974, 32'h430327dd, 32'hc39a9dd0},
  {32'h44c25520, 32'hc2a3e738, 32'h42cb9b34},
  {32'h4383ebb3, 32'h44d4e1a7, 32'hc4d549e8},
  {32'hc3cbb580, 32'h44c6750f, 32'h444525c5},
  {32'hc3fb3bd3, 32'hc476241f, 32'hc41265a7},
  {32'hc50c9208, 32'h449164dc, 32'h4402bc81},
  {32'hc2ea9220, 32'hc441a5ce, 32'hc4c3ce06},
  {32'h4485b9fe, 32'h4485996c, 32'h43c8b4b0},
  {32'h4450d45c, 32'hc3e6570a, 32'hc43b959e},
  {32'hc4c8d088, 32'h42e5e13f, 32'h43a2e187},
  {32'h44accf36, 32'h43012cfa, 32'hc45fa012},
  {32'hc42f3a8c, 32'h4447db6e, 32'h448c9001},
  {32'hc2c603db, 32'h450e96e9, 32'hc4da5cbd},
  {32'h41268448, 32'hc42072f4, 32'h449df8d5},
  {32'h44b14f06, 32'hc4afcef0, 32'h433cd42f},
  {32'hc3df3ab4, 32'h43869c0d, 32'h4328bf10},
  {32'hc3a0e258, 32'hc2cc247a, 32'hc3b0d8d5},
  {32'hc3c3bd16, 32'h43a03a39, 32'h45702942},
  {32'h4491e20d, 32'h43e20353, 32'hc49edf7b},
  {32'h447998e2, 32'h43af0963, 32'hc337a58d},
  {32'h442262de, 32'hc54787ce, 32'h43d862c2},
  {32'hc40e611c, 32'h44c8af13, 32'h4290d61f},
  {32'hc39e8c2d, 32'hc38d15d8, 32'h43411dbe},
  {32'hc3a88d68, 32'h446bd8b7, 32'hc3f0b7f4},
  {32'h452b0b76, 32'hc39a1289, 32'h43461cc9},
  {32'h43f8c5fa, 32'h4496ef9a, 32'hc2e58796},
  {32'h4551ae9f, 32'hc2cbb804, 32'h43bf2e54},
  {32'hc5276a44, 32'hc420fd59, 32'hc2dba2a4},
  {32'h44977e95, 32'hc3488eb3, 32'hc3c53dc2},
  {32'h4158a260, 32'h4385b877, 32'hc26e5751},
  {32'hc3fa8c08, 32'hc283f8c3, 32'hc480797d},
  {32'h45288b6d, 32'hc208f84f, 32'h43c38b79},
  {32'hc50934ea, 32'hc383daa7, 32'hc2fbbb21},
  {32'hc33b9a50, 32'hc55e838e, 32'h42a246ae},
  {32'hc55de776, 32'hc1d0d24c, 32'hc1eb087e},
  {32'h4343e434, 32'h41b7805e, 32'hc3a9f96c},
  {32'hc47b1d53, 32'h44c38e78, 32'h4281fed1},
  {32'h445a4a0b, 32'hc4f075ad, 32'hc3deaeea},
  {32'h42c7d898, 32'h438d6b99, 32'hc429571d},
  {32'h4388e8a8, 32'hc38822e2, 32'h43e0b248},
  {32'hc4a280b6, 32'h4410744d, 32'hc4c3a749},
  {32'h429436fc, 32'hc309d81a, 32'hc4bd16b5},
  {32'hc15f75f0, 32'h4500c6c0, 32'h44054e2e},
  {32'hc3497c8a, 32'hc37e500e, 32'hc55b7aac},
  {32'h443a8283, 32'h43b0e8bd, 32'h4366b816},
  {32'hc392fa46, 32'hc49b7029, 32'hc3a425f0},
  {32'hc3aec492, 32'hc17001aa, 32'h44e7e100},
  {32'h43df79c3, 32'hc386c270, 32'hc254642d},
  {32'hc48e93ab, 32'hc4d735a4, 32'h44e6e2a4},
  {32'h448f5e11, 32'hc41d2c87, 32'hc4b5e795},
  {32'h43acf3c4, 32'h448126bf, 32'h4416bd6e},
  {32'h44546ca0, 32'hc478e1f8, 32'h42d7bdc2},
  {32'hc496c8a4, 32'h44c8dcf6, 32'hc369ba33},
  {32'h43ed6e6c, 32'hc499d32e, 32'hc377da3d},
  {32'hc4be51e2, 32'h4412f980, 32'h44c064ff},
  {32'hc2434850, 32'hc4db9b07, 32'hc43413ed},
  {32'h44a6c8c4, 32'hc340330c, 32'hc2c53734},
  {32'hc5795ee4, 32'hc1ff9b00, 32'h440932b0},
  {32'h439d9606, 32'h44424171, 32'hc46145e7},
  {32'hc418eca0, 32'hc4d5d86a, 32'h4343450e},
  {32'h448b9c61, 32'h444596a5, 32'hc35db53b},
  {32'h435e878c, 32'hc45d43e1, 32'hc3c45b79},
  {32'hc38ef0de, 32'h454afc13, 32'h437f4d18},
  {32'hc50e5f70, 32'hc454f35e, 32'h4437b958},
  {32'hc48c6445, 32'h43efb3ef, 32'h43063918},
  {32'hc451f660, 32'hc3d36d51, 32'h449dc873},
  {32'h440bac6c, 32'h43a0a360, 32'hc3b953cd},
  {32'h4446f24b, 32'hc2b41592, 32'h4387d02b},
  {32'h44565cae, 32'h42d6594d, 32'h443e4e7f},
  {32'hc4e9e9fe, 32'hc3e6b52d, 32'hc283be0a},
  {32'h44fb8fef, 32'hc3a4666f, 32'hc28165d2},
  {32'hc37afc64, 32'hc4f25879, 32'hc24f664a},
  {32'h442ac59c, 32'h44cd59f9, 32'h438867e7},
  {32'hc44e14ae, 32'hc40a6bb9, 32'h43ffe9ff},
  {32'h44ed0559, 32'h445f130f, 32'h442c1650},
  {32'hc52ee203, 32'hc29a376a, 32'hc3a4313a},
  {32'hc4c34e44, 32'h422a6021, 32'h413fa66e},
  {32'hc5183c0d, 32'h43ea954d, 32'hc447ef1e},
  {32'h443eff6a, 32'h44aa8e1c, 32'h43e7873f},
  {32'hc48c4292, 32'hc3087a4f, 32'h42eabe07},
  {32'hc321e42e, 32'h4488d38c, 32'h443afc66},
  {32'hc4c13e00, 32'h434a6178, 32'hc4bec252},
  {32'h446d2e5b, 32'h447ea8bb, 32'h43cacef5},
  {32'hc3899685, 32'h42ea3f40, 32'hc419b763},
  {32'hc4ab6090, 32'hc4020e59, 32'hc2a40b8c},
  {32'h4422dc23, 32'h4505c4e9, 32'hc1a60bb8},
  {32'hc4d16180, 32'h43c3966b, 32'h440595ce},
  {32'h43f09f31, 32'h450d4668, 32'hc3a08a9a},
  {32'hc542df21, 32'hc441507c, 32'hc1c54445},
  {32'h45462c5e, 32'hc34e2f2b, 32'hc41421b1},
  {32'hc4467dfc, 32'hc31258d7, 32'hc387ef06},
  {32'h4414756a, 32'hc3ba19ed, 32'hc3662f3f},
  {32'h430cc711, 32'h435d4e6d, 32'h4457a88a},
  {32'h44971d24, 32'h4425f55f, 32'hc38f8fd5},
  {32'hc5358036, 32'h3ffe1640, 32'hc2f94884},
  {32'hc4a813be, 32'h43e005ae, 32'hc36a9d1b},
  {32'hc44434c6, 32'hc492ec08, 32'h42b95e50},
  {32'h40c54b70, 32'h44a1e87b, 32'h443bf3f7},
  {32'h448ce148, 32'hc2407e61, 32'h42c5f889},
  {32'h4333b8b4, 32'h42903ac7, 32'hc523b78f},
  {32'hc513d9ad, 32'h4102f8a7, 32'h417f0ff5},
  {32'h43b2391d, 32'h446e1bfe, 32'h430d518c},
  {32'hc3940b18, 32'hc4e2800a, 32'h4426ad53},
  {32'h44aff8ae, 32'h44c994be, 32'hc427c579},
  {32'hc4879020, 32'h434c7e3e, 32'h43cc2ca4},
  {32'h42f639cc, 32'h452ecce7, 32'h43064ff6},
  {32'hc500a8b9, 32'h43c3372c, 32'h42cc3006},
  {32'hc36cc167, 32'hc2377f7c, 32'hc3243e86},
  {32'hc40d2bd8, 32'h432a3d1e, 32'h44d3d648},
  {32'h4434b0bb, 32'hc4264271, 32'hc4ddd980},
  {32'h42b2aa80, 32'hc4d57e70, 32'hc27340da},
  {32'hc3d18b8c, 32'h4449fb2d, 32'h4389899b},
  {32'hc4cc1808, 32'hc3d346e1, 32'h4309ccb9},
  {32'hc45ac19a, 32'h43820694, 32'hc389d1f1},
  {32'h44b29d14, 32'hc32b13fa, 32'h44004498},
  {32'h44ce6734, 32'h43c9d458, 32'h42afb7b2},
  {32'h4522c25b, 32'h43c66d92, 32'hc3ad658f},
  {32'hc4dc8fc0, 32'h445ad59c, 32'h44833537},
  {32'h4459c2f6, 32'hc21f3d7c, 32'h40e883e8},
  {32'hc3c45f6c, 32'h442a093b, 32'hc4bb68cb},
  {32'hc28d4808, 32'hc55341fa, 32'h4404a605},
  {32'hc3bec7eb, 32'h4430634a, 32'hc31d98ec},
  {32'h44ec03ea, 32'h43b9795a, 32'h448ec8e9},
  {32'hc4e3e42d, 32'h445762a3, 32'hc453e7c7},
  {32'h418d9eec, 32'hc428d474, 32'h440281b1},
  {32'hc53c41fc, 32'hc395d475, 32'h440499a3},
  {32'h44a43af8, 32'hc3cd008a, 32'h43184424},
  {32'hc2958ee0, 32'hc3c2053c, 32'hc4871348},
  {32'h43a07092, 32'hc5270cd5, 32'hbeb36d40},
  {32'hc49c32fc, 32'h443f14ff, 32'hc43f7dbc},
  {32'h44b2ef03, 32'hc388d8b7, 32'hc308e1f0},
  {32'hc356b118, 32'hc23c2493, 32'hc40fe4aa},
  {32'h44b8815e, 32'hc2d74744, 32'h43da161e},
  {32'h443f30f3, 32'h4006f8fa, 32'hc3bd6f56},
  {32'h451b4fbf, 32'h434b479b, 32'h43acb991},
  {32'hc5405f75, 32'h43240018, 32'hc3c8486b},
  {32'hc401decd, 32'hc40378b3, 32'h43deffa2},
  {32'hc46dfc04, 32'hc460f83b, 32'hc43a9b72},
  {32'h43b296f1, 32'hc4d4509c, 32'h4506eaa9},
  {32'h44662f6e, 32'h43d04c57, 32'hc3a79ee9},
  {32'hc41cc48c, 32'h439ff82d, 32'hc43f46fc},
  {32'h42a31da2, 32'h43bdf9ad, 32'h4518f3c6},
  {32'hc40027b1, 32'h43219a5d, 32'hc3ca7bb5},
  {32'hc3bd0024, 32'hc30e1bac, 32'h43a04643},
  {32'hc38b9e30, 32'h45514a96, 32'hc32c7e80},
  {32'hc082c100, 32'h42ad2ee6, 32'h453f9961},
  {32'hc3868892, 32'h44d66030, 32'h451da54b},
  {32'hc4c5a6e9, 32'hc4750211, 32'hc43018a2},
  {32'h44f80e58, 32'h41e5771f, 32'hc3cf5abc},
  {32'hc4c49067, 32'h4204a7c2, 32'h43a8a561},
  {32'hc1cb7c80, 32'h44a576e4, 32'hc44e4de9},
  {32'h4404b7f0, 32'hc4ef1d21, 32'h4383e916},
  {32'h44949c82, 32'h44246de0, 32'hc38e67d8},
  {32'h450af026, 32'hc40abbce, 32'hc310b896},
  {32'hc44b1d25, 32'hc21e056d, 32'hc469635f},
  {32'h45813712, 32'hc39adac3, 32'hc39ebeb0},
  {32'hc5129240, 32'h43bdb747, 32'h43773370},
  {32'hc3d9edd0, 32'h440a4050, 32'h43e63825},
  {32'h41fae1fb, 32'h44de9a96, 32'hc36eaafb},
  {32'h44c409f0, 32'hc4a08bd5, 32'h444c9740},
  {32'hc51f60f0, 32'h440b1e85, 32'hc30f0f78},
  {32'hc4b98f9d, 32'hc3a8a364, 32'hc3b18787},
  {32'hc4765d1c, 32'h44b9a238, 32'hc3730b14},
  {32'h43911118, 32'hc50dae1a, 32'hc1dc2625},
  {32'h43d4210b, 32'hc3c80eb6, 32'h4448b5e1},
  {32'h40b50e80, 32'hc41b0ae4, 32'hc48378d6},
  {32'hc470dd9e, 32'hc25a7eb2, 32'h441c952a},
  {32'hc50ff664, 32'hc4362db8, 32'h43921d3e},
  {32'h44c633db, 32'h43e3981c, 32'h429e4238},
  {32'hc523bac8, 32'h43575b37, 32'hc2c70aed},
  {32'h44222845, 32'h43e99166, 32'hc4ab4acf},
  {32'hc4344bcb, 32'hc33622cb, 32'h44e5b2dc},
  {32'h4485299d, 32'h44310c1c, 32'h43ad7654},
  {32'hc3867e4e, 32'hc35c592e, 32'hc485287b},
  {32'hbf763018, 32'h43e398a3, 32'h44fd288f},
  {32'hc2e96f7f, 32'hc4ead2af, 32'hc4dd5b64},
  {32'h440e04d0, 32'h44531fb4, 32'hc34c8394},
  {32'hc4223d44, 32'hc4ae0e14, 32'hc1d9c5ed},
  {32'hc40db298, 32'h43b01a68, 32'hc485a23b},
  {32'h4304bdae, 32'h439a9c1c, 32'h4452fb02},
  {32'h43f96945, 32'hc1d17211, 32'hc50992bc},
  {32'hc3aa4a4e, 32'hc4dd3b6d, 32'h4298421c},
  {32'h455e87de, 32'hc3601d31, 32'h430c2154},
  {32'hc4920672, 32'h440c131c, 32'h43936fb2},
  {32'hc392e4fc, 32'h43a03bc0, 32'hc3ea5583},
  {32'hc497963d, 32'hc222a2c6, 32'hc3449eae},
  {32'hc33188ba, 32'h4514a34e, 32'h420e6bae},
  {32'h440382c5, 32'hc41b1d64, 32'h43960830},
  {32'h44a7b7de, 32'h43af24f6, 32'hc26cb27f},
  {32'hc4ac064e, 32'hc31af583, 32'h436b41d2},
  {32'h44bda82a, 32'hc2a7fd2e, 32'h4309ce1e},
  {32'hc38170cc, 32'hc32b1409, 32'h440a2580},
  {32'h4334e196, 32'h43305144, 32'hc4d47e3d},
  {32'h4461d72c, 32'hc449df22, 32'h4454c5be},
  {32'h433e7e79, 32'hc41c9fe8, 32'h427c58f9},
  {32'h450a4c1b, 32'h43833982, 32'h42886667},
  {32'h432c06f1, 32'hc400af2e, 32'hc4e4308f},
  {32'hc33934fc, 32'h445dc6df, 32'h438adcec},
  {32'hc4d09f1b, 32'h42867fad, 32'hc3d6162f},
  {32'h4508ebc9, 32'h4412c1ad, 32'h443bc493},
  {32'h43766ad4, 32'hc4675da5, 32'h428779db},
  {32'h43d222c2, 32'h44c10cb9, 32'h421a5ec9},
  {32'hc4244492, 32'h4365f722, 32'hc4b7497b},
  {32'h44a6e4c3, 32'h44085eb0, 32'hc3232116},
  {32'hc425207c, 32'hc457cf58, 32'hc3cde3d2},
  {32'h439f1253, 32'h453e1cf1, 32'h43c206e4},
  {32'h43849710, 32'hc2865be2, 32'hc4b69b19},
  {32'h43beb944, 32'h42a05712, 32'h45411a17},
  {32'hc3cb5bd1, 32'hc451191a, 32'hc579bbad},
  {32'h42efa67e, 32'h44f38c61, 32'h4410cbd1},
  {32'hc49faf93, 32'hc5066d0a, 32'h42b14f2f},
  {32'h44f67524, 32'h44cf59d6, 32'h431de349},
  {32'h448d5048, 32'hc3c5354e, 32'hc3ca2761},
  {32'h4386b9ae, 32'h44bab54d, 32'h41c07eba},
  {32'hc2cc1600, 32'hc482e44f, 32'hc3fed40d},
  {32'h45294ee3, 32'h42c3de2a, 32'h43daa86c},
  {32'hc531cffb, 32'hc37af59b, 32'h435eb733},
  {32'h450abe0c, 32'hc488d749, 32'hc2f85816},
  {32'hc3c94b45, 32'h447d3972, 32'hc41cd83b},
  {32'h438c0771, 32'hc49db4ba, 32'h44bbfacf},
  {32'hc3cd4289, 32'h43426ef4, 32'hc4278983},
  {32'h43f33288, 32'h440f4fad, 32'h45263fd6},
  {32'h44e1564a, 32'hc416a536, 32'h43f5fcf7},
  {32'hc17c7cf0, 32'h4449e8ab, 32'h430994d6},
  {32'h43b2a6c8, 32'hc46fc838, 32'hc4c6b7a0},
  {32'hc52c91a6, 32'h43c4dafb, 32'h4402a0e4},
  {32'hc39e9258, 32'hc4342791, 32'hc35e1f70},
  {32'hc354e5c0, 32'hc2b6b2fc, 32'h4496120d},
  {32'hc3c7a0c4, 32'hc3985896, 32'hc4063b4e},
  {32'h43e2bb21, 32'hc3a9c45e, 32'h446eb9ec},
  {32'h43be3765, 32'h4315f35e, 32'hc5234bce},
  {32'hc26fa91e, 32'h43a0608a, 32'h4310784d},
  {32'h45093d32, 32'h44049957, 32'hc2856d9c},
  {32'hc30cf007, 32'h445a6da6, 32'h45657f6d},
  {32'h44cc0e10, 32'hc457c4c3, 32'hc3ecf917},
  {32'hc3bdfb54, 32'h440ecfdb, 32'h43c82c8d},
  {32'h452e6b73, 32'hc43622ae, 32'hc2f8b50a},
  {32'hc4d389b8, 32'h44a4eacb, 32'h43cd6ada},
  {32'h44893978, 32'hc40af843, 32'h439ddedd},
  {32'h43768ab6, 32'h44eb80f2, 32'h444a4480},
  {32'h453db21c, 32'hc407b0df, 32'h420a4e21},
  {32'hc409c583, 32'h42b10db3, 32'h44518953},
  {32'h450787a5, 32'h437ebe1c, 32'hc3623625},
  {32'hc58a04ba, 32'hc329160c, 32'h435730c4},
  {32'h444568db, 32'hc23798a1, 32'hc38af40d},
  {32'h44ed0954, 32'hc39f02f5, 32'hc2d6c0dd},
  {32'hc512c862, 32'h433be34c, 32'hc3224143},
  {32'h44b859c4, 32'h42f0a05f, 32'h44890704},
  {32'hc336295d, 32'h43827146, 32'hc3b071ae},
  {32'h44f7d373, 32'hc4a47bbe, 32'h4072ae14},
  {32'hc426c370, 32'hc2d10e24, 32'hc32cc773},
  {32'hc4379002, 32'hc41219be, 32'h42136864},
  {32'hc398d230, 32'h45523609, 32'hc34a3ec3},
  {32'h450d55cd, 32'hc47cb58b, 32'hc36abf2d},
  {32'hc512e284, 32'hc269b3b9, 32'h4362de4c},
  {32'h4399a86a, 32'hc45cb07b, 32'h4534b7a6},
  {32'hc43988e9, 32'hc333180b, 32'hc49ecd62},
  {32'h4422ac60, 32'hc39bb631, 32'hc318d231},
  {32'hc4a5b3a5, 32'h4384cf4c, 32'h43949434},
  {32'h440cd9aa, 32'hc2d13eea, 32'hc4d0d19b},
  {32'h44a806d1, 32'h4093c358, 32'h43556f1e},
  {32'h4107219d, 32'hc5255e18, 32'h42f7d29e},
  {32'hc4eaa86e, 32'h43618fcd, 32'h436fab82},
  {32'hc4fa7dbf, 32'hc34b2e52, 32'h42fb67cd},
  {32'hc59190a2, 32'h4393d348, 32'h438be6ce},
  {32'h44dcbe3f, 32'hc487eaed, 32'hc4a3a466},
  {32'hc38d4450, 32'h43ebfd17, 32'h42d7071b},
  {32'hc2bb3038, 32'hc52202b4, 32'h42e9fcdc},
  {32'hc40db3ac, 32'h43196265, 32'h44d90dcc},
  {32'h44e76340, 32'h431831dc, 32'h429e1eec},
  {32'hc442df24, 32'h443f3d3f, 32'h448caa8d},
  {32'h427cdf00, 32'hc4a9955a, 32'hc4d55e89},
  {32'h4552775c, 32'h4292297e, 32'hc3783145},
  {32'hc4d7544d, 32'hc375d232, 32'h44e1c803},
  {32'h44a4ae18, 32'h43ae3b57, 32'hc315c995},
  {32'hc30a2506, 32'hc38dabdc, 32'h43956d64},
  {32'h44ef9f40, 32'h43254daa, 32'h43f2ff64},
  {32'hc508ea24, 32'hc1f78090, 32'hc30aeaeb},
  {32'h433237c9, 32'h4527e2eb, 32'hc328841a},
  {32'hc55b4d48, 32'hc3ed5f24, 32'hc44acd4a},
  {32'h444fc7e8, 32'h431819b6, 32'h43f75486},
  {32'hc42324b7, 32'hc42482a8, 32'h44845004},
  {32'h44801896, 32'h43c8e1e1, 32'h4276eeeb},
  {32'h44f22568, 32'h41125a9a, 32'h41ccddc2},
  {32'h43b32028, 32'h4535ac9f, 32'h43020b45},
  {32'hc47fd1e2, 32'hc4470415, 32'hc490a736},
  {32'h42f1f063, 32'h44957cf5, 32'hc34c6188},
  {32'hc3d00cd6, 32'hc36d40b8, 32'hc5083b15},
  {32'h4359d01c, 32'h443925f4, 32'h4362d392},
  {32'h44cbbd5f, 32'hc2c92258, 32'h436aaa86},
  {32'h44fc132c, 32'hc3be4872, 32'h44a6465c},
  {32'hc5694268, 32'hc3b5962a, 32'hc3665805},
  {32'h453973d4, 32'h43c161df, 32'hc3e29fc1},
  {32'hc3065ab0, 32'hc4b64484, 32'hc3e92bfe},
  {32'h43b21740, 32'h4380082c, 32'h4462fcb1},
  {32'hc2a2991c, 32'hc482e8f7, 32'hc400cf59},
  {32'h4487e20d, 32'h44b946fe, 32'h440c52b4},
  {32'hc50cfc30, 32'hc1def551, 32'hc447de83},
  {32'h453b15bc, 32'hc2b4c6a0, 32'hc4413e3d},
  {32'hc4c34ae7, 32'h432d2c4f, 32'hc38715c0},
  {32'hc4191039, 32'hc4ec9d31, 32'hc3dbb0c9},
  {32'h4466f78f, 32'h44b56097, 32'h43d34a66},
  {32'hc51339b3, 32'h42aac871, 32'h430bdf7c},
  {32'hc32a2158, 32'hc274d7be, 32'h435b1975},
  {32'hc51c3035, 32'hc441a7dc, 32'h43afab64},
  {32'hc4ad755e, 32'hc3818e1e, 32'h431e157f},
  {32'hc559fa2e, 32'hc3059539, 32'h43542af5},
  {32'h454ee4ad, 32'h43e75627, 32'h44130fc6},
  {32'hc5230da2, 32'hc40d2db5, 32'h43b4cf6d},
  {32'h44458a2e, 32'h446aabf7, 32'hc38bcc3e},
  {32'hc4d675e3, 32'hc3975b57, 32'h44246a77},
  {32'h44488c4c, 32'hc3183f5a, 32'hc47917f7},
  {32'hc4e4d6e3, 32'hc3c1171d, 32'h4369def0},
  {32'h43c43530, 32'hc34c7e2e, 32'hc339b456},
  {32'hc493feaa, 32'hc3bdf3e8, 32'h43f24a77},
  {32'h4503c439, 32'hc30b752c, 32'hc20d6fa3},
  {32'hc525fc64, 32'hc23132f1, 32'h434ef7b4},
  {32'hc4100691, 32'h43c99f4c, 32'hc4204d61},
  {32'hc4975e18, 32'hc449aeb2, 32'h442d36d4},
  {32'h449e3df8, 32'h44c2454c, 32'hc3a80054},
  {32'hc46e0a0d, 32'h43df97ed, 32'h41f99229},
  {32'hc2b14540, 32'hc3de5e9b, 32'hc538d8a8},
  {32'hc48ea681, 32'hc47650dd, 32'hc399f348},
  {32'hc39af49a, 32'hc2dc8c4e, 32'hc3b36007},
  {32'hc40fce98, 32'h44420ba5, 32'h444af143},
  {32'h43b54b70, 32'hc3a91abe, 32'hc48121d2},
  {32'h44472012, 32'hc50b70d5, 32'hc4032de8},
  {32'hc4abc999, 32'h448e9238, 32'h442d01db},
  {32'h42911d90, 32'hc4494827, 32'hc2dbfb01},
  {32'hc526019c, 32'h44023be8, 32'hc44044ab},
  {32'h43d687c7, 32'hc485d35f, 32'hc3f87d55},
  {32'h448041d8, 32'h42afc9df, 32'hc33bcbba},
  {32'h43fcfae0, 32'hc4cf1faa, 32'hc49fdf12},
  {32'hc4c39778, 32'h43c34c85, 32'h43a1898e},
  {32'hc462455f, 32'hc4261d52, 32'hc3d36799},
  {32'hc519bfdd, 32'h438dae28, 32'h441fbf64},
  {32'h4414436a, 32'hc486cba5, 32'h430b542a},
  {32'hc4786d12, 32'h4406e2fd, 32'hc427d37b},
  {32'h455b8e3a, 32'h43bd0d49, 32'h42c4b94e},
  {32'hc4b427f8, 32'h44b6096c, 32'hc1fef5c9},
  {32'h44e305d9, 32'hbf421000, 32'h439b8032},
  {32'hc48ac08e, 32'hc2ac57a4, 32'hc3973f87},
  {32'h44ed1086, 32'hc3f15c9a, 32'h42cfba34},
  {32'hc488a0dd, 32'hc35af7b0, 32'hc41da558},
  {32'h43693faa, 32'hc53825ae, 32'hc3081534},
  {32'hc4c091ea, 32'h44a0b383, 32'hc454482d},
  {32'h4561f91f, 32'h43f4cc0f, 32'h42ccf468},
  {32'hc480f1ef, 32'h44f90747, 32'hc2917d85},
  {32'h44126506, 32'hc30555aa, 32'h44e6c1fc},
  {32'h43cdc525, 32'h431dede9, 32'hc423fe5e},
  {32'h44e0cd47, 32'hc2945a36, 32'h44161445},
  {32'hc5224c95, 32'h4424d0e9, 32'hc3b8458c},
  {32'h440d4c31, 32'hc29b6eff, 32'h434998e1},
  {32'h43527045, 32'h429f41e2, 32'hc52f154a},
  {32'h4341bacf, 32'hc3c87c98, 32'h45391ebe},
  {32'h4377987b, 32'h443f1c56, 32'hc4beb941},
  {32'h44ecfe67, 32'h443ac66e, 32'hc36bd816},
  {32'h454963b8, 32'hc3a8521f, 32'h4400ef14},
  {32'hc4b4f923, 32'h446b4148, 32'h4371f703},
  {32'hc40cd8dd, 32'hc31c0b31, 32'h433b26b0},
  {32'hc30d6f6e, 32'h44df517e, 32'hc4786fad},
  {32'h43c59ce4, 32'hc410d910, 32'h44f3cddc},
  {32'hc4879a9f, 32'h4345811c, 32'h4436d706},
  {32'hc382228e, 32'h45149512, 32'hc4d390b4},
  {32'h44bede2c, 32'hc38f56df, 32'hbfe918da},
  {32'h44e89668, 32'h4381aed2, 32'h432f86b6},
  {32'hc42f371a, 32'h44c8b7f6, 32'h43f339c4},
  {32'h44ac6d3c, 32'h42530a8c, 32'h44270a77},
  {32'hc2b213eb, 32'h431a14b2, 32'hc4c4ad3e},
  {32'hc2a263bc, 32'hc4e64877, 32'h445cd9c4},
  {32'hc35093ac, 32'h45037e31, 32'h42e6be42},
  {32'h451a6c8c, 32'hc30354b2, 32'h43330d3a},
  {32'hc5838441, 32'h4344c681, 32'hc3b0f58c},
  {32'h450b0ba2, 32'h44279f9b, 32'h446b73ae},
  {32'hc4f66a40, 32'hc2e3c41d, 32'h4387f31b},
  {32'h442a76c9, 32'hc4b41b8a, 32'h442828da},
  {32'hc32a6300, 32'h432c5054, 32'hc41b9a4b},
  {32'h44490f41, 32'hc31dd521, 32'h423c6861},
  {32'hc3ea2b5f, 32'h44bd1dd6, 32'h432b3999},
  {32'h44a259fc, 32'hc4b23a35, 32'hc41b3840},
  {32'h43ffbd17, 32'h446247b9, 32'h43c4092d},
  {32'hc1d0a812, 32'hc4e6d038, 32'hc496b054},
  {32'hc4be4924, 32'h440312d9, 32'h44373295},
  {32'h43af13b6, 32'hc4bbe66a, 32'h447d194c},
  {32'h42cca190, 32'h4500d2f3, 32'h4370baf5},
  {32'hc4649eaa, 32'hc2f08050, 32'hc29ac3c6},
  {32'h427cfd00, 32'h44cc2488, 32'hc3b2fff6},
  {32'hc4ca1631, 32'hc40ab682, 32'h447afbef},
  {32'h43f8a700, 32'h44323425, 32'hc33ffb92},
  {32'hc46ec8fa, 32'hc436e720, 32'hc0209c2e},
  {32'hc403bef8, 32'h44d21d4d, 32'h44999de4},
  {32'h4395c4b3, 32'hc321911a, 32'hc4924103},
  {32'h45371293, 32'h4413144b, 32'h42d54075},
  {32'hc4202816, 32'hc4005cfd, 32'h44bcfa2b},
  {32'hc35d2349, 32'h44a08b68, 32'hc3c5dda2},
  {32'hc41bca47, 32'hc4f00a21, 32'hc37a1b0b},
  {32'h444f62d4, 32'h438a3d9a, 32'h43027847},
  {32'h4374feb8, 32'hc2e16e52, 32'h43810af3},
  {32'h453cf88e, 32'hc3c31e55, 32'h43534287},
  {32'hc445f275, 32'h431e7fb1, 32'h447a7d37},
  {32'h444033dc, 32'h43babd21, 32'hc123ae60},
  {32'hc4430e6c, 32'hc48b7e09, 32'hc314b6c5},
  {32'h439068f2, 32'h456dc81a, 32'h432de052},
  {32'hc335336c, 32'hc496fef4, 32'h43cba964},
  {32'h43a3041a, 32'h451014fd, 32'h427b3da4},
  {32'hc5411e00, 32'hc01f07e7, 32'hc284ad35},
  {32'hc478e28c, 32'h44855110, 32'hc3b75667},
  {32'hc3a9a40a, 32'h4485bed3, 32'hc2831de0},
  {32'hc477c92b, 32'hc461225e, 32'hc358e8cd},
  {32'h4483101c, 32'h43f04921, 32'hc2df180f},
  {32'h4208381c, 32'h41fb46e8, 32'hc2208175},
  {32'h42fae46c, 32'h43d3a101, 32'h44c16e18},
  {32'hc455ada2, 32'hc42c44ee, 32'hc40924a1},
  {32'hc41521f0, 32'h4389d360, 32'h43ae5870},
  {32'hc46a9e22, 32'hc20593ff, 32'hc4920670},
  {32'hc38b42a0, 32'h437154e0, 32'h44dddb09},
  {32'hc45af2f4, 32'hc35545ca, 32'hc117c422},
  {32'h43840522, 32'h450984f4, 32'h43459a09},
  {32'hc36919cd, 32'h449d9018, 32'hc4b9ac4e},
  {32'h4413c9f0, 32'h449fdd58, 32'h439ad5aa},
  {32'hc494607c, 32'hc3c7d94a, 32'hc3c9d32d},
  {32'hc28ae0c4, 32'h43a9939d, 32'h44bd7822},
  {32'h43dd52e4, 32'hc44a37b9, 32'hc385ad34},
  {32'hc3c2bfee, 32'h4509885a, 32'h44e8cfe2},
  {32'hc384ada0, 32'hc40104b9, 32'hc4268534},
  {32'h44254d84, 32'h4340844a, 32'h43ccfae3},
  {32'hc53277dd, 32'hc3ab10dd, 32'hc32061e6},
  {32'h43b43fbe, 32'h4561e5e8, 32'h43565aae},
  {32'h430ab89c, 32'hc4076b98, 32'hc3d4f594},
  {32'h41b9b940, 32'h450ab8bc, 32'hc3815f0a},
  {32'hc4414559, 32'hc4410ebc, 32'h42d79f51},
  {32'h44f54b40, 32'hc23f1988, 32'h44086adc},
  {32'hc43d1a6e, 32'hc2d5f507, 32'h41d28b12},
  {32'h44857a82, 32'hc411a3e5, 32'h43dc64cd},
  {32'h433142ab, 32'hc48bc727, 32'hc4039033},
  {32'hc4880771, 32'hc3753ca2, 32'hc35e1756},
  {32'h4464bb7d, 32'h437bd83d, 32'h436756b8},
  {32'h435b4730, 32'h452c0e79, 32'h41c13d1f},
  {32'h43cd9b3c, 32'hc437371a, 32'hc4ac8a95},
  {32'h44350bbc, 32'h43eb6789, 32'h410aecf1},
  {32'hc3f4d878, 32'hc4c9d929, 32'hc4f46d83},
  {32'hc380809d, 32'h446cb627, 32'h452b7fe8},
  {32'h44c00c5b, 32'hc3c2fcb1, 32'h431c426a},
  {32'hc4c1791c, 32'hc29f148f, 32'h447796f4},
  {32'hc323c330, 32'h422ea615, 32'hc493c504},
  {32'hc3b30932, 32'h441dc866, 32'h43face40},
  {32'hc36525c4, 32'hc474feb1, 32'hc3e58860},
  {32'hc53145be, 32'hc228b774, 32'h4226e1ce},
  {32'hc3086a10, 32'hc4b3f9d3, 32'hc3ad28e2},
  {32'hc50308f5, 32'hc214d669, 32'h4282fbdf},
  {32'h429f6b28, 32'hc496baea, 32'hc49b5002},
  {32'h441cce34, 32'h41d6feca, 32'hc3ce9dac},
  {32'hc3915dd0, 32'hc4950c1c, 32'hc3bae544},
  {32'hc51a9bba, 32'h437c5da2, 32'h438fdebc},
  {32'h4508d05a, 32'h43981a05, 32'hc0dd6787},
  {32'hc44a72c2, 32'h4452228c, 32'hc435213a},
  {32'h44b53228, 32'hc4cfcdb9, 32'h437c5d2c},
  {32'hc538dfd8, 32'hc2adc62f, 32'h429364ec},
  {32'h44a71364, 32'h43a8f79f, 32'hc3c124c0},
  {32'hc45dfd88, 32'hc3e078d2, 32'h43bb38fc},
  {32'h449e957b, 32'hc40166c0, 32'hc35cc13c},
  {32'h44e45a66, 32'hc36a1333, 32'h429e0828},
  {32'hc4e0d19e, 32'hc2a78acd, 32'hc4870229},
  {32'h4300e2c8, 32'hc35aa2e4, 32'h4390dc26},
  {32'hc508eee8, 32'hc34765d1, 32'h42b7ed78},
  {32'h44d56827, 32'h4414312a, 32'hc33825a5},
  {32'hc18ef145, 32'h455063e8, 32'h43a7f57a},
  {32'h45453979, 32'hc1e3c6a4, 32'hc2351f47},
  {32'hc53cab4c, 32'h43421052, 32'hc38747fc},
  {32'h442f89ae, 32'hc500ce37, 32'h43a7f232},
  {32'hc3473664, 32'hc38f89f3, 32'hc327d3c5},
  {32'h442e27bf, 32'h43d1b4ce, 32'h44f3bfdd},
  {32'hc3d33ce2, 32'hc4959990, 32'hc4ea0ea7},
  {32'h44010416, 32'hc328ba4c, 32'hc341cd66},
  {32'hc3427984, 32'h45025524, 32'h43d93593},
  {32'hc1e390f7, 32'hc34fbc60, 32'hc4a6027f},
  {32'h445d58b3, 32'h4391ad4c, 32'h449c963d},
  {32'hc38eb758, 32'hc492948d, 32'hc4140653},
  {32'hc4122cd2, 32'h4420f5e1, 32'h44e8ac5e},
  {32'hc4ef28f5, 32'hc409b661, 32'hc2096eb8},
  {32'hc506bbb6, 32'h444a9f74, 32'h4445bf1e},
  {32'h44b640d5, 32'hc479de71, 32'hc48c7efe},
  {32'hc444ae7c, 32'hc3e073dd, 32'h43e428e6},
  {32'h4470b34d, 32'hc48c201c, 32'hc42e7636},
  {32'h42d39250, 32'h428fda2d, 32'h44f94b9d},
  {32'hc3ddb38e, 32'hc4018c8c, 32'hc372c7cb},
  {32'hc402e001, 32'h4492e658, 32'h4507940c},
  {32'h451690cf, 32'hc3e526d5, 32'hc3f847b5},
  {32'h447172b4, 32'hc3a229ff, 32'hc48593a5},
  {32'hc5295736, 32'h425404d2, 32'h44442fc0},
  {32'h43086060, 32'h43ed3757, 32'h44008cb3},
  {32'hc4045664, 32'hc44d6a33, 32'h438e8ce8},
  {32'h44b5d100, 32'h448f354e, 32'hc2ad8f3d},
  {32'hc4f4228b, 32'h436e4089, 32'h41181e0a},
  {32'hc20e0560, 32'h45086050, 32'h422042de},
  {32'hc58c23b1, 32'hc3927bd7, 32'hc40d41ec},
  {32'hc461d1c8, 32'h44180e92, 32'h42d9231f},
  {32'hc51ce08c, 32'h4296a498, 32'hc3b8dc32},
  {32'h4534bd5b, 32'h431ebfb2, 32'h4383c143},
  {32'hc4d80d6d, 32'h4356b524, 32'h42fc68f4},
  {32'h4451da2d, 32'h422b49aa, 32'h44fd0a45},
  {32'hc45cb358, 32'hc4da0615, 32'hc4493a35},
  {32'hc23dd794, 32'h43908b5a, 32'h4457e426},
  {32'hc33daa4b, 32'hc521c61c, 32'h429bd01b},
  {32'h42907a6d, 32'h43b0da1c, 32'h456aafb0},
  {32'hc2c9760c, 32'hc40629a5, 32'hc4a2874f},
  {32'h4476228c, 32'hc3efd793, 32'h43e35353},
  {32'hc53750bb, 32'hc317d94a, 32'hc39ce7e9},
  {32'h446d8992, 32'h43c40c03, 32'hc3252ece},
  {32'hc4f64424, 32'hc2d97b3f, 32'hc462aba2},
  {32'hc396a31f, 32'hc29fb772, 32'h453624c7},
  {32'h441d23b2, 32'hc4b892dd, 32'hc37cf34b},
  {32'h4415eacd, 32'h4424708b, 32'h44882bc7},
  {32'hc5344b62, 32'hc329d3e4, 32'hc307b61f},
  {32'hc4680c5a, 32'h43e06977, 32'hc3612d4c},
  {32'hc222d62e, 32'h44c41ecc, 32'h43d790df},
  {32'h435218fa, 32'hc50d41e0, 32'h4261fe27},
  {32'h428774e0, 32'h45026419, 32'h438c505a},
  {32'h43bfaf7e, 32'h422d8cae, 32'h418c3610},
  {32'h4515df28, 32'h43aa6157, 32'hc411b3a4},
  {32'hc506afc2, 32'hc49c1905, 32'h425cf372},
  {32'h44388b57, 32'hc21053f3, 32'h433012a4},
  {32'hc58ce588, 32'h43876dd3, 32'hc3da0226},
  {32'hc395fc80, 32'h4411bead, 32'h43d8f609},
  {32'h43f4bcf5, 32'hc49af224, 32'h434fa7e0},
  {32'h43028e42, 32'h45214807, 32'h42092878},
  {32'hc4f2a9f0, 32'hc401b7ee, 32'h434d8691},
  {32'hc3cd7ca4, 32'h43ca37ff, 32'h428f6f04},
  {32'hc505501d, 32'h438998a2, 32'hc2d4e69d},
  {32'h452e8084, 32'h43d383f0, 32'hc2926f7a},
  {32'hc4a9d8dc, 32'h43f29c4b, 32'h426a4884},
  {32'h443a979b, 32'hc41fd54c, 32'hc4610ec9},
  {32'hc3a0d788, 32'h44210646, 32'h4547ca74},
  {32'hc3879858, 32'h443dc41e, 32'h433e2f0c},
  {32'hc367c19c, 32'hc54b6ed0, 32'h42c0e1b4},
  {32'h45421d12, 32'h43c3e130, 32'h430b0910},
  {32'hc2ef7db9, 32'hc3823287, 32'h4493bf08},
  {32'h419b5d40, 32'h450f3029, 32'hc3f53f7c},
  {32'h431a3f6e, 32'hc50c9ac8, 32'h43ca5624},
  {32'h43525832, 32'h43db7c12, 32'hc48b7933},
  {32'hc43adbc0, 32'h42d27d37, 32'h441338f2},
  {32'h457f6f71, 32'hc42161bd, 32'hc35d0b5e},
  {32'h4520c54c, 32'hc3a9769d, 32'hc44e602e},
  {32'hc4fb6df6, 32'h43bb848f, 32'h427926e4},
  {32'h44819537, 32'h42a37ffa, 32'hc41b8da4},
  {32'hc471bd5c, 32'h44e4a906, 32'hc3c2fc85},
  {32'h4528422a, 32'hc308e48d, 32'hc3920e5f},
  {32'hc38c2fa4, 32'hc226ce60, 32'hc3adb488},
  {32'h455383f2, 32'hc32f506e, 32'hc40e1702},
  {32'hc45df758, 32'h426be8ac, 32'hbfc65718},
  {32'h453bc4c6, 32'hc2b246dc, 32'h434cf599},
  {32'hc52dcfe0, 32'h439d813a, 32'h443c395c},
  {32'hc393a8dc, 32'hc4ee1051, 32'hc39a7401},
  {32'hc3a3f3f0, 32'h42ae82f2, 32'hc38333b6},
  {32'h4359eab2, 32'hc3cdfa2b, 32'h446f9197},
  {32'hc5148cf5, 32'hc3f98ed3, 32'hc4177ed8},
  {32'h4380b190, 32'hc3ca701d, 32'h4358c559},
  {32'hc3b32b6a, 32'hc39a4919, 32'hc51345d4},
  {32'h45181ab1, 32'h43821ac0, 32'hc397cc2c},
  {32'hc50c5e76, 32'hc113a072, 32'h41e0b15c},
  {32'h44cec0a2, 32'hc48ea551, 32'h42b35068},
  {32'hc4466036, 32'h453702b9, 32'hc3a88c33},
  {32'h43aba216, 32'h41ac125e, 32'h4433a5b8},
  {32'hc4b8533a, 32'h44a9bf21, 32'hc3a54f4a},
  {32'h449b5958, 32'hc4a728c6, 32'h428cfd9b},
  {32'h42b6ed42, 32'h449120e8, 32'hc406bc21},
  {32'h447c4aac, 32'h448ef213, 32'h432f3744},
  {32'hc569adb8, 32'hc2981996, 32'hc2dc4eec},
  {32'h4429af18, 32'h43b77758, 32'h448042ce},
  {32'h4412acef, 32'h432adf5f, 32'hc4b54a1a},
  {32'h419c91c0, 32'hc3313732, 32'h456b63c6},
  {32'h44b1c321, 32'hc399f732, 32'hc3bee3d6},
  {32'hc505eab4, 32'h431da0c0, 32'h42d01441},
  {32'h44f19164, 32'hc4998ad9, 32'hc335c1f8},
  {32'hc22d41e0, 32'hc382d4f2, 32'hc48c5ca8},
  {32'h43cde394, 32'h43b85503, 32'h44bd01fb},
  {32'hc55a1548, 32'h436bc2c5, 32'h41b95cab},
  {32'h44b23275, 32'hc4041978, 32'h43843269},
  {32'h44ad4680, 32'hc1d68671, 32'h43aff18e},
  {32'hc4b218d8, 32'h44b7d40e, 32'hc4aeeef2},
  {32'h4511289c, 32'hc30ef0a6, 32'hc4975ca9},
  {32'h44e72a75, 32'hc33da54c, 32'hc3804fb7},
  {32'h43b8a1c8, 32'h454f7be2, 32'h43cce8ae},
  {32'h45193779, 32'h4352faaf, 32'h42b2474b},
  {32'h4484f3f5, 32'hc306768c, 32'hc49f5152},
  {32'hc39bf020, 32'hc3dc275c, 32'h4486aa24},
  {32'h415cc6a8, 32'hc2d67be4, 32'hc4e850b3},
  {32'h44b4cdc8, 32'hc2b3297e, 32'h447cc8ce},
  {32'hc5842b41, 32'hc3a0f9d0, 32'hc344bd9f},
  {32'h44900d8c, 32'hc4210076, 32'h4346fd85},
  {32'h43b566bc, 32'hc344fb61, 32'h43668c31},
  {32'h43cf59f2, 32'hc5101be4, 32'hc464b419},
  {32'hc4d2ce83, 32'h43a020ac, 32'h42c64880},
  {32'h44bc1744, 32'hc4146e34, 32'h42aff51d},
  {32'h42ba1de4, 32'h456dd2e8, 32'h438bac7d},
  {32'h442bf10a, 32'hc4d8f476, 32'hc412fd44},
  {32'h43efd005, 32'h44ac70a3, 32'h44862974},
  {32'h43e0043a, 32'h44cff741, 32'hc489a82d},
  {32'hc3710350, 32'h4445095d, 32'h4549c68b},
  {32'hc32742a8, 32'hc5225908, 32'hc2c25513},
  {32'h42318112, 32'h4381aa2a, 32'hc4b982f9},
  {32'h437cfd9e, 32'hc48ad63c, 32'h43048efc},
  {32'h42b7e190, 32'h44fd1983, 32'hc498bf29},
  {32'h42c94320, 32'hc458da09, 32'h439ea61c},
  {32'h4475a548, 32'hc39b0545, 32'hc45e1104},
  {32'hc2a4bc0c, 32'h44315592, 32'h43b7eb3f},
  {32'hc48c8eea, 32'h440b779e, 32'h442bcb28},
  {32'h451b7af7, 32'h4300d85c, 32'hc43124f0},
  {32'hc313da1c, 32'hc36474c6, 32'hc4d74f5a},
  {32'hc3a3416e, 32'hc386d3cf, 32'h4442a122},
  {32'hc47093d6, 32'h441ed1ad, 32'hc3bd948b},
  {32'hc485dde0, 32'hc3d45cb5, 32'h44765688},
  {32'hc3577294, 32'hc2bb06db, 32'hc562a0c4},
  {32'h45023aaa, 32'hc327cf28, 32'h43853c50},
  {32'h42171700, 32'hc3a4a69f, 32'hc45f46f4},
  {32'hc5968a3a, 32'hc36b7de6, 32'hc4140032},
  {32'h45254bb8, 32'hbf7f2bc8, 32'hc374cfa7},
  {32'hc55dca84, 32'hc30b14c8, 32'h42ed23c2},
  {32'h41c40878, 32'h45599086, 32'hc26adb42},
  {32'hc5343de2, 32'h4304e415, 32'h43a0434a},
  {32'h44adcf0b, 32'h44f9c4a4, 32'hc3b73acb},
  {32'hc53ad9b4, 32'hc40faa02, 32'hc35d061a},
  {32'h44497119, 32'h42cd85a8, 32'hc24c4bf7},
  {32'hc4214d60, 32'h44c03d69, 32'hbf8e23d0},
  {32'hc415f1d8, 32'hc50e66d0, 32'hc3f8fdbb},
  {32'hc3d72b16, 32'h44096f02, 32'h441fb07d},
  {32'hc1f642c8, 32'h427feba0, 32'hc4b71d08},
  {32'h440e004d, 32'h45089eb3, 32'h448141ef},
  {32'h42c82dee, 32'hc4ed5e9c, 32'hc2d03edc},
  {32'h41627f30, 32'hc38e6fd7, 32'h44c8b44f},
  {32'hc50134d0, 32'h43212804, 32'hc3edf616},
  {32'h42fb7ba0, 32'h44d3dac2, 32'h44d7e8ff},
  {32'h43f3c2c4, 32'h438dae34, 32'hc43513aa},
  {32'h4445440d, 32'h44cb23a0, 32'hc38ff90b},
  {32'h43f8c233, 32'h43bbcb43, 32'hc507843f},
  {32'hc3777801, 32'hc3734645, 32'h44ca8430},
  {32'hc4824c28, 32'hc4a51e94, 32'hc2351672},
  {32'h44ab7500, 32'h4400632e, 32'h4390d3e7},
  {32'hc3cb1018, 32'hc3d19c6f, 32'h433ddb34},
  {32'h43ff89e4, 32'h446ccdab, 32'h442f02c7},
  {32'hc4c1e370, 32'h430db2a7, 32'hc48fdd4d},
  {32'h452f75e2, 32'h42f0931e, 32'h43012506},
  {32'hc3d08760, 32'hc573fc8f, 32'hc3c6d756},
  {32'h45018c08, 32'h4441946f, 32'h436fdff4},
  {32'hc5345ea9, 32'h43fe85ae, 32'h415e933e},
  {32'h4361e1ae, 32'h44967630, 32'h44079221},
  {32'hc42b572b, 32'hc4c9f9b4, 32'hc3e5b6a3},
  {32'hc47f64b9, 32'h439dd1cf, 32'h433d1866},
  {32'hc40cbab0, 32'h436fcb42, 32'hc40e911e},
  {32'h44f790cd, 32'hc4055679, 32'h42716c76},
  {32'hc36315ae, 32'h44fd3672, 32'hc4e31e9b},
  {32'h42c9a8be, 32'hc4df72f1, 32'h44ab3a45},
  {32'hc4021f63, 32'h43bbad88, 32'hc4113c86},
  {32'hc4808920, 32'h43f27f82, 32'h449df6cf},
  {32'hc28f6268, 32'hc4e303b9, 32'hc481c33d},
  {32'h440a5309, 32'h42b5228b, 32'h448cf4df},
  {32'hc0a45000, 32'hc4215ab3, 32'hc4decbd7},
  {32'hc461f564, 32'h4426535a, 32'h44ae9b4e},
  {32'hc414b9f6, 32'hc44e510e, 32'hc39bd6bf},
  {32'hc4923ddd, 32'hc2bf0b96, 32'h4433b570},
  {32'hc34874f0, 32'h44b948a8, 32'hc50d58e8},
  {32'hc28386ac, 32'h447148c7, 32'h430dd292},
  {32'h4495048a, 32'hc2f3c4d1, 32'hc43a1494},
  {32'hc3a4b458, 32'h4442b4a3, 32'h438b9846},
  {32'hc39cb6e8, 32'h42ef6b42, 32'hc4ce1ae5},
  {32'h4452b5f7, 32'h44a8d959, 32'h450dee29},
  {32'h43b6a4ec, 32'hc40c97ba, 32'hc4fb5141},
  {32'h416d1048, 32'h436296f7, 32'h43833505},
  {32'h42dcea74, 32'hc57ca208, 32'h43913315},
  {32'hc4ede0c6, 32'h44c72bb9, 32'hc357615d},
  {32'h4495dbe6, 32'hc424c4a2, 32'h431596ce},
  {32'hc40c21a9, 32'h452316ef, 32'h43332021},
  {32'h44ac8a18, 32'hc2b53849, 32'hc3c745d4},
  {32'hc3452358, 32'hc3818ee1, 32'h42bee241},
  {32'h44eb5992, 32'h4410ad54, 32'h43e4f8db},
  {32'hc54b936d, 32'hc3056a16, 32'h43962ab4},
  {32'h454f5fd8, 32'hc35a40ae, 32'hc408c122},
  {32'h45010028, 32'h42422936, 32'h43f730dc},
  {32'hc46b419c, 32'hc3210937, 32'hc5021144},
  {32'h42d21814, 32'h43f0a4cc, 32'h45541779},
  {32'h44fa3694, 32'hc38d7064, 32'h42ced10c},
  {32'h4438608c, 32'hc4e2960d, 32'h436a570d},
  {32'h432303a8, 32'h45084ef4, 32'hc3a03dcb},
  {32'h453def17, 32'h43b7fefa, 32'h434ab6b9},
  {32'hc5625512, 32'h43e35f71, 32'h43511d47},
  {32'hc2c6fac0, 32'hc48d92bb, 32'hc3ec7e35},
  {32'h4200dc88, 32'hc39af0d5, 32'hc49db22e},
  {32'h451f2a3b, 32'hc34cb356, 32'hc2583787},
  {32'h43239488, 32'h42925740, 32'hc3e64c62},
  {32'h43e612f4, 32'hc3952daa, 32'hc2a3ce84},
  {32'hc37e01d4, 32'h44a724f3, 32'h442820fd},
  {32'h44d2598f, 32'hc401aad5, 32'hc3ab379f},
  {32'h44e7d699, 32'h4268fa03, 32'h42d2a81b},
  {32'h453fba91, 32'h42148714, 32'hc324b2b5},
  {32'hc4bc4eaa, 32'h435715a1, 32'h432bdb56},
  {32'h43cacab7, 32'hc340f621, 32'hc3672a65},
  {32'hc56291ef, 32'h430c382e, 32'h43ef825b},
  {32'h4235bb40, 32'h442b693e, 32'hc41862dd},
  {32'h43818753, 32'hc2bab8e5, 32'h43540266},
  {32'h44292b98, 32'hc4968ed7, 32'hc495e27d},
  {32'hc4816370, 32'h43a80012, 32'h43b5bc68},
  {32'hc487a204, 32'hc3c0dc84, 32'hc3c8db4e},
  {32'hc3fb1557, 32'h432932fb, 32'h437b1f06},
  {32'h429ea7e8, 32'hc43a4899, 32'hc52b1e44},
  {32'hc2ff233a, 32'h43347058, 32'hc529d3da},
  {32'hc4a36b30, 32'h42fb7780, 32'h450c6da2},
  {32'h441780a6, 32'h426a9e45, 32'h4354176c},
  {32'hc45a6eb8, 32'hc4b17001, 32'hc384fada},
  {32'h450c6723, 32'hc316d4ab, 32'hc406d64a},
  {32'h440aee81, 32'hc2a7726e, 32'hc3e2af94},
  {32'h44a7ac81, 32'h4491ceee, 32'hbfb9dda0},
  {32'hc5504c06, 32'hc423cc9e, 32'hc43ca18f},
  {32'hc2cb6e10, 32'h44b54d32, 32'h43c96d7a},
  {32'h4375c8d0, 32'hc44c3381, 32'hc3a8ea83},
  {32'h44058fb4, 32'h4474aec7, 32'h44559f9e},
  {32'hc3b61256, 32'hc39a01aa, 32'h43c679f1},
  {32'h43bd4c79, 32'h450f1e44, 32'h44073eb0},
  {32'hc49275da, 32'hc43f9d5e, 32'hc4a241cb},
  {32'hc38d4d48, 32'h44ccc118, 32'hc0b2fc96},
  {32'hc277ea96, 32'hc5311efc, 32'h43d10285},
  {32'h431b999a, 32'h44d88f7f, 32'h4454f5a4},
  {32'h44cea5ef, 32'hc426c749, 32'hc3e5555a},
  {32'hc26ba590, 32'hc466e0da, 32'h444c5a3d},
  {32'hc53c1b93, 32'hc38c5d5a, 32'hc3831763},
  {32'h451210cd, 32'hc3c8dd42, 32'hc3c3788b},
  {32'hc3993f36, 32'hc3969613, 32'hc506efaf},
  {32'h42edf79c, 32'h44e588bd, 32'hc2422897},
  {32'h4339261a, 32'hc4e67c5a, 32'hc387f6ff},
  {32'hc262d8af, 32'h4412acf8, 32'h455c0790},
  {32'hc3d7b0c2, 32'hc4efebc8, 32'hc201fd36},
  {32'h44033dbc, 32'h44a355b4, 32'h42873151},
  {32'h444136c0, 32'hc31bcdec, 32'hc40a82a1},
  {32'hc4911176, 32'hc467b634, 32'h438e1795},
  {32'h43845d23, 32'h451409cc, 32'hbf0b4184},
  {32'hc4b49505, 32'h40a31727, 32'h420cf350},
  {32'h44dcae2f, 32'h42bd8f0a, 32'hc24acb67},
  {32'h438cae7c, 32'hc52f47c0, 32'hc392394d},
  {32'h452ab479, 32'hc3b8bfed, 32'hc424b98d},
  {32'hc4600514, 32'hc42e6ab2, 32'hc3d79208},
  {32'h4424f33a, 32'h44816eac, 32'h44849b1a},
  {32'hc3b5af98, 32'hc2fe8a81, 32'hc29856ea},
  {32'h445a73c4, 32'h43ee62b6, 32'hc392d2f1},
  {32'hc4c2012b, 32'hc3b20960, 32'hc35d9684},
  {32'hc38a0164, 32'h4415ca6a, 32'hc0c8c2ac},
  {32'hc1563b98, 32'hc33558da, 32'h44d244ad},
  {32'h44f6b247, 32'h443c8694, 32'hc325a42f},
  {32'hc4a7bcf3, 32'h43dc0a75, 32'hc39dd4b4},
  {32'h44dd456c, 32'h4352e3f4, 32'h42b233fc},
  {32'hc31db390, 32'h41a35578, 32'h41b18c36},
  {32'h42d88e80, 32'h44185a68, 32'hc422f973},
  {32'hc3b485b5, 32'hc4ee20d2, 32'h441b2973},
  {32'h43fdedf8, 32'h4562223e, 32'h438c1952},
  {32'hc4e74157, 32'h41fd8cfd, 32'hc1a7b98c},
  {32'h44ae9c62, 32'h42d7e6ba, 32'hc5030523},
  {32'h439c9576, 32'hc42ae942, 32'h44f724fb},
  {32'h44669816, 32'h430cb781, 32'h428899ef},
  {32'hc4c292d6, 32'h44001021, 32'h446087a9},
  {32'h44a9123a, 32'hc38bc888, 32'hc49b66aa},
  {32'h44a6ecfe, 32'hc502be74, 32'hc38ec4f6},
  {32'hc460c642, 32'h44b2b6ef, 32'h43f6eeb5},
  {32'hc3be60e4, 32'hc4cf552f, 32'hc343c106},
  {32'hc49b4e29, 32'h407668fa, 32'h4432c3b7},
  {32'h43b463ac, 32'hc445d94a, 32'hc35c74a9},
  {32'h43876ef8, 32'h443917ce, 32'h43197245},
  {32'h44cff348, 32'h440853f2, 32'h42e02982},
  {32'hc47905d1, 32'h438dc3d5, 32'h43d765a4},
  {32'hc4ec148f, 32'hc38a83bb, 32'h431141c0},
  {32'hc3b7971e, 32'h44926235, 32'h41896ebc},
  {32'h4221ec74, 32'h44956b06, 32'hc4f1178b},
  {32'h43ef736f, 32'h438870bd, 32'hc427976b},
  {32'hc3b932df, 32'hc41d1f9e, 32'hc3b47635},
  {32'hc31c5912, 32'hc3851161, 32'hc5024706},
  {32'h439c15a6, 32'hc40fb540, 32'h43f77c9a},
  {32'hc1337558, 32'hc3676129, 32'hc4e24320},
  {32'h435b7d00, 32'h43d35749, 32'h44f5c06e},
  {32'hc4601f10, 32'hc31be07e, 32'hc3cf18d9},
  {32'h446b293f, 32'hc514640b, 32'hc3ae5605},
  {32'hc2dfb9c0, 32'h4416685e, 32'hc4f21f17},
  {32'hc4378910, 32'hc38c706e, 32'h441bd24b},
  {32'hc2fe7020, 32'h44b17d04, 32'hc4133e07},
  {32'h44879340, 32'h43652a78, 32'h441a128e},
  {32'hc32fa1a0, 32'h447121ab, 32'hc394b722},
  {32'h40809200, 32'h441b143d, 32'h44ecff9d},
  {32'hc526eec9, 32'h43a0760e, 32'hc28d742b},
  {32'h44cb8a2c, 32'hc42fc164, 32'hc2f7a0f2},
  {32'hc37ac6b8, 32'h44813385, 32'hc4e2a0d3},
  {32'hc31a7594, 32'h445c35a2, 32'h44b13c64},
  {32'hc487ad07, 32'h4466bfd4, 32'hc42696f5},
  {32'h44740a0d, 32'h439c88a0, 32'hc469f551},
  {32'h44b14c12, 32'hc48f24f3, 32'hc2856fbc},
  {32'hc3037a28, 32'h4522846e, 32'h42f3824c},
  {32'h43ac4a0d, 32'h439476e7, 32'h4492e7c4},
  {32'hc5225174, 32'h43964378, 32'hc1020c89},
  {32'h451ca38f, 32'hc3e19c70, 32'h4367ba06},
  {32'h44186f60, 32'hc42439c5, 32'h44d9aea6},
  {32'hc42c8ca0, 32'h4498caa8, 32'hc494dbbd},
  {32'hc4077e72, 32'hc485e892, 32'h441cd553},
  {32'h440a5886, 32'hc452d4c8, 32'h43083100},
  {32'hc47fe852, 32'h445cf406, 32'h42c5b115},
  {32'hc3792e2d, 32'hc5372caf, 32'hc397eae9},
  {32'hc4893e34, 32'h44090b87, 32'h43fb1183},
  {32'h450d00b0, 32'hc3b9ed0a, 32'hc35f22a0},
  {32'hc39eb280, 32'h4516eb51, 32'hc1a9681d},
  {32'h44b06650, 32'hc3d8a7a6, 32'hc2408e4a},
  {32'hc543e73b, 32'hc30ebda8, 32'hc3f2d6f2},
  {32'h44f1a636, 32'hc2cc6caf, 32'h43fb4cba},
  {32'h447eeb8f, 32'h44a8bb3a, 32'h427058ee},
  {32'h452dbad7, 32'h43073cdc, 32'h42a6e03c},
  {32'hc554b19d, 32'h43f0f33d, 32'hc386a4e2},
  {32'h445b474e, 32'h443c8832, 32'h43b70c52},
  {32'hc49d399f, 32'h450d752a, 32'h43164c62},
  {32'h44b0d4b2, 32'hc3b4821b, 32'h43869d97},
  {32'h447bf19b, 32'h436c2c9b, 32'h434c6be3},
  {32'hc2e469c0, 32'hc4a716bc, 32'hc491d009},
  {32'h41972da0, 32'hc3e2a0e1, 32'h44a40bf5},
  {32'hc49306cf, 32'h42cb9124, 32'h442b7720},
  {32'h42985cf6, 32'h45418347, 32'h42953467},
  {32'h43a0bbf0, 32'hc342e57f, 32'h44cf2437},
  {32'hc3275f7e, 32'h441860ee, 32'hc4a692ab},
  {32'hc55154e1, 32'hc4035000, 32'h43a26c18},
  {32'h44e470f7, 32'hc39c3ad7, 32'hc28cc315},
  {32'h42bc843c, 32'h42a3ca16, 32'hc463807a},
  {32'hc4020906, 32'hc394975f, 32'h43efbd8d},
  {32'hbf83f800, 32'hc39f3499, 32'hc4d5427e},
  {32'h42b71909, 32'h43210c45, 32'hc5166f3b},
  {32'hc3a4ae2e, 32'hc421c8c7, 32'h44213dc3},
  {32'h44a76861, 32'h437ddcdf, 32'hc420e9c9},
  {32'hc5082d23, 32'h42116d96, 32'h443a959e},
  {32'h43e96078, 32'h440cb8a5, 32'hc49a9fc4},
  {32'h440a39d1, 32'hc403bfca, 32'h4398715b},
  {32'hc22b4248, 32'h4345dcc7, 32'h44277cb9},
  {32'hc3a92b7b, 32'h4468836a, 32'h43a24073},
  {32'h4504923b, 32'h4361ca42, 32'hc3468598},
  {32'h42b0100a, 32'hc5444397, 32'h43863535},
  {32'h44699f6e, 32'h44ee3c1e, 32'h438c6e3f},
  {32'h4508594e, 32'h4265d78e, 32'hc2dbf310},
  {32'h44da1d80, 32'h44a1c5d2, 32'hc35ee84c},
  {32'hc4a73172, 32'hc4d88714, 32'hc38eeb24},
  {32'h4523ce6e, 32'hc432b25c, 32'hc3c0be52},
  {32'h447899aa, 32'hc452738e, 32'h439ffe9c},
  {32'hc50a5b29, 32'h427af078, 32'hc2ca0b00},
  {32'h44f8d70a, 32'h429efe1f, 32'h4403aa91},
  {32'h43af55a2, 32'hc3bbd9da, 32'hc4067b85},
  {32'h43e8259a, 32'h4424af51, 32'h4423407c},
  {32'hc39059a1, 32'hc49035fc, 32'hc44f9d02},
  {32'h42e726c0, 32'h442a9824, 32'h436a8018},
  {32'hc3956d54, 32'hc461798c, 32'hc4f44bcf},
  {32'h443e2832, 32'h43bf7d94, 32'h453b5da9},
  {32'h42b242fc, 32'hc31f4fa5, 32'hc3eefb86},
  {32'h436830fc, 32'h44886376, 32'h444d989d},
  {32'h4316aee8, 32'h44e6f6d8, 32'hc52073f8},
  {32'h45414676, 32'hc3a324f4, 32'h437eb009},
  {32'hc27967e0, 32'hc4cbde7e, 32'hc4542300},
  {32'h446b417e, 32'hc19deed7, 32'h43e98251},
  {32'hc4e187d5, 32'hc2c9c250, 32'h43b65438},
  {32'h446fdfb5, 32'h43c5c450, 32'h44bcda6c},
  {32'hc3a03efc, 32'hc4b7ef78, 32'hc49eade0},
  {32'h4514b7f7, 32'hc393514b, 32'hc374e666},
  {32'hc4460cac, 32'hc33f0a5e, 32'h4205e0ba},
  {32'h44ade419, 32'h44a6ee9e, 32'h4434f695},
  {32'hc53608d6, 32'hc32e54b2, 32'hc33e42d0},
  {32'h453b8abd, 32'h42fc5043, 32'h43a459c2},
  {32'hc488746e, 32'hc4b37709, 32'hc2b80627},
  {32'h43397ff4, 32'h43c5bd05, 32'h43c66e30},
  {32'hc48ffd37, 32'h4453a583, 32'hc487b213},
  {32'h45661600, 32'h42b6ed24, 32'hc377873d},
  {32'h4289c910, 32'hc42ea8d6, 32'hc3e39e48},
  {32'hc4655374, 32'h416949aa, 32'h439e91d2},
  {32'h43b576e4, 32'hc4a55c9d, 32'hc3f63347},
  {32'hc48088a5, 32'h440a7b63, 32'h4488c7cf},
  {32'h44c4dc4e, 32'hc3a6e515, 32'h42f1be09},
  {32'hc39392ea, 32'h43e5b000, 32'h43c5ba47},
  {32'h44dc9509, 32'hc3895ef1, 32'hc48849a5},
  {32'hc3eddf68, 32'h43f179d2, 32'h452fb4d4},
  {32'hc46492d7, 32'hc395e16f, 32'hc4c1e603},
  {32'hc4fd0795, 32'hc3e854f5, 32'h44628cca},
  {32'hc2dcbdde, 32'h42523dd5, 32'hc4d757ad},
  {32'h431a769b, 32'hc4cf8378, 32'h4457160a},
  {32'h43915044, 32'hc4054f4d, 32'hc461eac2},
  {32'hc2cfac08, 32'h4014dcc0, 32'h44709de4},
  {32'h43d45b85, 32'hc2f942ba, 32'hc45f22f1},
  {32'hc46787d6, 32'h44a0a55b, 32'h448ebb57},
  {32'h43663c7e, 32'hc3d333b1, 32'hc55a02e9},
  {32'hc4e7dd26, 32'h43f8b338, 32'hc34b65dc},
  {32'h4527944c, 32'hc42b2c86, 32'h43db68b8},
  {32'h427ea2e6, 32'h45656ecd, 32'h439b4699},
  {32'h438fdd24, 32'hc4d1272a, 32'hc25ba8c5},
  {32'hc546057e, 32'h4343f326, 32'hc2d61cbd},
  {32'h451e2a30, 32'hc41cad32, 32'h43857010},
  {32'h446e2625, 32'h43bbcf0b, 32'h4324590f},
  {32'h44ac0e74, 32'hc3677101, 32'hc3acb1fe},
  {32'hc4428742, 32'hc3c4094e, 32'hc3b7f3c7},
  {32'hc4fc254a, 32'hc3574e98, 32'hc41033af},
  {32'h44934e69, 32'h43214f73, 32'h44bf9d5e},
  {32'h41da5140, 32'hc24870f9, 32'hc559805d},
  {32'h44c95583, 32'hc3a7d2b8, 32'h4487f5ed},
  {32'h436904ec, 32'h440bcffc, 32'hc40b3ca6},
  {32'h450c77e2, 32'hc404254d, 32'hc1e0c15a},
  {32'hc441da4e, 32'h44b96e80, 32'h42529548},
  {32'hc47050a0, 32'hc40c7663, 32'h4382ec85},
  {32'hc50bc452, 32'h440797a9, 32'h42fc97af},
  {32'h44e015fc, 32'hc431158d, 32'hc3a1d662},
  {32'hc494eb67, 32'h4300fea5, 32'hc2c10153},
  {32'h450463ff, 32'h404525c0, 32'h439a1f6c},
  {32'hc5167f1d, 32'h43fa021d, 32'h440bf70a},
  {32'h43630749, 32'hc3ac0ae9, 32'hc4c414e6},
  {32'h42cbe409, 32'h44ebb672, 32'hc1175a62},
  {32'h442c3974, 32'hc35d72d3, 32'hc308f209},
  {32'h42327570, 32'h437d1e3f, 32'h44756819},
  {32'hc3bbf492, 32'hc4dfa070, 32'hc3e061c6},
  {32'hc3e7eee6, 32'h44b42592, 32'hc3025a6b},
  {32'hc38ae23f, 32'hc38dd541, 32'hc184f277},
  {32'hc4d6e411, 32'hc411d9b1, 32'hc27ff835},
  {32'hc38ca988, 32'hc49812e4, 32'hc467b0a2},
  {32'h44adf653, 32'h441442c0, 32'hc1a28d21},
  {32'h44f06d68, 32'hc405af68, 32'hc3db43ff},
  {32'hc4b40711, 32'h4439aa9e, 32'h44664b93},
  {32'h43fc2a0d, 32'h4330de61, 32'hc361723e},
  {32'h4350fb37, 32'h44d16803, 32'h440852d6},
  {32'h443d0390, 32'hc45faf01, 32'hc4ea7444},
  {32'h44de93ca, 32'h4318084e, 32'hc489e3cb},
  {32'hc508e9b3, 32'hc37eb286, 32'h43f6c9c7},
  {32'h44b79cb7, 32'h43b5ad5c, 32'h431c662e},
  {32'hc2da53cc, 32'hc47d92a3, 32'h436348c0},
  {32'h44d3811f, 32'h4405a6b1, 32'h43790fc6},
  {32'h42d76198, 32'hc3abbdb8, 32'hc44a77c4},
  {32'h451999b5, 32'h44915c54, 32'h4335c103},
  {32'hc460caae, 32'hc4956e35, 32'h43a0908d},
  {32'h444d511b, 32'h4457f4e9, 32'h43141a52},
  {32'h436cdd08, 32'h4389a5b8, 32'hc47dfe36},
  {32'hc3d475c4, 32'hc42f8f64, 32'hc5173cc8},
  {32'hc3025b3c, 32'hc2f6effb, 32'h43c83ca1},
  {32'h451421e0, 32'h43f541cb, 32'h4292b638},
  {32'h42a7e6a8, 32'hc5510dac, 32'h42d5c697},
  {32'h41d119f2, 32'h42bcc56b, 32'h44d803c2},
  {32'hc3dd6b35, 32'hc4733d8d, 32'hc450656d},
  {32'h41a0b300, 32'h44388022, 32'h449c0b84},
  {32'h43174626, 32'hc485b9e7, 32'hc2e73d51},
  {32'h443445f8, 32'h44765abc, 32'h44218a0a},
  {32'hc441dd2d, 32'h439e190c, 32'hc4beaebc},
  {32'hc37fdb95, 32'h440130be, 32'h422e6d68},
  {32'hc51f4e34, 32'h43acbd1a, 32'hc426c3fb},
  {32'hc322cd60, 32'hc309ac4d, 32'h4521ec69},
  {32'hc32d9dc7, 32'hc4868826, 32'hc3a25e51},
  {32'h4346b1e6, 32'h4514284f, 32'h43652a17},
  {32'hc555ec72, 32'hc3e1f56e, 32'hc3ae872f},
  {32'h433df2cd, 32'h44177729, 32'h445799a3},
  {32'hc4b4f88a, 32'hc3cabbd8, 32'hc3b43ef0},
  {32'hc46138ae, 32'hc47853ed, 32'hc3852529},
  {32'hc3393640, 32'h450bbac2, 32'h4434ea56},
  {32'hc51a1260, 32'hc3882889, 32'h43a8f4d6},
  {32'h430036d8, 32'h452b8272, 32'h428354ca},
  {32'hc5214d6d, 32'hc33c1bc7, 32'hc31f89c7},
  {32'h44bd6ad8, 32'h439edd73, 32'hc3bbc97a},
  {32'hc3cad38c, 32'hc3a501fb, 32'hc31b15f4},
  {32'hc4056028, 32'h43e50c46, 32'h43eceac8},
  {32'h43b92564, 32'hc413ed63, 32'h444e5b89},
  {32'h4376b766, 32'h44f4ae47, 32'h43831568},
  {32'h42a0f216, 32'hc52b10c5, 32'hc360e906},
  {32'h44b47f76, 32'h43a5f102, 32'h43076e1e},
  {32'hc43714ea, 32'hc503d524, 32'hc381a575},
  {32'h448d90c8, 32'h44839b9e, 32'hc40aa4d8},
  {32'h44a036c4, 32'hc2211eb6, 32'h43613f86},
  {32'h44de4004, 32'h438d169f, 32'hc333d76a},
  {32'hc48cef11, 32'h41a45902, 32'h441ce726},
  {32'hc16a639a, 32'h441ab17e, 32'hc38e14c6},
  {32'hc43107a6, 32'hc489fb79, 32'h44ae51bf},
  {32'h43b01057, 32'h4559e04e, 32'h430af2e1},
  {32'hc3839d8b, 32'h42fe3e9e, 32'h44c2ba36},
  {32'h428caf20, 32'hc30b9d73, 32'hc44249c0},
  {32'h43a3c2b8, 32'h41913cc7, 32'h451ef010},
  {32'h425ec08e, 32'h43f87064, 32'hc304b1f8},
  {32'hc4f228d6, 32'h438988c8, 32'h445bc756},
  {32'h454343ac, 32'hc3a0905c, 32'hc48d6c98},
  {32'h43f06420, 32'hc50f9cc2, 32'hc21f3d74},
  {32'h4338d3ea, 32'h4524e838, 32'h42a681ec},
  {32'hc24f2d58, 32'hc43f826d, 32'hc3d1eada},
  {32'hc499f3ba, 32'h44af73d5, 32'h437fe086},
  {32'h44f042c7, 32'hc41343f9, 32'hc309f5f6},
  {32'h43e04dd2, 32'hc3043ae4, 32'hc2a202b0},
  {32'h44c411dd, 32'h4427f068, 32'hc32883c5},
  {32'hc568d6d7, 32'h43aa94ea, 32'h440f6243},
  {32'hc4951d70, 32'hc393958d, 32'h41ea1f3c},
  {32'h434eb384, 32'h42d2d79c, 32'h443b396f},
  {32'h448c834e, 32'hc3995d98, 32'h44974b13},
  {32'h442dcab9, 32'h4130ed44, 32'hc35c3fba},
  {32'hc3a5a3a2, 32'hc481cfb6, 32'h44452f75},
  {32'hc3ff1a70, 32'h44b77275, 32'hc305a18c},
  {32'hc4845aa7, 32'hc446e74a, 32'hc39df21c},
  {32'hc429986e, 32'hc3b57e73, 32'hc482e47c},
  {32'h446ee236, 32'h42b5c886, 32'h4491e4ff},
  {32'hc46637a2, 32'hc30c6f22, 32'hc471ecc3},
  {32'h44831e25, 32'hc43a3faf, 32'h448e312b},
  {32'hc30162f0, 32'h4504139d, 32'hc44c77ee},
  {32'h439e44fd, 32'hc44ec057, 32'h441e14a4},
  {32'hc3d6d397, 32'h452c3a8c, 32'hc32be95e},
  {32'h451ab2bc, 32'h44067e66, 32'h43c28161},
  {32'h44ba7260, 32'hc38f2503, 32'hc349da80},
  {32'h44c46081, 32'h4303049b, 32'h44e35c68},
  {32'hc49e9644, 32'hc42e6afd, 32'hc505820a},
  {32'h43ed67e6, 32'hc330529e, 32'h43bda153},
  {32'h4193e8da, 32'hc50f1c30, 32'hc4dde25d},
  {32'h43b4a07c, 32'hc5118973, 32'h44b60c6b},
  {32'h44c33f10, 32'h435e67f7, 32'hc44a34fb},
  {32'hc435cbb0, 32'h4335aa2b, 32'hc3a56078},
  {32'h453bb652, 32'hc42b192b, 32'h43c98bc5},
  {32'hc44ec532, 32'h4205d838, 32'hc4614bcb},
  {32'h452b3b00, 32'h43fe62bd, 32'hc41102f1},
  {32'hc4032153, 32'h448320a6, 32'hc527a36e},
  {32'h4461d523, 32'hc472c366, 32'h43ea8d3d},
  {32'h44341df5, 32'hc42c13f0, 32'h44991905},
  {32'hc418f13c, 32'hc40dabec, 32'hc495d09e},
  {32'h440f75b7, 32'h43ff77ec, 32'h43485260},
  {32'h4460ff25, 32'hc42027eb, 32'h4381efc7},
  {32'hc4b799fa, 32'h43e29d89, 32'hc3ad6066},
  {32'h4424bf18, 32'hc473b44f, 32'hc3736f0c},
  {32'hc42ccba0, 32'h444b0778, 32'h43e8ba9c},
  {32'h451b35bc, 32'hc3b8ae9c, 32'hc2c67816},
  {32'hc324710a, 32'h44225fbd, 32'hc4c61961},
  {32'h449cd8ab, 32'hc3e1c569, 32'h433b51d6},
  {32'hc52d2100, 32'hc41c1acb, 32'hc37bf556},
  {32'hc3972e87, 32'h44021549, 32'hc324f96d},
  {32'h43431e07, 32'h44f4c8c4, 32'h43b5a862},
  {32'h438d7152, 32'hc5762c8f, 32'hc2291074},
  {32'hc4ac0e83, 32'h449450d0, 32'hc39df4cf},
  {32'h45507f2d, 32'h4340556a, 32'hc128346e},
  {32'hc4acf53a, 32'h44bbc144, 32'h439d3edc},
  {32'h43ec7b9f, 32'hc4a1a78f, 32'hc352b1fb},
  {32'hc3b8ced4, 32'h429e9fc5, 32'h440199cc},
  {32'hc39e4b28, 32'hc4882f6f, 32'hc53e5a04},
  {32'h43045398, 32'h448d5da4, 32'h44e5e6cd},
  {32'hc37887a8, 32'hc2d9e4bc, 32'h43df5d24},
  {32'h43762274, 32'h44dff5c8, 32'h41be6216},
  {32'h43808b18, 32'hc322b3f4, 32'h44610d63},
  {32'h44bdd7e4, 32'h4464f8e4, 32'hc432355c},
  {32'hc45f2c54, 32'h4323b0f3, 32'h44635201},
  {32'hc323a116, 32'h44c0fa81, 32'h43ccc0b4},
  {32'hc3a9f66c, 32'h438eccf2, 32'h4333a5f4},
  {32'hc3ae6b62, 32'h44a598cc, 32'h44b9965b},
  {32'h4205042d, 32'hc48d220f, 32'hc512fe3d},
  {32'h442cf7f0, 32'h43c2dbd2, 32'hc4872883},
  {32'hc408e17c, 32'hc50d26db, 32'h43258e6d},
  {32'h42ce46a3, 32'h42e59aad, 32'hc4fbab85},
  {32'hc3ec67ce, 32'hc405d5dd, 32'h448b6d33},
  {32'h448369c0, 32'h449bd900, 32'hc3f373b1},
  {32'h4453f01a, 32'hc3bb1fce, 32'h443cd597},
  {32'h449c50ee, 32'hc2491002, 32'h439c85bc},
  {32'hc518f371, 32'h4399d301, 32'hc27c8ed3},
  {32'hc4ce9a94, 32'h43cff4f8, 32'h4373b324},
  {32'hc4750e5a, 32'hc49c8152, 32'h43be0e94},
  {32'h4500d588, 32'h444a522d, 32'hc2bc94b7},
  {32'h423e82a0, 32'hc4312691, 32'h438a7051},
  {32'h45565584, 32'h4408e0bf, 32'h41f5cebe},
  {32'h43c893f4, 32'hc57291f2, 32'h431f47d2},
  {32'h43b58b3d, 32'hc293f430, 32'hc2f2c532},
  {32'h43c82cc4, 32'h4301f284, 32'hc085947a},
  {32'h43d4d76e, 32'hc4b24a39, 32'hc28b9397},
  {32'hc3ca0d84, 32'hc4e7b590, 32'h44daef82},
  {32'h43dea0d3, 32'hc3009aef, 32'hc42bcdf8},
  {32'hc32e9756, 32'h455c52bc, 32'hc2082d21},
  {32'h42ea24a6, 32'hc5127b90, 32'hc2f8f44f},
  {32'hc3fdd7ae, 32'h43bac676, 32'h4398f239},
  {32'hc46752e0, 32'hc41197c3, 32'hc4d2d2c5},
  {32'hc418893a, 32'h44534dc3, 32'h4568c851},
  {32'hc3c495ce, 32'hc428ea72, 32'h43592839},
  {32'hc306f09a, 32'hc502876e, 32'h44a626df},
  {32'hc444a624, 32'hc4678cd7, 32'hc40f889f},
  {32'hc1ae2670, 32'h4442c7d2, 32'h441cd8f8},
  {32'hc1d0345c, 32'hc5229f6d, 32'hc3c9b56a},
  {32'h44f1e852, 32'h43a6b4ce, 32'h4393eb84},
  {32'h444079e3, 32'hc3a6c623, 32'hc4409ce3},
  {32'h451fb95d, 32'h43887ab7, 32'hc2647202},
  {32'hc4a8a456, 32'h42009b7e, 32'hc44e9baf},
  {32'h42783f28, 32'h44b77c23, 32'h4346c851},
  {32'hc3902260, 32'hc509b7c5, 32'hc3acbad6},
  {32'h44ee4ff3, 32'h446c6178, 32'hc30bef91},
  {32'h44599b16, 32'hc34df5cd, 32'hc3a9dc6a},
  {32'hc3275e0f, 32'h453dbc34, 32'hc0d123b0},
  {32'hc40074aa, 32'hc5824eb2, 32'h43ac5589},
  {32'h45215e99, 32'h4434235a, 32'h43add475},
  {32'hc4cab750, 32'h43513cda, 32'hc374fcf3},
  {32'h43240628, 32'h43390a01, 32'hc3d3b928},
  {32'h4343a660, 32'h43e0f845, 32'hc4a52bdb},
  {32'hc31c2062, 32'h45058214, 32'h446ec787},
  {32'h43c546cd, 32'hc2913c74, 32'h43a94ae7},
  {32'hc30c4049, 32'h443bde2f, 32'h445c489f},
  {32'h4371672d, 32'hc50e6a24, 32'hc3cfc28a},
  {32'h422abea9, 32'hc41f9f27, 32'h434efb33},
  {32'h4545f598, 32'h4263d911, 32'hc37a20dd},
  {32'hc4e94305, 32'h4401740d, 32'h443dbc97},
  {32'hc4b706ca, 32'hc39d0c05, 32'hc3a4daab},
  {32'h42422bf0, 32'hc40351f0, 32'h44a8380a},
  {32'hc22826c0, 32'h4503dfd9, 32'hc4e1ee9e},
  {32'h43dfe2ad, 32'hc3447d8a, 32'h440cec37},
  {32'h4542ae80, 32'hc3fa9ef1, 32'hc05985bc},
  {32'hc4c45a04, 32'h430d3c3e, 32'h447c962d},
  {32'h4195dd14, 32'hc49f8d37, 32'hc3bd3cef},
  {32'hc3d718bf, 32'h441fa60e, 32'h44e43aa6},
  {32'h4497fba6, 32'h443818f9, 32'hc459b8cb},
  {32'h44202dc6, 32'h445c8afd, 32'h44978e2e},
  {32'h45020e37, 32'hc4170b00, 32'h41f7a7a1},
  {32'hc4fd5420, 32'h43c7f63f, 32'h44510326},
  {32'h44513734, 32'hc3c3ad46, 32'h43e7dd5c},
  {32'hc50e06b2, 32'hc34534f0, 32'h419c38b2},
  {32'h4459e14c, 32'hc4a3411a, 32'h4304d8f5},
  {32'h44b29a88, 32'h43a7eaa1, 32'hc09a48f0},
  {32'h44de2690, 32'hc35af503, 32'h436d59e7},
  {32'hc54dc1d5, 32'hc3249947, 32'hc40ef301},
  {32'hc451090f, 32'hc3a62e94, 32'hc3e7e151},
  {32'hc425f5e8, 32'hc3a8c9f9, 32'h44a15679},
  {32'hc4aed68b, 32'hc34b104a, 32'h435ffdd6},
  {32'h449ca568, 32'hc2b1cffd, 32'h43d95df3},
  {32'hc3a3243e, 32'h447e651c, 32'hc3911494},
  {32'h444be8ed, 32'hc4d573ae, 32'hc3a9a514},
  {32'h4126a500, 32'h43ea8ce9, 32'hc4208411},
  {32'hc4d71f6a, 32'hc365cc70, 32'h421ab0cd},
  {32'hc4a63023, 32'h44944a79, 32'hc350e51a},
  {32'h445eb070, 32'hc4826f01, 32'hc2a9f8bb},
  {32'h43fa326e, 32'hc1275746, 32'hc49a14a8},
  {32'h442f7bf2, 32'hc3c41a4b, 32'h450cddb5},
  {32'hc4ff7987, 32'hc404fb82, 32'h43c54377},
  {32'h451b9678, 32'h43a41d3c, 32'h43aa4cfb},
  {32'hc3809358, 32'hc373227d, 32'h450e08b7},
  {32'h4484cef0, 32'hc478b08b, 32'hc390e831},
  {32'h42cf5eb2, 32'h4508e845, 32'hc31b33e6},
  {32'h449c5e30, 32'h444f04ed, 32'hc4375df7},
  {32'hc4bd6bf7, 32'hc2494c9c, 32'h449c1e78},
  {32'hc4d00a20, 32'hc3035c43, 32'hc3d6c95f},
  {32'hc51a7ebd, 32'hc3302bfe, 32'h4403586b},
  {32'h44364b10, 32'h44768e62, 32'hc3a45493},
  {32'hc32496a6, 32'h44e871c7, 32'h4381e227},
  {32'h42f3aed0, 32'hc4665532, 32'hc41acd51},
  {32'hc50e092b, 32'h42299db7, 32'h43de4712},
  {32'h44d85115, 32'hbf721cc0, 32'hc2f3bdd7},
  {32'hc31aec58, 32'h4499d626, 32'h44a8da1b},
  {32'h4498f563, 32'hc4be1452, 32'hc40427ab},
  {32'h45146026, 32'h43b897ec, 32'hc459b08f},
  {32'hc4b3316a, 32'hc320c377, 32'h44b9a70a},
  {32'hc1844133, 32'hc1f6f80e, 32'hc44bd897},
  {32'h41f59566, 32'hc552f555, 32'hc3bbc3b2},
  {32'h447d1c05, 32'h44bce943, 32'h43b384ce},
  {32'h4467d4eb, 32'hc401d005, 32'hc35c6493},
  {32'h4325c69a, 32'h4493c8ea, 32'hc2621fd0},
  {32'hc506c1ce, 32'hc4450a20, 32'h43757da1},
  {32'h4335534c, 32'h44920fde, 32'h440d3f60},
  {32'hc2dc9f80, 32'hc3e870fa, 32'h4462f40e},
  {32'h44045da6, 32'h40ea473d, 32'hc499c425},
  {32'hc45962aa, 32'hc3ec6fd6, 32'h44a50436},
  {32'h44ac955b, 32'h4341e9e0, 32'h44d2414b},
  {32'hc446a735, 32'hc464789e, 32'hc3a4dc0b},
  {32'hc2c327c6, 32'h432a2600, 32'h4497db9f},
  {32'hc215b080, 32'hc5382234, 32'h43b6b011},
  {32'hc17dda10, 32'h43c5b4c2, 32'h453fc6b5},
  {32'h407d4ea5, 32'hc48697b4, 32'hc40b1292},
  {32'h4528dab1, 32'hc3577ba4, 32'h4250d383},
  {32'hc4af2247, 32'hc495ca73, 32'hc4b624db},
  {32'h44803cc0, 32'h434648a1, 32'hc388e4ba},
  {32'hc431cda5, 32'hc3d75d5a, 32'hc4094c6b},
  {32'h42d4cd14, 32'hc3cf2d34, 32'h4414c55f},
  {32'h44b6f399, 32'hc2634768, 32'hc3b68524},
  {32'h44f8f2ff, 32'h43cb0315, 32'h443f344e},
  {32'hc43c3901, 32'hc351ee0c, 32'hc542de7c},
  {32'h44ebff84, 32'hc354e131, 32'hc33e00f0},
  {32'hc49e6ada, 32'h43d72b2f, 32'hc34bb191},
  {32'hc51e8287, 32'hc345d81b, 32'hc21e114e},
  {32'hc2a15a8e, 32'h43e39ba7, 32'h4489621c},
  {32'hc4669678, 32'h436444b0, 32'h44203ed9},
  {32'h440a4c10, 32'h4496b1c8, 32'hc43bad72},
  {32'hc49d2008, 32'hc4d1039b, 32'hc3caef37},
  {32'hc4659d9e, 32'hc2e5be1e, 32'h436c5090},
  {32'hc5563738, 32'hc336ef51, 32'hc33f10f9},
  {32'h44ae1254, 32'hc3130499, 32'h443be37d},
  {32'h44564a0e, 32'hc1c68966, 32'h43c1f203},
  {32'h425cbd39, 32'h452e1f03, 32'h43bcd74d},
  {32'hc409be43, 32'hc362516c, 32'hc408367d},
  {32'h435c4cd0, 32'h44b41773, 32'hc3ab0514},
  {32'hc4c57e9a, 32'hc3eed23a, 32'h436b26d3},
  {32'hc37d73b8, 32'hc2eb3cde, 32'hc51625aa},
  {32'h44dbe3aa, 32'h40e31504, 32'h4303395e},
  {32'h4442b044, 32'hc3a227fd, 32'hc50b521d},
  {32'hc4877226, 32'h42d947bc, 32'h448e7a22},
  {32'hc48eaf03, 32'h43c2d958, 32'hc2acf0f4},
  {32'hc446205a, 32'hc4b2afac, 32'h43cd4440},
  {32'h44f28b16, 32'h43f259d3, 32'hc472e11d},
  {32'hc46e71a2, 32'hc2301fbc, 32'h433b4a96},
  {32'h445c54aa, 32'h445f121a, 32'hc404bc70},
  {32'hc2147166, 32'hc516a59b, 32'h44160b8d},
  {32'h453b254e, 32'h43d5481e, 32'h4287ad28},
  {32'hc3d14438, 32'h43842d87, 32'h45280063},
  {32'h454957f8, 32'h42df7cff, 32'hc45655ec},
  {32'h4412cbf4, 32'hc4503c4b, 32'hc4751520},
  {32'hc44fa38e, 32'h44bdc529, 32'h43cbadf6},
  {32'hc491cb44, 32'hc4162e5e, 32'h431cee75},
  {32'hc4dd7d19, 32'h441a809e, 32'hc3440268},
  {32'h442cf61c, 32'hc4f19832, 32'hc343f9ac},
  {32'hc4b83c79, 32'h43873cc3, 32'hc32754d2},
  {32'h44481434, 32'h42f1d130, 32'h4384586d},
  {32'hc4e533de, 32'hc46d2bc4, 32'h43f1d1b2},
  {32'hc4ac3129, 32'hc258ae4a, 32'h4377d590},
  {32'hc405ae12, 32'h4405b80d, 32'hc3ce2974},
  {32'h4394f2f8, 32'hc30f7f1d, 32'hc399cfe5},
  {32'h4358b00a, 32'h449a0bc4, 32'h43a1cb46},
  {32'h4424a2c0, 32'hc4948e58, 32'h406c5020},
  {32'h4352593d, 32'h45304f0b, 32'h43d0eefa},
  {32'hc3abe187, 32'hc4baa841, 32'hc3543058},
  {32'hc4bca438, 32'h436935df, 32'hc20802a5},
  {32'h430dc4a2, 32'h4313be48, 32'h4472adf5},
  {32'h43540ee4, 32'h4432d910, 32'hc2a1d50c},
  {32'h42320005, 32'hc540f0a7, 32'hc42e0bf3},
  {32'hc47c8868, 32'h41af8c84, 32'hc3aa623f},
  {32'h44f3c85e, 32'h435d2f95, 32'hc3b03637},
  {32'hc46add7f, 32'h43f5f9db, 32'hc506802d},
  {32'h441123b6, 32'hc4465bbf, 32'h440e0b96},
  {32'hc515c7d9, 32'hc1b6f612, 32'h435dff40},
  {32'h44a92d39, 32'h422d03db, 32'h4483420a},
  {32'hc41b9e53, 32'hc4046982, 32'hc531e85c},
  {32'hc3ec7392, 32'hc306f3de, 32'h43e7a245},
  {32'h4275fdc4, 32'h438bcc08, 32'hc49c37a7},
  {32'hc47764c8, 32'h43890e07, 32'h4420dcb3},
  {32'h433cc310, 32'h4453327e, 32'h4327d1bc},
  {32'hc4048903, 32'h439941e2, 32'h42023e23},
  {32'h4463e402, 32'hc37f08f8, 32'h4486ba53},
  {32'h436668b4, 32'h451ce2c0, 32'hc250250b},
  {32'h43d2862c, 32'hc4b556d8, 32'hc38eff22},
  {32'hc48f7479, 32'h43ce4624, 32'hc4a4a2a7},
  {32'hc3b51388, 32'hc3822acd, 32'h455c2a09},
  {32'h43a51ec0, 32'hc47bf873, 32'h44fb46bb},
  {32'h4382a104, 32'hc50f8593, 32'hc4ac74f9},
  {32'h43e178d8, 32'h435cc140, 32'h44463d7b},
  {32'h42093f74, 32'h427e3286, 32'h44da12b3},
  {32'hc39883d4, 32'h44c6e024, 32'h42b05df9},
  {32'h44f07aa0, 32'hc33576fe, 32'hc3c180e6},
  {32'hc41737ea, 32'hc37f8fd2, 32'hc4a8076d},
  {32'h447add62, 32'hc48cc78a, 32'h4422d5a5},
  {32'hc46da05d, 32'h441a73f8, 32'hc455c405},
  {32'hc4c2983e, 32'hc3c14a3b, 32'h42be10fa},
  {32'hc4c510bc, 32'hc489b045, 32'hc461d143},
  {32'h449685b2, 32'h4337b703, 32'hc39b8f7f},
  {32'hc4963320, 32'hc3fa46d7, 32'hc095000e},
  {32'hc374bdd0, 32'hc5498298, 32'h41e1b3d1},
  {32'hc5091f73, 32'h444c6446, 32'hc3ae41f0},
  {32'h43ce7852, 32'hc4c11bc3, 32'hc22d485a},
  {32'hc58f04ba, 32'h4197a144, 32'hc382e5d1},
  {32'h454a078d, 32'hc4288c5a, 32'h4323e904},
  {32'hc340e10c, 32'hc2e4ff8f, 32'h439f0ba0},
  {32'h43066c9c, 32'hc42b08f8, 32'hc4dfe281},
  {32'hc4a2436c, 32'h4407d526, 32'h446cb1d5},
  {32'h43b850d8, 32'hc48c572a, 32'h44a0f6ad},
  {32'h44ad93f4, 32'h43fb74fc, 32'hc3de8f90},
  {32'hc4b992be, 32'hc401387f, 32'hc31695f6},
  {32'h45151f81, 32'h439fb50c, 32'hc1b89ac6},
  {32'hc515b36e, 32'hc310b0ef, 32'h434facd6},
  {32'hc45b3c4e, 32'h4122f538, 32'hc49bdb46},
  {32'hc4027f98, 32'h443bbfdb, 32'hc41019e0},
  {32'hc487cea8, 32'hc43dfbb5, 32'h44b90e1e},
  {32'h43bce575, 32'h42921efe, 32'hc49032ea},
  {32'h44f58f90, 32'h43c5f7a5, 32'hc3244acf},
  {32'hc530e4d1, 32'hc41aede4, 32'h4325d4a3},
  {32'h43a7bbed, 32'hc1aa46ee, 32'hc4b9805f},
  {32'hc33cb0fc, 32'hc4caa888, 32'h4460f433},
  {32'h441d32f5, 32'h4367abff, 32'hc4e37aa9},
  {32'hc391695f, 32'hc45b2fac, 32'h437e1374},
  {32'h444cc766, 32'h441a2519, 32'hc00a9156},
  {32'hc4bf3592, 32'hc365e9c3, 32'h43d14a61},
  {32'h454f4a44, 32'h438e571e, 32'hc1e0a218},
  {32'hc49f5664, 32'hc4ad457c, 32'h43b32d35},
  {32'h44651a21, 32'h4428e1d5, 32'h41f873d9},
  {32'hc4728ae2, 32'hc3ddd6b3, 32'h4366e25d},
  {32'h43da0044, 32'h44a2e4b1, 32'h43c164d0},
  {32'h43ce4738, 32'hc5504e86, 32'hc3154a5e},
  {32'hc4a98290, 32'hc36e10ba, 32'h4374b05c},
  {32'hc421409c, 32'hc408806d, 32'h43cfd3ac},
  {32'hc1c8fe80, 32'hc3c7c7a7, 32'hc4484b31},
  {32'h44b863af, 32'hc4004e39, 32'h440488c1},
  {32'hc3481bd6, 32'hc3a12c9b, 32'hc24c5b9d},
  {32'hbe4cd000, 32'h42e9c422, 32'h45001af7},
  {32'h41e20f90, 32'hc3a441a7, 32'hc5449214},
  {32'hc3500ca7, 32'h443cc344, 32'h449148d7},
  {32'hc37f9c76, 32'h433be052, 32'hc48b648e},
  {32'h448a45ee, 32'h44601df3, 32'h446647bd},
  {32'h43eea406, 32'hc4337e57, 32'h416d06a6},
  {32'h43a634b8, 32'h4502c070, 32'h43e5dae2},
  {32'hc406f280, 32'h4358d214, 32'hc49212b6},
  {32'h44a63b10, 32'h41b82292, 32'h43b9d713},
  {32'hc406948e, 32'hc37ae32f, 32'hc4ac3a68},
  {32'h44d1820c, 32'h42f7a4de, 32'hc2fa130c},
  {32'h44b65cfb, 32'hc2b83ac9, 32'h435dfabb},
  {32'h45624cf4, 32'h42e98776, 32'hc2635c06},
  {32'hc424f706, 32'hc45bbb31, 32'hc3d66bc4},
  {32'h438d9c41, 32'h44579c7f, 32'h4362556a},
  {32'hc55da966, 32'hc43b11cb, 32'hc316ddd0},
  {32'h446034fa, 32'h45012de4, 32'hc38761aa},
  {32'h44bbb2c3, 32'hc0abde33, 32'hc27d5644},
  {32'h44023979, 32'h43ac149c, 32'hc3c982c3},
  {32'hc431f49c, 32'hc40a6533, 32'h42cada0a},
  {32'h43af4a41, 32'h43339eeb, 32'h4396c631},
  {32'hc570db03, 32'hc325ecb0, 32'hc421e885},
  {32'h45809617, 32'hc3c9d8ca, 32'hc236cc18},
  {32'h443ee87a, 32'hc509f95e, 32'hc46bb548},
  {32'hc4d30307, 32'hc3ff0df4, 32'h4430db65},
  {32'hc40cdbcd, 32'hc2540384, 32'hc3f74385},
  {32'hc4c1de4d, 32'h4230abce, 32'h43a23625},
  {32'hc377e7aa, 32'hc451ccb3, 32'hc45ac0f7},
  {32'hc308fb60, 32'h43547a54, 32'hc2a1f419},
  {32'h4375a028, 32'hc48390b9, 32'hc4a8b1d7},
  {32'hc4bc2360, 32'h4427c972, 32'h4456ca04},
  {32'hc3cf1392, 32'h4397eaa3, 32'hc35fd94c},
  {32'h4472c23e, 32'hc4e6a37e, 32'h450de0d5},
  {32'h450dd2be, 32'h439edf59, 32'h43baae9c},
  {32'hc4ed70db, 32'hc3a3e109, 32'hc357f759},
  {32'h431bd3d7, 32'hc51f3a5a, 32'hc4814de1},
  {32'hc41101ac, 32'h45117a8d, 32'h444694f5},
  {32'h43c6aa64, 32'hc418406b, 32'hc3af8931},
  {32'hc382d6df, 32'h43dff7bb, 32'h44c0dbc7},
  {32'h42fa5420, 32'hc3492dfb, 32'hc4a64319},
  {32'h42ece3d0, 32'hc37ffb1f, 32'h44abc8aa},
  {32'h44f522bc, 32'hc495f958, 32'hc3b7a214},
  {32'hc4ef9300, 32'h449a7e14, 32'hc351897b},
  {32'hc18abf60, 32'hc48abad0, 32'hc3cd219f},
  {32'h433694e1, 32'h43e7d4fb, 32'hc3a2f679},
  {32'h45127fb7, 32'hc43fd307, 32'hc29fbd2e},
  {32'hc444d0db, 32'h441b919b, 32'h4381a9c0},
  {32'h434419f0, 32'hc3e42c24, 32'hc3d56d9c},
  {32'hc410527e, 32'hc1e98d88, 32'h4190b524},
  {32'hc4eb3f7e, 32'h42003de5, 32'hc21ce42b},
  {32'hc3b6ad6c, 32'hc40b4bcb, 32'h432e5480},
  {32'hc5117216, 32'h432fb025, 32'hc45dc2fc},
  {32'h43059570, 32'hc36ef687, 32'h44db9f89},
  {32'hc50b19e3, 32'hc3fb850f, 32'hc22584c8},
  {32'h436845fc, 32'hc3bc8852, 32'hc352eae2},
  {32'hc523e65c, 32'h445b9ba2, 32'h42b5ecc3},
  {32'h45402ab6, 32'h44187716, 32'hc4002ad8},
  {32'hc50f9cab, 32'h434b951c, 32'hc2b21e21},
  {32'h44023eef, 32'hc5278c34, 32'h434a1095},
  {32'hc4c10ae9, 32'hc3bff6fb, 32'hc3d4074f},
  {32'h4431ca3b, 32'h418253ae, 32'h4503f128},
  {32'hc43b5b8c, 32'hc2acd4b9, 32'hc48ed9f2},
  {32'h4422e284, 32'hc439cfa3, 32'hc44282a5},
  {32'hc451d9cb, 32'hc377c1c2, 32'h44406c62},
  {32'h443520a1, 32'hc4727ddf, 32'hc42c4cf8},
  {32'hc492583d, 32'h4443e8dd, 32'hc347f437},
  {32'hc3b5f8ec, 32'h42e51773, 32'hc523226e},
  {32'hc43d026b, 32'h43b57937, 32'h44a59347},
  {32'h454faa42, 32'h438934c6, 32'hc3fad62f},
  {32'hc4e6642a, 32'h44262d3f, 32'h448776d7},
  {32'h44b1c2d1, 32'hc292aab2, 32'hc41a8cf2},
  {32'hc50bd7f2, 32'h43a64ad6, 32'hc3e8397a},
  {32'h43e889ce, 32'hc5284be6, 32'h42a63a7f},
  {32'hc380f5b0, 32'h44cd9efc, 32'h43d5c6e6},
  {32'h453378c4, 32'h42a3091b, 32'hc3173fea},
  {32'hc2bfe3a3, 32'h4542c9b2, 32'h434651d0},
  {32'h439f8446, 32'hc4d6e2f1, 32'hc34f9665},
  {32'hc366778b, 32'hc2031cdb, 32'hc514941d},
  {32'hc4272330, 32'h42965cb7, 32'h45326005},
  {32'h4549fa19, 32'h438276ac, 32'h43f485fc},
  {32'hc3acba47, 32'hc4e573c3, 32'hc394ce13},
  {32'h44e4222c, 32'hc22b96f2, 32'h4241c976},
  {32'hc3afb20c, 32'h43702ade, 32'hc36b4c82},
  {32'h42e5b550, 32'h450b39ab, 32'hc38c6d27},
  {32'hc249fa90, 32'hc52ce4fd, 32'hc3eb3716},
  {32'hc39422e3, 32'h44de77ec, 32'hc3895030},
  {32'hc497bbcd, 32'hc3521d7d, 32'hc4299b80},
  {32'h4539f4a2, 32'hc3533738, 32'h433206db},
  {32'hc4af0902, 32'hc400cb08, 32'h439d1ef0},
  {32'h4351deda, 32'h4513f3ac, 32'h441ae418},
  {32'hc47ad9a2, 32'hc4088870, 32'hc526a5be},
  {32'h40ebcc80, 32'h4443845d, 32'h430e51d2},
  {32'hc4429df6, 32'hc4cd999b, 32'h42a88867},
  {32'h430e7659, 32'hc16222fa, 32'h4491d98a},
  {32'hc3cb568d, 32'hc4804ca2, 32'h43bf9ad5},
  {32'h4543e2fc, 32'hc3144f1b, 32'h443ef705},
  {32'hc4ff0811, 32'hc2e3e6f4, 32'h4135a635},
  {32'hc485f703, 32'h43907058, 32'h430bab15},
  {32'hc4f5412b, 32'hc49b010a, 32'hc279d9b7},
  {32'hc2e57390, 32'h432c7b54, 32'h452afe60},
  {32'hc2b412d6, 32'hc396b311, 32'hc43a6903},
  {32'hc3112d2a, 32'h43cf0714, 32'h450e1efe},
  {32'hc4123b2c, 32'hc2d192af, 32'hc53d83fc},
  {32'h453a67c7, 32'hc328f814, 32'hc3b39422},
  {32'hc4337e0c, 32'h44818041, 32'hc367a7be},
  {32'h4386decc, 32'hc506c0df, 32'hc2bb31cd},
  {32'h44418d54, 32'h44be1ed4, 32'h444186e6},
  {32'hc53cf9b9, 32'h43435600, 32'hc2a80a6b},
  {32'hbd080000, 32'h4460ab2e, 32'h442c75ba},
  {32'h40809200, 32'hc56042ec, 32'h43b5b64b},
  {32'hc37e84a8, 32'hc304e440, 32'h43b50cef},
  {32'hc53e135c, 32'hc2b075a2, 32'hc381f5f3},
  {32'h44d887d8, 32'h44147b92, 32'h43e5b01a},
  {32'h43876bae, 32'hc4995dd0, 32'hc35a344a},
  {32'h44db0873, 32'h43d22fa5, 32'h426d39ea},
  {32'hc4cba350, 32'hc3768df5, 32'h43c9add9},
  {32'hc34c3ed8, 32'h43cf68be, 32'hc50f4027},
  {32'hc4a8a09a, 32'hc40e85f4, 32'h42d831fc},
  {32'h42b3a350, 32'hc19b835b, 32'hc4bf3510},
  {32'h44df7721, 32'hc3439f1d, 32'h43930532},
  {32'h44290c7b, 32'h431ab6a7, 32'hc4db0c5f},
  {32'hc3234ee0, 32'hc49c9733, 32'hc433d9ff},
  {32'h44944f66, 32'h441e5c00, 32'hc38087ad},
  {32'hc4198652, 32'hc480ab4b, 32'h441097ff},
  {32'h441fe399, 32'h453547be, 32'hc2883d3f},
  {32'h44680706, 32'hc436e723, 32'h42660fcd},
  {32'h45189ab9, 32'hc3d55a77, 32'hc3518f26},
  {32'hc44e2c90, 32'hc4031922, 32'h4415e3af},
  {32'h45556b89, 32'h434072e0, 32'h43c4a2c7},
  {32'hc413d1e4, 32'hc2296a66, 32'h44981d56},
  {32'h454a22d7, 32'h43b40311, 32'hc418f658},
  {32'hc3260f8d, 32'hc551c94d, 32'hc408c961},
  {32'hc4a975a6, 32'h44ff9f23, 32'h4227c9a2},
  {32'hc3c587b2, 32'h434ae3a3, 32'h436f2dff},
  {32'hc538f199, 32'h44388288, 32'h439c23fc},
  {32'h43987fe9, 32'hc4de127b, 32'hc2ceba93},
  {32'hc4e73f22, 32'hc395dd92, 32'hc35963fc},
  {32'hc201ff9c, 32'hc42acb7e, 32'hc3ebd4e9},
  {32'h40bf2008, 32'h44031fd8, 32'h445de10e},
  {32'h442e5b07, 32'h42c51bb0, 32'h439976f5},
  {32'hc3b4a2f3, 32'h443da35f, 32'hc5192bcd},
  {32'h4209cd60, 32'hc50b630f, 32'hc2a4bf56},
  {32'hc3c30b00, 32'h43f6b270, 32'h432f8ad6},
  {32'h450f5daf, 32'hc4408b95, 32'h43c1586a},
  {32'hc4d1ae07, 32'h42b815e0, 32'hc49766d4},
  {32'h4511494f, 32'h43b11e43, 32'h43af16aa},
  {32'hc4a3dee1, 32'h4360d856, 32'hc3b44f80},
  {32'h44a5ad9c, 32'hc43ba28e, 32'h441b5c06},
  {32'hc1a89a00, 32'h4455853f, 32'h43e038a3},
  {32'h440d3db2, 32'hc49c102f, 32'h450a6910},
  {32'hc540a3b8, 32'h442a2bda, 32'hc31ba574},
  {32'hc409d8bc, 32'hc421bfc8, 32'h438ce52e},
  {32'hc52dab5d, 32'hc20166cd, 32'hc488907a},
  {32'hc2cfb168, 32'hc3fe38d3, 32'h453091a4},
  {32'hc32de2b8, 32'hc3d033c0, 32'hc4d91a2b},
  {32'h43bdc4b4, 32'h44626174, 32'h452eb7f9},
  {32'hc519777f, 32'h4299dbf5, 32'hc4475e30},
  {32'hc44d84e8, 32'h436b4252, 32'hc37cadf3},
  {32'hc373bde0, 32'h448af54f, 32'hc4c7d4a3},
  {32'h4502a38e, 32'h436a4aff, 32'h435a5119},
  {32'hc3c58aee, 32'h42b153de, 32'h4438564b},
  {32'hc3dc1be5, 32'h449f26a9, 32'h433c738f},
  {32'h43a22dd6, 32'h42fca535, 32'h441d741c},
  {32'hc3a63d4d, 32'h42017288, 32'hc4efab10},
  {32'h450b4b50, 32'h4311cf19, 32'hc38d1269},
  {32'hc441cf7f, 32'h4505e268, 32'h439fb871},
  {32'h421f98e0, 32'hc4fd3f8f, 32'h443a6f1c},
  {32'h42420810, 32'hc4cdf9b7, 32'h44e5126f},
  {32'hc298738c, 32'h4492044b, 32'hc4ff6888},
  {32'hc46e32ac, 32'hc300c802, 32'h4393658e},
  {32'hc26a3621, 32'hc2f9218f, 32'h41961030},
  {32'hc3e82044, 32'h44fc3786, 32'hc316ba15},
  {32'h4516ad94, 32'hc3dd9684, 32'h43c90b7c},
  {32'h43978e30, 32'h442f9aef, 32'h4365cf0f},
  {32'h443dd96c, 32'hc45defd6, 32'h4306da8e},
  {32'hc50678df, 32'hc24b686a, 32'hc31dba44},
  {32'h456d9056, 32'hc41b7667, 32'h43ebc335},
  {32'hc4fe3a33, 32'hc40e6159, 32'hc1f3786b},
  {32'h42c429c0, 32'hc3a2b8fa, 32'h431ef34b},
  {32'h43928547, 32'h44c43e64, 32'hc3af1d44},
  {32'h44d656a6, 32'hc4799521, 32'h43fa4498},
  {32'h424feaa0, 32'h45325bbf, 32'hc30f0e17},
  {32'hc4a37d63, 32'h4323a6d4, 32'h437847f0},
  {32'hc40e0e19, 32'h454bf6f1, 32'h43fa0c24},
  {32'h44c11d3e, 32'hc4a2dc48, 32'hc3540ce1},
  {32'hc377a83e, 32'h449fc8f1, 32'h4358bb09},
  {32'h448e9388, 32'hc322d971, 32'hc3948909},
  {32'hc3342a21, 32'hc514e075, 32'h44abb571},
  {32'hc444d7e3, 32'hc3229ad2, 32'h44e5f4c1},
  {32'h439799a4, 32'h4520aaac, 32'hc31c3a6c},
  {32'hc4257e98, 32'hc4a817d6, 32'h431dda4c},
  {32'hc0c3f9fc, 32'h4532a7df, 32'hc3082bd3},
  {32'hc395d35b, 32'hc4abd103, 32'hc306a310},
  {32'hc087f696, 32'h44d1e355, 32'hc3bb5fa5},
  {32'h444f1b0e, 32'h43e4b48a, 32'h42adda56},
  {32'hc3ac322c, 32'h44a873cc, 32'h44f6efe8},
  {32'h449ce196, 32'hc40389ab, 32'hc4066420},
  {32'h4459782c, 32'h442e7d6b, 32'hc2871261},
  {32'hc4380f35, 32'hc50d742c, 32'hc31b47b0},
  {32'hc3a23bb1, 32'h44610ddf, 32'hc43d7bc0},
  {32'hc4045c2c, 32'hc4db28e2, 32'hc308c9f4},
  {32'h4542e0d6, 32'h43503150, 32'h41158e28},
  {32'h438b6a7c, 32'hc3fb1467, 32'h43732626},
  {32'h4485c7cc, 32'h43d29c84, 32'hc3d8eb81},
  {32'hc4fdf340, 32'hc256dbcc, 32'h43200014},
  {32'hc49e108b, 32'h43902917, 32'hc39965c6},
  {32'hc4a28b51, 32'hc49fb982, 32'h439bb2d1},
  {32'hc289e3e2, 32'h44b816ae, 32'h434a9d18},
  {32'h445717b5, 32'hc2f2d079, 32'hc1f095b6},
  {32'hc2eebefe, 32'h45331678, 32'h43614cec},
  {32'h431a096c, 32'hc5502748, 32'hc3655c4b},
  {32'hc4912451, 32'h43c86e6c, 32'h438f89fa},
  {32'h449703fc, 32'hc40eb8fb, 32'h431a4983},
  {32'h4449a132, 32'h44cfa5d1, 32'hc487e183},
  {32'h451889c6, 32'h43ea7187, 32'h441f06f6},
  {32'h439bf826, 32'hc3d6f2d6, 32'hc44cd394},
  {32'h44316c95, 32'h44114b60, 32'h44968a8c},
  {32'hc3bf1494, 32'hc39b2db3, 32'hc454946d},
  {32'h439a71c0, 32'hc2831874, 32'h43b43071},
  {32'h432ae2a4, 32'hc4cbe125, 32'hc524f598},
  {32'h450d1d59, 32'h43807eaf, 32'h445b23d8},
  {32'hc2aaffa8, 32'h4480a5a4, 32'hc3aff53b},
  {32'h42c70d86, 32'h442e5e8a, 32'h43b0679d},
  {32'h40ddd6a0, 32'h4403c570, 32'hc3843d27},
  {32'h4418343d, 32'h42a47b61, 32'h43f7fc91},
  {32'hc5040112, 32'hc2c9b5c2, 32'hc32556f0},
  {32'h44549730, 32'h448d915b, 32'h43ccf512},
  {32'hc4376b7f, 32'hc464451b, 32'hc34a68a2},
  {32'h436980be, 32'h44cb7b3c, 32'h448cb2b1},
  {32'h442051b1, 32'hc498f240, 32'hc53ad685},
  {32'h44f99e1c, 32'hc3a8ab25, 32'h43ef2b60},
  {32'hc3993b20, 32'hc57ef78c, 32'hc30d7b01},
  {32'h43a394f8, 32'h453a3d58, 32'hc2b42830},
  {32'h42d7fa98, 32'hc442cecb, 32'h4357a787},
  {32'h43997e40, 32'h44358b79, 32'h43f77d25},
  {32'hc4d21a55, 32'hc3b6d0e2, 32'h43a9295d},
  {32'h44946b14, 32'h4411220f, 32'h43928a8b},
  {32'hc47939a2, 32'hc40fa465, 32'hc3084073},
  {32'h43ec5450, 32'hc4189404, 32'h43b9d89d},
  {32'h4386adc2, 32'h44a8bbdd, 32'hc518b7e1},
  {32'hc3da21f9, 32'h442a27cf, 32'h449331ef},
  {32'h44bf09d3, 32'h431111e0, 32'h43810828},
  {32'h43c99970, 32'h45028ef6, 32'h4486e95a},
  {32'h44155d09, 32'hc48f96bf, 32'hc2b64713},
  {32'hc423a8e8, 32'h442c0e84, 32'h4308fc35},
  {32'hc384f69a, 32'hc4009df8, 32'hc540a443},
  {32'hc51bc03c, 32'h43bbaba6, 32'h42478fa6},
  {32'hc4430381, 32'hc4414e11, 32'hc4c5bfa8},
  {32'h42bb83a8, 32'h44971609, 32'h43f30c23},
  {32'h441b2aa2, 32'hc527ec69, 32'hc420134c},
  {32'h44679f5e, 32'hc39d6aee, 32'h41858390},
  {32'hc2681530, 32'hc26c83a8, 32'hc5367d29},
  {32'h438515a6, 32'h43aa1eb0, 32'h44989608},
  {32'h43d72af8, 32'h421132f5, 32'hc44427cc},
  {32'hc512dc71, 32'h43847181, 32'h437857c4},
  {32'h45476ddf, 32'hc38ca362, 32'hc3b81005},
  {32'h4343ba3b, 32'h431269c6, 32'h42e4455d},
  {32'hc38f890e, 32'hc4e11c5c, 32'hc39de78c},
  {32'hc571575f, 32'h435c419e, 32'hc30e016e},
  {32'h45024db4, 32'h442cdc82, 32'hc349a67d},
  {32'hc4a26b13, 32'h44ea639b, 32'hc3540f53},
  {32'h45257832, 32'hc434d5d9, 32'hc2e5f900},
  {32'h44647400, 32'h4437bccf, 32'hc10c3a3e},
  {32'h4536abbf, 32'h41ac3f19, 32'hc3bca38a},
  {32'hc46fb634, 32'h44000e78, 32'h44023fb4},
  {32'h45142098, 32'hc3dfff70, 32'h431c79c5},
  {32'h4470ca49, 32'h42b8c78f, 32'h44f77196},
  {32'hc496b766, 32'hc36b4c5f, 32'hc261685d},
  {32'h4545a101, 32'h41f16487, 32'h4384b701},
  {32'hc3b2fcdc, 32'h44144bd2, 32'hc2f83c00},
  {32'h448e3184, 32'h44245269, 32'hc39b2631},
  {32'h40e3c100, 32'h45163cbb, 32'h4295d540},
  {32'h451539c1, 32'h43ea9dc9, 32'hc3dbc1ef},
  {32'hc397eade, 32'h45160137, 32'hc2cbba97},
  {32'h442d4ed0, 32'hc4734a94, 32'h43d081c8},
  {32'hc4cb5abc, 32'h42c20cb8, 32'h43726ec5},
  {32'h448019d0, 32'h443920f5, 32'hc4444839},
  {32'hc41ecfbf, 32'h41f02960, 32'hc51b6108},
  {32'hc3262e80, 32'hc315c9db, 32'hc391a076},
  {32'hc3a2deed, 32'h4380ec48, 32'h44b79487},
  {32'h44844752, 32'hc3586d91, 32'hc32a4d3f},
  {32'hc3fe50e7, 32'h4380f6e8, 32'h445a4c7f},
  {32'hc2eec174, 32'hc4758d56, 32'hc4ddc296},
  {32'hc3ef1d58, 32'hc3d05ff1, 32'h44e6fff0},
  {32'h4418544c, 32'hc3eee4df, 32'hc32b5004},
  {32'hc50cdc94, 32'h442aa1d3, 32'h444b6fb1},
  {32'h443d5882, 32'hc43953b0, 32'hc4abd940},
  {32'hc48738d7, 32'h439b9289, 32'hc2bd0035},
  {32'h44460992, 32'hc46c3a5a, 32'hc471c7ca},
  {32'h43157a2c, 32'h450af698, 32'h444ff233},
  {32'hc43b0195, 32'hc41f05fd, 32'hc3d63769},
  {32'hc41a4d2e, 32'h43755958, 32'h450de150},
  {32'h45367196, 32'hc40c52a8, 32'hc450b421},
  {32'h43a8f365, 32'hc3e282c2, 32'h422cd816},
  {32'hc56b0da5, 32'hc3cb3911, 32'h43db61b1},
  {32'h426751ab, 32'hc33cfd0e, 32'hc43c191f},
  {32'hc4616c54, 32'hc4d76aa4, 32'hc38336a8},
  {32'h453d5752, 32'h4352e797, 32'h440022b1},
  {32'hc50db773, 32'h441172e1, 32'h43f80f94},
  {32'h442f5d4e, 32'h4490ca20, 32'h4332bf0e},
  {32'hc44dc9a3, 32'hc4cceb68, 32'hc17321da},
  {32'h43fe5a4f, 32'h4486e0c8, 32'h43b1acca},
  {32'hc4f3a7da, 32'hc3ab7b44, 32'hc3106f42},
  {32'h4305f345, 32'h43a919fd, 32'hc325864e},
  {32'hc50b492a, 32'hc3227212, 32'h439d54a3},
  {32'h45496fd6, 32'h43e3ad26, 32'h4301bac7},
  {32'hc4b80e2a, 32'h4210b4cb, 32'hc39035d4},
  {32'hc3ad0a4d, 32'h43a570d3, 32'h4401e5fc},
  {32'hc5352a08, 32'hc3a86b8b, 32'hc28d47f3},
  {32'h44519b89, 32'h44f1316b, 32'h4402a14f},
  {32'hc537fd7d, 32'hc3abe6f3, 32'h43493165},
  {32'h4460398e, 32'hc44a7293, 32'h4469f43c},
  {32'hc533e4e3, 32'hc38259e9, 32'hc3d40dc6},
  {32'hc3f25764, 32'h41e48726, 32'h434e4a56},
  {32'hc3a5c1e9, 32'hc4aeb2ca, 32'hc4682838},
  {32'h423c6947, 32'hc3d8b043, 32'h45238b76},
  {32'h41be1ca8, 32'hc4c66943, 32'hc34e8202},
  {32'hc3285094, 32'h45046915, 32'h4438a249},
  {32'hc1f1ca3a, 32'hc549e8a2, 32'hc216a68a},
  {32'hc39960cb, 32'h44af248a, 32'hc32f3e4d},
  {32'h434a0ca6, 32'h450175a2, 32'h43a862a4},
  {32'hc514f8c1, 32'hc38e6283, 32'h437bb78b},
  {32'h44b4c957, 32'h43d4eabe, 32'h444467f7},
  {32'h42c2f49c, 32'hc4bdf847, 32'h440d0fca},
  {32'h40382700, 32'h4552bbc3, 32'hc321f826},
  {32'hc53b9687, 32'hc0e30865, 32'h435845ab},
  {32'hc4577bee, 32'h4390d11b, 32'hbfc4ad1b},
  {32'hc4b35bba, 32'hc3f0da1d, 32'h42f5d843},
  {32'h45230e50, 32'hc0b7266f, 32'h440710fa},
  {32'hc415dd99, 32'h4427b5b4, 32'hc35e3053},
  {32'h4422d83b, 32'h43863531, 32'h43897464},
  {32'hc43a902c, 32'hc2474876, 32'h43904651},
  {32'hc24f18b8, 32'h42380ce8, 32'hc3d35e99},
  {32'hc4462f75, 32'h43419a32, 32'h448a546b},
  {32'h451d9547, 32'h435aaa06, 32'h436bcc10},
  {32'h448bb01f, 32'hc24cb5dd, 32'h428ed260},
  {32'h4521b456, 32'hc429c9ac, 32'hc291da18},
  {32'hc48dace0, 32'h44189af0, 32'h44b37051},
  {32'hc3c5e65f, 32'h448a22d0, 32'hc216eab3},
  {32'hc55961c7, 32'hc40daf07, 32'hc22c200f},
  {32'h446ab33a, 32'h434e1967, 32'hc370595c},
  {32'hc3833daa, 32'hc342b525, 32'h450db964},
  {32'h4560e43c, 32'h441a0c09, 32'hc3d382fb},
  {32'h42340fd0, 32'hc3538946, 32'h4536ee81},
  {32'h443bbf0c, 32'h41019dda, 32'hc47dd1d2},
  {32'hc48e6174, 32'h44003a0f, 32'h44fc7e4d},
  {32'h42edf040, 32'h440e1de7, 32'hc481c850},
  {32'h44028798, 32'hc4076bfd, 32'hc4258d7b},
  {32'hc552b8b6, 32'h4370de34, 32'h43715fce},
  {32'h43f71d2c, 32'hc4b4e25b, 32'hc302d447},
  {32'hc4b8d460, 32'h44c05526, 32'hc2d61f9e},
  {32'h4471bf9c, 32'hc299b3ba, 32'h42e87082},
  {32'h445185e4, 32'h4412b983, 32'hc395c909},
  {32'h44fed722, 32'hc42a7a4c, 32'hc43924fb},
  {32'hc514cb47, 32'h4140be70, 32'hc313dcf6},
  {32'h4559da97, 32'hc22f994f, 32'h43ec9a96},
  {32'hc488eff3, 32'hc2b17b34, 32'h4425cef7},
  {32'h447ea502, 32'h42803a42, 32'h43b7027b},
  {32'hc2d852b2, 32'h43f8f770, 32'hc4cfcb7f},
  {32'h441ea2dc, 32'hc4dacd00, 32'h416a57eb},
  {32'hc5054db2, 32'h4399ccde, 32'hc4054047},
  {32'h4381a91e, 32'h42e5f9a6, 32'h443e751b},
  {32'hc52d1748, 32'h4111f90b, 32'h43489912},
  {32'h4414f789, 32'hc3da3483, 32'h442680e7},
  {32'hc3fefd13, 32'hc37074da, 32'h43c39389},
  {32'h432d81d0, 32'hc4c518b1, 32'h451000fe},
  {32'hc502962b, 32'h4430279d, 32'hc4667cd5},
  {32'h44535748, 32'hc473db57, 32'hc4019005},
  {32'h432a3040, 32'h4466836e, 32'hc4f12f75},
  {32'h437fddbb, 32'hc2e29d1c, 32'h452c0bdd},
  {32'h435ed428, 32'hc41ad451, 32'hc504c8d6},
  {32'h4530b2b8, 32'h43b4c388, 32'h437d2973},
  {32'hc4efc3a3, 32'hc3efa60c, 32'hc4e071d8},
  {32'hc422495a, 32'hc42605b8, 32'h43760db4},
  {32'hc32aa590, 32'hc322476a, 32'hc4a7ec99},
  {32'h43b7d333, 32'hc4b5ef3f, 32'h44f093f9},
  {32'hc4bbab24, 32'hc42a0588, 32'hc1980a48},
  {32'hc2389af8, 32'h44e07b47, 32'h4204bdbf},
  {32'h443e4f4d, 32'h429f1e19, 32'h44f59106},
  {32'hc345afec, 32'hc335ecca, 32'hc4ffcd6a},
  {32'hc4189273, 32'hc2cfb65c, 32'h447cc1f9},
  {32'hc540ceac, 32'h43eb4091, 32'hc2dc0a6d},
  {32'h4524e9d7, 32'h433b4713, 32'h443133ba},
  {32'h43b149c3, 32'hc32be8cb, 32'h450ce43c},
  {32'hc4ddc370, 32'hc297dd78, 32'hc4268ef0},
  {32'hc43b66f8, 32'hc2a378b0, 32'h4451de1a},
  {32'h44f23ae4, 32'hc3bc1ea9, 32'hc3a396e6},
  {32'hc3a691fb, 32'h4459d680, 32'hc4b483ba},
  {32'h44ebee35, 32'h4396690a, 32'hc20b7fe3},
  {32'h44ae9979, 32'h4417fd55, 32'h4190d558},
  {32'h44bb13f5, 32'hc4586060, 32'h42ec9e9f},
  {32'hc44362aa, 32'h4438282b, 32'hc364e69f},
  {32'h45156cc5, 32'hc375b68b, 32'hc1f1771b},
  {32'hc562486c, 32'hc20c8ed8, 32'hc3bb2608},
  {32'h42012f40, 32'h448468ef, 32'h4416311a},
  {32'h44e91cb6, 32'h4363acf6, 32'h436be26d},
  {32'h44619354, 32'hc44d49ea, 32'hc32cf8b6},
  {32'hc409ad7c, 32'h44a7c499, 32'hc3053fde},
  {32'h440a4b46, 32'hc3bf086c, 32'h43161098},
  {32'hc5624bcb, 32'h4254c15e, 32'hc3719ed2},
  {32'h45455b0b, 32'hc40a4ac6, 32'hc22147b7},
  {32'h43d74f34, 32'h43efc960, 32'h44177d69},
  {32'h44295711, 32'h449fbbfe, 32'hc42c6cf0},
  {32'h438d66f6, 32'h4472c002, 32'h4536c209},
  {32'hc4b695dd, 32'hc371de3d, 32'h431c3689},
  {32'h453b2752, 32'hc1a97f30, 32'h401f95ba},
  {32'hc490f52a, 32'h404faca0, 32'hc22bad48},
  {32'hc3e76fb5, 32'h43bb10f3, 32'hc453d55e},
  {32'hc515c061, 32'hc42537c0, 32'h43c7dee4},
  {32'h44b9cc89, 32'h440a1e12, 32'hc2d9a45d},
  {32'h42bcb73c, 32'h44658c56, 32'hc2a644f8},
  {32'hc4cf7988, 32'h4254b588, 32'h42d28d58},
  {32'hc39c2f9e, 32'h43d2e869, 32'hc4f97b6b},
  {32'h44cd986c, 32'h44004b51, 32'hc408c364},
  {32'hc347247c, 32'hc43cc2dd, 32'h44897fbd},
  {32'h43bc1b61, 32'h44d657ad, 32'hc3f63697},
  {32'hc38558e5, 32'hc40de694, 32'h44c049c4},
  {32'h450808c8, 32'h43bd9332, 32'hc2a98350},
  {32'h42eb1a16, 32'hc32bd5a0, 32'h440b9e78},
  {32'h447f5b12, 32'h4200d241, 32'hc3310d47},
  {32'hc5912248, 32'hc31ed3e2, 32'h4341ce07},
  {32'h448dee61, 32'h43bd72b6, 32'hc341f693},
  {32'hc3d3f628, 32'hc5060cc0, 32'h41a17cda},
  {32'h44a75e53, 32'h44bfb9e9, 32'hc242cf55},
  {32'h44c31880, 32'hc3a7dd80, 32'h435db186},
  {32'hc2dc8aea, 32'h4570b921, 32'hc38fad29},
  {32'hc52acd06, 32'hc441b7cc, 32'hc3f4928e},
  {32'h446d8b96, 32'hc31d43fc, 32'hc2f91082},
  {32'h444c34b4, 32'hc3b96682, 32'hc3cc34f3},
  {32'hc3c351d6, 32'hc5116cf9, 32'hc4408971},
  {32'h4477d554, 32'hc20c5eb9, 32'h4458fb16},
  {32'hc5124382, 32'h440a8d15, 32'hc32a8678},
  {32'hc36976ca, 32'h4451374e, 32'h42af2702},
  {32'hc28b92d4, 32'hc53668d3, 32'hc2d5b5be},
  {32'hc4c0e2f4, 32'h43c51d71, 32'h43ca7248},
  {32'hc53a60ce, 32'hc3a72f12, 32'hc4484f5a},
  {32'h450928fb, 32'h43fc5446, 32'h442c1db8},
  {32'h431e2ba6, 32'hc4c885d0, 32'hc32fa8f6},
  {32'h4385b69e, 32'h442cff55, 32'hc141410b},
  {32'h42f044b6, 32'hc4547723, 32'hc4884e4d},
  {32'h44c74e2e, 32'h438a9481, 32'h43827965},
  {32'hc4943d49, 32'hc33890a2, 32'hc42ac758},
  {32'h4495160f, 32'h44a4e8c8, 32'h4309007e},
  {32'hc42b8e5c, 32'hc1048cdd, 32'hc421e664},
  {32'h44ba9055, 32'h435e4b96, 32'h43e424f7},
  {32'h43eaec8e, 32'hc499957f, 32'hc520ebc8},
  {32'h4215a366, 32'h448a6c47, 32'h438edf95},
  {32'hc384f7e8, 32'hc530e303, 32'hc42f853b},
  {32'h445f6a3a, 32'h44939625, 32'h4418f223},
  {32'hc3970112, 32'hc4b80f89, 32'h428ae49f},
  {32'h4560ca3d, 32'h438b9e00, 32'h43d28045},
  {32'hc53ee5b3, 32'hc3044288, 32'h430ecc41},
  {32'h45673e87, 32'h43a93f00, 32'h43a1d134},
  {32'hc564b1b8, 32'hc2449259, 32'hc4425804},
  {32'h437fca7e, 32'hc3f73466, 32'h438c3225},
  {32'hc3912973, 32'h440f5f8c, 32'hc4f3a3fc},
  {32'hc2e69ca9, 32'h440a455f, 32'h4264438d},
  {32'h44160c00, 32'hc34f80a8, 32'hc37077c9},
  {32'h4277ddc0, 32'h43e3ae4c, 32'h453518d1},
  {32'h43f0aeb8, 32'hc0314f0e, 32'hc50d2e00},
  {32'h431eab78, 32'h43d9b3ef, 32'h4334f582},
  {32'h44d050fa, 32'hc47c9cbb, 32'hc49cc34a},
  {32'hc30b9fdf, 32'h442ce93d, 32'h4559bedd},
  {32'h448d49bb, 32'hc423dad5, 32'hc1ad69de},
  {32'h4346adc8, 32'hc1ff7b0f, 32'h44d7a0ba},
  {32'hc2ae8674, 32'h44480cc1, 32'hc4eae354},
  {32'h4409f312, 32'h444e77ae, 32'h43d83a79},
  {32'h43ab1d82, 32'hc43cb2c2, 32'hc46f440b},
  {32'hc4612a22, 32'h44016766, 32'h4485dfce},
  {32'h44a22f06, 32'hc32046c2, 32'hc39da310},
  {32'h438d637a, 32'h4508dba8, 32'h44975761},
  {32'h44d0512e, 32'h43f01fb0, 32'hc395d51b},
  {32'hc32cb38c, 32'h44399376, 32'h43c16c5b},
  {32'h4505e4a6, 32'hc43bce47, 32'h4280b44a},
  {32'hc4a9022c, 32'h4447622a, 32'h43fc15ff},
  {32'h446a234d, 32'hc230b29e, 32'hc3bc6f74},
  {32'hc514cdda, 32'h42b24a38, 32'h43765b46},
  {32'h44424b34, 32'hc4a3328c, 32'h4303be92},
  {32'hc46c52b0, 32'hc3cbe367, 32'h427a1805},
  {32'h45646895, 32'h439e9b3a, 32'h44277292},
  {32'hc589447d, 32'hc1145a6c, 32'h43491b3e},
  {32'hc38edea4, 32'hc3f9a7a2, 32'hc4173043},
  {32'hc4919288, 32'hc3260652, 32'hc35bb8ba},
  {32'hc4beb86b, 32'hc2019e1b, 32'hc520bb96},
  {32'h44883a0c, 32'h4314b82d, 32'h44eae35f},
  {32'h43ba93d2, 32'hc2e2aeb3, 32'h43be3ff6},
  {32'h451cfa15, 32'hc4692c4f, 32'h42b6209d},
  {32'hc466df88, 32'h440e64fc, 32'hc3273e22},
  {32'h43563be1, 32'hc1c2ffc0, 32'h423078db},
  {32'hc3a61a80, 32'h4553a2d4, 32'hc2d3b8a4},
  {32'h45101007, 32'hc3cd3251, 32'h436a0d46},
  {32'hc52c4d7b, 32'hc3d35db8, 32'h413c7b38},
  {32'h4522ca50, 32'h43180fbb, 32'h41a431e7},
  {32'hc4a2f938, 32'h44a8399e, 32'h4420a630},
  {32'hc49fa20e, 32'h441e8feb, 32'hc3ae258e},
  {32'h4390ba36, 32'hbf8e86d0, 32'h4501f0a2},
  {32'h43ba4de0, 32'hc4538309, 32'hc452f121},
  {32'h44024dcc, 32'h42b0df2a, 32'h44de78a9},
  {32'hc485611c, 32'h42b7f712, 32'hc551c3ef},
  {32'hc53ea41e, 32'hc3eb0748, 32'hc302505a},
  {32'hc3a9adb6, 32'h43a851f5, 32'hc49a92f8},
  {32'hc4c9c505, 32'h43a65128, 32'h44a2a4ee},
  {32'h45178bad, 32'hc2d89878, 32'hc40c9f68},
  {32'h4435558a, 32'h423beb1f, 32'h42fe43d2},
  {32'h43f87b68, 32'hc240c9f5, 32'hc52db499},
  {32'hc4d6de8f, 32'hc317e4fc, 32'h441f82d3},
  {32'h4337e562, 32'hc38ea0fc, 32'hc4a8c0ba},
  {32'h423093d0, 32'h44529172, 32'h4520e16e},
  {32'h4545556f, 32'hc3758897, 32'hc406a965},
  {32'h451bc131, 32'hc32adcb1, 32'hc4a905db},
  {32'hc3a8b96a, 32'hc3517198, 32'h45483d39},
  {32'h44cff586, 32'h42623012, 32'hc2c9b0fe},
  {32'hc51a6e4d, 32'hc41dd60a, 32'h4316667e},
  {32'h4403b564, 32'h448fced4, 32'h42bd4770},
  {32'h450844ef, 32'hc2aed66c, 32'hc37a548a},
  {32'h43bb08ac, 32'h456d1402, 32'h432fe34c},
  {32'hc474f9f8, 32'hc48e3d57, 32'h43ea49c7},
  {32'hc41f85ef, 32'h448954ed, 32'h43cb3093},
  {32'hc48caec2, 32'h43c2ec88, 32'hc49687db},
  {32'h42f790b0, 32'hc190f77f, 32'hc52a81b5},
  {32'h445a6182, 32'h43ba6f82, 32'h43b1d802},
  {32'h451d2248, 32'h43bc23b8, 32'h43b9408a},
  {32'hc5227618, 32'hc368e865, 32'hc3499218},
  {32'hc3e91555, 32'h429725e2, 32'h440cd1b9},
  {32'hc2fb6600, 32'hc4af1289, 32'hc3d80d13},
  {32'h44155c14, 32'h4444cb70, 32'h44b1b59c},
  {32'h4364d2f0, 32'hc490a01c, 32'hc458c0c1},
  {32'h44e3eec8, 32'h4408a768, 32'h4345a56b},
  {32'hc52cd2ac, 32'h42f841f4, 32'h423de678},
  {32'hc4baeec4, 32'hc29a2206, 32'hc1399eb8},
  {32'hc3f49ce0, 32'hc3b7ec68, 32'hc48da875},
  {32'hc35aa070, 32'h433c3b8a, 32'h451b0a58},
  {32'hc2834716, 32'hc3ffde33, 32'hc45bd29d},
  {32'h4521b2e3, 32'h432f4187, 32'h442ae6a0},
  {32'hc53a5f1f, 32'hc3e3a689, 32'hc397cb94},
  {32'hc43da2aa, 32'h441f0ca0, 32'hc28dd035},
  {32'h440a49c8, 32'h448b35a8, 32'h4320bbbb},
  {32'hc4b5c554, 32'hc413e1a2, 32'hc2e633d7},
  {32'h453dafbc, 32'h43404d0e, 32'h43dc7f8f},
  {32'h4492eb60, 32'hc4388d6d, 32'h4281b59e},
  {32'h44b744ed, 32'h441ed204, 32'hc46267d3},
  {32'hc212035e, 32'hc51bd7cd, 32'h432717e4},
  {32'h43ea8b28, 32'hc31ac999, 32'h427ae3e2},
  {32'hc4671b6a, 32'hc457462c, 32'hc42da5bd},
  {32'h440c79e0, 32'h43fcbd89, 32'h446ed97c},
  {32'hc527c2d7, 32'h432de769, 32'h42cc2daf},
  {32'h442add37, 32'hc3edc201, 32'h44b2293a},
  {32'hc33ceb58, 32'hc4eb6dda, 32'hc3964024},
  {32'hc3cbbf06, 32'h4408b6a2, 32'hc3a38d02},
  {32'hc3fcb05b, 32'hc4a71aec, 32'h43669112},
  {32'h44b3c978, 32'h42256886, 32'hc125796e},
  {32'hc44dd843, 32'hc32e57b9, 32'hc1b4e475},
  {32'hc0775580, 32'h43834ac5, 32'hc52b3873},
  {32'hc4a120e2, 32'hc3834533, 32'h43102cb8},
  {32'h44d66bc4, 32'hc32457f8, 32'hc3d16dd2},
  {32'hc54a78cc, 32'hc3c9c7b7, 32'h42f54bb2},
  {32'h44fe0b59, 32'h446fe2f8, 32'hc380237a},
  {32'hc4cb5949, 32'hc35674a4, 32'hc3685b85},
  {32'h43e6e442, 32'h450da3ec, 32'hc3191c2b},
  {32'hc4b6a1eb, 32'hc1fb8dfb, 32'h440a8386},
  {32'h42d69966, 32'h41b4fb26, 32'hc4425cc1},
  {32'hc53852c2, 32'hc340205f, 32'hc21561ac},
  {32'h43b8fd10, 32'h440c26d0, 32'hc4c755f6},
  {32'h44191323, 32'hc4f82952, 32'hc3ca6b50},
  {32'hc579dbd4, 32'h436ecf76, 32'h44141742},
  {32'h44e16bae, 32'hc32042f2, 32'h43a2c348},
  {32'hc42fcdf3, 32'h4457a081, 32'h441704a6},
  {32'h43583c08, 32'hc4ed263a, 32'h4312bec7},
  {32'h448bf9af, 32'h44a8abb7, 32'h4318fed6},
  {32'h43bf513c, 32'hc3e644df, 32'hc1f0b295},
  {32'hc54eaecf, 32'h43889f61, 32'hc3c9e0f6},
  {32'h44dc1728, 32'hc3d3163b, 32'hc3a31ddb},
  {32'h43fdd5f4, 32'h44584d94, 32'hc4b665e1},
  {32'h4456a8bd, 32'h43c58ec6, 32'hc4280a44},
  {32'hc34d3165, 32'hc32bd6a9, 32'hc4b91245},
  {32'h43be57e1, 32'h438cbbb0, 32'h44e4b007},
  {32'hc4af8478, 32'h44583194, 32'hc3998bcd},
  {32'hc4ae50ff, 32'hc37dcb7c, 32'h4364f2d5},
  {32'hc4c8c01a, 32'h434602bc, 32'hc42838d5},
  {32'h441ba986, 32'h430a4e54, 32'h44079b4a},
  {32'hc3a44b84, 32'hc39c841d, 32'h42801558},
  {32'h4409b6ee, 32'hc5423db1, 32'hc3e612b0},
  {32'hc3f02bb8, 32'h454d048f, 32'hc394f9f8},
  {32'hc306b098, 32'hc2b6eefd, 32'h4499480b},
  {32'hc43ca3d2, 32'h438ec8a5, 32'hc3a3dca4},
  {32'h44272a2c, 32'hc20c4e8a, 32'h44c04864},
  {32'hc471c41c, 32'h417e12fe, 32'h4345c56f},
  {32'h44df260c, 32'hc306a8fd, 32'h4450f567},
  {32'hc493089a, 32'hc36b355d, 32'hc2f3372b},
  {32'h44d6e15c, 32'hc3cdd306, 32'h4387ed31},
  {32'h42983e59, 32'h43b166af, 32'hc51b1c70},
  {32'hc4c489f5, 32'h43cc1415, 32'h449c073e},
  {32'h438f48dd, 32'hc36088ab, 32'h440bb6c7},
  {32'hc403b66a, 32'h42e80b5b, 32'h43587231},
  {32'hc3690055, 32'hc551200e, 32'h42697cc0},
  {32'hc39f2e71, 32'h44a1c649, 32'hc3fa87f7},
  {32'h4509ba2e, 32'h438f4c9c, 32'hc24100e7},
  {32'hc4997d2d, 32'h446435cb, 32'hc391883f},
  {32'h4491b6a2, 32'hc3386bdc, 32'h4480a307},
  {32'h44cf3f30, 32'hc43925f6, 32'h442d6433},
  {32'hc39fdd0a, 32'h44986eb6, 32'hc4b6b925},
  {32'hc388ddbe, 32'h4489c3f5, 32'h4486d5f9},
  {32'h444e42f7, 32'hc30884d8, 32'h4454a00a},
  {32'hc3f8a3e9, 32'hc30bef1e, 32'hc4bb28cf},
  {32'h43b74d48, 32'hc504b1c4, 32'hc347ead9},
  {32'hc29cd058, 32'h44815ae8, 32'hc157f11c},
  {32'hc3cf9359, 32'hc2d8ed07, 32'h42b4e06a},
  {32'hc3909050, 32'h4408cd7e, 32'hc50e3082},
  {32'h437294fa, 32'hc3fbd7aa, 32'h440541c0},
  {32'hc50ccf20, 32'hc3b69067, 32'hc438d5f7},
  {32'h44e2ff82, 32'hc3d437dd, 32'h4429cea7},
  {32'h44e6267d, 32'hc35cc2bd, 32'hc39fd020},
  {32'h4543efa0, 32'h44269590, 32'h420f417a},
  {32'hc5174943, 32'h42ce912c, 32'hc3250d74},
  {32'hc2887086, 32'hc4b2e2a7, 32'hc41edbd0},
  {32'hc350ba8c, 32'h456e83f2, 32'h430d7709},
  {32'hc308c1d8, 32'hc524d91d, 32'hc3fa76c6},
  {32'hc3a3b122, 32'hc49b8413, 32'hc2b8c0fd},
  {32'hc38fbf9f, 32'h4483f8d1, 32'hc4d25cc7},
  {32'h418b91f2, 32'hc38533c4, 32'h4465a12e},
  {32'h43356900, 32'hc495ae05, 32'h4437ef3b},
  {32'h4405fd03, 32'h4549b46f, 32'h43f9c5b3},
  {32'hc50c3023, 32'hbe00b5c0, 32'hc4053d53},
  {32'h444c7f7c, 32'h4428fa85, 32'hc49feaa3},
  {32'hc500c639, 32'hc4630351, 32'h43148031},
  {32'hc42474cb, 32'h44178312, 32'hc3fadae1},
  {32'hc43ac376, 32'hc3d49a6d, 32'h41cad42b},
  {32'hc52e727a, 32'h42f8e466, 32'h43a26c80},
  {32'h44827148, 32'hc35853ae, 32'hc4500265},
  {32'h439aa2d1, 32'h450e8d3e, 32'h42a0d7ff},
  {32'hc46400e1, 32'hc4dcdee3, 32'h433c0a82},
  {32'h44290597, 32'hc3623538, 32'h42ad6556},
  {32'hc23f4b55, 32'hc4015f40, 32'h42aec574},
  {32'h45223657, 32'h438ba335, 32'hc3be2ece},
  {32'hc4f87bea, 32'hc40757bc, 32'h43cbad48},
  {32'h4421fcc8, 32'hc1cf54de, 32'hc435aefe},
  {32'hc57fd6ca, 32'h434b04d3, 32'h4103c548},
  {32'h449dbe2f, 32'h43fbee03, 32'hc1f2f3f2},
  {32'hc4438100, 32'hc343cae9, 32'hc3e8a883},
  {32'h43f7f370, 32'hc34429b5, 32'hc3d1c6c5},
  {32'h4468ec25, 32'hc3a67e9c, 32'hc3a5440f},
  {32'h4403f5e0, 32'h44b00e99, 32'hc421dde3},
  {32'hc404f54e, 32'hc4dc0314, 32'hc3de6e86},
  {32'hc35d33a0, 32'h43db8cbf, 32'hc41aa5fc},
  {32'hc184e500, 32'hc4c62840, 32'h44977178},
  {32'hc49814f6, 32'h420e180c, 32'hc457ba0f},
  {32'h43a17342, 32'h4510b215, 32'h441c5e61},
  {32'hc30e1d42, 32'hc4d3aaa5, 32'hc360d5df},
  {32'h455e378c, 32'hc3548001, 32'hc171e4d5},
  {32'hc4015c68, 32'hc314280f, 32'hc518b1b5},
  {32'h44c0c260, 32'h44372887, 32'hc2aabe3d},
  {32'hc43cf816, 32'hc2f0597a, 32'hc4870be1},
  {32'h43a11662, 32'h4502ff09, 32'h446e051f},
  {32'hc43b47f9, 32'h44bd5a50, 32'h42978764},
  {32'h4380bc7d, 32'hc3d43cba, 32'h4380f9f2},
  {32'hc43daf8a, 32'h44ae05c5, 32'hc4fd3c53},
  {32'h447d2228, 32'h43a9dd59, 32'h4257eccf},
  {32'hc448a3c8, 32'hc432c230, 32'hc3b9a41f},
  {32'h447bad80, 32'h4461fec3, 32'h446eca3c},
  {32'h44d8396e, 32'hc3b198e5, 32'h42e88a0f},
  {32'h44b050d6, 32'h44274c33, 32'h441fceaa},
  {32'hc4e0bdc2, 32'h429cb256, 32'hc49955c4},
  {32'h44406eaf, 32'h43ae9445, 32'h435a32ba},
  {32'hc54aa362, 32'hc3b36fda, 32'hc29786de},
  {32'h445e3cc6, 32'h44bd7cc0, 32'h4449f064},
  {32'h4412e593, 32'hc464a62e, 32'hc3c51174},
  {32'h452e8c02, 32'h43bcef59, 32'h433b0ccc},
  {32'hc542cb27, 32'hc3391c79, 32'hc2e2fe61},
  {32'h4505b107, 32'h43db1ef1, 32'h44152b09},
  {32'hc57282d9, 32'hc35575db, 32'hc3be3b6f},
  {32'h4512b3ee, 32'hc36d9718, 32'hc2cb4ea8},
  {32'hc3b9f673, 32'h44bc8e7e, 32'hc50037cc},
  {32'hc43afd28, 32'h41bd679f, 32'h4316e2c8},
  {32'hc4749854, 32'hc37992ad, 32'hc30a4122},
  {32'hc0a64000, 32'h4389eee5, 32'h450f3e68},
  {32'h45318085, 32'h42c6480b, 32'h432d8bcb},
  {32'hc5195bc7, 32'h43cb113e, 32'h42e3d827},
  {32'h44171cc2, 32'hc4b80db8, 32'hc4a09402},
  {32'hc4020f09, 32'h43929faa, 32'h44c5a7f3},
  {32'h41881aff, 32'hc4a66641, 32'hc4a4aa1f},
  {32'hc420b46e, 32'hc42368f6, 32'h442b9832},
  {32'h444e38ee, 32'hc2aed71b, 32'hc2a51675},
  {32'hc4216536, 32'hc47fc502, 32'h449c638e},
  {32'h4480a3ae, 32'hc4094f9d, 32'hc4631fc1},
  {32'hc408e507, 32'h436e49ce, 32'h428135ca},
  {32'hc3cc5546, 32'hc4d0048b, 32'hc14893ca},
  {32'hc4116a80, 32'h4489242d, 32'h449ef2a3},
  {32'hc40d705c, 32'hc48828fa, 32'hc56e6bb6},
  {32'hc4f00f32, 32'hc3480428, 32'h43e8fdf9},
  {32'h44919082, 32'hc4a9ac25, 32'hc3b8fa2a},
  {32'hc486ac0e, 32'h4485b052, 32'hc2f7ad90},
  {32'h44cf6a22, 32'hc3996d3a, 32'hc335d8df},
  {32'hc3634f40, 32'h438abc46, 32'h4367c6aa},
  {32'hc233bcc7, 32'hc56c3383, 32'hc3c053e9},
  {32'h4476809b, 32'h4440d46c, 32'h4087b488},
  {32'h4418f274, 32'h44967121, 32'h42c3260e},
  {32'hc52cea91, 32'h44607517, 32'h4411a4a5},
  {32'h453a2e36, 32'hc357fdc4, 32'hc3d1272b},
  {32'hc3cea005, 32'hc3ec4b7b, 32'hc37b9f27},
  {32'hc420b505, 32'hc3279201, 32'hc404a901},
  {32'h44d8f860, 32'h43aa1250, 32'h43e5b043},
  {32'h43298b4c, 32'hc32330cf, 32'h440edb1c},
  {32'h450131c5, 32'hc327cfd1, 32'hc3053fcb},
  {32'hc4c6d7e4, 32'h44ad7960, 32'h43cc0c29},
  {32'h45558a92, 32'h4420f389, 32'hc3cfb19a},
  {32'hc3e9aff6, 32'h45192bda, 32'h3f1b9b95},
  {32'h434e73a5, 32'hc566895e, 32'hc3888013},
  {32'h446042ce, 32'h438a2218, 32'h42bf49d0},
  {32'h431c0580, 32'h436436a4, 32'h43732c1e},
  {32'hc3bceacd, 32'h442dffca, 32'h446c8090},
  {32'h41527400, 32'h4392db7c, 32'hc2f6e2ef},
  {32'h44018b5b, 32'h4415922b, 32'h44a0046d},
  {32'hc212b184, 32'hc44516ed, 32'hc319ec91},
  {32'h43592cce, 32'h441cbdb2, 32'h44280259},
  {32'h4482ec47, 32'hc4825d72, 32'hc43443ea},
  {32'hc4a1f758, 32'hc318347d, 32'h4430752d},
  {32'h441a659d, 32'h436d4d59, 32'hc435658f},
  {32'hc530cfe8, 32'hc4634eec, 32'h42f25c4e},
  {32'h456b70f5, 32'h442e9c04, 32'hc1b22508},
  {32'h43857afc, 32'h43f0ffb2, 32'h44d5a98e},
  {32'h440d54b9, 32'hc505b0bc, 32'hc1f1a571},
  {32'hc4216ad3, 32'h44b157e2, 32'h43746516},
  {32'h4420f4ee, 32'h42a2d00c, 32'hc4a4d812},
  {32'hc4a2a688, 32'h4410f305, 32'h449b1f09},
  {32'h4411472c, 32'hc4a63cb3, 32'hc42e2020},
  {32'h43bd2ed7, 32'hc36d5d1f, 32'hc49a262d},
  {32'hc553156e, 32'hc306e8d8, 32'hc27e36c1},
  {32'h4542af86, 32'h42acf647, 32'h43dee982},
  {32'hc46b9531, 32'hc48868d3, 32'hc2cfbe54},
  {32'h4459d4e2, 32'h449b2732, 32'hc2d5496f},
  {32'hc31fd2f8, 32'hc4a68349, 32'hc2cb485a},
  {32'h441d9864, 32'h450d33ca, 32'hc2c94340},
  {32'hc540214c, 32'hc431674e, 32'h412e2e60},
  {32'hc471ac9f, 32'h4431ee3a, 32'hc32f3c14},
  {32'hc1bad580, 32'h43be340b, 32'hc466304a},
  {32'h4415ee4a, 32'h439b5dc9, 32'hc4ab523f},
  {32'hc31c8d50, 32'hc39a4b38, 32'h444fe910},
  {32'h42e71d10, 32'hc2e9bbee, 32'h4542122a},
  {32'hc4140037, 32'hc25a6a26, 32'hc55e7265},
  {32'h42d21544, 32'h44880461, 32'h43f6d74d},
  {32'hc2ccd94e, 32'hc4ecc75a, 32'hc271e5df},
  {32'h42823475, 32'h44025130, 32'h4529975c},
  {32'h43fd1730, 32'hc41148cd, 32'hc4072c69},
  {32'hc379da93, 32'hc41afe08, 32'h4472d5a6},
  {32'hc538aa90, 32'h428616ab, 32'hc38525f0},
  {32'h43fc9e0b, 32'hc33ecbf9, 32'hc3e72f4b},
  {32'hc0c9363f, 32'hc3ec5da9, 32'hc46a4006},
  {32'hc3874c18, 32'h44f7346f, 32'h442da418},
  {32'hc407a53f, 32'h428e9214, 32'hc390e27e},
  {32'h4422081e, 32'h440cd753, 32'h43a6c4ed},
  {32'hc343adaa, 32'hc514d5d9, 32'hc4036c80},
  {32'hc41a6a6c, 32'hc0c83b2a, 32'h44019e7e},
  {32'hc28bf744, 32'hc21e470e, 32'hc3e1c533},
  {32'hc29c58ba, 32'hc4fca412, 32'hc387d59b},
  {32'h443186e6, 32'h44a2e98c, 32'hc387809d},
  {32'h40989250, 32'hc3e012c9, 32'hc2f7b7ca},
  {32'h44e39e47, 32'h446f9c31, 32'hc2447a04},
  {32'hc48d488b, 32'hc39c9808, 32'hc405e429},
  {32'h44efbc21, 32'h4397e0c6, 32'hc2ca6c9d},
  {32'hc4e896fe, 32'h43d765de, 32'hc33175b9},
  {32'h45123652, 32'hc3b15b02, 32'h44613a8e},
  {32'h44515379, 32'hc3c2d4b5, 32'hc34a1132},
  {32'h45094492, 32'h433372a2, 32'hc2da2ee3},
  {32'hc38d45a6, 32'hc4836b8d, 32'hc399f7fe},
  {32'hc494b722, 32'h44407e8f, 32'hc290d188},
  {32'hc49ff262, 32'hc3be7405, 32'h445e8d23},
  {32'h43930eaa, 32'h4532215c, 32'hc21c8f5d},
  {32'h440a963b, 32'h43920d13, 32'h43aa0aa9},
  {32'h443bcb46, 32'h440664b9, 32'h42e7e746},
  {32'hc4d287a1, 32'h423c93ce, 32'h43dfb496},
  {32'h43c91f77, 32'h438df1b1, 32'h43ae711c},
  {32'hc506fc1b, 32'hc3d3dc1e, 32'h431eba99},
  {32'h443d46d0, 32'h44cb55e7, 32'hc4804a47},
  {32'h4453e60f, 32'hc27ebc39, 32'h42927c01},
  {32'h440976ee, 32'h443828cd, 32'hc4b91b4e},
  {32'hc2dd9bd0, 32'hc443160d, 32'h445d2bee},
  {32'h44ad0499, 32'h42ee985f, 32'h42815096},
  {32'hc4f4ba4b, 32'hc3a1d4c3, 32'h4493705e},
  {32'h429e1bf2, 32'hc4125c9e, 32'hc579a656},
  {32'h440de411, 32'hc50772de, 32'hc3887be0},
  {32'hc4141e68, 32'h44d47f6d, 32'h432260f7},
  {32'h449fa1db, 32'hc3f04b57, 32'h43059419},
  {32'hc47a588a, 32'h4501f4dc, 32'hc275cdeb},
  {32'h44ce275a, 32'hc46b180b, 32'hc24fb451},
  {32'hc4b6a1d0, 32'h43eaf43e, 32'h43a6ba51},
  {32'hc3d1d226, 32'hc3cb8b38, 32'hc38eae89},
  {32'hc512e44c, 32'hc3fb7168, 32'hc1fe9956},
  {32'hc4399c2e, 32'hc3537b14, 32'hc231c634},
  {32'hc28be6e8, 32'h449bd466, 32'hc507761f},
  {32'h4443bad8, 32'hc3a75014, 32'h43ad0884},
  {32'hc36e3a10, 32'h444268c1, 32'hc396e6b2},
  {32'h4379c5b0, 32'h414fee80, 32'h452e38c3},
  {32'hc1ec5bd8, 32'h44135a46, 32'hc3afe392},
  {32'h44f4de73, 32'h431bc582, 32'h43a3de5a},
  {32'h42057810, 32'h44351775, 32'hc4074142},
  {32'h4353e39c, 32'h4332e09e, 32'h449cb782},
  {32'hc1e29546, 32'h43b1495c, 32'hc42b00c0},
  {32'h45299255, 32'hc3992b5a, 32'hc437bc53},
  {32'hc3c88276, 32'h44c19fea, 32'hc504fe85},
  {32'hc36807bc, 32'hc33c18e3, 32'hc25d0885},
  {32'h427f1611, 32'h43a2b915, 32'hc42f5655},
  {32'h432265c8, 32'hc506b5ce, 32'hc3aaf8ed},
  {32'h4354e0e4, 32'h44b0f738, 32'hc3c4b9e7},
  {32'h44b181ec, 32'h41f10073, 32'h44573dc2},
  {32'hc3d9f958, 32'hc32de80d, 32'hc57d3aa2},
  {32'hc4a9dbdf, 32'h430f20fe, 32'h43401bfd},
  {32'h43087027, 32'h448fa552, 32'hc4ad93ee},
  {32'hc36ad40b, 32'hc4243ae6, 32'h451b94e7},
  {32'h43b3e315, 32'h443eae7c, 32'hc3d30bea},
  {32'h448ec556, 32'h4401ae51, 32'hc401f23f},
  {32'h45122af0, 32'hc359cf5f, 32'h44813ae1},
  {32'hc32e1a68, 32'h41ac515c, 32'hc5113492},
  {32'hc4bb65c7, 32'hc3ebf76f, 32'hc345e0c8},
  {32'hc501afa1, 32'h43953b95, 32'hc38699a5},
  {32'h452713a3, 32'hc4159b33, 32'h445784aa},
  {32'h43dec8a4, 32'h43ed5e3d, 32'h44b52399},
  {32'hc481362e, 32'h4412e0de, 32'hc496b855},
  {32'hc3758ba3, 32'h4486c889, 32'h449e1df1},
  {32'h443d159f, 32'hc2689ae0, 32'h43ccefbf},
  {32'hc3c026ee, 32'h42aa0166, 32'hc50635b0},
  {32'hc10e3e00, 32'hc44d967d, 32'h442c1807},
  {32'hc443b0ca, 32'hc3b2dff3, 32'hc4215b88},
  {32'h4464aeda, 32'hc46f0528, 32'h430bbb85},
  {32'hc3b71705, 32'hc37b2992, 32'hc50dac05},
  {32'h4519ba77, 32'h43a6ced8, 32'h42428bda},
  {32'hc4e3a3e8, 32'h44149892, 32'hc39ade85},
  {32'h4502e16b, 32'hc3f82218, 32'h4399daf7},
  {32'h440119fb, 32'h44275dc7, 32'h4253a1ff},
  {32'h440f143c, 32'hc50dbd4b, 32'h430c49a3},
  {32'h431af2f7, 32'h455f937a, 32'hc1e5e947},
  {32'hc3d7230c, 32'h4381d401, 32'h4213bcdf},
  {32'hc4efc957, 32'h44c12907, 32'hc195e5d0},
  {32'h44c214e0, 32'hc4a26079, 32'hc35e33c5},
  {32'h43d13354, 32'h44299738, 32'h44270b4b},
  {32'hc2f84b22, 32'hc486bbfd, 32'hc46b84e7},
  {32'hc39eb1ce, 32'hc4f8a5ef, 32'h45066660},
  {32'hc544a992, 32'h435e73dd, 32'h416d487c},
  {32'h44e3903a, 32'hc38e232f, 32'hc45cb632},
  {32'hc46fd830, 32'hc42ec846, 32'h41915e89},
  {32'h45264e74, 32'h440728ab, 32'hc409bba8},
  {32'hc47dfff0, 32'hc4acfb62, 32'h43c0eef6},
  {32'hc365740f, 32'h44b51271, 32'h42001571},
  {32'h431a26e9, 32'hc38e58ab, 32'hc4f1e2ec},
  {32'hc5111ee1, 32'hc2b2e8a9, 32'h44aaffcc},
  {32'h43678c62, 32'hc4c7f5ed, 32'hc503c210},
  {32'h442e44ba, 32'h448326fb, 32'hc3ffde8e},
  {32'hc4e6fbf1, 32'hc347a01c, 32'h44139e20},
  {32'hc4958c5d, 32'h4349bced, 32'hc37f7243},
  {32'hc40bfeaf, 32'hc29059a2, 32'h451fadec},
  {32'h4483a6ef, 32'h443ad774, 32'hc3c5d0bc},
  {32'h42bff6c8, 32'hc3c4ad9e, 32'h43f5cda6},
  {32'h44d8b0b4, 32'h43f29a36, 32'hc2828f98},
  {32'hc55087e0, 32'hc28db5f7, 32'hc2b35f93},
  {32'hc4a3647b, 32'h41ca85a9, 32'hc281b818},
  {32'hc4c9e929, 32'hc4b454b9, 32'h42b865c4},
  {32'h43a7aff4, 32'h44bfe6c2, 32'hc27c79bb},
  {32'hc2a5606c, 32'hc5070c86, 32'h427e8601},
  {32'h44da1240, 32'h44a70c02, 32'hc41df846},
  {32'hc46e6ee4, 32'hc4de057f, 32'h43a1762e},
  {32'h45466a65, 32'hc44033c9, 32'h424123f4},
  {32'h43b2efa9, 32'hc4cb6750, 32'h439f1573},
  {32'hc3b66849, 32'h43e1bc05, 32'hc4f0f378},
  {32'h44551ef1, 32'hc2ccf4da, 32'h443fafa4},
  {32'h43f57ef3, 32'hc333e449, 32'hc3521480},
  {32'h4368b9e8, 32'h43bbf41e, 32'h453f63b5},
  {32'h4243e346, 32'hc4ebf117, 32'hc37a280e},
  {32'h42959771, 32'h44a40712, 32'h44804e34},
  {32'hc3dcf990, 32'hc3fb6fd0, 32'hc4c417f1},
  {32'h44fc25de, 32'h442e7921, 32'h440031a7},
  {32'h44a0ac7f, 32'h440ac5b8, 32'hc37dcd25},
  {32'hc312a2fc, 32'h451277d5, 32'h43a2a417},
  {32'hc407a199, 32'h443ff5c1, 32'hc4c31a3e},
  {32'h438f51c4, 32'hc132fc26, 32'h44c18590},
  {32'hc28baf48, 32'hc462a926, 32'hc4567be0},
  {32'h441d5ea3, 32'h43913abb, 32'h450f7198},
  {32'h44e2b840, 32'hc40d60ca, 32'hc1a74b92},
  {32'h44b9c465, 32'h43a4b5d1, 32'h44bdad6d},
  {32'h43f1782a, 32'hc4af6398, 32'hc51df7c1},
  {32'h453dc3be, 32'h42f36b85, 32'h43bcda21},
  {32'hc4d1228e, 32'hc46f50aa, 32'hc38d809e},
  {32'h44f9c7f8, 32'h44a2ad9e, 32'h441a7855},
  {32'h445a4950, 32'hc4e127f9, 32'h432f7a6a},
  {32'h440934f6, 32'h44ddb1d2, 32'hc3a0ea15},
  {32'hc39601e0, 32'hc58461b4, 32'h434f49c1},
  {32'hc41a33ca, 32'hc1c4cdfc, 32'h42831180},
  {32'hc5730741, 32'h410ef44a, 32'h43cf285d},
  {32'h4534d455, 32'hc254b812, 32'h444f8140},
  {32'h44f4a5e8, 32'hc44cb038, 32'hc4804233},
  {32'hc4c27569, 32'hc48c0849, 32'h44818a8a},
  {32'hc478b04d, 32'h43ca5658, 32'hc32741b5},
  {32'h438ad5ab, 32'h4516521f, 32'h442757b3},
  {32'h44588d00, 32'hc4a0b157, 32'hc46531a7},
  {32'h4398d0e6, 32'h42157657, 32'hc0865841},
  {32'h44388bf9, 32'hc3c52634, 32'hc4dc6613},
  {32'h4404519d, 32'h44203d94, 32'h44fb1bdb},
  {32'h4535011e, 32'h4353a338, 32'hc2bf2d65},
  {32'h430b725f, 32'h450ba636, 32'h438f6208},
  {32'hc32b7411, 32'hc3b947b2, 32'hc4a076d6},
  {32'hc3ad2ac6, 32'hc3eb68cb, 32'h44c33cbf},
  {32'h4236f0c0, 32'hc4be38c6, 32'hc4900a48},
  {32'hc4a26117, 32'h44ada7af, 32'h430213c2},
  {32'h4432d30f, 32'h42c2cd7d, 32'hc45818fd},
  {32'hc29b2888, 32'h44d71430, 32'h45098fa2},
  {32'h4524cf32, 32'h43d084bf, 32'hc396936a},
  {32'hc5295224, 32'h43817e77, 32'hc3086252},
  {32'h43a53213, 32'hc5719985, 32'hc1528ab1},
  {32'hc3faebaa, 32'h4474990b, 32'h43073215},
  {32'h42f28ff0, 32'hbfa439d0, 32'hc3f43d78},
  {32'hc3aa8676, 32'h455deb23, 32'hc333d44e},
  {32'h43ea79ea, 32'hc52aca50, 32'h428e6715},
  {32'hc4b3faa1, 32'hc1393512, 32'h44178358},
  {32'h44232950, 32'h44847693, 32'h4392c858},
  {32'hc581e534, 32'hc1bc38da, 32'h438ded35},
  {32'h44a7e05c, 32'hc29cf0eb, 32'hc3835a7a},
  {32'h45313cc4, 32'hc3293697, 32'hc3c9788a},
  {32'hc48cbf5c, 32'hc358ba9e, 32'hc3f9dc6d},
  {32'h443e36e4, 32'h43d06799, 32'h443e8b3e},
  {32'h44419b58, 32'h44b43158, 32'h41819ed4},
  {32'h43ce5215, 32'hc539a1e4, 32'hc3ce04ed},
  {32'hc4200254, 32'h44eef9ce, 32'h43c93b2f},
  {32'h435765fe, 32'hc3d8300c, 32'h4420db4a},
  {32'hc56a4806, 32'h43206668, 32'h42ae1cb4},
  {32'hc31cd67e, 32'hc42c5cc5, 32'h4402a0b5},
  {32'h44a05cea, 32'hc3a298c0, 32'h44191392},
  {32'h44082d39, 32'hc3b83f18, 32'hc2d2048e},
  {32'hc39a5dba, 32'h42f269b0, 32'hc489bd74},
  {32'hc33003cd, 32'hc3c802e0, 32'hc30e3d2c},
  {32'hc41e64f1, 32'h451965f5, 32'h44378130},
  {32'h438f5148, 32'hc51d7442, 32'hc2ead37d},
  {32'h4378cf92, 32'hc2ea44c4, 32'h450e2633},
  {32'h452dbbd8, 32'hc2f426d9, 32'hc42dfc11},
  {32'h42bedf33, 32'h41564028, 32'h4503c451},
  {32'h44b006ff, 32'hc4129893, 32'hc403164f},
  {32'hc42f712a, 32'hc45b803c, 32'h44558712},
  {32'h44638d96, 32'h444b01f4, 32'hc4d6a72a},
  {32'hc39cb926, 32'h44fce854, 32'hc1494408},
  {32'hc3aee59f, 32'hc368d15c, 32'hc4f5bbc2},
  {32'hc424ca81, 32'h44701235, 32'h43bb9af5},
  {32'hc4b28f92, 32'hc3d99f86, 32'hc4010d6b},
  {32'hc3f51710, 32'h4445b385, 32'h445bfa7f},
  {32'h440afdae, 32'hc3cf3000, 32'hc52da125},
  {32'h44023a6e, 32'h42b232b7, 32'h42d8537c},
  {32'hc3e25c90, 32'h43b9cbe5, 32'h442706df},
  {32'h4481d11b, 32'h43f27eaa, 32'hc3264cc4},
  {32'hc4972ca8, 32'hc4a7e516, 32'hc3d3f574},
  {32'h452045ea, 32'h432219a4, 32'h43d94746},
  {32'h449f7ed7, 32'hc27848cf, 32'h3fc9da60},
  {32'h43f44c22, 32'h45006b49, 32'h4405000d},
  {32'hc2e5c720, 32'hc54af19a, 32'hc385f354},
  {32'hc4560f2a, 32'hc2b534cd, 32'h428dec37},
  {32'hc437d18a, 32'hc3b0e5a1, 32'h4464cb79},
  {32'h43ba2ba8, 32'h438d45e6, 32'hc4750f02},
  {32'hc487652e, 32'hc3c06441, 32'hc3e6233c},
  {32'h44af1b17, 32'h447f7c70, 32'hc03d5fe0},
  {32'hc461da89, 32'hc4a94609, 32'hc416dd9d},
  {32'hc405e233, 32'h3d80df80, 32'h44de5a23},
  {32'hc404b40f, 32'hc3441ca0, 32'hc50f876c},
  {32'h438e3940, 32'h433bfbdb, 32'h449b0a34},
  {32'h42d370fd, 32'hc419771a, 32'hc37fb736},
  {32'h450ec090, 32'hc43a3978, 32'h42d6f76f},
  {32'hc3b735e6, 32'hc335b6ae, 32'hc4b511ef},
  {32'h4532a6b8, 32'h434f87f8, 32'hc3df9081},
  {32'hc53cc9b9, 32'hc3f76a65, 32'h438a7111},
  {32'h429a0627, 32'h449a94be, 32'h4444a8d8},
  {32'h4250e8d4, 32'h431c99a7, 32'hc4306cfa},
  {32'h44d19a80, 32'h448c7c76, 32'h43f392e8},
  {32'h437ff1aa, 32'hc4c225fa, 32'hc4be2e64},
  {32'hc3139ff8, 32'h433f4252, 32'h43c65ad7},
  {32'h43a19a3a, 32'h44c9c96a, 32'hc40caf2a},
  {32'hc53611f8, 32'h42de29c8, 32'hc3a877a5},
  {32'h4469f686, 32'h44b7bced, 32'hc19c4b92},
  {32'hc335961e, 32'hc4de159e, 32'h4396ec2a},
  {32'h4493444c, 32'h444a4338, 32'h42874cf3},
  {32'hc4f730ae, 32'hc44c403b, 32'hc194c5c9},
  {32'hc4cc4504, 32'h42de9fd4, 32'hc3aa7da1},
  {32'hc4962820, 32'h442828b6, 32'hc403b429},
  {32'h44396a3f, 32'h434eb57d, 32'h43da4c36},
  {32'h447b4c83, 32'hc229f4fe, 32'h430007c1},
  {32'h432bb674, 32'h44a5411c, 32'hc230b6ef},
  {32'hc3d5b31b, 32'hc2dc7300, 32'h440e1bda},
  {32'h44608a19, 32'h4451abd0, 32'hc49436ca},
  {32'hc45510aa, 32'hc4c00aa4, 32'h435a4637},
  {32'h43c70f94, 32'h4461e9e3, 32'hc43ab6b6},
  {32'h43db58f2, 32'hc0aec6db, 32'h42d1e2d9},
  {32'h43fdbf3a, 32'hc39a4b6b, 32'hc38ca2c7},
  {32'hc481fbc6, 32'h42ce6eae, 32'h430e558e},
  {32'h440dc124, 32'h43fa9cbe, 32'hc4aab5f6},
  {32'hc5358eb9, 32'hc1bd17ad, 32'h43c02dc8},
  {32'h4550e035, 32'h4369090d, 32'hc414ce2f},
  {32'hc3eb931d, 32'hc4b431dc, 32'h435b016c},
  {32'h43b76bcc, 32'h4517cc1d, 32'hc2fc57a1},
  {32'h4396b943, 32'hc3b49c08, 32'h4502d2b0},
  {32'h41d1029c, 32'h4117792f, 32'hc3b45fc8},
  {32'hc48c3133, 32'hc36a31f9, 32'h446aae9e},
  {32'h4517b4cd, 32'hc0bc1528, 32'hc3cc08ea},
  {32'h440fc898, 32'hc4cb6a91, 32'hc336dcab},
  {32'hc53ed3fe, 32'h4392cd0d, 32'h42f318c1},
  {32'hc496341f, 32'h43ccda0e, 32'h4357ebc9},
  {32'h43a6aa91, 32'h456d9d69, 32'h41ffb375},
  {32'h44e96718, 32'hc31ef33e, 32'h4403a66b},
  {32'hc51e0c60, 32'hc18ddcae, 32'hc38cd148},
  {32'h44a6833b, 32'h440762c8, 32'hc402c2f0},
  {32'hc58acd9d, 32'h43c89db7, 32'hc421d5bb},
  {32'h4522cb95, 32'hc1baab41, 32'h43b171fa},
  {32'hc292c56c, 32'h4379dd4c, 32'hc2fb7b04},
  {32'hc17d8d80, 32'hc48631b7, 32'h446602f1},
  {32'h44e1cd32, 32'hc2940111, 32'h435c0b52},
  {32'h43967334, 32'hc50eb37e, 32'h42f997de},
  {32'hc403b7e9, 32'hc3f73152, 32'hc48955fb},
  {32'hc4961ba6, 32'hc2a6a330, 32'h43add875},
  {32'hc415afb2, 32'hc3c29bb5, 32'hc519e83e},
  {32'h44c47500, 32'hc1d56e9a, 32'h445dd45e},
  {32'h449f9cd3, 32'h43a429e9, 32'hc47393e7},
  {32'h4245e400, 32'hc4e93e58, 32'h43e14c7f},
  {32'hc4a023c2, 32'h44ddb74c, 32'hc3c8ee40},
  {32'h45242ea4, 32'h418aa9a1, 32'hc338aba3},
  {32'hc428da03, 32'h451cd22e, 32'hc3715787},
  {32'h451f740b, 32'hc41f500b, 32'hc189ce32},
  {32'hc47e819b, 32'hc26b7a5e, 32'hc3027684},
  {32'h444d14c4, 32'h43cf2375, 32'h4510a517},
  {32'hc5344bcc, 32'h43b8b0a2, 32'hc44e4360},
  {32'h42b1ac3e, 32'h43cde022, 32'h446f7bd2},
  {32'h438d511c, 32'h441bfb95, 32'hc556f3e0},
  {32'h445e092a, 32'h43802f5e, 32'h44282365},
  {32'h42b7d70c, 32'h44887b63, 32'hc4c894b5},
  {32'h43ec8dba, 32'h445e6fd4, 32'hc40745c9},
  {32'h4517e308, 32'hc4294149, 32'hc363f3b5},
  {32'hc4699693, 32'h448282b7, 32'hc4264871},
  {32'hc395c424, 32'hc3e278d5, 32'h409b0980},
  {32'hc50fc7a2, 32'hc1e555fd, 32'hc43206f9},
  {32'h442251e4, 32'hc503cf8b, 32'hc3af4bdf},
  {32'h44b0dc01, 32'h4309bd23, 32'h448fc420},
  {32'hc4d74b99, 32'h43871d5a, 32'hc3790f16},
  {32'h451a4297, 32'hc3c1a8e6, 32'hc38cb031},
  {32'hc455e1fc, 32'hc3c8e24f, 32'h4331c941},
  {32'hc3f4fce5, 32'h44f5302f, 32'h42cf4c5d},
  {32'h44851815, 32'hc4b2e021, 32'hc2ed3a4f},
  {32'hc453a66c, 32'hc3e10b6e, 32'hc4646a14},
  {32'h4406e52c, 32'hc4fa6e1d, 32'h3f4c9380},
  {32'hc448ea9f, 32'h43fdb790, 32'hc41c25fd},
  {32'h438575a2, 32'hc28d4a67, 32'h4470a538},
  {32'hc56b2928, 32'hc3f3f3fb, 32'h43ac6d4e},
  {32'hc315ac20, 32'hc3826a4d, 32'h437b5873},
  {32'h44890145, 32'h449bc1a7, 32'hc3b72fd5},
  {32'h44132060, 32'hc5246884, 32'hc3c49b02},
  {32'hc3d786c4, 32'h42bbb4b7, 32'h43b57dcc},
  {32'h44cbb89b, 32'h43cbfea4, 32'h43492378},
  {32'hc4f562d1, 32'h4481620f, 32'hc403b9c9},
  {32'h440f3f39, 32'hc53c586f, 32'hc10c7620},
  {32'h441fd86a, 32'h43aa271e, 32'h41db9131},
  {32'h4420b605, 32'h4345fc36, 32'hc3954690},
  {32'hc4acfe84, 32'hc3c23ab9, 32'h43cb7a48},
  {32'hc48e3625, 32'hc49ade6f, 32'hc308fc80},
  {32'hc360753c, 32'h42ec82da, 32'hc4eea3b6},
  {32'h4433453f, 32'hc487c4fd, 32'hc2642ead},
  {32'h4469e869, 32'h44961621, 32'hc406f425},
  {32'h43ca49b0, 32'hc4363634, 32'h44dc74d9},
  {32'hc428cd5a, 32'h4493a3fa, 32'hc2d4d8b0},
  {32'h44435dc1, 32'h440fbba5, 32'h435d5fc9},
  {32'hc5250aa2, 32'h435d5632, 32'h44084113},
  {32'hc2c3e984, 32'hc2ce113d, 32'hc53f2c2b},
  {32'h43d0aa1e, 32'h43ac9996, 32'hc4a6f927},
  {32'hc338a450, 32'hc39260d5, 32'h44fc8a1a},
  {32'hc49e0b4f, 32'h4351b7cb, 32'hc3880df2},
  {32'hc4318c0e, 32'hc4f36e16, 32'h42fbaffd},
  {32'h439bdf32, 32'h43b23a1c, 32'hc43c4285},
  {32'hc2b73480, 32'hc19076b0, 32'h429e4bdc},
  {32'h44cf09ca, 32'hc32fc96b, 32'h4250889c},
  {32'hc4c86fb6, 32'hc382cecc, 32'hc40e6291},
  {32'h4520d71a, 32'hc2aba113, 32'h42fd52cf},
  {32'hc4f378af, 32'hc487774f, 32'h435b5c66},
  {32'h454cda7f, 32'h4378b912, 32'h43496767},
  {32'h44a977c2, 32'hc39187a0, 32'h42ba9178},
  {32'h4377b080, 32'h453da7cc, 32'h43e724a6},
  {32'hc4b06ca0, 32'hc484ff74, 32'h43542b91},
  {32'h4205232f, 32'hc33cb230, 32'hc4043c2d},
  {32'h448e1d71, 32'hc4b66b09, 32'h43225e41},
  {32'h438bc659, 32'hc478146e, 32'hc3d103f1},
  {32'hc245f652, 32'hc5007426, 32'h450c529b},
  {32'hc48f48a8, 32'hc39029cc, 32'hc380d58b},
  {32'h443b23e6, 32'h4300b5a2, 32'h4502fa38},
  {32'hc40bb1c3, 32'hc4e1d1cf, 32'hc2bc6cbb},
  {32'h439ef3f6, 32'hc17c2690, 32'h44946136},
  {32'hc49627fe, 32'hc33e7fde, 32'hc4849af8},
  {32'h44d79103, 32'hc299845a, 32'h446666ec},
  {32'h43f9d45e, 32'hc4bb726c, 32'hc36879c1},
  {32'h44bb0dc3, 32'h4413124f, 32'hc117a3c8},
  {32'hc3e6e74f, 32'h440bd982, 32'hc4d572f7},
  {32'h4251937b, 32'h44456b53, 32'h435f82ac},
  {32'hc481688c, 32'hc2e2a7f8, 32'h426fb760},
  {32'h444f61fc, 32'h4394387d, 32'h44f678dd},
  {32'hc4066659, 32'hc379f7aa, 32'hc2a3cb60},
  {32'hc480dfb7, 32'h426ff569, 32'h43871d1f},
  {32'hc113938b, 32'hc4c917fb, 32'hc50d8def},
  {32'h43eac07a, 32'h44a6dae2, 32'h43abb91b},
  {32'hc43726b4, 32'hc4690f70, 32'hc4280f62},
  {32'h449e0d09, 32'h44dfab1e, 32'h43e55179},
  {32'hc48cefe2, 32'h432026bb, 32'hc378ca7e},
  {32'h44277dee, 32'h42186ded, 32'hc382d558},
  {32'hc45ebf18, 32'hc4ed07d0, 32'h42c4469b},
  {32'h447084f2, 32'h43c314af, 32'h43d677e9},
  {32'hc463e5bc, 32'hc194a831, 32'hc3f40cb8},
  {32'h4476064c, 32'h42bc0411, 32'hc3bc8f58},
  {32'h446169c2, 32'h44557fd8, 32'hc4fef58c},
  {32'h415d0d40, 32'h440743c7, 32'h44969a38},
  {32'h4381c8ec, 32'h449d54f6, 32'hc417f1ff},
  {32'hc48575c6, 32'h4474f1fd, 32'h4481c176},
  {32'h44025dad, 32'hc441b121, 32'hc49525e4},
  {32'h4453bff6, 32'h4395ca56, 32'h4454cf9b},
  {32'h43bff4f3, 32'h415ee64e, 32'hc49376c0},
  {32'hc4b408ae, 32'h438cd343, 32'h44c92265},
  {32'h45025879, 32'hc34faa9b, 32'hc240f19d},
  {32'h434ad0b3, 32'h432fd856, 32'h44c34662},
  {32'h44efc9f0, 32'h43086bd0, 32'hc3aaf9ff},
  {32'h4288092c, 32'h4489c1c8, 32'hc3873f48},
  {32'h451f1f6a, 32'hc3bd7916, 32'hc372e2da},
  {32'hc3b7793a, 32'h44023737, 32'h451067da},
  {32'hc4f0aa7b, 32'hc25bd948, 32'hc2469dfc},
  {32'hc37f87c8, 32'h43fcf14f, 32'h45194ca0},
  {32'h422e96d8, 32'hc3b7cdfd, 32'hc4844775},
  {32'h44a80a34, 32'hc2630728, 32'h43b54ba7},
  {32'h4421b842, 32'hc549eaf2, 32'h409d89d4},
  {32'hc4c7dd7e, 32'h42c15e31, 32'h43f40eb3},
  {32'hc4a461b9, 32'hc3fca824, 32'hc3290849},
  {32'hc41e04f6, 32'h455dd948, 32'h43094f4c},
  {32'h43c17568, 32'hc4de82b4, 32'h430d88de},
  {32'hc3ff223c, 32'hc4580275, 32'h42ad6e4d},
  {32'h445e9900, 32'hc376c140, 32'h43bb2701},
  {32'hc55af9f8, 32'h4405a6d6, 32'hc3e6524f},
  {32'h44b9ef3b, 32'h434da19d, 32'hbfb493c0},
  {32'hc4ad8444, 32'h4308c45c, 32'h43b738d0},
  {32'hc4d6fbf8, 32'h43231439, 32'hc506b9be},
  {32'h433fbce0, 32'h44143a7d, 32'h4265ee72},
  {32'h445fec32, 32'h43a66dd4, 32'hc3999280},
  {32'h449b8a54, 32'hc4a0cdc5, 32'hc4051894},
  {32'h436618e0, 32'h44944cf0, 32'hc303e89f},
  {32'h4548877a, 32'h43a7bed6, 32'h43c27d24},
  {32'hc573a394, 32'h43822494, 32'h434b936d},
  {32'h44bdf274, 32'hc4bfde88, 32'h43cafd03},
  {32'h44124f2e, 32'hc3258dce, 32'hc3e67274},
  {32'h4405a5b8, 32'hc49db452, 32'hc471b25d},
  {32'hc46459fe, 32'h432d6f32, 32'hc4c450e2},
  {32'h43188a2d, 32'hc488c432, 32'hc3989051},
  {32'h43c68fbe, 32'h43a6527d, 32'h449849b6},
  {32'h441ff1b2, 32'hc3cace69, 32'hc53e3e11},
  {32'h43b69d84, 32'h42c2d69c, 32'h44972f9f},
  {32'hc3a66f71, 32'hc380098c, 32'hc50de804},
  {32'hc3badf0a, 32'h44689204, 32'h4493488f},
  {32'h453b1b27, 32'hc3192d5d, 32'h43e0034e},
  {32'hc54615c2, 32'h4372d1c6, 32'h417ce101},
  {32'h45335a22, 32'h43d8dfa3, 32'hc337c958},
  {32'h42e7cd7a, 32'h41d59507, 32'h43b1a32a},
  {32'h43a2393a, 32'hc3ddbb76, 32'hc3cc591d},
  {32'hc5144d22, 32'h430bbb44, 32'h423d83f4},
  {32'hc20e3a40, 32'hc45f3532, 32'hc3bbc9d9},
  {32'hc4df1603, 32'h43bd2d8c, 32'h448cf31d},
  {32'h44fd91fb, 32'hc31a89be, 32'hc437cac4},
  {32'h43ce4a94, 32'h43819fb2, 32'hc367dd7d},
  {32'hc53c0d7e, 32'h43810644, 32'h413d7a7c},
  {32'h42e9df15, 32'h42cd8998, 32'hc2d6d368},
  {32'hc41a5a68, 32'hc3a26132, 32'hc3c10f8c},
  {32'h44556eb9, 32'h4485fe51, 32'hc2da2c74},
  {32'h4402cbb9, 32'hc4dfe9ad, 32'h4378d2bc},
  {32'hc2b64ef0, 32'h456f16d5, 32'hc3765d47},
  {32'hc3df18c1, 32'hc50d63ff, 32'hc45f20ea},
  {32'h42fce7f2, 32'h4339e5f1, 32'h439cadf6},
  {32'hc500a80b, 32'h42c28f7d, 32'h42ee6b8c},
  {32'h45489413, 32'hc21c826f, 32'hc2452c84},
  {32'hc3dbff6a, 32'hc37e23bf, 32'h43d86fef},
  {32'h439ee6a4, 32'h45050ec3, 32'h4427d8cd},
  {32'hc440420c, 32'hc41ae8e7, 32'hc4ba0a5d},
  {32'h448d57ea, 32'h431006a4, 32'h4381eeff},
  {32'hc50e83f8, 32'hc3e83b9e, 32'h42edb504},
  {32'h430c8752, 32'h438ff576, 32'h4500e942},
  {32'h448ecc75, 32'hc42bcfac, 32'hc3eea1fe},
  {32'h44991f2e, 32'hc4889724, 32'h44d94ebc},
  {32'hc58bd84e, 32'h430606bd, 32'hc363ac24},
  {32'hc4bae1b6, 32'hc34a9695, 32'h43205f1e},
  {32'hc31d5db0, 32'hc4b7e148, 32'hc480c805},
  {32'h4318c712, 32'h44066a8b, 32'hc3bea14c},
  {32'h44859b7f, 32'h43797153, 32'hc40881db},
  {32'hc20f5fe0, 32'h453445ea, 32'h4326b3ff},
  {32'hc53ff2a0, 32'hc1fc0322, 32'hc323dd98},
  {32'hc29ff65e, 32'hc3b8ce77, 32'h436d82c9},
  {32'hc3b4c98a, 32'h4505da6c, 32'h43d23903},
  {32'hc4e5efd8, 32'hc4079189, 32'h43e2f062},
  {32'h45042be4, 32'h449afb75, 32'hc29e38c7},
  {32'hc44d4450, 32'hc445a581, 32'h4411ae2d},
  {32'h433d2fb4, 32'h45832253, 32'hc0f9dda2},
  {32'hc3f6f635, 32'hc3ed5be3, 32'hc3cc52b1},
  {32'h454a4a38, 32'h4388c74f, 32'hc280a60a},
  {32'hc507d38f, 32'h43aa3a83, 32'hc3ae4ff8},
  {32'h44bd3c48, 32'h43ca1738, 32'h438f0f81},
  {32'h43b0141b, 32'hc4df0a03, 32'h422abe52},
  {32'h423f621f, 32'h4519d84a, 32'h432038a5},
  {32'hc379293b, 32'hc401aec0, 32'h450a8fae},
  {32'hc4a8bd5a, 32'h43ac565f, 32'h4376f155},
  {32'hc4499311, 32'hc4a52f1d, 32'h43d5a5aa},
  {32'h43ffa329, 32'hc2f10548, 32'hc533d06b},
  {32'h43767948, 32'h426045a0, 32'h4448ecd3},
  {32'h443781b1, 32'h4450d46a, 32'h434d0138},
  {32'hc401e4aa, 32'h43d132cb, 32'h41d81480},
  {32'h44e3738f, 32'h4421029a, 32'hc3323670},
  {32'hc3d19860, 32'hc4b6c7d1, 32'h442f1f20},
  {32'h45101c81, 32'h44596717, 32'hc41e6032},
  {32'h4464a257, 32'hc457ea67, 32'hc42acb5a},
  {32'h4309bbcb, 32'hc3ad6511, 32'hc53fa705},
  {32'h4315c600, 32'hc5438405, 32'h4219254a},
  {32'h44e0286a, 32'h438d6301, 32'hc3d97143},
  {32'hc501b6fc, 32'hc352f90c, 32'h447bc7fd},
  {32'h45017100, 32'h4370dd8e, 32'hc47cf0b3},
  {32'h4402eb30, 32'hc49fce1c, 32'h42e99d25},
  {32'hc3cc7f20, 32'h449bbb74, 32'h43a9f8b8},
  {32'h44e9a386, 32'h43bd99b9, 32'hc2e3731b},
  {32'hc3b31f40, 32'h450b09be, 32'h43f18f4b},
  {32'h43d6bb86, 32'hc516eedf, 32'hc3029a32},
  {32'h43f12a2e, 32'h4524c4fb, 32'hc2d55fce},
  {32'hc1a17900, 32'hc42e458e, 32'hc4955727},
  {32'hc42d7480, 32'h44365d88, 32'h43f8801f},
  {32'h43fb962c, 32'hc2752b33, 32'h43908a0e},
  {32'hc3e6e3f7, 32'h440afc1f, 32'h4284a614},
  {32'h442277c4, 32'hc32487e2, 32'hc4453a79},
  {32'hc40af55a, 32'h4467de8b, 32'h431706dc},
  {32'h444abbe2, 32'hc4ed35e5, 32'h4022c052},
  {32'hc5126a05, 32'h43b19892, 32'hc427325c},
  {32'h447da066, 32'hc3e01eb7, 32'h434f3bc3},
  {32'hc3dc59d4, 32'hc3d109ad, 32'hc502d2c7},
  {32'h452ba7df, 32'hc45b33d8, 32'hc3210150},
  {32'hc2fddb18, 32'hc30a1d4c, 32'hc48cb098},
  {32'h452e758e, 32'hc3737c77, 32'hc39fa359},
  {32'hc401f050, 32'h449cdcc8, 32'hc52f2a00},
  {32'hc404a650, 32'hc450aee0, 32'h437cb9fb},
  {32'hc3af4c33, 32'h44920a46, 32'hc381a0a4},
  {32'h4319da80, 32'hc492d0a2, 32'h42d0f366},
  {32'hc53dc248, 32'hc173b791, 32'h438f0765},
  {32'hc2c975e2, 32'h4407bb79, 32'h4548e5cd},
  {32'hc50165a3, 32'hc418ee52, 32'hc4a4204d},
  {32'h44030c1d, 32'hc3b789c6, 32'h441f76b7},
  {32'hc403163a, 32'hc4b16ded, 32'hc4c8ec27},
  {32'h44cf78cc, 32'hc2eee6a0, 32'h43a01794},
  {32'h436686df, 32'hc400c655, 32'hc4942e92},
  {32'h432e1902, 32'h43b83f81, 32'hc4bea276},
  {32'h44ded53a, 32'hc48a1b36, 32'hc38baf14},
  {32'hc48d43cc, 32'h4310eff5, 32'hc3ce99b9},
  {32'hc3af27be, 32'hc3a8175c, 32'h44782c5e},
  {32'hc39c8987, 32'h44536071, 32'hc456bc5a},
  {32'h44190db8, 32'hc40cfc34, 32'h44e4d26e},
  {32'hc3d118db, 32'hc4df5440, 32'h450a796d},
  {32'hc5042042, 32'h44384f8b, 32'hc4829aa3},
  {32'hc456f982, 32'h440d891b, 32'h4407ab4f},
  {32'h420316f6, 32'h435981f2, 32'h44d63709},
  {32'hc31eab67, 32'hc3cbb19c, 32'hc3d5f337},
  {32'h44080cab, 32'hc3dc5e8c, 32'h442daf45},
  {32'hc503efe9, 32'h439008cc, 32'h42cf81bf},
  {32'hc317e6ba, 32'hc50e66c0, 32'hc40430e9},
  {32'hc32cd91c, 32'h424f6249, 32'hc36e120d},
  {32'h4554165f, 32'hc431cce9, 32'h426a59e9},
  {32'hc462ccb8, 32'hc3d1f0fe, 32'h43cff378},
  {32'h44b9f61b, 32'hc417b67c, 32'hc212e297},
  {32'hc5161694, 32'hc3b38859, 32'hc39f4534},
  {32'h43b03798, 32'hc42eeca5, 32'hc39db26e},
  {32'hc48b787a, 32'h440f5cc1, 32'hc13c0996},
  {32'hc46a7b5e, 32'hc3d69ad7, 32'h43074506},
  {32'hc3705290, 32'h4500eaa6, 32'h3e82321c},
  {32'h4446a450, 32'hc4986246, 32'hc030b11e},
  {32'hc42ce828, 32'hc3ecfb0d, 32'h43136ccc},
  {32'h43e06767, 32'hc4314642, 32'hc46aa32d},
  {32'hc271d5f0, 32'hc4b8718f, 32'h44b390d4},
  {32'hc4d6c27d, 32'hc271c6f5, 32'h43a8392d},
  {32'h44fd048c, 32'hc2380c0b, 32'h433197c3},
  {32'h448689b6, 32'h432e3112, 32'h44084810},
  {32'h430e40cb, 32'h4514b9e6, 32'hc480dada},
  {32'hc2a5fe5e, 32'h42f4fb51, 32'h45381811},
  {32'h44380e90, 32'h448e8178, 32'h43a39e55},
  {32'h4366f6f4, 32'h44507f1b, 32'hc3afba7e},
  {32'h43dd8128, 32'hc50f03f2, 32'h450f2c05},
  {32'h44656428, 32'h443d66f0, 32'hc47ffad0},
  {32'h43ee2381, 32'h4534d474, 32'hc3155842},
  {32'h43062aca, 32'hc3e495e8, 32'h44ec1010},
  {32'h43eaa2a0, 32'h44d87bba, 32'hc36ab45a},
  {32'hc5280428, 32'hc3eb87d2, 32'h4450c9e3},
  {32'hc29d4980, 32'h421f9fb0, 32'hc53c1588},
  {32'hc50ecd3e, 32'hc3bdd5e4, 32'hc2b8d155},
  {32'h454ca183, 32'hc3609fbc, 32'hc368cec4},
  {32'hc4e2ae5c, 32'h43220ebb, 32'hc3e1623d},
  {32'hc421bf02, 32'h432e83e1, 32'hc3a83f3c},
  {32'hc260a2e0, 32'hc573c97a, 32'h433600ed},
  {32'h437692fa, 32'h4531d6ea, 32'h43bf5fcb},
  {32'hc306313e, 32'hc4f38180, 32'hc2d770ae},
  {32'h453192ec, 32'h44260e77, 32'hc37056fe},
  {32'hc3ddcf74, 32'hc5190c7c, 32'hc3595b03},
  {32'h43276903, 32'h43a793dd, 32'hc3ae5512},
  {32'h42358ab8, 32'h43fe0e2a, 32'h4338a16c},
  {32'hc3d34444, 32'hc502ea63, 32'hc3811a3b},
  {32'h4397d3dc, 32'hc3cf6360, 32'h44a9eb3b},
  {32'hc5160194, 32'h44011a46, 32'hc3c80b46},
  {32'h4416ce9c, 32'h4420af60, 32'h447824ef},
  {32'hc5377955, 32'hc2d230b6, 32'hc413a246},
  {32'h44893b43, 32'hc2ddd9da, 32'hc38f92ee},
  {32'h42ba746b, 32'hc3ddbc87, 32'hc4fb99d7},
  {32'h4521adc4, 32'hc0060c7a, 32'h4355ed68},
  {32'hc335ca53, 32'hc48b0c10, 32'h4258b6b1},
  {32'h440d2dce, 32'h44bc4cb5, 32'h440a1953},
  {32'hc4538f78, 32'hc3850cf1, 32'hc3a5c6d6},
  {32'hc47ef5ee, 32'h4304c514, 32'h44080ed7},
  {32'hc43f0ab0, 32'hc4c3258a, 32'hc3947323},
  {32'h440ce032, 32'h42b47103, 32'hc251cb6d},
  {32'h44fccb60, 32'hc3695991, 32'h42850886},
  {32'h4492dc02, 32'h43dde1c5, 32'h44c41312},
  {32'hc4ae4b38, 32'hc418c27a, 32'hc4422c56},
  {32'h44456116, 32'h4489af06, 32'h43450170},
  {32'hc4600782, 32'hc51d2680, 32'h43833c00},
  {32'h4491c5ec, 32'h450be442, 32'hc261c1a6},
  {32'h435e3234, 32'hc3924862, 32'hc3ceba1a},
  {32'h44922f45, 32'h44c5934c, 32'h440035f1},
  {32'hc3b19340, 32'hc52abd0b, 32'hc31111d5},
  {32'hc4839592, 32'h42cf7bbe, 32'h435194d6},
  {32'hc484a8a4, 32'hc3bd0f88, 32'hc4115124},
  {32'h456f9bc8, 32'h437662f8, 32'hc3b4f30e},
  {32'h44ca6fc0, 32'hc45cde83, 32'hc30de288},
  {32'h4398bf23, 32'h44dac62f, 32'h4404bab3},
  {32'hc32a5c8e, 32'hc29b5822, 32'hc3d6a5fa},
  {32'hc504a9cb, 32'h43f0c3a2, 32'h43db5386},
  {32'hc392de90, 32'hc491af73, 32'hc38012c2},
  {32'hc479e4aa, 32'h426d3fb0, 32'h43088686},
  {32'h41f38600, 32'hc5084568, 32'hc4f5a1d8},
  {32'hc2459730, 32'h44dd320e, 32'h44c7eca4},
  {32'h45318c7d, 32'hc2a06714, 32'h42d1e058},
  {32'hc304fe84, 32'hc4e42a10, 32'h450fd57c},
  {32'hc3ebb1e1, 32'h446a09b5, 32'hc55464e6},
  {32'hc109bcf0, 32'hc31a3a67, 32'h4497c8d2},
  {32'h448728bc, 32'hc3e28ff0, 32'hc16e39d8},
  {32'hc3352fe7, 32'h43494369, 32'h4564aa1c},
  {32'hc427d40b, 32'hc4c909ae, 32'h4214e906},
  {32'hc2598444, 32'h441f504a, 32'h444e3fe7},
  {32'h41836d20, 32'hc0684dc4, 32'hc559873c},
  {32'hc31e49e0, 32'h43a71841, 32'h444d3b35},
  {32'h4402aea0, 32'hc4fff0a7, 32'h4411cfa7},
  {32'hc55aaa8a, 32'h4284bd3c, 32'h442ff2f6},
  {32'hc48d8417, 32'hc2b68048, 32'h4315b03f},
  {32'hc414fd14, 32'h450d76ef, 32'h42c710dd},
  {32'h44f082fc, 32'hc4b4cc4f, 32'h439333a2},
  {32'h45033bab, 32'h42ba9a13, 32'hc321a8cc},
  {32'h4568baf5, 32'hc31da737, 32'h4391f0f1},
  {32'hc49e893a, 32'h437cd515, 32'h42e50b35},
  {32'h454a9702, 32'hc3b5fd14, 32'h41a2dab0},
  {32'h440c01ce, 32'hc339e2ff, 32'h4518ba3c},
  {32'hc45c088d, 32'hc272a7aa, 32'h41b01328},
  {32'h448ca77e, 32'h440187f7, 32'h43c53e1d},
  {32'hc4b23723, 32'h43686d48, 32'hc410f188},
  {32'h440358a4, 32'hc45e0ee4, 32'h43106c60},
  {32'hc3935150, 32'h44fd274e, 32'h4253e10e},
  {32'h44add532, 32'h43ed4d67, 32'hc4070ffd},
  {32'hc4510088, 32'h4417efca, 32'hc3e935f6},
  {32'h4459253d, 32'hc4f3b18f, 32'h438d5a7a},
  {32'h449734f9, 32'hc35b9629, 32'hc3cb45bb},
  {32'h421bcf20, 32'h43b67b86, 32'h449e31cc},
  {32'hc49b2879, 32'h43ea0bbb, 32'hc4c0bf69},
  {32'h44c6ae7e, 32'hc2f42f66, 32'hc0829cf7},
  {32'hc464ec22, 32'h44a7fbbb, 32'h43b8890c},
  {32'h44760ca6, 32'hc3e03092, 32'hc46ae5f8},
  {32'h42152fa0, 32'h440181d8, 32'h44dbbf52},
  {32'h43c21108, 32'hc4d53255, 32'hc20a3e39},
  {32'hc3db4ca2, 32'h442d6065, 32'h44da9e5b},
  {32'hc4a793c2, 32'hc2eef9ec, 32'hc3bf8942},
  {32'hc3c0e318, 32'hc4986a29, 32'h44cff173},
  {32'h452d4783, 32'h435c2946, 32'hc42fc94d},
  {32'h43acc9c6, 32'h434234ac, 32'h4391f010},
  {32'hc374d263, 32'hc4987025, 32'hc4bde286},
  {32'hc3363168, 32'h44352f61, 32'h449a0255},
  {32'hc4b1fdc1, 32'hc3d4b729, 32'hc3a9d2bc},
  {32'hc4ed8736, 32'h43a71ad0, 32'h44a1574c},
  {32'h44bf98dd, 32'hc4091ab1, 32'hc4f59235},
  {32'h4516e0bc, 32'h4352b4fd, 32'hc457d511},
  {32'hc3a005d8, 32'h434fe928, 32'h44dd679c},
  {32'hc4926bde, 32'h43406199, 32'hc1fd767a},
  {32'hc46f7bb1, 32'hc4403b69, 32'h436a01f5},
  {32'h4403e0b6, 32'h44fcb224, 32'h42bc1b8d},
  {32'hc3dcf399, 32'hc45e4c8d, 32'hc3179306},
  {32'h43bf1ca0, 32'h44a68db6, 32'h43a83a4e},
  {32'hc444dfec, 32'hc507be2c, 32'hc43cc810},
  {32'hc43d4958, 32'h440352f6, 32'h44036ccb},
  {32'hc4c64abf, 32'h438621c9, 32'hc335f0fc},
  {32'h45179c92, 32'h41426237, 32'h42a894bd},
  {32'hc33c6bee, 32'h421133bc, 32'h44ac08fc},
  {32'h44978d64, 32'h44a34618, 32'h435092b2},
  {32'hc40b8890, 32'hc1cb13e5, 32'hc47fbc01},
  {32'h40f5f800, 32'hc306d590, 32'h44042477},
  {32'hc422002f, 32'hc21b7b43, 32'hc4c9fadd},
  {32'h44f58b2a, 32'h438dd564, 32'h4254bb34},
  {32'hc51a7cdd, 32'hc3b80a8b, 32'hc366b6fb},
  {32'h4492e8a0, 32'h430cafbb, 32'h4386df2a},
  {32'hc52fb5a0, 32'h42638766, 32'hc1dd815a},
  {32'h44433205, 32'h43ac0756, 32'hc422906e},
  {32'h43696d2c, 32'hc4ce4c7b, 32'hc3191838},
  {32'hc295a88a, 32'hc2cc964d, 32'h453cf252},
  {32'h44b5a212, 32'h428428f2, 32'hc392a1c7},
  {32'h4425b2fc, 32'h44db4bb3, 32'h427ad4c3},
  {32'hc5117b86, 32'hc402fb8c, 32'hc413ca72},
  {32'h44a78ece, 32'hc3e0d899, 32'h4326ab75},
  {32'hc2bd8179, 32'h445041f5, 32'h439d73ee},
  {32'hc53ee146, 32'hc386aa0e, 32'hc34ba2bd},
  {32'h430b8af6, 32'h452881cc, 32'h443ec503},
  {32'h43200586, 32'hc425c5c4, 32'h438d0ba3},
  {32'h44635101, 32'h43d9b8ac, 32'h43cb03df},
  {32'hc3a8b0f0, 32'hc4e4beb3, 32'hc2b526e1},
  {32'hc31935fc, 32'h445b3834, 32'h43bcb967},
  {32'hc4aeacaa, 32'hc4b8de7b, 32'hc4908907},
  {32'h450ad72e, 32'h44375e2c, 32'h4455db9d},
  {32'h43b4ac38, 32'hc3c2116a, 32'hc32a757e},
  {32'h44f9e124, 32'h4310016a, 32'h43f7e1e2},
  {32'hc421176b, 32'hc442d7f0, 32'h44a450e7},
  {32'hc480b046, 32'h440d2c5f, 32'hc2cdae9e},
  {32'hc4c8a457, 32'hc286deb6, 32'h40c013ee},
  {32'h443a47b0, 32'h44a5f563, 32'hc45df49e},
  {32'h4490be4a, 32'h43948771, 32'h43b0f4ca},
  {32'h43e6899c, 32'hc2e7a52b, 32'hc4a1163f},
  {32'hc5183a9f, 32'h424d680b, 32'h4290e9b0},
  {32'h448eca0f, 32'h42b0aa5d, 32'h41278084},
  {32'hc44ae638, 32'hc464ca7d, 32'h44f3924e},
  {32'hc3e318d0, 32'h446fa828, 32'hc3bf92fe},
  {32'h43e3f723, 32'h439ea653, 32'h448f11d2},
  {32'hc2974078, 32'h44b7a87b, 32'hc436fd6b},
  {32'hc3bedc34, 32'hc276e0fa, 32'h453155d2},
  {32'h451faa4e, 32'h43b5d0fa, 32'hc3372901},
  {32'hc50886c8, 32'h441f8225, 32'h44f1e7d1},
  {32'h4401a508, 32'hc452b4fe, 32'hc4c808d8},
  {32'h44bfd6ad, 32'hc44e0a37, 32'hc4109262},
  {32'hc4c1f0f0, 32'h44824fd5, 32'h43196dc8},
  {32'h434a28d0, 32'hc4322d55, 32'hc32957e2},
  {32'hc407b0a6, 32'h4506e6be, 32'h436546ef},
  {32'h443f13f0, 32'hc501d697, 32'hc2be5ca1},
  {32'hc4fdf352, 32'hc3944354, 32'h42dd597e},
  {32'h44c397fc, 32'h439b20c0, 32'h43fd0346},
  {32'hc52511d0, 32'h43d05425, 32'h442749b6},
  {32'h449bdb2c, 32'hc3c90a66, 32'h43896059},
  {32'h43ec27ca, 32'h45445834, 32'h4391eec8},
  {32'h4478996a, 32'hc426f407, 32'h43069c17},
  {32'hc2f65334, 32'h44d5ae19, 32'h43612c4d},
  {32'h44a210ef, 32'h42875465, 32'h44504b09},
  {32'hc401029d, 32'h44c7f59d, 32'h41b05ed8},
  {32'h427e5421, 32'hc45484b5, 32'h43ac28ba},
  {32'hc505b7f7, 32'hc326da2f, 32'hc466be50},
  {32'hc0ce5940, 32'h43fb107e, 32'h454e9077},
  {32'h4457b622, 32'hc34dbd4c, 32'hc43efbbd},
  {32'h44fb92ee, 32'hc442e387, 32'h43839cf0},
  {32'hc483c365, 32'h44929bc4, 32'hc36904e3},
  {32'hc4bcde3a, 32'hc3080288, 32'h42c5b42a},
  {32'hc2c5043e, 32'h450c0eb7, 32'hc2cfa9d5},
  {32'hc3146cdc, 32'hc4402986, 32'h4508e9a9},
  {32'h449831ce, 32'h4494f992, 32'hc2fd081c},
  {32'h45851484, 32'h4404633e, 32'h42fd0fc2},
  {32'hc4d07eac, 32'h43a912a2, 32'hc4986714},
  {32'hc258dc80, 32'hc407d11e, 32'h446d945a},
  {32'h43b9b3f4, 32'h442095d7, 32'hc53ed273},
  {32'h4413e78a, 32'hc4a1dcce, 32'h441f2cf6},
  {32'hc33b045f, 32'h442d867c, 32'hc466be4e},
  {32'h438637d8, 32'h438e57f2, 32'h43294fbe},
  {32'h442e24d3, 32'hc225e600, 32'h45040f47},
  {32'hc3d341d8, 32'h44048c1b, 32'hc4c60727},
  {32'h4273708f, 32'hc4b1e2da, 32'hc393c994},
  {32'hc3876d38, 32'h42c2dba4, 32'hc5268cbe},
  {32'h43fc8e58, 32'hc47bddbc, 32'h44feb18a},
  {32'h438d0982, 32'hc4309bdb, 32'h44ea38a2},
  {32'hc3686786, 32'h44f40a48, 32'hc4f3b732},
  {32'hc264d106, 32'hc40f17e0, 32'h449e7e62},
  {32'h44a34765, 32'h43a601f3, 32'h434c9c60},
  {32'hc52d9050, 32'hc34c0293, 32'h4392235d},
  {32'h44cb9337, 32'h42d2cc2c, 32'hc3adf5f5},
  {32'h43514ab4, 32'h448f8493, 32'hc3176a01},
  {32'h440e9da3, 32'hc47d550d, 32'h4497247b},
  {32'h437fd008, 32'h442fd30e, 32'hc3ab2ce7},
  {32'hc4259292, 32'hc352c8f6, 32'hc32658fb},
  {32'hc53a9473, 32'h440268e0, 32'hc41d69f3},
  {32'h453ffae6, 32'hc30692f2, 32'h44129475},
  {32'h442bdc37, 32'h42dcf283, 32'hc41bbfd9},
  {32'h43d02b7c, 32'hc52438ec, 32'hc44ffef0},
  {32'hc37cfb86, 32'h4569c847, 32'hc23e291e},
  {32'h437a8868, 32'hc4c3afed, 32'hc41c0f7f},
  {32'hc4537fa6, 32'h4454eda1, 32'h4362ce9b},
  {32'h44b9b786, 32'hc4c20f29, 32'h441e0ee8},
  {32'h44106c45, 32'hc2b823d0, 32'h4431310a},
  {32'hc4393ea4, 32'hc4424e82, 32'hc5169f6b},
  {32'hc38bc9b6, 32'hc23ab2ad, 32'h45322c1e},
  {32'hc528998b, 32'h42dc5440, 32'h443d3b4a},
  {32'hc2ccdb14, 32'h44973d84, 32'hc25771d2},
  {32'hc50b9376, 32'hc21c8840, 32'hc38a5d01},
  {32'h4413ddfc, 32'h4400b562, 32'hc4bf89dc},
  {32'h423d5160, 32'hc50ed21a, 32'h4414c838},
  {32'hc36dd5d1, 32'h43505209, 32'hc41752bb},
  {32'hc21e229c, 32'h44c9c480, 32'hc3e5b9f2},
  {32'hc38f0560, 32'h431975e0, 32'h4511ac2c},
  {32'h43d9694d, 32'hc1a98590, 32'hc4e9769f},
  {32'h44762ad4, 32'h4395df44, 32'h42b13934},
  {32'hc4d191f3, 32'h435c8c73, 32'h4463bece},
  {32'h44956ad6, 32'h4300382e, 32'hc45a126c},
  {32'hc41854a8, 32'hc28d4fb0, 32'h452be053},
  {32'hc3b139fe, 32'hc30a520b, 32'hc53fe493},
  {32'hc422e026, 32'hc2ffe11c, 32'h4362c862},
  {32'h44f5d775, 32'hc2128734, 32'hc40e246e},
  {32'hc3ae702a, 32'h444f5a51, 32'h44202edf},
  {32'hc41e1ec7, 32'h4381c3aa, 32'hc33af690},
  {32'hc43de9f3, 32'hc40789fb, 32'h442e142b},
  {32'h45784410, 32'h40c62478, 32'h43804e61},
  {32'h433fe9c5, 32'hc4557207, 32'h436875d2},
  {32'h448295f4, 32'h44d417c1, 32'hc3d41b0c},
  {32'hc4eed761, 32'hc46c63ee, 32'hc36312ec},
  {32'h43550881, 32'h4170ec1e, 32'hc27141d1},
  {32'h45054411, 32'hc43eebea, 32'hc413b922},
  {32'hc3a49ceb, 32'h434be276, 32'hc42a26de},
  {32'h4447dab4, 32'h440e7d1a, 32'h4469503a},
  {32'hc43a66fa, 32'h43a4400d, 32'hc1af8478},
  {32'h429831bf, 32'h45493431, 32'h441c20c6},
  {32'h438f74ca, 32'hc50d8506, 32'hc478cc00},
  {32'hc410cfc6, 32'hc3d305a5, 32'h43e601e8},
  {32'hc4fdf5fb, 32'hc3929d0f, 32'hc4a04c1a},
  {32'h44905598, 32'h4364bb9a, 32'h44c9ac0c},
  {32'h44019e3f, 32'hc40bdff2, 32'hc488fcde},
  {32'hc465a186, 32'hc39b8c9d, 32'h445f68d0},
  {32'hc469420f, 32'h43abc667, 32'hc434ce9c},
  {32'h44d13579, 32'h43e7e722, 32'h43a07ee4},
  {32'hc462d658, 32'hc459dc00, 32'hc31828b9},
  {32'h43844a9c, 32'h4516e67a, 32'hc33bedc4},
  {32'h44ffcb3d, 32'h4268949c, 32'h42b14aed},
  {32'h4489051e, 32'h43ea9421, 32'h436c5d0e},
  {32'hc3269960, 32'hc3cc3f97, 32'hc564e01b},
  {32'h44818b64, 32'h444039d9, 32'h43d1d31e},
  {32'hc43d8228, 32'hc5310baa, 32'h40d56ea0},
  {32'h442c20c0, 32'h452caafe, 32'h43ebc9ab},
  {32'h43d2fa3d, 32'hc4a7e99f, 32'hc3f8da04},
  {32'h45329ac3, 32'h43d2ae5b, 32'hc32543df},
  {32'hc41a4224, 32'hc500a19f, 32'hc4053061},
  {32'h4443cafd, 32'h43342675, 32'h43f01d4e},
  {32'hc5697cb8, 32'hc2b9e56c, 32'hc1ad449c},
  {32'h42972550, 32'h43788f13, 32'hc37661a1},
  {32'hc35ad482, 32'h43dc985d, 32'hc519bee6},
  {32'hc375afa9, 32'hc483c2ff, 32'h43a12a1b},
  {32'h441aa469, 32'h42d68717, 32'h41636aae},
  {32'hc40a5744, 32'h44fdd9a9, 32'h43344042},
  {32'h442dbc06, 32'hc4c6ad7e, 32'hc37ec919},
  {32'hc315d0e0, 32'h442ddf1e, 32'h44cff034},
  {32'h44a0b644, 32'hc39c475b, 32'hc48a6fd9},
  {32'hc45b0430, 32'h44b1dd5a, 32'h44bdd632},
  {32'hc3c83a2b, 32'hc204cda2, 32'h431b2182},
  {32'hc306e0f2, 32'h443fb8a8, 32'h4489312d},
  {32'h41d6120d, 32'h43c666ad, 32'hc4fa88ad},
  {32'h43b5a520, 32'hc3ceea52, 32'h44f653a0},
  {32'h432823d4, 32'hc50afe79, 32'hc32a0d17},
  {32'hc4badd18, 32'hc2def352, 32'h44790d9b},
  {32'h44555a86, 32'h43a1a192, 32'hc40d26bc},
  {32'hc35e29f8, 32'h42ce14e8, 32'h450a85d1},
  {32'h43f5079e, 32'h430e8273, 32'hc49ffc38},
  {32'hc353ac1a, 32'h448c25fe, 32'h43cb06f9},
  {32'h454197c4, 32'hc385474d, 32'h431ff0c6},
  {32'hc4f2a707, 32'h44dbef42, 32'h4328dd8c},
  {32'h42763ae1, 32'hc1dd89b1, 32'hc2cff06d},
  {32'hc43ea91c, 32'h4518d437, 32'hc34f9e98},
  {32'hc3d034c1, 32'hc5129805, 32'h438a0247},
  {32'h44a6fc80, 32'h43e45581, 32'h41ab5e6a},
  {32'h4534d396, 32'h43e6b819, 32'hc2b3032f},
  {32'hc4b80b40, 32'h43d83cc9, 32'h43b20dd9},
  {32'h4504ed1b, 32'hc4088682, 32'hc45149c5},
  {32'h448152c6, 32'hc3ec37f1, 32'hc3f114dd},
  {32'hc4da8594, 32'hc39a6ed2, 32'hc3bffdc2},
  {32'h450ddc70, 32'h43b4c187, 32'h449c36be},
  {32'h439a06aa, 32'h44135f67, 32'hc3829115},
  {32'hc3241b7c, 32'hc56a1170, 32'h43a1e19d},
  {32'hc482e96f, 32'h44be27bb, 32'hc38f0e2a},
  {32'h43d12c2a, 32'hc4264943, 32'hc0561570},
  {32'hc4e3af28, 32'h4485761c, 32'h42e7da22},
  {32'h440ce090, 32'hc4fe6bdc, 32'h42fae965},
  {32'h44943d56, 32'hc281235a, 32'h42abc235},
  {32'h44988f38, 32'hc13a26b6, 32'h4466899c},
  {32'hc3ec8635, 32'h43e6b1c0, 32'hc5340372},
  {32'hc42c906c, 32'hc3b1c78e, 32'hc28ef2af},
  {32'hc429be18, 32'h43a52a48, 32'hc326acc0},
  {32'h44308ae8, 32'hc4bc7673, 32'hc452b3e3},
  {32'h4487d9a8, 32'h43a25e2b, 32'h42c29f06},
  {32'hc318d560, 32'hc3918652, 32'hc4a7ba6d},
  {32'hc4821866, 32'h43f817ee, 32'h449feb72},
  {32'h4537c5b9, 32'h42f4b337, 32'h43a2d19d},
  {32'hc53bd719, 32'h42e2390f, 32'h433ef13b},
  {32'h43e1d5de, 32'hc47a6b1e, 32'hc4c6f71d},
  {32'h439ff66c, 32'h43bd1025, 32'h443f14a4},
  {32'hc3ee20a2, 32'hc5435aaf, 32'hc423a054},
  {32'hc3ddeddc, 32'h4432978e, 32'h448044ad},
  {32'hc456715e, 32'hc42708b0, 32'hc3bf1d14},
  {32'hc54fafa0, 32'h44091f5a, 32'h4380f25d},
  {32'h44aa7bf2, 32'hc4443853, 32'hc48af837},
  {32'h44ada1e0, 32'hc32a397a, 32'hc4f40161},
  {32'hc5519b8a, 32'hc355ecf8, 32'h42995d31},
  {32'h4502a5d6, 32'h441e6b74, 32'h43f561fe},
  {32'hc4fd84dd, 32'hc4a51b1a, 32'hc448f116},
  {32'h4507f492, 32'hc3da9d5a, 32'hc2322d08},
  {32'hc467ee2b, 32'hc422fc96, 32'hc303d729},
  {32'h441ad910, 32'h44e8f0fb, 32'hc29b43d7},
  {32'hc5180e7c, 32'hc428e535, 32'h43a717bb},
  {32'hc2b0462c, 32'h441a79b9, 32'h428ad578},
  {32'hc4f0ee80, 32'h42c67a7c, 32'h44108c2b},
  {32'h44fb4316, 32'hc382884a, 32'hc4aa8519},
  {32'hc50738af, 32'h4309c559, 32'h434bba4a},
  {32'h42de76f8, 32'hc2c6f858, 32'h4502654a},
  {32'hc4c62edd, 32'hc452b51b, 32'hc49d4c46},
  {32'h428af05b, 32'h44af454b, 32'h44059547},
  {32'hc3526ab5, 32'hc4ee9957, 32'hc41e67dc},
  {32'h42db5ced, 32'h43ba3117, 32'h454a5399},
  {32'h447453be, 32'hc38f2164, 32'hc44100db},
  {32'h448b9a0c, 32'h4414102e, 32'h44494230},
  {32'hc4be80e1, 32'h446e0fa4, 32'hc4899e68},
  {32'h4486b88d, 32'h43c01b36, 32'hc33ead17},
  {32'h43815992, 32'hc41af9ab, 32'h436d5169},
  {32'hc2a99450, 32'h4344705f, 32'h4510f271},
  {32'h4384a804, 32'hc4620ea1, 32'hc35df50a},
  {32'h4214bc8c, 32'hc20570e0, 32'h44d69b88},
  {32'hc4167d02, 32'hc32a9860, 32'hc54b9df0},
  {32'hc3cbba73, 32'hc1c894e1, 32'h4402aecc},
  {32'h4494e074, 32'h430e6640, 32'h41a6535e},
  {32'hc4f0bdda, 32'hc3ef1b62, 32'h43e299cc},
  {32'h44546e11, 32'h450d12ba, 32'hc370e8d5},
  {32'hc52e8b6a, 32'h41b5ce08, 32'h43f48775},
  {32'hc31d7029, 32'h455d33fe, 32'hc2c43792},
  {32'hc3071e70, 32'hc42b54ab, 32'hc30eabc7},
  {32'hc42b2716, 32'h428933dc, 32'hc3a256cd},
  {32'hc4c631ae, 32'h44085901, 32'hc1c6fcba},
  {32'h45565733, 32'hc3931304, 32'h4435012d},
  {32'h42bc8f59, 32'h43456b58, 32'h41fdae5f},
  {32'h4499b1a4, 32'h44237600, 32'hc301b790},
  {32'hc4839b74, 32'h4245168f, 32'hc463488c},
  {32'h4506c416, 32'hc364a690, 32'h42c64394},
  {32'hc4474700, 32'hc3761eb5, 32'h44937698},
  {32'h443522a5, 32'h44e075b9, 32'hc30c3800},
  {32'h43ce6e53, 32'hc28d73c0, 32'h44891f0c},
  {32'h44c8f5ea, 32'h42258518, 32'hc480fc65},
  {32'hc3b611be, 32'h4405f647, 32'h4525b691},
  {32'hc345eb72, 32'h41398a6c, 32'hc480c14c},
  {32'hc4155ff4, 32'hc494017a, 32'h44638af4},
  {32'h43e20548, 32'h44e6bf38, 32'hc415a0c4},
  {32'h43e56970, 32'hc49ee494, 32'h42ad5f66},
  {32'h44ecc899, 32'hbd0d9300, 32'hc38a9794},
  {32'hc4243b61, 32'hc4cdbf5f, 32'h43432f59},
  {32'hc4d97653, 32'h435d7746, 32'hc201d2d3},
  {32'hc43484dd, 32'h4433b8fc, 32'h44c59a31},
  {32'h445551f4, 32'h4364438a, 32'hc35c822d},
  {32'h429dc5ac, 32'hc5319263, 32'h427c86f8},
  {32'hc3d61965, 32'h4546597b, 32'h4386096b},
  {32'h44597418, 32'h4203122d, 32'h43da2b53},
  {32'hc494c3fc, 32'h44a8069b, 32'hc3db0feb},
  {32'h43c07072, 32'hc29f9501, 32'h43f7e89f},
  {32'h44d2408b, 32'hc3321249, 32'hc31913be},
  {32'h44614954, 32'hc44d6b34, 32'hc4af6a98},
  {32'hc4fd90cd, 32'h442bef62, 32'h445f4d4a},
  {32'hc3b3c862, 32'hc30c3dd7, 32'h42d86a02},
  {32'h42b31de8, 32'h441c964e, 32'hc409c542},
  {32'hc236cd60, 32'h4450f30f, 32'hc4c946c5},
  {32'hc4ed81fa, 32'h438e5725, 32'hc41ba04e},
  {32'h451a061c, 32'hc2e5e330, 32'hc3906008},
  {32'hc4fd2060, 32'hc300f6c1, 32'h4057d45a},
  {32'hc4eedcdd, 32'h43c92e9f, 32'h41395e9e},
  {32'hc4bff3ca, 32'h43439cc2, 32'hc3e49f2b},
  {32'h41f7e180, 32'hc43ba104, 32'hc3874d2c},
  {32'hc3d5e5fc, 32'h43225a5c, 32'hc3b79a60},
  {32'h439a9798, 32'hc51a6619, 32'h4391fa86},
  {32'h432e4b28, 32'h4526a20a, 32'hc3078f54},
  {32'hc4689e09, 32'hc4360418, 32'h446b259c},
  {32'hc4fa613d, 32'hc0392f93, 32'hc46743ad},
  {32'h441e0e94, 32'hc526f825, 32'hc2baf75c},
  {32'hc4eb662a, 32'h43ba6069, 32'h430242f6},
  {32'h44ac98c6, 32'hbfc97ce2, 32'h441044e5},
  {32'hc5245cfd, 32'h40ae9959, 32'hc4a4984b},
  {32'h4501ad65, 32'hc3d36684, 32'hc3a3264a},
  {32'hc4a57897, 32'h440eaf43, 32'hc4276979},
  {32'hc3bbe345, 32'hc46ed9ae, 32'h44dd70df},
  {32'h448a6652, 32'h43eac4a7, 32'hc3e873f8},
  {32'h43d8d17e, 32'h43a784bc, 32'hc3c32fb2},
  {32'h4434558f, 32'hc46f3ece, 32'h43a7109f},
  {32'hc2ef5de0, 32'hc3ace09b, 32'hc4de2559},
  {32'h448b75d9, 32'hc3e57c29, 32'h43943535},
  {32'hc3bf12f0, 32'h44cdfcb8, 32'hc469ad35},
  {32'h4302444d, 32'h426770f7, 32'h4534401d},
  {32'h42a63800, 32'h4486ab17, 32'h44e41af8},
  {32'h41cc7e88, 32'hc4233091, 32'hc523e3e8},
  {32'h447aa560, 32'hc3b9fefb, 32'hc22174e1},
  {32'hc43c3df2, 32'hc321aecd, 32'hc2eab315},
  {32'hc10cb400, 32'h455cac0a, 32'hc32e09c7},
  {32'h43181924, 32'hc368c096, 32'h45330646},
  {32'hc4fb7886, 32'h4333cc9d, 32'h440505c1},
  {32'h4451e934, 32'hc3ba1651, 32'h44364669},
  {32'hc3b5396c, 32'hc446f432, 32'hc51133e0},
  {32'hc4478060, 32'hc4481f5a, 32'h42a73be6},
  {32'hc5399dfe, 32'hc3189604, 32'hc3bf0635},
  {32'h454c9088, 32'hc408b9b7, 32'h43820ed7},
  {32'h42c0639d, 32'h43574800, 32'hc3fc0668},
  {32'h44af53f8, 32'hc3c68b8d, 32'h4365784b},
  {32'hc34cc252, 32'h451ac4de, 32'h4331a12a},
  {32'h44e37394, 32'h4094d9ec, 32'h43b3f037},
  {32'hc482b69a, 32'h45229ae0, 32'h4326baca},
  {32'h43ee90a4, 32'hc4cc85ed, 32'hc41ee42b},
  {32'h4351d514, 32'h42dc167d, 32'h4480bd10},
  {32'hc4224b08, 32'hc4d71d6e, 32'hc4cfa9c4},
  {32'hc3a70571, 32'h44a8a537, 32'h4499f5ed},
  {32'h416f0900, 32'hc420902a, 32'h44793cb7},
  {32'h4410ae9e, 32'h4557d4e8, 32'h4429359d},
  {32'hc2d2d330, 32'h43939a73, 32'h44a40613},
  {32'h429a3e40, 32'h4493aea7, 32'hc512ec85},
  {32'h42eeb4f4, 32'hc51858c7, 32'hc32a2142},
  {32'hc4e763d4, 32'hc16695cd, 32'hc3bf4520},
  {32'h45069bdc, 32'h429e74a6, 32'h4401b84c},
  {32'hc40a77c9, 32'hc2543367, 32'h44dda2ed},
  {32'h447f690f, 32'h43561bf3, 32'hc48b07cf},
  {32'h44191029, 32'h447af393, 32'hc40e1580},
  {32'hc502a662, 32'hc3e24015, 32'hc2fa6261},
  {32'hc41df71e, 32'hc174868c, 32'hc436f32d},
  {32'h435c3842, 32'hc4e228cd, 32'h43403003},
  {32'h4303a313, 32'h44b54d6f, 32'hc46233d1},
  {32'h41806a20, 32'hc3d82eda, 32'h44e69762},
  {32'h441d2580, 32'hc3459eb2, 32'hc441528a},
  {32'hc55495aa, 32'hc3288619, 32'hc402a5c9},
  {32'h45545995, 32'h4343a2c2, 32'hc364c7ca},
  {32'hc504faed, 32'hc446dd84, 32'h43f60ecf},
  {32'h44eff542, 32'h43d93946, 32'hc36fe30b},
  {32'h44a0fab5, 32'hc41f2908, 32'hc2162507},
  {32'h44d25e0c, 32'h4448d4a6, 32'hc38628e8},
  {32'hc4c5bbcc, 32'hc47cd4b0, 32'h42befdca},
  {32'hc397f8be, 32'h44455a80, 32'h43671d65},
  {32'h444b78fa, 32'hc3fde843, 32'h441cfd28},
  {32'h41a63746, 32'hc39281b3, 32'hc4e76e75},
  {32'h43556482, 32'h448bb310, 32'h443a78ef},
  {32'h44d7970b, 32'h41219918, 32'h42d50a58},
  {32'h44074112, 32'h441ed402, 32'h44b0839b},
  {32'hc4388d61, 32'hc4585f66, 32'hc4c2926d},
  {32'hc39aa9ff, 32'h42485f82, 32'h43270348},
  {32'h43132f1c, 32'hc4f5d0f5, 32'hc4db2037},
  {32'h442eb776, 32'h44b955a4, 32'h44ad43d9},
  {32'h44aed0a5, 32'hc3fd8768, 32'hc339deb7},
  {32'h43e5b3f2, 32'hc4daa70e, 32'h44e3e358},
  {32'hc409acd5, 32'hc496327b, 32'hc3e9d827},
  {32'h44feb255, 32'h42370e3d, 32'hc279b226},
  {32'hc40c8e6e, 32'hc51e1aba, 32'hc3b76d23},
  {32'h43641e4e, 32'h4473cb03, 32'hc2fa0b69},
  {32'h440995dc, 32'hc463d331, 32'hc4b34210},
  {32'h44a83bbd, 32'h42901a31, 32'h4430dea9},
  {32'h436a9ad0, 32'hc215e8f0, 32'hc4a561c9},
  {32'h451965df, 32'h43ba74e9, 32'h4381a1ee},
  {32'hc4c86ed3, 32'hc3471dcf, 32'hc222fd61},
  {32'h448cac5d, 32'h44ecfb56, 32'hc38a57d0},
  {32'hc4e1e517, 32'h4185d884, 32'h42803f78},
  {32'h44d4679b, 32'h44af0d13, 32'hc257abbb},
  {32'hc46fee99, 32'hc4f70d37, 32'hc23e3330},
  {32'hc33b17e8, 32'h438c8a48, 32'hc27d67e5},
  {32'hc51f4948, 32'hc42568fe, 32'hc27cca1e},
  {32'h4544b61c, 32'h434bbb5d, 32'hc399fdd3},
  {32'hc39a206e, 32'h4506a993, 32'hc4c9fccd},
  {32'hc4801355, 32'h4395edd8, 32'hc2150e90},
  {32'hc2e831c8, 32'hc44b6264, 32'hc2a15cef},
  {32'hc3ed70be, 32'h451a980a, 32'h443b8b7b},
  {32'h44418c70, 32'hc44f7a28, 32'hc215b14c},
  {32'h4326b15a, 32'hc2974110, 32'h440ab77c},
  {32'hc2418d68, 32'h4352f2bb, 32'hc4c0983c},
  {32'hc3f35d74, 32'h44537360, 32'h44804b00},
  {32'hc3266987, 32'hc42e06a1, 32'hc306f0d8},
  {32'h42773bb6, 32'h431c3ac5, 32'h44ea150f},
  {32'hc4b3a06b, 32'h448c1bfb, 32'hc4a9f1d9},
  {32'h4405fa38, 32'h448c5848, 32'hc1931323},
  {32'hc37ecf70, 32'hc501c9a0, 32'hc4044184},
  {32'hc43870be, 32'h44ae0d90, 32'h44293855},
  {32'h43923e54, 32'hc2eb8b5e, 32'hc488e38f},
  {32'hc459cbea, 32'h439aa82a, 32'h44c95b4f},
  {32'h4470f16b, 32'hc46d68ab, 32'hc49ebe77},
  {32'h44048259, 32'h444aa58d, 32'h4448f64b},
  {32'h450a90bd, 32'hc44c641f, 32'h429416f8},
  {32'hc5351260, 32'h44634aec, 32'h422e8dce},
  {32'hc410036b, 32'hc3d276af, 32'hc36e199f},
  {32'hc3cdfcf8, 32'h44e867f6, 32'h43bde29a},
  {32'h4429ec0e, 32'hc3d0289c, 32'hc371c0d2},
  {32'hc38c6911, 32'hc273df33, 32'h42c8da8c},
  {32'h439dfd70, 32'hc3d18d61, 32'hc343048c},
  {32'hc4edbace, 32'hc2750de6, 32'h432011cf},
  {32'h449d3b8c, 32'hc321be10, 32'h42b7e530},
  {32'h449c23d8, 32'hc2a4c8b5, 32'h41abf17f},
  {32'hc48424a4, 32'hc2f4b14e, 32'hc2034d51},
  {32'h4474bd8c, 32'h411c34f4, 32'h452269b7},
  {32'hc382a2ce, 32'h44227148, 32'h44225a72},
  {32'h44613fcc, 32'hc5211e73, 32'hc3018f7c},
  {32'hc51ed851, 32'h444b5fdf, 32'h43762053},
  {32'hc4ac360e, 32'hc3cd28b0, 32'h42a3e19d},
  {32'hc46f2e2e, 32'h4510616c, 32'hc38ca708},
  {32'h449a559d, 32'hc4cb4b35, 32'h42a4759c},
  {32'h45043336, 32'hc2459d01, 32'hc1b3ffe1},
  {32'h44416c67, 32'h438e724d, 32'h41eb9828},
  {32'hc4054fb6, 32'h437966da, 32'hc4260185},
  {32'h445499f2, 32'h41e20a00, 32'hc2e590f1},
  {32'hc454232a, 32'h441e065a, 32'h44812ca7},
  {32'h446e7f3a, 32'hc4b11e91, 32'hc391d2fa},
  {32'hc4f89392, 32'hc280e00e, 32'h42a203a4},
  {32'h452c9c30, 32'h4125a014, 32'hc2e85595},
  {32'hc4973707, 32'hc41357ed, 32'h43c870be},
  {32'hc41c2a49, 32'hc401f865, 32'hc3b28032},
  {32'hc52f6af5, 32'h4390fe5d, 32'h43bd589b},
  {32'h4274b780, 32'hc3190b0d, 32'hc3a78090},
  {32'hc42db1cc, 32'h43cdea34, 32'h4394c5f4},
  {32'h445b95ff, 32'hc4d3a6a4, 32'hc32a3594},
  {32'hc439a452, 32'h44d4243a, 32'h43fd6ca3},
  {32'h4518a6f0, 32'hc3d45cca, 32'hc33dd6de},
  {32'hc2ed86b0, 32'h44daac5d, 32'h44c0677f},
  {32'h42b0bb26, 32'hc4ab459a, 32'hc48594d3},
  {32'hc273ad40, 32'h43df247b, 32'hc390ee36},
  {32'hc43745e4, 32'h4185ff4e, 32'h438b97bd},
  {32'hc46087e9, 32'hc2104aa5, 32'h4356a4ea},
  {32'hc4d7a89f, 32'hc2f1efa6, 32'h440c8fec},
  {32'h435149d4, 32'h453cd4f0, 32'hc28a9680},
  {32'hc4d978b5, 32'h42c1ccc1, 32'hc329b5af},
  {32'h45566d22, 32'h4442bfbc, 32'hc3d3fc25},
  {32'hc48360a4, 32'hc4c4e510, 32'hbf146288},
  {32'h44d2ea89, 32'h42891868, 32'h435f5d8a},
  {32'hc5081955, 32'hc3b18554, 32'hc38e0c48},
  {32'h43a5badc, 32'h440043f7, 32'h442b8098},
  {32'h43ac5ff5, 32'h42d755f8, 32'h43372291},
  {32'hc2867669, 32'h43eb0108, 32'h44e566f5},
  {32'hc4fdce46, 32'hc430c1a2, 32'hc4371009},
  {32'hc2c2f966, 32'h42f43457, 32'h450dcdc0},
  {32'hc194be00, 32'hc42793b4, 32'hc495d180},
  {32'h453a5f10, 32'hc16eb58c, 32'hc2cce0df},
  {32'h4360fac8, 32'hc3e7b031, 32'hc44c1829},
  {32'h452959cc, 32'h43c9f2c9, 32'h4403b67a},
  {32'hc5859aa4, 32'hc39a0ca4, 32'h41fb2712},
  {32'h449f9aa7, 32'h444e0b69, 32'hc35b87f0},
  {32'hc35d0d77, 32'hc20ff5ac, 32'hc4bef954},
  {32'h44364031, 32'h4421db73, 32'h431b65a7},
  {32'h43ce8a2e, 32'hc382538c, 32'hc406a96d},
  {32'h44edf53e, 32'h4421e18e, 32'h440c68b6},
  {32'hc450935a, 32'hc4fb8ec4, 32'hc310d360},
  {32'hc27930a0, 32'h43ee1b2d, 32'h42ce118a},
  {32'h4517a888, 32'hc46ab2d8, 32'hc383f0db},
  {32'hc27fab40, 32'hc4dc6d62, 32'h42820753},
  {32'h44f46664, 32'h4447b6c6, 32'hc3d0b35d},
  {32'h44150485, 32'hc383203b, 32'h43465211},
  {32'h44b86cb4, 32'h4468cae8, 32'hc30d91e3},
  {32'hc3f2cb14, 32'hc4f10769, 32'h43fc4cb9},
  {32'h44f00d73, 32'h43c495b0, 32'hc306f26a},
  {32'hc4eb6914, 32'hc4936407, 32'hc46fb461},
  {32'h449719b9, 32'h44699f24, 32'h4454c41b},
  {32'h44bd3100, 32'h440c63fe, 32'h411fd2bb},
  {32'h43915b34, 32'h44de6db4, 32'h43bf4608},
  {32'hc43eb3ac, 32'hc48383f1, 32'hc42c2a3a},
  {32'hc387329d, 32'h44711e7c, 32'hc3127981},
  {32'hc51b08ab, 32'hc3bffae5, 32'h438b6a57},
  {32'h4456aef6, 32'hc272620e, 32'hc38358b3},
  {32'hc3df5a2c, 32'hc333b26c, 32'h43b152a2},
  {32'h44104181, 32'hc48e6325, 32'hc52f3407},
  {32'hc5373179, 32'h4426ed49, 32'hc35daca2},
  {32'h43c4e302, 32'hc21900b5, 32'hc49d75a0},
  {32'hc362d490, 32'hc48dc52a, 32'h444ff45e},
  {32'h45097b11, 32'h44a255dd, 32'hc4055f9f},
  {32'h429ebc70, 32'hc4bdc07d, 32'hc4120165},
  {32'h44df00a8, 32'h43116433, 32'hc4bc430c},
  {32'hc4a58e75, 32'hc45c5f20, 32'hc34fd4c8},
  {32'hc366571a, 32'h422d0aac, 32'hc492c81f},
  {32'hc3bb1448, 32'h449405e1, 32'h44e74502},
  {32'h44e98682, 32'hc4076238, 32'hc47bcd06},
  {32'hc1bb7400, 32'hc547617d, 32'h4291f4c6},
  {32'hc4b3df2c, 32'h447126d6, 32'h43c28f8f},
  {32'hc4223cf6, 32'hc43b32dd, 32'hc02d1260},
  {32'hc400d74d, 32'h450466e5, 32'h43ee93f6},
  {32'h45241624, 32'hc327ae82, 32'hc3befe8a},
  {32'hc46fb5ca, 32'hc38c13ca, 32'hc3844642},
  {32'h455bdaf4, 32'hc33c8d90, 32'hc4485e2e},
  {32'hc5862d34, 32'h4345cf51, 32'h4412a3a2},
  {32'h443bd279, 32'hc246432d, 32'h439e378d},
  {32'hc3976072, 32'h442b8093, 32'h4197be49},
  {32'h452bab6e, 32'hc2d46063, 32'h43a5234c},
  {32'hc4b5fcee, 32'h43436f3a, 32'hc22f16c9},
  {32'h43031f36, 32'hc49a8e9f, 32'h42fb61fc},
  {32'hc4660b4f, 32'h44aecef7, 32'hc07bbbe2},
  {32'hc4a788f5, 32'hc3f06d13, 32'hc3cb8799},
  {32'hc4186a0e, 32'h4309ff4d, 32'hc4afe347},
  {32'h4405787e, 32'hc3073ddb, 32'h44ecff21},
  {32'hc510315d, 32'h435f3ac2, 32'hc3491e5a},
  {32'h44a7a2cc, 32'hc4833e31, 32'h4473d2b0},
  {32'hc3aaba9e, 32'h4448ed39, 32'hc4a68c0f},
  {32'h441f6051, 32'hc3daeae2, 32'h43e5d39f},
  {32'hc370f138, 32'hc0d64942, 32'hc4454db4},
  {32'h43f80233, 32'hc3ae9b4b, 32'h442fb4dd},
  {32'h44a7c822, 32'h4330651f, 32'hc3f39b42},
  {32'h43d164c0, 32'h432870c6, 32'h44981c49},
  {32'hc3ae2789, 32'hc2ddd061, 32'hc5056d5f},
  {32'hc41879df, 32'h4405cda0, 32'h4493f2fe},
  {32'hc396ccd6, 32'hc4910f12, 32'hc480573f},
  {32'h4423715a, 32'h43bb201f, 32'h44ca27ea},
  {32'h435f891a, 32'hc46f2591, 32'hc38c1684},
  {32'h43e0444c, 32'h43baea74, 32'hc407671e},
  {32'h441f8115, 32'hc4fe6a31, 32'hc1857d8c},
  {32'hc45be3ea, 32'hc30b585a, 32'hc49b1ff6},
  {32'h447b6eed, 32'hc38565b5, 32'hc1e276bb},
  {32'hc42b644f, 32'h43bf4329, 32'hc53ab9a1},
  {32'h44895b70, 32'hc477f18f, 32'h43b171db},
  {32'h420dc5f8, 32'hc4c74bb7, 32'h44f11751},
  {32'h42efd707, 32'h4464b5b5, 32'hc50585f1},
  {32'h4407a22d, 32'hc389becf, 32'hc31cdf88},
  {32'hc3829603, 32'hc4a8a50c, 32'h40994099},
  {32'hc38203af, 32'h4513477d, 32'h43f490be},
  {32'hc23a9280, 32'hc51f154b, 32'hc3ccbb25},
  {32'h44e35d37, 32'h43986999, 32'h43b3dbdc},
  {32'h441486ae, 32'hc4830ab0, 32'h440aecae},
  {32'hc30280e5, 32'h4316f8bc, 32'hc522206f},
  {32'hc4d5934a, 32'h43d63527, 32'h43c0083f},
  {32'hc4b98be2, 32'hc47eb8b5, 32'hc3d269a7},
  {32'h448530d0, 32'hc32cd014, 32'h43f13214},
  {32'h44e2f05f, 32'hc34e49d5, 32'hc3c8250d},
  {32'h43204f5a, 32'hc5192874, 32'hc39919b8},
  {32'hc4572536, 32'h44dcecd8, 32'h439e8426},
  {32'h44438f43, 32'h4385d253, 32'h4309be79},
  {32'hc2e73488, 32'h44ebc951, 32'hc3e86af1},
  {32'h450e41c8, 32'hc43caeed, 32'hc2dbca8a},
  {32'hc4cc9d39, 32'h42f1f908, 32'hc383bf07},
  {32'hc386c3cc, 32'hc4853586, 32'hc4eed8ef},
  {32'hc448c260, 32'hc2997efc, 32'h449f128b},
  {32'hc4371faa, 32'hc4073167, 32'hc17d259c},
  {32'h439540b4, 32'h43af36c5, 32'hc3e04639},
  {32'h433756b6, 32'hc50006e3, 32'hc3176162},
  {32'h43cac1de, 32'h44b0bf9b, 32'hc442bd26},
  {32'h42bd51ee, 32'hc41d9d02, 32'h4499bb4c},
  {32'h43719f04, 32'h43bbcbe4, 32'hc3158680},
  {32'hbf098e00, 32'hc42d2a10, 32'hc47e2b17},
  {32'hc4bab276, 32'h44b90802, 32'h44a93697},
  {32'hc2eed537, 32'h44134f45, 32'hc5385ee1},
  {32'h44143e3c, 32'h4508b99c, 32'h4317dece},
  {32'hc2d85cfc, 32'hc4306450, 32'h44498d57},
  {32'h4525d0c0, 32'hc3b6867a, 32'h42b9bb9e},
  {32'hc41f638c, 32'hc36c8832, 32'h448c6a89},
  {32'h44dad37d, 32'h43efba18, 32'hc2e4c5c9},
  {32'hc3c4f6ce, 32'hc409e95c, 32'h43bbce9e},
  {32'h450e5755, 32'hc385d66d, 32'hc345be6d},
  {32'hc50feca3, 32'h42181512, 32'h44301b39},
  {32'hc4af2915, 32'hc3365db8, 32'hc3313d6c},
  {32'hc4b64c0a, 32'hc466e1bd, 32'h4418a66a},
  {32'h42e23232, 32'h457d43a1, 32'h43bc5570},
  {32'hc500132b, 32'h42e83666, 32'h43d5d91f},
  {32'h42b9bf87, 32'h454769ef, 32'hc31ea82b},
  {32'hc535da36, 32'hc47390d2, 32'h42004027},
  {32'h44ef1ffa, 32'hc3fe11fe, 32'hc226d680},
  {32'hc3d30054, 32'h4467a575, 32'h441f6e44},
  {32'h4371cc48, 32'hc41cff74, 32'hc224ed88},
  {32'h442d8df4, 32'h449fbac7, 32'hc1ed1cac},
  {32'hc3e33564, 32'hc3db2979, 32'hc363ea0b},
  {32'h4504163a, 32'hc34e8d9e, 32'h43907afc},
  {32'hc3d3ab88, 32'hc47fe48a, 32'hc3e8c730},
  {32'hc178a490, 32'h43bae5cd, 32'h44809b35},
  {32'hc34a6eec, 32'hc3c0a75c, 32'h43306f59},
  {32'h42bbcc30, 32'h44f5546b, 32'h44c28e42},
  {32'h43e66a1b, 32'hc4c403e2, 32'h40ba8232},
  {32'h44763f16, 32'h44306a15, 32'h43f67140},
  {32'hc3967f4c, 32'h44430a71, 32'hc49e815b},
  {32'hc41e42e9, 32'h4231e3dc, 32'h4436e978},
  {32'hc38ae1e9, 32'hc209466c, 32'hc54b7267},
  {32'h450a4e4c, 32'h43f90c25, 32'hc3c603cc},
  {32'h43bf0ffc, 32'h420f91e0, 32'h439c8531},
  {32'h44665912, 32'h41f799f8, 32'h44ce02f0},
  {32'hc53da2fb, 32'hc282e10a, 32'hc31f51b8},
  {32'hc4090b11, 32'h441ec288, 32'h43a53c4f},
  {32'h41afaf90, 32'hc572c12b, 32'h43af35dc},
  {32'h44e9f0f0, 32'h44bdf1f1, 32'h44449e2d},
  {32'h44ca6099, 32'hc40acb18, 32'hc3314c31},
  {32'h44b97d7c, 32'h43502e51, 32'h44008efe},
  {32'h4240e49f, 32'hc56f1d28, 32'h4276b7b9},
  {32'h44b43740, 32'h4361bee2, 32'h441841f6},
  {32'hc4f0a1ad, 32'h43e7f5ba, 32'h44157394},
  {32'h443e7350, 32'hc403626f, 32'h43b3e084},
  {32'h43387a28, 32'h448601eb, 32'hc505cc4f},
  {32'hc38c9c86, 32'h45214b3f, 32'h440330bb},
  {32'h43f45d41, 32'h42c5c4c3, 32'hc2d9ed8c},
  {32'h43804fa3, 32'h4456306b, 32'h45011b99},
  {32'h44820cc7, 32'hc480648d, 32'hc3b824c9},
  {32'h423bf300, 32'h43b34066, 32'h444e40bf},
  {32'h4383acf8, 32'hc4a9b5ee, 32'hc4c0b0df},
  {32'hc43cb054, 32'hc33c0f5b, 32'h446ee503},
  {32'h44d787c6, 32'hc1e0dcc2, 32'h43747a23},
  {32'h440677eb, 32'h4508c8b9, 32'h427c7cd0},
  {32'hc3c41c59, 32'h445d28c5, 32'hc4cea7c1},
  {32'hc40022ae, 32'hc47b1bfb, 32'hc2d11e34},
  {32'h43e0782c, 32'hc4a69703, 32'h438f6e00},
  {32'hc52c874a, 32'h43ff36d4, 32'h424fb46f},
  {32'hc39d9dcc, 32'hc3161ac4, 32'hc3923514},
  {32'hc2860a74, 32'h43e70c9e, 32'h455495b8},
  {32'h42867618, 32'hc3aa4075, 32'hc4492c89},
  {32'h43f20747, 32'h43bdefb5, 32'h44ca1e4b},
  {32'h44ed6d97, 32'hc479ed57, 32'hc40c2815},
  {32'hc1707880, 32'h4536fccc, 32'h42a93478},
  {32'h44c54940, 32'hc3b74306, 32'h43696bbc},
  {32'h4206ba2b, 32'h44a53cf3, 32'hc3df2a43},
  {32'h43ceea3c, 32'hc58858ea, 32'h4288c652},
  {32'h440c82d5, 32'h42c66f94, 32'hc37f3f16},
  {32'h44b68f57, 32'h433bf979, 32'h43913a5d},
  {32'hc42e50d0, 32'hc3802dd7, 32'hc4093afc},
  {32'h4460affd, 32'hc4243720, 32'hc3850a25},
  {32'hc4810232, 32'hc2835a58, 32'h43459e4d},
  {32'hc489ec5a, 32'hc39181d6, 32'h43688658},
  {32'hc3cc31b8, 32'h443b10e3, 32'h43ea258b},
  {32'h43aa0290, 32'h3ff55a60, 32'hc3ea091d},
  {32'h43e8e1ae, 32'hc5524a86, 32'hc259c385},
  {32'h41c1d5b0, 32'h453df759, 32'h43c935d9},
  {32'hc40cd3ae, 32'hc2ce7fb2, 32'hc33fc803},
  {32'hc4ad33de, 32'h44a8a166, 32'h42bc7f08},
  {32'h43e28ac0, 32'hc4980c44, 32'h43bcac8f},
  {32'h44c05726, 32'h4269fe2c, 32'h42fdd109},
  {32'h445c35bc, 32'hc35e7efd, 32'h43afd180},
  {32'hc50f9807, 32'h439349f5, 32'hc4449636},
  {32'hc4527dbc, 32'h43055e17, 32'hc3e90918},
  {32'h43cdd0fe, 32'h432101de, 32'h452054d9},
  {32'h44adc30f, 32'hc4454fb0, 32'hc32e6627},
  {32'h4436e690, 32'h44031fea, 32'hc40250ca},
  {32'h44689e40, 32'h43d02702, 32'hc41fdf3c},
  {32'hc4880f32, 32'h4415b6eb, 32'h43f2767f},
  {32'hc4b37652, 32'hc38994d2, 32'hc3c71a3c},
  {32'hc53061bc, 32'hc4885406, 32'h4461681a},
  {32'h45191e06, 32'hc3e0a2b6, 32'hc47272c0},
  {32'h44d105d0, 32'h43d86bc8, 32'h43a05064},
  {32'h441df035, 32'hc48353ad, 32'hc3cb1c6b},
  {32'hc4a2ec6a, 32'h444f3ca1, 32'h44807b38},
  {32'hc410b27c, 32'hc0afdf40, 32'hc39ea959},
  {32'hc37aa7bd, 32'h44897a20, 32'hc270e806},
  {32'h454f074e, 32'hc3e5929a, 32'hc21921e8},
  {32'h43e23294, 32'hc3084956, 32'hc4a15b2f},
  {32'hc4827598, 32'hc05bede0, 32'h438a9423},
  {32'hc46c1b12, 32'h43a3e4ef, 32'h4339e309},
  {32'hc50d3cd4, 32'hc4b547be, 32'hc42061d4},
  {32'h451c0cee, 32'h41957c8e, 32'hc406c040},
  {32'hc3365862, 32'hc2bf7f3c, 32'h435814fa},
  {32'h4552a6f6, 32'h43896828, 32'h42cdca64},
  {32'hc401fea4, 32'hc547f4fd, 32'h4375a789},
  {32'h4486b28e, 32'h40a665d8, 32'h42bc0623},
  {32'hc3f8e622, 32'hc46768da, 32'h4507f31f},
  {32'h44d77440, 32'hc419de41, 32'h43e836ab},
  {32'hc51a0785, 32'h43ae7939, 32'h432746da},
  {32'h44a5faac, 32'h44727240, 32'h41d77bc8},
  {32'hc3973349, 32'hc3c5f113, 32'hc4771424},
  {32'h44243805, 32'h43ca4b06, 32'h42831c04},
  {32'h431138e3, 32'h42bd66a4, 32'hc51d8315},
  {32'h4394e474, 32'h445cdc4c, 32'h449898f0},
  {32'hc494eb3b, 32'h4357f397, 32'h439702cb},
  {32'h43fe3810, 32'h4453ab4e, 32'h44572608},
  {32'hc5170063, 32'hc3b70eca, 32'h42e617fb},
  {32'h45227e58, 32'hc3985c67, 32'hc3ef9ea0},
  {32'hc4fdf34a, 32'hc4112812, 32'hc494f639},
  {32'h44635464, 32'h43e1fcdb, 32'h449d9509},
  {32'h4352edd1, 32'hc3715ee3, 32'hc45a703d},
  {32'h454e44b8, 32'hc385c83b, 32'h430f056f},
  {32'hc486a26a, 32'hc43f8086, 32'hc3d8ab3e},
  {32'h4443f712, 32'hc3a14cc2, 32'h4416c88d},
  {32'h430d4674, 32'h43bf4ffd, 32'hc30c8795},
  {32'hc37bce38, 32'hc4acee13, 32'hc3d521ea},
  {32'h42f5f590, 32'h4546dbe6, 32'hc283b64c},
  {32'hc49ab978, 32'hc40e2a09, 32'h4081181e},
  {32'h4489fa35, 32'h449653cd, 32'hc432b9f8},
  {32'hc409a1ac, 32'hc3042296, 32'h43999952},
  {32'h44c1b624, 32'h432d8702, 32'hc39d0ed3},
  {32'h431edeb0, 32'hc4b8c84a, 32'hc487ba83},
  {32'h452c41c8, 32'h4319384b, 32'h42404b49},
  {32'h4323512e, 32'hc4b10c65, 32'hc31763f8},
  {32'h449bba6a, 32'h434d05dd, 32'h43ee5d85},
  {32'hc38fff22, 32'hc3e7c92e, 32'h450931d2},
  {32'h4452f867, 32'h43cac260, 32'hc3b87eec},
  {32'hc4d1dc25, 32'h41386d14, 32'hc2686252},
  {32'h442b56d2, 32'h43f37315, 32'hc387dea5},
  {32'h449de0b6, 32'hc290efac, 32'h433fbceb},
  {32'h4520cb0b, 32'h4372034d, 32'hc2a6362f},
  {32'hc5481668, 32'hc2e640b2, 32'h438e30c4},
  {32'h450e12e8, 32'hc3904206, 32'hc2d1e79f},
  {32'hc51571e2, 32'hc3fdda71, 32'h449146db},
  {32'h4411aeb6, 32'h45252116, 32'hc1e99fa1},
  {32'hc448cd47, 32'hc4c1bd1c, 32'hc45bc126},
  {32'hc37ede80, 32'hc402a0c3, 32'hc5127076},
  {32'hc3befa80, 32'hc42f0863, 32'h444fb3a2},
  {32'hc4d59ac0, 32'h42fabd01, 32'hc31e1c16},
  {32'hc5582645, 32'h43d47398, 32'hc2f979bf},
  {32'h44a781a5, 32'hc3c95c17, 32'hc4dbe6f8},
  {32'h45182544, 32'hc3acd742, 32'hc3fb56df},
  {32'hc47bddef, 32'h44dc2ee9, 32'h43f702df},
  {32'hc2a5a61b, 32'hc2302698, 32'h442d2df4},
  {32'hc3e6a43d, 32'h44da7db2, 32'h4406530f},
  {32'h447a452c, 32'hc4d23acf, 32'h43eae42e},
  {32'hc46e90b8, 32'h444ac2b4, 32'hc1220902},
  {32'h4441585f, 32'hc4816cd8, 32'hc49fc7b9},
  {32'hc4f08d1a, 32'h41410c69, 32'hc388558e},
  {32'h45322f76, 32'h43674070, 32'h43efca57},
  {32'h42cc6070, 32'hc22d7c09, 32'h445e6073},
  {32'h446f19dc, 32'hc46254bf, 32'h43a9ccc2},
  {32'hc50e4cfa, 32'hc1b1ee40, 32'h4319c75e},
  {32'hc3c74a81, 32'hc44e5a06, 32'h448e28ec},
  {32'hc480e775, 32'hc38f462b, 32'hc4c92954},
  {32'hc4ec07c9, 32'h42f2da2c, 32'hc1ea2c5c},
  {32'hc4936368, 32'h43c1153e, 32'hc3f78fa2},
  {32'h4498e228, 32'hc3fc173d, 32'h44656c7a},
  {32'hc3e7a56d, 32'hc3824501, 32'hc4c04eba},
  {32'h43497a00, 32'hc4b23e6c, 32'h44fc67f5},
  {32'hc3a6cc5d, 32'h44f18deb, 32'hc43d71b9},
  {32'hc4a2e67d, 32'hc39118c4, 32'h40251c33},
  {32'hc356b560, 32'h44be29c8, 32'hc3fcc545},
  {32'hc2468a1c, 32'hc3e1f3d7, 32'h451eef6c},
  {32'h44f6b45e, 32'hc3d15e90, 32'hc32d0011},
  {32'h44727dbc, 32'h43fdb71c, 32'h4505833f},
  {32'hc57b9b7c, 32'hc116e1ee, 32'hc473ed2d},
  {32'h44779bd4, 32'hc3a306e0, 32'h438d2fe0},
  {32'hc4a95e32, 32'hc48df60d, 32'hc45a9880},
  {32'h442fa722, 32'h43c15117, 32'h44709a23},
  {32'hc503b61d, 32'h42f00898, 32'h42233089},
  {32'hc43d5477, 32'h433c4250, 32'hc2db113a},
  {32'h432a0fce, 32'hc5375110, 32'hc3837e14},
  {32'hc47f7ad4, 32'hc3a74744, 32'hc427eac3},
  {32'h451a1454, 32'h442a02e8, 32'h42d4b140},
  {32'hc4de8adf, 32'h438663d0, 32'hc48f350e},
  {32'h43e2dd79, 32'hc3c30d37, 32'h44abbb18},
  {32'h449a7062, 32'hc3c549c9, 32'h4496f0a7},
  {32'hc42fcc2c, 32'h44e1b4cc, 32'hc506ffbe},
  {32'h43465d38, 32'hc3fc9a0e, 32'h446fdfcb},
  {32'h432118b0, 32'hc488aa2f, 32'h4217bd96},
  {32'hc48238a0, 32'h440ea318, 32'h43e4cdc1},
  {32'hc12a54c2, 32'hc45b34fa, 32'h44ac7d76},
  {32'hc43f7ce7, 32'h432c2998, 32'hc378b8ca},
  {32'hc3c99f40, 32'hc4c05a04, 32'h43805eb8},
  {32'hc40b103c, 32'h44a21ac8, 32'h41a1d42c},
  {32'hc4a519a5, 32'hc2460d30, 32'h43125124},
  {32'hc501e849, 32'h43ddc7c0, 32'hc2c0c8a7},
  {32'h45736f1d, 32'h440427ae, 32'h433f4c01},
  {32'hc41b4721, 32'h440178fb, 32'hc1dd5652},
  {32'h4482d9a5, 32'hc50ba1ca, 32'h4400bd99},
  {32'hc4038da8, 32'h4540c5c0, 32'hc334a3ae},
  {32'h436efebf, 32'hc3648c0b, 32'h4389d8a3},
  {32'hc4e90daa, 32'h44cfbf58, 32'h435f2059},
  {32'h44bd9048, 32'hc49c7eaa, 32'h428c80f3},
  {32'hc3d632a0, 32'h43726634, 32'hc37c4a16},
  {32'hc3c23d05, 32'h4420db2a, 32'hc5511a6f},
  {32'hc313e19d, 32'hc4a8bcc6, 32'h452d2041},
  {32'hc22ec9be, 32'hc5012a6b, 32'hc2f3ce68},
  {32'h4337bd1f, 32'h449c4bfd, 32'hc41114da},
  {32'hc49fc7f8, 32'hc391e1a4, 32'hc2cf98ce},
  {32'h44c9a745, 32'h4404622a, 32'hc40139b6},
  {32'hc44cd4e6, 32'hc41f7515, 32'h443650d1},
  {32'h4423f16e, 32'h440ad034, 32'h437c790c},
  {32'h43a2a181, 32'hc2275718, 32'hc4ce5b78},
  {32'hc56c4bfe, 32'h42100874, 32'h4416f0cb},
  {32'h448b2f94, 32'hc4b5ab72, 32'hc43ab714},
  {32'h4537949c, 32'h42bf84ec, 32'hc3b4a3e4},
  {32'hc404a7b4, 32'hc50681d7, 32'hc25646a3},
  {32'hc4a545f4, 32'h43bf251d, 32'h4353cac3},
  {32'hc28ac549, 32'hc50ad894, 32'h40d79861},
  {32'h428a4d96, 32'h44977c30, 32'hc4da7b14},
  {32'h433d6f03, 32'hc357ecb3, 32'h44e4cb67},
  {32'h452cddf4, 32'hc2e6ccf4, 32'hc3dbaa6d},
  {32'hc520cdd7, 32'hc2ebafe2, 32'h44073ef0},
  {32'hc48c3979, 32'h4352e09b, 32'hc323a7ea},
  {32'hc39c1b44, 32'hc5633609, 32'h425a9747},
  {32'h449aef58, 32'h44197ebd, 32'h43074908},
  {32'hc5469c91, 32'h43f10491, 32'h431b1915},
  {32'h42c406c4, 32'h4551731f, 32'hc3e04c72},
  {32'hc5345a10, 32'h4409b60c, 32'h43246874},
  {32'h44161639, 32'h4312da8f, 32'hc3895eef},
  {32'h44c09db8, 32'hc3a8ab77, 32'hc39df147},
  {32'hc4eeb380, 32'h43593435, 32'hc3969d76},
  {32'hc32b839f, 32'h43df0d2a, 32'h44b925ca},
  {32'h41946850, 32'h431e703f, 32'hc4e789a9},
  {32'h450af2d5, 32'h4410c85f, 32'h43eaf33e},
  {32'hc4a68bf4, 32'hc431d970, 32'hc3c3f5c6},
  {32'h3ea13c00, 32'h44ceb718, 32'h43a3a271},
  {32'hc396b018, 32'hc429f326, 32'hc4ed08c8},
  {32'hc21cb400, 32'h44bc27d8, 32'h44b049d8},
  {32'hc2e9c68a, 32'hc488870e, 32'h4329054b},
  {32'h43df52f7, 32'h44f58d87, 32'h42f07a16},
  {32'hc4f020d8, 32'h425ba448, 32'hc397c316},
  {32'h4459c465, 32'h444afb5a, 32'h439e49ad},
  {32'hc500675f, 32'hc3ea14a4, 32'hc2b6bff5},
  {32'h4502c9d7, 32'h4377fd8c, 32'hc3d7b8cd},
  {32'h44ff26e3, 32'h42d66fe8, 32'h43663dc9},
  {32'h448f1edb, 32'h4403766a, 32'h44c837ab},
  {32'hc46a79f8, 32'h42952df3, 32'hc3d1b3a7},
  {32'h453825f4, 32'hc3aab94e, 32'h441133d1},
  {32'hc4060716, 32'hc4e86e16, 32'hc2fcb58c},
  {32'h42489930, 32'h44a905ca, 32'h41a556ef},
  {32'hc3ae5afb, 32'hc3b17993, 32'h42017871},
  {32'h452a0c5a, 32'h4395cd03, 32'h430d3283},
  {32'hc50ddbed, 32'hc43759af, 32'h42d68244},
  {32'hc4f9d714, 32'h4322f582, 32'h43464530},
  {32'hc49bba22, 32'h444bb9a3, 32'h4359270e},
  {32'hc3dd4070, 32'h42a4e0d7, 32'hc381199e},
  {32'h44ccda25, 32'hc3e7a2a1, 32'hc4952278},
  {32'hc3125790, 32'h44995b45, 32'h4490796b},
  {32'h448aa268, 32'h439f42d8, 32'h43655506},
  {32'hc32f464b, 32'h4394e9b2, 32'h451d97ea},
  {32'h45002c44, 32'hc47b3aa7, 32'h43bf4879},
  {32'hc4a84a7d, 32'h43206368, 32'h4395b647},
  {32'h44237762, 32'hc427ea0b, 32'hc5073430},
  {32'hc4887f68, 32'h44a9b9eb, 32'h4435d3bd},
  {32'h4497ee31, 32'h43a13dac, 32'h410141f4},
  {32'h448030dc, 32'hc4eaed10, 32'h44df1abc},
  {32'h4395c910, 32'h43bc993a, 32'hc4b1e0b5},
  {32'h4265d22c, 32'hc4449675, 32'h43eefa83},
  {32'h4483b6f5, 32'hc4237ce7, 32'h42f47ebe},
  {32'hc48c4279, 32'h43d6c9b6, 32'h44abadc3},
  {32'hc3a3bc68, 32'hc398efbb, 32'hc414da5f},
  {32'hc3e09c7e, 32'h441b2218, 32'h44abfeac},
  {32'h4475e5e6, 32'h43af0c61, 32'hc412f8b1},
  {32'hc4aa66aa, 32'h442211f1, 32'h43580a5b},
  {32'h44198e68, 32'hc50cc478, 32'hc31f0727},
  {32'hc4fd47aa, 32'h44467822, 32'h440c6c88},
  {32'h44b89c28, 32'hc314b81f, 32'hc3ad9b4d},
  {32'hc4b11b8f, 32'h44e19eef, 32'hc2786e1a},
  {32'h4344a2fd, 32'hc57ec10e, 32'hc3c4f0e8},
  {32'h44ef98b5, 32'h436ec320, 32'h412a2ad8},
  {32'h44c8c216, 32'hc336644b, 32'hc3f0281c},
  {32'hc597aea2, 32'h4319862a, 32'h43a18aa0},
  {32'h4444e3c7, 32'hc208d7f9, 32'hc34c0d5a},
  {32'hc405709c, 32'hc3265f7e, 32'h44921462},
  {32'hc4fc9835, 32'h4393cba4, 32'hc40b67bb},
  {32'h446cf2b2, 32'hc28ccb99, 32'h44aafac1},
  {32'hc4c20493, 32'h436be2da, 32'hc4275c16},
  {32'h44a0cec8, 32'hc41c71a8, 32'h43a88ebc},
  {32'hc52bba49, 32'h44234501, 32'h43958e16},
  {32'h442c8278, 32'hc3a8f344, 32'h441bace7},
  {32'hc46aaaa1, 32'h4528c6d7, 32'h4311c42d},
  {32'h44390a95, 32'hc52e493d, 32'hc076d7f6},
  {32'hc51491e6, 32'hc3453d4c, 32'hc2c044a1},
  {32'h4400a7a6, 32'h42a3804c, 32'h44aa7df8},
  {32'hc353a8e8, 32'hc2640f23, 32'hc5157ea5},
  {32'h446e2d32, 32'hc36d8bdd, 32'hc381e482},
  {32'hc546e15f, 32'hc3a4dfbe, 32'h43000298},
  {32'h441d112c, 32'hc44446fa, 32'hc37cb23c},
  {32'hc438ee93, 32'h4423ee7e, 32'hc38f971e},
  {32'hc3b7e8ad, 32'h42abfed9, 32'hc5649fa0},
  {32'hc48ce7fc, 32'h40c71c8b, 32'h44b8affe},
  {32'h4490caff, 32'hc33f8a57, 32'hc361e06c},
  {32'hc593b60a, 32'h42a234a1, 32'hc32bc0fd},
  {32'h45454314, 32'h436cdf64, 32'hc44f57c1},
  {32'h431bce82, 32'h43935d2e, 32'hc20a41b2},
  {32'h44042cab, 32'hc3ab2819, 32'hc4273127},
  {32'hc3fbfb8f, 32'h449f8a2d, 32'h428f9db5},
  {32'h42f2991e, 32'h441a60bd, 32'hc4c1ddfb},
  {32'hc5047f61, 32'h448cd82d, 32'hc22db4d1},
  {32'h44e32178, 32'hc42eb72f, 32'hc4c4584c},
  {32'h442bce26, 32'h4433680c, 32'hc4eeb82c},
  {32'hc552bbf6, 32'hc36863c6, 32'h44692838},
  {32'h435a9854, 32'h436fa72f, 32'h43b1240e},
  {32'hc4024e64, 32'hc515f676, 32'hc30dc708},
  {32'h44c77a9d, 32'h441902dd, 32'h43eb6431},
  {32'h449a70c1, 32'hc24086be, 32'hc3278b32},
  {32'hc333d144, 32'h45298aa1, 32'hc39f5668},
  {32'hc555d734, 32'hc414bcdf, 32'h43aa8bb4},
  {32'h44598fe2, 32'h436dbbc3, 32'h429dbca4},
  {32'hc4cfe68c, 32'hc3f76232, 32'h438e3a14},
  {32'h452ac64e, 32'hc3b892a8, 32'hc201ec33},
  {32'h44eb9198, 32'hc3fb0a6a, 32'h43bc31e6},
  {32'h43724832, 32'h44e11adb, 32'h43fec077},
  {32'hc4201046, 32'hc4a0f83b, 32'h4328b476},
  {32'h4415a7af, 32'h41938252, 32'hc3c2f68a},
  {32'hc484fb1a, 32'hc43f8fbd, 32'hc3318792},
  {32'h43a9426c, 32'h43bb9051, 32'h4480d0ae},
  {32'h41e21240, 32'hc472ca47, 32'hc3fda2b0},
  {32'hc3e48853, 32'h438c1813, 32'h43ded9de},
  {32'hc4f8884f, 32'hc4198352, 32'hc45ddabe},
  {32'hc4c54f0a, 32'hc0d62098, 32'hc3008293},
  {32'hc44ce939, 32'hc3133caf, 32'hc3c6ee94},
  {32'hbfce4d00, 32'h4386392a, 32'h44ff92da},
  {32'hc30f2141, 32'h42a21f86, 32'hc433db47},
  {32'hc3c9e8cd, 32'h454454e4, 32'h43b7fd68},
  {32'hc411755b, 32'hc49cdafc, 32'hc38a5908},
  {32'h44ace792, 32'h422e973c, 32'hc3936997},
  {32'h44182bde, 32'hc16ef620, 32'hc43366b3},
  {32'hc4f705f9, 32'hc3197f42, 32'hc367eb7a},
  {32'h40fa9600, 32'h44682745, 32'h44610f44},
  {32'hc54e44c0, 32'h4410d9a6, 32'hc2ac2598},
  {32'h43c2e906, 32'h44fd556c, 32'h41cbbe4e},
  {32'hc4884947, 32'hc4f0afc9, 32'h439fa6a5},
  {32'h455fde73, 32'h4390d102, 32'hc37986f5},
  {32'hc4160e34, 32'hc403afa1, 32'hc2cf1a39},
  {32'h44a7d2f3, 32'h43d6655a, 32'h43a81952},
  {32'hc49c8780, 32'hc36ada4a, 32'h43357aad},
  {32'h451702d4, 32'h43a57b9b, 32'h428ae5ad},
  {32'hc1f05980, 32'hc40a7e8b, 32'hc1a5a57e},
  {32'h43c8567e, 32'h4467956f, 32'hc1a48892},
  {32'hc4a71c6f, 32'hc422ffa7, 32'h430cfa03},
  {32'h43927fff, 32'h432d20a6, 32'hc4e4393f},
  {32'h4467d9f0, 32'hc24994cd, 32'h438f6dee},
  {32'hc354c07c, 32'hc435c972, 32'hc50bfc20},
  {32'hc425ec0a, 32'h438cf06d, 32'h4515122b},
  {32'hc4b9057e, 32'h443bc388, 32'h42e467c7},
  {32'hc5120e51, 32'hc4614bb9, 32'h42f8bf05},
  {32'hc1f3dd00, 32'h44c62caf, 32'hc45ae024},
  {32'h435c5aa0, 32'h437f9f41, 32'h44254ffa},
  {32'h438b5774, 32'h44997e08, 32'hc45615f2},
  {32'h42b3bf08, 32'hc5303992, 32'h4389e401},
  {32'hc4b4f71e, 32'h416e4be8, 32'hc3d9eb04},
  {32'hc4886f49, 32'h4423d1ff, 32'h44bfcfac},
  {32'h431294a4, 32'hc39aae47, 32'hc53f3685},
  {32'h449a2f17, 32'hc49011d5, 32'h4398b443},
  {32'h43d099c8, 32'h45487356, 32'hbfff2dd1},
  {32'h4439d06c, 32'hc3b0729a, 32'hc3a56969},
  {32'hc3ddf1c3, 32'h451564cd, 32'hc3d5fdc5},
  {32'h431bead9, 32'hc54c0b5b, 32'h43c0c243},
  {32'h44ef729e, 32'h430f3f75, 32'h42807e4b},
  {32'h444c0dd0, 32'h42ed502d, 32'hc38ecc6d},
  {32'hc4c06160, 32'h446d2e9e, 32'h444801fb},
  {32'h450cf275, 32'h43217175, 32'h44124c57},
  {32'hc4a63de6, 32'h4370e539, 32'hc14c3ab8},
  {32'h4496da8f, 32'hc2c816cc, 32'h44530c2c},
  {32'h432d240c, 32'h4416a9c3, 32'hc4323b98},
  {32'h4360248f, 32'hc5292f2f, 32'hc29ee8a2},
  {32'h439a8f93, 32'h4482bb84, 32'hc43b35e2},
  {32'h434f912b, 32'hc46edbff, 32'h41cf1564},
  {32'hc45e9e38, 32'h448154d6, 32'hc250f484},
  {32'h422d5080, 32'h427a3bcc, 32'h441ae1c6},
  {32'hc5049c74, 32'hc312ead1, 32'hc3216bc3},
  {32'h44d20801, 32'hc4a88279, 32'hc378b448},
  {32'hc49bd45c, 32'h44cef7a8, 32'hc46a0a1d},
  {32'hc0baf420, 32'hc3ccbb9d, 32'h43ad848d},
  {32'h42b6e231, 32'h45212e7b, 32'hc3363fc9},
  {32'h44cf3ff8, 32'h43a0436d, 32'h43bb7587},
  {32'hc54316d4, 32'h42c84799, 32'h43ad04f0},
  {32'h4423ed20, 32'h424bc797, 32'h44db6d7f},
  {32'hc4c745e0, 32'hc48791f2, 32'hc47b3269},
  {32'h44903969, 32'hc27b20a9, 32'h43cbea64},
  {32'hc1265a34, 32'hc4d5aed8, 32'hc4ff7623},
  {32'hc4c5d5fe, 32'hc41fe2f1, 32'h4490ab4c},
  {32'h43523b19, 32'hc48882f5, 32'hc40d2ce2},
  {32'hc49e4bd0, 32'h43f98fa5, 32'h43cbe43d},
  {32'h43e2e6fa, 32'hc48200e9, 32'h444d22b9},
  {32'hc4945db2, 32'h44902ea4, 32'hc309f2b6},
  {32'hc43ef0c4, 32'hc34307a7, 32'hc2233f76},
  {32'hc47a8556, 32'h4404b15a, 32'hc47c03f7},
  {32'h44b99fd5, 32'hc416660b, 32'h43e9eb0a},
  {32'h43b649d4, 32'hc40b6a8d, 32'h44e521aa},
  {32'hc3ca6535, 32'h450b82a5, 32'hc511238f},
  {32'hc3d0d35c, 32'h44316769, 32'h44ddb0f6},
  {32'hc303ec38, 32'h42bd8e01, 32'h43f40b57},
  {32'hc30b5a3a, 32'h448259c1, 32'hc3049ec3},
  {32'h4511d73a, 32'hc38c5297, 32'h42fde39b},
  {32'h441fd6b5, 32'h43c93bbc, 32'h4418fc8c},
  {32'h44e591e3, 32'h42f0021f, 32'h44740d64},
  {32'hc4b0b0e6, 32'h41968afc, 32'hc105e5fc},
  {32'h44c21024, 32'hc428cd32, 32'hc2da5299},
  {32'hc34e26d8, 32'h4039d79c, 32'hc43bd50c},
  {32'h447c03f8, 32'hc418148e, 32'h440d78ac},
  {32'h45132c7e, 32'h4268c253, 32'hc211d6a4},
  {32'h442f7ff5, 32'hc51aaca5, 32'h43b919d3},
  {32'hc4799754, 32'h44ad23a0, 32'h431e6abd},
  {32'hc4a87e76, 32'hc37b53b5, 32'h43c4adeb},
  {32'hc3af0d3e, 32'h4563e5ff, 32'hc381c478},
  {32'h436a7f4c, 32'hc56c3e7e, 32'hc2f1d1d0},
  {32'hc44c5370, 32'hc3a99ed6, 32'h4373ad46},
  {32'h450d6e11, 32'hc2bb1787, 32'hc10e33ba},
  {32'hc29397b8, 32'h44762394, 32'h44cc21b5},
  {32'hc51d6420, 32'h43f7b481, 32'hc1a43916},
  {32'h4424dd4e, 32'h442c6996, 32'hc3b30585},
  {32'hc52d716e, 32'h41e48d1d, 32'hc36f5f61},
  {32'hc2b86148, 32'h439c5e6f, 32'hc51d862e},
  {32'hc3a982c8, 32'hc54d5447, 32'hc3bc9959},
  {32'h4500c0c6, 32'h43d18ea0, 32'h4368aae0},
  {32'hc2bac718, 32'h4445cb20, 32'hc2222ea3},
  {32'hc18f1536, 32'hc3fb46cd, 32'h45489dc9},
  {32'h434746a6, 32'h44acbb45, 32'hc4ff1293},
  {32'h436d8666, 32'hc2036bdd, 32'hc51cf63c},
  {32'hc4fa69ad, 32'hc3d3a302, 32'h4302d0ca},
  {32'hc22302f0, 32'h4435fb8b, 32'hc280d5f3},
  {32'hc46d1152, 32'hc49dc23f, 32'h4359afe6},
  {32'h440ae754, 32'h43a27700, 32'hc4e3ec05},
  {32'h44a2c5dd, 32'hc3684c18, 32'h438293b6},
  {32'h4420d4c8, 32'h43fdc6a7, 32'hc406aa53},
  {32'hc48a64e2, 32'h42f396c8, 32'h4443703f},
  {32'hc410b2bb, 32'hc2ee58b1, 32'h40ac73d0},
  {32'hc4970bee, 32'hc40b6d3a, 32'hc2d46490},
  {32'h43be6018, 32'h45172874, 32'h443c28ec},
  {32'hc4de14de, 32'hc3819879, 32'h42980292},
  {32'h4522f325, 32'h447d2845, 32'hc3ca0cf5},
  {32'hc465d4cb, 32'hc4d55fe1, 32'h422c4d50},
  {32'hc4b87955, 32'h42e73a8b, 32'hc42166cb},
  {32'h42e7ce83, 32'hc3cc94e1, 32'h445583d3},
  {32'hc3920e0a, 32'hc4563bf8, 32'hc48abaaf},
  {32'hc2f07c4e, 32'h44204100, 32'hc322ff53},
  {32'hc421cc54, 32'hc2809557, 32'hc341c216},
  {32'h44a806d9, 32'h428f6b24, 32'h44b37a7a},
  {32'h43679c02, 32'hc511bdf6, 32'h433dec98},
  {32'hbe127200, 32'h44b25cb4, 32'h4450e5c1},
  {32'hc3a49768, 32'hc392d191, 32'hc4f0dbf4},
  {32'h4516cae5, 32'h42c27d78, 32'h44735af6},
  {32'h42d1187a, 32'hc47db099, 32'h4430a2ce},
  {32'h44e3f674, 32'h43749752, 32'hc38d025d},
  {32'hc41d9f9d, 32'h43d9fc3a, 32'hc4bced27},
  {32'h4555bfa2, 32'h4377cadb, 32'h430d9f8c},
  {32'hc2d57870, 32'hc328924e, 32'hc514a116},
  {32'h433e46df, 32'h45491da6, 32'h4432c1de},
  {32'h43b23e10, 32'hc458b77b, 32'hc4b33147},
  {32'hc3d4f60d, 32'h43cd1550, 32'h455191e2},
  {32'hc40aba17, 32'hc4efb6c0, 32'hc4d32ec8},
  {32'h43aa28a3, 32'h44023be4, 32'h43e9268c},
  {32'hc3ddc640, 32'hc4a49733, 32'h43ecb6a4},
  {32'h43e0d978, 32'h4555e041, 32'hc30d83cc},
  {32'hc4ad6df1, 32'h431fc956, 32'h4384ab1d},
  {32'h452f94ff, 32'h4327d6b8, 32'h431c71df},
  {32'hc3c8fe90, 32'hc3e7ec4d, 32'h43a056ba},
  {32'h44dfe847, 32'h437d3fc5, 32'h4400d3f6},
  {32'hc4a6342e, 32'hc3859ef5, 32'h42eff67f},
  {32'h452d296e, 32'h42d9fca0, 32'h4324246b},
  {32'h42fb22a0, 32'h44833c88, 32'hc5062867},
  {32'h43fb1880, 32'h455a6e9d, 32'h443d2928},
  {32'hc41fc381, 32'h449a1867, 32'hc3226a8f},
  {32'hc41e5059, 32'h449ff2ec, 32'h44c8d2e8},
  {32'h45031889, 32'hc326027d, 32'hc3b17ead},
  {32'hc4992830, 32'h42fd29b2, 32'h441114e4},
  {32'h4431af16, 32'hc42cde88, 32'hc440795e},
  {32'hc48726b0, 32'h42816296, 32'h4494c676},
  {32'h44cdad64, 32'hc42869e4, 32'h41fd618c},
  {32'hc34299c0, 32'hc3f137c0, 32'h44d54c38},
  {32'hc1f45678, 32'hc49f63c2, 32'hc3ee7f79},
  {32'h43ce60d2, 32'h443c4fd2, 32'h43a7b2a2},
  {32'hc343aa37, 32'hc48eda6a, 32'hc415af36},
  {32'hc4a34977, 32'h439cd5bf, 32'h443a632b},
  {32'hc4d99298, 32'h4189ca88, 32'hc35e2e60},
  {32'hc42bdb6f, 32'h445ae10c, 32'h44a970c7},
  {32'h44304680, 32'hc30ebda8, 32'hc3a31169},
  {32'hc457cdd0, 32'h436de670, 32'hc3270744},
  {32'h4301aae0, 32'hc5603a44, 32'h432a4c60},
  {32'hc43addc9, 32'h44624651, 32'hc277273c},
  {32'h450d4149, 32'h4211ba2e, 32'hc36c1229},
  {32'hc4f393f7, 32'h446b6ff3, 32'h41bc6aa0},
  {32'h4531b93c, 32'hc4326cb7, 32'hc38810ec},
  {32'hc3a7e795, 32'h44d9559c, 32'hbe2969c0},
  {32'h450fcede, 32'hc2847e51, 32'h43c94090},
  {32'hc48946b2, 32'h4346d796, 32'h431c6a06},
  {32'hc4a799b0, 32'h42f6173e, 32'hc3fbc132},
  {32'h45370656, 32'hc32cc088, 32'hc2811e34},
  {32'hc34de798, 32'hc280b39d, 32'hc510d107},
  {32'h44090028, 32'h4381a1c3, 32'h4526d1f9},
  {32'h44e5ac24, 32'hc3a62cbe, 32'hc33954f5},
  {32'h438a6b6c, 32'hc50d1aab, 32'hc3ba60ca},
  {32'hc4b0e308, 32'h44597ae5, 32'h431aa94c},
  {32'h4427070f, 32'h43267256, 32'hc302c6bf},
  {32'hc5011af7, 32'h43d25636, 32'hc342a7b8},
  {32'h448b625e, 32'hc4e49b1a, 32'h4311dd1f},
  {32'hc3a05557, 32'h43d63606, 32'hc080520a},
  {32'h44368cac, 32'hc3d1f2a4, 32'h41951dd5},
  {32'hc493c374, 32'hc42bb6c1, 32'h4383af26},
  {32'hc2dbfc44, 32'hc49ed7eb, 32'h4333c021},
  {32'hc2e59f70, 32'h444baf5e, 32'h43866829},
  {32'h43e0e1a8, 32'hc4858837, 32'hc3ccbec1},
  {32'h440a62b2, 32'hc1d9f77c, 32'h43d7486d},
  {32'hc3bc1e93, 32'hc4885dab, 32'hc44be62a},
  {32'hc463907e, 32'h447c8235, 32'h4247f42d},
  {32'hc3bf69c1, 32'hc2ac81ea, 32'hc44108b3},
  {32'hc46c640c, 32'h4430b077, 32'h44b0a5d3},
  {32'h4549ef5b, 32'h433ba6b0, 32'hc44a1457},
  {32'hc389d2ea, 32'h4407133a, 32'h44251fd6},
  {32'hc2ceaa08, 32'hc442339b, 32'hc4a9d185},
  {32'h43997b20, 32'h4500e393, 32'h431682d8},
  {32'h44ce7c50, 32'h432d6175, 32'hc3b7eaab},
  {32'hc2ada4a0, 32'h44177dd4, 32'h44d13769},
  {32'h44407d15, 32'hc4b5db68, 32'hc411acd1},
  {32'h44cdb631, 32'hc3dad93e, 32'hc45db682},
  {32'hc56b1a3a, 32'h436ff892, 32'h43acbce8},
  {32'hc4a7f6ca, 32'hc29371e6, 32'h42dabdc0},
  {32'hc5520797, 32'hc3f61635, 32'hc47eb844},
  {32'h43d0f2e2, 32'h45071827, 32'h44266dea},
  {32'hc19e6cb2, 32'hc4f5d2dc, 32'hc1d551b8},
  {32'hc3966533, 32'h45294c31, 32'hc2e964f1},
  {32'hc3947d02, 32'hc5136c78, 32'hc3198e33},
  {32'h44b4bc97, 32'hc3d4073d, 32'h42f5ab4a},
  {32'h430a0cc0, 32'h4337c200, 32'hc34728ec},
  {32'h442c1de0, 32'h429f6554, 32'hc5093ed9},
  {32'h4421d97e, 32'hc36cfb13, 32'h4397f4e4},
  {32'h44db702a, 32'h43bbf1d2, 32'hc273aac0},
  {32'hc3d6edd6, 32'hc445308c, 32'hc53256e0},
  {32'h43f32c23, 32'h4482b34a, 32'hc33b0978},
  {32'hc493fe43, 32'hc41584f3, 32'h439dd9b8},
  {32'h434a7a12, 32'h4443946a, 32'h440acbe7},
  {32'h450870b4, 32'hc3983572, 32'hc3e27748},
  {32'h43fd40e0, 32'h43ec08d4, 32'h44b7a749},
  {32'hc40980d0, 32'h442f3ccb, 32'hc41d5943},
  {32'hc286acbe, 32'h43487a2d, 32'hc3552617},
  {32'hc2842ffa, 32'hc42e1d11, 32'hc4aabd75},
  {32'h42ecfd54, 32'h44802d86, 32'h43ae467a},
  {32'h4448e367, 32'hc40e58ba, 32'h41890309},
  {32'hc39015c5, 32'h4558308b, 32'h42b8f3a0},
  {32'hc4d6fdbe, 32'hc4520e31, 32'hc3566697},
  {32'h420133b2, 32'hc33f38f8, 32'h4505d928},
  {32'h44386934, 32'h43ec9550, 32'hc407fe46},
  {32'hc361b2ec, 32'hc50fee48, 32'h4321dd34},
  {32'h443fda26, 32'h444f5273, 32'h4443e6e5},
  {32'hc385a708, 32'hc4f3077e, 32'h43b4acd3},
  {32'h44655e40, 32'h4439444b, 32'hc335623a},
  {32'h4274bff8, 32'hc576e00d, 32'h43b57d0f},
  {32'hc46c8402, 32'h44047f06, 32'hc3d96cb6},
  {32'hc48d430a, 32'hc4b3c65e, 32'hc49033f9},
  {32'h42d432cb, 32'hc140bce1, 32'hbfca0289},
  {32'h4446d775, 32'hc3f16e06, 32'h443526f8},
  {32'h444cabc9, 32'hc3255ea9, 32'h4469d809},
  {32'hc46aa9f8, 32'h43834b8a, 32'hc48035db},
  {32'h44a39c47, 32'h4436af3c, 32'hc1c4854c},
  {32'hc4d66710, 32'hc31929fa, 32'h43cd4855},
  {32'h44dd7e57, 32'h43c72227, 32'hc4195ebf},
  {32'h446883c6, 32'h437ec970, 32'h435a96ac},
  {32'h44ab0f71, 32'h43e6b0ac, 32'hc48ae161},
  {32'hc1f43d60, 32'h440b85d0, 32'h4539148c},
  {32'h42374d8e, 32'h43d951d4, 32'hc41a7752},
  {32'hc4cb97d1, 32'hc47b2088, 32'h44a9c08c},
  {32'hc3a57200, 32'h4500b691, 32'hc4251ec2},
  {32'hc48c9a9c, 32'h43700662, 32'h4401c157},
  {32'h44d37f4d, 32'h431a8e54, 32'hc3fbc962},
  {32'hc49dee07, 32'hc5097766, 32'h43fdeadb},
  {32'hc48da64d, 32'h42adced6, 32'hc31b85a7},
  {32'hc5027e63, 32'h41e2728c, 32'h43b4458a},
  {32'hc3481670, 32'hc218edf7, 32'hc52c3153},
  {32'hc2b018e8, 32'hc55f9757, 32'h439db58b},
  {32'hc49eb623, 32'h44de8d8f, 32'h43a6b3e8},
  {32'hc4d31e1a, 32'h435c10c2, 32'h43a55161},
  {32'hc43f8b52, 32'h451b22e9, 32'hc31778ae},
  {32'h444986af, 32'hc4b49fe4, 32'hc33b60b1},
  {32'hc371c48a, 32'h445990fc, 32'hc3543e2c},
  {32'h43ff949a, 32'hc314b83a, 32'h4304d51b},
  {32'hc519735c, 32'h42fba0b2, 32'hc388315a},
  {32'h4533ff27, 32'hc2061be6, 32'h43c7fdc7},
  {32'hc50be408, 32'h44239fb9, 32'hc46a1ecc},
  {32'h44bc38a8, 32'h4425da55, 32'hc41a4941},
  {32'h430c62ce, 32'h43545b92, 32'hc3ffd5ce},
  {32'h43557111, 32'hc5244d08, 32'hc20ce7ba},
  {32'hc490c668, 32'hc2baf985, 32'hc33ee96e},
  {32'h42f9d876, 32'h43ac0523, 32'h45135081},
  {32'hc44e3ef2, 32'h43fa678f, 32'hc40338cf},
  {32'h442cae49, 32'hc3d4dcab, 32'h44156d2b},
  {32'h43d8f6b1, 32'hc3701842, 32'h43f30830},
  {32'h456202a0, 32'hc430fc1d, 32'h43741173},
  {32'hc375e386, 32'h4513974c, 32'hc3ba1719},
  {32'hc3b472e5, 32'hc4928b18, 32'h434481b6},
  {32'hc4493ccd, 32'h4411c9b8, 32'hc43b132a},
  {32'h4321ba14, 32'hc3c87fbf, 32'h45091f2d},
  {32'hc4f3fa45, 32'h44132556, 32'hc38ee454},
  {32'h43c2d608, 32'h447607b2, 32'h453e2b54},
  {32'hc54f9ffd, 32'hc2b65b4b, 32'hc391ad95},
  {32'h44892526, 32'hc28838c1, 32'h43a9f667},
  {32'hc422ec75, 32'h44d06f0a, 32'hc503e349},
  {32'h4506bf92, 32'hc2523734, 32'hc32aaa66},
  {32'h42b77b12, 32'hc3a7731d, 32'hc454ef4a},
  {32'h41e4d854, 32'h44d2ce71, 32'h432b8b68},
  {32'h43df9215, 32'hc49f448b, 32'h43de656d},
  {32'h43a2eeac, 32'h44ec0f59, 32'hc2e7bee5},
  {32'hc36327db, 32'hc3eeca92, 32'h435136dc},
  {32'hc5351d01, 32'h4410d528, 32'hc375b158},
  {32'h43716d94, 32'hc411cf8c, 32'h44f0778a},
  {32'h4435d014, 32'h437f9add, 32'h44af4bcf},
  {32'h4410ebcb, 32'hc4be8da5, 32'hc53178bb},
  {32'hc2b5bda2, 32'h424750dc, 32'h44795b43},
  {32'h446e4844, 32'h40dfde2e, 32'h412749bd},
  {32'h426e816e, 32'h451d0e13, 32'hc38cd7c5},
  {32'hc401cbe1, 32'hc3b6baf7, 32'h44f662fb},
  {32'hc4a4eb6f, 32'hc29bbe3d, 32'hc371292a},
  {32'h43259808, 32'h44174aef, 32'h45513706},
  {32'hc363c714, 32'h431c00d9, 32'hc49173cc},
  {32'h4413bb7d, 32'hc418b85c, 32'h43712d44},
  {32'hc5718369, 32'hc3ba69f9, 32'hc30c8a47},
  {32'h441c197c, 32'h431be5b1, 32'h4439c1cd},
  {32'hc3805fdd, 32'hc3ab3cd4, 32'hc1dcf4f1},
  {32'h450abb03, 32'hc30a30e1, 32'hc2e04424},
  {32'hc47a708d, 32'h44bb0106, 32'h42ad9ae4},
  {32'h4456b9b0, 32'h43805593, 32'h43e49d62},
  {32'hc51212a0, 32'h443d6012, 32'hc30de878},
  {32'h4402d473, 32'hc4ae7490, 32'h41945171},
  {32'h43b1abe6, 32'hc4aa1ce3, 32'h43e2378f},
  {32'h4433c1a6, 32'h43cf2a70, 32'hc4240d2f},
  {32'h43fc9150, 32'hc387e884, 32'h455ef325},
  {32'h438602ee, 32'hc49db46a, 32'h44846a0d},
  {32'h4523de89, 32'h42a8e08b, 32'h436e9c7b},
  {32'hc3970e53, 32'h43c35fdf, 32'h44b2eb59},
  {32'h43d24bdb, 32'h4488be8a, 32'hc45be4d0},
  {32'h44030a14, 32'hc4ce4667, 32'h44835100},
  {32'h43fe472d, 32'h4234ce25, 32'hc489abf1},
  {32'h43deb240, 32'h42d8d16b, 32'hc40b6123},
  {32'h438592b7, 32'hc522395c, 32'h44ee81df},
  {32'h44e8e4f7, 32'hc3f3aa98, 32'hc4603300},
  {32'h4427f807, 32'h43e5d833, 32'hc48fcd94},
  {32'hc30c4953, 32'hc37e4cfe, 32'h4523b66e},
  {32'h44a959f2, 32'h430df36a, 32'hc3c6dd6c},
  {32'hc3af1b65, 32'hc50da3bc, 32'hc387559b},
  {32'h441e9376, 32'h44ddc831, 32'hc119ffa9},
  {32'hc4d730fb, 32'hc44f7d20, 32'h42eddfa6},
  {32'h45580010, 32'hc3f3f400, 32'hc30f84ab},
  {32'hc5037e01, 32'h433253f9, 32'hc39f85aa},
  {32'h44da7ee1, 32'h4242fb80, 32'h4321fc68},
  {32'hc4a7e16c, 32'hc48504c9, 32'h43442d61},
  {32'h441d3327, 32'h4512572d, 32'h42ad930e},
  {32'hc47c5ce7, 32'hc417b5fb, 32'h439e4c44},
  {32'h45583f45, 32'h442ae3da, 32'hc278006e},
  {32'hc3c165d8, 32'hc51eb3aa, 32'h431ebf7c},
  {32'hc4f1f2a4, 32'h438a3404, 32'hc38181b4},
  {32'h430b378a, 32'hc45287bc, 32'h4427ab04},
  {32'hc3c12ebb, 32'hc40519df, 32'hc4968361},
  {32'hc3e09877, 32'h438ac250, 32'h4464a3e3},
  {32'hc52e5cec, 32'h43a5b316, 32'hc2a87d65},
  {32'h45114f76, 32'hbf8c0928, 32'h43dcd0d8},
  {32'hc4a50464, 32'hc482ea8e, 32'hc2978391},
  {32'h45188a9d, 32'hc2d94d61, 32'hc34066cc},
  {32'hc4a733dd, 32'hc437b24e, 32'hc4b1b4b8},
  {32'h4482507f, 32'h440c6bbe, 32'h44c76f04},
  {32'hc4bc04eb, 32'h441f4624, 32'h43a5685d},
  {32'hc41dafc7, 32'hc4918b9a, 32'h44837cfd},
  {32'h43daccf0, 32'hc451ba06, 32'hc2c01206},
  {32'h4402abbb, 32'h44f4aeec, 32'h420c5094},
  {32'hc3379c8d, 32'hc4884433, 32'hc47cc9d6},
  {32'h446a5ddd, 32'h42a389e5, 32'hc3061cd0},
  {32'h4442eca0, 32'hc3a62640, 32'hc142f875},
  {32'h441acac0, 32'h437add92, 32'h44a3686b},
  {32'hc44c8c6c, 32'hc2ba9da0, 32'hc4d413f6},
  {32'hc486b4e2, 32'h439cd5ad, 32'h43028e67},
  {32'hc50b52bc, 32'hc3955111, 32'hc325c31f},
  {32'h45313764, 32'h446dc2f6, 32'h4419f6b3},
  {32'hc4073341, 32'hc3cd57e5, 32'hc4684739},
  {32'h442ada8c, 32'h44ec6d82, 32'h441c8c26},
  {32'hc4cb6fb7, 32'hc4674f7f, 32'h432ec9f8},
  {32'hc4ab6c9c, 32'h43667e3d, 32'h441af32e},
  {32'hc54d64d5, 32'h43320475, 32'hc389fa84},
  {32'h4510ea2f, 32'h40fc1e46, 32'hc41b1712},
  {32'hc2f0c690, 32'hc43b8864, 32'hc44d901e},
  {32'hc275d0c0, 32'hc4bf2b09, 32'h45063486},
  {32'h44c100aa, 32'h43cebecc, 32'h43850489},
  {32'hc424a807, 32'h451330d5, 32'h442198ea},
  {32'hc4243b55, 32'hc27724a9, 32'hc5728ccc},
  {32'hc408552a, 32'h4439038f, 32'h43a574f0},
  {32'hc2c73c98, 32'hc4152327, 32'hc5384c06},
  {32'hc3ceb098, 32'h44180dd7, 32'h450765b8},
  {32'h453ef26c, 32'h4339f1e9, 32'h43854454},
  {32'h43fc4f14, 32'hc4711301, 32'h4523195d},
  {32'hc40aace8, 32'h446f8dc1, 32'hc51b3ae2},
  {32'hc3ff3530, 32'h44965865, 32'hc28ce9c9},
  {32'h448e681e, 32'h439853d8, 32'hc4959ef6},
  {32'hc3c6133e, 32'h44c0cebc, 32'h43a3e74d},
  {32'h428af670, 32'hc36d7a7c, 32'hc4857974},
  {32'hc2839e12, 32'h4481cb29, 32'h44ac54a7},
  {32'h42c7ea54, 32'hc439da6b, 32'hc555027d},
  {32'h44464999, 32'h4470ff11, 32'h43f3246a},
  {32'h439fc1fb, 32'hc50723b6, 32'hc392e1ca},
  {32'hc4f7f5ba, 32'h44475a8e, 32'hc36aa844},
  {32'h441d9161, 32'hc31bf04e, 32'h42db9e18},
  {32'hc486e63e, 32'h440dbe0a, 32'hc37722d5},
  {32'h45358a41, 32'hc4005746, 32'hc34fd81e},
  {32'h4433253f, 32'h442e9c56, 32'h429a06c2},
  {32'hc3e59260, 32'hc3d0529b, 32'hc3d1f9a9},
  {32'hc594f99e, 32'h435e286c, 32'hc3bc85c6},
  {32'h456ccef9, 32'h43aeaaf3, 32'hc294b17f},
  {32'hc4a41938, 32'hc341bdc9, 32'hc326bfbd},
  {32'hc5423e9c, 32'h430f34a4, 32'h43601b0c},
  {32'h43aadc7a, 32'h440804bf, 32'h451da056},
  {32'h4419730e, 32'h44b425f3, 32'h430f0cc7},
  {32'h441e19bc, 32'hc537a583, 32'hc23e3016},
  {32'hc4c91b0a, 32'h44158b46, 32'h421d3875},
  {32'h447beaa8, 32'hc363d5c4, 32'h443f3510},
  {32'hc48e6125, 32'h44afa26f, 32'h43bf31f1},
  {32'h45323a2c, 32'hc40a2dee, 32'h43087b06},
  {32'hc408793b, 32'h423f4d77, 32'hc4330f6e},
  {32'h451d44c6, 32'h430b730e, 32'hc29a30a8},
  {32'hc5042aac, 32'h4389af18, 32'h424f1436},
  {32'hc33e7710, 32'hc38b3d03, 32'hc36f5774},
  {32'hc336aa72, 32'h443f18cc, 32'h44185910},
  {32'hc3974542, 32'hc5279bbe, 32'hc39402a6},
  {32'hc3d24a84, 32'h438f5c78, 32'h44144f58},
  {32'h4327dbf4, 32'hc51e5896, 32'h42ca00f7},
  {32'hc389b9cf, 32'h450f139d, 32'h437bc6f9},
  {32'h453f3568, 32'hc2deffc5, 32'hc34028c5},
  {32'hc48b9ad8, 32'h43c00633, 32'h43fbc587},
  {32'h4499edaa, 32'h436a265f, 32'hc4902a54},
  {32'h3f28a200, 32'h44fd311a, 32'hc25fe4e8},
  {32'h44df37fe, 32'hc3854217, 32'hc3d7a818},
  {32'h43190e42, 32'h45480170, 32'h438753e2},
  {32'hc2accb96, 32'hc433a952, 32'hc41c5dcc},
  {32'hc4014815, 32'h442a7282, 32'h43e46b1f},
  {32'h434e7af2, 32'hc4f71a6a, 32'hc404a75f},
  {32'h45167d6a, 32'hc345a312, 32'h438772a0},
  {32'hc51ed47e, 32'h4346429d, 32'h43efdfae},
  {32'h44857b6a, 32'hc33223bb, 32'hc3ba0570},
  {32'hc3f54a28, 32'hc539feea, 32'hbfb159a4},
  {32'h44898d46, 32'h44664758, 32'h42811d80},
  {32'h445c9f42, 32'hc387a219, 32'hc405c2e8},
  {32'h450d87d6, 32'h44bf5994, 32'hc1bef7f1},
  {32'hc53ce69a, 32'hc3ae0ef4, 32'hc184390b},
  {32'h4492c0f9, 32'hc4191a07, 32'h4312d348},
  {32'hc4b4bf5c, 32'h43bdd178, 32'h4432cafe},
  {32'h446d6591, 32'h43df956f, 32'h42703f6c},
  {32'hc403d301, 32'h42fb0f18, 32'hc37ae24b},
  {32'h44fd5384, 32'h42e317a1, 32'h44a73e81},
  {32'hc1042368, 32'hc50f1fd4, 32'hc48e2980},
  {32'hc428a2f0, 32'h432e7bbf, 32'h439d77d1},
  {32'hc4b7adca, 32'hc49b744b, 32'h42e70268},
  {32'h4491b943, 32'h44110224, 32'hc38f71e1},
  {32'h43da3358, 32'hc33382a1, 32'hc4aa893f},
  {32'h456c4fb1, 32'hc41a238e, 32'hc187bd4a},
  {32'hc4a7028a, 32'h44262aea, 32'hc47060b3},
  {32'h451cf2ae, 32'h424f2214, 32'hc413a030},
  {32'hc5380b73, 32'h434528e6, 32'hc3a9b514},
  {32'h44c87546, 32'h43dae8aa, 32'h4313c577},
  {32'hc534edba, 32'h437efb77, 32'hc34942f0},
  {32'h4481e6b4, 32'h44b1a7fb, 32'h43c760fa},
  {32'hc4cef3b1, 32'hc43992c4, 32'hc35d01bc},
  {32'h429d8048, 32'h44b06d06, 32'hc36084ae},
  {32'h431cbd4a, 32'h44fcf96e, 32'h42456fef},
  {32'hc5216018, 32'hc40e140a, 32'h437b9670},
  {32'h44746a3c, 32'h44c319c7, 32'hc382105d},
  {32'hc4ffc41a, 32'hc1946882, 32'h428f244d},
  {32'h451ac29c, 32'h440d97ac, 32'hc40136f5},
  {32'hc4973083, 32'hc4bcc490, 32'hc38150e7},
  {32'hc444381d, 32'hc1ab9f62, 32'h4359345a},
  {32'hc5545822, 32'hc36ad77b, 32'hc37dc3ee},
  {32'h449fb094, 32'h438176a1, 32'h44389e01},
  {32'hc46f0426, 32'hc3ba9530, 32'hc2a4ba84},
  {32'h431d77a6, 32'h44b6c967, 32'h432b6058},
  {32'hc3f0c1d4, 32'hc3dc1c5a, 32'h44a1ed5d},
  {32'h44e293f2, 32'hc2f2b8ee, 32'h428ab352},
  {32'hc4f125db, 32'hc3cb5ded, 32'hc10f7edd},
  {32'hc3f6149c, 32'h43c877f6, 32'hc509f53d},
  {32'hc4a3097a, 32'hc3ee94f5, 32'hc30855ff},
  {32'hbf3b1800, 32'h44a96091, 32'h4483e582},
  {32'hc4fd34ee, 32'h423d9b8a, 32'h436c20b7},
  {32'hc414fb94, 32'h41748286, 32'hc3a44861},
  {32'hc4931ce7, 32'hc4e5e764, 32'h431afaae},
  {32'h44f0efa6, 32'h44437c5c, 32'hc41ed72b},
  {32'hc3051460, 32'hc3bb3552, 32'h448468bb},
  {32'h44813a54, 32'h43dfffd1, 32'hc4410dab},
  {32'hc42c9f56, 32'hc4cf9d3e, 32'hc3d69a65},
  {32'hc327cb90, 32'h436c6bc0, 32'hc3e7ec58},
  {32'hc525a6d0, 32'hc39823f4, 32'h41e01b34},
  {32'h436f81e0, 32'hc3e4ddf0, 32'hc547d585},
  {32'h451bc906, 32'hc1c30db3, 32'hc4106a1d},
  {32'hc3a09612, 32'h45212726, 32'hc26f0fad},
  {32'h45256e78, 32'h42d064b7, 32'h4301400f},
  {32'hc4170146, 32'h44c6be63, 32'h441e08ff},
  {32'h454601e2, 32'hc30181d2, 32'h42d5a0dd},
  {32'h444bb203, 32'h43ad0071, 32'h43b31903},
  {32'h4509b2fe, 32'h4404de98, 32'hc3a60c1e},
  {32'hc471b450, 32'h42ca25b1, 32'hc217940c},
  {32'h43da0235, 32'hc3a93005, 32'hc3ac7256},
  {32'hc45ba5c8, 32'h441e8214, 32'hc34cd6b0},
  {32'hc2948000, 32'hc4509d04, 32'h4494719b},
  {32'hc49c7a92, 32'h43bc516c, 32'hc413c434},
  {32'h44255308, 32'h43056d8f, 32'h44c62ef0},
  {32'hc45cc5c3, 32'hc3db3281, 32'hc5089395},
  {32'hc49865e7, 32'hc2d5fe4f, 32'hc38318d0},
  {32'hc4956e22, 32'hc3d75a67, 32'hc4ba1b30},
  {32'h44d7e4d8, 32'hc4868529, 32'hc32ff810},
  {32'hc424f3b4, 32'hc37d4fe2, 32'hc384036e},
  {32'h44ccb32d, 32'hc4245bac, 32'h44782464},
  {32'hc3d2c758, 32'h450e646c, 32'hc3e052bd},
  {32'hc492119b, 32'h423eb0d7, 32'h420e1fbb},
  {32'hc4fe8455, 32'h43dd7991, 32'h434ee9c0},
  {32'h43ad411e, 32'hc41df995, 32'h44b05cc7},
  {32'hc44a25bf, 32'h4409f02a, 32'hc36ad68b},
  {32'h450b4afe, 32'h43ddc8e2, 32'h442cdb92},
  {32'hc56264a5, 32'hc3c058a2, 32'hc4190089},
  {32'hc388ef08, 32'h412eef59, 32'h4413fb21},
  {32'hc3092aa2, 32'hc233cbf0, 32'hc4890afd},
  {32'h4299de24, 32'hc42cf9cf, 32'h447043c9},
  {32'h4416a8da, 32'h448bdddd, 32'hc4694b65},
  {32'hc422649f, 32'h44b1c954, 32'hc2c86fb4},
  {32'h4426bf32, 32'hc4ac9d5c, 32'h43b4c196},
  {32'hc4419b32, 32'hc40de3a4, 32'hc4d7cb6e},
  {32'h442f4236, 32'h425a204f, 32'h444efe2b},
  {32'hc3fd9bf8, 32'h444aa793, 32'hc4ac8843},
  {32'h428470c0, 32'hc49a5298, 32'h44a087b0},
  {32'h430c7804, 32'hc4f158e8, 32'h4500dba7},
  {32'hc4d5ede9, 32'hc48fe324, 32'hc4103fb8},
  {32'h44bb835b, 32'hc32aeea8, 32'h43347a11},
  {32'h44bab320, 32'h444eef38, 32'hc22bda7a},
  {32'hc48ac622, 32'h438078a8, 32'hc32a55c7},
  {32'h40f42300, 32'hc4d63286, 32'hc3ca6c63},
  {32'h439e350b, 32'h41a2edda, 32'h438dc8cf},
  {32'h43c8a484, 32'h43bb18f7, 32'h452eb6e0},
  {32'hc4d09273, 32'h41e5fc4d, 32'hc3b91385},
  {32'hc4aa5684, 32'hc4066d18, 32'hc276b998},
  {32'hc58f0541, 32'hc426405a, 32'hc3f7db2e},
  {32'h44e8128a, 32'h43b12620, 32'hc35ab203},
  {32'hc51b17e8, 32'h435d0cdc, 32'h44039fa3},
  {32'hc3906cd6, 32'hc3d58861, 32'hc23c9ff0},
  {32'hc557d131, 32'h44007e79, 32'hc3ad4a17},
  {32'h446b6d44, 32'hc3a45e6c, 32'h43ef7ae3},
  {32'hc099b000, 32'h454ebde4, 32'hc3b7609d},
  {32'h44b7b78b, 32'hc4bf4d04, 32'h434b3b67},
  {32'h432b0cac, 32'h442ec35b, 32'h44268342},
  {32'h445f9817, 32'h440d182d, 32'hc47def3b},
  {32'h43b1a075, 32'hc26e33f5, 32'h454bc09c},
  {32'hc4062b19, 32'hc3c55f9b, 32'h43c4d864},
  {32'hc33dc708, 32'h42048387, 32'hc4bb4ce5},
  {32'h43e864af, 32'h43ae8467, 32'h4444f361},
  {32'h44ce2cb6, 32'h44153df2, 32'h4294442c},
  {32'hc3ae4b50, 32'hc4e378bc, 32'h4417293c},
  {32'hc4b7dff8, 32'h42432008, 32'hc447a9ed},
  {32'hc41c3171, 32'h4467ebb1, 32'hc1ad2ae2},
  {32'hc4eeb39d, 32'h432e0e0d, 32'h431c70c9},
  {32'h445406fe, 32'h43dd58b7, 32'hc4b2e384},
  {32'h444b5cf6, 32'h44b894d7, 32'hc3d70a89},
  {32'hc444c953, 32'hc3fa0705, 32'h4467b6b4},
  {32'hc3b96bf3, 32'h43bffb35, 32'hc3c25dd4},
  {32'hc443b95a, 32'hc328ade8, 32'h44bb66e0},
  {32'h438c3a50, 32'h44fa5de0, 32'hc4109f8c},
  {32'h43de9de3, 32'hc425b7fd, 32'h435aaff8},
  {32'hc4049d09, 32'hc397f1a8, 32'h4376be23},
  {32'hc55d7012, 32'hc2908d08, 32'h42384cac},
  {32'hc43a2e79, 32'h441461c0, 32'hc2789abf},
  {32'hc466e708, 32'hc50a8bfb, 32'h4385a03f},
  {32'h44ce4bc3, 32'h4431da3d, 32'hc348fdb9},
  {32'h4397d454, 32'hc392d68a, 32'h43a3b9d4},
  {32'h444a9ab8, 32'h44dc4e91, 32'h421dffa1},
  {32'hc5367bf9, 32'hc3c78d03, 32'hc3486994},
  {32'h45578276, 32'hc44c449b, 32'hc213710a},
  {32'h43b3633d, 32'h449ede12, 32'hc3086dcb},
  {32'h4287da3c, 32'hc4a96913, 32'hc48e0fab},
  {32'h41d7abd4, 32'h44c98d5b, 32'h442d7cce},
  {32'h43875ee1, 32'hc3bacf0d, 32'hc40e55a9},
  {32'h43a605d3, 32'h4534aeb9, 32'h430de0fe},
  {32'hc408e8b6, 32'hc5002185, 32'hc3cdca3f},
  {32'hc4514787, 32'hc29df807, 32'hc2cf0048},
  {32'hc4895c81, 32'hc43c4980, 32'hc3afbb4c},
  {32'h41bdb27a, 32'h43b9527f, 32'h453f9dcd},
  {32'h436b5555, 32'hc1cc2003, 32'hc48ac09b},
  {32'hc445b154, 32'hc509249d, 32'h44ac22b3},
  {32'h43e51bd5, 32'h441d7c67, 32'hc4ddad0b},
  {32'hc37bd0aa, 32'h422f63c5, 32'h44719546},
  {32'hc52f06f4, 32'hc3e39a49, 32'h4397f41e},
  {32'h4473d86c, 32'h4507467c, 32'hc2a966ba},
  {32'hc28bf286, 32'hc49dee44, 32'hc3b8776c},
  {32'h454789ba, 32'hc3b6de2d, 32'hc3e98f3d},
  {32'hc47cbbe8, 32'hc4b871bc, 32'hc4292657},
  {32'h451a47ff, 32'hc34b412b, 32'h4368af46},
  {32'hc453d26d, 32'hc5112878, 32'hc2eb8205},
  {32'h43ef0563, 32'h450336b9, 32'h41104f70},
  {32'h44e5a11f, 32'hc025bd96, 32'h42f3cc75},
  {32'h4437f692, 32'h44f138d4, 32'h4353a18d},
  {32'hc4743a1c, 32'hc496f1a2, 32'h41a42f4e},
  {32'hc3724a86, 32'hc2f9b082, 32'h43a2936b},
  {32'hc57ac5be, 32'h436c8e44, 32'h438c1af8},
  {32'h45258eb6, 32'h435e240f, 32'h443879c1},
  {32'h44566e84, 32'hc48aa406, 32'hc40d0ef8},
  {32'hc3078518, 32'h44eff993, 32'h43d3627f},
  {32'h447e640b, 32'h4108cc9b, 32'hc23b4901},
  {32'hc4884191, 32'h4506c0eb, 32'h42af7bd7},
  {32'hc3faa569, 32'hc3d53516, 32'hc53ef62f},
  {32'hc3e28435, 32'hc311ff43, 32'h4467d0bd},
  {32'h447b45be, 32'hc4432794, 32'hc467d05a},
  {32'hc491d857, 32'h448043a3, 32'h44544412},
  {32'hc43bb84d, 32'hc392e912, 32'hc4b0b8aa},
  {32'h439e4d86, 32'hc4bd017d, 32'h44d05b67},
  {32'hc3d50559, 32'h44858a1c, 32'hc4e33041},
  {32'h43171312, 32'hc4b0b7c2, 32'h440f93c6},
  {32'h441e5c1e, 32'hc431f0e6, 32'hc44c52e8},
  {32'h42da00d6, 32'h4363d3b0, 32'h44fcdf14},
  {32'h4425a20c, 32'h42a39fe5, 32'hc3c8672e},
  {32'hc3eb8af2, 32'h44aca330, 32'h450183b9},
  {32'h447cd590, 32'hc4dc9d02, 32'hc488eca6},
  {32'h4456eb26, 32'hc3f0713f, 32'h4419dc82},
  {32'hc1dadc08, 32'hc54ed8cb, 32'hc38de0da},
  {32'hc535c53b, 32'h442428fb, 32'hc17fccd3},
  {32'h438efd0d, 32'hc0949482, 32'h438dd034},
  {32'hc3cf57d4, 32'h44b33f64, 32'hc385ccf7},
  {32'hc2dc3a74, 32'hc533870f, 32'hc3ce6964},
  {32'hc39bff38, 32'h44177100, 32'h43a963c5},
  {32'h44bf7584, 32'h43c5db34, 32'h4383e98a},
  {32'hc512a1b6, 32'hc3520d03, 32'h42e601b9},
  {32'hc326323f, 32'hc30a4a99, 32'hc3de35b0},
  {32'h438298be, 32'h436915c7, 32'h449e7160},
  {32'hc327dffe, 32'h41847799, 32'hc4f0c8b0},
  {32'h45201aed, 32'h43c0ccf3, 32'h44be2599},
  {32'hc5146c1d, 32'hc32114ce, 32'h42187bb9},
  {32'h4200fe00, 32'hc5304f7e, 32'hc382e3b3},
  {32'hc52e0fe3, 32'h43507e09, 32'hc1efef0f},
  {32'h450f3e2e, 32'h440216c6, 32'hc361fa3f},
  {32'hc52b522c, 32'h4453bfc8, 32'h4328efc6},
  {32'h439fbfc2, 32'hc4833884, 32'hc40ec721},
  {32'h44787799, 32'hc2ae75e0, 32'hc43fa0f1},
  {32'h452f6e6b, 32'h42325d5c, 32'hc286f004},
  {32'hc50e22db, 32'hc3c5c4b1, 32'h43a6de78},
  {32'h44152bf2, 32'hc3806260, 32'hc462934f},
  {32'h433e8194, 32'h43d18053, 32'h45163e66},
  {32'h44408029, 32'hc35ae955, 32'hc4e8aa83},
  {32'h42a39763, 32'h44d70cca, 32'hc2f68e10},
  {32'h4342b71a, 32'hc4f751b5, 32'h4239cfba},
  {32'h43ab700c, 32'h44d557a2, 32'h445aeb1e},
  {32'h45357ebe, 32'hc33d1f72, 32'h439b5fe0},
  {32'hc4a3ba78, 32'hc387b9c4, 32'h42de34e4},
  {32'h45087e3a, 32'h443b0c17, 32'hc48066e5},
  {32'hc4cdd49f, 32'h4348dd31, 32'hc3a9168e},
  {32'h41dfd894, 32'hc4a279c2, 32'hc44a11f8},
  {32'hc388d358, 32'hc225c38f, 32'h4518d265},
  {32'h42dec171, 32'hc4a2a4e7, 32'hc2991258},
  {32'hc3f7045d, 32'h449d44d0, 32'h439863a8},
  {32'h448ef179, 32'hc49234f1, 32'hc3f0ab00},
  {32'h4537606c, 32'h432bc451, 32'hc3e4a4d0},
  {32'hc51ce90c, 32'h42bd7590, 32'hc35b2ba9},
  {32'h43c9b5e4, 32'h4407a611, 32'h43ada6c0},
  {32'hc46cc992, 32'hc4e9ae5e, 32'hc3f4769d},
  {32'h4461830c, 32'h44a7fd3f, 32'h431ea11a},
  {32'h42409557, 32'hc515e929, 32'h438d911e},
  {32'h440429b2, 32'h450ff1a5, 32'h411c95ef},
  {32'hc49c1c84, 32'hc37b7154, 32'h43e4e2f4},
  {32'hc28a8f30, 32'h44c7e583, 32'h42da267d},
  {32'hc4e0f245, 32'h43e61e99, 32'hc47646cd},
  {32'h45110845, 32'h42fa15dd, 32'hc44b1742},
  {32'hc520a7fb, 32'h440ed023, 32'h43204bbe},
  {32'h4415d0eb, 32'h448805e6, 32'h438a77eb},
  {32'hc4b6c1fb, 32'hc4a64a86, 32'hc3da1bc6},
  {32'h4481b40a, 32'h430eacea, 32'h4406bada},
  {32'h43272177, 32'hc3822a63, 32'hc3fca41b},
  {32'h446424fa, 32'h443c6cb5, 32'h44560a64},
  {32'hc4a879ef, 32'hc487f031, 32'h43bc0e0c},
  {32'h44faac18, 32'hc3972075, 32'h4473a8eb},
  {32'hc4a538a4, 32'hc28b44f2, 32'hc351ecfe},
  {32'h45345d38, 32'h41dc8013, 32'hc43baea9},
  {32'hc1e106e0, 32'hc4fc7727, 32'hc3d8cf2d},
  {32'hc2f5e884, 32'h44f2a482, 32'h43510fbc},
  {32'hc2a057bc, 32'h4370dc4a, 32'hc4f8712f},
  {32'h446b4c06, 32'h44385a19, 32'h44c8d404},
  {32'hc4e49fcc, 32'hc42fd03e, 32'hc4a2fb95},
  {32'hc4923e41, 32'h434592df, 32'h437c51ff},
  {32'hc4b40642, 32'h44306d26, 32'h43e62262},
  {32'hc539435e, 32'hc2d7012f, 32'hbedbe180},
  {32'h43218cc4, 32'h454298e8, 32'hc3b64a2f},
  {32'hc4d4d806, 32'hc38bed76, 32'h429d5ed8},
  {32'h44e21a38, 32'h448014d6, 32'hc3ba2d92},
  {32'hc48b92fe, 32'hc49e6085, 32'hc36a8a75},
  {32'h448bdee6, 32'h43ce64e1, 32'h42970c6b},
  {32'hc4bd13da, 32'hc32d4cd6, 32'h430ebdb2},
  {32'h45000933, 32'h436f1c90, 32'hc297b637},
  {32'hc5156072, 32'h43aa904d, 32'hc39006cc},
  {32'h4439ce7e, 32'h436ce110, 32'hc29793c4},
  {32'hc4c72e8f, 32'hc3dd2245, 32'hc22e837c},
  {32'hc38fd3de, 32'h4360c8be, 32'hc380dcf2},
  {32'hc3db3d68, 32'hc4978862, 32'h4485f301},
  {32'h43b7860a, 32'h44fa3539, 32'hc34be9e0},
  {32'h441e4480, 32'hc2ddf1fc, 32'h43acd71f},
  {32'h452ecdb7, 32'h42aebb11, 32'hc277af8b},
  {32'hc493373c, 32'hc37bed03, 32'h443612b5},
  {32'hc4ec1bc1, 32'h43768c36, 32'hc2981bcc},
  {32'hc579c4ab, 32'hc4031c27, 32'hc339cddf},
  {32'h44b69db0, 32'h44d999cc, 32'hc421a6b9},
  {32'hc3cbb786, 32'hc467ea38, 32'h43e35024},
  {32'h442f8612, 32'h4381487c, 32'hc50b7478},
  {32'hc440d001, 32'hc0ebf037, 32'h4458a1aa},
  {32'h44997e87, 32'h43b3c944, 32'hc310a7c0},
  {32'hc3d1299a, 32'h4439541d, 32'h456f70ac},
  {32'hc30591d0, 32'h43b3f611, 32'hc4298276},
  {32'h44444333, 32'hc4a94e56, 32'hc42fc48b},
  {32'hc5552b53, 32'h43ba28d7, 32'h43960716},
  {32'hc3e18373, 32'hc41f8dd3, 32'hc20cf0ec},
  {32'h428bec13, 32'h444bb57c, 32'hc42692f6},
  {32'h450c9a55, 32'hc36b87f0, 32'h43c87a65},
  {32'h44584229, 32'h433c45e7, 32'hc206a434},
  {32'h454fc996, 32'h425dce20, 32'hc4028258},
  {32'hc4f4fecc, 32'hc38aeeb2, 32'h43b252fe},
  {32'h452f87a4, 32'hc3672a7c, 32'h44327353},
  {32'h4312e897, 32'hc3c63644, 32'h440c04a2},
  {32'h4439265f, 32'hc3c7f871, 32'h44cea5ec},
  {32'hc37de630, 32'h448e9529, 32'h43015e17},
  {32'h4412e81e, 32'hc1d85236, 32'h44e94c57},
  {32'hc4d35b32, 32'h43297ab0, 32'hc4a92e23},
  {32'h44408313, 32'hc3160f18, 32'h4416fb34},
  {32'h430b7414, 32'hc35e1a92, 32'hc5222682},
  {32'h4542b28d, 32'h440f9f09, 32'hc36ec111},
  {32'h44f97b0d, 32'h431f16d1, 32'h43b0332d},
  {32'h44e565d8, 32'hc495954b, 32'h42abfeb7},
  {32'hc427bc2c, 32'h44409136, 32'hc4a55d96},
  {32'h44de5ae0, 32'h43690e49, 32'h4341430f},
  {32'hc5403d9d, 32'h43961790, 32'h42ad0084},
  {32'h43cd26b5, 32'hc3301947, 32'h440c27d7},
  {32'h4389cc08, 32'h442230d2, 32'hc3ad371d},
  {32'h4567998f, 32'h4410f31f, 32'hc23cfc7c},
  {32'hc4dc7814, 32'hc2eb2c88, 32'hc45c464e},
  {32'hc37f003c, 32'hc35128f9, 32'h43d9d6e9},
  {32'hc4217cc0, 32'hc4fcdc39, 32'hc4833242},
  {32'hc3bb74a2, 32'h4432252e, 32'h44ae4583},
  {32'hc4f113ca, 32'hc37bc718, 32'h43202a58},
  {32'hc51ac980, 32'h43ba4965, 32'h4231afb0},
  {32'h43a272ef, 32'hc466a26a, 32'h447edf8e},
  {32'hc29d5452, 32'hc3bdffca, 32'hc49c5ff6},
  {32'hc3a07e40, 32'hc2364c81, 32'h43553ec9},
  {32'hc55b5567, 32'h43b203c0, 32'hc34c8aca},
  {32'h44bd14dc, 32'hc427764a, 32'h43b727b8},
  {32'h434b3de0, 32'hc3ae9c10, 32'h44ddb312},
  {32'hc30987ae, 32'h450fdc8a, 32'hc4dff500},
  {32'hc4b3b165, 32'h42873b1a, 32'h4331b85f},
  {32'hc3082ebf, 32'hc2a5dfe1, 32'h44d32305},
  {32'hc4fb5d36, 32'h4212d5b2, 32'hc481cb1b},
  {32'h4390c784, 32'hc43a1238, 32'h43933962},
  {32'hbfe99f80, 32'h429992a0, 32'hc50c15ef},
  {32'h440f133e, 32'hc49f9c57, 32'hc3890091},
  {32'hc45d6a61, 32'h448c7970, 32'h42840c68},
  {32'h44900b4e, 32'hc305bd00, 32'h414215e8},
  {32'hc4751800, 32'hc455f1ab, 32'hc3a02239},
  {32'h4551c807, 32'h437e1801, 32'h43aef33a},
  {32'hc527f282, 32'hc3517ccf, 32'hbf2df65b},
  {32'hc26ea218, 32'hc53649f9, 32'h43b68a39},
  {32'hc487cbd9, 32'h44091f0b, 32'hc33be794},
  {32'h44cdc6d5, 32'hc285a669, 32'h43d2e1f3},
  {32'hc46bc448, 32'h450c26cc, 32'hc418cf94},
  {32'h44a9d3ad, 32'hc49b94a7, 32'h4463151a},
  {32'h43a740c2, 32'hc2599bf8, 32'h44b0f9ec},
  {32'h44760a63, 32'hc2d26421, 32'hc4775466},
  {32'hc31e8bf2, 32'hc4bcabc0, 32'h44ce3876},
  {32'h42b22b5e, 32'h42ebb1ec, 32'h451ac7f4},
  {32'h44b3a46b, 32'h43caefa9, 32'h437523c6},
  {32'hc4f79305, 32'hc3b6afcd, 32'hc30f9399},
  {32'h4475af4c, 32'h42a40fc3, 32'hc4dfdd17},
  {32'hc2966c64, 32'hc55be0dc, 32'hc3e68a7a},
  {32'h44d579da, 32'hc43d0adf, 32'h43841f96},
  {32'hc2b8a4e4, 32'hc4059808, 32'hc415ef40},
  {32'h441bce8e, 32'hc4870c53, 32'h452eb993},
  {32'h444b67f3, 32'hc2ed5ca8, 32'hc48b150c},
  {32'h44eeeecb, 32'hc1e7e2cd, 32'hc395a531},
  {32'hc37b5714, 32'hc53e8f96, 32'hc41de8ba},
  {32'hc42ee9ad, 32'h42f0495f, 32'hc41f935e},
  {32'hc32e3c09, 32'hc4c2aaaf, 32'h44a58561},
  {32'hc3c26431, 32'hc388f23f, 32'hc55c48e1},
  {32'h43cad926, 32'h43aff466, 32'h44a10772},
  {32'h44c25876, 32'h436d0b6c, 32'hc3b21431},
  {32'hc55f6eb4, 32'hc321ec41, 32'h40d91f3c},
  {32'h439a26d1, 32'hc0eb8645, 32'h42e00fbe},
  {32'hc40ecb5c, 32'hc4d4101f, 32'h410c2272},
  {32'h4519b952, 32'h43e6308a, 32'hc42791c0},
  {32'hc2d25378, 32'hc33f6623, 32'h4433a38f},
  {32'h442452e9, 32'h44944225, 32'hc36eea8f},
  {32'hc528fa74, 32'hc444a5a1, 32'h43196c7f},
  {32'h44eb7548, 32'hc385458c, 32'hc3c327e0},
  {32'hc3ff4b55, 32'h441b2e54, 32'h4346d360},
  {32'hc0f9098b, 32'h440d98f4, 32'hc5103e07},
  {32'hc432e992, 32'hc4a24ebb, 32'h44f93678},
  {32'hc1e529ec, 32'h440f066a, 32'hc4fd875d},
  {32'h44300c9d, 32'h4475b9da, 32'h4243f3de},
  {32'h43babe27, 32'h42066e5c, 32'hc51fca00},
  {32'h43f7c646, 32'h43473257, 32'h43ee5ecc},
  {32'hc32e60b9, 32'hc3c45292, 32'hc5188428},
  {32'hc257ccf0, 32'h43beb4df, 32'h44d1a2cd},
  {32'hc3b4ed62, 32'hc3f30959, 32'hc1af2bb3},
  {32'hc3e5fd05, 32'hc48706fe, 32'h45166f07},
  {32'h441194fb, 32'h4435cceb, 32'hc517f65d},
  {32'h42cf5c76, 32'h442d771b, 32'h432b0cb8},
  {32'hc0d87a21, 32'hc546d60d, 32'hc328ef77},
  {32'h41d322c7, 32'h448cde02, 32'h45036d51},
  {32'h448c8cf8, 32'hc2acdf5c, 32'hc4b9c022},
  {32'hc39e36cb, 32'h4443d330, 32'h45670b21},
  {32'hc3d8add0, 32'hc4b87ff5, 32'hc47b7c6c},
  {32'h4252753b, 32'h443bd804, 32'hc31eaf3a},
  {32'hc4e615a8, 32'hc46a0d94, 32'hc3ab5967},
  {32'h4457461b, 32'h44c32f8a, 32'h438938f5},
  {32'hc334258b, 32'h43158c50, 32'hc3848bd2},
  {32'h4577fe47, 32'h4383a530, 32'h434dae49},
  {32'hc53c39b4, 32'hc3f368ed, 32'h424b162c},
  {32'h44c99fdb, 32'h440bf9ab, 32'h440b8dd1},
  {32'hc42fd600, 32'h42451502, 32'hc4177975},
  {32'hc37e1370, 32'h44052d4b, 32'h43de631e},
  {32'h44806c6c, 32'h42da10cb, 32'hc3c56696},
  {32'h445911ea, 32'hc49c974e, 32'h450185a3},
  {32'h4497cf6b, 32'h442a966c, 32'h439075e3},
  {32'hc451c99a, 32'h44245d60, 32'h4419cdbf},
  {32'h455d864c, 32'hc1cb578e, 32'hc3bfc5c2},
  {32'hc2b13db0, 32'h44c4e20d, 32'h441a4b5d},
  {32'h433ef0a0, 32'hc4ab3cca, 32'hc4cf6751},
  {32'hc5125337, 32'hc3da304e, 32'h4463c586},
  {32'hc3aa33f9, 32'hc47488bd, 32'hc3639b21},
  {32'h43873fea, 32'h451154fd, 32'h43cf1fa9},
  {32'h44bafa7c, 32'hc38020c4, 32'hc39d22d0},
  {32'h4400c4f6, 32'h44c20971, 32'h43bfea48},
  {32'hc2ccfafc, 32'hc2a2f3fe, 32'hc53cc67e},
  {32'hc44cf076, 32'h43abf528, 32'h4502c096},
  {32'h44a3cc1e, 32'h42df8c63, 32'h42a2d53c},
  {32'hc4156cd2, 32'hc2b1802d, 32'h450d1297},
  {32'h452b5ec0, 32'hc3970f86, 32'hc32415b3},
  {32'h42a2367e, 32'h44d6f1d3, 32'h442364ef},
  {32'h457b18cc, 32'hc4098752, 32'hc38dbe83},
  {32'hc49190e6, 32'h4503cc4d, 32'hc2e8cd74},
  {32'hc4b72f68, 32'h43685d8e, 32'h433c5468},
  {32'hc50ad826, 32'h4466da2f, 32'hc389b98d},
  {32'h4450609f, 32'hc53eae9a, 32'hc38fd332},
  {32'hc545f120, 32'hc34b2d42, 32'hc233eec6},
  {32'h45474441, 32'h43c3f07a, 32'h43c2fc23},
  {32'hc5207721, 32'h440e0670, 32'hc29f0fab},
  {32'h44650076, 32'h438c9bdb, 32'hc3b6d938},
  {32'h442ad110, 32'h43095901, 32'h4168943f},
  {32'hc53fc97c, 32'h431b338c, 32'h4293e99f},
  {32'h43f6ec26, 32'h4408b4dd, 32'h452f9dbd},
  {32'hc4619c4d, 32'h4339a858, 32'hc3de3511},
  {32'h4560e482, 32'hc355e62b, 32'hc3e6318d},
  {32'hc4989b70, 32'h448d404e, 32'h43eb239c},
  {32'hc4cb0929, 32'hc2ebb3b2, 32'h43205373},
  {32'hc50b2354, 32'h44388ddd, 32'h43bd3e53},
  {32'h42540555, 32'hc53ad612, 32'hc32a8ccd},
  {32'hc40c03d0, 32'h431db831, 32'hc3ef35ef},
  {32'h42995740, 32'hc3c481ec, 32'h4476ddbf},
  {32'hc4de9476, 32'hc3cadc30, 32'h43850ebf},
  {32'h450f7313, 32'h41ee1318, 32'hc315b907},
  {32'h42b8c599, 32'h4485375a, 32'h440ae24e},
  {32'h440311d2, 32'h4238baa0, 32'hc3b17cc3},
  {32'h44b13710, 32'h43080b55, 32'h424ff5f4},
  {32'hc3427d34, 32'hc50b4df0, 32'hc30a076f},
  {32'hc31c6d68, 32'h4403f776, 32'h44a6eb82},
  {32'h450b4cad, 32'hc43f1bc9, 32'h429af7fe},
  {32'hc57a6afa, 32'h436f1aac, 32'h43b8b9c3},
  {32'h44baf6b2, 32'h43c50060, 32'hc4611ecf},
  {32'h43d7d923, 32'h44178bba, 32'h43aebf18},
  {32'h43ec6248, 32'hc403eb4c, 32'hc4c51ba4},
  {32'hc464a69d, 32'h44978d02, 32'h4444a9dc},
  {32'h45306d0c, 32'hc3b03358, 32'hc3148421},
  {32'hc1cc6c00, 32'h4487bc5a, 32'h44e5f824},
  {32'hc2601532, 32'hc54b0689, 32'hc2e952d7},
  {32'h44768ecc, 32'h43eeff95, 32'hc511fd18},
  {32'hc373fb78, 32'hc39a5385, 32'h454250dc},
  {32'hc2b3b65f, 32'h43984c0f, 32'h429205ed},
  {32'hc52219bc, 32'hc3150435, 32'h430fbe2a},
  {32'h4433d564, 32'h4498c528, 32'h438ccbd0},
  {32'hc36efb5c, 32'hc465f187, 32'hc391d96f},
  {32'h43fd0134, 32'h452c0673, 32'hc29c8c8d},
  {32'hc558985b, 32'hc467731f, 32'h44336369},
  {32'h441b019c, 32'h450ebb40, 32'hc24b74de},
  {32'hc4a3364f, 32'h439a8cb9, 32'h443ec38c},
  {32'h44b130ea, 32'h42fbf438, 32'hbf319ec8},
  {32'hc4ddb21a, 32'h42fe4746, 32'hc3341925},
  {32'h4430b707, 32'h4533fa1b, 32'h43bd2ef8},
  {32'hc460b0a2, 32'hc4ac7656, 32'hc3225e33},
  {32'h440d07c3, 32'h437f26d7, 32'h44919b1f},
  {32'hc2a14748, 32'hc512240b, 32'hc3c5d6cd},
  {32'h447890aa, 32'h448bc965, 32'h4492a44e},
  {32'hc5404f40, 32'hc3e28bdb, 32'hc36cc3ba},
  {32'h451c9261, 32'hc3f59857, 32'h42a641e3},
  {32'hc4813b0f, 32'h43cfeaaa, 32'hc4362602},
  {32'hc3a2575e, 32'h42206ee9, 32'hc2d5cd86},
  {32'hc441b4bc, 32'hc40413ec, 32'hc3e01eed},
  {32'h4483dd32, 32'h42fe785e, 32'h43b0134f},
  {32'h44674f8e, 32'hc4808c4d, 32'hc28b8c1b},
  {32'h43e0ec50, 32'h44ad533c, 32'h43aad75a},
  {32'hc4cba7c0, 32'hc4a9e256, 32'hc43c5264},
  {32'h4529ca7c, 32'hc2de281c, 32'hc381545d},
  {32'h44bc52c3, 32'hc38db1fc, 32'hc287c223},
  {32'hc4c94338, 32'hc42f5a41, 32'hc21b6c84},
  {32'h4417a870, 32'h4425527a, 32'h43c0a31c},
  {32'hc4be46c0, 32'h4437eace, 32'hc372f4fa},
  {32'h415a5900, 32'h44b6c3a6, 32'h440f7ba2},
  {32'hc4c32af2, 32'hc4816e23, 32'h42be3276},
  {32'hc413b9a0, 32'h43ae6c70, 32'h42ef3ef7},
  {32'hc574bffe, 32'hc39a3763, 32'h43609801},
  {32'h455cbf5d, 32'h4400c89d, 32'h4444a029},
  {32'h4296df14, 32'h4369d6fa, 32'h4120cdda},
  {32'h4511b1d2, 32'h42ce6362, 32'hc1a0e991},
  {32'hc45d65e7, 32'hc494d42c, 32'h43943840},
  {32'h42171688, 32'h4444ba6a, 32'h43403060},
  {32'hc341b469, 32'hc4bf776d, 32'h41be99b3},
  {32'h44178be4, 32'hc2884a0f, 32'hc4bb7144},
  {32'hc3bbf98f, 32'hc3a52a83, 32'h43759a6d},
  {32'h441d0663, 32'h4426381e, 32'hc311d66c},
  {32'hc403eecc, 32'hc39a7310, 32'h44a69940},
  {32'h4520d4aa, 32'hc3b48a14, 32'h3f90d9fa},
  {32'hc46a8d4c, 32'hc41b7065, 32'h441f0747},
  {32'h430c45b9, 32'h45284f36, 32'hc3ee6157},
  {32'h42d5ed24, 32'h42edeeda, 32'h4443aed0},
  {32'h451d4419, 32'h44122ac5, 32'hc39c31b3},
  {32'hc54504df, 32'hc0ca7eb3, 32'h43541fb5},
  {32'h4362b3cc, 32'h43a04164, 32'hc42fd374},
  {32'hc4c70558, 32'h43e9fe3d, 32'h4474e60d},
  {32'h43a3e630, 32'hc41f62b4, 32'hc42f34e6},
  {32'h4405f274, 32'hc5197541, 32'h41be1ac2},
  {32'hc51969fd, 32'h430c5817, 32'h440d6f4b},
  {32'h447a3649, 32'h441b6ff3, 32'h43819f34},
  {32'hc4cfd49a, 32'h44a02274, 32'h4421c60a},
  {32'h434e9c6e, 32'hc5182d56, 32'hc236edeb},
  {32'hc5171c5a, 32'hc23e2e33, 32'h43620de2},
  {32'h4565dd22, 32'h41eef57c, 32'hc3cc609f},
  {32'hc4c06776, 32'h43264759, 32'h439e3696},
  {32'hc3fe2c21, 32'h432b3c94, 32'h44096c9d},
  {32'hc38d82d4, 32'h44ef9cde, 32'hc2041720},
  {32'hc2e16c1e, 32'hc46072f6, 32'h44c6747a},
  {32'hc4abb13a, 32'h43bc6496, 32'h42d76877},
  {32'h429e5c78, 32'h43eb8a22, 32'h45163b0c},
  {32'hc44fe05a, 32'h451d6ca0, 32'hc3a2e6d0},
  {32'hc19bca0c, 32'hc2b9e9a7, 32'h44942dfd},
  {32'hc45bc0ec, 32'hc2d3fcd8, 32'h42a51fac},
  {32'h42d0d4c4, 32'h441cbf09, 32'h450f5480},
  {32'hc523b957, 32'h43c17c52, 32'hc158c4cc},
  {32'h43155e48, 32'hc4acf653, 32'h44d05203},
  {32'hc50c55d8, 32'h44508330, 32'hc42207e4},
  {32'h44b733e4, 32'h42367994, 32'hc335c5fd},
  {32'hc44703e0, 32'h419993ed, 32'hc4d16c30},
  {32'h4527dc20, 32'hc3ac518a, 32'hc1f1960e},
  {32'h443a3c1b, 32'h44736417, 32'hc3aaaaeb},
  {32'h442faf3a, 32'h432ceb22, 32'h4433620a},
  {32'hc46ef082, 32'hc39f8ea3, 32'hc5370f33},
  {32'h45454369, 32'hc17a7f58, 32'hc3362641},
  {32'hc2c61288, 32'h4455e815, 32'hc4f451f2},
  {32'hc2d12778, 32'h44b7417a, 32'h44ae5e39},
  {32'h44d5ba67, 32'hc3e2568c, 32'hc32c9f91},
  {32'hc5155bed, 32'h43ec829d, 32'h434f1077},
  {32'h4423c45c, 32'hc49d9b23, 32'h4353114c},
  {32'hc48a156e, 32'h43d3abbf, 32'hc3c0d264},
  {32'hc33f4ff8, 32'hc2ec32c4, 32'hc1842852},
  {32'hc4476050, 32'h44f7efe9, 32'hc45f45cf},
  {32'h43802f52, 32'hc452f251, 32'h43ee86da},
  {32'hc34797fc, 32'h44890b06, 32'h44eb0a71},
  {32'h430e7798, 32'hc482a27b, 32'hc4f29ab2},
  {32'hc3a869cf, 32'h43b65054, 32'h44df6c7f},
  {32'h42534d80, 32'hc3ca6f0c, 32'h44a0d747},
  {32'hc2fbd628, 32'h447324af, 32'hc42a03c3},
  {32'hc3d7f8a8, 32'hc2d61a53, 32'h45673eda},
  {32'h44b5e6cb, 32'hc2305094, 32'hc4639e30},
  {32'h4390be13, 32'h43a340c3, 32'h44e55dc3},
  {32'h41d730c8, 32'h42cd7622, 32'hc501bde5},
  {32'h457427a0, 32'hc3b43aa4, 32'h43f6574f},
  {32'hc539be3b, 32'h43cf1627, 32'hc4377a97},
  {32'hc3fc620b, 32'hc306c89f, 32'hc3e1e05b},
  {32'h44f88048, 32'h438638e5, 32'hc2448de6},
  {32'h44bc207e, 32'hc44dafab, 32'hc3a4f64d},
  {32'hc4738064, 32'h4478fc05, 32'hc35ee650},
  {32'h44aefb3c, 32'h43414772, 32'h43478b96},
  {32'hc4922fa0, 32'h451395dc, 32'h43a4e680},
  {32'h43e385ee, 32'hc4bd0765, 32'hc2cb34e9},
  {32'h44de6e01, 32'hc3e84a46, 32'h413c9c00},
  {32'hc43ed57c, 32'h4480600e, 32'hc51e5b34},
  {32'hc3d699e1, 32'hc3547b1a, 32'h44e267fb},
  {32'hc3e696e4, 32'hc49f0c31, 32'h439d8a34},
  {32'h436f0218, 32'h44e7fb51, 32'hc32df4ee},
  {32'hc41dbbd5, 32'hc39d6bff, 32'h4407e1d3},
  {32'h4526c023, 32'h446b6d87, 32'hc3a17828},
  {32'hc443b02e, 32'hc49d51fd, 32'h441a5a4a},
  {32'h44da9770, 32'hc303b2ce, 32'h4425cc40},
  {32'h44037a3c, 32'hc494f111, 32'hc34ef46b},
  {32'hc48ca9c2, 32'h44cb8f93, 32'h44ba7fc0},
  {32'hc33387da, 32'h44b0abca, 32'hc4d38d97},
  {32'h441ba4f8, 32'h43e04dc5, 32'hc4910838},
  {32'hc504c4db, 32'hc410c0bb, 32'h435ad707},
  {32'h450eecf0, 32'h437fe1c4, 32'hc24f5d90},
  {32'hc4b428ca, 32'hc4342964, 32'h443947a9},
  {32'hc32f9c20, 32'h4511294b, 32'hc38c1130},
  {32'h44f4e04a, 32'h40c8f154, 32'h43f6914d},
  {32'h440cbb34, 32'h439a2320, 32'hc40becc1},
  {32'hc59b8563, 32'hbff94150, 32'hc39fb1e9},
  {32'hc4def8b2, 32'hc242c048, 32'hc3979b05},
  {32'h42cb7bc2, 32'hc53ce9ec, 32'h43c10b90},
  {32'h449cec93, 32'h4395ec79, 32'hc34e7830},
  {32'h438454cc, 32'hc4be6274, 32'hc3f78cac},
  {32'hc139ed80, 32'h455178f1, 32'hc28d47a6},
  {32'hc450695c, 32'hc4ebdda6, 32'h43ab06be},
  {32'hc2c1615e, 32'h435cfecb, 32'hc3d0d438},
  {32'h43a546cb, 32'h43ac5172, 32'h44b42e81},
  {32'h45033ebf, 32'h442ce5d8, 32'hc37dae20},
  {32'hc318ccce, 32'hc44b0044, 32'h4485ae7a},
  {32'hc48eeec9, 32'hc3b03dff, 32'hc30eefd8},
  {32'h43f79685, 32'h44db9705, 32'h43cfc253},
  {32'hc44e89c6, 32'hc47f2980, 32'hc379ad3f},
  {32'h44059c82, 32'hc3cc4e0d, 32'h4493fa2e},
  {32'hc4084f20, 32'hc48de205, 32'hc49ba286},
  {32'h43df3ea0, 32'h4461c257, 32'h4524a04d},
  {32'h440e9d0a, 32'hc40fd8aa, 32'h43541b05},
  {32'hc481c809, 32'hc4f40a7d, 32'h44c920c0},
  {32'hc4aced25, 32'h4394ce9f, 32'hc4418900},
  {32'hc3cf0611, 32'h434ea833, 32'h4483f29b},
  {32'hc3969800, 32'hc45ef221, 32'hc3e25161},
  {32'h4400ca84, 32'h4377b0c1, 32'h44802fb7},
  {32'h4432a218, 32'hc3c10580, 32'h437f08b3},
  {32'hc2c7ae38, 32'h43b00630, 32'h4527c689},
  {32'hc527108e, 32'hc2767184, 32'h431bc44d},
  {32'h44073bf7, 32'h44ba7099, 32'h42f0d586},
  {32'hc522fa59, 32'hc448a55d, 32'hc3113456},
  {32'h442a04ae, 32'h4512b6fa, 32'h4219677f},
  {32'hc2e25c7e, 32'hc4a665a1, 32'hc3fb65ff},
  {32'h42fb5e1f, 32'h43e669ac, 32'h439dc18e},
  {32'hc3e6a29e, 32'hc52dd637, 32'hc3aae5a8},
  {32'h442b6b16, 32'h439fdb47, 32'h4403591e},
  {32'hc51d9cae, 32'hc3e2eb45, 32'h422d8731},
  {32'h439a8195, 32'hc41c1cb5, 32'h44005926},
  {32'h43488098, 32'hc4461c1b, 32'hc3ea2590},
  {32'hc30009dc, 32'h446e26e1, 32'h449528dc},
  {32'hc4061a1e, 32'h4433d93a, 32'hc4492d9e},
  {32'hc4811cd6, 32'h43b3e217, 32'h44740155},
  {32'h45179840, 32'hc337686d, 32'hc3292a56},
  {32'hc302a316, 32'h4508247a, 32'h433105c8},
  {32'hc291ee04, 32'hc41dd5d6, 32'hc5387c10},
  {32'hc4f32a6f, 32'h44934e7c, 32'h439d8d7a},
  {32'hc3b0e5aa, 32'hc468e603, 32'h42803f3b},
  {32'hc0376bd0, 32'h44097bf0, 32'h4482fcd5},
  {32'h44110931, 32'h4442484e, 32'hc44d14b0},
  {32'hc3a32130, 32'h43f1fc69, 32'hc1cda28b},
  {32'h436354d0, 32'hc10fc28c, 32'hc4763a9b},
  {32'hc45c6c26, 32'h426bbb19, 32'h44ab0bba},
  {32'hc3db8418, 32'hc407c30a, 32'hc2f7f80f},
  {32'h433923d2, 32'h44b887f1, 32'h44c703fc},
  {32'hc4760450, 32'hc426b07e, 32'hc5322474},
  {32'hc5235349, 32'hc3ba88c1, 32'h43aeed2a},
  {32'h44eb5a36, 32'hc48957f8, 32'h42c960e1},
  {32'hc4b4559f, 32'h449d63ca, 32'h440911ef},
  {32'h44341a70, 32'hc48b843a, 32'hc2508e08},
  {32'hc4668a6c, 32'h4484e715, 32'hc4053f0c},
  {32'h44f7e00a, 32'hc4830e2b, 32'hc3a48b19},
  {32'h438f891c, 32'h44d25b68, 32'h4317a91b},
  {32'h452f712e, 32'h43db5f05, 32'h43dede7a},
  {32'hc501eb66, 32'hc3a07639, 32'h435425f9},
  {32'hc49a8184, 32'h43454299, 32'h4306869e},
  {32'hc4cce798, 32'h43e269a2, 32'hc2f220b1},
  {32'hc4a86a0a, 32'hc32389c6, 32'hc46c9ed9},
  {32'h43f6aa80, 32'hc3e3bb56, 32'h44b243df},
  {32'hc31e77dd, 32'h43ead966, 32'h431681d3},
  {32'h449f3538, 32'h44060ca6, 32'hc1882812},
  {32'hc3d2c88d, 32'h433665cc, 32'h441a3c85},
  {32'h443d609f, 32'hc3331f7e, 32'hc34537cb},
  {32'hc4eba073, 32'h4487e91c, 32'h3df14685},
  {32'h4404325e, 32'hc504e43f, 32'hc1360d48},
  {32'hc45c6f4d, 32'hc38d47eb, 32'hc47df1c2},
  {32'h45193fe3, 32'hc2d3c864, 32'h43d47d1e},
  {32'hc3e9ba65, 32'h4428ba22, 32'h44258156},
  {32'hc48eb1c5, 32'hc3a734c8, 32'h42e7aa8e},
  {32'hc42228c5, 32'h41be7342, 32'h44b07cc6},
  {32'h4528fbea, 32'h434b13bc, 32'h419392fc},
  {32'h441ec2cc, 32'h439711c3, 32'h44069d97},
  {32'hc3ed7c98, 32'hc2448f24, 32'hc4fc3dee},
  {32'hc4226f38, 32'h44b444b4, 32'hc3397d25},
  {32'h44bed943, 32'hc404418b, 32'hc25b0fcc},
  {32'hc566c289, 32'h436fdf4c, 32'h42c0d741},
  {32'h442f83cc, 32'hc486930b, 32'hc4d830fc},
  {32'hc525e9c2, 32'h44093e27, 32'hc42e57ba},
  {32'hc322b90e, 32'hc564a0fd, 32'h4380c5dc},
  {32'hc231ce25, 32'h4532c630, 32'hc2152adb},
  {32'hc4234204, 32'h434e36fd, 32'hc3d1b6d3},
  {32'hc4a11a2c, 32'h448a0626, 32'hc3906dc3},
  {32'h453c337f, 32'hc467314d, 32'hc4793968},
  {32'hc40b5d17, 32'hc3bfbb16, 32'h431b6721},
  {32'hc4d9529a, 32'h42a97ea2, 32'h4424e01e},
  {32'h433e7b06, 32'hc41bc906, 32'hc488f7e4},
  {32'hc4743f5a, 32'hc402bcf0, 32'hc3420b90},
  {32'h453aaa6c, 32'hc3cc5386, 32'h434f9485},
  {32'h44880785, 32'h42333398, 32'h40b41b2b},
  {32'hc33b1fd8, 32'h450ada42, 32'h43914387},
  {32'hc515f3c1, 32'hc4995d24, 32'hc30e76ae},
  {32'hc48bfbdb, 32'h43e043d3, 32'h430b71fa},
  {32'hc4fcecfb, 32'hc35ae47d, 32'h42238ee1},
  {32'h45218724, 32'h4346a6e2, 32'hc3328804},
  {32'hc3897b9e, 32'hc18a6abc, 32'h44a347f0},
  {32'h44c08deb, 32'hc1117ae0, 32'h445d26b9},
  {32'hc4b244f6, 32'hc463e63a, 32'hc347863a},
  {32'h44fca858, 32'h413df069, 32'hc3a9f26f},
  {32'hc48e2556, 32'hc3ec8c0a, 32'hc3ca732d},
  {32'h4440f9a4, 32'h44944d4d, 32'h4428a691},
  {32'h438c66f7, 32'hc2ebf792, 32'hc4aadf49},
  {32'h42837000, 32'h4425c7cc, 32'h449e9921},
  {32'hc4b87510, 32'hc2c50405, 32'hc4100025},
  {32'h433b9aae, 32'h43ac7db8, 32'hc31635f7},
  {32'hc381e1a0, 32'hc4896248, 32'hc4937b1b},
  {32'h4322bcac, 32'h45559740, 32'h42a868e6},
  {32'hc4fd5bc7, 32'h42836972, 32'hc1d468c8},
  {32'hc3353b78, 32'h4502326a, 32'h43a2e19e},
  {32'hc4c5c27d, 32'hc3a1549b, 32'hc4d42a8a},
  {32'h43b2f560, 32'h438d05c7, 32'h43e3b441},
  {32'hc481aba4, 32'h44a511e3, 32'h43d3fe2d},
  {32'hc41802bd, 32'hc487b945, 32'hc2ad32d4},
  {32'h43d44109, 32'h452b7dfd, 32'hc3869c66},
  {32'hc50cfdc4, 32'hc32b88ee, 32'hc1ff39aa},
  {32'h44844efe, 32'h44a7e63d, 32'hc3b8e147},
  {32'hc47998b7, 32'hc495ea03, 32'h42c4a738},
  {32'hc4e342e1, 32'hc23e55ea, 32'hc2a1f8f1},
  {32'hc51c45c2, 32'h4322dbc6, 32'h4189d1a4},
  {32'h451f31fe, 32'h4395e3c0, 32'h442c78fa},
  {32'hc32b1d0c, 32'hc4c58ae2, 32'hc3f1a77f},
  {32'h442ed46d, 32'h44304ee3, 32'hc44956e9},
  {32'hc455a3c4, 32'hc3af0758, 32'h440e3fc2},
  {32'h445afc9b, 32'h42c7c80f, 32'hc2d1dc9f},
  {32'hc495462b, 32'hc44415eb, 32'h42a99089},
  {32'h44f4be2e, 32'hc2d5adf6, 32'hc422deec},
  {32'hc4fe2c4e, 32'hc3b0c770, 32'hc397ee4e},
  {32'h44a2a667, 32'h440aaf1e, 32'hc3d91371},
  {32'hc36876a0, 32'h43c896b6, 32'h45479b3c},
  {32'hc463cda0, 32'h44422345, 32'hc2f81de3},
  {32'hc47d14a6, 32'hc47e549b, 32'h443e9cfb},
  {32'h44a13c4b, 32'h44d5c6d2, 32'hc324d60f},
  {32'hc47a2928, 32'hc31ab505, 32'h4249fd06},
  {32'hc23e61dc, 32'h4029b08d, 32'hc531eb16},
  {32'h4208ffd0, 32'hc3f126a8, 32'h44c081e5},
  {32'h44adf034, 32'hc330ceb2, 32'hc115aa0b},
  {32'hc4a27e78, 32'hc374eaf1, 32'h4481ab25},
  {32'hc1834500, 32'hc31034eb, 32'hc4ed10d8},
  {32'h446f1cf8, 32'hc3df5d07, 32'hc482a90a},
  {32'hc48a0bc0, 32'h44f89741, 32'h439092b9},
  {32'hc3a8655e, 32'hc3534caa, 32'h440761bf},
  {32'hc551758e, 32'h43efe4db, 32'h435c695d},
  {32'h449bfb38, 32'hc4691b1b, 32'h435c8e6e},
  {32'hc41c50b6, 32'h42f8b6fb, 32'h431f51ad},
  {32'h4485d826, 32'hc44bf6bf, 32'hc4560716},
  {32'hc590451c, 32'hc35f181b, 32'hc3ad1cb6},
  {32'hc0928f00, 32'hc1d16937, 32'hc288ba2a},
  {32'h41e69740, 32'h4446a456, 32'hc4d8b038},
  {32'hc42aa0b7, 32'hc4cc240b, 32'hc4102ea3},
  {32'hc46b94bb, 32'hc30b611a, 32'h428d3f0c},
  {32'h43b26806, 32'hc3071cb9, 32'h44ab6ede},
  {32'hc4b0a624, 32'h44211e26, 32'hc3da7cc5},
  {32'h44d0ddfc, 32'h433a4394, 32'h41bd5847},
  {32'hc4f7bd36, 32'h42991520, 32'h425f076d},
  {32'h44bd7a4c, 32'h438bda85, 32'h44976d52},
  {32'h40a4fe80, 32'hc39f3865, 32'hc4f99dd1},
  {32'h44bde29a, 32'hc4635e50, 32'h43b17384},
  {32'hc3cdf124, 32'h44f008ee, 32'hc44bb22f},
  {32'hc4b327b8, 32'hc36d8e00, 32'h42602c10},
  {32'hc50f1d98, 32'h43fa8a35, 32'h43795e61},
  {32'h431951a6, 32'hc219c320, 32'h450122cb},
  {32'hc4489d50, 32'h434ca92c, 32'hc3e5a1dc},
  {32'h42dd7cc0, 32'hc318aece, 32'h443317a7},
  {32'hc548c9aa, 32'hc3deae14, 32'hc3612516},
  {32'hc4aae397, 32'hc2d2b043, 32'h431d1832},
  {32'hc4c86ea8, 32'hc41e8b34, 32'hc44aa963},
  {32'h4455e6d8, 32'h443b5b7c, 32'h443b3fa1},
  {32'hc44476ad, 32'h43d4657e, 32'hc3a8ef43},
  {32'hc41111fb, 32'h448b7f07, 32'h42f9ba2f},
  {32'h444a86ed, 32'hc33b1b5d, 32'h43ad8741},
  {32'hc3c5e8f7, 32'hc3028572, 32'hc4419b9a},
  {32'hc3cde3c1, 32'hc384ae30, 32'h42b6f9c6},
  {32'hc531ff98, 32'h42bdd8d1, 32'hc3f090ce},
  {32'h430670f0, 32'hc3eaaf6f, 32'h44693661},
  {32'h43a2cba1, 32'h449de2ac, 32'h449a5cc3},
  {32'h4281369c, 32'h44359fe4, 32'hc526befa},
  {32'h43a56cfe, 32'hc4087cae, 32'h4399ae4a},
  {32'hc19fd9d8, 32'h434274f2, 32'hc37a1b65},
  {32'hc37b4bc6, 32'h43fc39ef, 32'hc4d591ee},
  {32'h436acf50, 32'hc4806f70, 32'hc3b2b603},
  {32'h4467cae1, 32'h43f0e2c7, 32'hc411b414},
  {32'h429be042, 32'hc1f3f8ad, 32'h44fac93d},
  {32'hc4c3dfb2, 32'h43b3ed59, 32'h42195371},
  {32'hc49b2295, 32'hc2a883c1, 32'h430d184e},
  {32'hc3d224ec, 32'h443a2682, 32'hc38f3a7f},
  {32'h43af1961, 32'h443708ff, 32'h442d76c1},
  {32'hc4c3205d, 32'hc304d902, 32'h433fa136},
  {32'h4529ac97, 32'hc3be9b70, 32'h43f1ba4d},
  {32'hc5245a62, 32'h43bc1861, 32'hc28930ee},
  {32'hc33424d6, 32'hc47dfec4, 32'hc3aead24},
  {32'hc50ca67e, 32'h44a289cd, 32'hc3b165ff},
  {32'h453a2d62, 32'hc479b1b9, 32'hc28da818},
  {32'h446f832d, 32'hc331f47f, 32'h441e2cd9},
  {32'h44ad100c, 32'h4237db7a, 32'hc40385ab},
  {32'h4361a22c, 32'h445e9e80, 32'h452b4cbd},
  {32'h43f64c25, 32'hc4086ab2, 32'h44f09699},
  {32'hc3d9669f, 32'hc3ecc813, 32'hc52df6a1},
  {32'hc512775e, 32'hc3c3db24, 32'hc335212a},
  {32'hc3af30f8, 32'hc186a17c, 32'hc54e75d9},
  {32'hc5002c03, 32'hc4327680, 32'h42a73300},
  {32'h45086fbb, 32'h43339f13, 32'h440ea3de},
  {32'hc2028c2c, 32'h448f4e5b, 32'hc3d30e85},
  {32'hc53c2b43, 32'hc199daa9, 32'h43288bd0},
  {32'h4522041a, 32'hc40a1c63, 32'hc47b053c},
  {32'h4513cb2b, 32'hc2f7a04b, 32'hc38d2863},
  {32'h428d39a7, 32'hc43ff183, 32'h44d3933c},
  {32'h440a27cf, 32'h41f280d0, 32'h434a1cf2},
  {32'hc441bbe8, 32'hc50236e5, 32'hc22bd292},
  {32'h43d69a24, 32'h43dc9e2b, 32'hc4abc3ca},
  {32'h44cb4d4f, 32'hc3eac697, 32'h43953296},
  {32'h44860a8a, 32'hc44ba62a, 32'hc275def3},
  {32'hc3aeb200, 32'h44331d8d, 32'h4328d3f0},
  {32'h4388213d, 32'h43bb06e1, 32'h421927db},
  {32'hc437ad20, 32'hc49057e2, 32'h42a183e8},
  {32'h43356796, 32'h44c47223, 32'hc35eeddf},
  {32'h420a4d88, 32'hc4e50623, 32'h4112c241},
  {32'h44d899e1, 32'h449574dd, 32'h43867eb9},
  {32'hc4e364bb, 32'hc48aeae9, 32'hc39b60c5},
  {32'hc101c190, 32'h440ea726, 32'hc3cf1981},
  {32'hc3119982, 32'h4256c2be, 32'hc3583d4c},
  {32'hc37e1be4, 32'hc4dc87f0, 32'hc4168d07},
  {32'h449297b7, 32'hc32b9d67, 32'h443fc465},
  {32'h44921a3f, 32'h4359da7b, 32'hc42a6e0d},
  {32'h43dc0a51, 32'h43c35c25, 32'h44cf4e2a},
  {32'hc492b880, 32'h42c4f210, 32'hc34d95df},
  {32'h42e19515, 32'h441f2581, 32'h44d3fdcb},
  {32'hc4c3f28a, 32'h434493fe, 32'hc4629143},
  {32'h43643ae0, 32'h44182454, 32'h4529a208},
  {32'h43c8083e, 32'h44b169d6, 32'hc3b6ada3},
  {32'hc46e9067, 32'hc48dfd90, 32'h44fd6fa4},
  {32'h42988a9a, 32'hc53549cf, 32'hc3da4fb1},
  {32'hc460a96e, 32'h43c89446, 32'h4437dc12},
  {32'hc4c8b2b8, 32'hc3e10364, 32'hc3ec2013},
  {32'h440ab29a, 32'h43c4b16a, 32'h452ea39d},
  {32'hc485894e, 32'h4301eb27, 32'h43248771},
  {32'h43fa5a78, 32'h44a8e5ed, 32'h446022d7},
  {32'hc4c4420b, 32'hc3da73b6, 32'hc423156f},
  {32'hc4ba22be, 32'h43ba1219, 32'h4399f5ff},
  {32'hc52be465, 32'hc48d97de, 32'hc3cb8a0c},
  {32'h444f1d8c, 32'h44a1dfe8, 32'h42643c6c},
  {32'hc3634c02, 32'hc4d35677, 32'h43cad436},
  {32'h440d4a50, 32'h4458e50d, 32'hc4270b50},
  {32'hc2b487c0, 32'hc4d9105e, 32'hc367e464},
  {32'h45465046, 32'hc2567131, 32'h4376de59},
  {32'hc48e2359, 32'h43326412, 32'h43225f96},
  {32'h42a0dde1, 32'hc4574767, 32'hc3090654},
  {32'h43f3d2f3, 32'hc52244c0, 32'hc43b818c},
  {32'h434605b8, 32'h44edeec7, 32'h43fe01eb},
  {32'h42f19a86, 32'hc4aca60c, 32'hc391f101},
  {32'h4364db23, 32'h43bec36a, 32'h44b0970f},
  {32'h426aca40, 32'hc5062b37, 32'hc21db1ce},
  {32'hc39a06bc, 32'h441bdc58, 32'h44038801},
  {32'h44b64c2d, 32'h416558d2, 32'hc4270b5f},
  {32'hc403ccfc, 32'h44e33619, 32'h44e49ac2},
  {32'h4348b298, 32'hc48fe596, 32'hc36b417a},
  {32'h438311b4, 32'hc3f99292, 32'h44a1c3a0},
  {32'hc34a6ace, 32'hc42527e6, 32'hc296f286},
  {32'h43f2a233, 32'h42a435a8, 32'h428d86d4},
  {32'hc36832e0, 32'hc5317ddd, 32'hc2736d80},
  {32'h43070777, 32'h450b0e49, 32'h43229c3f},
  {32'hc4262173, 32'hc40f4d77, 32'hc4089ebb},
  {32'h43750c1c, 32'h4487ffba, 32'h44b576bc},
  {32'h430bce60, 32'hc365247d, 32'hc4c3ceef},
  {32'h4425d0a8, 32'hc358dc5e, 32'hc3cb3e78},
  {32'hc3ab5570, 32'hc4b73c67, 32'hc334c885},
  {32'h42c5bb60, 32'h454038b1, 32'h43bebf69},
  {32'h441eda9e, 32'hc4ee10d4, 32'h43347190},
  {32'hc42bdafc, 32'hc3939711, 32'hc334c862},
  {32'hc2930420, 32'hc4da8406, 32'h438c3f2a},
  {32'hc35c4050, 32'hc3321f92, 32'h4307387f},
  {32'h44f89252, 32'h43382c02, 32'hc2de73cf},
  {32'hc56a4839, 32'hc41241b9, 32'hc3727c19},
  {32'h4573aeb0, 32'hc30348c9, 32'hc43c04b6},
  {32'h44351e5d, 32'h43a91441, 32'h43f8ee4e},
  {32'hc52afd65, 32'h44605aed, 32'hc402ae77},
  {32'h450a548b, 32'hc29459d8, 32'h43f94cad},
  {32'hc3135609, 32'h44857271, 32'hc41fea9a},
  {32'h434c4198, 32'hc4bdbe45, 32'hc37913f1},
  {32'h4338b542, 32'h455f67fd, 32'hc2f98a75},
  {32'h43f73c5a, 32'hc4a7d9a8, 32'hc35e1c85},
  {32'hc532b5ba, 32'h43e47271, 32'hc2d19d58},
  {32'h42158e20, 32'hc54da5c6, 32'hc3db66d2},
  {32'hc4cb35b2, 32'h4334bdea, 32'hc2983bac},
  {32'h44699b48, 32'hc368c42e, 32'h44943309},
  {32'hc4d3db97, 32'h440c3bea, 32'h4348a816},
  {32'h45372787, 32'hc2d4d3c1, 32'h442ba61d},
  {32'h42db36b0, 32'h44ea92da, 32'h44150d56},
  {32'hc2638440, 32'hc50e52b6, 32'hc320491e},
  {32'h420b2f78, 32'h430e6321, 32'h44122ac8},
  {32'h450e3943, 32'h4400e4fa, 32'hc44d8f44},
  {32'hc46bc121, 32'h43bb0f1c, 32'h43b13868},
  {32'h4548c2f3, 32'hc44649ec, 32'h43193552},
  {32'hc3bde6a8, 32'hc4873611, 32'h448ab339},
  {32'h449ce5b7, 32'hc3b81169, 32'hc448d5c2},
  {32'h44ce43a1, 32'h440a1661, 32'h4382aba4},
  {32'h43945c80, 32'hc454c165, 32'hc4f34985},
  {32'hc4b6a693, 32'h440660cc, 32'hc3abfc55},
  {32'h4144466c, 32'h412ad9f1, 32'hc4fb80d8},
  {32'h43803e3c, 32'h449c9b42, 32'h4492f195},
  {32'hc448f488, 32'hc4cbd47b, 32'hc483af21},
  {32'h45000641, 32'h41fa3270, 32'h4261e66b},
  {32'hc4a582ba, 32'hc3a23110, 32'h444bb0db},
  {32'h43a9dc2c, 32'h4431fcff, 32'hc4292ba0},
  {32'hc51a53c5, 32'hc46a3fda, 32'h433ba564},
  {32'h4423eb7e, 32'h44ab7590, 32'hc355b5e6},
  {32'h42ec68d0, 32'hc424c390, 32'hc46990fe},
  {32'h448b23ea, 32'h44c15392, 32'h44086d1c},
  {32'hc52dc866, 32'hc404d917, 32'h43238751},
  {32'h44c87658, 32'h4404c767, 32'h440ce06e},
  {32'hc4e5d0f8, 32'hc414709b, 32'h43fa94b0},
  {32'h44207709, 32'h441d4d74, 32'hc4dec01e},
  {32'hc503c3cb, 32'hc3c19740, 32'h41c35510},
  {32'h4407eca2, 32'h4499fecc, 32'h44333723},
  {32'h42886990, 32'hc410d0ae, 32'hc4aec87f},
  {32'h44435899, 32'h442690af, 32'h43ff6e2a},
  {32'hc3a2d584, 32'hc37a4e82, 32'hc4a45875},
  {32'h442e46b6, 32'h44b98f44, 32'h43579d98},
  {32'hc3610a68, 32'h410c9c91, 32'hc456e42d},
  {32'hc4083c50, 32'h430d899d, 32'h4364dce6},
  {32'hc50e2c66, 32'hc40268e6, 32'hc488b268},
  {32'h452a1e25, 32'h43ba1803, 32'hc3d1b59a},
  {32'hc39c51c6, 32'hc47464eb, 32'hc45da67d},
  {32'hc3c86f7a, 32'h4514a661, 32'hc35f624e},
  {32'hc4f38db2, 32'hc2297b53, 32'hc34e1eb7},
  {32'h43c779f8, 32'h44df958b, 32'h445088cf},
  {32'h43755e8e, 32'hc5032769, 32'hc471be3c},
  {32'hc34ac6bc, 32'hc213b208, 32'h430fe4c8},
  {32'h452d65fe, 32'hc4440566, 32'hc2457900},
  {32'hc5524c7c, 32'hc312739f, 32'h43898638},
  {32'h4327bd10, 32'h45104237, 32'h441ae5f5},
  {32'h43ab57d1, 32'hc43a2578, 32'h439b5bd5},
  {32'h446b242e, 32'h4491a731, 32'h43ff6454},
  {32'hc48d06a2, 32'h43630274, 32'h43e20030},
  {32'hc4aeabea, 32'hc3ab3657, 32'hc34f1607},
  {32'hc44fce87, 32'hc4106f25, 32'hc3fabcdc},
  {32'h453efd8b, 32'hc2e77a20, 32'h4409e410},
  {32'h44e6e861, 32'h437805d1, 32'h4141569d},
  {32'h44aa95ff, 32'h44091dbb, 32'hc181086d},
  {32'hc3a1ecf0, 32'hc216074e, 32'hc3f0a691},
  {32'h4407ae98, 32'hc2434f90, 32'hc453edec},
  {32'hc37ac508, 32'hc4cca0aa, 32'h43ae8394},
  {32'h4341750e, 32'h43e9a46e, 32'hc507f017},
  {32'hc4fc1a41, 32'hc2090ed2, 32'hc3a52d87},
  {32'h44dd73dd, 32'h43c75ff9, 32'h4394fbcc},
  {32'hc35ec4e8, 32'hc47aff37, 32'hc3ebdbac},
  {32'hc4854716, 32'h4331c8d7, 32'hc3a19129},
  {32'hc52cd9db, 32'hc463abe2, 32'hc33d8eab},
  {32'h4460f368, 32'h447c4aab, 32'hc4d04346},
  {32'h43aa38fe, 32'hc0623796, 32'h43b2b25d},
  {32'h4332058e, 32'h44bdb262, 32'hc39c7148},
  {32'hc276fd23, 32'hc49509da, 32'h410878d0},
  {32'h422a820c, 32'h4018a90f, 32'hc351812a},
  {32'hc56267b2, 32'hc42c3398, 32'h43cecd9b},
  {32'h457a578a, 32'hc19bd1e0, 32'hc3eb15a3},
  {32'h4328bfd3, 32'hc4608d4d, 32'hc3ee795a},
  {32'hc53b89ef, 32'h43e0638e, 32'h43561b77},
  {32'hc45325bd, 32'hc4272373, 32'hc06d4478},
  {32'hc2bdb3e6, 32'h45729e16, 32'hc3373437},
  {32'h4514c4fe, 32'hc41443f0, 32'h41c72d38},
  {32'h44b1078b, 32'h4362fdab, 32'h4261551f},
  {32'h454341a1, 32'h43b5b140, 32'h42bcc54b},
  {32'hc5586e63, 32'hc34ed557, 32'h4381e8ca},
  {32'hc483c472, 32'hc27c0377, 32'h43b06a7f},
  {32'hc42feabf, 32'h44c131f6, 32'h42a44062},
  {32'h43a05e80, 32'hc4139418, 32'h4457c225},
  {32'hc379cc3c, 32'hc40282e6, 32'h44071c55},
  {32'h447e144f, 32'hc3174a52, 32'h44a88b2f},
  {32'hc2edb414, 32'h438e95ba, 32'hc4c32a3a},
  {32'h4433e936, 32'hc379c2ed, 32'h42a6320b},
  {32'hc399611e, 32'hc3b8b45a, 32'hc51b4929},
  {32'h443178f8, 32'hc37edfeb, 32'h44885483},
  {32'h4401a2db, 32'h43b917ee, 32'hc21d9801},
  {32'h44dc9189, 32'hc45647ef, 32'h43302a16},
  {32'hc529fbc8, 32'h442e37d4, 32'hc4199d9a},
  {32'h44f05a4e, 32'hc35b8d64, 32'h3fa4a500},
  {32'hc27a3ee0, 32'hc2f4c8b4, 32'hc51183e5},
  {32'h43e76f6b, 32'hc5572e0d, 32'h42b7c4b3},
  {32'hc4558390, 32'hc39133cf, 32'hc3bf0c43},
  {32'h453247a8, 32'h43880581, 32'h43cdb197},
  {32'hc53865fa, 32'hc1651254, 32'hc4b4a5cc},
  {32'hc3d6af6a, 32'hc26d73a2, 32'h446a8549},
  {32'hc3c0db4e, 32'h448dfe88, 32'hc40bccc3},
  {32'h44255a4a, 32'h44963d62, 32'h4433c595},
  {32'hc4bd3683, 32'h43be2c9a, 32'hc390d803},
  {32'hc4036198, 32'h42dca52b, 32'hc2eabdad},
  {32'h45132c1a, 32'hc378d3eb, 32'h444209a7},
  {32'hc47daa6c, 32'h4034e1ba, 32'hc3b4b385},
  {32'h450e99b4, 32'h43a180de, 32'hc2c66861},
  {32'hc44a7026, 32'h439a82cb, 32'hc42a4c30},
  {32'h45042050, 32'hc3c351ec, 32'h43ccbe0c},
  {32'h44a11130, 32'hc4017f8a, 32'h444224fa},
  {32'hc49c8df8, 32'hc4ae581d, 32'hc41a3b20},
  {32'h43e48a56, 32'hc3a35b98, 32'h433c1d8e},
  {32'h43e311db, 32'hc2c9b7b2, 32'h44d806cc},
  {32'hc4c3658c, 32'h42572ac3, 32'hc4693f74},
  {32'hc379f9f4, 32'hc3beeb66, 32'h453fe6b8},
  {32'hc23711d0, 32'h43b6ec6f, 32'hc4b7ea01},
  {32'h43f9b088, 32'hc50a44de, 32'hc2e0c06d},
  {32'hc4db8c50, 32'h4305a508, 32'hc4928d77},
  {32'hc4f7907e, 32'h43894ecd, 32'h423226dc},
  {32'hc4bd7f2e, 32'hc22ad0c0, 32'hc43ecad6},
  {32'hc3915954, 32'hc2ac2888, 32'h430dfd29},
  {32'h442a8992, 32'h40ff5d8e, 32'h42fb77db},
  {32'h442716c7, 32'hc265831a, 32'h43636abf},
  {32'hc3afc52e, 32'h45417020, 32'h429a987c},
  {32'h44e26f02, 32'hc272a8ae, 32'h43a05f81},
  {32'hc4c15fea, 32'h44154a90, 32'h43a5f358},
  {32'h43bb2790, 32'hc520e895, 32'h431e46da},
  {32'hc3ae49ec, 32'hc40755d2, 32'h43147b1f},
  {32'h44b9641b, 32'hc35cb18f, 32'hc436348e},
  {32'h43098f75, 32'h45097dfd, 32'h4496d694},
  {32'hc412b59a, 32'hc4a2355e, 32'h4435e56f},
  {32'h440a1a6c, 32'h441e222f, 32'hc46e9943},
  {32'hc505d6e6, 32'h43ad9a8c, 32'h40f5f41c},
  {32'h44ca7b92, 32'h44804b05, 32'hc3c2c7f1},
  {32'hc474f14c, 32'hc4979b54, 32'h4391f96f},
  {32'h4422dfa3, 32'h4454fc74, 32'hc31c71cf},
  {32'h43a2c421, 32'h449b28b1, 32'hc3537a68},
  {32'h43a689bc, 32'hc45ebc8b, 32'h44ea2f26},
  {32'h431b3f34, 32'hc4c37253, 32'hc4db5bc6},
  {32'h4254eab2, 32'h43f9bbd7, 32'hc4b04b4c},
  {32'h42cd842f, 32'hc4b23ee1, 32'h4308f131},
  {32'h44a9ce16, 32'h43aa363c, 32'hc41f55d6},
  {32'hc4a99035, 32'hc3409390, 32'h44c19826},
  {32'h44df6cbe, 32'h437da445, 32'h415938a6},
  {32'h43a491f6, 32'hc3a82ac0, 32'h44d5f1ff},
  {32'hc210f998, 32'h4400aa9c, 32'hc36e985d},
  {32'hc48a215d, 32'hc40eccf4, 32'hc24e925b},
  {32'h438acea8, 32'h42d093b5, 32'h4203c1e8},
  {32'hc4e3ac0d, 32'hc4832eed, 32'h42b8e2e1},
  {32'h44013a68, 32'h44f03a0c, 32'h42ebce48},
  {32'hc4ec48e5, 32'hc2e4aec4, 32'h43b103d3},
  {32'h448ad092, 32'h444e3df1, 32'hc3243aca},
  {32'hc42cdf22, 32'hc4dd728a, 32'h43a5b6de},
  {32'h453fcd66, 32'hc3204993, 32'h4211fd06},
  {32'h42eddc5a, 32'h4447ab0d, 32'h432c2458},
  {32'hc337ece8, 32'h448c8105, 32'hc48b06f1},
  {32'h43593164, 32'h4554dca5, 32'h4438568e},
  {32'h414de800, 32'hc26fd181, 32'hc4b97b62},
  {32'h439b5e7a, 32'h44ee8a37, 32'h43d7d15a},
  {32'hc4901b4f, 32'hc42636a1, 32'h438e6ae9},
  {32'hc4339852, 32'h43425c62, 32'h43a1a783},
  {32'hc3effea4, 32'hc06bf0ae, 32'hc483b1bd},
  {32'h445594c4, 32'h449fb3f2, 32'h444cad35},
  {32'hc4bf7818, 32'hc3f0ba5f, 32'h41ac9516},
  {32'h43cefb7c, 32'hc417651d, 32'h443b4435},
  {32'h43d7b47c, 32'h43b7bef3, 32'hc4cf43d3},
  {32'hc3bc5f8c, 32'h4487b04d, 32'h430896aa},
  {32'hc4d12fb7, 32'hc3e5e51d, 32'hc3075e16},
  {32'h446c89ac, 32'h43a2e560, 32'h4203efcc},
  {32'hc394df46, 32'hc3184153, 32'hc49c0eec},
  {32'hc2940d2e, 32'h43bff9fb, 32'h450010e2},
  {32'hc4a90ee7, 32'hc3ddaca6, 32'hc3ff4121},
  {32'h44af8467, 32'h44018a8b, 32'h42d1b448},
  {32'hc459141f, 32'hc518650c, 32'h43c06c6c},
  {32'h44b1269e, 32'h44bd9314, 32'h41fb2b18},
  {32'hc50f9d99, 32'h43acf413, 32'hc3a6f395},
  {32'h443f56b8, 32'h44c4d0d9, 32'hc20cb58d},
  {32'h42495e98, 32'hc54084f6, 32'h4159c799},
  {32'h441352e2, 32'h4385265c, 32'h4386a635},
  {32'hc590b36a, 32'h4353915d, 32'hc3cc3f1d},
  {32'h42756980, 32'hc3ce0125, 32'h440f92cf},
  {32'hc29df5d6, 32'h426fec02, 32'hc4e48f22},
  {32'hc3a1dc9c, 32'hc358d27a, 32'h4405975b},
  {32'hc3f667eb, 32'h4292056a, 32'hc3ad4103},
  {32'h43bff620, 32'h44018bef, 32'h44e7bf66},
  {32'hc390f4c4, 32'hc101d95a, 32'hc5681021},
  {32'h448498ee, 32'hc3464cf8, 32'h43d90028},
  {32'h43dd2736, 32'hc3d7c786, 32'hc53795c0},
  {32'hc507a33c, 32'h43f2a3a6, 32'h430605fd},
  {32'h44b4c000, 32'hc3dcc165, 32'h42407132},
  {32'hc424ec93, 32'h42d6d33f, 32'h43e9344f},
  {32'h437123e8, 32'h44af24a9, 32'hc495b459},
  {32'hc3e0c812, 32'hc27191be, 32'h4420ad2f},
  {32'hc2d7596b, 32'hc4ae95dc, 32'hc43effef},
  {32'h4316cffa, 32'h42f4f3f8, 32'h450bb08a},
  {32'h44832858, 32'h41a5c688, 32'hc45b558d},
  {32'hc393d0e9, 32'h43e40f10, 32'h450a60c2},
  {32'h451c1335, 32'h4388cc74, 32'hc2c82c72},
  {32'hc5088434, 32'hc2c59b66, 32'h43c75a43},
  {32'h441a1e94, 32'hc508f094, 32'hc3a1535a},
  {32'hc50832f0, 32'h44ae3019, 32'h42119e06},
  {32'h45042a0e, 32'h42943714, 32'hc3e110ca},
  {32'hc3e06ad1, 32'h452c2719, 32'hc39afd66},
  {32'h451ed334, 32'hc3e0d78b, 32'h4304d41b},
  {32'hc2e1d237, 32'h445a384c, 32'hc31e36a1},
  {32'h45132b98, 32'h42fa6777, 32'h43aebfbb},
  {32'hc54e384b, 32'hc37cd35a, 32'h4343f3b2},
  {32'h45755c35, 32'hc3907f61, 32'hc2a72575},
  {32'h44db313e, 32'hc0f87ad6, 32'h43175015},
  {32'hc47408d8, 32'hc3c60469, 32'hc462b332},
  {32'h446ca1e4, 32'hc3082f80, 32'h44d7d9a3},
  {32'h44f4bf6b, 32'h42696243, 32'hc2dd5a3e},
  {32'h440a3356, 32'hc52e3c44, 32'hc314a3b8},
  {32'hc48e078d, 32'h44bdc56d, 32'hc0f6d5bd},
  {32'h43a39ab2, 32'hc3a98781, 32'h4350d593},
  {32'hc4f0f8da, 32'h44a505c6, 32'h42c7dc64},
  {32'h44ac3344, 32'hc4422e89, 32'h44013907},
  {32'hc42f94c0, 32'h42b1f879, 32'hc1a6f476},
  {32'h442e941a, 32'h439986d2, 32'hc4159b39},
  {32'hc49396bc, 32'h444f4bf5, 32'h44215e26},
  {32'hc3afd90f, 32'hc3156f7c, 32'hc3e18cc8},
  {32'hc300d6dc, 32'h43d304ec, 32'h4505220a},
  {32'h43c947ad, 32'hc38265b8, 32'hc5011a0a},
  {32'h425b6180, 32'h442d1094, 32'hc34271be},
  {32'h448b64d4, 32'hc3abda6e, 32'hc41cd131},
  {32'hc3948ea8, 32'h430056a4, 32'h4181b10c},
  {32'h454018ba, 32'hc33790aa, 32'h41abfd80},
  {32'hc515ec4d, 32'hc47028b8, 32'h44b204f7},
  {32'h444ac90d, 32'h43ee6436, 32'hc4c0ec5a},
  {32'h43563614, 32'h44c2d4d0, 32'hc31dea05},
  {32'hc0f3c560, 32'hc525b148, 32'hc43fc1c8},
  {32'hc4692616, 32'h44a220ff, 32'hc29bfc06},
  {32'hc496751e, 32'hc33a55c6, 32'hc36e3475},
  {32'hc4377422, 32'h449147ad, 32'h44339c09},
  {32'h44c1845f, 32'hc33cf07b, 32'hc491a3ff},
  {32'hc287fd20, 32'h4313e086, 32'hc52b4773},
  {32'hc4a38275, 32'h42bb1d6c, 32'h44a1ceb5},
  {32'h44830a6f, 32'h43aab2a6, 32'hc408292a},
  {32'hc3150438, 32'hc4f432e6, 32'h42c6413a},
  {32'h4531dbb3, 32'h43141dc9, 32'hc2c62e76},
  {32'hc50d785c, 32'hc39942b0, 32'h431fc204},
  {32'h44b474a4, 32'h4436c645, 32'h4331f1cc},
  {32'hc47f486c, 32'hc5026ffa, 32'h423851e6},
  {32'h4500aa69, 32'hc43cf778, 32'hc38d5fc4},
  {32'hc3f7274f, 32'hc406b961, 32'h44a2cf1d},
  {32'h41edd68a, 32'h43db7730, 32'hc52e74e4},
  {32'hc50ebe67, 32'hc2fe6534, 32'h4385ea9b},
  {32'h4281bab8, 32'h4497d57f, 32'h4404a725},
  {32'hc50bf1e8, 32'hc42fe4fe, 32'hc430575f},
  {32'h43047f31, 32'h44158e2f, 32'h447d1121},
  {32'hc461ebc0, 32'hc371c639, 32'hc4d774bd},
  {32'h44f22656, 32'h442c2206, 32'h4405d196},
  {32'h42e1ed82, 32'hc32bb47d, 32'hc49903fb},
  {32'h43bc8dd5, 32'h433b135f, 32'h44be2d8e},
  {32'hc502c416, 32'h43a2480a, 32'hc3b46ade},
  {32'h453ac46c, 32'h4306cbe2, 32'hc4612979},
  {32'hc34d3563, 32'hc50b34c6, 32'hc3ace2c3},
  {32'h436d3b73, 32'h43f629fb, 32'h44adb4a5},
  {32'hc43d2b77, 32'hc4414cc7, 32'hc3dbba60},
  {32'h450795cd, 32'h440037e9, 32'h444bdb39},
  {32'hc35cefa8, 32'hc42bc6b2, 32'hc559ba35},
  {32'hc185d788, 32'h433e2f7f, 32'h44884728},
  {32'h44510a87, 32'hc3f6c491, 32'hc348613f},
  {32'hc4b3ce20, 32'h4405409a, 32'hc49d353a},
  {32'h43988190, 32'h445c1725, 32'hc1476908},
  {32'h44c960f3, 32'hc3a8707a, 32'h422eec6d},
  {32'h44ae19ee, 32'h44984ee4, 32'hc382f20c},
  {32'h4364a1f6, 32'hc52219fb, 32'hc34087ee},
  {32'h45316cd3, 32'hc331b68e, 32'hc3024952},
  {32'hc54d6c51, 32'hc31fcc93, 32'hc36fbef9},
  {32'h436113f8, 32'h44a9ca52, 32'h4493ad5f},
  {32'h44242cad, 32'h429aa5f9, 32'h4373a8b8},
  {32'h4055ea00, 32'h4495af64, 32'hc50c7cbc},
  {32'h42c2ea51, 32'hc4df58a5, 32'hc29f0fe1},
  {32'hc4811a56, 32'h43c07cac, 32'hc3541689},
  {32'hc44178e8, 32'hc4a292b0, 32'h43e7d6e3},
  {32'h44b81072, 32'h440310ac, 32'hc40526b3},
  {32'hc49ff147, 32'hc43738c8, 32'hc24a5c22},
  {32'h44848c62, 32'hc239aeb2, 32'hc4671082},
  {32'hc4c57661, 32'h4267faa8, 32'h447d3fac},
  {32'h43e92500, 32'h438a882e, 32'hc3befdd6},
  {32'hc3d77404, 32'hc5632ab2, 32'hc3c231fe},
  {32'h4484bf42, 32'h444f260e, 32'h431aa7c4},
  {32'h42aba72a, 32'h43186172, 32'h41838312},
  {32'h4504c83b, 32'hc35b9248, 32'hc4a101b1},
  {32'hc4beae3c, 32'hc3b8d907, 32'h4226ff69},
  {32'h44d2c755, 32'h44029aa0, 32'hc0bfc3fb},
  {32'hc41783e7, 32'h43d973b0, 32'h45429d0f},
  {32'h44b7b7fc, 32'h4368729e, 32'hc443dc08},
  {32'h42b952c0, 32'hc52b7a48, 32'h43a3e3fe},
  {32'hc4cd7d70, 32'h429bb7f9, 32'h4427352c},
  {32'h4386a09b, 32'hc4c51bba, 32'hc28c050d},
  {32'hc55cc072, 32'h43fe18f6, 32'h43f815f1},
  {32'h44c92d35, 32'hc3970dd2, 32'hc2e75a5d},
  {32'hc33b1834, 32'h4314fbba, 32'hc3035115},
  {32'h45200494, 32'hc3be2e98, 32'hc4102b9a},
  {32'hc4c722b2, 32'hc335e8c9, 32'hc3f09f4f},
  {32'h4478793f, 32'h439ba1f6, 32'h44279e47},
  {32'hc39e2674, 32'h433a1916, 32'hc3b913a2},
  {32'h4496432e, 32'hc31a6172, 32'h41290258},
  {32'h44b58f83, 32'hc1f7b870, 32'hc3dd5416},
  {32'h44317a59, 32'hc4d50e33, 32'hc2ca5bdb},
  {32'hc43d0670, 32'h42c9c364, 32'hc4b37939},
  {32'h43894126, 32'h430f9e4e, 32'h44507b6a},
  {32'hc4bb02af, 32'hc26c2053, 32'hc439f082},
  {32'h4377dea0, 32'hc432ac06, 32'h43af933a},
  {32'hc4a9499e, 32'hc27dcb06, 32'h43772253},
  {32'h44b2d100, 32'hc46cfcb8, 32'h4413d692},
  {32'hc4db7dd1, 32'h44c786e8, 32'hc3089e1b},
  {32'h43a0fb46, 32'hc39455ef, 32'h43a01d93},
  {32'hc4ae7f80, 32'h437fe0d4, 32'hc4ec869f},
  {32'h446d5aa0, 32'hc3e4a155, 32'h448a38f6},
  {32'h447e940a, 32'h413983a1, 32'hc4197d51},
  {32'h449290dc, 32'hc3d0b1fa, 32'h438b0f48},
  {32'hc43ee7a6, 32'hc39affca, 32'hc560fc42},
  {32'hc3aff5eb, 32'h42257f01, 32'h42a7d30f},
  {32'h44219958, 32'h44005fa2, 32'hc48202f1},
  {32'h4170a800, 32'h44d68372, 32'h44c2c4d7},
  {32'h44b7dd14, 32'hc3e1d9f9, 32'hc39576d6},
  {32'hc3a517b5, 32'hc379c4f8, 32'hc4cbd3c7},
  {32'h43a4b068, 32'hc4aa212e, 32'h44454730},
  {32'hc4b4e983, 32'h4029d741, 32'hc49ce244},
  {32'h44531c5e, 32'h42356ae4, 32'h43fe2b11},
  {32'hc300d6f9, 32'h44fabbe5, 32'hc39f48c9},
  {32'h4423dd99, 32'hc4252fbf, 32'h44eb311c},
  {32'hc2248d1f, 32'hc43f8c9d, 32'h4522ae4b},
  {32'h41f1f4ca, 32'h451640f3, 32'hc504a672},
  {32'hc3535e5c, 32'h42c5b8a8, 32'h44937dee},
  {32'hc4f52bc2, 32'hc3cfbf7a, 32'h42f12aa2},
  {32'hc4e52d8e, 32'h42d83eca, 32'h44128ae5},
  {32'hc0f2cb40, 32'hc25a1afb, 32'h453eddae},
  {32'hc4d7720c, 32'h43c8696f, 32'h43f40d55},
  {32'h443e4d12, 32'hc2684b59, 32'h450e317e},
  {32'h43e8d0fc, 32'h44624695, 32'hc4257490},
  {32'hc4892d91, 32'h427574dd, 32'hc1bd9749},
  {32'hc5849a02, 32'h434bdd40, 32'hc2a01bd2},
  {32'h44aab27a, 32'hc282ac2f, 32'h438cd6a4},
  {32'hc5055ead, 32'h40a6ebf0, 32'hc3469dfa},
  {32'h44ab630e, 32'h42b4776a, 32'h43d15e68},
  {32'hc4512d1a, 32'h44be7fdc, 32'hc31df6e2},
  {32'hc42d843c, 32'hc386d613, 32'hc2905439},
  {32'hc3d5d64a, 32'h4501ddd2, 32'hc34d59f0},
  {32'hc3359ad3, 32'hc57470d7, 32'h42a4ace6},
  {32'h440a71f6, 32'hc41cd8cb, 32'h4337f77e},
  {32'hc36a6e5e, 32'hc509b821, 32'hc4ab71f6},
  {32'hc2940da9, 32'h4443dec2, 32'h45031db6},
  {32'hc4ad820f, 32'hc4252b76, 32'h42dbf76d},
  {32'h44586b14, 32'h44441b8f, 32'h4289b93b},
  {32'hc45fc586, 32'hc49226af, 32'hc2c26a07},
  {32'h44fe021f, 32'h43fdb16a, 32'hc25e7dd9},
  {32'h42ed3c48, 32'hc47c7973, 32'h444d5d7f},
  {32'hc42c8bdc, 32'hc37493bc, 32'hc24b03a8},
  {32'hc417994e, 32'hc30b9c2f, 32'h42d5c20f},
  {32'hc45ec74d, 32'h4409f98b, 32'h43bf0aad},
  {32'hc1247630, 32'h445202bc, 32'hc5180f42},
  {32'h43a1088c, 32'h449b6aea, 32'hc3c3b18a},
  {32'hc403dddc, 32'h436e26b7, 32'h44c45fcc},
  {32'hc48c53af, 32'h4390bf76, 32'hc37df169},
  {32'hc3f8494c, 32'h43ae2200, 32'h450e4513},
  {32'h447b9698, 32'h44318b0c, 32'hc430ef0e},
  {32'hc48506e0, 32'hc3ed479e, 32'hc29e4c0c},
  {32'h452c9441, 32'hc39a70a9, 32'h430409dc},
  {32'hc55a985e, 32'hc337d33d, 32'h420aae50},
  {32'hc48f2c19, 32'hc23445a0, 32'h430946c5},
  {32'hc417315f, 32'hc4956015, 32'h433117ae},
  {32'h43daf668, 32'h45178486, 32'hc261feb4},
  {32'h43a3a407, 32'hc43ef3eb, 32'h41a8a0a6},
  {32'h43b27f0a, 32'h44257f9e, 32'hc37ce108},
  {32'hc5730ad9, 32'h43e5054e, 32'h43cec7e5},
  {32'h44bf5dcb, 32'hc23de29c, 32'hc33b3631},
  {32'h445b7e7e, 32'hc47c1009, 32'h422c66e2},
  {32'hc341d701, 32'hc51dc497, 32'hc304fa82},
  {32'h428c4ab0, 32'hc4bbff14, 32'h44d8a9d5},
  {32'h444fe07e, 32'hc3e6b00b, 32'hc117c4b4},
  {32'h44d129ec, 32'h4282bf74, 32'h448540df},
  {32'h42c64d69, 32'hc51976c0, 32'h43371c85},
  {32'h44daaf9d, 32'hc39afd70, 32'h43544230},
  {32'hc4882336, 32'hc422143e, 32'hc3204b1e},
  {32'h449ffb61, 32'h43fc2277, 32'h44c4f9be},
  {32'hc5144cd0, 32'h439fc7cb, 32'h442dcda4},
  {32'hc3371e37, 32'hc4831b85, 32'h44931d4d},
  {32'hc331b3e0, 32'hc2a848c6, 32'h4314b449},
  {32'hc37360bf, 32'h44972644, 32'h432cf24b},
  {32'hc42e6f5e, 32'hc4df6e27, 32'hc38f38a8},
  {32'h4232f299, 32'h42737de9, 32'h447f2ad7},
  {32'h43755611, 32'hc460fb35, 32'hc381cea2},
  {32'h452d622c, 32'h4300e4ac, 32'h44075864},
  {32'hc377ffeb, 32'hc4a415fd, 32'hc4956802},
  {32'h43e7adf4, 32'h4361c558, 32'h44447634},
  {32'hc563628a, 32'h432d6b2b, 32'hc27f372f},
  {32'h44c43368, 32'h44bd5e54, 32'h42d846fa},
  {32'hc502930f, 32'hc39766aa, 32'hc27a4797},
  {32'h432be574, 32'h453139df, 32'h4406346c},
  {32'hc43cfdef, 32'hc4cf8901, 32'hc3a5a94a},
  {32'h44db0c4c, 32'h437ceaa4, 32'h440bf636},
  {32'hc588c1ba, 32'h434b31f9, 32'hc2416202},
  {32'h456ebe9a, 32'h438143f6, 32'h43ce22bb},
  {32'h447d8740, 32'hc3775ba1, 32'hc48c5856},
  {32'h40fc88e4, 32'h44938cd0, 32'h4302881e},
  {32'h44541aed, 32'h439d6f2e, 32'hc2f1b468},
  {32'hc4cb70e4, 32'h4407af69, 32'hc2b656b0},
  {32'hc3cc2122, 32'hc3e86951, 32'hc51c18fc},
  {32'hc4846115, 32'h44456ac2, 32'h4429e809},
  {32'hc2ce878c, 32'hc41ea4bf, 32'hc5203f24},
  {32'hc3e6dca5, 32'h43736f2a, 32'h4524fb13},
  {32'hc3fd2918, 32'hc3e7d610, 32'hc45be098},
  {32'hc3f2cdde, 32'h448b3393, 32'h4481b275},
  {32'h43fca75e, 32'h442d8044, 32'hc4971e1d},
  {32'h4419b8ba, 32'hc1598f49, 32'h4385efed},
  {32'h440f3796, 32'hc3a38e2e, 32'hc44d47b4},
  {32'hc4043979, 32'h4520ce80, 32'h432241c0},
  {32'hc3886eee, 32'h43fb5bfc, 32'hc49619c8},
  {32'hc523ba7e, 32'h4240a659, 32'h43854dee},
  {32'h44972ba4, 32'hc416c559, 32'hc49c7153},
  {32'h443687c2, 32'h44283778, 32'h4386bd50},
  {32'h44095a44, 32'hc4ca5552, 32'hc3581421},
  {32'hc38cca4c, 32'h45095530, 32'h43fc9ab6},
  {32'h44a1c1ea, 32'hc391627e, 32'hc3c1c7cf},
  {32'hc51d6a02, 32'hc3d19cdc, 32'h44017fb7},
  {32'h4510a964, 32'hc2549d58, 32'h411eba6a},
  {32'h44d91bdc, 32'h4166c254, 32'h432cc2d7},
  {32'hc30bac00, 32'h43943419, 32'hc3a36f84},
  {32'hc539b65a, 32'hc3ce92b0, 32'hc0cbfc1c},
  {32'h441f7cf6, 32'hc442f73d, 32'hc38b282e},
  {32'h44d2a806, 32'hc30d2044, 32'hc403a94e},
  {32'hc39e99ac, 32'h445b583d, 32'hc50876e1},
  {32'h44c84f2c, 32'hc3233b17, 32'h44c0ea36},
  {32'hc4d26e46, 32'h436abb92, 32'hc340f63c},
  {32'h43d38c58, 32'h434ecbb9, 32'hc3805a97},
  {32'hc53e2862, 32'hc204ab9d, 32'hc278d34e},
  {32'hc3925b8e, 32'h40b011f0, 32'h435bb14d},
  {32'hc4e5f482, 32'h448d0551, 32'hc19779a1},
  {32'h45082552, 32'hc3e856ed, 32'h42b486df},
  {32'h44fe144e, 32'h43e01afe, 32'hc2ddb08a},
  {32'h452f7c1b, 32'h42b0fa25, 32'hc09a53dc},
  {32'hc48f2261, 32'hc28ca4cf, 32'h440fb011},
  {32'hc4d6caa9, 32'h41bc1a8d, 32'h436f0171},
  {32'h42d1228c, 32'h425b42f0, 32'h44dce274},
  {32'h449b2c5d, 32'hc41f6ff5, 32'h4181fa26},
  {32'hc3968d74, 32'h449d3fa8, 32'h4440efab},
  {32'h452d15ee, 32'hc3bc2f1b, 32'hc3124a9a},
  {32'hc5047858, 32'hc3ce1fdb, 32'h43f53f53},
  {32'h43d2b834, 32'hc28f3da3, 32'hc423c94b},
  {32'hc4fa0546, 32'h443d6419, 32'h4454db34},
  {32'h4432da9c, 32'h438e93cf, 32'hc4b11e58},
  {32'hc38abb01, 32'hc2b831d6, 32'h44950cd7},
  {32'h43105426, 32'hc50b1106, 32'hc42759fb},
  {32'h43ed65fb, 32'hc2ca8c9b, 32'h452e7a50},
  {32'h44ef125e, 32'hc2c798b2, 32'hc2701298},
  {32'hc4fb6b46, 32'h4466a6c4, 32'h44558fdb},
  {32'h4389051c, 32'hc51cb042, 32'hc3935aa2},
  {32'h44b317be, 32'hc3d5e234, 32'h43a345b5},
  {32'hc570b4f9, 32'hc2f2705e, 32'h441ca766},
  {32'hc27102a7, 32'h434594b8, 32'hc43f44d4},
  {32'hc44628b3, 32'hc4a24607, 32'hc3949bd3},
  {32'h442dc8e4, 32'h4414bcbb, 32'h4336b35e},
  {32'h44909157, 32'hc49ea425, 32'h42fae127},
  {32'h4560740a, 32'h4405b2ad, 32'h43070669},
  {32'hc3e62376, 32'hc56db841, 32'hc380ac47},
  {32'h443bc7ee, 32'h43252e83, 32'hc17797b3},
  {32'hc47cd54e, 32'hc1a84c17, 32'h4506b406},
  {32'h4462a3a6, 32'hc3c20281, 32'hc34b2548},
  {32'h43623384, 32'h44399304, 32'hc48094dd},
  {32'h44019100, 32'h4487a33b, 32'h42dec1bb},
  {32'hc4108a6a, 32'h41f43b12, 32'hc52882c7},
  {32'hc326b680, 32'h4439d03f, 32'h434dc238},
  {32'hc3bcdc4e, 32'h4123ddfa, 32'hc5259fe9},
  {32'h43101d00, 32'h454d2ff4, 32'hc3d2acc6},
  {32'h4460d945, 32'hc2b8aa23, 32'hc15d7ecd},
  {32'h450fe0f9, 32'hc34c865b, 32'h44341391},
  {32'hc58e633b, 32'h44017aa9, 32'hc293dfec},
  {32'h432e7b9a, 32'hc22f5374, 32'hc31d0954},
  {32'h435078cf, 32'hc53c63f1, 32'hc36bf1cb},
  {32'h4345eb36, 32'h449f1e32, 32'h44177d03},
  {32'h44410dd0, 32'h4336d06f, 32'hc423f7e7},
  {32'h44658852, 32'h44ad78e4, 32'h42ce04be},
  {32'hc54771de, 32'hc06284eb, 32'hc3490f24},
  {32'h44cfe614, 32'hc39057f2, 32'hc25aa55c},
  {32'h431fec91, 32'h4482704b, 32'hc4293758},
  {32'hc513e7ca, 32'hc2c81808, 32'hc2bb0e7c},
  {32'h450d627c, 32'h44035bb8, 32'h44082fe2},
  {32'hc1a66116, 32'hc497cc17, 32'h431149d3},
  {32'h455baca8, 32'h42c2c345, 32'hc40758af},
  {32'hc214236a, 32'hc5507f86, 32'h4303cdae},
  {32'h430b2394, 32'hc17c85f8, 32'hc43ec9e0},
  {32'hc552c284, 32'hc2e0eee9, 32'hc3bb75c9},
  {32'h4527c4d4, 32'hc4315750, 32'hc281d7c3},
  {32'hc4a647d2, 32'h437c4f8c, 32'hc3a6e9dc},
  {32'h4417bebd, 32'h4479e20b, 32'hc29568c4},
  {32'hc3785d90, 32'hc3f6cfa8, 32'h44c919d0},
  {32'hc48e31e8, 32'h4186ae04, 32'hc2eafa5c},
  {32'h43a0b140, 32'hc38563de, 32'h451e0aef},
  {32'h442dc64f, 32'hc3217750, 32'hc52367b3},
  {32'h42af6968, 32'h42d051e8, 32'h44c1dbb1},
  {32'h44335cb8, 32'h44a0dae6, 32'h446ce72d},
  {32'hc4858c5f, 32'h43aacc46, 32'h44f3e639},
  {32'h448dd1e2, 32'hc36d38c4, 32'h4446ea1c},
  {32'hc5080985, 32'hc429c81d, 32'h437aca3f},
  {32'h4477d030, 32'h4480ea7e, 32'hc489e5c8},
  {32'hc5396c8a, 32'hc2b4c1ad, 32'h42116a32},
  {32'h439da790, 32'h44ce94b7, 32'hc42074ca},
  {32'h42a611e8, 32'h42af8e6a, 32'h44ed1d13},
  {32'h43b9d0ce, 32'h42717168, 32'hc47d69ca},
  {32'hc515a94b, 32'hc2a44462, 32'h44201fb9},
  {32'h44d1d192, 32'h42a4b485, 32'hc49bf2cb},
  {32'h43fb56a5, 32'hc4de2516, 32'hc3943978},
  {32'hc43efa22, 32'h4526ee1c, 32'h43880979},
  {32'hc33aef9c, 32'hc31cd50c, 32'hc2ded5b3},
  {32'hc4dd765f, 32'h44aedfd0, 32'h43c465f3},
  {32'hc26a1ec4, 32'hc568d383, 32'h431cad5b},
  {32'h44845033, 32'h4317ebe6, 32'hc16d3300},
  {32'h450d930c, 32'hc41edaa0, 32'hc452baec},
  {32'hc519a9cc, 32'hc33cc7d2, 32'hc164661b},
  {32'h44c93416, 32'hc32d5d2d, 32'h445fcba3},
  {32'hc286d1b0, 32'h4444edcf, 32'hc4b9e4a7},
  {32'h43f7833a, 32'hc52a3fef, 32'h43d8a33a},
  {32'h44d5ab7c, 32'hc1c5cc9e, 32'h437de0c1},
  {32'h44cf2fe1, 32'hc3bb6b40, 32'h44913949},
  {32'hc39bcad4, 32'hc37055a6, 32'hc4fb8ae0},
  {32'h451882a6, 32'h43c9d7e9, 32'hc18c9f21},
  {32'hc3317517, 32'hc39557ff, 32'hc5471f39},
  {32'h43cfa698, 32'hc389b4cc, 32'h44b39fb3},
  {32'hc31554c0, 32'h4353929b, 32'h441ed0a5},
  {32'h447248c5, 32'hc4203d2b, 32'h44e5735b},
  {32'hc58a3b8a, 32'hc2dd0540, 32'h42976c67},
  {32'hc4423ea4, 32'hc3c9809f, 32'h43c6a63d},
  {32'hc4976b95, 32'h43d18e56, 32'hc4c4757b},
  {32'hc0c87fc0, 32'h431978a5, 32'h448ad591},
  {32'hc44dba31, 32'h44337098, 32'hc3ed9931},
  {32'h447f53d2, 32'h43aac366, 32'h45062458},
  {32'hc43a4d56, 32'hc28e3c2e, 32'hc4ad4281},
  {32'h455e0955, 32'hc3a1b840, 32'h42a77461},
  {32'h440b0fd4, 32'h44ce557b, 32'hc513cb91},
  {32'h439eeed9, 32'h429005cb, 32'h4427268f},
  {32'h440d9563, 32'hc4768595, 32'hc3354f07},
  {32'hc50bf815, 32'h431a6611, 32'h433771d8},
  {32'h437fe8ba, 32'h42eae642, 32'h4502d012},
  {32'hc4dfb136, 32'hc1126c7e, 32'hc4188484},
  {32'hc4c99f98, 32'hc3699c13, 32'h43368da6},
  {32'hc51023c8, 32'h440362e9, 32'hc2b2eb73},
  {32'hc3d31ef0, 32'hc44a4ef4, 32'h4372038b},
  {32'hc18dd9de, 32'h44123269, 32'h44fc06ac},
  {32'h4324ae9f, 32'h45135f1d, 32'hc4e94a68},
  {32'hc3928484, 32'h444ac39e, 32'h44c83f1c},
  {32'h43ce5910, 32'hc2aa5216, 32'h44a248b7},
  {32'hc554e202, 32'hc3882a5d, 32'hc1e3b5cb},
  {32'h451fea76, 32'h44231e6d, 32'hc33184ce},
  {32'hc343c6cc, 32'h445ea5e4, 32'hc3f317c0},
  {32'h44c535ca, 32'hc3ff65ba, 32'h44610fa1},
  {32'hc4690f1d, 32'h446ab839, 32'hc3d85d04},
  {32'h457cd867, 32'hc3a7e5fe, 32'h422fd63a},
  {32'hc4696866, 32'hc46ee316, 32'hc3d05835},
  {32'h44ff0735, 32'h434152f3, 32'h444a37a5},
  {32'hc4918f5c, 32'h43d708a0, 32'h43525e03},
  {32'h43b68e08, 32'hc3523d64, 32'h43c17479},
  {32'hc4441b64, 32'h44d14878, 32'hc3063a9e},
  {32'hc3afa401, 32'hc3f44c39, 32'h433f39d3},
  {32'hc5346c49, 32'h447e482e, 32'hc2c93081},
  {32'hc12a3e00, 32'hc4c320cb, 32'h4426be7a},
  {32'h443dfed2, 32'hc3ee6c55, 32'h44480398},
  {32'h450a0b14, 32'hc25bbf9d, 32'hc385f39b},
  {32'h4247f520, 32'h450e1b77, 32'h44dbee7d},
  {32'hc33c9280, 32'hc29fa236, 32'h44fa07de},
  {32'h43b4b528, 32'h449de98e, 32'hc3384c62},
  {32'h4234a7c6, 32'hc320513e, 32'h450284a3},
  {32'hc3998875, 32'h451d7b03, 32'h4384c132},
  {32'hc47ea3d4, 32'hc39d22d5, 32'h44761009},
  {32'hc4f0bb99, 32'hc304c257, 32'hc38ddee7},
  {32'h4498ec30, 32'h43442db5, 32'h42c777c4},
  {32'h43a435dc, 32'hc2b77c86, 32'h453b3008},
  {32'hc282dae0, 32'hc2e18655, 32'hc4db63c0},
  {32'h4410f00f, 32'h44d0a4a6, 32'hc320a42c},
  {32'hc43232be, 32'hc42707a6, 32'h44856eaa},
  {32'hc2e4a507, 32'hc31f32a7, 32'hc3d9da45},
  {32'hc4af262e, 32'hc3e3bc96, 32'h43dc3d6e},
  {32'h43980a8f, 32'h4183ff5f, 32'hc4e51044},
  {32'h43d5da34, 32'hc40d4b54, 32'hc1a4ac32},
  {32'h4487d3ec, 32'hc1d5f7d9, 32'hc37443f6},
  {32'hc58a7ce5, 32'h42d20a24, 32'hc31c007a},
  {32'hc49ea72c, 32'hc3112da6, 32'hc35c0210},
  {32'hc367a864, 32'hc4bc3e9d, 32'h42175df5},
  {32'h43d9529c, 32'h44d11b3e, 32'hc38be7c9},
  {32'h44ef92fb, 32'hc39f4117, 32'hc3006762},
  {32'h44eb951b, 32'h43b8cdbb, 32'h431af32c},
  {32'hc56c549d, 32'hc1f08ca1, 32'hc3c04449},
  {32'h44fa8e7b, 32'h440a6281, 32'h43876837},
  {32'h44b61a4d, 32'hc382448a, 32'hc39d52da},
  {32'hc35788c2, 32'hc4f68658, 32'hc309b973},
  {32'hc3824bc2, 32'h42170b55, 32'h4468b7bc},
  {32'hc46e49af, 32'hc3976776, 32'hc3eb6bc8},
  {32'h445b68fd, 32'h42b1cde5, 32'h44c6d66b},
  {32'hc4a9c3eb, 32'hc1202894, 32'h42916478},
  {32'h44905ab2, 32'h4360559c, 32'h430166a6},
  {32'hc50a2ce0, 32'hc3f0c8f4, 32'hc429ba4b},
  {32'h4440b4aa, 32'h428234bb, 32'h44f2ddeb},
  {32'hc482b31d, 32'h443a48c1, 32'h43a7d4f3},
  {32'hc3822ef2, 32'hc4a5446b, 32'h446e3edd},
  {32'hc3a0fdec, 32'h4477810e, 32'hc475de8a},
  {32'hc235ca18, 32'h43dc5c4f, 32'h42e84a35},
  {32'hc3bb4949, 32'hc343ddb5, 32'hc5101d93},
  {32'h43f99568, 32'h450d9176, 32'hc3ae7957},
  {32'hc3b0a6ac, 32'h42e46f34, 32'h43322c11},
  {32'h442cc3d1, 32'h43da74e0, 32'h44ecab84},
  {32'h43e79d92, 32'hc4b8ee46, 32'hc4c2045b},
  {32'h43abdb4f, 32'h449c98ca, 32'h43b84308},
  {32'hc4803151, 32'hc47ee4a8, 32'hc41c994c},
  {32'hc3863579, 32'h45659a63, 32'h43883981},
  {32'h4263da20, 32'hc3a5f387, 32'h430ada53},
  {32'h44433ea8, 32'h43a7ceb7, 32'hc40969f3},
  {32'hc4a852b6, 32'hc41e3f97, 32'h438fe5a2},
  {32'h44720c57, 32'h44349d2b, 32'hc2b8be0a},
  {32'hc3971884, 32'h443425f7, 32'h440008bf},
  {32'hc2935cc0, 32'hc4465c9c, 32'h43c4ed26},
  {32'h43995624, 32'hc49dfcda, 32'hc3a052fc},
  {32'hc4a96626, 32'hc35e8ff3, 32'hc284f19d},
  {32'hc354c96e, 32'h4305fd90, 32'hc41087e7},
  {32'hc4d3a2e2, 32'h442417ba, 32'h4432cdd9},
  {32'h43cfd9c7, 32'hc3c791c1, 32'hc512683f},
  {32'hc5113249, 32'hc3b859fa, 32'hc27cf748},
  {32'h436ae3bd, 32'hc4508dea, 32'hc4ef5e23},
  {32'hc4c2be0f, 32'h43cebf15, 32'h4499a224},
  {32'h4441c876, 32'hc4510e9b, 32'hc30c96c5},
  {32'hc28dbf48, 32'h447378a7, 32'h4448a7f0},
  {32'h433be672, 32'hc50c3601, 32'hc43320ec},
  {32'hc3de3e30, 32'h447e7035, 32'hc3d5d9be},
  {32'h42ab247f, 32'hc42b40b4, 32'hc45145d6},
  {32'hc4992d8c, 32'h431d0d78, 32'h44b18578},
  {32'h43b357a4, 32'hc3e3e3cd, 32'hc4eca91a},
  {32'hc30f8efc, 32'h443fd832, 32'h4405964a},
  {32'hc40ab127, 32'h43051151, 32'hc3f1ae07},
  {32'h4426739c, 32'h43ddcce8, 32'hc3817aaa},
  {32'h43cfdc98, 32'hc524e451, 32'hc41a7b8a},
  {32'hc492017a, 32'h45060ec0, 32'h4395e7ac},
  {32'h449038d6, 32'h43853ce4, 32'h432b4658},
  {32'hc50e0220, 32'h44a67046, 32'h43cd4d20},
  {32'h4423c417, 32'hc4278b43, 32'hc392e338},
  {32'h4457c46e, 32'h41c9bb0a, 32'hc2c9aec2},
  {32'h4536cde3, 32'h4405e437, 32'h4400eda6},
  {32'hc5234d7e, 32'hc3d3cab9, 32'h4291eaf7},
  {32'hc455bafb, 32'h43145058, 32'hc371fe11},
  {32'hc46d82dc, 32'hc320d6a4, 32'h42e03abe},
  {32'hc41b6268, 32'hc1987ccb, 32'hc46e0f5b},
  {32'h43ce4984, 32'hc42b91bf, 32'h44a0e3f4},
  {32'hc3982536, 32'h43ef29fa, 32'hc3daabb1},
  {32'h454f7c89, 32'hc31bcefd, 32'h4300d45a},
  {32'hc4ca5b4f, 32'h43f0ab92, 32'h42c74f5d},
  {32'hc41f3689, 32'hc37670ae, 32'hc3a0ffbd},
  {32'hc46a565b, 32'h44d8f7e9, 32'h428700c4},
  {32'h4535fb60, 32'hc3c9ceab, 32'h43a3dad1},
  {32'hc48e3e37, 32'h411d87b8, 32'hc495f0bd},
  {32'h43dcef78, 32'h439bab6b, 32'h44bf1660},
  {32'hc3e36c39, 32'h4382d366, 32'hc42f2678},
  {32'h45295cf4, 32'h43548ea7, 32'hc32e2f79},
  {32'hc412c866, 32'h442a2ae9, 32'h432546a6},
  {32'h4352b444, 32'hc512f884, 32'hc403e489},
  {32'h4338e430, 32'h44395785, 32'hc392a28c},
  {32'h43a6d230, 32'hc4ab5e0d, 32'hc356b0c0},
  {32'h428a4680, 32'h4500e845, 32'h4384f908},
  {32'h451c3952, 32'hc3b1079d, 32'hc296b125},
  {32'hc5638c4a, 32'hc3a298aa, 32'hc3447162},
  {32'h44dde3bc, 32'hc3c9116c, 32'hc4667735},
  {32'h4416ef9e, 32'h44411751, 32'h43be3167},
  {32'h4491882f, 32'hc40323ba, 32'h4380cbe0},
  {32'h43897db6, 32'h452aaba5, 32'h3f0ad180},
  {32'h455d3425, 32'hc21cf7c1, 32'h43c24bc6},
  {32'hc51a87b8, 32'h44c059cb, 32'h41bc582b},
  {32'h43e5f0f2, 32'hc4f6720d, 32'hc321a243},
  {32'h44bdad58, 32'h43ff6f56, 32'hc3d5e009},
  {32'hc51d7214, 32'hc2a6e1bd, 32'h42b8adbf},
  {32'hc4838df4, 32'h4412caca, 32'hc40569ac},
  {32'hc4054df9, 32'hc49d9e2a, 32'hc29ad664},
  {32'hc3108fac, 32'h452965ba, 32'h43a41e97},
  {32'hc3487e05, 32'hc4f08154, 32'hc43027b3},
  {32'h444da51d, 32'h44d5a6d8, 32'h43b8638a},
  {32'hc4c1e22c, 32'hc4755286, 32'h43daf763},
  {32'h452103c4, 32'h42fad6af, 32'h43e531ae},
  {32'hc448f47a, 32'hc3fad23c, 32'hc3aa966e},
  {32'h4480bed4, 32'hc42b4cfc, 32'h43ba21c9},
  {32'h4415e66a, 32'h42cc97b8, 32'h44344fce},
  {32'h44307a61, 32'h441e01d5, 32'hc1873185},
  {32'h41e649c0, 32'hc467b694, 32'hc2d49639},
  {32'hc39a812c, 32'h44fff716, 32'h432823ac},
  {32'hc444ba28, 32'hc406bffc, 32'h43d37953},
  {32'h45051c6a, 32'h442df0d1, 32'h43051064},
  {32'h44bd9252, 32'hc429d5f2, 32'hc411daca},
  {32'h45172083, 32'hc3ef6eaa, 32'h43c46ae0},
  {32'hc41fa14c, 32'h43a2f9bc, 32'hc497c39d},
  {32'hc4d2bd88, 32'hc3872be5, 32'hc32065d7},
  {32'hc05f9400, 32'hc52b3b70, 32'hc338f42a},
  {32'h43fd10de, 32'h441eeb0b, 32'h4475aa5c},
  {32'hc3dfd45b, 32'hc3e4ffda, 32'h434bbae4},
  {32'h44167cb3, 32'h44b38d61, 32'h43817dea},
  {32'hc4354554, 32'hc4bec934, 32'hc417466a},
  {32'hc4267ec6, 32'h445fc697, 32'hc2463497},
  {32'h4527b0c8, 32'hc32c298e, 32'hc3717f23},
  {32'hc4ab8915, 32'h425eec5d, 32'hc4439e31},
  {32'h42835d83, 32'h454ce928, 32'h443c945e},
  {32'h432a61fa, 32'hc41d3f2b, 32'h43107565},
  {32'h427a6786, 32'h443c4adc, 32'h4384b3e9},
  {32'hc4348e6a, 32'hc53f8b71, 32'hc1c71f6c},
  {32'h44f9122a, 32'h438597c6, 32'hc41bd545},
  {32'hc58ebe74, 32'h438652df, 32'hc4008554},
  {32'h442776da, 32'h430f4431, 32'h43f47310},
  {32'h4463c804, 32'hc42a8425, 32'h43148d8a},
  {32'h430446b0, 32'h45114e90, 32'hc19bffa8},
  {32'hc492be20, 32'hc2a6e75d, 32'h4240f27d},
  {32'h448186c7, 32'h44549c5f, 32'hc32d6130},
  {32'hc46180fe, 32'hc48e743b, 32'h4327532a},
  {32'h441da630, 32'hc2ca1283, 32'hc4991857},
  {32'hc4a4aae3, 32'hc1e3d8ce, 32'hc1bf6605},
  {32'hc1b9cfc4, 32'hc32f3442, 32'hc53847b4},
  {32'hc2e7f1a6, 32'h43fa8ecc, 32'h454b81be},
  {32'hc25373c0, 32'h4451551a, 32'hc3100d68},
  {32'hc4c79ea0, 32'hc4b0ad9b, 32'h448e01e9},
  {32'h440afc16, 32'h44d91310, 32'hc42c1a9d},
  {32'h44ad85a2, 32'h420e9fa0, 32'h439ee1e8},
  {32'h44204c58, 32'h42f39799, 32'hc532965b},
  {32'hc40ef491, 32'hc2fb4bc4, 32'h42c2ad62},
  {32'h4516ce06, 32'h4194e6ac, 32'hc3a8eb7b},
  {32'hc4d19bc7, 32'hc346950a, 32'h43d5faf1},
  {32'h43dd9962, 32'hc3707857, 32'hc483bca1},
  {32'h431992c0, 32'hc51c86fe, 32'hc34adc60},
  {32'hc4149e1c, 32'h4492b893, 32'h40b94bb4},
  {32'hc32ff52c, 32'hc2765636, 32'h442e778f},
  {32'hc5375dc6, 32'h43cb07cd, 32'hc4603e17},
  {32'h43a5f5db, 32'hc4e685ea, 32'hc33c9fa9},
  {32'h44885cb4, 32'h438e2d16, 32'h4390af26},
  {32'h4506b451, 32'hc2def2a7, 32'hc44cd5a2},
  {32'hc5331135, 32'h43f2ef52, 32'h441fb80d},
  {32'h44a68087, 32'h43bc41e8, 32'h43e41d79},
  {32'hc3925c24, 32'h443dfa92, 32'hc38f8bd8},
  {32'h42dd9c14, 32'hc5354d25, 32'hc307e820},
  {32'h4404083d, 32'hc388ec64, 32'hc25a34e6},
  {32'h4529e111, 32'hc328dd2c, 32'h43b74fa6},
  {32'hc367bf7c, 32'h423228a8, 32'hc5124e8e},
  {32'hc30b9146, 32'hc480cfbf, 32'hc2fcf01e},
  {32'hc5307736, 32'h40dec8d4, 32'h42ebf26b},
  {32'h4431a214, 32'hc4645532, 32'h44025ceb},
  {32'h44f54b95, 32'h4401ba67, 32'hc40ebdee},
  {32'hc1734800, 32'hc50fd692, 32'h43a0576a},
  {32'hc4fdc882, 32'h43f59fbf, 32'hc3726171},
  {32'h438fcd03, 32'hc25ac492, 32'h433089f9},
  {32'hc44222c5, 32'hc2d90119, 32'hc54f58df},
  {32'h43b51d20, 32'hc492a86c, 32'h449db6b6},
  {32'hc4c3858f, 32'h43e986e0, 32'hc4090242},
  {32'hc382f880, 32'h444a3d76, 32'h44cb6f63},
  {32'hc579b56e, 32'h42d88270, 32'hc2e61b99},
  {32'h454c94be, 32'hc3cf5b76, 32'hc32cfdf4},
  {32'hc24bb54a, 32'h443cc50a, 32'hc4ad9683},
  {32'h44880ba1, 32'h444cbbb8, 32'h440710ce},
  {32'h44ec4aac, 32'hc35c88e1, 32'hc3983186},
  {32'h44a4cf9a, 32'hc2b0f5fc, 32'hc0cf0274},
  {32'h43b27b38, 32'h430983a2, 32'h450fa841},
  {32'hc32b4818, 32'hc388e339, 32'hc458e505},
  {32'hc060ed40, 32'hc4dd5b49, 32'h4391929c},
  {32'hc4c78830, 32'h42684dca, 32'hc496fb5d},
  {32'hc40635f6, 32'h430ad6b5, 32'h452b1400},
  {32'h44a13373, 32'hc48187ae, 32'h44da44bd},
  {32'h433c8a65, 32'hc50fd555, 32'hc4af1a95},
  {32'hc215d353, 32'hc4bae17c, 32'h44337959},
  {32'h4387f4aa, 32'hc3ce1a84, 32'h431355fc},
  {32'h438127d8, 32'h44195c83, 32'hc389c7e7},
  {32'h43b0e08e, 32'hc4d7ffa7, 32'hc3ce9598},
  {32'hc3839a62, 32'h443527c7, 32'hc414401f},
  {32'h44f70d5a, 32'hc365099a, 32'h441bce7d},
  {32'hc3ad7102, 32'hc4598caf, 32'hc4e842b7},
  {32'hc3e715da, 32'h4391a11b, 32'h442b465f},
  {32'hc58a51cc, 32'hc3e753ab, 32'hc34f1519},
  {32'h452ffd19, 32'h43a396eb, 32'h44400a4f},
  {32'hc4cf96b2, 32'hc38ad282, 32'hc216014d},
  {32'h43786f62, 32'hc55da3c9, 32'hc182035a},
  {32'hc31d75e4, 32'h4525f617, 32'h43b738a7},
  {32'h4523320a, 32'hc375a101, 32'hc36f9c1d},
  {32'hc50bcb22, 32'h4490db9e, 32'h43879140},
  {32'h43945494, 32'hc544e671, 32'h43776d1d},
  {32'h449d155d, 32'h4311c81a, 32'h431a1f83},
  {32'hc3875d1a, 32'h44351ac0, 32'hc52de8e7},
  {32'h43ebafe9, 32'h435ef94e, 32'h4527952d},
  {32'hc43ed08b, 32'h43adf3be, 32'h44b3cacc},
  {32'h438b6770, 32'h4452911f, 32'hc44f3727},
  {32'hc3a759da, 32'hc41cc2d0, 32'h43ca5aa6},
  {32'h442b302c, 32'h43d799e6, 32'hc40c89ae},
  {32'hc5097490, 32'hc20ab988, 32'h446274e1},
  {32'hc33ec1c0, 32'h44a10f83, 32'h425c3b3b},
  {32'h44c1d7fa, 32'h4222fba8, 32'h43f345b3},
  {32'h4261d3e8, 32'h4457f935, 32'h44f14004},
  {32'hc224e574, 32'h414de57a, 32'hc545239a},
  {32'h448a5eba, 32'h44637329, 32'hc3790740},
  {32'hc44a8dec, 32'hc3317ae5, 32'h451b398d},
  {32'h43efa6b5, 32'h43ef4c06, 32'hc3efbd73},
  {32'hc48e302c, 32'hc48f1be4, 32'h4429d18e},
  {32'h447668ea, 32'h43d76c79, 32'hc308d58c},
  {32'h4472879e, 32'hc2a8a74a, 32'h44093eea},
  {32'h438743a4, 32'hc41b95e0, 32'hc349505f},
  {32'hc5891f60, 32'h42e047ea, 32'h426d2e34},
  {32'hc41c1a8b, 32'h42c1325a, 32'hc2e43e16},
  {32'h43418f07, 32'hc584af40, 32'h43410b2b},
  {32'h44bdf759, 32'h4428758a, 32'hc2e12ace},
  {32'h44e4ab81, 32'hc171303a, 32'h436dd894},
  {32'h4308e57c, 32'h456761a3, 32'hc2f3de7b},
  {32'hc4786874, 32'hc4c6e07b, 32'h43c60bf0},
  {32'h45145063, 32'h41f99518, 32'hc3967308},
  {32'h414d7b94, 32'h44b3ec90, 32'hc2806ca2},
  {32'h4402953c, 32'h44c0328b, 32'hc4b99b63},
  {32'h4300055f, 32'hc487f0bc, 32'h448a3102},
  {32'h42cb4b9c, 32'hc38a0298, 32'hc2249c96},
  {32'hc31b7c08, 32'h441f707c, 32'h4499bfe3},
  {32'hc4b4b679, 32'hc38bd92d, 32'h43eaa9f7},
  {32'h440460fc, 32'h43fd56e6, 32'h40e6a034},
  {32'hc3e87836, 32'hc4c50325, 32'hc4dfbf10},
  {32'h4484aab1, 32'h43954eca, 32'h44035a7b},
  {32'h44408ff4, 32'h44a95d9c, 32'hc40811ac},
  {32'h43f83294, 32'hc447da35, 32'h4480ae1a},
  {32'hc45e8f59, 32'hc2970f4b, 32'hc41df034},
  {32'hc3c433a8, 32'h437564ea, 32'h44a06bf4},
  {32'hc4d4accb, 32'hc3ca209e, 32'h42c68ea2},
  {32'h43bf46d9, 32'h430ed4a1, 32'h44ec5a0b},
  {32'h447c7d70, 32'h433c3158, 32'hc489352b},
  {32'hc36a837a, 32'h449224af, 32'h4534257b},
  {32'hc4265944, 32'hc3515f10, 32'hc4fd7cca},
  {32'h44d51e09, 32'h42199b45, 32'hc1b0cdf7},
  {32'hc535e35e, 32'hc42fc358, 32'h41e51ec3},
  {32'h44669a74, 32'h448125d2, 32'h44382236},
  {32'hc30c1100, 32'hc3e3a4a7, 32'hc36e98e6},
  {32'h452ebc24, 32'h43e31a74, 32'h41823e0a},
  {32'hc41c9950, 32'hc481a609, 32'h3fce66a0},
  {32'h454b2198, 32'h433a204c, 32'h4400811a},
  {32'hc5434e61, 32'hc18d11b4, 32'h432101f9},
  {32'h4579901c, 32'hc2939f92, 32'h42a0928a},
  {32'h44351eb9, 32'h421e8834, 32'hc3e0bf7c},
  {32'h439277d6, 32'h4387463d, 32'h449468a8},
  {32'h43fa9512, 32'hc39a3282, 32'h43eee038},
  {32'hc363d0b0, 32'h4523abc2, 32'hc1c2bd56},
  {32'hc3598608, 32'hc3cb0516, 32'hc4f66df0},
  {32'h418bd3d1, 32'h44239b9b, 32'h44f9dec7},
  {32'h444d98b6, 32'h42931c17, 32'hc487e0fc},
  {32'hc55a3b26, 32'h4339d31d, 32'h43e4fb30},
  {32'hc36d8f66, 32'hc452a5f8, 32'hc4ade878},
  {32'h4342d888, 32'h451decfc, 32'h441e066c},
  {32'hc3c2fe72, 32'hc50ed858, 32'hc47cefc1},
  {32'hc4b7bf6f, 32'hc32af62f, 32'h43413062},
  {32'h4472c488, 32'hc4a32af7, 32'hc3dcfc36},
  {32'hc4d40c25, 32'h4447ac06, 32'h4386e8c3},
  {32'h44a1301c, 32'h43814db5, 32'hc31fb152},
  {32'hc5386bc8, 32'hc2b98009, 32'h43960191},
  {32'h4329dd3a, 32'hc3704f0f, 32'hc4a9d4c4},
  {32'h445a6f89, 32'h434a7e20, 32'h43ac4c50},
  {32'h44a043bd, 32'hc4af76f2, 32'hc37758ae},
  {32'hc47669c4, 32'h44dfd1ee, 32'h437265da},
  {32'h4527b3c5, 32'h43d23c14, 32'h43027cd8},
  {32'hc48d1762, 32'h4502c0fb, 32'h43e7a358},
  {32'h41beeb63, 32'hc53e9e8b, 32'h434dd7f2},
  {32'hc536b922, 32'hc3c91f2e, 32'h40837430},
  {32'h4408aaee, 32'h438ccf82, 32'h4249405e},
  {32'hc580adac, 32'h43a1e269, 32'h43bb1bdf},
  {32'hc4537866, 32'hc20ddfb2, 32'hc403473c},
  {32'h4489faf2, 32'h43a7a59d, 32'h4412a8e1},
  {32'hc4b2dfd4, 32'h430c309b, 32'hc46dbd1f},
  {32'h4533f5ea, 32'h4328b45d, 32'h439d470e},
  {32'hc4656c17, 32'hc1eadaed, 32'hc24dfc04},
  {32'hc2adcb80, 32'hc53e7cb0, 32'hc22cde02},
  {32'hc3c68eb6, 32'h434ef302, 32'h432de5a4},
  {32'h450ed67d, 32'h440a3958, 32'h4368af83},
  {32'hc4c9cccd, 32'h44a8d0a9, 32'h4222ffc2},
  {32'hc1999000, 32'hc571ad71, 32'h439c94a4},
  {32'hc5327c1d, 32'h4365e848, 32'hc30cd0cc},
  {32'h43f3c680, 32'hc2588c55, 32'h444f8ccf},
  {32'hc451c790, 32'h4379fd5f, 32'hc445e484},
  {32'h455309c4, 32'h434b9f9f, 32'hc20df641},
  {32'hc46ccf4e, 32'h4350032c, 32'h443dadc6},
  {32'hc3c4d109, 32'hc4917d4f, 32'hc4b9509b},
  {32'h4446a246, 32'hc3644cfd, 32'h430f32dc},
  {32'hc3915a48, 32'hc49a0d70, 32'hc3d8d31b},
  {32'h42ea6050, 32'h453984dd, 32'hc37b24a1},
  {32'hc4887e06, 32'hc4099136, 32'h42f655b8},
  {32'hc41bf844, 32'h42b40d1d, 32'h43b1b462},
  {32'h45131c81, 32'h438ff318, 32'hc47f44ce},
  {32'h439b2e16, 32'h449c9a6c, 32'h43950366},
  {32'h4230b418, 32'hc52ec0fe, 32'h41441fb0},
  {32'hc4e3a7c2, 32'h4361237f, 32'h43fed5f1},
  {32'h449b4688, 32'hc416fa71, 32'hc3a38ae5},
  {32'hc512c410, 32'h44ba03d9, 32'h43795ace},
  {32'h4327cacc, 32'hc429ddb9, 32'hc5513227},
  {32'hc3047160, 32'hc35b4c1d, 32'hc440ae0c},
  {32'hc5042f45, 32'h43305720, 32'h44c3bf12},
  {32'h44f090e9, 32'h43819a84, 32'hc3c99ef3},
  {32'hc33697ea, 32'hc50c64ed, 32'hc3e32e44},
  {32'h4551fb25, 32'hc3d1d709, 32'h43c46c7c},
  {32'h442f6247, 32'hc3bd4c4b, 32'hc335285a},
  {32'h43588230, 32'h450b57f8, 32'h4405785c},
  {32'hc4a4eb5c, 32'hc50b5dc5, 32'h42b9deb4},
  {32'hc3f43410, 32'h44c09429, 32'h436cae3e},
  {32'hc4643e30, 32'hc32e714d, 32'h4506f1ac},
  {32'h445b80a5, 32'h43263a27, 32'hc44f2d12},
  {32'hc3a61ad0, 32'h4218e429, 32'h42cadf54},
  {32'h44bef81b, 32'hc3b4e9ef, 32'h43a08c0b},
  {32'hc424eb1c, 32'hc4d0a516, 32'hc436f788},
  {32'h43226baa, 32'h431c56a1, 32'h44ec82be},
  {32'hc4c04a78, 32'hc46e7370, 32'h4283295a},
  {32'h44b6a1c0, 32'h43ce2e63, 32'h43bb4221},
  {32'hc3bf6337, 32'hc4478a66, 32'hc4759e8d},
  {32'h44af4a26, 32'h4458afc3, 32'h4402a0ce},
  {32'hc5034053, 32'h4426c7b9, 32'hc47e6ab2},
  {32'hc44bdf18, 32'h42f415cd, 32'hc342c313},
  {32'h42366240, 32'hc43886c5, 32'hc501132b},
  {32'h45176545, 32'h43f885dd, 32'h43c680ec},
  {32'hc3ab1fd4, 32'hc445237f, 32'hc32b8fae},
  {32'h441b66b2, 32'h449b21a2, 32'h448c1c2c},
  {32'hc3bcee5a, 32'hc50d1ddf, 32'hc428725a},
  {32'h450986ee, 32'h439c7fcb, 32'h42c9f4a2},
  {32'h451e359e, 32'hc42931c6, 32'hc3673dc4},
  {32'hc4a88c3c, 32'hc45944c9, 32'h43ca6603},
  {32'h441dce5a, 32'h44014080, 32'h4411d0b2},
  {32'h428e233c, 32'hc4971753, 32'h43508cf4},
  {32'h437cf7d0, 32'h444eb514, 32'h4449c9f6},
  {32'hc420c172, 32'hc3b503f3, 32'h443eb7bf},
  {32'h452ee5a8, 32'hc3976278, 32'hc4062a29},
  {32'hc4ed1bae, 32'hc3f35428, 32'h434f78b0},
  {32'h456ee8e0, 32'h440918e4, 32'h445148ed},
  {32'hc36ea0ec, 32'hc47ba8f2, 32'h44997d41},
  {32'h43b7ca31, 32'h43d4dd5a, 32'hc46e7539},
  {32'hc38820d8, 32'hc405b7b8, 32'h44b62fe2},
  {32'h42606ac8, 32'h444db9ae, 32'hc2edb888},
  {32'hc399dbb0, 32'hc4a0d1f2, 32'h442f1705},
  {32'h444d091d, 32'h4412a930, 32'hc506c4c0},
  {32'h43fbc739, 32'hc3611c79, 32'h44bb0caa},
  {32'h449d33d4, 32'h43384955, 32'hc42033ab},
  {32'hc44453f2, 32'h43738d1e, 32'h4475ba94},
  {32'h4488285e, 32'h446dba1a, 32'hc3b108e2},
  {32'hc4461a15, 32'hc5145ad7, 32'h433d7d11},
  {32'h4401ced6, 32'h444b5e6d, 32'hc48fa254},
  {32'hc4cab0a4, 32'hc3a13779, 32'hc13e9e04},
  {32'h44f32d8d, 32'h43104cca, 32'hc44bf892},
  {32'h43da5034, 32'h434a6584, 32'h451ed1f1},
  {32'h4528baae, 32'h43a253b4, 32'hc37e7e81},
  {32'hc48c2b16, 32'h4313c557, 32'h44ccf8c8},
  {32'h45636411, 32'hc4267e77, 32'hc47a1dc0},
  {32'h44702049, 32'hc474a53e, 32'hc39008ce},
  {32'hc4949d5f, 32'h4311b57e, 32'h422128fc},
  {32'h452c67f5, 32'h440e1eb4, 32'h43db536b},
  {32'hc3af9260, 32'h43805556, 32'h43160c52},
  {32'h43feedc8, 32'hc4b01ed8, 32'h44131f49},
  {32'h44819902, 32'h4438898b, 32'h412f9bf9},
  {32'h4556d7e7, 32'h4297ed04, 32'h4309944b},
  {32'hc54f0e12, 32'h43c61de4, 32'h43af2bec},
  {32'hc4d2a932, 32'h42e214f7, 32'h4290ca5c},
  {32'hc3523f98, 32'h43a975ae, 32'h4416b4a9},
  {32'h44900a9e, 32'hc44dde25, 32'hc213d69e},
  {32'hc49ac42e, 32'h437382e6, 32'hc2d7e12a},
  {32'h44c038bf, 32'hc3e46bf6, 32'hc15c2160},
  {32'hc4552c30, 32'h449759f5, 32'hc4268ee1},
  {32'h43fc65ba, 32'hc457608d, 32'h428c4bbb},
  {32'hc3bf1df0, 32'hc39534c8, 32'hc4dbf106},
  {32'h454dffaf, 32'h440c3513, 32'hc3fe1118},
  {32'h44984be0, 32'h439c4ff2, 32'h440da9b2},
  {32'h43a8af42, 32'hc48f8038, 32'h44235533},
  {32'hc52f748f, 32'h4392b3ec, 32'hc2369600},
  {32'h4560e545, 32'h43e30629, 32'h43264dee},
  {32'hc37d2ea0, 32'h44108ab6, 32'hc41d6a91},
  {32'h44851a4a, 32'hc4519719, 32'hc3e013c5},
  {32'h44b870dd, 32'hc2a0450d, 32'hc248ccac},
  {32'h43f11a32, 32'h42ca3e8e, 32'h44f8d80d},
  {32'hc4ee26fc, 32'hc40adf19, 32'hc4c0a8db},
  {32'h450d3277, 32'hc2b537c7, 32'h43c33b30},
  {32'h416b34a0, 32'h44b5d77b, 32'hc4e05f03},
  {32'h4383b216, 32'hc4a2b3e7, 32'h443bb606},
  {32'h44324196, 32'h42282064, 32'hc43184d3},
  {32'h44c7acb9, 32'h43b6a58c, 32'hc35b879c},
  {32'h448e142a, 32'hc4b754af, 32'h4411964c},
  {32'h42f681f0, 32'h4383bb5e, 32'hc5018370},
  {32'h44018bad, 32'h43d8a790, 32'h44ecee8b},
  {32'h42cf436a, 32'h4543a0d7, 32'h43e8876d},
  {32'h4143ca80, 32'hc4203867, 32'h44ea7651},
  {32'h45021664, 32'hc2b08004, 32'h449d1700},
  {32'hc2606650, 32'h44875fe7, 32'hc4d32655},
  {32'h4462eb3f, 32'hc41e4f18, 32'h443eca06},
  {32'hc403b33c, 32'h43260175, 32'h442c9d67},
  {32'hc38a1faf, 32'hc2b7598b, 32'hc4c9cbd0},
  {32'hc3850436, 32'hc4db831a, 32'hc1859538},
  {32'hc3371c61, 32'h43fd8575, 32'hc4a29198},
  {32'h450f3067, 32'h4323ab76, 32'h43f6e7df},
  {32'hc3cd0cfc, 32'h444daa40, 32'hc4ca8fa4},
  {32'hc44c667c, 32'hc3beee2a, 32'h43859691},
  {32'hc578e496, 32'hc315cb1c, 32'hc3a6f94b},
  {32'hc380a27c, 32'hc2d58ab1, 32'h434047a8},
  {32'h418e6859, 32'h44306d30, 32'h41d844f9},
  {32'h448e647a, 32'hc4f58107, 32'hc3a92284},
  {32'hc458bb67, 32'h44a103b7, 32'hc3d0661d},
  {32'h445fe53f, 32'hc4b3f315, 32'h42b34536},
  {32'hc36254a0, 32'h44e639cb, 32'hc37bee00},
  {32'h44317390, 32'hc4abaf17, 32'hc420ba8b},
  {32'hc3dc3834, 32'h442c9603, 32'h44335ed5},
  {32'hc33a1ce8, 32'h450b96ef, 32'hc4e68f3e},
  {32'h42a20bb9, 32'h439415e7, 32'h44964379},
  {32'h4307cb98, 32'hc54255b4, 32'h3ffce530},
  {32'h4330d250, 32'h44c719f0, 32'hc1c01d7a},
  {32'hc333ea70, 32'hc416561c, 32'h430d6028},
  {32'h439e4f8d, 32'h43dfd02a, 32'hc453232f},
  {32'hc4716d8c, 32'hc4980bff, 32'h43c749d0},
  {32'h4337b256, 32'h433c5ac8, 32'hc3e72b96},
  {32'hc34419cf, 32'h442d5ecd, 32'h435631d1},
  {32'h43958644, 32'h43971b6d, 32'h455c7ad8},
  {32'hc36e05fe, 32'h43abd501, 32'hc51d539f},
  {32'h4489dc04, 32'h4483bcf6, 32'h43116200},
  {32'h41f18320, 32'hc493caf6, 32'h43426b16},
  {32'h449a3678, 32'h4408c4dc, 32'hc318b841},
  {32'hc40f8ca2, 32'hc4dfedee, 32'hc3b9140c},
  {32'h43cd6298, 32'h441300d4, 32'hc319ce2a},
  {32'hc4ded97c, 32'hc3d7fc16, 32'h431fdb50},
  {32'h457cf59e, 32'hc345ab13, 32'h4288de7b},
  {32'hc4983649, 32'hc29afab7, 32'h44023814},
  {32'hc49d0f6b, 32'h438a8715, 32'hc38c5a18},
  {32'hc4bfc515, 32'hc4da9b9e, 32'hc2527689},
  {32'h456234d5, 32'hc1d09c38, 32'h43bae9eb},
  {32'h43bf1cc0, 32'hc4994ad4, 32'h430bd23e},
  {32'h430d6d78, 32'h457a884c, 32'h42ff4aab},
  {32'hc52c81e6, 32'hc4024eb1, 32'h43a6414c},
  {32'h44f1ba2c, 32'h43210e6a, 32'hc42e6613},
  {32'h4427d73c, 32'hc49410b8, 32'h449b0c9c},
  {32'hc3161b36, 32'hc30656a5, 32'hc49cd8f7},
  {32'hc40bed0c, 32'hc0c96552, 32'hc397874e},
  {32'hc44cb99a, 32'h43ff6c0b, 32'hc27b90a1},
  {32'h453d1f32, 32'hc309b05f, 32'h442346ea},
  {32'h44335b82, 32'hc21c0ff1, 32'hc5209fe3},
  {32'h45433fdd, 32'hc35f9992, 32'hc396e99b},
  {32'hc5478ce7, 32'hc156bd6b, 32'hc30ceb19},
  {32'hc34657e2, 32'h44914eec, 32'h451b5a36},
  {32'h442e63ec, 32'h4478d167, 32'hc41d2867},
  {32'h4486c82e, 32'h433f7594, 32'h4285f258},
  {32'hc418c70a, 32'hc38b65b8, 32'hc4c012c7},
  {32'h42beb360, 32'hc302a403, 32'h4407e21a},
  {32'hc42e708b, 32'hc3ccdf28, 32'hc49d75b7},
  {32'h44348078, 32'h4472e102, 32'h43be626d},
  {32'hc370637c, 32'h421d0811, 32'hc26523e4},
  {32'h42acba2a, 32'h424b8acd, 32'h44894a37},
  {32'hc4729e49, 32'hc3ab497e, 32'hc4f04c5d},
  {32'h447fcbc3, 32'h44389524, 32'h434dd61e},
  {32'hc4f8c6d0, 32'hc488d1b9, 32'h42ad626a},
  {32'h44c05ee5, 32'h44802f5f, 32'h42530afe},
  {32'h4423db51, 32'hc3ecddc7, 32'hc2a6b211},
  {32'h443bfec8, 32'h44aba179, 32'hc33ecef5},
  {32'hc49440e3, 32'hc49271b5, 32'h43e2a826},
  {32'hc44c418c, 32'h43e66101, 32'hc2321adc},
  {32'hc52a5302, 32'h4423cd25, 32'hc44e50d7},
  {32'h43e24340, 32'h43b0429a, 32'hc3c94fbe},
  {32'h445beee6, 32'h4436ca94, 32'hc496509a},
  {32'hc37b0348, 32'hc2892184, 32'h449ad026},
  {32'h43be312d, 32'h43a6d66a, 32'hc3bd9e5e},
  {32'hc3a6e5e8, 32'h44251dbe, 32'h44e128f6},
  {32'hc3ecba84, 32'hc3b8afd7, 32'hc548fca3},
  {32'h4281eaf0, 32'h4376ca14, 32'hc27087e3},
  {32'h43c146be, 32'hc4d2778b, 32'hc4b7036c},
  {32'hc570e38d, 32'h438fbf4f, 32'hc3277ed0},
  {32'h43dac42c, 32'h43a2e635, 32'hc4a45a3f},
  {32'h44183b0f, 32'hc48239df, 32'h4501b9dd},
  {32'hc3715566, 32'h450c0abe, 32'hc515bd93},
  {32'h434c70d8, 32'hc469a162, 32'h442e033f},
  {32'h4365f4ce, 32'hc3dc125a, 32'hc51fae46},
  {32'hc513de25, 32'h43d1e181, 32'hc252b090},
  {32'hc406ef8c, 32'hc408e4ac, 32'hc44ad4c8},
  {32'hc4b0519e, 32'hc199ce1c, 32'h449df62a},
  {32'h44a7b998, 32'hc4174dd9, 32'hc493b75f},
  {32'h44f03954, 32'hc2ecfa72, 32'h4349b684},
  {32'h44c6b848, 32'hc4b3d556, 32'h429b367f},
  {32'hc555ab7c, 32'h4416eb7a, 32'h42d4df9e},
  {32'h43f8340d, 32'hc33b04cc, 32'hc3eace35},
  {32'hc33fe9c0, 32'hc298a991, 32'h4328d8f7},
  {32'h444e83d8, 32'hc4d26375, 32'hc3b10e79},
  {32'h4447eabb, 32'h43c4e9e8, 32'h4378e154},
  {32'h450ccc16, 32'hc18f0c99, 32'h436f505f},
  {32'hc5399745, 32'hc2bd510f, 32'h43cf42b7},
  {32'h445bcd77, 32'hc438d319, 32'hc32a75b1},
  {32'hc3e970d3, 32'hc3e68545, 32'hc36c9c96},
  {32'hc40f818a, 32'hc3009ed1, 32'hc51bba8e},
  {32'h45318680, 32'h42a90dd0, 32'h4365f763},
  {32'hc3da3880, 32'hc2ab632e, 32'hc0393aa6},
  {32'h44734e6b, 32'hc483ad58, 32'h411f3b33},
  {32'h42ec3586, 32'h4547c2f7, 32'h4388c881},
  {32'hc3eee8d2, 32'hc4925d9c, 32'hbf1b9a00},
  {32'hc56607a5, 32'h43bb1bf3, 32'hc254b4bb},
  {32'h44934dff, 32'hc49e56a9, 32'hc40372a6},
  {32'h44a901ee, 32'h4453073e, 32'h432e692f},
  {32'h44a95e2d, 32'h4369bdf6, 32'hc2b95995},
  {32'hc514d8b8, 32'h43e5efd6, 32'h42a5eef4},
  {32'h42b85d4a, 32'hc4999fd1, 32'hc0aa8348},
  {32'h44354e07, 32'h4441e84d, 32'h44dee7e9},
  {32'h43c28e13, 32'hc47cf012, 32'hc4619827},
  {32'hc32f6ff8, 32'h43c4b82e, 32'h4398859c},
  {32'h43f54c6f, 32'hc4709ea0, 32'hc3514052},
  {32'hc4ad97ca, 32'h4385bc9d, 32'h4438083c},
  {32'hc49ee77c, 32'hc2ac5346, 32'hc374d5c1},
  {32'hc499c190, 32'hc2364b87, 32'h44865e8f},
  {32'h4529d82c, 32'hc3c329ef, 32'hc42a8bb3},
  {32'hc4b4b38c, 32'hc33987b5, 32'hc058861c},
  {32'hc3eb9c98, 32'hc4a4dcac, 32'hc3c48013},
  {32'hc5113284, 32'h43b296a0, 32'h437f336a},
  {32'h44e26072, 32'hc2c3fd0a, 32'hc3a93085},
  {32'hc51d2a8c, 32'hc297567d, 32'h43b9f729},
  {32'h43e53678, 32'hc4fac885, 32'hc32e316f},
  {32'h4553c025, 32'h43061587, 32'hc459fc4d},
  {32'hc506bf3a, 32'h4219247c, 32'h4434734a},
  {32'h4388995f, 32'hc4522dfa, 32'hc4a3e719},
  {32'hc4e33bbb, 32'hc4969bcb, 32'h41345a6f},
  {32'h44e88c8a, 32'h4404de96, 32'h4364f51d},
  {32'h41860c78, 32'hc51530f1, 32'hc3bd41c9},
  {32'h442331c2, 32'h450b1938, 32'h43d755c1},
  {32'hc2370f4c, 32'hc4ee39ae, 32'hc346b29a},
  {32'h44ce45f9, 32'hc2f66d09, 32'h43720aef},
  {32'hc42993d8, 32'h43ba84a1, 32'h445b07a2},
  {32'h43b18bd2, 32'hc40f9a9e, 32'h44165624},
  {32'h439ef3eb, 32'hc27aa037, 32'h4357d01b},
  {32'h4376b492, 32'h43ed34c7, 32'h43d88202},
  {32'hc4a9dc26, 32'hc4801ac0, 32'hc4af8e75},
  {32'h42dafa80, 32'h4386b022, 32'h449dd896},
  {32'h42de3138, 32'hc4b29b5d, 32'hc4691609},
  {32'h449ac7b8, 32'h441846a9, 32'h443091ac},
  {32'hc385c60a, 32'hc4afef6e, 32'hc3f05f76},
  {32'h42e9ccc0, 32'h430dbf61, 32'hc307a291},
  {32'hc4f17422, 32'hc269e5c5, 32'h41ad7611},
  {32'h451434f4, 32'h4293ca62, 32'hc4020264},
  {32'h4421f771, 32'hc4e32a6f, 32'hc26cc796},
  {32'h43aca46d, 32'h42cb66cd, 32'h44ce309d},
  {32'hc184a730, 32'hc4ce2671, 32'hc381309b},
  {32'h4311f5c0, 32'h4515fa07, 32'h43d4d9a3},
  {32'hc2ba1768, 32'hc4a3f87c, 32'hc4e2bf62},
  {32'h4329e352, 32'hc3519c48, 32'h446720ad},
  {32'h44252ec4, 32'h44d7175e, 32'hc3dedbb5},
  {32'hc45f92cc, 32'h42054df9, 32'hc4c201ec},
  {32'h44addaf6, 32'h447b6078, 32'h43af1db4},
  {32'h44f80659, 32'h42d81334, 32'h430c5267},
  {32'h4528fd78, 32'h43602125, 32'hc3711ca7},
  {32'hc4805068, 32'hc43c8217, 32'hc37ded34},
  {32'hc4f8b179, 32'h42a3cb60, 32'h430f389e},
  {32'hc3b501e0, 32'h43285173, 32'hc39e59bb},
  {32'h44468fe4, 32'hc2123cbd, 32'hc2e6de29},
  {32'hc36ac8c9, 32'hc2bd1117, 32'h44336844},
  {32'h44c5aba0, 32'h442c991f, 32'hc325f602},
  {32'hc505213c, 32'hc350bacd, 32'h442259b1},
  {32'hc4acbf4b, 32'h44012a4a, 32'h43232662},
  {32'h40f79ab4, 32'hc48afb80, 32'h445c77b9},
  {32'h4367dbdb, 32'h4521a782, 32'hc190da14},
  {32'h44997734, 32'h4218d517, 32'h43313722},
  {32'h44ae034b, 32'hc2980d79, 32'hc49c287b},
  {32'hc4d11e71, 32'hc21a346a, 32'h4389c06f},
  {32'hc3021bbc, 32'h434002d8, 32'hc41268eb},
  {32'hc1893e90, 32'hc490d21f, 32'h4402f6c7},
  {32'hc3d89920, 32'h4480929e, 32'hc4c19477},
  {32'hc537a576, 32'h43c824e1, 32'hc082e9cc},
  {32'h4317f19a, 32'h440f45a3, 32'hc4931652},
  {32'hc3880151, 32'hc2bd557d, 32'h450ab2c2},
  {32'h4496540e, 32'h43d231f9, 32'hc3c78f2c},
  {32'hc4b9f2f4, 32'hc20d394f, 32'h434c3697},
  {32'h452251e6, 32'h43f5aaab, 32'hc4017916},
  {32'h450ed070, 32'hc43780bd, 32'h414076a5},
  {32'hc42ffac9, 32'h44c04e73, 32'h429ca7d9},
  {32'h4502fcbd, 32'h43848695, 32'h432c8854},
  {32'h42fca03a, 32'h457d221b, 32'hc338282c},
  {32'h4437853c, 32'hc3b1a323, 32'hc351953b},
  {32'hc506ee0e, 32'hc33dcf15, 32'hc2ca7661},
  {32'h44a942f6, 32'hc436413c, 32'h439e5e2e},
  {32'hc536acaa, 32'h44488fab, 32'h43e4cffb},
  {32'h44d3d96f, 32'hc444450d, 32'hc3248c31},
  {32'h42dedff0, 32'h442f755f, 32'hc508439a},
  {32'hc40cfcd7, 32'hc51bba5c, 32'hc4107ae9},
  {32'h43e749b4, 32'h449d0759, 32'h42169a8d},
  {32'h44901ad7, 32'hc39c51b1, 32'h4466e3b0},
  {32'hc3f0efa8, 32'h42abf972, 32'hc40ff343},
  {32'h43515ad0, 32'hc4e0d3f8, 32'h3f108c59},
  {32'hc48cb844, 32'hc2b5d53a, 32'hc50b9bce},
  {32'h43b3ced1, 32'hc35a91cd, 32'h448be683},
  {32'h44cc3588, 32'h429edac6, 32'h437fc158},
  {32'h43175300, 32'hc51caff7, 32'h42c672d0},
  {32'hc4cc5f0e, 32'h43c18176, 32'hc4533192},
  {32'hc31f2e19, 32'hc3d8073c, 32'h449ec5fe},
  {32'hc4925070, 32'h44539d70, 32'hc3e8b9ea},
  {32'h445484de, 32'hc46105d0, 32'hc3c537c1},
  {32'h441c0b8e, 32'h412acbb6, 32'hc43e1d89},
  {32'h44b71b4a, 32'h4397172d, 32'h44ab2bb4},
  {32'hc5103b8e, 32'h43f02162, 32'hc4809c8d},
  {32'h441de073, 32'hc3ac08ad, 32'h44119854},
  {32'hc489ad3d, 32'hc38d49fb, 32'hc3e6966a},
  {32'hc49d0212, 32'h44424f32, 32'h44a06e98},
  {32'h44436bf3, 32'h4451e6f4, 32'hc3fc24b2},
  {32'h4445f174, 32'h4075b458, 32'hc41159d4},
  {32'h44e4d395, 32'hc414b8a3, 32'h41886274},
  {32'hc4eabf74, 32'h433791fa, 32'hc37c0e13},
  {32'h43db50c7, 32'h4119e5cc, 32'h4360147f},
  {32'hc4fc0bca, 32'h444ffb90, 32'h42279aea},
  {32'h434795fd, 32'hc4c4c47a, 32'h44d84bcf},
  {32'h45371e72, 32'h430621e6, 32'h443866b3},
  {32'h4410a800, 32'hc4a740c3, 32'hc4e5cd34},
  {32'h44103a58, 32'h448e697b, 32'hc3ab2146},
  {32'hc4854fdd, 32'hc2a77c66, 32'h44275180},
  {32'hc31e214c, 32'h4310a971, 32'hc5021cc1},
  {32'h43652318, 32'h41c02e20, 32'h44c79d4e},
  {32'h44aab798, 32'h4423bf6f, 32'h4292d6a6},
  {32'h45364ac5, 32'hc1e07c92, 32'hc1b08055},
  {32'hc45107ba, 32'h42ebd23e, 32'hc483480a},
  {32'h4521a2d0, 32'hc3ee9f6e, 32'h440e9e36},
  {32'hc5734aa5, 32'hc42dd58b, 32'hc397956c},
  {32'h4433131a, 32'h4407e523, 32'h437fa31d},
  {32'hc4badab4, 32'hc41347de, 32'hc31999a5},
  {32'h43b52882, 32'hc4dc7299, 32'h4374b166},
  {32'h4267fad4, 32'h454e8157, 32'hc2a4c84d},
  {32'h44c50f4f, 32'h44254c0c, 32'h43a04e03},
  {32'hc485857a, 32'h44bb9a5b, 32'hc41472f8},
  {32'hc3669500, 32'hc5625b95, 32'hc39d6309},
  {32'hc1f59b10, 32'h449ddd39, 32'h4416614a},
  {32'h451db7a6, 32'h425baea6, 32'hc0e7a0f7},
  {32'hc404d332, 32'hc4fc2e54, 32'h44dc274a},
  {32'hc526dbd4, 32'h4389b6c6, 32'h44421da8},
  {32'h44dec269, 32'hc382c58c, 32'h42c70816},
  {32'h44b2a343, 32'hc32ce956, 32'h427032b2},
  {32'h439819b6, 32'h450858db, 32'h42afcf32},
  {32'hc32bdfee, 32'h43a20da0, 32'h45319ed8},
  {32'h440f25d9, 32'hc38888ab, 32'hc3cfcc08},
  {32'h40dd6d50, 32'hc48da9b3, 32'h430f6081},
  {32'hc2dddf6a, 32'hc4f4878b, 32'h44e41e8c},
  {32'h446b53ec, 32'hc4965218, 32'hc49b3ae1},
  {32'h424727f3, 32'h43172d00, 32'hc52f9db3},
  {32'hc0d62e84, 32'hc4dc9977, 32'h43602b92},
  {32'h448bc3ee, 32'h4450ecf3, 32'hc27fec34},
  {32'hc4237e4d, 32'hc4dd8a1c, 32'h43f36e63},
  {32'h42eda01c, 32'h450f3104, 32'hc2e49f3e},
  {32'h44cc5559, 32'hc3fb6ee2, 32'h440e8c35},
  {32'h453ced56, 32'hc34ada97, 32'hc283aa5a},
  {32'hc42371d6, 32'hc3251b30, 32'h43caa534},
  {32'h4587fe70, 32'h433a8961, 32'hc19247ec},
  {32'hc459d60f, 32'hc5001784, 32'hc38c6848},
  {32'h44a7ac22, 32'h448cf167, 32'hc381624f},
  {32'hc3843e5b, 32'hc48ecba5, 32'h441487b2},
  {32'h44b7b23d, 32'h446bd63d, 32'h43d9c140},
  {32'hc532a7c0, 32'hc43943f3, 32'h43f07282},
  {32'h4508e2ed, 32'hc2c804f3, 32'hc34c81db},
  {32'h42f635e3, 32'h44e48bd9, 32'hc371cb0e},
  {32'hc50ee949, 32'hc2b506fc, 32'h42a1b112},
  {32'hc1affb68, 32'h438f36d1, 32'h44a9df96},
  {32'hc3584464, 32'h42c56731, 32'hc45d9011},
  {32'hc12e7d20, 32'h45456f14, 32'h43a545ec},
  {32'hc4c07455, 32'h43a78442, 32'hc496a606},
  {32'h439e0c81, 32'h42a3a0f1, 32'hc1d39649},
  {32'hc4fde92f, 32'hc480b126, 32'hc4a17450},
  {32'h428d57c0, 32'hc2feead0, 32'h44b83c20},
  {32'h43f2538c, 32'hc3d0ac60, 32'hc34f74f7},
  {32'hc455e391, 32'hc3a13a17, 32'h451530fb},
  {32'hc3dc99c5, 32'h44d51de3, 32'hc50597c4},
  {32'h44b5aca4, 32'h438a26e7, 32'h440ddbdb},
  {32'hc3cadb94, 32'hc427c607, 32'hc3e58c45},
  {32'h44abea9c, 32'h439cb5cd, 32'h4453386b},
  {32'hc50bca6a, 32'hc2b74892, 32'h43530b3d},
  {32'h44c8be2c, 32'h43ca7f14, 32'h421d8fe1},
  {32'h4434ff0c, 32'hc3e437e9, 32'hc53dc8cd},
  {32'h4510a40c, 32'h43c005c2, 32'h4229da8c},
  {32'hc43fb2b8, 32'hc4dc8d11, 32'hc44dc231},
  {32'h44da7d48, 32'h4494a67d, 32'h4390f89b},
  {32'h43af860d, 32'hc4edd216, 32'hc351ddb9},
  {32'h452731a6, 32'h42d6f046, 32'h43802aa7},
  {32'hc417591d, 32'hc54f05ad, 32'h43908845},
  {32'hc4c60a94, 32'h435725d8, 32'h440d686b},
  {32'hc53b5201, 32'h43c024ac, 32'hc3a3056b},
  {32'h44ac3fec, 32'hc125151f, 32'h43ff44bd},
  {32'hc38163d7, 32'h4372a66d, 32'hc5052bf7},
  {32'h435784ef, 32'h45225c0f, 32'h4367cdf9},
  {32'hc3b63ec3, 32'hc2f7bc62, 32'hc3b8f87d},
  {32'hc3491578, 32'h409f567e, 32'h44faf2c8},
  {32'h444b2ab8, 32'hc4385435, 32'hc3682e2d},
  {32'h436ee9f0, 32'h44214523, 32'h4201819c},
  {32'h4546216c, 32'hc384557a, 32'hc3ec0faa},
  {32'hc5273fb2, 32'h432296e2, 32'h4414133a},
  {32'hc4492d6e, 32'hc4121ec3, 32'hc3c5c809},
  {32'hc49092e9, 32'hc313a849, 32'h446348a0},
  {32'h427b3fe6, 32'h4309420a, 32'hc42fb352},
  {32'h4340306a, 32'hc4910d30, 32'h44c68e4d},
  {32'h44218ca7, 32'hc3c78940, 32'hc213f5db},
  {32'hc51643e6, 32'h43988b24, 32'h431f5443},
  {32'hc47405e6, 32'hc140c484, 32'hc2aec186},
  {32'hc49a9580, 32'h43e332ea, 32'h44453da6},
  {32'h44d0c7e5, 32'h3d09a2e0, 32'hc3d3d474},
  {32'h438380fd, 32'h44140dae, 32'h4493472c},
  {32'h454f2137, 32'hc44b1cf8, 32'h431eed48},
  {32'hc48fe25c, 32'h4464f6cc, 32'h440ce046},
  {32'h439ca7f5, 32'hc2b92536, 32'h43958dfa},
  {32'hc4ad5157, 32'h44eb7dcc, 32'h4396242a},
  {32'h4509a698, 32'hc2147d60, 32'hc3ab3f9f},
  {32'hc3902fdc, 32'h44931d76, 32'h41ea9525},
  {32'h45586edd, 32'h43c30395, 32'h42993f79},
  {32'hc58a20f0, 32'hc27f66e6, 32'h42dd46d5},
  {32'h4210b69b, 32'hc406dc9c, 32'hc36c6a67},
  {32'h443feda5, 32'h42130e40, 32'h44406b8a},
  {32'hc49a840c, 32'hc19fbbaf, 32'hc3557dc8},
  {32'h44d7fcc5, 32'hc2221fbf, 32'h43d5a90c},
  {32'h44917530, 32'h43ab4d23, 32'hc3066954},
  {32'h44db4264, 32'hc4941843, 32'h4261bce1},
  {32'hc49e8a09, 32'h443a2554, 32'hc1066a41},
  {32'hc3917dda, 32'hc4740222, 32'h422739b2},
  {32'hc569d744, 32'h439d5cce, 32'h431bb111},
  {32'h44f7e514, 32'hc4bdbf7f, 32'h4313bf80},
  {32'h44c86d20, 32'h437b8ef2, 32'hc3dbc6a0},
  {32'h45078f5b, 32'hc323fd94, 32'hc37efdb9},
  {32'hc51a16a2, 32'hc40555ef, 32'h42f5ceca},
  {32'hc36d3d74, 32'hc496e09e, 32'hc2f335fe},
  {32'h433cef04, 32'h44ba52ee, 32'h4471d0cf},
  {32'h43f0eb4f, 32'hc4642f01, 32'hc497cd79},
  {32'hc305b51e, 32'h442197f6, 32'h43b15582},
  {32'h43fdf6db, 32'hc3d14eb0, 32'h4225fca1},
  {32'hc3d3e938, 32'h445a979a, 32'h449d2841},
  {32'h42e429c0, 32'hc2cb90d3, 32'hc40bea03},
  {32'hc50dbade, 32'hc405aff9, 32'h44a0b1c6},
  {32'h44a555ea, 32'h448c55bb, 32'hc445849b},
  {32'hc4b3e42a, 32'h438c3e60, 32'h4311c887},
  {32'hc25dddcb, 32'h423d04bc, 32'hc4f1d3b3},
  {32'hc3e7eb07, 32'h450e1bac, 32'h44129bc7},
  {32'hc328d775, 32'hc2fb9d07, 32'hc490bce4},
  {32'h433b6160, 32'h4481b7cd, 32'h44ed5245},
  {32'h438428e3, 32'hc4c59108, 32'hc441fb9b},
  {32'h4442cf4c, 32'h4466cb4d, 32'hc531ff41},
  {32'hc4608fea, 32'hc3abe075, 32'h45181b85},
  {32'h453f4d3a, 32'h42f03823, 32'hc16ad7ec},
  {32'hc51774b0, 32'h436ebbfc, 32'hc252f4dc},
  {32'h4459b2c0, 32'h44607450, 32'hc3881415},
  {32'hc459d2b2, 32'hc4a0e68f, 32'hc30f285c},
  {32'h451a98c3, 32'h4479bf4e, 32'h41499f98},
  {32'hc49da862, 32'hc4add43d, 32'h42415eda},
  {32'hc333ef95, 32'h42dca8d6, 32'h43dc203a},
  {32'hc4fb91cf, 32'hc13268f8, 32'h4362fb9c},
  {32'h44de26be, 32'hc2a60e35, 32'hc44591d2},
  {32'hc50d8bd8, 32'hc3ae3ee7, 32'h42c3f6e9},
  {32'h4389c400, 32'h44ac2219, 32'h4469a5c7},
  {32'hc50199ff, 32'hc438cebf, 32'h43147278},
  {32'hc366c5e9, 32'h43ef2862, 32'h432cc392},
  {32'hc4ecee76, 32'hc3b7e6c4, 32'hc3e7ad95},
  {32'hc394a142, 32'h43df0e5f, 32'h44cefc07},
  {32'hc23430e0, 32'hc3e8535b, 32'hc490f635},
  {32'h450fc93a, 32'h443ca6a0, 32'h446485cc},
  {32'hc498e612, 32'h4433eef4, 32'hc34a02fd},
  {32'hc2f0c418, 32'hc391a91a, 32'hc3be24b6},
  {32'hc5019ebc, 32'hc3e3b880, 32'h420e4eb0},
  {32'h44c9e10a, 32'h4403cbc4, 32'hc2824889},
  {32'h44856e14, 32'hc2b14684, 32'h42d08748},
  {32'h436c687d, 32'h448642ea, 32'h450f4391},
  {32'hc4d2fca0, 32'hc44ae769, 32'hc3cacbb2},
  {32'hc2a951d5, 32'hc3732f76, 32'h4501b864},
  {32'h438ffd17, 32'h43c557b6, 32'h440c2dbd},
  {32'hc501ef91, 32'hc3c33ea2, 32'h427e14c9},
  {32'h453b872b, 32'h43a5e814, 32'h43b257dc},
  {32'h42ebe100, 32'hc2d589bf, 32'h424a7bf8},
  {32'h45421b36, 32'h43cd58cc, 32'h405ba938},
  {32'hc42f0487, 32'hc5267ca3, 32'h43a258b7},
  {32'hc42f37b1, 32'h440c5bc8, 32'hc38d5474},
  {32'hc56d0e1f, 32'h43addd39, 32'hc3355e92},
  {32'h4544456a, 32'hc2da9a44, 32'h43fee25b},
  {32'hc390dd6b, 32'hc431a1df, 32'h438fda06},
  {32'h4372caa0, 32'h44837c17, 32'hc48be5c9},
  {32'hc41fc7b3, 32'hc413bd1a, 32'h445d421a},
  {32'h43dd6720, 32'h43ed6894, 32'h42e943cf},
  {32'hc50a286b, 32'h439a05d0, 32'h41133c5a},
  {32'h44a6bd63, 32'h4438efc3, 32'h43199297},
  {32'hc50ce1a8, 32'h430d1978, 32'h4308c0bf},
  {32'h424e67a0, 32'hc39dff0a, 32'hc4e523c0},
  {32'hc493dea6, 32'hc3975d40, 32'h432d7844},
  {32'hc48c060a, 32'h438b76be, 32'hc3324096},
  {32'hc4331218, 32'hc4912725, 32'h44e23122},
  {32'h43758e68, 32'h447a4c1a, 32'hc4eb4f4a},
  {32'h43928c60, 32'hc4861371, 32'h4388a9e4},
  {32'h43e24670, 32'h446bd30e, 32'hc4814741},
  {32'hc40b0284, 32'hc4adc086, 32'h430d79d7},
  {32'h44a71d4a, 32'h434f304f, 32'hc0ed4d00},
  {32'hc49a2bf9, 32'h42bb1d3a, 32'h447d3c8d},
  {32'h42c9dfad, 32'hc2169341, 32'hc44366c2},
  {32'h44469a32, 32'hc4cdebf1, 32'hc3968638},
  {32'hc5252c32, 32'h43b00b77, 32'hc38e72a0},
  {32'h44eba5e9, 32'h436da3e0, 32'h441056f0},
  {32'hc4342351, 32'h43431f50, 32'hc410092b},
  {32'h43348098, 32'hc4699520, 32'hc3f4385c},
  {32'hc2fc0ced, 32'h44e706db, 32'hc3b4dd0f},
  {32'hc301610f, 32'hc39a5921, 32'hc381ffa8},
  {32'hc4d3096c, 32'hc21f2393, 32'h43a8a60d},
  {32'h450e51c0, 32'hc4329bc6, 32'h432751de},
  {32'hc470af74, 32'h44549842, 32'hc42cd91f},
  {32'h4412688a, 32'hc47e2722, 32'hc38d8be8},
  {32'h448e4b46, 32'h42806e2d, 32'h441e0f0e},
  {32'h4359ee30, 32'hc4ccc723, 32'h4356ecc2},
  {32'hc2c39285, 32'h455311e5, 32'hc3ac1870},
  {32'hc45a585f, 32'h4355deaa, 32'h44e2d2f4},
  {32'hc5115c28, 32'h43aa5d1e, 32'h43fb792a},
  {32'h4454b336, 32'hc1d7203e, 32'h44b34952},
  {32'hc3f021c0, 32'hc3c4da82, 32'hc443182b},
  {32'hc3a635c0, 32'hc4a86174, 32'h442c50be},
  {32'hc5418102, 32'h438027fb, 32'hc3362a75},
  {32'h4363338d, 32'hc4c479e7, 32'hc28677da},
  {32'hc3a845a4, 32'hc36fed90, 32'hc4b3b039},
  {32'h430794d1, 32'hc2d45e8f, 32'h453f65e3},
  {32'h4488edd4, 32'h44032bd7, 32'hc37aefdc},
  {32'h44d5015e, 32'h426727a3, 32'h44656fbe},
  {32'hc4773bd8, 32'hc40c3666, 32'hc5122d4d},
  {32'h45052de2, 32'hc225eeaf, 32'h425d208c},
  {32'hc2faf520, 32'hc42e17dc, 32'hc4cd736c},
  {32'hc409b974, 32'hc47a855e, 32'h44c7ea67},
  {32'h44e3b8ef, 32'h43ba24f6, 32'hc3c51a21},
  {32'h42defc3c, 32'hc0f29920, 32'hc43b442f},
  {32'h4449e5f5, 32'h42eaafb7, 32'h43d84b71},
  {32'hc4bb50ed, 32'h44743be6, 32'hc2c12d3f},
  {32'h419451f0, 32'hc3b8bb3d, 32'h449bb763},
  {32'hc2fd384c, 32'h43d040b2, 32'hc4c05c5a},
  {32'h43513ce8, 32'hc3374805, 32'h454e6d08},
  {32'h44b5a265, 32'hc492df15, 32'h4476f253},
  {32'hc315d620, 32'hc34f7a2b, 32'hc4ab28fa},
  {32'h4488e3ac, 32'hc39fdc43, 32'h42a346e5},
  {32'h4307ef57, 32'hc4bb28b2, 32'h4312902f},
  {32'hc3ce6cec, 32'h44bb9844, 32'h44052743},
  {32'h43b11ee8, 32'hc20ef88d, 32'h4519cb6a},
  {32'hc4365a59, 32'hc22477ae, 32'hc38029c6},
  {32'h43d431f0, 32'hc33f39d0, 32'h44b0772d},
  {32'hc3e6f18e, 32'hc368d2f6, 32'hc4be5175},
  {32'hc48294cc, 32'h43152c8a, 32'h440d35d1},
  {32'hc3fd1a20, 32'hc3f6965a, 32'h4325142a},
  {32'h4419348e, 32'hc3bbc4c1, 32'hc2b6fd4a},
  {32'hc52816a9, 32'hc3c6669b, 32'h42b5e7c6},
  {32'hc4267b2e, 32'hc505dba9, 32'h40c6e610},
  {32'hc53eda80, 32'h42564214, 32'h43bda7b4},
  {32'hc300e1a5, 32'hc49d107f, 32'h43b47ca4},
  {32'hc32fdbb4, 32'h456f3a50, 32'hc3b31fa4},
  {32'hc2c2ba40, 32'hc5667082, 32'h42b37d9a},
  {32'h442fbf08, 32'h43b1c9bd, 32'h4508526c},
  {32'h439f9fd1, 32'h409d32e6, 32'hc49a583f},
  {32'hc32706e4, 32'h43fa671c, 32'h44d4468f},
  {32'hc353ae0a, 32'hc33eae96, 32'h4540f908},
  {32'h44512d70, 32'h43c620e3, 32'hc42c07c3},
  {32'h444df61f, 32'hc32b3160, 32'h439a4592},
  {32'h452cabe1, 32'h43f15e90, 32'hc404d894},
  {32'hc3bbd674, 32'hc5249172, 32'h4283d58d},
  {32'h443c15db, 32'hc3915474, 32'hc49f5ddf},
  {32'hc41ddcbf, 32'hc4499b36, 32'h4330e753},
  {32'hc42f185a, 32'h4433b692, 32'h44d861dd},
  {32'h43b17902, 32'hc499681c, 32'hc4c32fa3},
  {32'h44a9d141, 32'h44317229, 32'hc3bb4cff},
  {32'hc490acce, 32'hc42ffb50, 32'h445fe47c},
  {32'h452147e6, 32'h438bb236, 32'hc3385aa9},
  {32'hc4f82510, 32'hc39913e7, 32'h448374af},
  {32'h43b94c20, 32'h448a1ffd, 32'hc402486e},
  {32'h43eac3d4, 32'hc1adba9a, 32'h44887ee5},
  {32'h42a24280, 32'hc42554c2, 32'hc43f7443},
  {32'hc5827c10, 32'h42f36ba3, 32'h439c43e2},
  {32'h44fc4890, 32'h44525c4f, 32'h408672c8},
  {32'hc4b561b6, 32'h438d9365, 32'hc38d5b89},
  {32'h4336f931, 32'h450af4b7, 32'hc39012b3},
  {32'h43459c1a, 32'hc4c71bf4, 32'hc11a248d},
  {32'h42f771d0, 32'h44cbef75, 32'h4220cc06},
  {32'hc4ff4244, 32'hc4703895, 32'h4275157a},
  {32'h455ad780, 32'hc44eb5a4, 32'hc36e7088},
  {32'hc4012d80, 32'h4348913a, 32'hc281a847},
  {32'h445cceb5, 32'h441a00fd, 32'hc3b05b13},
  {32'h44124204, 32'hc2387b19, 32'h44831c6c},
  {32'h441edeb4, 32'hc0dba72c, 32'hc3f02884},
  {32'h43df4d03, 32'h452c7ea3, 32'h422555bc},
  {32'hc50f9674, 32'h43ff00bc, 32'h43c73ed1},
  {32'h433f855b, 32'h42ffef7a, 32'h44a69950},
  {32'hc2a0699e, 32'h4392d175, 32'hc3662511},
  {32'hc3abfe80, 32'h44160bce, 32'h45385598},
  {32'h4402a47c, 32'h4336d1d1, 32'hc3c007d5},
  {32'hc4376761, 32'h43bf6a9a, 32'h437ca62f},
  {32'hc28ac8c6, 32'hc4f0b478, 32'hc4384151},
  {32'hc5006cc9, 32'h42cbe808, 32'hc1fb55d5},
  {32'hc52cb93a, 32'hc39dc88d, 32'h431f3634},
  {32'hc3cf1428, 32'h443a7eed, 32'h44b119a2},
  {32'h4415dd8b, 32'hc30fe5d1, 32'hc505fe19},
  {32'h42e9f150, 32'h44a0a0da, 32'h44d7eb06},
  {32'hc49e2218, 32'hc3813a6d, 32'hc414738a},
  {32'h4522c610, 32'hc3c0b9d0, 32'h43eec992},
  {32'hc4a49500, 32'hc494f9cf, 32'hc3fa7176},
  {32'h454db32a, 32'h4411a998, 32'h4396fae4},
  {32'h445fe51a, 32'hc46c0396, 32'hc2df881a},
  {32'hc36f9969, 32'h4586d9d8, 32'hc36c43f7},
  {32'hc4871f15, 32'hc50a00bb, 32'hc3122ef0},
  {32'hc4b6c21e, 32'h43fe43a6, 32'h43cfe095},
  {32'hc40e93da, 32'hc3c057ef, 32'hc40a0a35},
  {32'h43e64f60, 32'hc4222b2d, 32'hc39b2c53},
  {32'h43595b64, 32'h44b14954, 32'hc4eb5881},
  {32'hc0b781cc, 32'h43ecc70f, 32'h4383f51c},
  {32'h431af042, 32'h422d1a99, 32'hc4cdc797},
  {32'hc464bf74, 32'h44865528, 32'h44982446},
  {32'hc1a36020, 32'hc47db711, 32'hc42a56b8},
  {32'hc35223ee, 32'h44eb5d66, 32'h43d58d56},
  {32'h4539ce68, 32'hc31fb190, 32'hc3f53fe8},
  {32'hc45167b5, 32'h44be423e, 32'h446adef4},
  {32'hc4bdc4b4, 32'hc40f110b, 32'hc2dbedba},
  {32'h441a114f, 32'h44ccab9f, 32'h44206202},
  {32'hc4cb65da, 32'h44340387, 32'hc426cb12},
  {32'hc4d4007b, 32'h43473146, 32'hc37d9b9e},
  {32'h443ca3cc, 32'hc2ef72f0, 32'hc48618cc},
  {32'hc349102c, 32'h43aa5b3c, 32'h4500f34d},
  {32'hc44bdfad, 32'hc28843e2, 32'hc2f9fb19},
  {32'hc41d5eed, 32'h4426c6d2, 32'h44226cdd},
  {32'h44002f7a, 32'hc2c8ba13, 32'hc4f4f913},
  {32'h43c9cd24, 32'h44a6548e, 32'h445df4b6},
  {32'h450d75d0, 32'hc456ae96, 32'h4309d42f},
  {32'hc475cb6a, 32'h450648d0, 32'hc373b2f0},
  {32'h451bccb4, 32'h442101a4, 32'h4311853a},
  {32'hc45d5c98, 32'h4504610f, 32'hc31b299f},
  {32'h43a1e898, 32'hc4d6fa5c, 32'hc3f453a0},
  {32'h43b41435, 32'h4190cde2, 32'hc30b0b9b},
  {32'h452866bf, 32'h43f8c4fb, 32'hc2816f37},
  {32'hc5866c65, 32'h44070104, 32'hc38f720d},
  {32'hc43b7c2c, 32'h43ca6678, 32'h428a4250},
  {32'h44b40363, 32'hc3d400fd, 32'h43129688},
  {32'hc555063f, 32'h429e59be, 32'hc31f5d5e},
  {32'h44e87244, 32'hc297df92, 32'h445906c4},
  {32'hc543c5c1, 32'hc2ca7330, 32'hc30d10ba},
  {32'h43bd1b01, 32'hc5344307, 32'hc32afa4e},
  {32'hc4347fda, 32'h449a066e, 32'h42a00eea},
  {32'hc4e7345b, 32'hc2a6d90e, 32'h4390ca13},
  {32'hc45f0f50, 32'h449fdc85, 32'h438d485c},
  {32'h4520fd1d, 32'hc3befced, 32'h4282ae99},
  {32'hc41d092d, 32'h440be63b, 32'h3f8edf20},
  {32'h44193b30, 32'hc35b6c2d, 32'h44d9b3c3},
  {32'hc2fa8a30, 32'h433fa0c5, 32'hc434e55f},
  {32'hc22ebb7e, 32'hc2b0f505, 32'hc4a1db2a},
  {32'hc5041a93, 32'h42f7318a, 32'h42b35a21},
  {32'h44815592, 32'hc44c196f, 32'hc3834aa4},
  {32'h44a65a40, 32'hc32b7424, 32'h43bea824},
  {32'hc3f8f098, 32'h424a71b2, 32'hc529e0d6},
  {32'hc2ce7ee0, 32'h440dbf37, 32'h42ce6ba2},
  {32'h431a4f10, 32'h43a4da70, 32'hc393351c},
  {32'hc53bc75c, 32'hc415a223, 32'h431a159e},
  {32'h451a6317, 32'hc29d612f, 32'hc43a5100},
  {32'hc4372746, 32'hc360b8a2, 32'hc2a26277},
  {32'h4511e8c8, 32'hc3e07318, 32'hc2dbe05e},
  {32'hc38d55d4, 32'h44d86f38, 32'h440eec7b},
  {32'hc34a7360, 32'hc3046976, 32'hc509bf53},
  {32'hc4e5d8ad, 32'h4442d1ac, 32'hc39167c2},
  {32'hc1bbee38, 32'hc462075b, 32'hc3d4af7f},
  {32'hc38fb864, 32'h43257a74, 32'hc4ac75b8},
  {32'hc53c135c, 32'h4395db25, 32'h43e99214},
  {32'hc39201e4, 32'h4349244e, 32'hc3b32fbb},
  {32'h4214ad94, 32'hc50ff51c, 32'hc3587e78},
  {32'h44a0eeb6, 32'h42a6f6b8, 32'h42c34a2d},
  {32'h43905239, 32'hc529bde1, 32'h42a8b54e},
  {32'h4538c55d, 32'h445fd0f5, 32'hc33c0a5b},
  {32'hc3e6144e, 32'hc497caba, 32'h4423b1e8},
  {32'h451ecd37, 32'h42f64b04, 32'h439cdd29},
  {32'hc4f12914, 32'hc4454657, 32'h43928b0a},
  {32'h440fe60c, 32'h43b6b642, 32'hc492eb96},
  {32'h4429d9c1, 32'h3fea06e2, 32'h436453c8},
  {32'h44215644, 32'h43886911, 32'h4310a882},
  {32'hc400eee3, 32'hc414b235, 32'hc537b92b},
  {32'hc416611a, 32'h43222f52, 32'h443421fa},
  {32'hc526ac8b, 32'hc301035b, 32'h425c427f},
  {32'h42de58e2, 32'h44e6d014, 32'h43959003},
  {32'hc38fd8c9, 32'hc13f2ff6, 32'hc4038dac},
  {32'h45084de7, 32'hc32b31ad, 32'h441d4bde},
  {32'hc50b6adb, 32'hc2b0ac81, 32'hc39af005},
  {32'hc36ecc50, 32'hc41e344e, 32'h43409e8e},
  {32'h43cd6faa, 32'hc42328a6, 32'hc51b7729},
  {32'h44c1459a, 32'h445dec66, 32'h4417eb8e},
  {32'hc4194083, 32'hc43e00a3, 32'h428801d2},
  {32'h44866538, 32'h42e6aab4, 32'h43a3d54e},
  {32'hc3c4bfbe, 32'hc3027de2, 32'hc4b2e2c6},
  {32'hc39a0939, 32'h44989793, 32'hc365c350},
  {32'hc3a2824c, 32'h4354e19e, 32'hc4114a44},
  {32'hc3cdfecd, 32'hc529a8cc, 32'h42bdf294},
  {32'h4421790b, 32'h44fa678a, 32'hc377cb54},
  {32'hc400869e, 32'hc3d2056c, 32'h42f3e4c5},
  {32'h4389f714, 32'h4531d08f, 32'h4269aca5},
  {32'hc50b1b11, 32'hc4451901, 32'hc39f3b6b},
  {32'h456f6582, 32'h43b289b2, 32'hc36f193d},
  {32'hc52d32e0, 32'hc3efb594, 32'hc36dc5eb},
  {32'h455fe59d, 32'h41097aef, 32'hc3523221},
  {32'hbf048dc0, 32'hc40487a2, 32'h44afe536},
  {32'h4441c362, 32'h43a178c9, 32'h436ad58c},
  {32'hc436a04c, 32'hc3dc0cb1, 32'hc3ca23c1},
  {32'hc3de3eed, 32'hc2b88305, 32'hc4b722e9},
  {32'h42100530, 32'hc4397005, 32'h445f7c54},
  {32'h4489f708, 32'h42934164, 32'hc4b815a2},
  {32'h44bd75e2, 32'hc2907b10, 32'hc2df59fc},
  {32'h43d7120c, 32'h43c24345, 32'hc3d87efb},
  {32'hc3b3a724, 32'h41a03bf2, 32'h44bd6f97},
  {32'hc3397c30, 32'h44a5a67d, 32'hc2f46fce},
  {32'hc5151eb8, 32'hc414e3e0, 32'hc3782e0c},
  {32'h4522267f, 32'h441b1a3c, 32'hc47e9079},
  {32'h43e87c42, 32'h433f8af9, 32'h4492f142},
  {32'h433f9140, 32'h444ac208, 32'hc467fdbb},
  {32'hc41919f0, 32'hc49b9cbb, 32'h4492c706},
  {32'hc499e389, 32'hc31e7a24, 32'hc341c31d},
  {32'hc40fa286, 32'h4444921c, 32'h454e94be},
  {32'h4513e4ce, 32'hc31ff340, 32'hc473b825},
  {32'h446025ea, 32'hc45f1fed, 32'hc446eb76},
  {32'hc4a3dd32, 32'h4450d22a, 32'h410b7fc9},
  {32'h43ca1cfa, 32'h432b3daa, 32'h4395c762},
  {32'hc4bd851f, 32'h448b3ffe, 32'h437a3111},
  {32'h437d41fa, 32'hc4c5bced, 32'hc3c10640},
  {32'hc406cfa7, 32'h43d4ba23, 32'h43498ccb},
  {32'h4540e714, 32'h437c7877, 32'hc34b98a3},
  {32'hc4060eb4, 32'h44928a13, 32'h4477dd55},
  {32'h445fd13a, 32'hc2b56a54, 32'h443b280a},
  {32'hc33a052c, 32'h4482a91e, 32'hc49b82bc},
  {32'h44881066, 32'hc4153596, 32'h44981a51},
  {32'h44235cda, 32'h43ae8294, 32'hc39e3c52},
  {32'h43911418, 32'h43028bc4, 32'h43fd54df},
  {32'hc440d0b4, 32'h43c4c585, 32'hc4888ff2},
  {32'hc452c0a7, 32'h43955cf8, 32'h43a38a48},
  {32'hc4605a31, 32'h42e368c9, 32'hc49e80d6},
  {32'h454cadba, 32'h4402817d, 32'hc2fdc324},
  {32'hc3d7dde4, 32'hc381c13a, 32'hc48ffd3b},
  {32'h441b2988, 32'hc4ba15bd, 32'h44236270},
  {32'hc4c23b13, 32'h43d843a5, 32'hc403c26d},
  {32'h43b48bc0, 32'hc4497bb1, 32'hc3e60975},
  {32'hc429f96f, 32'h43da5c43, 32'hc4b33bdb},
  {32'h4342f470, 32'hc46b7a07, 32'h445cee91},
  {32'h42598606, 32'h439337b4, 32'hc5037788},
  {32'h45242e0f, 32'hc29246cb, 32'h4469902a},
  {32'hc4419524, 32'h42f1995f, 32'hc4e68102},
  {32'hc47b554c, 32'hc30cf0f4, 32'h429baa0e},
  {32'hc2d6c544, 32'hc437eec9, 32'hc54a9dae},
  {32'hc3d60a1a, 32'h442d2817, 32'h440b2656},
  {32'h44564982, 32'hc415cdf2, 32'hc40e3940},
  {32'hc4551a97, 32'hc28d86b1, 32'hc3ab1d26},
  {32'h44455eb3, 32'hc49354b3, 32'h434a5e7a},
  {32'hc3e0dfec, 32'hc3d8d251, 32'hc516c6a6},
  {32'h442aedd2, 32'hc361d204, 32'h42ae5d95},
  {32'hc32de040, 32'h4519ac95, 32'hc3a8fd33},
  {32'hc32fd8e8, 32'h43671189, 32'h4584c316},
  {32'h448f0130, 32'h4246cba0, 32'h449e22b7},
  {32'hc3543fcb, 32'hc44771fb, 32'hc4c8d65c},
  {32'hc3889d37, 32'hc410edcc, 32'h43c90944},
  {32'h4494095b, 32'hc3eb5796, 32'h434a2bbf},
  {32'hc4b2f326, 32'h43c6260a, 32'hc38e0f31},
  {32'h4476580f, 32'hc4763136, 32'hc3768221},
  {32'h44d32700, 32'hc3825784, 32'h43b20b83},
  {32'h451c41ee, 32'h433d7282, 32'hc3faafc5},
  {32'hc4a9eec0, 32'h439686b8, 32'hc41c7c62},
  {32'hc5059632, 32'h419f7762, 32'hc28116b0},
  {32'hc5930b61, 32'h42852c3e, 32'h40b330e6},
  {32'h4584b99b, 32'hc31dd0c6, 32'hc38f986e},
  {32'h43c0c09a, 32'h43223081, 32'h41a070ee},
  {32'hc317a0f6, 32'hc57e0d68, 32'hc3b5eb33},
  {32'hc4f287bd, 32'h44197ff8, 32'hc310596e},
  {32'h445a9cc1, 32'hc4e14876, 32'h4324d062},
  {32'hc444127a, 32'h45708b72, 32'hc31031f9},
  {32'hc3a95578, 32'hc4d61b42, 32'hc30d6af0},
  {32'h43c14250, 32'hc4d77ede, 32'h43f89eef},
  {32'h43a9ff7a, 32'h42dee1ba, 32'h430d189d},
  {32'hc4a0dd8c, 32'h4478414d, 32'h443f348a},
  {32'hc501b16b, 32'hc3e681b6, 32'h442e8be7},
  {32'h45076d6c, 32'h430f449f, 32'h430b6e39},
  {32'hc3856b4a, 32'hc4491ae3, 32'h44878546},
  {32'hc1d83218, 32'h449d2740, 32'hc50e8dcd},
  {32'hc20fe672, 32'hc358baf5, 32'h452b418f},
  {32'hc28915ac, 32'h432f2201, 32'hc4009e24},
  {32'h431a28d1, 32'hc39774b9, 32'hc48acf80},
  {32'h42c1760d, 32'hc48a56d2, 32'h44462141},
  {32'h450a4f50, 32'h43efbf47, 32'hc444d91c},
  {32'h4412e990, 32'h43afadfa, 32'hc4ac8819},
  {32'hc3b16d3a, 32'hc51f3dbc, 32'hc3087ff4},
  {32'h435e98eb, 32'h430b3916, 32'hc4c5a135},
  {32'hc49421b4, 32'hc4aec0ab, 32'h439e55f4},
  {32'hc32c2cc1, 32'h43a6a214, 32'hc5133f58},
  {32'hc5004f64, 32'hc33377c9, 32'hc33abd0c},
  {32'h44dbdcf8, 32'hc4117f52, 32'hc40a325c},
  {32'hc58fe691, 32'hc28ea99c, 32'h43a22994},
  {32'h44fbdaa4, 32'h4347065c, 32'h4339ff48},
  {32'h43b9666c, 32'hc542b151, 32'h3f031460},
  {32'h450c5464, 32'h442d63de, 32'h40c0656c},
  {32'hc507518e, 32'h43a52341, 32'h4239211f},
  {32'h4509115b, 32'h44534cd2, 32'h43bb099e},
  {32'hc4d6acbe, 32'hc499a7ef, 32'hc1eedfff},
  {32'h4530a6c9, 32'hc11d3f0b, 32'hc39225c6},
  {32'hc06aefb8, 32'hc3b467da, 32'h4434007b},
  {32'hc4346f61, 32'hc2952ebb, 32'hc3d100ba},
  {32'h434491d2, 32'h4504ac4f, 32'h43f8e319},
  {32'h4420122d, 32'hc37be825, 32'hc380b49e},
  {32'h44d82361, 32'h43e54be8, 32'h44924fc5},
  {32'hc374af74, 32'hc5281a2c, 32'hc3f2a0fe},
  {32'h452697f8, 32'hc3d5c2ee, 32'hc382e8c3},
  {32'hc556c943, 32'hc39b1b54, 32'hc3d627d2},
  {32'h44850690, 32'hc1aa582e, 32'h44246a39},
  {32'h4347bf40, 32'h436a47a9, 32'hc4ba9dd4},
  {32'hc38feec6, 32'h4347a5ea, 32'h44874b48},
  {32'hc33ba6b8, 32'hc431af49, 32'hc4bae5bc},
  {32'hc3cb482c, 32'h42d3dadc, 32'h43963229},
  {32'hc43074da, 32'hc4e79904, 32'hc419484f},
  {32'hc330285b, 32'hc2d0e79d, 32'h45150c58},
  {32'h44b41174, 32'hc4458d54, 32'hc3af30bc},
  {32'h449e3c05, 32'h43c6c888, 32'h43b677d4},
  {32'hc42ced74, 32'hc43d749d, 32'hc46a9783},
  {32'h44fe8a59, 32'hc120130c, 32'h448e948f},
  {32'hc4355e5a, 32'hc52ddcc3, 32'h4333bd0d},
  {32'h455e9be1, 32'hc2e7936b, 32'h438d960a},
  {32'hc54721df, 32'h435e76b6, 32'h42de25d8},
  {32'hc29978fc, 32'h4538c8ff, 32'hc25e7af7},
  {32'hc484061e, 32'hc4a9c610, 32'h439e07c2},
  {32'h44d8c592, 32'hc27fb4a6, 32'h43cc0c5a},
  {32'hc59482fc, 32'h43682d23, 32'hc30a7e57},
  {32'h45127f10, 32'h42c7d835, 32'hc36b5c5c},
  {32'h436c8370, 32'h44124239, 32'hc4a0b1de},
  {32'hc3acf2cc, 32'h438a0717, 32'h44b25b7c},
  {32'h41f2f7c0, 32'hc380691e, 32'hc4483cce},
  {32'h4133647a, 32'h44c24835, 32'hc1ce2e29},
  {32'h45335392, 32'hc39d2dab, 32'h420f699a},
  {32'h44b03f64, 32'h4325271e, 32'h43b38f30},
  {32'h44266db4, 32'hc3495254, 32'hc48325ef},
  {32'hc516ba69, 32'h440c945e, 32'hc2cd42cc},
  {32'hc36674fc, 32'hc435a51c, 32'hc3764d29},
  {32'h43f5c8e4, 32'hc3cdf1e0, 32'h4510926f},
  {32'hc3a52f08, 32'h44575e3f, 32'hc5197293},
  {32'hc48cd535, 32'hc3637f85, 32'h43cdaa8f},
  {32'h43efa3d8, 32'hc4ede3bb, 32'hc29d7324},
  {32'hc38db43a, 32'h43b4937b, 32'h44d8e72f},
  {32'h438e7c6b, 32'hc105f04f, 32'hc4d2d030},
  {32'hc4b32cbb, 32'h41a0f682, 32'h442dbf85},
  {32'h44641b85, 32'hc48f3f99, 32'hc4cfa2bf},
  {32'h44120cd2, 32'h43921ad1, 32'h43444d70},
  {32'h449a4700, 32'hc4ba7df1, 32'h42f4118a},
  {32'hc2f7ab44, 32'h4518ff4e, 32'h433d050a},
  {32'h43b0a63e, 32'hc389f285, 32'hc3f14060},
  {32'hc49ee31c, 32'h44db08e6, 32'hc288a925},
  {32'h4383fe04, 32'hc4d54d3a, 32'hc39ddb6d},
  {32'h449430e7, 32'hc35990cf, 32'h440cd4db},
  {32'h45171416, 32'h43f981c2, 32'hc3038be3},
  {32'hc575e41c, 32'hc1a7c06d, 32'hc3a95ddc},
  {32'h417e5d03, 32'hc4124fd4, 32'hc38dc609},
  {32'h44fd5993, 32'hc360df5a, 32'hc24224f1},
  {32'hc5113b12, 32'h42806c83, 32'hc4308da0},
  {32'h4443a20e, 32'h43baeca0, 32'h450a8fec},
  {32'hc4525aa1, 32'h445bd39a, 32'h438e08b1},
  {32'h43889070, 32'hc4d8663c, 32'hc28683fe},
  {32'hc404b0f6, 32'h44e07c1b, 32'h434c63d4},
  {32'h44d54a2f, 32'h43083329, 32'hc2d78c15},
  {32'hc3c12218, 32'h44f3be8f, 32'h440ec63b},
  {32'h43f07900, 32'hc460cded, 32'h43bebe19},
  {32'h4386a2c4, 32'h42f614cd, 32'hc386c4e2},
  {32'h4459af68, 32'hc4677cb9, 32'hc3b4c167},
  {32'hc504227e, 32'hc3064fcb, 32'hc4237815},
  {32'hc4646712, 32'hc2fe3c3d, 32'h42d78d7c},
  {32'h43bbddac, 32'h44a0d871, 32'h442d230f},
  {32'h4505d35c, 32'hc3a77c89, 32'hc34c456a},
  {32'h438e788f, 32'hc380f19f, 32'h4497994f},
  {32'h431f6578, 32'hc4074c14, 32'hc4da89ce},
  {32'hc543e3e7, 32'hc40c54b3, 32'hc30dbab4},
  {32'hc4891cdf, 32'hc3c14fcb, 32'hc379d4e2},
  {32'hc4682134, 32'h443d9d90, 32'h44b1489e},
  {32'h44953de0, 32'hc3cb1225, 32'hc4511a93},
  {32'hc30d8440, 32'h44d27fca, 32'hc3c8fe28},
  {32'h424a4048, 32'hc42282f5, 32'hc4daf55b},
  {32'hc4e14d69, 32'h43a95d7e, 32'h447b1d9b},
  {32'h441c0e22, 32'hc410daa5, 32'hc430d573},
  {32'hc4c36ce9, 32'h42ed378a, 32'h446a2b4c},
  {32'h44ec95f3, 32'hc43666f5, 32'hc4439a7b},
  {32'h440d326f, 32'hc18e24e6, 32'hc4d7ab2a},
  {32'hc38eaeba, 32'h43966682, 32'h45201722},
  {32'h44a05707, 32'hc2766b94, 32'h44221c5a},
  {32'hc41e1374, 32'hc5105f38, 32'hc309a4c7},
  {32'h433e4f4a, 32'h453a511f, 32'h433b3526},
  {32'hc2c08078, 32'hc4a112f1, 32'h437f72f4},
  {32'h4301a59d, 32'h4587fb93, 32'hc33302fa},
  {32'hc4b8ab64, 32'hc48d3ee2, 32'hc43639b2},
  {32'hc419d4da, 32'h4391a00b, 32'h43f4a272},
  {32'hc52f4e72, 32'hc3ff7ea0, 32'h426efb1e},
  {32'h4341be36, 32'hc3f3abca, 32'h442bf425},
  {32'h44af1eb2, 32'hc39b701e, 32'h44407ea1},
  {32'h439f3570, 32'hc0f71d00, 32'h44800c41},
  {32'hc4da3f0e, 32'hc41f6c60, 32'hc4b5f384},
  {32'hc48956cf, 32'h43e581ae, 32'h4413f42e},
  {32'h411d3720, 32'hc34bff87, 32'hc5593aa6},
  {32'h443c9f4c, 32'h442783d8, 32'hc392abd8},
  {32'hc50bd18f, 32'hc399955d, 32'hc3967bf4},
  {32'h44d8476f, 32'h44135739, 32'h44195b86},
  {32'hc59df860, 32'h42bef571, 32'h42da8989},
  {32'h4533701d, 32'h42bfbc5c, 32'hc3e05c9c},
  {32'hc38045fc, 32'hc25a7446, 32'hc5208617},
  {32'h43574fe2, 32'h43e99708, 32'h44a04d8e},
  {32'h43950b10, 32'hc32b7400, 32'hc4516aed},
  {32'h433f7a48, 32'h4480a8e6, 32'h4510a3ed},
  {32'hc4cafca0, 32'h4286c2b0, 32'hc4ac79e9},
  {32'hc3815620, 32'h44891fb2, 32'hc4168687},
  {32'h4492061c, 32'hc30d37a7, 32'hc3fab015},
  {32'hc38bc328, 32'hc485d8e8, 32'hc430ae22},
  {32'h446c5416, 32'h44ba1f69, 32'h43c67287},
  {32'hc4e5d331, 32'hc370dac5, 32'h42900b66},
  {32'h44984ab0, 32'h4451eded, 32'hc24da4f9},
  {32'hc4f5e40c, 32'hc4297472, 32'hc303a1af},
  {32'h4538fccd, 32'hc35c7fcc, 32'hc4030bed},
  {32'hc58adccb, 32'h437e5b3c, 32'h43f9e318},
  {32'h456c31c8, 32'hc3e58b0a, 32'h40454740},
  {32'h44c7d79a, 32'hc397b9f8, 32'h43e33bad},
  {32'h430edc40, 32'hc4083b85, 32'h4487739d},
  {32'hc30ee6dc, 32'hc509bc73, 32'hc20b38ee},
  {32'h42238083, 32'hc386f012, 32'hc4bb2014},
  {32'hc50d5587, 32'hc3c7ecf2, 32'h4357ef74},
  {32'h444354be, 32'h43b374b8, 32'hc41bc4f8},
  {32'hc3ae45e0, 32'hc37f843f, 32'h43825217},
  {32'h45296b10, 32'hc46cbb71, 32'hc2bf084b},
  {32'hc505c8bc, 32'hbf16c67c, 32'h441049c6},
  {32'hc30e4fae, 32'h43d19d6a, 32'hc41653de},
  {32'hc49da2d5, 32'hc465e4f0, 32'h44b153dd},
  {32'h4507ed24, 32'h44617593, 32'hc462bb02},
  {32'h42285e7c, 32'hc4040db1, 32'hc3499cc5},
  {32'h44210b45, 32'hc23018e3, 32'hc4b4a324},
  {32'hc40f5264, 32'hc4b89bc1, 32'h44350cfb},
  {32'h43bbe44f, 32'h430c8920, 32'hc3bd7f13},
  {32'hc5602956, 32'h43d6a866, 32'h43af7a5a},
  {32'h4385deb0, 32'h435bbfce, 32'hc38a4b37},
  {32'h44b6d6f1, 32'hc4a82f01, 32'hc44623fa},
  {32'hc4d93dfa, 32'hc2e130ca, 32'h44a881fc},
  {32'h44aacb9f, 32'hc410c290, 32'h434d1adb},
  {32'hc4caee1f, 32'h444a6eb8, 32'h445092cc},
  {32'h446fe200, 32'hc4de4743, 32'h42aeb4af},
  {32'hc3a584d4, 32'h4407ffbf, 32'h437b9a3a},
  {32'h43dad19e, 32'hc38fa52f, 32'h437b1625},
  {32'hc48dbf10, 32'h4371d55b, 32'h434e99d7},
  {32'h44a3e282, 32'h4303331e, 32'h44280342},
  {32'h4411833c, 32'h44b1a98a, 32'hc3844bc5},
  {32'hc3f657d8, 32'hc501470a, 32'h43f6812e},
  {32'hc4702aac, 32'h43e74bb0, 32'hc2ad7f6f},
  {32'h43e9f27e, 32'h43261430, 32'h4510ef37},
  {32'hc4238477, 32'hc0bd5461, 32'hc50d585c},
  {32'h44627030, 32'hc1f8fbc6, 32'hc175768a},
  {32'hc396b2dc, 32'hc402729d, 32'hc5154254},
  {32'h45038227, 32'hc3ec63df, 32'h43c7084e},
  {32'hc4b5cb6a, 32'hc306592a, 32'hc41f7fbe},
  {32'h4439ac86, 32'hc47fe53c, 32'h44a1815a},
  {32'hc51f2582, 32'h44a4dff2, 32'hc3aaf5d7},
  {32'h44aa6b86, 32'hc3bc2d06, 32'hc2997950},
  {32'hc4a6cfb1, 32'h3f68d064, 32'hc3ea5256},
  {32'h452b1fd0, 32'hc40d85fb, 32'hc386c4b5},
  {32'hc2052130, 32'h44e96abc, 32'hc3a65c76},
  {32'h4518133e, 32'h4359b8cd, 32'h4417c691},
  {32'hc4100b96, 32'hc4000386, 32'hc5461b64},
  {32'hc4a5089c, 32'h41f62ff9, 32'h43521854},
  {32'hc465ec9a, 32'h448db7c6, 32'hc4b5ec64},
  {32'hc3459801, 32'hc4bf623a, 32'h44eb1ca5},
  {32'hc2b227f3, 32'hc2c37cd9, 32'hc21f28c9},
  {32'h4326d42c, 32'h43c1744d, 32'h42011b7c},
  {32'h4440d1b0, 32'h4255e67e, 32'h4321a22e},
  {32'hc48f169c, 32'h442fddf6, 32'hc3b103ef},
  {32'h4382da64, 32'hc3b6a4e7, 32'h41ee38d0},
  {32'hc5401837, 32'h43b11a6a, 32'hc3cccd5c},
  {32'hc1511740, 32'hc2272bf1, 32'h4548a695},
  {32'h44813b4a, 32'h44d101ca, 32'h4496ddc9},
  {32'h4433c5c4, 32'hc441621b, 32'hc4fc6418},
  {32'h44123fce, 32'hc3dac0af, 32'h43d0561d},
  {32'hc42fd58b, 32'hc41daee8, 32'h4384f9f9},
  {32'hc408812a, 32'h4287ed76, 32'hc4df3237},
  {32'h445ef235, 32'hc3112f4c, 32'h44d44e3c},
  {32'h44f74a21, 32'h43fbef71, 32'h434b2e58},
  {32'hc14762dc, 32'hc41edb61, 32'h4493cc0b},
  {32'h3f73ad00, 32'hc26e4aea, 32'hc541ac38},
  {32'hc3e85b69, 32'hc3635b8f, 32'h4369aa2a},
  {32'hc3d9b948, 32'h425be927, 32'h4352ccf6},
  {32'h44ff3bdf, 32'h44424199, 32'h44026df2},
  {32'h433c2560, 32'hc2c9b009, 32'h4378aacf},
  {32'h45223524, 32'hc44b6b7c, 32'hc3cb80d5},
  {32'h426915e5, 32'h45430fa3, 32'hc362a0ac},
  {32'hc3e61b4c, 32'hc3bfb37b, 32'hc3358093},
  {32'hc48066d1, 32'h44bc2c88, 32'hc4047c9c},
  {32'hc218ef86, 32'hc52541b8, 32'hc3d818e4},
  {32'h4413c915, 32'hc46c8c54, 32'h44039d4d},
  {32'h44de4824, 32'h4472ed97, 32'hc43152d7},
  {32'hc40bba88, 32'hc505e13b, 32'h44acdc14},
  {32'hc3ad9e2c, 32'hc50b5890, 32'hc23d2778},
  {32'h43c570dc, 32'h44d28bd5, 32'h430e1312},
  {32'h44be616b, 32'h42abfb07, 32'h43e64e55},
  {32'h4439247c, 32'h43510d4d, 32'hc4bfe5b9},
  {32'hc3a0335b, 32'hc3dd36ce, 32'h44f58895},
  {32'hc4ba45e4, 32'h43c170f6, 32'hc3bb7016},
  {32'hc40a48e5, 32'h440f2dad, 32'hc3cdc6ca},
  {32'h41e3e3e0, 32'h43b53b23, 32'h453dc1e1},
  {32'hc377dec3, 32'h4427ea86, 32'hc4e5ff42},
  {32'hc28ef9f2, 32'h434508fb, 32'hc5048f8c},
  {32'hc4947faf, 32'hc44f0c21, 32'h439d14a0},
  {32'h44fd6f8b, 32'hc2ad0c4d, 32'hc32f01bd},
  {32'hc3d15ab1, 32'hc48114e5, 32'h44aa628b},
  {32'hc284c8ea, 32'h44f1f3cf, 32'hc2a3366e},
  {32'h42d4fd1a, 32'hc489250d, 32'hc3d4c9aa},
  {32'h45414fd8, 32'hc3d4471a, 32'hc35f0c86},
  {32'hc558a7df, 32'hc388f0e2, 32'hc20999e0},
  {32'h4401652b, 32'h431e9ee9, 32'h4200a804},
  {32'hc45f544b, 32'hc4d55753, 32'h41e91841},
  {32'h44ce27be, 32'h43975bc3, 32'h41c3dbf1},
  {32'hc392e3d6, 32'hc324520b, 32'hc19c2cfc},
  {32'h44d26f6a, 32'h44c4ef28, 32'hc30aa4f9},
  {32'hc22fa2d0, 32'hc5300283, 32'h43ce321f},
  {32'h45476f70, 32'hc3ad4149, 32'h43b8cfff},
  {32'h42d48670, 32'hc4cea6e1, 32'h4411a982},
  {32'hc4611382, 32'hc40fac95, 32'hc42ab99c},
  {32'h430a8614, 32'h445bc9dd, 32'h4438d7b4},
  {32'hc49fb011, 32'h428ee6a9, 32'hc3c1efe6},
  {32'h411b1304, 32'h42b53549, 32'h45179658},
  {32'hc44fa0af, 32'hc4b00b23, 32'hc4223c53},
  {32'h447a3a9b, 32'h4315ecff, 32'hc28e2d32},
  {32'hc49b9872, 32'hc418692f, 32'hc4b64b52},
  {32'h43b81517, 32'h4451d9c4, 32'h455785a6},
  {32'h445475f1, 32'hc4120560, 32'hc33b07c6},
  {32'h437e5239, 32'hc5068b22, 32'h4509173b},
  {32'h43972823, 32'h44a12049, 32'hc44d0f8d},
  {32'h45233fd8, 32'h41d86d7c, 32'h41cecde8},
  {32'hc49fba9e, 32'hc3ddf3b2, 32'hc3d87026},
  {32'h43330bd4, 32'h43465998, 32'h450f2392},
  {32'h44ca36ea, 32'hc436b78c, 32'hc415662c},
  {32'h455f7437, 32'h43f1fca1, 32'hc3f4ffbb},
  {32'hc53a4ecd, 32'h4205d874, 32'hc3f29163},
  {32'h44bf3c60, 32'h442e0948, 32'h4353ff0c},
  {32'hc48f656b, 32'hc4745665, 32'h43dd95de},
  {32'h4317ad80, 32'h450ee5ad, 32'h44532f8e},
  {32'hc35b84bf, 32'hc4b20aba, 32'hc31c4909},
  {32'h4501430d, 32'hc2474aec, 32'h439cacc1},
  {32'hc44db6ec, 32'hc4bd047d, 32'h43a79fcc},
  {32'h4522b4f6, 32'h4399d090, 32'h436dbd3c},
  {32'hc3a97e84, 32'h4479dae6, 32'h42618bd7},
  {32'h44125208, 32'hc3a6e798, 32'h44090cdc},
  {32'h431e9cb3, 32'hc48b0f28, 32'hc3423b8e},
  {32'hc4e97832, 32'hc2aa3b37, 32'h445d82de},
  {32'h4331f3c6, 32'h4426ca4a, 32'hc4543128},
  {32'hc0ed9680, 32'h4429a9f4, 32'h451a4bf9},
  {32'h45216ef8, 32'hc31ce14b, 32'h441b1dd8},
  {32'hc48939b2, 32'h43b3f902, 32'h43ef2195},
  {32'hc29a63fd, 32'hc4c28d63, 32'hc4cbdc29},
  {32'hc4da2834, 32'h444a9b4e, 32'h441c1a89},
  {32'hc4ad8abe, 32'hc31deb7c, 32'hc21782ac},
  {32'hc48a932c, 32'h44a5cfa3, 32'hc3d75729},
  {32'hc30b8de4, 32'h44775480, 32'hc4cc86ae},
  {32'hc1db6db0, 32'h44e4cefb, 32'hc2ceb604},
  {32'hc333eb68, 32'hc4bfa574, 32'hc40c6fd7},
  {32'hc25075b0, 32'h44b05fc4, 32'h44b013b6},
  {32'h43b470be, 32'hc3153457, 32'hc465fe2e},
  {32'h448f4390, 32'h446ab203, 32'h454ad2a4},
  {32'h442e30b4, 32'hc3927bc8, 32'hc43c2600},
  {32'hc51fa587, 32'h42be5f34, 32'hc3db5c3b},
  {32'h44a9ebc6, 32'hc495842f, 32'hc3421ebc},
  {32'hc5410870, 32'h42e2a8b1, 32'h442522e8},
  {32'h42c4f430, 32'hc486f378, 32'hc3dc7238},
  {32'hc318f890, 32'h457b123a, 32'hc25e879a},
  {32'h44ea07dc, 32'hc41b787d, 32'h43ad98a3},
  {32'h439af4b4, 32'h443403f4, 32'hc288fa02},
  {32'h44bab7bb, 32'h43b3a785, 32'h43d90fe8},
  {32'hc49fa5a3, 32'hc3dae021, 32'hc1fc86bc},
  {32'hc4b010cc, 32'hc339a42a, 32'hc3a9f1d7},
  {32'h3ffd7750, 32'h431dec94, 32'h44c8abd3},
  {32'hc4b86998, 32'hc0e93d5b, 32'hc4b81406},
  {32'h449a5d65, 32'hc28f8492, 32'h4428ea43},
  {32'hc4fdc80c, 32'hc3b0942a, 32'hc3f51cf4},
  {32'h448bafbf, 32'hc4a04f09, 32'hc2a55c8b},
  {32'hc4f33274, 32'h442daf53, 32'h43974d3d},
  {32'hc4262c0e, 32'hc42eb269, 32'h3f22eea8},
  {32'hc44604b3, 32'h450197af, 32'h437c2393},
  {32'h449658c6, 32'hc4a22455, 32'hc404b024},
  {32'hc4a6a416, 32'hc3a1eef1, 32'hc3dcc00b},
  {32'h452aa583, 32'h4319e7d2, 32'h42023210},
  {32'hc22127f0, 32'h448642dd, 32'h4494cb28},
  {32'h43471220, 32'hc392e034, 32'hc4868ac8},
  {32'hc2742c58, 32'h438a0d48, 32'h43965fda},
  {32'h437d7351, 32'hc534b640, 32'hc388b225},
  {32'h44563580, 32'h4362d4ff, 32'h4383486c},
  {32'h44a1e203, 32'hc48bf490, 32'h4337e7d6},
  {32'hc5085f48, 32'hc3eadc9d, 32'h44283844},
  {32'h44a7617a, 32'h434c42b6, 32'h43fc99ed},
  {32'hc580c016, 32'h4293440e, 32'h43207cbd},
  {32'h440875b0, 32'h44507673, 32'hc4e10d2e},
  {32'h44b56362, 32'hc201b6ce, 32'h43f58b5e},
  {32'hc359561a, 32'hc50f6459, 32'hc46b234f},
  {32'hc5019e81, 32'h41f53526, 32'hc2b5bd26},
  {32'h4260a8f3, 32'hc4054e3f, 32'hc4717475},
  {32'hc528ab30, 32'h441ecbf7, 32'h439fafb6},
  {32'h44e5b631, 32'hc366c968, 32'hc47b0ed4},
  {32'h43a7c26c, 32'h412c1101, 32'hc4c009b4},
  {32'hc5625b00, 32'h431cb37d, 32'h42f00442},
  {32'h44f38f2c, 32'h439ae2eb, 32'h43e4f058},
  {32'hc51fb99f, 32'hc3d7f757, 32'hc36e9b90},
  {32'h44e18a42, 32'h43befecf, 32'hc3be57b1},
  {32'h43adc4fe, 32'hc40efcc2, 32'hc2a28c85},
  {32'h443ff4e8, 32'h44eb48dc, 32'h429f5e32},
  {32'hc55f1bc2, 32'hc30e2c8c, 32'h43345384},
  {32'h43ed16f4, 32'h44c54328, 32'h43477d3f},
  {32'hc3e72b88, 32'hc3eaf22c, 32'h43be0afd},
  {32'h4460f1c8, 32'h4421d975, 32'h442e7949},
  {32'hc4becb12, 32'hc2be5391, 32'hc167e7d2},
  {32'hc197c980, 32'h4422be46, 32'h44ecd5c1},
  {32'hc473b0a4, 32'hc2ad6970, 32'hc502e050},
  {32'h44342d50, 32'h428e179e, 32'h437ca8a2},
  {32'hc4b8a053, 32'hc3c2238c, 32'hc4ac3879},
  {32'h43a5b1ac, 32'h452e3aee, 32'h43f12d3f},
  {32'hc3d2b48f, 32'hc3084979, 32'hc41626e3},
  {32'h442d44a8, 32'h440c1e11, 32'h4431e1b4},
  {32'hc5672a94, 32'hc2f6ff3e, 32'hc358c362},
  {32'hc4e3e648, 32'h413ea5b8, 32'h3fc0b780},
  {32'hc374e880, 32'hc4a9e100, 32'hc3a73b42},
  {32'h436e3b7e, 32'h45300ebb, 32'h4293ed86},
  {32'hc44500e8, 32'hc3fdbeb3, 32'hc40c7916},
  {32'h440608c6, 32'h43f120c7, 32'h44dac23c},
  {32'hc4aee930, 32'hc4649e47, 32'hc43f30cd},
  {32'h452446a4, 32'hc3a1b4ff, 32'hc34f910d},
  {32'h4426f180, 32'h43bbfb0c, 32'hc4093032},
  {32'hc48a7bea, 32'hc44decf4, 32'hc31fdc6b},
  {32'hc1e27160, 32'h44ebaf4d, 32'h440546d8},
  {32'h44bb9e44, 32'h40a324b2, 32'h43bbee4d},
  {32'h44e5b477, 32'h43f6e136, 32'hc3920ada},
  {32'hc5320eb8, 32'hc395bd81, 32'hc31a58fe},
  {32'h44921f06, 32'hc2a45a46, 32'hc4478382},
  {32'hc4947642, 32'hc386e718, 32'hc353bd67},
  {32'h4503d731, 32'h437f96cc, 32'h425d0768},
  {32'h442345ae, 32'hc2b395b8, 32'h4390e307},
  {32'h44ef5317, 32'hc32bc0ce, 32'hc3d30d30},
  {32'hc4fd41d1, 32'hc2111e44, 32'hc36c63fe},
  {32'hc3b8540c, 32'h4445ee2f, 32'hc28d025e},
  {32'hc32b0617, 32'hc3f3b208, 32'h44d8e65c},
  {32'h433e5922, 32'h436c6c98, 32'hc5270bb7},
  {32'hc474471c, 32'hc3266c6b, 32'h43f67850},
  {32'h4493b818, 32'h43c6faff, 32'hc4f4e6b6},
  {32'hc4190f52, 32'hc40f76c4, 32'h44348bf6},
  {32'hc3fa2790, 32'h430f574c, 32'hc42b9719},
  {32'hc416ac76, 32'hc4a0c3ef, 32'h443cfe42},
  {32'h443a179c, 32'h452217db, 32'hc1311392},
  {32'hc3b303fe, 32'hc33a6c85, 32'hc36bfc2a},
  {32'h44ed8b1d, 32'hc326256c, 32'hc3f3f134},
  {32'hc2f2b93c, 32'hc549a3ef, 32'h4343d88c},
  {32'h454f28db, 32'h43238ede, 32'h403035d8},
  {32'hc5143e3f, 32'h4401c3c7, 32'h44601c6e},
  {32'h44a0d326, 32'hc3e1758c, 32'hc4fdade8},
  {32'h44552952, 32'hc3a0f344, 32'hc46ca77d},
  {32'hc5598d40, 32'h426cd482, 32'h43add5de},
  {32'h43ab4d3d, 32'hc5274da8, 32'hc22e1e1a},
  {32'hc48346f8, 32'hc390c80b, 32'h41a804c6},
  {32'h44f4dae0, 32'hc35ba175, 32'h42130ca8},
  {32'hc454aef9, 32'h4418688f, 32'h43d93a54},
  {32'h454fc56b, 32'hc2e62446, 32'hc41604f5},
  {32'hc505f493, 32'hc3886c82, 32'hc2a01b9b},
  {32'hc44f9c97, 32'hc3d5e079, 32'h43e08040},
  {32'hc4b49172, 32'h4375ca6e, 32'hc2f501df},
  {32'h45190f7d, 32'h432c9ca8, 32'h438d0fa0},
  {32'hc3fd4052, 32'h4394e6da, 32'hc405290a},
  {32'h422f6b73, 32'hc39b2315, 32'h41c07a92},
  {32'h41f58dd0, 32'h440d283c, 32'hc48a164f},
  {32'h448ea772, 32'hc18d6d9c, 32'h43e518ce},
  {32'hc51b9338, 32'h443b96e1, 32'h43984720},
  {32'h443abade, 32'hc40f8a84, 32'h438ede82},
  {32'hc4169e89, 32'h43ab0d11, 32'hc3b9e0ff},
  {32'h4315debf, 32'hc4aa8e70, 32'h440e1c26},
  {32'hc56772aa, 32'h439d9c27, 32'hc3798522},
  {32'hc2f49a42, 32'hc475117e, 32'h42729bae},
  {32'hc3852f0f, 32'h430d8626, 32'hc54350fc},
  {32'h454adf84, 32'h443afcbb, 32'h432ab576},
  {32'hc3c4dfb8, 32'hc20cb4cb, 32'hc2e57286},
  {32'h4460b580, 32'hc2e27ec2, 32'h44aed44d},
  {32'hc5493b05, 32'h424989b3, 32'hc445b717},
  {32'hc44b1e3c, 32'h4232cd91, 32'h43e14962},
  {32'hc516a274, 32'hc40ed568, 32'hc3bde2ad},
  {32'h438c0144, 32'h44f611fa, 32'h44b8dd19},
  {32'hc4bbb567, 32'hc439eb31, 32'h4328a200},
  {32'h437428c1, 32'h44a80139, 32'h433e8b03},
  {32'h42bf2f8c, 32'h43651984, 32'h450afbe2},
  {32'h438f56f2, 32'h4547f3a5, 32'h43b32c5a},
  {32'h43ce3e91, 32'hc456f182, 32'h43e2663c},
  {32'h439b3cbd, 32'h44f0f61e, 32'hc4320aa7},
  {32'h44b13864, 32'hc2a27744, 32'h445813fd},
  {32'h451402ae, 32'hc3d1c80e, 32'h447b1efa},
  {32'h4339e758, 32'h4330e58b, 32'hc5169f94},
  {32'h4486804a, 32'hc3bd97c2, 32'hc3910a15},
  {32'h442a0ed9, 32'hc467e197, 32'h44467f75},
  {32'hc4847ac1, 32'hc332b1a5, 32'hc4bf832a},
  {32'hc14d79d0, 32'hc389ee1e, 32'h452b6610},
  {32'h43b81046, 32'h44472237, 32'h42c16a15},
  {32'h443f1c1f, 32'hc439f587, 32'h44bd730b},
  {32'h439900c4, 32'hc3aeea06, 32'hc553b864},
  {32'hc4b7c125, 32'hc34bf87d, 32'h43b031d8},
  {32'hc4e270e7, 32'hc2ad5694, 32'h42a7db84},
  {32'h4211b040, 32'h435992ea, 32'hc3442b01},
  {32'hc51ba0eb, 32'hc399bd6e, 32'hc3d6a28a},
  {32'h447102d4, 32'hc4bfac7f, 32'hc3567c48},
  {32'hc4cbcec1, 32'h443de6d7, 32'h42b29bde},
  {32'h4403a960, 32'h42e65bd2, 32'h42818d7a},
  {32'hc568d7ca, 32'hc3b4d8a3, 32'hc3b4df94},
  {32'hc3a58cce, 32'hc522fa96, 32'hc2e588c9},
  {32'hc4ab8d14, 32'h41111e54, 32'hc33303b5},
  {32'hc1130438, 32'hc42a2e76, 32'hc4c103b2},
  {32'hc4dc2f52, 32'h419843be, 32'h41284bf3},
  {32'hc3a3a390, 32'h42bb894c, 32'h45061492},
  {32'h440bb9c6, 32'h454eac64, 32'h440e54a9},
  {32'h40beee80, 32'hc2aa7a9a, 32'h450753f4},
  {32'h44531284, 32'h43d1dfa6, 32'hc4a0f1cd},
  {32'hc5455f92, 32'h427168cf, 32'hc16679c3},
  {32'hc48c7880, 32'h4217892a, 32'hc4207a32},
  {32'h440fed29, 32'hc3b8bab8, 32'hc40d7afe},
  {32'h42b74608, 32'hc4c0db55, 32'h4547d28a},
  {32'h42183240, 32'hc4a8c8ca, 32'hc4d939aa},
  {32'h44496490, 32'h44426f1c, 32'hc45193da},
  {32'h3fc83100, 32'hc3d154e0, 32'h45492670},
  {32'h44796460, 32'h4442e874, 32'hc4267ee4},
  {32'hc5421dbc, 32'hc3079fb6, 32'h41152b30},
  {32'h415d6e00, 32'h4499fae5, 32'hc3d731f2},
  {32'hc4d00cd7, 32'hc29e4d33, 32'h431c3d5b},
  {32'h44b53aed, 32'h43ce0dad, 32'hc35dfc71},
  {32'hc558c610, 32'h433b38d5, 32'h4316d14e},
  {32'hc4f6f7de, 32'h4313c0e2, 32'h411d4a3d},
  {32'hc43925cc, 32'hc48d0f0b, 32'h429ec564},
  {32'h4247f0d6, 32'h4550c289, 32'hc2a7857c},
  {32'hc3508d3c, 32'hc4b26496, 32'h42748390},
  {32'h44afeee6, 32'h4463a7b1, 32'hc35b9b16},
  {32'hc2c1a5dd, 32'hc53ad327, 32'hc329079c},
  {32'hc2a87fad, 32'hc33fe7c0, 32'hc3b5cad9},
  {32'hc3320d7d, 32'h444756f1, 32'hc2e531e2},
  {32'h43fb58e6, 32'h43b01393, 32'hc4c38e49},
  {32'hc2be9ab0, 32'h4371ad8c, 32'h44bc85a4},
  {32'hc0288e00, 32'h4264b41e, 32'hc4e3db88},
  {32'hc40704cc, 32'h423779dc, 32'hc2b28ab5},
  {32'h433d14bf, 32'hc48f9826, 32'hc470dc6d},
  {32'hc49f76be, 32'hc3112ca7, 32'h43761ce7},
  {32'hc4ce0730, 32'hc4217261, 32'hc424f53f},
  {32'h43081b20, 32'hc3a57476, 32'h445653df},
  {32'h42657e40, 32'h442d29c4, 32'hc3a877b8},
  {32'hc43a4dd4, 32'hc470c0c0, 32'h44fba496},
  {32'hc43050ff, 32'hc341bd12, 32'hc46a3c19},
  {32'h43e57731, 32'h4441dff8, 32'h437a06bd},
  {32'hc4961dcd, 32'hc46cae4f, 32'hc395e890},
  {32'h441d6810, 32'h438b408d, 32'h45171448},
  {32'h44316399, 32'hc4182642, 32'hc4c7e5fb},
  {32'hc4074630, 32'h450123c6, 32'h44f4669d},
  {32'h4292219f, 32'hc1daafdf, 32'hc536d325},
  {32'h42961e10, 32'h441588f6, 32'h43d86739},
  {32'hc4d6ddc2, 32'hc4af80cd, 32'h436c7849},
  {32'h440e606f, 32'h45230f9a, 32'hc3a4b348},
  {32'hc3800b94, 32'hc4b516c0, 32'h43efb7cc},
  {32'hc3989b00, 32'h45850dd6, 32'hc207e0e7},
  {32'hc2fe5938, 32'hc5365ba7, 32'h42fb0b9b},
  {32'h44ced869, 32'h431ecc9a, 32'h42d69cf4},
  {32'hc58152ca, 32'h42143122, 32'hc2802ada},
  {32'h451ef627, 32'hc31e5785, 32'h44369ac5},
  {32'hc33414cb, 32'h43c5d3cc, 32'hc4f6f593},
  {32'hc3c681ca, 32'h42ec9c77, 32'h447d219c},
  {32'h435c0bb4, 32'hc40dcce2, 32'hc3589a72},
  {32'hc432d4b0, 32'h40889be4, 32'h44ea0a7f},
  {32'h4520ef26, 32'hc39408c3, 32'hc25fa6af},
  {32'hc3484b95, 32'hc378d186, 32'h4425bbdb},
  {32'h44878b2e, 32'hc459a358, 32'hc4b57a80},
  {32'hc421e566, 32'h4445ece3, 32'h447b365a},
  {32'h45318ac6, 32'h411506b6, 32'h42423552},
  {32'h42d7bd8d, 32'hc3bf46e0, 32'h44f1cdd6},
  {32'h44222d63, 32'h43c7e7e7, 32'hc3c8976e},
  {32'hc4e7324d, 32'h43ffd63c, 32'h42577518},
  {32'h44f5f751, 32'h42ebcce2, 32'hc33612b2},
  {32'hc30dcb0e, 32'h428b0bf3, 32'h451554dc},
  {32'h4504d59d, 32'hc3838407, 32'hc3e776d3},
  {32'hc4ac711e, 32'h4412b592, 32'h4438fa6f},
  {32'h4428fafe, 32'hc308b57c, 32'hc4044168},
  {32'hc500cd04, 32'h43cbe766, 32'h43635c1f},
  {32'h450f32df, 32'hc420c6d3, 32'h42a613d9},
  {32'hc45e0988, 32'h451d1a17, 32'h4391bdd2},
  {32'h442f5f87, 32'hc35054a2, 32'hc385753f},
  {32'hc325a8b0, 32'h435c7808, 32'h42bf13a7},
  {32'hc19fdc4c, 32'hc501ae77, 32'hc2736810},
  {32'h4279de40, 32'h449871b0, 32'hc39a9e07},
  {32'h457636d8, 32'h43e737da, 32'h4231e1fd},
  {32'hc4edbce0, 32'h442eff7b, 32'hc3421e83},
  {32'h441d7b68, 32'hc33c22ed, 32'hc3a8edf7},
  {32'hc4d0e1c3, 32'hc32b35fd, 32'hc21b6e7c},
  {32'hc49bd4fe, 32'hc3924a9c, 32'hc499fd21},
  {32'hc3482390, 32'hc42a31e2, 32'h4486a0c8},
  {32'hc4b45a0b, 32'h437743be, 32'h4303b3c7},
  {32'h44a1c287, 32'hc4d6452d, 32'hc221e5c1},
  {32'hc3af87de, 32'h457112d3, 32'h4392d42a},
  {32'h451e8e63, 32'h420acd10, 32'h431f2b40},
  {32'hc4ba6c2d, 32'h44d656b9, 32'h434e8a0d},
  {32'h449aab49, 32'hc4b8bbaf, 32'hc21408fa},
  {32'h4355f7e0, 32'hc3f9b692, 32'hc3c37f30},
  {32'h44c32b53, 32'h437df3c4, 32'h43343a0c},
  {32'hc4617af6, 32'h43e375f6, 32'hc49dd79b},
  {32'hc3710630, 32'hc2c64f06, 32'hc46ba840},
  {32'h4397b49c, 32'h456381c7, 32'h43bffc45},
  {32'h44550336, 32'hc311b3bc, 32'hc41067a9},
  {32'hc46050dc, 32'h43372538, 32'h42ba4688},
  {32'hc3f857c0, 32'hc1361d56, 32'hc520d960},
  {32'hc3d62f76, 32'h444f6ff0, 32'h4494b5d9},
  {32'hc4b47b5b, 32'hc3842c63, 32'hc32eebad},
  {32'hc51f83a8, 32'hc447cb72, 32'h42ae2644},
  {32'h449da0db, 32'hc1bc7636, 32'hc44e0cba},
  {32'hc3fd5d72, 32'hc3ebfa50, 32'h437345af},
  {32'h4510263d, 32'hc20d65ed, 32'hc41c5881},
  {32'hc43fb064, 32'h44093e64, 32'h43ec26d7},
  {32'h4398ae0a, 32'hc15d0894, 32'hc3275dbc},
  {32'hc15c0cc0, 32'h44434688, 32'h4503a021},
  {32'h42d9ac28, 32'hc3f106a8, 32'hc511007d},
  {32'h443573e0, 32'hc30ab51d, 32'hc48166bb},
  {32'hc5288071, 32'hc3770c9e, 32'h449f6a29},
  {32'h4432f554, 32'h40c2b0b9, 32'hc4417cbf},
  {32'hc43a0dac, 32'hc4f2f0a4, 32'hc34e3507},
  {32'h43dcf9f4, 32'h44d73b28, 32'h433ddc6b},
  {32'hc49eca45, 32'hc26c7b9f, 32'hc33181b7},
  {32'h441a760a, 32'h4529336f, 32'hc29bd298},
  {32'hc3e79e49, 32'hc530ba7c, 32'hc346f6ba},
  {32'hc3bd7390, 32'hc2834a5d, 32'h427269e2},
  {32'hc4c3c78e, 32'hc3f31d59, 32'hc28a2a4d},
  {32'h4448ff49, 32'h437dfa20, 32'hc47b19a0},
  {32'hc46d6948, 32'hc3670a72, 32'hc2bef64b},
  {32'h43bd64f8, 32'h44c4e707, 32'h43e44465},
  {32'hc3c6bd56, 32'hc53ced2e, 32'hc3863c88},
  {32'hc30eb573, 32'h44c90aeb, 32'h42b6c813},
  {32'hc3e33f76, 32'hc3157686, 32'hc54f53f2},
  {32'h44c676b3, 32'h44670f6b, 32'h44222a06},
  {32'hc2682b30, 32'hc4a52254, 32'hc3a9833d},
  {32'h4450ff06, 32'h44817a5c, 32'h4495ac98},
  {32'hc4707a1a, 32'h448351d1, 32'hc3eaf7fd},
  {32'hc31fc4fd, 32'h4470af42, 32'h43963248},
  {32'hc51acf28, 32'hc449b65b, 32'hc320f8c4},
  {32'hc24c2810, 32'h428cdaed, 32'h4521c37d},
  {32'hc5157c66, 32'hc39e2241, 32'h439f889b},
  {32'h42c002ee, 32'h4526a270, 32'h436c2e61},
  {32'h43a93c68, 32'hc5218f19, 32'hc323c31f},
  {32'hc42edb66, 32'h42a9a7de, 32'hc3998d78},
  {32'hc4b22ebe, 32'hc39c6cbe, 32'h430a9c68},
  {32'hc42d8abe, 32'hc49f03c5, 32'h43df1c08},
  {32'hc1d5f838, 32'h456a7edb, 32'h4365804b},
  {32'h448956df, 32'hc4194a55, 32'h43834520},
  {32'h43b6beaa, 32'hc31751ea, 32'hc3a64866},
  {32'hc535ec94, 32'hc38758fc, 32'h431b0220},
  {32'hc47f968e, 32'hc390b642, 32'h430a7926},
  {32'hc50c2704, 32'h442e5164, 32'h42968c55},
  {32'h4499fbbe, 32'h4454983c, 32'h442b2b6f},
  {32'h441f1036, 32'hc417b03b, 32'h44001bec},
  {32'h451595e0, 32'h43f1d104, 32'hc2662e9f},
  {32'hc33860f7, 32'hc4e88786, 32'hc1c7a152},
  {32'hc2bb3058, 32'h43b4c5fc, 32'hc3dfb88b},
  {32'hc44ddd9d, 32'hc3d48dfb, 32'h4445e25c},
  {32'hc3d4ac24, 32'h44673b78, 32'hc499e0d8},
  {32'hc3a960d6, 32'h42dd0741, 32'h443f1382},
  {32'h44f0e84d, 32'h42cf10e3, 32'hc1f9f6b0},
  {32'hc433532a, 32'h42a10600, 32'h44b5918f},
  {32'hc28b4abf, 32'h440d89b5, 32'hc4bd539a},
  {32'hc422ecb0, 32'hc4f5b2a9, 32'hc38d4bc3},
  {32'hc2d55558, 32'h4510f765, 32'hc37ba285},
  {32'hc43895e6, 32'hc2b477b6, 32'h440f637a},
  {32'hc2fa07ea, 32'h431bd6ec, 32'hc51d291c},
  {32'hc433f411, 32'hc4fe1e4f, 32'hc432b744},
  {32'h44b1041a, 32'h4398786e, 32'hc455c874},
  {32'hc5964d64, 32'hc38a925d, 32'h43b78a1e},
  {32'h44eadd83, 32'h42602fbb, 32'hc481c486},
  {32'h431d2708, 32'hc5394ef6, 32'h4285f72c},
  {32'hc36bb730, 32'hc386c486, 32'h4501f0e6},
  {32'hc48afb10, 32'hc40f5615, 32'hc32e1002},
  {32'h42b21d2d, 32'h45210401, 32'hc3249b60},
  {32'h448302d6, 32'hc4d39a32, 32'h42063949},
  {32'hc5045913, 32'h42f7a566, 32'hc3c246b8},
  {32'h44e4109e, 32'h443ace48, 32'h427e3524},
  {32'hc56e310b, 32'hc311c5d4, 32'h43d416b8},
  {32'h45619dff, 32'h43545abe, 32'h44156b2a},
  {32'hc4a90ab9, 32'h4448ba4f, 32'h41a25319},
  {32'h44b80b6a, 32'h438d875f, 32'hc4037df4},
  {32'hc442972d, 32'h4357854e, 32'hc48a7333},
  {32'hc201a5b8, 32'hc541c484, 32'h4325d6df},
  {32'hc2aa5abc, 32'h453d16d4, 32'hc398a4d0},
  {32'hc39a00a7, 32'hc4a351bd, 32'h43b0db35},
  {32'hc43fd7ab, 32'hc34abd50, 32'hc4e78b78},
  {32'h44aa3595, 32'h43351587, 32'h441bf9ce},
  {32'hc5305ed8, 32'h443439c1, 32'hc2b25c4d},
  {32'h43870b2c, 32'hc42241ac, 32'h45084ee2},
  {32'hc56f7e2c, 32'h434ad350, 32'hc390644b},
  {32'h4295253a, 32'hc4a0353d, 32'hc1c5eeea},
  {32'hc2ce38f0, 32'hc37e37c9, 32'hc54944aa},
  {32'h450dc955, 32'hc42bfca7, 32'hc405cb3f},
  {32'h43b2102e, 32'h43c6c8c7, 32'hc49ac98a},
  {32'h44eb9da7, 32'hc1c0d41a, 32'h446cb8c0},
  {32'hc48129ea, 32'hc350c8af, 32'hc544a4d8},
  {32'h446c3384, 32'hc28f53f9, 32'h441314ab},
  {32'hc3611bb2, 32'h440215bc, 32'hc4a4ea92},
  {32'h44916a8c, 32'h4445abab, 32'h447e3f00},
  {32'hc40844e2, 32'hc28547dd, 32'h43829355},
  {32'h43ac60d9, 32'h44508b5c, 32'hc3e314bd},
  {32'h45372c77, 32'hc39b29fa, 32'h4429de44},
  {32'hc34aaab4, 32'h450be92a, 32'h4407263d},
  {32'h44770806, 32'h42069882, 32'hc345ab9f},
  {32'hc415608c, 32'h44e771be, 32'hc49286ed},
  {32'h43168eb7, 32'hc390b154, 32'h443eab75},
  {32'h43e5841a, 32'hc487b4d4, 32'h44d5b137},
  {32'h44167a88, 32'hc443d337, 32'hc4cd3b97},
  {32'hc3aba89c, 32'h41ada468, 32'h43c945a2},
  {32'h43da1ab5, 32'h437b0a4e, 32'h449ceb38},
  {32'hc3b39cbe, 32'h4498ce72, 32'hc3ba16de},
  {32'h441074a4, 32'hc3ff5c16, 32'h420b1028},
  {32'h441ea15b, 32'h430bc635, 32'hc3f262b9},
  {32'h451461dc, 32'h42db0668, 32'h44319417},
  {32'hc3161300, 32'h4402e09f, 32'hc40ca83e},
  {32'h455fdb2d, 32'hc3f65593, 32'h44319695},
  {32'hc4b301a7, 32'hc296340a, 32'hc3f0dd2c},
  {32'hc427a204, 32'h441b139d, 32'hc2c2ac5f},
  {32'h44a3064a, 32'hc36c78a2, 32'h430dbf72},
  {32'h4494a35e, 32'hc47e9689, 32'hc428e691},
  {32'hc4c66af0, 32'h4437633e, 32'h43460ac9},
  {32'h44a1d06c, 32'h439a51db, 32'hc35310ee},
  {32'hc5880f4d, 32'h425a6269, 32'h439ccfc6},
  {32'h43ab467c, 32'hc5483b27, 32'hc3f40865},
  {32'h4474b074, 32'h44836030, 32'h43e27032},
  {32'h4180f820, 32'h449ff43f, 32'hc4a3f585},
  {32'hc3b0e3c4, 32'h43e95406, 32'h4483d148},
  {32'hc4a9d8e7, 32'hc384b324, 32'h442559e9},
  {32'h45116c8e, 32'h43ae0860, 32'hc2a72dd8},
  {32'hc25ab668, 32'hc49d8d9f, 32'hc35cfeb0},
  {32'h4417d936, 32'h43f86125, 32'hc4a69409},
  {32'hc3c11106, 32'hc22cfcc3, 32'h4523c2c3},
  {32'h433353ab, 32'h44381b59, 32'h4250662e},
  {32'h439fa7d5, 32'h444ea0a5, 32'hc3b75748},
  {32'hc426bf01, 32'h43018b24, 32'h44b52faa},
  {32'h451ede37, 32'hc2e27ffd, 32'hc481bcf0},
  {32'h43be38ec, 32'h44408fba, 32'hc3d06c92},
  {32'hc4818fce, 32'hc435b661, 32'h43acefe8},
  {32'hc34976d8, 32'h41f0375f, 32'hc43f39a4},
  {32'hc3e89425, 32'hc398938d, 32'h4524d684},
  {32'hc24300b0, 32'h45277fe1, 32'hc3dcc138},
  {32'h43d909ab, 32'hc3d6eaf3, 32'h44e6f36e},
  {32'h44673f74, 32'h433266a8, 32'hc3fecbe3},
  {32'hc53b3358, 32'hc12d89fb, 32'hc363ef70},
  {32'h436bca84, 32'hc3adc0f3, 32'hc3e04907},
  {32'hc5294707, 32'hc4515b84, 32'hc14d148b},
  {32'h45329d1d, 32'h43973784, 32'h436e93df},
  {32'hc4856242, 32'hc3a3e04e, 32'h43ea761b},
  {32'h447ef808, 32'h44bee2ca, 32'h4373dd6e},
  {32'hc5888496, 32'h42cfb0ad, 32'h417e1d7e},
  {32'hc3afeb32, 32'h43bb108b, 32'hc3eff3ab},
  {32'h41a62718, 32'hc43fc848, 32'h44c2240f},
  {32'h4390419f, 32'hc4cb79e4, 32'hc31a648a},
  {32'h43ef9090, 32'h44bd34ac, 32'h43d20269},
  {32'hc502187d, 32'h430f1663, 32'hc30cd527},
  {32'h44d8a9e6, 32'hc3385efa, 32'h4413d4f3},
  {32'hc48fdee1, 32'hc38d5fca, 32'hc4249f95},
  {32'h44acc5f7, 32'h443aa293, 32'h4322256e},
  {32'hc4067d68, 32'hc3e2822c, 32'hc4ded5b1},
  {32'h44a5e950, 32'hc2ea0a1c, 32'h448a102f},
  {32'h42caf387, 32'h44a8f46a, 32'hc384fa11},
  {32'hc3a8f1de, 32'hc2d6e5f9, 32'h44b8e6ac},
  {32'hc42960a7, 32'hc3bcd0c4, 32'hc484a774},
  {32'h4475a2a2, 32'h43a7a9c1, 32'h4386e2d1},
  {32'hc4d9292f, 32'hc41ed041, 32'h41b01bee},
  {32'h44b1deef, 32'h44248565, 32'h42f81035},
  {32'hc486c805, 32'hc395c7df, 32'h437343fe},
  {32'h44faebba, 32'hc2c980a3, 32'h430fde3a},
  {32'hc53553eb, 32'hc3aad8e9, 32'h413010a0},
  {32'h43ec64df, 32'h44bd51a8, 32'h428047e6},
  {32'hc52137a2, 32'hc3a05564, 32'hc342a2bc},
  {32'h440894ca, 32'h4519e49b, 32'hc3962a3c},
  {32'hc4d709d3, 32'h4226b065, 32'hc3bc86a4},
  {32'h44aa5061, 32'h448fc751, 32'h42fd89c5},
  {32'hc483d0a5, 32'hc4ac0f3f, 32'h421ab18a},
  {32'h4288a15c, 32'h43e56d4f, 32'h43b857be},
  {32'hc57dee6f, 32'h43840f32, 32'h4326204a},
  {32'h42bd9313, 32'hc2beb564, 32'h43f3facc},
  {32'hc336ca16, 32'h442f1808, 32'hc3cf24e0},
  {32'h41589bd4, 32'h43b68006, 32'h44d9bb0d},
  {32'hc44976fd, 32'h4449429b, 32'hc41ec22b},
  {32'hc41974b5, 32'h42258d5a, 32'h450b2885},
  {32'h4511bc84, 32'hc36b805c, 32'h425fea8d},
  {32'hc45a4f06, 32'h4393c1ca, 32'h441394dd},
  {32'h40ea8300, 32'hc43bacd9, 32'hc512b707},
  {32'hc3e779b8, 32'h431f9b6c, 32'h449f3396},
  {32'h4528bb65, 32'h42b38228, 32'h434acd50},
  {32'h438892af, 32'h44e15aa2, 32'h442abcae},
  {32'hc3b685e2, 32'h449e83e0, 32'hc4d37b53},
  {32'hc1010284, 32'hc4c2efba, 32'h444d83a4},
  {32'hc3738962, 32'hc34ecc7e, 32'hc52623df},
  {32'hc4cdb4d8, 32'h43b143a8, 32'h4323875c},
  {32'hc24aa161, 32'h43492b85, 32'hc48d8a8a},
  {32'hc24cd7be, 32'h4335003a, 32'h4510aec1},
  {32'hc3e82dbe, 32'hc325a75f, 32'hc4a962d5},
  {32'h44de4858, 32'h40f8d2d8, 32'h434beb59},
  {32'h43ce8db0, 32'hc4f87d42, 32'hc3b22a63},
  {32'hc5110167, 32'h441dbd34, 32'h42bae4c7},
  {32'hc419c906, 32'hc48d31f3, 32'hc2078f86},
  {32'hc40ac34d, 32'h44b22d09, 32'hc37ab612},
  {32'h43aa7b28, 32'hc48be26f, 32'hc3c5dba8},
  {32'hc533b188, 32'hc25cf66d, 32'hc2c837b0},
  {32'h451bedcc, 32'h43ed9f14, 32'hc2f4a197},
  {32'hc5235177, 32'h43f27daa, 32'h4436c352},
  {32'h45576fc7, 32'hc2bcb5ef, 32'h43b716b8},
  {32'h441f71bc, 32'h42b8f06f, 32'h445e314c},
  {32'hc5351c74, 32'h42feb560, 32'hc3593ed5},
  {32'h43d19cda, 32'h43251f3a, 32'h45336834},
  {32'h4472051b, 32'h440fce17, 32'h4376c55d},
  {32'h430643e2, 32'hc51cd28f, 32'hc1912bd7},
  {32'h41979200, 32'h44d49537, 32'h4406e5c9},
  {32'h450760b4, 32'h4411aa5e, 32'hc23b50d5},
  {32'hc503dbd9, 32'h43c9e774, 32'h41a37f39},
  {32'hc1a749c0, 32'hc569e7c8, 32'hc37ae3d1},
  {32'hc52071ba, 32'hc24097b6, 32'hc2001228},
  {32'h4440b202, 32'h444510f5, 32'hc49a9b6b},
  {32'hc487ad4a, 32'hc1edd7c0, 32'hc483ca01},
  {32'h438d603e, 32'hc3952658, 32'hc3b1179f},
  {32'hc400b18a, 32'h4336884d, 32'h438e9c9a},
  {32'h438aed58, 32'hc450d1e9, 32'hc3dbd5bf},
  {32'hc409e9fa, 32'h43afb7e5, 32'h4338ba1f},
  {32'hc4113b7a, 32'hc3c922da, 32'hc4d51ad6},
  {32'hc3066011, 32'h453b3018, 32'hc3481d8c},
  {32'h449c4e8e, 32'h42eb53ee, 32'hc412f707},
  {32'hc334eca8, 32'h4434db8c, 32'h4485ebf7},
  {32'h454184f1, 32'h42934834, 32'hc3df1241},
  {32'h439fae93, 32'h44d6dba8, 32'hc39696ce},
  {32'hc40abc88, 32'hc290bad6, 32'hc51f85ed},
  {32'h42bf1120, 32'h44067b35, 32'h44cc9337},
  {32'h4474e934, 32'hc4115290, 32'hc3b87c96},
  {32'hc516c06a, 32'h440b32e7, 32'hc1e1cc15},
  {32'h43f2911e, 32'hc4dce4e9, 32'hc44d85c3},
  {32'h44f020d3, 32'h43318512, 32'hc43badd2},
  {32'hc506de01, 32'h4316f2b8, 32'h448651fe},
  {32'h43f409fa, 32'h447436d5, 32'hc495d4b8},
  {32'hc4a97f18, 32'hc48f20ff, 32'h410d54ec},
  {32'h4546089f, 32'hc34cd6a2, 32'hc3876605},
  {32'h433a11c5, 32'hc514f319, 32'hc3c55b1a},
  {32'h446c8950, 32'h4517007d, 32'h43e0bb09},
  {32'hc4d2e2bf, 32'hc49430b8, 32'h4413930f},
  {32'hc4179ff6, 32'hc356b288, 32'h439111fa},
  {32'hc467d9f1, 32'hc2e89642, 32'hc3cc9cb2},
  {32'h446b6620, 32'hc33036c0, 32'h4426787d},
  {32'hc37a0210, 32'hc4357774, 32'h44bbcbae},
  {32'hc2df10b6, 32'h435bbe8c, 32'h45058d4f},
  {32'hc35a97c3, 32'hc4d5daa2, 32'h43278bf3},
  {32'hc5108f76, 32'h42df93ed, 32'h4310ed5a},
  {32'hc4d5275e, 32'hc38f658a, 32'hc43cfda2},
  {32'h44e59892, 32'h441c4895, 32'h43f51f07},
  {32'h44a70422, 32'h4344d217, 32'hc42ae333},
  {32'h45307190, 32'h42033b47, 32'h43af4de0},
  {32'hc56a6fb3, 32'h428f0eb5, 32'hc3d5f6da},
  {32'hc42e01d7, 32'h43ec27a3, 32'h429ac588},
  {32'h42a358f0, 32'hc449acbc, 32'hc40a74e9},
  {32'h439bab5a, 32'h4397377e, 32'h442b27e2},
  {32'h446930a8, 32'h429c21e4, 32'hc4421f6c},
  {32'h43ec1c78, 32'h44177cf5, 32'h444bfd84},
  {32'h4383adcc, 32'hc3ec9a16, 32'hc547af1b},
  {32'hc322a596, 32'hc341f6d7, 32'h43ff7184},
  {32'h44ab7036, 32'h41c41198, 32'hc3b5a687},
  {32'hc381eca6, 32'hc4ebc2e9, 32'hc3a774d5},
  {32'hc279f800, 32'h44e45014, 32'h4443a414},
  {32'hc2b4eec8, 32'hc403007f, 32'hc247849e},
  {32'h43b748f9, 32'h452a5a54, 32'hc33b258e},
  {32'hc3d0d39e, 32'hc5595f20, 32'h43b00aa4},
  {32'h4541ad18, 32'h4395a9d8, 32'hc2f1ad8b},
  {32'hc4e3243c, 32'hc4932445, 32'hc4711b85},
  {32'h437fa170, 32'h440bff94, 32'h43d15d0b},
  {32'hc49f7f0d, 32'h42a48a81, 32'hc1c76770},
  {32'h44dfce61, 32'h43819005, 32'hc3663042},
  {32'hc468fbe4, 32'hc40890e4, 32'hc38fb87a},
  {32'h43ca850a, 32'h450510c1, 32'h42225a01},
  {32'hc49142b2, 32'hc41ca470, 32'hc1bfc569},
  {32'hc3a8d79c, 32'h417e057c, 32'hc54f2f17},
  {32'h44a77411, 32'h429ff7ce, 32'h428a8479},
  {32'h440dbce0, 32'h43515bb3, 32'hc4443082},
  {32'hc3bc17b5, 32'h436af5eb, 32'h4487daa7},
  {32'h4511a6d3, 32'h43db04ab, 32'hc4044533},
  {32'hc51aef57, 32'hc3a0f7cc, 32'h4465b769},
  {32'h44d5fa03, 32'h447d2316, 32'hc3b02a40},
  {32'h43af7f3c, 32'hc4a751f9, 32'h442168b4},
  {32'h44e2ba9c, 32'h43e70d92, 32'hc4786b28},
  {32'hc3f033e0, 32'h438fbf82, 32'h452fd5c9},
  {32'hc429988e, 32'hc2b079c9, 32'hc457d95a},
  {32'hc5428464, 32'h43afcea5, 32'h43f08632},
  {32'hc3430809, 32'hc2dfe52c, 32'hc584e409},
  {32'h44559c43, 32'h44664e94, 32'hc4ff9a05},
  {32'h4383ea0f, 32'h4572445f, 32'h4283da69},
  {32'h4407d5a9, 32'hc2928cf4, 32'h436e3193},
  {32'hc3f885f9, 32'h452c7547, 32'h43a976fb},
  {32'h444b6f75, 32'hc4c22714, 32'hc38fb6a6},
  {32'h44f0e8da, 32'hc3858307, 32'h42451635},
  {32'h451c63b0, 32'hc35224ff, 32'hc435ac09},
  {32'hc4e9cc41, 32'h44356b95, 32'h442b65c2},
  {32'hc3f1b4a6, 32'hc41cffe7, 32'hc35285a8},
  {32'hc43f6530, 32'h44c3070c, 32'hc39ae7f2},
  {32'h444221f8, 32'h43579c6f, 32'hc435a1ad},
  {32'h439bc4a9, 32'h443724f0, 32'hc419b354},
  {32'h4522d8b4, 32'hc42d9b7d, 32'h42c21471},
  {32'hc4d43757, 32'h44159647, 32'hc3c024ba},
  {32'hc2959e66, 32'h444827f0, 32'h44fa0104},
  {32'hc232c640, 32'hc37a4c0c, 32'hc5030088},
  {32'h44e94f0a, 32'h43b226e9, 32'h44193aba},
  {32'hc4da2ade, 32'hc2347f02, 32'hc3a59453},
  {32'h45675db0, 32'hc415f886, 32'h426f16d8},
  {32'hc4a3d076, 32'h43e5aef5, 32'hc37ce035},
  {32'hc45ce3a3, 32'hc46629ed, 32'h441617f1},
  {32'hc26d7884, 32'h4536ca3c, 32'h42f6c699},
  {32'h43a5ccd0, 32'hc342b2e4, 32'h44dfd1de},
  {32'h42a42de8, 32'h44368677, 32'hc3d2c0ae},
  {32'h4555591f, 32'h436f4956, 32'h43e50710},
  {32'hc450a694, 32'h43a60090, 32'hc422dcf2},
  {32'h448fe1bd, 32'h41980b6e, 32'h43c042cc},
  {32'hc4b0c540, 32'hc2eaca57, 32'hc4394772},
  {32'h416552dc, 32'hc2c05168, 32'h455759ac},
  {32'h437b9407, 32'hc4a20173, 32'hc3a38cf7},
  {32'hc488942a, 32'hc393e8ed, 32'hc2a449e8},
  {32'h4319f272, 32'hc54aabcc, 32'hc37c9375},
  {32'hc421d3ed, 32'h44462b22, 32'hc44fb7ff},
  {32'hc4714430, 32'hc35b8ce8, 32'hc2d127ee},
  {32'hc53a3016, 32'h4321edc9, 32'hbdcb1100},
  {32'h44a788de, 32'hc3e7aa36, 32'h442b7515},
  {32'h448155aa, 32'hc3b91113, 32'h44c351ee},
  {32'hc508eb5a, 32'hc43280d3, 32'hc4182014},
  {32'hc4255ffc, 32'hc2b4ad8e, 32'h4476d738},
  {32'hc3fadc29, 32'hc44ebab4, 32'h442da79b},
  {32'hc33b0a5d, 32'h44cf6248, 32'hc36a169e},
  {32'h4517a16e, 32'h4426afef, 32'hc28f750e},
  {32'hc49d21c8, 32'h4382156c, 32'h4210a1de},
  {32'h45304344, 32'hc2014ed4, 32'h438724c4},
  {32'h4412f5af, 32'h4555c702, 32'hc21d54a9},
  {32'h44a2a006, 32'hc413fa61, 32'h43291e77},
  {32'hc4bab7b5, 32'h43a498cb, 32'hc4181b05},
  {32'h450afe14, 32'hc2f3acbb, 32'h43cbd110},
  {32'hc458ed50, 32'h440db2de, 32'h4216e076},
  {32'h428f37b0, 32'hc42be174, 32'hc3aa6424},
  {32'hc48049d8, 32'h4447f7b6, 32'h426e99c5},
  {32'hc3fe0130, 32'hc31301c6, 32'hc268536a},
  {32'hc5181a51, 32'h4454506a, 32'h43891055},
  {32'h450ba003, 32'hc48fd469, 32'h43f64276},
  {32'h44f90f4b, 32'h4306f6ab, 32'hc16c4e27},
  {32'h4448d971, 32'hc3dd9ea1, 32'hc440fa20},
  {32'h43886478, 32'h44defdf9, 32'h4505da63},
  {32'hc3a78ff1, 32'hc48b2012, 32'h43ba9a29},
  {32'h44457c13, 32'h445af79f, 32'h43252c3a},
  {32'h44c1bd93, 32'h436ce30f, 32'h43bbcc0a},
  {32'h438ffa21, 32'h43fa54ce, 32'hc457b1b4},
  {32'h43ef870d, 32'hc420ea05, 32'h446568a6},
  {32'h453e48e9, 32'hc3e1698a, 32'hc3129682},
  {32'h44ac0bcc, 32'hc40e719b, 32'h43616c7d},
  {32'hc385f263, 32'hc496054b, 32'h44d86da7},
  {32'h42f51039, 32'h4498b4cb, 32'hc4acd1d4},
  {32'h449fde76, 32'h446d1c86, 32'hc42488ab},
  {32'hc3d48bba, 32'hc45a3f8c, 32'h448b872f},
  {32'hc45968ab, 32'h444eb085, 32'h43e8d0f0},
  {32'hc4c58cee, 32'hc43c4841, 32'h43b0d425},
  {32'h439ec601, 32'h451b33b3, 32'h42280f37},
  {32'hc38353fb, 32'hc4c99768, 32'h42a4ca00},
  {32'h44dbdc8a, 32'hc3c72ea8, 32'hc3e47514},
  {32'hc57abb1d, 32'hc3a93977, 32'hc3fbb120},
  {32'h44ded9d7, 32'h4330f032, 32'hc30da0da},
  {32'hc3da74ec, 32'hc4338b68, 32'h41bf4704},
  {32'h43abc26f, 32'h44adeab3, 32'h4334b7c5},
  {32'h44ddd3f0, 32'hc2e30347, 32'hc2b0d1c8},
  {32'h4538a134, 32'h443ea910, 32'h439d8301},
  {32'hc569653b, 32'hc3682b2e, 32'h430905c0},
  {32'h4383afbd, 32'h44090a2f, 32'hc409ff91},
  {32'h43ab1436, 32'hc462161a, 32'h42e7b348},
  {32'hc42d7468, 32'h440961b6, 32'hc4615a88},
  {32'h43cdbea8, 32'hc45ca044, 32'h44a6514c},
  {32'hc319daa0, 32'hc33ecb34, 32'hc47f68b2},
  {32'h44fbe234, 32'h44061605, 32'h44204241},
  {32'hc3f9a87b, 32'h4394fb28, 32'hc4300d63},
  {32'h41d1f960, 32'hc31b491c, 32'h447856dc},
  {32'hc49d93f1, 32'h436d2bfa, 32'h430fc3a4},
  {32'h4501f8dd, 32'h42e0a770, 32'h4408cba6},
  {32'h44617fe4, 32'h4466a6c8, 32'hc35612c2},
  {32'h448fc2a0, 32'h44103336, 32'h43aee156},
  {32'hc3c9ab2c, 32'hc40de155, 32'hc4718328},
  {32'hc443e1fe, 32'h4405c839, 32'h41a0cb34},
  {32'hc2b79770, 32'hc4881299, 32'hc45fa3a4},
  {32'h43093937, 32'h4439349a, 32'hc340f946},
  {32'hc526c0fe, 32'hc358460d, 32'h43c27e58},
  {32'h4450786e, 32'h43f2a0e1, 32'h45186242},
  {32'hc3a7d2e2, 32'hc4a4abfa, 32'hc497d65f},
  {32'h4419b591, 32'h44446184, 32'hc18df822},
  {32'hc3ec9857, 32'hc576d59c, 32'hc29c908b},
  {32'h444dda9e, 32'h44bd4cc9, 32'h4466e450},
  {32'hc3a8e4c2, 32'hc34bf32d, 32'h428d4dfe},
  {32'h44b40372, 32'h438e37e5, 32'h43c2845c},
  {32'h4326ee27, 32'hc5777143, 32'hc38ecaa7},
  {32'h44a3543a, 32'h4299d135, 32'h43d84256},
  {32'hc568c89d, 32'h43e88f60, 32'hc3d3eafa},
  {32'h451f8973, 32'h4373dfc9, 32'hc32ca4c8},
  {32'h43cd1512, 32'hc5064caf, 32'h43846f04},
  {32'h42e8d7a3, 32'hc42aa83e, 32'h44b8cb2c},
  {32'hc40bdabc, 32'h44315ea6, 32'hc3efed36},
  {32'hc54eb708, 32'h437c6855, 32'h43436d59},
  {32'hc42954b7, 32'h423c68dd, 32'hc56ae6ef},
  {32'h440e252d, 32'h44ddede9, 32'h41e8a6f8},
  {32'h43bf1c4a, 32'hc41d8b67, 32'hc4f09ecd},
  {32'hc46926fe, 32'h43d517df, 32'h44c51194},
  {32'h44117706, 32'hc4969adb, 32'hc39e3fe9},
  {32'h436cb975, 32'hc3fdbaf9, 32'h44d21a97},
  {32'h43e4a17e, 32'h439221d7, 32'hc4908199},
  {32'h43dfd979, 32'h4368c314, 32'h43ff4b07},
  {32'hc1fa1df0, 32'hc4c83708, 32'hc44dca15},
  {32'h43136b0a, 32'h449c6bb3, 32'h447ef14c},
  {32'hc33da9dc, 32'hc3be9676, 32'hc369d357},
  {32'hc50ccc12, 32'h438b3be4, 32'h440bff38},
  {32'h43496720, 32'h4315d400, 32'hc43b1d63},
  {32'h44356de1, 32'h436aa40f, 32'h4406f630},
  {32'h4498a234, 32'hc4a27df2, 32'hc3f4381b},
  {32'hc48112bc, 32'h44843cce, 32'h43f9ae04},
  {32'h4438fd8b, 32'h41f33690, 32'h433f5f51},
  {32'hc49bb7dc, 32'h447d50e2, 32'h44667692},
  {32'h44efe15a, 32'h43658300, 32'hc3970e28},
  {32'hc3ef71f6, 32'h441b7f34, 32'h43d65043},
  {32'h449b9f88, 32'h43c3de4a, 32'h42b545ce},
  {32'hc57b8cee, 32'hc2a9c79a, 32'hc29c8dc3},
  {32'hc4b86506, 32'hc3556b81, 32'hc3142756},
  {32'hc316ff04, 32'h4274b710, 32'h43b59d9f},
  {32'hc57af3a4, 32'hc3526132, 32'h440617a5},
  {32'h44225788, 32'h43878550, 32'h44de63e6},
  {32'h44a779d6, 32'hc031fb32, 32'h43a03ca8},
  {32'h44ab3e8b, 32'hc449c15e, 32'h43230751},
  {32'hc4005286, 32'h45310c5e, 32'h411f1a39},
  {32'h4513d987, 32'h43a28d73, 32'hc3d27475},
  {32'hc4da1ca4, 32'h44be816d, 32'hc1a77210},
  {32'h44290c74, 32'hc51a25da, 32'hc3acc599},
  {32'hc475c87f, 32'h4366e1b4, 32'hc47f40de},
  {32'h4449c36f, 32'hc3766b18, 32'h44ef7247},
  {32'hc3f0ff52, 32'h4371fae1, 32'hc512ef31},
  {32'hc40631de, 32'hc35636da, 32'hc35a32f4},
  {32'hc52846d4, 32'hc2e9b0fd, 32'hc28c474b},
  {32'h4422d9fe, 32'hc4f37210, 32'hc3422162},
  {32'h44804d6d, 32'h43e04651, 32'hc159ee56},
  {32'h44764409, 32'hc4915133, 32'hc44de28d},
  {32'hc3b82987, 32'h4388745b, 32'h44a9e0cc},
  {32'hc458b35e, 32'hc3e15d70, 32'hc26ececb},
  {32'hc3644220, 32'h4361ee07, 32'h4426707c},
  {32'hc3eeb698, 32'h447ab3ab, 32'hc4b8d561},
  {32'h4398ddf1, 32'h44e2121e, 32'h43840229},
  {32'hc38f1800, 32'hc47db3ac, 32'hc4dd2cae},
  {32'h42bf4f75, 32'h442edafb, 32'h43b35241},
  {32'h43f680b0, 32'hc47a7a3c, 32'hc2d725c8},
  {32'h434ba484, 32'h453409bb, 32'h4346e86d},
  {32'h4509dde1, 32'hc3b85651, 32'hc49cde66},
  {32'h447af3d0, 32'hc1ccd964, 32'hc49c130c},
  {32'hc559153e, 32'h4326e2ac, 32'hc315f5a5},
  {32'hc2b6bb5d, 32'h437f5432, 32'h4405f465},
  {32'hc42a26f4, 32'hc44602d0, 32'hc3af69f8},
  {32'h450eb44e, 32'h43867046, 32'hc1e80efe},
  {32'hc326d982, 32'h42e891e9, 32'hc40914ba},
  {32'h446842ce, 32'h452828af, 32'hc3202255},
  {32'hc4b5ce7e, 32'hc4afd419, 32'h415d339a},
  {32'hc48223d5, 32'hc310f27a, 32'h4407212a},
  {32'hc33d0060, 32'hc3844e4e, 32'h44b1c69a},
  {32'hc3505380, 32'h43228716, 32'h43b9d3c4},
  {32'h446bb668, 32'h4271a7e2, 32'h44186947},
  {32'h438c76e4, 32'h42f300f5, 32'h45465263},
  {32'hc342dc50, 32'hc35a8b36, 32'hc4130492},
  {32'hc4dd04a7, 32'h437d1bf1, 32'h43a5264d},
  {32'hc370d4bc, 32'h4267ce9c, 32'hc564203c},
  {32'h44102067, 32'h444ac880, 32'hc3495422},
  {32'hc213faf0, 32'hc440039b, 32'hc3f0f540},
  {32'h4508a4b6, 32'hc25ba95a, 32'h445960b4},
  {32'hc504c8f9, 32'hc4538695, 32'hc43ad40e},
  {32'h453b0fe2, 32'h43116b37, 32'hc41f21aa},
  {32'hc4ca840e, 32'hc4827a1b, 32'hc4762fe8},
  {32'h4392e76c, 32'h44f8872b, 32'h433a757c},
  {32'hc4f8fca2, 32'hc381769f, 32'hc316fd10},
  {32'h4415c174, 32'h44e2faf3, 32'h43fbc038},
  {32'hc4b620d0, 32'hc43e1a1f, 32'hc4cc518f},
  {32'h4320eee7, 32'h43c75949, 32'hc3c3085e},
  {32'h43116bf0, 32'h44caec13, 32'hc10edd48},
  {32'hc424df25, 32'hc4b4f04f, 32'h43a6121f},
  {32'h435c42d9, 32'h4520c45b, 32'h4474d023},
  {32'h430800fc, 32'hc3bf095e, 32'hc2a38b25},
  {32'h43b21f2e, 32'h44fcfb1f, 32'hc3bd2592},
  {32'hc33ee31a, 32'hc57ab9eb, 32'hc2ce42bf},
  {32'h43ac90a8, 32'h43303508, 32'hc4171c1a},
  {32'hc53307ed, 32'hc3b87f76, 32'h42db68b8},
  {32'h44bc087b, 32'hc40aee6f, 32'hc39c4194},
  {32'hc375587d, 32'hc2729607, 32'h44866fc7},
  {32'h43e5afca, 32'h44c1342f, 32'hc3e037f8},
  {32'hc2eb6978, 32'hc516f792, 32'hc1b3d7fe},
  {32'hc4d0657e, 32'h43a83e7c, 32'hc2ede8da},
  {32'hc3d32e86, 32'hc40454f9, 32'hc284ccd2},
  {32'h434aa7d8, 32'h43b7ad4b, 32'hc51ea94b},
  {32'h4482f04e, 32'hc2807d16, 32'h43d01986},
  {32'h445551c0, 32'h43ddf579, 32'hc4832150},
  {32'hc42b2676, 32'h42869697, 32'h450ae29f},
  {32'hc36de38a, 32'h44cf6cfc, 32'h42f8389a},
  {32'hc40d23b8, 32'hc4e8f03a, 32'h443614a6},
  {32'h44ffe4bd, 32'h44505d0e, 32'hc4aed56e},
  {32'hc4332e63, 32'hc213748b, 32'h4315766d},
  {32'h44af942d, 32'h4491706d, 32'hc2a3fc73},
  {32'hc35bc718, 32'hc3b18044, 32'h449d67a5},
  {32'h42f9d189, 32'hc3b434cd, 32'hc5143a0e},
  {32'h42b32a20, 32'h426c2848, 32'h4500e948},
  {32'h445644e6, 32'hc3c22edd, 32'hc4efac5f},
  {32'h4519bac1, 32'hc4480b07, 32'hc4630d22},
  {32'hc310cef0, 32'h45312a10, 32'h436d9f98},
  {32'h450ba001, 32'hc19ca21b, 32'h42dca5de},
  {32'h4169ad9c, 32'h4583cca4, 32'h42c5da2e},
  {32'h4423e6b2, 32'hc4b143fa, 32'h425ae31a},
  {32'h44a32194, 32'h42b4bbfb, 32'hc2d76a7d},
  {32'h430f9d10, 32'h43475ed4, 32'h43659f38},
  {32'hc453d57a, 32'h433b56b2, 32'h437197cb},
  {32'h44622953, 32'hc39247da, 32'h441459e3},
  {32'hc47bdebc, 32'h448cf0e0, 32'h431800b0},
  {32'hc3cc7bb1, 32'hc52e90c8, 32'h43b2d67f},
  {32'hc2a3543f, 32'h43ca77f8, 32'hc40ee03a},
  {32'h4460f5e6, 32'hc342ab9c, 32'h44c762c5},
  {32'h42cc6e50, 32'h4536e19a, 32'hc3cd715f},
  {32'h44fdc7c2, 32'h422e18e5, 32'h43c974c4},
  {32'hc4a97788, 32'hc2cf2df2, 32'hc4f0760a},
  {32'h4425c64d, 32'h43bf9fc4, 32'h44e68a99},
  {32'h450ebdbc, 32'hc2858a6a, 32'hc3b0c65d},
  {32'h440606df, 32'hc48394ce, 32'h444a0f01},
  {32'hc4f33e15, 32'hc20a5510, 32'h43ff1b64},
  {32'hbe92df80, 32'hc4cf2440, 32'hc3b43c5a},
  {32'hc4e836e0, 32'h4484f02c, 32'h43a897b6},
  {32'h43c6f8fe, 32'hc3880e5b, 32'h44f8f2bc},
  {32'hc357d3e4, 32'h4444c7c4, 32'hc3bca206},
  {32'h444b8f45, 32'h431be162, 32'h44bd3658},
  {32'hc3ee9744, 32'hc2b6c8a2, 32'hc50565e4},
  {32'h444d9531, 32'h4255e71e, 32'h44641ade},
  {32'hc42a16f5, 32'hc3d2cd7b, 32'hc4973434},
  {32'h436cd4a4, 32'hc4b0d7b8, 32'h451e4e0c},
  {32'hc5039a88, 32'h43361c1f, 32'h4341f8ed},
  {32'hc4c93f9e, 32'h43429719, 32'hc3f69b0b},
  {32'hc31749d0, 32'hc5381518, 32'hc22fac73},
  {32'hc41208b1, 32'h44860b1a, 32'hc39af731},
  {32'hc2b17152, 32'hc42ddd48, 32'h434d7694},
  {32'h4381af10, 32'h453cf69c, 32'h4369eb48},
  {32'hc45f3ff4, 32'hc4fc42b3, 32'h42b577d5},
  {32'h44acf950, 32'h44276df8, 32'h448aeea7},
  {32'hc4a9662b, 32'hc481fa73, 32'hc40b452c},
  {32'h444e6904, 32'hc46f75f0, 32'h445f5c08},
  {32'h433df4ad, 32'h43107f96, 32'h45096756},
  {32'hc47b5d6a, 32'h4400c410, 32'hc2af38ed},
  {32'h44ad2385, 32'hc332a39a, 32'h4393c97e},
  {32'hc4a16b6e, 32'h4308da7f, 32'hc30562fb},
  {32'h44250b03, 32'hc4bfdb17, 32'h43c82042},
  {32'h43e3eabb, 32'h45303602, 32'h41795fa9},
  {32'h446e90e8, 32'hc446fef6, 32'h434cc414},
  {32'hc4474b24, 32'h440eed86, 32'h439ef0ce},
  {32'h45257797, 32'h432ce61e, 32'hc40eae54},
  {32'hc50746e2, 32'hc2eb8eba, 32'hc2a2cbb0},
  {32'h44a4ecb2, 32'hc3f3b8aa, 32'h426d97e1},
  {32'hc4db8f2b, 32'h43acfe40, 32'h43b2acd8},
  {32'h43b7816a, 32'hc50892bc, 32'hc3aa446d},
  {32'hc480d03e, 32'h452518e0, 32'h43db81ed},
  {32'hc172ec3c, 32'hc56254d0, 32'hc40e1706},
  {32'h443b3244, 32'hc40c3a30, 32'h43ef2e70},
  {32'hc3cebd6f, 32'hc3be05a4, 32'hc54a23e3},
  {32'hc425fbfc, 32'hc307f7cb, 32'h4444d616},
  {32'hc40a71c6, 32'hc3b65e0c, 32'h444289cb},
  {32'h43895680, 32'h43f7256b, 32'hc4d66a6d},
  {32'hc50b9d36, 32'hc3445663, 32'h41ae9b4a},
  {32'h443ee741, 32'h43e047b8, 32'hc48c9b56},
  {32'hc480f4ae, 32'h431be4ac, 32'h45053892},
  {32'h440f3bb9, 32'hc3b503da, 32'hc41af2ef},
  {32'hc473f7a6, 32'h44398e7d, 32'hc1c1ea3a},
  {32'hc5198b79, 32'h43d325b6, 32'h43c243bd},
  {32'hc4914aca, 32'hc1d37e90, 32'hc41a75a0},
  {32'h44a6ef36, 32'hc2b47c0f, 32'hc376b2ca},
  {32'hc3f827db, 32'h4272b5fd, 32'h44c69f18},
  {32'h447b6db8, 32'h44440376, 32'hc404da77},
  {32'hc444383a, 32'hc48b534f, 32'h442dc1c0},
  {32'hc37d647c, 32'h44d6bb29, 32'hc47452e3},
  {32'h43d5230f, 32'hc23f8522, 32'h44b4f02c},
  {32'h43895270, 32'hc45599bc, 32'hc413d375},
  {32'hc526f41a, 32'h42e22379, 32'h42b0a368},
  {32'h43e5002a, 32'h43b6210c, 32'hc3824043},
  {32'hc51ce0d9, 32'hc3ef315e, 32'h437b6ee8},
  {32'h4569d8d4, 32'h43c10e55, 32'hc39230c3},
  {32'hc260808a, 32'hc3b5cd7c, 32'hc2aafa1c},
  {32'h4501f9ad, 32'h439094d6, 32'h4327cb4b},
  {32'hc38905f5, 32'hc52165f7, 32'h42dac4b3},
  {32'hc49c04f0, 32'h44172687, 32'hc39ac94d},
  {32'h43590372, 32'h442b48c4, 32'hc2956ac7},
  {32'h432e16eb, 32'hc2f0aef1, 32'hc48ab308},
  {32'h4370eac0, 32'hc4e58459, 32'h44b090a5},
  {32'hc51fccd0, 32'h43f9d486, 32'h41a34a03},
  {32'h44b3d67f, 32'hc1e20967, 32'h43e51959},
  {32'h433d8f4a, 32'hc4b5e7ea, 32'hc3ca3c1b},
  {32'hc4833d88, 32'hc14eadf4, 32'h4347d1c8},
  {32'hc3fb4160, 32'hc471b574, 32'hc4f5f3eb},
  {32'h44fac3fa, 32'h4381ad50, 32'h43bbfe7c},
  {32'h442b6218, 32'hc36f706a, 32'hc40c761c},
  {32'h44993b56, 32'h42cc0ba2, 32'h434f914f},
  {32'hc427b3ab, 32'h44cf82e2, 32'hc4b2fbf7},
  {32'h45046bf6, 32'h43e709a6, 32'h412fb828},
  {32'h42b15a18, 32'hc5425e36, 32'hc408af59},
  {32'h417d50a3, 32'h435abece, 32'h4552eedf},
  {32'h433fd482, 32'hc4a70bcc, 32'h4307eeee},
  {32'h449576ba, 32'h44396fb8, 32'h449b1072},
  {32'h43abff60, 32'hc48ebf92, 32'hc4f0b528},
  {32'h44840f7c, 32'h44396bc3, 32'hc2de558a},
  {32'hc4b80b16, 32'hc412be5c, 32'hc38b7e6a},
  {32'hc2b5e0ee, 32'h45073cd4, 32'h4454af10},
  {32'hc48c6e63, 32'hc36cff92, 32'hc3db8733},
  {32'h4499e463, 32'h431bb52f, 32'hc3997285},
  {32'hc3910080, 32'hc3cae75d, 32'hc2ddf0c4},
  {32'h455159ce, 32'h43cef4d5, 32'h44477d2e},
  {32'hc51ede12, 32'hc2957355, 32'hc46783fb},
  {32'h44af99a4, 32'h439e2055, 32'hc2c81afc},
  {32'hc1b56e30, 32'h4490fe0d, 32'hc458e099},
  {32'h429c64e0, 32'h42bc1426, 32'h44a2f636},
  {32'h43064978, 32'h4374ffee, 32'hc482ff81},
  {32'hc474554d, 32'h43b17a3a, 32'h43dfbcd2},
  {32'hc2416662, 32'hc3f0f599, 32'hc4dc9b6d},
  {32'h4492d900, 32'h43a0a8bf, 32'hc3c38cde},
  {32'h43eb8068, 32'hc4a89295, 32'hc4cd8271},
  {32'hc54d27d8, 32'h440dc850, 32'h4333a80e},
  {32'h447b3554, 32'hc44dfbac, 32'h42f6ed49},
  {32'hc30f00c8, 32'h4437db8f, 32'h4426b706},
  {32'h43dea37c, 32'h43df7945, 32'hc46d718a},
  {32'h438975f0, 32'h43bab6b4, 32'h43c62d3f},
  {32'h42008d00, 32'hc2a90f5b, 32'hc204c5a8},
  {32'hc4ba7ce2, 32'h43cbe705, 32'h436b12be},
  {32'h440bf3af, 32'hc3a8fcd1, 32'hc3c93752},
  {32'hc4e62d91, 32'h43c2ecea, 32'h440af258},
  {32'h440e7955, 32'hc4149abd, 32'hc300c8a4},
  {32'hc4a6cb71, 32'hc19a6c84, 32'h4004b767},
  {32'hc368c670, 32'hc4e93d7f, 32'hc33511e8},
  {32'hc3d3caa4, 32'h44b5cb84, 32'hc23a0baf},
  {32'h4538483a, 32'h413517f0, 32'hc3c9b10c},
  {32'hc53def59, 32'h43d7459d, 32'hc31284be},
  {32'h4540df39, 32'h428b8a79, 32'h43013d92},
  {32'hc3a2014a, 32'h41edc266, 32'h4299ad4a},
  {32'h44db9cf5, 32'hc3ba4e0a, 32'hc292f595},
  {32'hc49d1e04, 32'hc3f40f86, 32'h43b66836},
  {32'h450f9724, 32'h41b91ab7, 32'hc3955317},
  {32'hc218ede7, 32'hc0724120, 32'h44b2a185},
  {32'hc47cd516, 32'hc324e2fd, 32'hc51041d3},
  {32'h441aeb78, 32'hc38c12eb, 32'h427b5fe2},
  {32'h442bb8d2, 32'h4451694d, 32'h4399b516},
  {32'h43f792ac, 32'hc51add86, 32'hc381850d},
  {32'h4307b881, 32'h45236334, 32'hc2878fe5},
  {32'h4347e8b9, 32'hc4045c65, 32'h43b2b5e7},
  {32'hc4e9fdd4, 32'h447a686c, 32'h439513a0},
  {32'h44d9c4ae, 32'hc4901e38, 32'hc368731c},
  {32'hc4a5758e, 32'h415913e8, 32'hc3dbdd59},
  {32'h45069a38, 32'h4323642a, 32'h431d17ba},
  {32'hc34a1fd0, 32'h422f0194, 32'hc4a2ac11},
  {32'h43d1dd11, 32'hc3dd8680, 32'hc3d89cc8},
  {32'hc2de955d, 32'h44ab5b0a, 32'h4409f924},
  {32'h43f2e058, 32'hc49296d5, 32'hc3ae95c2},
  {32'hc2cb20b2, 32'h450f4a9e, 32'hc2479da9},
  {32'h426097f8, 32'h42ccfff0, 32'hc4d737ff},
  {32'hc246dc4c, 32'h450e9450, 32'hc3c69d14},
  {32'h4487a7b3, 32'hc340f093, 32'hc3a646a0},
  {32'hc42006ac, 32'hc3d18af5, 32'h44018acc},
  {32'hc1f7aee0, 32'hc441ccb8, 32'hc48c0102},
  {32'hc476d72a, 32'hc3ca4b82, 32'h4228e748},
  {32'h4395cb5f, 32'hc40a3190, 32'hc3bc0428},
  {32'hc4385d11, 32'hc0c4baee, 32'h44fb9a04},
  {32'h42f777a0, 32'h4381f16f, 32'hc3c3d42c},
  {32'hc50917c9, 32'h44b006e3, 32'h43b4e407},
  {32'h4363ec80, 32'hc424ce56, 32'hc50c88b2},
  {32'h442c7811, 32'h42855b1e, 32'hc4a919ff},
  {32'hc4c3dc1a, 32'hc352aaab, 32'h44bcb189},
  {32'h4508f85a, 32'h438b934b, 32'h4386650d},
  {32'hc5374b00, 32'hc4503403, 32'hc3aed2fb},
  {32'h44bac850, 32'h4462cdb2, 32'h43f9ad32},
  {32'hc41771ee, 32'hc32407fd, 32'hc3c28f00},
  {32'hc341ab00, 32'h44cc63a5, 32'h43884bb5},
  {32'hc565b465, 32'hc2f25646, 32'hc3d2b4f6},
  {32'h45140433, 32'hc3cd83f8, 32'h43280f2e},
  {32'hc519d127, 32'h4353057e, 32'h4346a4f0},
  {32'h44d6c1ff, 32'h43eb369c, 32'h4437ca1f},
  {32'hc404e668, 32'h43667566, 32'h442ced53},
  {32'h444a9773, 32'hc2bc5da1, 32'h44863e01},
  {32'hc3f49002, 32'hc55aa36a, 32'hc35b053d},
  {32'h45165332, 32'h430b238c, 32'h41a8c33b},
  {32'hc39ddd10, 32'hc423e16c, 32'hc44850a4},
  {32'h436e93b3, 32'h43391ab2, 32'h453189d0},
  {32'hc536808c, 32'hc3f6053d, 32'hc2e2fd84},
  {32'h41a97d10, 32'hc420b1ab, 32'h44381fa2},
  {32'hc5392bec, 32'hc3be8aae, 32'hc3a6c6b0},
  {32'h42aa2a30, 32'hc3cb268a, 32'hc37a866c},
  {32'hc39757c6, 32'hc4ba65ca, 32'hc4ae71c5},
  {32'h42d13c35, 32'hc0232194, 32'h44e4aea6},
  {32'hc477e56c, 32'h435b66c2, 32'hc452fce1},
  {32'hc35e75f1, 32'h453216b4, 32'h432f1fe4},
  {32'hc2a6a88c, 32'hc43516f8, 32'hc51b2e48},
  {32'h45031a6e, 32'hc3b98b0e, 32'h4370c003},
  {32'hc3293dcc, 32'h4488fc7a, 32'hc416aa9d},
  {32'hc2c1c3c8, 32'hc5396a43, 32'h4305252f},
  {32'h45158a8f, 32'h444ab8dc, 32'hc2e6388d},
  {32'h44dd5177, 32'hc2b9c1ca, 32'hc1d2d3d8},
  {32'hc2e62410, 32'h455a93ff, 32'hc2bf19c4},
  {32'hc4c59859, 32'hc4869c8a, 32'hc2bb0e3a},
  {32'h44215174, 32'h44085cc7, 32'hc185d8fa},
  {32'hc5683d96, 32'hc402bb5d, 32'h438dbf2f},
  {32'h44cedfb4, 32'h440589b0, 32'h43c8ab57},
  {32'hc4c44a7d, 32'hc3e330a1, 32'h43ac5c76},
  {32'h4521b40e, 32'h439e3125, 32'h436c454a},
  {32'hc4824c28, 32'hc3ac4aaa, 32'hc3590286},
  {32'h44447dd6, 32'h43b686b2, 32'h4392bfee},
  {32'hc4365841, 32'hc4082378, 32'h4405f3b9},
  {32'h44ae96bd, 32'h43e2fd6b, 32'hc2daa892},
  {32'hc4fd5b5d, 32'hc2ba22af, 32'hc3c82455},
  {32'h445b520c, 32'h437c4f15, 32'hc3c17423},
  {32'hc49ae187, 32'hc46befdf, 32'hc3d48075},
  {32'h440bf2b6, 32'h43f7c0df, 32'hc391cc44},
  {32'hc4926389, 32'hc4a5674a, 32'h44f94439},
  {32'h43819c08, 32'h4489082d, 32'hc48509c0},
  {32'hc3857d71, 32'hc40b75db, 32'h44967233},
  {32'h401754c8, 32'hc1fd00fe, 32'hc51eeb07},
  {32'hc4257cea, 32'hc310d284, 32'h448b7aa8},
  {32'h449fe093, 32'h436cdb70, 32'hc4768ceb},
  {32'hc487681c, 32'h42a0c932, 32'h44073d4b},
  {32'h4553bf3c, 32'hc4335949, 32'hc43e1972},
  {32'h43871692, 32'hc55b1d69, 32'hc20d2ab4},
  {32'hc4a5d970, 32'h43f776e6, 32'h426c072a},
  {32'hc4638e84, 32'hc265ecf2, 32'h43eb14d3},
  {32'h4108ae00, 32'h4569c732, 32'h434eadb8},
  {32'h451eba3a, 32'h42627b69, 32'h43d51340},
  {32'h42bdb2bc, 32'h445df529, 32'hc2599752},
  {32'h44a732bc, 32'hc3e6de52, 32'hc455afcc},
  {32'hc4201602, 32'h446045ea, 32'h4460a1d4},
  {32'h45377db3, 32'hc2a405de, 32'h439b2d27},
  {32'hc52044ce, 32'hc30874e4, 32'hc3e32b84},
  {32'h43a6504c, 32'hc3bd1ebf, 32'h4293b783},
  {32'hc504229a, 32'hc2edb944, 32'hc42155ff},
  {32'hc239a8d3, 32'hc4dee8f1, 32'h442e7eaf},
  {32'hc37de3c9, 32'h43a07842, 32'hc52adee0},
  {32'h43a179b6, 32'hc3ad26a2, 32'h43a26659},
  {32'hc51b15d4, 32'h435c5b96, 32'hc46bbd6c},
  {32'h452e1bc0, 32'h4402d351, 32'h4183c151},
  {32'h4284d6c4, 32'h431101e2, 32'hc4bc07b6},
  {32'h450abff2, 32'hc43f7214, 32'h439c3a01},
  {32'hc4850e61, 32'h4531a627, 32'hc2944c4e},
  {32'h44bbe548, 32'hc2bd073c, 32'hc38bb7d6},
  {32'hc40596b2, 32'hc155fa93, 32'hc4d0d37e},
  {32'h44c88c57, 32'hc231ed3e, 32'h43a13922},
  {32'h440e31ad, 32'h441d28fa, 32'hc4f8ff8a},
  {32'h44d1c2af, 32'h429ec0d0, 32'h43c3f5bc},
  {32'hc4b7cc9c, 32'hc42b55a4, 32'h43327d7d},
  {32'hc4c0f789, 32'h43312330, 32'hc3f3d6dd},
  {32'hc28673b8, 32'hc3ec49f7, 32'hc4d47ee1},
  {32'hc2820100, 32'h43a53c76, 32'h44278435},
  {32'hc476123b, 32'h445aa34d, 32'h40a2add0},
  {32'hc5399822, 32'hc188fd91, 32'h432f9a4c},
  {32'h448aa1ef, 32'hc49ec36f, 32'h43b14037},
  {32'hc524be03, 32'h43253bae, 32'hc3d05918},
  {32'h43745163, 32'hc47d726e, 32'h4242b22d},
  {32'hc53a61b0, 32'h42e8e46a, 32'hc210da27},
  {32'h4279ef00, 32'hc4ca5b4a, 32'h44a5e280},
  {32'h45370360, 32'hc2a762bf, 32'h4478391a},
  {32'h4443987e, 32'hc2b68226, 32'hc4826a8d},
  {32'hc46d23aa, 32'h4243f241, 32'h43eedc3a},
  {32'h43d6e926, 32'hc4cb678b, 32'h4380660c},
  {32'hc430f8c7, 32'h41bfde6a, 32'hc49c4793},
  {32'h4486c7cd, 32'hc40d01b1, 32'h444ca960},
  {32'h44a9b5f9, 32'h44135ec8, 32'h40c63914},
  {32'h442adffe, 32'hc4bec94f, 32'h4464ec11},
  {32'hc4f8966a, 32'h43195354, 32'h4201856d},
  {32'h450c2e9c, 32'hc3bd1395, 32'hc198194b},
  {32'hc59249e2, 32'hc30d1db8, 32'hc1feb80b},
  {32'h452fc01a, 32'hc3ced419, 32'hc2a8f8f8},
  {32'h4431948f, 32'hc3449fa2, 32'h43393422},
  {32'h451ecc8b, 32'hc3f38668, 32'h4231ae69},
  {32'h434ccaa0, 32'h44dd79ca, 32'hc41c8687},
  {32'hc4b35987, 32'hc3e52e58, 32'h40ac7454},
  {32'hc532323c, 32'h4421fe91, 32'hc304d4ce},
  {32'h45002388, 32'hc47961bd, 32'h439fca59},
  {32'h43b3f11c, 32'hc49abe7d, 32'h43e2e455},
  {32'hc424a47c, 32'h44fc2666, 32'hc4b3c201},
  {32'h42131380, 32'hc506e2b8, 32'h44af3011},
  {32'hc3dafe9a, 32'hc2809d99, 32'h43c9b511},
  {32'h4380adf0, 32'h43317c4f, 32'hc4b0c99c},
  {32'hc3ffa70d, 32'h43c15769, 32'h43f14ed5},
  {32'h4449add9, 32'h444b702e, 32'hc4a6d4e1},
  {32'hc474ad93, 32'hc349cedc, 32'h436bc28e},
  {32'hc4436155, 32'hc220680a, 32'hc476afd2},
  {32'h44f38376, 32'h42090188, 32'h4416c0f1},
  {32'hc3364fcc, 32'h4483ec92, 32'h44d82411},
  {32'h4416a927, 32'h43ff51f2, 32'hc499a5ef},
  {32'h4442a188, 32'h450785ac, 32'hc3c46ce5},
  {32'hc4f4a5ce, 32'hc40d0b2f, 32'h4395e531},
  {32'hc50d7667, 32'h42d19ba0, 32'hc324f864},
  {32'hc505b241, 32'hc40c7ca0, 32'h4472398b},
  {32'h44a3dd9a, 32'h4392f08a, 32'hc318759f},
  {32'hc4661bee, 32'hc20855d5, 32'h43a9973e},
  {32'h4515cfe2, 32'h439b5c63, 32'hc3b83597},
  {32'hc5789935, 32'hc303b55a, 32'h428fa6b7},
  {32'hc4dd2486, 32'hc35acfb6, 32'hc23cce3c},
  {32'h43063518, 32'hc567f8b3, 32'hc39efe61},
  {32'h44df065f, 32'h446c7eb7, 32'h43278c24},
  {32'h45088b91, 32'hc373e58e, 32'hc3790a06},
  {32'h44a654ec, 32'h444a0380, 32'h42a07e5a},
  {32'hc39476c4, 32'hc5222cb6, 32'h43906534},
  {32'h44cfb02c, 32'hc3d0a8be, 32'hc3fe8037},
  {32'h43c8aacc, 32'hc3124869, 32'hc3163d5c},
  {32'hc2a321c0, 32'h44af557c, 32'hc492f437},
  {32'hc384a2ec, 32'hc508fbdb, 32'h44bc8769},
  {32'hc3f060d7, 32'hc17479a4, 32'hc465f67b},
  {32'h41c2bc84, 32'h450a9b3c, 32'h4228cad2},
  {32'hc531e222, 32'hc38a701a, 32'hc3320c1f},
  {32'h43e37d8b, 32'h428ddbe1, 32'h4409e9ab},
  {32'hc3e64fbe, 32'hc4eb46f8, 32'hc4e0b139},
  {32'h44f3f44c, 32'h4414d7e4, 32'h443b3ccb},
  {32'hc371c351, 32'hc44840ac, 32'h43dbdd7c},
  {32'hc381af8a, 32'h44c30cab, 32'h43bfceea},
  {32'hc39c1d42, 32'h44a2d380, 32'hc4c341f9},
  {32'h4313a0e9, 32'h44a2f992, 32'hc1a3524c},
  {32'hc51bd9fa, 32'hc33dfd34, 32'hc37bea3b},
  {32'h44c154b0, 32'h43ac471b, 32'h440618bf},
  {32'hc4ac2634, 32'hc41067d9, 32'hc2390a78},
  {32'h4350530c, 32'h450c4085, 32'h44dbcf38},
  {32'hc43b249c, 32'hc4795b05, 32'hc5056084},
  {32'h44387a63, 32'h4293b7b3, 32'h43ebb6d2},
  {32'h430148cc, 32'hc5813463, 32'hc1c7eac3},
  {32'h44e35bdc, 32'h446587c5, 32'h443fd1c3},
  {32'h44d2c32f, 32'hc2f752c7, 32'hc34dfd5b},
  {32'hc33d314a, 32'h4517bbb8, 32'h43797273},
  {32'h423cc940, 32'hc583016a, 32'hc36acc08},
  {32'h428a883e, 32'h4325b656, 32'h43d5b538},
  {32'hc51201cd, 32'h430f677a, 32'hc30607a5},
  {32'h449e2edd, 32'hc4257bd5, 32'h4431f3c0},
  {32'h42f816c1, 32'hc496cb27, 32'hc3fefca1},
  {32'hc4102098, 32'h44af18de, 32'h43d6a0fa},
  {32'hc405866f, 32'hc1941f66, 32'hc3aa8e76},
  {32'hc2b30f20, 32'h45455aea, 32'h42a0d463},
  {32'h42d60e90, 32'hc4a4a594, 32'hc4cfbf19},
  {32'hc366fafe, 32'h43b1a406, 32'h44c8581e},
  {32'h451f9aac, 32'hc337c92d, 32'hc376fbd3},
  {32'hc56b1d01, 32'h42725949, 32'h42a9ac88},
  {32'hc480a2c6, 32'h419967ce, 32'hc31900f7},
  {32'hc341faa3, 32'hc400b677, 32'h44a89167},
  {32'hc388b01b, 32'hc3983646, 32'hc4ab14f3},
  {32'hc2b49ae8, 32'h4507a145, 32'h434fe0c9},
  {32'hc293f680, 32'hc425f120, 32'hc30db7de},
  {32'hc4c4949b, 32'h444febc4, 32'hc3598fea},
  {32'h43dcafdc, 32'hc3037d26, 32'hc4746746},
  {32'hc48db0f3, 32'h43154f36, 32'h445f000c},
  {32'h42fa0620, 32'hc38e2a54, 32'hc55c3940},
  {32'h43baac9e, 32'h4396216f, 32'h43d4943d},
  {32'h43a384ee, 32'hc45d2b35, 32'hc40864b8},
  {32'hc43bede8, 32'h45260ff7, 32'hc20f652c},
  {32'h43baa468, 32'h4359ca58, 32'h430298e5},
  {32'hc4fef04a, 32'h445d0753, 32'h4338e7ec},
  {32'h4331547c, 32'hc546089f, 32'h43965cd6},
  {32'hc4d82dd9, 32'h442d1d3e, 32'hc262deea},
  {32'h45261bca, 32'h4391959f, 32'h438449f9},
  {32'hc58a4be0, 32'hc22a6dea, 32'hc3b3e287},
  {32'h4508a906, 32'h42565b10, 32'h42cd0183},
  {32'h44cbfc69, 32'hc2f32152, 32'hc389f42f},
  {32'hc419eb76, 32'h433c51b7, 32'hc4be2184},
  {32'h44f88c90, 32'hc35882da, 32'h44856a1d},
  {32'hc421c9fa, 32'hc3011fea, 32'h42850cca},
  {32'h453e2175, 32'h433143c2, 32'hc3068947},
  {32'hc20459a0, 32'h4541aebf, 32'h43e4cf61},
  {32'h4406e194, 32'hc46da2d5, 32'h439e3cb9},
  {32'hc50c773c, 32'h4465c630, 32'hc13cc0fc},
  {32'h440ea77c, 32'hc4a98907, 32'h428e71b8},
  {32'hc4a2c06b, 32'hc3900cb8, 32'h410151e6},
  {32'h448ac2ea, 32'h4394ff98, 32'h4381fc1c},
  {32'hc521046a, 32'h4329bdba, 32'h42be3b3f},
  {32'h4398776a, 32'hc4ed4803, 32'h42efa62a},
  {32'h42408cb0, 32'h4488f183, 32'h4490494f},
  {32'h421ca9c8, 32'hc4d046c3, 32'hc49364bb},
  {32'h442c14d6, 32'h43a91fae, 32'hc1154ef8},
  {32'h444be4dc, 32'hc4398162, 32'h431628d3},
  {32'hc4393764, 32'h433bf65a, 32'h436d5bef},
  {32'hc4a31210, 32'hc414f293, 32'hc2d3b2c8},
  {32'hc574dd5b, 32'h438c5058, 32'h4306b1d2},
  {32'h4469a884, 32'hc4015e16, 32'hc4b80a51},
  {32'hc2eb1628, 32'h4387c784, 32'h44bacf49},
  {32'h424c5c48, 32'hc43dc253, 32'hc4f714d6},
  {32'hc4ca4cfd, 32'h430b8cb7, 32'h44555a50},
  {32'h44b226d2, 32'hc40b19e8, 32'h4201f33b},
  {32'hc49afd3a, 32'h44c82cbe, 32'hc33c61a6},
  {32'h4417c964, 32'hc35c1723, 32'hc559fd89},
  {32'h44e772ea, 32'hc18e99ff, 32'h42420614},
  {32'hc571e30a, 32'hc3d8e63d, 32'hc386b012},
  {32'hc1b694be, 32'h4474b607, 32'hc4b2d643},
  {32'hc5013dc2, 32'hc291c1f2, 32'hc268159e},
  {32'hc388e033, 32'h454736a2, 32'h43aeb047},
  {32'h44068a6a, 32'hc3c99b5f, 32'hc40db353},
  {32'h453fd355, 32'h4452aea8, 32'hc38f670c},
  {32'hc308dd00, 32'hc55fa345, 32'h43bc7e2c},
  {32'hc3eb9bd3, 32'hc3cd5410, 32'h432ce73e},
  {32'hc48c8d8b, 32'hc3d4aa2b, 32'hc38a3e7d},
  {32'h4524761e, 32'hc335e237, 32'hc2a15123},
  {32'hc393d5fc, 32'hc2a41347, 32'h449bee4a},
  {32'h4477753c, 32'h4443569c, 32'hc26d1993},
  {32'h4367a008, 32'hc52a45e9, 32'hc3e3b40e},
  {32'h43aa105d, 32'hc37d90f8, 32'hbe20c200},
  {32'hc3a33e30, 32'hc496eba5, 32'hc36120b5},
  {32'h41804e40, 32'h44c792c8, 32'h436a60ea},
  {32'h43b7d452, 32'hc41d707f, 32'h436f5757},
  {32'h44ef7ebe, 32'hc299dd5c, 32'h449968af},
  {32'hc48c4349, 32'hc47e1792, 32'hc49b7923},
  {32'hc496c9f8, 32'h4341e173, 32'h4372bd7d},
  {32'hc50d2e44, 32'hc431507f, 32'h41afe3bc},
  {32'h45214538, 32'hc2274afa, 32'h4399988d},
  {32'hc304d140, 32'hc337686c, 32'hc398a24e},
  {32'h4525dfbd, 32'h438ea2f2, 32'h437eb87f},
  {32'hc3dcf6c8, 32'hc4b2b2d0, 32'hc43d6c3b},
  {32'h43409ac6, 32'h44921d49, 32'h43cd5ad0},
  {32'h4485349e, 32'hc3533141, 32'hc3a305c4},
  {32'hc4073e34, 32'hc539df6b, 32'h42fbaea5},
  {32'h451b2caa, 32'h4391ae54, 32'h44075246},
  {32'h44b88c88, 32'hc3b52c96, 32'h4390d09f},
  {32'h452e4920, 32'h434c49fd, 32'hc3020f7a},
  {32'hc4830734, 32'hc492ea9e, 32'h42efade4},
  {32'h44e30cef, 32'h41aa3eb5, 32'hc42bd590},
  {32'hc590ab75, 32'h43a6d191, 32'hc3ab5ca8},
  {32'hc29cf040, 32'h42932f31, 32'h43ed2887},
  {32'hc522b9ac, 32'hc3b3939f, 32'h431b0f06},
  {32'h4235d660, 32'h418d64c0, 32'h441ee61b},
  {32'hc5126dee, 32'h4262f6be, 32'hc396731a},
  {32'hc1b13f76, 32'h4512e92d, 32'hc299d9c7},
  {32'hc377d4e4, 32'hc426e6f5, 32'h44be3aab},
  {32'h44e42ef4, 32'h43b84e3e, 32'hc35b7c53},
  {32'h44d4d96a, 32'h432afef1, 32'h4322e77a},
  {32'h41b4f6e0, 32'hc46b18c8, 32'hc518f5fe},
  {32'hc3f3b28a, 32'h42d5aeef, 32'h44b3b3f3},
  {32'h43d30ab0, 32'h44ac6a75, 32'h420859f3},
  {32'hc56f4d0c, 32'hc38ba5f5, 32'h43282618},
  {32'h418f2110, 32'h449663be, 32'hc5100c1d},
  {32'hc5389795, 32'h434309c5, 32'hc2c141dc},
  {32'h44c7840c, 32'h441c4c7d, 32'hc33eeb4e},
  {32'hc2366800, 32'hc51754fe, 32'h4386c9ae},
  {32'h44a7f865, 32'h43865ffb, 32'hc4aacc51},
  {32'hc50f6304, 32'h412f61c3, 32'h44933c8c},
  {32'h42673400, 32'hc3611e09, 32'hc474e39a},
  {32'hc273a56b, 32'hc5445cfc, 32'hc3384516},
  {32'hc31c07b6, 32'h453435a8, 32'h43f2d009},
  {32'h445b6f43, 32'hc4608b62, 32'hc14a42f8},
  {32'hc3b862be, 32'h44d43193, 32'h423d8472},
  {32'h44e5524d, 32'hc36d4e92, 32'hc35e4ae3},
  {32'hc468f6a5, 32'h41a85ce8, 32'hc2d80575},
  {32'h4534bdd8, 32'hc3dd0c71, 32'hc42d2f2c},
  {32'hc425f92a, 32'h43fb5745, 32'h4414fd42},
  {32'h44ed16ea, 32'hc3e3f03e, 32'h43d27ace},
  {32'hc3839eb2, 32'h43fd3f28, 32'hc50e7a38},
  {32'h431a1f0d, 32'hc4f10bdd, 32'h44836884},
  {32'h4300e210, 32'hbf103ce0, 32'hc35d8e38},
  {32'h430712a6, 32'hc4c412c5, 32'h44388f1a},
  {32'hc4fbd188, 32'h43f71f1f, 32'hc46626e4},
  {32'h45023e04, 32'h42ca4798, 32'hc3a37810},
  {32'hc38df6f0, 32'hc3e3bf53, 32'hc494fe22},
  {32'h450332db, 32'hc3e650dc, 32'h43a86e2b},
  {32'hc3fe57e8, 32'hc39c810c, 32'hc4c9d09f},
  {32'h43021608, 32'hc54ce7c2, 32'hc3092b8b},
  {32'hc4a33cb9, 32'h44833f6b, 32'hc50c429f},
  {32'h437f6899, 32'hc4059cd2, 32'hc0c6e735},
  {32'hc3eadbd6, 32'h454430b1, 32'h43178821},
  {32'h45139519, 32'hc4065219, 32'h423e788c},
  {32'hc4d3be20, 32'h43c91e39, 32'h438bafba},
  {32'h43976140, 32'h4403c47d, 32'h45347e1e},
  {32'hc4f15c37, 32'hc41bc920, 32'hc49838f7},
  {32'h456aaec4, 32'h43c35800, 32'hc40b610d},
  {32'hc47c3e51, 32'hc49e6c68, 32'hc480e89d},
  {32'hc199b2c0, 32'h43879101, 32'h4530f6c8},
  {32'hc3017b48, 32'hc439aa11, 32'h42b1e8d0},
  {32'hc3af0fe7, 32'h44c9965c, 32'h42e81453},
  {32'h42ebec1d, 32'hc39af1f0, 32'h435663cc},
  {32'hc33bf35a, 32'h44ba18d1, 32'hc3f086e8},
  {32'hc3f3790e, 32'hc4893fee, 32'h4311c754},
  {32'h4361ce84, 32'h45174392, 32'hc3ae526d},
  {32'h443c9866, 32'hc35364b0, 32'h44a7b644},
  {32'h41f9ad94, 32'h44fe8146, 32'h44c33392},
  {32'hc4a8029b, 32'h44ac31fd, 32'hc4ba2742},
  {32'h44a7d21e, 32'h43cb4465, 32'hc3f9b9c8},
  {32'h41808420, 32'hc45ce7d7, 32'h41a6425b},
  {32'hc44f0358, 32'h4480c613, 32'h432b6eb5},
  {32'h44d42146, 32'hc287c16e, 32'h44094901},
  {32'h443614ae, 32'h4490d3ae, 32'hc2fad893},
  {32'hc24b1b68, 32'hc53e4297, 32'hc3892aaa},
  {32'hc3a200d0, 32'hc34e700b, 32'hc52534e5},
  {32'hc495b5c4, 32'hc3eb89be, 32'hc36a973d},
  {32'hc4abb8ed, 32'h43adc286, 32'hc42662e8},
  {32'h4522bd74, 32'h43b4d1da, 32'h418a80d8},
  {32'hc48c5c1d, 32'hc365c734, 32'hc28ec7d7},
  {32'hc381c532, 32'hc560cfdc, 32'hc3299d91},
  {32'hc38d7180, 32'h44c167e5, 32'hc31ce586},
  {32'h44b6959a, 32'hc42ce727, 32'hc2cf2cf6},
  {32'hc38ec784, 32'h4549ae4b, 32'h43a8ff4e},
  {32'hc23c9480, 32'hc4ff0e62, 32'hc3e68ca5},
  {32'h44b3c73c, 32'hc37ebd5f, 32'h4397f1a7},
  {32'h42d901b0, 32'hc43a4859, 32'hc4d0ae9f},
  {32'hc3135ed0, 32'hc38f2770, 32'h44a86ba3},
  {32'hc2f79eb2, 32'hc4ade5ed, 32'h4326b124},
  {32'h41d5de37, 32'h44ad39c6, 32'h4336c605},
  {32'hc382f0c4, 32'hc4205f2c, 32'hc3b62ce0},
  {32'h448e6178, 32'h44c6f12b, 32'hc33827de},
  {32'hc39b3510, 32'hc45151d4, 32'h440bf407},
  {32'h435dec2e, 32'h43dc28b5, 32'h430ffa1e},
  {32'h439c304b, 32'h4495d395, 32'hc3a39824},
  {32'hc4456d10, 32'hc48c270b, 32'h44cd7003},
  {32'h448b62e7, 32'hc43025c9, 32'hc4a9c2a9},
  {32'h43e9697e, 32'h4433edd5, 32'hc45fb3dc},
  {32'hc5246b5f, 32'h43286437, 32'hc2cc1cd9},
  {32'hc43c5d3b, 32'h42e40587, 32'hc439f49f},
  {32'hc5033bba, 32'hc441778a, 32'h43d7a9d9},
  {32'h423e6148, 32'h4413a2a1, 32'hc528bce7},
  {32'h431bbbc6, 32'hc3c4185a, 32'h43729c1c},
  {32'hc1c21780, 32'hc469a21a, 32'hc40bee4d},
  {32'hc5219d32, 32'hc1bcc194, 32'hc1910b48},
  {32'h4528e46d, 32'h4302466a, 32'h43ad4f9a},
  {32'hc4d708d0, 32'hc3c9c6e1, 32'hc369510e},
  {32'h44bd1988, 32'h43d29dd3, 32'hc31ffe6d},
  {32'hc401f192, 32'hc3fe1c0c, 32'h4286af27},
  {32'h4465e6fa, 32'h44bf66b5, 32'h4404658b},
  {32'hc3bd45ac, 32'hc519eb45, 32'h4346f083},
  {32'h444d900f, 32'h43ef1aa6, 32'hc40ef6cf},
  {32'hc4bb6573, 32'h41f46686, 32'h436fa281},
  {32'hc308be2e, 32'hc3e2ccb0, 32'hc488ef67},
  {32'hc3ba1a58, 32'hc4bb4b57, 32'h44d3b2e7},
  {32'h4399c23a, 32'hc424754d, 32'hc2eaf2f4},
  {32'h42cf44c0, 32'h45328ca8, 32'h43f654a1},
  {32'h42ec49d7, 32'hc40b6213, 32'hc4a0103f},
  {32'hc3179980, 32'h44943e43, 32'h443e1882},
  {32'hc427f228, 32'hc40ef4e4, 32'hc4e4659a},
  {32'h440d1cc6, 32'h44a6f5f9, 32'h44a1c4b9},
  {32'h438646a3, 32'h43e5581a, 32'hc4f6c6ce},
  {32'hc409da38, 32'h42f3c792, 32'h44ab7e15},
  {32'hc3932ca2, 32'hc4d7da2d, 32'hc412748a},
  {32'h451b9b81, 32'hc2b37359, 32'h438db9c8},
  {32'hc558b81e, 32'hc40dc5c3, 32'h43820b73},
  {32'h444ae5cd, 32'h447976e9, 32'hc3d59cca},
  {32'h4394f462, 32'hc4b825cf, 32'hc43cc1f1},
  {32'hc39074bc, 32'h44a98ead, 32'h4502f064},
  {32'hc4fe4ac0, 32'h41da6ceb, 32'hc383d462},
  {32'hbf32a53c, 32'h44f3ebdb, 32'hc38c9096},
  {32'hc5201cc0, 32'hc433da6f, 32'hc2046c50},
  {32'h42cbc6d6, 32'h45681b2e, 32'hc36d72df},
  {32'hc4832105, 32'hc31b7744, 32'h4399f55f},
  {32'h4386c9cc, 32'h438bbf46, 32'hc4456379},
  {32'hc5111a78, 32'hc17975b8, 32'hc3885e22},
  {32'hc3c5ca88, 32'h4387e620, 32'hc1b842c7},
  {32'hc4e177f0, 32'hc3acd1ad, 32'h41a3f385},
  {32'h43a26998, 32'h432ac263, 32'hc2a74d97},
  {32'h43303a1f, 32'hc516b6d1, 32'hc4598f25},
  {32'hc4fd7412, 32'hc4415c21, 32'h4408202c},
  {32'hc3bba8b3, 32'h4491affd, 32'hc3eb1350},
  {32'hc526f023, 32'h4463b7c5, 32'h439eefb1},
  {32'hc3cb37f0, 32'hc458fd7c, 32'hc4d62fbe},
  {32'hc32b2008, 32'h44c6e0d7, 32'h427c9fe9},
  {32'h44aa9617, 32'h427b652d, 32'h41bd7284},
  {32'hc41567c0, 32'hc37c7dae, 32'h443ac13f},
  {32'h4418c745, 32'hc41ea4fe, 32'hc36b97b7},
  {32'hc46152f6, 32'h445d6dc9, 32'h43fe5251},
  {32'h43605920, 32'hc437a147, 32'hc4777837},
  {32'hc4004caa, 32'hc37a8107, 32'h44a2ef39},
  {32'hc3be44eb, 32'hc4d6df3a, 32'hc3e3d61e},
  {32'hc4a5e5b4, 32'h4386d6fe, 32'h4493f7fb},
  {32'hc3c9e3c9, 32'hc48a1c31, 32'hc3756821},
  {32'h438682b4, 32'h42381500, 32'h450991d1},
  {32'hc2bef5ce, 32'h42b80dcd, 32'hc4ce683c},
  {32'hc415d8b0, 32'h430be9c1, 32'h4244a7e2},
  {32'h44b89ceb, 32'hc4ad2f2f, 32'h43c78844},
  {32'hc53344b1, 32'h443da3b0, 32'hc2973149},
  {32'h453fc9ef, 32'h4416ed9d, 32'h43b504fb},
  {32'hc537bac6, 32'h4366d5c9, 32'h42fa29f3},
  {32'hc3397bdc, 32'hc512020d, 32'hc40112d4},
  {32'hc4c288bc, 32'hc281caa9, 32'hc309e6e4},
  {32'h453c46ef, 32'h44006382, 32'hc213af07},
  {32'hc488185b, 32'h43bb6b00, 32'h43e73851},
  {32'h44f0e7fe, 32'hc2dd1ffb, 32'hc2f2a511},
  {32'h44a1a2bc, 32'h434ae54f, 32'hc22b2a84},
  {32'hc4330992, 32'h4347aefa, 32'hc4b830ea},
  {32'h4413ae7e, 32'hc4278eb0, 32'h449c4f56},
  {32'hc355a768, 32'h4429f3de, 32'hc35d9aeb},
  {32'h44e1c7f5, 32'hc3f71d76, 32'hc3521420},
  {32'hc4d5dda2, 32'h443b4e97, 32'h42d6861b},
  {32'h4458445a, 32'hc4009322, 32'hc320fe82},
  {32'hc481c71a, 32'h44b83e6e, 32'hc10393ab},
  {32'h44be008a, 32'hc4d913a5, 32'hc1c3994c},
  {32'h43916579, 32'hc4400f80, 32'h42ff73ae},
  {32'h44ea0c3d, 32'h4298df19, 32'h43b1c779},
  {32'hc4ce49d7, 32'h43942ccc, 32'hc3571581},
  {32'hc383f368, 32'hc3f0be4e, 32'hc3e90ffb},
  {32'hc428b954, 32'h441b4792, 32'hc2c1648c},
  {32'h44b007ca, 32'hc324b298, 32'hc43531a9},
  {32'hc31b64bc, 32'hc24da515, 32'h43a8bc36},
  {32'h4086c900, 32'hc3290577, 32'hc50232f5},
  {32'hc4880456, 32'h439654eb, 32'h44fcb01e},
  {32'h44f3e84f, 32'hc3c9786d, 32'h4333a277},
  {32'hc5578a14, 32'hc3100c9f, 32'h43e94ac8},
  {32'hc34373b0, 32'hc28cb9dc, 32'hc423018c},
  {32'h442b4822, 32'h443ded75, 32'h435fb6cc},
  {32'hc3162fd8, 32'hc404fa8f, 32'hc50ec5ec},
  {32'hc4580c73, 32'h44a28951, 32'h4493d2f4},
  {32'h42f898ac, 32'h41ef7c3c, 32'hc43e5cdf},
  {32'hc4c19886, 32'h445b7059, 32'h43a08acb},
  {32'h4407e29d, 32'hc4518219, 32'hc4e21b2e},
  {32'h43fe6890, 32'hc375f027, 32'hc4de4912},
  {32'hc46c47ae, 32'hc37bc975, 32'h452cd2f6},
  {32'hc497a6ec, 32'h42c7b002, 32'h43a82de1},
  {32'hc47c9684, 32'hc4a56094, 32'hc3ca9b02},
  {32'h44272e52, 32'h45135d0a, 32'h43f4a00e},
  {32'hc3f03f48, 32'hc424fcc6, 32'h43a4c715},
  {32'h45072eea, 32'h442fd0e5, 32'hc3b99489},
  {32'hc4512617, 32'hc456ffd3, 32'hc233f67b},
  {32'hc2648353, 32'h44c15fe7, 32'h42dde512},
  {32'hc474e04c, 32'hc3e364a9, 32'hc3bcf91e},
  {32'h44508641, 32'hc1d54154, 32'hc5148c09},
  {32'hc42f974a, 32'h4281cfce, 32'h44605123},
  {32'h450a6238, 32'h43bea7e7, 32'h43aac046},
  {32'hc428ac9f, 32'hc3a63f9c, 32'hc5429214},
  {32'h448ff950, 32'h44504618, 32'hc26f8f91},
  {32'hc3dde7fe, 32'hc501d0f1, 32'hc4476dd2},
  {32'h451e8bd7, 32'h421e2d67, 32'hc28b33d8},
  {32'h424aa35a, 32'h42929393, 32'hc4f2fc4b},
  {32'hc3dba3d5, 32'hc1663cca, 32'h44668023},
  {32'hc4e1fd0c, 32'h43b9f5c2, 32'hc3a0ab9a},
  {32'hc4a1021f, 32'hc3587d92, 32'h42e5db5d},
  {32'hc3e50cc8, 32'hc4b99cb6, 32'hc3d2db83},
  {32'h431dfd38, 32'h43a5de0b, 32'h44c90feb},
  {32'h4421294b, 32'hc40cc633, 32'hc410f85f},
  {32'hc3d744a5, 32'h42a6fe2f, 32'h453c12e4},
  {32'h42a52208, 32'hc2257b51, 32'hc560f8c5},
  {32'h43d37e92, 32'h44443c1b, 32'hc2ca2409},
  {32'h4521d94a, 32'hc3911e9b, 32'hc2133c88},
  {32'hc4df8d48, 32'h42f8d192, 32'hc44d4a58},
  {32'h44ac64c1, 32'h448a5bcb, 32'h44245c2f},
  {32'hc4de3750, 32'hc2d3e6f8, 32'h4363baf8},
  {32'h44f0410b, 32'h44ab0e5b, 32'hc2ce1e50},
  {32'h43db0d38, 32'hc53867b3, 32'hc2992880},
  {32'h45286098, 32'hc2d1c601, 32'hc40486da},
  {32'hc55bd016, 32'hc2d1dd4f, 32'h438e23fa},
  {32'h4570198d, 32'h43d9f743, 32'h44327b50},
  {32'hc4532c98, 32'hc39ff1fb, 32'hc20b99e7},
  {32'h4427c294, 32'h44929b72, 32'hc2e4d62d},
  {32'hc454c452, 32'h4482c021, 32'hc4eb0cc3},
  {32'hc3972c1e, 32'h444afbc8, 32'h42989be2},
  {32'hc49bfa11, 32'hc37a5ec0, 32'h43ba906c},
  {32'h444e652c, 32'h4406aab6, 32'hc485fc4f},
  {32'h4389ea8c, 32'hc352b80a, 32'h44cff69d},
  {32'h44bf0a60, 32'hc3c12971, 32'hc3d05721},
  {32'hc306c0f4, 32'h43b9f32e, 32'h4566122d},
  {32'h4487b071, 32'h4417686a, 32'hc38c5096},
  {32'hc4639249, 32'hc490b63c, 32'h43cd3843},
  {32'h43a5404c, 32'h445cf78f, 32'hc49b0adc},
  {32'hc50b7497, 32'hc38097bf, 32'hc39f307c},
  {32'h4280c70a, 32'h45082562, 32'hc43613fd},
  {32'hc47eea30, 32'hc406b1b8, 32'h44a22e3b},
  {32'h44642ce3, 32'h42bcb5fe, 32'hc31dfada},
  {32'hc1933a60, 32'h441cfe07, 32'h456ced5e},
  {32'h43927ca2, 32'hc42dec2b, 32'hc517b338},
  {32'h453b1c7d, 32'hc3ef07cc, 32'h4310d378},
  {32'hc4728e20, 32'h44c3f7b8, 32'h437b3928},
  {32'h4428a91d, 32'hc39faa7e, 32'hc10a90a0},
  {32'hc341fdc7, 32'h44201cb5, 32'h43fd4ca6},
  {32'h43ca2246, 32'hc2974667, 32'hc44c3330},
  {32'hc4cddee3, 32'hc38603ad, 32'hc3760acc},
  {32'h44e65b79, 32'hc400b5ca, 32'hc3ddeafa},
  {32'hc5896702, 32'hc3245304, 32'h43fccee5},
  {32'hc4d2433d, 32'h404f2fbc, 32'hc301e6e7},
  {32'hc48021d7, 32'h42028075, 32'h43f8fa3a},
  {32'hc13c0c60, 32'hc4f915ba, 32'hc29a55c3},
  {32'h4324e156, 32'h444ca7e0, 32'hc3696e3b},
  {32'h43d1dee2, 32'hc3d12547, 32'h44f24bd8},
  {32'hc3d1b2fa, 32'h45129e33, 32'h43a4b413},
  {32'h4408cab1, 32'hc4271cb6, 32'h441909a7},
  {32'hc4ff5f64, 32'h42a11a38, 32'hc29d179c},
  {32'h450d89d2, 32'h438e7269, 32'h44033a11},
  {32'hc48f617a, 32'h42b1fd12, 32'hc4079d80},
  {32'h44362f62, 32'hc51003cc, 32'hc393d8e8},
  {32'hc503630b, 32'h4408dd64, 32'hc4574a42},
  {32'hc41cd5ad, 32'hc38cf446, 32'h437e5ca8},
  {32'h3f368800, 32'h441df8f1, 32'hc4db3551},
  {32'h43c9f919, 32'hc4d61506, 32'h43b1270d},
  {32'hc4c11487, 32'h423f77c0, 32'hc3b6f7eb},
  {32'h448336f9, 32'h43efedc8, 32'h447a64de},
  {32'hc4c6a9b4, 32'h424b1c28, 32'hc4c0665b},
  {32'h43baa3d0, 32'hc33440dc, 32'h450f189c},
  {32'hc37c2da4, 32'h428fb2a9, 32'hc4856b8a},
  {32'hc2d8e01c, 32'h44c95208, 32'h44ebc6b3},
  {32'hc2401ecb, 32'h42a8feea, 32'h43a739bb},
  {32'hc5195fba, 32'h423444f1, 32'h43963949},
  {32'h44105307, 32'hc46d0f71, 32'h445efddd},
  {32'hc2e99c9c, 32'h4432f9c0, 32'hc46b2193},
  {32'h44c048cb, 32'hc38c0378, 32'hc3249e6c},
  {32'hc4d92fde, 32'h44984d34, 32'h43853895},
  {32'h44e7c538, 32'hc479457a, 32'h44090d43},
  {32'h43b8a700, 32'h44832a73, 32'h44924f34},
  {32'hc315c2cf, 32'h4510b266, 32'hc4fdad1d},
  {32'h445a9d71, 32'hc4114c43, 32'hc39d61a3},
  {32'hc393da46, 32'hc4a8b85e, 32'h42f8288f},
  {32'hc516fa15, 32'h4343fb2f, 32'hc3ebcd50},
  {32'h441695d7, 32'hc358ad9e, 32'h43867132},
  {32'h433565b0, 32'h433ff572, 32'hc3d19c15},
  {32'hc36620ea, 32'h42db4e1a, 32'hc32a9f7d},
  {32'hc2c7bcb4, 32'h4508c366, 32'hc318663a},
  {32'h44e3e381, 32'hc3351821, 32'h4183ff00},
  {32'hc50dd2e0, 32'hc470350a, 32'hc3f41552},
  {32'h44bd86dc, 32'hc3db1777, 32'h44521eaa},
  {32'hc48f7e0c, 32'h4407abb0, 32'h43a0712f},
  {32'h45783295, 32'hc38d58b9, 32'h4288487f},
  {32'hc4a57b74, 32'h44744557, 32'h438dc00a},
  {32'hc41bbcaa, 32'hc3ba05c2, 32'h42ac8187},
  {32'hc5554d2a, 32'h43f465a1, 32'hc407029d},
  {32'h43cc501a, 32'hc4eba112, 32'h43ce8e55},
  {32'h441fedee, 32'h44d45b80, 32'h4353e1d6},
  {32'hc334f625, 32'hc44a39ed, 32'hc4c47276},
  {32'hc290aaac, 32'hc2cb1022, 32'h450717bf},
  {32'hc31a4f15, 32'hc48d88d3, 32'h42c67893},
  {32'h433e5320, 32'h44000ae2, 32'hc4258fba},
  {32'h4430b1e8, 32'hc4510236, 32'h42d8bb2d},
  {32'h44ef9e01, 32'h43ec50b6, 32'hc4132932},
  {32'h42161538, 32'h439ce3fd, 32'h45527109},
  {32'h45321b2e, 32'hc3d052fd, 32'hc325cf77},
  {32'hc48ce563, 32'hc432e3d9, 32'h4305777b},
  {32'hc4806289, 32'h4482362f, 32'h447f0207},
  {32'h4406e2d5, 32'h43236688, 32'hc4b8d918},
  {32'h43cc8ea3, 32'h44491ad1, 32'hc1ca3487},
  {32'hc3b06597, 32'hc4b08eb7, 32'h4405e726},
  {32'h440e24f0, 32'h449a0b61, 32'hc4972bf7},
  {32'hc4327d25, 32'hc42ebfb3, 32'h44e7dd47},
  {32'h44dd237d, 32'h435cefc8, 32'h4212c0b8},
  {32'h43d26a0a, 32'hc495f5a8, 32'hc2ca3f59},
  {32'h45822969, 32'hc3b36be1, 32'hc36ae708},
  {32'hc59c4715, 32'hc2b8f26b, 32'hc3c96d4e},
  {32'h44fd98e0, 32'h43e26acc, 32'h43121329},
  {32'hc382785c, 32'hc5159124, 32'hc2dc9063},
  {32'h448ef1eb, 32'h449047bb, 32'hc39c47db},
  {32'hc3228e80, 32'hc3654804, 32'h440e4a39},
  {32'h441b1de6, 32'h452192f2, 32'hc3d5dcb4},
  {32'hc5694edb, 32'hc37d7bfc, 32'h40cafa7e},
  {32'hc2c793ff, 32'h44e6bd60, 32'h42d4b5d2},
  {32'h44c61e6c, 32'hc368cf40, 32'hc3f3b9a7},
  {32'h438e27df, 32'h449c7696, 32'hc4fe432f},
  {32'h4405c363, 32'hc4b93911, 32'h44bf5a26},
  {32'hc40af0d9, 32'hc320d8aa, 32'hc41602d6},
  {32'h442406c8, 32'h419b09fc, 32'h446eb294},
  {32'h41d76a7b, 32'hc3a001c6, 32'hc482f6c2},
  {32'h4533c5ca, 32'hc328e91a, 32'h43e2086b},
  {32'hc4866a40, 32'hc4c0562a, 32'hc4d7d370},
  {32'h437d6242, 32'hc3ae9096, 32'h4460afd2},
  {32'hc2bfc699, 32'h44863cee, 32'hc4c6b70d},
  {32'hc4a0fc85, 32'hc44e4a43, 32'h4525d46c},
  {32'hc3d72fee, 32'h450b8b37, 32'hc4ff16d9},
  {32'h435064d0, 32'h44b0edc3, 32'h430a1cfa},
  {32'hc38382ec, 32'hc280bc5b, 32'hc340000a},
  {32'h43f12528, 32'h455209ff, 32'h409d6f6e},
  {32'h43487e5a, 32'hc4ab95ae, 32'hc47a7917},
  {32'h42249600, 32'h44f072ed, 32'h44e43e22},
  {32'hc3f5b1f4, 32'hc41846be, 32'hc5154892},
  {32'h450d78d0, 32'h42fef756, 32'h4331de7d},
  {32'hc498f021, 32'hc48d821a, 32'hc3fd1a17},
  {32'h44f752d6, 32'h44760ae0, 32'hc38a5f47},
  {32'h4501de2d, 32'hc30f8169, 32'hc34059cb},
  {32'h44f18a0e, 32'h42aeb764, 32'hc3b0ff9d},
  {32'hc4fa9272, 32'hc4086dcd, 32'hc25013bf},
  {32'h427fc1c0, 32'h41cae6f6, 32'h41b6b074},
  {32'hc4f19c47, 32'h4337e9af, 32'h4400de66},
  {32'h4559ad59, 32'h421e0904, 32'h43440996},
  {32'h443bd582, 32'hc4624e9e, 32'hc4441e76},
  {32'h423cabd4, 32'hc4ab3deb, 32'h44bd9d66},
  {32'h43666506, 32'hc15fb5ce, 32'hc34257bf},
  {32'hc43b349e, 32'h44ee211c, 32'h41815eac},
  {32'h43a0fef4, 32'hc42267b4, 32'hc419678c},
  {32'hc3fec208, 32'h4250eadd, 32'h448b4386},
  {32'h41b77d00, 32'hc3b6b1a1, 32'hc53ad6c0},
  {32'hc50eea3c, 32'h4359f7f1, 32'h4481b60e},
  {32'hc40c9d60, 32'hc4012a80, 32'hc27410d7},
  {32'hc3c4e9ab, 32'hc4253705, 32'h445ea2f9},
  {32'hc2905132, 32'hc4c01662, 32'hc409c546},
  {32'hc3e6041a, 32'hc49f13d7, 32'h4437861a},
  {32'h43722ed7, 32'hc4fac360, 32'h42cd5ddd},
  {32'hc3ec2100, 32'hc13332be, 32'h426468c6},
  {32'hc4d168b1, 32'hc326b25e, 32'h4266a3fa},
  {32'hc51b2e8a, 32'h433853a0, 32'h43882e80},
  {32'hc3d666cb, 32'hc405db36, 32'hc53b59de},
  {32'h4260b9be, 32'h44a34f11, 32'h444321ba},
  {32'h43304078, 32'hc44661f0, 32'hc43dfc5e},
  {32'hc4926fa7, 32'h448aedcd, 32'hc34d8df0},
  {32'hc215c26c, 32'hc4b9bfac, 32'h42902c03},
  {32'hc40c1210, 32'h4534b8b1, 32'h43b25a0f},
  {32'h44dafd6a, 32'hc480d6a4, 32'h4381ebe6},
  {32'h44ce38fb, 32'hc340bc8e, 32'h41973697},
  {32'h4495947d, 32'h439053b8, 32'hc2514fa1},
  {32'hc52cdc91, 32'h433a36c9, 32'hc2bcf592},
  {32'hc3a36322, 32'h4302200a, 32'hc412615e},
  {32'h43f890c4, 32'hc1649eb1, 32'h438143a4},
  {32'hc466a2f8, 32'hc3887b09, 32'hc489dc8d},
  {32'h44ea7c4b, 32'h43d6dba6, 32'h43d95adb},
  {32'hc31fb340, 32'hc386f108, 32'h43ee0082},
  {32'h450fd6f1, 32'hc4034fc8, 32'h43a55229},
  {32'hc35873cc, 32'h45671d2f, 32'h440d151e},
  {32'hc4ab4450, 32'hc39922b1, 32'h40b8aa48},
  {32'hc54f7287, 32'h4213603b, 32'h436aa429},
  {32'h451eee7a, 32'h43879807, 32'h43f1a45a},
  {32'h4462287f, 32'hc263d844, 32'hc44e2eb8},
  {32'h44c4c66e, 32'h4371fe47, 32'h43a586ec},
  {32'hc4156331, 32'hc3e6a255, 32'h441802b0},
  {32'h451215d8, 32'hc36bfec4, 32'h4319a728},
  {32'hc4e38048, 32'hc30ad215, 32'h43bf4469},
  {32'h4330e6f4, 32'hc5236030, 32'hc36371dc},
  {32'h444aa4ec, 32'hc3c81524, 32'h442aeee5},
  {32'h442223dc, 32'h43e37e6d, 32'hc5077913},
  {32'hc413b0a0, 32'h4496f397, 32'hc31bc8e9},
  {32'h4442472c, 32'h42f91e50, 32'hc45ee9da},
  {32'hc5865d72, 32'h43800b56, 32'h42909736},
  {32'h452ab0fa, 32'hc36a230b, 32'hc3bbd18f},
  {32'h43a9a9ed, 32'hc3061d4a, 32'hc33779fa},
  {32'h4462c814, 32'hc49c1476, 32'hc48fc808},
  {32'h4285dc5a, 32'h45055377, 32'h44ca505d},
  {32'h4549be3e, 32'hc328fa23, 32'h43151166},
  {32'hc4c2c322, 32'h43af91a6, 32'h44408cd3},
  {32'h45210e0b, 32'hc4461b7c, 32'h4281209a},
  {32'h44f66fc8, 32'hc3c94c64, 32'hc45b269e},
  {32'hc5132caf, 32'h43cc96e4, 32'h443dae6e},
  {32'h4460fbd6, 32'h44808238, 32'hc2ce35a0},
  {32'hc5427fd8, 32'hc47251d8, 32'hc44917ef},
  {32'h4484e39d, 32'h44696abe, 32'hc191ea73},
  {32'h43a86282, 32'hc4b0f38b, 32'h43faf9c9},
  {32'h42afe840, 32'h44eafd77, 32'h43c75396},
  {32'hc51383fd, 32'hc3b6b743, 32'h439a672b},
  {32'h44ed91de, 32'h4344e46a, 32'h44237768},
  {32'hc50a63ad, 32'hc4116f56, 32'h4334ad7c},
  {32'h45282cc0, 32'h43b3f482, 32'h43878ab1},
  {32'h44a34308, 32'h4398e16f, 32'h43579508},
  {32'h42ae68c4, 32'hc37f85a8, 32'h4551b06c},
  {32'hc2988810, 32'hc4c3ecf6, 32'hc3364bfe},
  {32'h43b29bfd, 32'h446dbde8, 32'h44128109},
  {32'hc3a82088, 32'hc351d150, 32'hc5524181},
  {32'h43b8e33c, 32'h4490466b, 32'h442f2a0d},
  {32'h42ea592c, 32'hc3dd25f9, 32'hc467ff63},
  {32'h45127caf, 32'hc3df4d67, 32'h434235ce},
  {32'hc4d40fa5, 32'h40f673d8, 32'hc2abe271},
  {32'h43f41abc, 32'h442ba1e8, 32'h41d25ad1},
  {32'hc3ee4e80, 32'hc3fef68a, 32'hc41e7394},
  {32'h44bda23d, 32'h43bc08e8, 32'h442406ac},
  {32'hc444a714, 32'hc3fd0069, 32'hc40b22aa},
  {32'h4533fafe, 32'h438ec56b, 32'h43679770},
  {32'hc478f4f9, 32'hc4adfacd, 32'hc43308d5},
  {32'hc49b3df0, 32'hc305a622, 32'h403acf08},
  {32'h4283c048, 32'hc21e918a, 32'hc41da8ca},
  {32'hc3eb3154, 32'hc4a4ef94, 32'hc3339157},
  {32'h43b03c28, 32'h449adacd, 32'h44545f58},
  {32'hc435777c, 32'h43a96530, 32'hc35bbb9a},
  {32'h455043fd, 32'hc2531f3f, 32'hc405e7ed},
  {32'hc4663f4e, 32'hc4490f96, 32'h437d9918},
  {32'h452e658b, 32'h43c9ca2f, 32'hc3ce472d},
  {32'hc4b5dd83, 32'h44642148, 32'h43026480},
  {32'h442e0d80, 32'h43aaeaae, 32'h44436a9e},
  {32'h433ccb50, 32'hc45c59b4, 32'h441078db},
  {32'h43a6293c, 32'h44049573, 32'hc4b1358b},
  {32'hc4499098, 32'hc46bfffd, 32'hc2c3495f},
  {32'h44626273, 32'h442a5fc1, 32'h4338e26b},
  {32'hc38062bd, 32'hc37dd2f8, 32'h44e29191},
  {32'h443ca19e, 32'h452b0b86, 32'hc3cf8fde},
  {32'h4331ac01, 32'hc3329690, 32'h44f47f7d},
  {32'h45027b09, 32'h4405a2ef, 32'hc348faf3},
  {32'hc3dd06dd, 32'hc2d7fab1, 32'h4453d417},
  {32'h430e0a8a, 32'h44b0519e, 32'hc272d192},
  {32'hc50eaf1c, 32'hc4866cfb, 32'hc17f47ea},
  {32'h43b3fbe9, 32'h445d2796, 32'hc4e4803e},
  {32'h43be32ad, 32'h4339bc76, 32'h43e76008},
  {32'hc349911c, 32'h4516aa83, 32'hc12c2a00},
  {32'hc359621e, 32'h42f1d225, 32'h451a4444},
  {32'h4514113e, 32'h438cda58, 32'h4373217b},
  {32'hc579a49a, 32'hc3169787, 32'h421b3d24},
  {32'h438871a0, 32'hc4006184, 32'hc51352f3},
  {32'h45046ba6, 32'hc4518998, 32'hc3c81350},
  {32'hc553c053, 32'hc2c742e2, 32'hc3a4184f},
  {32'h43c8867d, 32'hc35c701e, 32'hc1af4837},
  {32'hc4e73562, 32'h42a116d4, 32'h43ab32ed},
  {32'h448a609a, 32'hc4903050, 32'hc3974cfa},
  {32'h4414dac6, 32'h421f0eda, 32'hc325e6c0},
  {32'h4536545a, 32'hc3980bcb, 32'hc3c32e66},
  {32'hc57ec2dd, 32'h4405ff2d, 32'h414ffd6c},
  {32'hc4b98d5a, 32'hc305f1cb, 32'h42c7e181},
  {32'hc3678100, 32'h445ec50e, 32'hc43e4df5},
  {32'h4470eb72, 32'hc49ae7f1, 32'h4396fb37},
  {32'hc3065aa4, 32'hc1c29f5e, 32'h43c132f4},
  {32'h430b4afe, 32'hc40d53c7, 32'h4308a96f},
  {32'hc233c0de, 32'h44aa09f4, 32'hc351a2be},
  {32'hc3ada976, 32'h42f45f40, 32'h44d991cc},
  {32'hc4b37e58, 32'h44814914, 32'hc35ad148},
  {32'h450d6558, 32'h43d92963, 32'h4382b563},
  {32'hc48d311e, 32'hc21ad443, 32'hc431c8c9},
  {32'h4525b651, 32'hc402635e, 32'h43151650},
  {32'hc5647aea, 32'h42c76d35, 32'hc33be268},
  {32'hc3c65455, 32'hc411f940, 32'h442a0e9b},
  {32'hc38c9f21, 32'h454fcb14, 32'h42b689bb},
  {32'h43ed6f58, 32'hc46ffa74, 32'h44c76f3d},
  {32'hc5095a10, 32'hc36f3b0f, 32'hc385dd9f},
  {32'h453044ae, 32'h433a0c2d, 32'h442d5a8a},
  {32'hc4b4bb80, 32'hc3608bad, 32'hc5080bb3},
  {32'hc4ac3163, 32'h438adb72, 32'h42a0c269},
  {32'h4325bcc0, 32'hc50cd13c, 32'hc5028e2a},
  {32'hc4efb10c, 32'hc311c43b, 32'h42fee96a},
  {32'hc482cb57, 32'h442e244f, 32'hc45cad8f},
  {32'hc4f5e4c8, 32'h43de624d, 32'hc2c085e9},
  {32'h44d28b68, 32'hc2b5fe1e, 32'h442cca0f},
  {32'hc4c48f9d, 32'h436202d4, 32'hc411fb3f},
  {32'hc4497546, 32'hc41c206c, 32'h438aba62},
  {32'hc42e6196, 32'h447e7ac2, 32'hc4d3ea19},
  {32'h44df349f, 32'hc41694f9, 32'h442427ab},
  {32'hc1a541b8, 32'h44456bb6, 32'h44d946c8},
  {32'h434098d9, 32'h421d5c68, 32'hc53806d8},
  {32'hc3c8933e, 32'hc41a64dd, 32'h4401d453},
  {32'hc44717da, 32'h43f5062c, 32'h43d5f2b3},
  {32'hc51f3a62, 32'hc353f304, 32'h4203c398},
  {32'h440a716c, 32'hc40b8622, 32'hc1eb0b2c},
  {32'h44d123d5, 32'hc39b6b94, 32'h43b2794c},
  {32'h440bfd90, 32'h4320900c, 32'h450d4f9e},
  {32'hc2b486cc, 32'h44c035f1, 32'h40d6b150},
  {32'h439b23d9, 32'h4320a7ba, 32'h4158094b},
  {32'hc3d76b20, 32'h4317cf5b, 32'hc4755e69},
  {32'h44d956fa, 32'hc3f16992, 32'h432c70dd},
  {32'hc3ba1312, 32'hc290371c, 32'h43117f45},
  {32'h4537a92d, 32'hc435773d, 32'hc305823a},
  {32'h43b2a33a, 32'h457373da, 32'hc2ec7022},
  {32'h43a4c5ca, 32'hc4c39da2, 32'hc3b37d11},
  {32'hc512c077, 32'h4486beec, 32'h43720eba},
  {32'h43748d02, 32'hc4a283c7, 32'h43c7e1a2},
  {32'h4417c96c, 32'hc30f6e41, 32'h4506c092},
  {32'hbfdc4700, 32'hc4ba0fbe, 32'hc481429d},
  {32'hc3ee5854, 32'h4404cbb0, 32'h44478d71},
  {32'hc48cba48, 32'h4400b644, 32'h44686711},
  {32'h430b5409, 32'h4507477c, 32'h40efa07e},
  {32'hc487d9be, 32'hc4fc101b, 32'h431f6c40},
  {32'h42b2fad0, 32'h4493ef2a, 32'hc4be511d},
  {32'h435b0090, 32'hc548bd53, 32'hc1b8aa8a},
  {32'h44af0b76, 32'h43f82d94, 32'hc3b19e41},
  {32'h43e428c9, 32'hc3e88ac6, 32'hc3b090e2},
  {32'h43ddb9c0, 32'hc3b759c4, 32'h45521289},
  {32'h42b27572, 32'h44dba017, 32'hc4fd72e8},
  {32'h4396cbd8, 32'h43750b81, 32'hc502cb20},
  {32'hc509f271, 32'hc3fd1017, 32'h43d15875},
  {32'h43ec2a26, 32'h451cae31, 32'h4310bb39},
  {32'hc541471d, 32'hc264ed3d, 32'hc1fa0a6b},
  {32'h42f7c2fa, 32'h45114814, 32'hc468ae7f},
  {32'hc3ae180b, 32'hc3961035, 32'h442f650f},
  {32'h453d073a, 32'hc1eeb0f4, 32'h441e27dd},
  {32'hc5046ec2, 32'h43d303c0, 32'hc4191639},
  {32'h45129365, 32'h432aad39, 32'hc3890d44},
  {32'hc3fb2b1e, 32'hc5283317, 32'h432f53ab},
  {32'h447a040e, 32'h44e46bcf, 32'h431209d2},
  {32'hc536f633, 32'h43514889, 32'hc3b42321},
  {32'h446c8995, 32'h44aad955, 32'hc4296261},
  {32'hc42fcc90, 32'hc4f088ee, 32'h432292a3},
  {32'h43d7aafc, 32'h44cc71a0, 32'h4360ab9f},
  {32'hc3e1f003, 32'hc3f38d7a, 32'h436a5c4f},
  {32'hc3b7d809, 32'hc423221a, 32'hc3f37f53},
  {32'hc3ab73d4, 32'hc4f7920a, 32'h449cb00c},
  {32'h43736b28, 32'hc39111a5, 32'hc46df67a},
  {32'h453bfac5, 32'h443c0a33, 32'hc3c7c2e2},
  {32'hc55ecd60, 32'h411b4b23, 32'hc16b2cc2},
  {32'hc2b97b28, 32'h42f64463, 32'h44b8a985},
  {32'hc40d78cb, 32'hc5082413, 32'hc4e73b5b},
  {32'h449c6e4f, 32'h440beb6e, 32'h44aafe63},
  {32'h437cd410, 32'h440fa83b, 32'hc409ba4a},
  {32'hc3997b20, 32'hc51c116d, 32'h45071c39},
  {32'hc3510f4f, 32'h449bf710, 32'hc49fef97},
  {32'h447ef3cc, 32'h43317125, 32'h443104c3},
  {32'hc46da297, 32'hc3f4bb17, 32'hc4730757},
  {32'h44f5d141, 32'h44098eda, 32'hc40e5699},
  {32'hc33b3e74, 32'hc48777ea, 32'hc4bb1d26},
  {32'hc22d53d4, 32'h447555c8, 32'h455fcde0},
  {32'hc2e35334, 32'hc3b9be88, 32'hc5673cd0},
  {32'h4443713d, 32'h44627c08, 32'h438f4d65},
  {32'hc4830a01, 32'hc49b8327, 32'hc40673ed},
  {32'h448375da, 32'h4500aa07, 32'h42e51d14},
  {32'h44551b66, 32'hc47517bd, 32'hc3c2ece8},
  {32'h44dec365, 32'h43721216, 32'h43cfe43a},
  {32'hc4a325dc, 32'hc4392fe3, 32'h42b6a3fd},
  {32'h44fccb3b, 32'h42e139ef, 32'h43a15635},
  {32'hc4b77d88, 32'hc40c2a60, 32'h4386fc8c},
  {32'h45864edc, 32'hc3fe1fcf, 32'h40be1a34},
  {32'hc3bed964, 32'hc48e826b, 32'hc40d350f},
  {32'hc48f528b, 32'hc2c49d07, 32'h44a7dd47},
  {32'hc2810982, 32'h43c62b11, 32'hc48a2fb9},
  {32'hc4f09006, 32'h43d797ef, 32'h436fd1ec},
  {32'h44940587, 32'hc358a4ba, 32'hc3e3fb40},
  {32'hc501ed6e, 32'h43972271, 32'h43edaa51},
  {32'hc3d89605, 32'hc44d9455, 32'hc4d3c56c},
  {32'hc4ff052d, 32'h41dc5c69, 32'h4461d8c0},
  {32'h44d3494a, 32'hc3dcbd30, 32'h439c2a1a},
  {32'hc4222e7e, 32'hc38ce79f, 32'h43e6d93b},
  {32'hc353b3d1, 32'h43cec6f0, 32'hc5167c85},
  {32'h43c2028b, 32'h4512a6d3, 32'h4337e764},
  {32'hc2970858, 32'hc4ebe6af, 32'hc38313b0},
  {32'hc43985a4, 32'h453f23a1, 32'h437a9d82},
  {32'h438ec65a, 32'hc3d7e25d, 32'hc3e4f151},
  {32'hc3de08f8, 32'h445577b0, 32'h44fd43af},
  {32'h43478560, 32'hc5104062, 32'hc4d4f579},
  {32'hc4a6c4d1, 32'h4426190a, 32'h434b96be},
  {32'h4334fe8c, 32'hc4c50992, 32'h43b5176f},
  {32'hc4f167bc, 32'h45081444, 32'h42ed8f6e},
  {32'hc4c5dde1, 32'h43986a27, 32'hc29a4825},
  {32'hc433b502, 32'hc2bedc33, 32'h44642714},
  {32'h44928853, 32'hc42fdb84, 32'h41b4f0d0},
  {32'hc4dd4c20, 32'h43952b52, 32'hc251d252},
  {32'h445809a0, 32'h43825baa, 32'h43fca0d1},
  {32'hc43b4b81, 32'hc328566c, 32'hc34d44c8},
  {32'h44c7ce53, 32'hc3df4baa, 32'hc323d2da},
  {32'hc406dd12, 32'hc3631ff1, 32'h444d0dda},
  {32'hc2f31c64, 32'hc26a682d, 32'hc53b92a1},
  {32'hc3522eb4, 32'hc32266cb, 32'h45121fc1},
  {32'h44834ba2, 32'h4441e172, 32'h434f0710},
  {32'h452d8d70, 32'hc415f6a2, 32'h42d5193b},
  {32'hc2dcfda2, 32'h45442d35, 32'hc24ee51c},
  {32'hc4bab2b9, 32'hc3ba518f, 32'h431aae19},
  {32'hc56548de, 32'h4426aba0, 32'hc3399ba2},
  {32'h446e8334, 32'hc4ab667a, 32'hc2939670},
  {32'h43e235c8, 32'h43c6fdfc, 32'h43bdcf26},
  {32'h449b9b1a, 32'hc0269e85, 32'hc42bde3b},
  {32'hc5130b2d, 32'hc216444b, 32'hc3be8ad5},
  {32'hc494abe2, 32'hc232cb5e, 32'h423384cc},
  {32'hc4ce503d, 32'h42f9dca6, 32'hc3f20c13},
  {32'hc1a25a94, 32'hc401fd72, 32'hc536c612},
  {32'h4414d191, 32'h448729cc, 32'hc3b4b2b8},
  {32'h431efed1, 32'hc475e568, 32'hc40a1ebd},
  {32'hc4eadc46, 32'h436fb6ad, 32'h447b4aac},
  {32'h43b208e2, 32'h44583195, 32'hc47327ee},
  {32'hc566ff94, 32'h43ddd2b3, 32'h4400aaaf},
  {32'h44ebdee5, 32'h44783502, 32'hc40293c1},
  {32'h42f646e0, 32'h4224d113, 32'h44bbf9d0},
  {32'hc1ada7fe, 32'hc4fde837, 32'hc4a36e91},
  {32'hc512a0cb, 32'h4394fa73, 32'h445ef952},
  {32'h43b02438, 32'hc3b747a3, 32'hc40cf026},
  {32'h42f48d50, 32'h4526e660, 32'h4404975e},
  {32'h440b6d72, 32'hc4d32326, 32'hc3abbd32},
  {32'h44f4dca4, 32'hc29214c9, 32'hc412e2ea},
  {32'hc51470ab, 32'hc35ee591, 32'h43ff660f},
  {32'h44c9c87c, 32'h43d1feb9, 32'h4409a2bf},
  {32'hc56847e1, 32'hc32cc1cc, 32'hc428854b},
  {32'h44905b89, 32'h446b1f00, 32'h42629304},
  {32'h43cafbd9, 32'hc25c8ee2, 32'hc3a501dc},
  {32'h43c2e660, 32'h45218b63, 32'h43081543},
  {32'hc52d5a6a, 32'hc3e9cade, 32'hc1ab0cd7},
  {32'h4452a842, 32'hc23f91f2, 32'h42cbefc4},
  {32'hc48bbba6, 32'h44009f3b, 32'h43ddac10},
  {32'h43c1c2bd, 32'h439b4a5c, 32'hc5058cc3},
  {32'h44bfe5fd, 32'h43f3fc66, 32'hc3970237},
  {32'h4541843d, 32'h43ba933f, 32'h42bfae2d},
  {32'h413b7b80, 32'hc4dd7280, 32'hc48d0a38},
  {32'h450c13c6, 32'h438cb747, 32'h434def07},
  {32'hc486a7e0, 32'h42bb9102, 32'hc4eb46a4},
  {32'h449b49ce, 32'h4409e5a5, 32'h4496a3c8},
  {32'hc44ec4f4, 32'hc42a2c76, 32'hc3438c66},
  {32'h45491c98, 32'hc3a80003, 32'h43674fbc},
  {32'hc57bfb65, 32'h431013f6, 32'h43340842},
  {32'h444a699d, 32'h4481d3c6, 32'h4397c418},
  {32'hc4471848, 32'hc4125a30, 32'hc3b2c4ac},
  {32'h441ca104, 32'h44ba9141, 32'h43fc0879},
  {32'hc455597e, 32'hc42c0298, 32'hc3dcf090},
  {32'hc39d2b28, 32'h4563e43a, 32'h4396e655},
  {32'hc3cd2f55, 32'hc4319640, 32'hc526d580},
  {32'h438bd6e0, 32'h446363b3, 32'h4400bfd8},
  {32'h44a94b6b, 32'h42390686, 32'hc3fb45e1},
  {32'h4329e9a0, 32'hc507854a, 32'hc2c50b10},
  {32'h44d81ced, 32'h437bf24e, 32'h449002c9},
  {32'hc5278aa7, 32'h4389e6fd, 32'h435e279f},
  {32'h4331829b, 32'h458ad771, 32'hc0b99988},
  {32'hc3f426c8, 32'hc4a1fb34, 32'hc1cf0db8},
  {32'h450ccb91, 32'hc2917420, 32'hc3d33bc5},
  {32'hc56fac5d, 32'h43a8cc5c, 32'h42283fc9},
  {32'h45409a52, 32'h4232505b, 32'hc1d22277},
  {32'hc39b7d7b, 32'hc3ba9621, 32'h42e44e23},
  {32'h43860d78, 32'h4478d1c4, 32'h42c70394},
  {32'hc37d1b06, 32'hc4d81fca, 32'hc108b783},
  {32'h43fc03bd, 32'h44e16206, 32'h43162f93},
  {32'hc50e8cc4, 32'h439a95de, 32'hc297b953},
  {32'h43ebcc46, 32'h4362c678, 32'hc4d7cb97},
  {32'hc48d6fac, 32'h4338a54f, 32'hc400113b},
  {32'h45206497, 32'h44162c26, 32'hc16b6406},
  {32'hc4436fa8, 32'hc2c328ce, 32'h44f07d6f},
  {32'h4459cdd9, 32'h43328674, 32'hc3ef1af1},
  {32'hc4ae147b, 32'hc3c41b37, 32'h444a5198},
  {32'h439a8cb0, 32'h4474c64e, 32'hc5052dec},
  {32'h43c1a64a, 32'h40476b94, 32'hc324be85},
  {32'h43c6adee, 32'h451ac612, 32'hc3347e6d},
  {32'hc38c1291, 32'h43bc587f, 32'h450693bc},
  {32'hc2c25070, 32'h438de8fd, 32'hc377a345},
  {32'hc50696a0, 32'hbfc4d128, 32'h43b332bb},
  {32'h43c867ca, 32'hc24f1bb9, 32'hc45b4c9a},
  {32'h4336b588, 32'hc4a84d9d, 32'hc3dc84c5},
  {32'hc53e05cc, 32'hc231c924, 32'hc2b8627f},
  {32'hc4639d22, 32'h43b8d12c, 32'h4189d582},
  {32'hc37093ec, 32'h4544639e, 32'h4323a0fb},
  {32'h4546a9ec, 32'h433f2815, 32'h42258297},
  {32'hc3470508, 32'h430071a2, 32'hc402960e},
  {32'h44e19de6, 32'h43d93082, 32'h41b6c214},
  {32'hc563df01, 32'h43ae1d56, 32'hc3005348},
  {32'h453ca66c, 32'hc2931807, 32'h43e3c4f0},
  {32'hc387191d, 32'hc37b9dd2, 32'h4437466d},
  {32'h4522c4e6, 32'h42921fd1, 32'h43f8fb11},
  {32'hc4bfbaa0, 32'h43a3da03, 32'hc307e164},
  {32'h4337ce50, 32'hc42cc527, 32'h4420e1ae},
  {32'hc54c106d, 32'h428aeccb, 32'h4315a1a2},
  {32'h43956dcb, 32'hc4a0686f, 32'h43cb3d55},
  {32'hc485e008, 32'h44c45bb4, 32'h4454b87a},
  {32'h445d5172, 32'hc3ac00d7, 32'h448f4c0f},
  {32'h44d05289, 32'h4224288d, 32'hc41e94af},
  {32'hc2b50e28, 32'hc52aa75d, 32'hc3aca2d7},
  {32'hc556cc9c, 32'hc3666fd7, 32'hc2ebf390},
  {32'hc34d6e9e, 32'hc3c0dec6, 32'h420edd6f},
  {32'hc4a30767, 32'h44256458, 32'hc4839efc},
  {32'h448bf514, 32'hc41677aa, 32'h43fd8dd1},
  {32'h4488c0ed, 32'hc397d1b1, 32'hc4ae0b8e},
  {32'h42dc1f91, 32'h43c120c6, 32'h45546a55},
  {32'hc52c86e6, 32'h4355bdcf, 32'hc43fb86f},
  {32'h4361c130, 32'h43f4c8a4, 32'h44156ae4},
  {32'hc3189a38, 32'h44aa9b58, 32'hc4c8a61d},
  {32'h442cb489, 32'h44b93b1c, 32'h44a930fe},
  {32'hc2f2e87e, 32'h43de9007, 32'hc3ee0103},
  {32'hc516241b, 32'h4380bf94, 32'h4319eec0},
  {32'h44f6ee9a, 32'hc36a6f7d, 32'h441fc30d},
  {32'hc4ae7f54, 32'hc314e49d, 32'hc3ff24f1},
  {32'h4468c13a, 32'h41700df6, 32'h43efb31d},
  {32'hc304aa64, 32'h44163786, 32'hc4d0228e},
  {32'h448898a1, 32'hc4864c99, 32'h43a04098},
  {32'hc43222a2, 32'h44b34f1e, 32'h451e57ee},
  {32'h43d2d340, 32'h44e8b2dc, 32'hc50724fa},
  {32'h44e6dcf6, 32'hc377c76e, 32'h42161478},
  {32'hc43dd1bf, 32'h43316e14, 32'h4472ff81},
  {32'hc30fbd90, 32'h42f3ea86, 32'hc4a87c9a},
  {32'hc40c6474, 32'hc3d20b6a, 32'h44580a58},
  {32'h4281efe8, 32'h436a987c, 32'h43210701},
  {32'h43d89f84, 32'hc40b5539, 32'h44b60bc2},
  {32'hc5021d29, 32'h3e894eb1, 32'hc4077b34},
  {32'h4553e774, 32'hc34fa531, 32'h431b2056},
  {32'hc5484965, 32'hc39f83c4, 32'hc411a90e},
  {32'h451f680d, 32'hc2e3ec53, 32'h443e49de},
  {32'h4485df1e, 32'hc3881473, 32'hc2bcb31b},
  {32'h451c295c, 32'hc4053c1d, 32'h441f79a2},
  {32'hc4c89968, 32'h44aa3dce, 32'h43b3dc50},
  {32'h4343d637, 32'hc498a742, 32'hc324f99f},
  {32'hc4cce8a6, 32'h44e5aaea, 32'h4369e0b2},
  {32'h44266358, 32'hc4303c1a, 32'h44231283},
  {32'h43a8b133, 32'hc424d655, 32'h4483de92},
  {32'h4518e460, 32'hc264a17f, 32'hc3d6f3df},
  {32'h438acf3e, 32'h444bca6a, 32'h4537b6f6},
  {32'hc532477a, 32'h439a48db, 32'hc2352368},
  {32'h4438087f, 32'h4490e952, 32'hc3280b31},
  {32'hc3cae642, 32'hc4039293, 32'h438568b3},
  {32'h4414b3d6, 32'h436f650a, 32'hc4e7c13f},
  {32'hc3f4ad10, 32'h42d5b4fd, 32'h4510d28f},
  {32'h42b1e23d, 32'h44c129a7, 32'hc3a96e0c},
  {32'hc29a7596, 32'h44708934, 32'h429a5608},
  {32'hc3e07c6c, 32'h44dd076d, 32'h44cbd957},
  {32'h4427d22e, 32'hc3a1568c, 32'hc49243d8},
  {32'h43081634, 32'h4501fc51, 32'hc3536149},
  {32'hc3986a6a, 32'hc463e6f4, 32'h4424f598},
  {32'h44e1fa80, 32'h43879736, 32'hc37db386},
  {32'hc2cf2d3e, 32'h43ce4aba, 32'h4560f50f},
  {32'h447c2933, 32'h442f93ed, 32'hc3ad7543},
  {32'hc42a6c5a, 32'hc429bd67, 32'h419a3fec},
  {32'hc380a650, 32'hc400af2b, 32'hc3dd831c},
  {32'hc4e2ce72, 32'h433afe38, 32'h4391c307},
  {32'hc45cd1a8, 32'hc276e91b, 32'h42cd204c},
  {32'h4325a448, 32'hc5200ca3, 32'hc34f260c},
  {32'h4429cd60, 32'h44d77399, 32'hc3502e68},
  {32'hbf169c00, 32'hc4da8eef, 32'h43bea125},
  {32'h440d8bef, 32'h44f47317, 32'hc416cdff},
  {32'hc4aa128c, 32'hc4841524, 32'hc3154f17},
  {32'hc38899c6, 32'hc2e833ae, 32'hc372af72},
  {32'h445a2954, 32'hc2e6381a, 32'h43dcd07e},
  {32'hc3e65944, 32'hc3872388, 32'hc41e774a},
  {32'hc3b0a727, 32'hc38ec668, 32'h44b0daea},
  {32'h42365485, 32'h43616b23, 32'hc4cbe652},
  {32'h44ce6fe5, 32'h4465789a, 32'h4330f5f8},
  {32'hc253b17e, 32'h43948ae4, 32'hc40e7152},
  {32'h44394f26, 32'hc31cad04, 32'h44080c21},
  {32'hc3c07106, 32'hc3be67f1, 32'hc56329ef},
  {32'hc31ea7a4, 32'h44af9692, 32'h4507dbe0},
  {32'h437a6d4e, 32'hc3e2a999, 32'hc3e49b58},
  {32'hc3ebfad3, 32'hc468bd34, 32'h44a77437},
  {32'hc43e6c1c, 32'h41cde406, 32'h42d298ee},
  {32'h44bf5bb4, 32'h44059fdb, 32'hc258549f},
  {32'hc41eecdb, 32'hc37a0693, 32'hc4c8d59b},
  {32'h44c64b0f, 32'h442e4899, 32'h43e02ad3},
  {32'hc2204488, 32'hc4906427, 32'hc341f137},
  {32'h4546f446, 32'hc335bff8, 32'hc31da915},
  {32'h432590e5, 32'hc20f8a38, 32'hc5525c92},
  {32'h4474fd27, 32'h4449c444, 32'h43fc2836},
  {32'hc3282256, 32'hc535a703, 32'hc3a9637f},
  {32'hc352bfb0, 32'h454932dd, 32'h42745f46},
  {32'h445ab872, 32'hc3b0a265, 32'hc359099c},
  {32'h4435e340, 32'h44d53389, 32'hc4072345},
  {32'hc40f303f, 32'hc36e22d8, 32'h42c49e17},
  {32'h454a50a9, 32'h4410cf90, 32'h43bddc1c},
  {32'hc50817eb, 32'hc3ba4613, 32'hc4438e5e},
  {32'h454a2ece, 32'hc1fddd66, 32'h43a18bf6},
  {32'h43093398, 32'hc4ccb022, 32'hc3bf3a53},
  {32'hc46ee383, 32'hc43d18a2, 32'h44bb256a},
  {32'h43a341f3, 32'hc2fa7410, 32'hc22a8ac2},
  {32'hc3585700, 32'h4403e525, 32'h44c257c8},
  {32'hc4162cfa, 32'hc520a734, 32'hc3ba9d69},
  {32'hc3cc769b, 32'h43abf328, 32'h44f3252a},
  {32'h43daefb9, 32'hc447e18c, 32'hc4d89f16},
  {32'hc4314442, 32'h44367750, 32'h4510b526},
  {32'h447208c5, 32'hc4216286, 32'hc427033b},
  {32'hc41fe407, 32'hc1c0677a, 32'h44334e30},
  {32'h43a6d4d0, 32'hc39506c8, 32'hc488b306},
  {32'hc498d5b0, 32'h431cf6fe, 32'h4364b256},
  {32'h44fa9b0a, 32'h4365c6f7, 32'hc38f3887},
  {32'hc420e6f6, 32'h4432f818, 32'h446387cc},
  {32'hc35658df, 32'hc4b4f52f, 32'hc366fa87},
  {32'hc380c888, 32'h44ec922f, 32'h44e67524},
  {32'hc34eae48, 32'hc443a629, 32'hc513a33f},
  {32'hc42015da, 32'h44baaa9c, 32'h43969b7e},
  {32'h44b03fc4, 32'hc48e716c, 32'hc33565cd},
  {32'hc49bc4c6, 32'h44589de4, 32'h4291a70a},
  {32'hc49edc4f, 32'h4392e3a4, 32'h436efe47},
  {32'h42f698ac, 32'h4225f0a9, 32'h429e6cbb},
  {32'h4152e000, 32'hc54f7a6f, 32'hc379fa20},
  {32'h420b5260, 32'h44a3fde0, 32'h42f2be42},
  {32'h44de4c17, 32'h435d0e89, 32'hc2c42427},
  {32'hc4adf0fa, 32'h43d30323, 32'h42eb545f},
  {32'h452ea490, 32'hc2238995, 32'hc2900ce1},
  {32'hc33fab4e, 32'hc38e469a, 32'hc3278a31},
  {32'hc523efb3, 32'h42d551da, 32'hc2183e1c},
  {32'h430cc85c, 32'hc310f5cc, 32'h44211ec5},
  {32'hc4fcb852, 32'hc3957125, 32'h43484967},
  {32'h44cc7859, 32'h43445bc0, 32'hc37896c3},
  {32'hc465ef48, 32'h4507eba6, 32'h43008008},
  {32'h444195b5, 32'hc42b6e07, 32'hc3937f4a},
  {32'hc5365a2d, 32'h41edec18, 32'h43765c82},
  {32'h43f56232, 32'hc518dfee, 32'hc331efb7},
  {32'hc52637b7, 32'hc3b48069, 32'h4326cdc9},
  {32'h4533552c, 32'h4342a0e0, 32'h434b644b},
  {32'hc41c995e, 32'h4498781e, 32'h449b704d},
  {32'hc3cddc22, 32'h4211bd14, 32'hc27045b0},
  {32'hc4c82086, 32'hc243542e, 32'h4413e19d},
  {32'h431ce557, 32'hc42bd650, 32'hc5540393},
  {32'hc53b8e4b, 32'h4358b391, 32'h4325bf90},
  {32'hc38f6158, 32'hc34e96d0, 32'hc50e4cec},
  {32'hc506be11, 32'hc38fd600, 32'h4405558b},
  {32'h4534f94e, 32'h43f90ffc, 32'hc434a98e},
  {32'hc5086696, 32'hc44e30af, 32'hc31abc68},
  {32'h43a88838, 32'h4423ad6e, 32'hc4a8a572},
  {32'h445d26f0, 32'h43ed33ac, 32'hc2d46b0c},
  {32'h448c8322, 32'hc469000c, 32'hc2a78b3d},
  {32'hc404f9de, 32'hc34c754d, 32'h45617504},
  {32'h451eb80a, 32'hc3ce05c4, 32'hc3228a18},
  {32'hc0492300, 32'h448d0ab0, 32'h44fcf215},
  {32'h4278b8c8, 32'hc41f0a0c, 32'hc50959df},
  {32'h44522fc3, 32'h431072da, 32'hc4873b24},
  {32'hc4e126c9, 32'h437c3b30, 32'h44f3e340},
  {32'hc290f052, 32'h43b55ea4, 32'hc17312d2},
  {32'hc52704c7, 32'hc41edfc5, 32'h43001400},
  {32'hc20554c0, 32'h42b7d26b, 32'hc42a933c},
  {32'h433969b2, 32'hc4c56afa, 32'hc3353420},
  {32'h430a4ab0, 32'h45373e2d, 32'h43d7d9ff},
  {32'hc4da15ac, 32'hc4c4198f, 32'hc42e1543},
  {32'hc47593b7, 32'h43e76029, 32'h43c4d4df},
  {32'hc52175f7, 32'h42fe2e91, 32'hc265a5f4},
  {32'h44e81da9, 32'h42066a2d, 32'hc4860850},
  {32'h438dfd72, 32'h4306a662, 32'h43836cf5},
  {32'h435e8c1c, 32'h4388d7cc, 32'h452fc126},
  {32'hc3543dc0, 32'hc553f4d2, 32'hc21cf3f6},
  {32'hc4d24179, 32'h42d47452, 32'h439259fa},
  {32'hc4c5994d, 32'hc3e41106, 32'h4318d6f2},
  {32'h450f2ee6, 32'h44066e77, 32'h43a7ac4c},
  {32'hc47bf66d, 32'hc4ac1437, 32'h431d75c4},
  {32'h4342bfc0, 32'hc38e4459, 32'h44180000},
  {32'hc4c62448, 32'h4354ca58, 32'h430d93e8},
  {32'h455748ad, 32'h4387adb3, 32'hc31c1c98},
  {32'hc497de65, 32'hc308f714, 32'hc4e89e53},
  {32'hc2b1e147, 32'h4517bcd2, 32'h436074c1},
  {32'h40e47b30, 32'hc4b538b9, 32'hc3c0d3a9},
  {32'h450da921, 32'h445896ce, 32'h43afacda},
  {32'hc5253cb9, 32'hc3a4181b, 32'hc24a288d},
  {32'hc3c015a6, 32'h44171816, 32'h43fdde22},
  {32'hc18d5852, 32'h450cd0ea, 32'hc3cf210b},
  {32'hc5604eaa, 32'hc25fa200, 32'h435a319d},
  {32'h43a3a8e8, 32'h4493f065, 32'h43050a4a},
  {32'hc38505c7, 32'hc47ecd5e, 32'h42a46835},
  {32'h4355482e, 32'h4513134b, 32'h4141e79d},
  {32'hc53ea382, 32'hc4086cbf, 32'h43c6c662},
  {32'h44d8bcd4, 32'h4377c8e5, 32'hc40433e8},
  {32'hc54ea461, 32'h4342a944, 32'hc406f2e8},
  {32'hc30d6c60, 32'hc3af532c, 32'h4404fa5d},
  {32'hc49c08eb, 32'h43d1c694, 32'hc346b149},
  {32'h438a3a38, 32'h44696043, 32'hc4b914d5},
  {32'h4338657c, 32'hc52ea51c, 32'hc347c276},
  {32'h4337daeb, 32'h44042adc, 32'hc4a05090},
  {32'hc49a2b5a, 32'hc412ec82, 32'h44078544},
  {32'h444003ca, 32'h4340ca9e, 32'hc4be3e15},
  {32'hc4d9332e, 32'hc3e5a07c, 32'hc19267ec},
  {32'h428d1b68, 32'h44c38f38, 32'h44ae624d},
  {32'hc4c34dfe, 32'hc3a83d3e, 32'hc307747e},
  {32'h44a78ca8, 32'h43b63edd, 32'hc3119b13},
  {32'hc3060c46, 32'hc4b994b4, 32'h4317aae4},
  {32'h4552af4b, 32'h440adde3, 32'hc3c7dd4a},
  {32'hc46e4525, 32'hc4297351, 32'h43182ce2},
  {32'h4533673b, 32'h4387e17a, 32'h439519c3},
  {32'h43072e80, 32'h435cb3f1, 32'h44a46970},
  {32'h4556bb05, 32'h44291697, 32'hc2dfd516},
  {32'h42e9b470, 32'h44a5b37c, 32'h4522bef9},
  {32'h44db8123, 32'hc418572e, 32'hc48fd1a4},
  {32'h438b8eb4, 32'hc4731a9e, 32'hc2a66667},
  {32'hc3dc0150, 32'h4546f1e3, 32'h4413a44c},
  {32'hc460cb38, 32'h4312fb5f, 32'hc39577f2},
  {32'hc33e23dc, 32'h44203798, 32'hc34381a7},
  {32'h43b3e3f0, 32'hc55db428, 32'h43922679},
  {32'h44374aae, 32'h4379ae86, 32'hc342f61a},
  {32'h451eb683, 32'h4421b1de, 32'h43956afb},
  {32'hc48b7822, 32'h438abe9a, 32'h40180e7e},
  {32'hc488af23, 32'hc34f14ed, 32'h43e271d8},
  {32'hc28e23d8, 32'h4345e36e, 32'h43e8cea4},
  {32'h43c3e40e, 32'hc5047356, 32'hc1207c9a},
  {32'hc33fcd14, 32'hc2e2ddbb, 32'h4275d97e},
  {32'hc389e626, 32'hc5162991, 32'h43f878dc},
  {32'hc512f6fd, 32'h4416e82b, 32'hc2a29618},
  {32'hc4517928, 32'hc3b0d943, 32'hc343f04b},
  {32'hc4bad03e, 32'hc3644976, 32'hc49a1036},
  {32'h43a718a0, 32'h43b8e606, 32'h44a45f40},
  {32'hc50de720, 32'h44118663, 32'hc1da969d},
  {32'h42be6ae8, 32'hc437fc0f, 32'h43ba261e},
  {32'hc397ccf9, 32'h44893276, 32'hc4b8829c},
  {32'hc41edf4a, 32'hc462a357, 32'hc2ab78b6},
  {32'hc4663725, 32'h43926fb2, 32'hc4f8d3a8},
  {32'hc3848d86, 32'hc46d0fea, 32'h44d07d7e},
  {32'h441c9e2a, 32'hc33942e2, 32'hc302ee67},
  {32'h44f343c2, 32'hc2b991a0, 32'h4479756c},
  {32'hc4181828, 32'hc43670d5, 32'hc3c346c3},
  {32'h444e3211, 32'h442ecf6c, 32'h443fbc73},
  {32'h41127908, 32'h42932a9e, 32'hc4cc60fe},
  {32'h45007275, 32'h43d3f805, 32'h43d1e8e8},
  {32'h43a7fe0b, 32'hc46137fa, 32'hc49d9fb6},
  {32'h449d74a5, 32'h4390ee30, 32'hc3804dd8},
  {32'h4419ba1a, 32'hc47767d8, 32'h44e99358},
  {32'hc337c815, 32'h455c7f31, 32'h440ec7f1},
  {32'h4397f6cc, 32'hc4a20ce8, 32'hc3155a15},
  {32'hc43af588, 32'h449eb0cc, 32'hc3b94634},
  {32'h4489e902, 32'hc1f243d4, 32'h44ac5bc1},
  {32'hc291e3cb, 32'h45006854, 32'h44c2b88a},
  {32'h4212e958, 32'h4425482b, 32'hc50a8e1a},
  {32'hc44a9c00, 32'h438faa04, 32'h448fd556},
  {32'h440eccfe, 32'hc35fb81c, 32'hc31441ee},
  {32'hc508f259, 32'h439e8030, 32'hc2c1e3d0},
  {32'h442a0d4a, 32'hc20ff341, 32'h44c1e69e},
  {32'hc401f356, 32'h444ee3f9, 32'h43b135ff},
  {32'h444de5f4, 32'h4385ecbf, 32'h4400fc9c},
  {32'h4403df2d, 32'h4516d8f3, 32'hc42aa3f2},
  {32'h4249c250, 32'hc4680f32, 32'hc0cb875c},
  {32'hc37fd0b0, 32'hc383630b, 32'hc3ff4cf2},
  {32'h44e7f4f0, 32'h433214d6, 32'h433acc02},
  {32'h43a2f120, 32'hc356a4af, 32'h41dde381},
  {32'h451a8e63, 32'hc3fb729c, 32'hc38d294b},
  {32'hc4580558, 32'h438a0808, 32'h43796a33},
  {32'h45126de4, 32'h438f6e34, 32'h43aa0771},
  {32'hc533f0fe, 32'h43ede3b8, 32'h42494c07},
  {32'h45013039, 32'hc4be0f3d, 32'hc355dc12},
  {32'h43d1c8ca, 32'h442921e1, 32'h43987d9a},
  {32'hc404ae1b, 32'hc42cd29d, 32'hc5348b8e},
  {32'hc43b50b2, 32'hc4cb4be8, 32'h44b639c6},
  {32'h43d1e49e, 32'hc4489f09, 32'h44d495a6},
  {32'h430bd19a, 32'h43861a73, 32'hc4b74b98},
  {32'h44c7ef97, 32'h4389ed39, 32'h4392cd94},
  {32'h4421e436, 32'h43d41fff, 32'hc49fa412},
  {32'hc508c5fa, 32'hc4317bc9, 32'h4382d6a7},
  {32'h451ca910, 32'hc251de9e, 32'h44154777},
  {32'hc3574c5b, 32'hc42ba9bb, 32'hc47a9d44},
  {32'hc4b4d107, 32'h43c8f977, 32'h449c1913},
  {32'hc29e57c0, 32'hc402d763, 32'hc4c64d0d},
  {32'h448d5207, 32'h442d6a3f, 32'hc3ec3fe0},
  {32'hc3cfa86a, 32'hc1d889e6, 32'h442870ac},
  {32'hc48a4520, 32'h43db6413, 32'hc3d24c75},
  {32'hc37770e8, 32'hc53585a9, 32'hc36852de},
  {32'h445956fb, 32'h43514227, 32'hc4593f96},
  {32'hc3f0895f, 32'hc33226d0, 32'h4351d44c},
  {32'h43e02ef0, 32'hc353c7f5, 32'hc40de748},
  {32'hc4b557e2, 32'hc3f85169, 32'hc1c2c374},
  {32'h45130b2f, 32'hc3274c8e, 32'hc38799b6},
  {32'hc50bb6a3, 32'hc42b6899, 32'h43ab4fb9},
  {32'h44f0ad4e, 32'h42d68542, 32'hc25753f3},
  {32'hc4a367fc, 32'hc3b35437, 32'h432ecedc},
  {32'h44d5ef68, 32'h44b0840e, 32'h43be0689},
  {32'hc55a561e, 32'hc3deb994, 32'hc3e60f90},
  {32'h451fcdda, 32'hc437b017, 32'hc26d202c},
  {32'hc38ded4d, 32'hc3b9bc84, 32'h43beb27f},
  {32'hc3e7d9d0, 32'h4421921b, 32'hc4852c63},
  {32'h43c23345, 32'h44bc5818, 32'hc3b17fee},
  {32'hc3d4e2b3, 32'hc34f9b47, 32'hc358f024},
  {32'h42f17054, 32'h44e91dc7, 32'h43e8361f},
  {32'hc436660d, 32'hc241fb6a, 32'hc4175cda},
  {32'h43923bab, 32'h43364b51, 32'h44811aa1},
  {32'hc53251d2, 32'hc384d948, 32'hc35ba6df},
  {32'h426c5750, 32'h44df3a40, 32'h44dfbb17},
  {32'h44166477, 32'hc206086a, 32'hc3fb5d57},
  {32'h44843366, 32'hc1eea3c3, 32'h4380feda},
  {32'h4148d130, 32'hc50c0616, 32'hc3ec8be1},
  {32'h4513d292, 32'hc2cb8729, 32'h439f6018},
  {32'hc4117dc0, 32'hc4f23a13, 32'hc39c25dd},
  {32'h443e3d52, 32'h449fcb83, 32'h4334e5ca},
  {32'h4403063f, 32'hc33c9c5d, 32'hc3bfdab1},
  {32'h44bfe8cd, 32'h42b6fb0a, 32'h42cbd530},
  {32'hc4938cbf, 32'hc44eb19b, 32'hc410f811},
  {32'hc50b9029, 32'h439993bc, 32'h42da0aad},
  {32'hc55897d2, 32'hc2cf5708, 32'hc38fee92},
  {32'h4531abcd, 32'h43a7a642, 32'h43a2fef1},
  {32'hc4a4d6fb, 32'hc37a474b, 32'hc273818d},
  {32'h44d2d6d7, 32'h43b15782, 32'hc2e41b69},
  {32'hc310ae60, 32'hc4d777fb, 32'hc371cc7e},
  {32'h4501e104, 32'hc119243c, 32'h43af70ed},
  {32'hc4a26d4c, 32'hc421de0a, 32'h438b35f6},
  {32'hc30e9ee0, 32'hc3c97f9e, 32'h43a25c48},
  {32'h43d4fbcc, 32'hc4b3e3ba, 32'hc490d4eb},
  {32'hc28715e0, 32'hc50e51b0, 32'h44ba184e},
  {32'h44728f16, 32'hc20e25fc, 32'hc2dd7487},
  {32'h40b5ab60, 32'h44fc2bc6, 32'h4471a0f0},
  {32'h43d1dee5, 32'hc4ff4908, 32'hc36ac212},
  {32'h42d46410, 32'hc296c857, 32'h44caf90a},
  {32'hc04a72a0, 32'hc4626771, 32'hc52cf25d},
  {32'hc4b5769b, 32'h43511615, 32'h446cb795},
  {32'hc423642d, 32'hc3d80c75, 32'hc46fe6f6},
  {32'hc4887a80, 32'h448c4d09, 32'h43a198ce},
  {32'hc403b53c, 32'hc53b2e05, 32'hc40b8029},
  {32'hc45972d6, 32'hc38d11fb, 32'h436909cf},
  {32'h43a23d25, 32'hc3bafa0c, 32'hc3ac0ebf},
  {32'hc53bb9c3, 32'h40f2f930, 32'h4369f20f},
  {32'h44d63de5, 32'h433eb9c9, 32'hc3df47ec},
  {32'hc4b8fc0c, 32'hc206a055, 32'h449d3c06},
  {32'h4515d714, 32'hc480154b, 32'hc2c3cb21},
  {32'hc4278fce, 32'h44bb1dcb, 32'h4395a1f4},
  {32'h452648a7, 32'hc49015a9, 32'h439a6ae6},
  {32'hc0d9b2c4, 32'h453c1958, 32'h43167e1f},
  {32'h44c3663d, 32'h43948917, 32'hc1b19acb},
  {32'hc4e07c83, 32'h45042fe7, 32'h43747aa2},
  {32'h444b44a9, 32'hc575ca72, 32'h43db23e6},
  {32'hc4af149d, 32'h4387a00b, 32'h430d964d},
  {32'h451c0a8a, 32'h434d6f4f, 32'h43ea6515},
  {32'hc51f2b23, 32'h43ad8a46, 32'h43f217cc},
  {32'hc380c02a, 32'hc2e94746, 32'h44083473},
  {32'h45296db6, 32'hc387f287, 32'hc38e7d2c},
  {32'hc3aae41d, 32'h443b1e38, 32'hc50f4b23},
  {32'h451a0042, 32'hc401fdbf, 32'h44435b7b},
  {32'h440b2fe9, 32'h43847653, 32'hc3b5eca1},
  {32'h4500a7ce, 32'hc3e43dd6, 32'h4397a9a3},
  {32'hc409473c, 32'h443db052, 32'h43e1cb9a},
  {32'hc4d7094d, 32'hc3345c30, 32'hc3817f36},
  {32'hc567c21e, 32'h4418b4b8, 32'hc31ebccf},
  {32'h44f99617, 32'hc41d928e, 32'h4143f094},
  {32'hc461a81b, 32'h40a4eee1, 32'hc3f00c7b},
  {32'h440216f4, 32'h430a6203, 32'hc1891003},
  {32'hc4404a4a, 32'hc35d5fb4, 32'hc4d9949b},
  {32'h4423f5f4, 32'hc31e872b, 32'hc44d434c},
  {32'h4359014c, 32'h42cab29b, 32'h450ab19d},
  {32'h4387006c, 32'hc42e3803, 32'hc4cb9a3c},
  {32'h42e67a3c, 32'h45141818, 32'hc237b68f},
  {32'hc3c24392, 32'hc252b69a, 32'hc529ec00},
  {32'hc4290f86, 32'h4484bcde, 32'h4371eed0},
  {32'hc433277c, 32'hc3049fd6, 32'hc43292ed},
  {32'hc51fe2f6, 32'h4411cb91, 32'hc12eb633},
  {32'h44ea82d2, 32'hc438d92b, 32'hc442d509},
  {32'hc24a7b8c, 32'h437b43df, 32'h45024fd6},
  {32'hc40f68c7, 32'hc3bc265f, 32'hc4cc88f8},
  {32'hc306b03c, 32'h45453547, 32'h41e3d3aa},
  {32'hc416a101, 32'hc31173ad, 32'hc38003a0},
  {32'hc434fd36, 32'h437efc64, 32'h4463e0d5},
  {32'h4495bb04, 32'hc4cd4304, 32'hc3fb9f9d},
  {32'h43cf6db0, 32'hc423f9e8, 32'h4292e2e4},
  {32'hc3819112, 32'h436326a0, 32'h44db7968},
  {32'h439a225a, 32'h447d62b1, 32'hc422a810},
  {32'hc41473ca, 32'hc52a4ad8, 32'hc4100bc8},
  {32'h445e5aac, 32'hc2c4043a, 32'h42e83212},
  {32'h441cc576, 32'h42b2f2dd, 32'h42ce76b1},
  {32'h44448324, 32'h44ae7b21, 32'h43456312},
  {32'hc5064f06, 32'hc454f23f, 32'hc332caf6},
  {32'hc4cc6f73, 32'hc38f1691, 32'h43db9410},
  {32'hc4225ffe, 32'hc248aee3, 32'h44ab5bc7},
  {32'h44083f96, 32'h43d465cb, 32'hc43168f5},
  {32'hc3f64724, 32'hc12ff687, 32'h43a2957e},
  {32'h447d0120, 32'h4428ffdd, 32'h4491e713},
  {32'hc4201216, 32'hc3d99859, 32'hc3b76bce},
  {32'h438d2174, 32'h4399cac8, 32'h44803bac},
  {32'hc4c6be71, 32'hc3add67b, 32'hc16839f9},
  {32'h441163a7, 32'h440327ee, 32'h4413b7aa},
  {32'hc4ab4778, 32'h4099d86b, 32'hc385b8ea},
  {32'h43413350, 32'hc452601d, 32'h44c2fccd},
  {32'hc4ea754c, 32'hc40d9eae, 32'hc4b7aab2},
  {32'hc38d9357, 32'hc32d6dd5, 32'h434b62ce},
  {32'hc39e5300, 32'hc4f75b12, 32'hc25612a7},
  {32'h430e37ac, 32'h43e89152, 32'h44d796b3},
  {32'h4483a637, 32'hc438f7b3, 32'h429fe83a},
  {32'h43b65258, 32'h44e34c7f, 32'h4405e3c2},
  {32'hc0553600, 32'hc53d8820, 32'hc31fa8ce},
  {32'h440a0d8e, 32'hc396dfbe, 32'h446596b8},
  {32'hc2e53c9c, 32'h437ea1c8, 32'hc429c441},
  {32'hc49b3712, 32'hc37b20f7, 32'h435ce935},
  {32'h43ab577c, 32'h44b92690, 32'hc39495b1},
  {32'h448584f9, 32'hc4230127, 32'hc357223d},
  {32'h449a0901, 32'h44b2c7e4, 32'hc37cf00e},
  {32'hc449144a, 32'hc50a1033, 32'h420362c1},
  {32'hc4c04503, 32'h43b06251, 32'hc269eb45},
  {32'hc3dde81c, 32'h440d17ab, 32'h420fcb9d},
  {32'h44675130, 32'h44857346, 32'h448256cf},
  {32'hc4d1d1be, 32'hc1d6c43b, 32'h43b21d47},
  {32'hc18943a0, 32'h4498c701, 32'hc5069512},
  {32'hc51e557b, 32'hc2e892f2, 32'hc37b001e},
  {32'hc2e1a2a0, 32'hc26e262a, 32'hc4d12105},
  {32'hc45d1d3d, 32'hc3cc22ef, 32'h44530dd5},
  {32'h42b92ab4, 32'h451e355f, 32'hc420bf23},
  {32'h451003c9, 32'hc3011975, 32'h41b19eb3},
  {32'h4391b85b, 32'h421c395f, 32'hc48e911e},
  {32'hc3c99df4, 32'hc3b405da, 32'h4494aba1},
  {32'hc4ce2382, 32'h439f70ad, 32'hc39270e4},
  {32'hc3b6a9c0, 32'hc5070c59, 32'h4432112c},
  {32'h4506572e, 32'h449fb836, 32'hc42188e1},
  {32'hc4cb2107, 32'h41cd9606, 32'h431c467c},
  {32'h429eff90, 32'h44e07c5b, 32'hc43022da},
  {32'h4349c428, 32'hc4f7b8e7, 32'h4479e3fc},
  {32'h440e8a64, 32'h440cae1d, 32'hc394ad18},
  {32'hc5171018, 32'h43d57a41, 32'h43be7c02},
  {32'h445ac6a2, 32'hc3a46dda, 32'hc4a89d79},
  {32'h4482fb90, 32'hc42fcb1b, 32'hc44acf43},
  {32'hc4623f32, 32'h44fb74fb, 32'h43fb2f41},
  {32'h44ed4ae7, 32'h43398732, 32'h43fdcb95},
  {32'hc5262439, 32'h43439c38, 32'h4422d880},
  {32'h4518158e, 32'hc38e65e0, 32'h43ecffe0},
  {32'h449badad, 32'h438ebd43, 32'h438e3a07},
  {32'h4540c826, 32'h43865265, 32'h4265fa83},
  {32'hc50fff18, 32'h44121549, 32'h4434ab02},
  {32'h452afa50, 32'hc2fe89c2, 32'hc3265d99},
  {32'hc51daaf2, 32'h439525d1, 32'h4331bd16},
  {32'h435b5368, 32'h42655958, 32'hc3d4e072},
  {32'hc43a3f9d, 32'h4343f726, 32'hc3fce5b1},
  {32'h44b9034b, 32'hc33ba6d8, 32'h4376a4ec},
  {32'hc4238dc6, 32'h44d006cc, 32'h42e3a93b},
  {32'h4500be14, 32'h412a5838, 32'h437cee0e},
  {32'hc3293442, 32'hc3ed83ac, 32'hc54b7794},
  {32'h44f31076, 32'hc3e402c5, 32'h442dfe70},
  {32'hc50e86dc, 32'h43c5bfdd, 32'hc0ff246f},
  {32'h449a2abd, 32'hc45b548a, 32'h44245236},
  {32'hc533ad19, 32'h440266cc, 32'hc427afbd},
  {32'h44879a5a, 32'h432f7c76, 32'h432fbe97},
  {32'hc48154fa, 32'h44997fcd, 32'hc44089be},
  {32'h41b6bbca, 32'hc290815b, 32'h45207ee8},
  {32'h43ad322a, 32'h43e60795, 32'hc47937d7},
  {32'h4394d00a, 32'h447334d2, 32'h45168d3d},
  {32'hc4c2459a, 32'hc2ffbfa3, 32'hc50ce148},
  {32'hc4b24144, 32'hc3936eaf, 32'h437a17fe},
  {32'hc40c12b4, 32'hc5044f23, 32'hc4b4dadc},
  {32'h436b0dae, 32'hc4ffcbc4, 32'h45073b0a},
  {32'h420438d8, 32'h433d690d, 32'hc4960573},
  {32'hc4b27b32, 32'h43023b70, 32'hc2d5fabc},
  {32'hc1886080, 32'hc51b56c2, 32'h4409693e},
  {32'hc4b026d4, 32'h43d4c4a9, 32'hc3cd0098},
  {32'h44fc7f09, 32'h438aec54, 32'h43c37eee},
  {32'hc3c77474, 32'hc3251738, 32'hc55a2c8d},
  {32'hc45d26d4, 32'hc4c6de19, 32'h435508cc},
  {32'h42af9cec, 32'hc47263c9, 32'h450a0d13},
  {32'hc3f7e140, 32'h44eafe10, 32'hc4e2ed24},
  {32'hc4803afb, 32'h429003cb, 32'h43776472},
  {32'h425eed40, 32'hc4092b06, 32'h4457067a},
  {32'hc347c31c, 32'h43bcef71, 32'hc416232c},
  {32'h449f4edc, 32'hc3c2f068, 32'h4364d716},
  {32'hc2dad708, 32'h43490cbb, 32'hc4ef6c1c},
  {32'h44c10dc4, 32'hc4436ec3, 32'h43f7c6e8},
  {32'hc5003a0b, 32'h41c06222, 32'hc34bc622},
  {32'h44a68ed6, 32'hc41aeb96, 32'h4320b664},
  {32'hc47c0e1d, 32'hc42cc56c, 32'hc314828c},
  {32'h45761017, 32'h441b1efd, 32'hc35efceb},
  {32'h434cff2a, 32'h44929638, 32'hc2696a12},
  {32'h441e4cb7, 32'h438e754f, 32'h43c253bc},
  {32'hc4073044, 32'h45170abb, 32'hc3b4e8a9},
  {32'h41158e80, 32'hc3cec346, 32'h42eb109c},
  {32'hc527a5bd, 32'h44612ff7, 32'h4414c0ba},
  {32'h435660b0, 32'hc52f3f89, 32'hc3f32759},
  {32'h4485a994, 32'h444202b5, 32'h43bc8a6e},
  {32'hc2d92007, 32'h44216eaa, 32'hc5467e53},
  {32'hc38d33c7, 32'hc46fd06f, 32'h44541a17},
  {32'h42e5edf0, 32'hc4771c70, 32'h44b2bd63},
  {32'h455aaa87, 32'hc396cf4c, 32'hc2e62045},
  {32'hc2e0c6e0, 32'hc43b5332, 32'h3e89ea80},
  {32'hc13e94a6, 32'h453d5a45, 32'hc42496a9},
  {32'hc4e72325, 32'hc3f57c6b, 32'h4385510b},
  {32'h442abd88, 32'hc3accb39, 32'h432f46ed},
  {32'h4510afb8, 32'hc24467cc, 32'h43b10295},
  {32'h43033a5d, 32'h44d57f7a, 32'h45056032},
  {32'hc2f148e0, 32'h44b2659d, 32'hc4a32ec9},
  {32'h4435fa65, 32'h43917e59, 32'hc4a678a2},
  {32'hc3edf1d5, 32'hc452a5e5, 32'h44634a2f},
  {32'h4431b94d, 32'h431553d0, 32'hc4a8e9e1},
  {32'hc4814076, 32'hc48a7176, 32'h441642f0},
  {32'h436ac6cc, 32'hc458d9be, 32'hc515d7bf},
  {32'hc4ae4baa, 32'hc37f68cf, 32'hc42f51d6},
  {32'h450c1ca4, 32'hc39106cb, 32'hc2acbcc9},
  {32'hc5047ec8, 32'h425a255c, 32'h4445156e},
  {32'h43c781bc, 32'h43a78b78, 32'h4256a0a0},
  {32'hc4582a4c, 32'hc508556c, 32'hc376252c},
  {32'h43c94690, 32'h433d030e, 32'h42c5fa8c},
  {32'hc53b83a4, 32'h439281f9, 32'hc3cafbcb},
  {32'h43673ba4, 32'h4513367c, 32'h4406739f},
  {32'hc536a588, 32'hc3cbb1f2, 32'h43b8ee2d},
  {32'h4537a243, 32'hc3a3775d, 32'h43a5b8a7},
  {32'hc3dd57a8, 32'hc3bd11d0, 32'h4354363f},
  {32'hc21e558e, 32'hc35002a0, 32'hc4279af4},
  {32'h444d6efe, 32'hc3e0f030, 32'h435f5f92},
  {32'h4349db02, 32'h419aab47, 32'hc4c7b01e},
  {32'h4507ad2b, 32'h4218ffca, 32'h435d070e},
  {32'hc42dda40, 32'hc43361a5, 32'hc3d323f5},
  {32'h44167762, 32'h428230b0, 32'h44c5695f},
  {32'hc3e71ca4, 32'hc42bd2be, 32'hc531db63},
  {32'h441b42c1, 32'h446da456, 32'h44ed3c42},
  {32'hc3c7d105, 32'hc4574b6a, 32'h42ba88b0},
  {32'hc41908be, 32'hc2cadf61, 32'h45026bf5},
  {32'hc3516f8d, 32'hc4a49334, 32'hc4289b10},
  {32'h43c4bdea, 32'h445f5af5, 32'h43a527ac},
  {32'hc41ba764, 32'hc3fa101e, 32'hc4dd6535},
  {32'h445a5ed2, 32'hc2565e30, 32'h4362330c},
  {32'h4410bda8, 32'hc1bc034d, 32'hc41be91c},
  {32'hc4131435, 32'h445d57ce, 32'h451c5c8b},
  {32'hc3dc934e, 32'hc43e8157, 32'hc5809431},
  {32'h44466f25, 32'h43f5b8a3, 32'h4351350b},
  {32'hc410df20, 32'hc4bdfdcc, 32'hc3808516},
  {32'hc363e2b0, 32'h44baf519, 32'h446181e0},
  {32'hc37a44f9, 32'hc4b8c526, 32'h438ac553},
  {32'h44e278ad, 32'h439ec4bb, 32'h43aaa7ac},
  {32'hc43279c8, 32'hc4dcad89, 32'h42d08131},
  {32'hc3947aeb, 32'h43ae4980, 32'h424db9eb},
  {32'hc566bb4d, 32'hc2ff423f, 32'hc3bf7abd},
  {32'h44ae5c9d, 32'hc48b5fa2, 32'h435d8175},
  {32'h43a8e708, 32'hc481d326, 32'hc461b06c},
  {32'h43bf0dda, 32'hc4655516, 32'h4506be3e},
  {32'h43821906, 32'hc4dffaaa, 32'hc3c3d5e8},
  {32'hc4823117, 32'h4399e753, 32'h42fd7eab},
  {32'hc3a4d1c4, 32'hc4159a7b, 32'hc4dccea9},
  {32'h4461b0a2, 32'h445baea9, 32'h44542eb5},
  {32'h43456864, 32'hc490750f, 32'hc4ebb69b},
  {32'hc4d2e4c6, 32'h4443b37c, 32'h44487676},
  {32'h4412e2bc, 32'h4389ccb0, 32'hc4fb112b},
  {32'hc3d4a08a, 32'hc4eb5a5a, 32'h44ddb644},
  {32'hc26b2c10, 32'hc2302dcd, 32'hc4a303f4},
  {32'hc3ffb1f8, 32'h44451323, 32'hc38fc193},
  {32'h448b472b, 32'hc4ac466c, 32'h4340fab5},
  {32'hc4970830, 32'h43587b86, 32'h43b47556},
  {32'h43fdc57f, 32'hc3a90d91, 32'hc48bd297},
  {32'hc3bbb8ac, 32'h44e38f02, 32'h44e0f4a8},
  {32'h437191e0, 32'hc4ef6163, 32'hc50cd812},
  {32'hc4d4b730, 32'h43b456b5, 32'h429023bb},
  {32'h44b5159d, 32'hc482395c, 32'hc26b1350},
  {32'hc57e99fa, 32'h43cee040, 32'hc271843a},
  {32'h4499b931, 32'hc37a9f9b, 32'hc3d1dc5b},
  {32'hc373b628, 32'h44e8cd7d, 32'hc2e6c781},
  {32'h44d1af96, 32'hc452ed28, 32'hc3b5008f},
  {32'h43d342fb, 32'hc35f14f2, 32'hc37fc0b4},
  {32'h4529dfe3, 32'hc28c87e3, 32'h43eb9182},
  {32'hc535ed66, 32'hc3073a0a, 32'hc38a5a7a},
  {32'h455cfc72, 32'h43a18f9f, 32'hc3e9e825},
  {32'h44126f6b, 32'h43ce647e, 32'h44f9a242},
  {32'hc3f92f60, 32'hc3afaffa, 32'hc3272864},
  {32'h4297b803, 32'h44519a8e, 32'h43992dfc},
  {32'h4481f7be, 32'h435b10de, 32'h41e2a852},
  {32'h4534bd71, 32'hc3dc3a2e, 32'h41af8c9b},
  {32'hc45563a4, 32'h43ca386e, 32'hc3e538d7},
  {32'h451f42ac, 32'h43d75c09, 32'h3f08834a},
  {32'hc4a6f94b, 32'h44b51e4d, 32'hc38522c9},
  {32'h44aa1186, 32'hc4ba7089, 32'h43cb87d8},
  {32'h43d22224, 32'h444e6ac1, 32'h415b904d},
  {32'h446570a0, 32'hc41ef586, 32'h42101897},
  {32'hc44ccec8, 32'h43bf740b, 32'hc501ee4e},
  {32'h43d5a3c2, 32'hc28b4b4b, 32'hc317b1a8},
  {32'hc53be250, 32'h41d1baff, 32'h42cafd25},
  {32'h44c749e3, 32'hc389c20b, 32'hc33edda9},
  {32'h4372a076, 32'h44afbd9b, 32'hc26d7506},
  {32'hc3b19f87, 32'hc4ddda4a, 32'hc397623b},
  {32'hc49c4e17, 32'h442c7fca, 32'h432dd4ab},
  {32'h44563345, 32'h44158b70, 32'hc43042e6},
  {32'hc4af5fa4, 32'h444f6aad, 32'h44899fa3},
  {32'h43dadce6, 32'h4401a06f, 32'hc49d0792},
  {32'hc47177af, 32'h43789c96, 32'h4296295e},
  {32'h432723ce, 32'hc4eb4c24, 32'hc4670631},
  {32'hc2bad276, 32'h4535637e, 32'hc23c02b3},
  {32'h432f5d54, 32'hc2445a8c, 32'hc4dcdc14},
  {32'hc499c3a6, 32'h44e1b970, 32'h4385c6f4},
  {32'h44fb87d8, 32'hc488768e, 32'hc4781bc7},
  {32'h448b5b12, 32'hc3b7f4f0, 32'hc4c26547},
  {32'hc4afa389, 32'hc2a4c21b, 32'h443aa98c},
  {32'hc22d1f53, 32'h427c1f13, 32'h4412b214},
  {32'hc5622f38, 32'hc1d2f865, 32'h433f65e4},
  {32'h45112f5f, 32'h4360d767, 32'hc409ebd8},
  {32'h44836764, 32'hc42586ae, 32'hc314b361},
  {32'h44aadb2a, 32'h447ccfde, 32'h43808a8d},
  {32'hc4079aee, 32'hc4d82bf3, 32'hc3280438},
  {32'h43bb7c8c, 32'h44a47c78, 32'hc21041c0},
  {32'hc52503c0, 32'hc0b65143, 32'hc1a1f58e},
  {32'h453fb58c, 32'h42b21484, 32'h43276888},
  {32'hc3e69dcc, 32'hc3460ab8, 32'h423558d2},
  {32'hc2287800, 32'h4473f28e, 32'h44b0d15e},
  {32'hc5511c67, 32'hc402654d, 32'h42b77119},
  {32'h44cdb798, 32'hc4204cc8, 32'hc2c648fc},
  {32'hc3f2c876, 32'hc21f593b, 32'hc50240d1},
  {32'h447f9f7e, 32'h442e5be0, 32'h4479425c},
  {32'h43e42515, 32'hc4701f2f, 32'hc3e66b5c},
  {32'h41d7647c, 32'h4330725d, 32'h44a56817},
  {32'hc3fb5eec, 32'h44c1facc, 32'hc4b971f8},
  {32'hc4822952, 32'h43a950e9, 32'hc315d320},
  {32'hc508440a, 32'hc4271c13, 32'hc3275fbc},
  {32'h4331d5f4, 32'h433abf0e, 32'h4487c2a9},
  {32'hc3784970, 32'hc471f5b9, 32'hc3958c75},
  {32'h449b73b5, 32'h448aa354, 32'h43a09b3e},
  {32'hc4ac2c95, 32'hc39836be, 32'hc4881456},
  {32'h43db636a, 32'h4456028f, 32'h431ca972},
  {32'hc44d6123, 32'hc327af9a, 32'hc38f3407},
  {32'hc5378c35, 32'hc3b7931a, 32'h4373690d},
  {32'h436a8d70, 32'h44028ac1, 32'h444b27de},
  {32'h448c525c, 32'hc3f745aa, 32'hc1fa3aee},
  {32'h44f13f30, 32'h440d1749, 32'h42ad0baa},
  {32'hc50a9217, 32'hc42e2872, 32'hc18fdbab},
  {32'h44e977ee, 32'h43d007f4, 32'hc38866ea},
  {32'hc58d79c2, 32'hc3daa005, 32'hc2168f63},
  {32'h448b2690, 32'hc02ec960, 32'h41a53d14},
  {32'hc4dd90e6, 32'h4361de7b, 32'hc38bcde8},
  {32'h448101e0, 32'h444bfee3, 32'h43833ba0},
  {32'hc386d20f, 32'hc5268a9b, 32'hc38084b7},
  {32'hc0b1d840, 32'h40a0688c, 32'hc2a49090},
  {32'hc48fe42d, 32'hc3ea407f, 32'h448f01cd},
  {32'h44ee83fa, 32'h42868930, 32'hc4054f3a},
  {32'hc4cb60ab, 32'h43728480, 32'hc24b250f},
  {32'h43a805f8, 32'h4484a419, 32'h43cff924},
  {32'hc38ed5f9, 32'h4455c36c, 32'h451911c2},
  {32'h45426f3d, 32'hc383a573, 32'h43b47ecf},
  {32'hc4eb3c7b, 32'hc4537641, 32'h44c77f5b},
  {32'hc2ff2181, 32'h455ee829, 32'h439acd28},
  {32'hc325e5f2, 32'hc3b5f851, 32'h44292c96},
  {32'h4521839b, 32'hc2808df6, 32'hc404e870},
  {32'h4292583f, 32'hc5330658, 32'h42a4eca6},
  {32'h449eae2f, 32'hc193d65d, 32'hc431def5},
  {32'hc559c3cc, 32'hc3e0ffa8, 32'h43f6a204},
  {32'h441b69ce, 32'hc2593520, 32'hc5195ec7},
  {32'h4431c35f, 32'hc4c0657c, 32'hc280c8ef},
  {32'hc52362ba, 32'h4347c171, 32'h41030241},
  {32'h45225a7a, 32'h43755058, 32'h42ae00fc},
  {32'hc4828632, 32'h450fa724, 32'h4313338d},
  {32'h43afb474, 32'hc3ac023f, 32'h444e4504},
  {32'h4294bc3a, 32'h44438e97, 32'h435a6299},
  {32'h452c3a12, 32'h44098c76, 32'h42d826c8},
  {32'hc5543b50, 32'h4284b97f, 32'h4397ec7e},
  {32'h450bc056, 32'h4278e872, 32'h440fd538},
  {32'h42e38354, 32'h4468d4c4, 32'hc4b341f7},
  {32'hc0c7da00, 32'hc4b2acc4, 32'h441699c7},
  {32'h44b90cac, 32'h441e0bec, 32'h43045720},
  {32'h44d36d4a, 32'hc4251cd3, 32'h4248c628},
  {32'hc21b3c30, 32'h44a85b77, 32'hc4153594},
  {32'hc4c337f1, 32'h42ac642c, 32'h42fdc2a8},
  {32'hc542994e, 32'hc3ae7af6, 32'h439a8290},
  {32'h4528c3d7, 32'h44316425, 32'h4359b722},
  {32'hc5067f10, 32'h44251c2e, 32'h441e2345},
  {32'h44989928, 32'hc4678efb, 32'h43e17fde},
  {32'h420533e0, 32'h454472f4, 32'h4309fb17},
  {32'h43c94aec, 32'hc3bcbf2e, 32'h44afb62b},
  {32'h420888e1, 32'h4508f824, 32'hc3d1f10a},
  {32'h44616cca, 32'hc4c0bf05, 32'hc3bade8d},
  {32'h44067230, 32'hc3158292, 32'hc4598541},
  {32'h44dfd089, 32'h441bce77, 32'h446557e0},
  {32'hc444c8f6, 32'hc2ee32c9, 32'hc521a106},
  {32'h437bfb20, 32'hc3ede895, 32'h43eb5e0f},
  {32'hc3dbd490, 32'hc46ef85a, 32'hc499f596},
  {32'h44b20ea6, 32'h44350201, 32'h43cea3f6},
  {32'hc492c79c, 32'hc3d64935, 32'h43f1945c},
  {32'hc410acec, 32'h43ccae86, 32'h4362299d},
  {32'h436aeea8, 32'h4384a1b0, 32'h44a196de},
  {32'hc4a2b956, 32'h44826a2c, 32'hc360591c},
  {32'hc386cd5e, 32'hc44987cb, 32'h439535a4},
  {32'hc3e62ed8, 32'h4465607e, 32'hc52054d0},
  {32'h44ea178e, 32'hc3461f16, 32'h441bcf6a},
  {32'hc22043d4, 32'h4254a8d1, 32'h45088dad},
  {32'hc52cf728, 32'h43fa0243, 32'hc3c20ec0},
  {32'hc1c75e22, 32'hc4f9b209, 32'h442d396e},
  {32'hc4884d4e, 32'h43cfcc39, 32'hc30ed482},
  {32'hc45d4893, 32'h431adae7, 32'hc47bd129},
  {32'h441035fb, 32'hc383ae1b, 32'h44a7fff6},
  {32'h43c8b9b6, 32'h44a68af5, 32'h4172f260},
  {32'h436f7be5, 32'h42c0b8e0, 32'h44faf9db},
  {32'hc3232596, 32'h45113a2e, 32'hc3a78453},
  {32'h453bf42e, 32'hc4399cc9, 32'h4399817e},
  {32'hc52b1459, 32'hc4613c50, 32'hc4125e15},
  {32'hc3a84502, 32'hc0c3302f, 32'h43e01465},
  {32'h43dc05f7, 32'hc3c40f47, 32'hc3898ac1},
  {32'h44c6c400, 32'hc4573f1f, 32'hc2275449},
  {32'hc503afce, 32'hc273f432, 32'h438f8b43},
  {32'h44f34542, 32'hc34cd26e, 32'hc2c28628},
  {32'hc41ac512, 32'h451b6b8f, 32'h43caaaaf},
  {32'h43291778, 32'hc53ba7a9, 32'hc3b47f11},
  {32'hc49442d7, 32'hc383e173, 32'hc083ea80},
  {32'h4371c3b9, 32'h432de3e0, 32'hc4d4a0e7},
  {32'h4493d206, 32'h43abfba0, 32'h43d3989a},
  {32'h424953e0, 32'hc2df60a7, 32'h4516ec3a},
  {32'h44431044, 32'h431c9982, 32'hc482bcb6},
  {32'hc29b80c5, 32'hc3694860, 32'h43c5ab2d},
  {32'hc3138df2, 32'hc377ad1b, 32'hc569cac9},
  {32'hc4f72bb6, 32'h438239d8, 32'h4463ba6b},
  {32'hc44bfb56, 32'hc3257d44, 32'hc130d2b4},
  {32'h4408b088, 32'h4418d475, 32'h41d440e6},
  {32'hc431904d, 32'h434e5d1f, 32'hc30db45f},
  {32'hc3bf8b2e, 32'hc39c571e, 32'hc502d872},
  {32'h42697507, 32'hc42e7368, 32'hc53c8f0f},
  {32'hc45c6c46, 32'hc47c9939, 32'h43243edc},
  {32'h401faf00, 32'h44b81d90, 32'hc315ea8a},
  {32'hc512dd80, 32'hc3da98d0, 32'h43b01fea},
  {32'h42cc1f80, 32'h44050de8, 32'hc5158a70},
  {32'h44d583b1, 32'h43cba380, 32'h43f55477},
  {32'h44b93b23, 32'h4357373d, 32'hc35a8672},
  {32'hc509532c, 32'hc3b8bd85, 32'h434fd6cf},
  {32'h442ae039, 32'h43948da6, 32'h41fa0f18},
  {32'hc4c6f4ce, 32'hc44efa98, 32'h41e40a2e},
  {32'h42f7f100, 32'h436d8869, 32'h42f20344},
  {32'h442b27c6, 32'h433ce6a7, 32'hc3312e5f},
  {32'h45365127, 32'h4428e1df, 32'h429329d0},
  {32'hc44dd7d8, 32'hc4d560ab, 32'h43626611},
  {32'h43fe9563, 32'h4409cd49, 32'h42c39c4b},
  {32'h41916e3c, 32'h43e00b81, 32'h4467e5d3},
  {32'hc420bfec, 32'h451b49b5, 32'hc4b2c667},
  {32'h449c0236, 32'h43aee29d, 32'h445ad294},
  {32'hc3b21656, 32'h43846325, 32'h4349b6c8},
  {32'h440caa9b, 32'hc2f5b1c3, 32'h4504306e},
  {32'hc2e3424f, 32'hc507a820, 32'h41fabcd8},
  {32'h4540d7e6, 32'hc3c5bde8, 32'hc37f5f62},
  {32'hc3b7ca37, 32'hc44c1afe, 32'hc504a6b4},
  {32'h4318b542, 32'h448fb197, 32'h44b5dd9e},
  {32'h43d98f4c, 32'h446434a9, 32'hc43c3ea3},
  {32'h42d1583a, 32'h4527cbc0, 32'h43b1cb5f},
  {32'h439a7107, 32'hc4112a14, 32'hc46b17a2},
  {32'hc09cf92a, 32'h43046e6e, 32'h44e55cca},
  {32'h42ed65dc, 32'hc5103b21, 32'hc3ec108c},
  {32'h44183139, 32'h4480526a, 32'h4403e0bf},
  {32'h40bea478, 32'h428410d1, 32'hc2daa9e7},
  {32'h44012600, 32'h44c5ee34, 32'h44587e65},
  {32'hc338af14, 32'hc4837601, 32'hc514d8bc},
  {32'hc4b23cd6, 32'h431a51b2, 32'h435c16a9},
  {32'hc4ef9441, 32'hc41dcbca, 32'hc3b985cc},
  {32'h43c25ad0, 32'h4493e167, 32'h43f34de0},
  {32'h43b56e6c, 32'hc4ea6872, 32'hc411abc3},
  {32'h439c6a29, 32'h454ce657, 32'h440dee32},
  {32'hc4d0b173, 32'hc484d3fe, 32'hc35441d3},
  {32'h4420c21e, 32'hc2e43402, 32'hc2fc14b5},
  {32'hc4cf78bc, 32'hc3f239f6, 32'h42e3c33c},
  {32'h44f6e2b0, 32'h4358b4f6, 32'h437b31fd},
  {32'h43171d80, 32'h42d790af, 32'hc4f74e09},
  {32'hc2caa56a, 32'h44c29b61, 32'h43d2dd1a},
  {32'hc2bbc458, 32'h4324eb44, 32'hc48b27d8},
  {32'hc412c130, 32'h4519ccda, 32'h42de65ce},
  {32'h44416dca, 32'hc411a49f, 32'hc3fd9a16},
  {32'h4369b2e4, 32'h43b7f804, 32'h43505aaa},
  {32'h4397e71a, 32'h429cb984, 32'hc374890b},
  {32'hc4a3432b, 32'h43c591e4, 32'h4488f7c8},
  {32'hc3fbaf62, 32'hc3ccfb3e, 32'h43c45573},
  {32'h4336e690, 32'h44d35c1a, 32'h44505261},
  {32'hc2c46eac, 32'hc4dfa2ec, 32'hc4046571},
  {32'h4426d35c, 32'hc412eb61, 32'h443c19ad},
  {32'h450e356d, 32'hc415131a, 32'hc1596fa2},
  {32'hc3c381fe, 32'hc3b95531, 32'h4525f557},
  {32'hc3768c6e, 32'hc471dec2, 32'hc3f4d104},
  {32'hc50dee58, 32'h425c7c6b, 32'h43b5e978},
  {32'h442ba5fe, 32'hc4580d8a, 32'hc4b3f934},
  {32'hc42fa550, 32'hc19d6980, 32'hc18c0d02},
  {32'h44c6e81c, 32'hc4ad9478, 32'hc2c06392},
  {32'hc49a72e0, 32'h449301fa, 32'hc34ae8e5},
  {32'h446c9bd1, 32'hc3226805, 32'hc2805317},
  {32'h432ff502, 32'h44351bff, 32'h43444141},
  {32'h4509794c, 32'hc4b685af, 32'h4388ff96},
  {32'hc4d42bf3, 32'h43a0f9f4, 32'h43190104},
  {32'h451123d4, 32'h43dc2b8e, 32'h43e0294a},
  {32'hc55e476e, 32'h439340d7, 32'h4332dc68},
  {32'hc50834d3, 32'h432b8347, 32'hc377ae8b},
  {32'h4426629e, 32'hc445e4b8, 32'h448be70d},
  {32'hc5684674, 32'hc0a7499e, 32'h431afbf9},
  {32'h44faac7e, 32'h3e87186a, 32'h44ad0996},
  {32'h43ff19a2, 32'h4411c916, 32'hc3018632},
  {32'h43f7b77c, 32'hc4f06d86, 32'h42a0cdf8},
  {32'hc41c5304, 32'h44575467, 32'h43fc83ce},
  {32'h43539898, 32'hc49197ef, 32'h4319d204},
  {32'hc588d96e, 32'h437e05d5, 32'hc3af693f},
  {32'h43bcc0e6, 32'hc51e29b4, 32'hc365c8e0},
  {32'hc437f886, 32'h437731de, 32'hc2cd353c},
  {32'h44f639fa, 32'h43172804, 32'h43993a39},
  {32'hc32a8a46, 32'h434dcdb4, 32'hc38e55b9},
  {32'h43c9a6fa, 32'hc33bb8ed, 32'hc4161445},
  {32'hc4b6bb5d, 32'h43e07ef3, 32'h4317b078},
  {32'hc1f2d9a0, 32'hc5367fb4, 32'hc2341076},
  {32'h43488178, 32'h44077990, 32'h4507e844},
  {32'h44e1db20, 32'hc44a3eb0, 32'h431324d5},
  {32'hc50e0465, 32'hc359a7f8, 32'hc34c90eb},
  {32'h44d6c678, 32'hc41f5c97, 32'hc3775df3},
  {32'hc55c96b0, 32'h43e84749, 32'h441a6d0c},
  {32'h453b73c3, 32'hc318b690, 32'hc42d763d},
  {32'hc3f3a863, 32'hc38e640c, 32'h43876b90},
  {32'h43d76e10, 32'hc4d7ab45, 32'hc365d4f0},
  {32'h42283622, 32'h453faa4f, 32'h435443f6},
  {32'h44d318e6, 32'hc39f42ec, 32'hc3e00ef2},
  {32'hc56750f2, 32'h42645654, 32'hc2daf442},
  {32'h426ed480, 32'hc4c24c13, 32'hc4cd598d},
  {32'h446a552e, 32'h435c7aca, 32'h428ebcb8},
  {32'hc5044076, 32'h437de70e, 32'hc208dc7e},
  {32'hc3ad8ce0, 32'h44289eae, 32'hc498c7da},
  {32'hc3e72e4f, 32'hc512ba59, 32'h411b952d},
  {32'h45316bbc, 32'hc1a72f58, 32'hc3ecfb87},
  {32'h4401e17d, 32'hc4904c12, 32'h42be4980},
  {32'h44df7116, 32'h449a77aa, 32'hc3e3acd0},
  {32'hc4eddea3, 32'hc4b8d5c6, 32'h4352bcb0},
  {32'h435938d2, 32'h4515fb3c, 32'h435561b6},
  {32'hc44ae222, 32'h434099a6, 32'h44d7d71a},
  {32'h45026a71, 32'h43f7dbb5, 32'h433a0140},
  {32'h440a885d, 32'hc309b643, 32'h434d6c76},
  {32'h44736088, 32'hc2af65cb, 32'h4491afd0},
  {32'hc52e5560, 32'hc402cd4c, 32'h42aaee90},
  {32'hc4582619, 32'h448639e8, 32'h43aff524},
  {32'hc49599e3, 32'hc31bea67, 32'hc30432b4},
  {32'h44709a9b, 32'h43e96035, 32'h44b0a7f7},
  {32'h4500ead1, 32'h41313306, 32'h44009def},
  {32'h44867416, 32'hc4a3645c, 32'h44db1000},
  {32'hc58b91cd, 32'h42d79d98, 32'hc2e31f95},
  {32'h4515d5f6, 32'h435023b0, 32'hc4030f03},
  {32'hc26feabd, 32'hc5417de4, 32'hc48b0987},
  {32'h439befe2, 32'h4380c34c, 32'h448886b6},
  {32'h44c22905, 32'h42ae1dfb, 32'h438e9bcb},
  {32'h4325a73e, 32'h4444b5d5, 32'h446ce648},
  {32'hc3616cbe, 32'hc5325132, 32'hc2aa34c8},
  {32'h42d94a04, 32'hc2f9fe16, 32'h44968192},
  {32'h44d5f5b5, 32'h4221729b, 32'hc296003c},
  {32'hc3b32426, 32'hc382683b, 32'h43201e40},
  {32'h444d7388, 32'h44d354e7, 32'h440e56c9},
  {32'hc48c0aaf, 32'h4341f136, 32'hc31518b0},
  {32'h44d79769, 32'h442896d8, 32'hc39faac0},
  {32'hc4ad09d1, 32'hc48ec2e7, 32'hc27c0492},
  {32'h44a34ef4, 32'h42af5802, 32'hc3530980},
  {32'hc4071bd8, 32'hc400d2fc, 32'hc39fa270},
  {32'h43ec85c8, 32'h44585115, 32'h44893f32},
  {32'hc421021e, 32'hc0dbccf2, 32'hc3415126},
  {32'h4449d9a6, 32'h447b517a, 32'hc412b743},
  {32'hc5037c55, 32'h41c56cf4, 32'hc407489f},
  {32'hc404b47b, 32'h422d9a0e, 32'hc4fb7068},
  {32'hc3b6b6fe, 32'hc51331e8, 32'h43365538},
  {32'h44356627, 32'h4480fe0d, 32'hc4aff027},
  {32'hc3699440, 32'h42ba56aa, 32'hc3f2f5c3},
  {32'h443e3409, 32'h430a4aee, 32'hc458545f},
  {32'hc4a0f010, 32'h41e20b34, 32'hc338bcd0},
  {32'h43ba73b5, 32'h444e78d3, 32'hc306a8d0},
  {32'hc4171288, 32'hc4cfbe87, 32'hc38137e1},
  {32'h449be2a6, 32'h443f57be, 32'hc4bb05de},
  {32'h43b58793, 32'hc50eb79e, 32'h439a7c19},
  {32'h44b5b696, 32'h42a7037b, 32'hc38918b9},
  {32'hc52a6b9d, 32'h43f64c1c, 32'h42bf01ed},
  {32'h44804253, 32'h42d11ae5, 32'hc4b73228},
  {32'hc513833c, 32'h439320b4, 32'h4480ece4},
  {32'h43ae3717, 32'hc3a77a7f, 32'hc5671e9f},
  {32'h44587714, 32'hc49aaa12, 32'hc391f914},
  {32'hc51023cc, 32'h4450e934, 32'h43a6ebde},
  {32'h44a3ecd0, 32'h43070e3b, 32'h441a4a17},
  {32'h4199c5a7, 32'h45849929, 32'hc21b9920},
  {32'h442fe167, 32'hc5096273, 32'h43706cce},
  {32'hc5307410, 32'hc3b74384, 32'h43030789},
  {32'h44f3df0c, 32'h43a664bd, 32'h42079555},
  {32'hc5531cd7, 32'hc437eecc, 32'h43941c85},
  {32'hc4ad85ac, 32'hc3755f6e, 32'h4341131e},
  {32'hc46a0223, 32'h44414960, 32'hc4ed8ada},
  {32'h4449ed24, 32'hc42ea45f, 32'h4414fc7b},
  {32'hc39c93e2, 32'h44cbd842, 32'hc231a033},
  {32'hc1c130b0, 32'hc4d923db, 32'h44288b7e},
  {32'hc257f259, 32'h434c5c41, 32'hc4f27578},
  {32'hc3afccdc, 32'hc4b548dc, 32'hc3dac6f8},
  {32'hc477534b, 32'hc2cebc64, 32'hc3f5259a},
  {32'h44af5cd4, 32'h438acc0b, 32'h44751d6f},
  {32'h44986ecc, 32'hc34b4881, 32'hc427bc5d},
  {32'h43e3a378, 32'hc49926ce, 32'h4503d9e6},
  {32'hc4237d34, 32'h44e140af, 32'hc4bcfe24},
  {32'h448872df, 32'h4376c8f9, 32'h41ccf0bf},
  {32'hc501b20f, 32'h446d73b6, 32'hc3b14df4},
  {32'h4499f268, 32'h42958eea, 32'hc3c50bbb},
  {32'hc53f1012, 32'h4303a86b, 32'hc3af0082},
  {32'h4200f580, 32'h4272008a, 32'h445aa54e},
  {32'hc44564b6, 32'hc40d2a30, 32'hc51c0c49},
  {32'h44181c75, 32'hc4015a17, 32'h42bcfa4a},
  {32'h44812231, 32'hc3946889, 32'hc42d49dd},
  {32'h43968899, 32'h43287fa6, 32'h4511ca76},
  {32'h44b89708, 32'h42b49a1e, 32'h42f00029},
  {32'h44231616, 32'h4454c6a4, 32'hc41b051e},
  {32'h44316fcc, 32'hc29b54a5, 32'h44de9c8b},
  {32'hc3f4e3e6, 32'hc3acae3c, 32'hc4b8085f},
  {32'h45299d81, 32'h43756f4c, 32'hc3d73cf8},
  {32'h43847079, 32'h44f754c7, 32'hc40f5308},
  {32'h44645664, 32'hc49d44fa, 32'h438dcf7c},
  {32'h44f74308, 32'h442ba178, 32'h4434b189},
  {32'hc41f7c15, 32'h42a2827e, 32'hc497da04},
  {32'h424f061c, 32'h446d23c4, 32'h437bf9d7},
  {32'h44efb148, 32'h436b6855, 32'h42cff465},
  {32'hc2c45380, 32'h42e4cb91, 32'hc4c6a82c},
  {32'h44a42d41, 32'hc315387a, 32'h44474a61},
  {32'hc434eaf3, 32'h43656175, 32'hc420fba1},
  {32'h44a97602, 32'h42713251, 32'h44804e4c},
  {32'h4384025e, 32'h42a549f8, 32'hc4fbb30f},
  {32'h44144204, 32'h440d5e67, 32'h43d561a8},
  {32'hc48fbb10, 32'h4427c72e, 32'hc4199a5b},
  {32'h439a8c20, 32'hc28922ee, 32'h43485c96},
  {32'hc3afcc5c, 32'h4459922c, 32'h438995b8},
  {32'h427dd67c, 32'hc55ac81e, 32'hc1c024d0},
  {32'hc4b3fa23, 32'h4449b803, 32'h43291a86},
  {32'hc2758790, 32'hc4791082, 32'hc381baff},
  {32'hc54df095, 32'h445a2f85, 32'h44406b22},
  {32'h43a7ed7c, 32'hc4927245, 32'hc4232599},
  {32'h4440e6f6, 32'hc3418c7d, 32'h44c92500},
  {32'h43cf45f6, 32'hc478cb21, 32'hc4a180c8},
  {32'hc3728f47, 32'h441587b9, 32'h452d7759},
  {32'hc37a93f4, 32'hc4378530, 32'h44c4bbe2},
  {32'h44782b6e, 32'h4465b308, 32'hc34c3519},
  {32'h43bf1732, 32'hc26e1bc7, 32'h43017e87},
  {32'h445f3ca8, 32'h4469d431, 32'hc47fd56e},
  {32'hc438a415, 32'hc4f254e1, 32'h43915c62},
  {32'hc3c706e5, 32'h442719b8, 32'hc4ae65ed},
  {32'hc0d00798, 32'h43bfef48, 32'h41979d0a},
  {32'hc340a1e2, 32'h43419a08, 32'h44a4268c},
  {32'h44fb56e6, 32'h42955dc5, 32'hc4447a0d},
  {32'h437cc6c0, 32'h4447f746, 32'hc31bf920},
  {32'hc4806eb2, 32'hc3a50480, 32'h438b7713},
  {32'hc3c5b466, 32'h43f5269f, 32'hc4985da8},
  {32'hc4954c94, 32'hc44627ff, 32'h44315906},
  {32'h451be88d, 32'h43c09841, 32'hc3e8aa6f},
  {32'h44a8bb99, 32'hc3d836f8, 32'h4107d2c8},
  {32'h455fe0ee, 32'hc3a5f5c6, 32'h42571887},
  {32'hc4c7fe2c, 32'h44464d11, 32'h445ead30},
  {32'h4545eca5, 32'h438d5385, 32'h42ad2a31},
  {32'hc3d8b152, 32'hc5195a8e, 32'h440c080f},
  {32'h44fe7505, 32'h448034a0, 32'h437b9758},
  {32'hc52dad11, 32'h431e1dbd, 32'h4380165d},
  {32'h42b52520, 32'h450ddecf, 32'h43d53e5e},
  {32'hc490510e, 32'hc4d6601f, 32'h40e63c48},
  {32'h43dd71d8, 32'h43067b0f, 32'hc3d3ef97},
  {32'h4376e774, 32'h43c39fdc, 32'h443c21e3},
  {32'h43b60ba4, 32'hc48e2e71, 32'hc1e41b80},
  {32'h43a5d9b7, 32'hc43bf683, 32'h448c3917},
  {32'hc262cf28, 32'hc23e0498, 32'hc4cf0104},
  {32'h43a04cba, 32'h4498d66a, 32'h444b2291},
  {32'hc4505086, 32'hc3eeaf92, 32'hc44c05fc},
  {32'hc29c72e0, 32'h43aafa11, 32'h44125322},
  {32'hc4430951, 32'hc4d63e70, 32'hc49ca865},
  {32'hc3c622b7, 32'h448fefc2, 32'h453e0bbe},
  {32'h44053af5, 32'hc3093c9b, 32'hc421febe},
  {32'h43279a84, 32'h423b6ec9, 32'h44997a3c},
  {32'hc5000a20, 32'h40f24210, 32'hc3f56255},
  {32'hc35ffcbc, 32'hc2c1e00f, 32'h44c4418c},
  {32'hc508f493, 32'hc264740e, 32'hc381865a},
  {32'h43ed3810, 32'h45391f5f, 32'h3fc6a466},
  {32'h44ef7725, 32'hc3a25945, 32'h42c2c03c},
  {32'hc2e38480, 32'h44a55749, 32'h44a0c33c},
  {32'hc4b73149, 32'hc4050029, 32'hc40d16c9},
  {32'h426d3084, 32'h44cab8e3, 32'h438a5f2e},
  {32'hc50727d5, 32'hc3f541d4, 32'hc37793c8},
  {32'h43b4a149, 32'h457d14c4, 32'h4236cd7d},
  {32'h449ecfe2, 32'hc431c5bb, 32'h428e34d6},
  {32'h450ada12, 32'hc290ed84, 32'h438e0096},
  {32'hc3da9080, 32'hc525f1ef, 32'hc25c59c8},
  {32'h43833b35, 32'hc23df170, 32'h43608310},
  {32'hc5815854, 32'hc2f3f740, 32'hc3c74c31},
  {32'h44c8f011, 32'h43511317, 32'h44334bda},
  {32'h442fa937, 32'hc3ccaf99, 32'hc4b240d9},
  {32'h43e10208, 32'hc3db4ad1, 32'h4501f0fd},
  {32'hc43896e0, 32'hc388f8ad, 32'hc3f1429c},
  {32'hc3203ba4, 32'h43667bc0, 32'h448757e4},
  {32'h44d02c39, 32'hc3e4541f, 32'hc4798ca8},
  {32'h44ce8dbe, 32'h43e96556, 32'h3f886064},
  {32'h44fa03dc, 32'hc44b7ea3, 32'hc3a4976d},
  {32'hc38d8e1e, 32'h4424b670, 32'h45838fa3},
  {32'h444472ae, 32'hc490ecf8, 32'hc2edc357},
  {32'hc430e36b, 32'hc384e8b5, 32'h4487a642},
  {32'h40624408, 32'h44bfa689, 32'hc50fa87c},
  {32'hc4dd013f, 32'h409b97fa, 32'hc26cedc5},
  {32'h441bfa01, 32'hc47f0b7e, 32'hc2e04840},
  {32'hc418fa98, 32'h43025218, 32'h44772cf9},
  {32'h43de1349, 32'hc472fea6, 32'hc1b79a27},
  {32'hc396d69c, 32'h4459842a, 32'h44a13b32},
  {32'h4401a4aa, 32'hc4f4c3e1, 32'hc4bb0a09},
  {32'h44e8f53b, 32'h431583e5, 32'h43d889c9},
  {32'h4474f8ce, 32'hc4b3fe83, 32'h436da05e},
  {32'hc315a660, 32'h44cd6ff0, 32'h4457afd7},
  {32'hc514db58, 32'hc2d54219, 32'h429e0504},
  {32'hc52e81f2, 32'h4439dfe3, 32'hc2db9385},
  {32'h431f5db0, 32'hc54c6d8a, 32'hc3bed4e2},
  {32'hc50a6112, 32'hc255205c, 32'h4432e3c9},
  {32'h453158f2, 32'h4370d153, 32'hc373d96a},
  {32'hc4c81c70, 32'h44122c90, 32'hc21ce44c},
  {32'h4454d84a, 32'hc30c8aba, 32'hc307a9e3},
  {32'hc4e2c224, 32'h43626ca5, 32'hc20d3f88},
  {32'hc46e18da, 32'h4293e17d, 32'hc5341145},
  {32'h44a2d3b7, 32'hc39d1ec0, 32'hc29ba0ac},
  {32'h44b3229e, 32'h4301cdc9, 32'h40c9d2ec},
  {32'h440f3efe, 32'hc48635c4, 32'h42963d6c},
  {32'hc2a19869, 32'h45088e6c, 32'h44335b1a},
  {32'h44eef0ee, 32'h441e35d6, 32'hc3e5d204},
  {32'hc49d1c8d, 32'h44ed9525, 32'hc2eb876c},
  {32'h44bdfda8, 32'hc49ca97c, 32'h442efedc},
  {32'hc52378d7, 32'hc3585f50, 32'hc2551772},
  {32'h443e5eae, 32'hc4190198, 32'h452624e6},
  {32'hc51cc798, 32'h4355f4fa, 32'hc2948dbe},
  {32'hc4196e9b, 32'hc438ea8e, 32'hc3972843},
  {32'h435869f6, 32'h452cc522, 32'h43b42661},
  {32'h4395dc9e, 32'hc527dfe2, 32'hc35c9f7d},
  {32'h43c17122, 32'h44170cc9, 32'h44eae1f6},
  {32'h44b6f676, 32'hc0b96c40, 32'hc39e068c},
  {32'hc2ccec44, 32'h44e7b957, 32'h4321a065},
  {32'h444d2b47, 32'hc277133a, 32'hc4192fad},
  {32'hc428f399, 32'hc39ddc00, 32'h44c2440b},
  {32'h43214380, 32'hc413de19, 32'hc48c58c8},
  {32'h439ba1df, 32'h4266623e, 32'h44884b5c},
  {32'h431332d9, 32'hc41b3e0a, 32'hc4689002},
  {32'hc4a8e3ab, 32'h44618dd5, 32'h41beb9be},
  {32'h439f528c, 32'hc4e8d53a, 32'hc198af7e},
  {32'hc57229bb, 32'h4355ec6a, 32'hc38d32ae},
  {32'h43a3c015, 32'hc5078c7b, 32'hc3d068d9},
  {32'h4417e1dc, 32'h437b79a3, 32'hc513c038},
  {32'hc4435e56, 32'h43947a84, 32'h4504d143},
  {32'h42cf8774, 32'h446e8cd1, 32'hc4a8b1ed},
  {32'hc3b0200e, 32'hc4b33db2, 32'h427d3df5},
  {32'h44682af8, 32'h4326bd1c, 32'hc3e36c1c},
  {32'h44ed64e0, 32'hc2aec918, 32'hc31ae56e},
  {32'h45142de8, 32'h443cbdc2, 32'hc381cdc9},
  {32'hc3f72741, 32'hc55c8fd7, 32'h4318a90d},
  {32'h43e1e8b6, 32'h43cd420d, 32'h41ab2c8b},
  {32'hc4476326, 32'hc42971e2, 32'h4407f3d2},
  {32'h4388cd08, 32'h43f91888, 32'h43868b08},
  {32'hc4504794, 32'hc3f94e52, 32'h440c8268},
  {32'h451c8c56, 32'h43373919, 32'h43dcc34e},
  {32'h42e378f8, 32'hc540dcbb, 32'hc3b770f5},
  {32'h446dbbb8, 32'h420f1491, 32'h4307a607},
  {32'hc443306c, 32'hc467218f, 32'hc3f52e4d},
  {32'h4468af52, 32'h4476dd40, 32'hc062bc0c},
  {32'hc333e8bc, 32'hc43b9acd, 32'hc44485e1},
  {32'h445b845c, 32'hc48efbdb, 32'h44156bea},
  {32'hc5730c7b, 32'hc2bd5558, 32'hc380becc},
  {32'hc49b0cd6, 32'hc3afd012, 32'hc30ddb54},
  {32'hc4606e76, 32'hc4ab2c45, 32'hc4009056},
  {32'hc2f82670, 32'h44ec5602, 32'h443f8ef5},
  {32'hc11f3bbd, 32'hc33d10ac, 32'hc486e11f},
  {32'hc3497ad7, 32'h45345b8f, 32'h43a308fe},
  {32'hc50e0386, 32'hc4025d26, 32'hc23cf858},
  {32'hc3c7b4d5, 32'h436dc5b4, 32'h445d78ef},
  {32'h43f81a87, 32'h44a63db1, 32'hc3e77138},
  {32'h4285e120, 32'hc52b8aa3, 32'hc395f83c},
  {32'h44fc668a, 32'h443388aa, 32'h44005d04},
  {32'hc3da4f98, 32'hc4810e81, 32'h43b4b511},
  {32'h447892b4, 32'h44e8af52, 32'h4282f496},
  {32'hc51f79f3, 32'hc39a2b35, 32'h41b286e9},
  {32'h44d1efdd, 32'h43917ce8, 32'hc393d595},
  {32'hc37859e0, 32'hc4533d7c, 32'hc42bc627},
  {32'h444d6c9d, 32'h44939457, 32'h44929d71},
  {32'hc3cdf3fe, 32'h437ef4b5, 32'hc32e3cc2},
  {32'h44a1551c, 32'h4418e7d6, 32'hc4615c62},
  {32'h42d39692, 32'hc425bb4b, 32'h44b77126},
  {32'h44a3ed2e, 32'h438412a5, 32'hc35a73cf},
  {32'hc4a64db5, 32'hc3f9dc4a, 32'h43d2fbfd},
  {32'h4483d422, 32'h44093f61, 32'hc3026e96},
  {32'h44390dde, 32'h43983ff3, 32'h447889d1},
  {32'h44b3efa7, 32'h42effb78, 32'hc3bd88b1},
  {32'hc388a5df, 32'hc3e4e97d, 32'h448bf049},
  {32'hc4908535, 32'hc1f8acc5, 32'hc4117b4c},
  {32'hc5037f56, 32'hc42bd847, 32'h4398c002},
  {32'h44c404f4, 32'h44b71088, 32'hc360cda2},
  {32'hc5322745, 32'hc1f03a22, 32'hc346483d},
  {32'h44faf948, 32'h43d4b81e, 32'hc3aaa07a},
  {32'h443aa26d, 32'hc51718b8, 32'h43aabb16},
  {32'h45323ea6, 32'h42ec24cf, 32'h4287abc7},
  {32'hc49bc3f0, 32'h43b750a3, 32'h44887ec4},
  {32'h445e3385, 32'hc396410a, 32'hc53949c7},
  {32'h450306b4, 32'hc451ba1b, 32'hc311b4b0},
  {32'hc4a4e559, 32'h445940cd, 32'h4368ca11},
  {32'h4261c107, 32'hc3e26dea, 32'hc41b6693},
  {32'hc214a755, 32'h453b6381, 32'hc3931497},
  {32'h415ea51c, 32'hc55600e4, 32'h42b63810},
  {32'hc52dd294, 32'hc2e52463, 32'hc3e6b1c8},
  {32'h4427bd71, 32'hc3cee040, 32'hc39578d1},
  {32'hc4e6d3f8, 32'h442573fd, 32'h44200930},
  {32'h44871d17, 32'hc4744da4, 32'hc3c057a3},
  {32'h439ef299, 32'h45262f0a, 32'h4403c57d},
  {32'hc34571f9, 32'hc5191333, 32'hc387c426},
  {32'h440df48b, 32'h436a45d7, 32'hc4cfb156},
  {32'h4453403c, 32'h438d3758, 32'h45000b66},
  {32'hc4ef40b3, 32'h44060236, 32'hc2ffe1d0},
  {32'hc4bb1e4e, 32'hc16f8500, 32'hc31dbb00},
  {32'hc4e33cf2, 32'hc3ba0f2c, 32'hc3e64414},
  {32'h4427b8ef, 32'h44126b0e, 32'h44f4a9ab},
  {32'h44d27f39, 32'hc20719af, 32'h4391b95c},
  {32'h445cb8f4, 32'hc4bb0bc8, 32'h43fc74cd},
  {32'hc49a8f87, 32'h44dd0ec6, 32'hc38cbd84},
  {32'hc3e39b54, 32'hc318e008, 32'h4474ce45},
  {32'hc423e440, 32'h44741c6e, 32'h42679fd2},
  {32'h450b3b9a, 32'hc3cb98bf, 32'hc11a555c},
  {32'h44104b6f, 32'h42bb3077, 32'hc4126f7b},
  {32'h4448a128, 32'h4387e4b2, 32'h44c8addb},
  {32'hc41a84fc, 32'h43a8652c, 32'hc475707b},
  {32'h43ea23e7, 32'h442b047e, 32'h44d2a9f5},
  {32'hc3107cdf, 32'hc4d07f57, 32'hc50cb4c9},
  {32'hc417e693, 32'hc4062825, 32'h431611bc},
  {32'h4101bd6e, 32'h441e6624, 32'hc40cc6cb},
  {32'hc3614f69, 32'h4309c2d7, 32'hc48d8f64},
  {32'h450f80ee, 32'hc44daff2, 32'h434d5188},
  {32'hc52a0b1c, 32'hc2c18e13, 32'hc3d27fe5},
  {32'h43c18d40, 32'hc429d580, 32'hc302d9b2},
  {32'hc49aadaa, 32'h43bfc967, 32'hc424cbb4},
  {32'h44876ab5, 32'hc33a2f23, 32'h449f3de1},
  {32'h4438d4ec, 32'hc4e17bcd, 32'h44f97cf1},
  {32'hc5444841, 32'h43099cef, 32'h4402cde4},
  {32'hc42ab0c9, 32'hc3803794, 32'h4426867a},
  {32'hc4f32d52, 32'hc39848f0, 32'hc40d4b7d},
  {32'hc3990ac0, 32'h450aa8b1, 32'h44249891},
  {32'h4378a94e, 32'hc39e1e08, 32'h45310a20},
  {32'hc4f6dbea, 32'hc3a1926e, 32'h434c1209},
  {32'hc29100da, 32'hc33599b3, 32'h4543c2c7},
  {32'hc41e5c2e, 32'h43b4545b, 32'hc4c768b8},
  {32'hc3a90bf9, 32'hc4174cd3, 32'h42cacb0b},
  {32'hc49a3d4a, 32'h44179842, 32'h438ceebc},
  {32'h43e56240, 32'hc3d1a920, 32'h441ebf5a},
  {32'hc4796bac, 32'hc31955cc, 32'hc3ed3fae},
  {32'h44b03bed, 32'hc4b6336d, 32'h43a96ca2},
  {32'hc54e73ad, 32'h43b934b0, 32'h42b7ce7b},
  {32'h4478ef9e, 32'hc4b33897, 32'h42cf0941},
  {32'hc41a6f32, 32'h45334d2f, 32'h437d8b92},
  {32'h4524ad91, 32'hc437ef83, 32'h43932365},
  {32'h4454195d, 32'h4215cbfb, 32'h44eb9db2},
  {32'hc361ce72, 32'h451df5b0, 32'hc4dbe8ca},
  {32'hc4bcf1ee, 32'h43c9ecc5, 32'h44097a60},
  {32'h43372c84, 32'hc534fe92, 32'hc0bd0b80},
  {32'h43de43d8, 32'h443adfa5, 32'hc428c02c},
  {32'hc4c9b946, 32'hc42b081f, 32'hc22eb7bb},
  {32'h44ba45cf, 32'hc2045ae6, 32'hc4a6a8a0},
  {32'hc3aa1dde, 32'hc52074c0, 32'h4359526a},
  {32'h43b6e578, 32'h44355d99, 32'hc26a779b},
  {32'h44c99a51, 32'h43888b07, 32'h43c1e99b},
  {32'hc4097972, 32'h44938739, 32'h4497f568},
  {32'h426d7558, 32'h436d45fc, 32'h4300c3b7},
  {32'h4492ad74, 32'h426b91f8, 32'hc2fbbf83},
  {32'hc3998aa4, 32'hc50da0ab, 32'h431d87d9},
  {32'hc4304521, 32'h445fff8f, 32'hc2667a4a},
  {32'hc4ee1401, 32'hc31b8903, 32'h440122b3},
  {32'hc303d3b2, 32'h44a2dc6e, 32'hc32fc2b7},
  {32'h42900597, 32'hc20a1a9f, 32'h438bbc29},
  {32'h4502e49b, 32'hc2f1b0a8, 32'hc3b1fb09},
  {32'hc47dedee, 32'h43ceb293, 32'hc21234df},
  {32'h44e9a1d4, 32'h43bb49a1, 32'h42da0b11},
  {32'hc3d11150, 32'hc4df0217, 32'hc322e04d},
  {32'h44c28017, 32'h443cc34e, 32'hc1c66dea},
  {32'hc53f017e, 32'h4343a59a, 32'h43098171},
  {32'h446fc8e0, 32'h44be688b, 32'hc412195f},
  {32'hc4d7597d, 32'hc44b0bf8, 32'hc1c07abe},
  {32'h45055227, 32'hc3f40ce4, 32'h42dd0c99},
  {32'h42552a1d, 32'hc28092a0, 32'h433790db},
  {32'hc2a6c055, 32'hc5235d89, 32'hc3129a2f},
  {32'hc1d751f0, 32'hc43ac98c, 32'h44e3bf87},
  {32'h44a05a4b, 32'hc40a4513, 32'hc218714c},
  {32'h4447b3d0, 32'h4487a4d4, 32'h43d5dac2},
  {32'hc392ddf3, 32'hc37e2597, 32'hc490d819},
  {32'h4509f4f9, 32'h41905bdf, 32'hc307cbfc},
  {32'hc48cb9cc, 32'hc4f47b79, 32'hc4e40590},
  {32'hc378e4b1, 32'h44d729b1, 32'h450f4000},
  {32'h4414870c, 32'h42dbafe8, 32'hc40538dd},
  {32'hc397e10b, 32'h44852716, 32'h4417ad89},
  {32'hc31de8c5, 32'hc3dab010, 32'hc462f509},
  {32'hc301b7f0, 32'h4351f408, 32'h444b5994},
  {32'h435c74e2, 32'hc463edb0, 32'hc4eff3c9},
  {32'h44b1ffc1, 32'hc2ff3b13, 32'h442fdde4},
  {32'h44319fd3, 32'hc4a27451, 32'hc3d998bd},
  {32'h43980dee, 32'h448ded43, 32'h44caa785},
  {32'hc48fce9b, 32'hc485e5be, 32'hc43a7f3e},
  {32'hc4cf517d, 32'h42b70b73, 32'h438f47ef},
  {32'hc0ecd100, 32'hc4d0b946, 32'h43423db8},
  {32'h431aa9d0, 32'h4514ceab, 32'h440d5c63},
  {32'h43aed5c2, 32'hc48885c4, 32'hc3eb9cd2},
  {32'hc3b5cc3b, 32'h456970a5, 32'h43e0fbb6},
  {32'h426745fe, 32'hc532175c, 32'hc1d12370},
  {32'h43d5d206, 32'h4290f2cc, 32'h43e64290},
  {32'hc57a8aeb, 32'hc3f2dd8a, 32'hc3268937},
  {32'h449c9bbd, 32'h409397f8, 32'hc38c5e2e},
  {32'h43d4ccbc, 32'hc43999f9, 32'hc4b55dcc},
  {32'hc441211c, 32'h429c1d18, 32'h43e412a2},
  {32'h438d0c0c, 32'h44425d0a, 32'hc3de3b5d},
  {32'hc3c9fd75, 32'h45157b1c, 32'h42c7a11e},
  {32'h42c0d514, 32'hc5463508, 32'hc18429aa},
  {32'hc2fa2c60, 32'h43e4ad9a, 32'h440f2e45},
  {32'hc40cbe7d, 32'hc3028829, 32'hc472e8c1},
  {32'hc3eca056, 32'h44cb4f19, 32'h44d9b774},
  {32'h440a571b, 32'hc3820d47, 32'hc4965289},
  {32'h4371ffac, 32'hc357b517, 32'h44fc9f06},
  {32'hc3a8a151, 32'h44e1a177, 32'hc4f9a16e},
  {32'hc2b047b7, 32'hc49d670d, 32'h438bec85},
  {32'h431a0857, 32'hc3674619, 32'hc4c808be},
  {32'hc4a392f4, 32'h4490fbfc, 32'h43b7563b},
  {32'h427f7a50, 32'hc3f8f89b, 32'hc3741ece},
  {32'hc35a7740, 32'h4323b44a, 32'h44e4db17},
  {32'h45151fb6, 32'hc2ed8f14, 32'hc38713a6},
  {32'hc31ef108, 32'h431ab1eb, 32'h43d17be4},
  {32'h4405a58a, 32'hc4a56303, 32'hc33506c1},
  {32'hc5214c14, 32'h442ce37c, 32'hc38115e1},
  {32'h44de817f, 32'hc02f5fe9, 32'hc3abafd8},
  {32'hc42ca29b, 32'h42b6ceee, 32'h440b63f3},
  {32'h444af904, 32'hc4a3aa97, 32'hc21104d6},
  {32'hc376dadd, 32'h44df54d4, 32'h42092917},
  {32'h452ee56b, 32'h440a498c, 32'h42b090e3},
  {32'hc516a2be, 32'h437fa54d, 32'h443be279},
  {32'h45244955, 32'h41772f07, 32'hc3088a15},
  {32'h44485640, 32'h43abda37, 32'h443b78ea},
  {32'hc4de7d5d, 32'h436dc0b2, 32'hc42dad97},
  {32'h445379ac, 32'hc341a186, 32'h453ef24a},
  {32'h447e1527, 32'h42abd0f2, 32'h44116eea},
  {32'h4508674c, 32'h43b029e0, 32'h42dd0b39},
  {32'hc4ee25de, 32'h447f808b, 32'h43cd751c},
  {32'h44cc90e1, 32'h43b1677d, 32'h43a4d10a},
  {32'h43327154, 32'h4572d033, 32'h4319ae35},
  {32'h4444b3dc, 32'hc4ef37c8, 32'h42e68d73},
  {32'h448436d0, 32'hc3adffe8, 32'h44234f65},
  {32'h44b0032a, 32'h428e0171, 32'h446d5dd5},
  {32'hc3c7552e, 32'hc3b561dc, 32'hc4fb31e4},
  {32'hc26d3af0, 32'h41fc9301, 32'h430b837c},
  {32'hc3c45a4f, 32'h42a73be3, 32'h447d77ca},
  {32'h436f3d7c, 32'hc412c358, 32'hc4ada33a},
  {32'h4428346c, 32'h43fdb4a5, 32'hc32aa4f7},
  {32'h440f123e, 32'hc45542e5, 32'hc497c639},
  {32'hc2e15702, 32'h45051d35, 32'h40ded1f1},
  {32'hc48b616b, 32'hc2e08964, 32'h41ce7a3a},
  {32'hc58ba4f7, 32'h41a3ff44, 32'hc399d87f},
  {32'hc31f3020, 32'hc4973612, 32'hc4a7d59f},
  {32'h43ba6c55, 32'h4410ad8c, 32'h4474be56},
  {32'h44695076, 32'hc49b767b, 32'hc491a8db},
  {32'hc4602b67, 32'hc034c99b, 32'h4439e100},
  {32'hc4d3bcff, 32'h4204dbfc, 32'hc3345376},
  {32'hc4764ab8, 32'h442502bd, 32'h44cfb950},
  {32'hc2175fcc, 32'hc509752d, 32'hc400a9a1},
  {32'h447682ac, 32'h43f7e9e4, 32'hc4a8437c},
  {32'hc5621147, 32'hc28f3219, 32'h43517c5b},
  {32'h4541c154, 32'h435f7322, 32'hc17bf744},
  {32'h415f9d60, 32'hc45765d9, 32'h42745bf7},
  {32'h44202f1f, 32'h44b74b29, 32'hc32e32ac},
  {32'hc540343f, 32'hc349b0c6, 32'hc34b51ed},
  {32'h42ffa620, 32'h448a7a34, 32'h435d6856},
  {32'hc317a0ec, 32'hc560afb4, 32'h43aa7d70},
  {32'h44b4db00, 32'h437788b8, 32'h43d63bd0},
  {32'hc4bea40f, 32'h4399fe94, 32'h44002e19},
  {32'h4485d841, 32'hc3be4546, 32'h43ba0b4b},
  {32'hc5077c47, 32'hc0d3f548, 32'h4328c871},
  {32'h44ef0a9a, 32'h43d9b0d3, 32'h43ed66ac},
  {32'hc532f31b, 32'hc3c1ba0a, 32'hc3d4aa21},
  {32'hc4a3d11c, 32'h43043386, 32'h43815e76},
  {32'hc3e68d32, 32'h4303070b, 32'hc5049cd6},
  {32'h43ee301f, 32'h451bbf04, 32'h4433f50d},
  {32'hc496e759, 32'hc434a802, 32'hc3c17d8b},
  {32'h45463dd6, 32'hc392f8b3, 32'h43643f7b},
  {32'hc4f033e0, 32'hc3f84ad2, 32'hc480206b},
  {32'hc4bf6b98, 32'hc33196bb, 32'h4243e704},
  {32'hc5222577, 32'hc3de3d01, 32'hc32d4f74},
  {32'h442d8d0f, 32'hc361d93c, 32'h44d45f89},
  {32'hc3412240, 32'h4323fa34, 32'hc38c1384},
  {32'h44f0ea68, 32'h43db0790, 32'h4432a426},
  {32'hc4b5bb0f, 32'hc48ac104, 32'hc430f98a},
  {32'hc448dfd3, 32'hc052c040, 32'hc303f945},
  {32'h452172b7, 32'hc3d16be5, 32'h427568d6},
  {32'h4348b5bc, 32'hc50bc4eb, 32'hc27efa61},
  {32'h440a8e4d, 32'h44f0a350, 32'h43372171},
  {32'hc546270b, 32'h43e1d849, 32'h43badc9b},
  {32'h454bca9c, 32'h4392c3b4, 32'h42f36137},
  {32'hc4fc24e8, 32'hc46bbf48, 32'h433c1d6e},
  {32'h44451357, 32'hc34090a9, 32'hc465f063},
  {32'hc540ce9e, 32'h43add4b0, 32'hc302d9c5},
  {32'h44c22eb6, 32'h41c790b3, 32'h44055320},
  {32'hc49a97b4, 32'hc2e22893, 32'h4319b2d8},
  {32'h451a9a6f, 32'h4323d951, 32'h4330375f},
  {32'hc4572379, 32'hc32ec4da, 32'h438c3fd2},
  {32'h444d19aa, 32'h4489892f, 32'h419e0ac0},
  {32'hc4acaf12, 32'hc303d48f, 32'h43f589d7},
  {32'h44fc5f84, 32'h43ad709f, 32'hc3df9005},
  {32'hc50594bb, 32'hc0cf1a8e, 32'hc3d72d1a},
  {32'h42631600, 32'hc3b5f169, 32'hc49b3439},
  {32'hc518704d, 32'hc2d57a28, 32'hc221719c},
  {32'h4393e373, 32'h44a4faf4, 32'hc2d8effe},
  {32'hc493b472, 32'hc4a9272d, 32'h4506d804},
  {32'h43a9c2e9, 32'h446ca151, 32'hc4c14bf8},
  {32'hc3dab625, 32'hc4efc632, 32'hc44f5f11},
  {32'hc3b1bd60, 32'h4524ec3d, 32'hc39f8cc4},
  {32'hc440f5a0, 32'hc42016d8, 32'h438c22ff},
  {32'hc36a0b64, 32'h43acfb66, 32'hc257c9c8},
  {32'hc49f02a8, 32'h433a7c22, 32'h44796c3b},
  {32'h43a274ef, 32'h4367289c, 32'hc5299e0a},
  {32'hc3cb6fb8, 32'h43e53e00, 32'hc4c04924},
  {32'hc4a2f9fc, 32'h44c1ceea, 32'h41e5aa8e},
  {32'hc4c27309, 32'h43aa1d16, 32'hc2caa3e1},
  {32'hc3322fe0, 32'h44cdd545, 32'hc2f30895},
  {32'h44d0f044, 32'hc41231a3, 32'hc3b0aaac},
  {32'hc47dfc1c, 32'h447442c4, 32'hc309e038},
  {32'h454063c3, 32'h41dee66b, 32'hc19accc8},
  {32'hc562c7a9, 32'h43c50647, 32'hc3dc143d},
  {32'hc32fcd2f, 32'hc3390ec2, 32'h443da574},
  {32'hc39f6b3a, 32'hc3ad53a3, 32'h4471b8fc},
  {32'h4217e240, 32'hc491c549, 32'h43e0b59b},
  {32'h43d79734, 32'hc1dd4501, 32'h4416ef3a},
  {32'h44b05996, 32'h4350eaa1, 32'h444665f2},
  {32'h43300970, 32'h44896f48, 32'hc420776d},
  {32'h44509d97, 32'hc4121bca, 32'h44039b4f},
  {32'hc3c8928b, 32'hc3415f48, 32'hc5037750},
  {32'h45453faa, 32'h42c2f2d7, 32'hc27655a4},
  {32'h44d8480d, 32'hc3960a59, 32'hc3836ae9},
  {32'h44e4cf16, 32'hc4813eb7, 32'h439711ed},
  {32'hc4b5d604, 32'h44b938d0, 32'hc420c2a4},
  {32'h44684e9d, 32'h43a9cf93, 32'hc319aa8c},
  {32'hc39729c8, 32'h452018a0, 32'hc26d1f27},
  {32'h453b4e09, 32'h43f38ebf, 32'h44148eca},
  {32'h43e7849b, 32'h44c7ecfa, 32'h43f6b067},
  {32'h443f8828, 32'h43c0bdb4, 32'h44bd412b},
  {32'hc4638b6d, 32'hc276f0e1, 32'hc45dcd5e},
  {32'h4506503f, 32'hc3f0c231, 32'hc2a8e2a0},
  {32'h4303fe00, 32'h43236bec, 32'hc5220ea9},
  {32'h44a69696, 32'h4440814c, 32'h44700760},
  {32'h43a698ab, 32'h4474e050, 32'hc4373df4},
  {32'h44d1a84c, 32'h43a16eff, 32'hc31b6705},
  {32'hc24abb58, 32'hc4fc3bc7, 32'h43ab5f7a},
  {32'hc4d482f3, 32'hc2bc8dda, 32'hc3f5004b},
  {32'h44050db9, 32'h431edeb6, 32'h4294b644},
  {32'hc499b70e, 32'h442b6d70, 32'hc49a3b23},
  {32'h451bb45b, 32'hc472e53a, 32'h4447bb88},
  {32'h446cdc4e, 32'h4387e561, 32'h4440f44e},
  {32'h433992e4, 32'hc3731bc3, 32'hc5389b62},
  {32'hc4681604, 32'hc458a8e9, 32'h44329a01},
  {32'h4342faa0, 32'hc4ef74ac, 32'hbf7dd780},
  {32'hc4c6e085, 32'h432b3dba, 32'hc411db51},
  {32'hc2e03990, 32'hc520d917, 32'hc354f44e},
  {32'hc4d56660, 32'h440a9be5, 32'h442b5b19},
  {32'hc2bd7878, 32'hc51ec00d, 32'h42a6c0bc},
  {32'hc4c3dfd5, 32'hc2ae3540, 32'hc40c4409},
  {32'h451a56a1, 32'hc4335794, 32'h43e26477},
  {32'hc5254b68, 32'h431de6c0, 32'hc4523b4c},
  {32'h4502790c, 32'h44070c75, 32'h42c30987},
  {32'hc4d3f93e, 32'h43b40a4f, 32'h43b9a617},
  {32'hc29b4442, 32'hc560abf6, 32'hc401a203},
  {32'hc494af16, 32'h44b2637c, 32'hc3ce5bf9},
  {32'h446b291c, 32'hc0499b7b, 32'hc3910316},
  {32'hc4c79630, 32'h44e09c41, 32'h43a8d8c8},
  {32'hc2331920, 32'hc4fbd126, 32'h43fb2a91},
  {32'h4410ebb8, 32'hc3826085, 32'h44acf6a4},
  {32'h449824a6, 32'hc3f6eda2, 32'hc38f2e49},
  {32'hc49c84aa, 32'h444a4ce9, 32'h43dfcb91},
  {32'h43a117b4, 32'hc50b4b59, 32'hc215dae3},
  {32'hc3606098, 32'h450c2afb, 32'hc2977348},
  {32'hc4b1f906, 32'hc42d00a8, 32'h41fd2ec1},
  {32'hc18970b6, 32'h44b5f117, 32'hc516a903},
  {32'hc52b6b56, 32'hc3800540, 32'hc2cab41c},
  {32'h44a80141, 32'h442d5574, 32'h42aeba1d},
  {32'hc392b4bc, 32'h405fc0f2, 32'hc40b90d0},
  {32'hc45dddc4, 32'h4493892b, 32'h446e94b0},
  {32'hc3b3f561, 32'h444847d8, 32'hc53d4bef},
  {32'hc291a80a, 32'hc38f3304, 32'hc51fe83b},
  {32'hc43331f0, 32'hc42f3c79, 32'h44906510},
  {32'h43ed56c3, 32'h44a4de8c, 32'hc41470b4},
  {32'hc4202f59, 32'hc50b2640, 32'hc2b70d33},
  {32'h44f5d7e4, 32'h43487b92, 32'hc3cf96b2},
  {32'h442c2fa8, 32'hc42b06e1, 32'h435d8925},
  {32'h45456b82, 32'hc3bc88b0, 32'h42e24567},
  {32'hc51bcf69, 32'h404d9134, 32'hc2ead2e4},
  {32'hc4af6c36, 32'h43a16b75, 32'hc30636e0},
  {32'hc561b8d8, 32'hc271df90, 32'hc36f3c04},
  {32'h43e5fe3a, 32'h450a2469, 32'hc305b1dc},
  {32'hc4517100, 32'hc3113bbe, 32'hbf6abb00},
  {32'h4483fb43, 32'h446953dd, 32'hc3ec449c},
  {32'hc50ce857, 32'hc4867461, 32'h440d685b},
  {32'h42e8d579, 32'h446fa334, 32'hc38e80ad},
  {32'h440dbe30, 32'hc45075c9, 32'h43b39922},
  {32'hc41b4e10, 32'hc48b142e, 32'hc3eb6dbe},
  {32'hc3c1b0e8, 32'hc50e0bc6, 32'h44a5a989},
  {32'hc3991b26, 32'h426b5147, 32'hc3bf55d8},
  {32'h44230992, 32'h44b4e468, 32'h44607ade},
  {32'hc4cb072c, 32'h4116de14, 32'hc46a7668},
  {32'hc48d6a51, 32'hc392a88e, 32'h4380ee49},
  {32'hc3e2cfbc, 32'hc4185ab1, 32'hc50fe4a5},
  {32'h449f5c4e, 32'h4301f2d8, 32'h44ba3df1},
  {32'h433446b6, 32'hc4af43ec, 32'hc3177671},
  {32'hc48504b4, 32'hc451bad5, 32'h452b99dd},
  {32'hc47cc852, 32'h4327582d, 32'hc30724b8},
  {32'h45155cc0, 32'h42dc146c, 32'h436481c3},
  {32'hc460d8da, 32'hc44627b7, 32'hc3cc57a7},
  {32'h42f13008, 32'h439dd921, 32'h450d6d3c},
  {32'h44651190, 32'hc2a998b9, 32'h43282aad},
  {32'h44b14f52, 32'h4480ba91, 32'h443e38ff},
  {32'hc4b97b2b, 32'hc40eafff, 32'hc3c37051},
  {32'hc4067bc9, 32'hc1a64e16, 32'h43fa89c0},
  {32'h42fbbe90, 32'hc5394d2c, 32'hc2e70894},
  {32'h4401e376, 32'h453a1c22, 32'h43b8c398},
  {32'hc48425c4, 32'h437e0ff2, 32'hc33bdec2},
  {32'h4469fa34, 32'h438368e5, 32'h423e6fc4},
  {32'hc41a320b, 32'hc52b5fb0, 32'hc30a6a90},
  {32'h456b17ee, 32'h4431306f, 32'h434e3185},
  {32'hc55f24ff, 32'hc218c112, 32'h420e7332},
  {32'h44259ab4, 32'h439da81e, 32'h442231f0},
  {32'h434e1628, 32'hc4a0f8d7, 32'h43c61fb2},
  {32'hc322c068, 32'h4508c956, 32'h43e5db93},
  {32'hc12e5e50, 32'h43e6eb9d, 32'hc435428a},
  {32'hc5012131, 32'h431660e6, 32'h431c0d9c},
  {32'h418b1a9c, 32'hc4499423, 32'hc471a34f},
  {32'h4432c182, 32'h42e672f2, 32'h44cbff22},
  {32'hc38fe284, 32'hc4337e08, 32'hc5142d39},
  {32'hc48be052, 32'h4327d100, 32'h44d0acc9},
  {32'h453ed056, 32'h43a69891, 32'h439dd2ec},
  {32'h436a5308, 32'hc4a26e4a, 32'h44e69185},
  {32'h43fb43f0, 32'h448662ca, 32'hc48eabb0},
  {32'hc3b9b908, 32'h43f22ad1, 32'h442c90d6},
  {32'h452bd130, 32'h435ff93a, 32'hc3330d2c},
  {32'hc4ad7137, 32'hc3329b03, 32'h44c605f2},
  {32'hc4ed902f, 32'hbfa6eb80, 32'hc2cb0b72},
  {32'hc35cc754, 32'h4496e8d4, 32'h454393bb},
  {32'hc3ad0635, 32'hc4720fa3, 32'hc4cd3f9c},
  {32'h42014d44, 32'h4320f5de, 32'h44e113e9},
  {32'h43f0e5f8, 32'hc50e2e31, 32'hc36443a2},
  {32'hc45ec2cd, 32'h449fe50a, 32'hc33c5d10},
  {32'h44739061, 32'h4396cd7e, 32'hc3634ea8},
  {32'hc4db5aba, 32'h445e8f96, 32'hc2ebd026},
  {32'h4521dd90, 32'hc392afa8, 32'h42ccbdb7},
  {32'h44706ab6, 32'hc3e1f0be, 32'hc218f840},
  {32'h4494c11c, 32'h44206498, 32'hc3b170e9},
  {32'hc578203e, 32'hc2874be1, 32'hc3d61be1},
  {32'h458b5ed9, 32'h43a3afa1, 32'hc36ae338},
  {32'h454e45a6, 32'h42cc45a9, 32'hc4387c92},
  {32'hc4ad6f90, 32'h41652e88, 32'hc470c382},
  {32'h4470f3e6, 32'hc30fd8fc, 32'h450f2989},
  {32'hc45b9062, 32'h41fda57d, 32'hc4076a48},
  {32'h44ebe026, 32'hc40db8c1, 32'h4361a169},
  {32'hc41c287a, 32'h44ee69df, 32'h428d1d1d},
  {32'h44abc5c0, 32'hc1817dc8, 32'hc37fff19},
  {32'hc48d1859, 32'h44f8da02, 32'hc282d648},
  {32'h4320fe7c, 32'hc577e30e, 32'hc360ccf3},
  {32'hc4f2170c, 32'h439aaa49, 32'hc385dec9},
  {32'h4537b150, 32'h4291f008, 32'h4301dada},
  {32'hc4d9f518, 32'h434bf239, 32'hc3a39240},
  {32'h44450bec, 32'hc3c794d6, 32'hc3ab8d10},
  {32'hc2ecbef5, 32'h44c1861f, 32'h4472f7f7},
  {32'hc3ac1874, 32'hc4e3ff09, 32'hc435c2e7},
  {32'hc2f3f1d0, 32'hc329fd0c, 32'h4390fb37},
  {32'hc30f7b10, 32'hc41e0c4f, 32'hc4531927},
  {32'hc39f779f, 32'h44cb7957, 32'hc3501cc0},
  {32'h4505071b, 32'h43c95a37, 32'h427c2506},
  {32'hc56e809c, 32'hc332744f, 32'hc250bbd6},
  {32'h44b1a8a7, 32'hc407bf0c, 32'hc484ecb8},
  {32'hc4ce9272, 32'h41618481, 32'hc3a16130},
  {32'h451b288b, 32'hc35f55ef, 32'hc25fa33f},
  {32'hc3390910, 32'h44b4aea8, 32'h446f0eb8},
  {32'hc418f3c8, 32'hc3c38519, 32'hc487aa72},
  {32'hc39529eb, 32'h450c9642, 32'h4437f6c5},
  {32'h42d223d8, 32'hc4ca0513, 32'hc42b1004},
  {32'h45560f98, 32'hc376c8e7, 32'hc414517b},
  {32'hc407e5bc, 32'hc2d34b3c, 32'h450235a8},
  {32'hc4a30dda, 32'h43a2cc09, 32'hc399a56d},
  {32'hc4b5f88b, 32'hc4ad13be, 32'hc3eb2b0c},
  {32'h44c6ceb7, 32'h437797c9, 32'hc3e9b99d},
  {32'h44cde0bc, 32'hc3a9002f, 32'hc3957afc},
  {32'h44c9d87b, 32'h448c96db, 32'h433b7d58},
  {32'hc572bfdf, 32'hc3119141, 32'hc20607e5},
  {32'h44ff12a8, 32'hc2135d67, 32'h43342315},
  {32'hc32aff7e, 32'h44432bc5, 32'hc4b5a7e6},
  {32'hc31d7349, 32'hc400772a, 32'hc5376f31},
  {32'h44f32806, 32'hc362c5eb, 32'h439952cc},
  {32'h4469210d, 32'h43e4da85, 32'h44c22d1a},
  {32'hc430f240, 32'hc0d4cd38, 32'hc4bf0b0c},
  {32'h4419fa4c, 32'h43d7b59b, 32'h4369677b},
  {32'hc3162e71, 32'hc506e43c, 32'h438eec9a},
  {32'h446bba1f, 32'h444b2063, 32'h440569a9},
  {32'hc1671fb0, 32'hc4bfe177, 32'hc3633b30},
  {32'h450d2020, 32'hc4052b77, 32'h44b266c2},
  {32'hc4c85086, 32'hc41cf027, 32'hc49b1d8a},
  {32'hc3f4d5b5, 32'h43723ed0, 32'h427cb27c},
  {32'h43ba658e, 32'hc380dd14, 32'hc526bacd},
  {32'h4386cbdc, 32'h451b5e32, 32'hc230d827},
  {32'hc463f4e4, 32'h42c63f84, 32'hc487e023},
  {32'h442a94b6, 32'h4341e172, 32'h44e64a62},
  {32'hc4eded0a, 32'hc316ab6a, 32'hc3c20176},
  {32'hc14ebe00, 32'h440b72eb, 32'h4391a623},
  {32'h450cab2d, 32'hc2e0c534, 32'hc3759cc5},
  {32'hc313962d, 32'hc554ab86, 32'hc216bf0d},
  {32'h446f21d8, 32'h43647ea6, 32'h44969a79},
  {32'h435ac2e5, 32'hc48a85c1, 32'h43ad12dd},
  {32'h44897d14, 32'h449d1541, 32'h401658e0},
  {32'h43307b2d, 32'hc585aa2d, 32'hc204314a},
  {32'h4488a4ed, 32'h43d899e5, 32'h432e9a9c},
  {32'hc4326126, 32'h43a8761b, 32'h421b86c7},
  {32'h44f182a4, 32'h440c8a3b, 32'h448594a2},
  {32'h440452f8, 32'hc45cc58f, 32'h40841f68},
  {32'h43fc0aa4, 32'h44b3f404, 32'h43f016d4},
  {32'h416b3c70, 32'hc40825e6, 32'h4442e91a},
  {32'hc3cde758, 32'hc39f0a6a, 32'hc3f47d49},
  {32'h42b6ade8, 32'hc495ff3e, 32'h44373e9b},
  {32'h44ad31a6, 32'h4432ddae, 32'hc480f495},
  {32'h4408cb53, 32'hc3565b3e, 32'h4447567b},
  {32'h44fe3c13, 32'h4132e2e8, 32'hc3d12790},
  {32'hc4250d5f, 32'hc1863adc, 32'h44a7f1e6},
  {32'h44a472c2, 32'h428ec122, 32'hc47c8e6d},
  {32'hc5120525, 32'hc3eb257a, 32'hc33611f6},
  {32'h41d26f80, 32'h4525b77a, 32'hc41261be},
  {32'h44391a58, 32'hc4b21a38, 32'h42c014c6},
  {32'hc3158c3a, 32'h44e46ab5, 32'hc3fc4495},
  {32'hc49e981c, 32'hc31cb8f5, 32'h448b57ae},
  {32'h455c0298, 32'h440c311b, 32'h433b7a7d},
  {32'hc501f9fb, 32'h43a9898b, 32'h44650b94},
  {32'h450f607d, 32'hc371c64d, 32'hc4a203ee},
  {32'h4516406e, 32'hc481c968, 32'hc314981e},
  {32'hc4711ff2, 32'h44cbb7c2, 32'h43900a16},
  {32'h44d4c2f1, 32'h42395063, 32'h4424d4b0},
  {32'hc4fcf4ec, 32'h445e5e90, 32'hc3cc799f},
  {32'h44e55912, 32'hc4733744, 32'h44140f64},
  {32'hc124be56, 32'h448f42f2, 32'hc34c2f9b},
  {32'h45471fc3, 32'hc410827c, 32'hc438198b},
  {32'hc5830a06, 32'hc3956d11, 32'h43aee9d6},
  {32'h452a6aa9, 32'h42ac15bb, 32'h432f4e9f},
  {32'hc507dc1d, 32'h41bc7ba2, 32'h442bdae8},
  {32'h43c37000, 32'hc3cae7d9, 32'h43e38ad8},
  {32'h44cb1907, 32'h41417e69, 32'hc31146dc},
  {32'h43d201ac, 32'hc517cb2e, 32'hc2cec5db},
  {32'hc36c6b64, 32'h431bb787, 32'hc3cb95dc},
  {32'hc4c55892, 32'h430e9c33, 32'h43b4778a},
  {32'hc527c938, 32'h416617f0, 32'hc43662cd},
  {32'h453761e3, 32'h43bb6faf, 32'hc3ca11fb},
  {32'h4310ee36, 32'h42f1bc85, 32'hc47ee778},
  {32'hc25342e8, 32'hc4f0cfd1, 32'h44328e3e},
  {32'hc3686e30, 32'h4554ea2b, 32'hc3c2e177},
  {32'h42bc0aee, 32'hc48c874a, 32'h42775a56},
  {32'hc528dfc0, 32'h4391f9ec, 32'hc2cfb136},
  {32'hc2144bc6, 32'hc548d72e, 32'hc31c42cf},
  {32'h44838b83, 32'h434a6d1f, 32'hc48b93e3},
  {32'h449ff167, 32'h443415b9, 32'h45455fc0},
  {32'hc3087238, 32'hc3e221f7, 32'hc42d971b},
  {32'h448e3248, 32'hc3ce712c, 32'h439b0a35},
  {32'h4319e697, 32'h44830cf6, 32'hc51f9e60},
  {32'hc2b930f8, 32'h44b0b410, 32'h44a945a3},
  {32'h43b4a670, 32'h447ca03b, 32'hc4a84a85},
  {32'hc4404239, 32'h44842eb0, 32'h4373adca},
  {32'hc093eb80, 32'hc52e6170, 32'hc183dae9},
  {32'hc39e38d0, 32'h443031d5, 32'hc4878344},
  {32'h440f2374, 32'hc4120169, 32'hc367013c},
  {32'hc425a5ba, 32'h44128bca, 32'hc48bd9fc},
  {32'h4367cde0, 32'hc43c7da7, 32'h44be9ca4},
  {32'hc31481b8, 32'hc4405a82, 32'h45391164},
  {32'h42ca5614, 32'h441e391c, 32'hc4e3cb8a},
  {32'hc3b5c019, 32'h4400e134, 32'h44a025c3},
  {32'h44e4704f, 32'hc2f4cbce, 32'h435eb519},
  {32'hc30ef168, 32'h43af1dc5, 32'hc4e8b221},
  {32'h445c7c9d, 32'hc0114db8, 32'h44a2d22f},
  {32'hc4bca5e4, 32'hc2e15a0a, 32'h42d7d086},
  {32'h44a11635, 32'hc39cce34, 32'h444a8085},
  {32'hc53aaa6e, 32'hc2992462, 32'h41e21a0c},
  {32'h44681244, 32'hc3bf79d2, 32'h4369dbe4},
  {32'hc5037d14, 32'h430aaf0a, 32'h43de94a7},
  {32'h43868273, 32'h43b7c578, 32'h43b06e93},
  {32'hc32d1a08, 32'hc20110f4, 32'hc2eec36b},
  {32'h455c3f9d, 32'h439ef570, 32'h43896c74},
  {32'hc48908b8, 32'h445972e4, 32'h43202fc8},
  {32'h43f67c29, 32'hc50fb571, 32'h438d92cf},
  {32'hc5311240, 32'h4421fe8e, 32'hc1dafeb3},
  {32'hc3da7ccc, 32'hc579d546, 32'hc158d220},
  {32'h447c6710, 32'hc3db4ef4, 32'h4325af2c},
  {32'hc2d226d4, 32'h443c424c, 32'hc494dfeb},
  {32'hc49cb1df, 32'h4444d40e, 32'h44786f0e},
  {32'hc43bad22, 32'hc4e806b7, 32'h43950d4d},
  {32'h416a2ee0, 32'h44c4bf76, 32'hc33987bd},
  {32'hc4059a92, 32'hc38342d7, 32'hc38956ce},
  {32'h4500be8c, 32'h42eb8165, 32'hc355e5c0},
  {32'hc4438e8a, 32'hc4b6b16d, 32'h44964fc6},
  {32'hc4b2012e, 32'h44056ff6, 32'h41d8a774},
  {32'hc3fcc87c, 32'h42a5bd34, 32'hc409611c},
  {32'hc3bd96bc, 32'h4370159b, 32'hc330a575},
  {32'hc3a863eb, 32'h44b79a88, 32'hc4ec3009},
  {32'h44162096, 32'hc349d845, 32'hc4c08eac},
  {32'hc5236aba, 32'hc343ad19, 32'hc3772c46},
  {32'hc33e4234, 32'hc3802624, 32'hc3be92fc},
  {32'hc44d2abc, 32'hc484c5e3, 32'h434597fb},
  {32'hc2a7507e, 32'hc34d8b22, 32'hc49ed2f1},
  {32'hbdcaa500, 32'hc3dfe04e, 32'h44f2d74b},
  {32'h450f52e6, 32'h440ce583, 32'hc337c26c},
  {32'hc5619d24, 32'hc305d24b, 32'h43f8423b},
  {32'h44decbe8, 32'hc3a1ded4, 32'h436461b8},
  {32'hc46eb97e, 32'hc4c94d5d, 32'h41cc04a3},
  {32'h449ed3ec, 32'h44068144, 32'h3feeede8},
  {32'h442cf18f, 32'h41d2500d, 32'hc2990b44},
  {32'h44d916aa, 32'h44793667, 32'hc3911bec},
  {32'hc3e7c8de, 32'hc50bcb3c, 32'h43ec6d5d},
  {32'h42a587bb, 32'h436403d4, 32'hc1eeb297},
  {32'hc38acc30, 32'h43a45975, 32'h431a08e0},
  {32'hc4306b1f, 32'h4415daf5, 32'hc453a330},
  {32'hc3992c32, 32'hc50b176e, 32'h44cca088},
  {32'hc4bf4454, 32'h42e2e619, 32'hc33dccd2},
  {32'h44af95e2, 32'h4407adef, 32'h448679bf},
  {32'hc48a87cf, 32'hc2a73811, 32'hc4ab6c2b},
  {32'hc4a45e36, 32'h43199737, 32'h43139bd1},
  {32'hc5022aa6, 32'h431746c0, 32'hc3eb7dfd},
  {32'hc2d3007f, 32'h450b49e0, 32'h44ddedb4},
  {32'h43e3eb70, 32'h44b9d0c2, 32'hc3d8c143},
  {32'hc3418f18, 32'hc4b808c4, 32'h44e31bbe},
  {32'hc35fe2d0, 32'h443599b7, 32'hc4dfa129},
  {32'h430a45d2, 32'h42c3de27, 32'h443161ca},
  {32'hc19e48e2, 32'hc3b5ec02, 32'hc538753e},
  {32'h41a3b8c0, 32'h440320ed, 32'h44f6842f},
  {32'hc3dfd828, 32'hc465d2c6, 32'hc35f5686},
  {32'hc2ac2e40, 32'h43ad477a, 32'h44ba64be},
  {32'hc3374685, 32'hc3fdf64b, 32'hc57de269},
  {32'h450b029e, 32'h422eed38, 32'h4288d0d2},
  {32'hc561ee96, 32'hc327adbe, 32'hc339f7fe},
  {32'h44737a08, 32'h4502fcd4, 32'h43febc35},
  {32'h44b002c8, 32'h4183ec00, 32'h434233c1},
  {32'h43639d93, 32'h4339e23c, 32'h4184b005},
  {32'hc3e150be, 32'hc4aeb85c, 32'hc38a82ae},
  {32'h43ccb1f1, 32'hc385392d, 32'h42d85a9b},
  {32'hc527c510, 32'hc3b31fb2, 32'h43059482},
  {32'h44c6cf36, 32'hc303b293, 32'h4206977b},
  {32'h4383e4b0, 32'h44c332a8, 32'hc4997fb6},
  {32'h4270fec4, 32'h4535b74f, 32'h445cb91f},
  {32'h44eb566e, 32'h43b5edf1, 32'h4331fb27},
  {32'hc40f888a, 32'h44869394, 32'h440070f9},
  {32'hc28ecb00, 32'hc45cb8cd, 32'hc5291370},
  {32'h44112fee, 32'h449eb7a7, 32'hc314c2ae},
  {32'h43c61f9f, 32'hc44f9b83, 32'hc497bc50},
  {32'hc4bc6912, 32'h4449f64d, 32'h43f384d8},
  {32'hc38498a5, 32'hc3fc853c, 32'hc4b9af85},
  {32'h43a36f3d, 32'h4202d50d, 32'h44e2b1fc},
  {32'h4499949c, 32'h43ebf576, 32'hc41a090a},
  {32'hc3ea6e6c, 32'h441fb4cf, 32'hc3c487dc},
  {32'h44536392, 32'hc2f15425, 32'hc441ca2a},
  {32'h4336ea2e, 32'h4363d04b, 32'h42609c29},
  {32'h44c0ecb0, 32'h4332a674, 32'hc22c4cc6},
  {32'hc32fff2e, 32'h3ffebe82, 32'h441b3fc6},
  {32'hc40e729c, 32'hc490d760, 32'hc5398e2b},
  {32'hc443a5cb, 32'h4495c45d, 32'h4331cd2b},
  {32'h44bf3a7c, 32'hc4b79c57, 32'h420f11f4},
  {32'h42570074, 32'h4525c7fe, 32'hc14dc120},
  {32'hc4510517, 32'hc42473c1, 32'h42986ff2},
  {32'hc26daa78, 32'h454a057c, 32'h420d4c6c},
  {32'h452bfa10, 32'hc2b99800, 32'h43782c6d},
  {32'hc4fbbb7c, 32'h434b9e54, 32'h41e66670},
  {32'h449e2756, 32'h43d2d75e, 32'h42a6c56d},
  {32'hc597542c, 32'h41e9e87b, 32'h436a9aea},
  {32'h43ab8806, 32'h43a327ee, 32'hc277966d},
  {32'h43e2ef85, 32'h43f4c026, 32'h4448396f},
  {32'hc5216279, 32'hc0a397e2, 32'hc42abf4a},
  {32'h447ef02e, 32'h43fc8f83, 32'h4472b48a},
  {32'hc4d47903, 32'h43423d1f, 32'h43ae3b39},
  {32'h441827c6, 32'hc51e60c0, 32'hc32cf108},
  {32'hc4c55951, 32'h4488e051, 32'h44126308},
  {32'hc303d7cf, 32'hc4d44b82, 32'h4287b7c2},
  {32'hc57b52e7, 32'hc16cc091, 32'h43391a8d},
  {32'h4405a012, 32'hc514d9b2, 32'h43545c67},
  {32'h43f49df6, 32'h439e509e, 32'hc4d7a707},
  {32'h44135803, 32'hc35277ee, 32'hc2e4c517},
  {32'hc50cdb30, 32'hc3d9f1a7, 32'hc2f82f8e},
  {32'h4496f8b1, 32'hc4074ac9, 32'h434ad458},
  {32'hc3105a74, 32'h4500f943, 32'hc288ccb3},
  {32'h449966b9, 32'hc1b942ac, 32'hc3a785ad},
  {32'h4455bb00, 32'h43b43d79, 32'hc347079c},
  {32'h43b0c7b1, 32'hc47b35e9, 32'hc33d9759},
  {32'hc39a8b98, 32'h44a5a374, 32'h445a54fb},
  {32'hc48c7910, 32'hc41632de, 32'hc3cb80e6},
  {32'hc584bf6b, 32'h43ae8834, 32'h4063b1e0},
  {32'h44d93108, 32'hc3e447d6, 32'hc495ecad},
  {32'hc433291a, 32'h430890aa, 32'hc0c41988},
  {32'h41c47140, 32'h439a6950, 32'hc51e6a74},
  {32'h43dc4d2a, 32'h4521aabc, 32'h44120d8d},
  {32'h43f1167e, 32'hc4346c23, 32'hc422ec07},
  {32'hc25952e0, 32'h45006ec2, 32'h443b3b14},
  {32'h43a4e58c, 32'hc4bb1af0, 32'hc4c372d2},
  {32'h44ed179a, 32'hc28e0399, 32'hc5003ffa},
  {32'hc52a87d7, 32'hc16eb780, 32'h4436236f},
  {32'hc483a704, 32'h42baed12, 32'hc3a008c1},
  {32'hc2486ebe, 32'hc5586f7f, 32'hc39efb88},
  {32'hc3857c57, 32'h4562db90, 32'h436c75a2},
  {32'hc415f85c, 32'h421c5449, 32'hc3133e48},
  {32'h448c5b50, 32'h44156c34, 32'hc40ed6d0},
  {32'hc468aa3c, 32'hc52732ac, 32'hc3f062ad},
  {32'h412c0920, 32'h435856fa, 32'h4432058f},
  {32'hc42d81ad, 32'hc34b0642, 32'h44546baa},
  {32'h44f33e0a, 32'h43dc9760, 32'h43a98af8},
  {32'h442f0d5f, 32'hc4237ade, 32'hc29b2f9a},
  {32'h447deade, 32'h4462a6c8, 32'h4412d3f8},
  {32'hc5367870, 32'hc25f384a, 32'h41dd20d2},
  {32'h44eb959c, 32'h437a7210, 32'hc1d1b7a5},
  {32'hc2fe88c3, 32'hc2d2ce59, 32'hc4d9b04d},
  {32'h4410d5a6, 32'h42a7c694, 32'h45017ab1},
  {32'hc53d8dfd, 32'hc30650f8, 32'h4246c4c0},
  {32'h456a68fe, 32'hc2fd01d3, 32'h434e1279},
  {32'hc533c9d0, 32'hc2fefe5c, 32'hc3c3f2d5},
  {32'h4473b829, 32'hc3ff3363, 32'hc3d977b8},
  {32'hc1dd36f0, 32'hc4c1e215, 32'hc32ac137},
  {32'h42218cb2, 32'h44b075e3, 32'h44134b11},
  {32'h444f3eea, 32'hc0682728, 32'hc43a436b},
  {32'hc3c8ddb0, 32'hc2a9d31a, 32'h44ed0b47},
  {32'hc519ad76, 32'h42830f70, 32'hc3f99e3b},
  {32'h43e36eea, 32'h4465a566, 32'h438f25eb},
  {32'h44a8eaf6, 32'hc3f2b600, 32'hc25db965},
  {32'hc54cfb8f, 32'h43293ebb, 32'h4323128e},
  {32'hc0969700, 32'h4516b8c0, 32'h42f56e38},
  {32'h441fdc46, 32'hc406c52d, 32'hc086c4e5},
  {32'h44d7a2a0, 32'h44873e5c, 32'hc395de29},
  {32'hc45257d4, 32'hc495601d, 32'h434c5a39},
  {32'hc4af9f7c, 32'h4372ff7d, 32'hc2eb350e},
  {32'hc538fdd0, 32'hc34ba8dc, 32'hc313c1ce},
  {32'h441bc8b0, 32'h44450e1a, 32'h44654dd7},
  {32'h44c9f93d, 32'h4454f786, 32'hc3c81e12},
  {32'h44af7b97, 32'h4404ad0c, 32'h437dbc6d},
  {32'hc430851f, 32'hc440bbfc, 32'hc39c210b},
  {32'h4427e7b0, 32'h43e17395, 32'hc255ad4d},
  {32'hc30d6476, 32'hc170d146, 32'h454740d6},
  {32'h446161d9, 32'h435fa622, 32'hc427c822},
  {32'h44b95440, 32'h42fcd962, 32'h43973917},
  {32'h4225941e, 32'hc1cb7a90, 32'hc5442940},
  {32'hc5498df4, 32'hc345070f, 32'h43a9265b},
  {32'h42d455ff, 32'h44d9fa37, 32'h42207bf8},
  {32'hc383b36b, 32'hc487ebb2, 32'hc35638da},
  {32'h43d7e75f, 32'h45146bad, 32'h426c96ca},
  {32'h43beaede, 32'h43997e8b, 32'h447d35b9},
  {32'h44429ebc, 32'h44052fcc, 32'hc3db367c},
  {32'hc4f7b01a, 32'hc48209ac, 32'h438c1ff4},
  {32'h43e63740, 32'hc3847073, 32'hc5054fa4},
  {32'hc43d4f8a, 32'h42f936cd, 32'h44e02051},
  {32'hc3ce1cb0, 32'hc43e71e0, 32'hc35f2a58},
  {32'h41a32a80, 32'hc521c862, 32'hc204fb58},
  {32'h4326b15f, 32'h4558789b, 32'hc1643f67},
  {32'hc468756d, 32'hc476d160, 32'h421acc6d},
  {32'hc380584e, 32'h4549b0f5, 32'hc21b5b2e},
  {32'h44c27445, 32'hc40837c4, 32'hc3bdbdd0},
  {32'h43851092, 32'hc1dac66f, 32'hc38eb2ca},
  {32'h44bdf738, 32'hc3ba505f, 32'hc25474d0},
  {32'hc53f84e0, 32'h44596ef2, 32'hc29471b8},
  {32'h45042fa7, 32'h439ed910, 32'h43af720c},
  {32'hc479c0b2, 32'h4453ae3d, 32'h4404d5f2},
  {32'hc38d600a, 32'hc4d60a9f, 32'h4433a476},
  {32'hc3740fb6, 32'h4484f924, 32'hc3f9f4f5},
  {32'h42c3b1f0, 32'hc407a77e, 32'h44649238},
  {32'hc3f3f280, 32'h4472c693, 32'hc3c31c73},
  {32'hc4a99692, 32'h43f1bb4b, 32'h438c8903},
  {32'hc508d750, 32'h42aed7f2, 32'hc4523aaa},
  {32'h451dfad9, 32'hc443e9ee, 32'hc3a80a18},
  {32'hc40fddef, 32'hc3b7dd4e, 32'hc42b94b1},
  {32'h43b12894, 32'hc565a66b, 32'hc204674a},
  {32'hc57891cc, 32'hc29c57f2, 32'hc3e61b0a},
  {32'h448a7ccd, 32'hc41f122e, 32'h440ee2fa},
  {32'hc4c78a2d, 32'h43327652, 32'hc3f303a4},
  {32'hc3b66524, 32'hc393b2b4, 32'h45105b16},
  {32'h44918534, 32'h44027661, 32'h43e14eef},
  {32'h44314802, 32'h43a19808, 32'h450b0db9},
  {32'hc49e5a6c, 32'hc1ddd6c5, 32'hc4adb87e},
  {32'h44c0020c, 32'h42d02e3d, 32'h44156535},
  {32'hc41e986b, 32'h43f7df18, 32'hc4406be0},
  {32'h448df4ca, 32'h43280f11, 32'h448e3bb7},
  {32'hc3bcb024, 32'h43bbb958, 32'h42b603b6},
  {32'h43dad5f8, 32'h43c953cc, 32'hc41054b7},
  {32'h448e845e, 32'hc4186546, 32'h44b5e3c4},
  {32'hc2b9d3c8, 32'h44ae58d1, 32'hc347ebdc},
  {32'hc44ab1db, 32'hc39ccd02, 32'hc3044812},
  {32'hc3e030fe, 32'h44f5b03c, 32'h423dbece},
  {32'h43c72cd2, 32'hc500f702, 32'h44680c24},
  {32'h444af808, 32'h44a2f675, 32'h44891f5c},
  {32'h43bc5e6e, 32'h436ffb73, 32'hc508aae7},
  {32'h4396d49d, 32'hc3673775, 32'hc3d63ded},
  {32'h4400099e, 32'h44067dcd, 32'h44269cb6},
  {32'hc4a3da20, 32'h4287cabf, 32'h42debdf7},
  {32'h45094216, 32'hc42f16b1, 32'h41eb6eaa},
  {32'h444d24b8, 32'h4490be97, 32'hc210317b},
  {32'h445098c9, 32'hc466da0a, 32'h444c0bd1},
  {32'hc3380760, 32'h43240635, 32'hc47cf723},
  {32'h44f08d64, 32'hc32fe6d6, 32'h44404a23},
  {32'hc584b43b, 32'hc379a55f, 32'h43945f23},
  {32'h4556c74e, 32'h42a24bdc, 32'h43773bfe},
  {32'hc38da354, 32'h429699de, 32'h43c162e9},
  {32'hc0f1cfc0, 32'hc5101b11, 32'hc2d78802},
  {32'hc4f4a0ae, 32'h43b8f9bf, 32'h42b5d55f},
  {32'h443d8b3a, 32'hc43d6d05, 32'h430ae542},
  {32'hc30e8fb2, 32'h453daa6d, 32'h40c40feb},
  {32'h44b24c6d, 32'hc48ef588, 32'hc1e9c859},
  {32'h4433873e, 32'h43203ec4, 32'h44c5ea21},
  {32'hc3d18a40, 32'h44be41c5, 32'hc4b54436},
  {32'hc408549b, 32'h4485728a, 32'h44a3445b},
  {32'hc4070510, 32'hc4aa3a6b, 32'h43aceff7},
  {32'hc32f7390, 32'h4352ccc5, 32'hc527da59},
  {32'h43f5fa4a, 32'hc3c40a1a, 32'h418b9b0a},
  {32'h44f635f3, 32'h43fe4812, 32'hc40c99c8},
  {32'hc53f5607, 32'hc3d367d5, 32'h4384d39a},
  {32'h44a401ad, 32'h43596594, 32'h43a987a3},
  {32'hc47aff70, 32'hc413248a, 32'hc2f5bfdd},
  {32'hc41ed0f8, 32'h43ddd44d, 32'h44d59c2b},
  {32'h4489e5ad, 32'h43ed9573, 32'hc4ae4a9d},
  {32'h444176be, 32'h441659c2, 32'hc43400b6},
  {32'hc5014207, 32'hc4225115, 32'h409ea9cd},
  {32'h44a45a4b, 32'hc2e5c2e4, 32'hc3b93c1a},
  {32'hc406855c, 32'h412e7682, 32'h44d433da},
  {32'h44a0cc7a, 32'h4433e5b7, 32'hc39cd1c4},
  {32'h442b1687, 32'hc39b0c42, 32'h424f8734},
  {32'h440d18f0, 32'hc3f45f84, 32'hc3f7c26c},
  {32'hc513c979, 32'hc2fbffc6, 32'hc353f631},
  {32'h417036bf, 32'h43afbd94, 32'hc31b1905},
  {32'hc48ab163, 32'hc4a0a118, 32'h43d16036},
  {32'h44fc946b, 32'h43824362, 32'hc199c208},
  {32'h44e2187c, 32'hc320fe51, 32'hc308f171},
  {32'h452f51e4, 32'h44587b98, 32'hc320ea2e},
  {32'hc4830952, 32'hc4c9c4b1, 32'hc3b3bdcc},
  {32'hc339f07e, 32'h444a9e01, 32'h432bc14f},
  {32'h43aed0dc, 32'hc4b9a5d0, 32'h4286ab7c},
  {32'hc32431e0, 32'hc47d3a90, 32'hc48e2413},
  {32'h431778b0, 32'h451d3576, 32'hc3743c2c},
  {32'hc50e3168, 32'h430b1ca7, 32'h4334360c},
  {32'h4418b906, 32'h44c45da7, 32'h4470370a},
  {32'hc4850573, 32'hc397a838, 32'hc452addf},
  {32'h44057753, 32'h4433ce12, 32'h43f962c5},
  {32'hc41f8310, 32'hc4514033, 32'hc4907c9c},
  {32'h434fb960, 32'h44c0d67f, 32'h44a10f8f},
  {32'h439d16d4, 32'hc3fad8c2, 32'hc1a03488},
  {32'hc21aed72, 32'hc373c8a9, 32'h43e6e893},
  {32'h441be375, 32'h43cc87ab, 32'hc520561e},
  {32'hc494dab8, 32'h4307394f, 32'h442f6d9f},
  {32'hc272f7f0, 32'hc3fe96e2, 32'hc4d5c9c0},
  {32'h4467e38d, 32'h44a2c49f, 32'hc14e191e},
  {32'hc4b9a54b, 32'hc03228a8, 32'h438f2c47},
  {32'hc3927f36, 32'h44878c1f, 32'h4573676b},
  {32'hc54e9ad4, 32'h418ff4c0, 32'hc3e247fe},
  {32'h406c2840, 32'h44dfa10e, 32'h4368aaeb},
  {32'hc511b2fa, 32'hc4984ced, 32'hc3cbcc39},
  {32'h448127b3, 32'h450be235, 32'h440ee5b4},
  {32'h436a7bcf, 32'hc49e37b6, 32'h43402b28},
  {32'h441aa867, 32'h44ce588e, 32'hc37e32bd},
  {32'hc443c35e, 32'hc49c1d6a, 32'h439b18e1},
  {32'hc4db9212, 32'hc1337495, 32'h42d020e1},
  {32'hc49b22ce, 32'h42ccd049, 32'hc441402c},
  {32'hc31991a0, 32'h43bc0d50, 32'h43be8dcd},
  {32'h433566e0, 32'h42d532d2, 32'hc4e11d52},
  {32'h4379be58, 32'hc3e936e4, 32'h44ac5381},
  {32'h449bb350, 32'h439b8e74, 32'h41d0949c},
  {32'hc2c30430, 32'hc2e73e9c, 32'h4540dd6d},
  {32'h43cb7e46, 32'h417a4fee, 32'hc4f30d84},
  {32'hc516ba06, 32'h41d95358, 32'h4422aa08},
  {32'hc380eb7b, 32'hc35babeb, 32'hc5630430},
  {32'hc51d572e, 32'h4414cbc3, 32'h4415530e},
  {32'hc4bf8d39, 32'hc3c2762e, 32'hc358c57f},
  {32'h43a1b394, 32'hc309a55e, 32'h44154c4c},
  {32'h4394fbde, 32'hc53cb5ae, 32'hc44697a6},
  {32'hc48d89c0, 32'hc3ac1de2, 32'hc2cc7722},
  {32'h43a3125c, 32'hc38053c4, 32'hc5172f8c},
  {32'hc4514180, 32'h444c28f8, 32'h443eb775},
  {32'hc34a9e31, 32'hc3d79d5a, 32'h42e945cb},
  {32'hc4d2439e, 32'h43c18175, 32'h441d33eb},
  {32'hc321fcc6, 32'hc4dfd467, 32'hc4e0d9e1},
  {32'h4416e72f, 32'hc359f0f5, 32'hc373b930},
  {32'h44f55035, 32'hc40c3ee5, 32'hc3f51768},
  {32'hc415dc58, 32'h44e7cbcf, 32'h441b3032},
  {32'hc3a44488, 32'hc4a3bc83, 32'h43967215},
  {32'hc5038c80, 32'h44ad28ea, 32'h43847a49},
  {32'h4497511e, 32'hc4452f80, 32'hc3092d0a},
  {32'hc52ce6c4, 32'hc2702ee6, 32'hc19df5af},
  {32'h4516fd30, 32'h4390a23d, 32'hc3e341a8},
  {32'hc5848580, 32'h43a64329, 32'hc3b0b2a3},
  {32'h4526d1fa, 32'h42b5bb99, 32'hc315dd6a},
  {32'hc35ff17d, 32'h433c618b, 32'hc1779911},
  {32'hc544e512, 32'h4383cefb, 32'h4308806b},
  {32'h4433238a, 32'hc3b321f0, 32'h45161c01},
  {32'hc46693bf, 32'hc30ccfbb, 32'h43822465},
  {32'h45483463, 32'hc3621264, 32'h4395baa9},
  {32'hc3004620, 32'h447d23dd, 32'h4302ba70},
  {32'h44f98e1e, 32'h42c6a927, 32'hc3566bd8},
  {32'hc4ac792e, 32'h44d6c4dd, 32'hc3ab6158},
  {32'h4401bc14, 32'hc458a67b, 32'h440169c3},
  {32'h444ec2fc, 32'hc33dc8f0, 32'hc40dfd16},
  {32'h44a08342, 32'hc4068887, 32'hc37b33b5},
  {32'hc44ded7e, 32'hc36e6973, 32'hc3a101c3},
  {32'hc501dd50, 32'hc2ca2244, 32'h43019cd4},
  {32'hc420c462, 32'h440a0309, 32'h432b9e7c},
  {32'h43a63c2c, 32'hc3daf706, 32'hc51400f5},
  {32'hc405a2f5, 32'h44a0f7d4, 32'h442556b2},
  {32'hc3e515cc, 32'hc45513c7, 32'hc3d956ca},
  {32'hc484cf92, 32'h43c2fcac, 32'h441a685b},
  {32'hc482c1e0, 32'hc3e9ab90, 32'hc3f54e9a},
  {32'hc469c6d0, 32'hc3c16886, 32'h42ab0626},
  {32'h456032f4, 32'h42c3e608, 32'hc441a7ef},
  {32'hc5088031, 32'h43ba29c1, 32'hc2c0d24f},
  {32'hc2b041ac, 32'hc31975be, 32'hc34ecf36},
  {32'hc2f63073, 32'h446abe83, 32'h447351f3},
  {32'hc45ebd54, 32'hc2cb9a86, 32'hc3a0bb08},
  {32'h434bef37, 32'h442e8acb, 32'h4527f4e2},
  {32'h43941da0, 32'hc42171fa, 32'hc5179616},
  {32'h4518efa4, 32'hc31ed822, 32'hc4075a0a},
  {32'hc4405364, 32'hc19ccbba, 32'h450ec0da},
  {32'h446ac460, 32'h438cac2b, 32'h440320fe},
  {32'hc5212ddc, 32'hc3b869fc, 32'h43dc69b6},
  {32'h433570e4, 32'h450a1f63, 32'h42137b7b},
  {32'hc4168b25, 32'hc4af53b7, 32'hc2f6cde5},
  {32'h44b7bcfa, 32'h44eff630, 32'h4300e356},
  {32'hc3d528bc, 32'hc56ba81b, 32'h43ba7327},
  {32'hc2db8933, 32'h45102aa6, 32'h43902565},
  {32'h41723a80, 32'hc41af61d, 32'h44ada901},
  {32'h43cdaf8f, 32'h430cf62e, 32'hc4e22f86},
  {32'h4383527c, 32'hc3c134f0, 32'hc30a1228},
  {32'h4406c146, 32'h43aafaaf, 32'h450646fb},
  {32'hc441f054, 32'hc395715f, 32'hc4f6a4d1},
  {32'h44251bf7, 32'h441e24d7, 32'h43a93936},
  {32'hc295cda0, 32'hc41e5625, 32'hc4506657},
  {32'h43c619a0, 32'h43a00641, 32'h4440a6b6},
  {32'hc48abd1a, 32'hc4500910, 32'hc0197ec2},
  {32'h456bf008, 32'h44163ed6, 32'h43f47578},
  {32'hc52cf20b, 32'h430524c3, 32'hc3d2252b},
  {32'h4540369d, 32'h42dc0292, 32'hc3823a6a},
  {32'hc397059d, 32'hc5153993, 32'hc4756fa6},
  {32'h44a5a274, 32'h44125148, 32'h425176f8},
  {32'hc5004686, 32'hc2e08fd8, 32'h43863b52},
  {32'hc2ac37bf, 32'h4362ffdd, 32'h44a0d1fb},
  {32'h42dc6499, 32'hc50856a3, 32'hc481fff3},
  {32'h453cab73, 32'hc307b1a5, 32'hc41e97b1},
  {32'hc3991912, 32'h431f9192, 32'h4122d976},
  {32'hc296b7ae, 32'hc502454b, 32'h434b3cf2},
  {32'h4406b50e, 32'h441f44b8, 32'h44c8c0b8},
  {32'h43516b84, 32'hc479e647, 32'h438786c2},
  {32'h451c46cc, 32'h438bdb72, 32'hc395e456},
  {32'hc3aab3a9, 32'hc567c6e8, 32'hc3164c22},
  {32'h448274c7, 32'h43cdcb80, 32'h43646709},
  {32'hc4c8b160, 32'hc1c8eeb2, 32'hc38a38af},
  {32'h44e8acfe, 32'h42aa4842, 32'h440f879c},
  {32'h43f66697, 32'h4398b57a, 32'hc2aaef12},
  {32'h4488c84b, 32'h422e2f86, 32'h43708842},
  {32'h42316dd2, 32'hc50846f8, 32'hc222c822},
  {32'h4394f120, 32'h44071637, 32'h42080230},
  {32'hc32cb2f8, 32'hc539f6ab, 32'h4402e191},
  {32'h441c77d1, 32'hc2776a6a, 32'hc23987be},
  {32'hc4c97b77, 32'hc3a0fd82, 32'h429a5b80},
  {32'h4315b7e8, 32'h44400a55, 32'h42dfd3af},
  {32'hc5205bb2, 32'h43d9d537, 32'h4399332c},
  {32'h431093f4, 32'h44d16826, 32'h43184af0},
  {32'hc5093fb0, 32'hc43e8a4f, 32'h431508c6},
  {32'h43ee5b07, 32'h4520a7ec, 32'hc33c2595},
  {32'h43ea46e2, 32'hc345deee, 32'h44b8c40b},
  {32'h4385b92e, 32'h4367b3e3, 32'hc32bb7b9},
  {32'hc4a5252c, 32'hc379fcc4, 32'h44811f23},
  {32'h44e7f583, 32'h42180c51, 32'hc29ea457},
  {32'hc42a8868, 32'hc2c42635, 32'h43f9b3d8},
  {32'h457a0104, 32'h438311e6, 32'hc4174743},
  {32'h4529974d, 32'hc3c22a5a, 32'hc40b668f},
  {32'hc32637b4, 32'h4510f478, 32'h441ba7b8},
  {32'hc3ebae49, 32'hc48c8b40, 32'h436fb4c3},
  {32'h439c5392, 32'h450d1b4b, 32'hc311a957},
  {32'h448fec1e, 32'hc4c49f2f, 32'hc4441cfb},
  {32'hc54d5e64, 32'hc3acefa9, 32'h424ece72},
  {32'h44c49f3a, 32'hc3e0bf7c, 32'hc4151dad},
  {32'hc5441b67, 32'h4436670e, 32'h43a6dc07},
  {32'h449e76b0, 32'h431ca2cc, 32'h43dffaf4},
  {32'hc4db7044, 32'h441539f7, 32'hc490cc86},
  {32'h44e06cfa, 32'hc317a7de, 32'h43a6b38b},
  {32'hc49c3d80, 32'h43c7c9f8, 32'hc3950457},
  {32'h44582e58, 32'hc3280850, 32'h43b70afe},
  {32'h430039e4, 32'hc36bf122, 32'hc4f9a06a},
  {32'h448562b0, 32'hc382937c, 32'h441b76e9},
  {32'hc4d1e1c2, 32'h440dd1b1, 32'h43f5e27c},
  {32'h43cd5742, 32'hc2262f2f, 32'h44fcda26},
  {32'hc41ea808, 32'hc3666039, 32'hc42bc114},
  {32'h451aba6a, 32'hc4286ab4, 32'h42a37970},
  {32'hc4147c76, 32'h446b8752, 32'hc5388c16},
  {32'hc4f3c461, 32'hc200c300, 32'h413e68fe},
  {32'hc34c068f, 32'h43fb664c, 32'hc50729be},
  {32'h4441d710, 32'hc4982236, 32'h437d828c},
  {32'hc54fa080, 32'h3facbdc0, 32'h43e348ab},
  {32'h44c77d80, 32'h42e76cf4, 32'h441a22a5},
  {32'hc418a10c, 32'hc300ee50, 32'hc5627211},
  {32'hc4b079b5, 32'hc40347bd, 32'hc347b0b6},
  {32'hc2b0bc78, 32'hc4a8ead1, 32'hc5372152},
  {32'h43ac181d, 32'h43b16d0c, 32'h43d6cdde},
  {32'h4414e262, 32'h4460309c, 32'hc3f73749},
  {32'hc06f6440, 32'h42bb9192, 32'hc285159f},
  {32'h44b2979f, 32'hc38daddc, 32'h44c822f2},
  {32'hc4601e82, 32'h448e8942, 32'h4396ac87},
  {32'h4405a054, 32'h438043ac, 32'h44aa4742},
  {32'hc41bfc91, 32'h44ae5333, 32'h42996e24},
  {32'h44825e90, 32'hc2e3d8f8, 32'h443db292},
  {32'h44ece9ec, 32'h44152162, 32'h44a25bc3},
  {32'hc49903fa, 32'h44b29dd2, 32'hc466a843},
  {32'h4413b6b7, 32'hc488d9c7, 32'h43832e3b},
  {32'h44b85832, 32'hc289dd2e, 32'hc2bbf8d3},
  {32'hc32f273e, 32'h44b4e4ef, 32'hc3e37062},
  {32'h448e4954, 32'hc33c07d8, 32'hc174e326},
  {32'hc362655b, 32'h440b0861, 32'h43df8baa},
  {32'h44047e62, 32'h42b747d6, 32'h450a4fe7},
  {32'h433cde5e, 32'h44bb68eb, 32'hc42a71e7},
  {32'h453f0e0c, 32'hc30c6936, 32'h439af558},
  {32'hc4362570, 32'hc40a09ed, 32'hc4233e19},
  {32'h456a8a34, 32'hc357e33d, 32'h441194a7},
  {32'h4410fc42, 32'h448086a2, 32'h4404d48c},
  {32'h44bcfa00, 32'hc339756c, 32'hc3ebb959},
  {32'hc4101c84, 32'hc23d8e10, 32'h43136c18},
  {32'hc496e4cd, 32'hc31eb5ab, 32'hc38b832c},
  {32'hc4234fef, 32'h4510273e, 32'hc3988903},
  {32'h443bc7b8, 32'hc4e719ab, 32'hc28bb27d},
  {32'h4513bf3a, 32'hc39465dd, 32'h4378d492},
  {32'h42a106a0, 32'h43ab6859, 32'hc4ed8b9a},
  {32'hc3f6d688, 32'hc4cbe680, 32'h44ddd9f0},
  {32'hc4c67c1d, 32'hc3de1537, 32'h44128595},
  {32'h44df766e, 32'hc32bf2a6, 32'hc45becd6},
  {32'hc422e518, 32'hc3e9f11c, 32'h443759ac},
  {32'h4503870e, 32'h44907039, 32'h42f660b8},
  {32'hc4ce1157, 32'hc475263f, 32'h42b846ef},
  {32'hc3b4c168, 32'h44217c14, 32'h431d8796},
  {32'h43eede20, 32'h44d2fb19, 32'hc419282c},
  {32'hc4f1d5ba, 32'h444e15f1, 32'h4480afb9},
  {32'h444b1047, 32'h43f86222, 32'hc49dfdc0},
  {32'h44eebbea, 32'h443e2165, 32'hc30fcc8e},
  {32'hc3fe0c3d, 32'hc416f28c, 32'h44e130f3},
  {32'hc4c5161a, 32'h4284e0ae, 32'hc38e935b},
  {32'hc4c8907c, 32'hc406d6f7, 32'h43a3fd22},
  {32'hc379491c, 32'hc3bc8e01, 32'hc57c0546},
  {32'hc413bbad, 32'hc4538f0b, 32'h43f154f3},
  {32'h44aa7989, 32'hc33e61c7, 32'hc31c2fbe},
  {32'hc56eebf6, 32'hc37cf5ca, 32'hc1eb91e1},
  {32'h44b5ca88, 32'hc0ed6b38, 32'hc3420f21},
  {32'hc403b0ac, 32'hc48cdaa3, 32'h42c56452},
  {32'h44add30e, 32'h448cd3ec, 32'h43bdef8c},
  {32'h44a17e3b, 32'hc408854a, 32'h43a85e02},
  {32'h44a63688, 32'h44de5e06, 32'hc3d1c26c},
  {32'hc49aab00, 32'hc471c471, 32'h4335ee94},
  {32'h445a694a, 32'h435b9ff2, 32'hc349a9a1},
  {32'hc2ecbe3c, 32'h4462ab3e, 32'h4436ad6c},
  {32'hc35e1c76, 32'hc50cfd0a, 32'hc3ef054b},
  {32'hc35f579f, 32'hc3971726, 32'h45096904},
  {32'hc4460cda, 32'hc21e79af, 32'hc40a4fd7},
  {32'h437e3298, 32'h445fc2f8, 32'h44169ddb},
  {32'hc2ca2fb0, 32'hc4ba12d6, 32'hc464bc77},
  {32'h43808fba, 32'h44c162c2, 32'h43b67cd1},
  {32'hc3e3e0ea, 32'hc31742a8, 32'hc50688b9},
  {32'hc3d4de4f, 32'h4499258e, 32'h45266558},
  {32'h43c5f662, 32'hc40d3f7f, 32'hc21e013a},
  {32'h43b75808, 32'hc3ea7f75, 32'h445f6f87},
  {32'h43217de2, 32'h42b49cd4, 32'hc4efcbb8},
  {32'hc3540aa4, 32'h44525c34, 32'hc31b9fa4},
  {32'hc3b24c58, 32'hc280fd68, 32'hc41dc683},
  {32'h4388619b, 32'h44a7a1c0, 32'h43e756ad},
  {32'hc359feac, 32'hc28b0644, 32'hc4ea28f3},
  {32'hc26c9f20, 32'h43d1cd8a, 32'h452152ff},
  {32'h429284c0, 32'hc3aa7cbb, 32'hc55c0a49},
  {32'h41944800, 32'h44d8b80c, 32'h431cd29c},
  {32'hc412dd87, 32'hc52e28dc, 32'hc1649c1f},
  {32'hc19b35c0, 32'h44a7df84, 32'hc1bf5fe1},
  {32'hc4ec2acc, 32'h439f9233, 32'hc398f91d},
  {32'h454d22b4, 32'h43be1af9, 32'h42fb9088},
  {32'hc3e52aa5, 32'hc55ad5cf, 32'h42fc421e},
  {32'h4527adf6, 32'h43a11f20, 32'h428e0652},
  {32'hc508f9e2, 32'hc394b691, 32'hc39b568f},
  {32'h45350603, 32'hc1c072f5, 32'h436fa297},
  {32'hc360d5d9, 32'hc50eff2f, 32'hc2d994c1},
  {32'hc32e6073, 32'h43bc88bc, 32'h44558d83},
  {32'h43a8e904, 32'h43494b97, 32'hc3bd2de9},
  {32'hc45604cb, 32'h43dea7bf, 32'h449dbe61},
  {32'h420a6860, 32'hc2e33aaa, 32'hc4799bc4},
  {32'hc438a411, 32'h44263ba2, 32'h449b4edf},
  {32'h42b26a84, 32'h431a7caa, 32'hc496042c},
  {32'hc5297ab0, 32'hc3e1a82f, 32'h43e77212},
  {32'hc2b900e1, 32'hc3ec01c4, 32'hc517ab3f},
  {32'h43e28e8a, 32'h442fa47f, 32'h4479269c},
  {32'h44986370, 32'hc39c08f5, 32'hc40220f8},
  {32'hc33504bc, 32'hc3684dc4, 32'hc206586e},
  {32'h45305171, 32'hc397e62c, 32'hc2190bb7},
  {32'hc4a04a08, 32'h43d20a0e, 32'h4418b26e},
  {32'h452688f1, 32'h441ee3d7, 32'h42d538fc},
  {32'hc4fb8bb7, 32'h4405bc44, 32'h4401b730},
  {32'hc2c95788, 32'hc491a091, 32'hc574bbf1},
  {32'hc44b82de, 32'h44969539, 32'h42fd08f7},
  {32'h43fba25a, 32'hc515cd38, 32'h437e4d1e},
  {32'hc5586b22, 32'h441e5eea, 32'h435a17cd},
  {32'hc5051207, 32'hc2921b78, 32'hc2769be4},
  {32'hc4cf5652, 32'h448ae88d, 32'hc41771e3},
  {32'h417c68b6, 32'hc537ea07, 32'hc030e5ed},
  {32'hc21c4e20, 32'h44d0acd5, 32'hc21e3298},
  {32'h44ecb95e, 32'hc2a0c7fe, 32'h420c9aea},
  {32'hc501da85, 32'hc3ea5230, 32'h415b3016},
  {32'h451c89b1, 32'hc41df913, 32'hc4175603},
  {32'h452d9792, 32'h4387377c, 32'hc3bf2705},
  {32'hc53ab1bb, 32'h4437be22, 32'hc441dc24},
  {32'h4429ecb8, 32'h41a2cc18, 32'h437dac7a},
  {32'h44d48ed2, 32'hc3ce72b2, 32'h436ba8ac},
  {32'h44b550a6, 32'hc2b75a66, 32'h44149195},
  {32'hc2e70ff2, 32'h455734f1, 32'h431360d5},
  {32'h43b7bd9a, 32'h41f40092, 32'h436f94cb},
  {32'hc50ce99d, 32'h44a1e850, 32'h4374fd59},
  {32'h445f77cf, 32'hc5099b2a, 32'h42d3290d},
  {32'hc5097c0c, 32'hc3a645e4, 32'h4342d1c8},
  {32'h439ef922, 32'h434bc5a9, 32'h45480705},
  {32'h4321d50d, 32'hc4ce5eef, 32'h44ae681a},
  {32'h42091d14, 32'hc4eb2ce2, 32'h4299899e},
  {32'hc18ef0d0, 32'h449fb9ad, 32'hc293eabc},
  {32'h44f2c6b8, 32'hc3e40b9a, 32'hc38cb13e},
  {32'hc47a8bac, 32'h43a69fee, 32'h42703965},
  {32'h43995a7f, 32'hc349ce43, 32'hc4d786a8},
  {32'hc5102c79, 32'h42866df4, 32'h43eb9d55},
  {32'h4402c48c, 32'hc4408d71, 32'h43394eba},
  {32'hc4d27a0e, 32'h43a76d82, 32'h44632ad0},
  {32'h441f9726, 32'h443af93b, 32'hc4b1976c},
  {32'h42c8b1f0, 32'h44dd2ebc, 32'h43500112},
  {32'hc3a9c33f, 32'hc51512b8, 32'hc3be50f6},
  {32'hc357142b, 32'h41a2c5a1, 32'h4544caa7},
  {32'h44a36671, 32'hc3c73873, 32'hc3a8dd68},
  {32'hc428d64c, 32'h43412896, 32'h45097916},
  {32'h42b9dd56, 32'hc522884b, 32'hc3497fba},
  {32'h444b6518, 32'hc20b583c, 32'hc4a6d5f4},
  {32'hc5615d61, 32'h41890df4, 32'h42d26d28},
  {32'h44e7019d, 32'h4378d5ee, 32'hc0fa0d3a},
  {32'hc4475a18, 32'hc4173be4, 32'h43c0a30f},
  {32'h450a104a, 32'hc3a95904, 32'h43f52924},
  {32'hc4907f13, 32'hc38dd566, 32'h441e8764},
  {32'h4535b946, 32'h4404d735, 32'hc31a0837},
  {32'hc44f3f4c, 32'hc544a9e6, 32'h431b8a22},
  {32'h450bf47e, 32'hc4122860, 32'hc36da857},
  {32'hc45014c2, 32'h43c731b2, 32'h44c13dfa},
  {32'h42adcac0, 32'hc415d61f, 32'hc4ccc71e},
  {32'hc475be92, 32'hc31a2bbd, 32'h43ed4c82},
  {32'h4357a31c, 32'h4496fda7, 32'h43857bb5},
  {32'hc4f75daa, 32'hc3d89299, 32'hc4156510},
  {32'h44dcd359, 32'h42882108, 32'h3ff97f4d},
  {32'hc44f4456, 32'hc39f043f, 32'hc4d6f4d6},
  {32'h4524a502, 32'h411c8058, 32'hc2212834},
  {32'h42bfeac8, 32'hc489ab27, 32'hc40300dc},
  {32'h43c1f0c6, 32'h44841102, 32'h44bd5d5d},
  {32'hc56d5e49, 32'h42272697, 32'h43216221},
  {32'h44ab74eb, 32'hc2e2810b, 32'hc41ecdd7},
  {32'hc4413172, 32'hc51742ee, 32'hc32083bb},
  {32'h446c8f96, 32'h44d4f8c7, 32'h4409da92},
  {32'hc3a7cdfa, 32'hc41b38e4, 32'hc36e7391},
  {32'hc31d3a59, 32'h4559853d, 32'h43565335},
  {32'h430e8a12, 32'hc4626adc, 32'hc4fe0ca3},
  {32'hc274b4e8, 32'h43eaac23, 32'hc3d25f76},
  {32'h43f3e2cb, 32'h4255b680, 32'hc363e35f},
  {32'hc460c849, 32'hc4a5443f, 32'h44078b9a},
  {32'h44f7635e, 32'h447bb9b5, 32'hc2e77fd0},
  {32'hc54a255c, 32'h440e21b8, 32'h40e45795},
  {32'h4542e93f, 32'h437441b6, 32'hc27d4acd},
  {32'hc4581338, 32'hc46965f4, 32'hc32367fa},
  {32'h44ba5445, 32'h437761ba, 32'hc33a2122},
  {32'hc4c9ab7a, 32'h4364292c, 32'hc37edd2f},
  {32'h452eea80, 32'hc3878c28, 32'hc38394c0},
  {32'hc4fea986, 32'h438e6dce, 32'h447339d0},
  {32'h434095be, 32'h4337fb75, 32'hc4624458},
  {32'hc2861941, 32'hc51f3cd3, 32'hc359e8b1},
  {32'hc4b975ce, 32'h43a7d738, 32'h4282650b},
  {32'hc3fa641c, 32'h4348d712, 32'h44a6c1d2},
  {32'h44bc1290, 32'h43af2688, 32'hc417d3d2},
  {32'h435e093d, 32'hc3884aa9, 32'h4358ac2d},
  {32'h452d6f97, 32'hc28928d2, 32'hc1a1b0af},
  {32'hc3ec6171, 32'h4458e21e, 32'h4523ad16},
  {32'h44bd7f68, 32'h437d2741, 32'hc3f9ada5},
  {32'hc43d5380, 32'hc49bbde6, 32'h43ec2fcb},
  {32'h4389a4c8, 32'h44915780, 32'hc4bd9b86},
  {32'hc36e2110, 32'hc4671037, 32'h4423e107},
  {32'hc36915f0, 32'h44805f8c, 32'hc4b5f940},
  {32'hc436fefd, 32'hc5255fee, 32'h43b204ef},
  {32'h436987ea, 32'hc382043e, 32'hc51deb9e},
  {32'hc552d775, 32'h43b165f6, 32'h4365cf4c},
  {32'h447fad10, 32'hc3c0afdd, 32'hc4f4a107},
  {32'h44d1921f, 32'hc4a14200, 32'hc4384523},
  {32'hc33fdd4c, 32'h45359a7c, 32'h41a6acca},
  {32'h43cdea10, 32'hc42869ee, 32'hc380e201},
  {32'hc51ebed1, 32'h444f0a86, 32'hc443e809},
  {32'hc33eaa03, 32'hc543fda0, 32'h43452a7b},
  {32'hc41eb1ef, 32'h43f077bc, 32'hc2a9e345},
  {32'h4430d84d, 32'h442362ed, 32'h43810889},
  {32'hc48ca4b7, 32'h4431fbda, 32'h440ea244},
  {32'h4434855b, 32'hc2fef6fe, 32'h424393ad},
  {32'h42a0ba66, 32'h44ecc74f, 32'h43b2b3d8},
  {32'h44b219a4, 32'h43699093, 32'h43430e05},
  {32'h44d8cd55, 32'h41ed4b5f, 32'h3f8a4800},
  {32'h4517191f, 32'hc26c9fbb, 32'h44003098},
  {32'hc50ad20a, 32'h44010f5f, 32'hc105187b},
  {32'hc31f7a22, 32'hc4f4c79c, 32'hc218bf5c},
  {32'hc43cb58e, 32'hc366ca0f, 32'hc4ee208e},
  {32'h44b411df, 32'h440e8634, 32'h448023a9},
  {32'h4508257f, 32'h42f16d36, 32'h4409e1fd},
  {32'h43e2b580, 32'hc50caaac, 32'h3f4ec096},
  {32'hc3cbeebe, 32'h446b9a5b, 32'hc42eb40d},
  {32'h440e85a8, 32'hc413a27a, 32'h4305220a},
  {32'hc434b7ef, 32'h44eaf20a, 32'h42722ba7},
  {32'h43864e39, 32'hc336b2d1, 32'h45295946},
  {32'h4420d907, 32'h434e1ee8, 32'hc360fca6},
  {32'h44d2a337, 32'hc23570a2, 32'h443372d9},
  {32'hc485634c, 32'h43a66d88, 32'hc47f7089},
  {32'hc403ac36, 32'h434562f0, 32'h44001f61},
  {32'h44309c7c, 32'h44a36720, 32'hc510d521},
  {32'hc1234740, 32'hc4517721, 32'h4491d85e},
  {32'h449123fd, 32'hc4287e52, 32'hc3b73ad8},
  {32'h44b7f8b7, 32'hc203e8b7, 32'h435f4e91},
  {32'h42c8fb8b, 32'hc4cb62fc, 32'h4397e30f},
  {32'hc4b71aa9, 32'hc1cde39f, 32'hc3c2fcd8},
  {32'hc379f107, 32'hc49d4f35, 32'h43448e4b},
  {32'hc480cfea, 32'h4397fb09, 32'hc4706303},
  {32'h4481597b, 32'hc487cd1d, 32'hc2d96597},
  {32'h429f2d74, 32'hc49b8d62, 32'h4508aca9},
  {32'hc36d8aee, 32'hc4be2a7e, 32'hc50378a2},
  {32'hc46688ee, 32'hc4b7a500, 32'h444f8c90},
  {32'hc4b70083, 32'hc3811be4, 32'h439eaaa4},
  {32'hc50e041b, 32'hc32769d7, 32'hc3c202c1},
  {32'hc2f87ff0, 32'hc3e39b22, 32'h43b39686},
  {32'h44bfd7f9, 32'h43c3f774, 32'hc37632d7},
  {32'hc36e582e, 32'hc38eb789, 32'h449d4585},
  {32'h435809b6, 32'hc1a50d6f, 32'hc54b0a54},
  {32'h42c0acc0, 32'h43c28f1f, 32'h433bba6e},
  {32'hc5859a3e, 32'hc239ad61, 32'hc3c9c5b3},
  {32'h4550f288, 32'h43c6740a, 32'h43a9438b},
  {32'h430b04f6, 32'h44c89ec7, 32'hc3a1d999},
  {32'h43eaec45, 32'hc563308e, 32'h433ce79c},
  {32'hc39a4503, 32'h44923891, 32'hc3171545},
  {32'h41a05040, 32'hc431a7b5, 32'hc2802a28},
  {32'hc3bdc345, 32'h452891a6, 32'h43c58a43},
  {32'h45323894, 32'hc466414d, 32'hc3598fd5},
  {32'hc4043554, 32'h42061e5e, 32'h43e78c39},
  {32'h4462ded6, 32'hc4348d67, 32'hc3ea459c},
  {32'hc49031ce, 32'h446a8afe, 32'h448b6d0d},
  {32'hc398395c, 32'h431184ed, 32'h4518bb77},
  {32'h44973bd6, 32'h43ba9871, 32'hc3a9d04d},
  {32'hc4f2bf68, 32'hc3a40e55, 32'h4286d871},
  {32'h4339514a, 32'h439473a2, 32'hc4b5403f},
  {32'hc30b4518, 32'hc4cb40db, 32'h4401c1e9},
  {32'h452b99f3, 32'h4210af67, 32'h440b07a5},
  {32'h444d23e0, 32'hc3f98596, 32'hc2cfa851},
  {32'hc547a02d, 32'hc3276e83, 32'h4455ca00},
  {32'h4474734b, 32'hc311627f, 32'hc4b999e2},
  {32'h43710918, 32'h437e6253, 32'hc5002c7b},
  {32'h42cc4808, 32'hc3b97896, 32'h43107f3c},
  {32'hc4881b06, 32'h4426b1c7, 32'hc3993488},
  {32'hc45f5ff2, 32'hc48e4860, 32'h436605e8},
  {32'hc3aab344, 32'h445389f9, 32'hc415e9b1},
  {32'hc5059dec, 32'hc2165a54, 32'hc2db25bf},
  {32'h4394624c, 32'hc4173dcc, 32'hc42230dd},
  {32'hc48e0c3e, 32'h43c1a8a9, 32'h444a99a4},
  {32'hc4c3ed61, 32'hc363f0d7, 32'hc253f3d9},
  {32'hc2b38e58, 32'hc45158d7, 32'hc384528e},
  {32'h43961946, 32'h45392f95, 32'hc3124d90},
  {32'h44d76505, 32'hc26f1d39, 32'hc22fbc45},
  {32'h44d801cf, 32'h44981443, 32'h43c0f307},
  {32'hc41c7d4e, 32'hc509643f, 32'hc3c527b3},
  {32'h454d1d5d, 32'hc3dae12a, 32'hc2bfeda2},
  {32'h4386fe9b, 32'hc4b48411, 32'h44121a4f},
  {32'hc438d690, 32'h44de958a, 32'hc4ea0a14},
  {32'h4506616a, 32'h4428c386, 32'h440a3bd6},
  {32'hc27395ee, 32'h442fc45e, 32'hc41dd793},
  {32'h440e5079, 32'h4447628b, 32'h4472584c},
  {32'h434b2e8b, 32'hc4efb031, 32'hc29e3063},
  {32'h43eff51c, 32'h436858ee, 32'h4432159d},
  {32'hc564f424, 32'hc21a9a62, 32'h40d3da56},
  {32'h4489ca64, 32'h42502906, 32'h449ae944},
  {32'h439c5dde, 32'h449acfab, 32'hc370bc23},
  {32'hc2edfa07, 32'hc43bb353, 32'h44b9cced},
  {32'hc3c74d16, 32'h44b15b1b, 32'hc4ae2a89},
  {32'h44f826f2, 32'h43261c3f, 32'h439fdffa},
  {32'h42b6b204, 32'hc49d1567, 32'hc452d7c1},
  {32'h440e8088, 32'h450f7f34, 32'hc3238ae7},
  {32'hc3df07d2, 32'hc414bb31, 32'hc42fa801},
  {32'h4557078e, 32'h438a0549, 32'h432ccb9f},
  {32'hc4a4440f, 32'hc3a0dcae, 32'hc4005740},
  {32'h44c4058f, 32'h43d54a81, 32'hc2854e9e},
  {32'hc5477157, 32'hc415edb0, 32'h43562623},
  {32'h455cafc6, 32'h4336e871, 32'hc448535b},
  {32'hc32ad0b4, 32'hc3a1c2f0, 32'hc39e1db8},
  {32'h4528cff9, 32'h4361629d, 32'h420d383d},
  {32'hc2ecaa08, 32'hc530cbec, 32'hc3932e40},
  {32'hc4c7dab2, 32'hc23a1bc6, 32'hc3b4dc23},
  {32'hc47e5c60, 32'h448aef39, 32'hc465387b},
  {32'h44b5aaa6, 32'h4321849a, 32'h433ccefb},
  {32'h4492a72d, 32'hc3ce2a43, 32'hc43dd758},
  {32'h44155aa6, 32'hc40a2c7c, 32'h44f6b641},
  {32'hc4934ed7, 32'h43c47f8f, 32'h425d8fad},
  {32'hc514c45a, 32'h441327a5, 32'h43c65774},
  {32'h42b695e4, 32'hc4c86dea, 32'hc44b60fe},
  {32'h43b146de, 32'h44dd9235, 32'hc3587bb3},
  {32'h44bc9509, 32'hc4277322, 32'hc49eaa6e},
  {32'hc4061519, 32'h444574f7, 32'h450ea9f7},
  {32'hc39f3810, 32'hc4826dd1, 32'hc3af4f73},
  {32'hc41d179e, 32'hc2c59f48, 32'h439b6ff8},
  {32'h43e21f07, 32'hc3eb3f0c, 32'hc4848d12},
  {32'h43c6e85b, 32'h4256fd02, 32'h43c6b312},
  {32'h44f1d539, 32'hc0048850, 32'hc433b901},
  {32'hc5633c50, 32'hc3f122f4, 32'h4325717d},
  {32'h42a04ed3, 32'h43aded87, 32'hc4e2344d},
  {32'hc50ec4b3, 32'h438f1e52, 32'h43c1957e},
  {32'h446e4016, 32'h42aaf7c8, 32'hc485474a},
  {32'h443e6650, 32'hc22501de, 32'h4439304e},
  {32'h444bd11c, 32'hc5149eef, 32'hc2c6f328},
  {32'hc5600723, 32'h43be42d5, 32'h43303384},
  {32'hc454fc87, 32'h42a01bf0, 32'h4214167b},
  {32'hc4212f6e, 32'hc3688f74, 32'hc403f899},
  {32'h43ee233c, 32'hc4b7bae2, 32'h439df91f},
  {32'h44383515, 32'h4446c069, 32'h433c3633},
  {32'hc3964d61, 32'hc0b4ba82, 32'hc36d87cd},
  {32'hc587a011, 32'h442e2686, 32'h43a0b5b1},
  {32'h457d36e6, 32'h43aea6bd, 32'hc411237e},
  {32'hc41f0628, 32'h43b28d92, 32'h42c5b3c2},
  {32'hc4b9bf60, 32'hc3937a00, 32'hc3e36dc0},
  {32'h453a4c74, 32'h436be2da, 32'h43a8eddd},
  {32'h450003d0, 32'h43374664, 32'hc29d8779},
  {32'h44ed6127, 32'hc3e57326, 32'h4343c118},
  {32'hc52dddfc, 32'h432a8f97, 32'h441656fc},
  {32'h4456939a, 32'h42f92800, 32'h42b9fc81},
  {32'hc412c2ac, 32'h44d1686e, 32'hc3b4a521},
  {32'h44bc1a6e, 32'hc4d148bd, 32'hc3849179},
  {32'hc4d9ff3d, 32'hc364b59a, 32'h438693b4},
  {32'h43f97a78, 32'hc341fd40, 32'h43fdc460},
  {32'hc37b04b8, 32'hc44cfe30, 32'h442c3dc3},
  {32'h448d6e53, 32'hc30bf389, 32'h43a610bb},
  {32'hc2a75900, 32'h44699e5f, 32'h449600e7},
  {32'h43c8555a, 32'hc48bcf0b, 32'hc2631076},
  {32'hc4b09711, 32'h4283c139, 32'h43829287},
  {32'h43316b82, 32'hc3a47f61, 32'h4400d527},
  {32'h42da9f38, 32'h444323ef, 32'h44abcf89},
  {32'h449b8c8d, 32'hc4595f47, 32'h422f2084},
  {32'hc41c651f, 32'hc46c35d0, 32'h439e8718},
  {32'h4535e450, 32'hc38eb5f0, 32'hc48cf4b3},
  {32'hc39468ae, 32'h4325bd95, 32'h4373683a},
  {32'hc3e84daa, 32'hc54b2f7d, 32'hc4257cea},
  {32'h42d17795, 32'h4551962a, 32'h41154379},
  {32'h43c5f9e4, 32'hc3f3e5a1, 32'hc383cdaf},
  {32'hc493ae0f, 32'h444a224c, 32'h43e057d0},
  {32'h448bcf0d, 32'hc4a3a39e, 32'hc47edb8d},
  {32'h41ebbbc0, 32'hc3f64837, 32'hc173fc7e},
  {32'hc501fef4, 32'hc358158e, 32'h439489e4},
  {32'h44396c5d, 32'h43c85620, 32'hc3c18018},
  {32'hc50fb126, 32'hc4b5085e, 32'hc3acf9ba},
  {32'h44b1a3d6, 32'hc3456f35, 32'hc294c5f7},
  {32'h446dd4e4, 32'hc4823c7c, 32'h426af397},
  {32'h4504a2d3, 32'h445e70f9, 32'hc3d5d9e8},
  {32'hc3af4a58, 32'hc4e31607, 32'hc1dd3bc0},
  {32'hc34db1c0, 32'h446866d1, 32'hc2fe9187},
  {32'hc4e2c594, 32'hc3ffee89, 32'h43e28f8f},
  {32'h44f038dd, 32'h44061812, 32'hc2dc0910},
  {32'hc4c8ac12, 32'h4338f190, 32'hc3e5ab51},
  {32'h4478dde4, 32'h42278943, 32'h4401b621},
  {32'hc51087bd, 32'hc3bfd51c, 32'h43343d17},
  {32'h44b27e79, 32'h4350d985, 32'hc2a8709c},
  {32'h438a947a, 32'hc433221d, 32'h433ed21f},
  {32'hc31b711e, 32'h4532f577, 32'hc386743d},
  {32'hc31115c9, 32'hc3eec0ff, 32'hc4ca4967},
  {32'h42dfa2f0, 32'h437622db, 32'h44736ac6},
  {32'hc530b708, 32'h437a6ebc, 32'hc25ca71a},
  {32'h44525f90, 32'h42ba38be, 32'hc3d5cc9a},
  {32'hc3cfaa49, 32'hc2aac6f3, 32'hc518d7f5},
  {32'h446a91e0, 32'h449ce716, 32'h445e7c70},
  {32'h40f886aa, 32'hc429c24f, 32'hc3c73d47},
  {32'h4432e28d, 32'h43fb8564, 32'h42aad61c},
  {32'hc4d67f13, 32'hc394d476, 32'hc3c2707d},
  {32'hc47e815e, 32'h42d18018, 32'hc2174103},
  {32'hc279eaa0, 32'hc39a9370, 32'hc2a793c2},
  {32'hc42ec0a0, 32'hc504e09d, 32'hc30af66e},
  {32'h44b764ed, 32'h43d708ce, 32'h441780b6},
  {32'hc40b1740, 32'hc48df813, 32'h4410c69b},
  {32'h44dfa487, 32'h4414d590, 32'hc315e3c4},
  {32'hc32dd390, 32'hc4ade190, 32'hc1f51dd3},
  {32'h45190b58, 32'h43e18abd, 32'hc3a4057e},
  {32'hc55c9d2a, 32'h42ccb1b3, 32'hc3e26e06},
  {32'h43fc305d, 32'h444da2a6, 32'h4451871c},
  {32'hc4576c73, 32'hc286b90d, 32'h43f8032f},
  {32'h433f935a, 32'h4555f725, 32'h43baaae2},
  {32'hc5225769, 32'hc22e7f50, 32'hc31c2f6e},
  {32'h449eb16b, 32'h43ca8248, 32'hc26afb60},
  {32'hc2a497a0, 32'h41594caa, 32'h4513aed7},
  {32'h433f9407, 32'h43d3d42d, 32'h43e32d32},
  {32'hc38d5edc, 32'hc3be3d4f, 32'hc3eed591},
  {32'hc2be09ae, 32'hc3933014, 32'hc54f8e1a},
  {32'hc3f10479, 32'h4425aa2a, 32'h44ae99d9},
  {32'h43ea3912, 32'h43ce2f21, 32'hc401ed72},
  {32'hc448d79a, 32'hc47cf3cb, 32'h4446296c},
  {32'h452f1d19, 32'h444cc550, 32'hc3c4adf0},
  {32'hc381cbb9, 32'hc50c633b, 32'hc46a352e},
  {32'hc3ef0607, 32'h44f89542, 32'hc403fafc},
  {32'hc4a70b89, 32'hc3fa0097, 32'h42996893},
  {32'h451b1730, 32'h43ef40db, 32'h4288f1f5},
  {32'hc51c461b, 32'h43d7e53e, 32'hc3c4113c},
  {32'h44dbf336, 32'hc3e276b9, 32'hc497f2a3},
  {32'h443e7d9d, 32'h43c63a95, 32'hc4ce14d2},
  {32'hc3e7f1e9, 32'h450827ee, 32'hc1f06a02},
  {32'h42a53968, 32'hc504339d, 32'h439dd449},
  {32'h43b2de10, 32'h455bf2f8, 32'h4309c9ca},
  {32'h453fa25b, 32'h42ca37bb, 32'hc41ab43e},
  {32'h43e0df3c, 32'h446b85bb, 32'hc320c214},
  {32'h45130c28, 32'hc41c99be, 32'hc3642f7e},
  {32'hc56240d6, 32'h3f5d0618, 32'hc28bce51},
  {32'hc4c7171d, 32'hc2505a0f, 32'hc30cb5dc},
  {32'hc483b936, 32'h4279d3e0, 32'hc4569ede},
  {32'hc316809a, 32'hc4c343c6, 32'h43eca503},
  {32'h44464b59, 32'h439054e9, 32'hc49676c8},
  {32'hc3ad6670, 32'hc42cf558, 32'h44949371},
  {32'hc4924048, 32'h44287ffd, 32'hc3e05410},
  {32'h439167da, 32'hc492abf2, 32'h43a342b6},
  {32'hc37fe629, 32'h44b78342, 32'h44a31ac6},
  {32'h446cc24a, 32'h42e02c2f, 32'h44dd544b},
  {32'h4277f3f5, 32'h42db4b9a, 32'hc4b6cde3},
  {32'h441b0c52, 32'hc4e368a5, 32'h43c7db36},
  {32'hc45c0ff8, 32'h4403d25c, 32'h432b0698},
  {32'h44c50658, 32'hc2fda505, 32'h441353c5},
  {32'hc47cd133, 32'h44e20e22, 32'hc1356156},
  {32'h4424d735, 32'hc381d7a5, 32'h44a6beb6},
  {32'hc30edb8c, 32'h4463092c, 32'hc2a39069},
  {32'h455d134d, 32'h4395bdb1, 32'h430519f8},
  {32'hc36f1a58, 32'h43025256, 32'hc50c5f7a},
  {32'h4539f57a, 32'hc3ed7d64, 32'hc32e048c},
  {32'h444f9efa, 32'h4492434a, 32'hc5154dca},
  {32'h42147688, 32'h43ee66a5, 32'h45054425},
  {32'h43b173f7, 32'h4448dda5, 32'hc452ed67},
  {32'hc31eacd8, 32'h445f85e0, 32'hc36fcc3a},
  {32'h44b1290e, 32'hc47e0b84, 32'h4452e911},
  {32'hc3763688, 32'hc39e8fa9, 32'hc47bbed0},
  {32'hc343b650, 32'hc4148f13, 32'hc3992f1f},
  {32'hc43c9358, 32'h43824e20, 32'hc4bc3fc8},
  {32'h4526aceb, 32'hc3b819d8, 32'h4463fead},
  {32'hc4024b9d, 32'h4486a0e0, 32'h45299f6a},
  {32'h441460a1, 32'h4349f128, 32'hc4f15a21},
  {32'h447d0720, 32'h44375a7c, 32'hc2d4d8ab},
  {32'h4532fcd8, 32'h43b0d418, 32'hc3e63849},
  {32'hc40c6e9f, 32'h40b5a832, 32'hc4cbb9d5},
  {32'h41886e4c, 32'hc4e33cc8, 32'hc3b66fa1},
  {32'h441bf202, 32'h43dade66, 32'hc3aa07d2},
  {32'h42bfd134, 32'h408c665f, 32'h4510efbf},
  {32'h43ad6286, 32'h4546cde0, 32'hc298d6c2},
  {32'hc4e46ab0, 32'h436ebc50, 32'h434a0e83},
  {32'hc4788011, 32'hc44c15d7, 32'hc4393234},
  {32'h454bd3ef, 32'hc370706a, 32'hc416cf44},
  {32'hc4562b66, 32'hc1bf0c34, 32'hc3feb888},
  {32'h4515360c, 32'hc410984c, 32'h443123bd},
  {32'h43485550, 32'h445d3377, 32'hc2ace961},
  {32'h45372d86, 32'h44136007, 32'h43040e5c},
  {32'hc4ce2904, 32'h4496a262, 32'hc3fd518a},
  {32'h43c924f0, 32'hc4936296, 32'h410e2073},
  {32'hc4fb0f4e, 32'hc3aa527a, 32'hc36a0854},
  {32'h43a2e88a, 32'h441434ac, 32'hc4ae6667},
  {32'hc46e215c, 32'hc4443668, 32'h438e62ab},
  {32'hc515a15a, 32'h418ccdd7, 32'h435506f6},
  {32'h44c057e4, 32'hc28d2af2, 32'hc2186d49},
  {32'hc531e368, 32'h4239a2ab, 32'hc245ff58},
  {32'hc36eaee0, 32'h45334ca7, 32'hc24e7124},
  {32'hc380f564, 32'hc4ec42c1, 32'h43ed89b7},
  {32'hc2a795d8, 32'h43188c17, 32'hc4bb487b},
  {32'h44c90b16, 32'h4308e572, 32'h43bd0202},
  {32'hc4ab3650, 32'hc4c88454, 32'h44d6b9ab},
  {32'hc2b25e82, 32'hc40057cb, 32'hc4cbef15},
  {32'h450b882a, 32'h441e90da, 32'hc423148e},
  {32'hc4ca5f50, 32'hc4bb6cc0, 32'h436df3bd},
  {32'hc2bfb2d2, 32'h439d8b33, 32'h442163e4},
  {32'hc45f5d07, 32'hc3606532, 32'h450ebd99},
  {32'h4481b0c3, 32'h44397aa9, 32'hc2a68de6},
  {32'h446a7653, 32'h43325150, 32'h445991f4},
  {32'h45083a6f, 32'hc40de397, 32'hc2804d22},
  {32'hc55e86fe, 32'hc340bb73, 32'h43702d3f},
  {32'h4311ea42, 32'h42f24205, 32'hc2996ec7},
  {32'hc427aecc, 32'hc499403a, 32'hc34e8ee6},
  {32'h443d6dd6, 32'h447efe98, 32'hc327af1d},
  {32'hc496c7e3, 32'hc404b6b6, 32'h42e6d6fa},
  {32'h4375065c, 32'h4544be75, 32'hc40f258a},
  {32'hc3ad46cc, 32'hc4bee7af, 32'h438db97d},
  {32'h44181e12, 32'h4382eb33, 32'hc37e1af9},
  {32'hc1c92340, 32'h44bbd5a4, 32'h43203268},
  {32'h431aaeba, 32'hc4534b00, 32'hc3acfcd2},
  {32'h44ebd506, 32'h445bc5c1, 32'h43f034e2},
  {32'h43dda527, 32'hc4a38870, 32'hc40bdd3a},
  {32'h4537efeb, 32'h44260c78, 32'hc1dc4dbf},
  {32'hc396d4b4, 32'h4391d5bc, 32'hc42cf204},
  {32'h45166e25, 32'hc341a2c4, 32'hc1d5089e},
  {32'hc46bc4bf, 32'hc4887d25, 32'hc48713b5},
  {32'h4487d1d8, 32'h443cc96f, 32'h44402539},
  {32'hc39e0fcd, 32'hc494d26c, 32'hc2981212},
  {32'hc4a285e5, 32'hc4d4e374, 32'h452b4ee5},
  {32'hc302a130, 32'h44202c97, 32'hc5266913},
  {32'h44569ef5, 32'h427aa4f9, 32'h4476e7b4},
  {32'hc44eaf8c, 32'hc48ef251, 32'hc3ad29b6},
  {32'h44b3371b, 32'h4479ab78, 32'hc3772115},
  {32'hc4bd966f, 32'hc3653377, 32'h438ad1ea},
  {32'h43f53768, 32'h43cbcdc1, 32'h43fefbe6},
  {32'h43f30866, 32'hc3c8d155, 32'hc52ca33b},
  {32'hc39caa2b, 32'hc2cc8096, 32'h4402581c},
  {32'hc5157515, 32'hc456b618, 32'hc2ebbbf6},
  {32'h4398bb04, 32'h454c358b, 32'h42e59a7f},
  {32'h44fd23af, 32'h432d8077, 32'h428d14e5},
  {32'hc266a810, 32'h455307b9, 32'h4387a40e},
  {32'hc449d4c6, 32'hc4a20a16, 32'h42d28001},
  {32'h44e20783, 32'h4362d7a1, 32'h4404e5ac},
  {32'hc512f590, 32'hc39bead8, 32'hc447d783},
  {32'h43d3c3e0, 32'hc30de2ae, 32'hc44d492b},
  {32'h43bb8386, 32'hc5057a97, 32'h438b482e},
  {32'h4328c867, 32'h448abd6a, 32'h4411e45b},
  {32'hc3cd50bd, 32'h42b71050, 32'hc4364800},
  {32'hc4ea96ef, 32'h44502ec2, 32'h43836538},
  {32'hc308bae4, 32'hc3cde345, 32'hc53ac623},
  {32'h441b802a, 32'h44722855, 32'hc389d5ee},
  {32'h45363446, 32'hc43f8a00, 32'hc3db032c},
  {32'hc517041b, 32'hc283bc2e, 32'h43d59f12},
  {32'h4326f360, 32'h4344a9f3, 32'h4357d5dd},
  {32'h4351b916, 32'h43ac53c1, 32'h44ae8c64},
  {32'h44091a6c, 32'hc2c05d91, 32'hc47c1a2a},
  {32'h43fecc26, 32'h44ba7e20, 32'h43cf2758},
  {32'h44465052, 32'h429ef072, 32'hc4b69df4},
  {32'hc37a612e, 32'h452042cf, 32'h42f0c081},
  {32'hc40e3e10, 32'hc401a3a7, 32'h420f217c},
  {32'hc3491d2a, 32'h4496f986, 32'h44aaf3b6},
  {32'hc4a18c8f, 32'h4277e18d, 32'hc451bc27},
  {32'h443b19c6, 32'h43fcb84b, 32'h4443f8bf},
  {32'h4481447c, 32'hc4745a41, 32'hc42be246},
  {32'hc44494d4, 32'h44d34ff5, 32'h4409c23c},
  {32'h443f0b20, 32'hc4412d53, 32'h4336f1d8},
  {32'hc4a203ca, 32'h44a4e33c, 32'hc2fe41e3},
  {32'h4414c592, 32'hc3bf2f47, 32'h439b1aef},
  {32'h44195453, 32'h44779392, 32'hc2e7f65e},
  {32'h457052f4, 32'h43f2e428, 32'h436d3671},
  {32'hc4bf9eaf, 32'hc3c13c77, 32'hc4041cf3},
  {32'h44cb1b10, 32'hc2b7255a, 32'hc3470a71},
  {32'h44adcee7, 32'hc3c220d6, 32'hc40fdd55},
  {32'hc45117a6, 32'hc29a5abc, 32'hc3a0697c},
  {32'h452aaab6, 32'h42af71d5, 32'h443ff3a0},
  {32'hc4573969, 32'h43b844f9, 32'hc438ce63},
  {32'h4524fb9f, 32'hc382c278, 32'hc31deb98},
  {32'hc424dcd3, 32'h4506763d, 32'hc2e33343},
  {32'h452be056, 32'h4406456e, 32'hc34b5253},
  {32'hc3fa05c4, 32'h44b480ae, 32'h42c632d7},
  {32'h44fa57f3, 32'hc48d6d48, 32'h436526f9},
  {32'hc3936010, 32'hc36318fb, 32'hc44d801a},
  {32'h44ccf437, 32'hc38f420f, 32'h439c3e30},
  {32'hc3c6ebc0, 32'h4391f970, 32'hc546888b},
  {32'hc28d590c, 32'h433fffba, 32'hc480e67e},
  {32'hc34b8ae6, 32'h451cd35e, 32'h41284435},
  {32'h440792e6, 32'hc38d3178, 32'hc5305fd9},
  {32'hc358f214, 32'h4336a94e, 32'h44d4f9d6},
  {32'h44efabc2, 32'hc3962188, 32'hc3c45a84},
  {32'h41994780, 32'h44a1dbf1, 32'h442f31b5},
  {32'h45253a56, 32'hc42acc3c, 32'h41aba9e0},
  {32'hc48efedd, 32'h44a8200a, 32'h449e9d0a},
  {32'h4537b63a, 32'h43900039, 32'hc451eb3c},
  {32'h42ebd0aa, 32'h446cb715, 32'h43a1c462},
  {32'h442acc14, 32'h428aa8f8, 32'hc39b14d4},
  {32'hc307cdb8, 32'h447782e3, 32'h448662ce},
  {32'hc327d908, 32'hc42ccf41, 32'hc414f903},
  {32'hc445a98d, 32'h451943b6, 32'h42fa446f},
  {32'h44b40091, 32'hc43c8548, 32'hc3ceda4d},
  {32'hc33689b9, 32'hc38dbc1a, 32'hc4d5c39e},
  {32'hc47b7290, 32'h42a83242, 32'h431de14a},
  {32'h450d2355, 32'hc2f98068, 32'h4418cc1a},
  {32'hc489b7df, 32'hc4d11e8d, 32'hc3b06942},
  {32'hc394319e, 32'h45116de2, 32'h43daf4eb},
  {32'hc4ef41e5, 32'h4380a578, 32'hc29f6e06},
  {32'h45197ee7, 32'h44288b1f, 32'h42050cbc},
  {32'hc5936fc4, 32'h4305d6f6, 32'h43d2c4cd},
  {32'h4445f9da, 32'h43ce7912, 32'h432c2f4c},
  {32'hc4a347ae, 32'hc3c9f375, 32'h4472ede6},
  {32'h4519a5b2, 32'h43ba9935, 32'h43613515},
  {32'h41a07a55, 32'hc3c58c40, 32'h44825e03},
  {32'h441dac56, 32'hc2a626ba, 32'h45189512},
  {32'h437af1de, 32'hc4cf0000, 32'h43997401},
  {32'hc4cc6514, 32'h4313ffb6, 32'hc30988aa},
  {32'hc4efcc0e, 32'hc4531492, 32'h4378d50a},
  {32'h449348cc, 32'h443aa918, 32'h4376a166},
  {32'hc38ef53e, 32'hc501b1e3, 32'hc3f24203},
  {32'h41839800, 32'hc4194e14, 32'h448068bc},
  {32'hc53bffcd, 32'hc2ef170b, 32'hc3ecfe29},
  {32'hc49b64a8, 32'hbfead588, 32'hc362dd66},
  {32'hc3362a9d, 32'hc5097c22, 32'hc3e9eeb8},
  {32'h44e50376, 32'h43310995, 32'h43c61567},
  {32'h423948a8, 32'hc2797841, 32'h4312a2e6},
  {32'hc385f06a, 32'h45257662, 32'h43eb926f},
  {32'hc40b991f, 32'hc4c30de2, 32'hc371b5c4},
  {32'h447ac202, 32'hc339f6ab, 32'h4438a61b},
  {32'hc3cc828d, 32'h443dd5f3, 32'hc3fbcf0a},
  {32'hc51289a7, 32'hc33dfee0, 32'hc29e38af},
  {32'h4424b1f7, 32'h4509fa43, 32'h4462a6ec},
  {32'hc406a39d, 32'h4257a5f4, 32'hc279cced},
  {32'h44c385c2, 32'hc24ddefb, 32'h43a07ace},
  {32'hc3bae5f3, 32'hc5718b34, 32'hc2eb5e72},
  {32'h44b5df1c, 32'h43a1e4d5, 32'hc3b61f68},
  {32'hc4d6a76c, 32'hc33fbb06, 32'h429d077c},
  {32'h43cae36a, 32'h44aa11a0, 32'h44926c64},
  {32'hc391b048, 32'h41875115, 32'h44705bc1},
  {32'h439c3195, 32'h449a3194, 32'hc5038ebb},
  {32'hc45f66f4, 32'h4400f505, 32'hc4960f9c},
  {32'hc4006fd9, 32'h44516faa, 32'hc3a5f4aa},
  {32'hc3fa3ae7, 32'hc4709f8c, 32'h441d4e87},
  {32'h452016a1, 32'h4283d1dc, 32'hc1beed0a},
  {32'hc51f5049, 32'hc3a31790, 32'hc2bdf09e},
  {32'h44fa0c19, 32'h4251561b, 32'hc41692d7},
  {32'hc5052002, 32'hc3923f21, 32'h431624af},
  {32'hc449d048, 32'hc2b061bb, 32'hc42b6c7a},
  {32'hc41c887e, 32'hc53f7419, 32'hc3c5423b},
  {32'h42725450, 32'h4458a062, 32'hc54870e8},
  {32'hc3833a19, 32'hc3c1b47f, 32'h4497ace3},
  {32'h442ac4e2, 32'h44e1bfe4, 32'hc437ff50},
  {32'hc3a77aeb, 32'hc36f4ca4, 32'h4503a6aa},
  {32'hc463f70c, 32'h43ced3dd, 32'hc281fee2},
  {32'hc57525a3, 32'h441021a0, 32'h43148ead},
  {32'h454f733a, 32'hc43be11f, 32'hc40a1e9b},
  {32'h43856e79, 32'hc54c1a0a, 32'hc2bef33a},
  {32'hc3f0e607, 32'h4401a868, 32'h42bd478c},
  {32'h444f79b5, 32'h44388a08, 32'hc4818f8f},
  {32'hc39cb858, 32'h42a4770b, 32'hc3d574d6},
  {32'h442002ae, 32'hc4e7b128, 32'hc3dcb9ce},
  {32'hc519f6fc, 32'hc38b2b4f, 32'hc2808997},
  {32'h428c8e80, 32'h40ee887c, 32'hc1e63006},
  {32'hc57a2839, 32'h432c847b, 32'h44139add},
  {32'h44825fdc, 32'hc3b26ee2, 32'h44118772},
  {32'h43391840, 32'hc41af1a3, 32'h448abe1a},
  {32'h4389d97c, 32'hc4675512, 32'h4468bf0b},
  {32'hc51ff77d, 32'h42a0b985, 32'hc3d8dfde},
  {32'hc3be6718, 32'hc528e842, 32'h434f4d1c},
  {32'hc2c032ec, 32'hc3cc5e28, 32'hc50a9d12},
  {32'hc41d463d, 32'h4402dbec, 32'h44af27af},
  {32'hc32936d8, 32'hc353ede1, 32'hc50a7168},
  {32'h43dac347, 32'hc3c54610, 32'h43a571a9},
  {32'h43518e62, 32'h44065a2e, 32'hc3720960},
  {32'h4257d9e0, 32'hc4c95f18, 32'h43ef51e3},
  {32'hc452aa9c, 32'h44e0f24c, 32'hc46e4ca8},
  {32'hc473a5b8, 32'hc2b91563, 32'h436afd30},
  {32'hc37013f8, 32'h449746e9, 32'hc4cf9473},
  {32'h442b52f6, 32'hc41b4e6e, 32'h4493ed56},
  {32'hc4c34d0a, 32'hc30f0e0f, 32'hc33261b1},
  {32'h44568cf8, 32'h41b9921f, 32'h44840ff0},
  {32'hc57b734a, 32'h43fdfb64, 32'hc3602c8a},
  {32'h445d1366, 32'hc315f005, 32'h44142884},
  {32'hc303d0fa, 32'h44f57970, 32'hc4db2411},
  {32'hc35b49f0, 32'h4511569b, 32'h44f91ed5},
  {32'h443239f8, 32'hc3cf9e28, 32'hc349a45c},
  {32'hc4684576, 32'hc3a111fd, 32'hc340874e},
  {32'h44fe648d, 32'hc3b6c821, 32'hc2867120},
  {32'hc5295dcf, 32'hc22b23aa, 32'hc3cf60f1},
  {32'hc4d1e412, 32'hc340078f, 32'h41bf2ddb},
  {32'hc35f044f, 32'h440faf6c, 32'h42777d3a},
  {32'h4522fbd6, 32'hc3a93863, 32'h441eba07},
  {32'h43e67d49, 32'hc38bc568, 32'h440ccc54},
  {32'h43f8176e, 32'hc37fad6a, 32'hc3ad38c2},
  {32'hc425db82, 32'hc49f5551, 32'h4429c3ac},
  {32'hc29d6f98, 32'hc3d08349, 32'hc3e48730},
  {32'hc48471a4, 32'h4411bc85, 32'hc48d3ee3},
  {32'h42e4c770, 32'hc1e7f3be, 32'h445da596},
  {32'hc36fa11c, 32'h43f72045, 32'h43b5af73},
  {32'h44e4a1b6, 32'h4340cac5, 32'h419ab117},
  {32'h439d3fd0, 32'h448825d7, 32'hc4bf7716},
  {32'hc4e6409e, 32'hc39816a6, 32'hc288027f},
  {32'hc511ad10, 32'hc3ff7a8d, 32'h439d8a41},
  {32'h45430e2b, 32'hc3c95b78, 32'hc4103ac0},
  {32'hc50d9bb1, 32'hc3570056, 32'hc3004dab},
  {32'h43c78dae, 32'hc57f4846, 32'hc29fb576},
  {32'h42ae747c, 32'h4551a1ec, 32'h428706d5},
  {32'hc4b3698a, 32'hc4194aef, 32'h4328beca},
  {32'hc54446a2, 32'h41104ed9, 32'hc401dbdf},
  {32'hc30583b8, 32'hc5339a75, 32'hc40a091d},
  {32'hc3f238e7, 32'hc48deeaf, 32'h43b762d6},
  {32'h4356693c, 32'hc32fbea8, 32'hc4985d42},
  {32'hc3c22532, 32'hc4f7f1da, 32'h4504dbc8},
  {32'hc4fc3f6f, 32'hc43c5433, 32'h4346d36a},
  {32'h42804f48, 32'h441690e7, 32'hc3f2e043},
  {32'hc1a15458, 32'hc35e5d41, 32'h443b1aae},
  {32'h447df818, 32'h44d7338b, 32'h438ef8d2},
  {32'hc4bce39b, 32'hc479fea2, 32'h44426dc9},
  {32'h425353f6, 32'hc27b7236, 32'hc4f3940c},
  {32'h446a5d1a, 32'h43f0611e, 32'h431dac50},
  {32'hc4b6e90e, 32'h440f8968, 32'h44a9964c},
  {32'h4513478f, 32'h438b2235, 32'hc451540f},
  {32'h4424a9ca, 32'h44909b77, 32'hc406dc89},
  {32'hc51e2393, 32'hc358c855, 32'h43b88b25},
  {32'h452d9664, 32'hc201a109, 32'hc3b67b8c},
  {32'hc4fd4a88, 32'hc43fad6b, 32'h4401ae4b},
  {32'h433a91ec, 32'hc24cf323, 32'hc486769a},
  {32'hbfe31010, 32'hc408d302, 32'h44a15c53},
  {32'hc32ea986, 32'h43d6ca9b, 32'hc4325c9d},
  {32'hc5a141ab, 32'hc34cfa80, 32'hc3a6ef74},
  {32'h451dfad8, 32'h440e3acf, 32'hc334c9c9},
  {32'hc3f2dddc, 32'hc45179b2, 32'h4344462a},
  {32'h4494554c, 32'h44c0a88e, 32'h4385afd1},
  {32'hc422981d, 32'hc4587d5a, 32'hc1a840dd},
  {32'h439348aa, 32'h45047f40, 32'hc3a6aaae},
  {32'hc58280d8, 32'hc39433e0, 32'hc396f1cd},
  {32'hc4b6a30e, 32'h440ae234, 32'h420d9978},
  {32'hc32af880, 32'h4425fb8a, 32'h41eff6d9},
  {32'hc4004a38, 32'hc3861d60, 32'hc455adb8},
  {32'h4440ec00, 32'h44a44506, 32'h4431edec},
  {32'hc5127537, 32'h431da21d, 32'h430e324e},
  {32'hc1482e86, 32'hc41f46c4, 32'h44e2397d},
  {32'hc34e6fb7, 32'hc368ab8a, 32'hc53063cd},
  {32'hc3594375, 32'h4420e754, 32'h44583651},
  {32'hc34935b0, 32'hc38dcd59, 32'hc4aff505},
  {32'h4488c216, 32'h42f923dd, 32'h4418792c},
  {32'h435dafe4, 32'hc2c4817c, 32'hc470a9d8},
  {32'h44df844a, 32'h4394ce0c, 32'h438f0da7},
  {32'hc40d56a6, 32'hc3a5f7fb, 32'hc412305b},
  {32'h43d01a9f, 32'h4456d35a, 32'h42a5e9dd},
  {32'hc284d50e, 32'hc2e3cb51, 32'hc4833a00},
  {32'h44633287, 32'h44d1ea2b, 32'h4323158f},
  {32'h43bf830e, 32'hc3b74c0e, 32'hc52513bc},
  {32'hc352ffc0, 32'h448bbeb4, 32'h44cec6cd},
  {32'hc4ad2130, 32'hc345b3f0, 32'hc47d6a77},
  {32'hc4e35dfd, 32'h43d63d3c, 32'h43b9f90f},
  {32'hc50243ce, 32'hc3efff08, 32'hc100e6a9},
  {32'h44ae9bc6, 32'h45036245, 32'h43a6f583},
  {32'hc402b019, 32'hc43c90b1, 32'h42bf6409},
  {32'h42f67810, 32'h453ae4cc, 32'h43ff35ae},
  {32'hc488ff61, 32'hc4270991, 32'h42d4232e},
  {32'h44b0088d, 32'hc3199db5, 32'hc2f16494},
  {32'hc517c107, 32'hc3a5e486, 32'hc36138ce},
  {32'h451f6038, 32'hc29f2fd4, 32'hc337b190},
  {32'h433dfff8, 32'hc43424db, 32'hc49c1b8c},
  {32'hc4d0bc3c, 32'hc3958712, 32'hc338c188},
  {32'h433dbe8b, 32'h442358d6, 32'hc476e750},
  {32'hc405e955, 32'h4478ecb9, 32'h449e1a2d},
  {32'h450b3e47, 32'hc30cce28, 32'hc22739ef},
  {32'hc4ced882, 32'h424beb17, 32'h439f1d7f},
  {32'h44981a39, 32'hc39c5aaa, 32'hc4b4f42b},
  {32'hc5577308, 32'hc1817ef8, 32'h440e42f4},
  {32'h4522d3a6, 32'h4374e7a8, 32'hc309ffa0},
  {32'hc50e992b, 32'hc34d15c2, 32'h4418f364},
  {32'hc39e4e40, 32'hc47ae8ac, 32'hc3a982fa},
  {32'h43143b8a, 32'hc4df6e04, 32'h444bc6c5},
  {32'h44fc4350, 32'h4349f09b, 32'hc3e67aab},
  {32'hc3fcc966, 32'h42dc592a, 32'h445176f3},
  {32'h445c32f4, 32'hc399432b, 32'hc3d5ef42},
  {32'hc08545e0, 32'h440e04eb, 32'h4562a973},
  {32'hc3a1d495, 32'hc45a2221, 32'hc440793e},
  {32'h432c5210, 32'h442fbbe3, 32'h44d1f3f2},
  {32'h43a31f10, 32'hc495f8a4, 32'h4379304a},
  {32'hc3f09756, 32'h44c95ff2, 32'h42a215b1},
  {32'hc45ae109, 32'h430ddd7f, 32'h429b9ada},
  {32'hc4f59b3c, 32'h44c80012, 32'hc2ed16a0},
  {32'h44acf189, 32'hc4d67c4b, 32'h438a5efb},
  {32'h43ca061e, 32'h44330cdf, 32'hc3b16a7a},
  {32'h456a76ea, 32'h43ff0496, 32'h43a6ec9e},
  {32'hc502992c, 32'h433eca65, 32'hc2ed20cb},
  {32'h44eb7d13, 32'h4345b193, 32'hc3a108d2},
  {32'hc38e109e, 32'hc3bf67f8, 32'h4413b7e9},
  {32'hc41d4838, 32'hc35ad717, 32'hc4f99228},
  {32'h452ba174, 32'hc281d1f6, 32'h43effbd2},
  {32'hc0e7bbd0, 32'h450eeee4, 32'h436ed004},
  {32'h449add70, 32'hc40052b0, 32'h438cd5ef},
  {32'hc4fe224a, 32'h44117799, 32'h439a836d},
  {32'h45239164, 32'h44015a7a, 32'hc2a1766e},
  {32'hc4197a94, 32'h450436a5, 32'h438d0a3e},
  {32'h44aff2ea, 32'hc4bbd9be, 32'hc34f80d5},
  {32'h44d199c5, 32'hc370b13b, 32'h42f44e89},
  {32'h4480cb6d, 32'hc358fae2, 32'h43970f61},
  {32'hc48dbe03, 32'hc42fae55, 32'h44709cb1},
  {32'h430c6547, 32'hc494376a, 32'hc387d391},
  {32'hc2ca7cc4, 32'h4471397e, 32'hc22dd24a},
  {32'hc3212bc8, 32'hc41806be, 32'hc5229800},
  {32'hc46cd7e4, 32'h439e9c2e, 32'h41f583cc},
  {32'h451d478e, 32'hc395f6ae, 32'hc3cfa133},
  {32'hc392fd5b, 32'h445d1194, 32'h44b20e49},
  {32'hc239c530, 32'h432eec9f, 32'hc257ea53},
  {32'hc42b064a, 32'h444edc19, 32'h44a0b2d3},
  {32'h44914217, 32'h420627c6, 32'hc4afbd69},
  {32'h444cbf46, 32'h41c5f35c, 32'h43ed0355},
  {32'hc3bc0a28, 32'hc42bed66, 32'hc4c7d769},
  {32'hc43d8309, 32'h44b3c268, 32'h421db37d},
  {32'h44d45191, 32'hc370d7a4, 32'hc367e3d5},
  {32'hc5131ab8, 32'h4459feef, 32'hc28db208},
  {32'h4551b4f3, 32'hc3e72234, 32'hc404a236},
  {32'h44920360, 32'hc2577ab1, 32'hc356398f},
  {32'hc459d104, 32'h438e22e8, 32'h44fb592b},
  {32'h452495e5, 32'h42a00b11, 32'h441d2b47},
  {32'h4215f300, 32'hc546c29e, 32'hc3f61739},
  {32'h44961a27, 32'h446802f0, 32'h42a6bdee},
  {32'hc4ee41a0, 32'h423f4292, 32'hc327d623},
  {32'h449af792, 32'h44cbd462, 32'hc31b4586},
  {32'hc42912b2, 32'hc4c9220f, 32'hc41b9d47},
  {32'h439ae203, 32'h4425c2bc, 32'hc1231d83},
  {32'hc4a758bc, 32'h4321b348, 32'h4371cd14},
  {32'h44f5a6ad, 32'h41ca0c7f, 32'hc4805844},
  {32'h441cb328, 32'hc4361b7f, 32'hc35a4624},
  {32'h4384eb3f, 32'h43c41b7e, 32'h44db2017},
  {32'hc486b2e8, 32'hc3c49928, 32'hc1c039d1},
  {32'hc302fb88, 32'h4432106a, 32'hc20bf287},
  {32'hc49bbc57, 32'hc42b1eda, 32'hc4bc8d7f},
  {32'h4514d6e6, 32'h439cfe6e, 32'h41977a1b},
  {32'h43780e4b, 32'hc3469f84, 32'hc4c77384},
  {32'h4555ad36, 32'hc34fc87b, 32'hc09d9524},
  {32'hc54e58f6, 32'h4377c2f4, 32'hc2a2cab8},
  {32'h44bd9b8b, 32'h43838117, 32'hc2f82af9},
  {32'hc40c9b28, 32'hc41171d3, 32'hc480f039},
  {32'h44f19f85, 32'h430f2166, 32'hc12c3947},
  {32'h448fbbfa, 32'hc38468bf, 32'hc30500ce},
  {32'h449ff100, 32'h448220d0, 32'h445d9768},
  {32'hc53fe9c6, 32'h438473d9, 32'hc40b85bc},
  {32'h438a2154, 32'h44d8e760, 32'h4213ae3b},
  {32'hc40d9ab3, 32'h43ed2cb2, 32'h43e670ac},
  {32'hc39df9f1, 32'hc50df778, 32'hc2892ea7},
  {32'h44f97ec4, 32'h445f3819, 32'h4418de58},
  {32'hc4ed7432, 32'h43f87678, 32'hc3763cd8},
  {32'h4466b1e1, 32'h44928739, 32'hc40d5597},
  {32'hc45c2cd1, 32'hc2b34d99, 32'h43d22e2a},
  {32'h4521a2f2, 32'h43557f24, 32'hc32ef462},
  {32'hc492e491, 32'h43e9b24e, 32'hc27aba67},
  {32'hc36fdbe0, 32'hc39884f9, 32'h43cb659f},
  {32'h440cc79d, 32'hc4472e8d, 32'h433f0069},
  {32'h43567b1f, 32'h444a108d, 32'hc514e464},
  {32'hc4cd834d, 32'hc3983545, 32'h4457acf7},
  {32'h44561e24, 32'h43857b42, 32'hc21c8c0f},
  {32'hc404e336, 32'hc4ea415c, 32'h4444746b},
  {32'h43897616, 32'h437bacea, 32'hc470a1d4},
  {32'h44eade19, 32'hc21be304, 32'h43440ed2},
  {32'h4414d348, 32'hc3edbd4e, 32'hc45495cc},
  {32'hc4267847, 32'hc4836ece, 32'hc42134c7},
  {32'h4423bb35, 32'h42760ba5, 32'hc3e2d4cb},
  {32'hc4de8bf2, 32'hc442eb72, 32'h4403582d},
  {32'h43c48de2, 32'h44388fc4, 32'hc487e198},
  {32'hc353bd6a, 32'h4210cc2d, 32'h445d8a10},
  {32'h44c1de2c, 32'h445edb29, 32'hc36038ce},
  {32'hc42a1b19, 32'hc4b83b7e, 32'h438a3774},
  {32'h453c9cf8, 32'h43ad7c0e, 32'hc3d977db},
  {32'hc58c4920, 32'h42c85530, 32'h4305b68f},
  {32'h455c9d23, 32'h4414c70e, 32'hc34e5a91},
  {32'h44befc94, 32'hc45f36fc, 32'h418d52f5},
  {32'hc5024e7b, 32'hc2d0030e, 32'h440f9d45},
  {32'h43988952, 32'hc35baca0, 32'h441082cd},
  {32'hc300e2cf, 32'h45498787, 32'h43119db4},
  {32'h43d5a831, 32'hc45f02d2, 32'hc2fb5311},
  {32'h4384677d, 32'h4509cb73, 32'hc3579bf3},
  {32'h44996bc7, 32'h4321c743, 32'hc352f6e6},
  {32'hc3c43ff0, 32'hc14792eb, 32'h439b3125},
  {32'hc492590d, 32'hc3991128, 32'hc1835ef0},
  {32'hc49616c9, 32'h44408b4a, 32'hc450722f},
  {32'h42e64ca0, 32'hc448ad20, 32'h44f262ed},
  {32'h3ecce240, 32'h441f1d1f, 32'hc19cda3b},
  {32'hc394a6a7, 32'h40e9a89d, 32'hc34c229f},
  {32'hc39a7f8c, 32'h44c309d0, 32'hc36b53a2},
  {32'hc4a60cbd, 32'hc280aad4, 32'hc2c07656},
  {32'hc354094c, 32'hc3bea666, 32'hc56cd262},
  {32'h4463e9a2, 32'hc44ac69f, 32'hc3940e53},
  {32'h45064349, 32'h42b79e1e, 32'h439f6185},
  {32'h433cc4dd, 32'hc52cc6db, 32'hc388c0eb},
  {32'hc3b8aa00, 32'h44e4810a, 32'hc460804b},
  {32'h450854c4, 32'h4430e7ea, 32'hc2a9ad12},
  {32'hc500fe15, 32'h4394b794, 32'hc48ebd9c},
  {32'h449c7140, 32'hc23a60fe, 32'h441229c8},
  {32'hc4f235f3, 32'h42edb5c8, 32'h42974422},
  {32'h4480d14e, 32'h4392cbf3, 32'h44c1d879},
  {32'hc538d70d, 32'hc396ba3b, 32'hc484c946},
  {32'hc4588c19, 32'h433b1c24, 32'h43bc753e},
  {32'h43264675, 32'h445e1c00, 32'hc4f13d1b},
  {32'h440db77c, 32'h446bd501, 32'h44abb72e},
  {32'hc3a0eff2, 32'h4407d1c4, 32'hc4631766},
  {32'h4409a282, 32'h436e590f, 32'hc49342e3},
  {32'h4494a513, 32'hc4e814b9, 32'h438b133a},
  {32'hc3890d8b, 32'hc2ed3c62, 32'hc4fe423b},
  {32'hc323d398, 32'hc3909430, 32'hc331d03f},
  {32'hc4533a82, 32'h438d8211, 32'hc4bf4d12},
  {32'h4472c2bb, 32'hc4538509, 32'hc3ff9085},
  {32'h44a7b1d7, 32'hc385c439, 32'h44abcad2},
  {32'h439e5f3e, 32'hc441269a, 32'hc529cb44},
  {32'h438b0c32, 32'hc4a2ac3e, 32'h44717bf6},
  {32'h43b88890, 32'h42b06e23, 32'h43a854dd},
  {32'hc4f238bc, 32'hc2e7f183, 32'h429d05f2},
  {32'h44fe7d15, 32'hc2ad9b21, 32'hc3e11b9e},
  {32'hc3d65aa2, 32'h44be8a6d, 32'h4383bf43},
  {32'h4550bacc, 32'h4196b7b4, 32'hc365cf9a},
  {32'hc457820c, 32'hc255f788, 32'hc4cdbe7d},
  {32'h448b155b, 32'hc40ef5e1, 32'h43a782be},
  {32'hc550ecc0, 32'h424989e8, 32'hc3fb7b9b},
  {32'h44fcda91, 32'hc37b95f2, 32'h43c9606f},
  {32'h4426a19f, 32'hc3762f82, 32'hc38ca858},
  {32'h45335d42, 32'h43875026, 32'h4394ea05},
  {32'hc4ae1070, 32'h44b1f50a, 32'h4395aec7},
  {32'h44869a81, 32'h4185e019, 32'hc23ee4a9},
  {32'hc53a0b8f, 32'hc2538bfd, 32'hc3ef4d2b},
  {32'hc41d1e04, 32'hc5015c81, 32'h432613c0},
  {32'hc4b7030d, 32'hc3791380, 32'hc3c7b9c6},
  {32'hc349bb93, 32'h44e19335, 32'hc4d4d026},
  {32'hc4349fbe, 32'h44b8510b, 32'h4438dcf2},
  {32'hc4d99ec4, 32'h4412fd27, 32'h443a4ba0},
  {32'h43bfe6fb, 32'h45355eee, 32'h43e6467d},
  {32'hc4b622c0, 32'h4299bc6d, 32'h43a8efe1},
  {32'hc3519f20, 32'h452e26c7, 32'hc38f77cb},
  {32'hc4c4d8f6, 32'hc3c910d6, 32'h441c9f49},
  {32'hc42a62c4, 32'hc2d9ce14, 32'hc43aab78},
  {32'h43c0d6e8, 32'h4480bdcf, 32'hc37abb8c},
  {32'hc47fc0e8, 32'hc3ecd4c6, 32'h44738aa5},
  {32'hc3d0acf3, 32'h44b47767, 32'hc5056c9f},
  {32'h448c3860, 32'h43fa2a62, 32'hc427f05f},
  {32'hc4a0d90d, 32'hc49343ee, 32'hc3bd58d4},
  {32'h43f2d792, 32'h446b0bbc, 32'h436f8442},
  {32'hc4517327, 32'hc4065412, 32'h45003eb4},
  {32'h443ddc1b, 32'h44acb1f9, 32'hc420f4bc},
  {32'hc3af7474, 32'hc4c8fc42, 32'hc257f0d2},
  {32'h4518058c, 32'h428dbbfb, 32'hc33f98d1},
  {32'hc532311b, 32'hc311d5fc, 32'hc3014e68},
  {32'hc49f8294, 32'hc1d46a7e, 32'h4354f9d3},
  {32'hc4d125f3, 32'hc4aba95f, 32'h436b0faa},
  {32'h4390e740, 32'h4285fd73, 32'h42d50648},
  {32'hc513b296, 32'h432817a2, 32'h43963354},
  {32'h43493920, 32'h4509f9bd, 32'hc366917f},
  {32'h427826f0, 32'hc52c44aa, 32'hc3378e34},
  {32'h443c147a, 32'h4385d3e0, 32'hc3f016ca},
  {32'hc4685d1f, 32'h439c1a81, 32'hc25e3fac},
  {32'hc502da0a, 32'hc39360a0, 32'h430fd820},
  {32'h43eff73e, 32'h448138a5, 32'h43b6b931},
  {32'h4488e17c, 32'hc2c53215, 32'hc34d3694},
  {32'h445ca397, 32'h4332bbfe, 32'h4445164e},
  {32'h40275700, 32'hc3e485f4, 32'hc4b3ae7b},
  {32'hc4109333, 32'hc35c855a, 32'h4442ff50},
  {32'hc40d7802, 32'hc423c532, 32'hc503539b},
  {32'h44258a33, 32'h43cb4ffb, 32'h4518ef2b},
  {32'hc3abb565, 32'hc4eed7c0, 32'hc36a8aca},
  {32'h438c8dbc, 32'h43a052d3, 32'h43872c2f},
  {32'hc47794c5, 32'h42d5b449, 32'hc46c64ae},
  {32'h448d14fc, 32'h440585f6, 32'h42fca961},
  {32'hc4f748b0, 32'hc3c9fb4d, 32'h4386e4f4},
  {32'h4369413f, 32'h43309e7d, 32'h4507c70d},
  {32'hc435086f, 32'hc463ebe1, 32'h4208af3c},
  {32'h43e871ef, 32'h43e97b9a, 32'h442fe65d},
  {32'hc3defdc7, 32'hc419262a, 32'hc4ca0806},
  {32'h447876ec, 32'hc2ca246c, 32'h41ce2c16},
  {32'hc3e91ea5, 32'hc501af01, 32'hc3a851b9},
  {32'h44175196, 32'h45693071, 32'hc3970b2f},
  {32'hc4413d71, 32'hc337081b, 32'hc3ba5b87},
  {32'h454c5938, 32'h4416c268, 32'hc3202eee},
  {32'hc49ac3d9, 32'hc4842e24, 32'h434206a1},
  {32'hc38ffa48, 32'h43d3a4e0, 32'hc39fa31a},
  {32'hc4ebde0b, 32'hc379d323, 32'h433b06a6},
  {32'h4589d2cd, 32'h43a68e20, 32'h438f243a},
  {32'h42ece1a9, 32'hc5015129, 32'hc3a1caa5},
  {32'h4335086c, 32'hc3beaa1c, 32'h44f263fc},
  {32'hc40a64f3, 32'hc4bbc197, 32'h43184bc1},
  {32'h431ef26c, 32'h4164cba2, 32'h44c4d23b},
  {32'h446c0900, 32'hc3596cd4, 32'hc407a1a9},
  {32'hc512b34f, 32'hc3419602, 32'hc2e981d3},
  {32'hc3a6474f, 32'hc4f0b62f, 32'hc4ec1552},
  {32'hc42ddee0, 32'h442b85b2, 32'h44adb43e},
  {32'hc36c8fc0, 32'h4268bdd6, 32'hc4e5abbb},
  {32'h433065dc, 32'h449c337c, 32'h436dd716},
  {32'hc3b0936b, 32'h44d13b3b, 32'hc4cefe47},
  {32'h433968a8, 32'h43427d26, 32'h42b02ce4},
  {32'hc123d400, 32'hc4bbd87a, 32'hc44a3a42},
  {32'hc1fa8780, 32'h43cc61e3, 32'h4528b1a0},
  {32'h43a06904, 32'hc3923078, 32'hc4aa0129},
  {32'hc442fe06, 32'h44854d06, 32'h447441ee},
  {32'hc39a5ac0, 32'hc4ac6327, 32'hc56a1739},
  {32'h4489942d, 32'hc34dfb66, 32'h4419cbf6},
  {32'h42dd365d, 32'hc545c3ba, 32'h41d48324},
  {32'hc403656c, 32'h4512d820, 32'h436934eb},
  {32'h449b5004, 32'hc372da53, 32'hc0964ccc},
  {32'hc41227a6, 32'h454b6076, 32'hc3332ae9},
  {32'h44accbad, 32'hc53a5f53, 32'hc3971770},
  {32'h44246ed6, 32'h448bfe0c, 32'hc0f88aa4},
  {32'h4521916c, 32'h43296402, 32'h4312744c},
  {32'hc508c68d, 32'hc3afe271, 32'hc2ab6d40},
  {32'h44909499, 32'hc4058974, 32'h4298eb82},
  {32'h448f14b4, 32'hc2f3c93c, 32'h4401cd25},
  {32'hc496b7b1, 32'h43e1e9d4, 32'hc4b6cffa},
  {32'h45039c7d, 32'h43c16f6b, 32'h441f46fc},
  {32'h44e3f033, 32'h43b0db55, 32'hc2fe3058},
  {32'h44468e18, 32'hc51be480, 32'h4290c494},
  {32'h41440a00, 32'h443366b7, 32'hc3645f5e},
  {32'h4462b508, 32'hc340924f, 32'hc3e16220},
  {32'hc524548b, 32'h438a2962, 32'hc22d763a},
  {32'h44a08527, 32'hc41a405f, 32'h4458e275},
  {32'h44c25062, 32'h44476498, 32'hc3609614},
  {32'h43c5d394, 32'h43721560, 32'hc40a3c70},
  {32'hc526ced0, 32'hc2917952, 32'h4400ea13},
  {32'h4421ff3c, 32'hc4b358d2, 32'h4380a91d},
  {32'h42828d48, 32'hc3be7be4, 32'h45461fc8},
  {32'h432b9500, 32'hc51daba7, 32'hc15e0564},
  {32'h439000bf, 32'h43627be8, 32'h44213487},
  {32'h449a8378, 32'h440784ba, 32'h41ad1f33},
  {32'hc39defa6, 32'h44b9ed4d, 32'h43455161},
  {32'h444cf26a, 32'h41b29b47, 32'hc31da465},
  {32'hc4bbd49c, 32'h40141406, 32'h4424ffcf},
  {32'h440722a0, 32'hc41e0f7b, 32'hc4c24566},
  {32'hc53782f2, 32'h438b8c63, 32'h4336519b},
  {32'h4358eb8c, 32'hc4f8f320, 32'hc32e5edb},
  {32'hc3e00a18, 32'h450a2745, 32'h44170c1b},
  {32'h44d359dd, 32'hc0ac22f2, 32'hc37d1ec8},
  {32'h41945ea0, 32'h441eb2c0, 32'h4544fcf4},
  {32'h44648f4a, 32'hc4b309ad, 32'hc3db6bb1},
  {32'h4492018c, 32'hc37a6eec, 32'hc4692492},
  {32'hc433ee80, 32'hc36498e2, 32'h45140f1f},
  {32'hc41fab13, 32'h430b8a76, 32'h420e6a2a},
  {32'hc2ef2ae0, 32'hc41f5129, 32'hc2d2ba94},
  {32'h447b2236, 32'h444ed64d, 32'h43f50aeb},
  {32'h44a0b966, 32'hc3ded8d9, 32'hc2bd131e},
  {32'h4546c064, 32'h43ec1512, 32'hc31c635a},
  {32'hc4a25a64, 32'hc4540dfa, 32'h4395f1b9},
  {32'h445a8078, 32'h4484e888, 32'hc375e647},
  {32'hc410f30b, 32'hc2eaf8f5, 32'h447f1f67},
  {32'h45022bb9, 32'hc3e9ffd5, 32'h43033441},
  {32'hc48e6743, 32'h4450067a, 32'hc459b0d8},
  {32'h43ba46e8, 32'hc20c4b04, 32'h452f15d3},
  {32'hc4ed25cb, 32'hc401fe04, 32'hc3d0c32a},
  {32'h42f75b48, 32'h4430acea, 32'h4320d401},
  {32'hc5029c29, 32'hc3adf85b, 32'hc4587dd0},
  {32'h44356e4c, 32'h43ef39ef, 32'h44dc0362},
  {32'hc413efc7, 32'hc35b1a98, 32'hc2d0da4c},
  {32'h448f9606, 32'hc4083290, 32'h43196685},
  {32'hc28be080, 32'hc32dc951, 32'hc4b2cad2},
  {32'h44d87edf, 32'h4423adfa, 32'hc3ff0ea2},
  {32'h42eefd18, 32'hc401c3c2, 32'hc52daec8},
  {32'hc2f48e88, 32'hc3e56a89, 32'h451bb6d4},
  {32'hc4c0bd37, 32'hc40105eb, 32'h43887c0f},
  {32'hc4027a04, 32'h43daefd5, 32'h445f58db},
  {32'hc4e961e6, 32'hc4a63086, 32'hc3bfb653},
  {32'h43243eb8, 32'hc21ee011, 32'h44f519d2},
  {32'hc4449345, 32'hc39c223c, 32'h439abc7a},
  {32'hc4911b76, 32'h42d726a4, 32'hc491fdbe},
  {32'h42a37100, 32'h450f4012, 32'hc3496aca},
  {32'hc52d36c3, 32'h43860491, 32'hc30bb2b2},
  {32'h44236e22, 32'h4301b402, 32'hc34d1667},
  {32'hc401456a, 32'hc5018cb4, 32'hc392b34e},
  {32'h44c8bc0c, 32'h42f9ed1b, 32'hc426059e},
  {32'hc52feb5c, 32'h435d1d0f, 32'hc3948c87},
  {32'h43d34d64, 32'h445e4968, 32'h43fb6546},
  {32'h44dcf38f, 32'hc38c2a86, 32'hc32b25f2},
  {32'h43de2a70, 32'h441262ba, 32'h448b5d3b},
  {32'hc487d1af, 32'hc40c4645, 32'hc3c377cf},
  {32'h44953d76, 32'h442a22c8, 32'h41511e8f},
  {32'hc35e35ec, 32'hc46b6f5b, 32'h44565959},
  {32'h43621ba6, 32'h45091703, 32'hc39a29dd},
  {32'hc403d40e, 32'hc387bff8, 32'hc3e51102},
  {32'h448a0a34, 32'hc3e0bb8e, 32'hc41ad06a},
  {32'hc4e5846c, 32'hc260f1bf, 32'h43628cf9},
  {32'hc4215af2, 32'h429ec2f2, 32'hc445824f},
  {32'hc4b3a752, 32'hc41f00e0, 32'h443212fa},
  {32'h4428472d, 32'h439803dd, 32'hc5156e9f},
  {32'h4448805b, 32'hc41774ea, 32'h4365eded},
  {32'h44f36082, 32'h4401f2b1, 32'hc46501fb},
  {32'hc4a99e80, 32'hc3b72b69, 32'hc0e2b6fa},
  {32'hc4ab141c, 32'hc1e2fd46, 32'hc38ba2d5},
  {32'hc38acf35, 32'hc209e17b, 32'h452655a8},
  {32'h44923430, 32'h4353d6fb, 32'hc4d4f982},
  {32'h444e4f98, 32'hc50a270d, 32'hc324e4ce},
  {32'hc5334056, 32'h440e0576, 32'hc33cd5bf},
  {32'h45145e0a, 32'h427abff7, 32'h4326dc7a},
  {32'hc4e1ca87, 32'h449e3906, 32'h442ba015},
  {32'h445bde08, 32'hc4a5543b, 32'hc3dec6b0},
  {32'hc39c01f5, 32'h442b0513, 32'hc3a90038},
  {32'h44ff077e, 32'h429963e6, 32'h43a5c9a7},
  {32'hc5167850, 32'hc2f7861f, 32'hc28393bc},
  {32'hc4552616, 32'hc44a6fe3, 32'h42bde4ca},
  {32'h4287e738, 32'h44eec3e7, 32'hc41110dc},
  {32'h43ecd1e3, 32'hc34bbcde, 32'h44b487f0},
  {32'h430fae24, 32'h4381febb, 32'hc4d1af32},
  {32'h443c7100, 32'hc49b5538, 32'h443820b7},
  {32'hc4ad5a98, 32'h446d7754, 32'h41f66546},
  {32'hc43d5b41, 32'hc4210dce, 32'hc3b1ae5a},
  {32'hc3f2717a, 32'hc3495c81, 32'hc4c793ca},
  {32'h44c1dfd9, 32'hc49d76eb, 32'hc44daab4},
  {32'h44cb3242, 32'h44259ddb, 32'h438d4702},
  {32'h45062572, 32'hc4940f0e, 32'hc3b0fc99},
  {32'hc39e7bf4, 32'h4493c1b8, 32'hc5458482},
  {32'h43960de5, 32'hc4c0e834, 32'hc30cd16f},
  {32'hc44ca1c2, 32'h44c616e8, 32'hc41a77cd},
  {32'h43b74b7e, 32'hc37ed619, 32'h44b6cc58},
  {32'h4403bf0e, 32'hc23450d1, 32'hc49a7171},
  {32'h453721ee, 32'h43120c3c, 32'h43d91442},
  {32'hc5069d6d, 32'hc357e03c, 32'hc444147e},
  {32'h450ba042, 32'h4221b725, 32'hc23ad5df},
  {32'hc4edce2a, 32'hc3d458f7, 32'hc3a5fac1},
  {32'h445d5269, 32'hc4a7197f, 32'h44995248},
  {32'h437dcfb2, 32'h43d95b20, 32'hc429b18b},
  {32'hc4c98172, 32'h4387dd08, 32'h421b2716},
  {32'h440f812d, 32'hc39571b7, 32'h4541a53c},
  {32'hc2ed496b, 32'h450cb98d, 32'hc4075791},
  {32'h44b269fc, 32'h42dd3f1e, 32'h43f1807d},
  {32'hc4310f4c, 32'h439226fa, 32'hc5475f35},
  {32'h4494fe32, 32'h4227fce2, 32'h446f2b1e},
  {32'h443182bd, 32'hc4219cbf, 32'h449f3405},
  {32'hc4c5d4ee, 32'h43905eaf, 32'hc414af99},
  {32'h43beb907, 32'hc4e28db2, 32'h43aa26bc},
  {32'h43776dd3, 32'hc4af33b1, 32'h4423b955},
  {32'h42ac7ee2, 32'hc115d8f2, 32'hc533c4c3},
  {32'hc353ee50, 32'hc2a30e36, 32'h44922be8},
  {32'h4492d73e, 32'h440a3e20, 32'hc23ed2da},
  {32'h44289c74, 32'hc32c74ca, 32'h44cc3186},
  {32'hc2eea308, 32'h42be21c5, 32'hc50e93e8},
  {32'h435eed88, 32'hc106c75c, 32'h440f1d13},
  {32'hc4a18a09, 32'hc422e5b8, 32'h430cbf0a},
  {32'h454764ae, 32'h4437dbf4, 32'hc38d5818},
  {32'hc4a4cf18, 32'h43b69222, 32'hc41e1439},
  {32'h438162b0, 32'hc5043481, 32'hc3ada5b0},
  {32'hc38035b4, 32'h45001b6c, 32'hc09142e4},
  {32'h44d2b359, 32'h43f963db, 32'h43f6b1d0},
  {32'hc4f9a84c, 32'h44a8a0b1, 32'h426f847e},
  {32'h44f51fea, 32'hc4365645, 32'h43d23c6a},
  {32'h440cb1fb, 32'h44079e1f, 32'h441ff3b9},
  {32'h44fbb1f4, 32'hc391ff4f, 32'hc0858dc0},
  {32'hc4944cc5, 32'hc453ea6b, 32'h44433b5b},
  {32'hc41c7617, 32'hc44e7c35, 32'h43dc1ef7},
  {32'h429e3e00, 32'hc2b6a735, 32'hc52487b9},
  {32'h433e379a, 32'hc4c700bd, 32'h41a5c485},
  {32'h435b5c9f, 32'h44fb303a, 32'h42992585},
  {32'h42f7be3a, 32'hc5201f00, 32'h437ea20d},
  {32'hc37c762a, 32'hc2b9bfa9, 32'hc4dc540a},
  {32'h440cdf5e, 32'hc3cd5102, 32'hc31e514e},
  {32'hc48b7a50, 32'hc4b56110, 32'h4491812b},
  {32'h4347e900, 32'hc41b54fa, 32'hc5188475},
  {32'h4442436c, 32'h44413779, 32'hc3b12c22},
  {32'hc49c8ab6, 32'h4239659b, 32'h438e8698},
  {32'hc4997417, 32'h43a2147c, 32'hc43c097a},
  {32'hc3ec077a, 32'h4232bfff, 32'h44206fc7},
  {32'hc351739d, 32'h43890246, 32'hc4b002f7},
  {32'h44a2a547, 32'h42dcc1c7, 32'h43d9e927},
  {32'h449a877a, 32'hc331ec71, 32'hc3032330},
  {32'hc507e5aa, 32'h43258cb3, 32'h4440ed00},
  {32'h44981b5e, 32'h43b0db8e, 32'h436f7f12},
  {32'hc41c37de, 32'hc4914524, 32'hc40f9a62},
  {32'h4397cbad, 32'h45487938, 32'h433ed419},
  {32'hc5050228, 32'hc31af7e1, 32'h43deb8cc},
  {32'h43befd70, 32'h4504ccab, 32'h43832af3},
  {32'hc50cad73, 32'hc47281d5, 32'hc2ee157e},
  {32'h4238606a, 32'h43ec3d30, 32'hc38bad76},
  {32'h436a9d56, 32'hc4401754, 32'h4396a2f2},
  {32'h429d10f1, 32'hc3b12d0d, 32'hc4bea788},
  {32'hbf9dd000, 32'h44af7573, 32'h445dde30},
  {32'h43b0d82c, 32'hc3765ab9, 32'hc44e927c},
  {32'h43dc84d2, 32'h43508bb0, 32'h44bfe1ca},
  {32'hc3dd320d, 32'hc4cec9e4, 32'hc381f519},
  {32'h42ba60ea, 32'hc37a20a1, 32'h45061998},
  {32'h4194048b, 32'h4310cb1f, 32'hc514bec5},
  {32'h45247941, 32'hc1a92f15, 32'h441c6efd},
  {32'hc1f6adae, 32'h438206f4, 32'h4315fcf5},
  {32'h42b638e0, 32'h44a084b4, 32'h4456f59c},
  {32'hc352f7be, 32'h45065658, 32'hc4c24d5a},
  {32'h450403b4, 32'h42ff054f, 32'h4310216d},
  {32'hc41ef5dd, 32'hc3b0ab44, 32'hc3f06890},
  {32'h430f2328, 32'h440840ac, 32'h44c6e911},
  {32'h42bcafe0, 32'hc38517c9, 32'hc5043ff0},
  {32'h4420407d, 32'h448d931d, 32'h43fc29e3},
  {32'hc44e7cba, 32'hc4856e97, 32'hc4a19b7d},
  {32'h4461f255, 32'h43b41a2b, 32'hc2069ee7},
  {32'hc54d5ba9, 32'hc3953c8a, 32'hc2b4c173},
  {32'h446b4190, 32'h44ac480c, 32'h43bc75ad},
  {32'hc3af0aec, 32'hc493d45d, 32'h4308e2be},
  {32'h4544b0a0, 32'h438c2b97, 32'hc2d49d2d},
  {32'hc44b8202, 32'hc4ee19dd, 32'hc2d70a39},
  {32'hc4bb23a8, 32'h43002c50, 32'hc3a200d5},
  {32'hc5137a06, 32'h42e097ea, 32'hc384480d},
  {32'h443ca6dc, 32'h43b3d6f5, 32'h42b8b6b6},
  {32'h43da0a79, 32'h44302c33, 32'hc4b957f8},
  {32'h43dc51b7, 32'h4561495d, 32'h4416ee3c},
  {32'hc3e535be, 32'h41cdd325, 32'hc42d1cde},
  {32'hc404f30e, 32'h451640d3, 32'h43499a01},
  {32'hc2af842b, 32'hc4d870ee, 32'hc4566009},
  {32'hc4f8a668, 32'h4216b90f, 32'h43a360fa},
  {32'h4440b03f, 32'h42c0dd6a, 32'hc462af70},
  {32'hc3d53c9c, 32'h44f7a622, 32'h44c23dd7},
  {32'h43630ff6, 32'hc4a47dd2, 32'hc36a8af3},
  {32'h429bdc90, 32'h4477716f, 32'h4424fea4},
  {32'hc4525f6c, 32'h44a44127, 32'hc5313602},
  {32'h4456611b, 32'hc1a70450, 32'h42e57738},
  {32'hc341feb0, 32'hc34ba0fa, 32'hc0a1dec8},
  {32'hc3ae6cce, 32'h44e575d3, 32'h43f2b791},
  {32'hc45f28b2, 32'hc4853e8e, 32'h4222eec6},
  {32'hc3826f50, 32'h433f441e, 32'h451fbfba},
  {32'hc3d1e42a, 32'hc4829ec3, 32'hc456be0f},
  {32'h42b52ac8, 32'h429c950f, 32'h450754c0},
  {32'h44a0fbc4, 32'hc4a9b8c4, 32'h43e93fd7},
  {32'hc527e8aa, 32'h447df2ac, 32'h4350257a},
  {32'h44ab452e, 32'hc2b9a723, 32'h438799a9},
  {32'h42dbc3d3, 32'h4580caea, 32'h41ec9042},
  {32'h4550fb8f, 32'hc28f9be3, 32'h434677b5},
  {32'h43e6f672, 32'h44cf4e3c, 32'hc307797d},
  {32'h45259d75, 32'hc3a78186, 32'h42b0d4eb},
  {32'hc4b05a17, 32'hc3a60c2f, 32'h438e84e3},
  {32'h451284f3, 32'h42e8896f, 32'hc3b36814},
  {32'hc32f557f, 32'hc31bdb8d, 32'h4447ce0b},
  {32'hc3eda8a0, 32'h431d2c9c, 32'hc5051f5e},
  {32'h44c26cce, 32'h43c77bc3, 32'h4473948e},
  {32'h44725a5c, 32'h434daaa9, 32'h4134f366},
  {32'h43e01418, 32'hc4b9ecde, 32'h43b77727},
  {32'hc2e1f4ec, 32'h453a8470, 32'hc2d852e6},
  {32'h44bef23c, 32'hc0e9f8f0, 32'hc3d35a36},
  {32'hc522c88c, 32'h43f2a19a, 32'h4381c92e},
  {32'h43c0ff10, 32'hc49c6427, 32'hc3c8062b},
  {32'hc43ba587, 32'h416c81d5, 32'hc4195a8b},
  {32'h44858374, 32'h42d81a32, 32'h441b2aea},
  {32'hc42765b1, 32'h4453b02c, 32'h4480d8bb},
  {32'hc12cb000, 32'hc4b36e4e, 32'hc319bede},
  {32'hc51b9d35, 32'h430fc7d6, 32'h40ff47b6},
  {32'h4503b495, 32'hc20a74c7, 32'hc396c2cc},
  {32'h4409f644, 32'h433f56ac, 32'h43b492e7},
  {32'hc39f381a, 32'hc519245e, 32'hc3b58264},
  {32'hc4b90799, 32'h4220d134, 32'hc2841a83},
  {32'h441bfc6b, 32'hc3e8d160, 32'hc3c23987},
  {32'hc502e1eb, 32'hc2ffe7bf, 32'h44554e21},
  {32'h45245b5c, 32'hc38b24a4, 32'hc43c52b4},
  {32'h421ecb38, 32'h444b2e82, 32'h440cfc9c},
  {32'h44b90b38, 32'hc418996d, 32'hc3c99257},
  {32'h43b15d02, 32'h4502d02f, 32'h4448df3c},
  {32'h44a6d258, 32'hc2b05c75, 32'hc3be61ea},
  {32'h430ed31a, 32'h440ad551, 32'h452bd68a},
  {32'h44717b05, 32'hc44992bb, 32'hc4c566c3},
  {32'h44ea8a82, 32'hc37493d5, 32'hc42f2f92},
  {32'hc4886bdc, 32'h4375b769, 32'h44fa3f3d},
  {32'hc444ea62, 32'h43e8c872, 32'hc3383b35},
  {32'h4158f9a8, 32'hc4b856b9, 32'hc296cea8},
  {32'h44563727, 32'h44853041, 32'hc3d91d99},
  {32'hc48a30f6, 32'hc43e49ae, 32'hc3bc8c4a},
  {32'h43056678, 32'h453744d8, 32'hc3136327},
  {32'hc485b610, 32'hc4f60e2d, 32'h43041fd5},
  {32'h43ec2ffa, 32'h4461a58d, 32'h43b39aa9},
  {32'hc48a808a, 32'hc45d07b4, 32'h448542d4},
  {32'h4515689f, 32'hc3a3edda, 32'h431adf37},
  {32'hc4953333, 32'h43767451, 32'h445eed25},
  {32'h4446bb33, 32'h442067dd, 32'h440a8c71},
  {32'hc4ad8c12, 32'hc4b95e55, 32'hc3f1c2b8},
  {32'h441ee1ea, 32'h44305b22, 32'h42be1293},
  {32'hc4362a3c, 32'hc32daa59, 32'hc47c1a1a},
  {32'h432be72a, 32'h4403dd3d, 32'h45328718},
  {32'h44ebec52, 32'hc3e33565, 32'h43778b82},
  {32'h43ffbfd6, 32'h443e29a6, 32'h44a92226},
  {32'hc57ef51e, 32'hc3189108, 32'hc1361c28},
  {32'hc4a9517d, 32'hc2b7b499, 32'h432aaf3e},
  {32'hc40196e5, 32'hc4ec52b1, 32'hc44c929d},
  {32'hc393ec27, 32'h45128161, 32'hc3a7c315},
  {32'hc4a1e707, 32'hc408014d, 32'h43a06c56},
  {32'h40331300, 32'h449ec78c, 32'h44678b82},
  {32'hc4f590d5, 32'hc46df550, 32'hc4415b6c},
  {32'hc4d720f6, 32'h43a52007, 32'h428c2f85},
  {32'hc465bd32, 32'h443074a3, 32'h43af2540},
  {32'hc51bca40, 32'hc38c3f09, 32'h42dec7af},
  {32'h448d8a55, 32'h44853adf, 32'h43be41ea},
  {32'hc4fb530e, 32'hc343978b, 32'hc31e68cd},
  {32'h43f3a07d, 32'h44f6efe0, 32'hc37d7ab1},
  {32'hc4d05c98, 32'h42e28208, 32'h43890580},
  {32'h45559d6a, 32'hc4027ff0, 32'hc3d9d4ed},
  {32'hc48abdc3, 32'h43d6980a, 32'hc3329b2a},
  {32'h456006bf, 32'h43c68fcf, 32'h43fc2c19},
  {32'h4378335c, 32'hc447e3b1, 32'h43d17073},
  {32'h4458c5e0, 32'h44902a67, 32'h438f97aa},
  {32'hc486254a, 32'hc38d6ec0, 32'hc3a9cf20},
  {32'h448c06bf, 32'h44158bfd, 32'hc4330fa8},
  {32'hc4405cba, 32'hc4059877, 32'h43d76105},
  {32'h44eeb7f8, 32'h442413b1, 32'h42eb3d81},
  {32'h44055230, 32'hc2c18712, 32'h44823f16},
  {32'h4521bd54, 32'h42f96592, 32'hc11f1755},
  {32'h42a6ccf6, 32'hc312b085, 32'h44d4954c},
  {32'h45296327, 32'hc2588884, 32'hc39fbe34},
  {32'hc425f1f0, 32'hc48214ff, 32'h44e57a10},
  {32'h447f001d, 32'h448e676a, 32'hc5000eeb},
  {32'h422d61d0, 32'hc4480c24, 32'hc45d784b},
  {32'h44271fb4, 32'h4518100d, 32'hc1a08997},
  {32'hc4e23e39, 32'h4341f15e, 32'h43ba613d},
  {32'h45647dbe, 32'h442436b4, 32'hc374c42d},
  {32'hc488de6b, 32'h4465a571, 32'h44e4bce2},
  {32'h428ce6dc, 32'hc38b272c, 32'hc51624f2},
  {32'h431a7d14, 32'hc54883a9, 32'hc3a7f350},
  {32'hc281bafc, 32'h44c6d457, 32'h44130ffd},
  {32'hc4b218cc, 32'h438c38a1, 32'hc3815995},
  {32'hc4442a19, 32'h451efab4, 32'hc30b8ad4},
  {32'h44a2dfc4, 32'hc2f53485, 32'hc39cbea2},
  {32'h448684a6, 32'hc391b5f2, 32'hc30e37f5},
  {32'h4355345c, 32'hc42688f0, 32'hc385a579},
  {32'hc5332550, 32'h43c40616, 32'h43db38b2},
  {32'h44c205c4, 32'h43d0eb8f, 32'h440ebab5},
  {32'h43b67600, 32'h4474b302, 32'hc253b807},
  {32'h43543a90, 32'hc5251b47, 32'hc28043ce},
  {32'hc3680254, 32'h43697efb, 32'hc4b33fe1},
  {32'h44a8ed06, 32'hc43ec5c2, 32'h43c534a2},
  {32'hc3c21f3f, 32'h4384b12d, 32'hc48fce91},
  {32'h44588ab6, 32'hc3f43fe4, 32'h43e29a84},
  {32'hc4990c26, 32'h441d3c84, 32'h432dbb96},
  {32'h432c1564, 32'h432f3f39, 32'h4510ac0f},
  {32'hc4f6de84, 32'h43a3815a, 32'h42b72f98},
  {32'h453ba356, 32'hc43dad24, 32'hc4171819},
  {32'hc48bb382, 32'h44156d1c, 32'hc44c8678},
  {32'h44b0a254, 32'hc3d222c0, 32'h44057142},
  {32'hc3c999c8, 32'h4529338b, 32'h43716b59},
  {32'h451e5e3b, 32'h43940a99, 32'h4361a9d0},
  {32'h42e7f9ef, 32'h432a3972, 32'hc44b7e44},
  {32'h439c4868, 32'h43591355, 32'h4514c940},
  {32'hc55bf212, 32'hc351bd02, 32'hc206e812},
  {32'h44e3181a, 32'h4199e809, 32'h432611e6},
  {32'hc46ca080, 32'h44066921, 32'hc37c3e58},
  {32'h3fe77d9a, 32'h441df4bd, 32'h452db6df},
  {32'h44738e02, 32'h439036e1, 32'hc40c4cfe},
  {32'hc3777268, 32'hc2b40501, 32'hc4bf73b7},
  {32'h44197fa4, 32'h434b19ed, 32'h449feb32},
  {32'hc4b61155, 32'h434fc194, 32'hc44a2a21},
  {32'h43d7a4c1, 32'h43a599a6, 32'h44c85153},
  {32'hc4f32d2e, 32'h43a221e2, 32'hc488db94},
  {32'h44b819ee, 32'hc43deabb, 32'h43d6f47e},
  {32'hc317f83a, 32'h44dbb189, 32'h44e25beb},
  {32'hc50c49cf, 32'h449f817b, 32'hc4927e7a},
  {32'h452a2dec, 32'hc2c4cda2, 32'hc4310805},
  {32'hc323ac7f, 32'hc3c12863, 32'h44290a44},
  {32'hc27bb569, 32'hc2965afa, 32'hc4e6a846},
  {32'h43f7ab68, 32'hc48d8e44, 32'h43f4854e},
  {32'h44e1eeb3, 32'hc3f0a04f, 32'hc3296bfd},
  {32'h43d5da80, 32'hc4606ea4, 32'hc429ad15},
  {32'h42d0847a, 32'h44c03697, 32'hc4050a16},
  {32'hc4eec9ee, 32'h43a9a5e1, 32'h43de25b5},
  {32'hc51c6563, 32'h43d80a55, 32'h42e07b74},
  {32'h453bfb0a, 32'h4400a68b, 32'h43aa6188},
  {32'h43d16c0a, 32'hc36f4353, 32'h4334448b},
  {32'h433044f8, 32'hc4f91179, 32'hc2858c91},
  {32'hc30dc51c, 32'h455a25f4, 32'h419375cf},
  {32'h42fe8160, 32'hc468b749, 32'h4384cb94},
  {32'hc4e26f46, 32'h44832fd2, 32'hc409f901},
  {32'h443cfe80, 32'hc4d65970, 32'h439d2b73},
  {32'h443f7644, 32'hc488cb51, 32'h43d6c24e},
  {32'h430ddfce, 32'hc4636c99, 32'hc44ca487},
  {32'hc3bf637e, 32'h443160c1, 32'h44dc10a3},
  {32'hc3d3fde2, 32'hc490d128, 32'h43c53f98},
  {32'h42d59c1b, 32'h45358bf8, 32'h43219876},
  {32'h45120f88, 32'hc2bcc399, 32'h42ea650b},
  {32'hc2da555a, 32'h43967211, 32'hc4bb4943},
  {32'hc353b750, 32'h42d6be55, 32'h4519bb6c},
  {32'h42018188, 32'h433afb50, 32'hc4f7b1da},
  {32'h44ebb4ca, 32'hc391225d, 32'h43109f57},
  {32'h44093a73, 32'h440e1c72, 32'h4532c975},
  {32'h440e12b4, 32'hc4c8893a, 32'hc4e10df6},
  {32'h4457181a, 32'h43c7844e, 32'hc4aa0af6},
  {32'hc294d2b0, 32'hc5121df5, 32'hc210db0c},
  {32'h43b8f610, 32'h44b2b69f, 32'h434bdffb},
  {32'hc38a5674, 32'h4448b637, 32'h452f93ff},
  {32'h452b5e3f, 32'h434beace, 32'hc2613d1c},
  {32'h441a2716, 32'hc41b3fee, 32'h439423de},
  {32'h44d0fca0, 32'h43433b7c, 32'hc422d6d7},
  {32'hc5774360, 32'hc36d1ae8, 32'hc2c22a50},
  {32'h4559ffb5, 32'h4397ec59, 32'hc35d2bae},
  {32'hc40b42f8, 32'hc48a16ce, 32'h42845a33},
  {32'h4581f252, 32'h42ffcad3, 32'h43d96f97},
  {32'hc4352d43, 32'h432440a9, 32'h43cb84f6},
  {32'h442cb315, 32'h452877c4, 32'hc3472521},
  {32'hc42d3dfe, 32'hc4b4a786, 32'hc3b7ba98},
  {32'h43aeb7da, 32'h44bca0a2, 32'hc35994e8},
  {32'h448c7d8c, 32'hc4a41de5, 32'h439e362a},
  {32'hc43b5ada, 32'hc2aa60cc, 32'hc4a6b8c3},
  {32'hc23a17a1, 32'h450e0ba1, 32'hc38da892},
  {32'h4337c185, 32'hc38aa691, 32'hc4a17bfb},
  {32'h41b3a2e8, 32'h45119ef1, 32'h41987377},
  {32'hc428cf29, 32'hc447cd71, 32'hc4d34d04},
  {32'h428c0b50, 32'h433beacf, 32'h448342a0},
  {32'hc4c4d866, 32'hc3ef8407, 32'hc35fff24},
  {32'h43b6d734, 32'h43efd850, 32'h448bfb66},
  {32'h443c764e, 32'h43a7f63e, 32'h430db1bc},
  {32'hc26bca05, 32'hc2262d18, 32'h445c676a},
  {32'h433b78e3, 32'hc411bded, 32'hc3e8a5ec},
  {32'h43695c71, 32'h44e20ea8, 32'h428f43c1},
  {32'h4368f050, 32'hc4568b68, 32'hc1cabc96},
  {32'h438bcb18, 32'hc3e9de75, 32'h4414dda1},
  {32'hc4d6e34e, 32'hc33f0efd, 32'h4301a850},
  {32'h42dbd629, 32'h43fa4f4a, 32'h450cb81e},
  {32'hc15bc900, 32'hc2aa8daa, 32'hc486545c},
  {32'h4409c949, 32'h432775a4, 32'h43c74380},
  {32'hc5322e69, 32'hc4614697, 32'hc35549a1},
  {32'h44ac74ac, 32'h4489e635, 32'h43e52ff9},
  {32'hc46bf50b, 32'h43320fd9, 32'hc3abaaf2},
  {32'h441b14fe, 32'h4504041b, 32'h440309ad},
  {32'hc49344cf, 32'hc44be8f1, 32'hc2b302d1},
  {32'h44a54336, 32'h43d9210a, 32'h43b2172f},
  {32'hc4c131de, 32'h422ba2bb, 32'hc2c70fdb},
  {32'h4352baa0, 32'hc2b84920, 32'h43afe5f9},
  {32'hbeb66000, 32'h44a08d84, 32'hc51b59d1},
  {32'h4437cc03, 32'hc4cae697, 32'h44b8fe8d},
  {32'h436fd2ce, 32'h43e31559, 32'hc487a1a6},
  {32'hc4d45d29, 32'h43b5299a, 32'h43b81c6c},
  {32'hc3ef9d68, 32'hc434c56f, 32'hc5179223},
  {32'h44f20632, 32'h431da61a, 32'hc1a8d6d3},
  {32'h443df75d, 32'hc3fd462f, 32'hc5131507},
  {32'hc4272df1, 32'h44003ee8, 32'h44eaa717},
  {32'hc4259755, 32'hc274322f, 32'hc4cffba6},
  {32'hc4b27950, 32'hc386e90e, 32'h4476cae4},
  {32'h4285c148, 32'h438d6d6d, 32'hc485ed8e},
  {32'hc398b187, 32'h4434f9fd, 32'h4415b9b7},
  {32'h42dea0d8, 32'hc4ee0247, 32'hc35646c9},
  {32'hc3649789, 32'h44c721f3, 32'h43fb2a00},
  {32'h4481ed58, 32'hc30f991c, 32'hc20b52d2},
  {32'h42413938, 32'h445bfd53, 32'h44fb5cd6},
  {32'h43b7c1fe, 32'h41b453a9, 32'h41d93c70},
  {32'hc4f15363, 32'h413b9fd7, 32'hc2827ee2},
  {32'h42ab8be0, 32'hc489459d, 32'hc2f98ba8},
  {32'hc547b1f1, 32'h4463c58a, 32'hc362447f},
  {32'hc48a6eb5, 32'hc3640ad7, 32'h42bdea10},
  {32'hc491e45e, 32'h44581cca, 32'h445aff84},
  {32'h4483875f, 32'hc4d81751, 32'hc3d3a2c9},
  {32'hc4033566, 32'h4406d5c1, 32'h44064c26},
  {32'h44b9c163, 32'h42c4c812, 32'h42b4ec84},
  {32'hc424b000, 32'h43af1203, 32'h44237be9},
  {32'hc4b50d8c, 32'hc39afd81, 32'hc3bbde12},
  {32'h44dc9c40, 32'hc2e17fdd, 32'h42ed36ae},
  {32'hc488ac7a, 32'h437c7956, 32'hc3547439},
  {32'h45481bb4, 32'hc33c5f28, 32'h43ea4d48},
  {32'hc4bc96ec, 32'hc2ccbbee, 32'hc34970a7},
  {32'h42c80fb0, 32'hc493d9e6, 32'h42ed01b9},
  {32'hc3bad02c, 32'h44a56891, 32'h4124b56d},
  {32'h445e4ce6, 32'hc40ae3ab, 32'hc32dc147},
  {32'hc43485b8, 32'h44921e9b, 32'h425a9351},
  {32'h440e34b4, 32'hc500d84c, 32'hc1bbad8a},
  {32'hc5303792, 32'hc3ae87a6, 32'hc350b7c8},
  {32'h44e1c12d, 32'hc3c674b7, 32'hc3036cf8},
  {32'hc52ee7b7, 32'h43e35115, 32'h4344f2b4},
  {32'hc322b6e0, 32'hc21230ab, 32'hc3f70b62},
  {32'h424b3fb0, 32'h4316bcc2, 32'h44f9e81b},
  {32'h43998bb4, 32'hc4b2e826, 32'hc3a7f22c},
  {32'h440119f1, 32'h42adff42, 32'h440c13d9},
  {32'h449190f5, 32'h438dbf88, 32'h42cfd812},
  {32'hc0a670d0, 32'h44cbe8dd, 32'h4406bc95},
  {32'hc4d55a62, 32'h4323aded, 32'hc3cec0fb},
  {32'hc5459f0d, 32'h43f9c6ce, 32'h446b19d5},
  {32'h455e9162, 32'h43fb913a, 32'hc4175dd1},
  {32'hc2f2d15c, 32'h4506217a, 32'h423cd597},
  {32'hc35f2f8c, 32'hc4ec621d, 32'hc3899efd},
  {32'hc46903d4, 32'h44656349, 32'h4338f756},
  {32'h43096ef8, 32'hc4b6f3c6, 32'hc34f1029},
  {32'hc4c2348d, 32'h44811c78, 32'h44a1a9ad},
  {32'h45075270, 32'hc31b0580, 32'hc447ae22},
  {32'h44824fe0, 32'hc3e9c0ee, 32'hc2ed179c},
  {32'hc57f5752, 32'hc3bd0cca, 32'h43ddeb10},
  {32'h4523a05a, 32'h440b3f56, 32'h43bca74b},
  {32'hc42f891a, 32'hc39ef24b, 32'h44266e1a},
  {32'h44e577f0, 32'h4438a4ef, 32'h4434b62b},
  {32'h44997a59, 32'hc38828b5, 32'hc337cfd6},
  {32'h4412f806, 32'h4553df8c, 32'hc1dd0994},
  {32'hc439ac3a, 32'hc5348ec6, 32'h4305383a},
  {32'h447a05ad, 32'hc2a261ad, 32'h434975c3},
  {32'hc19e1f90, 32'h43a84376, 32'hc413f269},
  {32'h442cd9c2, 32'h4417d80e, 32'hc4f7e5a2},
  {32'hc3edc756, 32'h441f250c, 32'h44cd2bcc},
  {32'h412282b8, 32'h4497fc4b, 32'h43d868ea},
  {32'hc4d4bf4c, 32'hc3d52066, 32'h4354c2b4},
  {32'h443ac350, 32'h44033d85, 32'h43aa0064},
  {32'hc42b31d4, 32'hc2fbf96a, 32'hc5005371},
  {32'h43c8569c, 32'h440e2c08, 32'h45018815},
  {32'hc3b4667a, 32'hc49d1279, 32'hc2881858},
  {32'h45056cee, 32'h43e272ad, 32'h448456f3},
  {32'hc471259a, 32'h438e97af, 32'hc4964070},
  {32'hc4b14bb1, 32'h437095f3, 32'hc3089ded},
  {32'h42cc8a8d, 32'hc502a1f4, 32'hc429c51b},
  {32'h444044e7, 32'hc2a89f7f, 32'hc1973434},
  {32'h43763739, 32'hc504e178, 32'h413525a5},
  {32'hc35f63c0, 32'h45398e9d, 32'h435a258c},
  {32'h430aec9a, 32'hc4ca5419, 32'hc3503521},
  {32'h3f19ec80, 32'h44ead31b, 32'hc2e2a76f},
  {32'h42b9ce57, 32'hc3f928c4, 32'hc1c3d378},
  {32'hc420ecaa, 32'hc4a5e999, 32'h43ada833},
  {32'hc1718c3c, 32'h4548a6cd, 32'h41979eec},
  {32'h43746c6d, 32'hc30972e5, 32'hc1d3554e},
  {32'h4355895f, 32'h4525f93b, 32'h3e5d64c7},
  {32'hc4d60751, 32'hc472b253, 32'hc2229316},
  {32'h44ef96dc, 32'h43c71fd5, 32'hc35d5533},
  {32'hc572c449, 32'h440a61ad, 32'hc2253fef},
  {32'h43d61c88, 32'h44340399, 32'h44037dd3},
  {32'h4193151c, 32'hc44048e3, 32'h43ab3cf2},
  {32'h428e2536, 32'h4502e7e9, 32'h43bef303},
  {32'hc40ba7aa, 32'hc4effb39, 32'hc2c098f9},
  {32'h444b4382, 32'h43da05b0, 32'hc1a06048},
  {32'hc45b0e50, 32'hc4ac1076, 32'h433ec94c},
  {32'h439f8480, 32'h445f403c, 32'hc3bba284},
  {32'h441378ae, 32'hc3977338, 32'h444c7d3c},
  {32'h430368d0, 32'hc36d027a, 32'hc4e1b134},
  {32'hc489c190, 32'h43d7dfbd, 32'h4491bf6d},
  {32'hc4e141f2, 32'hc3169797, 32'hc38ed658},
  {32'hc4f0ad88, 32'hc438f4d7, 32'h43d2f1b5},
  {32'h430d800b, 32'h45193675, 32'hc3bb0078},
  {32'h43a1b51f, 32'hc239d9bc, 32'h43d8a7ee},
  {32'h44fb4844, 32'h433de889, 32'hc37ae64b},
  {32'h43daa975, 32'hc488123f, 32'h44831aee},
  {32'hc378335a, 32'h4404abe2, 32'hc3645860},
  {32'hc54cc724, 32'h415648cf, 32'hc4158b6e},
  {32'h45387148, 32'h436d5429, 32'hc3f172c6},
  {32'hc382c624, 32'hc507c269, 32'hc2d6cdee},
  {32'hc3ad92c5, 32'h448e398a, 32'hc2ca4aa5},
  {32'h439f30ca, 32'hc4c0262e, 32'h41a9a339},
  {32'h42ca48d5, 32'h455bf2ce, 32'hc247e458},
  {32'h439fea8c, 32'hc3a450cb, 32'h4338f1b6},
  {32'h444e3736, 32'h4390104a, 32'hc2313b81},
  {32'h45497c0f, 32'h42e365b7, 32'hc33e8e84},
  {32'hc5071799, 32'h4475c6c6, 32'h4434b4d7},
  {32'hc49406cc, 32'hc42e32d0, 32'h42e911bf},
  {32'hbf990480, 32'h44bcb8d4, 32'h4399108f},
  {32'h44db901e, 32'hc08c16b8, 32'h4273cb40},
  {32'h42e4e15c, 32'h445b592e, 32'hc35b0782},
  {32'h44daee10, 32'h432744c4, 32'h445eedd8},
  {32'hc40d11ce, 32'h44522fc6, 32'hc414417c},
  {32'h4433dee4, 32'hc3f6cca8, 32'h433bc9b9},
  {32'hc48a6d74, 32'h4336f3d1, 32'hc473cac8},
  {32'h4377c198, 32'hc3bef45c, 32'h4440ccbc},
  {32'h4425a44d, 32'h43dcded1, 32'h442e584b},
  {32'h44a02fac, 32'hc4274c13, 32'h44757916},
  {32'hc3e262ee, 32'h44470aed, 32'hc43b2256},
  {32'h44ab7480, 32'h43a23ac1, 32'h42c4439f},
  {32'h424137e8, 32'h456a9b02, 32'hc1ec1cd5},
  {32'h435c2816, 32'hc38f5afe, 32'h44917186},
  {32'hc467344a, 32'h43ae2864, 32'hc30a7b58},
  {32'h44842aae, 32'h444341c5, 32'h453f2ce2},
  {32'hc45e909a, 32'h43c91426, 32'hc4b23542},
  {32'h44ba093b, 32'hc3a9355b, 32'h43b6d8d5},
  {32'hc4a46a49, 32'hc421e978, 32'hc41eacf4},
  {32'hc3485af0, 32'hc4bd22b5, 32'h445e961a},
  {32'hc4bc5c20, 32'h441d9591, 32'hc39f87c5},
  {32'hc4348e94, 32'h42d66fdb, 32'hc3074304},
  {32'h43f089f5, 32'h433ac008, 32'h440449a8},
  {32'hc3c9bf3a, 32'hc3d5cb10, 32'hc4f1c18e},
  {32'hc23dfa65, 32'hc45793f7, 32'hc2113c39},
  {32'hc55676c7, 32'h436b12ae, 32'hc4038508},
  {32'h4412a60c, 32'hc3a4c2f8, 32'h450b050d},
  {32'h4464728f, 32'hc499bec4, 32'h44ced385},
  {32'hc4137d7a, 32'hc46b053a, 32'hc4b23407},
  {32'hc4c75193, 32'hc2fc44c0, 32'h43b154fe},
  {32'h3fbc4a20, 32'h42c980c3, 32'h4492f2cd},
  {32'hc4ef0e27, 32'h42eeea94, 32'hc3ecbd81},
  {32'h44fbaedb, 32'hc22503be, 32'hc0d89937},
  {32'h43c22c67, 32'h43efd5fb, 32'hc4ebde48},
  {32'hc3249ac2, 32'hc55e6c67, 32'hc3849d53},
  {32'hc406fad4, 32'h44d9830b, 32'h4199d1a4},
  {32'h44d3c0d8, 32'h428459ed, 32'h4465e461},
  {32'hc582ef9c, 32'h4395c23e, 32'hc32b9306},
  {32'h456b75dc, 32'hc34c5264, 32'hc40211f6},
  {32'hc51424db, 32'hc3060651, 32'hc3ac5488},
  {32'h44d53428, 32'hc4af12d3, 32'hc34ecf0c},
  {32'h43bfb828, 32'h44fad41f, 32'hc38ca09e},
  {32'h44ee26ce, 32'h4391d816, 32'h43e18be5},
  {32'hc49dac45, 32'h44dc68c4, 32'hc3811e7f},
  {32'h44f12dd8, 32'hc484461d, 32'h43b59628},
  {32'hc49fa6a1, 32'hc3ee6bd3, 32'hc38df178},
  {32'h43e8053d, 32'h44700b92, 32'hc4a17d0d},
  {32'hc38630e3, 32'hc4bebe47, 32'h4481e6e6},
  {32'hc5285952, 32'hc327d05a, 32'h440a96a1},
  {32'h43c66820, 32'h44d1b6b2, 32'hc40ecc45},
  {32'hc4630f3e, 32'hc448e559, 32'h42bd7544},
  {32'h44d763c2, 32'h435cf6dc, 32'hc465e60f},
  {32'hc44f23fd, 32'hc4e30ade, 32'h438265d5},
  {32'hc391ddf8, 32'hc266bfc9, 32'hc44387ac},
  {32'h44b50da3, 32'h420c1eef, 32'h43a2db1f},
  {32'hc45cf11f, 32'h4398f248, 32'h44853da4},
  {32'h439b69d0, 32'h444d2e67, 32'hc4bfb093},
  {32'hc3a8309e, 32'h428a6333, 32'hc48b10ca},
  {32'hc4c9c59c, 32'hc4095d51, 32'h434c91d8},
  {32'hc1789340, 32'h4374627c, 32'hc4e6400b},
  {32'hc4812a1c, 32'hc496fcde, 32'h43aea031},
  {32'hc2aa65ea, 32'h44b62ee6, 32'hc3ef56da},
  {32'h42e4ac70, 32'hc38b63e1, 32'h43b6c223},
  {32'h4446183a, 32'hc162368c, 32'hc30d38d6},
  {32'hc56bf94e, 32'hc415efc3, 32'hbfc23b80},
  {32'hc50a1d54, 32'h41a782fd, 32'h402853d0},
  {32'hc4b28f9c, 32'hc49410c1, 32'h43a9e18c},
  {32'h4484bd08, 32'h44c81121, 32'h44053845},
  {32'hc5099224, 32'hc338ab9f, 32'hc1a84abc},
  {32'hc3b978d6, 32'h452db2ee, 32'h43fc8357},
  {32'hc409e5ca, 32'hc4ef2dfc, 32'hc2e93842},
  {32'h44814f29, 32'hc1f0cf9a, 32'hc243277a},
  {32'h40e7cc40, 32'hc4ad0b5d, 32'h4498baae},
  {32'hc2db5590, 32'hc229f51f, 32'hc417c9c5},
  {32'h43f93924, 32'hc310d99c, 32'h44509033},
  {32'hc3c6ab0e, 32'hc43db0e6, 32'hc39b3be9},
  {32'h44559c12, 32'h41867ea4, 32'h43ac9ee6},
  {32'hc31e1222, 32'h4303d548, 32'hc4c8732a},
  {32'h449b5297, 32'h4286a1ea, 32'h44312c7d},
  {32'hc3689df0, 32'hc492b4b1, 32'hc4c4059c},
  {32'h44ef77f4, 32'h439016ad, 32'h43294635},
  {32'h43336591, 32'h4491075e, 32'hc403a728},
  {32'h442c3578, 32'h43ea13a8, 32'h44479e69},
  {32'hc334237a, 32'h443caa1c, 32'hc534d75f},
  {32'h448a82ee, 32'h433371d1, 32'h42c33ae1},
  {32'hc32b99f3, 32'hc4213fa6, 32'hc53d1de6},
  {32'h4468bfe5, 32'h44a34734, 32'h43ae06bc},
  {32'hc499f19a, 32'hc3c8d82e, 32'hc22fd9c3},
  {32'hc3847221, 32'h450dd163, 32'h44d94f41},
  {32'hc384f37c, 32'hc28f4865, 32'hc55541fe},
  {32'h443d0d14, 32'h43e9a304, 32'h42f4061f},
  {32'hc51b149f, 32'hc390f319, 32'hc325e67a},
  {32'h454f9f6f, 32'h444a88f0, 32'h43961a57},
  {32'h44bf40da, 32'hc3a22a76, 32'hc378d191},
  {32'h438f6724, 32'h446226aa, 32'h4300fba4},
  {32'hc3ff0e88, 32'hc587e0f6, 32'h420c9b24},
  {32'hc4c6e900, 32'h437b113d, 32'hc38abf54},
  {32'hc579a790, 32'h42b86cf1, 32'h42d94563},
  {32'h4571f630, 32'h4353d488, 32'h43d981d7},
  {32'h449eb3ac, 32'hc40a0dfa, 32'hc4069a42},
  {32'h43cbb79e, 32'hc38681d2, 32'h450ac671},
  {32'hc3614b00, 32'hc3848eab, 32'hc40c5e0b},
  {32'hc3c2432e, 32'h4511b75a, 32'h423913b1},
  {32'h44a3e67d, 32'hc4899a27, 32'hc2bf622d},
  {32'hc42486b2, 32'h447b3150, 32'h4431cd94},
  {32'h43a1f8c8, 32'hc3dbb3d7, 32'hc5425cf0},
  {32'h40392570, 32'h44df8fa4, 32'h450ebfe6},
  {32'hc48bed72, 32'hc3c4df88, 32'hc4833313},
  {32'hc3e4666c, 32'hc4a87904, 32'h44af07aa},
  {32'h44b97dc6, 32'hc35b75ba, 32'hc4069158},
  {32'h443b6c4e, 32'h442a1974, 32'h43a8034d},
  {32'hc2dcf112, 32'hc4cf7147, 32'hc3f46058},
  {32'h438af5e7, 32'h44cdfd94, 32'hc27dc5ba},
  {32'hc401ef5b, 32'h42a5a162, 32'hc43c4cc9},
  {32'hc39edb90, 32'h44a9c0ba, 32'h44cb6f85},
  {32'hc361c5a3, 32'hc4d0084d, 32'hc4624064},
  {32'h43f301e4, 32'hc30b13bf, 32'h43c701b1},
  {32'hc1a26e29, 32'hc546f787, 32'hc3fd7e86},
  {32'hc53d4c85, 32'h449cb4ca, 32'h43912a1c},
  {32'h43e245d0, 32'h408fe1dc, 32'hc3ad5e32},
  {32'hc503148b, 32'h44a1fd8d, 32'hc36f9402},
  {32'h44f51b12, 32'hc477378b, 32'h4390c23b},
  {32'hc40a2909, 32'h4416ac33, 32'h43a48554},
  {32'hc3f60332, 32'hc418ef01, 32'hc4025a36},
  {32'hc54eeb50, 32'h436acacd, 32'h44419a6d},
  {32'h45171641, 32'h4338a6e3, 32'hc3ab6d24},
  {32'h44fcdd16, 32'h434cfe59, 32'h42ade1a0},
  {32'hc5427f23, 32'h42c85365, 32'hc36ec1d9},
  {32'h453b70cc, 32'h43ce36a9, 32'h43ce2356},
  {32'h441a8c12, 32'h421e509d, 32'h43c05d12},
  {32'h440bcbaa, 32'hc520e1c7, 32'hc39368fa},
  {32'hc4ca0102, 32'h4459a6c5, 32'hc225c124},
  {32'h43a57d5d, 32'hc3dde1d4, 32'hc1c5ec97},
  {32'hc42c5a09, 32'h449cb533, 32'h436120e2},
  {32'h43fd8886, 32'hc4c754d9, 32'h43af1058},
  {32'hc4d9a9c1, 32'hc3097b70, 32'hc3b07116},
  {32'h4485c2ce, 32'hc3994534, 32'hc283550d},
  {32'h43607218, 32'h437f39ac, 32'hc48f14a9},
  {32'h431ee5ac, 32'h41b22966, 32'h43ee2121},
  {32'hc40941c2, 32'h44814e43, 32'hc38e92ef},
  {32'h4484a946, 32'hc4710ab4, 32'hc41f48a7},
  {32'hc4675854, 32'h42d2fbbe, 32'hc356c9ae},
  {32'hc40117fd, 32'hc4437afe, 32'hc2819ef7},
  {32'hc3acb812, 32'h43879f72, 32'h45470708},
  {32'h45684179, 32'h435546dd, 32'hc35f2cca},
  {32'hc57836f0, 32'h431c391f, 32'h4412fb08},
  {32'h44069942, 32'h441426e0, 32'hc4af399a},
  {32'h441bdc12, 32'hc295bf1f, 32'h43ab761d},
  {32'h44c1dfa9, 32'hc42bca60, 32'hc43055f9},
  {32'hc315679a, 32'h44a4e2ef, 32'h44f885e8},
  {32'h4446f034, 32'hc3280f4f, 32'hc4639a25},
  {32'hc50d966a, 32'h4462e527, 32'h42648638},
  {32'h436a5590, 32'hc4e4b490, 32'hc2d7983d},
  {32'h45041ded, 32'hc30deaa5, 32'hc33964d9},
  {32'hc41d914f, 32'h43ece90f, 32'h43807eef},
  {32'hc3e8f270, 32'h43d20c62, 32'h4373cb0f},
  {32'hc5367d98, 32'hc458fdd7, 32'hc43a3dbe},
  {32'h44210591, 32'h44dd4534, 32'h436a5f76},
  {32'hc439f346, 32'hc0a579e1, 32'h42b2b1c7},
  {32'h44f29af4, 32'h4447e4fe, 32'hc31c1daa},
  {32'hc46de5e9, 32'hc4d92f93, 32'h437ae94a},
  {32'hc47205b8, 32'h441c31f2, 32'h43d515d5},
  {32'hc4ca84e0, 32'hc1cc774f, 32'hc43ae15e},
  {32'h44764a37, 32'h443b577a, 32'h444f55e5},
  {32'h438bfe24, 32'hc2d673e9, 32'hc2dda55f},
  {32'h443b2a8e, 32'h44aafe9b, 32'h441118d3},
  {32'hc478d39e, 32'hc51b26fe, 32'hc379427a},
  {32'h4511ae4a, 32'h433ca4e2, 32'h42b24db6},
  {32'hc3ee0f48, 32'hc3cb2d40, 32'hc31bcc47},
  {32'h44083e1d, 32'h44d197aa, 32'h42622846},
  {32'h43aa784f, 32'hc4a6accd, 32'hc3b7a2b9},
  {32'h455a65ed, 32'h438a3339, 32'h4302ad6d},
  {32'hc42163a6, 32'hc30185bb, 32'hc4013138},
  {32'h44605078, 32'hc409ce4d, 32'hc358588f},
  {32'hc40230a6, 32'hc3949537, 32'hc4757aea},
  {32'h44f4417b, 32'h42a54a2c, 32'hc2eeb199},
  {32'hc205cf02, 32'hc4ee7761, 32'hc3afb549},
  {32'h43f29588, 32'h44aca9a9, 32'h4456de01},
  {32'hc3cb075b, 32'hc3657f55, 32'hc48dc3b1},
  {32'hc4630e8b, 32'hc36cd2c0, 32'h437172c1},
  {32'h443c7635, 32'h441ef9d5, 32'h4315d6e8},
  {32'hc452e528, 32'hc497bbcc, 32'h43830491},
  {32'h449dc444, 32'h4452f992, 32'h43ab065a},
  {32'h43655176, 32'hc419f7b6, 32'h4106bfd7},
  {32'h442fd94e, 32'h4436c4bc, 32'hc35ee2de},
  {32'hc3cc7a29, 32'hc5679d53, 32'hc3170a4f},
  {32'hc493e51c, 32'h4413cb8a, 32'hc2706610},
  {32'hc534c6bc, 32'hc3da526d, 32'hc311ea65},
  {32'h4352ff38, 32'h44968ada, 32'h44559530},
  {32'h44938647, 32'hc3ee69d2, 32'h4246ef3e},
  {32'h44515326, 32'h43acda8c, 32'hc3ffc1e7},
  {32'hc4983632, 32'hc3f2b896, 32'h42d1a557},
  {32'h4543738d, 32'h438865e8, 32'hc39e5a0a},
  {32'hc400ef49, 32'hc5506c3f, 32'h43c25771},
  {32'h429fa640, 32'h445ddbd7, 32'hc4ecc54a},
  {32'h4468758e, 32'hc40fb605, 32'hc39b811e},
  {32'h44ff394b, 32'h41249b7c, 32'h42ea8d1d},
  {32'hc4393bf4, 32'h436d557d, 32'h445b633e},
  {32'h4360c2f8, 32'h3f1d6e20, 32'hc48d6b1a},
  {32'hc48c1dbb, 32'h434541d7, 32'hc20d40fc},
  {32'h43647e95, 32'h45257760, 32'hc380a8c1},
  {32'hc48845b8, 32'hc4812d42, 32'hc437d995},
  {32'hc3a01309, 32'h445b171e, 32'hc49dfbd6},
  {32'hc4c63176, 32'h4246b602, 32'h4480fef1},
  {32'h44e98e86, 32'h43d7e276, 32'hc3abcdfd},
  {32'hc4c34bd9, 32'h4429a622, 32'h44d6eafa},
  {32'h4410cbbf, 32'hc3497032, 32'hc4f9e74e},
  {32'hc29f28c4, 32'hc544dd0b, 32'hc3e80b1a},
  {32'hc51d2d31, 32'h448a902c, 32'h4201f461},
  {32'h44bf1437, 32'h3feb0d20, 32'h4322df41},
  {32'h41b3799a, 32'h44bb3908, 32'h43551de5},
  {32'h449cfd58, 32'hc4afa0f0, 32'h4415b384},
  {32'hc44d1c18, 32'h4407ae38, 32'h42505955},
  {32'hc37228a0, 32'h43501fe7, 32'hc462c994},
  {32'hc5918111, 32'h443e75ac, 32'hc422b43e},
  {32'h451380ae, 32'h43518b10, 32'h43e19012},
  {32'hc3874120, 32'h4428c39f, 32'hc4cd6c65},
  {32'hc3c67f4f, 32'hc3fbac25, 32'hc4823616},
  {32'h4307159a, 32'h4497f902, 32'h40df4bae},
  {32'h4504d87e, 32'h43d4e789, 32'h446ce698},
  {32'hc3fd3bcb, 32'h446471d9, 32'hc3e74ac3},
  {32'h44d50546, 32'hc2638902, 32'hc1cd276f},
  {32'hc48af079, 32'h42ae40eb, 32'hc449f1be},
  {32'h427d2258, 32'hc2d91378, 32'h44bb89df},
  {32'hc521082c, 32'hc3a2a45f, 32'hc1329968},
  {32'h44476294, 32'hc4a49c8b, 32'h42b1ac3f},
  {32'hc4d4c638, 32'h448534e9, 32'hc46a52f1},
  {32'hc47f8916, 32'hc3dbc9fc, 32'h441bfea3},
  {32'hc3d8e433, 32'h456cbdc3, 32'h43462b66},
  {32'h4530cf9f, 32'hc35eb4e0, 32'h435bec96},
  {32'hc49dd09f, 32'h4187a74e, 32'h436acc7e},
  {32'h4425e5a4, 32'h43de2a84, 32'h45125c08},
  {32'hc43aff05, 32'h43ebdac3, 32'hc48c6cb7},
  {32'hc2bad84c, 32'h4396fb1a, 32'h449b5f23},
  {32'hc50cd06d, 32'hc39cd31e, 32'hc3c817d1},
  {32'hc2261bf0, 32'hc4f4f2b1, 32'h44981b29},
  {32'hc32a0535, 32'h444c4773, 32'hc3b88d2a},
  {32'h44bb6621, 32'h4334b051, 32'hc3683405},
  {32'h442230c8, 32'h43516f02, 32'h445c03c9},
  {32'hc4c0395d, 32'hc3e723d4, 32'hc48efd0e},
  {32'hc2b69341, 32'h43846761, 32'h44eedc03},
  {32'hc44d05a2, 32'h448c6f2c, 32'hc36dcd2c},
  {32'h43794ae6, 32'hc5168a70, 32'hc3aad7a0},
  {32'h41d12ea0, 32'hc3cdef63, 32'h44f80175},
  {32'hc39e9bb4, 32'h4463d41d, 32'hc49de21a},
  {32'h43ab4a8d, 32'hc20e537c, 32'h441ff270},
  {32'hc3b72897, 32'hc36f1003, 32'h44282f50},
  {32'hc473831e, 32'h44957f82, 32'h43065c61},
  {32'h43e3749b, 32'hc40bb921, 32'h4487e467},
  {32'h43795a00, 32'h4491f28a, 32'h4375923d},
  {32'h43d16068, 32'hc4c88bbf, 32'h43e3af4a},
  {32'h425de69b, 32'h44dcb13a, 32'hc3960c5c},
  {32'h4539ab34, 32'hc41bf02e, 32'hc3085be0},
  {32'hc5519074, 32'h43416baf, 32'h437aded5},
  {32'h451308dc, 32'hc346f241, 32'h43c073b0},
  {32'h44fcb8be, 32'h43917e2f, 32'hc1d359a3},
  {32'h452031bf, 32'hc38283ce, 32'h44123b46},
  {32'hc40cc8c6, 32'h4467d35f, 32'h435ea770},
  {32'h442b27f5, 32'hc3866972, 32'hc3c529e5},
  {32'hc4cc2502, 32'h4465b03e, 32'h43abc4a3},
  {32'h44a0319d, 32'hc482f6ac, 32'hc2348ba2},
  {32'h42d92246, 32'hc39e542e, 32'h43d3d0e4},
  {32'hc3d1bcd0, 32'hc4884e70, 32'hc54f9ab9},
  {32'h4292477b, 32'hc49bf9dc, 32'h4492f6ea},
  {32'hc4fcab62, 32'hc39a1bc7, 32'h42fa825e},
  {32'h44765314, 32'h43b70132, 32'hc458e32f},
  {32'hc50cf3d2, 32'h41e8e411, 32'hc3a851bc},
  {32'h439678fe, 32'h43ecf0ca, 32'hc49480ee},
  {32'hc44ade44, 32'hc485f930, 32'h43f4695d},
  {32'h43034dd4, 32'hc2a6a17e, 32'hc4f5948f},
  {32'hc49792f0, 32'hc1b11ad6, 32'h43b7e65e},
  {32'hc4e54f0a, 32'hc351c1c9, 32'h43e6abd0},
  {32'h4439b76a, 32'hc4634f64, 32'hc424c4a1},
  {32'h43f66466, 32'h438716a6, 32'hc480017c},
  {32'hc481515d, 32'h42d51e22, 32'h4467a680},
  {32'h44a68e2f, 32'h43459a15, 32'hc353e752},
  {32'hc44022d5, 32'hc391f93f, 32'h41ee7797},
  {32'hc2d10b50, 32'h450919a9, 32'hc39424d8},
  {32'hc4fb1953, 32'hc3df2521, 32'hc33c0488},
  {32'h45797dc4, 32'hc3ec7b24, 32'h439dbfce},
  {32'hc593cd02, 32'hc291ce3a, 32'h434c16d9},
  {32'h452ca8a0, 32'h42ff614c, 32'hc31be210},
  {32'hc50b9ecd, 32'hc45b0e42, 32'h41d97cbd},
  {32'h42613bcb, 32'h45272d83, 32'h4318f7f0},
  {32'hc54de800, 32'h43962b37, 32'hc358a228},
  {32'h43a2eeec, 32'h45042f85, 32'hc3fe5573},
  {32'hc528b288, 32'hc2c3466f, 32'h43f81572},
  {32'h447be1ef, 32'h42a4fe72, 32'hc40c11fb},
  {32'hc2c6e084, 32'h44a2434c, 32'h43c42f44},
  {32'hc39c2d84, 32'hc51baa17, 32'hc4210aa6},
  {32'h443c6537, 32'hc41033e3, 32'h447aac7d},
  {32'h4350c9fe, 32'hc4b454dc, 32'hbff547e0},
  {32'h43d10102, 32'h439146c7, 32'h452b348b},
  {32'h432500c0, 32'hc504385a, 32'hc43032ba},
  {32'hc3267e4e, 32'h4301faf5, 32'hc39968b5},
  {32'hc44d1046, 32'hc478fc5a, 32'hc4cb2a61},
  {32'h418ec610, 32'h44a3dc3f, 32'h451dfa9f},
  {32'h4337733d, 32'hc4dd1c18, 32'hc2f8bd4e},
  {32'h43838d36, 32'h43c8e636, 32'h4399b4c0},
  {32'hc489dc29, 32'h4404d3e2, 32'hc42e713f},
  {32'hc4ba65a5, 32'h4359c41f, 32'hc2194f08},
  {32'hc52b5fc6, 32'h43ae6fc5, 32'hc21afcc1},
  {32'h445e1bf1, 32'h446bbd2e, 32'h439b6d49},
  {32'h44a85368, 32'h4337fa71, 32'hc32f9232},
  {32'h451ca3ae, 32'h436a4469, 32'h43afe653},
  {32'hc2a9d9ae, 32'hc3c08737, 32'hc534eb1c},
  {32'h44a43e44, 32'h44397eb1, 32'h433dd7c9},
  {32'hc4c6a3cb, 32'hc4411008, 32'hc41f8646},
  {32'h44ac60b2, 32'h44b44d62, 32'h44116912},
  {32'h440f0dae, 32'hc4225f39, 32'hc3b3b211},
  {32'h4451b95f, 32'h44be6343, 32'h44206cbf},
  {32'hc49ba64c, 32'hc4b06e4c, 32'h42f8070b},
  {32'hc4961e33, 32'h4232bdce, 32'h43b0b70e},
  {32'hc4015660, 32'hc35bc237, 32'hc369e31b},
  {32'h452a2da6, 32'h41edf960, 32'h42e7f876},
  {32'h44c20408, 32'hc3cf6619, 32'hc43f0d7a},
  {32'h437db6d8, 32'hc3ea9e21, 32'h448b35fb},
  {32'hc3139d86, 32'h43ceb82c, 32'hc4c374ce},
  {32'hc4d3aef9, 32'h448f9a6e, 32'h440bde2a},
  {32'h45050784, 32'hc2adaa57, 32'h43ddd97a},
  {32'hc41615e3, 32'h423870fc, 32'h44eff626},
  {32'h43147c78, 32'hc468bfd4, 32'hc4da3790},
  {32'h444c3bb2, 32'hc33fc4e2, 32'h440eb679},
  {32'h437b5dac, 32'hc4aed32b, 32'hc361ed28},
  {32'hc3a474c6, 32'h44918d35, 32'h440c3034},
  {32'hc3e91340, 32'hc4dfd3f3, 32'hc46e9176},
  {32'hc4eb50e0, 32'h43a76090, 32'h41151164},
  {32'h43b41221, 32'hc32ee6a1, 32'hc4d28d77},
  {32'hc37e67aa, 32'h44e2fa3d, 32'hc260d118},
  {32'h43e5f13c, 32'hc1573968, 32'hc4e5f061},
  {32'hc4da5bb5, 32'h43b064a6, 32'h4434cbc1},
  {32'h44896225, 32'h42316b18, 32'hc415ce78},
  {32'hc3ae6dde, 32'h4113054a, 32'h4448618f},
  {32'h430c4be0, 32'hc5730f86, 32'hc3e8b54e},
  {32'hc4593cb8, 32'h446860b4, 32'h4404ecb3},
  {32'h4338c281, 32'hc4d3db0c, 32'hc2947770},
  {32'hc5076d2a, 32'h443dae35, 32'hc3899452},
  {32'hc2644680, 32'hc4c4e0e3, 32'h439529bd},
  {32'hc4106f1d, 32'h4469ed7b, 32'hc36db4ed},
  {32'hc30c4de0, 32'hc41baea5, 32'hc3baae3b},
  {32'hc54cf82a, 32'hc402907c, 32'hc30c6b0c},
  {32'hc38f7c9c, 32'hc3f68d1d, 32'hc3b23864},
  {32'h445f0b41, 32'hc400038e, 32'h4497df88},
  {32'hc508edd4, 32'hc1b1e183, 32'hc3633135},
  {32'h430b645f, 32'h43a4bbf3, 32'h449f9f97},
  {32'hc3e17870, 32'h44bc816b, 32'hc33e3aa0},
  {32'h452891d4, 32'hc39419bc, 32'h432bd063},
  {32'hc3b58822, 32'h440812b4, 32'hc444540f},
  {32'h4486f246, 32'h43837602, 32'hc3dca3fc},
  {32'hc511f428, 32'h443a3a40, 32'h427187c5},
  {32'h44eb1232, 32'hc3d852fa, 32'h44241db7},
  {32'h43d7d0cb, 32'h4310dcd1, 32'hc3c584fc},
  {32'h43b21bc6, 32'hc35fc73e, 32'hc1ee3175},
  {32'hc399439a, 32'h437b74c9, 32'h439d768a},
  {32'h44490a48, 32'hc3073526, 32'hc47ebdde},
  {32'hc3bcdd5c, 32'h444bab0f, 32'h448a89c7},
  {32'h43ab2873, 32'hc50bf805, 32'hc3292deb},
  {32'hc4c44d3e, 32'h42fe6a03, 32'h43fe8a33},
  {32'h4448e782, 32'hc4d8a7d7, 32'hc1a5ace0},
  {32'hc412883f, 32'hc21c2fcc, 32'h449b2599},
  {32'h43a5241c, 32'hc3cb8e19, 32'hc3c4d9ce},
  {32'hc536fd8d, 32'hc43120dc, 32'hc25a4350},
  {32'h454374fd, 32'h432f193f, 32'hc45aab30},
  {32'h443b5345, 32'h434b5ba6, 32'h436cd7ae},
  {32'h43cafc1f, 32'hc3cb8897, 32'hc52d0204},
  {32'hc3adff88, 32'hc2939ea6, 32'h45302a31},
  {32'h439f8d47, 32'hc46958b4, 32'hc3af323b},
  {32'hc40b1ff0, 32'h442f61a1, 32'h445c7689},
  {32'h4505064e, 32'hc48ed4f3, 32'hc3c61f49},
  {32'h4381d538, 32'hc3c28f8e, 32'hc55f8fc0},
  {32'hc4823208, 32'h43969332, 32'h44a41619},
  {32'hc4affde9, 32'h4266590b, 32'h4393ec79},
  {32'hc4af26be, 32'hc3f24d13, 32'h43382e53},
  {32'h4562cf6b, 32'hc2b2b9dc, 32'hc33799cf},
  {32'h4332069c, 32'hc4c28006, 32'hc416987a},
  {32'h44633f58, 32'h45142132, 32'h441589aa},
  {32'hc3b41078, 32'hc45d9197, 32'h43d0ec28},
  {32'hc4897c30, 32'h441b4490, 32'h43231fff},
  {32'hc464bfab, 32'hc40b79dc, 32'hc3f53f5d},
  {32'h450c8588, 32'h4413c908, 32'h4310750b},
  {32'h44632b23, 32'h43b2eefa, 32'hc3b5482c},
  {32'h44621026, 32'h448e44c4, 32'h43d952cd},
  {32'hc3297dc6, 32'h43377cc3, 32'hc3f82da4},
  {32'h44541394, 32'h42be8dc4, 32'h441d9ad0},
  {32'hc31ffb42, 32'hc4ca7c0c, 32'h428855b4},
  {32'h44040488, 32'h44c4fb72, 32'h44a19c0c},
  {32'hc301281b, 32'hc5000980, 32'hc3728ec2},
  {32'h4523515f, 32'hc3d3f14c, 32'h440a9259},
  {32'hc5007854, 32'h442a93f3, 32'hc465ee19},
  {32'hc3950e13, 32'h4337db1d, 32'hc285627e},
  {32'hc41949cc, 32'hc37f0054, 32'hc49dd494},
  {32'h438f74f4, 32'h44f13ccf, 32'h424e5ec7},
  {32'hc4107dff, 32'hc437a1d5, 32'hc42d98d5},
  {32'h4315aa20, 32'h449acf2d, 32'h447b32d4},
  {32'hc4e7c652, 32'hc3f4773a, 32'hc482d0cc},
  {32'h4499ff9a, 32'hc3387a47, 32'hc3e943f8},
  {32'h4449a196, 32'h449164c7, 32'hc3b75684},
  {32'hc448704e, 32'hc4975ce5, 32'hc3043fd5},
  {32'h449223b5, 32'h436466f3, 32'h441e3d19},
  {32'hc537960b, 32'h430d6a43, 32'hc3794b8b},
  {32'h4448b7ca, 32'hc1f999ca, 32'h44188341},
  {32'hc50a1746, 32'hc2e3ef3c, 32'h4294f346},
  {32'hc4e437d5, 32'h4339fe5b, 32'h4335cc99},
  {32'hc50dbdfb, 32'h4339da5c, 32'hc39de683},
  {32'h445cfd20, 32'hc2b54350, 32'h4345d28a},
  {32'h439584b5, 32'hc4a77231, 32'h430481af},
  {32'h45030d4d, 32'hc2c6d002, 32'hc35e33dd},
  {32'hc2af277a, 32'hc505f77f, 32'hc295b697},
  {32'h430a45d0, 32'h448f3770, 32'h438e5ca5},
  {32'hc3a49fef, 32'hc5242548, 32'hc119aaba},
  {32'h443268c9, 32'h44a4da87, 32'hc3248999},
  {32'hc47374f5, 32'hc38af19b, 32'h43a9dd45},
  {32'h4373974d, 32'hc1036182, 32'hc4ab9519},
  {32'hc4850189, 32'h43407104, 32'h43f916c1},
  {32'h45131e8f, 32'hc3c7c170, 32'hc484e7aa},
  {32'hc57ce759, 32'hc3c48ee8, 32'h42ce0992},
  {32'h4427f0fd, 32'h4533b3cc, 32'hc239adb0},
  {32'h44d568ad, 32'hc254aa39, 32'h4386599e},
  {32'hc3a96831, 32'h4523320c, 32'hc3826a6d},
  {32'hc401c1b0, 32'hc446d257, 32'h445ba5e3},
  {32'h45753bdc, 32'h4404646d, 32'h4369a193},
  {32'hc46cd332, 32'h43cdc518, 32'h446baa8c},
  {32'h43a1835c, 32'hc3f00c64, 32'hc526f12e},
  {32'hc286c620, 32'hc5553760, 32'h43b1b60b},
  {32'hc446f2fc, 32'h43e77f57, 32'h449ef5bd},
  {32'h432cce3b, 32'hc45a583f, 32'h42cbd6d9},
  {32'hc49ee433, 32'h44bc28c0, 32'hc41175e0},
  {32'h44cd4a1b, 32'hc4526972, 32'hc3872849},
  {32'h4219a4c8, 32'h4513c58d, 32'h42ecc59d},
  {32'h44660368, 32'hc47615e6, 32'hc39ba46b},
  {32'hc50e8c34, 32'h43f2e437, 32'h433120e6},
  {32'hc221e4ad, 32'hc3bedbd2, 32'hc2cf4602},
  {32'h433e1c59, 32'h41986738, 32'h444b8d45},
  {32'h440a4029, 32'hc4bb7c7a, 32'hc346773e},
  {32'hc47b71c8, 32'h422bcfb2, 32'hc2e884e1},
  {32'h44ace4c8, 32'h43bc2cd7, 32'h44b9c06b},
  {32'hc0d170aa, 32'h452314a1, 32'h4361a79a},
  {32'hc388cc28, 32'h430caec4, 32'h44d6d4c6},
  {32'h434085c1, 32'h43e3824a, 32'hc32389a4},
  {32'h44c4f6a2, 32'hc476354a, 32'hc3ba3dbc},
  {32'hc42ee3e2, 32'h44402f9e, 32'h437c9d54},
  {32'h4412b6ca, 32'hc4e218a5, 32'hc14c763e},
  {32'hc4b92b53, 32'hc317294c, 32'h4247e7da},
  {32'h45033b12, 32'hc2c552d6, 32'h428e3eb8},
  {32'hc5243d2e, 32'h43af9198, 32'hc35656ea},
  {32'h45045104, 32'h43aa1894, 32'h43ac0eb7},
  {32'hc446c472, 32'hc36bbfda, 32'hc48019fa},
  {32'h42f5df60, 32'hc360b54e, 32'h4469a873},
  {32'hc4f8fcfa, 32'hc3bea287, 32'hc50dc79d},
  {32'h4524051e, 32'h42a99dc2, 32'hc3543c26},
  {32'h43650a90, 32'hc4403a59, 32'hc55f701f},
  {32'h42a9848a, 32'hc4245314, 32'h453ac85b},
  {32'hc37b35d7, 32'h446859cb, 32'hc3f4f0d3},
  {32'h43e54163, 32'h43a1c350, 32'hc481598f},
  {32'h44f89c0e, 32'hc4246b94, 32'hc2894d81},
  {32'hc206bfc0, 32'h4355c916, 32'hc4adbbd5},
  {32'hc343db4e, 32'hc3a95069, 32'h4486dac4},
  {32'hc4e417ed, 32'h449879ed, 32'h413c230d},
  {32'h428449ea, 32'hc4c8bab0, 32'hc388f227},
  {32'hc3e92fac, 32'hc302737f, 32'h45598b65},
  {32'h42dae9e0, 32'hc4b47e19, 32'hc489a42d},
  {32'hc3a858ef, 32'hc305333e, 32'h449bcaea},
  {32'h429e203e, 32'hc3be9627, 32'h448ceb17},
  {32'hc4b90f64, 32'h43734be8, 32'hc40c6cfd},
  {32'h43f60fa3, 32'hc47dc161, 32'hc3f826ce},
  {32'h430ca4b4, 32'h4203316f, 32'hc3f15587},
  {32'hc3b69d46, 32'hc53b4065, 32'hc31ffe04},
  {32'hc41c3957, 32'h43a81e79, 32'hc1571e22},
  {32'h4331d2dc, 32'h42a18e20, 32'h43ca854a},
  {32'hc561ce36, 32'h43e62af7, 32'hc3ce6071},
  {32'h45033ac7, 32'h43b36ed6, 32'hc357b509},
  {32'h442cd203, 32'h44dc7569, 32'h4370f636},
  {32'hc3bd286b, 32'hc588eaed, 32'hc33b403d},
  {32'hc51f66e1, 32'h43c3a699, 32'hc3112673},
  {32'h443b6704, 32'hc4287bd4, 32'h42147ef9},
  {32'hc3260870, 32'h44cee667, 32'hc4036bd3},
  {32'h445dc5e8, 32'hc409570b, 32'h44039ee4},
  {32'hc2f51b98, 32'hc3201b93, 32'h431814a9},
  {32'h41209f18, 32'h44a6bfab, 32'hc4d05bb4},
  {32'hc30eb450, 32'h42951e31, 32'h44ae3c56},
  {32'hc54111c2, 32'h41927bd3, 32'h431f774b},
  {32'h4554de34, 32'hc3921bed, 32'h440291b1},
  {32'hc3f2517c, 32'hc426ee27, 32'h42efcca0},
  {32'hc3d2d87d, 32'h4538492d, 32'h3ee4edc0},
  {32'hc463a7cc, 32'hc502f68e, 32'h4319847d},
  {32'hc48bf924, 32'h4289d0b3, 32'hc43ed730},
  {32'h441f8a1b, 32'h4492dd1b, 32'hc43f5ea5},
  {32'hc3b9bb5f, 32'hc31ec90b, 32'h44c09b62},
  {32'hc31ee804, 32'h43cdb269, 32'hc4d255d7},
  {32'h43842000, 32'h43c5063b, 32'hc4bbeeca},
  {32'hc51d8f7a, 32'hc38bb9ab, 32'h43bcf47c},
  {32'hc409d91c, 32'h44890006, 32'h4206bdb3},
  {32'hc3a296f2, 32'h4344a2c2, 32'h44d318d4},
  {32'h439c81d2, 32'hc3b1715c, 32'hc49e2870},
  {32'hc2fddd7c, 32'hc4b8c429, 32'h43325c11},
  {32'h450d290f, 32'hc39223d9, 32'hc3e3f408},
  {32'hc593b6a7, 32'hc17c5c1c, 32'h42b1bce3},
  {32'h4460cd16, 32'h43491b6f, 32'hc353d522},
  {32'hc2e65538, 32'hc55083db, 32'hc3292910},
  {32'h44a6746f, 32'h441fc461, 32'hc30793ae},
  {32'h4460aeb0, 32'hc41d9c4b, 32'h43045faa},
  {32'h44f3a012, 32'h44862bc8, 32'h4193140b},
  {32'hc47f05ae, 32'hc51b182d, 32'h43961d8f},
  {32'hc21f4188, 32'h44d863a0, 32'hc1ad7b90},
  {32'h442adff2, 32'h43452e75, 32'hc36eeeac},
  {32'hc3bdcea5, 32'h43390c6f, 32'hc486de71},
  {32'h43776922, 32'h44502b61, 32'h44a0c172},
  {32'h44dbb59a, 32'h41c18019, 32'h42eab888},
  {32'hc36b70c8, 32'h441ddb5c, 32'hc41babb0},
  {32'hc4816efc, 32'hc46ea627, 32'hc39b65b3},
  {32'hc3c7e96f, 32'h44820257, 32'h43ffcede},
  {32'hc54572e6, 32'hc2fa06c3, 32'h42d29507},
  {32'h4317420a, 32'h42b98382, 32'h4439bee8},
  {32'h42f19832, 32'h44521518, 32'hc4b60379},
  {32'h430eab96, 32'h44cec594, 32'h44150ac4},
  {32'h42615720, 32'hc448a733, 32'hc490e378},
  {32'h453af8ef, 32'hc31808fc, 32'h438d6512},
  {32'hc472b452, 32'hc42062f6, 32'hc404f37e},
  {32'h441b7b7c, 32'h440949fc, 32'h44dcdadf},
  {32'hc4239772, 32'hc2c3873f, 32'hc45eaa8c},
  {32'h437cee4e, 32'h43828db4, 32'h45605eb2},
  {32'h41864a66, 32'hc40a9e5c, 32'hc4a01750},
  {32'h4446afbc, 32'h43136983, 32'h4433ea3c},
  {32'hc4b55798, 32'hc4aa61d9, 32'hc3b63811},
  {32'h44f68b64, 32'h4472fc1e, 32'h42a42cb8},
  {32'hc4e1eeae, 32'h43e5eae6, 32'h42be45eb},
  {32'h44ed1cc0, 32'h43bf82cd, 32'hc3ab7be5},
  {32'hc45ad926, 32'hc529b05b, 32'hc2e33d74},
  {32'hc4882f70, 32'hc20b87da, 32'h44113cf2},
  {32'hc50e1b4a, 32'hc22c3c0e, 32'hc487b998},
  {32'h456e2502, 32'hc357e310, 32'hc3b23332},
  {32'h440d5dc5, 32'hc3fe123c, 32'hc3e40717},
  {32'hc428ca3c, 32'h44f10075, 32'h4301191b},
  {32'hc3c039a2, 32'hc411ec47, 32'hc3bf7313},
  {32'hc3567c01, 32'hc0282f10, 32'h451c3009},
  {32'hc3bf383c, 32'hc3ef7388, 32'hc5267320},
  {32'h43f64554, 32'h440bd04f, 32'h44a18d4a},
  {32'h449f35f2, 32'hc4263ad9, 32'hc45448b1},
  {32'hc381761a, 32'h446003f7, 32'h45087eb9},
  {32'h440027b3, 32'h429bb793, 32'hc3cf13a9},
  {32'hc3da4e4d, 32'h43453e4d, 32'h44919772},
  {32'hc4e1b140, 32'h43ac8d81, 32'hc48fdd1f},
  {32'hc3828c1c, 32'hc4293d8a, 32'h447907ce},
  {32'hc329b93d, 32'hc3928a8d, 32'hc516e7e8},
  {32'hc411fb54, 32'h43951219, 32'h442ee8e0},
  {32'h44e9b7ca, 32'h43ee64b1, 32'hc37d74a2},
  {32'hc42c63aa, 32'h430a21f2, 32'h43800e4b},
  {32'h45350c8e, 32'hc3986ed0, 32'hc1ce3210},
  {32'h447b9ba6, 32'hc2f6f3d9, 32'h43bede67},
  {32'h44276590, 32'hc4f13e21, 32'h4387c221},
  {32'hc55236b7, 32'h4275e888, 32'h437dcf83},
  {32'hc442298d, 32'hc435cf90, 32'h41d71a97},
  {32'hc51b6bf9, 32'h443bd43c, 32'h40c93c31},
  {32'h45764d4a, 32'h428134f4, 32'h43cb7338},
  {32'h4450736c, 32'h42a34587, 32'h431290db},
  {32'h44a1b96d, 32'h4449af57, 32'h429a4bd6},
  {32'hc534bd8b, 32'hc3f003d9, 32'hc3997d18},
  {32'h42f7fca3, 32'hc3f5cee7, 32'hc33f395c},
  {32'hc4768605, 32'hc38489b2, 32'hc2cd3a2f},
  {32'hc42b6332, 32'h41bf1dc0, 32'hc52e5b29},
  {32'h4525c56f, 32'h43098332, 32'h444ab32d},
  {32'hc380953e, 32'h44896923, 32'hc311a74c},
  {32'h448e6503, 32'hc49c03a3, 32'hc3422469},
  {32'hc413714b, 32'h44a7feb3, 32'h438f2948},
  {32'hc32198c8, 32'hc438cd6d, 32'hc3861594},
  {32'hc53215de, 32'h42e53d80, 32'h426e2b4b},
  {32'h440d4bfb, 32'hc517670c, 32'h42419877},
  {32'hc4284e53, 32'hc3d22167, 32'h430a9d2d},
  {32'h4420a9a4, 32'h438a62c5, 32'h44a98ed9},
  {32'hc4f876a8, 32'h43b399ef, 32'h43ece4b0},
  {32'hc4ee19d9, 32'h42b32b55, 32'h42cd42b2},
  {32'h41967b00, 32'h4419f233, 32'h44db8125},
  {32'h43cee55e, 32'hc42e8634, 32'hc4d6304f},
  {32'hc4c5673d, 32'h41825382, 32'h439de9d2},
  {32'h45354d80, 32'h43d2e6ae, 32'hc2f78584},
  {32'hc531aabb, 32'hc3efd319, 32'hc2a3bcd7},
  {32'h445eeb51, 32'hc3a210ff, 32'hc3d96111},
  {32'hc554da45, 32'h43230f24, 32'h43abb2fe},
  {32'h4484864b, 32'hc40a2ace, 32'hc48de57e},
  {32'hc43176e0, 32'hc18c3799, 32'h44b3f8c4},
  {32'h44bf8320, 32'hc3b681fc, 32'hc45efad6},
  {32'h42aac9fb, 32'hc2ac53b4, 32'h4521f471},
  {32'h442451f6, 32'hc3b84348, 32'hc3de6d8b},
  {32'hc3163e87, 32'h44251b2f, 32'h45043703},
  {32'h448e62e0, 32'hc439ad5b, 32'hc4088de2},
  {32'h44b87ef3, 32'h43b0ff00, 32'hc4898acf},
  {32'hc4045628, 32'h4299dc22, 32'h4493d598},
  {32'hc3fc42d5, 32'h445d7e97, 32'hc485ecf9},
  {32'hc4176014, 32'hc47e50c6, 32'hc3d57c53},
  {32'h4505ae6c, 32'h43188b2d, 32'hc38abc40},
  {32'hc489a408, 32'h42b101f6, 32'h431170a1},
  {32'h43a29e98, 32'h456cbf7e, 32'hc3c43ab7},
  {32'hc4a1b228, 32'hc4a69f60, 32'h43be47b8},
  {32'hc2619d94, 32'h450ceaf9, 32'h42735810},
  {32'hc2c023a8, 32'h438281b1, 32'hc49ac8b0},
  {32'hc2eabd96, 32'hc3e774aa, 32'h443661f5},
  {32'h425c56c0, 32'h4310b631, 32'h443fcc30},
  {32'h438b3885, 32'h44030378, 32'h45233552},
  {32'hc475fd70, 32'hc3eea5c0, 32'hc432e9da},
  {32'hc4cde820, 32'h43dc07d7, 32'h4410f3d5},
  {32'hc3d79109, 32'hc50e2b2b, 32'h42c80bbb},
  {32'h453c98d9, 32'h4373a7d3, 32'h42b77041},
  {32'h42e6776c, 32'hc49adc05, 32'h42c534fc},
  {32'h45480dbb, 32'hc38cc3a5, 32'h4229b9f0},
  {32'hc54a6629, 32'hc3a5dbdb, 32'hc3bd42f4},
  {32'hc470e88a, 32'hc2253cef, 32'h42c6e484},
  {32'hc4e5d764, 32'hc3ac708b, 32'hc4671cc4},
  {32'h43b9f312, 32'h4458aafc, 32'h44199ddf},
  {32'hc5225632, 32'h4172d6ee, 32'hc3232bd9},
  {32'h4508fd3d, 32'h445a52af, 32'h440527db},
  {32'hc43545b0, 32'hc4b25db3, 32'hc30c95ae},
  {32'hc356d8fc, 32'hc2902dcc, 32'h448cd7be},
  {32'h4494d386, 32'hc3cafb30, 32'hc3842812},
  {32'hc53c4569, 32'hc31ba962, 32'h43cd22ea},
  {32'h452f23fd, 32'h4407e859, 32'h43011aaf},
  {32'hc4d47f21, 32'hc34a5fa5, 32'h43dc1b57},
  {32'hc2892720, 32'h44bf1180, 32'h43ed6295},
  {32'h43870106, 32'hc5493fec, 32'h418b5802},
  {32'h43cff4e8, 32'hc31c6878, 32'hc4492202},
  {32'hc507e7d5, 32'hc417d943, 32'h4255a493},
  {32'h451dbeba, 32'h441036f9, 32'h440116dd},
  {32'hc5024676, 32'h42f89c9d, 32'hc4191a0c},
  {32'h42b73ba4, 32'h4295da7f, 32'h43400704},
  {32'hc4a39ce2, 32'hc2fa5dc3, 32'h44805d57},
  {32'hc2c9a1ba, 32'h44dc0745, 32'h42852f3c},
  {32'hc52ba6da, 32'hc3f0b186, 32'h4328d7b6},
  {32'h43d9ed78, 32'hc12950ac, 32'hc4610665},
  {32'h42fbdc07, 32'hc12094a6, 32'h44c146c8},
  {32'h4486d6ed, 32'h4380b92d, 32'hc4a246d3},
  {32'hc4054c12, 32'h42944344, 32'h44133a64},
  {32'hc4197903, 32'h44610e9a, 32'hc31621ca},
  {32'hc4adbbd5, 32'hc4d16179, 32'h45230662},
  {32'h42dae6bd, 32'h4457d2c8, 32'hc51e0f9c},
  {32'hc41a7e7d, 32'h410de288, 32'h43f877be},
  {32'h4481e447, 32'h43a13991, 32'hc401758c},
  {32'h432697c8, 32'hc43e9f68, 32'h44a81ad3},
  {32'h43b43c5b, 32'hc386514a, 32'hc4fe908e},
  {32'hc55360f0, 32'hc37ac7ba, 32'h438eafae},
  {32'h4464d8e8, 32'h4265a30d, 32'hc4f0c170},
  {32'h45220aee, 32'hc429396c, 32'h43b25bcf},
  {32'hc3fc5d70, 32'h445aad9c, 32'h4072e186},
  {32'h44b9f38c, 32'h43abd488, 32'h43fd85e8},
  {32'hc522f88d, 32'h44491b4d, 32'h44063f83},
  {32'h454ade58, 32'hc370e681, 32'hc33763c5},
  {32'hc4fd9542, 32'hc39f9e4b, 32'hc2d02448},
  {32'h442fb2c8, 32'hc3f81819, 32'hc47b9adf},
  {32'hc5870a81, 32'h437859cc, 32'h41f168fa},
  {32'h43fdaf80, 32'hc30e1695, 32'h4360623b},
  {32'h43cd3ba5, 32'h4462e2ff, 32'hc2b5ad2d},
  {32'h42b8fb3c, 32'hc4fdaabc, 32'h4270f8a0},
  {32'hc50706bd, 32'h42b2f9da, 32'h43781cc8},
  {32'h44400fdf, 32'h421e59df, 32'h4361552e},
  {32'hc36ebf22, 32'h431775bb, 32'hc49b55bb},
  {32'h44d48194, 32'h42c12d74, 32'h43070811},
  {32'hc4403c65, 32'h43347c70, 32'hc48b647f},
  {32'h45595d8c, 32'h4364d855, 32'hc3edfe07},
  {32'h447fb79a, 32'hc3846185, 32'hc3c2f098},
  {32'hc2d7486e, 32'hc4c7aca1, 32'h448ef4b5},
  {32'hc47f9094, 32'h43faa5bf, 32'hc49b732c},
  {32'hc411dd22, 32'hc3350551, 32'h43926314},
  {32'hc386acb0, 32'hc2bf5d4e, 32'hc50b42d1},
  {32'h44b33fbe, 32'hc48ca968, 32'hc3badaef},
  {32'h4400a484, 32'h4416b406, 32'hc43d5adc},
  {32'h421b0981, 32'h441c3399, 32'h44e43079},
  {32'hc56073da, 32'h424066b5, 32'hc384c150},
  {32'h4381c024, 32'hc360a7e6, 32'hc3ac6074},
  {32'hc4538870, 32'h446ab9d5, 32'hc35981f2},
  {32'h44c76e2c, 32'hc3369734, 32'h44192b32},
  {32'hc45494bc, 32'h442b247b, 32'h444cfc74},
  {32'h4405ad52, 32'h4352dc9d, 32'hc34245b6},
  {32'h43d759a2, 32'hc3c55bfc, 32'h44fc4ce1},
  {32'hc3a89ddf, 32'hc3be1044, 32'hc535b633},
  {32'hc2ae172e, 32'hc4e75e8b, 32'h42cbdf76},
  {32'hc4fc14fe, 32'hc27c94a8, 32'hc3ac0150},
  {32'h414dc54a, 32'hc3e9af31, 32'h45100555},
  {32'hc40808d8, 32'h44938a7e, 32'h45131a4d},
  {32'hc327e276, 32'h4387f42c, 32'hc538b114},
  {32'h42239332, 32'hc4bf6637, 32'h44588c3a},
  {32'hc3481472, 32'hc47e5d80, 32'h440d0fd0},
  {32'hc551fc11, 32'hc34a69a2, 32'h43912675},
  {32'h44823281, 32'hc2028731, 32'h44b0d270},
  {32'h4255bea4, 32'h441e8be9, 32'hc3c31583},
  {32'h410bbc80, 32'hc549d810, 32'hc3a3104b},
  {32'h44244df2, 32'h452eff81, 32'hc2c5cfbf},
  {32'h443ca982, 32'h439439cc, 32'hc201e633},
  {32'hc506d19c, 32'h43ce5662, 32'h430d6ed3},
  {32'h458050ed, 32'h43464d14, 32'hc3c7553b},
  {32'hc40d6701, 32'h4461fd96, 32'hc3db18f7},
  {32'h45198070, 32'hc44a489e, 32'h4353795a},
  {32'hc4396054, 32'h40a1d0a4, 32'hc38f194b},
  {32'hc2da26b3, 32'hc4344bde, 32'hc3b38a53},
  {32'hc4b41e12, 32'h44b67e9f, 32'hc425e274},
  {32'h44a27342, 32'hc4d7d7d8, 32'h438efe7d},
  {32'h448eae8b, 32'hc358032a, 32'h437141b3},
  {32'h4392e14a, 32'h428f4dee, 32'hc4ab816f},
  {32'hc422fd74, 32'hc4dd924d, 32'h44b10ba4},
  {32'hc4aa7a9f, 32'h431877ad, 32'h448360b6},
  {32'h447dc520, 32'h440f98ba, 32'hc2ac2488},
  {32'hc347625f, 32'h4381d482, 32'h4468d63c},
  {32'hc3917c76, 32'h4426977e, 32'hc542a2fb},
  {32'hc452b910, 32'hc4a68244, 32'h443acbd5},
  {32'hc30b018e, 32'h44d51e26, 32'hc238b740},
  {32'h42517808, 32'hc35ffafc, 32'hc43ae43a},
  {32'hc4e00b3e, 32'hc449d9e8, 32'h44f1bfa0},
  {32'hc3073f10, 32'h447d725d, 32'hc50f612a},
  {32'h44208bef, 32'h44552c44, 32'h43c2845f},
  {32'hc3488cb4, 32'h430d9608, 32'h445bddbf},
  {32'hc43c7ad8, 32'h43dd9f2d, 32'hc3ef71f3},
  {32'hc4c32679, 32'h418595ff, 32'h44145d2a},
  {32'h44db35f6, 32'hc2924e31, 32'h4310aab9},
  {32'hc39d7138, 32'hc4ca778f, 32'hc2a8c28e},
  {32'h4548bff1, 32'h42c8422f, 32'h428f0436},
  {32'hc59d1048, 32'h4379f71a, 32'h421ae006},
  {32'h438c1730, 32'h43a10737, 32'hc38b079c},
  {32'hc4e09d44, 32'hc42ab8ac, 32'h4359a474},
  {32'h44e64fba, 32'hc22e7ab7, 32'hc29055e5},
  {32'hc3cbd03e, 32'hc4e2374c, 32'hc2332ffb},
  {32'h425016f3, 32'h4562990f, 32'hc2d3f2d9},
  {32'hc42f129a, 32'hc3e11f5a, 32'h4377fd43},
  {32'h44b113b4, 32'hc3125227, 32'hc2200c77},
  {32'hc4b603a0, 32'hc39ef998, 32'h43133101},
  {32'hc37bc228, 32'hc4936708, 32'hc42f0e2e},
  {32'hc2c39d4a, 32'hc4b61765, 32'h44d71650},
  {32'hc3af9f73, 32'h41de9238, 32'hc4889c83},
  {32'h43f33b86, 32'h4496513d, 32'h44a7f0d0},
  {32'hc43031d8, 32'hc4dc8406, 32'hc3084118},
  {32'hc2b2f3c4, 32'h44257b01, 32'h43dede18},
  {32'hc5168cc9, 32'hc3c170c1, 32'hc4313082},
  {32'h4519f5fd, 32'hc2fa4395, 32'h439277f5},
  {32'hc40a74d8, 32'hc3beb630, 32'h42b000fc},
  {32'hc3d27672, 32'hc49fcf8b, 32'h450f82f5},
  {32'h43db8ccb, 32'h43976c14, 32'hc43a7db6},
  {32'h4462db4b, 32'h439a0757, 32'h43886e79},
  {32'hc312427f, 32'hc3f07666, 32'hc52dffff},
  {32'h4478b671, 32'h44e1d8ec, 32'hc21879e2},
  {32'hc33b3b64, 32'hc499bea8, 32'h42ca0520},
  {32'h43ae6618, 32'h442a70e4, 32'h44b90752},
  {32'h4433a114, 32'hc304f348, 32'hc544fb47},
  {32'h4491f45f, 32'h4442c6e4, 32'hc3ab654e},
  {32'hc3da204c, 32'hc55b5024, 32'hc3587f98},
  {32'h44be2cfb, 32'h44a0cfcd, 32'hc38c85c8},
  {32'hc4ad1b49, 32'hc25351b0, 32'hc270f678},
  {32'h4455eabf, 32'h44a6c20e, 32'hc30cab98},
  {32'hc5081d45, 32'hc418dd38, 32'h4321070c},
  {32'h45624e91, 32'h430df687, 32'h441126f9},
  {32'hc32264d0, 32'hc3977d25, 32'h440534ff},
  {32'h446d42ca, 32'h43da4db6, 32'h428ee43e},
  {32'h44ae26d3, 32'hc38accd8, 32'hc3d5f601},
  {32'h42a0d824, 32'hc4b273dd, 32'h43cb74dd},
  {32'h435e1eae, 32'hc415dca4, 32'h43b693ca},
  {32'hc4983237, 32'h44bb3f31, 32'h42ff6366},
  {32'hc3b99aea, 32'hc5172653, 32'h41d60238},
  {32'h4227b036, 32'h433a04d3, 32'h442e8cf6},
  {32'h44bee462, 32'hc49e97a4, 32'hc481915d},
  {32'hc4a6df46, 32'h43b8e88f, 32'h44e358ce},
  {32'hc2a51532, 32'hc4b718f0, 32'hc382765b},
  {32'hc2097f90, 32'hc4019a16, 32'h44a660b2},
  {32'hc3083c4f, 32'h4528c6d8, 32'hc4ed0df1},
  {32'h442e6078, 32'hc45336a3, 32'h4401034e},
  {32'hc3790855, 32'hc46c7ea1, 32'hc4579f4a},
  {32'hc4f8c034, 32'h43cbc517, 32'h439cdbd5},
  {32'h440924e3, 32'hc4343ce1, 32'hc3df05a7},
  {32'h43ac25a8, 32'h449882c4, 32'h44b35f6e},
  {32'h4522fa59, 32'h43c26546, 32'h42148aa6},
  {32'hc4a02f16, 32'h4469af70, 32'h43871702},
  {32'hc31fca88, 32'hc510e211, 32'hc41348e0},
  {32'h43bacc8c, 32'h458332d4, 32'h439b9a34},
  {32'hc36c560c, 32'hc48a50dc, 32'h423572b8},
  {32'hc516594b, 32'h43e205e0, 32'h4415c5e4},
  {32'h44eb6436, 32'hc429f856, 32'h43186efd},
  {32'hc4a055ec, 32'h440f8568, 32'h4397de9b},
  {32'h444c0394, 32'hc36e2cc5, 32'h4322b169},
  {32'hc54a6e92, 32'h40822400, 32'hc15a09e2},
  {32'hc4ce85e7, 32'hc4132887, 32'hc40e7333},
  {32'h43c1c166, 32'hc2d85b82, 32'h431615fc},
  {32'hc57a0013, 32'h4253ed9b, 32'h435040fd},
  {32'h4511f5a6, 32'h4319b0eb, 32'h43c8d9af},
  {32'hc4cac0b0, 32'h4382b605, 32'hc37eec9c},
  {32'h42a1aabc, 32'hc4f9b70b, 32'hc3b17994},
  {32'hc4bb54e2, 32'h447ad04f, 32'h43f573de},
  {32'hc47c124a, 32'hc434a38a, 32'hc3ca863d},
  {32'hc47538ab, 32'h450ac7fb, 32'hc3039c76},
  {32'h44c0eaa3, 32'hc4d51b3b, 32'h43858351},
  {32'h44fea692, 32'hc308df83, 32'hc2227846},
  {32'h452b7e74, 32'h42843a3b, 32'h42072cef},
  {32'hc4f0d93c, 32'h44630a8a, 32'hc38517c9},
  {32'hc49185ca, 32'hc296a90c, 32'hc0881130},
  {32'hc3734a04, 32'h44cf48de, 32'h44219d6a},
  {32'h44628641, 32'hc48a80bd, 32'hc3eaaa5e},
  {32'hc2514694, 32'h44b7c994, 32'hc33e9056},
  {32'h41b1e6c0, 32'hc3809f2b, 32'h4335cbf7},
  {32'hc50d4bbc, 32'h4211db25, 32'h44573533},
  {32'h45457c5b, 32'h418abcb9, 32'h43c7a7a6},
  {32'hc4498d45, 32'hc3c5e20d, 32'h442eb3f0},
  {32'h451329a9, 32'hc3230a04, 32'hc45208ee},
  {32'h44566979, 32'hc0bf1fd7, 32'h43b225be},
  {32'h44d057a8, 32'hc44a3d55, 32'hc4406e06},
  {32'hc44faef8, 32'h44ad7dfb, 32'h43800986},
  {32'hc308cdfa, 32'hc31c8341, 32'hc473afa1},
  {32'h4281d870, 32'h441c56f8, 32'h44ec9cda},
  {32'h43bef4c4, 32'hc4e3d108, 32'hc4491d17},
  {32'h44943422, 32'hc2f3485c, 32'hc32ebea7},
  {32'hc4a8189a, 32'h4410abf7, 32'h437b2418},
  {32'h44f58d53, 32'hc1ff9b1d, 32'h43b688f3},
  {32'hc485b21e, 32'hc49e4183, 32'hc32289b3},
  {32'h4305f8e0, 32'h44048c1c, 32'hc305b599},
  {32'h448dc7e2, 32'hc30a0c0a, 32'hc3e29e40},
  {32'h4486c404, 32'h44ca2ab1, 32'h433643ac},
  {32'hc47359cc, 32'hc48cfd20, 32'h43fbad90},
  {32'h443d4e27, 32'h447ffe14, 32'hc2495339},
  {32'hc5121f22, 32'h43bbb73e, 32'hc3cdb833},
  {32'h4418e612, 32'h42757c4c, 32'hc3bfc35f},
  {32'h44826e99, 32'h401b3f2d, 32'h44151967},
  {32'h43c12650, 32'h453e1637, 32'h43d2564f},
  {32'hc3e9f1be, 32'hc4394868, 32'hc49c56cd},
  {32'hc4008486, 32'h43341323, 32'h44f5c90a},
  {32'hc5396415, 32'hc366cf55, 32'h41fe92ae},
  {32'h440f1a43, 32'h44a61347, 32'h44a457ed},
  {32'hc3872ada, 32'hc4fb0672, 32'hc20916fc},
  {32'h434c69b0, 32'h437e8986, 32'h44a77912},
  {32'hc434af0c, 32'h42b91dd9, 32'hc33fda76},
  {32'hc4734e6e, 32'h431067cc, 32'h4350a31c},
  {32'hc4a320dd, 32'hc1812228, 32'hc4bd929c},
  {32'h444d0b3d, 32'h44b209cf, 32'h43416092},
  {32'hc517e7b1, 32'hc382c03b, 32'hc3368d92},
  {32'h43f0685c, 32'h44fed1af, 32'h43c36312},
  {32'hc489c9b5, 32'hc423b2e5, 32'hc4909c72},
  {32'hc462f0d4, 32'hc32571c0, 32'h43b59445},
  {32'h43bb567b, 32'h45172037, 32'hc3ca53ed},
  {32'hc4973890, 32'hc48b79fb, 32'h42a78414},
  {32'h43b9b4a0, 32'h44961334, 32'h442c82a1},
  {32'h41eca210, 32'hc48e94b1, 32'h41ed3064},
  {32'h44821533, 32'h44815e80, 32'hc33ca8c8},
  {32'hc3d59932, 32'hc5129c44, 32'hc2318d4e},
  {32'h451389f8, 32'hc28fa074, 32'hc3c87fae},
  {32'hc50c418b, 32'h4307cc50, 32'hc02507fe},
  {32'h44c556ba, 32'hc42b754e, 32'hc2a92dd0},
  {32'hc4882ac5, 32'hc3f34c24, 32'h44090593},
  {32'h44bbdaba, 32'h44418c48, 32'hc3e20feb},
  {32'hc50dbb0c, 32'hc3a3888d, 32'h429abe15},
  {32'hc4225e33, 32'h4479bd74, 32'hc2f400fc},
  {32'hc5095e2a, 32'h43ae8dd8, 32'hc3a0babf},
  {32'h43d7700e, 32'h453159db, 32'hc2e54ed0},
  {32'h43ed7344, 32'hc09e3a8a, 32'h43d76da1},
  {32'h44921d9c, 32'h441341ea, 32'hc1e6fe98},
  {32'hc40fb0e4, 32'h43be8e8f, 32'h4503a379},
  {32'hc3ede15b, 32'h44ad4edd, 32'hc2b9cbf2},
  {32'hc4e16396, 32'hc49601ba, 32'h4383d1d3},
  {32'hc1588c00, 32'h450aa87e, 32'hc42f191e},
  {32'hc507663f, 32'h43ad5094, 32'hc3267c28},
  {32'h45069902, 32'h437ad0f4, 32'hc41fbfd2},
  {32'hc54c16e9, 32'hc3cef6fc, 32'h4378588c},
  {32'h4386044c, 32'hc339a032, 32'hc4c4f0ca},
  {32'hc47c6e86, 32'h42b6997b, 32'h44aced19},
  {32'h4550d2e8, 32'h40f1b8a2, 32'hc43b3490},
  {32'h437a7090, 32'hc5132c4f, 32'hc14f9cca},
  {32'hc3c9d4d4, 32'h450d6ec4, 32'h42229131},
  {32'h453ae5d5, 32'h42b93253, 32'h437d8bdf},
  {32'hc4fb253d, 32'h44264331, 32'hc2f116d2},
  {32'h4495b7a0, 32'hc4361c1c, 32'hc34df253},
  {32'h4417aa2c, 32'h432ad0d3, 32'hc20b4313},
  {32'h4509e898, 32'hc45a629a, 32'hc41f5bce},
  {32'hc5058ad8, 32'h435debe1, 32'h422bc614},
  {32'hc4e9720f, 32'hc18faea8, 32'h42e9145c},
  {32'hc4a856c6, 32'h439936e6, 32'hc3db6dfa},
  {32'h442b0a1f, 32'h445d5758, 32'hc47493b6},
  {32'hc49186ed, 32'h4327bbf2, 32'hc0d9827e},
  {32'h43d148a4, 32'hc3a58227, 32'h44ea1cec},
  {32'hc3092bb0, 32'h43aab4fa, 32'hc4e83d18},
  {32'hc39886a2, 32'hc4eaf811, 32'hc399f436},
  {32'hc28a195c, 32'h4271d4d7, 32'hc4a8817e},
  {32'h44e7f165, 32'h440aeb84, 32'h4380f96a},
  {32'h43f9ddfe, 32'h4388b4b6, 32'hc49fccd4},
  {32'h42c41100, 32'hc45a7000, 32'h442ae48f},
  {32'hc4cdeeef, 32'h44693328, 32'hc4fe7776},
  {32'hc4abe914, 32'hc1f4f37e, 32'h43451774},
  {32'hc478235c, 32'h44a69407, 32'hc3fc6c91},
  {32'h43be6822, 32'hc3cb1c5c, 32'h4510b091},
  {32'hc2a14cda, 32'hc12dda09, 32'hc2d81454},
  {32'h4414ad3b, 32'h42f5eef7, 32'h4490152e},
  {32'hc4c0ef15, 32'hc422bd22, 32'hc513d086},
  {32'hc46c19e6, 32'hc4214ef5, 32'hc3652aba},
  {32'h42478c98, 32'hc4a4dbce, 32'hc4e4be01},
  {32'h438e3d36, 32'h447def82, 32'h44b1bbab},
  {32'h4259f1cc, 32'h445dabfc, 32'hc4872197},
  {32'hc4ac4c3c, 32'h43626835, 32'h43371b12},
  {32'h4512ac37, 32'hc3b37d07, 32'h42f56391},
  {32'h43cee40b, 32'h45154712, 32'hc3b75bf7},
  {32'h4256c2bd, 32'h438a7ab3, 32'h4396885b},
  {32'hc4c0244c, 32'h442507f2, 32'hc3a15aaf},
  {32'h449fd2ec, 32'hc464f648, 32'h447d2df9},
  {32'h43eaf1c4, 32'hc4c5d855, 32'h450fe567},
  {32'hc51804be, 32'h4454e768, 32'hc431f572},
  {32'h446fd906, 32'h420cbe52, 32'h42998d4d},
  {32'h42c94f08, 32'hc4134efd, 32'h440e0942},
  {32'hc388e667, 32'h451ae2a8, 32'hc3cb8cdd},
  {32'h4378637e, 32'hc4cb73d8, 32'h426cda47},
  {32'hc3e49e30, 32'hc188ee65, 32'hc43e9c34},
  {32'h448d4a80, 32'hc386ff81, 32'h44a15e77},
  {32'h42494b22, 32'hc31cfa6a, 32'hc521d82a},
  {32'h4510807f, 32'h42831435, 32'h4446dd86},
  {32'hc4bdd0a4, 32'hc3a8653b, 32'h43b63a1b},
  {32'h457344b9, 32'h42dcd868, 32'h440fbad1},
  {32'hc3bfe324, 32'h44c94cfb, 32'hc266a21e},
  {32'h44cc2ef9, 32'hc4bc31d2, 32'h437e3685},
  {32'hc4db7500, 32'h44197966, 32'h42f32b8b},
  {32'h44db9fa1, 32'h4438827c, 32'h438cf7b1},
  {32'hc32531d8, 32'h44aa1d61, 32'h43d06aab},
  {32'h44aa9f1e, 32'hc4db7e06, 32'hc394fb47},
  {32'h44bef9a6, 32'hc3b0d9b9, 32'h43b045f4},
  {32'hc373ffca, 32'h44acf00c, 32'hc4da8b4b},
  {32'hc3a58300, 32'hc4c7c0fb, 32'h44c2bef4},
  {32'hc4a1b9ae, 32'hc392a590, 32'h44abcabb},
  {32'hc154e510, 32'hc3ed7bd7, 32'hc4f1e465},
  {32'hc4e89f9c, 32'hc37df0ea, 32'h43848450},
  {32'h44c0d4a6, 32'h4382ac40, 32'hc377a505},
  {32'hc24b8d60, 32'hc4bcfc17, 32'h44555f4f},
  {32'h44fbd34c, 32'hc273b00c, 32'hc4563050},
  {32'hc2df61e0, 32'hc49cd28c, 32'h426eb653},
  {32'h43ef2855, 32'hc3d99d04, 32'h4526a862},
  {32'h432008b1, 32'hc4f28951, 32'hc4b6a9fa},
  {32'h44a002eb, 32'h445a7fe3, 32'hc404e7e2},
  {32'hc40e9e4e, 32'hc3999a1d, 32'h444f5dde},
  {32'h4361df26, 32'h44a61d48, 32'hc30b4286},
  {32'hc45df7fe, 32'hc4197460, 32'h449d6aaa},
  {32'h442bb142, 32'h450b5438, 32'h40e62c60},
  {32'hc1c403f1, 32'hc38746e4, 32'h43e5cf13},
  {32'hc3b4c935, 32'hc3ea50e0, 32'hc3d23db9},
  {32'hc527b183, 32'hc1e8be57, 32'hc3baae8e},
  {32'hc348b24e, 32'h425a5fa1, 32'hc34fd3a7},
  {32'hc45693c0, 32'hc515802d, 32'h43c88cce},
  {32'h43a3a5c8, 32'h44eace4e, 32'h417c84c4},
  {32'h4335c88a, 32'hc4ddbb5a, 32'h430b631d},
  {32'h454d5aae, 32'h43f14e9e, 32'h439d0544},
  {32'hc5246af5, 32'hc483efa6, 32'h439ee628},
  {32'h44e690fa, 32'hc36be2aa, 32'hc32fec62},
  {32'hc3b212d1, 32'hc42f5e5c, 32'hc338398c},
  {32'hc37ad32f, 32'hc3741664, 32'hc426501f},
  {32'h443c7c8e, 32'h4452dac0, 32'h44911b5a},
  {32'h442b0906, 32'hc035e253, 32'hc3d08efe},
  {32'h447b154b, 32'h43cc6724, 32'h4498c47d},
  {32'hc2cfbdc0, 32'hc53eb9fc, 32'hc2b53910},
  {32'h424c0e61, 32'h42fab6a8, 32'h44cd0773},
  {32'hc5753f3a, 32'h42d7ad59, 32'h431b35a9},
  {32'h45308938, 32'h43ce388b, 32'hc313fc0a},
  {32'h43e22786, 32'h44eee8c5, 32'hc41000dc},
  {32'h447ae42d, 32'h437c4939, 32'h434e923a},
  {32'hc2956858, 32'hc4e96c4e, 32'hc4074f10},
  {32'h44136f39, 32'hc220e29c, 32'h432caa58},
  {32'hc3344801, 32'hc461836f, 32'h43088220},
  {32'h44c14e8d, 32'h43df9a9b, 32'h421a9a71},
  {32'h432fc954, 32'hc3933054, 32'hc51a9817},
  {32'h44612c2e, 32'h440c9529, 32'h44ba2267},
  {32'hc51f8b49, 32'hc3eba5eb, 32'hc2f06f69},
  {32'hc33ce2b0, 32'h43b41008, 32'h4290fa9e},
  {32'hc4802138, 32'hc51fe54e, 32'h408589f5},
  {32'h443f9a1e, 32'h44cc63fe, 32'h43adc69a},
  {32'h412238c0, 32'h42b7bc2a, 32'h440a5315},
  {32'h447cc4a0, 32'h448371fe, 32'hc3d3ef69},
  {32'hc42f79f8, 32'hc53341c5, 32'hc347df54},
  {32'h419d5230, 32'hc323dad7, 32'h41bde621},
  {32'hc530995f, 32'hc34c8fd6, 32'hc42fd582},
  {32'h43c75230, 32'hc345c15e, 32'hc39ac606},
  {32'hc308a2ca, 32'hc48a7d61, 32'hc46ed811},
  {32'hc434c480, 32'h446c2467, 32'h43d792a2},
  {32'hc451ff9f, 32'hc4abb880, 32'hc2948bd2},
  {32'hc38949aa, 32'hbd1a3800, 32'h45315986},
  {32'h449c9810, 32'hc27ee22e, 32'hc3ecab7c},
  {32'h41267d24, 32'h43742b0d, 32'h44a437d5},
  {32'h41984f68, 32'hc3a9602a, 32'hc5401e51},
  {32'hc43522fd, 32'h440c6ea1, 32'h45194c67},
  {32'h444c8a7e, 32'h4408014f, 32'hc4fcdc29},
  {32'h438f1e0c, 32'h44769b9c, 32'h443c343f},
  {32'h4417f129, 32'hc385be1b, 32'hc48cbabd},
  {32'hc1ed9100, 32'hc46621e6, 32'h44365015},
  {32'h443cf833, 32'hc334d045, 32'hc4cdff1d},
  {32'hc45c7aec, 32'hc4070901, 32'h45129a4e},
  {32'hc3923cad, 32'hc4c53c3a, 32'hc2919e58},
  {32'hc3e80c98, 32'h448e3b4d, 32'h44a01cfc},
  {32'h4456f21c, 32'hc3957288, 32'hc35d6f5d},
  {32'h44195ec2, 32'h443c8833, 32'h445910e2},
  {32'h448d3b10, 32'hc4d18997, 32'h425b5258},
  {32'hc3d17ce0, 32'h45043346, 32'h4396d78d},
  {32'h439c8773, 32'hc4120a86, 32'hc39928ed},
  {32'hc52ae2ef, 32'h43b7b8b9, 32'hc2cd0261},
  {32'h44195ed4, 32'hc490de1e, 32'hc335a13a},
  {32'h43438890, 32'h4484c939, 32'h4185132a},
  {32'h44e68b7a, 32'hc3b5e495, 32'hc402e20e},
  {32'hc54bee22, 32'h442d2773, 32'hc38695c4},
  {32'h454537b0, 32'hc308b086, 32'h4062cdb8},
  {32'h44f2838c, 32'hc3ec1642, 32'hc3c3237f},
  {32'hc53a71b2, 32'h4347c292, 32'hc382b2ad},
  {32'h44df8166, 32'hc2a3bd8b, 32'h4487c6a1},
  {32'h44d2767c, 32'h42c45efc, 32'h43851036},
  {32'h43af1761, 32'hc5012f59, 32'hc2c4783a},
  {32'hc420979e, 32'h44e4dd8c, 32'h43941c4c},
  {32'h449349e9, 32'h42f9517a, 32'h4294ddce},
  {32'hc34d97b2, 32'h45734b44, 32'hc330d1e6},
  {32'h43bce610, 32'hc54be5cc, 32'h43359ee7},
  {32'h43baf25c, 32'h41975564, 32'h42f70ac6},
  {32'h43c8da42, 32'hc3cd0b12, 32'hc41e1f88},
  {32'hc34d2a67, 32'h446242a0, 32'hc4ff2f77},
  {32'hc3fe1a05, 32'hc482db4b, 32'h4325ccf1},
  {32'hc5016cb8, 32'hc3235444, 32'hc14a9019},
  {32'hc41d0ef0, 32'hc4c913d7, 32'hc48b4611},
  {32'hc4d95f79, 32'h3e9dfabc, 32'h4398a762},
  {32'hc2bba480, 32'hc475aed9, 32'hc4598a86},
  {32'hc47dd344, 32'h44374972, 32'hc35c209c},
  {32'h44f1bf2c, 32'h439a47ff, 32'hc43927ec},
  {32'hc4aa2844, 32'h43e0ebfc, 32'h437810b4},
  {32'h4549904e, 32'hc386b178, 32'hc43e9abe},
  {32'hc4c095da, 32'h428f2ff2, 32'hc23e4117},
  {32'hc2081f76, 32'hc4117704, 32'hc5165a30},
  {32'hc48e196a, 32'h43532759, 32'h44fabdde},
  {32'h4485bfbe, 32'hc350c818, 32'hc46401a5},
  {32'hc481fcfb, 32'h439e09ac, 32'h4406f2c8},
  {32'hc2e9551c, 32'hc50c4dff, 32'hc483a739},
  {32'h44bca103, 32'hc3c969e8, 32'hc3b25248},
  {32'hc3d4e372, 32'hc386d2c4, 32'h4513f24a},
  {32'h442d38b1, 32'h43474c48, 32'h4422e292},
  {32'hc52a6c7d, 32'h438a3a43, 32'h44016adf},
  {32'h43c52804, 32'h450d662d, 32'h43874b3f},
  {32'hc3e2ce0f, 32'h412aa231, 32'hc359e4ae},
  {32'h4429b470, 32'h43d751bb, 32'hc3ea4071},
  {32'hc392a014, 32'hc526a2d7, 32'hc3013a53},
  {32'hc34141dc, 32'h4362b3d2, 32'h4387dcbd},
  {32'h429528ff, 32'hc3431e05, 32'hc344af17},
  {32'h434430f8, 32'h4338cab9, 32'hc396ea12},
  {32'h44d54063, 32'hc3e29d13, 32'h4408ddd6},
  {32'h43ad2c1d, 32'h44f908d0, 32'h4380f3e2},
  {32'hc3dcf56e, 32'hc35eed50, 32'h42d8dd6b},
  {32'h43e15d9e, 32'h440af564, 32'h438cba10},
  {32'hc3c3403a, 32'hc3c9b71d, 32'hc522fbcb},
  {32'h4402c9da, 32'h4393c5ac, 32'h4529ed4f},
  {32'hc474a71a, 32'hc3d07dcb, 32'hc3618efa},
  {32'h44501dd8, 32'hc45c1495, 32'h43c3d450},
  {32'hc48e0854, 32'h44360386, 32'hc33a47c6},
  {32'h4505ad61, 32'hc2cebe8a, 32'hc41c2f9a},
  {32'hc363df30, 32'hc4e439e2, 32'hc402fda3},
  {32'hc281e510, 32'h4458ddcf, 32'h44893ef8},
  {32'hc49287cf, 32'hc427920e, 32'hc3b4f6ef},
  {32'h44cb6a05, 32'h42eeffc6, 32'h44907adb},
  {32'hc4ac379d, 32'hc476b58d, 32'hc386495d},
  {32'h453dfe8a, 32'hc3c36cd8, 32'hc3cec599},
  {32'h453d4bf4, 32'hc41bcaa9, 32'hc41d3ebf},
  {32'hc5674bca, 32'hc2a7d12a, 32'h432ce6fa},
  {32'hc2b39d48, 32'h4506aa9b, 32'hc319e09d},
  {32'hc25c3dcd, 32'hc38eb688, 32'hc30738a3},
  {32'h440f0ebc, 32'h44093b28, 32'hc40e6111},
  {32'hc39ee392, 32'hc4f56dbc, 32'hc39c0249},
  {32'h44a3d309, 32'hc386189e, 32'h42b45dc9},
  {32'hc584d084, 32'hc33580d9, 32'h43aaf0ca},
  {32'h457153a4, 32'hc12708cf, 32'h43265273},
  {32'hc2da690a, 32'hc4bba8bc, 32'h4318d0ab},
  {32'h43cf942f, 32'h43aca4a2, 32'h4330423f},
  {32'hc2858fee, 32'hc4281d87, 32'h44290841},
  {32'h454bc27e, 32'h428afd04, 32'hc3678cf2},
  {32'hc4ae56ec, 32'h42e7cd7d, 32'h43ab2f31},
  {32'h43822a5a, 32'h4435806c, 32'h439b0785},
  {32'hc33a6871, 32'hc3a3f5cb, 32'h449c843f},
  {32'h448e915a, 32'hc08c8fb6, 32'hc4b8cefd},
  {32'hc3bd016d, 32'h426ce335, 32'h44017a6f},
  {32'h43de1f0f, 32'hc38c8b39, 32'hc42818b5},
  {32'hc50b8478, 32'hc4a1ded1, 32'hc31b0c3a},
  {32'h441951a0, 32'h451b94f8, 32'hc3ec66fb},
  {32'h43c26cb5, 32'hc42f86f8, 32'h4437a23c},
  {32'h42abc515, 32'h43aec39f, 32'hc3a42e12},
  {32'hc3c66467, 32'hc521ddee, 32'h42ceb4cf},
  {32'h43ec61be, 32'h4413ae96, 32'hc2e0888b},
  {32'hc5800d0f, 32'hc30a9721, 32'h42c65a6a},
  {32'h441dfe79, 32'hc38b87e8, 32'hc53e8f71},
  {32'h43bfa438, 32'hc5149219, 32'hc33cd429},
  {32'hc53f83c2, 32'h440fc2e6, 32'hc24dca3f},
  {32'hc32f1396, 32'hc4dc5129, 32'h439427f4},
  {32'hc49215c5, 32'h44d0f26c, 32'hc3fcf690},
  {32'h42b2c873, 32'hc5427bfb, 32'h433e88bd},
  {32'h440410f5, 32'h450b9332, 32'hc3137bbc},
  {32'h4505e64a, 32'hc40f4b95, 32'h425211d7},
  {32'hc4487ce8, 32'h44104b3f, 32'h43de1bdf},
  {32'hc4a08630, 32'hc258fe80, 32'h43f87548},
  {32'hc489bff4, 32'hc3e4897e, 32'h44b78416},
  {32'h44bfda38, 32'h40d1fcbe, 32'hc38ca0d3},
  {32'hc41ea882, 32'h43aaec2b, 32'hc416621d},
  {32'h443cf6c5, 32'hc4c04d43, 32'h443ead49},
  {32'hc44c1017, 32'h433e2f6d, 32'hc3d325c9},
  {32'hc30e4888, 32'hc4d4c9de, 32'hc343ef79},
  {32'h414c3560, 32'h4496ece1, 32'h4460c313},
  {32'hc313cac4, 32'h4386a92f, 32'h45543e1e},
  {32'h44b7f083, 32'h4389121c, 32'h434785b7},
  {32'hc0990300, 32'hc53f383b, 32'hbc718400},
  {32'hc4767bb4, 32'h448d0ed3, 32'hc4c58284},
  {32'h439e51dc, 32'hc38be605, 32'h43337f25},
  {32'hc2a5c0f0, 32'hc3a28d56, 32'hc4ed5b5a},
  {32'hc2f9c110, 32'hc47ca3ce, 32'h445adc88},
  {32'hc3d98074, 32'h4416c010, 32'hc4dfbc32},
  {32'h44884b23, 32'h440560a2, 32'h44c95a9b},
  {32'hc507e814, 32'h4320ee4d, 32'hc50008f3},
  {32'h451b0744, 32'hc3f3c710, 32'h4308359b},
  {32'hc23ffd30, 32'h43cf620c, 32'hc5026d81},
  {32'hc3a93910, 32'h4486dc4d, 32'h450b6d6d},
  {32'h447d305a, 32'hc303a67e, 32'hc2e06b5b},
  {32'h44408811, 32'h4464d1aa, 32'hc38c3716},
  {32'h445a377f, 32'hc2174057, 32'h44cd8bed},
  {32'hc47bfc4d, 32'hc3e2d149, 32'hc3e0ed1b},
  {32'h43577cfe, 32'hc31d05c9, 32'h44185fb1},
  {32'hc485d25e, 32'h4491da64, 32'hc4981745},
  {32'h44949599, 32'hc427edc7, 32'h448162e3},
  {32'h42ab05d0, 32'hc315a73f, 32'h44e55762},
  {32'hc52ba263, 32'h423ca990, 32'hc30f8375},
  {32'hc466c134, 32'h43adcce7, 32'h43680515},
  {32'h4404b8ee, 32'hc491ff89, 32'h43c0abc7},
  {32'hc41e7f3b, 32'h43b21b71, 32'hc3615f43},
  {32'h44a0a833, 32'h41bfd813, 32'h44877b7e},
  {32'hc3a9ffeb, 32'h442ca036, 32'hc30fbd96},
  {32'h43d84679, 32'hc434e986, 32'h4499482d},
  {32'hc40515ba, 32'hc45c9cfb, 32'hc4cbf335},
  {32'h45697da5, 32'hc332a5c5, 32'h440bcfa5},
  {32'hc53409b6, 32'hc38bfada, 32'hc3acdc61},
  {32'h43eba630, 32'hc406b2f0, 32'hc418d3e8},
  {32'hc4e76514, 32'h42ec7f17, 32'hc35fe356},
  {32'h452969ac, 32'hc44581a6, 32'h42c710dd},
  {32'hc3cf7594, 32'h44d85261, 32'hc223ceb3},
  {32'h44cb9f04, 32'h43bc197f, 32'h43b791f1},
  {32'hc523fa12, 32'h43de0806, 32'hc0120820},
  {32'hc341f92c, 32'hc53a8b78, 32'h43865d72},
  {32'hc4eb5d01, 32'hc39aa116, 32'hc2e16523},
  {32'h42dac990, 32'h4487da97, 32'hc4a2ce5f},
  {32'hc4120381, 32'h44c02393, 32'h44871556},
  {32'hc1d5a980, 32'hc53a67f2, 32'h42b97175},
  {32'h441bb88a, 32'h448e8915, 32'hc07eb65c},
  {32'h43e02c18, 32'hc4d666e5, 32'h40821598},
  {32'hc2262ca0, 32'h44dfc5e1, 32'hc4101edd},
  {32'hc506d23c, 32'hc3b40e69, 32'hc19bdce8},
  {32'h4201df28, 32'h41d8f830, 32'hc32121d6},
  {32'h43e7ce48, 32'hc393ab13, 32'hc4174768},
  {32'hc3b973d7, 32'hc5230770, 32'h44dbde00},
  {32'h40cfa380, 32'hc4063a32, 32'hc4be1342},
  {32'hc322198b, 32'h44fd0db4, 32'hc2f133cd},
  {32'hc4d2ccc8, 32'hc3e4252a, 32'hc2961419},
  {32'h42219f60, 32'h433558f9, 32'hc4cd6753},
  {32'hc4f6be5c, 32'hc39c3530, 32'h43298cea},
  {32'h431913e8, 32'h433dd606, 32'h4169f4f1},
  {32'h4368c213, 32'h43570db7, 32'h45078dd4},
  {32'h44f5e080, 32'hc4027fc2, 32'h43ba24a1},
  {32'hc5088543, 32'h43060391, 32'h42c8bac2},
  {32'h44b833e4, 32'h43ef234c, 32'hc38f8e72},
  {32'hc47939a0, 32'hc4929be2, 32'h42b954e2},
  {32'h45132100, 32'h4401bee1, 32'h439c9470},
  {32'hc1a7ced8, 32'hc4aa307e, 32'h440a6349},
  {32'h44d8278b, 32'h44b70c16, 32'hc3e133d7},
  {32'hc43b4610, 32'hc4d4858f, 32'h43943bf9},
  {32'hc338d24a, 32'h4414351c, 32'hc3a37116},
  {32'h42a41037, 32'hc4a1f629, 32'h436f5e23},
  {32'h44994c55, 32'h44303a0f, 32'hc420b236},
  {32'h44446365, 32'h44306f18, 32'h440a03ff},
  {32'h439a83f3, 32'hc3d9cad4, 32'hc4630eed},
  {32'h44f5648d, 32'h42b3495f, 32'h43a14819},
  {32'hc32eb571, 32'h423f9fba, 32'hc4d156aa},
  {32'h44fe6fc6, 32'hc3bf12d6, 32'hc3813a34},
  {32'hc380af7f, 32'hc2d70924, 32'hc514048d},
  {32'hc23ff8a4, 32'h44391894, 32'h44e8d1fb},
  {32'h43ae5880, 32'h448c4ca0, 32'hc409aa36},
  {32'h433565a4, 32'h44c381ec, 32'h441243b9},
  {32'hc39d0440, 32'hc52c7a4f, 32'hc3d7f56c},
  {32'h42a959c8, 32'hc38eae32, 32'h43283c15},
  {32'hc40ef104, 32'hc4eed140, 32'hc330c3e1},
  {32'hc3127c8c, 32'h441a3d3a, 32'h453d332b},
  {32'h4337bf78, 32'h42c94ae9, 32'h442a1d74},
  {32'h43991b8b, 32'h44d116e5, 32'h4434dfce},
  {32'hc457faae, 32'hc397ef06, 32'hc430cc97},
  {32'hc48d1c60, 32'h43900e51, 32'h43063c2f},
  {32'hc49c273d, 32'hc496edbb, 32'hc4225610},
  {32'h430f3cd8, 32'h455d29b1, 32'hc30a770b},
  {32'hc41649d3, 32'hc456284e, 32'h4358d501},
  {32'h415626c3, 32'h457fc108, 32'h4302e144},
  {32'hc4ccdfaa, 32'hc490ed5b, 32'hc1899527},
  {32'h4531affb, 32'h43515999, 32'hc2d916cf},
  {32'hc567e07b, 32'h438b3320, 32'hc2c28e24},
  {32'h44da4caf, 32'h42cc4f87, 32'hc2bae25e},
  {32'h42d0cfe9, 32'hc2d08c25, 32'hc4b77e34},
  {32'hc45a226c, 32'h4382d35a, 32'h4378500a},
  {32'hc29878c0, 32'hc42f99b0, 32'hc393d470},
  {32'hc4ba82cb, 32'h43e31731, 32'h43ad3abe},
  {32'h43b64d00, 32'hc406c7f3, 32'hc47f15d1},
  {32'hc204e984, 32'h43d55801, 32'h43b7c17c},
  {32'h4421ec4e, 32'hc43b4d58, 32'hc4edd461},
  {32'hc49f8db6, 32'h432abf6f, 32'h448be24e},
  {32'hc308204f, 32'hc429bd5e, 32'hc35ccfae},
  {32'hc465e5f3, 32'hc3c96d71, 32'h4472564d},
  {32'hc3aeb3e0, 32'hc54487b2, 32'hc3fd7d0a},
  {32'hc137a120, 32'hc4b29b0d, 32'h43c354eb},
  {32'h42edf20c, 32'hc53236bf, 32'hc386a91f},
  {32'hc3f1c067, 32'h4502ac17, 32'h43d459e6},
  {32'hc45bbf15, 32'hc415f8f5, 32'hc2e9b091},
  {32'hc442410e, 32'h43fa9d2e, 32'h44d4b18a},
  {32'h44c8fdcd, 32'hc38ca20e, 32'hc42aead8},
  {32'hc51211c4, 32'h432f2e0c, 32'hc1da81be},
  {32'h431627a0, 32'hc4b3a6f8, 32'hc3b01358},
  {32'hc45d1ca8, 32'h4463e26a, 32'h43b0aa59},
  {32'h443cab7c, 32'hc3193bdc, 32'hc33752ea},
  {32'hc4ea5288, 32'h44976648, 32'h42cd49b9},
  {32'h448a0422, 32'hc4a7c546, 32'h419396b7},
  {32'hc438b3de, 32'hc3edbc43, 32'h430265cb},
  {32'h457cb299, 32'h43e9b2a4, 32'h4440530c},
  {32'hc53e432f, 32'hc3d448e0, 32'h42b2550a},
  {32'hc4950a92, 32'hc385813c, 32'hc3941eaa},
  {32'h4528cc10, 32'hc3ae409a, 32'hc4130166},
  {32'hc53a1aef, 32'h4363dc67, 32'hc3a225c2},
  {32'h44950bfc, 32'hc3d61a78, 32'h43711b86},
  {32'hc37de940, 32'h44f939d8, 32'h420bec9e},
  {32'hc09ead00, 32'hc51c5dd4, 32'hc25c32f4},
  {32'hc527d319, 32'hc205cb68, 32'hc23d9c53},
  {32'h451a645d, 32'h43e62926, 32'h43a8d028},
  {32'hc45aa9ec, 32'h447292d9, 32'hc2a0afea},
  {32'h44dbc99c, 32'hc44da604, 32'hc36fb20c},
  {32'hc1c83ce0, 32'h42b1e594, 32'hc47fdf9e},
  {32'h4422cdee, 32'hc318c78f, 32'h41ce8a77},
  {32'hc4f6d07d, 32'hc2998662, 32'h44198b7b},
  {32'h4410b17e, 32'hc4069017, 32'hc385bff4},
  {32'hc4a75756, 32'hc3f14c3c, 32'h438d8c4f},
  {32'h448a502d, 32'hc3e39485, 32'hc4c5af6b},
  {32'hc3a5f55d, 32'h4384003b, 32'h441d8a72},
  {32'hc4407b17, 32'hc50c569f, 32'hc3a2a88b},
  {32'hbe73b800, 32'h44da8d90, 32'h43baa464},
  {32'h448714e4, 32'hc41ef196, 32'hc366d210},
  {32'hc4d46be0, 32'hc3d70b35, 32'h43f57aed},
  {32'h44e31e28, 32'h41deb8a1, 32'hc45b3a83},
  {32'h43f6a91e, 32'hc358e648, 32'h44e1c346},
  {32'hc3f32a32, 32'hc4816139, 32'hc3700c29},
  {32'h42ad9b40, 32'h44b7d52b, 32'h44307bf4},
  {32'h433f8f62, 32'hc4bb2362, 32'hc330e351},
  {32'hc39b2142, 32'h450c8669, 32'h4420d75c},
  {32'hc323ac22, 32'hc49559ba, 32'hc4e73985},
  {32'hc25054c0, 32'hc28819b5, 32'hc50cdf16},
  {32'hc412e9e2, 32'h43ab9996, 32'h442a2d75},
  {32'h44ac6c72, 32'h42417c7f, 32'h43a88c1f},
  {32'hc42897c6, 32'hc46395b0, 32'hc2a7f46b},
  {32'h43f6ad68, 32'h4500248d, 32'h427f02b8},
  {32'hc51b8edc, 32'hc339c35a, 32'hbfc008fc},
  {32'h453dda63, 32'h43fb6f82, 32'h4380f847},
  {32'hc4497198, 32'hc51d9f76, 32'h43d1b3a1},
  {32'h4535620f, 32'hc3d1b0d2, 32'h43202a51},
  {32'hc4d41762, 32'hc45d0f35, 32'hc43e5252},
  {32'h455761d4, 32'hc18f174e, 32'hc30effe5},
  {32'h4429a468, 32'hc3e8b52b, 32'h442c5479},
  {32'h450fed94, 32'h43bca566, 32'h43bdfb1e},
  {32'h43c0b6d6, 32'hc4ceffeb, 32'hc492e0c8},
  {32'h43448ab5, 32'hc293855f, 32'h441ecac4},
  {32'hc2f17380, 32'hc40a5cd8, 32'hc4b132ad},
  {32'h4429f289, 32'h4384d7b5, 32'h44fa8c14},
  {32'hc513a924, 32'hc4201312, 32'hc27f82f5},
  {32'h44d46308, 32'hc39eba1b, 32'h443fa44c},
  {32'hc532e362, 32'h430ff95a, 32'hc331df2c},
  {32'h44fd1159, 32'h436a725f, 32'hc3e3a816},
  {32'h42c6a020, 32'hc5599037, 32'hc38b4996},
  {32'hc3387f6b, 32'h455fafca, 32'hc2825bc4},
  {32'h422fb29d, 32'h42ff0b6a, 32'hc4b8a1c7},
  {32'hc418f944, 32'h44a7a8a5, 32'h44801160},
  {32'h429257fc, 32'hc3bb16d8, 32'hc5290b9a},
  {32'h4349a224, 32'h43ff9f72, 32'hc346a1f0},
  {32'hc49aeace, 32'hc2d6532b, 32'h43450854},
  {32'hc49021e2, 32'hc4903b13, 32'hc3a1f175},
  {32'h440262f2, 32'h4417f1cf, 32'h446fd8dd},
  {32'hc2fef343, 32'h43aa5bca, 32'hc279ab1c},
  {32'h450c5f46, 32'h41ac1846, 32'hc3681821},
  {32'hc462321d, 32'hc3126897, 32'hc42ec77d},
  {32'h44311a87, 32'h43a42f51, 32'hc45195a6},
  {32'hc48cf18f, 32'hc42ce09d, 32'hc342e38e},
  {32'h4510605e, 32'h43cea3f6, 32'h442365bc},
  {32'h4425a97d, 32'hc364f2d7, 32'hc4085185},
  {32'h44aab847, 32'h4404bed8, 32'hc4afa587},
  {32'hc4c46fa3, 32'hc2e517b3, 32'h439fbbb9},
  {32'hc421c04a, 32'h43d5a820, 32'hc18419f1},
  {32'hc4ddeef6, 32'hc2c6769d, 32'hc369a706},
  {32'h44611679, 32'h4398265e, 32'hc4f4c369},
  {32'hc310b9c6, 32'hc35d5918, 32'hc278b0c6},
  {32'h440c9634, 32'h44008e9c, 32'hc392f498},
  {32'hc4a01e9b, 32'h41184415, 32'h44c2f94d},
  {32'h450ac688, 32'h42e725fb, 32'hc3b77572},
  {32'hc378fb90, 32'hc53fa6dd, 32'h4385de90},
  {32'h4497e7ca, 32'h4401b443, 32'hc4550d8f},
  {32'h43852b0f, 32'hc4510b35, 32'h440ed267},
  {32'h43ea4690, 32'h43021f36, 32'hc40ee613},
  {32'hc288bc58, 32'hc50bb8ad, 32'h423ddff5},
  {32'h456e638f, 32'h4374df6f, 32'hc212535b},
  {32'hc512bbee, 32'h437c23f1, 32'h43ab1b89},
  {32'h42ce21c0, 32'hc392f92a, 32'hc4a211df},
  {32'h451bfe10, 32'hc42d6966, 32'hc38f61a2},
  {32'hc4760ee4, 32'h43e15520, 32'h44038e66},
  {32'h43cfe714, 32'h441535e0, 32'hc45d4959},
  {32'hc4d7f1c2, 32'h448ddbc0, 32'h4384fb0a},
  {32'h43988a90, 32'hc48aad25, 32'h44471284},
  {32'h44d18712, 32'h433aa23b, 32'hc2f8325e},
  {32'h453c9734, 32'h43fd8446, 32'hc30679e7},
  {32'hc48bed7c, 32'hc2581baf, 32'h41760e6c},
  {32'hc463b102, 32'hc2911d7e, 32'hc294921c},
  {32'hc4058c32, 32'h44c059b8, 32'hc405f430},
  {32'h44714538, 32'hc47228ba, 32'h44cba815},
  {32'h420c4cc6, 32'h44ecc097, 32'h42cbfb18},
  {32'h42c0c28a, 32'hc550dfb6, 32'h430bc3c2},
  {32'hc40cf104, 32'h439a9d9e, 32'hc4ba7035},
  {32'hc3ca3cd3, 32'hc491bc36, 32'hc396f9df},
  {32'hc4541647, 32'hc2add538, 32'hc42fbbc2},
  {32'h4477fd0b, 32'hc21be3c1, 32'h44839967},
  {32'h44af3f76, 32'hc40f4022, 32'hc43c4337},
  {32'h445d0cf7, 32'hc4a48458, 32'hc38f330c},
  {32'hc4325230, 32'h4534f90a, 32'hc2ed238e},
  {32'hc3184124, 32'hc49782ea, 32'hc32599f5},
  {32'hc3449420, 32'h439ca9ae, 32'hc50d39ae},
  {32'h44830326, 32'hc333cd57, 32'h440d416b},
  {32'h44dc54dc, 32'hc291ddcc, 32'hc2241f68},
  {32'h456140c8, 32'h43ea4461, 32'h439b09b2},
  {32'hc4bc9b77, 32'hc35e1350, 32'hc50d5a20},
  {32'hc446a634, 32'hc3077114, 32'h441347da},
  {32'hc4898cc5, 32'h43e1b233, 32'hc48ae25f},
  {32'h43edb2b5, 32'h44392c76, 32'h44e1009d},
  {32'h4259de35, 32'h43ab4ecd, 32'hc47dd1b7},
  {32'h4400460d, 32'h43ccc19a, 32'hc44f9d51},
  {32'h449eccb7, 32'h42d9d878, 32'h4489c84f},
  {32'hc37a60e3, 32'h44d07e69, 32'hc300c3bd},
  {32'h43d5f5b6, 32'h43a42125, 32'h44df3130},
  {32'hc400324c, 32'h436d2592, 32'hc4a5f8ab},
  {32'h433655b0, 32'hc5051f7b, 32'h43b6fa03},
  {32'h4459c6b0, 32'h4320fce8, 32'h44a07d87},
  {32'h4399bebc, 32'hc4c6707b, 32'hc506f5c5},
  {32'h443fc6d9, 32'h439c54d2, 32'h43d4aa35},
  {32'hc432c887, 32'hc4367a75, 32'h43eeddb2},
  {32'h4390707e, 32'h453e44d9, 32'h4401f463},
  {32'h450cb939, 32'hc302d76e, 32'h43efdf72},
  {32'hc388eb0e, 32'h4482e0de, 32'h43f9741b},
  {32'h43f2e83c, 32'h43ad6379, 32'h44e30fe2},
  {32'hc470db8c, 32'h42844ef2, 32'hc459675e},
  {32'h4538127e, 32'hc383120d, 32'hc2a587e7},
  {32'hc4ffd9ec, 32'hc25eb65f, 32'h425cbc8b},
  {32'h4557acae, 32'hc3335a2e, 32'hc21420dc},
  {32'hc3ecaa80, 32'h446f3ce2, 32'h441ddaa7},
  {32'h4373ae14, 32'hc5047abd, 32'hc334af19},
  {32'hc445fe23, 32'h44931116, 32'h43c52a59},
  {32'hc4c162b5, 32'hc2893204, 32'hc3f8e94b},
  {32'hc4850cbe, 32'h44a9b33d, 32'hc403f20a},
  {32'hc2ed5fff, 32'hc53ba885, 32'hc33e4d23},
  {32'h43ddf036, 32'hc34a1bb6, 32'h44c80a41},
  {32'hc3913d71, 32'h44a3f2fb, 32'hc501acfd},
  {32'hc2c3a2d0, 32'h423f0258, 32'h4562b995},
  {32'hc2ab8675, 32'hc2e284db, 32'h44b87c51},
  {32'h4466b4b2, 32'h440f8a92, 32'hc3e788dd},
  {32'h44c4c96b, 32'h4311f73b, 32'hc211f942},
  {32'h4374c9b0, 32'h43b4481a, 32'hc5081ba6},
  {32'hc48fde1c, 32'hc39939b4, 32'h439f365c},
  {32'hc4097286, 32'h44b6d349, 32'hc254cfae},
  {32'h4420d91d, 32'hc3d2cb86, 32'hc336e7cf},
  {32'hc4296ec2, 32'h44396c36, 32'h44ed8cc2},
  {32'h4448601c, 32'h4475a0bc, 32'hc4c529ff},
  {32'h4398d4eb, 32'h4422c00d, 32'hc2f63357},
  {32'hc50db038, 32'hc3f4dd77, 32'h429e4536},
  {32'hc4a1cab7, 32'h43f3cbc9, 32'h43097fbb},
  {32'hc439529b, 32'hc43eddab, 32'h44b27358},
  {32'hc3afb5ce, 32'h44e77f3e, 32'hc3ccb0ca},
  {32'hc4550a46, 32'hc43a8de2, 32'h43e18cca},
  {32'h4554d6ed, 32'hc1a15626, 32'h43bb5a94},
  {32'hc58f378c, 32'h43845e6b, 32'h4270133c},
  {32'h457f1e04, 32'hc33fe39f, 32'hc3d9b0a2},
  {32'hc4791e1c, 32'hc4da2593, 32'h43452c63},
  {32'h4481b2ec, 32'h44f6fe94, 32'hc30ca30c},
  {32'h43a38051, 32'hc498c0a4, 32'h4334995b},
  {32'h43dd9e9c, 32'h4503da0b, 32'hc4301006},
  {32'hc3da704e, 32'hc52468e9, 32'hc237c110},
  {32'hc1ba8600, 32'hc0b90534, 32'hc3cb3f21},
  {32'hc24875d5, 32'h42634565, 32'h44512150},
  {32'hc492ed29, 32'h440957f0, 32'hc3996f42},
  {32'hc3a739f2, 32'hc43de639, 32'h449e51b4},
  {32'h42fa0e4a, 32'hc4364576, 32'hc36fa75c},
  {32'h45380e3f, 32'h4425369c, 32'h40b6cee6},
  {32'h4415ad26, 32'hc3d2ee21, 32'hc4e43be7},
  {32'hc3f8be08, 32'h448bfc16, 32'h43aa0784},
  {32'hc309767d, 32'hc3912cf9, 32'hc530c79c},
  {32'h454441b8, 32'h42cb9bb2, 32'h434ed069},
  {32'h44b38920, 32'h448b9847, 32'hc3f0a193},
  {32'hc37c271e, 32'h44b1b07e, 32'h43ec05fc},
  {32'hc45ff706, 32'h421476f1, 32'hc47525d3},
  {32'hc4847ac6, 32'h42c02e53, 32'h44039a1a},
  {32'hc39bab64, 32'hc4c103d6, 32'hc41a9945},
  {32'h447f33aa, 32'h43732165, 32'h4480d938},
  {32'h446d4ae9, 32'hc3cc42a2, 32'hc4bc1932},
  {32'h44c70bb5, 32'h43759539, 32'h44a97d89},
  {32'hc354d840, 32'hc48c3307, 32'hc4602687},
  {32'hc4977947, 32'h44264044, 32'h4382ff27},
  {32'hc4106326, 32'hc4b84f9f, 32'hc3ab1fae},
  {32'hc34ee940, 32'h45505b2e, 32'h44106885},
  {32'h42da32b0, 32'hc3e186e7, 32'hc3c321a6},
  {32'h42b1d4fc, 32'h451dfa31, 32'hc30b6595},
  {32'hc389c9c8, 32'hc43296f6, 32'hc3397084},
  {32'h450aedf9, 32'h43539ae7, 32'hc2662a4f},
  {32'hc5540a14, 32'hc330f400, 32'h42f4ea8f},
  {32'h4555ac90, 32'h43835acf, 32'hc373a115},
  {32'hc3106f9b, 32'h4505f021, 32'hc4aab887},
  {32'h3d26cc00, 32'hc3cb1a9a, 32'h44bf5aa6},
  {32'h441d6259, 32'hc4ecc0f5, 32'hc36a17e7},
  {32'hc3b0b3f3, 32'h43c16753, 32'h4481af7b},
  {32'h43625b96, 32'hc468287b, 32'hc4bafb4f},
  {32'h44bbee60, 32'h4433f75d, 32'h43c9d78b},
  {32'hc3d5ba7d, 32'hc51623aa, 32'hc4de1d0b},
  {32'hc44cdd0b, 32'h4446527e, 32'h450055bd},
  {32'h4412abe9, 32'hc3b708a9, 32'h42511a10},
  {32'h438856a0, 32'h4428f920, 32'h449ed8fc},
  {32'h4428cf00, 32'hc309e790, 32'hc3aaebc2},
  {32'h4400f7c2, 32'hc41dcc26, 32'h442f2edc},
  {32'h44bc00b4, 32'hc2d741b3, 32'hc387f3cf},
  {32'hc4b1ca24, 32'h44826afe, 32'hc3168530},
  {32'hc3ddc9e2, 32'hc41cb4f7, 32'hc1daba65},
  {32'hc43ba0e8, 32'h448e0b64, 32'h44916dcd},
  {32'h4505c0bb, 32'hc43dc37b, 32'hc3cde3b7},
  {32'h4283e240, 32'h4430f734, 32'h440a4416},
  {32'h455c848a, 32'hc3d9f055, 32'h440ee402},
  {32'hc1e293f0, 32'h4556c60e, 32'hc29d8306},
  {32'h43c8e9df, 32'hc3894946, 32'h413c0968},
  {32'hc512e6f8, 32'h44bad155, 32'h439718a3},
  {32'h446ce3a4, 32'hc3dcfadb, 32'hc39ee8af},
  {32'hc437e93c, 32'hc3cc9490, 32'hc131aec3},
  {32'h44d9a172, 32'h439e2078, 32'h43139f57},
  {32'hc4978e3c, 32'hc35ae135, 32'h438fdc72},
  {32'h4311c73d, 32'hc3814a58, 32'hc3aa5391},
  {32'h45013271, 32'hc39b87aa, 32'hc3abb191},
  {32'hc572445c, 32'h41dc46eb, 32'hc2f3e2e8},
  {32'h44a1a0a8, 32'h430ffc8b, 32'h4494e8a7},
  {32'h44aa2798, 32'h4434398d, 32'hc2f464f1},
  {32'h446bdedb, 32'hc489eeff, 32'h44006fd3},
  {32'hc3dd4364, 32'h45046178, 32'h42c61c7e},
  {32'h448fa713, 32'h426a3d86, 32'h438e87e8},
  {32'hc55b4ac5, 32'hc21a6684, 32'hc2b16d07},
  {32'h443c80c0, 32'hc5260415, 32'h4303021a},
  {32'hc3e582a6, 32'h42c4fa2c, 32'hc3989f19},
  {32'h43a73573, 32'h42e8c5eb, 32'h4431c794},
  {32'hc4e855c2, 32'h426d5428, 32'hc4370785},
  {32'hc37e3596, 32'hc30ec728, 32'hc4892f79},
  {32'h41c50e37, 32'h440960ef, 32'h443752e7},
  {32'hc391a13a, 32'hc4a26ec4, 32'hc51ae304},
  {32'h43296d8b, 32'h44dfdba4, 32'h429253d9},
  {32'h423e8ae0, 32'hc4a385a8, 32'hc28a86c8},
  {32'hc4ddd183, 32'h43375f17, 32'hc33d71dc},
  {32'h44498f9e, 32'hc4155d80, 32'hc3cf2aaf},
  {32'hc5044e32, 32'hc4105018, 32'h43bddae9},
  {32'h442d6372, 32'h4355b1a3, 32'hc3f3565f},
  {32'hc366173b, 32'h442e9638, 32'h42ae3573},
  {32'h42c05eb0, 32'hc4da998a, 32'hc3fa6110},
  {32'hc531670e, 32'hc2332372, 32'h42998b64},
  {32'h441be567, 32'hc4859aea, 32'hc1f94109},
  {32'hc44903f0, 32'h45451cea, 32'h435fca7d},
  {32'h44a4fc7d, 32'hc3e03b53, 32'hc4fdb02f},
  {32'hc3066580, 32'hc2d5c2b8, 32'hc53974bb},
  {32'hc5685054, 32'h41bf72a0, 32'h430c5ac6},
  {32'hbf8d8400, 32'h43d96c66, 32'h4113ba70},
  {32'hc4a6d39c, 32'hc388e6e2, 32'h43fb5bfc},
  {32'h449b3084, 32'h43e50680, 32'hc387a181},
  {32'hc4290c86, 32'hc414edba, 32'h440f2081},
  {32'h44502da7, 32'h4552c16d, 32'h4422a15e},
  {32'hc382adbe, 32'hc4b0b164, 32'hc3c5a2c1},
  {32'h432dab57, 32'h4500081b, 32'hc3472023},
  {32'hc2625770, 32'hc1f97d91, 32'hc315352e},
  {32'h433e0ea0, 32'hc460b5b6, 32'hc5055331},
  {32'h449e9e34, 32'h439b582c, 32'hc155c788},
  {32'h43653afc, 32'h44da0724, 32'h431465b1},
  {32'hc4e1e4e4, 32'hc38a169f, 32'hc44ebd88},
  {32'hc4923e5e, 32'h44191603, 32'h4396e1dd},
  {32'hc44feda2, 32'hc3a51d77, 32'hc450b627},
  {32'h43bc6a0b, 32'h4481960c, 32'h449306f7},
  {32'h440235e8, 32'hc473a645, 32'hc4612dfd},
  {32'h440e6d64, 32'hc3bb91c7, 32'h444f89ff},
  {32'hc4fb3582, 32'hc4825188, 32'hc42f0257},
  {32'h45672375, 32'h441923ac, 32'hc24541c8},
  {32'hc4f1fa78, 32'hc3dbfed4, 32'hc36435b8},
  {32'h447d970c, 32'h42ead5af, 32'h438ba5be},
  {32'h43264a8d, 32'hc31d4058, 32'hc454e4f5},
  {32'h43252f20, 32'h450fad25, 32'h43d41570},
  {32'hc4872635, 32'hc3e5d00a, 32'hc4db68e2},
  {32'h44ca3ecd, 32'hbee4185c, 32'hc3a5e0ac},
  {32'hc3f07a12, 32'h4474789b, 32'h43bd3bb1},
  {32'hc4176158, 32'hc4b57c9f, 32'h4284546b},
  {32'h44948eb7, 32'h44a408ac, 32'h43ab5161},
  {32'hc2755920, 32'hc484aaaa, 32'h42a2749c},
  {32'h44de64fa, 32'hc3f084e6, 32'h42c504ee},
  {32'hc460a370, 32'hc4f7dc7a, 32'hc3b153a2},
  {32'h42cda63e, 32'hc31a5e7b, 32'h428582ad},
  {32'hc5848d3e, 32'h440c0e7e, 32'hc3d0d5c7},
  {32'h44792b64, 32'hc3fbfd83, 32'hc3926c4b},
  {32'h43ade479, 32'h43898ed8, 32'h449a4279},
  {32'h432f1104, 32'h443164d9, 32'hc420f918},
  {32'h4380c2b6, 32'hc52a6524, 32'hc3052d57},
  {32'h4521afdc, 32'h437b22e8, 32'hc3e27254},
  {32'h42aef01c, 32'hc386eb7c, 32'h4509d987},
  {32'h44b1ed51, 32'h448e5160, 32'hc2579848},
  {32'h4500c866, 32'h423e15ab, 32'h42bb7c80},
  {32'h449f03dc, 32'h3f668990, 32'hc4973699},
  {32'hc47076a1, 32'hc2b3aa9a, 32'h4475a4ab},
  {32'h43e6d79b, 32'h4469d8ce, 32'hc389e580},
  {32'hc50b3119, 32'hc383cee6, 32'h42d7e843},
  {32'h44467648, 32'h44f7f308, 32'hc345c133},
  {32'h4485baee, 32'hc43be78a, 32'h437ad38f},
  {32'h44f1a596, 32'h43ed442e, 32'hc3fdffc4},
  {32'hc1a063c0, 32'hc4bab4e8, 32'h434820d9},
  {32'hc4da617c, 32'hc3429072, 32'h42e57b4c},
  {32'hc4beab73, 32'hc3e597e8, 32'h43eccec9},
  {32'h4565ba1a, 32'hc2e36360, 32'hc490366a},
  {32'h43d4db68, 32'hc2fd9132, 32'hc485e699},
  {32'hc387e069, 32'h45187c77, 32'h438188e7},
  {32'h4329524a, 32'hc479ceeb, 32'hc3f055ab},
  {32'hc34d6060, 32'h45148491, 32'hc36a4aed},
  {32'h44ee0f26, 32'hc29b2796, 32'hc2a3e28b},
  {32'hc42cfb7f, 32'h4446d166, 32'h4358b47e},
  {32'h438a4033, 32'hc47c1c8e, 32'hc4bd5fab},
  {32'hc588f3f2, 32'h44161457, 32'hc29f43da},
  {32'hc455e1c8, 32'hc445c344, 32'hc3740585},
  {32'h426879ae, 32'h440befef, 32'h42871d31},
  {32'h438234d9, 32'h43b98b6d, 32'hc4578665},
  {32'h448b4424, 32'h439f2e00, 32'hc445d14f},
  {32'h44020f8a, 32'hc4245686, 32'h431571c7},
  {32'hc3810028, 32'h44544fb9, 32'hc45ee5c4},
  {32'h44204009, 32'h433bdbd4, 32'h438cf4af},
  {32'hc292e816, 32'hc3e59215, 32'hc55198f8},
  {32'h442e9f44, 32'h43093cd8, 32'h4493efab},
  {32'hc482bd82, 32'h44206c1e, 32'h4356dcfd},
  {32'h42cc9fd8, 32'hc4f9eb6d, 32'h43d82404},
  {32'hc4850210, 32'h44ec8f43, 32'hc41e88b2},
  {32'h43bf8420, 32'hc4249800, 32'h433fee36},
  {32'hc4390519, 32'hc391e91e, 32'hc4f29e5e},
  {32'h45020dd5, 32'h42a7b50e, 32'h442cf2bb},
  {32'h42e7a494, 32'hc381966a, 32'hc4345a51},
  {32'h4509fd38, 32'h41535bec, 32'h443bb3c3},
  {32'hc490d2e1, 32'h4397435f, 32'hc4d87fbb},
  {32'hc4fb31ba, 32'h4056a02c, 32'h43dd8502},
  {32'hc300dc7d, 32'h44e280e2, 32'hc4e84872},
  {32'h448c127b, 32'hc463a91e, 32'h43275ceb},
  {32'hc44c3b57, 32'hc4928430, 32'hc29bdb12},
  {32'hc4fabd1f, 32'hc38cce02, 32'h414fc45b},
  {32'h44034a74, 32'h41ef819a, 32'h447f8c86},
  {32'hc446543b, 32'hc2e88d13, 32'hc50059bc},
  {32'h42d6bb09, 32'h4381d9ab, 32'h44eb8ffe},
  {32'hc4b8cc32, 32'h43ebbcc5, 32'hc38b09ae},
  {32'h438fb19c, 32'hc5226a20, 32'h4436fb65},
  {32'h432b5060, 32'hc40d31d0, 32'h45047332},
  {32'hc3e1788c, 32'hc4e90646, 32'hc40f3c30},
  {32'h43ebb1ef, 32'hc3831826, 32'h4388f846},
  {32'hc3cfa94b, 32'h436e2bbe, 32'h44652bad},
  {32'h42f82d38, 32'h42ddeef7, 32'hc4f75744},
  {32'h4491d2f7, 32'hc4c7dedf, 32'hc31f0ce1},
  {32'hc3b832b8, 32'h4399e87a, 32'hc40d7061},
  {32'h440c8589, 32'h43a2710c, 32'h4529c5ed},
  {32'h4389c220, 32'h449e7ce8, 32'hc428e44a},
  {32'h45802e5f, 32'hc37eb06d, 32'h42c15f66},
  {32'hc57462c3, 32'h43dee4bf, 32'hc39eb1ec},
  {32'h451653b9, 32'hc1f97c42, 32'h42b4e94b},
  {32'hc54d1777, 32'h42f15439, 32'h424dd734},
  {32'h44f96add, 32'hc4aced13, 32'hc34fc4d1},
  {32'hc49bd584, 32'h440a3fe6, 32'h436e9836},
  {32'h435e5660, 32'hc4e26bea, 32'h42bec5f8},
  {32'hc4fb3d41, 32'h445a81cc, 32'hc35d015f},
  {32'h452b4452, 32'hc496ec12, 32'hc3bc9a78},
  {32'h43b2cede, 32'hc274d91d, 32'h44642fdb},
  {32'h43779f18, 32'h44136d28, 32'hc4b308a6},
  {32'hc3e377a5, 32'h439ed4a8, 32'h445c0fdd},
  {32'hc4cbc93f, 32'hc47dbdc0, 32'h43bc6701},
  {32'h43c08997, 32'h43dfe8e5, 32'hc4b95eed},
  {32'hc471724f, 32'hc4415ea8, 32'hc30c59cf},
  {32'h441de966, 32'h4417458c, 32'hc51efeac},
  {32'hc4967619, 32'hc40a4781, 32'h4434f4a7},
  {32'hc4553f84, 32'hc348384a, 32'hc4255a32},
  {32'h43e6b658, 32'h4358fe1f, 32'hc502c12f},
  {32'hc4dec43f, 32'hc30e2f76, 32'h4403f3cf},
  {32'hc3f05c54, 32'h43fac740, 32'hc538180b},
  {32'h43c03811, 32'h43beb83e, 32'hc4b96ed7},
  {32'hc27010a8, 32'hc5393389, 32'hc413cafa},
  {32'hc48ead83, 32'h4333c9fe, 32'hc3f4b18e},
  {32'hc46889d9, 32'hc429ad73, 32'h44612eee},
  {32'hc3db4020, 32'hc3120780, 32'hc4ed9f0a},
  {32'hc422424e, 32'hc3f078d7, 32'h43157d87},
  {32'h4543529e, 32'hc3e15bf4, 32'h435a491e},
  {32'hc4f7aa39, 32'h421aa8bc, 32'h413dfe84},
  {32'h4535db07, 32'h43519046, 32'h4380aba8},
  {32'hc42291dc, 32'hc4a77bae, 32'h432726dd},
  {32'h44c4a5df, 32'h44330a98, 32'hc1b88f78},
  {32'hc513e995, 32'hc3846e8f, 32'h4200ee43},
  {32'h43173862, 32'h44f366b2, 32'h4402e2f5},
  {32'hc416f316, 32'hc4c1a81f, 32'h43dda6ab},
  {32'h449fcc18, 32'h444998d3, 32'h42a31d26},
  {32'h44a436be, 32'h41ce468d, 32'h434815bc},
  {32'h4225877c, 32'h447a38d0, 32'hc50eb8a7},
  {32'h4427427a, 32'h431259de, 32'h44a1b333},
  {32'hc4563d82, 32'h42953d18, 32'h43f315a5},
  {32'h4558db20, 32'h4260fdad, 32'h444a0afb},
  {32'hc48f2e70, 32'hc393b10f, 32'hc3fbfa9b},
  {32'hc409c6a1, 32'hc35ad4a0, 32'h444e34cf},
  {32'hc4f5fe58, 32'hc436dc15, 32'hc4b301c8},
  {32'h451bcb0d, 32'h4406c375, 32'h43eff780},
  {32'hc26e96b2, 32'h42dc5565, 32'hc2ec58ff},
  {32'h42b6b338, 32'h4500d73b, 32'h42d9515e},
  {32'hc49aa13c, 32'h4351cf6e, 32'hc440670d},
  {32'hc37ec785, 32'h44afe68f, 32'h428404d3},
  {32'hc54c4ff2, 32'hc30fa317, 32'h437aafc4},
  {32'h451a3bba, 32'h4414a880, 32'hc29ae546},
  {32'h44a1a524, 32'hc44f06fe, 32'hc387777c},
  {32'hc3ddd973, 32'hc3bc6ea0, 32'h43c3c33b},
  {32'hc376b580, 32'hc500c577, 32'hc4b1b0de},
  {32'h452c6c06, 32'hc3f66729, 32'hc1f6582e},
  {32'hc3f0d1b0, 32'hc425e458, 32'hc1a22c04},
  {32'h44de1a16, 32'h4488abf1, 32'h443369e9},
  {32'hc3739f24, 32'hc4bcd548, 32'h431b4244},
  {32'hc412ef0a, 32'h4565d2c5, 32'h42307d5d},
  {32'hc42883eb, 32'hc4b14cc1, 32'hc38656a6},
  {32'hc348e348, 32'h41bb8206, 32'h424e4b51},
  {32'hc445c370, 32'h440dbac3, 32'h43afc8a3},
  {32'hc4000b98, 32'hc40acd21, 32'hc434daa2},
  {32'h43b1bea8, 32'hc3f2a0c5, 32'hc46d4505},
  {32'h42166798, 32'hc4f65f88, 32'h44c27f09},
  {32'hc492fbfa, 32'h4429a986, 32'hc475ee39},
  {32'hc48e0c66, 32'h42b29abb, 32'h43b5f4c9},
  {32'h44429ec2, 32'hc4b895f5, 32'h43b42889},
  {32'h44202d79, 32'h44dc41ca, 32'hc343224c},
  {32'hc2c23e97, 32'hc4b54dfe, 32'hc4b1e043},
  {32'hc466216c, 32'h43e07075, 32'h450cbf5c},
  {32'h452c887e, 32'hc225f553, 32'h40b72a91},
  {32'hc405f968, 32'h43968a7d, 32'h4481951f},
  {32'hc380f31d, 32'h449aae35, 32'hc4fe572a},
  {32'hc311cb66, 32'hc4a2e956, 32'h4399aaa6},
  {32'h433bbdb4, 32'hc5355380, 32'hc29f58aa},
  {32'hc40756c6, 32'h44c0c69e, 32'h442bef95},
  {32'hc1bf4a06, 32'hc3864635, 32'hc2a931f0},
  {32'hc4881e0c, 32'h446508cc, 32'h44604d8b},
  {32'hc2a7c78c, 32'hc4f0a747, 32'hc521811d},
  {32'hc4f621f5, 32'h43776b17, 32'hc35757d9},
  {32'h42e38a54, 32'hc55ca33b, 32'h43659038},
  {32'hc299a7e4, 32'h45294709, 32'h4401c808},
  {32'h44b106aa, 32'hc3a87959, 32'hc3abb867},
  {32'hc41593e0, 32'h44a4a740, 32'hc30bd5a5},
  {32'h449bd817, 32'hc4c4bbd1, 32'h42db4079},
  {32'h444eac23, 32'hc39a5a75, 32'h44280cd9},
  {32'h43d2ff44, 32'hc2710d5f, 32'hc3626167},
  {32'hc402e6ec, 32'hc3276e9d, 32'h43cf74bc},
  {32'h45627e3c, 32'hc2f9e907, 32'h4313e956},
  {32'h45015768, 32'h420138b3, 32'hc3b7b801},
  {32'hc5867f50, 32'hc3ac9b0c, 32'hc2e7487c},
  {32'h4512aab3, 32'h4380bb29, 32'h43038e1a},
  {32'h449d79cc, 32'h4374aedd, 32'h439d45b3},
  {32'h44498b82, 32'hc53a00e6, 32'h428c6a8c},
  {32'hc463d5f4, 32'h439bc344, 32'h43849761},
  {32'hc43ae2d8, 32'hc469209d, 32'h432e9fa6},
  {32'hc39196be, 32'h452e7b99, 32'hc2fabd7c},
  {32'h448d306e, 32'hc4301523, 32'h4154704e},
  {32'h45053a49, 32'hc3bf7ceb, 32'hc239b092},
  {32'h44faacf2, 32'hc316553e, 32'h439fd730},
  {32'hc3ed80f0, 32'hc3931e09, 32'h429d5fc8},
  {32'h4503fc80, 32'hc387e88a, 32'hc2d02460},
  {32'hc480772a, 32'h4371014e, 32'h43b873ed},
  {32'h445b58e4, 32'hc41d6a1b, 32'hc44fb481},
  {32'h43a2d6d1, 32'h44154c07, 32'h43d60e5a},
  {32'h432c5579, 32'h443081ce, 32'hc50c19c2},
  {32'hc2699470, 32'h4422a04c, 32'h4508c556},
  {32'h4519f219, 32'hc2efc670, 32'hc392030b},
  {32'hc57a0f98, 32'h42a2baf6, 32'h43b4a6cd},
  {32'h432051ce, 32'h443953d1, 32'hc4a493c9},
  {32'hc445358e, 32'h4335119a, 32'hc3810647},
  {32'h44a53244, 32'hc3fa66a5, 32'h43518f85},
  {32'h43dac38e, 32'h452f001e, 32'h433b270d},
  {32'hc459f0ea, 32'hc3bfbbae, 32'hc438f3e0},
  {32'hc38b4eda, 32'h44aff69f, 32'h437c01d7},
  {32'h4526d4bc, 32'hc355f612, 32'hc34e3496},
  {32'h45148e86, 32'hc395aa8d, 32'hc44f1f50},
  {32'hc5181b4b, 32'h425fe135, 32'h442275cc},
  {32'h4456ed73, 32'hc1be0099, 32'hc4812175},
  {32'hc451a82a, 32'hc4848f2c, 32'hc3fc836e},
  {32'h43142211, 32'h4522edcc, 32'hc226aa48},
  {32'h442a42e1, 32'hc50053fd, 32'hc0a38e00},
  {32'h42c08010, 32'h43f8adbf, 32'hc35f4cb7},
  {32'hc22b3d5c, 32'hc57d34d8, 32'h4317b6db},
  {32'h4476b017, 32'hc2b3c25d, 32'h432c2ad0},
  {32'hc51c53cc, 32'hc325a28d, 32'h43388ef5},
  {32'h44bf01ea, 32'hc4536331, 32'h4425cdb3},
  {32'hc4f329c7, 32'hc245cc25, 32'hc1aeb970},
  {32'hc35fa08c, 32'h444f5fd8, 32'h4493e275},
  {32'hc41d5e4b, 32'hc38839c9, 32'hc56d0839},
  {32'h4453ce93, 32'h43e37c3e, 32'h420bfc3b},
  {32'hc34cd7d0, 32'hc4b2a75e, 32'hc385fd46},
  {32'hc32aca60, 32'h446cfc7b, 32'h44b26417},
  {32'h443de835, 32'hc4181ca1, 32'hc3af3475},
  {32'h4521d819, 32'h42d17b22, 32'h43dd731c},
  {32'hc581d7ba, 32'hc2cd54b3, 32'h4147aa84},
  {32'h452ae54f, 32'hc3300918, 32'hc41802f9},
  {32'h432061fb, 32'hc47db432, 32'hc5031f0a},
  {32'h44b0b37a, 32'h43913734, 32'h4334ff7d},
  {32'hc4013b94, 32'hc37fdbe5, 32'h431d75cd},
  {32'h428a69a7, 32'h4436f56d, 32'h443871e4},
  {32'hc4d48028, 32'hc3d748aa, 32'hc3e8a1b4},
  {32'h447468a2, 32'hc373e5b4, 32'h43030dcc},
  {32'h44d18ba8, 32'hc2eee8f0, 32'hc3ae6fd8},
  {32'hc48f132f, 32'hc480f31b, 32'h441a942d},
  {32'h43b024de, 32'h4501bb67, 32'hc337647f},
  {32'h42972af1, 32'hc42b1b9a, 32'hc2b3d9be},
  {32'h4522ca83, 32'h4336e618, 32'hc38a2917},
  {32'hc4c45df5, 32'hc44223d8, 32'h42a12379},
  {32'h4449aa34, 32'h43e62239, 32'h4159e3c8},
  {32'hc544a9d6, 32'hc3e2bed9, 32'h4316adf6},
  {32'h45579a1a, 32'hc3a5c45a, 32'hc3110c52},
  {32'hc484350b, 32'hc34f4fe9, 32'h43b02dc2},
  {32'h40c27e00, 32'h44994b6e, 32'h432261b2},
  {32'hc4ede87b, 32'hc3611bb6, 32'h42b5d491},
  {32'h44fa414c, 32'hc26bb07f, 32'h40379488},
  {32'hc3c19f2a, 32'hc4db235b, 32'h43eaf6c8},
  {32'h434f92c4, 32'h44b1526e, 32'hc481a29c},
  {32'hc5321304, 32'hc36b8e35, 32'h43c46ee4},
  {32'h455c936b, 32'h43cbed58, 32'hc3f1be56},
  {32'hc4a6f485, 32'h43cb905a, 32'h4483855f},
  {32'hc497a590, 32'h42df7fa0, 32'hc3c3c7a6},
  {32'hc4bc6c3b, 32'hc493e986, 32'h43ea9856},
  {32'h45106481, 32'h4488e273, 32'hc3c79764},
  {32'hbfee2800, 32'hc332400a, 32'h44184cdc},
  {32'h4394ae70, 32'h44d12969, 32'hc393f86b},
  {32'hc2f86860, 32'hc4c4b370, 32'h448020e5},
  {32'hc4817994, 32'h430371fd, 32'hc28411c6},
  {32'hc504ce13, 32'h42211e89, 32'h44b4a82d},
  {32'h4549a7a8, 32'hc3119af1, 32'hc475aebd},
  {32'h4538555f, 32'hc424c1a8, 32'hc43cac93},
  {32'hc5795a46, 32'hc19c5c6e, 32'hc38b4373},
  {32'h45257bf2, 32'h437c124b, 32'h437d11d2},
  {32'hc50863f0, 32'h44650b9b, 32'hc2682fae},
  {32'hc386badc, 32'hc501eac9, 32'h441390eb},
  {32'hc53e5535, 32'hc3ec2c55, 32'h439c9525},
  {32'h44f26a4c, 32'h443c7c01, 32'hc31fd02e},
  {32'hc58378e3, 32'hc2cab704, 32'h42f5eeed},
  {32'h451efbdf, 32'hc30367df, 32'h44029551},
  {32'hc5126a34, 32'hc3c0f94e, 32'h42d4d053},
  {32'h436ab390, 32'h43f6cf19, 32'hc46b3f1b},
  {32'hc44582ae, 32'h447224ae, 32'hc2c8949f},
  {32'h450262fe, 32'h43c5088d, 32'h446bb508},
  {32'hc412c0a3, 32'hc384565f, 32'hc4ecdd30},
  {32'hc3d90315, 32'hc34a33f0, 32'h4250adf5},
  {32'hc3a3698e, 32'hc339d826, 32'hc487f23b},
  {32'h4544ba97, 32'hc408bf5d, 32'h409d83ec},
  {32'h42eeee88, 32'hc39012c3, 32'hc449085c},
  {32'h4468d258, 32'hc450079a, 32'h44a5fdb6},
  {32'hc34ece5b, 32'h447d4b6f, 32'hc536b719},
  {32'h453143fa, 32'h43a20f4a, 32'hc409a6c8},
  {32'hc3281acd, 32'h433f8ab2, 32'hc505bf56},
  {32'h42ea4558, 32'hc4f9ac06, 32'h43d13923},
  {32'hc53962cc, 32'hc1a62039, 32'h43a21212},
  {32'h45471bba, 32'h42c9b938, 32'h41f28108},
  {32'hc50cf661, 32'h4317315d, 32'h43225138},
  {32'h455aacea, 32'hc342c408, 32'hc40c120e},
  {32'h41d7a910, 32'hc37361fe, 32'hc4326cb5},
  {32'hc285ec2c, 32'h44efe64f, 32'h44c08929},
  {32'h44844842, 32'hc201492e, 32'h44060c9f},
  {32'h4400f850, 32'h44cfd19a, 32'hc3abd713},
  {32'h4511a30f, 32'h42a05701, 32'h42f18521},
  {32'hc4034fef, 32'h43d2c36d, 32'hc4074517},
  {32'h44103207, 32'hc1ce0754, 32'h429bbe32},
  {32'hc5458bcd, 32'h432c959b, 32'hc453914f},
  {32'h434dfb7f, 32'hc4927de3, 32'h4410355d},
  {32'h44be4a1d, 32'h43fbcf7c, 32'h446d8726},
  {32'h43007148, 32'h43527536, 32'hc507c215},
  {32'h448180b8, 32'h436ce1a4, 32'hc19bcdb6},
  {32'hc4e52f44, 32'h438230e4, 32'h429bfb43},
  {32'hc54cba74, 32'hc3772176, 32'h433e8b47},
  {32'h44e3f6a7, 32'hc3161444, 32'h42a96138},
  {32'hc5201c70, 32'hc3040fc8, 32'h4334b076},
  {32'h44b275e3, 32'hc4770b12, 32'hc3ba8313},
  {32'hc3b958b4, 32'h4471a367, 32'hc425bb85},
  {32'hc4b77e3f, 32'hc228f97d, 32'h43c9975e},
  {32'hc59387c6, 32'hc3a90a45, 32'h4349e44c},
  {32'h44fb4f44, 32'h441ada53, 32'h44075333},
  {32'h448377e7, 32'h424522e0, 32'hc4174d9f},
  {32'h430c3954, 32'hc4ca9763, 32'hc321bc3f},
  {32'hc52713ad, 32'h435b623e, 32'h43ba8c1e},
  {32'hc376cc0c, 32'hc49754dc, 32'h4282eae4},
  {32'hc5217ce6, 32'h446bbc69, 32'hc3988fee},
  {32'h43852869, 32'hc5208e5a, 32'hc3a71daa},
  {32'hc48995eb, 32'hc44e43e9, 32'h438af059},
  {32'h4501e40f, 32'h43cb20d1, 32'hc406ceb4},
  {32'hc4d81a3d, 32'h4486bbd4, 32'h4430157c},
  {32'hc41ae19c, 32'hc23baca4, 32'h44611243},
  {32'hc3824fa2, 32'hc34badd5, 32'hc531c82e},
  {32'hc38ded84, 32'hc4720490, 32'h42870990},
  {32'hc387380a, 32'h44793fed, 32'hc3c603ad},
  {32'hc51f7a80, 32'hc306244e, 32'hc3760f57},
  {32'hc31c4ed5, 32'h430b4783, 32'hc2982ede},
  {32'hc3d62667, 32'h4490a93a, 32'hc286d426},
  {32'hc44f1979, 32'h43546354, 32'h44dae958},
  {32'h450973b6, 32'h4469b46c, 32'hc4a4db66},
  {32'h4183ce80, 32'h43535ec0, 32'hc4f057df},
  {32'hc3854cc0, 32'hc4861012, 32'h44269ce6},
  {32'h448c61cc, 32'h440c1a86, 32'hc4069611},
  {32'hc48aee3a, 32'hc4896fb5, 32'h43b52c8b},
  {32'h4403a832, 32'h43bfb192, 32'hc42e480a},
  {32'hc1c27640, 32'hc30a1b56, 32'h44056e96},
  {32'h43c23c9e, 32'h4305d9c9, 32'hc40c0852},
  {32'hc517b19c, 32'hc2d28b4e, 32'hc3715702},
  {32'hc4bf0697, 32'h436b68e8, 32'hc3a123b2},
  {32'hc51fd0a1, 32'hc3f44f77, 32'h43b125d0},
  {32'hc3c9a740, 32'h44d5619d, 32'h437f18f3},
  {32'h42f489e7, 32'hc16f7d5f, 32'h4117027c},
  {32'h431d9474, 32'h45644b7d, 32'hc39e826b},
  {32'h414627d4, 32'hc54d62ee, 32'h43932cac},
  {32'h44f477c5, 32'h441cee5d, 32'h43216db8},
  {32'hc2bbcb84, 32'hc4163764, 32'h448fb6d8},
  {32'hc4fe9f4f, 32'h43681dec, 32'hc3f0ff4e},
  {32'hc3c5e58b, 32'hc4f50c1e, 32'h44ce5793},
  {32'hc48a3051, 32'h430d7866, 32'h416865d0},
  {32'h428111de, 32'h4515065b, 32'h440de2b5},
  {32'h435bd733, 32'h4375fd8a, 32'hc4f8bf0a},
  {32'hc3600b3e, 32'hc3a1e4f2, 32'h4425fd0d},
  {32'hc4e7a867, 32'hc485e996, 32'hc4c37c19},
  {32'h43452588, 32'h43e86f63, 32'h44a66af5},
  {32'h42962296, 32'hc49598db, 32'h43a44a99},
  {32'hc423a9a4, 32'hc279910d, 32'h45050223},
  {32'hc3abab5f, 32'hc4144d91, 32'hc3d23418},
  {32'h44809e9a, 32'h442e1308, 32'h43b7819d},
  {32'h42c00605, 32'hc3a8bba7, 32'hc4ee0795},
  {32'h43ed0c34, 32'hc3004d9f, 32'h41ecbda8},
  {32'hc4978346, 32'hc3d6f108, 32'h428a2a32},
  {32'h44fd74de, 32'hc1dea134, 32'h4430d1cb},
  {32'h434b8390, 32'hc41de4f3, 32'hc48a10c9},
  {32'hc4aa14ca, 32'h4377d04b, 32'h4185ab28},
  {32'hc50746a7, 32'h4387ab76, 32'h4298d629},
  {32'h4282b332, 32'h4545c98f, 32'hc31a4f79},
  {32'hc4a303c7, 32'hc2c8260c, 32'hc404938f},
  {32'h44b3d94f, 32'h44088db5, 32'hc30059d4},
  {32'hc50bdcee, 32'hc407bed0, 32'h431c25c1},
  {32'h44fe23aa, 32'h432d7bfa, 32'h43cf699a},
  {32'hc513b804, 32'h43c11e2c, 32'h43ebc012},
  {32'h4549ccf9, 32'hc37849d6, 32'h43d09f72},
  {32'h4427995c, 32'hc52962f4, 32'hc4065948},
  {32'hc33c48c6, 32'h451186e5, 32'h4399dc68},
  {32'hc16271e8, 32'hc49cb6f7, 32'hc3d9d8e3},
  {32'hc40ecc80, 32'h44501492, 32'h4460152d},
  {32'h43bd3f93, 32'hc4d39aff, 32'h42cbf412},
  {32'h431a1e17, 32'h43f18003, 32'h45027df8},
  {32'h451bac82, 32'hc3957361, 32'hc345c625},
  {32'h4263b09a, 32'h44843bf9, 32'h44a25fc7},
  {32'h43f9f330, 32'hc3c761e3, 32'h4242c5e3},
  {32'hc4791b9e, 32'h441d7050, 32'h4255f74b},
  {32'hc31608ce, 32'h43ad61b5, 32'hc5093b56},
  {32'h43b07929, 32'hc0753938, 32'h43eae776},
  {32'h4549af20, 32'hc171952b, 32'hc1f7e75e},
  {32'hc4c24fce, 32'hc3052d06, 32'h449e8c48},
  {32'h452b7310, 32'h44510d19, 32'hc15489f8},
  {32'hc48a21e4, 32'h4302cb15, 32'h44a4b36b},
  {32'hc2e8c260, 32'hc3acadc7, 32'hc50aa603},
  {32'h43982176, 32'h449c4e32, 32'h43fa4c2b},
  {32'h44e6b1f6, 32'hc49373e7, 32'hc37f1a6b},
  {32'hc4386dde, 32'h45220acb, 32'hc2290b7f},
  {32'h45081cbe, 32'h44360840, 32'h4206cbb4},
  {32'hc4347635, 32'h45327b24, 32'hc20004b6},
  {32'h44c54f5c, 32'hc4c91754, 32'hc2a2b2dd},
  {32'hc4007949, 32'hc2e65643, 32'h442f510c},
  {32'h4401cde8, 32'h4409f17f, 32'hc3e81696},
  {32'hc4444fc8, 32'hc4080fce, 32'h43d6913d},
  {32'h4427e49e, 32'hc397b27d, 32'hc4002537},
  {32'hc456008f, 32'hc3c53132, 32'h41916f90},
  {32'hc5764d6a, 32'hc38dcd69, 32'h43c88819},
  {32'h43bcb87e, 32'hc360e496, 32'h44df5db7},
  {32'hc444d19f, 32'hc299f53e, 32'h43943780},
  {32'h4419f5b8, 32'hc4cbc597, 32'hc3eff657},
  {32'hc4989a48, 32'h423f8bba, 32'hc3e9830e},
  {32'h44a4fbbb, 32'hc313cfe9, 32'h438abed6},
  {32'hc4a37e78, 32'h44b4622c, 32'hc3d62e0c},
  {32'h44bd6446, 32'hc4ccfb55, 32'h4343fa04},
  {32'h44c27445, 32'hc2a6f732, 32'hc42a92a7},
  {32'h44af20bf, 32'h41d63f56, 32'h4339acc0},
  {32'hc5422123, 32'h43897d1c, 32'h42b53ea6},
  {32'h44c0a195, 32'hc401b5ad, 32'hc38db1db},
  {32'hc4b45f97, 32'hc2b490eb, 32'h440ec691},
  {32'h44eece0a, 32'hc38e2446, 32'hc3c1e5b2},
  {32'hc377b439, 32'h44970f84, 32'h43f07eaa},
  {32'hc3721588, 32'hc4aba7f2, 32'h417e3333},
  {32'h43c20808, 32'h450b44e8, 32'h43df27ff},
  {32'h448ace35, 32'hc4530d94, 32'h4352ab79},
  {32'hc48c667c, 32'hc3b9648d, 32'h43dbb31c},
  {32'h4430c3a0, 32'h43f9b530, 32'hc481ebe9},
  {32'h432d0da1, 32'h44508114, 32'h443b78d2},
  {32'hc364df94, 32'hc547af58, 32'hc3829a37},
  {32'hc3c45f78, 32'hc3781ff2, 32'h454628d0},
  {32'h44cd5ba7, 32'hc3f05569, 32'hc210e352},
  {32'hc140c480, 32'h4455e633, 32'h45405c6b},
  {32'hc1c83b48, 32'hc4f4e4bb, 32'hc41d88ad},
  {32'h448b32bc, 32'hc38445c0, 32'hc42394e3},
  {32'hc40f64ec, 32'hc32c181e, 32'h447ee94c},
  {32'h4523bce3, 32'h43b5bd5c, 32'h43b404ba},
  {32'hc4f926be, 32'hc4a0bccc, 32'hc24b0069},
  {32'h45475123, 32'hc2848776, 32'hc30a4c3d},
  {32'hc4f9b69e, 32'hc16f1901, 32'hc2fa3c7e},
  {32'h42c94fc0, 32'h45205fc6, 32'hc233f362},
  {32'hc54c32c1, 32'hc3fad640, 32'h44161d81},
  {32'hc339a938, 32'h44c85f3e, 32'h4339cd7c},
  {32'hc4b619f0, 32'hc44ffa64, 32'h44100e3b},
  {32'h43f5adc1, 32'h42515ec4, 32'hc1e37a0e},
  {32'hc432164c, 32'hc3120c3d, 32'h44db403c},
  {32'h44dda19e, 32'h440115fa, 32'h43836d29},
  {32'h439e6f24, 32'hc376ed0d, 32'hc286e57a},
  {32'h45054524, 32'h430917b3, 32'hc1824a5e},
  {32'hc3723a6b, 32'hc4a36772, 32'hc3c7ddb5},
  {32'h446fd622, 32'h445f995d, 32'h4416645f},
  {32'hc38b249b, 32'hc4d596e0, 32'hc3bcff2d},
  {32'h44f04404, 32'hc43d7ca6, 32'h445870d6},
  {32'hc2b10790, 32'h44644969, 32'hc4c2ad0e},
  {32'hc316a6c2, 32'hc27a98b3, 32'h42852115},
  {32'hc4486e3c, 32'hc4a7ca71, 32'hc3f56996},
  {32'h44b1f3e3, 32'h448d0b3b, 32'h43cd3615},
  {32'h447edd6a, 32'hc431b299, 32'hc2aa97ba},
  {32'hc3f36d3c, 32'h44122079, 32'h4500bdc3},
  {32'hc4176e6f, 32'hc47bef0c, 32'hc428a5d9},
  {32'h438bcb6c, 32'h45080947, 32'hc36cf8bb},
  {32'h44270e66, 32'hc3c31bbc, 32'h43a65148},
  {32'hc543f166, 32'hc0f16b90, 32'h438a23ef},
  {32'h4493ca48, 32'h448061a4, 32'h43d200f2},
  {32'hc2add7e0, 32'h434d5a8d, 32'hc2303798},
  {32'h42a4e044, 32'h454e7005, 32'h42efe950},
  {32'hc43dc042, 32'h421bc27a, 32'hc1158d35},
  {32'hc3786e1c, 32'h42d61ebe, 32'hc2bd1afd},
  {32'hc58d3707, 32'h42f47ebe, 32'h43649e96},
  {32'h44d14a22, 32'hc3edf488, 32'hc34ade2c},
  {32'hc3fcd36e, 32'hc46327e1, 32'hc3a4b207},
  {32'h442eb80d, 32'h43362c22, 32'hc49c5997},
  {32'hc3ff3f26, 32'hc4829b30, 32'h4488fcc9},
  {32'hc3a0d85c, 32'h43c8a7ee, 32'hc502d294},
  {32'hc492c960, 32'hc3c32c4b, 32'h43a69c5e},
  {32'h450f4d22, 32'h433f92c2, 32'hc287a226},
  {32'hc4648c3f, 32'h4381b311, 32'hc37e9604},
  {32'h4431a57c, 32'h43bbdb86, 32'hc49412db},
  {32'hc4bb802c, 32'hc3b6931e, 32'h4427a170},
  {32'h44b113ac, 32'h429fe356, 32'hc4286d75},
  {32'hc4db824e, 32'hc45171b6, 32'h42c046ea},
  {32'h43b9d068, 32'h442dd731, 32'hc44b59f7},
  {32'h4489a937, 32'hc3a86e16, 32'h43a4f004},
  {32'h441bbd49, 32'h44656900, 32'hc39385a4},
  {32'hc53c7111, 32'hc3ccba1e, 32'h43690645},
  {32'h454f3738, 32'h4397eeff, 32'h4243ec40},
  {32'hc46e38e4, 32'hc39f2874, 32'h44a9d5fb},
  {32'h44bdc770, 32'hc28a2f70, 32'hc43f6502},
  {32'hc39d5b67, 32'hc5500e9e, 32'h41c5fe09},
  {32'hc3a99c9f, 32'h452510f3, 32'h43c083af},
  {32'h444acf8a, 32'h43e09348, 32'h43e5a3f2},
  {32'hc3f2d2fe, 32'h44f0c6a9, 32'hc3814c73},
  {32'h45089f00, 32'hc372375a, 32'hc3c078a4},
  {32'hc4c1141c, 32'h4311384d, 32'hc40fc0f7},
  {32'h44a15d78, 32'h440d569f, 32'hc2c5e4e8},
  {32'hc4b8b57a, 32'hc2828456, 32'hc2467210},
  {32'h44b3c724, 32'hc3ac027b, 32'hc354237c},
  {32'hc3ace9bc, 32'h4406a0d6, 32'hc3928cf6},
  {32'h45047dd2, 32'h42ebc199, 32'h4399adb3},
  {32'hc4410738, 32'h434928b0, 32'hc3d30403},
  {32'h43a4666a, 32'hc4dd8870, 32'h43afd2fa},
  {32'hc5540698, 32'hc3c5faea, 32'hc33c2cc5},
  {32'h44412d39, 32'hc4549a6a, 32'h436aaba7},
  {32'h41636a40, 32'h435a26fe, 32'hc458e616},
  {32'h4480ef42, 32'hc321c0b6, 32'hc2cb5930},
  {32'h43478375, 32'hc401aca9, 32'hc4a76274},
  {32'h4497c1fe, 32'hc4a59ab9, 32'hc2852bb2},
  {32'hc207b350, 32'h45444fc8, 32'hc0a7e448},
  {32'hc4b4cad8, 32'hc36a2a20, 32'h43424fc4},
  {32'h4366c2a3, 32'h4466ba31, 32'hc4993149},
  {32'h451333b4, 32'hc392f82d, 32'h43384866},
  {32'h43c990b3, 32'h44a79169, 32'hc31644c8},
  {32'h448eebf1, 32'h4469c985, 32'h44bfdef6},
  {32'hc554c8ca, 32'h43308abb, 32'hc43babd3},
  {32'h438a06ba, 32'hc38a58c2, 32'h4508f26f},
  {32'hc470048f, 32'h445da74e, 32'hc40ca357},
  {32'hc33fc190, 32'h4433acca, 32'h44f3b66c},
  {32'h43415699, 32'hc4570954, 32'hc3f2ffd9},
  {32'hc4dfb1f5, 32'h4306180f, 32'h42ef0077},
  {32'h435c13c4, 32'hc401e31f, 32'h4556482a},
  {32'h4322fab9, 32'hc42bb1e6, 32'hc5473671},
  {32'h43994510, 32'h436b77d6, 32'h440df045},
  {32'hc4054599, 32'h42e5bd2b, 32'hc5606f5f},
  {32'h43e66fdf, 32'hc3ab34cc, 32'h44a20bcc},
  {32'hc2c94364, 32'h44e5f3db, 32'h44c1ac72},
  {32'hc3b6f884, 32'h45046a24, 32'hc50925f6},
  {32'h430af2a0, 32'h429d540e, 32'h442cab5f},
  {32'h433b23cd, 32'hc4faeead, 32'h43690c65},
  {32'hc3fffde9, 32'hc178770c, 32'hc4b0f6e6},
  {32'h44385006, 32'hc32147a1, 32'h449f5ff1},
  {32'h4372358a, 32'h435d06c9, 32'hc4d2d4f3},
  {32'h44b0bfb8, 32'hc45d78a5, 32'h4400b7d9},
  {32'h43808a86, 32'h44f1a1fb, 32'hc40dd03e},
  {32'hc4eb5d29, 32'hc34e5815, 32'h43cb0052},
  {32'hc59db27a, 32'h43941d3a, 32'h42471192},
  {32'h4513197a, 32'h43e72b0f, 32'h4479cba6},
  {32'hc46cdd04, 32'hc3a9215c, 32'hc187ce08},
  {32'h44c9b180, 32'h435a9302, 32'h438ba6e0},
  {32'hc408cda4, 32'h44ff6de0, 32'hc2f19bef},
  {32'hc473689b, 32'h430f2ada, 32'h441974eb},
  {32'hc3dd308f, 32'h456fcd43, 32'hc3ab867d},
  {32'h43b89ff0, 32'hc534b57b, 32'h43eb8f1b},
  {32'hc4456cca, 32'hc2f3d481, 32'hc261c342},
  {32'h42fdd3e4, 32'hc301b9ec, 32'hc537c208},
  {32'h42cb9916, 32'hc429f015, 32'h45328c7c},
  {32'hc346eb46, 32'hc527f36d, 32'h42fda025},
  {32'h42b89ed0, 32'h4372bd9e, 32'hc4d66ae3},
  {32'hc35bb6e1, 32'hc4e8ead8, 32'h4321ddae},
  {32'h43a869f8, 32'h4525cef4, 32'hc3b43e48},
  {32'hc4723cb0, 32'hc4687596, 32'h44e2f182},
  {32'h450e5044, 32'hc2d3a2c3, 32'hc3e64039},
  {32'h44fb9b2e, 32'h43815315, 32'h437a6353},
  {32'hc513c332, 32'hc470104c, 32'h447fd979},
  {32'h42335600, 32'h44149ce6, 32'hc4b2e0b5},
  {32'h441622d0, 32'hc3ddafdb, 32'h43ed47a8},
  {32'hc409245c, 32'hc3c61c44, 32'h44223833},
  {32'hc41b4018, 32'h44a8c1ce, 32'h435fbfaa},
  {32'hc482cf98, 32'hc411a819, 32'h441944ce},
  {32'h45449cfe, 32'h430d02ce, 32'hc345eee4},
  {32'hc4f46ef1, 32'hc3eb486e, 32'hc353b6c8},
  {32'h44c925ac, 32'h43e016e0, 32'h43437035},
  {32'hc444ee68, 32'h44010e6a, 32'h42a1ebb7},
  {32'hc4e56298, 32'h4187b296, 32'hc3334fed},
  {32'h4383b6c8, 32'hc570a368, 32'hc2cf76d0},
  {32'h4312dac6, 32'h45577c3b, 32'h43cb3f95},
  {32'h44150199, 32'hc4746787, 32'h4418bdf7},
  {32'h45517e98, 32'h4385204b, 32'h43a894b5},
  {32'h43a87c02, 32'hc5752021, 32'h41f19796},
  {32'h44e10685, 32'h43c1c946, 32'h40c06ad4},
  {32'hc3bacc02, 32'h442bd722, 32'hc266b896},
  {32'hc4c08783, 32'hc3b53077, 32'hc345fbd1},
  {32'h4429a317, 32'h44ab7a94, 32'h439e9b44},
  {32'h429231a8, 32'hc4c6a13f, 32'hc3077102},
  {32'h43918c38, 32'h44b24e95, 32'h4459744d},
  {32'hc550bd26, 32'h43d830a6, 32'hc3c1938b},
  {32'h43fb4261, 32'hc3138725, 32'h4494e7f8},
  {32'hc4b74858, 32'hc4a6b478, 32'hc48fdaf3},
  {32'h44f3a410, 32'h43b9ef22, 32'h4429fbc5},
  {32'h4396cf67, 32'hc41140cc, 32'hc382695a},
  {32'hc413e49e, 32'hc437a4f8, 32'h44aad12c},
  {32'hc2d38720, 32'h44908398, 32'hc4e830c7},
  {32'hc3a5e95e, 32'h441404b7, 32'h4499ed76},
  {32'hc35103a0, 32'hc525c943, 32'hc333b07f},
  {32'hc3314340, 32'hc3b69772, 32'h44039a33},
  {32'hc386030c, 32'hc488970b, 32'hc2bb60d2},
  {32'h44a85789, 32'h438c696a, 32'h44a64b77},
  {32'hc4cf3c85, 32'h42902e2e, 32'h42e61291},
  {32'h45364a43, 32'hc2dfef84, 32'h448cfd44},
  {32'hc57d1464, 32'h427e4b97, 32'hc2f3587a},
  {32'h444a8a9d, 32'h44978a67, 32'h42cd7975},
  {32'hc4f753da, 32'hc12533b3, 32'hc357c873},
  {32'h448bfe25, 32'h445c64ec, 32'h439b3b2e},
  {32'hc4cbc42a, 32'hc468430a, 32'hc31e4f34},
  {32'h44f7a8e4, 32'h43596b9e, 32'h4397d764},
  {32'hc59a7064, 32'h41c96a4f, 32'hc3a8edbe},
  {32'h454bf3ea, 32'h426f3054, 32'h40b467d0},
  {32'hc2da910c, 32'hc486626f, 32'hc4988c1b},
  {32'h43032626, 32'hc4bd2725, 32'h44fd2f7e},
  {32'hc393a387, 32'h43168af0, 32'hc419129c},
  {32'hc52780d2, 32'h43a05bcd, 32'h437055cc},
  {32'h4500981e, 32'hc3428882, 32'hc44d2d21},
  {32'hc2826380, 32'h43de2e84, 32'h44247601},
  {32'hc3b8edbf, 32'hc4d843df, 32'hc4d890dc},
  {32'hc4025dc9, 32'h442b4a5c, 32'h450a35c2},
  {32'h4495de98, 32'hc42b19ff, 32'hc31a69bc},
  {32'h43a52908, 32'h44bcf82d, 32'h446fb287},
  {32'hc2183a7c, 32'h4420570d, 32'hc49ab71e},
  {32'hc310c584, 32'h43a40244, 32'h4409716a},
  {32'h437961f6, 32'hc3ce7951, 32'hc198297a},
  {32'hc5135ce7, 32'h43bb0a91, 32'h4312a611},
  {32'hc49e9193, 32'hc38207b4, 32'hc390d311},
  {32'hc435968d, 32'h438e74ee, 32'h4512eab7},
  {32'hc3955ce4, 32'hc5104e90, 32'hc4ec119d},
  {32'hc2ac68ba, 32'h42a757c8, 32'h44ed8dab},
  {32'h4344ccb0, 32'hc49bb9f9, 32'hc4698024},
  {32'hc4d54311, 32'h44896ecc, 32'h43aa0fe7},
  {32'h4541a05f, 32'h41f408c2, 32'hc3051054},
  {32'hc2abf620, 32'h4563d921, 32'hc31698ec},
  {32'h445d2e7a, 32'hc52a7659, 32'h441230c3},
  {32'h43856fc0, 32'h4405c2ff, 32'h430b6676},
  {32'h4563b2d6, 32'h439a9dcf, 32'h43f26b62},
  {32'hc5491bf5, 32'h4397e390, 32'h44094b98},
  {32'h43e0500f, 32'hc377614c, 32'hc3893fe6},
  {32'hc3e3df89, 32'h437800f2, 32'hc398f194},
  {32'hc4803d9a, 32'hc39ccf92, 32'hc508a1a1},
  {32'h44ca9930, 32'h43a27e89, 32'h44578c91},
  {32'h4257c2de, 32'h44532ded, 32'h42de809b},
  {32'h44aaefa6, 32'hc41e67ee, 32'h4102dd16},
  {32'hc33c2e82, 32'h450f5bf7, 32'h4321a36f},
  {32'h451ef579, 32'h43667f2a, 32'hc36c16a0},
  {32'hc385b068, 32'h455b8708, 32'hc366c2e9},
  {32'h43331d50, 32'hc54ff192, 32'hc336c23a},
  {32'h44f59f4a, 32'hc1bc5dcb, 32'hc4108845},
  {32'h4406ece0, 32'hc45e5e71, 32'hc4009f88},
  {32'hc3479088, 32'h447296d0, 32'h447b08f8},
  {32'hc424e8ca, 32'hc40989b1, 32'hc37fe311},
  {32'hc4cb8a80, 32'h443674de, 32'h43687832},
  {32'h4471caa4, 32'hc3c42135, 32'hc3ce6153},
  {32'hc15e51db, 32'h4392330a, 32'h44f46dc6},
  {32'hc3675e48, 32'hc3254432, 32'hc48236a8},
  {32'hc35eeab8, 32'h44345bf8, 32'h44c4cb5b},
  {32'hc4e69fd1, 32'hc3c6ec91, 32'hc2ba3d77},
  {32'hc5658b7e, 32'h43d2ed03, 32'h43684b41},
  {32'h4553c559, 32'h438fa82b, 32'hc3be8b6c},
  {32'h44e893fd, 32'h4393a5ad, 32'h43a38d45},
  {32'h438f3168, 32'hc4d8d653, 32'hc3eef551},
  {32'hc3b03d0a, 32'h44e7a786, 32'h44eeab4a},
  {32'h451f60e4, 32'hc34b1a6c, 32'hc21ca1b7},
  {32'hc568097c, 32'h44543939, 32'h43237ca4},
  {32'hc268403a, 32'hc56a7e6a, 32'hc2780f50},
  {32'h44b9302f, 32'hc154eb29, 32'hc4c53619},
  {32'hc5552f9f, 32'hc401c12d, 32'h42ae2de6},
  {32'h4466ea02, 32'h42f40024, 32'hc3099753},
  {32'hc3dc8030, 32'hc441b639, 32'h43dbf8d7},
  {32'h450bd047, 32'h406fab4d, 32'h42d46725},
  {32'h43d5994a, 32'hc3aab939, 32'hc2942fc2},
  {32'h4530af6b, 32'h449271df, 32'hc31254b6},
  {32'hc3e74a0c, 32'hc509f710, 32'hc429d8c5},
  {32'hc46286c9, 32'hc37610f1, 32'h445d4eb6},
  {32'hc49d982b, 32'h4193142c, 32'hc32d6406},
  {32'h43870ec7, 32'h4465529a, 32'h447a40dd},
  {32'h44d07608, 32'h43d7eb47, 32'hc2af5458},
  {32'h44440204, 32'h443acce0, 32'h43a98cbf},
  {32'hc392e510, 32'hc480e679, 32'hc436b947},
  {32'h44bf55c2, 32'h4330935c, 32'h426a0dd2},
  {32'hc346b9a8, 32'hc480d4f7, 32'hc4baea9b},
  {32'h42661432, 32'h450cd8e3, 32'hc34dbaf2},
  {32'hc4174241, 32'hc41061af, 32'hc4984511},
  {32'h4415a150, 32'h4445081e, 32'h44bc8aef},
  {32'hc3bac408, 32'hc34ea1b0, 32'hc426ab35},
  {32'h447f6e0e, 32'hc29da4ef, 32'h43394719},
  {32'hc46b7ffc, 32'hc38c5af4, 32'hc4a3d35b},
  {32'h4471fc88, 32'h43107482, 32'h440ca138},
  {32'hc529f14d, 32'hc31ca711, 32'h43e6c3bd},
  {32'h439963c0, 32'h4462d9df, 32'h44a90ec3},
  {32'h43b8c488, 32'hc55d9cf0, 32'hc31d3163},
  {32'h44cb7001, 32'hc33ce041, 32'hc3098bf5},
  {32'hc4d76d00, 32'h42c2e162, 32'hc3efbd1c},
  {32'hc43e4c8e, 32'hc4d48773, 32'h43154f42},
  {32'h432fb320, 32'h44e69d33, 32'h445f1c54},
  {32'h44a70184, 32'hc3dc1c63, 32'h438a8c99},
  {32'hc374f7ce, 32'h456bebee, 32'hc3508448},
  {32'hc1e16c80, 32'hc51d2c00, 32'hc2c6c63f},
  {32'h4417a81b, 32'h43cb1d23, 32'hc382f82d},
  {32'hc57aa356, 32'h43cd7f7e, 32'hc3e2f763},
  {32'h438c6e70, 32'hc34b1349, 32'h4399ecae},
  {32'hc3d48d64, 32'hc311957f, 32'hc2fe64d7},
  {32'h440d50c5, 32'h447dd593, 32'hc4b499dc},
  {32'hc4f61661, 32'hc3fda169, 32'h42e49e31},
  {32'h44485391, 32'h41603457, 32'hc3325691},
  {32'hc374f5fc, 32'hc1f49364, 32'h451f683a},
  {32'h449a6662, 32'hc2a0b20a, 32'hc40afbb1},
  {32'h44893615, 32'hc2d5ed86, 32'h44225864},
  {32'h449a69b8, 32'h44412bc6, 32'hc3c00f94},
  {32'hc32bfb90, 32'hc48532c0, 32'hc1e97e8a},
  {32'hc2b72fb9, 32'h44f7ba96, 32'h427ea92a},
  {32'hc4bff975, 32'hc4804956, 32'h4507785f},
  {32'h446698a7, 32'h4486becf, 32'hc314bceb},
  {32'hc4c6e696, 32'h44108d43, 32'hc3a0f5b6},
  {32'hc38af43f, 32'h4524efaf, 32'h430c2171},
  {32'hc4720456, 32'hc1ac6f57, 32'h430db6ab},
  {32'h44e70648, 32'hc09357ec, 32'hc3346899},
  {32'hc46bca51, 32'hc1b1b451, 32'h4431169f},
  {32'h432cf5b8, 32'hc2062dae, 32'hc524599c},
  {32'h43831638, 32'h412ce138, 32'hc492f5a7},
  {32'h434eadcd, 32'h4557ff8d, 32'h43c7b9c1},
  {32'h451414ff, 32'h43e38519, 32'h43949d9f},
  {32'hc5219434, 32'h41b14660, 32'hc2bc6aee},
  {32'hc3f4319c, 32'hc5610a45, 32'h43a19f09},
  {32'h444a3f57, 32'h44c06e9b, 32'h418f2ae3},
  {32'h442f1290, 32'hc3ee9603, 32'hc4303cc9},
  {32'hc510479e, 32'hc2b1dff4, 32'hc3f50648},
  {32'h4510fbf9, 32'h43c94067, 32'h4380af77},
  {32'h43795c68, 32'h44bb988d, 32'h43a67ea8},
  {32'hc3432b48, 32'hc48e774d, 32'hc4984acc},
  {32'hc3d488a4, 32'hc3ab9324, 32'h43d2160c},
  {32'h44c0048f, 32'hc35a111e, 32'h447f8e7e},
  {32'hc3b9e7ae, 32'h44c94f4a, 32'h42cd7ab5},
  {32'hc336b6e9, 32'h43578aa4, 32'h45228e54},
  {32'hc45617a8, 32'hc0e05790, 32'hc4acbcdc},
  {32'hbaf40000, 32'h4412250a, 32'h455dfde6},
  {32'hc403ae14, 32'h43ea5c57, 32'hc229a412},
  {32'h45245d78, 32'hc4071ab1, 32'hc31d6fba},
  {32'hc40def3b, 32'h449c0696, 32'hc366d2c3},
  {32'h4506dfbf, 32'hc1e09a88, 32'hc2d19db9},
  {32'hc48c8c2c, 32'h44e791b4, 32'hc11bfb26},
  {32'hc38746fd, 32'hc48c1476, 32'h44b3dbda},
  {32'h44eb25b6, 32'hc323678b, 32'hc2c61a80},
  {32'h445e20f9, 32'h449292af, 32'h44b2b54a},
  {32'hc3c11d49, 32'hc28dc7b5, 32'hc52c7495},
  {32'hc33c7c2e, 32'hc22ffd93, 32'hc3e957e8},
  {32'hc4ce3040, 32'h4223c379, 32'hc3dbe138},
  {32'h4417996a, 32'hc458dec3, 32'h4504ffb8},
  {32'h4440a546, 32'hc2174567, 32'hc404a0e1},
  {32'hc4895280, 32'hc34869c2, 32'hc2b237ea},
  {32'h44935ef2, 32'hc48ec1e5, 32'hc3330069},
  {32'hc43d2034, 32'h44a89102, 32'hc3658c48},
  {32'h4483b960, 32'hc39df695, 32'hc35743f2},
  {32'hc43bb9a7, 32'h439571de, 32'hc542b798},
  {32'h4454ec4d, 32'h42471189, 32'h44945a66},
  {32'h42f6d558, 32'hc222e276, 32'h4507f387},
  {32'h3f0bd000, 32'h4460a484, 32'hc50af5e5},
  {32'h450b4b20, 32'h43dc4e4f, 32'hc2c42eb7},
  {32'h4446b829, 32'hc435bd46, 32'h446ddeb0},
  {32'hc40bc85c, 32'h448514fc, 32'hc3a7ce9b},
  {32'h447cfa48, 32'hc4bf89b1, 32'hc3f0d937},
  {32'h4330f208, 32'hc35c7e57, 32'hc3993d40},
  {32'h4400685a, 32'hc4d2f841, 32'h43eb8ab3},
  {32'h41725c08, 32'hc3a1d7d1, 32'hc50383b8},
  {32'h44a4f0ba, 32'hc4187113, 32'h42a9a723},
  {32'hc4c94c42, 32'h435597d4, 32'hc4274f4e},
  {32'h444a002a, 32'hc089ba84, 32'hc3deb788},
  {32'hc3be775c, 32'h43cb5735, 32'h43cccb24},
  {32'h44b093de, 32'hc48fc20c, 32'hc23203c5},
  {32'hc2f627e2, 32'h450aedbc, 32'h43ea79ec},
  {32'h44e35c99, 32'h440e6983, 32'h433d94d5},
  {32'hc4533cf6, 32'h44c89b56, 32'hc3fce949},
  {32'h455c5700, 32'hc4349a98, 32'hc31ac3b3},
  {32'h4410ecb8, 32'hc40cc69d, 32'h44b4c8a8},
  {32'hc2ed3e00, 32'h450b9284, 32'hc49eb5a3},
  {32'hc2e89223, 32'h443ae7cb, 32'h4490a77d},
  {32'hc433810d, 32'hc3cb5bf2, 32'h41a63d6d},
  {32'h44f35734, 32'h423c1ebe, 32'h43ab3068},
  {32'hc3f53a3e, 32'hc4432781, 32'h423f2644},
  {32'h4450c797, 32'h44231d7f, 32'hc46c30cc},
  {32'hc426d49b, 32'hc53394a0, 32'hc2d6aaca},
  {32'h4347aa82, 32'h44ad6922, 32'h43f0d309},
  {32'h452d4a8a, 32'h438be204, 32'h442009c4},
  {32'h43928b2e, 32'hc482d39e, 32'h44f748df},
  {32'h452f5470, 32'hc34dfe11, 32'hc43741a2},
  {32'h43575dc6, 32'h413577ce, 32'hc511f33f},
  {32'hc4228d0b, 32'hc45a53dc, 32'h435277d6},
  {32'hc48302ef, 32'h410aa5f4, 32'hc3caf729},
  {32'hc50b3fcf, 32'hc45023f7, 32'h43b4a318},
  {32'h43e8eedc, 32'h432e4fb6, 32'hc4687a91},
  {32'hc5040274, 32'hc38a49a6, 32'hc2047a65},
  {32'h43ac81c0, 32'h4418703b, 32'hc4208fdf},
  {32'hc56d0a7c, 32'hc3eae88f, 32'h444d77f4},
  {32'h4583aa24, 32'h4382828f, 32'hc262365b},
  {32'hc27fdc26, 32'hc5884c2c, 32'h43927f7d},
  {32'h44069fa0, 32'hc2c8f9cc, 32'hc3dd6ca0},
  {32'h43a1d811, 32'hc3851866, 32'hc345bcef},
  {32'h44e79200, 32'h446782b6, 32'hc3e04446},
  {32'hc534da9c, 32'hc42791fb, 32'h42d553b2},
  {32'hc504ccbd, 32'h42e92728, 32'hc393acde},
  {32'h4489126f, 32'hc3431d93, 32'h41acbc2b},
  {32'hc2a4bef4, 32'hc3364e1c, 32'hc3c63103},
  {32'h444e85df, 32'h44a047ab, 32'h44276af8},
  {32'h434ab163, 32'hc2a45511, 32'hc3f93676},
  {32'h450121fd, 32'h44886b88, 32'h438a9803},
  {32'hc49753f1, 32'hc384c93e, 32'hc4812275},
  {32'h44396e8e, 32'h4321699b, 32'hc38e4e73},
  {32'hc45574c8, 32'hc4845ba5, 32'hc4e29366},
  {32'h44441a48, 32'h4413f3dc, 32'h44d2cf00},
  {32'hc3b5a51f, 32'h43207264, 32'h437642c6},
  {32'hc434e5cd, 32'hc292ae72, 32'h43ece2a7},
  {32'hc42d3c0c, 32'hc4899a07, 32'hc4194e7d},
  {32'h43fc04a4, 32'h44b3857d, 32'h43c45ff7},
  {32'hc3c8751d, 32'hc3c007b7, 32'hc4f8487e},
  {32'h43fe631b, 32'h451a3fcb, 32'h443f7f68},
  {32'h44f9cb40, 32'h421f3e70, 32'h4359cca3},
  {32'hc4179163, 32'h44d0c1a5, 32'h45150d0d},
  {32'hc519a179, 32'hc37874a9, 32'hc2fd7810},
  {32'hc3828bb8, 32'h44b2d77a, 32'hc17d813c},
  {32'hc23e8680, 32'hc5750335, 32'h42fdcab8},
  {32'h44529f65, 32'h451c66ea, 32'h43f3c374},
  {32'hc54a59f0, 32'hc3bdfc5f, 32'hc2fda8f6},
  {32'h44c89858, 32'h42bbfa97, 32'hc374455b},
  {32'hc5166237, 32'hc382fbae, 32'hc31a0ed7},
  {32'h446bdb6e, 32'h43f4f330, 32'h43afc395},
  {32'hc550ee2b, 32'hc34b95b7, 32'hc383dce8},
  {32'h44aea814, 32'hc34cd9b0, 32'hc3f274ea},
  {32'h43fb484c, 32'h434404c1, 32'hc42cc65a},
  {32'h43828e2d, 32'hc421c90f, 32'h44e737db},
  {32'hc43698a0, 32'h4433b01e, 32'hc49ad096},
  {32'hc31f7293, 32'h4439bf27, 32'h412dea22},
  {32'hc32b659a, 32'h411051b9, 32'hc52ec3e8},
  {32'h43152b2a, 32'h44a4369f, 32'h43d44ed0},
  {32'h44d573d3, 32'h43d70364, 32'hc460bb48},
  {32'hc51d17e4, 32'hc24a34e8, 32'h43d4d438},
  {32'hc3430e68, 32'hc1114d3a, 32'hc4399443},
  {32'h436ac81c, 32'h434b6b8b, 32'h44a40c33},
  {32'h412be830, 32'h450f9049, 32'hc4d283e3},
  {32'h4360e2e3, 32'h45172d55, 32'h40aad228},
  {32'hc23ec950, 32'hc4be3951, 32'hc3993119},
  {32'hc49e36a4, 32'h449527ec, 32'h43bb561a},
  {32'h431984f7, 32'h43d3e873, 32'hc4dd17d1},
  {32'hc3eb0f50, 32'h44f87910, 32'h44d029af},
  {32'h441c723d, 32'hc4ac3e25, 32'hc41d95d7},
  {32'hc39b5a85, 32'hc3eb7b92, 32'h44c22679},
  {32'h449cb6dd, 32'hc487b955, 32'h4337b326},
  {32'hc3db8c47, 32'h45492fbd, 32'h432f5291},
  {32'h43429de1, 32'hc4a1805e, 32'h43ac7d4a},
  {32'hc500a978, 32'h449e56fe, 32'hc3275300},
  {32'h44d98b49, 32'hc4211ec4, 32'h44052e73},
  {32'hc41d80bf, 32'h44465ca5, 32'h42b03655},
  {32'h444866c8, 32'hc3d2360c, 32'hc32f1af0},
  {32'hc596ced3, 32'hc3e38b16, 32'hc3a8b114},
  {32'h4549b5f3, 32'hc39f82ab, 32'h4399779f},
  {32'hc4a9b31f, 32'h42985615, 32'h43fc42f2},
  {32'hc55b9058, 32'hc3bc5af3, 32'h42109c7b},
  {32'h4422ba14, 32'h43df1dc8, 32'hc30c8aba},
  {32'h448daef8, 32'h43f32ea2, 32'h433e055e},
  {32'h420c4e00, 32'hc5072e41, 32'hc28681f7},
  {32'hc4a77b9d, 32'h448765d5, 32'h42dfc97a},
  {32'h40b2ba20, 32'hc4d7486c, 32'h43ae27bb},
  {32'hc4ce28db, 32'h44ae426b, 32'h42cb2bae},
  {32'h4391d14e, 32'hc507f59f, 32'hc3ef780d},
  {32'hc4ad38c4, 32'hc41846ad, 32'h436308fb},
  {32'h44533e42, 32'hc22131aa, 32'hc40570f0},
  {32'h42d45520, 32'hc09c640a, 32'hc4c64cc9},
  {32'hc3fe68c1, 32'h439ffb72, 32'hc430a6b8},
  {32'h44331c55, 32'h43a85266, 32'h4518fc2b},
  {32'h44e0038d, 32'h413a0e6c, 32'hc401f8cc},
  {32'h44883558, 32'h42b7b915, 32'h43c48a8b},
  {32'hc36607c8, 32'hc48c3c82, 32'hc416133d},
  {32'hc42b8ef3, 32'h4405a722, 32'h441351f5},
  {32'h44706566, 32'hc3d43418, 32'hc3932e56},
  {32'hc58d5941, 32'h42cc052c, 32'hc259a614},
  {32'h45284c33, 32'h440a0c44, 32'hc44b649b},
  {32'h441cf641, 32'h43fd5e8c, 32'h43bad960},
  {32'h453c02a9, 32'h439835ca, 32'hc3c672ff},
  {32'h421f1ef0, 32'h451479c8, 32'hc1b26867},
  {32'h42c43adc, 32'hc0805d40, 32'hc4f5e0e4},
  {32'hc392be80, 32'h448c4c0c, 32'h44ab06d3},
  {32'h447196da, 32'hc452ad56, 32'hc476309c},
  {32'hc39d204a, 32'h42c61eb2, 32'hc4c05aac},
  {32'hc54b5324, 32'hc0b76bc8, 32'h433c5b69},
  {32'h44fcbf52, 32'h441017bd, 32'h44128423},
  {32'hc49c3d01, 32'hc4b8f1f3, 32'hc4321fa4},
  {32'h44c8f63d, 32'h43ef3d45, 32'hc3d026b7},
  {32'hc41abdb4, 32'h439e74d8, 32'hc35beefc},
  {32'h44efc476, 32'h44c3cac1, 32'h43d0c684},
  {32'hc52f55ba, 32'hc3fd1abf, 32'h44110678},
  {32'h443459eb, 32'hc3afacb9, 32'hc305ae56},
  {32'hc45d31f3, 32'h420cd6f7, 32'h4511e28a},
  {32'h44f1c60c, 32'h429a7c2e, 32'hc487fd49},
  {32'h42a2535c, 32'h42d8101c, 32'hc3a549dd},
  {32'h43054c00, 32'hc0919119, 32'h44d88297},
  {32'h429fe1d0, 32'hc4293115, 32'hc4043f2b},
  {32'hc314b336, 32'h44e5c81e, 32'h42ebc3e6},
  {32'hc4feb6b1, 32'hc318757c, 32'h431dedea},
  {32'h43e8e618, 32'h444d280c, 32'h446c7f67},
  {32'hc48cbdbb, 32'hc486ef85, 32'hc3a3bcc2},
  {32'h449e0dd4, 32'hc29433a3, 32'h44ac7ade},
  {32'hc40dd926, 32'hc4261784, 32'hc4bf99ca},
  {32'h43f45782, 32'hc38c1708, 32'hc21f91fe},
  {32'hc49e2587, 32'hc4c18cd2, 32'hc32366cb},
  {32'h43d04f1a, 32'h4528f2be, 32'h4398aedd},
  {32'hc3d0fe67, 32'hc401b051, 32'hc41aa1d5},
  {32'h450b3ebf, 32'h43f76cee, 32'h4339d1ff},
  {32'hc4c27a91, 32'hc453294e, 32'hc40efabd},
  {32'h433bd550, 32'h43480640, 32'h444ea30b},
  {32'h4427e105, 32'h4405a9ff, 32'h42cd6fc5},
  {32'hc536a2a5, 32'hc385d272, 32'hc30051db},
  {32'h438e1b4c, 32'hc3b7fb99, 32'h450af0b5},
  {32'h4493af09, 32'hc4025cd7, 32'hc34e2a7d},
  {32'h42b43878, 32'h452d73ca, 32'h42d93d37},
  {32'hc381ac22, 32'hc567c0fc, 32'h42d9376b},
  {32'h45532d1c, 32'h42a181e6, 32'hc28a5d04},
  {32'hc4f8ae0b, 32'h41cfb33f, 32'h42d62710},
  {32'h44f3df48, 32'hc4485d87, 32'h42e04ce9},
  {32'hc50eb9f2, 32'h4407d741, 32'h4448b387},
  {32'h445d6d00, 32'h41cb0f34, 32'h443d0a8b},
  {32'hc45be7d8, 32'hc44887d2, 32'h44c34bea},
  {32'hc368875e, 32'h4326a36c, 32'hc491ab35},
  {32'hc401b2f8, 32'hc4e19344, 32'h431b8f8a},
  {32'h43986e07, 32'h43066523, 32'hc4540f9b},
  {32'h449d1a64, 32'h4215a5c0, 32'h43a77d72},
  {32'h441540a5, 32'hc2c833b2, 32'hc5039e50},
  {32'hc481b120, 32'hc391ff01, 32'h4413b571},
  {32'h441f047a, 32'h43bef829, 32'h42a7e1a1},
  {32'hc446f026, 32'hc4c592ba, 32'h441fa538},
  {32'h44602b22, 32'h451d5d1f, 32'hc3834ac5},
  {32'h44929f14, 32'hc2a7c40b, 32'h4412e1e5},
  {32'h441069e2, 32'h43a2acb7, 32'hc490be23},
  {32'hc49d35b2, 32'h4368276f, 32'h443808e4},
  {32'h4493b29f, 32'h43db1c80, 32'hc3704256},
  {32'hc4cedbaf, 32'h434a2cf8, 32'h4459f99a},
  {32'h44dbc3ec, 32'h42859f4a, 32'hc434f0f3},
  {32'h44e7d017, 32'hc4752d50, 32'h42afd28e},
  {32'hc54b04ec, 32'h41724feb, 32'h442f2597},
  {32'hc4adddc2, 32'h431ab45f, 32'hc2acbb3d},
  {32'hc2e7f7c0, 32'h44c9ec93, 32'h41d78397},
  {32'h44921e60, 32'hc475ac44, 32'h438618e2},
  {32'hc4a507f6, 32'h43c1bfd5, 32'hc28a269f},
  {32'h44eb5e86, 32'hc396c2ed, 32'hc44fedbd},
  {32'hc53d0420, 32'h43cbfcdc, 32'h4254f207},
  {32'hc4a3f700, 32'h432571d2, 32'h43745875},
  {32'h42435190, 32'h4513dc40, 32'h428da358},
  {32'h4525d44c, 32'h432af121, 32'hc3662b4c},
  {32'hc22f4120, 32'h44a3d54c, 32'h43d4cd53},
  {32'hc39a3091, 32'hc4d45f94, 32'h441d0961},
  {32'hc3bf8af6, 32'h4353bf49, 32'hc5475137},
  {32'h43c9d838, 32'hc41b7280, 32'h43cedaf3},
  {32'hc4572da4, 32'hc359f8fd, 32'hc4e40bbe},
  {32'h43e4b193, 32'hc2bcd6ce, 32'h4408c156},
  {32'h43f714f6, 32'h438dc06a, 32'hc43f2e19},
  {32'h44a6c57f, 32'hc4b58586, 32'hc3bf07a3},
  {32'hc4225ab2, 32'h44073b82, 32'hc4bb38c2},
  {32'h44b23d36, 32'hc3e42216, 32'hc326c7d4},
  {32'h4268f77a, 32'h44a79d2f, 32'hc48b27fe},
  {32'h445cd14c, 32'hc42ac331, 32'h441e44f1},
  {32'h43a804eb, 32'h450b6adc, 32'hc3eb4e19},
  {32'h44d132ca, 32'h42e15247, 32'h449c19d6},
  {32'hc585bf79, 32'h4337e476, 32'h43b3fcdf},
  {32'h44e2de05, 32'h42764bac, 32'h425bd461},
  {32'hc41b15b4, 32'hc48b4566, 32'hc4cb5b5d},
  {32'hc35ec22c, 32'hc4621e4e, 32'h44f6ccb8},
  {32'h4370e38e, 32'h449b7ce4, 32'hc4c8cf4b},
  {32'h448cfe33, 32'h43088018, 32'h439a86cf},
  {32'h43e15944, 32'hc28341a8, 32'h439ed219},
  {32'h426e0edc, 32'h44f3074e, 32'hc2288e77},
  {32'hc3b101f4, 32'hc380cd37, 32'h42887004},
  {32'hc517e3c4, 32'h43841f87, 32'hc250b800},
  {32'h452b7f18, 32'hc2fd71fc, 32'h43c2591a},
  {32'h440a1f34, 32'h44aab0d0, 32'h447f1d54},
  {32'h43773598, 32'hc485c7d8, 32'hc5332737},
  {32'hc413f472, 32'hc2ab37e1, 32'h42602a04},
  {32'h4424305d, 32'hc2cfbb0a, 32'h43871c3d},
  {32'h438af78d, 32'h451c6766, 32'h426327ee},
  {32'h43fd5b94, 32'hc41b868c, 32'hc3d1f15d},
  {32'hc50b649a, 32'h43a81482, 32'h4410a4f4},
  {32'h44a32aab, 32'hc2a37d88, 32'h4486db6b},
  {32'hc45b44b6, 32'h448dea3a, 32'hc3fcb5de},
  {32'h455ceec2, 32'hc3c371db, 32'hc19134f5},
  {32'hc480d309, 32'hc17763a6, 32'h4419d30a},
  {32'h453ec981, 32'h4353f883, 32'h441f880b},
  {32'h442d1b00, 32'hc3a233d4, 32'hc0a66235},
  {32'h4495c46a, 32'hc47437ea, 32'hc427eda8},
  {32'hc38223a7, 32'h445984c8, 32'hc3134074},
  {32'hc4dce109, 32'h412a4ba8, 32'hc237e9ae},
  {32'hc3c1f4e8, 32'h4556a731, 32'hc3bb9240},
  {32'h4488ad19, 32'hc4b64547, 32'h428e24cb},
  {32'h43da45a8, 32'h448d3d41, 32'hc30c90cb},
  {32'h4475893e, 32'h435504a9, 32'hc463f083},
  {32'hc3d5bb11, 32'h44dd5e93, 32'h44ba3882},
  {32'hc1cd156a, 32'hc4cb42b7, 32'h433f96ee},
  {32'h43d88e88, 32'h45245d0b, 32'hc2aa6f04},
  {32'hc3b56638, 32'hc4988f08, 32'hc38ea135},
  {32'h4374b4f8, 32'h42fe714c, 32'hc4fc9964},
  {32'hc3c24ad5, 32'hc40d0294, 32'h440c8a2a},
  {32'h440e2b3e, 32'h4440af1d, 32'h43bc30ea},
  {32'h43f9594e, 32'hc418bdb5, 32'h434733cb},
  {32'hc428a68a, 32'h44f66d6f, 32'h44bf7b63},
  {32'hc3d5b670, 32'hc4d49048, 32'hc4d9caea},
  {32'h436c1b40, 32'h44159317, 32'hc421c7d0},
  {32'hc3bb0823, 32'hc1428682, 32'h450c2c5c},
  {32'hc3370f07, 32'h43327f33, 32'hc2b8fd15},
  {32'hc3e8801c, 32'hc51bbb7c, 32'hc3ad5ac6},
  {32'hc2b56abe, 32'h45336b7e, 32'hc22e43ce},
  {32'hc1e69f1e, 32'hc40c5fa4, 32'h432910ec},
  {32'h451e77e2, 32'h430115fe, 32'hc28e916e},
  {32'hc4642118, 32'hc3284ac6, 32'h440af228},
  {32'hc46df8de, 32'hc3a1bf3d, 32'hc37deaea},
  {32'h428240f0, 32'hc52ceb4c, 32'hc34502e2},
  {32'h453062a3, 32'h43d84e8e, 32'h44039a7e},
  {32'hc280d390, 32'hc4d55e1b, 32'h43e70381},
  {32'h4556871f, 32'h440a2335, 32'hc3347418},
  {32'hc4b58bc5, 32'hc49f9a9f, 32'h440e3876},
  {32'hc4449d6c, 32'h44241a80, 32'hc3e7f065},
  {32'hc4192c84, 32'hc248f3d7, 32'h438e5aba},
  {32'hc3c50cd4, 32'h44d84c54, 32'hc48e9bb2},
  {32'h448e48d4, 32'hc384d6af, 32'h448215e2},
  {32'hc40a2d7e, 32'h436f5a02, 32'hc2cfa3d0},
  {32'h41a95a11, 32'h432a7b46, 32'hc3331f6b},
  {32'h434e75a5, 32'hc4cd0fd9, 32'hc344b906},
  {32'hc2998c5c, 32'h43849c02, 32'h437f1950},
  {32'hc4969622, 32'h43d4dda1, 32'hc49efc21},
  {32'h4402b0a0, 32'h4383e2bc, 32'h44fa4320},
  {32'h438302e3, 32'h43716007, 32'hc4937944},
  {32'hc409d9da, 32'hc4eb5aa1, 32'h4504b124},
  {32'h43c270b9, 32'h448bf9fa, 32'hc49cc338},
  {32'hc3ab2a4a, 32'h43c88800, 32'h443f4917},
  {32'hc2023278, 32'hc3814649, 32'hc5193ef0},
  {32'h4481cf1a, 32'h43a232b9, 32'h448817f1},
  {32'hc4e4d374, 32'hc38be86d, 32'h438d3a60},
  {32'h43760048, 32'h448ba767, 32'h442739f5},
  {32'hc2c98946, 32'hc494d852, 32'hc49b430e},
  {32'hc3bf629e, 32'h447dfaee, 32'h43cbce6f},
  {32'hc4165e0f, 32'hc5019375, 32'hc46aadc2},
  {32'h4314db70, 32'h44f5ff35, 32'hc2067f7a},
  {32'h448bf2a1, 32'hc418bf61, 32'hc3bad4a9},
  {32'h44085e76, 32'h44be07c5, 32'hc3cb4252},
  {32'hc47803d4, 32'hc4c1690f, 32'hc3de3445},
  {32'h456970a4, 32'h439e54ad, 32'h4451c867},
  {32'hc4b1eed4, 32'hc30bd1f2, 32'h43a3b2c7},
  {32'h44a5b71c, 32'h433cca1e, 32'hc39293ff},
  {32'h43e9c5ab, 32'hc4bddfb9, 32'h43273709},
  {32'h433289f2, 32'hc1edfa5c, 32'h4498aab2},
  {32'h4390db63, 32'h44aee9f0, 32'hc3e98896},
  {32'hc3b24050, 32'h4378daab, 32'h4402b8bf},
  {32'hc204e5d2, 32'hc4c3d861, 32'hc49db75a},
  {32'hc23e1bce, 32'h4350ed87, 32'h451dded2},
  {32'h4504449c, 32'hc34714d8, 32'hc40ace8e},
  {32'hc4c0ce50, 32'h4440e91c, 32'h40a0adf0},
  {32'hc387d7dd, 32'hc44ad742, 32'hc4b46f6c},
  {32'h44b389f2, 32'hc49fdbe6, 32'h450bec3f},
  {32'hc31e8b14, 32'h450d4482, 32'hc5150225},
  {32'h4418c1dc, 32'h410611cc, 32'h439cd44c},
  {32'h435e405f, 32'hc4982784, 32'hc493c1a8},
  {32'hc4f94ed4, 32'h443a4a6c, 32'hc328e92a},
  {32'hc4215a4f, 32'hc3d6024a, 32'hc42949d2},
  {32'hc3c9935e, 32'h44953849, 32'h44a2646b},
  {32'h453ed5ca, 32'hc2f064dc, 32'h422a7752},
  {32'h4425bde2, 32'h444c96a6, 32'h444de15e},
  {32'h448e57b6, 32'hc4a352e5, 32'hc02804c4},
  {32'hc54085e8, 32'h43f83dc5, 32'hc36304d8},
  {32'hc2eb7180, 32'hc4c3f3a7, 32'h43830c27},
  {32'hc50893df, 32'hc1554433, 32'hc36b1cc7},
  {32'h43c639d8, 32'hc46c08f4, 32'h439055b5},
  {32'h44d201ef, 32'h43b3360c, 32'hc33cdd64},
  {32'h4503b143, 32'hc33fd9da, 32'hc2d660f7},
  {32'hc565b00c, 32'hc3b81c2d, 32'hc30fa8fd},
  {32'h45350f73, 32'hc3e20b72, 32'h426d23e5},
  {32'h4532b667, 32'hc35354b4, 32'hc38ae8e5},
  {32'hc5085d5a, 32'h430f7dfc, 32'hc3a44baf},
  {32'h445bb14a, 32'hc34d5d24, 32'h44ee29c2},
  {32'hc436aacc, 32'h445d5a33, 32'hc2e0fa19},
  {32'h42a5fb60, 32'hc547f78a, 32'hc38f0c0a},
  {32'hc4a6efb5, 32'h44b40f9f, 32'h422f48e1},
  {32'hc276ac38, 32'hc4bc41ae, 32'h430b3659},
  {32'hc52dcbbf, 32'h43868dd2, 32'h4388d89f},
  {32'hc26ff456, 32'hc54eeddb, 32'hc267c7be},
  {32'h44da0488, 32'hc2d982ea, 32'h437f6a62},
  {32'h453e45fe, 32'h4293ad79, 32'hc2469ae9},
  {32'hc4a14b1c, 32'hc2469d74, 32'hc4a8934b},
  {32'hc478d50a, 32'h43f3dee5, 32'h418263d4},
  {32'hc48dd601, 32'h43c9835c, 32'hc367349e},
  {32'h43a8e87f, 32'hc3a57771, 32'hc4e2805c},
  {32'h446ec99f, 32'hc3785849, 32'h43571c4d},
  {32'h4476eba6, 32'hc428c1ff, 32'hc42f2f36},
  {32'hc325c5e0, 32'h444cf1a8, 32'h44bbd3dc},
  {32'h45398166, 32'h43d57a7f, 32'h43d794ee},
  {32'hc4a2fbac, 32'hc4427032, 32'h44093083},
  {32'h45608ea5, 32'h4382bda8, 32'hc43cce16},
  {32'hc4f491c3, 32'h439ee097, 32'h4342515a},
  {32'hc3cb26a8, 32'hc4888b64, 32'hc31be3a4},
  {32'hc3649f63, 32'h44f7853b, 32'h44bd6cbb},
  {32'h44c7cba1, 32'hc282aa66, 32'hc2ada518},
  {32'hc4065554, 32'h44d7844e, 32'h4289c6b5},
  {32'h4550f573, 32'hc3b7db93, 32'hc423d5b5},
  {32'hc1bc8b80, 32'h433d7664, 32'hc420ec5c},
  {32'hc492d8a1, 32'hc2723922, 32'h44dc02ee},
  {32'h4432dd10, 32'h4368a87f, 32'h441a361f},
  {32'hc3ba7114, 32'hc5052692, 32'hc13c4f35},
  {32'h44ce24e0, 32'h436f9391, 32'hc3a6b079},
  {32'h449a3942, 32'h43645054, 32'hc3384701},
  {32'h448fd3e2, 32'h4504daf0, 32'h43c62769},
  {32'hc44d9740, 32'hc50b8a50, 32'h4360b7e3},
  {32'h4457d3be, 32'h43adce80, 32'h439444fb},
  {32'hc39fd900, 32'h43811880, 32'h446ea8a2},
  {32'hc35c4da0, 32'hc34b46ed, 32'h443fb910},
  {32'h43a7e7ee, 32'h41c1cf09, 32'h434ab6e0},
  {32'h4345d2e4, 32'h4400a433, 32'h43cd0efb},
  {32'h439e4ca4, 32'hc4c498a1, 32'hc4babf6a},
  {32'h4450846c, 32'h440a6bf3, 32'h434b4a73},
  {32'hc35a8670, 32'hc4446a7c, 32'hc4075379},
  {32'h440a0518, 32'h440aa2cf, 32'h447a866a},
  {32'hc1b3955a, 32'hc1ddd3f2, 32'hc488bfb9},
  {32'h453c2e87, 32'h433000db, 32'h43bfac29},
  {32'hc5809776, 32'hc3a09189, 32'hc330f3ff},
  {32'hc4ab2d7b, 32'h42fea8e0, 32'hc3c656da},
  {32'hc5404a33, 32'h420ae282, 32'hc36a8eed},
  {32'h44bcf756, 32'h438d828e, 32'h443695da},
  {32'hc4cfe5b5, 32'hc3ab60d2, 32'h424309c5},
  {32'h4436c35a, 32'hc2f67f5e, 32'hc2701d28},
  {32'hc49e509a, 32'hc387700a, 32'hc5008568},
  {32'h43c26912, 32'h42affc9c, 32'h44fcc679},
  {32'hc413a94b, 32'h43e446c9, 32'hc41e8d08},
  {32'hc41308b2, 32'hc479a80f, 32'hc436d02e},
  {32'hc3ad0a0c, 32'h456491e6, 32'h40a0d984},
  {32'hc5258508, 32'h433ab076, 32'h440e0a5e},
  {32'h43fdb9bc, 32'h44789ef9, 32'hc4144d6b},
  {32'hc48bcb08, 32'hc4b44a98, 32'h435b05c7},
  {32'hc2798860, 32'h43f4223a, 32'h42269ed8},
  {32'hc5274c27, 32'hc35e1a58, 32'h4343b39a},
  {32'h44f9747c, 32'h43548c24, 32'h43373ea8},
  {32'hc516290f, 32'h42f00a22, 32'hc319121d},
  {32'h439edb08, 32'h4465b14a, 32'hc4949f94},
  {32'hc3e52530, 32'hc51835a5, 32'hc2d7d919},
  {32'hc43e116a, 32'h43a7d8eb, 32'h40a91a10},
  {32'hc5019cde, 32'hc3df1d6b, 32'h4376f9a8},
  {32'h446a456c, 32'h44818558, 32'hc32c1fab},
  {32'h450c2bcf, 32'hc3a7173b, 32'h4231db0d},
  {32'h44ccb7d2, 32'hc2da15f6, 32'hc4400059},
  {32'hc3ae207f, 32'h4401e031, 32'h450a2125},
  {32'h454a542a, 32'hc35da9fa, 32'hc435f132},
  {32'hc38d479c, 32'hc3d4c70c, 32'h44ad9b08},
  {32'h4487691c, 32'h448b21ac, 32'hc40b58c5},
  {32'hc4395e9f, 32'hc45e06ef, 32'h4385b5e3},
  {32'hc25ae990, 32'h41e67422, 32'hc528fa9e},
  {32'hc4681564, 32'hc45b5abc, 32'h420ca92b},
  {32'h450ece96, 32'h43f969b2, 32'hc2e3d8bf},
  {32'hc4e277f4, 32'h439f4a04, 32'h44917374},
  {32'h443df26e, 32'hc36dbd04, 32'hc5391dcc},
  {32'h45104708, 32'hc4210311, 32'hc4119e8c},
  {32'hc481d812, 32'h44c0a6ce, 32'h43ebe7b7},
  {32'hc496e38f, 32'hc396b4ac, 32'hc23d7f84},
  {32'hc398ea10, 32'h448b7a6d, 32'hc3e45ac7},
  {32'h452bde58, 32'hc3af6a00, 32'hc20f3b6c},
  {32'h444bf650, 32'h447c6520, 32'hc263d2da},
  {32'h45067e61, 32'h43ed554e, 32'hc34480e8},
  {32'hc54298a8, 32'h443ba795, 32'h4389428c},
  {32'h43c8a74c, 32'hc32fa9d6, 32'h442022b5},
  {32'h43540608, 32'h43cdb936, 32'h44282c2a},
  {32'h449d95fe, 32'h441c92f7, 32'hc3d3f012},
  {32'h449b0d79, 32'h429f0c3e, 32'hc428445b},
  {32'h448186fd, 32'hc34f1f3c, 32'h435d2a1d},
  {32'hc441ccaf, 32'h443e9fc5, 32'hc44fe018},
  {32'hc3aa161a, 32'hc2c3af2b, 32'h4317499e},
  {32'hc4ae0f96, 32'hc2b0d71e, 32'hc481fb39},
  {32'h44fa740c, 32'h43a4e24b, 32'h42f1c55e},
  {32'h44c4caa1, 32'h43a45d24, 32'h44101b26},
  {32'h456883c2, 32'hc3e3e58c, 32'hc3783593},
  {32'hc409d817, 32'h449c502d, 32'hc2e7300b},
  {32'h4494dd70, 32'hc3ad813c, 32'hc3adb71b},
  {32'hc3d0373c, 32'hc41d3b82, 32'hc5494f46},
  {32'h43485ab7, 32'hc50d5e6c, 32'hc198a13c},
  {32'h44dcf752, 32'hc37c2af3, 32'h42e996ae},
  {32'hc33354e8, 32'h44786c44, 32'h455c476f},
  {32'hc40b498c, 32'hc3a0975c, 32'hc4cdaa65},
  {32'h4492670d, 32'hc38e835d, 32'h441c8d6c},
  {32'hc3c16854, 32'h4465b755, 32'hc49163e0},
  {32'h44e350f0, 32'h43fa107b, 32'h43b21db6},
  {32'hc401bb56, 32'hc385e879, 32'hc406f4e0},
  {32'h44a6939b, 32'h43091575, 32'hc41c9d66},
  {32'h451de500, 32'hc39ffe80, 32'h43b0770e},
  {32'hc495bd8c, 32'hc37b04cf, 32'hc46620a7},
  {32'h43c1a199, 32'hc4af340f, 32'hc30cad4c},
  {32'hc4f3023f, 32'hc21e970b, 32'hc45b52ba},
  {32'hc1759fe0, 32'hc495f977, 32'h4485d469},
  {32'h43a50400, 32'h43f7928e, 32'h451193cf},
  {32'hc551b7a0, 32'hc3113bd2, 32'hc35fd418},
  {32'hc1a663ba, 32'hc4ea1a54, 32'h44881d8c},
  {32'h443addba, 32'hc218dcf9, 32'h44e2f1cc},
  {32'h4257b4a0, 32'h45077dd5, 32'h438c41f2},
  {32'h43fd5169, 32'h433ba878, 32'h453e9748},
  {32'h43bd3c6e, 32'h4434e49d, 32'hc43d5adc},
  {32'hc3de09d0, 32'hc49220be, 32'h444e9c00},
  {32'h437a811a, 32'h42d5e9da, 32'hc514f3eb},
  {32'hc215e200, 32'hc41515c6, 32'h437336f2},
  {32'hc553e93f, 32'hc1f7fc41, 32'hc3b15884},
  {32'h449ffa66, 32'h438a0c2c, 32'h434183c6},
  {32'h44b75f65, 32'h446d1c78, 32'h41d6e136},
  {32'h45515b6b, 32'hc37a9e3c, 32'h43826b8b},
  {32'h4399a2d0, 32'h44c2e263, 32'h4423e971},
  {32'hc47e64bc, 32'hc2da91fa, 32'h439550cb},
  {32'hc56c2b4e, 32'h43376536, 32'hc3eb4b65},
  {32'hc2448440, 32'hc4a5ca1c, 32'h439086d8},
  {32'hc41418b9, 32'h44276d57, 32'h42b83339},
  {32'hc4d51ed3, 32'hc2d5c5b5, 32'hc45c8570},
  {32'h422b9122, 32'h444afc76, 32'h44d7cc25},
  {32'hc34e7172, 32'h419255a1, 32'h452ac423},
  {32'h446c49f8, 32'hc0da458c, 32'hc46d62d1},
  {32'h42eb874d, 32'hc50a84ae, 32'hc3bffe3d},
  {32'h44891082, 32'hc2d7b2fa, 32'hc4c5027a},
  {32'h438e4ac0, 32'hc4822f9c, 32'h44aa464e},
  {32'hc394a87e, 32'h442405c2, 32'hc2869625},
  {32'h444068d7, 32'hc499d608, 32'hc30cecaf},
  {32'hc401dd37, 32'hc5185874, 32'h44ed7f1c},
  {32'h448af40a, 32'h443e41cc, 32'hc492ac3f},
  {32'h43e1e9b8, 32'hc39ab8e7, 32'hc4fb2968},
  {32'hc4a061e1, 32'hc3060453, 32'h449d510a},
  {32'h43b5681e, 32'h41e14cbe, 32'hc2a6aaea},
  {32'hc3eaf072, 32'hc38e0d36, 32'hc22d0092},
  {32'h437b8cac, 32'h433cb53a, 32'hc41ed839},
  {32'hc39718cd, 32'hc4ec7f2e, 32'h3fa07910},
  {32'h456432e2, 32'hc3e001a6, 32'h43be36ba},
  {32'hc4a991cc, 32'hc3193388, 32'h4468fa95},
  {32'h454893ac, 32'hc2be1b64, 32'h4349e740},
  {32'hc2a38a8c, 32'hc5723c90, 32'hc31757d8},
  {32'h43ca5f0d, 32'h44f8f34c, 32'hc2b5a731},
  {32'hc5310888, 32'h429f5d2d, 32'h43375dfe},
  {32'hc139a3c0, 32'h45245c45, 32'h43503e83},
  {32'hc4dd39c2, 32'hc455bd2b, 32'h428b85c6},
  {32'h45037400, 32'hc41c464e, 32'hc3ae6c4b},
  {32'h439bb858, 32'h441d1ff1, 32'h42115a4e},
  {32'h43c234b7, 32'h44e29bcc, 32'hc50dd178},
  {32'h420d0dba, 32'hc4a4cacf, 32'h4516c04d},
  {32'h44fc68fd, 32'h43ae8f15, 32'hc343efeb},
  {32'h4438c01e, 32'h44d777be, 32'h445c388b},
  {32'hc4d2b858, 32'hc38bb2de, 32'hc36b2552},
  {32'h42456d64, 32'h425b23c3, 32'h44c4af42},
  {32'hc3289da6, 32'hc48e6dc0, 32'hc520af2d},
  {32'h43a913f0, 32'h447d8bee, 32'h44d0b327},
  {32'hc284d608, 32'hc398c58e, 32'hc3f5dbda},
  {32'h435d1965, 32'h431d7329, 32'h44a2b456},
  {32'hc39beb2e, 32'h44d2b11f, 32'hc4b6d072},
  {32'h44df83d9, 32'hc2fa63e7, 32'h42eadcb8},
  {32'hc3689369, 32'hc3bc6f2b, 32'hc4d7bc62},
  {32'h44f41e3c, 32'h4302411f, 32'h43a6324d},
  {32'h448e1dee, 32'h42ac7c55, 32'h4327b465},
  {32'h4502c094, 32'h421fad86, 32'h43b18258},
  {32'hc543cdbc, 32'h42b69ce9, 32'hc3b2725a},
  {32'hc3933d3a, 32'h4469183e, 32'hc2bfcc06},
  {32'hc57e8c37, 32'hc3d63de9, 32'hc1e8b806},
  {32'h45040681, 32'h445904d2, 32'h44514f7d},
  {32'h4316ea89, 32'hc3c580dc, 32'hc382bb2d},
  {32'hc1d2e044, 32'h4507ebdd, 32'hc3a48866},
  {32'hc32e2ba0, 32'hc51b851b, 32'hc40ca481},
  {32'h44d95077, 32'h43865481, 32'h43efcbef},
  {32'hc54bd01e, 32'hc38cc159, 32'hc3647509},
  {32'h4524e483, 32'h43ade27c, 32'h420d3111},
  {32'h448ec924, 32'hc3d7fd85, 32'h434a14fa},
  {32'h437b2d75, 32'h43b9f8f8, 32'h438c3646},
  {32'h44595fc7, 32'h447b45f4, 32'hc256627a},
  {32'h434d43f0, 32'h44706739, 32'h450ff7f5},
  {32'h442d7a8a, 32'hc4cc84a6, 32'hc40059c1},
  {32'hc49f00b4, 32'h4256c16f, 32'h43d4daa7},
  {32'h44d76030, 32'hc466ee0c, 32'hc4435984},
  {32'hc50cacf4, 32'h4393af50, 32'h445c3bfd},
  {32'hc4790905, 32'h43b3a9b9, 32'hc4b7a9f6},
  {32'h4430e147, 32'hc45f7a09, 32'h450cd40a},
  {32'hc3fb66f3, 32'h44c9eb4c, 32'hc5054ab9},
  {32'h441d7fec, 32'h42eb71b7, 32'hc2d47f1e},
  {32'hc3e6c01c, 32'hc50bf25f, 32'hc42e341e},
  {32'hc4329697, 32'hc390c327, 32'h450bd509},
  {32'h4398debe, 32'h3fa2e91a, 32'hc483d6ca},
  {32'hc3710869, 32'h43d16eb8, 32'h4414629f},
  {32'h43dbb577, 32'hc1f6b272, 32'hc540c478},
  {32'h44852f5c, 32'hc3b70d56, 32'h43af63c2},
  {32'h42c0b84e, 32'hc4fab4b7, 32'h42076683},
  {32'hc527a6da, 32'hc357fb91, 32'hc2a29688},
  {32'h44b867f8, 32'h41be22ed, 32'hc39acc80},
  {32'hc520b444, 32'h44221bc9, 32'h42cdf62d},
  {32'h438a6890, 32'hc46e5024, 32'hc2afbed9},
  {32'hc4d29985, 32'h441e2c03, 32'hc3152d49},
  {32'h456e1c00, 32'h438dd48d, 32'h43e7a158},
  {32'hc5423fca, 32'h43925556, 32'hc17fac44},
  {32'h45524392, 32'hc403d0ef, 32'hc37659b9},
  {32'h440c9069, 32'h433b0e22, 32'h44d539ec},
  {32'hc4e5b597, 32'hc3bb595f, 32'hc3c920c3},
  {32'h44a27108, 32'h4296ef7f, 32'h451b0d31},
  {32'hc49871f3, 32'h43cf031d, 32'hc3094160},
  {32'h44edda7a, 32'hc4c3bf6b, 32'hc3891558},
  {32'hc5022abe, 32'h438fb5da, 32'h43b4d9d1},
  {32'h44397674, 32'hc431354b, 32'hc3611f6b},
  {32'hc390d614, 32'h4565c54a, 32'hc33ec201},
  {32'hc2b62520, 32'hc4960185, 32'h43cb2286},
  {32'h4471c6b8, 32'hc38c933b, 32'hc465031f},
  {32'h44ab9dcc, 32'h4434f59f, 32'hc3745911},
  {32'hc519ae57, 32'h43a1939e, 32'h43e10771},
  {32'h43363d15, 32'hc496f968, 32'hc4024289},
  {32'h43bdf85c, 32'h44afe519, 32'h43fdb434},
  {32'h4529ed50, 32'h4363de9f, 32'h4203dc44},
  {32'hc2b93930, 32'hc376b957, 32'h4206dd90},
  {32'hc2a25990, 32'hc3b25b71, 32'hc4a1adf3},
  {32'hc51da2cb, 32'hc3ace859, 32'h42c7d281},
  {32'h4498ed33, 32'hc2732331, 32'hc30884d8},
  {32'hc5453930, 32'hc2a81756, 32'h440f2d89},
  {32'h450c853b, 32'h4439dfcf, 32'hc389bfa5},
  {32'h42208d3c, 32'h43cc175d, 32'h441b18b5},
  {32'h44e87dd6, 32'hc456bcd4, 32'hc25cae04},
  {32'hc482030c, 32'h440638fd, 32'hc244f3aa},
  {32'hc4770244, 32'hc35ff971, 32'hc3f4907d},
  {32'hc34414d4, 32'h439621c0, 32'h451c4af3},
  {32'h434e4ab0, 32'hc4582340, 32'hc53f9f2e},
  {32'h44d18401, 32'h433379b8, 32'hc4d6ca3f},
  {32'hc4ffbf76, 32'h41974093, 32'hc019f025},
  {32'h44658544, 32'h43901d80, 32'hc40417d0},
  {32'hc4066ead, 32'hc5129745, 32'hc408536e},
  {32'h43c0b280, 32'h4525d6e4, 32'hc1454026},
  {32'hc4463ba2, 32'hc3903cd7, 32'h43931007},
  {32'h4491468e, 32'h44ff1523, 32'hc30c221c},
  {32'hc2a887d8, 32'hc584353f, 32'h42a7714d},
  {32'h433d8cb1, 32'h4500810b, 32'hc399f570},
  {32'hc2b2d236, 32'hc430de3e, 32'h453c63c5},
  {32'h44aa27b2, 32'h433b4a3c, 32'h43b9af61},
  {32'h44884271, 32'hc2e916fa, 32'h40b6bb52},
  {32'h448241fa, 32'h448fb615, 32'h44210740},
  {32'h43b85d12, 32'hc4b9c0e9, 32'hc4cd311c},
  {32'hc45a82e0, 32'h440c3c03, 32'h4407ee85},
  {32'hc2271330, 32'hc341a939, 32'hc522c73d},
  {32'h44ee356c, 32'h43dc438e, 32'hc2fb0cc0},
  {32'hc33ac5b3, 32'hc4335332, 32'hc40f6b0b},
  {32'h448e2d6b, 32'h4411eeed, 32'h44b50c42},
  {32'hc215e300, 32'h43f147bc, 32'hc4a598ae},
  {32'h454dbc5a, 32'hc380686f, 32'hc432e006},
  {32'hc3598bb8, 32'hc4ee6f02, 32'hc3e2b8dd},
  {32'h4498fe06, 32'h4435149e, 32'h4436a676},
  {32'h442f97d0, 32'hc396129f, 32'h43b8fb55},
  {32'h44b2fec4, 32'h43e03887, 32'h4479d6ef},
  {32'h4324cda6, 32'hc4ded2e8, 32'hc4a26d65},
  {32'hc4bbe72a, 32'hc24d6b87, 32'h43932f03},
  {32'h44196861, 32'h449458c6, 32'hc364eec0},
  {32'hc41b7a42, 32'hc494b900, 32'hc3af68b7},
  {32'h450b64e1, 32'h44306830, 32'hc3102cc7},
  {32'h44ad906e, 32'h431fadd9, 32'h43009ac1},
  {32'h44f918d4, 32'h445059de, 32'hc33c0aba},
  {32'hc4947f7a, 32'hc4444d7e, 32'hc1c21fdc},
  {32'hc3c2ccb2, 32'h43a846c0, 32'hc3800cc3},
  {32'hc5066f42, 32'hc394a0f7, 32'h426cae71},
  {32'hc383d440, 32'h43fd98fb, 32'h444590c4},
  {32'h44b5f40d, 32'hc3cc8026, 32'h4432893f},
  {32'h438c0202, 32'h4493e878, 32'hc4110cfe},
  {32'hc49a35c2, 32'h418759e8, 32'hc43531d0},
  {32'hc49c94fd, 32'h435aa123, 32'hc3a56640},
  {32'hc3620228, 32'hc422d117, 32'h448b27dd},
  {32'hc31248a4, 32'h44097238, 32'hc46b6875},
  {32'h44520522, 32'h420d050e, 32'h43fcec62},
  {32'h435cfc58, 32'h444be364, 32'h4477e4b9},
  {32'hc3cee5e2, 32'h43ccaaf2, 32'h4544a84f},
  {32'h4288565e, 32'h442b03bb, 32'hc4bfb626},
  {32'hc4198af3, 32'hc495f6fb, 32'hc3753710},
  {32'h44ec27ea, 32'h44972248, 32'hc352dd7a},
  {32'hc4a8f31f, 32'h43c7a7e2, 32'h43934fe1},
  {32'h44ba362c, 32'h43ca2239, 32'hc4a494c5},
  {32'hc5251031, 32'hc2179152, 32'h441f0a55},
  {32'h44d269e7, 32'hc283c582, 32'hc443bb41},
  {32'hc28e22d1, 32'h43e85b01, 32'h455873fa},
  {32'h4505986f, 32'hc42736e9, 32'hc4993085},
  {32'hc3e42428, 32'hc2f4a651, 32'hc4ab0551},
  {32'hc41bcaee, 32'h440b39ac, 32'h448e692b},
  {32'hc49a422f, 32'hc2cc03c9, 32'h435573c7},
  {32'hc4ff1270, 32'h43c2eed8, 32'hc150a82e},
  {32'h4551c7ed, 32'h4397378d, 32'hc0bcdb80},
  {32'h4501648b, 32'h4317d4df, 32'h4199d71a},
  {32'h4441a7b3, 32'h43c0ae3d, 32'h41f03201},
  {32'hc4d0797c, 32'hc302d617, 32'h41b0e1b1},
  {32'h4555149e, 32'h43b5b5b0, 32'h441e8b96},
  {32'hc4fe42a5, 32'hc3a6aaea, 32'h440ff724},
  {32'h438a182e, 32'hc407b234, 32'h44d8685a},
  {32'hc4c01884, 32'hc1afda2e, 32'hc449eff5},
  {32'hc3c373e5, 32'hc4dbbbdb, 32'h44338df7},
  {32'hc3b1119c, 32'h44a522f2, 32'hc3e58f49},
  {32'h4400e414, 32'hc3800cf0, 32'h4453e22e},
  {32'hc0c54cc0, 32'h4472aae1, 32'h444551a1},
  {32'h440c282e, 32'hc1145218, 32'h4291bdfd},
  {32'hc505119b, 32'h439ea8f5, 32'h438a0185},
  {32'h44eb6b08, 32'hc3f8e9db, 32'h43b4fc1e},
  {32'hc5090f12, 32'h440f2244, 32'h43fabec9},
  {32'h444cfcf2, 32'hc46ffa52, 32'hc1a0f1f4},
  {32'hc3edf2a1, 32'h44f59794, 32'hc24a8de8},
  {32'hc3af7f7e, 32'hc45fa9bd, 32'h448c96b7},
  {32'h43aeb20a, 32'h43c00f50, 32'hc3d0147b},
  {32'h44713752, 32'hc182b9f6, 32'h44ac5560},
  {32'hc2d58fa0, 32'hc36b823a, 32'hc4b95120},
  {32'hc2ebfc8c, 32'hc43ca14a, 32'hc22a4eb8},
  {32'hc3ad998e, 32'hc4fa323c, 32'hc487bd70},
  {32'hc3f6f30f, 32'h441536f1, 32'h44a21d42},
  {32'h439dbdc3, 32'hc4a948f5, 32'hc3fb993e},
  {32'hc4ac7b0b, 32'h43b7ec06, 32'hc21c0bc7},
  {32'h44baf911, 32'hc30a1a36, 32'h449bb6e6},
  {32'hc2ba2748, 32'h44e0bab7, 32'h438b1ba7},
  {32'h44dc9c2c, 32'hc3d60a76, 32'hc1d37514},
  {32'hc4e0f9ce, 32'h43b0b47f, 32'hc4695137},
  {32'h42136f50, 32'hc4822216, 32'hc281bccc},
  {32'h432f8a7a, 32'hc482b281, 32'h4500ac9c},
  {32'hc42f28c9, 32'h4488bf2a, 32'hc4ae64f3},
  {32'h44a938ed, 32'hc3e7cee3, 32'h42ffe468},
  {32'h42b1a100, 32'hc36b08f4, 32'h43da6357},
  {32'hc2a52c28, 32'h44717e78, 32'hc4231224},
  {32'h44d4d90e, 32'h43d3f539, 32'h435b3225},
  {32'h43b082b4, 32'h442034e6, 32'hc46efceb},
  {32'h443f0249, 32'h42d5f8b3, 32'h44ec18cc},
  {32'hc327a40e, 32'h453ae2f9, 32'h43831260},
  {32'h45634f09, 32'hc41b2c8d, 32'h43bfc2db},
  {32'hc59312a5, 32'hc3e15ae1, 32'h423ea006},
  {32'h456fd13c, 32'h444e5dd7, 32'hc4024f2a},
  {32'hc49774cd, 32'hc238e5ad, 32'h4380e115},
  {32'h447f480f, 32'hc50d47c8, 32'h4417a4da},
  {32'hc5436b81, 32'h42635c0c, 32'h43f0166a},
  {32'h4234d2c0, 32'hc50b92f8, 32'hc2d79df2},
  {32'hc3996f27, 32'h455065a4, 32'h43ffd939},
  {32'h4519ba39, 32'hc4830826, 32'h43142174},
  {32'h4362386a, 32'h44d0cc8f, 32'h43e8f086},
  {32'hc367862e, 32'h44d1d7a2, 32'hc498dc4d},
  {32'hc4bbf259, 32'h44099bae, 32'h440e5293},
  {32'hc3ed5b02, 32'hc450a937, 32'h4405aa08},
  {32'h44abd1dd, 32'hc334ea9e, 32'hc4ad6493},
  {32'h44c177a3, 32'hc38f73c6, 32'h43788502},
  {32'h43f57d22, 32'h4421a062, 32'hc3e09e0c},
  {32'hc4e589d5, 32'hc43a5ac4, 32'h43e1d83a},
  {32'h4498a999, 32'h438b91ca, 32'hc455784e},
  {32'h441669c3, 32'h43bbeeca, 32'hc29a2a3d},
  {32'h43becf90, 32'h441930db, 32'h446ec08e},
  {32'h421a9f68, 32'hc43c4a81, 32'hc514f1c0},
  {32'h443b8b00, 32'h44250f76, 32'hc4067d4a},
  {32'hc314e48f, 32'hc2fb9415, 32'h45687b4b},
  {32'hc4516081, 32'h43e99654, 32'hc3f832e4},
  {32'hc389c898, 32'hc4f9f0a1, 32'hc148bbba},
  {32'h440732d2, 32'h43a2fad0, 32'hc44a05fd},
  {32'hc3a5d70e, 32'hc4a88c75, 32'h43bd558a},
  {32'h44e964a6, 32'hc418e9ca, 32'hc20bcda8},
  {32'hc4903940, 32'h42ab0744, 32'h44248f86},
  {32'h455c546d, 32'hc2b32bfa, 32'h4350b261},
  {32'hc5247699, 32'hc42737e0, 32'h4216968f},
  {32'h43d7d1f4, 32'h44e43a1d, 32'hc2ad9de4},
  {32'h444616b2, 32'hc2fd2691, 32'hc30afd96},
  {32'h450813b8, 32'h4451be6a, 32'h43c237c2},
  {32'hc460e9b4, 32'hc4c42d74, 32'hc2e3bfb2},
  {32'h4483ea10, 32'hc383f119, 32'hc4332759},
  {32'h408bee00, 32'h43bc3352, 32'hc0b8d11d},
  {32'hc50e29c8, 32'hc29d9728, 32'hc41a184d},
  {32'h42ac45d4, 32'h44c12fe5, 32'h445f3e6e},
  {32'h40191e00, 32'hc301e58d, 32'hc39537b0},
  {32'hc2c92891, 32'hc2b8d711, 32'hc366d499},
  {32'hc304b2fb, 32'hc326b7a8, 32'hc5534f00},
  {32'hc02bc8e0, 32'h44cd549c, 32'h43c0ad5d},
  {32'hc3ff2417, 32'hc3e88bca, 32'hc55fd064},
  {32'h44626085, 32'h43b2b01a, 32'h452d03d3},
  {32'h430f5e73, 32'h442530ec, 32'hc3bc3d03},
  {32'hc328c6b9, 32'h42502a36, 32'h445400ef},
  {32'hc2ff1c8c, 32'hc4fbe930, 32'hc42f6ced},
  {32'h43d57e38, 32'h43f36dad, 32'h445c18e2},
  {32'hc3bc67ac, 32'h42e527bd, 32'hc5268286},
  {32'h44197c93, 32'h4406b213, 32'h448c7de2},
  {32'hc50bc7f2, 32'hc2df540e, 32'hc1973764},
  {32'h44c7e303, 32'h42a7e503, 32'h433452c6},
  {32'h43be2f42, 32'hc4845fbc, 32'hc50ef716},
  {32'h454e689d, 32'hc3aee25f, 32'h43859eb4},
  {32'hc5193589, 32'hc3f73a49, 32'hc3bc66cd},
  {32'h4480c261, 32'h449bca98, 32'h4274525d},
  {32'hc3d534ce, 32'h41bb2b28, 32'hc33ee2e8},
  {32'h45579f9e, 32'h419e36e4, 32'h43e21fb5},
  {32'hc47429ba, 32'hc3f5b85d, 32'h44190595},
  {32'h4394bdeb, 32'hc3589ff3, 32'hc2e15a2e},
  {32'hc4df8138, 32'h4213d3d1, 32'h43b7947e},
  {32'h44fcd92a, 32'h42f6d143, 32'h4297abca},
  {32'h443fd378, 32'hc491a3d1, 32'hc464c30f},
  {32'h43a203fa, 32'hc51b5a09, 32'h44bdfac4},
  {32'h43209a0c, 32'hc3b1b4ec, 32'hc3c9c84e},
  {32'hc344cab4, 32'h450b9cca, 32'h43c0356f},
  {32'h44140361, 32'hc32a78cf, 32'hc4c45148},
  {32'hc4199729, 32'h4474d009, 32'h42f70ae1},
  {32'h4233fd80, 32'hc3c90d46, 32'hc4a6f4cc},
  {32'hc3a2821e, 32'h440b09a2, 32'h453b4f87},
  {32'h43b07497, 32'h424955c4, 32'hc5176db0},
  {32'hc50e5c78, 32'h42a6c7e4, 32'h44202e7e},
  {32'hc3a0d3c9, 32'hc46acd9a, 32'hc470b3eb},
  {32'h4454682d, 32'hc30960ea, 32'h434e5fae},
  {32'h3fc54f80, 32'hc3514fcd, 32'hc4db6e1f},
  {32'hc44b9cea, 32'h44a9d805, 32'h441803a4},
  {32'h4425f836, 32'hc330163d, 32'hc391e70d},
  {32'hc3583848, 32'h447e8e58, 32'h44d704fb},
  {32'h44e658a2, 32'h438a0507, 32'hc46d3e64},
  {32'h43d8770f, 32'h4465b3cc, 32'h44126f37},
  {32'h43b9b856, 32'hc559dd46, 32'h432314a7},
  {32'hc3e357be, 32'h4533fd2c, 32'h43a250df},
  {32'hc4b39ea5, 32'h428b5db4, 32'h4342a6d8},
  {32'hc3daa558, 32'h4520ee9f, 32'hc002f2e0},
  {32'h447ed018, 32'hc4ce9863, 32'h43445d2a},
  {32'h43e67d76, 32'h44065325, 32'h432850b7},
  {32'h4546639c, 32'h440a76f8, 32'hc3029da3},
  {32'hc51ea2bc, 32'hc3a3b15e, 32'h43a6ac02},
  {32'h454b21c0, 32'hc2a8b45a, 32'h4374543f},
  {32'hc4611a7d, 32'h42e9fcb6, 32'hc29ada9d},
  {32'hc516bfac, 32'hc281e5f0, 32'hc28d7d39},
  {32'h4503c8aa, 32'hc2e8441a, 32'h4483ab0c},
  {32'hc3766d3a, 32'h43ae13d7, 32'hc331a30d},
  {32'h44bb739b, 32'hc4c0757e, 32'hc2b1a311},
  {32'hc3b7e033, 32'h451e5aae, 32'h43cb746d},
  {32'hc4b4479d, 32'hc304962c, 32'h43466bf3},
  {32'hc4227004, 32'h452243ca, 32'hc2debd56},
  {32'h44f3a43a, 32'hc48a041e, 32'h42d1d4ee},
  {32'h44ee0587, 32'h439fc1ff, 32'h4337ef8d},
  {32'h4541c694, 32'h42754a69, 32'hc3859402},
  {32'hc46389e6, 32'hc356fffe, 32'hc37abe29},
  {32'h45218c62, 32'hc3065850, 32'h439a7499},
  {32'hc50ffbd5, 32'h441a4990, 32'hc2398c7f},
  {32'hc2f241c1, 32'hc504d4f7, 32'hc45e1024},
  {32'h4414f6d5, 32'h440dc2b4, 32'h44e239d8},
  {32'h44db9c17, 32'hc46139b2, 32'hc3ad6186},
  {32'hc3b34270, 32'h44ab8590, 32'h43b4d99b},
  {32'hc44c993b, 32'h42c78fde, 32'hc39caa9b},
  {32'hc4e03d51, 32'hc46436cc, 32'h43b7462a},
  {32'h4350eec8, 32'h43aa4034, 32'hc4a99901},
  {32'h41012ee8, 32'h44f395bd, 32'hc3c4f516},
  {32'h4460c1d0, 32'hc40374ff, 32'hc424d07b},
  {32'hc39f4047, 32'h443b6ff6, 32'h44d2d8fd},
  {32'hc1e68370, 32'hc49bad05, 32'hc39277eb},
  {32'hc47fd0c8, 32'h4435ccc1, 32'h44f359e6},
  {32'hbefa6000, 32'hc3dd8582, 32'hc5224995},
  {32'h451d904c, 32'h42728fe1, 32'hc45904f5},
  {32'hc513d210, 32'hc2d65ca6, 32'h4405bf80},
  {32'h43a62888, 32'h44765b5d, 32'hc492d732},
  {32'hc3a4d54e, 32'hc4aea7f6, 32'hc1d228e3},
  {32'h43bbb096, 32'h44f1e07c, 32'h4280f1d2},
  {32'hc41ba734, 32'hc3f32834, 32'hc2d7acc0},
  {32'h4169bf00, 32'h44653457, 32'h439c3953},
  {32'hc336bda0, 32'hc505f141, 32'hc42193eb},
  {32'hc41e7d4b, 32'h43ee7d9c, 32'h43b59346},
  {32'hc46557d8, 32'hc3cd4138, 32'hc3513d90},
  {32'h45380622, 32'h4310daae, 32'h43d29a3c},
  {32'h448dbfb8, 32'hc1fc86aa, 32'h435f24a5},
  {32'h44c1b39b, 32'h442fa1f3, 32'h43893f4b},
  {32'hc35f86e8, 32'hc2a3e310, 32'hc34cc9f3},
  {32'h422b89cd, 32'h44a5dc88, 32'h42c412d9},
  {32'hc481adae, 32'hc3dd9daa, 32'hc2f835ed},
  {32'hc1c55430, 32'hc2db73a0, 32'h448332b7},
  {32'hc4e7007a, 32'hc34fad64, 32'h43932c6d},
  {32'hc2a178ee, 32'h443c7387, 32'h445905e1},
  {32'hc48e7b68, 32'hc443e446, 32'hc478dd89},
  {32'h451ed8e5, 32'h448fb8d0, 32'hc392946b},
  {32'hc32e1e3c, 32'hc471456e, 32'hc4ca7b69},
  {32'hc3a3cd83, 32'h438926a5, 32'h45340765},
  {32'hc4b659de, 32'h41f17080, 32'hc3c49eca},
  {32'h43ed71a0, 32'h44b05aac, 32'h44065bab},
  {32'hc3b2f04a, 32'hc52aa609, 32'hc38036ee},
  {32'h45089fc4, 32'hc28e8d08, 32'hc403d455},
  {32'h44543e05, 32'h43b74224, 32'h40a1dddc},
  {32'hc49cc7ab, 32'hc457fc0a, 32'h42cf8a5d},
  {32'h44bd62e8, 32'h44acca47, 32'h41d9d1e5},
  {32'hc4edacd9, 32'h43b61665, 32'h43b6fead},
  {32'h43232eaa, 32'h45070886, 32'h4328701d},
  {32'hc51587c9, 32'hc3864ac9, 32'h42f6a026},
  {32'h44f35a4d, 32'hc23ec200, 32'hc34d8eae},
  {32'hc585cc93, 32'h43ab9826, 32'hc3440f58},
  {32'h4555c697, 32'hc406b989, 32'h442be5b3},
  {32'hc402ac41, 32'hc3f13e37, 32'h4347ef19},
  {32'h43f2c5a1, 32'h440bbc91, 32'hc3b1e037},
  {32'hc16f3914, 32'hc4f274ce, 32'hc2d22cf7},
  {32'h45494ee8, 32'h43ea6a2c, 32'hc305c658},
  {32'hc46e3f17, 32'hc4537f15, 32'hc2281db2},
  {32'h441fd4ef, 32'hc2e32701, 32'hc4eebd56},
  {32'hc39dc4cb, 32'hc34dd891, 32'h44b43e05},
  {32'h4549c7b2, 32'hc3bae737, 32'hc39a5673},
  {32'hc49d6702, 32'hc3eb6f2a, 32'h426bdd41},
  {32'h44bd0f32, 32'hc2f37f29, 32'h440244b1},
  {32'hc4a2bf5c, 32'hc4b0caf0, 32'h4311356f},
  {32'h44de6fdf, 32'h43e08355, 32'hc3f487d8},
  {32'hc466defa, 32'h42edd5df, 32'h43b43887},
  {32'hc3a4c053, 32'h43628c82, 32'hc5262f85},
  {32'hc41b9c52, 32'h439c619d, 32'h44bf07b7},
  {32'h44c2a5be, 32'h41c51501, 32'hc3a11b2a},
  {32'hc528d44f, 32'hc2e30286, 32'h446b0b42},
  {32'h4521f06b, 32'h43171064, 32'hc42cf4f7},
  {32'h43b4b044, 32'hc502f9f7, 32'hc2b245c8},
  {32'hc4ba16f0, 32'h44e9ded0, 32'h42e93691},
  {32'h442827c1, 32'hc23540ac, 32'h413d0bff},
  {32'hc3c486f2, 32'h4515e777, 32'h4320a6aa},
  {32'h44b63c7c, 32'hc434756c, 32'h431d9b21},
  {32'hc4d3a051, 32'hc38a2b14, 32'hc37b5f01},
  {32'hc3d9a67c, 32'h43e6d358, 32'hc27dc5fd},
  {32'hc4b67120, 32'h4420a590, 32'h4415ddf1},
  {32'h43b1191c, 32'hc303ad0c, 32'h43c0f4e3},
  {32'hc481a06e, 32'h43b822ca, 32'h42d79711},
  {32'h44c266b0, 32'hc390ded6, 32'h435cb51a},
  {32'hc40bffef, 32'h43c411b1, 32'hc45c5d69},
  {32'hc286c118, 32'hc50e08e4, 32'h42aecc96},
  {32'hc478abad, 32'h43e67064, 32'hc4b0792f},
  {32'h44f5243f, 32'h43d0b1af, 32'h4296822d},
  {32'hc4a07a24, 32'hc35f2c96, 32'hc4d2d6c8},
  {32'h45322e96, 32'hc39b5563, 32'hc21242c3},
  {32'hc3a1457e, 32'h4406664b, 32'h43c3f366},
  {32'h45278fd4, 32'hc4163fd8, 32'h43526907},
  {32'hc48fab42, 32'h4489c388, 32'hc5158ec6},
  {32'h42b49d0c, 32'hc3ab7b6a, 32'h444b7bfc},
  {32'hc44d51da, 32'h43a7f74e, 32'hc50bd882},
  {32'hc31c965e, 32'hc337e632, 32'h452f09a7},
  {32'hc369c676, 32'h44cb18fb, 32'h43a9d599},
  {32'hc21efc46, 32'h43aef0aa, 32'h453a5531},
  {32'hc527d3e0, 32'hc3c13400, 32'hc4d2c624},
  {32'h44d8219d, 32'hc3ae54d9, 32'hc2814927},
  {32'hc2facfd4, 32'h43e17147, 32'hc47e14b2},
  {32'h441cd7f8, 32'h449c7f64, 32'h4486b626},
  {32'hc4c15f35, 32'h42e388b4, 32'h42e2db2d},
  {32'h44cba674, 32'hc326335a, 32'hc32cfbba},
  {32'h44775277, 32'hc3f4a141, 32'h432ed3de},
  {32'hc4ac8439, 32'hc1e9fa78, 32'hc3e01b8f},
  {32'hc4b1a625, 32'h442ae27a, 32'h43b24fc8},
  {32'hc496bd2d, 32'h44b91145, 32'hc39da268},
  {32'hc1ec6670, 32'hc532d3a3, 32'h438b3916},
  {32'h432dcb4c, 32'hc4c3c08f, 32'h452cbd72},
  {32'hc50cfad0, 32'hc4150ddb, 32'hc255cf61},
  {32'hc3bd3a09, 32'h4001b680, 32'h4500ff70},
  {32'hc315fed4, 32'hc31c11fb, 32'h44a56bb6},
  {32'hc54dfbbc, 32'hc3372248, 32'hc3455af5},
  {32'h448dbc07, 32'hc300fa39, 32'h44b8876e},
  {32'hc51f876b, 32'hc24dfda0, 32'h3ffc3d10},
  {32'h4493cb0c, 32'hc2e2dcfc, 32'h44307236},
  {32'h42c40e60, 32'h4495d39e, 32'hc442d6d1},
  {32'h456ee1be, 32'hc3893e2b, 32'h428ddf15},
  {32'hc59bdf43, 32'hc137c608, 32'h42ab79ae},
  {32'h454c3cec, 32'hc2abad3f, 32'h44025af3},
  {32'h441ed052, 32'h43487bf3, 32'hc420a9c7},
  {32'h44dd046d, 32'hc3fe262b, 32'h42b75a91},
  {32'hc2838858, 32'h45312d34, 32'hc38afbaf},
  {32'hc42d658e, 32'h403131f0, 32'h432316a8},
  {32'hc3208170, 32'h44afc773, 32'h442e0cbe},
  {32'hc2a693b8, 32'hc51bdb8c, 32'h41a2d88f},
  {32'h449fd341, 32'h43fdd2f1, 32'hc280f8d4},
  {32'h4390a705, 32'hc484a0b9, 32'hc4081d09},
  {32'hc3a2518b, 32'hc5171317, 32'h448ee8ee},
  {32'h42b3f670, 32'hc509ab0c, 32'h443f8017},
  {32'h4350adb0, 32'h430b07d8, 32'hc4ab05ea},
  {32'hc433ef85, 32'hc238ae4d, 32'h4469a20f},
  {32'h44af5216, 32'h4381b963, 32'hc3c81025},
  {32'hc491c252, 32'hc3b9810e, 32'h4348bbb7},
  {32'h43b6c3f4, 32'hc3478f28, 32'h43962948},
  {32'h43b297b1, 32'hc4aff051, 32'hc3a4f280},
  {32'h441d2a13, 32'h43df0f9f, 32'h45400e3d},
  {32'hc3857a60, 32'h43f8c22f, 32'hc51e4ace},
  {32'h4252bacf, 32'hc314f2b6, 32'hc50370dd},
  {32'hc519515b, 32'hc3ab5135, 32'h4357b84b},
  {32'h447ea7bc, 32'h43cf9218, 32'hc3a50c43},
  {32'hc4f0b1ee, 32'hc1fa3be7, 32'h441498b7},
  {32'h4281c5b8, 32'hc3895a19, 32'hc526fda8},
  {32'hc3feccd0, 32'hc45fb0c2, 32'hc285c9e0},
  {32'h44b5d77c, 32'hc36461de, 32'hc335814c},
  {32'hc59afdca, 32'hc40678fd, 32'h436fe8dc},
  {32'h4527c946, 32'hc3921e83, 32'hc28f2ca2},
  {32'hc40c1b5f, 32'hc519afc7, 32'h43afc2e0},
  {32'h44315d78, 32'h44ae9f71, 32'hbfc65ee0},
  {32'hc526becc, 32'hc1fe9389, 32'hc2dc25a9},
  {32'h44afebf9, 32'h44b9b7cd, 32'hc3e74f85},
  {32'hc432092d, 32'hc4cc55ef, 32'h439dcd65},
  {32'h43371a62, 32'h44907378, 32'hc0fbfc91},
  {32'hc2920cae, 32'h440f7c1d, 32'hc31589c5},
  {32'h436f1d60, 32'h4424b023, 32'hc503c43a},
  {32'hc38b665c, 32'h44346fe2, 32'h4469d0f0},
  {32'hc4be38e4, 32'hc3390a96, 32'hc2ce4f23},
  {32'h444c0f29, 32'h44e2ac2d, 32'h4380991f},
  {32'hc4c63605, 32'hc4276570, 32'hc29069c7},
  {32'h43aca852, 32'h446390dc, 32'h43e1c040},
  {32'hc3c9a720, 32'hc2d4491b, 32'hc496d0b5},
  {32'h43fb284f, 32'h43f31433, 32'h4544d67c},
  {32'hc3f874ea, 32'h44910d59, 32'hc389892f},
  {32'hc44be4f1, 32'hc4b730f6, 32'h44e0b0f5},
  {32'hc3094750, 32'h4384ebb8, 32'hc29a88d3},
  {32'h4529a3ae, 32'h429f8149, 32'h43c04cb4},
  {32'hc517b325, 32'hc4001f1c, 32'h42f6aac2},
  {32'h43ac17d3, 32'h450d4c18, 32'hc40232e9},
  {32'h43cafa3c, 32'hc4550c7b, 32'hc49df9a9},
  {32'hc400ac2b, 32'h44a75de4, 32'h450cc7cf},
  {32'hc4d52c88, 32'hc38cb1f8, 32'hc495fb7e},
  {32'hc400c8b1, 32'h443d3147, 32'h438c06ff},
  {32'hc4c6a3c2, 32'hc49973f4, 32'h41e9b225},
  {32'h435a4bab, 32'h453ed325, 32'h4305b75f},
  {32'h4413736d, 32'hc39144f6, 32'hc3781265},
  {32'h446b9a52, 32'h442b6fd6, 32'h441ce36b},
  {32'hc3f99dee, 32'hc556ac09, 32'hc3957d9d},
  {32'hc4e9443b, 32'h42e73fb9, 32'h3f4d2a9c},
  {32'hc589e20d, 32'h42961a59, 32'hc2fe8e77},
  {32'h455214af, 32'hc29d60b2, 32'hc32d918d},
  {32'h42f9872f, 32'h448632d3, 32'hc498d1c0},
  {32'hc36c102d, 32'hc37b1a1f, 32'h443d631d},
  {32'hc46039b5, 32'hc4e41bc4, 32'h42830750},
  {32'hc4078560, 32'h443856ce, 32'h43e58c9f},
  {32'hc311483c, 32'hc46c12c3, 32'hc494d1c1},
  {32'hc4844145, 32'h439196c3, 32'h445e879c},
  {32'h44511b52, 32'hc4b2d590, 32'hc4b49ec0},
  {32'hc51f4214, 32'h42e92eb2, 32'h4422bf44},
  {32'h45139ec9, 32'hc342d0b0, 32'hc30fee99},
  {32'h440eb87d, 32'h452efecf, 32'hc2a86b2f},
  {32'hc348d472, 32'hc3c964e7, 32'hc49fd958},
  {32'hc3d13de4, 32'h44b3798e, 32'hc3137bda},
  {32'h444f4a02, 32'hc34dd573, 32'hc4a61b12},
  {32'hc49c183d, 32'h44a3dbf1, 32'hc30cfaf3},
  {32'hc4959674, 32'h43264621, 32'hc2a80dd8},
  {32'hc2763a64, 32'h44970c35, 32'h45613126},
  {32'hc2851fe0, 32'hc4c11e59, 32'hc4b291e8},
  {32'hc51bdc28, 32'hc31f3575, 32'h4380407b},
  {32'h4492b396, 32'hc4a24444, 32'h43468ae3},
  {32'hc52008a8, 32'h44157b72, 32'hc3b5c65e},
  {32'h4489ddc9, 32'hc3a99ab2, 32'h43e9cbe9},
  {32'hc50ee7ba, 32'h4432c88a, 32'hc20d7982},
  {32'h44c15abe, 32'h42aa6728, 32'h431ee0fc},
  {32'hc535d83c, 32'h42c7ecf9, 32'h433aab28},
  {32'h451e6440, 32'hc307fc3e, 32'h43aa11ac},
  {32'hc489913a, 32'h42b1151f, 32'h4405c851},
  {32'h43ce1ca1, 32'h41cf085f, 32'hc3cf9893},
  {32'h44bf803b, 32'hc347e082, 32'h446d0251},
  {32'hc501b062, 32'hc2b59278, 32'hc1abd0ae},
  {32'hc38b5910, 32'h442818b5, 32'h43847361},
  {32'h42a36a38, 32'h44ee1a06, 32'hc3198460},
  {32'h4563e764, 32'hc313d8dc, 32'hc2187ffc},
  {32'hc423e4d3, 32'h44c9dc21, 32'h43243a28},
  {32'h44029204, 32'h430adc79, 32'hc3b9c19f},
  {32'hc388caf5, 32'h4528cc45, 32'hc20887c5},
  {32'h4473d7ec, 32'hc460e3a3, 32'h43c1a8c8},
  {32'hc32c1b29, 32'hc3cef172, 32'hc4d1a765},
  {32'h43dda16d, 32'h43961d22, 32'h44374974},
  {32'hc47c7470, 32'h43351ace, 32'hc4e39327},
  {32'hc4f358ca, 32'h43d7ffcb, 32'h438a2757},
  {32'hc31501b8, 32'h43c2eec1, 32'h44cf8b68},
  {32'h43352b3e, 32'hc3acd6a9, 32'hc51b1988},
  {32'hc2b3d8e8, 32'h42c875ec, 32'h44bf086a},
  {32'h43bc6771, 32'hc51e878a, 32'h42efb10a},
  {32'hc2bc2eaf, 32'hc3b05b40, 32'h450bf222},
  {32'h448e2a7b, 32'hc3cec20f, 32'hc36f549a},
  {32'hc4e242b3, 32'hc3c6fa20, 32'h43930d26},
  {32'h454b0032, 32'h43b611ed, 32'hc40af305},
  {32'hc4632ca7, 32'h440a36aa, 32'hc22bf41d},
  {32'h453f1c54, 32'hc41806b4, 32'h42e0193d},
  {32'hc453611b, 32'h4444c6ab, 32'h45047c52},
  {32'h41501701, 32'hc50668c6, 32'hc4341b72},
  {32'hc54670f2, 32'h43056e3a, 32'hc3c50017},
  {32'h440dd16b, 32'hc4b58ef9, 32'hc4c369c0},
  {32'h453a10e2, 32'hc3fabab1, 32'hc3cda1a5},
  {32'hc4d5548b, 32'h41e04d4c, 32'h448d4db9},
  {32'h44ff52ce, 32'h44099748, 32'hc2903b9c},
  {32'hc1e4bc88, 32'hc53c0afb, 32'hc40579f6},
  {32'h44992a20, 32'h42e3936a, 32'hc2546e95},
  {32'hc3d3a67c, 32'hc4a97543, 32'h44174dd4},
  {32'h452ba798, 32'h4472c812, 32'h43353b8d},
  {32'hc4dc5c5e, 32'hc493b656, 32'h41ac99d6},
  {32'h43113d24, 32'h44b26599, 32'h42247c4d},
  {32'hc4117700, 32'hc37deb67, 32'hc318be57},
  {32'h44911fc8, 32'hc38532e2, 32'hc401d59c},
  {32'hc4edd87e, 32'hc3e3f575, 32'h4316f938},
  {32'h4427c68c, 32'h455f9a13, 32'h434bf12e},
  {32'hc3c8d3ae, 32'hc5120e51, 32'hc49963b4},
  {32'hc36afafe, 32'h44a7b990, 32'hc2527464},
  {32'hc4370fee, 32'hc3245e42, 32'hc51e8611},
  {32'h43a8290c, 32'h44ff3d84, 32'h43a8bb42},
  {32'hc3dbcb85, 32'hc4ae2492, 32'hc2950668},
  {32'h4448545b, 32'h439f34b8, 32'h4489bc63},
  {32'hc5053836, 32'h438f4ea4, 32'hc317bf23},
  {32'hc40eb730, 32'hc33b21fc, 32'h435628d6},
  {32'h42b569fa, 32'h430f71d4, 32'hc534f163},
  {32'h448df574, 32'h43eb505b, 32'h42fbe9e4},
  {32'h44e5eca9, 32'h42274f8f, 32'h4359fe86},
  {32'h4373e653, 32'h449bc59d, 32'h450b7a7a},
  {32'hc441c27d, 32'hc4b77cf3, 32'hc42eefc1},
  {32'h427d0020, 32'hc3505753, 32'h44cac81a},
  {32'h446d2ce3, 32'h4375e7c9, 32'hc3e2e18a},
  {32'h435807ac, 32'hc51be667, 32'h43bcccbf},
  {32'h4198ec60, 32'h4531360b, 32'h41bd7495},
  {32'hc37faf00, 32'hc3c1ee15, 32'h43c35a8b},
  {32'h43fbb109, 32'h44f00129, 32'hc399fba6},
  {32'hc52fb951, 32'hc4280b29, 32'h406b8740},
  {32'hc434aec1, 32'hc310223b, 32'h433461ae},
  {32'hc508cc5c, 32'h42e667e8, 32'hc3524555},
  {32'h449f9d77, 32'h43d637e0, 32'h43f5235b},
  {32'h43ec9b3e, 32'hc42f9c4f, 32'h43e8066f},
  {32'h4516d749, 32'h433be97c, 32'h42880fc8},
  {32'hc417c093, 32'hc33b7ef0, 32'h43dd4180},
  {32'hc4121e24, 32'h44b71d1b, 32'hc356fc1f},
  {32'hc426682c, 32'hc494b224, 32'h44419a50},
  {32'h44104540, 32'h44dcde06, 32'hc41ed86f},
  {32'h438044a8, 32'hc3e1da1c, 32'hc397f450},
  {32'h43af42a5, 32'h43b450f1, 32'hc5092a80},
  {32'hc50068a8, 32'h4343f6aa, 32'h43df13d6},
  {32'h44e9ed82, 32'hc3648ef6, 32'hc370cf87},
  {32'hc4638934, 32'hc51d9a64, 32'h44271750},
  {32'h4451d21d, 32'h447d891e, 32'hc2cff0a4},
  {32'h43d8b3d4, 32'hc51846bf, 32'h41b88473},
  {32'h43f6475c, 32'h44a42421, 32'hc402484e},
  {32'h423de5e0, 32'hc3c0707d, 32'h4513c296},
  {32'hc4348118, 32'hc3c30657, 32'hc491cce6},
  {32'hc58623bb, 32'h43291b27, 32'h412c9f59},
  {32'h44430eca, 32'hc32aa732, 32'hc4a1e31f},
  {32'h43cca692, 32'hc4f901c5, 32'hc3a34533},
  {32'hc3d3488c, 32'h44d922f3, 32'h43e1e5d2},
  {32'h43b007f4, 32'hc51f243b, 32'hc29e2a24},
  {32'hc2d0a423, 32'h450eba3a, 32'hc37a0358},
  {32'hc2e87ee0, 32'hc4bd9d1c, 32'hc3fb501b},
  {32'hc41c5948, 32'hc3297cb1, 32'hc2685268},
  {32'h45691c7b, 32'hc254d887, 32'hc3d51e30},
  {32'hc42ca7f7, 32'hc3dcc1db, 32'h440457b0},
  {32'hc3fb9328, 32'h431fd0fa, 32'h433b5c34},
  {32'hc41ca357, 32'h444f2590, 32'hc499ee14},
  {32'h44562838, 32'hc3b8d94b, 32'h43a94ce5},
  {32'hc3817f2e, 32'h44848aa2, 32'h43a14d13},
  {32'h454a4e39, 32'hc3ceb5b4, 32'hc225fcc2},
  {32'h43a3cf4c, 32'hc29a08d5, 32'hc3b4f8fe},
  {32'h45017047, 32'hc2be7d42, 32'h43af1750},
  {32'hc49fe5ae, 32'h43d8d17d, 32'hc41a80fe},
  {32'h44de6c34, 32'hc32cd9a9, 32'h444f7d57},
  {32'hc524573e, 32'hc267b0e8, 32'h433fe53b},
  {32'h42dffa40, 32'hc4a176c0, 32'h44e0900f},
  {32'hc410be1a, 32'h44ac327e, 32'hc4c4969b},
  {32'h452a5bcf, 32'h432e7279, 32'hc376294c},
  {32'hc3d90777, 32'h42d0713a, 32'hc52595c9},
  {32'hc31e09a8, 32'hc47d5c88, 32'h44168ed6},
  {32'h44798548, 32'hc2533ba8, 32'hc44dd067},
  {32'h4392a988, 32'h430b0e46, 32'h44327712},
  {32'hc48249d5, 32'hc3f2225a, 32'hc507e82c},
  {32'h426ff1de, 32'hc2bd3083, 32'h445f8885},
  {32'hc4b2fe92, 32'h42cf49d9, 32'hc3f95f28},
  {32'hc497b373, 32'h43d15422, 32'hc2aa9b71},
  {32'h42395c2a, 32'hc41e11d7, 32'hc4bd4750},
  {32'hc31027b3, 32'h43a0531e, 32'hc2adc1e7},
  {32'h45030c1a, 32'hc375689c, 32'h449f6e3d},
  {32'hc398430c, 32'h41dacf29, 32'hc4686481},
  {32'h421241f4, 32'hc4c18263, 32'hc3c6e97c},
  {32'hc35a6983, 32'h455d8d4f, 32'h42c7c502},
  {32'hc32c8073, 32'hc56f919b, 32'hc1f1c989},
  {32'h440474f8, 32'hc48d3a8d, 32'h4546091a},
  {32'hc4adf726, 32'hc4636d44, 32'hc3930b5a},
  {32'h4506ef55, 32'h40eab610, 32'hc401d0cc},
  {32'h44c83ea1, 32'h42e9c875, 32'h42f5efdb},
  {32'hc4233400, 32'h43ee405a, 32'hc3adc713},
  {32'hc30b1c02, 32'hc4e617a6, 32'hc3383705},
  {32'hc21ff2a4, 32'h44c98d6e, 32'hc3915def},
  {32'h44da04f8, 32'hc31f7206, 32'h445ba056},
  {32'hc3d37716, 32'h44766092, 32'hc49b09e3},
  {32'h45547561, 32'hc3a23c04, 32'h438467bd},
  {32'hc4ce6215, 32'hc285c64a, 32'hc2a2a67b},
  {32'h457033bc, 32'h43bc88c1, 32'h41aac8f8},
  {32'hc4c01a3a, 32'hc2ecf00b, 32'hc23cdea0},
  {32'h41ec0020, 32'hc572db1f, 32'hc380506d},
  {32'hc4c75a58, 32'h4485c2fa, 32'hc3c8355d},
  {32'h453bafd8, 32'h43b906ac, 32'h426a934b},
  {32'hc3928020, 32'h4580c6fa, 32'hc3dd56cb},
  {32'hc4048772, 32'hc588e34e, 32'hc232086f},
  {32'h44093113, 32'hc4be36c9, 32'h43ee710c},
  {32'h41c4ef90, 32'h43b93526, 32'hc519186f},
  {32'hc5271cb1, 32'h43cac130, 32'h4339944e},
  {32'hc43485b9, 32'hc4ae73b8, 32'h44336663},
  {32'hc2ddd74c, 32'h41e3d82b, 32'hc4f6f5de},
  {32'h44f0c812, 32'hc23bd788, 32'h43921b56},
  {32'h4298d698, 32'h449d0ddb, 32'hc41dbb73},
  {32'h4267bd80, 32'hc488b599, 32'h44a01349},
  {32'hc3907998, 32'h44135835, 32'h43a69ca2},
  {32'h4440616a, 32'h441d2272, 32'hc33287e3},
  {32'hc473e256, 32'h437cc1c3, 32'h4486dc1b},
  {32'hc12e60a0, 32'h44eabbce, 32'hc49bfb27},
  {32'hc2866fe8, 32'h44e1d6b1, 32'h43ee2f7e},
  {32'hc4b55270, 32'hc3be927c, 32'h427d4494},
  {32'h4400d4c9, 32'h41af8b4b, 32'hc4bf502e},
  {32'h42b87719, 32'hc4a09ef8, 32'h42495cb4},
  {32'hc311f8e6, 32'h44e6e586, 32'hc38eb2aa},
  {32'hc3ffad50, 32'hc44681ea, 32'h43d24d0d},
  {32'h44d1c778, 32'h4366966d, 32'h428e7a9a},
  {32'hc5992bb8, 32'hc2ba5a32, 32'h434d10bd},
  {32'h4511bcb6, 32'h43ebe721, 32'hc371f826},
  {32'hc4773911, 32'hc4bdd630, 32'hc1ebef1a},
  {32'h458599c4, 32'h43ba1a6d, 32'h437ee925},
  {32'hc451f8e0, 32'hc3adacdc, 32'hc1d9a27f},
  {32'h4562d00b, 32'h441be5fb, 32'h434ab2ba},
  {32'hc3e028cc, 32'hc4f0874d, 32'h40e8940b},
  {32'hc4492820, 32'hc3296687, 32'hc4115187},
  {32'h43f3ba39, 32'hc4de59f2, 32'h43e0e698},
  {32'hc44c0a80, 32'hc380e2af, 32'hc4910a30},
  {32'h4421e70f, 32'hc4c578b5, 32'h4499af64},
  {32'hc2c7b93f, 32'hc2a4bd92, 32'hc4bae769},
  {32'h445c510d, 32'hc2854a91, 32'h44dff7e1},
  {32'hc50d9edb, 32'hc45b3584, 32'h42240a46},
  {32'h449e7bae, 32'h447a3c1c, 32'h436598b3},
  {32'hc3da7ffc, 32'hc50a0fa5, 32'hc4b0f8cb},
  {32'h436e926a, 32'h4405daee, 32'h454637d5},
  {32'hc43a2448, 32'h44230e08, 32'h434b29f5},
  {32'hc492ef60, 32'hc4ca537b, 32'h44ef30a5},
  {32'hc3960d36, 32'hc48e3c6d, 32'hc4588e5b},
  {32'hc438d656, 32'h4366d782, 32'hc3b97aa2},
  {32'hc51c409c, 32'hc39f0271, 32'h41ae1338},
  {32'h447e05b4, 32'h431c6b8f, 32'h41e0e937},
  {32'h4481532b, 32'hc4681fd9, 32'hc396da4c},
  {32'h451556b6, 32'h43bd4f0f, 32'h439c2e30},
  {32'h43e8d74b, 32'hc4dae1a9, 32'hc4a08800},
  {32'hc3b66e88, 32'h4439ed0b, 32'h4391d9dc},
  {32'hc4427e8d, 32'hc51efd6c, 32'hc39b6d5b},
  {32'h451d748c, 32'h44502d4a, 32'hc439627c},
  {32'hc3e73967, 32'hc35ba602, 32'hc41b5e88},
  {32'h43008bd8, 32'h45522955, 32'hc2557869},
  {32'hc4207a4f, 32'hc4b22c12, 32'h432a5a90},
  {32'h454ced43, 32'h42b2e3ae, 32'h439748d4},
  {32'hc54564ba, 32'h43dd4574, 32'hc42b5dfa},
  {32'h4471166c, 32'hc41819ce, 32'h431aa274},
  {32'h44a9fdf9, 32'h4405dccf, 32'hc4b034f2},
  {32'hc3164410, 32'h4495a56d, 32'h443c4c88},
  {32'h439fdb88, 32'h43495891, 32'hc483b64f},
  {32'hc3b8eda8, 32'h43a24077, 32'h43894110},
  {32'h43d348de, 32'hc5072af0, 32'h437ebffc},
  {32'h42ad96f2, 32'h44b69c08, 32'h441c4bff},
  {32'h44feb97e, 32'hc42ee0dd, 32'hc48164a1},
  {32'hc467bd58, 32'h445cecac, 32'h449dd487},
  {32'hc31586e0, 32'hc43564f1, 32'hc50415c0},
  {32'h4188e3d9, 32'h45013158, 32'hc32edc87},
  {32'hc40994fb, 32'hc4c9b835, 32'hc42297a5},
  {32'hc2ac5aaf, 32'h4483ed56, 32'hc0d56473},
  {32'h449d5ffb, 32'h432fe1b2, 32'hc418e191},
  {32'hc44c2474, 32'h43ee522d, 32'h44e24678},
  {32'hc2ca6129, 32'hc48d9ea3, 32'hc36c4ca1},
  {32'hc3f7ac56, 32'h448dc852, 32'h44fb3bb9},
  {32'h4410b5b6, 32'hc4e2eea2, 32'hc45edd48},
  {32'hc4e12765, 32'h4221e0b2, 32'h428b5bc3},
  {32'h442e4948, 32'hc534b17c, 32'hc3ee8e45},
  {32'hc565c652, 32'h4408a0f9, 32'hc3c6b499},
  {32'h4218b2c4, 32'hc4eb8a43, 32'h428bf74d},
  {32'hc380aec8, 32'h451e6d83, 32'hc3ddfe29},
  {32'h4498ffc0, 32'hc48f3e5d, 32'h41f0d839},
  {32'h440ae2a2, 32'h448c460e, 32'h439eb8b0},
  {32'h44a03d4a, 32'h43afc54b, 32'hc3149fcf},
  {32'hc4bf7824, 32'h43dba0cc, 32'hc36bf94e},
  {32'hc34a0a39, 32'hc3f5e78d, 32'hc3f56dd2},
  {32'h4340957a, 32'hc3818cb2, 32'h4451e5d8},
  {32'hc56b59a8, 32'h41ca4ec4, 32'h439ec224},
  {32'h4553fbdf, 32'h427e0673, 32'h43f7cd6d},
  {32'hc5574284, 32'hc2cc1108, 32'hc424e6d5},
  {32'h452ac3d3, 32'hc366e4c6, 32'h42f149ca},
  {32'hc527479a, 32'h43c3cbb3, 32'h437f8c13},
  {32'hc4184d53, 32'hc350a600, 32'h438d66d4},
  {32'hc56961ec, 32'h43b53666, 32'h42fcf6b9},
  {32'h43dde7f0, 32'hc52c3649, 32'hc1c7b856},
  {32'h447d4e86, 32'hc38047d1, 32'hc389b491},
  {32'h4482b696, 32'h434c121d, 32'h44438fbc},
  {32'hc4659d19, 32'h43c9bc63, 32'hc3e2be44},
  {32'h430492b8, 32'hc4a1e574, 32'hc316d10f},
  {32'h43027080, 32'hc1a23935, 32'h44e9044e},
  {32'h43f18dfc, 32'hc4d83002, 32'hc4545f83},
  {32'h44db213f, 32'hc3ac9d37, 32'h4380c6b7},
  {32'h44e4291a, 32'hc3c006ca, 32'h4203b064},
  {32'hc2d6701b, 32'hc2d47e5c, 32'h44b332bf},
  {32'hc49ba19b, 32'hc2a11967, 32'hc409d54f},
  {32'hc4fbd6ee, 32'hc49397e4, 32'h43ac6e36},
  {32'hc38f7838, 32'h4496cefd, 32'hc43ae322},
  {32'hc37f3fff, 32'hc35a8d84, 32'h42188b1c},
  {32'hc3b171a0, 32'hc4f96d9d, 32'hc33a14f1},
  {32'hc4a7b4e3, 32'h4414ac75, 32'h3fae26dc},
  {32'h42b5a2f0, 32'hc457ad38, 32'h438c125f},
  {32'h420b5a60, 32'h44b1908d, 32'h44f76775},
  {32'h4409a1d0, 32'hc424b32d, 32'hc500b220},
  {32'h44e05d89, 32'h41ee2e92, 32'hc45e98f0},
  {32'hc4aa1cf7, 32'h432af4db, 32'h42ec8760},
  {32'h44d905cd, 32'hc43061ab, 32'h42896468},
  {32'hc42997ac, 32'hc4e6aca6, 32'hc41b7654},
  {32'h4419fa75, 32'h44986308, 32'h43ac54d2},
  {32'h44c37600, 32'hc3087f7c, 32'hc22da2cd},
  {32'h44d46b2c, 32'h44e01bf7, 32'h43d0adb1},
  {32'hc5973ca8, 32'hc327ff44, 32'h42acb10a},
  {32'h4414804f, 32'h44422070, 32'h43ac0d62},
  {32'hc1fb7f80, 32'hc41e7f32, 32'h4337a8fc},
  {32'h43e631a8, 32'h43cad8df, 32'hc45e318e},
  {32'h4513efe9, 32'hc38530df, 32'h43576e26},
  {32'h44fee388, 32'hc23386c9, 32'hc0e55cf8},
  {32'hc4061ea4, 32'hc41b2258, 32'hc4a6a5c7},
  {32'hc3d4fedd, 32'h44d1e926, 32'h43b9bc36},
  {32'hc44cdf92, 32'hc4e5edbd, 32'hc35ebf7a},
  {32'h4401c1c7, 32'h4403988d, 32'h44f8605f},
  {32'hc51a49ce, 32'hc35535f6, 32'h43801e9a},
  {32'h43e12e7c, 32'hc41de501, 32'h44bade2f},
  {32'hc425918e, 32'hc392daf7, 32'hc3d4fd30},
  {32'h44f573a8, 32'h4263bab4, 32'hc3a21bc5},
  {32'hc4cf4e6e, 32'h43a5900b, 32'hc2a87a55},
  {32'hc3d64271, 32'h43ce9aa4, 32'h4481bdb6},
  {32'h43e6ebab, 32'hc4957f99, 32'hc3472df4},
  {32'hc41d7478, 32'h44dc2c24, 32'hc1904298},
  {32'hc2c2fb40, 32'hc4da8a38, 32'hc2ce7280},
  {32'hc4696001, 32'hc292d02f, 32'h441556fe},
  {32'hc31343ee, 32'hc42d78a6, 32'h43b1fad3},
  {32'hc2e55d94, 32'hc5708695, 32'hc3afa9f8},
  {32'h43b32544, 32'h4469e7c2, 32'h443dab7b},
  {32'hc2b81d83, 32'hc3be63af, 32'h4312be46},
  {32'h41c95820, 32'h453c9423, 32'hc3be10cb},
  {32'hc40e0060, 32'hc545f1ae, 32'h42e0ba1b},
  {32'hc388bb84, 32'h418ec03c, 32'hc3ca2fb3},
  {32'hc4edbcb6, 32'hc48af67e, 32'hc3e3c785},
  {32'h44068358, 32'h43ab950a, 32'hc3a71d01},
  {32'hc4d201fc, 32'h4206f4a4, 32'hc385bbe8},
  {32'h4400548f, 32'h44c044f3, 32'h42075b14},
  {32'hc46a1f7d, 32'hc3c7615b, 32'hc3a7dedf},
  {32'hc4bd3680, 32'h43a8731f, 32'h43071d74},
  {32'hc403aba4, 32'hc46b1f93, 32'h43ba01a7},
  {32'h43c29ad2, 32'h44e91fea, 32'hc39228ec},
  {32'h44802dc8, 32'hc388afd2, 32'h4291af3c},
  {32'h43a493d6, 32'h42884a5d, 32'hc418f71d},
  {32'hc3d63490, 32'h438c96f4, 32'h432c8261},
  {32'h43ded2de, 32'h444c339f, 32'hc3847bfb},
  {32'hc4e18977, 32'hc4756ed8, 32'h43ba1c9e},
  {32'h43deb238, 32'h448f5f40, 32'hc5003cea},
  {32'h4399e064, 32'hc28080f6, 32'h44726b87},
  {32'h43a41164, 32'hc29e0968, 32'hc4882c02},
  {32'hc4855f90, 32'hc3c96c6e, 32'h4421ca84},
  {32'h42c8fdc7, 32'hc3eb9cc9, 32'hc4baf197},
  {32'hc54522cf, 32'h4309a795, 32'h445a1302},
  {32'h4493f552, 32'hc31350a9, 32'hc42b5327},
  {32'h43e88aa2, 32'hc496fb21, 32'h41fa2741},
  {32'hc4ab7afc, 32'h446fc1b1, 32'h428b1a5a},
  {32'h4408b07e, 32'hc3cd9942, 32'h43f9b8c2},
  {32'hc517a74c, 32'h440c5a6e, 32'h43c5921d},
  {32'h4543bd55, 32'h42fb8a72, 32'h436bf7bc},
  {32'h438868c2, 32'h44965ad8, 32'hc28d4039},
  {32'hc3098940, 32'h44295602, 32'h42d0739e},
  {32'hc557cf9e, 32'h43a645fe, 32'h43cdc573},
  {32'h4504b690, 32'h431d2169, 32'h43a7c5ed},
  {32'h435299ae, 32'h43f8ad20, 32'h4406ed1b},
  {32'hc3e600c1, 32'hc45c5cdd, 32'hc21ce7f0},
  {32'hc34e2f58, 32'h43baa9b1, 32'h4390c243},
  {32'h43a11969, 32'hc48b8585, 32'h449b9018},
  {32'hc511fe40, 32'h441da03c, 32'hc35d8cfb},
  {32'hc4454635, 32'h431bc8e0, 32'h43de3e92},
  {32'hc45ac3be, 32'hc374eed9, 32'hc2a31128},
  {32'h44118059, 32'hc3a9ba5f, 32'h418065f0},
  {32'h428ff28f, 32'h422b3f0e, 32'hc45e63e9},
  {32'h44a1bd50, 32'hc4ea8580, 32'hc3a97e1e},
  {32'hc40855d3, 32'h449bb6ad, 32'hc38984af},
  {32'hc4cd9ad0, 32'h42068a37, 32'hc3ba4504},
  {32'hc47d1792, 32'hc276ba5f, 32'hc4da59f3},
  {32'h449c5917, 32'hc3b4251a, 32'hc34ed3d3},
  {32'h43abdcae, 32'h44f9c378, 32'hc38d00b6},
  {32'h447ae495, 32'h443193f7, 32'h45368b8b},
  {32'hc56b84f8, 32'hc395e0a2, 32'hc32b686d},
  {32'h45130c88, 32'hc3b3dac0, 32'h43a3957e},
  {32'h438cb89d, 32'h44361264, 32'hc5489a5c},
  {32'h43aeda64, 32'h42ff8dda, 32'h451f354a},
  {32'h43899ecb, 32'h441f601a, 32'h431e2f5f},
  {32'hc52a59c0, 32'h43bdedd2, 32'h42a4249a},
  {32'h4314c38c, 32'hc39ff4f6, 32'h44a2bd9f},
  {32'hc43972e4, 32'h44431115, 32'hc4435559},
  {32'h449ef331, 32'hc39caf54, 32'hc387cd7b},
  {32'hc48f8ecd, 32'h44a45397, 32'hc384b580},
  {32'h4312b327, 32'hc48edd5c, 32'h449241e7},
  {32'h414533ca, 32'hc401d262, 32'h450c3299},
  {32'hc50b390d, 32'hc3518b73, 32'hc3e905d2},
  {32'h44d57659, 32'h43ac7de9, 32'hc46f2c32},
  {32'h44741b1e, 32'hc2f2f9ee, 32'hc25f96d9},
  {32'hc44309c0, 32'h43d13259, 32'hc4101b82},
  {32'h4326be82, 32'hc51d70db, 32'hc3c5290b},
  {32'h43b48854, 32'h44e0a428, 32'h4348ed89},
  {32'h41c9ca88, 32'hc52f5b47, 32'hc310a9a0},
  {32'hc4e6c257, 32'h43c11ebb, 32'hc4104a62},
  {32'h451d868b, 32'hc1d005a5, 32'h437a2331},
  {32'hc53eef20, 32'hc08702dc, 32'hc3d4fcbd},
  {32'h456b6816, 32'h42f50fab, 32'h433e952e},
  {32'hc23e40d6, 32'h44d0eb8e, 32'h43f4c099},
  {32'h45734f3f, 32'h43c69862, 32'h4268ca41},
  {32'hc3858394, 32'h44848fc7, 32'h4338ef33},
  {32'h430ed362, 32'hc4b8b121, 32'h43835d33},
  {32'h43dd08bf, 32'h45576225, 32'h433c47d7},
  {32'h4555ce85, 32'hc40d77e3, 32'hc2f0eb46},
  {32'hc4db48ef, 32'h424023c6, 32'hc332fe6f},
  {32'hc4107cb6, 32'h4406653d, 32'hc537d80f},
  {32'hc484db5d, 32'hc40252d8, 32'h442e3639},
  {32'h428bf4f8, 32'h4215a3ed, 32'h452a8ed3},
  {32'h4411f03b, 32'h447a6638, 32'hc4957e57},
  {32'h44cbc37f, 32'hc1adfb4b, 32'h43993308},
  {32'hc33813d5, 32'hc19432f7, 32'hc56f6d76},
  {32'hc4bcf050, 32'hc4886f8a, 32'h43866555},
  {32'h4341275f, 32'hc32fc9ea, 32'hc4316b75},
  {32'h44240628, 32'hc443b435, 32'hc31bd3e0},
  {32'h43c2a000, 32'h415e431d, 32'h44c83736},
  {32'h40f49e00, 32'hc46112cd, 32'hc4f8beb4},
  {32'h44336f75, 32'h43ce71bf, 32'hc49dfa02},
  {32'hc3872aa2, 32'hc51b3e8d, 32'hc39da336},
  {32'hc49300c5, 32'h43aceb8e, 32'hc2db45c2},
  {32'hc4775ab4, 32'hc4731670, 32'h42b10899},
  {32'h44a6aee1, 32'h4362d137, 32'hc4052cf7},
  {32'hc484979b, 32'hc42b974a, 32'h40f523cc},
  {32'h44b9848a, 32'hc42de960, 32'hc3cb0414},
  {32'hc534e3bb, 32'h432d0260, 32'h4443a372},
  {32'hc48dc4bb, 32'h43b568ec, 32'hc30b7b02},
  {32'hc549644e, 32'hc4502aeb, 32'h430c3da2},
  {32'h451a022e, 32'h4439d2ce, 32'h436a5fb8},
  {32'h44932128, 32'h42866d68, 32'hc2db9bed},
  {32'h454d8e72, 32'h43de3e8f, 32'h42b9d52c},
  {32'hc4079b5c, 32'hc4d7a064, 32'h4341ae74},
  {32'h44664716, 32'hc33d5e87, 32'hc44ce16f},
  {32'hc4b69330, 32'h4385fa9b, 32'h435a9c9a},
  {32'hc497173c, 32'hc425b672, 32'hc2db039b},
  {32'h43bb107c, 32'h45009caa, 32'h4406f4ed},
  {32'h4390e713, 32'hc3a67c63, 32'hc4925208},
  {32'h42588a86, 32'h453702d4, 32'h439ebe88},
  {32'hc474a100, 32'hc44e1556, 32'hc3e99816},
  {32'h423e2bb8, 32'h43f63be6, 32'h4397ccca},
  {32'hc434b463, 32'hc3899fbd, 32'hc3b9823a},
  {32'h4415eb33, 32'h432c0311, 32'h44f63a54},
  {32'h431d588d, 32'hc3f230bc, 32'hc3baf36b},
  {32'hc4545830, 32'hc46b1ae1, 32'h45072ae9},
  {32'hc395eff5, 32'hc34b4ca1, 32'hc4b42312},
  {32'h44c81611, 32'h440752bf, 32'h43239757},
  {32'hc3be5614, 32'hc4ec23f0, 32'hc29cb501},
  {32'h44b05652, 32'h4401365a, 32'h43a29e54},
  {32'hc4ce55a4, 32'hc3f3f69a, 32'hc34c4cf7},
  {32'hc34911d7, 32'h449a91dd, 32'h450efc5a},
  {32'hc0e9f480, 32'h41f53348, 32'hc4b8a37e},
  {32'h450e4c69, 32'h4246889e, 32'h4220d986},
  {32'hc41c05ff, 32'hc54f736a, 32'h43ce27b2},
  {32'h440be024, 32'h44e31fa5, 32'h428c14ef},
  {32'h43dbe980, 32'hc2404394, 32'hc35c276f},
  {32'h43b5c5ae, 32'h4512ed1a, 32'hc0ba0e94},
  {32'hc2da28a0, 32'hc4a4d159, 32'hc303c296},
  {32'hc4cc59a1, 32'h41b6f99c, 32'hc42b1d5b},
  {32'hc58ab403, 32'h40a51808, 32'hc38a038a},
  {32'h457da074, 32'hc3b1dd87, 32'h43222d60},
  {32'h43a447ca, 32'hc3d18dfa, 32'hc3d4058b},
  {32'hc367507c, 32'hc4f9f496, 32'h44dfdcd8},
  {32'hc400b310, 32'h43988064, 32'hc45e49e9},
  {32'hc38df6cc, 32'h4424ad54, 32'h44ce30c6},
  {32'h44cb8eb4, 32'hc2d547e4, 32'hc446b523},
  {32'hc2ce9f8c, 32'h44e3be7c, 32'h43a51cb7},
  {32'hc4011596, 32'hc3ec08ff, 32'hc42cf6d6},
  {32'hc4f115de, 32'h43060f59, 32'h446548d4},
  {32'hc35b2c1f, 32'hc4b80a90, 32'hc467ad70},
  {32'hc4e08a46, 32'h43b9ed3f, 32'h4385621b},
  {32'hc3e81e58, 32'h44989342, 32'hc51df00f},
  {32'hc4b61f38, 32'h43c1dfe0, 32'hbfb4b428},
  {32'h4449c9c8, 32'hc3bd944e, 32'hc469ca59},
  {32'hc412b360, 32'h444dde3a, 32'h442ee651},
  {32'h440f1757, 32'hc3624e2b, 32'hc4e9dc6e},
  {32'hc445b5cc, 32'h43ea8acb, 32'h44c59527},
  {32'h42cfa870, 32'hc4b3e064, 32'hc45d4b09},
  {32'hc3f8f024, 32'hc375811b, 32'h4485f890},
  {32'h44b7ac0e, 32'hc4ba7708, 32'hc2d64a1e},
  {32'hc4cd5188, 32'h44bb58ce, 32'h436d6822},
  {32'hc48a7bcb, 32'hc29e1c55, 32'hc358d85a},
  {32'h427701b0, 32'h44894153, 32'h4323f2e4},
  {32'h4445167c, 32'hc4a24d48, 32'hc27f134e},
  {32'hc42abc16, 32'h44382910, 32'hc16bde05},
  {32'h443f35a8, 32'h408654f0, 32'hc40f8305},
  {32'hc3edae80, 32'hc180fc06, 32'hc3079c7c},
  {32'h452d5f30, 32'hc3016979, 32'hc3ab1118},
  {32'h4493f8c3, 32'hc3580bc8, 32'h44980435},
  {32'hc56aa58c, 32'h431df5bf, 32'h43ae33e9},
  {32'h44a82477, 32'h43edc9e2, 32'h44b91584},
  {32'hc3dc72fe, 32'hc33e876e, 32'h424823e2},
  {32'h4493f61c, 32'hc477fa63, 32'h43b7bfeb},
  {32'hc480d29a, 32'h44c9436d, 32'h42db7654},
  {32'h447f0294, 32'hc4063f79, 32'h43747568},
  {32'hc46408d4, 32'h451297dd, 32'hc315b4e6},
  {32'h4518c510, 32'h4237fe83, 32'h43b2386f},
  {32'h45001dcb, 32'h4385a6fb, 32'h42d41769},
  {32'h4431535c, 32'hc4753158, 32'h45168ab4},
  {32'hc471ea16, 32'h43ec2c91, 32'h4340a633},
  {32'h44f3c464, 32'hc3395fbc, 32'h40767150},
  {32'hc32ed62c, 32'h435b6644, 32'h44e29fc6},
  {32'h437a54d4, 32'hc52f1b13, 32'hc3a26610},
  {32'h428ad6e8, 32'h43c26f3f, 32'h44536f8b},
  {32'h44f932f0, 32'hc4351d44, 32'hc417b5ee},
  {32'h420e63dc, 32'h44dde179, 32'hc1a01e6f},
  {32'h452f1fc6, 32'hc3d59017, 32'hc25fb8a1},
  {32'hc523ad66, 32'h4410df65, 32'h441924eb},
  {32'h4495add8, 32'hc40d8ec7, 32'hc46691d0},
  {32'h436cccab, 32'h4394243b, 32'h44bfc18a},
  {32'h43dca358, 32'hc4331755, 32'hc49eff1f},
  {32'hc37bd2a4, 32'h452be78b, 32'h4473bf7a},
  {32'h42d413a8, 32'hc31b9e1c, 32'hc3ad2d4c},
  {32'hc53246e1, 32'h441b1d22, 32'h42f672ce},
  {32'hc3ae58cc, 32'hc50e1b5c, 32'h42a6c884},
  {32'h443c5fe0, 32'h4496b903, 32'hc520ee03},
  {32'hc4075c3b, 32'h440fc91b, 32'h43883a01},
  {32'h44c05e4d, 32'h440402a1, 32'h437b99bf},
  {32'hc429557a, 32'hc45dae8a, 32'hc29b83ae},
  {32'h43f981d4, 32'h4485a98c, 32'hc32ff4ee},
  {32'h43ee30dc, 32'hc4b7708e, 32'h4369e5c0},
  {32'h44a8d0a8, 32'h449e79c5, 32'h431833d2},
  {32'hc4408dcb, 32'hc525f255, 32'hc3dd31fa},
  {32'hc4138e86, 32'h449726a6, 32'h433028c4},
  {32'hc4bc83ac, 32'h42355f68, 32'h44a64a7b},
  {32'h44968f20, 32'hc404233e, 32'hc3afbd7d},
  {32'hc4608aa8, 32'h441bd3db, 32'hc41b4107},
  {32'hc392b10e, 32'h444d064a, 32'h4391e786},
  {32'hc4ccf21c, 32'hc44fef09, 32'hc4af3fc0},
  {32'hc4937de7, 32'h43f187da, 32'hc2726cae},
  {32'hc5234204, 32'hc40c029b, 32'hc2b23f44},
  {32'h43db99af, 32'h4492c6ac, 32'h44891f99},
  {32'hc4bb8cbb, 32'hc36f2874, 32'h4431e1aa},
  {32'h42f8c5c0, 32'hc499a4bb, 32'h44e6c790},
  {32'hc560a4d6, 32'hc36d5b44, 32'hc39c39ba},
  {32'h4442acca, 32'h4412c45c, 32'hc32a0f5b},
  {32'hc3a1ace0, 32'hc40bffd1, 32'hc4d4b299},
  {32'h449cf2b6, 32'h42a91271, 32'h44820636},
  {32'hc480536e, 32'hc412bc65, 32'hc3d23882},
  {32'hc3244310, 32'h4522c54d, 32'h442362e0},
  {32'hc41f4838, 32'hc3f8ef1b, 32'hc4e7669b},
  {32'h43be4c42, 32'h44ae335b, 32'h43dff0df},
  {32'h4525b96d, 32'hc3bc8d8e, 32'hc403c9bc},
  {32'hc424db62, 32'h3ede2760, 32'hc4a64884},
  {32'h4453c40a, 32'h44b0e741, 32'h43f83de3},
  {32'hc5375f97, 32'h43ec3c4d, 32'h4297fc40},
  {32'h454d33c8, 32'h437bfcf4, 32'hc2856599},
  {32'hc4ce0de9, 32'hc447023e, 32'hc2116224},
  {32'h449b11c9, 32'hc006571c, 32'hc4305cbe},
  {32'hc4a5040c, 32'h4410d8c5, 32'hc32c1173},
  {32'h44d71b6c, 32'h4394a889, 32'h41ddc94d},
  {32'hc4ba048f, 32'hc2e19694, 32'h3fdb1e64},
  {32'h44197521, 32'h441cab82, 32'hc43022e3},
  {32'hc45d8a67, 32'hc3b97e9b, 32'hc1758ec7},
  {32'hc2c2717c, 32'h450018dc, 32'h433fedab},
  {32'hc53f03af, 32'hc2da9dc2, 32'h43966b30},
  {32'h441119cc, 32'h45494751, 32'h41784bdb},
  {32'hc41af862, 32'hc2577900, 32'h446fed39},
  {32'h44322ee2, 32'hc4889c06, 32'hc50c070a},
  {32'hc4e3d775, 32'hc44b8c0d, 32'hc38c8f75},
  {32'hc40e712f, 32'h43a57892, 32'hc1790ab8},
  {32'hc4588e0e, 32'hc4b29b6b, 32'h4480e189},
  {32'hc3b46700, 32'h4481c769, 32'hc308b43d},
  {32'hc4960fc3, 32'h41d29e1e, 32'hc39d51ef},
  {32'h42f90aec, 32'h4557e82a, 32'h41f8f45f},
  {32'hc44e2b7c, 32'h42cf3392, 32'h44ee9556},
  {32'h454304b9, 32'h43a1f58e, 32'h43f4c28f},
  {32'hc3fafe30, 32'h4364b848, 32'h4484faa9},
  {32'h44e323d6, 32'h43ab16e0, 32'hc4948cf6},
  {32'h44045548, 32'hc434ff3c, 32'hc439be42},
  {32'hc493e6e2, 32'h44b0ffea, 32'h431351bf},
  {32'h446d0121, 32'hc310c415, 32'hc2ae81c9},
  {32'h433f0d30, 32'h457df5c8, 32'h4337b779},
  {32'h4349f68e, 32'hc48c6460, 32'h42864c0f},
  {32'hc4cb3002, 32'hc35db683, 32'hc2b62d8e},
  {32'hc333b6bf, 32'hc38f6bdd, 32'hc419ac11},
  {32'hc4f77e3a, 32'h44016181, 32'h435e0e66},
  {32'h43a0f2ff, 32'h43e11b22, 32'h43b7ec89},
  {32'hc32ac3c2, 32'h448eba47, 32'hc20ad790},
  {32'h44406bb8, 32'hc403df7c, 32'h4494a145},
  {32'h43ab2027, 32'h4488d762, 32'hc487f56f},
  {32'h445dd073, 32'hc4bb7842, 32'hbf0d7427},
  {32'hc4d7b0fd, 32'hc28b7705, 32'hc445b5b2},
  {32'hc44ac74c, 32'hc1fd35fb, 32'h4412e0ea},
  {32'hc23df8c0, 32'h440f88f5, 32'h437dc774},
  {32'h45066301, 32'h436d58a0, 32'h433bc1a4},
  {32'h43b2b2de, 32'h4419fe98, 32'h43e2f989},
  {32'hc14f2a80, 32'hc4b1bf0d, 32'h4495a522},
  {32'hc4c9af81, 32'h43c1655c, 32'hc48aa93f},
  {32'hc44bfdde, 32'hc47755c6, 32'h4395527a},
  {32'hc48d524b, 32'h43254216, 32'hc4e1a849},
  {32'h44f2b12a, 32'hc40c4d0b, 32'hc3549ba2},
  {32'hc4a1faa7, 32'h43a5ef3c, 32'hc398f322},
  {32'h44d7e40c, 32'h44007737, 32'h44306e03},
  {32'hc4bc3960, 32'hc39d3c32, 32'hc341d27d},
  {32'hc4e7a53e, 32'h43934eb2, 32'h4366d14b},
  {32'h4366463c, 32'hc4428136, 32'hc44d6a68},
  {32'h452ca7bd, 32'hc3133c3b, 32'h4218ccec},
  {32'hc1c1fda8, 32'h448456f8, 32'hc45c4a27},
  {32'hc31f88a2, 32'h44ee4ffd, 32'hc2fe7be8},
  {32'h44c372c0, 32'hc43109bb, 32'h428e9d57},
  {32'hc4cbf5c3, 32'h43ca0fb0, 32'hc3e8962b},
  {32'h43cf0327, 32'hc168471d, 32'h44018233},
  {32'h435afdcc, 32'h44efc51e, 32'hc43391c4},
  {32'h448ccaac, 32'hc49d830a, 32'h442f3585},
  {32'h432df639, 32'h4363542d, 32'h44f60894},
  {32'h443c82ad, 32'h44a94369, 32'hc452db50},
  {32'hc31f9e51, 32'hc44749aa, 32'h447187b4},
  {32'h42de58a9, 32'h4182bebd, 32'h430ba453},
  {32'hc40ce264, 32'h44cbbc68, 32'hc3559418},
  {32'h44e6352a, 32'hc2ac6ce4, 32'h43c4ba28},
  {32'hc4fe8b84, 32'hc34dc822, 32'h42483c72},
  {32'hc3699ad8, 32'hc1c14665, 32'h44f4cb3c},
  {32'hc3938ff6, 32'h44d1cd8f, 32'hc3b83477},
  {32'hc4ddbd53, 32'hc3a50c35, 32'hc2315562},
  {32'hc50150b4, 32'hc2914159, 32'h42e39634},
  {32'h4520d63d, 32'h440897c6, 32'hc33b1bb5},
  {32'hc311ee53, 32'hc31507f0, 32'h434a7c15},
  {32'h4478771a, 32'hc4e43ede, 32'hc36b5601},
  {32'hc538bfc2, 32'hc23d5108, 32'hc2981c7f},
  {32'hc4d0d270, 32'hc2d330be, 32'hc40a8bec},
  {32'hc370c4a0, 32'h44cbca9a, 32'hc4134676},
  {32'h451ca0da, 32'hc49f04f7, 32'hc2dc330b},
  {32'h43a5a144, 32'hc4aa4680, 32'h439fd8e4},
  {32'hc3963cc0, 32'hc4cd9057, 32'hc4db7666},
  {32'hc2a5b397, 32'hc50eaf85, 32'h44a46f5a},
  {32'hc5425fb7, 32'h421791d4, 32'h4389e7e3},
  {32'h441029dc, 32'h4393d327, 32'hc48d334b},
  {32'h44337529, 32'hc45f07eb, 32'h41c8a483},
  {32'h44832004, 32'h4418a725, 32'hc485a335},
  {32'hc4808a10, 32'h43c8b815, 32'h44e15159},
  {32'h439c94a8, 32'h44572784, 32'hc46a4fce},
  {32'h427af803, 32'hc4bca5c9, 32'hc402ecd9},
  {32'hc4a5906a, 32'h43106c6c, 32'h44b1d4a0},
  {32'h439ccbbf, 32'h44156ea5, 32'hc4fce77f},
  {32'h4447a37d, 32'h443c079e, 32'hc493ee63},
  {32'hc40d6b60, 32'hc412e550, 32'h4516bd9b},
  {32'h43d16189, 32'h44fc71a4, 32'h429fe8a8},
  {32'hc514be9e, 32'hc3c57977, 32'h43b86263},
  {32'h447f80bd, 32'h44dc35e3, 32'h4311494a},
  {32'h43ef2e04, 32'hc415ece4, 32'h43407466},
  {32'h457b1bea, 32'hc3d15cf5, 32'hc380b0c1},
  {32'hc539b738, 32'h42eac81c, 32'hc4071b56},
  {32'h451f1557, 32'h41a90eee, 32'hc1317e2c},
  {32'hc44e007c, 32'hc49052d2, 32'h42390a78},
  {32'h43ad11d4, 32'h4433cc23, 32'h4207a1ba},
  {32'h44c00e86, 32'hc3d257ef, 32'h424d9ca7},
  {32'h449956ae, 32'h44a3ad79, 32'hc4222692},
  {32'h41aa5dd2, 32'hc533ac41, 32'hc3c3a967},
  {32'h42d43102, 32'h4386041e, 32'hc43ef200},
  {32'hc2bbcd55, 32'hc3fa0a84, 32'hc3922310},
  {32'hc42b1c36, 32'hc3cd8371, 32'hc381acb4},
  {32'h44eee249, 32'h446c78ff, 32'h4400b783},
  {32'h440a6fea, 32'hc459cba0, 32'hc151200a},
  {32'h453cb5e4, 32'hc388cecc, 32'h4445c9d0},
  {32'h428569e1, 32'hc5039468, 32'h4351556d},
  {32'h4447a462, 32'h43030a7f, 32'h42922874},
  {32'hc4a18c7e, 32'h438d07b1, 32'hc3f45326},
  {32'h44f2cc82, 32'h43db7eae, 32'h4486cb9d},
  {32'hc4b6da2b, 32'hc2537c70, 32'h43671af6},
  {32'h444b8cb5, 32'hc4d2c004, 32'h44d9782b},
  {32'h4428d00b, 32'h43be3611, 32'hc51c13a2},
  {32'h4254ea14, 32'h44be4f36, 32'hc2933d43},
  {32'hc3509508, 32'hc3b51226, 32'hc507d502},
  {32'hc21c6890, 32'hc3132c1e, 32'h44a7150d},
  {32'h423b58a8, 32'hc4838bc5, 32'hc4a03605},
  {32'h42e25e67, 32'h432dcbf5, 32'h44ea64cc},
  {32'hc455e32c, 32'hc461a37c, 32'hc40b6fdd},
  {32'hc4754f87, 32'h4406918b, 32'h43cd1ae4},
  {32'hc3a88e43, 32'hc56ee082, 32'hc3c454dc},
  {32'h455a35d0, 32'h4354026c, 32'hc4554eab},
  {32'h43d87252, 32'hc4c19b18, 32'h43a22f21},
  {32'h45004b81, 32'h44342003, 32'h43ecdcca},
  {32'hc4bdb998, 32'hc34409f3, 32'h43e2156b},
  {32'h4542bccd, 32'h4417c3fe, 32'h4382520f},
  {32'hc3e7cf6c, 32'h4397db2a, 32'hc29779c3},
  {32'h4482edfc, 32'h43b2d1e9, 32'h439c145a},
  {32'h43780678, 32'hc50cbbd5, 32'hc416ef6b},
  {32'h431fbd86, 32'h4547f8cf, 32'h44242604},
  {32'h43986c3e, 32'hc3f267f0, 32'hc449640e},
  {32'hc3bf4170, 32'hc3376436, 32'h440ab64e},
  {32'hc39addb8, 32'hc44c958a, 32'hc5059f96},
  {32'h43c7e4d2, 32'h42ff8d5f, 32'h44fc351e},
  {32'h451645ee, 32'h4390673d, 32'hc4020af5},
  {32'hc48bc73e, 32'h448d22d0, 32'h448364fb},
  {32'h44a868d9, 32'hc1f51c6c, 32'hc3094be4},
  {32'hc3af759d, 32'hc48a2b72, 32'h44af1a3f},
  {32'hc38e48ea, 32'hc4fa43fe, 32'hc3921d80},
  {32'h3e622000, 32'hc35f8828, 32'h44607967},
  {32'h43b45420, 32'hc3bacb9a, 32'hc4a4dde4},
  {32'hc504aed0, 32'h3f588640, 32'h42987fe2},
  {32'hc4a1d73d, 32'hc3974e2b, 32'hc2880e51},
  {32'hc4207118, 32'h442fe576, 32'h44610e7a},
  {32'h440f188b, 32'hc4ee3bf3, 32'hc4ac0747},
  {32'hc2e9a6d6, 32'h430d59f9, 32'h43a37f00},
  {32'h44097572, 32'hc5578669, 32'hc2471849},
  {32'hc4f415d2, 32'h44fa2718, 32'h43c85a42},
  {32'hc2566755, 32'hc4ae8bc2, 32'h438cf488},
  {32'hc5423631, 32'h43abd2dc, 32'h4304126d},
  {32'h43e6ab59, 32'hc5555b5b, 32'h42e74eaa},
  {32'hc4bb9200, 32'h42c0b5b4, 32'h44651b08},
  {32'h44c8640f, 32'hc3956d96, 32'hc3c7d607},
  {32'hc4dc4ded, 32'hc40254f3, 32'hc2dc676f},
  {32'h445f158b, 32'h427ff04e, 32'hc416dc45},
  {32'h4532064b, 32'h439b1c7a, 32'h41fb4982},
  {32'hc414aca7, 32'h43d1e52f, 32'hc51c4243},
  {32'h45434aa6, 32'h43476f9c, 32'h441764bd},
  {32'hc43e05ec, 32'h435becf6, 32'hc26fb3cc},
  {32'h44bbdb57, 32'hc4b1e437, 32'h42b5d8cb},
  {32'hc4b71329, 32'h44c3610b, 32'h43f34b1c},
  {32'h44eb871e, 32'hc2a8c375, 32'h4358671d},
  {32'hc47666f6, 32'h44cbd0f5, 32'h4386fb7d},
  {32'h446b4246, 32'hc505369f, 32'h428820c5},
  {32'h41839d05, 32'hc3b7c34d, 32'hc49fc5d1},
  {32'h45011a17, 32'h42fb5b26, 32'h43c3120e},
  {32'hc291eb80, 32'h43af991d, 32'hc546fb20},
  {32'hc4a201a5, 32'hc3640b4e, 32'hc3428a40},
  {32'hc475cd5c, 32'h4474d304, 32'h43ce34ec},
  {32'h44e0e435, 32'hc47b6515, 32'hc33de8c1},
  {32'h42e7a054, 32'h43c0a34a, 32'h442067bd},
  {32'h4403db25, 32'hc4d96b15, 32'hc2e7fa01},
  {32'h41543ae8, 32'h4497e701, 32'h445d4ef7},
  {32'hc49f0956, 32'hc31e2688, 32'hc36d8ab9},
  {32'hc4a9bfc8, 32'hc4367691, 32'h440c38c8},
  {32'h4263ba00, 32'hc24fc719, 32'hc4120677},
  {32'h432269bd, 32'h43f4b411, 32'h449c09a1},
  {32'h44bb7000, 32'hc3f0111e, 32'hc3d4d00c},
  {32'h439330e2, 32'h44fd0e2d, 32'h4364cf60},
  {32'hc48f04ba, 32'hc2f6d22e, 32'hc41f5db1},
  {32'hc3853a88, 32'h4503d992, 32'h44162dac},
  {32'h4502e9a5, 32'hc460dbd8, 32'hc4678d6b},
  {32'h4500abb4, 32'h437a0a8f, 32'hc47f7460},
  {32'hc43c36ec, 32'h43a0076f, 32'h440ce31c},
  {32'hc4989681, 32'h43add096, 32'h43b762b9},
  {32'hc34f82cc, 32'hc51bcf74, 32'hc3d8b42e},
  {32'h4524872e, 32'hc02bb888, 32'h418efe40},
  {32'h42dbcfb0, 32'h43211023, 32'hc42fa5e4},
  {32'h44882900, 32'h45198ca3, 32'h4414b499},
  {32'hc4f854f2, 32'hc49a3adf, 32'h43e527bf},
  {32'h452da4b0, 32'h4417e182, 32'h43f7e97d},
  {32'hc4c37735, 32'h40fe5058, 32'h43f9c3c6},
  {32'h4527a4e0, 32'hc3919afc, 32'hc2b0f499},
  {32'h4408c2d0, 32'hc3ce76cd, 32'h4394500a},
  {32'h4385ecdc, 32'h44e0e874, 32'h441ad1bf},
  {32'hc4c1c016, 32'hc49eea37, 32'hc299898c},
  {32'h43a572ab, 32'h43d3ba1d, 32'h43d65da0},
  {32'h4332999f, 32'h435a9099, 32'hc55bfeb2},
  {32'h434c8f1f, 32'h43c362a9, 32'h4546fb73},
  {32'h4209ddf2, 32'hc2bf4001, 32'hc4e388d8},
  {32'h45069293, 32'h44774b65, 32'h43d8096a},
  {32'hc555e791, 32'hc32db4ce, 32'hc25af644},
  {32'h45524c84, 32'h42e54271, 32'hc4145d49},
  {32'hc40f823c, 32'h42753521, 32'hc5120cd3},
  {32'h433e2d60, 32'h43f8f28e, 32'h442fe1cf},
  {32'hc51ea273, 32'h43a0bc86, 32'h4462fa52},
  {32'h448f4f37, 32'h441e54f8, 32'h446aefe5},
  {32'hc4735730, 32'h42b3338e, 32'hc51ce1cb},
  {32'h44f09012, 32'h437b6516, 32'hc3d5a10b},
  {32'h44a04068, 32'h42316346, 32'hc407a70e},
  {32'hc46e7a85, 32'hc4b6a42a, 32'hc3bfed6d},
  {32'h450eb2bd, 32'h4421eaa4, 32'h44705e7d},
  {32'hc413a42b, 32'hc3b71d6f, 32'h4386eb78},
  {32'h43b0528e, 32'h4529526c, 32'hc286a998},
  {32'hc468322f, 32'hc48c5164, 32'hc338a0e1},
  {32'h44309d5d, 32'h44350c58, 32'h438d48e8},
  {32'hc55d9f99, 32'hbfa56328, 32'h43c767b4},
  {32'hc32b7660, 32'h437361d9, 32'h432fe412},
  {32'h4415dc92, 32'hc4bebfdc, 32'h4385b69f},
  {32'h44b54e38, 32'h44500846, 32'hc3e4164b},
  {32'hc31c142e, 32'hc508cfd0, 32'h417dbce3},
  {32'h443e1202, 32'h4445f349, 32'h42f24736},
  {32'hc499bff0, 32'hc39a7913, 32'h433e85eb},
  {32'h44833552, 32'h44c5a9ca, 32'hc34f661f},
  {32'hc518e3c6, 32'hc3410d58, 32'hc3c52bfe},
  {32'h44f4de58, 32'h434686d5, 32'hc44149bd},
  {32'hc4ecc9e2, 32'hc3bd2a1f, 32'h43bad957},
  {32'h44b91e44, 32'h43b5bc70, 32'hc4485e7a},
  {32'hc37310aa, 32'hc53bb496, 32'hc2e46f29},
  {32'h42a85cc0, 32'h452fa256, 32'hc386bc54},
  {32'h44e292f0, 32'h435a54cd, 32'h437f2219},
  {32'h41cf85c0, 32'hc418414c, 32'hc53785be},
  {32'hc38fe205, 32'hc2bd4033, 32'h44cda4da},
  {32'hc4191480, 32'h41e2a46d, 32'hc41ae3e8},
  {32'hc579f40a, 32'hc3820518, 32'h42c44852},
  {32'h43911060, 32'hc38fd185, 32'hc5302c47},
  {32'h4409266a, 32'hc52ecc86, 32'hc3f755e3},
  {32'hc2da76a8, 32'h44f99523, 32'h439df8bb},
  {32'h449dc286, 32'h42d9f20f, 32'h43318852},
  {32'hc4458ce1, 32'h4434fc63, 32'hc3c17ad6},
  {32'h451ffaa0, 32'hc3e2da33, 32'hc37d3bc8},
  {32'hc4ddac1d, 32'h41a32ba5, 32'hc096c05c},
  {32'h44117730, 32'hc463a1ea, 32'hc3e96eec},
  {32'hc432d604, 32'h43d00be7, 32'h443737cf},
  {32'hc309ae8e, 32'h422ce05a, 32'h4416a648},
  {32'h43af059e, 32'h43c36423, 32'h4295571b},
  {32'h4440da26, 32'hc4e42ba9, 32'h4373f127},
  {32'h44717d93, 32'h4444c146, 32'h4330292f},
  {32'h45161d38, 32'hc41d259a, 32'h43e0951e},
  {32'hc42bd1db, 32'hc11ca271, 32'hc5653063},
  {32'hc4bad19e, 32'hc354c5a3, 32'hc31752ea},
  {32'hc4eba202, 32'hc2638d5e, 32'hc455be3a},
  {32'hc191e0c0, 32'hc403d9e7, 32'hc3970b97},
  {32'h439070a6, 32'h43ac0fd7, 32'hc3895284},
  {32'h44bc4ade, 32'hc4a83530, 32'hc2966142},
  {32'hc527506a, 32'h43830040, 32'hc4038cf2},
  {32'h4558d155, 32'h436ce573, 32'hc2021eb4},
  {32'hc4b916c7, 32'h44911b84, 32'h42740535},
  {32'h441854f2, 32'hc521a7b2, 32'hc32ccc00},
  {32'hc398581f, 32'h4430402b, 32'hc41051b4},
  {32'h449b3964, 32'h434d0a79, 32'h4500071a},
  {32'hc54b3f18, 32'hc406700a, 32'hc428a386},
  {32'hc3ca7f10, 32'hc40b12ad, 32'h42f61f4b},
  {32'hc3830d34, 32'hc4265f3f, 32'hc4b8469e},
  {32'h42d27a5a, 32'hc4ca7950, 32'h44be9c24},
  {32'h440af73f, 32'hc40c2bd8, 32'hc4852452},
  {32'hc2ead043, 32'h438a5bdb, 32'hc3ae894e},
  {32'h43aa37f7, 32'hc1df282d, 32'h4405f0fe},
  {32'hc2989120, 32'hc3e5d5ba, 32'hc4c5bec5},
  {32'hc44b40c2, 32'h42dddfdb, 32'h43350243},
  {32'hc4c7a2b9, 32'h43ce450c, 32'hc38bd9fc},
  {32'hc33f53cb, 32'hc55d3a89, 32'h42d452b3},
  {32'h453cee6e, 32'hc26f6a60, 32'h4421a4e3},
  {32'hc38be056, 32'h4509ed8b, 32'hc4ed0f8e},
  {32'hc438d39a, 32'h440fb80c, 32'h4351494a},
  {32'hc4605c26, 32'h43501898, 32'h447033d7},
  {32'hc45c82b8, 32'h427fb5f8, 32'hc47e9fc3},
  {32'hc2c2ea80, 32'hc3da3aa2, 32'h445789fa},
  {32'h42f37c5b, 32'h43fcab79, 32'hc400647a},
  {32'h43fce9ea, 32'h436ea784, 32'h43d6348f},
  {32'hc3f38d60, 32'h41fa2f01, 32'hc3b279ce},
  {32'h450f5cf4, 32'hc4154c9e, 32'h4422bc92},
  {32'hc5556994, 32'hc449ffcb, 32'hc402e2c2},
  {32'h43879d6c, 32'hc3ffbe52, 32'h43e535b8},
  {32'h440a56a7, 32'h443264b5, 32'h441143ef},
  {32'h43d0e464, 32'hc4a4ddd9, 32'hc39e3892},
  {32'hc3c748da, 32'h4575e72f, 32'h43bcab03},
  {32'h44a6120a, 32'hc30d0429, 32'hc270d711},
  {32'hc49b8775, 32'h44b74066, 32'h43847ee2},
  {32'h4507ca51, 32'hc4886663, 32'hc10088dd},
  {32'h44907187, 32'hc46bdd02, 32'h4291ad81},
  {32'hc4011da5, 32'h43add46d, 32'hc4f1f85d},
  {32'h43fdcf64, 32'hc3574487, 32'h4560615b},
  {32'h4475c080, 32'hc5559740, 32'hc3b84a72},
  {32'h432b540c, 32'h44897b30, 32'h42ccb687},
  {32'hc50286d1, 32'hc376b32f, 32'h431c8342},
  {32'h41817e80, 32'h44e878f3, 32'hc3f4a1da},
  {32'hc4dc42d6, 32'hc3594a0d, 32'h4474a759},
  {32'hc38972f5, 32'h44bd0dc0, 32'hc2eed566},
  {32'h420dab55, 32'hc40a5d76, 32'hc40d6553},
  {32'hc227b66c, 32'hc410c75d, 32'h4552a82b},
  {32'hc3f007fa, 32'hc44a6f0d, 32'hc531d398},
  {32'h43d59132, 32'h45217e5c, 32'h42dee70d},
  {32'hc483a830, 32'hc38d5d30, 32'h44545e07},
  {32'h449e345b, 32'h403c8454, 32'hc36fe165},
  {32'hc4bf55f4, 32'hc3c897fa, 32'h446bcf7d},
  {32'h442883fa, 32'h4401e0b2, 32'hc495a564},
  {32'hc29a90d2, 32'hc38ea381, 32'h447a15cc},
  {32'h450779ac, 32'hc3b83c10, 32'hc3a1fc76},
  {32'hc47e9c04, 32'h4409ba09, 32'hc35a745a},
  {32'hc3c8a814, 32'h42c914fe, 32'h42a97388},
  {32'hc38a6433, 32'hc5324c32, 32'h438d677b},
  {32'h43534598, 32'h45654ef1, 32'h4336dcce},
  {32'h43f358ad, 32'hc3593274, 32'h43f91d35},
  {32'hc2b58da4, 32'h450d9925, 32'hc4285f9a},
  {32'hc5159970, 32'hc3e58559, 32'hc33da4ee},
  {32'hc3374739, 32'h44e6ef7c, 32'h429848e5},
  {32'hc2f7ee0a, 32'h43de6dc0, 32'hc2d2f8e9},
  {32'h435c4212, 32'hc47794d2, 32'hc4922eec},
  {32'hc3a4d45f, 32'hc3f0fa2c, 32'h45008067},
  {32'hc30bb0b6, 32'h4324353b, 32'hc442a471},
  {32'h42c59987, 32'h452e6822, 32'h43bdaf2e},
  {32'hc36926b6, 32'hc468c080, 32'hc507357d},
  {32'h43826dbd, 32'h44888164, 32'h442ac937},
  {32'hc3c530a3, 32'hc34cc48e, 32'hc51185e0},
  {32'hc37429ff, 32'h44360432, 32'h4544721e},
  {32'hc11f4708, 32'hc481c04a, 32'hc4000863},
  {32'hc33beaa3, 32'h45330258, 32'h43be9697},
  {32'hc1d73fa8, 32'hc427b505, 32'hc47317c3},
  {32'hc409c138, 32'hc393f27c, 32'h43a68612},
  {32'hc243c160, 32'hc40f5a61, 32'hc5386750},
  {32'hc3cb5988, 32'h451df48d, 32'h425ef17c},
  {32'hc4921890, 32'hc1857b7e, 32'h43ded8f6},
  {32'h4487c438, 32'h442e8599, 32'h443c3cb3},
  {32'hc317aca9, 32'h420c6f69, 32'hc4e2c951},
  {32'h43fec706, 32'h448a7ae3, 32'h429d1c55},
  {32'hc4436a20, 32'hc500ec34, 32'hc38fbea1},
  {32'h4419a3f8, 32'h452c591c, 32'h42cb5691},
  {32'h44365369, 32'hc0ea63f6, 32'hc35f61ce},
  {32'h44137f96, 32'h440eb05f, 32'h43bb8a76},
  {32'hc53f4a95, 32'hc3278730, 32'hc2a0b227},
  {32'h451f1dce, 32'h43897281, 32'h43f522f2},
  {32'hc3933178, 32'h42f72ca7, 32'h438d0f54},
  {32'h443f8d17, 32'h42e7f34c, 32'h431fe083},
  {32'hc46246bd, 32'h4485842a, 32'hc4ccacd0},
  {32'hc433c442, 32'hc2bd9897, 32'h43d7820c},
  {32'h4229ad33, 32'hc3419c62, 32'hc411fcc2},
  {32'hc4dd4d6a, 32'h42efc758, 32'h43e15628},
  {32'hc136a200, 32'hc46e5838, 32'hc4498ce0},
  {32'h43f7c81a, 32'h44ab234a, 32'h41cefdf4},
  {32'hc2fd0408, 32'hc3cadc81, 32'hc5650fda},
  {32'hc31780a2, 32'h43eaa7fe, 32'h455ce85d},
  {32'h44483bb2, 32'hc3c47f79, 32'hc36839de},
  {32'hc468159b, 32'hc45da417, 32'h44982653},
  {32'h44708fb4, 32'h43a2a001, 32'hc33d5f18},
  {32'h44720f1f, 32'h434fc4b3, 32'h43aa27e0},
  {32'h42565910, 32'hc3382d8e, 32'hc43b09d7},
  {32'hc3fc5dd5, 32'h4374f1c6, 32'h4465563c},
  {32'hc4356569, 32'h42590d3c, 32'hc389b0f3},
  {32'hc4519d6d, 32'h42a43f03, 32'h44cd017f},
  {32'hc202ee8a, 32'hc4199948, 32'hc4935b3b},
  {32'h44cd9f62, 32'hc39252f9, 32'h43502df4},
  {32'h441ea619, 32'hc56fd4a4, 32'h41c5abc0},
  {32'hc4e58cdb, 32'h44a9b2d2, 32'h43d5fe76},
  {32'hc468313c, 32'h41392edb, 32'h43066e50},
  {32'hc45ccfaa, 32'h451762b1, 32'h4221a34c},
  {32'h446afabf, 32'hc4d42d1c, 32'hc2b0a2ea},
  {32'hc24cea50, 32'h44b34bf4, 32'h437ea2c7},
  {32'h453b27ab, 32'h440eac8b, 32'hc2e9e287},
  {32'hc52b6b24, 32'h447b04e9, 32'h429e46a1},
  {32'h44b500b7, 32'h41aafd5a, 32'hc1936b5f},
  {32'hc412feba, 32'hc35f50a0, 32'h43b9f505},
  {32'hc305f7dc, 32'hc47ee026, 32'hc52b8678},
  {32'h44bb9c6c, 32'h43b892d8, 32'h44b2b435},
  {32'h44f40dde, 32'h43a1f8c8, 32'hc350585c},
  {32'h4559907d, 32'hc3aaf16f, 32'hc3ff73c3},
  {32'hc453b4a4, 32'h444aa088, 32'h43d29d27},
  {32'h43b88887, 32'hc4732475, 32'h40697745},
  {32'hc4af4fbc, 32'h44a6a08c, 32'h43589b63},
  {32'h451528c4, 32'hc478d948, 32'hc14faf3e},
  {32'hc501a6cc, 32'h4281e4da, 32'hc3240cd5},
  {32'h43d0b480, 32'h42cdf3ee, 32'hc3f20e8d},
  {32'hc43c3490, 32'h40c24384, 32'h43740ed2},
  {32'h449e1668, 32'h4360332c, 32'hc3c0d92d},
  {32'hc41c088d, 32'h4199804e, 32'h4300b1e4},
  {32'h43fab644, 32'hc4489547, 32'hc50ac065},
  {32'h44f99def, 32'hc2eb6148, 32'h43aadb11},
  {32'h43a42482, 32'hc4fd4a41, 32'h42922352},
  {32'hc40a4d74, 32'h4328c1f0, 32'h455bb85b},
  {32'h45204caf, 32'hc30b3694, 32'h43d2a0ba},
  {32'hc53dd394, 32'hc398a78a, 32'h43a399b2},
  {32'h442a441e, 32'hc40f9bc1, 32'hc4b7da3a},
  {32'hc3948038, 32'h42f0fb4b, 32'h4504686c},
  {32'h435eda21, 32'hc3ab2b4b, 32'hc53958c7},
  {32'hc5224a84, 32'h429dd3bf, 32'hc3349c12},
  {32'hc2a9e760, 32'hc38f5fc2, 32'hc4bfa040},
  {32'hc2b5da93, 32'h4538d972, 32'h43bd28e8},
  {32'h44ef5ec0, 32'hc43d970d, 32'hc4b2a582},
  {32'h429c46c0, 32'hc4227ffa, 32'hc4247a7d},
  {32'hc49596d2, 32'h4291710d, 32'h43bc691d},
  {32'h44d76791, 32'h434d8850, 32'hc2caf5e6},
  {32'hc50ca9f5, 32'hc488a503, 32'hc3f8566d},
  {32'h43568e78, 32'h45055e3f, 32'h42570e91},
  {32'hc51161ff, 32'h433957d0, 32'h439718a6},
  {32'h44f581c0, 32'h44335ed8, 32'h42543c43},
  {32'hc3afcccc, 32'hc505c8da, 32'h43cf3672},
  {32'hc4d55ee4, 32'hc36f10bc, 32'h43e740f6},
  {32'hc4567ef8, 32'h43952ea6, 32'h44a63197},
  {32'h440cd8e4, 32'h43f3d8c7, 32'hc30bd95c},
  {32'h44ae11d1, 32'h43e05c68, 32'hc2dcbbbc},
  {32'h451df79f, 32'hc2741b34, 32'h43d22904},
  {32'hc3dc66bd, 32'hc45c5995, 32'hc4b8b569},
  {32'hc42cacab, 32'h44650ffb, 32'h43b0ddac},
  {32'hc3cd2d00, 32'hc51b837f, 32'hc356d1dc},
  {32'h451f288b, 32'h4344bf9c, 32'h423c8f7a},
  {32'hc3a52804, 32'hc3427b5e, 32'hc41d8f4d},
  {32'hc368bb80, 32'hc43e8884, 32'h4409be4d},
  {32'hc5328f1e, 32'hc3ddc5c7, 32'hc402a39f},
  {32'hc4133956, 32'hc4677b48, 32'h4404f5a4},
  {32'hc3dbf230, 32'hc4871bc9, 32'hc49555ad},
  {32'h44964860, 32'h44ac030b, 32'h4386e3ce},
  {32'hc3d7b654, 32'h43b41bcb, 32'hc4468d59},
  {32'h43f2317c, 32'h449eb470, 32'h43c0ebcd},
  {32'hc4f31077, 32'hc465f83a, 32'hc473dd2c},
  {32'h4390a855, 32'h44ee5e7d, 32'hc36a7ac8},
  {32'h44ab2cf1, 32'hc3efba77, 32'hc2c68beb},
  {32'hc580f0fd, 32'hc311c035, 32'h423401ed},
  {32'h443cab46, 32'h449e30bc, 32'h4415426f},
  {32'hc4bea50e, 32'h4381ef64, 32'h42d9a220},
  {32'h4481a1f0, 32'h4488508b, 32'h42bb47c2},
  {32'hc4739524, 32'hc4a43928, 32'h42d9cdea},
  {32'hc3eeb781, 32'h43d60f1d, 32'h428d1962},
  {32'hc399d1a0, 32'hc4cefe93, 32'hc48143da},
  {32'h4433f888, 32'h44342c54, 32'h441a6338},
  {32'h44ef1e17, 32'h4400b543, 32'hc3785773},
  {32'h43276f3a, 32'h4498e897, 32'h41beaa2d},
  {32'hc4f41e27, 32'hc33ea99d, 32'h43f44d94},
  {32'hc3bfd7e8, 32'h440fc112, 32'hc38b4eee},
  {32'hc3dbb4dc, 32'hc437e4a2, 32'h44af3340},
  {32'h444665ca, 32'hc3b2483c, 32'hc3be0262},
  {32'h447a9fe2, 32'hc3792d0b, 32'h439161e6},
  {32'h455f26a9, 32'h43f148bb, 32'hc3f664df},
  {32'hc4934c21, 32'hc46062b3, 32'hc33d997c},
  {32'hc3e1e75c, 32'h444f6819, 32'hc23b0062},
  {32'hc50ed59a, 32'hc446d38c, 32'h44193a39},
  {32'h437e06d0, 32'h447c7d36, 32'hc3bca4ca},
  {32'h441f8d4f, 32'hc468ab63, 32'h433490d8},
  {32'hc2db72c4, 32'hc3b6772d, 32'hc5315a30},
  {32'hc45c06de, 32'hc41dd427, 32'h43864e7e},
  {32'hc3442107, 32'hc1aafaac, 32'hc499a205},
  {32'hc4c66ac2, 32'h4318632c, 32'h440ab014},
  {32'h4579856c, 32'h4409cdd0, 32'hc325c7f1},
  {32'h448f0193, 32'hc4a41cb3, 32'h413a65f3},
  {32'hc4499d38, 32'h4495df31, 32'h44509d86},
  {32'h4319c920, 32'hc5186e86, 32'h428b18c8},
  {32'hc332b4e0, 32'h44652a23, 32'hc3b6e0d6},
  {32'h44c5f21c, 32'hc35b2931, 32'hc3b8f2e6},
  {32'hc5046460, 32'hc31bf6d7, 32'hc290fc1a},
  {32'hc3ba6e4a, 32'h438d43f5, 32'hc2ab2b2d},
  {32'hc554d310, 32'h4367f2bb, 32'h4390b437},
  {32'h45590f5d, 32'hc27b37a4, 32'h4423d8bc},
  {32'h43afb002, 32'h44a79511, 32'hc3d8ef53},
  {32'h440854bb, 32'hc3f784c1, 32'h442cb218},
  {32'hc4ea38b2, 32'h43ebeef6, 32'hc1b958f0},
  {32'h45275ad5, 32'h443fa348, 32'h444aaf9c},
  {32'hc53834c4, 32'h433bf651, 32'hc1bad499},
  {32'hc40fc66e, 32'hc3686735, 32'h42b61d1d},
  {32'hc4c392f2, 32'h43a2d0dc, 32'h43fb8d15},
  {32'h44cae21a, 32'h43abaff4, 32'h449afe6d},
  {32'hc4b33f48, 32'h437a2ee2, 32'hc4378270},
  {32'h44895396, 32'hc43dd296, 32'h43331a4d},
  {32'hc489e4dc, 32'h44b5dea2, 32'hc4e73d97},
  {32'h44da1e42, 32'hc397f0a2, 32'h439963da},
  {32'hc48bf734, 32'h42897aec, 32'hc4321afd},
  {32'hc3c0f1f2, 32'hc4ac60cc, 32'h446708f5},
  {32'hc40656cd, 32'h4333b847, 32'hc300488b},
  {32'h44a1032e, 32'h4382c118, 32'h44d03ff3},
  {32'hc43c7fb4, 32'hc3bd9ea6, 32'hc5342483},
  {32'hc4bfc06a, 32'h4379a597, 32'h436ce084},
  {32'hc393df44, 32'h442b2bd3, 32'hc4b6a190},
  {32'h4375a5fe, 32'h44a6cace, 32'h449c4f61},
  {32'h4300e107, 32'hc45dac0a, 32'hc40887e0},
  {32'hc3b2fe87, 32'h44f15e3e, 32'h433a3d3b},
  {32'h4432fe83, 32'hc5238912, 32'h43a02f8c},
  {32'hc501887b, 32'h43492240, 32'hc3555494},
  {32'hc41e0fd2, 32'hc38abc2c, 32'h448d0d66},
  {32'hc3e6d94e, 32'h441ddbe5, 32'hc4e7f46f},
  {32'h44966ff0, 32'hc4ad0560, 32'hc32c25e7},
  {32'hc3169997, 32'hc3a25dac, 32'h453bef24},
  {32'h44237dfe, 32'hc43b4559, 32'hc5174148},
  {32'hc46b5a00, 32'hc3c444cf, 32'h4440731a},
  {32'h443947c0, 32'hc443a83c, 32'hc3bcfad0},
  {32'hc558ced0, 32'hc353e76c, 32'hc201bc2e},
  {32'h45135ece, 32'hc407fa82, 32'hc2ac176b},
  {32'hc4405a46, 32'h43b6ba18, 32'hc3d453f2},
  {32'h4361b82a, 32'hc515c58f, 32'h4230a79d},
  {32'h4388edba, 32'h43dc9be2, 32'hc4414928},
  {32'h441f6ac4, 32'hc411612a, 32'h41d9f84a},
  {32'hc3c6f6f4, 32'hc382ca55, 32'h43c110ce},
  {32'hc39cc4c5, 32'h42c8183e, 32'h42fdda39},
  {32'h440025e4, 32'hc3a21cb0, 32'hc2bcc4c8},
  {32'h457c97d5, 32'hc3c9ea9a, 32'h438792cf},
  {32'h42ddca80, 32'h4543394a, 32'hc23dc3be},
  {32'h43c04c9a, 32'hc4c36777, 32'hc36da599},
  {32'hc527f7bd, 32'h4423c2b4, 32'h432b63e3},
  {32'h43bc26ae, 32'hc4ed6c64, 32'hc43e5cdf},
  {32'hc502eb30, 32'hc2d1e15a, 32'hc344d72f},
  {32'h445611d6, 32'h44a433c5, 32'hc421cfe9},
  {32'hc493616c, 32'h42afeb65, 32'h44970269},
  {32'h43861275, 32'hc36cb619, 32'h44aeb6cb},
  {32'h43f6f033, 32'h453871db, 32'h4373713c},
  {32'hc43f9b29, 32'h43596d8f, 32'h43a6aac2},
  {32'h43f71991, 32'hc360f9df, 32'hc53f7b40},
  {32'hc3be7179, 32'h43632d80, 32'h4539259f},
  {32'h411b5100, 32'h43a4c0a5, 32'hc48e4d9e},
  {32'h43a667ee, 32'hc2adf782, 32'hc4cb64e6},
  {32'hc3e25778, 32'hc50c219a, 32'h44e57218},
  {32'h44522d16, 32'hc4fdbbd5, 32'hc4989a89},
  {32'h44a2b316, 32'h43a290b7, 32'hc44164d7},
  {32'hc3b7d2f8, 32'hc2a84993, 32'h455bb7ef},
  {32'h43815c25, 32'h4361b9c2, 32'h431a2b4f},
  {32'hc4809249, 32'hc45f9f57, 32'h433909eb},
  {32'hc34e7902, 32'h43d10428, 32'hc520ac15},
  {32'hc2ea8598, 32'hc4b2e55d, 32'h44234302},
  {32'h44527670, 32'hc2f42a65, 32'h432a9faf},
  {32'hc56621ca, 32'hc2a594c7, 32'hc40a9b1a},
  {32'hc4c21348, 32'h42357d2a, 32'hc2c84161},
  {32'hc50a1bc1, 32'h432586ee, 32'hc219d9f6},
  {32'h4515d74e, 32'h43cc1506, 32'hc354d8e6},
  {32'h4499bbbf, 32'hc3ac5e9c, 32'hc2ca4d6b},
  {32'h41483580, 32'h4521bdb2, 32'h43acc16a},
  {32'hc49bc31e, 32'hc4a2e511, 32'hc3cd2d32},
  {32'h439415b4, 32'h4439b98f, 32'h4317620b},
  {32'hc33483b2, 32'h442348e1, 32'h44538a09},
  {32'hc48cae2b, 32'hc258ebfb, 32'hc362f659},
  {32'h448e9c4e, 32'h4490c198, 32'h44044d4f},
  {32'h440e1860, 32'hc47c206e, 32'hc3804633},
  {32'h445002c4, 32'h44482049, 32'h44afa48d},
  {32'h43204e4f, 32'hc470fd3e, 32'hc482e19a},
  {32'h433a26f1, 32'h442e5c62, 32'h44cb3884},
  {32'hc4aa4dce, 32'hc356a94f, 32'hc490bbf9},
  {32'h44e22492, 32'h439329cd, 32'h44453739},
  {32'h423a2090, 32'hc4e8ff15, 32'hc2af3e11},
  {32'h438b0cc5, 32'h446a13f2, 32'h4476e639},
  {32'hc4717a4c, 32'hc43d03b7, 32'hc410ac1d},
  {32'hc3e86d5c, 32'h438aa2bc, 32'h449439db},
  {32'hc29470e8, 32'hc4f29059, 32'hc3d77327},
  {32'h43ae50cb, 32'h43493340, 32'h4507c036},
  {32'hc2f011e0, 32'hc28948d9, 32'h430e19dd},
  {32'h4519016b, 32'h42a0c588, 32'hc3a2a856},
  {32'hc31a84a0, 32'hc48733f6, 32'hc5735460},
  {32'h450cf6ab, 32'h4398a826, 32'h43841160},
  {32'hc52634c8, 32'hc4716eb7, 32'hc3f4ea15},
  {32'h45783cad, 32'h43baa1b4, 32'h437ca0fe},
  {32'hc3b7f7d7, 32'hc37fdc69, 32'hc2f75692},
  {32'h43b8fbd8, 32'h450f0839, 32'hc3e62d62},
  {32'hc4c4fcbd, 32'hc46677f2, 32'hc29189bd},
  {32'h4495612d, 32'h43071316, 32'h441ba0a7},
  {32'hc4c8fba7, 32'hc3ef8b8a, 32'hc41c85fe},
  {32'h45292706, 32'h4366930a, 32'h44486981},
  {32'hc1a39150, 32'h44af43bb, 32'hc4d87393},
  {32'hc467daa4, 32'h444ebfed, 32'h438c3a69},
  {32'hc2d2c86c, 32'h41bae989, 32'hc4b2a0fd},
  {32'hc43d41c4, 32'h44cf9f59, 32'h439d5de2},
  {32'h44ef16bc, 32'hc40b2f23, 32'hc326d38a},
  {32'hc5380c49, 32'hc3071b12, 32'h42e22093},
  {32'h44dba5cb, 32'h41b74ca3, 32'hc430e5bb},
  {32'hc547f521, 32'hc3c7c982, 32'h42b20c75},
  {32'h428ecb32, 32'h43525a3b, 32'hc46c54a1},
  {32'hc2feda2c, 32'hc4be13ed, 32'h452c6eed},
  {32'hc41d7c6c, 32'h43fb3ddd, 32'hc4c27470},
  {32'h43a947d8, 32'h447b1c63, 32'h43bdcd08},
  {32'h40ddf270, 32'hc4264a4a, 32'hc4271f1f},
  {32'hc4076f62, 32'h43af5dbc, 32'h44d5addb},
  {32'h443870c2, 32'hc4321965, 32'h40979bf1},
  {32'hc4765bc3, 32'h43f125ff, 32'h44601ac6},
  {32'hc309a9a8, 32'hc45e9bff, 32'hc49f9942},
  {32'hc522698d, 32'hc29e45a6, 32'hc2406720},
  {32'h45092aee, 32'hc40c697d, 32'hc33242bb},
  {32'hc3af8d82, 32'h4459fe9c, 32'h4425f7da},
  {32'hc3aa546e, 32'hc4227472, 32'hc236abf2},
  {32'hc4a5d1c0, 32'h44be4f21, 32'hc2a9ed7d},
  {32'h45366f70, 32'hc1c33db6, 32'hc1f7e077},
  {32'hc41122b7, 32'h439e0f07, 32'hc26417ce},
  {32'h450962a8, 32'h431285c5, 32'h43accc23},
  {32'hc5462186, 32'hc3b26a29, 32'h4399bbc1},
  {32'h456de039, 32'hc344a192, 32'hc36bd1ee},
  {32'hc41ef595, 32'hc201f9f7, 32'hc3dd6def},
  {32'hc4b77795, 32'hc2f2d9db, 32'hc4f38e80},
  {32'h44fb6cca, 32'hc2c2d66e, 32'h438bf018},
  {32'hc3065a53, 32'h44c2c784, 32'h43af6ec6},
  {32'h44c008e0, 32'hc4ad76cd, 32'hc4012f6e},
  {32'hc47d9af8, 32'h4486f35a, 32'h43b7a632},
  {32'h450988db, 32'h43e50fa0, 32'hc30f2421},
  {32'hc44dff5a, 32'h4393fba7, 32'hc3f80b7a},
  {32'h44162a56, 32'hc5131998, 32'hc18732ae},
  {32'hc4a0a0b8, 32'h4251fdd2, 32'hc323275d},
  {32'h43074b04, 32'hc1c1df71, 32'h45533025},
  {32'hc2907da0, 32'hc4247436, 32'h4414e313},
  {32'hc39e7348, 32'hc1bbb5e6, 32'h42e6db7e},
  {32'h41d762a0, 32'hc38ccdf8, 32'h452f0af4},
  {32'hc39a8216, 32'hc48f5d80, 32'hc5105f42},
  {32'h4333157a, 32'h441446b0, 32'hc387088b},
  {32'h44ba7697, 32'hc477d4e8, 32'hc411b161},
  {32'h43354999, 32'h4405b69a, 32'h44a2bbc1},
  {32'hc406496e, 32'hc2c0d53e, 32'h437bdf6f},
  {32'hc3f2daf8, 32'h435773b0, 32'h448414b4},
  {32'h45024291, 32'hc397559f, 32'hc46918c3},
  {32'h43ade038, 32'h444c2423, 32'h4466eda9},
  {32'hc34facee, 32'hc57a55a9, 32'h434278d6},
  {32'hc44ba2e8, 32'h449d42c6, 32'h4422ec97},
  {32'h453c930a, 32'hc268e887, 32'h42ee4a3a},
  {32'hc3377c76, 32'h439053ef, 32'h45251d9f},
  {32'h44b35a14, 32'hc46ac757, 32'hc4c11958},
  {32'h44a197be, 32'h433dba71, 32'hc50012da},
  {32'hc52c245c, 32'hc23f273c, 32'h44a22b6d},
  {32'hc4455d94, 32'hc2bb5eef, 32'hc4347885},
  {32'hc32e9ced, 32'hc5260dc9, 32'h42a3f8d8},
  {32'hc24120c0, 32'h45117900, 32'h43e8d50f},
  {32'hc3852962, 32'hc479d919, 32'hc24098a3},
  {32'hc2d406e0, 32'h452f41f6, 32'hc37560f7},
  {32'hc57545fa, 32'hc30f3aa0, 32'h434cea0c},
  {32'h43ff47f6, 32'h43cda2b4, 32'h4402265b},
  {32'hc40cf188, 32'hc40bbab8, 32'hc3d393e9},
  {32'h43ff40b3, 32'hc2111603, 32'hc3dd0999},
  {32'h448e1e87, 32'h43b62e9d, 32'h438d0d61},
  {32'h447da24c, 32'hc2c2230b, 32'h445ec377},
  {32'hc47584dc, 32'hc43e99c6, 32'hc4e046e8},
  {32'h43292f08, 32'h43a3cc2e, 32'h43f899f2},
  {32'hc39ead38, 32'hc43e16c7, 32'hc4eb3b0b},
  {32'h43cb4024, 32'h4493b423, 32'hc30b34bb},
  {32'h440666d4, 32'h42d29a0a, 32'hc4820239},
  {32'h4561fc1d, 32'h4360edbe, 32'h443dff11},
  {32'hc517ff90, 32'h43f3478a, 32'hc42b1ccd},
  {32'h44e0bdf6, 32'h4448ae2e, 32'hc229f30c},
  {32'hc1a67e00, 32'hc4993943, 32'hc47249a8},
  {32'h43af3560, 32'h44823bdc, 32'h44569d9b},
  {32'hc39b05e7, 32'hc4034988, 32'hc38d8c43},
  {32'h42bbf2dc, 32'h44d1a49e, 32'h434ca64d},
  {32'hc427c3e1, 32'h42e29124, 32'hc5585338},
  {32'h44af5068, 32'h43cc18b0, 32'h436814f0},
  {32'hc42e03e6, 32'h44615a40, 32'h43a85c47},
  {32'hc4922ffe, 32'hc4a417b8, 32'h437dd56e},
  {32'h4359cd16, 32'h452db929, 32'h442277dc},
  {32'h44bbc0e1, 32'hc3c963d3, 32'h428ba046},
  {32'h448e293a, 32'h44612880, 32'hc22ef30e},
  {32'hc3a6a84c, 32'hc4e435c5, 32'hc23f1002},
  {32'h44e99be6, 32'hc32523e1, 32'hc3bab452},
  {32'hc49eeed0, 32'hc3d846dd, 32'hc332fc88},
  {32'hbfac37c0, 32'h443028ed, 32'h44150d04},
  {32'h44a65e19, 32'hc42093a4, 32'h43788ea3},
  {32'h440351e1, 32'hc1e27229, 32'h43cc6f0d},
  {32'hc50611b8, 32'hc36aa211, 32'hc3293409},
  {32'h4443636f, 32'h405ff614, 32'hc3f698b9},
  {32'hc3ede95c, 32'hc3d1d5b2, 32'h44feaaed},
  {32'h44d4a1e8, 32'h43908cb6, 32'h4219ff86},
  {32'hc5351e73, 32'hc1d4c502, 32'hc3e7a9df},
  {32'h439aaf4e, 32'hc3bd9677, 32'hc4a836f2},
  {32'hc42287fb, 32'hc2471489, 32'h44f9a994},
  {32'hc34ba953, 32'hc25d2b4a, 32'hc4870be4},
  {32'hc49fe346, 32'hc497a6e3, 32'h450f56d7},
  {32'h442b2754, 32'h44e20dbf, 32'hc399c6c7},
  {32'h43bca4e1, 32'hc50240e4, 32'hc436939d},
  {32'hc39542fd, 32'hc38bd7b3, 32'hc54c41c4},
  {32'hc51a0e94, 32'hc3d5671f, 32'h4391f996},
  {32'h452d2a86, 32'h42233f20, 32'hc2e2c2cc},
  {32'hc4914340, 32'h43b56721, 32'h446a67b1},
  {32'h4423ec30, 32'hc3ccbf6e, 32'hc4dd20fa},
  {32'h4501e097, 32'hc48a34a2, 32'h43e7cd35},
  {32'hc580e3bf, 32'h43305d05, 32'h441cf51f},
  {32'hc3181356, 32'hc4f51dad, 32'h42ec14e6},
  {32'hc5082c73, 32'h444b039e, 32'h441b14a8},
  {32'h43a7f7e6, 32'hc51d668c, 32'h43cc412d},
  {32'hc5307dc4, 32'hc3074cc0, 32'h429395e5},
  {32'h44e8698f, 32'h433813f0, 32'hc3b12153},
  {32'hc4283439, 32'h4436ddc1, 32'h4459bd2c},
  {32'h443e18e3, 32'h4241c1a0, 32'h44100a5d},
  {32'h43ca3f58, 32'h44841e05, 32'hc4931c55},
  {32'h439579e0, 32'h42029992, 32'hc37f015e},
  {32'hc34e8830, 32'h447379ff, 32'h430e1134},
  {32'hc305bf24, 32'hc551fcd5, 32'h4210ac67},
  {32'hc4507f60, 32'h44237c78, 32'hc4004d62},
  {32'hc48c66c9, 32'hc37f8d81, 32'hc339911d},
  {32'hc4cc6977, 32'hc3818b9e, 32'hc47fcd0b},
  {32'h42e89da8, 32'h43295de6, 32'h4514e508},
  {32'h44e6769c, 32'h43e8ee00, 32'h43a899f1},
  {32'h4413bd5f, 32'hc4b6a8e7, 32'h449251c4},
  {32'hc5825051, 32'hc3281f92, 32'hc2f56e88},
  {32'hc3ff44dc, 32'hc2d02ede, 32'h41eccd5c},
  {32'hc3d7f588, 32'h4503cea1, 32'hc3ad2c00},
  {32'hc3924f67, 32'hc4061df9, 32'h44977bb2},
  {32'hc481b9f4, 32'hbfe9780c, 32'hc0ae1ec0},
  {32'h44d1884d, 32'h44312be7, 32'h4465acc1},
  {32'hc5863610, 32'hc37f2594, 32'h4338059d},
  {32'hc4d789f4, 32'h4290f0fa, 32'h439d2b71},
  {32'hc30e561a, 32'hc358e8e0, 32'hc3e15fe5},
  {32'h4307693b, 32'h4498b43c, 32'h44fdb1b8},
  {32'h4300ba41, 32'h4497223e, 32'hc4c22fe2},
  {32'hc4621169, 32'h43fa145c, 32'hc41311a7},
  {32'h43d19bc9, 32'hc42280b2, 32'h451f7c83},
  {32'hc4a10d1d, 32'h44520242, 32'h4374703d},
  {32'h43ae99d2, 32'hc3a046bf, 32'h4473dcb2},
  {32'hc47ab738, 32'h42c15554, 32'hc51c996c},
  {32'h453b47ef, 32'hc2ffe668, 32'h435ded69},
  {32'h431fd0cc, 32'hc50c49a1, 32'h44e4fb85},
  {32'hc510a2ac, 32'h412ae9c4, 32'h444062ec},
  {32'hc4311595, 32'h4436a34f, 32'h4455da69},
  {32'hc3e3fc28, 32'hc474d9e8, 32'h440d27c8},
  {32'hc3a2af04, 32'h4459aa43, 32'hc44368a5},
  {32'h44a294c3, 32'hc2af7910, 32'h43a1af25},
  {32'hc3c3ae5a, 32'h4296bc0f, 32'hc3ef0156},
  {32'hc3a85818, 32'hc4c43c5c, 32'hc4223efb},
  {32'h435bb612, 32'hc33af982, 32'hc4f83f58},
  {32'h449b115a, 32'h43ad9d14, 32'h43a3311a},
  {32'hc3826b20, 32'hc453a144, 32'hc430cad5},
  {32'h44a3aa7d, 32'h447ba57a, 32'hc381d9bd},
  {32'hc497bb83, 32'hc1ff4233, 32'h41816d44},
  {32'hc30869f6, 32'hc55ee5ec, 32'hc3cbc817},
  {32'hc552ae8c, 32'h42e5a2c8, 32'h42884b55},
  {32'h449419c6, 32'hc1a6a864, 32'h43f17419},
  {32'hc457fa20, 32'h45131d22, 32'h43302472},
  {32'h44665255, 32'hc4ccdd4b, 32'h43beef7f},
  {32'hc4605b18, 32'hc33a8bf5, 32'h43890b02},
  {32'hc3fc07db, 32'h44f5151a, 32'hc4cb52d0},
  {32'hc4afc2b6, 32'h4251e291, 32'h43497fcc},
  {32'hc46bd216, 32'h43f064e0, 32'h44ac6c11},
  {32'h44e420b4, 32'h43ed7e53, 32'hc308dc66},
  {32'hc307a32a, 32'hc43dff82, 32'h43e3d57d},
  {32'h4379013c, 32'h45461055, 32'hc41ea634},
  {32'hc4547004, 32'h43ba3427, 32'h450750f3},
  {32'h44b75924, 32'hc3a68304, 32'hc44bdbfa},
  {32'h443c9606, 32'hc464e5d2, 32'hc389a88d},
  {32'hc38a8ff7, 32'hc3201a72, 32'h4400b17a},
  {32'h443fa976, 32'hc4b83640, 32'hc4b2437b},
  {32'h44d70569, 32'h440fc66c, 32'hc413bfc6},
  {32'hc38a85fc, 32'hc4063276, 32'h44bd483f},
  {32'h41e570b0, 32'h4396544c, 32'h42a6e94d},
  {32'hc459a5a0, 32'hc3d6c075, 32'h44a5d22f},
  {32'hc28a47f7, 32'h4448a37f, 32'hc440acda},
  {32'h4409b295, 32'hc33d5aa3, 32'h448e44b3},
  {32'h41a28300, 32'hc305fc22, 32'h43e20ea4},
  {32'hc5599741, 32'h420fa408, 32'hc3b7ecce},
  {32'h452e9b04, 32'hc205c541, 32'h435b494a},
  {32'hc43caf16, 32'hc4f3c175, 32'h43ee7e0d},
  {32'h4557ff2f, 32'h439acdfc, 32'h4390e06d},
  {32'h446e6e06, 32'hc420bdff, 32'h437da174},
  {32'h43d7ef53, 32'h44c7f57e, 32'h43a07e95},
  {32'h428b1c30, 32'hc57db83d, 32'hc33c63d6},
  {32'h440d2118, 32'hc1b4a7d3, 32'hc3bad2df},
  {32'h44c9f719, 32'hc39a63d5, 32'h43d9ed5c},
  {32'hc39c1605, 32'hc5637f16, 32'hc3752789},
  {32'hc1c9eb20, 32'hc390404d, 32'h44b5c7fa},
  {32'h443c86bf, 32'hc360dbb4, 32'hc3457654},
  {32'h452b5ece, 32'hc274ed9b, 32'h440ef562},
  {32'hc52ec6ce, 32'hc4126b77, 32'h44243242},
  {32'h4518c9ec, 32'hc39bd345, 32'hc319255c},
  {32'hc3797c93, 32'hc415763b, 32'hc50dde98},
  {32'h44d1ed33, 32'h439e4802, 32'h44298e9f},
  {32'hc354ccd9, 32'hc4651fd7, 32'hc24d22ff},
  {32'hc4365294, 32'hc3c6ad29, 32'h44cc0e1f},
  {32'hc4dcb66a, 32'h4259ba56, 32'hc4016c3c},
  {32'h43148e52, 32'h44ad7ea7, 32'h433a5f3d},
  {32'hc2d020d8, 32'hc53e2bf8, 32'hc2926083},
  {32'hc389c8d0, 32'h443e16f8, 32'h45256c24},
  {32'hc4d7d237, 32'hc0208ac0, 32'h42042166},
  {32'h44f2ef05, 32'h43720afd, 32'h4488cd36},
  {32'hc3c5725c, 32'hc2932874, 32'hc4ffe5f2},
  {32'h446c6136, 32'hc2ae809e, 32'h43ee3852},
  {32'hc29f3804, 32'hc569d73e, 32'hc2dc5b69},
  {32'h436cc898, 32'h45796967, 32'hc21c40b2},
  {32'hc4f5ddaf, 32'h4356032a, 32'hc2e0a7b5},
  {32'h44e7aa21, 32'h442ec1b0, 32'hc36891fe},
  {32'hc502f236, 32'hc3f06b6f, 32'h438a857e},
  {32'h451ec808, 32'h43cb42eb, 32'h43828a93},
  {32'hc51bb60c, 32'hc3ccb4ee, 32'h42f37eac},
  {32'hc1d47f00, 32'hc2966ff6, 32'h44353d7e},
  {32'h43a9e8d2, 32'hc3950d0e, 32'hc4d53232},
  {32'hc4a98c32, 32'hc30ff1f1, 32'h449f11da},
  {32'hc4805538, 32'hc389b7ec, 32'hc1997b6d},
  {32'hc544563f, 32'h4385d734, 32'h426b6a8e},
  {32'h421bfd00, 32'hc4bcf871, 32'hc48f72c3},
  {32'h42480300, 32'h43a3ae9e, 32'h42ca691e},
  {32'h4535494e, 32'h4360e0e2, 32'hc3e86088},
  {32'hc265ad30, 32'h4500d647, 32'h44b1f047},
  {32'h446a6f3d, 32'hc40c80fd, 32'h41d2e9b6},
  {32'h435fcc72, 32'h440ac815, 32'h4461a95c},
  {32'h44c3dc53, 32'h43ba6023, 32'hc40834e8},
  {32'hc436ab16, 32'h44025945, 32'hc3a2c7c4},
  {32'h44adf5ce, 32'hc2e7f643, 32'hc405ced4},
  {32'hc19d0de0, 32'h44f1f9bf, 32'h43454f72},
  {32'hc2e37208, 32'h4377892f, 32'hc47c6255},
  {32'hc43fb13e, 32'h43e97149, 32'h449caad3},
  {32'hc2a104fc, 32'hc4df1260, 32'hc503c3b0},
  {32'h44f9da58, 32'h437a4eb4, 32'h43d3f262},
  {32'h44dde26c, 32'hc448e56c, 32'hc3d82371},
  {32'hc3bd564c, 32'h4449b4f2, 32'h4422e765},
  {32'h44888a0a, 32'h41e4649f, 32'h43851d92},
  {32'hc44a7ce8, 32'h451e62be, 32'hc29dbe13},
  {32'h44de23f2, 32'hc4964c38, 32'h43988d98},
  {32'hc37ba99a, 32'h444f78bc, 32'h429ada0d},
  {32'h45630e6e, 32'h43312165, 32'hc38c7b8a},
  {32'hc37882d0, 32'h43d5a400, 32'hc3a6b957},
  {32'h4502476b, 32'h4202c516, 32'hc3c9b553},
  {32'hc446bcbb, 32'hc26aec74, 32'h4430106c},
  {32'hc545fabc, 32'hc347b411, 32'hc373b950},
  {32'h4411d83c, 32'hc36216f6, 32'h454ff059},
  {32'hc43b8ac8, 32'h42692171, 32'hc3d7b2bd},
  {32'h4516e474, 32'h44042c18, 32'hc3e0a575},
  {32'hc3d67414, 32'h45086f8f, 32'h43c819bc},
  {32'h441ae102, 32'hc4164fad, 32'hc3f3c612},
  {32'h438b9c60, 32'h458634b7, 32'h42829f5d},
  {32'hc35c7562, 32'hc5725eb8, 32'h40b2c652},
  {32'hc4913ccb, 32'h41ab07c8, 32'h415ebfc2},
  {32'h444a11e8, 32'h430957e6, 32'h4363546f},
  {32'hc3833ae0, 32'h4380af18, 32'hc48339b3},
  {32'h44c75eee, 32'hc38d4166, 32'hc39c4054},
  {32'hc483c965, 32'h42b76bbc, 32'h43b4edca},
  {32'h44acac7b, 32'hc336fe47, 32'hc439541a},
  {32'hc46dfb9f, 32'h438be3c6, 32'h43c3bc76},
  {32'h44d92bac, 32'h443d1a2a, 32'hc42333e3},
  {32'hc34aadfa, 32'h4481f4d7, 32'h44a9327d},
  {32'h457dc010, 32'hc2db9676, 32'h422cd94d},
  {32'hc421a918, 32'hc238ca5d, 32'hc1a1ec54},
  {32'h44a8fcbb, 32'h444d5c5b, 32'hc497d9fc},
  {32'hc107e1ad, 32'h4402bbc8, 32'h44b3d1aa},
  {32'h43fade68, 32'hc4824df3, 32'hc42a5744},
  {32'hc2f274e0, 32'h43ce7641, 32'h4505f5d1},
  {32'hc3df532b, 32'hc3cc3572, 32'hc44e7e45},
  {32'hc55026f2, 32'h439cff60, 32'hc244ecde},
  {32'h43721518, 32'hc4222f72, 32'hc554139c},
  {32'h446576d4, 32'h43741c9e, 32'hc41fdd17},
  {32'hc4072eec, 32'h43211f29, 32'h44ae8bfb},
  {32'h42f28db0, 32'h43d58da7, 32'hc189591d},
  {32'h418ff480, 32'hc5001168, 32'h421da724},
  {32'h448af24c, 32'h433193ee, 32'h435c89fc},
  {32'h4513d67a, 32'hc2c778c4, 32'hc2e9ccb8},
  {32'h410f5800, 32'h44925e2a, 32'h43d831da},
  {32'hc3a86efe, 32'hc5666254, 32'hc39d4b68},
  {32'h4546848f, 32'hc3215ce6, 32'h43de9b96},
  {32'hc2c87120, 32'hc455e325, 32'h451dc38f},
  {32'h43fca034, 32'h42102b5e, 32'hc479f1d4},
  {32'hc415f3dc, 32'h41360224, 32'hbff04c20},
  {32'h448eb4c3, 32'h437c3df6, 32'h44123145},
  {32'hc38441c8, 32'hc4bf4f5f, 32'h432505b8},
  {32'hc41a1846, 32'h440e40d9, 32'h43a23c7f},
  {32'hc3f8151e, 32'hc3e931fe, 32'hc34f5c46},
  {32'h439287ac, 32'h4503606a, 32'h41489564},
  {32'h44a09952, 32'hc4275e8b, 32'hc399b5f3},
  {32'h44d06082, 32'h445abb7b, 32'h443430f2},
  {32'hc54aa209, 32'hc0f4cd91, 32'hc35e8148},
  {32'h456065e5, 32'hc393ca03, 32'hc363d9c4},
  {32'hc38875b4, 32'hc36ab7f5, 32'hc53d5d4a},
  {32'hc236ca30, 32'h43ece36a, 32'h4520e612},
  {32'hc3e9bdf8, 32'hc3e6a14c, 32'hc3764745},
  {32'hc382b42c, 32'h44985f91, 32'h44bd4474},
  {32'h43e87192, 32'hc549f100, 32'hc2dc1d0e},
  {32'h43521fd7, 32'h428ca377, 32'h44a3a97d},
  {32'h453b02de, 32'hc3a2be0c, 32'hc42050d5},
  {32'hc5115114, 32'hc4202022, 32'hc1e2b5d6},
  {32'h4522a088, 32'h43a7db63, 32'h43f0c165},
  {32'hc4500715, 32'hc3c6ee8c, 32'h435e76d8},
  {32'h43b6b87c, 32'h45114b73, 32'hc2403526},
  {32'hc3a47ce8, 32'hc52c2aa2, 32'h43df1a78},
  {32'hc4f4b8b4, 32'hc317dca7, 32'h429f31e4},
  {32'hc53d1b02, 32'hc3d8480b, 32'hc38330a6},
  {32'h44a130b7, 32'h4467c406, 32'h4453eba4},
  {32'h42b3ebd6, 32'hc49f2e01, 32'h420d2005},
  {32'h4445b927, 32'h440edbd4, 32'hc425eaf9},
  {32'hc3dafb84, 32'hc509ed1d, 32'hc3562765},
  {32'h42e90978, 32'h44a48040, 32'hc41bf0bd},
  {32'hc42737df, 32'hc40a0e2c, 32'h44d063b9},
  {32'h430da0a3, 32'h43dd1728, 32'h43e9aa76},
  {32'hc458156f, 32'hc30fe5f8, 32'h3f106d00},
  {32'h444d1cf0, 32'h41a604b2, 32'hc4c52361},
  {32'hc47a76c7, 32'h43d16f48, 32'h44bf96b3},
  {32'hc3cbec1d, 32'h42fdb9be, 32'hc458c37d},
  {32'hc56b334e, 32'hc391cab3, 32'hc1eeebaa},
  {32'h4318688c, 32'h44a0cebe, 32'h425e211a},
  {32'hc3da244b, 32'h42c36297, 32'h441d3b14},
  {32'h444881d2, 32'h446bccb1, 32'hc3c61740},
  {32'hc21354aa, 32'hc3e69134, 32'h44c5764c},
  {32'h440f1136, 32'hc3593fc6, 32'hc4a5c57c},
  {32'hc3c27120, 32'hc2d1a1dc, 32'h43f56383},
  {32'h45052b38, 32'hc12f82b8, 32'hc4912979},
  {32'h4533578c, 32'hc43b442e, 32'hc4054245},
  {32'hc490c163, 32'h43649f9b, 32'h444805fd},
  {32'h43a52ac8, 32'h43870208, 32'hc125367e},
  {32'hc30ebfb0, 32'h4542d776, 32'hc3599558},
  {32'h44cb0275, 32'hc424a4d9, 32'hc35c6e7a},
  {32'h44bf49b6, 32'h4369c3af, 32'hc20fcd7a},
  {32'h456fef24, 32'hc39bb470, 32'hc3b81303},
  {32'hc543e6e2, 32'h43d02b91, 32'hc2e8c946},
  {32'hc4b266e6, 32'hc3087638, 32'hc37c33b4},
  {32'hc5229ee4, 32'hc422c5d6, 32'h434c406f},
  {32'h429ba5c2, 32'hc45a75e9, 32'h449d809f},
  {32'h434d1544, 32'h43c63950, 32'hc3650cf5},
  {32'h42ea842a, 32'h427df4f7, 32'h44deaeb1},
  {32'hc3e415a4, 32'h42dfce5d, 32'hc4dde6b9},
  {32'h4358f83c, 32'hc2389066, 32'hc19488b4},
  {32'hc40ac80a, 32'hc3052c16, 32'hc48a36c9},
  {32'h452de73c, 32'hc2ed6554, 32'h4343679c},
  {32'hc4927578, 32'h432307ca, 32'hc3f9e780},
  {32'h44814b1c, 32'hc4752f6d, 32'h44dc27ec},
  {32'hc4602b7e, 32'h44ddcba9, 32'hc3afc221},
  {32'h40af4a00, 32'hc33d3996, 32'hc3524863},
  {32'hc407a4fd, 32'h43631d8e, 32'hc528c11c},
  {32'h44ad3fe0, 32'h41c734a4, 32'h44046745},
  {32'h433de337, 32'hc29127dc, 32'hc4a2e6f3},
  {32'h44142f77, 32'h44750874, 32'h45181e0e},
  {32'hc4d2c0db, 32'hc46837b1, 32'hc411f567},
  {32'hc4e8643a, 32'hc36896b0, 32'h4326e40c},
  {32'h43c025c5, 32'h44c5278d, 32'hc48b8fe6},
  {32'hc3c4bad3, 32'hc4b41c49, 32'h44c16404},
  {32'hc361e6ec, 32'h44b326cc, 32'hc458bc3d},
  {32'hc43ab9e3, 32'h422876aa, 32'hc30a9096},
  {32'h42a09f68, 32'hc251ae65, 32'h4532f9f3},
  {32'h43254d10, 32'h452a66c3, 32'h43d3f9b8},
  {32'hc4df2bc7, 32'hc2c872a3, 32'h4281522a},
  {32'hc44ed656, 32'h44b3dcea, 32'h437ec23c},
  {32'h429d06cc, 32'hc52eb953, 32'h43c24746},
  {32'h444a42da, 32'h44cdb82e, 32'h447365c8},
  {32'h439088bc, 32'hc408693f, 32'hc4e6be9f},
  {32'hc29632f1, 32'hc336fda1, 32'h4402f0f8},
  {32'hc4678101, 32'hc28919f7, 32'h43c0dd1b},
  {32'hc402c756, 32'h4399d3a4, 32'hc3f323a6},
  {32'h42a4c3b0, 32'h43a9fda1, 32'h4515355a},
  {32'hc4b8eb2e, 32'h43cd8990, 32'h442dda6d},
  {32'h444de707, 32'hc488acf2, 32'h444de1b3},
  {32'hc426ba50, 32'h4380d653, 32'hc4d049b4},
  {32'h456524fa, 32'hc3e02d3a, 32'hc3a54696},
  {32'hc518a653, 32'h43d092af, 32'hc3b8fc0e},
  {32'h4581bab1, 32'hc2da58d2, 32'hc42b3398},
  {32'hc31112d7, 32'h44f2632d, 32'h42f9833f},
  {32'h44762518, 32'hc48dd9a2, 32'h420e490c},
  {32'hc5119c3e, 32'h43374690, 32'h3f8061e0},
  {32'hc4b097a9, 32'hc3aa4692, 32'h40e81107},
  {32'hc406d037, 32'h454cd05c, 32'hc2ca445d},
  {32'h45397750, 32'hc41860fe, 32'hc3f48c10},
  {32'h4289c1c2, 32'hc31a3e42, 32'h43d87714},
  {32'hc3b25f11, 32'h44bd665a, 32'hc507f8a1},
  {32'hc3b9ee58, 32'hc4920f54, 32'h44fdf3ae},
  {32'hc48827cf, 32'hc393e874, 32'h4309be9d},
  {32'h4497f46c, 32'h4338eb9c, 32'hc36b455c},
  {32'hc3661895, 32'hc3bf8192, 32'h44a9997c},
  {32'h43de5348, 32'h44f46046, 32'hc3fd0e95},
  {32'hc42c15b9, 32'hc2d7eb17, 32'hc09516d0},
  {32'hc503cc03, 32'hc4042b32, 32'hc2996a4d},
  {32'hc44b270c, 32'h428b8eb1, 32'hc41784ab},
  {32'hc3f34a91, 32'hc51be5fc, 32'h44a962e3},
  {32'hc0de2140, 32'h441bfe8a, 32'hc4e6bdf4},
  {32'h43339b18, 32'h424b9642, 32'hc53e8f55},
  {32'hc39e6c1e, 32'hc4532d78, 32'h44340a51},
  {32'hc15adb80, 32'hc3968f12, 32'hc460e538},
  {32'hc49c5926, 32'hc3f673c9, 32'h44853b82},
  {32'h435b73bc, 32'h44fcc9a3, 32'hc3d2e29c},
  {32'h43c65afa, 32'hc45057a7, 32'hc1100f59},
  {32'h45522e92, 32'hc36d6995, 32'hc09b3269},
  {32'hc41f188e, 32'hc3d774ab, 32'h4450fcea},
  {32'h4566ad39, 32'hc2bbd294, 32'h43ad6bf8},
  {32'hc2c4747e, 32'hc58062ac, 32'h430ffa73},
  {32'h446bc55e, 32'h43f94d86, 32'hc404d879},
  {32'hc4643a5a, 32'hc3866eb4, 32'h4420fc56},
  {32'h435074c6, 32'h44fcacec, 32'hc2aad71a},
  {32'hc444d5fa, 32'hc4ed40e7, 32'h4378cdfb},
  {32'h44c469fb, 32'h44015e7f, 32'hc2a34109},
  {32'hc4405702, 32'h43e49027, 32'hc3aea42c},
  {32'hc47aa106, 32'hc3821799, 32'hc364f998},
  {32'h418db980, 32'hc4e6584c, 32'h44f0fc44},
  {32'hc30eb3d6, 32'hc2018fe6, 32'hc4ae7f89},
  {32'h44ab305e, 32'h4373ef8b, 32'h4411ee16},
  {32'hc4a11033, 32'hc3d6f0ea, 32'hc400b751},
  {32'h44268017, 32'h43775fbe, 32'hc38485c8},
  {32'hc4953438, 32'hc407d025, 32'hc406521f},
  {32'h445ac545, 32'hc1fc124e, 32'h44823a0e},
  {32'h43db4799, 32'hc213451c, 32'hc31c2b2b},
  {32'hc3322491, 32'h4429cb4d, 32'h438cc49d},
  {32'h42c03c28, 32'h44f68111, 32'hc4cc24f8},
  {32'hc37fa2b8, 32'h44703fb6, 32'h43664940},
  {32'hc44c4d2e, 32'hc261d89c, 32'hc441271c},
  {32'h44490f7a, 32'h440d41df, 32'h44d96e59},
  {32'hc28624e8, 32'h42f26c9b, 32'hc4bab912},
  {32'h4413c832, 32'h44821685, 32'h44304e03},
  {32'hc4a913de, 32'hc38ae738, 32'hc43319a5},
  {32'h44c19c9b, 32'h42927f47, 32'h4356c598},
  {32'hc4c2f966, 32'hc49c8f57, 32'hc375833d},
  {32'h43d8ae4c, 32'h4533cfbf, 32'hc34078e3},
  {32'h44041106, 32'hc4d2e306, 32'hc3284192},
  {32'h4345c1dd, 32'h455f583d, 32'hc29673f5},
  {32'hc3afbb5e, 32'hc54febb7, 32'hc4122479},
  {32'h455c782f, 32'h43cdf81e, 32'h43c52dd7},
  {32'hc4fa1223, 32'hc39cd9f0, 32'hc3c44550},
  {32'h44f4674a, 32'hc269232d, 32'h43b2d08b},
  {32'h4417eb6c, 32'hc54e679e, 32'hc3b4922c},
  {32'hc5376a04, 32'h42929197, 32'h4346234e},
  {32'hc3b7f586, 32'hc457b6ba, 32'hc2933a81},
  {32'hc416f572, 32'h43eff8c6, 32'h4513f67b},
  {32'h4452f08e, 32'hc400cd35, 32'hc3c20196},
  {32'hc3cc0763, 32'h4371c2c5, 32'h44f6ca17},
  {32'hc2d43a45, 32'hc3fd1de3, 32'hc541e68a},
  {32'hc4b8efdd, 32'h44b103b9, 32'h4486c6d5},
  {32'hc1601580, 32'hc3c26bd4, 32'h43d9630e},
  {32'h440f3622, 32'hc410a7ce, 32'h4414f18a},
  {32'hbe473800, 32'hc361040a, 32'hc4b3cfb3},
  {32'hc3208dde, 32'hc3d3ef03, 32'h44575a6d},
  {32'h443b57ac, 32'hc31c9d57, 32'hc34b7212},
  {32'hc44b63ed, 32'h44552d6a, 32'h4451e3a4},
  {32'hc2b387a0, 32'hc4a0e0d4, 32'h4352d72e},
  {32'hc4b6fdc7, 32'h43455d8d, 32'h449de027},
  {32'h409ebca0, 32'hc43e9179, 32'hc484163a},
  {32'h4464ca71, 32'h429d2e2c, 32'h43a222b9},
  {32'h4412f710, 32'hc4f19314, 32'hc355454c},
  {32'hc3b850ac, 32'h454c529e, 32'h43495c8c},
  {32'h42f39ccc, 32'hc4deface, 32'h42684b2a},
  {32'hc52e66c2, 32'h42cc2e80, 32'h42c93679},
  {32'h454f1350, 32'h436100ca, 32'hc2e21b35},
  {32'hc51c7d67, 32'h438331da, 32'h438d7574},
  {32'h44c9e4de, 32'hc3277c6a, 32'hc2185163},
  {32'hc53a9d67, 32'h44256f32, 32'hc20c334e},
  {32'h4537482e, 32'h42a9701b, 32'h4287feed},
  {32'h44ec600c, 32'hc223f28f, 32'h42e1e654},
  {32'hc5214186, 32'hc39d2ef6, 32'h4325ca48},
  {32'h44c89300, 32'h43b6b2ae, 32'h44aac4c0},
  {32'hc4a8530e, 32'h43991f9e, 32'h432c1602},
  {32'h43eb27d4, 32'hc4c584e0, 32'h43b74e06},
  {32'hc3c87708, 32'h44ca537b, 32'h438b92ff},
  {32'hc389caee, 32'hc421ece4, 32'hc428db40},
  {32'hc4a4d30a, 32'h44accdf5, 32'hc3f6019a},
  {32'h43facbef, 32'hc4d5caae, 32'h421111d8},
  {32'hc4c9c4d7, 32'hc3334c1f, 32'h43a3ca6f},
  {32'h4414ef92, 32'h4296275b, 32'h44eb73e0},
  {32'h42a54400, 32'h43a5f651, 32'hc5422262},
  {32'h44c8e98e, 32'h420e56f0, 32'hc38fba32},
  {32'hc35f0a0c, 32'hc1823a6d, 32'h4486520e},
  {32'h43a01b0c, 32'hc3a13dbb, 32'hc50ec334},
  {32'hc50c9653, 32'h426fb026, 32'h42f9139e},
  {32'hc1e2b434, 32'hc52aff9a, 32'h43779970},
  {32'hc34352df, 32'h44ed0f42, 32'hc375f4c7},
  {32'hc495aabd, 32'hc3527b14, 32'hc39c571d},
  {32'hc51aaf13, 32'hc46e6fe4, 32'h40c36000},
  {32'h448bf096, 32'hc310ae89, 32'hc46ac20e},
  {32'hc3e76e49, 32'h4405a503, 32'h43add88f},
  {32'h43b15adc, 32'hc4239272, 32'hc47997dd},
  {32'hc4c06bf2, 32'h44836f2b, 32'hc3803ca4},
  {32'h45566b55, 32'h41ce41fd, 32'h41c9070e},
  {32'hc4b8f6a9, 32'h4486233c, 32'hc3ab4394},
  {32'h43d0c3b4, 32'hc4dc3599, 32'hc3983c8e},
  {32'h4469f760, 32'hc3383526, 32'hc4e2981e},
  {32'hc4006128, 32'h4321194c, 32'h43928560},
  {32'h44ed9546, 32'h423bfc92, 32'h42bcebda},
  {32'hc3a7768f, 32'hc5396b96, 32'hc190d3fb},
  {32'hc2cf201c, 32'h45279a94, 32'h43585263},
  {32'h44f18881, 32'hc28edacc, 32'hc3392fee},
  {32'h44ab5734, 32'h44c87b47, 32'h430fe4a5},
  {32'hc4c029b9, 32'hc4905caa, 32'h43c262fc},
  {32'hc2063f3e, 32'h416cc456, 32'h43e88270},
  {32'hc4af2cdb, 32'hc413520a, 32'hc11c56d0},
  {32'h447945b0, 32'hc242a7e5, 32'h41fc2446},
  {32'hc2e7a896, 32'h4272461a, 32'h448da83b},
  {32'h42a5bf35, 32'h440752ed, 32'h4537718a},
  {32'hc408f1ba, 32'hc4eef8ad, 32'h432b154c},
  {32'h444c3766, 32'h427b14af, 32'h43aed6b2},
  {32'hc4d1dd2e, 32'hc33f88bd, 32'hc453c9b3},
  {32'h449c603e, 32'h44817dfa, 32'h44199f02},
  {32'h44d39dd5, 32'hc3f719d9, 32'hc3a4b469},
  {32'h44f66ff8, 32'h4452e094, 32'h4493b11d},
  {32'hc567f09d, 32'h43444d86, 32'h42e6a857},
  {32'h44ecefcc, 32'h44545fa8, 32'h431c8257},
  {32'hc505f06c, 32'h4379fd86, 32'hc4631284},
  {32'h42bd79fc, 32'h451fb4f9, 32'hc3252292},
  {32'h43988584, 32'h424fa282, 32'hc4394da4},
  {32'h4174f970, 32'h44339de5, 32'h45437f39},
  {32'h43b5b2d8, 32'hc46d8b09, 32'hc4b8d899},
  {32'hc285f686, 32'h446b6aef, 32'hc338f887},
  {32'h45162aee, 32'hc42ef8b4, 32'hc3bb1588},
  {32'hc4906384, 32'hc43fed3e, 32'hc300481d},
  {32'h44baaffd, 32'h4434011d, 32'h42ad5f95},
  {32'hc4dfb7be, 32'hc37b8282, 32'h4288d832},
  {32'h43fb55ad, 32'h43022a9b, 32'h44157e6c},
  {32'h4306fb91, 32'hc5254bb0, 32'h4355c2a9},
  {32'h45526ea9, 32'h431538d8, 32'h429bc30e},
  {32'hc5153c61, 32'hc41b8f03, 32'hc3765e24},
  {32'h440eed72, 32'hc356439b, 32'hc2c26dbe},
  {32'h44266ce6, 32'hc4ca0edf, 32'hc2c48c94},
  {32'h438cb8c4, 32'h44956c88, 32'hc324d4e5},
  {32'hc400620e, 32'hc4e27625, 32'hc2249ec6},
  {32'hc3552725, 32'h431de25b, 32'hc44b4c9d},
  {32'hc4afab12, 32'hc3a1959f, 32'h441549ad},
  {32'h44d8716c, 32'h4480c9c0, 32'h423e6465},
  {32'h42b468e0, 32'h3fd872f8, 32'hc2a53eec},
  {32'h4413f4bc, 32'hc303cc7a, 32'hc2948532},
  {32'hc4f3acdc, 32'h431993a4, 32'h43a54535},
  {32'hc48cd7e0, 32'h43ca2049, 32'hc42c10fb},
  {32'hc431a0b3, 32'hc512002e, 32'hc31fc541},
  {32'h441dcc54, 32'h44a0e37b, 32'h422c18f0},
  {32'hc36efbaa, 32'h42025311, 32'h43ad471a},
  {32'h448a3adf, 32'h44915875, 32'hc4250520},
  {32'hc4410ebb, 32'hc533c3f7, 32'h43d1c2da},
  {32'h41c5dfbc, 32'h4291ab31, 32'hc22ecf53},
  {32'hc53d7e5b, 32'h43def731, 32'h43baae2c},
  {32'h4485ca70, 32'hc35eccf7, 32'hc50770cd},
  {32'h450e09da, 32'hc3ce420c, 32'hc409f3af},
  {32'h43669312, 32'h4537f428, 32'h429f5b8e},
  {32'hc4d7a1b3, 32'h430f4a0b, 32'hc2151d21},
  {32'hc40884f3, 32'h450c2fad, 32'h437e6ca1},
  {32'h44548858, 32'hc4326490, 32'h440f8f73},
  {32'h43e78f1c, 32'h4518ee41, 32'h42fe2c31},
  {32'h45225fe4, 32'hc4130f1f, 32'hc30df376},
  {32'hc5813978, 32'h4285eb4e, 32'h441a9249},
  {32'hc452772a, 32'hc34b15df, 32'h41dc5505},
  {32'h43d05256, 32'h44afd8c3, 32'hc32c21ca},
  {32'h44c2d402, 32'hc40c4c70, 32'h43bcf72d},
  {32'h4366ade0, 32'hc388f5de, 32'hc3c6cf66},
  {32'h42ab6a8b, 32'h43d87545, 32'h44733df3},
  {32'hc3691720, 32'h452ec9f4, 32'hc186bb04},
  {32'hc32e4446, 32'hc4bc8aa2, 32'hc306b825},
  {32'hc269e420, 32'hc389dcc4, 32'hc46ec587},
  {32'h44ae8190, 32'hc3bacbb8, 32'h440e1f5d},
  {32'hc504fccc, 32'hc33d846c, 32'h422339a3},
  {32'h442c0824, 32'hc3fda1a4, 32'h44e1bdbb},
  {32'hc54bbd25, 32'h439ee31a, 32'hc42742d2},
  {32'hc394a5dd, 32'hc4252246, 32'h4348ae42},
  {32'hc4540f2e, 32'h4379ec4b, 32'hc3e88362},
  {32'hc36641ef, 32'hc4f0c1ac, 32'h443a5d52},
  {32'h43d813ce, 32'hc3b3696c, 32'hc479143a},
  {32'h4182d400, 32'h4405de3c, 32'h448cce2b},
  {32'hc4d161d8, 32'hc40be60a, 32'h421d17ba},
  {32'hc30e3874, 32'h43622d1c, 32'h4452cb62},
  {32'hc3a46f92, 32'h43ede6ef, 32'hc48a61b9},
  {32'h423182e0, 32'h44e571f2, 32'h44bc248b},
  {32'hc505e922, 32'h429b4d88, 32'h44021f0b},
  {32'hc3ed87d8, 32'h4342349d, 32'hc4952ad8},
  {32'h4365a211, 32'hc501ec27, 32'hc35a2e85},
  {32'hc3432f50, 32'h43ca54cd, 32'hc4273f21},
  {32'h4509be01, 32'h43ab9e62, 32'hc2601c9b},
  {32'hc3ec7128, 32'h4426a40c, 32'hc485ee37},
  {32'h451c5192, 32'hc3a57bbd, 32'h4420be11},
  {32'h450f400e, 32'hc3d8900b, 32'h442f9585},
  {32'hc54c0cdf, 32'h42845ff3, 32'h43361291},
  {32'h428997da, 32'h448db2ca, 32'h43aade7a},
  {32'h4513e751, 32'h442c3795, 32'h43083250},
  {32'hc55691c8, 32'hc26c8918, 32'hc3bbabb8},
  {32'h45003e4f, 32'h43b5b165, 32'h42bb4a7e},
  {32'h4488d5a4, 32'h431c93cd, 32'hc440fd87},
  {32'h430dd6d7, 32'h437ec4f2, 32'h452bedea},
  {32'hc5147ff6, 32'h430816a3, 32'h428ed3f3},
  {32'h449712dc, 32'hc43c401c, 32'h43348c7e},
  {32'hc521eb88, 32'hc36cc476, 32'hc431fd8e},
  {32'h433ddb00, 32'h434ad594, 32'h43bbff43},
  {32'hc410a9e2, 32'hc3b86534, 32'hc3af251b},
  {32'h449c8f7e, 32'hc48c788e, 32'hc42bf70b},
  {32'h42030a40, 32'h440f7b3c, 32'hc1ac2426},
  {32'h4440cce4, 32'hc4abdc70, 32'h428157bc},
  {32'hc22065c0, 32'h44c404aa, 32'h4312b71d},
  {32'h4494b79e, 32'hc4b4d901, 32'h439f90f2},
  {32'h43386fe9, 32'h42c3354e, 32'h442e10d8},
  {32'h4404603c, 32'hc388a4ca, 32'hc43f47ed},
  {32'h42aaaf1a, 32'hc49bb6c8, 32'h4539090a},
  {32'h41f46880, 32'hc41ffd83, 32'h44b39b9a},
  {32'h446ea08f, 32'h43a8452b, 32'hc438a999},
  {32'h44cdac86, 32'hc3f63ead, 32'hc3b7122e},
  {32'h4477da9e, 32'h449f9251, 32'hc412e57e},
  {32'hc4285872, 32'hc4d4b110, 32'h43ce3f63},
  {32'hc4cc3d04, 32'h43141fc1, 32'hc39472bc},
  {32'h429f7ab0, 32'hc38da034, 32'hc3bae3b2},
  {32'h43f2fad8, 32'hc47cf87a, 32'h453b550d},
  {32'h446d78b1, 32'h442aeb35, 32'hc43f85c5},
  {32'h44196808, 32'h45102d63, 32'hc2d4f878},
  {32'hc487dfe2, 32'hc3bcb708, 32'h4423280a},
  {32'h44f6a01a, 32'hc3aa76a3, 32'h43652b44},
  {32'hc4d46e79, 32'hc3710994, 32'h4485ad86},
  {32'h44885c61, 32'h413c19a8, 32'h435bca62},
  {32'h44995814, 32'hbfa240f1, 32'h4323893e},
  {32'h445cf055, 32'h421049f6, 32'hc3f8fba9},
  {32'hc43d938e, 32'h44481568, 32'h42de2da2},
  {32'h4573c248, 32'h43dac9ff, 32'hc297f56b},
  {32'h43803878, 32'hc5406c50, 32'hc2957084},
  {32'h44566ebb, 32'h44b87f86, 32'hc28ee4ce},
  {32'h4475edb2, 32'hc41ae202, 32'hc2d296a7},
  {32'h42d996e0, 32'h4520a271, 32'h41e4bdda},
  {32'hc4b3865f, 32'hc4015696, 32'hc2e67686},
  {32'hc3ebc116, 32'h43baf2db, 32'h437756b9},
  {32'h42cd4414, 32'h44b1a9cd, 32'hc3072a6a},
  {32'hc3db50b0, 32'hc4bc27f9, 32'hc421a67d},
  {32'hc46ab709, 32'hc49b6180, 32'h4496728a},
  {32'h45010b5c, 32'h41df628c, 32'h42c67634},
  {32'h447b7669, 32'hc39f969c, 32'h44775f7b},
  {32'h440116cf, 32'hc4b36f3e, 32'hc4129704},
  {32'h45167b46, 32'h43de2619, 32'hc3c9b8c7},
  {32'hc41b1b84, 32'hc4727378, 32'hc4c94c38},
  {32'h440e9ed1, 32'h44b14b20, 32'h448ee10c},
  {32'hc3fcc016, 32'hc407136f, 32'hc3157536},
  {32'h42eafc3c, 32'h43eddff2, 32'h449c93ba},
  {32'hc2c196d1, 32'hc52c9866, 32'hc4124808},
  {32'h4437e32c, 32'hc212fa7a, 32'h44e89831},
  {32'hc49d03ba, 32'hc449754b, 32'hc3fe6e80},
  {32'h44288804, 32'hc203d1d4, 32'h4477785e},
  {32'hc4bb2e41, 32'hc3a71380, 32'h436a9673},
  {32'h449adccc, 32'h440e98a2, 32'h44b0a155},
  {32'hc349cf00, 32'hc505b8c9, 32'hc4dfb74c},
  {32'h44dd76c6, 32'hc306f6a0, 32'h43ec8291},
  {32'hc4bcbab4, 32'hc482a0dd, 32'hc318d6c6},
  {32'h423997d4, 32'h4557f3b9, 32'h43905d72},
  {32'h44d595b1, 32'hc1aff6af, 32'h3f7b5b44},
  {32'hc20c2839, 32'h45198123, 32'h441fe003},
  {32'hc4a3ddb2, 32'hc3990260, 32'hc32aaee4},
  {32'hc4d4ad44, 32'h434abf5a, 32'h432aef54},
  {32'hc4f07045, 32'h41e4d145, 32'hc311f3b0},
  {32'h44c25492, 32'h42c458b0, 32'hc346d1d2},
  {32'hc20755b7, 32'hc56fa6db, 32'hc310e850},
  {32'h41cde502, 32'hc4f337f9, 32'h44f1dc2c},
  {32'hc31772fd, 32'hc2577d9a, 32'hc3fa14e0},
  {32'hc3e4010b, 32'h44f85d9b, 32'hbea46b30},
  {32'h447e8fa9, 32'hc4a1d4ca, 32'hc40d5689},
  {32'h44a7a8ef, 32'h42f12a9c, 32'h43abb6a2},
  {32'h43644658, 32'hc4564dbc, 32'hc4edf8c1},
  {32'hc52e321a, 32'h433e73dd, 32'h43eaf648},
  {32'h4403abc6, 32'hc406f4e8, 32'hc376d8d0},
  {32'h438a85b0, 32'hc49ce0ad, 32'h44cc0f02},
  {32'hc23e3a0b, 32'h440a5b37, 32'hc4c23dcb},
  {32'hc3b6c19a, 32'h42111c1c, 32'h4486407b},
  {32'h422dab94, 32'hc4d610de, 32'hc42492ec},
  {32'hc562e121, 32'hc38d0b21, 32'h432014e5},
  {32'h41a03d81, 32'hc2424640, 32'hc4929d6a},
  {32'hc4a808ce, 32'h4408534d, 32'h44529624},
  {32'h43f3d7c3, 32'h4364d731, 32'hc48ca916},
  {32'hc42b8100, 32'h4335dfe8, 32'hc453356c},
  {32'h44436970, 32'hc4b14723, 32'h42847b28},
  {32'hc4dece26, 32'h42ed154f, 32'h436f84b1},
  {32'h451a686c, 32'h444b1b72, 32'h435c7306},
  {32'hc4a94b77, 32'h439af7d4, 32'hc402ab35},
  {32'h4318ac22, 32'hc56c465d, 32'hc374f7ba},
  {32'hc509361a, 32'h430bc9b9, 32'h43a69ac8},
  {32'h446dbbce, 32'h439a5eb4, 32'hc2a8a494},
  {32'hc4543890, 32'hc11248d8, 32'hc3409c0c},
  {32'h447f183e, 32'hc2af9cb5, 32'hc3bed005},
  {32'hc4000be3, 32'h43509ffa, 32'h43a57b7c},
  {32'hc4810dc6, 32'hc3aa7e78, 32'hc4f3bdf8},
  {32'h446b9d76, 32'h4296711e, 32'h452f5882},
  {32'hc518d9f4, 32'h433ffa17, 32'h42b7fc50},
  {32'h442bc828, 32'hc5188834, 32'hc3b54e70},
  {32'hc48391ce, 32'h439022b2, 32'hc3da7136},
  {32'h43e7bced, 32'h4307d2d7, 32'h439ff374},
  {32'hc4a5bbf7, 32'h44aaffbf, 32'h4381cb9a},
  {32'hc284a240, 32'hc4a4aba6, 32'h42b158e0},
  {32'hc4b9ef22, 32'hc33202c3, 32'hc42d5a8b},
  {32'h42b5d090, 32'h4367223b, 32'h44eb2054},
  {32'hc50a0ac6, 32'h43310aca, 32'h44079c40},
  {32'hc4a52fc6, 32'hc39a2286, 32'hc2dad95c},
  {32'hc48ff0ef, 32'h44a4a3b5, 32'h43d9a7b1},
  {32'h44ea7038, 32'hc3b5320a, 32'hc38c67a6},
  {32'h449c499c, 32'h4204c624, 32'h4391b433},
  {32'h452b1a73, 32'hc3a027b6, 32'hc33b9c72},
  {32'h418dda60, 32'h449d6bfe, 32'h443fd80d},
  {32'h4532f82b, 32'hc2b2a20b, 32'hc345c078},
  {32'hc4b1c9e6, 32'h44a36c64, 32'h448d2d2b},
  {32'h44ec1cbe, 32'h42785d9f, 32'hc47abccc},
  {32'hc4657f04, 32'h43678553, 32'hc2a509b5},
  {32'h43a844d7, 32'hc50815ca, 32'hc4371941},
  {32'hc2a134e0, 32'h44cc5e62, 32'h432eff41},
  {32'hc4ca47cd, 32'hc3238ec2, 32'hc40e37e3},
  {32'hc40299d3, 32'h439593c8, 32'hc209c870},
  {32'h436f28e0, 32'hc4d451c1, 32'hc39db076},
  {32'h43c484f0, 32'hc3037041, 32'hc4b14c0b},
  {32'hc4201086, 32'hc35d69cf, 32'hc3496474},
  {32'h44528fb6, 32'h43ebca6e, 32'hc2fece92},
  {32'hc4a74e7c, 32'hc4b030af, 32'hc3c9786d},
  {32'h455b07c8, 32'hc39c8a54, 32'h42c34ccd},
  {32'h445b1a43, 32'hc311924e, 32'hc2c7c7b6},
  {32'hc140c5c0, 32'h457913d3, 32'h42cb28d0},
  {32'hc494a442, 32'hc440f6cb, 32'h44001e20},
  {32'h4422c73a, 32'h43e4234c, 32'h440a3cec},
  {32'hc4f88e2e, 32'h43a4e8e3, 32'h443001ce},
  {32'h45176d96, 32'h4072a339, 32'hc436898f},
  {32'hc42700f6, 32'hc2b35d08, 32'h4501d7e9},
  {32'h421d9780, 32'h4450b804, 32'h445cc86e},
  {32'hc493ad92, 32'hc36007c6, 32'hc3590687},
  {32'hc44a04ea, 32'hc2b0e935, 32'h4496ef8f},
  {32'h421e2450, 32'h4314d2fc, 32'hc471e9e3},
  {32'h43cde7cb, 32'h452e3cde, 32'hc2f92d85},
  {32'hc47be362, 32'hc48f7772, 32'hc44004c5},
  {32'h45283e17, 32'h442eddb2, 32'h4436bec2},
  {32'hc4a19e62, 32'h43041e47, 32'hc4af89ee},
  {32'h44cd2a2a, 32'hc39d8a6c, 32'hc3c0d9fe},
  {32'hc40774d8, 32'hc422e44d, 32'hc40ca18d},
  {32'hc0a44f44, 32'h44a11bff, 32'hc36e85f1},
  {32'hc3a28e7e, 32'hc440ec0a, 32'hc3f536a4},
  {32'h44b4871c, 32'h442d6383, 32'h444e4c8e},
  {32'hc47064d5, 32'h43447e38, 32'hc3b6879e},
  {32'h42a0a76d, 32'h44cfeb63, 32'h43c3d476},
  {32'h4282cb3c, 32'h443e5b31, 32'hc40ef8a7},
  {32'hc43eaade, 32'hc49639c8, 32'h439f05c0},
  {32'h448bd491, 32'h44977b3f, 32'h44149872},
  {32'hc50874a9, 32'hc384ce06, 32'h44132235},
  {32'h450e6431, 32'h43a9a020, 32'hc3c2e222},
  {32'hc1ea4a80, 32'hc52db784, 32'h42c14e22},
  {32'hc4926805, 32'h43f8a4c8, 32'hc3b9cfc0},
  {32'hc4c45c48, 32'h43dfef94, 32'hc35395be},
  {32'h44d33091, 32'hc411c2ef, 32'hc3d6dab7},
  {32'hc485e268, 32'hc25df26b, 32'h434c087a},
  {32'h43a47b6e, 32'h4466558d, 32'hc29ca593},
  {32'hc2a0ad02, 32'hc44ba84b, 32'h4454b9a6},
  {32'h42c14b68, 32'h434a3790, 32'hc4787418},
  {32'hc3883130, 32'hc4f5ec2e, 32'h442d14ca},
  {32'h4485f0b0, 32'h44a6e804, 32'hc341211e},
  {32'h443f2735, 32'hc355e17a, 32'h4447933a},
  {32'h44b5363f, 32'hc415b402, 32'hc41d6e6f},
  {32'hc48f66aa, 32'hc2e26cf7, 32'h4415640b},
  {32'hc490ba45, 32'h4418d395, 32'hc2be387f},
  {32'hc3c27a80, 32'hc5214554, 32'hc3b72cad},
  {32'h44802d0e, 32'h43ba618a, 32'hc4c0f7db},
  {32'hc4efc292, 32'hc2599932, 32'h4196f040},
  {32'hc2ad8190, 32'h4396e454, 32'hc509b4c5},
  {32'hc3f64965, 32'hc3ee527c, 32'h444db657},
  {32'h45432ca4, 32'h43a9db80, 32'h3ff30200},
  {32'hc54174d8, 32'h426fe2f6, 32'h446478ad},
  {32'h42966310, 32'hc4477101, 32'hc4b34488},
  {32'h44ac2bf2, 32'hc4818b84, 32'hc335dd23},
  {32'hc47c8dbd, 32'h4220eef8, 32'h4441ed1b},
  {32'hc481d23c, 32'hc3f9eff4, 32'h437f8de4},
  {32'hc424e422, 32'h44d88e9a, 32'h43ae4fce},
  {32'h441990af, 32'hc5031425, 32'hc28e1c64},
  {32'h43abef98, 32'h44a0d86e, 32'h430c0746},
  {32'h42e22440, 32'hc405d51a, 32'hc38b176d},
  {32'hc493bf97, 32'h43d86107, 32'h437142c0},
  {32'h454f3f1b, 32'h43ace828, 32'h4429abb3},
  {32'h43ec3f40, 32'h448d69f6, 32'hc4136042},
  {32'h445325b4, 32'hc44d5dcb, 32'h44133fb3},
  {32'h44918f8d, 32'h44721fa4, 32'hc3a844d9},
  {32'h4067c320, 32'h4351a6bb, 32'h45446601},
  {32'hc350c18b, 32'hc2f3296c, 32'hc5245590},
  {32'hc41ccc0b, 32'h42fd03c9, 32'h44735c15},
  {32'hc4c745e0, 32'h43e5cf24, 32'h43c63cf6},
  {32'h42f349e6, 32'hc341b7bd, 32'h44514d53},
  {32'hc5308198, 32'hc2ed16b0, 32'hc283ac16},
  {32'h4408c631, 32'hc4dee4bf, 32'h4381a86d},
  {32'hc45f45b8, 32'h44a2dd82, 32'hc3cc4942},
  {32'h436e04f2, 32'hc40a2c39, 32'h4384cac3},
  {32'hc52355cd, 32'h442a3bae, 32'hc17a9584},
  {32'hc3a23f33, 32'hc49b08cf, 32'h44047550},
  {32'h44886d87, 32'h4407c994, 32'h43020359},
  {32'h433550b0, 32'h4007eb54, 32'h4423b79d},
  {32'hc3d9a023, 32'hc3827a6b, 32'hc5676eb5},
  {32'h4481c145, 32'hc2d46c44, 32'h4407799a},
  {32'h440d59a4, 32'hc48e0d86, 32'hc4da32ad},
  {32'h428294a8, 32'h442fe3e1, 32'h44267b9f},
  {32'hc3e2b5dc, 32'h43ed8018, 32'h4285ae9e},
  {32'h43e92076, 32'h43e0109f, 32'hc4992f48},
  {32'h453246a4, 32'hc2c93c84, 32'h43b9196c},
  {32'hc4c49908, 32'h402075f1, 32'hc43c0e37},
  {32'h446c57cc, 32'hc33ef4b5, 32'h42ba13a4},
  {32'hc4ad00a0, 32'h4484792d, 32'hc40b9a6d},
  {32'h4406b34f, 32'h42e45914, 32'h43de4355},
  {32'h444a589e, 32'hc45bfd9d, 32'h44b56210},
  {32'h41cdfb3a, 32'hc1480787, 32'hc4c2d04a},
  {32'h44bef760, 32'hc3ab6209, 32'hc381a3b9},
  {32'h43e6f38a, 32'h4338100a, 32'h444ac226},
  {32'hc2d79026, 32'h444782c8, 32'h42ac31ae},
  {32'h42ba9798, 32'hc50b3512, 32'hc405fc7c},
  {32'h43fb291d, 32'hc3f171e5, 32'hc4f37a5d},
  {32'h43b30eee, 32'hc3e0c3db, 32'h448730ae},
  {32'h43e2baa8, 32'h43fbc9cb, 32'hc43d7b0c},
  {32'h453e24e6, 32'hc42b2b14, 32'h433dd417},
  {32'hc53a1a24, 32'hc33c483f, 32'h4360ca06},
  {32'h4498bba5, 32'h43d747e7, 32'hc2c10180},
  {32'hc44944d3, 32'h444b8c7c, 32'h441036c0},
  {32'h45015129, 32'h439d39c9, 32'h43dcb4a3},
  {32'h4252e780, 32'h45457718, 32'h4397ac59},
  {32'h455135aa, 32'h439085df, 32'h41f752c7},
  {32'hc4d854c0, 32'h44aef148, 32'h4417eeae},
  {32'h43fe2cb4, 32'hc5179348, 32'hc371d8c3},
  {32'h4401a198, 32'hc318f778, 32'h44b3ebe6},
  {32'h450e8a71, 32'h437c44ba, 32'hc2f4a1fc},
  {32'hc3e120a5, 32'h44dc97b0, 32'h449e13bc},
  {32'hc3c781d0, 32'hc44e1a6b, 32'h43d9f839},
  {32'h43b84d38, 32'h448656c6, 32'hc33601e5},
  {32'hc1890e38, 32'hc3365c5a, 32'h44fb779a},
  {32'h43891219, 32'h44f90a97, 32'hc3121cbb},
  {32'h420aa3dc, 32'hc456f225, 32'h447e213e},
  {32'hc4af2e6b, 32'h43f60406, 32'h40e8b635},
  {32'h43f16a0f, 32'h44c0e5a8, 32'hc3a3ccfa},
  {32'hc3a2b675, 32'h429e2851, 32'h4503321c},
  {32'h43230912, 32'h448f7640, 32'hc5000839},
  {32'h438611b1, 32'h44a7a179, 32'h42f37f65},
  {32'hc5133ab3, 32'hc3a74ad9, 32'h43f0e6dc},
  {32'h43c91f46, 32'h44344466, 32'hc49eedce},
  {32'hc3765cfb, 32'hc4ef0552, 32'h4389c64e},
  {32'h44dcddc3, 32'hc2b4793e, 32'h42c7ac17},
  {32'h44ff6b10, 32'hc38e61d5, 32'h41e73233},
  {32'h45809bab, 32'hc37beb0b, 32'h43a5d28a},
  {32'hc597f376, 32'hc2bbec6f, 32'h434b6e20},
  {32'h44234240, 32'h441cacdd, 32'hc39a3b3b},
  {32'h42c98e80, 32'hc514c1d5, 32'hc39cf77b},
  {32'h44bae0bb, 32'h43e01958, 32'hc3d1423c},
  {32'hc4637c0d, 32'hc3388d0f, 32'h42968a91},
  {32'h44d2b7f6, 32'h44b98247, 32'hc3e8f53f},
  {32'hc5456420, 32'hc37bf892, 32'h43cad40f},
  {32'h453759c2, 32'hc426cc3a, 32'hc433a2c0},
  {32'h44e2224d, 32'hc36ab637, 32'h4317ac3d},
  {32'hc304be00, 32'hc4349531, 32'hc423e34f},
  {32'hc2ee6af8, 32'hc39dbf0f, 32'h44f04a0e},
  {32'hc4ef6688, 32'h430a2698, 32'hc2cdfcf2},
  {32'hc28ca97f, 32'h42cb10d2, 32'h44d5d742},
  {32'hc4d075d4, 32'h434bc4f3, 32'hc487af45},
  {32'h4495cbc0, 32'h438c0953, 32'h43f6bebb},
  {32'h43aa239d, 32'hc4de1b9c, 32'hc52df773},
  {32'h4412c0d4, 32'h43da4ffb, 32'h45305c3d},
  {32'h44077d37, 32'hc3a2c47d, 32'hc3f367a7},
  {32'hc3fca880, 32'hc3ba6249, 32'h43ececd0},
  {32'hc3c1c97e, 32'h44d2b125, 32'hc4d37314},
  {32'h4441ffbb, 32'h41454e43, 32'h44b48aa5},
  {32'hc4e27743, 32'hc39850ba, 32'hc3d2ee1f},
  {32'h43bb81bf, 32'hc2a6aca2, 32'h451096af},
  {32'h44dafd4a, 32'hc3e835c2, 32'hc36d1895},
  {32'h45083f79, 32'h4286f27d, 32'hc2fc421f},
  {32'hc33dd5ac, 32'hc50a59a6, 32'hc5148661},
  {32'h4561bf65, 32'hc38f3707, 32'h44245bcf},
  {32'hc44f72cc, 32'hc4b74b8a, 32'hc3abeb64},
  {32'hc3b5f138, 32'h45620117, 32'h4429cf53},
  {32'hc47c8268, 32'h4387230d, 32'hc378385a},
  {32'hc18a2b40, 32'h45312484, 32'hc332d6e8},
  {32'hc4f6a97b, 32'hc36a106b, 32'h43876ae3},
  {32'h4478dee5, 32'h434c01c9, 32'h43aa4e35},
  {32'hc4630798, 32'hc4107be3, 32'h4233a202},
  {32'h42e24983, 32'hc39b181c, 32'h43ef3b1f},
  {32'hc321f344, 32'h42a2d81a, 32'hc4d82a29},
  {32'hc44bd5ca, 32'hc49da85e, 32'h44abe4ed},
  {32'h43ad12cc, 32'hc497ad68, 32'hc3dc194d},
  {32'hc324ccef, 32'h44390027, 32'hc11e9a29},
  {32'h44dbc8aa, 32'hc3b27e38, 32'hc28dc2f2},
  {32'h4339a3b8, 32'h44f54ad8, 32'h43b88b49},
  {32'h440b4ffc, 32'hc41d75f7, 32'hc4d5b00b},
  {32'h4212d674, 32'h44c304a5, 32'h4501fd4c},
  {32'h43881852, 32'hc3d5c693, 32'hc404614e},
  {32'hc34e5182, 32'h448490a8, 32'h442cfbd7},
  {32'hc25aef04, 32'h40f29fb0, 32'hc33ee4df},
  {32'hc3e99779, 32'hc487cefe, 32'h43b6ada1},
  {32'h44eaa370, 32'hc36cd13d, 32'hc3e04002},
  {32'hc40f7398, 32'h442ff091, 32'h430e7c66},
  {32'h44eac03a, 32'hc282500b, 32'hc410f5db},
  {32'hc3cb68f4, 32'h448974f2, 32'h451bd8f8},
  {32'h450f99d4, 32'h43bcff4e, 32'hc3c9db2d},
  {32'h422d2f7c, 32'hc39368ad, 32'h4461cd66},
  {32'h41f05240, 32'hc4eca1b6, 32'hc46aa369},
  {32'hc4cf9264, 32'h44535f47, 32'hc3768531},
  {32'hc3ca750f, 32'hc4d0e1af, 32'h43560272},
  {32'hc3cf1b3c, 32'h452024fe, 32'hc2017c87},
  {32'h450c882c, 32'h433a7d80, 32'h4284f706},
  {32'h4515c510, 32'h42ace2f4, 32'hc2ce016a},
  {32'h444cfc30, 32'h4449a69a, 32'hc3fe124a},
  {32'hc59e273c, 32'h433ddd59, 32'hc395efa3},
  {32'h44da3c07, 32'hc43decb5, 32'hc4276865},
  {32'h43c2d222, 32'hc42583e9, 32'hc1db17e6},
  {32'hc517a1f4, 32'hc3c6bca2, 32'hc2ce483a},
  {32'h45487963, 32'h42d99cbf, 32'h43ef9468},
  {32'h450590f7, 32'hc2f6813b, 32'hc20f7b7e},
  {32'h44e3eafd, 32'hc4bf9d17, 32'h42b71cc8},
  {32'hc3a85e1a, 32'h44df91c2, 32'h441c8738},
  {32'h44ff6dc9, 32'h439eed8a, 32'h43c79b52},
  {32'hc558f682, 32'hc163cee8, 32'h431daa75},
  {32'h4417dad5, 32'hc4d65e89, 32'hc3ff42d2},
  {32'hc2d1eab8, 32'h43be03d0, 32'hc4c8a085},
  {32'h43d64c8c, 32'hc223bc06, 32'h4409ed97},
  {32'hc51773b2, 32'hc374d487, 32'hc1c17c28},
  {32'h447409ba, 32'h430b49aa, 32'h436d0564},
  {32'hc2346ce0, 32'h43b87516, 32'h42b28a96},
  {32'h441184fb, 32'hc429669f, 32'hc50d8bd0},
  {32'hc3d89464, 32'h432c0c8c, 32'h4358f654},
  {32'hc3d62a70, 32'hc46886e4, 32'hc4966b68},
  {32'h432e6a10, 32'h451cab4c, 32'hc1bf7578},
  {32'h44fcf80a, 32'h43dc5f26, 32'hc46231d7},
  {32'hc4e73323, 32'hc4c571c6, 32'h44d1499b},
  {32'h432ea608, 32'hc400c5c3, 32'hc44e4a2d},
  {32'hc4974e1a, 32'h433d7c1c, 32'hc37c0e98},
  {32'hc2eeffd6, 32'hc53dfe83, 32'hc30476f5},
  {32'hc3c94e06, 32'h44d85622, 32'h431cc282},
  {32'hc32ffb0c, 32'h433c459a, 32'hc40a643b},
  {32'hc49e7f71, 32'h4410ca06, 32'h44b393fc},
  {32'h443545cc, 32'hc50d6e9a, 32'hc3c1e20d},
  {32'h44db04c7, 32'h43926b4d, 32'hc43ec210},
  {32'hc50adad9, 32'hc36c2224, 32'h44a2ee5e},
  {32'hc4533cf6, 32'h43e790b9, 32'hc43467cf},
  {32'hc3cdcce0, 32'hc5091c2f, 32'h4211d40c},
  {32'h444f01b0, 32'h441db746, 32'h440a7eac},
  {32'hc510dabe, 32'hc2176ee6, 32'hc360b97b},
  {32'h43562508, 32'h45604935, 32'h3e1b21a7},
  {32'hc4cccbc6, 32'hc46c6957, 32'h43d3cb5f},
  {32'h44f64d6e, 32'h433514cd, 32'h442579ee},
  {32'hc3305e88, 32'h44497b2a, 32'hc4289a4c},
  {32'h4470672e, 32'hc3472411, 32'hc40aa5e3},
  {32'hc29ee09f, 32'h40b47cae, 32'h44e9bcfe},
  {32'h43e3f069, 32'h44edfcfa, 32'h43f0037b},
  {32'h436c5fe2, 32'hc5011a3a, 32'hc39a1416},
  {32'h44c02972, 32'h42818394, 32'h42b040cd},
  {32'hc3ee315b, 32'hc4fe4543, 32'h42a49d50},
  {32'hc340cfeb, 32'h4559d7f6, 32'h43874ce2},
  {32'h44ea82d6, 32'hc4185367, 32'h433897db},
  {32'hc33bc340, 32'hc458baf6, 32'h44439e69},
  {32'hc4ba7138, 32'hc33d4673, 32'hc4089184},
  {32'hc4126bb6, 32'h4369a47d, 32'hc2b28b16},
  {32'h4416c769, 32'hc396469d, 32'hc4979309},
  {32'h4485163a, 32'hc3c4ed28, 32'h4425ecbd},
  {32'h4463001e, 32'h430659e1, 32'h429ade96},
  {32'h44c854f4, 32'h4477d9d1, 32'hc31fd8b2},
  {32'hc3ff9bf4, 32'hc4b2ef03, 32'hc42a6750},
  {32'h45132f82, 32'hc3b91b12, 32'hc3912d85},
  {32'hc4f03b20, 32'hc3c9bf47, 32'hc2ffdb2b},
  {32'hc4f77d7a, 32'h41cae182, 32'hc3c209ee},
  {32'h452be775, 32'h433d22a8, 32'h44181218},
  {32'hc509263b, 32'h441e8fab, 32'h40d65280},
  {32'h44a4fb3c, 32'hc365c8cc, 32'h42af8a2f},
  {32'hc251d5ec, 32'hc556bf16, 32'h40e3e013},
  {32'hc4296af0, 32'h4361345f, 32'hc39b272c},
  {32'hc592b315, 32'h439bb786, 32'hc306fb70},
  {32'h4568b7ae, 32'h439cc3f9, 32'h43db8047},
  {32'h43a58d42, 32'h4244f1de, 32'h448bc46c},
  {32'h4443ad60, 32'h44d05512, 32'h4217f51e},
  {32'hc4a19f4b, 32'hc40bd5dc, 32'hc3da981e},
  {32'hc4c694fe, 32'h4404b18e, 32'hc147d3e7},
  {32'hc3cc35cc, 32'hc4906efd, 32'h44621c35},
  {32'h4401d316, 32'hc20bd3a2, 32'hc44634a3},
  {32'hc2c4b8c0, 32'h426e44c2, 32'h442b117b},
  {32'h421c4370, 32'hc23cd2d2, 32'hc52eca87},
  {32'hc512a1f2, 32'hc3aa83a9, 32'hc336ee57},
  {32'h4444e50a, 32'h431fe3d8, 32'hc49dbfd8},
  {32'hc48757e1, 32'hc4c07f1d, 32'h448a5a2e},
  {32'h435aa0e0, 32'h44cfed96, 32'hc42af769},
  {32'h44d0f470, 32'h4272ebda, 32'h436c35c2},
  {32'h44693503, 32'h444f7043, 32'hc4061234},
  {32'h42835cb8, 32'hc5464d98, 32'hc2b0f02b},
  {32'hc47c8c65, 32'h43b2b47a, 32'hc3243934},
  {32'hc438f2c4, 32'h44056172, 32'h4556a114},
  {32'h44c9ef10, 32'hc36eae47, 32'hc4e6dabe},
  {32'h4520472d, 32'hc47e2adc, 32'hbe943544},
  {32'hc1690700, 32'h4501ed09, 32'hc2240aac},
  {32'h450f625a, 32'h424067f8, 32'h43c94543},
  {32'hc518a824, 32'h449c72fa, 32'hc3eee5ca},
  {32'h441aeab4, 32'hc4504be8, 32'h4212dd30},
  {32'hc4846cb7, 32'h443ce5cf, 32'hc3e6f1cd},
  {32'h44d906e8, 32'hc4ad0fb5, 32'hc480f524},
  {32'hc40d2440, 32'hc4293f7b, 32'hc39fa756},
  {32'h45534a4c, 32'hc28a4943, 32'h4411e2fb},
  {32'hc493982c, 32'h43302736, 32'hc2ef9d5f},
  {32'h44f9adcc, 32'h42a8fc89, 32'h43c24365},
  {32'hc4bde6d7, 32'h43006566, 32'hc3842d9e},
  {32'h434df895, 32'hc4ba49b7, 32'h448a3a43},
  {32'hc4e412d2, 32'h43eec758, 32'hc32379d8},
  {32'h438274e8, 32'hc4058ab1, 32'h447bd675},
  {32'hc4eeefd6, 32'h41fbfd2a, 32'hc408844c},
  {32'hc28dc362, 32'h43f1a398, 32'h4582157f},
  {32'hc3324390, 32'hc3eba574, 32'hc4c9333a},
  {32'h446abad1, 32'hc497ee45, 32'h44acc021},
  {32'hc5048eb9, 32'h441ffe67, 32'hc470be63},
  {32'h44bfac0a, 32'h42f8fb24, 32'h43602b51},
  {32'hc50199ed, 32'h436f1e1b, 32'hc455ea78},
  {32'h45100557, 32'hc34f23e6, 32'hc336cd48},
  {32'hc3faf9ba, 32'h43effe88, 32'hc44e5d7a},
  {32'h4489284e, 32'h4405e36e, 32'h44c11e87},
  {32'hc545b953, 32'hc3cdbb86, 32'hc429c67e},
  {32'hc5036a2a, 32'h434442f9, 32'h426b07b5},
  {32'hc44d22fc, 32'h44829fea, 32'hc4899d7b},
  {32'hc223ba40, 32'hc4d5acfb, 32'h44c30e54},
  {32'hc3736b08, 32'hc45505c0, 32'hc29cfcb7},
  {32'h43de9590, 32'h437a2933, 32'hc4cfb178},
  {32'h4406e602, 32'hc46acbd4, 32'h44c312a5},
  {32'h4127c1d8, 32'hc319262c, 32'hc52000cb},
  {32'hc2b25d08, 32'hc4a79f82, 32'h42bb4cb0},
  {32'hc488bb30, 32'h441cb738, 32'hc466425e},
  {32'h44224039, 32'hc4597ec4, 32'h4490ffc7},
  {32'h4344b454, 32'h40c2e533, 32'h44c6d505},
  {32'hc49e66ca, 32'h449d3396, 32'hc4905068},
  {32'h422b3634, 32'h42f147e9, 32'h44118b92},
  {32'h44a0c274, 32'hc3f5539a, 32'h43e3ea5e},
  {32'hc402bfb9, 32'h444f5d2f, 32'hc4ae69b2},
  {32'h430de36e, 32'hc4fa2db9, 32'hc01b7f30},
  {32'hc4cb223a, 32'hbe82f890, 32'hc244d8c1},
  {32'h42b56016, 32'hc444cfb9, 32'h44a6ed18},
  {32'h4374da40, 32'h4517a95b, 32'hc16c1a50},
  {32'h44f47aa0, 32'hc424c0e3, 32'h441c5d69},
  {32'hc586854c, 32'h43ec91b6, 32'hc30eb449},
  {32'h4531b430, 32'h439a4494, 32'h43fe759b},
  {32'h44ba858a, 32'h4473b381, 32'hc3bc2a32},
  {32'h44a68d43, 32'hc42022c8, 32'h43f3a317},
  {32'hc49e8535, 32'h44e85595, 32'hc2900b38},
  {32'hc407da99, 32'hc3a58fa6, 32'h43877f36},
  {32'hc5594352, 32'h42cc2166, 32'hc3ba6c4d},
  {32'h43d61e69, 32'hc49d65db, 32'h443f3c10},
  {32'h444ed587, 32'hc2084058, 32'h43da857f},
  {32'hc43498b6, 32'hc494e729, 32'hc51b6a5b},
  {32'hc4af83f4, 32'hc45e5983, 32'h443a02b9},
  {32'hc4ddf91a, 32'hc364e5be, 32'h42dd4554},
  {32'hc3143f5a, 32'hc310b2d2, 32'hc535d421},
  {32'h4397c9b8, 32'hc2e2c28b, 32'h43c9ce97},
  {32'hc2f7be0a, 32'h41e72ea7, 32'hc4c35cde},
  {32'h43973589, 32'hc1f235a0, 32'h45444fc9},
  {32'hc29709c2, 32'h44866e94, 32'h43445b61},
  {32'h44d76a45, 32'hc3fa40f7, 32'h430718a0},
  {32'hc52cf2fd, 32'h438ea0a1, 32'h4480f3ea},
  {32'h411e4eee, 32'h43b94a2e, 32'hc5243a7a},
  {32'h449b2948, 32'h421e946b, 32'hc3d87098},
  {32'hc38dafde, 32'hc49ce00a, 32'hbf893404},
  {32'hc238c149, 32'h44c59141, 32'hc39184f7},
  {32'hc4856a3a, 32'hc1d35327, 32'h44e35140},
  {32'h446bc9f9, 32'h44115028, 32'hc2d71a30},
  {32'hc43454d2, 32'hc30b972e, 32'h441f0983},
  {32'h454c1ede, 32'hc3165854, 32'hc1d6dae2},
  {32'hc588b9ae, 32'hc288bcca, 32'hc402419a},
  {32'h4409850a, 32'h43b386b5, 32'hc2870ce6},
  {32'hc5556454, 32'h43834970, 32'h4200e3e8},
  {32'h45238d65, 32'h43924c09, 32'h4270d587},
  {32'h44e2eac0, 32'hc29d5493, 32'h4355d96f},
  {32'h44da47e2, 32'h4445ae87, 32'hc383232d},
  {32'hc4fca702, 32'hc41b905c, 32'h43937ebd},
  {32'hc4958f05, 32'h44374609, 32'hc41f43a3},
  {32'h438b702d, 32'hc3c17dfe, 32'h42f2bc32},
  {32'hc487ebda, 32'hc45d8905, 32'hc3c360b8},
  {32'h43a1b8a0, 32'hc40bc871, 32'h44a9063e},
  {32'h44710eac, 32'hc1d85a56, 32'h4307b279},
  {32'h44029934, 32'h451351f9, 32'h43a0d09d},
  {32'hc369d42a, 32'hc385aa05, 32'hc485a020},
  {32'h44be5afa, 32'hc349ba12, 32'h42e1e6d0},
  {32'hc50abd97, 32'h41b436b9, 32'hc41e1700},
  {32'hc41c6fc1, 32'h444eee44, 32'h44f94755},
  {32'h43bb7944, 32'h446f4a8a, 32'hc40caf54},
  {32'hc3446106, 32'h451c678c, 32'h435390ff},
  {32'h43c21dca, 32'hc3839652, 32'hc49724a5},
  {32'hc4d36b60, 32'hc2a14630, 32'h43178fea},
  {32'h4361b49e, 32'hc4ff3a64, 32'hc42e5ea8},
  {32'h4527fd57, 32'h43ab6add, 32'hc367f159},
  {32'hc4b96d2d, 32'hc28db903, 32'h432eb085},
  {32'hc46410b4, 32'h44383e72, 32'h453c9f8e},
  {32'hc3315c78, 32'h4213183d, 32'hc4e2e7ef},
  {32'h45506aba, 32'hc3b5a797, 32'h43c1e385},
  {32'hc484ce0c, 32'hc5189197, 32'hc4435898},
  {32'h440144d2, 32'h44e800cd, 32'hc2c487d6},
  {32'h4491bce1, 32'hc34bc010, 32'h3f8eb540},
  {32'h44a3cb20, 32'h449e311f, 32'h4438c47d},
  {32'hc3f8c578, 32'hc55fb56e, 32'h423dca19},
  {32'h450373a0, 32'h43b4d515, 32'h4319b424},
  {32'hc4a15948, 32'h43b68f3b, 32'h43a3835d},
  {32'h4508199d, 32'hc3b4f70c, 32'h41294f8c},
  {32'h44f88caf, 32'hc3226652, 32'h40c84bbd},
  {32'hc50fdae9, 32'hc36002b0, 32'h43e37b6f},
  {32'hc1f551e5, 32'hc4b560b5, 32'h419acbaf},
  {32'hc462a714, 32'h445ef900, 32'h438de350},
  {32'hc3d5b2d0, 32'hc3d63dfe, 32'hc4a63527},
  {32'h450f3761, 32'h4315c6cf, 32'h43c2e7ec},
  {32'h452d76c7, 32'hc1beed36, 32'hc40fdfe0},
  {32'hc4b58a38, 32'hc40a88f3, 32'h448be01e},
  {32'hc4f93c79, 32'hc3c73fa2, 32'h42a7fd5d},
  {32'h41d31e40, 32'h450e60a0, 32'h43d097bb},
  {32'h44f57ab1, 32'h43b06569, 32'h4360c781},
  {32'hc3b2d54c, 32'hc40d188d, 32'h442b0b78},
  {32'hc3883489, 32'hc317c05c, 32'hc2ddf08e},
  {32'hc3fcc538, 32'hc2fd9561, 32'h43a79274},
  {32'h437aa84c, 32'hc38ffca1, 32'h4221b3ea},
  {32'h43af294f, 32'h4417c6f8, 32'h451142c5},
  {32'hc3654d24, 32'hc461eae5, 32'hc4f99b54},
  {32'hc52222bd, 32'hc2edae29, 32'hc3c389a1},
  {32'h4403838e, 32'hc52eade0, 32'hc4191c9c},
  {32'hc42804aa, 32'h45173f37, 32'h43fbb85c},
  {32'h43c6acf7, 32'hc4f99e8b, 32'h42a92ed4},
  {32'hc3232044, 32'h44f06aa9, 32'hc300835c},
  {32'h42e6b168, 32'hc4f21682, 32'h40d50c58},
  {32'hc2b51708, 32'h449f4d47, 32'h42b8f1ee},
  {32'h456706e1, 32'h42e4fdc1, 32'h43cb94f4},
  {32'hc4650ece, 32'h41be9317, 32'hc223a3f4},
  {32'h4586d53f, 32'h423e58f6, 32'hc31e0853},
  {32'h442f9153, 32'hc3f5b05e, 32'hc3b86577},
  {32'hc4e562d0, 32'h41c61b14, 32'hc3e97bfa},
  {32'h449c321e, 32'hc34e3cff, 32'h4460042b},
  {32'hc3536148, 32'h44c45410, 32'hc40f7a3a},
  {32'h455e72da, 32'hc319c4cf, 32'h43da8a79},
  {32'hc4b11d19, 32'h4454e8ca, 32'h422c5390},
  {32'h45351dfa, 32'h43e7c786, 32'h42598436},
  {32'hc3b84a28, 32'h4500539e, 32'h4322e2ca},
  {32'h45316b05, 32'hc451bd7b, 32'h43b9db00},
  {32'hc3a8b6b0, 32'hc3bbf00e, 32'h42538cb1},
  {32'h442296f7, 32'h43d68b83, 32'hc4599886},
  {32'hc3e8dacc, 32'h441ab7de, 32'h41b6122c},
  {32'h443bc22d, 32'hc46da6cc, 32'hc460d405},
  {32'hc430efdf, 32'h43910c67, 32'h447d3e04},
  {32'h421ec1d0, 32'hc45633f4, 32'hc4e1e404},
  {32'hc48ad1f9, 32'hc36c50d6, 32'h4345988e},
  {32'h43a33882, 32'hc4d4eac7, 32'hc3c577ea},
  {32'hc3be8988, 32'h43cefe80, 32'h45349101},
  {32'hc4ad18af, 32'hc34fd429, 32'hc3e1bf40},
  {32'hc3b5dca8, 32'h443ff902, 32'h444cbff0},
  {32'h4307288a, 32'hc45d56e1, 32'hc43f6a63},
  {32'hc378366b, 32'h449d6b4c, 32'h443ff979},
  {32'h413309e4, 32'hc5256488, 32'hc3145bea},
  {32'hc361a378, 32'h42ce3e67, 32'h45369f17},
  {32'hc251c0f2, 32'hc4892b4f, 32'hc3d45807},
  {32'hc533da36, 32'h44103b5d, 32'h43769cba},
  {32'h44477f94, 32'hc4868613, 32'hc48e537d},
  {32'h42e4f280, 32'hc3d77820, 32'hc52d222f},
  {32'hc536a256, 32'h429cf142, 32'h41a2d6bd},
  {32'h445ff203, 32'h43fc9995, 32'hc2802de7},
  {32'hc483c7be, 32'hc4af3cc3, 32'hc2cc38e2},
  {32'hc2a31a48, 32'h450bf9fa, 32'h4332ba08},
  {32'hc4481781, 32'hc474ec5b, 32'hc3ff8a8e},
  {32'h44ae9949, 32'h445afe2d, 32'hc3a045b6},
  {32'hc453ddfe, 32'hc40875e1, 32'h440c40e9},
  {32'hc4d9d55f, 32'hc2b936d4, 32'h42b38d63},
  {32'hc38724ce, 32'hc4aa1690, 32'hc497264e},
  {32'h435808dc, 32'h40d0a6ac, 32'hc500f15d},
  {32'h43b40e37, 32'hc3bb29eb, 32'h442e5d66},
  {32'hc36a662f, 32'h44bed867, 32'h44454da3},
  {32'hc44a4698, 32'hc4c86b8e, 32'hc4c33cde},
  {32'h43cc5275, 32'h43a521d0, 32'hc22b7f4c},
  {32'hc324d53b, 32'hc44e5f89, 32'hc4b6c6a9},
  {32'h43edac9a, 32'h4497ba16, 32'h4463ceb4},
  {32'hc45e00f6, 32'hc4365dfc, 32'hc21f1f70},
  {32'h442ea7f0, 32'h42e34dfa, 32'h4486fac5},
  {32'hc5524eda, 32'h43da05cb, 32'hc34b43b5},
  {32'hc49d006f, 32'h43402542, 32'h4347d992},
  {32'hc4cf0ae7, 32'hc39de932, 32'hc4669153},
  {32'h409d5000, 32'h4419c5ee, 32'h44adf7ae},
  {32'hc413525d, 32'hc49cda2d, 32'hc3c397c1},
  {32'h4388ed2b, 32'h44d538c8, 32'h4367896f},
  {32'h41d39c08, 32'hc4258154, 32'hc5303fce},
  {32'h448cefca, 32'h4429e892, 32'hc3bff843},
  {32'h44a6dbd7, 32'hc1daa434, 32'hc3cce61e},
  {32'hc484af03, 32'hc42bf611, 32'hc44be668},
  {32'h448cbfc1, 32'h448c3bd2, 32'h42b8df2b},
  {32'h44c640b4, 32'h425f0ad1, 32'h43431392},
  {32'h4427a124, 32'h44f2fe1c, 32'hc2945334},
  {32'hc4c0316b, 32'hc4a00117, 32'h431d5ff0},
  {32'h45423eae, 32'hc40433f3, 32'hc42ba800},
  {32'hc55019b7, 32'h432aa279, 32'hc3c9ea93},
  {32'h4521a0fa, 32'h44795b54, 32'h444623a6},
  {32'hc3df4118, 32'hc414e929, 32'h44062a57},
  {32'h42fbec14, 32'h4517f81e, 32'h41dc99cb},
  {32'hc38fba53, 32'hc4b1e3d9, 32'h4434c8b5},
  {32'h4524924c, 32'hc2b32fb7, 32'h4255b3a2},
  {32'h4392511b, 32'hc37fa586, 32'h4530c60c},
  {32'h44f71dd9, 32'h43b5096e, 32'hc20ab883},
  {32'hc3b4ee64, 32'hc2d631c8, 32'h433f04f9},
  {32'h4419b3aa, 32'h3f251e50, 32'hc4922c77},
  {32'hc425a0a6, 32'h430e7f6b, 32'h449a3e74},
  {32'hc4cd18bc, 32'h42597bbc, 32'hc39c316a},
  {32'hc4b62d8b, 32'hc413773a, 32'hc3ad878e},
  {32'h442afb35, 32'h452d1dd6, 32'h4378ac20},
  {32'hc466c4f9, 32'h421c37b6, 32'h4311793d},
  {32'h444ec846, 32'h43bc0fae, 32'hc503dc38},
  {32'hc5256aa1, 32'hc427e843, 32'h430f722a},
  {32'h4484e9ee, 32'hc3605075, 32'hc416f38f},
  {32'hc52f6250, 32'h439f38ca, 32'h444ed616},
  {32'h44b8f58c, 32'h43511898, 32'hc4d0278a},
  {32'h44712888, 32'hc4343e44, 32'hc438d291},
  {32'hc4dcc6aa, 32'h4472fe04, 32'h42ad08c8},
  {32'h449dcc86, 32'hc2f3e876, 32'h43f2cbd0},
  {32'hc49cf8ce, 32'h448a56bd, 32'hc3d8ae15},
  {32'h44557e6d, 32'hc4ff8deb, 32'hc2f573be},
  {32'hc3303dfd, 32'h430b3f09, 32'h42d19497},
  {32'h44ab33b7, 32'h43b0cb97, 32'h430a6e41},
  {32'hc543ddf2, 32'hc321ba55, 32'hc0bf2479},
  {32'hc4a5b802, 32'hc2257f8c, 32'h4383963e},
  {32'h43a7aefa, 32'h451b4766, 32'h43d8f15d},
  {32'h426c688c, 32'hc4323ecb, 32'h44403d68},
  {32'hc52fa382, 32'h421e53ce, 32'hc3c020fc},
  {32'h43a07dfb, 32'hc3b0c76b, 32'h45283dac},
  {32'hc37b8664, 32'h4441b862, 32'hc44a7aa9},
  {32'hc36092f8, 32'hc3cb2d6e, 32'hc216ffc0},
  {32'hc437b47c, 32'hc39e6bbe, 32'hc4e36fc7},
  {32'h447541eb, 32'hc3c3640b, 32'h43d8c58d},
  {32'h449a0329, 32'hc29e82ea, 32'hc385b990},
  {32'hc3946d9a, 32'hc4bc8839, 32'h44bc86e5},
  {32'hc53834fa, 32'h439b1f43, 32'hc3c9d544},
  {32'hc3ad2c7a, 32'hc45688ef, 32'h43b5509c},
  {32'hc44615a1, 32'h450c59e9, 32'h437afc73},
  {32'h4501e9eb, 32'h4386801c, 32'h44106dd1},
  {32'hc47f7db8, 32'h43fac7eb, 32'hc43ea361},
  {32'h453a3092, 32'h436cd4c4, 32'h43fbfe1d},
  {32'hc403cf1d, 32'hc344bb38, 32'hc5289f02},
  {32'h44b0bf6d, 32'hc3a521c6, 32'h42fe737a},
  {32'h435d708a, 32'hc481e37e, 32'hc4833ab3},
  {32'h42aec41a, 32'hc44c1765, 32'h44a46151},
  {32'hc37acb0b, 32'hc3cfb2c8, 32'hc3e8285c},
  {32'hc4b736ec, 32'hc2a4e788, 32'h4337384b},
  {32'h440ea076, 32'h429823f6, 32'h4502b223},
  {32'hc3c11116, 32'h44c56a65, 32'hc3b49472},
  {32'hc21bb2c0, 32'hc3aea4de, 32'h44a42892},
  {32'hc372072f, 32'h442b154a, 32'hc43edd87},
  {32'h4465b55f, 32'hc402211b, 32'h42e66338},
  {32'h448af493, 32'hc4e634f4, 32'h44e33e99},
  {32'hc50cffc8, 32'hc330f29a, 32'hc442a72b},
  {32'hc327016c, 32'h440a85e6, 32'h43bea407},
  {32'hc3cb64d7, 32'hc459e434, 32'h4393fd08},
  {32'hc445afe8, 32'h44005201, 32'hc4b6528f},
  {32'h45090ad0, 32'h4409656b, 32'h43ce07ef},
  {32'hc4af79a7, 32'hc33fe4e1, 32'hc3179926},
  {32'h4492da1c, 32'hc2f9f198, 32'h44a658ae},
  {32'hc328906c, 32'h43225180, 32'hc4f8712b},
  {32'hc413c144, 32'h42c05b54, 32'hc3068a0d},
  {32'hc58bdd96, 32'h43615353, 32'h433cfefe},
  {32'h4450a20e, 32'hc29d2810, 32'h44817a83},
  {32'h44e66e37, 32'h4406c813, 32'h42eb792a},
  {32'h44945d9a, 32'hc5035382, 32'h44133c9a},
  {32'hc4b77d16, 32'h441b8945, 32'hc399a582},
  {32'h45185ba1, 32'h43f22cd4, 32'h43ddb6b1},
  {32'hc31231be, 32'h45745de2, 32'hc35612e2},
  {32'h44260cfc, 32'hc4bb5704, 32'h439de26d},
  {32'hc48586e3, 32'hc30f5a38, 32'hc3935e84},
  {32'hc3b5eb77, 32'hc3834aca, 32'hc52901d0},
  {32'hc3c7a20a, 32'hc13bfb58, 32'h44904875},
  {32'hc3db26c1, 32'hc4dec36c, 32'h4419d00e},
  {32'hc3456b79, 32'h452b9b60, 32'h424d8f55},
  {32'hc41d11a8, 32'h43632e9a, 32'h4503e534},
  {32'h4421337a, 32'h4260e000, 32'hc5264954},
  {32'h43bb068f, 32'hc43233ec, 32'h451a048e},
  {32'hc44a2940, 32'h445cbc2d, 32'hc3b26655},
  {32'hc2a817c2, 32'hc43b4013, 32'hc46c8c82},
  {32'hc4d861ec, 32'h43c8b637, 32'h44580d10},
  {32'hc24688e0, 32'h4276844c, 32'hc515cdb8},
  {32'h436adb40, 32'h444dbb98, 32'hc367a08b},
  {32'hc37763af, 32'hc49893c6, 32'hc313e407},
  {32'h448b8fcc, 32'h439ec1d8, 32'hc2d7c77c},
  {32'hc403fca3, 32'hc4c28bf3, 32'h433c5011},
  {32'h43a67577, 32'h44de22b0, 32'hc4a15f97},
  {32'h4485d12e, 32'hc2d6b5f4, 32'h4372da08},
  {32'h4525affa, 32'h424dcc9e, 32'h4373e75b},
  {32'hc4cbf99c, 32'h43e04e6d, 32'hc3bc316c},
  {32'h45119bca, 32'hc38619e6, 32'h440891b4},
  {32'hc55ea8ea, 32'hc3b7d53d, 32'h42d4a410},
  {32'h4436a557, 32'h4500517d, 32'hc3a5c165},
  {32'h430d5db1, 32'hc434ae14, 32'h439636b2},
  {32'h444ec24d, 32'h44d2181e, 32'hc39087ff},
  {32'hc5160a2a, 32'hc42b3093, 32'hc2359d37},
  {32'hc3e37dce, 32'h4464f7f4, 32'hc32b7008},
  {32'hc43a50a8, 32'h44a12a3d, 32'h4389d83c},
  {32'h441c9c14, 32'h4459f83b, 32'hc4df38b5},
  {32'h4380343b, 32'hc34381fa, 32'h44daaa75},
  {32'h447fee4a, 32'hc40e62ba, 32'h41aa8c1b},
  {32'h4427c0cc, 32'h44f45537, 32'h42d6c704},
  {32'hc3959dd8, 32'hc32c7a30, 32'hc5004afc},
  {32'h431baab4, 32'h44c7f923, 32'h4396d78e},
  {32'hc538c0b5, 32'hc395fb50, 32'hc30f9c3c},
  {32'h41d44e60, 32'h43f81b46, 32'h45543a7f},
  {32'h4361aac4, 32'hc2588f7a, 32'hc455b0a1},
  {32'hc4398d04, 32'hc4f3348b, 32'h4503d4b9},
  {32'hc46c5f3f, 32'h421adfd2, 32'hc39a25ac},
  {32'h4210c7c4, 32'hc369da9b, 32'h440a16e1},
  {32'hc2de5fa7, 32'h40e7902e, 32'hc51f26e2},
  {32'h44420b2a, 32'h4470967c, 32'h43756a8c},
  {32'hc482999e, 32'h437b1746, 32'hc035c9a0},
  {32'h429aee31, 32'h43f67fa6, 32'h4565fb95},
  {32'hc3d274bc, 32'hc4998131, 32'hc4703e43},
  {32'h43826507, 32'h448a10ef, 32'h436d7f31},
  {32'hc3ee82be, 32'hc4bca987, 32'hc22f0470},
  {32'h454ab998, 32'h44653e02, 32'hc38de01c},
  {32'hc5153a15, 32'hc21bac9b, 32'hc1b79ac2},
  {32'h4480a73d, 32'h446a78d6, 32'h444d320b},
  {32'hc4584b99, 32'hc475b07d, 32'h43702199},
  {32'h448af522, 32'hc33234e8, 32'h44130d48},
  {32'hc58fe356, 32'hc39a7524, 32'hc3a7f063},
  {32'h43d80e58, 32'hc2cdf478, 32'h437746eb},
  {32'h417e03f8, 32'hc3d337fc, 32'hc4227beb},
  {32'hc469acbf, 32'h44d022e9, 32'h429671b9},
  {32'hc1f0e7f8, 32'h448abc02, 32'hc4076b8e},
  {32'hc46e215b, 32'h45060ae0, 32'h430bd1f0},
  {32'h44459a94, 32'hc44d42c0, 32'hc373c754},
  {32'h450e7074, 32'h419f5334, 32'hc38ad75b},
  {32'h43dcba66, 32'hc45d0d37, 32'hc5004df0},
  {32'hc317d8ec, 32'h443d3fed, 32'h451c9a61},
  {32'h4315b71c, 32'hc4336e8f, 32'hc2adae0b},
  {32'h43f99170, 32'hc4b1e10a, 32'h4516a78e},
  {32'h43b47c8c, 32'hc48c6115, 32'hc42691f8},
  {32'h43c5b705, 32'h44c2124c, 32'hc3983582},
  {32'h4407e424, 32'hc35bb7ae, 32'hc49adbed},
  {32'hc535d1a1, 32'hc30ad3e4, 32'h43f05dee},
  {32'hc37e5c4e, 32'hc48d5c6a, 32'hc3017696},
  {32'hc48a69aa, 32'h430cce85, 32'h446f9aab},
  {32'h445304b6, 32'hc49d79af, 32'hc48184ad},
  {32'hc4a0d049, 32'hc393dd01, 32'h43628866},
  {32'h45342621, 32'hc485571d, 32'h43ec5d0c},
  {32'hc2b423d0, 32'h447bc6ca, 32'h4416af6c},
  {32'h455a8cc0, 32'h43904885, 32'hc419d295},
  {32'hc448c710, 32'h452f6525, 32'hc3ab1c5a},
  {32'h4514a3ef, 32'h43a1ad14, 32'hc383ec52},
  {32'hc48f96ea, 32'hc34a80fc, 32'h439d0f52},
  {32'h45113721, 32'h435177d8, 32'h441a2a92},
  {32'hc53bca7a, 32'hc3ac279a, 32'hc35a2b96},
  {32'h4577322f, 32'h438849cd, 32'h43c73856},
  {32'h44dc61ef, 32'hc385f31e, 32'hc38a80aa},
  {32'hc3d6dee0, 32'hc3a2eb2d, 32'hc4437df9},
  {32'h44d0a06c, 32'hc39c463f, 32'h445f2322},
  {32'hc532253a, 32'hc45968d8, 32'hc3c1f62a},
  {32'h4334c350, 32'hc4a58da6, 32'h42b88992},
  {32'hc4974400, 32'h4477972b, 32'h43781cee},
  {32'h44642126, 32'hc49b6354, 32'hc070b0ff},
  {32'hc5549f86, 32'h432308af, 32'hc203849e},
  {32'h45114327, 32'hc49040b8, 32'h429328f8},
  {32'h438b9ec2, 32'hc390e378, 32'hc48364ea},
  {32'h4488e518, 32'hc3aad182, 32'h44945645},
  {32'hc4849bbf, 32'h43a45f9a, 32'hc453413f},
  {32'h4535f9a4, 32'hc16cc7c0, 32'h41992cbb},
  {32'hc5142ee6, 32'hc27e2ad3, 32'h43d52690},
  {32'h42a7ac80, 32'h42b404e2, 32'hc50a5372},
  {32'hc3d2a572, 32'h4274ce3d, 32'h4474579a},
  {32'hc3429f9a, 32'h43181850, 32'hc53a5724},
  {32'hc438f80e, 32'h43e72a58, 32'h451ab795},
  {32'h45111080, 32'hc26ffb50, 32'h43ef76cf},
  {32'hc54750cc, 32'h443c6a6b, 32'h43c7b72e},
  {32'h4538522a, 32'hc3baac90, 32'hc4345cd8},
  {32'h4412c226, 32'h4337eae7, 32'h44eb25e0},
  {32'h44131d13, 32'hc3979f16, 32'hc26e181a},
  {32'hc29cef14, 32'h4483f038, 32'h446cca41},
  {32'h450477cf, 32'hc155c9be, 32'h42b09c33},
  {32'hc3023ba8, 32'h44f4cadb, 32'h4482cebb},
  {32'h44a1f2ba, 32'hc48ac5b4, 32'hc478b9a0},
  {32'h4552438a, 32'h43571552, 32'hc389d036},
  {32'hc4e64967, 32'hc2f58088, 32'h4427b38a},
  {32'h453a9f53, 32'hc1aa4b0d, 32'h44540141},
  {32'hc379fdd0, 32'hc4fd8a72, 32'hc38f6672},
  {32'h43e3448c, 32'h44c06a6e, 32'h431b7417},
  {32'hc5180fab, 32'h420cf18f, 32'h429c39d3},
  {32'h44ee25f8, 32'h44aa38a7, 32'hc3572620},
  {32'hc49d7fca, 32'hc4bab90b, 32'hc459b330},
  {32'h435dba70, 32'h4353db40, 32'h44190b32},
  {32'hc4c57464, 32'hc2867cc4, 32'h43701672},
  {32'h44c34528, 32'hc3c9e9ce, 32'hc2ef1090},
  {32'h440a2f46, 32'hc31c0b3e, 32'hc31ccd95},
  {32'h437bec86, 32'h44b0a7c5, 32'h444af08b},
  {32'hc44b5bd8, 32'hc4497b0c, 32'h41e5e632},
  {32'hc1b63f60, 32'h440d5b20, 32'h43a5eb67},
  {32'hc2eff300, 32'hc40de2c2, 32'hc45221d2},
  {32'h43cef45d, 32'h42fecc1f, 32'h451daef8},
  {32'h4506a120, 32'h42cc3cb8, 32'hc3f915b0},
  {32'hc3c1e9e2, 32'h41339983, 32'h42986a82},
  {32'hc55bd9d0, 32'hc20fdc7f, 32'hc2c7f76a},
  {32'h454e29f5, 32'h43439c5b, 32'hc432f380},
  {32'h43a45483, 32'hc5638156, 32'h4285a391},
  {32'h4418a3f2, 32'hc3c83ae0, 32'h44d17a4e},
  {32'h4473713c, 32'hc43ebbeb, 32'hc2669138},
  {32'h453211d9, 32'hc29ea7c3, 32'h4364852b},
  {32'hc47fb04e, 32'hc33a736a, 32'hc535798b},
  {32'hc335ad76, 32'h43501d39, 32'hc3e3bf08},
  {32'h435bff34, 32'h44b9f3d0, 32'h43bf573f},
  {32'hc4afebc4, 32'hc40fe9c5, 32'hc35abae8},
  {32'hc3326ce8, 32'h451e2f3f, 32'h4431b367},
  {32'h44ead56b, 32'hc3d9ab4f, 32'h4351f936},
  {32'h44092061, 32'h451e25f4, 32'hc1fa5f1c},
  {32'hc2af3150, 32'hc49059a8, 32'hc3b7b0bb},
  {32'h44ea9fc2, 32'h439f72f1, 32'hc39ca6d5},
  {32'hc44dd36a, 32'hc4eefa8e, 32'hc4c56e31},
  {32'h44fc4c1a, 32'hc3e72f44, 32'hc3038ba8},
  {32'h4493f252, 32'hc3204631, 32'hc3b9d1fc},
  {32'h43b0908e, 32'h446697dc, 32'hc35fcd7c},
  {32'hc36c37f8, 32'hc3f99c8b, 32'h42d51f6f},
  {32'h434cf922, 32'h44c7aa65, 32'h439ded55},
  {32'hc3bb4014, 32'hc3fa21dc, 32'h44cad2b5},
  {32'h4448b6ca, 32'h445e6a4e, 32'hc4a06ff8},
  {32'h443fffed, 32'hc36fdbd1, 32'h44577c66},
  {32'h43b700a3, 32'hc3f1213a, 32'hc4c2910c},
  {32'hc253f67c, 32'h43fc1898, 32'h448f84af},
  {32'h434263b2, 32'h44877922, 32'hc2385fce},
  {32'h434b8322, 32'hc4507c16, 32'h44491c2a},
  {32'hc39fd8f0, 32'h44b8dbff, 32'hc2a7be43},
  {32'hc3cca414, 32'hc2c123bf, 32'h435845c3},
  {32'h441d35f4, 32'h44094cd7, 32'hc4112292},
  {32'h41af2c78, 32'hc4ae7e59, 32'h4450d42b},
  {32'h45664364, 32'h4465cbbb, 32'h3fe32120},
  {32'hc4a6619a, 32'h4422d50f, 32'h44c2ec8f},
  {32'h44aa902f, 32'h41963ba3, 32'hc4d45d6e},
  {32'hc27eb545, 32'hc49cf41e, 32'hc44d9178},
  {32'hc3f48dbc, 32'h455dd239, 32'h430fa6c3},
  {32'hc3ef796b, 32'hc363ab44, 32'h4412d1e9},
  {32'hc38b77e0, 32'h453a8cc5, 32'hc37be824},
  {32'h44cf76a8, 32'hc48028d8, 32'hc2adb2c9},
  {32'h44a4e9b5, 32'h4436e163, 32'hc3b36f9b},
  {32'h451bfd87, 32'hc3c3aa10, 32'hc22837c8},
  {32'hc4962741, 32'h430a3181, 32'h43079c72},
  {32'h4547a727, 32'h42c315f5, 32'h43807a92},
  {32'hc4b7d2d0, 32'h4062f4fa, 32'h41e01f3c},
  {32'h430bb35e, 32'h44906d70, 32'hc4cf95fa},
  {32'hc3aa377c, 32'h4413b306, 32'hc4957c8f},
  {32'h451d9004, 32'hc2fffca9, 32'h44208d9c},
  {32'hc410e4b0, 32'h40b90d41, 32'hc4d99180},
  {32'hc200d9d0, 32'hc4e3bdcb, 32'hc3667a3d},
  {32'hc4e029fe, 32'h431b9997, 32'h430f9fa1},
  {32'h4296c430, 32'h4391b202, 32'h453989c7},
  {32'h44b53b52, 32'h442611c6, 32'h43b3dd99},
  {32'h44ae8268, 32'hc423ebc2, 32'h4491540f},
  {32'hc3e33040, 32'h44b58b3e, 32'hc4ba86a4},
  {32'h444c9fd4, 32'hc38359ef, 32'hc20e8951},
  {32'hc391b994, 32'h4454ed8c, 32'hc4136247},
  {32'h44c78408, 32'h4302ed72, 32'h4400f636},
  {32'h44127c36, 32'h44c6c995, 32'h43d3d5ac},
  {32'h43a24528, 32'h444d293c, 32'h45428838},
  {32'hc56fc41b, 32'h4384e9e0, 32'hc41bf470},
  {32'h453fa745, 32'h435f4e97, 32'hc3c5678f},
  {32'hc38ea50f, 32'h448d81d8, 32'hc4c08683},
  {32'h42406b3c, 32'hc4c56985, 32'h451c9aa3},
  {32'hc46c242c, 32'hc4117ca2, 32'hc380dfb0},
  {32'hc41e1a72, 32'h447a58ae, 32'h42d945a0},
  {32'h43d1d350, 32'hc4cb923d, 32'h441ab123},
  {32'hc4cc666a, 32'hc30ecd7e, 32'hc478bb26},
  {32'h43f110ad, 32'h434ccd37, 32'h44b9a8c6},
  {32'hc496c83e, 32'h44523509, 32'h41a04d07},
  {32'h42d6c2e8, 32'hc4dd36d2, 32'h4461c800},
  {32'h443a1f5a, 32'h438e6b0e, 32'h449aee4b},
  {32'hc18cc044, 32'h435a3087, 32'hc533cd78},
  {32'hc2873543, 32'h4483c3ca, 32'h43661a22},
  {32'h4497095c, 32'hc3852fbc, 32'h442ba148},
  {32'hc3ab85bf, 32'h44809cc0, 32'hc2542d6b},
  {32'hc3a1957c, 32'hc4ea20c3, 32'hc34c3ec4},
  {32'hc52ed65d, 32'hc2d7b702, 32'h417b653a},
  {32'h4517e12e, 32'hc30dde14, 32'h4416960e},
  {32'hc43ce83e, 32'hc2b9924a, 32'hc424f6c3},
  {32'hc48af86c, 32'h42f82a11, 32'hc31020dc},
  {32'hc3c90af8, 32'hc3dc4447, 32'h44037b83},
  {32'h44d40dd4, 32'hc3848b05, 32'hc3b9d465},
  {32'hc34f6f13, 32'h44a9a6d5, 32'h43e281ef},
  {32'h454512b2, 32'h436047fb, 32'h438edd0d},
  {32'hc3b6bb58, 32'h451a1b24, 32'hc33e676e},
  {32'hc444fff0, 32'hc3df436d, 32'h441158fc},
  {32'hc4e2bd1b, 32'h446e0d18, 32'hc41efdd5},
  {32'hc33a696c, 32'hc578d39e, 32'h43665e21},
  {32'h447bee04, 32'hc373e57c, 32'h43b555c2},
  {32'hc36ee089, 32'hc4f7e7f0, 32'hc4c66ec1},
  {32'h44944a23, 32'hc313deec, 32'h445bd728},
  {32'hc22adf40, 32'hc49174ad, 32'h442d2ee6},
  {32'h441a56d6, 32'h44ac2ee4, 32'h430a0306},
  {32'hc5077320, 32'hc38a1170, 32'h40efb20f},
  {32'h439542c6, 32'h447ae033, 32'hc44e6185},
  {32'hc4a4b04c, 32'hc3bfe9d0, 32'h43ad5e93},
  {32'hc31493c5, 32'h44911d6b, 32'h43b445f1},
  {32'h4452ff1a, 32'hc4054d27, 32'hc455146c},
  {32'hc47d1ad1, 32'hc3907b55, 32'h44df22e9},
  {32'h450970aa, 32'hc30f06a2, 32'hc452e019},
  {32'h449439e2, 32'h447230ca, 32'hc3145ade},
  {32'hc3e9a737, 32'hc380a072, 32'h43a3e2bc},
  {32'hc34ae3e0, 32'h4313b233, 32'hc423b56f},
  {32'hc5072549, 32'hc371cfae, 32'h43d96c33},
  {32'h4503c806, 32'hc28e69c1, 32'h42da3a16},
  {32'hc4783a84, 32'hc38d8ea3, 32'h43e9392a},
  {32'h451ddaca, 32'hc425ae82, 32'h42b8a164},
  {32'hc491c474, 32'h40e24b0c, 32'h43b94e18},
  {32'h4564dec2, 32'hc39fa356, 32'h44028b54},
  {32'hc549b176, 32'hc341242f, 32'h42e34262},
  {32'h453060b9, 32'h43f04d2a, 32'h434a1f63},
  {32'hc49d7ae6, 32'hc381f8b5, 32'h4309ab36},
  {32'h4530121a, 32'h44472f83, 32'h43318f8a},
  {32'hc4307d9c, 32'hc5184b44, 32'h43e868c9},
  {32'h4409417e, 32'h42e46210, 32'hc334407e},
  {32'h42631d9c, 32'hc2098c0c, 32'h44378ab8},
  {32'h43239670, 32'hc2c24717, 32'hc4b32211},
  {32'hc387c44c, 32'hc495da41, 32'h4509f978},
  {32'hc3596c5a, 32'hc34a4e49, 32'hc4f79471},
  {32'h441d803f, 32'hc33ad006, 32'h45435196},
  {32'hc2ce7e21, 32'h420e8cb9, 32'hc3fec952},
  {32'hc2839558, 32'h44989a62, 32'h44155fbf},
  {32'hc42b524f, 32'hc32d9b8d, 32'hc53770be},
  {32'h43ffde22, 32'h440b8c5f, 32'h447382ca},
  {32'hc4d567af, 32'h43c8c0a8, 32'h43c63ee1},
  {32'h4401c5a4, 32'hc38077b8, 32'h43c60566},
  {32'hc3dbbea8, 32'h4393babc, 32'hc4a68e13},
  {32'h450d033c, 32'hc1ab9f2e, 32'h42d80d5c},
  {32'h43188a58, 32'hc52b8141, 32'hc3ffe8aa},
  {32'h45118eb2, 32'hc2772a4c, 32'hc2588f4c},
  {32'h44376a71, 32'hc40d6036, 32'hc44313e1},
  {32'h42a01039, 32'h43c4130e, 32'h454039eb},
  {32'hc401984f, 32'hc4aab1df, 32'hc4a7326a},
  {32'h450e5080, 32'hc329de7c, 32'h43aaff99},
  {32'hc4da45bd, 32'hc4cdca49, 32'h436acc0e},
  {32'h4527824e, 32'h447f771c, 32'h42d643d4},
  {32'h44db0885, 32'hc38a6862, 32'hc3f4371a},
  {32'h4469bec7, 32'h45040110, 32'h442be761},
  {32'hc4191ba0, 32'hc55db43d, 32'hc3b6d057},
  {32'h45384d7c, 32'h443082f0, 32'h4246c01c},
  {32'hc52f3dfc, 32'h43ec0d69, 32'hc4815428},
  {32'h44aebacc, 32'hbfa0ae18, 32'hc2c75a22},
  {32'hc3d39d2b, 32'h44832a2c, 32'hc51e0075},
  {32'hc3cd2456, 32'h44ff4d47, 32'h41da6514},
  {32'hc2d86ec5, 32'h41fc6b77, 32'hc4603d11},
  {32'hc1749f80, 32'h444598ad, 32'h44a6de07},
  {32'h431a3eb3, 32'hc4aec46c, 32'hc49d4539},
  {32'h444908ce, 32'h4292a86b, 32'hc37b9385},
  {32'h448dd39e, 32'hc387cc52, 32'hc4bc7b51},
  {32'hc4f511c4, 32'h440b0ee2, 32'h43dfa78a},
  {32'h447df8e4, 32'hc46ea9af, 32'hc342ae58},
  {32'hc43225d6, 32'h4500614e, 32'hc3b0deba},
  {32'hc401795c, 32'h448ababe, 32'hc4fa68a2},
  {32'h43e6eb56, 32'h42a8905c, 32'h44a05e36},
  {32'h43ba00d8, 32'hc213b8bf, 32'hc4d9ceb5},
  {32'hc3826862, 32'h4363d662, 32'h44e65e03},
  {32'h4370ae74, 32'h4277083d, 32'hc4479b91},
  {32'hc395b4e6, 32'h43a969e7, 32'h4430700c},
  {32'h4534fe96, 32'h43ccd73d, 32'hc33d8783},
  {32'h44b7f3dc, 32'hc31bc8d3, 32'h43b555d5},
  {32'h44162e7b, 32'hc54be29d, 32'h43d05dd2},
  {32'hc4aefae6, 32'h44f1debc, 32'hc2da5554},
  {32'h4406f136, 32'hc408d459, 32'hc31f2e26},
  {32'hc36d63ad, 32'h45575c11, 32'h405d4d94},
  {32'h441b52cc, 32'hc4c203e7, 32'h4346f748},
  {32'hc23b63c0, 32'h4435510c, 32'h4301ccb7},
  {32'h4529f108, 32'h431e9206, 32'h4425cb13},
  {32'hc2e7eec0, 32'h42f9f738, 32'hc353b250},
  {32'h45278ebe, 32'hc2a6015b, 32'hc373601c},
  {32'hc4bf8888, 32'hc379647a, 32'hc200abcf},
  {32'hc542d95e, 32'h4383b338, 32'h4322ebe7},
  {32'h423f5180, 32'h43c5c2db, 32'h443f9c7c},
  {32'h43338f02, 32'h44f25f01, 32'h42df8b56},
  {32'h442c7373, 32'hc48038b8, 32'h439145ba},
  {32'hc4bcdc33, 32'h448edeb7, 32'hc202631f},
  {32'hc3955451, 32'hc4905273, 32'hc1fe0602},
  {32'hc39d9c14, 32'h4502666f, 32'hc406adcb},
  {32'h453dd665, 32'hc34b05d8, 32'h43c2a65a},
  {32'h43f5cbb7, 32'hc3b290e3, 32'hc441abc0},
  {32'h43c0d0e0, 32'h437077d0, 32'hc42c4703},
  {32'hc43a1351, 32'hc4077b91, 32'h44258e3c},
  {32'h44943d9e, 32'hc3004e67, 32'hc3a224de},
  {32'hc2f07d33, 32'h436314fd, 32'h44a4fac4},
  {32'hc224f8d0, 32'hc4538ff8, 32'hc47b845d},
  {32'hc379f61c, 32'h43ea7626, 32'h44089312},
  {32'h438f2e55, 32'hc421f1ca, 32'hc4734300},
  {32'hc416586e, 32'h44c087fd, 32'hc35d563f},
  {32'h41817f70, 32'hc3a10a1f, 32'hc3bee387},
  {32'hc5256e60, 32'h4441073b, 32'h444ed156},
  {32'h43b8c6ee, 32'h43d4fa61, 32'hc497d84a},
  {32'h44046da9, 32'h43097c00, 32'h44de5d6c},
  {32'h4381a67c, 32'hc42b87fc, 32'hc4f27529},
  {32'hc44adb8c, 32'h43758fc1, 32'h44339937},
  {32'h42cfe6e8, 32'hc2b31e82, 32'hc4f8b146},
  {32'hc2dd7a10, 32'h4496085c, 32'h4437ce32},
  {32'h441242e8, 32'hc3ac7394, 32'hc4f0f6d8},
  {32'h4526369c, 32'hc3441836, 32'hc434914e},
  {32'hc4703500, 32'h41769a1e, 32'h44a2ec42},
  {32'h44cc02b6, 32'h4395b82d, 32'h43dcb9ed},
  {32'hc4ad434f, 32'hc4413ea2, 32'hc31faf49},
  {32'h4409b837, 32'h44bba369, 32'hc16847bc},
  {32'h44654aa1, 32'hc3b7caac, 32'hc2b54459},
  {32'h448e7e90, 32'h44b764f6, 32'h4351724b},
  {32'hc4718a6c, 32'hc4ecbec1, 32'hc24d30ce},
  {32'h448d13fc, 32'hc3d0cccc, 32'h440bbc16},
  {32'hc440519b, 32'hc384dd5c, 32'hc2a6143e},
  {32'h44b29c55, 32'hc3353f23, 32'hc4027a9f},
  {32'hc5389006, 32'h429c737a, 32'hc2888f9a},
  {32'h451f298a, 32'h438e417a, 32'h4431a9cb},
  {32'hc27c2250, 32'hc457f63e, 32'hc4b67e7e},
  {32'h442f9a8d, 32'h43224758, 32'h436eef17},
  {32'hc4e83857, 32'hc3996879, 32'hc46dfcf9},
  {32'h44c5f828, 32'h43af122e, 32'h43fd64af},
  {32'h43cba93b, 32'hc20bbc28, 32'hc467d0a5},
  {32'h44b9fe59, 32'h44687304, 32'h44c3149d},
  {32'hc58993e6, 32'h433eba52, 32'hc3d37b4b},
  {32'hc3f7a62c, 32'h438eb3d9, 32'hc319c69c},
  {32'h42bc0e8c, 32'hc51f705f, 32'hc437c87a},
  {32'h44db6a06, 32'hc1a68cbc, 32'h422a4a56},
  {32'hc4a26646, 32'hc3e1fe0b, 32'h42e0dd15},
  {32'h4347e1a0, 32'h44d7b9ff, 32'h44395bf5},
  {32'h42dc30f8, 32'hc5107720, 32'hc43470ed},
  {32'h43d8c0a2, 32'h44c4ee07, 32'hc3f56b79},
  {32'hc4a65ced, 32'hc388305c, 32'h439c6e5e},
  {32'h40262240, 32'hc55bf726, 32'hc38f7acb},
  {32'h4446cec6, 32'h44db3cbc, 32'hc38918a1},
  {32'hc215562c, 32'hc3a28054, 32'h41a35016},
  {32'h445c6a40, 32'h44b2161e, 32'hc3b37d70},
  {32'h428d14e0, 32'hc53f91a0, 32'hbdab0910},
  {32'h44bd5196, 32'h43adeae5, 32'h42d4fcd7},
  {32'hc4517bc6, 32'hc3b43ff1, 32'hc34dd290},
  {32'h45778865, 32'h427e820b, 32'h43fa0a73},
  {32'hc233d5a0, 32'hc418c8c1, 32'h438c381a},
  {32'h45018dc9, 32'h436177c4, 32'hbe14da12},
  {32'hc30dd470, 32'hc4375944, 32'h441efc07},
  {32'h435f3519, 32'h445f4282, 32'h4208c682},
  {32'hc398d8d8, 32'hc51a2a3b, 32'hc174bbbe},
  {32'h433ed323, 32'h453c2c55, 32'hc4060eab},
  {32'hc46af9f0, 32'hc32a43f7, 32'h431a087d},
  {32'h4511928f, 32'h431f2e29, 32'hc3f5f84e},
  {32'hc2b2ccb2, 32'h43bebf76, 32'h45486bab},
  {32'h44247934, 32'hc38c03cc, 32'hc2768290},
  {32'hc500c7b5, 32'hc3f32102, 32'hc39c21f5},
  {32'h4423d323, 32'h44808d7d, 32'hc516e74f},
  {32'hc553d759, 32'h43989d70, 32'hc2e7e77e},
  {32'h449eec72, 32'h439cad1f, 32'hc3a66ddb},
  {32'h4295ecf4, 32'hc231f920, 32'h453b7643},
  {32'hc455a24f, 32'h43347477, 32'h428db23a},
  {32'hc3cdea40, 32'h4393716e, 32'h44a5c5a6},
  {32'h43b5e170, 32'hc2c02a5c, 32'hc53a22db},
  {32'h4281be74, 32'hc52a38d3, 32'hc29d1c26},
  {32'hc38125dc, 32'h453e0a3d, 32'h43924da4},
  {32'h4521c205, 32'h43bcf1b5, 32'h439f3477},
  {32'hc40c738e, 32'h44f4e848, 32'h44399e40},
  {32'h43eb02b6, 32'hc52eb96a, 32'h43eeba5c},
  {32'hc3220b98, 32'h42bcfa66, 32'hc315f215},
  {32'h45500da6, 32'h434506c6, 32'hc27a1cdf},
  {32'hc41382dc, 32'h44acd782, 32'h448d6cf3},
  {32'h455d3f14, 32'h42c53d1c, 32'h438c409c},
  {32'hc4bf902f, 32'h44553e15, 32'hc3aaeb24},
  {32'hc328af5a, 32'hc5025b2f, 32'hc360195d},
  {32'hc4a130f4, 32'h42bb6325, 32'hc419eed1},
  {32'h4527a2f2, 32'hc330c6d4, 32'h43eb5e99},
  {32'hc4209e9a, 32'h43fe5af0, 32'h431e6d4a},
  {32'hc4b999b4, 32'h43ebc43e, 32'h444c2b11},
  {32'hc3b20e14, 32'h4221240a, 32'hc4815e94},
  {32'h4542fd6c, 32'hc412c7a3, 32'hc2ad6be8},
  {32'hc4b0eb42, 32'hc36753e6, 32'hc3d53dea},
  {32'h441c39f9, 32'hc419f741, 32'h44db0fbf},
  {32'h433b8d5b, 32'h4545353e, 32'h4233ad52},
  {32'h43931210, 32'hc49f696a, 32'h44b3b097},
  {32'h430d62f5, 32'h441b89ee, 32'hc4a11ce7},
  {32'h43f475ee, 32'h43b363fe, 32'h448f60ca},
  {32'hc41bf67d, 32'h43d85dd9, 32'h42a6e5e2},
  {32'hc4080b77, 32'h4307bf7d, 32'h44888e7e},
  {32'hc54cdcfa, 32'hc2c43fe9, 32'hc4732a84},
  {32'h44e61268, 32'hc3d5aacc, 32'hc38fc7b7},
  {32'h440431cc, 32'h44b8ad4f, 32'hc539f5ce},
  {32'h4451f8a2, 32'h43a5e62a, 32'h44741500},
  {32'hc33aa01a, 32'h449547f1, 32'hc3b3609e},
  {32'hc48bd3e6, 32'h42a921dc, 32'h42cd8cab},
  {32'h444657f8, 32'hc32586d2, 32'h45029240},
  {32'hc541cbc3, 32'h43462cf7, 32'hc192b5ad},
  {32'h4406dc6c, 32'h42a0f6d4, 32'h448bf3d0},
  {32'hc287d2de, 32'h44f6933c, 32'hc3b69a41},
  {32'h450713c5, 32'hc3c1d96a, 32'h441f5772},
  {32'h44045a7e, 32'h437b8d02, 32'h44a3a727},
  {32'hc4b05118, 32'hc4bfd54b, 32'hc48a8807},
  {32'hc41ba404, 32'h4331ccbe, 32'h44ce96f5},
  {32'h44070d07, 32'hc480c037, 32'h42e3a9a4},
  {32'hc53967e0, 32'hc3b65abc, 32'h42ddeb0f},
  {32'h444bb34c, 32'hc3a93ebf, 32'h43e9e343},
  {32'hc4a94471, 32'h40a55170, 32'h4197cb30},
  {32'h44726e4c, 32'hc4197a2b, 32'hc3de475a},
  {32'h42cb4636, 32'h41b6770a, 32'hc5136458},
  {32'h4499324c, 32'hc3fc604e, 32'h4383d30f},
  {32'hc4f0a156, 32'hc468ae28, 32'hc3c1ef0c},
  {32'hc45b49d0, 32'h42b77000, 32'hc3a88a8a},
  {32'h44d15328, 32'h439ee72e, 32'h42472bde},
  {32'h4428b0ba, 32'hc545c0cb, 32'h439db3fe},
  {32'h43e50f18, 32'h457a2c98, 32'hc374f101},
  {32'h454dfe76, 32'h43bfd7c8, 32'h43671060},
  {32'hc4fae68e, 32'h44aeb3f8, 32'hc29f9215},
  {32'h4556603e, 32'hc4429034, 32'hc3c2ffbf},
  {32'hc31102a0, 32'hc4b51db4, 32'h43fefd4a},
  {32'h4502e5bc, 32'h430f1e4c, 32'hc3a7c84f},
  {32'hc3f6c1ee, 32'h449bb015, 32'h449f81d3},
  {32'hc316c670, 32'hc40e858c, 32'h44cd56c7},
  {32'h43f039a8, 32'h4461c28f, 32'hc314fe37},
  {32'h444ee4bf, 32'hc3327ed0, 32'h421605e4},
  {32'h446e9886, 32'h44eeaec2, 32'h42c3d22f},
  {32'hc387bc70, 32'hc4c17be1, 32'h4435c011},
  {32'hc4745718, 32'hc102638a, 32'hc33af500},
  {32'h43c43961, 32'hc3ac30bd, 32'hc49e50a8},
  {32'hc2dbf300, 32'hc42fccb8, 32'h44eadb58},
  {32'h43e6eda8, 32'h44afd6e7, 32'hc4c79558},
  {32'h44ffd858, 32'h440b4ff6, 32'hc335a351},
  {32'hc50fe502, 32'h42a5ed44, 32'h42e2e730},
  {32'h4425ef01, 32'hc12a8db4, 32'hc44954cf},
  {32'hc48d9c1f, 32'hc3db159b, 32'h441c5c4a},
  {32'h439c57de, 32'h43a8d007, 32'hc5091630},
  {32'h44407962, 32'hc364b3c0, 32'h433fbe96},
  {32'h44988b72, 32'h429795c0, 32'hc394122f},
  {32'hc59d0bd6, 32'h429be1db, 32'h42d346fc},
  {32'hc427e5c8, 32'h43e55d1e, 32'hc3c1e921},
  {32'hc4d7fb3a, 32'hc47edff6, 32'h41d121b7},
  {32'h43bbcfde, 32'h450ebe11, 32'hc30ce3bf},
  {32'hc4dde655, 32'hc3b29082, 32'hc28a080a},
  {32'h44a20591, 32'h4494b235, 32'hc35ed91b},
  {32'hc2b06b83, 32'hc51b040a, 32'hc3af2a58},
  {32'h42223480, 32'h4487c104, 32'hc371ab2c},
  {32'hc35c4a74, 32'h440114ff, 32'hc3bcce9e},
  {32'hc4fe9b11, 32'hc219dcc4, 32'hc3874ccb},
  {32'h418e2d24, 32'hc40835fd, 32'h44bcf653},
  {32'h44c455c8, 32'hc3f4897c, 32'hc389433c},
  {32'h44c5aaf6, 32'h448a71e5, 32'h4331232c},
  {32'h4353b250, 32'hc46b8e98, 32'hc48479d6},
  {32'hc4686868, 32'h438c3ade, 32'h43400b71},
  {32'hc3e51c80, 32'hc3cbea86, 32'hc51759d1},
  {32'h43c2a878, 32'h44b07578, 32'h44a72120},
  {32'hc43402f6, 32'hc3732534, 32'h41d2724d},
  {32'h40b3ed68, 32'hc50cce43, 32'h44ec50cc},
  {32'hc47e891b, 32'hc2683c50, 32'hc46db244},
  {32'h4449170d, 32'h4448febc, 32'h436a3ff6},
  {32'hc4a51b7e, 32'hc2f95875, 32'hc4859472},
  {32'h43a7a57e, 32'h43b6ba28, 32'h452a8dfd},
  {32'h44266b6a, 32'hc47bb6a0, 32'hc204e6fe},
  {32'h44ca1f23, 32'h42e35857, 32'h4484b27d},
  {32'hc52a5d98, 32'hc3035e8c, 32'hc4851dbf},
  {32'h45275576, 32'hc3e371e0, 32'h43a147ee},
  {32'hc54ee5c0, 32'h432369ac, 32'hc2cf4818},
  {32'h44d8fabd, 32'h448f5613, 32'hc31e0237},
  {32'h42fca2b3, 32'h428ed7fb, 32'h413584db},
  {32'h452205dd, 32'h438e97d7, 32'h43fb25c5},
  {32'hc265b614, 32'hc54008ae, 32'hc3ddde6d},
  {32'hc3d78f72, 32'hc293eced, 32'hc192b145},
  {32'hc56ca98e, 32'hc35361ff, 32'hc35696f2},
  {32'h449ef268, 32'hc37e846c, 32'h42d93d19},
  {32'h43892eeb, 32'hc4c88777, 32'hc471c83e},
  {32'hc29e78c8, 32'h4527996e, 32'h44308ebb},
  {32'hc4528293, 32'h44973123, 32'hc39736ac},
  {32'hc4c9d1a1, 32'h447c9a46, 32'h4426e4e4},
  {32'h43994d18, 32'hc4f2fd61, 32'hc452896e},
  {32'hc394cef8, 32'h44c249b4, 32'h4402106c},
  {32'h44735488, 32'h42b2d00a, 32'hc46448e1},
  {32'hc2f2c5f0, 32'h44bf2e9d, 32'h44e8dfe6},
  {32'h44620b6e, 32'h4389de11, 32'h4238bbce},
  {32'hc3a066f4, 32'h3f9a2950, 32'h439f0d88},
  {32'h428872ca, 32'hc4d37fb5, 32'hc47cf44b},
  {32'hc5000c19, 32'h4374ee8e, 32'hc2f23f1e},
  {32'hc2c0d420, 32'h41ced2ca, 32'hc41903c3},
  {32'hc422c303, 32'h43857ce3, 32'h44a98f4a},
  {32'hc4d25a61, 32'hc20ff2a9, 32'hc2d3b692},
  {32'hc44f108e, 32'h43c64d01, 32'h44a925a4},
  {32'h450b6cae, 32'h4327b0cd, 32'hc4235ce1},
  {32'hc3db7ab2, 32'h437c69da, 32'h448c277c},
  {32'h44f6d8b4, 32'hc48c78c8, 32'h41072f63},
  {32'hc4bf1e89, 32'h4495376c, 32'h40e7a202},
  {32'h43f31adc, 32'h4372b3a3, 32'h442b5e7d},
  {32'h42edd8ca, 32'h455edf20, 32'hc31846fd},
  {32'h45634899, 32'hc2ac474b, 32'hc37cdebd},
  {32'hc428425e, 32'h4414127a, 32'h4345eab0},
  {32'h455af8bb, 32'hc2084056, 32'h43b01592},
  {32'hc5346386, 32'h43ae2c5b, 32'hc33722fd},
  {32'hc479ebdc, 32'hc3a8a1d2, 32'hc1785bd9},
  {32'h450b06a4, 32'h43878f74, 32'h423ff4fd},
  {32'hc4d9958b, 32'hc25f03d7, 32'hc309663a},
  {32'h42f2d630, 32'hc3918ada, 32'h44ef9822},
  {32'hc4acab5c, 32'hc3b910e2, 32'hc31eda3e},
  {32'h44aa8379, 32'hc4bd8835, 32'hc18a1d30},
  {32'hc4365f14, 32'h44668671, 32'hc30a2f0c},
  {32'hc4237a3d, 32'hc494bb2b, 32'h436fb793},
  {32'hc4842d1c, 32'h43faa90a, 32'hc334a2c4},
  {32'h4481afdb, 32'hc4c8443c, 32'h42930b90},
  {32'hc416cbf8, 32'h41a3dc67, 32'hc3c95ab3},
  {32'h4385f12a, 32'hc4332a8c, 32'h4520d68c},
  {32'hc3dc69f6, 32'h437d2f0a, 32'hc38e66ca},
  {32'h43e26eca, 32'hc4ae41ed, 32'h4218ef75},
  {32'hc4a35ef0, 32'h42ea891e, 32'hc2dc07d9},
  {32'h450391b6, 32'h4307f6b9, 32'hc3d55120},
  {32'h420122ac, 32'h42b65544, 32'h44a9119e},
  {32'hc39d325c, 32'hc4771503, 32'hc398bdcf},
  {32'hc48cd423, 32'h43d2e0c5, 32'h44ce3db7},
  {32'h44eda7ce, 32'h4251dcdd, 32'hc400229c},
  {32'hc56f733b, 32'hc319df19, 32'h41c314da},
  {32'h451ab175, 32'hc2280d2d, 32'hc436c2d8},
  {32'hc3869d16, 32'h427aa3e3, 32'h4429853b},
  {32'hc2b568be, 32'hc4d20ca4, 32'hc4a67bc3},
  {32'hc3f3da29, 32'h41c0c48a, 32'h44d17266},
  {32'h427a2820, 32'h4229604b, 32'hc4483c55},
  {32'hc3d742a3, 32'h444fccc4, 32'h44595ee6},
  {32'h4443e8d2, 32'hc3ac218b, 32'hc5453e1b},
  {32'h43a40844, 32'h4137d42a, 32'hc4b51fd9},
  {32'hc466be98, 32'hc3f9dd2d, 32'h452fcb7b},
  {32'h454b1497, 32'h435a22d6, 32'h43d0e99d},
  {32'h417a03d8, 32'hc5514814, 32'h41b096a6},
  {32'h443f0e38, 32'h444cfd0f, 32'hc26f2323},
  {32'hc5223a0a, 32'hc38900fc, 32'h43cc7166},
  {32'hc4034f6d, 32'h439bb768, 32'hc4191cde},
  {32'hc5080948, 32'hc466482e, 32'hc4602f76},
  {32'h4521f0f3, 32'h439c881d, 32'h43ba0f35},
  {32'hc51f49ea, 32'hc3edde65, 32'h42b9ad3d},
  {32'hc2551992, 32'hc1d09b7c, 32'h43803a68},
  {32'hc4e38d08, 32'hc352d4de, 32'h43d709b2},
  {32'h43787757, 32'hc363d945, 32'h44fa9520},
  {32'hc3b50cd4, 32'hc5595b8e, 32'hc39d8141},
  {32'h41bcca05, 32'h44d4c0c6, 32'h40d7d3e7},
  {32'hc3c9dd43, 32'hc507ba01, 32'hc271217a},
  {32'h442c4718, 32'h4386ec2e, 32'h44cd77a4},
  {32'hc36e8eec, 32'hc4e2d0fd, 32'hc25c91f3},
  {32'h429f8042, 32'h43fcd3b3, 32'h4314a173},
  {32'hc481ef64, 32'hc468fd2f, 32'hc4a9ceb2},
  {32'h443a371b, 32'h43b92da1, 32'hc377bc07},
  {32'hc2f26e16, 32'hc4e53e84, 32'hc3a5decf},
  {32'hc4184561, 32'h45492da0, 32'hc3894886},
  {32'h44c61ce0, 32'h41cdce7f, 32'hc3e06d02},
  {32'h4400ee97, 32'h44d99eea, 32'h439f509a},
  {32'hc4c22f50, 32'hc38b0fcd, 32'hc4e7f50f},
  {32'h43bd0ab7, 32'h450c6a59, 32'hc3e968d1},
  {32'h450c417e, 32'hc40238cb, 32'hc2610d98},
  {32'hc4aaa334, 32'hc42532e1, 32'hc2a05c15},
  {32'h43f74ee0, 32'h44a86194, 32'h44347fdd},
  {32'hc3c702e8, 32'hc3a5f259, 32'h43b358ce},
  {32'hc1d717de, 32'h458a1347, 32'h426909ea},
  {32'hc41aa4c5, 32'hc35f5f84, 32'h3d39e38e},
  {32'h442c6b58, 32'hc3091d6e, 32'h4335556c},
  {32'hc5107fe2, 32'hc4436ae6, 32'hc30b9236},
  {32'h44529148, 32'hc33f0f40, 32'h4318b82e},
  {32'hc362fe80, 32'hc41e91e5, 32'h43c00b94},
  {32'h44e56c78, 32'h43831549, 32'h43810207},
  {32'hc3d464a5, 32'hc444aead, 32'h442f1332},
  {32'h3e920c40, 32'hc3a0379e, 32'hc473a91e},
  {32'hc22a798c, 32'hc5292238, 32'h433b9cee},
  {32'h43cff9c8, 32'h44720f2f, 32'h4400f65c},
  {32'hc45da5d0, 32'hc37f20ba, 32'h42afb86d},
  {32'h437f2028, 32'h44851e37, 32'h4455e0ae},
  {32'hc4bc164a, 32'h42c67588, 32'h4412e980},
  {32'h44b5a3a9, 32'h4263cb32, 32'hc46f0f4e},
  {32'hc50ae2a8, 32'hc425d625, 32'h430bd0d5},
  {32'h429d2c0f, 32'h4525cb3d, 32'hc39b35d3},
  {32'hc33504cd, 32'hc452a209, 32'h441b2151},
  {32'h450d8133, 32'hc3d43a2c, 32'hc3904842},
  {32'hc49a8b81, 32'hc40c7ee8, 32'h43c6a0d6},
  {32'h45195b07, 32'h4376847c, 32'h420a428c},
  {32'hc48237b6, 32'h431d5c54, 32'h44d8d94b},
  {32'h43a8aa50, 32'hc3050920, 32'hc4d549e2},
  {32'hc3ec702d, 32'hc565265f, 32'h4254447c},
  {32'hc398a482, 32'h451f6a50, 32'h42804673},
  {32'h441bd034, 32'hc3d500f7, 32'h43ce1a75},
  {32'h42f8f840, 32'h4537618c, 32'h42e3c447},
  {32'h44b25f5b, 32'hc4940fde, 32'h43c60685},
  {32'h427736e8, 32'h44093ee0, 32'h43c21aaf},
  {32'h452d3cc2, 32'hc2f9edf8, 32'hc430be62},
  {32'hc41f0040, 32'hc420c3f0, 32'hc1e04ca5},
  {32'h44f3dd41, 32'h414c7b70, 32'h43fea978},
  {32'hc4d113a7, 32'h43e93dd4, 32'hc43137e4},
  {32'h4447535b, 32'hc4debe54, 32'hc3a02e21},
  {32'hc38cce4f, 32'h405ef95b, 32'h43023c70},
  {32'h439a450d, 32'hc302513a, 32'h44f73ff3},
  {32'hc42a6d12, 32'h43f42992, 32'hc300e6c3},
  {32'h4507808b, 32'h43435c0a, 32'h4286041c},
  {32'hc3eaab7c, 32'h442cc42f, 32'h4413e33b},
  {32'hbf3451a0, 32'h44268bd7, 32'h456cd7cb},
  {32'hc50b9a5a, 32'h41d5a11c, 32'h43ab0914},
  {32'h4392b91f, 32'hc43c20e1, 32'h444fde6c},
  {32'hc4c9a29f, 32'h44b129b1, 32'hc4139b80},
  {32'h4525fab2, 32'hc22e0ed6, 32'hc3a894c4},
  {32'h43696893, 32'h448a7563, 32'hc4739bec},
  {32'h44e4aac8, 32'hc464629a, 32'hc39c1a0b},
  {32'h43528506, 32'h4427979f, 32'hc3bf430b},
  {32'h44c2925a, 32'h431e6c05, 32'h445c24fb},
  {32'hc4463340, 32'hc3a4b73f, 32'hc386498e},
  {32'h455f5097, 32'h3e945550, 32'hc40c123e},
  {32'hc50156af, 32'hc2c48ac2, 32'hc3e066d5},
  {32'h437f2fb0, 32'hc3697004, 32'h445ebfe9},
  {32'hc48901eb, 32'hc3b0dfcf, 32'hc3a37d0d},
  {32'hc3ecf065, 32'h44aa21d7, 32'h42799b14},
  {32'h447d17a1, 32'hc3176a8d, 32'h44f32e84},
  {32'hc3c4148b, 32'h445b4b7e, 32'hc4565718},
  {32'hc242feff, 32'hc40e3bdf, 32'h4490ff51},
  {32'hc4dc652c, 32'h4363b4e9, 32'hc495219c},
  {32'h4208a140, 32'hc4fd040d, 32'h442155d0},
  {32'hc214cb6e, 32'h44d10a88, 32'h44d43205},
  {32'hc5087bef, 32'hc4523606, 32'h42a0d37f},
  {32'h432aca2e, 32'h43323b9f, 32'h4395a761},
  {32'h4499a86d, 32'hc3e0f952, 32'h44318475},
  {32'hc4fd5829, 32'h433dd618, 32'h42f76264},
  {32'h4387b842, 32'hc4d0c5d5, 32'h43a21b7b},
  {32'h432727db, 32'h44c5f799, 32'hc280b15a},
  {32'h44011459, 32'hc3288f75, 32'h448e4335},
  {32'h41df2260, 32'h43d0bea2, 32'h42ca3e39},
  {32'hc3870b02, 32'hc3eeafa0, 32'h431904d1},
  {32'hc4b28954, 32'h41b9c6f3, 32'hc36cd0b6},
  {32'hc32373b8, 32'hc40c2e14, 32'hc4017907},
  {32'h4505f99a, 32'h4393bd00, 32'hc3e23150},
  {32'h44e4baa9, 32'h42c15e4e, 32'h4303abf9},
  {32'hc3f7e166, 32'h44fb86cb, 32'h43522b86},
  {32'h447ddd7e, 32'h43a6c79b, 32'h43887fa2},
  {32'hc5509bee, 32'h43eaed59, 32'h43c39fd1},
  {32'h4327e0ee, 32'hc463c3e6, 32'hc41d2319},
  {32'h424fc213, 32'h43eac0e7, 32'h44666d4d},
  {32'h4447a5fd, 32'h44eefac8, 32'hc4584704},
  {32'hc37c6e74, 32'h446449ab, 32'h44f8c4f6},
  {32'hc39760a0, 32'hc2dd6de7, 32'h451bf41e},
  {32'h4506f3f3, 32'hc2db37d2, 32'h422c8486},
  {32'h4478adde, 32'hc39f3208, 32'h44107984},
  {32'hc3b8f801, 32'h4493ffde, 32'hc3f9d384},
  {32'hc42d6aba, 32'hc4371acf, 32'h448d1a0f},
  {32'hc34eeae8, 32'hc33041ec, 32'hc490854e},
  {32'hc2b87582, 32'hc4173fdd, 32'hc4895e81},
  {32'hc42491e6, 32'hc504dfaf, 32'h44b372bb},
  {32'h4421bf90, 32'h448d5a87, 32'hc43bd17b},
  {32'h442f6359, 32'h43a721ab, 32'hc4a4ba48},
  {32'hc49f5a34, 32'h41c80278, 32'h44131c08},
  {32'h43fe0504, 32'h44a6f730, 32'h42288896},
  {32'hc4539794, 32'hc381c038, 32'h44bad5d4},
  {32'h44bd0d1a, 32'hc3c21c4c, 32'hc3bb1600},
  {32'h4364f7b3, 32'hc3342bbc, 32'h44e0864a},
  {32'h44a0ddb6, 32'hc3cbe414, 32'h439ab9fe},
  {32'hc480187f, 32'hc2af64fe, 32'hc3f90061},
  {32'h430dd640, 32'hc2f17cea, 32'hc2f00673},
  {32'hc3ecf76d, 32'hc5506c84, 32'h42e1c770},
  {32'h4499fe12, 32'h4474b2f1, 32'hc1894388},
  {32'hc39c9d5d, 32'hc40c4354, 32'h437da94b},
  {32'h45529705, 32'h44162840, 32'hc30a53c0},
  {32'hc5833a73, 32'hc32764f2, 32'h4281c1c3},
  {32'h4528682d, 32'h432a0bd6, 32'h43db06ec},
  {32'hc3e1391c, 32'h43b9664c, 32'h432d22df},
  {32'hc3979d04, 32'h445d2f98, 32'hc4540d80},
  {32'h44bffc94, 32'hc38fa6a7, 32'h43af6616},
  {32'hc4a0a4a4, 32'h4375d145, 32'hc35cf24a},
  {32'hc3958710, 32'h440daf3b, 32'h44bdc03e},
  {32'hc42d554e, 32'hc4c0ed7c, 32'hc474c7ef},
  {32'h446e9424, 32'h43b6a1d9, 32'h43852a00},
  {32'hc4caecef, 32'h43ccfa95, 32'hc3c6c109},
  {32'h447adf88, 32'h44a78319, 32'h446aa5a0},
  {32'h442f3a64, 32'h43df2b6f, 32'hc42c3713},
  {32'hc2a8fd76, 32'h44eb1607, 32'h43bb32d8},
  {32'hc3a0e0b8, 32'hc4f66ff8, 32'hc3d243e9},
  {32'h44d1802f, 32'h42f20363, 32'h43b666c2},
  {32'hc3149026, 32'hc4525a9c, 32'hc4e53f4b},
  {32'hc3e24de4, 32'h441ee2a2, 32'h444efd26},
  {32'hc428893c, 32'hc2440d09, 32'hc411353f},
  {32'h445b385b, 32'h4383b61d, 32'h4527f850},
  {32'hc1944a20, 32'hc345a301, 32'hc52936b1},
  {32'h447ae786, 32'h43f928ac, 32'h4422c370},
  {32'hc468b06b, 32'hc51127e2, 32'h43a69e1c},
  {32'h43f49f30, 32'h45149bc8, 32'h4451c9fd},
  {32'hc506beee, 32'h4394a415, 32'h42914691},
  {32'h44917402, 32'h448e9ba1, 32'hc3d4d51f},
  {32'hc5080cf9, 32'hc3f6f45e, 32'h43398d96},
  {32'hc269954c, 32'h441bc2f1, 32'h4420e8f9},
  {32'hc5867165, 32'h42b790bd, 32'h43831674},
  {32'h429f2fb7, 32'h43c3d169, 32'h44106500},
  {32'h43aa4da4, 32'hc3a6c5fc, 32'hc4612ed1},
  {32'h42d8f50e, 32'h45168899, 32'h42b28c5d},
  {32'hc446f025, 32'hc4de19c5, 32'h43371521},
  {32'hc4d0a6ae, 32'h44593d29, 32'h41e350c5},
  {32'h43fbd1d6, 32'hc1aa917a, 32'hc4edd988},
  {32'hc420edee, 32'h4325c504, 32'h445e0d6a},
  {32'h4460e86c, 32'hc4de90c0, 32'hc4be184e},
  {32'hc51469ec, 32'h442d0bfd, 32'h43e88248},
  {32'h448eb92b, 32'h437f9141, 32'hc47fe081},
  {32'h43279174, 32'hc4339876, 32'h44bb4cdf},
  {32'h42594fd0, 32'hc4982c80, 32'hc424875f},
  {32'h43e8f01b, 32'h434393f2, 32'h43eac50a},
  {32'h43545f70, 32'h4313fff4, 32'hc518fa29},
  {32'h430de382, 32'h43b9681f, 32'h44150710},
  {32'hc41559a2, 32'hc46b8ada, 32'hc3c47aa5},
  {32'hc3daba13, 32'h446ae861, 32'h4543a2d3},
  {32'h43f9892c, 32'hc3f4713b, 32'hc4cab808},
  {32'h4474c507, 32'hc320f73e, 32'h43c1c9d1},
  {32'h44ebf897, 32'hc4a2c465, 32'hc2cfc2a3},
  {32'hc486e4dc, 32'h448f1ed5, 32'hc31452ee},
  {32'h45582389, 32'hc2afbfaa, 32'h42795891},
  {32'hc3468866, 32'h4466dc9d, 32'h42720f91},
  {32'hc399551a, 32'h434f5b33, 32'h434aa65f},
  {32'h445b4300, 32'h4422acd1, 32'hc28714c5},
  {32'h453e4936, 32'h439f2395, 32'h428abd9e},
  {32'hc537a6ab, 32'h44408964, 32'h44155a93},
  {32'h437dc75b, 32'h43942e45, 32'hc3e16907},
  {32'h45467e2f, 32'hc2f34ebc, 32'hc3b51c5e},
  {32'hc4fa401c, 32'hc295113b, 32'hc34fd3fb},
  {32'h455359ed, 32'hc2652d73, 32'h42cbbd20},
  {32'h44d2173b, 32'h4286aa4f, 32'h4202a8c4},
  {32'h43c2c674, 32'hc54e0fb8, 32'hc2a69778},
  {32'hc21ca1d2, 32'h44943b41, 32'hc408658a},
  {32'h42fcc190, 32'h40700700, 32'hc2938089},
  {32'hc43e4c70, 32'h4415010a, 32'hc276b0d8},
  {32'h453c9916, 32'hc361331f, 32'h44058af9},
  {32'hc5045b50, 32'h42c15602, 32'hc0f7afad},
  {32'h43e2102c, 32'h42d7f905, 32'hc3c78444},
  {32'hc4c940d4, 32'h40dfc2a0, 32'hc1ecfcda},
  {32'h45065bfa, 32'hc340c007, 32'hc273dca4},
  {32'hc2d92404, 32'h4485284e, 32'h448089f3},
  {32'hc31133d6, 32'hc336c04e, 32'hc4834d61},
  {32'h413b6680, 32'h449f989b, 32'h441bf848},
  {32'h44744fa6, 32'h43d9a44d, 32'hc419a31a},
  {32'hc37d0af4, 32'h44bf03ef, 32'h439043d9},
  {32'h431513eb, 32'hc2ed0f89, 32'hc3cb8cdb},
  {32'hc50acf27, 32'h445d5825, 32'h43c06818},
  {32'h44249b84, 32'hc4013807, 32'hc4b18f75},
  {32'hc3cadae7, 32'h448f1231, 32'h436b6cb0},
  {32'h45367e61, 32'hc42db335, 32'hc3a3fbe7},
  {32'hc501d6af, 32'hc2a7772d, 32'h44358c66},
  {32'hc2c57140, 32'hc427c930, 32'hc355212a},
  {32'hc3a5ebc8, 32'h4517784e, 32'h43f939c0},
  {32'h44ce1b6a, 32'hc32459b5, 32'hc4a685c5},
  {32'h43e94872, 32'hc36ddf67, 32'hc3108e18},
  {32'hc481448c, 32'h43af2852, 32'hc32156ee},
  {32'h44e0176c, 32'h429780da, 32'h4368f7ba},
  {32'hc5059aad, 32'hc4b20bff, 32'hc405de61},
  {32'h448480a0, 32'h44911eee, 32'h43bf3c4d},
  {32'hc4921c72, 32'hc263531b, 32'hc0ec6788},
  {32'h444eebbc, 32'h454baba3, 32'hc312788d},
  {32'hc4c2f81a, 32'hc4913f67, 32'hc3877634},
  {32'hc50c5f3a, 32'h42b09d8c, 32'h42d3fb88},
  {32'hc44f63c4, 32'h43b6c125, 32'h4487a54f},
  {32'h4489126c, 32'hc2d3bbf3, 32'hc411b5df},
  {32'hc50def1d, 32'hc3ac5ec1, 32'hc28fe6ba},
  {32'h438d4db3, 32'h432aa36c, 32'h45335106},
  {32'hc4a53b39, 32'hc436ad05, 32'hc499579a},
  {32'h42ba3626, 32'h437cf6bc, 32'h44a523de},
  {32'hc4d7964a, 32'hc4183791, 32'hc4491459},
  {32'h44a49aea, 32'h442c4789, 32'h442a0f4d},
  {32'h438bbdb6, 32'hc345719a, 32'hc4902d25},
  {32'h4445ec4a, 32'hc3afbae0, 32'h44948e11},
  {32'hc498af67, 32'h4490e41a, 32'hc49f00d4},
  {32'hc336808b, 32'h43969eac, 32'hc3934f82},
  {32'hc3abe958, 32'hc50887ba, 32'hc42d8498},
  {32'h439fcab4, 32'h451b07f3, 32'h43e50398},
  {32'h43993362, 32'hc485470b, 32'h42e22014},
  {32'h4357cc44, 32'h44a8970a, 32'h442eebed},
  {32'h43983232, 32'hc5478d06, 32'hc3431d4b},
  {32'h440ec0a4, 32'h44843b5d, 32'h435cf942},
  {32'h447ffd53, 32'h4346a41a, 32'hc404d7c3},
  {32'hc3bf7f54, 32'hc486ed3a, 32'hc4648991},
  {32'hc2deed70, 32'h43f2fad4, 32'h44932cbc},
  {32'h433b5c33, 32'hc3e44465, 32'hc31216fa},
  {32'h442f96b5, 32'h44e5ce48, 32'hc3f93ad7},
  {32'h4257e19a, 32'hc53fc0d8, 32'hc37db5e5},
  {32'hc3ab20fb, 32'hc363bf61, 32'hc29f09f0},
  {32'hc545dbec, 32'hc3c0b719, 32'hc3a57781},
  {32'h44488860, 32'h42e289d4, 32'h42b9eb2a},
  {32'h43973d3d, 32'hc30e3bec, 32'h44100823},
  {32'h4435ccc8, 32'h43321100, 32'h43f02068},
  {32'hc3b24084, 32'hc4d9dfdc, 32'hc37ce1f3},
  {32'hc3eba92f, 32'h41942936, 32'hc4d8fdb4},
  {32'hc3a4fad0, 32'hc41570a8, 32'h44435840},
  {32'h44ba863a, 32'h43b24884, 32'hc3985bea},
  {32'hc4dda016, 32'hc350ea8e, 32'hc39881b8},
  {32'h4498feb9, 32'h43297086, 32'hc401198d},
  {32'hc43ca542, 32'h440bf7d2, 32'h451dbdae},
  {32'hbff9ea00, 32'h4469a81d, 32'hc31e6340},
  {32'hc469046a, 32'hc482c761, 32'h43c740b4},
  {32'h45135033, 32'h4431d480, 32'hc3939e44},
  {32'hc3bc467d, 32'hc3225941, 32'h440e7669},
  {32'h43855f86, 32'h44f72e2f, 32'hc388942f},
  {32'hc4d5a4ff, 32'h434f3041, 32'h423c891b},
  {32'hc47e1167, 32'hc35d5046, 32'hc3585c60},
  {32'hc5319b84, 32'hc378b32a, 32'h43ad0388},
  {32'h447eb99e, 32'h41923bfd, 32'hc4fce4c3},
  {32'hc2c11800, 32'hc4f4126a, 32'h4396a228},
  {32'hc4ea5314, 32'h44822cb5, 32'h43383bb4},
  {32'h44cd669b, 32'hc30ea679, 32'h43be97ef},
  {32'hc443d764, 32'h43b7a6f2, 32'hc432cc4c},
  {32'h44fbb7e6, 32'hc3873bfc, 32'h436b759f},
  {32'hc3b7edf2, 32'h44b42ab1, 32'hc39bb4fd},
  {32'h4485597e, 32'h43c50b93, 32'hc480eb19},
  {32'hc4fe4520, 32'h44307a68, 32'h430f034e},
  {32'hc2779a0f, 32'hc23640ef, 32'h4339bfe2},
  {32'hc3824fc5, 32'h44c70601, 32'hc384bbef},
  {32'h450902fa, 32'hc3104e5a, 32'h4372c3bc},
  {32'h431dae84, 32'h44cd1fc0, 32'hc276b229},
  {32'h43d74af6, 32'hc3dee644, 32'h4369968e},
  {32'hc51e4aa2, 32'h440406db, 32'hc3717541},
  {32'h4505807c, 32'h43a49c2e, 32'h43542a8d},
  {32'hc3a1b3f8, 32'h431f50b5, 32'hc4b0e2c9},
  {32'h44b44d1d, 32'hc35a0fbc, 32'h4383c0a5},
  {32'hc2cb24ee, 32'hc43512cf, 32'hc4faf5a2},
  {32'h426303c0, 32'hc4d688c3, 32'h4478c891},
  {32'hc4c8f016, 32'h4500c0f3, 32'hc40256cb},
  {32'h4437e610, 32'hc469aeaf, 32'h44a84c17},
  {32'h4309f0c8, 32'h446a86e4, 32'hc458e18b},
  {32'h44b2b5fe, 32'hc49a53bc, 32'hc3288b96},
  {32'hc2dd68f7, 32'h4349a7da, 32'hc4e23c99},
  {32'h4568dd0a, 32'hc2fc3888, 32'h44087afd},
  {32'hc51e050b, 32'hc40e0df5, 32'hc448889a},
  {32'hc3d26566, 32'hc2ca722f, 32'h43aebeef},
  {32'hc227d98a, 32'hc50d4ac7, 32'hc4d6b70e},
  {32'hc3099e84, 32'hc4b9263c, 32'h4518fab7},
  {32'hc4eff1ce, 32'h439e3266, 32'hc3742de0},
  {32'h447016b4, 32'h4396d761, 32'hc2332838},
  {32'h44532e39, 32'hc47a0bcb, 32'h44b05b88},
  {32'hc2ed2742, 32'hc31d0ee9, 32'hc50c5a93},
  {32'h44d1f7a8, 32'hc394a794, 32'h4385b78c},
  {32'hc4571c1e, 32'h439dd49d, 32'hc52a5ea0},
  {32'h4505e027, 32'hc3b2f39d, 32'h43c7c683},
  {32'h43c25766, 32'h44815cc7, 32'h44844ed3},
  {32'hc439e286, 32'hc3a70aac, 32'hc438db4c},
  {32'h44c654ca, 32'hc303beb7, 32'h43620c91},
  {32'hc4924c60, 32'hc4066f1b, 32'h42e1955e},
  {32'hc43231f2, 32'h44be2aa5, 32'h4409bd8c},
  {32'h445b78a2, 32'hc3cefd41, 32'h4131c930},
  {32'h42737b30, 32'h4205f110, 32'hc26d99bd},
  {32'h43a7fbac, 32'hc4cf40b9, 32'h43c0fa29},
  {32'hc42034a4, 32'h44c30a7d, 32'hc21435fb},
  {32'hc496f6b2, 32'hc38499ca, 32'hc3459132},
  {32'hc44cf288, 32'h4098ce70, 32'hc40a218e},
  {32'h4580bfb6, 32'h42e966cb, 32'h43aa67fe},
  {32'hc4f06244, 32'h43540ae6, 32'h42a5d125},
  {32'h430a2b80, 32'hc3e1374a, 32'hc3d0f503},
  {32'hc4a40240, 32'h448e1991, 32'hc2a38cef},
  {32'h437c1086, 32'hc4ef9a22, 32'hc32aa9d8},
  {32'hc407016e, 32'h43285e4f, 32'hc335d2bd},
  {32'hc388ec50, 32'hc4934fbb, 32'h4403ef4d},
  {32'hc4b05ddd, 32'hc200db00, 32'hc37ccb00},
  {32'hc35a6a06, 32'h43cfb0d8, 32'hc50c37a6},
  {32'h43a96367, 32'hc46a5bee, 32'h44bdf2ed},
  {32'hc3fc4335, 32'h43b9d084, 32'h44db0c3d},
  {32'h44d4faae, 32'hc2f623d3, 32'hc36df345},
  {32'hc44fe215, 32'hc4938386, 32'h42f1853c},
  {32'hc2b50fbe, 32'h44f17419, 32'hc47073ef},
  {32'hc40a78cc, 32'hc50f3715, 32'h435c2226},
  {32'h43a3a180, 32'hc1373aed, 32'hc4f7ed54},
  {32'hc3e0d306, 32'h44650ea1, 32'h41eeca17},
  {32'h438a1fdf, 32'h448c4c5c, 32'h451b015a},
  {32'h43104e9d, 32'hc4a0488c, 32'hc4c2141b},
  {32'h43848a11, 32'h4407a939, 32'hc4923ed4},
  {32'hc369e9a0, 32'hc41c9b01, 32'h445d1a95},
  {32'hc248f638, 32'h4388ecff, 32'hc4090ac7},
  {32'hc44e72d8, 32'hc47b6950, 32'h440bc334},
  {32'h44320e68, 32'h43f678f2, 32'hc3d1fb02},
  {32'hc46bfa13, 32'hc35caf2e, 32'hc4601211},
  {32'h452ad0d4, 32'h42cbd958, 32'hc3cfc9cd},
  {32'hc4da1b14, 32'h43ecc5d3, 32'hc3d25f9e},
  {32'h444fc0be, 32'hc274a207, 32'h43c8622f},
  {32'hc38ec4eb, 32'hc43b173c, 32'hc1c74654},
  {32'h443dfcdb, 32'hc338a1a2, 32'hc2822dba},
  {32'h43a784b5, 32'hc283f015, 32'h4323d91e},
  {32'hc1ce7340, 32'h4558a2cf, 32'hc3278df4},
  {32'h4398adbe, 32'hc56d0f5a, 32'h4288b581},
  {32'h443afd62, 32'h44a44249, 32'hc327f770},
  {32'h43c01ca9, 32'h43b2a303, 32'h43ae5be8},
  {32'hc4654ca4, 32'h44a51d43, 32'hc4630dda},
  {32'h42aa808f, 32'h44af9c30, 32'h4464a8ff},
  {32'h45141c7c, 32'hc2fe5265, 32'hc296b7c2},
  {32'h445c7b08, 32'h44a2ff50, 32'h44660ef9},
  {32'h43a2505f, 32'hc4ca31f8, 32'hc480ea3a},
  {32'h44f6c614, 32'h4251ebf6, 32'hc388efb4},
  {32'hc402de54, 32'hc42a5463, 32'hc53202b4},
  {32'h446067a0, 32'h4402e685, 32'h44a8b6f9},
  {32'hc3f71719, 32'h43640fe7, 32'h441eeed1},
  {32'h43f97c68, 32'hc455ebfa, 32'h448eb415},
  {32'hc4dffc3c, 32'h4263ab23, 32'hc36db20f},
  {32'h45295654, 32'h43444a18, 32'hbeaf27bc},
  {32'hc4d21c4a, 32'hc3a36017, 32'hc402991a},
  {32'hc2f99f2a, 32'h450dacea, 32'h42023752},
  {32'h4465114e, 32'h43946d1b, 32'h418ab27a},
  {32'h44b626a0, 32'h43c37a84, 32'h44b21253},
  {32'hc262b0fe, 32'hc393c50f, 32'hc5493e7c},
  {32'h443f12af, 32'h44999b3f, 32'h439f7120},
  {32'hc4f8eb0f, 32'hc487ae69, 32'hc256c0f4},
  {32'h44888189, 32'h4509fc17, 32'h415ff8e0},
  {32'h43f07673, 32'hc4802127, 32'hc398e912},
  {32'h444b573a, 32'h44d75987, 32'h4429a388},
  {32'hc37a349e, 32'hc5883903, 32'h4283ba23},
  {32'h4543eaa8, 32'hc10370f4, 32'h428a27dd},
  {32'hc57ea857, 32'h41a9e0ae, 32'hc3ba1b7e},
  {32'h455f3c69, 32'h42e05987, 32'h4388be41},
  {32'h449de418, 32'hc493bcf9, 32'hc4151e4a},
  {32'h432bfc2d, 32'hc5048f5c, 32'h44c47942},
  {32'hc36fddfe, 32'hc391db2c, 32'hc46dd328},
  {32'hc4c2e002, 32'h439d7d0a, 32'h444c0234},
  {32'h43ef64ed, 32'hc377f403, 32'hc503b3a4},
  {32'h4483767c, 32'hc33d458b, 32'h436a6978},
  {32'h440be254, 32'hc1a7ae92, 32'hc520a6c7},
  {32'hc4473b74, 32'h442171c9, 32'h44910fb7},
  {32'h430fe06c, 32'hc40135bf, 32'hc3a44b01},
  {32'h43b0107a, 32'h45122c55, 32'h441fce08},
  {32'h43d197aa, 32'h44052bbc, 32'hc4bc2186},
  {32'hc247987c, 32'h441be7d6, 32'hc3c89b9c},
  {32'h4437b56b, 32'hc3310414, 32'hc45129fc},
  {32'hc3b4f303, 32'h44fb4c9f, 32'h436a6f92},
  {32'hc409863b, 32'hc385d32e, 32'hc42a2d9c},
  {32'hc388d690, 32'hc11d14f5, 32'h4535df1d},
  {32'h44f70a50, 32'hc41fb247, 32'hc27c7fb4},
  {32'h439b4c31, 32'h44809e15, 32'h4411c223},
  {32'h441298ac, 32'hc5207c2f, 32'h4381416b},
  {32'hc540770b, 32'h424aa5fb, 32'h4282c0ee},
  {32'hc48f86fa, 32'hc22af154, 32'h4328edfa},
  {32'hc496ea4a, 32'h44363d77, 32'hc434cca4},
  {32'h4491d418, 32'hc4c0ea15, 32'hc3b103e0},
  {32'h44afc584, 32'hc1297dc6, 32'hc33d4518},
  {32'hc35ca500, 32'hc1de449f, 32'hc26276fe},
  {32'hc54e1da9, 32'hc3d53994, 32'hc386c516},
  {32'h4509ce4e, 32'hc3cd34d0, 32'hc2e603b1},
  {32'hc440141b, 32'h43c3544f, 32'hc374b531},
  {32'hc40aff0c, 32'h4309e1a5, 32'hc4f57040},
  {32'h4550d29c, 32'hc2f4c015, 32'h4399faca},
  {32'hc33d49f1, 32'h44b79d81, 32'h43ac9f6a},
  {32'h413b1b80, 32'hc48b75b0, 32'h428a43c5},
  {32'hc50352bc, 32'h427815f4, 32'h430cd0ac},
  {32'hc4a95f0e, 32'hc3fd82c5, 32'hc2fcd41d},
  {32'hc4620977, 32'h45234998, 32'h43c2d12b},
  {32'h446c8662, 32'hc49cb7fe, 32'h43b89623},
  {32'hc4c48205, 32'h42ea9e99, 32'h42bdf46d},
  {32'h4527ae73, 32'hc183ba2c, 32'h430a7705},
  {32'hc31cce20, 32'h4376770a, 32'h439c754a},
  {32'h42c3b6ba, 32'hc363f686, 32'hc44fe770},
  {32'h43dbe9d8, 32'h44849de3, 32'h441333e0},
  {32'h442e4ca1, 32'hc421c8b2, 32'hc44d6b51},
  {32'h422aa51b, 32'h44735957, 32'hc35e2ba8},
  {32'h42bd5015, 32'h434cc124, 32'hc4f2e7a5},
  {32'hc383678c, 32'hc3860d14, 32'h451464e6},
  {32'hc4000c2a, 32'h422d21ed, 32'hc2ee49fe},
  {32'hc3cb08fb, 32'h439a44e7, 32'h448add5e},
  {32'h45112354, 32'hc3c9899d, 32'hc46225aa},
  {32'h43d26bdc, 32'h449bb4a6, 32'hc390a7d2},
  {32'h43504356, 32'hc32720d4, 32'h4399f992},
  {32'hc41a4059, 32'h446c7a7e, 32'h44e98ab9},
  {32'h4327f30f, 32'hc4de2b24, 32'hc455a75e},
  {32'hc4ad3647, 32'h44deace5, 32'h4431d277},
  {32'hc24d6546, 32'hc5369a61, 32'hc334820b},
  {32'h45602842, 32'hc3a4faf6, 32'hc3186a56},
  {32'hc4a33e82, 32'h431fa8af, 32'h4481e3cc},
  {32'h44e572ec, 32'hc1ceb77c, 32'h4435c0fd},
  {32'hc45cd663, 32'hc27138c2, 32'hc40a6476},
  {32'h4485fefa, 32'h44b7bf58, 32'hc199ce58},
  {32'hc4df233c, 32'hc31bb877, 32'h43919008},
  {32'h454150f0, 32'h444c0fe0, 32'hc3adeec8},
  {32'hc42d91a6, 32'hc53caa42, 32'hc3c55520},
  {32'h4489c434, 32'h4356d3be, 32'h435af5cc},
  {32'h43829ec8, 32'h43cf7869, 32'hc48d45d7},
  {32'h452553c4, 32'h429cf730, 32'hc23b1932},
  {32'h449709d1, 32'h4344aac1, 32'h4351c851},
  {32'h4466e7de, 32'h43acef56, 32'h44665582},
  {32'hc4da4003, 32'hc35ca4f5, 32'hc435269a},
  {32'h439f12df, 32'h4486b240, 32'h434102fb},
  {32'h42880f30, 32'hc4512d4e, 32'hc47d59d6},
  {32'h43ce02de, 32'h4526ebaf, 32'h4294f39a},
  {32'h44cfe01c, 32'hc3b61abe, 32'hc2db0202},
  {32'h4514eece, 32'h447379db, 32'h441d5996},
  {32'hc58ae590, 32'h431f66fb, 32'hc3b9eec5},
  {32'h43d32c1a, 32'h4361312d, 32'hc298bddd},
  {32'hc3b9bd5c, 32'hc40ef3be, 32'hc48cccc0},
  {32'hc1f3a320, 32'h450f6091, 32'h410501d4},
  {32'hc4e25b0a, 32'h42bf278b, 32'h418a86b8},
  {32'hc3a8c92d, 32'h42720cef, 32'h4508eeed},
  {32'hc40af09c, 32'hc2d505f6, 32'hc53da8a8},
  {32'hc308df24, 32'h44c1092b, 32'h43de62dd},
  {32'hc4ec7ee6, 32'h43b6cb30, 32'hc2f186e6},
  {32'hc414551c, 32'hc45d414b, 32'hc39d4c6f},
  {32'h43c7e54f, 32'h44fe2ae1, 32'hc310483f},
  {32'hc3f3026c, 32'hc3bf030e, 32'h438bda2a},
  {32'h44cf23b1, 32'h44aae904, 32'hc363e4d6},
  {32'hc51e737c, 32'hc398ae56, 32'hc220a700},
  {32'hc2bf1398, 32'h43b6bf92, 32'hc332eadc},
  {32'hc5416461, 32'h433b557b, 32'hc2553f69},
  {32'hc16f6890, 32'h448da6d1, 32'h44659d27},
  {32'h439654d4, 32'h43802147, 32'h44a38069},
  {32'h43d486bd, 32'h43e0a90a, 32'h433b0049},
  {32'hc3447f39, 32'hc439ca7f, 32'h42e8b259},
  {32'hc483cc80, 32'h43dce2a9, 32'hc29a3b18},
  {32'hc2df3f51, 32'hc4dd55bc, 32'h43bd67d5},
  {32'h44280735, 32'h43fb9bd2, 32'hc3edf74d},
  {32'hc528d495, 32'hc3bc31fc, 32'hc2daceb1},
  {32'h4499d830, 32'h43316b14, 32'hc4401e31},
  {32'hc460fcca, 32'hc449748c, 32'hc408929e},
  {32'hc42f7008, 32'h446d9119, 32'hc2eef3fc},
  {32'hc4deb9ae, 32'hc45d085d, 32'h44310c8e},
  {32'h44451f2d, 32'h44b18513, 32'hc51925f4},
  {32'h4404b011, 32'hc50009ee, 32'h434f6fe4},
  {32'h4477f12f, 32'h44a599aa, 32'hc30bbc0e},
  {32'hc2b6227b, 32'hc3eed196, 32'h44907dcf},
  {32'hc37887ac, 32'h42b5775b, 32'hc3f06ae3},
  {32'hc4aca1a0, 32'h42b58709, 32'h4536da78},
  {32'h435d201c, 32'hc325751b, 32'hc56cafcf},
  {32'h4537e436, 32'hc4799fc7, 32'hc402da86},
  {32'hc5282461, 32'h44078737, 32'h42e4b581},
  {32'h44258070, 32'h4386fdc0, 32'hc3844a54},
  {32'hc418030e, 32'h450e011c, 32'hc3f0d702},
  {32'h411d2200, 32'hc51ebbdf, 32'hc36aa293},
  {32'hc412912b, 32'h44b4b205, 32'h42e43780},
  {32'h453b5f08, 32'h43e2cc31, 32'h434ec185},
  {32'hc4ae9e72, 32'h4496f9e1, 32'h44817e70},
  {32'h43a11022, 32'hc446865d, 32'hc3570a80},
  {32'hc3f1b77c, 32'hc408c041, 32'h44a73b0b},
  {32'h4514fb7b, 32'hc3589e6b, 32'h43b313b4},
  {32'hc492777c, 32'hc33b7e31, 32'hc38dac23},
  {32'h44245091, 32'hc2d9dff0, 32'h44eeef47},
  {32'h3fd0d780, 32'h4508ff13, 32'hc4229712},
  {32'h4503ad46, 32'h43b84e91, 32'h42af2e94},
  {32'hc2963440, 32'hc3c92a72, 32'hc5288831},
  {32'h451a7afa, 32'hc469a5dd, 32'hc3caab31},
  {32'hc454de43, 32'h439e2fe0, 32'hc434acae},
  {32'h43d22679, 32'hc4a12e40, 32'h44ab3270},
  {32'hc4a0264b, 32'h44554d14, 32'hc50ea997},
  {32'h4500af9f, 32'hc38c6d18, 32'hc2aa407c},
  {32'hc44c3448, 32'h4430eb02, 32'hc4f9694c},
  {32'h43cc73fe, 32'hc42797e0, 32'h44d080a1},
  {32'h43d33888, 32'hc3192464, 32'hc501207e},
  {32'h44d63a28, 32'h435fd62a, 32'h4467b2f0},
  {32'hc5884e4d, 32'h42ee0adb, 32'hc427eb1c},
  {32'hc486a166, 32'hc3a53288, 32'h439fe43f},
  {32'hc3885ea4, 32'h44b467f0, 32'hc4c61bae},
  {32'hc3fb0134, 32'h44fafba0, 32'h450f947a},
  {32'hc5118eab, 32'h4367653b, 32'h43e8a5a7},
  {32'hc525831e, 32'h43026057, 32'h42de7aba},
  {32'h4484949d, 32'hc468cc0c, 32'h4449e274},
  {32'hc2e97740, 32'h449f9144, 32'hc46aa55a},
  {32'hc2d2bd36, 32'h43b332e8, 32'h44e2e740},
  {32'hc40e8a25, 32'hc33767f3, 32'hc369f28b},
  {32'h431be96d, 32'hc47f0c0c, 32'h450bd0bd},
  {32'h43cd4542, 32'hc4e85629, 32'h44b70c14},
  {32'hc41f4f25, 32'h439e8c28, 32'hc4949049},
  {32'hc44a285d, 32'hc2c3b36e, 32'h4462d159},
  {32'h43fe4d3d, 32'hc465b1da, 32'h439ac42a},
  {32'hc4c151b1, 32'h433ebbb9, 32'hc325bedf},
  {32'h43a2255c, 32'hc3102eb8, 32'h446cd950},
  {32'hc085c0c0, 32'h438ac302, 32'h42da3cc1},
  {32'h4412273e, 32'h4356d209, 32'h44f7a411},
  {32'hc40bd74a, 32'hc1debaf2, 32'hc4e3ef09},
  {32'h453dfb45, 32'hc1f68f61, 32'h44545639},
  {32'hc5015ca1, 32'hc39fe47a, 32'hc436f73e},
  {32'hc33db910, 32'h42a1fee1, 32'hc2e180fd},
  {32'h4384a771, 32'h44e88b59, 32'hc2f1b620},
  {32'h4501a726, 32'hc455a02f, 32'hc24642af},
  {32'h42837020, 32'h451c2fa0, 32'hc37d3123},
  {32'h431c8f9e, 32'hc4e645b5, 32'hc2d12e02},
  {32'hc49102ec, 32'h45103b67, 32'h440c9053},
  {32'hc299d9e0, 32'hc4cb18cb, 32'h4387625f},
  {32'h438c55f2, 32'h44aa8b8e, 32'h44a8f258},
  {32'h42dc5408, 32'h44142592, 32'hc48995cd},
  {32'hc3cce927, 32'h44ff2d17, 32'h4472405b},
  {32'hc4c099ff, 32'hc32cf373, 32'h41dc9c33},
  {32'h438f6354, 32'h44e94c67, 32'hc2ea9555},
  {32'h44951bdb, 32'hc2770f72, 32'hc305ce9a},
  {32'h44d0c322, 32'h44ac85ff, 32'hc27e9d9c},
  {32'hc50a2348, 32'hc46af9fd, 32'h443c8abf},
  {32'hc5010435, 32'hc266fcc0, 32'hc3d9cf21},
  {32'h42716da8, 32'h422a43da, 32'hc472cb97},
  {32'h446de4ab, 32'h43b27875, 32'hc39ad6a5},
  {32'h43915d64, 32'h44b15bca, 32'hc4e27236},
  {32'h44c8d2d3, 32'h42744bbc, 32'hc364fda6},
  {32'hc4412de0, 32'hc3cc45c2, 32'h44a821c6},
  {32'h44442fbb, 32'hc12cfc0b, 32'hc43bf76a},
  {32'hc3babab0, 32'hc334eafc, 32'h44d763be},
  {32'h445433f0, 32'hc456ba76, 32'hc44f2314},
  {32'h43dca4f6, 32'hc427db86, 32'h42b28409},
  {32'h456c41ea, 32'hc2c05e55, 32'h440d4011},
  {32'hc4abb76d, 32'h44132839, 32'h43c980f3},
  {32'hc49b85a0, 32'h43bcce22, 32'hc30e4da7},
  {32'hc390b640, 32'hc5265ae6, 32'hc3613027},
  {32'h45113eb1, 32'hc3998169, 32'hc0bee094},
  {32'h44cd8660, 32'hc2fd150e, 32'h43e32c4b},
  {32'h44e357e7, 32'h44490f0d, 32'h433ffba6},
  {32'hc4061770, 32'hc4edbad6, 32'hc28a43d8},
  {32'hc42759d3, 32'h44562933, 32'hc338d1f4},
  {32'h433fdb90, 32'hc38d2ca4, 32'hc2b63d4b},
  {32'hc43febce, 32'h43c2a4d1, 32'hc4a3aae0},
  {32'h43a97290, 32'h449bc47f, 32'h4448ffeb},
  {32'h43c1b25a, 32'hc393b187, 32'hc3bf256d},
  {32'h4461244c, 32'h44eca6b6, 32'h42088817},
  {32'hc4276eaf, 32'hc5028c76, 32'hc38574e9},
  {32'hc332f26e, 32'hc3c8e56a, 32'h448b7875},
  {32'h41858600, 32'hc3ea5143, 32'hc5285f37},
  {32'h440b9331, 32'hc3412791, 32'h44a1ee4e},
  {32'h43a5832e, 32'hc4315ad1, 32'hc41d5a87},
  {32'h449782ce, 32'h42a92c5d, 32'h43a7e000},
  {32'hc32432e8, 32'hc4b623ac, 32'hc48120d0},
  {32'h4540a574, 32'hc3868bdd, 32'hc2a80564},
  {32'hc3afc9f0, 32'hc50dc126, 32'hc41351ed},
  {32'h44115390, 32'h4393d437, 32'h44195eb0},
  {32'hc34c0750, 32'hc40c8498, 32'hc2891be0},
  {32'h43588466, 32'hc05cfca8, 32'h453c1096},
  {32'hc43e04ef, 32'hc414716a, 32'hc50b14cb},
  {32'h4479a8db, 32'h447fb70f, 32'h4391dd37},
  {32'hc5837704, 32'h42ba2aa2, 32'h432f8c2a},
  {32'h443ce3ad, 32'h452ad375, 32'h41f669f9},
  {32'h44bfe5ad, 32'hc2723306, 32'h4326ef41},
  {32'hc29ba0a6, 32'h4581d194, 32'hc26fdc86},
  {32'hc32a41e0, 32'hc4264b70, 32'hc299d033},
  {32'hc43a115e, 32'h41dbcff9, 32'h43c6132f},
  {32'hc56ce6b5, 32'hc3510a79, 32'hc3441fee},
  {32'h457ce1dd, 32'hc2074fb9, 32'h438be317},
  {32'hc35dfd4e, 32'h4411af47, 32'hc51ea2fd},
  {32'hc4674f1d, 32'h440e0570, 32'hc3266192},
  {32'h43e01658, 32'hc3b71efd, 32'h440bc723},
  {32'hc343ad68, 32'h44e76f54, 32'h44b5a609},
  {32'h4372bee4, 32'hc5163560, 32'hc376f3c0},
  {32'h44ab536a, 32'hc2e429c4, 32'h4412bfa6},
  {32'h44f44a23, 32'h42a705b2, 32'hc46fdad4},
  {32'h42411c0d, 32'h44839ef7, 32'h4509045b},
  {32'h444d6df0, 32'hc397c29b, 32'hc4d1b100},
  {32'h43af1883, 32'h4506b67c, 32'h43b47f4f},
  {32'h445559da, 32'h4447e504, 32'hc444da3e},
  {32'h43baa108, 32'h448b5edb, 32'hc1e70de7},
  {32'h45559792, 32'hc34761b8, 32'hc02a05b2},
  {32'hc4162c2d, 32'h44c23ae8, 32'h4428d884},
  {32'hc411c5f3, 32'hc4511cbe, 32'hc3d9ce63},
  {32'hc1d830b8, 32'h43987144, 32'h4572274d},
  {32'h4496d593, 32'hc4b991eb, 32'hc433dd4e},
  {32'h4418b502, 32'h43750fc8, 32'h4404d960},
  {32'h4496faf3, 32'hc4d18064, 32'hc3bc17f9},
  {32'hc4edac40, 32'h44a1ffcd, 32'h4389fb04},
  {32'h44c52fdc, 32'hc33b8e42, 32'h413ce6a8},
  {32'h433c63e4, 32'h448a52f3, 32'hc417c804},
  {32'h440e255d, 32'hc563ad94, 32'h43068a2a},
  {32'hc507fea3, 32'h4199f874, 32'hc104af67},
  {32'h442ca8f0, 32'hc2c4dbd2, 32'h438839f0},
  {32'hc4c385ca, 32'hc3fd92cc, 32'hc4103678},
  {32'hc47665f0, 32'h434fea35, 32'hc39d0a40},
  {32'h452fdd8e, 32'h4367cde4, 32'hc3374b5b},
  {32'hc4b8ccbc, 32'hc21573fe, 32'hc3c55c07},
  {32'hc33dc920, 32'h42f0765e, 32'h44c96895},
  {32'hc516b13b, 32'hc427dbb1, 32'hc43355e6},
  {32'h44d33581, 32'hc4b2e249, 32'h430ba67c},
  {32'hc49f14ad, 32'h423822e4, 32'h420f7d08},
  {32'h4317b8e2, 32'hc35c3738, 32'hc326ee4d},
  {32'hc3a48000, 32'h4579b3f4, 32'h438adb2c},
  {32'h43206a0e, 32'hc5023b77, 32'h43d1ef0e},
  {32'h44e1a036, 32'hc434f22a, 32'hc336a1f5},
  {32'h448385e8, 32'h43138f52, 32'h43c399aa},
  {32'hc3c8ba04, 32'hc48a938d, 32'hc502dc51},
  {32'hc2ba0aac, 32'h43051709, 32'hc413e4e9},
  {32'hc53b6f7d, 32'hc34dd100, 32'h439de2da},
  {32'h43e6aaa6, 32'hc4328d6b, 32'hc54c41f8},
  {32'hc49632c3, 32'hc289d1f4, 32'h431c5106},
  {32'h40c98d80, 32'hc51b2931, 32'h434fd161},
  {32'h43add885, 32'h44b5cfae, 32'h44761f71},
  {32'h45162bd0, 32'h42a4fa21, 32'hc433d55f},
  {32'hc54ba878, 32'h43480c10, 32'h445d4678},
  {32'h44ed58d7, 32'h43a378d5, 32'hc463b2ac},
  {32'h430a85b0, 32'hc39a16ce, 32'h44c925e9},
  {32'h44107bd7, 32'hc49388a2, 32'hc3834a0c},
  {32'hc424b91a, 32'h42af4312, 32'h446756f1},
  {32'h43cf86b7, 32'hc4b9d0ec, 32'h41f7e8d6},
  {32'hc556cf71, 32'h44963958, 32'hc2d1ff59},
  {32'h448ba4e2, 32'hc4422633, 32'hc45641d9},
  {32'hc3f70398, 32'h44731ea7, 32'hc513f0ab},
  {32'hc55f5bd5, 32'h440f3a0a, 32'h41dd45c4},
  {32'h43aa6f55, 32'hc4034544, 32'hc4a7c1b6},
  {32'hc475fad9, 32'hc501ed3f, 32'hc345ba54},
  {32'hc29cdce2, 32'h44ee42cb, 32'h4247b7d2},
  {32'hc550328e, 32'hc2915334, 32'h4362ff35},
  {32'h43a56ca2, 32'h455a4ed6, 32'h42c25d86},
  {32'hc3f8edca, 32'hc5329f1e, 32'h43d06eb0},
  {32'hc49a309a, 32'h42224e0a, 32'h43675a30},
  {32'hc465c9b1, 32'h43c20907, 32'h42e3c8dc},
  {32'h44de488f, 32'hc3f122ad, 32'h43de37bf},
  {32'hc4d78f5d, 32'h43834694, 32'h4320b6c6},
  {32'h43a4a160, 32'h42dcbbc4, 32'h451810de},
  {32'hc494add3, 32'hc226974d, 32'h42b79f48},
  {32'h44d42b21, 32'h43cef057, 32'h41d43d16},
  {32'hc3dee120, 32'hc38886f4, 32'hc3d6afc7},
  {32'h44987342, 32'h4421ee78, 32'h436fc512},
  {32'h42954734, 32'hc3a0a99d, 32'hc4b1c978},
  {32'h4515411f, 32'h4426f781, 32'h43a26863},
  {32'hc46851fa, 32'h444d5278, 32'hc49ebed3},
  {32'hc507ee34, 32'hc3430ced, 32'h4313abde},
  {32'h431922f8, 32'hc55fe565, 32'hc303536a},
  {32'h43933ad8, 32'h43e4ba25, 32'h44bcbe3a},
  {32'hc2591b96, 32'hc4820e46, 32'h438774c8},
  {32'hc3b8c9e1, 32'h43923247, 32'h44c4cd9e},
  {32'hc439ba1c, 32'hc3ee4b73, 32'hc3bec247},
  {32'h44a53fbd, 32'hc3bfaede, 32'hc33ae5bf},
  {32'h44b2cc96, 32'hc2a248d0, 32'hc2cbb3cb},
  {32'hc4432252, 32'hc1fc5528, 32'hc49700ed},
  {32'h41cb41bc, 32'h4554aa48, 32'h44020178},
  {32'hc5061058, 32'h4390f47b, 32'h427407ff},
  {32'h44080dce, 32'h451ff2d3, 32'hc28be738},
  {32'hc4725573, 32'hc4be58b1, 32'h430e73c8},
  {32'h4553e48c, 32'hc36cae44, 32'hc441da3d},
  {32'hc50fd1da, 32'hc3beb34f, 32'hc34be677},
  {32'h44878502, 32'hc3efb320, 32'hc2aa3b45},
  {32'h44c0e353, 32'hc40d0cfa, 32'h43ca51f8},
  {32'h4380b8a6, 32'h450a155e, 32'hc2c3cd8a},
  {32'hc4b8dba5, 32'hc31ef985, 32'h44429063},
  {32'hc31941d9, 32'h4300f3a5, 32'hc3de7f8a},
  {32'hc3da8710, 32'hc402da40, 32'h42ca1d98},
  {32'h43ac613a, 32'h441121d1, 32'hc4d00b1f},
  {32'hc4e3164b, 32'hc1542b8f, 32'h43f5edc9},
  {32'h43b20ad0, 32'h43fc4377, 32'hc3567152},
  {32'hc307723c, 32'h4294b566, 32'h451d9ddb},
  {32'h450ebcb3, 32'hc3e072fc, 32'h42efb490},
  {32'hc445a626, 32'hc3ea2274, 32'h44b04b1c},
  {32'h4326fd90, 32'h44a26d0c, 32'hc4f2edad},
  {32'h44a1b5d6, 32'hc41563a0, 32'hc3fe31f3},
  {32'h447ecaa2, 32'h4330cfe9, 32'hc3f3acb6},
  {32'hc54edcfa, 32'hc39aa95f, 32'h42c150f9},
  {32'h4482e3e3, 32'h435946cc, 32'hc42756c2},
  {32'hc4fa9102, 32'hc3ffcdaf, 32'h442ff0a5},
  {32'h42ef02bd, 32'hc3bfb887, 32'hc53a194a},
  {32'h43f51468, 32'hc3232216, 32'hc4918092},
  {32'hc36a82d0, 32'h4547591e, 32'h43d5b272},
  {32'hc42dab02, 32'hc452c216, 32'h43a72691},
  {32'hc28715c0, 32'h44c86e7a, 32'h439c7f81},
  {32'h4446a5e0, 32'hc446991d, 32'hc1df3ef8},
  {32'h433f38a4, 32'h44aaf8c1, 32'hc3a3d240},
  {32'h4540787a, 32'h42b61dad, 32'hc3ace8bd},
  {32'hc495cf4d, 32'h43419ec8, 32'h4186c1e5},
  {32'h455ffc6f, 32'h440dc80a, 32'h444eb12e},
  {32'h43d7ae8a, 32'h451809b1, 32'hc2ae67f8},
  {32'h441d6f6e, 32'hc309ae00, 32'h443c039e},
  {32'h43393770, 32'h442359de, 32'hc468896c},
  {32'h44fa051c, 32'h43c04091, 32'h43fa7474},
  {32'hc508a5aa, 32'hc3870070, 32'h4192ff2a},
  {32'hc47a8d4a, 32'hc33f29ba, 32'h44883efb},
  {32'hc47875dc, 32'h43f902fa, 32'h439fc6fe},
  {32'h44f26e5b, 32'hc45b95fb, 32'h4296993b},
  {32'h4507509f, 32'hc2818aff, 32'hc38057ca},
  {32'h44c95fc6, 32'hc43c2ea0, 32'h44cfdc45},
  {32'hc48c5aac, 32'h4445c766, 32'hc4c05a0c},
  {32'hc3300217, 32'hc3fe24cb, 32'h44ce0f42},
  {32'hc4d17610, 32'h441f71f9, 32'hc41aebed},
  {32'h42b7bccd, 32'hc52a7205, 32'h43df7272},
  {32'hc47b7e6e, 32'h443855ac, 32'hc3cdde2b},
  {32'h431a4800, 32'h448d4c97, 32'h4350b8a6},
  {32'hc4567829, 32'hc459e5f2, 32'hc4295fbc},
  {32'h456703fb, 32'h42955a49, 32'hc47ed810},
  {32'hc36fb902, 32'hc4ebc659, 32'hc4e12733},
  {32'h4469d2df, 32'hc324e840, 32'h44050630},
  {32'hc321d472, 32'h429f87cf, 32'h433a0cce},
  {32'h44b71e1c, 32'h3ff8e98a, 32'h4317b085},
  {32'h434e3020, 32'hc4a82e9c, 32'hc2cef514},
  {32'h43a92e38, 32'h45201734, 32'hc31020b9},
  {32'h43841a83, 32'hc2bc6e52, 32'h4473424d},
  {32'hc4628a76, 32'h42ed9f9c, 32'hc4ac0e0d},
  {32'h446e81b5, 32'hc4ba1cf6, 32'h442864c1},
  {32'h43d8753a, 32'hc3db6018, 32'h4514e628},
  {32'hc389e216, 32'hc4784fb1, 32'hc502a2ce},
  {32'hc22d64d9, 32'hc3e97651, 32'h448e8f19},
  {32'h43cdd08e, 32'hc473ce00, 32'hc3363965},
  {32'hc42c8274, 32'hc3020639, 32'hc4b66adb},
  {32'h452b063e, 32'h42a5d69f, 32'hc33b3d69},
  {32'h44f7c5ca, 32'h438185cb, 32'h43077abe},
  {32'h439fa7fc, 32'hc45b626c, 32'h440cc820},
  {32'h433bf176, 32'h454088d8, 32'h43666a62},
  {32'h4382d51c, 32'hc42f328d, 32'h445553d8},
  {32'hc4edd8ac, 32'h4284c2b4, 32'hc30d0e1d},
  {32'hc3b33ce0, 32'h43a02b78, 32'h443b426e},
  {32'hc3dd18d0, 32'h445b72a6, 32'h436fbbea},
  {32'h452e8626, 32'hc43cac44, 32'hc2e1d773},
  {32'hc501cf36, 32'h4335473a, 32'h440c00b7},
  {32'hc4d7a681, 32'h42f65cf9, 32'hc2b7fd02},
  {32'hc4958aa1, 32'h44bfb4b1, 32'hc351b5aa},
  {32'h44252d17, 32'hc50d89af, 32'hc3b60a83},
  {32'h43db2cde, 32'h432f741c, 32'hc2e41922},
  {32'hc4088568, 32'hc4887d9d, 32'hc5067f60},
  {32'h43045d33, 32'hc472be57, 32'h44bddf9a},
  {32'hc3f29306, 32'hc49d5368, 32'h440b0d47},
  {32'h44c0eb6e, 32'h43ba05be, 32'h42cbe6b8},
  {32'hc393ac40, 32'h43c709dc, 32'h422ac4f6},
  {32'h44c3698d, 32'h440ae42d, 32'hc42acfd6},
  {32'hc31c5708, 32'h432b78a7, 32'h44f1c819},
  {32'h446664ab, 32'h438522e8, 32'h43d13ce4},
  {32'h450ab132, 32'hc31990e4, 32'h436aef8d},
  {32'hc417c4b5, 32'h44238de8, 32'h44008ce8},
  {32'h44180dad, 32'h4435efa0, 32'hc4b9610f},
  {32'h42e0a097, 32'h41c409b3, 32'hc521a986},
  {32'h43042360, 32'hc4d8ff69, 32'h41a5c8ba},
  {32'h4454798c, 32'h43881622, 32'h420bca1f},
  {32'hc43769ea, 32'hc4b4dc94, 32'h42f1dbf9},
  {32'h453ff756, 32'h4387d17a, 32'h42f7c62f},
  {32'hc42be8cc, 32'hc42e7e43, 32'h4333a7a5},
  {32'h44ffd6ea, 32'hc2ef2733, 32'hc39bc7be},
  {32'hc4e70f87, 32'h43190e07, 32'hc33ee902},
  {32'h455cee46, 32'h43535322, 32'h4380e77d},
  {32'hc4d009e4, 32'hc4e450a9, 32'h43b0e996},
  {32'hc2626014, 32'h4570e4a7, 32'h439f67dd},
  {32'hc52807bc, 32'hc3b4e594, 32'hc19d26ba},
  {32'h43dba580, 32'h44f42864, 32'hc38e4aaa},
  {32'h43078c68, 32'hc542418b, 32'h429b17b8},
  {32'hc44a9831, 32'h429f8b47, 32'hc256d4c6},
  {32'hc35691c4, 32'h42c350b8, 32'h4465c029},
  {32'hc3ef83fb, 32'h444e33ea, 32'hc50230cb},
  {32'h42803a0e, 32'h44881edd, 32'h43d7ef22},
  {32'hc4999906, 32'hc2aa9030, 32'hc3b33b4e},
  {32'h440f5108, 32'hc0c37858, 32'h4469ec42},
  {32'hc43566e7, 32'hc2c728c0, 32'hc4af600a},
  {32'h4515d869, 32'hc2c63f1f, 32'hc35f6d44},
  {32'hc3b30eb8, 32'hc405691c, 32'hc52b6907},
  {32'h44159d68, 32'hc3ed7cd9, 32'h4476763d},
  {32'h44138245, 32'hc171f728, 32'hc2ff845c},
  {32'hc2acce17, 32'hc51be788, 32'h44e64310},
  {32'h4123c560, 32'hc5092eec, 32'hc382484d},
  {32'hc407d6db, 32'hc273d713, 32'h448c9206},
  {32'hc0acb8c0, 32'hc4ebdea6, 32'hc43ed303},
  {32'h44b2e8dd, 32'h442ebed3, 32'hc20feff4},
  {32'h432c7e1a, 32'hc32d1a69, 32'hc321e28a},
  {32'h438d1184, 32'h44c7ed75, 32'h44491b97},
  {32'hc30ef5d4, 32'hc3979f54, 32'hc51df4b5},
  {32'h434f9f9c, 32'h44882e9d, 32'h42df5161},
  {32'hc53e9123, 32'hc4262ad6, 32'hc3a902d1},
  {32'h430cef40, 32'h453dca4a, 32'h434aafe3},
  {32'hc31c5b57, 32'h42a999ca, 32'hc26bf791},
  {32'h43b15f47, 32'h44081ff0, 32'h43e348ab},
  {32'hc505f939, 32'hc41ee7c7, 32'h43245a40},
  {32'h45661d0e, 32'h443d77f2, 32'h437594f7},
  {32'hc5120efa, 32'h44014aef, 32'h43e8b24d},
  {32'h451a7790, 32'h432a506a, 32'h435de561},
  {32'h445109ae, 32'hc226f898, 32'hc46d3024},
  {32'h43a744d2, 32'h439e1ea9, 32'h44ba3f42},
  {32'hc424b942, 32'hc3727622, 32'hc383117a},
  {32'hc4d9133e, 32'h44368c19, 32'h44719fd5},
  {32'hc414280e, 32'hc4c5db0a, 32'hc4313b4a},
  {32'hc4c9e78a, 32'hc3845c85, 32'h437fd582},
  {32'h43d60f40, 32'hc483f2c7, 32'hc49f2fd2},
  {32'hc4200c3d, 32'h44033a3e, 32'h44dd08b8},
  {32'hc372ca8c, 32'hc39788cb, 32'hc3c82749},
  {32'hc4e6298e, 32'h42ef3daa, 32'h443ac90b},
  {32'hc3377db0, 32'h44ee6afe, 32'hc4facf86},
  {32'hc472727a, 32'hc3bd6e95, 32'h432a8e10},
  {32'h43829e90, 32'hc4878b19, 32'hc4884e2a},
  {32'hc48886c2, 32'h43c8829e, 32'h44275de6},
  {32'hc3a1b889, 32'hc5005d6a, 32'hc20ad8b9},
  {32'h44138334, 32'h448c8c5e, 32'h4536671d},
  {32'h4500f4db, 32'hc473671c, 32'hc40759a1},
  {32'hc40111e8, 32'h449bbaef, 32'hc1e5cbcd},
  {32'h440b8218, 32'hc4bcd5e6, 32'hc4819d4b},
  {32'hc3952158, 32'h45372812, 32'hc30a562a},
  {32'h44a5cd30, 32'hc377e06d, 32'h42da92a5},
  {32'hc42df202, 32'h454dae7c, 32'h4400e149},
  {32'hc10ade80, 32'hc54daa77, 32'h4393b4fe},
  {32'h44930978, 32'h4424eccc, 32'h432da76a},
  {32'h4368ac20, 32'h431c8f46, 32'h4284f124},
  {32'hc4444118, 32'hc4673502, 32'h4234bb6f},
  {32'h4554e051, 32'hc2543735, 32'h42bf42c0},
  {32'h42a77ff8, 32'hc2f0ea4e, 32'hc28b2fce},
  {32'hc4111ee8, 32'h42f3900c, 32'hc346e897},
  {32'h44f33adb, 32'hc28ab23e, 32'h43b1accf},
  {32'hc3d42806, 32'hc2d987de, 32'h44037951},
  {32'h452c9189, 32'hc37276dd, 32'hc3bd59aa},
  {32'hc4d42015, 32'h4417cc50, 32'h42a71e4f},
  {32'h4531aa7b, 32'h44287a02, 32'hc31f98da},
  {32'hc41a02ca, 32'h4521988a, 32'hc36eeeb2},
  {32'h41ec8d90, 32'hc5509589, 32'h42810b55},
  {32'h44a5c127, 32'hc3bdc0c8, 32'h4422644b},
  {32'h45198224, 32'h430d7b6d, 32'h40a647f5},
  {32'h428a9be0, 32'h438cf1f7, 32'hc43623c9},
  {32'h4507dce4, 32'hc28bb613, 32'h407dfa19},
  {32'hc2503f0e, 32'h44852312, 32'h449609e9},
  {32'h44835f34, 32'hc3a054ba, 32'hc3b97562},
  {32'h439365b5, 32'hc355d088, 32'h44e98cba},
  {32'h44a1f6e7, 32'hc3bb9d0a, 32'hc4bc148e},
  {32'hc4f18156, 32'h43783a86, 32'h4488499a},
  {32'hc3c9e1bd, 32'hc411949c, 32'hc3e7a817},
  {32'hc579a126, 32'hc38f92d1, 32'h440cb8c1},
  {32'h4540ab6d, 32'hc391ad37, 32'hc45551bb},
  {32'hc4d8bc85, 32'hc42008bb, 32'hc2367500},
  {32'h43d39b7a, 32'hc42abb4a, 32'hc4951d0e},
  {32'hc4e9f44a, 32'h43f84e10, 32'h4307fff4},
  {32'h44a876ea, 32'hc346ba39, 32'hbb920000},
  {32'hc4abf94c, 32'h44faee45, 32'h432f6f62},
  {32'h44d16e00, 32'hc3e355e9, 32'hc4b8c601},
  {32'h4496ef3e, 32'h431b2077, 32'hc4a4af4b},
  {32'hc505e873, 32'h42b4d3f1, 32'h44b6e8a3},
  {32'h44cd0d8c, 32'h433ff3c4, 32'h441fbf61},
  {32'hc4351eb3, 32'hc4bf0dcc, 32'hc384432c},
  {32'h444b4344, 32'h448b7107, 32'h4200100e},
  {32'hc4ae13d8, 32'h42508441, 32'hc3dd2e05},
  {32'h44a6669c, 32'h4504e2db, 32'h43b2294a},
  {32'hc4729cd0, 32'hc483944e, 32'hc3ba5fec},
  {32'h4426302a, 32'h44867858, 32'h41f4994c},
  {32'hc39fb03c, 32'hc47a44f4, 32'h4507d354},
  {32'h444e5922, 32'hc2c671ed, 32'hc4c4dbc8},
  {32'h4408c146, 32'hc36d95c3, 32'h43b258ea},
  {32'h42b7e020, 32'h44a0eea5, 32'h4462ce67},
  {32'hc4edcd95, 32'hc3cf7082, 32'hc3a0448d},
  {32'hc46cf263, 32'h42832036, 32'h4443135c},
  {32'hc5104167, 32'hc2f7db07, 32'hc42c856d},
  {32'h43beb020, 32'h43fd2062, 32'h45085515},
  {32'hc5072594, 32'hc41dccde, 32'hc3e7fd50},
  {32'hc39c9faa, 32'hc3106ccf, 32'h402aada9},
  {32'hc58a4f12, 32'hc2f90547, 32'hc0a186d8},
  {32'h45530e5b, 32'h43ed6cd1, 32'hc3ea5cda},
  {32'hc3fdd9ed, 32'hc50a7f9a, 32'hc4411f6b},
  {32'hc40d1365, 32'h449285fa, 32'h440cfbdb},
  {32'hc4834b2f, 32'hc41be914, 32'h42ac374b},
  {32'h42ecec30, 32'h43f9d940, 32'h452f2706},
  {32'hc3ced5b6, 32'hc504c2fe, 32'hc47939c8},
  {32'h446356ba, 32'h4499a84c, 32'hc3264406},
  {32'hc3960708, 32'h438c020a, 32'hc0a4ab90},
  {32'hc41dde73, 32'hc4c6a9e0, 32'hc39d832e},
  {32'h45477399, 32'h43bfbe55, 32'h43b02dd3},
  {32'hc482086f, 32'h43bbf61c, 32'h42b530e0},
  {32'h44f924ba, 32'h440b4284, 32'h42dd7b37},
  {32'hc37668ef, 32'hc504f6ea, 32'hc2eb56cd},
  {32'h43e3a1a6, 32'hc321348a, 32'hc309e363},
  {32'hc56ca73e, 32'hc2015648, 32'h42da364d},
  {32'h4515a26c, 32'h437f82a9, 32'h44a4d0cd},
  {32'hc2851862, 32'hc46a81f2, 32'hc3aa0e1f},
  {32'h44b5f383, 32'h440400de, 32'h432001c0},
  {32'hc1ad82d8, 32'hc44a122e, 32'h439ab913},
  {32'hc4e14cbf, 32'h4420aea0, 32'hc2b6f576},
  {32'hc3acbc10, 32'hc5111686, 32'h4431ff01},
  {32'h441210da, 32'h4482698a, 32'hc401c2df},
  {32'hc519c82a, 32'hc393f8bd, 32'h4296a341},
  {32'h4413285c, 32'h43926535, 32'hc3ca4d0f},
  {32'hc4b32d74, 32'hc3b59854, 32'h4424b3a0},
  {32'hc49db28d, 32'hc280d6b3, 32'hc4253328},
  {32'hc4403156, 32'hc47633a6, 32'h4492ce4c},
  {32'hc2eca9c0, 32'h44a7a92b, 32'hc492e637},
  {32'hc1072d98, 32'hc4865866, 32'h444be572},
  {32'h44a0bb13, 32'hc397bb58, 32'hc417ca93},
  {32'hc534f240, 32'h4386712a, 32'h4222750b},
  {32'h452cfc84, 32'h4320dcdd, 32'hc3a03350},
  {32'hc3fff68e, 32'h446e0eb0, 32'h452b682c},
  {32'h448f0aeb, 32'hc3d6d18b, 32'hc42b008e},
  {32'h437d4ee5, 32'hc50388c8, 32'hc333a689},
  {32'hc450f404, 32'h44a7dd93, 32'h432e3220},
  {32'h4409fb2a, 32'hc507e377, 32'h43bbadea},
  {32'hc3aa650c, 32'h43581dc7, 32'h43cb9025},
  {32'h43aac0d7, 32'hc55a0fc7, 32'h434dfeb1},
  {32'hc346062a, 32'h440e9e52, 32'hc291c86f},
  {32'h440df274, 32'hc3804888, 32'hc293069f},
  {32'hc500b8a9, 32'h438a53c8, 32'h428484ac},
  {32'h41f77440, 32'hc429221c, 32'h43d68f55},
  {32'h434a00a0, 32'h45289982, 32'h438e2217},
  {32'h4504a386, 32'hc30d221b, 32'h3f88e25b},
  {32'h449af90a, 32'h421b5750, 32'hc41af99d},
  {32'h43d817e2, 32'hc3e7eed6, 32'h444551b8},
  {32'hc516ba4c, 32'h43ae319e, 32'h42179bac},
  {32'hc34b14ea, 32'h444baf76, 32'h450cefbd},
  {32'hbfbcc800, 32'h438a4f09, 32'hc4377ccd},
  {32'h43e30c48, 32'h43307b34, 32'h44f25960},
  {32'hc451adc5, 32'hc39fab53, 32'hc422e0ec},
  {32'h42e2f798, 32'hc520e3ec, 32'h43e846e3},
  {32'h42b16d80, 32'h453bd6b9, 32'hc32be064},
  {32'hc48a379e, 32'hc31318d6, 32'hc31bd52c},
  {32'hc3dde6a7, 32'h44b6b25c, 32'hc458612e},
  {32'h43b74aea, 32'hc380893c, 32'h4487bb60},
  {32'h4421e205, 32'h43a41734, 32'hc302d12b},
  {32'h448307ab, 32'h443484c6, 32'h4535fbf4},
  {32'hc4ac74d4, 32'h426d84e9, 32'hc50ef831},
  {32'h43957290, 32'hc2b2e8d2, 32'h43086ab2},
  {32'hc27d192e, 32'hc469c65d, 32'hc50936ca},
  {32'h43d35cd4, 32'hc4c6e72f, 32'h448cebbd},
  {32'h431d67d4, 32'h434cdb16, 32'hc4429016},
  {32'h43bdf476, 32'h438f3797, 32'hc482dcc0},
  {32'h43c8fb2a, 32'h4284b056, 32'h450352aa},
  {32'hc3eb190b, 32'h4492be90, 32'hc44abf02},
  {32'hc4ac4457, 32'hc390758f, 32'h4463c19c},
  {32'hc4981665, 32'h43f61dcf, 32'hc44ae82c},
  {32'h44556eda, 32'hc4ec397d, 32'h43857b9d},
  {32'hc40436ac, 32'h43c640fc, 32'h4520dccb},
  {32'hc54a1236, 32'hc2e3b827, 32'hc3892348},
  {32'h445482f6, 32'hc4260c37, 32'h437fc9cd},
  {32'h4516e855, 32'h4373352c, 32'h42c7c041},
  {32'h433bbce0, 32'h44954326, 32'hc4590b46},
  {32'h452b42e4, 32'hc2ca6216, 32'h43c18d57},
  {32'h419d5a18, 32'h44b70a28, 32'h42f643ec},
  {32'h44f37d62, 32'hc35be344, 32'h445774c2},
  {32'h43b6285f, 32'hc2a40af6, 32'hc512c990},
  {32'h449afb9b, 32'hc41f800a, 32'h418d17d4},
  {32'hc38e5b34, 32'hc48c9181, 32'hc41eb073},
  {32'hc386c7f3, 32'h44453b7f, 32'h440bab48},
  {32'h43241a84, 32'h44f66133, 32'h4395f5de},
  {32'h42986064, 32'hc56d9425, 32'h4379edb5},
  {32'hc472282e, 32'h451ac602, 32'hc31d389d},
  {32'h436f4ae8, 32'hc49d2c3a, 32'h43504933},
  {32'hc24d9490, 32'h452986db, 32'h4337a72a},
  {32'h4404f32e, 32'hc4f6d863, 32'h424e499a},
  {32'h43769d5b, 32'hc34b3865, 32'h43c70835},
  {32'h42b67133, 32'h447ad9f2, 32'hc4bcacf0},
  {32'hc395f138, 32'hc3f3e1c8, 32'h44879502},
  {32'hc5161598, 32'hc4010a19, 32'hc31d9e84},
  {32'h419a55e0, 32'h43364433, 32'hc4cb4481},
  {32'h43fe4cc8, 32'hc4508069, 32'h4339fab4},
  {32'hc3c0752c, 32'h433ff351, 32'hc50bb52e},
  {32'hc3fc3130, 32'hc3ad52be, 32'h44c958d7},
  {32'hc2a5253a, 32'h44e21b4a, 32'hc31df813},
  {32'hc49abb01, 32'hc300a47a, 32'hc38a9887},
  {32'hc3467f54, 32'h43ca5a38, 32'h452b5ab9},
  {32'h434f4c55, 32'hc2d05fad, 32'hc4b1a84c},
  {32'h440d7e11, 32'hc2ff64b5, 32'hc48b0bda},
  {32'hc34e4cdc, 32'hc4b585ed, 32'h43a46e61},
  {32'hc4d9ea2c, 32'h427253ed, 32'hc2e40353},
  {32'hc39c2381, 32'h43c23bc4, 32'h419f0d6c},
  {32'hc367f143, 32'h44755d57, 32'hc4b6ef55},
  {32'h44fab0ea, 32'h43aa3455, 32'h43dec848},
  {32'h4502ef6c, 32'hc301336c, 32'hc40ab275},
  {32'hc52eb5a7, 32'h42be76a3, 32'h442a70ee},
  {32'hc3af5668, 32'h4361f1e3, 32'hc211d0a1},
  {32'hc4fdf798, 32'hc43cfc4b, 32'h438dc569},
  {32'h454b2e45, 32'hc383c638, 32'h40d32b1a},
  {32'h447a403c, 32'hc3bf782b, 32'hc26fb338},
  {32'h44fac22e, 32'h449e1a08, 32'hc410f686},
  {32'hc5392c58, 32'hc3a828c4, 32'h43b9236a},
  {32'hc4a7f0d4, 32'h4257b7f4, 32'hc365f2a0},
  {32'h43a973d1, 32'h42e37132, 32'h435c3159},
  {32'h437ee5c8, 32'h451356b8, 32'hc4e3777f},
  {32'h44bbc72e, 32'hc18d93b4, 32'h445c1e60},
  {32'hc3e7da65, 32'hc2a5a5e4, 32'hc3fdb8bf},
  {32'h445ee72d, 32'h438c6e2e, 32'h43b9d70a},
  {32'hc4fcb636, 32'hc3a1e6f6, 32'hc380715d},
  {32'h44109cde, 32'h4381fa7e, 32'hc3836e8c},
  {32'hc4fac3e5, 32'hc31400bd, 32'hc4b07dda},
  {32'h431f8d0a, 32'h442484b5, 32'h45334916},
  {32'hc4a755c0, 32'h43a3c1d6, 32'h429369db},
  {32'hc3daf6e7, 32'hc4989b88, 32'h44e4e875},
  {32'hc32c0f56, 32'hc49b3fcd, 32'hc48b0cea},
  {32'hc41f3170, 32'h4299f130, 32'h4444ebcd},
  {32'hc2b4a47a, 32'hc3c16499, 32'hc51393d3},
  {32'h4445a990, 32'h43a1aec5, 32'h449093a9},
  {32'hc4e0d6f5, 32'hc2793f04, 32'hc2d7842c},
  {32'hc392ada4, 32'h44d068cc, 32'h44d1badf},
  {32'hc3891a6b, 32'h437c7bf1, 32'hc516255d},
  {32'h437e670d, 32'h44f7f9e8, 32'h4406660e},
  {32'hc5127509, 32'hc41ad89f, 32'hc3900cb9},
  {32'h44f83cad, 32'h44b2f6c5, 32'h42ec3625},
  {32'hc49613a8, 32'h409a2de5, 32'h43810520},
  {32'hc323a740, 32'h45817a2f, 32'hc3cbd3fd},
  {32'hc46707b5, 32'hc50fe5d6, 32'hbe949dc5},
  {32'hc4849434, 32'h43afe2b0, 32'hc3f7d0b0},
  {32'hc5287385, 32'h445e18b8, 32'h43a04702},
  {32'h44f8393a, 32'h42a3e069, 32'h42d0a0f3},
  {32'h4498cd7c, 32'h4477ff36, 32'hc4ab99d7},
  {32'hc412b569, 32'h4314eb60, 32'h43fa61a8},
  {32'hc40fcbf8, 32'hc2c0fbe0, 32'hc384165f},
  {32'hc3f323bf, 32'h43429217, 32'h43df772d},
  {32'hc3221749, 32'hc362fc45, 32'hc51296b9},
  {32'hc499ba5c, 32'hc2009e34, 32'h42638445},
  {32'h4494984d, 32'hc420a57e, 32'hc48a9d8a},
  {32'hc45cef6c, 32'h43df9a6e, 32'h447e3894},
  {32'hc4af6891, 32'hc3af572b, 32'hc3e356da},
  {32'h420df330, 32'h443b5bab, 32'h44ad8a77},
  {32'h43cba5d6, 32'h44c2ef32, 32'hc4cf640c},
  {32'h437d2d1d, 32'hc4583929, 32'h44a81b62},
  {32'h42d9b612, 32'hc4bc19e5, 32'hc3d52864},
  {32'hc2e68586, 32'h43c75d2f, 32'h453ace49},
  {32'hc2892da0, 32'h43025ae6, 32'hc39f2e77},
  {32'hc4a532a7, 32'hc3e0d146, 32'h442621d6},
  {32'h4413dfac, 32'hc20703a3, 32'hc42a896a},
  {32'hc52b9658, 32'hc38b41a4, 32'hc3f81e0b},
  {32'h43ffe462, 32'hc4bd303a, 32'h4147d054},
  {32'hc5658aaa, 32'h43aa3357, 32'h4301df47},
  {32'h4479a01c, 32'hc46d553c, 32'h42e719a3},
  {32'hc4bfa644, 32'h448f01fe, 32'hc42bd6a5},
  {32'h43c692a2, 32'hc579e74d, 32'h42d9ab47},
  {32'h451168fa, 32'hc35c195b, 32'hc3076769},
  {32'h4486bd22, 32'hc12f54c6, 32'h43b7102f},
  {32'hc562c284, 32'hc409881f, 32'hc409dbf9},
  {32'h45752d3e, 32'h41cdf2ba, 32'hc419fcad},
  {32'h44a5cca5, 32'hc32d1044, 32'h41a4eb87},
  {32'hc5284809, 32'hc33d9e4d, 32'hc3993b61},
  {32'h451b41c6, 32'hc350bce5, 32'h4376aef7},
  {32'hc2d12786, 32'h44a47e98, 32'h41fe9de2},
  {32'h433f5778, 32'hc4479f83, 32'h42cc2b98},
  {32'hc46e9fa3, 32'h4448cb95, 32'h42fbc72a},
  {32'h442f4c68, 32'hc1c40686, 32'h41f7f838},
  {32'hc4b93a14, 32'h44454a32, 32'hc3a5f436},
  {32'h445bb52b, 32'hc51995e9, 32'h3f67df00},
  {32'h44771428, 32'hc39ad13b, 32'hc364056d},
  {32'h440ee552, 32'h439c6c99, 32'h44b90492},
  {32'hc462907f, 32'hc2d47020, 32'hc35853f0},
  {32'h44a6f169, 32'hc36217b4, 32'h42c1da85},
  {32'hc50c5f9c, 32'hc36d6ad1, 32'h43bdd959},
  {32'h44264ace, 32'hc400144f, 32'hc3db3640},
  {32'h43cd2578, 32'h429d528a, 32'h44ddc87e},
  {32'hc4450ac9, 32'hc40c1ad1, 32'hc43ce1d5},
  {32'hc435331e, 32'h440257c8, 32'h45309c42},
  {32'h453646be, 32'h427cc58d, 32'hc29cbf1a},
  {32'hc3cc91a6, 32'h44a5e55b, 32'h448d6105},
  {32'h42af6420, 32'h44916a69, 32'hc49a26d9},
  {32'hc3745c11, 32'h4397d4bf, 32'h4435dacf},
  {32'h446f411a, 32'hc4ba634b, 32'hc415e06d},
  {32'hc46a3cf2, 32'h42f2db33, 32'h4388120e},
  {32'h441f484d, 32'hc4288f05, 32'hc4070979},
  {32'hc41707b7, 32'h450119ec, 32'h436c7fc3},
  {32'h44e2381b, 32'hc4a06ab5, 32'hc3d43fc9},
  {32'h43262720, 32'hc42d03ff, 32'hc3c4ba30},
  {32'hc4dd747c, 32'h42972db9, 32'h42d9a8f1},
  {32'hc447b53d, 32'h4440b7c8, 32'hc4529582},
  {32'hc1601400, 32'hc442aaa7, 32'hc3e934a9},
  {32'h443fa343, 32'h44b2ce8e, 32'h439fe871},
  {32'hc41bf963, 32'hc3a4fb78, 32'h437a7912},
  {32'h4510bfa8, 32'h44ad95d8, 32'h4258c314},
  {32'hc55a1a90, 32'hc3e8b8cc, 32'h438eaac9},
  {32'h4252c508, 32'h451535f3, 32'hc24231eb},
  {32'hc365c1b3, 32'hc31b1cb9, 32'h44e5d0b0},
  {32'h443102b0, 32'hc43fcdbd, 32'hc4bc93a9},
  {32'h44fa5ea7, 32'hc38c449b, 32'hc25c2312},
  {32'h45027934, 32'h43cf1cf7, 32'h4230a35e},
  {32'hc3255e77, 32'hc43ed85b, 32'hc4a91d8a},
  {32'hc44afa60, 32'h42cf096f, 32'h4438c277},
  {32'hc3b7c4d3, 32'hc31ac9dc, 32'hc54157a7},
  {32'h44893d47, 32'h43c41b32, 32'h4492da79},
  {32'hc45a1fe2, 32'hc41f218a, 32'hc2bf70b9},
  {32'h4341c7a8, 32'h4407ddbb, 32'h43996c50},
  {32'hc51a97ae, 32'hc3d4081f, 32'hc3cc679a},
  {32'h452a0116, 32'h4411a225, 32'hc3c5d07d},
  {32'hc448c15a, 32'hc4c48a4b, 32'hc31872d6},
  {32'h45083fdf, 32'hc2ee990f, 32'hc2c631b1},
  {32'hc483164e, 32'hc3dd15ec, 32'hc1ab1dc2},
  {32'hc36571d0, 32'h4481d971, 32'h44c0ac24},
  {32'hc4d4aa88, 32'h4381861b, 32'hc42f1acc},
  {32'h43cd6104, 32'hc3443169, 32'h4404895d},
  {32'hc36a79f8, 32'hc3f7ccec, 32'h4301dd38},
  {32'hc4f45388, 32'hc37c3618, 32'hc32c557a},
  {32'hc31d27a0, 32'h448c332b, 32'h43c7d7e1},
  {32'hc410aed4, 32'hc3d2f342, 32'h43ae6464},
  {32'h449c7347, 32'hc3490e38, 32'h42f88b3f},
  {32'hc4f01de6, 32'hc35fbefd, 32'hc199c548},
  {32'hc49d7ce8, 32'hc3be47a2, 32'h435772e0},
  {32'hc5016fde, 32'hc276d740, 32'hc30ee25e},
  {32'h44a54483, 32'h44670214, 32'h4468679b},
  {32'h44d46f31, 32'hc2980fe9, 32'h43c4d377},
  {32'h44036094, 32'h445f3ac2, 32'hc2e9502c},
  {32'hc407db60, 32'h438d27ba, 32'hc4768b91},
  {32'h44b82062, 32'h4364d111, 32'hc31cbe1e},
  {32'hc3708750, 32'hc3cc0b8a, 32'h44e29efc},
  {32'h43adf516, 32'h4530d17e, 32'hc43c0cf9},
  {32'hc4e0ed30, 32'h4195703c, 32'h43cafbde},
  {32'h448629f4, 32'h43f97ed8, 32'hc4ee5862},
  {32'hc35adeec, 32'hc4c264d5, 32'hc4ad1781},
  {32'h44e8dc52, 32'h43b63150, 32'hc41b5469},
  {32'hc46ae558, 32'hc341857e, 32'h449d9bb5},
  {32'h447af2b3, 32'h44446293, 32'hc4e73a61},
  {32'hc4fc7b89, 32'h4256b934, 32'h437afd77},
  {32'h433f71ae, 32'h439ca5fa, 32'hc517ab5b},
  {32'h43412a17, 32'hc44769c2, 32'h4487a180},
  {32'h42f79320, 32'hc2a6b66a, 32'hc437277e},
  {32'hc44d6a07, 32'h440bdef2, 32'h45064dc2},
  {32'h44c96ad8, 32'hc35e1a8d, 32'hc509db04},
  {32'h430b0920, 32'hc493dbd8, 32'hc3f0e656},
  {32'hc4e6d328, 32'h4491e197, 32'h43bd5bfe},
  {32'hc49ce60e, 32'h43d71c33, 32'hc3816d61},
  {32'hc506d0f1, 32'h44878c39, 32'hc3928d3b},
  {32'h45129289, 32'hc3388c50, 32'hc2fde0ec},
  {32'h44b2b586, 32'h437e136f, 32'hc2bce986},
  {32'h444f9590, 32'h43d53293, 32'h431c5676},
  {32'hc464fea8, 32'hc37c7b55, 32'h441adaf6},
  {32'h45509c0d, 32'h41a3a8e8, 32'h43b3739b},
  {32'hc3caf38e, 32'hc2c977f9, 32'hc4648047},
  {32'h445d6bab, 32'hc443aaf2, 32'h4391bb32},
  {32'hc48b05aa, 32'hc340e0c6, 32'h43156b4e},
  {32'h430c77a6, 32'h40034809, 32'h450d1c63},
  {32'h43a9d03e, 32'h4443a66d, 32'hc4269c6d},
  {32'hc3cb00d4, 32'hc444bdfd, 32'h43ee911a},
  {32'hc50e03d1, 32'hc1c3eed5, 32'hc390384e},
  {32'hc350a853, 32'hc25f9965, 32'h44dbee97},
  {32'hc42acb31, 32'hc3e051c3, 32'h425017df},
  {32'h44d6026e, 32'hc47709be, 32'h42b311a4},
  {32'hc464990a, 32'h45369816, 32'hc3df1004},
  {32'h4263c5b0, 32'hc2bf4874, 32'h43949fc1},
  {32'hc30a5203, 32'hc388137d, 32'hc531abc0},
  {32'h43a310a7, 32'hc5186489, 32'hc3888ccf},
  {32'h4292a8b9, 32'hc3131dea, 32'hc3bc24e8},
  {32'h4509fec4, 32'h43810605, 32'h4417bf86},
  {32'hc57f56ae, 32'h43275c06, 32'h4380c24b},
  {32'hc4acd970, 32'hc3154486, 32'h43bb4476},
  {32'hc4d54ecf, 32'hc3d5587d, 32'hc404cc5a},
  {32'h4515e24e, 32'hc2671e26, 32'hc33372b2},
  {32'h42bb8c10, 32'h42e6705b, 32'hc3b4588e},
  {32'h44fb45e7, 32'hc35c6637, 32'hc24781da},
  {32'h4288e7e0, 32'hc4b0159f, 32'h43cfe3fb},
  {32'hc39859d8, 32'h45233bb2, 32'hc14db2c7},
  {32'hc4c9cd9f, 32'h4290366c, 32'hc407316d},
  {32'hc4abbe32, 32'h445416a7, 32'hc4284e53},
  {32'h444174ce, 32'hc4a8bf0d, 32'h43686392},
  {32'h44beb065, 32'hc2c63147, 32'h446f5c06},
  {32'hc4f6a208, 32'h449fb1fa, 32'hc3d48fc1},
  {32'hc46ef9b1, 32'hc41461e1, 32'h445d8abf},
  {32'h4437bb05, 32'hc3c31b5b, 32'h43c88a9f},
  {32'hc3d0bda7, 32'h44b48e22, 32'hc3414a2e},
  {32'hc40ba034, 32'hc4bbd6e8, 32'h44443ff3},
  {32'hc3269d2c, 32'h44e59a1d, 32'h4362bc76},
  {32'h44d189e6, 32'hc42705b2, 32'h4302782d},
  {32'hc53441da, 32'h41655006, 32'h43554c6d},
  {32'hc4869bb4, 32'hc3304a82, 32'h434dd799},
  {32'hc5381124, 32'hc2be27c5, 32'h4326de25},
  {32'h43a602d0, 32'h4473db04, 32'h447d6db9},
  {32'hc3f8f015, 32'h4468942f, 32'hc2527a15},
  {32'h456a8cd0, 32'hc409910b, 32'h43c47c73},
  {32'hc3c312f6, 32'h450f6470, 32'hc3420c78},
  {32'h451ee47e, 32'h440350c4, 32'hc360ba33},
  {32'hc5047390, 32'h449a1a36, 32'h4380d1f6},
  {32'h44bbe271, 32'hc4c1a14c, 32'hc38a30ef},
  {32'h42b43c58, 32'h4314e2fe, 32'h44743119},
  {32'hc3ba046c, 32'h444ab411, 32'hc51b7f32},
  {32'hc38d951e, 32'hc4c7b0aa, 32'h44fc7868},
  {32'hc4a75fd3, 32'hc44e83e8, 32'hc32fab95},
  {32'hc3b8a9a7, 32'h4246ae82, 32'hc5591b06},
  {32'hc421772e, 32'hc4632d02, 32'hc166c216},
  {32'h43b2b838, 32'h44fb571e, 32'hc3f327f9},
  {32'hc57b2a52, 32'hc3a16dab, 32'h4386888e},
  {32'hc4b13cc0, 32'h43fa8641, 32'h414abdb6},
  {32'h434103b3, 32'hc491f1be, 32'hc3e8d8c0},
  {32'hc5000f8d, 32'hc45fffb1, 32'h44e2ac0c},
  {32'hc3fe0672, 32'hc4920d02, 32'hc51f52be},
  {32'h442fb18e, 32'h44f13dd3, 32'hc3d109ca},
  {32'hc473b71c, 32'hc51926a4, 32'hc324cb37},
  {32'hc20aee00, 32'h439bc474, 32'hc3ecb104},
  {32'hc44fe209, 32'hc4852939, 32'h4352d92f},
  {32'h452995e1, 32'h43329d87, 32'hc38fe10e},
  {32'h434407c4, 32'hc3b9edbe, 32'hc26ef33f},
  {32'h45492460, 32'hc375c3ac, 32'h433b2200},
  {32'hc5136228, 32'h43c74771, 32'hc4075e56},
  {32'h43ecb09a, 32'h438f16aa, 32'hc391d750},
  {32'hc4e796e8, 32'hc44b7dfd, 32'h43e0f4c1},
  {32'h44118328, 32'hc21f5839, 32'h41d1328a},
  {32'h43d9f70e, 32'hc2361a33, 32'hc32b8648},
  {32'hc310cd36, 32'h454e8f49, 32'hc340770a},
  {32'hc3ed137c, 32'hc5367b59, 32'h4310403b},
  {32'hc1b5ed60, 32'h43770907, 32'h42d387ff},
  {32'h4411ce76, 32'hc3c51612, 32'h44ad6839},
  {32'hc43a9e10, 32'h440cce64, 32'hc48f811e},
  {32'h4364a1f1, 32'hc4e5c19b, 32'h44a47045},
  {32'h44d4899c, 32'hc3d73b40, 32'hc27b3157},
  {32'h43c55013, 32'h44145a35, 32'h44916a43},
  {32'hc42004c3, 32'hc46f1b01, 32'hc46233de},
  {32'h4467d9b8, 32'h4460db95, 32'h429faacb},
  {32'hc509a0b3, 32'hc31930e2, 32'hc40a096a},
  {32'h43c2510c, 32'h44760abf, 32'h4539fd53},
  {32'h449b78d3, 32'h41b6b792, 32'hc3a98555},
  {32'hc3b382a4, 32'h44a1b09c, 32'h4405da2e},
  {32'h43974b75, 32'hc4b81c19, 32'hc370ada3},
  {32'hc4158d8f, 32'h446eba4a, 32'h41e85657},
  {32'hc49a1b51, 32'hc3fd9bc5, 32'hc3351219},
  {32'h43e13ea7, 32'h453f293e, 32'h43de5770},
  {32'hc2a583b8, 32'hc3f54d86, 32'h439a58d7},
  {32'h44bbdeec, 32'h4281b576, 32'h440bd4d0},
  {32'hc46c14fe, 32'hc213db88, 32'hc42e6322},
  {32'h43e77444, 32'h43232794, 32'hc0a1f1cf},
  {32'hc4f28313, 32'hc481cee5, 32'hc387dafe},
  {32'h45619e5d, 32'h420f09d6, 32'hc3e90918},
  {32'hc51df3c0, 32'h44511b56, 32'hbeb02375},
  {32'h42232fa8, 32'h45236cf5, 32'hc3553352},
  {32'hc3d7b4ec, 32'hc53095c1, 32'hc28efde8},
  {32'h45500b2a, 32'h43f5c91e, 32'hc2f8f616},
  {32'hc596fceb, 32'h42821705, 32'hc37b92ad},
  {32'h454a8c7c, 32'hc34ffc3d, 32'hc34d5e85},
  {32'h43054853, 32'hc5074e08, 32'hc2a1b923},
  {32'hc25eaf64, 32'hc4eb4952, 32'h439f6835},
  {32'h4319ed40, 32'hc4237561, 32'hc404d663},
  {32'hc299acea, 32'h455cca02, 32'hc30a7440},
  {32'h443e0bf2, 32'hc48e9716, 32'hc339b4ba},
  {32'hc416315f, 32'h43c4cbfe, 32'h4461e237},
  {32'h438961b6, 32'hc482f6ba, 32'hc49223e8},
  {32'hc4addbbb, 32'h43f6f126, 32'h44b567ab},
  {32'hc31202c2, 32'hc440cb2c, 32'hc5012f2a},
  {32'hc3c40b33, 32'h44bd0d94, 32'hc38d096d},
  {32'hc446ae28, 32'h444cfed9, 32'hc4e4023c},
  {32'h4409e038, 32'hc3e1032f, 32'h440bdac3},
  {32'h440773ac, 32'hc45a4e6f, 32'hc4460112},
  {32'hc52b8f06, 32'h431abf94, 32'h432400fb},
  {32'h449a7d52, 32'hc33044f5, 32'h42dbcc42},
  {32'h4481c52a, 32'h44bff74e, 32'h4512459a},
  {32'hc334b0eb, 32'hc3c9637f, 32'hc5560469},
  {32'hc3396652, 32'h443228a8, 32'h42bbb4f4},
  {32'h4569f601, 32'hc412b9be, 32'hc22f05d2},
  {32'hc4668980, 32'h44a7d6f9, 32'hc12dd7dc},
  {32'h4419c5b1, 32'hc46167d0, 32'h427db136},
  {32'hc195c900, 32'h448bbea8, 32'h43ecbe6d},
  {32'h424ae8e0, 32'hc4d466b5, 32'hc1e9cd6f},
  {32'h449afc4e, 32'h431372f3, 32'hc38e8734},
  {32'h453eff4e, 32'h431f2c41, 32'hc3d44092},
  {32'hc4b5ce3f, 32'h4356baea, 32'hc1e27b17},
  {32'h44f73e20, 32'hc3cbb226, 32'hc39be0f1},
  {32'hc479a3fc, 32'h42928082, 32'h442973a4},
  {32'hc39ae43c, 32'hc4237074, 32'hc5518bf7},
  {32'hc30f1374, 32'h4434f31b, 32'h43b45ec8},
  {32'h4469e378, 32'hc3009d6a, 32'hc2d14c87},
  {32'h44512cf4, 32'hc404a814, 32'h4327500b},
  {32'h420f7500, 32'h452377f7, 32'hc11c20f4},
  {32'h45372de0, 32'hc20be733, 32'hc31b6e6c},
  {32'hc36ef9a6, 32'h450d0fe6, 32'h439509c0},
  {32'h4456eace, 32'hc48f4412, 32'hc39ce2ee},
  {32'h4479402a, 32'h43adb0f6, 32'hc4601884},
  {32'h43adf724, 32'hc2d65590, 32'hc4517031},
  {32'hc41dfd6a, 32'h43858bf7, 32'hc43a177f},
  {32'hc47d9439, 32'hc417aa58, 32'hc36fa726},
  {32'hc4ebec73, 32'hc35198a8, 32'hc28c8b9a},
  {32'h43a63c94, 32'hc4e158e5, 32'hc3c76ddb},
  {32'h442bd534, 32'h43be16e1, 32'h4358a49f},
  {32'h438f5000, 32'h4398caa5, 32'h41c7ebd4},
  {32'h426e8200, 32'h446ae370, 32'h4487f862},
  {32'hc2509a80, 32'hc41e13a9, 32'hc2ca823e},
  {32'hc3a2ba5d, 32'h4359fd69, 32'h446e7e2c},
  {32'h44a9a29a, 32'hc336a4c3, 32'hc4678653},
  {32'hc4832aa5, 32'h431b4c2d, 32'h43831f53},
  {32'h437d14da, 32'hc4645915, 32'hc50d6367},
  {32'h43630229, 32'h45435daf, 32'hc25c8c7f},
  {32'hc119c56c, 32'h43d5b9a0, 32'hc3d19020},
  {32'hc586b89e, 32'h43b80f18, 32'h43535f10},
  {32'h4500417a, 32'hc4670bd8, 32'hc43fefc6},
  {32'h43583856, 32'hc3434cc7, 32'hc56b880e},
  {32'hc413fcbc, 32'hc2f80f85, 32'h442c24cb},
  {32'h43f5e734, 32'h448eca5d, 32'hc4b17c54},
  {32'hc37047c8, 32'hc531e4ac, 32'hc36c1e98},
  {32'h455c9b4f, 32'h43230960, 32'h43af4c1f},
  {32'hc4cc3632, 32'h4360fe48, 32'h432d48fb},
  {32'h451ff01e, 32'h44405b4a, 32'h42637c7d},
  {32'hc51859cc, 32'hc42b7946, 32'h433bc7e6},
  {32'h4545d810, 32'hc2a4623a, 32'h44091789},
  {32'hc44c681a, 32'hc3869ed0, 32'h43dc77fb},
  {32'h43f6e250, 32'h43dfd20d, 32'h43d871ea},
  {32'hc41f20c3, 32'h438088e7, 32'h4396b10b},
  {32'h42b3bda0, 32'h448098cf, 32'h44c9e0d8},
  {32'hc423042a, 32'hc36e1f7e, 32'hc5594fe1},
  {32'hc3ad7d1d, 32'h442f0a02, 32'h42ddf7ad},
  {32'hc41ec4ea, 32'hc4c034cf, 32'hc2db4801},
  {32'h4402565e, 32'h4486f137, 32'h44331a0a},
  {32'h43c3e29d, 32'hc4951707, 32'hc35a09bf},
  {32'h44a227ca, 32'hc413f67b, 32'h44c018ef},
  {32'hc3dc9281, 32'hc3c3b987, 32'hc497bf79},
  {32'h452b88cd, 32'hc2ea1b95, 32'hc42f83ef},
  {32'hc314198a, 32'hc5285e79, 32'hc4849a4f},
  {32'hc202ab8e, 32'hc2bc6763, 32'h451acf6e},
  {32'hc30ab1ac, 32'hc4c2ee39, 32'hc338a102},
  {32'hc08cb9c0, 32'h44f4d220, 32'h4449be50},
  {32'hc471fb61, 32'hc3d8d0d3, 32'hc53d6aef},
  {32'h4476fba0, 32'h439156ab, 32'h435bc2de},
  {32'h4459cee2, 32'h431e0bb5, 32'hc2f39262},
  {32'hc4c15daf, 32'hc4523497, 32'h44119559},
  {32'h45098a4f, 32'h43e39c7b, 32'h3fb659f4},
  {32'h4499682c, 32'hc2c6eeda, 32'h434192c9},
  {32'h4452955b, 32'h44ec1d01, 32'hc23a3217},
  {32'hc4db1077, 32'hc2f23ec4, 32'h43631510},
  {32'hc435b903, 32'h442e4530, 32'h425a0eb4},
  {32'hc5694b7f, 32'h4140372a, 32'h433f2494},
  {32'h45117989, 32'hc2dbd795, 32'h432d4143},
  {32'h44d3b7f0, 32'hc3e6615d, 32'hc2014c73},
  {32'h43ff6828, 32'h44685f37, 32'hc4dd9a99},
  {32'hc4cdd119, 32'hc33f0bd7, 32'h43ad7226},
  {32'h43bdab4a, 32'h444b1a69, 32'hc3d31552},
  {32'hc4078680, 32'h42e687c7, 32'h44a1d632},
  {32'h4431fb00, 32'hc19d6b9c, 32'hc4e1da9f},
  {32'hc44287d9, 32'hc38ed52c, 32'h434a7743},
  {32'h44966a15, 32'hc38f70da, 32'hc46f7e1e},
  {32'hc4fcc756, 32'hc39ad41f, 32'h43c61f58},
  {32'h442c87c6, 32'h428e37d6, 32'hc4359259},
  {32'hc49caff0, 32'hc5086e0d, 32'hc34d9749},
  {32'h436ef3b8, 32'h4494ace1, 32'hc1afad4e},
  {32'h44ace9a6, 32'h431a7e33, 32'h43410d19},
  {32'hc34ce045, 32'h44261138, 32'hc4cf3e7b},
  {32'hc492cb26, 32'h42887522, 32'h449a07ae},
  {32'hc462e7b6, 32'h439c770f, 32'hc28f47ae},
  {32'hc53ed066, 32'hc337136c, 32'h4418a3b4},
  {32'h448c32a7, 32'h43ae3811, 32'hc4d963e5},
  {32'h44ac3f40, 32'hc4ae2f25, 32'h3fb21ffb},
  {32'hc541ae22, 32'h4412019d, 32'h42109242},
  {32'h447e18b6, 32'hc43c9b66, 32'h424bf9e8},
  {32'hc50f6bd3, 32'h4483fd68, 32'hc3c6def0},
  {32'h45484a86, 32'hc2d49eea, 32'h434fd51e},
  {32'hc3674709, 32'h446c3941, 32'h43a08804},
  {32'h445ecdd6, 32'hc35fdc46, 32'hc492f93e},
  {32'hc4d3cb21, 32'h42b07d57, 32'h42ad1603},
  {32'hc4c82b16, 32'h43511e85, 32'h43508ad6},
  {32'hc4310e8c, 32'h42db20b9, 32'hc49aa37d},
  {32'h4402cc89, 32'hc4495ca2, 32'h4333346a},
  {32'hc307606c, 32'h435d337a, 32'hc4b04ae0},
  {32'h431b27e5, 32'h4322a3cc, 32'h44895c44},
  {32'hc4bd47d1, 32'h4399cc7f, 32'hc46e886c},
  {32'h4378410f, 32'hc4a414f9, 32'h43522fc0},
  {32'hc495cb8c, 32'hc399b653, 32'hc4a43664},
  {32'h43e6a666, 32'h438deafb, 32'h44e4c79f},
  {32'h43247122, 32'hc3aaa776, 32'hc4b74ef5},
  {32'h4492135a, 32'hc4bc439e, 32'h44548193},
  {32'hc4fe6036, 32'h44388bf0, 32'hc48344bc},
  {32'h444c8f2b, 32'h43528370, 32'h4460bb9f},
  {32'hc535f0e2, 32'h4390ba97, 32'hc3029434},
  {32'hc2e03fdc, 32'hc5092932, 32'h4447d319},
  {32'h443d9a4e, 32'h432eeb7c, 32'h42cb5f9a},
  {32'h451ff7a2, 32'h400c71dc, 32'h442a64aa},
  {32'hc4121315, 32'h42a2daca, 32'hc4cc9096},
  {32'h4158dd00, 32'h42178150, 32'h4404149a},
  {32'hc49020ac, 32'hc34ccd83, 32'hc43dc7ca},
  {32'hc3febd01, 32'hc3ace395, 32'h44844ef4},
  {32'hc49a56da, 32'h4491477f, 32'hc4833310},
  {32'h44323c44, 32'h435ef560, 32'hc2e22f2f},
  {32'h44924095, 32'hc4ef7f65, 32'hc3ae183f},
  {32'hc39499a9, 32'h44c37aa8, 32'hc2ca8d70},
  {32'hc37ce62c, 32'hc352a4c5, 32'h4136f8f2},
  {32'h423ec080, 32'h4406e0cb, 32'hc42874d2},
  {32'h4400a54c, 32'hc41865a8, 32'h450fae90},
  {32'h43f00b50, 32'h437795e0, 32'h44ab5064},
  {32'hc4ca230f, 32'h44184b61, 32'hc4a00a87},
  {32'h42b9036b, 32'hc44d49ba, 32'h446241b2},
  {32'hc4ac35e0, 32'hc3f948d9, 32'h43487a24},
  {32'hc39f068a, 32'h4392d2d8, 32'hc4369c6e},
  {32'h44c09fd6, 32'hc47ffa87, 32'hc3a1e764},
  {32'hc400bd5d, 32'h43229b1e, 32'hc46c4bb5},
  {32'hc21a66e2, 32'hc4d558c5, 32'hc360fa27},
  {32'hc4ecfc5b, 32'h43ae559b, 32'hc40fd6b0},
  {32'hc4cfaa3d, 32'h3d8a2a00, 32'h43645edb},
  {32'hc5231b32, 32'hc4184be4, 32'hc422bc0f},
  {32'h451c932a, 32'h4379a0f7, 32'h4401562b},
  {32'hc49b3823, 32'h42e99f66, 32'h439a947a},
  {32'h43855a67, 32'hc54b8051, 32'hc363f8bb},
  {32'hc42424d7, 32'h44df85bd, 32'hc2a9e2a0},
  {32'h42091c13, 32'hc4c45724, 32'hc3f4a6a0},
  {32'hc5913ae1, 32'h4219a1af, 32'hc34b5a38},
  {32'hc38bd471, 32'hc50bb13b, 32'hc387f36a},
  {32'h4405488e, 32'hc449a5f4, 32'h44896260},
  {32'h44b87e6d, 32'h422c1575, 32'hc3f80ac2},
  {32'h4286032e, 32'h44bb4066, 32'h4498ef8b},
  {32'hc393cc84, 32'hc5073bfb, 32'h4412a5a0},
  {32'h440635ee, 32'h44828787, 32'hc478ee2a},
  {32'hc4e9c9f1, 32'h438b7eed, 32'h43189e43},
  {32'h43760c6e, 32'h449f2fe5, 32'hc4bd57e9},
  {32'hc4ca9c0a, 32'hc34f8dea, 32'h42f1de88},
  {32'h433b7b38, 32'h44781a15, 32'h4298be4f},
  {32'h42894017, 32'hc32e17e3, 32'hc3e47f43},
  {32'hc32ead78, 32'hc4875180, 32'h44b9bb63},
  {32'h44cddc98, 32'hc388a919, 32'hc451b7a2},
  {32'hc0d0b4f0, 32'hc3893279, 32'h42ce4939},
  {32'hc407ad92, 32'hc41d10ca, 32'h44322a9b},
  {32'h438ec2a0, 32'h427d1a8f, 32'hc4139bdd},
  {32'hc40531ec, 32'hc4f9a54c, 32'h4331096a},
  {32'hc29a0963, 32'h452d2d50, 32'hc325ed76},
  {32'h439eecdf, 32'h429008f1, 32'h450072e0},
  {32'h44157fbf, 32'hc3d83d02, 32'hc3ffa623},
  {32'hc4818e46, 32'h43b60c4f, 32'h428e30b0},
  {32'h454e4722, 32'hc2a1e446, 32'h421847b6},
  {32'hc488765b, 32'hc3a027b1, 32'h445452cb},
  {32'h43928591, 32'h4561dfc3, 32'hc2da093d},
  {32'hc417883b, 32'h42c45785, 32'hc301627a},
  {32'h44b9ad76, 32'h44a6748a, 32'hc35bc659},
  {32'h42b89428, 32'hc53b9bc7, 32'h4348c5be},
  {32'hc4d05e62, 32'hc331d6d0, 32'hc3d0849c},
  {32'h4487b3b7, 32'hc4478c39, 32'hc0e48660},
  {32'hc33c0050, 32'hc4679f9f, 32'hc3ce4fd0},
  {32'h41fdeb94, 32'h42af4d6b, 32'h4421f5e0},
  {32'h442ad777, 32'hc4119182, 32'hc44ce64b},
  {32'h44b1cc86, 32'h44578369, 32'h44865d64},
  {32'h40048980, 32'hc4f3420d, 32'hc360026a},
  {32'h44085e41, 32'h430d20d3, 32'h44fcca6d},
  {32'hc35ebab4, 32'hc41011ab, 32'hc51c4bd0},
  {32'h426a96a8, 32'h4402eeff, 32'h45649bf7},
  {32'h4305050f, 32'h43cca0b2, 32'hc3e83ec7},
  {32'hc3fee022, 32'hc529b0ba, 32'h44b13713},
  {32'hc3cc108a, 32'h43ab3791, 32'hc407e456},
  {32'hc4a57be8, 32'h42ca05d5, 32'hc292cd00},
  {32'hc2d301ac, 32'hc10f2dd6, 32'hc4e087e1},
  {32'h44a59e9e, 32'h444fe5c9, 32'h4371d89e},
  {32'h4435e246, 32'hc496e521, 32'hc410a5dd},
  {32'h4319d482, 32'h44af0450, 32'h44d76f60},
  {32'hc46b95e6, 32'h434d66f8, 32'hc39f3707},
  {32'h45191228, 32'h42a8a874, 32'h430c6270},
  {32'hc4800d39, 32'hc4a5c5e5, 32'hc3bcae2e},
  {32'h44757d52, 32'h45205dd4, 32'h41d31146},
  {32'hc50fd6fb, 32'h4411366f, 32'h41e43453},
  {32'h43ea48d0, 32'h450ecc2a, 32'hc30e2435},
  {32'hc431af28, 32'hc4c7eb66, 32'h415dfd86},
  {32'h45504aec, 32'h4332a32c, 32'h416f884c},
  {32'hc513a7ff, 32'h444e4c56, 32'h42e1e6c0},
  {32'h4509e4c3, 32'hc39dc7d0, 32'hc118f438},
  {32'h432780b0, 32'hc567c674, 32'hc3b889cd},
  {32'h40bafd0a, 32'h449cda02, 32'hc250bd7a},
  {32'hc07e4f40, 32'hc36f2f2f, 32'hc3d85b23},
  {32'hc4e3514a, 32'h42058adb, 32'h440a90bb},
  {32'h43a80c9c, 32'hc51c5cb7, 32'hc199bcf1},
  {32'hc4ecea10, 32'hc4007124, 32'h4407c1d4},
  {32'h451598b0, 32'h43800b2c, 32'hc3ec3f76},
  {32'hc3afc2b6, 32'h441e2574, 32'h454e9aee},
  {32'h4474049c, 32'hc3a596e6, 32'h43d33815},
  {32'hc41233e6, 32'hc3d206d0, 32'h44857f4b},
  {32'hc3283f80, 32'h452c448b, 32'hc4e22dc5},
  {32'hc2e150f0, 32'h3fc0f780, 32'hbdb96400},
  {32'h4236cf20, 32'hc40ef9f6, 32'hc40aaa58},
  {32'hc4b083ac, 32'h4351ff1e, 32'h44205995},
  {32'h440dc313, 32'hc22440cd, 32'hc4e44749},
  {32'h44243180, 32'h44b71af5, 32'h452a27f6},
  {32'h44b38a5d, 32'hc3b9deda, 32'hc482ca96},
  {32'hc42997e5, 32'hc2d51d15, 32'hc40238a8},
  {32'h45081c0c, 32'hc423cd20, 32'hc40d48bd},
  {32'hc4b58ddf, 32'h43f6be19, 32'hc291fb55},
  {32'h42fc5cdc, 32'hc3d4717a, 32'hc25802dc},
  {32'hc5237d68, 32'h448c419c, 32'hc3976e04},
  {32'h434d9996, 32'hc56ee232, 32'hc3a43140},
  {32'h4409e357, 32'h440b3692, 32'hc1d65685},
  {32'h457718f6, 32'h43ef3991, 32'h439956a8},
  {32'hc4c2af8c, 32'h43b8cb68, 32'h4430e3a4},
  {32'h45426039, 32'h43fb987c, 32'hc3868d1c},
  {32'h452c0a0f, 32'hc2cd3344, 32'hc3b70f3a},
  {32'hc4c71752, 32'hc0aba6a0, 32'hc4f73e6f},
  {32'h441fb890, 32'hc31a7ae0, 32'h455da848},
  {32'h449d41e5, 32'h4478ea09, 32'hc1ba570e},
  {32'h4378f0a6, 32'hc55882aa, 32'hc3486ea3},
  {32'hc39040d0, 32'h44b2841d, 32'h44199c5f},
  {32'h45636bd1, 32'h441bbafa, 32'hc3bc4dee},
  {32'hc3db5e26, 32'h4474fcae, 32'hc3a82c77},
  {32'h44615222, 32'hc47ea8cf, 32'hc344c886},
  {32'hc4b1f55f, 32'hc39ecb08, 32'hc28a3866},
  {32'h445366a4, 32'h43682266, 32'h442f867e},
  {32'hc4ce5045, 32'hc3019efb, 32'h4277040c},
  {32'h4456a89e, 32'hc3a21d45, 32'hc3b85bea},
  {32'hc2c95014, 32'h43869350, 32'h44e64ae7},
  {32'hc396b563, 32'hc4839624, 32'hc5040f5c},
  {32'h43efd3de, 32'h43e53617, 32'h4390aa11},
  {32'h443c1a2a, 32'hc380934a, 32'hc37866a9},
  {32'hc336d4b0, 32'h44a834e5, 32'h4443f7ae},
  {32'h453ee4d5, 32'hc11b1ed1, 32'hc3853a61},
  {32'hc43a3cd5, 32'h4440f827, 32'h44cfa7d9},
  {32'h4489f863, 32'hc2d6a0b5, 32'hc49f2fe1},
  {32'hc3ff6864, 32'h44b214dc, 32'hc3596d96},
  {32'h444fa46c, 32'hc4a9c257, 32'hc3b8d890},
  {32'hc445f4f4, 32'h449a4b06, 32'h44094511},
  {32'h4378deba, 32'hc3744d68, 32'hc4d94915},
  {32'hc38d1e7a, 32'h4361071d, 32'h448305e8},
  {32'hc384d14c, 32'hc3b2e891, 32'hc56d5b1e},
  {32'h43138c3c, 32'h40ddd2fa, 32'hc53212bb},
  {32'hc4cc2850, 32'h435ada43, 32'h449f9dd7},
  {32'h4471f9a4, 32'hc288f11a, 32'hc4387f7c},
  {32'hc556001f, 32'hc3d15181, 32'h41edd384},
  {32'h4260bfae, 32'h452d324b, 32'h43568017},
  {32'hc3e4b594, 32'h420b79e2, 32'hc3476610},
  {32'h453d6a03, 32'h44828133, 32'h424067f0},
  {32'hc503da32, 32'hc49d9a01, 32'h440b640b},
  {32'h4433d334, 32'h44827a85, 32'h4281b2c6},
  {32'hc500ca29, 32'hc42d8064, 32'h43a057d7},
  {32'h44d61c3e, 32'hc328d7fc, 32'hc4cda3f5},
  {32'hc509f5d9, 32'h434d33f5, 32'h438c11e6},
  {32'h40bafb5b, 32'h43ca3d45, 32'h42d1076c},
  {32'hc4bc4729, 32'hc4c36bfd, 32'hc4415457},
  {32'h42e9e47c, 32'h430f2706, 32'h44ee9398},
  {32'hc4b11c80, 32'hc492c6e8, 32'h434f2670},
  {32'h443205fa, 32'h44581e20, 32'h4483f671},
  {32'hc4c3578a, 32'h422efd9c, 32'h442a1292},
  {32'h44ce1ce0, 32'h44a3453b, 32'h4419fe11},
  {32'hc535e332, 32'h434465b8, 32'hc4082da5},
  {32'h444b9523, 32'h41f49cbd, 32'hc13e371b},
  {32'hc4c633ee, 32'hc23374d3, 32'hc44039aa},
  {32'hc32811a1, 32'h44a31d21, 32'h4499693b},
  {32'h45049551, 32'h422fa618, 32'hc2c2958b},
  {32'h440eca10, 32'h447d9d55, 32'h43a81acd},
  {32'hc45864f3, 32'hc4af6a57, 32'hc42cd573},
  {32'h4485ad10, 32'h448715a5, 32'hc3865dbe},
  {32'h43c33d47, 32'h447bd5eb, 32'h4156f872},
  {32'hc3b35eee, 32'hc477fbd8, 32'hc38a580f},
  {32'h438eea95, 32'h4525d0a6, 32'hc2a138a4},
  {32'hc400e914, 32'hc4735ac1, 32'h43cbf181},
  {32'h4507dbc4, 32'h443c9c62, 32'hc3beecb5},
  {32'hc497889a, 32'hc4f64fce, 32'h428113ff},
  {32'h451ed649, 32'h4394c2aa, 32'hc389ffa0},
  {32'hc55b8bd5, 32'hc2f2daa4, 32'h434d468d},
  {32'h43cd4d5c, 32'h4442cd93, 32'h4475ef35},
  {32'hc44bccfe, 32'hc4282a36, 32'hc275a4af},
  {32'h44cfc156, 32'h42c1f72e, 32'hc2bd37a8},
  {32'hc31cb1d0, 32'hc4db57d4, 32'hc2d64e00},
  {32'hc2c73f50, 32'h43f02e57, 32'h42880e36},
  {32'hc39120da, 32'hc48c93e2, 32'h441d99eb},
  {32'h42b3a170, 32'h4505eeaf, 32'hc437c2f5},
  {32'hc3da02d1, 32'h418bc42e, 32'h45013d0f},
  {32'h44ab5bf1, 32'hc33cfa56, 32'hc4779355},
  {32'hc43616be, 32'h439006b4, 32'h44fa16c3},
  {32'h43a2f011, 32'h44a1eb77, 32'hc3959a45},
  {32'hc576ce86, 32'hc32771e9, 32'h4380887b},
  {32'h43a5a393, 32'h45533461, 32'hc21f431d},
  {32'h43a1d198, 32'hc3433c40, 32'h444b0eba},
  {32'h427e3ee0, 32'hc38663b0, 32'hc4cb9de4},
  {32'hc3540f04, 32'hc43e3855, 32'h4432ce1d},
  {32'h44c4f10a, 32'h438ddb57, 32'h4301d309},
  {32'hc473b448, 32'h43e19835, 32'h44c756a2},
  {32'h43153d14, 32'h41885b84, 32'hc4ca4a52},
  {32'h4461c9d6, 32'hc4d77851, 32'hc3f8f2a3},
  {32'hc5242d9f, 32'h4204d243, 32'h43e66cb3},
  {32'hc3a59d73, 32'hc2eb95d7, 32'h42247bb6},
  {32'hc4e608a5, 32'h4452b806, 32'hc3c2e4dd},
  {32'h45488cce, 32'h4333b337, 32'hc333ca1e},
  {32'h44c83c56, 32'h430f569f, 32'hc39cf4d9},
  {32'h44a6ce72, 32'hc3ee3de9, 32'hc40fc804},
  {32'hc3b23734, 32'h44916fc8, 32'h44754c62},
  {32'h453b3a74, 32'hc39bf6b8, 32'h43bb628b},
  {32'h433163a4, 32'h4495f0db, 32'hc421f953},
  {32'h4487ce59, 32'hc4648f00, 32'h44ad11fd},
  {32'h44b0b6eb, 32'hc2ddc90b, 32'h425c0cc7},
  {32'h45173054, 32'h4405e4df, 32'h4400364d},
  {32'hc41f32da, 32'h44a59653, 32'hc32b876c},
  {32'h4248ad34, 32'h43517bd2, 32'h4498b4e5},
  {32'h42f3e2ce, 32'hc317df14, 32'hc4d3dae8},
  {32'h431104c0, 32'hc23b5af0, 32'h447363a2},
  {32'h44ef21a3, 32'hc3565b26, 32'h431dd956},
  {32'h44f256c9, 32'hc3d7313a, 32'h44b51451},
  {32'hc4959010, 32'h44426877, 32'hc49cdc53},
  {32'h44b49828, 32'h421a1f27, 32'hc389d7eb},
  {32'hc421a6b3, 32'h44a1cce1, 32'hc468b083},
  {32'h44a1c4e8, 32'h43438d4b, 32'h43beb424},
  {32'hc202d700, 32'h4464a04e, 32'hc49a0a70},
  {32'h44c131d7, 32'h43ed6235, 32'h43408e3f},
  {32'hc4aa6c05, 32'hc4689dfa, 32'hc4c57a63},
  {32'h45545254, 32'hc3e05825, 32'hc470d5ee},
  {32'h436b71a8, 32'hc469e397, 32'hc4be19f0},
  {32'h4443cf78, 32'hc4689ea1, 32'h44a23cf8},
  {32'hc52a2cee, 32'h439a14bd, 32'h430bcc91},
  {32'hc326f366, 32'h44131b7a, 32'hc43eded6},
  {32'h44639b89, 32'hc344a14d, 32'h44f11483},
  {32'hc3ad0de1, 32'hc38503ab, 32'hc4d0f364},
  {32'hc2f9a31f, 32'hc44dfeaa, 32'h444789dc},
  {32'hc490e38b, 32'hc302590c, 32'hc5251667},
  {32'h433134bb, 32'hc2ed42f0, 32'h44de07db},
  {32'h452fceb0, 32'hc3eb6b09, 32'h43e73bff},
  {32'hc4a0400e, 32'hc4f66524, 32'hc4364e3a},
  {32'h444b2661, 32'h43930540, 32'h43fd40fe},
  {32'h44dfd157, 32'h428fb678, 32'hc320f2d8},
  {32'hc4a5e9ec, 32'h43323b71, 32'hc442552e},
  {32'h4466ede8, 32'hc3a05c15, 32'hc3bc8bef},
  {32'h42e83e58, 32'h44f4bd38, 32'h42898e14},
  {32'h44c2d752, 32'hc2809dd7, 32'hc3397af7},
  {32'hc21c7205, 32'hc3bcc644, 32'hc562eb66},
  {32'hc4fddb3f, 32'hc2dafa57, 32'hc2933018},
  {32'hc5028159, 32'hc425f528, 32'hc22cb829},
  {32'h4523fcac, 32'h441a9965, 32'h43c5be44},
  {32'hc556f87c, 32'hc40dcf08, 32'hc289451b},
  {32'h44a82999, 32'hc4b9dc58, 32'h4428b804},
  {32'hc15f3c50, 32'h44f370c9, 32'hc36d60d3},
  {32'hc431a58e, 32'hc3043749, 32'h42a78a4d},
  {32'hc555c780, 32'hc340f6b1, 32'hc3ece72e},
  {32'h4465818b, 32'hc4c0ce09, 32'h42a41e95},
  {32'hc4266da6, 32'h4222fdc2, 32'hc30e54b4},
  {32'hc36c7b00, 32'h43dc6ea5, 32'hc55881aa},
  {32'hc382b736, 32'hc3bb3a55, 32'h452d2070},
  {32'h42c0fc48, 32'hc2fb98a9, 32'h4482079e},
  {32'h43e080da, 32'h449a828a, 32'hc36606bf},
  {32'h43d874b0, 32'hc49e7822, 32'hc0e8585a},
  {32'h43afb13e, 32'h44144b4e, 32'hc53d35bb},
  {32'hc5183faa, 32'hc39e929e, 32'h43c0a9f2},
  {32'hc3d699fc, 32'h44a12880, 32'hc2fff5bf},
  {32'h443d4447, 32'h440c9497, 32'hc0db8f77},
  {32'hc23f6e93, 32'h44dce210, 32'h44d96bb1},
  {32'h449c41ec, 32'hc2d4eec4, 32'hc3ea106d},
  {32'h44488b56, 32'h44d01fd7, 32'hc3afc2d9},
  {32'hc5467893, 32'hc341eded, 32'h42840476},
  {32'hc46dd90d, 32'hc08be392, 32'hc450fc79},
  {32'hc4b5ef9c, 32'hc403c0d0, 32'h444f9e75},
  {32'h44597a53, 32'h43a9a086, 32'hc41d3c7b},
  {32'h42a05a26, 32'hc2661946, 32'h44fc3e4b},
  {32'h4560c438, 32'h416c55a0, 32'h4434fdca},
  {32'hc544f2d0, 32'h42e73f42, 32'h42a474f5},
  {32'h45292f0c, 32'h435f95b2, 32'hc30c898a},
  {32'hc30a706a, 32'hc509d552, 32'hc3838d8b},
  {32'h451b2ee7, 32'hc0609b40, 32'h4323b05c},
  {32'h4404188a, 32'hc468fc20, 32'hc38b4944},
  {32'h431f6e60, 32'h4553687a, 32'h4244c0e5},
  {32'hc51d1c4a, 32'hc42f2f8e, 32'hc354193a},
  {32'h45169203, 32'hc2f694d2, 32'hc33e6a98},
  {32'hc3d1e8c3, 32'hc31eb745, 32'h43ecb361},
  {32'h43e92468, 32'h43814813, 32'hc42362a0},
  {32'hc1b4c800, 32'h4477ceda, 32'h447ba9d9},
  {32'hc42d4b6b, 32'h432b3098, 32'hc2c2de70},
  {32'h447df52e, 32'h444ad103, 32'h43b23cf6},
  {32'hc3a22ccc, 32'h435da593, 32'hc4c27cc8},
  {32'h444b2554, 32'h44828d85, 32'h42d44354},
  {32'hc51d2626, 32'hc4169c48, 32'hc447ba40},
  {32'h447dfdfb, 32'h443d58dd, 32'h448f6ba5},
  {32'h43c2337f, 32'h446662df, 32'hc45de488},
  {32'hc39f1c6c, 32'h44a4f354, 32'h437bde9a},
  {32'hc4d3c3ec, 32'h4393883a, 32'hc2272c78},
  {32'hc351984c, 32'h4488a12c, 32'h41609efd},
  {32'h4188a000, 32'hc409ca40, 32'hc4f95d1e},
  {32'h448a086a, 32'h44bb5ed5, 32'hc39fa822},
  {32'hc50ef7bd, 32'hc3355c51, 32'h43a8b7ee},
  {32'h4440e35d, 32'h442130aa, 32'h45087020},
  {32'hc439f390, 32'h41f689fc, 32'hc4617051},
  {32'hc483fe4d, 32'h43ed492b, 32'h43557f68},
  {32'hc45575a4, 32'hc5255df4, 32'h4321c7d7},
  {32'h445866f2, 32'h448c2807, 32'h4227c869},
  {32'hc47bb48a, 32'h4381a8c5, 32'hc29f716f},
  {32'h448fad9d, 32'h44c4cf89, 32'h442a4064},
  {32'hc4d80f7c, 32'hc470608d, 32'h41338650},
  {32'hc3441ebc, 32'hc0c2c810, 32'hc1ddadf6},
  {32'hc4994d73, 32'hc3705cdc, 32'h4345bae1},
  {32'h445dacf6, 32'h423cebc6, 32'hc3de5d49},
  {32'h42f22596, 32'hc3a87dba, 32'hc4c8b5bb},
  {32'hc321058d, 32'h4482c8ed, 32'h4467f896},
  {32'h42854f98, 32'h4303d459, 32'h432e4ba7},
  {32'hc36faac6, 32'h439a4052, 32'h451d81e8},
  {32'h4138d420, 32'hc53b0eb4, 32'hc3c878f3},
  {32'h4482add6, 32'h43a35424, 32'h439aac24},
  {32'h450216ab, 32'hc3bd67b5, 32'h43281644},
  {32'hc30c764c, 32'h44143cd4, 32'h452a5616},
  {32'h450f1ccf, 32'hc00c9f20, 32'h43a93afa},
  {32'h43ec3f85, 32'hc4a3529f, 32'h44fc3b52},
  {32'hc363c2a4, 32'hc4d2b366, 32'hc45f4aa8},
  {32'hc481b1ee, 32'h43fb4178, 32'hc28d82a0},
  {32'h42b535e9, 32'hc4d4446f, 32'h412f4d3f},
  {32'hc4956b87, 32'h442bc704, 32'h4429113d},
  {32'hc3cf184e, 32'hc412f15e, 32'hc3026990},
  {32'hc4e99044, 32'h42e76ef8, 32'h43ccb6c4},
  {32'h4344e3c6, 32'hc468bdd2, 32'hc4d1712d},
  {32'h448a7323, 32'h43b06bc6, 32'h43b781b8},
  {32'h4469dd74, 32'hc4e8f80e, 32'hc3de922d},
  {32'hc44fd7c0, 32'h45464076, 32'h43bfb4ae},
  {32'hc496c4bd, 32'hc42c7fbb, 32'h4393912c},
  {32'hc34d8883, 32'h451a4eeb, 32'hc2edac3d},
  {32'h44ea35f8, 32'hc463c763, 32'h43d02893},
  {32'hc41b3028, 32'hc2fda5b8, 32'h4399f09a},
  {32'h454bddb1, 32'h430fcf9d, 32'hc20726dc},
  {32'hc51d17ea, 32'hc42b0445, 32'hc23deecc},
  {32'h4552b189, 32'h43bc5036, 32'hc3e2dd93},
  {32'h454d571e, 32'hc3087f4c, 32'hc414d1d5},
  {32'hc409f83c, 32'h42329cfd, 32'hc457e29c},
  {32'h445cb7ed, 32'hc3b10673, 32'h44abb0f8},
  {32'hc421e802, 32'h44ac82ed, 32'hc2e2378d},
  {32'h42b30900, 32'hc2da3f0f, 32'h440f5152},
  {32'h438f143f, 32'h453e085f, 32'h43bb1d89},
  {32'h40198ca0, 32'hc47a0c79, 32'h4324da49},
  {32'hc50f4a6a, 32'h4456b9e6, 32'h424bbdf0},
  {32'h43414aa3, 32'hc53d5684, 32'h43e0a556},
  {32'h44914d2e, 32'hc3464bac, 32'hc47a1fda},
  {32'h4296c338, 32'hc28ac478, 32'h44d87d60},
  {32'hc42a0a1b, 32'hc32d20c6, 32'hc48271a5},
  {32'h43753846, 32'hc419205a, 32'hc3987a68},
  {32'hc38fbdb0, 32'h433f392e, 32'h44103f00},
  {32'h438d10a0, 32'hc383b9d1, 32'hc48ec765},
  {32'hc3817a24, 32'h4385aff2, 32'h449539dc},
  {32'h44a0ebb0, 32'hc2e5bd5a, 32'hc4a95269},
  {32'hc400ad78, 32'h43a1f57d, 32'h44debc67},
  {32'h4520e7ec, 32'hc2560d57, 32'h44113a9b},
  {32'hc53cd8ac, 32'h43e683f0, 32'h43e8df8d},
  {32'h44eda475, 32'hc3e43c63, 32'hc4472d75},
  {32'h44f020ee, 32'hc309bd99, 32'h439d4ffe},
  {32'h4485ceee, 32'hc4a1bcf9, 32'hc459860d},
  {32'hc46da55a, 32'h448cad35, 32'h44c105b5},
  {32'hc438936a, 32'hc3803144, 32'hc447c203},
  {32'hc4e05c1a, 32'h43de4bd5, 32'h448c2233},
  {32'h4229567d, 32'hc564dcbd, 32'hc2dba999},
  {32'h450c2172, 32'h4390d35d, 32'h415417c1},
  {32'hc527f73b, 32'hc24131cf, 32'h448b14a6},
  {32'h43dd8ca6, 32'h4485d320, 32'hc4971b5b},
  {32'hc20ac3b0, 32'hc54a0ef2, 32'h409fbd81},
  {32'h448fed9e, 32'h441d814d, 32'hc3828a52},
  {32'hc36a1d05, 32'hc4d95108, 32'h43326866},
  {32'hc3ac8c58, 32'h458250fe, 32'hc36f46ce},
  {32'hc4929e6c, 32'hc4a348b9, 32'h43a0aac7},
  {32'h44ef6aac, 32'h421c6cd8, 32'h43504e21},
  {32'hc476026c, 32'h4416428c, 32'hc447e662},
  {32'h441338cc, 32'h439ed278, 32'hc432e4b9},
  {32'h42505ae0, 32'hc3072520, 32'h4347ed5f},
  {32'h44b55c88, 32'h43ff4fbe, 32'h437855d0},
  {32'h4229b7b0, 32'hc469f307, 32'hc4bc5e14},
  {32'h44d38f9e, 32'hc395294d, 32'hc2ebe99f},
  {32'hc4b0cbcc, 32'hc3f78f4a, 32'hc4b7777b},
  {32'h43bdf070, 32'h4483b587, 32'h44e06e2d},
  {32'hc38a8624, 32'hc432768a, 32'hc32aa411},
  {32'h44c630ce, 32'h4368d4df, 32'h43da6f92},
  {32'hc44b8d21, 32'h41c127cb, 32'hc38fc217},
  {32'h45459f31, 32'hc39ee439, 32'hc3852810},
  {32'hc44facc1, 32'hc10f421b, 32'hc50445f7},
  {32'h43eaba8a, 32'h44f3add1, 32'h446b519b},
  {32'h434f4780, 32'hc3ae2310, 32'h43e874cd},
  {32'h42c39390, 32'h44bd3a20, 32'h443b18b4},
  {32'hc3f8e640, 32'hc1a88ffa, 32'hc5531cbe},
  {32'hc240c5c2, 32'h4448f266, 32'h442b64db},
  {32'h4431434b, 32'hc171011e, 32'hc3ace22a},
  {32'hc5788232, 32'hc2738554, 32'h4432fc4d},
  {32'h45034807, 32'h43f4db8d, 32'h42968498},
  {32'hc3becc0b, 32'hc3567271, 32'h43855aa2},
  {32'h4453779b, 32'h44b55702, 32'hc38f9731},
  {32'hc3be595e, 32'hc5140931, 32'hc322ac9d},
  {32'hc4117f55, 32'h429e57c5, 32'h43a5bff3},
  {32'hc560bd32, 32'hc329efed, 32'h4410cef8},
  {32'h441d7028, 32'h447fb349, 32'h4405672a},
  {32'h44e8d510, 32'h42b46ca2, 32'h4399d5d4},
  {32'h42d4e52b, 32'h453437a6, 32'h43296ee5},
  {32'hc3cbe828, 32'hc3c3c2d6, 32'h44ece828},
  {32'hc40d8844, 32'h44616082, 32'hc366cc00},
  {32'hc4ab06ae, 32'hc4604c41, 32'h428e1a02},
  {32'h4512845c, 32'h442971e9, 32'h429a85bf},
  {32'hc4e6f472, 32'hc2ff4e0d, 32'h429a5132},
  {32'h43a1f90f, 32'hc366a4b8, 32'hc4c314e0},
  {32'hc3fe003a, 32'h40c43ac7, 32'h44bbf028},
  {32'hc4e1d6c3, 32'hc290f1de, 32'hc2e69cbb},
  {32'hc41c0ced, 32'hc4c252ce, 32'h43829fcd},
  {32'h451c6e90, 32'h447b9dcc, 32'hc3a0899a},
  {32'hc51a5c41, 32'h43d72539, 32'hc30b94c4},
  {32'h43411650, 32'h44032ea4, 32'hc508c429},
  {32'hc38d4ce8, 32'hc5650316, 32'hc0ac771a},
  {32'hc4393a14, 32'hc31f6e83, 32'hc3ae88cc},
  {32'hc472727c, 32'h4391c0f2, 32'h44b7415e},
  {32'h442ea088, 32'hc33c27dc, 32'hc5186def},
  {32'h453a4d81, 32'hc44b714e, 32'hc31f87fa},
  {32'hc32df724, 32'h450045b8, 32'h433aaddc},
  {32'h4509bd98, 32'h42ffcaac, 32'h43fd18f9},
  {32'hc4ca7591, 32'h43df94a7, 32'h4444f30e},
  {32'h4504a106, 32'hc3d39853, 32'hc3bb46ee},
  {32'hc40e3ac3, 32'h4416dd67, 32'hc36320fc},
  {32'h4493e8de, 32'hc451111b, 32'hc4113bac},
  {32'hc5129c7f, 32'hc419db0b, 32'h42581043},
  {32'h44e09e94, 32'h43d6658d, 32'h441fca7c},
  {32'h441be58a, 32'h44cd5e66, 32'hc2ce0938},
  {32'h4468eb64, 32'h44357806, 32'hc438d00a},
  {32'h44b5055b, 32'hbfea0fa3, 32'h4403b0aa},
  {32'h4456dfde, 32'hc4b94689, 32'h441f6888},
  {32'hc43c4320, 32'h44cb811e, 32'hc43699ef},
  {32'hc463a5d6, 32'h43dd4846, 32'h442e886b},
  {32'hc17af900, 32'hc335b950, 32'hc50b9a3b},
  {32'h43fa384c, 32'hc4b0e306, 32'hc40e26f6},
  {32'h42fa12e8, 32'hc23686c5, 32'hc4a51631},
  {32'h43350e35, 32'hc4d5ab48, 32'h447d62c2},
  {32'h41a3de80, 32'h44e8deb1, 32'hc4528918},
  {32'hc3b85aa5, 32'hc3065e4c, 32'h446ea96e},
  {32'hc492a495, 32'h44a46711, 32'hc43c4c8a},
  {32'h44acad44, 32'hc39ef347, 32'h42c8964b},
  {32'hc3e968f8, 32'hc2dfbc9f, 32'hc33a668c},
  {32'h441128bf, 32'h441284e3, 32'h43979b0b},
  {32'hc5302425, 32'h437d74b9, 32'hc418a4d5},
  {32'h44fb2b5a, 32'h4392ca8c, 32'hc34dc9c0},
  {32'h439c3327, 32'h42a3fc2f, 32'hc56df933},
  {32'h440e68a2, 32'h4429c432, 32'h448de256},
  {32'hc47bcfcf, 32'h42e93813, 32'h44121c5e},
  {32'h4459c504, 32'h4385e805, 32'hc38a5129},
  {32'hc2bd5570, 32'hc5612b8f, 32'hc3a40bea},
  {32'h42b9e139, 32'hc404204a, 32'hc526bf12},
  {32'h440a5e9c, 32'hc42451c1, 32'h42c2976b},
  {32'hc509358e, 32'hc30914e9, 32'hc47971f3},
  {32'h440de3cc, 32'hc4221ff4, 32'h446d77c7},
  {32'h43d7a1d0, 32'hc4c67bd3, 32'h451073d7},
  {32'hc30a8818, 32'h44f6f235, 32'hc4b9738f},
  {32'h44a79c04, 32'h44088eed, 32'hc3d55d8a},
  {32'h4441d302, 32'hc4418e72, 32'h430f66fc},
  {32'hc4c88324, 32'h43088e16, 32'hc4793202},
  {32'hc33188c6, 32'hc3f4c978, 32'h446f36ae},
  {32'hc426a65e, 32'h42aeb2c2, 32'h421ff398},
  {32'h42659bbd, 32'h431caa92, 32'h448b8cc2},
  {32'h42978c66, 32'h44f31f5a, 32'h418da408},
  {32'hc4d8b4a6, 32'h439dd378, 32'hc21e9810},
  {32'hc54e3640, 32'hc4064e37, 32'h436c8222},
  {32'h446c97cb, 32'h4369c80a, 32'h438be3a3},
  {32'h44c3e6a6, 32'hc34185b7, 32'h42c22be2},
  {32'h43966c70, 32'hc49c318f, 32'hc3f7bca9},
  {32'hc40403e2, 32'h4501795a, 32'hc3756af2},
  {32'h410e762c, 32'h42b8be26, 32'h4334651e},
  {32'hc41ea908, 32'h450659aa, 32'hc41266fa},
  {32'hc40c7cb8, 32'hc4ddb603, 32'h43fdd9ea},
  {32'hc429c9d6, 32'hc3519c5e, 32'hc2761f23},
  {32'h424bcc82, 32'hc398d170, 32'hc4d5dc86},
  {32'h439954f5, 32'h44d12f73, 32'h45015b9a},
  {32'hc50ce818, 32'hc3ee1383, 32'h43283654},
  {32'hc4073007, 32'h427d8559, 32'hc542ff39},
  {32'hc4ff6d1f, 32'hc3e2dade, 32'h4338450d},
  {32'h42f300d0, 32'h4184baf5, 32'hc50c6c75},
  {32'h437b0a8e, 32'hc531daa3, 32'h43fd3faa},
  {32'hc480b7ce, 32'hc2887e13, 32'h42b49cae},
  {32'hc1daa7f0, 32'h443bfd94, 32'hc398d975},
  {32'hc50be5d6, 32'hc49da4d8, 32'h44cdd674},
  {32'h45277b41, 32'hc371558a, 32'hc422abfc},
  {32'h439f54b0, 32'h4369ef49, 32'hc45b1860},
  {32'hc45fcf2c, 32'hc3af9bf4, 32'h44e63940},
  {32'hc486ac12, 32'h4396890f, 32'hc3355b0e},
  {32'hc41ef99d, 32'hc48bc930, 32'h44262a53},
  {32'h44ae0c34, 32'hc29959b5, 32'h4288bc13},
  {32'h43d69cf9, 32'hc42b3fc3, 32'h445d71c5},
  {32'h4480036d, 32'hc44a555b, 32'hc3447c7b},
  {32'hc5087160, 32'hc2a3ad54, 32'h44008147},
  {32'h447760a5, 32'h42354859, 32'hc3b83986},
  {32'h4399dafa, 32'hc5805ad5, 32'hc336b0f8},
  {32'h452f2254, 32'hc3045dae, 32'hc28909b7},
  {32'hc40feceb, 32'hc4a0d77b, 32'h43661ab5},
  {32'h450e16f8, 32'h446cabf4, 32'h432e317f},
  {32'hc3862233, 32'hc4de0cb4, 32'hc3c98235},
  {32'hc37d56be, 32'h4426d1d5, 32'h431b5bc4},
  {32'hc3c63dde, 32'h438fceef, 32'h4401eb1b},
  {32'hc381e094, 32'hc41b3d95, 32'hc4b2427b},
  {32'h44860a5e, 32'hc3f01496, 32'h4470c8b5},
  {32'hc3aa5140, 32'hc4199f26, 32'h42914d76},
  {32'h44e59b28, 32'h42a13691, 32'h4493fa94},
  {32'hc3c06b89, 32'hc40575e2, 32'hc417f214},
  {32'hc4d132bf, 32'hc32c7837, 32'h42238ec8},
  {32'hc50dd3e6, 32'hc3cfa40e, 32'hc48a1f23},
  {32'h43feddd8, 32'h42bac3d1, 32'h44ec3129},
  {32'h4380b7f0, 32'hc4b880e6, 32'hc188ad66},
  {32'h4311b7d7, 32'hc37f3c29, 32'h44c5abd2},
  {32'h44466aa8, 32'h446ba7ab, 32'hc4db3c2c},
  {32'h44c403f0, 32'h432e7e47, 32'h43d43dda},
  {32'h43b0f9e3, 32'h42ae49e0, 32'hc4afaaa8},
  {32'h44a4a1a8, 32'h4382e94b, 32'h4491f4e8},
  {32'hc3f82d28, 32'hc44406fd, 32'h437101c9},
  {32'h452a9be7, 32'h43d5b6c1, 32'h43d21f23},
  {32'hc4146fb6, 32'hc30ce64f, 32'hc510cdcb},
  {32'hc3ea45c8, 32'h4432035e, 32'h43be9409},
  {32'hc48e0296, 32'hc50b8b52, 32'h43a19894},
  {32'h455f640e, 32'h441127ba, 32'hc3d46f4b},
  {32'hc48ad290, 32'hc3bc54b6, 32'hc3c39112},
  {32'h42b5ec31, 32'h454fdc80, 32'h43e7873e},
  {32'hc4457473, 32'hc526fe34, 32'hc0892a0a},
  {32'h4556f4eb, 32'h43a38f24, 32'h439693ca},
  {32'hc56f2b1a, 32'hc140e9c4, 32'hc3f4ba9b},
  {32'h444ee0e2, 32'hc3dd5547, 32'h43f3cdb4},
  {32'h438b6aac, 32'hc46e0725, 32'hc49f8ca2},
  {32'hc3c57d29, 32'hc4580999, 32'h4470488b},
  {32'hc3b33c56, 32'h4185e18d, 32'hc436f3e5},
  {32'hc4d88a14, 32'h436c9a1e, 32'h440b88ec},
  {32'h44e81169, 32'hc425b9e4, 32'h42bcd5df},
  {32'h429485b0, 32'h44b590f6, 32'h4481c3b0},
  {32'h4104d600, 32'hc3919243, 32'hc53c86a7},
  {32'hc52f797a, 32'hc399b7ef, 32'h440ff024},
  {32'h44be63a0, 32'hc3a6be50, 32'hc3e82f1b},
  {32'h446d53c0, 32'hc4a53c41, 32'h452249de},
  {32'hc42f6304, 32'hc32d29cf, 32'hc33fb3d9},
  {32'hc4f7b859, 32'hc3790a67, 32'hc39bcdc0},
  {32'hc37da3da, 32'hc3c918dd, 32'hc4bcc32d},
  {32'hc4673cda, 32'h449bdcf9, 32'h43e58cc8},
  {32'hc2c62e0d, 32'hc4d9975a, 32'hc38638da},
  {32'h43d4b21e, 32'h42c88c22, 32'h455012dd},
  {32'h4382d4c6, 32'h41800b3e, 32'hc50d1577},
  {32'hc4d97de0, 32'h42a0774c, 32'hc3169805},
  {32'h43b0d2b4, 32'hc4fce5e0, 32'hc16feb24},
  {32'hc53af95e, 32'h44580b74, 32'hc3308499},
  {32'hc39b7682, 32'hc50bfd18, 32'h4347ba58},
  {32'h432e636e, 32'h453047b1, 32'h442572df},
  {32'h450054b8, 32'hc3aeacd4, 32'hc3cbb8f7},
  {32'hc4c501e2, 32'h4358d821, 32'h42f6ef23},
  {32'h430289ec, 32'h43c9394f, 32'hc3c0753b},
  {32'hc51a8853, 32'hc3e26374, 32'h44255998},
  {32'h453faa74, 32'hc3d1c81c, 32'hc44dd140},
  {32'h4437716b, 32'hc3ccae6c, 32'h437a48f7},
  {32'hc571a0be, 32'h436ea511, 32'h4306ba2c},
  {32'h40b36900, 32'hc32e67a4, 32'h4545fc7e},
  {32'h44bf5a58, 32'h439e6365, 32'h424a6cc0},
  {32'h445830ce, 32'hc490b45a, 32'h43297a17},
  {32'h43654aa6, 32'h45607d68, 32'h43dd2107},
  {32'hc39b1804, 32'hc48f053e, 32'h42f2cd15},
  {32'hc400c82e, 32'h452b09e4, 32'hc36da88f},
  {32'hc32429cd, 32'hc45b8a4b, 32'h440261b4},
  {32'hc515a699, 32'hc2b669f5, 32'hc2116684},
  {32'h432eb540, 32'hc40237ae, 32'h442eb7cf},
  {32'hc2df39a6, 32'h43639f80, 32'hc4a47d83},
  {32'h4365884c, 32'h43081446, 32'hc4aa32ef},
  {32'hbf55f000, 32'h43baabfa, 32'h4443556b},
  {32'h43f81638, 32'hc51b94a6, 32'hc43cb03d},
  {32'h42bcf532, 32'h44d9c353, 32'hc196c3a5},
  {32'h4480c507, 32'hc4a37b7c, 32'hc3ac7d35},
  {32'h43b7c8ee, 32'h45006f94, 32'h43044233},
  {32'hc41ad0bf, 32'h4235f32d, 32'hc3d6c972},
  {32'hc53bc158, 32'h437b0a39, 32'h44027d22},
  {32'h43f23500, 32'hc44e4cb4, 32'hc4cb5e94},
  {32'hbf374920, 32'h44639540, 32'hc3a1c311},
  {32'h44d6ff09, 32'hc4016bcd, 32'hc398a96f},
  {32'h4304cb43, 32'h453a9a50, 32'hc1f41815},
  {32'h449328b1, 32'h4266f5d7, 32'hc47419f6},
  {32'hc4169063, 32'h44a97021, 32'h4371d3f9},
  {32'h43f5ebd5, 32'hc45f2c56, 32'hc4f410d4},
  {32'h45469fd0, 32'hc33516fc, 32'hc45336f7},
  {32'hc550564f, 32'hc427482b, 32'h4395e3c2},
  {32'h449281ca, 32'h434937f1, 32'h42edae75},
  {32'hc418540a, 32'hc49adea9, 32'h430f7f37},
  {32'h454634ce, 32'hc248024d, 32'hc3ef34d4},
  {32'h44ddd1be, 32'hc32c1aa5, 32'hc3b1ded7},
  {32'h42e6cde4, 32'h45122b87, 32'h44021150},
  {32'hc43e85d0, 32'hc50d0be6, 32'h436adef4},
  {32'h44ca07ac, 32'hc3775039, 32'h433a1df7},
  {32'hc4f8f626, 32'hc3b77a52, 32'hc2f4977b},
  {32'h44820c8e, 32'hc3e88bd2, 32'hc3d7414d},
  {32'h43cc8c92, 32'hc3bf0c17, 32'h44068921},
  {32'h4436af58, 32'h43f43310, 32'h44cd849a},
  {32'hc2d35d77, 32'hc51a2b8b, 32'hc3d9084d},
  {32'hc38550f8, 32'h42b18e78, 32'hc3d11092},
  {32'hc51dfce4, 32'hc4116713, 32'hc2241e51},
  {32'hc26d445a, 32'h45020cbd, 32'h4388268c},
  {32'h432e92b9, 32'hc49a7439, 32'hc3bea9cf},
  {32'h44e4bc46, 32'h432d4afb, 32'hc15656f8},
  {32'hc457fa02, 32'h446b1402, 32'hc491efd7},
  {32'h4513160d, 32'h43795bb0, 32'hc423fe48},
  {32'hc481d977, 32'hc44b66fa, 32'hc3a9ab85},
  {32'h452a6745, 32'hc3e210bd, 32'h43594788},
  {32'h44922f63, 32'hc1cf9eac, 32'hc415bc54},
  {32'h450bcdaf, 32'h43ffe564, 32'h4452688d},
  {32'hc4ada6f6, 32'hc2c22bdb, 32'hc3da8023},
  {32'h444c304c, 32'hc3c27e44, 32'h44625561},
  {32'hc47390fa, 32'hc3406f0e, 32'h4385383f},
  {32'hc4e6d80e, 32'hc4315436, 32'h439fba98},
  {32'hc2381840, 32'h45494371, 32'h4285e224},
  {32'h4275a5c0, 32'hc3f42fc0, 32'h433eb60c},
  {32'h453a7d3a, 32'hc1a95082, 32'hc1ca1aa8},
  {32'hc416e4ff, 32'hc4d30ee1, 32'hc31bce0a},
  {32'h45650431, 32'hc3a53f4e, 32'hc43fe234},
  {32'hc3d77654, 32'h4429ceae, 32'hc20b860f},
  {32'h447c9faa, 32'h441d5200, 32'h44518acd},
  {32'h44eba30d, 32'h4400c49f, 32'h42b0d147},
  {32'h4432c956, 32'h43fbf92e, 32'hc417c7a0},
  {32'hc449854c, 32'hc30e3f32, 32'hc3b8a63e},
  {32'hc420869a, 32'h418672dd, 32'hc40da378},
  {32'hc5414a19, 32'hc3f3a072, 32'hc3a9e5a3},
  {32'h4360f317, 32'hc305284d, 32'hc42477d5},
  {32'hc460464e, 32'hc3192ef8, 32'h43584bce},
  {32'h44efc816, 32'h43bb573c, 32'hc2c691aa},
  {32'h4026ec00, 32'hc338bee4, 32'h440ae1b5},
  {32'hc35d4d38, 32'h422079dc, 32'hc410e71c},
  {32'hc5335c53, 32'hc4007b55, 32'h43becf17},
  {32'h43ce39dd, 32'h456bf4da, 32'hc379f341},
  {32'h44e6a824, 32'hc3318eb1, 32'hc09b571e},
  {32'h454eb7a2, 32'h43bbdf3d, 32'hc3ef8bc1},
  {32'hc40f8763, 32'hc189cfbe, 32'h44aa4b00},
  {32'h44c284b2, 32'h4409f2ac, 32'hc302ac5e},
  {32'hc35fc3e0, 32'h4468453e, 32'h455e36af},
  {32'h4444b37d, 32'hc395eb91, 32'hc54fa2f7},
  {32'h440a1b55, 32'hc52329e4, 32'hc34555d2},
  {32'hc486d754, 32'h452fbb66, 32'h439b7548},
  {32'hc4437f58, 32'h434c6cc7, 32'h43f1f88d},
  {32'hc3f49268, 32'h440538c4, 32'hc434d5e0},
  {32'h450e922d, 32'hc3a3c439, 32'hc23c886f},
  {32'hc4d42696, 32'h42c3c564, 32'hc3aa99c6},
  {32'h4398d8c0, 32'hc48bd5c2, 32'hc4aa89a5},
  {32'hc54aef99, 32'h42e1ce47, 32'h42d06ec2},
  {32'h456ae15e, 32'hc2fc6f55, 32'h43516e2e},
  {32'hc477879f, 32'h44e25f58, 32'hc2d42bfe},
  {32'h44b45fdf, 32'hc4279840, 32'h44185b12},
  {32'hc34b18f0, 32'h448c9848, 32'h433bf26a},
  {32'h43d5c191, 32'hc50dbe8a, 32'h428a45e1},
  {32'h439a0aca, 32'h4381de09, 32'hc4a5751a},
  {32'hc47f28b4, 32'hc39d16bc, 32'h445d53eb},
  {32'hc3f23c68, 32'h44b22f29, 32'h447d2fb5},
  {32'h448c9cec, 32'hc38b6d43, 32'h444ef3d3},
  {32'hc51f1e82, 32'hc2aa9c36, 32'h43327284},
  {32'h44b111a3, 32'hc47e11fa, 32'h42ac054b},
  {32'hc437ee16, 32'h44ccbe2e, 32'hc4215f53},
  {32'h42ec4d98, 32'hc4dce795, 32'h429956c3},
  {32'hc2bbb7d8, 32'h455e7708, 32'h4315c0ce},
  {32'h43482768, 32'hc4b914f5, 32'h442c8f02},
  {32'h43c82a7a, 32'h444ff323, 32'hc37acd39},
  {32'h40563940, 32'h424ce9f0, 32'h443c7a33},
  {32'hc58517ca, 32'h428f0df5, 32'hc433981a},
  {32'h42786730, 32'h42a8d6ae, 32'h44c2b80b},
  {32'h438f8834, 32'hc4b379d1, 32'hc4b8ca3d},
  {32'h43628b68, 32'hc51349de, 32'h44cfeb28},
  {32'h44260542, 32'h4393457b, 32'hc333a478},
  {32'hc42ee3e5, 32'h439b3c03, 32'hc3777c6f},
  {32'h44d7f7a0, 32'hc4204010, 32'h4482085f},
  {32'hc302c35c, 32'h450d3b0f, 32'h43f83d1a},
  {32'h4357486e, 32'h42b7e300, 32'h44e8a015},
  {32'hc36d5270, 32'h44943928, 32'hc4d3491c},
  {32'h43a73836, 32'hc4258888, 32'h44926741},
  {32'h44610f02, 32'hc48e2165, 32'h44bcb5ec},
  {32'hc50711cc, 32'h441748a6, 32'hc41efb16},
  {32'hc3863004, 32'h438b0201, 32'h43e63066},
  {32'h45149c13, 32'h429f323d, 32'hc2d20828},
  {32'hc39cf3af, 32'hc3ad36cb, 32'h433d842a},
  {32'h4484c8c2, 32'hc29f5ba3, 32'h4381986f},
  {32'hc4504117, 32'hc317d27a, 32'hc46b1253},
  {32'h4317cfb0, 32'hc4fbe71c, 32'h42c9d6d0},
  {32'h4345a5f1, 32'h44ffbb0a, 32'hc3e92475},
  {32'h442f781d, 32'h4344b918, 32'h44168d9f},
  {32'hc4da9538, 32'hc41b5fbd, 32'h42908050},
  {32'h44662f48, 32'h432a6b79, 32'h449ae6bf},
  {32'hc5117bbf, 32'hc3013376, 32'h42d71aca},
  {32'h44119628, 32'hc49fea13, 32'hc38e3466},
  {32'hc4929905, 32'h43a95869, 32'hc1a29d53},
  {32'h44c920ce, 32'hc27b8926, 32'h426fac43},
  {32'hc48f39ab, 32'h44e4e93a, 32'hc3edd02c},
  {32'h4524a3e2, 32'hc4411ce3, 32'hc2d63e58},
  {32'h439a6961, 32'hc4e71235, 32'h43dd5901},
  {32'hc3c75c18, 32'hc2c7e1ff, 32'hc2858e96},
  {32'hc3a200c5, 32'h42c1e36e, 32'h448eb291},
  {32'hc38a36ce, 32'hc45011be, 32'h446fbbea},
  {32'h42bf8298, 32'h43f775ee, 32'hc48f34b3},
  {32'h441310d9, 32'hc4bec599, 32'hc39a4cd3},
  {32'h439c9993, 32'h433c8adc, 32'hc41acf12},
  {32'hc47dfe08, 32'h43a84a40, 32'h45075021},
  {32'h437d96db, 32'hc20244ef, 32'hc4735bb3},
  {32'hc4942635, 32'h43ba61a0, 32'h4392d182},
  {32'hc47686d4, 32'h44a60d2c, 32'h44bc523b},
  {32'h442a4faa, 32'hc3f77421, 32'hc48a330e},
  {32'h4396038a, 32'h438f45d8, 32'hc5345066},
  {32'hc4a78dbe, 32'hc488ae1f, 32'h442f64ec},
  {32'h44abf076, 32'h439c77e6, 32'hc3047ccb},
  {32'hc408fa40, 32'hc4b13bed, 32'h43a7f919},
  {32'h43ddfb64, 32'h44a06602, 32'hc4192027},
  {32'hc52adbd1, 32'hc3662860, 32'hc32f5da3},
  {32'h441b38ef, 32'hc44d2b1d, 32'hc4109a4b},
  {32'hc3a28478, 32'hc4186133, 32'h439e3a16},
  {32'h44d8e7f6, 32'h4321e8fe, 32'hc351a283},
  {32'hc503de3c, 32'hc4477fb9, 32'h430895c1},
  {32'h43425caa, 32'h4502beda, 32'h42f139d6},
  {32'h447b042d, 32'hc3762502, 32'hc3ac03fc},
  {32'h438b7cff, 32'h4535068b, 32'hc406d8da},
  {32'hc4f10fa4, 32'hc4370fc7, 32'hc2a3ecfd},
  {32'h4509f624, 32'hc3cd27ba, 32'h41819b28},
  {32'h44beb50e, 32'h40b3ac20, 32'h431cd799},
  {32'h43a7747c, 32'h44f8cf29, 32'hc4abdb55},
  {32'hc28841bf, 32'h41ce333b, 32'h44e77374},
  {32'h43d29e0e, 32'hc47912b4, 32'hc411de61},
  {32'h44907d49, 32'h4396b845, 32'h44263ade},
  {32'hc5213920, 32'hc455120c, 32'hc2025ac4},
  {32'hc4ce0967, 32'hc2d57c64, 32'h43a7cc1b},
  {32'hc50c7d93, 32'hc45232a6, 32'hc48853a8},
  {32'hc3b71476, 32'h4476ae89, 32'h44c70ffa},
  {32'hc3e65aa4, 32'hc32162b6, 32'hc348f57c},
  {32'h439bbd18, 32'h4433b334, 32'h449524fc},
  {32'h42931a24, 32'h42e269e8, 32'hc44cc6ae},
  {32'hc4f23a9d, 32'hc1f64580, 32'h439fa9de},
  {32'hc44e9392, 32'hc48c1621, 32'hc3ae8434},
  {32'h444b946a, 32'h44d3d89f, 32'h42b5b1d9},
  {32'hc4ab9269, 32'h43483a6c, 32'h43a62d57},
  {32'h4296c458, 32'h44a0a89d, 32'h448f3e72},
  {32'hc4f11478, 32'hc3f4ab08, 32'hc3efe6b6},
  {32'h437ffab7, 32'h44bd5c78, 32'h432f61df},
  {32'hc39c14f5, 32'hc50279d6, 32'hc3659ab2},
  {32'h4489eb54, 32'h44ff5032, 32'hc3c6b086},
  {32'hc310ba94, 32'hc4d8548c, 32'h42dd3413},
  {32'h44e682c6, 32'h4444479b, 32'hc3326029},
  {32'hc2d49640, 32'hc5394868, 32'h42bfa526},
  {32'hc4523fb4, 32'hc0b07eb4, 32'hc38cdc38},
  {32'hc2f64d80, 32'h4431286a, 32'hc469ca40},
  {32'h43aa4398, 32'h43bb43b4, 32'hc2972ce4},
  {32'h44431556, 32'hc4a371b9, 32'hc48b5cba},
  {32'h42cb7ea3, 32'hc3b10329, 32'h44cb361a},
  {32'hc4b4ced2, 32'hc24312b7, 32'hc313ed89},
  {32'h414647e0, 32'h441ab5ea, 32'h442c1bbb},
  {32'h444f0ea2, 32'hc405aeb0, 32'hc3c4b5d0},
  {32'h45071b1c, 32'h423c0af0, 32'h4346309c},
  {32'h432f7060, 32'hc3ec2f53, 32'hc543cfef},
  {32'hc4d7754a, 32'h43acf1c5, 32'h4463631c},
  {32'h44509b9b, 32'hc34c87e8, 32'hc3b008d6},
  {32'h435fdebf, 32'hc3f66fef, 32'h45034c43},
  {32'h44a2bf16, 32'h4413a0ce, 32'hc2e78b93},
  {32'h42f55c1c, 32'h4289f44c, 32'hc3649ab6},
  {32'h44022ec2, 32'hc4427816, 32'hc4882129},
  {32'hc425837d, 32'hc33268dc, 32'h4347ca44},
  {32'hc15d3703, 32'hc44068e6, 32'hc4171892},
  {32'hc3d1a9e8, 32'h43466792, 32'h449afe0b},
  {32'h43ae1bd8, 32'hc3e027a2, 32'hc500e2e1},
  {32'h43cb5e7a, 32'hc2d5f635, 32'h432e5d77},
  {32'h43aad836, 32'hc514e39a, 32'hc2cc45ce},
  {32'hc3a84061, 32'h453a8d8c, 32'h436d8607},
  {32'h4390442c, 32'h4342c162, 32'hc3a89d71},
  {32'h43e18040, 32'h445903a2, 32'h43c26e6c},
  {32'h448af2a3, 32'hc506a734, 32'h41c536bd},
  {32'hc3c56d3c, 32'h43c9bb47, 32'h4348ae3e},
  {32'h44a8d2fe, 32'hc3c432a1, 32'hc41763f3},
  {32'hc5142d2b, 32'hc4287f1a, 32'h4284607e},
  {32'h44307ebd, 32'hc36083d8, 32'hc3111623},
  {32'h44eb5c50, 32'h3fb173f0, 32'hc289b1d8},
  {32'hc41d4b77, 32'hc330de13, 32'hc4864458},
  {32'h4496fccd, 32'h43d04aab, 32'h43d81874},
  {32'hc3c8aff6, 32'h4480b4b7, 32'h4178fda5},
  {32'h454cb6e8, 32'hc3a835d0, 32'hc20389db},
  {32'hc451ab80, 32'h44fc8d75, 32'h440ac21b},
  {32'hc4b089af, 32'hc3b83a66, 32'h438268b8},
  {32'hc4f327f7, 32'h42f02ba9, 32'hc1dbe58c},
  {32'h44985212, 32'hc4611b3a, 32'hc3229386},
  {32'h4389ba3c, 32'hc40fb1cd, 32'hc4fd4c4e},
  {32'h44ad8cf0, 32'h4327def0, 32'h443e6926},
  {32'hc4ca02a5, 32'hc431fce4, 32'h436f923b},
  {32'hc383a08a, 32'hc49d7151, 32'h4352611c},
  {32'hc4b0dd1e, 32'h440001b5, 32'h43d98c62},
  {32'h43df3ccc, 32'hc4acf11d, 32'hc40df176},
  {32'h432a5662, 32'hc3919255, 32'hc353e0ea},
  {32'h44b7e0cb, 32'hc494b805, 32'h42411920},
  {32'hc45fbb72, 32'h42da85da, 32'h44c64400},
  {32'h45158e7e, 32'h438ac78d, 32'h43d01bdd},
  {32'hc47f8f1f, 32'hc43402d6, 32'h4410fc61},
  {32'h451e0369, 32'h44106712, 32'hc40cee15},
  {32'hc3248bde, 32'h43cd874f, 32'h42c15667},
  {32'hc0c90a70, 32'hc484a3d4, 32'hc477681a},
  {32'hc4cced4a, 32'h42851efa, 32'hc2555565},
  {32'h441ba4ae, 32'h43b1a7ad, 32'hc491439f},
  {32'hc48c083e, 32'h44018f52, 32'hc29936ee},
  {32'h4413f290, 32'hc4e14570, 32'hc31c1f2c},
  {32'h44cbb47e, 32'h43575f8a, 32'hc51033d8},
  {32'hc493715c, 32'hc38d9fa9, 32'h43bab5b0},
  {32'h447b425d, 32'h43a19589, 32'hc31ce0cc},
  {32'hc4e7f3ee, 32'h4382c01f, 32'h43081b06},
  {32'h44e2cf52, 32'h44196553, 32'h436ec3da},
  {32'hc4ab8bde, 32'hc331f08c, 32'h430b6aca},
  {32'hc3453cd0, 32'h44b8967a, 32'h43605098},
  {32'hc24b8550, 32'hc5053bb6, 32'hc2fb7d86},
  {32'hc44de078, 32'h4386875b, 32'hc1bf5fa3},
  {32'hc0eec200, 32'hc461ef19, 32'hc43b992b},
  {32'h441955a2, 32'h43ec9e54, 32'h40cf4da6},
  {32'h43a6f52d, 32'hc249821c, 32'h44895955},
  {32'hc1c1293c, 32'h44f5cc76, 32'hc30d27fb},
  {32'hc443e8d8, 32'hc4404920, 32'hc5132aa5},
  {32'hc362d7a0, 32'h4478b1db, 32'h43d9c785},
  {32'hc178bab0, 32'hc472fe85, 32'hc3dee1ea},
  {32'h435a43b6, 32'h4513aeb2, 32'hc11064a2},
  {32'h42f4a160, 32'hc3ac92ff, 32'h43fc7a96},
  {32'h457b3033, 32'h422ccc78, 32'h43a26514},
  {32'hc513dfac, 32'h43e5f78e, 32'hc4457159},
  {32'hc49eb34b, 32'hc2ad7484, 32'hc256f296},
  {32'hc3cd3306, 32'hc516f5ae, 32'hc463557f},
  {32'hc24041eb, 32'h44f7b52b, 32'h42130a4d},
  {32'h448c7919, 32'hc3cb8abb, 32'h4249035d},
  {32'h43dd7678, 32'h449fc791, 32'h45084d93},
  {32'hc4a59ddc, 32'hc426ba04, 32'hc3a3ac6e},
  {32'hc4400849, 32'hc359261d, 32'h43313b97},
  {32'h421368d0, 32'hc2a13b14, 32'hc395f95b},
  {32'hc441d016, 32'hc47b0917, 32'hc2525560},
  {32'h4433a088, 32'h44c32c47, 32'h4396d50f},
  {32'hc3c10ec2, 32'hc498e30b, 32'h4412e191},
  {32'h43b31280, 32'hc32ea8a4, 32'hc20b2a9e},
  {32'hc42f78f4, 32'hc5225cbc, 32'h42e90c7b},
  {32'hc2792b38, 32'hc2a3dd18, 32'hc448da96},
  {32'hc598632b, 32'h442f4217, 32'hc3dcf579},
  {32'h450d44f4, 32'h42f84f5f, 32'h42684555},
  {32'hc3879f2a, 32'hc431d50f, 32'h43b746cf},
  {32'h43abb0cd, 32'h4516a0d9, 32'h43271b21},
  {32'hc3f9c4fc, 32'hc4b225b6, 32'hc3ba62aa},
  {32'hc340823c, 32'h44b09159, 32'hc3962ed4},
  {32'hc4d0fdef, 32'hc36fea40, 32'h43c2e824},
  {32'h44c90606, 32'h4325c0e3, 32'hc3beec1b},
  {32'hc1f0baf0, 32'hc32e05ba, 32'h44dba049},
  {32'h439c0c24, 32'hc413ef29, 32'hc4db23be},
  {32'hc4a1e94c, 32'h43dd144d, 32'h43bab82f},
  {32'h44ab08b2, 32'h441bdfc1, 32'hc3a5514c},
  {32'hc3684510, 32'hc4ed75ac, 32'h43dd21ed},
  {32'h44dbc146, 32'h44b58360, 32'hc398c801},
  {32'hc49fd0ca, 32'h41d55da6, 32'h43c6b65a},
  {32'h4503ec12, 32'h445078eb, 32'hc35925e5},
  {32'hc2f6afea, 32'hc5296e86, 32'hc3d6d42d},
  {32'h44ede0f8, 32'h439956ed, 32'hc33eddaa},
  {32'hc4e21797, 32'h43d4928d, 32'h4333a816},
  {32'h44dcba3b, 32'hc31c84f7, 32'hc445877d},
  {32'h4480fa8c, 32'hc49ef169, 32'h41ff97f5},
  {32'hc538dfd3, 32'h4405713c, 32'h43b58b72},
  {32'h43f95eb4, 32'h4310a6ce, 32'h4424b17a},
  {32'hc50e25ba, 32'h4422c5d3, 32'h435733f4},
  {32'h4552ce0d, 32'h43493ba0, 32'hc1ecad16},
  {32'hc4e86828, 32'hc13d2bf7, 32'h41e672d3},
  {32'h44bdcb92, 32'h43480382, 32'h4219e4bf},
  {32'hc5855d4f, 32'hc335ea1b, 32'h4347fd58},
  {32'hc4c98139, 32'hc2b4826a, 32'h4401e4a8},
  {32'hc4075900, 32'h44714320, 32'hc4d0184e},
  {32'h44327bb1, 32'hc3b6ee81, 32'hc402337f},
  {32'h44bde167, 32'h438f38e5, 32'hc429582a},
  {32'hc2e5afd9, 32'hc5571ee3, 32'hc2102278},
  {32'hc32b1438, 32'h41002448, 32'hc44b1cab},
  {32'hc2c1c664, 32'hc3ac75bd, 32'h44bf0943},
  {32'hc3d2a608, 32'hc2e23285, 32'hc420bbc2},
  {32'h441576e9, 32'h439a3bb3, 32'hc424b135},
  {32'hc38c7728, 32'hc36cf2af, 32'hc49d6e65},
  {32'h43a988f3, 32'hc52885d4, 32'hc39792a6},
  {32'hc42030fc, 32'h45000883, 32'hc38f3a3d},
  {32'hc4990bd3, 32'h413b608e, 32'h438de037},
  {32'h41dd6830, 32'h44d7057b, 32'hc361772a},
  {32'h44de7960, 32'hc3c62412, 32'hc3e513b0},
  {32'h44cd6040, 32'hc1bba196, 32'hc2831c50},
  {32'h44f17a82, 32'h43b2e7bc, 32'h4474b51f},
  {32'hc4cf1372, 32'hc3feb77d, 32'hc4ce0897},
  {32'hc437533a, 32'h4386821a, 32'h440f6d17},
  {32'hc1d4b580, 32'h4487bffd, 32'hc4d155be},
  {32'hc2d3da78, 32'h4490130d, 32'h4519fade},
  {32'h42510758, 32'hc3bd8f23, 32'hc3b5b1f7},
  {32'hc48be237, 32'h4254f306, 32'hc31d9234},
  {32'h44a463aa, 32'h421d1b0f, 32'h432d0d54},
  {32'hc3a3eb5a, 32'h4487ce82, 32'hc4498307},
  {32'hc461c991, 32'hc406f7d4, 32'hc3667055},
  {32'hc4923c1f, 32'h43f0060a, 32'hc46c548c},
  {32'h440630e5, 32'hc491962c, 32'h44c44fd6},
  {32'h42985428, 32'h44b3dc81, 32'h44c24445},
  {32'hc4ca2b90, 32'hc218d216, 32'hc4eff6b7},
  {32'hc2c8e886, 32'h43106247, 32'h43212308},
  {32'hc242d4c0, 32'hc42c38c3, 32'hc29767b0},
  {32'hc3160cf4, 32'h43b61bbe, 32'hc5308c96},
  {32'h43923ea8, 32'hc5129b60, 32'hc38adf29},
  {32'hc385c088, 32'hc1abc983, 32'h435fffbb},
  {32'h451f0caa, 32'hc32d6811, 32'h44178d58},
  {32'hc46425f5, 32'h436b7718, 32'hc4aee71c},
  {32'h4529eb9d, 32'hc3f9857c, 32'hc3630dd0},
  {32'hc529d494, 32'h43dda696, 32'hc3a7d14c},
  {32'h4568167f, 32'hc3c5f03e, 32'hc3c50c62},
  {32'h44458184, 32'h44bc10f9, 32'h4395d436},
  {32'h437fc650, 32'hc54a329c, 32'h431c5d28},
  {32'hc2d89b0a, 32'h454b5bf6, 32'h42c10a28},
  {32'h44abd17e, 32'hc4005947, 32'h4317da9a},
  {32'hc56b1d25, 32'h43eb6d25, 32'h43d807bc},
  {32'hc3822b68, 32'hc4dd9b9a, 32'hc2e9a396},
  {32'h43e0d842, 32'hc2a0f317, 32'h4470c37c},
  {32'hc0760221, 32'h44477f9e, 32'hc4e1f349},
  {32'hc2e68c88, 32'h435c9dee, 32'h44df3b90},
  {32'hc424cde3, 32'hc4eb750d, 32'h438daad1},
  {32'h45334d95, 32'h43057bab, 32'h438b5c30},
  {32'h44d51f87, 32'hc4431065, 32'h4212696f},
  {32'h43857916, 32'h447bf66d, 32'hc4be479b},
  {32'hc5276f58, 32'h42bc839c, 32'h40d1b330},
  {32'h443a6248, 32'hc3849b8b, 32'h43e21c1b},
  {32'h44601692, 32'hc327d3b5, 32'hc407509b},
  {32'h41d275f8, 32'h436d3c09, 32'h44f92b8b},
  {32'hc414525c, 32'h44c5e84d, 32'hc508aea2},
  {32'h44dde8b5, 32'h4457e130, 32'hc3bf667e},
  {32'hc4bfc914, 32'hc445b3e1, 32'h440224b8},
  {32'h45029fa5, 32'hc28d12bb, 32'h41bd07d6},
  {32'hc46a133a, 32'hc3f91e01, 32'h451a46cd},
  {32'h43538a4e, 32'hc3b68b4e, 32'hc4d20f37},
  {32'hc41e4677, 32'hc487bec9, 32'h42542ce8},
  {32'h439587f0, 32'h420c5c8f, 32'hc4436c32},
  {32'hc53e648a, 32'h42e6e18c, 32'hc236a149},
  {32'hc4df4b4a, 32'hc3962ad0, 32'hc328fbae},
  {32'hc4de5170, 32'hc48170bc, 32'h42537596},
  {32'h43b7fe0c, 32'h448b07b2, 32'h43c0e579},
  {32'hc513e13a, 32'h425a4268, 32'h44096603},
  {32'h444f9fa8, 32'h442e9112, 32'h445d399e},
  {32'hc3bc364c, 32'hc4c2c209, 32'hc2826b00},
  {32'h42f7f6b3, 32'h444e4aa9, 32'hc40fd0f6},
  {32'h43bfb010, 32'hc4a41ab2, 32'h43fe33be},
  {32'h433bba70, 32'h4430d3af, 32'hc5173311},
  {32'h44119720, 32'h44388644, 32'h43c07bcb},
  {32'h43a352a0, 32'hc403fc5b, 32'hc40a20c4},
  {32'h43a8bbe6, 32'h438e2059, 32'h4441de7e},
  {32'h4366c5ad, 32'hc41f9498, 32'hc4cde315},
  {32'hc3190b1e, 32'h4406ccea, 32'h4405e822},
  {32'hc397c398, 32'hc43ed17b, 32'hc488d8ef},
  {32'h452980cf, 32'h43c2a169, 32'h4422d9f1},
  {32'h43e1042c, 32'hc40ae986, 32'hc3c5c3fe},
  {32'hc290cc7c, 32'h44597c1f, 32'h44608964},
  {32'hc476b398, 32'hc2981fd2, 32'hc42249c5},
  {32'hc21a4d9b, 32'h440a70ed, 32'h43354f29},
  {32'hc4b06085, 32'hc401f654, 32'hc433976c},
  {32'h43b41f26, 32'h44bef222, 32'h435b4b93},
  {32'h448a83cc, 32'hc4256ef9, 32'hc3a887db},
  {32'hc406b508, 32'h44dd1191, 32'h4506b3b3},
  {32'hc3b22730, 32'h4220e6bd, 32'hc3839840},
  {32'hc43f7708, 32'h441951a5, 32'h4317cedf},
  {32'hc4de8424, 32'hc49d1bd9, 32'h435282e8},
  {32'h43af5f70, 32'h4568dc53, 32'h42fa57c8},
  {32'hc5178830, 32'hc2b25be1, 32'hc2ab22a5},
  {32'h446bbf1c, 32'h4464fe45, 32'h441cd77d},
  {32'hc4505f4f, 32'hc44d119a, 32'hbf0b4380},
  {32'hc4b2bef4, 32'hc182a3a4, 32'h43b34633},
  {32'hc485684e, 32'h44639dd1, 32'hc31b8272},
  {32'h440e9857, 32'hc38373ab, 32'h43d1e7c3},
  {32'h4392b8ab, 32'h449c9a14, 32'hc4855a11},
  {32'hc2e1a6d4, 32'hc47a2f72, 32'h449b6de1},
  {32'hc3b69e0f, 32'hc4844176, 32'hc317121a},
  {32'h4326a5fb, 32'h4520523e, 32'h43f4acf9},
  {32'h42b59f0d, 32'hc5513d95, 32'hc36ab266},
  {32'hc4c01432, 32'hc3223f5e, 32'h4241c163},
  {32'h431b2760, 32'hc4f2eb40, 32'hc4c8c97e},
  {32'hc426847c, 32'h445831ed, 32'h44916af6},
  {32'h44b26a14, 32'hc41e7032, 32'hc2698f65},
  {32'hc33b77aa, 32'hc48f7a7f, 32'h44bb1149},
  {32'h44616846, 32'h440c0642, 32'hc431c65e},
  {32'h434ee7c2, 32'h4343bc07, 32'h43e06b4e},
  {32'h4419c8d4, 32'hc3f4f574, 32'hc43796af},
  {32'hc523bc2e, 32'h43dd8884, 32'h423697de},
  {32'h44547ff4, 32'h41b8ecaa, 32'hc42d27e8},
  {32'hc40fd832, 32'h42cb50fc, 32'h449a20ce},
  {32'h447ef414, 32'hc3800ba5, 32'hc4b92990},
  {32'hc28f2efe, 32'h42b2c94e, 32'h4498cf1c},
  {32'h453e3239, 32'hc3eeb7da, 32'h43619a97},
  {32'hc4308cc8, 32'h4452d6f6, 32'h4427fb7c},
  {32'h452d23b2, 32'h446522f6, 32'h443d5ed3},
  {32'h43c07e0e, 32'h456c2972, 32'hc286bf94},
  {32'hc362adb0, 32'hc400281c, 32'hc1ea013c},
  {32'h44049633, 32'h4492eba0, 32'hc382d64a},
  {32'h42d08aa0, 32'hc33cea31, 32'h4324c102},
  {32'hc46fcc50, 32'h43f620b3, 32'h438eef10},
  {32'h452240eb, 32'hc3f0bfdc, 32'h42dc4660},
  {32'h45188bcd, 32'hc382fc62, 32'hc39e4b5f},
  {32'hc336f738, 32'hc1f849ec, 32'hc4b02645},
  {32'h442bb5d4, 32'hc1fc4922, 32'h4546fb07},
  {32'h44d632ab, 32'h438f2f73, 32'h434ce057},
  {32'h455b8a28, 32'h42f5b189, 32'h431c26df},
  {32'hc36b02a2, 32'h44653082, 32'hc36a5a9d},
  {32'h45292745, 32'h42860fa6, 32'h43296bd5},
  {32'hc486f547, 32'h444685eb, 32'h432aa419},
  {32'h43ad71ea, 32'hc55e3cee, 32'hc0908976},
  {32'h44dbf6cf, 32'hc1956362, 32'hc3f17265},
  {32'h43daa40c, 32'h42b3b46e, 32'h449724f5},
  {32'hc4557caf, 32'hc3ad5e59, 32'hc38b1848},
  {32'hc3987122, 32'hc49ea162, 32'hc10c3036},
  {32'hc3d34422, 32'h44392e3c, 32'h440071cf},
  {32'h44399e69, 32'hc426dc7b, 32'hc49b5969},
  {32'h44a60876, 32'h43d3934a, 32'hc297ffd0},
  {32'h45083290, 32'h438966ed, 32'hc3b31245},
  {32'h43fdaf22, 32'hc415430f, 32'h43e02076},
  {32'hc49030d1, 32'hc3fa9d3b, 32'hc30f7311},
  {32'hc51cd0f9, 32'hc4751cc7, 32'h44177d90},
  {32'h4503b858, 32'h4403c889, 32'hc4530671},
  {32'hc49e77be, 32'h42a44ec1, 32'h431286b4},
  {32'h43f40d90, 32'hc42b1662, 32'hc43a7ef9},
  {32'hc387e7e7, 32'h448a1bf6, 32'h43a352cd},
  {32'hc38171d1, 32'h43bd0416, 32'hc477a796},
  {32'hc4551928, 32'h44ae8864, 32'hc3eeb1bb},
  {32'h44778a32, 32'hc4870bc4, 32'hc4dd8c77},
  {32'h432eee10, 32'hc3c5ae32, 32'hc52de943},
  {32'hc420293a, 32'h44d359b4, 32'h4515580d},
  {32'h45096d5a, 32'hc355c3c4, 32'h43c3ccc9},
  {32'hc23313cd, 32'hc543af87, 32'hc43a9525},
  {32'h44d77036, 32'hc149ef10, 32'h43d9865a},
  {32'hc506b100, 32'hc40179eb, 32'hc22524b8},
  {32'h44012fce, 32'h454f03dc, 32'h4379390f},
  {32'hc50f77c6, 32'hc45f03e3, 32'hc28f95a4},
  {32'hc2f1a1bc, 32'h43dca377, 32'h42bf4eb7},
  {32'hc3db9e5c, 32'hc41dcf44, 32'hc404b160},
  {32'h44435690, 32'h4462e81f, 32'h446c4af2},
  {32'hc48a0da9, 32'h43708643, 32'h4487614d},
  {32'hc232decd, 32'h439abffa, 32'h451662be},
  {32'hc4032530, 32'h429fafac, 32'hc4456352},
  {32'h4484267a, 32'h43a1c91d, 32'h42e45d65},
  {32'hc3843bca, 32'hc54cef88, 32'h4383f59f},
  {32'h441950c2, 32'h4505cf3b, 32'h447457b9},
  {32'hc5071d68, 32'hc08f0809, 32'hc3c1751c},
  {32'h45433f28, 32'hc41d91c0, 32'h43313cca},
  {32'hc5169c58, 32'hc3fc3cc0, 32'hc40c1c6c},
  {32'hc44cd871, 32'h43531ee0, 32'h431c808e},
  {32'h43824860, 32'hc3e5bca9, 32'hc544d81a},
  {32'h42bb92bf, 32'h44f12a14, 32'h44c45955},
  {32'h438f1440, 32'h42b04a98, 32'hc49d59af},
  {32'hc2e873d6, 32'h42f6ac66, 32'h452228e1},
  {32'hc5200234, 32'hc1cc4ae4, 32'hc39c0689},
  {32'h44930b3c, 32'h4466e572, 32'hc3cb0530},
  {32'h44b346b2, 32'hc446e4bd, 32'h41a48b4e},
  {32'h431b0457, 32'hc5197b7c, 32'hc3a65852},
  {32'hc39b0ed3, 32'h4532199f, 32'h42596720},
  {32'hc40eff50, 32'hc437393f, 32'h42e44d54},
  {32'h444ef080, 32'h44dc1534, 32'h4339f229},
  {32'hc5214a80, 32'hc386a1b1, 32'hc1c3186b},
  {32'hc4f7ffa8, 32'h43569bf8, 32'h429723c0},
  {32'hc44c9df7, 32'h43d38327, 32'hc4808872},
  {32'h45495c92, 32'h42c6814f, 32'h4420c0f6},
  {32'hc40dd922, 32'hc430e74e, 32'h43d16fe9},
  {32'h4441c4b9, 32'h444659b9, 32'hc50178a9},
  {32'h42ea987c, 32'hc4a7903a, 32'h43a75890},
  {32'h449ce12e, 32'hc1eefb36, 32'hc3f367f8},
  {32'hc3b369e0, 32'hc47ab9bc, 32'h439365df},
  {32'h44c64bf6, 32'h444fbef8, 32'h4323a121},
  {32'hc40f75ab, 32'hc3a6c863, 32'h4410eef8},
  {32'h44918239, 32'hc37b3c10, 32'hc48345cc},
  {32'hc50ff258, 32'h41c50447, 32'h42dff410},
  {32'h449838e7, 32'h445ed634, 32'hc3bb5903},
  {32'hc520907a, 32'hc3edaa6f, 32'h42c29f53},
  {32'h444e07d0, 32'h44abb8c9, 32'hc4afcfed},
  {32'h4063e940, 32'hc3bd0e3c, 32'h44c58be9},
  {32'h4306cc12, 32'hc3847722, 32'hc4c531f4},
  {32'hc380d504, 32'hc4542223, 32'h43b46afc},
  {32'h4466671c, 32'h42c7c9b6, 32'hc4278bce},
  {32'hc11fa600, 32'h434a888e, 32'h451589a0},
  {32'h450158a6, 32'h433aabc5, 32'hc3f50d66},
  {32'h432d03b1, 32'h44055ffb, 32'hc4c52901},
  {32'hc4caf2a2, 32'h449a33c3, 32'h4312ad11},
  {32'hc45722d2, 32'hc46bf2fa, 32'h43a4b95d},
  {32'hc429ff6a, 32'h44de8857, 32'hc3c88f06},
  {32'h44f41cc9, 32'hc4717044, 32'hc3d2cf32},
  {32'h43cfb675, 32'h44f30e56, 32'hc3340ea7},
  {32'h445ad118, 32'hc3e34aa4, 32'hc3729d23},
  {32'hc4c16e36, 32'h43b2f953, 32'h439c4a62},
  {32'h42e6c88c, 32'hc45e5f79, 32'hc416736b},
  {32'hc4a6f3f2, 32'h4383e0e6, 32'h41b12c97},
  {32'h4488f8b0, 32'hc249a3a3, 32'h446cc852},
  {32'h442b411e, 32'hc2539ccd, 32'h43b54248},
  {32'h45784555, 32'h435dda33, 32'hc299309e},
  {32'hc38e07a5, 32'hc2a11396, 32'hc40c516c},
  {32'h41be6578, 32'h432d5a36, 32'h43f74f96},
  {32'hc5116d30, 32'h439e0f87, 32'h4414e1c1},
  {32'h44a93b03, 32'hc47ad532, 32'h434b0f22},
  {32'h44f20cef, 32'hc2eecdfb, 32'h43524e4b},
  {32'h44fd302b, 32'hc3c5e47f, 32'h44b7fde0},
  {32'hc445621c, 32'h448ccfd9, 32'hc4b5c7f2},
  {32'hc4952e1f, 32'hc3998572, 32'h43a0cf16},
  {32'hc21ad5a0, 32'h44d57e09, 32'hc41d833b},
  {32'hc2a5a687, 32'hc4f75240, 32'h443c5e31},
  {32'h441be514, 32'h430cff57, 32'hc3246d72},
  {32'h45681d0b, 32'h3fea97ee, 32'h44295212},
  {32'hc4a4ce2c, 32'hc43abb83, 32'hc43af592},
  {32'h450b820c, 32'hc30a4879, 32'hc2ddd9c6},
  {32'h4308e508, 32'hc504718a, 32'hc4ab19ed},
  {32'h448035b3, 32'h44128f0a, 32'h4488ed4d},
  {32'hc40f39cb, 32'h43b84b38, 32'hc437ca83},
  {32'hc3958563, 32'h43b2e4e5, 32'hc33c66bc},
  {32'h450dcadd, 32'h42342cc9, 32'h43bc8e53},
  {32'hc3e9ae22, 32'hc3e6bc5e, 32'hc49f0762},
  {32'hc4dfbe38, 32'h43b094db, 32'hc3f6f357},
  {32'hc4953b1c, 32'h445a393a, 32'hc3ce0e1d},
  {32'h44f29271, 32'hc21c994c, 32'h43e6baa1},
  {32'hc3a20afa, 32'h45066809, 32'h4508829b},
  {32'hc2a164a8, 32'h43a30acd, 32'hc536a8aa},
  {32'h44e0b768, 32'hc408e89b, 32'hc36f5e9a},
  {32'h43d238b2, 32'h43fac257, 32'h448d566c},
  {32'hc3cf30de, 32'h4356a81d, 32'hc4eddc97},
  {32'h43059093, 32'hc4eb4c27, 32'h4254418d},
  {32'hc5006692, 32'hc35a5cfb, 32'h43a79b00},
  {32'h4302f310, 32'hc4d14d96, 32'h44560999},
  {32'h42b865a0, 32'h450713eb, 32'hc335ae48},
  {32'hc40c7c0b, 32'hc41439b8, 32'h431c551b},
  {32'hc284b138, 32'hc37cb932, 32'h43881da4},
  {32'h4423d4f8, 32'h43f2adb9, 32'h449c238e},
  {32'hc50c6550, 32'hc35c4cc9, 32'h4406eb6e},
  {32'hc2bb228f, 32'hc556e339, 32'hc2787163},
  {32'hc5225363, 32'hc300c49f, 32'h43d379f2},
  {32'h4545916b, 32'h43e3f565, 32'h43c4f7f0},
  {32'hc515d3b4, 32'h4427e251, 32'hc3a46939},
  {32'hc3a857dc, 32'hc52c1226, 32'h43d290de},
  {32'hc4b53b54, 32'hc38e77cf, 32'hc2e8a35e},
  {32'hc4a96483, 32'h431d78c8, 32'hc4916f5f},
  {32'hc2c7c4c4, 32'hc31c2a4a, 32'h44bfed1f},
  {32'h4363073f, 32'hc3f53796, 32'h45336b07},
  {32'h4391a56b, 32'h44c63a3b, 32'hc39ab60a},
  {32'hc40adf2f, 32'hc2b0a1c7, 32'h450378c2},
  {32'h45032c2f, 32'h44027d1e, 32'hc3b603a3},
  {32'hc2708230, 32'hc4f876da, 32'hc1bfe284},
  {32'h429fc3ae, 32'hc3855fb5, 32'hc3e0dd12},
  {32'h41057bd0, 32'hc2ba7e9b, 32'hc48e2a8b},
  {32'h438ceb38, 32'hc410d56a, 32'h44f895b6},
  {32'h42591040, 32'h44aa80e1, 32'hc507a98b},
  {32'h4384465e, 32'hc38b435d, 32'hc51a0c43},
  {32'hc3ff5e70, 32'hc4d130b5, 32'h44128258},
  {32'h4485e95a, 32'hc2d963f6, 32'hc3da592e},
  {32'hc3e520d6, 32'hc4bfee12, 32'h439b3a39},
  {32'h428d5a08, 32'h448f7008, 32'hc41d10a5},
  {32'hc29a6c05, 32'hc45a2a6b, 32'h429b63c4},
  {32'h42bb45a3, 32'hc449e653, 32'hc3d0c31b},
  {32'hc4c46886, 32'h433a297c, 32'hc33b95fd},
  {32'h44769b71, 32'h43c5f6f1, 32'hc2804f17},
  {32'hc49a3430, 32'hc48f4b35, 32'hc390ea00},
  {32'h4437da4a, 32'h44566988, 32'h43d0aa34},
  {32'h43dd92e2, 32'hc48b7993, 32'hc2e5c8fb},
  {32'h453d691c, 32'h44274163, 32'h43cd92ad},
  {32'hc457748b, 32'hc4b20e22, 32'hc40d4b90},
  {32'h4397a844, 32'h418b67e9, 32'h42d4aa7e},
  {32'h43475f68, 32'h43876748, 32'h4415b292},
  {32'hc3846284, 32'hc4b88ddb, 32'hc3fcdbf5},
  {32'h40f93f80, 32'hc4cc8093, 32'h4511f235},
  {32'hc2e30cb7, 32'hc38b3571, 32'h4250aa9e},
  {32'h448e8ab6, 32'h43b89d87, 32'h447ba2b4},
  {32'h4088bed7, 32'hc43c9c7a, 32'hc4a434d1},
  {32'h4362a31f, 32'h44aaef96, 32'h4353b01f},
  {32'h4403d7fd, 32'hc4923885, 32'hc53dd42f},
  {32'h44238c3e, 32'h43d811e4, 32'h443149fa},
  {32'hc38bc063, 32'h4458a013, 32'h42bb6142},
  {32'hc46dc6de, 32'hc3d1cfda, 32'h4508f368},
  {32'hc45a74b5, 32'hc4820e6b, 32'hc36ec323},
  {32'h42d744aa, 32'h449a25a6, 32'h40f034fe},
  {32'hc4370697, 32'hc3942f0d, 32'hc494531c},
  {32'h43b6d5ec, 32'hc31de90c, 32'h44eeaff6},
  {32'h4446c2b0, 32'h43ab1d76, 32'h429d4c3e},
  {32'h44e3f200, 32'hc14d5fde, 32'hc305fca5},
  {32'hc32ec808, 32'hc4ae347f, 32'hc5427162},
  {32'h444b60ef, 32'h446e5569, 32'h4309e792},
  {32'hc4b3be32, 32'hc4b8b8f9, 32'hc30bd7fb},
  {32'h44c23c31, 32'h44abf1f0, 32'h43881dad},
  {32'h44d52400, 32'hc2be8322, 32'hc34d0290},
  {32'h455319dd, 32'h43eb6eb8, 32'hc1f8324d},
  {32'hc48893ac, 32'hc4a36562, 32'h428c776b},
  {32'hc48149a8, 32'h42be271c, 32'h43a3fd42},
  {32'hc4cb351c, 32'h4450d789, 32'h43183804},
  {32'h44d55a56, 32'h439be450, 32'h44325e82},
  {32'h44744798, 32'h44350c59, 32'hc4d440a4},
  {32'hc511715d, 32'h441b610f, 32'h444ed02b},
  {32'hc27e6b84, 32'h449fd249, 32'hc40c9de7},
  {32'h432eb1ce, 32'h448c96c0, 32'h44f1c32b},
  {32'h430dfdec, 32'hc419e83f, 32'hc492a5b3},
  {32'hc5189235, 32'hc36241be, 32'h4237f012},
  {32'hc1749480, 32'hc394355b, 32'hc5504737},
  {32'hc5031a90, 32'h43bdb246, 32'h448eda9f},
  {32'h44fe9a10, 32'h437cce26, 32'hc4777d65},
  {32'hc3c1826a, 32'hc4cfc612, 32'h44dd5d29},
  {32'hc2442842, 32'hc20e5f52, 32'hc420428e},
  {32'h44196cba, 32'h426988f9, 32'h435e372a},
  {32'h450da5ff, 32'hc47fa475, 32'h4395efde},
  {32'hc3c73a50, 32'h44f1f108, 32'hc39c50ab},
  {32'h44718917, 32'h43776a8a, 32'hc42ec018},
  {32'hc490a1a2, 32'h449db681, 32'h445aa475},
  {32'h4353381e, 32'hc3a569ab, 32'hc4cdf969},
  {32'h432d8307, 32'h4405f06d, 32'h44324d6f},
  {32'h4576cbb8, 32'hc40cfb63, 32'h42aa93a5},
  {32'hc529f104, 32'h4389a432, 32'hc13fdd7b},
  {32'hc45daa3f, 32'hc3a3218e, 32'hc3430240},
  {32'h4259cc65, 32'h4507e093, 32'h4419eacf},
  {32'h43b041ce, 32'hc4f3d3c8, 32'hc3ca4735},
  {32'hc415556c, 32'hc45f14f2, 32'h42ddd4c3},
  {32'h438c3478, 32'h4457cccc, 32'hc432a5a9},
  {32'hc40918a8, 32'h43f12f17, 32'h43261868},
  {32'hc423bfdc, 32'hc3affd77, 32'hc3cdb649},
  {32'h44b4fb5d, 32'hc30830df, 32'hc38fa63a},
  {32'hc4dfd485, 32'h402b7bf3, 32'hc2a57454},
  {32'h446db2c4, 32'hc3e0c509, 32'h447a5e10},
  {32'h44bb8b9d, 32'h422a565e, 32'h4394e025},
  {32'h44e3a431, 32'hc362a3d7, 32'hc3799a63},
  {32'hc5071b76, 32'h4405f3bd, 32'h4364e834},
  {32'h450b96ef, 32'h43fcc331, 32'hc375fa66},
  {32'hc5652a56, 32'h43b281fa, 32'h43571107},
  {32'hc2059900, 32'hc4565b40, 32'h43a56d93},
  {32'hc3d0121d, 32'h44627a89, 32'h439955b8},
  {32'h43ef0d12, 32'hc201abbc, 32'h4537e2d8},
  {32'hc4cbcdd6, 32'hc421e613, 32'hc41a01ac},
  {32'hc492bade, 32'hc3dd8c62, 32'h42581173},
  {32'hc385d185, 32'h443a494f, 32'h448f5fbf},
  {32'h436eb2d0, 32'hc422ef26, 32'hc447c8e4},
  {32'h4490be32, 32'hc2b6d244, 32'hc2a238de},
  {32'hc21f1518, 32'h438b4b08, 32'hc54a585f},
  {32'h424114c8, 32'h435405ef, 32'h44efac6a},
  {32'hc4cbdedb, 32'hc3c35f93, 32'h41c4c570},
  {32'hc4889e36, 32'hc42c53ad, 32'h43d78461},
  {32'h44e584aa, 32'hc41f3152, 32'hc47d9b24},
  {32'h43d1b505, 32'hc36856af, 32'h443e6f3b},
  {32'h450535f6, 32'hc428f579, 32'hc3e31561},
  {32'hc3c5b94f, 32'h451b6177, 32'hc30dc355},
  {32'h44b6bd99, 32'hc1ddb47c, 32'hc427d7a7},
  {32'hc3975cdb, 32'h43bc1442, 32'h4535c820},
  {32'h450c036e, 32'hc3748698, 32'hc3e3469a},
  {32'h45314f73, 32'hc4141604, 32'h42981ffc},
  {32'hc583d5da, 32'h423040a9, 32'h4429e89f},
  {32'hc46ba8ac, 32'h4398891a, 32'hc2b4e60f},
  {32'hc4fbddf8, 32'hc4450d45, 32'hc21c4fa1},
  {32'h4409b57c, 32'h44c1421f, 32'h43e1950a},
  {32'hc460ae84, 32'hc41eb79a, 32'h43feaaf4},
  {32'hc3408bd4, 32'h44b6e6a0, 32'hc2969923},
  {32'hc4836b89, 32'hc406d98d, 32'hc40cf886},
  {32'h44a127fa, 32'h43b5e52b, 32'h43b3661b},
  {32'hc44157d6, 32'hc3be7fba, 32'h44d360ac},
  {32'h445c1aa6, 32'h438991cb, 32'hc4c2b590},
  {32'h44ee8b33, 32'hc21a5725, 32'hc2bec3b7},
  {32'h43dc02ec, 32'h4492fece, 32'h43362d14},
  {32'hc3aa3d5c, 32'hc5574491, 32'hc328de86},
  {32'h44cee6d9, 32'h41b310dc, 32'hc349a631},
  {32'hc39bd165, 32'hc328e6e6, 32'hc4cc8d52},
  {32'h43d5d624, 32'h44541fc0, 32'h4510b785},
  {32'h44566c46, 32'hc46188e9, 32'hc40cdd34},
  {32'h4442d890, 32'hc38042c9, 32'h432bcea6},
  {32'hc40bcf8e, 32'hc43e1eb3, 32'hc4a986f0},
  {32'h44b868f4, 32'h4480fb6a, 32'h4380d68c},
  {32'h439c580d, 32'hc3d19207, 32'hc52f53fa},
  {32'h451d5e6d, 32'hc38dfed2, 32'h42fcf160},
  {32'h4412ef70, 32'h4389aa06, 32'hc4a9e03b},
  {32'h44676424, 32'h448f069e, 32'h44f39431},
  {32'hc57d0fb8, 32'h438c6bbd, 32'h433fa829},
  {32'hc3be0f77, 32'h44761fc4, 32'hc3f68fe0},
  {32'h4477ff38, 32'hc37c21a8, 32'hc33483f3},
  {32'hc4303586, 32'hc4cd34bf, 32'hc38e777c},
  {32'h4495112a, 32'h44dee8a0, 32'hc388e34e},
  {32'hc3e9bea3, 32'hc3d06540, 32'h43db9a7b},
  {32'h42fe0138, 32'h451b20e5, 32'hc2e74840},
  {32'hc53257df, 32'h41615774, 32'hc2888912},
  {32'h430aa0d4, 32'h4284ae51, 32'h423e3ace},
  {32'hc56bbef8, 32'h43c469c0, 32'hc2fb861f},
  {32'h445a6c49, 32'hc1adcc18, 32'h43140f9b},
  {32'h4306e4ac, 32'hc4aa39c2, 32'h44c246d8},
  {32'h439c58bb, 32'h4484e3aa, 32'hc4bf7056},
  {32'h41a9b668, 32'hc4fd89b7, 32'h41fa095c},
  {32'hc367a99d, 32'h43b05d1d, 32'hc208f4f6},
  {32'hc32b2165, 32'hc50b604d, 32'h42d206c9},
  {32'h43a9972a, 32'h446f2ac6, 32'hc3373c9e},
  {32'h43413393, 32'hc3187abd, 32'h44c5e1b0},
  {32'h43b4f1a8, 32'hc3caf08e, 32'hc524a442},
  {32'hc43daa2c, 32'hc4668462, 32'hc2a27b3d},
  {32'h4448cb48, 32'h4398d026, 32'hc3b95b03},
  {32'hc26e4980, 32'hc5521ebf, 32'h430ab7b1},
  {32'h455b43c8, 32'h43561444, 32'hc353de57},
  {32'h442513d4, 32'hc4d42be0, 32'hc435e381},
  {32'hc30f9af0, 32'h43309bd8, 32'hc4c5dfbf},
  {32'h42d6c2d6, 32'hc55c917a, 32'h437585f3},
  {32'h451f2002, 32'h439d103e, 32'hc3bf7e2d},
  {32'hc5415b00, 32'h4379687b, 32'hc36d8ad3},
  {32'h44ef4094, 32'hc31c345e, 32'hc4a842cf},
  {32'h42b5a5c8, 32'hc5057fd7, 32'hc36a8f0f},
  {32'hc40f17ba, 32'h44ddae56, 32'h43d98279},
  {32'h4385c477, 32'hc391a62a, 32'hc39fb169},
  {32'hc31034d8, 32'h454bcc77, 32'hc2233db7},
  {32'hc3d56b05, 32'hc558d609, 32'h43afcf4b},
  {32'hc47e4eb2, 32'h420f6a2a, 32'hc384f821},
  {32'h4440dc20, 32'h4183675e, 32'h430eabd8},
  {32'h4302aec6, 32'h44af1def, 32'h44b211f3},
  {32'hc3076886, 32'h41527845, 32'h423bceab},
  {32'hc4b8e256, 32'h4461c8e9, 32'h43884c51},
  {32'h444af930, 32'hc41eb243, 32'h43e6ae75},
  {32'h44cca428, 32'hc2a76e9b, 32'h41b3c471},
  {32'h445aea57, 32'hc4031b4a, 32'h44822807},
  {32'hc3c88897, 32'h44adb887, 32'hc44006e6},
  {32'hc12533c0, 32'hc3a710e3, 32'h432c81f2},
  {32'hc3ca8e6b, 32'hc2a49f90, 32'hc4062a3d},
  {32'h42b12be0, 32'h441a4c1c, 32'h45388482},
  {32'hc40e8fca, 32'h4478c5a1, 32'h4420d3e4},
  {32'h45157eaa, 32'hc473757e, 32'hc28ed9ac},
  {32'hc4db3f98, 32'h44e1f052, 32'hc4153c56},
  {32'h44e24612, 32'h423c4008, 32'h433dc2a7},
  {32'hc51803b2, 32'h43d6dca5, 32'h43a5a43a},
  {32'h444485a4, 32'hc3930956, 32'h43d6834e},
  {32'hc4ae3d13, 32'h43d98202, 32'hc2de682c},
  {32'h432e7694, 32'h44090d72, 32'h452c804f},
  {32'hc3e0f9cf, 32'h43502d72, 32'hc437a54c},
  {32'h443ba8b4, 32'h438ba4f1, 32'h44ca97ea},
  {32'h412b81d3, 32'h420c2f8f, 32'hc4dd025e},
  {32'hc3c85f7e, 32'h4502e1e0, 32'h44e71f91},
  {32'h438c9028, 32'hc3fa3f4c, 32'hc2f9a328},
  {32'h4397bce5, 32'h42f378cc, 32'hc4364a4e},
  {32'hc311244c, 32'hc3cc76d1, 32'h441c853f},
  {32'hc3dbc498, 32'h43434156, 32'hc4d4dedd},
  {32'h42224108, 32'hc49eda26, 32'h439c2f12},
  {32'hc40ed578, 32'h45040cd1, 32'h41ded2bc},
  {32'h4485bf55, 32'hc48c2822, 32'h440a6d73},
  {32'h4523483d, 32'hc38f672f, 32'h44392d1f},
  {32'hc43c4dbb, 32'hc503f6ea, 32'hc45c30c8},
  {32'hc3a6de40, 32'hc408aa36, 32'h4397da47},
  {32'hc4b7ffb8, 32'hc3e119fc, 32'hc451da8e},
  {32'hc40f4c4c, 32'h43684464, 32'hc3d057fc},
  {32'h4111d25c, 32'hc26f9540, 32'h441039ff},
  {32'h44cef74c, 32'hc2b019c1, 32'h414841e1},
  {32'h43b6d90a, 32'hc115b51e, 32'h44e7b495},
  {32'hc2a8cf0c, 32'h44aaa122, 32'hc4885cc0},
  {32'hc4584d73, 32'h41ccc5b4, 32'hc14f3c0a},
  {32'hc51fdeb0, 32'hc1d064fe, 32'hc225e60e},
  {32'h42fa5954, 32'hc4009a48, 32'h43e2a5a5},
  {32'hc4b6549f, 32'h4305768e, 32'hc3fbd80a},
  {32'h44ba9d1e, 32'hc30caa21, 32'hc3cf9fc3},
  {32'h4286c168, 32'h4540a180, 32'hc29f4fd5},
  {32'hc418f857, 32'hc4748def, 32'hc3faa4fd},
  {32'hc3eb2302, 32'h45121724, 32'h43b3fcdb},
  {32'h4541fa23, 32'hc43b20d9, 32'hc3a27186},
  {32'hc4127cca, 32'h4345e3d8, 32'h43a85d52},
  {32'h41aed9e0, 32'h44b8ef60, 32'hc4e5efff},
  {32'hc4221699, 32'hc398743a, 32'h44acb09d},
  {32'hc1643260, 32'hc2d4d6f5, 32'h43ac2439},
  {32'h4225c7a8, 32'h42ab231b, 32'hc4d78096},
  {32'hc489a127, 32'hc3ceea01, 32'h42ca76a2},
  {32'h448011a6, 32'h437a746f, 32'hc4d81166},
  {32'hc4a8dbf3, 32'hc4a4b1c5, 32'h41f15b5a},
  {32'h4513bba9, 32'hc312553a, 32'hc3bdf46e},
  {32'h439f941b, 32'hc380388d, 32'hc4042cc9},
  {32'hc39bd038, 32'hc4c5c3d7, 32'h44cbb566},
  {32'h43c3d7b0, 32'hc482d780, 32'hc4c3dc32},
  {32'h451c18de, 32'h43aab2d6, 32'hc445a674},
  {32'hc485e892, 32'hc432958b, 32'h442440c6},
  {32'h438dcf96, 32'h42f73773, 32'hc35817e1},
  {32'hc3c069ab, 32'h41b4b01f, 32'h44ad899b},
  {32'h440e1a89, 32'h4448a562, 32'hc3d28b5c},
  {32'h44c0d0d5, 32'hc2d1f307, 32'h43ba1389},
  {32'h4570d2d4, 32'hc4043a51, 32'hc39966b3},
  {32'hc5546d17, 32'h4358791c, 32'hc41624b7},
  {32'h448421b2, 32'hc2dc3847, 32'h43e8d0fa},
  {32'hc4b3b946, 32'hc3ed81e4, 32'h41378896},
  {32'h44076729, 32'h44bed94b, 32'hc3e9fdf4},
  {32'hc4ac6a16, 32'hc3a3383b, 32'hc2a62484},
  {32'h43229118, 32'h4524c097, 32'h4170d37f},
  {32'h441599e0, 32'hc57feed7, 32'h4320637b},
  {32'h455951c2, 32'hc4693f72, 32'hc382e2d4},
  {32'h43eeac60, 32'h42d98a06, 32'h42ab5696},
  {32'h43566f92, 32'hc3582415, 32'hc4ae7526},
  {32'h43e93498, 32'h44f714aa, 32'h440c8054},
  {32'hc47c9ba7, 32'h42a40414, 32'h41df1516},
  {32'h44715024, 32'h44ae209b, 32'h440f8611},
  {32'h4389c0ec, 32'hc4fdc2ef, 32'hc46646ab},
  {32'h44f55994, 32'hc35036a7, 32'h435ffb36},
  {32'hc51095d8, 32'hc37d3c5a, 32'hc3a24428},
  {32'hc339e1dc, 32'h44a7b176, 32'h4539d545},
  {32'hc4361702, 32'h43d2c32a, 32'hc347af9e},
  {32'h433cbdcd, 32'hc3de2f2a, 32'h444824bb},
  {32'hc2f3415c, 32'hc490b475, 32'hc3eb0f64},
  {32'h44e906b7, 32'hc25461e0, 32'hc38ff43f},
  {32'hc50bce26, 32'hc3ce691c, 32'h42ba4973},
  {32'h4396997f, 32'h454fd98a, 32'hc3d45de6},
  {32'hc36f5400, 32'h426b9d83, 32'hc33a5298},
  {32'hc353664e, 32'hc2d706de, 32'h450e8c88},
  {32'hc3308533, 32'hc2ca8c36, 32'hc4c45000},
  {32'h44d1b49b, 32'hc2078e23, 32'h4379fb02},
  {32'hc4b63984, 32'hc4a48342, 32'hc3f5e0f1},
  {32'h443b7d95, 32'h4497bcf1, 32'hc2b8c840},
  {32'hc4cd168a, 32'h44132103, 32'hc3739ccf},
  {32'h44031778, 32'h4516f750, 32'h43176fe1},
  {32'hc39f2544, 32'hc4dcb24f, 32'h4284b480},
  {32'h445dcdc3, 32'hc3a15d27, 32'h43e30663},
  {32'hc5031ac0, 32'h42da951f, 32'h43500774},
  {32'h43a0b01c, 32'hc46e4201, 32'h43e201d5},
  {32'hc3b82812, 32'h4477c839, 32'hc515d241},
  {32'hc3f37404, 32'hc3e03726, 32'h44ae8452},
  {32'hc43d4927, 32'hc3a57093, 32'hc3be0ebd},
  {32'hc3aecf70, 32'h452469cb, 32'h41fa8af6},
  {32'h4427574c, 32'hc41a8a9b, 32'hc41cac76},
  {32'hc477021d, 32'h43509789, 32'h4419e411},
  {32'h4403ffe3, 32'hc4d74326, 32'hc4a86e7f},
  {32'hc571ba5e, 32'h424cb8b2, 32'h433c734f},
  {32'h4507893d, 32'h42ad529f, 32'h437ce21d},
  {32'h43830a9d, 32'hc5072b99, 32'h44fe1ae4},
  {32'h4480678c, 32'h44921174, 32'hc43adb5f},
  {32'hc43249b1, 32'hc3763706, 32'hc17144c6},
  {32'hc277b050, 32'hc4838a3d, 32'hc4a3fc8f},
  {32'hc3778508, 32'hc2baddc1, 32'h449f6ec0},
  {32'hc4713c01, 32'hc2bcda54, 32'hc3ba3e69},
  {32'hc49fa467, 32'h44089037, 32'h4454f75a},
  {32'h42814207, 32'hc3a871d5, 32'hc42d7085},
  {32'h433c3656, 32'h43883e8a, 32'h44ad343b},
  {32'h4522856c, 32'hc43fa0de, 32'h40ef2fc8},
  {32'h4352031f, 32'h45670c7e, 32'h42d00f6f},
  {32'h44e73fd2, 32'h438482bb, 32'hc0b50140},
  {32'hc3c991c6, 32'h4533ab57, 32'h43cf205f},
  {32'h4438bf50, 32'hc49ee90e, 32'h440ec68d},
  {32'hc4e5e054, 32'hc400834c, 32'h429c271a},
  {32'h4410dbf8, 32'h430830a6, 32'h437a4770},
  {32'hc54c9310, 32'hc3e3a7e0, 32'hc3905928},
  {32'hc4c22da7, 32'h42bab986, 32'hc3dd8942},
  {32'h43f41c60, 32'hc15a19d9, 32'hc3a7c3c8},
  {32'hc51438b6, 32'h441de05f, 32'hc3883a83},
  {32'h44caafc0, 32'h430571c1, 32'h449c6104},
  {32'hc4c6ef2b, 32'h3f29da00, 32'hc42aedce},
  {32'h444e7cd8, 32'hc44fd9df, 32'h429a89c7},
  {32'hc5113695, 32'h440e23c9, 32'h420418d8},
  {32'h4546cf1b, 32'h444141bb, 32'hc3518e30},
  {32'hc4f12a05, 32'h4426e2ec, 32'h441fc07a},
  {32'hc30c6eb0, 32'hc504886f, 32'h431230ca},
  {32'hc4b17675, 32'hc1d30dd4, 32'hc28aaaeb},
  {32'h444f5313, 32'hc38712e6, 32'h448a8d64},
  {32'hc3d67b3c, 32'h4280e917, 32'h43cfd35e},
  {32'hc30b42fa, 32'hc459fa94, 32'hc4440be6},
  {32'h43889a05, 32'h44b9055c, 32'h443b6b44},
  {32'h440cd58a, 32'hc33e9f36, 32'hc4603183},
  {32'h4489d830, 32'h42d88039, 32'h436685ac},
  {32'h43f6e055, 32'hc3d37702, 32'hc4fc6918},
  {32'hc2983ba8, 32'hc3be347d, 32'h4510d301},
  {32'h44cdc5c6, 32'hc3d2d9aa, 32'hc191255a},
  {32'hc4b9da65, 32'hc0df98ed, 32'h43d6af80},
  {32'h44edb1c1, 32'h440a5468, 32'hc3e6dfb5},
  {32'h43bb2163, 32'h43c45270, 32'h44c4eda4},
  {32'hc34d2514, 32'hc45de76a, 32'hc4b3910f},
  {32'h42df46e4, 32'h454fac2b, 32'h43376ca0},
  {32'h44ee0801, 32'h418a920c, 32'hc33677de},
  {32'h4256daa0, 32'h44991e07, 32'h44ada51a},
  {32'h43d926a8, 32'hc5067836, 32'hc416da51},
  {32'h4463abce, 32'hc3a57b8b, 32'hc4878da9},
  {32'hc54af908, 32'hc2677e9d, 32'h44712870},
  {32'h45078d35, 32'h4317bd73, 32'h42335ead},
  {32'hc38d6c90, 32'hc43e45a4, 32'h43b479ff},
  {32'h44113efa, 32'h44f37823, 32'h42b31a3b},
  {32'hc51cf9a0, 32'hc3b56f78, 32'hc2d5455b},
  {32'hc32820f5, 32'h458a2ac0, 32'h43dbe1d8},
  {32'hc3968b78, 32'hc48b363e, 32'hc40fd4bb},
  {32'h444bf70d, 32'h447a6546, 32'hc29c13cb},
  {32'hc4d566a5, 32'hc3423b08, 32'h42d785db},
  {32'h450c3182, 32'h42ee1c6e, 32'hc40ae1c5},
  {32'h4374f3d0, 32'hc3b1908d, 32'h44bd34a3},
  {32'h44077c3a, 32'h44910f63, 32'h435f9abb},
  {32'hc4d986dc, 32'hc48069ca, 32'hc3a647a6},
  {32'h429aaed7, 32'h44b1bfb3, 32'h43cd2c58},
  {32'hc29ddd18, 32'hc416b370, 32'hc501b751},
  {32'h439bb124, 32'h43ef1aaf, 32'h454b371f},
  {32'h44018439, 32'hc4aafd2e, 32'hc380917f},
  {32'h44f2601e, 32'h433d99f8, 32'h447009ae},
  {32'hc3bd8240, 32'h445f7e3c, 32'hc4aa1bf8},
  {32'hc4c29523, 32'h43790cb7, 32'hc3745fc6},
  {32'hc54d367d, 32'h438a33e8, 32'hc303d9ce},
  {32'h43e69735, 32'h4473c8ca, 32'hc1b2a6e8},
  {32'hc47874c0, 32'hc41e5e17, 32'hc3ea4281},
  {32'h44e49fe8, 32'h441cb6bf, 32'h446f58eb},
  {32'hc4d63944, 32'hc3fad817, 32'hc4a915b6},
  {32'h44866660, 32'h439f7602, 32'h44146957},
  {32'h4514ea47, 32'hc442e9bc, 32'hc357d096},
  {32'hc4bee2c3, 32'hc3bd1ced, 32'h43224851},
  {32'h446e1563, 32'h44f3b03b, 32'h439abb5c},
  {32'hc36e059c, 32'hc2e35139, 32'hc359b47b},
  {32'h4423104d, 32'h4498c5ee, 32'h441ed58d},
  {32'hc5218765, 32'hc3527b5b, 32'hc1bd83d3},
  {32'h44c3312d, 32'h43d0051a, 32'hc30ba7f6},
  {32'hc4d72108, 32'hc2cd0efa, 32'hc32b2378},
  {32'hc24aa480, 32'hc461774a, 32'hc30942df},
  {32'h441afa38, 32'hc4327201, 32'h423124b0},
  {32'h430dd638, 32'h44963da0, 32'hc4ba3bcf},
  {32'hc34b8f94, 32'hc4b95f34, 32'h43e6eb37},
  {32'hc446c445, 32'h42d066d7, 32'hc3f6a437},
  {32'hc008a440, 32'hc5059008, 32'h42f35afd},
  {32'h448fcbf6, 32'h40b43e88, 32'hc3b1f058},
  {32'hc3d14f3c, 32'h438df640, 32'h4361563b},
  {32'h445230d5, 32'hc3a1fff3, 32'hc4faa68c},
  {32'hc546a27b, 32'hc2edcf74, 32'h43836809},
  {32'h43834f51, 32'h44c37875, 32'hc2e119c8},
  {32'hc404be2a, 32'hc49c187c, 32'h450dcbbf},
  {32'h44b3056d, 32'h4471d140, 32'hc4f672a9},
  {32'h42c7847c, 32'hc4899f31, 32'hc3feb6e9},
  {32'h4321bd68, 32'h445d5e6c, 32'hc422c0ba},
  {32'hc2cb5ca0, 32'hc5056343, 32'h43b6d0f3},
  {32'hc4b7ba5b, 32'hc12a0b1b, 32'hc31da89e},
  {32'hc48755f5, 32'hc223853e, 32'h43e2b226},
  {32'h4459a49e, 32'hc3b551ca, 32'hc520ed8b},
  {32'h44e06fa6, 32'hc43a7c3f, 32'hc411f482},
  {32'hc4108e33, 32'h443ddbb3, 32'h3fcca482},
  {32'h42a4f13c, 32'hc4407fff, 32'h43a1f226},
  {32'hc31c8d74, 32'h453e7ac9, 32'hc3c50559},
  {32'h453d63de, 32'h42ef8877, 32'hc3bb330f},
  {32'hc4510a40, 32'h4389599d, 32'h4336136d},
  {32'h44358842, 32'hc4c863fb, 32'hc4bde0b2},
  {32'hc44a632a, 32'hc3facbe4, 32'h434b41e7},
  {32'h44bfb732, 32'h4278a423, 32'h445f0d5d},
  {32'hc4b9e2e9, 32'h447cd3f0, 32'h438baf14},
  {32'h433c9c00, 32'hc4189264, 32'h450cadb6},
  {32'hc50943a4, 32'h4269e589, 32'hc364b183},
  {32'h43c26902, 32'h42b59907, 32'h44bac7ff},
  {32'hc4822403, 32'h43c5405d, 32'hc3a8639b},
  {32'hc49e3106, 32'hc31f9f2d, 32'hc3608242},
  {32'hc498e3cb, 32'h44007a49, 32'h42eafabe},
  {32'h428392ec, 32'h4398e0ac, 32'hc42e4136},
  {32'h44c58865, 32'h4273531f, 32'h43ad2ad4},
  {32'h436795b0, 32'hc4963f58, 32'h44afc976},
  {32'hc42e0448, 32'h452654af, 32'hc2c27ed1},
  {32'h44997ad2, 32'hc2f62de4, 32'hc326e09d},
  {32'hc3c2c5b8, 32'h44b7b7fc, 32'hc2ac3e94},
  {32'h441996a6, 32'hc3ca38e3, 32'h4491208d},
  {32'hc5458734, 32'hc302bb82, 32'h4392b788},
  {32'h44855a3c, 32'h435bacae, 32'h4417d7af},
  {32'hc4ae179f, 32'hc342f1f8, 32'hc50d1a70},
  {32'h440bd22f, 32'hc3a4b14a, 32'h4211cc2e},
  {32'hc41b95b3, 32'hc4d3183c, 32'hc47d1c9d},
  {32'hc370d65c, 32'h448814a3, 32'h452a5d3f},
  {32'h43704dc0, 32'h4477efbe, 32'hc4260b68},
  {32'hc4dfd771, 32'hc366fee3, 32'hc1989bb3},
  {32'h42e6f630, 32'hc330131e, 32'h4544fb07},
  {32'hc3ed4f72, 32'h44eeff03, 32'h442b504c},
  {32'h432b47bc, 32'hc42df8a2, 32'h439aed4b},
  {32'hc40b461a, 32'h452fb569, 32'hc19e15b2},
  {32'h431d24c0, 32'hc4d1396c, 32'h43e64b22},
  {32'hc34f033e, 32'h43d4b794, 32'h4390be82},
  {32'hc50c5ece, 32'h4409c1aa, 32'hc42e65f6},
  {32'h45001cb9, 32'h43823123, 32'hc3f4d3fe},
  {32'hc4fce1bc, 32'h43ec3ecd, 32'h40e5f3dd},
  {32'hc451c171, 32'hc33c47b4, 32'hc4f98565},
  {32'hc3983c3b, 32'hc30327b9, 32'h453b8d99},
  {32'h43d25c68, 32'h44ecdbe0, 32'h4337487d},
  {32'hc2ac8257, 32'h4402fd8a, 32'h45398018},
  {32'hc25af160, 32'hc38107c3, 32'hc5313acf},
  {32'h45181477, 32'hc41f041c, 32'h4318da00},
  {32'hc53e9483, 32'hc3ff33c3, 32'hc41f8ccf},
  {32'h44ec34be, 32'h432dfe4c, 32'h448e4c66},
  {32'h43a5228c, 32'h44401ce5, 32'hc419ded9},
  {32'h448a8718, 32'hc401a877, 32'hc3849d1e},
  {32'hc53013ac, 32'h42d617ba, 32'h439f4246},
  {32'h4348bd66, 32'hc4b3a631, 32'hc3a82bd4},
  {32'hc4cb9e64, 32'h44afe232, 32'hc2a1d2cd},
  {32'h4423fa80, 32'hc43aa35e, 32'h439cd37f},
  {32'hc4c74f6b, 32'h436f7b2d, 32'hc20a64f8},
  {32'h44b81c36, 32'h44997498, 32'hc42a2628},
  {32'h437b36d5, 32'h43e48df7, 32'h452a9365},
  {32'hc3bd1b4b, 32'hc483874f, 32'h444c69a3},
  {32'h4395d550, 32'h44db9cec, 32'hc3d2bd62},
  {32'h44e800b4, 32'hc3eb218c, 32'hc2c028e5},
  {32'h43c0270c, 32'hc31cf9d0, 32'hc535408b},
  {32'hc3aa684e, 32'hc2a81f67, 32'h45010a66},
  {32'hc42e8a37, 32'h443d9dc8, 32'h42ac9d2e},
  {32'h43cd4515, 32'h44bd4094, 32'hc479e917},
  {32'hc4cf3a54, 32'h43f75ba0, 32'h4473c22c},
  {32'hc3966989, 32'h449ad081, 32'hc5106191},
  {32'h41274241, 32'h45027579, 32'h43cae3eb},
  {32'hc406dea4, 32'hc518961c, 32'h41eaab2a},
  {32'hc34eee70, 32'h432c8d90, 32'hc3bbf480},
  {32'hc381d235, 32'hc5479511, 32'hc40d2641},
  {32'h4421a999, 32'hc1999ca6, 32'hc3b6be73},
  {32'hc3f2ecc3, 32'h4303fdc2, 32'h4330e958},
  {32'h4510f4f7, 32'h43c1d1c3, 32'hc23dc399},
  {32'hc4642a39, 32'h434b4927, 32'hc3bb7af8},
  {32'hc3569caa, 32'h4407c986, 32'hc314a076},
  {32'hc3761708, 32'hc4e2671b, 32'h42c954a9},
  {32'h4189e460, 32'h45412a32, 32'h4287f3f4},
  {32'hc4e8bf7d, 32'hc331deff, 32'h43e60199},
  {32'h448c9376, 32'h44feedb4, 32'hc35cc275},
  {32'hc4a263e0, 32'hc4ccb586, 32'h424064f3},
  {32'h451dcc3a, 32'hc37648a7, 32'hc2ac19c2},
  {32'h44791636, 32'hc4cdd828, 32'h43d4024d},
  {32'hc20634d0, 32'h4508b518, 32'hc4830364},
  {32'h4169aba4, 32'hc4ce74d4, 32'h44728bef},
  {32'h43fe946e, 32'hc415fad3, 32'hc17d4cbc},
  {32'h440c5ed9, 32'h44a87f6c, 32'h4495f085},
  {32'hc3717fb0, 32'hc3d89cd3, 32'hc462beb8},
  {32'h43db6f84, 32'h44acb54b, 32'h43637345},
  {32'h43a06d3c, 32'hc45eb3ac, 32'hc51ebdf1},
  {32'h44144f27, 32'h44b6c81a, 32'h44b96e3a},
  {32'h446ec3d3, 32'hc3078f5b, 32'hc23a35ed},
  {32'hc43ac389, 32'hc2be6adb, 32'h43987e28},
  {32'hc456df69, 32'h446efb12, 32'hc49c15f3},
  {32'hc49dbb72, 32'h4399c4d8, 32'h43419c78},
  {32'hc3c1dded, 32'hc3cb6b05, 32'hc4d676dd},
  {32'h44e14d5d, 32'h43834cd7, 32'h438c071a},
  {32'h44a5047e, 32'hc4204690, 32'hc3f136d6},
  {32'h4321ec52, 32'h44184f91, 32'h45275ed9},
  {32'hc4e32678, 32'hc301d38c, 32'hc3c85006},
  {32'h433f70cb, 32'h4483c4c8, 32'h430eb3b0},
  {32'hc495f7e6, 32'hc4a32378, 32'hc22b5c0a},
  {32'h4510409e, 32'h44710539, 32'h42de03ee},
  {32'h441ff4c9, 32'hc2ee6d0a, 32'hc3a38151},
  {32'h4522fa3e, 32'hc37105fa, 32'h43471026},
  {32'hc3c877e7, 32'hc53410d2, 32'h43786880},
  {32'h443a4430, 32'h433e0abe, 32'h4409a502},
  {32'hc58262b7, 32'hc25cb29e, 32'hc2c0cd6f},
  {32'h4502847f, 32'h433ac2d5, 32'h4127a8f1},
  {32'hc378b7a2, 32'h4407767c, 32'hc3f6d88e},
  {32'hc31030d4, 32'h449bf358, 32'h43fb019d},
  {32'h4112d3c0, 32'h434589e1, 32'hc44b1ca2},
  {32'hc4fe1011, 32'h43fc00f9, 32'h4299ea89},
  {32'hc1e7f208, 32'hc4db9298, 32'hc38d3764},
  {32'hc3fa8856, 32'h4461b778, 32'h44258454},
  {32'h44d92799, 32'hc264772d, 32'hc488ff90},
  {32'hc3770c40, 32'h447eb912, 32'h449b3c41},
  {32'hc290fc10, 32'hc22da41c, 32'hc416225a},
  {32'h439471a4, 32'hc513498b, 32'h44f68064},
  {32'hc42d425f, 32'h445d4f94, 32'hc4061848},
  {32'h44a105cd, 32'h4328d1ad, 32'h4346b726},
  {32'h44d3213c, 32'h4363e628, 32'hc43ca5e0},
  {32'hc4021982, 32'h43950d3a, 32'h44db2de4},
  {32'h44ed0438, 32'hc38a9f63, 32'hc30bea6d},
  {32'hc478b8c2, 32'hc3acfd38, 32'h43ae1053},
  {32'hc3a5e990, 32'hc4a993c9, 32'hc4ba5e3a},
  {32'hc4542d60, 32'hc2853fea, 32'h434bfc0a},
  {32'h4418aa70, 32'hc4528c6f, 32'hc43efbc3},
  {32'hc4929bc8, 32'h44c69228, 32'hc22531cd},
  {32'h440b3972, 32'hc48ad7ea, 32'hc36aa224},
  {32'hc4823202, 32'h451688bd, 32'h41aed38c},
  {32'h43b04dfb, 32'hc56b2227, 32'hc355234a},
  {32'h431e23a8, 32'h44aaeb67, 32'h43927fc8},
  {32'h456af9d9, 32'h43d29c21, 32'hc2afd2bb},
  {32'hc527b467, 32'h443bbc4d, 32'hc3a7bc7f},
  {32'hc3e3137e, 32'hc3920bb2, 32'hc15e4c2a},
  {32'h41d0efe0, 32'hc36dd72e, 32'hc38f4772},
  {32'hc472c97a, 32'hc3d30860, 32'hc438ef2e},
  {32'h4504b793, 32'h42b6f9fc, 32'h44763d61},
  {32'hc30e17b0, 32'h409098e2, 32'hc388349b},
  {32'h42cb13b4, 32'hc4e9ad6d, 32'h427950b2},
  {32'hc52a955b, 32'h43f83e13, 32'h441af3e0},
  {32'h41867ec0, 32'hc4908df4, 32'hc2d475de},
  {32'hc3377437, 32'h45621351, 32'hc388285f},
  {32'h4505274a, 32'hc39dbf04, 32'h43b4ff1c},
  {32'h450d0667, 32'hc3de7ed5, 32'h41dd4a8e},
  {32'h43f08012, 32'h4395b37d, 32'h4355b6e2},
  {32'hc483950d, 32'h43bd713a, 32'hc4c1fdae},
  {32'h444abf5c, 32'hc3e2befa, 32'hc45c56f6},
  {32'hc470261c, 32'h435532d6, 32'h443cf8b6},
  {32'h437f887c, 32'hc4764d3f, 32'h3ffea464},
  {32'hc2b9c3e8, 32'h44ed6dbb, 32'h44163c62},
  {32'hc3971e5e, 32'hc3168540, 32'h4158ce86},
  {32'h435696db, 32'h450de9fa, 32'h438539d0},
  {32'h44e9671e, 32'h42a1c4ac, 32'hc43d80e2},
  {32'hc3a11f90, 32'h443a87e1, 32'h44e9c843},
  {32'hc24490f0, 32'hc1abe9bb, 32'hc3d38f21},
  {32'hc391e843, 32'h44c01367, 32'hc3c7300e},
  {32'h449d6133, 32'hc4321c7d, 32'hc3b10772},
  {32'hc2f56c56, 32'h4495a82d, 32'h4512287e},
  {32'h43f569e6, 32'hc49152c0, 32'hc153fc30},
  {32'hc4af048e, 32'h42d9eb5e, 32'h4494652d},
  {32'h44626a43, 32'hc4d46af2, 32'hc403478c},
  {32'h4515bf94, 32'hc3b6e6a8, 32'hc44093ca},
  {32'hc505afd4, 32'hc1285b92, 32'h42a39c4c},
  {32'hc3891698, 32'h430ba2f6, 32'h42cfe24e},
  {32'hc37497d0, 32'hc4dd9167, 32'hc3b1de5a},
  {32'h4281ee68, 32'h4501a2ce, 32'h43660cf4},
  {32'hc53a4188, 32'h42cc6dfd, 32'hc354090a},
  {32'h454a1898, 32'h43faa9dc, 32'hc23178ea},
  {32'hc3dcdd68, 32'hc513fc9c, 32'h4399525f},
  {32'h4438f922, 32'h42d186de, 32'h4368c77b},
  {32'h4325cdc0, 32'h439cc12f, 32'h4330a2ca},
  {32'h4313a45f, 32'h43abd244, 32'hc5296b92},
  {32'hc47f3732, 32'hc23e3611, 32'h42ccc9c5},
  {32'h4364ccf0, 32'h44978959, 32'h44046635},
  {32'hc4cca2d6, 32'hc3f994fe, 32'hc43e390c},
  {32'hc371260a, 32'h42b839d6, 32'h44baead3},
  {32'hc5241ee7, 32'hc3053646, 32'hc468e6fb},
  {32'h44c67600, 32'h440e1142, 32'h444c763a},
  {32'hc464b1fe, 32'hc404fc7d, 32'h43c1e4ac},
  {32'h447af5a0, 32'h44055b14, 32'h440c1ea4},
  {32'hc583e34c, 32'h4365095e, 32'hc325d7f7},
  {32'h45393be8, 32'h42da57dc, 32'hc427ac4d},
  {32'hc47902ff, 32'hc3b36c9d, 32'hc483000f},
  {32'h44b5e5f1, 32'h422d7604, 32'h4346e8ad},
  {32'hc3194d24, 32'hc3bbc2e2, 32'hc4319826},
  {32'h44ccb566, 32'h436971cf, 32'h4438d9a9},
  {32'hc4489b24, 32'hc48d5d48, 32'hc4e33924},
  {32'h44fb76f0, 32'h435512d5, 32'hc394fcfb},
  {32'h445315bc, 32'hc233269a, 32'hc3832f4e},
  {32'hc51293f0, 32'hc3a6a636, 32'h44032e94},
  {32'h43b7177c, 32'h443689ce, 32'h448f2411},
  {32'hc3432085, 32'hc4dc3989, 32'h43b16a5f},
  {32'h451b665d, 32'hc387a636, 32'hc37944c8},
  {32'hc4b078a5, 32'hc419fc3d, 32'hc084525c},
  {32'h44bca856, 32'h433db8dd, 32'hc3d4fd03},
  {32'hc5310c28, 32'h42b44308, 32'hc408820f},
  {32'h43581268, 32'h44964d9b, 32'h44659489},
  {32'hc395da06, 32'hc49abcb5, 32'hc14f24fc},
  {32'h43205880, 32'h44970aa7, 32'hc3aee6c0},
  {32'hc48142d6, 32'hc34af811, 32'hc3e990fd},
  {32'h447f24fe, 32'h442a38e4, 32'h430d0b50},
  {32'hc473ac8e, 32'hc364452e, 32'h448647fd},
  {32'h44949962, 32'h42a4557d, 32'hc30384fa},
  {32'hc4d5c74c, 32'hc2c27843, 32'hc29ef040},
  {32'h4436c604, 32'h43ee343a, 32'hc2b7654c},
  {32'hc32b24a4, 32'h43e9a0b1, 32'h4535ee43},
  {32'h443c2ddb, 32'hc3e975b4, 32'h42e1c734},
  {32'hc420b700, 32'hc51642c1, 32'h44070f30},
  {32'h41a26573, 32'h442cb8ee, 32'hc4a3e635},
  {32'h449cb400, 32'hc449e6ae, 32'h4294c427},
  {32'h4484dbde, 32'h444d764b, 32'hc49621c9},
  {32'hc483792e, 32'hc445eec8, 32'h43d84436},
  {32'h446bd29d, 32'hc36b9ea2, 32'hc4a45786},
  {32'hc549df14, 32'hc3f2cddc, 32'h435645f2},
  {32'h44bc8ddc, 32'h43740197, 32'hc43aafb8},
  {32'h43bbb594, 32'hc459aed0, 32'hc41a5c8f},
  {32'hc4ba3eaf, 32'hc2daa0e5, 32'h442f147b},
  {32'h43df08b1, 32'h434a172c, 32'h43b8f6d5},
  {32'hc4a0a390, 32'h438bec5f, 32'h42750c5b},
  {32'h436117b0, 32'hc41904c8, 32'hc3b027cd},
  {32'hc4b686a4, 32'h4220bfdb, 32'hc3a3272a},
  {32'h43e4364a, 32'h438890c5, 32'hc43a8255},
  {32'hc500ce34, 32'hc3039069, 32'h43a0e957},
  {32'h4539669c, 32'hc3e2ff58, 32'h43e379dc},
  {32'h435e1f74, 32'h44122015, 32'hc4394a64},
  {32'h4446ba06, 32'h4489f116, 32'hc496e6b9},
  {32'hc4ee2838, 32'hc2fe559e, 32'hc3107cff},
  {32'h44a95524, 32'hc48ac59e, 32'h44422823},
  {32'hc42fa7af, 32'h44243e9e, 32'h43873102},
  {32'hc4ba0f12, 32'hc28fc424, 32'h43167721},
  {32'hc4939cbf, 32'hc317abf1, 32'hc4b35a2e},
  {32'h439ee2d0, 32'hc37e9b9e, 32'hc11c22db},
  {32'h448b04e6, 32'hc3b28bbe, 32'hc3f0f9a7},
  {32'h43737fb0, 32'hc5024be3, 32'h43628a18},
  {32'hc5532969, 32'h43c69bf7, 32'hc36097ee},
  {32'h41acccb0, 32'h435294d6, 32'hc2f2c9d0},
  {32'hc51437f3, 32'h44753ae5, 32'hc3135299},
  {32'h45622c48, 32'h444d029f, 32'hc3f4c122},
  {32'h4366acc6, 32'h4426248e, 32'hc3534400},
  {32'h453d7083, 32'h43e6a787, 32'h43a15d27},
  {32'hc52305eb, 32'hc29f111b, 32'hc4a4cdb8},
  {32'h457300c1, 32'h432edbaf, 32'hc3941382},
  {32'hc1e597a0, 32'h449705f7, 32'hc487e67b},
  {32'h448f7c25, 32'h43cb9564, 32'h44050471},
  {32'h44045ef6, 32'h42991766, 32'h4457582b},
  {32'h43d726c6, 32'h425fec36, 32'hc4c50b4c},
  {32'h44141402, 32'hc43d5e3b, 32'h44e6fc1c},
  {32'hc3330df2, 32'h449623dd, 32'hc41ce4fa},
  {32'h45012d32, 32'h43389b2f, 32'h42dc923f},
  {32'hc42585ae, 32'h4505df28, 32'h43ea8fea},
  {32'h4249297a, 32'hc405bcb8, 32'h44fe390e},
  {32'h44d537e5, 32'hc1bac214, 32'h445ae60c},
  {32'hc4228913, 32'hc4a55990, 32'hc4b51c66},
  {32'hc4546714, 32'hc4908876, 32'h44035798},
  {32'h429adb50, 32'hc390686a, 32'h449a6734},
  {32'hc37d7f1b, 32'hc3d6cb78, 32'hc530f417},
  {32'h4443e92a, 32'hc3b9a9e4, 32'h447a2416},
  {32'h44840630, 32'h445c1b2a, 32'hc1e5f1e7},
  {32'h44c61598, 32'h4079c411, 32'h43c04a7b},
  {32'hc31a36dc, 32'h42552864, 32'hc46a67c8},
  {32'h44bf04e2, 32'hc3f9d63d, 32'h4231dfea},
  {32'hc4e05240, 32'hc3a5fa78, 32'hc3897fba},
  {32'h4551f2c4, 32'h428fe04e, 32'hc46104d3},
  {32'hc53a4be1, 32'hc4091d6e, 32'h432ef902},
  {32'hc36672b0, 32'hc5271115, 32'hc3145c65},
  {32'hc4428b65, 32'h452d3424, 32'hc2f98cb4},
  {32'h45211864, 32'hc3fb8162, 32'hc356ec37},
  {32'hc3381908, 32'h4516a678, 32'h429aa3f9},
  {32'h438be9d4, 32'hc5238b15, 32'hc31df2b7},
  {32'h4462229b, 32'hc3276ac2, 32'h44736750},
  {32'h43196d36, 32'hc4027b99, 32'hc4b11828},
  {32'h4407cedc, 32'hc3832b92, 32'h452bf3d8},
  {32'hc466dba8, 32'h4412df06, 32'h44c4b92a},
  {32'hc396d820, 32'hc3526150, 32'hc51ed1fa},
  {32'hc4fb59aa, 32'h4206c85e, 32'h42c522f4},
  {32'hc1b14328, 32'h45676333, 32'hc3811ea8},
  {32'hc2a348bc, 32'hc4a7db26, 32'h4419262c},
  {32'h44194701, 32'h4367c594, 32'h43415109},
  {32'h41ce61f0, 32'hc433dc55, 32'hc3d8bb54},
  {32'hc3f2f2ec, 32'hc5020e40, 32'h44abf44c},
  {32'hc35f3bed, 32'h444919d6, 32'hc4e69d79},
  {32'h44cdc5ac, 32'h446aa635, 32'hc375e09d},
  {32'hc37bb33a, 32'hc412abd2, 32'h44a6c45a},
  {32'h443918ea, 32'h3d699320, 32'hc43ee43e},
  {32'hc3ee93c0, 32'hc2ab7bea, 32'h44edd964},
  {32'hc18835a0, 32'h44ed75fb, 32'hc30af07d},
  {32'h4412c3f7, 32'hc1f2c24c, 32'h447d8de8},
  {32'h43161700, 32'hc460e253, 32'hc417d844},
  {32'hc50b601e, 32'hc38ba6ee, 32'h433970c2},
  {32'h431e4a89, 32'h4422ef89, 32'hc3d1d5ba},
  {32'h4226afa8, 32'hc50921d1, 32'hc34c0baf},
  {32'h42c63854, 32'h4566a0b8, 32'h43dd2950},
  {32'h43f5c9e0, 32'hc4653396, 32'h43a275dc},
  {32'h449315a6, 32'h44caf8de, 32'hc3538424},
  {32'hc4eb1116, 32'hc4a98cf1, 32'h434a47fb},
  {32'h44e37565, 32'hc3f370eb, 32'hc1a42088},
  {32'h430e8064, 32'hc2ff0898, 32'h43cf3174},
  {32'hc31aafb6, 32'hc4c5bb68, 32'hc3c58ca4},
  {32'hc25588ba, 32'hc33c2f38, 32'h44a24983},
  {32'h437354e0, 32'h417bebe1, 32'hc4a15835},
  {32'h43cdf62d, 32'hc3a9a9c0, 32'h4247ef14},
  {32'hc2dc9538, 32'hc4f25de1, 32'h429899c7},
  {32'h44263110, 32'h42a0ed1f, 32'h44054176},
  {32'hc4406c7c, 32'hc32691fc, 32'hc496a9ba},
  {32'hc3279790, 32'h4334e7cb, 32'h446ba29a},
  {32'h44ab53ad, 32'hc385e5e0, 32'hc3b026b1},
  {32'h443e48ff, 32'h4412613a, 32'h432651d2},
  {32'hc507c7f8, 32'h41e52516, 32'hc3d737cd},
  {32'hc3357a0c, 32'h4492f159, 32'hc299c6fd},
  {32'h43d9b39f, 32'hc49b9f53, 32'h42773548},
  {32'h449edfba, 32'h448011c4, 32'h417b54cf},
  {32'hc47a7fc2, 32'hc3bb8d1c, 32'hc40fa63a},
  {32'h42fe3ef0, 32'h44ab551b, 32'h44cccda9},
  {32'h43fe440f, 32'hc3ac1bf2, 32'hc526dedf},
  {32'h4551eedd, 32'hc374b07a, 32'hc132762a},
  {32'hc4996b43, 32'hc4bf673d, 32'hc4053cbd},
  {32'h450ae1cd, 32'h445287bb, 32'h4320747c},
  {32'h444cf522, 32'hc4dd9771, 32'h432b330b},
  {32'hc3a8f7fc, 32'h4587b006, 32'hc380f5ce},
  {32'hc47dd2ad, 32'hc4f8fd8a, 32'h4392f681},
  {32'hc41f2a58, 32'h439bf8e7, 32'h428e1039},
  {32'hc52ba3a8, 32'h43f1c84b, 32'hc409dfea},
  {32'h457b8214, 32'hc220ef2a, 32'h420a4c37},
  {32'h44835571, 32'hc31d2ec1, 32'hc2d067e1},
  {32'hc38344a2, 32'h4450051e, 32'h436a1192},
  {32'hc397e20f, 32'hc49ebd76, 32'hc3ad8fa5},
  {32'hc45c7002, 32'h451c67a8, 32'h43b470d6},
  {32'h433e5e2c, 32'hc44f427b, 32'hc4e51207},
  {32'hc391e380, 32'h44a65ca1, 32'h431e46e9},
  {32'h44ae7bf3, 32'hc3ba72ec, 32'hc491b790},
  {32'hc4deefd4, 32'h43a3b82e, 32'h442043cc},
  {32'h43d6cebe, 32'hc3af94ed, 32'hc4888e99},
  {32'h441ae68d, 32'hc47950ff, 32'h450341fe},
  {32'hc3cce66f, 32'hc540b983, 32'hc4519ee4},
  {32'h443aaaa5, 32'hc3df3d85, 32'h43f5a221},
  {32'hc34639b6, 32'hc434031a, 32'hc47c1c8d},
  {32'hc480f9c4, 32'h4504408f, 32'h43b27d2e},
  {32'h43ad2c15, 32'h43c9ea8a, 32'hc48d4b7b},
  {32'hc46db381, 32'h42285e0f, 32'h44393a66},
  {32'h445ceb2f, 32'h43c8fc92, 32'hc4a08148},
  {32'h443f6f34, 32'h43b43004, 32'h445c3569},
  {32'h4318d030, 32'hc5256422, 32'hc4073f9c},
  {32'hc43e43e7, 32'h45190799, 32'h42c11cfc},
  {32'h4541512f, 32'h42918b67, 32'hc3ed5145},
  {32'hc422abe0, 32'h4510c6e2, 32'hc2b5b818},
  {32'h453e5fdb, 32'hc3dd47e7, 32'hc36146b2},
  {32'h43c58b8c, 32'hc414cca7, 32'hc2d68819},
  {32'h445b40a0, 32'h4395f2b9, 32'hc4039361},
  {32'hc4e85f44, 32'h42832e4b, 32'hc4057994},
  {32'h430b431c, 32'h42434fa6, 32'hc3b0acb4},
  {32'h437b2af4, 32'h42c97e97, 32'hc308dba7},
  {32'hc561118e, 32'hc314eb9d, 32'h42cab888},
  {32'hc3fbfc00, 32'hc3962fac, 32'h442d2521},
  {32'h44e0fcfe, 32'h42ab6b9c, 32'h42f0701e},
  {32'h45368682, 32'h43a4b16e, 32'hc28272b9},
  {32'hc4628b50, 32'h448e186d, 32'hc2b720b3},
  {32'hc3318d7d, 32'hc4e48031, 32'h424aa625},
  {32'hc438a97d, 32'h451901ab, 32'h439fc3b6},
  {32'h447a7972, 32'hc4a1cd48, 32'hc3137043},
  {32'h4424c32a, 32'h4420571f, 32'hc4af5c1e},
  {32'h451f2784, 32'h4202ef36, 32'h43b1f661},
  {32'hc51cd404, 32'h437adce7, 32'h424bde6e},
  {32'h44d6cf63, 32'h415d70ce, 32'h438c2b6b},
  {32'hc3f67e66, 32'h43c76b3e, 32'h432349c4},
  {32'h443e357c, 32'hc442042c, 32'hc4420e45},
  {32'hc530cc16, 32'hc30621a3, 32'h43800131},
  {32'h4468babf, 32'h42831060, 32'hc4c6a0fc},
  {32'hc49e4582, 32'hc1da7d9a, 32'h446c3d39},
  {32'h456dd194, 32'hc3c237c8, 32'h436eb6e6},
  {32'hc529727e, 32'hc425abca, 32'h4347a95b},
  {32'h44dde997, 32'hc3ed2b99, 32'hc485082f},
  {32'h433b9378, 32'h43bf409a, 32'h44f4b03b},
  {32'h4481c486, 32'hc29b7443, 32'hc41035ec},
  {32'hc2fe8e60, 32'h42fdb026, 32'h441c4d4b},
  {32'h453b853a, 32'hc3868f3f, 32'h42c19d7f},
  {32'hc5666ef2, 32'h435324cc, 32'h44322e6c},
  {32'h44b5dc44, 32'hc49dc202, 32'hc40c7690},
  {32'h4533ad37, 32'h42dbd78b, 32'hc27fffc0},
  {32'hc37d2634, 32'h43fdf5f4, 32'h45464c64},
  {32'h451e6fe6, 32'hc2bcd458, 32'h432ceb62},
  {32'hc540db6a, 32'hc43580e2, 32'hc449065a},
  {32'h4391f6ca, 32'h4526e832, 32'h416d3bc2},
  {32'hc431b8ae, 32'hc2ff624d, 32'h40d799b1},
  {32'h43abc578, 32'h4502d8ef, 32'hc3314069},
  {32'hc3fc2de1, 32'hc4850811, 32'h4343ce87},
  {32'h4308f336, 32'hc3e03f9f, 32'h4403c594},
  {32'hc38e679c, 32'hc47980b3, 32'h4504352f},
  {32'h42fbf680, 32'h43a1f36e, 32'h43b97a20},
  {32'hc49aee8f, 32'h43179692, 32'h4449400f},
  {32'h43fe6499, 32'h44dda846, 32'h441df4c8},
  {32'hc48dd640, 32'h436cc90d, 32'hc3f5a98a},
  {32'h431f214f, 32'h44a3b021, 32'hc1225aba},
  {32'hc23fe05b, 32'hc5236b6e, 32'hc4016c41},
  {32'h4455b496, 32'h43b918ef, 32'h44ac4964},
  {32'hc3d95cf6, 32'hc504dbf7, 32'hc35a7169},
  {32'h446f0648, 32'hc44b2c5b, 32'h440a6209},
  {32'hc579127c, 32'hc25cc0f5, 32'hc3951524},
  {32'hc4c89387, 32'hc327e2e2, 32'h4315a115},
  {32'hc405b365, 32'hc4d798d2, 32'hc47667c6},
  {32'h4415aec5, 32'hc382265a, 32'hc3da371e},
  {32'h44be407c, 32'h439e5b60, 32'hc3fc5151},
  {32'h440b213e, 32'h44a7946b, 32'h440bccfa},
  {32'hc17ec200, 32'hc40a6b97, 32'hc4c0f185},
  {32'hc336a91a, 32'h44109ec7, 32'h4477fb25},
  {32'h449dce2b, 32'hc305071b, 32'hc39302e9},
  {32'hc24149c8, 32'hc55d1cea, 32'hc297af48},
  {32'h4340f8b0, 32'h44dec11f, 32'hc3c7bcfa},
  {32'hc47a6acb, 32'hc3080da9, 32'h428d55f8},
  {32'h4555b5d0, 32'h43156ffb, 32'h420e6816},
  {32'hc4e61387, 32'hc45bd8b8, 32'hc3c2987d},
  {32'hc41ceeaf, 32'h432f08ba, 32'hc4055233},
  {32'hc522083c, 32'hc3863b8d, 32'hc38afbb5},
  {32'h44e26816, 32'h43579412, 32'h44914382},
  {32'hc4f02330, 32'hc39c8d0a, 32'h423ede9a},
  {32'h4426c3d6, 32'h44821437, 32'hc4e0f86b},
  {32'hc3692476, 32'hc47f482a, 32'h450b2118},
  {32'h43b20ea7, 32'h447781a9, 32'h4353244e},
  {32'hc47fff8f, 32'hc2e6cde3, 32'h443bb228},
  {32'h447d73fa, 32'h43c56b62, 32'hc3fd9759},
  {32'h4482760b, 32'hc35f1890, 32'h4425aa3d},
  {32'h441dbcf1, 32'h43883afb, 32'hc3f7f911},
  {32'hc3def216, 32'h430e9a27, 32'h452b25f6},
  {32'h450f17be, 32'hc3d5055d, 32'hc43f4b95},
  {32'hc4362894, 32'hc48725c3, 32'h4469dc6b},
  {32'h444870fb, 32'h443a2739, 32'hc4ec3fd1},
  {32'h44961f6d, 32'hc35f2dfd, 32'h43eaf66e},
  {32'h44d44d8e, 32'h440c5807, 32'hc4088e35},
  {32'hc4362d9c, 32'hc4556e9a, 32'h44c491ec},
  {32'h4503679e, 32'h435bd0f4, 32'hc32b578a},
  {32'hc4e667af, 32'h43a5ff09, 32'h446ce751},
  {32'h4521f122, 32'hc1c86652, 32'hc4814374},
  {32'h440ab8d5, 32'hc47d21f9, 32'hc400e0e5},
  {32'hc4d457a1, 32'h4467057c, 32'h4406f223},
  {32'hc393e63a, 32'h4240a8ab, 32'h43e2c274},
  {32'hc527d1ae, 32'h43f39fd3, 32'hc48607c0},
  {32'h43b74f74, 32'hc5221f9c, 32'hc30d6910},
  {32'hc246c640, 32'h4369d6cc, 32'hc33fec5e},
  {32'h44abfd02, 32'hc4a8a501, 32'hc45336c0},
  {32'hc4095bee, 32'h44252272, 32'h444c07a1},
  {32'h45006868, 32'h4314300f, 32'h43b4114e},
  {32'hc2701500, 32'h4428e36c, 32'hc32358f2},
  {32'h449d2aa8, 32'hc4403b17, 32'h4418e3df},
  {32'h44a0e4da, 32'hc33f0723, 32'hc2f78a18},
  {32'h44ecc7a5, 32'hc38ec1c7, 32'h431d195b},
  {32'h4401aba3, 32'h4509e7d7, 32'hc1e6b061},
  {32'h449ea09a, 32'h4212d692, 32'hc4060687},
  {32'hc1e184d0, 32'h4419dfe3, 32'hc3112b40},
  {32'h4417432c, 32'h42d367d5, 32'h44a4f620},
  {32'h42229d76, 32'hc3516535, 32'hc51c874f},
  {32'h44473f76, 32'hc4f8ea6b, 32'hc342cd4e},
  {32'hc2794340, 32'h44195e59, 32'hc5030210},
  {32'h446f7c1b, 32'hc39af763, 32'h41f76023},
  {32'hc4013591, 32'h44da205e, 32'hc48b4693},
  {32'h43d2c40c, 32'hc4846ab2, 32'hc2d36332},
  {32'h4504aacc, 32'h43cc1911, 32'h43a2d66f},
  {32'h4331f9b8, 32'h4480625d, 32'h456183b4},
  {32'hc556d00f, 32'h43ee7c41, 32'hc3150bf0},
  {32'h4379f255, 32'hc2f6cea6, 32'h42b0001e},
  {32'hc4276ce9, 32'h42a305b0, 32'hc41543ed},
  {32'h419bc1e8, 32'hc4ee5236, 32'h450d1a99},
  {32'h43f58448, 32'hc44e8f94, 32'hc3cf2ca0},
  {32'hc3d9c1ab, 32'hc2bc2ddb, 32'hc471c978},
  {32'h435c1bbe, 32'hc494f654, 32'h4440ebe6},
  {32'hc436819b, 32'h441e4787, 32'hc461cdf2},
  {32'hc409b220, 32'h44070e72, 32'h445c4331},
  {32'hc4205f60, 32'h44920be0, 32'hc516cc3b},
  {32'h41bf5c88, 32'hc4c1df91, 32'h41eb66d4},
  {32'hc45b120b, 32'hc386e2f3, 32'h44f78ab6},
  {32'hc3d29d41, 32'hc3dbe53e, 32'hc522e1e8},
  {32'h44c7a324, 32'hc39b79a6, 32'h4321e183},
  {32'hc3b94307, 32'hc45ceb2c, 32'h438cbb4b},
  {32'hc4de01b2, 32'h42a56b30, 32'h43421949},
  {32'h449168fe, 32'hc3a918c1, 32'hc32be120},
  {32'h4228c678, 32'h4482e694, 32'hc48355bc},
  {32'h4445f70d, 32'hc2f1a523, 32'h44a0a9f2},
  {32'hc45094c5, 32'h446896e6, 32'hc2c3513c},
  {32'h4534418a, 32'hc3c73538, 32'h42a624c3},
  {32'hc46b581a, 32'h43aac134, 32'h441a6793},
  {32'hc3140206, 32'h4269d680, 32'hc386b601},
  {32'hc373efc7, 32'h444365bc, 32'h4345164f},
  {32'h44031d48, 32'hc4abf813, 32'hc3e822bc},
  {32'hc44dc11c, 32'h44f3d7f8, 32'hc3023af0},
  {32'h454e9fbe, 32'h43a776c4, 32'h4386d753},
  {32'hc5741cf5, 32'h440719e0, 32'h440458af},
  {32'h452e16e2, 32'hc42e2465, 32'hc3e7c51a},
  {32'h444d0f63, 32'h43de0169, 32'h43898063},
  {32'h4428f0e9, 32'h44b28e9f, 32'hc458cf32},
  {32'h433adf76, 32'h44adca5d, 32'h45002126},
  {32'hc3a3293c, 32'hc4834af1, 32'h43a9abce},
  {32'h4353d940, 32'h426c2bef, 32'hc4857216},
  {32'h4486bf70, 32'hc48171a2, 32'h4234582b},
  {32'h44a97e1a, 32'h444fd16f, 32'hc38db07c},
  {32'hc4071fc3, 32'hc3ff0d45, 32'h44d14654},
  {32'h44628f44, 32'h446a7f99, 32'h43cc4e21},
  {32'h4440a593, 32'hc37f0036, 32'hc39ac4d9},
  {32'h438d5bf0, 32'hc4c5956a, 32'h44f6673d},
  {32'hc2f76fc7, 32'hc4eaa5ee, 32'hc4f78083},
  {32'h4431b06e, 32'h4412bf34, 32'hc4832a54},
  {32'hc4aef63b, 32'hc4769321, 32'h43997fa0},
  {32'h44f381a7, 32'hc301efc5, 32'hc33cfe82},
  {32'hc418f50a, 32'h439a7a2f, 32'h4525057b},
  {32'h4120e300, 32'h43d9a0c6, 32'hc524b645},
  {32'hc374f254, 32'hc4319904, 32'h444e853c},
  {32'h453f9326, 32'hc3269404, 32'h4387e451},
  {32'hc5105281, 32'hc20537d1, 32'hc3852ea2},
  {32'h44b3072b, 32'h4368c98c, 32'hc2ee557d},
  {32'hc5078418, 32'hc49d60fd, 32'h4369cc35},
  {32'h45668a32, 32'h437c5fa2, 32'hc2ee1c6c},
  {32'hc236db20, 32'hc4e1a9a0, 32'h42323d66},
  {32'h4386a98e, 32'h44bdc074, 32'h42508247},
  {32'hc51823b1, 32'hc42a6d24, 32'h41974f22},
  {32'h42473e2b, 32'h43853f97, 32'hc190045c},
  {32'hc3d7b8ab, 32'hc41a066d, 32'h43a0cfdb},
  {32'hc3342170, 32'hc50f40a0, 32'hc40713fa},
  {32'h42d006fe, 32'h424279fe, 32'h44e11926},
  {32'hc3470ea6, 32'hc4ca7df5, 32'hc2f43747},
  {32'h42a49ef4, 32'h43be95eb, 32'hc3890190},
  {32'h4260b958, 32'hc48fed56, 32'hc4cba2ce},
  {32'hc4bcd6c7, 32'hc2d6cccb, 32'h43940ea7},
  {32'h437fbebc, 32'hc48dee6a, 32'hc50ac012},
  {32'h454a555a, 32'h43270287, 32'h4429c8b4},
  {32'h43dca330, 32'h441224bf, 32'h41f7eec0},
  {32'h42537ab7, 32'hc3662789, 32'h44905663},
  {32'h443c6b05, 32'h44b7b5bc, 32'hc5222673},
  {32'hc4e59574, 32'h431bebd9, 32'h42af1f56},
  {32'hc4cf818b, 32'hc3c7d471, 32'h4231b979},
  {32'h4492f64f, 32'h447e5ed6, 32'hc380a69c},
  {32'hc493ce9b, 32'hc35b4082, 32'hc411fcba},
  {32'h43637890, 32'h447a5197, 32'h44fd3457},
  {32'hc2c069ec, 32'hc4e8dd20, 32'hc4e468ee},
  {32'hc490f415, 32'h439d3102, 32'h4382b563},
  {32'hc4855e41, 32'hc50ee02f, 32'h440e654e},
  {32'h449fdbd6, 32'h44f02b8a, 32'hc14e8ca5},
  {32'hc426076c, 32'hc4342d9a, 32'h42d94cea},
  {32'h44c73a5f, 32'h4292813b, 32'h40bf2428},
  {32'hc45bd4a2, 32'hc4091731, 32'hc303b560},
  {32'h45525e56, 32'h43b6f8e3, 32'hc388d35c},
  {32'hc49f92ab, 32'h43003a84, 32'hc279bc32},
  {32'h44f04610, 32'hc21bc9dc, 32'hc1b65f84},
  {32'h441e8a61, 32'h436395d2, 32'hc49b5d90},
  {32'hc5333405, 32'h43ba21af, 32'h43a17ec7},
  {32'h4330d65e, 32'h449a8305, 32'hc41731d0},
  {32'hc49a9cf9, 32'h44dedbc4, 32'hc208fc57},
  {32'h450e375f, 32'h4305ad44, 32'h42b5543a},
  {32'h44d7df7e, 32'hc393b362, 32'h4279d678},
  {32'h45066cb8, 32'h41057770, 32'hc462b8bb},
  {32'hc5503b86, 32'hc3b2093a, 32'h43b6b929},
  {32'hc3fd66b6, 32'hc42cd8f3, 32'h42de7043},
  {32'h42cf05ac, 32'hc4a9ad94, 32'h44c4862d},
  {32'h41f81ef0, 32'h44a78505, 32'hc5318913},
  {32'hc42119fc, 32'hc40edef7, 32'hc27e547b},
  {32'h4407ba26, 32'hc43a1191, 32'hc41d5487},
  {32'hc394ad76, 32'h450a8cd4, 32'h446751fa},
  {32'hc4d95bd8, 32'h423fee56, 32'hc307f3c8},
  {32'h429b9f70, 32'h44eaec00, 32'h44a69359},
  {32'h4433b970, 32'h432ec45a, 32'hc49bf351},
  {32'h43e84744, 32'h422c9842, 32'h449f7780},
  {32'h42462350, 32'hc586518d, 32'h42fc9469},
  {32'hc55ad2e8, 32'h4439ab90, 32'hc370659e},
  {32'h450f4898, 32'h43d04565, 32'h4382c685},
  {32'hc1c02ec0, 32'h44ef9b14, 32'hc408c564},
  {32'h42fb0250, 32'hc53f20e9, 32'hc3ecb678},
  {32'hc35a4c63, 32'h449ee44b, 32'h42c78db0},
  {32'hc336fc88, 32'h443aba7d, 32'h4340d54f},
  {32'hc54df262, 32'hc18d7544, 32'hc3a52b52},
  {32'h457878d1, 32'h4250d203, 32'h431919f7},
  {32'h450aa226, 32'hc3847100, 32'hc38cf458},
  {32'hc3e0e698, 32'h42b6bcd6, 32'hc3cad812},
  {32'h44ee7f2f, 32'hc2aec0b2, 32'h4483a91f},
  {32'h4448e311, 32'h42ef99fe, 32'hc31f9695},
  {32'h44ef7116, 32'hc4b6b61f, 32'hc2bdb56b},
  {32'hc46d0cb9, 32'h44b17e1d, 32'h43a045ab},
  {32'h42b3f224, 32'h42e5b5fa, 32'hc376fe05},
  {32'hc1b7ea0f, 32'h4573a84f, 32'h40d9353b},
  {32'h4506ce8c, 32'hc413c67a, 32'h438e319d},
  {32'h441c4cc6, 32'hc3c31c4a, 32'hc3a3144a},
  {32'h44529dd8, 32'hc39f5ade, 32'hc40afd48},
  {32'hc3c9306c, 32'h4363f466, 32'hc52b40e2},
  {32'hc483876e, 32'hc2930f70, 32'hc266b1d1},
  {32'hc3953006, 32'h44db8eda, 32'h43f9fe52},
  {32'hc392838b, 32'hc188b431, 32'hc5366550},
  {32'h4220b35c, 32'h43f1db7d, 32'h44db306d},
  {32'h44faceeb, 32'h42352d13, 32'hc03892ac},
  {32'h433b47ba, 32'h44d57008, 32'h42b5ff57},
  {32'h4525385d, 32'hc2e9734c, 32'h436b6148},
  {32'hc2d2e068, 32'hc44db63d, 32'h44aa0b29},
  {32'h447dee4c, 32'h44280d9e, 32'hc49ba3fa},
  {32'hc47b246b, 32'h440e9714, 32'h4283aa0b},
  {32'hc2cbadca, 32'hc37d1218, 32'hc51eb02f},
  {32'hc4f16e67, 32'h439af0ab, 32'h43f6339e},
  {32'hc3ea3e75, 32'hc3196192, 32'hc411fc38},
  {32'hc5510d48, 32'h448afd2a, 32'hc2af8520},
  {32'h4405b4c8, 32'hc50d3b22, 32'hc3acb8ae},
  {32'h44c0fc32, 32'h4343aa64, 32'hc51c2cb0},
  {32'hc35b530e, 32'h4387f38b, 32'h455fe83f},
  {32'h45069b63, 32'h403b932c, 32'h42ba50df},
  {32'hc492f6f5, 32'hc4642225, 32'hc1633bc3},
  {32'h44838924, 32'h44920f4e, 32'hc35675c6},
  {32'h4448c953, 32'hc30e3221, 32'hc3f23fd8},
  {32'h43120cb0, 32'h4494cf71, 32'h43b2fd6f},
  {32'hc11048a0, 32'hc5215734, 32'h42179584},
  {32'h44bc5b7e, 32'hc329caff, 32'h4390d52d},
  {32'hc4bdbc9a, 32'hc3393ae4, 32'h441241cf},
  {32'h448c9294, 32'h43a21de9, 32'hc3313cc7},
  {32'hc535e3ae, 32'hc1130a82, 32'h4365ca11},
  {32'h45428b43, 32'h4295ece5, 32'h43530e1e},
  {32'hc40b8f97, 32'hc405d994, 32'hc4d03d21},
  {32'h426eadd6, 32'h44c3562c, 32'h437285c4},
  {32'hc3d884a0, 32'hc4d93c6b, 32'hc38fb914},
  {32'h43ac3364, 32'h4474c102, 32'h44a4148f},
  {32'hc4b69311, 32'hc433c5f2, 32'h4316249b},
  {32'hc1ef06b8, 32'h42e75d09, 32'h44b1c8d0},
  {32'hc494b4a4, 32'hc41d7fc2, 32'hc38a47b2},
  {32'h454f0a15, 32'hc3195ef0, 32'hc313976a},
  {32'hc4e1cdcb, 32'hc4632df6, 32'h43325ff1},
  {32'hc3231069, 32'h45433140, 32'hc391a4ff},
  {32'h43a5a17f, 32'h43c93b64, 32'hc29a487d},
  {32'hc319a18e, 32'h445a0928, 32'h45596344},
  {32'hc5030d6b, 32'hc3c676e1, 32'hc32b8326},
  {32'h44e54d30, 32'h435d39af, 32'h42083b7d},
  {32'h447360bc, 32'h43a53e9e, 32'hc3d66140},
  {32'hc40c9ec3, 32'hc4f792b5, 32'hc3a4e380},
  {32'h42679444, 32'h452f0dea, 32'h44393f7d},
  {32'hc43ebb05, 32'hc3b8963b, 32'h42dee99f},
  {32'hc3411722, 32'h455a06c2, 32'h42bc2090},
  {32'hc56239a0, 32'h42985582, 32'h434382a8},
  {32'h4532a414, 32'h43f33d58, 32'hc33884de},
  {32'hc4ace85c, 32'hc42091cb, 32'hc43a8d3f},
  {32'h454bba5e, 32'hc0837c8d, 32'h43499c11},
  {32'hc4550c7e, 32'hc382cb7d, 32'h44101b1f},
  {32'h442a578f, 32'h44b1258e, 32'h4165c9e7},
  {32'hc530d7c4, 32'h3f644c20, 32'h424bc541},
  {32'hc24f6ee8, 32'h450f89e7, 32'hc2d22ac6},
  {32'hc4efaacb, 32'hc415d005, 32'h430dbf1a},
  {32'h43278330, 32'hc1fc73e2, 32'hc4fb18f3},
  {32'h44d36da8, 32'hc1b2f23a, 32'hc29fad7a},
  {32'h443d56a0, 32'h4497de02, 32'h444818d9},
  {32'hc4b3cf7e, 32'h4309c17a, 32'h4427a6a3},
  {32'hc4ecc9c0, 32'h42576144, 32'hc3835852},
  {32'hc3d0e99c, 32'hc4966e7b, 32'h450318ad},
  {32'h43368990, 32'h44e6e4dc, 32'hc4063a35},
  {32'hc45b85c1, 32'h415b08b2, 32'hc3a56575},
  {32'hc404feb3, 32'h453fe1f8, 32'h4305c282},
  {32'hc3a45600, 32'h430eac9d, 32'h44eed9b0},
  {32'hc466d50a, 32'hc2551854, 32'hc2a6c72c},
  {32'hc4044b96, 32'h4437a8ba, 32'h455b4a2f},
  {32'h43b430e0, 32'h42e3c0ba, 32'hc31bb453},
  {32'hc1255a80, 32'hc4e28bcb, 32'hc3ddc6a4},
  {32'hc491c34d, 32'h44d16464, 32'h43b16273},
  {32'h44656186, 32'hc4326b94, 32'hc3ab0520},
  {32'hc4ac1e4d, 32'h44b5dfb2, 32'hc3a4ea6d},
  {32'h43aadfc2, 32'hc54e7bb6, 32'h431c4dcf},
  {32'h431420a8, 32'h43afe6e2, 32'hc256db43},
  {32'h44cf4373, 32'hc462490e, 32'hc4589aa0},
  {32'hc4b1ee88, 32'h44ab3502, 32'h448b7612},
  {32'h44a07bf6, 32'hc26ae812, 32'hc1631271},
  {32'hc4a75970, 32'h44016252, 32'hc4a647eb},
  {32'h44453ef9, 32'hc35991f4, 32'h443ce15a},
  {32'h448fde65, 32'hc3935f04, 32'h43b5cf0f},
  {32'hc364a546, 32'hc4905540, 32'h44672055},
  {32'hc4422dac, 32'hc422de9d, 32'hc54fa4f3},
  {32'h443de219, 32'hc478c1d0, 32'h42a4e8b3},
  {32'hc4306dd6, 32'hc364d3d5, 32'hc4fd9859},
  {32'h4514e901, 32'h433e9c11, 32'h434f7df4},
  {32'h439fdb1c, 32'h43c13f75, 32'hc4e1d2f0},
  {32'h451ce61e, 32'hc419cb35, 32'h43e3d41d},
  {32'hc343f395, 32'h43f6d13c, 32'hc5214def},
  {32'h4530aa9c, 32'h430bff2d, 32'hc4088e1b},
  {32'hc302f06b, 32'h42fa7bd4, 32'hc5102eea},
  {32'hc3e9cf7f, 32'hc46bc6db, 32'h43e23b39},
  {32'hc512e63c, 32'h4258c403, 32'h42a243b2},
  {32'h4488f097, 32'h430ac358, 32'h44cd5a59},
  {32'hc4bd5c6e, 32'h4440bf65, 32'hc43ffa9b},
  {32'h44ead9f4, 32'h438f9307, 32'hc3226f35},
  {32'h44666e8a, 32'h447649fe, 32'hc50bfedd},
  {32'h44d21f4c, 32'hc3abd581, 32'hc36362fb},
  {32'h4393e00f, 32'hc4043d07, 32'hc48a6daa},
  {32'hc463f997, 32'h442a74f7, 32'hc32597bd},
  {32'h4400630c, 32'h42c6a346, 32'h446e22da},
  {32'hc3c29514, 32'h448fcc20, 32'hc31d2024},
  {32'h44d1ae86, 32'hc10cbbb8, 32'h432ce04f},
  {32'hc5486d89, 32'h428817af, 32'hc3a4ae14},
  {32'h43a2be7a, 32'hc4ee22e4, 32'h441706ae},
  {32'h4406563b, 32'h44efc899, 32'h4492f0ff},
  {32'hc198f810, 32'h4327d98c, 32'hc52de5ea},
  {32'hc38f09f9, 32'h42255cfc, 32'h43b87c14},
  {32'h44c16931, 32'h43b92ae8, 32'h4215b01c},
  {32'hc367b25c, 32'h441e7eb9, 32'hc47dbd28},
  {32'h4391bb58, 32'hc3e248ed, 32'h44cb9e93},
  {32'hc4bfdab5, 32'hc3ebc5b7, 32'h42a3e3b6},
  {32'h446984f0, 32'hc3c6f29c, 32'h44a8c445},
  {32'hc3634c2c, 32'h44e42e50, 32'hc48b6d53},
  {32'h453283ea, 32'h42014d1d, 32'h43f47a45},
  {32'hc5962ded, 32'hc312f1d1, 32'h41b812f9},
  {32'h45482783, 32'hc2b58719, 32'h44112409},
  {32'hc53a3975, 32'hc3d2a03d, 32'h41758b18},
  {32'h4451eed4, 32'hc4600177, 32'h44366224},
  {32'hc42359ec, 32'h44ba8e0c, 32'hc40290a3},
  {32'hc44c5e7b, 32'hc3c8f636, 32'h425ed91a},
  {32'hc456b74f, 32'h448bfa08, 32'h4344108d},
  {32'h450db8b9, 32'hc42fa3e0, 32'h43f2c3e0},
  {32'hc42ece72, 32'hc488a6b1, 32'h44115f8b},
  {32'h43e21064, 32'hc400a344, 32'hc42c9aaf},
  {32'h43a0efde, 32'h43c53975, 32'h454e8578},
  {32'hc4a7d0cc, 32'hc44fb25c, 32'h437c030b},
  {32'h42ad1adc, 32'h45380c2e, 32'h43e8de37},
  {32'hc4554452, 32'hc207da85, 32'h4423b65a},
  {32'h42e71dc0, 32'hc33569f1, 32'hc520aaf0},
  {32'hc3c1881a, 32'hc3a0486e, 32'h45036b0a},
  {32'h44d4ce82, 32'h4343be5b, 32'hc3a39546},
  {32'hc4c9b169, 32'hc2940d73, 32'h438b3c7b},
  {32'hbfd57900, 32'hc49c5cfe, 32'h450c1604},
  {32'h4359ed98, 32'h44aef9ed, 32'hc4da3dc6},
  {32'h43f234b0, 32'h4527a1ff, 32'h4307d368},
  {32'hc44b6353, 32'hc31c5beb, 32'h44a6c827},
  {32'h4489c5ff, 32'h4398a495, 32'hc460ae0b},
  {32'hc3cdeeb5, 32'hc47e3c9b, 32'h43a4eed8},
  {32'h439eab9a, 32'hc3bff4c1, 32'hc51699be},
  {32'hc3e8c909, 32'hc4a27ece, 32'h437a013f},
  {32'h4415969d, 32'h427aa17b, 32'h43b72774},
  {32'hc55973d5, 32'hc26e20df, 32'h427cfde3},
  {32'hc4a1e9a5, 32'h4389a300, 32'hc2bc93a4},
  {32'hc4c21266, 32'hc4675231, 32'h43586048},
  {32'h44e34fb8, 32'h43d65ecb, 32'h4407d998},
  {32'hc4b6250e, 32'hc4026a74, 32'h43a0cd39},
  {32'h44550604, 32'h44bbd836, 32'hc27f6740},
  {32'hc44b09d4, 32'hc4d45e36, 32'hc3e8f969},
  {32'h41a2b825, 32'h449efbca, 32'h427cf921},
  {32'hc3411210, 32'h434d3444, 32'h439d029a},
  {32'hc39ccf5c, 32'h43e771b9, 32'hc4ab6f58},
  {32'h4108ab00, 32'h437de2ca, 32'hc3aef806},
  {32'hbfc72500, 32'hc4ad31bd, 32'hc28916e1},
  {32'h43d00854, 32'h4482ee45, 32'h448b8981},
  {32'h43ae6dfd, 32'hc3ae23bb, 32'hc5286241},
  {32'h45312581, 32'h4363bcc7, 32'hc337ee40},
  {32'hc4451770, 32'hc4fdaf65, 32'hc4e438d7},
  {32'h43876f7c, 32'h450a5d77, 32'h4487e760},
  {32'h42d2f726, 32'hc3f8c361, 32'h4182ac3a},
  {32'hc27f6729, 32'h4287798b, 32'h445701f4},
  {32'hc41e6637, 32'h4370e7df, 32'hc4137a1a},
  {32'hc3803c29, 32'h448bde20, 32'h43fe8e7e},
  {32'hc47a5858, 32'hc44bf8a8, 32'hc29a8d9a},
  {32'hc1d6aca0, 32'h442036f8, 32'h4543f8a0},
  {32'h44a31a52, 32'hc4170d50, 32'hc48de7d7},
  {32'h44b079b9, 32'h426b9736, 32'h444288b3},
  {32'hc478e1c3, 32'hc40a1968, 32'hc4c4b71a},
  {32'hc4def5f8, 32'h439d191f, 32'h43f2b2a3},
  {32'hc30a6784, 32'hc5619fcb, 32'hc2543952},
  {32'hc3278e67, 32'h457ce405, 32'hc225bcaa},
  {32'h449766e7, 32'h420626ba, 32'h4278454c},
  {32'h443ca8c9, 32'h450b52d8, 32'h43c93051},
  {32'hc50b874e, 32'hc41b08d1, 32'hc1272b46},
  {32'h448774d6, 32'hc2347501, 32'hc2bcf2c4},
  {32'hc52db6c2, 32'h43390b6f, 32'hc3c357d8},
  {32'h448763e0, 32'hc40fe99a, 32'h4422a29b},
  {32'h4421401c, 32'hc4896b6b, 32'hc47afb94},
  {32'h42ee023e, 32'hc490335d, 32'h44b1b350},
  {32'hc426cf30, 32'h43525263, 32'hc45d3905},
  {32'h42ce1c40, 32'h44193557, 32'h44b2ade1},
  {32'h4443cc2e, 32'hc4487257, 32'hc3912593},
  {32'h43b66a5b, 32'hc3941e0a, 32'h44387d76},
  {32'hc319cd42, 32'hc50b3da8, 32'hc4ebbb46},
  {32'hc2b6b5c8, 32'h447fdaed, 32'h45320ee1},
  {32'h44be4217, 32'hc324804a, 32'h4356ea90},
  {32'hc4804496, 32'h4454e020, 32'h436e56ed},
  {32'hc36d567e, 32'h43f445f6, 32'hc5111a76},
  {32'h42c9f781, 32'hc47bc0d9, 32'h444108d3},
  {32'hc4124731, 32'hc40ae443, 32'hc4e88baa},
  {32'hc51169ac, 32'h4295bf4f, 32'hc2840b36},
  {32'h450e557e, 32'h43a7c912, 32'hc40a0fde},
  {32'hc49fc4be, 32'h42902108, 32'h4498e6d0},
  {32'hc47030f9, 32'hc31436c7, 32'hc4c02161},
  {32'h44298f3f, 32'h44261632, 32'h43c48b88},
  {32'hc37b6bf0, 32'hc504fbe9, 32'hc46c6ab9},
  {32'hc4871124, 32'h44974100, 32'h43086100},
  {32'h4532711b, 32'hc31718dd, 32'h416b434a},
  {32'h4200f550, 32'h43ac0072, 32'hc41eb274},
  {32'h43bf21fa, 32'hc503a142, 32'hc3af216c},
  {32'h44f25f52, 32'h406f6977, 32'hc30ebc03},
  {32'h44e9bf52, 32'h43227d96, 32'hc2f756b9},
  {32'hc5866a7c, 32'h4232428a, 32'hc34640d6},
  {32'h445087c0, 32'hc25a4c49, 32'hc3d455ec},
  {32'h44dccfdf, 32'hc3796e58, 32'h41d42978},
  {32'hc4ef8aac, 32'hc413eb54, 32'h43806e68},
  {32'hc20aab80, 32'h43728ad0, 32'h452a32ef},
  {32'h42848df7, 32'hc3330743, 32'hc398902b},
  {32'hc182aa00, 32'hc33df7be, 32'hc40b3b9b},
  {32'hc3c81b24, 32'h4511cf19, 32'h43a864a6},
  {32'h451ed51f, 32'h4403a4ef, 32'hc2dc0339},
  {32'hc249edf4, 32'h45850aff, 32'h42a573b3},
  {32'h430d1c76, 32'hc43af309, 32'h44081de9},
  {32'hc3b2f38c, 32'h43947503, 32'hc432c011},
  {32'h450f82b6, 32'h42e5a8c0, 32'hc297c5cc},
  {32'hc4adb9c9, 32'hc31e2295, 32'hc1a23ac8},
  {32'h44f35d86, 32'h425bfe7f, 32'hc30e30fe},
  {32'hc3f39604, 32'h4394297c, 32'h44669795},
  {32'hc2c9872c, 32'hc520c9ab, 32'hc38f952e},
  {32'h43ad7064, 32'h43d079a9, 32'h44d307b2},
  {32'h452da3a2, 32'hc2e75a73, 32'hc3ac3105},
  {32'hc4547289, 32'h4454718a, 32'hc2823d1c},
  {32'h453e3c22, 32'hc38026f3, 32'hc26322f9},
  {32'hc5315ec2, 32'h43ddfe74, 32'h43abb92d},
  {32'h455faa31, 32'h43236b20, 32'h4180c00f},
  {32'h44636199, 32'h4233b350, 32'h448cbc44},
  {32'h4539bd52, 32'hc448796c, 32'h434803ae},
  {32'hc380ee81, 32'h444914a8, 32'h452be7d3},
  {32'hc1f1ec26, 32'hc487aacf, 32'hc3a5e7e6},
  {32'hc4833a6b, 32'h43c7393e, 32'h44835d37},
  {32'h44b1ea26, 32'hc4a7b5de, 32'hc4642ee1},
  {32'h452f599a, 32'hc327c2b8, 32'hc3f43a51},
  {32'hc50c14fa, 32'hc365ec3a, 32'h44a7b072},
  {32'hc49a8f1c, 32'h433ffba1, 32'h41b373de},
  {32'hc3c08548, 32'hc3aabb64, 32'hc384bbb1},
  {32'h44ebd1dd, 32'h4435c340, 32'h43b5c814},
  {32'hc382cf19, 32'hc50f5013, 32'h435f9f9c},
  {32'h4491a726, 32'h45155fa7, 32'h426b13cf},
  {32'hc58b9448, 32'hc292714f, 32'hc3d6af58},
  {32'h42135110, 32'h430db727, 32'h444d2a81},
  {32'hc40c61a6, 32'hc4522043, 32'h44a6fd74},
  {32'h43b3f0e8, 32'hc2010ff4, 32'hc5059491},
  {32'h4238f942, 32'h4296cb64, 32'h44372e39},
  {32'h441e10e3, 32'hc28bdcd6, 32'h44d0c835},
  {32'hc4a61b16, 32'hc356a910, 32'hc46d69d7},
  {32'h4443f7d7, 32'h446e0a8a, 32'h42644e12},
  {32'hc324698a, 32'hc4433a51, 32'hc464f4b9},
  {32'hc3948e02, 32'h4470ddbd, 32'h43a74088},
  {32'h442e8c60, 32'hc36b9508, 32'hc39aafcb},
  {32'hc1225500, 32'h4415dbbd, 32'h43a747f8},
  {32'hc523ffcc, 32'hc3611ea8, 32'hc3d2c8bf},
  {32'h439610f4, 32'hc37f5fd9, 32'h422bdf5a},
  {32'hc490c1dd, 32'hc3ef4df6, 32'hc4a5357a},
  {32'hc37be9da, 32'h43efb57b, 32'h450bbe49},
  {32'h44127e92, 32'hc2c2fe45, 32'hc2c0b1b4},
  {32'h4347095e, 32'h454bb3f5, 32'h4334ffe1},
  {32'hc3fe1751, 32'hc3efb6a0, 32'hc4ded5f2},
  {32'hc2c9e6b4, 32'h44d4ae44, 32'h42120ef4},
  {32'hc4021ff6, 32'h4362436f, 32'h436d4270},
  {32'hc3432d64, 32'hc4e5fe98, 32'hc3139519},
  {32'h4414f7a7, 32'h4510a12d, 32'hbfe71260},
  {32'h4410782b, 32'hc4300bf7, 32'hc321d2a5},
  {32'h4404264b, 32'h446b72c1, 32'hc29f74dc},
  {32'hc4eda193, 32'hc45d4096, 32'hc3810428},
  {32'h4509bb4a, 32'h43422ade, 32'hc39c5a00},
  {32'hc44f86ac, 32'hc3d83bf7, 32'h424e9e9b},
  {32'h44bc9b06, 32'hc1413d74, 32'hc36ef484},
  {32'h43ce634e, 32'hc40191ed, 32'h4435c07a},
  {32'h43c40106, 32'h44f48ace, 32'hc2b264ac},
  {32'hc43bb8a9, 32'hc44c47a9, 32'hc314c365},
  {32'h4450b0b9, 32'h44749af9, 32'hc3a1b04f},
  {32'hc4c0464c, 32'h40d2da4c, 32'hc32f8778},
  {32'hc398e3de, 32'hc20b5564, 32'hc53331f2},
  {32'h44956451, 32'hc266f291, 32'h42b95a83},
  {32'h454077da, 32'hc30e8596, 32'hc3316a23},
  {32'hc49b9f49, 32'hc2f8ac0f, 32'h4432119f},
  {32'h4432c866, 32'h448c29aa, 32'hc3a14097},
  {32'hc4f138cc, 32'h41ce389b, 32'h440192f2},
  {32'h4480ffd0, 32'h44a8a525, 32'hc4a3e941},
  {32'h4491de45, 32'h42f35c40, 32'hc0cd1c68},
  {32'h4387a964, 32'h4425a937, 32'hc4b41869},
  {32'hc52f2293, 32'hc3b76f51, 32'h43768001},
  {32'h450676f6, 32'h4396a6e6, 32'h43dd10bc},
  {32'hc3e7c4b8, 32'h441a4dbb, 32'h452c3ea2},
  {32'h44720ada, 32'hc41f97df, 32'hc4736c39},
  {32'hc3a66d18, 32'h4286adde, 32'hc49a93fd},
  {32'hc4837ff5, 32'h43e88831, 32'h446c6798},
  {32'hc429f058, 32'h43e779c0, 32'hc3aa77f3},
  {32'h43ed7074, 32'h449c63c0, 32'hc41a91bf},
  {32'h44c32f8f, 32'hc49572f9, 32'hc393ed72},
  {32'hc4f6a7c8, 32'h43a89110, 32'hc3ec1b47},
  {32'h4205e600, 32'hc394645c, 32'hc1e32736},
  {32'hc586b720, 32'h4445fef6, 32'hc3baeba3},
  {32'hc2bbe18c, 32'hc400177f, 32'h43768068},
  {32'h43a03bc8, 32'h44b32793, 32'h4380ae6d},
  {32'h43c6a882, 32'hc443e40f, 32'h43ecf913},
  {32'hc471c863, 32'hc17237e0, 32'hc4544b7a},
  {32'hc33197f8, 32'hc4a586ca, 32'h43e04759},
  {32'hc53d5c8c, 32'hc363d284, 32'h4363037b},
  {32'h44f89648, 32'hc305bfac, 32'hc10927aa},
  {32'hc490d336, 32'hc3ccd249, 32'hc4d0faf5},
  {32'h4377e630, 32'hc3f25256, 32'hc3ccfb2b},
  {32'h440167fa, 32'h444b194a, 32'h43274579},
  {32'h437ff2fe, 32'hc42f80cc, 32'h44d38fd8},
  {32'hc4ca0579, 32'h43f61471, 32'hc398640b},
  {32'h453e3c89, 32'hc31455e7, 32'hc398582b},
  {32'hc4655866, 32'h44a1cf03, 32'hc2fcc156},
  {32'h43317150, 32'hc3bff007, 32'h44dfb06c},
  {32'h43052fc3, 32'h4449379f, 32'hc3b89ef9},
  {32'h45259887, 32'h4443cc8a, 32'h441516ee},
  {32'hc5448fee, 32'hc345ca7b, 32'hc3c5aa1e},
  {32'h4401e84a, 32'h43532593, 32'h439e97cd},
  {32'hc493b8d5, 32'hc4b7861e, 32'hc45378b1},
  {32'h44deb072, 32'hc3a13f98, 32'hc308ad01},
  {32'hc4444230, 32'h44428aa3, 32'h437eb9af},
  {32'hc3a40dbe, 32'h44e248df, 32'h43aabe71},
  {32'h43cc5c28, 32'h4049f77a, 32'h4514dd22},
  {32'hc3d25a58, 32'h44c8c70a, 32'h42c4ffd5},
  {32'h44cd93a6, 32'h436b06fe, 32'hc0e13c08},
  {32'hc38eb3e2, 32'h4502d628, 32'h41ee12bf},
  {32'h43ff15e5, 32'hc50d8f29, 32'h428f16e7},
  {32'h44850046, 32'hc5164d50, 32'h44f9acd4},
  {32'hc3d731df, 32'h44daa85f, 32'hc49d7987},
  {32'h441ba36e, 32'hc2e39bee, 32'h43307013},
  {32'hc29c39dd, 32'hc3177225, 32'h44de5853},
  {32'h4333dee0, 32'h448942ae, 32'hc4506301},
  {32'h44a0fdaf, 32'hc4c27445, 32'hc4219a93},
  {32'hc4047730, 32'hc182ba69, 32'hc48bb0c6},
  {32'h449ce1fc, 32'h433374eb, 32'h441bcb71},
  {32'hc4b027a7, 32'h43cfb5a2, 32'hc3ad09d3},
  {32'hc4824946, 32'hc3fd3b51, 32'h4301a074},
  {32'hc4e9c494, 32'h43e0603a, 32'hc3ef2759},
  {32'h45206ef5, 32'h4409c05e, 32'hc35c32ec},
  {32'hc425d97c, 32'h4456bdaf, 32'h4338860a},
  {32'h44deb5c1, 32'hc2f08fdb, 32'h4222d489},
  {32'hc4fe5c82, 32'h44146457, 32'hc32cce64},
  {32'h44912f76, 32'hc445b8fd, 32'h42cf69de},
  {32'hc4d9b576, 32'h44acd81c, 32'h43bce24b},
  {32'h443beb81, 32'hc50e30dd, 32'hc34d68be},
  {32'h43ffae1e, 32'h449fe00a, 32'h43f17c1b},
  {32'h42a4158c, 32'h411d56c4, 32'hc574b50e},
  {32'hc310ef1d, 32'h4485b84f, 32'h4543fdc8},
  {32'h43a57192, 32'hc2ab14c4, 32'h45426e85},
  {32'h4479fe76, 32'h4423f7ff, 32'hc429db56},
  {32'hc48a92c3, 32'hc501121e, 32'h430832db},
  {32'h43f0c368, 32'h44df0457, 32'hc4026688},
  {32'h4454b6eb, 32'hc492ea4d, 32'h44971608},
  {32'h44dbd0c6, 32'hc3a47d25, 32'hc43a7511},
  {32'hc23e8b12, 32'hc48a8f11, 32'hc423d2dc},
  {32'hc42f68b0, 32'hc4c75330, 32'h44e1a5d1},
  {32'hc3bd1cb3, 32'hc4937cf5, 32'hc52176a2},
  {32'h45131504, 32'h43d3157a, 32'hc3be6c13},
  {32'hc2e03334, 32'hc4213026, 32'h445a172d},
  {32'h438b2f8a, 32'hc2e0b28a, 32'hc4958830},
  {32'hc3a548fd, 32'hc2f83dbe, 32'h44373b85},
  {32'h44a82b2d, 32'h442a1061, 32'h42ec7d5e},
  {32'h44b793cd, 32'hc31a7174, 32'hc2781408},
  {32'h455af590, 32'hc3fdff89, 32'hc2db6227},
  {32'hc583bc2d, 32'h432df5d9, 32'h4315f942},
  {32'hc4b31aa4, 32'hc2dbcddf, 32'hc2af1c22},
  {32'hc4ee379e, 32'hc44a41e4, 32'h43a396d2},
  {32'h44226dca, 32'h44f293d9, 32'hc3cecdf8},
  {32'hc4f05526, 32'hc405832c, 32'hc16d9214},
  {32'h4520fb46, 32'h442e0596, 32'hc38abbeb},
  {32'hc4d83dd4, 32'hc446c17e, 32'h43eaf2b2},
  {32'h44845175, 32'h4295006e, 32'hc3306dd0},
  {32'hc473af8c, 32'h43265390, 32'hc38acff4},
  {32'hc38d1cdd, 32'hc49b1125, 32'hc41e3673},
  {32'h43620290, 32'h444c8f07, 32'h44b17211},
  {32'h44e7b914, 32'hc2901bf7, 32'hc1aee516},
  {32'h440f26cd, 32'h450c4c7d, 32'hc265a818},
  {32'h42c71885, 32'hc4f134a5, 32'h4222d1be},
  {32'h447ec934, 32'h43dad65a, 32'hc290e746},
  {32'hc54f7ab6, 32'hc3ca63e6, 32'h429cdeb5},
  {32'h44b92388, 32'hc02e3654, 32'h44724da8},
  {32'hc2a14d1a, 32'hc3cdcd4c, 32'hc394f593},
  {32'h448c1e5d, 32'h4493bcec, 32'hc3abf32f},
  {32'hc40523f5, 32'hc4999443, 32'hc3c54b86},
  {32'hc182c38c, 32'h43391551, 32'h44562363},
  {32'hc3b31c69, 32'hc561d295, 32'hc3dd1622},
  {32'h4486daa8, 32'h4482b608, 32'hc2646f15},
  {32'h43b38a67, 32'hc4a83ae5, 32'hc44d8a8c},
  {32'h4519ab5f, 32'h43a81f72, 32'h4430d760},
  {32'hc40f4c18, 32'hc39042d5, 32'hc51f412e},
  {32'hc40ec588, 32'h431a8995, 32'h43bf3498},
  {32'hc48fae1a, 32'hc4ab1041, 32'hc3c0e3ea},
  {32'hc38d14d0, 32'h447fc42e, 32'h43988b48},
  {32'h43babefc, 32'hc48f90f4, 32'hc3e49bec},
  {32'h43cd8274, 32'h44e4b88a, 32'h430e1470},
  {32'hc42964f7, 32'hc41803f1, 32'h43687342},
  {32'h42606360, 32'h43974ab8, 32'h43793fac},
  {32'hc56cc40f, 32'h43a2e9cf, 32'hc402bb32},
  {32'h455a5684, 32'h431e5b53, 32'h438ae634},
  {32'h45169c5a, 32'hc3fc35e6, 32'hc4637dc2},
  {32'h438d4cbd, 32'hc40b94b1, 32'h44e8429b},
  {32'hc382b7a9, 32'hc33bde22, 32'hc39b7e39},
  {32'hc3ba081c, 32'h45002e61, 32'h4321b96c},
  {32'hc39afd33, 32'hc41a75bc, 32'hc4f965d3},
  {32'h44320801, 32'h42958c29, 32'h44050c14},
  {32'h42b485e0, 32'hc4ee5aaf, 32'hc501d56e},
  {32'hc48107ad, 32'h441f20c9, 32'h449934eb},
  {32'hc3806e5c, 32'hc37c6ea1, 32'hc5114f43},
  {32'h43b93ad2, 32'h452480d6, 32'h43ba91ff},
  {32'hc1db0e6b, 32'hc48958c6, 32'hc494bb6d},
  {32'hc3461f84, 32'hc30080ff, 32'h4443a735},
  {32'hc3ce0e70, 32'hc42783ff, 32'hc476591a},
  {32'hc425f314, 32'h455fb8bf, 32'h42acd037},
  {32'hc38529b0, 32'hc195ba4c, 32'hc3e11a28},
  {32'hc4708c7b, 32'hc0817309, 32'h448774e2},
  {32'hc30f0247, 32'hc367d80a, 32'hc4071433},
  {32'h441abee6, 32'h41622e60, 32'h44ba44b3},
  {32'h43dc2d2c, 32'hc50912b3, 32'hc33f24f6},
  {32'hc479b368, 32'h4481ec5d, 32'hc2e6c730},
  {32'h4503bd0a, 32'h44384670, 32'h43d79eb0},
  {32'h4396dea4, 32'h444ef0a0, 32'h44228b72},
  {32'h44ca7a44, 32'hc35d214a, 32'hc34f71ba},
  {32'h442d012a, 32'hc184dc50, 32'hc1be65fa},
  {32'hc2129922, 32'hc290ef86, 32'h431aa13c},
  {32'hc549e9a9, 32'hc340fe1e, 32'h43b711e2},
  {32'h44ae2e69, 32'h43053ec2, 32'hc40269c5},
  {32'h4315d01e, 32'h43d12d8f, 32'hc3dd4d16},
  {32'hc424123c, 32'hc450394c, 32'hc5337ca7},
  {32'h44d4ede4, 32'h43f148e6, 32'h436ed40c},
  {32'hc4fbc9aa, 32'hc35c66eb, 32'h431d2063},
  {32'h44741d84, 32'hc5209cc5, 32'hc312b37f},
  {32'h4367c0cb, 32'h4566672a, 32'h43239337},
  {32'h44eed81f, 32'h43ef6d42, 32'h42e24cf2},
  {32'hc27525d0, 32'h44a896a4, 32'hc350b3c9},
  {32'hc1d86680, 32'hc50f76ae, 32'hc39302e3},
  {32'h43aa4f6c, 32'h44610c21, 32'h438b28df},
  {32'h443985be, 32'hc4228bad, 32'hc4085426},
  {32'hc4196e38, 32'hc2b1b26d, 32'hc4a86dda},
  {32'h43b39417, 32'hc3468473, 32'hc47dc743},
  {32'hc485622f, 32'h447ba8f4, 32'h43faa833},
  {32'h446874f3, 32'hc39e85e6, 32'hc4cd9288},
  {32'hc4d8df8e, 32'h4409ff93, 32'hc14116ba},
  {32'hc3635df6, 32'hc551ca05, 32'h43f3d3dd},
  {32'hc42d1ac0, 32'h43ed495c, 32'h44f00802},
  {32'h443b4668, 32'h434bb138, 32'hc477060b},
  {32'hc4e45d0b, 32'h4410ca4e, 32'h44ad9a3d},
  {32'h43da3e98, 32'h44171537, 32'hc4021d3c},
  {32'hc23a2d78, 32'h44121a50, 32'h4480f3f8},
  {32'h43e98439, 32'hc482bfed, 32'hc4ec9342},
  {32'h42a52458, 32'h43470c7c, 32'h4518d172},
  {32'hc40a5382, 32'hc39995d2, 32'hc4258aab},
  {32'hc2b883c8, 32'h444a1861, 32'h44ffd5b3},
  {32'h43d02b5e, 32'hc3a61397, 32'hc4bf7e34},
  {32'h45019fce, 32'h43d6a49d, 32'hc344954d},
  {32'hc5257d4c, 32'h420ead95, 32'h43d8ba2a},
  {32'hc20377a8, 32'h427e9ba3, 32'h43c5d216},
  {32'hc2374a00, 32'hc44b4dd9, 32'hc3376125},
  {32'h441dbe7c, 32'h4383e253, 32'h4206c278},
  {32'hc538d065, 32'hc3241e50, 32'h4304ca29},
  {32'h442668aa, 32'h452c3534, 32'hc36cb2dc},
  {32'hc550d090, 32'hc38fd30c, 32'hc4382e18},
  {32'h4316aad3, 32'h44f9dab8, 32'h428a9701},
  {32'h413895ec, 32'hc2c9645f, 32'hc2a6c7bc},
  {32'h4532faeb, 32'h4275a7e2, 32'h434ad271},
  {32'hc3fa27be, 32'h43fa05f7, 32'h448bc3b9},
  {32'h4404b8fb, 32'h4438c8e2, 32'h44acaf2a},
  {32'hc40438e7, 32'hc4460238, 32'hc4959acd},
  {32'hc50b87aa, 32'h42b0b0cc, 32'hc2a11c48},
  {32'hc450ef41, 32'hc4212c45, 32'h441a3429},
  {32'h43451937, 32'h43e7bb25, 32'h451302d9},
  {32'hc2717e00, 32'hc364c66e, 32'hc35adedf},
  {32'h44bbe1ea, 32'h43917bf2, 32'h44a14ecf},
  {32'hc532f6b3, 32'hc3a18eee, 32'hc393cc7c},
  {32'h44b94a05, 32'hc3aa140b, 32'hc390cc94},
  {32'hc2a032a1, 32'hc3de7337, 32'hc4b376c3},
  {32'h43fbe4b5, 32'h449c0877, 32'hc21b2198},
  {32'hc3b97c2d, 32'h4173908a, 32'hc4ad41b5},
  {32'h456e851a, 32'h43a23ae4, 32'h4438b224},
  {32'hc44c0ab2, 32'hc4048e67, 32'hc529d57e},
  {32'h44cff75e, 32'hc2c89675, 32'hc36533f6},
  {32'h445e34a5, 32'hc2f00154, 32'h435336b0},
  {32'hc41a1510, 32'hc4d1519e, 32'h435d9226},
  {32'h448bc545, 32'h43e36338, 32'h447916e6},
  {32'hc38a2557, 32'hc4617682, 32'hc307c5c4},
  {32'h45527cdf, 32'h4321b729, 32'h408c8492},
  {32'hc50402a2, 32'hc49725d0, 32'hc126fe1e},
  {32'hc4a3c6f7, 32'h438ff93f, 32'hc3bd8432},
  {32'hc50b1b39, 32'hc3fd4da2, 32'hc3bcd0df},
  {32'h4493e4c0, 32'h43fcce6c, 32'h445ad33e},
  {32'h4386cce3, 32'h42c61c46, 32'h447c5f7b},
  {32'h42cced63, 32'h443223df, 32'hc48182b3},
  {32'hc41478ec, 32'h446a7d3f, 32'hc4d47278},
  {32'hc358353d, 32'hc34b5b89, 32'hc381c0d6},
  {32'hc3b6399c, 32'hc5118198, 32'h4251eaa8},
  {32'hc1401f20, 32'h442e1c0c, 32'hc272aafa},
  {32'hc4469360, 32'hc40f8405, 32'h43f2b2b2},
  {32'h41995d80, 32'h43378009, 32'hc374a4fa},
  {32'hc407d238, 32'h42baaa4c, 32'h441327cf},
  {32'hc4bdd760, 32'h4348163a, 32'hc387aba0},
  {32'hc366ca40, 32'hc3ff5a4d, 32'h44a07b4a},
  {32'hc3293a78, 32'h44869997, 32'hc518451f},
  {32'h448c7f56, 32'h420a2456, 32'h43de0537},
  {32'h42fc3660, 32'h453423ac, 32'hc3b6a778},
  {32'hc489f7f7, 32'hc485a849, 32'h4350578c},
  {32'h455f122a, 32'h437af133, 32'h442099b2},
  {32'hc4330fd7, 32'h441dbd2d, 32'h45090b48},
  {32'h44a4e37a, 32'hc3d3dfa1, 32'hc51630c5},
  {32'h44e269e9, 32'hc43d2495, 32'h43c394d4},
  {32'hc3ad6a45, 32'h453e6f6a, 32'h43dac626},
  {32'hc4bf6ef7, 32'hc30bf08d, 32'hc38f9165},
  {32'hc2f0132c, 32'h44f91edb, 32'h433fbbb4},
  {32'h440612d6, 32'hc4e797a2, 32'hc3b8183c},
  {32'hc4346a76, 32'hc2226613, 32'h411fead8},
  {32'h44554750, 32'hc3929c42, 32'hc41667f5},
  {32'hc32f2ba0, 32'h447b57c7, 32'h4447045e},
  {32'h453b4ce8, 32'h42bee16a, 32'h441767e4},
  {32'hc40b5e9a, 32'h44954f03, 32'h43c73657},
  {32'hc3d9e1dc, 32'hc54b5b60, 32'h41ccb0ba},
  {32'hc4901292, 32'hc2f70ee0, 32'h43741cd2},
  {32'h44d26cfa, 32'hc4919d01, 32'h42dfe15a},
  {32'hc41d455b, 32'hc3d46ba7, 32'hc5089748},
  {32'h441f7de5, 32'h43a606fd, 32'h43c9033f},
  {32'hc4dce3f9, 32'h43b54310, 32'h4318febb},
  {32'h4460ffd4, 32'h43e86035, 32'h43b18c8c},
  {32'h441aa740, 32'h4301485e, 32'hc4483c7a},
  {32'h44c4da34, 32'hc3f9bd77, 32'h439bff60},
  {32'hc4be9cba, 32'h43aeaa0d, 32'hc402f7cc},
  {32'h43f398b3, 32'hc3df2697, 32'hc3379ed1},
  {32'hc4c7c04d, 32'h4493b548, 32'hc3a89c6f},
  {32'h44b369ae, 32'hc3fabe7f, 32'h4381e58f},
  {32'h42b72ba5, 32'h4346e0a1, 32'hc3f185d4},
  {32'h4435ee7a, 32'h43bba352, 32'h4500dbe9},
  {32'hc4102b44, 32'hc48ba808, 32'hc544a276},
  {32'hc429c5ea, 32'hc2b97e70, 32'h43dc45c3},
  {32'h44248242, 32'hc43c0ee4, 32'hc4d09842},
  {32'hc32b026b, 32'h43745bc1, 32'h45311c7c},
  {32'hc4965381, 32'hc315e3ef, 32'h4404b258},
  {32'hc423b8b9, 32'h4365bc0d, 32'hc2e8ab33},
  {32'h45531d0e, 32'hc3f1f8c4, 32'hc36beda9},
  {32'hc3d07a02, 32'h4492b108, 32'hc4444dba},
  {32'h44fbe9dd, 32'h435961da, 32'hc0e028f4},
  {32'hc4150739, 32'h4368a93a, 32'hc55dfa90},
  {32'h449f165a, 32'hc38ce027, 32'h4448a3e8},
  {32'h43260921, 32'hc4edd022, 32'h44e14fea},
  {32'hc4fbf8c2, 32'hc1830374, 32'hc4af6855},
  {32'h4435bed9, 32'h42eabbfe, 32'h440c6eb4},
  {32'hc369e66e, 32'hc4845d04, 32'h43a82053},
  {32'hc44831dc, 32'h445edcf7, 32'h437777a1},
  {32'hc3a4be9a, 32'hc3ce1295, 32'h45533cd2},
  {32'hc1304230, 32'h4496097e, 32'h435db621},
  {32'h438e392c, 32'hc49b279a, 32'h44b4fd29},
  {32'hc3343320, 32'h44144003, 32'hc45d3da2},
  {32'h450324ca, 32'hc38dd0df, 32'h441297a8},
  {32'hc5678af1, 32'h42f4ba24, 32'h438bd937},
  {32'h4521db30, 32'hc38a7c52, 32'h4445d420},
  {32'hc550f4da, 32'hc3a9c8a7, 32'hc2f94fd6},
  {32'h450f880c, 32'h43c71f44, 32'h441a3d44},
  {32'hc4118eb4, 32'h44bf9777, 32'h4389c26c},
  {32'h449cf026, 32'hc443e5e2, 32'h4228e619},
  {32'hc440f01c, 32'h44b5c434, 32'h43e30621},
  {32'h433951a0, 32'hc570371e, 32'h43b2d4c7},
  {32'h42fa7ef8, 32'hc4a7bb3f, 32'h43af08be},
  {32'h429c2d3a, 32'h445bdb24, 32'hc4db0c72},
  {32'hc312010f, 32'hc48a7ef2, 32'h45451555},
  {32'hc3c30e7c, 32'h429f7d56, 32'h44230362},
  {32'h425e70a0, 32'h44873b8e, 32'hc4219a4a},
  {32'hc351c190, 32'h439379c4, 32'h44c490a5},
  {32'h444a4190, 32'h44174d9b, 32'hc486b8d4},
  {32'hc353f310, 32'hc4c311ab, 32'h4323b268},
  {32'h450bfa4d, 32'hc3c521e2, 32'h4418e481},
  {32'h43d689a4, 32'h448aaa26, 32'hc37dfd84},
  {32'hc42dc0f2, 32'hc319978f, 32'h44c9700a},
  {32'h4367af08, 32'hc46d16e5, 32'hc4d9d97a},
  {32'hc18c49bc, 32'hc30bcf68, 32'hc533959b},
  {32'hc3803675, 32'hc3cf85ab, 32'h4530c867},
  {32'hc393634c, 32'hc3c8be85, 32'hc4390da0},
  {32'hc28822f7, 32'hc527a8e2, 32'hc2f948a0},
  {32'h4420b642, 32'h446118a8, 32'hc426f36a},
  {32'h44c625dc, 32'h423c1691, 32'h443c72dd},
  {32'h450878d7, 32'hc3d29031, 32'h43a43ce4},
  {32'hc535ded0, 32'h42fdfbfa, 32'hc3482168},
  {32'hc36dd3b3, 32'h436f0bdd, 32'hc387fefe},
  {32'hc4c6b682, 32'hc495e39b, 32'h43aa239a},
  {32'h44e49485, 32'h4477811c, 32'h43765b0b},
  {32'h44ecc2a1, 32'hc30aff40, 32'h43bbe1a0},
  {32'h453aaf99, 32'h43f9491b, 32'hc3a87926},
  {32'hc4483390, 32'hc523394b, 32'h438d4a8a},
  {32'h44e0fefd, 32'hc1ddda21, 32'hc3f3e291},
  {32'h43aa2a5d, 32'hc4a1abc3, 32'h443440ee},
  {32'hc52c07d9, 32'h437b81a3, 32'hc2858d1e},
  {32'hc2097350, 32'h44b119c4, 32'h444c7b5e},
  {32'hc35499ae, 32'hc4aef008, 32'hc30db82c},
  {32'h430f65f4, 32'h438e0ccc, 32'h44e1cc97},
  {32'hc30d3a90, 32'hc42991da, 32'hc4297328},
  {32'h4395b287, 32'hc30ac06b, 32'h434521e8},
  {32'hc45ea588, 32'hc426d3a1, 32'hc49f6566},
  {32'hc384ef88, 32'h44d11cf4, 32'h45087b3a},
  {32'h43822e48, 32'h444e9157, 32'hc3bfc051},
  {32'h440ddb92, 32'h44b3afad, 32'hc2ca493c},
  {32'hc43c7b8a, 32'h44bb378e, 32'hc4acc59b},
  {32'hc498a04c, 32'h43be176f, 32'hc2a5b831},
  {32'hc4128550, 32'hc483bd89, 32'hc3dca43f},
  {32'h44900a94, 32'h44a02f4e, 32'hc2bae7d2},
  {32'h43cea84a, 32'hc38782e0, 32'hc52260c7},
  {32'h4532b104, 32'h437617aa, 32'h440bd0ab},
  {32'h42503764, 32'hc3d065fa, 32'hc4999a7d},
  {32'hc4b68530, 32'h43d9c535, 32'h43ba9a0a},
  {32'hc3b3965a, 32'hc5513f49, 32'hc395edfb},
  {32'h44de2963, 32'h44b4af17, 32'hc2e6715a},
  {32'h43da01c1, 32'hc4a75d6c, 32'hc4069816},
  {32'h43332dc4, 32'h450cf9d2, 32'h4321cfe1},
  {32'hc4f48338, 32'hc3ffdba2, 32'h428b799f},
  {32'hc4827667, 32'hc34db71b, 32'h421615c4},
  {32'hc5628634, 32'h437989e0, 32'h43a9b760},
  {32'h44b17854, 32'hc408b0c7, 32'h43ba08f3},
  {32'h41465240, 32'h43f92634, 32'hc50098fd},
  {32'h43bd896c, 32'h44d5bc52, 32'h445148ec},
  {32'h41b66d20, 32'h44258996, 32'hc3dbb68c},
  {32'h428dcdce, 32'h44e3871f, 32'h444b43d2},
  {32'hc1506c00, 32'hc4ac62e5, 32'hc3704901},
  {32'hc34e497e, 32'h4500d32a, 32'h43b709b3},
  {32'h43f37024, 32'hc481e9bb, 32'hc4d0ffca},
  {32'hc515941b, 32'h44163855, 32'h4423c314},
  {32'hc4745002, 32'hc4213b2b, 32'h4351fb5f},
  {32'h41fecede, 32'h449c9bfc, 32'h445f7d7e},
  {32'hc0b5e330, 32'h43a70b5e, 32'hc50fdd55},
  {32'h446c3f84, 32'h43c06694, 32'h43fa8fe6},
  {32'h43fbb450, 32'hc4214947, 32'hc4860f86},
  {32'hc30799e0, 32'hc336a66e, 32'h43b3403c},
  {32'h446d664a, 32'h42b3b894, 32'hc2878319},
  {32'hc2524af0, 32'h44a9d895, 32'h452e375a},
  {32'h44b7ed30, 32'hc2abfccb, 32'h427955c0},
  {32'h44e0eca5, 32'hc318fc8b, 32'h4338eb25},
  {32'h4372c7e0, 32'hc4e1f626, 32'hc39e3aca},
  {32'hc52afeef, 32'h43a09929, 32'h419e2e47},
  {32'hc385f253, 32'hc4878fd5, 32'h426f726f},
  {32'hc49c5376, 32'hc26921bf, 32'hc3b2aa15},
  {32'h44ab5e3b, 32'hc36fdaf7, 32'hc3d20383},
  {32'h44292aae, 32'h4416208c, 32'h43334e5b},
  {32'h44fec7a2, 32'h43460669, 32'hc228e1b3},
  {32'hc57ae36c, 32'h43cb4cb3, 32'hc3f01c60},
  {32'hc5014602, 32'hc2528f67, 32'h42a2a85c},
  {32'h44bcc968, 32'h4386c70b, 32'hc2d9df29},
  {32'hc49209c9, 32'h43b55fe1, 32'hc501b476},
  {32'hc2fcbe7a, 32'h431462b7, 32'h44bd86f5},
  {32'h44644cb3, 32'h41380569, 32'h4356320b},
  {32'hc3142368, 32'hc5370282, 32'h42e2e7f4},
  {32'hc40b1d60, 32'h44f45632, 32'h43cbdce6},
  {32'h43bbf967, 32'hc2e8c911, 32'h43466267},
  {32'hc58d36ef, 32'h40894075, 32'h43070310},
  {32'h44f22ece, 32'hc49aafe6, 32'hc3866b9d},
  {32'h44c56b2c, 32'h43053ca4, 32'hc4721326},
  {32'h4509c005, 32'h419707eb, 32'hc2a5dde5},
  {32'hc501cba5, 32'h44328aaa, 32'hc260245a},
  {32'hc3df7d10, 32'hc475a7c3, 32'h4235f71a},
  {32'hc3f2770b, 32'hc2a731ad, 32'h449af097},
  {32'h44bf1506, 32'hc29714f5, 32'hc4242085},
  {32'h430c4e46, 32'h444234cb, 32'hc314e651},
  {32'h438cdb18, 32'h43852811, 32'hc50f042e},
  {32'hc3c663f0, 32'h44713568, 32'h43d15a2b},
  {32'hc175fff8, 32'h40da6ae7, 32'hc40a4a0e},
  {32'hc4cf3042, 32'h442195e8, 32'h44756bfe},
  {32'h455439f6, 32'h43e6bfc0, 32'hc428943a},
  {32'hc3a45c77, 32'hc32313f0, 32'h443fb795},
  {32'h44d33335, 32'hc3a2b88c, 32'hc50332ef},
  {32'h443f4d51, 32'h452e9fb0, 32'h4387613d},
  {32'h431b0067, 32'hc4d72587, 32'hc39ca07c},
  {32'h42f24428, 32'h44da7fd3, 32'h4485e5ea},
  {32'h431102c8, 32'hc4663ac4, 32'hc51262da},
  {32'h43925f68, 32'hc3ac46c8, 32'hc48a7921},
  {32'hc4de7598, 32'hc36e8ac4, 32'h43da0f0a},
  {32'hc2ea83b0, 32'h437991a3, 32'h434be932},
  {32'hc3abc8bb, 32'hc54dbe83, 32'h431fc3b3},
  {32'h4489b9ad, 32'h43b615de, 32'hc3bd7be6},
  {32'h451d2fe4, 32'hc2a1ec0c, 32'hc3865acd},
  {32'h42f05a40, 32'h452c7117, 32'h42eb2bc3},
  {32'hc4d44d35, 32'hc490e57b, 32'h41af0f4d},
  {32'h4468a1ff, 32'h43d13840, 32'h43e8e6c3},
  {32'hc33bba28, 32'hc40047d5, 32'h45129df0},
  {32'h44f6e1ac, 32'h42ceace9, 32'hc42f6224},
  {32'hc134f9a8, 32'hc13483c1, 32'hc36372a0},
  {32'h41fb1e20, 32'h44f243e4, 32'h43c6d572},
  {32'hc44bc964, 32'hc442408e, 32'hc5243418},
  {32'h446c8f0f, 32'h42fd5773, 32'h441bafad},
  {32'hc3d2463c, 32'hc4e3223f, 32'h434e9be9},
  {32'h44953dfa, 32'h43ce826b, 32'h43fe594c},
  {32'h4451feac, 32'h432ec89f, 32'hc4564841},
  {32'h453bcc54, 32'h43f25ca4, 32'h43fb77fe},
  {32'hc4d120fe, 32'hc4342980, 32'hc4339656},
  {32'h4193cfe0, 32'h42df841a, 32'hc2916448},
  {32'hc36ab228, 32'hc4b2cce5, 32'hc4b0f953},
  {32'h4488fcc0, 32'h44879b51, 32'h43463b72},
  {32'h4463a04e, 32'h435da33c, 32'hc41452a8},
  {32'hc385ff4c, 32'h45365245, 32'h4386b292},
  {32'hc56a504a, 32'h431c0df1, 32'hc399e1db},
  {32'hc29e17a8, 32'h435a5c9e, 32'h42bcbe7e},
  {32'h44422f87, 32'h44294387, 32'hc2b229de},
  {32'hc3e78334, 32'hc4235807, 32'hc43d9338},
  {32'h449a3fc8, 32'h4418982f, 32'h43a9c00a},
  {32'hc492726b, 32'hc330fc65, 32'h41a59567},
  {32'h44db7b5a, 32'hc29372f1, 32'hc3bab555},
  {32'hc4eef26b, 32'hc47cf2a3, 32'hc2cbfb0f},
  {32'hc4a7c647, 32'h438e8a4e, 32'h41e22152},
  {32'hc4057a40, 32'hc4b35bff, 32'hc4a96be3},
  {32'hc355ffd0, 32'hc423f020, 32'h43957be4},
  {32'hc4eaffb0, 32'hc39f8454, 32'h43ce4729},
  {32'h43300190, 32'h444926b1, 32'hc4565981},
  {32'hc5273745, 32'hc22cf55e, 32'hc32b42ba},
  {32'hc4206948, 32'h43159310, 32'hc3858df4},
  {32'h43926ee4, 32'hc3c7dc81, 32'h45202547},
  {32'h44148ef2, 32'h44aeb3ae, 32'hc3dfd264},
  {32'h444b4a4a, 32'hc31da2cc, 32'h43b54faf},
  {32'h4495ba91, 32'h4363534e, 32'hc3ea3ed4},
  {32'hc41a434b, 32'h431abfcd, 32'h44df98d1},
  {32'h44aff54a, 32'hc3a4c826, 32'hc3f09454},
  {32'hc4d99e84, 32'hc482f57f, 32'h441f5032},
  {32'h44267294, 32'h42911282, 32'hc2a771eb},
  {32'h4511c1ff, 32'h43bc4a9c, 32'hc3240075},
  {32'hc3df7e8a, 32'hc292d930, 32'h4516a106},
  {32'h44e8b27b, 32'h43849223, 32'hc1b3f2ba},
  {32'hc51350bf, 32'h43c1be25, 32'h44c2dead},
  {32'h453831f9, 32'hc3f0179b, 32'hc48b6762},
  {32'h4344c318, 32'hc51e184d, 32'hc2a9faa5},
  {32'hc487a256, 32'h444ec40a, 32'h43fe4c6e},
  {32'h4501ee4d, 32'hc2369444, 32'h440d0939},
  {32'hc4498770, 32'h450df350, 32'h43ebafd8},
  {32'h449da5f9, 32'hc347e874, 32'hc3937958},
  {32'hc4ee12cf, 32'h42700738, 32'hc3ad01da},
  {32'h445ab718, 32'hc30310bc, 32'h4192100b},
  {32'hc58aee9a, 32'h43469c68, 32'h442eba29},
  {32'h453f1788, 32'hc263fb28, 32'h439969d1},
  {32'hc3223657, 32'h44409fcb, 32'h43597057},
  {32'h4482a9e0, 32'hc42161be, 32'h44732975},
  {32'h44686af7, 32'hc3c1d910, 32'h42171927},
  {32'h43b11f0a, 32'hc2756616, 32'h45083586},
  {32'hc479f361, 32'h441635b2, 32'hc37334f2},
  {32'h43f08bba, 32'h426905b8, 32'h40aad044},
  {32'hc4db3d78, 32'h42d7f144, 32'hc3c8f971},
  {32'h452a8508, 32'h43c851e6, 32'h4360ec3a},
  {32'hc4e23159, 32'h439d5033, 32'h43b39ed8},
  {32'h450f2390, 32'hc4264d31, 32'h440be7f0},
  {32'hc2d8ae44, 32'h44fc7eb6, 32'hc4802ed7},
  {32'hc3860465, 32'hc42be54b, 32'h4409e120},
  {32'hc381b492, 32'h4496b283, 32'hc3067b44},
  {32'hc3ce785c, 32'hc486d8ab, 32'h43e30911},
  {32'h43a45b2c, 32'h42b3fcd7, 32'hc2e8000c},
  {32'h44e403a6, 32'h437aae8e, 32'h4474cc3e},
  {32'hc4fb8c77, 32'h440e9467, 32'hc44ca840},
  {32'h4553f3f5, 32'hc29455a0, 32'hc3e1e95f},
  {32'h43adcb16, 32'h44966711, 32'hc4b8edf1},
  {32'hc495a78c, 32'hc3a12d2c, 32'h44c37d34},
  {32'h43b54be7, 32'h4485d024, 32'hc45ce4b8},
  {32'h44fadf52, 32'h43a45948, 32'hc367cddf},
  {32'h44ad6dd8, 32'hc4dd04ca, 32'hc3e20a91},
  {32'hc44bcea9, 32'h445b0be4, 32'hc393ec7a},
  {32'h42a2b39c, 32'h4400e6ec, 32'h4500e5b5},
  {32'h41893f8e, 32'hc36be984, 32'hc5064f0c},
  {32'h4454b67f, 32'hc4dab33a, 32'h43afdfd6},
  {32'h44bc04f4, 32'hc3cdda41, 32'h446eccd7},
  {32'h43d81aed, 32'h44fe1b5e, 32'hc501089a},
  {32'h44a054ef, 32'hc3fd2b53, 32'h42ba1f88},
  {32'h43515e3e, 32'hc224736b, 32'h44b69a57},
  {32'hc3b3d9f9, 32'hc2088d47, 32'hc4d08d35},
  {32'h43e315d2, 32'hc3253cdc, 32'h4489d76c},
  {32'hc51a8746, 32'hc341a800, 32'h42ce3573},
  {32'h449e2795, 32'h4308970b, 32'h443369d4},
  {32'hc408581e, 32'h430021dc, 32'hc4a6a492},
  {32'h452c00a4, 32'h42239db2, 32'h440f1dd2},
  {32'hc550df18, 32'hc3b8ff40, 32'hc404e3d4},
  {32'hc373e200, 32'h43e093ab, 32'h43e4f586},
  {32'hc53c4b71, 32'h421b335a, 32'hc25b7c28},
  {32'h451516fb, 32'hc483b8c8, 32'hc36706e7},
  {32'hc4f89ab9, 32'h4389e7e6, 32'hc30ced4a},
  {32'h449fcff0, 32'h43cc4f56, 32'h43ddb9a4},
  {32'hc4642067, 32'h451fc75f, 32'hc3c74c3f},
  {32'hc19025e0, 32'hc55645b0, 32'hc3d2a364},
  {32'hc2b72964, 32'h43260e8a, 32'h4412522e},
  {32'h4340dfe6, 32'hc404cec3, 32'hc45dee36},
  {32'hc31817fa, 32'h43c2ef5a, 32'h44c94a32},
  {32'h42d3f238, 32'hc32c31c5, 32'h453b3de5},
  {32'h43a41841, 32'h44d5cf02, 32'h42b2d15f},
  {32'hc4d2376a, 32'hc43c3ff2, 32'hc334fcb0},
  {32'h43cbb014, 32'h42959599, 32'hc4abca52},
  {32'hc519b833, 32'h42be6bf6, 32'h42f36ddd},
  {32'hc2841a78, 32'h44b348d1, 32'h4308f056},
  {32'hc30c20b8, 32'h442bfc8e, 32'hc4a28b92},
  {32'h43a4e98c, 32'h439db95b, 32'h455421d5},
  {32'hc33f4064, 32'hc23658b4, 32'hc4bb94d9},
  {32'h431cc2b8, 32'hc3fb0215, 32'hc3cf59f1},
  {32'hc4448915, 32'hc390720b, 32'hc3e06d0c},
  {32'h444852a4, 32'hc3048ba8, 32'h42adaaa3},
  {32'hc33572a3, 32'h427e6829, 32'h44d92e36},
  {32'h449817e5, 32'h43b0bbf0, 32'h41ef4b2a},
  {32'hc502e258, 32'hc31558b1, 32'hc35fa374},
  {32'h45364bd6, 32'hc39297a8, 32'h4330b644},
  {32'hc4702dc4, 32'hc2a847e3, 32'hc3968d58},
  {32'hc4312fdf, 32'h41c07d48, 32'h42554a9c},
  {32'hc4aaf4ac, 32'hc4881a44, 32'h43ac6340},
  {32'h441b4f77, 32'h44fd98d6, 32'h43b608a8},
  {32'hc30b2050, 32'hc38d28f1, 32'h4289d928},
  {32'h41dabe60, 32'h45763231, 32'h4304ae4d},
  {32'hc4922f44, 32'hc4a5c8fc, 32'h432f2b78},
  {32'hc4e20e8b, 32'hc22ddfc8, 32'hc2e881e0},
  {32'h43cca05e, 32'h435e8516, 32'h441dcfd1},
  {32'h44081646, 32'h44d14e3d, 32'hc4c0d419},
  {32'hc37f9ffe, 32'hc4176ba2, 32'h44ff16ed},
  {32'hc1d55620, 32'hc49a6607, 32'hc3a5b9f3},
  {32'h42ab227c, 32'h453d010d, 32'h441d66f2},
  {32'hc335b8aa, 32'h43007766, 32'hc4972e9d},
  {32'hc1bcd220, 32'h42cfb405, 32'hc1d7186d},
  {32'hc4507acf, 32'hc4931557, 32'hc4179167},
  {32'h42dbf780, 32'h445b23b1, 32'h45206c5a},
  {32'h441bdc85, 32'hc46e88a7, 32'hc3c7549c},
  {32'h43008abc, 32'hc354b19e, 32'h449d4688},
  {32'h44179277, 32'h42f07bbb, 32'hc3f32c07},
  {32'h44ec8f42, 32'h4339aad2, 32'h4379be49},
  {32'hc42263ed, 32'hc311ab2b, 32'hc4d739f4},
  {32'h44bbd53f, 32'h444adda7, 32'h4271e123},
  {32'h44ba4589, 32'hc43641f9, 32'hc37a5754},
  {32'h440ca4b6, 32'h44b6bb03, 32'h447016ea},
  {32'hc22960d0, 32'hc3ee0136, 32'hc5656a5b},
  {32'hc28469e8, 32'h44d4b701, 32'hc3a10be8},
  {32'hc431dddc, 32'hc4b2c1db, 32'hc3f6558d},
  {32'hc3d95ad8, 32'h454f1c15, 32'h441bbea2},
  {32'hc4ab0c0b, 32'hc316199d, 32'hc1e66ccf},
  {32'hc32acd1c, 32'h454e9908, 32'h430e6d7c},
  {32'hc4fbfa6a, 32'hc40d2410, 32'h420706dc},
  {32'hc4e6e3cc, 32'h42261b73, 32'hc2a65a05},
  {32'hc53f30d8, 32'h43cabc08, 32'hc3f4ac65},
  {32'h45417d0f, 32'hc1f71244, 32'h43eb058d},
  {32'h4322ccec, 32'hc4b81fac, 32'hc4146755},
  {32'h43c05225, 32'h44aadacf, 32'h444677fe},
  {32'h420c5748, 32'hc34a0131, 32'hc3cb2a24},
  {32'hc4edbec4, 32'h445f4f47, 32'hc3417fc7},
  {32'hc3732686, 32'hc42002c4, 32'hc4d89941},
  {32'hc4d04d60, 32'h43b78b79, 32'h43db279c},
  {32'h441fa063, 32'hc11e2270, 32'hc4a0d86d},
  {32'hc4ac6c00, 32'h42126f2b, 32'h44824480},
  {32'hc3f01a58, 32'hc43fab12, 32'hc3174883},
  {32'hc347ab39, 32'hc4a6f67a, 32'h45151d95},
  {32'hc39b1af9, 32'h44adf4ef, 32'hc50c757e},
  {32'h43db18c6, 32'h44ca128c, 32'h43764bc1},
  {32'h4330d8d8, 32'hc4aa4f1c, 32'hc39c7b7c},
  {32'hc38a7910, 32'h44a01cd0, 32'h431d7f4e},
  {32'hc481e32b, 32'hc2e8c70a, 32'hc3732fa8},
  {32'hc2b1a0de, 32'h44591d64, 32'h44d9147a},
  {32'h446c7912, 32'hc37f510c, 32'hc41feffa},
  {32'h441a79f9, 32'h446422f8, 32'h443d0104},
  {32'h446b87b2, 32'hc5288f76, 32'hc2ef4f48},
  {32'hc4f02396, 32'h442c8ed4, 32'h4285b700},
  {32'hc05d2c78, 32'hc2452901, 32'h4377245c},
  {32'hc48544f2, 32'h450ff213, 32'h43206dc8},
  {32'h43fe9091, 32'hc439f303, 32'hc0ed1cf1},
  {32'hc4b920a6, 32'h441085cf, 32'h430a38a2},
  {32'h44bcbfda, 32'h4381c0bf, 32'h43ce71c6},
  {32'hc5782792, 32'h434e85f8, 32'hc3be8328},
  {32'h4510217d, 32'hc20ffd05, 32'h42df8c49},
  {32'h44b4e1b8, 32'h42931ced, 32'hc40cdf9c},
  {32'hc4bd3f3e, 32'h43521b69, 32'hc4308a89},
  {32'h455620e7, 32'h43746695, 32'h435af231},
  {32'h44550ef7, 32'h43ce1fce, 32'hc2cb9789},
  {32'h447d3636, 32'hc4727a1f, 32'h43bd7ba9},
  {32'hc4e11a6c, 32'h4463dbcf, 32'h435cb372},
  {32'hc3ce4df9, 32'hc444ff45, 32'h4311ab28},
  {32'hc4ecb5e6, 32'h449ac536, 32'hc2586e8c},
  {32'h4432fda7, 32'hc50fa756, 32'h438643fa},
  {32'hc43c453d, 32'hc2fa299a, 32'hc45db50b},
  {32'h45345bc6, 32'h4346c9dc, 32'h42a3eb2c},
  {32'hc4ea87c6, 32'hc44b51dc, 32'hc3891ab3},
  {32'h448b732d, 32'hc1fc3ff4, 32'hc3777fd5},
  {32'hc33ff7be, 32'h44fe4704, 32'hc2313709},
  {32'hc336a239, 32'hc503c13b, 32'hc47307ed},
  {32'hc427997e, 32'h44008f3f, 32'h43541046},
  {32'h449301ec, 32'h4394978c, 32'hc4e01eb5},
  {32'hc3bb6f35, 32'h443872cd, 32'h44d29caa},
  {32'hc47a6044, 32'hc3e9aea6, 32'hc207870b},
  {32'hc4ed1b87, 32'h43c757e8, 32'h445114ea},
  {32'hc3440550, 32'h449f7a97, 32'hc47e6233},
  {32'hc258dd28, 32'h44bd24b4, 32'h43a9a68d},
  {32'h42ab3231, 32'hc45047fe, 32'hc5193e42},
  {32'hc533f74e, 32'h42123c78, 32'h440332b3},
  {32'h4369710c, 32'hc43dfd12, 32'hc42b6227},
  {32'hc54f1840, 32'h447ee961, 32'hc2990d05},
  {32'h448d8075, 32'hc3a66634, 32'hc4ea8600},
  {32'h45597a14, 32'hc32e3288, 32'hc44bb936},
  {32'hc5653ec8, 32'hc2bb39aa, 32'h43219051},
  {32'hc44dce3e, 32'h443824fd, 32'hc42e2df6},
  {32'hc3b39d68, 32'hc4f15d71, 32'h42d6a3f7},
  {32'h44a2173d, 32'h44497b22, 32'hc3a01188},
  {32'hc4cb6a12, 32'h4386decc, 32'hc3cc6796},
  {32'h453fad46, 32'h44017724, 32'h43832437},
  {32'hc483d1c3, 32'hc4c70e1d, 32'hc057cae0},
  {32'h43989f72, 32'h41310e77, 32'h440f065e},
  {32'hc31b57cf, 32'h4377bb9a, 32'h447af697},
  {32'h4426e6c5, 32'h440063d2, 32'h43957cfa},
  {32'hc389f43a, 32'h43ddbb22, 32'h42fdd9ae},
  {32'h439abc02, 32'h43e9942f, 32'h452054b0},
  {32'h43545968, 32'hc42ecb5a, 32'hc4c397d1},
  {32'h44c3cfdd, 32'h43390b53, 32'h439adfa9},
  {32'hc479eb65, 32'hc1e47bf9, 32'hc4ecc1c0},
  {32'h442f0f5f, 32'h449724cf, 32'h44b26a3a},
  {32'h42c33662, 32'hc1ffb9a4, 32'hc4e25776},
  {32'h452a26b5, 32'hc402d996, 32'h438922a4},
  {32'hc513a5ab, 32'hc390796f, 32'hc411f10a},
  {32'h45483174, 32'h43d8170f, 32'hc3cb49a4},
  {32'hc31422f0, 32'hc4577ea8, 32'hc4b2f4e5},
  {32'h43352d7a, 32'h4504b58d, 32'h43ae9440},
  {32'hc4da85ec, 32'hc3589cfe, 32'h438bc66d},
  {32'hc2ad5eba, 32'h44b0a724, 32'h42cd471a},
  {32'h435729cd, 32'hc4a07b02, 32'hc4d8b85f},
  {32'h452218b1, 32'hc20c308f, 32'hc3b8b14e},
  {32'hc4edf5e6, 32'hc29fd150, 32'h42ec4021},
  {32'hc41a3bda, 32'hc4c86a3b, 32'h430a131a},
  {32'h42966e04, 32'h44e67bb6, 32'hc3b10b9d},
  {32'hc50139d6, 32'h428bcf9d, 32'h4359419d},
  {32'h44c389e5, 32'h44973504, 32'hc384b096},
  {32'hc51cca5e, 32'hc438c2fc, 32'h43a80313},
  {32'hc41dcf9c, 32'hc381b150, 32'h40b98e96},
  {32'hc53c8c42, 32'hc12f55f8, 32'hc33b469c},
  {32'h444f1262, 32'h441e4027, 32'h44840953},
  {32'h43e0f94f, 32'hc49a3c1a, 32'h44b21c86},
  {32'h449f7d8e, 32'h441a52ac, 32'hc326e139},
  {32'hc4c73109, 32'hc33857e5, 32'h432a53bc},
  {32'h449aabf5, 32'h43c22e63, 32'hc2523f7a},
  {32'h433ac8d8, 32'h4299c885, 32'h45612f1f},
  {32'h4447f88c, 32'h451b21bc, 32'hc3a7ee58},
  {32'hc4b4ef6f, 32'hc29cc578, 32'h4374456f},
  {32'h44ff2f38, 32'h43db7a14, 32'hc3783210},
  {32'hc47b6530, 32'h43d89491, 32'h43818f2f},
  {32'h451966b4, 32'hc3acd8d2, 32'hc3ab0d27},
  {32'hc3a59ad6, 32'hc4aaf549, 32'h4480a296},
  {32'hc4a705c1, 32'h42fb3151, 32'h412dac1d},
  {32'h44ddd6da, 32'hc310eeb7, 32'hc38ed99f},
  {32'hc354a073, 32'hc4ac46c0, 32'h43ad4d38},
  {32'h43d853ee, 32'hc2e9e5ed, 32'hc5081985},
  {32'hc48d2c35, 32'h43373911, 32'h44a67b3d},
  {32'h43c15a38, 32'hc3a294af, 32'hc517b191},
  {32'hc2619be0, 32'hc516f13b, 32'hc28db6ae},
  {32'hc3d25b36, 32'h43d2bcc3, 32'h44c7fb1c},
  {32'h44438e20, 32'hc3defdaa, 32'hc31f494d},
  {32'hc403f624, 32'h44923459, 32'hc400acc8},
  {32'h4419d302, 32'hc3a122da, 32'h437afa4c},
  {32'hc39ebdde, 32'h44a02c49, 32'hc2fe0142},
  {32'h43730dc0, 32'hc4a4f5e5, 32'hc483ae1a},
  {32'hc41ca144, 32'h44a079af, 32'h44a8dcea},
  {32'hc4acdcde, 32'h42e68c64, 32'h43864e9b},
  {32'hc4e51bee, 32'hc38ff117, 32'h427d2641},
  {32'hc29acf98, 32'hc4aa1d60, 32'h439bd549},
  {32'hc4a42854, 32'hc2befbc4, 32'hc3e503c3},
  {32'h44a53cbf, 32'hc2655e17, 32'h4424079a},
  {32'hc42a9228, 32'h43e60907, 32'hc443831e},
  {32'hc307cf93, 32'hc4ed9731, 32'hc37d5ba3},
  {32'hc3dca67c, 32'hc3fd461f, 32'hc444e77a},
  {32'h454d7ac7, 32'hc3d395a8, 32'h3f803a38},
  {32'hc4868683, 32'h41faa4b2, 32'h4386cd32},
  {32'h445e49aa, 32'hc49166c8, 32'h43739d40},
  {32'hc3ea2e55, 32'h445bec58, 32'hc4686a75},
  {32'h44625df8, 32'hc3637e79, 32'h447a4df5},
  {32'hc4217a43, 32'h43a19877, 32'hc4215300},
  {32'h44ded2b4, 32'h426fe868, 32'hc327e43f},
  {32'h448fcdcd, 32'h43b7f037, 32'hc45b8878},
  {32'h43037ab0, 32'h43e3eb9e, 32'h44d308b0},
  {32'hc544b399, 32'h43567374, 32'hc4807d98},
  {32'h44f8f588, 32'hc3c4eb1f, 32'hc36c765e},
  {32'hc3d5cf85, 32'h43fa36f4, 32'hc45db970},
  {32'h4484fbde, 32'hc4788046, 32'h43087ab3},
  {32'h44a23525, 32'hc403e65e, 32'hc3b8b91a},
  {32'h42facb2e, 32'h4364dd98, 32'hc4dfa69f},
  {32'h4355e1d6, 32'hc4953d8c, 32'h4441cc50},
  {32'hc407e57c, 32'h43fdb342, 32'hc48316d6},
  {32'h434606ca, 32'hc3b81ca4, 32'h44804bd1},
  {32'hc48ad0cf, 32'h4449dbf3, 32'hc3e5b8d7},
  {32'h441b244a, 32'h4384f080, 32'h446784bd},
  {32'h45131bba, 32'h444d1edc, 32'h4496946a},
  {32'h42f5e112, 32'hc5035665, 32'hc4ea6b2a},
  {32'h44d8dec8, 32'h433d0d28, 32'hc3545400},
  {32'h42eb60e3, 32'hc1dc3b01, 32'h45120ad7},
  {32'hc45a8dc4, 32'hc333cdab, 32'hc4462d08},
  {32'hc2b87320, 32'hc49882b5, 32'hc27fb16f},
  {32'h44b8428b, 32'h431eff96, 32'h43ce319a},
  {32'h44c051fe, 32'hc455db55, 32'hc2fa493d},
  {32'hc44a347f, 32'h434f06e9, 32'hc49ae9b4},
  {32'hc4191ef3, 32'hc4116e4d, 32'h43165176},
  {32'hc49488f8, 32'h42572f3a, 32'hc3c3b200},
  {32'h45231ece, 32'hc3cb04e7, 32'h439d69cc},
  {32'h4430fd7b, 32'h447ed364, 32'h43981e24},
  {32'h44e0cf5c, 32'hc2c90da1, 32'h43a1a074},
  {32'hc3357654, 32'h4529e08e, 32'h429700ed},
  {32'h441066c4, 32'hc49b0ed7, 32'hc3b70980},
  {32'hc350c690, 32'h4528f693, 32'h43571790},
  {32'h442358be, 32'hc4974fd8, 32'hc3b34908},
  {32'h448e7a42, 32'hc3f8dae5, 32'h44052606},
  {32'hc3d1ebbe, 32'h44ca21c6, 32'hc50455a5},
  {32'hc4b76210, 32'h43c01be0, 32'h43ae2241},
  {32'hc448a3fa, 32'hc4c1fc5d, 32'h436f1f88},
  {32'h43dbc00c, 32'h42c77f6e, 32'h4046c870},
  {32'h43475b9c, 32'hc413bab1, 32'hc28273be},
  {32'h44e1fb45, 32'h439f52d2, 32'hc43a0bf2},
  {32'hc487a4f8, 32'hc3f20ef3, 32'h43bfeb46},
  {32'hc3534efd, 32'h45000a39, 32'h4391982c},
  {32'h4449cf9a, 32'hc30777bb, 32'hc3ba44b8},
  {32'h4320ba23, 32'hc3348906, 32'h44d4b218},
  {32'h435ebdb0, 32'h44c37070, 32'hc4d997fa},
  {32'h43e12290, 32'h44adb785, 32'hc3479c21},
  {32'h4198dd80, 32'hc4977752, 32'h44082bc3},
  {32'h44507300, 32'h43663bc9, 32'hc3a432ea},
  {32'hc49f54d3, 32'hc48a0f63, 32'h4379e860},
  {32'hc33fddff, 32'h443e0d71, 32'hc51087cc},
  {32'h44c26e5a, 32'h43623780, 32'h4416d928},
  {32'h449ec533, 32'h4357a12c, 32'h41e2009c},
  {32'hc574dc83, 32'hc1f9af7a, 32'h408d43ce},
  {32'h442774e8, 32'h43948183, 32'hc3fd69ad},
  {32'hc23f0ee0, 32'hc5645732, 32'h4227dbaa},
  {32'h440719b3, 32'h453c1c1f, 32'h41c2401b},
  {32'hc4a702d5, 32'h42127316, 32'h4402e4fb},
  {32'h4489899a, 32'h44cafea5, 32'hc3304a94},
  {32'hc4831f60, 32'hc4ca649b, 32'h42bd1153},
  {32'h45562f94, 32'hc40331c7, 32'hc2ec5b42},
  {32'hc1f4f5d0, 32'hc4a224d8, 32'hc0aea980},
  {32'hc5011aab, 32'hc13b0234, 32'h437a4635},
  {32'hc2fc0d37, 32'hc448fd87, 32'h4484265c},
  {32'hc4de8e03, 32'hc211b78a, 32'hc394840b},
  {32'h441b95d8, 32'hc18d459a, 32'h45072de2},
  {32'h439557a3, 32'hc3f2dc1b, 32'hc4c25ac4},
  {32'hc49abee3, 32'hc35023ed, 32'h429ee6e1},
  {32'hc423d4dc, 32'hc4056aca, 32'hc4cff185},
  {32'hc38da539, 32'h443cecc7, 32'h4581543a},
  {32'hc4c6df2a, 32'hc396cb90, 32'h4390c813},
  {32'h44169a03, 32'hc427db77, 32'h43af61d6},
  {32'hc18bcea4, 32'hc5282234, 32'hc3f53096},
  {32'h456359b5, 32'hc26d1b6e, 32'h4277758b},
  {32'hc16f4110, 32'hc30fc3c3, 32'hc54466ed},
  {32'h42e97a58, 32'h44d37320, 32'h4403bde6},
  {32'hc42d2900, 32'hc239e6c2, 32'hc3775859},
  {32'h44c4562e, 32'h442005e6, 32'h438e8fca},
  {32'hc4433809, 32'h43a7980a, 32'hc4888c75},
  {32'h4461ced9, 32'hc31fcf73, 32'h43bb2adf},
  {32'hc4c9f41b, 32'hc4af24ea, 32'hc2d27a0c},
  {32'h449d1f10, 32'h44c24d88, 32'h44277aee},
  {32'h43242910, 32'hc4f535a0, 32'hc31942b1},
  {32'h43759890, 32'h451abd89, 32'h41cdb6c2},
  {32'hc40c1485, 32'hc51d81b6, 32'hc2f4cd50},
  {32'hc3f1ed22, 32'h42cf109e, 32'hc3c634a9},
  {32'hc56abe28, 32'hc27f2164, 32'hc3261ada},
  {32'hc2bca580, 32'hc41aab53, 32'h43a71616},
  {32'h43500380, 32'hc49fbdcb, 32'hc48ca832},
  {32'hc3ae85c0, 32'hc4cd206a, 32'h44f4484e},
  {32'h44306bcc, 32'h42a2dd13, 32'hc443a016},
  {32'hc42b92c2, 32'h43ee4377, 32'h40a26f1a},
  {32'h431c236f, 32'hc5386001, 32'hc4012c4d},
  {32'hc4fb3fa7, 32'h43b43c12, 32'h43e42312},
  {32'h428a9620, 32'hc3af2bf6, 32'hc51869e1},
  {32'hc250352e, 32'h442ccff8, 32'h454160ce},
  {32'hc3373cba, 32'hc48e3a8c, 32'hc44312b1},
  {32'hc4a316ee, 32'h44388e6a, 32'hc3732622},
  {32'h427e431c, 32'hc401198c, 32'hc4c188d7},
  {32'h44616ec4, 32'h4402fa1d, 32'h43ab8436},
  {32'h442be698, 32'hc42cffae, 32'hc46172fb},
  {32'hc3005d24, 32'hc305561b, 32'h45596dd2},
  {32'h4510bb97, 32'hc3677b76, 32'hc4159531},
  {32'hc4c5365c, 32'h441bc1eb, 32'h43c6698d},
  {32'h4209c334, 32'hc49d4f0f, 32'hc5001ef8},
  {32'hc40fc5cb, 32'h43930107, 32'hc3a51de9},
  {32'h4547b32e, 32'hc442b981, 32'hc2470281},
  {32'hc4eab0f0, 32'h44286de9, 32'h439d6087},
  {32'hc4755851, 32'hc3b78269, 32'hc3680f0b},
  {32'hc50677b8, 32'h44368171, 32'hc33f0e1c},
  {32'h453d55d0, 32'hc2ef19ee, 32'h43829fbc},
  {32'hc46ab8ae, 32'h441bf896, 32'h42488a76},
  {32'h4549797e, 32'hc3e928b0, 32'h41ee07ea},
  {32'hc4976c13, 32'hc38f92bf, 32'hc34e5949},
  {32'hc40aa1de, 32'hc3958148, 32'hc43b1bc1},
  {32'h453818a6, 32'hc36a951d, 32'hc3a50a33},
  {32'hc4935d3c, 32'h4329172c, 32'hc4800141},
  {32'h4528442c, 32'hc31b6afa, 32'h4421fe29},
  {32'hc494b382, 32'h429523c8, 32'hc46ba9c8},
  {32'h42a937d8, 32'hc52895aa, 32'hc3838ecd},
  {32'hc50cf869, 32'h428fa4fd, 32'hc2ee0ba0},
  {32'hc4d4da38, 32'h43092f76, 32'h4221622a},
  {32'hc4c2d56d, 32'h4495f063, 32'h4221de75},
  {32'h434c393c, 32'hc5463d8a, 32'h4008df80},
  {32'hc31d300c, 32'hc35a6fa2, 32'hc4d11152},
  {32'h4307a900, 32'h42dfa902, 32'h4409a704},
  {32'hc4432a2e, 32'h43a31212, 32'hc481d289},
  {32'h447b72b2, 32'hc37ec80e, 32'h4375ec0d},
  {32'h434eaf1c, 32'h44abfce7, 32'h448c990e},
  {32'h44b556e4, 32'hc402550d, 32'hc4807f7e},
  {32'hc4bc0382, 32'h43c38f23, 32'h43b7607a},
  {32'h4527184f, 32'h436ebd10, 32'hc332c6b7},
  {32'hc33e9195, 32'h4495150f, 32'h441e8395},
  {32'h4506c455, 32'hc20e6c5d, 32'h43bee4b3},
  {32'hc57559d7, 32'hc2bb959e, 32'hc30cac31},
  {32'h44963c38, 32'h445e275a, 32'hc4afa972},
  {32'h43dbc50f, 32'hc28e1ae6, 32'h4378ea16},
  {32'h42848358, 32'hc4a87492, 32'hc46634e4},
  {32'hc3cb6baa, 32'h435b86e7, 32'h446a0dc8},
  {32'hc35ac48e, 32'hc321eb2d, 32'hc4ddee6f},
  {32'hc3efc300, 32'h450fe5dd, 32'h4423a76e},
  {32'h448c2d71, 32'hc429ed40, 32'hc4a51161},
  {32'h44d8716a, 32'hc38f8fd5, 32'hc49f54bc},
  {32'hc48e5ada, 32'h431ca339, 32'h43af2438},
  {32'hc3cc5296, 32'hc22a7d5a, 32'hc4453dff},
  {32'hc3e544ee, 32'hc3f6483d, 32'hc3ded5af},
  {32'h44b5161f, 32'h4470df54, 32'h441b8559},
  {32'hc3f88f93, 32'hc3f85b88, 32'h4159f3d0},
  {32'hc33687f0, 32'h454e347a, 32'hc2936dca},
  {32'hc4adcfcc, 32'hc462a46f, 32'h43a8e6bc},
  {32'h43203e13, 32'h44db76ce, 32'h42cbf405},
  {32'hc3c7c607, 32'hc438457a, 32'h453564f5},
  {32'h443b4eda, 32'hc3479b16, 32'hc276d51f},
  {32'hc410565e, 32'hc1c954e0, 32'hc2fb04b5},
  {32'hc18317c0, 32'h43901f27, 32'h4532e119},
  {32'h42e4f518, 32'hc4261458, 32'hc44fa15f},
  {32'h44dd3438, 32'h43ce6f51, 32'h42adddde},
  {32'hc31160ec, 32'hc48e9a3e, 32'hc33c7bfa},
  {32'h44a439e5, 32'h444c6ee5, 32'hc2487239},
  {32'hc2dbe010, 32'h430fa2f7, 32'h428b30a8},
  {32'hc31ffc70, 32'h41e6d3b2, 32'h44128ae6},
  {32'hc45fd5e2, 32'hc395e9ab, 32'hc42e9b17},
  {32'h44d8e837, 32'h4474bfd2, 32'h42d068e3},
  {32'hc2fe6850, 32'h44001134, 32'hc53a0622},
  {32'h43b841b8, 32'h449c4ba2, 32'h446991c5},
  {32'h44039407, 32'hc3a715cc, 32'h43f35aa2},
  {32'hc342f100, 32'h4448a48e, 32'h44b11bef},
  {32'hc4bbca5c, 32'hc3501b70, 32'hc3db1b22},
  {32'hc3fce7ee, 32'h4396e2f0, 32'hc3ae826a},
  {32'h443ab86c, 32'h43ca423b, 32'hc3ed7d0b},
  {32'hc5391601, 32'hc3bcf822, 32'h437f84ec},
  {32'h441b290f, 32'h44be872d, 32'h443618ba},
  {32'h446d3558, 32'hc332149b, 32'hc2934fbf},
  {32'h45159131, 32'h435a4457, 32'hc365d2a0},
  {32'hc4026305, 32'hc4a9dd66, 32'h4459b003},
  {32'h445ad7f5, 32'h43845d36, 32'h4417e128},
  {32'hc563adf0, 32'h43ff4a8d, 32'hc3aafd40},
  {32'h455e65a8, 32'h4466491f, 32'h442c53e2},
  {32'h43cbb591, 32'h444d6194, 32'hc3b2a0f9},
  {32'h441db44f, 32'h43bd31b8, 32'h442c4203},
  {32'hc4b13fa4, 32'hc41a8598, 32'hc33555d7},
  {32'h430ea71e, 32'h42baf715, 32'hc4e8c396},
  {32'hc38f30dd, 32'hc3ef2eee, 32'h444ead86},
  {32'hc342694c, 32'h447d2bdc, 32'hc4a72d41},
  {32'h43a4a104, 32'hc310de70, 32'h43874365},
  {32'h44b240c4, 32'h44056ed1, 32'hc462d074},
  {32'hc3298460, 32'h42aca878, 32'h449faaf0},
  {32'h43f213c8, 32'h42928719, 32'hc48d9f8b},
  {32'hc56d8466, 32'hc22e86ac, 32'h416c1e95},
  {32'hc4542ba3, 32'hc3c7ed0b, 32'h43ee41e5},
  {32'hc2a90bd0, 32'h450927c2, 32'hc40abcdf},
  {32'h42fa5c83, 32'hc4c46ae7, 32'h445a5de3},
  {32'h438f4f6e, 32'hc3f5a780, 32'hc50724f2},
  {32'hc53b8ade, 32'h43c3a8ea, 32'hc37877c9},
  {32'h4321d40f, 32'h42dabe10, 32'hc2d81d09},
  {32'h43f519c6, 32'hc4d3e32e, 32'hc4275f5c},
  {32'hc38acaff, 32'h44a15d69, 32'h44596191},
  {32'h43fdb5bc, 32'h417f5786, 32'h443237b0},
  {32'hc3cdb4f0, 32'h43f9165e, 32'hc3e2a508},
  {32'h4381271e, 32'hc55189bf, 32'h433fa84b},
  {32'hc4c0b3ad, 32'h43b0ebae, 32'hc3977954},
  {32'h455575b8, 32'hc29440df, 32'hc40b06ca},
  {32'hc4b96971, 32'h4492662e, 32'h4485bcb7},
  {32'h45580ecf, 32'h4065c70a, 32'h44265c4a},
  {32'h444067ce, 32'h44f959bc, 32'h425e6d07},
  {32'h442ec9f1, 32'hc40e9ad2, 32'h44b58776},
  {32'hc3524680, 32'h439f8d06, 32'hc44edd25},
  {32'h440cb39c, 32'hc3486fea, 32'h4448cdba},
  {32'hc42616f3, 32'h42a7b8f6, 32'hc54824a9},
  {32'hc490ff10, 32'hc340fbad, 32'hc389e057},
  {32'hc4795b84, 32'h4421c7b3, 32'hc2c7b2ce},
  {32'h44464078, 32'h4332cdec, 32'h4488b4b2},
  {32'h441a2c5d, 32'hc30db002, 32'hc4bc4bf7},
  {32'h43a22c88, 32'hc52d244a, 32'h43896ee4},
  {32'hc2c6db54, 32'h44e59f5a, 32'hc4348bf1},
  {32'h43aa06cc, 32'hc41d1bc0, 32'h436b3210},
  {32'hc3999a64, 32'h45037ce0, 32'h420ddb36},
  {32'h43e19a52, 32'hc398d933, 32'h45051f8d},
  {32'hc0cb7acc, 32'h440fe4c0, 32'h42a5af8a},
  {32'h44157652, 32'hc370ea2b, 32'h43ffe8c8},
  {32'hc500fb8e, 32'h439c30c0, 32'hc422be6a},
  {32'hc409bf98, 32'h416cc004, 32'h445f527d},
  {32'hc469f05c, 32'hc3619fe5, 32'hc451e5fd},
  {32'hc2d9987e, 32'h4450bf20, 32'h45235bc0},
  {32'hc39a3ca7, 32'h43e9bdba, 32'hc3756756},
  {32'h4499fff6, 32'h44007351, 32'hc40f5bb8},
  {32'h43545394, 32'hc4b22372, 32'h44808284},
  {32'hc52729c4, 32'h43ed6a16, 32'h420e52cc},
  {32'h40ce5210, 32'hc4499f51, 32'h4413d2d6},
  {32'hc5328c53, 32'h438680cf, 32'hc38c84c8},
  {32'h443611ba, 32'hc4949519, 32'h44b97439},
  {32'h44056ab8, 32'hc48eb734, 32'h44f2462b},
  {32'hc47fa52e, 32'hc4455bac, 32'hc475efbc},
  {32'h443937cf, 32'hc4004817, 32'h43992468},
  {32'hc2ff9efd, 32'hc2b2b040, 32'h449038dd},
  {32'h42233fc0, 32'h444e90dd, 32'hc49b74fe},
  {32'h429f3270, 32'hc51e7a9e, 32'hc326c42c},
  {32'h4435285e, 32'h447f762c, 32'h430f7e90},
  {32'hc1ba3ad8, 32'hc54b3687, 32'hc3aab84f},
  {32'h43ac23e0, 32'h4439315d, 32'hc4654190},
  {32'h4432eb3c, 32'hc4210291, 32'h43288263},
  {32'hc5725d7b, 32'hc3b9fb7a, 32'hc282403a},
  {32'hc39c59b0, 32'h441b3f43, 32'h43b79d09},
  {32'h44cfcaa3, 32'h44347987, 32'hc2d2a1b6},
  {32'h450d5905, 32'hc420d3e2, 32'h442b445a},
  {32'hc4a41bfa, 32'h44771ae6, 32'h43b3c2e4},
  {32'hc3c97e90, 32'hc451eba0, 32'hc3344514},
  {32'hc4a9780e, 32'h44bb150c, 32'h42a4d16e},
  {32'hc38a5b1e, 32'hc5663a22, 32'hc29d4935},
  {32'hc4317286, 32'h41d1ec45, 32'h43d501d2},
  {32'hc302f67c, 32'h44849f58, 32'hc50dba3c},
  {32'hc518ef32, 32'h4316961d, 32'h43e07e81},
  {32'hc39e4496, 32'hc45c98be, 32'h4439be29},
  {32'h4535e2f5, 32'hc1eb1616, 32'hc241e70f},
  {32'hc4db0950, 32'hc3a67424, 32'hc3535122},
  {32'h451a9e2a, 32'h44439c9a, 32'h41b9cd69},
  {32'hc3089f78, 32'hc22fefaf, 32'h44e6fca8},
  {32'hc48fd560, 32'h44341c84, 32'hc2207f97},
  {32'h4449ba0e, 32'hc3ba3074, 32'hc3d63d1f},
  {32'hc44060e5, 32'hc4d0d636, 32'h442a890f},
  {32'h43c098c8, 32'h42fdc34d, 32'hc4e0f9de},
  {32'h4356894d, 32'h44fef47a, 32'h42bfd804},
  {32'hc405b446, 32'h4249337e, 32'h449a7970},
  {32'h438d7378, 32'h423644bb, 32'hc444af7b},
  {32'hbf96a580, 32'hc394c737, 32'h4431099e},
  {32'h455832cc, 32'h42101e16, 32'hc302f4d0},
  {32'h44b9d0f1, 32'hc31ee5a4, 32'h43ddbfa1},
  {32'hc36115f9, 32'hc4274ac1, 32'hc3a35c35},
  {32'hc5440a20, 32'hc1ecb289, 32'h42875086},
  {32'h437dabe2, 32'h43bb25a1, 32'h418fd3fb},
  {32'hc35ae855, 32'hc54a7cea, 32'hc2a1e4f9},
  {32'hc40ac730, 32'h44f966ce, 32'h43668e82},
  {32'hc36b1250, 32'h438cba8c, 32'hc347ce88},
  {32'h4506ef27, 32'h443ef7ca, 32'h433bf228},
  {32'h439f5f04, 32'hc540f021, 32'hc38070bb},
  {32'hc2187bc2, 32'h443b33c3, 32'h43197dc8},
  {32'h43dfa7da, 32'h43b412bc, 32'h448d7a0a},
  {32'h427ff598, 32'hc495828e, 32'hc40f0874},
  {32'hc3835fda, 32'hc45e0bd6, 32'h44a6368b},
  {32'hc32a55f0, 32'hc31e6396, 32'hc4d6466f},
  {32'h44cadb78, 32'h42fb1b59, 32'h43b2a975},
  {32'h43879f67, 32'hc25a34d3, 32'hc3decb57},
  {32'h453324ce, 32'h434eb6fe, 32'hbec9f500},
  {32'hc34aa134, 32'hc3196dfa, 32'hc51d33de},
  {32'h42d064eb, 32'h441748e6, 32'h453f9b57},
  {32'h4460e6c9, 32'h4452e5d4, 32'h43654bf8},
  {32'h42fa8218, 32'hc41019fd, 32'h44ae0627},
  {32'hc47c0212, 32'h4442d30a, 32'hc461d7f1},
  {32'h43aa88ac, 32'h44f4f4be, 32'h42f8c8aa},
  {32'hc4411ff7, 32'hc3c950f3, 32'hc49eef48},
  {32'h444b6d6f, 32'h450c1554, 32'hc2b8d6d6},
  {32'hc48b114d, 32'h43c6d217, 32'h431192d6},
  {32'h44cef1e5, 32'h438c607b, 32'h445c27af},
  {32'hc53586f9, 32'h4355f44a, 32'h417f8fda},
  {32'h4523b414, 32'hc30bb272, 32'h44a66e68},
  {32'hc4cbdd1b, 32'hc4ab4cbc, 32'hc4141708},
  {32'hc391f8ae, 32'h456ef1a0, 32'hc1b907b4},
  {32'hbea7b100, 32'hc3ba34ac, 32'hc3ebd9c5},
  {32'h44731d1e, 32'h44ec3829, 32'hc29950e9},
  {32'hc33e670a, 32'hc519eb76, 32'hc183281e},
  {32'h44cca32f, 32'h42de92c3, 32'h4356f66c},
  {32'hc58ff56a, 32'h408ab201, 32'hc3824e16},
  {32'h44625360, 32'hc435cc8d, 32'h441e979f},
  {32'h43a85298, 32'hc3ccdd44, 32'hc4820e51},
  {32'h42806639, 32'h42b0f830, 32'h44565a85},
  {32'h44b12ee0, 32'h44203b57, 32'h43da2c59},
  {32'hc45a943a, 32'h44c5f34a, 32'h439d4c39},
  {32'h4383b24e, 32'hc4ffb3c5, 32'hc4497cf2},
  {32'hc3cbb72a, 32'hc2000067, 32'h44bae447},
  {32'h42da2820, 32'hc497d544, 32'hc49b2adc},
  {32'hc457c13c, 32'h441a0b56, 32'h44e1343c},
  {32'hc397ec77, 32'hc48a8e77, 32'hc39157ee},
  {32'h42a40364, 32'hc4111191, 32'h44a8e262},
  {32'h4512067e, 32'h440e5448, 32'h43dc54fc},
  {32'hc498c98f, 32'hc42fcfb9, 32'hc28ef0c4},
  {32'h42d33990, 32'hc514e7f1, 32'hc42e9677},
  {32'hc40d6ec8, 32'h4509b964, 32'hc1caf41d},
  {32'hc4d6e73d, 32'hc2b390ee, 32'hc2f22b99},
  {32'hc4a42c46, 32'h4410b1ab, 32'h441a89b9},
  {32'hc3bc7c1f, 32'h438cf47e, 32'hc4a162a6},
  {32'h450127d1, 32'hc3c47457, 32'h4389a503},
  {32'h43d93e7a, 32'hc4e2591b, 32'hc363d93c},
  {32'hc44ec386, 32'h44617d92, 32'h44139b86},
  {32'h449807ba, 32'hc16c664e, 32'hc1a1c9d6},
  {32'h4309d816, 32'h45561030, 32'h41907e7c},
  {32'h42e2d294, 32'hc570e794, 32'hc39b0506},
  {32'h450e5b74, 32'hc2f175d1, 32'hc38bfd5e},
  {32'h44a66f20, 32'h420790b3, 32'h4374196a},
  {32'hc55e676c, 32'h40dfe6f0, 32'h42a2bac5},
  {32'h44d67c7b, 32'hc36eb924, 32'hc39d09aa},
  {32'h44dd13d6, 32'hc388b4cc, 32'hc41caa84},
  {32'hc51280d6, 32'h42c01278, 32'hc2c83cb4},
  {32'h4531422b, 32'h43a51452, 32'h44303d34},
  {32'h44af2f3f, 32'h439044e4, 32'hc2f9d23d},
  {32'h443d8c16, 32'hc537b574, 32'h430ab8a4},
  {32'hc489b8a6, 32'h44b91cdc, 32'hc318858d},
  {32'h441346ba, 32'hc4aea8cb, 32'h4363fcbf},
  {32'hc429b2f8, 32'h44b60288, 32'h435d07fe},
  {32'h4459626c, 32'hc49a3293, 32'hc34fd074},
  {32'h44f56676, 32'hc1c922a2, 32'hc1e1cdf6},
  {32'h44710d95, 32'hc40b38a1, 32'h4306ea04},
  {32'hc4234fea, 32'h4499b070, 32'h4480e1d5},
  {32'h440fc296, 32'hc4378775, 32'hc42dc276},
  {32'hc43607ea, 32'h44be2199, 32'h43e4aa39},
  {32'h43764e8c, 32'hc4a44fcd, 32'hc468174a},
  {32'h4410588c, 32'h43e580b9, 32'h42a894e8},
  {32'h444d9b42, 32'hc491b4e7, 32'hc2fdc968},
  {32'hc298b3aa, 32'h426752f8, 32'h454c4714},
  {32'h45276ae5, 32'hc394241c, 32'hc1ed2dd7},
  {32'hc593b873, 32'h4308ed4b, 32'hc36e68cc},
  {32'h453f91a3, 32'h437df5e2, 32'hc43848e2},
  {32'hc4db22b4, 32'h440145b6, 32'hc3bd70bb},
  {32'hc36dbc74, 32'hc31fcd6e, 32'hc5470a52},
  {32'hc475a842, 32'h4478f3b2, 32'h44d94ed1},
  {32'h44b72046, 32'hc3c4cf97, 32'hc40459d6},
  {32'hc3e45ec6, 32'h430a5077, 32'h42d0700f},
  {32'h43734b10, 32'hc4e46a1e, 32'hc3ee1955},
  {32'h44b10d7b, 32'hc1c8797f, 32'hc4313d24},
  {32'hc4fc2cd0, 32'h4189764a, 32'h43d70425},
  {32'h44e8a54c, 32'h43d8c77d, 32'hc3312c8a},
  {32'hc502c5b1, 32'hc415a3fe, 32'hc2fae12c},
  {32'h4440a49f, 32'h4496a560, 32'hc35c95a5},
  {32'h4520ce87, 32'hc2470cb6, 32'hc36052fa},
  {32'h447fac36, 32'h453dda52, 32'h43ec39d4},
  {32'hc49eed98, 32'hc4f6eb37, 32'hc3839a8e},
  {32'h4434616b, 32'h43932273, 32'h41c289ce},
  {32'hc4bb477a, 32'hc4110986, 32'h432e5252},
  {32'h442820c0, 32'hc315f22a, 32'hc301f258},
  {32'h44ce1ede, 32'hc4136603, 32'h43fd0e31},
  {32'h43828e70, 32'h43533720, 32'h451490f2},
  {32'hc4814d4c, 32'hc43437e6, 32'hc4a7ce4e},
  {32'hc47be224, 32'h428dfd9c, 32'h4413f05e},
  {32'hc51351ae, 32'hc3a21f09, 32'hc425d1de},
  {32'h44201290, 32'h441e161e, 32'hc3c75062},
  {32'hc4ad9c99, 32'hc422393b, 32'hc4620fcf},
  {32'h451ce6b6, 32'h440cd639, 32'h442317d8},
  {32'hc38ab12c, 32'h4475fb8c, 32'hc49fdd4c},
  {32'h44f67fda, 32'h43a9f426, 32'hc3a29b45},
  {32'hc3b00c58, 32'hc476b936, 32'hc421016e},
  {32'h44f7e4e9, 32'h4389de3b, 32'hc20294c8},
  {32'hc3356446, 32'hc3d2348c, 32'hc3846210},
  {32'h43375050, 32'h449425c4, 32'h4515befc},
  {32'hc5214e8c, 32'hc387c9eb, 32'hc1de9ba0},
  {32'hc2a50c66, 32'hc241c0dc, 32'h43d5167b},
  {32'hc49c758c, 32'h435f6099, 32'hc31420f6},
  {32'hc51e5910, 32'h43c21337, 32'h43c312d5},
  {32'h4195c788, 32'h45102e32, 32'h44449165},
  {32'h45045535, 32'hc3d7cca9, 32'h432694db},
  {32'h42a96e00, 32'h446fa050, 32'h443f1c5a},
  {32'hc510960b, 32'hc4500327, 32'hc37f74e2},
  {32'h4487a87b, 32'h43940da5, 32'hc3316649},
  {32'hc532d7d2, 32'h430fc5fa, 32'hc39d15a1},
  {32'h44fd3243, 32'h438e8504, 32'h4466f6f7},
  {32'h44b9c595, 32'h43cdfe1d, 32'hc39b28cc},
  {32'h43267a3d, 32'h45097f89, 32'h42288182},
  {32'hc4305958, 32'hc40ea6f6, 32'h44061111},
  {32'h421ce6c0, 32'h4485e537, 32'hc4279d28},
  {32'hc3fd882c, 32'hc482ae67, 32'h44621544},
  {32'h4406c7bc, 32'h45231c87, 32'hc422f176},
  {32'hc3e40204, 32'h41e0eb73, 32'hc3dc3685},
  {32'h44407403, 32'h431c3fc1, 32'hc475767f},
  {32'hc49a4d71, 32'hc4749811, 32'hc3cd7f58},
  {32'h45109dfd, 32'h42899957, 32'hc3846f72},
  {32'hc4e27814, 32'hc48a4f45, 32'h438714e3},
  {32'hc4853e8a, 32'h44207630, 32'hc1a3df7c},
  {32'h45503599, 32'h44249b1c, 32'hc3ce5320},
  {32'hc4fde517, 32'h43163b74, 32'h440a3cca},
  {32'hc3e0b446, 32'hc2e0dca6, 32'hc4bf7122},
  {32'hc3c77f08, 32'h428aa4b4, 32'h44ce99dc},
  {32'h44464eb6, 32'hc43744d0, 32'hc534f09d},
  {32'hc2a836e8, 32'hc5235be3, 32'hc3977780},
  {32'hc49987b8, 32'h44a6134f, 32'hc23932a7},
  {32'hc4c55e89, 32'hc38f81bf, 32'h42f17152},
  {32'h41d3b680, 32'h451e43bc, 32'hc3bb7dc9},
  {32'h4359ade4, 32'hc50ef13a, 32'hc3401eeb},
  {32'hc4a5abc8, 32'h4360b534, 32'hc2f82bca},
  {32'h43eae6f0, 32'h43186aae, 32'hc2abdc1c},
  {32'hc54efa68, 32'hc335a805, 32'hc38e89a9},
  {32'h43f54b20, 32'hc285d088, 32'h441ccd75},
  {32'hc3a6a952, 32'h450403e0, 32'hc31c44d8},
  {32'h44a407b2, 32'h40b82dc2, 32'h439ae438},
  {32'hc4c831d3, 32'h400c4b67, 32'hc32784ce},
  {32'h427a611c, 32'hc5169530, 32'h43332b93},
  {32'hc3d3d2a9, 32'h43f31815, 32'hc4905722},
  {32'h451931b1, 32'h438f395e, 32'h43adce82},
  {32'hc4d09ef6, 32'h443afd04, 32'h440f9413},
  {32'h452d759f, 32'hc3370262, 32'h42fc0163},
  {32'hc41b8614, 32'h423e035a, 32'hc3c20171},
  {32'h451aea4a, 32'hc38712ad, 32'h43896e44},
  {32'hc500bdb4, 32'h44bd1e57, 32'hc4770232},
  {32'h44197ef1, 32'hc40607ed, 32'h44861c51},
  {32'hc36afe98, 32'h44e5a358, 32'hc39db9f9},
  {32'h4401492a, 32'hc495c0f6, 32'h44351c86},
  {32'h438bfdff, 32'h44824833, 32'hc3b2230b},
  {32'h44ee9734, 32'h43a1636a, 32'h4450b412},
  {32'hc541919b, 32'hc3953b3a, 32'hc3f72f8c},
  {32'h4424c26f, 32'h4355dcad, 32'h44a88662},
  {32'hc4dd42b6, 32'h41deb3a3, 32'hc3d810d9},
  {32'h45190506, 32'h441a5a20, 32'h4385179a},
  {32'h4391c16d, 32'h444df649, 32'hc410bef3},
  {32'h444fc59f, 32'h4407f8fb, 32'hc3d6f901},
  {32'hc39e7a5c, 32'hc487d4af, 32'h442fe64f},
  {32'h431c3958, 32'h44733039, 32'hc41cc192},
  {32'h4471243d, 32'hc41a4d58, 32'hc202e315},
  {32'hc4647415, 32'h4482c0db, 32'hc44191af},
  {32'h4428a48c, 32'hc3b73ef7, 32'h44d8fdc2},
  {32'h4510e141, 32'h4471d059, 32'h4484498e},
  {32'hc4e43010, 32'h441bddd0, 32'h43ef308d},
  {32'hc3e17c39, 32'h4420ad23, 32'h43eea107},
  {32'hc4100dc8, 32'hc49a71a6, 32'hc39db5ba},
  {32'hc3ff5650, 32'h44051897, 32'hc3504f5c},
  {32'h44322f90, 32'hc3cdc380, 32'h42cf71a4},
  {32'hc3b876e0, 32'h42a27e94, 32'hc4941f8b},
  {32'h4424137d, 32'h44010121, 32'h44fdf069},
  {32'hc4b7d077, 32'h440f0f63, 32'hc3f731e0},
  {32'h44ea5eed, 32'hc42818db, 32'h435e6b67},
  {32'hc56d7753, 32'hc3e3c1a6, 32'hc3429f0a},
  {32'hc3828120, 32'h433f40df, 32'h44897ead},
  {32'h43644ad4, 32'h447c77e5, 32'hc3ce0b08},
  {32'h448b5c85, 32'hc4bd2004, 32'h43930b5d},
  {32'hc261b300, 32'h43fdacce, 32'h42477df5},
  {32'h44a542ae, 32'h44031053, 32'h43988fb4},
  {32'hc4983858, 32'h44ef435f, 32'hc2b3cdf4},
  {32'h43e956a5, 32'hc4d1d14d, 32'h42a5dba5},
  {32'h44385755, 32'h44b61890, 32'h44a72a12},
  {32'h44995738, 32'hc2c2f237, 32'hc461062c},
  {32'hc4b29329, 32'h44015629, 32'h43a83f4b},
  {32'hc4c13d43, 32'hc3fc5df0, 32'h440acf24},
  {32'h452d2b1e, 32'hc373d767, 32'h43805c42},
  {32'hc3eb2b35, 32'h42a0fd34, 32'h44db1d9f},
  {32'h454078c6, 32'h437075fc, 32'hc3a5ec69},
  {32'hc3f201f8, 32'hc4832f5b, 32'h443b97a2},
  {32'h4435b9ad, 32'h43dad199, 32'h436bbcb4},
  {32'hc4c35b65, 32'hc31d2305, 32'h43b5910a},
  {32'hc3ca9da8, 32'hc4a77e14, 32'h44da139a},
  {32'h424ff43e, 32'hc4bb038e, 32'hc4a5c015},
  {32'h4361f420, 32'h44ba5d98, 32'hc36cf38c},
  {32'hc46d64f5, 32'hc439710e, 32'h446a2ae5},
  {32'h43236f38, 32'h4494023b, 32'hc49a9be2},
  {32'hc4885141, 32'hc49723b5, 32'h442da233},
  {32'h44aed051, 32'h4464d461, 32'hc381a930},
  {32'h43476f53, 32'hc380ce95, 32'h44988803},
  {32'h440dd3c6, 32'hc4349398, 32'h43c1a93b},
  {32'hc5233946, 32'h4317711f, 32'h4455a139},
  {32'h455e4f52, 32'h43923d8a, 32'hc3cb13c6},
  {32'h431fdff5, 32'hc5814441, 32'h41d7b323},
  {32'h44b6be44, 32'h445f43bf, 32'hc35cd1cb},
  {32'hc2b647d5, 32'hc4c6b1f1, 32'h44123ca3},
  {32'h40209c5e, 32'h4525ef29, 32'hc3e7f82f},
  {32'hc49bb65a, 32'hc493dffe, 32'h4301841e},
  {32'h443a4ef8, 32'h4485ace0, 32'h42f0282e},
  {32'hc2771b50, 32'hc33ed6de, 32'h43a03f16},
  {32'h43553a0b, 32'h438f65e3, 32'h4219be37},
  {32'h4405313f, 32'h452a8f15, 32'h43d58149},
  {32'h435311aa, 32'hc4699363, 32'hc3aed2b0},
  {32'hc3e5fbcd, 32'h443d25d7, 32'h44ac3ed2},
  {32'hc2e9ec00, 32'hc4ddb1f5, 32'hc48b5516},
  {32'h44ea5478, 32'hc3797e90, 32'hc3a4c443},
  {32'hc40c709c, 32'hc4b38f8e, 32'hc4e8f30e},
  {32'h43cdbba3, 32'h43c04253, 32'h451517b1},
  {32'h441af35c, 32'h44d798c6, 32'hc4303292},
  {32'hc3b0df04, 32'h45133893, 32'hc4045df6},
  {32'h43263e17, 32'h44afd82a, 32'hc51cb10f},
  {32'h441b8c3e, 32'h446aa966, 32'hc164dc15},
  {32'hc40588e7, 32'hc367f92e, 32'hc492a013},
  {32'h44002c58, 32'h44957224, 32'h44982fc2},
  {32'h43e79924, 32'hc488d95d, 32'hc33df4d3},
  {32'h442b277c, 32'h43cddd3c, 32'h44332fff},
  {32'hc52cda5d, 32'hc37cd2f6, 32'h436ab057},
  {32'hc2f49efa, 32'h44c2d035, 32'hc3500780},
  {32'hc4ee15d5, 32'hc4711063, 32'hc3abcacd},
  {32'h44d62ec2, 32'h4499ea57, 32'h445563c5},
  {32'h44ab171a, 32'hc3d482e0, 32'hc385802e},
  {32'h44c879cb, 32'h4491c11e, 32'h441481aa},
  {32'hc4ed8578, 32'hc3f98944, 32'hc3086772},
  {32'hc4953aa9, 32'hc260d848, 32'hc4107896},
  {32'hc58db021, 32'hc249c703, 32'hc2a93afa},
  {32'hc3086b00, 32'hc415aa72, 32'hc385bfc7},
  {32'h44351e9b, 32'h449cb1cc, 32'hc4b6da4c},
  {32'hc4593b54, 32'h4409386e, 32'h438bc4dc},
  {32'hc41198b0, 32'hc49dff02, 32'hc3860cb8},
  {32'hc453ef92, 32'h4520a7f1, 32'h43444551},
  {32'hc38b30c0, 32'hc2e999d1, 32'hc55f46e4},
  {32'h44a971e1, 32'h430c694a, 32'h43d07ee0},
  {32'h44dd0175, 32'hc4bbde8c, 32'hc48b1de4},
  {32'hc46c95b4, 32'h43299178, 32'h44c1504b},
  {32'hc3ca0d8c, 32'hc4586d3d, 32'hc3eadd87},
  {32'h439a2221, 32'hc27d0f2c, 32'h44cc4eb4},
  {32'h44bf4e00, 32'h43f4d743, 32'hc3e67750},
  {32'h436e9246, 32'h437c00fe, 32'h438e45bf},
  {32'h44ae8420, 32'h431894af, 32'hc3f6c252},
  {32'hc49bd042, 32'h43848309, 32'h43ad7066},
  {32'hc3121c08, 32'hc436aa7c, 32'hc42b0bf9},
  {32'h44732c4e, 32'h447726a0, 32'h45349dd7},
  {32'h43e61c8a, 32'hc50b9971, 32'hc4afd4ec},
  {32'hc45fd074, 32'h441aad9f, 32'h433f81ce},
  {32'h4522702d, 32'hc49f99c0, 32'hc34019a3},
  {32'hc4e10dfc, 32'h4441bcfc, 32'hc33b7028},
  {32'hc497bea1, 32'hc289f2d8, 32'h4079e03a},
  {32'h43b49a88, 32'h44134062, 32'h4376018b},
  {32'h45427706, 32'hc38802b1, 32'h439d6c75},
  {32'hc37b31b2, 32'hc387ab7e, 32'hc3024efe},
  {32'h449fc6a6, 32'h43e6dd49, 32'hc22c9baa},
  {32'hc59253d8, 32'hc32133cc, 32'hc2b5b3b5},
  {32'hc33d401a, 32'hc39039f4, 32'hc3d924b1},
  {32'h44785a1f, 32'h416c0dda, 32'h4467f4eb},
  {32'hc531f6bf, 32'hc3909130, 32'hc384df1a},
  {32'h43ac5af8, 32'h427589ad, 32'h4345c959},
  {32'hc4a7895e, 32'h44121eba, 32'h42a40e92},
  {32'h452beeef, 32'hc3f69de5, 32'hc351cbbf},
  {32'hc3fa266a, 32'hc34b6437, 32'h4338617e},
  {32'h44980909, 32'hc3272483, 32'hc28ac000},
  {32'hc4138f94, 32'h453b5073, 32'hc3701e6d},
  {32'h45296538, 32'hc3f4a8c8, 32'h42a054b4},
  {32'hc4f7c7ef, 32'hc38d7907, 32'hc40a396c},
  {32'h454494e3, 32'hc2c6085d, 32'h43a38b5b},
  {32'hc328abb3, 32'h4393d49c, 32'hc4544019},
  {32'h44abe424, 32'hc3bd71b2, 32'h43744500},
  {32'h41843164, 32'h452d31de, 32'h43492816},
  {32'h44e26a5c, 32'hc24b415f, 32'hc3d5cc62},
  {32'hc4682cf6, 32'h44532c13, 32'h42bfa3c1},
  {32'hc4131986, 32'hc40535f7, 32'hc50abab9},
  {32'h441aa354, 32'h4363ca08, 32'h4419784a},
  {32'hc4fa3f53, 32'h432b5bea, 32'hc3034c0d},
  {32'hc4557758, 32'hc38fc824, 32'h43cec45e},
  {32'h44ced5de, 32'hc2495859, 32'hc4885d19},
  {32'hc4913fd0, 32'hc2862604, 32'h43dac746},
  {32'h448ad077, 32'hc43ab872, 32'hc411e1ca},
  {32'hc412f9e9, 32'h44836649, 32'h449efbd9},
  {32'h4265f453, 32'hc2c54d9b, 32'hc484820e},
  {32'hc3c049c1, 32'h433aeff9, 32'h442f8302},
  {32'hc2eec7ed, 32'hc413ca62, 32'hc55e27bd},
  {32'h45513350, 32'h42a3838d, 32'hc3a6aa2a},
  {32'hc51400c3, 32'hc3783c5a, 32'h44c343db},
  {32'hc3bbb7f4, 32'h4442587e, 32'hc3fd95f8},
  {32'hc4302f6f, 32'hc43409cf, 32'h43f7bdf8},
  {32'h432400f7, 32'h450b4e76, 32'h438c3042},
  {32'hc42e604a, 32'hc47e19f3, 32'hc3db12c2},
  {32'h44d737f6, 32'h4456b9f6, 32'hc35794a8},
  {32'hc4bcc786, 32'hc4d9f1a1, 32'h438eb8d1},
  {32'h43d14313, 32'h43778057, 32'hc214dad1},
  {32'h41afbb88, 32'h43bb816f, 32'h44caa138},
  {32'h44e1f91e, 32'h4255d306, 32'h42ac40da},
  {32'hc4428df8, 32'h4255df3b, 32'h443566c1},
  {32'h42a7a916, 32'h4490d3d6, 32'h448acec2},
  {32'hc390a408, 32'hc34ba7b4, 32'hc4f6df02},
  {32'hc2b208b2, 32'h43f3316e, 32'h448606e6},
  {32'h42ad5d6c, 32'hc48dacb9, 32'hc452b305},
  {32'hc2ae92b7, 32'h4486d75b, 32'hc33cb4fc},
  {32'hc41a464d, 32'hc3acbcbc, 32'hc191ab38},
  {32'h44e92c43, 32'hc48c8f3e, 32'h44cd7daf},
  {32'hc43f90a4, 32'hc47952cc, 32'hc4e42b16},
  {32'h44c4ccdc, 32'hc41d50f8, 32'hc40caebc},
  {32'hc4870722, 32'hc1c15bcb, 32'hc44f707f},
  {32'h447e0105, 32'h431ff048, 32'h44b60587},
  {32'h43af67e3, 32'h4202b13b, 32'hc49d35bc},
  {32'h4241c5b0, 32'h44c69a5d, 32'h447f0b6a},
  {32'hc44eef38, 32'hc50e92b7, 32'h400d9d53},
  {32'h434c9a0b, 32'h42cc3424, 32'h446b3c57},
  {32'h44f1a80a, 32'hc344d4dc, 32'hc3a03c48},
  {32'hc5111799, 32'hc38e2d61, 32'hc286bacb},
  {32'h4462e000, 32'h443149aa, 32'h4425065c},
  {32'h40e1587e, 32'hc45196be, 32'h437e5707},
  {32'h4448f524, 32'h44bea6a3, 32'hc3c06823},
  {32'hc433603b, 32'hc51c1e54, 32'h438b9c67},
  {32'hc3a42458, 32'h42fa080f, 32'hc3cfdce0},
  {32'hc40d3f30, 32'hc3111ceb, 32'hc12e3d1a},
  {32'h45201adc, 32'h4410bd3e, 32'h44674ed7},
  {32'h4148bc68, 32'hc40ff801, 32'h4416ea42},
  {32'h44a6ec76, 32'h43be7106, 32'h43ed3ccd},
  {32'hc3972440, 32'hc386b294, 32'hc4203812},
  {32'h44d8e1e2, 32'h438e82db, 32'hc24938c8},
  {32'hc3c086b4, 32'hc510226d, 32'h43196963},
  {32'h44683273, 32'h4398337d, 32'hc4618530},
  {32'hc4b436f1, 32'hc3ccc5f4, 32'hc386c457},
  {32'hc313dc97, 32'hc28f5440, 32'hc555150e},
  {32'hc40e2c1a, 32'h43e31a72, 32'h45289e4f},
  {32'hc32a017e, 32'h44fa5726, 32'hc3c32667},
  {32'hc2949e78, 32'hc55de6a3, 32'h43303c0c},
  {32'h441138eb, 32'hc504e28a, 32'h438c2c8a},
  {32'hc2534ec0, 32'h44a5ff31, 32'hc47e9213},
  {32'hc425d7ec, 32'hc399a11a, 32'h44420550},
  {32'h4499dc3c, 32'h43886de5, 32'hc4d34b08},
  {32'hc4987c64, 32'h43a8787b, 32'h4486fa43},
  {32'h43976ca0, 32'hc2d1ec4e, 32'hc4c78067},
  {32'h44c40b08, 32'hc46b858c, 32'h42a24a6f},
  {32'hc4234677, 32'h452e2a9c, 32'h435f2697},
  {32'h444ab30d, 32'h4360a5df, 32'h43b68bde},
  {32'hc1b01d76, 32'h4547cb35, 32'h4328be98},
  {32'h451fa1db, 32'hc3be1640, 32'hc3a9427f},
  {32'h439e420e, 32'h43bd0446, 32'hc323ea26},
  {32'h45160a1b, 32'h43d60f81, 32'h4315530a},
  {32'hc57c315c, 32'h4343b405, 32'h43fa7eb2},
  {32'h45142efb, 32'hc44b79f2, 32'h43c8972e},
  {32'h43659350, 32'h44952249, 32'hc4648bd8},
  {32'hc389aa72, 32'hc4ea62a8, 32'hc2bbbef6},
  {32'hc328acb7, 32'h44b4675c, 32'h42c12146},
  {32'h439ee02c, 32'hc18b1408, 32'h44fe9e70},
  {32'hc45de0de, 32'h4463acc1, 32'h4254b3cc},
  {32'h4402f813, 32'hc413df6d, 32'h440b4eef},
  {32'hc4355f09, 32'hc309398d, 32'hc4d1028f},
  {32'h45020efe, 32'hc43df88b, 32'h43054554},
  {32'hc525aa50, 32'h420ec886, 32'hc31e5596},
  {32'h450a7f82, 32'hc4720afb, 32'hc329eb7f},
  {32'hc4bd53a6, 32'h44d9e20f, 32'hc4176ae3},
  {32'h4537a911, 32'h439d34b9, 32'hc34ba28f},
  {32'hc2a418a0, 32'h449d465a, 32'hc41359d5},
  {32'h44834d20, 32'hc4f0d51c, 32'hc3ec7953},
  {32'h44ba3257, 32'h44017c2c, 32'hc35551d0},
  {32'h44ad6074, 32'h44027ead, 32'h44e2ac10},
  {32'hc574204c, 32'h43595def, 32'hc46e4992},
  {32'h44c94f9a, 32'h4280a42a, 32'h42b75b1d},
  {32'h427dd0cc, 32'h448dc923, 32'hc4c1836b},
  {32'h4474498b, 32'h43e30649, 32'h4494b1b7},
  {32'hc513e330, 32'h43a1c6a9, 32'h43b22b57},
  {32'h42ee44d0, 32'h438aa5c0, 32'hc4874002},
  {32'h4389545e, 32'hc3584f35, 32'h45326ebe},
  {32'hc42b357a, 32'h436e230e, 32'hc3b3677d},
  {32'hc0b64187, 32'hc34b5f2d, 32'h43c8b6f5},
  {32'hc47c2e8c, 32'h442a0063, 32'hc42d9b5a},
  {32'h44500d8e, 32'hc21798e6, 32'h44a47810},
  {32'h42e2da58, 32'h450d6dc7, 32'h44b3aa08},
  {32'hc1ca6050, 32'hc4590b64, 32'hc50a542b},
  {32'h4368f50e, 32'hc38cb11a, 32'h43d223f4},
  {32'h43f779ee, 32'hc400ebfc, 32'h44168b98},
  {32'hc4906a70, 32'h434e4f15, 32'hc46276f7},
  {32'h442b3a9c, 32'hc43262ac, 32'hc4112c16},
  {32'h44dc82d2, 32'h42d007e1, 32'h42f863c8},
  {32'h44ee2140, 32'h43384d73, 32'h443cd4fe},
  {32'h431d3442, 32'h45487302, 32'hc3d3def9},
  {32'h4512aa04, 32'hc416a7c1, 32'h42ac8954},
  {32'hc55571f4, 32'hc382aa71, 32'hc401e0c4},
  {32'hc3acf40a, 32'h43dc6b21, 32'h445c2f3a},
  {32'hc4b982f4, 32'h4296b9aa, 32'h433b17ef},
  {32'hc352edc2, 32'hc5793ba6, 32'hc3254b03},
  {32'hc53b5d80, 32'h42eee66d, 32'h434c5d2a},
  {32'h438bff1c, 32'hc518347a, 32'h42ab2c44},
  {32'hc3b58742, 32'h455e0fb7, 32'hc2a43e9e},
  {32'h44bee0f5, 32'hc4b3fce4, 32'h43a99a1d},
  {32'h451b78b6, 32'hc3a3b6cf, 32'h43949590},
  {32'hc3910ca9, 32'h449bd073, 32'hc4c5dd1b},
  {32'hc43b4af7, 32'h44462376, 32'h448899b8},
  {32'hc3fb6a12, 32'hc47bf57b, 32'h43911101},
  {32'hc2704358, 32'h44deec9c, 32'h43b2be6f},
  {32'hc48dd36c, 32'hc449dcd7, 32'h438a9913},
  {32'hc4106004, 32'h45322999, 32'hc147dcc2},
  {32'hc4ca4cf4, 32'hc46332d4, 32'h433e490a},
  {32'h42ec8de3, 32'h4495ee67, 32'hc183c786},
  {32'h43f2d13b, 32'hc42e9934, 32'hc290a415},
  {32'hc4e26072, 32'h429e7361, 32'hc316696a},
  {32'h4475fa35, 32'hc492fb8e, 32'hc4772d1a},
  {32'h44373b0d, 32'h44042ef5, 32'hc484c940},
  {32'hc3c2ddb5, 32'hc3a32acf, 32'h45448a45},
  {32'h44685104, 32'hc1d33ab0, 32'hc3a66d5e},
  {32'hc4479a34, 32'h432e8cf6, 32'h44ae8bcf},
  {32'hc3b84223, 32'h4500b0fe, 32'hc2a27e6c},
  {32'hc4b13ab0, 32'hc43b5ce4, 32'h441f9319},
  {32'h4526e9c0, 32'hc21df482, 32'hc319a10c},
  {32'hc45ce960, 32'hc213fea0, 32'h441e59f5},
  {32'hc466c01d, 32'h431371c9, 32'hc3217e18},
  {32'hc360ac7c, 32'hc5875023, 32'h430eff6d},
  {32'h44ffd494, 32'hc3c9e7d0, 32'h4294f00e},
  {32'h43446240, 32'hc4b7421a, 32'h4336098a},
  {32'hc2018da0, 32'h454dcbed, 32'h4319a4b2},
  {32'hc44c0ca8, 32'hc4ee79e4, 32'h43984e57},
  {32'h44a959ea, 32'hc398b7e6, 32'hc2f05e75},
  {32'hc2af28ed, 32'h44732281, 32'h4400af2f},
  {32'h43b33c6e, 32'hc489dce1, 32'hc3433c11},
  {32'hbff51000, 32'hc4ecc908, 32'h44db1817},
  {32'hc1acb03a, 32'h41c296da, 32'hc10144b3},
  {32'h439e3f51, 32'h4400b6a6, 32'h44edf662},
  {32'hc4ba326c, 32'hc45cb61e, 32'hc3852c2e},
  {32'hc4822050, 32'hc35c78aa, 32'h40c9ab70},
  {32'hc3c64427, 32'hc474c2dc, 32'hc4f06862},
  {32'h44e034b6, 32'hc34fd566, 32'h447f114b},
  {32'h44be0a7f, 32'h43b30a78, 32'hc35c636e},
  {32'h44f96b3a, 32'h43cb0b5c, 32'h43563e2d},
  {32'hc4e052c8, 32'hc37390c1, 32'hc3c00981},
  {32'h447a07ab, 32'h433e71fc, 32'h434bc159},
  {32'hc3ede849, 32'hc46588f6, 32'hc3ba9404},
  {32'h449092dc, 32'h444abae8, 32'h43083194},
  {32'hc4308ffa, 32'hc32272ea, 32'hc37f89dc},
  {32'h44415d8b, 32'h44106643, 32'h44e0d10b},
  {32'hc50fd6d4, 32'hc3fdbf56, 32'hc37e5c23},
  {32'hc4bb0fc6, 32'h436549c5, 32'h43f59e94},
  {32'hc3cc9330, 32'hc4f3dc45, 32'hc41116f5},
  {32'h44be6fa2, 32'h44b5aa71, 32'h44397ab6},
  {32'hc42a659d, 32'hc2c17028, 32'hc354a0aa},
  {32'hc426b391, 32'h4580be5d, 32'h43023ebf},
  {32'hc3f807fe, 32'hc4ef5ec2, 32'h4362800f},
  {32'hc396b483, 32'h43c8da22, 32'h42a4011c},
  {32'hc4c6cee4, 32'h412d33f0, 32'h42bc6d65},
  {32'h44cb3ce2, 32'h415c2814, 32'h426e382e},
  {32'hc2d07e79, 32'hc433b5e5, 32'hc4a97c47},
  {32'h42c44467, 32'hc4430e29, 32'h44b835d3},
  {32'h44766ef6, 32'h4370ac34, 32'h43fc0f41},
  {32'hc397a08a, 32'h42baff06, 32'h44fc19f8},
  {32'h451db16f, 32'hc39b6f9a, 32'hc3348d71},
  {32'hc392baa0, 32'h44905aac, 32'h44365303},
  {32'h439a3cac, 32'hc49f65b4, 32'hc4af7803},
  {32'hc3d6187f, 32'h439bdb98, 32'h4514d8ee},
  {32'h43c8ec5a, 32'hc48921db, 32'hc3f7304b},
  {32'h438ce503, 32'hc4f752cf, 32'h4508ef5a},
  {32'h432b21d8, 32'hc3a6592e, 32'hc46d479e},
  {32'h42cfcdc0, 32'h4349bc53, 32'h427ba28e},
  {32'hc1a24e08, 32'hc49a3fd8, 32'hc46c1d2f},
  {32'hc4285534, 32'h43c75238, 32'h447048a2},
  {32'h44611342, 32'h4335f0c8, 32'hc4568e96},
  {32'hc323f8a4, 32'h4451c964, 32'h4503014f},
  {32'h44846980, 32'hc4d50cfa, 32'hc471f4c7},
  {32'hc2ea2d88, 32'hc3e0b132, 32'h44ba3137},
  {32'h430156d6, 32'hc5014c9c, 32'h42d494a1},
  {32'hc5096203, 32'h4411ad10, 32'hc42380bd},
  {32'hc32e3a2c, 32'hc472e5a3, 32'hc392cf43},
  {32'hc4395112, 32'h4553a172, 32'h4322978a},
  {32'h4452972e, 32'hc5581ad1, 32'hc411709a},
  {32'hc4928d4a, 32'h44596b73, 32'hc1a6b5d6},
  {32'h44d522fc, 32'hc39f6fbc, 32'hc3f3961d},
  {32'hc51352ef, 32'hc2b6b2cd, 32'hc3597a03},
  {32'h45788817, 32'h41c631bd, 32'hc40c7893},
  {32'h446ae989, 32'h41c91373, 32'h41da58b2},
  {32'hc546567c, 32'h43838525, 32'h4123847c},
  {32'hc3f3fdf8, 32'h4440f1b9, 32'h43a5a7fb},
  {32'h439712f9, 32'h4519e8c0, 32'h41d8295c},
  {32'h43261dad, 32'hc530f798, 32'hc39879f3},
  {32'hc39dbf14, 32'h452600cf, 32'h43a8269c},
  {32'hc4b4c9c2, 32'hc3d5b420, 32'h4371da0e},
  {32'hc4eae521, 32'h448df6e8, 32'h43a9079e},
  {32'h44aad8d2, 32'hc4d11e75, 32'h43a394e4},
  {32'hc49aa11c, 32'h4415d88b, 32'hc392e51f},
  {32'h43a96eb8, 32'h420169c5, 32'h43cbd48d},
  {32'hc3dee0a9, 32'hc43b8d0a, 32'hc52bf8fb},
  {32'hc32a07dc, 32'hc48fe095, 32'hc2031f1e},
  {32'hc35d4235, 32'h4440f463, 32'h4391b5b4},
  {32'h44a4ae26, 32'hc410d867, 32'hc4026954},
  {32'hc49864dc, 32'h43bd5840, 32'h43b4ed27},
  {32'hc3c8abaa, 32'hc469420f, 32'hc3d5c511},
  {32'hc46db818, 32'h4370abf7, 32'h44f0a748},
  {32'h4409dad6, 32'h43d448e1, 32'hc296c617},
  {32'hc49063e4, 32'h4427de59, 32'h449824a8},
  {32'h44d8bf12, 32'h4483a312, 32'hc3d80856},
  {32'hc4892adb, 32'h440d10c1, 32'h433eedf8},
  {32'h44acb117, 32'hc43f2995, 32'hc3e983bc},
  {32'hc4fc571c, 32'h441fdd4d, 32'h42ccc406},
  {32'h431857bf, 32'hc4790991, 32'hc3d6e2b1},
  {32'h413f1b00, 32'h447b4c65, 32'h451cdaf5},
  {32'hc2b4d3e4, 32'hc4f1b6bb, 32'hc41f892c},
  {32'h44b3324c, 32'hc2e360ea, 32'hc500dd03},
  {32'hc43ee8c6, 32'hc345d205, 32'h44443d52},
  {32'hc318a540, 32'h44283252, 32'h43091a3e},
  {32'hc41814d5, 32'hc3a15f43, 32'hc3d2e2cf},
  {32'h43fc17fa, 32'h44b72718, 32'h4347822f},
  {32'h449c80d4, 32'hc24908da, 32'hc3817d49},
  {32'h4503166c, 32'h4480855b, 32'hc31427e5},
  {32'hc5328439, 32'hc2e37242, 32'h43c5ce1e},
  {32'hc329b781, 32'h44e36b5a, 32'h4371906e},
  {32'h43b21eb7, 32'h4248b578, 32'h4071edc9},
  {32'h443b62fa, 32'h418180a6, 32'h44226cd5},
  {32'hc3d3b444, 32'hc2eb24d8, 32'h43739569},
  {32'hc10156c0, 32'h44ac0cd3, 32'h4418ab99},
  {32'hc3a8be9c, 32'hc472e057, 32'hc45e901d},
  {32'h44f36a1c, 32'h440b9929, 32'h428bae33},
  {32'h40d0f588, 32'hc35cc72c, 32'hc5175176},
  {32'h44514a56, 32'h448c57e3, 32'h443e92fd},
  {32'h43ae76f3, 32'hc3822887, 32'hc49fd816},
  {32'hc3a0f98e, 32'hc30b9faf, 32'hc13c4d69},
  {32'hc556a3bd, 32'hc3a84c30, 32'hc37522b7},
  {32'h44e5b13c, 32'h4462484c, 32'h42e8fc07},
  {32'hc3d455e3, 32'hc4a12a19, 32'hc4274596},
  {32'h43fc9cf8, 32'h44af057e, 32'h43ccd1bc},
  {32'h44324a2c, 32'hc2df0870, 32'hc2e40f8e},
  {32'h449ff479, 32'h4491915b, 32'h449438dd},
  {32'hc463c4c1, 32'hc3474fe2, 32'hc53c8a2c},
  {32'hc1146bb0, 32'h44c933e9, 32'h43084c5a},
  {32'h44fa5045, 32'h433ec4a6, 32'hc3dc7b79},
  {32'hc430632a, 32'hc500913d, 32'hc3ed4c34},
  {32'h448c073a, 32'hc2cb64d9, 32'h44793421},
  {32'hc55dfad0, 32'h44556450, 32'hc2d506cc},
  {32'h442286dd, 32'h44ef495a, 32'h41ff8bd0},
  {32'h432753d8, 32'hc51454bb, 32'hc2c1f11b},
  {32'h446db2ec, 32'h42e565ea, 32'hc4267ffa},
  {32'hc587abad, 32'h4383e92e, 32'hc3a09630},
  {32'h44355e4b, 32'h44232170, 32'h4468c6de},
  {32'h44f95a9f, 32'h43bed695, 32'h439d7d41},
  {32'h423ae85c, 32'h451d70c3, 32'hc27c1854},
  {32'hc50be199, 32'hc3cc5ede, 32'h4377655d},
  {32'h4520043a, 32'h442c4978, 32'h4413f0f7},
  {32'hc40854b4, 32'hc4e0898b, 32'h443be8ed},
  {32'h44b46b26, 32'h4482b5b0, 32'hc2d33ba1},
  {32'hc43184bb, 32'h439ecc6e, 32'hc3702e61},
  {32'h448ec28b, 32'h435f453b, 32'hc4831818},
  {32'hc0c3fc59, 32'h4431869c, 32'h4544a4c5},
  {32'h441f4879, 32'h44975fbd, 32'hc37e1cfd},
  {32'hc43ed847, 32'hc48171d5, 32'h44413718},
  {32'hc4e6a461, 32'hc2c0c624, 32'h4302a323},
  {32'hc3f364c1, 32'h4522e3b8, 32'hc1ecefca},
  {32'hc4bef1ad, 32'hc333d730, 32'h446e57cc},
  {32'h448c943a, 32'h41900cfa, 32'hc4a5e2b5},
  {32'hc22d2ac0, 32'h43d4a083, 32'h45580583},
  {32'h44916731, 32'hc3290c29, 32'hc4d6a399},
  {32'h44199aac, 32'hc4cb7ac0, 32'h4300deb5},
  {32'hc4f89a2e, 32'h449a85fd, 32'h43cec316},
  {32'h451a9942, 32'h44108477, 32'hc26ba0eb},
  {32'hc52dd233, 32'h43cf0b33, 32'h43de1b4d},
  {32'h4480f93d, 32'hc4d17011, 32'h42bfc04d},
  {32'hc43b3023, 32'h446b180f, 32'hc39a4cba},
  {32'h44c4c2f3, 32'hc42d6a0b, 32'hc4214233},
  {32'hc587dfa6, 32'h435fcfdd, 32'h43c3b625},
  {32'hc412c8c9, 32'hc2a8f14b, 32'h43b82442},
  {32'hc5106ae5, 32'hc267ef2f, 32'h441b9d87},
  {32'hc19db7a0, 32'hc4993ecc, 32'hc334df7e},
  {32'h43c073d4, 32'h4421b05b, 32'hc34bd541},
  {32'h43f736fa, 32'hc3907542, 32'h4473f897},
  {32'hc380db2e, 32'h449c7dd3, 32'hc43895b3},
  {32'hc3cd837f, 32'hc50361d3, 32'hc1924466},
  {32'hc43391f8, 32'h4451a0f1, 32'h4485e96f},
  {32'h43f3fdac, 32'hbff367b0, 32'h44e968d5},
  {32'h4311643e, 32'hc3b410cc, 32'hc241b0a0},
  {32'h44ac876a, 32'hc48e58b3, 32'h4521802c},
  {32'hc3c0ff80, 32'h44cd44b0, 32'hc40c8e7a},
  {32'hc4433091, 32'h42a98706, 32'hc3aef8e0},
  {32'hc329ace0, 32'h44f019a4, 32'hc339126a},
  {32'h43340c7a, 32'hc420652a, 32'h448e5639},
  {32'h444365f4, 32'hc3d3518e, 32'hc5002db0},
  {32'h4536bcc8, 32'h43af873a, 32'h43b2fff6},
  {32'hc5955986, 32'hc1f532b4, 32'h42f9bfbb},
  {32'h45461e7a, 32'hc3e60df3, 32'hc40cd001},
  {32'h42d556ee, 32'h440d0577, 32'hc474c0a8},
  {32'h43253bb6, 32'h44ea9602, 32'h448a1697},
  {32'h433bc8c9, 32'h449d77f0, 32'hc44720cc},
  {32'hc46b2630, 32'h41c33cb4, 32'h4311a3ad},
  {32'h448c8f93, 32'hc3cb38e9, 32'h44941006},
  {32'hc4aaa9b8, 32'hc3e2d1d1, 32'hc417f460},
  {32'hc3e035de, 32'h42f2b280, 32'hc30f73f6},
  {32'hc3a702e4, 32'h4275b58d, 32'hc4b69db1},
  {32'h43196c58, 32'hc4188ec5, 32'h44ecfa00},
  {32'h4500c277, 32'h439e2b09, 32'h447da95e},
  {32'hc480cc3d, 32'hc46fdbf3, 32'hc3fac1f3},
  {32'h445296ef, 32'h43f1dc97, 32'h429d8142},
  {32'hc4497f0a, 32'h44008ff2, 32'h43b36ffb},
  {32'hc41fe82b, 32'h4390723e, 32'hc45d7faa},
  {32'h4391ae01, 32'hc4990749, 32'hc2fdb0d4},
  {32'h42033e76, 32'h4283ae66, 32'hc4f3eea0},
  {32'h428ce33e, 32'hc49e6991, 32'h4393eb98},
  {32'h438ce7b4, 32'h44acb44d, 32'hc48ccbfd},
  {32'hc49b3979, 32'h43554b3a, 32'h4300cdcc},
  {32'hc490f636, 32'hc3a5f851, 32'hc4690105},
  {32'h45010b65, 32'h4409a843, 32'h4380ca77},
  {32'hc4d4ad19, 32'hc2d7cf7d, 32'hc2bfa5e0},
  {32'h4305c1eb, 32'hc4a6925c, 32'hc3adc07d},
  {32'hc3190c84, 32'h442bcf12, 32'hc30a21c9},
  {32'hc3215a1d, 32'hc4b86224, 32'hc3ead884},
  {32'hc480717a, 32'h4515e8f7, 32'hc3c3f2ff},
  {32'hc218cb04, 32'hc56cf526, 32'h43c9a747},
  {32'hc3c1216f, 32'h4268ce57, 32'h443a1a94},
  {32'h4318088c, 32'hc45956b7, 32'hc4700d9c},
  {32'hc4a91654, 32'h4421d75a, 32'h442dbdad},
  {32'hc415cea0, 32'hc46d92d4, 32'h439a0e30},
  {32'h44110bf5, 32'h422895dd, 32'hc5017d2e},
  {32'hc3cc9a54, 32'h4258a911, 32'h449c5db4},
  {32'h4489e30a, 32'h44b0dc76, 32'hc411f3e5},
  {32'hc2813643, 32'hc4ed516e, 32'h439112ba},
  {32'h43f1d5da, 32'h441fa6c0, 32'h4403e39e},
  {32'h4287e512, 32'hc3e442d5, 32'h43c1d13a},
  {32'hc4841f4c, 32'hc3ad6115, 32'hc2bcc55d},
  {32'h44c05378, 32'h4450a25c, 32'hc420468f},
  {32'hc3e640ac, 32'hc2c131ea, 32'h44e76599},
  {32'h442623f1, 32'h4331fd70, 32'hc478616d},
  {32'hc498b7d2, 32'hc4bc733e, 32'h4401a2ee},
  {32'h44bb3f04, 32'h43b6ecac, 32'h42143c90},
  {32'h4486a306, 32'hc39047c6, 32'h447db677},
  {32'h4468332e, 32'h441163b5, 32'hc3eaf856},
  {32'hc5016683, 32'h43d3c179, 32'hc3a13ade},
  {32'h453aafae, 32'hc381998c, 32'h3f66d540},
  {32'hc3be5758, 32'hc41f1a86, 32'h43eebba5},
  {32'h4580f5fe, 32'h43238608, 32'h43d88c51},
  {32'hc5264cc6, 32'hc33df756, 32'h43b85a22},
  {32'h44ae2eb1, 32'h43dd5568, 32'hc3288fae},
  {32'h429f8648, 32'hc5425fb9, 32'h43b67749},
  {32'hc4e52238, 32'hc3e32567, 32'h43848c46},
  {32'h441dc311, 32'hc48a66c9, 32'h449d5a4e},
  {32'hc40088c9, 32'hc2ea066a, 32'hc480ebc0},
  {32'hc34b20b9, 32'hc39790f9, 32'h45094764},
  {32'hc42d9c4b, 32'h4341f4ca, 32'hc41b6286},
  {32'h44aaea30, 32'hc2eef61f, 32'h44a7ffc1},
  {32'h43a526ce, 32'hc1fb72c2, 32'hc5098805},
  {32'hc2b05df0, 32'h44687a35, 32'h4443cbfe},
  {32'hc3864808, 32'hc426f76a, 32'hc4f07e19},
  {32'h4332f758, 32'h44be8bcf, 32'h44da21c7},
  {32'h43a80cfa, 32'h4495b48c, 32'hc3a85b17},
  {32'h449dbb90, 32'h4395eac5, 32'h42dfde08},
  {32'h43420078, 32'hc4d51cec, 32'hc445029e},
  {32'hc4e7ec46, 32'hc222c431, 32'h43f07894},
  {32'hc405904b, 32'hc4be93f6, 32'hc1d0080c},
  {32'h44bbed48, 32'h4396e5ee, 32'h4401575d},
  {32'h434f42a0, 32'hc435eb0d, 32'hc4b563f0},
  {32'hc0726000, 32'h4404c0d7, 32'h450d20e5},
  {32'hc396b68e, 32'hc3e73429, 32'hc58895da},
  {32'hc49451ec, 32'h4386de5f, 32'h42dfa759},
  {32'hc58af7fe, 32'hc302560f, 32'hc2896540},
  {32'hc39029f4, 32'h448dcff1, 32'h405674b4},
  {32'h44a582ee, 32'hc370627c, 32'hc0faba74},
  {32'hc2320544, 32'h454e1011, 32'hc2184fb4},
  {32'hc482c9cc, 32'hc47b3b1c, 32'h42bb6a44},
  {32'h454292eb, 32'h43c8c866, 32'h4402954b},
  {32'hc58f64d7, 32'h4205be00, 32'hc3645b5a},
  {32'h45124278, 32'hc3977382, 32'h433cc727},
  {32'h44fca7ff, 32'hc33f775f, 32'hc312871b},
  {32'h439ec164, 32'h4351eac6, 32'hc22c5290},
  {32'hc3e0db88, 32'hc3293168, 32'hc4a84fed},
  {32'hc49c9271, 32'h43828f54, 32'h4385606d},
  {32'hc1bf8b20, 32'hc4b3ddd9, 32'hc4b0fa61},
  {32'hc37dd28d, 32'h43b815e0, 32'h44b7e3f0},
  {32'h44651942, 32'hc35d49e3, 32'hc40c25bf},
  {32'hc215fa38, 32'h443b291c, 32'h45248a46},
  {32'hc4854896, 32'h435fa0cb, 32'hc482f695},
  {32'h4226c5b0, 32'hc446dd7a, 32'h44887ece},
  {32'hc3f59038, 32'h445d2011, 32'hc545e026},
  {32'h41add6cd, 32'hbf4dac53, 32'h44ba2140},
  {32'h445cdfe7, 32'h413562cd, 32'hc48a95ab},
  {32'hc3f96712, 32'h44bb6a8d, 32'h438c8224},
  {32'h43a57e1b, 32'h43cec73e, 32'hc436778b},
  {32'hc3d5bf50, 32'h44a3b61a, 32'h449a91c7},
  {32'h438d7202, 32'hc41752ca, 32'hc4268ed7},
  {32'h442f57ee, 32'h44086285, 32'h443abf36},
  {32'h440b3c60, 32'hc456c718, 32'hc45d98db},
  {32'hc5379f5d, 32'h432f6bb5, 32'hc189138f},
  {32'hc3968f88, 32'hc1288862, 32'h431db9e7},
  {32'hc3dce63c, 32'h451f285a, 32'hc4164b8e},
  {32'h451621e3, 32'hc46b1f38, 32'h4168aed3},
  {32'hc53658be, 32'hc378f57a, 32'h429f8558},
  {32'h450ab607, 32'h43843be5, 32'h4407af83},
  {32'hc5878fb2, 32'h419af276, 32'hc3f9b78e},
  {32'hc50936d9, 32'h43858da6, 32'h430af982},
  {32'h42885c60, 32'hc3b00ffc, 32'h43be5751},
  {32'hc3d76dd2, 32'h44370176, 32'hc517c4b5},
  {32'hc1c39f00, 32'hc4055b33, 32'h448c5ca1},
  {32'hc531ccf0, 32'hc47045d0, 32'hc3fd7725},
  {32'h451dc37e, 32'hc406ba8e, 32'h422e5a6f},
  {32'hc4bacff8, 32'h4427d7c9, 32'h42336e08},
  {32'h4478657c, 32'hc4213d96, 32'hc3597c50},
  {32'hc4beaed0, 32'h43e2ee29, 32'hc38bbacc},
  {32'h43f1a9b6, 32'hc40ece32, 32'h421ec08b},
  {32'h44786687, 32'h43c9a711, 32'hc4354819},
  {32'h4429b4b0, 32'h4385bd57, 32'h44a37aa6},
  {32'hc5058cd9, 32'h4435263f, 32'hc27bed72},
  {32'hc4cddb7e, 32'hc376305e, 32'hc4039fcd},
  {32'hc4df45c4, 32'hc31d260d, 32'h44099cf4},
  {32'h42b8e02c, 32'hc4b40d3b, 32'hc4152764},
  {32'hc42581c5, 32'h43452a6c, 32'h43f77f78},
  {32'h427f6f60, 32'hc1d226e5, 32'hc52531eb},
  {32'hc438791d, 32'h42abcd8f, 32'h44eb412d},
  {32'h4494c944, 32'hc3888521, 32'hc381908f},
  {32'hc573333c, 32'h4396a183, 32'h426d25c3},
  {32'h454eec96, 32'h43c57da3, 32'hc4429b8e},
  {32'hc4901d71, 32'hc43f4a62, 32'hc405754a},
  {32'h43843c80, 32'hc51c3e54, 32'h42838acb},
  {32'hc47bee98, 32'h433daa28, 32'h439fdcd4},
  {32'h43093c86, 32'hc4b2d88b, 32'hc374028c},
  {32'hc33309d4, 32'h44f83183, 32'h442e96bd},
  {32'h43620cb0, 32'hc4a15e34, 32'hc49518e3},
  {32'h44605bae, 32'hc2b5e98a, 32'hc4813839},
  {32'hc403cc42, 32'hc2dbaa56, 32'h4538d29b},
  {32'h448f1170, 32'h42fe8306, 32'hc40e8752},
  {32'hc457964a, 32'hc3f2ac61, 32'h439f5b42},
  {32'h4478b15a, 32'h44770872, 32'hc3557855},
  {32'hc5019f55, 32'h43db4c25, 32'h4204f476},
  {32'hc2880bc0, 32'h45124fc3, 32'hc30a42a2},
  {32'hc3faf2c0, 32'hc426786e, 32'hc29c2020},
  {32'h452dce33, 32'h4359ab87, 32'h44469133},
  {32'h4345fd20, 32'hc40eb1c4, 32'h445ce5b0},
  {32'h44d3d4da, 32'h422a28f7, 32'hc4924046},
  {32'hc483eff0, 32'hc3e3bd73, 32'h439a180c},
  {32'h44b7cc1d, 32'h415a95ce, 32'h44aa9077},
  {32'h42820106, 32'hc53482d5, 32'h42a5b67a},
  {32'h44ad1d7c, 32'h43673a18, 32'hc35d730a},
  {32'hc39d8b47, 32'hc48128ab, 32'hc4be0fe9},
  {32'h43bb8840, 32'h43dac9e1, 32'h4530ebb7},
  {32'hc381e3fd, 32'hc4aedbc5, 32'hc2ffdded},
  {32'h441e4a94, 32'h4469a618, 32'h44b4285e},
  {32'hc54574cd, 32'hc30ba560, 32'hc38d517d},
  {32'h4497c3a0, 32'h435193a8, 32'hc400d059},
  {32'hc3cf2940, 32'hc4206b02, 32'hc487bf19},
  {32'hc37389e8, 32'h4535dd13, 32'hc35c3538},
  {32'h4441d6d6, 32'hc3a1fdd9, 32'hc4622874},
  {32'h451441a8, 32'h437c21d1, 32'h4406c5fc},
  {32'hc4e0ab6c, 32'hc481fdf7, 32'hc420756d},
  {32'hc3fb2904, 32'hc3064e7f, 32'h43440e77},
  {32'h43a580e2, 32'h438f93a2, 32'h44010420},
  {32'hc435eadd, 32'hc41b9dc0, 32'hc4203603},
  {32'hc3437cf9, 32'h450fcf44, 32'hc38473e9},
  {32'h4482ae5c, 32'hc302ec65, 32'h42f3df7e},
  {32'h44a3f92f, 32'h43eb15bc, 32'hc24621f7},
  {32'hc4988c80, 32'hc4c9dce0, 32'h438fbee3},
  {32'h44826e69, 32'h4395420e, 32'hc3ff5408},
  {32'hc55293ba, 32'h439588cd, 32'hc23d1cd2},
  {32'h44b86272, 32'hc4614316, 32'hc3db48a6},
  {32'hc4cebff1, 32'h43d9cb7b, 32'h4327c9a0},
  {32'h44410483, 32'h442173a3, 32'hc3f9bf58},
  {32'hc4249be8, 32'hc3d4d81f, 32'h44aa22b4},
  {32'h441a3074, 32'h448460c9, 32'hc2d6e293},
  {32'hc49ef647, 32'hc3c43f1a, 32'h440f0496},
  {32'h4497e34c, 32'h43e05651, 32'hc46d037e},
  {32'hc528acd8, 32'hc2aa285d, 32'hc3a875f9},
  {32'h44dff008, 32'hc211ced8, 32'hc3fe95d0},
  {32'hc41b78d9, 32'h43cc0ffa, 32'h433c6503},
  {32'h44074e3f, 32'h442da1bd, 32'hc4479c29},
  {32'hc425e39b, 32'hc4997804, 32'h448f9a45},
  {32'hc4f84bf2, 32'h432826c0, 32'hc3c07524},
  {32'h43a41f34, 32'h4358a557, 32'hc53a6ba6},
  {32'hc5476c2d, 32'h42819a6d, 32'h43a953b5},
  {32'hc4d9abae, 32'h42e89010, 32'h425407d5},
  {32'hc42e49b8, 32'h42ffd2d2, 32'h4518b1c7},
  {32'h42b05f80, 32'hc2bf5e6e, 32'hc30a6aef},
  {32'h4441c7bf, 32'hc5474067, 32'hc329cfba},
  {32'hc41afc34, 32'h446a58cc, 32'h4409ceac},
  {32'hc3b2723c, 32'hc4a051aa, 32'hc24b7c18},
  {32'hc5231244, 32'h43daffef, 32'h43de9ab4},
  {32'h4534f5c3, 32'hc3930cb2, 32'hc34f7da2},
  {32'h4401bbf7, 32'h4429e7af, 32'hc32b6a88},
  {32'h4505c695, 32'hc3e91975, 32'hc3f89d88},
  {32'hc500e26e, 32'h43c14b45, 32'h43cb291d},
  {32'hc3ffa11a, 32'hc294a4a3, 32'h432b4f2e},
  {32'hc4243145, 32'h44331eff, 32'hc5076a06},
  {32'h43aba598, 32'hc482ed84, 32'h44795739},
  {32'h4404f9b0, 32'hc395c18d, 32'hc2ef7985},
  {32'hc2cb0a00, 32'hc482d6de, 32'h44ca913a},
  {32'hc4606e1e, 32'h44d5cd1a, 32'hc3fa7978},
  {32'h44367f42, 32'h4218f9e8, 32'h44101b6b},
  {32'hc3ea5671, 32'h43f7d3c3, 32'h442fe08d},
  {32'h440a36f4, 32'h424baa6a, 32'h44d63ed6},
  {32'hc466125c, 32'h43b9c346, 32'h4403d542},
  {32'h44ea4d7c, 32'hc445f195, 32'hc4035836},
  {32'hc4a5843a, 32'h44b3a186, 32'hc4e25463},
  {32'h4407eb9f, 32'hc39da5a0, 32'hc35681b3},
  {32'hc2df51e8, 32'h44c3edd9, 32'hc40aac63},
  {32'h4498c27c, 32'hc2f8efc8, 32'h443230c5},
  {32'hc4f126de, 32'h43942791, 32'hc39b9906},
  {32'h43bc4278, 32'h439675a8, 32'h444426b8},
  {32'hc4e34ae8, 32'h44097922, 32'hc46c11ba},
  {32'h44c6d392, 32'h434950cb, 32'h4325a2a7},
  {32'hc3b41622, 32'hc48b1547, 32'hc44bb298},
  {32'hc3b45be8, 32'h449fed37, 32'h44e4da9c},
  {32'h44eeeafb, 32'hc3d4a61d, 32'hc31b58c4},
  {32'h44a7efce, 32'h432538c0, 32'hc1e39ada},
  {32'h44c407e3, 32'hc2996907, 32'h44766a83},
  {32'hc3953ebe, 32'h43463b32, 32'hc4c77361},
  {32'h448335e7, 32'h43b096b5, 32'hc1d1d5a8},
  {32'hc50c7b0f, 32'hc194ccd2, 32'hc3f48ef0},
  {32'h42b3d820, 32'h42136952, 32'h455db3ea},
  {32'hc4396585, 32'h44414bc4, 32'h4547a36b},
  {32'hc31c4e5e, 32'h442950da, 32'hc4ed63c4},
  {32'h4514ba05, 32'h428d3a5e, 32'hc1891926},
  {32'h450816e1, 32'hc3103107, 32'hc3250d44},
  {32'hc3585cbd, 32'hc30fd8d3, 32'hc42fe75d},
  {32'h44ff1e0a, 32'h4414aa8a, 32'h431cde3a},
  {32'h449998a4, 32'h446b215e, 32'hc37b1105},
  {32'h438d385c, 32'hc34fd96b, 32'h442939d5},
  {32'h42a8c79e, 32'h44d09e27, 32'hc46748a8},
  {32'hc48aeb2c, 32'hc383dcf5, 32'h42fb4c0b},
  {32'hc5991f68, 32'hc2b5aa34, 32'hc3cc87c3},
  {32'h44b7dba4, 32'hc408d96f, 32'hc36d7400},
  {32'hc4caefcf, 32'h431a2e57, 32'hc3925132},
  {32'h4471ba86, 32'hc4aaee84, 32'h43e2eb26},
  {32'hc4cfea95, 32'h4440c77a, 32'hc2e710fc},
  {32'hc411f9af, 32'hc3c47f54, 32'h4363b98b},
  {32'hc526401c, 32'h431bb9e4, 32'hc3ce110c},
  {32'h43a2c720, 32'hc49f581f, 32'h434379e2},
  {32'h44b7cc1e, 32'hc45bf272, 32'h43165b7a},
  {32'h443626ac, 32'h4481616b, 32'hc4276f9d},
  {32'hc464ba28, 32'hc4614107, 32'h444a3c8d},
  {32'hc309760e, 32'hc25f47b1, 32'h43ebbdf0},
  {32'h4338caef, 32'h4378489f, 32'hc1a5b567},
  {32'h412dae38, 32'hc48052bb, 32'h43e944b4},
  {32'h43e4c936, 32'h448d028e, 32'hc4a07104},
  {32'hc386d633, 32'hc527c4c0, 32'h43472bc4},
  {32'h44b898be, 32'h434474fe, 32'h43fbcc60},
  {32'h43d1cdf1, 32'h44d3b54b, 32'hc45d4923},
  {32'hc4152858, 32'hc340e6ac, 32'h44d58598},
  {32'h451b4ff6, 32'h43e91323, 32'hc3b4da55},
  {32'hc4199c14, 32'hc438f20a, 32'h44584bf2},
  {32'h4406f6f2, 32'hc29301a9, 32'hc46f0ea8},
  {32'hc4a1d900, 32'hc4470ebb, 32'h44254dc2},
  {32'h446097d7, 32'hc316af60, 32'hc3be56b5},
  {32'h43b1df23, 32'h425138fb, 32'h44c96b1e},
  {32'h456a2415, 32'hc2b397e5, 32'h43ffdeea},
  {32'hc4f864a2, 32'h431edf5a, 32'h44299ed2},
  {32'h44d9ae6e, 32'h43d2f931, 32'hc30cafb2},
  {32'hc4364300, 32'hc51ad3ce, 32'h430b89af},
  {32'h453fc5b0, 32'h42c5ea41, 32'hc39e1b57},
  {32'h43dc1f8e, 32'hc33f375a, 32'h43aaeef1},
  {32'h44a58fb6, 32'h44b7aa76, 32'hc369a9a9},
  {32'hc471cbfc, 32'hc4d029f0, 32'hc4017a75},
  {32'hc2cfe55e, 32'h44b3e4f7, 32'hc38ee477},
  {32'h433acaea, 32'h4286e58b, 32'hc34ea53c},
  {32'hc3a95c34, 32'hc45ae8bf, 32'hc4033243},
  {32'hc296d01c, 32'h41c8910c, 32'h44b87953},
  {32'h43047ce8, 32'hc21a412a, 32'hc505d13c},
  {32'h431770e0, 32'h446fb4af, 32'h4429f6e4},
  {32'hc3eb8755, 32'hc26bd764, 32'hc494b658},
  {32'h44302819, 32'h4421e6c5, 32'hc36d822e},
  {32'hc36a9790, 32'hc4122f78, 32'hc508b9c3},
  {32'h44edef6b, 32'h43c63e94, 32'h4410019b},
  {32'hc3f00830, 32'hc432ab02, 32'h42eb4352},
  {32'h44aaff3b, 32'h43877687, 32'h4316ef1e},
  {32'h4386aa67, 32'hc36d610c, 32'hc4aabe58},
  {32'h448f813f, 32'h44053c69, 32'h442ca879},
  {32'hc50e61e6, 32'hc1ed34fb, 32'hc3879fcd},
  {32'hc3a2b624, 32'h4421f554, 32'h450f852d},
  {32'hc5282af9, 32'hc397af14, 32'h43c0e237},
  {32'h440ceca3, 32'h4410c727, 32'h45038056},
  {32'hc30e7d1b, 32'hc4d631f2, 32'hc4e80b91},
  {32'h44a86118, 32'h440b15f4, 32'h42fef7f0},
  {32'hc4e8b6f2, 32'hc42d6335, 32'hc2f241c6},
  {32'h44198664, 32'h44df0c28, 32'h4416acc1},
  {32'hc5358344, 32'hc2865260, 32'h422dbd45},
  {32'h43fffc90, 32'h44769fd6, 32'h440618af},
  {32'hc3fd83e8, 32'hc4289260, 32'h420cad80},
  {32'h442ff54b, 32'h43c09538, 32'h43fc31fa},
  {32'hc52df875, 32'hc41c78b6, 32'hc2c027f9},
  {32'h44fd3211, 32'hc31125d3, 32'hc2bdd2bc},
  {32'h437d36ad, 32'hc42a1199, 32'hc49491f2},
  {32'h43612694, 32'hc37f91bc, 32'h4500818f},
  {32'hc2a991ec, 32'hc2d18c44, 32'hc3f46f88},
  {32'hc4f6a5da, 32'h4450acd8, 32'h43268f9d},
  {32'h45018e3b, 32'h42e7afc0, 32'h431c0a4c},
  {32'hc23938d8, 32'h45129826, 32'h43f93ae1},
  {32'h42f50390, 32'hc48599bb, 32'hc525502e},
  {32'hc33cf511, 32'h43f1ad73, 32'h455899d1},
  {32'h44976700, 32'hc42bbb54, 32'hc322289b},
  {32'hc4880522, 32'h41930b58, 32'h443c21f1},
  {32'hc3a14d22, 32'h44fcf1a6, 32'hc4a906e3},
  {32'h43638d9e, 32'h432c6e5e, 32'h4412223c},
  {32'hc35c82e8, 32'hc479886d, 32'hc4a91b99},
  {32'hc49ed775, 32'h43070361, 32'h43d6c1b9},
  {32'hc415f67b, 32'hc4817eaa, 32'hc2abb0d3},
  {32'hc52e112e, 32'h4297703e, 32'h4317ea4a},
  {32'hc384aad0, 32'hc370aa9c, 32'hc4daefa6},
  {32'h4422c384, 32'h43c97f5e, 32'h442694fc},
  {32'h449fd13e, 32'hc4a32a1d, 32'h425679c6},
  {32'hc54c2d6a, 32'h441dc142, 32'hc36eda7e},
  {32'h44d6dd42, 32'h43607ba0, 32'h4105129c},
  {32'hc4c306d5, 32'h448df119, 32'hc2525dfa},
  {32'hc31b21f9, 32'hc517a281, 32'h43b35262},
  {32'h44fe12f2, 32'hc275c6cf, 32'hc3ea4ddf},
  {32'h4498e705, 32'h43b95a47, 32'hc20b8d94},
  {32'hc4e1e7a6, 32'hc3e0298b, 32'hc36e686f},
  {32'h432c89fd, 32'hc4278773, 32'hc3a77e2b},
  {32'h43d90e5f, 32'hc3021ab5, 32'hc283ef28},
  {32'hc569c2e0, 32'h4397cf0a, 32'h43332960},
  {32'h451d5cc4, 32'h4322ad5c, 32'h4352e7ca},
  {32'hc3906988, 32'hc3909ccc, 32'h43b4d17f},
  {32'h43ed2b30, 32'hc5403281, 32'hc32b02ff},
  {32'hc4897076, 32'h444c58d7, 32'h42538452},
  {32'h43b2cd01, 32'hc47b4a88, 32'h4362b824},
  {32'hc530b943, 32'h440ac6bf, 32'h432097ec},
  {32'h44af091e, 32'hc4acfb2f, 32'h414da81e},
  {32'h443822f7, 32'hc1818452, 32'hc464df64},
  {32'h4513d2c6, 32'h420e6ef2, 32'h42dcf507},
  {32'hc5060d67, 32'h43fcad82, 32'hc3098195},
  {32'h42e7983b, 32'hc33babfb, 32'hc48fbf4e},
  {32'hc3265268, 32'h4495a2b7, 32'h447e45e3},
  {32'h4411e238, 32'hc41914ec, 32'hc47110c7},
  {32'h41ef3842, 32'h44f5b4b1, 32'h439781bb},
  {32'hc30a945c, 32'hc409659b, 32'hc423d030},
  {32'hc4e49577, 32'h4311ed21, 32'hc24a42ec},
  {32'h4513052f, 32'hc323a028, 32'h4355b188},
  {32'hc410d4e8, 32'h422d88e6, 32'h433d4210},
  {32'h443cd9e6, 32'hc4a8e182, 32'hc4e54074},
  {32'hc52ffa60, 32'h4339e3ea, 32'hc41987db},
  {32'h442e9f60, 32'hc45403de, 32'hc4914f60},
  {32'hc3b2753e, 32'h44303033, 32'h444bdbae},
  {32'h452f6a1a, 32'h4346771d, 32'hc3d2308c},
  {32'hc561b85e, 32'h44600eb0, 32'hc18ce0b9},
  {32'h42487aa6, 32'hc541685f, 32'hc3039bdc},
  {32'h449e354e, 32'h42f16458, 32'hc50b673f},
  {32'hc52c8610, 32'h41f30cf5, 32'h44157b60},
  {32'h4202f6f0, 32'hc28e9bc5, 32'h435b4c40},
  {32'hc302c370, 32'hc530ddee, 32'hc14e4005},
  {32'h43a172f8, 32'h451b0a05, 32'h433aebfa},
  {32'hc4cfd789, 32'hc366708e, 32'hc397b506},
  {32'h44521bf9, 32'h44ab9916, 32'h431f92ee},
  {32'hc551fc32, 32'hc4377e2f, 32'h43eb06d7},
  {32'h4460c29a, 32'h4453e449, 32'hc2e61bbd},
  {32'hc4aa8c0b, 32'h432a3b42, 32'h4405fb25},
  {32'h453d34b6, 32'hc3953c54, 32'h42842c42},
  {32'h44c6aafa, 32'h43a22bd1, 32'h440e1cca},
  {32'hc2ee5953, 32'h44cba3ec, 32'h4399ef99},
  {32'h43759f89, 32'hc4a950fa, 32'h43579239},
  {32'h44334528, 32'h4414175a, 32'h439f367a},
  {32'hc38782ca, 32'h424fddd5, 32'hc53403bc},
  {32'h441e737a, 32'h4488a686, 32'h44694fe2},
  {32'hc503d0f5, 32'hc3dc831b, 32'hc43ed30b},
  {32'h45214aef, 32'h4437b20e, 32'h446dce37},
  {32'hc48f759c, 32'hc4368bdf, 32'hc4b09d42},
  {32'h42c498e0, 32'hc313123a, 32'hc38a5a0d},
  {32'hc456db98, 32'h3ff672f6, 32'hc403446f},
  {32'h446d723c, 32'h43b75115, 32'h43185f75},
  {32'h44bafdc7, 32'hc22bfb7f, 32'hc387d2c3},
  {32'hc2f9316f, 32'h44af20db, 32'h44c614b7},
  {32'hc4a13f8c, 32'hc31b9a38, 32'hc4db0174},
  {32'hc28eb2ba, 32'h44b49483, 32'h44005921},
  {32'h444845ec, 32'hc4372abb, 32'hc37fcad3},
  {32'hc3c635f4, 32'hc4f39730, 32'hc325afd8},
  {32'h4336eabe, 32'h45503bb7, 32'hc3ac1417},
  {32'h429ad5e0, 32'hc4c24f93, 32'h42867884},
  {32'h450745ec, 32'h44355798, 32'hc3d27d87},
  {32'hc5251233, 32'hc4112884, 32'h4198adea},
  {32'hc47a98f3, 32'h438292f8, 32'hc332ef0d},
  {32'hc46f1745, 32'h44302d04, 32'hc282eb86},
  {32'h44658e28, 32'h4483158a, 32'h4487979e},
  {32'h432087ca, 32'hc284a1b1, 32'h44cd0e9c},
  {32'h433dcc63, 32'h448fd331, 32'hc3d676a0},
  {32'hc3673dd2, 32'hc3abf8a9, 32'h44fb6001},
  {32'h4120257e, 32'h44bdf42e, 32'hc3a7c0cd},
  {32'hc4bd11cb, 32'hc3a32e02, 32'h43f4cf61},
  {32'h44b299ca, 32'h41d2794a, 32'hc2ec87a8},
  {32'h441de8c4, 32'hc3588f14, 32'h4467aacc},
  {32'h44cd817d, 32'hc1c488d2, 32'hc47df5e6},
  {32'hc4a05813, 32'hc3274d23, 32'h441c2cb4},
  {32'hc4996bf5, 32'hc2e907ca, 32'hc43d0f6e},
  {32'hc434672a, 32'hc52b1435, 32'h444f4758},
  {32'hc35321c3, 32'hc208744e, 32'h40d07dcf},
  {32'h45075b26, 32'h4396ed5b, 32'hc36ba901},
  {32'hc508e893, 32'hc423ee49, 32'h44305217},
  {32'h441c2f94, 32'h43196cbe, 32'hc3eabfe1},
  {32'hc4880682, 32'h43162986, 32'h44d94a84},
  {32'h45159c96, 32'h43c41689, 32'hc43fe7fa},
  {32'h42f80616, 32'hc53333a2, 32'hc3149c3d},
  {32'hc32efb0a, 32'h443368f3, 32'h446f62a8},
  {32'hc3b1d3df, 32'hc4dcf506, 32'h429a9d8d},
  {32'hc504bcc3, 32'h4488de4a, 32'h4216e98c},
  {32'hc38d920a, 32'hc56c138e, 32'h42f05f0e},
  {32'hc5274317, 32'h4307a764, 32'hc30edb79},
  {32'h447c1048, 32'h43851739, 32'h4280ae52},
  {32'hc542d1d8, 32'h43811c13, 32'hc3177c94},
  {32'h44256908, 32'hc44e1bb2, 32'hc20ad027},
  {32'hc4455bee, 32'h440262b1, 32'hc493f69b},
  {32'h436dfd8d, 32'hc3f2fdc6, 32'h45166d4e},
  {32'hc404f643, 32'h43d8270d, 32'hc43e573d},
  {32'h43b245b8, 32'h42d79831, 32'h4513045c},
  {32'hc3bf1470, 32'h4346c6b6, 32'hc531c682},
  {32'hc38ed6bb, 32'hc499338a, 32'hc38ccdb3},
  {32'hc4c61396, 32'hc210f8dd, 32'hc446fe63},
  {32'h45095c36, 32'h43b3cf50, 32'h43a68a50},
  {32'hc51f064e, 32'hc28d4d88, 32'h438509c3},
  {32'h44320292, 32'hc4bf493b, 32'h43e6078a},
  {32'hc50599de, 32'h44bd22f4, 32'hc37d6b97},
  {32'hc41bf926, 32'hc439720e, 32'hc2542ef2},
  {32'hc3ba1680, 32'h439fc8bb, 32'hc513832b},
  {32'hc22fff10, 32'hc3c345c3, 32'h43edf663},
  {32'h439e7a55, 32'hc41a1ab6, 32'hc4faceee},
  {32'h44b143d4, 32'h4447a323, 32'h443c2de4},
  {32'hc4dd1cc9, 32'hc3993abb, 32'hc4a03127},
  {32'hc39dea90, 32'hc310316d, 32'h447ab166},
  {32'hc44cf1a0, 32'h4302598f, 32'hc44f8a5b},
  {32'h44160063, 32'h44968943, 32'h446ae494},
  {32'h43d21834, 32'hc3c8cb7f, 32'h3f740a60},
  {32'hc4553fd8, 32'h4335a6a6, 32'hc386d584},
  {32'h42ffd53a, 32'hc50699cb, 32'hc392edd1},
  {32'hc3e4131d, 32'h43df6fc3, 32'hc4b4db98},
  {32'h448fe92b, 32'h43e0042b, 32'h4113151a},
  {32'hc3bfe02a, 32'h44a355d6, 32'hc3c52768},
  {32'h450aa9ce, 32'hc3bce3c2, 32'h44320970},
  {32'h43a52946, 32'h447fd318, 32'h44a0a248},
  {32'hc527b073, 32'h44848157, 32'hc43139f8},
  {32'hc3fe7140, 32'hc2311a9f, 32'h44d14be0},
  {32'h4515f99f, 32'h43f0337b, 32'hc3ea2640},
  {32'hc35f7343, 32'h45158238, 32'h4399ba8d},
  {32'h440dd693, 32'hc4d494f8, 32'hc287db85},
  {32'hc39f5511, 32'h42dbc8a1, 32'hc5091b2a},
  {32'h43ae4c84, 32'hc507186b, 32'hc337598d},
  {32'h42268c8a, 32'h43903d21, 32'hc50f5fec},
  {32'hc41fa802, 32'hc3aa8bcf, 32'h431763cc},
  {32'hc44443cb, 32'hc1be2389, 32'hc46deb68},
  {32'hc38c24bc, 32'h4413336a, 32'h445d5214},
  {32'h42efe5d3, 32'hc30e1f6f, 32'hc38b5b42},
  {32'h4559eba5, 32'h44622162, 32'hc2165cc3},
  {32'hc4d21246, 32'h4448df28, 32'hc100e82e},
  {32'h454bf55d, 32'h433de8a2, 32'h42f8481b},
  {32'hc4e62ffa, 32'h4486e7cc, 32'hc3b5ec24},
  {32'h4404abb5, 32'hc4b57221, 32'h432aa834},
  {32'h43d67a94, 32'h43fd62cd, 32'h441d370b},
  {32'h4312e678, 32'h44050d01, 32'hc5273e31},
  {32'hc4240941, 32'h4442d5f6, 32'h447c5582},
  {32'hc3eddbfc, 32'hc2cb8079, 32'h44dbadcc},
  {32'h43d475f0, 32'h438f0f55, 32'hc4b46ec3},
  {32'h4401c933, 32'hc5020ebc, 32'hc375639a},
  {32'h43dae384, 32'h4529bd15, 32'hc3b6f155},
  {32'hc3d1e375, 32'hc4a55001, 32'h43e911d9},
  {32'h436bb9ec, 32'hc3475957, 32'hc26903e7},
  {32'h431ca734, 32'h446d77b8, 32'hc3c03831},
  {32'hc3c3e3d4, 32'h43f79f9c, 32'h44e71bf4},
  {32'h43dfe4f0, 32'h43b8670f, 32'hc4b76e00},
  {32'hc380306c, 32'hc4339e2f, 32'h44568bef},
  {32'hc50afb4b, 32'h42d1ecdc, 32'hc32f2cf2},
  {32'hc4435498, 32'hc2a54385, 32'h44be3502},
  {32'h4364c814, 32'h44742418, 32'hc457474a},
  {32'hc4fe0942, 32'hc28aace0, 32'hc2dc97f9},
  {32'h44f813af, 32'hc3acddc6, 32'hc3f65044},
  {32'hc51f9566, 32'hc292d4dc, 32'hc34ebacf},
  {32'hc4e3bab8, 32'h430c85f1, 32'hc237c146},
  {32'h43089cd5, 32'hc5815268, 32'h434479ec},
  {32'h45020c48, 32'h421294fe, 32'hc234624a},
  {32'h44df57fc, 32'hc2abcdfe, 32'h43bb5996},
  {32'hc266e14c, 32'h453a6723, 32'h41357cf6},
  {32'hc524b4d2, 32'hc40d589f, 32'hc36ab0cc},
  {32'hc45c439e, 32'h442b8838, 32'hc3c56c89},
  {32'hc2b315e4, 32'h43cb4754, 32'h4380f93b},
  {32'hc496eeaa, 32'h4461282f, 32'hc323d2e3},
  {32'hc31f2a7a, 32'hc2fe5dd4, 32'h449969e7},
  {32'hc3587c5c, 32'hc405283b, 32'hc26eb964},
  {32'h44123e30, 32'hc371bac4, 32'h45247f9c},
  {32'hc483c0ee, 32'hc283ef2e, 32'hc49243a4},
  {32'h4524eb54, 32'hc2e36ed3, 32'hc3343ebd},
  {32'hc33030e0, 32'hc42a5839, 32'hc50dfd3d},
  {32'hc3c6abeb, 32'h44948416, 32'h4538a7f9},
  {32'h4415fd44, 32'hc4a345ee, 32'hc35864af},
  {32'hc0a43380, 32'hc104d13a, 32'h44c97fd3},
  {32'hc3f6f5ae, 32'h44a07f5d, 32'hc4e5a2eb},
  {32'hc440d7fa, 32'hc2593bf4, 32'h4481e02f},
  {32'h43a84a78, 32'hc498c087, 32'hc2c9b17c},
  {32'h439f6f31, 32'hc36726e6, 32'h410dac81},
  {32'h439602a5, 32'hc443ac6e, 32'hc4a8f2ae},
  {32'h44c18127, 32'h43bc2d23, 32'h44861c43},
  {32'h43da0c08, 32'hc321e15e, 32'hc4b69932},
  {32'h4487de5e, 32'h441e4709, 32'h4413ed04},
  {32'hc56b66e9, 32'hc44d098d, 32'hc3b8f0ae},
  {32'h4502338f, 32'h446d20a7, 32'h4432b9aa},
  {32'h442945d8, 32'hc4952bdc, 32'hc4008cf8},
  {32'h4480e372, 32'hc14adfb0, 32'hc3474193},
  {32'hc4b69a94, 32'hc41ed1c2, 32'h439c27fb},
  {32'hc4854677, 32'hc3785718, 32'hc2d8aad0},
  {32'hc488493a, 32'hc403aba6, 32'hc20b4b0c},
  {32'h449d9643, 32'h438e9bba, 32'hc378c184},
  {32'h44368260, 32'hc4c4948a, 32'hc4848323},
  {32'hc4a6cfdb, 32'hc3d3df75, 32'h448006b4},
  {32'hc2e00c08, 32'h43f04993, 32'hc429bdc7},
  {32'hc4c77f3f, 32'h448a5824, 32'h43f7a934},
  {32'hc3e583c7, 32'hc41e83db, 32'hc50e656f},
  {32'hc342b96a, 32'h43c9e8d4, 32'h439c7fac},
  {32'h442756b0, 32'hc4630be3, 32'hc4a54371},
  {32'hc2dbfe27, 32'h44e26b27, 32'h44ce12e9},
  {32'hc419979e, 32'hc3b5edc7, 32'hc4ba9f1f},
  {32'h440d9a82, 32'hc4db04e6, 32'h4484e370},
  {32'h44282133, 32'h44813e5a, 32'hc49e9860},
  {32'h440bb057, 32'h443cca9e, 32'h435db257},
  {32'h4405c838, 32'hc380aee2, 32'hc456f9bd},
  {32'hc533c022, 32'h410c2391, 32'hc27dd34a},
  {32'h43cb4786, 32'hc37ffb84, 32'hc4acf5b9},
  {32'hc405950d, 32'h43cbb44d, 32'h44c965a0},
  {32'h43b55b7a, 32'hc4385609, 32'hc4a8b63b},
  {32'h44c92fe4, 32'hc359cc84, 32'h43653286},
  {32'h45237302, 32'hc47662bf, 32'hc2a7af5f},
  {32'hc53c165e, 32'h44685698, 32'h42f2bb7f},
  {32'hc437d959, 32'hc4a06ccf, 32'h4409b50c},
  {32'h42a0b82b, 32'h4503e461, 32'hc3efcec9},
  {32'h454b69a0, 32'h42991b3b, 32'hc32fc0ac},
  {32'hc372c4d0, 32'h44b073ba, 32'h4354875a},
  {32'h44c13266, 32'h4350c170, 32'h4261556a},
  {32'hc58b30d0, 32'h43a665af, 32'h43f1843b},
  {32'h457f89ad, 32'hc34b2df8, 32'h43d97031},
  {32'h44b6d6be, 32'h43197d83, 32'hc226edea},
  {32'hc54a53f2, 32'h440120c4, 32'hc3edf7a6},
  {32'h44326b5c, 32'h43ac2f02, 32'h44f1e60e},
  {32'h44992124, 32'h4325ba8a, 32'h43d561b5},
  {32'h44a1c904, 32'hc3b38f3d, 32'hc252f5e0},
  {32'hc51083c9, 32'h4435e138, 32'h43b5f1a1},
  {32'h44228be6, 32'hc395563d, 32'h4375e3db},
  {32'hc573b99b, 32'hc304f0b1, 32'h43271fd9},
  {32'h44a31cfe, 32'hc44fa91e, 32'hc29d46e2},
  {32'h44effd26, 32'hc34568e9, 32'hc30e9b9d},
  {32'h441ffb5d, 32'h4385e991, 32'h44b34f84},
  {32'hc3838fcc, 32'h433b8df9, 32'h439a173d},
  {32'hc0325f20, 32'hc225d716, 32'hc46000f3},
  {32'hc5157f75, 32'h43d5fa2c, 32'h42ea7c6b},
  {32'h439b96ac, 32'hc4c34594, 32'hc372035a},
  {32'h44180efa, 32'h42dd45d4, 32'h43f3824e},
  {32'hc37bf214, 32'h42b1491e, 32'hc4b9890e},
  {32'hc1d80f4c, 32'hc35b80a4, 32'h450e40ef},
  {32'h45480d9e, 32'hc24d74c2, 32'hc30ccb52},
  {32'hc3766840, 32'h4354b709, 32'h442d02a0},
  {32'h4462f894, 32'hc4947247, 32'hc4b13333},
  {32'hc50ebef9, 32'hc3012a2c, 32'hc35baa06},
  {32'h40cf2b80, 32'hc3fa5306, 32'hc54b32b7},
  {32'h43e1d23e, 32'h44be33bf, 32'h441d827d},
  {32'hc49fc458, 32'hc3279832, 32'hc3714f14},
  {32'hc484e8ce, 32'h43902c8b, 32'hc34056e4},
  {32'h4501dab4, 32'hc3e337ab, 32'hc4a6cb90},
  {32'h439f1780, 32'hc23cc284, 32'hc49982c0},
  {32'hc4308464, 32'hc36cd2bf, 32'h45414b81},
  {32'hc2bea0c0, 32'h43d117a7, 32'h43cd2958},
  {32'hc3009066, 32'hc54ae8fa, 32'h43f0a134},
  {32'h4358fb18, 32'h4549f934, 32'hc323e355},
  {32'hc4f6063d, 32'hc22ff6fa, 32'h42dad1c3},
  {32'h450e4df5, 32'h4483df2c, 32'h43438413},
  {32'hc4a22b7a, 32'hc46e12a8, 32'h4406d531},
  {32'h4530e1f4, 32'hc2f0da48, 32'h433837c1},
  {32'hc361e6c2, 32'h43d453cc, 32'h448b4f07},
  {32'h44520d8f, 32'hc3625faa, 32'hc42737cc},
  {32'hc5214c6b, 32'hc269ec52, 32'hc32a04ce},
  {32'h437bbf2d, 32'h441a06b1, 32'h44d51bd3},
  {32'hc44a2d54, 32'hc4c4b570, 32'hc4b779eb},
  {32'h44227d2e, 32'h4213a48b, 32'hc2d5f0a0},
  {32'hc30d87dd, 32'hc46a4f6d, 32'hc46fec2e},
  {32'h43b82718, 32'h449a4796, 32'h44a2051f},
  {32'hc3d9d164, 32'hc41645af, 32'hc3a2826c},
  {32'h44966de0, 32'h4485981d, 32'h44381275},
  {32'hc44079e7, 32'hc493528e, 32'hc4e5817d},
  {32'h4536f348, 32'h43aa0819, 32'hc4082373},
  {32'hc47ca1ba, 32'hc49f1d07, 32'hc3802cba},
  {32'h432d4637, 32'hc38cba40, 32'h44b02646},
  {32'hc33378ac, 32'hc3e085b2, 32'hc44c233f},
  {32'hc39be694, 32'h442b45c3, 32'h451333bc},
  {32'hc425571a, 32'hc4f394b8, 32'hc3ab5d0a},
  {32'hc423f07d, 32'h443d97fb, 32'hc3c8a12c},
  {32'hc40b36fb, 32'h4453d0c6, 32'h437832c0},
  {32'hc2da4229, 32'hc5092160, 32'hc3138b89},
  {32'h44f24d46, 32'h43a9c278, 32'h4334bb70},
  {32'hc3a275e8, 32'hc4b23496, 32'h43e2eedb},
  {32'h44106976, 32'h44fe1754, 32'hc2417332},
  {32'hc4f94420, 32'hc46efdcd, 32'hc38e0726},
  {32'h44995794, 32'h43feafc6, 32'hc3f4ba6a},
  {32'hc4717b80, 32'h43c28083, 32'hc45fa4d2},
  {32'h44b058f4, 32'hc3c964a9, 32'hc3a12534},
  {32'h43bc0ea6, 32'hc3375538, 32'hc4208b09},
  {32'h43b236ea, 32'h44678de2, 32'hc1838484},
  {32'hc457a41a, 32'hc3f68acb, 32'h42787845},
  {32'h45494aec, 32'h42d00493, 32'hc37d94da},
  {32'hc3987dfb, 32'hc51d2597, 32'hc2b1c9cc},
  {32'h44d30662, 32'h441f3e2e, 32'hc3df04bd},
  {32'hc5145edf, 32'hc30c1633, 32'hc383ec6d},
  {32'h4539dff9, 32'hc3bd06de, 32'hc3181805},
  {32'hc48d44d6, 32'hc402e218, 32'hc30c6570},
  {32'h451a9dba, 32'hc3cff7b5, 32'hc4181c88},
  {32'hc3e065f8, 32'hc4bd9bf0, 32'h44258ad6},
  {32'hc3d714b0, 32'h436b5494, 32'hc22c275f},
  {32'hc3289980, 32'hc451dbf4, 32'hc539f933},
  {32'hc49f28b3, 32'hc4bcd1ad, 32'h4409b630},
  {32'h4301ae14, 32'h436ef593, 32'hc3195c59},
  {32'hc46c6dd5, 32'h43d457bf, 32'h44be5c06},
  {32'h43b9c9d0, 32'hc2d4fa64, 32'hc4cae7ae},
  {32'h44187afa, 32'hc4af4e28, 32'h42dbfb09},
  {32'h427f217e, 32'h455554e0, 32'h431a6a57},
  {32'h440b1297, 32'hc4c8dcc5, 32'h43c16bb2},
  {32'h42bfcb98, 32'h45646f1a, 32'h42c03145},
  {32'h44bf18b6, 32'hc4397298, 32'h432e56c5},
  {32'hc39e3ab2, 32'h44d3984c, 32'hc400ea98},
  {32'h4432950a, 32'hc32a4a59, 32'hc34fe659},
  {32'hc485052a, 32'h43e269d1, 32'h441654a6},
  {32'h4534a43d, 32'hc3d9b31b, 32'hc1104638},
  {32'hc50297e2, 32'h428b69d6, 32'hc4065f2a},
  {32'h438bb820, 32'hc4c4b3a0, 32'h43c55cdf},
  {32'hc47ae526, 32'hc3b6f3f4, 32'hc0f627a2},
  {32'hc1b36d60, 32'hc452ec6e, 32'h44f59019},
  {32'hc2861a78, 32'h435c0437, 32'hc507437e},
  {32'hc2c01580, 32'hc424fdf8, 32'hc2a5ccbe},
  {32'hc3bfc3b0, 32'hc3e2430a, 32'hc42e7c0c},
  {32'h43ee11b8, 32'h43e0f972, 32'h4522992a},
  {32'hc3ceb8c0, 32'h42c9e24a, 32'hc41f9d6b},
  {32'h43e4936e, 32'hc480d5b8, 32'h443d0f1d},
  {32'hc548b105, 32'h4469ead2, 32'hc3c6786e},
  {32'hc3683038, 32'hc4b8b09d, 32'h42ff5e60},
  {32'hc4ae5de1, 32'h431333fa, 32'hc496b618},
  {32'h445af922, 32'hc4dab9f0, 32'h4404d688},
  {32'h3fad2f5d, 32'h44e56884, 32'hc3aaab89},
  {32'h4424f5fd, 32'h44371353, 32'h452a8bf9},
  {32'hc47e4f50, 32'hc47514f8, 32'hc4aabac4},
  {32'h441d7250, 32'h436c0a21, 32'h44b94343},
  {32'hc4b94e94, 32'h4330250e, 32'hc41f69b0},
  {32'hc3112f94, 32'h432323ee, 32'h455517a2},
  {32'hc2b3d1dc, 32'h43f32357, 32'hc4339bbb},
  {32'hc3a4c285, 32'h44ed9216, 32'hc32b86d0},
  {32'h43fcefd6, 32'hc2671472, 32'h45027e14},
  {32'hc4175b93, 32'hc3c4b28f, 32'hc4b9ac1c},
  {32'h450d767f, 32'h44212ee4, 32'hc32eca93},
  {32'hc55f16ff, 32'hc38aa07d, 32'hc07863d4},
  {32'h44d12d58, 32'h420e6855, 32'hc1a88cce},
  {32'h41c82e70, 32'h4504a9af, 32'h44c6a36d},
  {32'hc4ba81c0, 32'hc49e2fe6, 32'hc41e3b9a},
  {32'h437bbe68, 32'h4392a583, 32'h430d8daa},
  {32'hc4057ffa, 32'h433cbd65, 32'hc34a67d1},
  {32'hc50328dc, 32'h42b85c7e, 32'hc3e6e81f},
  {32'h4461ce80, 32'hc4a9275b, 32'h43825860},
  {32'hc446f3ae, 32'h422c523a, 32'hc1102afc},
  {32'h44b39b50, 32'hc452d3ca, 32'h442f8c6c},
  {32'hc4e84b34, 32'hc32d25e7, 32'hc3f3e818},
  {32'h44708437, 32'h437cefec, 32'h4459f383},
  {32'hc5004f0e, 32'hc44d8c4c, 32'hc41b4384},
  {32'h453c8cef, 32'hc303559d, 32'h43fc2d2e},
  {32'hc4df2d05, 32'hc29b3753, 32'h43f7f590},
  {32'h44f9d49c, 32'hc2bc6ef1, 32'hc35dc151},
  {32'hc493b81c, 32'hc2494352, 32'h42c2e2a4},
  {32'h4504c682, 32'hc38e8049, 32'hc1bd8ed0},
  {32'hc4d23b9a, 32'h44923635, 32'hc3d9df7a},
  {32'h4451f994, 32'hc50a99d6, 32'h437fbb39},
  {32'hc392a138, 32'h449d28b4, 32'h439baf3d},
  {32'h43e4df82, 32'hc3f7b960, 32'hc48da6f7},
  {32'hc4148ff3, 32'h4412733d, 32'h44d1febb},
  {32'hc2be5688, 32'hc5246155, 32'hc1212ef5},
  {32'h427ed2f4, 32'hc32abb18, 32'hc3e6b4a6},
  {32'hc4a024d7, 32'hc47eddb2, 32'h42c23018},
  {32'hc0290c00, 32'h444c2297, 32'hc44b1aa8},
  {32'hc536c8f8, 32'hc3b13a4a, 32'h43881aed},
  {32'h44530466, 32'hc2b1d25d, 32'h42f04a78},
  {32'h45056f96, 32'h43ee6be7, 32'h4405edb1},
  {32'hc254e780, 32'hc487caa4, 32'h44f082fc},
  {32'h42509996, 32'h4504d962, 32'h43bb2d03},
  {32'hc33bcc40, 32'hc4639e72, 32'h4450810d},
  {32'h452b6020, 32'hc31c29b3, 32'hc34a39f8},
  {32'hc4989e7e, 32'hc49c5b7f, 32'h441f8c0c},
  {32'h441731aa, 32'h43abd90e, 32'h4178caf5},
  {32'h43541353, 32'hc43c6797, 32'hc4257bb6},
  {32'h439b93d8, 32'h4368f8c7, 32'h42aa2f29},
  {32'hc55e301e, 32'hc327eb8f, 32'hc401640e},
  {32'h4393d1e6, 32'hc385da2b, 32'hc3a859b6},
  {32'hc3d9b4b0, 32'hc5828a56, 32'hc3ccd89f},
  {32'h43beeef0, 32'h442ed65d, 32'h4308631c},
  {32'hc448adf2, 32'hc3a100fc, 32'hc29946f4},
  {32'h40ad5000, 32'h4504faf8, 32'hc33fa058},
  {32'hc48f0fe6, 32'hc4bdbfe1, 32'h434b2352},
  {32'h45455723, 32'hc43bba93, 32'hc355f8b5},
  {32'h44283c57, 32'hc40eb8f5, 32'h43338327},
  {32'hc3396108, 32'hc3b8c055, 32'hc3d88a2a},
  {32'hc39e4d57, 32'h42fe48a7, 32'h430bbc58},
  {32'h43ac2b24, 32'hc2d103e3, 32'hc41eb1e4},
  {32'h44260e51, 32'h441ff024, 32'h44f949ed},
  {32'hc48037cb, 32'hc28343fd, 32'hc48613b3},
  {32'h44eaf75a, 32'hc3494866, 32'hc317c26c},
  {32'h436c8ac4, 32'hc335bbe5, 32'hc495e0fc},
  {32'h450fd65e, 32'h42e203d1, 32'hc21a7c6e},
  {32'h43ae0f0d, 32'hc5075204, 32'h43068afa},
  {32'hc3df2c8e, 32'h42ec7f17, 32'h448aa44d},
  {32'hc44987e5, 32'h429a1a6b, 32'hc46bb316},
  {32'hc4e6a353, 32'h436e77fe, 32'hc31b7782},
  {32'hc50a0cfc, 32'hc4351886, 32'h4291e411},
  {32'hc316a222, 32'h43660115, 32'h451ddf37},
  {32'h441d36fa, 32'h434b41fe, 32'h407ae35c},
  {32'h441b07fa, 32'h43a75f2d, 32'h44a40bbe},
  {32'hc35f1408, 32'hc37696d8, 32'hc5779a2b},
  {32'hc2cc6a04, 32'h44d68cd7, 32'hc3949563},
  {32'hc3a6a288, 32'hc584fbb4, 32'hc31967e2},
  {32'h44c1aed2, 32'h44aa66d9, 32'h44167061},
  {32'hc4d474c9, 32'h4384b32e, 32'hc3430c86},
  {32'h44e19bfe, 32'h446f36da, 32'h42f05097},
  {32'hc510d050, 32'hc3cab046, 32'h43d052e6},
  {32'h45625412, 32'h44083d03, 32'h438a6af5},
  {32'hc4420e7c, 32'hc40d08b6, 32'hc3d315db},
  {32'h444fa440, 32'h42d89e31, 32'h441720fd},
  {32'h43c7f828, 32'hc433b140, 32'hc43a31e7},
  {32'h431a500f, 32'hc5131c6e, 32'h44a7ce74},
  {32'h434e1dee, 32'h42b533b8, 32'hc4310be2},
  {32'hc50cb59b, 32'h43e151d8, 32'h43f2ebff},
  {32'h44c395dc, 32'hc44dac0f, 32'hc2e20f40},
  {32'hc55b7df4, 32'hc3a23d4e, 32'h43159f52},
  {32'h454d2312, 32'hc415bde6, 32'h423f8f53},
  {32'hc4ba13a6, 32'h4452edd2, 32'h442bce4a},
  {32'hc491103d, 32'hc35b2d41, 32'hc4529d5d},
  {32'hc4bc789c, 32'hc33a67b6, 32'h4406c20f},
  {32'hc3515ffb, 32'hc4188397, 32'hc494a73b},
  {32'h446f1e42, 32'hc34300ae, 32'h434cc0da},
  {32'hc35ec1c0, 32'hc50db886, 32'hc3a2bdde},
  {32'hc3d6ad94, 32'h4493b43c, 32'hc3d47bcd},
  {32'h43b0f858, 32'hc3044e2c, 32'hc4853b17},
  {32'h42bf1268, 32'h41d99500, 32'h453f8651},
  {32'hc40bd61f, 32'hc2ffc41b, 32'hc51cae01},
  {32'hc547298e, 32'hc2aafdd6, 32'hc3b92629},
  {32'h452dab84, 32'hc48f0007, 32'h4010c6d3},
  {32'hc5001e37, 32'h449e392a, 32'h4395783a},
  {32'hc481a1d8, 32'h431b620b, 32'h43121f8a},
  {32'hbfc77790, 32'h4559dad2, 32'hc3408920},
  {32'h4484f712, 32'hc45ad8ac, 32'hc3062fb8},
  {32'h43565d63, 32'hc3f1d148, 32'h430d4208},
  {32'h457c5c94, 32'h440fc1a9, 32'h444cbc6e},
  {32'hc585c022, 32'hc38d6f62, 32'hc388454a},
  {32'hc43b2097, 32'hc18850b8, 32'hc3f218bb},
  {32'hc4b3c041, 32'h42defa41, 32'h43bf91c4},
  {32'hc49d0ed5, 32'hc3a9dfb0, 32'hc26b8880},
  {32'h44d90ead, 32'h41fbd382, 32'h44bc7b95},
  {32'hc3d95fa4, 32'h43c093cc, 32'h435927ec},
  {32'h43a5386c, 32'hc5201ee4, 32'h430adabb},
  {32'hc43d6128, 32'h440493bb, 32'hc43ae73e},
  {32'hc461bb2a, 32'hc391a08f, 32'h43c83e21},
  {32'hc40865f2, 32'h453a7dda, 32'hc20f193c},
  {32'h450d0dcc, 32'hc3d84e3d, 32'h4345a931},
  {32'h44db47c2, 32'hc3d6113d, 32'hc2b1f175},
  {32'h43ee7620, 32'hc45eb4e5, 32'hc4172644},
  {32'hc43f2d06, 32'h43419a4e, 32'hc48a7d51},
  {32'h437db065, 32'hc38cd93d, 32'hc2e64e37},
  {32'h43455730, 32'hc3001bc4, 32'h45241b58},
  {32'h43ce8d5e, 32'hc439c55a, 32'hc51b037c},
  {32'h44961e81, 32'h435f9f36, 32'h439ffaf8},
  {32'h43c4ca22, 32'hc312fcbb, 32'hc50bfac1},
  {32'hc395b590, 32'h44f3d690, 32'h438d7325},
  {32'h44312a74, 32'h440ff47c, 32'h3f81779f},
  {32'hc569f206, 32'h4010b1c0, 32'h43ee3def},
  {32'h45417922, 32'hc2aa1565, 32'hc40c4d67},
  {32'hc4c436d9, 32'hc29a7b70, 32'h41089b86},
  {32'hc3ce9e48, 32'h441af0da, 32'hc53dc41c},
  {32'hc4017e08, 32'h43efec6b, 32'h44a68591},
  {32'h436282da, 32'hc38eb1d6, 32'hc51245b1},
  {32'hc3690505, 32'h45091541, 32'h4110b754},
  {32'h44e47b8b, 32'hc42de156, 32'hc4ce3cc3},
  {32'h44c1625c, 32'hc3c53560, 32'hc4bc3ee5},
  {32'hc45b525c, 32'h4361dee6, 32'h443004ad},
  {32'h44f831b9, 32'h42423a37, 32'h4335fbb6},
  {32'hc29ab790, 32'hc51bb2a7, 32'hc43300b6},
  {32'h440114c2, 32'h450cf336, 32'h43c0e3eb},
  {32'h4442ca4c, 32'h43577b07, 32'hc393c1e8},
  {32'h4412c890, 32'h45175acd, 32'h431b9f8a},
  {32'hc39e9ecd, 32'hc55bc3f1, 32'hc4035e3a},
  {32'hc17aac3a, 32'h450f44b1, 32'h430827ec},
  {32'hc51cba80, 32'hc363f4ea, 32'h4190defc},
  {32'h43e67233, 32'h43bac54a, 32'h43aaaeb2},
  {32'hc42c6d00, 32'h43a999a3, 32'h4408f04f},
  {32'h428dc362, 32'h448e5ecb, 32'h446d8305},
  {32'h42acd270, 32'hc4bea72e, 32'hc1431b46},
  {32'h449f30d6, 32'h42102ac0, 32'h42987bd2},
  {32'hc3c0e882, 32'hc50bf78a, 32'hc37c0158},
  {32'h4529cca9, 32'h43b9c83d, 32'hc1f19a1f},
  {32'hc4a003b0, 32'hc39fe48d, 32'hc39dce27},
  {32'h42d3c340, 32'h44050925, 32'h44ac8d32},
  {32'hc4676c90, 32'hc4421aad, 32'hc3db1394},
  {32'h44a9910f, 32'h447d8d0e, 32'hc41b4c1f},
  {32'hc3e81af7, 32'hc4bf5307, 32'hc43b46d3},
  {32'h43aa9a87, 32'h44c277a9, 32'hc2ede4b8},
  {32'hc308acf0, 32'hc2e660d4, 32'hc48777d9},
  {32'h43af9223, 32'h44a14fa7, 32'h44876fd3},
  {32'hc4f3fa71, 32'hc3742fae, 32'hc39a8a16},
  {32'hc387511b, 32'h43c8c7a6, 32'hc313a4b2},
  {32'hc4216ddd, 32'h43bd79cd, 32'hc41c5c01},
  {32'hc505999f, 32'hc35d8bb2, 32'h43011339},
  {32'h44496cdb, 32'h44ec59fe, 32'h4454e52f},
  {32'h426504a5, 32'hc48edf01, 32'h43d28e77},
  {32'h446bbcad, 32'h4486f175, 32'hc3b00cce},
  {32'hc3e5bd02, 32'hc4a47d3f, 32'h446e3d1b},
  {32'h446a7b63, 32'h4404e744, 32'h438f3c39},
  {32'hc58f84e2, 32'hc39e66fd, 32'hc21a2ab5},
  {32'hc3f28338, 32'h43f51e05, 32'h43c7c22e},
  {32'h436a5acc, 32'hc4bbebea, 32'hc2f1a3f4},
  {32'h4394ad55, 32'h443ec8f0, 32'hc5134c32},
  {32'hc50dbbd8, 32'hc381e33b, 32'hc25b301e},
  {32'hc412d168, 32'h44207de5, 32'h42b53a87},
  {32'hc3eea969, 32'hc48bd0bf, 32'h44356f3b},
  {32'hc2a1f5b8, 32'h42c5886a, 32'hc508aa13},
  {32'h44c058c8, 32'h42adbee0, 32'h433ad9fc},
  {32'h4426ada0, 32'hc3f1abef, 32'hc490f6f4},
  {32'hc39102b0, 32'h4326280a, 32'hc3eff0e2},
  {32'h446ee586, 32'h4399e7a3, 32'hc466b0bc},
  {32'hc4c5fcda, 32'hc4af84ec, 32'hc3bf1bf9},
  {32'h44e257ee, 32'hc3477a52, 32'h41535afe},
  {32'hc1556f08, 32'hc39895a2, 32'hc4e49d41},
  {32'hc3dc372d, 32'hc4b72840, 32'h4345ab6b},
  {32'hc50200ed, 32'hc2c1eb01, 32'hc1582f00},
  {32'hc5817b22, 32'hc386eee9, 32'h426f64ed},
  {32'h446650db, 32'h439c7b71, 32'hc5057873},
  {32'h44661088, 32'hc493072a, 32'hc40284b0},
  {32'hc42f95f4, 32'h44a79679, 32'h440c22ec},
  {32'h44e354bc, 32'h4412057e, 32'h430bdd1f},
  {32'h419a5140, 32'h452bd687, 32'h4340b2e3},
  {32'h45016bad, 32'hc35734d8, 32'hc335d6c7},
  {32'h43b91c7f, 32'h449e1ab4, 32'hc19c1b81},
  {32'h45434da3, 32'hc3ad2847, 32'hc3519b03},
  {32'hc5766939, 32'hc2cbdaca, 32'hc18f1c94},
  {32'h451b6981, 32'hc311ecf0, 32'h44375652},
  {32'hc4a9e823, 32'h445767ac, 32'hc37793c4},
  {32'h44ac78d4, 32'h43c0b69e, 32'hc4348577},
  {32'hc5124f02, 32'hc3016dd7, 32'hc29e3764},
  {32'h43eda190, 32'hc421f426, 32'h44d49de8},
  {32'hc3777346, 32'h445efed5, 32'hc401fd29},
  {32'h423d4d00, 32'h436f8570, 32'h4425a7f7},
  {32'hc4970ba5, 32'h4412673d, 32'hc3fc52e9},
  {32'h45052065, 32'h434dcd38, 32'h44184e73},
  {32'h43ec275f, 32'h4271d5c9, 32'hc468a96c},
  {32'h45023cb6, 32'hc3ef9acc, 32'h446a9028},
  {32'hc040fc68, 32'h45159324, 32'hc37f003a},
  {32'hc46a581c, 32'h42082024, 32'h4365c647},
  {32'hc19c5300, 32'h4468ddf7, 32'hc3c4e618},
  {32'h44def577, 32'hc4270474, 32'hc2ed33f3},
  {32'h43f916f6, 32'h402fd6c7, 32'h42693f19},
  {32'h44b54670, 32'h43895fd2, 32'h45140c12},
  {32'hc44ac098, 32'hc28b29f4, 32'hc577917a},
  {32'hc299f4f3, 32'hc2ab5502, 32'h44476448},
  {32'h429366f5, 32'hc4247c73, 32'hc514b6c2},
  {32'hc093922e, 32'hc40495a8, 32'h45253305},
  {32'hc449406a, 32'h442cb190, 32'hc130c410},
  {32'h431bd336, 32'h44869dd2, 32'hc38177bf},
  {32'h4526b279, 32'hc4325908, 32'hc409f8b0},
  {32'hc378d44c, 32'h43225550, 32'hc517ba79},
  {32'h440ab32e, 32'hc3408e5b, 32'h40c3a4c3},
  {32'hc3a83bdc, 32'hc26cc22c, 32'hc4b07700},
  {32'h42bf07d7, 32'hc3ab7dda, 32'h448ec31b},
  {32'h446c9c06, 32'h44ab18d7, 32'h44882c94},
  {32'h41df3340, 32'h44960f13, 32'hc4f3960f},
  {32'hc3ebf2a1, 32'h43d8fb75, 32'h42f22c8e},
  {32'hc4052fd8, 32'hc4990368, 32'hc399838b},
  {32'h42461bb0, 32'h44360780, 32'hc46fec05},
  {32'h44134f81, 32'hc35acc83, 32'h452aca0c},
  {32'hc3ad11a8, 32'h4423d4f2, 32'hc3f3d823},
  {32'h4369f690, 32'hc40c435b, 32'h44a43d0e},
  {32'hc3364a98, 32'hc3129798, 32'hc5112ccb},
  {32'h434a6f18, 32'hc43c6a91, 32'h4331387a},
  {32'hc4346a5c, 32'h43cb1c10, 32'hc3a1aabd},
  {32'h44b17170, 32'h420f520e, 32'h4474e203},
  {32'hc5143e9f, 32'hc3a334fd, 32'h438ecdd9},
  {32'h454aa774, 32'hc4057cc6, 32'h440bedae},
  {32'hc49cd22b, 32'h44c615f1, 32'hc34e49ea},
  {32'hc3894951, 32'hc2828da6, 32'h43b16fbd},
  {32'hc5776ec3, 32'h433a5caf, 32'h43d879a3},
  {32'hc057ca80, 32'hc510c80f, 32'h43729936},
  {32'hc4db4a51, 32'hc2c88688, 32'hc387499b},
  {32'hc34bc760, 32'hc4e8e905, 32'hc525ff4c},
  {32'hc3e0f56c, 32'hc16344d3, 32'h44d74fc2},
  {32'hc4136491, 32'hc4023fc2, 32'h4407946a},
  {32'hc3005cc0, 32'hc3254715, 32'hc44270e1},
  {32'hbef35100, 32'hc4959c4a, 32'h431f1043},
  {32'h423a9f16, 32'h4251a31b, 32'hc5662cfc},
  {32'hc456ad7e, 32'hc41d2da9, 32'h4425baa0},
  {32'h4515dc81, 32'hc3b6df13, 32'h43f5a802},
  {32'hc2934f9c, 32'hc4442a05, 32'h41fc401f},
  {32'hc502a7de, 32'hc28a989f, 32'hc3be7b55},
  {32'h44060566, 32'h4480cbcb, 32'hc27c948e},
  {32'hc39bdf2c, 32'hc3fec773, 32'h448b6005},
  {32'hc44abb7c, 32'hc26f628b, 32'hc404b2b6},
  {32'hc5481214, 32'hc29ec3f3, 32'hc1f4cb60},
  {32'h428dedaa, 32'h44b28812, 32'hc487d841},
  {32'hc461bfb1, 32'hc387efad, 32'h41f9a60f},
  {32'h451a5128, 32'h435fb404, 32'hc382f47f},
  {32'hc57902ea, 32'h42f0604f, 32'h42621a72},
  {32'h44e14fe6, 32'h4396ea8a, 32'hc2cef9e7},
  {32'hc4808b2d, 32'hc2002b4f, 32'hc3bc39e6},
  {32'h4327cefb, 32'h4522ff22, 32'h43b6d052},
  {32'hc38ef9a6, 32'hc38030f0, 32'hc2fedc96},
  {32'h44e11646, 32'h44023127, 32'hc3f0e75f},
  {32'hc387d8b0, 32'hc5168058, 32'h43423be7},
  {32'h448b815c, 32'hc384fe67, 32'hc3dba330},
  {32'h44b2d40e, 32'hc40a61e0, 32'hc335551b},
  {32'hc36697ec, 32'h42f13b24, 32'hc4e257b2},
  {32'h450f3af7, 32'h43ede391, 32'h441f2669},
  {32'hc2770116, 32'h41646582, 32'hc448dde3},
  {32'hc26f3a4a, 32'h44bd6e5d, 32'hc41b92e1},
  {32'h42e7032a, 32'hc2bdb997, 32'hc55ecf13},
  {32'hc4c89ec4, 32'hc3746b01, 32'h4225331c},
  {32'hc369b930, 32'hc4083874, 32'hc53ec8f3},
  {32'h44a74359, 32'h42a86444, 32'h449ec2fd},
  {32'h43e168ee, 32'h4489bf1b, 32'hc3908028},
  {32'h44646693, 32'h4358ee2a, 32'hc38b3260},
  {32'h4050cbe0, 32'hc3f61d10, 32'hc483cb71},
  {32'h45170ffc, 32'hc245ce1a, 32'h4326ce24},
  {32'hc2967dc0, 32'hc5375e51, 32'hc35f3dee},
  {32'h4511d19f, 32'h43e4fe2d, 32'hc408b042},
  {32'hc37de066, 32'h42048332, 32'hc3020201},
  {32'h437a9aae, 32'h44d33576, 32'h4481a889},
  {32'hc3da5ce8, 32'hc2fe3d71, 32'hc53a6bfb},
  {32'h440b4c02, 32'h4473be6c, 32'h43919eeb},
  {32'hc4fbbe7c, 32'hc487c69e, 32'h42162f3b},
  {32'h43ecd7f0, 32'h456742a3, 32'hc2e6103f},
  {32'hc52e50f4, 32'hc316d704, 32'hc3577857},
  {32'h425d4540, 32'h44e22a88, 32'hc38d5f24},
  {32'hc4a37330, 32'hc453fad2, 32'hc3485775},
  {32'h44f68f00, 32'h430ebe4d, 32'h4419efee},
  {32'hc56409fd, 32'h432fa85b, 32'hc3eef636},
  {32'h45239ffc, 32'h42e54fb3, 32'hc255f620},
  {32'h420301c3, 32'hc4a1222e, 32'hc3d01e1f},
  {32'hc465d2ce, 32'h43e9cc3c, 32'h439d2433},
  {32'h4241d25e, 32'hc24ed2f0, 32'hc49521cd},
  {32'h43e59340, 32'h44a6ceea, 32'h44cd6d78},
  {32'hc37d2fdc, 32'hc43afb7c, 32'hc4a11a16},
  {32'hc41c514d, 32'h42f6dd2f, 32'h446e273f},
  {32'hc392417c, 32'hc407caf4, 32'hc5370211},
  {32'hc5062a82, 32'h4411d985, 32'h43c7b49e},
  {32'hc2b57f20, 32'hc3f05edb, 32'hc4eb75e4},
  {32'h44197054, 32'h45183e25, 32'h438005a4},
  {32'h449cba4b, 32'h439becde, 32'hc44c3245},
  {32'h4409cf4a, 32'h43a7c873, 32'h43847559},
  {32'h4431b84a, 32'hc3f0799a, 32'hc43be987},
  {32'h43c6b498, 32'hc354e40e, 32'h45343209},
  {32'hc3d6e62e, 32'hc46c4769, 32'hc3938173},
  {32'hc4283318, 32'h445e2ab5, 32'h44a59a42},
  {32'h441749ff, 32'h44245e31, 32'hc4693c50},
  {32'h442b5ac9, 32'h43329efc, 32'h43955a64},
  {32'hc3637806, 32'hc4f54673, 32'hc46bd828},
  {32'hc53348f7, 32'h443c6b2f, 32'h42dfe629},
  {32'h4564e5b4, 32'h43b13b5e, 32'hc33ec6f6},
  {32'hc4af02ac, 32'h44e0564d, 32'hc3886788},
  {32'hc3284f9a, 32'hc51349fa, 32'h428c26f4},
  {32'h44de5d7a, 32'h435d9173, 32'hc3522ddc},
  {32'h44b6d3ae, 32'h432b7216, 32'h42fb32bc},
  {32'hc432f9be, 32'hc31add32, 32'h42ad5e56},
  {32'h4475a4c6, 32'hc3c8f583, 32'hc36fe37b},
  {32'h451424ce, 32'h41c89f8d, 32'hc3077a71},
  {32'hc49055f3, 32'hc338d236, 32'hc2341163},
  {32'h4414be60, 32'hc342340a, 32'h456347b2},
  {32'h4410f1de, 32'h42796013, 32'hc32ebd54},
  {32'h43d4e984, 32'hc4a64019, 32'hc329af97},
  {32'hc40149c0, 32'h45187a1f, 32'h43f58d6b},
  {32'h450b981e, 32'h43b32572, 32'hc3245db3},
  {32'hc39ac60c, 32'h45418dee, 32'hc35c2cba},
  {32'h441df074, 32'hc4cc618a, 32'hc3329651},
  {32'h4430ee3b, 32'h438656ed, 32'h43cbca98},
  {32'h44011dc5, 32'h44827552, 32'hc4aaa267},
  {32'hc51536b9, 32'h443cdeca, 32'hc394d0c3},
  {32'hc44cefaa, 32'hc3b72cfd, 32'h42aae045},
  {32'h4386e895, 32'hc3d253c5, 32'h4542e91e},
  {32'h4423d1c0, 32'hc4a458e9, 32'hc3866057},
  {32'h44b53a6f, 32'h4389433e, 32'hc3b63664},
  {32'hc2ae86a0, 32'hc49a0ed7, 32'hc41c5847},
  {32'hc482a4da, 32'h422d1527, 32'h44b45812},
  {32'h45366367, 32'h429eff31, 32'h437539c6},
  {32'hc54d4b7a, 32'h4331c0ef, 32'h440021a8},
  {32'h4523cce7, 32'hc3c35e5b, 32'hc456afd1},
  {32'hc30fecec, 32'h448195a2, 32'h446fa1fc},
  {32'h4521ae5a, 32'hc381cdfb, 32'hc3d0ac05},
  {32'hc512138c, 32'hc2670c22, 32'h43dd938a},
  {32'h4398a5a0, 32'h43f2970e, 32'hc3cd076a},
  {32'h431f8f60, 32'h442461de, 32'h45048ab8},
  {32'h44c22667, 32'hc42977d3, 32'hc4ad0f31},
  {32'h450eb76c, 32'hc3ac3a43, 32'hc4922dc6},
  {32'hc43974a3, 32'h44054a32, 32'h451e8461},
  {32'h44074acb, 32'h44680579, 32'hc4a2b1cc},
  {32'hc5252de6, 32'hc4192d9c, 32'hc2233166},
  {32'h449928e2, 32'h43b47cf4, 32'h423d6675},
  {32'h44b0e938, 32'hc2f8f09c, 32'hc41fc9f3},
  {32'h452418ac, 32'h446cb642, 32'h43af872e},
  {32'hc453205e, 32'hc437df50, 32'h44053943},
  {32'h44a02c96, 32'h439c427c, 32'h4415c529},
  {32'hc47afd14, 32'h43abcf2a, 32'h44b87365},
  {32'h44a7e7a7, 32'hc2bd0e56, 32'hc4316633},
  {32'hc4b51c9f, 32'h438882d5, 32'h43fdaba5},
  {32'h43e0c762, 32'h4491163a, 32'h44090351},
  {32'hc49569f6, 32'hc42147fb, 32'hc44d589c},
  {32'hc4ea447a, 32'h43b70183, 32'h43d638f6},
  {32'hc27b1ac0, 32'hc3ebfdb9, 32'hc4394138},
  {32'h43c40203, 32'h44d38ac2, 32'h4466d469},
  {32'h42820228, 32'hc35172be, 32'hc47f2be3},
  {32'h42697ce0, 32'hc3221a27, 32'h42213ee1},
  {32'hc4d3306b, 32'h4353bcfa, 32'hc284f9d8},
  {32'hc3a92f6e, 32'hc15fb991, 32'h42f28123},
  {32'hc50bf303, 32'h4302eee2, 32'hc41f12e4},
  {32'h4536e2f4, 32'h43cdb161, 32'h437f985d},
  {32'hc39529fb, 32'hc3fa0c58, 32'hc3da874f},
  {32'h446fb850, 32'h44a15033, 32'h43b33a8a},
  {32'h42c84ac8, 32'hc4e08ddd, 32'hc36d3d95},
  {32'h4532cb59, 32'hc3abca59, 32'h43939f6b},
  {32'h43979307, 32'hc381e422, 32'hc3cd9bfc},
  {32'hc44cb568, 32'hc4d1fb3f, 32'h431cec21},
  {32'h4435d6d4, 32'h44b8e358, 32'h43e5c98b},
  {32'hc46293d5, 32'h43462547, 32'hc33f9db4},
  {32'h4527e72c, 32'h4367ed1c, 32'hc3633d17},
  {32'hc40562dc, 32'hc53e69bb, 32'h4382a025},
  {32'h43a33842, 32'h441485a1, 32'h42f8a6c4},
  {32'hc57bc948, 32'hc1bbf3f9, 32'h4352be88},
  {32'h43b7d4c3, 32'h44773420, 32'h4482d0b6},
  {32'hc467636a, 32'hc42100c1, 32'h43fd9ffe},
  {32'h4411769d, 32'h44cfcfe9, 32'h4375790a},
  {32'hc44340d4, 32'hc34432e4, 32'hc36d2d74},
  {32'hc263a006, 32'h4476334f, 32'h4298e3bc},
  {32'hc480ecd9, 32'hc3cacb2a, 32'h43045430},
  {32'h44ff5522, 32'h43f9c9c6, 32'h421f67df},
  {32'hc481cd97, 32'hc3be83ce, 32'h418a5ad9},
  {32'h42e9ba10, 32'h43d3b20e, 32'hc4280135},
  {32'hc543736c, 32'hc2ca64e7, 32'h435cabc5},
  {32'h45502a8d, 32'hc3fa37b9, 32'hc35d88c3},
  {32'hc50ea2d6, 32'hc4174582, 32'hc357864e},
  {32'h44556dec, 32'h423880b6, 32'h3fe9bfa3},
  {32'h44882e73, 32'h44a0e925, 32'hc3dd4454},
  {32'hc4ada463, 32'hc451098e, 32'hc399fdfa},
  {32'hc488f9a9, 32'hc208aaa7, 32'hc336872a},
  {32'hc21f0034, 32'h43e27260, 32'h45527c20},
  {32'h4513f590, 32'hc39c05ba, 32'hc4a0c156},
  {32'h4488af52, 32'hc3cc7dcf, 32'hc46ce054},
  {32'hc45724a4, 32'h4409cdf6, 32'h44660255},
  {32'h44cfd578, 32'hc3472560, 32'h431f3fc7},
  {32'hc5454ad2, 32'h4306c8c7, 32'h442cbe76},
  {32'h453acade, 32'hc33edfcd, 32'h432fef8e},
  {32'h4479e06a, 32'h42f4798a, 32'hc3454db8},
  {32'h44b648ff, 32'h44130d54, 32'hc2b6afda},
  {32'hc4bd686f, 32'h42ad8ed9, 32'h43b77b26},
  {32'hc4bbd311, 32'hc3be61a4, 32'hc2a5f526},
  {32'h43b88ac9, 32'h451ad7b5, 32'h43d5fcf3},
  {32'hc30bfbb6, 32'hc376eef2, 32'hc408799c},
  {32'hc421fe4b, 32'h42b404d7, 32'hc4529b74},
  {32'hc2942504, 32'hc4c741b4, 32'h43957177},
  {32'hc3abe6cf, 32'h4512158d, 32'hc40e1850},
  {32'h437725b4, 32'h428ed47f, 32'h43c7cfc4},
  {32'hc50beddd, 32'hc30ef56d, 32'hc4117fdc},
  {32'h44bdb53c, 32'h43d4514d, 32'hc1f872d4},
  {32'h444b52b8, 32'hc3328601, 32'hc48401be},
  {32'h44604e1f, 32'hc4735822, 32'hc2702305},
  {32'hc515fcea, 32'h440a6200, 32'hc439b677},
  {32'h4545bc10, 32'hc266a038, 32'hc2ae2d90},
  {32'hc3b783f0, 32'h43b68490, 32'hc3f0bcec},
  {32'h45475eb4, 32'h43c7a4b0, 32'hc3fa9a35},
  {32'h431e413e, 32'h44091dea, 32'hc21cbfc6},
  {32'h441ce620, 32'h443a042e, 32'h45435599},
  {32'hc4c72446, 32'hc3b3c9da, 32'hc4d4f14e},
  {32'h449c93d9, 32'hc2709954, 32'h43ba34d2},
  {32'h41f6cc18, 32'hc4852980, 32'hc4ff9c0b},
  {32'hc3068324, 32'h4342d265, 32'h44d3a85b},
  {32'h44da8a5c, 32'hc309348e, 32'hc4296069},
  {32'h43ea59ee, 32'hc34cefab, 32'hc499eea8},
  {32'h453ed406, 32'hc3b3284a, 32'hc38e32d1},
  {32'hc425c290, 32'h43c2c557, 32'hc4263aea},
  {32'hc3e861fe, 32'h4407f574, 32'hc28f7e43},
  {32'hc429a51a, 32'h4514a8f8, 32'hc2d8e396},
  {32'h44307712, 32'hc3950360, 32'h44dcaba7},
  {32'h452750be, 32'h438dfb6e, 32'h4436bdf2},
  {32'hc3eda5a4, 32'h44b066c7, 32'hc46e455c},
  {32'h44e8460c, 32'hc3943ecb, 32'h43719941},
  {32'h44243f33, 32'h43715dfa, 32'h4407c6f8},
  {32'hc3b311c3, 32'h44bd4665, 32'hc3b97c58},
  {32'h43d84f36, 32'hc3cd3b06, 32'h44cf8e02},
  {32'h4351a5da, 32'h4469c3e9, 32'hc4763e47},
  {32'hc3a019f0, 32'hc30c673d, 32'h44f183d3},
  {32'hc4ba4b28, 32'h4212c096, 32'hc31337a4},
  {32'h44c75915, 32'hc42804b6, 32'hc2a4b676},
  {32'hc4628141, 32'hc485bffd, 32'hc4226e03},
  {32'h449d74ae, 32'h442a39e7, 32'hc3a9bc1d},
  {32'hc552fcf9, 32'hc370da90, 32'h41bb3e30},
  {32'h449dee79, 32'hc491798f, 32'hc40896fe},
  {32'hc4f08d79, 32'hc3eb4784, 32'h432422f3},
  {32'hc3f544b4, 32'hc3f3b4ed, 32'h43f4bd5f},
  {32'hc497bc62, 32'h44dc17c3, 32'h4362600a},
  {32'h455c7287, 32'hc41ac0df, 32'hc29934ea},
  {32'h448dbf4d, 32'h43483c83, 32'h434bf6c1},
  {32'h4381fa7c, 32'h43956eca, 32'hc4be0a42},
  {32'hc470e7e4, 32'hc32d20c7, 32'h442d611b},
  {32'hc44f755a, 32'h4397c156, 32'h44bb9c1d},
  {32'hc294d128, 32'h44a7f4e2, 32'hc44a8c54},
  {32'hc50928b9, 32'h435205a7, 32'hc359271a},
  {32'hc40d6522, 32'h439b4d3a, 32'hc46a4c1b},
  {32'h4300779e, 32'hc428a55d, 32'h44e67464},
  {32'hc4b9d63f, 32'h422b5154, 32'hc397b432},
  {32'h44e4a510, 32'hc3fd5cf9, 32'h42b42b9a},
  {32'hc3943981, 32'h4284c772, 32'hc300b907},
  {32'h430ce892, 32'hc473e358, 32'hc40ad360},
  {32'hc491c856, 32'hc43b9ef3, 32'h4490fcdf},
  {32'h449ca7c7, 32'h43b134c2, 32'hc45ec8a0},
  {32'hc4cda964, 32'hc465b9fb, 32'h443357f6},
  {32'h44a4e7f2, 32'h42b77a5a, 32'hc391fa14},
  {32'hc4ae97d6, 32'hc32817a7, 32'hc30d4b92},
  {32'h451263ab, 32'h4377bd3e, 32'hc349b2ac},
  {32'hc58fed3f, 32'hc2ce4373, 32'h435868ca},
  {32'hc38f2aca, 32'h401d8af6, 32'h42c1a8eb},
  {32'hc4404210, 32'hc4e4afe8, 32'h43584288},
  {32'h42f7d5e7, 32'h455db902, 32'h4350c29b},
  {32'h42a08a54, 32'hc4e1b128, 32'h43abc5d7},
  {32'h44a9c499, 32'h44d08dec, 32'hc3ab6d31},
  {32'hc3c24569, 32'hc4e9a40f, 32'h4381977a},
  {32'hc3cdf41c, 32'h442d7f24, 32'h41695249},
  {32'h41b70c94, 32'h447bed02, 32'hc280b82d},
  {32'h4454ec55, 32'h446e3e20, 32'hc4ee9e1a},
  {32'h4438415e, 32'h44ffd89a, 32'h4410c938},
  {32'h43890c9c, 32'h42b78b23, 32'hc4d60e87},
  {32'h43bb0577, 32'h4505473f, 32'hc240f560},
  {32'hc4361d45, 32'hc380e870, 32'hc496b428},
  {32'h42eb5c50, 32'h43cb6f93, 32'h43ebad83},
  {32'hc44028bc, 32'hc42a3f58, 32'hc4e46054},
  {32'h43bdb9a0, 32'h44e47e97, 32'h448b5fe7},
  {32'h4460525c, 32'hc38bd9ba, 32'h42f9a92e},
  {32'h44a99032, 32'h4389c276, 32'h41eb26ad},
  {32'hc40e0679, 32'h44e441ed, 32'hc4dfb2b8},
  {32'h45209fac, 32'h43271eee, 32'h40fb288c},
  {32'hc46d9c8e, 32'hc48edfb0, 32'hc3608154},
  {32'h449b8f68, 32'h448dda85, 32'h435be141},
  {32'h44ae4b8e, 32'h436bad2a, 32'hc3228315},
  {32'hc3122856, 32'h44048c00, 32'h451fed18},
  {32'hc48e7777, 32'h43191b03, 32'hc2f627f8},
  {32'h43bbe8b4, 32'h4385f17d, 32'h43c66d21},
  {32'hc51f711e, 32'hc1eee0fe, 32'hc39ad743},
  {32'h456181af, 32'h440e008b, 32'hc3f37cee},
  {32'hc49fa913, 32'h43bcfe90, 32'h43c8d2b8},
  {32'h4549f6ca, 32'h43e8d62a, 32'h41d6f5b4},
  {32'hc18bdde0, 32'hc48785a5, 32'hc396d465},
  {32'h453fa3ec, 32'h41611abb, 32'h4388ed1d},
  {32'hc4591246, 32'hc3c58a4b, 32'hc2f6d486},
  {32'h45758a33, 32'h41f46d16, 32'hc1d7dc3c},
  {32'h4117b8c0, 32'h44c67e91, 32'hc4f3ceb4},
  {32'hc2e55200, 32'h449985c6, 32'h444f7333},
  {32'h43bf7972, 32'hc423f796, 32'hc3e2367a},
  {32'hc12f71a8, 32'h443495da, 32'h4381edbd},
  {32'h430e7448, 32'hc476e2a2, 32'hc4e05171},
  {32'hc495ccbd, 32'hc35f6952, 32'h43243a5b},
  {32'h4486fc4d, 32'hc469bfd0, 32'hc474f38a},
  {32'hc5541759, 32'h42c9442a, 32'h43f866f9},
  {32'hc30da927, 32'hc4355bfb, 32'hc2cdff2c},
  {32'h43bfe3c0, 32'hc499bbac, 32'h45215441},
  {32'hc44093d9, 32'hc4a1a460, 32'hc31ee947},
  {32'hc50a6d36, 32'h435b2647, 32'hc2560453},
  {32'h43dfda22, 32'hc3f2ade6, 32'h43a7e520},
  {32'hc4b7e7dd, 32'h4428c202, 32'h432199e7},
  {32'h44fa1e29, 32'hc28c4ae8, 32'hc385165a},
  {32'hc5092ce4, 32'h43105d69, 32'h43d8ffdf},
  {32'h43b820a0, 32'hc31cd2aa, 32'hc5101218},
  {32'h43150e4b, 32'h44b40d63, 32'h4447b97e},
  {32'h44b90544, 32'hc493695e, 32'hc4041dd6},
  {32'hc32bf1c8, 32'h44429907, 32'h4414563f},
  {32'h45503335, 32'h42db7080, 32'h43e7657e},
  {32'hc4cd5287, 32'h44eca0fd, 32'h440e6efa},
  {32'h44ad354d, 32'hc4aca7ee, 32'h435a6cfd},
  {32'hc2e15352, 32'h44b021aa, 32'hc38918ae},
  {32'h451da967, 32'h43f24821, 32'hc30bbfcc},
  {32'hc55b93c3, 32'hc3e7d84c, 32'hc334ac06},
  {32'h447b1fec, 32'h425e486a, 32'hc3cc4100},
  {32'h453407c8, 32'h42dbd29c, 32'hc3254814},
  {32'hc5568820, 32'h42a0e100, 32'hc2de5f67},
  {32'hc2ad5680, 32'hc2bfd9a7, 32'h42fff27e},
  {32'h448f8f51, 32'h42d291a8, 32'h43dfc733},
  {32'h42b91660, 32'hc4b7cd8b, 32'h43971fd3},
  {32'hc47de601, 32'h4473ca06, 32'hc296adc1},
  {32'hc3a58fda, 32'hc4918bde, 32'hc2b20da4},
  {32'hc10f77b0, 32'h458aa9fb, 32'h4229e7c7},
  {32'h453012ba, 32'hc2980335, 32'h43e0e7ca},
  {32'hc51220fc, 32'hc3d1f6ed, 32'h432afcad},
  {32'h44c31a72, 32'hc382d214, 32'h43f68c9f},
  {32'hc41ed29a, 32'h429a372a, 32'hc541a5f7},
  {32'h42bd76c0, 32'hc3b38768, 32'hc43a59b8},
  {32'h42df4c0e, 32'h44806dc3, 32'h44f095d9},
  {32'h44202b64, 32'hc4430c54, 32'hc3f2b56f},
  {32'hc50e8f20, 32'hc2feb190, 32'hc363a8d8},
  {32'hc1d13f08, 32'h43775cdc, 32'hc556b764},
  {32'hc53f9a48, 32'hc20efdf1, 32'h43a0e10c},
  {32'h4544884e, 32'hc44b6146, 32'h43884c1e},
  {32'hc4b81696, 32'hc4334c7e, 32'h4400094f},
  {32'h449e9de4, 32'h4397c393, 32'hc4a12766},
  {32'h43dd89b6, 32'h43d0a6b7, 32'h44ba1542},
  {32'h4440fee8, 32'hc308a601, 32'h43243b26},
  {32'hc4866bae, 32'h448aabb1, 32'h435cb8d9},
  {32'hc0eaf0c0, 32'hc307a99a, 32'hc4a3984b},
  {32'hc449dcf2, 32'h451151c4, 32'h43dc6ed6},
  {32'h447ca685, 32'hc4992a4c, 32'hc399121e},
  {32'h453275c4, 32'h42e6289a, 32'hc3f5222a},
  {32'hc54fcc61, 32'h419ad162, 32'h4327a05e},
  {32'h446dd44e, 32'h43490875, 32'h44475122},
  {32'hc510964b, 32'hc47fec09, 32'hc401854c},
  {32'h4509abc1, 32'h428a5eed, 32'hc3e22ca3},
  {32'hc318c6c7, 32'hc48c9ac1, 32'h4390e646},
  {32'h44c9ebc0, 32'h449c9fd6, 32'hc3a11e74},
  {32'hc51d83b2, 32'hc46580bc, 32'h43a4872e},
  {32'h44d1695e, 32'hc28c6b5b, 32'h43811e18},
  {32'hc3fc7a40, 32'hc2696696, 32'h44ba3e6c},
  {32'h443aa07c, 32'hc295f02a, 32'hc4e84de0},
  {32'hc29754c4, 32'hc2e0f40f, 32'h44c99933},
  {32'h43855fa0, 32'h44cbf86f, 32'h44402485},
  {32'hc432fe34, 32'hc3a3d00e, 32'hc447389c},
  {32'h45025a1d, 32'hc327d26c, 32'hc341ca7e},
  {32'hc50d3695, 32'hc4223b5b, 32'h434809c9},
  {32'hc3a69fd4, 32'h43d2f288, 32'h44cbcc1e},
  {32'hc43546e2, 32'hc1869dd1, 32'h42f1023b},
  {32'hc2d653f1, 32'hc36a16bb, 32'h44961fa2},
  {32'hc50d83c8, 32'h436d8695, 32'h42f23399},
  {32'hc4802c84, 32'h41416176, 32'hc36679e5},
  {32'hc30f7e4f, 32'hc539e004, 32'hc27186c2},
  {32'h43c0e896, 32'h44f98c73, 32'hc282d3cf},
  {32'hc532220b, 32'hc31b477b, 32'hc2a6c55f},
  {32'h4367e684, 32'h44e3ccc4, 32'h445b8659},
  {32'hc4c46cb1, 32'hc488370d, 32'hc3996ae2},
  {32'hc19c3b30, 32'h44dca6cf, 32'h437398c1},
  {32'h44e0d84a, 32'hc46e5327, 32'h42f81a88},
  {32'hc431b138, 32'hc4c8c113, 32'hc2dea04a},
  {32'h43714fd5, 32'h449c9768, 32'h440c817a},
  {32'hc3ee142a, 32'h43aac781, 32'hc38025f5},
  {32'h452a455a, 32'h43caf875, 32'hc3727e6a},
  {32'hc4b1d43d, 32'hc4b77269, 32'h42f455a5},
  {32'h44340d11, 32'h43b08420, 32'h43c35208},
  {32'hc42f0707, 32'hc45a478a, 32'hc43c9258},
  {32'h453ce707, 32'h43b44ddf, 32'hc31e9da0},
  {32'hc3c265d1, 32'hc427ee2d, 32'h440957af},
  {32'h433f0d12, 32'hc3b0129d, 32'h44791bb0},
  {32'hc491ce82, 32'hc40d88d9, 32'hc3bd6c0c},
  {32'hc394589a, 32'h44231d32, 32'hc248ab8c},
  {32'hc45235d8, 32'hc37af670, 32'h447cf83a},
  {32'h428f9a70, 32'h4221372b, 32'hc4cfb063},
  {32'h44c9eb94, 32'hc34bc4fa, 32'h43332229},
  {32'h44cee2b7, 32'h4410ac0a, 32'hc42c6756},
  {32'hc4ff99af, 32'h434f292a, 32'h44146c67},
  {32'h44624780, 32'h439e9bbd, 32'h425c2aa2},
  {32'hc465f501, 32'hc45d5eb5, 32'h440f890d},
  {32'hc2e1e0bc, 32'hc2c87496, 32'hc2549f07},
  {32'h4383dc60, 32'hc3538412, 32'hc49ba7ab},
  {32'hc4f6caa2, 32'hc4759695, 32'h430552e9},
  {32'hc4c864f2, 32'hc20fde2b, 32'hc38fb006},
  {32'hc52d767c, 32'hc3a700e3, 32'hc38ee7ec},
  {32'h44c8807e, 32'hc4173750, 32'hc4aec8ed},
  {32'h442c3dae, 32'h43ee42eb, 32'hc4dfdc3e},
  {32'hc4c792d4, 32'h444a2cbc, 32'h43a321a3},
  {32'h452b3ac8, 32'h441b0e95, 32'h43fe43d5},
  {32'hc489b7d6, 32'h4508d6ee, 32'hc31138d6},
  {32'hc432b52f, 32'hc5185477, 32'h43fb627a},
  {32'h444b0131, 32'h4479afdd, 32'h43c23608},
  {32'h4516fb18, 32'h431a91f9, 32'hc1fe692a},
  {32'hc58f71a7, 32'h42380e44, 32'hc358b506},
  {32'hc48f78be, 32'hc3198d19, 32'h43edf033},
  {32'hc506f5d9, 32'h4397f9ce, 32'h4307403a},
  {32'h44c6dff3, 32'h42d492a6, 32'hc29b1ed3},
  {32'hc3a2d2b2, 32'hc32af5bd, 32'h437d80a5},
  {32'h448dcec6, 32'h435f34c0, 32'h447c3c3b},
  {32'hc4ddf368, 32'h44071846, 32'hc401d2c2},
  {32'hc4e3bdcf, 32'h43dbbf8e, 32'h440cd0e0},
  {32'hc41278da, 32'hc350e808, 32'hc4c3ceca},
  {32'h4499ae64, 32'hc4b070b4, 32'hc45ecaac},
  {32'h436392f2, 32'hc3f4e5c7, 32'hc49ec623},
  {32'h43e093e2, 32'hc4d2fc78, 32'h431c7df2},
  {32'hc4b00ab2, 32'h4454bc2b, 32'hc3dd5ee1},
  {32'h456349b7, 32'h43cef14a, 32'hc3592c4f},
  {32'hc4d85dbb, 32'h42654c8e, 32'hc4520d20},
  {32'h4491a501, 32'hc47ca8a2, 32'hc3210c9b},
  {32'h4381fbb7, 32'h44d5bad1, 32'hbf245ae8},
  {32'h444da0ef, 32'h434e3c4c, 32'h44b6182a},
  {32'hc4bb80d6, 32'hc2ddea0b, 32'hc51ca6dd},
  {32'h452e383a, 32'hc37d0f6c, 32'hc40191be},
  {32'hc43f86d4, 32'hc2d70eda, 32'hc4b1e9be},
  {32'h43831386, 32'h4421b798, 32'h450d0eb1},
  {32'h42b8df73, 32'h437ae14f, 32'h42445e9e},
  {32'hc489824b, 32'h448bbd58, 32'hc36de877},
  {32'h440a81ce, 32'h42f7d11e, 32'h45113311},
  {32'hc3b1f1c0, 32'h44d3ab48, 32'hc42f0939},
  {32'hc423957a, 32'hc416e1fe, 32'h431bfaca},
  {32'hc36aed38, 32'h440a1c0e, 32'hc50bd1b8},
  {32'h4303c61a, 32'hc541691e, 32'h4288d8a6},
  {32'hc43d7ef8, 32'h434cc440, 32'h454e8eec},
  {32'hc3818fcc, 32'h44bc5b52, 32'hc4c7f938},
  {32'h434b7c5b, 32'hc44070d4, 32'h43690d48},
  {32'h4523764c, 32'h4381279c, 32'hc361bbc2},
  {32'hc458554e, 32'h430f40c5, 32'hc49b6746},
  {32'hc4253a3c, 32'hc425200c, 32'h44aae4c9},
  {32'h44c4434c, 32'h42ab9599, 32'h439a3250},
  {32'h43fab530, 32'hc2298e3f, 32'h44f569c2},
  {32'hc4bdad75, 32'hc2094ffe, 32'hc45dabe7},
  {32'h44406acd, 32'hc4101ba0, 32'h435f50f6},
  {32'hc5855f53, 32'hc3b241c9, 32'hc32e0be7},
  {32'h44889f24, 32'h44857fe4, 32'h43925da7},
  {32'hc529e6fd, 32'hc3e4e59b, 32'hc363c84d},
  {32'h44cdebaf, 32'hc4a850db, 32'h43b76aee},
  {32'hc4c4358f, 32'h44391ddf, 32'h434efe9a},
  {32'hc48184e6, 32'h42cc605c, 32'h424d5373},
  {32'hc3b28606, 32'h45491275, 32'h4240b0c9},
  {32'h446f5cb4, 32'hc4ed73c3, 32'hc35d95ad},
  {32'h4507ba9b, 32'h418692c6, 32'h4397f984},
  {32'hc39abf7c, 32'hc4cf33ce, 32'hc50574fb},
  {32'hc313a8a6, 32'h444aff2f, 32'h44fc5a2f},
  {32'hc40a598d, 32'h42bcbe7c, 32'h44c93f47},
  {32'h4494b766, 32'h43326142, 32'hc353b19c},
  {32'h4383a986, 32'h42e26a16, 32'h448b6b9d},
  {32'h40743858, 32'hc324fc33, 32'hc55a2bf2},
  {32'hc2a85058, 32'hc4368f25, 32'h448618d3},
  {32'hc4a39aa2, 32'h43ed1545, 32'hc3b0b3dd},
  {32'hc3dee299, 32'hc492bb04, 32'h413bd92f},
  {32'hc3e7b664, 32'hc47339fb, 32'h44e58824},
  {32'h44285cf4, 32'h44a64ca3, 32'hc4128ec0},
  {32'hc39364f4, 32'hc4b0d3a4, 32'h4356d3a3},
  {32'h4518bd0d, 32'hc351fb18, 32'h42aec617},
  {32'hc4583cee, 32'hc44a5cc3, 32'h443a6319},
  {32'hc3aa4134, 32'h443a262b, 32'hc414f49b},
  {32'hc44a27ea, 32'hc41a238c, 32'h43afdc07},
  {32'h4532e2c9, 32'hc4114198, 32'hc2bd0c5e},
  {32'hc50b0e78, 32'hc3536135, 32'hc3337f77},
  {32'h45036cf4, 32'h4006189a, 32'hc40940f0},
  {32'hc4180278, 32'hc4898b6d, 32'hc139706a},
  {32'h4562c8b9, 32'hc41ccaa4, 32'hc266f7be},
  {32'h43ff2ce3, 32'hc47a082a, 32'h4283d736},
  {32'hc3b6f6a8, 32'h44cbc22c, 32'hc40d1da4},
  {32'hc548731a, 32'h42a28078, 32'h4385a5ae},
  {32'h42a28644, 32'h441d2d97, 32'h42f831d5},
  {32'hc472c516, 32'h4352a802, 32'hc2e9119a},
  {32'hc007d740, 32'hc47af97f, 32'hc3e11c30},
  {32'h4501fa5b, 32'h43b5c229, 32'h435abe35},
  {32'hc4b60ed4, 32'h440adce5, 32'hc33f5e69},
  {32'h45573174, 32'h41c9e7f9, 32'h43e46ed2},
  {32'h43b01b2f, 32'hc50ccaa8, 32'hc47d221a},
  {32'h4406d03f, 32'h42e9ccf6, 32'hc2df9593},
  {32'hc51dd52d, 32'h41daf78a, 32'hc3a5b1e0},
  {32'h454ca75c, 32'h43a3a419, 32'h439b69e1},
  {32'h441ce1da, 32'h4451a642, 32'hc30d9c20},
  {32'hc39baaf3, 32'h43f139fb, 32'h4477d4eb},
  {32'hc3c5e7b1, 32'h44a0dcbe, 32'hc5058712},
  {32'hc34ab3aa, 32'h42fc363a, 32'h4421793f},
  {32'hc34509a2, 32'hc38f882d, 32'hc503d275},
  {32'h440bfa60, 32'h42d68959, 32'h44890bea},
  {32'h447f8c26, 32'hc48b6a4c, 32'hc3fd41bc},
  {32'h43799a04, 32'h44b3f33f, 32'h4482c477},
  {32'hc28e70d8, 32'hc4f701dc, 32'hc4a9a503},
  {32'h452dfd61, 32'hc35c0d0c, 32'h4483ebd1},
  {32'hc2131960, 32'hc542424a, 32'hc3c29cb0},
  {32'h4568eb90, 32'h43a407a2, 32'hc3f11cd9},
  {32'hc54049d8, 32'h43953c8a, 32'h4266df32},
  {32'h43897991, 32'h4518e74f, 32'h4425c544},
  {32'hc4a8656f, 32'hc42dbd0f, 32'h43d3b48b},
  {32'h451acb09, 32'h4356f1a7, 32'h4386bbd7},
  {32'hc4c7ef6f, 32'hc3f2d4e4, 32'h43117051},
  {32'h4363eacc, 32'h438b4fa1, 32'hc3ea9f0d},
  {32'h43cc295b, 32'hc4d44b23, 32'hc48be805},
  {32'h42b33666, 32'h449f6053, 32'hc492b6d5},
  {32'hc45b2886, 32'h4460d448, 32'h440b7c4c},
  {32'h44043b78, 32'hc41f6cdc, 32'hc434e64f},
  {32'hc2b646a0, 32'h44653140, 32'hc1406ac1},
  {32'h44040e78, 32'hc49e1c06, 32'hc4d03666},
  {32'hc40380db, 32'h4509fd03, 32'h44bc8356},
  {32'hc409e87a, 32'hc2b1b36f, 32'h43ae4882},
  {32'h42b358cc, 32'hc3346d53, 32'h44a57cdf},
  {32'hc30fb6d4, 32'h44b056a2, 32'hc50fae30},
  {32'h442caf49, 32'h44aba48f, 32'h43bdaf51},
  {32'hc39c415d, 32'hc3a564af, 32'hc4e30ddd},
  {32'h436a89ec, 32'hc311ea9d, 32'h43a7988a},
  {32'h448065fd, 32'h42e957b2, 32'hc3b5571b},
  {32'hc3cd08ec, 32'h44971cf3, 32'h44ca0954},
  {32'h44c09216, 32'h43119f1c, 32'hc45a8a9b},
  {32'h442ed4d8, 32'h43a1af36, 32'h439f8867},
  {32'h44afa23a, 32'hc4f4349e, 32'hc2e6bea0},
  {32'hc3a40b57, 32'h453d5a27, 32'h42ffa9fe},
  {32'hc3593f63, 32'h437052aa, 32'h42aa63a6},
  {32'hc46331be, 32'h44df216a, 32'hc3ec8f36},
  {32'h4424b54f, 32'hc4ec3803, 32'h3f188ce0},
  {32'hc52f0534, 32'h42272809, 32'h42fbf723},
  {32'h45005e43, 32'hc3f246ab, 32'hc36da386},
  {32'hc4298b42, 32'h43195ea9, 32'h43ca9d01},
  {32'hc47c5803, 32'hc3e6ab46, 32'h431d75b7},
  {32'hc46a397a, 32'h43a27dec, 32'h44a737c7},
  {32'hc514a23b, 32'h44206d6e, 32'hc4757776},
  {32'h43ce9290, 32'h43dcb7c9, 32'h44e34c88},
  {32'hc4ad51f8, 32'h41f86124, 32'hc37afe0e},
  {32'hc484b08a, 32'h4443c2ff, 32'h43add9e5},
  {32'h44b8fcf2, 32'h42e67afa, 32'hc321a19e},
  {32'hc53165e6, 32'hc18fd811, 32'hc3d4a8f4},
  {32'h4413d8c4, 32'hc4b0a394, 32'hc1b4069b},
  {32'h4427e353, 32'hc36f3f6d, 32'hc434216a},
  {32'h44472de4, 32'hc414f446, 32'hc27fca78},
  {32'hc42960cc, 32'h43e1c4fb, 32'hc3ea0adc},
  {32'h43edc73d, 32'hc401464b, 32'hc3f51a1b},
  {32'hc53dc230, 32'hc4047cb9, 32'h43bbaabf},
  {32'h43fed8c0, 32'hc49ccded, 32'hc41027e4},
  {32'hc436f7ed, 32'h44647817, 32'hc38e386e},
  {32'h430b1cf6, 32'hc3330742, 32'hc4d91cca},
  {32'h43946551, 32'hc414f000, 32'h4499dae4},
  {32'hc447d196, 32'hc3372270, 32'hc41cb1d9},
  {32'hc400c5d8, 32'h4433d423, 32'h44b7d917},
  {32'h4504ddf0, 32'hc30c42c4, 32'hc4364447},
  {32'h43723b7d, 32'h4343948d, 32'h44988f88},
  {32'h447d5a10, 32'hc4eb2671, 32'hc3ecbc10},
  {32'h4352ad11, 32'hc3b2d1c4, 32'h453ec2d1},
  {32'hc4c69eab, 32'hc31bab75, 32'hc3c77507},
  {32'hc55bb8e5, 32'h43ccf003, 32'hc2e2bfb3},
  {32'h45555180, 32'hc41164ee, 32'hc402ec9b},
  {32'h44b06c67, 32'hc27bcc29, 32'hc50f95e3},
  {32'hc41b68e9, 32'hc3503ae2, 32'h44e77c3b},
  {32'hc4abd083, 32'h430f7f32, 32'h4393531e},
  {32'hc36559e8, 32'hc536bf6e, 32'hc2865612},
  {32'h443c5dcf, 32'h4469c98d, 32'h43f3f66e},
  {32'hc3acd95e, 32'hc4c99560, 32'h43b1cd1b},
  {32'h43f07c36, 32'h45279637, 32'h43701ffd},
  {32'hc3e05a4c, 32'hc5204796, 32'h43092e0c},
  {32'h4529f26f, 32'h40bcbc42, 32'hc1086fe8},
  {32'hc2fd35c9, 32'hc3cccc10, 32'h446b99d0},
  {32'h4470ffa0, 32'h4374352d, 32'hc3f8055b},
  {32'h44ce4654, 32'hbcea1d00, 32'hc1b716c7},
  {32'h41d4f3c7, 32'hc3a4a21b, 32'h455ba5b0},
  {32'hc515d424, 32'hc28c8d57, 32'hc1d6ce9a},
  {32'h44d72fcb, 32'h426c5e5a, 32'h413390e5},
  {32'hc463b671, 32'hc35a9931, 32'hc4c9e1f0},
  {32'h4492617b, 32'h441f0a8d, 32'h441d95d0},
  {32'hc3426170, 32'hc45bc58a, 32'hc3c9dd0e},
  {32'h438d0070, 32'hc4463a10, 32'h44ccae64},
  {32'hc5870e2f, 32'hc39ac25b, 32'hc2481aae},
  {32'h454e35c0, 32'h43554cd4, 32'hc453304b},
  {32'hc25e29b4, 32'hc4eddb29, 32'hc410f78c},
  {32'h44f8d5fe, 32'h4424668f, 32'h44013e78},
  {32'hc3da10d6, 32'hc425f055, 32'hc41315f8},
  {32'h439a52ce, 32'h44ee58a9, 32'h42331fbb},
  {32'hc4681c2e, 32'hc4bc8f6a, 32'hc498c0cf},
  {32'h43ec2893, 32'h4460b494, 32'h431b2b4b},
  {32'h45299c92, 32'hc42756a2, 32'h43465243},
  {32'hc49b838f, 32'hc442240b, 32'h42959db0},
  {32'h43dde0fa, 32'h452d71a1, 32'hc294ac95},
  {32'h42f30488, 32'hc3bd3dd2, 32'hc2aa7da8},
  {32'h44d8e019, 32'hc36a49fa, 32'h42636e1d},
  {32'hc3eed37e, 32'hc539959c, 32'h4398ee41},
  {32'h43b79bd4, 32'hc3821096, 32'hc33f7f21},
  {32'hc5785395, 32'h43988932, 32'hc30cc5be},
  {32'hc29088cc, 32'h449ae338, 32'h44762dc2},
  {32'hc50d5cff, 32'h42d2e37a, 32'h442a3b57},
  {32'h43428bd4, 32'h4531de2f, 32'h432499a1},
  {32'h4237ed4c, 32'hc51788ac, 32'hc2983632},
  {32'hc4d6b6e1, 32'h44282428, 32'hc1d07f7c},
  {32'hc3cd65ae, 32'hc4bdd21a, 32'h43260956},
  {32'h44e753c8, 32'hc2a15e62, 32'hc341f070},
  {32'hc50a806d, 32'h42e679de, 32'hc301b5af},
  {32'h4423e9aa, 32'h41421c90, 32'hc4bbbd50},
  {32'hc4dde095, 32'h43a93794, 32'h44042fb6},
  {32'h44cc0b01, 32'h42f314fa, 32'hc4304ac6},
  {32'hc4b3bfd9, 32'hc4b4b1d5, 32'h447a3650},
  {32'hc4572c5f, 32'h43814a23, 32'h42260c56},
  {32'h444ab10f, 32'h430befb2, 32'hc333485f},
  {32'hc4c3a142, 32'hc3d668b8, 32'h42b75dd4},
  {32'hc3b452e0, 32'hc395df92, 32'hc4c23f39},
  {32'hc58c6116, 32'h4382c164, 32'hc19a7b7c},
  {32'h445f52f0, 32'hc3b3670a, 32'hc48d528c},
  {32'h4461b694, 32'hc4be9b45, 32'hc3c7d4f4},
  {32'hc47da7be, 32'h45166e67, 32'h438358a2},
  {32'hc20da2d0, 32'hc48aae3f, 32'hc3acbd5a},
  {32'hc39bbaca, 32'h44c65d4c, 32'hc3a164e1},
  {32'h44f2aceb, 32'hc3fddf13, 32'hc3c6cbe7},
  {32'hc3f89165, 32'h44b9dd4e, 32'h430e20f5},
  {32'h451d735f, 32'hc43a7b13, 32'hc434ecf8},
  {32'hc55d4ca2, 32'h441a2561, 32'hc2025f55},
  {32'h430b59bc, 32'hc44ef43d, 32'h43937814},
  {32'hc4408bd0, 32'h445b1da3, 32'hc4d5ba97},
  {32'h449618bb, 32'hc341bfe6, 32'h444a754c},
  {32'hc40225ec, 32'hc2d51064, 32'h43921715},
  {32'h447d2bbe, 32'hc43efa00, 32'hc39fe185},
  {32'hc4066b93, 32'h440cd28d, 32'hc264814e},
  {32'hc3f5fd02, 32'hc3dcf664, 32'h4417a4c8},
  {32'hc30e1dcd, 32'h43fd2677, 32'hc3fa8def},
  {32'hc293b7f4, 32'h442302e0, 32'h453ef0dd},
  {32'h41e6c940, 32'hc1974b56, 32'hc489c748},
  {32'h4492a97a, 32'hc4ee2297, 32'hc3168d24},
  {32'hc4c385b8, 32'h44672451, 32'hc4524d80},
  {32'h428c5391, 32'hc50233dd, 32'hc4017c93},
  {32'hc31663b0, 32'hc27ec521, 32'hc48d7c08},
  {32'h43621df1, 32'hc2991700, 32'h43ff7b05},
  {32'h4304b48c, 32'h440c3708, 32'hc445601f},
  {32'h44f014f2, 32'h43b1d648, 32'h44abdd04},
  {32'hc2832890, 32'hc493cd77, 32'hc563f4d9},
  {32'h45316e38, 32'hc1d3be41, 32'h423cf7ce},
  {32'h44672274, 32'hc388ffb5, 32'hc525fb6e},
  {32'hc2b52088, 32'h44535e63, 32'h451f22a0},
  {32'h4419b512, 32'h43842543, 32'hc3dbe534},
  {32'h448c0ef4, 32'h4424356a, 32'hc3cf9fe1},
  {32'h44b010d1, 32'hc42f4550, 32'h44190b1c},
  {32'hc384c914, 32'h44fe35b2, 32'hc40f2cd6},
  {32'h4468bae9, 32'h43833383, 32'h44959a13},
  {32'hc3e33fc6, 32'h4473f4b7, 32'hc40c3333},
  {32'h4528edff, 32'hc1e178f3, 32'h44307d17},
  {32'h4452bc26, 32'hc413ac44, 32'h44c048ae},
  {32'hc33e5f7e, 32'h4281e583, 32'hc4c3851d},
  {32'hc3a33f36, 32'h41ccedfa, 32'h4313a6a4},
  {32'hc39fb99a, 32'h42b3a138, 32'h44cb6c55},
  {32'hc39cb239, 32'hc323193a, 32'hc5058034},
  {32'h436c1a63, 32'hc33697dd, 32'h450e1b7e},
  {32'hc4c06dc4, 32'hc379b8fd, 32'h438e0ef8},
  {32'h42f899da, 32'hc54a2d06, 32'h42541852},
  {32'hc4944c46, 32'h42f8768a, 32'hc48a7ab8},
  {32'hc4a54410, 32'hc39e6449, 32'h43a74fd6},
  {32'hc580715f, 32'hc387e260, 32'hc2cedcd6},
  {32'h457fdd41, 32'h43607695, 32'hc44a70d5},
  {32'h43902c31, 32'h442df365, 32'hc45d3c83},
  {32'h4280d0c0, 32'hc437934d, 32'h41e5a29a},
  {32'hc4fa6886, 32'h43ce3e62, 32'hc3ae2a6b},
  {32'h455526a9, 32'h43fb9985, 32'h41fd3558},
  {32'hc4a0647c, 32'h44da17c2, 32'hc27631fe},
  {32'h4528a3fc, 32'hc493592a, 32'h437f1bee},
  {32'hc32c49ca, 32'h44954d7a, 32'h41689b0e},
  {32'h42909f10, 32'hc4b5c0db, 32'hc4971533},
  {32'hc4ccfd91, 32'hc297e6f8, 32'h4333731f},
  {32'hc24e6398, 32'hc28420ae, 32'h44bd869d},
  {32'h42c253c5, 32'h43baf51f, 32'hc4ccd1b4},
  {32'hc455c2a4, 32'hc408c848, 32'h4480f644},
  {32'hc367ea63, 32'h44d1e3f7, 32'hc306c461},
  {32'h430c6f20, 32'hc377cf8c, 32'h4502103b},
  {32'h43ad06eb, 32'h44d56227, 32'hc2cd566a},
  {32'h42fd7c44, 32'h4412362d, 32'hc3882d99},
  {32'hc41801ce, 32'h44707b76, 32'h44e3445a},
  {32'h44d79a82, 32'h443c74f2, 32'hc20b1447},
  {32'hc51cbe70, 32'hc36df922, 32'h434cafc4},
  {32'hc47fe6a6, 32'h4380451c, 32'h4169157a},
  {32'hc3c206fa, 32'hc50abeb3, 32'hc3bd03da},
  {32'h4483a124, 32'h43ccacec, 32'hc32f4848},
  {32'h4358ef42, 32'hc3c9c3f0, 32'h4378bbce},
  {32'h4489f560, 32'hc2dc8853, 32'hc31ed9c7},
  {32'hc58e4f9a, 32'hc2af022a, 32'hc3b6e9c0},
  {32'h451c0734, 32'hc165e239, 32'h43ddd58c},
  {32'hc427376c, 32'hc4abbee3, 32'h438925ae},
  {32'h4411aa80, 32'h450aa698, 32'hc3df6305},
  {32'hc5300fa4, 32'h43302092, 32'h43a994f3},
  {32'h43d7bd9c, 32'h4472e610, 32'h44331636},
  {32'hc562c56e, 32'hc3a4dcca, 32'hc24e0054},
  {32'hc292e264, 32'h443dc873, 32'hc29a6086},
  {32'h448c3cd5, 32'hc43884b0, 32'h43abf324},
  {32'hc3e7a910, 32'hc4eec503, 32'hc3205436},
  {32'h447aed0f, 32'hc4799a94, 32'h442857b0},
  {32'h43058074, 32'hc371e299, 32'hc4854ab0},
  {32'h448bbef6, 32'h43d02d5f, 32'h44d04a6c},
  {32'hc2373ecf, 32'hc33b2479, 32'hc501cbbb},
  {32'hc3914809, 32'h44c3936c, 32'h43900a2d},
  {32'hc3725304, 32'hc433d078, 32'hc53ece69},
  {32'h43b846d3, 32'h44d7fa4e, 32'h445f9310},
  {32'h43ca4d91, 32'h44a55e81, 32'hc3c9e52f},
  {32'h439cd3dc, 32'h45227e90, 32'hc2d3fed6},
  {32'hc3bd4420, 32'h43c3eaf5, 32'hc479254f},
  {32'hc4687c87, 32'h441ce9fc, 32'h42ddea2d},
  {32'hc3a86038, 32'hc404f23e, 32'hc5104a43},
  {32'hc3179e2c, 32'h444b1ea9, 32'h451cf089},
  {32'h4490ac83, 32'hc3c42232, 32'hc29ddd01},
  {32'hc4208f36, 32'h44f65a5a, 32'h44d486c9},
  {32'hc3c8a0b0, 32'hc49be743, 32'hc42ad5f5},
  {32'h438132b4, 32'h4498f326, 32'h43914c5d},
  {32'hc4a3ab72, 32'hc49b3bcd, 32'hc3dbe6e9},
  {32'h445d6148, 32'h45066d96, 32'hc39b40ac},
  {32'hc3d0d1b2, 32'h435139a2, 32'hc29a750d},
  {32'h44cdabce, 32'h431dbc7f, 32'hc28a5000},
  {32'h421f1570, 32'hc52b1ded, 32'hc3bea64b},
  {32'hc494e914, 32'h438cb2bd, 32'hc3eb6441},
  {32'hc568a4d0, 32'h43791d5a, 32'h43d6a3ec},
  {32'h4421f043, 32'hc41ddad9, 32'h43a72da8},
  {32'h4483ad1f, 32'hc3cbf0f2, 32'hc45486e1},
  {32'h44d8af49, 32'h443a11e5, 32'hc3e325da},
  {32'hc21545fb, 32'h44909b39, 32'h44354186},
  {32'h4549c99c, 32'hc2f3ea12, 32'h44057d3c},
  {32'h448fbe8f, 32'hc35dc547, 32'hc2c55d74},
  {32'h43196b88, 32'hc4b1bc46, 32'hc49ba41e},
  {32'hc3b6bb60, 32'h4501938f, 32'h44cb62aa},
  {32'h44af36bd, 32'h4403d600, 32'hc432e708},
  {32'h41b94540, 32'hc4734ba8, 32'h44b44019},
  {32'h44dc89c0, 32'hc22b2dc5, 32'hc3cac566},
  {32'hc4651c54, 32'h4309d85e, 32'h44007bd3},
  {32'h4372aa5c, 32'hc5041dd5, 32'hc0ab2d44},
  {32'hc51c4a9a, 32'h418fcd6c, 32'h440745e6},
  {32'h444f0f66, 32'hc3ab34a7, 32'hc4016427},
  {32'hc3e76782, 32'h4422d19a, 32'h4503038b},
  {32'h4301f73a, 32'hc50ca8ad, 32'hc4f27bf4},
  {32'h43bb37fa, 32'h446706fe, 32'h43e7a0c8},
  {32'h44f55989, 32'hc46a17d4, 32'h4350c49e},
  {32'hc3c60850, 32'h45219b99, 32'hc37303f6},
  {32'h452d5917, 32'h43fb1058, 32'hc3c6187a},
  {32'hc489073c, 32'h45543dc3, 32'h438c917c},
  {32'h45352048, 32'hc36a6a8c, 32'h43840eb0},
  {32'h44fcaac1, 32'h438905aa, 32'hc358eeb7},
  {32'h44e51674, 32'h43e1bfd8, 32'h43692aa1},
  {32'hc4e06b46, 32'hc416d514, 32'h43515425},
  {32'h449c1dba, 32'hc3a3ed21, 32'hc3f298c4},
  {32'hc3247876, 32'h4380d4e4, 32'h437c274a},
  {32'hc527e990, 32'hc397fae0, 32'h43873273},
  {32'hc38799e5, 32'hc40439e9, 32'hc28ba59b},
  {32'h42fdc90b, 32'h45099215, 32'hc3eeedd1},
  {32'hc49da9a8, 32'h44a6ebc4, 32'hc182e235},
  {32'h4495245c, 32'hc25fe7a0, 32'h43904f63},
  {32'hc5897e80, 32'h4308febf, 32'hc18527d4},
  {32'h44ecf967, 32'hc4b70f67, 32'h429bd62d},
  {32'hc5092682, 32'hc2ca42c1, 32'hc226b27e},
  {32'h4425bdbd, 32'hc1adb733, 32'h43f46ed5},
  {32'hc5246665, 32'h43c7a5cb, 32'h43b80dd9},
  {32'h43383eaf, 32'hc319c92c, 32'hc40421ad},
  {32'hc3dadd44, 32'h450ad5a4, 32'h440658e3},
  {32'h44cdb943, 32'h42557b9c, 32'hc4046d60},
  {32'hc449dd12, 32'h4388afc6, 32'hc1f8e66c},
  {32'hc22b5000, 32'hc433d948, 32'hc41cc129},
  {32'hc453a9f8, 32'h44a3810a, 32'hc2fe9c9f},
  {32'h454470a4, 32'h4346bb64, 32'h4396ea50},
  {32'hc54f4c05, 32'h440eb572, 32'h4401f169},
  {32'h44b1f574, 32'hc35675fa, 32'hc44d6103},
  {32'hc41b0af9, 32'h4426c2f1, 32'h43035e09},
  {32'h4423be34, 32'hc49e0667, 32'h42ba4a33},
  {32'h4193d1a0, 32'h418eaf17, 32'h45110fb6},
  {32'h435bc780, 32'hc3337000, 32'hc4c76b63},
  {32'hc3bb7258, 32'h44435bc8, 32'h44bc0f5e},
  {32'h451be5d0, 32'hc4127df7, 32'hc4606e2f},
  {32'h450fd158, 32'h429f9aee, 32'hc43b51ea},
  {32'hc505ab20, 32'hc3566745, 32'h43b58ea8},
  {32'h4488abac, 32'h43de62d7, 32'hc391f880},
  {32'hc51c979c, 32'hc4a9637f, 32'hc445880c},
  {32'h4492b4a7, 32'h44621723, 32'h41c7d50c},
  {32'hc3b52947, 32'hc449ecc4, 32'h434f71a5},
  {32'h43ae350a, 32'h455498b1, 32'h411e4d3f},
  {32'hc4453d32, 32'hc50a58c2, 32'h4368dfec},
  {32'h4528006c, 32'h42e4d6dd, 32'h436224d8},
  {32'hc4c7fa3a, 32'hc303e4fd, 32'h44433454},
  {32'h44d9a20f, 32'hc3c39563, 32'hc1aa4bc5},
  {32'hc4c134eb, 32'h4351be9f, 32'h44062c7b},
  {32'h44d73317, 32'hc2148832, 32'h44718165},
  {32'hc5038a09, 32'hc39579bf, 32'hc4579e41},
  {32'hc4842b97, 32'h438e80a3, 32'h43acdd1f},
  {32'h42f27d80, 32'hc49e5203, 32'hc462f7a4},
  {32'h437e6e66, 32'h44ddc6ac, 32'h41a93c3c},
  {32'hc3230ce8, 32'hc43d8d79, 32'hc3bc907c},
  {32'h45233ceb, 32'h43ac7a52, 32'h4435a5b1},
  {32'hc569336f, 32'h4233360a, 32'hc3c230d7},
  {32'h444cbe3e, 32'h436e4ea8, 32'hc3c0f86f},
  {32'hc3ab2cb7, 32'hc42d04ee, 32'hc4f51aa3},
  {32'h45309930, 32'h43c227ef, 32'h43eac634},
  {32'hc499ea42, 32'hc426e25c, 32'hc2b61ffd},
  {32'h44a22cfe, 32'h43542eea, 32'h43ce5000},
  {32'hc4d0876e, 32'hc46ef6c3, 32'hc47013d3},
  {32'h433c597c, 32'h43ba98d3, 32'h430ce5cb},
  {32'h450b6d44, 32'hc2a5174a, 32'hc38f205d},
  {32'hc5535244, 32'h438b5f58, 32'h4395d85a},
  {32'h44142b12, 32'hc402e356, 32'h448f4a39},
  {32'h44561c7a, 32'hc3531426, 32'hc3601f96},
  {32'h453a07e5, 32'h43de4975, 32'h4327d979},
  {32'hc4a50e52, 32'hc451198f, 32'hc2093121},
  {32'h448df649, 32'hc33dcf23, 32'hc47f2f6c},
  {32'hc4ac1294, 32'hc40206ea, 32'h42ed104d},
  {32'h44f9fbbe, 32'h41b7d35a, 32'hc2392228},
  {32'h44cb9752, 32'h4467e954, 32'hc3c649c1},
  {32'h44c3f7d2, 32'h442e3e30, 32'h43084b58},
  {32'hc4bdd312, 32'hc3742045, 32'hc39ec909},
  {32'hc300b6ac, 32'h42c43a45, 32'hc491c2ad},
  {32'hc4f5563a, 32'hc2fffd1d, 32'h43513dfb},
  {32'h4435bf70, 32'h452c9165, 32'hc0338a6c},
  {32'hc3ee7348, 32'hc38aa52c, 32'h42865b32},
  {32'h45373526, 32'h43ab8579, 32'hc355550c},
  {32'hc51d2634, 32'h4315ea3e, 32'h4353e12b},
  {32'h44e34795, 32'h43cf6e98, 32'hc4806806},
  {32'hc50c850f, 32'hc42f5c84, 32'h438ce743},
  {32'h44b3abb9, 32'hc414f923, 32'hc34aa916},
  {32'hc192d800, 32'h4516e2d3, 32'h422ccfdf},
  {32'hc45bf092, 32'hc4a25e3b, 32'h42f422ff},
  {32'hc4ce891a, 32'h431097b7, 32'hc299cdf8},
  {32'hc53fbe9a, 32'h43753bc6, 32'h42752da5},
  {32'hc315b840, 32'hc381e618, 32'hc55a06e8},
  {32'h453a97ee, 32'hc3c4f789, 32'hc3bc371e},
  {32'hc51cba02, 32'h446d5f53, 32'h440d572b},
  {32'h44b3fa32, 32'h43575e90, 32'h4359c661},
  {32'h433156f5, 32'h455eacca, 32'h429536b2},
  {32'h44f4c547, 32'hc37d17fd, 32'hc2e182c4},
  {32'hc37f00f0, 32'hc2ca0e61, 32'hc34adeb2},
  {32'hc39a34b0, 32'hc2720148, 32'hc414aab5},
  {32'hc4173fce, 32'h4393702e, 32'h437f49b5},
  {32'h450ff4da, 32'h429c92f7, 32'h43d6cef8},
  {32'hc4a29ef0, 32'h445ad4d9, 32'h43e0cfcf},
  {32'h44b6515e, 32'hc3889adc, 32'h42ca6c0d},
  {32'h442a7c61, 32'hc3bb3320, 32'h43f473d4},
  {32'hc2b12754, 32'hc25671de, 32'h44faf3cd},
  {32'h41ec7e20, 32'h44de69be, 32'hc422c206},
  {32'h44123095, 32'h43b9b198, 32'h442bd723},
  {32'hc3696868, 32'hc435fe5c, 32'hc52558ba},
  {32'h43698cc0, 32'hc3a721a9, 32'hc0930b14},
  {32'h44095246, 32'h442a5b4d, 32'h43fc8dc2},
  {32'hc3e07f02, 32'hc49d27b2, 32'h441c829b},
  {32'hc4673697, 32'h448863fc, 32'hc34ab96a},
  {32'h44a135f8, 32'h42d26641, 32'h43b074d8},
  {32'hc44b1f18, 32'h4390076e, 32'hc3c43715},
  {32'h434145ce, 32'hc43b8583, 32'h444dff0e},
  {32'h42a79f56, 32'h4471e773, 32'hc4abef4c},
  {32'h4439cc78, 32'h44339fb4, 32'h45061fc6},
  {32'hc539c4c4, 32'hc32248d4, 32'hc4c6e9d6},
  {32'h44a7bee8, 32'h42513003, 32'h423ce8ba},
  {32'h3fc09700, 32'hc2e9d92b, 32'hc55a0c10},
  {32'h4386db9e, 32'h44890981, 32'h4481662e},
  {32'hc4336654, 32'h43b134d2, 32'hc41a239c},
  {32'h43ab1516, 32'hc349b5ba, 32'hc4ed2866},
  {32'h44266c35, 32'hc4e0877c, 32'h444027b0},
  {32'hc3ef8d23, 32'h44c79e02, 32'hc2e53af3},
  {32'h435e47ae, 32'hc49003ce, 32'h43efd30f},
  {32'hc4655e84, 32'h448595a3, 32'hc4f84e5a},
  {32'h445c8c15, 32'hc3f35dea, 32'h4449cfbf},
  {32'hc3ec0609, 32'h4502eef9, 32'h4517561a},
  {32'hc4aa2cd1, 32'hc3c2849c, 32'hc4316b71},
  {32'hc385f4d6, 32'h448cd213, 32'h4400adcd},
  {32'h4438ffef, 32'hc41a65fb, 32'hc327d065},
  {32'hc4b3243e, 32'h4356ee69, 32'hc4267012},
  {32'h42fd2b18, 32'hc5000a09, 32'h4257e640},
  {32'h44b7e238, 32'hc3dec261, 32'hc462361f},
  {32'hc2e86034, 32'hc4fa3a55, 32'hc2c887a0},
  {32'h40c36780, 32'h4376cad8, 32'hc5187fd7},
  {32'h45467fab, 32'hc30537d9, 32'h44588f77},
  {32'hc59310bf, 32'h4269a530, 32'hc2f20ce5},
  {32'h456e0dd8, 32'h444b9fb8, 32'hc3955eee},
  {32'h44d9da63, 32'h43fbdd40, 32'hc26c4de3},
  {32'h4465f11a, 32'h41d8af58, 32'hc3c89cc6},
  {32'hc3b353de, 32'h44de5dd3, 32'h43fab849},
  {32'h4523192e, 32'h43437ca7, 32'hc34e99af},
  {32'hc528d074, 32'h441f75af, 32'h40c75cb6},
  {32'h44ddf495, 32'hc48393f1, 32'h432b0d9d},
  {32'h4466153d, 32'hc4285d17, 32'h4102d719},
  {32'h44865517, 32'hc377ce56, 32'hc40a99da},
  {32'hc391a0ec, 32'hc5092bb6, 32'h44aa9839},
  {32'hc390c8a8, 32'h425ae928, 32'h440c242e},
  {32'h447cd563, 32'h44b4f1c5, 32'h433874db},
  {32'hc43e94be, 32'hc408a600, 32'hc39a9894},
  {32'h4491bcd6, 32'h4491ed42, 32'hc3974226},
  {32'hc3507b97, 32'hc48392af, 32'h444b4c6d},
  {32'hc4c1e404, 32'h44005361, 32'hc348cbec},
  {32'h445581df, 32'hc43a93db, 32'hc1ecaf82},
  {32'hc5282c68, 32'h440ce681, 32'h448133d2},
  {32'h44107ae6, 32'h43c8afc3, 32'hc4905728},
  {32'hc318186a, 32'h43ccb893, 32'h450741a2},
  {32'hc3f38b1d, 32'h43133a61, 32'hc4367516},
  {32'hc4a89c10, 32'hc408548d, 32'h446534ba},
  {32'h44332e20, 32'h43f52dfd, 32'hc3b52169},
  {32'hc4b3c3d4, 32'hc41e0bcb, 32'hc39a527e},
  {32'h457d54a0, 32'hc340cf80, 32'h42e14d66},
  {32'hc50092f5, 32'h440176a3, 32'hc3f48cda},
  {32'h44c864ab, 32'h44252614, 32'h4358e367},
  {32'hc5350282, 32'hc412bfaf, 32'hc33c1b62},
  {32'h44ec50e2, 32'h4290d5c4, 32'h4194de44},
  {32'hc49ad04c, 32'hc406361a, 32'h439016ce},
  {32'h42873deb, 32'h4558d1aa, 32'h4329162c},
  {32'hc467c30c, 32'hc4f60bb4, 32'hc39d7854},
  {32'h44810026, 32'h42e6b702, 32'h42dc2e37},
  {32'h43fa1eeb, 32'hc44f1242, 32'h438cfc08},
  {32'h433f2286, 32'hc42dae2c, 32'hc476c2c5},
  {32'hc3174560, 32'hc460818e, 32'h44e6a677},
  {32'h4485aec2, 32'hc42a22fc, 32'hc35d99fe},
  {32'h44ca6dd0, 32'h443b0dfa, 32'h4419e024},
  {32'hc4897ec0, 32'hc3a8707d, 32'hc425aec3},
  {32'h45091e49, 32'hc3843533, 32'hc149bbbe},
  {32'hc43dae0b, 32'hc5055f5c, 32'hc48f06f1},
  {32'h44c8f65a, 32'hc3ebb59b, 32'h4441094b},
  {32'h4430f11b, 32'hc23f8876, 32'hc3eea851},
  {32'h448aff14, 32'h43c21f24, 32'h43c73cd7},
  {32'hc236fae0, 32'h44e36df7, 32'hc4d276b0},
  {32'h43fbd068, 32'h446f70a5, 32'hc3a0a484},
  {32'hc4959064, 32'hc40bf4d0, 32'hc3a9c4ec},
  {32'h443823da, 32'h41462aa2, 32'h44ca6b7d},
  {32'hc4a8db86, 32'h438fd743, 32'h437bc7d9},
  {32'hc291cd70, 32'h445f1daa, 32'h44823201},
  {32'h4385365a, 32'hc22203f2, 32'hc437701a},
  {32'h44f0f9cf, 32'h43914222, 32'h42da526c},
  {32'hc500961f, 32'hc489c269, 32'h4349a61c},
  {32'h45163a6e, 32'h447406e0, 32'h43c34677},
  {32'hc396d5f9, 32'hc4ba9303, 32'h43fe3f11},
  {32'h443a471c, 32'h44de6f46, 32'hc3edfa60},
  {32'hc3f95ba8, 32'hc51b39e6, 32'hc3a69758},
  {32'hc42302af, 32'h43629305, 32'h43842212},
  {32'hc514c7be, 32'hc1fad70c, 32'h432cb7d0},
  {32'hc33fa3a0, 32'h4309b162, 32'h43d09b0c},
  {32'h44316067, 32'hc2be833f, 32'hc4544ad9},
  {32'hc2a36843, 32'h442af8fe, 32'hc4b34aa6},
  {32'hc434f19e, 32'h4393a612, 32'h446d1f41},
  {32'h44866de9, 32'hc4a90190, 32'h43a16ec3},
  {32'h449f6d13, 32'h44044739, 32'hc401a54b},
  {32'h44de32de, 32'h436a2b11, 32'hc3f8479b},
  {32'hc4d2c4d8, 32'hc31dd360, 32'h44668b5f},
  {32'h450406ba, 32'h42a5358f, 32'hc3ca0d62},
  {32'h43a28d56, 32'hc3ca944a, 32'h4500f368},
  {32'hc400c5be, 32'h449ebc8f, 32'hc523c237},
  {32'h43a399f3, 32'h44b826e9, 32'hc2c4a955},
  {32'h44f3fe1d, 32'hc4810e46, 32'h41a3fc0e},
  {32'hc295915c, 32'h414f227a, 32'h450f7c65},
  {32'hc479c901, 32'hc29c666e, 32'h415d12dc},
  {32'hc1e06bda, 32'h441a7edb, 32'h45044528},
  {32'hc43e33a3, 32'hc3418738, 32'hc5818d43},
  {32'h44232ee2, 32'h44730e8c, 32'h443183b1},
  {32'h43aa46d8, 32'hc4a9e273, 32'hc1d5ef31},
  {32'h42845f78, 32'h455ef5d5, 32'h42dc7088},
  {32'hc489c609, 32'hc32201ab, 32'h42322462},
  {32'hc43d7a53, 32'h431db56c, 32'h441bacbd},
  {32'hc3823594, 32'hc41fbdbf, 32'h4354d14d},
  {32'h44bab7e2, 32'h43aa84b1, 32'hc3e8d2ce},
  {32'h448315aa, 32'h42ace660, 32'h43d8e200},
  {32'hc4d9bc8b, 32'hc30228ac, 32'hc3a3c85b},
  {32'hc2e0eaf5, 32'hc404d209, 32'hc387398e},
  {32'h44093714, 32'h431714d8, 32'h4130aa04},
  {32'hc56dfa9f, 32'hc39021dd, 32'h43191d33},
  {32'h43046a30, 32'hc2b700f8, 32'h44f671bd},
  {32'hc3da58c4, 32'hc35a0c63, 32'h432bc80e},
  {32'hc306eaf6, 32'h452375ea, 32'hc10e3d7d},
  {32'h450cec52, 32'h42f83de9, 32'h43ece706},
  {32'hc46a3384, 32'h450741d3, 32'hc3810e7b},
  {32'h44063677, 32'hc51c85a3, 32'h433dd20d},
  {32'hc4bf82bb, 32'hc32b429f, 32'h42db7a34},
  {32'h445a752a, 32'hc2d3a9e6, 32'h443e1651},
  {32'hc3aa134d, 32'hc3df8067, 32'hc52d2640},
  {32'h4431942d, 32'hc3b9fa86, 32'hc31b3e5f},
  {32'h441694fb, 32'h43e22077, 32'h44c35338},
  {32'h4418d32c, 32'hc419b67b, 32'hc4cf9d1d},
  {32'hc3cb04a7, 32'h449d0015, 32'h44479cfb},
  {32'h448a4967, 32'h42759122, 32'hc2cdbeff},
  {32'hc3a984b2, 32'h4416e70d, 32'h44a8a208},
  {32'hc3a9c786, 32'hc43833ea, 32'hc3a6c16b},
  {32'hc5233258, 32'hc4706569, 32'h42bc2ca4},
  {32'h441ca770, 32'hc429958d, 32'hc4999c45},
  {32'hc53eefd4, 32'h43e5c231, 32'h41d2c0dc},
  {32'hc3ef609a, 32'hc3d1593d, 32'hc5481f7a},
  {32'hc3dbabe5, 32'h449d5dca, 32'h44036831},
  {32'hc3d01a1a, 32'hc1cd8d5f, 32'hc40086e4},
  {32'hc3a5f03c, 32'h45083f94, 32'h442cf762},
  {32'h42b27350, 32'hc54c00e3, 32'h4220ec06},
  {32'h44a46f30, 32'hc1392d59, 32'hc4a119d6},
  {32'h4297f750, 32'hc3920377, 32'h4537932e},
  {32'h449dd954, 32'h439ce039, 32'hc408b565},
  {32'hc4341e2c, 32'hc4f66ae7, 32'hc2a60700},
  {32'h44adf160, 32'h4439be2e, 32'hc3b8036b},
  {32'h42b58af0, 32'hc36a5039, 32'hc3c3ee7d},
  {32'h4474fd1a, 32'h44ae0ca6, 32'hc2cb3d1a},
  {32'hc54fa063, 32'hc4382321, 32'h4409e158},
  {32'h43877435, 32'h44e4ec67, 32'h4374fa75},
  {32'hc4ce5201, 32'h429de278, 32'h441cdbbe},
  {32'h4405f070, 32'h43db7c48, 32'h43e649d5},
  {32'hc4ba78c1, 32'h437247c2, 32'h43edd234},
  {32'h44fa7ad7, 32'h43a86b2c, 32'h44278353},
  {32'h42559684, 32'hbe1d5ab0, 32'hc44879aa},
  {32'h446af0ee, 32'h4311db2c, 32'h4201bb0e},
  {32'hc4d347c2, 32'hc2a0bbc2, 32'hc487ab06},
  {32'h442ce345, 32'h449ac60a, 32'h449ad30a},
  {32'hc37403d2, 32'hc44b18a7, 32'hc3ee1a7d},
  {32'h43f6702c, 32'h446cd328, 32'h448d78ec},
  {32'hc52a34e4, 32'hc3a317af, 32'hc3d51e49},
  {32'h445f3160, 32'h43215c57, 32'hc3b6b1ae},
  {32'hc2c41210, 32'hc51ffd91, 32'hc3071cea},
  {32'h43e8d2b4, 32'h4481895b, 32'h4447e226},
  {32'h43da7020, 32'hc47b1592, 32'h42ee19bd},
  {32'h42d2d480, 32'h449d1b96, 32'h428ea612},
  {32'hc4d4a228, 32'hc3b9b4b3, 32'hc4c086f2},
  {32'h4459b7f4, 32'h444659b2, 32'hc3e23215},
  {32'h441c041c, 32'h4370f734, 32'hc3ef5571},
  {32'hc39e4dc0, 32'hc4caa904, 32'hc3ab4429},
  {32'h4534cb5a, 32'h4448e388, 32'h43b20cda},
  {32'hc50a8dd0, 32'hc379382a, 32'h436709d2},
  {32'h449740b0, 32'h44311299, 32'hc35b78c9},
  {32'hc4777392, 32'hc2eb6da2, 32'hc297695f},
  {32'hc4e9e443, 32'h439657e5, 32'h42c34e41},
  {32'hc55c2c28, 32'h4420d91b, 32'hc3133940},
  {32'h452d1f9e, 32'h44806843, 32'h443a1806},
  {32'h43fb5c71, 32'hc2a83332, 32'h449a124d},
  {32'h43b9980d, 32'h44823310, 32'hc5051d11},
  {32'hc491de73, 32'hc4681850, 32'hc376c15f},
  {32'hc3f9b268, 32'h43a3988e, 32'hc37d1b4d},
  {32'hc3acf914, 32'hc43872c7, 32'h43a933ee},
  {32'h44bf5a54, 32'hc2f9b27d, 32'hc3df10ba},
  {32'h44a66812, 32'h4288d63c, 32'h4201bfb2},
  {32'h44c1be60, 32'h438db9c9, 32'hc4572508},
  {32'hc47c3264, 32'hc3451d5c, 32'h4447f47e},
  {32'h450e71ac, 32'h42438c8a, 32'h443e60b6},
  {32'hc473c1f9, 32'hc4b57d58, 32'h44691d38},
  {32'h445acd6d, 32'hc3c1c422, 32'h443d8ee6},
  {32'h4487f049, 32'h43e586c6, 32'hc4fb7a58},
  {32'hc4d206f3, 32'hc358832b, 32'hc36f65f2},
  {32'hc330a496, 32'hc2c08c11, 32'hc473ff0b},
  {32'hc57c17c0, 32'h421f2096, 32'h43b5d4bc},
  {32'hc3a24860, 32'h438cd370, 32'hc4b12dd1},
  {32'h45288abb, 32'hc354fe30, 32'hc416c94b},
  {32'hc48e722a, 32'h44b701de, 32'h43a5867b},
  {32'h44c0599a, 32'h430a13e2, 32'h43bd9d84},
  {32'hc506d872, 32'h4468f7b6, 32'h4120934c},
  {32'h4477f6b2, 32'hc4d48605, 32'h43992d43},
  {32'hc3bd4eb2, 32'h44bafa72, 32'h438d2a53},
  {32'h454f49b6, 32'h43a5c97a, 32'h41112536},
  {32'hc541af90, 32'hc28e9092, 32'hc3809841},
  {32'hc2a59e78, 32'hc3fe2643, 32'h4352b12e},
  {32'hc2cdf428, 32'h44875df4, 32'h440e4697},
  {32'h4479df86, 32'hc4270d58, 32'h42b61167},
  {32'hc499c8ea, 32'hc3d92a81, 32'h43b62c54},
  {32'h43a0e306, 32'hc48ec752, 32'h4403ffda},
  {32'hc42a2fc8, 32'h44d2c504, 32'hc374767f},
  {32'hc38eed0f, 32'h430e5014, 32'h44cde3a4},
  {32'hc49c7658, 32'hc2db81e3, 32'hc42a2ed3},
  {32'h44ff8844, 32'h4400c29b, 32'h438071d6},
  {32'hc4dc602e, 32'h42e453e3, 32'hc31380d0},
  {32'h449b6276, 32'hc4bd77b0, 32'h42efdc56},
  {32'hc4944561, 32'h44fa9b7c, 32'hc3222ac0},
  {32'hc48e5755, 32'hc3b19d37, 32'h43240a48},
  {32'hc4f50dce, 32'h43aa5af6, 32'hc3d91e79},
  {32'h44c7e268, 32'hc2b10978, 32'h431d3e3f},
  {32'hc3526a4e, 32'hc2ddff4c, 32'h433a0080},
  {32'h45106d6e, 32'h42c5d63c, 32'h44269558},
  {32'hc530a3e2, 32'h440e0159, 32'hc40183e5},
  {32'h44e57516, 32'h431024c7, 32'hc3ce9ff8},
  {32'hc4e181f6, 32'hc3656ad0, 32'hc4113b98},
  {32'hc4c6af1f, 32'h41776944, 32'h44ae5773},
  {32'h425276dc, 32'h43b74244, 32'hc4222029},
  {32'hc1c0df70, 32'h42c843be, 32'hc28855f3},
  {32'hc3608f64, 32'hc520a9cc, 32'h433da198},
  {32'hc4050f3f, 32'h4496660c, 32'hc40147f7},
  {32'h436d297b, 32'hc49e232c, 32'hc17dfadc},
  {32'h43ae7ca0, 32'h452b673e, 32'hc26686d1},
  {32'h448c1920, 32'hc4176e6d, 32'hc319aacd},
  {32'h431bb628, 32'hc4fdf878, 32'h451f3997},
  {32'hc315da04, 32'h44aab132, 32'hc484f127},
  {32'hc3da3345, 32'h4376a212, 32'h43b575ef},
  {32'h42376d40, 32'hc4aa2378, 32'hc2154770},
  {32'h42adfbf9, 32'hc5392eb1, 32'hc39c35ab},
  {32'hc31760fc, 32'h434d040a, 32'hc4f7a8c3},
  {32'h43f303d6, 32'hc4f7ad31, 32'h4399ecf1},
  {32'h42c99344, 32'h444d123b, 32'hc4e254a1},
  {32'hc4c59ab7, 32'hc397796c, 32'h439d318b},
  {32'hc470cdb3, 32'hc43ba0a4, 32'hc2fa2251},
  {32'hc3eb51bf, 32'h4409b136, 32'h429da1fe},
  {32'hc4d0a403, 32'hc30e8095, 32'hc371a12e},
  {32'h43772a23, 32'hc584807c, 32'hc317ade8},
  {32'hc48a3c4f, 32'h44a3da19, 32'hc3486019},
  {32'h42fc6f58, 32'hc423a421, 32'h4325e817},
  {32'hc3c2c15c, 32'h452f9d93, 32'h4396c4f0},
  {32'h3f99d800, 32'hc507f716, 32'hc30ceb2a},
  {32'hc46efbf7, 32'h43d030c1, 32'hc34b00da},
  {32'hc3991f46, 32'h450eeec9, 32'hc4e94d32},
  {32'hc4ee236a, 32'h42a7af0c, 32'h438c9f9a},
  {32'hc3d3b730, 32'hc48d62e1, 32'h436af5ff},
  {32'h43e53492, 32'h45330634, 32'h4394e28b},
  {32'hc3c0e158, 32'h4386a246, 32'h44b75f03},
  {32'h44029b1f, 32'h43eb478c, 32'hc4b15191},
  {32'h43a85c57, 32'hc52758f2, 32'h43b0cb2b},
  {32'hc495de97, 32'h442a8edf, 32'h42749125},
  {32'h446aa6f0, 32'hc471aa5e, 32'hc3136ad3},
  {32'h4395671b, 32'h44056b16, 32'h45318c12},
  {32'h435892d5, 32'h449ff2d6, 32'h434d0f7f},
  {32'hc3f15ffb, 32'hc3b0d795, 32'h44ce7cb0},
  {32'h448c4501, 32'h42c0814c, 32'hc382a800},
  {32'hc2fb6b01, 32'hc3169a3e, 32'h45307d45},
  {32'h44951d5a, 32'h4410ccd1, 32'hc3f5c334},
  {32'hc3eb89e5, 32'hc4829d86, 32'hc3819f9d},
  {32'h445850c7, 32'hc48bdfdd, 32'h432e4c99},
  {32'hc41cfab6, 32'h43c65e75, 32'h4337aaaa},
  {32'h45572af8, 32'h4340877e, 32'hc3f44aa1},
  {32'hc412d796, 32'hc404ede3, 32'hc2ebf516},
  {32'h43a1d42f, 32'h429028e8, 32'hc3c7500b},
  {32'h44efea3c, 32'hc3d017e9, 32'hc2ccfbc8},
  {32'h447d25db, 32'h44e05112, 32'hc4508792},
  {32'hc4b2a60e, 32'hc46fe8e0, 32'h41985995},
  {32'hc487c561, 32'hc2eba435, 32'h4390697e},
  {32'hc3debf76, 32'h43aa4707, 32'h43e8a6fd},
  {32'hc4f33670, 32'h4374adc7, 32'hc0033554},
  {32'h449da8bb, 32'h44a6f822, 32'h442b154d},
  {32'hc3a553b7, 32'hc3b1c84e, 32'hc4425b38},
  {32'h43135f10, 32'h453a3fb7, 32'h43438f59},
  {32'hc4b2321c, 32'hc38f0d2d, 32'hc4369c42},
  {32'h44ca5a9f, 32'hc38b865c, 32'h44371d7c},
  {32'hc4f92a72, 32'hc3e11b45, 32'hc3945c44},
  {32'hc333f580, 32'h448c6c20, 32'h44942c5c},
  {32'h421727f6, 32'hc4174f97, 32'hc40882c5},
  {32'hc42399b1, 32'hc4ce034e, 32'h451f67ed},
  {32'hc38ac961, 32'h43c91fdb, 32'hc406f200},
  {32'h440c0a1c, 32'h4436783d, 32'hc394356e},
  {32'hc501ae18, 32'hc3a2f5d2, 32'hc20fe0cb},
  {32'h44d3661c, 32'h43ee6379, 32'hc4092ec4},
  {32'h43875cc7, 32'hc3fd5a16, 32'hc500ba62},
  {32'h44a499d9, 32'h43a4e426, 32'h44321224},
  {32'hc410061c, 32'hc4c753e7, 32'hc4830b2f},
  {32'hc3771f9c, 32'h44086fd2, 32'h439e78a5},
  {32'hc44dddc5, 32'hc4b7815f, 32'hc42f3e9c},
  {32'h45059bd0, 32'h44884e69, 32'h441a3ce6},
  {32'hc4a4c6de, 32'h41dfb166, 32'hc2418308},
  {32'h431f4ee0, 32'h445ebc48, 32'h437b8b79},
  {32'hc4c65bb8, 32'hc48d9371, 32'h43b40d76},
  {32'h44f742c2, 32'h44171bbc, 32'h4338ed03},
  {32'hc5868c75, 32'h42b71792, 32'hc2a57090},
  {32'h44e3a730, 32'h4382c116, 32'h4406261f},
  {32'hc48a4238, 32'h4401b5e5, 32'hc4ca5f99},
  {32'hc318697f, 32'hc3196f8e, 32'hc41ba29a},
  {32'hc48e7f33, 32'h43e6fb61, 32'h447f7c2d},
  {32'hc3a8a154, 32'hc2b67a25, 32'hc565b74c},
  {32'hc3203b29, 32'hc2486a52, 32'h4467b012},
  {32'h44b18506, 32'hc33f53a7, 32'hc486734a},
  {32'hc4dc6c58, 32'h4464237f, 32'h424b5f1d},
  {32'h449cfa06, 32'hc2badfea, 32'hc31f52e0},
  {32'hc40b1c8a, 32'hc405d0e7, 32'h443346f5},
  {32'hc3ce6b95, 32'h43e671a5, 32'hc4a425e5},
  {32'hc37e3c00, 32'hc4b3d982, 32'h44705e08},
  {32'hc3c54578, 32'hc4d02af3, 32'hc3fa9b29},
  {32'hc4937a32, 32'h431f5786, 32'h44c48201},
  {32'hc40521f4, 32'hc470274e, 32'hc405e0ec},
  {32'h444a36a1, 32'h4482b9d2, 32'h452d6eae},
  {32'h44b6ff83, 32'hc49918f6, 32'hc450eca9},
  {32'h42f0cc53, 32'h440649c7, 32'h4496de08},
  {32'h43f9a4b4, 32'hc4a168d8, 32'hc487a5f2},
  {32'hc547ab3d, 32'h44539fc2, 32'hc21334a7},
  {32'h4418f3cc, 32'h41bceca8, 32'hc2e1a956},
  {32'hc439a0ee, 32'h450f355e, 32'hc27e9860},
  {32'h42ce86bc, 32'hc571bbb4, 32'hc20ff49a},
  {32'hc539dc98, 32'hc38828ad, 32'hc39e4806},
  {32'h433c9730, 32'hc3f891c6, 32'hc415c8b4},
  {32'hc5842a08, 32'h43704df4, 32'hc3c5c555},
  {32'hc4cd1fb7, 32'hc3d26770, 32'hc42bb36d},
  {32'h44962700, 32'hc2c79ccb, 32'h448342f7},
  {32'hc52bab45, 32'hc35f2a1c, 32'h42d9e6e2},
  {32'h45287ae7, 32'h42744fda, 32'h42b8db98},
  {32'hc5172973, 32'hc3a5a701, 32'hc3a6fcb6},
  {32'hc412cbd7, 32'h44d35793, 32'h43bc177f},
  {32'hc4c6cfcd, 32'hc3652dcc, 32'h43e33634},
  {32'hc450ef95, 32'h45327d2a, 32'hc2ef2590},
  {32'h446ab1a0, 32'hc4622f61, 32'hc395ed53},
  {32'h44131042, 32'hc3df3107, 32'hc4d99e6e},
  {32'h44109bc4, 32'h43f16c7b, 32'h450797c4},
  {32'hc4a89e76, 32'h44137303, 32'hc4c8f1fe},
  {32'h4484a8f8, 32'hc36808a7, 32'hc282f341},
  {32'hc526938b, 32'hc2909dfb, 32'h42b90c8c},
  {32'h44406ffb, 32'hc4a76d2f, 32'h410bdbe0},
  {32'hc53436c4, 32'h42a89f91, 32'h418cd90c},
  {32'h44897cec, 32'h441c5f8c, 32'hc49eea78},
  {32'hc42aafc4, 32'h44307c49, 32'h448dd86e},
  {32'h44dee220, 32'hc33de7e0, 32'hc2d39aa2},
  {32'hc48f67c8, 32'h42910429, 32'h4462ccb4},
  {32'h454a7908, 32'h4306e872, 32'hc3fde907},
  {32'hc4ec00e4, 32'hc3be7dd7, 32'hc266973b},
  {32'h4420b694, 32'hc4ce3fdc, 32'hc2421588},
  {32'hc249ff50, 32'h450509c6, 32'h4417795d},
  {32'h42d1e7fc, 32'hc44161db, 32'hc339629f},
  {32'h4357f13c, 32'h450b97e2, 32'h445fd996},
  {32'h4410ee5a, 32'h42b52913, 32'hc51733c8},
  {32'h45174083, 32'hc3509a8c, 32'hc3e80692},
  {32'hc4966bf2, 32'h439ed1ac, 32'h445e257f},
  {32'hc4bcb29b, 32'h437d7eab, 32'hc02760e0},
  {32'hc4c8999c, 32'hc42cb154, 32'hc43321de},
  {32'h4484042f, 32'h4495f8d4, 32'h43fb115d},
  {32'hc46bfe20, 32'hc38d581e, 32'hc43abe6f},
  {32'h4466f970, 32'h4498706e, 32'hc38eac22},
  {32'hc470ca7d, 32'hc5262c6a, 32'hc360933c},
  {32'hc488636e, 32'h43d7ce27, 32'hc3807ede},
  {32'h429eb9c8, 32'h4192f70f, 32'h43bd738a},
  {32'h43d3e96c, 32'h43cfacec, 32'hc4b7bf07},
  {32'h4408eeec, 32'hc3a4862f, 32'h443ad237},
  {32'h440275cf, 32'h445f92ae, 32'h43395ddb},
  {32'hc55c6e45, 32'hc3f93be1, 32'h43698af5},
  {32'h44ccfbf2, 32'hc20ddba0, 32'h439f6353},
  {32'hc2be32a6, 32'h41f03794, 32'hc55e9087},
  {32'hc2aa20d5, 32'h43d6de4c, 32'h4509ff10},
  {32'hc4e1caf8, 32'hc307d815, 32'hc31ceb01},
  {32'h453cf82a, 32'hc30f5063, 32'h441664b7},
  {32'hc4e8318c, 32'h43da02cc, 32'hc491e73c},
  {32'hc40e1a48, 32'hc2af2649, 32'hc3e18bbe},
  {32'hc33bde30, 32'hc40d2599, 32'hc507f6a7},
  {32'h42e82b7c, 32'h4512b021, 32'h433da93f},
  {32'hc478b5d9, 32'hc3149390, 32'hc2924e04},
  {32'h44ac8095, 32'h43ff0efb, 32'h441c0997},
  {32'hc5129dac, 32'h42d0fa52, 32'hc42b23bd},
  {32'hc386fb12, 32'hc382c3ef, 32'h443720f4},
  {32'h450a24ea, 32'hc3fac2ad, 32'hc3c554f4},
  {32'hc39bb700, 32'hc534d45e, 32'h434c699c},
  {32'h452c05f0, 32'h438985cf, 32'h43e5901a},
  {32'h44973d98, 32'hc366d1fc, 32'hc240663a},
  {32'h439a3bc8, 32'h452220d1, 32'hc3ab64f9},
  {32'h43a20983, 32'hc58967ad, 32'h4247b4a2},
  {32'h44259022, 32'h442c1bd0, 32'hc3f97a04},
  {32'hc402e108, 32'hc3f6da77, 32'hc43afe5c},
  {32'h450ab13d, 32'h4428789e, 32'h443d9b96},
  {32'h440db50c, 32'hc445f667, 32'h43db6622},
  {32'h43aa4366, 32'h442b5657, 32'h42dd0dee},
  {32'hc3ee24ad, 32'hc42b7c8a, 32'hc2d78663},
  {32'h450244b0, 32'h43ca0151, 32'hc337e137},
  {32'hc3a3b377, 32'h438167d3, 32'h44d2631c},
  {32'h441b456e, 32'h42da691a, 32'hc52ec06f},
  {32'h44518ef0, 32'hc334f2eb, 32'h44488a5e},
  {32'h438fc8fc, 32'h43b9b718, 32'hc47d86ef},
  {32'hc4291c67, 32'h43f39107, 32'h452a6d38},
  {32'hc3916fc4, 32'h440fdef0, 32'h42bee36f},
  {32'hc529e87d, 32'hc4004180, 32'hc2d547be},
  {32'hc3abbd0b, 32'h431bc3e2, 32'hc2b6b1da},
  {32'hc3294f42, 32'hc3786828, 32'hc51ffdf3},
  {32'hc48e96ac, 32'hc42358c9, 32'h4450152f},
  {32'hc3f15ffb, 32'h43c1db43, 32'hc20121f1},
  {32'hc32b7188, 32'h440edb30, 32'h456b5d1c},
  {32'h450e5c60, 32'hc320876f, 32'hc492a036},
  {32'hc30a0251, 32'hc547a55f, 32'h41a61059},
  {32'hc3fc0be0, 32'h4492e168, 32'h442f741a},
  {32'hc4926744, 32'h43b2749d, 32'hc38f0618},
  {32'hc535ad72, 32'h4462af43, 32'h43aa0f23},
  {32'hc292bba8, 32'hc537f035, 32'hc34ae145},
  {32'h4464c396, 32'h4307377d, 32'hc3a66ea7},
  {32'h44c7695e, 32'h43bcef7d, 32'hc3134469},
  {32'hc509fefb, 32'h43b9a642, 32'h435cf55e},
  {32'hc4d649f6, 32'h4204c4c6, 32'h438dadf6},
  {32'h43926534, 32'h443b14c3, 32'h44252c8e},
  {32'h448659d0, 32'h447a9630, 32'hc4761157},
  {32'hc4e4f5dc, 32'h43221a9e, 32'hc42a62e4},
  {32'h4448c184, 32'h4357b057, 32'h44a4f939},
  {32'hc42e0746, 32'h44b491f5, 32'hc403c67c},
  {32'hc2844e68, 32'h426e9f66, 32'h44291266},
  {32'hc4a9110a, 32'h441a437d, 32'hc1ec3b24},
  {32'h451559cb, 32'hc45d7fd6, 32'hc3bbcadb},
  {32'hc3e81aeb, 32'hc3a05b03, 32'hc4557021},
  {32'h45352b9d, 32'hc4870752, 32'h439db3d3},
  {32'hc52f9294, 32'h448fca8c, 32'hc3b9d855},
  {32'h44998739, 32'hc28ced09, 32'hc1564a8e},
  {32'hc398be2c, 32'h44e90eff, 32'hc3e2b842},
  {32'h444a221c, 32'hc414d81f, 32'h44d3d1ae},
  {32'h4459316e, 32'h3fa04af7, 32'h4387f96d},
  {32'h45080611, 32'h4221a767, 32'h444153ef},
  {32'hc3cd964c, 32'hc20d3aed, 32'hc54fc431},
  {32'h44ec24e0, 32'hc33e90a5, 32'hc30b412b},
  {32'h445728f5, 32'hc4b4fa58, 32'hc4b6146b},
  {32'hc329f8e8, 32'h4446d817, 32'h44b6fba9},
  {32'hc44b437b, 32'hc4ccd23f, 32'h406a3716},
  {32'hc45e3791, 32'h42e8550f, 32'h418d5b1d},
  {32'h44315074, 32'hc317b68f, 32'h4489430d},
  {32'hc40f02e7, 32'hc266c0e3, 32'hc4c207f6},
  {32'hc4b9f46c, 32'hc2b937d9, 32'h41cd783a},
  {32'hc4838f4e, 32'h43c9bbd5, 32'hc4554920},
  {32'h44927d75, 32'hc4454c5a, 32'hc3d22800},
  {32'hc44d98a9, 32'h43b7afa8, 32'h454e81d0},
  {32'h43be811a, 32'hc419704e, 32'hc508ee9c},
  {32'hc35929ce, 32'hc131b9d1, 32'h44b72343},
  {32'h43735df3, 32'h42607964, 32'h44e7b4a3},
  {32'h44c40b79, 32'hc335d262, 32'h4401f9f1},
  {32'h43c32640, 32'h44bd5cfc, 32'hc39db752},
  {32'hc2e26210, 32'hc30ec69c, 32'h43f33018},
  {32'h42af7be4, 32'h44237108, 32'hc4fe0cf5},
  {32'hc3c0b08e, 32'h42944779, 32'h43d49150},
  {32'hc59d8709, 32'h4300c9e4, 32'hc2829ef5},
  {32'h44c3844c, 32'h43954656, 32'hc38455b7},
  {32'hc4c963ec, 32'h42d0cd6d, 32'hc35acf0a},
  {32'hc37dd870, 32'hc5293cb7, 32'h41e5c690},
  {32'hc5330523, 32'h4389fbca, 32'h43f3bf11},
  {32'h45177c41, 32'hc27cd0f4, 32'h437ddb32},
  {32'hc44c1860, 32'h451a3885, 32'h4332066a},
  {32'hc29d21bd, 32'hc58072c1, 32'h432d5e89},
  {32'hc2ea2885, 32'hc3e89869, 32'h43cda603},
  {32'h444f786f, 32'h4317d478, 32'hc475be5a},
  {32'hc43199f7, 32'h43489003, 32'h448a4e86},
  {32'hc30f93a4, 32'hc4c1abd1, 32'h43682193},
  {32'h4442ec8c, 32'h4400a50d, 32'hc402a20a},
  {32'h4369ead0, 32'hc373dbfb, 32'h43e99ee5},
  {32'h44403728, 32'h4426316f, 32'hc4e5e713},
  {32'hc40f1b42, 32'h4335fd50, 32'h454b9fca},
  {32'h4311e935, 32'h4404fc0b, 32'hc4b036f0},
  {32'h44a31b27, 32'h438013cc, 32'h436cb72a},
  {32'hc3c4a8da, 32'h4504f8cf, 32'h44d21984},
  {32'h441ca564, 32'h440c9fc5, 32'hc4a9b7aa},
  {32'hc45f6e23, 32'hc49602ce, 32'hc110e4b8},
  {32'h43bc6e62, 32'hc2f32421, 32'hc43bd0d1},
  {32'hc3f303dc, 32'hc4e905c7, 32'hc3949303},
  {32'h44d40eae, 32'h427a6a48, 32'hc35c2e2f},
  {32'hc30503d3, 32'hc46dbf0c, 32'h43e43218},
  {32'h44e3ee2c, 32'hc3a1f630, 32'hc1990c52},
  {32'hc5496a15, 32'h42724d42, 32'hc364fe7a},
  {32'h4565106e, 32'h42fed825, 32'hc2e7cc5f},
  {32'hc2501f16, 32'hc4fd5d18, 32'hc35eed62},
  {32'h44c26b0b, 32'h4422b767, 32'h42adcc5f},
  {32'h43e11089, 32'hc31e5a5e, 32'h438c87ad},
  {32'hc3b20906, 32'h453d0a73, 32'h43df642c},
  {32'hc56ba059, 32'hc36b77a9, 32'h42482061},
  {32'hc4502435, 32'h442d8229, 32'hc391a7da},
  {32'hc3d4a516, 32'h445a7076, 32'hc2f68736},
  {32'hc30e7300, 32'hc4df89c2, 32'hc41061f2},
  {32'h4341a665, 32'h45115eb6, 32'h4323c0dc},
  {32'hc48d2fd4, 32'h41603862, 32'h430b26b9},
  {32'h43b832c4, 32'h447f16ce, 32'h448e6e9e},
  {32'hc31eb8a0, 32'hc389e9e8, 32'hc486593e},
  {32'h445bfd1c, 32'hc480fe91, 32'hc369072e},
  {32'hc55cacdb, 32'h41d55f35, 32'hc22e2f9f},
  {32'h43b413dc, 32'h44d6be62, 32'h445825d2},
  {32'h43aacb1e, 32'hc4600e04, 32'h43380234},
  {32'h441f62d6, 32'h437daa83, 32'hc398d63a},
  {32'hc40fcf80, 32'h44195835, 32'hc4c414cb},
  {32'h42bec4ec, 32'h44fe9c6c, 32'h4371eb20},
  {32'hc49a6442, 32'hc44f091d, 32'hc3a2f519},
  {32'h4505577c, 32'h4301642c, 32'hc40dd637},
  {32'hc4c67f71, 32'hc2ab00e4, 32'h43942820},
  {32'h453b60b6, 32'h437a5109, 32'h4403c86f},
  {32'hc4bc7026, 32'hc3aac0f9, 32'hc34beaa6},
  {32'h434511e4, 32'h44bfe18e, 32'hc2f2ebaf},
  {32'hc5432f12, 32'hc43c08a4, 32'hc3dde904},
  {32'h44ee2837, 32'h446f6580, 32'h4409d598},
  {32'hc48d1512, 32'h430a8feb, 32'hc2ef4bf1},
  {32'h447f4754, 32'h446e73e8, 32'h4417a200},
  {32'hc4aa0714, 32'hc4dd17ff, 32'h43508659},
  {32'h445237c2, 32'h4218a070, 32'h43616643},
  {32'hc470f034, 32'hc3fae027, 32'hc079ca10},
  {32'hc312c0f0, 32'hc4632d9f, 32'h4421aa46},
  {32'h4357a178, 32'h448f4792, 32'hc50bb37a},
  {32'hc4705fcb, 32'hc4dee1c8, 32'hc1ce84a6},
  {32'hc434a423, 32'h43039197, 32'h44b87f62},
  {32'hc0870d80, 32'hc44bba04, 32'hc4bee80d},
  {32'h441a9e51, 32'h43fe46a9, 32'h44cecd71},
  {32'h41ef3580, 32'hc4ecdac4, 32'hc5176c94},
  {32'hc317972c, 32'h43459956, 32'h4507b907},
  {32'hc3e7235a, 32'hc417ebd8, 32'hc2815eaa},
  {32'h43f7ef18, 32'hc4ebdb88, 32'h44e5f0b2},
  {32'hc407cd1c, 32'hc49a45ed, 32'h4393bd8d},
  {32'hc4ca6b6a, 32'hc39c25e0, 32'hc3547c6e},
  {32'h445e9d28, 32'hc28f5867, 32'hc3e4f90a},
  {32'hc3cc4167, 32'h441b8699, 32'h444bc7f0},
  {32'h43cde984, 32'hc3a8b225, 32'hc3544fc8},
  {32'hc4c57759, 32'h43cc6914, 32'h441f6ac4},
  {32'h42c9b278, 32'hc4332520, 32'hc427cb8f},
  {32'hc4546bc9, 32'h439be4d3, 32'h43951176},
  {32'h446d6190, 32'hc50551b3, 32'hc2d70130},
  {32'hc5012dfc, 32'h448fdcac, 32'h4378d8a5},
  {32'h441bc131, 32'hc500088a, 32'h43ffb075},
  {32'hc4a3e1b4, 32'h44c2af54, 32'h413320ff},
  {32'h43d3d211, 32'hc5880fe5, 32'h429ec21e},
  {32'hc4d49b66, 32'h4347d326, 32'h42a65bb6},
  {32'h44de1c42, 32'h436ed973, 32'h436ee1b8},
  {32'hc4ed3542, 32'h42f09852, 32'h425180ef},
  {32'h454c5664, 32'h41193c7a, 32'h438ef749},
  {32'hc2f63120, 32'h433fa31f, 32'hc1b8df48},
  {32'hc53035f4, 32'h4342cf13, 32'h431ddca9},
  {32'h44d19513, 32'h43144fde, 32'h44c3b241},
  {32'h4350da60, 32'h4418789e, 32'h441dda72},
  {32'hc48b72c6, 32'h4477af71, 32'h42c09d72},
  {32'h4528b1ac, 32'h43353fd6, 32'h43b96cf3},
  {32'h431338d0, 32'h451d6487, 32'h44121916},
  {32'h4452384c, 32'hc4caec09, 32'hc211915c},
  {32'hc496467a, 32'hc417d3c0, 32'h43f023b9},
  {32'h4429ef2a, 32'hc360fe5e, 32'h451c7a09},
  {32'hc48aa644, 32'hc3b4e940, 32'h43f54787},
  {32'h443fa6c6, 32'hc3b54f5a, 32'hc45253b9},
  {32'h4358be2a, 32'hc4f4e4ab, 32'hc37ed228},
  {32'h45082947, 32'h4333eef0, 32'h437902e9},
  {32'hc3a36dea, 32'hc44c27f4, 32'hc4484316},
  {32'hc3a1e7ee, 32'h448c61f3, 32'h44676ebb},
  {32'hc480058c, 32'hc41cfc50, 32'hc3131ba4},
  {32'hc512d28a, 32'h442e1eef, 32'h44830a5c},
  {32'h44fc9206, 32'h436aa0ea, 32'hc3896cce},
  {32'h437a70ac, 32'h449afdea, 32'hc310b3f4},
  {32'h424dbf48, 32'hc4aea59f, 32'hc4af85e2},
  {32'hc4f10034, 32'h4337118b, 32'h44780cfe},
  {32'h429359c6, 32'hc32c166d, 32'hc5179f91},
  {32'hc4bd42ed, 32'h44fff253, 32'h437ad3c3},
  {32'h44831e99, 32'hc43cda49, 32'hc4898134},
  {32'h44ec64fd, 32'hc19175c1, 32'hc41fab87},
  {32'hc4e8d6d7, 32'h42becd7a, 32'h43e6b88b},
  {32'h44222e17, 32'hc41c1bf8, 32'hc48aa5e5},
  {32'hc5280d40, 32'hc443c851, 32'hc360c326},
  {32'h44276fd0, 32'h447aa8fc, 32'hc2f2abeb},
  {32'h43a7ec86, 32'h43104b17, 32'hc28cf687},
  {32'h43d8e0a8, 32'h4564b494, 32'h419e9f28},
  {32'hc4016069, 32'hc518bf00, 32'hc2d85810},
  {32'hc33cbf4b, 32'hc38229aa, 32'h432bc462},
  {32'hc43ee562, 32'hc450bfdf, 32'hc4427fa4},
  {32'hc130a8c0, 32'h42a7f150, 32'hc530273b},
  {32'h44577986, 32'hc40dbd44, 32'hc2ea89c0},
  {32'hc29844e9, 32'h44fb75c1, 32'h4403e344},
  {32'h4327e74f, 32'hc51ae8ef, 32'h4363497f},
  {32'h45152536, 32'h43aa57e9, 32'hc2eb1c7a},
  {32'h426c88a8, 32'hc4993d7c, 32'hc47d77d0},
  {32'hc25064a2, 32'h44882493, 32'h4389dfff},
  {32'hc1ae51c0, 32'hc4c3e7bd, 32'hc350c01b},
  {32'h44b22e35, 32'h4432a909, 32'h44b576d4},
  {32'hc583b352, 32'h42767bf2, 32'h42d790a1},
  {32'h44ceb192, 32'h431b80d2, 32'hc311fe0b},
  {32'hc4e81cda, 32'hc3f482fa, 32'hc4868a83},
  {32'h4545c348, 32'h43b07879, 32'h438cf690},
  {32'hc49c59b8, 32'hc4083930, 32'hc28c009f},
  {32'h4565ade6, 32'h438433fd, 32'h4368e586},
  {32'hc381eb84, 32'hc42fd921, 32'hc556e330},
  {32'h440733a2, 32'hc3210bc5, 32'h431dd769},
  {32'hc3878ea9, 32'h4473f5b0, 32'hc3c487a1},
  {32'hc4b2b2ec, 32'hc3e8f6ae, 32'hc40ad4a8},
  {32'h452cedb2, 32'h438aa24b, 32'h4405cd03},
  {32'hc477239e, 32'h440669ac, 32'hc1993e56},
  {32'h43f5220e, 32'h44a80e3e, 32'hc36da696},
  {32'hc454ec09, 32'hc50776ac, 32'h41822c54},
  {32'h4512fecc, 32'h42216020, 32'hc3302254},
  {32'hc57bfa1a, 32'hc1bb3056, 32'h4382bbe0},
  {32'h4527ed70, 32'h434f7e14, 32'h436ce2f4},
  {32'h44875749, 32'h43af920e, 32'h42c67aff},
  {32'h449ea678, 32'h434a6da0, 32'hc3ad5795},
  {32'hc441e4f3, 32'hc4e23b75, 32'h430a5cfd},
  {32'hc400fec1, 32'h43c33d3c, 32'hc4187a28},
  {32'hc4288dfc, 32'hc47319fa, 32'h43e31b14},
  {32'hc3d60750, 32'h441834ee, 32'hc49a4bb6},
  {32'hc3e0d97e, 32'hc272c709, 32'h443f32f2},
  {32'h44437a8e, 32'hc15d86e2, 32'hc48861f3},
  {32'hc40090cb, 32'hc3a94aa3, 32'h43340496},
  {32'hc346856c, 32'h44e0e363, 32'hc35d33cc},
  {32'hc4e22730, 32'hc469b55e, 32'h4417d53a},
  {32'h4380fc60, 32'hc3046f23, 32'h439651e6},
  {32'h432ed331, 32'h451ffa7d, 32'h42299270},
  {32'hc41ec569, 32'hc30fc241, 32'h451c7332},
  {32'hc44b9776, 32'h43dcb6bb, 32'hc321044b},
  {32'hc418082b, 32'h43250d0e, 32'h45272b4e},
  {32'hc378ca20, 32'h432f4174, 32'hc4b0dc36},
  {32'h4506e210, 32'hc425b714, 32'hc427cde2},
  {32'hc49d6a56, 32'hc3b40c94, 32'h44d938c1},
  {32'h448adc2e, 32'hc40c2993, 32'h4175c446},
  {32'hc39ab4ff, 32'h43bfaa13, 32'hc357f23f},
  {32'h4550ef05, 32'h41c9fdf8, 32'hc3d74800},
  {32'hc2b33182, 32'h44bdbe7a, 32'hc380a276},
  {32'h4554194e, 32'h41e00fa8, 32'hc38fc8db},
  {32'hc5439bff, 32'h4413f1cb, 32'h438b5c00},
  {32'h454aca35, 32'hc282d9eb, 32'h44139bc4},
  {32'hc306185e, 32'h45251b6c, 32'h42d8ac7f},
  {32'h42e9101d, 32'hc48db3ae, 32'h43f39f76},
  {32'hc3407e39, 32'h43a1e5b8, 32'hc4ae08d7},
  {32'h443dab4f, 32'hc4a615ab, 32'hc10f101e},
  {32'hc4361cd4, 32'h4435b3e5, 32'hc481fb28},
  {32'h449beeb4, 32'hc3291a9a, 32'h410504ee},
  {32'hc3153f20, 32'hc3827f5b, 32'hc5291a2c},
  {32'h44fc6e1a, 32'h42ffa0dc, 32'h43251be4},
  {32'h41c753e0, 32'hc3abd26b, 32'hc4e7326c},
  {32'h43f16ebc, 32'hc2a43156, 32'h450ff5cb},
  {32'hc4d2c722, 32'h449d9a57, 32'hc40abaa2},
  {32'h44ef4e48, 32'h4297e22b, 32'hc384d7c8},
  {32'hc3c55e80, 32'hc335688e, 32'hc4a5bfe3},
  {32'h433ef3fc, 32'h41b66fa4, 32'h451b9658},
  {32'h44641720, 32'h4242ff46, 32'hc3539f77},
  {32'h44825d68, 32'hc38e8627, 32'h436b7462},
  {32'hc5019f26, 32'h43abe0b2, 32'hc49c2df0},
  {32'hc4b9dcbe, 32'hc3864498, 32'h43dc0cab},
  {32'hc4c955cd, 32'hc20ccc5b, 32'hc3f0538b},
  {32'h43b9d8fa, 32'hc4c2776b, 32'h450ce0b6},
  {32'hc3ff828a, 32'h4399ed91, 32'hc2f17492},
  {32'h449cd527, 32'h4305ed2e, 32'hc388779c},
  {32'h4483ed3e, 32'hc4b5b9e9, 32'h43d35830},
  {32'hc1af8398, 32'hc3bc26fb, 32'hc4dbd58c},
  {32'h4285d78a, 32'h42d20d7d, 32'h44c1feea},
  {32'hc4b94b87, 32'h448359c6, 32'hc3eccdf7},
  {32'h438c6f98, 32'hc47aa01d, 32'h451221e1},
  {32'h45205ef6, 32'h4430cb31, 32'h4480278d},
  {32'h4381d96b, 32'hc5256799, 32'hc4b5a8c6},
  {32'hc3af0716, 32'h448da9b3, 32'h43843227},
  {32'hc2532a20, 32'h432611ce, 32'h43e96d66},
  {32'h43105150, 32'h438bc065, 32'h445709cb},
  {32'hc4ed8952, 32'h4328ca6c, 32'h44101ffe},
  {32'h44024169, 32'hc5049d5d, 32'h4347b008},
  {32'hc4033bdb, 32'h448ceed9, 32'hc434cf06},
  {32'h4518a3ea, 32'hc40c8211, 32'h441009d1},
  {32'hc5583428, 32'hc3dd3dfa, 32'hc38bc22a},
  {32'h4556a8fc, 32'hc0db850e, 32'h441c83b3},
  {32'hc4e42377, 32'hc263664d, 32'h427faf99},
  {32'h44ce4217, 32'hc41370da, 32'h43d97f20},
  {32'h42bc6580, 32'h451b667e, 32'h439df817},
  {32'hc495ba0f, 32'hc37ee1c3, 32'hc391cbaa},
  {32'hc4210ca0, 32'h4537b048, 32'h40a3cac8},
  {32'h451cfca4, 32'hc48a9f88, 32'h42756d5f},
  {32'h42891838, 32'hc4c3fb2a, 32'h44616a48},
  {32'h44429c3e, 32'h432ef24d, 32'hc2d2370c},
  {32'hc4be0904, 32'h441b92d9, 32'h444f8701},
  {32'hc4b9edf7, 32'hc432744c, 32'h4323e22a},
  {32'h43a232ab, 32'h44e7eba5, 32'hc2b9e69c},
  {32'hc29322e0, 32'hc4700b39, 32'h443bd4e5},
  {32'hc143a380, 32'h448fa1a6, 32'hc4a409e7},
  {32'hc46c1b99, 32'hc49277ac, 32'h427ae2d5},
  {32'hc1f12638, 32'h44eba3f2, 32'h436f0e67},
  {32'h43e7b03a, 32'h448efd56, 32'hc388c47b},
  {32'hc4ac24c5, 32'hc283d5a6, 32'h44858703},
  {32'h448ab10e, 32'h44564a5f, 32'hc3e2465c},
  {32'hc390086e, 32'hc330794a, 32'h4547946b},
  {32'hc294589d, 32'h43400518, 32'hc4677757},
  {32'hc3ae6cc3, 32'hc4dc8003, 32'h43a949f8},
  {32'h432d026d, 32'h4500a8e1, 32'hc43244a1},
  {32'hc395d10c, 32'hc384499a, 32'h43c73c54},
  {32'h44dd51bc, 32'hc4101e9f, 32'hc3c70356},
  {32'hc4c86f49, 32'h431b7b01, 32'h422ddba4},
  {32'hc47d3aa6, 32'hc52b4c6b, 32'h42bd07cf},
  {32'h4580053d, 32'h4376e5ea, 32'h43e09d91},
  {32'hc189fca4, 32'hc3b78806, 32'h4399d9fa},
  {32'hc39eee5b, 32'h44ba573e, 32'hc36e2ed5},
  {32'hc4d4f658, 32'hc4506f8d, 32'h420f7cb6},
  {32'h45307b01, 32'hc40da5e6, 32'hc40c3e07},
  {32'h44a3e388, 32'h433ff93d, 32'h430f2a1c},
  {32'hc379ce86, 32'h4494ac75, 32'hc51304d1},
  {32'h42d27bfa, 32'h4299d3ef, 32'hc13ca52c},
  {32'hc37aa7a0, 32'hc41b906d, 32'hc3b63467},
  {32'h45185bf2, 32'h42a87a7b, 32'h44291b8d},
  {32'hc4595716, 32'hc47e5559, 32'hc389dd2a},
  {32'h45555469, 32'h42973b59, 32'hc248f0a5},
  {32'hc395ce40, 32'hc3e69754, 32'hc4e9691b},
  {32'h441fed4f, 32'h44c1d841, 32'h44bf9297},
  {32'h439b1dd8, 32'hc4f22176, 32'h439a3738},
  {32'h43a7c0fe, 32'h44555e0e, 32'hc3694ac6},
  {32'hc33e757c, 32'h449c0a74, 32'hc5434a83},
  {32'hc34de7ad, 32'h43dea0ec, 32'h44be8437},
  {32'hc3afb09c, 32'hc4c15dac, 32'hc2e54e2a},
  {32'h43aecb3d, 32'h44bdb37d, 32'h44533a73},
  {32'hc3da6309, 32'hc14b91c6, 32'hc460a128},
  {32'h44edbdf0, 32'h43caffe4, 32'h4428f970},
  {32'h4395e90a, 32'hc327dc64, 32'hc5304ee8},
  {32'hc4264165, 32'h4472d0d1, 32'h42ec8954},
  {32'hc583b2ac, 32'hc3454ca6, 32'hc30b4716},
  {32'h45178da4, 32'h445344cf, 32'hc36210b3},
  {32'h43134fd4, 32'hc3316f24, 32'hc3fa1acf},
  {32'h447e3512, 32'h44a1d7c6, 32'h43f16d8f},
  {32'hc5380b10, 32'hc3222383, 32'hc1a2819a},
  {32'h4530f6f3, 32'h44275e06, 32'h43834fc4},
  {32'hc50ddef4, 32'hc2d68453, 32'h422da5e3},
  {32'h444ecf50, 32'hc3c0e81e, 32'h4412c644},
  {32'hc3a7424b, 32'hc3592150, 32'hc3c9182e},
  {32'hc20e24e8, 32'h4496e3ac, 32'hc4088789},
  {32'hc491d192, 32'h442adbb9, 32'h43aa15e6},
  {32'hc3e452a4, 32'hc3ed5cbb, 32'hc4b8727b},
  {32'h43ff1689, 32'h4403b8db, 32'h43d85824},
  {32'h440231cf, 32'hc43148d8, 32'hc4e57f55},
  {32'hc4150077, 32'h4502c94f, 32'h44c96351},
  {32'h4514171e, 32'hc25ceca2, 32'hc2ee9c3c},
  {32'h43682264, 32'hc35da1c5, 32'h44f3b3a4},
  {32'hc411d2a0, 32'hc49e62ac, 32'hc2ee19bc},
  {32'h43521451, 32'h432a33b5, 32'h42cb4e90},
  {32'h43e08c13, 32'h425ff890, 32'hc4a8dff7},
  {32'hc482f31f, 32'h43d60725, 32'h444fe96d},
  {32'hc4de53be, 32'hc299e4ce, 32'hc25d390a},
  {32'hc39ca91c, 32'h44f6a103, 32'h44eb2f98},
  {32'h452e14c6, 32'h437f6b5c, 32'hc3590c41},
  {32'h44aa35b9, 32'h4382efa8, 32'h4426d4cd},
  {32'h42f12750, 32'hc4cd0d57, 32'hc246c20b},
  {32'hc447af0c, 32'h446de9db, 32'hc1ef0d1e},
  {32'h44c3e743, 32'h4368c6b3, 32'hc338486b},
  {32'h43e94510, 32'h443d479e, 32'h441641be},
  {32'h448931fa, 32'hc4b54e65, 32'hc203c5df},
  {32'hc53c6ff7, 32'h42216304, 32'h42b6d103},
  {32'h44538e60, 32'hc398d5b3, 32'h44202e70},
  {32'hc5194e2e, 32'hc42a2c06, 32'hc14b433c},
  {32'h4578d324, 32'h430214ba, 32'h42c54ef6},
  {32'h443de50e, 32'hc4823b9a, 32'h448b877d},
  {32'hc34d81f8, 32'h43269120, 32'hc55549a1},
  {32'h454e4b58, 32'hc3886d56, 32'h43c12f00},
  {32'hc431be19, 32'h444f1a97, 32'hc4593a42},
  {32'hc41e8c30, 32'h450bb959, 32'h426004b6},
  {32'h44bd3105, 32'hc1a79745, 32'h43b53796},
  {32'hc41e4277, 32'h4514085a, 32'hc2c65bc2},
  {32'h44e9097d, 32'hc43bca00, 32'hc33f8e46},
  {32'hc506ba37, 32'hc2005514, 32'h424fb1c2},
  {32'h4446acec, 32'hc2eb82dc, 32'h445ee55e},
  {32'hc40d11c6, 32'h441fcac8, 32'h4435629c},
  {32'hc387c0b0, 32'hc40727ea, 32'hc38e733a},
  {32'h4415d5ec, 32'hc4381cdb, 32'hc40741d2},
  {32'h43c3bf5c, 32'h441490ec, 32'h45168d0b},
  {32'h452dadce, 32'h437199a6, 32'hc3b0bd03},
  {32'hc3aa549a, 32'h45033eaa, 32'hc284b5fd},
  {32'hc49c8362, 32'hc371d75e, 32'hc3018593},
  {32'hc4916cb6, 32'h44669e22, 32'h44a0ec02},
  {32'h4456bfde, 32'h43a72b95, 32'hc4a25242},
  {32'h44ac2c98, 32'hc3ae0fbc, 32'h434cd012},
  {32'h448c2dea, 32'hc43e4c7a, 32'hc35ab872},
  {32'hc44668b2, 32'h4471bc55, 32'h433fe887},
  {32'hc3bd7bd3, 32'hc386502d, 32'hc476e5bf},
  {32'hc23503e0, 32'h44384b82, 32'h455c2866},
  {32'h45082bb6, 32'hc3412d2d, 32'hc448209f},
  {32'h4532ad86, 32'hc2ea9523, 32'hc47abc0d},
  {32'hc4d3bb92, 32'hc0a094cb, 32'h44cccd2b},
  {32'hc256fec0, 32'h43b626fe, 32'h440279da},
  {32'hc4435e16, 32'hc4b0cdc5, 32'hc372463b},
  {32'h43811954, 32'h44e87904, 32'h4399caf3},
  {32'h4480241c, 32'hc36dede5, 32'hc41e8f71},
  {32'h44e4d1f8, 32'h44483473, 32'h431e0e6b},
  {32'hc43931b7, 32'hc5068d46, 32'h4181a4cf},
  {32'h44559708, 32'hc2054ea7, 32'h4322c513},
  {32'hc3fc710a, 32'hc3931c52, 32'h44b42626},
  {32'hc28320c0, 32'h43c0ffbb, 32'h442989ac},
  {32'hc3a219fc, 32'h4363d62c, 32'h4441e353},
  {32'h439602f0, 32'h448cb79f, 32'h43b1e3f9},
  {32'h43d4caec, 32'hc4211aeb, 32'hc422cc9c},
  {32'h44ade9fb, 32'h43803442, 32'h42db7478},
  {32'hc2a7e619, 32'hc4d10d5b, 32'h4338f16d},
  {32'h43403156, 32'h4424bde8, 32'h45236fd3},
  {32'h43c2e817, 32'hc416f15a, 32'hc429b573},
  {32'h4535886a, 32'hc37a1f2c, 32'h4479f6e6},
  {32'hc569f66e, 32'h43a3f297, 32'hc3469c4a},
  {32'h45262757, 32'hc31ba1f4, 32'hc3f47769},
  {32'hc3579888, 32'hc3ba02a5, 32'hc51319d2},
  {32'h4386a61a, 32'h450a51c7, 32'h445ed850},
  {32'hc208998e, 32'hc4b0e9c6, 32'h435b0e1a},
  {32'h4153d940, 32'h44f6c1fc, 32'h4431cfd9},
  {32'hc4ae4986, 32'h4292094b, 32'hc4efec0c},
  {32'h44a9dce1, 32'hc37b75fd, 32'h4371b32b},
  {32'h44264ce6, 32'h43a1e7dd, 32'hc3af40ee},
  {32'hc52d4538, 32'hc3deacc9, 32'h42b593ec},
  {32'h42cf4d50, 32'h44e23d5b, 32'hc3b82633},
  {32'hc3c2e5a5, 32'hc499f699, 32'h4413d69c},
  {32'h43fbb768, 32'h4504507e, 32'hc1ae6687},
  {32'hc2c64244, 32'hc550ec36, 32'h43ca6f2f},
  {32'h45346459, 32'h440020b1, 32'hc2d1eae8},
  {32'hc5127681, 32'hc439c0ae, 32'hc32ee429},
  {32'h4509a8cb, 32'h440b2d1d, 32'h4481dd37},
  {32'h4321ff00, 32'hc4811ee4, 32'hc2b93a1c},
  {32'h438f3d45, 32'h45108f81, 32'hc298af5c},
  {32'hc4bc6384, 32'hc32f615b, 32'hc3a56288},
  {32'hc4be05c7, 32'h440ee7c1, 32'hc16ba804},
  {32'hc5471cb3, 32'hc2e7fd12, 32'hc3452c44},
  {32'h445a85ce, 32'hc3935ae4, 32'hc3e530b0},
  {32'hc47711ed, 32'hc44cd28e, 32'hc355fc52},
  {32'h44b95da7, 32'h43781566, 32'hc46c5eb9},
  {32'hc5219244, 32'h41dbdc1e, 32'h43ae2618},
  {32'hc3a228dd, 32'h4407c289, 32'hc3bb62b8},
  {32'hc4d38c93, 32'hc491200b, 32'h444c2aaf},
  {32'h44606c6e, 32'hc33d8364, 32'h4376c1f4},
  {32'h44250987, 32'h44c21573, 32'hc3c9b532},
  {32'h419233e0, 32'hc536fdf6, 32'hc1f09457},
  {32'hc47bd306, 32'h42b5648e, 32'hc36a59f9},
  {32'hc5736641, 32'h43e8d8c0, 32'h433130c7},
  {32'h4467ec15, 32'h43a33cca, 32'hc4fd85e8},
  {32'hc52a76c7, 32'h43c83e79, 32'h42c5ede6},
  {32'hc46a64e6, 32'hc3bb2eba, 32'hc2559b1e},
  {32'hc430405f, 32'h45073410, 32'hc4067f25},
  {32'h44743950, 32'hc1a1c80a, 32'h43c6a77e},
  {32'hc4d3b225, 32'hc2a4be20, 32'hc3cc3073},
  {32'h454a8100, 32'hc29dd9e0, 32'hc4139f47},
  {32'hc4fd9465, 32'h435c6f36, 32'h4290064d},
  {32'hc49ac349, 32'hc3d98843, 32'h43ae89c0},
  {32'hc4c78de4, 32'h4406a877, 32'hc4a38114},
  {32'h451a3ec6, 32'h424b31c3, 32'h43f20db8},
  {32'hc49940c9, 32'h4356df79, 32'hc43e6a88},
  {32'h44acd296, 32'h434b22bb, 32'h448afac5},
  {32'hc4d7d825, 32'h441945c2, 32'hc44d5217},
  {32'h4420ebb7, 32'hc3d4b3c0, 32'h441463b4},
  {32'hc3adcce8, 32'hc39315d2, 32'hc46b0d5e},
  {32'h433b1fb1, 32'h43ad5008, 32'h4517588a},
  {32'h4185f080, 32'hc34038df, 32'hc4abcf5c},
  {32'h452cbe5c, 32'hc3b056a6, 32'hc35e4dbe},
  {32'hc477af40, 32'h4475c8b6, 32'hc486c084},
  {32'hc36ba85b, 32'hc3ade804, 32'h4427de07},
  {32'hc3eb5e92, 32'h43333191, 32'hc5434a72},
  {32'h4525dda4, 32'hc405221a, 32'hc24de20a},
  {32'h43fb635c, 32'h436fddbb, 32'hc44be5f1},
  {32'h4397280e, 32'h44af8d34, 32'h450ef25d},
  {32'hc50e77fd, 32'hc28dbf19, 32'hc4449bc2},
  {32'h44cb0f06, 32'h430f1517, 32'h424c4f6b},
  {32'hc38e5a3e, 32'h44c6451a, 32'hc4c6b072},
  {32'hc2da3ea0, 32'hc4bff0b9, 32'h4506bcdd},
  {32'h4424c994, 32'h444badae, 32'hc401f992},
  {32'h42a8fadc, 32'h43b795d9, 32'h435b1cc3},
  {32'h449ddbcd, 32'hc341be7c, 32'h44b5f59f},
  {32'hc3712bab, 32'h42ceb1d5, 32'hc4817ee5},
  {32'h4457d1f0, 32'h4358dedc, 32'h44849ca2},
  {32'hc3ad2c4d, 32'h452b6043, 32'h43b672f9},
  {32'h4336d8c0, 32'hc49fd79c, 32'h45082a68},
  {32'h447e12f5, 32'hc45c0f74, 32'h449338a5},
  {32'h43257d2f, 32'h448b1101, 32'hc5257c75},
  {32'hc354efae, 32'hc2350bb0, 32'h4332187d},
  {32'hc38a8580, 32'h438b7456, 32'h44a6cf83},
  {32'h43b12f5c, 32'h4330504b, 32'h44788679},
  {32'h44112e78, 32'h449dbcd9, 32'hc2b8bf23},
  {32'h4424b4f4, 32'hc0eb5a78, 32'h44fc2a73},
  {32'h4346fb48, 32'h44d75ca3, 32'hc42246fb},
  {32'hc4b3a1de, 32'hc25df720, 32'h439e7d7d},
  {32'hc54d7079, 32'h43e678f3, 32'hc399bb7a},
  {32'h42c837a0, 32'hc39eddfd, 32'hc3815b0f},
  {32'hc4e4474a, 32'hc342bfca, 32'hc38523ad},
  {32'h44a0eea0, 32'hc4878b4c, 32'h43bb51e8},
  {32'h43891460, 32'h44aebd5a, 32'h441c4da9},
  {32'h455cde57, 32'h435643fa, 32'h42944ff8},
  {32'hc505fd8b, 32'h43e05c5f, 32'hc2de8041},
  {32'h4463f3e9, 32'hc4e2d5b2, 32'hc365f19b},
  {32'hc460ac38, 32'h4432b369, 32'h43491960},
  {32'h4502b145, 32'h43dc0829, 32'hc37ea070},
  {32'hc2837fb0, 32'h43eff943, 32'h44c5049d},
  {32'hc38543c4, 32'hc4a2fcfa, 32'h43d533ae},
  {32'h451f4721, 32'hc3fccd0a, 32'hc2e62b36},
  {32'hc4727394, 32'hc3567209, 32'h4423a6fc},
  {32'h43fd9ffc, 32'h44cae1d7, 32'hc4814c00},
  {32'hc4e7ce83, 32'hc48e8fda, 32'h42af73ac},
  {32'hc47e05a2, 32'h44568fa3, 32'hc3603201},
  {32'h439ee1a7, 32'hc43aa682, 32'hc3a393a0},
  {32'hc48f6418, 32'h44b03dd2, 32'h44ab68a8},
  {32'h441df01c, 32'h446e9e1c, 32'h422fdee0},
  {32'hc368b4a8, 32'hc3b7ce68, 32'h44f62008},
  {32'h4464cf7d, 32'h4355820c, 32'hc3d1c531},
  {32'hc475034c, 32'hc41ef76a, 32'h43a94a18},
  {32'h42191324, 32'h447ec457, 32'hc4348011},
  {32'hc3d4023b, 32'hc4ad0919, 32'h4200a2d7},
  {32'h44c42e74, 32'h43ef46bf, 32'hc35b7416},
  {32'h44b2f9e0, 32'h42e65190, 32'hc3bc0386},
  {32'hc2ea43f8, 32'hc505e7a7, 32'hc3bf3899},
  {32'h45297ffa, 32'hc33b039e, 32'h41a97722},
  {32'h440372ae, 32'hc46a2a2e, 32'h435cc45e},
  {32'h4421435c, 32'h44c1dfa3, 32'h4430b35a},
  {32'hc46a8c62, 32'hc4c3d6a8, 32'h439f7ec6},
  {32'hc1d761cc, 32'h44d4b223, 32'hc333ed89},
  {32'h44358601, 32'hc1cea808, 32'hc35e8a66},
  {32'hc25a5f72, 32'h4311927f, 32'hc4a78bf9},
  {32'h42c7ea4c, 32'h44a0e02f, 32'h43cf4311},
  {32'h43d815df, 32'h43164032, 32'hc44f6354},
  {32'h44036dca, 32'h44f13477, 32'h445584b0},
  {32'hc3577729, 32'hc573b0c0, 32'hc2ba0cb0},
  {32'hc3abeac1, 32'h444f6ec5, 32'h43513220},
  {32'hc51f45b3, 32'h42790e9b, 32'hc3595dcf},
  {32'h44365883, 32'h43bf7242, 32'h44ecf454},
  {32'h43f3d8f1, 32'hc4d43e53, 32'h432fa080},
  {32'h427c7db0, 32'hc43c2b01, 32'h449b8da9},
  {32'hc33cf088, 32'hc4d5644b, 32'hc3e099b6},
  {32'h442d970f, 32'h429009bb, 32'h437d45d8},
  {32'hc3711ef4, 32'hc331d356, 32'hc545f448},
  {32'h4427c152, 32'h456855b7, 32'hc349ac2a},
  {32'hc4d7173e, 32'hc3145acf, 32'hc2d3bcfa},
  {32'hc3820054, 32'h43a3a188, 32'h4510c48d},
  {32'hc33851ee, 32'hc4d29f3b, 32'hc4a9a46e},
  {32'h452413e0, 32'hc34f535d, 32'h42e07e42},
  {32'hc529ec97, 32'hc470e291, 32'hc410d0cd},
  {32'h452dacf2, 32'h44ac429a, 32'h43e8ae2e},
  {32'hc4d5a9e4, 32'h43c40650, 32'h42bc982d},
  {32'h422cdc98, 32'h452bd507, 32'hc3774b8e},
  {32'hc4d4f204, 32'hc498f2d8, 32'h43aef27f},
  {32'hc38bdfcc, 32'hc361ccd4, 32'hc2d85c52},
  {32'hc4326d42, 32'hc31b8062, 32'hc318a67b},
  {32'h450cc3d3, 32'h43876472, 32'h444b3da5},
  {32'h417016fc, 32'h43a7a9ca, 32'hc4b9c812},
  {32'h422dcc6f, 32'h44834ffc, 32'hc41b4dd6},
  {32'hc3f8e668, 32'h43b36fd0, 32'hc27da94b},
  {32'h437c6a3a, 32'hc3af2ecd, 32'hc3de0d4a},
  {32'hc489bf23, 32'h442ff607, 32'h43d8a67f},
  {32'h44d1b6d1, 32'h43b66b27, 32'hc417cfb6},
  {32'hc50083e0, 32'h43d67a7f, 32'h448468c8},
  {32'hc4f1c734, 32'hc3cfabdf, 32'hc22b3118},
  {32'hc2b1ff23, 32'h42441d41, 32'h440c5192},
  {32'hc43d734d, 32'h44ad97d3, 32'hc51d32b2},
  {32'hc3cab8c5, 32'h4424f41a, 32'h441688e3},
  {32'hc398bc6c, 32'hc49f8be4, 32'hc41704a1},
  {32'hc3e941a5, 32'h44b0ce2e, 32'h439ed6ee},
  {32'h44dea412, 32'h43c2bfca, 32'h42010bfc},
  {32'hc520269c, 32'h42d792c9, 32'h43406900},
  {32'h4449d65c, 32'h43b542f3, 32'hc2c9b322},
  {32'hc4a2de7e, 32'h444b6ea0, 32'hc1409c10},
  {32'h44a5cc93, 32'hc49318bc, 32'h436700db},
  {32'hc50f9c8a, 32'h4461c2a9, 32'hc39ab10a},
  {32'h44b69b00, 32'hc318b030, 32'hc3afe992},
  {32'h4210dfe0, 32'h4582eb91, 32'hc2391ff2},
  {32'h44634e4c, 32'hc4ad9205, 32'hc28c837e},
  {32'h450fd621, 32'hc2767b23, 32'hc2fc637d},
  {32'h450110d2, 32'h4403d77f, 32'h43cbd1de},
  {32'hc50b4920, 32'hc3eab0ae, 32'h43195ba6},
  {32'h455cf1c1, 32'hc28a01f8, 32'h43d7521e},
  {32'h442bcba3, 32'h42b8b6bc, 32'h44949e09},
  {32'hc58d56f5, 32'hc3b7b7c5, 32'hc264a397},
  {32'h40f01500, 32'h429fbc00, 32'h45275cf1},
  {32'hc437c18b, 32'h435dc9d0, 32'hc3e26525},
  {32'hc4bb20da, 32'h445f89ec, 32'h442c6a2a},
  {32'hc36163c4, 32'hc4b2c62b, 32'h41bfc6fc},
  {32'hc430ed08, 32'h44ae423c, 32'h4322c20c},
  {32'h44f3b641, 32'hc3ecb0d1, 32'h42bec48c},
  {32'hc39a536c, 32'h42d9f3b2, 32'hc3c68375},
  {32'h44ee1711, 32'h43b00071, 32'hc37fd5f4},
  {32'hc515ff19, 32'hc23e6442, 32'hc2161b0e},
  {32'hc3b96ff4, 32'hc2e450e6, 32'hc4322f56},
  {32'h44028392, 32'hc43e807e, 32'hc31ba93f},
  {32'hc4750c12, 32'h4281a30c, 32'h43a78e02},
  {32'hc3db6e49, 32'hc41f61f0, 32'hc4760af0},
  {32'hc3052d1a, 32'h44ba7985, 32'h441c0239},
  {32'hc41d7861, 32'hc41f4712, 32'hc2f2d4b9},
  {32'hc411dd40, 32'hc458fd1e, 32'h4452bf1f},
  {32'h427524b5, 32'h4442802c, 32'hc4cac1ee},
  {32'h4368ded9, 32'h4397823a, 32'h450236d2},
  {32'h44964a5b, 32'hc4812359, 32'hc3b40d99},
  {32'hc264da84, 32'hc487458f, 32'hc3165b8f},
  {32'hc4a2939d, 32'h4387f9fa, 32'h4484180c},
  {32'h42380aaa, 32'hc49bfa38, 32'hc48f162f},
  {32'h44ee2932, 32'hc2c45ec9, 32'hc4e9025e},
  {32'hc5061794, 32'hc3708233, 32'h4501ef20},
  {32'h44879b30, 32'hc0b682f8, 32'h443dd31b},
  {32'hc461c35b, 32'hc4eca770, 32'hc3228d23},
  {32'h45058092, 32'h43f0db55, 32'h442c5f02},
  {32'h44f0013d, 32'h421ddff6, 32'hc35709bd},
  {32'hc30c2cb0, 32'h457588bd, 32'hc4006d5e},
  {32'hc470dab8, 32'hc4f3d797, 32'h436729cf},
  {32'h4441e79a, 32'h41d9afa1, 32'h441cf691},
  {32'h41e5c678, 32'h4430f93d, 32'hc4f831e9},
  {32'h4405c3ee, 32'hc39fb514, 32'h434ea816},
  {32'h44bacd64, 32'hc38b1547, 32'h42bc1d66},
  {32'h451b9d54, 32'h44088efe, 32'h435485c1},
  {32'hc41b0ccb, 32'hc417e6b7, 32'hc5434de2},
  {32'hc43438f8, 32'h42ac8656, 32'hc18061f0},
  {32'h41ba0080, 32'hc48b0de1, 32'hc4154501},
  {32'h43ef45c9, 32'h451fa6a6, 32'h44344b89},
  {32'hc1ee9140, 32'hc28e46a9, 32'h43c6883d},
  {32'h452a9197, 32'h4418f4bc, 32'h44185f94},
  {32'hc573d1e8, 32'h43953b86, 32'hc2ff87da},
  {32'h4543bc3e, 32'h4383cdf9, 32'hc3d594b0},
  {32'hc3b5a328, 32'hc2cb5c29, 32'hc522733f},
  {32'hc31ee336, 32'hc3889b2c, 32'h45156abc},
  {32'h44a71fc5, 32'hc2b90448, 32'h42debaf0},
  {32'h4393b2e8, 32'h44c678ca, 32'h44bf6b54},
  {32'hc458a97e, 32'hc4eab7bf, 32'hc3691c52},
  {32'h438aca5e, 32'h43d56529, 32'h4199f13c},
  {32'h44b6d020, 32'hc46beaa9, 32'h434718d2},
  {32'hc387120b, 32'hc5254c0a, 32'hc4027c1d},
  {32'h45018355, 32'h43060faf, 32'h440f8071},
  {32'h43690b01, 32'hc3d31d21, 32'hc35f91f2},
  {32'hc287b5e8, 32'hc56a88a3, 32'hc32be267},
  {32'h44a1510d, 32'h43423b6b, 32'hc3ae7562},
  {32'hc4a66ceb, 32'hc3c2dc52, 32'h43706d13},
  {32'h4551e11d, 32'h445cab29, 32'h443c85ba},
  {32'h429432c0, 32'h43bbc6dd, 32'h44ef9a77},
  {32'h43aad956, 32'hc4153b4b, 32'h4450808a},
  {32'hc3cbd74c, 32'hc45b8984, 32'h44c69209},
  {32'h43073896, 32'h44c38ad9, 32'h43542763},
  {32'hc4e10898, 32'hc3f8247e, 32'h43edbeb5},
  {32'h44274811, 32'h452ef3e1, 32'hc2899432},
  {32'h44b2e33c, 32'hc3c4b329, 32'h43d26660},
  {32'h435d2816, 32'hc35dda02, 32'hc52b7cfd},
  {32'hc4bddabc, 32'h43d795b7, 32'h42fe8588},
  {32'h446649be, 32'h44519e79, 32'hc3b94709},
  {32'hc3169a7c, 32'hc51a31cf, 32'h430d1ca0},
  {32'h43153f42, 32'hc2586549, 32'h44de4fc8},
  {32'h43ddbc5d, 32'h450ce94a, 32'hc394c406},
  {32'hc4379b4c, 32'hc4c559cb, 32'h4340bb39},
  {32'h440d2394, 32'hc0bf1fdf, 32'hc3e68a94},
  {32'hc518564a, 32'h42bab5db, 32'h41ba2287},
  {32'h452e2159, 32'hc30a9d6b, 32'hc444d9a5},
  {32'hc3a735f0, 32'h442b332e, 32'h43c26d39},
  {32'hc4aa76f3, 32'h43402d5c, 32'hc1646a4e},
  {32'hc3103188, 32'h415c348e, 32'h4357d0a7},
  {32'h4479d045, 32'hc4bcaea7, 32'hc3b31a63},
  {32'hc3fcdb06, 32'h4486a7b5, 32'h436baeea},
  {32'h4504d9b4, 32'h4330e4b1, 32'h429aa833},
  {32'hc3771fbc, 32'h4468304c, 32'h446a683c},
  {32'h44cfd91c, 32'hc2b547cc, 32'h43fc3870},
  {32'hc4864254, 32'h449cc404, 32'hc2e2e37d},
  {32'h45033ef1, 32'h43d51933, 32'hc1dbe70f},
  {32'h43c21e28, 32'h4390e1bc, 32'h43c7a127},
  {32'h43c109ba, 32'hc517e212, 32'hc2b728fb},
  {32'hc409dffe, 32'h44aa5ba6, 32'hc2ad500c},
  {32'h44348094, 32'hc3be7505, 32'h43bdd600},
  {32'hc51493d7, 32'h43039f5c, 32'hc4254b6b},
  {32'h441568de, 32'hc43c38cd, 32'h441d93d0},
  {32'h44b37b76, 32'h42eb7816, 32'hc437fbf7},
  {32'h4471cb97, 32'hc4b26b8e, 32'h4388c433},
  {32'hc499b81c, 32'h449a9b08, 32'hc3a5ccb8},
  {32'h411d3750, 32'hc3cf2215, 32'h431958f8},
  {32'hc383f9e3, 32'h447e5abc, 32'hc4dad175},
  {32'h43892a48, 32'hc32b1d1b, 32'h44e5b214},
  {32'h4438d780, 32'h44a1355b, 32'h440528a8},
  {32'h438ea844, 32'h433e7545, 32'h451fc6df},
  {32'hc4cbb562, 32'hc3f123c6, 32'hc4c585fa},
  {32'h4511f0be, 32'h43d467a7, 32'hc3639212},
  {32'hc4574a7a, 32'h442b22ff, 32'hc44bfaac},
  {32'h43eed568, 32'h44404a5b, 32'h44d9dd64},
  {32'h43bd9705, 32'h448a517e, 32'hc4b39631},
  {32'hc3c0bf97, 32'h43b25a8f, 32'hc42393d6},
  {32'h447b7fb8, 32'hc469ca13, 32'hc0e0cf2a},
  {32'hc4016642, 32'h44a67fc1, 32'hc3469fc2},
  {32'hc38c2654, 32'hc1d7f263, 32'h43a0e9a4},
  {32'h42aa12b0, 32'h44f38766, 32'hc43fe00a},
  {32'h44f5c756, 32'hc41764ed, 32'h4408df47},
  {32'h43470569, 32'hc42fc447, 32'h45013935},
  {32'hc3498f7d, 32'h44f94e42, 32'hc4a9d392},
  {32'hc4894c1b, 32'hbfd90617, 32'h43ef2952},
  {32'h43368880, 32'hc4311730, 32'h428066b4},
  {32'h43a65c70, 32'hc4cb42eb, 32'h43006707},
  {32'hc528edc8, 32'hc3c5267c, 32'h43a6cff8},
  {32'h4467a872, 32'h428c663f, 32'h442af787},
  {32'hc4539d98, 32'hc2b155f4, 32'hc469b9d1},
  {32'h454f97cb, 32'hc3aea132, 32'h43afdfc6},
  {32'hc51f455a, 32'h43d00250, 32'hc31e607d},
  {32'h427dd340, 32'h445bc1ee, 32'h43e17e0f},
  {32'hc507459d, 32'hc3209a57, 32'hc37f12bb},
  {32'h4296dd60, 32'hc458f091, 32'h43aa6332},
  {32'hc518f361, 32'h436aecc4, 32'hc3807f32},
  {32'hc38f353a, 32'hc29be5bf, 32'h43a803fc},
  {32'hc4a18c42, 32'h45017afe, 32'h435a275d},
  {32'h450c3fc0, 32'hc48a4405, 32'h4213eb46},
  {32'h440a931e, 32'hc465bddd, 32'h44a28bea},
  {32'h43862355, 32'h4329eb65, 32'hc4dada17},
  {32'h41d34e80, 32'h44b2181a, 32'h4493aaf9},
  {32'hc460441a, 32'hc43f06da, 32'h4407f8f5},
  {32'hc2cdfda5, 32'h44b7e428, 32'hc1bc923c},
  {32'h4291e7ae, 32'hc40a6ca0, 32'h43cb2c01},
  {32'h4481529d, 32'h44a771af, 32'h439aa79f},
  {32'hc40662f8, 32'hc32970d0, 32'h44e386d0},
  {32'h436c595e, 32'hc2f6a33f, 32'hc4c064e5},
  {32'h43851afe, 32'hc4385270, 32'hc4b8fe17},
  {32'h437c7ab8, 32'hc50983c1, 32'h45017af4},
  {32'h4425fc08, 32'h44516721, 32'hc4277896},
  {32'hc25a5b58, 32'hc55278ff, 32'hc3d14248},
  {32'h438b5f2f, 32'h44d23e1a, 32'h42f9fa78},
  {32'hc2b6882c, 32'hc53473f5, 32'hc403c2f6},
  {32'h4328e0ea, 32'h44c3ba7c, 32'hc42a0a20},
  {32'hc37329fc, 32'hc4ade738, 32'h41d48b89},
  {32'h42de3c00, 32'hc42c9809, 32'hc422fc38},
  {32'hc477d5bd, 32'h43e4caa2, 32'hc3a152a5},
  {32'hc4ee9f4b, 32'h43a85e0b, 32'hc217db37},
  {32'h457a1372, 32'h445e5eac, 32'h4202e622},
  {32'hc518774e, 32'h42643880, 32'h43b05d91},
  {32'hc3eb0d03, 32'h454416a4, 32'h4417cf73},
  {32'hc4ae4339, 32'hc4923e44, 32'h42761b5a},
  {32'hc47ff7ec, 32'hc337ef8a, 32'hc32b1486},
  {32'h43f09add, 32'hc4b01d78, 32'h421245ef},
  {32'h439e7f9a, 32'h449ff243, 32'hc503052e},
  {32'hc35d175a, 32'hc4c6abff, 32'h44bc5a68},
  {32'hc498b358, 32'hc2f33f8b, 32'hc36ca849},
  {32'hc1b1576e, 32'h45512eff, 32'h41f181d2},
  {32'hc4f87b59, 32'hc4458366, 32'h439919b0},
  {32'h448bdd8f, 32'h44667f5a, 32'h4199d324},
  {32'hc401ae3c, 32'hc4d6b08c, 32'hc4d58449},
  {32'hc3ce8203, 32'h43b4ec2e, 32'h44fe7416},
  {32'hc3179c44, 32'h44a8e790, 32'hc481ee34},
  {32'h44b956f1, 32'h43613016, 32'hc2f99e2c},
  {32'hc412cb1c, 32'hc3e2f2b5, 32'hc44e3336},
  {32'h4393645d, 32'h43ef30b1, 32'h4035523c},
  {32'h43ab1db1, 32'hc4ba80aa, 32'hc34a2a7d},
  {32'h4519acb7, 32'h40130da0, 32'hc3ddc5e8},
  {32'hc5025a9e, 32'hc392aa8d, 32'h432ee98b},
  {32'h44b5f015, 32'h43ece6e9, 32'h438d88f9},
  {32'h43bf2a74, 32'hc3696903, 32'hc51eef93},
  {32'h4422d9b1, 32'h442e6b86, 32'h43e47385},
  {32'hc3e7777c, 32'hc50684dc, 32'hc2591153},
  {32'hc3ca2086, 32'h456c2f14, 32'h43cf4880},
  {32'h44a20e17, 32'hc3a7fd73, 32'hc3b93e47},
  {32'h4506dc37, 32'h4430e6bf, 32'h43d8da96},
  {32'hc4448817, 32'hc37e2a4d, 32'hc3916662},
  {32'hc44f9120, 32'hc2b4347d, 32'h43360d24},
  {32'h43d23410, 32'hc40e1f81, 32'h43c95c56},
  {32'h43e2ea6f, 32'h44bb1cea, 32'hc4800353},
  {32'h43ea1d5a, 32'hc3490281, 32'hc2a72dc9},
  {32'h43b62f6f, 32'h44d2e5a4, 32'h44962b55},
  {32'h43a92d10, 32'hc402828f, 32'hc48fa9dd},
  {32'hc3bc1eb6, 32'h4486d642, 32'h449076c7},
  {32'h447e78b8, 32'h4264fb1a, 32'hc4c01830},
  {32'h41f56e40, 32'h44b239a6, 32'h44ef81fd},
  {32'hc4ab5b36, 32'hc39e2795, 32'h4313bf21},
  {32'h43666e4c, 32'hc1c7c4cc, 32'h447b111f},
  {32'hc39fb8a7, 32'h443f0ca2, 32'hc51aad3c},
  {32'h43a2a5e4, 32'hc399eb93, 32'h43fa71b0},
  {32'h42eb5940, 32'hc2e2f710, 32'h40596f74},
  {32'hc45bceac, 32'h44afef95, 32'h436fd13d},
  {32'h44ac3f7e, 32'h430fa6a2, 32'hc3f1f6db},
  {32'hc4d81552, 32'h435b1a01, 32'h43dabaa2},
  {32'hc1ce1e80, 32'hc30a702f, 32'hc444d93f},
  {32'hc496662e, 32'h43a1509e, 32'h4216f6a2},
  {32'h42949854, 32'hc4505bb1, 32'h4300e97f},
  {32'hc3320902, 32'h4557a14e, 32'hc3117e65},
  {32'hc44e76df, 32'hc2b93205, 32'h43e3997b},
  {32'hc3962478, 32'h448bd8fc, 32'hc2a4c047},
  {32'h4485d478, 32'hc5068567, 32'h440cfea7},
  {32'hc502038d, 32'hc360a7be, 32'h431a4682},
  {32'h43e71fa8, 32'hc3c97d6e, 32'hc41081c5},
  {32'hc57b27f7, 32'hc3d92b9a, 32'hc1ef68fc},
  {32'h45372678, 32'h42dd0df4, 32'h4150fbf0}};
