-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
J4urr+tPku3zOKlAX75XVzV9yviS0lVc4LcfpRob60gekOWc1Xqx5nlvN5rd6gYO
0/1+0yQ+PZFINGuNOON5RCcAifyXojEBpBHiEFF37OjpSptpeteS7PzmUCpD9zZf
qZ2NuL3yIOecNq2pwRUK35eyqKowSMQtyX7XPOWDWUdqhu+Ob3quUg==
--pragma protect end_key_block
--pragma protect digest_block
zWeftGoHJum1WqsmBuBz8bNOcdo=
--pragma protect end_digest_block
--pragma protect data_block
K4KT0QFpAbmUlCucxMpLK+aV+FdhAd6C1loAxSYTJ9tqofPYBew5B8uoL4YCqP6b
JSF3MwS4cgxLdlaPo8ViUP+YQRS0BzODMB+F5VZ3+WeGLYkbgkYTB914UWVeYzml
vMMdWz6S2Gq2O16kcSxb7iNzYeg4jThvFFHpY3PYeiy0VDximgMmTVkXZ7OmUAop
StOfSUp6rz8c+Y+0sSYZ+uGxWozuFwsbGoFeLJ0MJafoK7Y3x6M7hCaQcmn0uwOF
94aHlsOM2a5gWid3As3rZRVa7NiDXpZFPbPoONS5BaYCJ669P/9v5+1+FT7ObNaK
ggN1y7bc8hAamvsXUwcdy0KJw3osBoA0tTYq+GzbRIX3j/UWopw+E+dq5Lv7/C0o
dHwx1y4xfwrbtAZNuy9ww1j6wOD+fjHUfvVqILMvoZuXOe6KsP/fyKVpOXC6giw7
P6Np2oU3r4ISm6G4U4qOm8MXa/LhTr5SCGHwBU8PAxgr9EYTLcOQdFkQCB/qc09m
Kbd2oqrFstIK+bdzKYSW+t7ui5h61FIAQjCQSJY9X3tqtaAmSEmVh4q4E+j3PhGl
/gmEDBws26EVAPttQomCs68NSjWR553llYz6RxPZxE2SaJiMMYOEQkcvkIgTlxXd
XWiVRWpDxi/kT6wg2VVMVPlD4jWKDLCZkuKExnr+oXvhi6LBB0X+aULTaTXmYL3m
kz3ssiNIt7tm7oKUiLJ+qGYBYE4fWqcacFml+JGSCdFfDl1vRPnBxpcjEF4m5C7n
8H7L8JlFw76/5g8mKscVMnwEuTbUIXJ/XrBi6NCySPHX8nxlD97pObbFLkuZd69I
0QwueVtWSOvFsvheg/BZ36jSrcS4I2OhfCCYwWUnFXMCxlVw249XiUoY/TrADHp+
gKsPT6bmj6E27io05Urbs2ZctjPZy3uP6+K6XpLSAEilB+rQfGvVLT7Uc9nWqa1k
UH9whLkGIjf4c1qCRbqPFYj7USIcgImqPu6OyBdWcWad3SISe8fE5eY+xwpE9b2t
MpE+g3CkL+pSijM3m5e2s3kaMdB3r2Y2hLUI7Ac8C5/TCtB3tzJtX6P87lDYM3nn
Ul1KytIzFcxAjWThR6BU0dB9jlFiTSkfnS+eC/en9jROWMaxB5n+DvUv5DXyyT9X
xfhj1bjxz0OSZAJ62pvy2+7U6B9JcmmveP9HitQZqxrpjfR6Ivw3LzovhCSLcdqp
2F4cdCiSTSQSvzB9T0nVzVXELLfbhkr4mrDUnKEs8so5LIbIVyGDfRyKR62Esivt
ZjOmyLNNuauwV67w1W1KxIJBU7Ql0hXBvAYX+UUbmWvS36bn7wCyt1mg8jeSVJ9y
zpxPn0fBtl7Nl2rOejfh9w2ejZDnb9gXioEkoSRSSuPEYWEnm4iylx2ZMoys33rl
LbIx88CTYjq2/p4FgdVjdbLrlAz3BI6jHxNlRMfP6hCgLJwV59zjo69KZSbgLdon
6wa98Co3Toc1pYBAHrW69Fh0ivTpn1C10jvSj2T6/uR4wzeTag4li+xagY2NUied
A4Oo+JH4Q89SFTey0g3GN9XCcrDcPVglOGSPXPZt1elXQ36e3kCi5/9Ud/YseviB
r607EUtcniEqKXpQPqaDyro6cadSicD9MeE7h/nEI7TBF9d8G9zKoEyojuzkUq6C
wltJVM2BerDxf6e/6v6gabNIpB7dHMzpi8mFa1pBxbKhN87wTsyJvA1PcQbrK12g
Xpy9AV6mRxK37zhmtaF+OZplEG9pca8k41x6624TTpuZTeNvC53CSB0hkaruCkXy
N1v+m0FykE+dAP3SyJ3TVR/1f7SwWG8B1c747h/JNjoq3AkjFinDxVr0roXsdWCr
kOkJx6e1lPSByhDzzcWixz9l6THkILOUfZx5/HK1SjRs9t1aAEfjtNsBfl3sxXj+
rK/pySLIcykAlPOFtVeokbKywn+vpR9Vht8rvH7Bc9TsTMCaymwRfEqFxbsjBirF
//VIzqQD3EJGJLmDlKs9111m5tYITWH+bYjxLidKEGqt0saOx59a5+uOfP+4wxMe
e5q6c9qnTgXGFexq9vQ1MmczsL7m2EgkeaGdaiUsH6hY0ZmLDPl7OqnG8WYHFbou
KrW/YuawDwKw6i7S8XlLvpsvRoFyn6rDqVchB44OAF5z1+UG/hxjyyGHzAdlAK2E
jxIo/sRQvDNxdFjBhyqWV4app/t5A+jE22g4yhOM2V9v+hNa2zDRDtOOOkqfFuGA
MRS2clMBT4dH6m0uAz5i9Aun0iOj4PkorfLleGhTUe3L0vU2Ysm2C1Zbj41OhqBL
bif0klPLVEdptprIFclRc2dZuRHpf2OlBaEtDSbyAB2ddw/i90atu0l3mHOAXyOn
+c2QNcsDKHm/UqlGB+HCcPBnO2tph2pC6lkroMaLpV7CYLrThLRdl19FTtE98vVI
Edn4/XG6nq5kWm0F6/CM4YnAcV0+coQ/L6HWPFKG8pAwhhXZaSz1rvp2UUo7531O
YpqVnZ+ifzCS7eH86n/isGAN8p2yULQWl9hIXFTW5hd1AH5fXHNpXWbGHZsBrKLQ
7uvI4S6wJdHfnsxPUKQmgeWCQs6NFPlYG0qE47WJe1qC33ojce7Pc1ga4+gGMDTl
WDNNiVySTvkKnyLu21iyb9g8lozAtOLpNqfN+43APi2GEndekt2xRcq9UOggwIhD
ehalnZJiXePhglutF2WldXbDSNjrh2gutXu+KF26M5k18x7GU45iB6k3LGt3n8uc
mW1ciJVuIvhqZDwiamqLQwZ0wT61lgLRPFLb3np7BVTHf029ECQ3m0U3/vBrVDUV
Ompd3MzZ8UeMjd9NW7eFVJxDx91s8Nwi96V2pS6f57+NwoEZ/mQHG7Ya5+x/Jogu
bEPOydbXeW2cin+wV8m0E/VL0hon3jTTlitRYeFLQUAfFeMI5pCFUAo6jDKorXA8
lSSA8BWMP+87FPRZxKt0r16F+2+HnfHbqe+Qw021xIgeQ9ZTbpaGYT0lTMg+xwe7
yg6UTvFtXm3tKMYWpRjRt56T2AqNjJpI8HWMfbrmLfsQ2s4RgV+tIvGxeHbcPnLf
2jNDXzi0T4VTOXNyIbik5uTociAR+v3YQaVp52ZVlvewL09O5/yfcN+ZxwO/h1qS
WI7oj/IIxKSpm1qXBvM0mxJTI8KNJwX0KI4F3hXuJ07/rt4cnwycXuiLugkvu1Lo
PFHZ8rDDhG1wSKrYAwORTIA0Y+P67xXP1vJqGEhVa346cXGrGll9U4INJF8DO6Qm
Bo3ii7fX7DLqGbZ7/ikeZenrB7MfnRfnfPi+JotYP00PgAPuifji4S7jYzgYBInW
SaeugF6qdvld76isKXnkXTL1NlgcvdK0GDkrMu+RGxCPYifouNdHhlxON4X21HwZ
Zg7fplZkzk6HCYvcjm6XY9n6LDIOGuqn+5MYebt0t6ZDTAM2TUnzWTCaT9I/AVip
PwDysAzoO+zJKkm9SUeMxswmM5c8xg7UCwZQkm6DLqXPnuLqdByh59ijST8j7fnr
aQOcO5O9a911uA/stIZwnj4BEWbk0Ca9dm78uDkbmg7u2O4lv7YyuX3pq23ht3eF
HU/RtoENa0FTBjRtmIQr3TRls8jtgsolu9BdUrFOkVoxcknCLqrje+urdg8/Lltj
g9dF+lTPzLVvAOgLoTcANzTclASiG4XK+fv+aunyE2h9Qq6z/r7kYj/v/GkMg15D
7LJyTl7MRMUo37Lu2+xnjKFQ6idu8vqvMRLnyFOYwKW0rOlnj0ul9eaZgzFWHJEb
Hv/GeMdUL//huSxVSPlQ3eE27RCjkhGOE0Cc+IS6m83VmTNx3h7wl+VtEX94/i8e
D6LuZegWPPxGR5jJ0pgGXC5EKV4oYngpQhalu/yPRTneUdeh67gGvyRfSZwOdLif
JcuLc1g2PJWBJuK9aEegGxhtHCnhRfhvf4WqjS9esRUcYlxzi9S1TAYhFfWnNFOx
cI0eextSMH6T7n7xRjxfcvw+Eo58cWsbp/wSPZzXUOcakJbGFAmfuCSiUt/12rNq
Xy2mpqq0sdubJq56lXlPyAGb5T8Kgtl78ynXersH7BHJwyRTJ9hXrN22Nd7hMI5g
G8b9zNYycMK6roWdOBdytC3pu3B+Ty9nhoxb1A96r1ZigdX6Lwm+86oXkd3S7c5o
fzR7YXT3Uh1Lvm2/CjGlnjZgdtX1+Tf984V2DQvP3x7w+q4+NJTrP266VXC8ZOuU
vFLKXz4WgSbuUWEF99A2RH0BzdguAv8S8JsJc7mCwCU9VFpyHMW+/HMI2jFuRyh4
BllzFPl5J5cz3TzogDmRtXUkUU3MrjnY5mJqiJ6exrJQtKRol262pN77EivSn4Sy
alF1D2BHDiUrWuCfL68A9JsYCwhV7WmGsCJEy0qy9wCUBcr4TgO3pNV56uHh9moY
81cQd/wxlmqOinBB3+cZTatR5d41Sa+iNJg4HyLYfkERUXWhE0vnFT2LgY/+2LRi
7DAyTHDGCFPZ1sG2RmHFdX3GW7e2Bhk6V5KyOosozxVNtHA7Aswe95BWcbpSJy5s
daZFzvEZHDi4ngXE514aTaS0n8jwNZO/es7YBqMekv1OrwnnK8sS/G8vDjNdLzaY
N6TOwX7c8x6fEIf2Mr7R3WiUPK3hUS8GihYVlvCoXIWIORbtXiZ7flHanFCi/Jum
vUY5TXIHM7pfp3DMeuZ2w6B4Ml44DBptCd+oW/Ms7hLHIvmVZ3YrhUjPUCAhemiN
lLiX6UpfRLZg67bJz+mA0lfKwC7yAGPycvyTNbNIxZw+sMsNTi3H7OOug9Kww8F9
nWdkLeX1uBQR8cx/oUM2NCxSw2QA57/gu6hcOZQi0mK3XPX734N2j+/FtmGJdJjn
0GxWDlaGqnnj9tATm7EGa8Wayn94u0yCFHRq9UnUBTgpsU9d9XERjm0W2+iuEK3G
CD4rBoekVTTAu9WInyFxjvr/C0gnWV0RsRYa+aYSBPg0sKfYH/24wtc6qwH7a/iF
OC4FUSOpFvbG3oZWEw5dZd10vxTfd0LHafjSEhNGj2u4MIF2jiojH6quLdjDrXZE
Jefl/QJ6OzxGzwPhw2r47PZQWB75eMIKijdL+nlnHiwFW2A4BXe//GcMyocd8hC3
3O26gRBWAiH5OtzRgzvIw3ibooyG56+DBbj2HsW7B9+bVE6wzBDy8m7qd4LMIkUr
84Ny2/zjygSEf+1fZD0QVOvMUmurkEMKLqmayv+6HgyljpX7AYX7CkqmBW8JkU9s
+n1h0bpVkZqH+n2+sSBphZ5WtqoI9MrWVgp5JtCEqVB73682WENfW0LhJ2zTLOJj
ltNdhTKk7uNfKjfc0V7S+sdQavwPNQuGjr/kfsRRSJidO90x//W4CNXIm+7+rdho
eLyNprOWuRF0BmcG/wjmnqqTjLpr2l+6pfbsd9I7rCXoYIJ53Fw1ZoIfTUfAmGo/
biZEFKQ8JeAWXLPLgd3wGmvyBgAb08TstSJK4nTWwmo6IYY3EmUfY1cTQAptsXZ1
Y8MIKMXQor6YvFu8T44J0Laj6xb/9VCiQKr2N+8u41zNpbJH0D/drvbM3SB3Wp0O
1hp+GdnUADG9Vv1wcpOZQTVy6eTpJWOJNs7ZSoe+A6hffhBIQsziMnTLGbxHI5xY
ReHsUo/Yv9hPKZyUsNzr+R7qjY43+7O8JjCn+jNLs5U4SXndQ2+dIM3Jkq36IBB2
sv10wUsfKdXYOcQXEA8GZRO1u49GIWX1awa9BSZSLBUnQlhTIyzJ/eI1lOpqTrEc
2Rjy6Ej+xP9Wk5wMV3wxG2xhUdPrQRp1ANX8+ROcpbVSwc5XU0E7u9NfImG2z128
OTI9Mn+A/ht8GTq1yznmiKZ6xyVqG+qJRx0sVX02CSWtVlsGgVYGcIYYLEGzYTgS
bVMV0VE1Si764XTOBbaWctjeunZcsoyxzaia+b6pMvn7cNpE4fW5eazqZz5j3B8d
89mgbMCT0Jc2xVqjmInZdmrstufX4P+Vf2jb5DzHcTlJyaJOavzGdH05JM2UV5mR
LhOPNiV/RUvjz5WbvHF0qJHucUWC/qxf7dlm5Sv/lxK50cvIDJOjiRvtVZITaiWq
lQbwZcjjSU88mwiPTOl92JhqcOb1MXJit2OlZYw8rz+0N8Ia+EOYvlO15RgZxeY6
itqJpMS9eDYJ4eogpfl61rCjGX1b7m3OI1WkR4dXnMcmat0rihuqnilOTpLug8l5
Ijs6zHLBAKqC6yyqZu+I4leIXVdkfCsaATCTfR/B4UIZEsvTBKtchSXsZ+FSV0T3
vFMvfQUTXG6XHYyIsOs1uLkrvW1KPuouoDSpQcu7407ipLI8K7K1Zk7TH3DPp8Tb
bQgBp7z4SL/000OosifC3FIzRHnOrjwjeiOpljP5RG0RGRkoYJUpYriZ8v+OuONc
cDwWQ7up1ixJLaqK065Yq2whz0d1mJoQJ/x5214vnbwdM1Pv0W03VNhq+nBPa7WZ
2h9b6a0wFJFRrlwyp4q2on5Ynh+5aE6a6K8In8U6xKKBYj6iRCsGDH0UPUq1Q5mn
uBrdIyG8KZT3hXjWGbrz7gvFAiP8ihesdTM1z4VI/S6botVqPg8W/4thk0Z1Lm+d
RbnS5hAJg4H4U4NQ/7i89ntiyKIyf7V2I+LjJ4NRolQjXH/uxGvZ2tJQcejK90NR
KYtBxeLPjy7QIq0qXXAMKQ93zWkfC/JbfO2vGlN1iR7BUcc5IRHjZL426j1rVQqJ
N6gTWry1GyN5JYkpAlu2B3WGV1yRFAltkTqqn0LScnaEMjxgZ21CTj2Tn+zRePSi
GMKnqJJ2weCnIpRhD9xJz58x/3jMbJqMSIVF6VBvkCHZIjn8VDU2HU32uvohSFD4
KOHXvXwZXmQ43LqDJDk+DzRaAkAX2qPVGHADzGUeKoLTNPgLJXPOe3peN+bVDUGk
7DVLGUTF+ejADUBjHrw3lbE+Ef0NHTVrRaf+Ti+cprAYrTZ/HgzJPPRBYWQimw68
CwOzevNyMOnfiF8W+99SipZGKlA238sx/lcxpzb3DiPuUzfy2HENG3r99NnyYXR9
X5ukOhisqdEu/K4Q0dmpZPVML3PXZAGCB5Zcq6LeSvGk52zZtWLyeM4vA3bBeTRM
UQ/b169aUawccVLan70A43Vx0LcBulaBrnwaSfiiwcKi7dOsqTvB+zxgGh8pp1Gq
4r1Pga9mli0m6hUkrQPTSpa3oldl+vAgGFNM7jxbIYh9Rvq/H1S3XeMx0/8VYHqn
2lwmXFHqmkwNQMKRbftfz/Wj/C420MpJKN2l9F5UitUE8Vej8DQpk2+3MZbCfztk
V17z+qp4cmF4506txCbETIB81ULs7Fi75yVHDX3wDISNhgyc7eM7Jp9BYsPxBBg0
zI/65JM7flxWdAL8NzJqz2C131L6w+Zg96MJUsAaq7rAwearMdB4+C7LXr87XDjl
4JlheSRJT5gDVO0AvWbojUfmHJLbC4ICk7XRS5eXWbNzZzADo+ZiYMpLcFb/P0Iq
DDttUT+zimaf+SpRAOaKP3Lgo1vLbj41Ihn/0y4BLslddtP+RA9xoW9fm1/6qK6C
jPmSBj9amtH7PbOaT52VVku7e7GWa6i01uyaTHt+7B/0EPJjwfPQ/jPlrGSDd0ua
G6i2Jp5naguelQGGaapQ8O77iocogd7hb/fTC4ZD4B5Qvw5g3YnSGsJv9rx0Ycnn
IErnnsBYn0sFBNFmH6s+98qtJSXTe25bKIztxHewwiQqUw6J3DE9B73CgxDX85PT
f+0JlD6HLTRP7Hm1F0JJ57xenYgov3xKrXdNLtv7xOLZ8s5IYAOpL94E6cmiMLDp
wbkHh4Rmd1oeS2q7Ln0iyW9h/20FLBVjZTBvOxX0bGZs2ceyyj+NOMnGLXNkASHD
qGeJqKUP+XESTmBuIHUGCa+f8durL9iE5nUc4hrJ9D9b4OeMwQjrxx0hst7man0C
oBkhtfB8VO3wjk3Ep4i5k7wqoqeAeWQuPu2Ym/re2omqPxwv5IyMv8gOjCRa2eGQ
S7Ev8yJwWFNVHuSRpnUoGbGln1zpZxSscbUl/OM/qH6j5b704WZg+/ibPU4rvoVo
Bunvhzq5kPufD+mhxXjpkl5yW7Jg1JqEVwzY3mWLdj12usOCN5uzGJHbpudPx3Tw
UQokfYjFUm8pFd5y5XDcPRoJIjNIZ1b+zenz126j5jdhMu/vwfS7gH5tF5ucCF6S
SoXjvMPTcKmAy8mUOeWB/XomcNft2yWjT/fQyNK8/nSLS0LQdqkQdrumoilK4wYw
KYH9M/yF9PVShkLaySrCldqQGJvQUiioLnIcv9VavAAPi/JwOAnt3zeKhl0nlJo8
0AI1+QRDXhf0giQVFprktHkT2HMdQpG5XM+L2EYwsS68uqSY8jGzYmJ078mADXuP
UfAakuLM7D3gs3AQle+wW5ei+21HX6p+WZm0K4rIzADJ6TdCEVNeqRoBpDx5WK0V
IZy/xCbsJt3qL/rYFy6aaEfgBCjf6z/UrICX6zhGKC83S+G1Yy/t1JpGsYYm4lHl
pQRDggIxOrTL7ygtZAzIjktgIzSBUla/uxL6TQIOvMIOi2F1ZG87IFUKsiyypvwB
jkdCQpfukiSFqsT0KaxS2yrn/DaHwdgzdO5WcYz1Josy++SrbDP9ACuHQlFTjq3E
HNZEZCbHJCk6x9HDl8ue8M3PP7mQMPopZ2Jm2fps45d4zW4vHJ6NzHmLiZl4k9aL
S5GzO1yb898p2wMZ+MH80KbqgIukndjWJhafKOMofFV/9ch5Ix7tzkyE1m7X3eZJ
0S/sany+ivS4cELwg339cLrzJJRuJJPf0aoyM8h3AkFOAPB3pzSoegnIO0uzHTUy
LSBajcrIRRmaC6LY/OpOZeMu/BGdQ/RAAwPopEHK9Y5TMhyo12Sx/kh81JYjfejS
z34frLqZLKvrnKbl+ewRffKujrtpsQ/cGms2xoFEbr+/qwyI9tha9qr/ragT6LpW
Hn1eCrz5qBV2ZSzJMxsvBSVQzpNHrAt49uo0Cg+DUGSUTI4WqbODVmTmjeIr/HPb
mQHd9ncCT4LTruAolftjogqsjrwQDeN6RQ2z6Z4wWMJWh/xPw134ND13x4Wqm0fS
6JtXR3jGgmPc2idgEA43+YSOEHt1a7Qr6+vW7hEmtH2OjB/XzoHwgn4w6SOp8YjP
CY+1Z3ylDEIkh+h9GhrhOuQjwbe/Bu3uMyRA9LGyiujFc0BAhuWOmnO0Gt4si4XC
GuE3pPJrSbF7FmvY1WZCulgQg/m+1tBKDF1u6sj17hxjo7mioXzAl31PVzVDMfWn
RgL8tTtEslBzf4Ph4Cpv1zLW6My0sv6vILAwbH9iA9s1+PTPiDT3p8Tr8ksSbKpK
fylMH8AaKfJQScaA88cWw+/WDoW6FNphfYwUd8hYuDUX1KrLSNMrJ4ZmdGkSXpqU
1g1owYuLQrPGvL+ZUX04y1qozaNwpFua+AMoi0db15eYnhdEPLToMXQ+/7nuZWFg
/AWvzEqgAL+onVkhbkyPOW8pTdfvUviJtkOrdVFzB9otDwhZqhmPWxsohWb27uMP
kU1bKDZUucJjNoTngqRtw0H6wQx2ShNOCOahsxSXJ4lHD4SbslBL/hX2sLltsBBp
kRomgiALfrhRB7zGvSTEcTvMWsBwbuH2kJywt8LsGKIR9r6NeBwGUdpIvz8GJR45
koPeZZLwCaWEUWl9WVTebzlLn5dGPveIQjIrxbgegA4kPrdR6Rd9HuLisizdwzRp
ipmFFWaPNPwG0xngHEPjwWWgOhV9kr1glYra/I+t/eRrCYrmthPul3zYbDKAsLOY
RMUksxzxKq1uDnI/tFaJSCz+W3iT3SAlzdVp4+1ppCdorfa7ZRKIWMmk653RUkPM
z8xAghpcZQhEd+MxTei//ctBwbTg8ywzrjCs8RQKloUjuVwynC7/h5ssf/xBv4AF
XRy8O9fn71SiEnrpud32IWcomXYlqh3wZSeV1mn5IpOau+xe8vylNXiDm3316OxE
js5uEjRLThoJMyvEPQWkU/eNctEAuQmOYf6/GaQ3JGuV00+ZD6xzRl8pdu33YU7q
lRM3wvTQeOXSVFHgtih7mj7zhi+m/jFPDtQSqnUx34+jcvkyfEX7hzrBYBWKJBIC
dyfd7LqPtvKHe2upxX+AylhYkgdwZIJn0qw7Ct5f80nFjhVdhTtxc7s1Xkyz3Bo1
Najs5msUAImNIegPGiK45C4ldoteMO6bDTeI5pMUyE0q4PfRWUzqkgU03vHf+hKc
syEs4IQ9X5dguQFh6rqkpeg00S/urir5Ddz/+vrurpHzFi81/ASabun2iid1swAp
TDjNGJ03ayEzCZ4BqXtlc2iIui2H0oJr2gC6cVwQ3WE0BzqIul8aXr+phvgK01LO
8SoYiRvP7EkNltDOCm2MK9bgg2PucFbD+iL+5lfnfFExAxdFepHXWBBD61YIztnb
eGO2guYASlFJ8pUk/JpPGy7Bg6YpYhtF4nOfZbFwjofqdxAEok2QhL1eEQNCg42s
M77z5j/JMxZJQ+2Tglv05trdTw2v5vsIVFRKmT3LrsVx/Ima894b2h/4pVTNzajZ
dHNcv2mus2MLVeuZ8VoRTdiBgzchy5WXGKLkcNSz91Gk2zsaGiBWpsXxdBVgvKbH
o7AsR8wIO2+Ovfo/bFVZz75mlvIcgX2IF7zLDw4UqZ2L1h3Syu+VLLjb3sPag84N
QKJuXVW0idxwfpzs9dOaN8Hi2D7MXD46i2HQQ5SGS1p2WinUBfbdniPxD3weFibp
wULgFiagHx/aZNDOafUrm37juWILdBc/UbmkidtIV9zn5bpj4GpJXUlRNAHL4/7q
5R42Tuz8lQJ81ylFT+PT8upIHlOd+peFUeFVwLOVLGzjazZ523M/x7NF9END9ghe
OPRRw7wRSHv675yyUdlV+44sBT7DPlbK3RxNz6l0mHBl9Mw4dFr5B5d72Iy8h+qQ
hmpe0knMWS3HueRFI316qoRJc2XJ7bW6H8rtG4KSp1JTN0QZXGA5Y71mQGbylcJb
9M4oOgZ5Fg7LcHSAqyYyv3xGPyd8o11645pjkbGv5d/N4Kj6iajdMX0K0SjmWbTp
zMAEAIdSse5eSlraTPLH0uaUYqx8+11Wtrj8fstpqYfTau6/l2z+PIJnfsD6s5oA
wjAPprqhcfGt8OJAje+jge2XYaYy9iaP2oEf8bPGvheIgWkCd1vTsZvpO7JwLrHA
mI0AvS407lQyrtTzhUXaagZSFatHsvoSL9iZgPgAbcVDuoMHLhXBSXPqYv6Wus3B
xRSLRT3biVHj1udQ44PwGjIaQ5t2nJyaYEJAfnZcI+7s6jP/lWU91JzUQVsv9q9C
+YHeF44jpNoAUlE+um3+6zou8tFmektwptYNvaMOdEuKByRgRFMc0JcJXmtIGFBr
NdC3xXRxpn64DTxdFQS+mJg5xv7z1tCWtYeCQa8tv+3KhxByHL5RsL08Y/W+kT5m
0GIXJCwvZd2ocVm8lrwsCLIi501qpUWUGNaI/XXymX2PkRZsgDlF1ydMUFwRRdll
Ec9GZPZWJxSrFcgsffyvyeOqyC40agryndJmdhv8BuKJF4aSpFuq7RyEEXgjCPIJ
mfu5lS9lSN/RMv1e8bAeF146Y7wHIiuY0Hi1ISCkFD/aD9CmXIkIjjKfmvyh9VNa
RldYrH5D5vY7fDr8j28irBNM4nO0/MCs2z8x4bIq9trw87eekPBtMA60S495RXfj
pxiPDXUgkoI6ZPldhSg4xahkYzPErvvzcOqIrUqsKFFEK5prAbwOvgi13SMryscF
Ke0LyK//guGM1MrVA/EWD1xBR9+Hg8j3o0H1Hcb1jsbl3bJ8qisjEt8eyxkBC5lx
8YF7T4Q6/FHofd1dKRBcN/jY1qUVA/aU04+F7fodscF8EOsK1SkrolnBFxQ0VKAJ
7R1W9MvokoS7O1rjCloOXbkd6kay3GPlBh0rNzE1GLw7esxjKDmPwVKeyh3uqdmE
+6ATxNGyq/GM1NA0Hysqohaa8ONzTyyyohp2F4hD08OdzTE7xNdlMAt8twEQr54r
iwVVNMJSQ6PsRVDHo3r9pAknQFdHcA+2j43lRU1dtsMO1ZPmQj1vs+ngSTtxLQFr
8wXdZu+XPm1OEbDHT1M8hFblISB2++75U6V7wGmDj2xnZ4ztXNbUXjz3Hzz1iWQe
Cu2JBwppvZ5Ia2d5WUTY7hbTLpeOyvvbNNIlfiU5hi//GYNCe3tESJq0m5VDifrE
zX4hUNF39r3EHJ8nL//C7Iew4SO8IOhWmFUAZnA5HaKK/z9tFFkTDva8Q1rJu3/T
0W9Qk5PkGL/Wd9lVf3Cjp9hbTXQKue/AwinJCkPwfStdhS/ClpDLcV+aRLrPIpWk
E0iFSUaq6/cLw0gGEzIwT9+F5IFcMutUV9TLc5D7zLmiYq+5X+DMCpS4G32RTMTj
U/nRzQTZf9vImj1moFC1oI2ivvC0rl+85vX2RzWu1qbfwJCGyXB/FJ3exJ2Oshj7
re30nPvb/bIqUXPVTvUxFW4RxhFIVVkibQi5Ks17hBX++uzW5gPLoYZZhfjmEA9L
5f5Le4zn0JUevw+SxEm/Tb0n6lecji5+WTWZXUfveQ0Ai5jSaEjvnYMPIx6JntuH
/M4d4ZP7l3/hFn8I+kjcRAlHz7yi9VBtQWuA5fUz3F1z/3OrQLHzzBsUgiTZzEnY
iSyscz7isIjDquMo6SLFebXL973h3a0wTbikTBwUtotbxEM6br/+Xp+0TKQlVAjP
s5IfOBmXnMEwevVnrWbIOJHMq/pSFH+DwjVHDCwaFF4TS1y8etoPi3bovMAOngbp
akqHsNmG4dlcfH8m4ve0RM4zl7JUsgAgBUmELR3zTFuiKkyPex1q5i7A5h5yhihK
smoZ6c7HSMnBNUbCLGKbh8YqrvTUvpaVM8fRsx+jOMVgIAcfA7HtmkfxC1pn8vuV
BtP/swvrHfzmNtBdV/ztyEMvBRne9OIoPCzAqPJqXtT3fhOEFquh3/FWKnujIdFK
c5XXBgYNmTMGqSCORaguNCEuVWKNVff64OMwbVNiS0YDHa9nuzPjDTVn1NQ0i6Fd
eyB1Pos6hx/imV5O5tpG+4xJwgSQveP8lpZPgI2hTrB/aWuxQ3ifERRUs96zQEWP
S+WQ/PMBKtp8deTgwJQzxz8wgyb0Iiw8E4KzdFIg+Dd+V/9iS6EUh04TlMYP333E
TcCnCZDGlTu5Bqw4EF/P2uvp4uE+dX/FcHaOLF5JHLiEHe9yOgz+PCt6I3CAr2HC
0QIvmgtAxoI7bLFh7Xap6a7dqK1wIGm8Cva3VYZbKL3XYYzhHb1lqGIiuBPBuRzX
Y0btui/PZdaUJygO/Sz3uQ+BRsIDBLiZVUvdAhVgJYphfvMjorni/nOQs6i9n7pD
M/T6yDWwA/pPcusSPBf/3afkVa9zDgVGuPH/y7Unq5sW8+aokUaxSBJXSqJLgNMR
0GOlObHmGcGyUPncJg5/e6z0FHkcxqXxB5i4/ArgW94p2ijGusgZzSbEnnPFXDcG
i4Ie4iaOMjLVjh0yhNHJuvS3MPxVZm4HEtYj5qvlXcv4FgyAXkJ+96DjObUjFbHn
9bXpU/tBlNxkCXyJA9FaFa+51M0N7xpQJGQGZZTtdxxZY0ZZx+zxSwOrc6YGsoyl
EvwNQMviUyyJdhyQsjhcsEEotFMxQFnh2l0lkHoy4U9Uf1BUYaUuNeFGe8mDWKAH
ImhmwwJW34Om3WuWMYQYCnw6ESdTqyihqdf/3wUV6311nJz8CvWsNR0fNefy1CDW
i9GaRbyUEltfO+fKk3fFmTH+wW5u6raKgVFyFJwbyUOY3vktckGB5ii4U1nqH5Ny
WGy7Y5K0oT2xQfzyxswZv8k3+f7Vho4r82zlFrYkwY9kkmnkLaUdMjevAufmt0v9
XnDOJB/qK+yHZH8XivwEiZefzNVNiCFprtJjMv6MFzJDuLN4Zn6TRZNcz5sMiZhT
QvReDUf5gJvy0OnLCOhso8ADf5geWD/z5dlusjSddEKr/JHP0j9xti+WDViMJYiJ
4k7tjCB8+HmlK6fPRY08sxSQPqtcKQnHDoyCg/PjBdtNWRIwZSrylHxsVoAkJo0C
pA/+2FBzpE//XUYcAJHYs9d+ISBkjZeNpxoHsejPDZaoCcfQFAbBPvQkEKWh3E6E
knEbBUAdpCo35PuHi72JXaZGrN0nb/wAa/cgxhpvFTNZXoUd5DC3qfu9WITeF1gB
SLUbJap8yl5AFC+ryXtOJKrZXsHNys2qAQCdE2P4nBN/q/ltm8jfhyD9S2V4S1su
OZROEzk+ROe88uVuyWmE5v9+uEksYsv0uMmvquQ920dAsoOZKCNTqyVQF0dqwQHy
s9FmZp/qYVcz2urqcN+7g/tHOI2eieQS6c2Dv1AGwbVI2Rd784heiySllPFivYjA
EIhRlj/qKtez4j027k+6i9k9I7PoWUEUjCxcMI0eHv4IH3Nj/zEOBylSy7P+3OcP
vZ7AwNcBErXV2DcHSluWgLxCuCfe6ZQksPfjiqHuui8Y/6EEbNS0IQedU/663mNI
Ap/qSPWZWdR4zs09gsZVGDPUfG/zY+OPjHgE9l+vo45b72W1iw11MxhXkmtiClCq
UFia9ncY4dWGs9rbgaK3gBrIjb7Wq2qg+jg82IyUm5iviTOC27yE8CuLk3Tc+z0q
7N3k+yNOyQ3KpaMAWnL0GsAkX4VvktPm6Stenh35VLYvlByHfTpOtTo2X8rEwzJg
Rvhm91TS1Cv22yfDeestnIDJNOgy8wYCRbmf7Gus0Up+fKzaafPYMcQGUrAxMLVp
kL0VuQWIdGcynYyO+rISSdqKPpxUcy9vuTLQfSvlu2HdyNODSfs77zPvFgHs8ANK
MAjaeAl/zaOidZ0QKq1f9y6P4yus0Q2h5UPdk7kJZdMLdVPYdVhGQtk3aVmUM3Wo
5xs5HBWPDSJKvUcrTUZA6diQC+rI9vQF04DSWehYSGq+sx+xCRCk13r19deI//Ag
9Hv2aI7NUQhoNAXnIp86Chp73AG5LKI3Z923t2jOvwrU3HMIOXtPc2VBKUWrs276
7fWbhIDLxPy/FPLa16xe5cLAuETiKR+xwWAZIFSorJQ+vSwUDZeooNW0Oe7Fv5Wm
0yY7BiYypV0EBzzG9UJtPzbrxMRF4qMGK7RDT0Vcyodstow4Qkzv3bmEq5oGQhm7
20aioxgyyZCdiTkP+mTiLPNBlJfnHfUmwrWY8/2cCUCGYGVs8wjHxapOq7w8aNwp
wi6MgAqBkYM7M0PStF8lre4odRglWce6+y5ZGHB0AJZbHnEGUYjCuZ+hcOvipvT7
Jn/dBR/OSKrFG4BMK2vE+bWrPZBFBE2UWtjbFROeOq8xyV+kTgpKeJ4uYFwxpzkT
VMLUWMPP0u19jFP7xtULSYhXGSDWLNnnnaEu1QX0S9fWHOIjRrBkjrngHDDTP3tD
EO7J7GLoCBTQPZTzyPqX8/E8j2qChnVvG9N1MvpdmjfgdmlIEJcvnT0ih3LN1nLr
E/8JJddSxBPNgCCNJJ5L1RpD+LNtTp69G95PN1a2DiJ/G/3y5k1x1geTLAvBav6j
tLfY9RtrEcTgbpPRq/y+ZWRCggMnb+La7YI3olrbAGJMTGXh3omGYQRRWP9gS6Xj
OGyycReIq1KefP39gRQLL9ZihZOhu5EULSXZXmVEO0OOI7fC9G8Va+KAPrsGkUjJ
QiNOXDk7PO9KaG5eQ3AOMN4q+++Ej2TMFAMGHZSnsPf1xqdCOFoHvAYWMzes852S
Hcs/xcOtQSc5K3mQRufgnvRNftVDMCS2kGYL6r4EIuLcNMhGOLKPa8rwyE24cioP
76A2YkNf4sm+mbRL37FImAMyr0+gKc5MyWmX2N5A+AsLFR3ptRuB/KkOncCWVkFV
kbQ5vB+6LIswK2isNidtjkslCmYw5bL6YS5nY8Mw7h09HbAKSMWJglunnlZaqPsh
PApl0pCwsDfrroINCaDI/igsUiDNo2Qkaf7INbY9l02khWarHV9CqE9eRyRh4q7G
3eQYUDC7a9vlsIwySDIoQ4ccLxmtS0UJ8xrjiLHcEEZroGFg9jNl/Fdjc4jlt8cB
RYvt+wRO83YDLc+zBdiFvKucCrYcCl0/T6JGLlEVnbvHkgqp1xpurtkh94p1k2Lq
sBlFLq7hy3M7u/qCeRdmhKnlqcvqFQFEWMLE6+GuC9ZJIDl8ehWRoiK+hNa22nKa
bCqX/hN0e6+W78rxSbF6C2aeNWsBAmA79nFdG6RIbYHLs0cHxXsGr1ysNJ2XLU3m
BIvhaJ6fb0zcbd+Ac9Ilh1AlxWz1ahajrvqXaf+hayL1u9s+MvrX53sU/ctV3zPu
FZaf28t6bUuH2o11fp1/2GlC+1hwHpk5u4lQHAussDJaPnIsz8XWNHHfuriXCl54
ZWv+evB2nr68PbBGApQ+ZHnIESIga2YfRbcTqxkpxzP6SUXm/MiLxuybsJkA1EPn
uP6rnNSEZUXa4xvTXIAf3VLAuAHjBeRgVHSKoCh8Xz5/WuO4vb/r1WiAdtXHJKNx
2FN+oZZl8xBnUGD447PXKjK9ZLzSNCEyW3iUFQJEnFpz9wssKW4bCjm3dHv4onii
NqLiA9yysYTKPnF7xjVU8paAjfICgkUAY0rjPDVTM02SZIvVNZEZMPKmPL6kSGYx
hfc2rbpOYc32mYjgMZERY0BgICuVKomcPB2dDSaN6pMvvO0LrsR/LC4F7GBdiwSt
qiCZp08BsLPFm9JSZezuhgoBXk9DqCIZSGSGSBOiTQhiZ7mfmTK6CRq1bVTM8A/D
7m+1jUD3HOlAtU5ES5tVk08iOWUrDnavYjFi3g1YRMCvIX00rqllctBToUoMC/wd
HS/FGUnkYj9EcXzFwOrBk46bNlmFHxOiKF9zdPNfTPU6KT843znqE7AuA0tSdCPw
J15thW3YzLJZyUTURbRmRhRcdtc0pCuITS7UOEN3bkIscgLcBWpRubL4PLpoKPWX
7RSg7Ru/Ch82G9GKvqNIakInxEIJs11sTxjpRHgMlzu3T/XpTEYY6AvWjoLDw2Gp
QUVpMrU4KV2OWMmMivzn6R4ZayhBdADGVR5SqeXIQc+AVzJf8GHkKo7JGZXiVtBD
uamo4v0EB4ru+IvJxQj+GyNefxGiBiAAFxs3/f6iVmQ4uvt/yivyryng2MX6fcXH
jBXJ+EZL6AUEdp5o0dzqpt2c5dSwc1JVxRhvVywf6fmsJkV6gRLSv7L8jV3Q0cLZ
fxGhaV2mUmEmrUREp2CBmovBkXtQl0YyFprHtRy5+H+AdZK+cvBXF79SIBS7KEtt
6VcvXiO+D5tAm/JARqP3U6Gq1PKm6EdHj5OLuu9WhvJLEZ0kXy38jr/DUGxDb6C3
6TFi9X1SAvBO5fgRQUDchPv9p7x/MNpnFKQpDEW6acQdVT3KKGp/aHiJ7a61q0sK
IAaktAVbMf2fA01ZmwoK4OP55JJCl+EPELK7QMfvmRI3eevQLFMwaD590Cn8WJo4
5e7FpiEFFCA3dTzL9e0HChCupvSH91NLMW+e8nuTvB/ASuXI9EaFOsTejwHGWKRQ
+WHEGrjIqoPXEf1UrCu85VrsG8yaySBjt+PuVmRhBCivpOgtNmbIPQXYTYVppOfO
26jXZs46vmiJxXHnDJyj/GNv0TDi2Qqeez5S1D26JDiyPeVCX0F8icxN7lfJdotp
9P/1NpmkR3nIxOMS79dJUXBiTTKoTJrkf4Z7gO49+0Khaq0J7MsL6r04fV/TiRwP
o7H0gzvMR58uzRKAVU3i51QS6nd9DzZWG7h66mHZ//B++wvVysQPJqnPs6lM1mGF
EPaOB5oO5/xIrnyZnnW2XqjTs7zObLwdPLi44C/3SYkehT4DZan34DsGmVPxHB3C
9kMGVmp1ge8VLV3Jasbl5cl+7KDePLll3cUEef5fEkwilNY8jogInLuRGzSbvm2Y
bh59WN18ieOwb1WocH/f2jB/7nHohEzgUrIcyPRlflU=
--pragma protect end_data_block
--pragma protect digest_block
ucfcOsVDFejN1tfpwwI+St3hPe4=
--pragma protect end_digest_block
--pragma protect end_protected
