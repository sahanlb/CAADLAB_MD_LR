-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
eA0Q3lYwOs6gh1Y4w+NiAUe5v1Sxrb3cDNZf6hLhzYcUPdjkjfJjlZzBpkTf4tdn
rnhypt0sa0uDd53s/Aj1mpSodlzNOflJahUFjG5wIGK2MmP2/EmgzEK7zxSkGWmM
wpU7O633w94vzL1Oiis/tYV2BHQojW6vs0TCYy9zyQM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7600)
`protect data_block
kakXw+pk1wEzlwEhFCI9RtGpJfgu+TaJ2DtVC9vImDCPg6wzGmkGa2mZvhumrxR6
3j1VNJUDpc+vl9TNH1oeimyr7XnJSNm2XrjMIXBC4hY08yq6duFiANocIWD8J+le
cOzLFtCL/obGEBqhT5/pt8RVGr3VFjT2845olcO9q3Xm+IjcA9CGcKqlbLaiPVh3
KpLH+Mmz5dh+6hN90AqOexN91j/vO880RhWSEZyYwshvwdlfSjDCKRkRCwg7rL99
lB3pxAOv0pmy1awXcjatLlTHQ3MURExr+3jYnG+uf9RqQHhU/9i4vrcUdamzV6dM
Y/moNQ1VMvrMBn3Al5WXQRFiqMxVezqKuQLOUV6tlWeToeDVjCxtzgnzv1zI/MCe
Jdi3zsc4+8tNImicbHhVJj5+UQIQoRdWqJn5d6sI+GPOtLHVQ83jyMAe6Q88+Yyg
KZxdX5rERL5b9yasevjLb3T38PU6Jo3Tk1mB7My+fulhAVYCqSQTuolmSHzlUqJ6
ElI7wdFrFvrpUxqZigVPA9LurJcIZqnFLWcJD0sCT1kycPX7BMjBdccRt9FyFrjF
rqNfTW+/E3stPaxzX53wxA/vYKMzTisD9NeOaSFJ3v4l/sD+JPwIoanMY94K1vYo
/huXxoUQosCklOqapzoAfXlJl04GA5j1zwXf+l98jnFwr2RggklPbKyGbxoeVchG
MYMwDfze9S4lqQs3xBLrUmEK2h6IkyhKPmO+WUCqI751qulTcsmlQB3Vv2Z9Ql8o
nizvFByJx/tYMtBbBDh/nKrGQxhsN4HYznfVZNCZYfZX4v88EvzN/N7b/QIk1APz
0Yk46he7lbqmOQJaGWdncNDktyT9/tjVs7AhE02ejYSAMuW4jqdcgsJ+j+DFwDIO
e//x+YGA7xVCjtmlySzydltQCKrb5vt3vXPp+u+lGMy+8HvKuS4eazkH+h8XuMcv
tb99HI7TFApMpz3eZEZb1cl5H6Mk8UyDCzHOGNEIqxKRCPr6plKRPSywMwsSb+Eq
R+DviC07kUa6zL1u+CmE8pGBk32zgs+CxNswuhkZuHn/L7Y82Uf8gBcpUXOV+d0J
E2sDgCTzuO4mRxSy3iepo0MDZCBPg2/2o3LN/MTlosnSqY89jhjiGdVcHnxmBsJK
1F1fNcTuJoBhBZcDwG74MuXVE9yp/tM0H4lT44XXwWB97WZa6RdJzrxrTr9mA8qn
f41KGd8KXhpY35nF9Q9wAc/8WseUMrAaV+eCFC08SyqtxG80DPQFytywagS1Gq7R
EomwAwT6UFOaW1B6ogKqWiO1yigxws+RV8jMHyQJVHk94BoACP0QgQd9EsCFwKpi
1CuWMSBytBPOggKnoVdrhzrp0sRVdc+olpk8KzwmrNyU1CkmuzaGOJ9nI4+g8CO2
dFRzkb76vVVNviEIpRG7DHyvwHhQ+F8zCtzVtzF57XRyWbVrGVrrIH+/5BNkzyUF
eY5vLLqq4/DdVHSM5PD2gl5FNIS/D+rAUhNuDZc5Hwjn04lfNOwCjZ2Q3WK/JXX1
YsVrAFUXRpb7YN6o1hwRz0hj8OlWKcznbuLxcNzEgmwppyCHgR9jnRk3QriQEjGU
1j6H6hsf8t/gERNIe/0bu8MgYg/HK6/accfxIzUp5cmDy+F9KRaW3ycKEi1Cbbdv
2sI259WotExi4vI/uyg0xCk/pQKYh10KBo0JXqq3v0mTER11lfr6o3/zGv3M8hiL
zv03fpsDHX1hkSglv8w5PciRkRSoZ6hJy2SrzWYTnqx9SSbVyx8o48jJSVPrOWJS
QRKo3I9/FnCCiS20CtCN2d/nGyet6Gv/RxIPEWgWSGPsz/S2T8QzctF4NSFaw4ih
TE+IadPdtZo/YQT/R+fdIX5beCkYowas/TMm83zPZBg8lhKTrBkLJPyPsKQEEjOO
4r55ARcJAVBwN3nCYkC/GzVljbRd8Jsrjcscq4n7tdeeMPIO8OIIhLeRM0o0XH5k
191ylGqBrB32G1DjF9pYikUKDwxBI6oSWzldfZxvWL+532DLhaPvznA1e2pwVDF7
V5jS+kIDgeB0SS26cawZovH3VdgJwxEXXzXACok880IVIhunoRYKvfyrTXUObM7i
Xs5ow4E7Vtdf5QEuemDQ+MuCvq7U/sG/b2SVv9gWCFJy418u+cM45B772HEde7WG
fBhBwKSvDKghwUcZKSdyJRH8oP4p4RpI5hhYj6S23W6fHzmZHpW88lyDyCXUqy9W
FsfoXtTk2GdMWLlLKdwEtEs9+eufeQL7H0isHtNmFNVgA+ofSwWMiF5+ncz8Wbbo
h65VlcJ8TVr92fsvcoGJqL9MOBxuTpAu3dklqSdN2gNjuYLyyE1qIePr4hBAahRe
BHCXMWLmS6AWNj6CWYfJgagCiEtEFYR9VRPOwBrM3JK7irmlSz4ql41i5NaBaCg1
rz6289wQHHfxuhNPddO/ge7JdiHdgs0MHtn9WYkspEnm6kJ/RJaHR0rFy7wJFwJ+
h5MvpmANL+yV2ot8A45V1Zhcq0XcDGZj+Nfxym9I6t6sHu4rByhDin9yJ9Cb5IdH
43eLF5Nbj9uPX+YCPh5Al0ttQgIG2LUb20a/IGFPnViv9b87QRfzw5mkn7AMg6Hy
/XD7JYM77Y6zzcnTb9DKKkc50xdQXsdGHHxIXk9fcn0c8Oq8OhKX2prszk1LNiuO
9Uxz6L5OiSB2rNvQB7dJSkvxCd9YESBeAu4AkVk3P6DOaa6Lsp744J/zy+k1C61D
mGWcW/xu3YUj072g167RR425a3dRVdOYD0dqTdJ76MsT5MY45anL5a3CRYOL7/Bs
hIYXg8iM8Ws/f470qbAsjbRh9JNKho5a565dWctsAgcjxTHqRNW6HrxzPqPb7vJ4
3/Vtga5C5MpQ3uE58xNirlNfDcGyB+nWsUwt2ryDNAc8Q4/I1DPdcY6yU65Bi51Q
gZnCcTYvHz+mzjKQDK0z5DGe82lizIxNIYyI65gzkU+m8pukA6zgfn5fcHTQclkl
84PKuWzgrPOaV9QexC+XP7LZpBQUEsiVtydzRB87M9tZjLQNRl0xsQAyM0akNKTG
akXUu7Mz0QkNbBaeUcDthHmI7CPH7Yiq/0lP9pjbcdqBcOF7AGLSPfWm8q2OA74o
TRObdOPrtS0GzFtzN7iIzfWp5v/hBUzKLu+TzEFCcWq+TsPLPS/cNM3ynptIftc5
XfNBX189G37dt9h5NJiZ/ky2/eAuDEa8a7dkMc20ijzZffZz+1wSTXu7Vg5lmppr
hNUbjUwhqd4rAzp606xUhy2RD5CdtzY+7ARxYSwWw2dLqxDDFrkc+N58OhxN97Iv
8TRRkpyagRBTy/LvdawfZ1sAMVeBLOgWWaHJJvvF8Gw8ZNURR+n7X71L7T/zAdTJ
or4FrUoK/1a0l5jfeejLPe+xZ4SOGtQwk/lUtVYzMSJR6Q7uGbTEQyHzFcqWkiW2
sZyEpiliXm0s/C77dsbIIO6P6dil+dbREx+mQem83pFmP3Opfh7OvIO68EdEPlHu
dB2PYG+XRXnwI/l0amiKZWaZfXcqnsPRoPNuOkOyRfP7ymMcMzj5TiK+I5C4E6op
IX3EVaHAg8a5hYunsqcchERqaLc9MbsbV2RQDRmlQHTijpKdpRaHgzd5WQqFz2tG
24nzminjG9TkdMxiIKTyzP1pOXzTCF75XEM+Gg31bbAskMb2cEt2/yWd4aMCPgMo
Sw8nYNjoZ46AuFoga5g50Satbdw+VCi7pp4f/hDhUSS7mbDBKOxoIUxFdhXWcLcA
FK/nzBNptoUIxMGJAsQlaErhm30NKIZbnOvjEzHDgkeY0y/++sI6Vfot4NpO+V4w
+Hq5atf1Anvs632nLahCrBS8kxU0TOykzhVButmIUAyDfYVAwWS3VgvsPFtjE93L
InmuJgrW0xVObk+WfoBKKmjQZ7PIeEEXPMmUqdqcXylp2pJG+t+TwmZ4OsrK+Tbg
rXjlldyonZ0+LHqlSbHx3zf/XIJsg8xv3ztXfJDOq/Zvnhiui53W3dHrXNi96Dcs
MBwlHdtEU9A9GPntoatEcvcSdu+nmY82BuKQ0oNktuJA2uYWLlEksxPIXVIUeMZf
uZ9mm3la9ZGshr2lnw1q02XU8pXJi5OlTuzPLMd7a1fNH0ZqbsWCl+NyFOEYpWrW
pyYSJgSs2R/cwtW4vGKT/7a33ftgsCWFJR7ma9qLKdiBkUeeqENzWAZwuuc5GkQA
TWMfnOeAprT3lhaD+o6ukO6uv1abhCjYfWWH9YWuFALI6f4V/E5mvcX+4JUwLmym
0dG1fBeDHFRB1YFxlndk8lXGA/Jn7bXZdQEC1RpTP6UNL3xVXmCsn/UuAZGzBFVv
JsDznopdd1isLfuOQpt5HOETYEBhLlAMdwvcUgeQmEHvGvyQ+oHs2zZB4C/+rD+4
b2xWXVPdXjIP8QUQZhsNLiSd/WlTOL47C3Kc4Ba3z+lTdSfOxKAfm8JYur3TUQcn
sGjlynyDaJrCVTGo+aSRqWCLXtQSO/d/wC3MZtgo1YjMxSUsxeK1vF00Pp4ca1qR
731+0Wz9MwR6X10dGOMnsijSi+pquYBneXI3W+IkpXyJAPQETfRZvjM/r67fRme7
GUh83Gkbp7EHohRoNc0tKfbNqgQrp3YCrLlqswys24upMDhJLyoArdYn0n+acHrH
vGLZ4g9d2WFmDXICwhEI38nvZNaPf0Fv7kj1aJcbNfXOgCQY1hlIRQL/cVrM/q5M
pxoL4RVoVLBnakYtOy/B8eVOAZJTE5rAQihwV+zc4fP7/VltbSicpPskdR9KMSGp
waG4tWx27I5cxR0c2+h8cfDADJXuWScQglg6DlJrRlIkgy/Oc0gXFFS1bQRViH4/
EqykkozQQ1cqvUtSfkUOS7Q84C1MpxmM1wRr3cGBrdHQRrgemqCYiLirLj/jSyx/
FNKLuGqmnwtROk+SGwKc+bEe+/t70wqm1VX49t5nQ4iSYLxtR5o5OVQRwYwUJS5z
xsymEBTytV1teqokF2d0bHjZePLvjVmJOaSQydx8Qb0gNxYdvcq/22MkesRqdLRy
zZ6GnB+6K5yYTF0qUt66U1ZhinUTAOjg7rpsPI658V/uDoMaqVQQTRMd8hhOZfrD
Gcc8LR3u9y40HnjFgjK70y/dThcujehCVl21VBerVWuoTppLREqYHfUf1ORsmzw1
36sUT6/iGYy1/QG0uhSMAlso+SFR2U5eDI5HzYnBnpP6FYzbDZYYreFhzd1G8wgJ
Ij2SJaeOkEh0bylGwVKi9Vm7MnBlD5UEFyr9NVC3D7gT3ge6c31KJtrYE7DVxzHz
T4S/SDIxHsmT/8fKjF+YOEG/hwKqzuD4OXVKrDLlQk2N1clV9vzymONXK6WCqKfE
ob6ssegq65rzEmzGXFz7xzhALzNGnNFxa3IrjpQ1F65dZsAH+UJ97a7qdWRQ5HVh
gVJjhJr3jQQOdUVfo4zN8l9QFKpv3ZR/EsuVzFzrKBRjCtLwY5j83Rpx4TuwbOek
NW1wWWyEKyIshaQzPA/PopZrN+ZFgxt8amx5P7k3Ko2KajeQGosr96TvOzR/upX6
AAVt1OJt3+9mIYeEPlwEjwOk609E1uvl+l/+d/u14c5T5g4oaX1ip0+W7IPM2DrV
r4kRG7beNbAudGysvis/aBXANrberidqQnuFesjWpPFdWt8lj8HJ0279a9OSFIXE
u+UT+/hGVpWauvwTbGyMrABPUYnhvvX/y4qCBFXVd3WSJXoygBmuVImdg5KOP2j3
LtJAjHrb4I5Sa6rVEmOkWjKOPBEPjFmIRSDQ72oE6u963Ddtzl542GwYI0rqgj2w
uDQOtp9Z3B+yiIk44wRJtVc+vuFtTKk713f5BNtk2zGs7J3pLwjx2RuHJb2e7/vZ
LSjfgODQzbXlsbJdPzjsvDk194rQp+NW9RsivRpZ7+wtpyGHgMc6U9CKto7p37f1
bjY4jImX8S9auuCPXoRSDu1LyQEYQl8WDqPbG7s6/vVFR7SsUfMmyUZhV0U7DGgC
OMGlnYiruqTnP99rdsMwK4iYAVAjysE0MxlWTnswzxTY4IcB2LTXl10JvjykCMNQ
bo3B5P1eLSzQdRbOWqZfFcFXcxrJlVTg3ulF5YHNPBOP3NiTMQQPkPDbUXdEbNGy
o3HfssChfVkMCLjgBiuU0BaTwbzGuY+DKGG0slILtJzePkluVGWkY1sa+oGBfKdW
QpQmz0NMx6rH5IJN4RYoo+YtBqryX/BTmv9yCRwgiFSIQwp3Z8DiMFzJyL0AaeOO
JYep8ApXupynPcYPtHYUvQtbu7DAw3I95/CatmzfWu1NAuzCkvsbrFck+ij6wHPz
ygYOzOALuLM0hIQ4AvKd6bM8PMILCuB+cturA1NX3smyWHnjZyAz4BSVqdYStKTx
g/3xuyEpH3+G1MV7S3s7PepmqGzFiE2Mji7hjX3PpoAYJXypM8ulZkWB66fxKXJT
oeU1slnmN7EA6frgBszC+6tXdbLL5Z0uKCYcCgo/JKpdZZdyNsPvBGHOyKspCqHL
QKmkTSYlnyMYxb3bdCgKvjVK7IywAnbDG0sdaRplNa6y+0pfB/ZrSHcez3SdbHf/
m2/aWINuL4+rr/hPKdwf6VRyCpbTcIbxUWiL8Jpemj/nAplMpCPSlmc3uTviw3pz
T4gW+mnM1U7vjMCipkqVLky0mi6vWuYZL7etbqLK0i7kCL/PkTeHUFKutM1gSCrj
XqHsK0X03Dv0vYlwkHG4zSNb5pULE6iO3pC2dA7ZAz8WsgunTroRpRx0fCEg2FVV
gSrJQfjghGnZmNCcgsJMGtqkRRG0xJQjaLD1HoEEjDKYeW46w/oB5Wfr8vTaw5XA
T9GoZIoFAyFUmwHpMV14rHDt1bFU7B9iEczNNqZ81IWzmikZqjUAloo1JzDATCJF
11WGgO0RUaa/6mqZ5qwMsT1PI8AF4oNt8s33BdVsCiQY03cme/DGNFbAwOd977e5
999vj/6LCbq+/K1wkf7aiS93dI5CDQ52WebyrCjRAhaEQd/Uqzxyq+Jr6nV8G7BA
Rwd6Rs6WOB0fFoHOnhDHWF8t0bsMTshlvKPjl5VxUtH+BdBz8Z12tMtykVILydD/
c/EtVEWaGYE72KuLbVZefPWYFv1j8NTFf7WBVZY8Ux3ooA+r4dIo8uwif4hFM2bP
awnAkG6jTrg+BQkYHrfTPcaHZlWvfJi6S/qlilPDvRHj79rJ6E0HF9d0NIDNXXe4
DVM3qkAqBGBJXjOpqOImKH6nWCNZ1lM5BhvEFjueWiVvGupIdZE9/Wp6YJgobXud
TNs5f/aF8jdYybFknMrjyccTbPRoMfcTTL08/mr7CrVShgRMzty/m3DnC5+gaK6J
nf/1Nz7IkrUsABAbqv4oKwdHWANhEulUeHBhSVtmSrhXwYXFM/3/Rvk/2NtOViVW
uQLBUEsk1SiwClz0yBaPcnjO6qBS1+I3FYwPxtKZhKt+8OexxBibiR3GYdGfpii6
zLrOCfJHlvx3won4Rcsn5GoDKHUhi8C6+BjoWK9Z5BaT7bRbWRs/9+86gj/8mswi
knaWAtZT2RdtDJz6TupizYDol3PT8BCGhL9xBtDWA/CPsPlNKvt0Ov/c0t6rhfql
ssOVQo5Uh56aikm1jJd/TKKr2tPArvEXQWfBuf4uOc0LV68AKUI4UpOAIk+JkR3Q
/lTjdJaCZztcUYQ5eRFQ6GqTxbtVUpTCd9bldw4MQTANcjA9vkF5H5KLkboBYrzx
HMnGcvyeuksiB2aVtu/HjeK7hxigfRm1FM1Bkvg2lLgkv4DemhrdpmdzBLkGY8kq
jlClrJrRPomYViWsOT60go5U1nlBYCl6HChCguNmmVNSXhkWWf9laqGkWNqiJi0m
61vU9JmUpjqVhdcdiwLtYJziLzvFJoKnqAmB5Xi/rnhvSmgE6cyOAuBkv7ViL5fD
HHNfNCE9rMJ0FHysAc4bGszQlxefs6yxFEzyD3O1ASd3ce0UZPVzZng9g9XGWOx7
34hwQq6Vp5J8vAgLODEHqiJc9jb4Qi/8ooEl/mhnSayJGkavegHBLQjFm3HbOmVT
WVEfO0EvdXNQ0ayrg+OaPcv/x3EHg4+5yM+A5Mi+Alpawe6icTN4YOfwKVx0mR9n
N2RwQK2m+bvzzBnJr5vIF/0RtIZIXZMMgvXQ5hGKjRhq3DfSKCWyIX0ZDwtxBFts
28ZUcIIIwVywkiMVC8iCv/j2bnKT5gY/1bQrXPSL0+dP4hpnUZew8/AaBRZqLOwn
Qczf3ahYT0+wUBrHFe43B4a0hSKWYZE1cfTZngjXuAhC7MbLnkD0JfnL1ZUqUK7h
He6PFzQ556ADwydPkdfu683lvW0gPXDRnnkfUdSrwmW11WWYdD5HO3aRIpNra0ln
7C/e2CNrTiARj4P7uwBYG5z+Gv6Qb5MkhEu7otFvPek3/m+XJSg+HfVEAxapmq4e
k6/86EIVRK8Ox6OQrGaI0fi9/9IM1BQZ/+ZHtQY/2DuxW3HGlzeJTigN9/oRkXmb
jyGdMB/ylhghYavVsEnFKggiv/pgi/c0FgkNAKxaupbPuOPhIfOYtRztcClin7py
k876rLUZM7lVZALOu8QO5MELrtgAAoFU9gp2nZ9JwcaHgqKYxecCoC0nepHujIQo
8QuRTfBmWnqeAeTbwJt8iTNMm4SMM+EW6Sy+RuOW6kvz6EgiAkzdaRUtdZm1dBzE
QMrOskY/1uv5AB8f8WodEnqrBOlaiP9vFv5v1i7oP19DmpQAlVarvHwKuR1E6RHD
DdCwe4vN5ifeXnU1tOie72TM2ciKghVWidd+88VZ3GWtvaicNE/U9HPEAVQGb8hd
ngNjjcpw3CgowDtRrQvBJ8W+dbXbrCyV3/J6Z5TwvupW3p6GivZ9mIx3dnGmHKWo
RQp/Y7Q25u6ZUyJi01qUuUjFonegIB4AJ66FPX1HGhT7ZYiSAdpmww57jNxMH5p+
TFq1SlddGpAceCgiGLQLmPKoDvAWGdlVT6yiFTJQJsDiIownnBjI21TCkOK7fZaT
j4fyZst8tsyqaE5wTAvaMLuWjyYKGYHU/7e/+J5buGikL8MYZI6WquMfDn4ExGhJ
6/RANzGjKrXZD1eYOgVVDMlyLLJoRhOj0WcswB+ByAtR52liS4BUbqtEOSzSdviV
8nm0vKP4Mf9W3jCiUYIhIYubtjL94/0sR9pfdS3UlWJ3bt43Wr2yjNcF6ru3AXZk
CxWwcK4qlbsgobvkmkvNzgQ60l686FOLOizo3eSo3981xFkW5UWkggDa13hHWFvU
8/YDRQi4DBJObqORACXa3C4BNrPortaETdYLPsgkk+hR2JVwC2hCY5oC/hCilTHD
QaIhw09U44Sl6edVWKBHBNJwtHP5HZ731R4pdn8H4o9Zth0qsC1E4rqf+RHFrCCC
2llPKLHTtu6Spz0Hv+GZMQ1DqiClauJ+pKtHJ2Ho+7aa8ZsnyH79Dmf/wcpxeXoz
lQA8jjxTn4L4hY0jMZdz2YV/EXzRS5kN8SIpjyMEaCk76pfoy91PkpykfhoFyqUd
GAklPIcUpqJR9p1QQL/f6ODst6HtZBsTwHR1oyGhYzbccGj+cDg0u4hIXu8Kb2Ia
YypzMJ26sWYFXRu8x4a2XBLex9QXkILFglkq1tobiqboYEK0djrygbFDlwiEMp5V
+WkP7H/RxMm4pe67dOzY4dbo5PlDPY7L8UVYJnECt5l6fqIbHrObe0B1iA5nYp4W
7SSHi1ioCW792V8/oS4RxsebSPVaQnSdhh5lqZ4S7x+If+ZyaTMYiZ8SDSD8VvoB
qLzXWwZ+2tcf0QEJSro2h7VXwyrt8R4mqdhmPdK+buoFuGPvGR/yuYK/Xt5DeP1s
j0BBq+JfTKzkPxq4/QvLpsdsW69IkGkw2+Uyqkv7IsufG3VL56tl6jAEiTjMrfF5
7XWHq9y6NhJZTiNYTPDMpcD/dPT7Nq2h6TjjIgpJYtb+q9JiG3+uLaP9IYiggs4t
R+gxTwFX5PZGC3THzaqHemCdWHvUgWv1GyxJRKLwdTEVc+TQIHmadOXcinKQrJKo
A9mpBa/UJfG19ZwWanXrq+LJ9S1BKhvkYdORAI4uVFsr02Om/DO1HeoVOpHTqgc/
rrirEH8/LmII8kw6qEWtDg==
`protect end_protected
